`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
CqVA2OrUEw3rS2L7wrnupzM2b8ryA3Bu+lnJvxgVgrjNcEfookBm3yP7nJiadlfzz4GXwIp9iz2p
s3/zJCpagw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
PGdlKzNiAp+RfljaUz/4qWu4UrsaDdcb5I8m2pHEh9Dw5NlzkSTUrehmIwXHdNZusEIuykWSAGWZ
/B64COg99vwXbChOMVOzpixzv2mQr+HqmujYKEqSPvVqZcYkaJU+XC13dHTzB+nF8v5xP9lv8O4r
vnd1MJemao4IqJNNJS0=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
O9C7HpJnOAPQ7vXXyALA4SPMh/k2S46Hh5XdLMUYWYp17VipkHtaPGZ/6KFccH6RFn58ICZGO3KG
sGL5WYBNemFQqBq0y8svyUk+CP71thqm1XgysiiwK+cLbzasmWv6gd72IZaDJ0Dm/koqglZz9rGr
Yy1oI9Hp83u8w0ZrJCUozxT9sRuP6Hk4NriTgdm1bEZtEe/2gsoRGZ4uypGCTZ83caU77u5XkSG+
sY0WMUN4I9JDArAXRZlcZzwLEYJek3pwzASxa3Ss4SHc2/ugyBQEnz0u03Ct8/oB8h+AKz/WBsKk
FtYCRL0FkFN7NG6Rp1n4otCijlZmPDy0sb+V4Q==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
UYTymsFhvRnh93jsBmiwdgozSwCEH1PzuBioTnilEvHeHSSg1Ob7Oi1NUv6bQneX5bC/xEpsrKCF
ZzOktRibPyX+3Jk6BpXtTU3T5z4D8X9+eQTazzRLlGFkOR25EDBRMKSnXfl6zR1c91u9+kYZpCtD
tT41G9m2iVNn0qwHADM=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
EKb6oPxzLBvAKIrzC7UNBK8eY5ryi5iGJ7/BdocCXYMaivf2xcPKTIiYIkE0Hv8PshEsJ9YIK1VC
T6c/GEUGhuDsDpN8XNAiNGvxpcj+TImzhi0UBgHdiDVLhkJAtmhW7fOxixaqronVrRDaXAhWqA6z
eRM9XDYWonBS/l0El/PUUSoDAWcnU5LoHeBeSG8Z1TM+qyUa7w6WDqALs5O4HEYB8EIMehKvTcBS
pzbXxQ5k2wT+39vCq7Vncv5YubiSbq19B/yvttj/idZ0/y9fFAXYHF6USm2KGjPUs3+CmdnaA+hm
Q9TgqJDQ8e3agIUv19cQIAqFNQpoClnjhD3haQ==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
VT15/X4T4V3jrHxVnZkn6UrAuaA2quR8EdrkmUFjWmWdJf2TkcB/YHt56tVEUMbBtX0cu4OhICAV
5m4ThUbdpGUSaVYCFzK9V/BGPk159BTr9sJRQ450Co5g/TE3faaAIaUcLrZ3NPDqDbB8RYHXBpv4
SzpcX46ohjmLqHyCiSUO9tAg3SQcUm6kjbRntvPdE/PWVqx8jie33+EUwa1OD+KsIwM3co577bv/
C4E0EyQrjR6YYD7VCJNxl2h7GqVjE2qMqA0zrYZxk7F6DpgH8zWoSyd32pPOkBTg3YVuftBqGZWi
Vb6Jg33JUZNlOQqE0SjOJRpR8BExFJ8BGHwy0w==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5824)
`protect data_block
yJR42fHc5CAsXyeEoKbA5GovJpSKCtWqsx2WJOFLjdcR2YchvlSTX1QH6Hs8adhdRDi7cAP+WD33
mgXogbn4Ob+6oh6ZDzCYEL6NJI8MANxseD3T3GYyruIRMcP73cIi7ycSN0wSjmP5r/2dbl7scd6g
c5ywghWd3Zw0P+YeFzRPmtXs6NYFlZ9frnDHR+a1m0to6/KP8jsf67hbr+1Z0zdUN7BJlR9dQa+D
6WFynYsZuBRqECjGbUEm8pkhm40nTaZbuwxc3MsAczlaEstcQnTw6yaKvAprMFlxV954dn8NwI1S
Jyb4r9M8pmvXTbJsEMzXEJHtEVDIfZuy5MX4Zf2TK7EYoVF/VuNvJv8pVNnjdSv7UgT+BmmYLnsI
Bb+rHvYkMyus8qn53aYnWw26ngTj0iJcjsuA80xMxXpUH1+dU9A1jU4+oCSOQhmW35rhdz2fjZXe
oVu32o+co2okxofWcJESdgMLpZ1AP6+QMZm2fZRhhZP55pfK1P/Uk3UAWF3hzKQ2iJjJsiLGQTlD
LWSI1Ku4iBBLKwUbnqZht+hu9ul46nfDvJPnWlpO2jJOJKJzTDE3p/snKt4ZIgG4dXl0dRzB1f32
exPDK2ZDtlw3zl83Xl76D4ZCkBQyUvEtYPDf6dcPZ62Dg48oEKSomJUo4tVAspO8ft6d81j8M36w
ji7vr+R94CkW13L55d+Fm6gKkxTRpTeEii47E0A2SQbKzKzGvUEdtMnBk4B/U6PHMrrRmygUr68z
ZAM17/dsxIv1ZFsk0HDCk4jIqMM+DHIoAFEEAn6bw938JmpCJhXWTRBmKLCpVf2KFP1w19HtZ6gF
DKp7C49PiTtTTpF6Azux4VVKyzBDfVqREjkYya8W75o1qRA0kDsBrr9Pp3f9BB2A3rwqkgIiIY3G
k7ti1O/ds7/KKv/x4l5uU6X16jU+tpn5RvJuatsZgKTGkbMQ5eZedBaULY7U3p4h685ksDfhAG5B
5N1rtb4NnsFq3AAYBQbT7qQ5XfPZemZ9DnZjtiGRw6hXIeR5KEzKMTA/kTgnyCWZLq1vMBt9lDBt
YVgIFDU/sovgdvJhgfhnDgwO5xJgnI1T14BEWluhz2M4A9DIChKlj8BrRE6OqnJ3dcKmGs3YTIrW
NCM4VlDXdMeq43285pm5BlnGSaqP0YLK/S8wnF6mLnlk9Crgyujxuq2sFPcW4J79WSuURoKp8UfA
b/9UYJefknEntCgt4JQNSZqPIt5RzTX/BdVzL0kmhnlfKlPuJhEd02/IqnyjSwwfRTblk1yVD3kL
qO0PTJEm4lFDpOKxqTXWbIPRIw6rZBV9cwxF3fGfw+4s/MEMF6wHkS+XrVT7vKz9Zli0SUFTkvfv
cxfcGDvRWFSC0dXcppgiPyMm7gaNMyW5ZN0LSz+8CESZsjslgSdY8POJPjsR0UNcCIStuvqCzJBn
xaiEb+RgvNUKACEKKFxj4SUWuVkhBkPgxyXHc8aX7pXQiZVZY9A9Sib6hoIgz2RMG04GXfSCzIcA
f1i5t50JmrChcSTIoduprU27Do51mkVk7B0f04UxfOHYSo/TH5EfC9OH75PkeuL016u5xpCkqomV
h82N1TEYT7Yz7YnMKkubk+hPO3YS7ukGUO1NccBD5r03EvTWJIkAuqHWbGGLaX0D3w6EmmlkgEGG
QKNqttS+Pf/tQlO+rZdtL/VE4dS3OZUI6hqpeaLl21Ft7rHqiGbExIGCmiG9jI1/VJmpjmvIsESN
oe1EKSqx7h4XsBPWunJ0kLNeddWX2RUzT22JmUa5kYq+FTP68jAUrjOPVG6U12g6QGgiQGZ+/957
LAGD5xrFwtwQpZc49TQc7RiNQMyM+YniUlOSaZxouOg7Fvhy3vRXsYnWQLXFaUKZmTqbCT1tHdTc
ULN7u/x5Y5fk2dGFUHULmtb+W7r2mb1lv3hisSQ/1QrSbYl5SDexOdbSifKCLbdCbLr5Adkh3JZ5
uNA7DBzP4EhjhErrxg0gQPjPLBxlkyfuUfHELFf2vh51nspToO5QjqpsdFVt9DUIdeam4lzCyVuZ
0uF8VMrusSXuq20yCNDMtgrKTTfrDTs56ymPewOH0LkpArz1pcgxzaeWFI8kK9dyW6BCBiaUKXL8
BXh/CWu/5xNdgdsNhabSOhxR6F5AHpDb/E+uVFt4OP+OCl/iypLU81XG/fJjOuaurdfkqQvzYrOe
zEMv51DM2537+eubZTCikAb2juR3ZnoqyWiojOScuOjMznJ3GMQ+kXSyTyR9YS9B6rz8MC+Jtaxb
19pVNc4GMSOD10QWFNsoLdEj8MFYXO8Ypezr9i4A8++QXi4eJUcvflmq6mxteCh0DsClBjGJU29S
JgVY/p99ozih8Blr1aYBZDkUGwL4XBWXXzHfN23uQQOjPJjcB6Zs3a8FTms6TD5TPtEQNYlhE7ma
o/OwHWGb1sfskK/Mi8gZWzpIQ4Lkq7c5b0I0PoR6HggbQ+K1/6Ocu5WsoWUNdfeZrjUwjqiyckvo
hnxtI2ncym40dlCZnLB2zzjfv3GjoEDBRxzL3wlwvnFOIVhbqnfQXqN7lXvXrsfFdB/+Ov7b30LW
JQgWdQ3+zpYQx0Lj8y3tqzM4tjvnwgTLBQXhVN7WP1R81OE4q7P/8HMhI/8BBMNqh4nGHHW2619B
JGidbjo1YUXI4drZcQsXTXh5KLauFFYs1X4j8Nk8EhNQ4SI9QeGoM5yOIiyZyyLsYLm5KOtShL28
m9gHOie6EJQ2zCL1ukVyGvlDe/GR3v2dTnoIc/2lugnvIn7jiIDd8xcjggW25paXac5CSjr4dxSm
PCVUGZlTbTaz6ZhUVFvIogFYGFyDQ8iCk1bEZY7n+yB5zSRpemmamX5+G3o7Xai4KW7my2D5C8+Y
Wgvy444ODPJyZcqPpAs5+9AzWu9Hu8Z9mXnHi2gAKBwalGouAWytKR1CFa2C0lPtfHhX63st5ZMi
/tiJU9EO1ZVA4eaEJ+yueC5E9dWDE89A6bMYmWjb4u2Lb7mHs/eiTYhP3zB3uz0nSnQRxZIrVFFm
dwaatPM1tyrdAOal4Mq3QTbxdPhyyBIMxhVBrVzvQM4tWj0MtiGJ72spBZQJFDokoaalut4ZLp0I
2TfkQiMW0z4LBo3J7VpTugMdD6W2iEFwc3/MdS3Rn+wNf9+Bp4wOxr7n2BLEMj0F081fufvcH2W5
i3mrFlFSUOq+RSdO4cFCoDiIyi7k1ZLQvCtsQr9SXjEAvBZnhEJVX09fDBrW4MSktDwP9svNObpV
kjkEjfvwvyCt9+FyLeBLuLWY9izaOAkkacz7lAtGY0TOJCS/ywHIkTDjIeTAe/crXBoSn1xMwRIY
6MOlFHettkQXrbmXh5fl5Pvk8WzpOyU35vua3U0iQOASkf1E1aRLt5eY1BBM2GQ8TzNMX7khBvp9
m7QqBqKTGZ5MaxfFeXos9/OXWJGuix0UwsYQTDC2LLejCIVeEMiSkJtwvCC5Z48ttOmAq0Jl060h
HqRAiesfoR7PiPRVqGgVjrehHJYlJqk1wWRQlcWy9ns8uAhS32WHWWAmfmdupPpSqzE6k7Irf0Z2
rj9A9X/XfgeR30c4OOneAqmGBAy4xhlU4ihgvmg/cfZlcP19IyHpt5cjvhv7/5ZejZOBkOMcVdOV
ChbLH/qTEbrg7Z89QiB1Kwg9fzPnNr9ocbKgqVnxbsXVCQiK8QQ730OESphG8zdENYdR+lkZY2U0
n47Z75c4l+4yVpkNE7Pmnp7TX0/79WqdjTWCRtoG5KNlxNDwTEHDKA/TNtTw7zpfzlL9puxYyoa/
l90scwydu2r2xUuiH4gFvXyItCdznbDb5jkPF/h2e96WUYqqnSHWr7hHijYgGpiz/D4Yu2hDz1sf
c0WmcEfOwgRWtNhINVRxrUlzHA9i353+kozqRiPgcZGAefBqov61ZBI49PAF9mTwZQKVgOrQTLX7
/XoH7XgageTR5aqtP9iCxjWmrmOztzKBKKmDeJgud3IoXKRXmIKPP8FVLO8bHiSzQ2K9QuErDj+A
7YrxQURPcjxVkDP+te1/1Wu2EtlVKf35xufVzPYbzskP2AkHrAORG0n3RWWoie8ihYX8UYXhbj5T
jITJRzShBWqU3GxZ3PYL99Jq9fKokPWSuABAFt6wsVkQzGHrAdeCuO00Oqlkpi9fDSgt1aTDEV46
n3g1E2f6eQiUa3AAZ//4G18m22vErl2c3aa7wnQopM+B3jrW8Q10yYVTJAfZ4HcWB8qjC18VH3/H
DFmCRsA+MywdoaLRD1l0Jdl960AfLZdOD+MN3XXBh8aJ9Xm4Pu2CV96XYicBc5T+bPGDJWURsVfF
7VEFTZQz+ZBsL8tnlYLKyrlZs3rzGEfcC0oCawOdxJJjgos4D0GkcTz1ygtYXtSFVo8pM5a9dqVX
6a+hKQS8/xD+ok5hLuN/3MJj//Ba9rL/p/j++Sk2ieHLc0x2d3f/j7Jkq3DH1QWSoiVs/mMrwTfX
k6Cb3aTAjSdZOvl9SXQ9ZQQ8dB7ryjtOns46/oTN25V9j/ztuLUgiu+Hninj1LZm/rCPJ4B6/l+0
4W3KNSEWOoa5ojxrHjZTc7tmgwEZAHYy7KNfLMGilvdARQNIX0UEYnvVYnAyrIh8cO3VKupDUJXx
UVdRze20kWVpvu9w3JIjyLKefDo7PigZ1SnEn/sNiKkXDayJSGJ8P1hPsJ+2lxedJqmRznIXum7j
Dwh74ZDEJ2+V+TFrhTZ8tzmruZbj3bY1YoBbd+Cx5QMH9GEs9acv4vIFkzY/8odQr8iiG2XJjXar
hS3+hZzQ97y1sJ+QzIL6GuaUzkf8hyQ9gHLMzm6fzKooXfzhnkqirk5CCefF4NbSIg7JOTR+PKR6
jYeAWQdl7vlQ0hJr9qCItMLoQOXX78+MTRRKQ4JY+PrHBALKPbVw7EBnYWlVmNtBpJbC1T7AITvB
AbBgfWcN6/lO3Zk4ROJryX256mN+mvrAq+cp2vwP0X1txs0gWKKUMNmdZIlS9w6BxK4fTaU4sWqG
SqddzSzJiQtiZwewIxjlVQSB/L8FI4FzaRpK1WOPe7cSCid5W6DPlJYLalzIXG/VoLYBTt+ySW8o
OYhiVrX15gNc01c5thw41SgZYjWMfz0qXTFrEKXKap24syOPwSbGQvRJPFyAy5rYkPLsBWtUiG1d
FTlbH5Fg0R/4/MTZKI0JbCj6baV4gFmSRCO8IE11amwD5wdGqAb7SplByfOtxG/b00+BTJLsw8Iu
mYQO76G8qJmbzq3+mcngSmIvLeaWALDnb8aosuLWXTSbHC6EqgtsDX/gwl5Adk3q2fS92JZ0bhT+
M+6X56O6KreSJ5QMIjRKDKvI/kOVjgxVD2nJjdhwcv83W99lASaU+B2kxtccDslHB6BMLJijvrTj
fSjoRghd97OVGeJEQr6h+PxcMasRXkfjVp2oK9Gdae5ajwJUTu0DcDEZF+imErMyczMlCkoERkpw
k3DacmCfmN7yH83/5QO+7pZbFVJCHQ+pGlTKvV7yXEe/7qj5yXPULK48XS3XM3nOiqRygKTYP1Hq
IEo9X5zTOeUNHONo6KZcXrFrXof9Xcn2swmaYPm9u3kB6ySleg880keK2ojgTmfMwpkjIW43WUFM
CWNTP7D7bfe7M6O5QO8t+HGCJKyHq/TbgSOmczUZiZdUa0VqenHnwEEN+p40zvRmIK82mn2+wT3U
9bVi4qGG79YwK5d10rq7p4ZmMvoXj1JeYfYJmRp63p0/LjhAeqMfMOpQv+O8Ne9v1qU2OyGHsN8V
03AM7yIAQ1E4JdhEoCmV4Zzgp7Xy7hR971xFc4ihPJGPbHX6sAi9r/oMfg7M6IJL3WCKZzhw3Yg0
aqEey4Ul5ObEWFlbb7Hw9JGN1GmQf1swqP3a4kV2fZzpSHwRcupI71tPdGhhYHXX4ISkD1f+Gj3I
46MGsFDkTTEa0PLGCS60vBCy95sNIzTI+LpSuIVyPgO2HrZBa3tCCVlsfO2XmpvSAy6+/09bVswZ
kKyHTXrZcH+OQ43aA9Oqf0C+yMPDyxwS/VKw+sIz/a+j74mvmZDfrI0WyIfgS8qAHgoTQmKipXOD
AdHc6heQlGvz18wFqCkPeSUp5qxA9gODZxLOm6kWN0m/C9bC24bXsGjFZ+G/XjzF6vfF4Mci6PUV
6sRJ0j/sQrpiUR98Ca/b80Fpn68NbPONfCRPdfkl6+EAOPTlCcMN5uYO+3JZuaoAjGofL0I2XDjC
eQaVM1xdeMXqc62UPD9PEYP6IbDLcOZFGkYhP+1hzqHSG+sX129TjgXGNagPkoRQMPebXUO6sUp0
p0RUttmS2JCq3m6f/YBVHUtkUFvAOUzz0abM+5F9nYtihrjQrvC4vV35plaJq4CpS57E0EOsxTG1
bC4mRZ/qN/KX15I6MgTQMIav9jCeHf9+pC8xfz1pZBy5xt5uZixwQnI8Vc9hqjfrI+M4WRxzXkIm
LTiV8f7O3HWkeNDYofbruD+uNEa/GRSi6NVJJm901sNz/V0B9SWo3Huc112CmPErYBmNA6AS8nxl
+HobpUATsjdHgtccSHcGhjNdNWF2XUe/lLdEi9WD18fJIWYejwj7R7uR9nIKmi3FqyhXr2cmmsBI
KOuhS23/+gDmi/eB5JZsHGjeHds5emdr68WDRc6wTBCAJU+pQy3loIY/bEA2i/fxHwG9+5KS+wug
YEDEKgekzvGWdZCXgLQ4yE0kgdRF3RqPxhAt5kQ+RpQaKJbgOsY5Qy4F0H1Rfdzm1oEn66HcfsBq
RFhxvgs1Cip/tiYA/Op3ISoPjn/xI6zChB9Eu1AiPIJnffzxpDj6368Dk4k7k0DJdaoRGfvkxg7B
W/XfaQxU0O1bjCwWewL2FSQ8LpXnAJ7t6BcCwZnv2di2qT8CE3ps9fDwB3KaKKTm9VPWKRmSG9v9
feiRZL4MBHl67v4gbtyWMrnBZwTeD44m16oMwYLcsPklN7Uns4doYCFS4PWaSf345cckHaXpjnJR
0Pp5Ip96QR0vko02AkyDXSeh91rtfQnNZVqcxoLolpaUp0FYUcxQ+iBgjk7HWW9Gsgx7Qegnxdn2
yO8H0YuGkYo9ZzOUlc3JlEn07nyRCgnh2Ll2LyoLXWpDjgi6FRTPDQRCGUWVTRmYTvW3xsIZm0k7
VVDc2UimeLX8OGVkkj10XVQI0erwMpQRJJql+GhUzB0U6bY9NU/ChaPrejUU6+tehHGjwhzung0i
5LSTGqyZJzaOEciIqeLYZRxfbsMNZ1qZk+xCMW4EVHB/qaJnys7oUx4iWn0KhmhE7CZzpi7p2a0I
c8lhJ6ONJEt6ackGrsCTHyJF8Y7iB76RcRmj7zR4BV4ac+RyGLU6Usbb+KJe7YwIMwH1DDcyc+k6
BHiO9Tor/phI0As9woblcPWhyj9VkoXPCAJyX5yLTcBL5ALm25t9s+TMJC0+s55cVYu6mm+0uedm
bS3r/5lxwgxlQXXtgYMNOutuYWCGM7GEd6GhCD3ldk6vjp4OxaHLCq8FSWredp1EPyY02R+IolMp
J3C3F3GdpuS9F2ji1hblG53OInHOLbbb6pHjH7c0aahMtDUzT6vcAsdVhiLqRE4hshJrVZ+s7ooA
3+wePYWIAlKLebsvuZtVwJbTe3dRIbWaumXeg2I+C68+OzGp/r0EepBUZNXh6Xc9AOqUcm0LHyul
Nb9v+WFclHz8WC8WBrUnsu4cQqiMdgtoIsCoNqYclX9IcVneLb4+A3trQgewA81+5bG0w7wjlfLi
/VWsFmwEPIaZiw==
`protect end_protected
