`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
K6MLXsHy1mE/e+BDKQWWCf+4ivx+zNnJ8O6cBeb3pUw6btsYq6X7MtHOz2Oz8HDGPA6q9x8lkpvp
HcdJOMY+HA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
P6xTgR8Sldnm8Q2SDl0KldP8Mxalhk+FQ8DKI5wS3in+vTjwT+0Qnq+F+NLFFYSjCVLQsvICID2y
uDTWUrzC2hBYfXhSogTyPkvWjKOEUhadOtQFmXVRiaRRmDsmYIP0VfzBDciE/+KgDZ8IlUPPc2cU
WqlOcJ/eLogYE6zQYMI=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
QdKj0eSWfm5SMookhXL5Mfkv6ZPZaxlVqSnBQx6Zt0SW9kTejDuRAfDQp4EiCm9dC8Y0Q5g8DAto
xJWkPZTunorz0KoMjqzfZLgIPVA5PGWbf1yF86jDL7ftFfK1/8E+/7kecMymdPwvYYkrdFLOrl83
j0kjqGJFjwWrjZ8CVV09XjFElDr4v/W+DOpUjCphuOH5LKetNJs0j1z+JTO6XyruGaCJzAbl5xfA
R3li4pGfWu8XeN8gITkQImYGrrJF42U+3XtYru5NbH2wQlg+/uqFprJWP947IwURkztN7oj5DsqW
VGP0FCt12yKYCT2AceNJcCSCSfsK4Pc0HB0raw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
mPUaOpmvmhBtVYCiUSfFBnEWc/b/39RU8W3MPTyFNUhf8hLULjpBea+PhKmrbx+gPsC6jLfNd/Xy
itAaLl+gJoHCpcTd0fHd0QVx5zBysFQ96p8lvwTAzlgiIf3KJfmwt8iSojdq84xPq65iSh5WwHu/
tEAPVBe9eTqEsegw5OQ=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
jrmiVyp7fll8pzeg0coNDePx3gVSGIxJxJB6Bfv2T7tlCbnb88FAvJzHLMoMUWGpWm5r2zw8eCKa
Re0+GzIsqFVL4pR1zaSSapK4xk4ypME+FriinPALL2yVdhs/1J+jPO4gjFoISVOsvns5g2dSuY3P
GJVpKqvQHiraQr52fdpU9xAyUKpykZT8l/DaSAGnjzaVdxVj+HEfd2wVvaJm2IxmKgnNA1zzVFzv
P08LRfOwoyCo4MCVekMYpFXSZriE/BwYHLhQ0uJrHSez7UD9w9riANFGHIoCRiRg998RhA8HIHyB
SviozKjzIIihOUGyb/M6tsh5Yc/fya86iklPYQ==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
KLs19GN1d72xAG6XSs7/+R2FVv4B0ae56gDUM2+UPaYIMAruFbPejUIaZmGcPW74627oECmrLsqv
yMhGuqy2Y0ZAH3mvlDb2l/KsIFLZJZNfnjHfIqdh2ln71HiLa9iLYqMfDqFpjbsNmlibkeIK6Ye1
6tjFbBzcYUfGzxxN86GVKIyqUC32+XUgV9CY07BtadF/xu9ANU8romdQ3zqjalL6iPbVHMGpO+ri
zswv6sMOd1tX74Na1ibUuhZG1Pyqcpbo+mRkfRQN/QptsqOS9K+PrfdE7Vhte7nW2/xYzDgGdjP0
IIGZJzDtIH+iqkAC+Hw6/elB7pBRqkRDetaGzA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1658064)
`protect data_block
m32k8HPm27Xy1sF3XgmUlhhdaxULN0v3NgSTxzON+3Z2mASsM4BptcgjLMnB5DQ88KbAh8F7Yafu
+YhW91jC7WTZf+DScWwFcR4dc85nCfeK77QuMp5btNH2/ZOzYXKYLBcFRh98o7+UDA8Gd4uXc1DD
NVjJzk3Y3WnRWUgA0HcroV35L5CtIVrxBOITIqOxwiJaqn6QpVbj90Mh5HUx2MYQmHemwLRWqINZ
1ygnpjummT9ak4WcJ/ihKPW/Yk/hX2kFC0E+jpPLJ4pGlHyO5KKSc4DnjEEW//hDsz8C+XxAeBA9
yZyl9UMji64VFpR/PQ/V8zZ/VmfIziP7IAPtigZc9ADvG1ZZ4rpaKK6R7BeOcEfXYYVaRh+sDXNt
/q6XWccAlM6VHsy6F+OGIGlEPvtdHkm+IKeiyh6e+F9tc406hVOA4u/4tHmmma2VUdCHCcl/T0ch
hW/rhKbarAXSNr4EfvBOVQwnGnq21gO1OxNKB/odM6DUk+Vc86RnVXeQR7owYKKLkk+QBMJaaQM9
3yXDg1oCzLqc9o/uS0WRKxPrDd/CvrWioA4BClkkBPXQNEX61KWYd08abDCSiUJbaAUxxa1JGqPs
BRx0F6LQtBnSZdopFIhl6aBxz0/zVEunEDQXdQP5zYBnTWGCK4X3XFYasR7EQXhMhQLizsbqKwGX
NMOW+sJ5cXYhMVlx7wuFKoCJUqPDm4C9QfuIoBRZGvDPJQzqsbwC0BcNfB14acwqT/vSXXZf+zDe
36uSoD29y6nlV2btY03j06Cye8NacFwZ7Vyl6izcvB9xcS9yzBGLA08OIXskV+Lc8QYJCa38SyZ5
IySFizxGZLuivM3cKbc1XanMH4c6+vl7R716ySsHIPkStDeqrVrnggCw97ecYalgakxcWaxJzhD3
pQFebis63xkqNj175DDhGflCZ+xmjI2uwPsif5fg1DBcALb8pv2las4cOA5OwKsX4BuY5iSVyuDm
Gn1gQGpq9mnZJOom6EcpJ+7S5ZCRAvi8lk9rkQQGD3m+F5fczpu59NuStUSxjfjKvfdyuXxipTkd
SLpXAnqkthcXJ1SfxyyInf0luzIG8RmocWJ85z0rWswbJSUe/tVIwAoEe/0VCp6dpC4KShfV2xIA
SIhWVpjdPxRAmqfql5X2DU3Jj6YSOMR9uHI7c3xdvqjSo6k1QJ0QJiOF71+GvjNPHQTkY4H1tYnQ
9Rtge11bByvapJ1UgWGn199u0Vl3uuJeC3/dfhTdmi2oPo93y4WkG13bdhE5pfxarYdKwiO8IKR3
mQdYsFh519XpHvy6IxSRqzdBsmSTl5mGfP0m0DdEvGtmmDWHeV7uMOpfX87HADJdPY1yqwsmhq2M
pYdjZnn3aLVYqbffv2GrYx46Au0AIU6oXHchw3YIpb19zmO+b8T7MYyMPvT1qPmj7HuoG8HUpYSh
37feP24Y6ZKoAjtleOUlFrZLfwip5DiEq/x9wMSXvbc4PoNGFeudmqEjJYTK7Jgyv4p7/2vPuWOR
8TUYwoiDeVH7ZNBuufR5rUACGCZYC2wZHE1S5Ks7DJVvV/4YUr7tKp8uQvkngTRKKvJYR/GX/YpE
SUdhYtU4gOi+iLFov/L2mBbhWPqXB8rMa47EpN7eSPXm3Z7z/+LltNIO1xq+Dt6Xn61uouahEtiW
xv+idnmfConFKDtlBwb6eP/bPgWKsE4L6ossUJbjx05POYE6Heltch6LABtkquyVQEagA4riQXQZ
EzMgrr9Ty4WxyjUnGjG+FCCx4K17HxSLEZoGJGVbGdCGSDTkO3TrJXaWpR4sTo+c2v8RPO5W7D/B
MoP3Os8GTO7KobuFkLyFRoZTdt5x49+kuRKMfSv9rqPDY9eu/floEcd4IhB52w5eDgyh5fhJulji
vxH+Fm54MRntOExZ1XJczxjfEi9hV367vaaQHyfT2mMf+PRGkYlOuHYOSAWNoxz4Bd0fwBF8MaU1
wUBVDHI8MsTJBGyu0ibfCkI9xVlh/IFZKyXP08SOmPuMM0x6aI804Z3Roqj2+bt9ZgfvmdTHl0UC
fgZT+xtHh5uHfp81pqPts+gHR1ixVmn1WalqBCt9V7pk9SIbRp/gbS3RMQFP+PwbVPxifF3XxN70
we9KQ6z41VMXLWXZE8QGuZWVd+63GhL2ZpP+6uzo1gtLimQQbxHzVW29U2OaU5ARSdFt8t+lTHXo
d+0kNroiTbqTaBncaMGebcdP8cVASyi+TzR+XN7gMHZ0HgS4TBtHG+PBk12zAlsKuhThxAXlBoMY
P/Gcf/ca42m2Rlgc36cZC1wtsQlUB1avo7DpD/e39I+bprXHS1GuUsZmX7m4yjEe9Ium+5/YfXbX
Re+RelJlbGOTNEvkVf4YVjAQl4J59LAwUhm3eIj55tLdvTeXdrxHtGWiTStaz1zdnZ1tKfi6SOvi
s6ocpy2VlvykpjvbFCoSGvlVSyLGBh16zlGOdmDJ4QDgjUrK0TbTLSVrNOAJzaisLTwkpER0kfiF
l51CPaEddyOI7SruN6Yj8jfomtP9qm67tcd4G/fh2+bM4dFWM1D4tj1HyQfSr5HGO0mBrVqw/1mK
ig7uND5xxk/HrakQwDNVIj/wbSIIcTQK+uUGVzoDhx/rsxabzjudMz1K26rH3oiuoWwBLtNQ2ILL
enTY+0kyzrTuXfYylpXJzUNF8L4IqMYyrcV5CZKPoWYQzEN2Yu7JM/PhcodTml2+jXxKpYIn6Qwt
X1C/V1OZCu/Zmxan/oVzeWIxOkKMvwzC9sCmDyi0dcO7SKKRh75cVIKDUnuRLWdI46S3TEaQOXsU
8bR8c+ZPP0/S8y8HP8JLcp+CHPNGvxDaaDvtiADMk5MUicMwcj/RAryfGCtFEVbimIpcGAokSaM5
oOTBp+SBHd6a16CxTyVvUHTn/Xi7RkKJLJgubPCE87T8/o/vSOvQJJVkc0XUf/x9P9H4Y/iQEj7G
2G/51qMjjqRaMex1n1xPOHGWLbhyfYifWjoBtY5H7Y9l06CFJc+ItbIU0GevjlJpjn8GPpKcBHVA
Ut3Ue/uR2DoTh8VICnN0ojBvi+WUjAgH4Ri+0bDSyZqRshwbqfxo5zl8M0lOEY2GWVYnI+M6Aj4z
J5zcYpTnQmAlMx2S+lAG1PtafbPRZZ3+FUAXBS9eEvclqO6OMV2Jvk+EnAzhMQQhjyAExBTXUpO0
pBfpo/t97nDOMnPorHXqrWnIKTUZ1/8CJBFUYy2/hu3l3gVvuQD22z6XoWzIvPXSczk8T+i+i2aZ
Mm8aQOj1LPFjf8mq+jwoapcF+jRiHcmIHtcD218e/KA6zUjVlhiqYoFW737B7XxSJNQZKlPcABpO
S+olnKPR2PAIOHKDgbrvP/JS6KYEO9j99HC8shXEQxc9YooMT5fVRpPfrNwGR+dFDKs/f+CuMz2R
Awv+v9J4lOL0ZG9ZYWVyW+bDRecaxwHHLlZ5JCysBb1Xd28bbp69jHcOfvgZVclgZoxcsDxFO2JD
jAPkq+n96oGo6rLYx5nXtHPAKCauvSJC203Jkg5RwlBc4Q7c75xCKNjoi4mENXmqYBvF4PEL1+Qr
l5bW4RroU6cI4drhNwMpcT8AdaA5MKZPHtFkzNv0EhVdP4oWv/Ozix/d6fHw2uvvCouAMZFPmduZ
6L3vQSmyLo6DwOsZPpdR7YEMF049ZeAaE2GaKoLpc7zYe1HdAzDfRneuzljGChvpreD5a2IB1f64
vMNcZgwV0ikEn33tn5LUf7iBUDgPodnn83WtqUjNTa6g6oFXcLHhegJzgXYBj3ABCHBLofidjuwX
ALX54dCrJV9S4ZDCbKnaikZW3Q7CLelFikycgqP7PwPWdS6Y8/IeuF5iJZot+ebMhhYIniX+yFas
dntdKuLTZhhDafNh2UKBkZWQZNN/n5O7GqUd4SifpcsvUQG1q5o7guUFRCYDgtJeeJgEJiDEHNoZ
cA8LxYlZ2sD+awcTCYuKM4AloQMW2k1cm/Ri0s/7uWf54q9QaZRDwCve3sZw09O0+SLxFUwfhk8n
q9Sy0d8A6y3FKt5yPa5/EwPuVkQ1W/lomj/w6eMjBf3T+qC3fPhw+GdThnVhaflWDCFt4nR5f4Bx
yeEKamd+RIt1alfUjINMMSJRHjzT5FySay9nutAXeErQN9vh0WrziwZD5/39/C9xaX3kEdRBue+X
oFRpR260GPXvggUqNRSMBzsrz2sWxnSSrxc159GatL/I7DFf4QQ/EQuxEPNq4euqMLMgXWUhNtLE
4kTQMeRSAu9JCgzYcm0nmPKzCnGLWYxjC88xURXk8ABN2J4yx7t5lKsKVxQdXI0Yo66amelc94An
M+PBSgmVsNK2HyaZ9hVftdbvhV1tjzKtIrBLEKqjZNuTM5rV5XgSyL2bH+IMIyap7AYuo+qtEi5W
Eaz+TpA5TOti7eVMxvmNpoezS4kFR0yc0ZHirK3zleoDbrATQiDJ9kSCZoA0XO6rAMsypmbyL/k8
ltyry+eLiQ+iJRAcNoNqKKuVbRM2q+ZXep3vUHu4Z5KV/GQql8k9teKnp/MwFnU7Y8BwAvQBlzfN
t92Z77pV+JGKIlEruPSNbUCqGV7yzuk328ExUZ9MqRgXh3/o2L6P7yA7J2p6ZT7w5WR2Af3ONhg4
JJV6Wkbq+TgWbgnFENQ2v5Vi2SjsnNSn4CVtSq5fofjRBWArjfljuKHRRyHzuJ5ZULhyRMUufCbK
s4KeWJ0ilW+eDUuT3q1sdPAQO7OjY7eJANmZo1ED//H89RcOqcsANJ2Gww/np+fcb39vPWmMjL41
e+RK1Cnnu4Y1yPR7zms7U9PX9rFodnAvWn/M/mkwqI5VpO1uKbZ0YljyKHLKSxUQQ1DZJN5Xa5Sy
XklBrYV87sVFvIFV48jC8KZrqZdmAADAFcuEh2xlTAfC5QvxiKvJ4sPnoGN4jvu7WmHuyPUcXwR4
gmZq7Fm6Ycm18DFUITqDzGnit0Mi9+0tkCljznLJ8B2PkFs5MRDsOIplRrlVgtr6DzpmPbbzMFlu
ep5qhd6TVdFBV8jPjoVazdtylERLOUx7F1FDk6T8RTSzOhfVwYeV8cUtpPuGdIPo/qZ562Qj67/7
8kQK9lybXOYs9CPQQzNuloo62XkdG+SSbllHq2m5zVwsUMgAEyyU9uwlWvjJaQH5xvUd9cvScBL8
oFBYx8BUTAMoEzIZNK55WyiLfpSh6r4garq6ZtmpnqpkNkovL6rNDZSWpukY0lXd72GuCj4AwUTw
PmqJd7p+bsc1HNQkwDLViLUUeGpOzFBkD36ujpxxANUxTSPISBluVcH10wkyHInNoE2+ntVH6tZg
ocN/QIeHC88Apqa/ZLmIkTx5LCYndLIl23AaFAuhN38k9f8zhbz1Y8/tF0rpy2qQD71ef6jW2kpz
Z7ASirJJeCgvQMo6WE0EJD2sFUCheci1bd1qrcSIUrxLSUhOqCmc83RM+WZShQQG+nsPvMp1Bimf
3KsnXcmyI4NzWLtacvsV1lPCx66Va9wByGYmgp+hHWkKMdTDn3VNax//JP0KIiw6fW2EyMB4hEuY
Zd/EMqtRYlp0ZRvRb3qCKsS/3jWud7girHnUB55EFV9UDD6edvUnIM0JOqyCGETehTXhNYqxK2Z8
6+s5DM0s+9eS/2K9JlOIlqmcIRnu7NkvLqq7W+tehMLd5yG4IBzqiyySI48KvVhbeSK7QoN/4MgS
n7QRPx+ZzSJFAtOIlMcN62BStGLph5VtuWdw4/4rvRX2dw2SYxqr3f8p3fa1rYCQqTQVaFHYK1xK
XrXtDGFUnVDPwEnJDg/OQO9g7tQvNx33qlZ6D7uTFcZlMK08mMQe6fSaS5avzJpsrDnATFZsTRVX
4NSRVSnZesObydyWb844O+dSAnGqQUiCV+RTayTiTEprALYu7U8RMcEarCT5ZFbJvA5kmglqOccf
ZCezyaEjjHZ3vwR4VoszrKBjVoKmxVas2FWo1umzZT4lUiEMa/DIKzju0WhewA/WmUO/2XuskZk0
KoEnr+Nz1uc3z+BbWc8aHFZKF/rIiRF6bErKFNrbjNPV8tdUwEJdRj1OOSJ+v+ZGZcSfe8xEM/9n
UjKAvX1ZSYWzvOCu4bGKpV7ZDVtblY5RjyN0DBWJzdzcBYOe4bjJ1mBeJvM/pTCSiwFcXzWblEDi
WDk3V8wzW4d8FXJOk/CUlBavu906VOTvbqbpDrvxBn9DN4W04J9kSiQ90mW7pio4mfRuAchphwkb
fJPYAOziWenImGznH3/6J+qbTGMeOP8lkgdWRlLVeuaSXqvyYagA6+vtv4ceS92gbakj9QtSr0F5
EMuAoM0cMWWY01mu+cyYdCwT24H0k+fZWe7LqDHPgOs8JIuJvyaWERZGeBllYCXJPQs1gDcTdJOk
QpsiKYb4S1Uti+7ChTHEuQFWcy7n7RzzZFWqw01DMus8iYPx3/UnTTOlw3B3bgyy/rpm2pD7+ESx
tUZGPXUArFZFF1gbGdlWLeX9Oc6AboUdWJnKNiFykaW5hrKZbsm2z4GWZIJLzQoa09zC0dZMFTk2
DvG/RPXYRoe8td/YvtSFKQk+3ULP8vP4laXfbtvCqXiwByvrRtbelfOF1/lNfnpUGFki6xr58Tmx
IjggIK02dflhpc0640721lsPzFF/gTiycHf6EgJzrjqEV8qderRl7RuOTG8j37bl7paZI1E3rdOg
Xw9+N66nfv5zN6IdW6vKzs5hCCV3MxY6Kq9D1NP95yZmwAyeuxYjl+9ZlMTMDzTVajc58vNmY6SS
8lYPLxE7Kn1xOLY0lPKZZsGyOJDQKdize6YGqe7nNiegzozBu+HkdNs3pxuJZS8McjcgKq3xLybR
qxoAzxxeX5NRV3zrPyakR5ReSkEfAAXSZbyqZmrw5FT3VDMPjzJjJEaQslrwjPxNCEFEnOo+Qi6w
pNiXCrXs7FI+Q/TPEzXkSD66Q8J6QMvU2n8L90jD1vkmPeRpfzGTjV0MQ5Zqr7+bJJ4MsTVd8G2q
3J+to04B/xd7TWAbRuaHWWYaruvJXksc2BZ/svqPtlOVNimX36CHtY/cdGNDaYuc76iFvCFFENr/
pHXWlWv0EdevGJhvcokDkjit6+DDdwSox6q0V4o6MnjOGkqinJlfjUYfWwjujaokbxEMAEfwGuwN
ErdMKqiaRM8u2Sj3hKttFBYEptiTbhgbuwdUMR7nLsol7rbE8mk0YMEE5muPvaTU2D15Zs2izm/Q
4pdZ/kEOlEnN0cKz/DY8yqPi39SstMKQ+ID6fqtvPHlUdtwaquCGd8Kpa9iXhFzlvAiWFfB5c4vH
mseZXNLhee0RERDALhUPMVAoE9NtH4zlgcm11/juSTMychhMP3UapzHo7Jbu4vZuXwjqzk7WVU7R
OdjBCpsQlGQ4dbzoKh2vHgMkz3GkAiKPo8+q6OZJyoWyvmgjnWAYx2xWrkTLwRYZwa2aJnINVH6c
OkZ0KN6b2uVXpd4C9ssW0b4wUTlvOk1PFiSz16xyksWuXbEF9G5GtYDb6KMD/PyfpCZuvIP3pWTd
+Ot8kppZR58LZFTTueCkSBAHdLXVFkWLhW23L6NrFFOSR3X2yLES/6wQjXDIWVee5EehyMCdrwwB
mMunN8gqqjCSG3TDLoWaNJk4n9/+kSGsFBMb+Itqyoowtqaf775w8smHaKoEEqjRBYAvX/kQJNG8
3nfO39NDM9xEbop4hyYCqSfSAkEJ7URfsHAwlES7usW/cgVARuVvRnNz6jw2Ehdo4NHRASPJDGEw
oKOgfUjIDglhv6DmgZ848Qvy4VXF+kdQHBH5+mnmjT8JL3vNApuwlk6rfarWeq4GqvRcnlpYusJ6
68R62Vfgdp+ujNLINop5VmXywzeaOEtXFqg8sQfA4KZqABe9bJ1htfEyuviX6PY+aXUxhxE7lZMQ
SGJU2fREeBvyL22b8UMO46ThhtJU3AbxcU+MxbwjTXtJ/mzKTlXKMl7ps5+F6FJdY0ARK4KGCfU9
X2t0yVdStm7Cn+m7F/IzOvTDssJnjmZMKTJzZYvAGM279zCtK5YB4THbrjlPSvoeQ8qXmQaq/yMJ
TsN0KArZH7ujjDV9Bhchy81W6wZ1ypauUUXxnFhB/WoB7IK0ADRBz3ZuM/ZaMMfaiu6Wcffd3FaP
1CJs/okGszbJAa7CyiI3gAY8kQW+65lRlGaJ4odi8EylTdG49qt8SzyOIcJOGkQiPYK2J0XW1OIn
g35c+u/DMjXtXKhYdDiKkcQR6KxJLZvr1w/vaUtv3WUE3zx2S41wEmwjAGcO3NoaIzAU38DXAUt1
RJrOimi6fkZQGvBk5esko80wKJoz0+D/8M+Kp+zfX0SyiCuCTh5cw1tLpS4PebjwNQBtpwmsoMlA
UpcYoPgaPvvrmCJ/weFxvIe3XJkIwX0YtyM4ZeCrTbzmabkQPEFG/S/g0LjdmuFCT08PcfJ52PsA
djLLPcVYnKy00YVoBZjNcdQbD00xff5XUDHoUNpCL+5i6SKNR8Ju0UkuwOfyUVwQjzYcOpDninxF
jE/iGgADM75c+gVvV0ND32wq5ehCg7/k9tT0s80+yQbdjdSZ6NMjaZGgM7GtD/Xw2IB8tCyXrdz+
A6+0YfKLrXcvLm+Dpe/tSyGfPO4+O+FQH9jTFDtxXg/cWv0S1r3LJDXZYVVqKV527WGV+kR8RPPs
urCqwAMh76QPTXCnc+D+SUtbJZVVsVYz8I7j5ZYAfpcY+Pk1AoNTsI7cwvgyHvh782dvkg1PN5Wg
CoW8tCDsl5Ih4fPubEI74cZdTSelcdeOeafh1UocgI50QCF3oQyXazE+O9bM/1E1ZtkFPkBrqcQl
n9flzEp/qPxJwaJjAtT6nqNbfeWaL1gvD5Zg80L77WHbdGdRmxSXzVbDrA2s53NEtH4Xiziwadhu
KR/5n9sg0nhPkq/zyQO5wOdgUc3yMIt6hVy3d9k7UF+eOxkA1iBDIwqalv3en9fubPhdDjcJGJz4
GD9uXrykfumORGHn8RujrD+ctP2MZj1ojlFv2EeJtV6XRme7R6+0/Q23GMdplEllenXoQrmHoKyd
ATnzhUiYn3eFc58qgX99vOw1PboQqbnOc+Ri/pF1STlFC66+Q5feU+LFNP2jmL1NVrr7JtuL/pVG
BXF4XdrgZQuN3V80SRXu2TBwKTbuvpdNCJBDH9Ao35dcBeWncUOb0YQtgyy4wGOX96EPKXnuzUDF
gWL029nEPDYvgUt/kn19Zv0mcHN5WcgzsBiq3RaBly46aoBrTiVO/WCGdsjHeLkGRnlQurnG3QsX
OLNr0Y2wVefjV167jDDisJgd2q4ZchaGqWxVeYmdWc97r3qfp/Gt9UCcF2svkjsmyGFzlE4EeEou
wzcgtLhWo8rcNxYw6iSSQcHnIe5en9lpV2Vvv/+ZXmkrfwujP4I+zXk2PP2ETY/qcgaSvrj/hnjM
gczte/Ci94MqPW97Zmxv7J0P6kRWk/md0OGG9OOA4HnhH9qjhFZMz9iDGXb/yB8z2zJ2576dCtTj
kKWPKrYcU/3J9BiWawoUtHisGptczVlsWja9gHmudxRs9Lq6OL+YrSDyYvLtaag2GVJBTb7ZJKHL
obPyxSbe4DjnbgjWd0g2p7PdkX43xCAxNB+g+SUQkbtQ7PJWqybpK/LTDAzW9NxSYuHBIpywuF6X
rKhLIq3IPeuBy/IG3vN+KKpb9xR4n0LS9pk50hMW+phQo1LnQ2P3UZxe63RsU3F8opBxWQCiHKBw
uI97iLGOWmCBgtG+O0FxE1ey5um1rftNfjobrXIelJRttBcGi2rYnDjNSx8V5LAuRdFvaBo7MvA7
+Tw4oGufUqFNZx+uOS29UFoaZO4jkG1AxB1e76Ugz/Svy3zMtKJzSon72OVezxcnDEGV9r1Gy2gw
C1hz7cYl9AZdU033c0wJWkNub4x+jZ+0+PqUz1egK9fajJoeYZjxOVKahqUCHVb9ysyyR42nOeiB
BxNCfgtd75ZQ0W5qWAheQDMsJLHAifYCMpQrslhs0j7nfrcLxKTjz3zH4MiVxb/ZKX3TVwxSBZpx
Qn1zvVDGFOaXX2MhuEnHpIEBVto2a+uPtTlZELR88kB294xaTzPiYQxwqod1dzKPvu7A1ti+QmtJ
KxveHmsR+pjM+fw+HesA59VP4Gdg9z8o1gtuRBk5GDGhjVcOue9Tf7d7zIso2l45JGLFm5DaeRyb
uBHeFfBEPu1w46ueLz0XcCCPyF34tAghcjst+DRPmnChz5Ux7shZ3og/FLpP0u5rFv14S9VkCmqo
7920apDXYM+DNq15uigkhQnB0wc/soO/+xk4M04nFMPsHkbvgh/xCIgLKeJPZPmV/6qLguEIkGi9
Eae6rKMq8kLudzqIXaXukjs5oAgws0gdTBVftYJB43oDr5d/fWdb8QYLORlTDnTx2Kl/SmHLQ+BS
NLSqnJHnAmv/0aHnxyC4g/FSHtfxtT0BXrcuvUJxHzX9dj+gyBOwmayuxLjXcTgXL3RzNqiGk+Ij
oCVsTS/H4HgtWQ8unPKF2yIHF2JNgWLLqZ3SjtRZv11K7v5eUscR83e72vxQfH5DBA7DyP0930a/
19dIpTmec5fohnUTDVD+qQIf3cQdtrhDdm2hEic3+W1M1qmyNl+PY0o6ldwAPHDFuzjTSfN+l/sV
yISowVj9xdWal9MLrFdCKr+ZEBuqwHE63ORA5ztZmkPosmsr5HRxkQ4V7ZSGUlZHWcZTPK+sCXH3
UiJBU9odOIy+QfNGCM8LtTTtdEi/E1rrOF0yAMHz6AFPeq9l5d3tkR+09JIydS5H7gfMVw3/IIbz
9oChn4Q3Pny+fFpVqX3UMPpYM/m0GsJZQZd7PCxG7+YN0GHnbEftOuY1X/E6OUuZX3wmNO2jGvLZ
POFW3ah1AgjFWYKm64VTwQMKAlPIo/WOVAP4hpGTZoCXGqF0te8HOtDvv13QHlyFWoMcfG4WL8UH
dZyvT69GMtKJB52qD5DVC4BuWoTo6RwF8jN0Jn5UWbQASTjutBpnpAq5Cpb66bSZxVlT1EzbawFC
u/6TT9BNZxrDB0JEKj0CjmRJIWWpRVDgo5HgUumOfDRzAkJ5Kc2OEKeYR/nZ4hZtBQQ3EIrQqjni
D+QMB0WYDdoxW5hSSXo4x2Pr8T4VnTiE1XT1BqKY6hCEwNq1O77gtmSY5d02yKS4GCToS8O+lwKC
7yKk8EgtB3L17M0IOZ9YgaXgSQ5yha66uc1LoYBMprtej18yP3/XOJHxrjCmhNvb4PMdU5bwFPh5
wF9BkdIzGuEL6/HjZEEAZZTu1RwXrYjpgJBTBgaLApv//mnD4v5nCanCO13yMo33dwRcyD21hIyp
kbklysRrrkW3YCy0OXgpGKDxRmr2A9OGkcXTSuv3+G9gcJh841ErlTshzV59Xn9Q2bN2uSW86CWT
4VIHZvN1BIy7/4lWRqz8giuHKaPZv1Emm4H0f2pgKVyiYc0z365arEeW3KXBMqN3qekEsOElPkSc
NOxO/lLQOmPApP5TOmaEKstihc+8ujjAH9J2no41Nr+s2QdTYNzaatN6HoiqbgBzuf4CR7sSGzAW
ZP7iD0Y6i2sQPdIrdkyZTgAp1kI1b5Vg/49sUC/m3BqAljUOsKUVvaHnOazQ1mpX6RPgoKHchTVY
b8uEdDfqUjWCu2p/svV/hP/BLung5sPaXdgdBewJY4xgEgDh1bODGwuYrB3MpqDxWVczx1+yfCG5
n6yuEVxfsl0snMXh6wj5+6rCKWWR9DIVsGtWs++ZrxAcqBgn5L2eRD6svtK76ekUYX3NKno2l9GU
UNYX5xdmnlxGOl3V2tGwsavW2YZV28G4GdtgUmxfYDm1BYW7OOOlPiynQCjyFscgZH0WqO2V+eHm
bRZNwteLyJsleyXW60cICASyK9G9x5x7tcaX1PGppDQqxzFn9Gxru8fmD2AmXvlwCGKNQSzDT3VK
CWA64zejOhyv1indys2pfIZPE37pkAhoCaUbu3Xm7zlwSzclErCcniK3w3QEmj9qwexhLggfpobk
JqRRKQpDoGfV5SuJxwpgiSXH6dQA44JYEgNo2JcVZDVAnaOiDTMYGgMz0kL2Uso/yE0Ef4MlUy0t
EJTK86HD/gQaMk/v9KTdoFvcqLDj2M0OiBdlpcjLgg/bz1yx30n4sZX5e6ZRPG2tcP7bKvqpzIUM
NxamYwK5qQGk1pvBfyZKibg3ESWltsuLNR6VNN3QQZUL4hVviKn/mehqB6U7pBfp+QtIIDhUn/Qq
pa9clJD9y3hCxOlzwsd0pogOGvguGn8Wzi/2uhlII6uqPBnkvr1O0j4eJz+ZnVYWjmWp9VbOUzxW
cn7WqD0XBgNaaktkPFsYtFrSeqWY/Yx9P9BqUA74iOCO6uE9wMJ8bjtITFvWNsTdJ+aT+UcHf70P
jx16CEz5lRLkTT5lAg+KCtqmK6Ms5N5I/JXvJ5ehBMq2CPDsGn1J/6LYXoHlWGuaB8aMpdreon/a
HFoZz6tx36AonmDmBgifsFQYAsbaaf0Mv35MFfZiO0wMhkHC6/or0IV6vtYUkwhOuFb1vTPwEr/a
wp0Pph8x/mEa5emKbAELSabL3oL7jDGCEARpcsU/LrfmTZRepFlVmq2UgYKH59PCz461rGlHw5Ma
+f7ZSR189kYX1vvN+bsbK7qXoK3IYx+6dOueaYtH7gLxsZq5J2IqDrn/WZOk0Ngcqsn+8S/LbZfC
CSUxm8yHUq1BO6lrxsbWz9InWnu1CZ6QZ0l0KVYji8G7bxasCyC6rd3GOVdqwOezuyXRvmf11S8m
LRIlIDpES0FfZqXfNxesA+D7UJo5U59MKsLN7eBT3EM1+OKyJ7iEvKT1x7lzYCY4Kl7BGQ1fNP/G
z28+y9lxgWAC56pSuXbE1xbtrOV20t9oJWBEBDO5aBUsYYG+e8Myxx+ckcPpqyIrsj+P13Q+MYf+
d43DSfYX8cWrauBG0+D4SNKOzZ6Y2NByD4dsnc9h8xJ//z4aEWKQGSSvjj4JdSaV59rXlU0T1c1T
3nqCEdHODrMRmkFuH/hp+fspVqfOEonZgYfBG78pUaPSCXhYqEqOslfP116T2dCRWfnz+0/6lABS
CxlW1nuhawP2Bqv21RpklfiYtbMkgeiBst189GSmPUqV0IehfeYtAQS013LbVj81yFpl4hSfjL2b
8k4nNpbkKMAhIdwdegtcjLs0nzhPdhQeOp7sBt9XUcbv9PTTMCqo2ra8ihtrxsgmw7IIhd/BlkVk
mVyFb7w4l5eDvH6KUUuvAR90y72EZvAopHhRefHs+HNwrnfwV1ny6/0BznSHjc+bTGYZ+Kw217Tu
m32ndIEgolovnuAlA5Rt4U9a2BWDwoWMIrGNgRjz56GXgb7Mu6hzWdlXzvfh4MWfAZjasvlTwVPX
y8ZH2z5bGceomqcwM0GNcPBhZpJ1NkMdp2dFZYiK68SdHHGXkhX4l4BSQ7N+22T5+5Pssehggn65
MXFaQPuCLF+LwB3ThufrwQxnBtw3NZynsgJNu4jfBepfP2yn70yiGotgUhXVq4FkqASv7HqhpVPx
tHuZAXdBmomqbuAmIeY7dzOpSbEBX7zmOKjsvGM1U54rMfIB874Reyzq6dYLs0E4+KkTaJEb77n3
lVatUD15RbPrRaE/NcwrUMzpLTS3TWr1xQBEPzBEh/szjtlbjhUTZmVNQEEEMnsU/dA5Zyf2KZd1
lFvA7IHo0Pof9aeUq+K84CJ+29dK2fobOSEVNaWNR88p1GcAhPqlDFd6uQH5F7IN+/LXlJTQ3M2e
Hd6MDiyoRq1M5jJhnDV0CUPyI4/iS7CBoaPct430WttjU1EfqZloUPGcuykQXEuzgQbNyUAlcblz
aRxPu5w2yvyzLohpRD6gSZemwqwWLCXLRWUEiHd6L5Sg253dppYw233bigXL6qHVRf27XxOKIc0Z
T1reHVOHd0/ZBvsdz4sbLKXLxZHhHwB+uv3eBFjiKtMYoSXfozw8JY68rx6+y3tl/7K8UMabhuQb
sttQesfocklgAOO1hvgZ98doGzjcMBq95SYPbFNPo3KYvuuPkMHCMotEINI8LmMMyKXzSv9nMk73
sD91lNWASiSiSQD1NXrh2oMeLygZsL2lVgMiskKBGPhqnNTKSJe8ophPaqtj6IIv5oN1mP9+sSdD
j5NJ4nqjrK5rSIMLlptbzTVBVMluLldLOiGXZcKDxHvGUEzelRwiqpjyLlTzyL4urSFvkYWJJvK3
Xp8sw3LIyhv7GTYKbLiVTs2VBwyikl7bMvODJhbwMYtbc+ROCc3rzDU/YNqZp/SlqzC8rGuNRx8l
UDwDnJYrDGOLeBZfNhuta6xSJVwhrtADVQ2E0OMqu/XkVJlveo+m2lfdxsZajB5EusgncMfffRoG
ehYp2pS3ggoLmYB2UBbY6l6cZSgSCdsp3RSr3TeBO8KkYn30AMI61GI4ctVMo6Tpt0Q272plLLEk
u0+RmKBvXUTQnq6TP9Q50SSr/KJWC79wlsgwg8eHm8GQsUj5yueF6T0vpUy3+jNB6tvGPrIjNDio
qteOKj06+C7JRIhg7JDDCez50jQ88cynYFeasqb6e2tiH8YxQNkAan5Iqz+kDd7vyuScawwPbAFI
XEB8DCTYvyV7ymsAQemkVAIKKnnTahbA2RvGTFo0jVwx9D/nhrRUMZD8BHiZ+6MMruI12zUkmopR
MLL3bD3jqWw59IcEirgT7E5BrU90yMC1CxRqorpUImSabffUekM0ZO90XUIA6azfXJgzWITU1eHA
crsS1Xr+W/pPbEmrKhuW4J2ITf/pTejmKIwT7vsWsqeI3RPZskyttdRYH6V6YZNAO02RHG3lAQlK
cWlwQKtqwd83yMW1A2N7wKdy84lIP0QjYHnT+NfehULjS4Org2P4ay1t96F5+vFaUWo7epD2Lbok
++CdhzE4pU4XBVZJrsrYnMiu/9IIcjx9iSHWYQ0xDJYJAuzkba5d8XCfszwInMTPRfS43D1p2E7w
liAetyOEucdlk5mPGjeJIWuUXpgSHfLzNxfe3JTaK9J2aDiU7P5+QOrBwvVfdTdlVOKa1sy5+A0R
5UzAHJgG7ZdGZcgpzBoQQrIOdx+0Ei7Vuh/mX4lHIjQes6WuFv1Znh8uBlWySdZBpM9yPlgAHFkd
HUXgw4At8NaNPu7F3iJqxindO1weDUrPpj1bxudiCCe6XlSQmOCkiFRcD0yGIkN45BjxwV2AJzOv
oM27F3wPUHj7hmAGZubx2yX9Qki23h8ff+eiBmoWa+JMjmTZYL7Y1ARx0nIXf2eFJlEeqReYGQ1p
tHsYvETKvAJadi9x2iwd9wkHaPZCN5Yg5R822jJoZNLr/g9XBZVAVFYEdAzpM8xS1cg2CZHdSdt8
1NCxfLK3aLIYHaoq7MPEIKtbfl0p6hTfZ4s3lQVFlz4WFkVg9vDoZHTnfkp8Cta7zcztLtxumPOU
esSFz5O4bBGtQk4WQs4tTd6xhjpsNDH0MV6rqb6Ma4eaglkyZIy32zTOUq3jH31bai4aVJHvtREN
EbBGahLrmM3EpEu1mPmoa17Ikl+Ri7UF3iesQsvVsz5XQO4b6qYV3EA42F/JYLxIJtBWmhduprF2
bG6a6RipaAeb4UBhF6IPhQHnhy7wI8FGCYmdfrtosODzrZZOH09j4jXNaDIhTnSp56BCrnP0kIJP
k6QhvyPralWRqJO7mbkFAyKL5UFyqVxrWOKCufFieAaD4dz9TvGumUmYbniOBfWODx98u95Yne3z
uukNZTi5Md4Vp4dcxgu8W1osHIpvInolARdi2cg5ptnGTBlh+WRvD9h14UK/5LLEuxe4I0GN+XZ9
m5JII/chEnFs6Cxa8dKs5iSH7CqEGG5j295h+LBuFjA4YzVTcd8Oz6TOAtmNB5+kO2iWpHMYgp8m
YwFtAL0nQdG0yx6PzSZEhuuWtRPaA5cbSvNeHSw9SGUGYfvBfkSGb21EX0HBeA4MuLn5GwSucY6b
bzaDWhOsviu7l2BVpNDPSk8oVGqE3aOIvoPGfasWXFypaRoiSrMTM+ERjWPp5rx4EYSqRDxy0xew
ZCilsfs4bgXPaMnHVFOIqhL7871nkjmc6Kpxaqlt8ZYTjOx90YGTm2JWIRDrXBCbiZNFMWkKaqYY
vHrHFPFR8ogV3137blrsST/tys2oqgq1Lh6R/viS2j6ZWND0d7jxC/7er/Bvy6c0lKitbZld+eeM
jm4qHioxJwwhkn46je53MaiVJ6sW3VEiYTHDfuAHq48U/LtTnVa+wvJYO+OF+LRKZAywii3eItCv
uUNsobjb081R8rmekxP85pHN0HYJsS2iwREwvJFmpHyHw2T5bYhjeUpQtyC2EBXSw7el4G/BkNfc
PRMOjoCvMXzHrIBrG7/UB0MxPKAZQ9QhZyqXqp1df7rOAplxw35Djig7Fl9MNm2uOuPqiVTRJyEs
qJWeT+b+77yVzbM40HcgTIJTStTcKtMF+Onnyge4DkkQ91rIBweOLDLRXLzzdmS+ctY5IWK+fyN3
zjOLkGu9D/o+p+DtKjTUbHPzDlq2ejlZgpxRT9t/VwSa4wPH9lAF7dN6cNQ7NxFybefq/Zyq7yM/
vC9n3RKJbXlbXEqPhvUziZlsd7xN8YBKUzQGhbctUgUMfcFJdSAoyHW3i5aNBRDSbkcOtSGvrltS
clqyx7A9oCPAlIuZh156+iHoX+3aOjvE7mdEr3DCfhAVWw9CXtl8UtYTjHMo9q37AfXHofRT4S0x
Zd639ooJ77fVgJQ1mz1dfah39Z6iP/CU61Sszi2TTfuZe1VbNlWkE2GrdEwCM1jQ4GhIcEVNIAgP
MtV2BZsSOAS1cAkuvnOu6KFub6usONtEe39ebSf2wQn5K3v2lm42uTq3/0djP5yPETeGQvjgcPW7
vYctsQP6JVhTMWSHZXYFy991W0jGoU61oGbF5v5uqXfg4Y/Q9jbWPaAs/LiBea2k8Ube2fUotCeg
W6s0/pgj/vMcl6HgSp8IovIlPDb0+9bAZ5S0EeGXSq59Wdyqqe9NDE7xsaN2dwrD4NbmomnZNL3B
3WdpCrKvsEWEpKWmQyWk2XaAuy9ATyYJGCbCLdPxx9LzLYQiN+ypkuRjgWnHb4Z5aKUkisw23pgT
rreQbAucV6LyT65CXyjtDzKNmWvnhgIDV+xXqTdiX0I7EJSCUvxdrEhKCR3pbQyt4VQPbgd1gLDh
Gm377t50wOvCmUeZlx2SKPjNn/wCetYxZ6jMFPLzPzOewAyy+LzG1eDl3VqUiqR9GZSV3Yd7bFZq
a1TqUJG/WzE9+RzUhV63u3Hf67S/2xjh3uFangRrUV9B0GSKhuRt6IVLTiImmC48Lc+s34ppNCOo
J9gRmz4VpAxbX1V/5D5Y5horGAIUJ8zTrjK3X9zyLA8/TVzK3yRKFTRNHCln3S+kGzkd7R6oKis5
SMz+VH3+UUYPsyqtQpCWLQLuDmConPQznSAu1SoF5qGY5oZ9OA3Z3LXUmUiL60aCduYCv0sX10Ec
eto+eXJMAsZCFUyZA7Rb6FHqHk6xCO3PrLHnEFu0p0GrycmjqFRJeP5zJsFKEpgqYXgpELpUNwgR
dfpqzjKdx/0kB21PA0Dv5KFKePy38tFl9QKIFjDjEtxPhrRv/rUozEW+YHDhOJbTNgs2Ua7MnS7L
VW1zHDLlbZPaLh/lfwmnflGHqGvGH8eevIeVvyZfalH7G8kWQ4MGYhDdOb8PGyb5OwU1g28yG2ny
xZyph4uY2fr6VeiC6ghZQTIw8z2cLSPyEFz+Hy31B0e/VZULAsFsRbUriIVJBMan3IiBZwl6IjMz
s1xMZRvOcOW1C5dF3Q1KU/1HQjHElF36mMjGAums0irfxu8vM2Swd/amJx9OjUGhqbHL82I2rDJN
bX//Xa2hcQutFGFnlrt8S9Ag//rnqV/pF37RR9VGmfz9Ob1KYQxOcvH3XVR1CYtsvNiHG0kfF+nu
h4iR6lmiG7UwO3p3BWq1zkANCenCnbVMz1bMan14LQVaf8PdjHGX8Lpt+ItAOaJhoKqui/rUhkwO
UwNJpLxzb/Rg9qx5HvU3zwgWmHt19aSE1F9AK2qdv4O9ATEZ7WnIQLfyY5v3MD/jCom9az/LeE39
DwpfIUw1A+auYhQ8CYF35EXGIOjXrFsmtcEseZhwirNL0dXsgBKaNcnlMM2WBnKPTf+yu7PdWeL2
0iVbsrKiqCMgUpufNyWy8HZAPPfpKGBBmtJU8N3BAFUgLICH4IWeMIy1CxUglcdd5dUY75AfgizS
89jHVdRXF+mzr1CW+h+ce3JFzW1qGv7ayM8S1kyS7Bz4QXm8Tb1UB8uHEe1c5wXu+jBctkQl0Taw
62Hi2Uzx8kapKJI8hQDjlr4OXIV6krfPFvDvVE8sRgkH4Zuc0LPL75fA1Gh/MOU2lKOEHXx0EV2E
zGnESvouQDUi+VH8W7yJInm+Y1mGz3LX3ZvJWgDrdjsfT5azknNzu34lrt+CEQBD5joS4o86Txqb
so/E+lksoGin1zDrmh5JsZG7ReRNQ+rnAfE6DpyDbkVUCYSFhA9lwtMJ2wn2VzFP8+5rNiassLAZ
/12chOqHjuyMDB8QZotL8ZHkW7Inax/wTlvG4I7Xn3C3MM2CCFKEW/xDNM8TNgE4FlB50REEa6Es
SUwW7EE5wsEJK/0bF5pHqtJUZDMsgG2DIxeeFxrcR8Mx7rdt71k8R7aZ19BbDStEv4004j6w/gJY
3p4txm1h4/qurQjtWLWBxcsntMYViF0dTz/Nxs9O6sSaqvg1Kpfk9fqxIF0reqAO2oLodPKDvJKz
7LAg9qioyZz967XrSIk7xv7nCp6HeUfli/kc2b74bpZ/2jp0nH2gf1gJMVND1YGVXZldZEvVq8mx
N44adZ/jLXd6PLn5G5mo4j/UrlNoiCpSqMpjVgNqhERYy/MF1vjXibJLpKL3u0xY5cLqox2LEPbp
zVL/DsOZKo5lBoa9U3Te/ZbV3XFl0hK3th8R7AjAr5B58gNTDWXD2Lcq6xoTBiSl/K5mZobCoJrG
9ulqG95pQNfTxSNmHxY0Sgvo+Nj9XcHl/enN0hAJnrdNURZ7xoH2idbahMRGI/k1aqyxqefxFKAO
bszS2Zx1xqN/UGU02CrzV4UwspylzllMtPEKfJHOu9red1nxhNs7I+8ETulgvemL0zNR4GA6OSM8
gOeca1qtaJ2f01hiKknrKKxiSZm+NmVRgb0E6lRpMlVw7KzrIxKNqn6goyCw7WAnemyLGT1v1Ejp
Q69O61usp3DK/SgNC+P+ebdrxfBUy53hXdKFukpXUo3H97du17ykRR29jn0lAjxnaxMfBMP4mFUk
B8EBODqCYOy6BynPIG21e6QC4E7HZhWsBoIIxTp1kd0cjomU9nTlEWU79iIQ8Z9MSkWy3BkBab1X
DJaZbTjBmmhMaca5a6TB4g9OPA2fh72eIYGXN9YAp/XHLxqCNbrByfnTk/NuL85ooxLSRpp3vzIu
rJqLVHP8AR5hzLCSUNNeVGq/TlR/aOnxEDnZFkn8h1ZaUv5X2TxK7duv7FxsVebfnVPeDWIwQ/3h
wfek6LH0mARHHQASkrqh0eU6Ml/e7us+hBN12WQ41JJcLat22TGeADr4johLZwwmLM4p1xd0rrja
F0omUxLlakY3B4RSHKK3A4UsnxJCj5mCZB8d8rbN0X04pU5bZk0CaNYXLY4IjqKeU0LnPnqvfU0x
RnvmvpD+mFsSIYFDMe8jPgs3mZrXKG0rPSuZo+KyYFV1s0mS7NlXDIzZd+PzpPoz6Y/lN4iIvnpj
bGi7QF7wsVZx3adWF0nHcAMBuIxXL5p4etpiTaqrM7L/50uHzGmv5dMG5HByYxC1eXL5ht8012gU
7fJsp+wzCJmdiyUf70Ss+VuuQq4mtotXx7n/MLhJMrli/EqrXkSMhM1uLb29k/zJMUYZtyVbxNhW
sfSESu6Sykv1c97LqbRxR0XUBnwqEOurfDZlI6YaDJSndOuyR1GarYsfr/hu9i3njUkKLQ9/3KvH
L+WIUfkYgbibh512FBaIzSsBQ0SCy9r9aDd3sC4xHEQ8y8vBTN2pnENNJy6BhFuBT8VQsQwOpFs2
P3HM2oKCGvus36Sr8y3+LSbUCKns5mPS/iBhxWXGbPuqthXE69+G1TaqQowLXaX2lUJC9Q2MgE8M
AdQMkpMCmriWyh5lDvYC4GcHugFQYohj9UeJ2PmOoZg4IOteI4aNQD6bmFoyyi23PXJwfYai3GIL
fAUeiWu8t/I5eTmpIy5bV0V8CnX6o04RwXBjYxkqmZWaRCBx1u6aymXDp6heTOX+y4sg91UcCW0d
XX1iHmmyIW7Ol0shhXzCX/r8+K4+03fbO8YRfAlh8EwAt0MC81oAYlaz0CNU5fgiOwR9AciI9RpD
QLsFNVbpZ9D/XanJaaV8bEybyt8oH6U3K+g1rbNnUOjtmGjdWZeWauHgYbVIBL2/yDM+oWOJy5qN
OmDj5ZqqR2JFYO03PAKQx+V9xO+6mrdfYhuF1fXVOf7iuJq93iMXZ3n0fyBzm42lrxV8Jz/+5zUq
5ZlawVwq9/inOE8yDnQ/k5GMrzl+1FGlUMA5PpQu4r5PSOON6pm4SnemM6MlmQSq2bEjzlAOvwh3
B4ODl54hJ+bybxMGYN1BQVEpiA0gNeWo4sUpX2m7e129D/NDefTauMw9WWZbHAlbPxxTqi7S+wlI
g6nhFJp0kdXjOJLq/b4Gwk7roIhsDpEtA3WWTCAJgmHOd3TVeuO56wvbdsVg2+d/yfL0g0OCLNoj
ZI5uyQsAfps0cV2G3XXquY0t0vlFTN/fLD/6pwx9jmeN5C8IHQ8HG8IQwP1TIoY3yg0sFpsl63qb
eWeXkrDr8mh4KIcUz+UhQhGV1cD5ErS+mF5q4QWh8kECIinGbs+uZpKt5/vccIHl8msMKu4uDj9h
Q5W6yWvVZ53Gn7jEuvbezi0Nmj30XZXnGaz0492OfAisseTOrh+Z8bYcsX5Z1bM8op5BtGFCeSnk
QEbRVXbe+FOH5bdCCSrN50/nwG6iFOUuSE1YPXnsfDTBw9+7mwp1mUOqxZ7zXghD1Pt7oq84XP4j
Cf1aNZ/s9fLbhRO3QpQijdmJd/DxSVM7QjhY5WWNDMb7C5y36kDkkU4KrpaXqhoyz3RqtdVQTfAI
KwPEscP/XRY/ccRquwg3AkzSeC2OUPjKLjDA6cJSCH0ZuExPnQlO31cIP12v9LqkcDC7RS9daOlV
/8oJm00tpjTIWo+tgTOqa85LMO/6HXdnUZQWJ5C8/nzEGRlrSdWMtkYGwAo3pPnDMvJEUucit2Yg
4+BFdUslBp9ZWThgInnZ5vtFq3lI6B0gJHPJ/ZFKldKgyxzSV4yFQg7bvz5Bcq3hzSiA9jIpBSQb
I529QG0tcJQ2QBGpibuEGbsijRvgqNoBiPZR6wq+s7mU3fglBxqOuq3+u342kVpzK2vWaFJb5izk
belm0YQyyQWlKOjOO3MlhO9zVCdL3EQNfpJPfd+kD6xp8+2v8W2vGWa44WpDuvDGH8tEefJ65p+2
BCe7gr5DrxNQPaDLU+T4Rq+zN3KM8yAkIylzCyTBMuwCAfy500dLaSGi3R3x+KnLW3gYcR6dVS1O
uHB4mWZ3Bw51x1Jh8mp+XIh2kHqcveyxs9yGos4/E9ZyimKWWgXt7D+3mp3oa2QCzPMo7dEggGiA
LGWRYoMv1AQty5RLCE+S/UyDyy+xY6jUoHNr8wO692X7XHHHNFdGe+sg629tDXrn8ICkRakhhFji
Pvx1OHOnRyVOleMWw11cLQ1D+qsXWv8qYjSvMT9/jIYyc8lhDelGZYgYV42rlC2E2Uwi2qNY98wJ
i796QgnMYDN7sJn7QgNGLW7ERE8d3+f+zkXaNs1IB5RyOpGUIQHW+tAGFtYQFxLfifTZEbKDy7Nw
d4mYnWE2+yVYilU78UdHKqsJhAFHXZ5HMbFZBzRyFtnlcF4BA6eZzZgmilTP/F3X+joFdaF6kr3o
K4Q4u1PwtPJ8l+aV5Sw2Tpw2QwETn9INljBIZE9jFObDxEz8okWMVs5dB89tqAOgSTWgYUbVOdQ+
oDNYQs5o332u/wf20WcM6nqbXTPd4eRna476clQEUkSH6gVXR/fLucuQperGO4f8ExoC401DVXjN
Ska252bTz8sjVCqWXswRzKCbKu7QVEI23yJpzOeRxZ5ImxgVQkKan5W8aMLZh4cCn1p8/ka3tNQT
pJvI/hg8SIPeMrqecOnJS3wynrasqcZsrdgUdjyMON/dSkNjpR/2dHgK0kKsswwGbnbratTeOe1U
fNrXR3FL+c4ZgXzWi33ilGeaXiDWtfX+KjEn+xIL+ByqfelNPIoYf6xkJcRl57O25R/ftCuT+fYz
9sSBFOlYhEY0/XgNlxoLRC7rdQSG9cCVFLtmm91YE86tSTOXi2oaN/pk78Mky7evgpzXee1QpBd7
+K1L7BNRi5nxf4QhnIRcf0zWhCG7ycwnLHG5O3Xd7KwwLIW05m9QEmXb0qIlE52bawoLShwIU+33
e3SumODpzbwgyWFsglIg+d3lYNoKQ2yRSgViRhwHR/ia2l1w0mawHH5NzK8a/FlK4fLLl7YwXhGY
9I68wFFvtQmWE8XtbdKn6kB11WMdo9PkytgFOlM7YZHYumqMfmYrGq9usjcj3BqOPs353rJuQpNq
tx1Z84e1JX50SXJEe3l8UQG497Vzr2tsB04FWp3+gfLyYdRTDYXcwe6kSVOJcRxCm8/X5imnjS4x
pY9DMctpfTdFs4uLN7bDtccrITuE7Eh1knYbaWl23814Z3ThtdlNvwhOH8qaLur3qQjoTOwAysHB
DpwWjGldT5bm8BnAeoDHJg2VW7mh5+0+bNNtvRKT5zGMz3JDHB+0jkAEKlsgw2Z1Om5gsU5ad0HW
5VyIOn3s3du0yv/rxxwVfyvrhqkMXuoQ76pkWFrXdQBO9KQC8Aj3eVcxMl0/kg1VVO9jx1L/C9r4
kHPilNchnvcJeZttkYqth3bXr9h9ZFzFP9tU2+K48Q+w2f7pNrhUsvGxk7p50mgAC8iCQ02KwkdV
Zf9ikW0Lw7bW6GHIpJRq8XiDky+sJWhq9rNI217l1uOQLWqPWnSmPho5KOkYMWCgHSS8uKw8hpMV
qu/yOPKr6pVj4wPOQfnSeSteGBQyoQoC1/di7RDFEltExRe0rqHqwv3btv6F22yxicRGaxV10w7W
Zp+1JsV5i33d9Oh/lTTYx6fxok6jrduZTs7ZuPCb+avTmtZwA6alCdkwSwkTnRP8YA+fP3Or1Q5r
Egco88NWLm+her3pdrMoMc1jG7MRpR4bGYyRhNoAbT8U7VauTg8HIsWlpVg747F3BSGeQkPfiFGe
X0ZSSlZypWfsjx4h0qW0CGzH9VNXKCS8FajcD49l970R6SdnPEI1GZ2FQvHwg2uyleRk44nCoIE1
aRMnPUjbhwz1tm46EIfyooTbmrfrXV0w3shNcgui1BPDDfWQUqH08olJMMiOtgBvc4bEiUQyMt6l
oaUNXibum+yXdNU0+vBkFPvJEV8Y39k2EYEWWs4Yki6odnNiTlKn0bymcLAH1d/zJsCeQMDJZusV
r+NR31E99NWsQch64tk68zDS892JavsGreOtKq3kbZiol09+2lqdZyn5b/jl8bvqEcxhITyB40wi
BY2tKQFWpE2/BRPXhHgjmAlsCA+onqw+gwcHPQ6h/qHSlkcZvySdQcFU8JYX3HFQ0QSF+Y0sybje
lxawOEx58nUyzSUJ/RwKm5DxSCZY7HWKO1Mckkbesfyrw3hhuw/I4UoAdxrRdjmoBjB9NFQ9SJiE
Kyf6kuf0CnKY56h+lpWPm7n1aqHMHjdr4TbEYyK/D1r4VxYPW+RNMnUh7Yfm1GwHNxtg9ikeAW/l
L7sGwvzd60j6XxIJRMP7wqmpslX/WkS1zeFr+uCtk9Pu5lqaoBMKHUx+9UsqPAfDfyN+//Mpo1EF
WdBgEcyMCRyyh5DxaumwyakiCeBcoZ4pypdlifUDNOZTrbgG3MITi8L6zZlsy3vn1GCpS9sOY6lg
QoDbNk6q/M7XDPL2MGpH713ogHJIwk4rTpy0L6xCiZNrhYJQP3Br/1ZevAlm0+8hZJ0mxyHHp7u6
EQPv5nofqCtzQR1WlyDqr+ceD/h/m8kjm1NeW/PiCR0c0QBY31Pv2LbYKWHpn910xMpGKmPWMjkz
yeHdVw3w1fs3y7vvAm1gRi95vpOTmAX8XsQwWnwR7kgW8ruudylj5xOHkOTkIl8SpxdXdZSlUEx2
V25tpZLjN1m3NZKL+gP2MZGqlH6V/or5zooxOw/UkLgnjzyDkSyfvwdxZCOkQLkradsWk00LK3x2
PMRTm27vjuWA2+ZsBYXbKjU5Zs5++R9Zl6jM3aBDPXnRSNHKB1eNmTMth1Jjtwv/tIazWn1q6pL9
eUJjRDmrXbScMBgBIE5YavFdQRziaQWbbwqk2Y5NywopUufjP/xRwZzC8CeGH4TPymsdbRVcWx9p
tZ44+eS5nZwZRxefrGjcrFd7KPyLrHwycerMXhkPd52yuYHdqA8N3+IJ8ki0lMsY0ndE/EyQvlzd
W34Y97YJ816aRQ9l1PreLjk0xVWb54xM7u7XhsYmuUrFKXRoULJVYeTJoEIGj81q291knRlpUfGG
4jhK3bxt5O5iRQ5QUVZbIqb2XLQ9lcXln4QxW/Q7dOq1+HpwEQ2+19jBm3I+BdcyuF5pujBlcToD
KqdO9xkxiAmSUoiiGlx/37FzfkMzGGm9qOAdNI7Tu4YQEslkxLYKUIfLMq64llfSMs1V52q2zubF
dfuJ+eoS4shfCi2eA9m0BP72iG9UtDuJiuihQNuWrCaN/R/QxR6pHr86fE3SlTUjpUEJpR0AIzmC
tcaRfUfhi5ULZYW8dhb60D6iefe6+T5TIe9bK6UwCrdaxRpTXanq9dagZBKveh2RPkDxUIOCbLjo
DZ9Gn4UENgU2L6KAHRFCZt1egiPcD9Wm3pAT5SZePZTC1GSTLdhw6VRab2Xwq0CWmBgVTjDDc+JR
IboYIuIpCnq8KUdenyuHJUf+VHjiFes2SLOctlBio8z3NsnblqVcFQfDCXFTCgpjuIXptX4HtSXz
jGj0AldNS5WNlvNuVwMcEVk9S9/ImE94kZV5dD0SPIOrGMSZ0A1pYEp75ZmQvNnyvXpLExVH56ew
eaXwU+tOLUbCPtbrF85N3hH6EQwRaZMVjsTvZADHm0P8ntKfoiTlGaRwkKl721mPwEs3QGj1r6wY
0J4duyVpAudIqcYaO1miTn3IMlCY25bCJiNFukI23HBBi5SH2csq2uwnYVbxIsFdl23drQsxobwG
r4kiZS42DH0qXMm5FlCcD+Ivq81orUj6/qcV7EUBOrslfVcBsdIKVO8ILFYl/MhSRrPvmAtr6mKa
jXaw4wmPxpT5FjdaSVBOdQpxoGYEELx6Zw0/RJQB1MCBJewJJweRLzVzUZdnkMV77A0N6D+KI+Hf
A0HEbPVgEnpKdnwJhvmdm2zRV6ZY9baqE56RkQAQkN0/jBQZBG6qkh6D+wXOUSK9nsiUrbJb2uRA
G88UsO7q32b88s/lEQiLRaz3lNDdcm1AO+6bwxYZ1FetuwWCmHQP28QZj2ZFxu7WYtoaKS6cb7ha
ckeh9zqUCELk/Fyvyx8HFxh4GSNhu3mWttdCSBSRN71kbX1MFKJw97ujKB8k7cfd99OvnqVjoIbD
EQhY2FtdTNCLqeMQt2ffBJflYu88n7rxy8MBQiVJWuRn62Wmi0pvIrcMI85fOTZD3+oOWmhC136E
EYvYPW91Cmn9rwoH8WfJLSHDLMjj2CDqbkkOBbCcZPvUGIpzCSW44BcHTQB1f4lrXdTWpS6jJTCt
ZlfcihvGtGC6rSxfEC5gp7mbYshxQ4CajNHdlqmbrruf3qKDgx8AWXkfjG9ZkU6e2Jee37sXk10x
pYV+RpesHe/PCGlnkF/rOJTa7+klydgCqM7caCytgNcJGy+puxAXLU8ov6FybGZHFoCePeFu6TNM
nINZGY2VYhZ3ZRiaxyV6wgAsPzEyzeeIQLsnpwzOfv6EOYDHeUuVwyeYRkt7VwVinAgX63N8EDjT
gcVfuHXUQtVVnMdCRWIepuMe/U1ka/dEYtiPnSNmFgtSHrUX39xis7VFPociAUQmSx/VBOCc9sqe
EOasCQvHqt/ZVKOv57kYBvhBrUVo98CMRo4NPWxhCdFVUQptgQDSybqKCEshPnWEhWA08IpvcuLC
WlKLe/4+bOcfsnhpg/ATkghJpNB227VrGngaO9yzE53osJDmLqJCKCiTvjwcExMAbteivG28NaT/
5egL3/mqjCgE9O1KWonfKyzltZSGAx8u3YydZwjPQvxFOGiYgUeOZZmXmPnmNxfVHb+6V2ystJfb
IplK7vZwgCLRX/17fMIH1gGFCkmZWFaQR8uZ11H2t85HcKMU8UJHxMUZZEy3Wt9E1JYa/FS3G6at
w8sMrAd8aB5pAfSLR8qop8afQzN+LZL8JkTGvLNzpuArUf8r/AfzQkJQQfqLfvScOR2gcj86sjjR
pg0aGSFERZhpTTBdPH8K5J8vSFsh3Gg20Xy4GcBlVhL7CGp+dHXSuIw2sDbaD2mpJ2gnlEPM0ih+
EUdoWScgOtbSkYAJZD9CKx718MpnrYEdP9tsV8oT6pJMd1ABaBwf+qc52xBPbBOPyimQ2GEuPY0d
fZBq5Q1eoXLK4fYVo/LT800E/2trUlkX3D8EmvWz1meHZYdxvHOg3IlEZK3yUK95qRlWUywmwd1S
IuPaQ7FSty5BF/YumbpH52qsF7zCwFMsBQ3XxyE9gBPY8P/A6D95hFFeL2fF2frivEC38J2iRAyB
Wr0mGQX0HJ6D39KRV+KHrxXl8hLoKnrWT8iOvr9MTl+Z7lnqTRMeTeriy50l+dAY7Cl03mysme4N
4QXbTiaTvYbzCzvdqxzKWja6ZhfpQsH1zmAu+s16eFn5SWabKM/IEX51vdStI2hjOmN8lGE5jRbs
0mCdi2jsbJTI0JpwQwcRj281plfzsLKZX5I2cF30dw3ElRN3uDqna/4K5VbBZ5D0E2BnRFpZ334w
Yk4dmys+AQ63KWyPfooE0Y9MpjP46Fo0lqTbeFdSZARlSVDl0K7V9wqCrEiH2Tz1fh75qzetlWu/
LWzpFA0ESFkwf9fvg61NXu7LBisTaEhryZRGOkWoUtH6Hbwj7GM5Tl41Vk87JPJK9BrpAg+Qu8Tj
QqhfvKAtVDMAAR/4WwumEHoWvOhVGvXbY9QHaJDZzEy/+XUe/DhSxY0dmOkFGIH9wZgzUe0CrBqV
Bm+vwDD3fpBCgVZt0d+XqKH7AvuqtgWyOscyu/EmKD+xVmH3wEH60egZPDj7ypgG2+guuKTLh/3M
3lfPhVUGHAys4Cj9Km046NJhDQ8xYEa9GtXRsCt/TeJLja/u9UTk4L3CNmhpaUJUcvN0iROAxamg
VUtFtaU+fZoG0njHjS8e6u+RowE2+HabWYJJ7z/+361ahYqnunEDXvorIpR740YYKz+/eNGmjpeJ
p2XF+p1I3v/p6QYR7mwj3tZknzv77mdRwjzjpPZ1EeObSVTX1gkZbwZOwi4NPufB+WEaH5A3WeHf
I4b3gVWikr01gJW5AocYpspRA8RBFglpAVZ65Tqsni6sGnzsAvNQIkMS84FU2Gj/6SGapxW0trpE
RqxEl6VH+G3dZpfMQ5inUXJ/hHxsa/tb5gghKoDOgOjFPeazJ4r9N6ABj6ecjS1uJY4BCTIcBiVw
KKTeoJyz4rONZNvDWRtj68oNxspadH8koX2FzdZ3aB6kUtpNBgN8dwwA1Ql7Aujt9+7OdUE0fgzH
vUP1D15ECuozJKOVO75J2c1WJO7qZNBS818jiHx+WoKWRa36nEznKj0gF8MoKS/2bynrA4ohNZJo
evO0vQvAOpRtYHY+AV+idSLRORCK/4fokwW3x5vbmDpZJfBXrhe7l56B1P9GR5AFn8OZXXikkZzp
gMWmSdnzYh40g9YOdXaqWdqCuzjYOyiLw9CvVsrhZMJ/djC5Ebj4ir75T18xaFJf+dFaO39alD+M
2n/ZZ752xNlaSalwxwzCvrXCHX4M/plgyinqCG0TyDBQJyqhD6NBm3oY0q5C/IU0mYImwfWHeXJX
IphxuoOAeUU/Rxm9gdjVm2m3tXd3f1yOqv6M3hHguhVBCPljEtK/QtgHxqBE5TTccQpEWgsAAQab
Zi/UZGAdFeXj8Soh8V+WN3WDKknj9nSGujf74cYygyleyt0xp/O+flncH8COL2N8uBPQCcQ/gEAe
5/pUS/LYkaTVoQsvv1k50hUQEblEkw2220xJHQFwa/mlnktUvDoQmzvIvUaKxBdfoeBi+qXKiShm
aXS2EBbM/mZAqDsT6G0q6oUR1DiguzlCVHZvqKulQKwQzzhAUe+d5D/rj8R+wQE6C/uRZf4cyZyW
vrXV3jreXUxoyNjmap/ruWDA5yXrLGSjl927uRuqxCRD2lfSPR5MMjjwkMGFGL2xjtEUzSmZkwNj
42QgrvokF5RArJcQeyNq7GCvUj7dbYwHKTcQV9DTBkh0/yItQczTwHt2AwB+lUpXqiaz10m2419x
Emj58k5wZ0hb9HDnbp1KGa433hehWqGSBIdyW+JVnCZl95sKs+7kTiBZNSe6DWoXvcTZ0VQlvTZm
xK7ltaTscYaFts3plZM4qVP4HwnluNWMVZNtrq7Wo8vqDz73Q0UXaKtnPH8ZKlO0f97UD4ZgxDNW
/us8+fzdLqb6P+pJOZBWol5YK/hsumEe13EhHav48df5jFoA2IjOKh6spMD+hQmgRjzJwB2cYyFO
sX1E0AQV09iwWXL2EHjEjYMc/WUHYk7YqzGhF1OQmA72HLOLx5coNLqrrEOhRcGV2G996zh3UKi1
igIM6l6+tLShmaJccBKqNqK+fdCJIuRsk+Mke3r2LeUjhss0xySbjlxTsTa43m8CHNGV3L2PEbYT
bioqijTNSC1BL+etescGtBLKLDNVYxeWhnrM3gtJe1jf1cTznDneP5H4qux3II+YubgCx58Ccwx6
tuGLta1OYrKWbkzibIszzOcFqvHcuohaZqZsgrgtL9FhBaR3H/QCP5pJErb0jFDesSm2g0K6D1s8
dynU8+IyoTHCXrxw30zySZcKj8cTO9ckmMi7JKGB5q5PuSsqGiepLSODvvz638RPLvbuFNWcv9sc
SDhWxw9UasknVsArTIT8FGy4WAfNjZUayiNc5x3MmGTh12/k0nv8kjQe+aBPzrv5kWJhkA8jrvlh
Sp48jtaZRWT/1DLDpFkM66sZ6SARlOo6tc/r0p8JPqLodnWjABcsPp1MiodtGV8TE9F1+l41DIwW
vHsnJNCscNF1m1K7uZYonQOi2yFaxvoo8E9M45nfntw/ZYjp8mbSVJpfzx9n/qv01b66PXKDu0VK
ylHtUlLmF0wNJBsnfiNiV/UCQVfbIZTWXc90BLN8Le41jYZMB2fzb1u7A188j9LhdYHpEqeu5g+w
kjwQ+MmZ/CxK9Zknbdv8y8ACFAQEEivJtp59hNjVnoIB/jxTnD17eupU7oXzfh+7FflCUq+ZPh1n
0f0Tof8L7E8Hjoz9RbFdgdim+MtnPSlJSPF/lZAqBK2jhabSErIfxjkQQLadw7JO22m4jXhkVy/V
39MCcRVeJeGOvsE7H+as8bV/ghvnAMn2TUFkZQgYeJkm9DbVtdmmn4zuRUMTNNQad+LRQUVwSTxb
U7Jco4wgHupmOoFil/Uxuz4DbArvW6vwV0IsxQ+TFjWaH1LIolZsvPlXzAGGwoA1Xlk0niWyfAZZ
JwIgX+wBWaQSmhDVppTLTdMJ++1BLY19uqlFP7W1rPel88/IRiPeyVSesQQ/Ijxw2NInRVcileU3
hh7aIHX189KGjnRxt73+Q/bBcj/Yl7lxxZ2Q8wKIsTH6uuNVC20rYZXyZFDyy4Fw5SBAYiiam8gg
b2SsQIdiJg6p/Cwr7XqWKTvGOjsvFihqkxsMykIN5XpTEeBKhcm0V+SbeyQu0hX7hU4GNlYD05id
Ey5U6TFXjOp9PCJ/mx8pm9xD1gqZpq7RU7gXuhuZQbAxFJSYRoH14GJUzyMBi9ErV1gmJNv8Npdt
c4JRzlRE53e7uuF7FuDMixTR4aOoG2SOE2OyMUivbsqq0KrcWjHzGsJs7GuV5fbQkh+/hOCN0U3Q
vXp8gYWd+mFbMWPS9uQeHu1tfOcG9z4+Ld/Cn82p+ULGrQeNbUDMqFShMleg+qbMA0mg8GenT/O6
Ocd0Td03aDZhRLYUiJ25N1LiS5wiwBtHeuf5ouLTOlwKL4WOVQYKc7vmJ2ydL/JR0sr/XAB9H+1v
eGD3WRFKn/QjkFgafRKGlN/Y70ffDRyGW5p48Wn5cLUq3KRcQxV86mzmidPcxOSYzqEK55A5CIqm
6noDGYoJQNCQPXM8AfJK4cOld7iLsZZxIHliAy7KOIvHyEUcKLBXpZbmWLvzr+lihX3CI9XBc1Nv
eQTxkSJcs1bdQjZ+X//Sf1pZ5ivvpLYjGsPONcugQ81/GwhviNW8RQm/alT+ifEk09xA60NlFnjo
P/ZhtfkNo0guOUv+PK/wcyr/a/EzWhL11I54Y651PZ9MD7E8wZwssVCBA1cx9oEMICpkRHBdPBi8
8NxHuSD/X8Zb4BANzzlukIz5zzDEHfws05LHLOXb/EAqpPahdBWtMcQkC/jNCtVjJtz4e1onEL4A
Xm34G9P1skB5gHzzNyqCjxs7+9isbg1ykRPIaQDkYZzpTGTWdjKl359xW1nw6gFyjQYMW4yKAWpN
NkPfD7c4YkqsM7ohlvTy4boEVLDD7zo79ebX3L+R9xei+eYdEnrbvIu9IMrV7/0I31DawdGjogMG
hQIzPSv9hRRUcGImQWuZBYyhWZx9j48g6r9DXoe3tqerp+JC+zkRXOucHGl+pKgsiVZjEVd6pEHR
MMvDrdfDc3FJPG/LNYWTjiTNOHt6gpUXQpz/vqJZiaAXeP5/HE5ZmX8PM0o7H+9WDedlOdMVGlZc
VGmXPhBqrYFZQleUgr6QR94FgmBYtfVfUcNz7zp3mGIHsGZy5QvKAyo53lbKzymYIOdPvAs1+lHw
Mz+3eUp1OOGWV7muRt6RcoFfjXtT3dNa4RxTMvxmP0bsvP/keW7QbLFZacsuE8XWQ0yVu6JynMp8
OHgvJvryabZc2UoryYyzKBDetF1bBHTZMWbyoeZYZcgzApkm71HR+GPcaBVOHuc1kxYDxYomrh5g
ndWsEPWyxYur7R2/W3ek44e4Z2jywvigxcmBq2rISAg6bfuO4lQuxmrCI/nVkXFAfJGViEonvt9b
+/nDQe4amol4MG4jjNYH4TRHrBTfYK+HuYtGBEdljWB8OKV17ex2bdHdb8hfIZUqKS8TvH9kcVzF
PmqzYij1kP25pZzZmvtf0stkkEY6jzpQvTmWv1ruKrZjeTWIv7k2wnojEd+ya5j8Ye9xT+fRFstw
RF4AqSEojZiagk+h1YqQbFCC9kRO26SMra9zfYGdS07uhBh/eaechHke2mwjqV61gmLuuE+wXRyt
eTPdtKvxYiN/JBMB6Dt4NAY5OjyWGFkZUhyErS1sgrh2yvBbTBcH1cEyZrXg9HZyHkZFfxo56Nly
wGFPDOUaB5xACv9LC2VX4DpBc09UzTKgauGetMK6dj0JlGclgH2Wzksg53LRSw+I7Qd4dXW43ZIs
TxqGIUCzsIUIXEjeJ2Tet3BinNmdYrwSySeCACog5Wgg2QdnMVezaWCwxmpTOyRaDgut0kvL9hYZ
9wLZib7q89UzHpRSPx5Rj4eoxAyvydaV8X/nR1/7EsVBSET7d4SykLb+/22wtJVcOHtWVI9udc9V
AKlQ3wuii+Rs7ZbDKGO22S6i8ZSe85dDUSuou9PuFDeDYvWzpEBhSiSl79aRq4AmqwsTQXEpWIfG
u7Jg9tXEts7sC76Xs/AZTh1ITPLaHMGokwnQqORUyIAnbjSTNrlotrDMcmgf7ums/C3fABxDN7od
qx0vUUAM7nWTvvzWfUDNs6u/RVZy0y2esAy80jxn+xKeGz7IJeHBPLSgZcWsjYKOYWW1JsIMQdxk
9itWyplYVmyj/wRydftI0p2Qcu5+DxFYtM7Yz/LwCHNZmhtZu9dUavIZJ1aFBkpTIC2Y3kE8dGuI
tKKpXzAVr4CvvFq+yInuS9MhY5Vg86LF3u5G5ljX0aLwn0uJQMLMr5GMNEIEbgHJVWyxVa8duDKO
OnfEh2PD9uXy3p97Axh1BjtFIDoV4r9la08iH8tphzuXux/2H5n7vgdvzwQxYWSMoooQPvKli71D
cRWCivy4hAfbL0CuJ0XKqWLKh4Q1wD3Po86BqYac9Ip57cjtWYkFlQ/s35YJFwaiBPa6UsJKjTTg
5BtB4GyJJvZMTYjlBa4heuOEyP5DIFP/SZ9NfSc7j44GozzHFp5lp3ZDz0q7FG/ByN9RHbWm7rxZ
Sj77bbZZ9FOxgpheYrO2OM0BZMrOCE4GDulTroDLORmy6/3fBCtVcl62DcEl8F+shsAHVzUoD+ma
K8lga0Xd5mVAVERx0ykGeTyUuj7DscCWDqDEAnUDYn33t7Qqerk3Qd4wWnmgiIADXxxKXGTU9dbR
96g+WHySxY3dZuuHCHXQufIJIRrKHCsCbzDKpct/IarGubQpPHUuoRJ2rOnd3If8vlZIghhGYdLc
s1C7Bkltw7IIrxMuRyfYotKloXVVpEr7E6NwzWpeA1dswaDjdHm1aOvwwDwx2dDs8f0Te+aN39b6
+XRXRgl0FATMJGmyeaM1MGtJuvdl0pae6yW7dnusn+wHlCzqJAoKFLeDq5Zb+CKsqM04jC2ASD1M
HJoOpTI4aC8AG8aYk2H+WmrWR2F9fG3PMfkMVUUEs5vJZpIeQk21JgTO4uNjyNWNihmUQeT1yUvL
6b4fpPiCETzYkABkc2aO6VJ/iTFn/Ec1N2+6PVyvBvwwGhMP2vJwsb2UsA5QPoCP1ihSWvA22r05
Z+N5c0KMNXalhkwKsgJTiVl7E+Xf/LfJCK7G3U0bZu1GodcKPUlAxz58gOqd9ZjIZth+2cE9GQbd
zp9aNWx4PH6GSAspODCuSm9eHdaXdZ5nezBU88ji27EG5cbqvH6l902gU+zmBppb2tLxb24na5RB
B0UF8npSEPitPwPYRU6VWkZhgKkWhO1lhslq2AcGlgQGEKWZzVT+Derwu6NamiXAVu3LHtYxIF3a
oQykKYUs6hb+3R0i8bzp+XvrEwOsU91bmjRPCOAmHaNo+MFpndDqqeeWCKnn7W49vavhHxHVRp0T
NPtVqSnEOe3mP1cxy1VINDp9zYR8gCejs+IFHCjX9ohndQKR6gzRsWlB0eX81huItKMvuayO99I0
1/Vfx8ahGo1fAELJbGiBMWY9AQFGmxacWxl2/kKzPnpQz0QrWJe8msekKh4kNqfDl+eFZvD80HmR
Te94Ts0rwbeXmkIiBMHFjQj+055jXZRhr4cJuqa5+vntJRpLiHOdZUSukm4ztoHwRUyUeAnkvSwQ
c7hlMgH/3LWURex6vGdz0Rn7D3nlVtRW9PIW097RAoA5y4DFatyaMeKFUBMoDSyvNlxr4+qaxEx0
LTv+HqEpAm7evLEFA9oDto5XuYUfbLwdGYWFP9q1E+2P0DjKCHRl2Hm66buLwmglZg3nSAGZ1m3k
uA6JVyGUq+1a7cXB2cXqPB4WeNvHMX/k+m4sBOV/0ETCyzGGOD6ZiZqTac2t3BZMqaU+EkTsoc3H
MZdjNsu6lTk579C2TW+8aCap0Ru7rzXt2eXxzc0e0z4+vFONa8Rx1+DviI/VqqrgEhAIM4r6MZD3
hDq5m7LVApkn7gYIT5oYIS1/5sXVy/4OD6K6Kc8ZbG+hzhTcPlQdOlxr34yK+UBrvhx/A/4CL2Mu
gOGL4YFQRGPrxDSlreSjThTd0dAEjodMW4Ocx8RymzJZ+OgG5b2TchJgUuOVrRY5nRJSfzLelbIb
pX8vJYU7ngqxTyk5zPudyf645Dmq0dCAgcl4rLhEBizntC6YJJZhV/+s4Dvs45rRFQRqFTXlfndI
6D0PH8tP48rMdb/Ad0AjEWigKqrx6rAkvOSirUxE7qfkWQbuh09JK1FjVh5egTUroreU4OMfP5HZ
lA1GFCSfanolPO2ZDtwpepM6ZwEysJ34+/7bCjOIufV3IQhCK18x0kvyXkRr/r8vHdgrMvZrZUm8
CWasM2qbrhO2sbyKlOD1oGJfYGe+BRZEbu2DmB2B0pedDrzjF1evmztBwHWgcajhpchvGkE7eqoL
gYWrpcL22ymMuzkzvAfDN4DOjAivUUamf9v3+oHBe/R/uJbzsPBnGlRdAeTjSdXLnqFsHtvlX/oC
q07dc1z5V0fUqnSnuSr86UMKK1JjaXDb+0QNeHA2PUE5gfdNjZxKib99S08p8TKWEcqeHWYQr/N/
MjCNDO/usinAnueetGpNRBwF/2Rf/5FuRoeQRfv71tK6UBGavDwAdxDrBxsErhz/xVl2vUQG36g1
PG7UWX48BunHB0GxJJGlXTPQy8cMkSQF0ZqBGRKOQsJOG8bL28VHRXErUeq9oy8LpBrFqwPIiZEg
1qkJFjnCi3SVupZHJsEgASm8E6OfKekSdBz3G5MODErWV8sIZfOnXfbm4oLnKTdlWjTXarNY0Il5
fqOjw8JaGEgMjNjCcCKPTn3X5R9M3HbVsQ5vDj+z+gGXp8W4G5EaVoBQPxTk6rGYmB4Mhax9sII7
uod39MsBoZ4Qc/1oQTfZu8Tc9gYWHNzTHuWGPTKGev/34+K4UrEGO1KdEhYkSojbV3ooDCYW0vpj
m66ePv0MRixnTa/GEpsdFfIKHdZIbvcaAqDEjLlRrcJKZPHcAzKRuhjQbhks2Xf6Wnb8RL8Fc0KQ
wvf9vQExbJ7QWfxxBL45K3aw5l5WuR98Cr9ZPhuPvMaLEZIIHR68XE/gu7jl1ScIOQKW4vOuvjpO
CIvgZT04dKDff3lc+9XwY275Mq7qPxkboKeVzu1tFgNtfp5KXMcEktGmmxtDrhiT7F27FdlbiZzn
i9uaWEB8WRM3nQR40d4hmAOJjdBTPZsh8rHsWvGG98cWc9b6hXgnbVmaTTskTXBr7ct2cKMEWe/r
H1PtBkSdj3rewx8ruUSS9aGObAIXbrc1LtoOj2O6+lsjJYSheTSZYiTo9TRlo3fuUpoB4OhP4oZc
wwNcxDEBytd7crjTanzmfRkRoiwLZxQz0C6reCsdR/uRILfc+i08lUdjxCIlxUFYIWrKGTRJSdTj
2d+ZUZaR4q2oaMSYTBWUgcs3no6Dc31ujnGBmYBON9dohX2jSu7BrfAxP2nbf7HrBWJEbgT6X4HW
2NS/VL1RqzXawrheHCo34NKLRniMeXfIDd3Gjfm0XS2eJnnBes8xw1x/IcTprxIotJfdozDGxxYC
T7idMqVEryO+GqIbZZ7GV4+AeYTqpl2ShpB6Bresp2QMsXrYh4MyEc/1JScPwPbjWpWCzuP5ywwF
/fI16ZeKU9f5Qy7/nxvqEk9pVVfvmwFbLszgKMhM55fruLLdqE9CiYUU71fLrU/SFmkqMCW3Sciy
fA+xuImNhxvAzBnRUJAxZnhKLfAn0+XdD29yBPSR+h5YwrTcIHKhLeBqKDdLatg7cLdATaek4fD0
4MW3zGPQ0I6oFy76OvuofKoKR4T95cH2MTVYSVSxSRHg4mmJY9JT89f3xMYMg3c/V12AUDDjbJnK
c9tte3KgFGlskc3118K1rHiSuDPmeSSjRbJgJsjtR5hm6zxgi6Shm+cTMVkiPHyzRfgR6Bsjk30t
KTk/DjlsM9E1utYMt5tR9jfhdavfpFyhVUgEW+bRP3CQVVpT7snZBKhMB+LuJsxca/OUevsQMF4J
HAqI0PiMetSoUa2+yPdGD3JM+h5U7d3fA9iyTZq9bHugV0MZkTxwE4RdYc0Dhyi15jsdV75RbRT1
S1evKgrwmzqtJ93utMmfd2aUIn3mzq0sn9rI9LJ0t1BvzawxpsNiBX//nXIGwWz5ROhUGkJYI2Tn
MuJcOzxRZU2YzQ/0id2omTxWS2JJ9vTBiPbG1Cl7nnkZUcD8TfGGyiOKgTDcvaABIhFAW1C5lj2M
9BjmaRJ0i6ixPsVYURevQuHfF0sJToLnPRlevmRxOpL5nKeUSsKIz9jPdu2nvrv/L4jXhjAcx6b7
QOZNXrwIIIZVEe6+Qx6V76ux/ffeu5C3QfEDC8Ydd5Y0DzlrcvhfUKuBfn6e8ci9CGxzrxBnfMQM
kxrf6xPH5AAj2+3FHyt8DlJZPBcx8yTNJsDjNgYGhuwvWWaiCprP8RkUzoTAyHHDwEDbaNjlNhhM
KWoVmZy35D+kszzr1w4bfR1mNru9mRepY1wTj/aTGgffNd/pjR2oGCKfD9Ndia76BAK71bjYowIs
axoK9J3UjCoTxEiGCWziB8B6S+FnUW0qMVAJna1UzUVjZ3IcAUAL6FWphVVEhajqZqqjM9XBhCY9
5BINGxdwTgU/6zDTffW951J0D59B+4EQy9/98bzNnYN59pThN2W68JckeU50Jwa7ywuUNdjKawSM
QqP4AXZH80lTCHayRLvyVf8Vmm8jvsqQANjQ0Xr+v0dePVVZS71KE+wlrK6LcdSr7ZyqUNDff9HF
l4mgtKLsDamotBwzT3fSpp8lapePagbC0twWM7hiKavR/YyEc/xkWqAso8eL16Kdu8oKDAPQG/3w
Ds1yGMcTW7eM9HpFyo770jR6XpyCHicRO02KfKK/40a0AXzGPOJRnjIODscH/QlxSntplaWxhD5E
b59XqujiL3fk575OGozP7+61F2CAhge7tPa2MVhRxhUFdK4XjgolUWHu2FIS4/12KGAShIESIX4w
sje/OHpM45idqkMTQYQA/Tp1BtBCXPbc81Alsruwx66agFgEX9qh4rjlqBkx33YDYlstNMrIXkBD
MpgO+2C/atjNyxOcNDgrDtMmSwkjUkW9wNO/VJ/1nXC6CQewXWqPN8uWYab/3c6vSZVv7t/WtGcj
WG1BG+r22qyge8yuPNYifT7MeB9ewHalGAHx339ZaS9EmZ8rJjhcRUaQrQZH4ssu71SN+t8gKxZE
VvB2ARcByzPXez2+MY+UvcSPV3sek1w7jlu+UnDjrF41sh5/tdWWg1K2JcWCmTuqQkm+OsIgD21c
7MYHoa0POJwViZQtVp6y5S+RPXMw7otxIybvhpBjbSCFJ6Y1nMT2iDsFcZmXt9u76d3Yg+RZtTMq
X9Wd4bOmzI7f71F7Fltk+G9x7Du1TVAdwwMZ4nV0pzwn3ONXqlbmeiKpDyLB8KJMvHPJQxbOVdck
juyhzavLJRHNzQt47SVqagy1TCdHatC+ioMYo5PA50t4n+jutCXefzC6AWfqWekiGf+GR0mLwxNm
BL8gt77Wo5v/ZsB4zIo9GVu/jMKTYE1qdKhsOq/IlWdRT5P/hRsAesXPUrqNB9F9VUgZWEl9auR8
dKUo71/NVLLpDtOfI6J7p4fNoiCAiPL4TYExEu1ORGnhWIpk+x4xSswIbqQWFgPk2/ZymO9SxmZl
qzk8AMZJLcrpQtrCosycFVpgdWWVW1TcsC5eRzP6ren4eE8aP6nFEQ56AhvYevjn2HhS/BUtqaGN
nkpek1UOMTG5guK5XZjpIou0t5KQuevLmSabiu31wmSIaTPHUssjz43x6BPvCbzWG6M94Hha0l4N
4R6Hd6AdMjAufozPmlYbA/bXi+nLyXPNuonD4BRoF4J05INhm9RyPWnlo0rz4Iwv3i4xUoIDLIaN
nJlczUDOJABYSq7iY7rA8Gv2HxB78bav2zzbZvu9w5thmc6MBnAlxf02cPnvQJCxFQz93EMjta4n
9deYY7xB/yumefGx0HRFs2FJ836Gwu1uCqTyDIPuMXOS6LYJwcyHG18AUH2FK3D/CtVkRkJMsEEO
h8FuqnGzAWZnvPzvQ+vrnzD+ff30zkg2OlPYlxCImbyYP2Ob+cdls/z7hHN9f1mCQSoJeAtDQNuY
j0wrejRa4DZZzHi70XaBHlvB+Kbd0ICXHUQq2tpTo2bfhz/f4r80aT9+93Zos0DnJSCMUTsObipR
/SafWj71eu8gbpht62jPyTPvELL4k0igswl7176++bQfOQ15CuefkJNzh1cEqFtDF3O08aSMWHic
kbrDilc0AIi2Z+fCbBIXRY1yDGg9GJXLQdXZgQ3RoIx32QWNpbKvCyFRPYsNfFe9fOHTSXgFDzvR
lc9g1KUHdHawCdGv/YyO6xp1dGY0GYlalJI3DlNtRP48gtvsjOSm9Z23XiVoCqs49hhrvr1Szfbu
5Q35qs3y/A7CKgiO65DPZfhMOQsiXomnl0972afJQ0W6ZJgr4AQZA8LSxtvfDz87woqNI2qzclj5
NJ+fOTl0gOvvpQbdV7bVglBSvy7PqKnX9ZGu5tr2QnAdFTdyAWAaKIhDGaYsszkY4Rj9esxc8MkP
Bck/bZA3sPYkGODnk6cJ+qIu3dQapGtO27dzXgI0p5FB2+2rm9kGatIxbHzM8CKpWXkV3PmO+GNx
2j+LsHGqlpyaDZFW3b0N8bXLPhfmsnGAVOLuZysMT4/5JryXwptySoSiKT/uzZ3EJmMhBH/ey/Ht
v2u47TN/VFQgky+gZTxsQc9lR0wnpL1YMr+cI3YzX+hlP8yh27KbgHzzG0e5BRGHEOx7vpJvmD2G
Y2p7/Q5v2c3ofPznp1XvJCvywdTstX3la4VWHw4y6jI8UhN0OdB6b9DM68InbouU3MLz1O6yS8TG
bNk9cZtzp1yGYbDuM4aQ08jl93m4MEd8XKcGq6mrqu1Aiwo+NLj/4DgylVVvpRsMUMK/wPEwZk5A
gZG2TxP7V+aSN1zLk0SWHSN7VxAeNNi8adZzUgyw3DmbtQFJ7oDg9uoDJR+kAtk28eITcowc2YLw
YAG3oi5rqI8OC/fPmj+gJk1A8QTGxLd5KjVV7zeZj+0qFFil/eF1HeipYDbckvWKFBC0nPaIVTbP
kFOlyz2nFzhpDNiNA5DQjctnt88Bz6Te9A1bDO0ppXYgtLcnKq4Bx7yE4M7Z4M1wt5KQRPI0d1SJ
/RA5kwx1vAj9ytUqOAl2TrWN1Rs1hfJ+cJi9QHWMxNP5UFL67BT/hH6feXCI9TULWCXrPsrUFQV6
Wv9cNBhIBekHjhnuT4AFE3fPFzbftVaZ6uqqMB/LhU0gzeEP77daCWJPTYYJVaUF6+214DgMlS0j
gy3lb0Z8354Z6xUsBZGSu/60CszD/51t5eqkfkkmGeNFchoU4auaZPGr4OuVfCxgD234h936CChh
TSiQKnW+f3oTapTIQDXMsZvONt1f1MQs7PHo7/RTQXYdgPi2S/4oVhkZFvFJ1O/hAiWWmaM3fOKN
5H4nLZFzJnmUf9G/xWZM3lThzc99ugO/ziK5dVyOl2SCO8gcefziNQG9YEJo5O0pVAi5xQdyw/gI
3Ce322cImPZmCbEJtH+mBg9jpbrecNbkWWJ1MhLtz+aX//FIi370nGyMawsqUREqTGiXeQZOHkgx
FlOVaKZTsf5O4nIwUlHd27ILsbVcLc7tGRziXZjG1uWSakiSvwItYiqK09TBeKvyKAS6+/+DtAt1
x82gMsgHgYJQPxE0TxBh14RYHQIPtw5InkguF+mw54UtDwJ4EXiFCaMCitkljt4l8KeXq444JxT+
SLI1wo3Tt7JtVQPtL19+G3AsmtQVIjXeSz9aLdN7mquyoBC5DYsEm2cM6+RIgDexqgAz1ncmla6r
a6rVuBbtOdCmBTLRn3YWQnNjMhHgNeXMrVHDfzw0/PQoFxfNmpxUYVKuy/tNjco5+Y+Uw1e3SKWS
Oj4QHJ5nI7O3E+8fL2HEK/xcHPRcrIp81AFvQxaP3mscmSbjpvpRXxK/06KvpiDSs/8vArvWpOnd
8t1Ruf43niCcNqdNeiIGgu6mxko2mBVelrnKppI5L8yapxNM3Evk+EO/t7Zu0FZMZOD1cVLTYN/o
6qnheXZUA1PbvvVQKIl/oA902EdC7Pa0J2zuEwStqnmDmohHvxVJpek/UKUE3nDbgZIDspGw8Fuc
ErF9PiL/gwdQbJ5CEIKHbE76joPBAPp/hPUVGhJE+SDgRypmUu8FGsBSnSy+JnNadiE//U4koK6y
MKrf09ZlDQLYUzoTf0EdDOSxGXzuu6ejD9OK9vLu1kIUDmehBuybkMsRLmpWncetg3XXAcrQJu5c
ssAxCUmRoC6P3/4QyItUMBihx7aur2oVciqyhBGd2QZuR8pk87Faa+MhdbUPzuq3LA85x9KDqqYZ
y+YXQ9fk4WKugbUZGSiQKeCb3E6MMBCllbeR4qFi3enoFbgMTacrH5/N+JMEoZqw3lNv78cqZx04
J8ym9UBrZdwkN3HWmlFncL8Px+gQz7nGL2cKtsaDvYzPU/svyqbFEjdJ4Q8IKN/h1V+mco4oTJGU
hsHCp2++zXa/cTWAqS+tgrnb4Fzrzo64PdCTaQtLVqmFow71bNL5/hLKJbLb2vfQo6Gk6gZkON4T
MKBXFnm3jn1jh4v771idu02ZXkvnqkoNZlsQmmmhc1WNLltze1tRkCxXdjOEJm1MYQCBWW0vgLAb
1f3FJRzbw1oPLy8gvyjCAG7th+nxEiVqqtPAMzqqvgrOzh4u6+YNeTvw/TjCfQ+7rLjay6Q90/Nn
doQy0nhMJKWMkw2zzzMIPfNy2m5rJYdexo5eDnhH9HmWIgYTfOJNPhu7a+nETJsDnzOViQvMEKkc
0b5OC+ler72mni1yjMZgqBk6APmt88rnjS2T5lRKbsP9ZINMttd7MOS2ZHQQDxACPahSSuBMRtWN
cxfolo78uyNBHqt9p2g6KxtUGrW7fGAX46UTPgkSIuTirl2xvuwPIrdvu3TlW5TemMLdvn57NluB
DI7s6qe+dnPayKmxucEJWtixCwbuSVkmQ9lRM8F7ol/72XiAz7DoF1AYq5k1DDL3pbQFJ2fHM/UJ
Ogc7TVX1AZzw0BFznBCHPvAAJBf3sziDuTUzqyx6yA0HmLxcZqLoA3NUdS65P8xY/vfepGy64TO/
Gxc9tqLUuDPoHQDdpAguGT2rUCHezsQ5nSiDFyuJ5426U/rh1SwIx6EuVeo2YI1xir+zEAt4UGky
fcXSe4zNCz3oNz9Gdx1FMrDU3i7Wiva6pX/Eh5qHGzKF0YpQLYccM085RS0VS3HcJJldeV1dWwXG
EjuX7vhHSCS8L8jA820tnaQm1E8YswEFHgwoYDHGDSBsFB/eInf71aURoyWgY001TOgOA9jz7qTl
hCCuiTfNXsAEFMiMBoLkc1DXXtKNWrePJLYFlyG1QDu9GXZEWkgRmMOfMs3jvctvtZ2GqQVy07lz
yQbT1ROAuKVz1P1mL/CUy1FroiOeK6hVmdvM28GgCbknITIAGt9iEbnVq7qyXV1CEhkBod97mnpi
cOrAhYlCbcbtDIE+9UeCrcWSIbQKUL0Xe1PXUUFQJDEC8weG+pmTmcpak3xAv8btEliXt9xnlBr3
cDgmWyg1muzgSw7Dr7wzkkTTjHpyxiQqbYtPlhEWBMnnygKh5vwwBulWw/9W3Fe470cVa7bUkUNw
1BVbfUC8A6+dlszsDli+jPJCQ1zEqBUSNobonpSktDmZ6JxdVGmTvXQS9kxcPqHGjslWtmRxsIAA
ErdtXy7FdwjYBAsQsEsiDR22iunFlql/0zfskD4frq/A1sKbDyDwMLkwqzKfzeYO9WCfA2tEIlHd
IpxKiYky25+uiabqHP/tYX0tzwWqHOr6a6TjTrCYAND7+OriPCnjpMXvYefpIK/LLlyqkDNXsfyU
zZ3cIx/ph+DS2Wvm4UI6BkaBW6lgK0R+mDSWCymIApddhHnU62K3FfLD1siH+TBJIILp2ZnS28FP
7EASHW+TkEXq5jDpNK0Iu5OikPdvzK4NBhTpnOP4NVFyi9ZaY2MF2da2abMKdPhJd7gdBjs94E7v
/g5/T9o+qnPTrM60H3pE8fsiCwOX80gFdRh1qcxUTAs5dvIMQ26v8iq8KV2ohZTI82x0KZm2LPxo
upIr13vDYknVPGoFTsdB3/BS+mbpX+EI9YRUl0dD4TEZSX4wc0/F4KfbXL4ke/w7PT6xQG9UVgz8
cxv7iHxyXYFpzDaIynzazUR2s0KD0eMKppu3lqWNWiFzDo5g3LxnLg2/gQiC8QI6n+8BS7XjQC/8
00UTvmRIfOD4Dz04gHUsLV3rRbdV+g/ebryrN4Th4zw1Ph6c2Zceu7k+3fy+7y54cop9Nakz4N0D
aQxIovvYihcAMstiuNi75eqdl7BzMtVzlRNQIUO9mLTcl0HCEo2JcdFRx1I8rE/4wdsj6/2waB+b
s+DGeGIF0gy0f2jfKfHtL9m0cqf1okfhQIiZ67LXe47kSgvLrbFjRW8SCmj4s20jjEC8hX34DUva
p2IjOtPVlolfgotIR5uZnwdjH0hrg3p33b8G098WUCXiNHuFn4UWAbeNvjFfLAz3ypty/qaqPPmf
VY4z8xq/hnB1y2PCI26VXqH/YptHciLXEtN13fPJ1g+NXhbqA8M3KY4niep4NwubCR6ea8p+8U8k
iPKGHhJgcM2puto9hILjeG+KAHIH07k7j0Pb7uPRn4vfdEL9gAWCDIxsa6EYIaWZrIbI4Z00KCmg
uUz7XQIXmWXJwBMeAQojYV3OVHb5DwC8jQ0AjSCQVJZzvB1f/CCqs1Go3gpOE+6Za4V2/EtXPA46
T/4tG8P6ePs4bP7rQmJ1tbWqeGV9tMlwDlAfvmPNxetCoxhuxa3Q2Wvm0mm7/YgSadZZo2z81D6k
5I0K6FSuHhUwEPAfx37FuncBE0ni4KrQictNqzLEY6U4MozoLdS8JZ0CP03qgzb5GALdQC+lO14D
cHeRNzsuEMrpNewiRhQtHGhLkhNl4bav7ys5/FHk0bkfYpP8V/tN5SDqPRQOqojii+kueICxDdUA
nAb0Fb26dKWnR7H0y+oJGStv6QE4jgYLoxDujjTE/ArDQlZJxevEurGjXN+Fr/rrerd5lYNRGeoU
kkeng4N45mSPBLa6YIm6EYgkXF2YOWGMMnH+os7MFSKDlrcFRLSjNQIipzHeozbBqMFAltaSIBHv
OUwMkRaDSB6l4F2JlLo0g0AqaI3S65HQxFmNoGnbKOuJsz5R9ZpDCnd0OdFq2v9O/EPHL4Q84rK7
L2IXKWQDqipourJvtVHNa+ya9ZktWFw3U/S8Hke+TJeup/E1Sj1Kn3/oxnJ/m2ceL8F1F2QyBzqk
hl2cGvXxdriqyPGnu9/dpAKZpbphAjVZjCFYEJLts6goh8Umtu7+FR99szCJ9/biyw/iC8N2mfgs
hMCfQMxPjh27b0RuD0j/WkPHGrOv8v+8iMvGmKl42waQJE3f5QDk+4NRJ+5BSrNO/yFSJdOgseKA
IvkIodDkf72DgVgc7QU2HlwLlcmvqSyydb+Iixvg4bXNRczIFLGspMYKIU7FOuPAVhpQ5UN+EGJ6
4aTLeBa9bj7Acv2dRLUiAPwBQwYQ5N3aQAKouMpw4cPsVTl+JRlhYvy5hjYfCQ/9Y46arbBHhAW2
0LBTxF5wcwUu1+os6B1fBYa0PG0yZjOaZmWGkskPSmkREv70uEOlTmdoeJcHNgJjpKYEOyoSyzjs
jbVcWs2QFHAtsI05M8Xl6/AoeyJldNKFdNnD/wjgto1y58Toc9UtCotB1z8ZmeFj+oeqy6Mog9kW
NpzEia6mkOaeUuRLuApHc3xlYKw7AH+iapxLNv4JkPbqJ+gyB+Hsa2wkxsXZUt7C2JW/0GORk20Y
V9QvIllL3z7q5i0q5u6Af33S2A3oqm6C6kwKT3Z3AEd0VP2d2db5pr7ubMw0rQzArsbphQopcXwn
e4dJmnMtafdgmUApHLjqbMbP54AhN9OEOUzEqp1rrHPtvS6a8JqkiAudrRumCGyrZZ/Eemz+RMz5
BlUUxff/SzUko/WbKt7wiw+Za3xc50c8Ci6+0MQzWOPAnW1rIfvaW8zWnQMOTIzs0Y8BYE36mEZR
aLoCjkKalt449m1cCV71dGdihhYh8FCZsCSlEoaYmWZFCOeWXjd3s+Jt/AcH78/hr7YnK0ioSL7g
Y/I9LuGmCTPiPRJ1Hznpme22o51t3I50MjQE4XVCuxugYpUl9Fx2F5sP8UQeUdWMNyTx0xon0RSB
BcJ2JzrAKfOCnj3+iwQ8AbiyGnNfUGxlpbN7VsOfC7We6NdJkS/h7NHkBAL41IVegvyQQTDdVJKl
7Pu989ql0os9GYoBvm8EBpQEUVUjSXdR2gdtOI+Fi4gaj2+NYPiix6GdJc57yR/LV0zYPRnZ7RKZ
mM58dWvdNGs3ctopchKzks5KltjRMU1klUog/0QX+cVs+lbjkSgbhHMd/4aBIndRI4HAuqLGmT+s
w51G6SbpI0wrt38xKAos86MdPwD2ZNpGRoKykInO8ZFpeRIoIev7PiSByYagoTBz/aeZy2ZvUCz0
sshVdGk1i0z7f5LTYTG5TkhElHYX6UmVvaSo37zk6TC03/IeMRrKNPu3AG1Io/RjI8Jc77UdXgNw
p0hPSuBRPsEt35F0tgTswLA9o16QPtzqiINorpxt1GmCM7OElwxBwrAA9uHkEshNacZsE6ckhTpm
PuheBV89BqCE0/IaOnBWXtkdlsdeDn/hTframa6pOHxNiDcgVnYVJlwkIPnSkoZuwUDT5xV/239A
4O/j+w/sExfxY4ppUqGxIn5ywucFwGtdR16xB3K95WUffH/8yC30fWUWNK0daRVNZcBs9+NacNbO
R28twkfaNeeuc7acv/GBXoZZ65op4S7vvDomflXWZOczyCAJmukev6q1K9XeV7sEsrhn3o0UfW/9
FSbFuDkShb1sv0wtb4p0bqjDmHDIRcmPU8jqvePvgQb3Y6Ae6mNwoTIoWDiX88qXK8fWPZHxtwFa
SmtAfc4JvvVp11Ktmz9d6TpFOFbJ83ZjCRTBcTkWNoEnXtc1ZyzOEf7uYn7u8m2bRxJNVlHcQwpq
yCjXxD1+XDHg2B8Yzyn8aFmnsVnQa/lysI5YhEKW2KC86NbzCQbVkj+jx4KIVc8fQFeGGZctiWyl
aLEQJTDcskQCwSWG2D1Uv6BeHiUxcvymvpbL5+BtwOIyhCc/7MyNVC98I8DUSNV2HbcMOyH0Ro2e
rk8v0naARD64uAC27yChfTwT66AoAQkORsbfvHXd59H8dvtjdJ10EAjt/60qeGqMd9T+Gs7u9rcD
ZZ1C1zLoCYfrDLCdkg+JbWArpKp2N4TmDhCae2U+xDtzWaYOq1wwmVSM/L7/QLOcFDg7mht6aW+D
5VZi8BIa9Vau//4qi2lWhAGLOWPkUlM8QF6/5M+B72Bw/645cQ6NU89/Y1txhdqIbpwpAEnAiRsr
AetRCLX9cmYQ40lNXlnknqQCoqm3PSxmm91lZB/HUI7s1VtCuHvghLc19Nd6230A818m4zz8JjKX
KgXznTjLn2pruWNN+A8htz8nInx0bngXz1uGambeymHGkWXZxOdwDvypxZa3dMaDmCexilMhLFOz
auc7YqpNUT7l7PmkfI8IWf6hABz0RdHt6KpocAfD4z8Or/FXdtULTJuqNrn6UV/laGAfBJ4HpcID
qn0MWdhZVR6TOkk2W+q4jeMgULThwOrMAqhCjhbWPwDISTYo+podzj+ZrVMUBk58UhxDNt6y6IPD
eO7D09BofmekiAtk9C2dBjizqsFtlqMfWW4g+N0tDw/Y28G/8hUZjOA6vmGV4Er+DSe6ppsiRryi
aCOqqAmnAjGsVL+nz1PHrmitzgOOi15eMk5ay71ST6ahOlHw/aDtM3t7w2+SWI0Kqab3YVV+3tBk
/pRdhTvX/soPFAq3VcnfD3pBqQrscvGZDOaeaE4+UsTeeCDPiTnenX9YFEdO+0RwoN4BIMC57LVy
jxXMjci8rBuUcH6wkZNaXq6ecIwaHo1BpJDm8P5cvtP8aC4e0KZSA432YQQ/ksvHKCvduVCTvMet
Dxpx868X63+CkgdA1LYNu9B5J0Gi9xa68JazU100fU7VQBPa9magxOwdmv3CX9k99CgfUZrz0sDF
Q1TjpjtiwBO+INmwpvvfjVHor6NQg7H9hy2cmhRqZbBuDvkI/09ycqIob49syKzLeBwbvq2Ea9rm
TOBXZYNwTIHpBv9p3USB/e2tAoEHjRGxE//PIOS3EKULyV6Da0IAKAcnPMmvGpy5BOZbdwCSr+PG
vkNgW072VTij2ype9OVpiFvhDIhU76IZwOa5vsiJ1v5jn06K9edFl2VRamGLAPYdFQ+7eWVazXzj
M6hGaLCNTIuN/S4x9RxytF6riE1Z8+kJRPGL6pqxCAXIAMdAEMymZAsQFEjFFlRKJPJY5bMj5slk
nhIGBbpcsLqnh68Bl10MProK31w/YN71bD493E7eszJwaykM6ZEO3HvEqjm50sYz8MK6p5hNRWVU
E/r/I9WG/U0T/tGfCg0UrfYFMBfQfqmyMwQPZeZETMAcLbg+U43cWUWU1o4A7Kt5m4wzx12ON/vV
vr7PsIQxmuvPM4VEUAwAV8OXyBJKxW1fsp+Z9C/Cp84CkkC+veN3kkByROx2IG9jDYMR55tPDNcL
LeL71SW0kLeyUIrLA3NZb+62augT7xrWND+i15RMJ2z/kd8uJRs0RdOorjPzrdsKBxrt0Mb0LPRc
fDL2xy6ozOCNkvMT+6NoniypVrJ8pxR7n2n9bgPcf6PupJNVQKrrIrYmfkm0uOR16/UJJJeAQfx0
+foY4pHuwiy+41m7TuobBHRDZm7/mCgPbY+xrUw1fY91Iw8PCQKPpBSWytHaDDQDY/SMOE32Iain
W7F/xET/tJMCLBto5v710ZdonDml2muEk2aSDBBAauAaEHqA2dTUQjTMqIhA6bwJH0f1QIW/fo/Y
HkiUBxAAGhlkmP84gPGa+fbTkbnviTo6U/YiGmZLb82tL+ytHJUs513QyZo0gMbDeDp5zlAw4Mkn
yljV2JsTT4Q9fXX+VKz3+7K5Zm9gFSQP39apWoJl+hWaISDr0GTaQtheRZrTkXFX9/c7B1l9RomZ
CYHygZVHEOKpOARoJgIMkCBCMUWUN68GN8Fylb0CKRNTUqCMt42w3pO1hy9WkefCYyhgTTCVssNt
H1hgvEuZ74IgBeoXPvo2DXNzsf9/FAeYFZ8etYJhGmh1f+k0eRL2zN6rPKDrfhWcn30HLUNhEX+G
S3IXI5h5nSnsOk5gBAcJiRuQS/RngWk5WLFdhcPlYvqFYjTmoOFwMHwdWHefqOAM7YQgJudr62r4
6fhLDZnztdocwyrs9co9BnN5r7LRZ6oJkP380IlKmd7AQcdCMo7wkwY6zVJMprtfgwS3q70ozcx3
2RGQI6cvzJaytLxJro3RYRKGcMznXDNgiwwEZa2bXWgKDhocg2i2YLkjAE1YSbIQisUnY0o4HnWE
sBdrUuJpPUWOpJZYJeTLfO5bnr+0tAWaKaMC4/xg19Kenj9L3EZUJ0wnGdUCnmzWO7jXSyHa+Ste
vFr57k//IveHgCgsS+MHu6SqbzD0DmyI3qi4tYqgur3kAgtmIxIvRheLUA3ztmCTOS+Dsnd0tvW5
KTW7cp0CIyEZmqo8TbYjvnIg3+3fUDwV3aBnjAkWYmiv4MAQo/xyJ7f0pK+BTIRU9K6W2DJ38U/u
kFE9/a7B+jzdxjJag8Hi+HHGThatQCzZ7skH92QdrJRk3RD1PSqNCUOCoBWW5d7p2fOSL/XqLwTU
do08PxVF1rvLnKRP+OXYcccP6owN1Ep3k+gePA3NzDDWfkYf33uKiLYm7iqqJtqoBdGwXD42qrGe
7K3+rllgEEj/s+ddCrb+ctZvZZsa1ZVBu1qUf9ZKJzYRABLbteTFZpsieF4rWzXLbQy4kK/LDulI
BNNWrvqZM5e2puNLNrI1MGbqP+KeCxeCpaXslGkJt/Pa7BPGViYSSNxETQA0yLfZqUt7xn6qIBrK
RFDVFs9x5ngdk0DCGPDsCixmAf4oU2LgI+8JXFFD5nEG5C9EQ/0fqUchARYOGKXeh9QuXALDA98q
kLOabbwlqdpK9w+y0UGx97jEUblPvIriqYwEAFdmTRuNN0FZyufYrGv2ayPj/EX8LVelmhoP9gln
W5jTnPvIbHgQfG4ElmfuNHFmFgYVCRRN0M+4h4rM3AnLZHBX/enTNRmRL2euvinHpU1vdcXawAcI
BgwChqOL+VG3RR9ITlV3O2rFc6M4etZ2H/hA2f+oHOwgNJ2KREm1WVjCwqxovaoJc7dVA9lDRUge
5E4s8eRfLTwQ8/6ua5pLUN1/OAVVKnuxMatfb0KJb2RbiWY0YHU5TPt5eht4n8D63rFz+OkOTTnX
sblZAFp0K+mBU2jO3brvGpYdrDymle8owIzEIsvZbVJ/KhxCN5QfFJvMnG0g8i4dv/uhBrVbgV1F
FgSD6ZWZ0Xd20LESjlTuFVF5OaoLYtsGbRhZS8sbuyQ4TFBa4sytCJ7gDfrLC8deaT+ezntFwF8f
3h72yN/j3QYR60qiWHbI7/hmsx1U4Nf69PVLLohZYwAKuP4z5ZhLcnxAaG9rOS/XH+XphMvREIoy
ngEn09V0Sq86LmWSVGsBydow7wpw5BmJU5BGTVVwBrzUnIlA0+kj5DUHbynMf6LKJ92ZwyvGUeo6
/nFG+2h91q+BOomYnHS4rpBecAoOtuOX7foxQ8Y4ouiAm2jLoH3Y3KrLmF/16F6hvdmMRt+2vV0+
f1a0z5SD7j+oSr8EidKRn7ES7Vi85iVSodkq5iiyaLHkxp52uufHzY1iYJki66eIAJLDVITATBiN
JISPyEOoMaTCsgwjFdQDYbYrgan9DPsO5Ty+3QfAh/PhjvW0uMgiKBWogR8TIfg/Y5z0UxYutKVw
+9OW59vE0ZFmIbExHx5hKW1JkjfFdeAn4bqfSusEKudlFUf3+2XGMA7qtxl/7BF9zIceYUHBtAib
cxr/fZUeRntqL0KjsFcTgH+ZIZ9GA6u7q/iJBgiwQbqLCzHPXTvzKgjXnpBBcWUHMt99kFee7isc
Oh60GNsqc4tQnNOJtYzqCyf0qs/G/MMXT7mugjd9nPh3wPIL9AwuirIFE79XyLzvcP0CrEhbL8zm
7Sj3dAG139EmwHijwzoYS4OVKlvpGOPnneTM/q55gmJ81aFwN+R79HszGyhDXVWprZcS/SH1fAvW
CeI+huB4K1hnEBpYYGp9S30rk+SAM5fGk5SjX5kyDt1i0H6xEPZFlhTos7HRusZJjKJy3l7F8eCs
cXVC/FxGmPJfeTGFCMQXR9gtneKnMTX1sc4TqzTvEZ+NYq2RU1rCBed7gbEFgeWyXjcSMIlP8OnJ
jiiUeadvBjWo5l+sJ/FEhJ9dS/0R6VwmjH1KptsKjk2tG+xIEERRWUTbINEkLbac9IB5tOZuc2M5
PkA8dSkPIijW/MYdIvl3JQaiuAzAUFyWid8OG+ya+gSI9kGrg/lRkILR6ALOwnqH/+sz+dy3tyo+
zB1gP+MV39ilzk3eAH7s+OruJZ4Z8fSwA34UVAIwNR9FV+m853tepNtMJoLBTotR4HDOs6e+7hBN
Zpuprc7brNzLbMiftedifU7q5z9C7fPY0OWFv5rdGMkt6zUuhQo/hlybCWKO8pe5xeF0DZGWi31N
EncXJMTa1ibsUSOLWOD+MJLYbkZk5HuO3wM2vvnTuHek7hGMBJUpo/d232qogIYodxkjD+xMt8/L
PAFMmiiKYefC3XnxPFXuDmSPMZuEkG4vLYTpAJSgvdbyk+TUdhGk2A/L+w5sqPZ28ZvVEXLwXz+6
1cIjPjGUV4K1Ipx2jOJzdMin+XAQSSd9s1chSGkSkjiwNMqsqgc8F2z6C6I20b82CiiBUwEWW6+5
iHg6LXnYN67zTYstkEvXDo8pRSZ0adeqMlPqRNfTkVOI3mYKVtcht9YsBrCQOKsFr/bsy5Kf/uTj
S9YZrcpoxT/BgHDFgDHLQ7R3LE8V3pLRjhHiOD9N3H0q8kwC7Fgt8eqn0mKaMw24/nupBzi/WAXW
T/UreyBV6n6ZKHruoYn8Yd0skKNZ252sMo50cUU+Qe6ls2CB1+YRqoElzAHlGi6O5SDyQKIjgMrQ
eAGGnVxk8FDmv9PIOt488HyAhol6lssg7hSSudpyz6/3KkdQNDliazFPK+IlrHKJmzJQhVINXlU5
J8IL7mhY6LPGIBaQBkc+fqrS0njGlqlrmi2/SJDtlXl5i+lXhudMVeW68kjeTBM5boATHquJGyU/
ypSFRH/SM1G7IhZdtLSKIWxiq4gM+me70rMFyzRh9dpCnnIBxIogmIY/hXwgZaQ1rpy3WPJrX4DO
ft/supYbxtmsM4W++ilX+zPELnKO7T6A3GSMDVnmlzp1ANwgSXgOFWXcQD3lg1gN4cVh07gGavPX
PEYbGp0wf9A3DOlsduYv1tJnATDHvesyU6/w2wgbYsVvuvICn5Vt5KpYj06Y3z8RPri7/1YBEfv1
gJOF+T0SgQMeL6GrSaMkVi+GC8Il2eZRqPyONQ9VD3XwVCS6voZ1qyQYtkx559Gj83QUhxiwSPRv
rceMIN93295/BxWrlbBqOQSmDsmEluqkL3bova6DaAZhQyGIGTGgqbOBlb3qSMbSV/hKJCz05KlQ
R32dJeUh06kCuWqiRKF5lckuRyiIn3hwS69w4F/SMP5ljt9xMNdr17NeKQVWGb+MARytV3a2AK11
t2TmoCDZASjDkCB646fvoPsZMSGxllEzefAt9KdG5izoBEkzSkdro4Tbkyt+NRaSowhPWseUIMFW
p8EW86kaywlgFT5qYRRFfcyodbdRJqxsU9Znz1Crke5p2z/AYrdC/x9EFaS4+3IySiXfoEgV//QN
QB2B47/n9aP0jUlnjIlLwzCRzXjzbKMvJ9FWeBf/ECKFu2FboFS1W0ZrikS/aI5zqvpsRXwzfKE5
cpLuyQqaYNt3BcoG3HeJGIRpEXEaNIKruM+8oo8G5pDSCNakEOxdES+Z8dm+Bav5yraNMTtpX+pP
UZ3BF9NcwLXaoBpT1NKizbYMPT1gZ/zpgruragvRuzaZ5UAnihAeS9n/qk01rjZgDja/fCbpxdNW
I6qgQpxDUKHUx2LTRrw3MjaJkjvLE3vlPAQ4BsoHyFIfoqAU3j7/B2y28aoWCN4vQE41QC5OTsc8
C9CI+wmcvQP4cN+ei38m3Ij8swBJcdfdlI1rGdX41nH5Uy0OGMHvZyqrBVLNGln0jPwq2pmoLxUm
ZD+oYNNs2ywtsXjEA42f6dT3vvtKJouuM5s+QC8pZmzNnwqytcWGvScEVYa5bKiQCnl4CFhM73MI
SLeIGwpCQjtZ1ZQbNFuWE8kRqkiPHvRYDb4BE/S8c15tJlt6aqHMXb+9GplI9j8DZJlFuXd0VSEO
/27WDm3f9DNtHDP/QAjYXOVES87ck9RDG5+WweXq6BHMqnSmMB9j3EuvPAUBhqiTmOmJiPPvI8TG
lYp2hsS0bYXEaMbhJDnWqUQ/1AG8CsRGqLL38cgsDzJcUhjv5Sx9v4l1fPgzdwl8wNXn1q/HC3rD
Yx8++VeyY2D3ccC+qv/K7hZXEoYRhv7Q+AeaBCTwvM/hfs4Ab6oUzNKRkqUppI8yWkgDr6TGS33g
xXQLLyVFIUGuyoZ8vxaLD8nPMk86lMX6RzFTKuaG5PjbB2DOqud+fqpoxXd95+BvuyS33oyFrP2K
0w2NTgzVMmYkci/lxSrP7MnDHAaKszkTRDZU0KdJ06krvGRtfuJez25LVOUctdLjtXzV/vjhfFnK
+hN0B16KrAWRn/M91cDHRcfwx88IPtlUCEO+VJ4eQCk9z55q9GAUuoFZ2hGKvXRpYtmYQ1/Oxsc/
exoZMe4pArLxtQP498haDSFheNkKoiHaBAS6xYoIJoa5bXmpcoC/ktoC/cWdZTC5dFDShAYStjzA
3r1FDxYwUQUUtyLpC3RGCj5ljGTBIwsZARS+GVQHNXfqZRrDtRBCdggENg/S7Hz3Qy0ZJJgYMYKL
rkGMVkTc3zYZvhCXdN/SDPZQRIFXMibqHCS1BCcwS9k2r2fTawIRYfEt7QyqUfMUSmJ1TWURGq03
fSrOQ6e9uuti6uFnRhOmyna8lign8wlaR97TU4WvdS1m8edRDuOX8cQOdi4GLooHiR7d3IXI9J0D
zyZHbW6ZRpzp5ao122QbxTDRZxF4kIH3pUCcBYmmsxkCHzK0Hp1NbyS1DMIh4CZ//bAPo1Qk5Gs4
UqWIwJeyk0aUsGc8GdASkocoYtmTVUIm3z/mmG1Nx4xRNp/jR2eYJ0JLuVW3MgfoblEFXs9tkk99
YK9/3t2w5yJnr4Q/yEClELfG1kApeuZSB5IQBnRLwQM1dXCh5ro+d4J1VmFv29sC2X91PuBJ4mYk
3Nqf5Tboi0lFjP88m4Qecp7oP8NIrQyXUugDjkdIqk0EmeQbQX2beb1TV/Gu+VaCypmOZzw7iZyC
ScExywnCeVJl5FN5FD6MbTSl/WhU+KnvoB0Opovp7IDVRffTV+npTNpsZ/mABqqma/U9DDfAH71k
U5NCn/JzkRKgUzQEPQmv7OjEhwCQKHjMie++mbpFKynPKIWOsgosEbPQO1i5Z4PDEHUkw56xwTSt
IoBjvPvUnfKuc2BQsNfiEvYmFXZ8BZEx5H7eK8kwih2KTZrg6xUFf8uzmHbN2xkBl2S+byHIAN25
aMQZL2czSjzzhRYAu8gcJvlPp9WoeDTCd3/V+GNg3ru+n9zEF/iibHnrENccVnwRwFtxhjqFcN68
jbPTBYE7hknWtaFI3fx5mj6/vm/DxL5RjGbGweazfhABvCxkMtZoFb/qVlsP0SteKs7Be6XyJu3N
lZ8y+I6TWdARglDqOMh8tcPibw3KGlV8Xhi8CUGPrzrHBWy2iwsspdX3fgYKwxFu0TkvSlocQe/j
l1Ymc3ODA2jl8dFYCN8xSOjUX2gfygbAiPxFFJ63IwGhUaiWiqahG125DyIv0rryU0wJyYy7eS8Q
HVplJCeGo1jMSi4XAbMFyg+4vZvKYpohS0YqSsVPFRCG75tYjFZKIm4w4J44725oHwdpRBL4ZJ2n
ApUZpp5bY1bLb+8bPer289F1Agmf9Rh5ZSHsx+Lvvsm9Apg5q6ijK1g6XDPt39Qkz0SA5NHkFeF0
s6O8HxmbYhmEptxcluZb4GqALY0sIxXQUmqhgEz2hKTXQHVS5QbXDYOyl9LOnWPZnDxs4w46aMCN
/EUdsakQD1tEa2GUfu1aMoI09NF/AgX/tC5DwByWedbi/U5SK9R+1HEGBJVsC6A0pNSntTtZjBwR
10SX9QLtt/o0yor9cgVSSpH3edUAepDY0yHlGIiHEPT2VkUvLaU08Xa2px7dqgwJFyDCt0cozN2v
HZQQoaeSLP5BIJ8HxaDERGy6Si4ok9VJJzkGiDtykEgQ6ycpa6T/FhA1AadNrIezziliKTTNA109
4ofj7p02wLbIRCF5mvMWDIi2EZKcViBjQreonazJbP6Pqm6h20sUaRUjz4WTpgM9SLE6YuW6g+az
fH+xAFehadrgWRiLCvl559nKX6U5DI0HNzs+OQn7es0PtHAIqoF4PhhtW556K6M4HXmhcbVGRbWo
gPvXZ4PuVYNiLFc51m2bEtcNn7mejx0XEPSwuQcCN3cC+z2Y8XciPSEZEdXPh8otD4XO3OG5GKLG
kzW2VGGu64RKEnuCDbNxaxVbgngAm6249B0JCbxMnI22rYvL94VKe9fxKU7n9YES7fECvKWfM9Xo
x4L4WZRkP08HWrCGBxTsmZdM11FrFweiYuB4YOHwZFWqIBokjiA5O1iW1z5QtGFKqxvyoEsFi2v2
fN0WyrXHSxM8EYI0cKfjT1/7jt8cA2qUXUFupTmT+MBwuNXWpy1VT8OGw97y+1UIlg3ns0xLBKHV
jyuERIvINPTxDCGqK9eeWfBKBiCSx46B9pS+e/WD7YeU5ORSfEay2B7/6HtyOYHPu/2gzqsiGj9B
hgi4hJ3NzHLU9Wdn0Unb2Kf2aEeLcMYoxrldfyLTii8ItInSZQ0uAKuFD4If3Hb4QgVZSE/TiDET
l/1RbvJgjcNLvsUoGYwDdhtg8dcnXrgPaZ7ePAyhkwEAzmZqF2QjidYvgNzF5WNesVjUSPWPuVXW
XRR2ENH7zSoJmwReVF6W+qfkUvM5W66iAcbfWFu/hSUYIdfjkzcvjegLmjs/4TStgpCFoK60iXxR
hitCwGXnDnhPwczzOwAkhgSr90DQtANzkIaScMVJYkHRd440diZ9HzrFD70ib7XsJfcyOjyrjK3k
/D7lgIdwuIPiNVKMwIsE5rMty8mPgoFNcncwAx9p3UngGU5veWw9KsrlViTL8DvyEWbOD20w6pCM
+YwGLXx3gsqo/4bUkn+3BP8TTWIL464k0fKGa3kLQA31Z47vksq1P5b0b9zCQeGBsBGabNSo75xc
Pi63Gg6+pfZ1C4AfWSXD3qpdU1ii+hXJVA1LsQocGIcfJRTCS5ecFAEekSgUEFtE2vm8kss0C4TH
3D9OT5MLPAaLSydhKO3xf7HSzf/r/0dxkjxXB3qgXQZG4NTcysWNJVieUDxHHuvs5UJnM26M97b3
OqgwfTHKjZ07YMhNETlmWzdxczq/LbaIGYHNTHA+yU0HhgXdZ2ocrsYEheEjlDwLEk7WRf8xYyAt
acVCoD2KP8IBmIYdjG5eLogFb+UctpsSXeE8uExJoEAndvBOMe4FcMHijzSyzFyBp/uV4w3mnla/
/kFKS+gBrGVfoanGSdEVrLr094xMvLQE8eaEkE0OLkfICf0oEQV16F6LPlGf2X/A4Ak4EhltRgAS
qZbMir7XBIbSpM3k7kRP0dCaUIAHOPbB4P/Vq2Cr/U/ERhOPkuS6BsJbClHUYa+CwfnAl74JGoTb
FLDxeII5GWjm4sM4N4N8FqPo6WZE8FjgH4UUZYm0r0oekGpwqZwvP29IDmvAIqHfm3YOTl5qvRHf
Kixz4eB/8NZkdXWzKf7Gfre1i6+OwrAn31dBoittGP6z0YU73OtgMB8Ilp3uQfiRIPsaDDX7r5CM
z3NhuNV0zVi1VPI3YIJ3elB2aBkj+MpwGCs8AVCXJpjmzV3XmZPF1znkc6iGjNoMOlvn6HZcfXsc
Ro+Splyej1tL7KadgysAzblVslInDkyf4juBvbcx7b4NhElgT2XyTLu04EK9NxtWb1fzB3tvk0HI
naQuO5AwiqNelqLslv7Th6YVnH/IYTgGFEn4LVIijHONdGUZWYQrraYzg/SoRJ6N94lQWYNDPDOk
KX0ecUVjhJ76069fDqe0FBKVswyBe/QhhretQzcRxfThX54pdB+ftHmXLmP55eAlScVY65thrBrl
9vs/7l6rqYznOZ6nS1AulgLicIU8tmbm/GDu+VS09ydLVOkda8E25IRZhitfxcN8Q4e9GXi0Zh2E
sbJ9Q5igpgGCVi5vclTt7g1TbdY+vgwPE4tNlDEj+waEQXU13nFfVjk7FHovzg/2lgXR8JJx8GZa
OxymQIDfhB0mfZQ/l8DdU16z0k/1oZiDDvZaNURDjOK8ieGTphUcxA3apZXOUOUrpWIj3NGiL9R7
lo4TN4HSHvG5zCynXLTkKg8MPQCoV7KyOnEaCbov9Tle9VjPw+xTfB4IKPnQOtpOE5FFZwuboROq
gm1NcxRXpV1HafvSX7p6lkF/Akg4Ap3X4AlpQnq+GozLg8e5fkcgzZvMCsShsPAIh856WSw1e2N6
RoXPea4XX0Q8owdQFjcG8nJ6cWSZ6Sqmd5u3P9PilYqC2pmMy8dq/bRs1lbCeKzZTv3GoOrq/nna
t37oF1Q4G443vJw3rgI4/qGX9jJLZygfF18Sb9zS5W29WyNQ0Dimqpn3svf+V4vJqiTfn7MrJnzy
Lo73t6zjK7BYKENcbCBmjAi86PTPuTT8PThoEVztSYP0OHgXpTZgVDMtFnIMdwbTfx+F3CTlsaIn
bJgLyG1DloUBFNAfrmJaUtcP6WJo/x6KY8KSUf87LVaI8Wb4wFVSRuVafz8dxx84aroa5eaCAeKE
MwZONiteC2oOq2RIeBuQMwiOLaNzuqskKn5+NuUU4+BOORudm/gymlkt49fNi/gmOGvuBilkLPBS
but04v5CTql0iVWonMCEjhf48dOqpL55II1g4niN3uw3vQfMmI/nwyzzBt439l4QIGRbwVkK/xGj
+fumZKp7DmVLNKDMBp6ap9/73VlhJuAnHifHyzQaq0GscuK81p3mfthpOrTjyhO+lL3j5wfInisD
4O2ieZA1iALw4yF6PJFu+g3sz3VoBD44CePB3xzPz1haiqXLWz52YSEQG3LaegYTwQA/wHVJZT/X
a/bLPltcpIDOM2URemd6ZGuKiugzQSfbni4Qf/wGpgwKTs5VmsUi/3y5IpTv6+n/FJ862MHIDGCh
nMMwup7+rXs50+lD/OUyNJwfZW+f7TUMjAdOd9fo0b7R5AlOPFTWItsbUhvGKOvRM5hhiV/Q0k3O
JEKa5YPIJNWdPX5rnFVd3l/GXuVxMKZ/8t+Ood5PGA8J0oatP+xef0AJrh5hhAk3/JpC8L5M1BD4
SU7p0kiiMzb3iOgiB1b9jyCz+KqJgQDDMZIFevxd9yYDCHeGX+dcRVYV7tvlNZIoEBnEAT21Iixc
nqQ/vN3DXZEod8Pdbi3U53nrvhIx08Wu0YT501ggIRFtFR4ppbinFgsc7/ufMTX99RmprSe3EuBZ
kOuAfTnCEAyKXv+K5BCVReONlEUEGtDsX/honX1NmgV2CsVwdXaG0cOj+C9EsceGsKweogq2slh4
buLw9jJHNBI0xFebiIruQKtSuJrPApFr1W3uzxzBqjwBeIU5BAGl2xCuMlVU5k7rszm8eIIYdo+5
oY9aCCtoLfhJVnm6s99jh+f6gPkghUP/oKVaA2mW2MF9CRC0DW0dl77gKRBAv4bzFvlSDUwfjVcp
YCwQ+JGEwqZ5eXxsDcKzdcxbR3s6MLLDbFChP9ie2EJY1/qOD4Ie6TGhapVE+I6OVxG7Qyl5k4k6
rHvBZ5rSISIRnX8eQGPwNhOQ62GHjARZCxnPUEZobJ8Z7S1pOtlv9g6kOkY+pthH3pPXvJQiKt+g
NwIEqyfi4oMOmux2/SK0kG78sCIlPDkv1BSKI4WdX4HHY5jDZgPrDed8sfREsGS9zYWWwSY0hrGu
15I2LV6a01QkQO2DLSxewpFvO+dw3CJcyfawq2TDZSicxOTff2qOjLpKMkKSmppDmpY/6ijSSVi6
11OSh3FD/iy7V1QBkJNcbJr5v0o4oeuNxRjrhpzHTh+zTdh3wAc7cbN01ESqX2+mfDBqGuzagUgH
j2NPiSepIBQDxAUI+JGPolWLEiHHvAM+3nZnkBPuqAbrg9hIZv3nMMfuGnKO5zvkAeJD/m8Cv3Id
DUnVITau+iMD5WlWOVwZ/YrkKxKUQFroT2pKVBaJl8berAMLi1+zFMZVI3MO5mI/lizHMZ94NKQN
WWhNFwaD8g3KwJsACeIP9Bcet3MN/Pzwl0GlZitDkR5uQJoDUfWtNhrCTHYkNlcrI491CJMF6Pox
iqm83zrTtH6JaMBffaSTCuf+PmRHUbxlMlzqeXyIA/UlTOyWh8xdLAUpPhdzrA2MtJbftCTKBD1E
LS+ADa+vtrpsCmPWbdhqgvhCrWL6sj8+4VX0OsJn3VKGJ95soakCFXrsFUzMBOYhI5vldunzA9ue
fZPOp0U5oSBwKDySr0C5jCPtWoxlqfcvpigNVBgGwCmQgK2uI86/dGGiebMnQR+zmS3q7nb78oXF
2Y48S61E4qEdNHsCHWL8HMLYBUrz9RszkbOSLxKVL+EegzzputW5O6KfmNIAJaX1NAqQkl2OaI9C
pYUShqSiiLfoMZmGHa07U0DzICK4pQqWl0TMGhX/OFzGyVUyFDHl4qQ44H6dlUOc5s10ILZwSCA/
dqeKZG1sfPsRb4mPoOH3e4YNHyzCQL648bDCqNMHQQTs4RAEHCNs2aEM1XozJpZ67Pl6L78SyGRS
U0EQsQZ1qAbcnWtBQriUnPx19x3o2qs0nIOnJKtJjbDpGYXWTwvURZqOl1AoQlkjd0Va74mAMBpW
KmuE6HKLvUDfbhLCdq/OuWcrIJcjGM1xITpqMx+ioZEbzXInICRRgDHFj1McOf7CNOSZKo7UdM6V
t2f6QD569W/Taq32C4rvwmJIqiynTnRoNDzCkoemToJapctOCzE0Q1HpIrVtujzlTloibCEt3blq
if6P85AJ+LAkq/Gm0/P685OqLiyYotMrMelvdLO2kQRfIlwjJkbJmjKHVgWNVXtUMlJ2iFUE1mWN
/GdDTd/pdfFhhCALkCqkX9zWgyXNntWd/rnRnzTlicwBbZuKkiPDYfBHvAX3VVesWKF3epzEtLZS
quURPYRfHC21G9cJMKmHLoXc2L7QNT0h8pn4dYPodnvTEykMVb2EtK8Rufst6yMLI/9zGMcbBIm4
N3wYZaISdOckMYescaTNMImtatDoP0Vyhf8CeuBnrHORONxCA5LNOHgA54Fr8pUouwTc7uT55eYO
KEi/YTIOboM0qNK+OTUSX61UCaJpkbf4tNsGNJn0lyNapSZnEQW0T886vdgSq3uUhLNTqaMmFofn
RKeONIT/wfqvEp1uOJAMheS+O47eBuHt2AgbiWhNemVmlO1nnAlMQ1Jlao6hmfds1AcUkEaEtfTm
oLAyubNPah37kPUZyS0a9uN9pBwWPbw5lGWU0TR5hyek9jDe6UfT9v/0v3Tg3SVeKvEn0P3oIPu3
USqmrhmJfhbbdJ7eU02qq1pDNgTJdcc1Jj2m5jLp7GqfDADJB99Yw+9E08wBvthvphITAA/ihNzy
Odt64MLDNmJEA0/MID+5xTL7iiKFWaK+O9tD+syIu/jbL/bZ/7gb1nVSeH4LA35L2KDdaJd1/E7W
/zfaO0FiBvwOX5snuw2ywndMZKUIyBfn4tT9uvI10AU73wL1KH+4TFWnPDqNHFofvjIBIWW18er9
ozMTDFJeffR3h7ora70vMGSFF5x0xAL/cY0crQNjn7f1sGOsoSMxZDqaUVeKpUnEp+rrbsF7Vn3c
l5CVsYFyv7RAIz+5/oF5CSOIGvKPTbas0sSn4CKIuMQmnUHiTMNCd7lwqVoJXZ7hYE38/LExjtz/
d/PD762zhqvY6kt3/lM9pQCQdwWGvBmiooeqmALB5BQLiZgPPKjMUGDriqiYzKujs0Nc0xIpQIFQ
Kdn6FhFTx9pYi0Pm9ikSzzecumL8vgTptIUrNX8uYmSRz7tscQ+Xw0FWewm9GsjXTQq9KtWHsCeX
RWZ+E0Om3N0qZPtD+PHCYa9hNEYYMl3P/AzM3eG8boEDgX/7vBl2W2qsKKLagfOcIfinxLW9XpB/
gjTsMeskmmTHbaBt/iFRx4NqNWMF6lmnWjOXhXimliFMmO/Nf6If2pUXlcvOsr/kal2kLBcNmSbL
Dz6LH7XKGSy2wUmAl4JCxPUENdkTVWQfJsccTGGNv3FzLcJF20PjRYKn+zlNvl/0WKxKed9Ssz4p
KTAIOM5DUpxmriixg5jsb6iqkMYF4vOZxGs2jo9Jsz2wfJ0kzKWT87pTGx/GyMnIZ3dJ29NXZ1WU
qCf2abeeaAjl7Vyaf2Orr9GSXTfwUz9/A2JvGFPpjgCA+LF6nhM+9RbkgG+7Rl7PKfD+HmaPnLbD
TgmlskBeAdFp/D9q2WDrtfosbE5iPE0hGeRYSwRXA6YF+vl+eu/tQaw6LYoU8MUcsUXkTHGBjCdQ
RM8CNI1J7Ocd5dO2A/NmmGSO7tMTTdujoveYsFuH5Jsoe7JyW/TPeFsQPxQuDBE1F1T9RBxJHfW6
T5ljoh6Xhrd3pi0FnmAdcKtK+ShuR5ZGn4yC7JmXNsbQMoVB/Pk3I9vYFEdEU9yWxf5gKm+f77xi
2Pm+8lR/Tx6quE7W3qPHvcZTpHhk+D7D+8CLhaHQEaDpFrmxkGXmIHRnGzBTTjOEUschlRkfKx1Y
+QajIip0j41te1BNhJcDHPrNrbicAYfnB7Atrl1ffdNM6iafoKqG/hmUPf7NnOAJ42kmbpaZ4vno
USwHkRlWCmavhhCUHxzOmghYHU2mNXvZbVvZFsYeo0lpKY0uZgJUQiwAn4AP8SWSJoaY8PIUJ2bg
lZF1ZeCdJUpK7ZWMMNpIze5/YLIKvxxFWxXK813bmVTFDy38S2h5NnB1bfQwsDBQ+bnKWD0wzp3i
pydKJ5YAKeLALC17DGEIBUC+dtAajD73puLvURiKVAwnFBTwFICGhEShwQ9tEqzcaTOww37gE6Ft
m/TjQJUh5cdKzlgNabiP4dx1JDZ5CgVQyQKNM6AcFpwJEOtN90vJFGIP6sMS/RnGOB/O98SHdfjg
ndzpCRIJIdafFF/2vjgbFUARy+v5JYUPbDGLalycpIWGYmVmOWsMw71rp9yL9paLxEHENdMAa6UD
1NweVNn88Q+kJubJcCrYYcCOiOG5UEOXW/a2uMZi43VF1GpCiX/j2eMkFmvwbGVsWONzmjzEnBdh
4yMZ9SljJ2gtOxqDVXyZX5j7CXBSofXrEboMnS17srScA1E/w143VMaeQKLB678uW1Z++HPFrqZu
u1heL/SfqQYUcqgdRbW6yB2klyn2NUjCWD1iiGZnt+74TPi5miBrzBEtcugwOYDIEO9PUeeTgDlF
IgsZbk6wKYqQVmhoU6CiyPHVJa1epYkvBbVRRPHSOoK6PWth84ALjOK0n7vfSW9ca/rEXZ8I7YW/
mFHKTb4kvaGt9PXFdJsZuF9FgxoMmA2AZiT7AxG/U6HOcLSq4zIDtjXfOKco5B9zv4wIC3dVeY4g
wzrU37bImpVS/V/wJlJVJ5rgI4K/yX8hgI5DLj9tjqMWuxml1i8gW3IzsxsCl4NBhnWtUVlP62qu
twwVw/ypy/0M03flT1HM6dWAXrPyC4i5P5tARhQML6pTZv1VPG4cvXOaZsEs8QILfcfb1djqZypd
VKzh6w9fVWtlkrCpG6zIIgfl4dqwV91QFlbJtj9Zxqpgb8KXIOpxMElTjrfUBgDpHj7wU4MI89TU
mjHMhPVaGxYUH/92IBNIrVtvsWEJJKiJI+Almr6i8YMMmiXNsZUjTg4HU4C5OxfqYMtYlCF4ngi5
RQmF9Jo08yWW8ncxbslL83JhDMojvV6Pt7gMU+kU3rxnMDo1rRL4SEMUJKaghLZlD2/yFlMIkVnL
dV38AX+jeIbluzbiLz2Rp44a5+ZfXinoF3n8c1u2aGtJwu7bMhPzft2NuTkT5KoymbBWaKHcS3zW
n0qIQWf1u2F37QETgpnyasJQVQ1d31plACFS55FaBIdkcq7QLiYNn4BZ967U1KID4thmruiPi/nQ
5i+9Buy/eFAg9L9e/YGHekkkVWY/rNDEAwNlklLYnMVfQzTQ1CSGKA/itSn2x2h4qND7niSikgBI
dwpLx6358l1A4KWLBjmOXy7Q0AHALCafVPrQxVfK7UYYsMR0LJI3N3mLC3Ite+VDTeN9pYBwHOHk
GS/PgbXgUucll5ctaWV5GDMp8dqK3xFPGVviuSbT7NtU6LQLRVHaeIZsTSwDM3icN0qQGtLi9l64
YaT6vWxkMA9pzyQgLGvycwgHAl0AQEjnp6T/8d5ILR2cGTK9sJr99wQzMXYTqyWs2SNE2xEJIpnD
DbXCFAC0kFqbZTfGPWQ+DOEfFFq37Brw4PeC7ttm5QVZZ45rXqlQFgS6PgX4zOIBPBAcy+tRNxyi
mWlG6VioQecjrTyZJreowIKkXop/0IXd7XUctCjDZkcxSoMijT1uwx8f/WRHmVVQk4ZZGEq+5s6O
5AMwdkAJ8qbc8bneqPRtnzhLlQKUo5vNCmIZSLt02d8SEvu5ZyY1SE8Si7ibpF15fe0oTmInIbz0
iBbinAzQpf6uZr4iNouAO6SXPx7Kfzu+REL86I7gTpR3u0Bva9UUIwu3Mn2fLnW6PJfLwO5720Ih
AEZcdu9k0BLUU9iKLifGlst/ZoTrPQ5uuMPQgdwudQg/5MrJ8D+RiIMJVOS1Ex6g5sQJuYqjv+nK
fbGJ6nS/fx+NotsTo8Hc9zOGNHrMcFdDh0oYrWnRFYOTm27HLvMygsjtliCKqjUGDsyHqiaHhwN3
qNfaTGxs49OCBtknoYUXXXx5ERbblFwh2lR9GaKhupRssoGeyXxXPDu5Tg0LQJ3YAiucoyGCJxts
aiSLtpjIcrP1p1Px0kPuT0i4xgap4IMMAoG2xnwYQMLqASGSpycU9Y+6H65BN/WN3VrmBE+iYwmi
IibBMifZARwSnoqNLfUP1GnrKWRXmQNCDVZP/W5IIOtrKJzB8iwhDXTn3xI56LNr/jq0mJltcZGP
UGS7+BH6tjwkur/BQcqcbqrF/I80UU6BsIAMtB8HI9wKu1KmnNiV3vCJDP7zsW3arIeNpBfC6xJ+
+DBz6/YfMVEyjG5nqPnt/i5YZvPYHny9P5u+4PEg1GZy9yR8t0KPqJnv0la1x2buNDNljPo9ZGWR
IpfwWQOWMs5mFlNpDgaVoqqWW8Ltl1fATPPe4icVIfxghHziynRoOtGns7AkviPvHPw4WwFcpqpc
5rJY6VVmI4CV67+4JYrrzawzmGZT45wB1wQGxUmvJwmaY6NVcou+VAmNbla+Hnq4vlorgQGEHApT
AtYhk4uoBkvVrC406TbgKy/J9V53mrZoF9ZcE6vluS+XnafeG/9LXFPHnTgO2eNOOVL8JlkNsDIv
Vna42RPtIr8BiUwDvJMkJ6n2uFOxuDBHWq0JKlCOYau9ur6rYkpfzMs0ARSieya76sHK/gh0iO1w
/hUnwvDqF4rUPbVielTa4fkLOpiaX9gNmzkpe2fVRmvoQNMvOXGTCry5TcdNMDIKzTI3k4UEhNtJ
UDyA8Xoxb2v6ZljWy5lZcYqwhugGHt6cL1Uihgv6HTdLAgnvQ/uTJAWE0it8DGjVt+FzdsgaQiTl
EsmxPNa5TvMIucCmJSBGaUaRp7zLtaSlnjA29+fzddwQ5AsnxxfnlBnKS5BBUyKWE4MDkoi0Bh54
b8D5QXhkdaqj/cOKn00l9lXW4g7YKpX3t9ThS6U+nK6UK1G2axW8u7/CVzX6I5J/CsTxkXorbKdb
Ain2+2k6w+F+YBd3AIELsqNnwTg/33rptjIuerfP0bZZJB9jnB5XI6+Nw4Y98KsALiaEbcM0EVZw
Y7wB9To4ZOmHcl6p4STU8PtjacjgsBP43SiGNEDV2xn7Ujo9NtHLh/0zOhIHoq09Ma231Slnbqhu
kmG76Bud0K2r8KQZ3/84WT0KmsxtZHLpvPR+WiWn5wdkBE6JM1w6Dcy1PbuOC3xTT0gsrfiH3kr5
ckNBHFQX3XbsrjTHMZF/dUih0OQjorDlyxEg9ck9R7wTFDL9qVdMN4xZ95gaAybUmUWxJ5YVCsc3
qpDXQB18yGifMxJfxnB6WljRf0Nkui/Fwp/5W1AkqVNnNYHFDsjIm3mFM4pt8TqdYe3qu6WFbXok
NHaNoyS4Ms+p9w16CdakhXECt27Wdm1ayzdFOwAIUvH+0KT5sljqCSEb5Rhm3UK7H43i6sWN+Frl
Si7ljRlyT+F20/sUKu+PtYLipw7ji6+2ub1wVOtNFaWnIe0+BHlPwbERVjWVpF4QHvg4xS3NmYUG
2ul/PVO4KqDRGrBjC+CEq9ojQLiqfsxcQEHCY47qLtPXRt5/bE7zBqo92ajv/ee+T5wl3p6IanaO
xHzXaHbWta/lSJ70ASLwv0OBa5wjDbHzz0UInmg5abbV4luQAF2g4tN3PfF451YSr+DfV7JF3Tla
gFXf6Uu7WmZ0f/qV4X5cBLgg/q9TeG/6XXtcZIWg9y9BLmEegVKZDNPDZN7TlyaWAnU0JVD2UXTO
qII3+sRdaPG66gIdFmaHmVuaJO0Ixh/uZkkt0PGzpzREoQWN3UEJLsKtS72C/gmxKbGWSmMrr1m1
+4eyCKgUTAa4Ejxkf0v3Kh0+FhvAbNy1/n3hOc69D9HbU28XvnQkWnBRRumYakThu+dO+6DDhXwg
YQvUch9d3uPOMttTlBI8Y190NKfPo51IuiunEcMCVZkQiETxws+9MRLUlA4c6TWoXiDluDNxe1Yy
fod7tY1+mDRzS7D+3yAcdqDF2KY/jT/OiIP2IaKIRyn8FP3H7UVKNp+Jln8kOlep6StXJ0G6uUQX
1lNtVIRMWzE1LljPlNjiOpvjuHNRdGVEHDgIvIG0m9uvLYXCSTE1KD2ovXSw9cLGK2OWlfNqEsI3
YSTXnKHlFMrjBbVTphsOqHnzPCgEx9TOaW36IQbWsWHGJ4Gsr4sK/uIfBk3ZBZxaGzb/MSzl/U5b
1w7DdcmHyUNWNZmDw5f3yYhSlLku8mH90uNm9D3aI7mIIPEr7V8CV2q5rFu0Uogap33n1rUQVFEy
MXOfcM7jnJvj1qcGxJuFkyYuLM31uwVEoYuGSz1sosiRFWBd/GiAu7iwJYv5xjgp1UGdM1evUyNO
ljYCjPcqYpm93z5KuP+EngHphnELidVuh4DA+DsFeda492wrbTSCTP/qG8WBuyI9bVZFBBgBT3w2
L6X9S1CtJZc4DxZe9jrL0ucKh3sAM1YjYsBD36Ij6UaKL2oZYyPatMNyx4SJ2Iz+/D5j+Umqa/dt
Uod3iw8o4kc4AuVEnGip5rkkAVhMWESXMLIEIWB2Q1of4wJ17bd8dPpqv9En4UFiyxRrF0puTU0K
mJJTOwSdDbTtIO5hMLLXumfYnT20zkca0yi4CgsP+mSZQ/NaveSSmBeYMoLpvkxyTJEwSWr/EHHp
vjO6ouujr1muQ2x0Jn540SejVJk5RySD514zYwyPlKL0AeQOpaFQXFup+Gc1lLErJMRLCYM5CcaB
f/uy48EPPoxg/NYrtmaPOl6Sh/Cqv2oAN9Wh2Oi009TOwEJ6ni6b4ImVi73FhzdrFN00AZ5GELbe
uxd9uc2p3p1diSsXlP24PnDTOrewjkC6sKjRchNCq10dPgac3DXkX5eBQ7Cwh7FQJnTdDa3Z4ysZ
rg3QOORgD8XmPP6k9uE/Lj/D9SdvCBQ+lLiG/nclQt+pZ5DstYQwLgWo/dS4nhjUf8lkZxAJnd9L
qiTO4iGvN/933kBrqqZc8NnD4xIfn1JB+tPBZKEzuBFFSTICbS+OKzFALktXFCUKgqTYLzo/rhIl
fPIeWx3Ao+fZU8ouf44udX4ASJ/dC9yS4HZ5arB2qv2YfeKvCovpulyyRjJF1JeWVk6grfOapRi8
z6WVslxiortmhLbiRUholzouEl166uSVoeYolcch/DGSQv0UPTE2Yd1fXB5klZTXJMjLBy1/wPS1
JNvnDZhhN48kbI5hM3Jm1RYxqFWEJTpXukyHT4MZQej6ht+LtuQfmAw9Se2D6DZsAsfeErUI/Yuh
uNO0e5eO/c2FHFYHJc7OOpVOVS2QXX6PTrYeGB7xk1y6r0xXKniYxazas4K90RFP4pbiEVsBkYuv
b7S6hQBJkDpJEYd6Dr9/PqoJfbNuqMAySUlKYP7Vm2tzIRyo3QTNbDRCwE17RmmU9FilZd7Lgexl
XJ4Gqbo8uVKAEUQYcgVJJTIxD9YxUPcbVzGrQAfHrUGcTNv3KUAQaYGk9MTHabsFsnFJwlbEIvW7
SYFwDpSTA+VbF3wbJCHPl5PGAeY7BJ/L4p8NjJWPVHZn7QAhb/PdFU2EsFgOfv3OSb9w2G6GXOVl
2Kejdjc+ycgMGjJXggi5zsma//8/sYNKbDadb9JGnLrp2AaE5YfScMUBM/wJyN2pSjKlSx8VgTzh
llD9hGX2eLnIiyoXIwXCSJ6qaMbm7r4G5hd4JwknU9v6w57z8SSHhgOX3JkQo6oGCmJaDw/Pt3FZ
YvJUWI+7pTYV5D2uPvc/4CY7i7VDkbgrFDu2xT9Zi/WORX+XZ8C67VvqoUpdOsDKRfH/b9S+UN8r
6avYyeUxt1rN78cqDb/GfYtsvP3ZNErdo1HjqzzFTgl6jqeTwB83YuWJnSnvotdhG1PJQgFnlN9P
Z4DrL9mthAdKEs7e3Q0uewSgFrG8JuOUjDXqw+V81AEvRJnyFILWtjwbuwrbQAzFzmP1xZhy8bRz
ayjM+nVf5YT5wO7Jn2ekOeqzx7MlZ5MbKkdPAZ6UIdqp1xwrmz2HSlFcr2xWW0sZKnA9EEDSpR+A
4BYpQnf79MEkmpXfDUf/Yk+PjMtecC+ckFDJlrGG0+XL0YiKeHySRyWCsXgQ2ue1wKWDxcLKYQ3C
lxpKBofQpSSP5fDLvTyXMk4wejI0DOiwHSV+e2vQYpg+JGh7ge3D/rCtfkV4zgvtB3pJeGXJ8DtK
aUywIaXQqR8NEVHTJbfAgtxGAAwQnb2PeK9zxyGU5SHBtWcksPBOBD+r6WCiL1aAh7F0ZbvFNRce
0+I4D5C8KxXruHFNADauT2SXpFVHFiQFcadzk4tXGjIlixtBcgCEJTVCk/u+AuxQ0/9HJtDYKEDE
Jsdf1ymktA0dEhPRU9NUmZi45aqoUynpKf0QPysYz7v6BRm85pffMjiyz50yUNMCiabC8KlXJ3if
c6OCWattUvm2LIduR33Rz2+WZqipjXk6zjg2ZJ3AzUBtIk/f+Hc4KE+MWn1MdqWOvVURnLkwrgm+
PEFesw+ikxN0rFC6cIp/1IZYvs2m5/s+5fQAT375+0FcvCalp1Xp4Ja1PTj2xqeU/s0UHouSCYGM
5LlyCMIRO7qi+YN7oKR6gDprXsPmjWJ0p0HclGHcbnZGoC9N81YCDL50MZzn/FrHXh+bRI5ZcEF7
8qTlFDtE0dp31rVBHuem8oiHpDAeQO1ztCiSlfmB/9YVVVFWAKQENwxOx78B+R6LRqAUzrD+xR/c
u1uIPi8xnTOCoZHzu41CD0Oqv+JPSK0ygrHYnXvTDi6W+37VT9L5akxIHl3Vlxl+MjMNi/OngGgh
ncjo0nNOmIsQ7iRhUDbZpSm9+oet+rYdKh7ICekwR11GEwvNRYalIvn63zFvgkZ03QaRm5OiBKhO
ozPkoKMrQfzY9JtISnQF76qkDe6g+OVOKWId/cgZla8KoMHdXBcLaP3JIa7hlyqeQsl+YtQpNuek
ahlbSarV/BnaiGHmNB6VuVKHjp7LLUCu/BCq7IpRTHPXSGG/XTDdaOK9QIbxBfEjqt5HrSKvyhK7
i0l6bUuuMWeY8ZeEa3+CZiGMAXgiEhCkPqynzQg1H9IT0S7qzaC+cCdJvS7P0nz5XOwlpQtPg20a
dGzes0BFVA+cx+RrlFABJ+BM230ZxFHVap4bkYmDgJ87k20pASLB2CzCjRdFyESoBpwUz9i9qjxH
AWV8HpJE+NcVQT0Ld2NaLTYfJu2vgxXRBEAFqiKE/TaXPM6NynPbL+429mJW7mQK8906z3ZZ8Z9u
to+WP8z2+SNYYfzibleHIIaoljyompd0jC577VGI3aGIR9BlYH6t0LSQBVwIELxb9Dt1AGftWm+y
p11lnAdOt701VZdkjIQio/jbksdz7H1KDNLxOHrQevwLqwfPEz3pEyMTxIxPvrpXyGzqTBSy7p7j
WBcaZUGk+o2jKFjMCoJT2h3fSXwWUI07iiwugNfDFbGgbk4/9Uz6HuBDT3CWbQnCA5OY0qn9drwB
p5ZDoA3cH3EbkY1ilGCcudnkbIqTF1MEjbThUZTnFYcSKN2+Z2LKxcRNB8kpTr6q334PVKe8yU/j
anXTgJIvGPP9TkqEn+9ZWH3UApOtZpTOP/T0TaidU7oK9wd6k5s48We1IwMC96Ep233yLlwv22Z0
Qoc25gtHd1U/rCRfuUytcNc9dCz9+dQYtDSm8/Z63rJY8xrt9UTVRLL8cBt8O6ON/a7iKLGNQRog
nXgXE+WG3vgor6OX/4eJp626Aa3WhDpdAqphZsVjWxBKyYcjoqRr1i9iHugZ9OtbmbMMf3I95PtY
d0eAo+EesIGFmzcVH3FYKwE6pMkLcw/XX8TMnjPbneCYGkqecyKkU/F6wULS0Gn2oWITJvxOgE1G
gr2RrpngqhJGGs68UjnPEkIE1hQxD8mggQMm8AWluJ0hJ4G6Ol9xzjf9LFkPThyevMUmv76ihECN
E/3k3Aa7OvE88mJnfSqYVhT903vITgr0lDln3LXEl5AS61rK/ISFWagUnxXNfVmSlYIUS87/5j7K
9u4NbWnkixq+uD5Hyrk5Ypw5AUUndVaiC2LhTB1qk76PLouB2yYoqeyl3a8M2B9vN79TUZzbJKFD
XBQq7/YM4Q+UypglyPPqhFUXrTL4OwUsdTCcriXkFk4hE2CI+nB8rOK7HxtXL+Vh/wZTuFaeyuS5
7W7zZI5FKzZWiBpVUHUQ7/tYuW8TWq6HM3kp+gatC5QElKGaHNL/H09gQHA11xZhGuayeOoxXfEq
1SijKn7Br4LuRXpMeBv+8w7lWgib7KxjLOgpZp1gIWWOARsSo4adHSsysFZH8q6GhQqlrloGnI+X
UVqIVCmM7uzgRMZcVC81pKhtnT7TlAJIOYflAUstOuBLMzIzuYtvxzRxr4gLR++LCoBRKnTEFHGq
1a/P/CNwHhruG86+BLWJP1bbvQQVlEQGyWgSfae31L7J5naGL6yHAhOLt1ON9uXfqr1i92IyK/mS
kp8Kzg6zAdog6l9xBcdOEboFD/QdwhSsOBqTlxFJ+88dEnMFSRET9ijd2iXccRQEYzj+ihG0gCnx
ZBq7F2jAByEfw1kIEUZcYFVpWOpH0Y1qXQSsbh8+uZVAfmIECO1/svdGf8P3IFqHpR8PULaO34ht
HqAjQGO/ohWf5ZwtDie2e6WI57diMVX+ZCpCHg4Zws9TiHwOfKfcT6mGL3eQ61hIOs7DHIVhaTK7
QX8/lbu6TyNzvQK5kFxawVLVCRlJ6zeBYuyKtTXM1BKf3LtlysRkQl4qLvZgIu0f6kkzBZ7o+zF8
G6Pm5xxWBCUhgferfxNV9iqLYP3grlt5bNFBg29Jp30EF2rrlosPvSkXiddQUcddR0ey3dhAyx3P
tvgSJb4Ylm66CsOIrPKEY5aQP5YB4cTfXaE0v7j1rX9IGfce2ayRQiafdb/cEnaoJ+CNOnVkSg68
F0JeKDp8p/yFUSbWTxHUEFf1dtnXY22MkhP6kzKq0qFvPht/Ir7FBG64qyBNtCkNCvw0Z0JoQufj
eDpB3kJKiiJlxSut2kBwTydY/9ivGQs8LNWDMHjTV75+3SgOc9/SJV0ek8KWXCKCzfTuDgLfiHXy
Drkn2Qxe8BfXuOeCFvLaaJmwXb71eIuefz7D8AD4iLzrgEmYmvenpu+OAcnJoKHCnYOGh5h0Oj53
9whh4JNf3KfveY+rzoqRh0e+ZEBDKPHNUVK5/c7Jb1Tmf4lB/6ettGKf2ZBhtRfQdOBd7fuhJtxk
ws6RZXrx53zJvGtJ6V7zZm671L7AuMqPreoK/I/uOoi/MOhh7yt2IM6twtkoD3eBEf15z9h8nz49
vW4IxMoBXkCpwUnZEPYjPQr7BZvJGunbnF7skGRhXv9TZevuekqtpoe2eiOYowaqtq7QXdWqTZzN
ACuSDTS9Je6rljpTSE+U/oKBkT6tMV56UWbIRuGsDH1QOQvoY1cRDxQg4rnrK6Z+08OZK73QiLoc
C3qXZwvDTXP1UAXXIN/mMKTlUYoAC5yAKiOOmNN5W57z4xRiB7fL1Aoac//Zy6C18/ZCpIk90g+j
Y4PLYMNW4iNC3hLyX7YIGwFIwgjuVdaKG7cgzBZCr0KPJJ1Z42VG2iE9vepN7tTDJJXEWP2CDZFL
Zh/015qjrwd8tAbiHztRjpHevYY/TPslJ2aFjHIXtuNuDe5INAKS5MqS4vZcO+EM8zx8bbUZruNm
ZrWb6OrpDdZblk/k3vYzDysCmJDFDBredY4ViffREIJVlP/8riBvMKM7Y6SOpG5b27Np9PFWolau
fyN6B3QqHmDyd/fIfi8+aGk75tJSNfLXMpZ8z0C/hVhoJ4U0QZlWDlj4JVkeOrtvXymxLE2rFQjk
8eyOAaG2wrme7cg83pxtFP+rSSyk4l7yH4Mwew1RMcbbopu3YNmdEprw0Rkks4FiJZdVT6bJGqT/
rx5eH/D6vAe3+LD4B7+U5YSUg93mQjBDIywxQ8HnqebRNfyQeaOzYTJvPbjWucw7DltR26WV1rLV
sAvashx5D7y5dyiSlS7RueppcqYHsT6OrHdNU157dPwNXLzupWamDLcnsDZc52tN15hHannrlg/S
aULV+GqDqFzG/4AAkFAAd2szDH5QF7sbp7+Qdi19DP9bL1ZN8C6Zvbx/mcenM2qpyFmGX6mD+4Aj
Om5yQsMi2aMnWrFQjJU/0PUiKhW1oaZu63qQUpiMT/soxdO+4SwmcgMsyNVuNknfvYELC0ozhV/q
S9jP7GTo+41DRVi8RGRj3qSRq/1zTru95brxiDRKuew9f33cv1qRyAwy33po+ERGNwBWElOoO43e
UayJrEmwQSj+2cCXLT6OKOljMYDwkV3NM4vTg0vn/YL3xpWCwz6+qM0/DUUZYMpUE2xlFWHWH15J
hi/AsTdttn2yoeEZfcRnHY2dHla+kB6Uh1DbPBL/u3raB2BASzflavsksX4kNiJsgCJZBftyA7Gb
G9YcvDJUkPSWcDC4i5dDyLjBLETw79I6+pB1pPSz4bdAJvBANkBlTkyoK7VBnuE1gPJgoNm/3WzZ
nMCMCU9qLrG018KcDYgnOPNX9ctVV7eryz7cysOp7JQl/YR2mxqx6Y2fJEqWWgwgwc2S1Ar1Iis1
tM1kEz1oyaTzcGDOdczh8JH0Hv4UHzchB6qZItyvSeh65M5cyBq/JIj21/AFDc7rJP6rsBXch04O
2o30WBtHDm9fQ7ysQJoJ5PsLnymB1Jod2yYLEbgC1QbLMsmL44h9gOG++wPqhpStRUJMSUFrlwLD
1DloTWzuk6ObX3fzTo/4UQKnhO7ZL2o6RnJNFckXzh6tgoeiB6ws1y9mDgF4FMEqXOaHASC932mC
MsDnme1G4Aqq5kf7m2/8M3E15dKAv4qWyduoFau6BPGJ5s7T6JF9gO1vzSdMNV04CiDqszyxvkuC
BD3YZzQVIt11pUO7zdnjDzXvt75ZsQsxxAn5r5i6X55k+5mKPd6DJl1JM5aVg6nu+IFA+qPY7Wzj
PNwFdT4+xCj05/LQovV13Mmfk/UT9KFcFcREcmElzb7qqGl5ebdJg+NvaXJLciaOFy4beriCPHyz
XnuMevy9OcZkx+BTKsVP86vGR9I704i/exYqrRswLmGs2Bb+JDdMECKU97qPHnln9kSqhxuL78ww
DLwMGISMR7n7lg3l8U/VRsRiV+scVDconRYjYlPkX9M2ruZwUHNOdHWVp7Cp9kN+Phmp6AbKlkX0
ltleL/AHKTleV59mZeYtlH1EiA0OPNfl/FF9lCvWXlh+nKl2WOVn65hBGRY800bI9KyPKPCqMW9y
kDSv14Vihf6FYESKWiJ7qDUddvZbcCvkv0DpaQ6x8mRaziKvp/zyo0cagw5HUvWDJxfS2fsR9p5K
5Rx3Ks6uiCDVodV++QVkgqwbW6XJPgIVBRhJ+E9Wy9T5y6zThgnrhmR9+PDCZ8Qetiyah7bE6g97
AY1j2QYljOojHAUTnp8rEHKDVRSiwKyD+UjvDVmSWGCxSV77SiBxm1lIkVfMhZLLbM5qlfbYj4o2
Ynwes21cz0zEynpnz29uut+G0JgLvpd68bOc39YUErLQjN6s5he1OHm++Pni5jsTaUwcgBS7u5M4
rrEjKmZuiyt/yBKMOgLUey8hSCZ0oLuljHwA6aDIKTwudYRxDZvHi76gVwSsTszLh8ruwecfBG/r
IMwsrzN1cJ6ysiBbMGUm6Sam5T+Kwl1U0/g6qvBjaMPRsTwglKe0INaw+zlWNmuOSSj0zJ0JEsCZ
DW9Ne5FFLetNR6zU2L9IqtAhxOUnE3CnHTP5L6WG7BaRSJCpy+hvX4OyqfuVwZL+4FT2CZHdnb9k
vXLcFyHveGGw8LS3wD/jhlVn6fG+uX4lzSDHzSU8pO39fpq0KXxZukrcTr4Hieqm9ijonrb4Fk5w
mu87LT2d41A38Xl0dZFBGL+l5wKaeCp7I5fRJmoRDIT1/9ZHwxlwiMkcsqhxhAlUWgfmydSpxBot
xvSCPzhTdAAzzd8JRDQLc+MrZef9p5gmfaBY5TWdoxiBWjR0kst8aXCU1odUi7aeS/lix7fsAlNI
GuXfqKGcunBedU16R+Mac3AvA0jbcT0UWBAONECTYniNRyCnnhB3kTFrIyaKBxhF3fZ/54ZtqZ3i
HVZLtp3wwzNsh3fBrdLWfbQIdeTNG3urKnYDprieMqeYRg+y/yTMtgA1gLZk7ZyVXENjwdc0LLuD
GW8zU6VM/9SPT6GiexqK4r7c4NLP9Y9Z+KzD+g92NdjUD9NPje7Mvcc5DC52cdbODCTh1nesIhKn
MEyufF8UBAT25UBzSFB6YFqz7BX8ap6vNiyn3tWRU5BjXvBhXZYEeXCy09+5CDGO2t0xn78VgpQf
i/5US6LcNCEgXd39232nVf8KrR/w2YK9Fsg+pR1ca22miXr+9ClR3lbu82uixNWcIkxI8redwvFy
+EbNj6u8FSgZzvRmbHhzvf7PzIUMC9PSqtcV1YM4QC5ffGmBXwrqmPKB0gIsE167GG3tbmOV1wEf
u80F2QFiBc8WX7ZhWAfMFufdkeUetiNzi+cfTbtqUyq6RJMkY21o847e5eyHljw7colCtx9pamOb
Y4Wc/1+6uDzQ5dxdXctBlHb8bPGfVT6qdMNCtCXaXbzr96C/dy6U7YAHSYnKP/tsOyx74GIyhg21
MFknHIlMF6OVYXA0Ueorn0Uw6G4kqcGtIRmgsCFX4Fg6tqPGojJjwcBzObwiG0lH+0ivNDRkRFlv
5IJa5sUimnGnPs6jn7/iQ/OPT0Ild3T+r699S5oDRCGzHrNY2LYLHSNGTnu27DF2X/3P0lM9JcCq
k4odtZQbpPzhe3UfvP/ukVTqk+WsDdHFLG49cyQLIAnYv7ZBTjHCqTm3asVou1X789U/wCk6RLJb
ojzeN1edHsA29eht+RGKX3Bgzn1BdxpW24xhicV2AQ1YHxkyIS1fJV6GAg3wXf/5lBogER2VE1in
fzYkRcqBFtqTchQWVtqil/dkr+glH7h9QmrF/b+m89+a08OXBVWJ6pMGnN2LKiKtp7cqauKNUTD4
0DRG46MuT6u50U68HR62v5n8/u1Ab/LHa/ozl7Y9meyR2V/M9Ss9EfGb3j6WKcpJUI5vacaryW/T
y6emJKITXH0wSLkQ7jmt52lL4I9TfbjELgs12/kqj85NVYt8ANRHV+omzwzzSms4tP+jzUL4SsNX
1Nok87ARUQZhbLaOiAM/2W6B7adu6du8QI2AhbbJhSFpK8HjyqGTgtw5Kjfuhh2bJHguokNkGad0
2luxs+moBAGVygsgyQ7IrnzUw/PcbCUS5OTVxqQPqUvBk+sXYRC5bddiPQeveiZdivUNayvg3Xzx
mq8lRpaQ2VQNodfpzcrZ/dmhbJ18NmVB3sIRum7sGk1FnzJ49kILH9cTpbH4u7Tdrqe1x+x+yKDY
IJ70+4ZLx4HBXt/Bpdw04XjXfCg6Eqf5R/Ofczj/sz9WLuwvG+qki+3h5PPHdQlMHb93LM4BPjtW
1IPsq9wik7Nz+WBeOP2IZFCwg+lr3wO/AIPG98yUc9G9nSoMo+ogOpoXExTE9bFMVtOZIQuNBANr
oI6gtLdsiuhhePudJIR4RwQqEW6HWm9FRucRqHU+6NEsMuPBPXhXY37hKvHufgciC1wbQOdygYwP
AKLARc2vahbBYDnVOjDFSVpyi7MbwAHLlPl2Q5xG+d5Mz/GZVWX6QRcaO6992rokseSj+Z08GXWL
IUDDQxaY/2oW43ti/F//dhooF7a8q+fFypcA6XsDE9UUA0ZF8T6IOUs63LHZmDZ8XOlypzgmgz5K
4cAg6iRkO9snOOAmdIhJQY94jaMp7R0XI3HBuhN7ZIPPMJgSP6SnbYe6xFclgVXqjWgZ2V6QUHZk
mwHEMPeAYG4ti3AbntW46D3/6pTpBFSrpmiDV0A/JQwhAeknwZ+7pMPKt+naXxwr+3TNOM2HcCVX
vEd63XpozBQDmo+3s+6ei458orfWb2WO9FE6s3TTwbDGeaqQr0Nf0J8OkCk2Ypg9hImAfXRxPMV4
wA0Tozpy6wL1ZMtPYzIZ5EleUSoVBN0OufXeq7HpHHsHQmQuSzsCyIoDe8lPjx5YfvhGsfEJT1yK
5Yh30dnchzOJSWj0J4FFyyTqVdLrmXL1OC/RFgAurscxkova/CAW+y1ukk2TtKGaWCl9ePN0XPPe
lNIVyHsdMutSKzcSpDtqRlvo6iE4yyU0iu0aJxTMpelSDQl4mgnK+rQxhhdnZ+curNKnRjt2taEE
fKWT64jCprXhcoYdz9VTc0rppYIE22ePbuzpQtqf5KFw2vystXTrhSM8AD4XZdpQLutvC3i/DqvY
6CN7kYM8+zPZ6SnojUs70+F8pAwLbGOMrHRuHb2YqiI3gIy7WiCi2E/Oq/ugVGAtlwrMwaSEZrx+
z7hegJzuAyFnC9EshcL/+azXG+alRj7UcB40n4aR86NSjCSBgllpTc8NU2eP9JGSGopmvxuboVwn
Z/x90q6Q15sBVFRI5Ohbhzkj7SaeiSOnXA/K52WhXuDaBu3Skr9UrbfzY/CvDuyKKrgRliBcs0lV
O3/WRgGLZoRvGZjLnd78Q+lJuAfxtWedUTaroLinFDz4KUNPCyZLTi2Ml/TS9hysrehhsObm9bYF
NGZlptacDLrj7cyCJ2CTzPD5uCLfKvfb1pbGtVxrJxESnGjXxchbL+bY2tgyCqvfbgGuHO8SRVi2
oh/yHWlz//JvaCwR/Krn8Y5A702BzQ9R3DYxjQsZNzb2rg6kCXI96kVOXLKdR2mSJqnwyfNpEpuP
uT2Q6AWZixB3EnjCSWQJ6u/kfB9lSIWJnRcLBxCfjuspl6/jb3iaTfJyQJmRAuLpwLkqoRrmlB5Y
vthYmBWv/+/K6yEom0HT/n3swYbgYBx2i32cSiakBnBCqGdXMhZBbpdSaJkaRcueTsAUSjgeJOt+
sZHLRlq6hrKCYen4cEHButrKw4IS1BvUyk7hFg5V6X5GQBOWzrtZjMaltuYywUK9vR7sOqaQCqnS
c/nesQVKXLqcVVJkB/CqhbUjQAbMnIouObh0WYbnegXsb+OqMKefPZGN+7aM7ott+c6gfL1TwQaD
nM9eh7yzGedonxIOM2p+UKIaZl0wDrQ7VHmh2Q8wj62DQvHbl8TjOyQBvYh4IDL0Jc/7uKvJsj6s
KxSps2DOFNi7cysY1TmtM+roGrJ9K6/42TVMlkpnupZXpmdqFUpSfR1VrVGcXB5+zu3ClWC0mquN
+hCHnNQL9paY3ODPBjlhvPNCxCBUoqYE8PZw2a+P0ij3LOJDU7vGY4N1emkINSYeHY18LtCgFmug
nSRlNctn3kOeB7Z3rbALHgJAjksK9yMCoQ1gtKPe6SWR8p25wdtiRAPP7XE70SMYT6nDHLl0Oj9A
JhA9JnlrbSEWQgY5GMKz+cY/T5ZZNW1Qm4NNLoUfbCY0fc69OjOQRrTQDPukr+YeG/Kf1un2x2AY
J9/fywYZ9DrKrUMNWoLYbTVVV4Lke1r0TwX2dMcRX8WxDy8VwvjJFgDA+92quRrfgNL10wl8jnKO
szth8ggfPFqLOR9joF1bVLWGFnXCL1GwXJENKDA/aZBHbFpTesSx16OemfRFJghq6JOY2xQaHR8+
/dRXYzDOOPxthaghKy5gJm90WYzB8+Mm6LLn4XJ/rsInEW1cunnxprWl5n7iXi05Njuzr84WFVHM
o4mTKDht/FVKMQRtgURRghquqejnloHIgvmgvE+XlFKZsZgIRI71YgFm397rKS2OQBCdBRGtI5Mg
pxMaAQF4tbqP8i5nurbNMWJHTOCnGLvjBYk6YadtK56t8vPdvveOpPpRP0rUociprKW5YI2NaF5p
PV/30+r9HP0TlWZOPchhspQOGB5fGi8dt8Rf6iHNjnlh9xA7zcXAXaGINsfGFzL+zqJSyZ8/SRJB
DMS8UafVHm/VptS9mssCHNAkw5495+avqeQhV5Vsi1+80QyywCs0pfUAnbLIW8Ah/XRzhDvBtBc+
G7C8TuHZ9TzS/pvLinidle5e3WlvSv7Gy5dHj9+Ea2ni8/O6B3X+wma1fkuD1dG3lZjYeTbBI0CP
QCmHdlLGlwACLSk9aL+FRRQJG+SH2O4PKJJeRZuUEWUFFoRLQ+UUiU0tgTYKuEFnd7c99Y5tJ+zZ
/8oBhW3REEkw6kG4TzV9mWLKdNNHmTpauMnbTV+4KaTKgwXi4rC5Nto31VBekqiumKN3vLP1wLKR
iiJxWrPrK4t+jZUbZ1+Bz2FWYvNbeUUgCjLNP3m1SPnMWwwH0Qwkm8ZbLGQpXexcGeBkiBEnBTuJ
KlYbdO2ZHeD++V9FeQsQUgTLF3nDF1SkW4CgbM1vdB6Vbt63jeQR9l+fO+EZ7xQHLPDGbLMy9pU+
ecl2EbxWDkhpReqi0xGg304rlNRZUoOcZGBb2iSMIh2uZMxIntIiTcgs0pxdsoAYMPtZZfvA598M
UlxBK4Ky5Azu0P0dkYinSMiAud+kclmTqJ16tVq0lPew9K/bQEJJp7l5ieu8ulePx8QGPymm3Sgo
OId6lVr/fKIA1GJwwtWHpUE3CjqmMfh6No0gGih22G8ezgK8Tt3kQmXvam7U3x7919jrT3EqoKsQ
A6NfXtXu3ESLG945I0Ogz55oBqHcNVeeEm1ggmIxZju2cJRbyAnxrlnBDoCSJY6LdppA4rpW5V8h
lc+YukK4PwsHJNsEjYWwAbyxQ1lbgQdytZ2oM6w3rJNTmXAsTiFlqgSl08ZMgP2/NQ+j7YoYEEut
nsgi5bThKZIBJpPCmRrXVzp88YwakTjRo7Ewh93gB4Mo7BSB1fA5RelxhSXTI4iy0fGyT356tXII
B16XddBl0tbBQKmoEftci19Nt+yOtYLQXwuhOOrMVZkFL1h/q2r6rq/4A1LP18rSU736G5fW6Q8I
BfdOmEFg1a+mj+2gEDvfC0BiVMzIt8qGyIpXslexS5rq1TdjNcX1VBCEuQN6L0DqMoUgDrQ1VWK0
scsNSK7ZC03CGdJ2C2xcR5uYQCj2c2dauUJ+nEcpx/yOk7ofiYlY/b1N+M4pUeJmHd/9oKm6JkCn
v5gPD0Iv4SjMwRLVnNil+VailNmEun1UvGEk/vmNXVzJe3+gR/GR9nsuhC08h42yFwLSpSfuCatc
Dm6UPAFO0IKq4FlWCFebUfkNVQmoTMEMCoaeV6SdAyft/CCI6KmsrB/P+jqxVBwBxFP8zVLc4hpV
Rn0SOSesv+ThVZnwGbml+tAB7/uUrUaoEnsICa0ilermezXJwgGaEA66EKnH1A3aZ0O5yKVWUu4q
5uw021Oe1m3bgyLuYkVqbzEb73htwB8o6TpTlXS6iGs4lStmFzYcl8DNAWWP9lJyTHvLOr9mFidM
iB6b/J/ih2X6GQiQxWkZUx06V2lt+KbPtpZzUz5jngCd8p0h7Pn9W27d61/5/QMjgSmjY37VAYJQ
7suaoI+QyMp8KH1gkNxUYayVbttS+gpTODhlKzYxhsVX+QSfCiOH1cnG4fJrBz6F/W34xxaUXcDt
jUYedTT20Y5KCdbhzuULvP6uCk5kOqjRiLgyednvNWJ30f6x3/vQNQZPzfUTsQmRLfP7VzxIj+ju
RabBTXVs+gVK1J1Zn816/DE3FVnb2KYyRR4IhZ21PMcwn1mhOtrc2Rwn35lT2irywH+T2NCaXcxS
SRACe2YzfaiXuQAM+Yi53Qv7VfI8CmfLXXFuAhsa+W6VoZxRn3cnksKb+7MleWD6Xrb/n5tf+eqO
UilQbgRvVVmaebwItTbYBBb72wLifjduXIrkeUuZzFzR2o5/b/IbnWR5ImvYQDPInRObtzT1iWiO
2SroJGDi1SpwiuOa/jPqZTgSS6Zc2FaOYq/X7n+KgpURjIGxIMnhqUBeALNo4KTGOkml2bfJZW4/
HVqWzprX+HPpvLZN59AIv3xciOyjIBav8N4fzttyGbNWx39XVnJRROixl26Q5sdFcEGdkhAmud/H
nbpqs5njVszGOFqECaUdJtvcbj5aFYD/Y3K/0KHaxVX9Q/JlBdMQQM2chS+5zGAUQq1WObkZ9seb
BFiJT2x+e12UY1xcCe8Ycu/tYLed5F89P1IRZJLTF/lhXPa4rZJO2WzlRb0JD2RJkyVVGJy0BSXB
3m4UoOAGfc6uqkrJGlgLhyWYdVeeQacYyfdUkNPfPS609zCflMWu/QXItWzsAobOksvn9Ybjema6
neZQE2g+nTIIsers2HT5pIRDs999ieypv7oZhw1m3XCza9uGeHmopMMdhtgS3wu68V4mYIA2coMN
iiMvM+F6DE0o3013nfvrnfqScYXcviXGcE/UwzjlNnzheFe3NEmxtvl+ADss5zbQh3rl0OHp8VUN
wWp40UbU/4OlZlmZneDxBg+t41h3pWUQZcA9a7PCse1hG9AIx7Ky3VGOGetFqoaVYQjP4QhOy3Kn
eC+VjL6bmLIX7ZwyKvFfp1j+TTlgNyOigwcGxiY0PkQZkSnlpoEWz8VL4PpgxS9c3spOnBc+BOvL
Xgb/PLejwkxbVXjBMqkD0BYr2FYJ/dVkskim3vCIBhHLWGTKRDHPPb0VcHO7Ao2iKoMqUkXc+Owd
lkhW94lVCAuShh/3uJbvjCuxwT3s67sT/rAfN0gXc+7/GfSwEmVVN7NTdGDUqRzd1EjLeyb84NXK
gRPeX9nUbXQrbLMKUz9OIjFcoSRjh5YEzMJYSxsAwMeYtBuuffQuszqcQRphe2YgG81ZUc9zEVPU
/EkpjrJDQUnb14YA5NRFD+BAwMKbr/pKtu7AebkllFVxWjCeXXjaiR7uh7yrCibHvKY7uDEDpBrw
DcagQp48j8ztmYyT+9Md6Rd6P77Vpqvvm12Ou+I3Kl5CnePdF5KFLI0YZjOf6ntMfTN1wOXx4T2B
qCWU5IEaphmoyz4Ck7VTB2P8tdH5bgvN8C/Mx/zPvsb+LkSaWSxNqwYWh9Vs9Ziqnl1PryKIaAAb
KcPqfeyE8MvXsE2pyih4sL7pt3/gE9bs6camzxngGvFzpjELmBHAiNGRq6bsvvcleVxCGsAScvCO
Te41aqZGbogpLmDVjsDBio17CyThkDkp8fJfiYZXciqVshhMM2jY+BYnuZUAaUFH4J7N3tMAC8Kx
VOZm9TytSf7bxt5+z8WuNkzxhWCQJy/rMZ9aNjOkjasMdbgCe3QHA37bJT3l70WHQuebE+3b0boc
Vn3K+PAlTj3lD1MYn8dv6LvcPjNjTTh7szvDw+E1jWTXa8TrzVhMKrxexLIfQl3znNzVa1hj5ZsD
+knLHSdD9SW8U76Zc0q6CwjKjg1Lu/2p71Fn4sdC/nEJJac9OnoO8TFkX4HMFW8HxtZzwjvI0Is3
f+v+6G4A+3T4WYzxirp2hnkCp3aNjhR760ldDnWbE73E5iKgwpq+J96rx2jdPgo+ZNrvAxAtcB63
WNDnU54LJ2yRlhFpWCQhqafBtG47tqlo/xTmbLfQuJi2rEv1z3pUvw0fj/VtUqoHvl1B/f4EN4mp
4/274WlfQ7LYLbZy++yN61RjDF/Bwh8QVBBAuqhMSyTxobHrxclin4k3ejmMWeo8tUMSL5sY9N4s
jLpCqQ36SViQCSB5LVfC3wJ35LpsMCbYHGlyYK7dJJv8aVWXI0TOi4Ht0mtUkeodp3y+og2/HvQo
o/DXjf5K6LopP4GLuhC4uS9mvRG0gHva7qRe71b2IM1IgAFWJj6zezWQ8xa7Db6hP49ObMgwwr7+
wIqOtD9H12GykjhDzZlfa9X+OQQVcLF+nV/Nu4567uX2r0BY+5B/2fUkC3tNDlY5kzV60tNrGWCK
jVmgTuXfOee3cjeHTRGTmwPwKtIFVm0C605UQSVU0s/taqSEi2Kh6czZd4BtUVx7JJexG3k0Yv7/
+cvYJUkBbBp2lsw8v11+GLz5LIedw/8k3qEBSp1aE2IS/GEgewt+JzmJvQYbSuLgEUy1XsIUw/K8
IhpJ9Xa0vGtsAfif3FQFfCTtNIWXsEFyiIKeNbQitIGgpXJYj1jNl2MKWgGxTNIPjdw4VBkz2Gg1
wg2b8pqXW+6CHMVfyOESfzYOlvHjkwQH0dfbypasKSbbdEicKeZo3VjoDAaoXBLknVsoD5ex+yJf
AUVB32MAA6neuWfGoTC9XaQVvRwwFSxO6Krx3ePMkRvu7r2DyLJJPEDTW3N8xktckIxuLxA6FIhs
WJKOtox8mAeYRSsVaabCADXgRsOvm4c4o5rWM/Cqh+myAAWOQ4H3Vs8KXHrTcI4z4LbCpfn0MM9U
UL0eq5wW7Ktx25nCWx7J/WxJctiw+Af08tVoGt0x7yKb1Mpn5JzIAy/esRCPCTb3crruoOZZFAPv
pfssY8CR5AOEg0HkM7OQjoGKMgU7Badn3V1ILTemvJnsvON7evT8uUMJpOoXxv61U/h1v2eOLVRH
AwTi+Y7Djg+R6KblaIaWmc9Vj0LPIT/rmouig8yu9LI5UeiVIZLkQnttNE0ri2pxK1MGq/BKwXwR
5kS8XUMwviuQMyDE1vaO2kYFk70RmM03onTYD4+RlCSmroOyeXT+fxRiEsF4ui+quBb9f3omOVAa
djbtrTWAzUnji00/Rd+UtH9fyv6syTlSzVsGBavU7pZxxZ5uk+2aUYP8dhj/eH7OY5q9ucboVt2o
eSrVHn9OMNVr9UiU2E1ahwsgMu/zmBsNf2RGiuolYIip7ZtiPweVJg1CYgrLfcRJe2a89jcSUQpy
lg3aeqjw8az7b6Z4RfYpP3Z6K7uD4mz+bD+FsW4ItV71jsO+itPtrYCMJ2gkB8tuGnMreJPdyBVz
F9R6rqVqpu9shY8oXzgaRomfqsO6+yqeE5ymLL04BGDb1do08ss5Kb25U4faMM4R99ot1X2vHvPf
yqFCvlx7U/is7x05/vZ8F/fMG99m9GCjbS38dPmcYDkHXzf2XmpjwG1EW41kLiTxKDnie2fSDt4q
I5R6glokWIqwEXYg1R7MesR1LJW+CKIEXjLZUDA6sNb3Sxjbw6TTGJ5xI+fXMLz2T1FJhuf/jf5o
N5maaoiFRt3Jc2f4tx/lOyfsSTYBJiNerC5DnBOvgV7O0mA/TVVgGVpxscAvz/mMRARqVXT19v4a
pSfEejLR41R1rKFY3rjjJVKRp3EEyGOp9TwAAF+k4cmbFuTaE4CKvhlR5cEDfojnfB/MX+QzbXWS
0D1Dc1MTal8uvWKI9JyGV2cJrwwwi4q79FrofxR+l3HeYvXJwQtLUb1WlHIVJ5RWn5UD74tUBFTK
O34fRVS1dysEELhVNElMDvC4GkVENVKwuKvtB9Tn1Qtl468nN+wt4rUjvOMJwidUIV8hb/UfxzDl
S3YL0X7aqBtvntzym2vB7pzCnOLr2ejaLsCOMW4dpyd2Fbedm9s/7NhRiqPShmKYE4S8xaWxXDyq
5xB1hFEAW5s4/Xrryo7kMMnKVQwJ6NKnHOONGQI2uuD+DFgyNeHP9Ddle3eSWfyAsZIPGbLV+C6x
xxewOeDBB/9f5dd26plNlgCsoHLi3KAT2qmThR7v1NevfYtbPw25QgRto5rK0yD2vItmKb6KBc5N
TBH/eutZl8VyxPGapxVJIMlYNiWwweRvXVLyaFbUC0go6x1YwW79NBdbGC/BrRCBARhbEeIEelcQ
FbXS2RkG+8i6381P4P8iXC/5TZqgRJgyvvGymPp939f+YktZh/ooj6TPo6Odz9VrmH/d9D6fyMhT
Kl5blaRSwPXQxO8eT0X1DnYc127BSB+o4GrJjwt3fS5a+xHPAGYPNr077X1+/7atSNPmFDjhelxY
W5S0GhmJCiDXhL7FfjCMj224QynAVP8U1c1DMzrJ+WmycBs++FNg9bv4tWUKIy/79D2UXkywaoxV
TYn4Uha8k/Py86+qABP9EQQRqejyWfvyMkFeHkB5vwSDilLBR/T/k6srE+X6PfQikh4LLfzM7jZP
LnsfKiXjDcmr8jDhP/2LucnOe8zzWbnUgw9oN8FuWhEgClgcI5vdqmAZ0pIcWaNoZzi/6AF82PBm
du/ye+kjYImluxZhx7ZumYhpxJewThptvCSUr7B0QD0djof7IkdkjYNH4cH/G0ZkirrGLUjssi7k
96xHMneHBBjT84swxFSlmtvgZNMPKTz+MTzAK7XvZ6dshzatJOVrGXTQDhYTudrbuYhxRHS5N1Pj
3LBwUo073+7rWbFctZWnSzWMGUJ1lwikJZFYePfGM6RjMQ3XUGkOA4YhYn/J3RUwcGqVEFdFLw0E
teJgXtG7ml3IdqFq32ZVSzGbjOzA5uFHL+/BxmoP4SBDzKNtpqqZpnRkFaYp0sKqwEmJDIfJkQLV
VEQ52rpOFVZoFKBFCZZxb+Rf87CmKHnRxN9eCJxfeADQ6T2i2VCjDOEWEU7R03W0towP1T40C/RJ
l9rlTMn6/2l4rD6My5vauw2YX7VOqZuMX6I+oGwOEDJEfckcgoRbWcSqyI0A1PcE3mYM4yzIgHVr
tIlZROxKg2wAiJh1n2+COh/URbwwo1YmRm/NrldD+IlhW/Gfy1FjrL8cUyF+tk+p6cipcccJsgNi
xhMtlrFGj7FB55DyBSKInhRlEJiGd1XZGHf3WblfM5z7LmB3AU5xzw67UJr+q+yPb2EaqLhcIQDJ
+D3siFN6lZrFBAQ6pASyjwTFMW9rmhXE5ilqXjJPAh0iusmog6rjMV5mr12tXXHKyTtnuuocM2qh
v+Q1rxzp4jpxaf6LDyux796E/9oxyS7YrZIxGXJ2hB7IBJKPmzzQsMw6qw1Owki0yI0/BJB9ofDm
jFRHWItEPZX3ml2LjaqxigVJOw2UC0i+tw6hJyXu25YEzN613fj9Sh/DtSQoj2+CbY6U4JXc8Uxk
ET2gJED86QQBK7g3B5FofyfV7u9gywmfa3pZmekmGO4cwpsLmytKEOI88+ZwhTaVckrbI0naMfto
Xl4P9BJt5Di7T8lz9c0cofqDYE5wiC7ddRy1h5TF3Pk7ZRB7oRGyQIp+aQPHPDvVHg31vCUAXwkW
Nh5GaE6fNA4n+V29oQ1/6aQ0e/M1amzuBkiLF8HXnXifGo70xZlHXYFecK6z3jpqG+S8imqkwYQW
WyAMm4whR8RV8rbGFceS9B59GfW7fzAXBv9cPgJarm45ABYMkd4G3nuzVzDsSInvefrVJrhPNZfs
Lvnk9OAR3pLn+mQBQxm0tE87/3PchFCHtqEF2hNxGpNHJY+6U3dzfc6tQQaYbHS5WlG+WoulMB8g
EVMdvEUOCDFaJGCoUtpftM7UQOeUXiMEJ/BelNa5q6K2NvwWZJKWMxGqhRdMTTIt8SvObD3MhWoH
HXxHury/eoaTFmEQinMYXWRl7yRP+tG34kHhGTG10dBL1nhXqbbT4guqDiatO0SCxZ8tvwx1Y14j
qWP5ft0ohruJ3RMBmFki+t2l7VzbKV71o2lmO5VxuQXgj+HFC5S6+5UqD7VokS7quoEv/lpIJV83
yLb/kyLrdXVW7HIuivYQ1jZZSuvkEgiXfAPH2Gu7T7hHsQvVMcHz75C3f+Z9su066oMS0e0OwC7+
07Ts7pAY3IKWb0gXACFRD9zk0zRGQS9RVo9eGGzeG0/JlkmEG0BT7FBTSq4EygAAI4DT6YK1TDj/
q11qOUU+JSLJ+i9qBCPsmvNpxog1mG0MJoUmlsfmMAnkPnf6X+WbZPu6zPr2HCLXayhg/qsEd8OF
dAaXSBMULPNIVMLkEJq6SHJcYifx9M683EPRTvXG5CV9koM/SpJGpnbQV0Lib7UPfeh+YmjkIpNK
UfxuqZWSNtPOnrWc8Mr3Ck7BPnSUnT9SAdYDzqDMWe+0Cqo+FYbLPTgBnBrM8K0Y3GM7Rw+pSXNp
qjcp2cclSED/6NzLFf59lSdwLR7quNzIApLxRr6mnkuWhndgTew3VfmQR8LAmU/t0cenNociXzR9
aEVCWco/maEJcdlI2GShDKZEX1c53o/Ca+XNab5eUT8YevQA/uAFl3fMv6fN0Ay2/eLUHI979ye/
FwHPgjYsg7AnXedZKFAigZWhenVP6dwuu2s+eOFjzEIrm1XBiTFurLiN0Mu8K6EAymG73SgHZ9ne
46baqClp+NsK2dNS2+xCpLLHjw+EuPfATchYipmByQAcNJ7kAKo2u8mZCJEEu3wH0B24i2qssQwx
zNluU1YrP5wCWZ9oTiP5YPaqm8/OKzrkkVNPJ3z6zVewj/t4HiXZ65LrAMi4Z21kVlJ+zyz+xwnV
XsNS3KCXdaoU9l6lOMHR8J8/fiJ88RS32p0nJkd2NBrba64iPfCTtlswESuROVlVJnSDfGtWfWhj
Of4eQnJsCVUOdFciMKwzMuduM6CmOgGumWTYUbwaDiHD7BFVHATVMKIc51TyqGOLvgv+jVxybnMK
gMZS9BSB4ZPM/spvL7Cq0oDsgP4aYFGLSnWUNy9d7SaeGUAKLkGgLPL2tOD9rZEHN1n4lZsF6aAs
n0TC53e5yrTQis+gcx/OYkKjqz5RR9uL+/1ne4+lWO6bglE6uEnV3QBsQ/LD29Yv7xtMXWNZXBPf
CAlMKJ+gw2Ylpg7jm6mVkJ3WyZa7Dtpnp3lP+Iae4Yvm1PkhPvm/Dh7ICnYl5B9vDrEnIH9KItQg
2hi4+YFRlgupFeVfb7EBS/xvd3hNnNjonygPvvKO0UOMyJyq+FkNXQkXA6tBohOF3MWFbnTmj+P9
LiwoPSorLrnM7iLQRSaM1dKD+PTTgUBDRSyqyxrgvWLZD21dy1kPBQFZ+28MukmD284AjZMwL6Zh
YNMakLSgR2DN6LgQ3iyqlZjBF91HtopCpigv9SWE5FDx2G1W6hmGhRZKzBJ+zhKXl6P+9/DBNDpt
C2lvVYp1Pnof/yQpD8fjLN4bXCtRgfYzonh7Wy8TO2yH3D4cfdSbe2EBrY/8KfKyvjKT8RDn9yTh
ccypHgf99YZAuez2RDl03A64hv5emyiXMUzhTkJQXIE65EgiDFG+Ii44O1GiJmjtGwm2oUMkQzRC
NvkVBXTXXEOmPf24EUDN6GgQ2wxADnfWouykf6N4CCNKdzRr14iS1Qx81hgIl8CLDu5s1HytLZVY
Gbty5V4iLzZF8k38OsXF69DlGCYacQGFzj5+66B8TnPoqhU88jKJc7C0bAVbLt7iSE+4NWDxxQA6
51UhTwGJkvRiOU4jC+X5N9eQXYYd774VjlNPPnb0He5mYiWGf2KV1sTKIrONdJ7UM5EuD8GbEOS0
V5ROA9Pp/Gbd2iIqUwMku866KeeeJEZXj50m8DQFzn9/7ApQOPvvayzCoW/wNQLeAJXLlr0IrqBu
0JtDBzMkqwxKxux8YA97zTxmV4Ftf1btj4ugRmjehPb8kWaIumus3N6+YxFhX/tHQEhtTMk62use
tI+KLxnhZ0xA2v5k2oYcqFkx3HdhXeGgo+7Izp4cvDEOzncmeQB12sYAp1bXJxUHQjzyOjzLlryn
omKEE350THMbiicGpq66N/uyQjKnsjq19FR6hVm8Aze73b/8EaA12Gk016nuNZnwHp9zgiV2e2z7
P8JqNe4HF2abBuPrxFfZIsrDhBzoGdjC53BUPoVyXbDofC21EHVYMdo1b0GsxgxcEdKKwx2Hhq+g
aaeEdoOL9WraXjQjK7lNzb+cxjdIrycATYLqFdx61AOA2wOmrQukVV5wJZXWfM7HF24hUcrYPwky
hEMldMloIF86maxY/Q0JInPTRPP2DQDz4jMGCHWnraDlGFJS0WKK9utmiM3S+DA0q826efYnx3z6
lHlLILMMZrN2JODTR0esJ6eVWchsB1Bk1MH4au190jsbQpemHIhe19vN3h40NrtqTBKAhouTM9AL
KdpeOYcFxjX8Acjb2XzameZHQDloss0H0LSvWIc/v5E75SCyFiDUyj9xd+NViu54phrO36sso+wB
wxWNzFN1ODiJCoURGUVvdo7TJwNhrSsl7W0EBQFUlZtmxgVaoihs8Uyiy2vOaY8MGdjekAePTbIV
7V/5d3lCESIT3xdRZJly95+y28tzYEcec33AqZqDw6pem4DHXYt6NT1KI80JjrOZLTKYI3I5lLDu
mERhpx0h4rp4WgqDjYeewzbdQcFayyl9YVuILMFDXWW+WDHBam6aDGHWDmTu7AaC6Cxzn6dnky68
bz+KqWODPO8I9OE/L66QDJoSwE/IHgAgaaQdzUKZj3vyGF/7pXgn5CiFroqd/G6FZSrg4pERaPQI
AT8qD6Tah9oF3l/x9KUGBrIONeZdIYlNwLLZ3wUnhZP6oZ5obv/kK08fjsE4PTWqVqfL+BC0/4od
/nVwmTFwWtdQLEtIkggeetjSZ2MgSSQAvwdtsOnA0hgnLSsD7UTndWGOiyy72Gv11c97B8WvEBr8
zT93lN28nazcdCze67vfbKJMGwFpguFqHHQSL0aQmgplYI7PlIPxq+TREw/pgfmtWQFW547QXrGl
G+EzFnRejJJ7GNff2N8ghRFNDRj0wkDrQG0vC/bt1BGacvgx4DaAgIqOhWaO8fFcWR+Ip5fUOoKE
wB0vQk2aGQ2tqbKM+U48SGVGHgy2zd+3XzY7xA/7g27LHpW9QDoXiOdKo3nb2uLhZBgmRAocp8O3
0d5D3JcI0noDrukHxfhIahdjH5QTK7zKhBjN/KyTvKeB/5sajIyzzJIIP87Y6Kh8SjUehXI374c3
YG0Xp7Li19yq7VYnbqG0TpynY3ixT4vWchawzVaiVFaZS6NMSgunxndXdRhgNC7X3Nxr6aL6eN4g
GA5Lh2EPW0DJV85FFjuCu2H6AlbaanjEdWo49acBrw5A0MQr3tkSOVy/cIPp4K8G2cYE5kvm5V/4
uQyBrdags67T4oXR7TvwRqKTS1FK5750t5DoLufrVJhM86C1Wats4CfZTfpzpjBXnH6dFHLUdbiu
zBgfCr7C85TKjnPRSzIT2t2EZOWj3TKILd4b43MN/pmzG1lwPz26b/4xH6vi6KHf4/MwFf1uHv9t
LYdJh7YN2G0QmPq9o3iumRsSW5M8GJzdghmtQHEKZ43d7Fd3I+6+la8srbxhtOr5KI5c85BvYs2x
5TIwAQopD2P8u401BLaiEiUf6SkR8oGisISQW9WC6FH/OlCE2i769NWscO5GmDen+5bexgdhdu6I
F+94DbVIiPZ8NU6YluEnoc+czdLJQUR+lwan1YYZn2l9HOgcuFu6i8RMYhsD2tpqAjyZPmIZQRMG
vspHDcl0M0R0F5OSg0ggesrzqKnROfMh0+V6BteRl9MczQG6Z4FC1K5mdGMiZ8VElcHqs1HZFW9p
G0OAEmcJ3HVlqO4GQuTyFdyoZF9/G/1AQHeswmk6cReYgBkz+VHRKbS/70bA2iJAfFUtDywaPdyp
a9EWy5eWVbFghRxosYPxepnd9DtCryCwwyXIHD3JeODGm7yYVAHa5DbuGTYHLygIsf//UbbQb9i2
JRPDzEvkDElRmNwEWzEjDv6jwRlpR9WUarIjWU5lE1n5t8AAaWii+4hljODRlVpukNeFkX/5eJPl
ZQhTFwIULDzeQ7KuHSiU36VDMOnmRUVU7icM+p35gJQ6U74dwVmc4UA8rs3HCDHC8HUX9QTuCskg
e6Z0shgpzAc3LK+6aYNamA0aBRKrWtedgmj9Ji43pS/UbisvmDrNcxE/HXYcETqFUOiaZhkpyjka
wpyTRI6Xz1UjmtyDQdhs+HDGAS5SlWLzFGxCMSW6EE6Y8lvkIGBBxxsaeYT0PClCldS5v/0nClvl
TWbxcNNvnvJWdM0R6RPfjEYjfcJGBd6PaSVF5T4qCVgbXg9pa0pSoPWWc5cLDlK6EMYmjG+rQYFq
bWP4aLB0OxC2AGKrT4BuLNtPtBq+DPTujuQFf1D/0AHSKm1X/Bg+pIuoeRs2S64ko/OBxqUA9mHA
gEzSS9nGrhWG227ga4zmhHRranaUq5F5YrKp9bS+NoKVVScjOgqYVvQ49lqCvlAw5LTjSmLkyFSQ
EykQ5P5o9BSsYr1yzOjRtthTTwpeatNc5MYo29axvP3TDyLIPfJ7/OxXW7cQ3YE+yR5vXFV/ZyeN
ewul4p+QfMuvMmHX7bqnIbyh/AT9FxQoASOr+TjHxLQDUzqAk1g6mcIeXlSq1h2hcG3DWmDwdI5G
Rs6HXojXolPhLK1ryHxrQuQZG+NV6JqiArp9dW8nwkk2Oims7z3N1rWoqBQm0BvIEezM4ZMRTSok
dKkwPUHmWFbRwseghJ5j6vJEffDtnCpyNaMyL3UFz2Fh21DByX1RApdaN4UEDhAtY2PXiAkdhoV9
qhUiwZxVrdXAcU5AysjwNNASDKcNkTU+tXNwIxnoV893P/NHXfMkmjPRqYgXDlqNM28zdCgHv01P
i7SLf/um5zU3Z/nTrgq6jWLw2Q6s1BLCvGaBxF2cW9RZAVj0i0kL5XSqtv5bC4zmc/3cBJuqqway
S3SgQhUEx21/cXzQeUCZcDa93dvIJVwdEdVa8pynX+a4Oh699PJIcVJOPFWGrE0DajPWIKD0n37e
H0VFjUqif/FHRivtcd50wbk88U4qodBqcP6VzohqmorFaPYtAzgAu3ramY/kOEBniDG+jckFcDYb
eW5mlzft0tbzgoUaG2Wj+vv9fEMy8hXPBpCSi001EeUrFpPt+XNaIQVrhoiqWHu8MQDzWYTcJ2wJ
jviifqG++QjMpJsxlRznsiBAM7P9Hh02e1R4bSqvTImeGLVnEq83sdEaSEvl3cQw8uZt+9JHSrd5
Uc6u8guIT8NvewgKsjQCULnJMnd9vO100dnulEn36ukPCftBsCmcf7ko3Q/bS/v0QsXJGjo8wGQn
klzG2SRj2dNcXm5/ayvq7zYaUXbtJ70fmOwuJuQfWq/HXRCYdIh8sObxPv/vNXNAn8dwGh4GUXGr
4RacWx/VmdvvAVNHv7m802qyNR8AOepelJW5VDT7ocwm/8nHEQMeSnlxjLQLHbCHDkkMmtn6fdbB
ocEuh68dH6NW+QVmx3010Gup45BKu2cux++3jv319esyEuk3DoF9DZhGPV8dn/npA4adXqlye2gr
9M/yww6GH2PwXDDxOMG1Gre9+IGQMvkP0FuQ71PcXjdNAH5i2A9Hd8zZ9rdy0Ft6dW/TCMqOE4xH
VwykV8FwciulVycaM1NLft5bb66Anbvqqs4Htokqbl2laNahe5NFQXn6gcgFR2NXc2YgqIc4DXq/
wR+7TdLOmeW5twNOu2PWa8pxtRoaGVBr4+XFpvWOMWKr+FCEBXH7jvKOOqkXgiqWT4uM7kHnZ62E
jM1wzpTxvx1c7NA21ka+9g7c1jWuS3r394HH5PdgNhXkTMaQ0OYjR+CqUE3aeMdVKpv9gwI+bVn4
b+5Gefxb7bgh/5Plr0Jyqoj63da2Gtkjt6fL6fQkVDkdd/+7p/omlHYJTyVihIkZjrUeyvjvZpa5
4P6/7ZY7a5hdjbO3C1tFfsZwLr18Giq36htI7CE1siMJF2g/usvYhWt7so36iQyZk0I8ndSTsPXz
HhS1degq+J3nTaoRCOBxz2DvqT276Fy/bfzUC6TEJiTzHfDxfMd+vS/t9qLqiNubez3ubwG9Q6bw
P/0Xd3TRMbykZweeVKwPEldSAB03Vrcbm1KznJGFnLqVyP+des155gaUT9XSmEDYb+g5DrsVTQSd
jzRU4yYxemPe7wOfA5u7VHW1nFuGUTfPg3iD/YWvVZDObpIsCe+rMFDxH34xPAyK1lbBTZPZpbXA
k1FLnvXc6ix7o8BMGMa/jrIj8XXUk87MsMX4W+j8vNiy0XIoBJ/blJdIDNCBEiJPKaTEuNS7Aruu
MNsLzT5Ubj1z5DPB78JYeOyfrlDXql+M/X3Xk/wLpXWdMmqTJeJLIFtT0Fv4vvIqSh9SQsRGK3TP
/OO328AFERmwpUjqqY98HUMnAQFBEJnwGtJY9j+oPLJNqZLCaaRsk3kQiy9ApOeLlKVHmK0hxvTa
MABCf2IjkgQko2AdLiV/BBKK2J5ccpe+nyuyBX8i88oxQmhOKF9ocD3r0stM44q+4q7rt02xxbLZ
FVwJktXbXG6i67QQpykmOxJesaZGTJWwwKUefc1E/S346BwvGyZnP44rPPf6T8yx+Rg+PoC6xHM4
inGM32gCGKSvJUMHO5pcsHt3TcvZEgbSKuMeG6Qv7dSIrRNJRdjYqPkUi7JChusEvkTQR2U/uSLt
5lckq+MjJ1XIzEgN/rb91oIy1hh9U0FdI4YhiWO9CH8lbRzqQORl0QRhIRylid9/gWiN0pZDlOlq
QCPV+gOUJL68iIk2F9UOvnTdAMAsJ5pYRsg5Ee+6YPayIRCN34OfRt7HOdxkMwbtmo3NyUbLzswz
ejdkyQ8b++0aTg7+W9UqXIfmVmJbGRRfrpL1+4ICK9ROZiUhZ1WwnWBwZNuw/Ulet1rGASbmyMu1
6iN6FH+MFvA8dZvcggbuWtYwnlwLHX7uxqRsTXQzQ+ztu7A2OjLTyOXptm4JYGfT0Faw5tamh25z
3sy5KiIda4aUlJh/SJmT16e9fuhDrdt0PSzsM7f/wIQOmChUMaz2LDJTsOeb5d7ITTc7DMfR2Mv+
E9CwMh63uSRqnfoLQysbqm23DxMFI+pdX5VD9TruF9SAEh+hRigC1dO2plimXBWUoO8iaE7XAqGb
zsMgfGfY7j3uBOe5R/F1mLOl32Z+IWV0jvsjQy9rBfOQJOZXS7GFzfqw2LE4twkkl+JjL+lgCXqt
JZwJmYscpOW1iIaw8jt3dNrfQyBTMdavk7YWGFTXUPC/miTm7XkpxtOoDcMmQx1b9ccJKIR2BNi0
tIqAFFhE+0H7C1KHTqf0zV2ASB6Y75+MX9jwYT1bUYqg2Xdse/O4IN6H5h1/BHJYHMXySpvFVrbm
yFkiJcMrJeccl59KsPA+MCj6WOBZsDcuX5W4C/SpZGYOBwtIqWXhAGm6vmBrKD/tySionq8oRCQ1
9FL1wOLCqyMWgzGxI19fVUUsCYrHjWYLn7zvSo3cZqno1/aEnmUahzAwUw04fhQ5JrpdavVkd27X
mIUMUl6wvr9oJUJL3bHMgfVcN5aNzg5dCU6fX1ERHUWwXIfj6e7PlLtcRJnVkdjEtQP4ZHdQZcdn
/q1VFduR8qgYbHT3KA0MpUIFo9NiKNHtj9Wn1Nyx6/imwl83WsfSBT4AhScuroMZjV2MpP67yTEi
K7SJbqSm1JffFQ2WEMwJPKwjUU9eAO6BGuEbTpkJWyWjX5U7pDWVXwousdf5JSQHp/Yi3KNa6Yb6
U01xu631LXHDCT+ndJCCFkwrevP+hN4gTBv45opO/r9TKiKggjTcl9v98mIwGSTqoGy3NWMSnRr0
Jn3TfJtC0eZJZ3KQDK4J9OvCPkkmNo7uFmBcjcB8OlczknmQPeFFvDT9auKPrv5mAXXOWOt/m88Q
+7iK4u5JZWKC5bzPwBCU2kMuFkaEbunNHKsNjydCS1WUF20ekbPmvdMqG1WOZ71lFGKQt2jnjpIw
hHBHyZVEleblpCNFmE9aTq9pROFKr6aKre17FVBW2huq/D0nK8NHCNYC2eTXmGs3MLsNUs7q5nSL
F/MWO3WF25M/A2QN+INmEkPb/2EN2WJgze9FueDZ+iJ6ss+leqKgxvTxJnSsmyH3MGbm517picW/
oU+Yn8A8xqUiueoAERvWk+NmOJ9O4hTI0LacR2Xj5M7SRxBhgVAe8gAgHuDTnv2PAlI90fYLfiUE
R6f/wETjjLQ+qtAi/kXmPcT9AqYnw26bu60yM1KINUFCapuFbmAsyU9ootl2zaNDQ0hFpZpbQPL7
SyGmYPsdlPY5ImWwIk9EsjZu6lgHDGrUqmh+hzD06Zp8gShpxDMeGPflLwqrL0VafojajX68VN0b
t+XWB+AQsclsBa63kq5JrjyAxWOL0Dsph6LifNUI5nvimiV0i4SfIFMhpT032LObACPatnOq+WoD
CJgNZHSD5UcP5QkjhzkR/hk/URVWHd3PRsnTpdJde/lKQilrdnp2Qr717mPVDg4ECELzUobmtk5L
h8+SWO9fRbGkHLkpqRUtUKZSbbvB6N7CWXV/iY/UElV+Bt0ebuBYGJLaVfZ2JHD5hd5DxkH7CI0b
yeLyop82RfjDr4QuhaN4UlwL2pmxrG0P7b6ly0JLMZkrNiZvm9lUjkK3SQLHZDca2NV/RGSdu1JI
4utuZrjGX/7EbcUMPBXVDGOEghITZscQMQrIuMsoNf7V6mSZzubBD18fyodpxy0tAmOO6CO39Kyn
eMuIl1Ew1+lmrb57hosqfVBYFlGOzHgybKQOEZXZqS/Ik7YxbpCzwKaQWOHLy2NfTBVQXHLhqQnA
DzPd6efSOluLJOO+7Mxphj6Nm7I6JhFEuMlRvf5Qg1AHMdEtOarQBiiD5aOaRbpcc+QwJdr8wWpB
xkw9nifpFdENiHUK0reFxBZMbx0pq5bDQ1olDTofN28wq1gRen7SFvI563KwMML2LdDhhxK438h5
ZEkquLfByJDpcwj/A5aQ4elXRHS1zBKgep8V4dVzREp4z265Ffn3+/DdsfOPBVOuEqOaR7rkptwy
UQo2cwq1ZPIkhe5H+e0P2t+1G43TYojRwMqQo2Sph0T65L1UoZ0eNJKQAZEfQOmSKStF8JfP3tV0
CS8n87oH2qieOIibTFPgq7zSKWjYLy4EJdmnAlT5h6JAphF+epi/h845PNzOrsucCsx6tpgo/h+d
ASsYnvPnXJhwhzIc2YJNP2nr2o7L/8Eb51jOUfJTbWlM27WHeXQVyutzUH1ZMUC1PcPsN2CkrBtE
RZzyYpOScXv75qY+Q7mAMRvP4IKf+wjim+SqUnEYJofJqkB1O6nmM/EzDIZDa+ccmzjiXnyzrN5Q
yZ8gc5sIPtS3Yw1AxsRWCuNCB2x8ZhHXNDuMgrsnOaqTtfbUBcYmGV7Kfutg/xQ1NUDf9oMujpCh
Gk5Iqtn0rnXYcAd4mIPmJpF5H6rs9ujGdbXsTu8fdzCC/9gOqZ4Yp0f8rjQSiW1DbY3WagGlwmhr
rIyIx9qNlgKhO23pD+0HwBPUe32Vv6gFCxbl07lcBT6stVRY6ip8Lkuc9xFXfQCy4mpECPMKTRI6
a54efXdeS49NwnkYdfA4r3mIy7KMzOnIAYptnFPQIA1sFZx7rvLPUhut461FMjCAHDTG36GnpbLg
B6UwZckufsqC0YBj+d3IfcAuU6ZNmE85YbGnnprlZKhETpqSAnyC4HIHkhykIhh6BGv/pa5iqB/S
UVyd5zBabu6fETLzV/ViUkHt5EKx07XLWV5Ir9OysEI6touSkUP6Fc7eez3RN2U8rh/CpbWlXZJO
Ys/IbCpWL30JdfxWGXhVam+9UZFPLwnfOedtQFIyLHp+/Xc1sfCPQnk8INraRzZUFSc1HI16WmgK
d1iQehUQIlBcPvO6Y0nZ5dkl4uacLVMUSfT9Np6w9XzgyL090kURnyOsPFELmjOMsw5PBR1Td85k
1Qq5pbLrwr61cG+vNK5RTPSbX6INL3ZUfF+mxZ98sNJU/0MbhY4yZhj2ckutNx6xrbEhZDKzeohd
ocyE8PJ7sTI9PcskLn9Zgxe0ETfDNrZu5mNwIUSFTNCswnkpC94tcKsFoAUUfsw472WYnV1xaAqx
y1GKGtKkSmAuQcEsaSgE7+zyxdoakZLZXJ0+ZgxGs5QsM8J8+Sy3XC8v0qw1d/FjWbfWJAIoK/cj
Rflq2SlxaRRGJxqW5235oBI0oCfTFGHs7SVW+ewLBtDOTbOzEJN19faMEx+fOwu2PwPlYGnm3mnS
qJDqxVfzCt7i9puqT15+Vk3IRR4GhaMP/Qu5BtJj7TOKm5GJAhVTmDGvzeJnYM2kpAgTLc1ZKuFr
t8EokTlxs+mEyAvWLB4nCp3SH2Kr1HB3vpBVPVIg4aCqQTjB8VNVbyX3sQtqLoSphs5nS0n2xD5Y
SAspsTVQ+KHBW9jMQudryUbc0btVM2jd6sz4Uwm2WnFGlWYHUWoLD4V2BAI+Hu0wEs2JRb7VjWc9
KwuvHjjvm4CGBblVntg63a4gL7e4q0HF+8spX3E/Xy76AKal9hTLIBfRWgV1XhpvY60GLpwOyCYp
voxzfuV4BqZUsC4RLkulsT1U6F4ylmTBS+VzcNv1qdnYH26hrrZeWIVESQOzXKQoxARhj0auNCgq
MIxr2r52eGMMpFP8wQIXXEn8wRPm5jkZ9FXUyii1wcMirWQMOJZyabmgWkuFqIZIyi6++wckHByG
2ZueIwIPBTnUkhz5t+Nk7yGbPs89qqRKFXUT/arr2LhiL0H1MxCKA/0VIFX6GmWpeE3pMgk59hp2
k8qgQshhaeLDGzX5Qf84VkinVRQgACQLUW1WtYrH+oYEA9W40rQnZ5+Ocb5Gmrlbn67SBR4Y5eDb
0h6QQ/1rjqxTrapdUn85PZ+7fXHYmJTyCKizNVus9xkAuIx5OMbszB0BmFrrj6rSd5Kq7tqABdk8
Gk9j4YwFJ47YlwnOYiiXaYdIlM2jwfhVCsl733ktMIPOdx/+935+sZJ1s2m6Cbzci2LCe4PhfOij
oqSEkN8k0QwcUEcYDo1S7imD1D7+gwZ/TtDRbKrQ1PjtEUEnOoJ7aascROLJ+ODsxYbDe/EGcaa8
ISuLoJ4w7TbSwg5MIRyaPw3cmQd0e6ajKVWsHewVDKzdSWYNzIzU2RMvSSk7690FDQjMHBQ1QhEm
M/yf2X9HdENagFnSyFHMHkOY2Q5F3o5Ehklky0TYf615zwtEu1zOHAGW0f+ztuUzk66ehz4Lfk0q
Oz5bwYfErjgNtqbAjR9Kj3d8DdKXyYqzoDHYE0aUJsExnKEqGz9xwDh2xpk0E4rRwthwVogTQSV5
v1mIDHFDTBNyeePOiyuiOSAWht9aZFGkmBIkGwDPqsSd/A/PwJjN2t4oTfIlkfF+N32r/zkSZVr7
6yRrjCdbjtuJ6ZiVrbJCxCKHbsdvSNeAUEEb2Hcn2BGxjk3Yn22s2t0bO3uBCVNduq3eovc0hi7m
aJGYneOlo3NI5uBMSqPYZgMrWyj20Cs70ckkc05j8ks62kaEAWm1OanjPRvKuHZMznal673Qonot
ftJkYaWf8AWj+3YvYX8sjY5N4ASjALfk28Bwt38roDG4vhMLAaWTP0IOF3ngN+6Ob204ULOPchOr
LoWPhsO3u0n/veaj6EBFNEjw2ifnlFMEdNWiIEnPSmTHC1p0mlSMSuNQ7WZqkDsUuimQIBYgrWio
iT/1zx6NuAruRssJ8PmuhfXJNsFnuCDJPXQ51ukwpWgiJcioaYIVWuvtlBu2KcOppte6lBk3lThe
Wr6238J2lzF6ebXuAKh8NhN/VWqsCFP08ZfeIhl6z1xnMQ02ZPbMNm+dpKNJbX1Me6DvjK0m21M7
RoPba/wvuAKJGlZlD5MBah/SiJwOhksm7QhS5twsSu2qEKuX8t2rX3jQDbFY1Dv2OPIuxXlqnho/
86EfTdOEMZQVl4nHwnkHACB533Q36S6oztyTBkPBjGDt/Oa4hz+88Veex/UCCnwiVfKzdab8z11Y
xqZzyfKQ6ezOAM17HRux9Za2yM9isPXX7yFETDon6YHXBqd8fiQNSukno+XyFE+dzqzcQRMFwhQ6
ypRS7x4/nRT/24j/W/ClsBG4KvPySCnYpx2MBNhkSai7nh/1Y4V2dT+mbyifwNhu9J0bAqIrSsXY
Uuy0UIoiIqx+bGGC0+9FF4I96epdl5zdVfPJflwiWy657CKkNBei+k5u+dAsGALxn2Imdm396pyR
hxPxlEcNPXdz/yff+rG7z0qlPQ3Cx3ywSFsP3FRzFoG7ndeCLjMGICCD4tc1aCk2y3MVYEvMacVi
2KLJa9v/E/fkxd4BgkhIBVKyCTBf9aUcq2cbvGV10+KlQ80k2/jOOgVN39zr691SheYPW/Zo/hsZ
kS+lS0igCQRYUs2/2PelWuJWLEgvHTL5C0F26KzlJwsr8DveSvQ1Te1to3dOjN4/dHEWmf8wwydJ
GQXmzRjvl7kW0vOkp5hwz0eSXGYsCYcvWmPG8FPfwqlSfSDh51nBgsUdUcI0H7s0zRLzUOYl9o6p
DPkwxZtmmzfsqCuePrJ/YMeJQQNW//UrnxaktU4ksr+XSJtb6Vj+jSazL15K82ZuVYkVzdAuGDaa
Hn9yKQWURVRMjTUvLYFLzzfXRdhR6H366IbGCmMz2eG74bMsqMA6GrujWAA+8Nw7iLNsc0yji8Bi
gmC8RUAoKdXntxSF9GzsZ29BBp7mEtyrQhQD0kgRDkNfZ48e6KGQPYAK5YPSc0w6GrBhTWi33os7
Qu0RFMoGexUnpr9oNiFaxCYYjnlP5hoWDJdM4mpps3YP1xK5D01C6sn6S5mXWNq07aktkwrZgBdw
6wMnEMHL3xXOJtSBrAlwWGWxeQyaqrXvZx/7YQxofPLHHZFYwkn1kExtc2DF4vPNpVz6MneonD32
gC8dnxvfkV0cSDWXKjorMwAEfIWFW7M0r7Lq+0sNC45lkBk9beyC6n7FM2M0ntUNVdS9FNHYiuk5
EU97fuI2HScpwUKoNynPklY/tOcERa6plTHGHoTiv82RiecZ/jDPNsU55B5jGDbU1LEoZZYlOey3
3JZfC4lohI53HeP+zn8W6QmCBjpg9fWUZufIAqZUBPHIbn4zZhSaiPqNZTFSYNzkatIFY6gQQ0wR
IWJtVW3++0IPTYyXBe7vPhJIPBG4u6RQrjwv3bDzhFNmPDD8Yfxv/lxae/aMpO0c2F0OO1uBD12z
gn08FbK4wjNGdb9Sxd4fxZgm0DcWaqJfOPPcPnN42FytpS2qniglrU+AzU4hN13d3oIMnfWLhYPp
fBmDy6lBubClsqu0S1fOjY7x+Zci+kZjp3bFslda/J3VNb8CkkukuPHlvOG8ehnyiJv+FvbkjW7B
7RuNHPUwm4rWd2eIWUgnJlICQ+dzuY5A3Kshdx+ikMbfdD8tUSjDOOs7VSVLzcAJCHVeJKpKTdtJ
/UKRtfAKl5WDGBxEaUH2BBJX8gsMK5kN8rOaBuMsw67BcPxgi7pGFtMI96/p793i9esVNujQUwin
0bnfoFv/Tb6g8CajJOBCokpk1BhmTANG8CRhv2FIzj0HFWffqbjB0ZKO2+G4tVx3cbTuuALNLwsR
7wZFEInPO+mcwK4acqsZj8KuF3pb8GHdN5mpwyyETCDwnyGEadC7VOmkSBUYB4KHGZCW1bnW7L9l
vJ6cFT7yjkXnZ/sJsPgi8QHJrEbomOweclKYb4nzWnO+ktUuibvBTK+FTPoAEpPn4KkxXgSriPbG
ZhhUN3tjcvSEF1fhn9KHMFNF0+k8QM/o7cqw/d1WNfzeVJ190BUKinDzpO3yGn5Hs82Lu8x2pgdU
/0L8fGGvHlxDAzupYWu7/pG6MKYCmWuf9cichuGJFxu+7aZCkzJU8NYxkuewsrCL2CredG/2d9m+
BfJZm8gDM3ph6hamRELcjXh2OBAZaH9X2nHtvJH85JFlAt+ZLl5V81ZeX90VjDfiA9t0C7evCAXT
azGzrAWziGFFYBXsbuigc8p8TKZeb9j91xjVGzjityolrmzBlEyYbIFBvI2KVJRT1SkiWo7+payp
kVh5/hnqzuyUK6w+qrPjPUOp9xfEPGcIuM028v8sNd9n6JhbkycGD8h0+Xa2iFwYjAF1g6YBFWLW
DLFN6nR6/K/TKH+3DBfn8oD08fqng8VdrAnhMAn+RvhjEhOYt+lbwyjGKl6lbQ6JMLJMMWQqThs3
Oe0xyIFzRllVvkM/Oj1pDZAWKmXJbt5+pz30kCr536kDILX3IrJ1moQZ2sLWx7YiawNCyEbq6IpF
hGk4Sy7IpBcQ+Uc9P2ZhlWykLG2YH1/blElAkQkhgPdzHLqATauyX9FG49mqIlYNzDy1pQEbiEi+
Ewc3fcNm7m3Y+GbIfkb5VjBzexRInJ24Jyr57JuCe93trWTdQyTfdhWQsQ+5T/j7dz56K8nmr2fd
Wqj4WT5VVV/M+nSr9X9i2K2WXHvRgt9PtmGeIVGJ/j7ZbobgztHqvTgqtvxM5bA59e8J3op0fZWo
xSNUE77QaCSnCbLgCZCPM30nEslb0GTVUYdQWOPRTTmJYnuxoKvnaJ7XDqPAp3x0ZkcP4aO4w1a4
yYkODXH721cJ5/B/bdbvE7VsuJil2gi6ZUsIwsAhwAyrhEZVv+sUN/qhF2boSVVRFYJ1fZFsDgw2
PJsxuOcqFUVospPq3K1ZtmDxLUr6+uURekELfP/v8VlvPoPY5QEmSjXeoqVuBu6fte/pLMI0XdPb
PqWoUxre5+HcaRWNyLc+DkDcyERBBxke5e4S794kJtwVB3rDs8RmtOYIR3NMnQh7DtB6DYWmPTnD
xzD7AsH4OoWHKkvaAQc0KnIapFZ7KhqdsgFWk5lYdlDGs3BCe4mDrouFViNZ5jO2kDCfoPPNRfHO
aMPZbKL5MWa1SehDBFMBe42fM/nd35ud0eEoWJ974CPycca2j9+RqBNi2fhII7Bykl43MtwvCPa/
5QEzodnnScjfRmMSxzlQ3DJRGSvuf/vWwmnJq0nGJQunrsopth1txxy9ENBvAnyIkWbhiDoRWhRC
Fj700NS8hhLfe7q4p7BkZUrJVsaqnmOjZhxiEaVUQp+AWKslj6cEF6dJU8kD/vxoL8Qncv6apQOM
9sszgCIUpZtngLj/RIyxAho3Cio2BggAQSnraSgD/8sIGuK6XueRlleFsKbnMTKtphqvmwzLA2zH
FFZyxfa5732x4oMF+01j3/ULbQAovUb3t79OqJWPG1ePKO8LbMw+p8+laoBwyGukhMEmmKvmWl6O
ZOJj1VgmvV3z8xEwNqfXPz/6TNWlWo76wmivwj18fYlwEdqGIMd3OhWqNNHoBqRSSo4XdMY4iX7f
6U5l4zs459Kkxz7kG9fDy7SvzYNqlNRrb8RSMJfZbqBLWYGyzI0sR12NE6sx/AeRCCLYGdcBN82C
SC7APCUlnJpGFAHHvNFkuQdFaHA0mZb336cuyAalh0ORIgpjYbnyZjYLk5mrqA9BI3HzNLBlkSna
RS0CAtPZRRRUFv/6yhQ2zJRipTAGaUZguiBIbiz6t6pSjNWN07uaV43KezXp+yZ7rOt56amtVVNY
VadmUwcKoCGCeNC++pBLHQveT3wj9oXndQuTFSeujUaCnVjbY8f3cM7363lRIfFK8MBI8OgE2bcQ
MSG+AXm6c81Ym8SgnzsgijU+0PiVHZnt3UjlJmbiIQ6EvLyCWciBSns8868fdB3ZN8FKQn7yQtEi
Rd7+6kyGZXGVaPhOr+Iexa3Goxsw2iZ7mkgHnby1Dgk1Mgww1r3fyOmUrTtToq9nF30HWAAonsZ8
WYcJ39tEC1TESam6AxbInkj+dwJCMX9bfERKElbMkXtzTZAiBX0Wze4QB/eWRjUk2MIyaGzxMk0v
138u+IwEboRJUhZ3Rf7jRpGj7aZmiFUwwheD80EXiwTB6HcA1z7HKryID3HhlQxFT8QyC36okSSH
FHyZez1pQwpn8B+BzU5WrQlW5SEM85q674xPFcL3hR6+8OhLQouNjTIzVhwz0VPsGqROMx/pN52q
sp5HQS/Hb2WNNm7mBCOAQeUUJHKE2/yQ4qJCKJe61Qmd/ohezWdkIimpOrd4b81X5gefQVsFqcb3
DU7bc95KTmZ+EyeiYMpF3iKPQaQNmgYHo4apzLBoKKzHpIZ35YM1ltGcFxYpF3ZkCEQ1rGeEcQhN
O85HHzOGblr4MJhqSgkZx0/i5GUEyKl2QEofPGyMYXb8/pPP5mPHfxx4LhfN+q6wH1NOkz2+gCJX
vgRYt9J0hkJ3dWdk2Ds5uLtvcT6DU+dPXVuL7C9nJjleR7hXqRl9NnppvVg+Lhhyl8mmqGj7Ww5K
yj9/mO6o/cLB+B82IvfkdAPlWpwvA7s7QZR/Yuxgsh4JrR6hUA8zPGiT0RfTKC9TXjq1JRtksyXx
hTqPYjwShPr2LBCeTGjNrot1D4YKTqAfE8UCz7gl4tIxwCZG03Uv8IQHUSf6oeOaPa5h5gjvecQV
QwjBcmfxfpvGjsUtGm6dEIkJePYZhANiP32k+pUb0Ky9cijoFbJ4jphOAZjcIOxfYK0LOWi7OxQs
s4LgYT3oY78CrOW+gkSDmXzIud/GFnozGw9YLX07Y2eb7DBkFwIvYyeJQcwNl+DZBMcqU2BU7TLu
FX5aynIzwBByVpbKEwS4d9XhN/kUtSDqa04PEIT9Pgr5bAv5RoPHf5mFxv2Xe3WBJb9pzdxw/fV0
3ai5kf3UQHLJqFtfHcRNvR8GmK1CTIvjUvT78gdBk8vIiMe7lwDa19c6jS1l7wbkmIeIs52MAL1T
2110U9kQL0kNTGCghs7elDGnJVrMS+ZFzO6PKr2YfKgCjYS16dMy8n4hmb0nGQS8h9ms9i9B/ItE
22ZW72Q2spOrPQVk1MDZGlcbE6GN1u2qfxF5ytEvb9CJUfv0uRBKh1NpLurZcN7Yx53eEd+GXME8
Sfqsvh9YOPsqPjFjqMzAP+NNiH2i7dhAdxBVb5GphEQSXaSfdLMRE/RyiwxSWbCNhNn6nEXR1S1K
dstZVoaTz+P4l4skv3o9axkCzgmx95xNkrlYS7a6qGKEc9kjRPiT9wtIb8R1vMk/EAf0HkLYZfhQ
wX6GdzhHLxOrjFVRQhOFlByEbxtA3GbUXxDww0fMYG5+5r8YM94oVtWhZNA+xPsqxnXjmD7X/Hxq
l6Gs+BUT4wWatY7u22y66HjbmXTIdzw/gpcsmhK7c6DJ68fIfLv4lApinUP1dJB0mQxqnshwl8ZS
A0ap0/Ff4Rorpj8IVRH5OVO57Q1JMpNmAqWFM/Vr5hrQf/oNd6jAUJc/YXVqj2KDqqrg/dsYv66c
PnF20Eop81jFcgZDx36/DhHiWl4/iALosrp+yh9kvnphxXbVk22zUN5olzGbX3ANOw/z5zYlwix5
Ci8ZqIWsRGqXWAKj4CeK5npcO1jEf42O+TAPf+aptTmsnyT2hiyYtuUUbmMq2JFPmkd0yE9Me0xp
vHs8OpwwZFbdJ0QOBsUTl5ROw1fkdY+ITj29q8kK8vf64Ks/xfLsqQ8W1QVw5NmtVJQ4LfxXXmVK
EkhMK4lHRk893qte4phQ+c6jmf7qzikqzTjRMBtvFjdt0M0vNPdujFTEa1ydYrh0jqB0F5Z0T+iY
1it6+Cz6z9Ndo6oBwlgAFnFAlZwg+/mfY93yDq2dMTpdGqWqMoenm8kmHN8WlVIYaI0mkyotDNGC
J31sZDuTTpluHPgHdn8/eA+6Q7y8XFelM8QmOt86Ad25WUWOEsNZDIJcIV1F+C1nHcer5sB2Hc1k
VLpHv7bgA8x63vb7GTZGWFhcgM+O752DagEx7222Qw/oQPhAg5JMSyqJk7lP/QhJgqyeIFvKUkVk
9PG4H9l4UV0oJqmRDwWd2Ba8YkfmvHqP+By+YcAqHYuZY2ga5iOkgqMGIQZK0LTzlELC2hzX+XUL
3fNS74hmQGyus8DCSf4nk9VVQ/FjXbVAeJZ9/pNJEFWRJOsD1eyXGTA89CKAN7bT/UdKa1R/3oq3
Jf/BpC3em0crFAjiHHMdkUyV3PcHKS2X4+MkEGazP7/oXg80d+f6EHby3Z8HTtuYJAzyyHRAP8GI
rq+lTv5cYPZhkXXPT1pw/X7cx9epxZOIeD5mQeQlZbvofnB0wx89C2b4a+ko73O/cCW7+p8A2F7z
e80qQEzTeZf438Ae3Nh3tUV9O7zRPNQFgQY7T+uE7llac2Us7YiVgoG2ayX2N5Kd34jSBw7Xn5Bi
wBkGgR1YJmOM9V7ufnh/D1EoG7KTYHee1kA5UsD4Yuc3FHjSxDZMiXPW8jlhXCXP8xgVaWn7/44y
DWZbOJ7Y8v5APu1cjCamk3lWOvlZPtssgHM+nmDN7msOjsQoZ6YZ2qQjDRLq680Zy68T2nINg9q0
e0/cfrIyRG0J1UsCw1brxIvZrFdZMoA21SFDoERSSXydyh8quU1OES+sPm85MOQLu3cDYWqa1NmB
nFIdUJzzsmR8sQ7n+hMMPbEOnN5Wl6CJUCr3mpN11hwfN1iOJTPAueFMyIX/jLv7XkF9AXMwUdkr
RsnGB/oyHa9JH6nlz0vaANKG8vsCTkHlXDw9M5Yzabala23ij70yTavJl4U4RX11pqGxLK3YgOnG
AVwAawIcswXVz5CfrddxCOi0JVZNClh4VeYCrWZcNY2zWwZ85OIF3ndQAcCUQpvraJ48KdW1HoLG
aHkATDEk6KoDITIFffXrMQHWIMBlJPPxksQxvJ0ivYtbFheM0xrO/g7cVF2tQA8J1HPrmtHA/w+X
7MPg0GmGtcWGFwTAkQODNEGh+1/+vuPilepcLIRnWWUTFsgbyV+2sYnqUp0KttCPcM9jsAuztj/F
D4/cOdOi03f72AOnpQUhuZbpXDvrhqSSM3yomuCeonbU5PTTxXxZE9saZ7Xfdj51bWWlAs8WSQeP
74Y3Br583ENYtp6nO+XOY2TmyWss7zutSWGBTX3ElUMIj/lbG1yHJ1js4c0R3xOZoLiB9nDU9vkr
NgRccwKglLZ/RmJPjNV4Ipts3CniX89SffBL7Y2F2ISrO6UMFYBQp4t1LbWPibjyrL+v9DmmX2vm
mq/7g1POj7uCH+vHEWB0FAzN/42m1ESr5Nt88dwZdyQ7RatO7BVl/yTW/IWmRDe7JX7DdeaKVbOv
VwQotTJp6xHKHc5rIooDjTZZ7LFcvPzuPd+oBWazwc+HHpJAwnGrQgAqGGmn8aOxLDf7ysZQ9rYd
6nzFewWJtam+8BROQLNfPvXtySLZBKeahYVjmaeQuBumStB0Ndnid/XRyIYwAdMsq0qKacv97EhK
HbjLNFr28O4E+YwY9+tLaAkDuslBPjjr5bOYpPkrLoDrmGpiExOmejamCn0dmFXlm7HbOvfsqbCi
KG3iT7gtIjk6Ppwt2w/UKbIQCovGXYPG4QSxSD1lKBiksdWuyoqlf14OC63fI7/9PIOlt6nUzPDo
Yj9lbxq3G8SdAVSV0AUXRqR/ywVmdrtDWYrlSyr/gd+/FqnSpn0qGA0ybLl1LzIn8vyIgeSRdwMI
zTSFODohcnJJLpmlxscEGDwv6Oo8UPc5zTphmOOTWSM8OjsCNnjy9XHsF6E2Cquu2Ezx7HmkKTcN
obE67zvu+6/jEDQXn5tA4meV3E0041BjXWcni++KKrcolnVSdTLsHOAqqUJaDzDJUZoMEqGbTFZu
L4M/muWUiHYi4OQYTZJkPTKCHNC0BwNQ7Hwgf0HrAHdvPmvVOxv002l86dsb1394JTr6imcU00Pb
BXLeHtaV0f+cRdMukMMwU3NuDTK4tJn3haAjBSDBgxLddzmgdWQHU9BlcIt7Nf1I0Pb65jRkJv/s
NnuAw3YmyJsJ+rlJCINOWzsm58Cji95GmBM0MaIsS4MKYMTAvpuzm77xn3S2Xk7CgWQT82cpYtvj
KelytE04LnEL+C36cgyfq+SpUONKe64aoC1eRKyB6M8R88NEgAhdx1zaGagkDhNu2SdDGuZkj80e
YJha64SxsWr2c09TmuaKJrwm/94H8XfVFT4HUYvvRihaqP2jD80DDNY+pdmhTJTpkvXrfcwwKeZp
dYIRXQhNH5n05Gko1j+WFe/LCQw/iJX3C7WcqlBjQuv+SWInPsWXuvBOxE3ThlFyk3QW36bP3lJn
5xUaJW8FKI3ektxM0ffvAlbGD9UUm+QW9jveALZsTra6AFNlMX087w2UMOm1LaTEDy2CcquM6aJV
MQ5dz3obpMvF1w1NFjrOItSMktc+qw7z0XMQxhmhRA7g1J+raEXXy9EZSaNAuQwcEpdk7GdzrsEC
4CEyu0rUM8yC3PJJbuTIF+cqr9PHLozwHdjtu8Uogvk02P92k8ntzSIYYCy6DN9gzxcStoJ3kvSx
P53nqGgm2yzl4D1o/fJM7T8chvabbcrvalPiKI7MRTN4tl8nBn+QUGLPZgBqTnhYvL0cN9bNASqg
7RGa/eYKshNGIPxDf5+uzGSAqb16r0Y/ReTSafJfdD6mv81WHoEWqGuobwrCXKZdUtLBIVTt19ra
pDNgkFqxl0Bk3gYKIxsCn6QuwGCi2tY6U8HKPit1wgAC006jn6yfNYivzfQ2waOaux/BSk4aU/rD
C/0ykx69Z4hEovOmO70j9ObsFY63dBnW/EvI7qHzkcqyzsKNO+4ayn937aD/dBsgIdiv+HI0Voqn
VzWGL81ZaqbArcDwpMWurTaicoIfP52YfLK3gIkmYfOXQM0WEx0P/EzqRQn6xEuQRfOBKakypKmQ
Xl0RGzAF/bdcyAtwHIOi724nzKK28oUudn72f1BLgFU60Knrwi5Le98Ooy0ZdYgJbSg1W+70In3m
82i33DP3og2lbSaYxf0Y+4IYDmoL4E49yqVLX7DIbb2fknBNQhl4H8IzSMi8nILoHYsSQzjaDZPl
BkpDdyZu5hVFNRu4ficWdqgJ0mc/0cfMLqcDaSnqTEFnKuH+j5hMyrILiZGrQXj03AaNdU4vlUGs
JqcaNBdjkgvUPeb9EvuN5VV6IoyIYxC/jAABkTy/MmGaDbE/50qmkDmDpzFzUNylr6+lAwT0b8sg
elphuHKrZneZ3Y+5tW8KI0Jun7OUHUz3HpeFQAQJXCR/qBdbcptr33EpsHIVBQGx7LU/7V+ZwiCy
/98XfwOxl9by1BGEuFlLZJAG6sFhEM1z0rjqnd6g7cvkkBq1h+SqA1tgMDjmashclpWZLhX5O1za
2jC2YXLEvlVqgl2zrZWLDVIsIn2SrjnK0d52pY0QPuPjW3E0jismLEhUVU6GICJsVqJuVtdMJkx4
KXHqKtH4NKdByj4rSiVZJNDtUr9FHB6/sqK7cZza8eefeGEuXn0S/4dLCJKsYsg2cln7Xr8XLBO2
wGBq7PNsyi/OWdxhmJd6oQUnF6WpIPP3JrxSe74ZmUnOxT/U7cWkVLdHTlEg11Muqz5fWnUSswnB
LvFyMRygSuJn63LwaNOMnkWChmIE6tCljblSTGFBW7NR34IG9wYIBNMAD9P+nDTH6II2qA4112BO
l3iwztaO4WYrpuUHugbG8T8H+LAGR8WvyH0W9KegtYDrg2ZuvP9IQSup38UXOoFc7e4WSM3W/VYJ
DqkeDT0Mif3FvEsyoEeyAE26rZpN/y+C2Y2EPCQ9YqzeSRYY0V+xJa0q90S0FDdnzqlEZ8qwFj8F
n5nV6J8QyisqQGvisG1OYMBk0bi8RBfUyziEbtT9UGzUaFgi5fpjqmSbGT+oofZMRrRhmBCh4eKH
XsK39gGEl07dtNs/ye2Dj3/B+viFLL1gAn7tOFAKaXihlKSN8SrEn+RT59e/e1C5Plnc57jB58Od
WEllTIEHgjJhpunowWAwH6EytFRAlmgCAzUIdfbUU4FtnKk4ZoGbWgU9V5NNpta11Z6N+7ume/hc
qXqhESI92+R6NMYfOGBGhMnoRbXJmTZxuqZ4XG5lMNdBOQPgcyEnamealk4sWs+7+1BGgcN7CkOZ
l2pjNG6EDQJnjH26ZnNRiI0sFdkw8ltPsHjI1jWhVWi93tK7O5srwTijQn3BCpD5I6QQyXx0Pq02
UdrZv74zZ+mnT3bZRRL2XciYVNChDIo7/ARlgQhjwr4w7zFYGW9GngRN6HDdmf8sXn0iMB0RvrPv
EcgfIQIKmNKUbl24nN35Lvwy5/isKoCHaJE4C1Y1NP1233cf7EwkXxiy+Qic77nLXHlZ5Fk7mZwL
wqycdogOmxjKbfayVeOvOk2PasghDZZ2Oi0+Y8j0zV6c++62Xa95ulvz3UV2leexNFB1jB7JwI53
Cul6cKX1MN24cyYDTpjCdWkScR6X7xzLyUz+sA524oETxog/y36oVGLACzHeSRt4JFNnbp1sLbJX
cXZQeDWlpZF2yJEr7nNwp2ZshSSDafTJwd/MQS4QlTBFCYb5J3YXDl+JI1CvhpXB8E2Hkvj0cQ1l
r8xnSmHNxSrJC8fJpPnDjM+E9ZyHkAIjJg0PGaDGF80lEA1t88Bs/+DewIJE0+C74iTiLlJhpfc4
oVewHME9j/1ITgMoxkMMgSHxlR+jJqJTVowCI9a4wBU069An6RW9z96n++eM4wUDS0cYOFGG1S75
Ec0pppK6x/KoTFzF6cXWSoiPzOLk4vMzC37rQhhlo4qPd2P4LgMIInWNK0YJjaKWDsahbszAmD5G
x5lwQ67esGCP7Ya5mdR6lNUC5PsSEXycgCzko5iJlZbEPa151LhdSesXyf+mgK9nqADTGZnlkNHn
yEIxH4PTuLsXugOZ4+i8B5WhhodkpXxzGWwo4fcvBT5W958aCnYXNZFVfZKcoG+wjpkijYiuBNbN
lv5kxhpxx7h3fmfa4/Vd69J7j+DoQCMawP4yoh2/4TDaoW0rjFaSFQmeknFea1vzLzZjlzjGeKzl
Jl+IO3j2t7xR2kAr7Jz2H4HicC8nhJHyC+PY3+T7RvCS+AhQPvFbyYrImU51XQDfdkYIT1zh8DW3
F3TII68jmtwDWEhTtRXcI1121rSihCE5apzUkXKvOa6p4CRvx8KejzZNrkQahbyfU1+ceecZQj6T
ZOKuqShdCwIwPQ+cQNAdImuIVlXzUngUdUXxrjZb7tksWHEikjdg6erI3q+VPst66E43W/rgtt6O
k3IuGM7CbOeNIT6CmvXosEmSeh1G/AklqEv8/NblCW7enKRSA+oal2lXOPdXFY04iFH20dZ32AZx
0XD+O2+2EVtRuUFwDATBWbIPiBcMSsMMnI1RLyOFDXja2ADONdj1b0xudgG3zMU8uz+1klVrA8jc
Uj4CBqU9ZTXorGwB34xmHRe0RuL9sTf5UWb7Smff6ambvbGyh+p5KvJ+C1y66c30SSNXncg0F+gY
1Pz4MAjJvD7g9YrW+P0ktcfxBnOl9EQ5XQnDfmIIvCOMp3vCmjV/2J2Glx4YlUs8AhihtbqUiZlJ
xHxcCRu1sz2yP5g9bkIjPnvB7J2S1wPa4Rzm2Xl1fB3HYgDvpeLckMsCtIise2fj+gRoN5MCxnU2
5MWelfw4xb3qYJFYw5pUJ58PA43LdN4SWV56vWQ7rejJS8HTgsLn6/dIwkufFK4NOX4TDXvOyU6g
ZZRjTw/odBT2QrRyuiJeOB+zcAh2AXVRbFrIbnQ3KB9rkoMLRKfTU57KzSJu6TZ1B6h+8FmMRsM8
Rj2naBbH91k7wVg3bmHOADPHpsQtRB4JfJVUEXPVKxpi9ZwlISC7iPvE8xmBLo6rBFIdyosT0hC3
DOghXLI5QVAYys5p9yY0OFlmxaxKTyFrzvXTpci1JeRqKWd9LSy1xvLkxhZ4yp8fFJfCr7IL1qGa
GdVArFs3XN+TqSzXtPTZljTi5jAW4WyaXBjK9MUwgZ1/OzmAKxwlGgtjZEkMTjlVUJlEWTtP8qKh
BnArFVr1EVG6afkrpCPL3PuH7tw1m78t9dcVZUzUaIj4acjUXtF9ZSuzQIn+BUwTQhFr9q0L8lZy
288iwC3EgKbZL0b99YDSz69hMF5POujJoAjPY/vm4WVWdrAO4g9EJAG3OvVGXu8qaoosw9LykU6y
NZeyvjBJLEtdAKb/7pKe5D0IqyJUBkZRF5Ff9yg5GGIVvMswB65RuOuLMt1HTmv/wPtUU1amESlk
VozH7INa0Qzm2ZpR/+dojlNS0sHS+zmHnJLPdxmuKlxTD6E/66gZ+XGVPJcZ/kec5QjLd5CxeysB
UZahrk4OQRTyQkiWUm+FAS0DM0Wx1EsW5U4wRh3H0kvIFlGpt1C8sVyNitNDDjcNq5j/DuCfx/se
LmItl39tpdQe6iudIXSaPyISrhL1zCD/TIp5llri68ufR0IGxuGWKClYFq7Acy0yptqaxJi34mU2
fOuT6b0G5novdpDUHdWofd/CLCFlBfeTLd0zeRycyG3c3XwPfsLSx2dmvAeKopkl98Ceegnu6jq+
WBBKRmFFj2AOECzulM+Yg5Vp/rAmbRDkk9hTpI/OlHcEDY0DBkT49TvD3nLkUkZrD/RYP2K2jxzu
ph/3wVMmiAgyr1l8GRD+F+4CPHuJBVBn8n5z6nYJco3g8CzI0W1PfWnZ2GbPIwCMMqGNvkYHFTpm
eVoHorB2uCjLNpdHoDq6TwsoX7PsfzQ2LKoGtGiX4rkim0S7CAVW4xKU9rddn4ZGMs4iY8re5Fyd
l50FFAXZ9cW6oURdLN1dWIsYIMHoOFWyTLy2vOkNjo3ldAoVilKqKsgQbInQKNRTG5Exs/gttE6P
wqmhd0nMPGYrmp6a7SOtYJY8Z0FUBgfwQCVxNJwGYp4ofOUaGXMWcjW6n6Hz/clkb+CcCt5GKZvr
KIzsRPLwbBkLhKIvDYEnFrJGgqBgxGQBGI01eCjuSri19jVemR2+gutbwIBCzWuXZwMfDe+6sY7f
DAj1tDuL5pPgdeVeSxYKM2wS5+qG8K8n7d+oyrhTDWMDU5vxvUbfTkeZqXnzhI7LaALoKUx7slNy
inWJv+HFoq9+NjnNfcu2SY4CJlXMEmKikckgze7HTV5wS4lBLaWjlhpBbMFSEBgq6tUxVULAQ9xE
+7A3gaoKXJk9+8tEWlqCYkGTLNd+tXiMIBlH4ND8NgyUPXfjedYkUQVPbpbjxpikrs2aiwon7wsc
pIBV3lY4DFqGE3JS1aBZE4C3lm4yYXRfVhtzixP1EueD1yRtn3vC5nj2R+AqSIUV1hzGRjrr7I4Y
0VdDsFSTfrRB3LKljp/sglfD+SsTVraqW8L9GHlvzsaNfjhGF6B1Y9FOOxC1Bk2MwWePjqPgHuvc
BhQB9AeEPNMiJZDPPYSMa/7hbo2D0XD+nVHrImWm/5t863NUq8mEq5QCLEUAS8vZ8u4Pq0bZuU0r
yM41QNro4QP8HpQtUe5H0KRr1m58o/pMi17O7FTsmqwY2R6W+LL42ndWWujQFpTvuMIJX3t4mKv4
R2wlQqMoVk4+hQo7FdphQpLSjNO+DRZJ8F7e2NKQ/JM5mUm/yNHdbeIdslW5XaLpmuGlPgSLtOLY
oTn8mn/eqLZ5HXJK1aBAvNm5KRDfARx0tvsHOkk2mRkkSmon9pYzwdDskL1+rm6llmGOdtAWeqB1
GJ5i6AaqzUvE9M+nJmMsg3NyRwxACwI/yt77m+Ot2suVHXVPzVTYOHODOeDjSFr1628EYLGct+VC
aF7s29GlXZCfpTni0Q0XbGot4FLjsXgpded0ZvzSy+Qatv9psN9T/h5G+/I3qPTISyS/DfUmqoXl
v2q6oiRyKZ3Ci606wxbe+wATWlxej6WZU5Qb3FyJgp0EELupi4D+dLxSoYF1T/9l8V6LjeiJL2GT
ot5LfPOpsdny7ELZZYPV9vnvsmIFXu049Cq7oJbi0xngXUqMInCkixUvR1KWJIsCc2O6pHhlXO8B
aqLuM85QIqmWzuta9mSTnrS2sz0/sDlYfRs56T0OByUEB3Z/GpCZTAcP/hYcFSqg0jLvPuV9A6ja
lx4wqtcxmX/KS6b33GmwwJBHPTovTM0SNTW4j8buJFfZ/5TcKVunxfmf6VQrc10qOHAtdK8zunA/
ixlvL0Z4B3DlzDefWlMaerHum6qBPvN4WVB94hfynYijrz34jAUrUVSd3sp3ZazF5wF7ozDKhthg
3DHpnFqMHos5k51WD28IBaVyKSit0Xt2g/qtypchgsj4yWagRTbHT3QP2Iu86q+D3rDvkvkSU59Q
nIvdwbUG4IZB85joqmlwLwN6EOFA1ZyJbytMgVMdroDGJjtBGBVlwHV/gbXbIH9U7fwJGhFw7Vii
kKpZBaQbYAieCEc2lr0/k8b0ffep/OrNGgXsgQFCLR3qBbR/qQDPB6GSlr1Zm8AHeyEe0T3BjF9B
TKhUtdFCBph7wRjzNFTPOMr81ON4cNsTHsf4r3LW2Zgn5Jza4ZzjoY3MlkFViFKkbHciRjueOKC8
NYZfMeJdc3/N39Pf8SakRM7XIgsVUxCuG7oEA9E97kTwo555Ohv3QFQr7LCRAOgbwd5g/OzMoar8
o61MDmXbdoUerWKO8MShnuGZqRoDH+QEtR8pu2dCwi33iCuUHaCGm6bz3HeF8G5Jq/00n/mowd+n
5BNDP+1FFZ0rajU/7oKEdByydrt7iA79I60Yh1EzPJui0sBbwXoL09u+oOb9lKv/wM8kNIKkEKyv
VKbin/yHMtpDqEdK3RG5zNAR1/TYF86/mCvfAF58Q1uhNVmObk1lsGPVR61J5MGTRtyLdgfrROPU
JDLWopuud1ahmwkLo0BWO4fI5mAF7IEZSxljGCSTUMet0zG/yEepRuTjjdaW38Yi6clmzAy5NEmE
a9RS7FKw27J6TjAnmP+DWbxMoSyrXOUe37vV0mwqRs87ocMePLxy/Ezty2N7aqrTyweNz8rUwrft
B2pRt/8o/OfG38b1EEbd+QWfKqnZNOLiWcd7ODvCKlwz7qPVCerbHWkmSFIs3J54DYiRkdJ324/j
C6wG+hAn/gy5J1MIVP+tWLUSOfUgpE/3PYvFuvH3ABvu0hy+ptH8jQfImWFdXr+NFvI0gAHL2bbp
OBURQbl7Xc4MmZCLQP67+icFsaFEYdVfT9Nm+CYyb5MgiKHtns7+zhVM08zLwZnmuxBQzWG1pqhg
PTvUtqmYCIxTntEPIY8zC8WsJ/XnFmGeIqMv0gr/dZ/4ZOfS5kJoVQwojYtkaYlKLHIOuNcLawpW
uHp+KquHhH4DrKqMeWfuv39vhLSaXlS55pGH+SDglu7n79ahecx0fnDxxU//LMtUxnoEQ/i8LeFV
g5bp6FStq2obsAPHK8UXvyhPdGf5LLRVkDr3Qzt9IeLUBNnie4SJ/3Qm55Rk/nDOvEdvcB3iDy5O
jJ0SNOIzSXG10S/Jp7suHuishEeAVRseC1zszuG8rCNGdJq20OZC0Rphs7zA4gwvriM3sG+SZVXC
UJk3PA3Am49GwAWg7QRhaEILJ376LnebF3konRoessSMXJzH0hEra88QZtTsY0R84UnYfR0XCCVE
m9KdEeBWmMpMTFL82fNG+AGXt6cMQj73xsFwhkKzsH2cI9ahCXOqRhUtpuKS1NXqxRzr/8lWyqmR
B8t6vC1CewRWM8aLZWnvqN18hp+A9A/eQ+VyZI28pmyZnYvX17uNf5LqKh3FVqJPiyCtgjrUNvf2
03Vm0pERRw3mPcYK+W6qXJaZuASQu4uFbUYfZQHNMyfNqMsYp2A9SnI9eC95UHw7h42CTBIB/Qb5
HVTAFgGnu/8O5mFrqc8ysotY2r4qurWC82PzcWk2/AEuMkelc1y2NwZzeW12c03AaFjU/qAait9h
aRojiJ442tBvxItKcqDzpkXfpJxM2kGnT8LMvkuQdsBG1eMXQh4cWFpHd/TvxpwpSW/MkZFvnUrH
Y4aejPidtQRyhNcJqIU58HngU+GUGbMrphG2VvgJOEAJuoM9mKLZZc8JngxiIEzZzE7kaWwJn8YN
Z/uywcztyq99OIuEd3iR9+Tu/Z3J7Rt/lAGbrjxsXqoNowEXvRCuIGWbfR4y1GX1LBYtl2VsUTwg
mZOuzVDU0Oo5yDSCLehea7zWZQI8Bic4YNiPuVXAhQSryqcxdvlO+J1q0NkCJ956GCOOEfYsVKqF
jJibwBFfAQWJL2PjMf/PHp42fv7rb6K3jE6voJ8o6WzWd7TpEycT57bd3QqQvCUhuV/t/N/4W/zD
qSIkFQt7hRPaZPL7X5ATbCPJ2CQAfe65+iPfEMSWXCyqoWNXN0K9Tpd2a1HQeRpQWPppC3OB9Ypq
c4hgoOzf2JBfCgONqPmDzh6iEVMJe+lXLJI6ZEg0ZGYnw4FNvnKz7MlQQNa+Umi4HjiKbDSDAl8D
2FLdB5o1fqVBjYJ2P6pgJ1kZgjgS7Z4H6pdF6w3gQPWC0FXs6qe76EtWJBnKbCj9z9/SmYbbaf3C
c50BOEmfUE7wZMSYsfdGulnF3Dj118yTdaNut7Db2lAYwkIbcA1oxcwyu3Tn9OpnNB1bSGnM5LbK
k5j/RaF4wtTo/KywlUMRQjYhJNOVc2pvt2QEKav7C5iMCHHPw2mzlds0WxPRiB+yx/ht/lQQlrt+
wCzzhvyAfv0RYhuTluEnSyub5kHw2hGlH97uMDMTh0Tij0yaRl2HWNKk/ll2OadTQxvy/b3INxcJ
ai688f4OT5JSniWBk8dV3s7NOmOb8bThb8DS05HOtWjyRNpbH1kRnG+aG/1rgkzSnQfGoATyND1E
Qc0KiFCXNZAE735kGjnh7WBYwAESh9FQ3zkP5m1hNOlTlg0h7yTIH9Nrbmcc8TlvSc6X1VFIXJw5
uwDz72MojPn/17/m2Tb0CkAgUhTxxpjRBYfEiyXjCxhbldgNmMe/rXc5V/eUY5iDrEQ5zRDJhv3O
x2JiWgk7uA2IWqFLNTnkR+F1kvPP7icB+BQelcHZ7OIvfmiH4M8GZUJbCv1jGgYnD6VyPOSInqVm
A4i6f1aT8oyUqYu0SGDgozlyso4XBJihYoizsIm45+XEQDwwtgm9Uh2hr2DJVsZJqmD6HZdwGE0x
0d/8Ui+cUSSXSHYqtoEt/nhD87+0Ia6F97hbrFFP0RSTAUaER5zy054vPWWbTw9dRBLO91UPdMGv
5wYGTjWsAtfp4pBYKhV7SbZusHSb4PmrSnRG9Ourmhk3sFSLjpfmEoAP24svaVnNQWpxISoeDF/2
YGFgVbbtF/JcBVLmDK6wQfRUpZ/cW6dP+W8cv4UOb2byF9mACMqtxlBFAUcJtWmqXtautCtkRna5
q5jUj5XnT9zO34ZXSh8nD8gc+F797M811AonTEj3iGbieCidaeD3bkvAoaucBMIoGrsClnFi7R31
3LSRw+sFISmpk2EUfTMCVD5Uw39CnQpavsrXaqf2vWtIf77Ixn6KU43lVR/d3nrgTrlrSb0/GVrn
qbA5OWuAql2cf2E5hJVmRSaZdrt/EpgiopNjsKVi0/H8kF17JqpGHKTthPP4RRdSryv8K1VJYxvB
1pUZiRchOtRMB1jVa3UgunsEJ45D0aau9NR38NvZi7aGnQsjmHHcDCdiDFfmdKb+wv6QEN86+efj
4mOtx0MuxQkAnaV8b6nilZb+zJq/v092qcg9t1F4rhm9IdrW+IAcUnc7NxZIsLjTt5WoN15hGuF2
vXe1ha3tIL48Mn3I5rkoRIkNE34WV1oMztxESfiTdalCZvTVIYF0H2xBj3hE0FExOOoDFtRxUjz3
3D9bbgkCx8h77QFsHNKZQuyoYrya21224bPpPGSmLGjfWQdM18NVLOuhaLKOTd4lv2HDQj7cG8x+
3v+YfEM884f4AtU36b/WHK0qAptCFTIQV6MtR3npbDs139DOArxT9FcbC4hLr7UXHAizucJ6UfwN
qFUFICW8f7WaazY8ZTcdgTm80nXNUMA+wtvHGt3fhsVF0K4NkraUfC6kJskM0Wpg5hmCZppq/BWv
tM1jOBz75HHwRf0yvIhcQmrzSjQTo+cv6azKjZZ2PIHnfKNOl0UnWHh6sTS/qGAmwQEnrkKGVEYU
va1veDmArogAKBdRtYlPNNTrbkZEKnZZ1eUcr0K6I9Sq8m7WUF4uTPHOpdaTZCXl1aeEGmXXgvV9
U/waXDmzUNWrjza5XRT2F0Oo2DN1iOaTnb14Ccff9kUrfG4eY0ZufDGsXLATbc0nZJAZACidy+Q7
FWTRdfCwD89OoPYeTRgZfSVrhSsqklWu4AYUsiTGc81pcJUi91RQNnxg84Et4qvLtrNwufTy9Rqe
CilBJb7lzIYluRqpkJvxUuKDeYdhA/XXF9SV7W/tJCYO5Os0t0sJK0kuL2UCfa7CZFWg2yoZWHIx
vAOBUdm50iu6JLuihY4J5g7Q9pjJ49WrRiF7RNk7NBjpkUQDV+xvSTiXP3W+8eqyRI8lc8oIdYHZ
A+62KgWzgL0VdBrfpNwYCh0wshoLU14y8Fp2Y+Nku41WBOdoCqDIYl1cmbIOISgjcm6X+B/jeDkK
EXqxoRnkbcomwN2ztoJRdzGIOpIllCR7Gqch8ZhBT7qavf9y3LB+hM/KrgXTQ74KGu4KMvwcKvR0
j1wCZ3No5dSFUeEphOIQHIRrPU4EeLldINo/aXJzT62XGQU98VCEfc6fyUcVU7huTT4/H7ufu3pQ
RVWqSpmu2zZSALzkd1beNQT29RAiq7kLFTwO/8fhR22MfYyQcCwcWz2tD+qfKXLYvmLwmGggvDXf
oCs7yhsvVJqdbkpecYJd+lWSvUbOal2uJwfjJP492JK/vXoLepyLnCsLmNrLiRsoBKbS578HWLJM
Zoi4Shmj5ShOK0L469jZ3z1oSfIeHd9Rlzi/qoU+kKH/eahvAWkWz92EUsGGmGV2cHvJO7ORnxzy
ASKdpvwQImDHckh+xx1TXvNlgGzIsFlMZ9nInat3TtqiL4BbjJfPjcJeDjtB4IDJuR5FeBl/sf4e
fU2GyZh3KwiBFaLx6N0GUFlWLJ9nd+MT9aC3vW6kRrZuXmgMdenuRSfn/dXlbFmyEmlj/Mntbuj5
t7jioqRh69e3Lm2/1ut6sG5NFBVmekIOH1CxZpF1Yu5RAgJ8PjN3QvOVGNeC2Z9DWz7hYxB5WVIx
Su/8vyLldz89wUifqlbYk1ls3mRzumzYNup7JDHRUinnsmvAehkNV5Ge2YTyEi6ZAKVKOwRRz7tf
K9IYnA+wkGkC4I5igvpmB1oADmKWBjmzVRxDzNl30rhOoZuzGX8SEKTIZbAGnTk3cBYIsgK+P7o9
/FkAPuumwlNBTh7yynXOYmf+3W7A5FqBrP1aidBX8GooqODMc8T1ggKEXNdsOC6QCIqt6WMGqaSr
JgZ46gp77oYtSnEdnqAqt+yOLeG2QtpN+7NALsxP1ks0tVPkkptL93t4TWHczy5vKEuVcb8faSUg
DSJQizgADA/BATyprqWZHGaRsHiUfFGkahXAxFbT9swXQe0+BYdCNW+rdwt5gmzpMG1TWgx4hokF
ATxzSvHzGHh4VpipDuXEbGt9IUSXzx1mBmIpeHVERWYFs2C+jSP9VxfHHCq52G32juMLwIft7R3n
4aS3mtdF0b/rGR5XAXonS9aqFePpGrNmX0vlJnua/dzYq+eZDrjZWBhWVq0QsMdxwwtlgG4a9q3o
PHXCE+oOzPpfon9RjZRK27+PmjMSK2zuKGjFAT6cJkwFTqB63Sjxt2pMtCOkGl4Lb2tg32YoIMYH
i4JXZCNPfDd30LURjvKsxll4B9Hj+dYIF1EVkM+PaZNYBwv9UlImTU5zZE8hoVaQmKCWltR+ww6/
KzbBirVku8p8/tDX2nGciv20AT9+Obg+HrrtZ+Se3FJwzDOEM/HtZ/fiySnZU33XIV/VueOvLsyp
hLNvdpnZj4EiQ55xpNi87XNd5tLP+3PhU4NW2H72uqfqObdkhK52FkQyzaruxskFX0LeIw5o3FOW
OBxtGVd3nFXd98Ivc7Vu00Q2g7wlwL0ADN84ofFPIE9IdskKpuUnngFAxQstBJcLEOoXTzGDPC/6
9mLa0bC9vWM6t80z641L3OY5pazpevaa9rL9834LBXN1/t13M5tAtMirAbPOBlH36uzjGuMADY5d
0Oi0WNdetIBLaqC8yg/6cDK6JSEIA4uyDqBsr06Nr70+1keuKgmabngCAb4DQJfwVKPIsYoGhBH4
jsBy/4YHA7lTzu9zDfp8NbN3qiee2QE28Zs+H26kQPHTpqtAPQRCV01ofdV+ZCzd48fmiZZvAgfc
aAmLfe9n63rvQffsk0gkhfn64buW5clp83dgDEyrM91dz9peqv4RjupDyTtzuVVdO7PkMDaiXioK
ggmlQ2zl8NRYxQ72CvaVjXeO4XWSyYw3LHfqi8mG+w5rfvMIV++LDT05BHo/8WZGTFOy9sZxbEDl
146LlFp/qXDloFjVnJ2zUq2KNeQKCIaeS9fnnnR8w5OLD5ualdASFMa+3SfcNb5RFWeAKl7mjuhM
nnvlFOGB1iEQe5AjBydq/b8ceFlY0d8/leDyt7DKzE/HM7LB0vN0lEfW3DjPzXS9DjRWUN78Rcm2
+a6D0iyN0Mo5StKV+zdHl/7xIA7humZdpbFX5OoCGvu4R9EJsPfXcxjC7NtUalUYdXjILc0THOrg
rPW/lPiWiSH4ZFK+FoDfpyZKbC6IamHpkWhZUEuno/1enSXcMSysNbYumxKtJ4HJWT1ge1nNBQQe
vrxtdYa2D5nTL6u5J07FLwvNiwU14wQohCIIRheSEW/bcUhhy9Hh7jTMofUbeK0fKy4Vm7mMRSAS
TmCT4OWm7Zo5xZ604Dm0mbc75bJ/xrVhIEHFFEbDwL8AfyaUzqWcG9gpe9py4xygid+4+CrISgqv
8gvSeQ+M7Li1A99VHVLG0PJzPTNt2O4fgqHfAPl6r9ZMjuUG3JoofY+axmS8ngMP7p2V45ZBGmy6
0V1OYTU2pu9tA7/VBap+VB7Hed+WEmhgIvs48ktkW6D2pGEOSEmeaysOjUYctwqTu36myZzkHIY3
lAfyMn+ULB5d2tnPb2GuTuSCYWi/g8qBGnzTXWPHHRicZCh9CSILBf/06B+bawKjYWrFAw7nX2Ff
hECWF29YfW9diE7w+aCdotmyrYaUMLZf5eRYZT6EBvBg8DcpiPIM8RJru3PoNK2aBdcBgLwpqDNy
2M/6r7YyBMZJ6z9H8yFk6Vea1OnKTzUAeMJbz13/qcuMwGJzeSPuEWwlDWMDVuM+Wy9ZafkCOmJ7
fT9bT3ieNhhsuOcsJmcNyYCsrBxhWnsd8pxO52LF2hpru8cgbjWuckVERozC3oKD4jwJ636JLr11
FKUjhncAsQTST92pAxD9oF4DAkfGcibVCo4573reKso6cxJLq15jPoQRdm/AReWfS7XcvgmLJYj3
GaARh5lh/aCbItDCzuVKy+qMXF/cVjWXdHkAmj9j/dY8C6Ii9PfbJbVRMq/56rPWwUYkKSa08ClE
ohqVcBvX/WGt2NgOojYG31cpy47RTF/DHOqKtk1pdXRPmuMgCruTCtXUws8DwX/YAnmymDCDak4e
G/ZsBZ/q23Ata/X6VrwET44YT6P2p+Vp+47U73R9hJszFiXM7zlSKhrjgiQBHApIER7xeF2PvZnY
5Uc+SsZ6Rn5VHIz03exxRhXBi4eYUj5UkeycoINuXdWpWcTU+9uRsYvDVOKK8NET5Lpwm5vHqckL
vbXlgQJqNHWjmVeEuY2PGTmuJLMgLTteIIBztRuCzdH6nbb0wO3jhPSErjBHGuPOuVJlXGmsXqc3
CtHzoXf8pUBVSpbM7p2BYhYKykNkP0uk1ebgS1erwelzjlF0f1DqscQdxA/WS5aQ5Y37dISXtlb9
vx5yE+t9wc5ZHZs79Kr/Bh+atNe5F00F9FCmXnJqg28w/lRe0UX537iRMcQq/c3XjYAQeBPQutvu
JbuccDSWef0hyhuHigDddnE5PFsltf0WG4hFASPWG1Xp67q4aT5qMs0nsytnYWdGDqH7ZPmMIP4y
NMcUgVTPZYybwj95AykS+4b0gZks8OyofxJ50YTtQrywenIkk/Raj4a3CmCFFh2OzwDqNIR846YK
QYIfBZ4qGdCU1fzKrCasal6ZyEVe99eqOzDXK7xHWFb4Dkt9T8mra99r8wy/IrKKDRayoQWbfaww
tFZr1Jx0cS1LDEN5I6dBE7rHionoPxVWPyLLlA1I3/n4fjEpvupmJd2jhK0flG0ThIAE+IVUnmZO
4praMbtlnnIo+CfQG6tX8w/RSsmhBF1jltRia+e0BDI4n6JMQNaYqYPpt8TDL7irnYnT7H9fjqaE
5VUYIWryK70ohiEFYj9u2LaVTSLRB/AHe6f/9hhf7AdWNtCEa3Ohcn64wPfv/u5VLG+GNlCoqt8a
T+FX12yChatRn8SqCOG9QYtInTmLXQY/obYZkAYZJPVBqmY2ufl3hOYmhrLFCBKNWB1DqquzcyDp
yoDz0dqReJmLQdWxoBJ/UNHM+/anD4wfdObsdplmjI4GC1bVhmWD+kyFfEG/7alsSEO5muixFmOV
MEmlWFTukM1u1OZXzuSDYBXYsirT1E/j33/jWdVUGhs3TWn47x3IPn5CtlPT6hhwZvKNH2Ti9pDM
/7daIV67AcJSsZWTXCCvD8LUuCx2NUA07JsRwaKjexgR+OS0FGIXQ+OjTC61vXr+s6hVZRJOWsnf
WzFecaofrUgk/EzSaPOg2WDAu90B3vceeDsTNPPMD6vyk5/i/WGZZMDKecQACs5ouKF6bIyvgPAE
gWCtLWpWwEx/GeED/VsE58C//hDrFHgxT4lo72q7TQvYLZVl+mdQths2xfHXgzB+81ATsDQNqcr7
dznMRjfd68t+jM0Upa53rqktgwrc2yYvYd0nOewMFsz7SOB7vZnTXq6Qn1LqQwLhPl7/hEsZ+bqY
WB2zvCMjBkAZ/33V/CRNRfoUImloNhDoOTeKc8fiZg4bwBTbC8a5HsXB+1ABROHKCBQoTWcRkHWW
ftHI3HyOXhlAJ7C4lPiIXXzEqolgvGsL4qigygshF2tsuiqf6ryJAZ/NTBWMGwH0CO8Kevifn5/A
rJOtiU2ENIsg28RSu2XVHnhK3ZlGUEXq3nKFBvyIHloPolv6QdnGfT+Sz+pcfu8EKgpkDSMJbK2N
jbzRuDo20o4leGEGHvzghV5AasUKAbmdsLSYxfZ9NwEq/x7lAcTxA6bzz3psbT3MLbUJgBlJUOQB
VWRlqKCw4nu+AJPp139wduTspWGw9mcG2TSnJv1oQB/HW5klakJIE7v2dh91n0uNq8e1MiF1aniX
QfvEBLCJUUnceJy6oVjVLXfbUt5zTVUO08zeaK3z+Jk/wX16QOVc2+ykqcuHn8uWxiQr4v9W8Exz
2zljZ9bhVvHLfk2Umt7Qq2eR24JeB4PvBqoPO9l7JLJrKJo+WHDggnQzJ5atum+o2OwwqwjgJTNX
KwcGR1/1987DVuumf55TQzHRqX/SnBtkd0e5bf0+BW5W3Rgutjmwg/tpfg1rATBxWx6H7Ovg4QVj
AQxIj2qPUQU11L294iik7rKB5/suVWkAcUDvapUTH8rEpgyqzx29GNAW7viSaeuIPbcsPXfO4Ong
2ftqpJ5DA5Hyd/72tqsQpvypyIRyyR7DM9A6PmSfrmFeRPF+VHhhZxp/rPS6nnk0HvQlp5HRG9cK
2h/mDk6mRnL2GHDaFTfyx3CYc8XI/vOlXRVQWvWyldGOptOKFzKnYbqnuIXlG/rJTJwpq5LaZ10b
i9f0qv/sqp+sObDLPbaIOM4Vn75aE5p1RWoMJGHAnQKYbJuKLkjrvLVL8fw0oO5iR98eVtAG6yg8
PG26RojLKUsXXsx4IadDjpgSebEVSRsF13Yl2DZFNxg6gnOvuC/JICCKGyVpva19kYWvOVnRQKeB
AhH426115sDDOaDY4Onj3jeklSIqvE/hiRdpL23swHjS0zWpmteHVgW8rM2nyNoaNH/Odc5paRQ1
S8QgbdXdtMJNCndcrmP9bap0Cm4ZTFaGc3j0qf2qEkeYltbgELMndW6TM9A33bsijT+Er6hNA/XZ
pZDCrlgCTSOulcDPVj9E9Soa/RXkEfkptCIRvii47QNUGZpKRQaJlzvZcmoYh89t1TapzoN6DJjU
Vbx6rrSaR6HnggOd4jCU/c5VAlfOQblsgPNmu/ITpg/tyrAki4MX/MmjtlhbCUzFbwhhNsvR/psI
RBfIARS3utNA3kzty/zpt6lxSE/ogMZHfXh33GyA4xxTopZgNf6JezGJFddnjIwBiQE5jcExiGpA
51e5BMZsNqwHoDQqZ8HDAJH4lkufGSBSrFc/kgleW3i4zvXKYu5TjesdVSNwBZkckfx96Hp6saFM
kDsEmWy3aHLOUskBO0VVkKGfT6H2CEa2MelmVhm6zy+f26KTQxK8l+15he2opGzxyz2s2Ii/LrFt
oDL/uoJwN9cqxP1EEie/koKzTbvujKngELFq5cLpYiuO9dUCzYXpOEabn183Lu4q1akG0WvYwPSk
6aHzGXP+KxamMIHxGAw+6mbrlqLKpmxGHwdgX1f54b5lJvWMV9fZE4R9o/FucK2GcHDcsC8DDNe5
JQ+eNt192EpnVV/hGXPhsL/sI12ZczyOGXqYRDneXgcdwBQXkED7KbnKkA/VC9+L33iKzhqS9O78
BdrpbSaDhKMVOn9sqhBLhwYLWxps6+1JLt2HjfzGw9kKEkySMWd1Y/uUwFHakgLlxoBrfCk/pgsA
a77gAGw1lfyPbGQC/zPWjn2lTuj6RkTgbznWtsjIHraWIF1v6VKyuPmreqdkuWuMSMRA/TLs5L1t
uwjxoFG3UM6rBP9BV/y6LEuy2EG7s88aL2A7FWA23kvdqMEMeRaW/9jHK0hQc33TJF7pZOMEI7aG
04wmmCnvkumAovBrMc82aoWRMx81FtK6UlVSFyZGpGlf8QICtDm71YS5aGkVvwfUzDvqZvzbzpWi
l2lmcT5AyOEr4tbVfMC1PBN8V6dSWooSLqgiQu0RZ7Izgixw0hoyTHZkHZKBLVAkx3xlXzVXfY6U
L5frTKPyrJZ7GCDMd4MVK3r/jq6kTKsnW3Fpelfw448Z96AxYAM6ICKz6pqyVRawyUX+GXoK6uqT
j9lmbYoUBQwU4boeu3oXPXycNx1dBlu7jUUz6lSvAs/dUeA3+I74oizco4rLsR4LnDyDeRkdvaGN
WLc3483pGRKcQr4LjVj21s2FpH9PVGhJknQXn1G9q8xwWilgxQ7G3g+KgaiIWogc8Q+ut4Dous8V
sYxGtaJ/oM1zjOgBfn9IMxUU7HnFwP8aUqgYI77dWWqveT3LteUn2dY9DtMx7gRZnW8KmwJ7VfVj
JM+BK4ZB++sF82eKkFY+MI/3tBqZNI819uLIyt1eUqlmbu+ujdRUAAOTMbIog2ifzMpTiG+5NCJN
Ph1/kRTS97xIgs08DoEshVAT1hxzUqetDz4kdtvfUguY4dl5AG0vao9BOvThAY7LO4UINPvub4Xq
UogBZvUcpR4uh+0+sn98bRY/sNppeqEF8waHdoPQaM1gnZcM6HwyO4GN48Nuk66SGFdCGHyWWbWe
zUoh1Bbz5brELEmaWd25Pgu/d5sNNaB329+Df4ISWgeSG3F9X3KeARCNl0nEYRgHvPEsPsl8YMfg
l0iy/xIfAi24egDRK+XvwSiIufhcKV/pdDxSBDpi0WsQMRWzjGkOx8UU4fWFoRj/4s/zMB8PDlJR
bbzuRmbtBXN+fdM9PxGPve4WyrIqmyctiVn913EgW9qccXjfuZE1WeRVvG26bKQpSMAOxNO+Hais
y6RCk9VoAuw7p4bnYx6TT1JVVfQuajR4fJWp0EDnaPtP8GAleU2ncSoTOtmdfQb6voIVTHGfBuFt
dMZznu6VZ62vvuelb2SB4aLqFCCPddP3wk0uGqVY/hDN19Q1+j68BTcOctACWjyXZ2FbtlPgXU3v
UCA5uaHmrYHSJyi94UWLD9HYh3LTRzBDbIp7kE9HwDFjoeBP+vyncNRbfMv3WyGpIzD6S9PtywwE
I0ANb0NyZzgx0EvpE/1ZrQe5HXUw0LU/wvBx0bS13Irj6gqdN23UtDPTi1Y7s5m9IxI03d8xevQ4
SNeI2aiEopz3H3rf6JLowKlb3NM9RJT950OuZgtIoOVmDVd5U9cWTnBAEhuGdY7v6jlJTfKN4Zrk
Uh45Vjj5F8+w/sU/UosSloBEze8i1vUyvKW3xEr6N6KXJhjGL73YUKuvzT0RO/bgTrmczJ3mbQ7p
0Jh4jWktQvRP3dbWdSAX/2dcTl5K07oNdyjZTPw2KSjXrHXoaCRUqQtB9K+/iB5iLk9fO+CKdCXL
XNiNTK4jiV52/KxQr6dQGgyfs79mRAJ2eRS2lmiGhq/CRT7mDUZPyMlI1AAochhgbliGf/ZID/g2
oLCSu5yG4+0yZ61aoNJiRsggB+1eW8nB6eFF/vbcmFlVHXX2sY5JWvC3FZzyuOgNpXmIjhG2OSqA
0m0jrm9n76n6C7TuuYULGIWaf04/135cLQzz5/g6fjoV1UNlxZoYLmfg3o7BoiX7qtTg3miwDidR
AUmc7NN5Y+CnBgcGtdZ/F4+/DWRzEZToOAoCNYbFpePGVBy/iqDRtoFfaM9/ScY9XvNcQF4naYtf
hXsw79ydFpIHTYx8fPazBzZtuuA1jeyG8qttaZj7G8dQPBpmQ/SFLYkARIojNXcwwEACUHnwSLBt
AoYxHo2Ee+Ht6MaGqTaDXlZzruLAQJjFRxoikV5uAIYDXkqxLi1TwwQ2pniXWBLe9sKQp2SL0nIz
VyTv8Tk2Gcivl3fE2GtLqBMJpGLLYkGWCE+/QNNerNk5JhQBQFLj7whP6AUt5HPi6PIa/S0YPI9Z
S/msbCbVGkq4u/xPIllfzO5/pol+dyVW7xU9XNdGWaWh80aFnJ/t9ETkEwlQI6q2FjwD3fptEXeC
K9GirWQHHy44ziv7BBEvOri7LQo051bKleCY2k7lFJexNVdpSojOGefWvgMBqEGT3mVlYCYPDfGp
PK4ULW1TPO/MiojyMnU2Ji5vmvwS/yKys2LdRNts5dcAs9m/Do1fcepS9YFOo4cRakIZ+u3wDhcx
mrGHg7n6BXDdSACfDWN3HsBA72G8r58Np3cLAUAKQj+VZmNlRdXWA8oKc72MblkAMFCrhFn4JKbH
pMZTrq1J9G4GfIPL3jLRhSLoSz10iTOvKOxyN2FvPqmsqvMrtKazZYBsDEPWs4OOSsVd6B+LQF/I
nbjefF+421n6BsnSB68FHc9NhXNgwLovPz++oLuGxc8fAPq4RJNGxxs91fkw67+oRnDq08MIFOea
vGgRfyBWhrIBwwhHRlrTs/KO6UfeUULXxm7JuHr7KeiHNX8J9+1UlATyQdCZ8PaQL05+D36oyZGH
EXbk+z8TDJeYa2YHpgizu/L8mm/YaVxoc1F9Fj+d2oYrXhut/j/SjfROsGG230U57Oexh6NJeipc
ENFKDGz4sM/Ly73HIVwB141M6ixAsVp2jO/ChXpe2n5B3mK9XdpcOvanBrb7cfebx1zfNgoxJIWg
wQBmMbkI7y8sbKQWkhcI2yg4/bRKUo+5IT9xF1rjRWKoK/zE4XrtsGco3hP7/MX/DG0Vf1TLkVhU
BBtteYIk0GaNz0thsXWstgUjx4ceROWChAYSA/46c4l+e1x3stdmw90+CEM0wqMze1uCokBSpdZD
ulvdBJDqGRNVcAnr5eD0eFiqgDGRONdxQ0JH2g8xopQNOx7VBR7UGVgbNQgvQcH2EdTWocMlLx+D
ocOmoJm2t90RYI/T91JzV+7TH71agsUEg6hk2uZEI3Re+7VZzhW4vqJlCQrf+skMBInecExT8vZL
xnC1bA5/7lYZUNwCi3CxG6juBedX4NfRMpY90jjfOsogO0/589mIGSoELj33cdqMszM9LEJGx3uz
Chbd3Vm2Ec71hE4AAa7mc2xJlbUdfGjKnhcOF4C3LcBKQjP1OnxAPCYX+ZTScUoWa11EiX8RW+Ob
P672TnoiNSdNiqCxOZyFTXHi9+cZQJmX10J+Mde0AV7oLgjWN6lqS3ljR/bj7baFrk1WkhGtwSQh
NEXtUOi9DZVkZJJCl0CS1zuiFLq96XNJIy4fVzHJ84RPZc3ABX9eQTniejOrJHtu0PR/1IyoWjZE
DTqpH8tbgWbb9vByRCG9L1T2iYwfRywgdlMrDlg3aAXz09w8Z+rP0xpvBtmWF8GfO2B/JwZi7DjJ
XZVaGCaegNDMR0P89BUhAw2I+8ZDUfUICtA7I9xe/hPHdqAhgHewwmpQ3hc/oCwGszinEFTHvb9a
4Cs+slys9u+u+TDuJVSY3I98Q6v1tNg76TzKivD60+6pGUJHhU5+SgwGq/fi+6l7hAC8cI7HKaVT
gVE3QdmAqHzcmF5uQsrV+kTjbCHpByI5MMTrkeEZ4SjVEj1w3j9YbRZEcAzrJ8yjFy1qeCtYb123
FZBN+erZKM9GrqvU35B+OTogmCFusGD0+giTxNLSQ4jep7etHoKUITiJJbWmkDzcuzE9ACL2XOvv
DPRmyaBYsGxrMg10f7CFpf37lBck9lvp1vfWxgZAjt2U+7of97T0/scfNXqXwKo03iQkAnXWt0p3
3c8cQsEf8W22gwUpzFZ2e5MxgYeb5xWcrsloxxqf5Y1zqIlrf+0pcxLtdeEQYXZLwBGYYGyc6g4w
k4S8wWs/udYLvlHgOf6LIKjdINZ/GSzAdzyPMo+l/kjp+Lop+yVYGJLyNuPTX3wXQogNvbkRJJvD
62iuq5lNP7R5XNHxWNKDyPYD+1ziepjlA90mjR+UQB1uwo4DGGP76y4vjpY8/d9WBH4hCjFo0gC1
FDmqJzq6FgD18vPb7dgZ7aGQq1aWd+dx8Z8+Pd+81cHymLTj9HmEdNoqGNG/2HA6EL+VwRSLZMXa
L/CddsSRDJ9c0c57gpAD/7kbYvFV9sfN9toUPmz16XzO6K/V9glPolPJQiaGJ3Uhf6nuGAsCexFf
mJPvI9Pzo1mhXR6jyhTKYE67a1NwhiMmZtTlMINHKaGfyPRCXauFxbXoqhblKUIWMuDs08TVdjKb
/kUcBqIIWWz6rbuRj56fzxpJ8e9HVnY+zJ6SdplO3pEpE9ATnt5VpwkZ+yWwrH7cKW+Vpt/ksIeJ
pb4Oq0pFg9jGiHTyH9rZnCfFVQqza0V5kNiKkGtQY2Md8J8YczUXdzUygQw5kzqc/nnGc0ZUz6VD
lAyO3NoapTBLKQMckLcEeipOy9vZwu069FOWhOFlcVVErYtbfIip2e2QzctBBppF5TfJiKjzqbm0
tyXez/sMXGbDQENh+l3tN4qnDI6/azyq7kfkyatP91kj1NYSGs1ZoSHRH9Y2Moij/e3yIB1+HjIk
2PaIl0/ZM1LxoZ6aPJnmiy9bNcm0ZYGpqnShitXCSJm/o1KNlT9AiStwQ6fxL7dzNMTe5VMX3AlA
qtgHA9oNjZXx2u1fma1mBJJe2gXPJ2ZAXG3kknXHJgHUHzBCsHdumx7GdxkGKGMmZ2VXYLmcIqHS
89eUemLntaY0jo8ROC4pbpyWPmGTsLtWc1wRpwHFpRHBI5Cdm59YY+cfUbz7E30jAJx6utrM9Ae0
HKiSB7Q6REkHtyGKEkrvOpHCdbs29EZcdROXtNqZPwOFA5E2obctnbit93V6Ubd6uwRnDpPzY4Cm
Hpor30RVXBgnT3wNaT0jtqOoWim+e/A3HQYULwGrzuxncgo3ZIdDAThK+EPl14tUEUJX/tAdvBIm
D0KA/rVEPe46s3t7CeQf9SHmMIu91M5XuVkgfJPi3LkT5zaX4JRkH/cZ9G9IyHz7eJZtA+jgTpS3
sTUXS2MDKxPV/tYfxFB4Y9OVOUStLOxD1wNuBbGQ5le0UnMJ9AMgQA2bWBkBDKXOtv3qILaIxAm4
iMRtmAko5xjtjxzH2id4gXrcDsiE83bScxmisx7jEcu/sVY2KzDEuBJMlcUhAHR7EnFXbXuzGl9W
wXTqCLbdko266ylNuWoKl2FCIpUZZ3DjXVPBOdvuGbjOpRKxBoe2f/G36IDSVH9C6xGbepKXh8sG
cicbCPnG2eC7ZsCiFCqGx4ti5gM2xr1TzuutiMRR7mh1qcLheXXpX0T+QjES5/nco3ywEDg5kcu9
f2d+5ZGBZIxLmajIJdQ/O2QENanSLc5jirdklMLW8hdLLIGCCQ3d1OclE/qQJ/rAp6SdVdV7Zrrf
pxbR9RdoTSme0wg4vAeJA4kD/Yidr1vu0tHEwnL25Z6SQ9XMw8QSwZbmPR3DwKyTI050i45OAouV
vnoWQZjYVOeoTXsreGXa60rncWtvr9Jk2weW00Cx/ZttA+ZG2t5WexrSJ8uGnjV9cr+Eq98QJDdj
o0RGaGAb7cH/eTulxXI85KMMmy8n9kNedxVWtrvQJKOGGP6HLrrA7SMbigr/zWYOFRUaWdxOfiIT
8kLDvjbC/K4Fi48Qd+3o+e/0uga0+KwlMtV7Mz3Y8HHhjAmAPjmsToekRCXc8SKtmBQE0KibC9+A
1a2FsHnusn482G7KKUwwINKQtIuf470EW1mTnKUpomH3wpx2Xkg2CqDqMchxjQHZJDKbgzj8hyy3
75A0+x3PiLf3gSbjvHF8nYEGmquH5lYE8x0T+RvUP6yHmGmKGj/rAvYp6U1ala0Xqtmw0ld7vcTk
q+PGPRtD4kvEq8Qix1turTC+83Rsrp/bLq7XZdMw+AkkX3OT6iaCvbu6ZpK8aCJEJhvTzt1YusK0
uk7wpZQFJM4RsUndo7BLtLnphNYYicxf3NJqnPLONWbZglwo3Q0E0nCAr5nBX9FrYPrLjJN89+gW
8huqmsede7P1FWXtiCoAAkhuGLIx+i8mmIwj49rGWTlq2P5xOMYEFTcDp2U6YZL/HMgQB8nP2Hj5
AsyEUKlWyFHEF5nV/1Cbk/FN6uOgmnZSMxw6HAmyZBWNI5xHqp0lNm4k2fAsjPSWjazGUbkdOdxv
nIxE37T8ensm9yEXXrOtvIjxpBddDzMTToqCQ4nvmcYfVKGGyLjegIEoioO9p5wjv/2U1ruBgq/D
/ubq0k2esPiUzBqoyhwDSi08CANBUoGkD0Ug4VzccYA2qApmFuiITCUSiNc470Hfxn6C8ZnFBMC7
c62aPhXZTb+a5de4uOkSK/nWb1jRfFKg8m+t2UtDEXXj4ygvl4n93A1LjAvfIEZAsdm6V9flaS++
l+GsGYG8fWMIBXxR00g2ySNjk9rLlSc1BBHjW2kQnCAb1fkwA9Ly1iHlgXesB9uZenh9rjOX/ZLH
AoDXr2rS0KinyXjnE9i9NZvZplMfcV3f8EL2bFFd6Mb/7gsEs8RDCtHyeK12Y68Qk4MQCKneN+sR
xyy+QPLa+bW734x6PV5UsF1pXzZg9H54JS1DjSZo0Y7NzuCYIq5CMBbY4xuhm+WpsR/Wvylnc2QS
Jpyr6BkmBJTbTL3ynH+XRxV3CuJwOAL1UqIObk5d/7R0qDibd0U++BpxOl0VaQKswrKjUT0GcROO
Y5V6Huex85M9aSkVODPcrN0aZEc8YCY1k/yEDVh2Sr4jiL8//h/QfmY25BuGCbhXsYSVM+SKrlV+
H/7AkCQVxkvrV0NGhtSatQ4N3nbBclv1aiEALZGT9aUMBAgYU08pyKhxLstBGTf8QwB+BwCzsrtx
88FqCQQwjIQa/HMISRr8Hbu09q1GtMDgMSQ5ZoTbLFnxasirUF89pzWxEqEM39mA+FWC630r2W7U
plWEPSHdme7pjFQUAUsqC+f9Sx/PYO4IGVIzoV5P/vMHCtrFixhLTV4zQQy8cqXyGPQRexZXEaMP
L3pdJejGrJ3/I86CUdVPUAjwzz02/rDtrom6n+GQU50BIR8inPsDA7Ia36YLIVAnBCwdRue9eGxF
gCWcE0GA2xXLUtTdcoxr31Dw3KYmgHFMQRtYXPsIAyOcX1POKNlYxroACnM7Chc8XMsKrMGAX7mv
oh6Br/YJ3hB22AdFC7fFrwjiHFx05YSWhSliy35ZexC0u8xgCoivYo7Qrc8/rZhR57RIAFWMD/aj
jLJy1Qyn5Rpb2u4E7262ETb8C46oChNzt3HCGKqUNqbM1mSm4fICfQMVN6qOqAOzUKhZDp0a9ccw
iJBaY3fnoB+GyuJ2jSYBZkeiDE9dWoZ6hmoxVgeMe2RZ9dPccQGOPANi6g2zgZFOhqp3kMMc6hnt
z3EjZK/UrkLxfYfzqH4LZI1dZIdplJtV65JKDnLr0cm3j4P8DklQxPOz8Kql16gTod3fO1rFk02w
HtD0EJqVeUdy4pM0GW5Hndvks4hPI6+e3WKm+AptPNKVntP+ozfTlqLjgvRRz4U5FeIRjn3ef82V
+zVHwlgLlNOZw6T9yLSsNDtmDvG6puvXFPNddgEuxN1M6iPBetFMzlDTYhlFFHdY08pCr4tCgMni
UuHGDBNzbFgD0RqkIe5OGRj14ZZw3k1/eN5uWkhv+/fzKRQFbn9RRcpCS4bJce8xk8b7QlNS7SFz
0cvItg4t6c1pwNFKhZmnKZG+XpI+UoNgG/fXAEzlwtmb9I/dVKPPoCrhvp9U4leP5L/tm6/6SLvj
pMwQFRZXnzMwSRNS9UcV7pGIYCiXuzgjiHeVoyJ5mQ2UWg37GJFHR2j6wrWEx7VvpmHYCCf5VMeY
bGcHOiSRMO1FUkNuiX9djTb4Fx4Jn+WWMu80UqO0W+Zns3blQhvv9oaM/qhwBd/aTbh/bphbfX3F
a/SeJDuQ4X4ow62JEMaGD9WXm/aEbW1MbY0CEu3nIjQp5yfhKskC8NEgKK5583Ip0AGRrE2kauvz
IvUSNMDSj63K+0/jQRKB1GghVhUmBMV9LAtDAbYwtZYkQigil0G1jd1meaHEIKOq/8tWRU8cuJrS
9ohsA73DG9Oow3nsQFy17Cpyntphdc7cjj8MERiRoZOnTo44ulsQtQT3K1LK6U1c0n37EOBeOq7W
HhQA3mcFgzrCJiDrMTbuomuF8Ifql1mVpzxq8tzhkkqpMMoaFDsf5Qdl6bGD0rCxdCXuJj9jqmS2
8NsdsTkey/3hyUtFYTnYJ00WU/ps10RbBjQcZsBn9eEW85cJj9QkYHcigR5VBszKyoK+ERiG3LQJ
YfwamJp6LR3Sbm2G0pqkaq8RKNeLXsSRTwx703OMH+vGJpTMx/glCg+SN+RGQzFhK57vQY88f7P7
6Tx6JF8oanBYdOa42Pan8NAtOdbSwxDiSilAv6ctLo7eyXAWoyxRpGC660HL+dqI5SSeyW7pHymX
GVK0MTEd+Wl6L/BZxUb4ZYuHBVdeIQ1jinvZtTcHnjdHA/1BQlk+4t5YXdjzyvMpRdybXWi8TnO7
pEwu1UqYO6zzyibmW0lh1BmzgRLS1eOAHujV5mtGowa1sxv4gWuXjvnXaZtvfG8Ez0I5W8WWtkiD
XMUY+pFOKxD3LaL04V9KxztXGRr7W34jh8yUydZeCmZUL4nWBghHdcGLfgLr0a22v0lRfvHgCK87
9Lb+kndwugA6lEQxoFRloOwSIGOibAB+Q5hK10s54CiRtpi1kTNlgrtMbDU2A6OERRdeAkWlO7fF
22PbXFStvJeDDS383Jy/8ltddLGPfCrwX/FE5cj4/MPIgE73WGxExcBzwPCwpiqBUw38sq/MN9kk
PaMocJYV2ImazGWVWIts7xVgoFZQAKAxJUB2396EKkylTLmjodwHUPMIO0vboFvGhuzLycv+CKyG
h6JrEMo+zZZsiWpi6Kup6Z/y2SFr7ThC4D5mGH1yzN2nw7kSpj+luXxeuLq/JNM5Hwz+/1qrTkiM
Jvcf+ALHJRJHOPKW3y86qFW5wYKZumsE/gxIeLxhwWV5jkqQNBEdavu0KxsSv09qwK+0HyR8LkH8
AMzD9K3GIwufL1uVCp4WsiMQejJvraqL8d83EgpFCTEbBcZRF9TjSGJSDkUO7OaDly2u+HLPwLoX
ntCbhBn7qikxKEMDsfsdCG1U5wySJFfWiiiCmMEUaioruZJT53UCAB258Jaqn2yMcGFAKPUlmIdY
YcpLCBUoBYADKoZlVVnou2ZsXmordwhTBKhAy4XD9a/UlPrZx1VBzYof6ngLKVFUQ3l6YCrtM/gG
N1Gh57c7Yz8Uc4ZfS19CVRO2ilfVoajILEBaUEnI1xqcJcGfxD1I3kJSVBW4W5PXHsSoakcPjc+M
U+p8g5mHRrzjgHPoAGDWxfAIDt27KfeQu0ryplL3coR/oXNeVGfpAcPM3Dk0FBFHLuPsffMuPAEh
Ng/aD9wzkyfZjVc5lWYOSCoVPMcCoISMXA/WMTSrJ0T3nGUadDqleJxDRqhcFdR1XszGtJhPLqO7
knbsQBvemn6Cj4t0up9/ydIBH7D69VRpBnqDJ9tGNBEvulD2xuLElbCzInkZ5TC0jMnfDAz9g3iH
emWyGCTGuwx9/Kx8gNNaKhJtw1SQ+kgaxCPpBPBawImqHkH8mlZN6OlXO/85UvFKfMIoUXnSy0dL
JTdUuLvpw4ZDn2UPTzyKroVjwdcVTaSOcwx/tnh8kPLtqWtANy0UGfjzdwbYxmdCqNYXqBuhyc/w
oUL/Z2SMxbk4rAgC+ibwQ8W9ohY8DM1TNeUDPaHK0681iHQ9Eb6IgyjqB0q1YT4gXnfcTiYWvmy7
upCq0x7cofjEbZ1bAwzEJpA+gGS/N47PEUcFLPmK3sq3vSv71elpdbTnDyR4vNu+PUNgpPr2/4Ql
0MGBdPtPs6yxPqYu2DEb03D/lEEYSZCRo33o99xTk6embzyOeGe4NMc8E6bwbBOOjoq3ZDHCF6Nt
dkGbX7TNzuhmY/jX745OlXnPALEbXflYUqgR2Ds0lyWbOma362Qv0xBUkI6F0EgDWcdE/0/wVi3O
9P4UN96FbyweOFprGBMr4Hu3X+lDSyY409Vf+xx4rJr2B7zjNHi3ETbwz08edAkPCa+vcwfDs4Jp
YYrz4C9Z1uPDcOhdbMMczkhSz5ZuNKGhSkXnGmmH0+QqihN7XEPgBGxyZQJfJLebheYQq0yJiCq6
g1oQPEWVDWbxxeE6KcMj9k9R9m7aqR6FdeQuEBVgfCaead0+MmEo2aK5W2xInImDFNzHH07QPswF
R1uV2T3irvPlZ3SCD/VMvm8BL2vWoNeiHGvJoG40GvS/CKKJTU5Qc20hfLNxf3kqCVmqqK9Uq2Gp
E3+e2xzzX//CZY/2BwbOZX7PmczUmBEHJ5WXjylAJEQiKJG1r1BKWnz7UxfkMNeSpHRk7mxZCS7Z
0dBicvIiFwMX+cN9tpkyIKUf/weMv9nMKDDLLZMR9/7yy9p9mSAF85KiOVfmk2F3e9PIZxnelcjO
xaUIHJ0WwT0lRRSQ0um6pv+T5WRfLZzvYHUbCnUbFG9JLT2NJmji6Y1zyaT0bCArRLWmART5db3j
PmqZkxcHkIMBS0xDo9hM+s7WKXRofLsZKOFqgWzs6bFVxHdiD18XLhjWFl9Ed8kjP5duKwi1Yjlr
jOAdVGhdfUWlU0mcZDFOJ9dtv57tf981n4q7KwWTDEjcmk9qw8qV2nVLOgIpcqO8tA8aMUSXdQTe
GvzfXo4osEB8GQA24IaQwddr01Klm9pMx/wU8qkyhTPiCNFpDRuegEXt+vp+m9wZZzsIOgwdXK8z
t+0uLktwE0knzoij72Mv8dwCkkbHrDjN2/TMVLhW7s78062CJfLjt7sxMeAN29+8YB5uFuLmfynn
SEbRIkA4WQJwDSHyjXGa4yWFFgkwCDPyG8lYEwpxeT5synIvu+JGTr+8GjwUaPD/AMz+7mBmUiHA
2t+7USAugPmx/7Ol6W3N3PHtotWJfkbJYqgOl5/qGrcA0zSzw1xnNk5CepuwjEh1pOLoKICmgxoY
CZ2z/g7ZpgVa96nrZ5RaK3Trlouotz3//P4b8uOS573Ve2X5uvsx8ePkRmgylwQaIm0/A450Kk/i
zxoplUqhRIpDpkhjEl27IbStOc32vG2ymkD8s4OMZLbABFB4oNS8NyKP8N+wmwEgCJXkp4qtj2zt
YuO7qjPX4V9i5k19kdPktViT1mSYFdrcYDRyiufuw5hldrqWdNqAdON7CiwHWnLv531grzVinXaJ
UkqLROjpcOha97QTr05nevt5N6BzUua7jzNAx+br0M1yN/O9PGShK++d9qWWJ2kvOpVTm/SMqKiV
KTatqzk7dBqMQuS8SPAUHCnCvXPKgXb1kckyE3KNbh+x1OW4P1FUBw0IRQmwjOVUm+mJFVVQDNO3
/1bT47OV84zxMhJPSQnU5pj8b6m9r1ykpY12LFKAtuV5aFeruhnOXwE9/0EN4ZH6I44N1HshYIrx
LmJNSX4HhKSOFJy0FJ0oS6ZmKnSQXK9/gNJQNOZkDb/6L4mEGRrTUo335WAO+zjDF5EoccIfw55+
Ga89u7DzQIMB2z/Hjofszww13+BtoqY3nwLomuwaXQ6Y+pr18a5Si32gowTrbKL9ZW/WI2hUoTfw
gQWarGbV1LCxO+sf/LtP/ORBxXKDAZjcN5e6eEG58xVR4IDwPGcLYks7VFfpixXVmynaCkZtKqCf
8nBp+1LFGuPlRvgxeBZEQC3rMZwnsZvPJk08+mtuze9mHEtTt+2fvQAeFaGpQs0wtkXt90Z9g5r5
4Mx/+P3fS9u+mRBVmfmyna3QLDAuLlkGE/Jjs3lm315U0lJtmxutVEx9//ccp1KY90YO9Dr9Mbbj
/PVF5HsL5AdETT2JHD/kY5bHLWcyD9ATxq0YafgCF+Ux3JMA+C/vibtUYxPlq5nRklCUa8VWF/Fz
vu2tWfUj9WQcQtOBvY0dHnolrUmfwq0OPxPPfNUXcp7vW4q557faIZnSV+ZaCKm3EoU3Zd8Cd7Jo
w15lRfRDZtam+IljYNDoGbAIEmy1zYegUpsxHhf+aZIHdVbM4PKgCtKekkE+etBoWeADfqbyOuE/
DsJkQIyBwfbuONwHPAcqHG1n/Vff/LDbq0hZgwb0amjPcIU3HO8JGWYVB1pjlebZ9VMRfH+Djap9
YGKJ+zuXAGo5DdCAkZlr6B0sK+1GKaKQ9x2kD5BciMk+3tEtz4XpZ4jA2oEP4lNXTdPct7wxihzR
CvfUXMGn/XxURT9kraal05N1zIH61dNamVLhPoewBTV8FuzFQKCXG4QrCmO5yZuwr/2AEAMKsOEi
Fuq5GbjDVGGZjxl2UGgqVesPGhxa3JWsyvUYZ+1wyyBF94E+hiNDGgueSb8MG78jJ9i/8XGXL1eR
raSctiuHGbBQXGlJLbhHokbkyFXFs8UtBAxNsw3gtuz/d3vXMjyc0YWP6t4hr81Y4E/c3UoMVlDD
JKOzv4T4DSoE53lmDRQ9W60dqaW4byHuyxDbVvQVWAPhkya6Z1K7PvWFuzE+PTQWDnJKZR81PIOY
Mq+aSEmlCLRZyb/GQEe7H31sZYLZosAWfAxtAhpSLOu6tSgK2wH2+V46kRfyiOySlsH3cEjCsmZc
Fv4a0UH/7qf49b/1+z9p6cgoLzSYaP4Du1pbcJRaXPRkXBs1E+18rmlcAysjC8yRiY15vzqZ+PJY
GwFtqKB4qVA+ZzYcEpp0hQceF2O8RPcFu9+PZ9G8giFWu2REDkkyCrJdD02YGnRsWajx+pvgdyxB
naqiYrqNF20Gl+ia5DRWba3mgqWnqgkNzWf5l0DQMezTAud/t12pKmB/4fu8pvy4q1+Qn7KKl98e
80V8+8Coer1cgDmM7aHv9ky7rFZ2L4Yb/TQPNBDBI8wPzxz8I7Ym6pKxgdv7Ahjxk0tYKIStYhwB
LgqIpO0ZYLzeZDXVWjfMG2elvYnlh+LN6243xVibt2UaLgg+27aHL5ICNaCSqHv/wtHSNneZCeCT
rH+PtiV6SubVrbuffBVw/I8KiGT9ZtidaJJIIZO03S666f6jMClYzR1+j29B96oqlCOwqkXOy0Ut
Oi4Q2rVvVPi4QmzEljbpjeqOrcLapnWVqdKew5G/ZsAC6AzNJVoWcY13LCXbaH2Dju6KjFY4Ax+h
lgfCpn8G8FV9TFvh2WCFHRGghn4TSIf/n+dkOFcsFgTXXk1GZqgdiqS9XMCGgiwV0YhvgVChqBKR
byDU7QuC2gYCgQ9M2v6nYkzrhPYzD65vVxWg59fDNV4tMQsAx023BEXP2Xinp5kFmB74jI5OuGCx
8/xGNXnUf72xx9izuiq7mRKXVK5plFLyVwuXlai/z68JEmXi0mrZmoKeVzqAIf6WPA2GKtKJgqiu
Xdz/5IxPlOvH4n0R76/xPfpAPJQK6mTo9WfFi6RfuJ+MpEjc2khXOiwdcxG1DzJHkYkaYP7hqMr0
gOeiAEJy+FIXydWyPQsysxQNlf3saXUXrYX/xKSZF2qU3OcHvsaqPEoQ1rnk9LsoC2lpskIytx3H
Xz2k2IKwf1Js1tmqtBCPrzH9VbHffXaxQ9TNmYA+yCHfzd49A4lxlcSCbYe/mvCW97yHt3rsKMTi
UxCzinWUy1xM86S0/vCXn4UIjAL3jQ0p92KmtrjjoLcB1dAx+pbm+sIqFN3oL+BFITABve9i1dUV
R77JpmMgqnQg2uaVQO8MwYcprZ+uPaZ7MwvmqCWvRun+jNgo2FoPprU694OORy+mt1jky8FWFkQl
I5jRXsut8V2l8ehuCJE5HKzNaQNB9EQljs3YvwuEcwvtoFGqXr2ttuZotY//KdexIu0xX4frRNlw
wHeihiFw+NuKCH3owtivScyXPIhv5EDA4xwibRmKopwet64JU9ADtj6KqtvDKjgNGSv0SUCUZ+Lp
N0PFXc6Uro/Jo4iY7xuz7FWrREsyGVhhPXsA/3rlCOQSjdlg8LRza+wuPFMK+tmknTJJnLfpHgx+
817DraeTLlHY1j3iZ+nqp6fh65omeMWSZ0S11CgMZsx40XcyEJDzljDSXofXpGxMjWFG8Vm1Mb/r
2W7c67iVh39Yxr2euc+9d4rjf54bnlhx/MzbIWpAQaA4a1ZFn9bprIIyJc/AwyzepU/Jq3dLZ1Cd
IrUqtxF3Rs42bHlPSEX/n23ZSeNCLOKONDIb2d8MvTBtZkU38LB0bGLRBin9bWUFni7BQBT78TjW
58NrxjMdUXRvAujDO87gO6Fe5WfkM1+4PFuVec9Yrzz7ChD19zEVwFUGBaTh1QMSRp1S4xyAhMSC
0Ggun/hmFBNNixFcsrPayPEq4KNh+a2E6d8umlJbF5RqaQncJV7fa1TIsvJD+q9M2tUk2udB7K+V
P3nG51vQkrXSuA8dHHn+GX1pQDAfQEFhmGsxRo89yEcXaSLUN08SvXkE9fIB4jfki4taoplJscCM
3iipqPt7K135EOBvkyM/6osgZh+tUs/1pCA7UbqhOtcbDCq63SmJjNmDGXaMu7/eHOiS7tX5Rukn
hvVAw2HHY6wHc2D6Q6c629cWYptGhD+xyIvJIxcJxKKLwv+U1kEr/9knkHoc5kTHH9AExxqys4lK
WywmZwDHFjXjG/KTJFISUvb9PurBODsqT2Ss2HZrjALqaZnkxsOAur9lhxrQ9h7SAHO0zjTWAHko
9HJpM2UnO+XbALde2crHMBj1ZYD0n5hpv1uubEm44spOACpaHMYAIhdWfSXXz1mmsRi2X8En9SFZ
mAmaey+O8X0+iVtH0y2SNp7FnW0fiX0HHmjeXPk/W1MZIAC0SvfV1Y2ynp0ni1BIoo2a1xT9yaj0
gHUQVHed0iSz5LrfCf2O57s+8E6c2X1LS2ig2Jm9I2TT/0eLmjdrCI99IVabX4lbGItPk4SOHN1s
79xOwI4Oj021An9ojC7DIe3ohfcFDIFk1I8jun0EYaUYt/ewVnMnwjNLKntDxd8x7YmNH+AUrLxB
BWQre6zUM7OjCoeTukfAQOkhWxLyMgP7igDPuz4u0QXQrF3FqD9eBK8sTlzTK4yeWVIQmyDs9eZq
TMv/mU+Zn7poiGAwyaMSTxIierC0ZtDCYNd+epNBkZIw8TILgPq4XJ071zLFKZV8uxvwi/Vmoa+j
mBXHk04etjru6KZBmzMDsRlXflqhwyxtnUp5JNGHg362vqDAuvmoqPNemQDrxinzEI1dUhQFEBR1
qtMA10eX32GyJ6CnN5s9KfcmuTd61Dr2e/bi0fTx1PfBJ0Ur23UuUehx/RTj4SDuWyAyJoYskMmQ
T2BFfsdFgrxqW/LHRCRu6OB17Sfrl41THMr7hkB2lkL1qiujdaD90zYf7P3R5E0OsEV6UIVW+L2I
4uZsWzUpE8GJQVDLPPYeCM1QndXnmdd7Ra486vemJWJ9WAB2+j14IHkvjDD7pcxKU+RoiFNA6Tte
zxu0lD937QYtjmEBJaym0IZoClyHGiaU68WIcydSWfazOVRd7oZ2gGZ3dT3J/TBmOqodQ5Mx3s1x
y/Wf0MKvamdhY8ZALFaGgo1Ur8YkCTBg0ybAdMzwK6gD7nzGe/YYBu/nNpLDFt1A4bFrx9/yrjzN
21rE5U5AclKUwsOrQcwJrUBebPxy8Cwk4MWR1JZL6UEVSh8kQEWZJPZb2DcykW4vkn0J8f1y9Crq
KoJTGnc3uSOHSugOvNAqQ+OiXVuPc3ExiRsEd+9QEBjA8A4lpDs4j0XLXGBAZD0cS26XvtfE7+Qz
ksGnUl91iUVvQqZdJHKAGmBUgkhHtrt7fFfcWI9dYIv79qlxnAURpcHVFBH4cONXS+ljn/FQaFK+
Oi9QCnhJdKTTQ9IxaK/InM0PzeVCt/0VW+3rrNo08+PFgZH8ipoOb01VMwFEf4Awlx+fTDXJn8eJ
4HM2WFCV2mtbNIKdS8unKkOi9+RxhPIkY3RswwZEQmh0R7goTofuvf3aTseBSP/ONF1+Tu+Dmuou
4tvMorTz1Rr6lqQf0Esj9X/K0ossXiK4Ix+hJ+fqt/kHBG4vl0gwxeg0rf8/Gj27dmXkTouWvsIZ
/c5InEGn6tDr7TJ3YzzLyVnjFeXJ3t4dS5Txf6Hv+BFBfv8nhzQqjmyIlJ6UY35eLp8n9CBqRfXZ
0wWkNtULWRxzHpNX4vVJJw/7GDGBSb1WocGvqh1H09AHP7PjRjfAaae+MoVHtDXLar23LcPle2xS
8lMyrdN763dhO9MSyaCGUA7zbttTwnnSBN00WgGgdDSq9PF1ad2cfbV8CkmdNZEhetcdrTmJ/fBz
JUxW5Mmb2HCcislkoPiBWo1U5ylHhl8ictqmRd4of5SkQUP5AmQy4mofxK80epE7lekKkwxHJsQM
tqk05LPCWV6VPQfoyq15HHMibOxMtRCCKmHlCr0c9qLJSqLxQOB1robW5wbZwVD7FMPkOXhWV9dh
H3zsP2d/AO8fw53YKkO4HN9zgXfPc62XOL/7dDuFta0R/JksaY408BN6vxFrSZJehCALukgkTw7r
EDIZcanxlXx9K7Zrb+k5yykhRtWvSOhUS8JyUlbP55RYdvELu3d5BjDwbk/rfrBHpmqWlccLtsYZ
WgXb2EPQxJDERQAjNdr3rgM7eRELHURLmTcl0y9mlXwKKISdYjHc9HtBec+qmPezq30++k2Nebwi
wduCMmXF+uaxGzsxza+6bZC7jjHhX07VqLFa/2vBFrIwQTPtdM2PcvkANxo5vsT3JmkWjw3uukPI
ta42Su2sbyyCtKNM9JWdbqpWjp/7yQSHYBPz4tA9SmlVSCSuY5ZkJu0TvXKntxuJahl1nCA2J99J
slGtgQo44ir314gfAK25P7Tx7gWCH00VmEbcUwpyqljLwUlN9HlmkBQgggNsaLUReHvbKdqPJCXy
ypqA/DC2A1VivC7QEVXsTgarggriBzAUVKDWWswELoFA38X+ATZBYyrSa9T3fa4L7jfUoOi0Jf+n
3vGvEtTPhD40jsrk0Ywhw5OWywKRVW1C+gPQybdpDdkHY25ALXCFM+aE6Om9SdrAoOeH1DDLAlxr
SuCfwBnVcEOuoCISZFxrg28dNS12McJQ/++/yMZb2iyEdZ2tzUFQbRwtFwDDrhxY2V0JUUKcvvWV
y2r6VAdVSld1h9dMlm/1UnrYPzStmBtD9limYsYsOhNb+7HmHsBZPNIjGlWQwy3ja4PLWalnn79G
WNbB1Q8IZeFg2CAOo2547+k4FSTc9wgQaZuVZ2n2Evhodg6ur/VhUQTDrJJ4oEcqNg4vBITuPRAf
08Fx2/m7Pm73doW4plwCxmKh3N9AIevSQV8KVW5kC3BUFbiJB+4v5ZflwNo1SPkEAr72BPxe6dSy
BLNSNd/GxQQivUe4E0jT8VyPe58w/7b6JYlbxHJTGr9m0h7DyPpuFQmpiz/ewzCAYLCKqrIph42Q
9pMcxe5yJNWSHrF3DHaIJn1SRuCajcdkvNzIUg9l4BTNs2Ah/4wNE0+Efp3rxUtpa+MxTcpds7A0
q7cQnVOzHwWM5XVVehhcO4itG+oF1cHYZIBlIQ8J2iRvgwUnrFbag7297VZIUm7/N639/pefnweu
OjiaIPTdoCJ91vHjJBL2Zijt8lsEpJXwikhBQOjjhUH7lS9xcwH3M6h2oZ69SNV5L7cB6ohjXiTI
sPLKegnEO4oWSzzUMibDf54Rln5oV3Jfa6ZaXV2WnXAPHMzkDAIxlreK/YbDy+sJUcL5orpdkC+d
WiP/Y2e/fAJ0zbhKMhRRHsFkV37KxVNuI0Lq/WvzkS9rC0Y39jLUu329iiQZf++hUE1Zzk97UM8w
vrPZtcJ9CniVxCozcH04SJHCj+KHcZjZZiTykyhKJDB1+t8YgvRGLXs8NBbUae1m6In+BYZfiLCy
hFY5r7FdG1IE/SULEVEGrcjwdfRblQtgzh0y42nvNN6vIyMIE6UyiPcSPoV83Xgy2dyWp2pMkiwg
xvcEp/fRXtj4ilPp3iZiWO/Gs91U92gkNadypK+iN5IQd25du4eaggjQBSAOjs2xKZgSUluef4CF
7xnBSNzU6U94ktC/tUtkAbD0Gl8c4GXfrpA5DDwE1LLDFCzZu9/1d4efucf6UCvq9Vhei2tQ6hvD
qCin7R5WPC2WWeEYsPSLh9AK2bCCaH2dNdZE0QVL2+UNWN9EUTInNwFKiePzfoSj+C3Ag/QhrhdZ
k9aqXqhpNOkNC9yK0wMiFS1SZq/iYplxGRE8CrPaHkt+jdtzw9HqAIDzJkD7gX4P+nyh/kvA/RfE
aKhmjJhyHi7K8nzSsiTDYP73lnQ+gwPPmZEjj2OeZE+yRPmGDK0WrzzmU0JaVdVzgwfhhO3z/D7M
/TdjCS40F7MuhpYQGeGE0LDVl2iU8Wwqmow3ca+VSMw38rQabKescnhJnRUYNOUGNVHR3HWZ2iCf
bQGtpcWBZer/YmqLZYCWZqMBa6nwpShlD7T2SRBWjWBE8x6yEQmU2Pcw6ApfK8qQ4DDHSrw34cfJ
yogfXinMfMjWJfYOYHUJDmKXy6dLZo2TYgBxQDeSc9SE2msLcHKjQCAeiAt2oo29AgwnELsW2Eps
BZaFTzqoJD9jVsebicS7+6zZiVZ5JnYe68vMdpYKT7MeTVnoFtppInzXoXXD2oh3CgUFzLqGcUbJ
bVZTgIYrTW47f6ED4ckywZYuHqteKiKQTsISOmJs4aF975PFnnZh0k44GHN7Z8N855JZg8rO+UEK
y8/7eco9z80tNh7EmUzdnl70Fl1xk1GkRfWI2zSsUdFshig8Gm/UvF4wqTYGYgiUPBIi+Kii7UtS
6nExkfdOW2cEp1bNFeHqNVpizSHEWcYCcBuwNTOXi0zbZDlDb04/j8vP/xT0t9tHMvLIUXkedJCf
dAjbuR5AxrSxsacu3MIsojWjYB5WOaZx91UnpxNZlIcmTtPS4zo3v7gu3U8qVz8V62orxma5apdj
FPiXQmffUDn1aMk9W6qAlXJe2sAr1Lq8ZJU1a/F5eqsRVDrcu/nyO4ik6AsQNX6An5wKCZuPbl2F
3enDsWnKTQjBAfWYG4fELmpruqyOJLyevOfVSa+8i6PocwvF4wODdbuRBY6B9Nf03rZTRcd0U0KU
a/mAEfyxTqr4JPh8+7q8LiMPG7uLRWQkBwRC5qxKzc9w9C9uJgqhVw3ABoWbO0J2H+A3u5YW8hX6
qdIMzyiDHL6mntFx5JmbrAhgin3B+7VMkn9YYWfdcOiPgpTaa8yGWqGVFs8CYrLR9GvFDSENUe1b
U7/+GCp35PwKlo7YadvMnExS4OwGoIQ/F0nmTmE45Qecs2+OMzXq45XeuCYfN+v79ysotvPTAUYI
FFTX/KLa4ugWj7wXsrDySZWMCu0xSIDEwVFXYkcwTr8hTt55ZAgGyLLyz8iFo9ri3ftpbFNqfkpX
tAu6gr40R3+e/EG7UsfW1DE3zL9p+LnlaEJ9zWqFNGNZhcUSVf6JtkOjzZLVcOgnS5D+tQ4mcauB
IpOQMDBXSyBsmmJv6IrEb41y+CHC2zeIT/+P9xICAF+OG2iDGXruWtqzbb9h5KZYbPDeect7hIIA
+gdPcTClquqBVD6lR7BttPcs12/8xysWnLx9e4LJ2RFuUbNcY8nZ1Vxl8EjC+Kk0xXLcX2J1Xye6
pckhAkErQk7pf0hkVUYeC0/24gkt0hX6ysxDiiQ0RGMEi0+yLGQfxes3WEy0lAMlLB85jg1wGahx
0pq4PhDMq/RJe50PwJ3G1tFjmeqj3NRm50mI+Uqyl3/uSh13nXtDlpbDfzctEDV3YA9T5pRwq1d0
eMDsj47Fks1We4BXofcak6tvYLSCQOjcxbwqAbGj3MadnnHrJZOm5QAXpiXqXvn6k3h18ANlcZYw
vMFduaEuVrR7qcH6cn12BTCFhBZpIDHoij3PpKS9xQYfjCdF20VaHV45s0VADt1J1yle8sE/QuQZ
Qz48BoGuKY9m379CYs4CMUKKC2alurkm6NB8WkAHI53Tz0D6b0xR/6F2FopBfP1qD6u0fxXJyJpF
3ACWCGt4XKDG7i4ZMGH75MOMLEUf5Ixq0Mpo20YG5BQW/QS0yED48cOndvAJ82G7CJDIIiCcK7Ds
NHyOksk/wPrhi8Wj4e9DBfsTi5kJrB9qr4mycodajB582s20KMglpGaDPKjn4dwdtCEDin6Etvmd
5W9hj6OM1ZDU8ssm8/0hx/kk+o4mcX8wWZjfgxVUXLQ8x0NTf/aO0P+FjvNGHPWWjB1NXYKF4pCV
OQ/ejXdpuGf1ujHCD4ENBegIPu/qmCVx6I7nG/TXNEJGOZbO8/ZSOFCl9/IxAabLyj00lwh1rYOX
l8aeMz8oa5+nn+wEe/bNTZCa37/ksc6GT/sAn2wSoZy4qMxMyHddn/Yy3aLplcRAhvttvg3dIEaW
qLn7BRQiVZ+50WuUHZNXHS7O4/kd2nFXiUZgK1spHP3BuQuwpFTvjL9RdCOlxdRrvnMZ5JdwDWbh
TnKzFDbkBoy7PHB+lciJMW3SN2JAVj7IGCzS288ctikh5Xz3kDVcHBFwOflkd0iATJpoXtZxniY4
a6w36aOKg20Z2gilZrP/H50ndJtDbN1CY7jMDHZ8hlGH80M3YEhqb2cR0vAFLnz6B2UwWg9L28eO
6STEPUBz82CtA9vlPwdCuhPsiQUGzfF5X8ADrSnXNvTZ5au3C/9iXpza70b7bWSL+dut98Zxf4hk
KDa6tVAfpu91eqs6QxFdBJCq4ShhFwMPXKEnbywrh7R6Qp0RBdFeblZTCVs5TCm84phtDcHtUsFs
fZQUnVND/O+eHH5OWEacbW24KnxiM8ZjQhshRzBlRgvp7m1hiIlo/D2dkogb6gZTRg+plAsjve2o
uFYJRxY6uQFP1yaFo3QQnuBhvsJfBNbAsaRxHbrCtQCmb2O6Go44ymeYedAG+niugN5CgAYcLhGy
9aHWuCvcOc4g/6/pVet1jikgbuR9JYwGJBBQ0/QD60l8YXAgr4IrECLet54OZmFQoi/1DTef/4uW
K25XcSn+w3L55hPERg6KPwG4IPMZOwjCYcdCMEDPu/d9iEXYSmTCYhXJiDVBIdoNN1bgLHEsvcV7
ZRwNlOLtMOLZPqwXZe0MFpXmGfnFT2gDMBw1Gs5Ls0BLEMP+G3VACIb705hae3Da4ATHVX3qdB4Y
22P8cnzGjMIl7XF67sZm92yAp9yrCN0sNzUN9oH2dZxh3AGWjc+h9eeqId+5M9grubHRsaTpSDxc
AGGNIpJeImWMpb9zaKj8qOvJBrnryDxblxS9duiLC5E6JWYYaoHLBsPUZwvhwokORjAt60sH7YFG
8Sl1CC4qnFys/sKctZJE0EKVUER0/TkBjIdTerGerz+G+p/Lq6a7BNwNucXcxXynNkcMjsaOe9ny
ff2qtmoZQPAqEGDQwq0uJv71L2AyjH0LgiZss1TX8I8Frf302pgypKa/w+K3rwl91gGY25SzJGXX
4IKESdwBI+gP21UnmV2VMUHeqZSJl/Rl4RQiKwyJo5vWCMl4r2b4nWaz999B4aBVOE2WYoUwEWlV
yEx4T12tlxpApxuNDntysnMWASQ1sBIdWdVug4ZjV4tZhcQVN2VvKBYcy7CXuLpJMx5vwvTfUIEC
8HqUTMI74k6xe48RMzVK6ZB0Qc7UJPbUYOID2ImLeC01ZZQz1UeiytxAtg+xEIZpOiyS0WLDSTpl
InzVf/dI8acAha41YtmfeI4J9YS2y2DJe+yohnHCwlq8fOWkQw+VGuNEuSgo+NXh6F4hbEt0cShG
zYR8I5fz15/YmmTeHm2gMJxnXyDdRKgS4ngFig5ftbugbSIML5i1WRxCTTZXj4R8VTZd2SM0kv6U
P6HdtbzpJn+KCOjlGJYuXowZBvBqi6BcTdfoQ3RiTJ3nsg7jw9Uf9AGNYAKS9W9I/Cg/3Mx9Qa1E
Xu5hYCzwAfrqKTzUJJjhBYAN4pnQPcwfY0CFglWx/n6adqOUwj2GlY/criHkCCTynjPh0AWvsyh0
IbMYj+RbRQfziocF0/jcbNvZ5tjzwvmMZkG+N8TeasqLXUExvWU3yJ4nHgoRQUdah5vQ2c/NSubb
QqonAlw7eJ0pWfPF7zVHlFIRyjqnrvSD/tPsxA0eH+sl+0Pe42qeolO0zbuswNFqa4U5nP22L7qK
SU6P+/2BEZ9OC9BQ5NHmmqeVXb+67K6V/nxydbQ0fHnx//H1UdLCz+zD2ar3FAhJOKfjN0JKzJXO
NH0gl/AlGhXZrohOi2thEmhoWnvWdtZ6mdfDgxj8T+WLzHVTEXFyDp8KKNxHI0zrIlU89XQTItij
ecTNF+6+QBMq7bdaLtaywH1EL3R5w2MbFSDbUhMzZpiSrL37WoOne8enAxL8znw0pvCSyU45v9++
Sn+jFw3I8+iBDBhQZ01ZshBo8MqBlbtgM+DxukZWgO0Ibj9XxspWeC+xHVqA/7Nq68dbLjnveqRl
jojhD+F+hUpqNoEN778PGrxud+lhBVVizbMAnKLT65zVSo10EPKA7+mwvYL1scm6PORy+fjc3BNN
OfmHCaRHqT+VtaDMHe8ulF1eZAEOAw30nxbQE4CpHV0L6mj780kqYjlgPdHkE0dTv5qXuenp2SBy
DXTLcquNw8hqe6oZ8qTqrx8pvwdWNRUKEilDN9Rxm9RP/dSd266j6aZouBMD21cM+T7xvmhojDzR
AZvCQ90y7blOO6ZkXwcpK5wrCXTXxlIZmcJ9REB97PWQRquliSGgVEicJbu2jM4pAWiAv5qBoM2a
OmyePdX8gUINGaqY3gK/yauz5CXBxS9wj54GbKmq286bslC/2wz7ZQZphIw4SjiMKd2UmZtPBgd4
Hgy7yJCk+6hatNlZV6RAPJo1d5KioCAJ8ATcZJVmxBlvq2pwFNsMx/DxIMf6UtI3xd4ac2eSvPv7
fJnth486v2Gnu5a0EADgXVCVYZaBeEe1wV72S0mSH7056p0lZMVtYeBupypYOHL4bFddjIu+TZoI
6H2LGh96kqOUsz6WzlC7Yi8p4o/94mmNLeGAUIsYUYEcXtwMAidghLqdH0z0kNSbCmTAbe6t6Arv
zgeCiuBuscj0CuD404oDkI2zhHH65oAThxrOUUS2SpwoMj4dhrRWpYDc6pxEnJsfm8ZbdrqzgPor
96CXzpQEuLw7P3PAnGgi+vvj1qeea2FOVoGdJjfjnfz6LAp1pP1CUSUH5pp2oClNFl9bJpsGCsaF
G/PnciJpoGzuI9jbGmQAmlsZYYUelvd3aPjvC4tucl7m9lDllWp68gveIHgtZeJmHwBD/MnFlFjU
mIWss6ffk61RdL74nCMalmOvCGRzM85YqMTCkAA3t/lUA78Ec5uOrIPh+W5fq7zLZyFGzZ2Wt/+9
pVH9X/2GfZzw/8FCYQ2ydH/VoB40HthhSPKGJtYmLqf2qaKSQE6XRJRYk2KDmhXmUi0wFPoy/cx+
MYCrL0oYfUpaPDUVarNiU2mdRgNg8saFzpf9JgCXrJOTJ/hX36aKD/UX2cGE5DNo13XMBNO+SPfp
Z5HEK4CuTTsrRV6TGcGT0gJHAUbXUwZi6od82y6ChQ7l4wwpf4Aa3tQY3BooxgAYp6Wb0NO2cEmP
2whKLF9cb0vf8UoRH1cs3nue7c6/+3ToRL2FpIroYQl4BKULB/GnegK8zUxDFw/MuRoFjzKg9zec
fb3PFL/CJ5zwfMZWSIGLNA/L8r+OKOfYwY4ZtLAnm60/6zbY2TbPcyZXzO4O0EyEUrmR9XBRJMGD
xq0fAHCRXoJ8USpCKq94XBCz9B6yFnj10ho65mZD3ICFqqp/78NtJL12dADEU4sr9PLJ9Zo/NiVZ
oHpF2eoseUN3McDU4+JoDzs5PyiFfJXvEEoo3ewP1aipsyssFLGa6denICcIyykX/SCbk7Le9Tlu
Q2OPki9+1p1OxrCkl/ZC08Jm0yrFuHZZxwkb0jNHQvcHUMwgIHAEHoX7z0wj0YCB7SfldPGdYwPj
gZXxtPZnUof5ZAUgHmNGFyM0/vwVrD4shLC2AtmlgiAdZ5Tm42KJW3N9rMf88UNjdzJqXEEWttf+
dSz0oMlSUB7moKdLOvJH3l3yaXtBc8uaM//VtPYPzMHxR5TxY2BgXVnpSOP5j2eR3UIcgfMjyWGi
1IsLoZaf0OMjvYfcZABgXbg9aAeTxR9VGomdMbRKN1iriLMoInUs0A222h+zaXh8uFnbYN3/fbc3
7MrgNxpj5eRjRcF3Iw2+LE8lZY603lHswTltfjBeI803u8gK99qpWUcEgF5Vgo+TnjMjlc6yh7cM
S3xGWzVbtlb7jEmdsKIybHD4triIQIs0kMTqnFAP3g7+zhvOP7IDYKSUGHnKOajVNw5wXpvsHgjk
PK1rkKXQslkrdQDMLKb0DVP6fn00Uqgr6BBng+/cCPBy39LV6JNJ8A2e1oA0zDQj9Z+O6EQ6Q7rg
YUbvj1aua1gM2Lylmu/LpqyBXSn8GsRiuGNgFlbzZnjj6B1Nxnyuar12HZmZykGnPDKFp4H2AB15
iSQsP4oTdLIOsfWO1LYC/tN63GHSMS+K0ewv7/oDtEee/lxpeU2y730tlgTj/bzklA50EPVyADKW
jheOgUoLd3qf45ImuxA3see4m3ya2yn6o0JiCp0UMsauscDyqAigIKGG+TrF4ckyzDvmUHyuFvL1
zhxTlchM4ByLRWF2KJByzs4B7u4cS5GCfluPKTTdOX78bTpl8LSkw9KxeU2VP48MW+Nr4NEbHK7v
NhpHlRbCLRgCQ/DsPxOAYcuFnohpGUNafv5+vh4s/H1gJ4/rpo1ZaYIfgSMfLjsc91fu0TdSffbP
w7z+WXqzyhphlCTc+cfEuqnOpE+m0FreFjFJ4Alz/m0bVgjY/dIC2BpFEL1nyGKcbXZ8ABX0D8mS
d78bLL1O7ngyvaIsm2mSzWz3Af62J/5/EV0j02F2U4jcZST0mhlCKxkQCL8PistDfceZJ4sdcAqA
FEsCeCTSru7OI9zcxrkZrn/td0tmYzcXb/t+vE9FEHazSVo3Uk/Q80S67ceLzUFB9nt8HUHB/9jF
aSxTDjTzmlNEjEsGNwJ2XNH0djeO6s+xdR030lnaOrbKF+LGx6G+eO0UXFRRyM7xbqg85DpvR00L
E5iSjW6+dfElizklyfk63d7tuzuIMhse3bHkNjPpQCOT2X2wVc5k65sVgViez/NTFKYofUb6vhR7
E647wMzuu1buInLN0t88aiJvH+zLTZhs8rDauTx1j1VHdfye7eXKhLJ6sC3+7GP9/BjbAepsYjZa
YPNY2KVPv97RFAEDIvE35oY1rYAHk0CDaoqYsGIqLaMIFPGV/COLOxhXrFJSoDp9QCbvj2s7LLPH
lff3QwrKKz9v7aLg9hCJsC7EPC+FN7IdXuLC30YxlOH9f8U0uZnELEUUBgZXGtiMEVvKRDBkEvD0
ckVrumiBF3pCKE8lSpLXsR/hglKAhN8Zttm8xG7GmL6M5RqYVHyX/BgeEeNSboW89Cm6nFyuGTbT
iqEID1Yb4ZXuie7OrBYjWt/HH8nbFcV5Y3YmoLuZqlumhDjsyw+YqE15rsTiGso4F2APdK0R7Ghn
tOEmHrFTejp4+AiDQtaebX3r6Wdp1vHIrdQUT7r6s+5esOpt/NHQPhmDtFGm6TEggfN+lBIKOgmE
QL9zFeSVh+DkthwITCxcjUOx99B2Tei8DJTYvLN8fwTXwKXG8iafav7FgYZI80hI6Us/fLpJGtnm
2Hc4LXKLvGkpS6iIk1r8xGo8HV2ko+gYgbYpknKmh1fk2MqsO8aciGBxeLZ9GW68ssqPtl4nz8xD
knkrSrjbhH1HsL/jDECO5C/im0sEwMQvraZQlsEhXS5qW9N+KsVlUwVMq690YmE/wgy3oJ+RQ6mL
wJqpM5Rxiv25rzQ44ZbjC4nBR3bI7k/AI4oxzQ/gdETEcDOVKEkQWbc51OIzKziu9BJLsO6RFFUP
Ez1lB5Rw5I4mGWjJI0QUigzxaaqUUZbfQH4ZdrSITWp+XhkLOjN3Y0kyveTAIcyzO/9GUh8+gPM3
KKJ052jEZUsYGmX8eTxKDYKuRbgPWcbZ/FwKpIeGpfFHaDOLyagEi3mQgWlN2yagfW9bYEhd8XHG
4YR7uCoYtXdADRuEDYp3MdGKJSGCfA3MbZzEyw4ra48ubM/UboZU5pqLt7t8kiaNahpyxubevhgM
AMapuhDkesQ5fGGCyOiONpDA9r5IyREC4G8FPFEGeLypqcICP7RG9awvucTNbo0MBIdlWyhgVARg
HkUQE+YVxl6tV8lvIIXSVdEIVL7kAerpzZpD/MaCqxkm4u/ewWhoN3gJFMD3Kx3ag0AGQ46ZS5JD
jbvfMUtcARSC73FpeVsar6Az8YoNf8gLLaC+KeS9fdv7FkaniIzElMiCkYADHHpXz6vbkiaPwyuq
iREqg1qCnhygIzAKPFb5RCfVBqKwI1FGV9S7+7SJE1JjsObvcrY3umSkW0c5LPN1NAJidtGkJrl2
40gg/noOW5qWuJGOrd+oPqOswvMCLtj1AOCJB9UhOm7Pb917uga53rQ0FgaQVI4OaFiCzR35BGjp
dxYF1tf13uOfDGYY4Bj/hC8O+spyeU8Jh8vl0SUdA62+9AyI86Tu+hc4z598C0hTcDixewS/rOzc
6d7mqeByI5fV2Pr6oc4GwH6/4Y+FwoqpsaFdu5uCHgnl5yBH1PRaRd/Y0RLz3cQ1RIchMLRuh76f
vvNAapOvM2+If5UYGyJTsVc1vMatbY9pVBRclILcZ3sC0F7XKQ6NSB0Fydt/dz5wi2c+I8bRhVQ3
pft8fSHhcUmUnzYN9v01RVPcw4PnUK2OZ6N2t7BircVElBXyYUS2d127ixvP2cNBg4gaCAi39mBa
HOkyM2JOzBUhT0QPYS88V6stJ4OCXbKK04YZxTAnUiv9fmEVMRwsMbiBWpTnZDhJ1qhOIVTPBp+S
98QPHr8pdSo0F5kI73mUHXY7SrN62mkc16hhlTw+N9YfACt+k09OMlhLiTi98vAS6okMWENF0d/5
iLeTBoXRw/BhgTd7T0vV8VkI4WCUfV6huPNX//5fQ0id9p+3dvHSI5hituuqVs1n8UHwtVnNsTLb
9pM6rOXEw4pqxy/KEiWSBk9I3Yj1fwb0835IKZautPXxkQZ+jMddwj3MCCRSm2J0ki/xEGKhG4JJ
4OgB+/CZWhYkWvXOpyNuZ7mHPberyz3i82aIdzh1mHNrWpFCkcbBYpEcuex7ba3gWTPlqdQ6IUdT
nA1tx8U08AnZ2txHsZWM/zUdGe1zUxHVATzb2n3nFb//Gyjde2UA6oUfiJL9KPqi7KGu4+Jp3bs8
dvCiT7e4BkIqPQyBy3okMDGDuoDQuN45U0n/qY0YnmQVM6cyYkqJ4z+j6C/EvGmpX1FIXH0dFn6Q
Bwf1RQGfmC9qoLGFm4qkaCnL0iGg07pPBO9s0GbIYm3tRiIplwZvaYeFHVctFw3pwtwZwuN/6mBw
HHiPvhaQNA1rkEzu3WFBrwpUaDxxJAEt/JlQvbWMoTaSuBtmDJ/yDSw5SyCX5koAH8B0ywf8tN0D
MuQ27BFG1YpCxHAcjX1xTrcMfM47e4IcFbeS9Z/gLNQJQkjeBuXycbLUU0tN3bFWGuFKwgcy47oa
i1/7zVBgRfystI4nrPFuFlFljhnsVYqUEH24fdykMkAMpSE9PdWD/BqWNjKLhgGuGdteu1QoHYDv
xNTlHMNvmnLrY2Rc0G/+EDkvTnNM9MrDUWRAEwuzQh+4dXbVJOwjiIE9TcVdMIBgHkbMw0WzEnIG
i0nSEJO7kOn0oZHzUDwCHPv1VE2+q8FNIH2RaszgOlThzngOJAfFGmMdVH3xuUIRxPdfuAJb34qW
tgB0visDUEIplEM4zWisumwxBjchR8C0P4xz9tLQLX0uYn4Z124xQWxKHV3a38KC7uMv8MEgBKNk
K211WwvKw9f/z8c9emk7dI5uaRZpvxT2mBSkoMazYBKLnTg0b22JiNPqZMrxSKpuoyfPecO3EKe9
4BbJQTIwYoIa9m2jUJdHKRiZzE4HH88qhLVFoHTF3RuaSgmAEwW6Xbb+EtvClvjGsWdrXxwvCAEd
s07iqtLFTqkmMEeEzv8X5Kq1wZeu5tkC+TaGtBw7qw4YVt7W8Qcxg/+NPMildNX/VgUcMIVyNhJ6
irRNRA9gR7ZUM0Y+CPakuowm2fP0nWF2MFhd6yDZuaf8XFUsEbEJw5AntwhlJpg6TRm4VfpCEHWK
R3Ki00/YsSK6gnnF88Pc7LIREyJkdxSFc9WGgfNAlzXZTkRIjHJzJnA8WaOTibJ/2KLGqxQORd9i
Dk1bY3lyDg2SMPorluofST3LWRKcsULvanNMnZP+dI8feKpJDxW2GilJM5nGGwbfRM6UCIQ2YezZ
CGwpnXyXil74qm9OTI9yfEARsNW9ugsRdzhJ/TG+Tf93x5LJPJI5CTJQLGC3hYnvri3v1DYQMPTr
Oq1A4/Rc2PUAsyrna8k9F47DpECfGZCo+dCQdLjPWjmKTg0KKr7LzQ9b0n18TxjiQKd5QxA4eE3/
QuZmrBjKPYwdKEPDbwJCUfWRF1Hrc6Q1eanAPS0Z8N7ri4xb/5LT5i8SiY9mOLPU069oJs/G2iN7
4F06yTIRxA1uSR2jQlXZ7lU/cKXjnM5JpbuA3J0Lyg1iaaTQjWdeqnnUVM5XO4Taj6Vv6jSkfZVT
sHOxW2W+OMl4EKJM2j09AK59pMabkU6dXpbqSWfljRAklf09g+krj3O65fRyF4ladN2DnwODD7I7
y3AKmZk5RImlWVnRU9LUVn8LlOm93kWJoAxA6MDVyFuJrDUWePOosmHBev0uURA6cZRdtn9SbiXK
Z9rt5xi3+wvk8LXmVAmVDymAr3D1x2KP6Jsv/0cSGcPqOZHCpGMY1k50F2pGD7ZnylyKAkAu5I/+
CpgG5u62LVaSiEVOE56Ih0GM9EtgFP5sm3lSxQ7BviNc/QGboN/pYWQreht/ldB872KqmoPRADYD
4M20bgWMtrWADNBMcm4CPytzjbCus2hubEWKi2UQ9PaHQhqYWZFxGhG63pocdXVmQ/CUlyMv67AL
lopfz5/tZMiRErXmAhP3Adp/nHIDX6HLpJWqC3ciV773CJLp+2/E+0jyokN2kap1VnjKwPSEMjdu
0MuDu9V7xVgmHzUW0G+fGUWVdKRO/4hEaySVG2YVWUH5ge9odLMOLKc2Q6mRP3BtTP6UMHsktH4A
onEFT10gxTjJic62ODMtgGCV3mCRQKldD89rvW65grmy8t3eOFYLXcHFj1RqtcqxQ+HSNKwkeGKJ
T+insJ9GeIDrREdh6AfK7P+c8220hYIjZX6WyhfXmJpuug3uMjW3UACPl6aEbXYC/fHjjUDMEPAE
dnyDZ32WwJorp3qHRwlRuPFDjLYd/gB7CgeLCqFhTtwk6OKzOCD+FPH2Ofy+DcLchtWPGd2oQv6b
gRS8xxiyN+SFIQGade7+b/+w6YglPgAWTvCxzNqImbW61A71GCe+NCfer0gNe+a3q1CXQWeNdJYO
tKjvYoFADRbd8cSSiLQWpK8mfGPdFKPwM8oPhw/pibjwZOOs+TDcgkqD0ca8Gxi4eF2BbuCtHmnq
FDBeXBmsZdSh6X0EKOxMQi/LLn7LdifiBoFp8t8JBmN9Tf2OsewnXT0/Ud6qD1qHn94jB4X9Jtei
SbB8uTQ21v/T1Nr2+xZ2X4rujKZRafQqayGgbk7Cd+59ylUBziv5f9ESyOuD+VisejQNpvuU3gG7
kGyr6huMizfInqLwhUOCUixnkJ8WxfU0ds8cLuo7cewNNcz6fXsBLVgGqGusTNCbwE2GJ+kqxDhS
xv3Wg8zeZGHxVkX3Zs4sS51RCE+ObH08yggcud/EuL+aAmWCVR57N5T4bUG78WF/sX2oovkOXxlj
N9hQ524UgmK1Q9NePqy8zZGSPH8wgm08w918C9Fx8T3YtuXdiOS8ge2Fkcvz+hwwjm7T6m5U5ktJ
Fpy+K/CDkeH7nOObc9ra7dqT3SjlTcRexlaLFk3tXM128fg7opHV3W+JPYbCfgsNQLjUd9P3kHJw
WHNaQlbeJtQySV7GWfL2JxBSLAEQZasiyKNA7FrZHouZk2ImUcxseXBT2hCxrmjlPMyR7DaSlHgk
q8EGyXb8fyXwStELFVXEQYjapNtqiUPqNsmXtupouzqfttKunzbjNYTIJ0AKTnI8KAx73M4HGDv6
7dLIdQkIHBhKNgX1Yp4LELAebJ2ZiuWJUbbYDBr5UBUSLD1myh2KBzZchi9WosK2+IPdXlLQ2Dw6
DAGqfk3hsaWGhNPt0kiZskiL+CZemXRv9yDlKcRegLk4b2LuiN6f3fCkL3qPb7hgnlcB9hJZx7vF
uCQfIYfgLeOjUPsZCKuRGFx1OMopYSnPbUkJRiqW1LzjDdYQhqhXd/GICEFXreFDY9Voysrmrjzz
ofGnc/zFUw5LQBZ+XiMARgDNx5hmPqBKwS9celfncTp267IDooLnnlJeswtzY9Y0KbLYehzWbnut
bJYuzMW36puddsLkbYA6I8aoHJow+DQH9XvnoCNXbZHou0VO5qaC0LYMdiemU+u/rPPQli/njFPE
m+mMsxG9pz7nEiPWut0dR5qmsaPuFabcJYe9XFZdCycxKVpBSPYksbnZOrNPpLLa1VoyeiSRztn6
cJWgzb+gNJFlnCNbaA+HvrbLuOaJE51wDArrrHFe6Cem4etJBFUQ01Vhgyf04sqHK+hM5ERmUNj2
rv6Ux5NneFqbUha7+2FfkAOaKlCN3v4f0a3IOsz6IuYEyhZahN59yksyjtRRDAFUK39i1tK/M/TZ
e7KzvdP7hiHkKVbs8sbaB2pPdKBDGF0owDJ8Dx2AJrEtCUGgCWygBikcJzjFWzQc0EYtURpfzc2q
oZ+OO7Ujpl0lrV7iidXb550TIdYrWvfxp6mHi77FlvBXCtmO+rOZlPOZLvDl+fekpyqAOpwLBTDr
jvowdScwNhXofByTq4x2zIZtC3ho6QHX8mmv3XcKfnW7UuhJpgOWQ6DKsibCe1+fQRdB6Ykg2/zj
XGGZRIULZXUUABRHaAAFmVWKK26ZZMUFBcMfxLejBFPYcBux7JCMruDE2MMo2jtSlTSJFS1hv5/5
juFo9//7Y1/Oah/KO7Zchx42HWfxs2YoC6CtTeET8UPD1NW4OsIcg/5NfbRTD4JPL/N43N+YhioF
2MyEjwApgJzJOg61m7ngP0LadK35t596PRgbX35HfZlc+IxSdICCoVtkVA1wjSGv7lIV7SiB8+O2
pXynA5yjAz2nbINda0E0cnLc+8kbIz2es7K68LGOlNLpazsdlDV4KQIXPtRVow/CN0bXwlIWM3LH
fk07rZNY+USQMVCULNyUujAhwQL/XPG5T3Ri+t8KLmIksKjS4/Havme+qsAETb6p1CysGOlRWA6Z
E0rclpnK54PmkDwLng7kEXK3h9mxSBs0ZPCTuUKdfgT5SHsCAy+rr0fQhXo5oCrQn6aK89itV/G5
iGvBqy59RQ5vDqGu2t54JOpbyz5cFDmkyNH4YLt4fCoCNF22AOvEc9Jzdy6b/Dk01T/RSAtJXrIx
BNCo/w9yW9pTqn+xSKzjJAvwCsHPD3c1ViFcTB3vM9OA3Saq19kCbF8EYBpQHFZ+fMQnIc2gIhg/
xQURCpoyym2sE79zh6yqGMiTk0mhNPRb69VsIuYJ3rBPi1KcsUKNRAQWrxiJuSwRM9qVm3umgYfS
/a9EfaWHfwpsnSgr2q+jR6xsMcYim2Q4JM+rvHOYzGGiF12X9ZnpH/S23End2MGM+mjt/wLWjdi/
Gxsf4kse8V245QW+w4sRcDU8W2nCQAnhditdXdegEuEbGhcSF8B8gqlZQl210iBNjX5djpWABcWV
xEwTfGcwsQCaaFjZplrsVIvUj0TzuZrn3R70LwhhJqddSHkKWrkVkhfhJmUphBVPW6Q94oykeWqB
zLXBzxIgnev0AN0vcmP9FVwIg5DdSsvr5tRStIyhsvabT2A2lm0m1ZxETANLzHGrvFkQFPMoFYzx
tXDwrAHCecWZF1HBtmINmvDDDEJVT8ANtgFnDy5JFYvafa7legCxYMfYhm/WB2CtEhlVz5M4Ld1P
bgUzbRK/tvW3i9xbH9zirad8TIjOfIFCabT+WgOiqFp6Xs7TnRzfIEZK4r+sKN8dSZbfXg7zDM/e
cPhh+PPtC1TACHVORT43OOFVQ3XiZBu7xJBnGd15nDOg6LOmC3n0+nGzIBi3f+D0n3sdtmP/26cl
Q6y5a/gKjvpXcOqxbW4Hz4kPHdaA9Cjekm94GcDTE/J3+My4mlYhnAr1QC1aPxLB0TooSGcdVfu+
6oP+vtsHQ8T7ARrqYIJdFiAztJL1XCJcvcZWkAZhm89MaHKpOtMSp06phN1+NV7E+bA4XA1E3Jzn
GmF56D5YiGMULq4Qd+Wz6jkXnAVWOv/l/Ja9e0Lr2srPpb9s8rep+ZlngUCKwjzSYs9qKK26mjxd
F7nqZ74EtAXVNBVH0Q6FY/TL7Dg5ccasLixg+npnjefUuTdD5HY4e5/gR5/lZsfJtgc0NQqiya5V
rKdDOzv/VV67KccTjvOIfpwFAjROhbSlCl2A6evkfEc11HyCh9Be48drmpONcxXqSMSszJPaTs9m
5VYXeCNB80ZqNF4emLl85eoGmXZnCzAq70AQ1kHm6nKPu8RYwT2uHoCa13L9P0R5VySHqNwL0X5b
FFeTqaw5tMCiWJWqkMaZLtKNnI9NaQcVzeIgcRaZ2ls7AHeiD+GbrQEAdh3wOd+ugnP21gsVnoLN
YvX9aGooQCZIXRHmhgLpoiUFqqk6yG+YNkpSu1JcvAHwkpwrFVcSJ6D5Dik61gYbqzKGLhoIO9He
9zZPjDKp2TGQCgGdoG7w5DA1uNb1ufgNP9WgO7jTSEmDnM/+0c3s1ST7i42yRKXE6YWy3kKsw1S+
YyJDJ3ujzNIXuv3N5ID4ftDYBFz6LVxeB3uf4RyIUF6srBBYvYuuRXCdOuUmOkFQ5N/vkfWfuhL1
n/IniA3In5q1LaMzGnRV/wQ1cFF2G/GfkhK4gnYPRKcLYLk/s779MqDxy8laL4GePjdaTBwbHAgg
SLLaiVqI+cGLerTp3gEaRurHiQ4kDVkvomwYYaMO5qoMHS6LsTggU+QL5QKEhd301yzgkrfr7Hd/
lMR1/+xyk6kIp9TdizqIQ230DU7kU31wn+Iix+ry2kLlFzNhE2t4VXvY30hIzHofWJCdlvtrrY4P
rPmLmDUjkbISg8sUvWID4rtosrukAPhmLiTaBPBZ6EUk/gvXXQDpq8oCs8DNFfV+ksHnxOQYZX+E
oovN5gpzWcRBFGr1AzBAGvq+/5B5vlSGvIMjzqnZnK/7crFayhoht+jBOLX/1FOpTkoIAFkS331h
gGUArD5qCmvm/KDrqpRnB9hM/Hd5+hU3JW7GPb8ACF1EJUd4G8WoZ0Xw5XgmiCQRr94W4Hg+ouzp
/+HLyML3rhR6d1meSJLQBdKUdWYXE1K1uGJsZFTtQzlIHdojoTH3xxWCB+n8L5uBwxK/uFnISPMJ
TQCjg6K5SX3eCN7qgWM5PlFDCg4hfQ79u1yLkMKGvkThO9ZgoFm3gxDw1PVoebyf1Ivhhp7g+0uc
inOP3vggRr0Xdn7R/bbIDxmKNJenYc1Xe2/i+5be2ePFoZ49uUni+tlMSrBEN9omVjDeq9kOiwVI
FXl6YUhHP86U8QOYW0b8SfjxnuTqapqbo3RoYq31xbSDg1r3TzpaQHR5Y3sIM0V4V73HKUnNsr9b
V77AQCGk19Ylca5oYNE2rTqdxkFoYyUvuG2xMGa9rsIw2IxyRsHuSe18kpevfceps3kKTzo6yml2
0qHYnd02bV+Vhdlc9KvlT29ortbk40WX5FJAgEVfsimgaeqAfX3V4z5Nrxk4A7usKF4bsCjlMKwR
9QwlfWYyzH3r0eiMdy+x0zzXFwxrqvP5KpHVG6DYUc773cCzX2yQAJxBntNBVOmUOMypuKdsSYwR
xVExK1b3srq2As63VQXOd0rVIaW5Zl/y48q08raaHDykHjsdLhh3+9hjT98qApONLNqshaevhefM
fDXvtykUzF3ydN2HUIB/AUagjMP7r+b+FZxRtu11uPKvklRCxAgm+sspgzmdeCVjpVSPX2Z+wdet
7qk6ajut+gs8g59eNbWT1/8vO0i2Xwe/tzDR8RQvB96fiXS5wIh44Lr/57kGfwei0/I7/inWY482
/X9yC/uyLPZcUBHU8wGEwWFoneQcQfNhBRthGwkuI08F//erp34RlvPXXLeCVEZcPi9JTBRuHi69
3YIW1oQdg027XiZg0WZB33by9BZ8jrE/BbEOgtL3XlmGoBDCzsxq+Yz6FayiuGga1vEWT6FFcP9V
2Lw4ZbV9yjRjXSqVs/8LOAI+RSYiHd695EAF+ymo8fs/bbgJv4ReY58ctchCxvlS0v4g5GTNjEv2
pttOJ1G/zxgeS0EO9JmkrgDxxw6OwEDMz0Kv2GLRRjF6A6kxHQySaESgjplHu379YWWnPmMt0K+v
4RP48bV9rKh53kYgzEm0zBX+7K2QcCf06dN8PSZeR7oCGG9aahv+afX2esYS645n0sMGkMtiyTIl
znuMrH7/oFsmTRtWnY0dFaNPkc3BrK7hEs1fX8BH//BcPo6m63Drk9BJZgJSTn24lVPAtL3xM9NB
qwFm9YfB7np6AR6dMQEe2KwUxvJKPTRjIgYXObh1j1VVnK0agAM6/WcAvJj/FKwI/yP0qWYLbOg8
XUdumeLD1nM6O1+3S8xQ/HlIt/I2Cqlu6SSBJ9shENPaZCuMVN5Z7kC4UuSjCRcUkCdHcZNY3g8h
nGs53gyiLlLSVPQZff4EbmrMaUA7oWta6BxEXU+Ual2X6sPZEo1hHcFKWYd0D6NxAyjGrhnHUKuM
gJo98KgH8bfPCbSjJkBO6dksyA0o8C0KvTdyhkLbBP4cOD9E6eVhfWU+Hdb0bK35MULu/MdE5Ttz
SJd7bzv+TxfCNAB6pHXnzzow54hGihM+2ao6h2jjXfqt5KxAiEucA1znxpKmL9UnX5aP2D1PjTt0
Krcp1QcKc/uzHanpDCZKU9RN40DE7UScjsJzGtMmTfJm/EE0tgAVZqUsUwLlFjnYYkLUIYM19Pep
/CKhU3J64i6TioQ8zLJpLUbCKGtwgJDKgNLUANeCrPqLigCCWheUgqZMnNoxFBJ7RX7osF+lpjYS
zQiBuKnLIM3eCfY0tF4XicBAAxWOAX6SaOrYPxZxtg+P1HUOe2lytIlHUjMrVQ7HNrBnATup060j
utrfjaoq6SGutXp3HJPJyQucrSajeH99yoBPnrFyk1875bUnwAQA3UlOpMoaODHka2OrCLdA2WfM
q9VbNa4U4+ZgNtu/g+skhdvtKPnNwo0MosOEuZ9bmgXF63kIMCqQxBnpfvDELMLrYvgS4LASgBV/
iUAZECkM8B/HF3BtzhvCIE/C7JdtjFs1UmNthOlPoBXS/7Kx3begN6q62rlALLR4DSeUIEGhy5gb
oqcbRdGqznutDT/Undh3u1ITYBqLoRykCyJyTRhO3xky2FXQivsscaq8ruWnRy1VBupfTXFvJ0x8
sf0WRjk6OipUuiosfNmpUKjjyLuMHVaFHBYxKAXPwfeDrrwHzLfcWavIotImgJGvszezDRUhTErs
LmU1suGHF7rBrd9hKa9RAkDxSgWHhPftvoo8SjlSl562XWMs8Lfsj69W0dAbZGtGFO2+yek6nDSq
piKAXFM5d0MZivgrJkDBCHaaH4E1EDMCFYYvcLleiy1MfkvomnuS7b1649h/rJuTlEJpaLP13XQT
Um4uusRHfheUkjy5MWR5jqjcNWILydJwTxfALPi6ILrvI1yZ3SU2Y/SKk6bQ+T4TlSKZACQSUZH5
hJZ3RekolViAEUQDd4pMaSaNODWYfiEAQ6fiO5g0JAvI08/VWB7GjhiTWR0iMxsa8bab7+j0Ay3I
RE568t1BMfVTdCU4NBqyIZw0kdyrdeB0BIj5gyFypyMIRXnMWd4rKupQRU3AzfMMaeq9jzLhzKiq
YYSbhewUbHIDKInWDOFdH36zsPgl0WK4Jwxxeo2EOGoMx2f6LWXqItgbuV61w2FdkSbO5G9dvMQ6
hXZKmPcNicq2tDWqmfunmxO06p40Icd8LGN9nj5qUBiE0FoToLo3Dy5HkIpP/QWZEJNN2TT4BuXM
NdAc0XdwgSzwA5IfhKM1bPhHoi4TaNrzCJPL8QvjgeOYyPy+U0cp2vkdAf/RGCIBv0QTzy1yS28g
N1onnFS3dKn39C8bc+k90Q7a1Yc1ZZbrCBwRYIDN054Yh4QPAPypJcR7dQO5ISb2i3bq2h3YZLrJ
mfhqGsEoqicV9hKeYjVLIOlSX2/A4cVvkrhSQh+TeFV6Ir04ptwucAbJJmzEJk0NHFu0jnLMmS2z
9mm30DjOAHHqmkCQCd2jXe295b8GfyGKYU3WSO90kphnlZDz7Av2yUlUOaIW91sWM3+bulAg76c3
9FumYUZIjshhIxMirbEBurSPaRNgVCxdsC/JthrBfriYu5H7o5TQI2a+wI3S60n468oJ8pTdbku/
B4FDkdQkI5yZr87NzaHS3GMKLkwLUD2Rtc63i0v1U52R0CfGbaIrJ3oqsZ0JgFh5PdPIUUeYyNgB
f5c/gxjoK2sDt7bu+FIQtjLVjLfJESbfEOLFsfaVHOCOtKUwuNqXeqOm4MupK2PUY+f2Dpx6glHj
SiJqSJEo+PVdBUYe1Utklrt5jHch0CbexdAOiKi0KcPZ5HCJt6p8DOd10XKzZnnCsnFAVjY+3WSn
gLPFTzp4tnvaz/B2NPOkO6v4cORi5xX2EcMpON0MQJkbhjT9XNefKFUSvoXCUGCGQQ+urPBgDmKV
xa2c5XGI12+no2hqv6AeahBxJEdVDpJ3Wuzr+q3U7zU5VmSiBJ6Ii+KnPZUWjDTuxXYQI/rmkOZT
hSDTVxlKx9Qgs3Yc0Ld1E0PRe3+t3quiucK0GP2rZKXcwkGkC9AyvAxgste4n15uHLmvtnNb9cTl
ZL2NLR1i9RjkWvHWCIqY0+T9fncD1lgotegOUQFnpdT3BZ8wZFOUjQLwO+dM+rTKP5II1LcBUx4e
hdCFHKAaY/FPTdz9x2fDPOGqLDoL3A/qy/psfH6Rnkk9eRll3wm7NkoFnfYd2fbPrOdcY0xduBfj
xS03Uqa/TuzFSg5Gvwz+HH6bmUWtQwq+xwJWoScqrjdAJqVe2a3lUKD5N+2bNcabaPU6BHDoDJK0
Qy/wcXM0Iqziq9fReD/9huc6p1BHEArS0kYX6RXwuTEDQcYoaNnROU6tS7BsMtwl06bcD1eJE5cd
DUSqF4C2x4vwfY8FpdnJkj9pQrXN1bYg7YGBKUiDJEN522+N+bTchNhhuvPJGPatip0qcfEGR9WR
hD8zrbldPf6T3+TXQLCR+Uf4a5dvsrYh1oEwcOndNpEnPzILgDTgrNQ1qHcdFBMDivRCRRBm53oI
QJDZL8mzG6f9XZ9k2lJzDbdUAbeT2bisVXJD+x5kKnVpwKl5l3mC67KRS+Tp+KfuvGLOvWEldz26
qhxg/7k7avdAxva7TdKpXr/vtjgq027s6BaB1BHHyGLSToZz7Y5bqCOVP9gfYBBxkOeNDGEib7Dm
K+N9U2Tn8qaR9EbokD0iLqoaKuwi6k0JgAYQOCVBgK4fvCzwin7HceYuakFGCXgi/I1ApCfKsiss
InCzcxTrqehjy1WFJoUsgSTE0stDvMsD4uvmIQec9q60IJhZu9ax8NWaIh5NpBzxhHAV1k7+fGwJ
tNYIzIRmuUTrtlIzruFcJms8OgtzXreOsRTlxr4Ffun9L4Uf0tSgH/2YaEwPOvBkpCap8rcdu+kc
QRkw1W0mF4ck9Vb/LFV7ycHJleyWaPbWRv1Zfiqu0TriGEiWZRpKwVpuYaAgEhkXNztKCynO09i0
8O6PQsopjF7c6hg+SJBE2Bp70eEi88snSUZU97hvTDgIMAuwRAzY93x0LhD6YA2HOwVWQ4KrzEj6
iHnzDj11K+nN50KYWWUastUH3ffStLRVmgrpxgB+w0+1EGrDPrQyu7PsLLFqw7MbFYx+qgWGgAFp
JoJoni/r00dfi6YvewRUIYMP3OQAwTtm4WlaUgwTlCVEZbjJ9grwqNDNtHmox+XWLEciFJT4fpfb
uwYZ9CnCeOfNovh8+4bgXivIgZnSgmDuurN3Ze6YzH7UujU0bkYM5q9KnNBcZqZAqhKT5I3x1Dy6
g5zq346fOwVrSQ68lGrHXURUg6C3w5IHndn4zfgtKlLJdjsn5FVFWh+Ce3GYQVTtomV9qET/F8lG
KVF8PeB4RSKyZe9/RvHoxMCywSJAgJqnDTB0n6FjgcbsF5vCbbWEdGrYhbIGBYyz5oupIM+B/tIq
0Ytj3o+QBh6ZzvcWRY5mLZO1Cq69r7RjcrLWzpbMZU132D5W5m8UuTb+nzsMHFvuYC0fIf8YQ1R7
+dmd+ovaXbzXi7NdsmsZ+TMixUbDF9vAkIVVLxuyENIa7kXELOgwwYRxNJqIMtIn43NVnqF9uXRZ
3ZfHaXbZI19shAuMHrdJ5mmtDzGKgjpUMHSWQw9wFItleJMOqGmuOkiOONor7kCJQEt6kHAXys13
BALxg3N+Uxa4jlei5qDLu2OUpPtlOWGcw+hPg+5orui+jnqUiggb6RvWMHb1RXs3vgS/XoMLJjMX
+lSXMWeSY61sYRJIXWyrKO6rRMUBhukWQ2plhos+SvmOJYyVdtT0ynN4OzxCGyXQ3kRDTL2u6s/o
IY0ttQyMKRqukHkc80Sfdel5OJe7vfh6TxdbM2B8Zj4s9xpLoOZOQKywOBTSqX4/hNOXx+KcuRj3
GHtw35r5tNzNSIkWDrj00uYjFfdwKI72l/4ddGpy1h96SrdDKxYEJXv6EIX2YDlRO+uLghdRo6fv
Zc/QAq8p+sm4To3HElBiu+FdRW27vDSMAOSCkHvZ0DlwIDGBEqAq5QgXwRyOou/NBVjndMPlshxP
2+7ppUwksCdRogPk+k1WPYZebIM1fSM1xJoNNsXVuNAXAeVoOd7tfRN0o422VON1sQW3V5Ub43YB
0j9zE6mY4fOXizQt3M+OiLDCDR175CgDKZXN5uUJJSW21jCWRTEGFqLYBFcNxS2I0prBUTYDBkqq
hZGOUgLJGVsMepEbyp52vnmgpUWUpWklFcc98sIoF35odfDs9LJOcJlaPzbuGBd/kXpswm95x+u4
Zj8sgFXUsZWTi/M/v2+tqs+ouLLRjJHuKu0tHJ9vyPDgXaWQtIhGZr3jAIQMcaeW/gT0u1rmPyI+
0cAFGG78QOrGhtDTpyEIILsTkI2KjXo7nIHIGeh6qE78oSvZsS5NRiAlhJU79flm3dRzDse6gms6
BuqHfDSD72Fd4J+NwXDAiHQRXpNdJL46dYF+u3C3bbd5bk+bxOffVDXQSv89MiogaUyPTvLye9kn
xLkptqYVLGWSTpIbb7rY4Ion6rpFRpEPKDDu797J/fq/l3N+Wsoa2WOpOK6CNvSu7dkXu/lee90G
jJmTxsR36EC0mih0j/LMqI0eg7f6f3hcX6GASN19No2/ErysUl1RhLlRHeCOV93UhXDYzPa5mFPp
1l+4xn7cOpgxvv0rHoPN7VCktifDHlR2q73alrIXhjB1Kl/KxpcoOf39GP+ruezYg9JmeoU5h34e
OJcz5h8oYhU8Qe0h5/L0Ch23wGL83+wHRgNo0x5OuCGXNO92qbkEpY4wcgdetGCOQlEJ5Ktg8eKo
lh5s18CIAIoIYLX80mSd3TPyBqC8KM1Q/EUf6+LNv9yCxzzCV25/fhji2wKakOmxkriBRGvZ+CCq
oXDKm7tw9+yvAVTgv/Umqm28TtkOpK40paf1FSW0qQNrMsurhtSBThI0+d+fEuInHWZVRzLeDNc5
aDi49VPw5jW4yzE81lxHWXi7tj8cP5woY5742FJiPIKcF1KW5w9Usn8tIsFxLaph9VOBVntHgMax
0CdoWvpiAuLwiOTREGw5lHPKlz8AwlpQPT8fLnSLi69gDJXaENomBm+KQogZPUvhWn0U7ADKI6h3
ReRcnDe/5H3JYDVvOlEw9KVy+EJeQYi7+p9oqzMUTdOn5uVSjU/kiD2RTgoahb9NJj2vVQey68OS
wiqDjmCmj9RKpFiwpOQZ0/A8mFeWQDByt0D/6OpLJL5NZcBwOpctNdlXof1lCsLH8k2XVACkZ5En
n0RR3Jy3C8Gn6rgMQkWHsAZXUbmWQO3JQSw8QF7n5ZSA3e4MVXDjKuoPXqe1YC009r62hWtbZG/8
5DuyBU6pAFxv7rWgnC68ePT22CJA0qopajulc9O78p7slMALmZmi2BZJrL70/YlyXRiBjQcG04/Y
aPnfEEf2jd1GRZWgd+SjPoDftqWSslPVgobuvummB9fQ+PUxnWBdzFuu+0E5+cgFrWd/cViOuzvs
qzsQvzmiU/o5iW4JH/EFGHw2AL83N93uNgpao3TeQnmKKjUf4NRP+oGQhPLpInWdnncq1ROACPov
vOh6afESjd/U31mrSoaJEA6aBB/uuxCoHyBlR23YLvBgI2qnAKOOQRqE8vOnW4ccrFUvAneczVpH
RnZHZvqg+pHYjbQLjvGcJwmQ2LcHMM+nCdMsHyOI3EnJWrHDZAlGKaHBrQbV0dat11h3WR/cu9Ub
wpzBzvWoIPFrFOoPS25WwFmBvulhFFwRkZwun3im2yNojp3zRj0oYk/QcCTXrpYh5TkaHf0+hMRd
niqu9JKvjCRhtX7XZ2MGs8XM6T7M5yK1TQETHW0Iho4ZGqtSBIYRfgu3fk6odTC6gsivbwOUcgF5
VmiT0KLIRzpmvkmsO5T5ew6frK4E0LpIrC2+mlvwij+834kzCQrdODH7/ybrpFNx9xNc8qQ7Ptzl
YDq15Hut/1rVW0WcOimoqk/1axHSJ/+GnC+A+7z0RGaFxLjvtE+Mi37SQ5r0KQFJyvnhhnd7P9Ng
f7dp/lNUFw1SLFv6cbrGUFuohIX3i/9uX1BsgGBsd17kVtH41y7P0uiL4ISijRF/Rvi2qtS6q6gb
LErdoglL0mH7aF3lOrBDt0ei3MYY8IZpWCbI6pxSbVwQm5h/tkbz57UNm8kopLgjhHHWo74B6sf8
HqqppLLmaibAhdtE2ChlTS4eBNl49fEb5wG56IPnTZEqiAjAttyCfDHw3hB0Efv2S+gW66O1yp71
/b82P0vfmBqAMaU7dKcQbaacyorpLgTyUFiAH62P175lrpRt9da3tQrHSBqYxJccfZMQtGD/pPbY
n8sF9mgph/go2AMgUDjaiWLa8DbYXYCrizDJ6JD5zGw0KGvjnF7AWmhSlyAeDksfyCDm38DoU6ou
JoQjuUgEu6u18oXf2eldjH8KCEaJ5zvWDPLBUuq2sOYUn5cTFOfaADWrivb/EHCvfZBT5CTb8Juo
EPfINGAQbQDekHU9eCWhby7MJJazpUIDuHl52NrHKBtw1PM3TsQ4Rn1wYwoCmt5ZeSajgPQr1VcB
0hW1JSVXNNuYk+kKRpgjYJk/FVSJUB/41PWGnr7ddvIORXswLbUZV7TDR6TWJBdJY0YO28Umh1G8
VaMAK/Rg7GcIIbsscWoIXZGc4e3yTh9v82d2XG6hyLAC1YtO7NJTsXSr5+IcMfm+mVrnqXw8qeY4
0D1YD9SbozdRZbCV0chZrYlQrQHfLTaSDjaK8lzdTihg0cSBdDxmOcijqXMmocNi2+hrJOHdOXjL
HNwRM3OJaW55sLvdlF85/dXyK6EtA9rv3Nnovm4pidxSJLVeygu6O5FOzHNInULBa17wPX04IgVC
/KQGpa+SoOVm51Jmo4/9QXBiYJKMLkLAiFq1zOxP60Mv7cyGURswJwTnLV/CY4ypYgrL482vXyLQ
VPswIt4wVOqCA+roLgfUs/htBDUnGcYEnl238RVfr6xaLf+i3FLEHwkkAI7CW6YnSHHDubEt8X5S
PXtQbeeLrqlNhSuuYKMP4wxnnqMLDEPChVBOiK7BsOMvfZ4KUW2oj9FYlnAtTH7e/d8m4XHFa3/M
PJDq7pSR9LcjaRr8K0ahqNHGSd7L3JzkegZdSaxWE+RmQUovh96g3+qf7pkPpkRCJHupeNz9K867
ppTDr1o7SvHxz5uEmtYsSbezlbI3UX/NuSotyRku0rsvxYkAS1Imqk3Er6RPNHCyppm4qPufkE4M
7oYLKA7j0e4smd86ixx1XvPYdIVbmJPn01jariBmsNUaoTYt52DkGWMS7gi+pB86qkPlYkNiVUHG
IsA3BuOJXltAF6nZFZkXFbJIEFlomL4+ai0pl0dHypJfbq0W8cKcadyzjPKlqFQIlbX+tx8M0Oxh
wRQR84r5004ptUJWaplQYe2BxZbJkPLDYkcxsABHIXKB33Jd1yy3GACyVXJwg24W98OUrXQmUgZ6
4V9QCF8VzW5mUbALmq2vf2RL7o6dnNfNPxFeyvfbcnZ0pwHwO/oQYXw1OCuhuYKM++xtDSi76YhZ
3QngAqU6b7a3u8VfMoC1FsZ+LLgPXR+IVe0lNb7U2Hql6lUwif3Jnu7I4YHxqkmUmTR2CoxKJHGe
f4HPvdMog80Ke5D620JTqacXhvO050FxIgxMqVGkwDZXUGvS3lx2kOFtcBRRGcPbuwWC9iAn0NQd
tjrt1nLkUh/kg7Yv+ZdroHhae3+CDcD0tUKttPHCLdwVY1Px9Ku9kax4FiCFExazsuDpyxTvz1Bw
aqC4qjU114KTr21hbROUO/hus3aPht72eCBd5arI7BCJg/l2XD0snJjCqlgzv9iUWEcIbX0FY9s5
gPY29SpTPK9bGT5LKF7XD9NLe5tcN1cMX9ixrNZR7u4V1dRAbaYbnPXXgTtTwhbGAJnVK1AxeKyW
34FCMwLJwTp4m1YQoc1bXJem+ZTAnVeO5zgjhp7WA/Uoj9UF+Jm9D3zURWfJoWstWFapre1CD4DF
nCaCDFcrT86tqUwiyFxlPSY3zSKC1+F4WiQ4Qga8xT43Yt/qx3GP293dwRmy4dEFjtm0gS+kPaxo
CkkgGenys7OS3p3+tFs8Cc+v5unO+0Tv7qTJGqCihHkVP8Rg65lwLmchn8fuaXSGG1aWfMKeGbJM
7OCLZtnV709JL6CQ36FMLRSMscqv0mfV4P87D8ACs3RI/OByWj/vqdBqP1/8LyV20iotObon3gZM
Bi4WGT3gBHjNwVn1XY62CcgHISj8zLoA6Mkr3+OJNuTb/W12NNpEfvhlzdVo9IQTlDYhRNGU5vSL
MQuZ9lAYntBugs8QXxbMN5yAjzFwB5JFRhS8s3SJg41yoogFX4l34sD5DNy8urD5l0VQp50biGhG
36I/dDLbzo/zvbIevVlb9laaroPm7qW0/VxiVkFK87WWtfsqCjAn6YXl9OqWIskcmFpXB/jP0zOc
5kYrz+6kcKJe1mgHxd0ghwd8tKSsNi2/Fiyjm4c2WyMX4n7wyz9hc1TKFvpOlvxjXFTBtUM63mLG
u4dfMFj8XC0xG+x4+8y3SZLxKpKfRVWTysmI0L/jiwXJjbZVxWDsKvSy/t+hjFBCKAKMSnfMUgUl
tE3sTz3qKGjvhtKER5WTbG3Sr0rP9wyQ1Aqu+ncsgP37oj0tL3hbBZOdJm6jSWXiZQKEeR59T2aH
IriixqZX1yASySTxflolRS96ZYVO/Ev13p2yhgE8EJDLAM35ANsMx438IDqaXMntpkSpWxYWtILt
QFpCxXctQS7yyvjM+6Kh6JEu1GMM3H70hSwwiocxMOs7Dwie7HJlnpEaTrLuiNmFYip9IYocXMC9
XLuZrrpWTRNuEk9aoqFu1OddwrIdQQocpb1pgg1ZkuNWIwKBHcTlDlEhPZw7UYWcWdQEuSXyAZhz
qp6V437tM6lkjgbWVbwARVNFaPTG8oYFfc+FXxu3Ct8q116vjJFDBS654flGJr73U669uDuLulWY
kFYL73sf6jHwW3hpDVU7l7+tHPfci/7hI/qsoVajrDcxDqAMBu4p7FQWzX2eH6CeMyyQ5NTLQbBN
8SMZHzKEsdUQYhR43DZQTyQ4Jdc7GcnFmlIaKNz5dMu/NB9BgdxVEjTEZfusAAgSHknHVCFi1mX+
nVz3iFFQ6lnyZzDtRpcuJ12AC6Dy7gcCIucPrz//zmNLfhDzBz1Xg3pD1qLnPl8EvUQSn2a79dYo
lzw2aA/0rupHw/gzJQVl1pSSpbXrEWNuwigeHmqlg9Cl6nn7JEcQfZACi4i+mlWxKAp3MUc+iI9G
JetKwpbef6M6wxhlB+5S0gS5d6Ms06olLj12F5ySikkVMlEBaHiP4jrdYsPPU0eISEbBqYdpuWU8
IwOTHQtRdhpyS2h5S3GT2URiOEYc87TJVcLrlzA76xEbtsTYo2t/kV4yYDoKz9dlXD2O9+9rHEkX
b31XpBtz5ZuKB/S5vUOgz0Q8pUjJaN9/EKtOvkuOjf6UsQhsyGePSV6/pULNUfEuLzQ9Qwp51lRY
/+9BRmgNFa/AHOpSSfQozBRWUawToRa+OiMmdeCmP61yILox3pGSyMfaLamn8jRD0Ha2r1Dkvi8X
rc0vWF9YkK+3iNH+YjoOQCtPZQCa3nVC02ZXKVmFnmI6hxobGf4791z55HS6RU5nLMwWro7oS7St
pTlelF2aKaThmqexNeeZRq0cUw1VFytkqaO1XY0gRpMdeCzOgJOJA8im2d+BKDKGe7n00XT5kS3D
M1FCz4tA6kMgZBz/VACZabSOwUgOqYaFLjuZZcWi8zWRT9LTu2wSUuq2N+paSbBiPuRqLItehViJ
FV3DbSSSkhzWGmsHPnJQJOspKaXWCM1rtLsVslIok8Wac8H29CZXyeeYOoQBgb5njRpPVyJdY7+G
7vxsU68PLrWBKszFK6TfKGFEuoJ2ORl63Krmod+YDOGLp/M48748oKAUbWUPRN4fuWjCbZmyQ3M9
nOwPtPhJISxH8DdO/Ma/D74Gmba7JlgIPxWHc8V7RTvPGuLImYF2LyQpPdJ31HB1Uqkq95tTKLaZ
GeFx7egr0uYu47RUg1gz9t1d18dpXTL5TsjDu1hBU+sTzgVoQ8rc3f29/V+K2AWzP547yJQQGhd1
p1rvhZK96xKFyUgqIxBF/mev7q02Vhdjhax5zPhF2xwHRoJtapAsq3LBMfZ4LJkPGmoY7Yer0qd3
hwk0yaHL4t8axbgUcgRMsArSXfuEBMqfm+OmKs8CWJmYH8o8ZTWs6PlFuycqHNh3iIK1hICioA3R
HQ6BY9my6tb8il+z1bt1O9EXJzTMIJbo+jov5a1DUx0nc47aYDX5Nixx8PVUq1kFRS0nIrF3TkeA
rdhqHjb/buIGH5PeFN9iRS/q6BeiFsBlJPqzgP0QP+Dhlis6Vv6m6VQmEP8dt4+OSAmo3UNCmoUR
OoXqKPmWHJRJiZjlqM5IJxkdvxNOqauS2DufH3QtKwDTLsd0Nmp5UqWgR5FDB/KOMcBFGsFD+DHE
2TYTX5/5ThbJFs2vpThsUhKQ1vnyR7ntvJJCxRwhakp9XWY5Hf0UOQ8Kyuh5F1U3K/bHu1VJn4+c
9XTKfzEND0qq3U1SHGQp9wgVDXgjNIJdw3x3d+jK6XrdGjNyfdX1+qqFm3YcvFumdT9BICAXTjXA
ZsINVZaYAk0mUbxryNFPNMKYJvdplLbwg/+UY6S4ZPBEGlbQNsSlIbO/hZX5LTLPkU89dG8DRSfY
6FVwiC/6ndfKOtxbVmZprs3dCXV3uBTRkTiZ8FALhf64Pobi0Fe0FoEU9k8l4KwheOqOF7scZQX5
6w3Y9Wqa4GUgOiSr0rrWOygnHRkS7ZY4KX1f4P/d5TpFBhMZfw4Hw54MWzkhx1sn2WLMN+TtVOvE
tehNCkVGF3mOYVMfVKS8JzLhGnSS5b5Xsm+0zEpCuehl2N0Te4gQABJI3dssJd10t5pfhDUsi1Y0
+p9OEhwaoLOFF8CnbgxVOa9aTMF86cZYLOpC1shE89X+OEse4Jt1cH4Q9FCEV5RcPwBiS3cMwlg6
HkSSYmCU0hd6vIyeLjawNenJIcaL0wAwcrg1/5PGa04s4sszdeZwVU/Icqz+5DiXKp3CQzFDP0QP
G9IHX5rfE9XnGe3lvCVhz2uplPhD1M3JIIpHst1a3qzfVtvfQGFGU4JNGZ+Yl9/SO0rP2lQRNRp4
op58MP8vxHQDXswAyyMeHRNYMbwqctfOmSSjhRtq/cVEloEF4FTVNcldNLt8+yyi4hhp4Zh8BYTp
sB+hxUpbSLibaAPjjqidsJo5Bu3vKR7VsGLiySxAFWSLczWqTNJEKEyAf+fFqLYzWjl2XCiUTYzE
EqlcRTrg4mjKWc4To2vObcor3ym3laO6ywLLx2w72RwfJa/1/Fz9gXxUoM5cIQ59vf9ooHZcRmeD
efuRr4bchHyZGJewjMumM2yWhBhZ889p+z78f5lfNspm/Bv4QpJVUxkyTfzAFodbilUO3Jmz321p
Rx/ry2O1lVd5Xic/WF//V2kYogJCoEW18gAXIRjhuzfqFKf1syxMT+F842yFGP9SXTuuZOXM/UG6
Kf3rJVy4wX+IBjdGkluCyme+SSd76KbV8ERMclLseoWYIkb/pB1fqC8fBkjS6xo5cWLiptcwuzxN
UijisjN/KJQccKR6ViPXQZJt9fYg9J0oF1+aQuFERZv8QmkELTw5Sxusg1TvrlqqNgTdwflOdZdv
4yWdsI2Wu1+aelAjdaHyQRtr3tKt/lc08nvHCtXBHHL9rjepd4eZwmvF98hpumrsPn82YtM3z9DP
8VrOMRuvWp8n6eupdYMWfOomx7ZnjD10hBsI8SJFb/UjhNmWqe8jZwk1qFjPENX61jqQRgQ3lzEu
DyRU4oRejT+3piqNC6Vzfv47z9/XJhbA6RT/2xiyzgYMZZG/3X1UMHf5R/QjoQsOlJKA9zWUD08J
YrmclxjF/W7YTjXnhx4NfxtPDasAgbb1jtZKaBd02+RowZCo1rDV+5V/dM0pMEG5h8BCvDK+fABi
lemRAi9F/AjkyJNlMZQKke2SqpND00mWk0wdky7r1nf//0iS/hvb1NPWm/WFxaVT9MLoqfq2QS+q
8xL7wbGHZNqgbABVVWY6Uq9lADA2Y8dlBYCaiqrrJMURK8/zNiPpNosfZos5XqGApHI+XfE0NKUH
VMmxftYx8oYvjmHF3QfD2f3j9RxMYJYULqVCEFt61yB3DYloozBs65aRwNU0vkz6LWAkowkeZXSm
0N8k5xWPzQywQRNn8yGPL+jdaVmH66+bHejxDA8JXOdYA4sNXL65t/qfLZ78QOVha2fJUH2Sm2cB
kFr6G+YNphAmE14291iioSJ61SPt2nyKSQSV0O0jeqFU4JrskPoM4011iY0j2FisuV4EFq2lut/Q
1Xe2oINGUPjebLchVcCqidvlri+hS29JBa0Gl1crVYGOhKEJnVSEfmTuCw+QJk9n8LMK7yVtFcNK
YRUHWspwSO3q7TL6TLvxS4qMlMvbJj9PlpGByhrIoo26liC47LtTTFy12HCrE39sv8MzKpQcJqAu
cXN8GQ92NFeAYjAecvcvn1Cal/pNsi089X/R3yyUUOUTLCKep8Fbjg5VWL4DGmNKs+iYTvGEJPpX
KMG8jV4EslsLChmJWsd8Ejkq0JltA/7PELbGJs2EO5mkJYnHjoJmR/X7XywJG51/+4VU9ocAanRk
WJOlM9cIB9wx+4TiHwUbjHg0Z445+JFPFTTeqhAoKPz+D4sGzeyRqI+HWNPSBiUYGcOkx6ovAEK3
2hEFPA6xuqIJ18bJ2wwHl5Z41iraHPK8S3aGkZWgvkjUg5hp59Tq0LD4DohsYOSC+QC5I7SMb5lG
ajvKPybYwjp5UZhOSviOEccJ9+OzaroTELrPJdDdQHepEC3YIRuZd8X//QK3XJoM5cBNYflAHXRu
qbGjMWGfyuvP/vaRNee3ZsC/RNWn6sFb3taoDW/9AM6Xe6o3ioL+i0LC8yJVTMoUbt6u9weXJQdH
5mV+J3NpzfnnWTcLqtBup3NEQY1dkW9wIOTePOnLpLF7+Y1gHhKl5gBdVo/wZUO1AOKEtJ8VnBdP
R4cEBuALtx5MBPcfkOskc4i2OPY+z71+C1toWbvZ7gqTeB+vTOU8JuWda3SyRVbCLGi3U+LVnCPL
FTC5xsFs2LFWItHxQEyh0RewR1G7kozt1egybREQ5/BFILWYqnE1zudzxx3t2tt2FmiCOGMoGxnk
VwyNiMdg+9k14WY5oKLjKWQAErJKF0SL+RxPUpNT+PAtTLGQxNAnrD2ZFsSRoEIvEsS7+38ziQZM
RM6KSOTWSpqb3y+m9RTeMl/5+d7+GsLRoB4SAvwhpbJ4GcdiH9ATZ0ctH3ih5LNSa5/eqOMZprja
W2P+nkLFMFcDGPIuaDikYR1jhG2KFIuXc8Xb6ZpnauPugAAd6gPcDnfjgyBAdQYRKfPfFfTgvd0g
Cr1KS9j82Tt4Ts7R7Ais3zPKM4cFScBNtd8eCArFx85FtdHmfl3ikyP17RbpCUrPiNcB+5FUqUGX
3oriXproTjpIW5H3bRlnNoaiZxuwuoP/ZgytGZDWwyk10llkgP1rkS0XT2Onro5huhFnMmDl6BGQ
hM1KkDIX+QuRsvCLcuRFoRXkvsrezFcrvfWGa0czaFL36n3slCFUwYqf7bEhAOl7IyVeD3HANKTv
Elv3j0WEe5EiZRxiqi80oF2GwMP6j268OhYfTXfHTB92tlgJOZTXT3uLXIQARtEMArrRmlCMzmss
oRCvDDIbNl7E+/Rv9WYMinxBFQXTxA1EjK0ceHHVsq6CYmf3deeq3Lh13fNues6d4ogovFKw/dnb
ClIFDS5FGWpJhjoEWWW4e1S8bimQ1cWdmoTYw2F5uhhhrWU6IxKHdff0PZBoOe0lMSJv9V7v9LUp
m8KFH9+yDW2e2syit58yFu0CSSfcCkfpEnVlGMu3UTgc5Y7jLzg/SMkqK06hMocJVs3wxSDzag6L
gJqz66LDe+XnDjpouiQU9Qa1ka8BDznBWaAehyRFl+gCkuAN7MDEHAGzfINrpwzMnfmK7bc+5ZwW
qJU8aEWnonoIMlW4PT5QNtGnhGr1yPkkfPPOxy4y73iztHusjljDTCTqMa2zLsjavO3KJB66KcNN
4A61/jPj6YWdnVURFvqyhGCXf0YlsdXmDG/ndbilXJ0yS/88YWfS7Sfml62yv6TyzEv7IG9U1sIp
VB3lIijhKrt9ej5sPvKMdGhOBMJMmyPzSIR0YAKwRDYXUQm1nX1t8alfVgzkVUGhADQILkawg4Dq
9c658sxRGA4U+/izzZiQfBSRGRgShEnP+fB42Y1n4gnjUGZu/zj2wajpVltfAkP4ySZSGT+MTfw/
w373BHWrLZW3aRp8yIiRnoKO7Tzr8OFaHY2faH43oWYZVuBtRtIixjfOQSXi7S4eI70JDwX7JF8I
k+ojsG+boLojkF3MVn/eGgFKdYFfpoGILZc0VcAYLQpERUAl0qaJLGLxg6WV6ssz9umkYUOLJP22
73D8uBvyiWO+ePFea9uUBzPfgj0jrg1oq74a6A57X21ca5r0lHE/hhLBALzNPWHNpGtAXH/8TFBT
vNBFIZLrgHTMN2BlXt/77UFITQfdJk6nxBCM5vJSG1knCe8tX8CmNVx3P8ZFYn0itMQkqdYNRrxx
VsGSmyybgdUK708BvqYE7uToF/rTAOe/cR2cNT9Dv9pXISpSGn10Eby1WlBL5HvwoO4PVac6m+vA
c+wG8SL1edf06Ywn/wydDY4mJMZKtH8bM6kneASCc1CUbmssEIzJtsA9mPlCe04YgKpxzz4NSKbH
og9CYxjs52XOHrbXeKjjJCc4Jctgre1KHrv/OkmOFEiKjnZ3fqZt6bIU8P+mr3vsjFHAUSN+EnX5
90qTMzFIJfw/LlZNwifhffF3hClC999mVcwxP+NoJ8AaBwLbwWD0dl9jDMc0YiLYzaQVQ/c/Fnx9
oyafeIOC4GYepAqm8ykZTWIFyaswy7MBIeH6qEPqwFxmMr4pe8ek8dZy0WiZae3OuCgTMeudHSPf
y47BCibZRD3UxvyHCprUXjJTrL1vshtIwWFJrABUNCQFCcfbPF5l4P7XP0H67rQGdBcxvPUBBE59
fCk8Yq07ZjiApaUdvilQdRyeGzZZ9IdeGYDCbSctQAGdDlvpHLO40z8Nj41sk+Jyk4XMLTdj88WM
aCdXDjTvH6v1N3DQBWxY6H/DslXJiqqHT7nGvvfawGDdN4uWx/xwTtk2sZIFSsgxLK7WD3zB8f3j
PD/QT2MmUqIXL4EuoAEMhEEOqb6ja0OGOlhwz2KTnRQB1Iy4m6VwS8airppZBenC55ftzPjwGudH
yX61G+mmXVhXlNqU9tMqFSrnf890s7EpzUr7plYGXXd34TwCqGd8qEtbajWgPy0YX+n+qr0KPi3m
a6NsvMOZZO/au2MJoEWHL4ccbuGeGsgoIIRm/46cSiUx7B+WowCQXhoV8/Z5XvXSfSikVDAO8m81
X49MF9rhNiCbqXDL/3YXMF/g6aq1Nqo9Ltk2/HZFIY+fZ5wm8mEyYXUvJ6KMjVzEriirQvU9s3sT
j6s6nWpkpquJO1EJuDriV9EXGojdQZCGNXIoSygg2Eb8E3q+Sz0K8OTb91bXyUln3rYH3gbFnQ0k
gweEPm/CGPTf7EIia5oBE8ItGzbXN5li+0dw4qCKbzpAPqWIAmUXZ3fO+NrRwt5yg0q7n/LBiBmU
QDaq+z4HcZTndqDbpUHcWsT4F87WNE2It80SfEiQ7g3UL/tR3OKHaOaZnkuQL2oGz53nohiiSfMJ
GzGXnqSAfG32kOflrSGz201zN8xGeNvivlwgSxyuZA+XE8vfYVeOkNfE1PRfbjks8okaO9xpQTfx
49xtBzruSh5j7qDVgRnPB1t0URobwgDzNc1rqZgQybimt+JMnNeDnJdWXpl4hpgbG0T0IVpWWojX
tlNV53phlG4+zKafzCuxyVZLS010G43KJq1p0zqcRllSBV/qvawaJw6r4/MGxkak6UJ2h+w39iMj
L+f5PRbd3ji8P9sYz++xOgErJlhKVvEilPOO01lJ9dd4EcKhbMFTuLnKOuj2rM1VzNGZDsDBfjTR
JI+MtXvHaOprEyXMijX+lbzlVKzPulPHwYU9BQEkemOPg3ha3WLmSUF7tQQx/tfVbSD7lvHZSNFj
NGirWBvK+0CMk09xkaAPNV9zjx5+mK/OX95MVYO6zxqtwLFgBk7+UOSki2PgA2LFP4Fy4yYovbMI
BMws3uiZLLBPn3vjZEktNbAp1gjtoBMKG/JeV6Yt4kfRh2ta0J5Bkkm4LfxaBmELQF6zTqVkQ4nb
QtGPYOVt24Wa66mNyxu+W1VXsbfHPGgDjE3huZ3n4b5/paTHvSmjyEJMxyiIleRQFT7svhPZf2kU
oXwndBtyKKjTY64OxXwPXz8D2lueRglZqwBMezQtD42Sp0H8S/lZ1/I2R5YQmslHSd8hzCseIEuK
D+aFZonIl5WTetxXsSpIjBD+8kpZU2qej1pXuq51qxXJvbprf4Yrb4rratUX5i4LquHMfDcdlCiM
fAQ5WngjfMs1NCFDh6gSSiR0kWkq1GFxAsPSXT4EuLWP7dI4bbu2eCz6529PDkrln12BcphZWxFQ
1fuuuEIEoO3fjFgKOK6XoLR2tUHI5VflW+EGhlAT0tyzXqO9sg8DDl25bBipcqZNbIxFsxDAEvEQ
1A/j16s9OaKMBb288G3JLdQviY8nL1DXYHR/eCIbqwYA69SMrDXmFh5brI9NjrO9Ydecb/Ibq99f
CgZUTS92ou+f1viOQ1I73FmhSzErmmiZCz0pS1zMOt65B+YABCKnjvYmt9ZCFacW/EkU8OPQ2PEw
guS0ZCWn8bAiyU+XVhKxkFnuCp8i+vdCuPsmkGs2yncIAs5d1SnZ+fz8rHnyHWap6OZY3yANaxqK
pXJOKbLijZgfufG9Q/pQqCFwft85dZJ8beKgjJGNee2J24KP/PIIimtI5CSD2maxVkvLmg5cudvM
O516q3WGN2jBIXLwHDYNAAt6WZLSwoYSA7NbOi6xbQHLP9iZo19iRs1MRacA2reToaebvdwcqxWQ
4C2YSp05O2I2AL+GlCi8VmZyK5KhNIfwegUMjjTc7RsJubiJo51RgxUPdp7ijHSGOGEMjdmW5ahh
hZeLTD+b8nuTG9C7DMnPw1xTYCvmyHvbpvfusp9MC+dNCxJY53qfYODUlE+iTOXUOTWhMVkyBRhK
t4ja96l6S4EW3dZQBhUPgX1i7vO22dqyiRmWSPEhxkYTFTCYeYmwScfd3udCktdKrp3LF9B4pUWr
qlDQ2Z++sE4W914QNOGJdbFsW32XLnLYs1uSoIGAbxWfuH96G1jiAJFdspkyVEmr0Ws1ZtQKaFFk
6GVFYjA/96duFf7XtdP5DJemBkm4EKQL7u3T26HQSq8LQ0pnKD/BiS+i1uUFsIpTPM/MW1GFTO91
5sWSQmSOVEa9Ima1Am/DW6QkSOaz4yZ6iU+OpAYYK6dKomECvHolJ+5ear4MI1srf/sglhpKNjq7
9YWzsLlvmQBiDN/cM2NMxcNOW+K7h1nGQZD/bP93zb3GLCdlkYKdR8veL7oXHv64cpCQmcrSL5m2
xSQvjg+sDMmnkE93STeouwL2sFO76v3tdv4+PAVZeRaTQYLztnElIk2opOFPkVod5poYz0mqtOKA
dhsJxZn+YcvHh5NI0HMrF1YJVM3T4w0+ag0mCMemzxK0di/tIMVdWbahXGm7e09Y+KGtdvHL3sqd
lHVInzfHeKvVunv30OjWMdSZwcPHzz/VObKje3sFjlagoikjgr/Nslufmoxr5Xi/pK41pVU0SWst
Jvr/2NWmagA1A4O1lXyV2qajidm8thS0lum22mgvDmfRg1hj7jhZ8hU6Gq6GDcX/TR70Hb1ZTLco
S+zAqyrqsTKg9VJUkv+logTGOG/C+X7/X6gBLXVgD2di40/Mpg13f6K1wV2kpfSgK9JCM22/U01B
rGWKLQMhrpojCeiisB6/tC1bPhCZQ4lU3tXoNWsl9+veZziUfWgL57ygWpUTVfor7G0rVb2eU5iF
DmvEXOiUCWvXO3z0JvYGPvDUIWcZedpoSXR6WlaIzDSzBk4OHc/h8bl5XvdfAe4UHUVT8KNybixW
ui8YNtd0SMRvKo8xqwy3YmNGZnb11j1+Cz1MFcutHK4dt7MUVF0QsXWBWLY13c+4sGv7ZYUvqna5
jEXbDOTAb27Dfi/uu8D7XPqXAsUWKpLnEI+WvKeb7GCO98do/Kb9/1gYWZ5HbrpcuROQonJRUPBe
KvV9F56p5UtP1jb0cctS0WE/BdVeJ0sFqxiVu0kQuBFFP1kWXL/Sv6PhqUYF3UAgRw4TwXtSzMzg
ZzmUuGGwA5fbLwEsMwTC8iuTEsad00MueXsVi/Qgd9mVYn3txwu66/ETH/Alf8SRctm8NE7PjuQg
DW6XqZpmIN3Vo24KSSVkiWNL7tamrvpYi5j2hW8chJODx+QVVNr7r+RXhKCshcHyvNUEjqE38EfX
7E0exLeB6006C8rJd8Nefa88wySGCFkmEoy2kc0ylLw8DEPOJi4TpiLfyhxIB6nhSbe7iRiK9KDG
fpf5aqjrLc7SkvIALk05hXHJIBpjGsImskyy2/4G0WQ+FvmurHCP+IrJAD/dc1qS+eNiflXeiGgF
agl9YmZGaT7bTqYcORGRtZabOxPjiiATccvAWE4T7VTamFLxhNyXCCEpcWdpDQeD5GtKQf9xPtYg
qodagpRK6gX/ais/t7f/hWCZX4gYDtdLNxB4cyDvbEQ2wWU8cxvtVVE/H+0OeHem4+RPgcbPb/yj
L5ERY61qboLmc9zhYNp+rD1f19yUL2f8jrSkn0QlVXkBsnoA0U7chCvJUX+VB26e/18roIxdm0Qp
nYWJKKp3ulcp9fnlDsCzwZgLsVWTkNe07LcJlX5fdy5pzJKwngrkzzDCUzuMtPkQGob6UfHppGQU
UpSOSi43gs1hp2VPqbhqonuOFPURbFASZJVXZ85kljpSPFDz2V7ebNpU83Af6aRZ1oSYgM3GIO6X
3E26/IjDE+ZlSZqLNUgf5L+QYMUvqL3RaPqXyU1EGrNkT9Ll3xxFbNLT8XZYZueZvBltYyA7kM7P
WFaxL9o7rD5hfOs40IwvZGUgfg+xIz7d1MdtbcuQiQpN3uL+UonKHHeEG/YKo7c226YpVO690HE/
6vxfJteUpBJLNhGlwhn56uzmcWr1wkAtIrqRiK8A0llRTiPIAEzsk30iTwPEsYOwgySSPikm8Q51
iGfqahFRnoZBW+syTMAGINTG4zu+8yOXpBfVWr7lYFFz5Yorr5TBiUWIRoPHDu0XC+9sEMi0LIrv
WWfeigJr+WQhYo2Z7GQ0aJtyJJo2g3iETlD28ZNd18yGuh3SZ4sNr4dU2Yoad9Gfi5XVRjEFmcbt
ShWSKikwBzQ39wT4ypEWsL36wSGS+0p2xuJUeg546jp6U5ZB4SS6J1+4pB/jmeGIB+mbBETr0U8D
hObYa5XI8//LKqvX6Qlhg3/ADg3At+0J+tsON98mWuR/0/x+Ix5zhO400/nJZUz92AeB6uuIyamk
z117ovRuYJJz8adeI6Q0FzFiau2Lkwnty0hpSDnnsgw392kuAju15HTirmFoQwG12AsfZ0XE4F8d
OhInRBRfeBn+Trpk0LbMot6dxenH83qtWHobU2v85OQYO6nqu765JytU3bDiXuYta0Vxbnhs0oX+
2cOI8KGAvQIomscsXnkl2O92CCr8dPiu3h/1o2KUcgZOp6/PRU0dQlxHhemlxVZmmYDf9MRjpBNv
xKj5CD6Bxny5Ag4iuybFxFDd1ujBN7CyD02hA1f2hqGtAbd2itlRkzuS/Wa0F9jGO2ejmRrxErJg
LGEkgfCmZHEOhJdefLHJyF18YiCYHu/e8dCalEcSBPAc7sjU34f4aOvbE+kyc6u13NCGTojnB8oT
L0rAe/H9h9rCAeag92TTPlwpDAX1q9aHTCFBTx6DacRpNyphMSZK/e2z0H6kRAOngYyOV/Ogxl6s
mqYeCrNiuQoyeEwKOiuPfkMGpGbHggm3jdn9xNm5wJec3kBurF016pW1ZMHzgPnlC64wpB6+OJb2
M7IEbgNaGIIYUw6eY/saCtTtC7Cb5uc6lymIZfVHf/Ou8B0xPwP3On1NVpI5qbZJ/3XmoqBaWvC0
d2luwund2oIEp8LNlOKdbfUQanlevnXb1b8yWrIR14E9I7tPz1s+rb6efcDyViTiL1eYotwpUrsR
A4XVAH8eAYPFyJYABEAu4Qy2t9PM/Q/rl7YZfoWdm01xKuHTCRSMMK4lO72gbznlMaFaB5n86oqL
BL4hFJL4DucN59sHVHjtZQ5bWSWIrU8KK5+izWGjfnbEM0XzEQqxE/8DH8rDMXjAY4ZW+8nGa6Kt
Q55xNzMHe58r7RzrSQghZFnYI4ePLhxaK4yNirrb3HHHjRPyplVVnNycQ25JzCMY8imDFVgcqbtx
t2tc/zsIq4LlVQ2lBwPvvx1ufgmGrT6uNYGQXj4BVs4wTMQyzyASM8R7yJ27bTE8NYW9aSnuBrVW
LgrbHy9XTvrZNUaekIuyhHFi/puCWTFX4bvufiG/Wfai4UYY+L69mkNjGTfoH7oL1g4FaGmygqrA
IbbhR36INq56KsLSR6F+yJr4/abgxU33l6K0UGguEr5Vc/yzi7J4n5/3SGbw7qaowyPBRdSSq0SM
u8ZKwgIx/5wECbjt8S4Tno6QrNwXWQvfTNqp/ux0EV9YpYkPwlI0epa1U4NwG35GKfkVSZLfZJfC
XkGgOeJ7ZvWFeL0SOTq7lRG9jE+EYwBI1sIcrf1xsVQXXoK06f5A8wrYYZmIA2Fsk4hHc76/Jyy6
iKhJoUVAtLGqZrvDT31vXv586/6knjokbiykrjDMHystcGG8GQksvjCqVhi2xLAS+okog1x5t9Xv
8FisZLYBnfrw0ZombwsNtOGuQKauZYhQPCBFqO+EHT+7Vj1Qabjv0f3OadN0Bxg1OjYZlqxNb9Lz
EYkkpRevVz0l2cnUJUojcuFU53G1jhHqNgXSz+0ebxMZvUtace7/4xDyBrI12GEQaLiEYfwIDa6y
qAPSf7V3UOF6z8fYK5VE1Jl0bJA6hrcZD3IgOXUeKW4FQ/bLYgQ4pWcrK5Jr1PbUbJgkmaom26+G
WlNbKBcmlhcuf5xzIVaQ0xs8GYAt3OLlvrFQ0zB+qHsdpUtwoAzgSrxKW36Tp+EpcJDPJR/ugFeN
Z0wj1PBZP9ngzLrrYazBm4TpaPyVVXTNqqJi84wlvQF4IOBrD90JEEKZmPO5vsH//iF/1yKaf/1N
0uho6ASNF9HI+8qRTgAyIpHXGzFENzs+40+j0Nz2aZ7LPIESh6LOdJQ+Pg1tFmK69Y6UxN2tg9EF
K/KnSPIJo9dmGhGn8BVMOscPC3hIRws7FF3mE6DTTMWUNmxwLy5FCTmq6FVmqqkXJQQRN3i3eWTT
ySttIipDVlE6bxgLaS2zptSsKvxrfOJKwOqaRf7dOLMhKj+xaUwnUTm4+SPpFZYoT3V9HHX/MuwT
voP2Uc7g07+ZmF0GkDmRGMZvreKSgYXeElvsT3RcgOhurgD/AifN1BwlZlg8S4qAIvOAGSQz66v7
znYWFZGuJ2dPjSlZzM72lXcJhecJs+1baax8q8wns30H/d31boaIcdx8eTLBy3+73p912DrPXjou
N0+1L9XaohrZaANH9UvvPmIUavq5K7frQaJ+NMx1Ph5pLkF/Ai4deIR2CPrlgO1EEfuoivEYF9kI
3YAkM2uSURxb6HyRJac0PnfL0yFa5s4uXhqNf/g3k0b/JQxvTiSFPKYQTdJLF+GLTotJRLGHf4rK
d3L9ybZe+9rwUA7lvHvk1LQB64rM6tR39DTfgE74HpyrTDUDbd8IMxf53/NRIRCNOXEoqnrLiQ6N
H/HI5T/lr3ctZbBuWs6hobcyROQMzGxDOwo/ci1FEXdgmH2hHEjcFfpbqFyR6PQ7VWqPgVZsZuic
7sJqpIufG+9nCr0uNxck0QwufZva/8Rko0/vNRuff0cYEkRifblQgegVdGycmoR0ts9UB7Djm40Q
17KpOBMNaEUc7F3/P82Uw7iniQ5H+Mp7+ah9Dzemko9GPMWczfLQWAooB4maxp7DL7+uve2q3drp
wSPSBteCqCdnfwvCNDc+xGWTcWHBrhqcT9UgIOoY9GPm3vKlzAmk5MHRipGPwS7ubf0Wcg6dlJw4
N8etJdrthO0y6m9v0MEB7vngYUiQjHNwnadDGEmmc+nDsoZ/1ltqmnbYSKh44mFjLHqVF9mouxoR
Q7ZDoBNW30s2HJ0RFTMVD7wl1PFBg8DfLfJXKRJXB8QqOWMuHg1MiXCAgkTIYkfb4QUSnevZy/j8
HigghklquO+NbhcfINdOuA0ZUbdMPRGdwIOo789XFjIZMw2ldd21WtKiHXs4nPwnmHTT4NwdT+RY
3bFdVtYDCGlTV49R6DUurbj0u4MFpoSVmzKRTQMlpCYyKavARRWPY38vmPlUGiBs/QBVtkzMeRri
APrxnC6kPmZizeSEeuGv9YFpA1VSgAMg95YPxrV0wUrDMjPMLuYni/jiSkvLG41IUHUHQk6Jhh48
N5fA9ZdZwjoCpMzNxm+v6Gi3BZi/rioSsmJEa9NwvnKkEShP4NDMvYkiVbtfselpYPzFKmtHWdOv
gAJfUzBbxHQbNlNV7y/3m5enkveZtr+WaoBCO2Wrbq1wgZYkZohtjn3+ja8yOu59JkbFj0W2pFEe
SC97IW6/5nIE0DCxhJAwA/R4OncxQNcL2vrsK6Ymz+hi4MgbL1QcixTG2jvdpcORRQsX0G0SG00X
cCU9UI3bSyDHw/Ww6gJcj4BmBubeSlwAu43noFGciFKU26codv1clEeuz5qNyfd9FjhjTW7ahWpN
NuZaT9JTDNpyoUDlcfXXQitzjYZXqEhONETkCvEllTuEkaY+3xaoKOFWVYzYb6BxiaXhQV5yHlCK
I3DO3jinGHLDTqEaV8BQ/F+DHQaNlQ9LZkX0bw3GycXsq0AScsFFkwJc8K2srFQQkWGmTXqLyxsS
IqEMDReKzEPAjcxJsARKXhM6o4KUaOWduK313UVCq3yrmovYPQoHy5tg2HrCwSiDfi2ADdFvU1Du
9lvT2aJm9by7VNSUkUCSD5EUzp8WKnguwTtL7O+xGc0rORTf6bPCKOEjnWEEi6/QowsidXmZwjvX
gkl4x73vh5REJSu9li3qcP5KLo19FjkQMCJm0as5aCA0CkpMGDXgNhdsbpLbFSfoFXH5Fys9tgAB
U5IkCk8NFHwP64Y3zSzWRWQkFQU2tgYYloOqv1kyeU5VJrIRy2yzOq9eTxhwxHXQ4VO5LwdkFMFb
lxHEv4Db9OTfrooCP9e4YzCUrDXnBm8bamiWjUz2Ap3oT/0ur/v736vPlmRbY7MTARSwCazHj1Q/
pl0Tq4/OSnKG64VVS0yORh/8WdjTsZyAFRSAPd/jFxjqkvBuIQ1oUJzut3OLeDBcJ6eBzpddhEdt
v6DqiGZirFF/UMo1FhySXGa/Gp2qJQV9xSA+5q6BPevcE7RrSOtAtdFLJE3zugKs3von5ourY/DE
vkhze1zneF5/Mumkzd87BWKcq5QjlKC9apnhK0pR3SFi0A7uQhcDj4deAgykdY8bzQ7yJfKIZB/w
9lDF4jtIwl7oVdnWZmUhtAAxyU2lg6T8MjaA7aKf6z8jp48E/zq/SYd42/HfzcSk5fnb5MQGbHcS
Bf1gu/4Q8NVLRrtdpDKjVG0vO2uXTlvQlS4kI6RZ3xhPEyQsNUb+s94VihnLcgqTiRz+JelrajE0
tfSNmy4ue6Ot5gorotcKnoOeXmQxYiwOGxh3uK5uTpvB1p0mgBMys+3S7KEiyKE0FC5B5AVK5vuH
HiUFk0guv76yVXWDLsFp51aMaskHG/2wYeFwwBDE9b9wdC2iVHN/boiQkRhwySsKuPQcSb1beU5x
Lhn6vziXZPbUQUgSsb9r5vF38FDiJAfL/27XsIdUBLj+PsFw3a4NA8I4lPjjuOULdIQIpz17WLLs
xfot+qU4crJXcEBFcVeY0sr5U446R6msX+x2iq4zG/WSOx5i11OJ+vZMBzdX9CwkdDIooNM337SL
JkucmL1cOo1i/nT47zYZsZwoWltioVS1SG0Xpwz0ZsF8JkwSYG+6f9aoVrNDchMO8p/2XbY9DIYU
UEHGRpAsIlhEXnodWnFAoHMZeYcezFiMhnvP13lmEhMt7p4cV+r5Wu9NBEiUdj7k5OSVKOGXEkdt
LFXUwKf2GnHsvK3qT5JjqexgVr0CrkDXjaZOymKMCs8MZiq4Z0oK++CtHXNpdyK6B53emb6jQWXW
Lco3H1Q+iC2YeIuLJw2VurUm5u1Ew3uwHvDhDyv7H3Z4XaNTEkJtN7ty1x/B6XxQpPuW0onRgmhS
ZJlXVxWZ7RlndPl4z03pDq+K7WifSTPhqsHAedT4QvJOZ/3SoyxdliA/uOq7EwEiBRtTUyvA6teV
7g/xSLTSAZp8pzoXj5U0PICULFKbDXYGDfEUO8fEa4mqEvgGom1lTkbW9AxW21iPaFFhay5iGn6e
hdc1PYnmxm7oOWklfJgDywr3RE7hHStw5/6Wc8lpJzRkRz+RLmoMHzLd25GRQBoQCoD/wNViymRV
ILHyg9d0KuSYzhNPUZDzRZTih03cFgzrUDO+lTKJN5H0sMJrIaHnaXGWg5xxPM+OMWlIGNe8iGEH
zjccWH0G5mliGjHpiCFmkxJwg35Q3YMrvOjz4kWT+rnMlbNo7WrUvzC8GgaVgAXW+8Umnh4gK9/P
MeYFrQhUGgqoOTdgrWgNkL5+QXim3t6ZkZwBriG38wSLhGaOwvk4xfi+nU1xPma8OHgImJ+Z3wQO
eUWaY/3xsn40gd3+LGBqiCTASjdDCw/hhOQNawlr+4rikx5e16eFhy7AKnq1Q7EP1RhFAiT8u6zN
bk7XVPxl3lCg6Ye/Gef3/rFmQWLAnl1kD3S9rqtY9MLboHwAJFb1sz/1+hGyl+tLBtWz7xwlv8Y/
PCkznImUZqulNgEoOkm5FlLpS1KP/C/OYuQ/Zmm8fBSpAmr74tMoVijfnJprWoCtigSWGXp8r0wS
a5qiehLgog6CQtG7MyQKhjslrNGc12cUw2EYgdlOY+SSalIgJMsqvgcGee/4dlkf4WVlNv3Ey30G
ILEnFBDYtlVvbznweNe49KuBHVj0cMxLySiYuogzbKfVCfb+U/y8Ki58kD1hPsixmIF3JPif0ral
G5xsb7QjHSJaPzhDAEcCvFfW0YGeJxuWiPGfyMC9uSr1IYXIOJ82TXtjujlreY3tnx9j4qxi++f6
pCdCSwq12zo5ueV8l4mioA8jb+O/XPFpuwFvysJR9YdyECtDA8ceII8P48A2MDlu2Z9pXlilo+z9
Tlioh/Sabq9RgbYH3desFajAVkK3m9YtqZ30ikdv4ZN0kScYjOB2/vQWkxT8QXPWTMLK9nCzxEhR
KFIg722aZNmPPh+5XBvsCjApCO+sRDC+/XCKdhYaEs4C4aFo26lTAZJcAzEzCnJp+aF5veUjkVgq
Y5yK//X4JQada/zO+6NFXPHs6zaOja0U5FvVqvtNX4iZmsSI8N2+uHZ5aQKVwQOq8qLH8jTtj3AT
LfH/+KL4PBDjefoNffaUXUt4W3xOuOUWtcQVH/H1enT2VOtoW+sVtt3o+zD84FEUfzvU47tlTq3O
Zq0pN/1CzOcv0WSCz2uuwPIEIo2BpaYJrfgYfuVK6SVk87fdBysMnmnNbfFFMf3dXoMo4AKFIkIm
FPizv2sW5UeOON/d6zT8cpzQj8XzJn+pNRIdxgoH/oJzuQTeM2hM52P+5e+VLtrERc2odknSxDk/
NKhrRR3A55gTd1g7Eq1B1Dn8EDRIcGDqnA9FsgpgpuluAvUQ0yJSu/k+DmVi89JgzH/UJFQi6MdQ
+gxTvVwBFsqFZKkVzo3DVTrc9KyvqR10MUqFkIGtEQ61f328pOBKQFVJoy/4EkUfBJwupfFi+UC/
YhpQCMr+TAspmn3hBFEh7NpyiuBbRdI09PWUDYobet4f76sKVXzOZwjH98Nlep7fIw51XdOEY9Q/
r/tm0IHKSSEOiCvx0RCjSpulgZyIT3Wke3KRi+6eDDAPa9Rrs6kVOV23TxALkQauR0DBFOCMsO2O
nGD3aLfhHzrkCJ/rYVUoDh31nK7RHR0qh3CR7CoYmVlp8T9gzFRPO29pWERmvKMmPWDp2FVVLrM2
JS5sVjx3jcNaOmVE9j8dBuc/m2usYMjIf8d9sLq2tszyzsDYdAPKSVQlKXGhxsg1QNDX/YtEkwGh
r+0k8Hf5CYgaQrAmCXj02zP8CKDnFmkW+nxnnQe10rNMjFollzoRD8sQjjjfnxFxed1ymp57Bybw
RHgcNLyxHGyA91je51a/aQRe6oVhuJigxbspPKxi3heK6TOiJhCrWnMNQBw9v2YT6tPVwHjawBVl
BFsSOCqBSv5VLJET4JZCY1pxTREd1b0RFiS9FXh8RjyaDugAq9Ovet53AfxeSv8Li9mDfN5sBGbX
pnRCbyGWXjQCEWxgpbA3oV4jtiW/Vg346kpTgsrbHikHJVG1KXRPrSTOruN1NpuvymVqj+ZdVaDf
EQBtkwJprl5AZfR3HlEWxbEjc6Hsecx+Yy94aFpebMnvDVzc3KQsvlpl2NOr6gw+phauCzpuyFfz
RL+YooM6TTcV5rv3BBFm0jjsG8EGOdoYGOMQWpBqozAjduDZD586s0jh7D74A2EguPPen89ObfMv
vMm9UVcgkKRKmoPYIrqCEtzVl4yY9ImHQuoVEHfU/ykSnFN11P1n7Y8KZ6Ij5ubUum7uAuoyZv4w
P5l4wYfyMrJpd6G2+PnqIVEn8lZA+pwxtIu2jsA0nWCnw3Ai0xDzIpAp+PXKQ0W/CzHGCmZg5+Yj
QNtG96k+sNcxtA1FNk2oQvFzM7FVx80WEqDGNLTODWqtA6GkdjjdyxoWAmgOYS0HiG3KfdlzAv2n
Toxy7ZPuk6+6x5c4GoJu880cYak5TbzaWrT4s7FFc4bhYYiAU/BQLvmfoQtVigSDbSaRk0VRrGUB
rPYJinD1Mir+fkN/W4yZD+oePvq8nMut4jWL7Sf0ownSVc1UzW60nlAkIPdEThpnrAwZsJObGr8W
DdkpGJNCBiPYpmXILiL7t6mWzhsBPRcU6BcFToeMFrLdExNbPDT4Y0ssdylUyK1RPJvPzjlmuFRH
zuWYAFmtMfsXR8ssEa3qyQHQB8OW5AVtFTK4wYZB8oJuws3XlLa+UE3tFjoL5O+JNBBonkrJkgck
UYXSgmeLysPXmlT+O1UtGSfI07ooghyEZcwiUCERdg/qDWY33zPhZOWXzTYRKDICByl6A1OvzCOh
XE2D7aWkdhHVmSlNwbhfqv/zwzlqe6E7GORvntyTELvOfSuGHlPmOHCUbw6T2Z88ATBaPT8Lt+q5
qE2TjI/HpqZ9wg5S8k4uhrzzFDKD92vuLGNYiMl3kpwfJSBAV5BQHjpKQt0/Y+Jwpw/2oMHzQ/kx
eeBGr23Kj7Oy+fNRIVbBaF8X6ttekU9Gb7ISf7oMt3tj6E8WQbQ9fwN6UtcSSRnmYrHhptNKQmyT
oY/XjmmZQcaZ/+03LMIpDlM8qhz+I3CfqQr/4qeQtGgjUdje0E/fvhs6q5/+SNJPZt9NGRPlGc9M
eAZ9bxHBijNbROY6LPZUFSjJRC1W0XWyum+8rTmug6BvRl7tdapA6tandJW04y3lOo7Ix4aubK1V
PwsHtw8P+LqLIsErP+tOkmKS7MmzLg2FnNNGR9W/YwQYW2Dk6kJqgX6GRqz/YneXxXoaQnbsGAW2
ZwkzY4vaQWhXxGf4TWX1tq9n8eGIGE4EpVkdS8DAs+dXIlviy822PgvQ2tAxkQv5n657+j1tfg3V
gRpHdlsWCGOn9oeU18m2bVwPj1MRoXGs7K2QrnIahW/3r1rysF/7fm6qVLTpZHGqw0zSEJVP7Ciu
5+5G1B6SvydiisRqej1HPagtwUk65l7v+8FfY9wuixBI0cDhVhxme5Vir1VCUH22O4W+rFtc58/h
RShadps2B2lPGfovnQnIfgM8OBvIZWp74Q3RXdua18gtlUIbXInjfD6zxJr9L5JdkUCm6//+MPdm
7ZKdCTWr1lNn4dzkswRq+/myCZ4gZfWvvcMojl2dcudUGnWS3I8qXe9hm6i5wEEhC7wKO3lNjrOv
Kx+LXhClrUfXvEtwqI9Y8qpz9gtuX7Cf5yc5GcGozd41kQc+pd3QCIcDlwiq3LuSVn82FFEAq5nz
oZUXxZggQlHf2zoXQcDLk8cwfF63h1/Ydy7B75bmuXwHPWo79Iqnpsj28BWo6Ux4r84Yyw51zqdE
Gjqo/7U90z8ojdAHaMWtieHyhms5N3MT9+4rzcfDjU9TyJNuT5bT/6BcJ7z9FUF2Yq2AfTupHmLb
F2+Cj3cZaZU+EetEoVTwPakFHmY7MEyrJX5aaZHKGPtW7x3XgRi4JGYnZHuKhn4RSD0/yrO4yEoj
qYSc3ThcuHuFeFsZOZNHvmkuRs++snAJ+TSwmvz5pQLRLovhD38T5KxkDbZ+L/yEuh7zoo5MOodi
HwhfJrnbdbFsQBDe2QC5Yq7F+2p8MdcBjZPA6fmngER1tnZ0Mh8ntkFmHO81wP3xNkkG5a5C+Ltf
oScuWa/zBZFZz4rD5YT7QbrBLGcX8Es4d5NNHjYLa6dYLeBRW4b8HreEn0Bn6eSmSNPCnyrUtesy
6GR8H43fk+LVH+btdSV7M256ZXPHJJnIsCE/HcW0pZwWvbr4QrvQsVqYlwGPqqOknAl/CcjvOZcx
MmvaNzyP/OXoDmY/6CpzBkV2PSW29qo+cFj89zhUg8Gtq1A0zLxmaJsx/Oj2K2vPRthERkXSi2iL
EzL+Zr8uAUzTjpDsP8jNkJDQ0pnfhzGY6b/mVdr8MNkNdHYLNvSbQSFkEK8XlHM8qRHJBgoX2BX+
K26V+MjOUVMQdhPOBArZfsr24tVFA5MJQ567JoWU+KQmFezwvMPdGmrWjq6vXqMxmaN59mI68aMD
UNI380zyi0wnxByeugHHD9iOFcVyVaHGKUw7pN7je60OPRAuuJDc2Yi666mCCnbvEvaNexZ3a2M8
3El6oXx8+/D27o7gVLH8/eD/nRVWrHdSAhW0xkX6LnF8j6rEmcZK+7sWOfQcxqmkoW/SfdnYUmQC
hvnEnLJ/mcoTEqm+LzXMBdhTD0SS9jEljy6TePTd/JI28dS/IQJ+hG7BxcsFYTweaX1m0JtMx+B4
9tpk+kPA2CDI0OiU56a3ykqrdN78po613ar68wPJT662fO4CUO1p46rTLO0ip8pvxXxDdr0K3TYj
Eaxo9hU3Y9HgBsIfBAEmAM/1Nw6usH11b5MOOP5u2WDyLxirbtCDtbRgbuSj60p4ksdpvOYuUkCF
OWInTIMzZQYoZy+e1Jhf/m/qrkKNX880ZowXg4RInvtT+jieHrhGJJl3iLgUYW2jkSJ76vO6GGKA
GTOtgkjZ/cTJ3WctRX6ngnyVvsxvzrQPmuUeKsLQuMItNjJZjW2iPPiEn2KyEeqc4qFQFHTvb0Hj
+gO9mpFMjIEzjD5mjaSXaKr28RhyXS7+KFGeN9TcgURt3XDnxEUOQBgvd8vVZGTfMPb7sB/T86hH
pJqHVafYlFtZZIHEx7uNOt9/sCLK5yszu2ENVtRhxb7thv0J9dHi+oDPK6Mp5kU6dPnFA3dlJM80
Zx1AxPNTm3jD+jiRbzsu+Uvc+j5ByNZjXOlndSzyZ8LUfdlB4bzGKGaamooP8wkqYz6o6PlkkJ3f
SEAthinzc4wH22mde+lAaiQrDkEUuxz6/SgFxCQjjb8M/zSp5GzxeQgzqT4yOwYs4OOw/lvcsuVU
VBGRYgB0Y3vKlAYa6Rp+YHzcsqnGHtEL2ykzm2xV8sjdSiwnW3w5XW2UHwbwGHOOUOM/GJ8QxAgE
zJUW6eHNyho9mLJQxq8/02CSO8duYdGIxoKQGsVvQud4+apN5zJ9FWPM0rrehARXHRtnCG0Xt61a
xpMby3T8ZW7nEY+hvWK3X3Bcq0iEDgq1ZwMkIUK9l4GXzWr/pLf3/5LXSRduUxzofCoyv83YtT0w
w6r4fAl/YabRVYOGpwinldLsqVIlzCOYyGx3MFwru6EEQkedfgJ8CpthjM1a7oRiD4sGiuX3lZr2
JgaqVEU8BVcsTg1wLY32zXsdr0A2hIJdXRH6AF8TJZ4xl7X/rR6tpf1n5IwpgB29XJwi694klhyF
8kauMfjeunAmjJHJAfb7FZn1Kch29fa/VG4GAgfINcXlYMgmaEh6tF7N31mUvqvY5HhWj5m9zFUx
zowKLQ4i6NZhx1U75D0CMpNcLcW+5hvThBBBsSP/fWpUT45nblKyM+I8qe6Q7rHKmXUNz9RJjCA3
Ha+adCCJPkeNMPLSi4VOaZdhuxaBtoG2yGy+GokR/GcF5yAYMCghp5gL25lE3FAMZatLVKJIQwiX
uf6uxewmK+U4P2hU1/eL5H7huDz7v15L2U/0l0elKa63pEw87rvsbAOEfY1/zVWAJEnIulsp1EJH
9pchGawLE2ipZzsiq73pa7fWkmZiPROQjdK7HUJ99sM5QliubkS01/f93XzAupwQghE69h8wHykD
FskSMgt40Pw1adVGxCwNTbA0PljjnmOcdtSXyltVLcNzkMDa3USSJbYuMY/02ozDkcA7UtqBd9/T
EmIQ80oaz+TFHJpcjEUsarlIOzaq70B8duOCFp3X8ViwRNUly8rSHpDRAZjPdQ5ZW+/dwJWwjR0s
jVhcb4UHEMvsztzwV2x2hQBYKaeXIJLgEiYBJLtdPuSZqe3zoNjcUlLbK3dNOb5ZOhJewN/LVx0C
uYXyBZiO5kIPsmlE4VWotmVnyyA6ADgNFptqubVNB1dfzylks+yTr0kRwKGaN1wFV0EvHYkY7k5o
tzf2MAg/dOG9ZgPTVW+cXb8EBf9OGXZZMuZcIQnJ4AzXdA6QTrmgbecsINCGgz4h1ZAmCMXSf0mK
kWLfoGydyb1JOeZrCqmecYJk2nRvtY6F9QmIXXSDGd2N5ezL8nmQpnqGp6pTh0kcRGloKt7hrIm0
wZRYtGC+QCQCiJCw+uMohf14B50UqiCdoYDAhzBhOhtGMrWvEyvT4f6rH6bnpBB35K2j6jbqcvtb
ajW6BBI8vaQW2BrNNC1oSruvuskXNMSqgOGxSUUF24bO1VCPP1TDFCPq2CGj2XfVkttgX6KTWhKC
7jzHXMZC7cj1C6/Nz96WD5l9INtczqcI5Pv7JgLqL85Evrwuvl/3QmtVQok+CqvCZXX5cSh+afTX
iBryiOsM/riefPh+jOqt3d1FyRC7XUCYI78BvsDmbcIUTCHLzi9M9/MQdgF6f3V1EHB0k4xJubqe
fraaeWem79yt8/Xn+2MX8TfIakWCWCJdy6wZCyPB4B6d+iS+Xn8B/cPGO2fwfSoqfVjIASWWD+fW
Tb/Z77TncbwH6wJHl7wgcBO2si3dlav/wjRi4SJzX+6ymlFUgBrpXIA8+o8crGv2MbR8cG10+OSy
DEoUCxaZl0AbxsV3y2RHwNlPGEzGlR7EWBsFSq0Y+dS5YVtvCAkS+1KMgWScnt6Gux5Skc08jJYz
mJTtm3PMQt+qZf0d1gHnX0DRtdsX/k92O904xuOCOJlxaXE8gE3uQ2bbhOFM6Gk0YRporaB06Pl5
cTx15NkVEmHr5j0g5G9ieAV6FoZub1ZrCiUPcnMdYg6XL0cf++du5DQZEi1AikfJyR7AhZu+ahz0
8eKMXxDnF3j/AzZ+rvdxldPygVzqn/hdSge+p8sqstCpkC9TReq8KwXNixoYR5poEIooMVHR3QsQ
NVhO9HFKzIwRYYcHUWn4BWBPJNrO6gQGI4CUtOiD9yFEzpa8cyfTDDyJicyvxTLoOzdPUTVXI8Xa
Lc2xyL4nEW6K9EZkXRi0sZMmxll2C3VtdCg/N65TX8eLF5aw7ChjmKAeVPfiXGpWWrq+AYL2Bcnv
j9mqSMeoZjGpPEBvTCBkK9+IOAB/Du4tKyvigKFTcnnTttF7YrRfDuS6W7TZX/5jGBnvSGCb7Fd5
lYWZsnB/pN4XniK41yZrI6eNvycVyR3GHJAvlwlHI7R+mL/IwkvgOLGV3kIfPs4LiW4RYyeWA6xU
t1EtlG+IErSFuLoFDu2RPmXXC9v6XMEHCopHV6uwoXfDXASh2fo9gr38q2CKBkkNxRqDP4G0loDU
REFrRiiiNiQIiAvcyVS/5l+XmOaLbaCvbEnZXa09FJ75oaXd0x1VLiyLUuszFU9q1IH1qicc1L9u
ij79RIX8P3DQ3hY4mOd/pcXT69L1Zk/2fZZgbxJ0UHz2jIH45Mh2MoAjPpb0hXFpYbJTp4nM7zJ1
zCdLQynrD5B5U91XZLXMYG74DsWkxeXa7+/vRr5yicmBVNV0sPSGir6FqDX5lxJ5POVp/iL+93ge
yuQTkQVEOBgep8foZrPzVLqfg5j1NduDEDtSTZVVmGwkJllcuzBzyirrEfYYGoa/5WT2EKP9myug
d+Fg1S7Xq+Y7ls3IS9aEiWpB9qjoTDy6QYlpw5IlbiMhrXV+Xmzh2ivNPTWZ2y3q6Wigox/cG844
GeFtng4clFXjDx9zkbUE7RC7+G54Md2qfPzWMVLxj0xjraO2M0lYLUkZT8Ek6C2soovd7dFxCORJ
/8y4a/r1zX2W/YqHhuLnvvVj6tON6AdRCoMp8off6wssiUPhnAw9EOFdfSDRp63m/Ko2zQDj9cvq
WJaTcNxjRQFG2LLCYR6694bpxolcLj7JmsI1emEp/BYB3Qs2HlZcnJVWV3lV7y3o+euXZEvM+l1O
9hfM0ljl5+z3o9B0aK59aJcUH1dOzUz+o0MGxLh9ZdWnyOIMNH4gYh1A3diTGoawLnB1a+WRmku9
tYuciBKohaC5nj0aSOzsYy6KZNsXuXhIwp0i4/fL7zCkkWpcVFDopZApRFc4a/WsxytA3faWT7R0
cAo7mfv4TyignuL6klv04IB+0Zrikesuo08tjJKkL9TVtCl9FdySaYxOIHesGjK9y1p8EkJrYBgf
U2cUPSJsrKnPIq38V2NrCwcVlIUeFGsjsUp+cFdORCBdXqCgdYM2OE/5nFVbvMk5TFvzMzyzmqxm
5r9nT70fWfHT6VcRTk3XozmkczB/oCI1SzxYqpKDdTYZMMNE3iQy1KGVdUoYTe+cme48pkYbGdB7
Atl/6vPpBXX5JVcXKjmhwczlL9Vk/9GVbmvSefYPBnZlpSJZDirE2c13geXjdkTeoaAX1TiFR9iP
B+RPtCa5AbqiRx6Kesf8xM24qg4PaFYb6rYLp1YkUlj3NYicNEUAAomrdatPQm25g2IpWZ7IeYOz
XaFfFYOkrDekJUZm9MZbg40XSEkyXnbfzr2o9v+cbIhrlTugnLOQD3zP+JOY2CoM2KCwVixZZ1ht
cenT/BnLF6poUl415iZB1fsNEDLDNt6U7AXh/maPHidBXIircVNQyWougpqLAnWoZp36LfgMohUh
7egBGVzdleMCaFgVVUnezuJc9CuhX1cxduXK656Qa9CMUCwEiCirO8bbR//2Y1OC2RsjNwJ3LRkj
oRay5Gj/CtLeaYPCefh62Td4KF6fhhYpHymKETBd3kg3WygdS3AyHZJo5K1zA1TpF67/iOKVGwu3
hHC2NYHwKJAW7bXpBzzpr3gzlG8g7dg2lzF1zxPWYVZVNNSiIWCYWzGey4u8IAhGeYCBAZPexHW3
LpoREVN4K4eun40AksVopjRSaMhyrPx4y31TfBJRMLppi+bk+E3T/wG8eQoB+RADL5ipO9fMVgGS
9PRzPFu0CgTiARYK6ncRFvmVmna5X/nUPih6sGQKdE21oJtPT8VkUSGGF2qGIOE4AxPCPQSU/3uo
jtA2vEolzn/oNBxfABzJoWc29tQhtL9jtRXwt/GZhCunEuKucOQoTm8HPaaac7qYj7XlIo07iQnu
/IphAvpgLfb7bRBFfHBMC+vTo+/jNW6MxBxfNTwL9eoCcGxovTJhD1WmgUlzrGNqWiwCQzTF89O0
Yk+mkB+DYPeIpmTrD9gR3YCq0R3zLsgysi0NPycbSAMuR2vTZ3Jho36/+Mw55kyRfrC+yHrDZcl+
59OKAeaexE/ZTgvtmByX6S4PKDBDwWYnkgYd5Fm3ti8yCpZEn5SZUtmH7ddOdZwtehDhEQTf9AZ0
aE8TJvXpJ0/rE5Gt+LMpGhWzvKyq489fklbsN89GlXTyppSPEYcN9TiX99UrtFv6DAXNlemRmoga
ILltCfCtrH22TlzSl5WPC5Su4xwUakPZD7cN0N/0ZFBokvxOjj55jSzzu/PLUlT1FlgSThKFFYzz
uJ54xNDiGj4ob2R6X7XG5FltpFp/kNAW8S+9F4R1ynJHUHd1jcGPJ9nrBB1dvl0nW1l4SQI6UzY6
d68HpeO5ztHXdiONepuJnyS2A71nnJUC3ObpJf1eB+th9sF5fMAAa94y9EexsJOkuSKMDCTL+b11
/00fTwp7eGzHqa8Wr4LGFfRgVkmgVMBN6fqfEom1LfzSX0c1eAXYlLVkJ2SdvzdwVcK2kB37IyNO
d/Aw0UjKiHWZE2cyS+KY+rGO+KtEV4j1XLsz/tHI9/m7Uh+zDHaK512h4XcHSMcHJHNsZoWAncI/
1n4wTOG5RM3XUCEOvxLJtkicZrxt6RGNqUNagCSFE2tXwmm5m52IqFMgrev9NFx+P0H4sVHBQsUz
4Cjb8yPbtrkTr0CXXoAUCJswX/0z3tZiK1xOcAHimDS6Y9015OwdDpDeUbtoVIVrS+J9oKl0utAK
9Gi1AGGO1gW4TAqLGAo3sNsO+2DuAxN9GqmJTVQKR9FS7vOgR7/Hk8worf6GkT7w9gQYspW4Zr7+
Os0Q8s5nRelb6a7Y3E2vuGPzJwKvX1SVkdhvER5a6MdJKHPN6J4wXJOS7m3+4WHvd/pyaIVV1R/L
7/IJJ2o8Ld2o4Ywgv3oBXBzexZRrBD31KdS3qGB2gfniUPliFGwZfkbs+znlm2toZ7/GWNZU0VKX
6zm8lVOePlCgXCDWKP66JVwqXQHKPdgAG1YjgDij9YSNjoz5t5V0dPWUZgHAwd/KxXm2yKFwPohQ
g7Z4us0xjmtg6HbRamfHDVHZjuUJgzZCl7hrThyU4WE7uG1SX5FyOUlHa/GFtHyTmYKVILKcj3H5
mhW/jVDI7KTw0owlyuOWg14nZXGdpzyATi91glpQk7sqKysy3yEPbaBwsJ5XG5N0j5HCV5JhxHE7
9J9exU33ONhvchus2brvFrpA9vvlJUMTAdxwJaq/yFOaQ5G3hEnKXlBkzbeO0SIyZwDloITMis7G
cCntNEhY7JTOCRpGXwVa6HuGqjkOn87cuZHm2xxWxAQvlwaETbaaRPM9nTcwctvxFdpTn5MR5pfX
+J0kjp6rvcHQwHBRX2hFkILTgHPMB0fxI54SLt+NanuLvxCTtj6Pc88kCoPoVh8MOXC/ndrJ6lND
dxmVWjnb6urioro7/ivazw8OpPXdbMJFQAW/5eebVhvM5DKsdH+cIwWgWZf6G9zzsaIZD3SNwXI8
xOA7fi7/jJjq89ShvpYHprrXuYTTkTdjkH/9EwvgYrQ0m9xfHGVcqgpzaZYSkHE1mApqo3kj0GaQ
NFyFWduRpStjgCVTmdq5LDIKN4jipK7ZngV6UNeYgetg2BqIkWYLXyv+CHxgj35Gt7CZYx0ZToNT
yfpanVnzQjz2Xx3sGd23eaypoK5mNwP2pVivzZ92FuTkkZzn74R5zwWiIzT7tkYdAs9mpuxG6YE4
CeWhCFhv85db8qGfbdfaffRf3U+YNkntprRAqUYlO1TmB1ZB3uIv4I5NJgBfDQt6i9yaJ4MRc4Bm
BLmiJSbppkx1LWStnka0Rb1DHq59QP7lAqTqmlTFwA1rgNljqNHcGOcbidJnzKZIBl9yUTpLvx1k
oNnT8i9+rZk+IyvV0KYvIVk2nokV0UpmtcASKQ3jjGENyywnDei6MyeaqtAgNRbnJ2lF5w+hpikj
fbSKt8fW9WGDSUKpFxoJu2b+wu5NgLCoSgCPedGDOXJmsOk3HWl6h2yOaPj28CH2FI7jXhLiMHOZ
3rpW7EH8ZHvICyKWLnWvHBPefkpu+Kq/iGZZoKEL9x8MFGLwue1Cgw/3CVxfTGpyevoSJQo/34OI
DfZS8vfVg5wGu6PfDahSyNHJGzyqhF4tefYNXHfI65ieljtfMV1YTAZ4DbKQGsDOeQqHxwcUL5w7
73jsHso/jF3D2FWNKyzhQ2Nk4h7LwOfmtl5Lh+4vjgWGBEItW2GgvIiwJqOu+6UxI2YhiczD5Xsc
Eb+OG20hxL8MjBkBE2cz8XfdUCGTOU7swLs5IeZeg2iLhDk06ci5HdScVYemf5gci1eX2IE54FAl
shRDeHw5t39qxOgf/HvMEvS547+Y9QpL/P+Xe45QCoUVmXNZG3287bWV/FaZCrh+cZM5LdQ+UkIJ
P4bMC/rGrPeOrLvEYBKKg15Bg/oIKcTMLSJY5UYVSNFU5lLyg+8OzY7oJJ9o+H4vGPQ6aGw39Hgh
tggYFCQd6XzlzCu6KwRjmiKf6sgbkKzLhKCutprZtRQks+JISTfBo1QidkiY2jJ8CU5KUIWSpifz
OF3Bd5LzE3nlroRLtuKAc9iST5ioZvGj+21UkAEqQ6uZwnodg83PT8OCLT6ebRI0JEuGYIfpswc6
1nWQOIKFJ+dHrS4nK0pxMW1U6q4ZBeFaCyip6jCfjABcbqqjICMixmn43tzTVB4lUZC7pnrCQi5n
8JrCfjM9OB3BccsAEVjCYJydklEqVl06KdRAblPwMi6PD49ssZWj4sGKqgay6ALioFFGn03Q7eb8
Ir85qsT9gzkaZORC96I2iDljV5WuvIz2KWs3/lkriieX7mcFWjJxQ08SO/O9vJzSL9HE0l/vo15j
ldy7HkeY/gyEK8fR6CRxVN+g2AYAv+WeI9iZEj5zp3/nqQn7YDS9AuJYoDf6lZB7S3815618Pfe0
O7d8YUhD0nCWYqwGXbhExRK4nmKIIBE2y+rdLUYAkpz/S6inDhgN0/AeeWjXz19IOBmY4iNKHBGs
HKTmQMJAqokkmPLWJv25c1tt5s42lHOquy8jTttlTIJXsfGREGH5qVzT6aVZknLb5KjHkKwTG/Hd
fJ8/IjSxo3WuhxmLXskDtUYskojIlTJuO3ZkOym+El2+krBi5B7X/kXcwwL54DNWhJLFwiE5kDIt
1tMqlFCbiXqqYPbFmHHtSk4IHEo8mdxt9P1J/WescMjlR4vVLV6ZSEfHN1dinTyOclLAxkS+OGdn
v5aXUf/nLvgg+M5BDNq8sZuz8JH8Lhi6QQByWGVdn9gQ64+GFarvYtDblR6+saUG3UOYwP6ZupqT
jmBFXGF8iHslT+avF8w8WL5NvjSYE9vbQJT/UDnuj2YvBeEVfuNoObzBSAMf4vIYD7nzGAlg208i
5sYt1MbR3A1rTTB+/0Gur0CFcSLwv9+NUGwpm2sa0IRdGard09Qo9E+ADXxwuA4m7DX3c8+Md9w7
GdvrpQ48Tr1b9P0+DEYwVCooCDLa7BMKAs6KQpJncz1IyJl9zq0vPxmudM+RNkSegSKCZrUKAeOo
usGV1H1JWp6itJyAOOt69s7qp5HzDAbqsOfjpCLOt8r/0n/dVSdakKxlR+kNKHKs7yfXP8e+mryj
ZwPQFYu9cn3Dal0CqHYh+GFMy7OdCYs8S4wIBERISbekArhpU/PklxN/9M/WZTluOQk/UaQBl6Nf
M8v62E1NdMx34jJh+mCwtDiUKD0dP6WPAltQ5iQ+CxZi/7606xPGsH+2AHIMRhmEG4gJoA1WcvTZ
TcN6HEWTwArkr7fnoZqrZe9DaquUbXUahObt1SWUM6u6BfTDOi3RYx4f709Nfdm//BWRtl4QQXvb
T4EqWApErl/6PWpe6nCJ7+/TXgamDFGzlKQKj73ymzKyvsZTPhp/LRNCOpXHMDpZkjb/qKAzXdJP
XNubsLHxLJFt0zXdZQy1A4OopM6xQ49mmbyuum6x1Wv/q/PNvdX+nK3dYilfG5vYqo3g4CnwFiMj
ucV1QOSCGhV2fxMoaCQh1rf3RBS8jMCxMk1i4xpSDAOsHQQvncK4qfw76ey0cL5FpayZvjwLe8SB
N9/D3ILyOvMZHxa+puJJps9FhCQAnty0vf7XZ+I6OTZQJf8PW/wosJzZtnDrzyAfruo0F85Vs+9i
NR2Y+f7fWngB2QjrZeVnlN1EjGypF9uw1lnB2rvd4tyFf30jByteSHwYJQCllmgER4NHNjgXNdEp
H1P2F2BaL7+7+Ud+b/4G5AatmpbY8hsJh+qlK2ckRZ/V03mUJqCPBWv3or1Ibl0YHeAAoh/dxb0C
tAWYOIwp+kkl7QUuSvYs9Ybe8ubelhaTS2jMOibJsUZSl7Yjv5uSj7oeox8tsNKOhinZH+xn+CD6
p0PCu12oEb8m6SxuU999lOu5k+50e7RJo6wARRUpcB3WF4aDFRgC66csIcVhfygGh1sNSi64oDIL
6tZSSpMW1PtMwhpN3K1Gs8cFmbgNy7/DvBYzCqpF0I2npmdBh56iH1sOqI6X+ezs8ENa0dPReViM
Vxyd329LEzxBKOWgKLX7ygWnMKbjP5C9VAuLxzN2dFehtRuA9pvaLVt/uOcd1ue1ZCZY0Fr/k5eK
cOJZ69uWQTt8ZtUlpUXgKTlD65kzXmKfM4nz4h2hMV8OBRVOfqIDZCXKI2VtgQ3t3RuVXJL0Nxd/
mXFnTUDpMctgJNVLWyxRcvnkeilHpiqVdSEP2qjNBAEtQKxgF2GfoefApcSQxqOeSivz3BtVyk5J
VGkquBMXoQBz0dkBRdXrrhmxEzxeO/Sr30G4V0JGByk4ci+WQsi8gDXHbQSv3Rg51uJzZBsaVzY8
eU9d1/AbtnSmIEbM68GGQa1HCBEDzDDb+I27TLqPsLySYIYKGTXxiYgtVdxquc2eKeZMv1dgxMyH
XZMW45lX4ECMfrsCfl3CmTHojo+acs7Yi0KdFuFts9R59B88b6AuSZEBKaT8ZDmuSaVWbLX5odFd
sf91Y2GngSafLXnpfOdwBhi3yBn3rm1xj1B1Hh7R4OnvBrcwvznzxlVt61SYpI79mMLSolwEvT5d
/3GksZ52GbRu6KhZpmWgZ2twdiskZAAjwjLTn2QbEFJby4HrsZfV+KjV1OJLrx/8aMPPz6d3d6Py
uPt1TTQRP2ZDrSTIHrOg0eCCkd6s9TXCnJPOvDsWSStd6gG5LhvF7yyYM5wKXwbsut2GY+kjoPqJ
PORBW83FeYyLZTorECIHlqsDTOq8uedlGJVJV+b3XPDSErJri9dDuc0161GO5bn4B4kvD+DCOAj+
09iAnEInoFlWvWVJYE64rPBBqvxggfWwnfeZD9t74QFyyE4S0uoPhBB/OKrbhy3y2PyiNfHhc57s
xHCFybkwzip7gk+TmpWn5lUBJfxeqFyCz6l0RkG6adbdhrh9EQX4eLi67qBIQ+o46ocJEUN6JAz4
jVHWo0PhVdSaXADCURjgA5DZue0JhY6jqJpoEem17fSo5nCS6CDLyzYrv+THJcsu6bKFqPhrC0EU
tfi2QcIpofz+rsZ7tl1nwX2Ak20PbnEMv4Hg1x8/mY0zmErk0ndDKOzubk82ch+cWcFq8A2ALaxJ
lnBTj2fjhhAlaXwNStgLSNJzMMaXN2ykEEKIvKWIxIlfNCMzvXXjSeNDivsjojtwvGC+o8BU46rz
xx9esI1FjnLqJe0Ys8wif4RGsQyzpRsH8Jlua3cPcI+gL4+eKTybL3GhE2/h67IH14yWgBfcRUnK
Jis94A57bEfGqAZBHYLPU1+npkClhayT52LPMTETDXbcA3p9suMlkJAuGuvPjYOycxiJK9h7OB6V
5pphRmkzCJE+xYzdbY1bVtlpCRGeMratciI5za7ZMXjllHhejK/JsZGPEWoMjDZ61iib/vxEQO9N
sFiKnAHFtCvTqbFI9k+j8CSCgpbq/2iE5qddKGs7TUoNnqx1qc6fH1D6ZbMbfkitxYlaMv8lx6Cv
YA3mYw3EHwiHX/QinygXMg0g1JqFM/vxKPILrXpYqU3RO3DqrnYM9NiBue79joTXmay1L3896B8r
6GE0o2jhyCy/sMnQ0anVEZy8lfFk3kUIlY+8IzYgykQ0S4g6zofu9rkOpGMzEpZv9KqlBHmi0Yuq
N5VteDVHa/k5m5OT6NXXB6PjTGqtSer7g3O8nctk2aFjIm6RSN2XJPCqBOLVt9t3rRP1TaV1HPLJ
bXWrhYATB4mm1uSXAisBKAUYyfLugm67Y4q+Fq+lU4zfgLo12Zl9wFEIUOOFo9RF/C8Nh5OzMkYZ
qUOwKRud9cOLF+COH9LNgcd4hU65r9MSwCI/mnp/m3vjSQIIwjqCJN+ukMn0LODE99N827iZoIE4
ibnsrHSi3eEa/nMDjVzqbONYx85YBmI8jDat+TMuzU4rhf0STC6fhO73JJXPPXQUP1HXuSxOH8NK
1fd+3Poqans4EOMZq17m1KZYTmRyJsG2/JS1/kuW7rD4G1fy1bzXzRJUdGuhTHfEUyudLqJ8V6fC
9z/u8W7rCCAySQEnkDW3jizn08A866ya1Qj+BKZ26xTK29TMHpQz4E76uu0lEfA6DjDxFVvoa9KM
HAVCRBQdZByLcYO42Ezq0q2PrOIiDGk2yot77aP+XB4Ci5RG+XIai36uNrdnQSlLR+I8SMQ8+oaj
KcVuZxmj7f9pWYXtU5bQ/SOvVF7hWf120gLwDgmS/t/FrpbX44xNK6gUtoZZdRWjQMiXgulXEvBl
eCUoZNz2vfuFEIy6Z24S4c57h9GNxCSfqXEbV6+/wfUqZBg60rK7qgorU6rqyVNvBxqWn6GWJOwS
mF4A9IZIQ7+4z9IfN4R/6BdaJ4OF5eQG4PoG8cRj0vDbie4jQVZlAtw7XDhdtcVJ8zUtYqQ6rI6t
JJ6SwlDbJ9xvepbwyrToChnYcVUIgaejFZfq+uPFXk/eGf0C5GZK1lo+6FJR0uhqTovxb1U2+HYq
0AtPxzPoRsyaAa172ls909dpbr4PnrbD1HWDYuvuT2r5KvP0Z0PRhMBaPmEr2bVBseFipVNfVfaz
LPJQCWF/b4TQiAQHfrOW5un79/pGWWq9igD80rcnxju6fCN5r2frvk6DCD+W8RZGyeavw+tzt6i6
ZJnngr74rpO4vchtp4BOQ4QF1emFKhKkxQLXJvVtYEifukqgWFZkjCjzUoZmOTRcYAYfFyOJ95K4
aimM9FX5r/9fR5vjtkkkrOy1FEh97VRL8Ct7gOnnXu/awes4LlPfgcxxBhNV2zpp1RdKiFVTvy02
0GWW951pMPI2j258VKmJYPfbvXN1jsMqOXskHlbz2aa4AOt4XPI5UWOpTqFPA+X0OJkGN9ce4bvF
C+uKixWboGoSg2+tjdNM1dFbasArdi3yoeP86dRDCisHOSzbBGf1ZT8o4N62PGpS7tKbUpesLWAN
MrGnxuCaUhaW/TGHZPUjmQ/0FrLBOBXYlNU5bpe8utg/zv/a8Gus4hhcBZktTd9IcqqkcZT+x2Fg
sk1utoU59gxlXHIXd8UZfjUrqx6X36OSOF65Zc0UlvCRIMtstLplh/OSbRQiO0vcy+q8C7ZMN0CI
VEWILOlbvfZwrR5yxsUj/6kmJ2I3vvMpZ82f5iN12ZrB5bhNH9PtjisvRxpz1JazSZPSJ1arAcn1
qkYl+c+IXWPdAHlTV3W/SoyeJrr84Nz/9t2Je6OQUrQvqZj/PZ4YLHgKCLPbB6clXZMZFyhA5Kv2
j7euGrIhPNTiEKlelMD3I0AoqYsYLD9kbMzaqWcL7ZxNtZRsQDHB+2KwcmcnWZy1eSc+cZ6Eq7hK
/aV1jkCjLNK5QMxnDZJU2Ei2OzMvBT14x5mUzs/NAwRPVcJJlKiovvP0v4i2ALLq2rpT5++9PYPK
/TZaQNBVvwI+f804WGrf2IyGRR63ZJMFI6mJOSB3hrzHiZ0cjoypy0tDJsyV9FRLUa5ZHoqf7GB+
aGlaB1CEWyslSNdGFYXII03z81DXgYKeRGn5lPA/LD+OL3VE5GdFTxuC/nGU4VXwpbaip1j4PtR5
JjQ0bq7VCAN8NN6F3bvOf6qTZALaY5r2GylG4YcNWZV7TGYCBrY7JTZjGeTeZL02hjG5h5t1bNxe
WaLr03d1mKfrIr/Uw8vbLuAnwBJSO0DasS6Dqio0WJRRkDe/DWqfWHENOC/DwksHkIjQyv8YskXC
tRDXaXVLAgUkWUZSOjntsg1LnWJggJDw/TtYG3EOpyzQ+z0+Nq2LzjfK/bzN4//s77zWy0heI5Jf
MlSHrGwmqzCNuYnw3+riIbnOcl/K7+F9oVpbfgxB4VaNF/Fdu71jz131Svyly9akO9hEfsDVwH3N
O+6Wq+/HwYd/DWa7hiWrnIktu5ozI9iP3Jr/im4JyhfKPtJgkbVJB/9Vm0FiL3vPtmERj1sUDCrE
q3FgqllcI+Jzk0usp462h4Of9MweF+VfNRtm2uafjQB0NUsO9eEr2YT/U62U27cWhRnnGQX3Lx2F
nlAPgk4GeEtq6U1FH1+5JbREC2UW5ivmlyamJ0aPg2RVlizF9zRMLLCGdm9F/B87DmosNzXHdgrv
fEyeZUm9vHGHJ9fo1Knq1KEjPp3YGUI3O/HfcTWJKAtuaAm2ZzpkxBLLmBGmMAROXl1cufP8vDC7
KIMHCfVCkOy51Esieh2qrulfQswIVXOQnzUPOBey48pLjypCIEgY66orxjsDnMf+eX2+71knLTAm
CLbHkXEnFETGc3pmI3rUYP1FO6coX2XGfTvP8kpev7jhLzzKHs7e76N7VSL2piv6zHxpYpBt+5Ez
6BkS1/+nDiffvPAi4xV2cPPCDunaNjTpQ3TBdz+j/N0aDUD/kcu3tgwa5mr28TeoPDx6PFTF1K8J
EbC23vk9Su5LqPQ2RreW/2R4+SoQXcSB8Eviw2Up41NouO+SxrZjCyU89ZsTRFQgKoZXLHMubvmj
9DHWlHF12fvKFyiMHJJljHmsXdYtPgIXpEDy4qOsIk3K5WEE2lEfw4gZfASlbG3Hr3lzyBHmVPa+
51FwfH468P6J/fEwjqcLSXQhpEmO+lVawaKIhTyebyA2ViNJlWUD9nzA5PdPjUpsj7+7Pw6P1wpb
bOAZR+RkOQqMAB+oEztprr6BcSh521KLPeVnamtzdQWCfB/9GXuItmW9SMLrmEHDcfW02ZJFaGzq
ulpp0yEcSGad+UJBqeDQjeLsg21orfz5tx6zsXbkG6T0iEl/n4dllRjipfzut35rtBrwG4Oew9rY
VP2fc4XdN7C3ECilz9surWQySKDtDMItFZL2h543bEhvudxs8Ls0GGn65hS1s4N6YP6VqRuVkDtA
kr9TLLWqbrti4wuHI4qTKrVdcWK/7ebrDDQIn3mrkG5RSG7DHyvbCmElGd2qPMAWDUWSB6mCvh26
DUiaKXNp9U9HrKYifqas/D94UIk2Yy/RlQoLYUy315MBySPDrjN28fGtEo2WObxOBhUS09dgeGrl
OPwJ2XKJRR2TWJ/6IT6UlZJS5K90twWdehBfokZFHSqIDwJLHrCCojlP20sWeZJKhn9WklE/DLuj
UPCxa9GYBrymOZu5istxm3LYIgaxFYila94p+cJKN+IFY7aO9fAAJJwMBOJfPO94JNi7MUiBk8Pj
MpwKJjuNNKWEckXI4LdDDfw5Fc2Xw/WawDh93sY460f2/n+WfhmuCgxOykSjR/cRTS3q0UXGI7T9
91bU9QIRAEttrkhp7p/5IzJMNMy3uIdpVNkHtiX0+c9J9nj0d9IE48amaZbpzxCHlEGJiovun6Dr
9i8HnLtR8Cvh8hJmXKgdcAOm20z/d9fFB04xlu5gg8F/Ip45q3S2WoH7gICAvSgn4RiY/LHgXtGj
VjeLr6Um3PRtJZrus898woluvafk8GnD6lEQPLuYbX962cZi1vrfXADPXC0sn4P3gkB5++dZkgP2
muIcejWB6+2QdvII7qZZ18RmtDqqjszmBZ6t4OgcILz3Od4W8r2bFgVEsPZhcrTY/lrR46ALCbgg
oPuxOrKYcUC2ZPW/BHqIJr0wpzXcVujdLdD5WRzpug8WhUxEzxaNGq6aofdw5/jP7k2GdU3asxya
y4HUtJWvx5LvprrbpjQhsW3cWrxX3rKq4IZNnCBgpF6bUOJVW4MVs1vKzR9Z/nCXWSfgCyGclyl9
6zu/GH+Qodp5Mow+UzWVuiKlA01MMWnjl2jiBBO73JQOwnUJfWRsf4KRDb/Kgg0sDScBI88NPDF+
dDItgKm1Wne1GPRkqA0dqnqriBgBnNjzfyZMuJAPOtlncErRdBu2s7fHb/PPR/7/X1W0wlAnaAcA
20vRvfACTZt+QJRjOGIFt3uz/N+yiMt/vN2qJxsBG0EXeKZB3WrFImCFswqpnaimjKErU5pA4LiV
tFwz/EabRy0GhkeWUIR0QGJRJz4WQCizZwr5RzjuUFQg003iKIRksUjV7fjL18Abqgsn7MAOjKcJ
EfKtFrcIeM284J/tKSK5CWNQUHHun2f09+OxCezbc7+fDJKoLsqhS4sDVM/P7qJS1KbshgSud33i
S5o7kqorV/DYPzAhr5UUF9DWRJxXZAKHf8zOgkfPA+oeq2Cd17fcIDdFsN5C7LKqBqwGVQYDztKc
fzfZ0y5QVe0rFi0DyeX1ncZrJK509JF68InFUKkCsDPGif2L1EwHWDxaP5k7K8chRCQ+KjjpHmNz
UPUM/GfoQ8NL1moz1RqN4LC2xGY/6Nv7L0+05WnyQp4z54roY5kMx4NC7bJZRAbOx1Y9H9PmXdj+
V0OqnFV6uLPJms//Giy7no5R/rOtAKbaLOCQkn/1EIQzTRnXcPVwNkqwBE9W2xJ6N89PqjomjWHV
MhnTp8xxn7n6h/b94YxlZ8ezvNxejNSKSwZ66e27EZrPruEhDkyZ5j8WSYft+KvoV9OVIlH7u1R9
rPHgrBMYKPZgDcGn7Rycz5j7j7VJf4Ofy1vvQ+De2RxfxrUVh3/Q5Yqv27swC9Y9hCf8+ZmrpeYB
198C+MhuIinPHEUcJHTneHSixPY3ZJngiAmdKklfxa1mV7ic7nsKRJ+ZuZFlYd4yvR/BbtwHjVkp
sc9NEFX5MzzmGsPeuhdT6wFu82MT16N4AlXaPxGOClmv66UxKemM8bPfqoqh0G34AiAKnALomKzM
D1odlbqrMCKGzreaTak9XqZ5/BgGWh0ivEz+Yxf4qrHNsnTMD/FYwFN7bM+d9mdOoyh5DC7D3oRM
Bqj7DL3DX1556QidEJkywWfkLrd4n4TB8xXuK8tOWuqPPIHjeG3587BuG7+r97MCCy8oToUqDdEz
MT3rhPB4RSYnjMA3AXwGC2Z99Ix5+ud6qZJB2Iz4lvJum15Yx0KeYjSln7e3dn7NDdWiKnr3HGTK
5V7LGoKW59S96aPCiiEuwUVSReQGUdPIpQ2Jhh72AWi5uK83VyNg7i4+O2izF78CuADZEUn7he/G
GVbm/iHmf//1JWX2P/xgIHLeHBlCinea031FkqgIBlb9kG+mGFa+yO4YfSz4rLsw7B5Ari2khDYw
2EZW+48pIyljuNrKLJNuTzrSyNNHXG49Jj/SgomMiQwFkJNQZbPMZYDlkkVBGKUkq+dUQvNJQSbz
SmmB5Kr3+YrOvr0YVIkIsCINcJ16t4igxrUxVg9QADzfW6VO1x82uPbLfYGb65VA2p19B55woVNJ
suHFdRkIxHgM2rbIms4VvKTXXVHxBSA22sce9LSKe4aAaUienk7L3d9ryTbPxHSuoZA6Gy2Pm2Bn
5U0kKcVJAy5LSvH2LbrbCyIFJAB+nCrSOZXL7BBp1FioOxT9ifLB/SGOaeJfZ7gTHN+7Y16Tke5S
8RQe/AQu853B/l+hvJFOkToZfTBXZUJEiiozJQVWh7B12mQNvpsXhD17Bdxq3LnyQBn9WWvoAF9i
z7qdWgJyl4M+ZIGuf7QznSNEBQxs2ZC2Gq8a+RBHc5lpU5OvcK0NvJS+61rxW+B2WnD2v/hGCX8u
ENZ5jfstMi2PhhP8XEuZXU5xIBARGY+usnS+/eERXoO1bWqt7y2pios4K6G3LZG2wKWIXhWExxmw
fahpeGC5AyQo5aUCxqhPImmsJzM+RzFRmVVaz61CGiio1jyBOq2fmDdarZWPkwcQuv05T6PfXO9K
ErDUCXL9eYbAu8WqVpcvYIBHa3lfp1e6w0NmtVwsTsR97qe8A5NWdeLtFSW1T5lhoJj0HVt+ebya
lcN+ibvbtoCI6yF4SVFvHGCRFMhLrD3f7ajGIhQ42Kzh9iOVhuxwtH95EyAY7pfoWVZLKxDmhwKv
3pzAjQ9JCQP3U60a6EhvUf4R27/g1CqMp0WYPoPx+OjdycuPTbW7CrlqeRKNm+wLqFoBQHfcBpcG
BSj6AXGqFkon0ninSQn6lUSEIarLDPHu4Pzq0qiSbBEfrjsjNB1lzhzLilguFeyNiqF+7PqxrwFL
xFuhbynQD+/uDjDqguiR/r0dqte2i3SC2IMU7R1NKv672ZwIPsC1agyZunW8jIv09UeeVuhnglrL
yFCnbHcc5ZSV+JYax7R5pJGV0MAyNgFApE8RAvhmZl0OABQmpyDdQalLm3ZoFLAV5WVXH5ERhMUf
MqzbgsYoCk8ueq9Gjn1iqlF/aydNdftEe2/ePkX6sTQ698VHT2erd5jYrD2Muh6IdwP8rtnRZ8oK
aN9ysjrzoFwnhfxaRfD9z8X5oClfaACo4mIhPHkXbF6Sd+X7JVjBnq4+hfP1momjTqssXlN7cDZF
/2W6dx6gTheraTa9cpgpmLOaUH8Niql8q4SNviTE4kFS+5mMXCIDzAWOTVhAMQZ5uPshgt04jbQi
RfpoWB5o0svv3WVHC8gZ1Uke0JGw0iexAnQ4RjubxiHp3bx3X+7haWEQa1n35WZ2929ZurnIbKhu
3NRMkPl6+wUSEJLFJzn1sLNHJk2sHaFf3WjDY5q62c4GIT7CY/bumF+CKoMXQyMaaxwVcKCd995C
YN5oiNNoKhIIQKaHPBiS5iZ0R9VCJHX4N7AZ+jJwv34VDrgGUeh+WhkZxtQhDPVtA5Hca8lf0CVo
hsrI0QJrqvm0R1ncMUinfwP+MNqLGiPP0eudYMX3zamh+8crnofZQvp4AVV5lXTXZLcr1wlipgYP
PSPb2Dmp/6HbuPStidQbjRksmiXkbC3khsnEPnw/tufxcpckaG7JHP5kXChq9pJ8TfIbWzGSbAt7
RnmpZXHtm2OLPMM3eh93E7UI2S2MniQEm0idbG+9wMQ3d4+dvTFjN9z9wrTENPCQEZMUiou4cLWb
JG6oDcJn/8hY5U12ITMw94Bp6IBVoqwgZJBEdAD/EBvm0isu6gKQZOdq3vIEfSgMqO+tt9YQuTrZ
x+IZUSVs5n6KrEl5eg0rmKFxxwxB/wPaF0ln6LmkQtXs7QnQJeeYD3n1QQP13ove1CjrHQGCo5YN
wfefKasQQkY17ioatwN8z02U1RUQG7gB2Lq0aUWUVkbmPVF/Xh9zkUrehyNWKzxTvmm8Ner6upuW
C4h3uxpXwo0G1YjG5qFtSiyJ9KeUeDoiYu+hcmEZw2iYtVb0uCiC/AjrwLPbT+7QlFZHbnAsF8uT
y8ohrHGkmKabQPvLFfg6dvB7CnvbgU4J+TciJvkwtr1m+OAJpoZqLphIHu46IgCO+eAF6Zd7PVmF
G0bo6xZU0SNUvvZjLVpcBUTwYLfd8tUKvbtT5mY/1+cgjOB5SqXEvHWM87On+tOkVl1VPdwDE5lS
6CME8dA4H2dUCpYBDyX1AB4HnZyIhE+NWXJQmCsJvqrFovqgUgVERFBGtJTRUxZbwvGZluEpTDZf
gy68Z/BMgSGyOi690068WdXrWJHBuYLTovhxniU1pUUZRm1EKIVRPmmbW2PQfV0ZmYaWvpCC92/7
sUbRfvnn6Msf+PBbwinflDpnxeqAwFX8tNmEBlqnb7QWYOd8VY51+OFVl+oDxaO2XZTZxWBswwJx
tlDwTM8TyJhOnGXLNCBnSSkvgilMYbKFverm8m/2A0kdOGBsVqcj1VSfqYM2p0x/WOTSkW40pv1Y
XqOwpv1YC4aeyehf3DsB7TTyaRPfRkuBaS3EoVbP+wr8Q+uWGSPQVXskPV0QfWachqPd1CfGI2nM
w5FkY6P6YroM2qdeKkKHCmZRbybtIeN/LMlxIwZejFEF3fNN809kALw6TQ2B9M4YHaKNFoy8BZlS
AwLbCXE6cQEpUcq54ZRaWINItti9g1yHYt/phy3irbkDEwUqsyf6Vburxa30wFVxvTcH8gu028MM
gcJ0CUjkZ0q7wh9ntlRWelCufjFEx+YK2Ydyo8xDpXe80cwcuaJZKYo0UuU3+cRXzzjlvw9kpSwb
nWCh+XykWyR/0egrvmBPG7BeckPh/lT7nMm+eRQDPnG4Vl2zjAL+Yjua9ICqPeh+JwkZN3h1ShZ6
/72AmhSw45A2qAkaJKhpFz8VW2hGz4vY262JJ/RotSlSiIxiAHCVSwU1mwQ12ZaR0U3MavXAaTI8
ZKoS1VyQwIxoHRa+jn5eFwlu1/yA7qTO02aPW3T9LsMf18Ge1/NgjRAiKmbFS6s+lwFuS7HJZFXK
SUOqNgfdyyEVZ/WCGSMlSLUUO4Hd7jJWiKbWJ0WPxvoRVyPpmRQMfp7P3nLIjJzSRcblZ0E/eGiJ
5RWey1nLHtb6qvzrfi50LEAkDuOiAtug41A4/B2JO0sW7iIl+8vLgkik9DxdItjKUGmT6iRC6sHf
qCL4481dKR1rjC6fM/l821gvzkBrx8gDC9aA6SScFwhAmjV8MnWGlSiR+O1k5xBAIQyoS2n+nBv3
AdAUGzlGG3HjNiYalACWnLhu07mkccTZLS1/W6bWPpczUka9V3pJhw6P501/DOPa6LNeBQfqJ6/1
40oDCmGLPfkObB97Xgfyy9gs7S9o5FCS99/soeRiLFfAAcox1gz5Y+qhdICRMqpCN1aOUT0+ekLg
pBtabhSdeFWRavKnH1a73pYCTyXUCYdKeO21C1484JofsWUPpbXP3FpPXgplo9ywPTddD7Epb54o
8VCWAkyVctBD12HxfftxJXjyO6/dDDN4H5tZxCBUKYV/Z8pLZB0+S1VP+yq8bQGmSSLYyDxGrm52
72/sJQghGoC/EgA2+1dfWUjhi6k1DpnyDh2raBcQjXmeJaiClOqQpIAoAzVPW9QjP7UCj2AQnurM
gg5uMQ8KfeGTw+HWBGhaq9FEpfwCmUenXhOXZ50Oc0JLw7hfjqpcUT6YsNmlo4oMvJOKcwt0SLAl
aIcIXnbS5CM58qLM7ZbW5YsnpsN/xrcU6E4jYClUQxRgQWFr3hAj+Mhd9I5cATETcijT3xt0w9bZ
GpezZVgbd4MPd6M8HGRp524AJq1t78/FAOuNpJww3jUMWVZM1OmQqI0Sd4zt2bCticKVnXPEKb2K
MGrnoYym0CuJAZw8BtgrJTqrxpiMzTplPFrXYkOQ+OTRVXEKkizmPe/zeH6pFBrfBWD9IISGWYzt
vJooWUiieQbMKT78tB83rzOAMbSckbTcIch/qDe6Bd70j6y2Ulhl0cDbbU97aRzxJ5tOBfSjFO4+
m1ZhP34MMKsgjA7anxStyTKsGOOV7rp36HqvvAWHbgSd4Oa1CxrSokz+UC35QkP68DPho4soAqEg
7XtVnOY7zaxr/XYdtZ91KejJ72saoQwbirv11LuDpmxlc2GDs09+KlJ2AG7rqZz0dzZo9T9ZpCtE
yLZ7T1UtCTrtTTuDWRSCgS00jOvkKVUzgmWllbd6MWVewud8jmpn7uQE8RsG9FwuWJBtwYAVz1HL
QbNtYGH3qz8XyG4J2mp6HZLz46zz2jKagcfzq5kzIPIyfno2nvd3iom7bigtrAwrObPtTvw054mA
B53eW6kuHkvAWyOBC7bxa/roLw66xyJMf0R0JhnY3+I1v9Px/xcN81mQWrkXf9TGbcBIWpnWhjzH
kfzKNZXI9VTocuBc02Agyp9IqqxLxr8TGpV4JXHEvdY+Zt4OOyHE/x3clHzBhpxLjtL/TN+ekyAD
ObppwqifZk05AnFIweLcVMMeZ0N47/xCaHDg/DhYnDqkDm/YiLtQeIc44ap0mVtk0AIffWMI32Mx
+AE52exqOMg1bSEd4o7qKf5WUnJ05ZI5Scf8ZGUY3PotIqKWp3wQ/uxsehv60ehORNFMwATXZ1fx
sjMVzslCFJYZbMyKkErO3aPnIkKVwYsx+vUoct31Huf5LRrWHJgmoDU8iEa/Bh+irUirO8mGL+5N
OxQhnfwZB2LdrZ9QoXrM9l+m5RLz/NNyXCqZx+rKpcsJiNU9ip6rj9q61aEeWymGVRI9/mxZ/Q8K
St55PAUVYvC9+l8iNe17l2XffxSM9DDe39vbH3Z2L0zCefWP+WkK/24DctIN1an9MS5W4vBkG0x7
Va0mQwEqlseF+vV9wdn4TujawCEVOrKaFhu+jCeLJDgw5snSGfug89lz8g0DEGpXtc155DJU4xCi
sXXtIYRycgijJtUuhHlld6lKWH1nIXIfhwu61LYQhAqwsh5tC6S2HCnFbLSsv/0OC5visKn9YYRW
DNDOwemnekQAA7LbgAu9XfLImgSBhTlvG3Ng5aJOm/Yrdut4+nRvAoo4439saGqokvDPj0NbQrsZ
unZo0aWMTTkaAwg/WXSgrMaJB9UyG1RVKeAJ3AytFYBaIfbsfFja8dv+wC83vOpZjup7AxUCUGKC
CcKFOoogrnA4+tNVwUe368nGxxLqfshqI5fcA1tLYUk0sx6QbSSD/+B1u71olJ45Q4WxrSpLjeOk
RH5P0EScg9iVowO5i0xWmXNF2mecx6O60Ong5Jdl98LThhiINodYU+GruXexLzia/N40NhEEKioE
jHRlRvp8FIoHzVuvqyaDSKTHCBi82lDGak//6h44Hdwdcx99PUZAMRH4F6DBdWnDnsyywLaR+Y3b
kZU36x305WzA4aKVYRyn7uwdeXPcv9wvrpXQnEMDXNKcskBAqX33VPDi1eW5A4RRj7Jbptbh5kw4
33vSSngmrSqGVZCvEuuWuCD2ZQ42maY4pFOo/HjQaJGpn1nK6Vp53/p6nZwRq3a/6q6G6K/b7irJ
F2+hN8O8KWnJwntaaniN494gVNv+NzZYcTlxobxQolpHxKZup5pw1kjYPKmrn5vTTFQ9oTO0QFLZ
0UHzjSfFgUBFJbCBmT0cbmjhrciIINdK0KIsyq/kcjyiMXdftY1RM48qvnrg1XUl/x7y3cfgLWu6
ThgKcbEMMBM4nZEkeFxAKutwzcP7bc2ZX4fc81+G0isBN4Cy/C9MIj4al3Aj0gDlc6JJ+4xz/zS5
01Yk7Tm6Ppl7FFENQgIwxcYa4KlYk4vPK5DyFjDQfeqj1kJu8SiN8BO5Puvp1TiVfJJWWlNfF5fd
02Gf66skQZUBGhazwByK92pk4kH+X92KAsz/EgKyoitTh1R3RM3NYjxkd+IvIOd/Cwn++BXY1lrW
uyl7+sc+qyNphMdtueFoBxbn00IxhBYQDIG2Q2ImuvME2BvNogo2XQeQdCKirbUrvSMPqV0BI5fA
XwYeLf9fhV2agkDSXIlSeEwi6egfD0yxuuCXSWHaDxHNaG6PABdUmweu2x9UzGT5kDLir1p9ofKD
baTx5MxnFPNDJGIpLo39+PZ5OFkSmHFAYs2cpxu7OvMaXjaGT5fO86kUh/m/GNBo2J4B+jRWg7b3
ksj6AVW8HqOLSh07wSCRxXtWOuU7stiLiqzCdStEpPnDQz4rukctVXLJvTfQpyYZ9G8Mrvilzie1
Nr4+MunXPbZToI2TTe45gMTYsyL6SwpvJ6d/KFhNHm+QVjTNvPX63YrZHY+qo9hm6ch/sJX4SG3p
ImR5dneyrldawjj+Cc+lr1idPCB8rvwK3AK5DqoEUZu2MFtMywQgGw6DKHp4mmoVysiIYNlZS15J
jzXzK+E8Rzz5IY+Dn7AOJEwk5yy7JiVJ9tpQLWn1q7OapdQLHokalAnws1vbOrclj8/mpFcOeJH9
43Sr8lBm8pPoeok5au/oHr/u6xJJZwVk4d7VLrHDi/kb6W8AoOpQysbmqJU24YnscM9z5hCSzFUb
YTPu+EvdsYDJK8elnddVUSPuMI2urDgk02ClnXyDg9pBXfPd0lcVmwDwsKPGcMCKSnOeP2fQZ78p
SrzKKGgqQ23SQF/2Hs4RM8M+PlkHQx7fcczeUU9v/7Q6LkoCaJj+C5k+Zyi7UV4GEX5p6YjqSLI6
4vy8scLJ/bzchyGahG2jsMJ3lxIqzCOx+LkXVywyQHPQWCVuWZHVAF5CK4ZqfDydYD8fSFhrVkRI
4NnM6iILEfd01OijCnswek6xp6tWsZDQF16ctjF4NOMA7EvLVn84blCp50d7XUA41GrS8dom1CvD
bZpeD8rA6gVtKE8vYZQWXOQ0bY5y7GjOobCY4DlHceDi56keUA+wy5WJKKAybRiPOEqR4JCf6XzG
I68rE/KUdrST67yXZ6d68dqqPpJ3RxSAJL8s0FLXSNqVif6K2ZmW1vP/AwDjvSuCq4EZ6GyE8pjY
ymLTwU2fktySBIxAz3FNLLOMCoGCMPrptv7mtojeMff6dreQAsBwHZba+KYm9xJDgSLII23SgBfQ
QW64IDvZEwon4R9eCPs7J0PNqFAZWMttjZErtUWwBCLabi0DBRXtJLfOJIddpme9ITdyuEMhmpyt
SXsvn7JZrtFVU0EvU3C7LCRBOaPrb8n2MX6TxpkKLDk/bQGbpa5Zf04soLCRyPIk/YuT8ducbYX+
2YnNfnItjFHGBOczqjdi3WX+M7nQJWwuNCXg/v/1rARWXbEPz9jxlCoznO+biWx/fCj3c036SMSK
hUzgSyDPYWurTaFFY/eMO3LlBCs08GidnYgLrU/rHP/scaRiKF/IKoi69IJ+jIouH/9pmGqnetHa
Crid4C8hg5nQs/iYV7kLqMIkKjz4wqUNJOJextuq4H/sHKZNk676mwPZ710ZmdLr0Z+W/hej1UCn
rzDSuzOQys0lmdkUMkCzILPCVoxU4GcvkEGoEJZajRlJ4tXBGTihQXwZaIh2Hfs+wSEXiY8dg5tC
8rEjaVHYbv0OiwNmopcJWm5I1i6z59o24BklpunakpUACRdZRSyvrp5hRmWkkRqzSkz2+O6noiaq
k6ptUtrTPwqA7ge090y7sSeeEgUkdSNpnyuAjFOukmyLBCeKZIbGEewrTEJZZMq2VdczaslMQlu1
1KvUqLazDEiZfMu7K9WMKZ905t1vTzsvmBtJDAxqv+fRoZLPJVRqLh0M1hR3IrHFMKZRXlJwyJRU
0M272W3HvR0oQwUhX6R+NQYFkBDwrjpOIZ4z7c0p7oPgDCq5K0RQ4TE7aXxAHNrF3iH+8ifH50IT
zJeSB1Io5XSUGzMJ+crWpC/ZLkiXcOdCN/a46qxcZD4Fx2mNkh5bW/nNChzSVCHlrqizexAadttN
4Ede5zrlAaZLn7Cpayxy0AWeRgHWETY9vkoL9qmDxTsvnYpEtatmk5+/ZjJmBN4nFclJ01caN5OM
9aL1BUvbt8v5Xx4xDS66eM0jVVqs+2iUdYBr0jp/6ccJ9DbjWh45fzc/zeqklQC+tNAo9JW+9bE0
8ufh4bGbSuPZDReV7kma0duecVW07J6w3p09PzGwz5MtChlKqB8GF8CK/DIZthiscRKKXrY10Kh7
f8y1BDgbsdfVfu5vCsBhSsd+lw2/f27xoru0PpTjUQqBw5AFM/qdDMuJqTqOAOqstvOxr35uibY3
ep8ec23DArOc0JuUmvL/4Wyj5cWVJQZN0uoijaGoh8YKrTWUTzum3PJeD2KrQ+NPY6lqVF1Qs2ms
RCit33jbxGTyA+I/K/DEgYBA7EoA9jqw+7vDi01pQoHYrvrr0T/LbzPZt6+/a6UqUmf01+yDvQ6A
eCwhnhUvxWJiIOunJvtyidxZZqfMg27N2j6taiMtEcqq1VSbglaw3xEdL7jKAIeQMl+4H1l6tFzO
zU6PncN4uQEwNJxBFk2iL0PlsEyYfJT8FKBSCkGcGwuBeDh5jqeWONoy04pTDck3e1Jm0kdLus3k
BeNsCtmuF79n/n8vbfRoojGu6nfW6xsi8FpdXD+F1GE2cigCyYY/asy3b7WAXK0pPGxNsrgSg0jg
lHWE6XGRvYds5BZbA1Iz04orRvZychySRkLbh4XzTTJwe+cpKAJDSmK0bpz/qnDyJRB3ICr6hdqN
6seVJySxsHWXDj4aQ9fvRLQM3Db+DwA4qcXHi1DQuHlM42+zGg3797qwZcG4qmu9i+J3ED2vwtMM
oLZSdMkqJuayiTfvaaN+hl2i2903fnLXKFxTHZTE2RVps4RZHL+JGJFwbg1wujBk0ymZfSk8yaNo
vCGUheztdufwV5Zjn9XvX1Yn52W4EEZfWf6sKVePt33lhTkmGUEaWnPD+aNE/2qmFV4/c4qs5f0G
02i4iuWIcBD3/WHNpWTgu1sm4viPMgMtbypHy05DDoLI3tVmX12/H5GOIaZ/jSnh8cRCvj0+s0fx
1oQg5VYyPqjPmwMkt4m30BdicOjrj4IUm6aqb7ziPp8SJKYGJ464FuDc/vVubhUc5ZjXmB0+qotD
MHp2vCzvXiPE+wD2VvP2bz+M1Gp98oKEUGWnp0nGsN8keJaGAUMLFTK+ebXxK/m4IyKTj0yI/fc6
x6S9WuhSsGW4brK4MGLV0aTpYHJQXduqT8O96gonPGCyon7cnU12HIUF0o5kiDoyRFYCtxMdBrWo
tBQwpbht4NfONgY7I8iDsmbMgwSpp2fTONKNSbjfEiY7FngknxrCEm34+v6XvQHL8oZmZ0iRzzHt
x27QebJPE7DUENX2/NEzDYqgh5srXe8lNyhbEriWcxZvuRrPQrLCogyb74TU5tnsq7RFXJE3ubEZ
kbmqBRLJH9lrIWaiyeo0wV9FTjpxWqfIKV0zNbSvRh6O11cQw77w1rykdp4QY47dUBdtunMvhC3L
wxWx8YaT9yPoh2t57QlR8nRXnSAdZo5KqgssxjBeGD+YerXH32Lu/fXUylLX0YJy05c8lxOwwL33
glAJOtMisWiOr6HR+1VDTTvaL5YL05/X3Knjap7B2e0+/UeuluYqrb0CA0i5LJS95imeG3DrunAn
o4wYhza+9q9mboe9mBshF5T3WC3+4VApSHngCG92Mwe2wl1S6yAt8h8XZDW7kQ1GFBdlx7LAKxfQ
4WQ4yX6JfC4wT9qOgrZVvEP4jP6rVMz0NfasAlxZDwVm1mHxoiwesYbAUxlo7Wt9YyHnO7Q39aRp
4/7s7SjJI26hBpAVlvB1sRERf1NO/qWXATpCqMydRCVJ4xrfarIM0nJfq3xIcfAh/zMVZaOxxU3Z
W2KekmliasoyJdPUMh690lm8B5rdF+9RoD3HlJo5kwhdr+vE9UEFdFyxPrdJNpaYS4Dcs7AllxYl
FXjPwqg/BIa9Iy3J2Igm71mJT3DTh+uGnrwI16PK8fdT05Ra8fG0ZHlF4jOk4+I0BPuuQTsk5gMY
3pctghmjiTAW2yK1BO+GkAEQMGPZvLRqXs0Zq87sPdJrTkH7wB8R5rFN08YMaf4TaTMX1P8XXH2G
d30gmMyJj/OGYe8F9Fcqle8xeocrnuENRiMr3qfplIjdBPudQJCeVNKA4Mvfrvd29ohuZmYi2cyV
5Dw8iHFCM7gtRo51BgZDPRbUXQHojWvVnupH7iHCV8p+Ip0ts05OJxAC0u5BdIBOYDU6MniE+IEX
S+WeIu1/9VMLrPUz6qog6/qJ7QnCKuKHGyJZ92gj0qFl9f2PyfY0L23qzbqDV1RETrsZwkxiIzN3
hcGPjknwW9s4DMgwekxMNmhkskPptZ7s8z+ayajadrYBETEGQ8dG3EHNjAdMjdZj5BJv9l8167vN
a9KntKT2qx2oa5Fn3Nh4eKL+kegDxIHDMNBkumcTrnX1PfU8JOwPI9EsGRlW/tFNbtlfryZJJYLS
/iZyvT2A62cRRSatRzjy5N4UpEZ30XYCtYoUsdQI/+ADvd/l+W+L3gCiVgwwnXc9bNuY3KK0J1UZ
o2CQHVy7y3/nHkH2HldO7YRMyDJ0ncCVXSZdZbrjXSlPqQyu1Jj0On7izcG7ZXLqsCWXqzDdQEnA
YbgiNB1o75QkvxjUHQmQOTdWfi2zRol6vuCNL8ftuuBl4DLbRhMYnrqofUEg/vw1irSGiNZE8NMp
Cxc61FLBxWd38jO4uuiZqeEHMnsQzMA4mEHmxHi31rjQ6VfgMeJlYK3jeOti20/iEWlSAHmaoE7F
2MPFuakDflJGQ7lHk6FZqBZI8ZYm7R4rAfdS6K+yMqqXUTotJK4tUz5FRR7pdRkO0n8SMqUdgZYU
Q0bSvEtTtajC6w6ZhU7+uoD3gnCp9gWg03N+eiqObu6PX3VW5N9oC4e4p97o8Qb5r/rjuY2LiW1z
IPTeT7EsfotfTaobAvnAE2Naa/KNufPGnby0XsIQCH9PsUWzrqwYQ8XLKomGBLcDtxaorIZ7GWNQ
1jf7T0b5YGzDclcmNyYVL2AffqvMwXeU2bdPW3rAKHuHRorQe+tgk7UnvgFSQqm0Q82pTy3USB/g
nJVY6dtjNdTle2kWUzHhg1/7XyRNp28wcN/f/YAV4QwCCj4Gn2UlMJDs5Ok6a6/+zthc0dCf6lwK
SnubnyxQstA7crogV63sazii2aDDanlycRu+71KwiJXGuXRl8wmHQQ+Py9noQTTJ9PO7Wc9LN6a3
Nje5xauLr6CJyWhKxwuyxZuCPh2ItnmPqzrhM9q/45HOUQKcwkyghBeJ8gczxrjwm96oZVcTKoZT
ztdQHm/wtlcQkJUiJNqZc2KDbibWfo6CRAnM3WpIUFYwEGKWNPoy5nyMgzMWBjWdeZdogUY2uVnm
aft0dd3HL35gL4JqIxFC3wi1CTT458LndBVNI/NMkKCuDU+HUsnhUmrOzabZPqXkUKMvWkpezNtt
1YqEnLIP4e3RmGJkY2rSqQXwtXtGGp/bqv+dKW726LTiHrIoMubYA5zmLY77Bthg/tx5+Z6UizaE
Ly3pnIYBx97/Kn5/bMa38xoYUD1jPYe6Uhrs7bOfnBXsYdQVQjIMSY94yPzera+hIXTupzB/t+Cm
XHWHHDsihlJ9hwf3T4cT0SnqTUS9Y5v+3LFCDER19bo1IMvfTa+KqFCl23oPnKB5nFy9UJZwLYjg
Q/7JVgjxTuw2UIDzni5oM2lr/tYePQGRO277SNdy6fX/m3WOEc72BiyiD58N2h7SqVO+QcMwBM9d
LPc9Y/trVof1fHG0yzkOrga9F2TV5iHPQsDS5KDZiSGA8fsL/gqPWa5ficfSwrGRqmmZaBzmsvxn
SlOpWS4GcWdsE4YX8AFCmVOz2BS6mDikUqxTBWJLB0Xm4dRTyU0ydUhQ4mJGo3V2YwDpQjuvVNyw
qAXL31qvDKDrjlDd2VjuB8uviiM8zdyZsC6FI9LjKVEav45D8+mWkNKLagttA474fkO69/kLjAN8
eh1vQU5mjYLNtfhbYpCe4TWYgE7WauW6w20N3G7jv0r3qFaeJlVCIZC01ntJXCIW2X1oYC++AnH7
qVDpO9fo4/sqc1tOpuzSvSYQaLKt5neZYaNMSRIyjwuu5sy+28eUL1uKslXwAyIvbF98livXC4jH
dGVrxMiX5G/IqxTg3cp9prqBw32X5dJ2BsBEaOgkGsexv2xWnr5ND1GnK95w3HGI8tKTNFw57rVM
UD5G/7uw1pjUAyXD7l+Wd4d+yzPFJhAXv0YH4irxWk3Y7xHrgzxx/l0PXFW/BJQrkfjd9tY0uo2j
c/s+pnt1B+agqi/Lyz2emT0Qik/vVrMecaNud6k+pPblVm38autcqp7ruCYHZNg2/vDTIEj5Np9p
aJ2w84o+AgP8MMm2jLzn6NoZb9qEkYskXFFiSyJ2jtUXRUggUAZfUWJXWynowo/XLx5HTUJIn2D0
YbBuOtKALbthExiiv8A5Tkn1pEVyJemm7f5qWUc0iSDeM2iXI0nd3ystLH1QWRuydZ7tFeIwzJNZ
gv/LA5Nc66Cbl2P3NMLvvEABCexq4Hbf4ox8IVcjYasSQNwcd3AUd9iD2tn4z6bW4GXrUBHp3nDX
tt8HPLDZuHeXJi9E6rCIvi/ktKKLtOAsORFVtSbBlq4YaIMwKa79CQRtw9IqiGMixL0Mmkfl4TCs
pnXDW/BpGzFhVehfooq5S2ldbQOE+9spoC1AsSUjSvst1q0xRNpihe/9e0j+eyUenz5nvUtCVYsD
eGAasjmPf8GveUqEFJhDXd/7tv9EsdvJOQ/2dKmTxVpgDERgfRQfieHyy+JPLYBgbm4/ta77R3UX
FL/MYk51P4NwP8OR6Lu4n7QSls2ESL+EfhGZSEDHQpHMn8mHH6jCO7Wh+4Ze77gpl4LnrFFnH2CD
tINZMYlhB1w6w5oUmtrHU3iMKVA6WfqK8UGAAgsCX+hN9iTcVKkWiNoE2Z4diMG/fZZ7M+Du1/Gr
iSc0HWm9EpxpM3vB04ycKRDO6IYERCxMFMCik9Z6k7Qt8s/fIp8HYjjUM87ndukQlIp5spuz3weh
mQ8H0Vks2cQlaly+LVuTKw9X9TRw8p0thw/tLiLStfYOkTKPwzcaM/ndsrQHUsrrLIB6KRkCVRzY
P9ye/rYDUNgbnF5x1a042puTD62TEBPoKSx6A8uRgKoGQ21zGg9YmlssBv4jf6zGLoekQcwB73nB
3mIylkN+LYrJUNNq5B16OfEni5aCUkGr5TS1yoTcXeQoyPwH+96ekhO+vsCYCRzaSI78xSUBDBUo
xqXIMQ209p/amQmwVd/W/+voCR0j12/zKW35AUqM6mU5UpG+73kr5ct4NsjEOknzVUseH0Qf/TfH
fONOvyn1TqBKH4xp+2K924OiHMmfEb9q4H5VAz1LpPp6Mi536o2k3GYJPQbLjFZy+s100eZ2ZtUL
me0rrDW59wiJBYIKz4yjUPekWkBA2VntN304vyRqoZu9QsClQVp54wI4cmJt7wt7EgumHnjAwG6x
ek4QffOAUcDJY49MXi3bcm27rM+NONhe/OXD6o57U1m2hzvgWba2l773oY4aUA+5+yMrh5ih29XD
tdEzxIfxGnIugGpHVnvf0zHUt06GAKXIgS2D6/6QEGYdOr47/MyX18lAehc9nLqEkKUVOva5/+qI
BA9mNfwehCLrLeVLunsTzYGWQ9L11jHQNxnvIhIhDSaJEvzoAnFKNoA+ivh/y0pIp6uAQRE0qCVS
v/QqKvpSd2QJFzQMpyKvrfiIzank3pOKg/EL4duhM2YlT5N6ym/imVGzjs28vlYJkT+3oxB9Qpc7
rBgeYegzvcPgPu5FvnCvLjHTjtcGqdJ9epYcVI/ib3NKjAC7O3r5rV5HY28YT+XHswL140DxXRkT
MRyIGdCJTXBt4Qrgfd2USrcnGbEP7SRDFRJvkdYnBIxA37mAI7tDtKOZfe9s34RHZISd4iPJK8D/
nYAgYyL2rl5NASnGWE+GFFJ+TxBdsWKUuP/zxagCAFRRAv6YKwVfajy+fV8yn6M18LVNT7lz7hJa
TwFvGrXVv3G7qrHPbMkgn48U7YXTvGMqTc8IIqTJXUwYiM8jyRcdp1rCct2oF0EJk6lpJl/x94Jv
jz0ypiDGfFCef2RaKv55jB0zzRd67yj069D7iDQJpJCCRrlCy6H5djPxCGVUj1Q6IH5mV6+vWcqO
s0UwbmF94ZFcg9VsDYQzVWoMkDkCpRLMRiF0ES4KzQgHzPw2SLSp/iFNP/lLjK2RJOF9nBxKZJYr
/uTDxOD1LoTutbKWmwoyyMbPgHsxNeplP64H9jYmEB2pEVJ9Om9hw6ZODhJbo/EXMH4wfg+OGhIY
DNybU6DKy7DMEVuGtKvZxuPptOD7nqwywIhoZhZjetANRtIc0dg6jpZZaAEIb/1z/RIiSo36WoV3
X+xfSW9rfSbtd2xxhlSDuTvK4Ko/PUAobwPT5JMP70wlKbGoJ9XvyeiBnYJJUL3xZvAUG/DTSnCC
avSqD/oGRcmOzXuWrp5mrroysLt9biICh30tfPVcGxz3SZEpFa/sq4/BgdXqN1zoDFDIuDWXKVaA
x+dni7LRExT0PwIJbnI8J1HZbW4kpdJK33gyryPp8LgR5bTFGeGIJxsm/924se+ej4lcwFEsHpNF
/RUrBfN/ZDiV3pm3bCQ7bucKhF82rp7ODhk8rLb6Nukf/E/I9WgCoIZcmshW88hEOSon7l+o6Q46
4sE9r6aO1Km0GaDmLLFm4wfwgTIwPga8T32y8ec6tHkmehewzTZEd3AHzQhWq3Kk3M3MGJDvrBtq
dGpvq4JhK2+ar6QpKnwiTHiCPffKsoLhCgrDy66SCZOlP5bQVpZkVDTI4jcBSOsGURyN9hJj1pqm
t8uZfc3/UkfeiaPRlrGno911S0VEehSRwsDWqhafGEONgIHFkr76p7Fgip7N20gjyK5lsgc6+q3k
RFd2kRTbVoi8wVtoQ/YQN5/K9iQHLuiIIF1WDK1X4JJckKYJiNGie20WMBUh67gYhtwKN0raJLCP
vMCgJOYuItqDsipFdU8wv6d9GMpP0Oq4aVV3Kl0U6fSx+oItvaaA7WTpWRtyCoY3iZkzpsNYObFZ
JIf+A+lSyy5z7LUAP/VOHEfjAVpjCBxOhn947OQ6DlREhqpMQzQkhPhpoLj0ScOQKNikI/Vfl3Cc
bchG7kcVX6wMkAa92hk9rG9gwo9ahB3hp6r2KmUyqmVcdqxQM+PtVo4cL+khukY/aCnc8lR8EZ6y
tezC+HEbmQ73zHmPmk9UCbdyr6AnS4n7pjXWnduIGG1fzgbM+yWfLeMDjxxAFjOL7bD2BJXSm7jG
LLPpGz202hohR1dUWZcMHpGTVlig4E7XXxND/SfIpxS7BcQE3r6uEZICp3zQGnQdLeSRdlqCuMft
vPfV9hW6eZyNeV4jLfa5l60Z60KMXtW1G5Ti6GBVunei3zRwPFxfFIU3EMNvXo7qgP8jDLH8+zMf
UyZ5XSTjZ1AMo2KMgAMUv9UPjc3S776MFVYk3w+YwFskOqcc5ZU3DMMKQe51Ql3EZPa+3eYx460f
zU+/lEtwOnvWuMTrm+hMI5m72jjGPGc2Opq1TTKdrPObOnIWW31zk6fPi/j1uLBYjMe1fyFEfzyP
6OpMY8YU2+fA3SsLXWwdRXgzfmM1wf8OkjprpJE8bopOMC0iDXuYsFbdFq9OyftMKEJzqWszh80C
FZ2WJCfGngPpMzd9HJIYPDNh3p6jxX8l5rkZpnHqqLMUl3aEX35xzgd98YKRP1Ln3VKrpxGb44Sv
HqqFhffKDaCdLdQx7FQteznltx5xtXol4kKFMsS/7kGPtN21u13pR3rNvxEJUxXE6DNgavZNKQyU
CJeQvflxNhaRnXOyv9BZk2yflaVWmgzaDk11/BK2lhMnVgfADuTa9HAvDWILZhV18VzuISMVHy+O
6zUrZ8AHWBo7FzQrCxhl3Qc6OviB+myTNDV55ZEJwtd74M6D+hujjRhHayyjgiTvx4HOSvLPY9m2
QZJ0fmtoykPHcX7ZWmuVZh/RP8b0RxmG7D9c17ACIQbGjzUse6FSWZieNJXxVHo+fcTscjvSMuBq
drhjYIB1HPkZXAM4igeXD7sba1odSNwcraCess+Oz3Y+/nucykSB/B+LzlAhlUP0Wx9scHb2Gmip
soF7SRyQfPxDFWGo4wQuJIx9Bs9QXGScwk/CrEuc9XuUg+0bINxq8Q5lLPVuxp1kMIbXuuY3BvOM
7A/gz5CWk4W3k2/OGowPoGebuT58x2C5DQi5+MXSN1b2K5c0s4xFHuh+123C/csV4kHInkROtDgn
wJuggTzOtjLAFDEGtexjmdz334QCOJwUR11AKVI3+tcmuSBn84NpmKU27z8Ar4ZHagACQ5Tfcltr
OhhYJmAy6kdWfei6fyxWmqwH/mCtj9W/xT2K258gKjiaJTfLp7CRJpHLwOjGnjN6mdtwHPSEkAcr
N6MfRRnCzM6J2cCIwzuR0c9emTV82VARqf2vPwCh6pADPxBS8+n61o5xgdJlqn+k3fW7Usx3SnkT
A2WUe7xjS3q+pUETimYR1vQ8tsHbX8UkB3czNQGzPCtfQBcxOyWC8iwJHY+GLXz5rZzsVulS79EJ
V03sVSPbNSG7A7xzBEZxrkrPu54OTa/nKQPxXnOyn8LPXGQjd1s5lPoN2gjPAiMt7CFwS4UJ44Lz
5op9vZGq2/0KD/MtSCd7SVF2GYLDbdSQ1fF6o6K2QMScAwX/hGlHyjSZ9B2KQ3mUQmXVlZLP+Ahl
nGazxT/EXM85mpFzysdeKRLjZf3Mt48H5Dti/ig3gNsyur75cISrT2lj1Xj2OlgFWzDOxdVwFPHZ
kQ1XKffIXnnjV/dUH7KTE8+LG4Jc0q8CJGU8FASJ40Ck2latrV2NxqIyhLGDmwT1qAZzVxYP58cn
5Gex1wgBovgdArhj0ziWpnupyiw9oZLZtuLzDMXHU2gG2ekGZmtXEAieT/GIMEYnpXraiP6tra5s
IXET10QY2Z/Qf3lYWdast2JyfI7wn1yBmsgeVtnepo4E4ln4GdIuadBvAlsWYiHO1FoRnjh+QS7a
vN3lYNIIHYMNi+TOUxb7zpjsjVlt3nkm61CBgXZSEMdWOJlZLBs9w5VZMi6QbyNwjo90jKHLmJpB
HcystCCxUDYYEsITlAUdgQvRb6BSBKIEHdNUYcmfDsG23pPFOJJH0SdXnABBIRtQi7z46HuGtzBi
P1lJ86U1+gwDhmyWUbb/UH/G68bXe7Qf2oXCbrsreyc75lFMUdh5qOpiPTPs+WWA/6Jl4js4J2vc
owH/CKsiHOdrmV5YoABNw1rVhf3lKTkjydbfuordMztabKu0KGNFK19OjoAsuUOxB8hD0eFaKgFD
n7KIhCcKTUlq08xASbxq1q0pEPtoSdoEKfVBqI8oYdDlfu9SseWss6XeHl/adtEgIx4kgR+axL71
FmkchMciZ6EhMCIXybUKjHofubTkiD7WoPsIufsw4SzIA4W2VJO3LmSgunDpXK/Z3OcH0vYZMEMg
4K006SVgcOZcTn+rUdnA5hw2ZxgwArRVd+XT4mf6GowlLB78bvJk4s0JtOMJ5RTYHmTlkOVasCst
jBWFU3sg0Oiu7v97bBQbv4TAC+fWgDMwF2RUBmjZXSCfEyh6crDWRv7JLrhaLSEX9hvrN90H8sLC
yAKwA/hNLaUSn+vL9FUpcO3upQ5k4NIHecw0CNYX72Mrqmr5ry6L7mV2TLu/tnZ0qVmd0TqSABJv
3mKgzh2bdjURfQwAQHVyRT6rCFBJ7zl50lw4+IfU2lmrW7UvzhD2YXEvtvGB/tGQ/HSigHN8e2Cc
NzcpBmWWNxxK0N69R8HEHQenCw5ERwUm9hjWc0KDQDokfnFDkkdjiTEIM3NOcuJDOvhqyybniY9B
2mePuR/1uXP28L8pgW+Q+unHH2yi224l90vrXq1hrFFm28+dlVpqTXwCUedf5/FWhc+ktBxRdnEm
tzIH3vpATJ2w4kwKNNIfgb8G68Dwt+qQh3cqQlKa/FOR4LX+BECu/BV6CY0dXNwnERQau5L/liMR
SiIE26IpP5nFhoULzNh5Zi/XVuniPqmIuUXFsrQVWIPLLte7sP7Tin3yMoBLO6BQXiAstJ5DhmBS
W8as0zXLwS8DqYzEY+GyAFUwpqfnkmZB2RiVSbPGTbZw48CxczOeZyEiwC0qZDR/IWvPYHvbd+Vp
kAEDvX+RLqYElTBdH4qXir9MOCXREm6i9yuCbG4+Jgxki9YkRJItQ6INouKLe1YEEBZ7r5x0cDfP
iYkFHDwBSYF+yeS3EIKN30bGyjjtqxkvIqPq16MDk7LRAIeOhp/z4AKdwbz4j2nbJ9dvf92wf9Fr
bsVWor6zXoGgXBkBLjyB0gwJxa0zU8Zw411kEeKH/rh2UtkjEQDuQlk5+JRPLN0JLFha7QCICLOT
xewzLHT0W4jPQgAzEwMhJDfy2qKogOkvLqtxhSn+ujTzykp4j7n5yWsaqjDHp4848eyJio9M/hYO
6+t5ZkYzt2AZ6jxv2OLA2nGpawLxRObDx64gvJBPs49MdfHkAHCEM2IDkJwD6k9FXY9n/Cnj+cSu
+xrVb+Q0XImLEcdcoA+2cInoRMxX63/AohxRpOiocxRLUF2gjnnjk2Z0FXLML2qekFbv0AfD1FTR
WophscqjuaP+L9x2N8LrDaB+kn5e2mK5eUVrn22hauVUlr5feBbAyIMv13SgV4lPiSwOV3dyB1XL
z7i5gQgnpGYxAG56FYqkwF8OCJdJwMhqw1uMI1Su9QaOBRjZhbwn+pwlEhxLe+S1Man7aYf2BP7m
snZBxs0Jl6+jj6wIFKrZCS1ZAxcWlF5tobddr7MMSkFx9AfmPFO0zTGDWd2g4mm6Jhbwa3IE8PsT
Yg3WPBwObye2iv4RVPtzCx2CPZS7L9uGAK3Md2IKIn8VQu5cdkAWup5ti0aSfWMC42Mie7FblmgX
xHEys+oVEhu0aJvPJM9i6YICFY1jIsoEeBPuWFl1+HyqRHQ+Pf46O0S1ElbiiY8fdEeAt6179At9
rnaV8spzXcW7AD9KLbJuOQ81+RSoSTA0Ooc+CgOhAHVB3/FQ/bYhtivBKGCAO1C3l22VfABp02LD
2X95YwTdLyJqRBTdajj3Klz9H4U1J+Hp3CTE5SEQaXcCGblySEuYUc2wKIV4FYYRGnaGSIfZ3GYL
fNtSKLxZPwWiiqtJjJd0IhPTATkZCEn/FiLdAL4fbdVj7KI64uJno99eEzYUJM1faXcVWOTejrgh
uWnlGnGN+e/THuDaDtL8Jtj17TdvYyK8zZB3070V64yK4kILeIZ8Iq0lLh2Ox58yfKULmMr/g2Sy
HT6NiEoxq4/i7oRYc2sKYIRmuGV0eNXvd7uup36VNlap1Jg0Jm+IPruSi6ZMEf2idnPjiNit/+Ve
dtEESUbMlTkTNljRe7KSdDo5nYCCse6SQaYzRlmUjJTBe+YNjUQkVLiP7qPNilw3dZxtexjJTgaB
KtiELCtS1EnAwgZGdhqRMznTXbLVlwU1evqRKFQVK/z7qbVvJfiWxsHFHFX5fCWxThWqwmyGe1zP
OJBiIZGASgCPA/JHQTQR7uaairC8mOY7pMqKsPsrZ4fJt0foG7NaSsJws8SZLlVv+CyzQPuYLJU8
Xuncr1CQUCeWaIOLJ14G/34aWTq9YilVVUxr/dzbxXMLGR7xMQ3lQY2PXTkk9ftGdxHnrawLKe8F
Lldi5QevYL11Iji8daN3Q2CtmdVB61eIZkY07nlpf1SHN1Vx1IBiO70o589vOrk2qzVavoPLF5Bw
rQttRmBip1t1KkZesXWBgtIry25EU/RL+ho1kS9EJYV6IFg/OSYrDcH1dHRYx/6i9UWmL8JYtHJH
yvHF/AtQy+e7uavHM3GNH1QlhshXHYU7EUVq94/EE9Gh3nLn8l9S0wYTtbsVvs9MtN/Wmsgtv+6R
tqa7JGs3beOfJXtkVUMGvFFX0UC87LER3wu1+2S/2vgfAwCtCP/rvRbGkVbIJ8+qIdcpYY17GSee
q8HByWVp5jGL/6asqiVsi+5hsWJGyHLfLVsgvcHmopc2+nV5j/gaxBor9wM+/EMilrkoOPy2z3BF
4ywjw/i6+A0uTLgxUlEBujYKwoKGILPAOn/J05+1JvdlnQG9bQUWO1WIQc9cqbbd1tK8I+nFutiH
N47f1gl2dO+KxQIaLNxUe28FQVnknHUjDfa9XXidx2keSo0y9qyzlZbDmw3ozKxTJTwbokhUocFC
L4kbPEW/6tHcq5wM93xTzi0jUbqZrXSNT+q8ky6go1nQwiNTYh7hIfQwX0QjiMUl+m9U64UoHqhR
ThxJsc4BVIzU8An7+8nlfiF0+pyECkJqqqTN25B/kGoS0PWhyw7XoE/6OlTu9hXaurA+jHsrIJ1D
h5AXsvOg8urcEbkDlL4wlYmpDIofpo6x8BuFr47LUgjZ5c+siWyH3Bu8RmJ/bO2apKCoMpuC0eMy
saUOd0uHALuWFIlJilVW56WWq5rGhmcvuQ2EFrc3RlEO4VGO3dyD0+A4YfjdYs0GG/wRTRy9PuqF
LJSsThjpitBMp4ttJal2ILBLhAJkEL+4ZZsNUnOvoQAEZDvmXRbn/Et1VbwcVnM2BuzQugJDXhxO
LZyQE0SJbCQNLFwqYhVIIdj4mb7qdRrx7yK9NgQOfv4g6hKcdcHI5iVlUKV4S+U3SUgBQULOn5Ny
ggRdQX0bkfdCkdLXESFfeGkTWEneSxSiTSQXeL9Zj73klJO8Y4LdubVEUOiJZCWJKrHW7hT4PUxh
hE6I6G0O/YZENJSoPpwQ2X3t3oRlEglSpEh5/e4sqIrac0r5JuM91NCOQDh4F1g2erZ9uIKB1sCO
q+B6scl1l+ySZ7QbMjJMKtCtWtKdzSbnhhB6ghCevq8xmuaxkEz4FWqSHgyKqMm6zPeHR9Og/nTK
Kl1eV62/kBo/6baSRcAkJ6pY8HSJ3ceNCdJW/LNDQkvQLzscjludR0Rr1cQj/u9rwpT6V2qdW6vG
cVoF0BfjYplTY6N5Ig/zBSN5lQTV+f+KbY2xcvhFINAjMttqkyXfIsoMpLNDzvgR6E3yQ5ZDD2/f
2YzyXupF0pUMw+hP2UYg0GHsJ0EUObIfGUqJglXjPMBi4BWDgAHuvZad0DfAA6a3ZRhr6/t1E7FU
KoC7ojolPQ48uANkCxQW8yj3ui6PLNLh84IlAlv+VyARHeO+yBMbZax8bKzS6rP1/wk3UYHT7GJL
2Hp4PpgSmlq65XeXb12mHI/RuAJH69QdLh50NALDPhqv1ykZ21Omtdz40M/zgYba8O2cSG1xHAcQ
Yw/SFo8hIyoqZFhtC4eu7ZOi43rfERuzi2l4VQHolcfRf2CM5I2rX87rlgcbFwbvwDo4QqXKdIiX
yHYXS/o3+TmJA2vsUb6JydGRQtRFsgIbxjhvUsX1vXuWvhrr33EVms6X6QMrjjqxLCeSS4hSmCR2
oxDyxpTeUxhFIQRp8kutNQdTNufbnk6uphxQIb/SpRjlP14hQE2ufPPBOh3zjdiWoMwVjDnLNcZ7
FnvOUzNraf2o/c5NZfLnf9iqs/FoEf7e33+2XNBNtgXHy4ym6viKtdJ+ctdW952wHTGbXTL+Aqpg
lx9u47cNRW8/v+ug21VFUwEKcpasDnOXQIMquO7UrCEQCDPX+KsWNK4GUg2pmiLJA4Y6UFxa5QNe
nUoNnyipSpw3sv0WFVktUNDh7QdFoZDHzpBm6GYpLzSDtQzcN7QG5sw73ojDyQBKgkq7iwAfwY8O
qo1qSypaZFgksCEvr9rPKYSQIHSdSPWeDXkhy68KJEOw5/3B15tiMJIDodGUFRSlJMoPWah17nPa
WUjxuCjqQ08Zu3+/9nc/CfEIiO/VfYoYCcagboMWLB4xihHY/81VRdqsZf3JP2voW2QGRVQi3cMa
OlKIK0dEPO6GAVKcmCFYEyWpqAfK3YwvCbmTyr94BTfJkhASswkMSksjhEGCWJMzHyzhcEa2UQIY
g+hCXgvu1ncXXI7O2zf3EXMRJRJVZPV4JfLpqIFivtGlEbmHnByWai+uAfw1plDZtKxUojTwwQ+g
3bcpsTaWUAws6KGC4rJNye16qoFPp6+9AK34B1pgJMLNa40LiH28j9MauzBQHs+eZW/Vd3ilDynm
i8nHXCroIEChUhTpOPW3r+3XPaBatscvEA5wrJ1g6kPZNBXPP75HtMtJgMEf4o9KXgnitNGGXysI
cKHBkTlOCPbyCS5+Pp8ZJ6nju1EACByJlyTzxZusg+1WFsAkfOm5DDx+IqM8G8LHo+pLcDbv4cXi
jE7vHb3/Csy5w8xM+mndK6Ssvky01Q7lKjuOJeUnDBDOYrb6uaRgJxYiyiSXtf20eMzaR4sxdyb8
EKEyF/XE/zSH04bnG9mT0xqn2lrMRnYig8YysFA5ir/Ue+N0B/DNojiG2YmWiHiKX0XnlVzdxpUP
R3kwi2GxxH/eMoV+uPEbGE1yNpoG0s82Uoli3/tdXgiddTR4gk7VtF4o5frh4sePM93j0hCPSETx
SeV8ecsq7Ve4a1/edsvSAkx7Hdhd3j06F44iR9Pwu4heO51XumgT+AcwUiPCbW349Ekamdpkctel
vWa8pV+an5b87IXokANoJxGRHag5L8rODUCSaoPETDUKTXxDOPYwsyWrzBG3LPFakRz8KmypCAU0
q6qc7KwpR7io23Kcto/dhcmQelBmowXwRYd0bVGM8dL3NahCNQD55w3fnhz8Ctv9hYUZl8Yqtc83
8TI/sff8jpXjV/pG0krBCdpdlk+Ciqci6zTTHhTqUryFiFa72XniI8PjBEm/uMg0X2N7qcIXYdZS
1zB7V6t0Cmi1p/UTBwCy1YAwxDv8kj1wkeKBzmrwiBxn3ot5seWOv1/8w7TaN/MBC0sk67Jw4E08
Om9IbayvzQw1UUDlisql4HiYrGDqXRLvYa5xyTpo/DfIL9el0xQ4YT75kWLDPyMUqAZQjLnCpuxG
mN9k8bsEE0RFYgZjHY7v2OiNXHczTeNKn/YWsqkl/qwxoQE9Zxu1cxN00ipwJCN+HcSErO3HGaLX
1WAJHFPO++DQyq1Mx380O+A5sRcBi8SC9b43lYqZiDUiqof7kxIGOEkXY125G2w1/OcTjBMk0pwW
Or0D5cc1ayiTydMWaBauPl40jonIvAKXQdTp263E/oLNdPbuQy0tB3Dvg0DwMlAPQAbwctetfBQw
7ng3EM7wltXzKlePxLRoGxTEMFaOaAMV3DawHm2OlKfyD0AcueVaM3l6cRCkfVlxvkR5sEGHORFW
7VAaEmYXD5ZA0NOQyTHdX285Wy3dD7PRMYTCiwmVD3UIJUZuAo1k7WjWacNHcsaqMN5t4XiLG3eW
t6h41hqGLtEVga26Dc9PjHphx9G4ZClGEq269g8miPoQyE+nfrc3UqECl7khzRfG6tbDQL9YABvY
FLINuOsGK5apA4B95QbA6aIblk0MV/uXsDdwG3+nEGxrg3e1lP6bvg8GxLFHtG5vLACKkXQ9w/eW
v1guClvPborAHJ4l72v9swOIHcLS8Ao+GLT/1PdpTuX578VCO9XrzWg3e+OPQMbtwE51Fmm1UTuW
bNJDiXvTe+YpvvPOtq/mqgEyVXSvzaAjw72kAAZnaFpAd5uNnw9tkQZPcLihmK4hM3En7bS8v5/k
/efd6cQOIZucs6DG1ch1eF3hdIUWnbEbPxVTirPtdz2Frxpe9Z558qyLMOHDOz0iQ+Uuliak92iB
/odhWdpTCdq+m20dheoqHgqmXlTokL4x+Ysv6v0AbiJA7gUYrS+4QPM7mAl0KQUH8pckf9xKB3oQ
Rp6ciUQFPwBY+Vz3fpqCC5plDkNavCrDt6BYHNlXtClb3uf6trBr0fPLnnB1q9zUIglgMOySRZqI
YPaDcMK+wEsQAkjdxOLTR3dJBxQS1kYBhXh5dx6nyLLNsd3BJYpdNaBtHiGvY1QzrHYI2NZxjeGh
srrSHza/9qt5PVOhFM/2T9j9AhIgtS5Qdr2b49qbcbekXfVP3ExFh/LmCVqBH2NYKdZc/OkS/5eW
wt8TuWTUyJTeyrxhIA5nArxor++zyQjT6po2PIeNDuPhXqWu3JV33ANA/U1yBS5zI9R4g5je7Dyv
k7kyksaQKFxtEHkyjl3YrZBMc1Pv3Y9TzQvKyTOvA/a7Pqop9d/Q1uLKnwvRXW+b3e99yyENfPsh
WfDK8GlH23JApnMoiEtXYkhoZ/ZcvqaTRIM3h52b6dljBk+LSakCR1Rmcg/AZqL4GFsDwcUh6Pi5
0lCtNjonCINY+pBKIjrCv6f6qyWVQJ4L47yMktZ6vC61FUsyiuu0ZA6QPSiei0t4tOvep7d1Jiwt
PUbWZ0Gygg9j3fV/A5RuejzOk7ybcrmVRwLfRp8sOROBBaGdJZnHn6yQFAyYFuoq4OIFUX5kK0oF
9AUMXhrhg8nEQ8RBl9vdCLv4bAK36wOvqqg5QKlNSD9DtA7attoPLsJIqcYWAWQMYlIVIWoNt29C
5ZVrymATArcZzQxjr1lho/Urj+2Duse/5eK3MCkxRuBHpCNKqiNrZnUQdksaxSRA+sB+eyvvGHC4
l29Yg92fEKRFhD0kcJfoUioAwbFCgtZdWT/2u3VXVJYpokQ7/+FT3C5HQthv6SxnJo9wi05PDQ/1
DXcmpV+83u6PepnXgsZN7U7fsCP5yTQ3/vXLwqe4Tjw7xTs2Plc7AHCVEvD6DGBuTyxMzlj+KyL2
ifCt2mT3eL+cucRIRX70aFIUpoEghxMOlH0J+36Ay+YUV06NAlFOd7PB1WCS3yr6O6PY0r5/Xg6p
X8Dgj6FDTyuvAnC6Wh3F7OwogdlCewTLLlbqyVgbFkmr8FFF7Wti8A1RYDC460EXt24UBdK8rymH
TmcrJ4JXHLwVrizxx+noH7s6Yv2XqezUL2+hoF0E2NvDuw/Zo9rIkTnc+Ruy6suZniSpAze82L48
D7zpWtV8EJeg6/EjhAS6GDKuAKmtNaDE0+Nvu8xLPUZ8VeefwGDYijsqhoC92t88e6jG3DbMmnQZ
bjaFOVVUOZPPMEhcwDjsrhfD03SVfFick1BlCdG/9F8L2OAEWI0qL1ow6LITdjjuop1mYGc3BNWs
qHoi8Jf4jZkzjxZQ0rAc5v9duJUEyHd0Gxz2DWm8vMgVHozHT3jUFfEEts+Iy1ofdeR5Gt36BkXf
aCR227EuGl0S7/VeRJsTHDwdQBus2ImRIebW1B6dfQM94USKxiXeg8eQN9ZHVpQ5YE3UOfPHZqA2
PxUG6+95i6J3GwO3RAdswR26dA6uPYAub3ut1Dnc/IHod3M5VJQH5AuCckmsBk3msDsmXErUp/Je
wT6qk2tn/g3FQAigFPz6W/zfM4cTF2xPu4OTUa8sY9u4wWsv1iHhaavc8tJOCgD3OsSZKK1cA0K5
BOyyb+zq1WsapV9c8v5p37x1ZqkIqsFPh1j80MehDO3OhwpJAjU15Sl/YAX92rFXNg3De7yEogxY
5Ic2aEIOHd6oyhDuL2e6EvBKFFsVYYlFN9G51zRtzBbGFToGAuxCA79eEHAFURRStYiOU6zA5LIh
FKEk4o2a8qGPWJOdY5lf8NsCuIZDqBqg7NKNdPlySgCXjRNabUUvwEqNuZXwIs02AiA25sdX/haU
BQ1kwuWDcx3Tml1GMIL4wxzNOzBxv4XBWeti7qn8Dztje1ZUPDh63btx94NuVr6a/T9b7wC8+N3A
TVpVdeh1+zb2/o1J6dakk4lAWpYPKmwBQm0z/nG6P5lEaI8GEbe93W4Uedy7BFVffuT9LpdjPRRR
uKCxaOUm0mArKsnhBVT2lLifC/OjoqySaDHivDiAK+rNHOD0YgwTWT4JCqgdUxEtevQboMQx4Em7
fVj9qRrVRakdHYU1IEjuVfO8lRXAkl4xr+02KFz02atJtY1vLYfMOVhQzOklnCQcG7LZV/0g/rf1
VjzVPbVA5PwQBaJNk5nLJpuCzmulhY1lAMwYt99wIGPuDCsgkrxPzHvgfy2Wg2JVIw7t0m0N3ud+
VA+paxt0vJ8N0cZNoWvzwE7vNnL6Zpwrpi58q5Rj+U1Kw5+QQToBNB4JhKcR8V94gBexzvFKHiea
KI/JPb/7PjGplSUZEusAeMExWQBSVrwZKw25wbnhIObYCqLLOOlwkUAYLTuWS0MKsIZRu6jSbvRU
+T1rKYT7IjtV6/nJVF8xARqhbkNMksoXnwRptGrEkPzgNhGfPCYBPzQIYjL9XMpQPOuTlvtnk8HG
DwJteaZFR4aimTN085iZqoO9pnYR9UCI1FU1wZpTWq0Z8gBIMqkBX51cxHXznnPa64Jjdhu11KRT
bjiK6rzPRQ2LzeOCPuAGK1tqJObjONQtF5XZfDe1JVkIMUeVEbpiHJJW1zTB/+fxOUQp3oBZI36s
HZxfxSl2bf7JC7pHyFNnO+TsbedYvVQWSXlP5ZqN/eSpWSUqC6az3A9PIiLBJrx6zs+XtyBrKpiZ
dmePpPCzJwde8KGPLRah+ZNl0+16JG4KyoEcWnxzgYbAHEpUjGiO9YkBeKdu35MhMTN1W65f95Ej
vBfdRsjgHvWDKWKOgVZYrkxD3QcUEarOmhLNHa/MqjPm6rrGFTNhQA7PBovagPMXQ6fnjW6CsrfC
M0e0FsTkY98nR4/dfxevT/zhJQ5BtTYohhc0U6AIgsjGO+Ak8eL6Yvh8XVFseoE3RL0Ney7SQtp2
0U6d8E4uec6SGg3EIiByvX0sOfFRc2yyyLYy/S0Ics75NSAAtewLC74qM4LhmN/J9C79fM4sH9zw
MBLlOrguXTE1MwCcio7E+UH4E3BiIrWIeI59HiNukBfH3Eg7OTPlKpFQefLD6pAYj76+NAJbypIZ
Kv7wz/mH821XAng9EAlK0/leOG4XD89FjidsjBRreXb2nFU4klOD3d/d7dmKUilqcZEtdxDBAAbp
tRnU7UD1st7RCmyp1J0mHZCQtytA9Nx9WpsAnZO/w1BlemER2Fu6XaCk69Du5b3hpf8fVrhTDXie
39GATGOK7lukYxMnRNCte5NJ4HCBucfiZHj6eHDXautmLHh9Z+DKHbGSqA/ImTyn2OrCLwlnXmTO
j7e+hNhbR2dIBDLqgx7qOQgThRm5oqBlFeIDSoxIN3vhTgkIz0FVBb7sMqzzAVkz5tGmgNq8/+pi
CjShmomUjAFo3DA4rwyEbZfKvlGFOqmYDE9V1nO5Ob4DL69OXtR/LzmhapASPhqh4ofPmTzCaLH0
9e/DvJxUtYgp3CwshfStNEFEMjcplEN2OOZl/FG8G74/WIsx/hAPPXPKnkmUHXro/YZ5m620fKMp
x36a9Iin3cM34g39wg349vIyFdZpDcrtiTvRiGlaj0G3/DO8TJBGRgGZzNBTcmXdRRnq9eS4Df2U
DfZvbrQvpDrdCjirjAgHcjnlObTIZsOHY1GMewDYVsAko6BXQR5Sv5JKH00KEcoTkPqBKmv/0x2M
bji14zda5lklsxnKU9I0WKXCpLSWLqMetBr5E/SRbTjb5WBY6JYud1fjFsV+GtMWq0JKgqZxVz/E
W0aFcmfuQdpojOB6QvzP1e0dzyF/VQpw7S4mXtBPvgMLTBFL5XjIuKi0G4KJnaOMLyQUIbThD+PX
9AzS0MAuJAx0+gl2H3fUMCFRejSOQ6OAVZZdPJUn4LYn0NLktcfhxqqKcY37d00GA9qQs2njmWJG
th+RBGXhPHZnUmqE9cweoXOqHmuCC1kOr3Vcb4R54lkpiqY+97QbDPO3EH2HA3uG0sHIYohV35mr
aWwrgU1fyIz3wZs7ePUzip/XkgfIdEOG9CZNXaAJQDnI6+Bo6kng/3THuHdQ38cdsA7HKQykPfem
otMAhll8O17G9Huo1FQMlxoRsX3rcRdQQpO86tzrW2pIVKxvn5BYzMhIdU0CnlSppFoMVnCcilzj
/CuRbN8SVib4Anq2CwG3tz0+wblCHQ1YdlaZxl/zh58oUd4E1iseXy9K9aNxro8gc3fGgm+299M5
rwYfpkHKfqd0no4nGRTeI56287HiZGLh+lDFvVdM61Nys9Rqn09Slxn2Uu7lV8W26rjVadrmhZky
Gd0yipZeq8kXl84VMFZdl6xMVhV6QbJ2AGfiGpivsNSmzL17yuKgTzJhN8N5dyU81y21SKUYqXCY
sKPi53JwIeXErdta0dqPOK52XLJfxhFjuBu7/VuYzCbG+IVjl5FD0W83cZuJdCk+DwRKEYLRQ0ad
mXcRPil9ZddmjXPBG32MaZyFciUODx9FEcrvVPmNqCf2FPG8GGq/PRImyya6wvWuiRM7jJTZOzux
Y35+zjF4A17YryEbHjfjHU43JXwJ7omTJTA3BRG6y5pNmz9DHWyEgoWNw5pryt1i7mik8Et8Gvtt
b6oYGEE8uRjLZI1hT/58BpoXzxSQgxmISPicbBMbAhC6wcW1zr8vFOUzMYD9DZYQWnke3FXN6DJ5
E2QCB0TtVHQYDAKog4TLi8i4mLL+i+3c2CuazlYOlABEbh5rbVlvc8zC34icXMSBX656EWWt5ds/
y5MR4SfmPQy90AMOzAJAXwdbC693OMroDAfZkaR6/fivOIb46aoEQqm0S3wypNOznGluMZJb4q6i
YZ4tpyfAXpOFgXhWwMrFNOYNR5imYFxzZ+38IHGdI7Sm2PDcNMTrjBUaUUVcYOqaEb4LoQbSwWn4
aIdHOCGCZu2KPgd5nL82m5QHUW4aeHJusFg6j0jE0A4ZtSBuU75/vmNTe5KZrfCRu3m4Z9Cdr+rp
5sWfMRnsVClRHdkquYKhoMJos0Ry1hK+QEnlhuFjMIpBqulF9jDOzDpglgL65psk2qDlia8POvrF
rZPHZP4tvbJUG6niIzTp408xiwvtCqDBkKJ5UKzBf/pdNN/zOjcr9vhv9jLgcrTm+W+GPteLs1HZ
0czMUb2Y2rdxALbdFFqOrR7Lq2OGTCNk7Sh9tZwTRE7bQvENtl30aGqjfYuGgHE7d5CQTQ57kSh6
Hu8R8+OTIu5FWUWaDnDjEdEqUEAl/8Zvd6nOoLWep5ulld4DbevKj6AEjC0iX8wGip9y8vfCgn29
KVpDRtZRTsnn7jxPDnetBOhvxoqj8/LQH/qfEoPnNYnRH9Tg72CwHWtf94hM3Ck9nLsRlbiOMKde
K0Ghbc49qSx3Ok8b//jZhPZpYD1F8HHEzEm8OdXS5LC/jFdHzRtC6fuAnxwNUQvDeUlxPvdiNlPV
HHPgaoWjin5MqzShnBPIUUXvswk+l7nHqVfZ8+PdWLu9miWi921dYMHNdKPeSxbO/WlvCPcDi3Rh
DxNecMuDdFUII5/Q+oYc4LnntTxomZV2WUF7a0IqU2f/tLOU6+O1w6Aj8GU7YWQ3oU401uMlfFBe
kzZDbt6H9b7BUJX34F4ooogSMNUNO1Wt59ABy39Xwl993qa0JhJnjB/pOxpn4zk66FfcJyGGVzml
nm8unhLO6plS7sa4rMQJxDn14fh0dnl0pc6QV5wA9UTYuQ9WqoO0rg0yMyiGiWDK6+1I2yu0AYNd
ecRucU1hyEp7NtevzANmNguiuM9CqSacE55s0mfVQZvBA90mB/Sh3BNrUn7hWcmW8kIR3t4IrnNV
/a9aVjJ062noomhBYbYVPR3mPZYCwBwR5CdB/z+gvI8mCyVzQmuzGccV4uEYMpaN88C60kz7ADcg
b2VON4+gchxtmlatCxwQ4dVfyb2M6CCKuKZiutOs6dK0qgnQ+31466zHLDFekmjsVulNpQphu3tQ
QFS4+JQfMpKpIUcnNq900d/SeeGkcqhaVvHmOqkAG0NTFIVvzBcBNl99kfILxb7h66WowFJjFIYc
/adUK9j2yIvleb0p3fejIak7R+njEqb8U9PvCJBpFu+3FOVEFtf3KIJZzhzuqIb3FfSjxbRvF3V+
hPaAPK0iak8J2R45Iym89yMoB7tt94ZocC5a656Um2jIDhBZ7BpBhwY+RpHHgGEi+WObRKBzYtO3
sro/x01Ff0k5nhxlZeWxyBkh/2mFUMTuJrP/dDma0cv6z/TbdaZfmN9X4QalFIAIUSGmMQN+0ym4
4El7Q/1qrE794qceNpTY62i/90zE9eW5zAXYYZh9bWdoO50izgVSROp8PYe0n0XXjuRv1zN07OGT
WwhEMS37S2nDHNae/GBLiGVQGfJ2TIkqWFTOZ11Xj/HW7+p65d+FTgFTRGV4qV2cT90p3EGw/Dgo
+fV/8CUEt4FF229hkLefv2ei5j8LczNSrPpBkn7mGlGEEtXP7+oELYeYlIZT9uDePCd1GXv6+QNW
lnccous9dfDElW5wfsdjdoHbUG6yn1HudVi0xY+nXVs7taj9jnjaw3F+YLzQB79xOaftVPjzeCmz
smHjyo9jklwzLBXv3kFP9csAmZjSn2T3wtpmem8DkmRaBdhSiHlK2YjeExjVnL+zraGPFTVYb4h9
nPQeL+KuytkwDlO5toyUbDnNYWRgWc1RgAxUPJrEAGA2WzMLM1tgV0eI24A85FOagksnFodMPhHV
sushnxXbdZmc5WNbYgmA0O0XIrqYfvPdBYfuVJsPohTdnJj1OdwxZmQSO+VK8i0qoO8Jwmh2ygR/
LUDBNIbpihiETXvDD6JDTDyLNZCWstZW/jhn6/u/+eZF8ANte7TBKLIQlQp3oGJvkW/ozSNSCqxq
KSpVE0f/O2ykPlzrwKIk9n6cIuqWtZvPerb6sapYc/NZkyoAnhF9X+s6IVbttm2lhJRjeApmUEG1
JzJ8MC83Y/XS354SzZeaKv6c9pYLEsoXBIsZ2zfGgV88TGBl/T3fruiUTupBzua+SmFIVQZSDLiJ
vBi7AQ1UVzGdEKHNN6l00eJR6uS0SW1i3s3/7gfvP+oGfsNxajLJlTo2Ep2tHM119oEp+Vd9MKMy
GIrhaF7iGWjFUtypkVXwSoMElzwTbdhpjx/Rp2yuGCdulGFE6RxSwHeGBe2w2CQksjEnNVywcxl6
/zMbNatoFiZrmAHGHW+z7BUl0dIZMTBtgrf+zeq0Cuc5krJheuTzV2yKW2WgEEhPNlDMreJsTglS
D6LtM1H4dYRvsf5QJdmV0x3THJbsGpXPLOuE0rp6hyhuWcEJG4CsYcXaVGasut2R5LdLyJQ48Aue
C6/ILLlZRCUk9ENZAVZWzV8lpf19XA/5SX8BCinIlWoHxQka0mSJ2Fcmvp0+nXbxtDZKX/nW4g5q
9sphcSdHjSmy5XFsiIsMFa51ZMMgFIjodtnDImrO5iYmO6MyYlWRhd3oF/r031DZ+Ps/kiTr3hCp
HTDRPVpSwAOaUT2y47vXyarDFGDmXOdpteqA/k5T5+xUMnU1trECyEgbxacXILYzlwp+xWBvoEOO
qG/lzsxS3xbzNjH7rRelXxvpDPsz9Kho8m8bniu1Q+1TFg6OA7aBUZbEYriSyEp7vDvtECF60lwX
RhFhgyRu8tzeBzxFpkiVWg42Nx0EEx7o1dOCinjDkXwHY44OJmc2Bp8oeVlDXr6kpqAyxvIi9tH0
TtTf0+c/M5mzlR+w3m9Qr/djggm2bB2Je0U3zyFEiFrvnIg/cLmmWz8ilW+U4s00MurNDiqFYaXY
6qKBDDtZ9goRMmFqaS+OB1KOx10aVsL91+1vSlfVQMym18O/zbCAkhPFZdaDy74opkUf5P/JaaGb
v775tkrwfOIiHIO1IMhS9+ztR7uVID8h5590+m62LT/paxMe/bs8Twk7DkDoRKK9K7/O2H4ryeUo
3cBWO0Hz9Q7vYg9PIidtYfcoxcYSSlGo4RyYBz9KI6OhnIANGkyFiYX/7z0jxAMyVr1fFK4ncO67
Pftxue16LfobdK4UWBUfOrXuK+CQFiAH+ohC2JziCdzoA/RBdyubdJldRZWrJVHoWgSQGR2WNDGm
nVH8lWwCwRWZPUmy+e5Q7q8/OcPXLOTknMPjuU/3cpjOp2/jpKn756CeuW34Dn2pLINTclZAKnwW
bd0ig25jk9DhhCo8rn3s4BH3lX5GbLypgVe/lGA1CU3uqSeJ3TEf9lj/IDJqqXwwsLy0u14IkIY1
kVBvil/rxR51T9XRGULNUTGsB+rer9ZSdwdo5OPLZm45E+Ov6Lys15Wb/TnC1fY97qvK63QME9iZ
7zKiKGWjqTaClTW+Ge4WqeKRhC6G/cgauLgNGNM9vtmBeshmUOVKDZmBxUNRmx8Zyj4jrt5/Lmm4
qp1N9JtjUyyuPtOpW9tRav2CUH9D5vqS4GA5aW1Aana35yQlW3qPbQsZ84ji3oeCNbueijg95LXo
v/uroGcBT4k9LUPpVF7qDH9JbVeQWB5V0wtOUG5zE3bAR81A86KDlvwQSlhtTUjTDzuTdOlY2lbm
vQVUeXgVcV/Bc21R5/LaU8x6rKx4wLmCnIAd4j43EP1xZRK3troQlz3ezAambLag3CoG8fF/pQsB
3zE+Ze/YkYlZAKdmk7AqxO2AK4pacr/oaIzZHwtRJQDXSeliZlS3IilUY7xO3RMR3uV0yn2Whgud
3QcvadMNoYQI7nLmMh3W6uxdhXw6vcMbnFu1MXqQyjEsD4V1eM097kI9Mx+btZMJ6uMUsGkX9mtF
7Ls6l+M61eFyDz/J0rKLkA2docKR1Kk79prMXHSC5+UfZ7rOUYemKPyQZIv7wH1+8Mnz8tTN5Yx8
5rrwBlHJ/EMW2iMtjElKzvfSqkHbX28pae5fYEaq3XfetQgQxnUqdA1T7+PoFm0gNabtXpOVHhJ7
c84/eqdk38lxTIU43UIA9bNEW9PaLLF7XZSUhUhKDwLF4jt2WqV0arcp2+qh3u0IcUEDAiAuS9N0
sT0juak92PuPzFc5mXMV2K2rG0nm34x3iFjGuCEGHXEyG+oDFyYBxv9Ksc2yOh4K5DK6m9Ryz0nc
8N19HL0WrF/ZJvd9wnvIt6m63QhZMgrLvAh6Nalz4ChsL1xFm1TyxMECOC63Ztb2ANqVqtDduxUA
sNQZp3zX79AL+5Y2/GYjT+tZbbe25dHSgOw5OamVGJ9nSSlTLnz7JDnRrSfUHiUZQ4PajZDAqVWE
7r9IHpA8bS4qTtUSTfAunwOYQIZgVVAqozvlv1r0c6NQo37QxaQTVcCZcEEPaTTCJuai3Ywij20G
8Nks21k3fUIBa0wPWefp1qzJLLwoO23Lgq72OGWkYAfH8oJ9MzkybRi7iQnAaoK+6Me24tc03+5s
BR1hDcR/wh44Aumn5BlxaAyrQ8U6W0Ttb6HPB6Z0x8+ujH/0vGOO+lrUlETlkmnutkRiMa+lXbnh
zIRxrrN1nx3BlkJB0TnGcTYjf2cFJJrtDSNukAwdN0k+tBOo8A6YhppkMa1sgMTSxyv17O3Hrv13
zwADtu/qss+shUt3RG6cVQ94zVoijYZE/BO5IianQHdXCfjeUgQQJ7se4ehsWeo7frBw0qorqUbG
xEJjdsEzLlDJWfSz4oA/mKf3Z694nRNcV2rfr20mmC2z6Hz40a/nmi2EP3SOfPRc015W4GyQbwZ0
J2v0eA/GAmtFMngF5xEpdNMoc+1ZnZMdLe+ow6mn2inJQqitqfhVaLtsV1o8KnfrzMJy1u1QANyx
GsJom84EhU+CGK0oUUC4eDwBcnXmHUTbrAlWLxdULhWbzT52yEK+ZgiUkb9wjOLEMbHlp6hZcrBo
DLPYtUp8a36Jdu0dLG4Ziu6+2xvO54fnPorvHQKmAVD/6YKn3KJs8Jh67tdBbi3WZWNcdfN3X7NR
ekPNatcsKsNFaSi6agPgj7RPR0ku8pGXOJ4GSDDTfOo2093f5yDABgc8PdSea1NiVDb+S89TQz+w
8FI6nIsCxTZstS44bqrQV9zh/XxWtGJS59eBkOt7CSsTql7Xo0JMEQACAlymyYV9gt5cn9u3EWYA
JHdwfkcnLmfefbX8liB/S78qL4kivlCea+hJmz7oQjPfxGleP4A4GnQwIpj3VbQ13OZN64ChXZoV
opM1s5vmh7Gpzgsh2LKWQVzLrF6yb0q+m3d4h0CzoCV9wrD4FL6YWCDq4pEyRhQ+Ns8Cr7Z0DhY5
AXLS0v3xLOIEuEUqOIi+zf5/aryNrBcAyYnUkN1t5wEpYyCiItsnJE6WIMFtGYRmkrjok0hDjfEK
j2n/u0KAd8VkmIXnTozAS7G8LFmqiqhUp7ZEH9/xmLWzd6JssuvgOsBm4Oq/DbFhMOZ/kTC0ksTM
MdFsuF3qUgM0cxgZdZqgztYMZY3xmRmFaMVs2cg9JLpN5RiVVU1lJiiAthDjnt/73rADMKxgA3uX
RpMi37HfePgSt5l640mFftkLCuXU6qvfFEZbMydvKusw0N5BN3xLQIgNpQk9OWbAxprZuaGYDfoF
Tr2n/XevLszjeTiqfWPDKbgqO3o/JmmyWYEKC6AHILRe6IkshcMd282r7s5YbByk6dYGmIEEiR2B
Fnpj3UTX1fJh2aVjfrCW9N1DYdlxgMy5LbaGmzJk5grCvJYmmqhHX8yjgfVCIRCU/Zql7Mce9jXy
8habzaFuBdtGVS9MRaugvNzfUJxQ7Bf7zEw4iFfJYKQoiT4HVGoXb9f1hsXE+robxbc+dOtOP6Yj
/YWA/6araPuEHXlElklQU55ASAXasD+zYNrKOSyWMaf2UZNKV8EDhF+TpGE/PfeMkruMrfipDZ4f
hjzKWPmeQ0EYj/gpkOXLBiSZo0byrNOXKhKxlP+5CPUhBuptKOs/UhMeR39XVXQDexvwarP5QWG4
ckXRdJFSb7oZmxiH0BIH6b0Be6r6lTj2O5hqfa9/COt9aDFrSgi9S+Da9pXMJERZ/D1nB2jO+26i
Mmx0Uc+p/O3a+yRUQbI99IgPOYlUHL1W/bxnpiNWdDEGPMnEoNBC7E7lOLfX/USjqZZSTQmnk8UA
UT3LzbiHQIkLFNun4n7Z3jpN7ihe3Ynq7bScPlfpA6FjSGdGTtTfTH6I2kFcXz0Nlsytu8pUB8td
uIPU9QjJy4oSAp25gw9ICDSatvd607PuT+10pAV01nVw2KRW6M2ACjtjf0/2AEEQJ3WXdULS+uSb
1MuQ+Jw7uri1rI9DZ9KGqkniYklxsPuZYpu2pWeTePy899W6Vi+Bi2oMa9VLfz0YpSLGrWk+mIi8
z6Trmm3ylYjbMyQRgCtuHCMczmftw02ncWYKIaDUMeZvyQTm3Ecx7v7U5rhIAdiHvN5u6gk3t0+3
4txSt/W/j6lBc0CsiOppr0Qo6kttXhYJQ2lA9CDXb2KW7DiHi2DXQdmwVmXM1YVbFaGWlFZtjllH
EE+WOXb0Q61ARaoHf/QWJiWmGnbjC6BcXDQxBavg6K2bdWgtSCojoMjLDqVlQvn+doCfbsRTQiSD
0lvm4nJmOzo+Yn51M3b2BCdEXghFpfzEXapQHFMC1+BIbGpP6PrXtdmgBZ6g42FMzlKX0g9nbVpi
tiDtHT11NA8wNWBTsv9JN6IQUlGpOG6jUEFyREwfng6eoy/aeLa/ujuqe2fUmSp9wdm6drt+CmDc
pj6vmZD4iA7A9cqQUiiApWVCIpT2LczferDCKDTL7xdU8Y1n7KGIXuRcDqx3V1NXxrgQheYgN+Yf
0ZiKzEUk0Ma3UbMm8TKTOwbwcwiqOTvz+4cYGJqNKR5zAYByMc6ZNS2F76z847Lbp2CaQCsIQtBl
qeLVV8DWG4Dxg+tY0OxW+43cDEC8yzRQGPV6/zJSsRxd94R2Dc7D7FEF42aEHE9Ot23Ew9EuEQwE
zMlsLhJQUbA371n3LRUmcWnVQtoR46D84hINCc3DjREsQMKqd3dO6xFWzgpt5YmjD+iUoOr+T9ZF
SP79Jtr/OK7xZwH02BBCsqhlY26Drzb8ejP2GmXfyX9kvf/EVwbiFsCgS5woCfeX241gfJMSLY/m
KNc64nTbK7Lkjro2aNfEtyDUfu2yHRBRI6k0oZ+zEPWbOJ+79/yYvdmWyVZKPqiQiQrG4wJtACfx
F9Si4tkIuZRJa9C/bIgSiEPlQHAZ3W3SxHXe+efcvFjimhtR0GMNJngOYonv25Edb71dbiolEz1/
d9JO0yHsonoH/NxbMocAWfZFW23vQ8lfOx+gT58kFswy8F7jDDDCyRv6VvhiF35YJGZfQ8f33Xz5
Km7CxnM5+NgjqCgv+lQG9/7c9GgkFZviGiDvgtMZ7LgQxu/LE3OKJe5zG8NRDSR9Rh5tpXf4n3U3
NmGOl9BYYE1DojLTbxNzczprHFHfI4RogDzdf0xZklPvdJHrrjk0sVPFnu59eYXFWy+EPzjZABPD
NeK0c7rHDrnijfQgMRNW/y7nJc+mIw6p8eiKyrt6ROjvhyczHRpND5ETGMruZDR4U30+ZUT2iAdq
OjNEzNcw7e5Hi5wejn5ntwzNZM+Ql8+VBJVSVIUrEr8WMb8Uq/Zl8t16PXxJLRHZfZM92lhfJ2sP
ymTmr7jd4gNI/btllNt3Fzt4VznSFkiEAnDkxQh7cLlgFdnyAV2C7j/ubq8awU7iXzPeoGhBqixQ
ln2tRjSfe6GXP3Wei0acurDl4Axkew7Gt/ubBRmwGae3BXfSpmwuF5M8jRQ2NLIw4B0xlJBlXShI
wmkOnIVgB1DwQxhrls2BiQZ2YHYwhSwhA3thlXOpPxnQrJn7jBNscAmYN1bcFNrD9Ww6/S56k3TF
WPdOHrhLh4dOE8LFsNZA/as8aTbWjEojt10BfrMR1kFZSdPCBbmSV6hAk8tTfIeAsAx7SVUoOAru
IzBkqBdQuMhyz6RDOeWcpGLniij406Rn12uoaxa0wAimlf+z8Kyw+r6nnYAiajwmLPwQoNnrproG
7zxVTyK77tBxIUf1ap72bYKfP2TO3RsCPK1JefN33p5mHs6UmxR1RG3fL/98z+G+qK3U2yG3eWdp
EQ3S94whC3Agu8jKpAjMfwYcMCteFafmu/KlIUmQn04JCUtUbN5dYC95CXTCwXYPYQnUA0+bdmbu
HXVBoVXqxMlTlBUvJEi/U5kh6sXRyUU1bMN5uLDHvX31vVoHT+AmuMXPEohin/QNoZv/4dCcNg8l
UdI/Ylq8Hp3XEIcbp5AIzoomTXdypVHmmlb9xmqzTiDhm5cxxczDRpmUC6/LTrJXMNBWXnEvTW0i
ArP18tbZnVqMaa6uz3EIErxVUtWA+d2yIvUAznQCoRr+FIaK2us0OWcPvAv8CxbUWNJaLZyNm2e4
uCTpHEvHkFAW/1SzOAMP4On/xcGKM01DFQIN2deIgFHH/bBhj8j9yGKdUfT9rKKLV5r3NhvgKdtA
FFuNzXNi9hqwYq9pJV/ifxEHQX3xjyBbSqv81lXlDpcCP4Ujtnx31ixZ5NZtxwsvhG7N7fTVy/0z
soRFHnCgOZ8m/rdkpFMZJPYqhTTylL+tkis03cvQOu4/Z+xI/QZpcxjniKF+OSs9TLYjzcFOYSwy
gQ5ywDNR+trRhfHQdn0W1aaty9QE0sLKHm5EyBwp82XSB1OPWJK/Gx+jmfGuqAylFyipa+pxcOUD
pL+RdGP/ezV5XbSHh0gLpUWMZeeLy1HMoisFKGCL2yqOrbWxQBpuPRTvHb1omHMG0GMiQ0QjSLI8
SjZtPTj8/pP0ZyH2G1NLTxTtNBL0fleKl9LqUK0UdHXJpgETE9p8zrYVkDBOo8ekvL533N+u1uDK
M9p7cHDGH32Xr5G3wz1LXnQJO03iOjOWYUzS05bwpotzG4Ji95QRBe97bOL42dtyyG0/cqdWXMNv
aTtBNIZqWVybjKslwmXYdQyYK+fhljJhGuYzv+hDOpWJu30oKY/a+BKpWqLjKorSuRWIp8oQczWw
PIlxP2aFbZySBV+iQ6RLJTUwwvX254j85AFHPrkbnml3OVj9SDz/SAmNutd2DC2wGyw9hHy00StH
xVRnvlE8nLpZ8/jJU/BkUcUFUgDHD9UuoVL6fhVYBFrcmMvDDimWtvhCyQ5nJTvcqBj2Sv0lahBc
MCaX2NwLN+Xw8H6cV2+ASw4yj32b3o3isRtEVwroHY6Xg+7FnL3KnFEwmnbZCNBPYpuNp4OhTRpw
z/Sh8N/8ARAXsq+cLy+DwXOkVBCh88JNVH3ZOgAi21W6fUh/Burwffy8obY4iomjHP8XqQs+FHiI
/D9OJlYemOcXUYdqPrqFq6is6zbcQtFC3x7mBbfnmozkxpUdv6qFwOlhDZCtWzykwbTFLtllu/tz
hNqIA/MnMetTgZ7J8CsuJcg8Otcp4bCiymNcZurE0aZ3vowdf75zPY30k6lJtC18jjlkE9tqz4Bm
FdApd538NTKFsPkueDdf7QOGCUp7nWAcPU+IA/GhmUR2GTmYwCGLG6rnb7Rngk7pJ+Q2xBUMpKJ8
LLW1+8MieJToDxfSxOFJuENh7W+SBaguswHfYFb4wwkqx0128i2kepoJ+pbOffkQruby6SOx1Ce9
DaIlCq5hv+iscgohNw7myl+R9n9jPLmbkfcTzuSAh9sPe+aN4djpzVSXbi7Ei96U1jpz8+xUtctK
1juddnO2SDwftSK6vDYcCKmGXGhcEkm9XZLYc9dByJK7a1rWDVV8hlPxPxPkexqu9dK0+Xojm2UW
n6ZhtwgzSOGut9DsMZvFJSEiMMsGIG2m/ghWeKy5OqPHMUefnSbjGuKpIZ10otC/y5QD8M4/90is
eLU1oz6KwBAe3eN8HiSwxL9/qZXhMtoM5IIh8ui5srVzO7rgyBIJvSrMvEVfM4w/oAsJM5VQiKsm
DPkRe2+xv/aPsUwwHHBxSAraN47XWMDM/zoSRL55DzZctvdOzy0MWQUDtLmXl1tZ6idz+sT5a1HV
A2eayLF+yifvQRpHCbM2uk1PFoJhVEcvOuoVgP5lW0EdDr5R8iNcpQ2ZavWFwGk2nz4AhtYqCZsf
vPvFQJIC/6OLEJEu4YC+L6s/SkU7TAqG8RCCFCd3EMWU50F9qDILg1WMTbkv70YP6yCEwanjs0LJ
pi68qXZFwGaRNbsixkI5GJq1cMXa1yUNP5M9wr5e4jjn62kTF49eSGveSQl2j1upT9WBaFlaNwrp
uJarS6j2AZSCwq39NFiFSaNkA1RmXxdKLIUwd4gTs9kzt9j/xyndhw5PBwwPLah7bn9igFm1SEis
KXJPxjuzsOzsI5Vw78RoO275PNn8KCU9rWxChxCy+vQBx6PbK26vvq2Bwket6u5GP2YFzboh7pHs
IlPeh+qox37Gw9RqopmQwU7l13pNuf1/ueop0Ik69+6QxGeFqOGzfPjFfcG28A/ZN/2jFkIecqSI
XwxiCLf5dF6mLNGob1MH98my+PwQszSCyGB5JKE5WT98TXzKmnnKXUVQa0SFcQsF3wG/XmbmG3gQ
ck2QD140vtfbL1SYXUoEM0EO/4FD8yqW0gncOgr2yOwzFvH7TnBEATC11xXqtl9XCLxbMTF8/sr3
8kLpGJZpD548YMBTeR/Y1yjgeiIb6c9RcYwJOxmcpN2TiQ6HjUHE7XsfAO5mBAciSraTMCIoI/ij
/S0BPacIGH1jWZdUFFzdk9GNEreMkT4MwKsqoWHlQjK3dVbAeQZ3ptfbBZaBTSZuIpyD3FbfINeB
hUUyFWBhfleId2TVIesMhDHhC4qPtMLekwoAeXKUaeUge+uYEH+XSEoCgdWCAbHOgAzLddEmdu4X
FHh1/wXBiaQEUiB7d3SBepI34Wn8EahXPYrZBfNrDM0joI/kzv5TYx5raTuykuJ1p3PFGQelc2CS
0R2S4BqdVJpsXVbmsgoERSKRswfCkfI2qvtj/0zcteGPPeWxD6KNjPsTrm9EgQnjgEqcXhU8YtHC
vpfqJfP5l4+3dNodH3mKRIv+jLlVdoP0qyFg36ikDG/gXiizcXIQpa6CqYxyhYpOaP5YLkudAZuY
GzueHkh/O6lqoztzYxt8JGVpFviZ2m6q7R5cbWjYLYzeK/m3trkKo897adHdjDXW8ulGnikEnc5r
iPDAlEbbk88ET351MBj9p9PHwmD3MleAHYtaJLHcevLV8xzpNIDTaIuCuuda1vd4EDctowaXYdZ9
AEyFlyoGq0Db5aAulMHXZElZv3yG1mZ/y66zh/FWypkUDCha16kKfIP9abrF88F6Jw4R8bkSAPM4
7QTUHMv8PZ6F5UPtoLUOL/JwIgXTlyxrWxsP7Coedyto9n6hvBvHdnlFYlH1k/VEX449/9M1DFdo
F3b9FdMndjE4MmyWQlhKL6D8nrXf5CxZDuSTVPi0ZExa1jNXx8jWO+7Tj0NWlHXbiVQTNDzsoTS5
KJ/lGCjUoeogqEsYEVedRKu5gH/f1fJt1AhmA/rl+hinTgiFcP2gE27vQCi7zX5mUTxZExGhGDzT
ZdMaZO7FIUhl4buNvPhFNF4k+f7R9H9jr4zbf06QAQvQONH5v2wGgAW6Fx2BqTK+tDZWFbv6IDcD
fcFOjCxanFTvcb+b7I8jufhYabfL5nzTM4/YgagU5Jq7x4L+FwjHJZ7wkisDPsei3nfHufjA6BNi
BklzBJcYtr5N/ZZiMHUe3FmxQS6lZ1VZGfQuiA8oXYcYHsR4tcFj3Ie9xoIGuiQhvyvAIHYCP+GC
UnlpA+z+F7qkpAE4dH+ye+ZHdLd2FNF/8IYy092DrR4zT2UCKWvL6ntm+e2+kd8hebdCrbDjlLKh
AH2ilguubbtZGN4jdjj1OKqLF6BZm9+0WFzVVn5SQsPO9jyNPlq5V1YYuO1URxGj22E08cqiQ59v
zBLbNPqLEusObiS/jaOJ3BwGegUexPtrorMXL88WMHyDJbtj6KbiCH9IZhC9L5KeyHQ+9S6UdHoo
1iFAjwYJPrtBQqERF1LL7/YvymqlG2al8ICH4+W+ktrCRfUZpBWNBPWQX91EBBYN8eWpFNfoYHAd
JxEARvF3niSt8sGGgYOVYJ47D+AmM3IknKq3zVXtevc6mxJ2hhBrqxmCi2lh8pal2MW7ITcV0aRY
qBLj3FkKFiCaHYGsUBmTztvu/n1ZD2fdZFB/gP31QJgaPidOUhFlx1lzf05q9AROCvMEOQnj2sEQ
hTGP7v42g1tTvxXLthEaY7XAoxyUE9rc/BwJcYnxJVCy3Nn0NoBk1FAz9H6XNHsi4nRix0R1hjlJ
zPSqmgANickHoVDJ1JxQHwTCngLZva6UNUAd7z1VW7rrswzC3abXtuo/RjiMtpOjOjciijQqv/ts
v928azn3T4dBh8wE/eqJEBg9dSB1JC3FtMbi5ajISYRL0fxQk6nzU2/YDocChULlKfQH5ttPT0rY
iGdmqRtBieOvfofS/vlnTm1UF1YTxEp8hr7sdIJ+NkNZaWnTzG8xeqcTeYRq6hk6ppIEBSO3XVha
v6j3tWLLnHCErpzLMIXuk/5R7GwDSUWobUJhJ0VbtS2R+sfjHasw60D2tjOLZMRZQkSTEjq2CUt7
F4MrrML1+95w4yNrNEmMdp42VbneOl9hVGIct3cf//cwf1I9QUorIegmxWISShP5hLZ8tXIe3Y6B
MI3/P7HRf6F2QSOXH2+5n6xWXhYay6fm2dDnpinHIlztyORK3+aJZsuLKe1IK1/zvZZJTB3b2P73
gYrEG8r//d14F7rKHESRpiE43ir8PNNBOnA9SSqWpWc95HkBO1mdXVdTZKHZnyoteIL72QJAUQDt
xPkCFtR+DSmxmMGzgWTdhy7qrK2GYT/Suohybbue2Miy1stGkjKBLKhZ+vqJsaubEKFB78beKBlh
kUPLTu7U3jj7Ls5LDoD/BFtzlJ3eE4t8itxQaMBZ7dY+Q3IuBNppqfS80m6355ryU1iSC57yailb
XCVynR6T7txKxx8C6yloh80WAJwkwOmXswvhkng8j0MAKn03nSytTDGs3t7wtId1YHUUGE21hLdL
ql9z8Sv5NQw0raLfhZ2geSsERerGahauJmeMxtNXb8SIXSAWgZHBZkWFEg6i7h/i5EjKWC5wi5ND
4S/twZvUvpvN2TX6lV8Z+CQIHkcVVG8XzyxcQr0cNOHUaqHLF4ThiLnnASNGpEzeWjhnEcee4hJu
uerc8eHfvbmsheJMnTH1LN26z0CsKyvfH7r4T0Q7/fCOKemt8sa9RuQszCI4aiieXfsc+g22sPrZ
Et48fMTD8QpqpuZAP0kMcyki6UdqSLajwTu2ZLUiguVpi0+ioOGyWBVdpVa4S0tUI/UD1IloRJoz
hi9FpXx2oNCjILXRKmTJNeCUCOLWvz2KAV3LrhZVohwZwH7mJlIw9iMSBBHP8Gs0Us6dCdnXBhcX
chTMX+26nXSrQrHlYXy7CRzv1OuBbUMdNY9NlHL9auMIE8QHwl8oeG9hyPalQt4agLdWqrkh9u0p
kxZpCEqWDnvBng6Mlc1QEeTjZw9GPfOTW1Oa8aqmmI36lz2tmQcIaFiHarjYfrJ5mpTNiHVW+vDE
jX6Py2QrNYBUgFQjSWlBjZFubRJbCMZ5E1TI2hrhOWx2NJFS4rcp/7ByDX523IIqd8vmdSEKx/YT
ft+GJaF39kb05ZEWjq8G3CFDHzz5Y7Qzvs/punXBsmrrNkb9XI/XC4X0hoxrohimjetMyj6elQmj
EafE3uMEF0mzOuSa5fbxhNONVZCc7LhVL+4Y3pvYaXncEAY/G86K8682LbQ1V7heG5H77jet92HZ
ZeQrl59zgJdgzwgolRRJAEX1jAtW4glCxGVqWHkCa0tRwqJf/LX+EeSut34H2hkGAbL3Yq3PWs/0
SLx8aADH+o4W0mS8X90XzVCtc3JK5CqvucTk/qxK+Bebm4k/eN1gHRQsqoQsjKiwqt3hKkwGiW1X
MN3UoUwuLSemB87+/VkH6s7T0+0V4qgqxJoruWR8ynAMJJO6+cR+jfzyNK8FAZ6qLdSh7t3QBxvz
UwQsRY8ODHUhCtOS+WmRSmjY97v7dNyieJvPJSmidZ0NsookGglbUI4NIDrEVGsi1JAfhNDPm2+G
z8ToZwZQz5y8/K4+QfpGm4yKL6xU1zSVfKrRUy+YbV6YGevV/lP3eZoGJuYYirGQccvfyg7hh1CK
/WFOaBTi+9VM65pWaPq/5uwvBvbpjdIQChVFnC78Xy5xwpjQOxw3+EDtmZNJCRjOFY0V8j7A0fGo
eo/kmGQIeNYuo1KjxwOSlLU9ciykfr0UZKfMwD+n4eJfkWEhvJAS5G9SaBO8vFVE3JVewDAU0H5Y
HL7znTqD4gpeDGAQB8o+EbybWKD4WC36Maz9s0sxjLVVMha6JXO8UpLpddB4QgU3xY/Ma+goOxu/
NSpVsYxrxIHLbAzB2E37sUREuIog2FCh8EHdDqez7sLw7FMGOELpPepkzn/hA8oLH6AP0wJYw7rB
Oon8BMwvClMiztdesxK9VrPoG/Mwb7fSWV2RCvk9IZ4MgoD5+1fOOWw0vdepsBCste4pYMI9TENG
SZRBj62sq4KWdbXDQe/cXAPQxPDTAYI7RhZ2qBQIWgE8yKSkZKHODwqIaiVt5uQSYZh4spJ9RJZR
rtKjjZNPW5GqvB2YhXiAHU06abUPI7Xwk4XyTBmie939tVc3yh94GJnDIodIMI+b14lYiyWpSXfB
+yQf3TUvQ9GTep+eqiUh8iiSyY3GMG25QoOKz9g8smm5rldJa5nUdrbaRnfqJbQ+DrdPo/Np1JMa
SbTBXopXhT7Wd+wVRR7tIKwj0OJNPORDLCM2zNxYO6YHoSD2+utRS4G1kdNnDwMq7h/TV/RiP0qE
NhxtrQ2qta5m87Qlf+AqKgaSuvKY//Jvp1WD2KDTJAq+Isnj4TZ4EDSug0PtRPvKJJbAvqZYc0LN
QM+LP0+AsES92uk3yctUuKHmCYol4ys2CFJ4ARugrNfVOTOyUGNlazNhf3ggqGXeDCf8AyBEIOR1
pPLQfqsuN60qXHSFOuG8o22+DSn7ME6HHR84jj5vMd6LTfwtiVRjOOvAF2JTtrNsIJ3SkPYlG8rT
s4qKys2mRAZFnCqvMV/7kstvn0WtZ856rd//8AmzFtGJWveykmHga1g33qvYmvkVTVkV/LS21ZGo
AWU5m0I5jQ65ol4as17mnV3pq/BrVwnnP8FEXT7Y4XrYAGd3EIufXz629wuCEd0fOelTqsrAt0/C
7ChI513ur7k9kFplhqz8l/zNsL2zZsc3iroeMpkOdNG0/ogf023CanwlSywSb6xleoru0h7xPcBI
dYu3mqOtXBfQg+EmW38je/o3pT394/K1NBvWDepNgGW7z0uLLN5WNflKHzJnI0V2Z++WDIu50EvZ
NTUDWC6PyaQdAgcAjSSJsuIQQTSscP/5CUHQJs57uulSca5UtuNJeGMrpFwu/2RCYCMektdVFNBK
33a4CxRQaUqy+zhulQPAjuaZaRZX5FXlJ5cQkQ5P2zTQx1q2cHmyP1zAiy6OtvkDqaBMZTdE5ZJU
3inggzlegBSqUuKvikxGdy2oO6Agarhklba42OXgE05LRjJLWAw5I7tXoQjgIALs9Wnt86GM6u1C
AJ0C60ms82LjOVg7e5Lzd8EJ7bFoeGuRsYzcKjcFRbyGwKUtCmrIqW+Y2T/Lie2R64EovmGoEf87
XTi/fgdbUMiCXIcjzi2bpVulPixpMjUCf0+FjsGHmKdlWa8pF6CNLq+M2H9jFWoAthZKpT+QGUAo
2y13DzSO+VBiRhxqYdm9rJl8ZT51tuR0KtmRdLyHUBo2u8svPptt/4hlweuiN87K/D16hRx3SEjr
dIUMfnPP5FIh/H6MSq61zYEA0XU3iiiK52KD5AjpfSznp9QKEn72SLxm/o8um1KBCp8LjDvxoD48
6D0jub5Fnu0muwvKQG90KrDia6gZf00Yc+ZW3yo+Hamk4nB58aje7P0ISzr5GndfNekzOOnJq93H
tqBSD/HR1zhfbX6jZSxjAONmU4l+oTCVUycHeKC4tcC1XE8PVvb+HVpeaigalmZIHdHzaIE8RuPw
RVt8RTthh+bBGh7Bkz1wtRDHmcRyoMf4IkR4tGrsSVYaZwlqSewSp2hnIp7dbpfzmqJB8AmcykPr
oLAOmgsUpE9kvBBln10mLKijbsSPB42d6EzWnqMyxJdpM9CW6LVtgm3vE155tvQWZnOaDy1F/N30
rYKIq2HIvcSDhXazQljFyoDlOauidhlQCRhEfOr8XcRqEyEtBkIj2HiKeT7ktTC2feQJL0TCX46H
T0d7UcTl3T0CWUiBucoiVrZiFpyzfrAB8w6PrW6uNU/NjL5t3u1J/FYVOpppa+rQmp6gSJE7/F5+
aOmkiGGCb3q3mNYK1Cl3cIrJqOwdA//WdyiPwueJO8Ps8/2RZgqmcjPgiEUd6C42s7/MT+u1I+Kh
cBPUCQTvkv8/egoR8WK1rrx2Z4ywCqUhen/8Ne/1LoyF7XynfsAPF/ai67USMPNobUSIpxkHSCC3
yJH7gmEgGaw8aKGpFCcpK0pQF2p2IdGxINEnop/iLuJV80GXiBuV1jamHreXXsHJYH2pkjVVo3ZU
4tOHrD8P7WPktAkbyT66eDj1HzwnX5JbeEMKCbnZzE0zv1/LfFH41MSTMY2yoLnrgdHJ9IsRZTrA
d44Vq5vipvjhrgi08fbVj7vBMcjw9c2nopHfMGTXDFcT9Is+fETUiM1qh3TdCiRZEVuGSEeTpCXf
4LKklw8yDupIOxBWuZON56AToGNI2QBugXEHe28K8WrQLIIBgm+hdu0LYQTpS5zvBEvNCvspQonT
d07ePk4dx+bHSTj8sXisx67GB4s+F4rLY8SwDMHVdc/bFJYNL547G1T7R5c5pOPFlpC6J1ZVoLMI
bb2Elgmj80HcuhpCXHHIwz2wgkUKNLAf4Zb8Y9MlXOLYlTAqk7OUdGoJwEdWQZBF5bCwhszx8zfR
/R/OIkEPK5/Wq7j0ZtN4oOzqqzMr0CaLBeGnlHOhDWLaDOoii8Q/ad3Xnm54BDwcbKlUwHV3kX1x
53PKkuYGcply/Uhg4OMd/xEatOu1gsYyHEuoEiT/6bQL/YYz1Zq/TJhDsWmySmlexFT4pjYxjJwM
pJN/8xt5u8cMnVTwhkez3BwDwyP9cGsuDXVHsmgu7ruorVHkajxRgd0/Dp0CjboesApIEfKR5s3W
nUjk3SYOpEjtHOJpj3zKSasGxCt53pBjEoF8q6bUqMCnYpBbbODDiSPkcgfIhRMM5cOLugBk9hla
MesRsNReRVjbzqhnl9UX1DCb2vB0vvHjHZjys22rliFUlxxJAFZ52HXKdAsmQp8kmcGlFmyR3R/+
UhNMkiBLl9AWqiD1GkqPBvRRgtUF8D3gp9RdRB1t2tmTOHTlXug4lZUJk8wgNulTMMahvN5SvFkm
9jQlStwf0qw1F/ESuvt2XC2tC8CJXLVzkqF1o92KkmPuQurcnjwHwOvotU0QsLCqMNf3p/vDbkQ5
BhvjNilPI2N4HlW9iCQ8gTSFPB1YOVu5VL+M69lDmzew0PAq7aSo5spXnXTdhHscsaqXPgLbpk3f
nhjVW5YZpAKWlzlUYvJBNgcO654iVEUCEfHNTciJIQVopFAdiR2hbFysW/CnAMeu53TLi8Kmja2H
RDugH8rFGAQe7mgYYV4kJg3nOu+P91oMtP9DFsyz5mI2O3mNqiqClgIPja+0puhPwp9UX28S7Dfp
0x1T93AU00SxO3NfAX+fTbTnAFZaqLf8Bocm/kTpdC3nRH4tDkv5fucXnCQBaXM8/Fv5ZIt8GMmy
mtCvdMtq1KmEhvmuD0GgXI2qRoK0nqaM4xV0f+26P0YTYHrn6pBRjhoccnOogg+dQtwF03wXgTiy
i43dwJzwy63j/xQDYS2dXMwnQxNPHhKS7sM/3v56EbUN0k1Nr3YYDFZRhY2QcjLyj57QkGIPWbS5
mRo5vYOB10uQ+4gaG0w9pe57+eWX9Ldp1JRlGdTC2bI5cGgz4EVbOVnciwwBsDkCpSxWaFgQxpon
jj8lMozaETemlaIipbilBIjmvPTGFbSHQDqcnQ240nE4vx74owtxqpWdy/cMe57rSGawHN80B/AT
JicLZCckvaZGYngUZKejkfEKyd43z+I2eltw85sllSNAuoMCZMsmMViFT5t8pIWvlVPnkN2nWLrn
yipJ4S/waUUHTFHWTw9wHgPrkoypS1f4HWe3iIA4mKXBaQHhphhwIthdu7GdE4Dq9qSf2zsY1z6+
5JTOBgg2NBS0wE4pt8AjKxeFHltuAQirQS1X5bzURITVxAC3HKfaqyzJf3Ey/J2AxeAgtrnA1KLU
dzHSmw5yl0eWgJz1eK3Fz3vfJkXUz+QN+ihk7u5hQDrOI5bi57DiJn/x9FYbfHRqFGoql/UtCFz/
Pg/TgwBCQfirDtrhk4wJBc0vIYjXZj1/SFor74rRmnVyvAiQ+6jGlQo0aWESocIOErWmlGs65hxz
ejKf+rHc8g1Tde5YXni0KsrNvBhhB7RFYDEXYEhOSDo3MZnzWptxG4LXbuSlQ4/o4zmjnBM5GnFz
U9c+2nvrLLSCBPRhrWHUddfroctZImY91EpRoQ2n8IH6g9TZIIQvw80F8krMBULTCqphKavpYhoM
atMCfKMXBxHP09cwExeq5MjBHN/An6D+saf8VCT1K2UnksL6W1+J7nQQWWBGrr5W19tdeJoCq2b9
QdzTaXWBPET/TwQQfeX/Lmhf6f31zr8bzyE8krF7iVZ32TQOBCgmiqkZeo3z+UmpNeLp91lnA1Yl
8UoDNxlrGaRI3aaSEVdy7v5gWRF96kdEkY1ngwd35QMN1xdokX3NspTEq1hqEWZ2iYMLmeMoU7Ll
uOuGmWYVHA3q+XNE8BbgIe7qEFUFdnANKEWFwOZ2sHTRyY1jMHxHoFie9xtnvniXWpcLnmNKMM89
v2gTtbf8gfbQ6lrfEne5YZ6hP+P5qzTLJO+h55guzLiVdSRli8sAPdKTF591VybrQEOCn98GuzYS
l6jwmwF9eYTD81FeSkl0MRi8C5uvH9m4pqeOIWntrrzj07OwzwwksyPc8pbunBvPonsQB+12o7t0
O5124C/qth6/aIFV7LIVXcOw02oCDK9/PFEwPUIOCPr0Z9dNUnGnh9B4w874liFFoc+4BFQ74PaL
/dQ0/KtWVCw7vGAqwIxmYJHNQPvfhg1DSoV+SOPW/8Qh0h+bb9LUq23AvMYyBynAabLd6u6kQE+Y
pS6Qy/V4bzPJZbJMoaOB7C7KZXgeo4WKTa66Z7EvPN2HL09LV+5nauCPHaLl1QYo6IUq3jHZIIW6
XcqxuRcOqsNdKX0gBxRBXe9dKMw9uyiBNgD7I2lN8Y4Cv/mmJzZDHvkVvRsa2rnXgltHdzjkudB4
LzySax0NhT7QGtZQ5wUVnCQ/FnQ/DAxP2QX+Fy72Num6QrQVfLvQVdHCr79pW12aNNrFvhDlEEif
SU6RHwxfgvLhGjsrHg68sIayQEQkoGQHUfIvZlEvis3e3RslurZb9FyMRilR9NoJqjQBkFLlIafe
boCCwrPTLoQY6Zy32WTfj2BiWstzha8TuwHrqFFU5E1gfjEsgFX5tVcjbGq9CPBNieIAVCJkWcLJ
57+K0sd9K2laT3y+qv1/2J1mve/tu4XP5Zwk6ZQJub8eHPAj2yLYO8y0ArtMiEygmoNIWGHa8GsJ
h0v6WoLsnjJWCUKvVfm+cb2X/I1iuHwVqsYifZANaiMAkn5Jqq3bvXpBa9ui3MEe6EJdk9+ykK61
ODAl/pbsOVk1WM1pVDFXcrT2nVSkZclvBkE/fnBZKtprRYUyhCYdgz4S3YIBQG+j2DFR/s6Gr+0D
m2oPpUwMva9zUUwLgJVKWWOlafinV8DtnToOPE3tViinXHpiDk9BwOH6LvdQQcAuusnpNJv6u3wr
e9zpmoAzUFHnUSaWE/Q+Sn1cdO/8Ncw6BeAGNogUadF4gYya+bxbsUGI0BRw30Ap0hS7WXaZ91El
NFg5Q7Cmb6xDD7EUT3SPxn+agfqIe0WxlgKkuH++oXSbfqD4pR5uS4/JUjfjcTrl0I6nI7EcCMwW
3C33ef8UTBQuAB1UzHv62ftIEtAYlPAtAhycSZSmOgBu80VlaVqx2n0HMXeeTaZBQ0HQfCo6SqXm
gTWaICg+qhq70iYnUOQQIBmwqnnLVLtf5pjGVRlnJtkUw0/SWAb9zaWX/F+GpVn1Ool3jPeUZweY
WSFBjm9E1j6l0Z2GZ/vaJTdt61LgwnAvMLu9vvYVKllJIa/RITEsSvW6Q9CURncpXUHYZMcB4trT
5sxhGA5JgRFQbcNRevynK1kSb2OB+pSP20Amo1dZyap8QideR1uDhAoguoEzk9QEDlt9vYEwK65W
vvATG3yunde9RBLtXQVLKwppnrRvkUxX4J0hXwk1yYtCSjwg/UXiFWFWnlDlMzllJSluUWdU+RgD
oOXXjoJHlcSiBiCsnxC7fp1ANeiHm6x7rOXNGTWi16pyNEEdXU5d/MFV7EJTOOGYYUNvBXIzaBM5
HaCADQxLbFg0jBwmfcvagZX9RRpksgVhbFHjN0CId3CLturK7WSVGHd9Ao4o89iYbMEYeGZ3XXlR
HbQGG4S3osZ36i6cG6lQzl7xl+8rZQgPN7yHGXHFv1gIxRsNlYnFvZtjRGS9DAw2ApmLcOPT2qw1
pZ/OO8fQTGbpGsJmIw4ko9q7f9K0WfxC1BhADO10l8d3eskdpaJjJ2Fdtp67jryEMTmygR9iG1oU
QMYngjKqCyJRGVfydI1XhGv9B+oqJxVHBWKgaipHRpZq0vXkLhHjNj1t65hvhXHsSt/j6G9IEXqK
kctdzKRTpW7F9yDHcLPKVYjeOySSpbjzjJjUUSVxDZgNqhJWIS7zyqoWatVOqcUPKOuJ+H6/lse5
iQb7EpQCCh4inW7RS/j/yiTWCWEF7ezq7xlDQeXUDQd8Xz7kAn2aACETNH0rs/5N/UNMu3eifUHM
G6QRQF3fDTQuwp5sefyhoXRxs/Byr1Maeaz0otv+GEPZJVKhYOVnKMRnmC8QtDMSEJgpvewHk3sn
W5hoLwRssuU87cmD1EYF7kWSryskENJ1mj09eaG4t6r9slvJ/lBY7Setbv/jEzR+Zxf+oQfp0zxt
QNvz4nqzWZNcKJihaRHDhJFi45df1NAFTIQLjF6MIOLWoeO2iu6p1N0G5B3lhvHGTOMN/SzxmdYQ
bwUbQlIeFI4ZKfnTWUqhBHYkmRfH/baiz+0fPzZgNbZriqug5CJADHs2urYZdcaDs8Zd9yuM3rVS
7w1fPv+igQ+Youppi287EuWW/2DmfVB27t7k1Jtxe6uYpQ9BOm9U69UoyJ7kQQySN6245uV12Vcd
zCOjAhaPiW08uuGKylJF+oC/l+gbVWDlpyed6c2Evhl5shtaLRgkTU8wyvuJiFAI3VfYE6cRslK8
E5TAAYklMa5VqKfp1P2E6O7QAd3nRo0w9LM2t3a41IIqHpZWnIgEhX0/Ej/jY87g1Ix7ea9r4Vfp
/DegwxiiDe/FU3UW1bcg9DAt+p2PZvKfj7REQ8d8Ye+dzu5dv8gZ1k5o5bHUyhrmrKOPIuuDttGI
u6pClalckJHSVPy0zrpDjOn8DjSq5Q5NMBe+LoBNWTWOu9l8UGgAkWnQ6yE5YcM22EOrwzyJE9ci
qxXy5fYCFGB2n6vyrlKoz5NTK46NCovjoq+A/niWuIScTN92XnQWzOMezIcMkRDdsV1+dlb5uhB1
7JDDRZukijfty049phmY13o67iAHty8n+AbRwkBLpSrXKQ9jnKUX7DDGdZ6GKQbljvZyhDX6+xwq
oLmp5lGYbznOx+Tz9Zy3tB9BZJG87UZGlCD0UbpD8GRVYVOZTJMI9NloG57TnljBYaPPSwYFKPdB
HQduLShR0ug8RUGoEYoV0l6mszPznm7wt2RwV90b+my3+U26kU4cR8iBtZ/wbM9oebI67xofhxKU
CS/aTcqVDhQTk2+7gzwj3f2f8BMU8nato0wWKhUoP2ZhENewovp472gCzwcms2Wk4OVPNb69J7/r
WAQoT9YO9oNFYwnFaFlihHYpvyzhDpITh2RxfVFFSJc3ujB89vuM7hNPo9f7JHrrbPYNT/qD56YZ
VEEl9RR2GSLNmEmj2CcbyEwlc+D7GHw15FAMdFOp3bFHiQC0whJTa8GDIel+e2WKtLFeMkYsner/
Ap4AaDHAAhuc9wr3KJCQstU/RMKC2e/R7KN7vLoNg6fUZ827zya6MZqhhDqkB95Kbpdfb/XhHOmw
DQv7iNwP0nA9GQOSbwi13aTSKKYsibY+N6jH/yBwBjjxe9zfa/JGiQ5fwmb1voEU+uC6f/ruF1gt
LhJQtnohM/1thmHt/SvjSeIUxvA/jM8kCDd9Oo/GZWM4yu7n0a4q4PkWLTNcs1xqw7AfnG6NU5i5
bAagRj+Zh9M4wIzNjAYGrMtvVYPZHn36b2z0NFWR6MLgQTv//w3elde8kU5lju6u2wAhUXpmB1wB
xgCPhuxSn3QBJDvoWSP3syiFX3uq4pXycPiHq4CJh0Ob7e3qNKsHpyA55g+lS7He33oIhvQuoPs+
5MM6aYuOdg6U/iC29iCJijJUiYQU9Gf5w1lgESOfcVxVeLe05p8pcg/4m89ZyfUrRnl0MWiY5DUD
XsbYkJmdgD35YTe1TR/542MRlwhJM5vMWKGNzSpW2xK0CM3sR98ksHIhPNRIQKw/KgJXGdBZ8afE
2lVsRl5zcMfxtQ+y+7ko3wt2Ci06zPdKXli5BkDg0YGk9LAMcacZvx45eQ23kLz/Z64Q02GFVDFf
6XRSg3r/UYuzJ/bppntr2ROf2Y4BGjZLldSwufzG/m+o1kfLuBnuE707IKv+tsOo4V2W9uG04xmB
mqJZ0S95CfrGOc4OtC5unNoSZRuLFiVB1CSyUk2RaUzWJMt9AwgxETz1i9bilLrsPIrv8dpcEGfr
mfFVln6LMI26Q0JD4amfWdc/qKj5faGXWZengvTFBtPDDiEwniUJeBf4V6xv8Y/QfcMyE0Z1sbYL
3sRsOvKg59knhc7QmA79ZKINNguk6bw6oCzf0G/cXn9kVGkbUfRNlde9eJHAaGdhFLDcGcKlmIsM
A5slDwZ6mchF9CXoID3npx+mGFvstbdH7JHudMNxvmSkQLRhIxWjGqdQNHV1Dng3KbkbKvi35NyC
lWLAsAyMO7tHDrRRQ8Sj/Jfg/zgs8qxZY+GppsjnQIBpNa+vV+PDsxhetWkOPHbNfC4cPPB5UMMq
emWD+atS4ad63Vm8sV0cE2gIjiFca8BkF0WGbLM4GsyGAKe9rjDfFoc4/FPqhFeIBag908gxQAwT
FOdU0+HC3+RcHMMABD2BVpR46Rpqq6aWxZ7uo1rDCsGohbGvpnq6L9+5HjK1MLm595G3Ui3skpRN
81RF7n7QPhIxp6WqNMdnUzwCf8peWcagz2L+f4FhMIVpkMdWhCUg9yXo9OXnEU9S0g7E0Epcvzo1
XIoMZI1gHyr9O8u3aBp/Lo5HozHT1TYtuvSGkSX5CiYUetVsNlWOSA39seVgLYxHSGJ1CqNFnPaq
a+hMek9JayEYg1ybqQgem3ojtkCNQ0VPBwnmkpJ9NY+kztO34jb23D4qdIzFzZkYXxSDHIXm/aIa
byWvHrQkTd0hXeUlcRO3FAJrWut7dGHHpvxieR3+thou98xnQsHN38uTBCG9XGaZbU8cAgURC01y
5ppguOfQ8vT4PSBUyo5EjMmx7HzcDdOH/T4A7Cxj4YeUtUYekp+IzESBTjl5y1VzatIuRZbs31Zn
IoMYND5n1VKwQ34EWEno90usX0emYrMnCcFzQWU2oxNxAIyqZciK6zv7rzFmjbF+L9/Nvctybdy4
XvcqCqcO+2mipMhnylr/Lw9Acrz5qDlkGRkGB37nzzFKUC9hu6+/CY+Z9V2k0Q56i6Et31rV0OXG
Y9ACwZ2XMzLK8hl3hvlaZPqM8VxiK8nuyhGpOxoKst0/M+0/TIycj1yioKdfB4XeDcjdA29S9Hhf
CUD/ava9VkUPRpkmhVNIpF3rfBucgiqLeecSdSQ9XXtYGZzjJptZOpZKxZ/WHV+1wj9+WtRkb5FF
p7JJjHalmX+cZTJnx4hWwerFXAzT52t5EdGwELmiH41f5RID8mUl6y1v+uCUfVrEe/03GaIWS56d
YkajttQSI1wNRQdEK7xN6bkhVQlSo6HyPLLoNz1lx9Vv11hPnCYqopzDgBSPZQ3FUhXlbpNJptV2
aLupzSxSo+g0TzhI5ZM+G/N90VjSbGq8R1S9ord7yzh+cAMB0xpJS4ktLmz7s9PJ3IhiPwTZJKuL
Ng+bHTHorxxaLJWVQos1wfEDGnBMp0Cn9uAtoWba44ASgFyqyJOKJlurpU6FwOI2rZTC1z8655GY
uk+VVLygkMNc+xVeXCgVV8EDIUz8UREOMBJ/5vDc1Q2gkenxhMnlbFxQhyid8KDd+VbB0Nc2fd2S
yBki4ttQeEwjlkH5StOpzzVKBt2A3C/bmFXCqs0dkoVwPOIGzWkDcjjy4rQFXXfhdxJSiJsAx4vk
7jF2rEXSZR8WRrQsmsvuVsvJVE1y5k0wGYQOVEswxkH9yuPehuyUVlnoqU4Ey01pk/dohMMe0mMP
3zVnTKo8o/9THNdlz0eg+rZAE/RXifT5RCm4p8jCoXic1rY6HvI/ochFtflqEJDJ+s6C0vn01nA7
GKMDxJ+L6EHeSe3NiUpVXRckh7/koY5u6mARfSTLTthlTnEbG+d8uC7lYj/aR5xkhzNIXcldWt6s
f3Db9AV3P1hjLPbfEkMTK/ROC63Wi1MR0C3/rJXPQWcJw3LXBeXzuOWD7L89MlZd77rpANAW+S1e
hluWdIBnzv//CTgnR8lTdbyBQ9SZ8PZKkAnt+gI2kFrV7xy14nYpTshHkXh+jMsKKf+roeKsGTON
v3drwd50DwhQ+Aolunh/N8uKSrGeKgWtEXEvtt9JO3ORAbhRmM5mD8t8eNt7x5e0sbcDVIB7YDYf
lhZYHzdlDsVz/edQZ65+1ozDe7jvrJZB+FSyFXu1uv0w+wDYkDffjRHcRtCOeK9XfxAvjIED4ipa
JRHf7FSkgPQFrFw2TdMoOp6LCdGX2X2ou7qWqGtDS2GhTXNadbf6/8vM2WG3LI8dPflvxIEPQtDI
3BB7c6NHvevOryHc6RvzUYLw5P24+cIW2dE27MErSTVi/bRZzRX/0QEXPXjbov/zJt6+9m9p3Dvc
Z5s957q6rVjF9G3Upx5Ao6nwxx5cdIB5WegPbrkx4q1XYsodqSRVeNhHcAJVO/zZP/55wsHHKYuR
mMeCaCOA4NCek/XNvGcz2AnXPcdYAS9lwxKQHSVujCb2Y1JPRNeW5zWr6+xO2LB1GfSs8gQ/R2dY
UZRSinp/lol10tOPlD+YUx96pPE75qyBWu7CLrofrvWdy5aWuB9EKDQnzZsQoGiELzxhYngYZch+
9njnzzeXhLAnxi2NzaguX7kDE4xvLpMvXzK2LrDQiUZomJk0VZbTuUDpbrxSxKEkzUHMD0c2xRBd
nOcjREF+rlJgeP4zwujvcpeX7B1h7uAKlRH29qrWhi8ZHJPqfEx1T2EVf6BT5Hz8zQynYC5KLF+d
5Oz4N28CotQl8bt67BIwKu4Pr6qlWGtSduLjHOyJgsuCgpSidt1D0OYbTvfiV7fhO3CXGH5rOM8e
IMzT6yuicROnQreTdomYSwo7GL9yAmSGrpTDKXRRqF6Jj/5GBxB9k0za0SYoW5KRy3KIsW6V0JDt
rTnmMuXZ7XuGZUlCxQjg0j7b9mRrNVNk3oHHjZbV568SJ2a5KZiFtv4qCsoa5xn7lB8JOR+nM2em
I8VT60zr1zbNe9YikTzXqZikknxY5b0z+hKgQJa+VE9AUpyBhJeKrnKa/dRme8GRbC4CsNWbaLBX
Etu3IPgQc8KSk+rKBV8F8fiqDYqLdUDSDl6wrEx4Nrpj/R7kCUpw0/CNvC9hxzqk2hUnpVx6LTKG
NIte74fqan5gdMSKWj2L4GnGjYPPCY8lMOUejJSZYOJFk6kLp+ZbXp7Xp3i6ikoR6wsu3HojQXF9
yCsqfUO5VlS0fNP1iA+Ir6eJqTkhmT/pOOKJYKa+acP7YfPnf7bm6hbfy19Qrnlw3fzjedPGhJrs
a5Xo+eM2ID88G3kcpCHhG56cH8Y7s/LWsn1ttBIbNnuzONxdozrFDpxFT+weGGg8g/pVuUSUk+m6
9g6Z3sCdIKpOg72F1cEhBQ4F+g1Gyq+6FVLBpI68FiATe/ohMM+0EXlJh3mx0XW9/s2qWq2XQ9Dg
CFmbyTe6eXXyaLCiuYZ+np3SHqX5Qhwu6HoQoS1/BrALnNyjzbyZ+kyqIlGSHEGyC1e+cqw9C9k2
Po1YLe0u9bOLddjtPZMxPPT439ZHV5YM/W4/60tpPF5D8tvQ5aLNC7uuoqCCNd0zcNV80Hnjatyi
WSab1AV9n67IXSfmRVUZNFmYM3Lxg8p6vvM60Ez9M0gCHGZ/PGxjlWj1qL9JSVTecQbavDj8aiDZ
HXhN+N/YVnwyCBS0J8kOtK2kFqfn2FaGfU1uVkFqin+1V9bzHS7kKIinIMxeRMbTZs8G6XxWt4xH
eC+b2Czw9ZQQDHExK9Y4czXJKIMY3M/O3oHFrbaISUTfc+t/43FOJVVOWSZiCd9y6bNH3pCNPsBB
ECGNb6owRGjb6EDgKvE60Hitppb1m2vMHVxWaJTSQCTl0VkENo1ecjl4PSYyD/CYJwtv4KZO5ne/
dGoFs4XYQEflZ7luLHTjVTWjpLNEpLv7GYYDe4KIyWDL71rqtVTR8juxZ4lZ9XGmalR1FOZTkY7z
02oCnEeu+HOCVCM9j2YZcjbH4G73TiBS0+PRX1ecjxIpQztHsHm5Uqs7fMqejPjlDorEuZMMGpeX
a6J3vRwEADv1y9WVsfwGMuMDkSHRr+tO2SpTWKvsCaMWAgQqFQAuTkkWrbU6VKYn1bUSToOrp5bS
hjL0OgowUu1hsbUnNz+ChzFIZjxporILv0Qc1kdz1Ke2TCotJ+JHpyPtjwOumDoMFNnTqbw0WbyH
JTLD4n2pdwJVSGksQzPEN+RWORBnW19u5QcSKFOvICU1hUWhJrZaNAFG9vLMqu5eO3UMOnSghiGK
ZG2Dgp0aluU9WJW6ke10ummWi8QJE0+Rkq5pv86CvfQNDzfqUV0YEw9VSWyxCXLhauP7Zql6DK/v
fW+U/mArQlQxRWejkr1N+JJGWdkCSCjXOnS6Wxvr2T7tjABhZ+BnGxNu3zSct9N9XUlO6oJ/1dkU
LYpPkYxzpknXv071EXDFRVyc2XIEOALS7vYyt9IUjxrTD0BpqIejovY5nlgi+O8eygpZfXIJpi8U
/Nu0IkeXJoSiitx/YPQHStLXN45DCC3rWuEtcLlDLPCHKdu1iwTCN3iveuDl0H9MUamO/ZYRNxwI
GcE+QcbwJWNR2JSiJ1L2YZolpCs2YrVBz7WIAqj4SR7nUq76yyrrM7K4FeM7xpH87+34XDmNv4QR
w95h7P3fKSEaWIvrYeoJSrf+0R5CDo27cXJ9p8O6FXI2FNzsEHnCP8abaA31haRBoaPcZgeWQ4Wl
5mAzVovbNVtUWNLfBjoo3RiUq1LTrMdDP7qBjjmjRLEmhne0JEIPP2q9BWWnD0oTIadaUAhSMAdd
UYHHJSU+RtyPHlMLpw/l2WN/gbHwsDQ/AfXfQWCSkg+hKY9S8LGGs/eXY9dXC5KByQKOdtawM6V1
dVxFj+XNgOnP461v3w7yTKcjNWNw6u2eVbDlVMQkKE1lizAp58KuU+MVkMzPjCMyTKA9/Sp6Yvjq
0NcdDGam3/+S8ZNWpNCbgxri2X7M3wrsh9SaHkz5vVF1zagNBdJCUSyKfOuDtbPJCHhX994l3PHt
P24A96TJQsbu8EXeSpgnm2yeQmN3Z+/0z8wpBfmKjKcKduD61NFVmcPJYTc+fyucNurjUtXl+UyX
kJzC8/6GM9dffEph9qvgc1QeWLcauiRTO0VEQoSlNYugg7mZRQFdQDqYQWjtjSqANoCyp5TXWvaJ
e7oDwEFYGUTPT+/VjQUy2bOz+oMt+r+BlKfRX9FJBnZJSrlxVq/MVRYn7RXkEUsQhRd6itHKyQYs
B776WomXbFVunHqEQY/2mWfl3UvcLTOqbHt4u8DvSZgVyZBAhvsT9XEc2cV89YQKM0BOxXbIJJn/
sgylcl72XarqXDaDa8XfiZt0E3gel2tasIdQQLYn2F4R1AK69/Ny/3+DNS6PILJbuDNrDPZmPjvx
1VUEPORJ3W4JH9gqVibwCduyGoVCC2Z4rjlD3YLxzVRoP5XDThi3n0w3RUnuc87aCuodqeXxwocD
jbx8/uTbmZ4a59zbAPjL3PRSR1SWoGu+zAgKwfIk7rW7h+s4lA9LDbs2I2jvemQWI/mBICN0wKTc
pFtVdIa/alxdPlk6TyDMat8eTO5QPay9ou0ys/zdJTzSf6OZz5f/RNNCXjzat23usGRff34eHHNy
E0UzMaInM+oQuAxRDTfCMB6sUDf9d86DduaMnbiWw5ab3d3fUtuUZbkehjPxVte+d+ph/nvZuyVh
ZXZED87+CzMI7WYm3fJZzVtKBYZAvra3N+vXeLzWyFMrTuD2ozIsUbJNk79Kn/BMKy1+VF2OzVVw
JlRHYoLOC/qlUsPMFgYmgYXBAwfc+L6ng9CDCZ84UnB/+YfC3wo80fqWmAtPfpwx7yooDA31jqIO
JkCtxZJgQv1FITqRE1PYWntx65sMQlwewLj87zR0coxDNNXuW50TvpslIKYzNE3IAIbdPnEBQZs9
gAPdoqfr9fuyu1DejXYu/4fJP84XBCig94iOsdaRNBjvy5hBxcst8XgtugKwf2PVAQ5igmevxZBS
/T0eullUVXC3fJsVu1OTyvISqFm3yPAZZjRGmBCudi+61Bp/sMnKzCS+3l67RXtzgRGyaJhdgtY4
a8639r7FIsVxJ6f1rxpcrmytKPbDHiaDX6O2DylbOrr/y1LYfRsK110Wz+POUaGU9OOpyphzJHwO
de3K9L+PLefY+aBZR+GFk8g/LqpA4lWLE1n4+vvd1y3KJeG6cn/YSOdJkHrSXLfe8pvZ1jKaBJr6
Ox1IjH3s6bLUrrkGIblfpkPJnoPx2HKsBct9OTtCGszKoEwnTKQnaBYYEFidjVest7OR4oWSo7Hp
mTESyAXVYCtfXlHPP06LMwNE7coQI4MoTa8fBKKMqFj0DTAn9sniJCarcvu0Nexo4idUp7RvTe0C
gYkAviVYwQ5lGJDj0yFqDMut76/Zc2dffPxAWAuyl9AIeM76Y0l1kfGntbBcPIkpKEtMGIgSTu+I
Yp0etTUYV+Sv2cVj6nWT4yqvIaW0mPL1u/k9iFhP0oLwoDPAw5gv/12pX9mGudqJxmVaklCzs4J0
H46ehsDnzd6MM9bBdcADa10niiHpu/wNDUwQ1KicvyjGPTwt4SeZ8QDL529U07cxsAV0joGs6o4l
HwvDrF9UTXPbImy6UFfxtAhtMfBrmTY5eiTnpSM58PNNlF/+eIeiHK+39f0i84+DgXCGQtMKVUxa
Y7fqxI07ijVU1pLLJj4NSs9MggmIyLwRn1k/FD9Y0qVk9RE+bpiq3cSciQQ396nbez+sp1VCTVr/
5Fe8UYM1L4UpCAED89wMyj0sG7aZRfzI0aOAniNvx6B8KlPY198RlugO05QuMDyuNVWK+tbEBWsm
8rbrfw5TSoDov3eSAx1AMmqdfAXoK2NAp1/um2WuwygoPSVtudrsWxkarZgdaRfUUS9XA1DQl+El
PNegj8uVw3aGn2SuS4NWQc/2DeXHdJKe+W94ON6F2iuuCW3WxMimseiGbGUlQ/QZjINKTCcZdwJJ
Ej6jivt+9O1sYyYb9JAOGC/LjZDag7rdNKkKkzaVrW6kX8lMcUkO1AJxf7LNQBZu6vTltc7MuLeP
WUDOsz2AzsMfGkxhlXzHp3DJphv7U0ko/Q4l7z4i7kjWCtlg/adrLMZkPhjaVSwxVZJZimn/iZo6
u+QF9AibjBvMRIREBGEP/SMr0dwfqJYELV0V9UcgH2mSNs7hCUmDZPeuBc8mA97ZkaW7dRk8Fwcv
E2wpdGYpIJY1/RB2UpGCFFtexD62gz03vdM3lHRBClok6IR4ETvbuWzAzNr8X0+MNoCKqvQjIXIF
ngXoxKkpil8OqFx8al2t7IDHBdewDYoCtJb4qJbaPiNj0ZiGOKqg/wAUWd1ZA7rVQbSCbRqR/0KI
BDA28S34MzKNk/dvfFXCf5s7hNizwl/YbV2zNXCOEtyEFlx2Vtoq6m+H3agORZf4RBp+L6E84tJD
ZQQYYLTttbycI4G2hPGgv19oKaoNxxWPbmyjY70D0e0ncMwo771qTwOdG8LTH4hFeAwnK9mYZqhA
U76KM5KT9ho/0WKivvIXLOHCWB4L6UYZKhWN7O4FZ82NNQX3TFW6q3SatkDWCvgFUY+Cfc0L3Y6D
Yf+AgEf4AldnAigocj4JWt/KK/wTcUFKINX3i/AQeLIVCuATj0O9QlW4/qWH8ukdAGU+PqdhbewG
J77mTxfSwWcXc/O5E9zAvhEI+NxHdCl+dwiTCoNP9D4HxsADpGLjQAa2F6cdcKEcwLUNCQBm8OZV
9sZ1BdVYlnotn6aek4Ry5zMXhnWfzIJ1NG2zNnHDWT2v186UhrsdsC24iHd8DmRFuwUm/LOXKGCV
yGZ90fmnC1x7q+EJZ52M9VRRldzMrsL8YY1Kfx+9+wcSV5D1IJomiAYzAtfwz5n3Nth1KI24uHeI
wPGaDNpnBvRf9FeUWqKWDbbg/Mk3QIggeg4ikFExMQffvd5zj0ROajJ0F8KiFOqk59D/+8hfa4IK
AUV0u2aMZgvBSNfYZjagcDGRMiyO2MB9H4ftRNHergvUGzIsGEWINxm20bf7oJSAthdb692UNGL/
0ao8qqKFxrvnnqFSI5LZpsF1X6NL+agaTOZxRXEcH7Rk5JSKQSlFgdWcpycs4CnhVY3xtiG7AfXK
u7W+K8LfjrbDDZMKyFulmK5tyer07wVJpI1TjMOlHaRVmQn6s8oKLqpfVmT1C5E5FMf1NCc1DA/M
OeuNKgZKy2hCWQrHqwgKIyIy/0V03f9OboQ83492GiMs9bvZXcVMFHuCH6JtTKTRs16yvG/Rh9K3
DOzdBKsYxrQ0scRRg81fxslzjo3zEL1BwY+aOa0j9PIqz5HFssYPZz3MXaF0H+Xuy6qOo5gcUrkh
QiplGdO4S3DToO6U+Yld+KTakqemPeRngcqSMvpxzZg6jeuPMJDXCidFiAAk/xbLiQOeFJ7MHKUu
zwmkLv/aEAPxks/ZOtXUT2IDYwI/JEtgyfYcy7cvAHfhpPV7YnhaDxSWci+J21w7LPalFD9xgDL6
PWmI7YAFFTMxXZF6m+E6dzguTP/qeH7ePtX/7oLl12jlcxPbRcvkI9tsNbmNkxfsCjkUaWoA2znv
YD5q3AJq3+DxxyTYa5SEDlgGRi5MIHqmOUVnepuFOY8/PXtovCw5aUNb12oxFFYnAYJ5F0UggnD3
XQU3/NFaP4zSVScULs3x2IucvQZWh/iB0Yq1aa5UCFr1w5k5icPQKSTbACPP7IhPPj1FOjR40L28
OSjTCY75Mxv4fy331T6xhEIZw/oMukiCl9vdJajy+N7ZheQXmAXZJ0td2o2oeTEKlajiRPodGsOw
NkI58+JrM701QWmHaz7xlfOrocFS7XSbLU3r1iHr2kj/IfYq0UHG7L/2igq31Jj7kEZuQqs3yPfq
WNSATnXnU0yUOVQyXm/dvwVMORN68xRnIRZaxPntiiIWOtfQXWGR6dmByR0AjV7xgfAcXygbnGWG
pt/pUFFWXJTmQP5pU1u2umFRdMDq3UpR3zAh/5ohMHQexxo+NN5vNGfCPu+DZ0JKZgTNMjXyylUZ
qysGV0VmO21i0czJNUdhotFgV1eNpWKWD3GUVyO3l/dl6IkEFHVIUg0gKin/habRCfihUkcs8FPQ
0t7SjGwZEUjm56nPAsm2ozE1TGJ13IeQbDUvLAwc8dwbQyYT1u6BfCPbxIwWRRyB6TGfX6hZcxzu
Snv88ziLJArE77R9qGNQlajleniyO2h6EHlUNjX8yF+Zdk78VBY5pQaFleWThQyKPzDgLseDL9jr
JUEO8DhXgp66E8DFkP78f8CtOaNxgB0aIXuv6d2bWIzP6v0oNv0Qf/o2mrVNwJNTebh9M+CJuE91
AMB4PmwdITgDKfTwQTwbrUqX/goTjTfM50P3JFsO+Ffd0q17noxODc2XoCPZxcmwF+r7jR8xVM1D
MJICUGd6B24TiiZMKNjV7Yzj8Hww63WjZYkV9Yn4eP4lELgCu9k3VZEdxV74NgZ7/vtLEcocI//1
JMqyzn1jvsUCv+/rqHylHoomyozTku9ktjU5meLFIzmjhggKCW74g387gW/zQnPFN2lpaSYqDL4s
uC7Jm47eBukdtdOZ4Im8rrQBfmHarRoHKrSB3jEmMPxXCzPzdyKnLqrJGXg6alx1li8ZGAv662eY
5om+7o9eqX/NJF0T+Cztxh/sulfCSfDeafjLo4hhusYizLFvpn64IcsM0LQj2p1OCxKTdccu4x+Z
gHHSkx4YgrZ1SM2teN6j5nZSGWhp2QZ5CuJH2bKB1zHnz9J9fKjlu4/aR+aNepwbr6fd5eryLAlI
x3eI6KcNN2BXCyCzkmoICx27Iqgk/WEcdlhD4yv2oqGl+Z8NKw0sLlP3BtzonP//+US1xZzewpin
PT4S/ZXaqenzsxsFYw2dql7iKKXJiQsO3M7TO0zeFkj3CTqlv9+rVOEHjYfFyeQc8EIX8aoQmSWL
oXBbiigeLK/Gms1OKL2axMKTXOar1davcZLelh16Z5pZVGOw3nztQIWkVoSZE9VokYgPoBUbFJm0
71r7QKhUQsj0R3KHARuxCYOrXGiL1m4DSHvDCiKOtZqB6xDRgVPwoMVwuwTpsUyc8XABiX7Llq+7
c7FMUO2AUlXtIBv6WHZVlxAX/SyyDlfnB4lw+/7I8b9iac1AwQCZN+eMv7LLDSfkbGz6FYj0HY1r
QaqQ/cDSpgv1o3ohBkFZT4l7NWDEvmNHqLZCBRJeUHUoIpKPhzAdEgM89R1VK/sprX3u8yxKsZ29
7Srp9BCSSVFpHM/zXCptnywnT/M0kHtcpKlkiJRnBX0kede7RL6tvFQRUXWBdgUTZSufHRAJv9zB
5dXBqEUkV67aPsMaNE+FjGr1eRtLSCqUJaAyCcdLSRGEsybOvbefbY4MOUgbTDv7OBwy4C4ZOWPD
6NBk4rPEt1pEHvJUfzXjnV3s55sSgTJEgF19BNXc9qjbRJx4DrLAMtydSdDM+tQvRWkMwLhRhRkm
rXTpxfeucxEmgQnYjgaIvDfeLtUW6rJBwLJxJ7jDct7zkVoShpEOYHNy/hBwawLkW6GLG0l1l1id
0Mg5nf/NU5akhBgvpdsN4Zmxv4+0RsNxubMRI1V3TRqI2FshVaOzSa+r4y7x0q9TfpdtAMLWsMsQ
v3nlsB9sq8F+Cm7hGHoqQcgmCqTgnYsE1OpAx32MsdeEdcBAdSrke4quKr6HF4RllndQWpXoqHaX
/j/K8o757hNZtYwzRjv4tp4kPCDvYMzjarW9S2jwt3zuxPKzcHuWjFUmTHvdQyBZFzo1YyTFNhrA
v4iNrb0CSr1F+UwLp0pAqogZix5QMdjNxaxssDC/dDYkBeG3r5fmIPqqTgfoncIqONMCS0NksxYp
68+IcVQQ7Ie0EmQ3USyRBxCdl2QJo/Vk76TAsU6mqvW6Bz6fN6IX6c1bidEqGuMc1XGigIQBubJ9
YquIyRnYfSl70KhkZhKXvKgihib/0vqhgZ1x9I6jZF2KD2R2/gQIGUuXaUwiPcZVKucZi9lG73Lb
b6GoA3+3hPEbLiwGetPeMyjEuaISn6ql6jBGeqEMPuZUYiFqnOcm3q2A3MsIp4p1uzqtRiAoK2hW
1t7KoPP1cgGlGLRaV7MI4Xp/r+incA/pxTI5cCAhk7YGok6gbmaKHG6iEkhJRUElnzCDPCjeZBdh
Mpj/35m3F6051/gB/OKnGmda+eJnyDRwoTWH5c+mlWbN8u8JxYohgjKtAIMCbfMck1ulHQhegReP
IYEnTSxTAGuSe8Sl0ooXvA+Hv2HS8y4I77X+guTSR+6yQ+3SUp/N/JMpS2cqdNmnYTT/1DOAY1NH
VNNHqVtlzkGfs/xHjILG6C3xUpq0c+xa3nOXdzvBD6Mbu6ewl2aUcBAPKBNUNsuw7p1oKDiW8DZb
nlqZYB/Non2/xaWgcdvw6ZuHZOTuECkYoWmcLim/+O49FqsXczOuSS5w25extLsartPILUlY0brW
O0lITaSy0AIRxTGaConPYjSujgGFAJIonf41R+t3e4tdmbnjHM5VH5e6mp1qHjnFrZVPFvKLLEeq
DOWiqIIvs7mLKy0V1xghF0NWMA5420uZ1lZEZ/XvWFvI1+8N8Imws0RkO6CLe4RQCeL9x1e6pD9+
R3ZTrZBZRR/+QlGYp25GBbBBK/iszkn2La7OiA/SqN4/9EFynC35r9+R+RrCHBEuRLGKx9hthxBU
BmGbsRWM6a9bL4+h7AbMr1W6b8vcJqYIz8cRAVlUbywBVzj+06O/n4RlnQJgRngqkkQPj044pt8t
hPho4Gv5kENeNRisy2N5yUmjCI6pVp/LypWivlrmWB+dBOYMWpcSHv4v2uA+e1YAjBC9nqaheTeI
U0gy8R57o5gvfi7B6UlhP1is67DtXnGG0AnmY3SGkvtPfhfitX/G3Cu6gFaRoWK8fD4wn8Evk1VE
AM5zuHoR6YcSZ69K9YcrGp2FDZBqJtQUJtAbY5nU8DzHpfVebZoCQwy+35k81ky5Pigs/1TQ4lCc
9Z7uz9d8qYmEwNPR+1FXPSTyoZhyItNBS8CW+w5GsnJza0jIMDj27N0YQN9j6Tp6bjFLSMElff9M
Gi+o8gi3hpYx6W7ukgUfLBkmYGgqWf7zaP98BMDb7YIoWl5/uQo8Ps/rdCALHL//s5Pw0HXtxjj9
V6LYD7L2xd+uy28GTIpQvsZFsS3PPPOPBB1LScr7FWwE0CKo3x/Ji5SCH5Cc8+ilClkINqMvAfK8
2a5dTPwNEVs9NNXGAp6xnuFqqzpmO0E41/2yMSKbuUgcCdy4swR5F6/A1rfQjao7vugDOLEXYZC1
LXav7l+vKf5dRfXap9+pqq4wW5rdHzU/ZxpMQ7jCbtLDlub0Yp6bRztrojtEMhT5+J9ZVzksCmXb
iT7iphemA387QDwmCTHAo749fqFIDka4x3I+NGZCVOvAfZJNg5c61hEHgju/KqVYs8wSG/mgMYAg
LyznK694Tv2ZcPGzRIJ+rRxg7mthJQBYuf4G1DhCz5B4+EvE/YO+uqcq7jxBzq2TslXa9OGwVRif
VnrA4sQ8B3/QmdbuSuaMYw3HB8TM1lOihwHz9qx7DB1p/frOks/wRN6YaOR9ZEvemqVT7rRV9+Vu
7DIaGU4UaAkNRD0N4pp7u0sXOmY4uAFE/bRAz2XQY882CEux9Ez1tyy6oUx9CcNqbUMhoZiBjBui
z3RhWeHvtTj+Ocmsb/2cRrG83FCR/JhSmLING46T0vPaV5vQ5L30ISmfjHHd1ragSDF9B9jl9CGL
67xjY76bDiVK5yPsRC/P7FMe70wXObi0ilps/VVQTe3tWFMgjY68ri19/dtmfqAL6OTjDYTwLWMz
on/ZeK2xLAECnWk5jrTYfiUB1GOKRpyq/1Fk+lpMH2Irqjm04mbSwDMwlpVrfCafyvcblUZ5ZTn5
ZsbxacxZw82WpRmlD+AcOvOqkB3R88+Hh8lFovMVN6I3Mmp8JULbjQ1Zi9/eXEXB1a2T8zTjJjyG
JlbuQ8+7kPSN9FPVtmRXp40hzlEElEPiiMLaEhasfUOXir5qQZA5GBnLZ0MBIFGDViy91rH0nR34
7DQCxcQ4NcT+FKjMFlQ6acoxuqLnzvf+mWfXFfMXmGgq9yClBVnFid1GDgjumQHUcSktGZ/7T7Fr
np3CZDKlveW1hvwnyrFFc8MDD5W/I0N9wXzdR2v+FY95vIcZAl4yRP9O9GFEfa8dVCbG6aQrsjlW
CfYDkkftFn3b8JHc0MprVDWhrvwcw74zbSlf5T9f9JCv3Ya/tAxB7fd48AxHIiPJjZzi0uIbiqh/
uEkb2kowSFET5y4rHTzr48Jx0SG8B1GrPixOwOujNuAR0ijkDon3HgyatPumnY49mM217Nhi1W9p
s8oJV2DnBHZZRonWWswYW/ixMMHRTFXIGGAbqvfs9rj5DsSvl60rJ73YvdA4MdKq5L8Gy7IKAu4Z
wWgJas+T3wZIPmUoGN8PhWjuFZzoWaYvyktNFcLBK40gprH6m7ZgH8pLfI/QvTcIaDwzH52lJ1Yv
a5AJpkTinaBLzOwAtyCwk8QLlY1/nQ5LErQfvRNtsQ2YjdJ7Qv29Qjsha5WY5zXS76/TKT+9hVW2
dwS2XxgssG2w7qyS8mkIJfXnlo543N0TAz1IhzibkosqQBKpxhbsDQZPuv3oFHOGMZ8oIVVFKaFI
y0kIs8S11RNWHSf5JMIuX+OMs+mH8+AEikxtIMiUKkiGIP7HAq7fo2NIe03U0QfcDIAST6kgpyFE
BUf2u9NbzzqNPgJxHzod+5HmTJqh9TAe/g0rhUlq4oNJIZaD80XowWfGdPbeGVl33Sn/lvhK0tSm
Mbm5HjY/wZFdF3Wr9inbyhgC2sd7cMADS+WmtDCWllNo1NAUMgUkpM1oBIk5LQa2hj67aQ+bFAsY
UnNOFnaFM4BpWKJIcLuZ8s0mmhNNChhR1B8xg2zoNMgYI/WCTCP7CAsmuEtcSSA++vaaM1F6csMR
T3I5+CYLSVIvjgIpmltAXVx1gTKj0XHSzf4JxE5n4W1IT0uF5nD/MMa8G4z7j6HJ8q2OgAA8qp1E
tyNmRxmrp8+PUrwGpYUpK63v0p+yCAewxB1epCkc2JSNv7T9s8i1EK8ptDn0nTzfsxbnZLKDEe6v
Y4w+KbgFp6P6fwb5I5M94tKLBAD6F3CSi/C4XmVNdro5jxgu4WIMtNM6B8MiMRtucBmWzga9jHCn
0lrHXivArtykprmFxwwFCYOprpQQpd2II3qTovOJ06ksgiIjETsH+a8fVPm6amXpsq0uwpNJS4+s
6AfuppaFjoT9gjffCBIWfD263o7Na6uDtf1Sc1EOWDitcErJ6MAPiGcSq01Rk35ZcWvNkkoykA9g
/PJ+VxjhKoCNDSJoUCaRAy4K5H3jEKdeY8NRHF8td9uJEhOfHNscBDn9JFrfqRF8h0nja5e91sW3
cH4XSLVHfiq/lcspaux+3C/8Pmt/YH0h8SqJow27awSRhE6svWoTm6oRed0tQ3dosia79PYNKnUE
g4fhW9wqNDaTSnzuUjlcPqLYJ0qnk3cxLiKoYC1IZA4ahQg4IE51nAYdV/8HNzu65Jbv7OZM5x9C
VDYSpA6bkxZLuF/Wyx92J8efC+0PoS2mOsu/ZzCPQ43oOqLNh27YCDf8qS424+F4uFvaSF8qx/d1
W7+7sp1wFnDRl9o+nbfa8E//iZhlXMvliYfeKDSlL3TsHDgIDMnXYlZ6/WsKrP/tp2AXgng+TOgI
t2cn0T9wMiMsPH36Ew8TZO4GTjlkloEKyUF2gUjwS3VXKmUkxS5bUQSLUxJv5BMLNjhvS0dWZ+NB
erD2mAGx96EavdVqe2iazFY2Rb2K6bVJp0JVMui63wojT7GTT0hf/Z3Xikl7cwmVtw1YPR0ubz6+
m5frz5MKfcWGPHAOlqz8sqx+IMzpK2JnV4e5F8hOvWLVGgl4EPKxqUsfPYmymPZe9PM58xl+PIlH
9IzMVVErUX0xea+jocDSfLgMCHTKK8+fWB8rB1+I8iwUPv4ST9K+ylsLutmlaQax5a85jrSDXohC
SHBHMBzVtr8gA7PCwhZybtstGHv+QgYnvtpVCzesVFfcwPDsrori+lRylNANBoDtH3Lkvi6sh7+K
GGPMxOyKeDrI7MtVo7BGQLLg4r2qRZ/Spm/Bhl1cUF0cS0xAhFaHakT0fPfq5UNIzw2pg/d5TwUF
aiGdz1D9vw8s1YBotO0wXQCUpbhLGc2HQjv+mqMh9zL+t/xgQz4RI64aKfc6n4I9uo+gPstsVqO0
ThhdaA/2B+PTM5kupx1/TEJ3yI2M3Z6CfM/QD/66tJbLg2mQWiw8YEmvZkhydwx7Tm429RRp8+aa
5pXlo0WWerpk9mx+sdqJ1ULW9ZfVW+O+40YBw/3Pz2tJeueHGsOrgEALvmdfEHsgAk4Nygk/YHr8
f9oKhdliMhmK5clF9YQOadjhLMn9/iz8iRNtpQk9eBGXBzn2a7/RZUGHPeEGMeHSPzZKZWEQR1uZ
c802v+W3bhdqMCVR6XmgZ+wtiq3/Wo0aRSeQh5uJQRuOdOdUunTG8hK8xRXz5r8pqQRRUr1eAJ6a
UtU7Eo07scdTiCGvjDfVCrJxFgSyJR/r5BCdLEqojl2oRBOB17/zaPls0ajzzpDgrOPgTh0x9Mjs
O2nhp3cK5uHFhrwrePRlnFOm1xxBtqp8djyM9HcJP+fRqARKVlgJog/ZdLTWmrOVOCr18ZIJ84ih
ALtcUd8lWhGR8ovPzvH4Q4m1BJXSMl4DjXgp9rlx5N3w/LcHuYjzOcbsHZqyAo42afG2oYA1yCBD
oCYiWwlsKxR60bgoOAuNiO+1ni7ZIiW+92mVluhckwZ537pptZ7oMTB9uUTGCvxbzMOe3KNiyhDh
Dff3IftDBbwCvJLhX+NgwSqJCozVGw9+FVyerfXd0QJdOeT0W1kzItd4pKiSMOD7kVTm398Jo82c
UpDrvBq4mLXsEfscAu9x3ti+BLdmw/BXnOl6J/8ylU9rEt0Ya5YPHwHD74sl6Ze/BwxN/HS1+fJN
1unlxCKNBtl9kL3kU8I9iLUXR/xYJ48j88NuZOQAfSbctm9Bgd+4VhwOrVwnJAnM1O5kesjLfoqU
kGuHd/Xyu0duns2H2iyIzNDxWefmElIS4qHOQLUl9V9qoUbkY+jRCmXewcGyE26g4d4zu1E75LtL
4kTYP/ToylmUmvVXjZ5Rh5jhR8qfon/jvdByvkwkwZ4rSvowfCENv0v+uHhPUbfJviHqWi2g8N4V
Nf9oWb2PtBOIJBF+9vcDviRrtlyXT9yU3zrZxaF89chDejaXIGvExdGVTSITZzewq49vLQRhEzvj
7qLabzHsavBVvtzBZUqbUxSkXLHW3Jn1hJW6LLJHeMi7iqxhrA/m3woWFdX6CywB+hpwFoLtzuO3
JvbXjhEo/GEAHujR74gVzB/l+H6UTtFbGzMIHIxLvt8/yhe/iLVR9WaegLaRadG7N+ckzUXwTYs0
9Ihcey+Z7zqD4mDgpCrRqhfzilTYnR4nMZJ3ByI/ID+86rlMGWNkAfnrrLz81b4s+PC5t6j90QBz
y0eFeh4GetJvzIW/ZzrxXSIak6j4cvrRa7QWouTNkRiQy/dg92b2xefMoi7SsaV88S8idRc3Dl6z
UOBJNyOHUgJDJWRyB7koaP8UcoWSqgYKoZXgstGcFy7KGR658WJoXMHGclF8uwUzLyidhAsFstnb
UaNpyq9KKK7roTeLOJWiD7r44Xtg+2OXr8IGjzX0BVseYIj84wf9qaUEH6FHgZV0dBnNGZlyR5MS
/348RgZlU5IWu9pZKLtU2idZzZJgxUOMBtUqSrrxZig+LJF8Kcov4uQN3HMxu4zWPnWdGsrNg4Xm
MJRyplDD/ObSMErDZtoYRa79quMwo30KJzh+1mgLxtnKAPOMQR/5tG0vskOerqqNQU1mvSrREaJV
8A8l5qfbJiyd8YUbB+YNkmkvIOEya3Of0rLpKbl3EMSqUOmwwg0+l1fVjlYlXGoJvyd14bhHQvLA
sQtFi5ieYw6V37itzzvXIXBrmtZfgyz8zW4GeowekZPPFi0mWB2qIQdy3BKMCObU6LmvCBZqtacB
DNUlQPGqIuWPd0DyA/WD5OeZU5+JHXoUoE1jNORtwyToyTJ0CQSONudmCW1iK6sbvJU3J5diYGMl
FgvqFjT/J30ht85AsrStNG3RqVJdFblUzvvqk9Fi81//WdqF9+NkJx6qD+VO5ZMrksWBYgWJlAyq
QyoieUxxYRcfj0CjyaXlm4Z1V40NabaqYZVBJdesC6wMUtXsyXnlSvmPyfyyqsvJx+FltiihVUDu
1s7ynUkptGfmw1QsumKUwPVr6oKbOU0C5D2EarhzZmm71OCF2xnMnN+xRjI3Yo8S6BKPDx6lDOhz
Rqio60J7t9iRcPGyA2Mbm36QaSnrm3NClMqpcKx68JcR6/gF4fEFlUgwnDWoLaGJ3ZOOYOxQ0gSZ
5o2qER1vMSfnYtZ3ijAie7adaH6CXL3dAMby6Nu13SVTQHNsGWZPfLbDXeZVjr43Tg8t1J7JzEQh
XG/UmneHMvJXZWcjKxqJ77oiY6YWsUu6BrUUOBLen+kA8JJm1vYMF3GofG3fHyGHPmU6exyZX88X
Td6PwbLJxGLLJd3bCqEYNhCKqNELAW8IHU39ru99J+n8rYqLb88+vNYsjvCxJIhU/cYubkwKgfMP
q2V55VKActhqhDXSh5noUOZpnUm2zPxrpI7YFcDH5v3sQol8hu8rI5T0wWhwb/G6Q7ASaT/6yKZv
WW1XrFuM0lD54C2FF7mkSpJcfKmhi4s1+ziyMP385VcJzwUbiKwZFSiiP18UBR8R3XUmgLn/BF7e
6R6N3HuqVUbjonL6V8rVcX8dPwjPd7fNcpo1bnBecsi0DRZ078da469Q1yJA1T2+7obNhyOUObs9
RgdUCJVHyBJaMlB3NtG54VFH114P6N92S5ZZ5/v0oXybeFFHOMGL/af9jZsRJYv7E6i8uukAfDM1
W/zTKBsYf9DeeNlZr9MKsweXe6dHVRee664WFeB/jO6rOrHpsLiZ9XNW3+0vDm+dLEn8uA4Fq4Zd
/1HRxTpDUkNr8IqY3ztJs8MiOpoo1rd9S+wvvPDrQo49RtzuAJVhh5dhi+2n8lkx0u0L1mgfqd9Y
07UF82Wp48yysG66d+4DSrImiLKElctd00Zujd45R8DzrwbkKjQKJmBouDaMJQcaecaT3ns7QNrh
UiGBG3B/eGwbtbhbSLADFo4PtoMPzH7FwZHaKoruECVId7vLTh1bIKF5TNq3C+kbc4/g/Pp+U547
PYs5A7HJWuF861wtaZYt8v8OLx9y25uCHW0PGmApJz/5u60LRKKBZJVlH9GfnNMi1EXNCpck4JEE
wI4jNE+6itIohdTc0DdQVJ38rsISoPidh8ZyTyQXdKjiZon8qcMei4y4v0ldgBCTm6MnOCqRkr5N
0fLre+tIsQI05usYBPzxJgTJ4kzefqn60zE+R7kp1PtrDsp7IBvefOm63OvhICgBKR1YIWxjvarl
XAM1lcmqF4s1wGs/WPhKDlKO7Hz+HsZGuF3WeL4Enf2bE3FYn9pXVqPKJVUL+wY7rpJzETUPrvYJ
u4A2+dFufkfnuYBwidvNzDI9w7vD0vyVbH+Hpca5jSLXkF+8Luzr7NJpCoreJcAez06FUD2KFzc3
O9H7RDAPUfJARZJukgM6nM2p6a9ICRO9a7km7/EYmPv5Gt0EdCvSPlnfumkOqbg0TmtQkVG2PLBH
/8GHXHUSb65WvvwY+m2OPA1inzAUk5hqd/nId86RGRtZEQETDfMSgPb4S6LoIkGrKo6Ik/+E52UL
SA9fhDM2Kx7BHwq1JcyGVMGOZOnbUyQdqXJrS4/f+t6Zkgi5OE4Cr8YPCfv7xdL8IqzgAAXlCUCL
eraRSS533kG77UpSBcQ/6jeDEbC0BRUWQfQrYUqMAhXGnjQQhP3J43BKoctB2Sz1fRDvlhkR/O/k
p+8GRP9uJhzhVDX66OqFnztxv5QbL2ek0b7Rb7WwSSGJcl85gasnKMHo1++23Ql/i7kDL5IQLSZT
29wEYfMRyUU8Yqt9MOZfgcLHD/9tFQXcgJmq7KMbuztcgwf5mp9gkp7UzLxwLffKJX45WKo3EF4d
UiimzZbaI1MMxKuZaoldD2Qohx5QbHxIRZdaKxf5WJ6Q21TZtSNIVFBk20nfvOPOGmvssljEMGvT
zMLi1QabCpauaBpkeU/oJHvBqCXAYJdjHrz7rNo6193MVpu3FGag2KcrkKYISo+tup6eqCjnhUfz
ZqPkLMfzQdLQB7v03630Tlls0irHbhHA7jNAz9PYMyTmeDyrOfGJ61q7nS/Ue+7djF+nlB4NbLOt
tqekYMqoqceYDinNWGhO1uNKZ3PZYGONrow3PxWe0bQsxlBPqmZnEQuyHYq/XLfXVlzC2ki3kwno
menKXX2uaS2XjH9JWV8lE+bIXWkC39s8AEH7pOkEXG/SCItEoRSLv6s804PKuuCSAqefiAuyCCs/
QyBjCKwPDDMAeKIIgIRNWlPZp7JWwajiQqfchTWQve4o9XG64KDikEMWpwFCmHMOvBcwklFN2uKc
G3LyMHeQbNRPD1FHpyxP/At1ppPZ0dKHEjWmPMTDOauUzWbpwaUcw17gY5MjpuRXcVkYEVSfw23W
aSLXLHvLOpF6hga/xdhr/gjLJVaQYkQLaJuGOjAsg1/k0GR0EWdjFz0GMrDdqLmQhNRPiU4dv6yl
9am5dnAc9smkYMBlm1Y5Zk4+ToJl7YTAqOmEzZCztrGT7bSU0JJd4W3hVvKrDNBdgDbdVLhsCAOh
iuFsqCdxP5kUxrzpC45ZurW5f86FcLx2cn42kEK/KnXsjpmHEEQrRwfpL9XAB+IxkAAdiEcODqZX
BXpAltop5C2OoPyTVMsb57z0XVbIcXwtpK3NF6MfIWgW+VDiy8l9Fsjwf+S5rvmt37vyCiH21yBD
tL7S3HWCwmoLEWgLb04wgS0HDwkzT32wyORuM3lvn8VY1wwqez1z0nxdyovpDorC9vEnfyC+vqYn
i/C9aYntVW/3RdjThYTaaIOQflRh3bZ2bDUks6OGz3fWKxrF3KM6WOV/j8nLWjCbQqDjgR5ZGH2Z
5Vfrs2tGYTNLREbMrJJbj7sNCAnlZKkUcJl7y3722d4KVGmILEcYX1X0av/iSS6P9kp/Yp0tde36
EkXGZoupqUcSweUeiJkI8L0R+bNIdpFq7wLad/0pUYXW1inxg+NdQoz3cfIUXmWtDtEpoyHEq57a
xyEw16EFkI73vxbGFRF3BZxAL4RUsFLSEf4ej0ypda17bmvafe+svfCl6NHYGhXet4JgfPI67M7F
AuR375q1pXTkepGVMddCb3V0UUEKqRW4yNN6MZ2TIgBWbuVzxU3a7rFTFxRgsYiqBjomBA3lA4dI
pqfpsnjz1VluFAmltVseYnhXvuxNQMNW39BgiNmllIGhdP6Yh7j3XYaJ2CrVCMTe/RqcNiPfhTAn
/p0CODmQg8NT0Y+Hx+KHjDGd8SvWmoZrwmFtiF2iZgsvwRIDEzA05/sjvyHMMltkugVfoDOK0NIg
0sKMXTZCcrR2ezetso0SZwMaewdY/x0BuMqwAn8BjMzZUK0wM001OZeg/kxDKj5JjogML3QAutze
ISfh+n0XiPb05Mr29WORkuTsId+JdWrXS31Suv6FXM/2DSDcS3RpEAo/AfO9RqN+1lDeH8O0b46w
l8Rn8jJxaCDDKVLJhjoFFoDhTJ0Qwoh7ye6YT3PpeBc5+NnFIgcteTZCaHuWBIa/kiiHD++4nqh7
UAF1AOmFtDfojB9AXmJL9MAQ90LXjqLdAjw3pNdfr6tqAXcLu6eWE6Z++da897DxMWcXx6FCx6GU
FHwNb/0yu+oKmuci+dEKXeggTM+aPmfJZEvg3NMUQ5zEEFtuEP6+Mz0BmrbKjzYEFmGgTnlqySxP
ifDoXBd8F4m3Rit2OYaJ3nCrHJ0HzpLiQHnkNcMi+TJTnD3SbRMlh4jMwWRgZbJ2o3pkbkx+R1DR
l7aQf5Mtx+yh0DpCfeG2Cgi0hkgX7JV6pWNsr6E8MmTO2g+zWmP7VDGrSkuy960PDn39RJeRSBW7
X+00rM5Jp8wVgvf3RaythUV0GQvYc8lm4OVcGrt4oCl328IeePHckcdPyE19dbIYHJGVeRQLe30M
fMtZGptg7BExNBCMUDdmNqzrCaRMzN/9plyElACXkAHHIdqWd25ehUzyj67c3Zp+dqecPlrubfXr
TuAgXpdqYH4b7pwLuaWUa1Ek/yWpnwf2TjGbuwzKRQAbL1bvdn5TQCfPZ2vyavetCfn//okPQpEF
e+51+adXc1/RIgzSHdulwbEwUTZKsEvD5ot3A6QfWtm7T39mnugbQZOnVsX3IN0q6WectmDmY1Cv
hOKkHgjN/vSmQQ6ZVRYs6gDo4fpTAcIMkW29xqJG9+zu+fBGaaUHui6WyPsSVrgtLjYutN8Nn6eI
aws42n5H9MdB4370OKzOYs3tkfk8QJS3ijEQWLavIYzVe4WvVSPEKjlceSRqbb+8dVzRxg0AvDNJ
BXlRaJE9k1RWpGCToUarbvMPi4TaePStQPIz55rxN4adix7l3rzRFvoBPLxamp5TUGgZGs0QL3ux
JmqE/IUm2b0FqAvtOHcaCrumvYBhJU04GL3Rmv9lFZHu4nJaU0Ik4vgyqT7Bw7WbArcvTwsCmVz+
2l2cNTlgKDTUizfq9C8eukMGtDVZ1J5wNQCvXjp+gwtvHOBE/78Fvl3RiP3uh9CRP3JDPJKeQT59
XecxdfPfwUQsewAbHHuc2U3SRwUuZ5PriAQZiSN3R+cGJW+SdtBY/u9sfWxP5GBaE8G9gzXkoqdU
u+8ksFU2mFlnZ/yNziromW45l9TW8lHCRokvLrLeXc8HUr4O6CvPPX+FCNNHAMwjUG8vZsKvmI+a
LMQ0EDivkPsf6lyHkOS3ilZ+EyMTnfcAO3Ao26hkSdOvKmjAhXB77eHoG7ElHXSJ7eJvBXt63z8b
+rNp9CBTDl5TPz1KTo5DQ1U4zFZtJl3bU5QUIFGBlHyvqOwpB07L1oW41ZR8PUh441gHP+dwL8O/
lgYJzS1VgCjnZKK3eQyn4UlwK5EhDIFL1icXd7mSOKHzJMdxZ7MB+QDBfIKFfPU50g8v47ZzHbjr
swikwHGeKdmwoejB9xWEYqGV5tLuEVkP9kdELFcZCOFRrV+w/xAgd20jiyY+PPT2JsUeaZwoyrJf
oqa3N+xe1qNR8vbFXEFKc0LWpcS6zTbTWLhj7MMkZ14oKQ/JEt6WQ4FebByU6EtYTmJchfJNbzXT
o7JrBlpda/OxhPg+UiPAq8BWNo5oYQbezgVx1bMjDyPKrHGMmAkzOHKVAXP1WdJHFptoh7rwOFGX
L6lD+PmrXbJ6ooZt9GW4XsGXaZXfPzDIUBxIwaWfZwYyp54OkurSEp83VWJwyIykHuvUPmCluh9y
qcO/GwGDS+HBh1NYNMq7avGOr34TDHAWpVgaY1ptTrljKyWWH3Q7mrUhQqA8E8dPLChiS+3Einkf
lPb9bEkOHmPTszeHHorB+0pWI7CqdDfVt798oSfxHLP21Ge02cFuqdqPeDlPcEQ8QLldAMaP+HUe
qAOkwnS/oZ0+2Xzlo6jG/RCrUPOuuA8dH0B085djTyRJlEBB8jpwtpX536DYZ59GHbYoW3XMpdG3
ulVXgAufbYqeAOoH6cdtJOvkflXWz/kb8t8ApGOZjxg/YFf7d7ndyNYuYj8J2J7x9d3CMJGRZHX/
jwiqIed1hwKnRgr0Xrt00zLkk8XI9PDjVtApnzTn4XdTd1xYuX6oqozpYuTuU83umk2kshZdXsBg
hGBJM0j1fchfhNnilfDxAddzDtarD2WdWG07DiDEfiwrjn+LjWVk7xR/BO4xcM03G7qpwqOCg/ue
9Uo+B0GvMlfjYMbh0bxhzfD9qDwR0VPgb1eJKe26pqLVUL/it3wjKHkHvL5+zLdZAtD6u4IiR7mE
yQy62K3plL4P34iYio5QAPMtY4Zu/9F1eWC2VbtavlJkwTXAC2aRni3Uq/0aCgLD+a07TgHrOQfH
U8XuoTHtV4L8jPxAiKdT/nX+Ofkci26Ja3FTz4gC/mY6NGs6tgwg20fKZUH9/+XVISmoJdz6ei8G
Q6Aznvp7Mvi9QgxZwPMKhp8wpjLOfen1Rn7/nMfUUsWYI/w7yw1aSXaMOQOpVSo249l9WjyNwCOq
7hLQPx0mM1IUtiMz07AWfCyREX0bvomlAUgxhc7266IZLZoW2saej5B13xu2r5maZkd7n10XKZZw
tBTNc2C92z1qKKgIasnkf9UDxJ4iP+q1nogCKz9t0NXkkiOdBoeZc9Io57uAUbYbtK7X/PZbBknX
oEhbXjmryXmMu//RtVhMOjnjvn/vFK/oY9Oe/ZS5jTrUbkC6Qii19EkK47LWA/F00vWurv6TjxcD
Fi1fWw6zVURkSO76PpWXUeAaXxTuWFd9qcm8sc7ihUfv+eEqL5OC9tCGIui7wrMoy9edZ2xU16SZ
pPdvLgsBRGYMriSSFUTY7yYrB3dJXndle8wajmN3yM38FP8PdvH+g++/Xxv2/7GFrfoira8NoZVT
FVpP4i5+U+doXqRDbvTrYfJEa+/h78PUueW16+vn8EoiFfoAkJgLKmvYTbVMYkOVGawFAZdWW7Rb
3VcWJ7ZoLgi55hXwXC1yjuPIAxcWen1Jc5W8MKXDAWC7DoHiY/nSnje3PchnPLc5AfIcOAxFBwxj
nVrX0Lor7lbNSPIbaNGW2TL54d/Voij8BAS1qzIX7TZISTcI2LlP2KdoaVNXVO5xVzIL9ajDzxpz
nYw2++W/NzfjJ1Ftx1DzDE+8bL6OmFbFWjPog+8oZN08Rnod6LU4yfyIE6Qu2bWQt4tGltWjN5tZ
iISJ3HDFrEOFNiLUR5vVPQkJEBzE6Rq7KN7SzHrZyv7l5PajX7OuNvCyF3SRq85fNKU+TGmhjiSd
EYdwgFkxA31OJE3ktOY/4fklM8BYsgeeU5CrUj1kdTwWieoea4QE957BxvJhDEAK+Hvteo2Ywn3L
ly51UHuCwmLNyXK+LA+h4uAtaFt8QQVX3ZSkxY7hfCinopj4/Xy9MX/880mKtb7q2nDd9zg7XEFA
+n0UwefxrPk89A8Ee6MyhxOaBDD9bi30sUX6NnHYRwM6iBAE41IWtP342fOfrGxLmk5F2V746Ofb
rFPlg2MZT85w/5R/5n3MNs0TD9sXd6cmPCikWOq6WIpAhlTjSmIdg0M6Q0fEfsOn11HBP2Gud6CR
742QTw1a1x+vb1Y/CTq3H7uW5xPln7CEcoiP6ZboGG12BezwCEF26Peq5WlffhMQO44yhbVhv99c
4zXqzXgfgnKeVE21JxwT8QR/cQL+7o55hYbvCn/2txLR5Q5sWOCfLg+s3E6nhoz/JaTpNqIdRC46
GIG3G/+2sb34HUZJ5eNRMWWZonzTjMTtaOMv0sYfoA5o8PahAddbKkajnh+jgeY+xubSffZ3ZEHL
ZDqPC5A8ACtW5O16sTy8gvtynzCxjo38dNW3Uqu6Pv387mSMXtaHou7qAJSyaBsfUT4p0Cc1o736
E1F7VqACKyQQ9NiurYRmnU8j8pFSbwMxE2Q0viuK38eDBwHdMsWfq2Vs9FA4wAuCZiZGRA4/scZm
p8pbZ0+5XtlKxUycWwT5jyVvMYaPfHZT/UF6ORdPPwCNtIX1lqF9A/O6mEF9ZSts3zpdGAb2cIBX
t7OdWKCk1YS2wLcDW1Rln/JxCNAlxxIipXnsdsFlPlpC1aV+7CE/EBBsXEIKmkFDRfc2wHV83YeC
iwvrb5O3/9/1ek7XCYTbjSopLfB6v5M88/zcwnrdn5w/CkGfIUEK6VVX6f30/o133tlieXgr7TP8
XpNkiHPF79S2TOzs5OOUWvMGgUq7wpht94L7wTLDOjwExu9WgF6bOJWoGi0qhuEyYLEjeClugkuC
Z2ae+wrpn4d2XcFvHAPFrdZq4Yd8RrtO6MMvP56Forq3Z5KdgX9LcSWsjpLPp0ZPqDsGKTPbcdT0
oQRdDJ338qOpoAuIrkPOnCt3c5oC3uVYNFRUCIBD5YsCpCY/J0fkPYYNFiduXpwo7FimB22UGqDC
sT+THDUJMPLlwAHBPQApVHa3fIVhz4CCg8LMT7VK01aoBnaqE5OcC9/gOiEAvMEoeXrGGKEUXy5h
kOIS2xihUXO83+Oe/mCWaKafWWCNxyEIAlpHYHAU0oNntd5neOFMtooraAnvU4Jzh38fb1brKBqR
Cucvl4irDT030reNVbqvFvrXlVMwOrgAQRzF2jhPFRzgwgt+DZILf68sxsi+hI8cmoFP4PXtcv31
VCwyO/D/Bj3TNDCDZA5OppNBxcFfxMMm9Qa30zh4QtXhRor66eEW0rhXgMplIBQ1w10XekudaBga
VnEqu8lNpu/srujGZPxCU/dOUQA2UMVdEzx2bwEuwHqbG8QzhLiCmqjxn9QYNXoGkTw72aej9Fch
qkQPpvS23KKVX1YQkf7vivESEIQ14vpzXiu/FDg9BKHPAgOfH1KKbH3JWbbt/ANq/kZvqXEA+Q1e
iyxLgToV0r1Hb8OT/+wWBX1otv/eqgUAtCtJtd1CH1N60hW0VUXWwy44RghEhrVnROiInS6vTX35
9gVlgaTaoAREOfOrsMp+wyIOdg2idSokKZ2cmHiDAqMgu+57S0NWhbfxZ+4DVWGzS+BLaee+Wa8p
VXGtl/iAXxLwUQaHYy2Xy0GYRG+R8HNIZ07Rv0S66spq2bZ0iWgUWnik2xmPK2UHMKQt/uUCoExv
xlTGK2n267/yM/JE55b55cMk/MirSAaQYPB6jBQTMCSauz21DTswWpYix2KpTXfNX6h9OL+dPX+j
3dtfuDdxDn0GzVbWmZM719+xYonZEIUZnAe6SNIgn/JCFTfre+4vOX8b+qMilZNy1hWjnmzBmOeE
9HIThpvORRglCBrLmxsd/ylALrMEgBzDplz7FnOo3kPVl2N5WByp+pujhXvLin7k0Frl1RFaQHMl
HXM8Mrl64urXvcvQP6HTp8wmdNsFgx+wtrAesiD+z4ywG6rAq/9/3UO8tt5IGms8ue4o+xVFPSXo
ur2TwaEYStOAlWOOG90qt4grgr+hbwRMsOZnvI8MZK0u5rQQFAW0u89iteWCL4ktKyyi5whPxK7r
eD04UKqhim8UaHizSS+XXPIW6EFG6NAMmmNGzW3GnhxqwJtaflAPONtP4GCMA8/3yILqMF5J+Thb
sFyg4PvybY//P1UP10BX9Rhrrd0XH9CuDj6MdEb5PC0GqRT16Yp0bfQRtJhKVAZtIpw56C6Xvb9R
Bg0kMEvzdNwbwa+4wG6eMQMo9qUKjcXa47yRco6xsNvAwG8lVbF9ZN/wAZts3VFVrvejP1xm8kv9
b+cqan+vMAK2B17sVt1kcRWv8yPyGqBXSVOyu5f01u5GID2rcsu11xgMoypcAwwJz0+RetZ9IcDj
UwxtqZscEhtyXDEULvNJj/UNF3GWOrEyCCJyALyRabzzfVUXtJGXitfRJLPNQD8U9a3JkbNdQzvn
+6fKWZ0jqqj4ltJDS3blZNZKwUxJPzkSik59jHhXVBgPj4K/2oiff4h+tTbRne4awf20zkP7jaXr
aTtPmVVpHz+00jjC+6Sh7HPznNrBRxWNqufEYcWyzxYh6XqR/WvZ+/0JVEuEDzxoumwpYCPPhznW
i8TLvi/y59RegOP7hqx/rO5/YyGN6tQfvLnAqpeXTUvq+GDhVekLbCjYV0fUo89bicpTsHGEI9M3
qbH0BDieofbtOUf+b3vbf2Rn5myz6KHWTVUq7T9LpYSTb/zcJVgXP2n0+623XtPsgUgODTmMKEMo
BqPgZQkm4vw8Ksx282UzoKGjoEZjuPYbvzS8uh+mSTDzbC3gIQiF9yUf6LkcXsMSYgL6LkjrKwy5
rZis5DLlBXk9sH9uPN6bd4KMjTCVZJZQm7gCYViQeuYYBDU3afCIJ3O0XI4nfZfkdLEYv8EY87m3
608tlVuGswpPbnDyIE21bJbjFHDLYuH0R/jRAg2G6PqMggBGYtBH8sYluWI7s+uvXGG31ZaYlFi2
S5H40h5bZAMa56ogViYeBy+R7CkleP9OC/e8RTJeKp6W9vjkT6q3CBf5uLacL+1ftsrAQLxrw1Kp
YiZJWMP4jJd3ELY9w0bdRmSMjDz9cZqRcNUCxX/vzj41wT1hyXRiciWxfKBhDdr2FY1jGGM3o1Sd
DySfVLB345lKKnwtONqgCOFDrXvWC1GZEoKjEBzH8Dyn7lukgu3v9lgEXxzK8hN8eMw55yIZkT+C
XhmjIl/ZYX87rG/gOYtF6ztEWFrBKP3zrf0S2rkVVU1QQyUHKXD7sn4hbzGa7uIPQlAue2qRhDqu
+lIuwV2Qfv/N4/diI0yDbEFRiQvoCR3AfH/hWh+Iwf3ZkAGsmHbfc5XEHeRmUh0KoQQMlrIJTkKb
qDPOk63eHOFVRpTZ5K4yn92rIuC/t9CDTm8y/9rSnxgLWd+wrlv+kGv1bSVoObDnFrM3IKZDxmou
0jDf2khlsq2PiQm6503a0j9VWe2qXQGYVNEZF3FalwW1J71S331mOm6w07iCCZxshcUlPW891/SL
ZpqyPM4shGs6vzWIiwIJ5G+9DFjlVACTQVXHlOf1+7wgXtjzQXLQYA9WrsW5bEAkULVleSS/9zTy
c9KIXLwDQfXPS+88PrZJt6VOw04BiKOmKNJmCWDtNdNKtEmyyvHEg795jz0CvN2YrhGyCNs6OjjV
uTDmiVOAC7t0+1MSn2etWIfAygbH6j+8uC62KFY9pTpj12IcvuV8amVjuYOmCSvT3yXj5dJI/hfx
DafgIsVCfLpjyEBfb7jzi4vsSm06YEXlhWB45M8cta7wjgZPW2ekdun+jlqOqVf/aa+u30C9w4+4
vfObxNaQgPueKSMAnoUBopYussHYCeOIS+w1vqCG8Z25o6fzW+0/gE0nueZvzL9lDV/mhxj9AAIQ
xuZHpYvSBYML9IuonUOq4DRpi3TkT4xbjCJtxkKIfUmyAl3Gey+Wc90haDvyKL0Xp8bsD8TZegmI
XiNKkgibop+cff4iXuUX3pO0ZFJZXvMoXBHQ7OqFBh9EPSQN6iEuYvf2K2G4P8XhpoG6t++uKqlX
EOVCV1sv0ooo9tMqauVg9X0KjLw0BCo1BJx/90lAS3xfJ6hi33Cz8OMn1eVvE7wQQi4thPp8xdzG
cBh/JTdCPgoZHS/aG2Oc7oQHNztM2/dBhjgmZ43hEpqsVoj+Ncn00evQON9n+pKNhsq8EVtFeUU+
VomBnL77kMOQ3CI5qUTuqQJRjLky7vfWRl6BrYj/8t0HAlmRKSlDBrzMVpdHRIQ/bvVZQFpSlx9L
LMjvA4CjY0NhF47w4hfrbf1hP9PQRB6W8kxt1t2jETHpqMZv6zzsxmuC27zjn473Qif0KUPuxDJ3
hGByQzE5HoKbsWhf2zN86NlbJ9edCvHUOQA+8iLnqo1LHfvUeheGdVP7UWUBpZKTmv+IEkCFAb38
/8EdbezLqu6RGbm+8KP6OuLdth3HuWjv5o43HKKe1u9yH71rKrXGD2IzlrI2PLiw+24Ca7XCiGKH
Esf+crj/sACNUvQFq0X7nIJhfOlVqheYI99uzqf46+WAVsQbDhUREe3wHnih45ZgNzu7hUcw372A
oKsPg83NlPYyCo2PsiR5JnfoArdhQiPf6ut/XZkPq+qPfVrsieb7MI62SoGxAaSlqWXF6EthUnXG
5ZIYAMdVsYBBYqrh80a1UUtnZml+PPSp4YYmgjR2xrqeK9z2L8a7kHHFw8zRaDkqH/5ytVPuoX1r
98JbbWtcGmdhBb2QcTY9g/6wWdrGGwhv8p0RrFAiG8+puGXjnJ0eKaKIduMWiRgA1vfIjxIiky+9
vNr/tVJLv8JZys8kINEvRk/sSA7aIs8TulF4SABTId3ibYrWknaXaBFsNYtqZLaW70tk/c3S8Nvt
hPOwF9000XUGAgMYHZz2CtZFoSh/E3IyzfRTAMX2DucIAf5rFlEo3QgePC+zORNNfypKr3HaSHqc
pcZVh6YSXwc0OV0K/Y4mUkpaGeq+pEiz25mBBJghuK4cldjrk30wR0aqAvzFZtcbNd97t29kmQCC
3vhZq2iqAgt5kpWE20pdAVZfV9XGMzbZIHpXFUyRDwBuXkdmSu0Awj0JEtMNncbexk+AxlpJAovi
uKVk/V5NK71diDkrYRzkqR2BsB9szG+tOob2yjX1EtmTePjaa8Iq8Fowz1Ez/L5GiHulAPszaSon
pnAbzm0fsnSW4PHH16g0DFxHd3DEc8X3nCumVU6HQ7tB8F22cBVP5lIF3NTA68vTGoCv1rB6VTlv
DRVYQVNdEUXURhlMsRLwh3FtuXm40AVkOeLFtp6h/mIsQAJgJFTJChxgN3B94ukglqgEcMPJi9Gd
6rUW9dFpjBHHy7u5T9zeTyVqkbt/tqFz7FFfKLb1zLRMRsnwOc7BWKpymon23frW6LgSF1clgTMF
xnqOl9AZbxU0aAY33Vnox1Xs29XsOQ6vbUxm3fAxdR0d1OKePGunncJR5YhzdzFHlauyV8w+a54R
rweW41GLBeKiC5p/HN76FBYMeSU7FKcYcylc1Af9WvJebI3PsKiEOX+Ine5lU8RVncqqrRb57nS9
IsP2hKaDgL7JG/VyoSXLuQZIuJe7Jm0gqfutMmREq5UPIJP2lIe2qftWXa7tY8cIeMnfvOEK3b2H
3uTVkQdCylFS2jiTyrpGuWOazZMnb56JvPGbUb6zvt+4WJcJGfgYwCCHK593NEZE/Jqo2vD11rGq
ni1sqz4HWhYASYOziqLZpVN2NXbHGzCSc3apcXsMEMPHv2IDYJ4EXNiPZRF6ZwiZyiegUseIKQrI
iKSZPk4G3V2TOLobTynnHJXoClBwQefsqERL+OQifdRnjyaYWi79TnN89Xjh5G+A/WyrmTMhaImm
bgUY3podtp9v93BvOoosUsQEUm/u+A+u1KNOGsVKYY7Y8oc5ZZHo2U/IlhYoZpKoaLG8R4O7iRo0
u+oF0MgCdzGBiANKeagg9q5JHq3iNIifghAgJOHoepreEL2BVHMbZ2letZM+wwH/u2XmnkrLNJu1
MaPg07WloEB5g0HJEEjitDkYWTLPWuoI5ngj8vjB4gecGMYIz8dHmtJDxLHH9XkEa6DMIxeQ7REt
IiYf4DVYQ2VtzqkMcz4oU56WOUY20kKUz/ZuwUevNeZR2MxUO5p8+FW0o4Giekca9B1ZjNvzSE49
UUkP62TTuC7FojnCOhnnvqiGbRpZdptHqify86dRENgWbcITIG0e+Wv6Z21vMRths/Xz0cH8mmzH
70P4B40xIJY0YMxvEKgUI5sWVKSekv5lTippYywYjVvzx1WuY+P5EdSAQWNkLH3Zzzjrqy91xkz1
10Ospw5/rlyfdrbOtwc8d4h0ql/bspCV3WKhYjjRORWLwxb3tWUxwDxnyq5+1hICVwejbI/d+Nnn
VgA/65m4JGjymKKRkYJxI0KA85PD7k7d/Rz4U7xGcGuIQ96kD2JF9KN2Yp/CUNzfHP2CjrekFutt
Pn5n0eHjVl6Idsx5jGPs5yyO07EAiIImo7NY4SoU7ifoAo+B9PWqVh0EZRSHr+evghNHbs7nTKJx
eKESfNZJHLwkExB2dtkmfLJgXjdb4k/WW5x6ghmsEnWkiEzlz5saKzYpydfu4I6ziMakmscJS6Dh
TeE2axiGddGEIyupP+BzYJAdu5MqIov/sE5Pv2oGVSbH/mE1z0QQ0UI8HxC0F6whx1v4KJXXN6XF
btnha31gf8FlN2GTEcecmLN2bfNFPbZdiww94mO8y0pZUCYKkOrq641hrIiMrXO94jY5W5AMP0pG
AFtw1OKjUKs6DzzTaWYknBLAGwLNsVkj4ZNeUs4re1DnLkKry+k0wyNitgduFmBZsJ+ncVGWy4kk
wuxyhZCZ+aJFj8+Sdk4qkUet3Cwmw6KRt4ZOGOztTW8Vw1yvnshr5ii4W06lY16hQXt55QzOXCDk
o7kP2LLwU8zX6o4hU8EO9D8md2f0vMP1/KEUgRiEp60eyBrf/ZpWMswtr/uFieisIypPg4Aqkla/
AKx/Bd3KQNTK8JBshc+cwQmr63ySA+k4govyogaaHZPYW/1GBFple6IdbjQnyiCttqxwADQelpQD
YAmqQMsbgfq8ZqCZ+quUPBKAmztwcHv3YOoLVrl+qf9CcKdjn+chpWpAYcSSNk5r8WH2o2E0J70l
24GFNR8oZEaqwQhMvYAXzXGJY+215Fx4s7vBbmBqQElANyI6/IkujSzbivIS0W2WuQpS4Ag4c6x2
JnhzDakJ7l4xX18U65Go/2V2mxCXwqoNgAvEHUvDhKuhNScF1Sa2x8okTKaltldap5OWD3tqI36q
L3+Lc7HCXkiyoyAqnCEu2qg0/Gd7iikI6N+i+fdiSKLWk1cRFdz6kI+3nr5G2AtBwWx8FlCie11C
unQD3ABpMSsXDtBV4Da3tZFbLz4yIUjfe+QAdYX/zGZLxTjLKM/AAKrV5s8Fo79gJQDGsqwlkEma
iOSrT9S5qt8EyItdPUguf5cZcthjXtDZwvqeidIw6TK9tKAK6uerpyeJr7Tf8Fb80JmwXFurZQxV
ne6ZqbIdcmVv/vGtaPjAZRPV2AEIGUL+/VY+QIlEFViONL93vQlJD+i1JYDgSh0jiO3zL/ffMQsk
wIO4xPQ1smMsYMzloD2Otgnbu4MUcgHsPRYqZ9zNm3uRB9reGDWxYPidNXqdoOKisQaf5C1tNymd
H9hJlqFmiKLPOqTy9B45RiFvLV8Az63604FWL75tIeVMmThnBcSMGm8oA5ptMXT6HIpazyLI2e+i
84bCtNIdcMc0U+0OviiNkDaJZ1K+9kDWdCDuDQONBd+9xzZMAOuP5lb2oyMiGmYqssxscfw/dUqy
HHrcfuoz8oXqk6SCLBY4BGEHTM6PYg12tOM2koOdFTKaVAWycH0T9ogXto+NbUM4nhU+5fZaShhO
vYONAnGqo3EgrDyG5HUM2yX+c5sHuSC+qExHuqtn5GeqWXyKlQbG3GbR82K+3C98NQ+LgNvByzOv
/RDTv+SpNKJxufcICzpSu37tVjp40fHICOJMQeTe9XIcC1uTN2zzg03lE27rMuDtFyJhV/N0GS10
WEOd9R+f+Bkaemd+P4TQYbkmoBL92Zjs678FmNEepuANvsKQZiBYoj/fvKhF38+YbForxAzJn5Cl
iS9bVp7wztlQdu2aIGBoKAaAw9Gil/eoS4AKV7ec+ejb4wY6uxuh5Pf9xLu+l3oNZPSh1rPimZ2n
pWGuKx5VIYjPHr0/+A9SjN0cm79COdGB/5Yu5iFO1lPvKLFDK8OF4jvhFM8VIYlyjsdHxmPpCQW7
RvSNr5GHp5fM2WlrPTKNwfkKTyPuifYUzygRJD+FNqlbEvQUx1/B0vAx3ao3pE3f2Cg6+BqPAAR3
n5MHs7HP5B5+TwqgdN0+AfjtDJ8/LarzYbKlFnrEfV9OipwiKMX9xEqw5yOLYy7cDdD2gUHPirY7
iUdW5Esu01Jl+jnVWttqkBuXEzbfHS7h/SnLMmOxHoahomsH2uOZeaprrrZnOB2Ph5wmBypdOMhO
jvTbbmVXjTM0UK5JmDTo1tJAadr9U4NnJJXxyns8kjNTPrtnIm7wGG1FfUvzh7O/ktpiDpkU312z
di8E8MLuv5Oip/IO0TvNY3Wl+RxANOtnvIq4TA4rd//egiQnzIz8W97JWbjwJMt5Ync+GoOHMeLL
jxBxe3mQ0sw0I9SZJZ8oqNE7rVpr2Mbbxin2kAQHNq/GowvaHtqQRyX8b86il00vJQA2bSh0HLlq
YLVxE3o/l3q+HIZLBmlDI1TJatKiERKwuMrDdv4y8ttW47+/1bOJ/CjraPlmsy6jxs8/bjBOjXyF
EIYjZy+s8C0HC7YfniyoAGLuaG2yi82qKF54V6pV7auD5uRZP70ggBpUodWSO5kWc4JYujf4rqIz
4K8MFnpqo+1cqlFZaTG2nlnYxSGyop/e3uk/jLJb+u0HsTAlwu0zouwTLhFIKgD08tFtstY1QuC0
oZ1pS/wDnyjPQdASLwR3aNwCXIKuJb7RJpPVId5i8XzKWgSiFIJIvDbFmsw49yvUkGoX4Q+jXXP8
s9FIdR2T1xKHUBT1tVbx2A2LLwWmmH3PWsLaNPptpX9THKkuB45RFyj/g75xRLrypMlj/CnJfvh9
rdhS2ei6fHeTQE6g6mNvj0+YQ1OLyxIbhyrvgnTWaevzpzZbMvuRGl/JZl1bduWJyvnlnE14/f2V
SNtIRZU8nGRF93myPBFcRGGG1cVRuTqdDWrqgLpQ+ooH3s9Mluj40GSZXYU15DgiBjdO1NeSOfeB
Pfla7dCETH0WWcb0DRBe37bs0z4o2O9QR+JCdB+UYZr3wEMifsXSXj0xvp2sgCMRrVZy+Z2DkTIt
PXCXF8yU/ZTCjuFS3sGbONFgVMwiiwGV8K4jqZ/pKYrVCBUvuXFNnMM579l7dT4TD+umDkeo5EJK
4V5pNn9KJR7NraFaXgGeFIr5bmLzHabhLaXy7fpupEeG9BV4W1QKJu2w5QP7LcJ12BobTH37ck7+
YkgNevabwgmGlgsyyHoQVQ7vTaSVe9hu69D82oCP7ntvGxYbhY88yHe5Tza48ZCxh4QTZGn5iP91
Jjlku+4bjMbyVSMrcuQfBqnbSzS3fxERCIvrOsW1Jgb07lJm/hxyXooFNz5VDvuQB+HOe54w6iYX
kYk/lhvSxShWAenzQT11Gr+SQgTIrXEUzGaBfe2rTuzz9FIaYL30e0KBtfo4lpwszM2VEuY/MBs2
QJP/YEK/jG6fF6uw4wSaoIidDB8um5eJtqvjMhdeUu/B7e2z/HAK1ZQj6ouusY2lYX4gZT9P8NEC
TwhSZ14I2SJp4RnXivrU/nuluu/yYHnaNbgK1XGLZdcQsdCLvvz3WNcK4E/SXp9OZbO2ythKpq8s
nh3WJbffDVnOejfwcc+1c4M1HJq3t6e5dfwBc4OQ2+bGUoaft0WB3epnceD0AfYvGAK3WTH6yPHw
sH5b6VqJnwaCY2ujkTTaqja+5Q2UtCTTANUNDS0b6AvTUYa8x0ZZwo8KBgvFrLWK3mZ71QoOVDRj
FMtqKsNjwR5J2YxT9qAWrK4nHnmCmCZNs8n4xAkIoNgE0Y+E3b8lCjTvfnbvJFJWihrccJ/HRXhX
6hqtPVrxhMvqt98SE9rNP8uPUTJ6Srtut2PMN8UOFqyGNd2lVndx3MTi4Z3mp553RazycUtUvLAK
wk1WEfc9E0zVEOm/aY7I41w64VzxiXr0jczDheYg6qEIKNlTaVxAeJ8e0e1b7uKcLCtlPiGMzozX
X9SAK1zvQbCbF9HrsKPjrqUFiN+FtkN2UcYKjUqQMzKLvyVnse9vMgKx0yO0lEgDRXJMAYraXIMe
ox228n5QJuu59NoHWEdRNbOhpJ0orj5OQtHtAULrbd7z63H1/SdHgD/5qNODPS27UplkNn1cb0s8
wkL5K0OLUwPHVtcXSG5EWpS/scwG1fy7uMaFINgr+aQeWwz6bgMN+kVaOE23OphTLFCvq5iuo9Hx
RCXmL7Q/O/SnkBNwKO6XiYmXr2GpYnW8dSLIaDAHUOGfxjH2MfIeKmToqAy30Y5yqLJm1DAkpxHS
Ltvni+Ixwevllopa2EDBuuhMrOYMKZgsCdVDyspI9G24/SSoWyiAAL/QuMdmXz9I67h3qLpJppCp
79Yopt0w1nPQ4iy8mNyfFeJHRnRBaMZmgxIOQ5wJEmjpYpaUCTxiB6LwaK4z7EfubVQx5Pu6m7Ym
vdf/UOLm2ub7VlcFBiZcXeWxSpqMqSPCVrsRu5nVwlhIzYa5+Rjhpw2/4SgGvh+WEMIe21NGfR//
RqK52qLzV4cTkeegZgZAeWGEQEWXBeAEjnyZEQxww7Bo6Wat5MDWCFuqUk64bbHPMVkv9yU2BWrk
HPeuSHUopp0IHWbF6Nbj+44Bc6ALXpPqmQRt9Y53315BeT9qt0ZoEG9EQk42R8vzBCpE5+6iGWaN
gKeSpDwYWeA95AwkuHeRTZhGmSMdPkZzZpHlpV0Iitv4/uAlGd5VP5i27V/mY8JHyUO7aGLkaS6A
dMLbQn1Q2WuxlfPFxbJih0qpW3Zf/pj4tBiYVoNbJRJ16ndQ334SAe0b8JJQQmXMI3A7HRhEYnPA
kEUPoaY8qeiUn0qPDxuN15pdvjCCEdsn1OqBL33CBcbjUUAc1PUui89hamRNyQZ5nMpQjXnMx3r5
Hxf6/Cf7FQGi79C9tHZrDMIQahXrXF7iHfxIObNk/cvH75lJNrGBcy1rZJpoX2b5K/LY0BOqVfqZ
VPsTV8mqPVOjktxbtQ/Epo5BJW2xGKLMDtEkFdMG0Q94x5plB0If3Kb++HswFVotgQXJ8ubmWZpn
1VL6+GapQz137iveP0jOU6aketF3wRxeH7XuwSHjX1iCevglLBF7ItJHTXQLVif3oe6lPGeF0eRY
NqSp6g9n2Qqo46FM2VB8NaeV9C2PIrXQfPpB62Yu9VvUqHuTLMLrCgfvbiswlH0zj87hGFq/ImsT
9GjIdQXGL2JcKkep2NFbgEDucndtV8vYarblWNMoG9cF/nTfcRPmXOR7CB5ip+Q49wDKZyDS3AP6
vidk9oCkRUikuc6BbXuG36YfnlWQhlm3DS83Oz+fThpO+1KgH+WwcdmCGMoBG0/CgvxrJpXYxgKo
ZFZVKKmEwWaCr/paVjEutGfwCvBw1ze0Hmpi0a0FxyuNdZzb092r58r3lyjxWGuvUH/gJysFmlu7
4AsDi1Zss7KZkGxP7bKl29O5GxsjmvCtLx4fe47OnEzUsi8Mi1aODYGc9F6WFFzqB+D9xHdvg3rZ
pyRo2h77jErFKy6H5HJ64bKugGEMAnF9k41s2wlbDtgCh8y72UzIVj0vvCRk5op/5cnl2YqDOa1u
KWSMmzD3cQEeifgLi1CmBHsXkoG/6RZPu6QaD7FbI7HWWJmOY4vGhfFhhQIxNiYXfUN6utNIu6RM
EcVZc/8xLSHFjEZzmGXN2K5y3IE2P3DFHJ0ANOVRO+AtiK0XQCagcaFf1T5JdaIzSuhja0UW+qqp
RAs4qOqLlY/XQln1gSLnQzByaRmYOxZRcr5+5wuFeH2jCdtEA/gKTMe9n2plubKSQb5CdZo0FF5B
zBVkixHd9Spr+P8Gns9gDMK+MnLtubArwFqLVyWRZrmXjnqUimIY/9ULY2Y1YmjueGNOIbMmP8Bc
lPRuBJSY9LH5M3W/5wYaADgcmlTLv/0/6ZdM6rEVYgduwXffsIPRmXeN0FaeD7KRv8GEtdhhpwbi
0419Ak9JCNhuRd61AIvLJfgJhHYE910bypwSKkvmzN4As4IWvnD6/SBJl7XrkNMaeTBSK7beDy7/
uZkUMmVyrERz1BYexb4tjf9QpmE6Uclv5ea8RanMbmPxLGLK1SypGXhD9HZ4p25VkTw796rP3ZRd
IZ+PrSvq+rlHLY/IPvnVJBHlYmLMWWqL4Mn7fQpoBEoYN0C7AMF4FObvviGkCE4nXiCGETEc0JAp
sXzACb3RO6lGKjbe0oxMGk0386ftMuS0M0nzDq+jfCEanZqtSnYJyJxc7jBMHakV7cWZkjNApt24
MlW9tbM8MouwxHolGXOk+nAvJkR1UgEeunbt2Bn/V7lAp3pGePJGm8dovo3Vx0xFZh1NTAfcYWFg
MLvGrfI+u8a0j/iIt8VXMOPxwoGB47UqUXsr/qd6pvvMMluiUczTKb4ZqylNFa13BBRAuYOE/iIT
8Ux9CqLa9yVb+mNsfwN3Gdy/T+KYe2nLLizF8h0tqlXsJmvLIjGdDwnIGsrw/ZghaFAEky7tnp44
Q7Cc5op4dSiciTCRpImZZuPYtupAtA3H17NEa+TBb1syWkBcW2D1Xok9hviekGJme+uYIyvshIQz
l+zAZoUcKvBl2pBkv7c+6a0lSsGQy+BZO+Y/qzi0SMFLLgpJ6EBkDMERg4rIpvJXw+1AoYQ1Zw44
PHEEBvYO2kULvBBBc0Ux+gJLgzR77BdVwmCoEVr0vFSddUpXcmdg4ghXhV5oDEi1i3DaDzQdtJ+3
5KK9r61MBjhLMzMVP+2z2P8aK1DojeyOm77GKp0ZQ5Z6RxGb1/69hvJy+fPv56ErETvxFO31MtTe
1oNsSNjRBO33uZUgtCyYAIRk48gaxf109sT3bkIc8BXSp6AqvQS43UhUZvTBWUm6K9ejBKzufo7G
ABj7zfTxN4JexSBP8aK9g21FcH+5Xf4bq+UjnM3mYo+TLjwddi2pGENj6a5QyB5J/MdXRRyNXuOU
N5PtD/lRQywjaW/naZPqDdifbEE5ENQEKdlDzySdnEaWsLlMZYqdxmKWSZYZem7zAuYLoAl3cFyd
EPv0gw9NEuhFSq9V2jXViSRAXT5KfkJirCobFLBn514q88Co5CXXz5B+7wfLGVNkQ7/2KaHpvdaQ
Sm4GNClMYCq6DbN86MDt8NHw3TwbsTl0kLhtYANOSIfetHiaCUCl3Ukk5AKMwcyQIsR4W3Z6VORA
NDfftUUOQcieyvQU/1lWgTht3WaUM8FfCyQr8yB+l724+E8vnEP/wMwlQbbmYguuvoMraaNfU30t
DhnU2B7WC1zX7ucjPAR6MeeT7nfQevC3dcmYMBiPAxa8d85lrnRhldN3ihNGI0Bqq4N7txB4Mr/x
3FHNPYruVJMfYObELG9T4MSuijIkvyJMlfwGI7b67xGql6uu1xi9uFbbuEF7h1jXt48xr7MJIruT
+IEwfue7xXSY1bVOPa185X/Ku8WZHi3+JYWVcXb+n5DAZlOUFmZ3aI0iDlEznjvwJesAzntTkeCw
a0H2MA4V30rn0x5tDmqkEG0bqsuziGl8jNWEYmW1YT9Lapll1noLmn8suUiWjCRHzZwo4d0v90y7
IX2tti7O/yqAPxofjVuLzloVJfA26OhERHYnQ+stt0Uacfr3dRWiPVZVs3xfij8lCQ8eshdmIXQd
K9BK7hsIt3Wagj4jigl6szL3AhiISpHfEJe9gqVrJ5k9wLtWmih86/+1BFWOWdeGJO6Qohvxr1zb
h5eLGckAd8MRi6ZqHtOij8BlgMkuUWC7geujEOjpguPxHoZFzInlokCisZqcS77SJQgCn/22xWEO
x+h0hdV9Artk9CWZAds1DQrgHrRTKiPUDJGimuRhlerRUihygc5Pt5Ne0XeKN4updmX6GyVhV5iP
J6NxEcr1KWZWrU/nmseMiWTjvyyyr7CviKV1WZq7C1/n1akMEplzDAkVdFrC2tYnCLk/OQY71RWw
m7sf9/AxVSaZiKunftUQun4PX19AySFrRbzxFXlBwJ3R6nsv+iAU24UrhPnLu7kp8+lnN/qaDrY8
rCMXtaemHnw8iSh3W1Xq4vyAYUahw2djIsdwidPIhndwmaTpbCG2Y5P835ONYEG3l28XC/IDhwwY
g+N5lMy0F3rJ5UI8vDwfnFn04TVjprQjBu09mvhW04X24mt7Rx+kC3IZzPZS5v+PJEndbGqi4+/r
aist9vPMtSIZ5vmvNRK+rcQRjok0lapIylVtYxuxGCl1KurdaYIgLld+QlUQcKhJybS+OPEnkDun
IoPopWjEHgYJEIDMBruFd4eWlKCt1CF1f6bGdHnlM/ySStzGDG5Jt2iucc+bDBE4lB+TNDuE1ubH
bfvz7nuqoczgkaZFrMSh5BOjuGaXajpt8VweQxGS+YW4ap3+WpPHvaVJL/sMFWX3U6RrNuiKLJvw
S7RuNVHdveiLypkGROTx+0RTQCuu+2ZvdBQMQkLQ7lqHEQMCPL5BnHdiLPvJ8Zh6i9SQdNzsq1h5
iGRTFs8Ri6sqAnbegdKW8pGo6c7POB92e0ahFOYAf0Gh7zzIPRud2THDj9UhAxRcM55V6AVl+o4H
drg5ujuA0hgUXaNmEozkcJlAS3CjosmQdaZNsGFYdogIHIh30NdBdWbllSBA1/I6CGAH9bcYraVj
QcDIKoyaiD01Jjjd0rLGhGmvgUSUmlo9Q7iNyg+heZk5AHqqPOouI+aixJCQ+Y9dOwXq/kWmmHxH
tnJmcw+YEOyNZkqk/U1lGo3vQqCrLHtXqHEU6z6Q140e0GF310xRbPC4+0Sl/ZjT3HSSB9IYAh6X
ByWBTxR+2U8fd+w5V+xRpZo8gZDRm8ZeuXUIUqUycJiCGIFz58cakWpyD2NVVee7pSLbPLOd2bfn
dus6uYYUaAUonaO2i7mYy5REz9Z1RFu0lgSMm5rWsGr/8GFVNZcxN7MXd6/9Soj8N5COOc/vOMmL
ZGB2wsUJDgw/yD3Iqbg3L5EqLdQkwasFhIxU/kX4PfAlIIJ/TRbngyG2dr5+dYHR8WLpKvxFR8aM
dpa8z44rd3tqbn7aAQeL7AwAhQ1SbomTzU/cXXtjbbWTHt2i6RFi5d8B3F6RtoQkI+hYYV5zLCNR
K9Qgtmvu6fpTsB4otSoZLoSsj4YVQtab3kq2GtInidSp6BjQw7f3YFdvF+mfPINhB4RhyD9UUaIt
rSOK2EQKLiLSoEJCBmo9/mTD5RejgwvgSXv1buFuvK/pBwlGWKJX0AdkkQOQmYsV8cNk7pOUneU5
ehy1x+mZnqq/WNQoIjPVHcz1z2rYNRyliQT/wcmjrNcrTpKkxt9Us1trwMs+E17GqsfBNEGqCjRC
/LGRgmtdyOuzN9JrmxaUiv8LSaO1QhJhG3BhdVQWI4ZY7DbTT5lHKxLuGfCA0M8PXzzvEAo9uu0x
h5G0YuU1zY2waLEBFS8wehoh45SnHViysO93DaMNGz2KXaz15ge7cHkwU8+7x+udDpldC6OcGH1g
4NCGlAcMQvQQtJgQxBMinEGwSS/MlCXdIr7pN1FGlPUi2AjEF40Htid6mvD6dIymYVNw0p/ANn2C
aG+dRYf5JWNvCpVqJMhfn2lT2DAfesLr3rva0OqQyFmgPzOJ9rI8F68HzaErm1o8fzlHjelE5P1A
nJQgFq/3L62VHGzXJwYOGFBvPiv/yub6bDCSNY3oi6q4afgW3RyOubUXLTwmhA3tkPLIZFeWHkWI
dk4iPSa58W8uedHF0iVyK+B1ifGtv7qsNFI7ZkPLED1oJpZFFurdnGppSJp2bUDgl3Kkay0FEKV1
yvxd8Ikg5YnLlqzNzzbQsIHlNYZHRDjBUSzDKm2iHQ8N+SIqnLr7u1c/934EHGRc26i8a/gW6TaI
w5BL+kJQg+mW9Ut5AnnNPF/evYM2h0FL+nJppJeIqIXmMnx0L2OGatfYSPPZu9nsqgLpJYRxpvXV
HSZiEuiC0uuiXf1Ab1hPmcrVw5Plb7evZoPtOOgOUemJuz9XtuzE86nFdprrKmhHeV9DPkWXgtNO
LWuK84Caz4Th4LOrzLz0Watykq8B2gJiuBaXyeGXMPeKkOgitbIlH+ZYbpnS9PIDdTY9zlqJt6dt
boXLQaGxd00KOWekHX/capM9yx9N4Cktd063rr8x18gPaj0mjf6OPogxOQaIWlXAs/RJvt+TKS9W
kDt/Dolo9ltOu7RQP2ndnHPBTRNHTrSSRKGVFvrYDQMkew3yyYaMgc7M7QRYo85VSoTb0BVm0Jwq
S6W3d+Fcu4GMzvVhcTB+GikNjVJdSbn+SCUmfb5A30sqtTqSP4z6/6+yBb2kqFIo0UQD+Pco59BD
utrC41+qjAKX/V6l4XI5nZGLsJG8Ffl5hiDoNGZm2wx0BLKFvckY16edaqt8IkXAzmDkKKQNTbZM
iqzGizJA093EKaWM7tX+J8zzYEfe1rwO01tQxfoafGiT9hCRcvMBC5GmIJPcSzABKYqUf5RMnk83
bXw+YR2VYwiA8x1tZd7lekSAH6CeNuAuX6Gs5kAmAlCXzPiMO00krk7IyEquIuPVryHN64jCWxhs
jP9HDPZRBXpftb048ItydZAtr2Ce38ghVsdZ0R3oHOmi8EXXNWS+R0AL7tIkQYsyCErvydLWK3lI
0ef7atSFGaljkXr1S5IuDOQ9J+i0n8xRZs0t4AXSI/ab7dlmTs5kdIruj/jT8fGGdRlGT+a2RSma
8F4Iyh3pj79ZJ+SVTniPgkpBBEG+fvC3M9Gh5hWJi9V7bE2Bhkg77bmmfmvizLX0Pfl4DCBEf9hX
kDEcDzm3a90uVhd+0MyJc/r43tONVgIAqYHTmPwE9UuLW0jr1ilPnVVHJXz9QW+Z57H7l2N489wX
gCY8fVQgeCYKKw2hNCua2OFaROOWpZiebMv3dscVWoqB4PIT1jqP7pkXhuFC7MujiJWjYvki2ksN
NcL518dtPYjXzVWk/C4A0OR0MBPP7K+BwhTYidZZVbTO2aghOnsZVs3U5G9LMrGOM8QhPROrwI4p
Ivk3DFvLpbR2Z6o7c7J8NIEXDMk2XHStseVG78+zxG46azE07ugEFThh/sXeu0cjvR1Z1U+jW9ES
w6BLa5SneB+ZmvvFOVIYLAvyW5oQrRQ9nUgznxXazzxPd0ePznBr2ADJush3AMjM/2CPP42Sr3ke
L0aE12Cai2MZwQY/mh7WjNXUfinyZ9yQ+k6t92VbpfbVPTIedm6uNopr50wlm1atawBUJzm0+AiL
8iVbER4Cm0dnx2S67VrFlJdH1pBmwrZjphLsw4BYResN5vw7zDqqwXak28q5Oo9g0iEIbk2eNamF
xAhI1Ptxb6er+ouw0pPSjsr3xl9TNr5/xsRXiY17AFHSptZwd20W7mk/MzBNbmFxyibJy2d1ysyO
8lVEz56KejZtOvSeYE5cpMA7uOO393UUQlM7BttAoioX+/6PKqrQz4lTf9Mp0U1atInD1hOcmlKX
MINyn+MSipO0oR5snMml+afEYDKKnM2YiZk/9MoDsK/eXwzOCc7NG8dwSxe7SN5qorjV0PeENVh3
dqqvw2LcvS/coJYARp7x0R19wp61fChoDmOBGzhxFCFo6JkJd2MdIylvKGpdsG0NJdTQflLGxYZT
LvNyW7aXyX9P+8a05tQ0U9CvGEHYi5xBFBtHYCQDIkTWzGfvp1dCl+eTl/q1IzkEMqPPMk8GIZHg
re4s2DVdJ2mh4oz+zWaaT/hLyol4nX30DDYsOtZiW/Zb5Ybei6xUJehcjenEe32NJg32k/5x0yML
5g2RgoovIz2sb9HlXhMQH9Q0SKbIhGVaNIAf3sKWh4OYIoQQU8vlE2fobmGH9r4vInZcC1aZ7ORF
WmkqSp+inhGbFTfV0s+TCuU6UPALc6DUQJzw5sAnND6qM19vggUQMD23am5Xn7vfTEalhqZjCFh/
1lZKvqkDuw8E+O9Fp964PsKHJjzzehWgZcZCdYWoXj9Uxp9wE0eqpCEMK8guMc6nHRCZEVF2cWdf
wwcN7Kc3g4reLHt6Vrknu+soEQwnWrxWTxctN+um9ZRAurYKVDbaT5/fGZqL6g+UN2MOqZidoVtB
jUZhWJsFo3I7noxwbBdaThPI7SRl4F8St7q18SUmde9ZRRH/nLO2vIfEy47y+cMyvXkihavW4G3v
MRDA5I2coCR8POEEks3Wb2eRO5zs/HuXaYnMaUijOCOJUNggO9Kjh+2Pz1lkH5GfyvMj44nrSxLd
6re8vYCKwafa7NUs2ygI+/kl8Rr/lclWDSrntBZqV7Jcbsuu8HxJlBgeWTSpXCWj+w1mUwLs2M5x
kgPsBzGwT/t4UckJMufnXPkPuz0MO0dFZf15Qgpn7Rrv55mz5Bu+fNcTGGC14V4fnPnCsENyVuuU
+F943ONxz+sX01DecE3iNwkgDuxWXmxfQEMo4sSzk6EVpdpbtRZMZr+DhL3FqW0y5OoaJrMIUbO4
ZNlPz85GW/LUk6ROsdkEFr0i2IKff003wdJPzaZsX3qG9ldNHgXpouc3qTvi7nPQPKZoNlrDaEMI
cgOIf7NeOkLetepNTwOtwzEEST0sUOPUrvhytkYC0pg9g++9hQhL9F5bjKkqgv24bNeKlh7Oi5cX
xuk2f11CKrFeU0avW1XSpHL8Jmiovsq8JuUN4f6g9AGEUl6NKN/g5+5MsaNt2ZmY+/t+sICcf2YT
/mKMzfZsWRQTCsD4BaVcVqKgpEarFeXUE9/4xDONu9QNKu6snt/IAcw3YPm3/yobEw41OG1346S7
tD8oo9NqazZt69DGntEDi+rOpf4tAdkMgpmvFZaJJLjdtLSNsAETYZ2peR2aD0t68Ampv1uoDUPO
AOR8edDnz4ani+ZWTZsLpGdlHAaioGZhcmDn/UvDvoWk5UEQlbJ+K9lkfBYPaTBJc8/a4GIkFIU8
Er5XXNz36YvhDj6nuA68F0hU1y0qanYnJCionFWNj0snqjNle7kmpmCfHmDwrJzzzXRHMQOlus/v
WS1AyBKIe4qooohEenGinhVn1tIVgeAnU/MQeBDAjRUKPCrPi1IKj/RaslaSsazgJ6q3rEy6Q+TU
b6DCBWhjJpLOjyBtEiKJJilkCY/gDJyEAqX9bM1/f+UjVoFXarjDrNBTPzf7gXCFIl49wmwbUPog
INYnNWSVEq6qtnD4CcEdVdgd3gpvaFZeJFRGu/wiXmimXP94fCrz79200hfKz+ZCsGPg5VZinT7A
S1p29Q/rMA6/S1cbVn9qyNLTaf/PbOyECD45RK7SDdOMh5pwcOhZZWc8Ahmh7D9+Woj6sM1XD3+b
d7rWdq9xZyGvu4SssDMWCNbQB6AP0Lqc7YBkML3sjyPykhB1RtjpTWsuNiBGbZvb5znDrPD35HYz
m42O1LwPeaxOcTvpr0zDQIwVW8bfXG1pE515VZ11ipuw1VLCEJeDgPuI5CDANMqng2vm//CgUoTv
/fkxRc1Y0UfFrnczpA6WGLHNyZweCf4swxhr+kC87bCvTLBQ0VHJzWXKODusinlTDYUeZviN41WM
TjhyjHzZoExjsV40EG1tO8KMoO88S0n6czwcHxu2Up0pnepv8FXU4YJXD9z8rhoMka83xSJGP/JN
QqoYZrYowSWdiJ0/i9y6+yAh5UJ3t7aSkyKXLc6mDduNT1hCMF+d5b0S3Zm5JlTDyJpiIOW1sYvj
G0D8B6I5FcUfoUlRnHi+daLJ4lo5zX0QHKZ8+kJu+/NF3Z8bmcwc0fBWDNctA84lMwsqHS0uvdED
eongDWWGqhycukx4B+KzrTX3WxwWG8yeZ+Z+6tGWhAwHBTmCDhPkJXIIhOtquBUu+UlxHgXkVm5w
WSyNwcGpd/GL4REB1BodiMPYESIHtb5DuDndcTGgRrjzOYiAwQGv9xuKRtt3xRq6cnWdxSVPBh92
yQRvdtjchWCxftesbwQ/gVXEUWq+GKsUOmNu4+TBLlSSBaJRp7FKDXrTbIygVOjRvYZ5Uj9HgnHX
ga+507FH+i1oaIvbsdjGp3LZrdFHEcipjYxq2YNq2/Oq/J7KuD/swCMjJ/nwb4khyaVfZfIb2htW
V1bT4F0w2rgr1HD9pMfvgX2H6OEw/m3bruigtNQxRz7Jl9xEgy84wrJutkwghXPHFWOfVwhPaJDo
KGggeU7O8u2fFPbrCJEt8sLK7XuG27wMWXqS85ifeIm8tGDKblgyB8QC9BZZ2zMbQHidJHWQ3GCe
j1R1Oa6NUJ/VAylroJOgpf6vT39izEvQkI1G9PBpxsx5G+It9k1lUm1y9onpjVwrD8k67AP7zNQh
LroMnKoGc7nZtM08xc7Y1eyensmzgJKwC9anEHTcVRJh1ugsy7BincebwpP5Rc6ugCX6NiCxBGXb
A7evnaDt6ynBUV6L5PI3R1pXgi9m4OW+iq2dWl3H7otdVmlxyAjXruuZ7m+/qM6mtmfPkl5cXrXt
rV2sS5WzMemiQh97csq0LNBitSCXNbvhVUZAtvFH5L7Uh6en/J3vIUkllIkqNeDF/VBpGYrIRl0n
r7JjINKuZ7Q5fM2xWHx8sibjTi1p51LTS9ZtMLNOhU+2uw/xP15YIscIYUYfZjPckKf2n9PDiUXz
GXZ07aTLkcQNYEagpFXva1GV4nXuubmKoR63J2ViwW9khKJGCJ8QrtzVvv4D0Tz+evf9GXrXGfdW
EnkufK21+KbKUaZk32hVsMYvrhUFUeP1gs2jI6wwMZKVyPqCVmYCqjxnQOeSXa3dqYoAfmoN6dQa
8d/fKAbNciT7uJ2xzDoXVnV6ntBRfFt8/uVk1qRpV6yugJoz6JJAfZqhtar0gyWdnLqBTQ0nfOJ0
7Wpr/F13WmaJJwgVIH96hWGMR6boNDcXROmnBkymYRQHh7P5eAPzGeDZGdiieD3QcRYBYHnQ7fvX
P4DlrHlRRXA66XENItpQEtQy3ZaufO6qFinn23+7kfuR3XdQYIXJDgRpb3Jr/PJV3irH6DcOZQHK
ihwfVXDaulYfnFNxRUkBpkKw2v7AvTgS87qXnRPs3gCMJif5RB3yuz8NNb8vJoxXe6Pla8sIhijo
t4bJUYmSXiHVS9VbG8kiy5btXY9HjqDL07HmX98ldJHIT3PwVtclbJ6RLI8Um3JjrK8rYk9OX4Zj
SjS3605klKGhXpWrkNzfkhuP7Km96MIWR2PcNWM6B0rphHu2Kz1mfPEolg4euuXUVkhHIHrOXjUe
/ZLZgZwbP5kX/zoedH2eVWeTjLdUADGhterb0CLf4idz2yi3ejiA8EBZJS6T+uyGDd/0pNgaXsvb
wpDNeZEw69xLY/hSVBRIKGEyX1hz6I62jkOcdVOk3BAiPTCQmZQmklombbJkUT/H3l1tBdXY9nXA
57MUjHav37eBdLH3PVQSBi9F7/aaARImu78symX5RI8ORsKvrfMOq1lmORAysHUseY8eU8rOZyLq
rBa57elUE92Ed4kZkgQzVLaoiLvtcduOd7g39GDMNijrHsFTZtXVmnZDpl4hVzqeen9bgOTyNrRN
kI0QYuBRRgzaXY84PlSJ9CHjkHWMpTMM8uYTY98XWnRV3mTV/lrSfUsZlNY/n/WlzEVOgeHY9ny4
N8/yRjrL081kQP49FfXyvRP7I294y6CRVf1gkBUVDcPgGcZNfD5NFV6zXlHQLxGjYM4ezNAYgzL4
UVXKj4FXQrxmAs8I3TXF+qD06S4XIFQbhjzpHvtIeYY9doMadaBwkeCiPNAM4aFkKt58NEPxxeuy
j7uLNH/GvlJLZTrQ6r8zGgVSbmtkdp/WdlFF/4kYv67HtcmFRn99Xotsd54bUl2elqq0mY44P1ub
IJBwnQYJQWwuAXkihe2i67duO6rv+C5xuzMI/K4hWV+6+Ccm4klzAlNifxDzYd5YlBEJEQLNlMKZ
V+5xubE62heIVJsxus2ZsBZ4VV3jwKcR4/CKCgkPfaLSB4I5cotzjhgPhjAeuKQzucqm/3SEoSA8
YyCwERq7lENSrmff4HXUWW9Dgrv4OScDGxRP390fWoUDzt1q+jnKApLMD43VbLqIVspZKxYGkvcp
SMmJMXuJ1dxymbN2WD4APiuV0dR4+TXd5uwpGLKsYoyMLhrrnRLQh+mV9bslnQIBgUDIvm2EoEau
bKwedVAsXHKM0YLoOG3qrs30xLVx0OiHX9yDsSw4hb1JCbUaYJ8ELLyd+vSjmLDevQeTinT89587
NRH6OVWoL+3e+J3Q3iUDIeqNTCrFiMu0dboRgP4rMnuo1lEDR1b7rY+2iFZfKIgRX4Ggi0snFq5y
XC/mL9nb1hqEj0uS3o4WwYX6MaciK++dtVSEK6TsIpPO2clo57g+75MTWhWdYZw/30qXoxK2gV+9
idOy76Vqkl8al7X71qFcsVMYYBF4yAxVgPbgR9maetsQA2a5Y/pAddDOshWY0m+kdwTkQUoSnVYT
Ak5p8QYr/P8TPF7jngh6GVVnbpfG+XJbP9cQ/PRn/OMS1PrwWTzYMcM+wrz0SFDKe5jiheXl7LVm
9NNslU0Yp1gNDQfrB27vMs//BWOSeVE0KuJCD/HvwmL1TlIzqR1mH3eMJkNgVXKJFA0mXQ0aWcU/
DwYdvpOVkck87fmhFh6M1iXIWErPFq27SCeSHmjr76I/ZmCP0siBUbbzJpgZJ3q8lJbGDSBT3V/g
nAk9fp2MNEzSRR602u2mAzghsrYj6JMQf/m13LbOttI51wW71/c0OunG7OBd2dywq55T5mJmFsve
j+WMZYEPLPHR3CoJ9cc0nzOGliFjTps8pfwuPb2hF4zBxtzgrgOdLfeqGbzLeJ64/NIYcYtsOjrA
3fR9MQm6vcaZ8ZocuXqFZW0dVJD6LGlmlGJSfY7h3X9itWOkIu8xCmiTSEbFXTLbabzlBZ2jWTYV
cHEYjd6yb95/adhnklusUFq/0oJsMovHo7HbvlqhDl6im+yhNcFKwGJ/wvGQfY81vQTjWONQwbiz
ccPLpYtipbgCAQoXXLaFlKRgMuXE6aCMoIRr8pfpmDKUKyDAy3KTnIZoq72OnyqFcUyK7G1zjBr/
4E3KrLWVzpRJHkJVTxzZlvx5KeCEdsP0tTS8TFBiIybYyB4CbyltSrd7Q90tli6McArV2Sk6OgoE
udELA/GjGCk8bsCaneTaAZFuuBCkNEFL+G6ydli2+h64XPjHV/Hgq14nWE7BxiRQZYY5vqxROSGC
2Xkk7fb4c1Igh/D7IuygsQo6xQ7DdkXxTocvw0ccSI5cjhEhXTEeZEY0MBCCppIxnNo3VVhlhhGd
mBhmsTnhzrwHYWKeNSzc6w7w6QOS+fIiAfSLUFWXTIw4+tS9fIe0/ebG36eMt4xeUpIfxgnDNBNO
0leU5MRhRAKcsaMs6siQJ0gm1jy3KG3uZyGOphcgsdanX6S97Cx1oAsSu+QlzqWN2mY28FO9Xvfl
4jTgVLljuOUbK4MODIpujTVJ3hW8nl8XotW6B701Eb0j2Z+DLcZc5Iu++mVJ74izV3hy25UXR/rp
Q3nMlfFJKLJH2/eeFi1cL8CcIJpmYKiCfFaGgFJKv5Y55NLiGxk+yvoCtKv4iLbbbaDKgE6zwfsi
6oTaOtl7f2iUrSZH0pUSC4jzW2zWCovNjAJ3SOhdEALB2WjTIoD9UVKq/zE2ZyJkzXCuGYdUV+0b
MXgmIMCvxyRkIgsqm4w6edS2IHn1KaHwkT7h3ahtt7VABLLxORjvefI6cV9AQnbgsw/YQgNQWcgB
Kh2syPumWGD5fy6ymhofnWnOoTRNCMbrmuTCNrp0SbY9pZoyHsgN3IjuWzvwdOZ8/EV0H5zHr7ZI
TDqJ9B9cShr7Dk8pOm4gcp4zOPM1jlxUyByxOkzAkwG1b2cWH340Zpw36Jv7BlhQCnrM8NLfA9HY
NQtQRuGfBmUyzOF5VgrWIBBpGWbFtxwLsPMmMNrqtqTYZ+QjlkRT/A6gm4yxygXpE/6ZfU4N6YKo
5bPvRXjyX6yhBGam/3yo16qigALl5lBiNd09OdTZ30Yl/Ht/ln2TEmjdGVUMdfTz7EVbqxShrQMo
SNVjAks9Jnk+No4V0sFdF2ABK8yE591NzlbBNUWNvBhtvIjty+JUKjwzPy//xhX9BRZpJycYdAxd
Lg82JFdNuHtmzbLq3VUNe3nH6XSKUhw4wTORZibUAYnGcgr0Z1X2MHUWu/Hodr0SSSfr1TtWpjcm
qdoqPt+CSReRrejnHzDJrG6BPZNhJ4vHxyr3slIaZ+O1V8Seg9MfU79aykmYkMisSBYjItQRV/Lw
vqrAGy63UHTTkOc5qur1wuC/mjIN68a9pKmYTSMjbCX7I71UoQzCOFARhT9g7CMNpLoVeJfRipcZ
00kSbc2k20VOpmSaD0jiwa5i5uVuMC3BYDQURDLK5abs6zG+KN8irPTlY4OPKjS1i1zDCEIsPi7H
lh98YobHCMsJpbwptyczP22iUoTWCWx1eZ29SZjYSi74PLWr124kAeaRKmXxVvECyL2FOhSzQ4rF
Rhwaw+kVKzyCmsAeJwkwHisHw2zoL5LOeC7/PjV5PFPt6ELx10oQiBG7ZNys4ThfqQyuLpwIkEgT
k9goxP71hUJmDQDUl0hLOp6XkPxI6BPBjVA6b2fiZ5YHU6CeOorkeLn94Dc5jBlpB5jrphqlAH9H
kknJVWWO02qMqyUWUZmwgkULDrOBWfYVVjzMNdaRaoF04vSVuOXysOHwX3xttheGgvzlh6ui0Vmy
JrFczXVAO8YkAakmsI0AKSiJKBmCZqF2TPIo2n1Z9SXTVtupE7C5lkU3geYqp+WiIBZgzSuLlv/Q
sru9kP9UoZojcd/IrHawu3kGOEV2q/9CWQ5l+qzvbqXyHtH+IG7R1uxN6R8s9qLiVr/wxa+xv6F4
y/r0cWGUQgWJ7eH5bsyf9USAwa/6VzcNb/ggD2G+wVejm955ZIeeuONS1lQsAKJRxNzgbHbquOOu
Tzu1fUyCUyoVw2ZmrkVbdR/bWzYEM4gvWJrCc5Pe0phGhtlqrA4AZcyU5j5m59imSY/GtFFRDT+D
o0fkUSNhh6wTuCK+HuE4botBT4NOX/7bUX7mpFmJDeTHJdhXyOSXLn6aRaUGspOytPHJYIKmuUA9
KGDXEANtMyYALMYHYsMpeljFLT1/BhZPSzPdFSo5EIl6b3O2OwAh4M3HV+NtL2TGqZKKt3VhSFax
3awmlLuIvEmVzrcERyySLJUyacLlkeH0Iz8WJz7c1C3xv3w1Ggl3/GTafboEWKJn0ih25z4223C+
gGHS/AXYC+/kFiAB9KRoC9v2pzFHmWa5iNm46zjoAJhXAMsJJ5vaacvq7NdwjzqLWR4xrXxQcxm3
zRCXSOZZovuWqlMwCCynvZqy9BtmaP0ejfg2A5S4Kqhl1+tThIuKmYGSWVHPY651HdwmUbfG7Ers
Q4aqKQcmaviyUmxckTZJPmuRfSNfhyJX1XFaLsKf7x5sgHHFeobLcDDN8JIej20JfqGiVeFrPa06
aCITKYJNFIAE/Fs+sKcbEFARNrQxcHJ16sYfeTOp+SjZfAx1bqaK+ujpJZNRbBlOlJxE1s6Jc8Lf
kTBCQaWz7zMPdkDn5I89IeLdsPxXYemaB06oa4206iYfViTjMxTOIDNswQtKJE7H8Po6XNusRWHY
hw1D+LIXYjzpKq1WZEVmwSPTaHjGm6VjnGWwrdxb1IfESVlkOuYa76MBPclNjzauUCVAZwGLFiy3
YuiuNiD+Jw3CRz0+RlVMxngLb7YeH5eYlGh7UwyrNiAt94XcKiNQ2isR5FDBt223Q59RYRpZcQiI
BmI2ozYX7jG02tizAyo9w5TzosQcT9Re7/05VC86a3nSEBUm+SZ2b+UIxLsUHZp0kvlhdZPGKkuY
pywy8twAGL/wCYyaSU0GihTX14n2cjd4/mMT/tbtO2hbiSKp4lkL3fft/gQqRqssR7DnkWuSrzAF
aZalLZCPOhY2GCmB5F9LM8wiKQEEZ7zQYN+STLwSytwUSSEiXXGq1Y8eTd/Ks5o4L6G1N7La729x
tEjaaz5lJsywDtyBpTB3o3SsYJ3Hl7M+5bLxk0gLBRPnzGPvWjzvaFMBIbY8M5oVOL9f7xHUBYNX
XiIwKlxFOoNm+mLaazZzbXLUVpPQbaWyKGsBBdMRmIaKNr0S/dMN3T2GXiqrnYMwDiBVhzscCWxH
lC/pWXo15AmRk01N1G8sq5e7jNUwiQW2cdx43PKgfCI+I4D/3YvVyQsBMflvZ6M4UmPLQ+J3MVfD
o4nqWZXWaJ+fidzegM7slQzvvlfCaLthpTlb68MI5cW8CrGLCKQsnlQ7C+JQ67RLyGLahSEa7PwS
FCvm5Ip3dWsxLsScfX8ip3gq3NMD4LeTwpbwdfvm6GfXmtZ2dJ8kZt20YaX4LkTTzqDUtIxF83ZY
I5xjSMvnDUsHyeAGjFvgfi8ALD3r4EC+k8JSmw6Wuf3UJ/QsiCRH/l65PLsduXLVpePQMDvvwka5
rADQ6N+sj6gx2A8ZuaomV9RUcQx1q4F47qUmHVkTDf/F5Jl9SGUaSLRc1kYv0c+zSY6lQ3lVX408
TQYi0O9+4cXdcWK2sc0XixKPpz/dj4KIQvjbGxfycl4qEe87FkC2HCIg8cUnOg3d2WwGMAWwM1Cp
WzAncEx/gmA1CiY35xDwTN6AXTgZFRuDka4qMYvykady2sd/D4wVZA4eLknRLwTK1tIk02dquqAc
9TBFBxNe3gUqju4knrYK6Z5jbtSGKhkLN7DseLaniY8rFf9PsG6vWaZ6KMnhSU6YxtI5Lsl6wxmg
A1fyC5tLYJqEV1h0qQXw03EOSrXA7mADuAaNlUWp/IukUX4HY/q0LF8Gy4MR/CLV/RZe16jMrPW7
HVl1u29RKpLHx/STfQKLK+Qku0CRuDbCw2Og835HC9o6NECPOMKyq7uMzYpQROQzgyrhcUDwllkD
tSumCIa/CXVEQ0zzu4S4K16U6yN9AwLy54FruUXlk4z5ckw9HQsL9V/hZGkem//hZwpDhqmA5BjS
EZDd2oER0Ub/QeYJ27OZPpoHjuKTHesjPlxrSotuAHtaDIhecq+9sttXpVftFJ0nte3d87UV0eBW
7qkFKiE6te08Ug5MNZe+Grc7wlocBGwHiZysWkPXwxQCiKiDLswahDvko/9mLq/LWzVwsQTwGgut
TKHjYlBU6B5hFqcbgOK7HvGafkiovOjFk0pg62R5u03aU0Rc5SM0tiCgbVT8BQwmJnafiw3kfqtR
hVCNMzUqHr4nqCporWLCAk6sUxuSCGYoZsw0UHj7tfEhVvR0Egh7jZYfyqfvMAvCtZwczkxZEGzJ
9egrdDsUoYZQVjT0mIgzjhcuGmoF8aDEFtMGhGsxBZhvAHDYFuivEARdG6wQSM2lUxqd7aq97VUr
cP++ggsAL5dAe3fcBvlUuxbveTtCT3nYlGz2OIDhtsgBipui7zgmfNydw1iJLv72tE+7k9et87Lw
2VY4KZaF2owsLiPWbkDywx5pwWVW0lipUfzlCYp8xf73yCyPA0YWUnGLbi/N7alMHtTZvaBewEI6
AmX7SQc0mmZta6XautKP72ntWnVJ+WkQwhM3qMlg1hpN4VElh7U56IACeQph2QmveJ3mC6s/f+u8
GPFtXXU0cgy7nAJt5RrCuvM6qdwfNqq3rTXDYfbgy3K5k/Od1O15fS8OqQm+yawSM+Z5Ra008K5U
s+rOQiVTRp57jiq/8+CZF9g6KLbMmjQgxeE1hEfnzwSzFvnrl3f7VP6UQ5ooxQ0zY8vLMV0yAtNY
vl1HXGvRPuN4qq8tnOsATlX39rd4c9zpJKaxxhJvuL6ZQA13SiVl1YBhesKDmwnk9HlHJX3X2w21
RKGQiZNAS1QKlUBufYAkR21a7poQI1UNAC9RCcfZvSQGpwzFRoztW63fUPQikoaZMbYAIagyqocI
SgqCwM8H/T29HyVQmvSq6/arWord3zuKmnj8g5SJpMEVOPlqupk19WXyYSz4u+MV/Pzww+ZI9ut6
E3ZVrnB8heRd1djwGM/6KrOK8SSNmkDy8aFD0jXq82EkvCASsFB203qSMaGxuv6EzEOpNa1+sF5P
FP1sAJPlgi6NOKmHoH3JHQzkLrhCPO1kvfm7mbGVgKsLCUWMV9UcFlvt/6gBvsEOquxWGXR2ErkN
HoRDFb05pUTSKQrAuljeaIXY5Gm6ZhmqhEiQ2xp/mcb3MUEcbrMv+/R7J/bQX4jfl7hOQqPn4Aud
plzu29cwxZwooxIulxH4WpksNIHHTEmS5xWMw3mofpgjzaFgdyOzx7dYE5mzJfrZhsUAmBAyoKJR
sa25/JUJzjp4Blo7YjFThkLGA35aNNLa1sKa9rslluMrU7umPOUX3XS/aN0wZL3ZOxcaS+gClxd8
Qc9bd+xReWIzfzbcU0iqkeEoJAIC0p11qzZFSEzScmtClE/CXVxVOGUJlRRvmzEXu7JPvgc+o/Z1
JfYhC2JL3TQDnxGBdKlXImJ0v83pyeb30oSRLuaY5c+aWHXOFpbwzxT5fKlKaHCZs+Bpdh7mTEJD
WMBSBafapm6pERQyU+Ei9srvLGmvvRMw1+AvnrSyFZ3rdVGkvTQKbLA3kOP2rea/P3ETm4ji2W4S
tEWoT1D/h9HhPU3BjXvsqcPsHtP4XU1fMDA3TrVwggm6PSmmtaGEFVZExajeepT1tDYrC3l1rhpL
9CG3zH90KjzRza7r2QedZ+7/qz/wvBtazvG2zFf3YNjz88/oc8LbQVs8UBXTD4F+OWmm62Wg7+J6
dXkl7Uq3OO30U8mLg5rC3fw3/WgQ7nLIH/L2oyl0AfEZ8WfKtyUJto8ylASN7gc/WaeVspB/laS/
mavVK+pwQXum/9fIaz6ZL2cerwPAV6Yw6VRMijtx1GR8XgR5lYIiX2ehinT5sHVDd6RE82EMsDDQ
fCZuBftuDMMh0In8qzc5nnxAspwbm6Bhn+slJ0WDxcRYjfx8s3HsNS64hYe9sHKTzXX+owu+nQL3
/Gs14yACHdUMztDcAjonixrfHLSkCfXH3H1GlyyhpgLCT7hAyf10DY4nZ3GhwKC+jMu+48Ocz7oy
GdgSMt+/RRzzRbyk92F6xDtJRR7U8Lo+boTHKnfBbWtz/biS6r6aKg4nFed4wCkBGXANM582D/KN
MYucAfEI69kZD8eEGBBsWgDuOtOBo5DVUCAylS9gNYHbvzRUlGqdFys3P8kNN0MOI9ObctdDa86n
fhJE5UPT1uxvX4jG1CJ60iqFTNDBOTG0YfLjIhQhfaUKMENPLQ6yHjBjMWy7wkj81Mf7DABw+yFx
GdAf6F2Jf8/X1ZS0+fKihGp4si46F+z8hg9XZwOI1QrRjM/HnTrk6h8hQUraI1cQg0utXtHbcvES
HKft0/bJ9MJRW2xY+YLJEwejRrUnBIeAVMya9bAwikXNSWaA/yKHDGJFIffysUie90B66dTrZXAS
LG5l3Tz0DVtJUMnWXEHB+Ten5EaX1/ZroTX1Bp5OqQDVsFvc3dFHWclx9zvrSTHGXgJZbVv4+eV9
mD29Vl0ecfwP96OzY5NY+Mg//kYJub6OrnvpzjFrfsZ9kr1ZLu7k+S8gdHG6oollCi1rW19I7V9b
nwmIWDz4pFREKdPAcf3a978COFLnLviS5TWyZE0dL8hjwPC1seBBrOp5NIp8x9/mO+uWsB1D0Ngc
P2EDdjQvRwCcSWJtchBSPx9w05bfzPE/gyE3hAYj22wlE7jklazqL1ZBPjUgA/xjSuK/d7ha0hX8
T6UXCZQy1EZx5xbcIeQFaSct7fxycFtAJUYyToMjGkUay9XS1CDcxLX41KpaLmIcblvElfFoYQ6S
bdjnNH2kcPbXG2Tuj/T3iYmbelxPSGnzIegBScGDy390RqTXoNkWF574ktXazKeI6f961nRMlQ6H
kEWEzQKkXu2c0leGFoknurPLoqP9iydy86HMQ0AiIXKLHF6TQW7BdylrkmOIotl/ZjiH+ImpK/ge
flvVQ2uZDTX7TD3vcGUnjd+mpujZBE6iNqtYQVYUu3SyeMAXuh03FfqYo4U/1brTfhGtsZaJ/W7F
93yXADTCNEaKhGive4qm3YwV99l0jYrpXuYjjwRuAMPu9kMB5fsT88RoZZ5Tog9COv2Hfz7y4WUW
dDN3uDsd3XqOxoyKR1pnUymG/HfsBzTPo4g3VMAX7L4R7bv8wblLk5J+VUMhwPSFTw/dXDjLRXTL
SlqIaKicLKXwGJRzyUehOLzd/KyrERbHiMt1hvCQ6EIGr949DqfZolgXS7WcSe3hUhQ/w7YrkMe9
vy84RnzuuPm59HLLahJ5LP8kYLqohCQC5AlGRD+k68x1vbpUeFNBqCE9Wgb1ewimCU3EoMHW1aO3
6evoAvWA0TP1AN9zwuX/1HGDtnvLmFnkV+uvlBh18FlyAisOFpM/B9ZC++W6rmE6vFt0IVKJwsaY
4l10zaBomYhCxdDDzQCuClIqM3y6hYH9Ruu8lPMW9+7bQo7pgT0kF8UoS5K5f1CLIuK4CDLk5V2R
FyScLdU/lUJQ4hJQ/n1Pa2sb56nuKYAu+iaAU3Tkyy3tpUQlhgOIRtIk5j19lB/+dW9uJqi4KcXB
U+fMOMiyqvTBMa79xbrDIAkQhlnTSjgAYs8l/FFL0Q0lDa05DPTFaCbm3JZKY6POy3rpGSYxvEA8
ziWDRShEkvcupgrW4y2HLrwogJAca5ka+FAZI4T0uNflnMd1CJp/POMTJg6eM+FTa1XTu/hPx0yh
rQLm3yswEOI+01tGyPhfJX6gNX2HAgR+yrIII9NCrny8neTVmPpzZ5KagzXEr0xu2IwG8Ej+7+Cg
clmYSkLis6f6XwtKMbL1088mlfAHyR/AudVUD5Xu/B119BZPpaHECJ6ymNbX95vWbWrEC9iqi2u0
XXwmDxYQAMAEPbUiKHQAGZ0ryXcH5wx/+nDeZHbNMlXQKyBcUCD2xuZN+fgPSn/q8Yp/OIqXd+cd
TT5Epdj4Ef6SrgknhIaaTTzUX8NThmMjzRvepIlaKuve8oD9h3DE3E23dbgiFPzq9gsYq45ivwcp
dMi/1wjjp56uoEF+q3iw4xcG36/HxzwGONEJL8JjnoGlLnNA+gY5sJ2fhcvV1AKq0psWOzjY8hFH
TgRCW7nAUxMlfze9Ta1+usYZCiXanJC4+ASwqCxRqtpy7tnaT8pU94WBCFWjlJ2kvv9Pd1Jf1YLH
YuPPbDNJsVRtTjuh5cmeiIA8+aTVB5Q+FUMU2oDeMlfYztDUA/t8c+iGskcpwSpCytN45RAKeaix
jsrlDG1LTiQ8yuSUSGu4zGairktGvm/nMyVL3dK2CCIjozcfcUOVbTG9dE1gZG2Huo26YuRAqWnc
3SKPAumMuT8IqZ4QSEhyX6jtnLz/p8tIZmkygOkkB0vaxHvqi8FwMvJVcZ2cAFZLiJJORFYNfpEN
QnpEaot38ogKaiWwEg8Ow0bLBQZWHwLu4L/pTN64PMLKZz4BdW4rqygQ5TYdjfN0ybdiWwZ/ORis
LQUH3NtS8vQYZC86s34AyNxJVx8QIVBbA4yCnTqjx7VxMYN3j/Lf+LSLMq7d1hebxJF1jMsWOBD+
6CR7EFv1bGFz/8MkHXE1OvqKMoONZdcOB2JQ9zhbASw5aHF6rbSG056dC/0L7M6hjKvDNhbwOUfQ
1ivs4Qmn2vXS1WsV4QGnixsjrI1w5yULicmDExl/2ZZJ0VcgCmCafllf8pmnnUF4Nv+v8hEOwkYl
JDxNuw3hd5ze/voFjPipgYqxDxer1KNL0faWPT92MRuGgqH4V28XCjen9DRBLdxXbnUtJhwlRqD2
9oB7XwqhzDgSbvqI7B89P+K4t6duppdnoUldCuU5vbZyz2KRWQw1raCVwvu3pHQV/aiw9+pATgt/
yJkGtPvNgnBnmJGIuVblDy4gPqR0FAZ0Eg8D6xg2M0WhUGuj89uHuFNlRm2lpJ7PQge/aA/Mi1Ua
vDNt9T+Un7n+3ME64O+cRwnrzzP8S/vqjYEMU+XyocRPOX5l+HwpCmCoIKUgk3+b8R0Xlg/hOgCz
CJZ/MJgq4lQJztWDropclf7PLhklCr9bm/GG6eAkyc675TdVTg7t89YDvbVDY7eV35VBdgxeo6K3
mQ3J4u32N4CsZMCWdJghcfLFCR9gdMXjNDapuosYMbb25G8J+7ZqOhBQzy/l96fyGwIuWiQ57laI
Bi0ltOhwnKoCW9/053DykJt2smWtt3+OfMWTBbvgylssjNUa21gp7rMetmhTd9qyWD0nOg43BHm0
zG2uwwxsfHRlTy+2VhMuocjyt5wnOgDQgXkNySMFGt2+zqvreYwthZNxsxmdi2D/YQ1cMV91UpX6
tKj8C+SiY5IVPDcsz0p9lALMXm8nnabJK6VzcQgGq6eSkWKnPssxJVZrmukwtIUl7t5B8nrwZLnQ
SzsquI26/TSoc8Ygth8R/UQfT6YzTPZ3ibDX+0Z7I4CpZqRYO+IM2yZ1rRp5pMNiQPR0UFQmMQi/
AHaUkMfPgBLRNfQlcg/TYw3XO4eG3Qa5bJrL9A0PDFAIzB4bGiEXVttRXNorYJTNRgyf6WwJ3bFQ
LkUEM7ky8mCtdo46Xmlm3+iQtkpiC9qfDnRmijKEC/o9GEgryyHCYZ5kYYE3Tblkt0wOyto13/3b
crMEzuDBMO4skmJXg2MYS2Vkg+/FNGAcUOD+S9VuKogQHEn/4CNnZWGj1w6nwByj3jaSOebHFqXv
OXLk5UYNVm/H+V98q6NsMrvie6vCFNdFPOH9PCfwhqlsqnJ+itiJjvnq61Tb5oV1cz2rkvZAGRLK
jPfaFAd5j+SWLiXcPXuWrK7f+dbPJ4Vr3VT6Ofwuu6QPIuvdx2E3rzXdC+nIDc1xgpRRD3CAIkLz
iM3m8xNa04EjjTp+XF9jT1r0QihwM/mxStxQVjd5qoRHaXSLV8gXwJZZrLqyRvupZJgz4ji3wj1A
kgDIiZjfPw1ZV+sG0Jqpd4+v5BJ14LDguqJRv06bTtUJCEqyFeP2JgFJcGRtdClYXKEHz5c94Q3D
qVfI2434UUzVjZfhiYaugok+fTjRI6QvAfQrMWqW4Z9vyz55mDOZHzY1EEVds4nre/zEdmPPlJvB
vMVjsMVbCqxuuT+viXfcUbh7ESR8iW6e0z6a/pdq5ApPvwXzZ/YcSDrNgu3mq+8Uq6q7+HRQ8ciC
CQcN8YiXpz1HkCt/BZZCxeTo7C1GRGnBD23495eM4I2EuDmuLuAOZNVy+GH8MOHY/c1OfTs8gMj+
43eu+qhe/K5nJ1pfCwxgMSQlPNP4GZhnh6VmltyCc2f9Fnchmi4YDYnxYtRBEd6y43ctpBFEucE2
bTw8qw42Ao7nb9d4Q4asQ8VM9xviR6+lUW9eLur4tIU7QWMSv9AziUmWhsoHEf0fOyDWX4lC3LTm
ORdce0JgEWCNUvybcQdMgZy+qC0FljjzA0KWV2KSKOHOcL4tqsjqpIS5EcgXcswbuetKdMHnhZgl
d+1YlATleV3YluuwGcLs/M3M70dD5lop3l8zANwzf2pbr0bQ1tTQu4HHX4ejMnSXdXl94EZmZtFk
tyS1o8pyCMK0kgA0Gvvn8lBsXBNoTXQ0zfKGg+qUFqQi1JxwxwgV46ZCePzK+gnzX94xS9QZzw3Q
vIb+2UDW+vMoJJQNmplCq1twFDyepeKUUu/7sd6Bm5t2RBXlWrh0fh/lkn0StlWXTm8Mb6cfNBdr
pg9nHsQGWZiDMUT9JCXlW7NlxcJUVKR1JGcg6xG6uQ736ejk9qgtxZWngc/C2iJd6C5QJMv+pW9O
qGQiHMLX6tV5vyxsEPGca5G3Qb4BEq8q6rD4lOIkjzihcTxt/t/CAR4NHHc2Di04nMaMOS9EdlAW
PupWmUNEoZvIUfSCaNZ1YW5XBNvpGYBi/qpzPIDqMeBDk0xa0r0hwpvQwN1qvHe8NuSpE+uyWKcW
XIA/z4rzw5etbe7EZ1WCTh++j/IdvUiuzr4wKY4OoLsl5AQn/p4OauOQBRvI5X7KH5BfT6q/KXrF
9lbc7ADsfQ9hGG6pPUVxqvg+L7fHdtba5tBpb+20hOyl7i0rEyPcZtIwPHKNp2FT+TK/wadCgP1a
qya5sV1keC6rFCh61KWMfI6EOeHrr8yOPYL70pO9itanqdPZQ/TWacyths+Ar47S22e82rzrRzu9
bjymdDRCPJvv6pwzbNu+TLYxFObVSPPHNIrTK9x744EdB8ITQk7zdPx3eZ0yiZDYhj251PZ8rvJN
Uv+/Ib8exdWVnJyANljPfWCzQ7o7CpM+2mmsjLlhN+uC4Uro767yhUnlIzf2W22wRlpInWRWkbYj
2cPyNQMbFHkS2W4Jh357mRtQ7I3ZHfP7bWoU2dWh+xMAQVAn3j6Cf87ursS/7QpE4RG4sWhULjVF
J+8puXJ4BWcVlj8G4dAFjqSvXIrFIDInwCu+wKX2HwV29ijIpcOB1OF/QEkVlSR3eoDFCyOcN8j5
a5YQwv1cg/Kt3+pHNmQht/2IzDFDTBoC5JGRxm+arm0PeXwE8ouNkFdmqICyRwK5JXBupLEE0cTH
jmBgDyI0K3i21GN9BldHh80Wy0D6HokDnWrCwCA1GoHawSYI3oml68arfgUwguzUpI8c2vPM6BBZ
1rmsMvyT4sNIK1mpS+PF1TJIwLC4mIkihGKHpKLLHbAok9o+IVtXYfsheNPuJn/f7c6YG90ooR3+
aQuJKMnIKd09uyiUTV88umUIQQDY5QYob12Y8xc7+jtnFyqHGx33o7k+FfQaU5Qupv2gYPzQ5G33
wT1uZrAuZ9P2awBNqqndbm5mg+FfFlK/ZYs09xvHJTlYyfJoGI9pgndvQAynPE0TYedemoJ1wIrs
qgYy4l+eFac7Env8CDmLJXUK73vVGiHX8FyCUmPCaKATSH279Eo2w5iMWLz0FgUcX5A/bVsY88v5
ZFzJiNUXvPNh1gA9hrW+mAUTYBnNEVBBsQeEf099Bej/la7aj4XIA0r065InxZbgUz0SiVtuWVw1
UJSDdBHSCN6qoi3mxUtb0r/aB7+oEvUsAMpygM+tn2ubuoLmaOmayxjL1yrbf58OeP4OMJrtkFe3
e83sJ0N6KLF/dao/pPZaj+PqSlgBMaKKl2PVPHYVgLPidzlF2Q6tp6MqmWjZRjlNC37dm/Oim0cs
D4fsMHChj6SB4N78ebe4BnKx5NF6VMOt43GI4sbZY4qcpbwS3LdyzoEdJdPR7lHnGAHnZpzaCFnJ
YRWOWd0252B3Ar6pK+/sfEM9Ouyt+JPdai5CT0yCtXBSQUzBr1kYDsWCjf3wZvk+Mb1bZDrJxqJU
IZagYeLo0HMOZkgP2ulp4sNQHklPvU548BUB/bGrMHNVpsourewe23vI9SiTpB4PCsoRAznjAQQJ
wfvf5a1YTQgiYUwIOKqc42fED9fISV5j8IYT+iPJO4iBhXk17DvY/VSfW8MS+qBoarI8llgZcum4
pt+cZjq5ykLKkcCa5iXr7yzZb2qS+XTRgaZvJ0esZXYOkXKKio8AG8t72/FQiYdPNr+kWF2IBixu
Pz0WwK3iszWvyObU11i/BejEvBhzfHsTc7vanAuezrSDKBTDG0sYGpWmzcNszlMSBPeihXA6H4GF
CfkuFJIR4r6yEqXWiaGfNs9BramSnm45+X+4IA6e7ooT1M8nWh1/KoEJyz9KPoDup1H/sS94mkW4
r9RLgULVgoMU18YFAOy+hbbAyBAQgUwsNkXgtnEFtI0U8uHxGIcfdkw/RQqShLP71ggZ1kS1u+RG
G5EYzt49z0ja3pm2wZA9yW4mwxoSMZKteF5WBQO04dhx6H7+6hzbkYluyYYFGgeOjdF5qvZnpDez
oI1R9GlpIWk7IrkKgteSfSIgj5V/TLqIlTvd1SAZOOgSrC1O2cP5Rt7ci3FjFLU39eJ+gxc0n8tv
bLqOwTnYnkA7HRy6Ed65lUWipNlDbDhOGgAFbq1TgnRChSKJMjkg+Q1qjpsWawYdJLu8VcevC3lZ
lyuG4oPRc/7Iymh257R76twT4ZVhNTxZtJiIHFNPw1xbWKO5TmV78fkLqt/R7JuHy3FbdkBj1CBs
ERq1ZNthG3H6WlPlJ7wDAejCB0jQTcb41iPWlMBhOjyc6+S4mqtomxFPlfhRvCdA6zDo1u7CDjLI
yC38IsttD1EILp0Hf/+TrlOT7co7PrMsG67zL3OLjBoI6wcTT8WSM7JlPxqrbeBvfelH8gb6Ji4W
XZS1cNmIJ21oxYBbJyy1lX7s+Hwv7tyv153arIa5MvaNj1otrEe2mQG9vnEkPvgkN6rMaSwGOugl
acRW3AfYO7324koEMSvxHs/SY5oMbnqdXMHnIzaRN2JIsXjA0BTwkKtLPDeuct0chRezstVn/joH
tL6fHo6hCAtqexm6vi8gJbQiSZgWvuv/ACM4c+i+LFXcPgN5Bwg8eoxGcZlwICVVJ7cxx8SUqOfZ
LqZqQPH+M5C+i/tDcJWbht6muSvQjLfjCqFdLPCbDOS7a2Dw6BACgpU435e82D0PgCzvmtjdQgtv
/jvfUO7F90Afn9uT52tnbH8nbaPBUGIICGprEfOIBfxooMvg4wlVxIqXGbKZChD4wUxbXHXcHOJ4
/pbdw+MjjBJ5XqxlfWKRd3CXje5yIwALdH14+F33WZ3Xwo2nNE3282HiXZ5fLnHxXNxsi9w1+njE
zZz2fPAYgKrjsvcRMWIF5/iwKasE0qbko7CpQ9iS4rB7F+L6rM1Zm1rKldI0EgXC3XQ6i9K4F9y1
cHkKnWzQmQAtcz1nOwWguQGADUFqwUoWL8a4wNacumKL0H2d0/kRiZ73pwjsj1UYIDww4QkLSZ/C
Mq7+m6K90a0ZPEL1Lj3LxDKK481ygYnW/odHaCI4b8kls20i1+klwKd9rj+YoVa71H6JBZqfs5to
OuuS42HPLEeK6VtJYzIc9kdB8d8VrQof3PoI8T5b6SMTcRLVNvZNaqhYkRw+J8qqWzRe3U9GZfCz
nOncfDpBGop5xQ6oA9izap6AVMrTDU2CLFhSFaJ2w8bDRe92ohe7kbFGYwcB04HVHRNq6ehaZ03Y
S+lXcdR1X1RqKxD9+nwBxVGya+33x/qg4R6fFoYSgBdkjaKub+UFdmc3vO7NW+av6jfp9Ev+JngF
Q4WDdcJhLbEtk+yebXuOXenwwkXUGRhptY7yNlCuEN7TFpuEo0ZnzftrOchUBIqatfiLfPVIKWCI
aYzDjueQKcbpzyNXLGjNoGC68Cuogd2U1KmgU8/kKjjjCzJjTjB8writU5h1/LV8S1UEv7RbOTus
AgAcTCLyvPSdWt7G5kdGqJoNzEXSQNOBWyayLSCUeoRXA4vmHfOHkL/Oxr7YxkFKLYashl36xvlw
+NuOc1awppBjybwmo4tWaJ8aKkjQ/Y0m9mG6ml8Nqjnc1IPwhOslanCAq2bWFdZ7R5ew+3IDJLX5
tPapCvSvNvHT3r/uRQU/baCY4EVQn4fqcTMDOYnbVs0FggrLxbFlTEVACHdI7ugknB067PbuslaL
Qk1JynlusZ2vz3Zz8F8gjzhY+Ppz5trOK6BowNUp56sZ6ACO9cCgt81t5Xu+0OheKAc3rAStGehr
lKGSYg7A8ujztC5q156UD7wE9+L1h3elCwz+WYAKtf5mOhulKaL9noGOb6ukj2spMrrs3UQaUSpE
xgvc7bsxB3tk4SR0AWFjzB9NRdVtgmq+w+CHvY33bDEs1FIbs4QPgl7rqVjbOyS+1KwtYCdeaXpE
1Vnnl/iLmsNLuLhm773kRMnXhzxYVCoG5sbXE8LonPwwUwqQu7TXOYGy5VZ9qQr5seGYRNr3Zynt
4mQSnu2qyY0vsTI+8qyjNYo9S1kviTYf4WOemd1HTjDFXfjfLHOyGizM1D9Snvf/mSKfN0GNOQo+
hm4gEWGdsFPIdOm0NBAPIr/19a3/rBILbTtnG+zPV57Uxm8GC/CFCnaXnymIv7TqeQ2oQTBsbCCn
gAyGkmSgpC60hfSJUFZZhCcEiCMEwNEuVckxS83uLBrpTWlF3/48PUSbA2pd0fua7tRaW4HqLb+c
OkREoGg0lQuSSlKJHFRFGXtPDBwVzZS55Bu78JYOS2cVPZAOckrrQLeRvVEVExXBXM3gEX9hmCj6
C77N1mMnliNEciPRfn6dmYBIBtueoexva0ZHx8wx0Hd0jYMjwfeyhvwBgPGfXNzN15YFqji2/aOv
fSSIzz/so+d3nB/9V0qjPXSjeRnif/2AJbpWH4pjQS3MP5zDTaRcHqA+2EX0+khtLA7mUWXyWlcA
5H7ie8JwBw1xwdUAKmu9tDZh4yhC9K6dKno4mI7qL0Dlz9a8DsrjJcIlFr6R3q6Zquks7mzPbXc1
G2zjkRmpTuH3QZ/veGoOZSEIrwyrrJd4e6vPRSn+BWTyoIgwww0YYVX6yX/5jlXcM7InReS6CO2I
mjYI2duxZvIfnR4Mqb7o3d1WicGR9gjABxnzSyBC4U+Aq5nYvvlpLcDhWZ3DR8j7Qrkgklu55m1S
DmZsroyx//1fJnaJG0u1xF2ZskKggHtgI9i8FYc3ldAZbcP1tx14afnPUIfLcDenYv8bv0BZqUg4
2xQeY3fk/7SWOqcWEZxj6i0GicdzvFO2EOkUUA+7aIxGEaZe2BmUtgtxh4akDH2i2UKADc9vUOqT
SNYsPSRNvUXM11Gx8uXKP8+thydEJ3Ot1X6vNxuZCCziAEwT/HkWnqLB2vdCqTs+gxPeNrCGzXoL
YW1zo0bq2SS9y7fD/G9gF3Myq0FPCv9WvgMoHBa/t1RTHrtII7ySLICRz1ghhw8xOKa+vG7dc9jl
O4/hFhOc22bYya5kBvViue1Jg0+iDkWKW8vFiTT2Y77FtXYArvmsy5fge1EBzfC8Eq/iZQPhFZ+1
tpMBbbvtmrx/FtKXi4fJs2SZjXLE57unpMJbsNMuGc3nGHtFVt9iv7+hl2DtAa24rhSGm+IKSQOg
nHBmgPDlzle1QO9w/6a6nP4q0AZ35D791G2BNuaUUUbKbGlrbNQip5XPgRN0v7xZdfd9Lwf5nEkc
NQ+IHyNC/2c/HZiYl8nT4+VMnTfUbOoEKlCKXs4sUCysSmbisdXda0x5l5dAumMy1eUeA+wIR11+
B4gd+OJusPGSFYBnnGgpfA+DnyrU+71GR1ffL4aOlHv3ArLzlY4u8N3Pf51OQOXftZp7recBzYZy
J3ATJAc8X1agZ4E5KNzWoF6QH4M/vZuwcovViYIX0VLSkXwPhC1f0WH6AL2ptlgBpvj2JqDUkFed
qa8VGsvrfnXGqys6atfT2S2cS+MRLnhMhj8TsGkikEn2nkm+lt6k3YUBGkKNPU9FwdbXMFXa/Rcy
LlmZqTPQmFMau8n8gb3JxAk5HF28DDthTdL9xdcPWZgEbE21tL7tuzVOKSjFy6JRx2bJ2++5u5n9
A66JLLYGCJifEdaQHRO1/+OEgKkFhGJMHtrxjv6CvRLC+VR7uhIpadzPAiF06J1e8spTM6GGJogq
G3mSZ6OA7QRs4w7p66m+Hyj2a9zc2Ch/6biV4igwz2gCfJBls2bkO/+T0E2HkM/cmdyhSYQ1Z7hM
QdWgHVngWaAL/69BvUqh2D9B9oKNH9CoxBbItsMfipUSk0aV6DF5N3eKUeBa8WQXO34cqdVOZmoL
yazhWK541x60oRPd8xFYwUX5tCpGHSfnREPoAErQBGDXPg1VZ6YaI/BbgyXfbpkEfR4a7jZqQ/eK
vV1shnKOm+Dk45m1L0saxw9ltWDmuYPLbyUmg4qY81NoQWj45K+0Ge9wEIefayg5WUHGS13oQ/aI
fMuSYHp2QtNCUSD3XSHUDtOOruRbUPU0+JxhoqdgY0zwcPaCBqkvpOPq+KgrRBkMTbp6MBHfzSpU
J7uWpUM4yLFhVJctyJQsZCxX9CJ9wIXCkzabFXswGjbvCgc/ubFMkfvtT1VScDcmIzus1We+WIgs
SjvZRPgY//pl4vfuGOe454QGZNwn2m1V/Z4tGm0LKSFoLX6agUCz0Vt7OYpbiUec/PjRQHLFbDYs
bNKAWGGr4e6G2CqtdP0IWqxFbam/vFkUuddMfwTOBkk+wgTceJNcw1sJ0At9ZPbSxRoqAFCjyMML
ZI6xLWwOWpTUT71E2WZGp+UYM+k8V5JtPcXRHR29kTbBYoIDyQAttd3tIMwB75ZTaFxG/Hn1Am4i
9b5USQRa2XyeGLtioraA5IiO/7V48e9PPTh/qGq14+xiSp0ujERrWMFXObOrMjUDqWogEZEOyhfG
YFQDAhCHyNPEGUOIb6NcWDfnhRmcHoSVRa4E9RwxirUrJjgxCFrVN6knsFhj/YBGqaNtbnE65AaT
y6jpzt3kzsJ0YYkvnp2elgNCYQHfleyqXJAIrug/mxU1CvonX0o4e3+BQsLBHdp+fj7rE5jFV1Xx
osf8fX/l2HTwTxMv+vCMmY73H8wP586LTE2zETYhNxX4P7+O+vqHkb8Ua53EkEETbuJvsPuOyejt
xS7ASPb1XMcQ+GqewwmEvpo7DWtZM8y2SYlBd5scCQbfm2VSamuTvfgyla4nIDEtkRPwVX+20JT2
fFxxoGEyGR+33bQjwzRizzKbXEvXmqDBz4p+qprMyFson2Cgpiy3z1h52IwckFUEuuWPlwtgmOo9
5/frw4deyCfixlohpaF+sMCAnXWxFXpl+P/IGjK90o89YtgZyjDnjs/Ps+OwBHwNZVDhj2x7j6Zm
jfG7tgg61hUZnKv/VcxnFj5yNgyjSqsY9I++HwFEfLpZ4siZYfSRe8mzTomnqje16suapqUUmDBe
yS1s9kmEz6oqmLfEaDtANSQMvG8v08XTg0GCT7GyG59CC0Ok0OFIiJGiy4772Gp+0ogTCEJzeY66
gALO1+mQFnp8qXT2A5TkyC4cFzepl8HmKKEL3tZW2Jzl7Z9kAucjIuuEmDfhC26WQ/R5zCvZGH5H
NNJ6OpvgMeoZDkyjAvmZTwEAPbddRwGHX4Br5UBhaPjfjtn+MwNEDj4BCMiyZJEyKqb+1bpasCbh
k4KRWpSDGAM2/gGK4UCAg4RCnuTet7AkjVPSFzXC+RNqtfxbDrwULIgsUZOThuDfN1AHF60Nwq8g
klwrJh0OJwjphW4q4Z9a7tLJ4QhZwbeSTReKSb1/hao673zRPVQjT1Gepuugmuppooze4HiLr9r4
JE5v2tSwJyuz82aRws43RlEHc52riseQZ9WkYeVC4bBiRbJkQ3cCm580mrXbKVmFOkMr8bZkfEd0
vfLDJ494iTQNrNmQVimxXNVdq1KNvCt6LSuuU6Fdqh0ATa1cOhzVPv6yxPyHXG1uAMWkBooQBjwc
lDKhlyhekoDzaDKIlOsS2oajoEaAyiIfkmXZdaOghaASlS8B49293yj+KOEpfui1LuT17+zf8mN/
BdZhuWXR1y3RVePkfZFjCduvcqQNk0IGcCKgNNGxHfvG+vcO3eDOy5jwppYeo0iG/lXtE8jkONKG
jkWuerr9jr5bUUB5HtdC7tUsVqSj88YzOOjsGHiAKV7Tk5UReukCmcLVmybSqgnHzB6L3dZSUb4I
rd17zJeS9bxCRPiDkDF8UJNVzZkCOict0BpvpeifQwCjL66S0EP68tGXwFj7t202hb5xz9O0qAs+
xpMDnyk5KS03rKYsoyB/KvC7pUYNxminmjnZ68H0nqv1+CwslZqG3ap4vuShro7FsC82y8YRxHcd
H9Z7fzHjaBlFGFHsCD5dlgJOLbo7wQyGuJ51AzdFdK+ERZnH8yBmYnCq88KjtpTIiXUPTuaFXo/z
vgh3UwiqIOvD9tDASv6DyroLfNrxphFKX2NPS7s/vH+c2S0/ohZxmClKX1W+pd9+CeWigtXGyWxz
opvoMCg7GDiZ8C1QeZWT30ePC2KvgVp1wixJnHZLevQgtn/hJ8pI4AAS4CCRNe8C7d5V5B7jceNm
Xsi9RbkaGjTEhMzOBa3Mi9T5TovLRT20JRiqc9D8m8n68bovbg3JLuN4hLGZ4y47dqxmpKSSU2U4
FYsB7iP2HJQYka9ApXgK8TGHQMxM8PRrQ4OIte2yVXu2VpMDmxjTiZLMSSxlf07he9hGQmn5uLAp
IZMXJaQSHQkwR6D4tG4DSmui1yQY5+jbvwNkCn7lR59fL850FzIMfxswY/48hCwalhgG49z5Fd2p
l8r+iJqgJXGAKW/6BTlIPOeakctHTFKqCzx/7woqokBJ4vjjss825gDbNW9zt3O1YpByZzQLGVfN
HdeXBp40oZNuyNNB2EMMkIw6dYknIFbYEADmZlSuUssPpjubTM8y/sm+5Wp47N7EPwxJIbmrqHxi
WG7UXHgE04rTKuPIr0ZJeLXfGUG2SWTt9NfAe2aNOuTBucJ9r116xmQnbvGo3VK7kp1VbU4xrahp
0eqcxzyiOoRqhUTeGmeVtX/MtlzmsbFu805r69qBnJLqQKIfLZLyGtwWYO1Vp2afCE+rL/NrNYGh
L0Xbbd+OIExifDtauSpwxIOew861tAnKtWg3sOxw6NiOl6OvGJyVPz3p5deLYwdKYPgpj3T/M6oM
8AoDbRBlTjhylGujOG8ZCAPuJzROOKPeuBWo3x1G5aLifKtrxL3hceM84Vc5sFOhZCTDgrGVXJoz
kKMHUcLyYzcOeE1XuOBOyYNteTkBXXQMk9q6bdLYUrK0FpDESawZS/0g8T5EOhWigKzGam91FGQx
TC6/KljgpXXQLjSBf52lt3diY09kGqG2t0ESpetsKsaDKbHoVjOfz7CLkMvKGCdtqNK2ou+tXpd5
jkFZFgJ/wzYmK07nythApjT6oFtBYBSHn3HkER3UolnnbRmXGNMnV8aqJQAWTWOvw756WH5BXEHI
oNVvQOXC9/syBPNP/C6MxEtBfqrIdoz52BFTt3DUHft79RMp9LRGCW0PwWvQ/9UNH6CWop9B2yLX
R/vPfjBn1RYxWeMe3HSMN03rLGucSCLS7LFXPWQMM5ehr5lfdmqN08ewXX0VOVZnC3TdOBChaMGr
E0Cix8LcKG1WIsqhiUbAYxvUSUqeLkmBLB1VYelCOP/72jf+8ebX6NVXhEbEzGp7jSl8qn3gKBzA
mLcxtB7thAB0lQG/pcPzknG+Y/SlODBb+Fzfc08kniKVxh0SMFF05wVbUeSlH/WQ+thq64mAwciv
EcAzy/TUj98+D8lj7wb2YSXzoOM/ZGz0XbOz35ojcYQTXOspxbbs5Tlovu2iYREzQfVrqCsEZcmg
QwcmUjzkVBwaesU2tM9NkuBMf4xREYVBC5f/6KbDatIgTDW9cDXd3/iKlBpmW+seY3cZXFp6NanC
m6iJCWKJorGJi8lMjwHuv3FkxidY42FyHAGUYBK5vXjnLngJkEfbJGGI149Q59mc+6v23Kx2Rw2J
RlXRK8QI84Y6tUFrmpgarmZNlhe6rE4RWBJyaTx4PxpPncNWhYimvxlNSpUgN472VljKshvHPAE2
Q6UvqxY3MQKrhBVe9hUprs60H5JM0l8nqKC6RSZqoxl0rtBanWU1ka31mLxe849DAFVlrdXvkDPX
ca3sA5FK7UlFoV9SjHaDH78+2CxghlCqdmV1Qwzg/ImQThbllB1CipWTwKgGE3GnCQC7Fg351xf4
ApAeIYvMNdCEorqlnmPk7052iBTUQKv2h7+byIjZhys6P3Wm2yRBvej0iEK+3YN+an2Q3t01BksV
FL821zLMwaYK0eyfP00s2XxGSQhtrSBPnOUnfCmx1BQd89VgPaR65C4tpLhRfw7kEkCNzuSVi/K9
KjHAofZ6G8aYNeF4JSzmiGtMkaXpOrTC2GFIJMioMMEknrNZMP5emvmgFkeHZzfNuc+mfwLA0qNP
/i4b+j7WYA7gD3Up0SL8eLxMloJWgFp54Zf/N7zzFUWWaj0fqKZ7FI3vyPFFhXNJ54anXJlHF9tj
rd1utXOCvD0MvE64UlCWeEduUQ59SLWvQJKV9o09aFGOzYz5WiYNEb+3g5bqvSG5tj0J9pmLhBoe
oyDNZTNYlNlmHfkZdWEBuEH8FX6NmH17205U4T7bwA/iVp0pfD9Cy2GNYxSZRw620HK1N9NpPTKV
Mw7sxj66c+LBrS4hiJv/v/nx1yaIVN/zQuWH6l1sPLZNv2wHair8bk3DK33biY4qD0s3HEwJRrSl
Ky1WZioShlTRkSwyZH3ypfkC5J0yrbJd1E5g9rej0Ww1nn0qXrCZAC8sDIoGRe+SZ/jZa0Guv41X
/RD30iEdnEttWTvZ9sBn4uCMvHzZOltPZADjwjow8Z0MmEdZFaC2UM9y58/oluA0SKMpd5a/x0ch
+8w/rvKkYIxyJDcBp2/o7Yho5dA5iMXVZbyuHNVomuy+r8p3KFDxSC3VD1ISErZ7CZLmKIj/PatI
j3jE1PfsuZR5/NhoVwoCJo36/+mDw4F9Z2fhtQEAj76wqpfSkSanCoOpl9chfhciyh0IsOwWNDfi
tM90VxrnIaCBx7/LPKiceZaGqbrkPVGFtiusoMRVD8ELm0UchvekP8EzGggvHO190XFJvi8hTikL
zt2YgIf2XfuRjn/fMXED7GK667o4Mlq0RG+HZ4tYY7uF9cVeU0+hvkHDKF8GjumQoHmbSbv+Bt3/
ks0eprL2PvpwLCmo+lPZlVJEwvmazeOP83jTLjpGsjyObz6PzfwaLd+IDUsUcTR0E6jqVt6UMG0v
RjJ7qudfYM7hCRkdwjnhG0P8RlKz0DmYR8TZKiSuXzFUlial+OzCfCAQ162GXdQP1VbjJOwth9Xo
4ZCX0wacnUKV1o8I8Gz0CpMk4L7LQqBUCgtyYtapBmNktTkiSeiaDU2aflQpcWpD201+WU1gWPcG
AnVI5FZAz2kY8ykrxUiuRvM7Qm7WMuTspwhioy3c2GN3zeaxUwvCeVeyiObvLDz28GdLoP+tLBnq
oaDo+VCqQlonOR3+/6rSIZU09KTQCWxmwWXPyllBuLHRTv7RGjvNPOUd5QkDszN0WBrt4Y2V4pKN
FX+flVfUHLgeN90LH90H53OCEt8YQvnzISAd+VfLeMR0SFN2/QtczptrVL4DhOTvPVahsX52Gv4W
BSiAlyqWKV+wAIZxkoDvU16VFRYGjV4KSTOil0A6wTDUDWeWyw0NQ12T/WBJTzMrzwm1b3ERbuNY
zOEzV74S+cCy7CpodLMbNLLnoRYjtWuICoiYCMmGvYcNT1+YwPyyEMvKAwR0NXhQumLt1vdxZVq9
lq5ugeD9ERQY1T9w4u5/ylMzbh3edrD7kiZs1iqDbtgOkJA/tCS4JtS3cNa1XO17vL8APZrNNGd2
783UOzm/6HrIgVGHkYgyj2g3HdGi5X5jJLddcX8SMSYBZ17TtRSpttdOpqplHacXQJRTJny2DwGT
p8c9zglxoYEfXefBphxMpEFN5Y++SLM/L310u5HviBgxIaMEnmJazAd4J13ey1huWWo647gymwt7
kt/mGqAZ61G8Mcf64s+CmxvQpTORkRb22ThPW50njcAy026n87FMaA9vCCiQYV7tjguVvQlo9xZj
vtWaVGqzbTMl92HVD8nXmWX7MpWlWroq6Yf3WyHr7zV+nMFkBwSF/9v1XltZTYu5ae1wVTULBzi+
agNrVO8M1UASu8+m7ef9xmLGJYXvQqypPpzrJ3iYi+2Pv4ba4CLwPvn9a1lGVlZiC0zb/bwwcmAG
VJapJlnjAF+ayHHU8cD+C752Cz2o/nT5UVR/FZFb8IXAdmOq5wxM0KbslBKITYKINQofJsXtJH/6
eLtlOAvp8m1IYupoLAw/+CQBIZFVQ+P9K1P9256wUCsDYEDw4cqw5ZwXgc/HMj9o0Xn00oxLaMT0
TlCuWPu1O+ihkwMdHYPtNXKp0fSRDyq0VZpxixmaeUNTgnTVQtLHcMydVQ2X5jghLlwcBBOdHKkG
xXjibqgEZZaJ8wuL+9i5VmD8+PsJuZrNBqKe53jhiceKTIqf2gVTHI/D+Jk7/oqPVA9N1xX46QJB
fo2UL+x5COX4n94LZfP1nHdSLAJzxZ7qJa7+KnAj9gkF3FX5+IRkfVtBlLd5okWkOm5NH3aVMn7S
m6RM03MG5NfURU8L9zm20cEUgpa+UsbpcZcFlz9t2q49yUv73Lj1EhIijezqVV5l5LzVqY90dmI/
App+Su1O+qRQuFmcP3f2EaCSoxQVsQWNIo5N3fZEkeFrQ0X3A0Xxsxo81nWmxx1G8r7UWdzt6tBY
OzRAdiwMAGzEmgaUq+dhIcV2VRNO70Pv4wuMOw3RtM7ocbIPrf4ZoAco5SDh1qlfOfrcnIQFk/Qw
ANAQtEybkphlooc/zpEeQr3cu1sc6GJL0KIEwHZRSLk0lFZXH6ZQFqGwbLZF3agRs+6iZN8PTp3g
rYRwZHrd4/hhlrAlTYigiKZPKLp72xVPvajSXn1DXYiha8pd7Y8/dgMz3pA4JPnk5Fx4UJjVg2Je
R0KslcXxCIIivWN9mE+6svollmXtfWP+usd2wG1xb5Ua8aaqJsnRpYM3nOcLkHxvxCbPXy6wP9Ad
fxhk4EptBXT7q5c4U5yIHe3djm5emGXLOKK4f2m0NnDbKBA295LHawD/5i8zkBVUzrEbPwq/qT/Z
oBcUylJTQCEc/lCvivJk6gU9geowmlwRMfL26+0vpeSML2OMZGlrcBrCMZRv2vcC6cVWsldXOqb/
EUkttUsC6bhUzqhmpIxhfKJ08Mx8bs4XKfzKd8pwDdI+MCNJB3u1JNzxCMDKbxcQoS5FzGP8hG1+
N0a7fyGICyF7NppluwT9Y8CrdTs/xt7tatv3x5ZS6tS2pq0E4Q3kimA6HZuIWFw+JCKGA0rdJH26
E8R2OIsPAZtjfhBrl+6tDIGjRJxYJGA6iheWckoe05HyMZauxDxzjfE5dPiTYebj4/MrGt/xrEP7
/YrVyHUuxhxvsBHDVAGYWmtV7VNsUZZjb3HlNl/F3dp6RYNiuD0ci9bPWf1V1rwrqNmue3qhyAPg
NBaRoLYpgJiXTqyg1G9xlzpb+X6A+F3PdtY0DHuc3cBdnvIq4VyrKmGllokUM06ovPNE3eDjyq3b
uRgEwYwr16dTLAllOE0RQZ3xBOdHECTFb0XWPHO0F4LaATj+Xth9OVLgPUq542jy71qoLQb7Gd6A
Rups0bMPHe3quqM4777MheBpWM7s65hya2wT30QBsPLUqChb29YPkvobctKbX8P6tWwM8yvjD039
s65Kmafwdz1uXzQFLMIQVeP7RZH0rSXRvMjGvh0IV0cenoLzW//ZApa1vDhltiL5w7kGqcLtzc52
ps3k9FWRk3gMCCu8K8lldEMycGK+AlfGCVq9VbSJc+KKG+Aj8d47XLCn/UngmBg+sbQ53u1ys8kS
vS6jhXOGZviLkf50/PsUTF6KthVwtV0edYYhFUc0MwzCiK5qx9P1V7WxKUIz90GugZjS4WDF6u6L
w9BWKKW0Is25+8YEZ1LgRsrdkADt0+k8/Zl/KIdm3sHZpB+BM67Wq2Ha35trqfr7aBZ6Gyr9dRTt
VE9oEENXVW4Usn1S6CW4FXxJMCiHSAeYu/W1XVBw609wBe8QpJGdpixQ89nhZHK9XqXMj9nB4Kr7
QK3Axiyij2XKQRuKCY4E6RoF1BuH/4WPyze5Jse2Ia4E930upTsX4Z/sotJmmj9lEWgkRd2bXoLL
5wKfBExrRVe2nPt7ieIrDoWbcJjk7k4JnpFEJBVu8YVTyGnmpV5a2rX7HJRTMAYwaXjhoq0ps4A+
RKzkgh9JTAVlLpGedUM8nG6K8ExbnIvX05B9j6CiHH27x1ePz9+VEPnSA4/wspya4M6x5ROWFV3M
3nBqig4b5eSV38PQGVuMWAyPRpsTylxtGtIp/cbiLxqD3N1U1Pk/oAmET2yKY+EjT8svINXIBFHR
S5hX8CX/3GCoEhlGSszG90MKjRg8Y2fpnD+noUITvVX98n67YFyK/Xs+bmoBqr9FHB2qjnfx7GEh
rBkb2pK99XXIJTRdqYx+NqkYdy6Vr192M9Iwii2fk0lZhld9muTGltu1QB7Sw7iIHfjqR0dmV3b6
igJ/WcTruhqG6XrdO9YqJet3r8opVP6/Pq0o60vQu0w5V6kc+KlNRATdk629xt+YehGBsguDJ9hD
Sw2ybUciBeIzh9bGOnwhPr0bMezeqvGs8MdoXZQcYDJGC7vhJRQQRHDGR9QCoIg3KIc9xQtg25m3
vmLMTQAuN6AYbb2hTc/DORpDJ/OlWyPg9txGv+cH7X9xKtgJ2L5C+eskbVk4uTaOsA7bpczna0ML
jDhzpPIwAnn1IAYkrbEnHchKUe3B0I7a0jwvoah7GAMz8BQi9CNYkgBbrY+j9F4vrEkX4ZG4lGBI
3C3PYKp/wipcCIquG2hb+bNLfadvHlnwAuOdaiOUmHPmar8Vc84Zp0+HPwi1Kopllc37OvFTNJkc
AWmlgnU6rX5OoeHMtWBpmxsH5KWxvKx666uDZVBdM20FHDhdLngcydpDNWGXkp/2L+IE/lR42JxD
RnrrV9pMv9Wz6HRkvD7w+0DNUZ+0lgTcXyD4IyS8ilcyxaImD/Rh47YB5GLoVeuG3k07/RkWXMG7
R7F2V6BZS07MgZo1rwgjLwknAOt8in5e6/DI6h714hc+e2q6O4hWCMJAEboOTBiOewLtdOipi4zk
pv2XBCBlvY9PObeauDA+2oevi+/+ulwP61FB9+LnE8CHDjYLbP+hn4qEaeAxzYHDSkx5e/DlXCj1
DXVH3PkEkJ/xImyO+jT4rrPCBKIrm3m9GoAxduIN5/dQrcKR5hGtkiy9pk+ZIiF1635Uv1eaB9F5
dg1C1T/ASaO8TLVjnBhQoI2Bdd83pRgA73B3U3QMhizQcRiSdbETRfyreEOk3itKQBf4hDc+SdGZ
evzQgf7+poLKEDzkDwglZJxn5xmZVcMMBQcVVbEb2mcFMs3m1vOWohL7acq22H/kfOyrysKHJhIt
We9Bxon6OHlX7Jv6aIyNv5baBdIA+AXv90W0chDc+HFIcvBos2t4ebPH42LpyhcZaVuYBkwpdrgG
k6K05KdAucWJJ08byEyXpT9iMaGFHwchUmcIM4nafTa3aWpm/zsdizowPWUQzxeeDz/KM9e2Ly8R
lDPZEIOnCtqpLqa07+ZrxKqP3Ucfiu2qRi91XqMi3N+C5bluNTVKEzo82KLvbxCku7BKLa+Vx0Q0
MPFg48EMvAezOmet8qPUPCureLbKVHEHx4nCkdKTKmZRsZmEBR9wm/c00o0obRsZAfFIMqclWTc0
9qxOgnw2t1/DvI5KG+eZ9/N5RJyJjbqyP5ZH8B9hauVkARNhxYgXXiPg9fMFNL68ktDa/nHHT3mP
tovczBknmlAf3UUsvEKZCnPcKWU598CB9Tb5LJz8t/MTw6MkF7zot4qYrvf16tND6QErhGJBBRr0
H9JTGTnFMGg+do5xSRRe2mysKzkcNfH8KkK1VDh6tda0PnvtNrc9z+wbhvRGx2bmSruoGgogTeWy
RWB2WYXpTJd0K4s/+LfXiHBw9km7MshS1siEk9iWsEsuyj+nYOaTnlY//5nv/nOwk0tIxl+IpI03
S9SsrtZTB+ZJcZciIgDyCw5ngzgktnrg+b3/ENAGnrHI0jTYkLqjMr25iCBEOCImXOuZFLB0P/Rw
IPDJUc9zprV6NKzB27kDEs1b1kxZbk8h10nvhGSnNVvqXPk6p8tLbK/Xc1wEyGq/lzFVE0d8Sskc
ggUUro+cNaJ92Z17QS/DAQ6NcOKhh/dw/EuE6lHD1XQHUFw1JvMaa6y9UU1o6/9G1E0QC5a+bTwO
28KsdATiEFFeXhPAY1BdVeAM5svCZGbKtKulRKUpjtwn/xP1lFP+ZR0iY/41pElhbNi+9oVDUWKk
DFmDFO4PeyQClqIDjjfdqo30PDeFyAsTBIW1+h+avGb0zWVquu8qP8IIJJeGd8uLoQbz8Y+cVNQm
B6Vrob9skYdiJiAmtzrAzNKUCrY/OsKKbH0FcveLSGYasZiEwPKvvXTlZnvAJRjiVCE10XR8MR10
KOaHF51eYQDYfXGWS6wdZmHapo/o992Wf+16ausnnBcBGewVZp5AYAwE8x2GCPYchhJeF8gW1vyO
vHmG2aLewptnSGoDDmtV/zHpi3/wkGp8XczHtCgVs/Q5jsEQ5dRM8oJY4OlALfOVnIPJXG0LTOfd
UG3/FHH6zjknIaUbyoxBwal7Y/cSmZcDJXhGJD3ZqD6lD0DGgTl9cs9vMHxHqulsFnEoxmjv8LIA
F4bJnRerpcbjk53C4nHfl2jj+4yXJhnCu2ESKvpB2Lnec2WYxrxbm9Zrj869Km9PzxhJ4EE/t69J
RTjcUZE/zCv1Pi+GDA7fPSjftEJMd1x2YCDf3MNFyaCO+5JQ0TihPttL2flWMCCiftVPhxJYPLhR
QX1nRK4yaKEzWW1yzztafbUX0ANAS9H7qI/NHa+Rp1wdpDwXobZkcdQwMK70/T5ayrM9tgNlaRuS
PEzkBV5wTo/n1wgRFAK3MuSffXFy6HS5kB9TLzm56w0B78YB7Qcf/JD+na3PmcCdf+Vhxi7Bdwg0
oJTJ3k+i4h5mGAT3r8bgffmmtB1u3sXCeyK0OZYTGtyCCKkOEvYFUoH8987hLEo98Eyx83sEuoGz
QXay7Rea2TKilv5mYxK2sqhlrje6LwH4GGihI8KUvmOduTLfjxsAVwY1nBNOgFKWRt0S1Bbklwdz
6ccMIXLIb1ybzr48KmYrgdqZUjlnjihflQTIMw9Oqdnr25KWZUJiaE5/xeaJ+pALbPDDP/WqyWml
gLswvTDKQerXOVNiVrjWW8N/77Ex4gzwCoq8+DceS25DppIBkP5UpfQSz5suoVB72EDuGG7tDMjX
RtUypcghbig9vZjcslzUISVeuSahoruIhFoEYdhTQAQn21yxwI2SdLtwJn+HRC/guWjJ60w0vXHx
tOGFFucobtBja23vu+ajT+R/EjAK6noBlrt016l/mNMYlcYwA7m6q6oxbXXP/P6sFSXweJ070Opy
bQvNKrVGKmDBQZrL5jNV3qZ1xqemOeGTXq5jwQ6FK8CFIUzU1GClm+VNiYr+u8CBIQ+WWmD1ZFRH
EAH/k8L53IQZ2MA/c0exHquQd7jufQn1lgQr0lWt6Mu7WU8cwD9VZpppesP5g7KNeG306yg6xSuz
T4+DZzGdcvcVLFSiv7fhErll+qK5Rp40dl6NGoEg7E9R3/a8IwjUgMMzZd+yRfpivbwnjhoHbhX0
TMrgUtJW4GYL22pWDWfXU+me0xIF535aiTGV1VhQDjJvjbv2yjk7p0wX4EtDp6GJt/5L8yFnJgPR
eTXT7xux0Lx4QhI51Wnoajl2pNlRiaE+tdhEb9gGFFBlXXS6bGwcZhhh42GfId5+8ZuduHEb1JYQ
zhTgDORao7JNsDKQl7sr4R9ZBOmeP9M1pk+SH/v9ZJ9kJpGNK6Xl7VYJG447JzD7d4njSEOFJwyU
miEor75VkPC33cu/s3SPaAMzCamAX5qciZQ7jVASjaRwdFsxg7vTkQDF3L0yJ7+m8rEfGmmT7MCp
yLFj9BvyIOUNWP2HSZJXpSTiSzA04dEZY5tGnmVqnHkLcoWYQrgB9XpU8G3V3ENDbloWTLk8yQ4C
/5Dauu1diT6UOyMFjBU7XA/zi4yWzg6FXkaSUyqBlV6x8ewPkpAMHzYCg/Q1OtjsruqfGKSZ9GEg
8bBPu2+WrL8t1obL6rjvbvCs5SMTwndFQDxK5OY1zN3UuJMQoJWgaopgdj6CPpn9drJ/4Mr+EQX4
7/mHkSa2wm3yFM+flK8ziKKjYUJXQTuyNpAFuc863nAVIXy+S+KZ/9+VDKeSQ3a0wz2dM24HxYJe
9vSGz5DErhtg//zbfrc9HgNz7zXzS/QUIL03mP04MWTK1dBVqc/VofXsT/C00/9WFgHJblVxV6zF
UVE4J5sbPX/mc27ukg8mFRNvOGkcpgHzYKE/syfpPF/5SM2V2uiKyMDKa+OVpqWdi8f2TVINKuMD
JTOQO0zjLZSgrPusQec7HROfeso2p+u/Z9+pvvkBZPDx+OHAAg7oybeSa+5RGoAqhGzXutCpBbIt
G5Y/huStwm7x8WIv/FmyOKVCcOJ+EvOkWQY6IAPqxFlMLaYwyC9mtmCRTOcbPNolwFw1KEoLYOSA
GP+cuwVL5AKFszCAhyDH3LPXEsd7mlz8NCXCq0cDYxlxnaMJ/hq3egaCkTI1LY8iAfHjzFxdEWUz
1FJXlvkD0iFlG0kgEqIpCrh8fntkM6AO24bEJcmdwtTMj5NjM7iiO6UVyx4GUhu6hcb1GTXHdhIO
1AJa3N180HO/MCNw3IsuBxcrEBP88Zs0HTn8/zGnDdbxTYLxCxUpIXxvMeJ3f9qIgecnYtpXgedl
0aM42mswG9egcS+8vjTN45DLeYFbtACSYK3738Iyih4P+c3Yh6Avu/+/yIrzEjUo7XSqFx7gnSvK
mzW77ys5Fsnv5nsfiB7x6GgoEwh/EvO3CLqgYvMVOvvIQChrtm3ebAn6FWATd6K9gFooiaitFunJ
y8h+NwWgV/B5V6G2Da5lhaVzCHXy9dQTMHcDVGZPaS8i569fyzqcSROSsFyHZbZrrM12IrOc+Pt9
HsW0JB2vaU0x9+ckY1cJuxED+lNjEPiYfhDSvLqZbpo9YrzKcsx2V0G1R8IkUYIls4R07ZVK/YkW
7lWKPNxpLv0YLjDfGrPNfF4gDQMIfBa9KROrbNJf8tsaFunUAUoWBPnqk66zcMSvJmvJhnGMAH4R
egSTzX2xVpYG0nME4El+qA7B/OKqZxB83BzDClKfXSdZxs5HYEVY72L9XdqqoH2gCDffvBx6q9oZ
2loij9R0d/YDI6LjQZezHzMWhXZrO0YioxbWvWqOGtXzW1BFLG2znSnreeqo2sozvttSI/cKJaJA
u6pZ+B9MMlr2MI4+gCVISg46kPbHVuc0lDSGRe9X93fSVf29KRAWviT2dZemVm2TVcP8wMiKAfCI
/86KABRGTfbibW7fG18nwPpLjUoMFyr5C1n91X/fpoZNWX+E9v6F//SSBZMJtgvI4m5JEn7/y1ns
q6AcFAjfcG5nOs35mKkOYAtgHxM/Idl8nnVm6y1ShHslsTSiQs4VQBEzNQkIqgTD8GCHoPI+c27C
APNIJaQRcxkORiAL13OfvHWO3FNj5ciNimHZFXLWmILzpz8ugUTYbmnufoi147F6FcyVhCOj6i99
DEnWwL8wSzO/kLfZ2pzwyc8xNLdU5IgZfeYZtOB8iuIsJlu4XkFnSj4yVhFUzdVbO8E7V5DRt2vz
fmUNc4J4pkWbVQBKQdRJepr2U5qYYj5pYRqJ+la/hiEhXffMDWK8r7TCLLHlDvpb6OcTTmDeOlUq
z3UxWDAyX+UwXRUW23g7rTyNsuVwOinEvp1bGyANwtEVn4Lb7RUiKA64vuOLfxNyYgW2wp30EvDp
fqryrunrilMVPn3Rietx5WF96oxtYZXrwk6ziRGnFOTlwqZhlw/GMW1kZWvSvZb0LnM1qCJtuC/1
DneBikjznGp+qgzf8/yp3KgZvF7WumECod+ylIhyYljvHQPO+XrcraD8YqHlk4FEMhCJXwZQmiEz
HuzxchUBp9lQnv+J245mA3+1hWuVDBs7lv8kkbXLVfMo6vBzI8LqARvqMWdjqNxiy6mKujIf5xI1
zrzb2oX9bpEjVLtNvlV0Qt21Rz9qFYjsNx/Ixhicd1qi3FPPt9H29MtFqVsmtxwC+CI0Q8A3e1I0
ZrcpkMoO3zHZs6rdWuNLliNGtOghboQtcKcfLloFEXW/g6Z6QOk6C7T3471ytownpI7sYDzIgw0K
5ZJw5JWmIH8VT4e4UhgWx5hUFG9KBSWSz/Uct/LLBR1p14nMDjjoaOHsUOk7Y+hMbyOLYlOPjaHA
QolMd2j2RiAAonY1S5lNpvzTF4YjOFyKzEsZideW/+Jvq2V+nMfiAbKCc+kvw96/Yvo9xiAGjp4e
Kicgao4xga/5MhH6gbZN0/M9um6DxCVfX1jA7f0YVqH0esAOAgxTzz3qCQsTxDlSBAXVKHmn3rBs
TIEXUgA+zsOChWEUMHGGAgoMt8OG+26vAw1LwFRQnX17mJ6SQe68xsZeld+AKUY2OsHAbdpyyaJm
yCSpCv3QXG7dSJFpXRlACFaT6KI2jIPe6Gr1IHeCAUZ6s8tp1fYMG8NoX8P2EvQ6uchrJEfCpYOn
KQWo3OxkJvdvaHorrVKlmiCm13nYAJwahxTTkg02e+2JeslGPkQqpQml8+/uDpKdVOYXhAfWKSUx
8v1i51p61bQ5zn5Hi6jJ80JoQNGiHWtSgTFxzyIg8kCQWN6ZnrAxw5fOJQZcSJ2CDPYw6inAzcn6
Mznc2ko0OfW9plT/W+gsax10ZHpt1rPn3KzPRVqqvViGgvaXsPAXwOyK+JuAMkkYcH/GWQ9/4ncz
2VXPMKO7ExUunNRSD+87g2hVnVbYqfKIFtRrgRO287CbtiEznlFgm0seLzeQHzQaIaus91kn0C95
XNNXvl5kDehUCMkI8EZoRXAIoZSNNIdYFr41nMSqygE1WkonlBJtc0I8Mki41kv8WiL9SmrZKtWj
KyTCgwOAe4SdD0Esjn+lXjdTf+0MXaLcNXZUOR0sPEmok02/5ITHrVtU7rnAcTLyVZuJHw1KcQpQ
cqaEQaLzdYAVg45/mHsjk2XOtxyxmCTaefxeWO80rUpzRyy66H3GPAD0KGZ9BoAyLFEEZ4w+FVtz
3z8esEawaewz2GwN0YLSNRcLvDa4dou8neg1PwERTgAIsQ5fQJ7mXBTTVCzwaBsSQgTS9VZQMuWa
Zx6m29RRdKKueMJO//FMnn8zhy/LRWpx5DmgzlnW+V8HjacRG+W4iosJd5+SYcKrUAJeNy1QI7x9
0+ic2l8Oe0UxYcWqPfNTVkkBGYNjyluBS/MraQ1U6znRAnksPDJJEEBgWcF9W7LdF7nnNXYxs97F
qsaEbKjK75Q8ry8bYM0wdxaSRVMxiElLiI7ySUCxTNJL785Hf1G16MwMIt2hkVbHBf1bZuTK6rs6
qIALrbmN0aNiTOE7B/OIXsLj1qFdRU6aCJGOOQ0ZXqNqX5KQzgxfdcP/Ene5zjqHrYDGbfLztb92
VXFO5RHwkhfm/CYTfTJHxus2deb2jzLVy1uATzDxtW9S5tgNGA+NNSuAut3mpaTM/1q+DV3M9pl8
TS7bltNsZ8+FGzZiHQOo8Km8RB2NN43glatKkZXMQ3smS+YSFAiHkKQxMLMfHvm5+59fL7KW2DIF
TURwyQhG9oxaQaWEWgd+dYwvLCZjFLF8R/dRWTs5CsGPYVQSzJUEa7q41vhqhHf1m/2Y73vqjo+b
vt7ciOfJ7unKbNg1Iihjb0svxMaCgpM8sa63HwnxFUERL4wlgyEVygGI0uDt7vdiujz3+/KgpS1x
tqL3NQe4s7gHtzDckpyYVzLtizA5FN4OTbipSCC4SrWSEa/phbC1SegtkzJYwhbdSuYQQN8igsoC
CpZXtTG0dKvWnt0k/fKcut8agZ4b6N6GYaEpH3UFfyi/WuqThHwK1X8m9qDN95g3zfTb79LMz/iz
YZzmXvAIsSebVJE6YI4vacS6A7SvR34I6MCcdQOT7xbpfJcfpSHyaSFLbvMkcFeL/DvZVE15qTQR
NsxXf3RLT1lqsn90lWMXVcuyLq3aKQsgtGQfSGNt0r7WPFl8qVxruTgmNVhWvoYprTTlVaHD+ATL
nMAygOQFEd8bVZaIfelU4+cHobdozp0MEpCneZ5HfElr7LtP8dF6kELU36UjpEt1i3k2tDs29XJR
wd/ylgj6ypUdk1T/BUgkoR9Og6Z5hTY6VqkWxPnK+ESkDyBDzYQ+ZImCHv6p90ZvveJ8oDO2XaOP
naDpY3KLUdSylqObaQZggh3zjgZnKowrgb5d4GxAMPyanRxLgSSMNp+9ucW3jnsJ1FQlLOkWL6qr
wtZSB6ZgQJICQJqBZJoRHWCZgVlHnmCnkb5OwP/vFR2SMGzHWlP7mgUghu69pPtfbqWdHb2kqfGc
hLlhUnsWYcXus+gw5gdEePPTKIh/DIiO93eg7TrIe0z43WYKK2X9HcbJs7f2A8b3NCta5yTRUjkD
uliP+iN1rfPT2gSGl9yrvAdK7OYsqDgMq9FCXejd1g6lNvmgAXT76OIwJuOqLP9aGAxUoXF7K3q8
D0jquyvf9VPjZA63Ivd4AaT+s9iNlrGySprQptpuI6iZKrH7Wj5ebKmYVai7T0Rnsr9+15CUaOH2
2SnZhlrJniiTEQeDLJx6TJrtjTwWMZaguYnyxgw+4Ex/T6z23n+Sx8g3O+qXU4drOBXNCPenn525
f+ZnjZ4Yu+ULGg2JPm7YFrgWMYXxaUd1MHxR8mrQ8YRy9SwzRQwtN/fxwGXL9JzD/YayUYh9FLlG
lLwDD7BsRpOQxFqNdbk4iJfRIHnfsg6KYJIcWilbJqApmIjSXkXLFoUa1r7KJvxw4E+FU5BA7kpm
HxD/Pia1EPc5Jz7xFF0IuYBBC3QeBM1WfVSfsbfyefSkcApIA8Uo1nvdWK1ip0FqwUN9khZvD28j
DhztJGTkIKdbuQ9+mpKKw/XctNriUYd5tub3kZb4rQjll0QNjStnhim9hh057Naohb/KRUc2m6pI
ulc3DB+ZtQ8imgiLetaJn5Q9jnciRKsXNRFsIIOg5Y6akyDxik1UBLP6CYmkdoyHWvwuoB5mvlfz
koaMKqmmkKDiC0qlZ4br3DDQNYdpPOZZJbjQGQviHo2Qz8+sipznkJVSYLmszy9OB6phkjTbNqcH
mgVjCPCESLBhLyFfI57K2Fivcv0DujjqqFul0d9iJTkRIXYnA7rEnYt/toELpsYTR3ZCecY0c6uE
+9PTLu9wP3iuuUjavtEzp2EQO8o6TN7XTGzqYnFBLC0y94HDSTvuDxBbN0KvxMvOPmfci8iIjuo1
Kk+on/U2+gA2OwHjZbICTA8/7gZqviPrkhuPE4SNWClDxP/3Ua69AN8du3Zyea0LoCiLI9Vt79U0
ovr/AQLqpISckdKsG9PcFJzPLk0TRycrGUd9ucXEGxldze9mjsM2FNyO+gKWWfI0JL/eNOcdH+AT
Y6+tjDqjI7ZWPJ9sbWYiugWVagB70IgyKSp4qLyn+SNbdd2kW3Zjtfy2GteSevIkTUVVVjv5CS2d
zdNT5z8X8SKQcOzlxCm1u3/mURsGxv5BAx4BtfsASm+4VAbNHgMMujdBTTmyjAgyDEKBE/6oylXh
sghwaFUkcErHoILGZYMFLPBoMSt5MSHde7y6Qv5cjmxzMGIeUzXD5m2YAhOBi7zsJU7soKyIXtbb
GcTquWSz3XpU+k4V9fjEsJ/HJGVcIXSyC5XD97fhGNjBAe9dw/8I1Oo0iYkz0Ls14CnVgAWQXcJU
g2pXQwaVLTWuh8j7/GtC4cDmhait8q7P6Vo7BQatypUHXrDc73wRqDYBXOfKPVex3xJuoHjSn/p+
aVTS7ME+fdRpK/rhI5fz/TLAnoikZt1gbQwXr7nvNMZh+FyiglPLytc4fPYKNSqUWeebUQdNRuma
fBW91DH0HLN2W3FSr4aFYtJ8pmOrpWQfBhuUKwIkntT5QgV8hw1/XJRBflYfy95XBTBivzykOIwN
Fn0k9e3Nl3M5QfA0Y9fWzmCdsM5t/iRwe+oQMtX2l1o/sjrA1XCU3DvPJK0+aw1oIXaRYWbhYhra
sNrwS1INHLy6UJA8OKcu7mNg7zDWNijoWxVxJAbylA8Pd1Ns+7kN/XodLY3TuLwIY/tl9YUl1i1w
raIOtSP/OMgTl720vBIXauRZjXKVnDVt+DdQ/nyMlVHk6evxz3PYBI2mcBc/Rw+KDWhWNJwIg0Wl
iNFEO8JEnXnL+nkOOlKtH0byEGPkeQYvXyO6nyYjrlnGqiYrFQBdjEPzDriFUz7BxvCIgn3KejBW
aNSZtldcwRCvvDNxJof+MIhurtgnrsjoQDxSeqszu79Vuu6tFIh8lGZdDmxSq586/uflqrepSdSw
vBWlEnDb326nleTprL53NY4P4SsaAGqPetmlfwzSEm+JBI7SAAKSPeGx6y917E55rToG1H9LNzOv
tBelnFXrZjLYeotqMWBTYOCcaotqW5386uns9b/4I3o2nr5gIp5rlqZMr0+xzHKtp1o+z5coEi/C
5lUhuKC7C/Gs1B1l1L0QxyGz4vlYs+ch/E6aIoewrCsFfxqohHNcXUL2fQS1CqaQ/kzkwBxp6esj
mqEPI0hKeNqhA4/pkmnHvJmN5EToxidAUSbp1ZzW5wddSlB0Zht+MGbSyGLwNoyoOX+9jrbpi9nw
7fABoEtuHrjYndkWBk0p70e6Lv9u3T1HhkuWVn1E+G1zxsdgkdXc7Bf6Q6snaG1MNrQ3+BEIedzE
G3GvH0qW2NHJh20D/mizRbnwO2eoqyxh3YZB3Npcuoz7y2x6Tt6DTqAi/dRh06KcBm6VqDshkYde
X0Sd1nF8B7ieDkrBkcTkLgLQUnlAYWOn5x8FaWfq0DsmUZ+fuCy3QBgSsPBJPCZkmu3BFwA13UVa
yYF3JB6Oo0MlKr71EYn38ql5h8sWY+h6dA6N+HhxSirVLTzMMXFtORXCxT0nXFSCCOw3z6+UVPNW
FUqsbngvL3jDea5cfhHRJBDsJ5QBzrurLrBdvx3pA4gMHuyNRZM3HQlzk3ZSaSVN87flq3MpbMjr
j8rIcqDo2xVkcuytsjnrycDPOiQLu1tVOlaTIOncrTLNCrMMsE9CnkyRxgWYB2WQvM8NBNBeF23L
XFljSNxqgowKFPwVXehSx3Bw79YIat6epROWpW942rdmVFNXdkjsfFI0YN2xcio4d8hbb6X5q5iP
9jKocJefM47Hmlo3AFyOHHqaJeqHzkr1hnJY+RVEf1DTQBwor+b2WwHiT9EBWZ6HymA5+cN8HHmx
qGdv5r+Y4Rz8JwHdR7Z0WWxOcFEkIw8cPpO5YjahmOZfpDxclXdAhxX+EOaLewK9wOYs3Sey2zR6
9sSOze1/4SvBmNMZKK3MgrVScf162/I7Jh91E+4EQAXPz7SRswOKjAQtnKlP20rLYD06YRKYjaOW
7xHtN5z7ZLPpFeU1doRDos26+TRi2x1itcI5gT4FmFRPub4/iMCN2F75dGfl393gxNulVB4J2Gjt
bi0QpvkRXpBmKMgPHi8SLffRWQuBgDhF3Au+PRoBvQtJEP62bf+n/GPvt7gfksSnkzYujgDH2CO/
ObqWvlJWtCmBS+eNTNWVN7cwMSvLlHFt309dgw+mFTZa0dheT+bWZRTFSVAzylt6oiDLLDGXSCpL
IRdEkwcvo7kxEaFp98be3QOwNo/pM8E2/m6J5Owa+s+x1G90rVVSMub3tPcTFPqNuwjUal2Rx/ok
1fJkyrKRaOIxP/8Ic6Y5mJWmipt75mzEPmC7vafVly6OH5XIbpFDjxhKfJElZ+kVn6cqXyY98Kgf
2yP9cIXA5oIVbUTfE5SGQlGsLQ7ylOdT3fGB4up6k/Vicn0x3jlvu27tLGPDO8qgXDHyqf491BIB
RmawKxyZy4StVIptpqHiTqGljn6jnoVnd9DlCfrxEYFa1PYEN4KCKm/H6xFjbTbqfczl4mjaQazZ
9VyK9JLIbW6CBznYSQ0LRmswd6H0AwWWTUU8WCphFs44YDla0EGQ7HJewQU/chRaJOV5Jv+t92np
BM1gC1M+4ZYJ2ZO/06OwYZEFnapfZR6C4Ibe2DLP6zUiJm7BXjW6i38YxNWM3QY8665H6zLIJXyr
8vit2uiITTPTT59n5RRGIF0fA+N9BRdDrNiOU5+1oNz10RPLHDJtBWGsVZjn7Bh8uG3brRCd/war
Wf9jm/90MH/aBYxqeObpWOtTyL7a6hjvEHGqCPfEDZmClK/TeWWUp5KNKIhLzgDgzT07Ojp9fT7a
6Lig0HV49fOMVOiyZh9AHBQONIYRDFfMk8XDZ6A6ddV0sf5nGlihzmCVbr4AlcijMmratSrLBWLm
IBUvUU15OFb1/8Jf0Sjqvhx6PKoeJ077+84BmZ9xiCKk63LMofW7ktFGaIxUoAKxA9TUiqex05aa
fUov1zfBQ/DhXjSaXw1tCfftmU5EEkS++ehxVBthn5WlabuhjBoJKcqEIYV/DtlGE0EyeG6J5l4g
y3Y0NKc97hRgjFVZ/Ld7vTU8PNxsPSkQAbpaFyk3fv54/68KccmqNYCe6fjgYLYCg2nr4/HjG1bn
2OriUUcD4GbxIhT8YPzl0S6r5/yJi9aE53/zPT3w3gkyae4LGLf0zJktBFrl6mFRNy4W/9PJ0Tp9
g6ave9Vrd2d0kD309QaO8aeY/HQmNtA3YmZ1vqhlpFJLxJeNw451Q190ybX/S7r7YB36rfajWEyN
TRoHpImuHLaOL7sUFT235zg7catHU40q+Mkd0PCenZPa7wdG/wEJoGGO93hOOIpEfBWnajPnJ6uB
5x5eTBY0twThugqZm3F4OYSmM7uIoA7uFEYkQMpwSLPW9/IJgFwo2rw2A+6MYT8ZQNKDRr3JU4Up
Alh5JfQdp54OWNu3v3tZj9NitmrHcBGJh0T/1EHr07pP9MGVd89UNOVk0NCRwTSpOeCcFL4Tn/Nd
Slh5MlYX60i+0LCzUfhhzOm/dTKe9qJ6Tfv/ZPeWgZRK4WOv7OkrxLABdEavkuyv+MMgQWSZdnxU
kXRJg22NDjCE8FoIs75FIsr5/5IYUHEfgn88WtBZKtOvY66ZgIbi11S315yO3QYNLekA+kEZZHPv
Y0poakzYCYIOKhd9KiaEdRf3Be+L3MqVY1IpJIir/A38k+xCsgl54Sdhli1YsN8o80BbPra6fYFa
fCDv2h3oet/PouN7g8IyrOemdZqyIJy5yCNjBG8BDAfTFSrrZAFVEXHofqheBpFMnm6SpvEAHv2t
yPg4WIlBU3omQsrd/zwDhBA+brHbIxQ8X5HpZyx/9I4dSJQwMXv42gveKOUH+5c+hG13II5f2EeM
jJBMvnlWVLbqC6PEuDZWuwQfammujsRP1MXv63Urs6liNXbcJD5eh3o+1szEKXjV8H3388qM16mQ
twm/Ei4z2y7tAMbh1X3NfauMHV/ScXMYv+9+aktF9GwLyPH4VE7HLm/s/qwz9/KeUN6a4nWE26K2
ze/6VjwmH4FMuwl9PCWLngVJTbPQ6+YeJSPJw+U5HwFJrJU3Jlo+a59WGwvxTrBsEHkx7DqytZfJ
arG2bE/1v0grtYMMQwfSV8YujIL52JvByZ0+RM2OJVCkls8WQwteuUEPIpHRHa9dI//UACmPtXxj
tVuLeYKwQq3X80jnmXs0sUpZtFn5HZIljMzHD9E0eAKkWCt0p41wX/TESFBQOSAHhC3ml9WvYFuV
VAHdz2GUXn+z3+zvWoF+byawMurKlbP/dy4SWKmDkv3OcXP3csgywzUK2IAN2UIWfi0rWUrC66D1
8OU5Qh8L1yo73nns0EbjahprB4S5fMxTPVtva/gy+EolYvJJT/TTEq5E/Cc7z+JQel3ffIlOIBqe
JwPUAy4RnZ0gHKas9fu9pBc2rQIwLAuia2+XF18LDf5FoIxh+25HhNEHW5XmmicUomg0bC3iOJZz
lJMuhjmBEaX+cOPotarf94d0pGcJZr5304ytz454A4URoTL0Jp0wuMn0sA8FGVfu9wXW+MlcghOf
m/2PV0xCWeL51fkDyKTaB21lYhwiF7UENN/CdxBaflrgBX27hFpSn7FNibDNhvs/s7F5gWOnKzcN
Tw40qZAa6g7iMxFBgEWxX03khVAkGAKOU110nW3SVXok71m9orevyZvwUTPsk76UElsMafeqOquG
PhxChevr+hNdnGF5BJZPSFSLH+oNM922wIgCEzLLkUEMpl8cS9v/g+hsHfBc1iNnts67+nAhfDmE
sLmv5JpQfqzPWhQmLJFHXGclmDCumZBjFflMh4j1e98MxJME4LRjBTzpQpZw6QRqKmNthdEZfh7e
gYuli4gaW0V1cN4+lWVQEaly56io+S2C478A2UmlXDZwk1pS1wLjrgcHBuaKRNtjU5ZEmmPz3u26
BBqE2UDmFmurSEEVXTk3W5iiS/iPYNjBUHfhTWlJ9MH9UFuNnHTH3abKLcRvy6SYX1P2ffy51UlH
r5Letd/GfsjPM1HiZ6KBiRuTXLkTOvBtNnZ3XtyzjDZAjgxNr0xq4GpbW+QnNxol1hEhsWayBmeT
6lg18ajUhftGHeSkcGtq3hE/JR+jXtoOcENxC3c9B/uOUKkjTUZjGcW5Op85kNCyMmYj5CXf9sOJ
VeiKpE4Ty4RvipI5HMGjQ0h8hWwFx1h6jD9m94w9rFCMnFbl6ODxvN+QMnVSMPKsvpsBGL/TELZO
EiV1Kenw2Nlo3v8ayZo7hLQU/3br7K5aZVQpwtpNUbO7n5aUeIqdb4hh6VYEdl8GWnyRnDFABAIC
BXhTbY5YoLxas4IPk/5wryi8UooIWQuem/xZVuzrMbfHMZehIio+gdsYwKQGnJEDNV/Up/DRYhyR
Uz2gytIafEbEfiv6x1An3BG8BqJY6pj7KMoAFnAXnQdnEJtqg5/CJunx4cRXPoWAHWwFE7BaLwhI
ZTGxleJF5w2VMNlrXvsxCbx21A2/AxyhN2d9N8Lfu2+EaQ1PwqiyEz6hbq5XAn4bsiu7y7d9Pa7L
ewukpUdmL65NIwuKIM9HEn5F9ooy7s1vC1dS4HF/n3Ryg9CRXUsB1mh8icu0Vlo1xNRqm1UMkmEH
AAH6Wo2gSI/gIgmIaY2mXLYp6wRIMO+em5qdoTh+96BYfl+kAuGWGifhkRuGNEqDv0jYBjwjAg8u
mLIaxaMO+CA5xlQv3bbyZ0P02+HPZZ8J+JgqpTVWrK1KDaPJVYFSrBGEf6hmVlkn35PkF+IZCskf
UMq34q4By+fELcVUprSDQ/5m3NuOCl8H0Kw0Dd9UVPd/5jeQSRVlI4FTlf6GRpWGnrZYJ2iIk8gz
IkFBYcgkHI4hmbh2LmuJydpccR3ZtqsntdF1VzeWKQ5XUlYEnAceTDBO+JU+ggF6vlTkHdnfDgsj
hHHR29FOem+cDU2K1xeJI3K+KpSymqueuBXbj5OCZAMsIsMNumXVktTfsUAZat6+Demt3uowzTQI
QIRNc3rMv24sBfFVUeBmC3ntAzraTi6CmY8VNUkeDXlBwejeclJTrXvPpOiQyCa47DrrD2stp+1I
DHjBk9RQE6RJM2ypva6pfn8O6FEIODwcA/E6vjQQZNnJHx5QTjsdcXj3zOaUDG/CAgHdf8utsVS7
MEENbyqzZ33Mc9+JcRS9AjVtBX2O+2W4Lbrp/pQvgBjFrkVot1lPLyS1PmjKT16Fwu3T5atFAtVr
LLX26LOohEQIrSNszfZr18lso1DSpyMcf8mYbyeURJ8nVK/lJlalsF78pSpX5OpxKycvWxX6w3r9
b57Jt70P7gSPhU1zBuCaOr7G4XJ/8ThyjKnKn0OhXVYGq5GEkqUFOp+PNl4/HlmZugVFpGmlZXAI
BzeriQpoBNEovstpZevhCDBVmsl5RRDnGrANIwke3D1uf9Uj2HO9yHEkmc3jQRN7YS9LzQ9hZOOL
73er5lSW5TRM5EWlNV16N571Xi9BUrnm50qJX7Z8IMwOFe8OdBqpCA8s1Ft1sw9zPFXfedbGpWT4
wBsJPYMhEd8KP4LIdRbNmi6+ZxPRfB+RFHDM5ttFLZGoiUdiZ46fXJOCxgUCpmJh2iJGP6DZMQ7U
pY4lZCtNHz150CCJaGIDfnz/Ao6UOPGEY3Fe+rsxjAydinT8Z9IInmD2lMG6sjjHUloY5UuyygwC
MAF1eIT4yo0QpO2A3rja4yRghSjqrIQ0ua9S6OhRrZ8pIwPOSj+zu/djv2ihXZUDDaKhLdML/5io
DRcfgpSMYA6HoxNMwrYwOgXGfLsjhwdxGEdJ5qkXtMHRvrDnDCuQlyqU4R+1PH5LftFqJvgJMpa4
A1oB68HPg4jEpctGBa9wCab6jlRBS3ljBBAXd7zpAoB2AuzDFMF3MCP10j+F2FwKHEDRlYfhkch3
zNmgitmT+IVFpBw0fkDqa2GYxqW7COaRj91xXfbT+XoE+oL644FgxvvXSDAeu5ZpDinG8WO2jj14
QV5GS7Awtd+SupI/3qMOUEb/rLF3ohRdnNsEKzlORYoJH6X4XHYQhgpv5Nxiu+9WDsl40FH+fAcX
nKiaaWjAkaxCx6eDoEo7fZi3KH/442hNUpmyoEqXomkH7lKoc5UfAx0fGVdKPB2aG9Hxf2ik9nVh
TEv3cBO671kka8mJKEPstXwXg9mE23LFv41zWAsIpHq+aj4Stw9jsH+Cy5CJoJ/FYyo78yHCYF1q
BLfZl6Se7n40sXlTmXcHEq/pljf2CxaW4AfGEIzE8y3+b9KNMN+6xYBKfWivCklufHtZwkHrcypX
CH4iMMm2N6IXivmeeoliseogJnhBhi36Pr2bCOkCHwucljkoZ3klbrcRNmUfGmSJOSWkWve9kspX
ZQ5Qw2yIL5xkBYZA1eJSIHHKbFOKTzPoHr/BOqyHujghzmAVgcr142Fr+CsJ24TPb5rmmKHdmBPo
kM5WbkUYdKQFaBjcP/ZmlizG1VUqkOPnn/4Z0x1uc5g49ojLcCYJFXuiezydnky+VWMOQi+hWQVS
z6UVf3WYXYvOQMW1rRZg3l2fcOHmtvShs0+arpq9vqXPgzfLIn8borOUuLzAQdvRoLjo3k3/Drmg
X3C3tvUrojbDJV0X3pDrkwFVrF4nSOp7lT3A7bb4RnLcOen3CzRro8Jut9aFZILMDb8lW69gJbj5
iNRqGmtF5tKDdjh9QAl6nAgKq3SlJHxgbb23qR7/9QtsRVeGSEqukVWoUBoPrKLl3LX12nDMWIuy
gPaDWAnAJMLS6dERoP429vyusXOlqkG3TAg7buuHgzlKntG4aPxkQf98T+vFcvHAFRSvh4LRMprc
Tnn0pSoM8r3UWE2psR7X5ies0hn8Y45xZpLYqLrME6nvYLfrDC/E/qyjc4YR2XBsFkaNfzgp/QNW
darwUY553D0ko7avcw/ZcNakqvLghqUlSaISTUTDrZAlLsDa1wyHIRT2JixRzUkida9ARHv4QWr7
QwBDQGX6yLTkkxkUzTO8S23Y4uUv+jAFIVil1sbtRvr0XumjkPZXq0c+f2zZoaGLFbKitqRQ6O87
ZwIyDJS999V8LvN1Ep94LKt5eLzC4hxsHywG9J0IauiBk0Li8nnnSR8hTtYUXEOLnn9fxpgaHdSp
ZAFsReb2bU/b0nQSnJPiGZ8SUR9xJEHdRnpuum4nPrukqzqGYw+aNX40yIFBx0KtwZe4fW2HXv8H
MKBqGX0pbJIUF8kPy6I8AORVGaVF9tv86BdZ/S2DPOh+rTJAuhLazyvXdmpsphUXzYcgANWVsTZx
D7ic9HDePnVqmRVvom8bpwM9+HBNA8OSx00H8+QONRWAn9HRUAs27/ixX/Qpz0JA4vAAf+boEOqg
lOHJU+rvWrKc54CKm85Z+piPAp6gcXYmSCUCm99zNrhbOyH2Aw9QGsNuqbpHnZAXapS+OvptWNPW
+tBj0hdHl5spRbHd5PLO37Cv/XSbbKkFancIEsZC8e4PwRjtFYk5zcyuS0nZpFdgq1lDi0tEEXBx
yzBZm5b2laEwek3ubNnIDUj97CKqyS+tlo2zdKsgxalCotcdU8GPydHatzH/SeuiC9F4DmQmqJft
U+NjCJxWAZg2L7odBjQ2zFZHkj111njf1fZjoOzzvOEetJaJX3TTTy+H2bBJ5qfY1isrn2TyZfmw
QCNeRANCrv7W34g8p4gmSpcnuavbvPHjSpEzo8JDqS95MCpsjLJ+dls3KrD572hkOG/6CXJzjv0f
LXjB6rRt1yybvmeeOZihJI/KhYGfJ8PykOnLdcjpkSpCuOzflUSwpKJDK6tTEVA0mZSzwcBpFlcQ
QdI5K4fTd/AHuyNhJeKsRkckgE4sG2w5JTa9ATQXLLR6vxbOz2nz8mu3by0+Wx6Z6bD9p2d7n0Xl
qHxrD0BnCR+jkBfpaSGZc4gikBsqeIFn49gu2tNuaKNnZgG21cO1ZDGPMu/b7mhwX0I6mUeGDhBM
9CFVKURN87LNzYIfGgNB6wY/rp0oea3QQV3JSVFAHobD4sg2VU7QPvhDzOPU9keRNT9Q4idbG/9S
45nGhGz8yWcdDZW9XK1vt1L6gnqCVz12RiAEEYl9TrKvMFRh5H8QvAgC8prCJHhpHc1tMLhDoP4D
xG56E82qqKNqngGRAj3UfAnWVuOpKqW3XZTZMO/3GAar70EYdp27uuBdAlG4ELQYkN+Qae0hPOZX
D3o6QCuJLqhaKQQYbRf9F5dm2lgO4kndmwRMSNZ0uAATGmFHqKmhW6u07OtzNAI2iMjtJRVwXSaU
HwlGhFGbyhMBy8Xh8OjBRKoEp5UrdmJL7I6PcH3lIsoxpjI523yi66cOujTcvgJnr+0Oz70/Ywrj
cgY5t5HcSg3JTPqpii3+uyiyvqQYM+jfwUrL4+fpBLdnAxduj5STe5w8sbWHcoPZwZOcCf+rpGaH
fCFAx3FOqhtWWRsoF4FMcbrMEoCUoOiQPb5AhTJU/U1S5PYtTPCiWAR31j9Vr/gtOwC1TMNejkwX
8y5n0yxszfwsuPqm7r93l32loIFjJWuH1FKp+7kTpatNFJ3poTHbb2fMsKfx6qg8DrRs7x/9uyDm
QM/zuNxxP6wBNB5O7ekCabEOYO0ZPcw1Riurl+MwE+J8DtORyL5Kp7FP59A3Jy19oPq02WBhdflK
vBIgaXbbJ2ILGyJly3ZQEsszmCg2J0ov208yI5TWerYYE5YrzS8UHoNsw/OKd8cw2VuVmCaDBrMS
TsoUzvdx16K6UkE5ugnKEDM788VSg3bHNC7cv/n+/e9VSeH6W7BS4Pnf8RQuGM0a+/azHTWjX0Js
wSIRKz+a/LRjodMgQAjDsvGpIYVhC11KsdnPvDBv6kLFoKcdfnZMklTtluM1Kr4gOaFTpgNx9/lg
bi8cqPhSfJmnJIGzS5Q3t2sQnrwZlxB1rl60px8bsYYdqCi1dycceaEkS6XLmNDgfO1kYeaqW6C5
IL8Mil/sh9Jbl8BmOBCvj0gN6GsCnySaWXNC29H++ispE0KFXdpfBRUiH2CrdKSYvgz7mZofdWuL
X0G0we5RSZhHLtmEWzu8Mm1YBpMGKLajHRwFbjjqXq4e/EMQDxvPKrbfHZkE9dm4y5uH8ODbAxki
9a2IRAzb/T7DZiVuV0KR+nTw7ugaz57GcMwFdxgk5Ag6kkFtruzAr5W4azlp9/PXlNRXjmKmmq7T
awYT56bfr2R5DRpXd8R8n+o3T26kXKUz3O2DeQcqOmKob4F266OJdrOynXV0+D81gi8zBn5vgMzP
V3MOsF+YIYUV04AE4cTuP62YBJnS0FxryCkGb76fhwufIcTlQTLKM/LntQTB/VfuDsysP8yztLm+
GT2ZNtD/Qo/jIO5uEUhfG75O/5QDl7aTL9sMyGF3Rn7ork3lh8pglGdTafWo4eC4CIQn6PgwS4nm
Veq0dWplSaglD5leTyPDlxJkJJfzl4clvMyOh1WEl4YAsusm/xQNvQHNj/R6P6/2v5IyI+XnnrTC
HE/lkTlLsEDHsAgYnzTuUqql5DP6TWG6wtD5g1GOSlIFGL1AJL8A5hx/iYdQrnSjH9VQY82mSiuQ
6sFzlOEtWFhoyEzPKVzL4PA+AMkfprkyoMN4p3W2v5eQtpd97hI4tDcuJxKz/pWs762JmMyLo4Gw
RKsh8HuKwequbrvhULgqLn+o2XEJB9VIxi+osgeVZqj/WtVNugUTDW8pSDcKnP/qPbHrroDsyoB5
xl8f90qxa99AQ9Dl8L6GBbkAwWa8BYTrbSodYuWTTxPqN+Qrtl+nH3K+xznrBUyZ1L8CjhVy9yL7
Axw7n0jHnGtWEn2cCI1BVCaerR/kRrXsaEDmJ93BQO6w4C8PdNYFwOiN/3FtOBp81TaG7Trqr7tL
ComkUA2hO8MviK81Oz+zERmRTToHIqJvy7wHFjhwRDZ9TOJD4Fv/ND74ajNr2EdpdIdWolMGnRSl
1ZpBg3yRvryfvRNSV4e/sJWncYaXx//eDc/Vex1cQBE6EslZnsmAlrOoraW2kgsBG4684qwVtoxc
xrfBt83diKgsg2Oqwr206DYXiJfK257sJluwsllwvZ5fO2W/Q7AUGqdg5BOATCvHv4tL5UeywmRF
SAGPn8lN5e00Pd3a2ys772FBNqkgfcrPtJtSV5iz2f7gsYjKSsHaO3aLt+D4AdCszYxAz5I2KLc5
QpMSHPeorVs/MwTN3QsM4qiM0JpH3rbRsWTIyFclE+FJb3iEn+u1Z0qOKKZRGtxeCnpKMreXF6Sv
UuIQwdloFy5qNgBDCLUq2ockv5RvyPzAEgnwAMFiay4QrJPzWqQUpwzl525L5awKYFB8W3FyyZAN
I1SQT1oTMOQzI2W43dInOuRyYYB17Jh3ZE9tX+nAnp6CB/98D0Ex1JjFX4iN07cicQp1s347MPyb
Ut0GyjRbaBte/Rez85vWqpAajhg0aj6Og30Yj70F9p0qklbA5rN6jdc1IIMD6RjL8gNGq8QmqF4z
g4JJnzl71Vyb+CsP7XaHwu6eyyysr13FIqzCzJO+Xu7FQPe5dtaDE9ACwLCSuckNdqsLQTK39fJx
eysBJvgdacfUnBU3NojdQs5MWc4VQSiqAY6JWZVDZdOdWcxbLnn7a5vFMXcxu7ukXe7OYsERjei8
Aee2ZtxY04yeSfZZl1cLl+KMaqllBFjypFYTnXTXsxvWIl8QlOu3LnM7yKui+r8kDgKDh0qn5808
/1pCOzwkBg/abPXiMDurnXVzcTsdLh+vVHUkgbzrSdBOmpfx9CyyqWcU5g/kMW6cXnQg0LZi4EWC
NTymt87g7JqwQ2VISbIQyxPMc6Asv5Tnx3kEkh7EcPmgWzM55U1WWVf7M10DsPAiIQV9630n6X2l
ZlA+cRZkd/RDdajThEIoWF8IHUrj07q18SvHmgGbTdvORZf6xQJTiofiBfALS/VWfKWmayCNkptO
toUj+eJSZYzjFOikTjY+n+N5ko8P72bfZQoSDGm8SopSss6/bkQVTqB2q7k9JQWHyQi4g+h0Y5yy
5Rml21MZQK3+J7EP62rKitOeqSl90z5mtcL6rQUNOlno1LCh7NHNNx8fe+kVh1WmwvVIEeUjrr1/
ULgsdxYutLQCse7JyvOrkfiESSHlBC5R6FZIHq2sKc7AzAODkvqDOwyY8MkgGsR7dMX25CL6gTC9
TMP67OTF6lCw5s/MYq1B8xth66DSCAZvKXYPUNzAB1pb7AQrrld47/MRchJaHNNSELxFpBMel/En
nHrFJUszhyvIejhyvUiYcHorh1BbLCikG7PGQwhnaoNIdsKRoaZMCR5Jj1925st9Tyww827sHmGl
Zu0LKon1y4+AmvczGn9gYux2Oywmsnhv0IdlxO2+q5ZwrUAGGVAuUrdCShwmhOyAwUm5QdGkqQdo
jaKF/sBNxPUOlv1HunVV1HI9nWYIVDhdVy3dMVWrvHPrj6jxg/wXgnR791jXpSrK2fm7PaHIMKk3
Rt4knpJfTo1Uz9GSm/Q4wrC1E/f78aillJ8/e65NSc+aXpU4PVISeynTstfGwMXglT2Q5czTRmu/
U9c+Y13teF9NqhhH2SJdOMZznUBEwGY6PYON3Jjfw38FAFrnaxetAEaslT+XL4JrkG2CyZ3Dk0O/
cen4+ll9y/8UAHx9W3JenZ+igmgGQv6tSHXHUc5GevSX9o2fBFtLNomTHu26TtwfyhJrgwZEIT5/
eRjq4SmPkf+hFUDmj3L9MrHbrWB8xgp7Vt8FSkBlOZgEeqED2dJjAvpOLbLe9lThtGKtX3Rfhuxz
zm4drZTOrjORSQZN92p7A9d6EkYrUSIrU6wuNS/T2U5zTiHOp/wcq/fRR4/doxY97rWeanjwQSA+
6acLISJHAd6cRnOYVZKHprY24SyTTsYr/rDDnFBIkrP2EbjluQUMgaIYy/F4SVRURFSkzAi6fn0t
+iLw9qID4jFTY9QLhua2W+YuUSAgEePrMrkuvLzBqYWAA37ovCuOIqWQwat2rTWQES7iwfkW88R8
AmPELoi1ZKiUZ9/hosTl3iGdjH6dHVtbW9a6kNItMnNFinPbx0RdoIiVEx/OF5O7+kobOiIScQ6t
fJFR0QYGTMMYns0APJwEcZJkXzpQa15S7ajbzgEnfMk0oH90lmECDJuArouh2qIC173cwLf/gRII
V+NB5yEd1MckdZcUmr3S0okJxp0VCbFoWFEsY/k5C59zDYy/b/YLlcAyMx9nFGvHHtPMPQYziRrh
hycRH8ttnTKajBp04TBef47Z+W8vHBjpv2ITHq8NMT+Z2vXjSkGNCfLqTZJqeVt+nIJ+fZRW0HKh
aWqDNeysU3H39rKNg93i2Ilqz1QZHa/ClFhtTcMkQm9fctvSM4zY6xcxWA/FWTealSvWV4o6eBmj
4TdVqZ547K/euADNyK+qu4sBkLI16QkamvZa7xnFWerzA+K+HwaN2NBCpk74YvTwqB/1v8XBrVfW
fbMS4Fv7F6GWHF94kZqMxLqcJe1vvKX/UtcpgA58yJ1AVFZtPJi3OdNZKlAcdswpP4oB6XlvK7JW
JgCXtZ6cpOAd5HJYCn+qVg4ctf2O4qreQ6Fh9XByTzPWYZzPgmS3qVfj42oNfxGVhJEv+iunFl3m
vSUhikkUN+A0aN9moM57v1x4V9f9vhnE8QLphatthSz4sfXp6BKxoA02iEvss0zA7CaWMrbbzpCE
1RtY+t3O6BSjhKZOM4c0lSWmc76thjdF/CN8MrqU+0VcceIkf3DGgoRuMXg/qZvbuoROzypPT3hQ
34VOCy/eEveM+ySWXcN3AvFmp9y8oDaspHH9vjC0IXBvy+yjaBdwjtvgMYepiSimL4UEJ1qV8i5j
5/GPDH89FSydVyqfpfkVsLdvtgXE34TZtkx2Ob8NGVkYPQGk5PI75wZrzbeye9MTAJYBQ4HSumkl
MEln+GYb6+q3DNZxnndGkxQCcLm/tf3cRdYx97Cbzx5D07hMCtpi0CqNECcBnAL03mQ9FL6KLeiv
Nbn37BihFQmGR5UB8cEsy0CIziBSDEK/fsE7m+aY+c6qm0App11Ijh032pNhCZWuVgE3qcQLNxvx
PwBurBXhgkFoZnvYyHt7hyN2PWrdXkxPD22QK+dqHG6ficaWK8Ich6dpBmpInNEfAOkgJcGakHOU
8ZPsZHX5JbiL3gZTM9AA0dMj5dGjja5lW+e3wem3wmIaBOwkOvVfooL3KBYYJXuCi8CSYdp6oIi8
13apFZB6uu7gG9TVNH7s8wjUBNYRINtY+BnWcpbaBm2X+JGBXcklUOOEw3XlKD0TwqKOZ55WxMnq
J0xi0sX7XbJX8vUiRgVMyD4o57ilCzNl0YlmLK7MfYrppB6DhaGfhnXz9Uz2veR0ZJzlNvxmdiCw
bRAOywA3dK4/Wk6KYobHOlaBcOzErUdJLNsOrQoDQcg/Lo540VPboS0mPLEWhoQvwpqQzNHGeeYm
xwYAb8I4B53lBr5GuUlxxKsl1vxG7bhcyxUWs3dy0SMqLm3D43aY9XgiYb3cmlGNUsep54WO6lYP
SQ/XRqAmWkBu0czdK07kq0JkWTvokRQtgKyIwRhwyQubikoRC0YqQ+asAEFpVclOueuFnV1uzqav
cVFucYCUguZnt/lqToFvkz6v/ieBf/GebDShM1jMlOH8TQhkBTUsYcFVqU8287seDHMONLBOh2Bw
OnUh/7/An6VYovA/bZ3F/OvQ0Fxj17OHWgnCgb6gYGgwqc0ND8AruR0mIqM4u3QHcPjP5ltiXDCz
W82i8Jg8f7EnT0I2elCb5LJmMzpCtjbsBiadlAdllhD41RBb/EbEYG8nIQZWTvZ59VkhIm7mbQsS
HmXgkJwmaHBHRmnYVkEgjd0MPOjseUTQENCXYo3ziNs9ybylkhOb1k6IUAUxFDotIOnZC/t9QZXM
8ufKDvVE+KAPTkYl9230F26j3m7hlceBgqMn0ckl/V/zX9a2QDZ8yN7EOYop4rZmeY4krXdeM16j
5blpicW+Dc/tfx6KazU4LAGKNwPbe21CS0DA4pUy8gsR2qwyk1pSPQORg4AdkzODFEl4RMdh/x3t
5DxSvtkjyyXVVxFekTeFpuJLpmfIt1E5ZaQgSXYDRfc19ibJR/3awjWu5G4XzlZcQQ4oAvlm8BlR
nHM07e6ahUHsULSxYFw5DMjY2RVLyeBMYLDsTDviJ976Ulg6TxlgHa7msYzmjHCwqrh9LYXy7LTE
7pnpwGz1B3a9JKitxk/sOPPCgcZR04JMQ1nEVUcAfUc26K9d57Al+vD81k70CdcKKPtFu4tHsgw3
8WZXOIsSiD6BTTkDoW4SZOm+nC4gLaGeMun/CJEkugq/YbYXTzvy2r6+srwXbTo9R4rCQidDY4mp
k2U1dcGWGUGbjzv5e30vr3OtRNKbhqORTjOlt9WZUCZx1j8Mgxw6BnDisPytbkbzd9ImGnSGDVh+
Ag0vw1oHaiwa1fYk/UlfCklcMmQd/DdNMi71nTSyKcm411oAvpsAEnUzS0vwgKJYzIoN1HOUBMsN
hwty/FxY40CFKTtjSDJe1xJmXPUCcWsoIC10sTpl2wyhLESEb7LquEMc8t5+YJpy28avYpoKr0Hg
SGknobqiev6LhUvRf9BTfe8czg+ZkjgEHsSSyAU7ZesxDEcTdEO4ImsHnGUWTnThLCDGp0FptlSC
09dfW/CTBCX+aPRityKuXWXCj0VolwjnoEiIBUyiaX6NWyaUpAIDU1EYmAkPzSJEV++aAqBYepkg
CcZRYwwEAFDoo4GR2uXk+uhrv8DgTnyu1m11UUfbe2jC5pAQ4vhn+SoGvdGVa8zbPJ3fkw8IAFd7
SnTKEGdzi7TOxd06f3S8aUxMGxpiwILsSN+JFB4iz29epj0xd0hmQdDguJJQNkMubEtbWSeOS1dy
AygPbFkquULoosPX1ANiS308qPBTjJjeac2QpNywQWsNd7wjxt7hrw8ypY0mTi9VYdfGxUDnapPc
YsjpwSbv4u9FAO+IRQEPjJI9FShnGP+kzNR8X7XKtJ/Wf6UelNQ5jTzNfFqOvTUfURRv2moaXHic
5d2WJiparc38Hmu3ulaWxbCcnPKDj0OhgtyLWEZ2zoDnwrAeSmV0yROhU3U2gBkjTVdSvrdw764Q
p+p0lVllH17/4FNQ4VwDiUEy2tW5L0LDsTVtVgY3xBmiX3RTptRLAo+mensGruxEiV0iQTZBTW3g
LNpv9ZE96mnfBDQMMsN2FWYuFO6K8A68QxbAc2StsMyIyQWivqw8/2tFzvrHLr1ZKqAnXjOu3Akp
J9AdLlRHC3Eso1F1vsG3snGVH7/Nficdb+OVBDrgdQEXTOIZ6Fc2SiLBnVmx3PsyfunevxsRfGI0
neFnvAxAQyh5So2eEyii1RL+72rcdqSCWm1Ym0t89vIbslbN1BUX6QAXu0cbZ0cM0lD4xHMpomuk
n5G9KwmKRAPZ24Kge3n1HY/gtpgopI3uXW9F1zJEh6Z6pSxawNh8s2InXKxPGJQ5vGKbjQzb+dg4
bgGoX0IAHTf7VtRtfISHIv5SaHhieYUaQYj5ZAX5FTbuNVkbyK7n75suBH3m3gq+0oaLsRKpmSF/
yliQR7r5xpFoECPDh19Hr/J+Xj6JjdlLMLKiTJIh3N4Pqzj3/UrLbaaS+vgbnjTVvCc5EOSr5FU2
snTX9cNtmJUeC6BuGYOEg3u/VDT0RKGhf9QOVufd87WVt82HDFsmt+rXW/9Y4KvS6WfTHbdV+OcD
Ejq+wyMpYwh/p6H6Hph17GdKysCedbwC5LpPzN+68rEg5Q06UlWnHrCyX5xiTbi0a+5vmXtsWqp0
VOjMU88GK3bsW/fhStJi3/aMcJ8sdAcnoLZUZwul405WUa931Qpm1fIoYKBJtZb4FYz1FFiyZQFc
DwEAe0AplM3JV0se3WgEQcEuF/Q+T6gtztp277ZrcHjboaEolf+CWDRSjW3vbWWql0SK2ImPu8BZ
TNddwmCfOYRUhTLVuxyR8b7lktnoCIGqBfaLp80Fjun0cFxBvhX6VCsiBqp90EO2D+WCtHAcbw21
FK+PzmaHDJGzFZrM0AwQqMzkEbiXo7TpJ/o/tBjG3wYNmz+JTTzbqUhLPhA8BI1CY3/U+GmXogdg
zfm+gK9nDo/INFUKSDWjFhKHrLM/zB2KyMxNisWzaO7lVHmwKe9VY+MeEET/JspJPhAa4vmHaloM
Xup9zGdlPn9rAtSslznf4r6gyJ8HiEYA5NYZ5CmjoBW1eHzT98BjaPZn93RpGu4lLyjzttGBoI3k
uhRAXi7Zav544AI70gRKEuOucwJzNdIl6M1Q/27+E9a85jtoeq7kM9y1ZyhHZH8ShRBnaP2pBrWJ
LKpwTCkyOS6oVp3tSuEYdjQcgzDgzbPEo3XTBR1iFw73ZQe8GMRvpEykdb362pgk0v0syo8/1gio
fw8R1MZzBNBhvLoStPusPWHO6qMv2ZlWLhdUix+BQN9tk1OK1AzsPVkYopJ2bSQKw4Iiemi7vNaX
g/pxBm18cn/HeYSeID9egDA+ImO5fXpzekAy2q6FAjGmdoIoYfPuTGZ89eUQ+MN1dqEQ8o9milI7
ODE0AI2722+sRfZHGhMOf1zVBE09Bb7pLxF94xaCY4OYuZyaVygKYvoGwDckJU3OaXXW+oEbAuf5
v1KisatUZ0UNkxv42hv8KdPkfkiHZD+zWkdum9vGiBMjB9/nzFQTK9R7gumPzNYmqa1l+vgfGfGP
8SeCOWUqViHSApS+0CXBQEfdfLkulcFnUjxFy8snrIrN37rdJkQLWrOmjJICGKbfwv8EJqj+XlbD
1tWj5b/3DRqm4KlSoc7qo8AU0p/dyzyktsm6RCEgmuPw059r/JxaQoTm99+DfjtI8+dWulwJEIZu
LbykMjIYwS1eUOdv9swRMNqGMtSxBc1mvPgpVvqZsZmrQbl2tLkVaGkjp0oCQhbyjJP33z7A02T/
LxTgdaNyzsxw3VtuvFSb00187y1T9GUu/sRFWBrULG6Buewcp5Rf7ozTqxmfBlzlVqxQPP9IU8hr
LKgD9iqQouQREKgB3GCYrJkjXMBvLEL7Y2RpH45owM91+RB46A0g1JXV826mTFk+sUmesNDJnvnZ
hjt6bcBMXoU03fdq9Pd51tzbT25ZJlW2v0ZgwvAz7NCLrG4F45xmfE0pVJ1oLqC4EO4tgT4ncTHt
2wXXPGqSBl0T5PFbdTIcgnkEJ1Q0OHrKQpVUI81yAUOJ7xMPRoM2DAJCL+5+PsdoQLkwUZ8ytOey
xRQZarbXIa0qRlGlIaCk+zCdFdsvdp45hzXt2iY0nD4hBNfVYwPtuQVNdqnm4gEl7ZqCzVkTwq3y
02Wi2g5XXFL4lD5jy+4WQDBfmJAFekfG8djA4cWSGakNw4Jb186Yj7VI4lpymK9bZa2ZtLCN9fNk
EjdeDdkTqylA/Xx2kTI2O98wmNh7bGhPiUV7wPqrTR5+JAZrncgHu+MZO2RFjLVY956JV49Nyydu
6A9R22adn+ui1guraJjxk+FzpUq8jt6zkQ+yvXSn4hiWzN70ATypIpyl+05Qypb81FSMQ3goAXZ/
WTjkks4wfkquJcO4RrIud7ZE/0cSQ9BAxZdW4RLt98in7yOmvhr69D3la4IcsrQ8IBuedV8xyKN6
SD9Cxkr7DJxicRWLonEq3gJnrmJ7UIBDFQZ2xfGk2Lqhq1e1pAfXBwwVYGi9YJnspBsS1vKyFHOj
qd3p/levC4Ibw5DCihIUD7sWetpj/EdrIJDInU7pt4V1q5XmLFXFX4NkubuYBu7PJVG8i3S0tAjl
5H3kON+AvFO1OrX9qHnnnR3onxoALdQ5XNrCn5yPDX+Zu3BVGNr/Ltx4SDZjzmKZFRuNo30Xp4hq
dFDuyzktI6Q82FeigmEbvrFX4ooSNA4cdQ+shHafBsCiRoR5xoNozS5EHgNIdd2Dl236HpTwfeEH
K+555dsha6mgI2DsVk7uD9Gk082/+woceepS/FTj/sm5PGEIv1fzuFYrBsiae5KC5lqId3gC24mU
Hif8RQVocYe6396srmvwBXfoGb2cnrH3oZbqtKdgSkxbPqbmooB22l7n5YJBLxk4h+ZiBjCVucYF
A35Xz09Qk0qZObbUUGcdILBgqLwjdr/MQQrNgh8klcazuKkyxjFzznT33LQD/M5I+98xdemWJ2Ud
n329cfFYlaZJzuHj7vFZ9xqaUgospsGjN/oOTMbmbP7iN0ttjFkZgjaEyC9kMSa62mfN1EKqGhIC
gMWcLQJvyijVyA/H16uuq2+Gp2TxhlHNhqTTxTiR/TNXHRVaEGxY5STuyKFiCNqzi7So37gLmrcC
DHOBKEZLiUi1aAIyGWLTTw87u1g8bxBR5gNMT3jUGkFJEk0gwgvdpF+q8wf9PC69SrnY4zxjVZMI
QcbTauUneJH7K+1yMmCOInqWeDHTZnxvg23iDc06k6g5Fd8HhWdVyYl5jNFS5DAW24zEeqAPwXxp
JtUzhJFjKWC59IXcvp/IhXatiEZ5KyVr9dIJCX7L2HIGPtDNncoUh/v5Vvl4RjDZuBwtGpWzWDPI
iVDRyOysGDpNO8fHolTaW6EwIBYOm/nVSXj/rRIwLcSSnudfHtJwklzttYCu+/a9jErr3YPgbdBg
9yM/Mbg3+u4gN8hCrj7cP2grqW4oE4u/4coElVietFCoSF7Xu7nsAo2kjjsSaCLCwRCns1tnbkss
Ayp95L07ixhxoXboGrL20nOCvUsXLSkrM6JCjrCQKoMHJte7PZGClBz+RgZliMtZ2U90htZhXlfJ
lufvPpW9FwN2otZCmBHJcywAAqNkOTqe7OG0cazQEH3tpZdvEtoRbWl9Sh5q26dBqvE35EViDr+f
xtZ1fYdRoIG/aqixoXoK9haMn8uj1tC9k9XAWuib6G1Y00f5oligHQt/T1yfTOeYpkFf5YPDzTD+
AvcESlDP4Zqr9ATzEJN1Y85Rwo3oNTDELqUn/glW45jfQAr1ZzbghCCHn4q2a/XC1nNaR3Xflu0G
d6XN6ErPMWjUn1ulDS0h9cv/LRNKdePbmn/FlAFmbXA4j+Wir1gGYGy5owd7yFswuimz/Umweya0
CckozXMLFK+xl6IJ7ytlX/eXUur6iefZwm2gjfieb8OSgdeTwq5dUHKtRIDV5yQbw0sbWvaCnaxp
Lpqyi7OTO0Rw4tNY3dJmlefTddAeJ43s0JN9fRVZlA3lw3P/BYzZwb/U9J37yG6b38MofMhYD2/g
TOVh7CwHUlgHSQBU/fLJQmqof3XrjxWeGzz+HeQds/0mpTKuNc00EtPhXj+KTlMGHmazOdYW/GvP
Prlgl0l+xv8cpeWqwbhrngidz8i7fQiVvYpuThL+lQh+9qP14y2xCsrPdvsASngrgT/1C+ZFlGbA
BqK+HQ+8pBkFSf+TwVyhhGY7HhGLktooU1XF3PuF76GzEiujLRg98Kt8EAGr1EsdfByhGtBOGxQP
yzyuUINJ7MIig3ZFK29Wkj3ql+7XiihnQpe6mgi41F4pH2YKlDrPOyf1iLAdta6ADKflfq9gokOG
FTE2BRYgul2VS9WykJZA3m5FPXpm49iy7eda2pE1acocWTilR16b5Rs3OVT4ph4V+2FzMFd+Vn6p
uFB0l/MwdoCqRbUsdrJ7Y/f5wriNF7ZTN/qTOZCOrUbJe4jOP+CQpw5gdIueGE31J1hIUy1bv9P+
TLSVH/s7s3iJMAWMKPo6bTxJHYEIivqgVsw6ayHByHgISz9SpRUpvPlB5Xgn6RTEvat2YvTpTzU4
N155A6LCHZAsALV3d3Le4uovM2YzaetoGghZnMgOocbgGWFfPGqtI9p+cRZjMoQrRDCKAAfHbkhL
/x6sETI51EhJ6forHUo1x7ob68lt7YrWpibBMwY1jqO3A7oEar1lS6RgL0LWeeoSNeokCs35PjQe
G0SxqnIGeQUBGFOp7WaQeti9jGvo5AeVWUR/uVtRvnofF8u9fyMlk93+bqDZ4lUJWGY1pzmtOUoR
cmz9hMusUbbdzXur46MXNcGv5hGKm7Z4AQ7xFZIufIT4/FNS/I9LBh12CrTwpxaqv598HWTPId+l
edhgFSp5cF4ZU9jNICnlUIhOl9CuX+b/OJrzT6icMe1B8QOW7OtbQ6Vgxy6w7a6QccXhKDy8/GzB
hbqQ09eIvQKVJeeauQ1uHuBXySPcFfvuB3SRzdsKTOzZs7pywI6d5bS5QN/Vps4toniTey1FDawB
dgnqlGn4KYGuoGYvEuWMJXfSxdPGlFpsuMClharIZJR28+eoOuO0A9bX6/5qcUXxT5gbvthOK44k
4xQoHcie9TCh7gaELwkweETgIyl11PlU0RBwpXD/WJ/7IP9ZggEcE7FNdxyofaUOZsomB+MApT3n
f3mF+9661kH7rpk5TluaflS4D/UkuS8DsB5bsUj1ZAyE0LP6l80s1thCVYE2m/0rG6+f8viDvnn6
UCUE9uYH5h6GIxc233O+XJZinwj53Bsz/HVpWZPRt4ApYkIno97Xv95cGUofiItW1lAONpoqtEE9
IaJNbZNL97AFuQ8p6cvFzoC4bD9AkIRkhSzT/r/n5I+fvB/YiR/5h6wjtCf1AaGWRSxiKoWkjKaK
DA62BYd9R+UYZHrSbOpg0z3Oedvlxp0RpbJmFXc256wAqrk4+ekSZUA8JNgVqppO3u8V3PoQ36qW
nGCKNpP6FzvXvtCf/hupHlpNl0Ib4LSwzzbMQbPgacCWoW4t7lHMPR0gqs3IAd3mpJyhFI/wc12G
+x3K5nGcxd67+F5p9mVnJuiOZPP0EbPVmgKQloZd8OjDSON9fxR7roMkpHqr25inh0Sy0LEF9Ol2
kXyCROyLJHbem/RYur1XkrT+OU07NycWs89T78q3DXlrQZxB138pvSTHDRj8xX0ne+VGJ3ZR0ndW
rt0gK19bqBKcYatyrswdH8Oo3S2lCNs+B8MelFY12IMFdTOT0ejniPYfuRHAyt3/as9hBc+PvWV8
pMFH+3e9JR53kae4StUn3yRoNx7NIfha4DSXd21XM/q+q/zgXSjvJJLef0/wNzcvxHk6+OJ4EFIS
8u3thdquXAL9tRV9E6/V2k0tiwyzqt1F0ziYKCv9wxbmfDHMU0gpMWUq7Wipp3FhusApW/+tj3LS
tNYD/agYaRZVzNfFv0FGLJMAMHIGBrd86qCutF1J+9Ojzwj8PTfdsJ4H+ZTu/mPEJR3BLRHrOVre
F5C9TITr+fqQ77RkuBBJkwTwud6ptPzPQxcT5fspOnBqKtdTJ6fOuyrrD/0m4963YJC9ZdIWGQlL
4PHrp/AKT9leRdDF+PgmmNXqhjFok7tJadhkgpq1cDUpLKcx/SYKBsWncnM8YmZG4gzmiMpIqXtA
z8WyqoMcFXCRAXORYzJGIvtePEe+4em+iA4G74hGaDZgZgDlDBXxkp5daNRV7IPVYjywILXUkmNv
ZJ3vi9QHKdivf2SN9VyMg3pJ6YfOxpvnGK0lp/qYgfqAEsGev/7gsYruf3ZxwqR5zety0X1M74kc
W11kwPtxRU7aU0EAIgYmzqzUWBKrsyr6+PBtNzkmRmY9DlCxKozF2lkPm4Lf8fX/HUVe/FAT4gYP
tnpeOI9U8pSvQJyJhPB/jFEE1NiwNFmRVBxangJZa/iEZfFbqOeuN3JsOxM3RHr/3l+hFMHJv8ok
0jXb/34Q9jc8vQKUiur8hmzk7cZAiB+Y2ta6G6ZdD6JXcenhpYBX/HaI6WEkjkxt1TV1Brdo88Lz
ipDq7b7FDhGb9FT98eD+FxVr92rCp49IrJm6sx9/ArMKhL6MYJV56DcHES+xVulVYD/DkhHKaOQ/
UB5hLQrfkESgIYT6blhSPu1TzUchc6owUqnOWwap+sTF91p9tC2p3q0konBIfC8Lrm3hkiDlk3aq
Cy4w5QsPmEsTGMPkT91brKYMG3veQJAz8SZOR8zDiK87UDP+dBpNL5lYb0IFNspV881WMJqt5/t0
0ld4T11DmJ+vx3iXe++fF3xGX4DiGYClv9U+VyfCmNnM9/DdusKYXJQ8y49qSqkGL0D3kfwLw7XQ
Ca+HIS3MWD6fDRERcCfRL40D2CR7L3GurUv9fRoWv+SfWY7zmkcQ5jW+xTNRFV12M5rcI7A40d5u
G3d6945Hl2RQc7cQU1UwUVe0jhg+B8ws10myioxPmU/b9XxlHLwxgxDKei8WimlKD27Ts1aE5iHG
x/Mj5UcvLJWrtyY9dPwM8FTYJrImVCLHWotprA3P4/4ZpGsUV27XTa+r1ZOxaYwDH/XaMlj+YK//
Ny05nwprZWG2AXQz9vEdrCjkHMQpHO5S/0Y+9Q490lNx6j7JAtpvXatV+lMWQctticDHxklJ1on1
XDRfDGwPE8g+e1sCA5DGAqwTW4dQM6Fu34qF/aKy5V0l/1dR4TIBE7XG0PyoaWCCA86/U4RfR3oH
h1Wsaw/90YLEyIteGM1I20eOoiKo7GKowkKoIteTkI+rV1v9UOOR8oGbXzFd3KzF4pj6Y+x6fTAJ
pvPP40V4PslaVxxVSph5E92jq8+NxyP6i3ick8XOvl53fcU7GgHpddmPKXhCVm2OeNZVNhQcLpkd
Z3sYbGPU7sY+PCTn2SDdBwWe5OfnLJT5nQy4KEh+Ll3pA7QPMbdIyGNa4JRAtM1R9PPFN9L3YRXY
ALy6NnB3cQPCEdVG0x9BGvF1uHcUMTOMjZKXaPOb7OKdHihwyyeGYpIsGhMbQvrYrv0tknrUqTNx
Y4AWM8dhacTV+B95NpDVT9hHF8TCHbLvfbheiHx5WCLvUndvwDnNxKJgLgoJctnTanSB/P96l+LK
YakT56Loi/Kwt7J3pFYtYkCZgifMiggDUFVFUdN0xvCESLYmhsNlsWPwMxgZTaEKPjVmgScWrt/r
uH0moQHVUnCCLEAaVJGKj2hG7kYQ2YPY47orZOZki1U9PnSllpZWB3SLQA1deDnYnNrnT83lxrX8
xPr98146Kboz/NVJxV1ua/Bu39JoBIANVsEzpVCNdtNYRfeeTrdj1RbmmuzWrQnXkrzc18XSklMk
sGjJIwkQK5HPnxyF5H9PKySAGuyuW3Jt9TEcyalAVjswUz/pSmA8VtGGq96c9TXKJ2JGtLYvo3+y
T/MS0BahYI0w3zVOAWPis9ewD4vNeuBqd0Og1dJ3Y5+ryIkdYsWJ4SofF8KdEQ3Tchu4rL6gf4sT
h8i7Nxl4xD2Chzlc65pqp5P7CHOg3OyEKoPGWDUKiJ1EEAmnikVRoc+gHWH6InN6lk15Oh+YhUD0
qqvRmgM2hgBpDKQfWqVTKUUfN9npe7pjPKhZBJmxEqkJLWxAEeSWwEA0HMWUhjZhnnFuK04qPXhZ
2VT+L3gL+5FVFpoCIAWs2eNtwzzm1cc9KrIn+mLzZ3DF3qJ2NDEa9y61+O7kNSYTT/32HwBvSCt3
ZPjv50MCQNa5v4TyOFX9FuRFZ2of29cvTx1O7EX6hO8r5ygdLBECpjs/F23uoco9qJQDuxQO+EYW
X8v5ozsY1sKcKEg9175oj5UnDkPmzHGlcbEmTpS3tGXAg74sJ1PtDMg3q8VdFePvWlYhAf5cxqLJ
2MFvOcY9MgfWKoUV5GAQ2dfK+C5dnmccGFDQWcqpaDcC0KZUnKfLtixNob8ECvfaIOb7opNQnisD
rM3DqLiZ3zWU3A8Ffg+XlWEyZ5sfIG8OoYclvJVe0vGAgKmETi3ICj0CvuwOl6mZnpyCbQrAlUsR
bfnoon/pl+kJ+4vIk3LLsAJHkBXGKG1j8Tri3GNpckh5sX+Fucq0WGfsKPk8Cv4OawDDjJ9eF67N
JGn7jdMyMY1wOeW+gGH/zMbdlYGm9xN3JDxYPcsYVs01YF1y13mxhEddO/od8Le56bq90UmCmMnL
pmQ4HG1ikWO6ta6bP+GiZMZz3EQzGhIOJZ8s3NJ52fMCkDFFIRcFvH2OfQSfe+zpufQglhsiLDG4
n6Twl3rscR39oLd3BUUiORvH8NVgvUnelmieJdQ/M+Xs/2gycA5aD2ylje04poRFr5+VjQFVKwNG
R3DCxcNDmEYU0g4jVqrwr6IjBuDt6JG7B3oG0DvAS4+UPfPyboxlEtWfw3sVox+J4f9DWAJG9TlK
FNtVYp5NqxnSt/9BdnSr5oubBvTlTS9VIbDCM59dYcJ/7h7YOOUP016vD69ylAIOen9SiBZvJYyV
U1Dpu/YPy6imAaXim1Bw8orAnyJWcgEC1nceCJ97W3DTou/v3f7vs1BujUJTtG5lzkvDAXEVt6FJ
IWBew4wInezTidQKZcV4KA0tB7MRg3XnbM670KeNjlTsn5ENtMmP1FyMZlk5SEMNeZ15IF1+V6WA
7USgKAVbdbB23R/kmaI6qVyCG1OpgzBTMavzdKdxwGiwRnSv5yGBPu2yXdQ0sE3hmLnjVr4mbJQQ
9LBfPxH7OIra13w71r1FSwcXjh3xAF2Yf0OgvIIk5ZxJNJBtoGxnmb7b58ZE53+shSOZm7c4D1rY
GbxBDCZfcrS5uI/grLRcSPZjTpV13SkeZ03hNzmJYOhp3EAVd+KfWOJDXCzyAbtrAlMqdtXJzZng
gSw3SHTEiemuOBdHtPDpcoKxV5DGGvfWIMjUXB7dFMvux4tNR4KotuEScwJ9s+sdlyMUBQG2UUH9
2d+Dk/NjzhpL4fSzzyrC+DVOy2KEbJIYDWk2vONFD24J/LhZpmgdP7l+qRDkWXivMagvSrsxizcj
CP92jF4FnC1JzWExSNNRQDjmNsdpv8RGV8GZ5aYpEyprrgnYLc2u3UoMJ5nl2t4se1kqn4s9fNYf
cB2ICOX+KcMvuZ0KehMQc8t9V8i6RagFGtiFE3sgIhDa1dZhCr8uSfJia+l8w/lT9HWzj8mzCuEi
UJHbnAiYqLgzix9kt9/efFmxD2w1qMYUsk84ShhD8+tgEXM9+m5Umv5DTQrEjsdbHm3pRGNHOLP3
nfgC5HnSvcEVvJgpj8T0aVrWyTkRYqAWGnmLQ1vEaYLrUWGU81dKr6pxAZudFpbtLyYFUN6ZiHNO
RWORv2PbjgOygxbBovt19sAGlNM1a8H6rj+NSQoyznjTg1S/77WMHFqKo1+X0+MZUKiKYtHFMfaj
uyaE9icMJNJ9skOWltUjsFiBvrNT/y5JLy/3I7gJn7W/K3YlHydp1du/AVLJCiWh17dBYv/SYVuQ
3HlnZ7UEGCGdEkCD83c7eoxmYFC5/6HDmkiJEgJE7lfmwRPxdHgCo1hsCWaR0q5/88FhO9z4v6YK
e0hu99+yMbOStUuDvLHAV/FNiPcH8K9DXT/U+n+hld1D2zKajlEeMrEglcepzkEjs0Fxq70WQWnB
N8jRGjZUfUxOGZxYKMxkEntWOVMcdaM1f59YUJWzVe5kOGJZ0YOLMvucYSxmDHeL1iQ72wbIeJ2/
WO0HWfkWLMMz0ROKDxtvZ1Sie0IHSmB1ETTFt16yBXD0cu49BPmGEngZ/TcIOeQT4abtf+YJJVMm
k6nVhs9CP7crJmnSgJwpJy/pEeF0URz0ElGytuS+idc+ybN7gG3SbLpiWCpBdPQrSv1/FSZCFwit
lE3TdnNqnEzh+IAhNbWTmUilOzogkAyMdvrsws+e+IEcmArrBb4xK3eF7mhbBsmjZpwUemFw06wg
R8H8S4HwJ++vDCxgCxh68lXmd2OsP9wwA3LyC46kRFYDGglSRKHxq3VZmHgMl++CjcLMH6PMqpqq
HmCxT2Exb/onLDk9X3mshI8J2n0fDINvx2dzse3xZ3JCXqkf+st9UWM50MI3WJKQkRbJkfsuYvou
YxJ+Yn4AGsqnvFV33MeyPAgDk5u6qqiU78g4XUrxPHzVebl6wVghSZ72e/vGa/GsohDsLIF1xZUI
7+SpuNwnnUVHTSb1uJB2M6t/l993gv2pZpeiVk1S/CvTzRJdzplga4Pbz7/kZ6YvfHJ+qrvTEhyK
/W7UooeI1VImrVEnBRJoqmLJRSGgy4fane7tZzMjsppjMEn4RSMo8xION9VMV/Mcvl+BttTde7g3
cPjM/EInNE3BliHr5XI+o9ceNvlfsvEGP5eItYLklXqbVYh5GuHfAs7TCrssLo6PdnAX+j5ah0DK
lXQwPwmbiTFYd4NDm/8k+72s4ZPQoRDvem8wYGockAySfP70hECWZfWy5Jsrnn1MownQGKx5LLch
CCgvMcH11sCmk/5oJemMe2k3OPEM2jjcv7R0wk/9znR3NKQS7le5KcppvKZt5/zspFLFHkbU40nl
QxLYpO18cNHTZvDRWxDKeMSDwPUBUSeMIc6R35ZYXlCaTK8/ETjyvoPJE+FNIo3zKc/jAo6WIOR6
bZJf6KXO+5EZBSiQDxUxE3HBrucqvT0nhpMsNRi+5xEWKRFJfIHoNcORw0GEOo9VNg7RAiqQLnv8
VpL8S6rKaiE+wyvgd674s39/Vs/aWbSsnhQfG9WhY6PUneWJUOGMeYdHpu0xWO4L04LJ+54WXSks
uM+g0cFW43XIP/crTTwNNbL0GzARO0Zm11bx2J+8eJWFiZEHcTCjBZ6v7vX2GjOvccJkz9UOxw4h
3EX/VKP/ifKLSiqhpMu5dBGP3f4TiUPc+5NtKsX9dn+dry9SxrD5PAoffAj/Q+S5AF5ygGGl0Owc
heSKnP+nm3pkwfc2sYGyeIUGxTyCrjgcCdAR9dN5rS6UJPByySMshpSEn2nYUjMhL6ykwnrdoCUe
oyyNrcbwIKBpox4TmfGoTpB368BympLe2GmyxHIrhmeC9EF1m2FKnlQb+sMAJ8niMT9ylRLSNF4y
jtQ8vyopTNqPJelfXNMUuMi7y/hBsuYJoPdqcaY931glVSSp2OcOXupJKf1HFmy/KIDXUkgz/+Jb
m3E69ELmv5dzK/rHbZi3+JNlo6tF969djgF5zhd1eOmvzFwzhK/xqwkH1oBTw+fdmEadfqZdAJON
QfGbrzX8q2q+hD33FXtYjInIyTL5quwiRabPyaoBDe55m5HZaaiZeRExTv0TOWBRze6wTp8p74YD
D/68UzUlAtfsa1JnZXr6GdYIYfgSzZkKT/VfPBrTdb1vGO55+wQzUtAPmcqiDLRoXnfxRuHcOH1S
TwC4IqJyCNdle9m9enn7b0SlujVEu4FgQUdHi7pFVUjPdSST1OYT6gRYeDg7QtgDUBgZzbTORbtj
9nbdnWFsc2pCA+epn16N0ySrkcqw6qKDT/5OkmHxUX5J6+FsDdUJEggL5vtHHqIb1qISad2JP1zf
Pt5B+oowFD+uL7heAQ7aDQNDf/2G2eddWoisrZhejwuaREkw0BekMtb6MFsMOUdlolYg2GrldQBA
Y/kN3gryHnYX2tfh/cas9yF5e9i24Yl3OcZWaNatKQGZCWdQF7qh8ENGAVYvdlN1+EIpQGXytAZf
YM7iofOfftb0R+cmIsY3+87gBZBvUUcKbvZT/vmWh2h5V7K0JulNeyP57G2Rr4jyNgjJ9z/PF7MB
y6y6BEJwHOlaHNFHlQpcfQ5QX/Wm5LDsDhoVIj9hhltp8irHxBHMzB/xoGgm7mFIPcpFgUdNSKoP
I1LMHXXWJG2UfKiHEzuhdpguYP08da83nQTjtROg2QdFjHswCLpIaI0VxdG6bnrHbJDZNMQ7//p0
YHUuDCOMPc79WbQZ54qWX0/oCm8cV0qEx0kJ2Km8Ew9c+BSf9VB9rLQf8KMIPZo/hUlausT2rXtk
kdvfRfp6iZbihpUoPXnnM2nWHJvWLGjslMEE47Q6FnMjjFN5OqwhefXkDh1fz1BUNrU1e7HoxqmY
cwery4gODZDw0Mfejjbrv30Bt9J+rE+NHw47XkGTnvFpyaFV2VxQs8AJxmzk2/tURlxxgGL8Bx4p
+hNQpxdLK145o1Gvuu3F6bt4oyDvWixuVxCCWIHqsTl8puRpCn/T+LPq4YxNkyZw2LRUfeap0/Ag
L+W58qewSblH9Elu02y3Ex91r7MPO2TrEpjkbvZVb9fbYYOI+V44rG9rw3ygI8u67ND7YSPNLNYu
HNrLFOsO5Uw8ABeNFWlAXD3paLk4UxsEErSLDA3cAV0pWFpCfpyf41REYPqY/4uZri0nqjSll5Yo
+dfMTVLMsn7qFpye2IYHbjzCbBKrWhFiNmK1FrN+8QKV2EfZY3j6wEWjoRQoCPA1QoIPASRF6xpF
QGBGQ6mabuODZHjNl9VM2+EKHWAi9fZM7uoEk09QJe51qpN9GQ4AaZaPIX3/F7SXHiLaq9lSfkZp
tS6fEgY+3MDza8ZbsmY+RIrvkRPq+aXGz9iewjiDgZ8MKb58JKlcWPe3VcbuQB1OSnyC0TchYS/z
jJGMFGU7+cBWPPDrJJ/t4hsMYKtjQcm+PIkI5h3eIEa4LsaLhBERbB9GYCw4mPXh8+8CUVIt9ezc
QJfPk0mFqqLWlOWUbJlaadiL5CV2aGk6if3BBrZh3eoWrkRb2TG2orcrEwOSwi0zIWNS5Rt1TESW
s4EBYlE5Ymt8wV0P0k68dKE2mgN9wRwqh6Gw3BAYb6cf70U7PjmcaDyyolZ5uePmicDrK1iZv2xy
UHK4uBP7nRhYYBitQejibMBfoQCpIkX+vsGG00ht2Pec2qZ3+EnwD17exMAzn/nM5tBtHOcDwGwD
/uL1Rddl0Of+UuS0rzdmyoS66SKYNYuYxr5P74FdGEsb/xQbOjonHwSYYxx3h7hP0gyCw09IyAjW
mIJ0BR6lBwmKHHgBJaiJXQb3NZTlhirBYc8EkjNSVioVyubsc8O3aUTqkJ7WAFqMP1/L5Y+rqC74
au+5CLDRJuHhv+9VEG5keu37OI/iJ2VbVizz/TOMBLUTvfvLppR5NoMrlZv6za6hFv3VSNZIcI+T
mY5pUvJx4r+QqvE+47KsqtcQC0pHg7zb+jolZZcrrTRCjN7zd+BWkcBTMWpNwJAFmKRbsbnsQHdd
A7B/ejVR30G4ivFznsRbV0X49HjrE4bOLFC6zdUwHQFZ5pQWefIkllFnXEWOdcXb0pJvX0AULAzK
COpKKvuyA5zvEjOir1PKyZ0vlw3uSbpb43/bCUF2cTwj+bW5MBe2Y08W5kzw31ZUOXFaB8hErOiR
dHN0cmB/InrYrY0kWVg6/0zUeOjI3qys6vlXZ4x71ZMS+ptdBPFDzG3X1k2vW7wwjSthdLJk4vIs
WLdvpXe8bROmatM9EQeyN60DCTSW9xkMCTaqiWTmipRUEeAw64MVd10xhthcipfDNEKTnYvdh+Bm
XkbWPHor5Vgj5ENbfY/ushYUByElcIwlvshKsC/b0Ypo2atIWCnmVF6qfX6VBzWsyzyCmkSwVaxd
QtO6veTExZDRkCngkRFf+nbcqS2yLJK0SBGhksF0hoUA5EpgFsx3py/n/f9OU9j0XYyo29yzq/xX
Ao8Xad97dbM93CiHDKN5DBU8qMtu0+hiQKkTamh1SmanriuKcPwALD+cYF3mkt964Rlj9pM14Lrb
aaUW3nVbppzsy/ubN1nFkvnzlLrBeDImY8pOnComJ3SOxtlH7DXjndXqoTksfIdEfMYGVFFoIMCb
Y26ErW0H3FpCyFVzG2KUnkxgxyVkdEUMbuBjsHa9ayCORahsvunCqy9u6onsRyIvUWaueBmhk1ux
2FNMvwDL0ewwZ/3pSQEGhL/uX0DGevsqpKVMGOqgg4zusdWtWwWX6Lwkda/IJTCmEX/ZZVVwV12i
MkqOiL0RbBwljd/Ja03pzVBmKKhmrjRz8f34oRpRrB+32mUvaQx+eDio3eqlRWf7h8QBp3APJT64
psT5zSiH0/nZgEVshYHWhyjszJspSS+roIN9BFMPe4QaQurUujr1+cS4j3QzDce/irs/+LYccMYu
0zd7etAg1bu5U5gmme80RPDMg0IZHSRrgGbAiySdaH8m/ctBYg4jxfYytFhX/2eFqTg267s8HAGJ
xk8JpwKhW2ad5dP28ise6W9Adxi790SR1qYrKkT04FPnLaKxlEOh9OdRAYyKDU7IA7v1s8OrRRtG
R9AxeMVYT45IK7SkRTfxJZFk7HSVx+jUcAyTaahR4Q6lThHs1DjeBndelhTKi2XQLYzPCmw3IcMe
8mn5jWG3RtB0QsBKFd0XSeKOhowInfYHgZsbeZ/2LbMxGbhz3QV2vZ4+jo1fSMv+/yrbU+mjsNka
lgbARf1DQX65kuzhgoq2s+ivZDhDZ2y3uDcATa9bc+OqWITnMzCZ2y6AaeBs6zJgXh7uhyzDT6/b
/+CpgW8fywdlVuXeIX37wUR2g/rexlHYd4TjCTb0aRia47deUkkgsuuIn4AQ1+15YDePJ5aRGAe9
O7dY0w/82wtSHMp6G1bj+n/ogsw8+jsCCRXdg8/aTOJJCnZOfiBPpyn/MFdSrBTd6sUkCEpfqglq
TFY2XMpU37xs/rObH58VZirbBRw0Wgz0XliH+bynZDEYxhMB14qsrSnQ3XqBXVafe9lHqJL6n0mT
a0dAyrXLCHjp0lpRTGwC3DUdQWCKHwvBtNafYIezA4uMc0D7zsbKKe88rnJ3OuAnStG3h/CGdgPN
R7hfyerCak1V5E2KOq+JOEWgTDF4pcojXpZhn/E+/jfb2hrVLWw3kN04ieQzhIsGzG7J1z9vtDf3
waYZUzOPOJIz5Juwec6W8zOaAL+u3GFrbVEwksEHRivy528+tMoL44zNmrAvgYdJd97tkzPIUjMl
Y7rkbQTMPDshaNiffXMVVfGe0FCaIqkUm3JBubHIcVhqNT7Iwx3pD58EIAP/stwnqvjFrH7amriZ
8mUyCQkFutkdi5tXomGfyjV9R2hrLUi5xNjuB+nK+z153diImY9hoQi82B/7JoqhpcYV4ungkhyg
Cww4O0rIileUd6+KodFW10hPYOQoIVksQSXBoCywIa0T5bLqQrqR9X5+6OpqwEkLH1t2cLpm+6D6
TJqnvwR9Mp2siJBQoHKyM2Xdeb5olZfwXf8NNmcR9FjqHrLDqXDL1J2ZzRiSbeqfxm3w/tCvKW1E
AHcmm6hf5YOtJN8f/1vVqVqnWjlUpiu1sU5XQenzYyWaydCeRCYiPzEhmb0aKW7qL27gmYZ2GVM9
7uNAiPyJvDY1RWznZrOomlbi5AwYK0OBohQfxoz7Q9GbWfh7u4ijojv3zIEq1STvzL1NwpfIenP/
mEf05iSAhck9N78Tho1NtHX6h6Pv9i6ZxMbBt5lZIxqyz1yRwzPqU9IOqze0wjoTlehp5G1xebn2
LYCynbws1G7pYKeUc5jSejN5kuyDDSk6VbXHUe6SZ5yPp7CfWUVK5FsSjs3zyGz1PVjaLAZ30t4S
QvS3MpmGcUYobt10pF6NihcqNDD9OKOPTH5qhu6mylvm3WkywnC2hviWlxbJf2XotPLKCTGN/weH
+aCSEl3KCwUdlzRqtimidPQDZZ7wLOSiQU2Kdr+BvJLAt2cUgEhKznhfdWnmbgVUt0nALUBVfUTF
HnViQKGD7GKRzKdOZeEbx+wRQCtFMfcAcHeMScvgivF0EItAueMsvEW9H8xc7jyKw5eJlHfXTUCR
//Fma2fX8Cx1bZGiSBnaPyYvZzNz1y2Ad0tFjS+kKGWYY3VJ0vYfy4EdRySXjVMhdjdxHlmyhjyw
aCJ4FAUshy3Y5hm/r/5eEKVb/pwNRTdEYp+17r1q2H9uLNa6Y/Uns9F2x+h1GFw3KihHciM3vNYE
zQ52l4SeGhZ24y40cWAXWdXTvgonvIXMKuM3eUPVlHhyQugDGa8mU9FU0cXBniNtMPHRefbbcgoS
v/9KWSafRzum4lxzOhagLTSI5T2TlGHqn/I4mmxKzMZyr6u1RNxQ/hAlbyRZCzQllr9gcSII8vJu
FHzTCs7CWkN2zbGo7DJNeUzy0zYhxNF3S7WotEwFl9CNPLWGAj7O13P8yC3Jos1oysCk22YylOYw
hzWjIbjveU+arAQCRVahEC5EnyMiSXyp9zmPUP0f5c9G7zREgCPA8JQIYv32DjApi8/lyVg4rsuj
CPehX8UqvKP6d9SoxTeGn77+Em9yYqBT7LkdzbqvafeedflVBUVrtdUe9z+5XEDxWOqWVaey3c5M
QQzvuwNeBfXGdraqpNjdz1fI6Qy6F5N+bJKrUYEzhg0hBUwJFt2e/VozkeCWqjOLCfe4rTNsAWQV
cAvXh26cgdUW0GpP1FsT9EYszaHIDe/VkYjzJiUnt3LJMywpigq6MP03ZR2pCAcAJAAPFTZJxDLi
vHci74GHzt1eWkVuK0E6vG5H9neHR033rFMmMFMNJb3T/72Zp5r1yE4LGLTF3v96qSsJye9oaNft
vl4sIfz2Y1RzKaRVolNsZKJHWHz7c6i1PbrZzB+aAZ6G4nOLgEwF8GgSUw9Rrmc5iDZGrMHvRM9q
FflQDWfOU1my0xh6MKvcZzUXxtfzlzZYbi8k/YENVUY+BT3lsLQYqrgToX9taLQnQ3lXXOkwZm/Q
0zrjYIB43cf4QqOcc5ZZunUjPalhzbW0Bv9z2oPJy2QbfqW+CxdpLP5XHfo6c0/0oblDiOgj5i0u
F2Q7nBLYIPvfahL+qceuXw9o642fFVW/9Al4ulRgvMFCgN9mpgsKv+EPlP8yD03gCWy/OEbK2sbT
JDgd9pY6FZ6WZ7MNf3J9dyAlgm+EinbjjczpriLle9AcbEUE0hhtADjXTlkB1/oZGtgs2GKQKfjK
KYL/H7CWuLCdwAo8L0yDYrrDxlXS0L6XmDzKMvnkKXyUjldX1245IxkzyxqycpdvrH/pyTYRXZ1W
9gNU4jsTo33Wy7klRM3Xl3AvxdHxJsVTYGw6snWUa6thxi9q4fd77KjCbI4x1eUxDhOFVNFE6r00
DnxyLffQoRSJqKjmYCqPdeE7bU8ZizqEtWYQalxKuUio2g2NnOUsy5fRdOsOPwrmqAVPAC75IY8x
+QTBqV7gswFHeF7iABAPG+ycwLAXG581mF7C/dvOqy/8twvSQc1ATDHOs8JgZ9I9tAHlEwvD06nY
cHPE5ihj4VyQGp/kRFW1tZh8bWg4nvRPo5zSgUaABt/RdJz3D0BPULg77TV3MPnY/NNdccDJlX/r
LR3L1iy2YqlzWO98alwxPHlhS4ez5Hp2/OQ6gVvt3peY9ZW0VBkkb6tm+K4astrJ2Il0Jp97q5UT
T2jx7fRimyIBSveX44DHAh7tE3L2Aw4/SXKVfaYrdbkSK7A4eFoJlVV2Jr9f/eyx1fsgAsb9B6jK
jz62KfItiJupnsRQjOE/Pgd3pnLneILDxy710XCOocr8/Pz9wkt3OgeC9JFMkSJUCsqjBxZoj9Ul
Lkq2K+7JDXcDkcMC6yNNtbw+hvpJXbmYBFsPtzhQXF8QxoD0jcSY/GRiyopTq8H9kFTu4RZDg7w2
g3A4MDLxIbgr4v2Vo/h18NaC2Jg0t+vCpzB6ETZM3JxBIR150en6t3rVAYZXl+DsRe7e5BuUccmt
mmEQApDQzrPQK7FXLCnDWz8nF8p4YV60rq4lChgF5WTa92IU+WLmzuirqlcoKpyuZ4hKvN7Y1QaQ
/+9X56dYSDBgxJlsxBzaptJ15pqp9aNAOcJIJDxfiF/m03we9cO9QL6i+s9Py/n0DlB9bMIRkmj8
6puC2LaG4vktW4Zuo+xE/Lrdfy2tZGia0pyR1M5c1TuJTGsIj92tcYuruNNzRAlBy9BtNN28DF7k
Rd2xZj+dEUdZwU1zFs9wmQ6fliYYOonyRXUeeIS6ws0GsLMMEvwNJSd7HpGcPaHXm3ijnWnaC0H1
tW00crborTyZ8eQCKG4HHzO0ndXYT93x6sT2jxXnM/Pd4xOlHPAKU6aXR2IFmERbcaRyaq5vGTDw
hR2qqY23QSZzQ6Cl1lNXv+ruNt6tcg8BGIl0Wr1PRW+KpW0sNBxTzCKDTikYycERMhoHtfFJAYlU
8dB7P8QOTHYrsQAdlcNjETFuhZ3pVR1RKzem6w14ZaHozBLYEsI/CX+SmwNU/r+hIuVwvM+m63/K
008x0tuK2nQGQdqE1ctARUvnd5itdNdU2oTLdfUZVw88xSHptvvfBQk6LKTdnkq3w7l4L+2lmWnz
Z/U73D1jTjQ3dXdYrVp0KvVvLk2f03xJuRN9XV9N1szlDGTGkYeQ9sth+5k5t7Bn0bT/7dHLKtmW
1QLM5o5dY/kZsX0hZKOkLAt8J5Cp+eupHUB3PZUQl8dlxpI6HSbhRgP4q65K23kZFj3q6970wgBG
nvULFz2Ii7oD7+pgawRHwngCTiCSigTNSxzMewRwEVJOxaYntzQqITFIrGo1t0akimnrf1HCNCmm
aiUIVLGjCvupHO+2L0SyxsOiS+Fu9nIgRbbsBYhQJ+5fAo8nF0CINSznjYKeKxHbufj7kG4vyAng
jYRfxJJbA05SkQRrRElCSpu9zyxdB/9zuowDZZuH31oXj37amfnAMhtyBGpEnphr1ypnNi+n3Gdw
4BoOOmOdIcspgANE4P/b+2FyEcDNX2wzxd6LYdZyGBiFIXHDms+/L8cURSCYCfo0T+NY/ggoZBBj
Tj7Bdv2/ZM6IwH8rfLUSQHm0TzXUZZtXujsVSzDa75ZTY4gH1w37869zXwZPzeCU90EMprlYM/Jc
fWUyMv2ClqjoBUIl36BQHY+9RpvDstxEW50YpTkznxcYL+In07mIbGGU+azVP2Swem/0tgO7oSV0
iVMsyODfhnluQjF7ExOPq5xPoSIxcn+M86s/IOdTbtM2k9jZs6K/4K9MxPTvBpDq1Y/Lo5+FtoCx
tQ525NoXIcPPZ4cbopFbPdvWeTeGVjtaTuh3Go1Q1lPEYG4qnGdTAVnmMZ+9587btiMZi9I5T1gN
B9BB1UyeXan1j/rSrxr/SyuUsaow1FZBwmFyTSVfgq4LeY66rPSQHbu6YmFfs9aBlPDoo6zHHgg3
sqE2B4hQf5MWP5xlPBecNJZQz+Py3E+LX/3ewBM7mYeH7MLh7Yvxw5DxmMnB2yiwpnhGwgtuAYKU
9JSe7mQlFfjXPx+AxzNxwqY+ScoTshmhcSKZNXkl4qEBEuDduSdwmsACMJn++/IqAhtRl/3duOEb
wwrlxWa9WlB0cXHWHFNKE/Ny+KBi5azCL8aW4r1S7RdpXAbV72Dgyo1JqCswC25QGqn0IpOtFR6E
jPlDLvwido4HKB93pwfkvgOz2hzdWliNmDcppnPn0Wm7HHoSn4pao48Ow3PezMo/xlPfLpAnYdeZ
fC5tygAwE+RMh+9ukon0i9voV4s+eLMYGHbuVU58yyS5qyn8kBAxnGEKO4x77HTRCPWITY2qPclZ
ANUHQqYvg/muGFpxqSgLa2Tt1tjNxbe2RFih/ePDfW1qwKpMVikRqqfdqaWu3SzRGgDjx90+rkQa
mUeuaVUVVA6bm0EjG07Qyt3ELVkZJK3CRf42jdfUdkhIiP94RenWAKcn+CWqBWufHQnlLMSiHgdb
ksNwLv/dmRL4pG3thkKji9hynOT7nTKvkNk5wq63Cyce01wMwzyAJsTiOyMpPgN1R+zNllFO+dKZ
CoZ/b/QDliKhsEZxUc+9Cbv1W+QBC2SPNxme3wb9gUhWUK6p73rh1btbgA8QeyDctZHB8ATrd+bb
h6iLXN8533pu4QaGGgBE7fDB81wAStFThXZn7RDn9xfTxZXH519Dvfq+5eq0yj1dA9QHGiYKU5PK
bciGQHJfTq5cRwI07YX/PU5UrAS145tFnmDcm+A/cSj1O0blwct9JVqDDgCxzxp09oQhnKTCdaUv
LdmXi1VXEmt3E6bBZfXeM/l1e+BOo1RGk8L+F4RMMYXeVXB0o/n3kRaqWd8PFQmU37VykWb0x7m8
VJfG5BbGXzWGBw10sUxM8m+1XiWsgBc9qfM0ulFWlM+0BQDxItQqoXxX2kBwSkkVLnWr0VkTEuz0
IkFuNGNcTauKy0fdSwnrbVgzb3Sc8KD1snBO7LK4UXLfFLNTiJ9VXOeRdZ19dImwP0zIzkBWoDFA
zA16Q0HfAzrPCub7v8lWNLHkoTE7SKCtQTMlbQLt7f4UUREjjtdP5NPj9p68zq2iri5oyF38/0ta
VGSrg90q85nHvYcaeyUOyhX/+zItzXGo4vrM02YTcbAgfiZDU+ac2Y0THio/MTU5WLRYtNDjEGGI
4R5p1pxMGfpjL+98F0h6QW9akPEnReCIcCf1MTco31XyW7XKWsegWja4GQnEZdFFEidAGze4PgBZ
J1fmIC0/icBSoqy+wnUEKlOyXyn/JkUeW3Izg2R2Z4DpkjkjfHP8KP0eJJUARR7PjaCfqeKwVxb+
grKpongEud7onmNbdJhkNtkIpeOLoAN0poxLD9Eum4pIo8GhGD/9genhL/I4+IXHmq7WZyVcHllv
XVRwDf9fF/VO30VMuZrNa9efnUEob2fqeilazPFguqnv4u4drKWtuyr9RCB+H3IZVYkHyy+q2O3y
/Fs0NuHURcKG1kYuaH819Uz9vgkSM6XVU6+XlTmFbOgSejRNMZtZZzSK2l9mTDjy0lv3qTeiYtGQ
x+jckUNQe5Qkr5ROVrSSAVuCjsznGISRK0+J/cvnuX6OJorTa7EdyaQt4eubZu7DcPUAuB2iNRXu
lIS3PAZMb7z/FgIHRU9jeKrP8HCY98mKLrdQZXkS57cvfcJI5oUyhYm8/YsNqZf/blo0u4qHmP3h
lUesFWKqxdifCowQ/xVKfSrzj14ndHW7ELHmLZECBAGlFT5uJvuIaMBXPvoeMo1Q0FDeyH1PCAca
H+DxZ8DAKUjiy/4nFmuAiowF/blIBTyD72D3XRgLb+iMiWuc2IkJLsYNXLTZs/vjzrYgqF9xPc4D
omNBjbUYW5g4EddsF4cfcZBO1GFB5h6GCDVUWMaqD/0/VY7g0Nkmjqfuqtw8ggVyL0EaMW6VHTsN
SnMe/xPNgrCCgF5sFj1EVi+4DoP7jh9im6CXiGcLuJvQdVloVH5uKOo9PcwFgJbSz0JMhw1XMeb4
EkRBwjLqrLTXcfrxDai+oczmZ9r0mHaQ0ibw9/RbhLPC3LTDJcZBmfiYP7IWsupabpIxanaTNmUN
8NwL0mo/CREpjqynI/U2UeQYZz16rKtcLiRUWE1KNciORufZOl/osmkVCiFaDArRLm2rnHFSe4eT
irYqBRe/wu2f2+205CevXNISbOwFLPmDrwS3+Utbn5p3E4y97IBj8c7KL+hqC/7WC8Un91620Vq5
5+XOy+qfYbfok7ZG5XkbId/LYmkG2fSb6ZMzEp5MndBGHg2YsfgDumPxbH9zFzlviMM1uHjP/dS7
mnT5cfnkd/v239TKovPEo+DNM3ieLNqyIpGOzBAcIJ1UHZgDwHtLl3/EQtBg8MIIsANy4XANVOTP
p9YEG5AEU3AveaKDJ3Aqn+uKSebvu8jkFYzC5KPPoFGBFu0f5SwNAZavOEYqD2d5BOHJK5Fg/3y+
rb6chMhRjEqLNe4A2r3v/Yg9vUxxPtJROBAMXcqPZWClO5eHpuI/FSkaY6ZATPciSysH/vsINgdm
yzpf2j3GEJmkQu7L6DAeINxFBGvASXyekT/9j6EoGZ8n0Ttpyutldyp9lqbj0n/yPoE6BgAm4Y8p
wNwSbwaiATI3RL2nmAcHJJM8Y42yLw89sroQ1+JaQaSPu7dghA4XO1BxVnzDXcJuQgL3IHf9Dy4c
ENWPF9Ns/JKO6d2NMLKH77oA9f6KD/fMcM4oAA3tJrApaX0NTSIiowtcF2+Odqt6zjKMdBjeYKlU
25ZBDGetQMlK7gdFjRmn+80qkoi0xJ6N4/e64dhPzIkYqD88Mxc6mYSt+3pmGTZlfrXWLNBaOpdR
/PmbKtWOWwCMm5RwYy8GYhjW99a+ZTDQDx3otyKUztvR7pSbOkMFMPT+tAxBGnb9QZjk55xX+s5k
TRkzyys/k0uTqnb39Tq2TF6mf18X8KfWqKxOW6c4eAUng+2bOn0aZ5qLefZdEzBts6NnFHdA0zM2
otAzd6u1WfDQDJwo5TloWwJzD3CcoUbM68vJX+qB80wZyBTy14TfxgnO2kygLlRqVJvtfsHGzmaE
UC5jER3DqR3VM2w0vK7PNjOz2pEiORUEBfjeY+InUA2lu/V4TyluRvZTTqTZn3TxE0urnFHMpmpp
Q/dJarnji05p/bVnNH+/JoSFhQThzn9Kr2yA6C2imZk/TC8yKyIQ/rlB8hJ0KZlDuk52onKWxeG9
gboLtt6U/dGsfXseT8BxDBba3zRzo2Eu5pA3L6VE50hr5JuXWltB12ZTq6z5JHbn8NC0pPvuLAvf
sm30zDtUhsaw2V1yvPlBClN0ozqhtsOCzX3DzTp5xHAbjcj9g8PFAMrM2lwDm4rgi744MmKlaWoW
8FBf4bUrNOUgL7RVZyfUmq/ZFZVjkcHiFp/gF8/BloPIlYu3sLgLJMxBqclk5cG/mQe6PYCqfpnv
lt08iHvz7QQcapDk6fm94DSywzZWh1aLlDfhofSd74EOfXBHuM8+onxBm24cPwWqS5D9BCN4ITf3
s4bOJyO7rYpzFP0r9HD2T8cy9RNxrL2TLEBW3xgAhcIAjUCe3+AU8tvTkwU3lN3M7B985HsY8Utu
HjGYIbmtVubuzYPWNZgjFErH6zNG4kzf7/fplVihnxSIPZaR9eV6hNT6DaWv2r3h46h6H/zXVEqo
00fiD9f56+Z7S4aTrLkhgnPtxDjcvREBG9gK+yCSeUIHcVh/zWRjv8AP61BJGIIdtUSyrSZN2qTT
JVCj9fkRq7TLkqGIX1WggyJQLWHI9MrM0l1uNvnuqQj7LCXLTyLtwTleMDPxcnq4mD8GfOEFwKwq
R2hzglXnnlndiGeQUbJGmPrMZP75790Y3Ts1oX/P+Jd9vi/yxxjALVfGPnBEKEYjFgISS30wj55n
qLcFrTDaelVzagPkrQrWlQXsVN82fgi32LKeqX/y62x3HtlJFZrOREUWsK4RO9yrDK9hdIarbPn5
ZlIU45THI2nU3HhEpaHf+X0KkNw7TxK/KzAf7/IuqkO1ZxmYxg35m4AF0sXxqEz/Cn5pP29BZJ6f
jS+Kg1tHnBipGjM38WLdQrj4U6olBz/6Ag32ghatkHmyeJvD5kArtL+XO0hxw0sHwd7rvRSlVkVM
GS9ULVKwjbaXl8HAEofp49pwlSmVUzpcn/mWfrUQ3E6JT2HeZIqge7e10arlo/scUloWyejx5bw7
pevWNy0q2Tpx8NvCGkwM0A2lgIZrbGfRbVMN3Vpv3ztDbvzuj7Uj3OxNK8r5vEI0Bj/GpIJVGS+a
QiUXosa5F1C5HNIPpbaq6jjFvnvX4YEk96b2mAQehVX6FoNUKMFrFOoz3D6Rc4EcfnvA7kDsY0jm
yMP9D2NF+du0qjxdorH0Rh1cyFK7nKxDPpXPEeduM+/V7sTDEULmrV7j1HPwW022tQeRcGGkE455
T1RE1uqGXKc4ujiaugJ3jsJfCN9KDJxO5zefFGGH+JFR/lR8z7ty1oICIGnTWdQe/NPxTsaYrB69
xGg2tYQjP+beokgWMHjRgadm/KDF+G6UYVPRPflXt0in3DS8q8QAvB/X7evkrjqhbKRp+DWMB8aD
YW24X91s7XceXrepIqZZZs9qQkgVultTDIL3g6K23/nNiCXZjtESW4IYBp8tZZkY945OLVZrUqfa
+XNh3j+quCRGF7zSnIm1ZuPxb//cIXxfsoX2+AbcPsKpfNwlAdoF6EcC/0ggofPYP7Daif/4dAPY
46Xj4PnPcJNPt06zAe9uBBMg9nfPB34Dk2A/5m3vaYvo84uajkiNchrUPcN2vKacSaVnoLFw1tMK
QEuOowJLSzz3CYLPg9/DZDzZkAVOlsZyt/zXxxKlk4aRqyhQXJ3doQiA4eKwPww12Yr642r0FKKY
u76yVSg4zlt9u1FFvN4+EUNuW6coFwg99TEfvvRqHpGtl4wbU6i2n/I5oXyeGxiCVOgUTc0Aa/qB
x4So/3+1m9A+Y379cWH6eW/mZleCTxG7HoZZPOPVx6c9bWorDldI+c5aYUJLXVjcoYKjbXYLLm1b
9vzjJuchSyZM2/NlnxdJo55dLt2u8SfU/UFpgfQUGhEW5gnrDdbcTsodMTwqHilTfSFJ5bwSmQvd
GBYZ/zWq7lLbcBZzQJirXzT5+DgRtgripm7060kAB9YUmX9RurTcttnUdxBm7/O+1lfCC1IpyCbl
WJv9WUBsn8jN2eFrBBVpGNi+zpvYAsaNrI9oM7ieIi206n25RWZMDOBWZAx/qFEpbc10yvhZfVH0
3Ng3sXRhIZZ5A4uNJ9uNq+PdhYHB+nY4i2dDIqz9Kg5OTQ3SEcwtiNBlh9qnRA2Eho578YbFNXiG
MqGLktIdNE7jc/XsTRYqGcXnPZMnN2oj/X0gKSqSsAunACm68a/U65xIBFnC1EC4SctovhVqIS82
AmPXMOJxgEbuAm8U3JAk1rKx/oFJgohOi9J1lYgcSESFwOfzDwGoaDfcJG54x5RUUAbsn5dIUNO3
qW9VRX10z/PsxhcuCeSAHiWI5xiaAqgiPX1NxxYdQzAMRGvl+22xGBNs0EyDWSvTEbQZ6xqs/f/b
GhF8A9w5N1NLauTd5njmOHSLN0njOOiypW0B1Q0t5wgTcbdPAPqEUViHn7mEN+ZjJxmjIrOhQZOr
+6/8iv1z+0xJAZPfFsJJ4FdoCZ0GpWn/zRsAM68aiNjpMByfjG/lQnBYfjxuDmK51kRaUv6mmwa6
un3agwbgLTPx7rWIOykHdWGndUS21vPkl7s9Bn7q5PGU+Fftq/r5DrOevGGdQV9N3XXojF89PNFm
1ZzHnWGugE+8I4HWxSFI2JUkpGoO+cUnOrYY+qwYnfpGtCoFbqVKSKGatgDsgF+OmhNaGEvQVjuR
wgNmGRHbKEimqC5kQj3v8n6WL+8kjIGzMvXHojHWcLWm7wXU2ReOKi9MVXQ5VWlbl3JC+RUvMiLV
9DWaBMiDiBbSl0EW4A5aKa2UiQI9rJnEiP0WiudwnMDYttc93XacjHfIqTOs6ozTxeENqqU5OrFj
Rz5IzRoaw9KJP2tMZ7kb1zDiC48rSYr9P+kgItSRs2VL5K+LLm3/Ay1RsI6DgDBa5oHIbLTyeMPn
SqZ6Gl/bYzz90/ViO/yyPs92dOTn8eNh4Xb9mG+H/LIN2cZv4yrxIzFdbqo/gJoJlcw6Lv5vpJtV
GipKlHb0O9T/ZAWmtGXWigdyBx4izXIl8fSCqlk3xIy+UuRjZLK02bk11ssWyYdGuWzT9N1c1yNi
QNeN+N1ZmCHfyjFQmdtKCi17TqFelPxsF08NYNg3zfN7Odt/4Rwz2XZBu6vxsXY2HFRowc9zVsYr
WR38SZFhGvmzDkM8StBUZiKUcryrK7y/kMwoh77lr5VZTDP0IlZQ+zvc+9bMahv6gAGUPvWVnr9D
D5lEX1rDio79crgweJQuVqiAj+7fsL9knRJYGzJgKqZ9I0fN2+8+XleHW3lS14bbXnxATRkUXbc2
9PuJIrECp+z8NMd5mj75KVSTli2BJS+7GlV0t6rThOITmEFqm1ONyR2iK6Nx9yi3RIR/gudcXPsq
ju7a0ncERTusILDsAxuLV5UPzBZL2iML5e8KBeDdke2thxZUj9OKtzTQC1POcLU6uq9EjxIebOtB
RDhLqR5Ki47oYX3pLzpRSKd5ukVmzXIl7lcaSQKlQdC7BdSR91fnrGKY0/pjIdBU6IaOo6YlBbv3
W2YskbDk/TNwyO1WWbPzgxfMzr2wMlOeT+DJIgJjr9I3F+AZmQrOZ+H/bXYGSYiXCna8NkRxFdh7
SbKoOh/7RwLvJP/4m9KXL1dj6kITVeA6kc1xPo4OpbdFBu597sa39bngN2luxyQ1vca4ccEoGDjl
b8Rn3EXkMpCxkzkh/vfnaxB2+9mvIEtwmdZZSPjtGVfEpMCN4y/coFVgcnVRYkf4WncjZeFY09TY
gdxixKaDmuR9cYGTpvQCshHoDmRpQWedLdI7AKDKlyzKabcQvl8h7ibUcGGOpCDSnTNeOIph3V1z
whpVDtKNoL9pDV9ZiD5srpD/dsGd8TLR3byvvZ0fS3q2yRomtEhQrQ6D/PbXalYVWQEIyG2RNcy3
TwPkVljbdefHQcUni6SqHkBKmI5ksqHHpvnhxGePjm68xyrL7jnnQvCPcK+RcyIZAzz0c/64ijbT
Bo2y+6pjCW7Hb7geRCEVauHLqmDtPmVJOK/90xQn+E39EyYykW1TnjsfCl28z78pYEJndo9mYrMX
AEAIKAsCZ7Cfm0x4gGqeN8s94lvlrB6hIX31KcjY792PwYAb09ySVLUwVOazJYbO+uDOgAyLE7fd
UUirXOReByOZ+3cTTIBMR5hsTlYlh7Eo5sf6gyuUaKg1UgLtzNap363md5PuqiLBM7WQCpI4zYfj
fo9+moY1oPXFQOgPyxFbSavEaFuocveO2OCtws5AgW7pSsX1n0fQrW6u4SodPpaKYmMBTNWja3BW
XadIvW5sDpDzRIuRTE9u1tYP9Vu1ZQkdRbptu21MJZB28Jz1LBCj/L2yQ/HnFjg5/u8Kpk6bdlvZ
nL5IxTqY8snCSEGenLxdHw5G4gEG2dTA/14TRq1JR/YP10IbpEYsembWR1JtCobGshXcKC2gmBKa
3v4nFEz2QxUHVD1tK43j24FmVZJ4ND7Zc42/f/oD3rp3gGcmZ5/pN0vuqGRiAxeMWd589bWIEmWk
B6DTRIudQaa7JdXgP93D1lkYWKHPXPOobDzZDzRSOaOLcMtJbkmD/GI/Gf1ARw4h8wTpmJqZOyBu
hH0IhHFxqf3uP3If0VEa+3QYHGPY+mV0Becb087ZSQRAN8gL5yCquDd0HdrHFudSroDGZUeiTmmh
nomPgwXlIuvioM2ScDnEyENF9m3xEZ2BKd9vzAknG8TFqrLITUU5qBg1sKIuhZdYFfX9SCys9nGH
alJ6abpGP9fjm8hPwarm+L9MTQ0sYOx4VHoTiPvTuclFmgxUC80tMGx77/mbU+TpI0jY8JYfyyIz
btky5hoyUEbgJGLZ+h7DK8J9VzMu2X42Z6V0JfTm41gVq6txp7zRUqDzmDh7Fnbi8nclK24YhwUt
ef5U2N5xLY7bzm7XYZITBJD2FY8RoHyP49v6vUELJzrchQLsBEGazIilvCfuNSA9J0UvX/Hp+tC1
uxGSc1l9lEAPaCm5lIXtfhPKuiy9agsLaX0oATil7I4M48aPJ8rhnuksTPIGkU36GJBI9At3ku4J
ehaDbirsCBdisH8XBhLMp2I9tx1Qfxt9+rQaUSS/Rwk69r3yEBBfcuXaII2M8OW0VpvTmICjqP/I
EyN8j1NOG0OtJfyWJR9aHKQBzig/1F1sbiZ4ozVkdc5Lp+cOmzpbXSVIi5c4C77r4Ez4jmzYjKdp
DMKdtpnXey5mZKBQZikIJi4GOtITqs7UKnPJ4nV1NWqOH0lFrl1zJUxNwRcczOe6xb7hcKOjbxQW
WF1ILm2de0ku/dOGbzFGDm6QF/VkIyc+HwSvIPyS0Dd9N1YRsEotOT7WaPZBuZ8LjSmZImcRf/Cq
+Jm9Vyjc1/sPsCXCLQxhFLHgPGmm25b5FClpK/R73NgTbLVy/NtUn0eB2Mv5yfySLNAn0Wg0T1I0
itq8fVlMnb85rQLXlYsK5zO3YByb07aGy2MJ8erWqUq/2zM4F2KHLb0plBTl48Uwcozun4uCCPDf
4voHifWcMctDGT5nPaBAYxGOIRI8HjvErij65Y672qPNdoySWUuz6v50DIY4LSRuGoGCSLsWqPNU
1I3Q2SPtLpORVciiAC+OQCFcw7FwK9OBL2CVsmj5KWvxZmfyYFvOOa4VAy/yuw3G0PLJiFdnzb8J
b6GSkTREA/gthf2J2K2aHRMcr7CxiqCzwRIvLbINCmK2XziXHliDvesBC0ExKJx41y6Fr+SrneYp
IAXqoKK+iu8VVDfPPRmZNVwECW0Ayd04/WCF/d3ebuflKT5E6SuLVnNlmqha7J9TB1/pLbGB21I0
NPtEHiLNzH37bFHxTnwM1GzGJfRTG4gCmLQYp5qUxMhxwYjAxaAJlT+EgO42eYuj2wMKVJm+N7Qf
AC3SlKyqyBSD90HpJzVD/AMJYzrbr5KOqFlSm1C73GDOE1+D7OYOMziyqBNm9XYfM4aIu0hMTsLK
/7DrP1vT5rweWY4QafZouxgGf6q9NTwJ8CmkdSCjcPh8/qKQzq8kdjhlF86KmFcT8us9dP8XprCJ
zIrq5TwNtKwhx4W8z7QTnj6IIpqO13DaRBBVLIsRQJlLXdsUhqEJ+EHY1v4sjNoFylQw3WSyOKE5
5GkfU3xCEe8vXlPDEIqWtjUxNLFu/wj1PzFU5p8TVMnaWRyN866O/k+Uvfx5s20A4njLhsjV30DH
dcOTtAiFstEcdKktWgG5EjbBPpmK8pf5FkSMOD0U0Ez99zvaXJIWQ8E4cUT+1Aam+aHw7vYmiU9f
N+WvhRqG7LO1UWShAjajLw2KwSG/NHoa3yqdsTq/b0IqjnwCIMH25HDebuQTKasWAkyeQQGVNZ45
iTYydswhxDY3/0tLcRhLv499q20kwpisAGjP8O5E2AFrPqsX40c+PA0uCX2ZEBwdKMc65rPOZYpz
brpcxfVwNW0BYHrcoUQ867k8QeZ7ENwJ3czl4O0H4IAy1NxfHfEJKzcxahapCWc/3lBL4glnNGnS
8s88FrH2xYeTNKZfZnpNieJJrLrYS3IjvReD4tLa1+btwMx1Sm8jhokMVMEvQWtk8XVsoiRFZduD
wdX0+ivGhkbhG/AhZwqiX7TzpXiPefDXLcWYRnGFVbd2UVwanEgMEXO5kqQZYt1wwgKISxFGqA8+
1Ve8MOxRC/lL2qtTi6yAX6mtt3NPMU1CkksxY8WVfvkr7t/5JlBMKh7nBsiQg9KfCmtDsl8087yc
/W1hL79qGirzK4DfZujDKKnD34D3LA2WJy/xHhma3hbftjgPuUX1tVTDUlyHMu/V/VWXGkLcEN0M
1wlaIDMILG+jqsn4wIC2FXQqAm7/v4YTKlxKHYUUuaOJ+EP8S6ATulpX0LJ5VYpNjEMuFN7+rzE1
TXm+zxpaR2XG8WPHcQetevQrOb4MhLh1eZ75nuYQjRYsKgNBflCBwcMaztPACSplV5aK2THxwVOw
K8BrDp0ca95lj7spLZRyWZa3xfDk9OfO3y3qBlxnWrHfmgqj2FBdFd03sRnmPctMHmcQEsEOW+yL
S8NcYWwMAGwIfPld9SUVFu3sVJQe6z3RzYcoBH8+LPCrPXLqsPz8usX6eQaACQ0Rhyr6iq8a4LCn
fy727iPUEf4Vps5MkucqFcgFlolT87JMqjkdtAcf7ZUl4DmXRgm4wA0xXyG23b1uKwxJWEBElBz/
kJkjmbCuiYQCk71Jzhg0cIqG7tpmK3wEK/ZLvXQkxPEbkn+ANUB4MJZNVq4X6Hijjb8/konGCVER
H8yHE1Oe5gvjICr4C3riaq1C/MbV7cmMZa1IeYehUwVOWhfi0kUfcWhIKj13FBunqlwKsMILgDZT
4d+S+V2OCAbHTFUPhACJRRfTS0TmrEMkVo2ezwN6tlnQOrVMLO84jYgLM5xKFXiI07COSb4QPv06
3ooNrzFbuZMlIAC7h2Izs3bLxobYB/P7x70ZFqdg35Ua/xo2fiVE/HPeyAQ6764E+8zYlVvcQgPh
xkCAXeSpJvi+XvxKTZ3feTRU0OvAqy0pc+U+1IZxiWdoin75bsqkECSnFsb8Xh/DXQc2TmxXaLrR
cWut6Td5ViFmDIhzAum09lvo0qrVwRC3RH2E6eA/I+tffgsp80E9Q94DKIsulcKolVWmod3Pj+0J
rXkiEDjk5uIBo758qWc1MgIr1MMWI4UHIhMSszQao2nl1MrXDbbTeJA8Y5uMiZmKzoavKFLG0och
sHicb+Gesn78wsT8JUApSKLnHdEa1+XoDaCdcpPHf2qnSeNWaq/zUMei82idOTqm0E6PwBJy61Ta
REf6rhwTzhQxT1aJ5u5yZunEuKzqq/Q14z7RJIKNG8klNLXYa+wnBdnY7MKJKWI2uvpLgm5zF+/F
pxYOx52v9WjMr4WRS0BfXNLlXtcQBVzJOhMQ35KTtQD4ickOHxzSZK6F5wKOvXbIKsDQL366VASF
wYaSyOZ3B3belC0nBV37ikLtFjcLvEdbBsMjtQDieX06t/udqWGK/vIexOAo5GT9GvuOzvd+72RC
YAtQZqoGAZzi0xNM+Zd8HimlbyKF2bByVw8CBznnNnzHX2mywCH5gAVnogtGFXRkdT7QXNrCBQRS
3LSbpHQ1eIYt4gs2Ue2yo/zdYDMxq/PHUboIFFobOG0eM1oM8zdQnnySV4pWcECChvCvixZ+uA59
4Hwol5eIsWafTez7F+kFuO9lt8vDktTQpoRRH/Pvymm7KcFbuNOdMjWD3YFC0hNzmt5fEE69r+0J
US6RCwfmS0RgWoV65FSlWcAI6R0a4y5JCRkGnwTEnkuk/cZUQ8Y1wuG2xMCHQ0r9GWhTEv6inrma
qJuLrZa9QWLd1mlDOY5mVN/F6KIYZJ6I+Z22Dw5UxH+YHUFT0gq634JgiWSJNsdSMQhz2poMS+Bs
cXt6CREiUR5cF2yrVThKlb+aleILbG0++ucPq1/z72/v5Kt1q/iD92LssocwqkySX/rB5aMKMFFT
tzfFYANPKdZIAet3FKBSoCbrjJrEIu/tKD1aZjDBAyTzXrF/9TtVf1EnPXl30bhn6dhBrHQfHJ26
PzyZTqjAH9lMQLoIjw9QrBU/LlNgPJP+ez1Ry1f4bwm1L9yUneG9FalDzvutOmLJoRy8LoGJXvZe
LrkYOI8tAYlPXDIescyUqalkMUj2yGp+uHbiNRjLSuIkvjKiYry+h8lvelJNcN3USBiBijwUfoe8
8IWM6W6fWofSXceeVVGWIuo3OHOU/24Tp9OnQ0WcQVsNqabDNNidcaxN9d0ZibsZJRTjKOZ3MYUG
kW2yzUsnADyFGWAOZTkiuHGGhkGfz4mkwRA9GxceWL4DnvRfu1BZFeLaHYp8H5k203ct0fdae4RT
9dhEYRXwRvP616vpF8MV5O3arVsFH+8PUsuRYp0FOPTh16sahB04IiAg98p5BA/TENv5+E/Nt5N+
KSsRkcTYZ8p/QdtOygFVZn5HWVLEC3VicJVI1Q0iNAePR/9MmK2Puy641yXuxCAV56dYQLRWHP//
lX6pQ59KCzKSWBR7rgHV0FP8CQK60w5wryf6O5Owk1nIU/FDfs651uv9ArMeBj1PxbDKK62IkA0D
QGa4jTW1nzvQHr7E4DI0mp8sdxCKvoiUQuxNZLeS8vFFD+ljtckYuCaMj4MEdVkyKIcxwCAjUJ1J
JkwRCdGwO5Imls5D2o4d41L1z7p4D2t1nKJpU/AcLGyOF0yhNYDSHFMjpJT58n7WEvoJAWxGNOpa
QYvjyISmX4YkGbyPqMChFiSKMMITsytNkPlDNVqdLOOf9RLjfz9ogusAwS7RN3LPqRIs5SGYOIH8
NMf+qHYCvJnlcT1yMK6P9Kwk2CeqWpWytmHNM181debVjqmQhkSo0BXxvMPBq54PbIHaVZu1tBqQ
qcH0ob0+iOIrbJ7TLx2qgO8XkSR8ahwPcFTSlrhQifjC2pUlBOO6lSo879zznkihTTudektAk5aT
/ahrp/Zdtw869Dv6ZPqaC4qnKjVJ5SwQ554tyqM5CJPADDJ4QQgs1stPeZqH+BrhYMIHsSBg1ztQ
zERqqSU/ZP2bmTbgaKBt0wr5CLPBFKFIaeIWvWXa70uRlWtdsbcCG1yWR+myDQ714cc+opM6bkfR
TLvOO/j/46+kEo7O1x5GmTL2A6YZ05xf1PJ5NT1D4mKs5By1XGDRQ2g+J9RXeq8Zl0gxhUHwU5XD
JvhW3pra/ri2ex5Gp8DH4S5vuj0KBTHCXupSjgqsn5ll1vprWysFXpjT2SMiEPeUvqL2PrrlX2pQ
DKGyk1akZkYSh9G4eNgnF7hxQYfUDhGX+I/o+YQPn77u8DdcLHltKpJV0L64E2YYqThYwlcy0XG2
ujbiGJctEkDqmKmE7O7aiQDyP030C29yG1b/oi28ia4bnMyGKSv/Zp5l6SHvy/cv4IVGvSiX/MzY
UkKAluz4Qxm3DU3xFCmTN5cEbteSEJ6rnGkWNGEQPpbakX8uyxt1fb/kx5EHFhcc02RUjrJXdXus
1azZ7L2YN7+JSHsT4M7JOEUVTmwZhyHcrKxezHjadD9oLo8ZqyECA5dYjzIZ//MOPiR801wRyY7B
zgfMq6GzywjZVxDjuzyiW+aS87Lts7pPQTZ8BF2euEhwd46z8LsIHFeFhH8ejXbd2e3d+kjomtFM
6u/Ctltqe5v292D/bjywZOxX5wCFRlp5WTZSosKO8CLLc/SYLE/NR1qo3ay6AxkLVs6eJbUTsUlT
HQ2K3MasDMJ5GfaaVcZn+OqfJiPIqb46Huk4OHL+59dXfOdrlkN7L1HMPqfoxGajehyahIoSFn+I
Uo2qpNnYh3/lV63pPLmmqXlW1qJ8TH0b8W8RZDo24FW4b8lVHVUsVCiSkvcmjqcbviZ0UcDyM/4P
tYdWZF5E4/vvo+ydvE7MtQ6EbqlWtKi52bCK51VqOm1TCoFmAUF+oMX17SDZcV2ycuNDTWIs4AIK
XfY42vQ4sTH7sBYnRF/F5+311W0LJzvt397eCoiY4NeS2Vy5XqKZBQE3PJvdeJByMb+8kLLKCuwE
GEGdWFm1zAmtKUdrsQnwcAwqxTjiyK8aavb4XKZZ6h9+66ZzOW3QUQ3gNC5n2mxveQgoBI6nD6I8
j0FXAwqVqpJjZhfyhl3shjjmP4nIgBu91PjEUTI01SDm0ycMjT4kkB/dkJ2TQ7kculZ442AabyBH
mqzjz5qwvxDeuEVxCJqR1EkQRW71Q695/TscxLlDEQLbqzBACZy+XwBs//gONMsmzj5lJdHx0NkA
nlubqWaZx5fGRe+fR/vSYVgi8z34lxbGvBoxlVSG6lWcx0VICaTnJLa2Y20T6M2KeW02P6arx+J9
axjMTmxo4HjQxr99SWPO4h1qCaXPPVhUof5xtuKSjnTHjZlctMSVtkU3r0B+WWyDsMaf/x7bWrEr
xSImd1/MfIJIDXHi9da5M2RAKPLqtGQRZv1kGChDpDGgTftwGageZRjDBF6zndyb4gW2H1yrNeT1
PGThC4WPmAz22orlcM4BIzDAUk9rbS+9hOTW068ulw31HXy+phnuTbTUH2oYiBp0aqQm849yICEd
SAQS3T/OL9Zi5/xpowgyneZiTCc3jsVkIa1ZK3jUa4xN6UiCNaH8miKfqydwRUBVZfktRvyJUJp5
HDNg7cArVpkawwRUM+v42gVdeerlt+EhFoN9AlO7VDRW68LMdJW8Nk713PWTQx7wP+DlR0q0ZJVp
1vaRUDw2btwywU2jgKSkyn0axwnNLO/GYJ0nq8U9C6dofaUGy8LGwkZ2ZuUuzrZFHRNn79Cu8FP0
+Yh3do6bEYepAd7a7TvjQ5ebnlMCE9FmRjMcvb4kH1xZQrWUYouG67e3dueKzoMwiRuu5S81egBr
Wor6DSqkBgIeZ1/1kP4yZuYerc6nS0hpuNakl7DtCfwgDygNLXEerq2Y+URSnPC1vpvTx4rLX8hx
gbYARU9+waDMSz5vaGechRJTr4QDW5tnL7PiY3sI/zY1Ffm3u0FhcgWuSm/OpwSGaJXm5rkSmoRU
cap9QWTt2PP8DZhqdr4xpjOl00yCAVuDARdTjYM2Bq87XsFeJxpp+stjhHbpHO7HuoM6qArsKciV
GuagMVhR5Fx32Ns197Tkwo5TwuKa0G1DooBCJxp/yXBpg4yxWcxdMPXMam2n0IddOxMMWIG5xak/
RDjkKt7KS1Okxp5ffYo3hjAs+Q1C3KPnxy1Y21hiZkzjtIl+3VuuHcOXrGit6zLj3it/XUAK/2k2
X419IAb/l9tMEg4JifswDjsHulXLEZcJn1+PYKgzAjKYjxOctjx+eAupt+AkW6lJpAzJHlLfoMyn
XQgWr1nxl6iW8YqQRNl638FWP9t8I7HePvxw1paK/0PEb5h5aADSHzsOGbYCyRJQML3oTLf5aX5Q
KQ2s3/Z/eo6mzMQ5c+fgURwcJivjy0ANgshOQyH5P/8Vk6pCJSO3C5HlmxjyU4fv/9pUapGiG0df
noj0j7ab+xQNuRr/qob6A99M6zfq6yvhr4B68kWfLBlPbefgZ37JfjPdFMyfgc6qYruWo06CsMcu
dYz/9nxAAC4Al7jpyE2dbzLW2JVox3OacWoKLUOF1MgzWGBkUyn/Dg7tR0NOqnyi9sdbzb8eiVDc
RGUl6Q/04ahgay9CDXZgSeHf8AZLXY1uLM2Qkkd4k6lf9trh2ly/xKUL0JdXwg4e7LjzKDFnZ1AU
6YSlPLx28ajqZnsVQnr/IpdVG4aSSCk2JKs1Nlqh/23TL9JNhBvvl4mYCSbPjG5ljHCS9hW7jgeg
Lsll8VEjN7Fe2GYcGnapgNZrDhOcFilWaYhUMxdDEw2SP12hc+qaXyGmwceWMHkJJ4aVSTpVtbns
KqwHvmW7EyEwkiNpP1A4Qw1ghkuBznLPyd17gK8sO3dVD+5ptsc1tBiywD4AFJ3F5o0cV/4JgWW9
tnhv5Mm8+rZ0+PF0ZJ8mGQ8vyYRy/FPVuwuZXriWG1B/KZijim9EYO4tGvmy0GbJN4FD/3udGRS5
kJz/l0yqn/tAFUNnvgWGYkrapdVfHOByOwl/Lg/7O8nFm1rnkmI1eyu7QFRDoEAqiRU1FwypfUmm
we6N34oyHTVjSueaZWAsg/9/n447LYAEcIbvC4F7RL7dGxh2pFYU53oc66EihHJckXTSdDm1lbYm
VFQkfEcz+7VRTQ3MFB/ra4rXxDUipx2JxtdVhgX0fRVxl7ufmMtKFhoNiQscBDNUjEnNfNtXrFIz
aGIcMYhLbutBPH/zJavJzHYrwXYAVEe0426CiUDR0fEuO678DkFXSfeuF2eOZ8WiY9NHiXBWyG2t
kqj0oi/IOQBMZanTGY4MoDQkwyxNu0rjebDXQRMJr+R4mqHwW5gJnknK6Iv7yrDAQ8+QGUM7G267
m/8gI1uLaZkPzT/5h/16OJsbCs9RXHUAiygzxVttjchqbS8pjARWuGxTH3b1ldr0jHex5kn6OdmG
n3QspU906tC85IBeJOYsXOEkPIrTkiKb26j8Gl/Z+bzS47InS3OLZNhvOPdyqed3UU5Bp9HbqKef
tb8XFwDrTpRk4veBP0ojdjAMeJ5uIFrTVI1e5x7SPwyuTDbZa3nKF/lMUxqlu9EvUnKtscxL3vc7
3I4OffUNrk6AG0xWdNN4m4XUZ/+KHOLnd6tSK5OthqcwbwfqQxwkZFHX5lx1Ca+HhG+jEe9VZvvm
YtZZSpqcUyG3aovi62pgkjcKRUCJooBJdmBVRNJftyIJea/duGVSK60cBJ+x2O2s2p0MHbvHjYn2
kaQjra34NCBFmwnBA0ZFm0XZAS3iLBBqvdRoR34xtBWnL36/m1mDcSvZaQ8l1B4fDOnf5oK1dA1h
qHTNRaVu0JFPxFk14tRFXeDoV8kKbeJwlY255CF813PjQ7P4PVs/xGOZr6xevlR7nKt2QmvMdpUa
qmhyINRFg5ZKC0yP02LlFOU6mffOmRDeS0PDzTtwpU/YHvxwJI+3tj5u9w9ykjHkLKjsnjtWrkMp
PVqWV+niJYtbJA2rC4SLNAEvuXSSFoQDLWDRCsrmE0iVlF5ITUSSb2yJPLNlEDpbG7rUqAxmBsv7
7/m0E/ryYaI6TV+x0mngoYlNNwdo9YDSnCHZDalftLxJe03pHSaHCUQvoWfZE20CaQBMKBrW0BEg
PHYG8FlgTjnNWxREjBUmVLwzfTZKwIYr/v+zu7Sat/VMiuOKFwzt8fhBU/6dqngUpJ+Dr6KZ4SX8
4u0J9YI9dn68Nnh+L/cAT2pWD1AYjIzVshc7Zx88lBIuYu4nQDjwdM/H64pLDGaTNGcFvsEO//Gv
BEnAtltueFgXYzTJ9GpMTzCtRdNax48d4ldLcybJV7Sje/C1ArPvzrxC2HGaGKkXsPlmXAfLhGtZ
XtdsE9GZuGrvAiK/NNGzmTcOTJ8PZEAKgOLGWws78099fwH7sUMbPu42AbbpT9WUs9riFPwdTyo5
5iv0XB5UavM97UtKy5/JlKAW3xOyk7wyb0K1t6YLKOWmY+52mEaR1Ikwt1YruRR8HACX9BDKEJga
XNaalKQe+wwzhFNxLId3Yq/aQVtCWbRUz1gn1h9hc5XS1+SYW37kViypN7WRI0uEBuRRdfqRtGCo
PNYFby2Dj3lrBqzW3D71vs851dA8Wrzwz7S4tntIUQOcMvAi/LZGCNuh1bqJG1nQ3twOCyA/2Enx
906W7vGkWD0l3y5ybmL+pE0JnujvPUNkMXv7NuiZ9K256LPQks4VJFFfngwMp2c3ORAdzQdSQgqq
WjCKCwOqM733Z6CNH2vDyNTDR2+KcYOGXM5B+UHKtUnzckMrVC8vl4ylVdayD6PEX2BJ3DDd6MJQ
N2+QsZreQbFnDTa3ehm4qYJKKCq4Yg5+1mqb13h2bMdVC9tPoSWnvpbkuz0Kjp9sHk7WrvrAW1HA
+iahL1GwaNvnAi2uRNc63S24UmMyfk5Ci5c3pkgMiHZfOsgexKQg+bd6E0yb/M4/ymYJp3scwdK3
R8gj7ec6ArN9OSHwtmwr1u6HwBPd6ozyEhQxbhP/ZolRm4Tt6TRO8MJjAj/gb/lpGWWawyIK7lB3
IbvRPiWyTLGfqELo/CqTYwZjGR+mBJgHGNcf7TDQP+Egdn3SqTRkBL8FiJTzhaOQnc1NjevQozBs
cLk3Oscgx1ReHpk8K3+Fo6dgvodVRFQzFNSJ0gL/o4Z5Tcgo5xkJMXYx81rBuyzvslKE777iqz9R
/8J10kpU5OKBJ6omKW7DHKTb4eOXRGaTKsdHNdOBk6+31RRhLgLsaqp7nGQzfjikIkMSxn6aIm3X
mNLlEfyF1/NUxGigxRsiAv08Evcf81+Sd9Iju6Z40ui0FiqzZZMNGc3ZHjWsDwerLWpx0yF/rfdk
m+jhxGB2xBr3GI1AUbNLswIP/wIAVecVv8aR2Cs5DJJEJ3O7pgfmOSsOxbLYfFG8JJlE+3ohT+dj
Rn35/8Dum1SvrPBrkgIzXt51VULbW2vZRvuOv97olq5E3jcrI5Tywx6spS1Zni1K8fP+RpzpG4Dl
sw+pCBQeh+YQrmMeF+yuwBUSBeaiAX1veC0hIvT7tOLvFgFk3n4H9Mng8cS7LrlbTyd8XZW88FCE
Fr9gKgDOvW8flycPbP9UrM2ub+fuan6/U4qH4nwR++RcAL/zta2OxOumOIa+mnSjYuUmsaIK7PSu
YD6cPDh+cfc7E7MBHhC+ETf6/8CG4GKcQGZuAsHRd3yfkoCjS3QQVN+87RKWNz5aRH7wYf8u4NSl
sNOW/QvEosJL/6GRMGvog+NirCjDs5r+wYYgrvvY10uGWFibRhsCq9dGMzZqw8rHUuEP5ydI46EA
SUYumKLIRg+jUPrRoyNFl7Em/OAp1AUiSTRWnbaWpweERgAiQK8Xitulj+UHf0YVIVL/qw55w48q
O0kNfLZk3Pr/lL0PpMzIg1VMcDknOg59qfD8YaXbxfCgQQxnuT6cJdpN4ESirMlKPD+ZwCI8c0yR
Z1YnoflGsp7KglMvNk7PvJbsTLTtgSQ0ENXgj/9M7RUtprmZSTLQ50JEMp9C5Ik3rldKq8g5iPe3
WohrTbtTM9EfncrQxUVsY5GN0jlRNXge8f9Q8sgFN3EiPenGEkjntU/a3vkn8nE5gksRW6hAgGGh
ck2yiwEwwgHbksuPMIwcYns/H3CJuYcKkUvs/C/BlQLBGbF4x9mV/2bKczqPZqGdxFwyTzqUkS7S
Un9CrlMQASrIb+kNK07ZUsDfgIHj+UXPYJmddQ+K9JRRwd2SmqAcycpnRbZmh+6LMDl89I6Ukden
8yf9dWPKvO5nKsVkiww5VhSjvR77km8lYopyhUb5tW46Xofi9Hbk1KuzVqoEfcdFssUC7o12RaUH
2Fez0Dqckw4RT7v2LgUVNB3/Ov0cAUXi+6VYPlCpAhonOZE0wpVNzjrUem7VEPYSn/eUeTzxa28D
s5+W4HDs9aAEJWFYL7vbuvKphYuDS1e513OoToAegMXmwiv0xN3XJ5jBxWBMlQZaL6hyKvPPak3c
gz8Q6I+lumwI+5TPrtRPXDb9lO8p1bixAQ5VOCHMUWZSV13glFk7WDYQF3ft8pWB8g5tKplF+k3A
G7iuOqpAayWzdDargHD73M8UvLg2+UfVWHg+Qks+/OkqY5NPPs4OM9hjeZGV/3zKJvGZ9avoEJIb
oC+BXI76OsF3WFOqxc2quCg24GSdEfYZb4BHu4wne2/dEm1n7GvuCo4dGHg43U+LV9vfeGiAIunL
pZjGsUrHQDGwenSIIku4hM3Slgab8Ns29jKkyCu9y+KnQFDr1BiWEYFNrcRwyNecpFgf3jPC/lsG
ZqQmH+h+BJio3tAdC0ot/8RYE5qiMjrfJUCW1ukUTh/9iIyjvsvDKn26JlvQNZodM+gYF9AQ4cAj
HPEeLuGLJhsX7j5ejY3Xi2rDmRxS3dS1XAzghiH/cQ0f16G4hkJcS7SCNaOCWLJWYpMf6scvJADa
AyUj4W8HkZIGP0kKS6lOWGi0DM6CCsbwEv7pwwd5TAwfwXkkCGEsTt1/fu0wEkrRFxsaznD90ykO
vHtgJoilkzFwg/tzmbND65BdWpkJeL0Y6paJ8DcxTKDwdB3RgMuFrFstyo5gwOdbyxAbmhHlUHEq
L8hK2eVGBXQGiV46itYoU9OD1+2SEA0LLEafmHU8+jmaT9ZP6jxTJAy9Nx8KhWkG9kUw0rw3WFuI
2pElrgp81SMqNnMiPBjV0iGCBe+O85XPWR4m3tqrT8AgDz19kSTVWvivNrkQ/k2B2p4SY8WxdbFZ
63cpGBDn5Pw1zD6shkFxB1nl59/LxmjPF4EMrYl5SpvnVd32mjCfXzQplKMI2jLMOBZvVA9fyv8i
+cnk8/07ckFMWjzveIawofnzdwBabvYfHAFYUW2veAL3bK4Q6FSvoU2kIaVWN70OUa0n/r2ArjGC
6UblqE0eSy1l6QvohsQfP5KzFcad1aYdpuxmMHUg2Ox6x30OcFgVmzWXfkRcylTJMRhfeQnzLhCa
sU30Ztx6DNxQPdHJ9kSyHF1ekNRGuUaLAqcPecdIzCtM2uP6i9dTGnJ6w6Zy2/HreIgf9hCmO0hA
8rsUex4zTkuDspTW0UwBiogJgYCoPw4XhJRlrfCUnuhSMsL0rD/ehSZEOJZ7NmE2GYZjvzwzyxi/
GSaYQRVpi7oL5Z9E7vfjSyntSEZHooJDxmQ4ywFfpxnfpTEIdNYUiHWDZvoGETpBNazmfzeGJPCu
ZLhbP6ExEJr2xDllNOESnsztfoA25vVzltIpc/jvo6nZjCQR1MqnZrbmCzz0nDCRjYcLUMM6DZIi
8pJNpRNWNq7iJXbwSNgD7dL1C7IequNY1LIxl+izwW+0mhFSd2k5G3N5ULBhqqKCF0w4RALKWWV7
0UaVXLXRg7BGxkt5/3Bnwj/QIalbjKIj3AHOZQfD0C4UUBNmwX1Lk7+nHLpWKcuno4ULqWd6Mtns
L1PGep+xkeSBc0eniVbUmSAyInlE4bYFxM29iwgWLnya5CqS/bXH0v+TDz89eH0XrLoosnI915hA
gKjZch7NGYIawTKPYnj4WqdyQ5WtF8ZaGq+NjUO/Llh0VNe6zegIhU/6VFl24QTZ/LME8gndrzrC
6hpWWSCf7N0G9J5p5Wq0eYeYfVO76J2rF783t/mIQNNRejekefIYhzV1OgtM7aZLpv8Ik6RKrys1
7JUgNinCICOy2RNJptmkOPDBayMOpVWLXm1u3xl9XxA+tONp4nqAuDmaNCrJ93MGqCJjFU+c0Ej7
jSF6ysiWCLxt0soQGh0qzoTjrnW1aOzcAzUwOgDhOH6oQwoY8hFii9b58+muQstb2c8NAlB71nBP
5iZqm4UQQzGu2xLnnqdP6QcNUIDeM25TZBnbICCyAfK99rvQ3lTvMdeVqorHZ/IC2e3kUl0QgSes
zsysUfThZvn/TaBPrtABYpEnSiDzdbBW8ydm6htcbCqD6r5KOUwvyeqzSVXtSib9bg8b+4ORgjA7
cqrvuOwQ3EFOji/ftXw64Nj4/P61EmiKRs3csaMzPjmGz9alGkBVNapJXe10eimYi2gK+kiwGPvD
WUQ4SidWSlhZhHvC6b4qvguiR25paV7jwX7rpaQ4pFU5kcK4oIkajGYkVGZCQq41sECgIVedTZNv
3BUQY45hDIPTVhCqUKjmCoSajgzhQJYkyz+Cty2lSJiVrIKJpHP66FEpBJhwIcKKdbxZza4JaI8P
1MNY7DViZu+iN/cWx0U5DxYh2SumDFuMN8MppbKKGS1MSbry0Efxjfj4yQS/gfpvhVuUzbp9nVxE
uZZUNhQLWD/nbD8wo+3PBc8ZR7zLr+Q5V6srRlgM5ZXbV8V5mlSL5Xj582rswrrN/+EAYTd85L7u
7oBAY4+s9shaoGvgKQGzS8pMlf/gWkkmgXKIIfY2he3EBUW8KeksIjCXFxJkNeE4lQNCBXlJNfi7
SDxJNfdQQ3xLZpKOy5rvVotk9Q3xYgUWsPESyMxlhenndeGFRD34F+t7Apb7oI+ZONzOZ0HSeJS5
imoKswOY8Mzl6S10jh6STZ4duUnIvd4FL1fyqwFyefqT+TKvD/rTgEAWU8wJoiktyyVuuFXAUdtT
5fIctPJOUgNf5oYWFh5YQHEGvajZadcJs7C2ygV0unKwNtHzV3/VHChQkp5By4f7uVycp4rpEBP9
VcRxPPglpXE0raKyIdecBt3/ZnN3oRCKFt2twoTcrW078TNYyRm5SjCR6s6IKDzRaFsaY5SDzeq4
J2pi45DRTzKcxSCQNNx58swapzutEVyjV2Ag612eKiezkrUZzdH1w9IgJBH6VbnxS7X3/saXMogO
dYgmJYPQ7Dmnrn5WKGLcEBHeBA+as9JvzNV6cb5s+lJztzI7L16afGlWpaA60GbC2TyE0hh9CW28
bniFtHGL5SdxKTx2HcRSSgteZSGQOUYlpzOlaYe9kWxC5Tw5WLopC8PUbmq394s03VxlRI4sIE6w
bkIXjHTVXbMC3Y+a4UfZhY6p06Yp/3b8QBoBgUJhnsbNiaCvD5IrNMpcBgKKDnSGEu0cWPyGI2Ce
GQm4tG2tqE40RuiabSz16hcqN+axFIvQnfP8zo0sMJ7RlBiN3E0S/8QLz4hsAvN5X97SNLMqHgKy
n1k7Ds+tCfGL41PrKnM08afS8werqHz8qd+yWnSBnkcNlZyOJfVm1yqCdBNotz27Zp9VCJWXYHQ8
Mu4WXl3+O+4uAPJMaEMcatL90An/9+PSURLpzytYWF/oMmLZ9Cso04Sms4RWFF5/KdfqWFbkpqZ+
sVqzIgs381b58wWd3fALb4tsk5ScCOAFvblZAGYfxcs1NFdXMEHrUnaFmZGfiOnNWS4VRc/pI1Jb
nZXqemcWLnI4kyYsafTzyq9pWa/8XQGsTPsC3nAgKw0MeIqW2eOGjv7bNqvSztzNVDlxcUl2yKzK
i1RlNdK261I08wXW5SowBafK5X5ajjrREeXxFVD1oz9e1sn0rcIMUTky5/iEd9TAX4agXnbZ5jOH
rSL/g8StxJ8/OxOwYa+1q9vKKA5YtWRpw/aJPm/bn1QaVGKRZt+v/6fyb2+oSgPM0Wnkb/+KPlFi
vCUfoM8xHV3dmQpz+tTsPvO56UGx8nez/NB9LO586fa8O5AX664S2C7Tu9HuWnlDOmyF+EiEpLnf
h4ejnOfxUj5CSEXOAPQqAjeyrPR04FK7dw1tEREA/7/DS8QwL1WepLk0yZIX/KFgVFVPbG4JRpba
7MO1ZOpQYLPVQ1M2f+TCpTrXBZ6bp0HQtyR4kjZ0OgcJUv5QqzP6yaTDmVMdypvdvWcX1ekPrFxr
HFFqIIHuoKfyV3UrmpC6woFCKQdPuLbM2cBkUvH8KV30vJ34GXslroE1roA3TsIZNOWBu1ioX8Hy
QQCrHv/ri54EbctJY4Ut1L57pd+SDk8ALxELd4UYlkBAPO093imghwNNyk1vcBM+C5HgYxmNZGXI
crn+lNDHbEixFU9PPYZOOJl59WHT9WvI6WQgqwD7Tdg3P9wMT5gGxdGKDxMKf4OLez5p1pvNWVkd
dv6iVdjcBIIQl2kqaFO+q8AAmCDFoov6nlpvOsLrptB9fF7DnlE76+EhPTB/bYR3I3o83rVx9dO1
IQjGHJWk25SOzALdZ7wyStbovkZaaAn/JbV8Y/qoN5+9te2Yy/Rihm9I5dOmcEoaHary88K2RmGS
4O8auVt1c3GAlvpXuIqH0oJIjxJ2YkLGi4dJDG28FtKtMe6OBw5jqxLddCIew4VUKKJyyaYEVHAI
6peX9S46qI5Fo1aike35VdOrzhIjSlPyYp5giaMHe10DSZsDClADdnLTjzqvTUrYo7mlA+iwuIwn
NVWajck1HeBIa7Ixa9LXTbA0rO817LzvUy8zZYi57It0cTg7YVZTvHrmBwmS9Hq4O8Lpca8eEsUi
w2IObT06OWi6dFcgpBdYYaeHVGbZsTOBI+Vz/noUhDT1OTurdnLAsYuAn5iyviLGnCdDu//PnloW
ssgCLK7OY9JfjUK7QkOt0E5Rnk+IdOPf07myONxoNH5LnT6hB6G8I5U1Gg2N/WItf6ok57QnFgB+
8y7+d0O3gis/z6evZnqJkA+n0v0oprokfK/hLX2g2EauASrONen+0D2aT7/+liFrk7YzFzKbmEU1
Nnc66VdAAPGIo8Xxb54HXB2dJw1VFii1YXesWyjY2Zu2Hei0J9M/p1lxZycCRT7slzoDt89pJWms
lK9GXbVHFqhgwbW7A523dTJglgvzgTdWfE+kXoxj+KViCxemDQY9k56KfDNyGL6ESw3QsYyVgRTO
Cw1XxklC2ZfJ+NOj28Zq7d7pXnnCthI06RbWWws2a1M460k6vtchJ1af44c3tmuWqH+qPoUJJJiA
HmMVcofDwaRM5Akyvsn7BiRESzBREb00/La2PD1x6BJkX4rI5Kf2v7cPNmraa4Qgesgdp/GHYaYf
8tm4AUXE7Swepd5UUviIQvWJ65NFKywX2TFG34LCy4C4J4+zrgDJvAQ6dFTqCledrz/Su6le5kyi
X2IL3exAZtASAPpKoQ1btByIPZtrjnEn76JmXGioEnKxNMHE11y1S/ObIh95HYb+nOL2YUL93xs7
DgPX4VZuRjfeGEDFdIJd4e2U01rWcMqWdaShAo3mzpSD21fQOQOp++8q+8J5dDZ4IJbCsdpWigQ/
nXvwZFQtrYKnt/U+HY1G3iFS0/2t2/d1sdixbGf0rcs4E10vVientE//2FVvTBzueKzgS5byTHDM
fTrtmKALAUII5Pz8r2TyLmg38sR7hyFcs+TBP9e73X6To6uVJRxV91s02BZW39QXZjvxVzH0jl53
VSk/NwIV80qnwUjdqIRROtUwAZH7tScwwVU5UoWJ41pOFTid4wot5kD+SyxY5bBqpmo5GPseGriB
sGE9vsO1REUpm/8a9QV7ij5NRDWJkPuQoQyD9cfmRtXl1z8rukFyYV8R1HToxdKigseyX4bKCiSm
Yl2VtzB54YzkOwDvtJJ+yxHjOMXJKjzl4SNAXRcGAQ5SmwaQDpfYgnIZmeVIwsivV0qbMfNZqljQ
N+vNnkPQZ+XrFEYXf/GEldxLCl3v/6W81D1nrWO+uCWgxnXrCbQNStGIpoVT7Uwe1ugn6gW10Xn9
5re/Lj0jwgB4EAst8xZm+u7G840yLNWQ5WpcWBXv+qcf9azZ+sw+LeYtrLiIpNcH1hbpU+wu0oEg
chSJAtQTYTdXnDNBpt6jcto8EfltJZQQjhE9VkqYXPDs2Sy+RzxV7zu9gQJwvETLm7XeVPExwmNM
sXXKEWsc421TCF7MZoXazU35UencQ9CJUsRWjaqyBCPec6I1R9k4ZD4G5fSGJEodtZcCIGFWDIer
PVlvkoUO6ZsFbe+LMEBlAAxRrGraRwngalMw4qRZawiOAoNO3Bh40G3szZMXYJbRcUQjG18rKl9V
jMolBoWt/7Mt5PU8Qr+PiShbk6pxe4uBa0CJ7aHx7dYOegNiqZCO21GzKwpCiDEdLD+ab4hGoL7O
3+UriAqyyjoehm1K96j2viZqxH/3UVjDXqlFFR0bpbX1O4eCrqNDvtd5ouMNpsbhS9AkKdLil1Cd
XVb+NgG3k+utbaoMcmpXwZ4gUiAgp+eiqyyGJK7NC8rZU7NPW7ejOMdEi3tOKG/kjGmaCXNZb+AT
sqoUbZ7ImzyDJtrWzdRIeTpi7/mbzAH5jPznQb443CdkTplJ+oSsNrPe4sSq6lOCqwQa1UFRoNIX
DZqt1UFEZlaEAuyYlFeSkBaJZSV5q/EVYqPoJEZrZgjS9PI4pWFlcmt2D58Su/ShEfmXu6k+JMnu
tOGhbNEq3mFcnxKxTXp4lxJ2rbVJaNEuvNYQUpateTX2fqMJ9mdkc+j9+kP7Go3UxdASUq7JZJCw
hAhE+RMXTjD84ef3p2Tm9zEKp1UDAlYErZ7mHUgmvk2CsVIOvCjXLiOsmnWAHUI60FOjQpwTAPrQ
GG5CHXF/90pt5xZfFd4Q//gWrXzSNk8sr0+crRd/xJioddrVE/SajTKIadeeQlGFaQkNNuzgZT09
I5LlX8n468Edfmlk++KHhXMsq22F8qzBpZzyQCfFQuFtW+cNzymdkJMG/2aCNJy5OJVrmRN6VkmB
VHXui14GY2ZhfYki2glPXEdt2zigtPt366S4FWX+2aD4D5rNSfc7N4U/2KB69hzE6uQWxlYLqaxg
/Ivc24VnI1+pN3jMz6k/HkEwByhJ+Ut/IhaCfG4rOt1DUE6RV9rDNdFEEwt5mBmgX1yOAaB4DLV4
UNlP4YR7cX3/TTnIIMwoCn+w/akviX2NUjEp+YGr2KMGPz8YpjbIKBvNIIvs6vNurMkH+h6YVsWM
eX6fw4xGqFqXtd4sYIv6QmvMIKIcvzMzJhM2lqA1FSyvfFA2GEmghbgV4hLxH1mrvOzXW/8NpZ1z
9xUlAi9WbnYXlvMwx+C8W+LDm7AbmQOM+/xsEkoSOcvuiNCODXKAyGfMhIxe77Bnea85pAx5LFf4
/6xGOvgvQyQadx09D9mOMvNNWrObvZDsN+Uv60Y2ffLODf4ZPMg/oATFN2GqkiHfMJaJ7xS2hJSl
hVce6jy9W0EuwmCljwco5/6JRrKk5Qd59HQsWap64JvxWWVXJgsTzbkh7otv+9kNXCW6aTn6mLkF
GJPhvBRwZW0V+48+9uVgJhrocxoHU9Kv/CTEMSUfp4fBc2m6huKb5PUFkgBNqX4Gs/dMGMRdHdI6
7F/ipq2NGHMMX9wtiW8rcyj7/jUNyeXkSqIHFp9uE3FETxBAmGzAIzrUnKywh/egv8urfl5Gx2Il
LJfMtl67rgDPkhMTSPPitGZhJ6b70VVLKrFLIqfFVA0XOeOxA+Am6FYDYIntA/icCNJpvVDTr74w
LIN51GE2VYO2pfpZoaMk5qDfnNWWX61j1Slyk2pKcIiBcop0EHK5EVENDfMAR/OrrwHIC6g9+q+O
N+NSq23NGSvDYsf05yFrPnh4v7D8Tb2NBkHxsyLndmNT8CGWDAaXNtfavB4UNqoBAfsZu/pyCaoX
tQFjqxWgn1z1Pyrzi/WZZwrlnH3HzR3rfq/itDSfO6Q5I8lI2YNvVhyNm/eipZbHYlHVULBtO0Nv
4/bHXahThFhRFvT6YMRNJxRwzG3DGLcVJCE4pP2AHVEaI2Jbx8nj0fxycMyIdxp8Xa2gEPBTXr+Z
FuoVb2L9aslY1OqO79iOOduIWyrJw7YZfrWd2c+dK9V8hy9EXPGoZkf7W1sSx0XODqZMINGGB8Zs
e79gpx9DitLaDL6u8iShk8yWkDQaCD6Cr3jkndCIC+jw3GfscfpAVl83YkRkNrXyOFhYCANT6BYy
z31lLO4S1Ga9AGL+cO1Hp5BQuwmVdNpkjCtkH+0Y0nl7Pxfff50bB7CljyifeI1ggFhEXmDqdyBM
4DzjcXxoytpEwmRgh1z34SZPpBX7S2nHxFGz94SO1sEi9E7z+4mDqLmkut37+GgyJMINkQG58wZB
RtLAgouMkbg6Zg5NAJ45yuk9KTtArt6TYZzeTPT2rqoAGZ/evz15tJCnRa/hX7YOfA7dwAUNGiJp
fIahryNLmOhf9AcFRsWK67MRM0ZtM2JvVSZUkQkK7DIGYRs5kvwsIK2cT0sKyZRxQwtelCqlIuBn
cvcj2QvHRUakHQIeXtvkKdTf/4TsWfPsg+bLbHdULyA+LlMfojRDR786o6lzxajggVycEJXYBQq6
nzb2x6w8hDtN951526aDuAIZYAgCrsO6iTzOrlwYyl8MzhwbEO8FdjWisLLWU1DDowmml8HT1oiJ
pCZ6S0KqE5ovJNB/4gZamtnp0TPd+NZo/iYvgC6vlcWdNL1Qv7sBv+V0pv9bXGODzVQigHSxQzmT
240Hqc4RjkL66PYXj+eTxQUWDO1tJ0q9Ve3WhAf8/Y//kFqlM4Es3XpZyyyz+6XyvzIZ/GaFHYx8
JT9ub5SL/idSW3Ljz4MCzycVJOBDk8z3tJsU/594Eftffzq12ZPhrqrcg41hp/40ULM0Y1otoryp
m+hvAMt034yuIdZm687HrWLZVKmyHgpMkkdWX6mQ5Pwuhp7p2ReYppOBUEYTxOE64+h/MGGGBqC+
MG/ZhiHPdQCCGgz2e3YZE1rpkIpdygkGngJdGM02UuS8UftwZl9IZ6eMwNkSEwisWFOwFAoTGtRA
/ja1Bc/LKqTYJEM7O1pPVEgfA2erTlO6nHaY8ygpi59i1MkvPI6zUu+oEdR4LBbyldnrqde1KzDt
xOKl/dBncOG0M+9OsgW8Qwhr2xuFeskeVRYo0xLlRA8ZO6fq5mgV4hcR1wKl1YY/9aXUfAQpkno0
sf/T81OUbLsHV9q5PJ5jEzVTbMfVW5lcWCGqnwrJWV0xDrmhKrdDI5MOaFSgIWe1z9zcSyI34ygn
W6zDZ/CIvPM/xgSrti5bK1PN9P1uhtwKGafuN4XbNjfESpyP6rXuKYK7S0yVQvFbymhNI4WIaCIM
h4uztEPpJE+NwSl0d4hwimo0R+JuS8jLF02OvI+KYo7SMu8BVHB7ksfZgeZNlmUpSQb0No2lWpGH
Lm75QZEsnvpbj2tx3gNxVv7/a4x+ffxGlxcbrBRNvTTlT0kVQC5OoYjzrVEhgwmheBjFxWory0qf
xVybcSY5PAjkLtzAVakzhU0dSveeHAnnZl4tkQAMFkF5btuPr2czBezVlWqzC6p65Vr59ORAm4qS
S1vW6xi600SFOh/ksSXfujCxwXy48rhCJTMoYQ/Lppfdp3veNEaPzbk5Sf2QhJV/WlhaFeNEIsbr
wZerSNsh7YAe7HJNduS5fYkY2VLhUu1WBgDqB1NqBfZMq4/llYLV4F26K3xJA+beyY9+9JgvAVUp
3CbKjuIT41AE7ukAddJQ6PGo+SqmiWM0bFRf8ACC2b5gm1cenfuGKwrQSKUQqoBwaqka1acf0nRg
AHoyqw+IB7NB8kmjPflGMtraRWIfuYyq7xRRU68LahEeBz4pZ69I6cfWZqOP1OCD1PuipAoy1y88
DtL0/Tnh4lcUR2g4AkR9GgnR0Z3Y7UBynEzRLXWtJiDG2kYycLTZbDeeP7lXN8WzVqRMMoCYPZ63
oqja4cgo/NJQQ36smhmLa9cQ+pSAojkf81h4kTDtSEtmkv9lcubFXTK+M2SElVoD6k07rp9gJn2q
cd1AihNGmrbcODWZkeninhGCArPsTnr3VJeiQ1T7bGbcbA1h0eKzCGvykTh3VqsVBKeKsINKuLBd
NPjFFoAc+553M4lmRnQ5cXjEVgCe9xXLsggpw7Ca8G8ofFs8Hc5agAXhs7vbsdbE5Rswr6wbRzZD
tuu4Ee7TuZGm45p2M/ZgXfznir0Ap9DeL5AQFHjX65XiaGsHmugqjTTgcKLmBHFo4ragRpTjg6gz
qNEo4CjTZ4A5WU1YXmOoTfqeoPkxUv1A9dXcgP74NAYMwukFa9NFbrpZnOttgWDl2A3+JFH608da
+lprId4C9yUgdLpGReZ45ZLtJHiG/5noQwiz/WzpfKQMuBwVl/e/0D1X6/F7eaYXar7PSXcKEj7V
dPxP5RCygBD6MfdDbypUqH4kQ040bF95uyXmmdbRZHazV0hrEGnE3HIazh4LNNgi2zyJmYBlkCMq
UREVLlpO3rakp5A6iU8jAQsdmdM5QFnVuMrWz+yLeccFVy43CjssMws94SUlE4+d+Fg4N0yRGoqF
C8gg2zSJL2E9yrHUUZvQbyyXdMIS9SVXj7ERJ5K7w9tDYqpx+dt5zQiSLuuuEnuWIenwci9e09xx
qjOB0xw3tHESfX09kAupWFOPM9T3VGfeggnMAdU+bwky5HubQbvmud2U24iPDH+p4q/1v7q7Q/eH
OEuCKwbcvjGsqBxu3gnwP5/FjzwBGehHEr03zeKId6ZE1JXNLvXyPsNYOS/NHaOHzpqBwHmf8TNn
n5dbALQRVrofuhV0M8P2MKVnglOhA4n/s6c86T2gWv3PEU6uXsNCKmZZw0na1fmH5WvzRJj/riR4
tQxY96nE7/kSs0inXj+A3kF7ygodeWbfd51u1cHSocXbvXaxq83/hv66TzEnRVAnOyeSKij4/noC
LFRMFIPMgKFgv6dPGWrYcS750ZY9QiEnNAY02HSoSo2pLQDEVasqSD4v1nz2DmxB64KjOANTIOur
ysCizm9Mllwx0HOSRtucfTT8Gs0M70BN56MCC1p/tv7JlFZic99bXe+pzQbKb7YktAPDnaxMxCPb
Yoxqqtt7lKuyQsOYOCZkkaRR2XXZPK6zu/Yh6qTYqrQ7+1iv12p/9EqGSSfT2nQFq+vb4lBtUb2n
jGPSDR6Naz5yBZpWROzjwzJ0pWN9RHm8Xg0wwbWtwdyarj3vp5Z/3Hd9n4Jy0Hh1kEdf0PHTW1u8
J40jGJMM/b6LcMmVnid6vrJ2ALEHrQ8o/+eADYjbL90R9RNgNVw1enHkwpc1b+t8OKOuts5EdqIq
AspEitINHVTfEK9ttPvq97Puy3c3XGR6DgIRdWpUhHM8lXfL3uQRGkyJa+xROrmRI0sYsZkKNUSA
bH+5ft+b2qvu3NVRor5sge2RGcn1YqMlufB0gtOENm/UkVQga3UCIMQsINfC5wPEVfhx/kZtUTr6
FqmnF6G4ycm5r+VgEVv8JxNo0QNB8+pqC+GKWKGMoywk7r/hv1QArDiSm2By5WNPIHkiNfQVN/Dw
49N9Zxfw+qKs5sg2O3JmIkmNeHICCs0dTZiEXdu3R611n6VIXjHX60mvV72DSEvTL2Eg2t+LGzp1
F7CRbiM0BYIZXZ3rFsEbYDLXBiWDIVTuunD7agjFO9q6+OpdbJkoM6pTXdm5Iwyt1DWwxywgXuDU
WIR04homO+LuVTdBchF1WfpctuU8GWU189sUssxlsbOpL6lH2aQA965/YQcklJNqy0UHL0PJLgRT
sLGHdgYqH8yoK8DLqVrVeRB94Yf3ICShJq6PaNOQlrxrSpGlm+AELqcIwn458rcZVqZxGu3LV/wv
tlAcQZbgE//eOQWQwN7dLs1uQG/MPXhqRUF2dwYRS4ULM8y2UXYgQmTsfKKct4Qoq7zKnDsxOFKL
HQzGvuK3HIJcVawL0HB8rL5f41nuslF7nMkVedgSi29TwMh3l/OhK0wq3zfu689JJFcq7NMjvXS+
LQJzpVXxZsdFrBXREmqBIQCv+Fu0Y4YyIwZ18wWbB20GW3Lp/RTO7pbNkF+TzVgz+EZdK41yd2V8
izzmlFg6/FV/Y1JBPYcWir8ea87vFmrk082PZOiodSqSm1yY8Lb57KZxiqpJ002i9iBXzNAiyokZ
KcTachs2v3aGr/r880YLFv27qOxq6a21Fd0P1g8pKIArfGgbr+ZO1wquDsFTwTmdBkVub6+1rfFc
OS/so2hKdYTgQ9xO6eX3y2K8cpZeqzTB/zP3Hu5kU2YnXQUklV3jRPmACkGIp5SEJ9J3nQGu/Gze
QVE0Yg75BeGNAgzzJwmPqafv4JnABpJvtJC5+heaHQALPRS4FSYexEYGZ7NNd2qmmJbMpUYofsCt
nKcTOrRDQXXQ0a56zSI0uMRgBKbWDUR77YCD3RvxatIMSyxZC0ZJNApA1T4wyh8VeZD9mDVc+aaS
TDkvE+2WKt0qsEchKqZd++LnlaYMQ94zCzWtOAz4Dc25wUCqt5Mr3i9iM60Y72SK+4wuIZf8aNT0
6b79jO3qGIKNL+jahF+cqMZLOpR7g8vS8ap9vdOGXXYeTyYtPKxQu6mXduCMYlKTLT3Vsu7CEXKV
YofyOr9IQtNUjb6oeKSrzfbYvvqfPs+0iF1hgxohF8EtmtrbhSxLWZj0TkxGFXFo2Yy682OMncDs
7DAhbB3lFjovH8hPe2f4FXeP+xXTiTsCZmrOI0ubC+RJhMyp9BmgS8I02nGB259dhhEBPeHfQsE8
URgAttPQ5YNFCIpo3kd6/BVXK0I3hOp1J18wIcpnSP3NkHX8gYQ7ecw6G84vQtXXn4ImY2hBitgT
J0qhmTcrYW3aC/KUOQSHAPizsXqcku3260J15ttpdsM6Y2C04Hmg8Dj9YWgnwkdL2HXQh2CIxu+j
hAkXJFA3ZR847LXwVR3rZ3gQIaov3G9eXOeB5S39JaYdUzUMtNHoOmokpGBYTInJXe4GInWIsTuQ
rF42d5CEu2M7HcjUOLBoRhKB7N+R3WIY+qTfddWS8rXCEqtHYxXeSJpsPtPWOclCYUil7EIWdaFZ
RiGyXpP7q9qjerfE14+6D8wDaEuzWFFJYXYrzaEE/mft0RGEsAxuLgkzV22cuNvlSA1KDSUl+xky
wV22sk/GnN+dM6WqFpy0kpGjxAhwBzYlI2wjTA/INwm9+5wsLn6WhDGxgJ1Nc9jcpZRzo9vWEoEs
Eshil2gxaXyZ8W7Jxx7DzUya2yEn9UZfmlv3TlJjaDWs6R6C8zgvHZNCqPeVtcXDn1iwsPcE++Ni
et0ezgPZ5zGrk+Np98vpEB5/WMbLR2VfW7AfNwglMcIe/p/ybZ+chMWl4Hw0hB/BYqq0ZR4Mv8DI
c4WuPrMAIrr0QjQ+Vee9QoAO+Xxq0IA5IPX8/yPSqqsVk0n7byUKCdTzbCgL8+FEgXnb4LxMDOb0
GSQSjRE30D49dijrA1+CGXglA5XROvup6Ow+UfDFJmo4kUxyKUWVmdKbMIakGTxHyplEspnc/FvZ
4Jwi/AukTMW/oXxHC1yEM+aHZM9V4Dsl1md8GZN5ixkkHgQBKsDqPiJTJdhyYHEdzldGKUQ9Dfqb
rlEPT0YI6Xu8l8zBbHgJs686n1J7FgZmHXfMP54h1Hk3WxW24ZGvGICXpbhidIfg1jHsX925t1Vj
TqTv4Ngw4thWeMpeo/2Igt6BubmNYq55xU/bLRFWpm5hlxbWxAIsj5tT/sssufBVVfjE74v+F+Zq
GMQwOVVrx3/4Lv4xCjHdYXT+sYQPh5tCmm03mputbAxq/3inyc6uFEreHr0BqNCejizKBwjBgwjR
CAr5tKU0ZISEjf0t+t7w9URgOH4iNQ7MjXR5zKXKWesRJDipNStT/w0eHRptPjRGnp9F2zY8xXXK
hJ8Tj3VmVI9kH4MQHRU+hmuBw9qDrq6VpNz4PPM1e0Vxe6Gjs2T+ODnzcPE2PiK0ZWWnin1sI24m
LeW83MGThwWlwB0B2UUafK7jj4jKyP4Q6H9PQiGXNf2e1WhnYNUBElvYpN+qkJ974X4RgGIqo+1Q
S5JEHz+km91JMSYqkb5uCOVd0a4HgFUqg+VbRS+K1LD9oT6p0q3ypn3jA/KfsCfKQznbbfnOf07n
idnye9Wzx/D4+lYrTpilXlBenREqbhfRvNqSDXqFRFmvn2r3bskhxYUuc+5AMpvZ273RmCOt6DGw
a1m2dBuJsqH+lbdWXgT8Jqot54K/3zpgH5N6CMbTgNoSwEkqFXt3/dsvVCdnQus/uFaDv329nm7z
QDQDSPVDQLVYGRwYyDqWFJnhc9f77W4hACBGNcMw1JqxbznHZrV+SzwiYqs0Nh47bEo2RtxVGmbj
PBIP0isSI4f3JsYLtkxXmdsdq2DFxxgE3oV3DK3NQx6D4g+QVWgWBpDFtrudn3sL2OsLPxlNK8KY
14ZjunnOb0Vf6lC+VvfEK5p/EojfI6sYdk/BrcOXc0KxIswfx8vtKSmNL5sMdRBaVJ6qF36J6V5j
OE3N9QJJTtUF4vPBb1uIZdmKLIlfRJ+cMNU871AOMIWoiH/w069fdIZXBXpHO+enQcz7DgUW5GX6
ue9JM1QQKws24v6U1A+xvBaVwym2DrsX/eEp2LpzPLaCTChzY1aP4K2QV9eqxzru3t0v4PvEfZsU
URmILk1/+RWs67B5xJ9HQUEl5KagXEtkDMUTY/DXWM4Df6rN9PgS6ogk1/J06ukE6PY0S1PL+Mkd
/E9rJTnvLsIjOd2cb7N4PsUme0/lytzX401GVOcjpjXvD+WO/PcsrmNTE6qUe+Ns2/sUFcNS9JLG
UeOdYv5VZ9/2GSpqCtL4XAn/4bXG00ohE434haFux3AVfBLiNYqMbU3vMcGLU20UXuDqhckGpO6N
QBvnmFasr6zHDKCNoq10mTQ7sRd5/XiP3mFskLl3unF4CGDS2szuOpPkCq9xNvl1U2FZaLEx30hW
gNeNAlZ0FiFldDwt8EWE92XPUCACbWCM9TN7rufzOwDhoQofx+X8l17BNQIx6TcbhkkgOTrA+NUu
fSRqps2Cj/W3i3AsD8urK7suvpd5qdxCJGQ3DFDszrz2B8fVCvKlrLCWyI+z9nofE7eK8ukAf7xL
iCkBGtDQNofIyjDZCaziGP8rL1MdYnYnF5tln5Ndo2EEN13INY/IuJW0XLj9rJpSZc75YnpIaJ+i
odwg3K7vh1NCaowNPbqm6+fR6IffqjYO7armRrYcdipC/f9AF2Fot7tnXvhgBd6Br2jxjhXp4Jgj
bvnmX+vGnbRyeQX2hqQqcBgkVLQCo5KwwbnUs6mwQoEgmbBAVAjU9gidFSAWiOoimqQwWXa5rc2o
OAqqulQNwS9XqHOPeB/6GJpMIUwF1TczEs4+YeJ2HVFOZCikJBCh0DOCk1juhnc4Ah1c6O4KQIGJ
d633Qx6lZsIfMjn9M50QFng8AuRks8MLBbGWsniljxZ+EqaLRvlFkUbUImTPyorBzCm9O6UsCQVi
fbjN5+YWiG34kxZ/4Mz+oZiheHtsDFM54IrZD1Y7niMSDbm4nKf/ko05TBm7Dbn366ADT5cnG5Q1
GEW0nBiaI34WL2k9QCffM4xIBoYZ+tPY6B32UodQoTpRJpP1TiO3y5j/GcmIWTcnA4ihOpGnzDsq
Nca5D2pZRFQzXLMJ35flNXamr4uipcuzvckyy8wYjJhfHYgqFsPoQ2qJNrDzQ7dCf82hMU9naptq
a9Sn1T55rI+5Gb16k2BZ3poQ13IbAukEYejSZjxCBo9sTd+gSPoS0W/LReecEG1vg4t4FVBDLW7w
omryDlx3nXxOt6kXjt+RV6+I63nnaz6aFI0D628//+rdDkik2GijW4/hENNbEkQZL+nuf85CMu0p
3Ln0ImJbsswIYlRgfmdtY3Hc86152eGFhia1qs+DAGqNxELMeEAAKsy+vqQTV7+11KSYye2KNJ/J
/A6Coj1XqiZtJ5gIB/bnCn9nOO7AzM4NnMij2hQJPd9mhHpHhekMnwOknLx6omldh69xMc2I2dkm
8ljj6NTpPPWmTUoYeeDpQRJcv/A0Km+jLdl1CymeISCu5ymGLtN53TU/M0x7hYrBkXAl6xkH00V0
JtKKjCxLCgfxCNmiYjpEKkOHYas5oCmt2BNIrWUyOmTL4RCEv2Com241B6YfmTtGxhDxvnGODIV0
KN5XB628CO+JKnPWDvImbZIDKoXRhJcbaA0e84pCdOeYic4vN5i+rLLuPcjcKUUhYCRoib++SUr0
S9Eh6WdKcu3kIy8GewQ8jg/4I1OBM5LsO/hRMKv2ctph8h4j87/ypvirR+wfrAmnhSAvGR6AwibE
Zd0KV7ENQey62LdCIve8sD5y28CnIj+yrkBDXf8E9a/Lcr4L+xHRVUQZiUH6j5CTMd4Ni8SDQquV
5l+/6Haiitet6IpQGIs3LemLYX9XGHSRcRvuRMITbxDVcfL8C0TVUk8Y8U9xDS2TP6v3vZi67fKU
MKwYEOX7CMmpmbvbrUqQt7JaYAQKGyfIsI1yItciVwKqTDwmmZv6JMfnJ1/MBg3qwTcpr3cZbczC
dMh9uwVsjB1FUINaMY0lDmO1fggbwEVHyx8lqPe0xCe1s5uvcfZefQ2/+G2Pl9rvt83gSChmDtjo
R/NUuD7UH5vg7KkzW4v7D/LJHz94aDAZV9hjgds5PKFLjyF00eFBPy8DcQqrfl4m+qQcXcmb6Vlx
71Xab4WduAP6HBJbjItiWopQ9NQtzQ8RDlbvGqg2Cz+fpFBQMiFlqt//wAzeymhpCSfgtEIcu+CC
lMjcCS/iDJbBarFnrp31YBhvUPnSWdP96E0WAQEVX6PgknriAnDmRB7JCbxHrR/toLz5SXPkWM9O
trNjgWJ/etw01Xq97mj8aenOYBD7AT0fEDk0P0wMzeiaBVNFVTtB4ylLhFz/oQYC+TlQwoxotrak
TrzI/6bktjNVuP593E84fv5Jj5H6LVtkKzl8UdMRit6o1DzlCJ4eAdvgGUCnBuT7fRgIaeNT+/hd
KEywEajGpasF1h1nb4YjeO17lE5d60vHehpzhOTmUGBjM9lBvzxfc6RFCYBkXpPBJNVxRXlpi8Aa
zqT0uPa5pwewsMbQbxTBOWMb+ETeBM/+nllJYzgPVo7XtwAwEUFQ1e9lHpLubWYOi+ibe+ezmSlx
Wc86TCl4BEoqpjX/HyXHR9xpL/ZZHUdU7uXpRlYkzB2VwRl0rO4FhNs7VC/IqHUwpDuX34GUEnlX
znNfNVYjGVfvoX6Pwat8lQAYuMWBpMSGW02kxgiKhzBgnugza0gfJ0m141g4vuO5RUPnEaiEZJQf
8JhDr/xbdlJ5+FsxEkeQLqfirwSAsI4IB1qRNO9ykKR959WG0zIqrycDRRR2BXnL9TfepTeNWDM5
Iy5it74G3URdUhNdILnTuvsxCqT4u4OttuEzQqE8f6IAIfjOGgOAqHRkPY696J0OCYOsphaGZxk3
A3qn6ce+zNCbhQ6WcmoLTaanv8HISWrMYP957IN6T2KxEg5vZIwJ1BuccPWpdNFLkP1IXhmNwzQ1
lkTQNWSJyghqtp5Q+fz0d/cmRaW5gom5xOwjN7IFPtnMbMSf4e2dpLkWaWokYpWtNGVdmLI1HDJJ
shcCN5a7F5bBlsK9DAJNj5qyDHj59lg3uoz/Zxo1VwB+2nhiqoJcGNsoSQDx3sISEiy808NnYX+M
NDaWniujkNn7IuR+Yvz/5fdVIxcvR0wFHo2WmcxZPybE1Zsv3WtZhtJhhud3ZOAMrKVKTYbvfJno
LEhKkilPIoQwhCjVHV4ANs+B7Mo10TwTgJ6RVPyANSSQh/9+i0HEgwzMI5vJ+cHPW/2izMH5FF4o
wHZh9A18eiiNLa0Z2TbvnGbQDOMDJfeKinyNU7hofhOEdUSBzBzSVhKKYMwRnUrOOHstuBAcPDuy
ATyCdrM3GbJ2v7LDEL998cxuCNMW3sTO8D6RWRgxL4gG/0cR//iDyr6SasOZ77wYtjq/sWL4+FLj
31aBQ2xnZtPD/lnyx/p+UpkTozs9G3/vO5eEovEJWAVrdAuzxWWqPMZZTz4eLQbqoz3lCI/RfxUj
lvmyMrTYQu87SfOzL6hT+iDZFQTdZprhPiMj2IsMfK7sCepPaZbzIluTcbBjMRKK2P5Sz6cegYbo
XFuLHLO853Gh732qujXupB4EnLQH2oYMHMMbfrArvi7/RSYl+S/RkmQdEazBFtM0kPzM8bVqRO6G
wRCw75DDjnO6jAc6srT0w6poJs56uvgAEs5Iv7L2Fm46uWYSdhA2WGdPNBOKt8IN/RD9pxIbDLhW
3AMMCYmQcfmSl+mEfwdEJE4eTkPRl/GRC7NaqxSErdE/XnGfVemuhwZEdjYGopxOqbAvykd2UAJH
WS2zzMfMg2oQSV4neqq1fm+eq4hLFXQoaH/cpFXJBn2Cogvlw7/zzwUqiYbASEkkSh/Jni1ssQ+T
JchNRacwkjrdkdAxwtzhd8OFhGhzxwC4wHL0uiUMm4vQUUc2lo8kY02B1eNQRg7jTG3RvFXeHp4F
j6HoNzaPCvZtyREXDvF+BRMezZ1x2XgyGXNNDuZDmHgSJ44WUXA9jE3JG7iQkMt8QFUElKPRFcCE
+ZRkUq30g8I7Z9f5EFCJ9LcJjwAj7a30KOqL26QEV59uGiVxgtjSP/p7nKwFxoynWgYp33bRVRnr
YMb6yI8eE42YQVFpE4JRjUXOPBOiLQHvdSKRcQoJZncE/kZci0u+ArVc+Ai1ilvb6nVT2604QoLj
D5YZHWkHX7lrIh7LbdWfJq/EWuYygHfu14VK53S/hlSc6WRtWx5F69wBe/95Xu1nYUojkRwtqHjs
43VsexLAiuEIGVMETLcOQ0swFO9FA5MPRj7NNU2hng8Ysx02JIvmQHzghxMw7NUtsFpdQdKUEzj5
sCXGF6mEuuaJHb1PYqBvapodQiTO2jJPJY41r8WElpoALwm+eL5hQ4TuifNoLI/qKP553zTQM/oj
h3mTUXRgMf/Yl3PCgvP/iX65WCtxuCSG5Mu/orJLI9i7SDeIm5CWozOWh0Rh72VaqzluBAVWz+My
oUuNjzMjWqCHYWxON2pZqgocKoJ7IcsqYIKTpSjHUqA7mmt7Uzw7LCvMuXsU6ylESw79JHx2nJ4o
lCDcbUfGCr5DaJ0q3m+uXkk9F3B8hwJM8gYqBgA7KHIn8Qb5+d2TfZpqUFtWtrHWxBl22zlwPrSA
C+wFtnGedtd0RjQIabTx2REAzVc2CYTJlJ1fsYEG9qMZYghyWUszKrLgR/UAY5eRn7jHgcuNGc/j
AtEyul85GOb4u90x+bMZ3JH+gexcGFssPyZcwYFhoRM4YEHH6uOI4bYOulYohnnCb1eM6LZY/T81
yytogmfqlCBT2VS3j+ALqI6HCUAlacmTO/9ic4eSdcQCX2pp9moXCOhQEiLCM5Ta5TQFgBeeeKOY
tOvmURP6l1GODyllOzWyfmfwCibChgtn4sO6NvtQJwDIjg4yv5SyUYigRJiPjCToRhSF8am1bb/+
B8oc2+MdsqFFEevPG0cxXAMDELrTIxt/Wua493khj2xR3g7zxKJulwSrjzb5IDyFXz4qSKarkaq1
ktIP/8BXB0+eMlqAeRjvWGXBmAIwKJigfUV4nxGaxgUpxelpuzt/1oYrJbk3VtUl78dEda3S36TT
dnGFrbcxmuQbMi0LzftXtPbwHtJ6A1pCYgVrKWNnNp2Tjep5fIWV3tjH1CA6dIwDDwcMa6u6AJG9
aB0DA2PYWx37w8LBAtTHUXGYCsaRzTlxukRPDRGc8jcv81cDL7aDCUizL8/+oiXI8Gu1DPAz91Xo
aomZty1mADG274iTsQFEIi2YZIh3E7EIB5sl7OVUMRhfdGFyvlY0RzWF78nhvvg36e91KoTgW92E
Qp4cbh+sLIlRGl14U8qx2BBjfd/DubebYvp+CWiG/l/YHfw7bQAptx1oo01PMERbjYcCkDHrqNkX
dJmYBr8PUNPIhQSHxcrapE4hCRjmjT2FO2wrPEh15zyEa9PikVOTo7tuKfNJomIoy1hreb0aNCfP
AswodCBwaH5Q30jsDVU2BIGYn41ldj+jmjQQQAsKHIXjc3ZcZsI7k94hg/BH60vHaa7dz0ufXTcJ
e3nELxAOObS8dK1HQfUzK7ptwDsOPCi08YGCfEWmJxCEg/YhCeTkzGDFghc0NRrjNNFq2QfOEOl9
tCojkDkEAilw8fUN36pPnPKsIQQATIzcN43ngysqrSWb05A5LDVGc+ZOxEjlyrWOh6RLHLfpUMdt
kle6RN3FLzMerAWmJHy53aXNNXq2T+M2kkH9rkLMEYWRWLX7XkCxLLA5TAQUUApMTjiLtwFhgNTj
1ZOzvkvDv77QQNAAQHhx9jVyTKC3Gd4cOFqOHSJaivXb3VPdLwca+Rw03Yi6iTZyK75hvc6QTbN/
BRzwvPAiwjLgRNZLhZK0CGoH2rihmMEmSN5YOrx2qVcvCRdZfph7QBjf74RBOXlMDh1YISWeSkSa
KT/bGiYD1T3PMpN2L88bjARfqlWUdKCisfTfdmnIW2DZteWv/Pjxc9ExB/Th3iiJ3r47JkBhySFi
QzqUvDdz5C3adL2rMHqwo+YKnSn1kh26QxKmFeDxLdgcAXCRLxP9O5alBMIzbCHVpm1tBdCexzoi
yl1BU+s9lbVy54AKpHJGepYYGnvB1BmdUJg3IXrvXaj+faTGrwskrOenpfNgDJGwEKulrAscoPBy
a6DPKOOXKdDGPoSANunsAU1uEFBVWKHUOQRHSlhwvhMXRSY+ttnMVzgHhktnno6JAWnpjpchIu+G
d9i9VzDML9OM7uvxokKRT6SuwIA46Q1hfns4Jqhd0mSxS+FGuxDZiOWEPfSZVnVM+/IVr42V95bB
HqezfzZndZO67DJuHOS93a3hSHUQExmiRXtmiGIxkvyriJGGxOktIGs8dwFMDodR3KHgE7Km7ukU
JwheSo+eeOwfbbFnEF7+L1yRBsWMlwwVFf5j4VmYzrN/1x28wI0zU5pGh7ib7e03qYaoz4uo7oHa
hc9JhjaHjVCiCB4l9ca8OJl+/k5wFVRIW3gR35/wIfPOhczWItsrqzOpgKEl36O+b17ex9m8SXHp
zmR+Eoepi2c5/jRKC+F5TOnh95dSRKQ0ZZ2js1fq8vGO2SAmcdtKkoj03xtPJqPWWte5wESL8+LN
dL94GGr3mAeyNmgF3TktD1FD7tsj6y8zznTGcr3dPsr9MqgkLBpJiiVk1bClbVTkq1EWXF1MGJvi
cj1V9RlqxuYcoNsK1MkCBOE9Eg06sPjsfVTum5NXlSgz42wt5L5FISNJ2mroFKjry+U/6GXb55LC
lEAX2J8uDAQyMivVgX3kPZveSWdRa41Bzeq6oKdHonAcjkuX4tvIgb3g2ZJ6S0jwtqtTD6BkpZgC
AN+sxxEEs14CHNCSsYqvdlzJo5NlrzWdPHSQEQrpKwbnerDkdDWBp5u4K9O0tytT8/NGPjtLO9YF
HB0BFlTII3nCpdfBOhUO4gcnWz/y+Uy5tin2jNizTL/ncvzBbi8NBVZ83KLWrNgsNNpUtAmq6h5T
utJDgprgDM+Ij/LbEomU8XMqLdMGGwHEzPt/U1gW0ml+c9emtatMvVj6avW282FXTjGQJNqsfGrX
OrH0sCqcdRVVVm4HNhGKnDXAErPXo2Rts/jcQifs33A8wh3I9HFPJ7g3+rGOvfchTKYkMjSu/kJx
k8i3nRWx1IZk5yNFX8+NiOsbJ1eEvAyJ6KKenRWWtYoggzysAlFi39O6DK/r6cXK45FPJ0CZ2+tf
E0wEgMlGPZzgse82KnopuG8i42JC3zmhzsRQ9z+CSpkNQKAFG7cCg5qe7jfi+6xaQ1icXijbf11H
g3O5Fmzq4xr0P+fQVFBd5ga31ZNNgXCGZvTILt+hOxVyBwLRrrOfKXk1xJsP/wiAK7epUjCeW3X1
E67DdKQOU2VXz+qWxxqux0IE+EdwNdzw+SdhgP+mjTrVdrU115JHA5B0v9xwjrbZ6j06ZC+XjUtw
O3/+5LEbUhaHqYnLhGOJ/ij6J6aS25eZCH41t16QklIyAQPFSo1kD585ALT+Xrtx4jOj5+V6jUVt
Ly7zruAS0s1AxNr+duQwXVPqWj0k9X+uhskATeOueaqES+33J2ir8v1dDjXEDGGciQYM/wIrQ56m
SEwtOfLfbrUEBu25BeTZAZ9W714XNAjfYIlWumYxTKtqPuLN44p2Dl2xC0cAq7cy0awm4P6/YBjt
pz9VXVGeB+XGL7pe+0w/F7mZhJco0MMzNqT3yEDpO0v3BWsuO7A565PuNXYEp+89cKRBC0XabuQX
cUVq5aI/vY6Xaol3YUJraUFuqvlF7x7kSxI5IAXYttvHD6T5YG3PNsqgFRwSWaOMCoj9KPQAdCtU
/dQJuj2lRFPg7ivT+Pw+AOLoStA3KHLapbI3ObA5cn7vCAa0xg1H8WpAcvPpJBdwydg+jT/+8BlE
ozrQYLTxVlXU0HvJYG0B6P/apWzES/oLS1JDEMzZxIwSfii6lVbII77enlwuld9qef3rLxnuLVMe
BXHiVmeWu0HKREEzURUugGLbjONr660zH4drNGCdKwbV0fd3/1jy+hssKsVRiFlaclxaDlokuP/U
lMweR4SYaBqfq/iPHZIjNMpoHAznQl/grrtQxFDPiShHDYpQDDYHxkWOfPkCwXyjx9qhT6we6QR8
MM/axqb4yg5f67nk51sJHNszeMjI0WQsFhgNe08ekkqNKhbOdk12hj/vrKJEr0Nvx/c7/Av4ysBL
UJKTvxI2XvNBCzZsbXRUCtC6HtJq0c0jSy8kKuEhU0EjmzjsDhK1P7SEz6LEzBGHrbIfxqblZotU
cy7MnaxIkozDGmVWBA0+7sQ74Vecf1WPuy6uxWEAaqUs5gNveMimYypj1ht2bKfrdK3+F2JCbPMK
iB77bro7paO1WV9jidc8CYa0i/VpsJeP96IU0rtLGG/Q48MuNsd8q0dwl3jFVmHjGHw7bgd6bb4C
1Z0m7xhadXVkwUF0UwYw3BxNudhbimieE/Svu+JpY2P/CqY1KoSrB3nUOqXMiJ3TLzhjK3sYcmdb
tgKQUSVfqQGZ5CGIu5tJNUV92CdBG8HxWEtNElAmLRkZNDNFmmhQecDAh7aYwsPENZ/adJHbvXof
papzKAydkUt4Sfx2V3MQk4mcXeH/arWlpd+NAt4E/65Jh48/zPdoUNxLVJWonpx255TBdQ48Jc0B
2oYUOfqIzv7O2D6o2BEX54rFnT///9t4WhCB8s3EkA6Fn0U/wk9A8rfscaPWK0a+cl5hCCIUgOAt
+OIORt6pOngP/K6SuUv98PRLw+Lp7vHtnqcklkwjvIXnrLGRDuMVJrzJXR+Jl1BGXED//SAREBPR
j/VblVM7x8dHs8hUoAp4jfQecy5zUXyLJi2+wW6dq98YqJIk+NiDm+lt8Ezt5WnqkUsOTj94b+Ek
jTtHZVI842VvKZdIPZi9oXadNPkmgkRdCA9xGTV7QGNtuNtqlsz0Am+Ft6dhZsMS+mJorl7ZVYmn
Hykbh4s2CgCdzzbHw+YEJaPGN1yffwiJ/SW3yfKQmdbk3PJ3DVl1+XdygQei3K2P2TdhoJwL62X4
N5SaFEHQluX2YD5tel9m0mm3/1xcQd8ECyUCNPRMeP9CqWvRYcaDUCZmLS1kgT3KZl6L/1Bam1c0
Ft8J/m7gmAfYJl/P+Icb7ppup2lzVvgjhU/Bhhkv0OYEHNTHoo1kT059GSOCQJAeXbbqhEZC3tsN
00C8dLJTf9TGrO5/4YaaXRrnvmkpZH2KMYOY0jkZ9GKX1dRwGyY4noAf1tVnYXfAsW/A621IVmPo
up0k+1NeDCXZxEcRm1aFl3kILTj0iBl+aPLHwPUD2ZHNLGdrjagrl1qAxkbHrx5eszcfFtOSI5gl
nOxNOcP6n5aXqIO5p2q2rNtm5ZUg2NfDQFAXKTMyz4DsPcPSW7tfmADogCQZgkphQaYNIpg0Bx/y
S2SObwmG6x3/AJAXpaZRwCTD76y9OXMUw17KuiII2C+3xxmi3qeadw0wbRMjJ7mBsSZarRYOZlP9
nKf56UnzCkpxJ3eUHCyHLelr9BNPPeAZUQW/eD0Rj9ulwlgUkZkcMC8hZIzKNZyVkltlwIPkbFmS
cGpTCc18L18KUfxgX/Pof0CVoL+tND22I2tyokU8sWichAnwGHuiMpto8gKYrZXPz5hFmQ11YV9R
Bqtyp8j8K1xkpxNSRjkfoAghuQPttIZxGrFjFrvPpJWbHNpygud9h2r//ujyFxeK7TbEp41hlnk6
KWPlpEw5ph5hri+SfZ6yNTwcdLPxOtWaGrdrYbYftQBS0Vu6u6ozNv4krThdHIzfzZuYowpyHcN1
+Tf2Jj0JTghSQ3p6yhpGEGr2DjCO5WnU0FVQXXkwzKpvd9uunqZ8AaOnfGPBGiafNsvnFJ4xwLhd
tuG7MD8/8WRV8TAKT/K8vbrHHrbkjvn8kkVtxd3SBEpf+n/L6ZurH/XDb3jCRR7nQ2fAOlxzjYAQ
0n2MuUspg3BHCJPEWaQhZNNWtlWJtpzmPO34UUlcFEADV1Urx4W5mtfryeEfdHWbaziesWKWMjhY
0qPeDDJNM7t8/94u8/Mx2/tE7o47r/MbPvFcSWCynwUlCQed9ZLA0OiA4QivQKTOcCVycB2gyhX4
PdLJmleS4pw8lCUN1oXEJnnZ0WNQt/txaUMb5LfkrrT7aoe+cnfq6Tt8OdNEejYLLjzTh7HQxMAQ
V1m/hwrqbnLhoOCbKmTAUx+Qtww49QJgZRS0ApMG43X4++xj5Lc7pfUe7fgDJF6/3vGa0dboFaKL
Q3XJpEGNp3VBvVp+RNb3rDpgdvQSR7KzOK0fvP4VhvHIaa9xX79S6kbsS7UkPIaohesE7L2Z4Xm9
DIl7pkQ6k1tqDH2koSpSxnjZ3CXT4FWQqhwxxb964towJLaHvH58AbQ79mdZggnYJxocuRvmDWME
YNEnyQ4bFyYAtXYGzJQzdBtpfPN9NWwjb0acEvanjngeaVQy67AhZ4hyNDTVDLqVDz5UxUf5wuA5
9PvVCMt3Zub7FRBf2WB8u3a2EbWeO9/+wrCRAtPrJ9BAAMatYr4mUYM1AnMsHM0iYYo709u21nUX
j6lzKDZ0wGVYqdCLfmSavy4IHyFrH0irNxLUiSmySwotVjrZqJbNvyADmNeIOxOsBuiAncxLXcKF
50RLNbK2knFtUUl6xG1PTFT5XWgqocFV/oZ4plvaLaiewqaINCP9vM7clL9zDxzfjCiZ07yVpOZI
kWwTwNExrRs8VEYP+AN/NDfROL5ZtTEOFKs+6BdjCrSZhyfmJV8XBuGUdrEbF3NBvBM8nefQaK6P
6CP9pPYA7J2SONzUhzdH7/gGtuu60yybRjY24ol/fUAm7zeCGBv94IkdA0ZXWV7SiEnq2f6johue
4ja9ADYbWG2CRdm/WJHk3NS2ConEZWjdA86QPxaC3WUuyQPOjlzlzPOyLd3rD5+ksyyWKWusAXky
8FXvRODyWUjrmQAjZNho02K2kXOcN1JWvvssvplyFTU/xfou1s53aTG889wQNMWzySJZj+J8+/Mb
kTt/A+VMxf94EVkMXEL4hj0aRdQIbU9fgGjgsA50a6hnHetkNGCWt5jYOFUMQpc5dxSckWbPy3xo
8hZFo1n/SMLxOK78v0so4gFJBd51LiJ4JeDkHUs28kDLfZPJNZOSyVXz5ChkGS31fFlLP3bHdj+Q
rMmoBQl83s3EPRohHe9qoQ2F37v35wb1vCc5TPGfXex+RsjDHD7TT152smWXg0+CvoJ5GAJoHSBc
1O5d3k73EmBvkxawht761B7/MTtV5XoODZ8VrUTX7W4zn0yUMmGt1F/buhdbhZB/xiwb9N35BqFJ
IgjwsFyrJDv1bx5oo6ai9qaCm/+55zv/XkLrL34f1oMPwth9fBfxVBHpXN/FRWiHlulxI6zq6/c6
3AYwcasCsb2xuCkp9j5EIs58L/qFCiSQ5+PDzHIRYSTkzMRsFs24+Gm9pfG0aNdpg1xfNDPvz4KR
mhQa/ojQRQ/gerVQOB+yOfAuYp81P2wsSJOKKkc6QHnsLkERGtblaG1n81DkN9yJvTYmQ+flwzHK
Lql3+ZVyLxcFsldLgMDq0hMFvm11p0pDiO/SSw/EX72dnr+VJbBQKEB/yV2vhCWoGnon32l1r2Vh
Hf6EjNFZbJ/daF7iDMpa2EuksAV0UOU9ReZqRu+gF7eF9Py0mEcRZ9hdrwrlObGWbNF0wDDVl0fs
WDilRTqXlBmABJk/1CUpw25XGhJa8f/zh1VSUpycNaqeSViVF77XL9RXeYA/iFptHD/LdcEksAxP
4OqjOJ87/wgAPtw8MIKCYdoyXzV5wlKeTJHLQfXEivQEzqeODIlS/Q7qhJvyuoY5UPi1jPw2mLk9
MyTQPSh2bRQ8kVCaXvQmEKdYUVw7BzR6R0pWqiE3d95LcOuJpC11EgpfAfaBZqsQAmhD6sDXGXpG
0v1wSj32rBjE8bYNYH9vzBhWFifPhFtQ7hmFlZzbI4U1T9MYYuZtRqzhMKaG0SsYrSAF3fSNDvUp
YpmPXecFqtukMUdAFPUvcZNXmjcPFiKKEb3Ph5ySE2Ym2BiwrPZk5P+j5nGbGHpwMUBnWionVm1Q
vUIBRTc53h+nGRvrbnPB/gUOGMj46+u0v7v/kbmeqigh4WrDhPe31xsdsBGoplenM6Bz69My28IN
mxtvyQv6i6odYqmbg4onYe9fPM9FZeVPP9/8BXE9CrBhYgfw/k45U9Zq4CYp0SEiYGtuQiCdzZY6
7kBRMvOraOx3ylfMFUQ+xCR0UHRRAHTh/65YKTveCjh970aaYpcog3hveeCyMfN+afu0GROZdm92
VnFU7V+Egc1oWgYy6wSfuxZ/ex/BM8n94ULjexx7oQw0tbdHVD8YIrvH3+SnGterA8OMaK2uIfGS
bu9Q3iaVVVt8vRYDORPHGiSCw3vLrz1QRrW/3GbyZ5h7on7Twelm3VsZPHK6kq9A4+6weOpYsbyd
wt/0mfZ3NlU1Obiweo+5hFhVZ0XnfxcS/c6z+ZuVoucHV1cYITOcf0ZWtSIuFc9qizLqGj5C5uL1
Dv7bvQeA++cXEdIhGuc1vXa2He2lS5RK77/YOLXmIPDq8Ypu4AilQfZBdkZocRnqfk9rirpT4CfP
B5e956gIa5kx9sxlUKWnQpD3G3mV1ddNAvp+fqGXdly+7+e4gmoaX4fiR1895A+CyqJmGqVYhKwq
hUyPKq3EijNe4m6YINQk2aYV8fix4il6ZT0Z2WGUWUYCohV34nAOcZ3DlyY6D978AKAD8Ly4JFlA
BLYkIuO8XulH2cO4lM9YtWtiko+NCJnAgnxB86MVSZgLqbrZueuas46+8ia+1i+BxjbLrbgmHz/7
6+XNIqthg1mafBgAFWwKVgDdhMjj2+r1qUgs1oBHlb92vtWYWhNQiKunSFz+XdkYkSbm2Z8ApoVA
W9o+bp+1IrdJgAx+UVp/JYzcpissCUUTn9QRdUetIPzXW5nqdYevorZ4nhzyg91GEnSsz6ctgQVL
NF4pkpgskw93yiisuSL2hF+TQjtDG69Q4Z53FzE27e5EwwQ+TOIBC2sBSSbSViHrahknA9AP55IW
PMMzftVCbAadMnpbTD5oCkIV3x8OcQSVQ81Ch1dI8TTxdc3Lz2CAOpANFcVfZVWVA9TFb4jOChrD
iBDZlhel1VEwXUlOE9RDOW4rMR/e6cnf1NMM+mh2X994X/tug1YAD3XPAYnUNxtCZa7OjK6rEH2I
EBY+W3dRbPjkO552oOO6SCY3Wix/mHanCSiR91aUnlZu7Rxu6Ly4gTEH28dTpYdK3ZG68WJKRT1U
0URRCY6+EudERzZ7zH60Hcj3tx/yWrl8wFQsDHkyUn6izVn9oR52OcPAB3L/QdagATUhXxcbe+YL
23j55r0epnTakKKUboRunAxEa350vQbi/FVpgBdM+T7oErWI1Y0ntea4TmJAXGOA+7TxgC8zdrsX
VKXiujkxttnS7pfrXfOkLI5qiK8rDt2FFSxWelr5gv98yK1mgvBpgA1zTiAfQp4SdoWNNdijhqXn
y3rsYwa0WuHIb6mtOZ1p4b+NqOBqGXMns5Fg5pgQEeMbSpZAilfJmrs5XgnJsmh3wupRiFSzJqZk
ioCnxmdxPri472P0Xz5rFMIwFJhdVHT5IZm5/nn35Wc2p5raovtTyVjLIpS6A4+h8JoEpZYOEjqL
AvLO5bWCbDJ79vGUIu++vmhdYDSfrSsF9gnb5ZtaBk8uffJRAg2AReAsss5QrEr5fgUOk0MPjxqH
lwJ7SkA0Hq7MJzcqeVnbEgSv7yS7Qbbcl2XGgY9maV/EQJOU9w9Rt8bU/1xhOCQ4UnLhNSEHlCqs
2OjYCjCaLivbp+bJaGx6O9etsInDcBuvmzQ3OjkEHb+fseLSzBvhJwk0TdRLw9k9pPaOtNPj0SBR
iUlLQUCce0eumAyD27A2n+JIpp3TzgraC4PD7gE6cxFORIHXbY1lGchJXdXa2TldrOP2qC6Z77d+
qDy6Tur4cXfKVv+qC8/NxxU16w9G7Fe/xAwqrN+uIW9kXddvpozJW3oaKZwW/gJ2Mf/L5xmu8zgt
ka0A+XsyIcI3H3/lviOevzT0P4ViwAdOxRcJguWqyh9f3Oq2VO3EbKwfiIrLOYB0jlAj8ZhVCeUT
E4XXjxtGKrtvd/JJc/RiJttWwrncyiLRm0g7bcvxlA+06NEZd8YjKK/xmF7GykURG9a/wRZDYyzs
3DJuUvwiqAfhFh2lnuWFDI+Xp3vqMoyo77Vz/TOFQFcGxD5bYKtgEPV+sFCUlT25n5Go3PK6SmxJ
Wol71NzeO+tfdn2D/ERTXX7U5HkoIHUmn256jYdz7NEW87X68DimK1bLRbjeq/ht1GI5Xz1Dba6S
bNIo1gfnzkdGb7/ZSgqRJk1OzPDnxDCuDd4kcZLs9EEPwicAnjcnRpPxtKLrGfTCJHEEWCi+UL+t
C9Bc//xnJXDYOyFCmk+50KKngjEfOYewWMCl4U/2LvFai6+yAAX+myoz9zyAqlqXYkF0moQWnila
tyqXAJVgWh2VZ5SLqvmILtJrSM9z2HRRV8sjXaesAB+mvTMnw8RnXaZNjlFYlGs2wcxO/lMToOgB
ZwjO4C4uZWcbupim1BCDEGyWRI0xq/kJAs6D/r6kfei+qI5oc08G4fpCKIm7RWhAC7S35SHWnYDb
TnLs28Q5XpoQYJP9tOqGzb7ozek2J5iW2Bf4oxFCWAV5CnsD3Gcp7+euMiVnMkjG8o7UTbSc+ldd
Dlwtp8CntpCXmM2B58DBjLZgE55kd9oQD7JjwfDRH9msHdw9tFk4J9/0xpXk17cJQMcVoV6ZRbHm
5y+rVD/GGzvlI1/ub5AEPTNJ1ipAgo7q6Bk1F8q9HUMdGzWsblQJHn2bFzJ3TM75mWDt4hsRF/YL
d+4uu5s+ukHo8hvGI2KqDHiRtq8lLVKyGBb2LzwgZ/9cM6OvphDqu1rxwAlSVrs+DT7AoOfwiXa3
Xg0DtOHhO2WlgVu5eFkVxhxiPZokp22KsQ6GFf/pp6BjaHP/E3GWx96si7+LM9l5QzZBfpjvelRD
8Ns14fBBmuAvlJ2up6KjZEWlnOu3TF5zX02TmpF9SPsdi+iZm/qG+P4uIO1U4gdt0nTaE3IhM/vX
rMkh8dSxxXObs7CsfQ0zLDlCqZgAfN4qFAZCJ3jiVmhDDUvXv55kSy3Xk1wDt+/AcSZ+i2qISwyu
y7SMIlNEfHy/o1OtnxJhvsWsXTzT6BYw6pqGRn+cI0Fup9hvBcJFhOFz0sba+b5X10Jk2amJs5RS
cpVj8WDQ9Ru8XPamy2UcNRnGowzFg/4Lo1myCFe6ovUggjRtKrVT7tLNUVaWyJR9jlFxVTps1FQs
4HLO7SFGFuvZHm8G3aJMPuI9l/ifiSiltqJ5aA+WSRwoVpIdBx+c6qrWwas4J/PAxCZVUETG/9sr
ZirdvJAYl/W90Qejjuu7ZnL9RrVs90L0iOfFMGPZpoVkuGnvGxXWBO65VXQpXuW1Riy+9srAYFzk
SIZmyELAlBOuQt7AZu+LNlt4e3ooOQbATubhHKi43vmnLx7McsgG6KJBjSmnb26VLRKgUfo61BcV
gLzrfLPwK7PX4JytqsFslOG8FLU/XHpSCqzr8+Uo5WqnEt0spnIRcgNbhF1qTyOkpTtdzPw890yb
jV32wXkDy0cvomPI7OOS21l2NkOE1zeNb2HKPdApIO0GxA2oJkq5/WtxLvAA7wY24AazSccT371r
p3PunIaq9XQEhP6wKDfLkvanOMp5GCLrsRXUXl9CkUtNJUb316XVhqc/V2nPpibSa/6LEecbo/gs
1FpjgMttedYeC0BdylDek/a+12K4dWalVg5RBXJ3al85ef44QxheoGgoEaXAsyaBXnUlh/dn8xod
i+uH0/9PZWRibNcXqqe4iv93Ej3K2Ge8MMPrl1i9Vs/S/2Y/YVOdJUGKJcDdlDfhtxh7bhdEmEDY
TtjIRn3ktqTFCJASSh5bzarZ4st3LZW05dXk9AzvpekeMHlMRRjCaQO+HhmGerG6REuQUR+FOb/t
lp58ouBAsHXZLGRHKhh4H6JU171Z/pighdLmnHDDNAUkzkhtDLHZc3Rk/p1gufLskJR2rROpQ7lu
Leu+7MdeWlqFU4IGwOh90OHK3CIMqAmDFhAVxWJ1yv8QYgNfZ0qcZeVpoE1AQAMLsoKEFfhAsutF
clyRnoD1Rv2v8V3fLyBSUyO/2h/46UG95YUmSfwnOZiqFt5mazhAIEiOwP/VPwPI2KLjmR+fWChE
v9ty1kmAV9xpZyrIqu9PXFw/3R0k+eiBJyn6rKAKE8VZau3tmIlFieOxZhNkl6Aq/PPI+4YoLEg3
yEsDjXri/iC/ArTRfAqVQ2wBSok173UKTVPpDHDonRqGV1WVjqlqcnKth8QW8SMZkHEvRbphaLhe
boY7/IRkl0gN0Po0vBDRzgxT28OV3NjJ7ceKji4zNnX2wvKoQpR9inyAPoKzL+2mlbIbky8nPmbF
ulq7eUvPXGwchphSZ8mA0ScHYXH4noIUx0yUn1kiraMUs4ZOAKXDQFR+4ZdX9IPJbeN1xn0ysqWP
8gck0qA0bL/UuVPEQHZdHNoes2iR+AyDZdMNv7kgX5pSJo6WZJyLjQs6dCGaaulOSHYhlJ4v7UZV
4w6n09nOWfXvRIyyExx4Qw2SkhYYTsqgyAHN2uatXd+cPpE3xXWlm43aN+oKY7ugYLPB8SAupYCS
TSeAaBQVPhRyy63FPT6qfiBKj6y+ltKSP4f2CFrfjBqoWW7uZf3CBZ5yvfJl65czfOtL5FfAq0cC
tYndQSKEBBVR7qaKa8qheXOCYVO+np3E0XSVbB1+z5ITZmQwh9EI5D7I3ZoEesOieYC+jK4QYrem
Ig2SlvvZpRtZe6O5R+/lrYW/9Y7qeOwgVEbyFT3VkI+oavHpsEGjh8YWEoiC1NnGiten/LvdGS55
hTDxgm03ZcvDlejSQbMf3rCkPJXaZ0exL7Nm83JVyXMo2AC8WzKL5ODWlFSo6+khEY6J1NJZkpJv
H+PKccHygIdVTXncvhKRjjJGsJotshPkb9JasKrpY/lVhRbfXl2Q/WvBoml9OEykWQY1sn8fejDN
/rYBFcz6SPwSzzsnlXFCcAUf5CocPZ41B2QK6j+viZeB8rEkNN+qN0F87ilRl5mg30ismExgHzVR
8QYcxTpYSe1rJJ7IsU7+75KYgwFo9zSZU0ioZhXgREstq44OBxHg5hKdONB2wJ6oHibV6MyhfKAA
79BMakrSzi0EDQ2huq35TYQDXEVC/ELn8/GwqyXuetU5XCw/9ZSuDzuNsfYcPZ68HRt5s0B1S7hT
/sq3W+Z6WIKArta71ppMGBGxFEzEsUF48F2ydjkD2azozHOzGto1/GWgNVcmpTfmykVI9CNOFn4Q
3l5bEcSHXl/Bt7/693/Fvt7MiHqgQ9Sb30R/ooIjT6XTah5kgYlE9CyrAWgbUm1F7+EKHIbjZDnS
tOmVnxV2sRm+O7MWE32mVk9Dc6t7O4FboqRAwXo5lLj3bhLpUc3Uy2wG05TmYUhLi2zI57fTuzUv
/PVKGhGpXV1glc3WgJSONNkBV8Izx/fH2oG5z319vpaapnj4AfAtFgQLpPlC4vhduv2iY0O0ypk4
qMwAdM1FwSdpv1c8vLO0JlxAzi0ForiVGp0BYoiN4uRa8nqJow51bKFwBgHJyvRqB1IG5Nxk0gg0
mvhOYXyJ3OlOboC1dXVnv7ElbehHIrj2CKwQdwZOHCBCF45L78tyUO0HjJKKMEiSkfsEqacyG/F6
fYFNrxEtfn1zmqDt5JOG9aFmFwXZiF6mLJjc7Xfsp5hJJ3eoz5YKPAJJohUwvjtTNMidJjXNYmrE
xYD3dtYQikKZnykDzD7V/qYDZ5+3mVEunEIPS8DJ0wGb/VpRMpFHxG9xz1Aa6/A4J842fsRYRTYa
MwT1RvmZpSJZD8D80oS09z4iOJuCZMFg1Fmh8k40EVNJp8uHoYy5i/qDl178UdncIWG9gddGOU7i
+UD90jtHsUJu84lQ938ttDCwWLeeBkaUehkC9wf+inqdovPrcpD1zLZiN7d7bcGnekBn0vFsG42C
EAsWAr67RHw5f1kaDL3bwAd7GWJEgBQC1d2d0MK7SFbJeVVqE3JwpChRauaVuJ4THx/aDTLjNuDM
gAZV3jVrRkKMxYflP7bP0Rvmkwn3mWGI0EZCsNn7fq57ePcNN/RHtTtw3b6+Cu7JubtE4Gf6c8hb
gHKYN1phvWAErm2nFW2K3vuNWQP17CiO7G+gzDn+OwJ+8ME7B0A8p1ycRUA5RyizrswKbIzdQFVs
qyfIt549++KId4DILALIVEbSNvuE13fAUBs3f/81G3kCrIPKk45Nors/2EDZ1Ke9h9afJAEVjKcX
XkmBjvEpuzJDcEhwKhg8PdZeHQGYXy3tQ5gt1ulCVjNVxvs/W7BGlUAE3akEZhJddOQsQSLlHbXG
ba+VRIxOpu2o98rcnEGNEj0+KtGTzZMDcxuDYxxcLD0WSNZIvTh5U09pqVfqNQbTuriECYgXlOTr
QtvCW1/wvNwV1nK3/f12C6sQ2TSGeyG44UdEpE9UBM8/k+cxj46XpB90lZGRPGCVJho9ENL6zUEJ
MGkN5LbmNPFJLG2hIjfekSrup90Ku19Ta+qhNdiHUneWYPvEBm2hEbo6MvSD1GrDnXGnEVztCiH1
huTdVFqvaRhFSaHk34mTTOUsjZK7hgl02iiZIM13C+IXJ1G+goLjk+yBdp7ARdPCfbGz3ppeA9Ha
ubGJrFciKrQ3V+WBXEnCmGyvvFRpz78OtFJkrGHZvIgo0Ks6gLEuR06fU0U1wMBhVb2lUToW6kEL
slj5fN2LXFLaHwltn/yL/TxBvjiSTjL0MxX6sIRxchB6B1LCbQ1CqPBkZqvJcun2bFH5A7B+7e+D
ecQgTYA21u4yA7SKTFglo1wDeqOkle/ECy9fbQYkkiLkfCyq3QjGLiKGdIPgUtn+rswqdE59Ur5P
WpXqW+5CLEF/JSgyU6nvztCFByUSGT3pfSfs3LmkY8iTwYgORfJC/qtUzTefH1D0XumisFkUtJa6
C55UPl+mJmUC0+tm9s+x3ARV0WuVfh9Y3ZYxY/MJaSWuKYjcpqt5CVgAtItRmGMW/T2tXNUjdsvd
HhOK91zgtwPooFhQjBiyMXdMM+BjJuZ6CsFAF89dllt3tTdMiqUMBY1K5NB1Gi5JdmYTX4T+8fx0
JDWdjuWMAMNCKP+nCj53nmWQ421/bvPkZpnMIYrGWxcdTKdK+q1V+JL9OoWgKM2S+lfwbaSKdPh9
oA83Z+oBMJ4lAfWiIgyzbreKvsekT6Glp6QAhAGtDDmEhkV0QrBUZ+BUO/reb4Bfrmw+I4rUpUNo
t+iaq3Wx2+OTcPizJJjXqIHCe6E4ExNPyE0ITEyjsy1e7lA2aoyzA23MtFL0Jli9zDU5rukRo/dE
69AxkcK0+Q0CZNN1YoOcMq6AWLD+KFUV1gcOZDdkVhahSi7kStF0mJxjqIctpUGE5E9pY1vvpmjr
2dwNLg518EbM4hmF8zVtEwGj8X2dSUyQZpFet8L/HNCIAFaCDO1yof0Qvp736pmzkawaaL7kQJRc
EbRnT9R/A2yPrnUkK0t7eKKw9sue3wcyS/xFJ3Z0HqHxOf+D5bsmPHjg8ecFW02+MxiFSDGjKbUx
Du22ZaJGbWOfAhd5dieREkNznpYRBgnqPjm1KhYU0vQb/HlwU2ufE6m5d+pjNSAmX1Ppm7ehVGhB
HgfcWmHCI1DBWQEP8Pj2mUrlGKOQqhNMPGbzNxOggueVmiVM6Bmm2zHIEzvp09LFegfd8iWNO1HS
SwQ5J/QJFSiiWqwn1diaH3FBnGGh5tlb/XdUzXDk2r34b1QWg9eZe23snoBYtsr0HTwKhb3r/peO
QxOvWbsMwAfcDtx3MSTDBXoAhP8fEpPrih+911hEs/4IxLF8/uCLYuLulOcRLBeroTv9RYkWGrEc
whKCuTFzfFk9p6KK5IlBfsm0ohQPsCMv4YtRQbAIDpcaaDEYh8Lm2gyFdVVRkhC5LxXPh6tyEXAh
QNU3mW2CkUl9f3BPe58hj3cijWQ7bF8Rq/TzGMHeDNQYOkSGsT49RiJJam5/9Y6OIq1nvbIGw/P4
QSRupXYlK7EcUCTFI2y5jWbUABJ7UIWPTISknZ54xprBTn6FGZQsXNxig89TJle16QwMtkTCUTB0
sOZOl0SamISnpqFVIlRUIaqXvYkLTEFG9rDl41+hYHgfrAajfKkM2tuLJzucNyTI47HZw4AVhJrM
VBP4bdYtNFyQymSrLjIkrQBeEPXyr86lzkx819VRn5X87SF2AHYahcEps2gVlENmNpIMH9CJQCIx
2HxL9zBke/bpdmNCuVppb4K9XAz53Xm771pQo4ly69Peq4sm1ADzblZdbhlXlvp0kgKeBUA3jCgb
BUHKzrCE4QPkONav4sSHM9svVbu0k1PBxM2nbI2k8E1xHX7vwRqz11xhB1fagERiJjg9+7/R1Agr
zNJ9hfSJLgalnnUYHvHlNR2Utkap7zB1+gQSj0jIV0Aen5c3aUrBOutcBPi5YKU7z8EW76guJy0f
UWlf993LkcDIQyQDEZnUjkmbN3Xay8IyR4/2BAcLqrsBo16otmKCrw7Zc+7o3uWWCF7xpQqFfeSW
TZ5Tp2LWGE2RFe/pwYbhz7LrD+UVvg+rtw2bqVBM3KF/FLW6Fl2QaxrJduDbpInZMcPM9Txeaes7
gwT7amM35lSRNTChu5c7CPeLH+mH1Mg7n/0b/Z6WMWgYFTVqopbJHAH3s/4iopbNd4frfZkDX42f
0OG0YA4zs94w+Es/Be/MCV4GztJHXbugNfEiK4WNEVVAqLGAl1+rOvkecrNA52lc+ly/oE5Z8b2u
9xS+xJSldH3WBU0XJ1STCGjjprmt1DGPC9Jw+NmtGs9YbdOQpI8uhQmA9Iup8g0WpWWJn3hLzgSJ
u2pfFSC3ExEKDeEoNSV93K9ensQyq1tVnX+IA4kiZ8B/JPOBnN4PQTB3VhTWAqj/lDr3bqURwBHQ
tIE9kGpv7PrMKaT4T308sI3p4Pn8cmmVQkg0KytW5nF1Zq4A8uxjWmjqgZtjN8G7DhUYgDotSX+x
urnFmjlIDmqUgCRT+zG1LUS9Tl95W9LHQkpjL6QIy/ObqRHqtPHBIlPQKJw2oBVk8qGc7/YcViM8
7jkEEfcXOff469CXVxZiw8f0GhYVGCkgVWs+80esg0ESQ7xC7vAnGh869zWGTxRcsTFfIX7YXF9R
xtAxGslzVBztPMXoLNCM63FSp1C3a9HZzIncF+7FS7cYycXbXj+vrfSKygZqgE4IzfqTW52PJu9z
ko2tktcpZjJudvSrw8cmfXunTbiEsEhBlX+ZLjMeXGsYupmCflmQXbJtNYPfURInqmaYKkXeCh7Z
5I5vcXsX+WNzmIQjWEgIt9ghSQu78EncyuyaFKR0TeSkOMxqup+3U8jXsIBFJFLEFTTSrJYVBtUP
VvkknuEW4XRUPnUzYK/ifRPEZoLkhxPgw9aVNH0v3ha56pfckGIKYa0d6agC0RyB+U7CHSxz5or0
c4MywbMHsCjhEq+bmAcI20/w/KcV/Svve3V/xdn84NQG4AL72ielKttow2Pk9VND1gb/FDBlXoTQ
YNNlpd346XYOjt5YvOnH3vtONU3rn2aSiYOW+iB7PSx0ALd3WD/y/MsjcVDbJ/LnkD9R/94lMLmN
RCLP52nJDzfBBxiyFYHxo9rzDqihVjqMl02vXCCPsheH711NPHUL6Efh8C27G5O8knEJ1ZjCCnEa
wg6o4ONscPb3VOsYfYzOkN9GeVxKiUa0kp4tf6v3i6GHbWT9lpPlJtVl8oPCq19H21fvlOpsLhTS
qlWxNF5/hIaG2bCCWLFpAMDdaPzSHPACZBiCa1705OtfQjkgy2wwf0M3rkIx4NONxn/rp+soCdNE
ET4JdYcnYJts8m5SRbjQk1iaKlYDb6te6JfJjj839FG9fn6pVAFYnNBRhFxrSYqXN4puGcl2Jqn5
/6N2cDiYsnisOIJ72LAlFGHZv36Dy0eWB524L6xizLDAuMMvMhHJlIuaaqtkeLjRiVHwY6whgyL+
7e7IscFbi1jI78bbFRJDJ4w/ptLgxpi1ptZsrDKZ5N+vYTyw8imqupuoadmVIQ8JO+P1P9RwiJOo
OniUHayW1QrLHj8z7EiFL9wPGFXemmSDHvM503aDBiBhKO2z/JzLHlN1M121vW7wV5GGb+c4Cucp
llWnUjBgabWeRW7kQzVTS7XGISGq8f30ufeOKSb9devSb2TZracU/Mjr6PcKorT/pwrwWsLjPRJr
Q1fCtIEbUx8Sz9niZ0/vHXj8wB4Xcp7zGkXocVXWo8/BfOVLhMkFa26Kx3+iR2XpVA04NmfN7HzK
hFyDz/FW1hpk3VOqPheygcGIsAcZddtRM5NdqvecjBIzDiTrKX8USOlzkRtZiWOx4VDUk8RVFuv+
cSUocWGaEyZICovKPKjduVVYhCQwh7Hmds6OIiL1TYJsS7ZMxDmj0UMRAUtYy5OXDjQsFGoGhnnk
a8JDpIM0en8e8WulbbnLvIMgTzFcVGu66NIXPYGAkEamdKDmlgTbnWsU0z0rh610+nJ3moYOPqnF
cVnzrWuoFkocwPxPahAImN/CsRxvArIDsdTd1JwcRIM/c0Mfi6ZsPm9I8H88xwksZZMOWQe15PJh
FmKpgzTiO8vDz3/a7JQenvEjMiJ07LM4Q4f+MCk19NbBA3N7oYfBBrlk2UIke5dZoIt1zLg3F+4U
ENoRCQkJMBzp9HBY+qRLe9tFtizNIr8VNFXDshSc5A2zk4JbxaDtGuujzwlo+EBpXggJNP4Zj/Oa
ZDdaLQKkpxdZmuSl7XuO08ZDBYXBnMPNLR1cDKvewDBT2esc3x0is+8yeLojADSEAv805uZL314F
qa0El1WTDW0t23bwbbUZgZzC7NmlwgTrcCk372Qhf2GDkftTK2l7oEH3UsNLLWfUItBTguQRP2A8
e9r0e8/sXiZ1Or9gu/L+yzc0BgNV4OPX7amcq8kZmvNDLb7AEfxwtcP6TpsmCVe3MN4aJhvX7Ece
iw41br4QVRCmlVXbLWQHyWk3WbofkihUphEgMzmJNf8L9cmg6PCqE7l2yUTQlcYemsKM/dDeD0Pf
bDPRRhbD2xOaXnYuBkmJ4j9lLSSoKsC5MlnBL6DYf0FPmrs+rhbz1Hcx4hE7ENCCs1DLlsiJSvUs
70WZk57MUfFuEejO/WOZ9UVFr5lfJV2ZnN6YtWnFVkc0r284EUA+gAe8FculsN/FewdIfjxG/DtD
POJgvpYm8jrlOe9aM9j/rthmGgR78Kf7M+uH+kiGAI1XQdn56rM5GdvgmYnJq6JSCeJWb5NYYtwR
NwNKENbUJ1kyLGk0tp+bFGSAVXBw1cbJwO97SKdr6pKuZWT4YvUniPGSz6h6XaBytcMAUi3hRiCH
62q3vvqGZ9NyBkCe9hc/tuc9Rfw7I7eJSQUykaNcrdBjaRWO2pdIVCpKJO8ECCjjdQ0ARjInbKfh
GDu0Vmx+YCcCLtx3zw5x6ZNxH/YSI5Ql49RmXGiy1cqFXZCqQtvuK0z9BQMe8jj6ikHLTo319b7j
3uxEXT5zwkYp/B4mbt0pTwcWyipQROq7g4WuvV/O9USWPrIjhpBcD66hq8MAvPnWNodEarzeO7n6
qMJ2nLY/boOxCtTfNsx4IQ0TroYfjsZ7XXT1gMwG0kZZlwpb9oZ1UyWKX5eNkRSVvSlGJnYG9WK/
CIxLQhurI0YUJzNl1jTF3bsZHGEsq3fI5fMeArd4h+tzGuylujYy/54H0+jxY3/vW15/4AU73xpf
e1XuZl9d/rj2QWU7ym5sGkYXb0jE0+ivd7s/xw0M5IaecqvkPQCBKb+zptl46XUZz1U5k70F7SyZ
IRozKr7j99Glgge/PO7i2ZOyQ1KuHkn9RcFxS7ER5cRuKGP3krQNWAnbm2GfMT+ZgpHahb/Ofh+O
M4+0z9vWYFQ9tRZTT1TTsisKto2xLZeruPWNhTrhxtIQFIaFeHQ4MjSENDkfzWhB+zgAadB+tmKg
9S6iVH6qeNPbL4YFIrvtauyFr4J46Yb8suNrQ+ZD0iKQd1D9JLNxHwvfXWgCbh+EHUZfsK6VIrrU
SL0zlsBCunaAO5zEyqgTxD5oE4JYPaq2P1Kp2zglbF0ji2d8ZsW2xouFFfKDecsesLx9piJZP7aG
+q7F/xiJbhYt6/98PIRbfSfoSpizl9/jCJCM+TN77tnqWN6+8xZCf7VF8yg9LhoN6j2dotbcEafE
aW5W56M3qDC8jjaIqqRX3KEkUmjrTJ0qGv4UchM3bMlrqr37JAqE6hHRC8W8eiHfvIZUNFovXc3t
W8oj4pYOPIfbdJ5sRrJqNiav44X8JrSZiUmcaQcN4GwiCg0uJpCTr7AhzM4lyOgh5yYV0Yv2DGeS
bOjkUohbq5L/Ua75eUirXy+j6bCyENyTF56Zf4wIf4HHR7QwQszNiLT/Pn175NC/A/TDbe1M6H/2
xxotoDhNLXZ2+DJViZCluzlVFAXnEqq04FSJNP77+KM8NSgiOb4jI/rJ+S1jjllvZLlhuSm6g3o3
1slP6Sh/MV/Svk3qEPiJLw3OmJfaxPiMKR+aVQIDVZKhcsQ7L4uKebrztXBb4NUk/1Aev+a696/z
f7KSMVHm8967kJG7Jexy+szoEhp+dAJCigABy08vjJrJRw6jxybxdKy13oBpXxmgl9DYCOxm85k4
ywR+8D3riXYlH3ROL8tgdoyGGeHOzvfhGkbu1MinoFzSBoKbrUZXGlCs1xqf6UVxyybnmYPWqiDZ
ThZGPSVS6FEajY90C5fDStH9eZz/c5822fE84oW7DHPTSyZlz4Ik4F2r4ueBgD8CeqgMgPh66MOp
ekwcNWYUovxLi6MQf/4iqyRXSreCf2Y6hODf3vseJyYcbpxXAIwbglNeoVD+GNKCyGu7zDlFlYXi
VExSFDXqHA0uq46g8E9XrYqG88nbn5B3kesnkprjgvG1w7cXIjTKUud/0QibvZqVqWgh3bg3bTh/
xoXOcmKTNn4FIa5T3BkknwV3yVs3JlGHRKOax5qSN/CB3pb2rDsNx/xwXXIxDlbjK7H9xT6006r3
7CdIQYI9LUuIi6lb0thHCYrPxEAmdktudeI+nmVLL/J2HPbtXOoNXF8TGNVie66eikJKTrfBQdr6
wJ8jhO+sgcvdoX1LboRgLHekVMjZoAgDkYkf87ZeKfL8S1UxIM7CT+lddUzQD4ootsZa4dk5fL+g
yhPSjwH8VAquhoHVXcrth11SALjXsP//OAcVuksMSubOf+xNjPEtRBav8KdtwoU8VfIt5XtdKagn
Pand47JfRMZA6rXaG+dWhltX9E6Lq/2/NhT9kyvqISe93mlYmsQdOP0L0a7/lKMpnn7HeybwMz9z
YJuAl9ArQY+NTLUAdeTN1n9Acg2CqXbRTt9zlKpQ5sX2y9earrvHrXKBq3xXwK+pclBUljlCqoZY
eXFKG+S0GJZBhpSzvDEHiyGOuRJjgeePYOYiZvUm1SVNQ1lZwZWViFG6qxdKvvRAvt5YiDNqI6E3
+U2eK0EtNK/qGQjlBe0KcE6LgxD5ugxh9UlN1SpN2gD/sfJkADEo70NR/RoMD0tm6+7WuONkUL58
gtI16tT75M3JIixiJUu6mTznfM2swHdnVbOc7hJzYLdXGgHmx0X5VwPI6EfUk39h/xV+1CuShxoN
6QWL7vkWYwA8k3RpEr3wgirsbp917O/3P0iSXXvuO1KoZv4o/qN6YaUhbzmp8KYiVWiUjPiFRKyw
BBVwbSNrD63b1QmszuCmKM1cLlLVRfj7XX4GdvUjrHSevD1r1Lan7HQ8pcjM+hw9VsQfyIICvJ9M
Sj1Rpw/O8dX1CChchOMpnxKcRudXhPvMR3JjHUABp+zG9fLIzSP3W7tZEbrvA6g++Fjckj7za1ZB
L09ehw/6REM7crmyEyOAksV3BHc6G0zh6a1gPViiu72HGDBum66nMWYrT0yuYhIdPr2d+2rwaXjl
uFVu6zIEzMHsMVm8D1GVpimjvng5KjfOVuAZyUohxd/3t0hKNSpMYc63glL7ZiXcrsWIfObu8hwr
5Mlmqs65F/HoH0tWE2JEQRg7BHSNMSr8Pajd1ZLDcladLmO56AkcIIfdYUwjHnU9hAdTLAfCDcvk
AwbeDkkDNuUnHtZmeT3FUzCAk4lKD7el/ZmJZ4INiMdqdxI3m/1uVnbjp6ri2gdDnnhyCaKDNopL
JskY0/UEY4VFEMYN+wmh4VecZo6DH8pUn2lr9lu7TUvbVwmGXzQVFKPmWLLyeD7PoUZmr/84GtRn
p5as/vlbCZa0fKautUT3exELSyQkaKeHyiktPRTH4tP3BNf9JLJCd79lN5McwNvv7h5fxCHVRemn
uIRm6D6/NwYe86NGEmsgNM79cHatkkxsCXEqLMdtPbswbWvgtD1Mmozsze+mEuL1kIrNnbukxAmJ
Nh5lsNfQMVkwsxc4QItiGm+qZur1bAVaIm/Yvf/kKaKh6qs9iWiPxcH+nDrsyHo6aH5VeP9sCTVM
Z8YCsvegd8GhtcF4fWi+F+3hx5HwdFtGrDQ2DIcnGATz57b1MP8jaMJzALtCzTOSVIe+qUTJkt7M
ArdCWBV8GnBXgT4mGt/YferMsWN+9M26GVoy8yWxO8uOFb7zE6Ul6s9VxSIlN/Y4qMcW79FXXoSY
QbQWxC+WJ27JevrY5/gZhhJJdDQ9Ov3wXGvpCMR7P2Fd0vy7IFG6pYFb4sngEPMycUupLuH28DsO
4ENVrsJY8/cZemhSh04UDcO+3TtY/NGlqXOQ0h/kqcyLgOPYHf8fLolXPR2uEuIY+3HVYsen97Nl
mrvcycompmZ1SRm+vEhPkPPk2yFLzrMAdAZhSJ8Hi/Edu0vqTVnHZUhyjiHNLqr90UWNXCFGeoVz
+rE+o0OshSvYK2ISq3B+cvWSRhFIygaujHHD/YnCgc8QH6S6nLDOOJFPz/VxKGi9Exg3yKAtXUOc
Z7f0/FPlxmCfQeZnC0h8ilxAoRxPfumXb4tUOCsMcFdyBSLvQCc+7fxB7x9zjAzd7BmXIU01vthF
hedcN5q9ZqLifmIDUXThHxhbMZKS4s507w1nfun2u4bbZ2K8XQdiqTV4comIsoD9axEfQQXWrnem
qmbXqWXaLT/4uhCvXpdjrTmFETi4qxrHxyjZKDj7XsK/pMAaAVZGsvGZjp6/9eFKIHyX/Od3Lx58
qhHtNenSIAu3PwidRGjTv+foyL8lO2aw/UMo0YjSjTrxxAWhDvZWB+/WH7Zb2Kd84ZI9wS40+qZC
ta5vmdcmo1Ye9lzrxtottaHbOAkkaIbzmVAel51ATuFDIwVcbp9eP6fw0u3TIfCsogdJ1lwR1SBl
lJ7EnO4kkdInbjo0hZiit4DanJaAXHj9UifYfP1u0NIxSDd2R9QDb+7OEBQ8O7r+f1MWB3jG3Vy/
PWY3PhFAhDtMZ/UU6Y4iTtZ2MRD+fcm5YBSVijOJPv9dOLDx1bp30CE/joycH3vRzjAc/rHm9it4
TTpsrevEujSvx2lY/lOwLrMe/rZylnXenQGecTRZyrNgPcMDr80/tKoNVGlk1couYSemL0KXZulI
QSpaROLOnXFvTjS15andKXigMdBoA9al9/5PczWWh4sBkMjSRGmtbjyFeLnWOZ7ZAlu4wncA9wiE
q5VeU1f4WjZaH23Nk92Bjpg1zFsmnJlkl/OTWlWx1PO3TjtSkk2q6bcbb9eMJj9vJPTAj7YzhCdQ
ku5JjREj6g2G7cxK0EV6X8Rcm58GIektnv9OTSr9NG0o2GrKjkI9pt6R2eOWBhOFAPpxbbdL3xP3
cQ1XnmySLEfQhoXRoSnljYmjoDLqqCUJ8WYaCx7ygsd3QTWhkpRPGE9GECoPsxCK8mkddhvvzeZI
8W4s66TnaChX1Va3nSaQuksTTy9gmjgoo/Z63dfTGXPvY8sDPqJfKw9AKbFh25QmpQRPF465EEn+
gSH5ValJy5vUbOPu/h7t2sdhMep3g6wA8KncsK6aeQvJ0n7sQViWGwNmZz0FHYcLXjnTlVUU1J/m
mMza2SNsJ3A1ZHR16LprnqiHewfjF8SIMPsVZTAgoQloB5wgaq62rRrbA/EN440al3LB9OLXQaxf
0C2VtF5gNrYPPMW/S7NlNDs8439ERErvz/5iCI0io79sGSF+5ocnicpIqmCyldYmSJV5FpIgUlc6
v7o/6QzZDXrL5e62vogKhPmZcLBbzBEVWf1C6Kw+sUKm3Vdj+TWrLvFvRsuhQ6TXC7n0i7KF9Jgp
f05ezEigi2rKvTVBn+nS0a8LuK3VmdV83Y1ZKC1dqmAjnhqa4u14tuwxHk8gv44dP4w6dIfzKWSN
YOQ1QA5L6sMTwWNj2LN/usRJyuWoVm5FStg5Oe7v7NgewEC8ELiM2431AL4wlRu5dKmp/urZwaMn
RmSNzXXA/HoloH7X+8jrrieKwANggXcndZ6r+b1YC5Bh8ac1G4ytGgFHWDvtGYpHJpUzzUqnH6Qk
I+q6GywVkSbrGCRmUugBgbPvnXLUO9l8KarqOicD5sgRJwksKzowWDfgV8seTcFOFmEYJ12PaDYl
i5/uHxxnOd+sDkpkwq5EP1SM58wz0DuKyshakzxtApOjUAMXiQNdcv3nvthD1Yf1IQIi/B1+bO2L
Mpa7tkcG+18v7IX/de30z4OJ9HF8uAqAUQKM7GfGHjRgpCTsxkd6SkxZmTkZ9Dly8PQV1EGSvapv
TwEx4C1TD5grB43IB2s139gzhrWvjHKdo6VdSNEq6jYc91qj2VrjwfjJ73zejp2758MXjLTCmqLB
9SIGsxSOwz6/G2WZojeyofPmEm2Q594zUH22sUOtjkGeh4EiWLP0ZvTL5YvIMfLC4PRTKU7hI2/i
UCzCwO3gEpoiV5XokunDqqCe2jNkEIv1YoRS2eckE9w5Nbuh1xPtuFk0rH3YigNXraQoGFAhVhc9
NMp68BbngEp5ac2pOMyABuENDwdXpxCP/zSIE6I5RzoezcT5fN/x6geCvKlw/+Fj1yahgpesnYCF
xZz1QeQUp7Bn/NMEu+MGydp0fv2Dy/qrBKj/9pPKaMriJ8udC587+TORmAuCADCaWIAL8I1M38V5
ghwuxLiuksEn4B9FW5kEPoBLPafR4eROpMma6Wceq4QE+cnpy0shSsAf9l5OV44HRhWnr2Bs6lfJ
oLeSxwBFTF4ik0/apTvyMHzGfu4mN9hUg1+dtR0XSgDGYQ1ZJ3KeqeUxAC+nQeRC5VN4Y76Ba7aI
d6FgILNTZdMv5wL3OLwShuGpvQVO0CpBFuc3anWnbksBXVY4fMnZtSbjF66AEZFP+gnI7Hk+pfr5
SHpS4TpX1RS+aesJW4AMqkvOpyIhOwD7P6KbTut+z71BKn/jlrtTrlrMlVQRkZGCeUugkP7qO3uP
Z/iBUSPFmZC1GPEIA4n3eaZczeUXLdcIgp7lGUZ72eY3GQ9igWy+D80knBZQVpm3ZYCjHuafX/sT
Ehe2EaqeM9Wto9W/wMofp0r6G6OPnB4AfGbrN9xoJ4JyIjI3dPYcsa5Qsi0TTWUvnUJzz1T/VQrI
USmNZqF/+k26gxxt9LRoi/+xhZBPp3dWK6L6WS5I4H1f29juwrN3/CSe/koJA26/sT082u0ohGgn
iuG34mP2WBIHPWGKZrwKAj2QHXNHpVhCx9zfrU+KuXt6lV2h1rSPQUUqcIkuhJW+2Zqz2GmWsk5r
P/lkni4GnytTVyiDyJWuPAOxDt+nAWc7EkAU8G/m7TqDFsA7FHMSer1B4EQ1zUofGjGaZaKz1T8E
NMNtOieoJU759m+LQx3aDiqSu45mMcBtwb9p9ZItNm4pdosNm51S2qc+sSI9LLtPYAoxSpgQkJtE
Tqs5D0i/DPUHXGhghvpp7twi5vBsJPORU/56BAhwOx2cT2DEIt1e+aMAjh399Gtpfed70gEQCCGU
jF4f7sp7tvroJ4xV8w/BdmXUHV0ZFC/k03YNtbglVZbrtYXyzOZrR+WIKYqtfkJikc1ikGJ4Bbho
p+HL19vN9A9tq3/VxSKefuHLdWDrSv7n4cl2Da9mOF6+5wGXoMRgI32KQ11vL8BvbUoww/8oNPSN
KHdNAjF+fPWf/TEcpBY86tvuLE1BoLgfN3tZKb9YzFRUyKbYr5UpCSpLS4XnNCrQCT4WGXIL0woH
o4A0vwFpJOwMsi3vdl696JANtaVw8DTxOsm0lEpinjAXuGmJWWJrobZyPbT/JjYYvmPuXSbiNBRS
qPp3qkEFiTs4qUFIptGUcnQN7AQn0bh/pH8k5sYoUW11BQatCgVEW76vU+1jKGVo474yt2ln+Fly
CZYk40UaDds2RUGdLNGNZVGlMLsjZMG6SxJ3JFCgF8sQ6fPIOySh3nMdQ6t+Oac0cU6ur0D+GQcW
nDXVZYHPIboaEFqeXRiK7LmSIY23OqcKbWfMnb2qsIq+F9SawtYRvwwYH/wpwVKke7FK9IirRF+/
e/VeuR24tXNL53gvqMBBsL5IGN5LmRWQx0++gOFptqM7YJZ5CDIle8Dnij+3gUNtQDAGfHIKI4SZ
ZRwWWJdEW3aFJAvH+tQihfbWdeBaqqBDAwSnsjxTeMeYBU9RA/mLftNEiFD1sdWXo9bSWhh3dkbK
2X3vKeqp4hQJmh1Owwmr1Whh6Rbt+mR0Fqlqn3kfsG9ZLbcilGmejWjETbUt9Ymu8WXirMb7V/+q
XNJJhh2HTo+YpMehuDQHV72UQkG2LrTB4+JzKTKoYvNeNf1zI37RA83zjC4WDDrgyawzflDpd4vZ
72xoTLk+qbyojm6BuROpeFedFg6tuPEzn0knaFWGSiFbU4Y8ZtVY7rQEyCYtfQRjKFIxnum51RZP
nKJTVv/GGCWo0lAGdm9p6nWoXPTRWJjW9W/tW2CVnEDDuFD2JYw21HivM5+nHfcXjydJ2jiBT4dZ
QC6QG5A+zPJtbj/zanhq4AkOn+vzZA/gyTSdoXhHHUPtqWdGtIh+0QlG8YJw6QqYzMHClVmjVGga
gxj0+wLpXT228f8Q2uUl5SBB6y4WD7Xut5STLCZ4a82Wy2XykX4chi9bi7K5otSEqDGIijkEh9zV
DSStR9IOujc2zTJU2WnQh2czYtyx/IVhoXse+SjDqSMfWy8fMPWTyVT9xB2sFwHvdVcZx7ktYA2o
woEPjj7wHqEVzTfuZ7ybJMLMHrqrFQmNdC47h48uIGIxFcWcjbT+DixjQkfEBP6lL7dAabMU6GBW
Gg3JifVFGL9NvOKYNcS6O4bTAG5/nEDlzdKSiWvc61KdpSNAvM2YAQKmGNqk1lHWgtBp8H29TJ8+
7KS1vc/lZVGkbPVTQDnfOzvEPjKdJBElJUK/vIuj9b1Ek0fcsu+m2be6Y7e2UvyAj1RBjJhYmEDv
U5ySCHruIn/0DlqXT4MhAPSkhJco1L9owmd44xFLhe9SEGhXj68r2udfeQPdOZhFztWlchsFBpeb
gXvf6rtzZlXfDyyB28w+pQyk/pqEm/FDz2Z3S1gtJuD7wXByxJBIusFun04znO7Yks+yprYbh+df
8RtMJyzbHQ+SMEjf64rRNrdB9JrHcmpTe1Atj7EWgZ/JjWR++o2IucZR5lpl9ns7J/M3mbfrMCus
N/UbaU+9N/KlEZCgO9/OReut1oZlUlQSkkoAE3q/rlhmyuh57rbGQcznLxSOPYBTGU7l7Ony2JHo
6gFDX4UaiqIPRot7nWEIaO+B26S+AStu28DeBXKy0TvcaN3td1PMb19W7eox5xrPn8tGC7TyH6g4
EHuamxCMBp/z5WIt6iy3YGu2HFpxAsjyExuOA7nuJReOukDNJ7NCw3POTBl3hcFcdlmJ41C3vkQV
hxR+HV1oF3I/OpSdtzwU/IvNNXtAXvZy9dkYm1tYYJsR6Q+rnTaILc2vVTw+xb9SXvMFFW9fLbcI
IV5d50775tIcnRszZay3EeVxzAKREBNWP2k5KZCTGmRRLrybG525iROkszstiR//WoTMfn7uEdGd
dk6p9DkHFCVZm2lss8lICe2xrhQdsXgVPzB9zvKOZfgGB1gFU4jzyGRxjzmEGT0vk5RT4PhzBRGA
E2n9Ts40Fs9h3bZx597j3nBL0Ug1VTwaRWJ971ywl5E8vcieHHVIXcy9TLoiukn1kvnAK0ddLa/B
G1IUSQ/Glfg0lgfeZjcoa5EazqSpIesjwTmtC2gcRXEiUOJI+DgNSmgI/qDbmKmcvN7WLLNozNzh
yKM1PMCM5JdpQ8Ons7NzW6VCtReLe+oacQW1Qw2+SxvK1mwHzp7v4D8RqvJJ7oIlTBiwuM8RyCUf
tRvlgJ8wRtR5pNj++m7zc3OGXp021kBcTb0cYkcOj45RpvEys/DxuLtuTPnUbpKRamOJ5QXtGFi3
sUZX/laD4qSZU6CmDq78yf5IdQEsRbdl/jAVSv55yWpKsbYb2/fJAoJzzXkDjDNs0AJZVY6UQzE4
V4ps2Jb+vhwN0Of6r5sF8xIbZZ+MHmZXp9EAK3NxLDBgr9Wbly8XR2a7iurmTkBklnAInRMLK6MT
99GoyI2e+zD69w0IbYmHD5wBKx/L+Zn6r8tN8h74V8nHBhCGpERiawQjaaoo5rXmXrGaKPbiACRQ
qWt8oiOwQbymx4/wEfyFeWH7sQ+m7dxwJfYVypb4umCNIoGhXA6+G7PGbRJ9eQpD4k607Racg+yS
H3Kh7Qh3BEK8clBJieEos4pv9cPhtyEd5MJlB5m5+6gjyxg9GjMEhZCAKeCt7AVouJcXTmi06nqL
yDgjZViOhVHMNxXAyN2rPAE1G25uDa/5v/Lil2nLxKF9Evu1tXYRS5gGys6vfBWVb6T+zaUDTkxE
ZdKDjDNBUfceyXX5HrnjiayBbSs+3xSU1K4CLBI+RP+Jum0iZ1kXf1CX0mUQP0tnsSrvNJ5GnB5J
ZOFbyULlNJUR3Ytp2InWTIsjyg6DgFqPaLethYd6+hNvwALDjWtkOnw7p0lH7sa15vMvBw9hMqf7
S+gbYdrRbJw6jmLGNxdMzOB3Gp1jecqYLEKbhkCvGp0w8DrkJQdemCYWKaYf1TBYoN8bUQiYMdQw
FQCFw1o+sCzK8JQvRlD6f6tELJKbUpVkxr3oAdue4qRVoGflfRceBVRrIH6n1rMY6sdbIN132DwJ
xrzIZJyk8Ttot5yYlBqYUQIaxsEc7YWXoFcP1Ax6D2F1a4k1U9aX5t4exrNHS1LIRlhg4xRyre6n
MlLyQLY1ukmq5cIRG/2bUDyZU4NKwB8WWpvPVS0KDjYRPQLgY0qQCPL9CtGdA003kp5QaahoV2KR
Lgw//1OQzmViKeWBeuij73Uz2xrY1zjvs0N6GCLWpE4jJa+s551dX8W2Kt9d7xFDocg1NuS7qu5q
0pvuBOoGYIdUbFjLhPCkPP0yZxckoaw3nBDQUFDgtYukxTMb6uZSkBzKDXr0Ju7tOF/6XMBfereb
xm7a/ZUBCe9I4hTjPkeN0B08TJ1PVYtLaLJS69veV95D670xkEpfQTpZ6RtF2FDgdVZy4w6A/ZQc
XicaUBmnQoFEOb7xnN4yBCIkPUncTKYsgGy6Pkn3xyvfraCDOklbKGkMZed+TV/g0flSCBgEQv+O
XBQkkZBFPgUJvjXaDmJml8SGpy3GPwNq8kXNP3j8wTZT3fdoK93KobaVKH/pCPPSUi4dnkKG/P38
2+M/z0UhMwdOTgHaoW02NpcTPsrykD2f37h3VCVsPapAomQ4vQya6wLGRDcJME8KuI0+SILo2pcV
svxIb0OnmwwUKRZiVSrnFUdNIOR0x1a2hQuVItXZwsEg8Tqx+WZXDiCw28y3MK5MEsT6pDOXOxlO
m5v2kK+YxzfvXSlmSo4AXdBGCXOcP7lubMA1y6p7unU72yKLkQ1x7b5p6reW7YBl44q9VGOOLtOP
XPcvbYWec3C7f/H/YLMUjHfkmWbGyTa5LKs6SvudQVr8nBGqogPEM0aVquigYi0FA02wxZN38UMY
vvddB93hj1Ogqqzpo/fVjCbfLAl6c3E8edtkM8LZhBwdcZ1qt6d9NjSBqKv67k/+jIADQrsW/Pnm
U0adWIypCH2M67Lk3fYHE9MXAOa+5thgWDiBRatQ8YmFSgMb5e9L0prWI9KCwdxYjOdoub2u1rhM
saCSMqcGOd1GRj0Y/XjgDrO56oEqyHpBetPJZunyeleT+Vwmb0WQXbGfNAlIxtOpT3xfQGxkEUgA
ESoPiukuOWo8582lclfJhAsGxWGbX3DmYMSEzGiQ1QZsVpo4J9aA/KZa6N3RsVyFecq5rD0KbTl2
l7W5QV9ynNTtUN+BeRDXU0NAYFuNEY2DgjMwVqXs15OmGfTUuDKvlIwQHQ62q8bwsKaS0HtysBrq
P5SaWzSxQH16hNDC2v99zlaT8p4uQ54VoHwEukb+y6yEFTlvkQ35o2u6TttIwOXapxhecT8C5lH/
SCKTavHImMwo1UhW7u7UjlRuyASgVn75BM2QRmLoGG5cpix5I0gBoUbczOS1yqslM7TLKNB4ET4b
B2gB9fYwW+KFeuGKqjkfBQb97Owuv/vCepzIH8aG+yNtVV0HTpWh0dGQNhq6dIRp/doL2zo2GKYO
TfFOAqk1Hp8t31kei2txhqQdf50+yqvvUSy+lEgPi2XlQ3CswjmgH8eJpPcFtfzLEqlfmqn+JIF8
l61IwC0izs4nCT5HMAfWBfF6mcDg90DaOLS906cK1+baSnV+7/jgzVsJRFtC1Yhiu41wAjnrYmLo
/2cJF29SirBqKoeFwyVxTwx3IMGS2NcmO/rWccZCKKrJiUr9bxRuNK4zIwpafnTJ4KzpqzVft0Uc
6gkaXru0H0wED1GuIspM0cXYP8W0MrjCX2D4VqakhcZ6x0qheyqZOhpOeFGiIXT/m8c+fLSkizFU
SVpKBnppgqmUST6wHOuFXFEveq0+kgayjwRA5VssmWtYz31kbYJWskvB35TKmAuqOKTRF/RbfUv6
QJmA3cUp/CDUuQ9XMRXs6KbdOTGigMPwaMQ0cizpQP8SVB5g1Py3mOBBwMYDmPtpmYcO7dQ+CSJu
K0kX5mr8PzJSjtrM84YY69ctssERqMCwZ/6HjgDZEyoYS+rHxEVpuNcmCS4RmsF0yYKK/byIiBIm
dT6p/TgKUyaIQlJQGJTHPQlIYRKt8L6VM87+Tsr4wbcKqdQ5dDJPZT9JIsooLHxrCzmsIgAMjYaI
WQ6HgxWLDC92f1B19qc80QKAemphpdvIr/kP8Gc8E8g+Y9/A72I4KdL2uDb77zAe+zmvrygVG0WI
9mX9zqr07Ma2PdfXkNntUKAvdSTRpZ5s0AWNdxicTNs362TPuWC93rhG9auw59kYf5djEZUSID4D
7Phr91N/bmkkl6AP/8NfT3YEZQ2PGJvMxarJiBzQ/428SCoOgQiXinwg/CNT3a9hO4zAwYtuKQq8
j64yWSyL7MZAhF4Tkfyae9dz8ognSNpIGAXo0+0rcpJd9bY5sG26QqTQ3NOREXKmb7TRA1ZZpTAt
qUhfKj6Frk17sky945W9BqEJdlyDEDLs5bMQvBbfgBVpeSb96aTq8NB0koONY9cmQtn+VUmaDYg7
RihTkcJCnIgtbq2gUMYv6jXp1Yxaje1Rb6ENMtpnm1ijR84V228tzK1o0hxQEqxgCT8Uka2edcYB
SgBZagbPejsSXrJYqTk4T6HfEVqXeC6fjK88cLxNOF5gQAYo1bmQvC+iOYFtrZYss2ZtFPNR7zFQ
d2Au0F83m5cwbCOqVIar9PLl8jAkm8ex6P+JopPdL7J57aT1wfGkNAItXj+yYsa/6OTwX2mmLYGC
PnFWdJ+jrwbpXmf3vaUto3kC26a56don/w1Vcsrbgw5sLqYiJ1uWl5ex8ZcX2wrwuUfJjea5Sffu
mtT4OPMJlsS1T/HgdcqRnDauc5dMsax49hnzTp5ZRHECI64Z4Jd140Fown0rnTN/dPikdxNKJeRF
o5L3z5s9cBwZri8VUIx7V8rcZUDDwKdo/g+Z+qE+5cuyn7qWqgM7IBy3ehc5nKwltx3v+KBQkyFf
8zPSq8xsGxz6wuLrA7yfWPOmuxyYCajVQCQ1oP0Cq5liMUmO9lhOOXBghsOHI/4CHs2m8HPQkj7Z
WEwWT5AjSqsm1pEspCeykex0j+Q+vAuxcOozenSzarwUMwcCQoY4SRzrrqgRdzk9T+CCOPQ1T3Sv
aqvAbl3WMcR9jdZuL2tiJeuuLU6443Qgu+hxkkpQeN0tw2BsRmh8fR5vef+lSz6Vz7D3Go7qppxh
y1lMeElRaA3+goHI4CSp495wfqsGu/YUX3+vntkXUwpLZ9DRokt0t2RO6q7amCKn/Wr3Y8418Go2
EZlxJQSTFBVjxvgYDHMqGURQJhwvwHYGvz3ICfpjp44teNVq0Ff+P6SJXc0JLqXDAibMp1T/c6OT
K4Pe0fzgFLocepYxE8dvZ7KX/vNir5MQ7vWXIDuSN+MYDi4RIMqZLmt2bfu3x2BAq3boQ7OAwKdZ
NpIzSjIAbnHkNSIB4ec8oQpccTojR8Hqq5rvNjiDBH4O7zrLR9pbwdcDLqjbd398eEVmtIzrMHPZ
bNXV04266juXkxlhrvrkJOgNrYa06WF2yn1+U/mv0tmI9rl+BEivZGLULB0IXhHr6jugtf/mhrFR
8pBNkZ9MF06OcaCVT/ZA9tnPFDF2RgfeHMSsLtKls0V5+6WXaAYlwXRvoMks3yNTjJqpiM4u1Hb0
RAE9kqVCG/2eHvJJ//g8yHnIxYuDKzGE41JCZQxbHzKOMHY25TVt2nKqZ58iQ0XoBdX6FkFrYZ3u
yWnVEl7Wktw538UyAM8DY52g5nD3JGI5mrb4c+c5exU12VDivJ6PMEdCC0ePMTHepXaqEhE9GMgj
ENaNHCHWhGc2vN2UebtV52KeLzcqLJZbFkkkl/u2z1Bjeaf+Kufjyli274oDY53nEsyVs1DPw8Dz
rW50XV5e8awyujQ6120iodiAS6WqTJDxH9yfRVaQrFiu5XnQJMDEwZ0PyAzIAPYKXD4obq8wpVXP
fmNupxnFJjRVRiXjTCwsGyyHNzIE5mhvOB1Qp04QkGFjBQb4Pm1lHljnQr5NyVv97fiERr+t6YAd
Oz5Z04WmTG2JKdkSdoQBfjOMjnAuPyB9q3QV4NZHheAO89nVhRKKvXyNftwQiUr/vnSqqhi5/Kri
AIYEXexw0os2WowjMFg3pg2yhf//Tkof5eWaAwYETxvQJtNU2RjUpnFx5WMaKwiqHpYL8KmeW4VT
+Jvf640M7aWlf8uXw2dQko/CnqW4J9A3Poku9XzqsSq1V3A9L/PW1ln6Uw95+20w3X91n3pCRqsx
vh5JMSII+QGC7IcbtmAvjFAbBtfQpu69RGeTdMZCa2II0HSIyPoiFWIC/imQ58r6XTnDUKOGoKIo
D1M1RpeTE6P5dXW89upTuUbRM9LyjmzxW0jvvnOKQdasU9Rb0Q9H5bee1KK/atVFqhLfOi7p3mgw
NPmxw/BdGLUYiXgKKV96b1zrw5NUpBKHAVVgG/dgS92qsGLHp5/BcB3TkVAs/lGlZ5IFBZyqqrXu
pg5GisMtDWR59IEKBNl/r75NM3E5kY1Vjgz8UodnTzxYw/7q1FdwnGgx1UWXXFJHhN5QsnHWUVNq
9v1TUutHjBBawcVEdTnLyKU5pR7ZPo8oa1erfqu1JFRrmjZB2BLY+isX5DFtPgiuyvocqNKaWv1e
e3ZrnS0aJEKPX7bQQuZW0ZbuNyG6NxpipGUHdhzTwKR56eFobAnTovw9v0an2ojNODzN2WrZJpHx
jSlAYhpysacqsE9Tyr8NCiUB+LmNYutS7AF8qYoDe7wRlO6Zn04I4mFimsODehuYm0BjwqfyQYz1
TWw5y/sH3l4rtRb6aERBw8GahAYWNigz+Ey3HhViUBXpBiWy2Lac2j/77ozHOdpqKB70uEKT5ynn
ULhijA6f4yoFcNX2tGc+fpgabpho6qkvBNTmusAXnzPXMeQh77V45ZffpmOevxJO3600dxuq645q
BpJJJXbFbpb++wrZJ/sS5lOsA1EELTfRmPAs4EIn0fnPU2F7YX14QLJxTBfGOhWQ/NhnPNeqOQHf
E4yJ/5H7AbhPYhYwzmmWaZye5lMdLsWROVQKVMy0T1fCfrkbm8I2yJmsLze26F2XsRltjqai3Krg
Bs0hZjSf+IXDyrpkATN3xzLBffbygC4IJiTA+MmBj5s6ArLVQNyPu/5gZzc6IVhoMNlstT56fqcx
9Gttkav9YOYUwkAmZszdxki6x8wuopKxFMNh2wYHyksuRHhLm8SGMAsZ1h0f24mxtk/E40jJ9kHb
PZqL/JL7WXtheH/XB5lzZ7NAVfKQCUMOjCMsTHubzHsfxB8DB6Iz4DbJIE0BhJOMqOKVxRum6//o
BNX3AAp4XFcfHdK8QAwkaRjZBVtEW9ES/Lvhcx7R2nWoVZ9C4HQ8WeChUQQiwZGuLtoU03YeBCU3
iJNcu21B1nwrVsoCRt3GpxRSsAA50weIVObafdiYSfbL7xy2+5OO6ZMmg8ZAMTu5QSdYX5Zmo8WJ
c5UpxfpOvk0+tGaut5x31c+nxT9rLWYAahz8d9niNVDAApnJhVdQSXu0JVmxKrCb7qDI4nfTvO0s
LlVHbY7oNBeAb+b8HE0LNmcnS2sqORN/3y0jUa5QPmozkYdG2eLhnN/cNJ1vhI/sr8RaP1HGBKyK
oB+Ie3/3HdAPtDbH62+9olHMFU2MoLU06s3RIDjL+wqqK6DIlSKJlw/iDu6JGLOeNumpBKgftwOR
4l1vsqYpaGvrSVXREpDBE2mel/UoW0GKB/LzzUVYJRfvY55JCBUWUE+Uzx9cbkRwt6ewYEbHOreq
Usx0mhG8uZ2m2nqayVrAZ3CIms45y7pRCa0aZTwvB2Tcnu5kbXA0DBbIv/izM8ck078jOO2ND0Zl
v+XsAiyGl7jt/cz6CsLJ7JJp5lHDkm5HzXdfmIZCnD6x6SUW8OO7wLsZ1+w92c/OSizQthf/oCCp
REqCEmQGnrBCyQL0VNu99HLjv50D3E9D4tbz/AyZFvMBmoUrRQTIgyoWt1yT/0kPpj6QEK1PiNcB
HUOWRWE3iT2+TXBdDVyhGFRU4nmB3tXUJtK8rU/+yI7Hp8RgUpkeDeLT84jV23VRNDwkKeBR0fQp
VFLfl/YypmwS8+X5/hEIzvC0SD+LaarkTiztXRPWXxcbZ1MiB97HpnDJOdqQj3PBtRk2+eOTDAPF
euaX9Ihc+PfjyZ5SaHLAR2HoO7Utmc1bCRITECv1F9xxNK/KNI2QcmGDZ7Y28v3+wOA9lexZW3sf
IwSZB3xCw6/nNl6zUJKtk8HPKeYpHBvBKntApntiltx5hkNU6dwzfGthpz2EkorLflkm5kXclB4F
etxII2h7aBE0HyoSbaAdfruk7+1i2yflN0yVgKvGSxrzAydcBZ4f0bPLHaD5DuCeecWyiZFfH+3K
eabJ5B1oAF2qW+U5ZOUmirGKPqNZ/HDAJX7vjnZ4lxj1GlhAPnv4JTpU6wflVDhTnDj8PVpaoDtV
nOsk2SnixcXSCbGl8fiMnUg4wEZswuzfXZx0B+/AIiYxt14gOUpRVOVvO7lpNG+QNhpTuwJ/nG4r
hOELfynysNgnUN+iRCr6abtuv5ddCnGJVsPJEGqCv39pWkwSv99xiF/96Xg8if+jLYurzy9Vol1f
+TICF0X9d5WsMup8WMZzbhqjFIODJnviVPnzp56DbPRRu2a10oLHJfiqH0Qiz2VmiNL6XN4nYKSr
MT3rKzNlpFgihDFeG9NGXitl0RkTNOfMtauWaQWrk+rYPZw0tV+vlo8SBW0ngVxJYKeICu9Msn6S
FyZXyZ67WZ8qMpCaz6a3bxoXyL8AUIkvWlAOLIajsdoTaBPGtAPIbjBBi/CvePpMjoipyZu37rXs
5wf1pMAr+S1XTqro+UiX2Ggl/AVkxOHCN4nXaUJKSxNeoNsECK6BO+Is1DReuUt867Z4vhY50Vz2
1k1huXctG3SRs2kjeeO9txzupBjN9U9E5LyWvUahqqh6nW4o/AeH5o8s3PCy/EDvO9UngumleEpW
J8XQab5L2cBelWKHN4Xpqg1/kVtj/8fvuL9zhV7B0Yw6mPgS+3YQOUlttcgnh6PpdgiS9B8wsx2L
wE9PqIT22+eUScmotN9MdNQeEgpe0cnRMFClbikXU34JLMkcJ5ZJNqa7zlwrL3ystdliTYEeZkc5
G8RC0V/K+xxjy6ZUm0ENWpEAyCdHxSbrSFnlhA4dPPnUQl7WUGWtD2HcsJvyXo7vJlgZqG+6oKsf
XQRHgvWiAxnNKKlnjrAZSSqLvCQidaabOzisQE3orIeTuJjrLeLp1hE2DaOpLbAd1tcihIXVqZbL
fMNvGg4VIMSekDvCQwmuhxIj0ryBsYqR6hooh37jnYNWh1zerCVpiEw0UBFZK85JiSseWHpJ570p
DxI7XwIDjUvZk8IW4NJm1POyOYFSlXiF2Qkvq7mJKlXABSP9VbuO9ln1P2+lPLdcKk65xZiXGkoL
+1ZlyEfPqAfINsV4MYOmFnNHjoCHdTP1G+DjdyNZpuWaRr+SzAz/7yZ1dXVpKB2CSsO0YSelTIhw
vXiSnJYY2LIbS/V7FdNyEqJgcktgGNuOjQfgFIXf/wfkSZ/ZIhDycG8ds0e0pCBlHuT3F4CBWrmx
rDWxtSFRGPNpihDX9uLM00Vp2vQTYkBvKQIYR4+nemMcONHU2rsoHuEMOpgzkHzXaWQSQeAkFmIb
0UArfBjddK7uTXaexiJv8SiJrF+nZ3Kz9z3W2js8Tg6DsclxP9LXEOApt/xqhgmDHTYb+umcFKlV
8mxqwdSFVRkzc8nsg3Xou6PquQZELw/pxOIwHED+QEOdnf5Sy8EvVZzVWlArfIjH9eM1Uy6H585o
dwAdGvmXoK8y3lE0MLEee1LOR98KBG5cdBtlGRwufNAqWDyTLTixNM9Q80X1u78399dzrH65wjH2
ituSk9HrGwptneiOqtec8FA+v0hSyhNeKmeyUV6/LfvGD90DIBCPm1mhFMF3oXDYaE6sf08jTK1u
YxhtdS3moP9+7dysF5lMSnyMo738kQbE862UNOFCyDLT0G71for6RMvude9nW+Px6wb1zEoGOjcO
zXLTy0b/BZM+b5HDcb8LsYT0NPraCGGpz1Mqj3kxr0RSPdNecA2ZD01B5d4bF0F5mgrzAtYyAtEb
+TxevrWT/astOKlCdLGvuSu27cRf19NcOCPl8kexWGR8AArJiu1l5wiIqJX1TN/ND1MzGQpCNR0G
hCjolDvkq30lXQJL+Y2J7yd+dqls0yRxwb0tB7fdcDHwtew/hUOEP/O/M6Fi9L91R8cWEXik9KDn
KSuOaPHGVqqAhh1eZjPxks2+WtgAqxE43Kk+4oThmZ1mLWOr49xl7po8nrbedA+IQUD/BYHWr8Q2
ft3d2t0pXZzBv+XxyYjJv18MwrDvi9e4xLKsflQTkTG8KQrj/ScgILJCRybgYjtfT7nuNomIKB9C
mmgbFxhcJPiI2tXd1j7pVZeMBUGs/UOkLjAV1jXX8OZeQZxUtsgOPKtg+W+4oizU5BBc8jjJ8dB5
uFtzxGwt4j2MlcRDtC/LZ+sO3G6LgF5Y2pRLR7KyM/hvbggEtNjqD17y/v15qpZqPXIwXCCHHLjo
JDapkQ1FEoiWwOaUTYvZ+BfMZhdqmDg8qmrcQMARpWEga6EBu2XIhJw1gcE6+vQKoOEwPiOt1ZqS
2XwszdLPIayjpg6VUOPPgz1MbgxTvgFxWYMsFR+3p2IFdeDW4rhmxLdgSBlX2r8vV5M6zk9qE5Vn
u+RsxpktgpXHgMclNgruAoNPakj4bqIoWG2/6VOh2Up7A3n3bur94PZxfbmUV39IMhyRyOQbUQy4
BTSD8UguH5puAZDwn9b4ygSDauVBdlbJ/eRH51ksM8bIEmJgxFlQW6XG1xmesNBh4/YhlAj7vdIO
idvEA6PTIelyRXNsuP1ia0X8eBFsAkDNASPhgSV0uru2+5KiHpwkyepam4tvK9KFi+Vi+ZVuOoDW
HsscvyQEsuGbE1OgQTRnlfihOl4apJelPjTgvRO3mn5XbXKglGn31qEZGdTONQz9/Ah36F/KomSr
Mgw3k74gS35mkKj4zAC9G+ArhRdKW+CJxhK+ggH4cpHQuvWuH5YqOAFQe3vlskHKV3Hdpw1heQAJ
XlmCjNbsr03T1h2hwlXRtztlCunUCX1RLqtLqy2qN50OvfTYsOSd4LRoVnXcqBR9iyf2pRJ9+cIc
oLt5J+9RMUNviLNsK17SlWTI4NI9DmQ8K5RoGeTSD1FvJlBXlcUGEQY4lN/cIWya5bk4RUx5xQoe
jE3EH6jSLWU8I5isvpemX8T7CYjwIvqb3nY7++PPWtAg1qF0n9hAVXk7dZBNGGjLvVSFRbHGcq4u
vOLP2dQJX3SdwGUQ3TFjw3oH24Ns4abh+WSL5oS+sBZrPscmJXLLNlBhyCIWnbqlWgFt87syQSNt
cM4d0dlTascxeJNuaZyIqXp+lqPV9w9veWRcA9wMkCQV9XBjRQqhNjlSC/vcgIzqpL0bB/jYYc0K
X8wrU49SZNSKnJwlIy+0vS/60gjw3l5FWtrUIYpVO2ctHosQ72FrgQxI5AhJ6nED8MB3hFD2VqXu
EDyHRPj2WebTBjLDgvahcIV5cLqc1YO0RhCJBf+t72+3+/Bs20xceLTVjZCbldnkmq75m3/Er/fE
m/1foeO5WfmeVSgREG1jzyK0jikYE/DTTRf6Q/VckYWBdvHnUpENGDF7v/EJqYnpcIT1FMqYi/FC
tlhdKXtxezISRdaoCIf7TtqXimh76YJC2wU8e7dO6J0j1HkoDldp5zyGmjOdqUKv5BCMQ+wMTiS/
5mUYGUVoKHJZoAgJTJRybYOoibDvvnH/s30habxlH6DPN1if2EAJleOIzNgIAmFtTEd/zHddlkzR
16zZ9PfBxqRdKnXUf1UUw+S2/6tkBZ4wFHR+kiwmrPnR+SX5ArQwaIec0Tw5J7xXHHPnkMh+SDvs
nF7Ezr23xoMC7VPZ3NfJfpayHC373xb/b5JqnrRPwSn5afx6GBw1DATeexCHvdt94EvvYNzEai98
mzfDd4BWIp/nuMzFTuDovvvucqg0h/4qctfOCSwaCCpUPjUaeyUQFgw3DYWkG28efaVY7egJwSo7
KuYt2+t0/l69K0dOE9yyAYsN7YxgRtXjDkiwV4RqT8ajiumcmq57JlpiVuNjXcgF8bcyMYE73d/p
9lyjw8kRaxrFZinpDtD9abyL+nvigzS7uyQEiOdAhDu4nb9oaq1Lo4Bc1y0qr1PgSkkNvEGet0xz
j6emYFJEYMroH/188lDf476YFWHoflwRV/APa9EjMGQwoix99Jv3XUjopRgGr8rRUQEfaQHko2pq
NpAndatYx/cITcA+bct20a+L2RaNpGTUEY2Xzpe337LicrM0Crw6XHDhIpw6ALWoA9lzrAEgEWns
3cXKAJceIYh2DHKWBE8LV5kgVzircwGLtILTIm5vD+KWUHtZ4Xbrt+YrY3bFOTEGklcjBeNK6kKv
cm3XjkeUh9mPLatCrtc3tuFCaJXdfRGtp+tckdoTR2W5yIz95noEsDZH/OEv7kwiIBAbcVkz3U7P
bNfeN37/PQhMlMFRgvU7plIUdRNZe7poDRDnp3xajumHKFp+9HdmGl7EB3zH+Hw+bzvPY3ECsXnd
NpsSfVibxupuKi780bX1ZaLOX/pHxtx+QYrxfvAcIPyj0n0Co3usT2jmuC7BfExhwvQadEjmzLgg
QGBohKjfYO27NGj5xrhQspG9J/Cx0CnH06KoX7Hrzs7q4u2jPKLMVacIDXJY7UYd0ElINa7vqO28
idKm2ivChfe+4LWK5FF3qP2xKJt2/Ro8KJgdu6S7Ng7u4usnRBxBo9kyhff8lE15LZce/32mSdYh
v0Xwl1yTSmAk6mvEd/nhOp3nTkS+2SYoCR0Pzx4iFHQybL2iIVogVzV2PndyxbGh5utk5N3AGz0y
kDAvHA51rjdH+VpnhchzN2uXAgUtHltVJPvjvietD3kuY9IFH4AzxsE6eezCPFq8RxuOfQYeUURt
rwRThJguMhXlIuemb95+8t8U26QE7/htt5T8TNmTEJnDqNPZZ73WZCASV3MJcbCwZSeyC2JU6rAX
wS9RTvBE9Ru8U2FC6wq8T86O6mZbZK1CqAUQQY0lus6u2EJEAGTNL9CxUP7LVsoGpF6F8yY32roi
aG6eggT9xPpEjG1M1unsGKvl2boRtqgGnty+9kRP118LTYb9A65ub5JyqmSVC0SeAdc61droL/8R
d/RhO9MGnf29DvcL4b44eTsu2Scmo7O7Fs4ijSkE68IrONHvPe9cVUU8zWs94sYkaBYF9aYdMX7N
wIq+No6cwkrjyYJOl6t0Jzsou4reuhcezn596viifG99vq2DO/ISai0wTM4MWyUXyj2HJm72btOF
8FX5NB70wWRMfwc41vQZykfPtWiLBWmupeZd+tCD2x//YrgSWHjluZE3XpsxZG3rltyrt0vkKNlc
2I+2ZPTGXHl6wRka6mRwznp3GsaXDYCMXrpwumrJMN6+EiPZzPtw2XhavAR9RwqFx3vKJX2CpMMT
2e4+znZ+452J+ljM2IssjvoiTOmw1rplLs/pyms7j8UtmP3K9vxVjTFDv2JQAA4ZcvWLrsSPC5xj
qIvrEGTjkF4tTVVoH9bDzi4s58Qr0df6h9IC0vCDn3lCgdnYBG5zn1b8KpbGCRNniF5uIK4/5A8L
uVAsCSXY93GIZQnCg2wn7ZOa23MuLzF6z6T3geV2uq7IG7cRI7tCt1Mtn3nydWu+8hAVrG4hTgto
NLdDUxJROOV6x1o2X8YO+aIZVCtVWGKyWTFbyCF5TJXoM6y1sKy46YjaOH0uVUGCcLg17tDvsWAP
NtS1hq/BwWt1p1Nu+nHbrfiGeFfZvACpO4KYRcV3IXrcssPtIoeMp012Ymg81e94eKaOfdf3f0Zl
ncxbFCNH3Arg/AkUaWLWE3E0WsbB2myIo+mdigUh1mWpFzoEG7dBCYTpNSfr3kqM99vWlPNBD61w
9D6b2DDO++4AojMjiDfKqHKcp4J15FtipW/ha5o5YjAKVYkzDul66IIpg4vRb4w0bjM9susG6AB+
LKXaMuxMAunrDO4L17TADWQLKX08zejtIwdF30mvS1/31ePF9xVCf6qmqj1oXJOMiUnlD9i7UFU8
qzwM4sWcIehGC4Y6NjD2y3xM3AxHp7rVKhUAZ2DOYptUWNYTfRK+CGeKM09aWY04RZtTBxcCBzIJ
ntrVQNypYlcSIdQdPbl03zfmy40NI3gJ7Pkv26AuLCA0sdAiLMoKOmJnqcsHY6/l98cr2NVQKHQ1
G8z1gHr+xIo6I/XYPEOZs5bKmKh3GrBZT09ZOwUiKjE/B7BLOWh5YG4y3vWZVz47JB6kx9jGvN2j
0nWD8BhWWsYzWNRL0usmUzd4DrLtHaHF+nKs09BMCaRhSNONJinYZ011eHGffeTHIjpf/7ngxHAn
uTF4Q00oN64Iwm/Bp2N65yR8CQREXNwvGYn41rIylnncgiBV0r4atHpMOg9MS64jp9Cah8Pf6Yod
8MlWkMtR8z5m9tSXBPaoA30R0305LjrvD0d6LbijKwJwERyBsrFWBfWqxEcdQhLYpa0TCxAQ2So/
qGeSaJwORCPpeJdsPAbJe79LaaVmhhBJaMPLdfL3OFoL2/3M5KtsbT4vwnf2/eN5wwgjQPbMEVwG
KE/IoF6j7+xTFK3BlV6S3s8OH9AtOXbv7h7R2h/floc9cusfO2NjJZqtpu7MWEZZyDB3qBqacgVx
NpZPIFD0FMJFvwCky21Hovr/qJZmVC027H9AB2h+z8EGma+dlvhCwqanoKDkArClf/yRKuGyHcij
7s2oKY8Xo9CUfCygfeOEMEY5Ph8Xt2ZDk+QL2O+eL2PhVVa4jmDkKc3dMVpEG1XF0BdlzIMPklw4
Nov09anw6Hj4q4mNhucFKjlTw1HM/luM3wQ3mMx4xCc7coloIQn3LknNqCYWfnGjtJ6UNqezUJEQ
gA35vf7KNHQ4cCKov0bwTQllTE3d77RYcYndyuzmi+biK2gv+Q6zDSqacCnZRd6hCRUmThqoaZCJ
AUkCd7H0e+IbJv5te/Yrjer5J02MCtX6vSzKx2opMgsNq0rMC8wnK0gct3pjWurLPcICnp51xHOG
AOR3zt/rgo0tWgUjQ52Hz1wzTT1s1OE50kQ9bLGHmvYKhYwWj3DIk4glmc9k+fQVbiM+WHDxh9+Z
kiKktuEEUyLnXGAXiMnfn7Jcj4L3uyCB/NVjLvnQLqvF80Teoaef8OpzT/MM9Ykt0NOgcsMluVMB
Z7tfelYwnaDBryYQvE5KMLMGqMe62DFJ2dtnJclqnCAsKBRTCQtniQ/lkwh3RxqG5VDGl197++6Z
ffYj/z/bKFMdB2KDetGPqQ2Jy5KByfY2koznWhH5aOobjINQVwJZf5sh2gaA6lCwodkY/ppWcSEO
IIPtAXnKechTaJp6AjndxQryFEnpVmUsSbpwoM8ouIH8tin2De9biqwlkwuRRR0UbC/C2GYg4fEs
DAYTI3hjA39a7DKU+TqXUzX/ZaHLzmxUvvQQNCCDZQl1S93XXAXJanU2SzpAL2a3qpM+3IjQkD5E
lAAujU1IhdiFMHQMMRoowJ/CLH1c4VMIAL7fEgvzSUT+/gWt4kGvAuGn7OZs/mmD/GfCJkgS9LAW
12gvMRhQXIkAv18haBqztuM5WIEKnSQ8lM2sDphYeWrPUaN63us5zTpaoICr3nH0zMFmXH2flF2q
MtVMmSSeJcZt93Qu+WG/XuaiSxU7fAiJIfmAeKUAwWutyIBjc3udToCI6oUiPa/nVQwi+39PHfTG
jQXSAfMRJYA76+sJAIrGSGr49ZD/9xAViMiuHtxPEs31iay5PZbshQRuHFCsi+0CHu5GSDJdSCnC
ljRZfx6YsoUh6FIZSchDcnQNcm5PhxC7JTO7LPxRup1XOe/VKo6Jr3Z+HsCY5L1gEKh4fsbjkBOm
oRYCwFuS+JfHa8n3eihE/EReIeKn2/vVmPsc551yUhT+/O+DrRxFy+THJj2xG1BlLxxXH8gkbuHV
nVO+rK32WEOZ+Gmmntw8DDgshf1XZOC2w1ZowId5lmoMkRO4AN9AsipDvwnWL4VMx0i6RZ29VsGl
zCHzYS6osDddMtGmF6062AZhFsFmiRKASXiaPM7O5aJwt9EYTNiLV1UYgAv4saWUzvnhgAmCq8Lw
ShuCTu4SEGKofmzgIen0VV8IJ84yNq2a9jWGMbqsn79fNi4Y6spLOJS5W2l+stcVkRwXPUghkIOJ
omCaNzHjLVzb8BO03z1RRzOWOh/SnOyYuDhyb3p/5V+TbiUIHA8xdNJWt7Dx+Y6wvv9N4QRvlOYp
3JTWpCNgEeBdCDgRIea0blMxwoaoOIgr8XnTgJak+h/+d7Hf0iFflUFLpq/hIGgOdkN1qiAcF4pe
XOII9eMqvekFMOqGYuzrbCW8GVNHt7i/23zQhwHZO+QFiSvpNYjetzc5AvtNS5vjzpNBsQ4SOY5g
sPpiUr9OIn99FPdm7NeoZDihYsYarN/YQRvoDCgNG7stLc0QId7EjmkJspkBUypgnu6/ku/q2sZm
yFyxVmAH6nvfF01dpGsyt94uFqS4WhnU248XoNCm6ya/21cHEMaMquTpRB7JikZztt2h0RWhTTFE
oi2QniOBypQ3ls0xDolWOnQYa9GGg831dE2gPw67pHx3ctkPyE5yVpA6vBoNk/DKvMPKHLyRaiF8
TKqiVtjqKWbYRaql9acISzC02tYL218b+GGFwXth2v+QvtqHXi1OjyhbFp800FVHeLGALL4kDoes
6m2ZTUcE9buJPxXr3z1tZX++VkkLaMwcy19nANkwIuWtYmQySZz7DDMfygrjV/PCkVA9w6CYy5+q
bPWtjY+jiuo3EXFfBz0SS+YVHY7jl+3zhca+N3rnYM3fCWb37S7Ak53Yye3eLT7EmcpQ7DiyB8DH
txaVjJQWsVVXnYBtWJXqH+bbMvsQrRxWhoedLP/gdao/k5U1rq/xUQ6rYivpaHPJM54JN/qETo80
xfKV62ud/JhnWRYplrt050YxVi2ixfF6T9tAkcgWH7wXMQYaD4G0j4e82TRT5oM673lXR7iiuVbc
IsKBHBkM3inqACiss7rThNh6XLu+PLTgwqFPOXxq48saxkEywnU3vh9tY+tsDagtknGukB/biMrx
8sPqslpyhHTsPRWY59aEu1ZqkwNhlP8QIUcEiQHmq/VmFEYX559OMR38NxX8JrzR08OOmp4Iryze
yblIX1Z4vfCPxd3EOeR86caBpzbUNhnRTq9oWBaA1vsUgL3O44hduoTjiQAr53dETGeiiBRSwLP6
+d7X0CHGe6bkMG2R9cNe64LljwLO/2D12hIskCf8RWlrYYEKMYYeVb3XzPlhRsXGRLgADWA55iPB
p+SA1H/lRhbb/ZwFyTXevMqfPNNjH+3pxY7DN44/tzwps9BzeakMc4yQ/0FecXTJIRcYuA7UQfXk
TfKy+8wHhVgEqMQUAuHceEv20ouObK0KIx47lQD5P+1ZMnI2Vyw+i6BIspf8JuZLya/WfjL6QIWJ
a92BrsHlATgW+iF1TyIyprP6mQJPew26Ce2b18uLELHlPKNb+m55j3kUPjtQ3RtgHswh88phn2+M
E5VosB4Dk5tp//INQp2Ocwyt6p3E+gchthCt4bJ7SF0Hek1bna7lk8AxQCS0zKaGwRbb/pK/dy3+
oB3KjoM3QBqjKi+0hM6xRKnliGlKqgBotwmY/9HCrRZjvPP3TTAu3I3c4KhiUDwHexMc0oXMc/bn
50rd6ymJ3A5AnaN2elyXpH7ye0sdVp68lEBZ0xx+uiDaOa6Q2lQxgyhI8IL+cO9g1/u+1JvsggbJ
/18E/ROri3+uOKnFhv9/XsfKQ3TMtpP/FGeShHvr+h4FYFnthRiWOlWHK/gkDXLT8q4U4mON0aul
yPFNQQgEDZJq91qJlHAxbqDx1+YeZySrdBfgS1rTtkj9nlolauEyPNbgQpmFzgr437IAFMDBi5Ek
id1sqMD7s7xE1GyhQzc/GAbrMP96X/HyFIKhP0SH7qPxywppdmK8fG+IqhnEKMUwLCccsoOv0zKk
nl4rcek48XaFq4aJNFSqNcJv7rAu4NzcomhQy0vTdJzXzGHQ0/ypoc6m6n/mv+z+cDnWDZtJSD5K
awRLUUexH9fFyp9N7OoLetRiQ7SqSEFDxRh5cb+WQ/QVX/VqV6Nlr3b0SnnjR8gKRNiO9mZmOe7A
O5P1vL+Y11i532/J1erTV5F0D4XbQNrSug1egc+gDjni2r0ggO/IfSV1f3W2Cw4we938MY/KDKtR
73y5FhEZigIaS05tTImjghSzuJ1cKDYHHWzFWk+a1niw/PbkEbyzFySqhLd6ZsXnRMY/E+XGSemF
KR8UEXFdkgF50eUGCxjYL3YermXVwVL/O2opAzJbqI0EVDrNZ4NXCUC05DRmdmuiDBtgQJJk8FC2
rfvD1jFfSz7QRQExg+GwSQ7mIngh+cTmXEdTjYEujMWK3CO+DtFLlik3DoIG4gChhM3g+qQQul8d
jR7j4LnmHjNOJSiWWwuo6eQz0hhuTR6E7dEeBfMvJCfDrqFOuSj04dhc3V/fBT5OBhqOadXslzWx
lMDtkC/uI2e97ygHsuw9K9X2m6k/oT+0g1KbVv7Jxuhr9ZruI56DQE6AruPKXwlDl4CZdsircHq5
fLHIaN/HO0YizRKqFJo1tz8dEVLK0NCaqpUsmuaVDcLTUIfeK1Fm8IP+tSTElPqVs9x42vXGfuMh
zOl6j8ze5R1REcNSntR43zRX5UZdsUFeZprEAjsAYK6A8CdZv5kMmSgT2yOxDDMJsQexGlnzydvN
TXH5np65JqFDSVqm/RYKFsY+Ct+P4ZXl5JwPXpmwWLEp5ZOK3JWn1jsuPKykw1DuimVec0ndTkhy
M5HMVG3fvPK3hPJu4/iNba1EW630cd5/77IWZ6Th5ifr8TujWyTJNvgYucnq1ebeAcccxF1qy2GZ
jZGYIywIgFPozh/TUDhbahhWzo22FKtl5nIT5Vy+eWHe6Srvporc6srf4iaoMOMPEetuav/17sbR
+1zb8uG2R7YLy444oNBBxCigW1v4vU7d5rwtqO6sSJA4Zv6RtU3n+RAxwMYOMGdUtiL4v6DYtuFG
JnXOArMDCsc6J/SUH8YQPRC8MbTBJyuqrDUSpzaMYQiWiQi6N/JWsSD3AHtuqa/oFOflWMLtHsUg
Ps9Dm4ynDtZnCi4vGTZByYlgMDN5hhF0bcKHhJ3/oHSXTP5lRka+DzT6UF138tr9Z+AhkQB2QUEK
PiTMJWWvS29T/5vuXPLdMT61aCGYfGPWJWv0cpe5WsAgwv2Ssi6rqLIdUc1FxsGzrnaqeUtIZAW/
iivHA/SWV6co7uGso5vIc7ruvXM2420WV4/uEIJNVxsg/w0YFQghB2D4OqHJ59sbJtiqKaOBREaY
/NSWMrOCTNdtO8ok3O8BIA/xfcYSTsP1GGOG2WWevkt1SN1S3aZmilLGzIY/6/P8Mc403+G9PtMV
f+V0tmL4LluSPi9ZSbERUY7mstbIp6NCcMqREbkn4otPTPymhGb7AoMR+ZppB0OxqTeTiqGx/rex
fJrpkp9PMhgHQCsVnBRS6Kl8lCesqRPVYPXUsYMrss5T15LPpspttiBLjdmi0+6kceCrB9OcF9IU
OXRYfkL37hpTvzC52k1DVCm3ZEwOyKkANZTV45urcXGykIJBEiOb/nF3TFa+BndBdCcZmg5vgPvB
OcV+2Lsmo7w6BvdpGCuzeZ8rbWkCzOIMi8f6kgA9zXu17gdr1idFtx5239oURFI5jzlVQUuXZpD5
NTC7FRYbRad2okA3yEer8PUTqSw+L8DZK2mZsIjfKKIJhzKNUioMlhOnFzbb5TwW5DXmd8JeTHwF
sjfCiAGeEBEtxnSblGIzCC81hUNa4up4rU3d+0UDFvoL8cAyIlHqlrr0sjwMj4BHdPeQAVm4EYdz
MXngCT0TdMkMJwAmsw1uJ/BcbWSKxRRf3ffR8nW/EOAlJzuMjfQz7atrrJmTdVfMOJcaOvxVmYZd
dy+Zt+ex/rIolvsm7qf4B4Ka2DVHouQn3vM4MtajwDobsaywPD1DneAkdciDYk1iKcOW0UJ7yQFK
EQ28p5u7NU2qER2pO6BwTSryJ4TWcced6FUAqXYAo4/C5WVnpdfJhJdIJX9np4HS0r/jURh6QY6U
Lw4mLPHD1cDwGBInhwQpUk75PLbxUMKyVWS8pvLy4whzQS3JpoagNW11FXy/WRs2We6tVlij4fUB
7T083TjBAgvxZGGmlGl39/bunySMaUnCyRSRhzfKyC0mnsfbqbuyHDsf5LLlu1anr7dog0qijh2s
o3kCVdng4c9j6ceLp2n334B65b/2kaklAcWC3stQunROATorOWY+oQnByKPY6Sd0ZY87A86EYBkq
glUUTaVvT68xEZdOMj4VO0rggI0tqbIVUzu6NX11XCiHam22Eg9SIExvOAGAKgnqzEqJcwF+b+5L
zcSR9nt8y9UFeA11HeriXnW49qpjESdLM0iITjhf3G9X+uCvgLTuUxG8f3DiNmEsleUG/pGo7+Kp
BEPkAw5CwNLb8vZtR4zoSHhxKQyyLBG1wjbgduJOTXuNt/9YGArEtn7Y7caLoFhoKpMKwtnLMftU
ZjK+AwJSjZi6ePgYTlA9qpfHdcHIlBUoa9MWmAmmjupg+Qu2IHade4WJp2sLbTTHVIv0jKO+TMdP
fGzyS6uviOyklYASvnUZSUVUlH6HpWNNnZmyB/dP9t57k3mDCyslZAwBgnDmXQXKcXEfuczKI9nR
bpuk4Lk5yK6ebsGcqYTgTuhaJcGeXR3Rg4qx/gpJl6CMLLXhBY3DG5Rzwe3a2dYWfeFIJ24yENdy
fCZKrB3BlEhE9XeU03M7sZt5PjtnMocTdZRsC5IeTxTQLQJZFrBOL/mck7xUmT/rtEpzRaKc1i3H
bXxuAHMCdXkkRH41cfx++sMiMvUXesflTobkIxc18EdHrnor3Z1CACgeBGbQO4eLfTqRbIh2jMOa
LXLmaE58gpMkkICEs/sPop0XPrCAnHHMWcvlk8orCZ0nQWP4QWgazqPvYq6HWG9e0g4x5q6zgLZY
NzTRKKjCck5KE2ihQIdlCCsLcaNvrvXoRm1x+SVj3jWIDoVh3dCDfp7fcuAN5lTcKDlw3E7wdhfT
ZNTHmyIJ0yyfSs/1EGbJRThvx0LQTIBmCbgX4G17YBjf4GkT1hHolAGYw5WaiAG18GJHznZTPFB4
lKywuUNnaWBDIjT/n5zDu5pGxczPw+9UyVE6lPP+HPARLpg517rgrgc3Mg2PcSP6fzl1pVUKI1P6
dtKw06YP6mwEOmL/OEICkDiIlxHTUHMLHelaWk4KSDrXvhmhpSilA7Ko01NY5dx15TCwYGPti/1P
5m9Tni50QteQNKg8AInHThsj1aeGFx7GXehr55dav7HHfuypSSJ8mj0maSYBdD0Y4/8ShS2uAKqQ
Up0ElKixtPqP+wdvr5Q7sMFGoccyWPY9GUoyB0u8vqbFxigGAsyBzbRSp//jy0Xzil5r9wVsdAiS
6dSYVbvjM5GJF13+lNRn0CPToSnnjsBDZnP+rzFfUHXIihW5aLFawvPqPtdyDTDIGDR5IZATmjNp
z34i2TFnf+xvVhor4EH7YLuSzYiXZdpabvW78rDfUbtqNm1Mf5TlbifULJjHmiGJP2JVgdSM2dlu
kjDG7MD1MsbOaLXFGxjNPRVWYfbPdGINVLHhh5JjvTT8yJAohxZ+fQ1fGKurigyHhhuH48oRBSSl
+fsr0r4W1oTt64ne3IlTlfY8tcilm+0Zm55/Yjhg726cu4YoX5nj7zDEKMG77UbJ3vxX6byt5b9J
xkff5TEWvZEtskfsn9SUqFEAy7vN6R9aDOeNIcIhlpsIixgjLTxP9sWcszNpfVJx9kM+pqTNxbVg
zkARnz05k4VsW7x1idUFeTYGJecC8y89WlbsOeJcG1NRL1qp+ILHYnmR8pZNupgjdoCouaLvzst/
BbzK1ZOOiiZ8+0bSm7C3NeI3jAVvWYU94h8nMiORYl/+NjJ8z8aRKOAv1r8DVVphcXE06YrlOUrB
e4XG2WVGpZn3MDEZVM4AcKV4E4mBsXsgaXLZ2H9eMJv3QqFsSTjGQHZce0YIP0kI1ZimLQuY1yIE
SJUSKJ+lq8YcTY+6DWZhUGrROP9FQDtCZqugywL3CraQpyq5QX1DNGLJKrhqB8PDdVsOs+8NX1xj
LSjcwsg3Lp/qiztSq/yI4I74gRpj1g93V+5rDxbjiLVN7I0iFb4W0PMBntQWENQOLWUag4g7/2HO
Vpj4vFBGw2o3QXVkqjGDhtQhgVruvEafFScoc3nvLWPmjqxuXd4h7bgLV0+0ruhHaNu7uIGrYrQc
mrDqW4HzeRBb6Wk3VV0+1sRxJ5akXyMKSu3ZnlWJUl1uOnkrFb2k+zF9gFmQOKR6ttWCkuWuqtHY
+8LJMJj6v/aeYZFdEbbszEIVvI0z9OHfHYIf5JaL2sEnPFtauuTWUsQSFmqy/1RXtb8KPtsp5End
3uQvFsZBQ45KpfrOmNQKXdfwKCDSXyljH/YxgCMB7bOSk3GgkQuAA6CqcasUCAtD9XHqO5/76P2c
0QEi0Nvc9ENZ/1BanY/1OIulybf0oYE8RIJKW/63z0NNPzY+ww6WcNz2HO52WFEM96Wr476J2F6h
c/fjJci1qvK2yLEdBy19wSsBkPyioUA0is7obF1GTV588S3rY9bjUhm1Jy+y3IXdgCdJ0FdDGwVm
TgYhj5Eaga3JB85DEQHkTyb3yXQYT/4U4A8m67iNaDrtgaio0r43Jz4rTc47HRe1weCCY/sbmpRB
hp3vcA1Hl5tLJ7WhNqKe/DYPRUD1PEsrCc97eiEtfDLG/9ZQvN0RQtc9E62+hZ2FVJcBSw60fdai
STNVPjxQi2Mxv4bBZEfBGmJX9+AYmiENcT2dkW/Vw7V8y/nq2vBuoPlOjPG6T1pb6xzHh3KC4KDb
NoY2H/fbvgVuDtiiWE/u74pZe3RbD1TnuU8d/76p/01GT7KZT8qftqS84FnGISSRsxLN1XC91xLQ
0qE7CMWDWeXDYeNdytA3gfYbzkfE0SNs7rtE4hmOVaoXmuZuVabCDXilEmrb873H8VBYgX7g9bSL
isL8/BQTfF82plw7i8FJ8I2k9R73yxlJ2975b3rOv9Ut4GvEqdvLIsDtgF1+vauHmeXN3544YDNa
ZUn2l7LJIkaDZ/T9NzY8soYTOu09ouHz8XlP6JvMEzmzJ9qi7vzDY/0Xc3bfS1HPmdXGru6OjaS/
RHC09tUBNoHmR4V5ajG6LtK3FmWRd76YhHl+Mxr4XmzY3D576oCQE1Er3XJ6pD/iQ17e7kmplMt4
T4LYBahNf8eFWwyX0Up9tqx3UGhJLvxQMFT0PXhAQGzLKhIhPBWGy0AtighHnJuQ5vDV8frWefHM
sV/Sg3YPZJvcy9vChJ8M8F5HLU3eN7HmIn69n8CTcby/Er3BePWvBPmGAfeR9/82s4wh7f32+plf
VXXTyjRC8/jLBIkSSdQeSWGiAWtHrwGUyhG+VYR/Tzfssn2ToOQzp5vJwcUsgAiEDpnCMKN4Duq+
O/jFuiWHwgUB/HQHYqUMxjp2BaHfkkBJqiqUMCtbqdnBGjGX6XwhhUNMdB/PFAeol3qBdX0m5eGx
cwV+5wVyVHzplTksawNlplDWsm+RvJIoWDnVDsA+eiox9pTjcDDRfcz050oXRUjKosM0C38O/SRp
8yKlqyUNGkeK9Iy3w8NsFkBkzL+XDSmS9nUlCV7W0XcVnbJ6s7N4yOtkitbhjzNstkk9LECp0nw+
XQTJgcEM/L79++SVIBkerY+Ie2Eg2mDGGSwbnBnq5z4rRDYv36J6ckqBUk3xgdIgaGyb3bwTLiUU
zyWazSAgFh1X9AcY6EuFVRc1xB5DsUvzTffVyKJFAklntehaPShk/GaTqBFJY5isjvRbEuSv3Xe1
n3SNl1/yVf0artH8aCMz6z1s0Aoh1iMJWBDIjIIyrQhiWqVda5CpE8WdDKqPpV9yrmXmhJw9ekUS
hdNCPR/Cjr2tEtLX80LxPazAtl5Nsj5YuqNBDXor5+VSQ1gQV2ibUAQoVOWvslcuIcTCmALPJrnZ
255J/8CVzbESh77V5ilPULwHqlBeqU6eakxqvr4Z/LIqSfuedEEv2zImPpnNFH70cxTT8a/V1wY0
rx6+inPWRESZtqz9E+OY/QKBvME86RurM++qm4ckJ9FwDd+urDO00/yTtn3gQH/Vcc30KmmmTvt1
+UAIwImO3VwyK6lf++AvUif+rXGhSXEPn68ke1kplso3CyfBvFSHwtiqkQ1Hir+ouA3kLTJM6Z7v
LTB5BXRw0LdGhOnrHsEi/AoftGNkOI/KV+pVnoCVJ25gJ/FZ7mbO0CFN+vmC1qn4VKcwEIss83gz
lawp8wzFaLGy2Dzj6LuyW4Z+sYxYODb0IuEXUDB7GJxiPkkUFsM4xzRjudHCPbl3FO12bcNtvAPV
Zl418sUacRn5T5sonL4uSAvQR007PyQZfuCCn6ysM925k5UhDJIhpYpF6M/Sik2h2q3ztdvjeRB6
BK9HBH5okGyuOp3juQ8HDqcQU82QONePt04IZda+XVkQ5wMeG3WoydWwMhpLZ3vxwLkWbZDystrj
M5oFIbKdmHPLFUyzhHKc0MZD31OvQnNG2+SzpsFiqbQT4C7rJahDMldgTSJw/S3AeXt2819IFGKK
z+nH/69NRdbylNmWTKvctUcdZow9ZujUWej5l0Ih/fVa//BZyYOzKNThCvgQJ7Qih4LBDolMJw9t
CxsHfolFs2BNHb5c3O9ljkE3D/+GJDGYRg66GTNi9eIwGs4hO+acfpdqBjM8S/ftGPDG4Gqktjf9
RIIO2n2pz5KUq7KLKbpxBXcCc2BsIw9uVqzsmtmctp0hz62GT7CkXyv3V5xI2TGGYhtmtW+kksnj
Hsaa3SoZwNgP4lfkHZLQwFlT56lvcA6d5wrL667MkMaWDWDF2QQFcWh9cUybFqOgNcdqdCRtZGew
i6PYWZ48xk6hogX1Cieo9MOCH7TY8TCQOUba9qB9U2HlEcjZ1v3mmHRQhBgxg1ojTLELRtMOfRig
Iq0e/XhcBltUGtEtv/kUwzicvsWvEWQx5FSj1PYK+U7y1aeEDdOcJOiGWLx5aTYooFUB+OgXVC2R
YP5kbz2zRN9UK/UsfILEyVJp3Mdxp/h7XUNyPtxwJO7p1g+ZAPvqX7ehf6WdiN1Db8Yosm4vHf2J
OdrpjejLiXQ1pdCrt4KbeySHGcwHIl3zEckbHPcZWHAXw0dNCRz6QM18u2L/6njpcCbIV7GSBPNF
zlPNW3I0glKVK33Jqdg5OlPE0+E90noahaJ8m+lWSk8YTItBZjvNauutPX7g5FbLKDtCDT/j24uH
vjAT+pAG3wLT91TuqzvvmxIpOT41hkXUve/ZF+BfsKYYAi5f4Fq7fDmWcuuw4xFkutrSmBzqHk+0
aOCmrnDUVwpOYpzNelqEd3qAjrIiWcB1RSxmq5JfD2aIFBHpAUPwwL409zCh4muCdLJ6ggDNPvON
5XgYeAVqiKYPWuaUFDEmKozB7dTwr+yI/GBJWGFqbxV03OohFLk7lg491g+u1ivEpGPs5HbAP63I
zvh5dS4pGKYegoUUNE0tcvC6mw4wwxYVaRoDb/4UDtQNPVkY8vnmGhU/S2C78dn86qQoTR2Hzrnz
mBhB5P3ie3xN0JKh4i1KsO+rgzdn4FSmiLr6ARsz/DnSLuwwaEZKM091jQUDFjZvwupS7O39jRsw
rI+9EBTqXGeKVfVqIoU2pObWNyekz1IflCpfaGyqUlv/Y9e/fgq053pkgNPbDiE3GtLxgbLtRAd5
xpLI2/UVhAipGSg3KrUFm2VjTu4jvN1xmDHGElLfDMxphNFcH9NTXv+VYjGrYig76DiM9m+GVsIq
u+OgMqMigByb55KmJZzOaOz1RRRkkqQT5BCc4eb9MnWsoSzdquofsR1TqnVRjxsoaf5BY53P/7S9
YoinevrRGr63x/RN/SsmLSJoEv4TArKCFQJK5IL+KxQScGz05y3JDejhyREWiXnqtibb0sxUH4KN
1JM4K9WHsH9R81bxynN31OvkFpbVwAYuHHgKGzGDGns5JG386W6SZB6phlY6gmeVxIDm4yOVuygd
ktc2OAVaFaK4N/Oj8FyUODU5nm2Av3FWbGMrhsIOC1pOhINy2mDC4yoyC08tmlMvDvs6hV7U98jt
bCfVVRgMNGDMpSGYoBwYmDAgXpZrqARC8o9JgA0SwjT9RLc9nDbA/eOOq0jgHfkDlr7rKkPxPptJ
KHHYk5/hqRCI9hMuc/VZui/iNI9OXEaflCebd5XB1fxYwSGK4acJTsWx3p5J5RvUMH0/KFBPMFnz
IH0toR+5bERnzMDKSCHjO6CvVZcFErl4fXqFoJFxCxodvjwjDgyyQkEnmdhJnd6Mp7ZyAvQGXYD6
E00iOoKMUwXt/07PXwS+zSjU0jfxB0IqUl2HoFGfo6EoL3/gq8LUGPQTkhDEGnMSKte3oqFQNSxY
YmaPgvdaa7COe/dyUoGT63lcDsuxrHsZ7TH+1VJtbsV6IysUuglefLJ2qfLcE7SAXLDkdvkgwuRC
J7iJ0o4BUU7WsiO1bItre0c5VkioKllSpIe+vZ+T4SPq2MeNvmqGbXNdbYfclA3bhDTQD5LCB/Lb
/lFDC+O0NajJOyM2WWgzhjzxitlZHfpeUXxPMVJe3yMDmLineznDXmlNGLa5MHehtk4rYVLw60CB
OfHhrPolETIcHdDU9pWCH1F0MReAj6XuZQnbQnA0iFWc4BD8MrvDGNJbJvLpBaeT2BACYbOKFxvx
QIsOLWNMhHNxRaWtGNTAp19jFTeD/sSLvum7ivnurdnUpHuG9HVH3ozEBG8fRr1EFSf4G3HJ2QEM
NRajR2pExCGnqIUXCAxVc6uE5tT5IxNOc5RXCpQfzw/Eqz51H8BkW/ap/y0D9ykdbiQy/lEI9VRV
H+7Mu2WqR/bpfh+Nv+x68fUEECE3tPipAL5vDCxhqaexHJY3QszDb1dehiycCTVdmvnFQ11vIPOO
M/OkD0y/OrPeoNItl00n8uqzPi15PKQFVaQZMPhyJBpB3bR4MswHCujWJwc+YNQ0tRE2hDwWzbu0
8N4BAxrVVL0e31qOxjNTr2anLzVTT8kjmQ8j3sjWywymDECLIDe/9sE8810BqNe+39qcrcYyZ8W9
4I7UPXjx9GwsEISKg0ErJiPYIsxl+cwRBR+++YxnTs/w6ytDh3Gu/3UaY3aeGMkWLL1WGvBg7lpp
ONl5AsqZWSmpcNU92QV6dDuyg6llI5qy7VmNmKqej9j8Orh5iApQ8lN2smqbD7f8qihxO31uNQyT
UgvxfWxZQqszEpOZDw93Q5s22+v/hD2mX7GSST4UnjRhGhViQt6jq4FaV5vea1Vrh1IDfEJcHkfY
quWhE3YjJSWGPwE7X9WGHwkmBfztqNcJD8GZLPmyPcya1W0BduyQk6R5+7G2WiJnKGv8jeToaq4s
nind9CVtjSBlz89iZQdpju5ej3TS5PR87YLjkrPfX+D1NjSO69QcxY+n5SofhMwHuqm4riRK8+bX
uNp+VMJ7evIxHw7eEJr+qYZ2OwmIKzBpyEvJbSY+m5yTLTZNxcUmW8nlOWBFD25/a+G50SnKK1KK
2fkU4y7czlSs9oijBWpLRkB0DMu2GJ9LzRi6JUt+TwCUoGBA9RZNky9hRh9Sr1vnSAz0PpGUosJt
UOYRWjMWRUBaWVBNmb8LfxCEk4EtaG+3eiGNLOQGP60ZK7s6+utogZG1UOYZdLKooUIvJ4fCa/lC
f2ZM3+EHXLLLHLsAYmyDnTVzqF5W0Nv+pC57JbxyDlDotp3x63sc7PlZLaHThzg/ECIampJhoEBA
KPCzpU8JQluPUohXpMBAFZuA6Ata1bHVkJctrUPP6pDTuf9NgKLGsncamsZ/aDLnY4gszZNClwIK
GNY4cGCUopcqRZr3g+WCqxqow9fflnM27P2pyv8ZrXWX63JKGsH6xs6x0gZNV+qDWLWxeCPaM9Qz
B+UfGDImoROgVFDYgeWnRN6wrGJrUQVIJ0xJrbIttq10U9mt7OR1n8GySuKtxOXlQQEpubBF5RnR
6+5lfi0Drg9xlMdXPa/12ZMbYQ60a4UttlXtQPTvELlMoYKC+SjqhwS9P3qXCd23l/sfBIwGLoaI
MyJzwNwzRbCrQaPi1lH1j5jZhFCU0HGYvmty4C3a7YZ6dATK9MH27zQMKDQWMCSUt4LCk0xudpwJ
esLsRebmKEN+jptlfnY/W+/0mZmwd3ylqI+e1dRNvFg/MXiZrSTMvqTXVzkfLE5CLNa3duSUPY/Y
hahr1p2iZpRvfD5WE1FLUJqUgHfNsMp9hy5IsDKrjD85h1UltC3oyu/fEkdClgemL1IbYsd3WB1o
QOlpO+OpylY+GgGh70q97EQV0+7lTXLKi8aExHfP6c7yG+F+DqW2deJU2ULa/NS7cmgFSOixV5PU
NKmfrjb1PaHv3ZKkus9amKvRPCi1mAZEBcQQJlErUZBvIky7OTbi9+SdOEeJZ/ndMkgLq8aCYDvL
5lg1+1ZaxrLw5TdAvDW2BLeqNR/KRNOSBkC/JrfCV5VWGvaeNBXKAH4Wp2i4mdwJlWeawRw0J9pj
hZeG8lGZbovwfp19JGZDHrSMqMQ1gdKyNGd9LbCYFIWCWNIQ6rBO6LAbh2fdD576dthG5DcAbDSJ
Gf8Q1o1UvC+9w7L1vmklpNE6BBks6KOr7ktn2KE4Z4OyvwBLzTuvdBfr6rMlW3tiAD1kmJOqqXOx
R2ojZlMXF12GT7DtM21VZ0EuRlgCr9zqpNnbN4cTh2yBnmRtt5n1kioOlMh9Myd62i2XB1B1feu1
rcF989htGzMEdh4ca/qsm//JZxCMLn9qpGM9dM1SH6hswEI9NS2mlmpwwIHFZ6mclndy9xfBK3/i
BxooMLuTnrxmM8VJiglRbqBUI3Z7H2rBykvh/+02gVigch015yEeOFTykNpb1ZdQM1vTm6l3gPIs
kA2yTRslaxHX6OywX0ad25sie6pBu2oN6DnJ//PaiM6xRvALkywzxFgnUAdif4LTRzZ6ppmsmHGe
cEQVK4Yuozwqcqqzg2NhkMtKwnJeEDq8uoS+Dsb5WEhLOCIdkYVh2axz6KGklQl+/N0crxMTNE7V
mk/6KLTvr8T2VxmkyghbKkbXmjUDGXElnB8Da6CgNv5FrezLtQB/ouNG77vURFxz8PWMU3xWpGXK
K5V1pGEk50Tzym8NW8pJ4N7vuDihW5IYatjC3o8+zJY3ib28g3kxxv/DN1V0oDVqkJe7cMg2i8LX
W2CHwuFFCPBysLf5f74/q4p2i0QJjGmwXNFzFPXvSnyLQoCZeV0PQosL8l20fpYMDRgyVwy8BYqW
TtTcZKQnSXyQf59XQ6on6ct24HOHiqbsJcaFZGuTD5uvOFkNTcGdGKVzY8i6gXis4I8FUZ1mKP3v
WhrdL8aBIhRcs7PJlWvwIx1KNGlZPpc6ugY2PrWivu76lNcec66/fUFU0a75WjTvdmb5d2Mh6k3p
1RvqJDRqAWqKJlZ8KOlYBClqBjRkUocqdbrwG2G7op/jDRKk/pwQJ5tFjzG1WFnHH+kQijIfKfCx
6eRF+nQKJeDTv7DQpliF+48trwegk7X9ZyWnJ214QPPphsRKovDiwBridC/QIEk2ioq8Oj9kJFT4
63xRxaKKDnFmgQx+/I8xcKh4TsxX1DbsN0S+XVXJObn6qgpsXp2DyUVyZterRvzwj4fnjXtPqzfL
M94aFt+r2162Ro3WRsFTSTPYlw4rQb/8pVsDwK7VIQj9/pH3VH+6g1O3PgEJjZfPO52a85k2/rS+
NO7PQT8/pF0IZ78U7X3qACRlnLNMvH+10tk6hfwMcEng+W/k2XJGXbtTnAKvQBEC79W3TAqhNyLz
3SM47IRjRcerV0e22F9PTsA3eNGC173rDw4flMnV50Ir8A/AlU9spJYz/qhuB5hEmbktcgM+T7mX
kW0k9kHjcxGHlhjkP7FgOUa5MGvTWMBRYfLEnLYCdyTOfmtVg4yg7CFwHhJTWzbH5NZQUueW33FO
h1CIzqfudi0Bnfsz/gRSD1oe8sgDFX7Ff6cJO18P9x2tXKtu7MJjwtO133rsBNS7uAud9BTR8m7t
FaDUkDA/mTrgCpa+id/EZmrrzbWADLO7zuRD6C4sblSu0omrrVBqhLjMQesMwd4Rwf4LP96fAazt
PZoFyC3cQhgaUeUQtIRBp5phYXTSv2KYTShB2JWeJCb8pw3n8QgNjPO7fedEIALyHZ7zJqqIHhhI
cjoGcBHjnm5cMoBoZiFUep+muV+BoT5BWhCIqw6nIoZE6F3XWrS3iS2NOdGu9Jy6jdTHhZCIJehH
bCF0aw+QxSswbeaNqT4CPhxy6MqBX68lWPSStP+xjhSIo/8eJ0Ue1t7SncjLxfTD1vah7Q0yzsuO
fkSriLouLGQ8/4XHccPt9ZOIy+p80sV2fN4lH4gV7jjGwQr/w/j7R/BIaBF4osbc0llm5Rv5ghP3
MAzHt+i4I0els6y9hbizIZh7L51hG/q1vvhes2JSgS8MKRCAKMWHq+QVi8ZY1LsfsnqyAYR+YE2s
1aEF6goZF4Ui2d5+eJip5Zs8YPBbT93BlkNcyKOFU7NUv/mfVCtdZ3Qs7n5mPs93VWxCz1x+g6r4
c7lZOOA2IpGODWM419wVx+bTdXwOkS4W/gNDmQcIfRE19kSVRxabUC8hTqbBp4LR3c35/Smyvfmc
oNQVyrIohvyOR67extAzNphrF6kBPEdyu5JhKOzFzpKnfGrc4zjQC9hQR8kFJ2XzXQCFCUALw480
x9I/DtCZEXwPGO4Z8ibqYlSSHIJJ1a0SAyKdjgiIz4JUiesdDLK+WQrb2UbkfA1j82kPKBKP3WC/
M2D0mbJHVoOJcJ3QD5+YbWgOS+nxzjKqBhdBG878yMGezl2A8VxXhsOGeJIwc37OH5rsJOyKV31R
A6NkxApRZH8L3q8xZlwCOYoOImptTlVWYUjgbg5QsuSP7GDf/fNeODhlamzrVXQhn+2t4LdVTI/3
565LzryGKEwGZYrHGsz39BKRhdhNZSa712tEEKxpuatZn1VXSQ85IsvlLeeS+6u3lzk1Nh1ljzDc
Rq+D40eEoO7+M6zX3ZIIGFJOqwApUjA5JanIQiECsvdtWk2TvGD4qo4cwMWI7lnqctMLSgVosIq4
I3qi3IxaZbOWj3avO58ArSVg5Kiw70mbKE/SFdwFAercqXJFeGXYbF3/UcjGDhTMx6qDiQAOGGkh
aCSTZCME9no+Ewf5TNOawKClQvUqxaovAtDzyDX4pQ5jzjrcpDJjDYUPMn+jsthWYQ8QaSKb6ksJ
2vF1ZalyMGg5oLYNIh/4QROgTBx1JTGAWTtTUW4IQSmM3JUJA1KStcUo1jeXDOH9rVvmPo4OjyxA
wh5Q0eBV8KZG+ndP9mHyfYtOyiHIsyz8bqQr6CliszyyJpMDnmBNOLQoM76CXOClHUc1ao0FfqHq
pfwHfBdhjvYGpcszAPHHOHUTS/8HQvZWGYjXL4nM1pyJIuRkAR2F/QNJQG57mZrjDEqepV1jMnII
snZLEP6o9kFHesL/fDxD0hlVeeydE7gx6wHm89+jaeBxOYgRoEkkbnGkfNALVRCM25Hb0lAx/WUG
SsErQ0wXat5NvUPTJBdK1W8nH6+3QuylsTxz3gDOqSvTn9WF9XsbXCEMvebejXgVTw81+gAFMd4t
M+Js1e1eBoE7U3u+j2ioAbOEvYyDtk40+ET5tRvbSgQMRr5F/Aq/sBGWZMcDa9qPdM3mEXM18v/P
X30XzwNlzarybius7nD9x9cJLTd501l3v+hbqNofeqb8oHqHKxBBhsbUOUieC0b2B7fqD6CgyRVu
Wb6UE/n3AnZxm0h/N81ho1WuIfTHm66qU7TT8QhO1bwDDRoe7gn0tBdpyWVsSbc3P+RrLMXy2PAn
SWK8Hz38/o6XK4rG7otg+AE0t1KgaPRVExqr0DxJbRqak/Zttx7Mkgl8pD10lcVRbA8S15vcJ6AB
G8HcA2+Noc8f7InaSwSbhELpM4C52KUBav2hEB2fFGvkAt2EZ1vv+0tXk0UZrCXCTOY6hRHQMrIM
5ApbskcvIsggpVYmZAsn11bqUhURE1hg3UAFklq48sKGDXNjyvHma2mJ2LPbeM34wv3Iqec0kgYB
9TunZXsGmDtATPU9yVcZIYDGKsVFnE5BqTFAKSvafAyWa7oCnPNjYZ67hUA/BPjMilkzz3H+dghn
RQcwNvN+Cwj2Bxi+3jkWJBxPbqbLuQ4hhA316znJLXR6IhXVJR9OsyAbWbJwivHaVEdu26ZhIN70
jLx8M4X54eMkv+KGfzYVhRCq2OQkB4HPpL34Vni80/JJJdSVCPVzmxPMBMDknCjGKjR7scZEz9/6
zeBS8gbp3ZuxHfHp1TFh4TQxBuxan+5g8RWpRkmdxBGpdybwbCchkTgKVEG5mRoXlTDjCjTwvaQk
kPzC/9dUTrozsCYaxjP9wka0Hf5Ybx1hBGrc0pWcQS0VgUixuwtaC3I8wDhmCQ2urmqXBqJhB6Bf
P7x2NH3ux6o4G0FRnltVocuke1sMnd2xNeg3L990sxWWGn66QbnkDraECanJXK0ECT6bkdxVXd+k
ER/KBkBKHz3o0/S+QENqyou4wtPhLx7OA+kU4ElxJHRqZZZS5RmO/gRxFZcg23MN+5AAZIigWkKo
mU8Vcl2x3RdxROJrq8Wuds2CDVJF2IehtiJc1HBB70pOEaybs65vjWPIMtb63KVYfj6CpfyDrjIR
hEpc3xhLryrq881FiaDXoJ1UFSuGvaNcDhtNyXqC4bzrAYmvjhJATbpYDUWTi9opRfcpC3LMGfnc
SZTLEWRmo54/bcnJ9kjSWI6GgWo5MG9sDyvvUjaYje0TKsVLscHwcx/iws9g2kG1Yjx079QY0uMV
APKsGSMEOWkZeY+8zMcbQBYuMalfu19BDh4979G5xD6lkbii9bQ5Ih8hpwHtg2i58J/1bPGcEuzh
sOIHKVSX2rlSZa3VpNS4gpYh7RJaUS2n6lu1wDdbjqE+rumPga8jAx0A3CtEjwi46j8lW349sPEa
oUjiSvKL5v8OokclYAAUuAicTd+MmpCWM12HtbOj5u6QZAzMyymbro+m43zQptADBhfyCTk3lQJe
i0KW7EiopVMl/OeLKH80l4U5EiZcCYUhc4kuRf+6mlBAPJhAoWfRTMSzw0Y+GLeOyja6W/zCZifQ
Jtr09ZcKEm9W/VG5UFAGTExKF6PC5l33PaFP4GpiMtRx9Qf5dlHN7hB462GfCw8plXRvI8NQPkn/
7MGdJAPBOgrSHyPW1eOfqYX8sxOTggkFUEUmU6MNfhkdDPwx9BipJqou0YD9rD0b+bZMbFeRneRV
L6NtCVnJf0/Bfn2Z6mBnpB86uT0fC7qCNdkwwHWSC0u3wnS1RxKmCHJrDBRyaahLrRjDEKHROxsu
mAre+GtR4U5bgKQzp4Yesc2JC4ZfHRKFU6UXPoLmgUm5CC5ICViIJkfld1IrgoytWk6CPcfsIYop
4fM15OLfz0+sNBT3NgchWl52xTmb0gGXMEvQkwBIKCnpGdxV6a6G92kxaeMxrQbqmApUI6j9pygQ
59Q8QuMGt0zOUjcjYWCOmyyrCfqCoiHYSxciPy6XzvNENkzRgEkwz/dueKFdB3In/XrFv0UAvVc4
YVk4gk4qYp5m8ozEx0FbAJZ2HLU1NL+kHAzGPkawFaVt8WoMRs/9JycBjqAJvBil9+JSzwJMY1U5
0hhnMgG+YFT1LtIit+lktikkWFgr/oj7cyiy/ohkKZKHm7k2lCgN+qvjeSZWsMBby8++E2qnvBVI
/Sz+t9Lhzh4IBRqA8y7osWOenkNjxE3a1bgGuUtEZ7BzfDzqrwfOECbAjFo/IETqLo26H+mDUMf0
6UzSV3L1Ut8V4SXyLYursietsAmdIJpwGHAj1AzrAAO1ojfVlyOUymTvLz10wnEGsckU8GQVkbdW
yYpOCC7nMrqSaUkwC4spp26iUiL+CUbDPVd8aX47+iWje7XxQ6lzU0XeCX34QK85FLKn3HSbQAfp
HtebFT9mUR0g3FmNNg3tnacG3T9faO+bNJxzZ009ZDOPTtzlK+cyD5Y6WGV6eVX/lfmBAoq448Rn
/+MbsGDx2S89IbCuUA6hGMN35GiQ/vPTE626+FT9SBvfuANLBNtEnBxU6klxpmR2Cv+zNsQuwhU+
P9pcxFc/EGIIdN/y3AfCuPAemx5CMUMFvg7/8Lfr2VgMjgoBrHlUT6I++PBi9c1ItXnddSA6wavo
IKOvrFpaEq2QtmTt7VfrGLY/ejOm6sKvLOZicfrD8EA2uFPMUeXTcboLAyxsf7pUVD6D0HmsHGGP
0d/nzQwu5AMUYpgNevAyZGFTzIo31j3Y+5UnwCgg0WHkegof/laFEW2D8GXyfkcNoTkTbI1cNSYP
2JmKsI4j1nNfmkTmEdv8aP41uIrVZmRdl8MuSOzif3kDqnt24R8BKKvn8UPaqDZ4Y4UX+UtaXJve
Yu2CG4KIPB26C8nwDlXNT8sSumAe0FgDck+wAmQaLycQGRQYEhHegOUMAhrLfORDMWb8H9HY1XXa
TUHULAxlqYZti1UsbD7AkhG8gBqdPMLsDllq3zcFVKm1xwD5FNHGjbsHfI+jTVcjxGisDkhENny8
5oTFNoobHpToaoHLFsKzBpUAEwkjxCO47UTkSMOg5AUI/skfUUjBfNwZqZcOPF1q4j0kT0NANITR
RMvCBJDlwQ1IRMHaDcOlC3LWWHXNIYFhUxoKsc9ZZE309FNlxiP9JUmh35ONneR1ZCF3RCU+fTLM
qJrhQFY06eZZ1zGDaTBfEdaGnQ7gRGTUUW39STaO9LLU1kGl4AsbaYjXVlIWR1J+xqB2StbpS8Hx
H6x1kdV7SILcVNaimQsPhe/ZtcQvAIkPp+z1HoNHIsBpvUmxEyz/2e2Da0/gKk6aOQoN+9JYwR0p
Ks02qk25i+Ri5ZaTT3qiFOhN+16NxfS2w/PZ2ct6zqtX0/efl8p4nvbjuMMNWRRDAOYjMssn8A6p
xHgNx1VUe3B+aOqjUT0DrK0EycktDxrrOPURm9lX+V3Yb/3gZyAWs9jbArzVOFJndo0XOd4NlExV
Fm4ulqphqpkyFfh+kbwOTrQ0vqmTsndL0b4frrWJzs2cPUzukprjorniskCILQOSC6om4RrZrwwS
OLypKDYeYOYOcuH6rGIjbPDjP+LeQGt4DlqLsyfWZgg3xOiDOxw57X0N00bvZovdheX8BIGSOaBU
9US2tVKP3jykF65Iq6w63/eSx1aeQSzgUa/l0z1Tq9niqaVbS/P/HIreda2Cnv1WvGHczcfVLgH7
imyJtXwR9Usp4rECcecrTVPoibmsQzOCCDzpZoUmVvSc7LZYnlNWOWXN4h92BOC68lzCN9XRuARl
3H75csiHsi/NWCQe+lde3f+oDcipBF8YKFSUyK2Yv8OLR0dzfBac5AqS8JWJPiij5jAGPraoNWeN
a0VrJn03gYIO/SdyKjMUufNNxPksYwFVoRpmUO58KztZAbbPXtxLrHxXiXfOJWEt8luUpWumHcnu
wTK/ytChGVZTtscsnQi7LIB02NHGLSbm/o72cMIPgAHhYnommc0emgj1sludtmOjNm1nPpEC0RrH
9V0Xs40SFqorDQHzlFO048CsZz793iRR9m/TuZ+GW0GckvEayEBtYzXi8z2Dd9SQfcHWVmvxi3R1
qgTHaOhlvnbeoC/pvDrBFnOBQt/aRTGDBGdvfaWxoNo7wB9mqh8W8pdK69chAwKJ/jy93F8GAEez
vY4H1J07K+mgDnOtl7/sFC4bT+PVkW481qGSXUwXlCoCJ/HWAKSuHZv51QfhE+ApwRMUGo4+LsxC
YpaP9YwpPDElIAFVudrt+/AZO89+uO0ZYL7JoyZIb5yf+T123kHoU3WOunwIrSy/FETwmn/zEKAI
oCRBOMBviSHDNSTULGUl7hmGVxEu0iCJRPfECN56JgKwOzLjMdggb9EoRWEheCoo832B9ktQCGri
aCnRiFZu23fK3Sq9Gc00Q1CTs1qHjKWhl4TKK4sBaoWGvM+WMSnJ5U1UjR8cMhWphPwyMvL3KtO8
LIxb+b9G5M2N+ANnt4pTJevCeqYUnRdB5t0FYOjr9inPbYX9c7TB9QtE6eH6Q3+6RuxdU3eBeRRf
oIyfpPKB96UPJdk7F856RbZP1ZaCkQYha/6cLzuRN4hWn4O0LdWXW85p9yezo8Eb7GE0mpNJKFj6
UBNJTL+pneqIOKCp5csDRxN7CmU6zEXIiUXdHmDIg0JMuoIDknxBn95LaAxsCAH+98AUUYz6Qbvm
L2DKupBVJVM2jnDJsedbDy8cj+G7jtQSrljxZi2TckJ2xwHTrFGQNlGO8lWkP9R9k4CM1fpIG3TA
FDKB7T8ShI4g33sUUSU7Hlz5Xu5b5cYdnXuWQ5qCxMQY6jffpdWpw04egiL+AK3blb1Pcsltz5fs
X61csQnHXWJrYbHAqJ/GjW5lI2CPyIr4YhnKblJX1z4+Qi+ZrE0lbr6x8tyxv8Wk716Tp09xhOVE
su30FqH9+p1IDTh48n3G5wz7cQMN16VVnm3G5PpHOgBJRZOhQmEbvaqi4cBQyITXWvejaBG6VIeJ
HJlOyVIYlRzaNHQa9vDnQfQ0hfvzY9xsatFQibTvleacYOeDd7bqNDvJF7qbBANMc24HqdR2DSzK
WKbsONKfVePMUsVJHfifTMIPPjY6V5L5JaGKyO8VTV7cnE1OnI4ZOrs7qBk9Xlnm6eOb7LZhOfrT
AcZ/hW86cZVL4PNJR/MGdMz2Qu4W2fQXGVJpbU9wxMA22RjeptSaoMy49qYRnpuCrO+VOe0dl1rN
cVlPPsm+ljOmZL8NwSjhRez+uTw51r3EAqgNyU+Bvrt+mkkW9IoVJXzAi1tHO3rDBBUEAStlvgIK
e7F27OnHhR/Eh5sOnOxDjrTXaroqxIU0jbLx03fVCjWNO0Idq8OJzRXosXUcnLv8auFmRvUE6P/R
WnG6AjHxV3OHGmMKv94cgXVUQ1ZkSEq9mujrn2sbxnVWLn/AJN4z+fpeimpexUUZ2mZMWw9jV5fL
M5qQRM6aiFqf2Mef/B9XKC6uwprnhpTKl8G3y5KuJNjNyr4bOskzu3ljj143PuJP17Uashj6jHPE
K5Y4e51IHHk9e1XUjONTpq2goS/Ye4Dtwrue1L9k+nAEkhQHbpXxjSQPQt4BhZsI2VhmNTDYQo1D
edYCYa8k7qsLaJbhqU8s47d9f4j7gazz+0+tmS4RHq4WuoD7JsKso2ye/BsojqUG3yVisgZKiyC7
ol8bVTUhWGzvDG/PGcfzModI+kV+4k6RksEZUcEnq4fx9KVRZNeJTzhD3chLwRjXnzCYWZDE07uA
Ae1AaKke+U4Cr3nou0EZpVslCMJqF9f15bk31OFTSZRY3S/EObCMck7aF9a8aBUBd3MfrJEGOBZA
Rf/Kqagc1wdebXLBDBNnqT5d3appV/KB5Fy40hLXKDtHSaxyNLYN9M6aRkW8A4kWhZyI9eI+Uitg
VnJW+BW+5KTLMnJJS3YBxpI+jGmtduF1D7N9gce/x2JWvGO2g0ndC1eu+3YjkPjMiCJ+F+PMlIxc
tulQ0HzFeUkYs+X//rG0sjeLEm6yqtyOmrJNSFToO3+ueQntgmdSMdzVdF8LM28Uf4Ed4pdmCDHe
gUfz6f87EsCa9VNHqH6OzP2yB2rb1r5ekASI1lhbtppKpv2SRXCtGX97KtxQs+XG6F9QkV8As3BB
SQFiLMIzPq8r5laV0gW7DYF9lfStk6DVH0O6F036X2VLJVtMy9uT6/i5TNv6r0mJoZga1LshW1gF
SJNNuPQyPoKcJfOByWK6/hque4oWrpAso/5t8tv1+EJEcL2vRs6kf+k5hnJikLvTKyF/iF7LNcNl
QiNk6aLr+BWT8tyGhvRvliMh4sM3N5eB0ZVPHWVpH+Vs/ZzVgESpIAfY0jj2+63/1a8u5mkS9nH8
naQZAhJblPsLRtGuVXj4FQifp6EwzuMHH/HyBdrfu0tqC4qko8i1RIH7tqOSSqWm0+4a04Zc74D6
3iLS7U2nO16W0gD5ujxzO10ERlMsdnTfx8nwoZ+vYMDnVPLaLIqXvluLN/CApRBl8jKykLa1lqNz
DZIxOcMmd49DB1u7Xw+NC98b2xWPJvuZKq7HD+37lyVeybjaGwmk2bLVLfnGrh/vNfqLLrQUnjYq
3PnAM4x6OKYTReqAvoH6Z8rQZyEBVbTuo3Fh+KEmrFh5NDgbK8Qbw8A9BfDpygom0+8LaEeq6cXf
S758mcOSxCQ9SLkZNZB/tHDVMjngMtaJpvMWeSe1FvFJJLTrqd632qPdZnV9FjX0CgxboCyfkYRe
+4upTBnlCgOcWri87NaZVPbVGy0OB28yKm6gE8V7G+8kGyonC8AeUMLn8FwC5r7lqtMay+ZRardG
WDYTEXtZtoH5kb90ewqWs+NFVNbaVlGJHeaNhtvBcgVXca4CvoWkjZ38LlCgd8U849oqA3B6Xdte
MfbRG+Sy3KHWgkzqQd28Ig4E4gKWxIEaek9tvIM2qYv7VaIZGTJjQZalU0GQILbqm1RfkNxb+5Wo
XCEIWtIYaKnMinpLwMUC5yYSxNeLaOWWOG/Q3xCqqnjBIZ9R+Xj2gi6Mar/R5savGJx/BHzm3oh1
Y2+0xHCkvX4f6zsVa69sQp52L24dujdx7Z0cspOysPsy9Twl2GdEmE8McR/7ITqTcns+dwf5p1Mu
HIutlb8Tb6GDyK37MlIN8IWBklExLZ/jloNByy8evnPkoi5w8jYi/U6znkIrS241B7G1gPOr/DlB
6qB8Rt241Tlmwz4dtwnE1AGL8xjBmlxto/Fn8GRPaGPBahc22ft8348UKADS8zdT1HMOadwcbrYx
MD0ibf9GvLq0HNFYZvWxjpIdQ+7YBwmy9hsSytcRJp+BUlxnHulEoGFLBYR9qXZskqkYriv8Adou
I6UXJlRbcRm6DXx+jI4YTCBsQ52cY3bdcRJ6rPTcMuIXJn35gHLcCN72cQa+RrEw/Z+oGxQMmkGv
Yzs9+k3hsCJuuk85XUH14KKe8UwzWRfDlzxa0eclBrXUTigeInEPDjYO3q/UnpJgmBJS9Y9fUv5p
kWcSKWqJTawMMcso++vP7017OkuHuGMcPKxYQ3mvg9eexeMBlE1MlksUvV+hNF+WGPwrE+Sq+H6f
BZAFbS7tLd1bK4smIdeQ9n/29Z93SmnYn19deXTBgqCJAxRUHVW5TizJuBR079F8OrjiqKXfIwzn
7Tnz4EG66TGuK84ddgAKIJ4H8aBl1IoDEiAffWoxWYhGs2TdWrdH4LwYn8jWWkgIJvaxafV4Ei13
NXrmjWWM0PXOmO/Q/idK+3W0+x/D5I077qohAtItFlUILMvGz8zOYOZX0WAgJ+JQeFZDtFeAjZJm
2FinCVOCmxQvsw1p5ktq3YMYlWGS8VfwUXq2e4Ax5cv1h+sKmdNRNVwh5rLsscE2QdLBex/wPUrT
TzWqYFR13ftHx4lvjzfDO+hkcPpjNTLFa46QcAXAzt5YX/JpZdqKFpm84SIJzZ06YuB5bozlEWp0
8/r81BqlRC70IdPgmMPSYNUUfzBNJa38hOdXGqfzZFisI/2KKpEUCKJwREeY4GrHguBIfzKWPAUj
mdgBse8HfuLXIPi1ts/SA8m6XYEHOWH319Qp7gAIJ2VWArvcrxdcEv1MtR/sck9aN+iQ8qN7VIpo
6M/xibYvV+rrKOqrWcI/6dNPzEYl9QmVf14kv3D4XL4AUVRiz27xiyg8C7Z678yJRsozWqzdqfdh
oiNDebipsuoCIf9mtUnmQz7FTrA//9unJKxDwq1kKDw6EKL8FnLNxl7a+KUdpECVd/hofzm3Bkrh
2TImMcjd+et8AojXRwXCYrEipwYW4sUk7/p1DOM8B5oGPWO/5Ex15TooirPxBYbfnN6FplJRuoHb
Sfmf01CV0c3i4h8Q04dFLRgBC/s0QKXwPVTSNc4SSsb0zfBHRUpiiscUrYPD6Itute1cnVUCyTFw
0Yag9F+2oFNp+voaCSBKppmhBwG26uhJ1BV+CzG1DwnDkQyr6RlcEM4dwyp08oCvqmkDK3eow/IN
eF2BMQc9iqlipETrk1y3ndRoE+QJOPTyp5EurPNO9T/mCJAi2Hjwbo03GPLjK3ZGwv+oDrSGQtge
iYfNVASptk77pYHrld7Er+lcoYwbXrIANcNkznuVs3YiQaR9YhUH1pWMEhUP451dGjszRX51g1+Z
mBhWfHgUgrX+syokKoduGlo1ZgTvhJVPL1hp7+PGeQfzQX0uz+VxmilzcCONzzsEzSFeRd1oI2QM
9LBQLd8aVk7rwLkoOtDS8Kv/7DxqzFIw7nWa5+QTcMJqZY3LLXNngpbw1uQ76BpHuvMgcvc5U/P4
JtNoUhAx3DhExtaAOUyTPR4ZrHjgulYdW8fEKp4Et54YbpqIJdt7xyyRIDUnUNtKKSo1QdJvLCC0
MYemyyO2KszrKq9lQJ9KImD15YNz7sn+iJKGTNkO6J7cGmEfwuUaUM4T3MfXV+Trqr7nfiaCkx4n
2vuFAeuqqRQVyj+mA3IFKJzc/EZf9vQW3fPHmFMT0Fzw/QtmAQFUYiuR+4HQQVOC4SaSeLXv/70f
b10g0hzTSPCUh8kItKu4qxkBRiQc8tilWyWUkqiBwyh/oI5z+ppbaWEMencrcTSULlSWTj4NS476
b2M0I6w5UK2kTRMedVt7gannesUfcT5HLv+945jDWl5lJ24pgHgouBD8vTwJ7X6KNBGxToeFKaE5
Ri+BGxigaPuRQpRKRlGT4DADwkLU9lCMsVUoIVOA8v1Zu3g+WOtTv90vCHnHG7qMG+HyX90Kdnmi
sXorL1ZKytycHTkPzd5OgdOPykqjcp+srsvEu+yShwb32iRLef0sz6L2npSihpi6gshxhke2aX6n
zoVpWT16JrVhBqs2iPllOT9/dOSoydQSm034SQiMPMO0+aCbmDr4st21yFw1wy4Lt1yfqUh3UhEZ
iCVdwcGIIk3bgR9UmemVvJ98YL+DGVvU6JZ9vQkNm3tgzfwOTV2ArOb0lrHJMzZ9ec8ejaLqvqpG
mMFGw7zhWTGp5IVj52nn0OOmBTcCEltw5jJsV/rRNqwdUOGsQl7St96eeARkTT8XMOkvIA97+13U
GYLoDoECT1zMQl/4LwMtZkWtW0ceLTASe8yG119n1t3nVl52iXnjz5mOPwaKWTbzaCweKJ8GMj62
tLusBbJop1KRt4M9SVds6o9Lc9iRlwnMoZT3B7VPkq/HKBobwek6lnUAM0wJploY0xWQal147PHE
+/EiS6tV7MEhutsc3r6FTqmaawhbL0jI0y6MnRWIBR/ps+l9DCZK7YkItBtWWcbxz0OOzkigw22R
fM1sNvlPJb7vHxwovNO3GSyNZUASJK67qKJk7pkJJsseRU3FpBtvvuTgZbCZwBrdYQeRf1yR1U8E
Yu3QSHD+LHXN3cW9o5DQ5QDngwVHNFdZKMbdWN38QdhldBiMoZstvh3687pQbwju9arlYO5h1TsM
XpME7D7LdOGcsu2SXP/+4ok5lD2NzEAYhQ6u0/VU9cqXGHUguxLy+/J/iFy+34lU5+o6qAjbdmo5
SQrafvlORlwDmq5aZk4tcYuwzheP650QGbUJZYsFHSxq+fY57uom8ChmUe+eIvrcKM6aP8soQcSQ
SThVR4A30Oa9bpz/uykFWKpXdl1ivwxZC77i5HrkfrRFDt3UzOjWd1JZEB7g07aeIHRfaMSSYjV8
97QsZOdEDpiNkCHYk91ho+Yiv2D36L0zAw+D/EZwl3M0ybTHwbl+hoJf7JNYMLOAytyXaqUE0for
GEISzNcH3BtQ3Ux9cUYuhN2aC/shktGfK70BMJdpqS7icplF/dM158nw+zZ2mxuOOqOOZ/u7Sred
DFq7QytvQy5N3hMKGWSyO4yJwyEfYZ6PfA4rdFupDYM/Ieti84B1+nEY7CIhn1XSmsA7SZ2KOpDB
+QxiP3vCqCDVWmAJ9zcVXXQnW7mXMdDRxDZEn9flj0/i68J5F0jRsnG9mJBiWVVZr7ZqdjrC8bMp
RosCusnfQDIPiA/Q6rqUIku+zNSP76Py2yQs6Uz3GPwXAjR6DFejmSR+mFy4/Ma8AVpB/EmYl1ki
6EK/RtDKBwAmMTygWBlHGJneS+wD5O1oU6eC9UzmmMkOHBR7vHqp/FusnPElhikCccbyf1X5GVNh
5/NPUOU7TZGjHTQDWDGzFIJDugFQNBHF8MOYq+l/skiVtGij/k/PAEirVCzYYCYSUYOowNxqTkpm
itArExrvjWaUbxKEihshFscT9vL8KUANUhwIZDBJDsIAo9yII/qcf7Giquaa51VZUp+Y13m+ztZT
r+bIRsXe8amq5XYF5HAZxP6AkPSFjRzYBegj+DBnQ3Xkx8nU8oN23EXWowLWGweRT4A52YUir1Vj
ZiP4DOlNNwFo6S31eflOw4iO7Ly882+NY0ks+2oSwmco7zmygdV219sTu18kN8gXbX9bFP2Wk0UN
TZjDoOPqAQnfE5QR0aEKHfAEoVSuZnvBNC50rFm3LaHxQFWD7A1KWm0VYSzdJlx2A1SyoDI5kR/G
rNytsxISQPeUb4iAlJPbKzjA4mifsgc6q44iXNTNeUviL4vgRvVsuL7b4TejVhA2w9rbHKaXimHt
IAUw/RKTHpRDHbT3XhtQcGpWfGJdl8ahYggM6+TGkpJTyzUQ7kguj3B+IkU8Ef3pULlEx3puKP5G
jcDGmtnJLqJneZY2vCRflYOaVO3YEm3dx0I/ks1kLhrGsmHvgEf5/ljEmNsELisrxjJGbu9ZbocJ
zHboZ9wpv3Y0O1xHJ6RDiI6mXZDX8N2OSXvGmxkyffy/uya6HlxnlW1ScWWuNLy7pGSNy+ThKcOa
VzJzzXPBloh12Pz6E1xU9rSZ5+UxhEXV8k90WzFFhDvxDuP3rXSQ6jO3BxNadjplJkxS8Nn8hKqK
+RUgMWY6AFUy+Uj+xCE/45uTFCVtdsSlr4MxJt3vTUTxd0C0n6LQrFpWNKH2RGVh19KU1Hx4fsjm
WkaTJxbBdt1wd57aaO6BnbXnbx7tOAr72Evn76BlicNpbO9wQFaR1gRI0BCKVVsR1XP8EjE75+MW
9wZwQzCHoV4wKhTZpbqtYrXub3taLc6bxWtSqxygzJAK3rXSq7vcnLIhMNDszM93nAlvaLZqF97U
ENRECBwQqGcKDuwSkT52YCuWTRtT0iHn4HcBDroKZn3sDeZb5D3QDuzyFNb0h08GnoQaumyYsVdd
s+7eUbYPY4MTUWaX80yuCC8JExWxkl9QHhim8MEnjZeo6BfUGme1tl+15UvZZrjk2n+BPEvVrUy+
njJkJ2BS7mUmLXGO3NJa5dboHDa5dO6Hv4tpf9446c1nHnd4yM/KG4Yueyp0ExQUtFbMuG+sJIRm
VOXqDuLH5flYtTHzcGtaKqXJk3fRMAcSofH2BPGeZY7ECN8Ap14U7JNRkXabWeRtSqcW8985zav2
qaM5JNBZCCuL5JUW4xlQmm5EkM0UNlxhOyyNR5i6epZghebIL2BtKSt5pRR2klAy19RVHbydbr4y
ArNYUYFjUyq6juwot75q79oPFYOg+uv3OqD0V2MhVh/YJTEt5elTuyDsA8hS0OevRXsQOItXlzz7
iKvSzhpKvdIykJLA1uvoE4H2dtulbMBCDYU8aViUX2fsHfAue5d6gSPpnx8KPShG7uXbgkx5RGHM
7HjoFQdp77TSYdrjvmY6U00rd/JhnvkryDpszZfPOAq67Lc1WlALejq7M7f13ecsNRmB2E+C2gn2
GWHQ4rLUCMHEw9X4OIK8vKNtY3V3EAMoFHwdbdhWZtwnV7RyBZD1xmV10rBi0NGvGy6nUqruSFJm
Wy7WovKLKB8Wnot56DCnCF13Q7WCDSFL6Sy2dBhltQCa17cMYB61x8B9RnxTJWQ6BkEPteVcGjWA
JZZxiNLtYyZMmJO4Fiz1EiIYvP9bgV5+eh1OJfbscG9veL2OMZQaNQ6rN/S2MUiLBLfMaH0lAYBn
PmUXrdmE90wi8/Xgo5VtOhlPTxtL9eEqc5ypCJNb279ar4aBSovUBGLjK7Z5sHuEn061lVohLeeV
Egmvc6kqDgFJrFxtToTgao+9/z0jpGeF+SmtlLW1KQxUUFQwdpWEJbeDlbhTSa0MspEgQ1w7Q2RA
dfE95OeNPWEz3d/tWbwuiEPnZKEzYhJQkZp+SAfaQ9gYoSsg/SpWEHOxyjdqSmVeycd2hcwRnKXH
O79xnfXG2SczmBJWrTGmMRrThVHW6/Xj0tr3IopZbpRVW+AIbkvnsQ4I9ds2bA0WOoWjSo6TJUT6
k8HimSwV7CArm47PVz/QQFoFwW6SaOCVJtYuQG+yV5weJFho+Nhc/Z83x5Sqs3yGkHQmrr9Nub/Z
fhU4Q0xy37se6K++NEfNYHf5jD0awEHLXOBWkTCe3jJERJQULHr3dnNzWazIF2EmBr58otFRbxDk
Kz8MZ1t48nFMf8JOYvXdMgNFy2G8WuWEpaa6JqRDxFdh5D+4sF9ZmTRZYk/XjR8IgDd2TbepfPeN
E971hPFiKa3twBN8TgyOhVScfIchdkGfamOSLShUynxRDsMtZyVpj7+7HuyMKGZJ2w8YQ3BZhpx1
3VeUScvecdAQmsNOW9KfyAZTaLvmYhwd0Ekrs6WoGAMTsyafkdQ0Y4xZRLDnHvP/ml6b/erBJto5
+i4UA40xP+d7B0tKL1gVcMe4rJGDwuuMrB0X1EYu2GXi9GUYm3e/rLGPPtEFWRcOzTGVxEbMiyVa
5LDMyookiVQ0CCu/u2g7X8vpyk0j2SLQUk9tT05pjiCnODjpPMbOpLuBqCcLHMcEFRndHUP9CBLg
HelOm0ajXSTct75epVpysiPLKoBEmJZ853H7YBQLF463bWomSzNl051PcUXWkIKLgT0S/Xrrpzks
5HBGKohk2c4KSoAHNRD7qVCOIS4SAjGDoe7sff3cEPD3mygPj1FWikQImvVsktURy/iF0W+AnTMJ
Cl9Ss5eFBfTX40dcXj8INu5VatcvlkLwtxajnaJEMsWSH1Xh6FkPdsd9qMDex3oHoVwwlBVJCcF2
gWJkv5tbt6qOa+pwxxN1eQiYH1PDJV5idwcOLDssV6BdNinUiWdlMwQhyrznUjpBb2JsVtVaqIP6
hgZmsnWf9wCkyM2WKU/8YoGlsSnvAt1Vxrf7VuyXtGZYHmOG6l7FXqcEBU84AvqM3H88AbLpl9+J
s1ZFDxbIaVDN6jWFVE1/LYb/MdyUKYCP0LzToY6b8U1aNEbKain0IWx2jVzJuTvIWG8LDGPODbA/
uWmeFeRIilpE6kx/HlrRB6UPVhbrK4Oxmf++EmggMkar5SLZoasUb0Su+seB9ifC/A6KNqKWF53D
l1AXbk1N1m3k6EwmL+FIxXiRjyfvhP+eg0ulq9EKDwEd3+qHHInL48E7eNeJNL5Q1nheQ4XZnBLh
4nF0IkNAsFL9xB9lJ0GvWou9EBFODhLqUib+7OYKhQJtSwMmmTNx5rsuQaZjL0WzlQwDSga4KYZz
pic3SuyUlhsgMAezSolVp3HVDoqqf3sSIzPiEGQ1g6aJiUJdUfaUiNEI4NIqLxSeimyW5yS7wq5s
zsINiN0DZpb0hDax0EvvRGAE8f6UMSk1c7EXfCJ1yIW6JUgekhKQ7AmNQ+XJVzjEJ8XVNnXQQiBB
Rb3NxdyOhIvdT/PS170GPC83hW8tpLvMcPXFBWdgwe0v4jEVezZVhJ6pRZDXLEetFIcjnWqSJswB
hkj1v5/hIcMwqx4kFttD/s7fsJf3ZnBswUW0s+4BjGHmFyfLe5yiKM7lK2axN1Eh0dPdCNtZpfrx
t8jC8ACd4awdfeFr3VNNfYRZdzLu9+ZOCnv4XsAFVpvYw7BIN38Dldoc0ym8NYu5YRwk4IuSjrpw
bDENSNT5t/Pq3m/Br6j0O3sgZDX3hzGHNNGCyILyT8BFgPoPMcO6qBw2RC1OQJ8OFUtQm7Vr47fm
FloJSWVfbtavfATcAlTFC1mzuCdYM87sdz8f+lZlws4qb4or8py0ZPLoP9aKO6eydZnkxjiEw+VV
IZSp58aLltzmrs8AHZLxnErkvc7tJS7XcEPXriehM+1jcSYusomOu0nKCrzilM83vCrp8CR9hH7x
aC7rBV/JqfHVsLOgWbGV6EFeGb5Kyn41eb+Zr25+WutgQ+AC3w3BB3+XzYivs0z/xGeLMkGuFiF1
FTE5CdhueA9kCwnEqAS9DuI1/HvRB9qzf2KPyf9R5kCi3J4+wBP3k3WnhRKiqM/yI3A3aFtbc9gd
o8nW2jkXQUj7zpsGviXmuAKeTF8z4J0FM8HqVu2+y6NBo4A0ry/dMVpNeO8DNsXOCN09fr7RSZwu
P681SQgsx/0p/RbiX2COuwTCgb6mBM/s/8Z5FqAY5m5NzuQq2GE0Vgk+30xuHzxtF7wDRiaBIFLt
/4d5weNKvWyaZuJLko2l7nXhbJRNv/nTN9gUQQQNaB6EzUne4T/F5NjqqN8bBwQ7Nn34C5k6MYcO
ruQN8FS5y047rPMo73Hrye6nOfX/BoWhWLbZMcSyxQOhUKzHlUIV1q1IIcCBg86vrR1yrXzUmNuF
PO5D1AXyJopfDwFm42YG0JTrmWX/PrMU9stgiyBOCJ5A6hhRxVUmcsX3gmM6KtMVYKrZ7xW7ZBHz
tikBPYFgCBkydCxDHz2b0B69Qiapw2pmNxYnTkhpEjCARDBSE4zC/1cG4ghmE2K3jbHGud8g4U3s
aW3gM0oMMmmwfcKnAhSVvkdNvdA+Zg1NrPt1WbeDp3rEObA/YsIsmEFQfc+NUPvEsohb8/4OXgBD
tOK8MKiqHu6a30JcYwP5NoOXjLj/l6eo7PMUSaJFaFeWKCzkWcNTGeCariOv877tidKxvOpduBAu
qwkgBUPlR/j/1gueZXldfJu8WPDYuhwraBWKKqr9iwnYIP/ZaMm3BmsrXDhM5u8rd6te+J3gfVww
LA99SDu2Gi8OqbnfdWrTpP5lGqjK3oIvC3ROVJ3AAzuXqbem+oJtl34Hg80NeHl4fATwzoW00g8g
/7YcG25rjOcM6oPlzqerRZNjMgTJN0zo2UAQKRAgDDLPpsy5KWAqyIIh536cT1JbOBiq+O4d+HuE
XiS2tKxqax8YiUKXDWm060qqcDjlhQkLuR6bl/4W8q/2Ew8kHLd77Zi29s7/KQLBt5YKsN1A5tQA
QrJ1OeajhYYAR2ihApNROQf/SfPvKKzRFScVS0WkXwKxcqdTIBHM1cJ91py4N2qsDeBD4EFnkvvj
I/Idp4yu7OqNu3+NbgZ8i93HuGX2xP9LPBHUd0Ul8e0wIVgqGJWXhrEDzRvaOUoWTQdvYqPYfmx3
6vuulJDLsx2lYM1XbwUnMmEWuXSPcG7b1nEhKf1OiIX9o3OzROBllh/CTIMNCJFpuR3ZDUFVTchb
QmBulxsx98H9RZJXtFS44kmSk1906riTRVfjm3+Ulp53WHTIjKAqvyaLtAwhxrHxsJAvwIkESDXX
rZYSxEvf68QGbmZ7Am1iKu3GsNZcf/GlQtvD8k3BhRfEefONlWIZ583Xnm9LpV+7MSYWjv2Qp/av
4gaowABMn8HYl1hLPayp3HipzUorLqRlnu9HvJZ06kkHX2wuo9ReUbqEBZZw+fdKrCk9A+N6GVj/
J4cKvPE7gD31enMoime5Zi2ydR+hOXXMeaSiATkrn1dTSI8rLminCIxkB+/OV6X4u9uZGdgnfU6E
ct1QiC3NAIWimgDmxIGO13gOn8L7Fh/3CK/hxOXbIv3v8jXRvBRd2a2g0GI8vgRNmn9FF/LJ1mJS
+zxgGh+MV/OkaJuY8bdd/3jdvh0latzF3fAIpykqerUuH/eRWK9Tyhvcdchv7nQZ5Ac1+htxXEBc
LPrxzUYfskkIZ05OWd9n1TPa3HCBT2zX3ipOcRX6d0Fw/qed6BcxiQnHg182rYs0/B9aB5OjPQDK
PCdMrFCiFtnbK88z7sQ50iuQgwFfxaLxr0UTAZRt8j3nZmticPc8iS0a9ujHcFj4IwUmHE+uybDA
Cn/VyWmkfugZI5NXD0d4GOeAG5fYi4WzTy1JzZS2hYRxOln/7TjC9KCojlh0E9g4hPs9S90x5S1K
c3O6AZSnr4HYkosDQCXBprROiOSPw7bDk69vKixI6agP/O/rnDG+pikxiixAnz3feUXce8sNiGJb
GR45e/Ka45CzloVuHom2OqYKpSXNRAXrGpyUHWHEp0/1XVHK2joKyI3BFVblbrlddBC63tMSY7fZ
zjxzBgBBqIGuSg+H85PoMwOusD6AKI15WNLdEq9lSSL0jcMQmJ4JsmqEgccjxumhXcg8YrIVfM4i
1XEdD6zc93u0SOsx1gMp0K9Wt5gGNBtj4dTFyji3/XYPjYQtJ6R/zXwHsNcqUv04tvMmcmTMhTDp
/q/I7gJU5mwwc2qxHVMzfMqC6zWvZpUcGrZ07cbB/KhcgPp+xa3mlQuqVuKFABnGJCsro9rnKBPt
o75eUWA4bF0W/HkJdMytBpGiCQHCucsBSbdw/zNn9wcVSituDS7HStsQSiT/MryrU6OOglanRTHC
5IkyY4PMWzpy79nv7wDmlmbUcSYNpRWusGXfCe1HgFLH8ZqnRf79lCC6oHRZ7bFpga16GT10XjCO
7Aarx5+vYU2mrwYHmqkeWmktSm2FnF9LIxwQYXJ1akiyYlTY2ds22bocdHUVKa94eyKSxh4eNoNJ
NqFsHdv4VjY7M8exZHrSF0SDR32bMqQGrLxjiSfed+FJVPmtp5UDEtTbr6hlnx+reNsPTnjcS3qd
CAXAeUbq/8xub6p5KJOPr0SH5fhzSX5N2jnErhBYfEmRnePEicyaZ8u0AGuXEHgM+0O79/K27WnJ
AgBsKgVzusNUrqkoPOqoRwTgK8JeTnqMIviWxyVGKEpPW5rhQdNBAOafkY5TswIjSq6SJ5IygK8l
0yoDb2CEFzbC+taoxD9gcb3FUsjc8NSr/E3r1L2L9/50JRBBBmXgV8uL25izrxNr86quAk6aO/57
/fJlfSn0J0WN9kCHyA7fzncDY98arlTQTEaL2vv9RktD0yGrahjg0id5/vnpX1kpYJmSQ7V9VEAO
8DQztU4vpKkhIIsvZPN4etI6UsbCCKpLha+zX6bfqUNXtXMiZRjppWGukfFy6E1/5bpLCceMKJLY
19XIyQuFZt6osafEzFa6gzJEAiqxD5TSEqah8GpdfD2chVXnpJsSlE8d0obuUvpHxUJAgQmEbze3
pypa8Q1rSGQ55oE8xEOo3qDWDGQ1u7CO7ZZ983TD88DS36vhIonx62ZSlW2b9l/j/wMdUyOdDDYM
Gao8BKCjc+dOZFaPS+pRADBAEqT3y/FuBZj4HCWRhlF8cOu0YcECMJ2gkC+jQ96HO/ixF56XmSzu
FO0oIdItpWe0HfsFH+BFhrZHR8hCG+UTyk43MJv/v1h4NOnO6YTb/0l3q0SgYJst6quLZoL26BPc
rIh/rw4vR/HKaq+NdBusEHdqO3Seq6sjO7moGdnoOasUIMR1uHxwMBrh6KIg4JIKTt4pIWBY70UR
2bSY+gufBwNk5uEa3A4jxYRLpKa13WHJ71+gFPojaJCaTF5gNgJ2gEsx3u0TcoGUKky46VUd6Qj/
WZb2OEheS4XSAWEgpnPobixbjYX/DgFxdlKcDUsMxa/N0hY13fU+R/9sGESgkVWsJgOVF050vMxL
A8jQN+xIvVJf2n2RNgesV5Op1hQu0PePEdwSCM8hIo2GR7UlTQwgOGHFcOuiCCHAA+FGVS5Xudvv
xumg0IfqANTkOJlUekrMT5y0IoQruYke+wsrv+10xndo58KLcMXMbuUh0gv6vyYnLeeHlwF9PYpE
9nUOkiDJQIQH3RGSx6GY32oPih/5wJdtg6hBYfkP6SmDAhY+pmxKNV8dnvVEdmI2f7TmwMToPzUL
vQGLjPimqb0fdvED2cU7ggTouMepTYedu+P+qmrh6C6MCHfRsZu8JkOmJtUbYx/675ouNJ05Ywz/
ERvOmMbK3atLcN6Mvl+S2sdPTg0bVxSbjuhpVeLXmrDzqXBpOXH/yre7EbHg7HR95mV0GUSapgxt
ccFQb0yqR8ehgzJcVdSIVs6+qV0+old23qy0hX0zh9laQGgj1noBKUG0TF5TlmDfPKP7ku1KG23N
M6dpbA5zWzkn4jZU4cTb4j3K++SZAj+qFON/Qejk05/ZCQ9SrMh3pC681HThSZ0oS+Deq5U3NLMX
jxbXamOw1H4dl5atkL5TArALdBQXM72s7sE9QfvoWRqRkq5+tCuW0pIXGiDBo0q8Ys6JHouQH9uh
CbYNhMI9CtZ7XJcMe/pBKcp5qo5oqrSGo9gGtANKAojLolxClHWfSMtzRsPXOe6ompqhDfub/huj
hfh1/5TpxBVh7l2w3+nkh/NlrLxVsdqlasGuwE1+Fsw7N37dIeTMn8gpEFe/3j50bqF6s4alxnUp
WcPrOtytm1ygGKeR4ELcqa6h9AGRtmRYvQw0aEL8YxYMU3FaS1n8VIYQe5lntP3TmLZZgKHQsF1B
BuUaNuLX4St8XjBtT3sP8yCZ6sw6KTMMAEXboA73qIS3U/4z1vDrOvlSJHxwkAGfZxLz3dmY/hOb
duKGX4+oXdbNNhbVQGrEfqTucZIrV5vvOjsbMo1eRARFTA2Xru1IzcXjGU0HexBcMsYKnGWeKm5y
xej7mCNQa9YPZgfxG3AtddHJHhuDMLrLVO0chEG6L7qqmS3UMac9Hb6E2PVzMZGOFFdOxo5TfqqB
mV5xSe/wZaz4+6wzLngvt2k/E6oUXxWMvbmSveDHGU/Gj1L5/quImF/eq4shMwF9mDOAFLbS6fMv
zJGsU0LTKVMD7NCXGUndisizyQiE7kzTqHTtms76GaTDQqX/7KL4ieL0Mri/KHjphZvOo7YhP5hu
hKtWksw7TmK/c/3eOMYDApU2i0nj3qDC4N6yHVpt3WoD2yu0VTTWxzlIPviFG2Szw+wRUXt/eJZ4
fYXYytxE3/sAQ7JjB8vPHbpj0d+PPDFdXTJ56wIl+gC4MHL54xpAPDCjf4nedsM+5hnDB9UJHhAB
i1TrLI87sxKSCQ7zrjU5B7ZWctVBUtuqcjWRVBqqX9PM0SJox9KTztbqdMWchV+p5scFEuHkntKD
MQhSUQYUAtaXbx0J49e1FTgpR/U2CNgap5MzvycbMdRo67kPN5zwuYWqy7u3bNjxjCt8xSfuRCb6
U6YU1AB7XUw/L/Dl5aUfLd2pxbgZ7wWrZcRr686VCGR0D9KAd225uvRg5oDO+gj9fGlmK7V1/vSD
cb7jeI9C6hetLovy13zeIlIuh8zUbTX03BslzCSrYBu4LSAcCmhjUEwClNwL8n3uA6Nd5LeXGiDu
h0yxkGC84sA7qmYbKyPhFdpqUw2wGKDaCY/DJOjQPP8UMK3LF1rnI2i8DqVsb0UUBl+rIlBYs7VX
QGTKj9BzwOD/vyY3Yznpin53uaw9M0MVNNJGRy0ViAO3uyCv8b+newui42QjRPJQT7X6Vg5AqGIR
as9n+/feV7P0je7T0AaFkvb0azqBclukzsDoVOZbljactObvpKPUtNmkuUtWFkkfisc3xeUEmXXP
DtWW7FRdeN2WC2xCDnRqMk9MO7DNjEMn6x7mcFJGZXDeHwCQ58EtKMaMPkA63JSnwKOeQgLOuRgm
Hl0bq827adezi3pHEIFla3WmSTrprZjT453aQxjkYn9XuIp8QAnLRR9ZEcg9jzRUtwvWQ9lqjPvd
FoLVfmjGtE9M9qM94sklBc8aGCXmL22ecSIqtrnX+9gAwFC/LwDv+vEp8wl4WOaiVtln+KLaf79a
QmDRNbXW57sVApiWVyLF249rJRwNzWXvqoPofyA0ZOEYUJxWvMVjqhwNj3a9Npy6K0P7xgMP0bKz
OvNzcdwJWu3JWNtb2q1EBjDP0mfyXA7uMx8sxVVH1qxrfNKu9eRDvtamBtdZKxGr4Gzr9Kp+pIQi
KpZwmzj12SP0e7lzQw3Q4AX0evFx9V08J9LvlvihKqM9nxWiQxuNRKjvfKiH0KE2oQuIzogExYLI
50X/dsEDlruYJ15+E07/exncXynt2IpuT8RlK40Mr7Z/VZDhMOKGotcB9uKc/Sdhu+pyAtpGE2v7
ipWkdMF2YyuAf+pFs96uFvad1jNuk0c7jRUVujKkC30Gz+tHkygZUTvYn6BdcJkzGTQ9uRmo3pzY
YsT46DppolhCcu0ZN0M4wX89U0gkBfr8iOQiKqpARE4XOWFXmT0S+qjvpazrohCGHQqNFgfo0GRg
DvMPCkooxNabNx/t4D4wnl9DclRYTls+hIaFEYFjYa2NhnCr4RXWye7lXoOOvSrSLzuNQa9mwMsf
ZsKp7a41H5QJ09I46ifW7taPfzKedjkdKawgGIZdfQuIkp5b7i4b6BMPYl70dgxK9zmop2Bw6SYh
2qF2iaypHwj+gCRJ4J/zNUbm+1ZK8tOrlN12mAgr7aEQedn+Vaz8Z5Odqcjpy1VZKbYtsaEO4NkE
j4MpctzsAQFxbZ6Y/2+Qr3p3wZmYG027RCQABichKX4kmNWcrg6GUtWyo+L0UOmnsis1h87Mi5Hh
EZugJT5HOQb1QAXixCHf1NIxpEM+/EOmW/SJDzn0YBe7i4S8RPw+0tQiCoYKLPI3vK9/59lEZ9U+
aBmVhdmzqsGN/INsmWg8x3YUeXua2rgAo+BbYufurRJn+TBdptOmWtMYRst3t5BoKbTSGiovDySn
C7YMLlg2K1kubJ7sykCS2F/lJvc4CTsPE4JJa0W/DxxsAhWEMwWvr3AErRQ8ds61kOqf4iqD9/pH
g9duCl3y/8/Ko/2wE1dDZVzX5ihV/ccN0h+QdlasdVdMuVFo9hdL14MAk9MqinkRxaPzBJ8XeqRS
8suImXED6jg5XDKdGGWkMINtwGNwGu4+7RENCHiKDTttgRszcgtoRWVV5nOQ9eGuDlb8ZD3P+c/z
V2Zv40piLfN4P+SKZR1r9+DFAeuuwSdcUrkWgbxpBHPopXZ7yry40/kHOrpiVw6z//VrL/bl08Wv
GautoKs6Vnm4zjGfp1SEvwEpaM9FWCv2f68/7lnC9ejS2QAfcxHVQjanjgWPFIwpkdYv1Fr1DVf3
qk6VNyZx6cLr8oJDwhFWZI+9dAuASU9Zg/lYMPGeM2u/t1+ZBRplMDUD5rCgchzHHQXctzBSYGZC
8Nc7EYUwEEQbptX4AdqxDfdVJhseR3L9TDlr53KX627wAkhwMtzVf+E2XG4BsZN1ATvEzNXu3iEh
GhruU1eVJyi/z3UIxA0lYLRtrGnYse+zwSXhRgxzhKCrA5gMTOdqxDzAcJqIehgek2NJydhhJCPJ
S5WnwBV8RyQXjhlyXNYYndNWF2abDBfuAHQlckEETYt+piDvJgkhfC8pwwDEDwAmq2HkNcZ7pcM/
EdVRl4HYVMraKt6tt8WwwyBp8hbcrk24DF1Cn22yoGKiTwFajn7z6YkR3qOe8a70rD1sZzh0gedu
DRFRFxJC5loOCF2X0i37AYfHOcPsP7pesicW8T2y16L4I6K08d5fnNJBfHCbK0Ux1F9FDRPsTd/L
D6CleIff1ZxhkHnuBtI1usPlwmi90mhFN0SJljtPb/4dFXzY0hkk2Z8pZUlsK6hwUlV4r7C8L5Ex
nGDDgFHFusceaE/sqHWRlbkH/y3jpFsEzpwteyZ+EDs+X4/HIE4aiU5QLZtjdfpOplCWatUr4jKC
JOP+PvK/OrBGsfcTreok0W/GCfoglWh518LRFieq1h/J66/Pt9oZJ4q97KrH6J7qyLxXMljaOC1M
UtrCk12y3m1SC5S8/vG0cbq4JJPBbYxqEa41Wd+1IbA3joinvnd2cu8j5kWs1rMAdX/UnRU53oJC
r+h+KRAHJo+AAotAhpjjh1jNZKL+31iTPQRYJsHke4DKgLqUh5mjLt9CvqnO+pHUnUFEwwV8d6Qi
GCjP2Yrc2lV/NUk/SvvhFM1uBDVGtZvNZuU8td5XyChXMxruaVFAW0Uglbd1dTGccspbo2Fm0jD1
4RNwxbf/jR15+Q3EObd0dLxq62b+S/khehmipoSI/NXogDKmKQ1VgcAWDSw7UKp76S9fq2mEQdxZ
nrmsdiPU2RMBt9gkhIJqdFD1c5lvzM9P7oOzLwDsOU7RrdaIDtRy97aHb7jL4K6QcxMjrpPkmr7F
l/roHTOWGvTVh10z4r2zXsax+dwoPTujAI0YNfvD0G5E+g+crEnIm4dmGvn4ozpssF4Zqf6I1apl
VWnfLDELvid6eX13ZRfr4eaiVU0e1vXehfaRM6xGJsYkCVtC5YG6Q2q+DBQ9WNqatFSsTnaf2PpZ
1a5QKqhmSoQtaWmRmZurbwg61NJC0DhT/Y5udMB5+8Vz5AyDclRCsUBQ51Drn+0U7PccYvC7wr08
tQhSiRT0S4Jsc84csoi6e4wi/UjcUIFTGje41sIBqsIepUC8HZoQfZ/6q8TY+Aza9LZvTcI/7ee7
MPtMTvudalCIkuCkd+TNuBB97N59xMPBRKk0QmfiFlBwWF8/7D+38vCldDOpt61KAcZXGgQKBSkh
6Ff6G4RfuGvaJaGJf2S3CnQNFIzlAYXm2qG1x5qdBm0l+XPHQVxrRqjAD17Ar1TS3uTJmgLMGgqJ
eFbMJC4jJEt6I+mOvySWM1HYmFx7xALUiBbP13PnAGyiAdjpyARRY6rrRsPRUxu1knxNn24u4UZD
mWHXMg6Ikl51tHaZcZ+kbDpd3o/fM04rntCnZGoMbMAWdWvRMJgPKFsqhjwCuj0ExIpERGamuNta
xFe2ow/XGnMdknbxDfeArc46Tn16RLf5fVebBCNsE7oAC4eN3OgGXrdhfHUer4+uzYYwZv1IJM13
XyaVGfPFk9a/BvriGnhfNu3c5PtLmUI95JW0H0s9Wcg04QHwFvOaZ4XFvjL8ACH23gYI4Nh2/yq8
3z8KLnFJSK6fPSgiTU6XgkEFIc7W2345RzxtqyY6PseYf0EvvpBElhOwEsCuSBPdL8UA58SPqcRN
m/seJKngvWwqVFnH6stAyefgKi6iQB+ynoTnx0aaxC6SvNybrrBLgZpmkpB2P7TlqMpETOr3eU40
af+HM9IOwASUqXA524bqT62BdmE0FXqanSD2vKxeKr0kTDaK3YmMJXzUJmi9qi+PgjQVgDf6o9Qg
Qin0C7JvLS607yygH53jWzy63bmI4rWIArN4m8BGIE/vHrK93G6vVCy06kYGIqH0JoIWOodXM/9w
YKTeljTDgQOu0Ip7oPVO7tw2NCxEBphVVqqji50bCzgcjNN5cAPxd64uYgGfb6UUioOSfz4E+eiE
r3a0lnWCDl39Ei5l7pRQbhtiJ/14TaDn0i8vkxqAVucOGHaKftGvbSg+LnthK2rS9Lo1Mfeg/Zp/
jP7BJvkfVSbbSgbkmvHspIbWOS0DeF4OCcgWxuDFqQcnr35iSxG1ki/tkFAA0R9xc4+5nXQvylu/
MfMJKcINgIbjBd+UiFj5kyretYQg8jb0i38OPs2U4C9SjKgM+psV64kEu/M3OkBUIXctVHcXuNER
UBvmFcqQIePKFULsyeTIhn4uCN1VYKbEJVyGb05IUmFHuBRQbdBsLcgZy+10NsCxRL8tWGuzYG83
7SCNqtW/2rKjBKHgTh1MSEwPTD+iXHd1AqIC1A0x1HAuCGowWnxRjZueBfexteCkfRbSdNvJVC/7
r1oO27YhOJ1ECVhH4NpcLdWbvcBF4xpqVlDrrRhoFA5Ilby1Kj5W8/ip+nQYimuY1JEwpxOlpxs/
Bm2dob6oCLOcW88pSC/lS6vea2wpnYmneM+sc25XtxjBWXhwCIO5rzvD2lMXTEAoKPQep2aIRm2H
UWTkFixj9O+KJserExw2o/mMcp7Wn4O1W0bpmV6Zkd+J8PIK0gGlPtn0ers5h8eetM1XNYUZpUnB
YPKNmnh7WOyeUwDXQd9s9XcmDvQlIgHKCmNAdjRxJjtuLaNNAjNeiOzmnbVC6qA0hJCMO7ht/fz1
ag20aeh0oZCB2MgxoEJi+DV6QHOstTFvPIWedTAqk52/WUs9ACjLuiwEvDUL2S2QfYU4j+blUv0i
ZtPuRpr1Sy7X6oW5nozcgorTtmAAX1D65ENHOCOAK2NKFCAiPRJBRY6pIS/shSjYUEKGTGixym3L
EkSkarUwYsKw/uYVNbvURW+wq9bzh66nm07EcXRcyrBmk9GsgBXAt05i2CO5KmLVokx3GN9oJ/36
xZsybuI6J+ceumXyX0YeB37ildJN0nmkDCMbEHSp3QlR2E+P4bGHTEgm1fosgdwiF7T4HhUh28e/
8sO+ofp6QpLYs7TSdG2OZjEFhrvBaUbyPHj4CV3t8dOQO13cSnt9lcK9OK9nrAqpg668PhZ+WtTC
WwBOoYci1zNF+bPdw+kGvxJbTl6wJWKJi+Ou05lox5TS0aGN/OAS8L9IBcfDYc6PI7czYtjB1EeA
ikuiRq6sNfMhprsnuRoJr4UhcQVmpkn8nnzn9ufp+/IWfnqLNXelarBc4yGBtw8/ky/2JZMvAd5G
mVXTQNd37QFppAowRH41nVtzZtKpyaqM5Ue492FfyWbGio6jrod9vRpJg3oCfytEFRyPJ5M4dAgh
3+G+8ShbcDD2dlvJ2N4ibVH6Ls34R/9LKV9A/raz64mZRc/MoOBOgtbhifAEF5sVXCqUXKUGWJVh
hNXW1Sz4q1kU6Gt2kEQjdWTCQkbw8b7YjJ4jeK/2zLNhTRTmlflKysamQaUgSs7mL+h2ZYyH6lFX
1WoJkdYtpW2pSbubh7iCwLZIv0/eFa9BokLp5VEe7Ebm4e1R1pjx7/OIXh4rsI69oQQuNbrsPasm
zNyFz1VdEw83KypO5xTjuPGs4Sb9vhqu/oYwRmPHqyMWWcBhJvDE3eM/oSQf91FA08LI5PZki7Ud
NDUFxjEXAL4jZlGvnj0vyGAxoeMXGTq6i2NPdDQoLe4442YS/wkpDiYatWEKKwWXslZZOOAlpPCr
F/AB0bx3QZ+YfpOYg/Cv+6caW3GOK0/xkhsEPxm+hxkkidpuGNJsESOBIhJ/Fggpt8u++f0T2Vjp
PDWVtMyBs//mNV5+s7nnN6oRXgizgSOjNmPHg5L3q7RQfe/UayPXGF/2f4Wv2h1BPnqVAqMg5X4M
mEU78aPLKY6V9zbXsdQPbTTYP6EPk0z3d6h8HezWM8ZmaJf+pYfSCwbkA/O0YGouHrvuL0Kd6bgs
Do8+kOYRNK24tgxYwLCMIO3rpLYmE0COE8HyDN5pTvuNbFWIVNkviHIhGGH6eBEK4VCRERF8ij35
ssFucItaO43bjSvnISWr7o6PTcwfcZRewOb7FaDzFnrOVFdwKDCXrKSkLMKYLZTFEunE1xCENvzk
PJgHKI5uv3l2eeZ267MgowNhmED/R2lBiAcQ1N/Xc7IV7R+jGofOUjNta5pH9R/ikAejSSiBMapo
x7f7fkj845/4J3XS3+KzCixfepCskrZHlleA2DmpDET3w37dTJ0Z837IlEGaBTfe5lTBwP9nDvbh
RKTlHu8IlbSnSpMlh0f9MqaV12c++wUgh4R6MliiWcdg4/J6YJtxuYEJ1uKHigzOJlaQ2X/TcvAx
zHCtGI2bpAmI5x19mzQyUcaz9ycVHkHzN80wItW84ypIWPyjCPwmeqSrAlzwLQp3gGQIfMH0HIjZ
d0Gq8CDu9Uk+UN288tcRmTp0dVkZWB+wZH5u3zPwpxwFBC1HtU2ArAPUNU4AOToHQpBn/+pEKusT
Jukvn7x9G2BFbceefM9iKv+5TWuPy3IueWaQOK7gK3sRKQ3jMHI3ZPCBy9chdU7hKlxpqK7o+rDR
epaRlOvdad4QKajI9y8mHsT20eGFnkaBhz+Sf0bAoXq/hMj00Obw9Tj1VzUobnUEv6GltZszrMBE
YecFjlngWXlIjL/uKLExp8ScCT6UAiiRVrt2TcA0tMXNoOP3lRuiogrXCWJ6s3Ope4lUnDTKqA4e
jJvFl7Ux1mGkeLD283uhCSFQtOhwWb+ggxNgpqpuknI+v68ishDiUwp0M94rhqHnntHeJUpbKox6
x3BQwZZxPlt/DfBOQtohisQzrcraQkIyvXbAif+5gBDgmYuClc8/bwQ3aWmCY/WGdZYFopEbTAEx
BfYDZg69E3CQ9xWBlfq+SYOSQXdHlooWVvu5Mey1BI/gYsuL4eH7+fMeYSwItjW4/nnfHw1yp+m9
Z0sTTQo+gJfJG3ijKepdIhfQJ6P2JC9WwmH/o0m6/T9D1I3NT8rz21P2zvXRPqMJ0Ul0hQ1AKLMf
7TbF0Rt5nH/ULySDzFQ2aWjxfa1tMO9ZZ/HAE37tlylF80Eunq2nYN/9URK9BngXQaYknm/yR9Et
Z+AC8qua4ixkiz7AC0FeRk9jPG/81viy11emfhMZHG5kQ4V96AemgsTvuwOEvN6+SJGpK4eXUyOT
nPOXFwV53Q6UrnO6G0XnFc4Q2cNrAOIGJnrDw8NwbG+xKpPKIZ/9MUOXUVGRrIVqdKcpYRWmIRtz
ssJ9YQPpwDJLDY2l9N8lD+SCijkEPvijBXqyKU9R1IK4FFdR+mU9us4+PChZWSdP1MedNOWE97/s
JxB5wP1oL8iVi1nyT6l8pCuHkBHhmjrR8s6W5BhTijv1j8gh7pvVHfRKoYEs/kYN27aesk81QVyE
XQmDYHieqwADmN1eeX0OOIH4B7tgXcXb+7/1rMJNso3r5d4gIrdq1FwvmqA2BO+sZhx9cF2HHOn0
sBJz0oQZCIt8GQJ9A4hHryEYYqjt7yQmJ3pqgE27X+JYioP7rWb3CHbsp7vtIus5KBqKCgbbl82F
kCtJOHszW0eHdljyRNtxqCRSjxXPC9bmtOeT2QQJ5fPg7HX3X2d9ynYNfnqjmjVmYLRQecbi/GS5
wfT07MpUezQvX2rnPk28KxWUFRx5FuVi9cNfCU7trD5oeBz79SjY4+bVQvivuOqJH46lcz9VWpb1
quBGi3M9d5MRGR9GQSP87oybUfFHh3FZyupZBlfrVF8ZjXxAWpvCi3z4IhLPFGM18KONcyNzIxH6
y7ZxIXBLyG3NKVJ4RbUtfMnM1rUf0LWOMNSqJANqwBWbZ4iWsroMsliwMTFr2tjXtoLo8nJpgi6r
53TKbbHAfLfh59aTW0uWi6JOwf1mGRAKAVQego26lTvA9GCWeo32nGE3oyb3/eTZcZLaIHsVGnCb
aa9bJNKyNfPdgvqpeD7eOEPKZOFa/QYt2ICgVRtAUVqB58jU+bW/RlWDUWz2pJb7tFdG4OHubyW4
faGKVFdO27poHklzvL6l1USefmI9d2zHCM8W5jJnqEXcucf6ZPZwXP2k2ee67solS365e0RhzYu+
ZmnNj5FyMGcHWx84vtb5DysFuSS9rBTxrCJJSeYgVd3Nm2W0ptNTn0NAwsFL9khBBVx4997xLz7M
jUXwXwghKsMm9ccw3uV9mXT8+xnJ4owu0VFvpR++ohLUhQq4Y8Z5bdDb8qoLD+DmqpddJX1LuZc5
TFAKN503tdI9nRz4VCUWpfERH+H2yN/ezrjh4GH7jRCrFflcr6AcsvHo3IxAKH2zVHB0YK2xWyKa
mGkWjIeOmGd9mvumYnEzBHLr/Zgmr4k7v6J9ZKGl2MY9Xr9B0tmiaI7jXUwSFlK22mQrHXBrC+bZ
Upm+OTcGwkV9uN1fvWEpKoE/MO7iVG8Q25XTujU75TsRLgNjo0TdYy4UGPMWWpm2w2KuLrqkBZYY
JOfvHuX1AEWDAFIaOMG0rXOJk1bdH4hiMkCZzB1tESb6PMaLJrvQbd04u+Z8ffh/ooMBfSE5iXhY
3OkjEcL5NveN1C0KTAsrfTB/pwOs7MMcwtWfeM4yza1J2EK/7E+Dl+io73zi/1N95bxdHq1RcJKg
i2Jrc5gM+jBqJH7+up3oOV8xfosYXp0xKu73buNMUO+XLj4SA/R5y6pbdHFJVRbRnSHrtrWpUZIU
V6xp1JXV2EbOr7QUGsgTb+gMqPA5ruJnfLTtpTLZe8r50Qumv57Z9oY06EtUGpD8ajbwwTNm0NIJ
dgTUKqCOsL2Ry239nqcFw7y4j3xvP1SnkpIiTmNYbqHalpOUxlfKfCV4xsfekQ3Wp9P6DW76V5DL
ojQnUcA36JNnwucbdC6ICpy+jyWH20doKsZbwQA6hsYahCpL3Z8l3VrNhRZuweJfS6rOqC6w6Nwe
pqHfnrNVGBPfOxq4s52UGL3yiiZhMiM6wkdb0LfB4Oa5pPzu8nIMh6GPlqU7z2BXmdndFd2d9VbU
g3hEtKBGiosjnHsPfqv4mdIlKmlnBbgGhh70YHYUmv+NTf6mFV5qv6D88qFUjYMfhgA3VXghRTiR
4jI3JECyvJEbNx/SjXSq10hOW5VHJOkpNpgodYl8dkdgZiZymbFOrE1Coi9XsnpMwZPY5Pp4dq3s
3lJSgfRWdRVAYyTB1wP5cDj7uwWIlaMkIzbGwZz9ImA9mO6zYzPw30m4Ll0eLV4LSnbOk1I9Kysf
Ycc1vvyYtU6uRAlScMEyJPR0I1jC2NoYhUR6KMLQu1wvG3QiH3/ZNrs1tCbOJx8fZFy3Hil/geGl
5dNEMSs9/iLnn9Je2ak83dQhbOFexHkwkuF5u0HIMDqu+dx0Pq6XIJ7LfEetAVIyCACx9MM9PWQW
CKEXmShrGRqPhO13i42DDF36qh0e8OyXH0YZTNfF9sLj8bmnsKLscP6YIppcpJRYxT00mpt9hBbP
f+hsiz/NqORKDt5d1W61dO18vTHfAF9pgffYxshRb0p63ft0eX4O0Rbv42cxoBLlI2UYv5XEsZNn
VxJ3jzmCVMZBxYYARUirpw5sXePl5M6nIvPVMSS8Qm4EFvdmZaC8AE5w98cDfdDCfdb7L57cMFQh
vNjz1V81dfMPDLFZf9ah9peN8klR56jGL95GNgKnJTMLUhOy78YwDpI/YQmi26VNyCffL8r91Du0
mfiygZJ1ej4ymdWYu+Z+rVmuW5kqI1PztTei+ryYRrxgg0u1nEXiySZXW31/daeSMeDvTum5ydNy
dZdZFPRZGvCjd/+q3tdjDntVrutyh+qxfy7Q/Z3OYJVBRZaYD8PKwJJURZM1VQOnklMh2DiqNDWE
fDc58F+0yR78G1hwubCkou9zTFlzKzGxw4n29y/iLkHTCb3ZRUf1apAUgdt59+qcWYo+8w1m60pl
lWiCjKv5TgQCN1GNh11uNApSgpZbkWQI+QEnMa26XnZ+1mc3gJzsndaRLjn0BfNjVD3WvNtlrkin
fSBxd13GtidxYA+lUxxZRxv7tHyUMl7YczZTMv+2CifA+wswnab8NPNhFsoULsdMfKmDM4dm2J9c
4z1699F9UrTYAMOtXmaZhtYo/UDsMNQTLWIJAn6RepAWYHOK8dArtlr0bgPRULqhl83iDuQJPOox
M3GCPCL2aGm1KalGecShLKVWQbZ4KChQQb/x5x1V1PKI0woyq3oyycwXh0DX6YoN4A3s4kj06wOS
+QsOXQrNWGWne4LbXDOE2LM775jn3XnkePY8kuYMNZM2qQW+la3eSDWoMcOELIYdijFNvMYyx7MJ
3uGPpAAaZ4l9xGcJRBy/VUt5+rEK7NedapNS70RFayU89HS8lT30zdhdSK7rQBsXrMXuC0gktMhJ
lvpClpNy1uCIApO7wLD+ZYm7+2qMVfI9AMdg5gaCZ/ZKH0cxo14+Jd+cxtDG+PjSf1ik4rFEQYbZ
CzBrcTdak2O32uurTMXuX45CXWJzUF7mLmqsd2N4moOTFJDpCOMMmXpwaF9Q3fTHJNtfIwn2ZKqM
h0ngHPRo7V9Jpz2SMTzyvASuv4T5kNsfguSeYNECDwLmS53INaDLimIxbva8GOL5tD7JPiZF8xGO
rGRuWOGNdd0oI0y4W2+VjFGImBpz/PWfQKC3RfLbf8MDk5aUv8YYLIJEODiAPPRpIdSXZbfpQi17
r4/Xcrpm7IX6R9pCxweIUhtt77Db/Nww5+vykO/svUgUwszWrHibeiulmjBlCbo8va3+RtaLi/cV
aMhiXhwocIMyXBQg64YVxMCyuNLVQoaE6eZN1pZagdxzQgf+YqVoraA+gbw+yd5m70eqhQXYA4uU
vij8lHw4XveiUsWGIYrnb8AIpiZTgVWVUQunvV+gONDjUOgTU0uWXvqhLPYtu7tuWVzLnXRTM56J
gDLgtFZNreglhlN0PaL0yiWd2vNuW93Kt0oVosbEv1B0WhsblhWM3TpNd0oWFjf8rJCE3WV+2ekr
SewzEibgBDhVm1UZkcSDpaC9XJSVHnoNAlEQwNTlysg79ESx3rerJCgLgKCzo+h5rwpnHzutuLy/
hXlar6W+0zOH7Tipc4OPxOG4/GXhhdXqJYqzWgkQ5OZvvlIIcyYX68RcuV7ZbKTgI3iLeH5jwZhm
xuRhuQG8jnO4fUSC6YBzp4zeg+w13TKEDlkD2T9Ov+mlt6/yzxkxehID1p7ZjICdmmKejTxxTtVp
Dtl8eT1jllbvfOCyAxDDb/Bbd3THTdiB6wqMk5fEWyeLSpo2yVSvpG8v2lKjGrMRn604xhXQA/Nw
zMDe8//vmIP47kg/IBjFGJ/nFTHQUATIv0yEHi93fuwzKI1BdfO853BYP5Gc33MPzRsONrBRy3zd
EZ42tdvaIMJGCBk9m0wO8RueT58jN0d3FbRSu+0PehFYhMkOvYdCBKDbZF3Y4+v+cxhslJID8fNe
KOISNzYoLWzzUJzyRzdlaFbdkeQkyhV6EonkpRI4yy/bZ0GwRgcl2ElRnx1FzvBazduyvSg6kLDh
enHvw0Hbjn8D/X32kBAe9W+BwwdmFKeooB1g2xU1gXf/trsJyvJTOnR11+y/2RVwY1nOD/Ttibay
qAjjTCHPal2iUk/Uumr27VQt1w9qJ92BHP2ceBlAEmV6Ml8/6DBXm/De0kPHiQhGiumLWNh8iJEA
bGgR+LSaAH4RZYP6SN7hG6B6bA6KYR8AgyFZ2+ZAxLG/3aXi8+euYfT3SNDrhL0fcZgA6tkgwmT3
eNas1HJZ6E+Gl806yQcADJ3BVAGq+Tfc8WRkcdhV2xHhjVVKFetzxM6oUOYQDA+DJXms/ONftTNN
h5Q/8pPcRaHJ+R0U/63WsHQ9j0AcHRgnaeNS7L+m4Oh/2eOViZLEslGJVcG+fbEcKqzG5lBFlU3f
fkhFf4yhhGqIfo+ZQhUWbde0jFKtJO7YRjMhihTsCZuP28xbsetCYTQv2qIuVVrvUEKlzuOvhow6
VdXEyaqRmX+8+7Tq+ej2hHcNIQlYsOeUmnNAL2HvNVPDbVRsSNIOLn4uRQppDftxm+PGtIxTwcN4
zqMkIUUTRzjQ3VJPzR76xR/4DqCHJmEfjTvNX6r8B1GohseVAD20JD3Cg7ouie9uB8v+WghzzIiC
KltjKBPS/7jqL711zA9G9/qPVvXy4jIGNCJrQg2keuu2ofSXLKXlbW+cz3LPWI3H9WBjQHDJxp+4
UOmJg240CVWXc/kZXx5iEhvBHjHbOlVAwRWbi4LH/NZwFtrt5NPZa2eaUrxbaLuiz8ebBBTezBEN
kADdp9WWru54QKog8xfuO/q6PpJM1UgSE4sC6rRS9BqOM0KPThBWjg5Qidshb6uXX9vEBeBt3tTb
ebMvUQVHuEdJKWz9epVwWiUfXhlMuP9T5gQyVeYrqrvuCn2tJL9W6reD6rJTajg/mD0TZTyUwMyt
SeZ5dIu3Skvt+KProICUU+WJeME4LW827Tuzd535HloHLL9LUgzCsrAL5zuXwZnSVulvud64NldA
TpW3SEuyMEdcLW4WvQdZ75acTjO/VqepoylSCHSPTsK1Sdjv1iHb3EfctvLJamwb5Rgmg4hp8gZv
ale+SCtEFFVibSdfyuQRu+jWoU1YtGWqiVnXBG51uUY+EbDJCDGB6H0HWNw7Pw/s7QqXX3zTPtUg
30wGqsVWoNvTF8R22zlaVWJuiid4lq3kp6Hc4RaM8jJlTk8bumfkIj2P1d0r+xkrtNjJ+zyqaykL
/r37DoHFwGkzs+oAb9hDmUEjzPPvFfH3fqhvx7HDJwBdWAFYsIFTwnVMQD+GioOkovzPE8kKWNn4
zU5DCIVcDXI5rVRgM1NGO/E/ZU1steG19wy44DHMZTCfMM498MmkO93DmLIj40e0ULVuemomWOtk
lL2faEqIvyF/RQW8FeXjiWncaEXCZgtIxKx95PFPTJqpZkf1auTMqS5up4l+bz/iS4G3xph5AI/1
WQJnvRoroduILQGsmQiQ1VV0s3NN/5gh45ywZDYMQtNwFF0mEu3oHs0frthcjeU48ep9rgBzs1Vm
zuwuklc0GWXA+17w082kV+o/MdDv1Z5eHSmQvvgvxodgRc5Jxua/jqs8g8YlEXlmX4QuIVaI71IR
0FjAvQVQzoPJasKkvsIZlFf1+K//dcHS4uwo6Z7QlLUa8o2+CCoCkfnIQc4aLZG+pNlk4JYCEpxr
A3wmdoUtDefeur51iHQ91zQT6VGtGsL2NTmSjOBaaSCXZNRsl/jN27RBwEBozIlzSuV0FluZ5mNj
XzXKndN9e4OmR0esfDKoNBqTZArX4HIMjU9RShGsckd9i6r3upooIcyBi/h71e1Se2o1kce/exw8
Uz6mbouB3z6BNU2dpGvGVNWg2aIVfraDgC4rwioOwAEV1FrKPqrAklxaUWlNv6keXqsV9N4OjIeI
UeqeQpz9YEnpYJTwd/Eqe9MwcTkcKsdxQywfjnM0EKg7BhHOP3Fkh3A3LC02ITkexX0gFPvSa0Ws
xzNjNKDngwf5lJdaq3NQPyuri0BxZG/3VPAQ3vco2KEj1TiC9NIE0RatcYycA3tU2aX9p0THlOHm
NLITAjCuhCiZXGiP8PmftealVNSen4e/860Lkn9LuTzm+Dz2w1wdg7jOwIgJrX3hGhiF44c7tN85
4mf0ycRVA9yZcQI9ggZmLjWOq4ULeE5+xKvP3TVtMwfz17xXUXHPmzlyYLPPXGGuL6QFF+PIHGUG
3Rzx9PAxOQtuMJhiBvYJdwOtvdF5IAYldkVUEjdjB887PnCUEHf4eZz5X/RI6sUjlIiYLT7iyBGa
tQovO4PTpZUS86S8yK8SV+ufoN9gakq+tVzUvrUrBdxtP3CU756r6SZmCkESOkFQ1TWCItkm27I6
0UVQOvkK5fis3wHj1rQYsjipVR4nPN5MfDQECK/EC0LLUbUpa263+/LDpGdpUp9T98snllwZTAKv
GeAwXFFwEHKC5yhrDbFITlt8h5/+lQwtHOzzBfFN8/ugb1xSKX5ANU7eIhkETzbml1DNz9VBov7V
1gxUTzK2CRluq6O9DILuxcBtAWJ+9rjOHG7+VgiDYt4BdGPIUPLB6/gUSLYVDZM6eQfjKfvx0R8w
3nRdij2Z73BveejBhytF2CgsnZ+zJNjs9d0obf9HGpFun5z0wkMrZhcR2l+LtYT43BE/zRmAbeFV
bcH+5b6eVBtW639SMa/WgM7R9lJ5z4v34DuerNcEdHhtkOn/IpzcC1sepqVGk1F9olEjLD7Rq6Hs
Lv9q4a6IVH6HGA2/qtauIV6rOaUuzteJsZFU4u2xucPh3wnpPVRIxXH+ZeX8CkIjzl7ZdlU0Ckfn
w5GiZSTgsq83mdjPeDVKOhnLbTp7l73yZ6VlNbnaR2/T9GGYETgJWLgAwlkGi5afZYDvdfN4Ggy5
yRUddZr4HspxyeMrxPxlZJgepn35JeYZxnHKJytoSriBe58TRo9nqRhEIGwMJO/3uf8mSPj3OBMH
qthe7TrUMfhcPoZK/fF8zsqekTtkQk8HCtWcF387hg6FvZHFBWP/zBEMbU9wmajJRcHjy93ryH4g
DqhzCfcsldxjQMldJ9Up4/dxoPCf/wff4S3XruoPN6+zHoCs/UfFwKEy8UGdZUx7T4zysIRLFc/L
zsldq9KGxvqRP6TiyEmjs9+2L5yU7A4hWqzNWO1RmXZK6ROPsONFgMXGUEIyP89DXJKEio1vjYs3
ps7uWL7YfDvfkzSIO/vLRmwC1BWvuJwfkiVaH6GZvLtcQVYVWCKrNHFXxThVki2u5SkhmqJIIyUZ
OPjjR4XtJV5uNWplUZ0wqHs7HxemEGsUGFHgYoNLGrlNRF9/doBgLuZDP1x1czgXTwqyT8XH3cvV
Yo9zM0FzsWeNxKuhK3EsdvQACThkvHMX+ymxhEgIFJwGmDNjGsOqKFxz2eF+UgryrDFv1PA+uMOd
cSHAOvcyUzfDM/GOBXfmW7aPx75hUxE9EIg/D6a7h9qJg55lWi7D9ROShCFw2Mfl5ZIVFCDLsrGc
rDDfXbvLe21ncRQHcQgqVWMDLNOjOfrxstlJhb0r8onWuLdQCWVyjlomOwyHEauC1kw3dTjacMZv
51v26brrSQtgHhfTYz961xqvwOkCNuQ05uwTpV3YpMN6Grkiw+BEwJzK+BlW/ZG7hOsiLijKJeJQ
1KIQUxTsmWjRKP70AAXdaxWVkjbLMJofgCaXTBfLwLJNCHBwcjVFN6TDxrTTFNxbiIKXsEOfVkyL
oVMrVQXM/XQjbq2GGzYyv6WcUF8fn3TOeeCbUCLlw+QH69K1IbNr4hsiNzXLuEMb5bS0PCrkHtQJ
KKpHJaLbq+Ns5+VkwlP5aV0zW9MI+NJNR7S1fckurWe6AO5vEeE0K5MF6pGy+L1xtG/US6JvCWh7
LIIhxgJx6Aesn5CygYqmEiVNJCEH9/iMcVhP70toLj2kbFaLL7b18fE+J0/MYZD4Q2gfxMVbYfRA
RQt4I1cvQHg4DAQsYEfFqYdzuw9B1fHnv4h/PrkIXS1jm4bfOytBDwcppRHq2CiOOl6hAL5YSNjV
g1LpV+isxjBC2ALkzF+B2CUltNdbQS98BKkRTmp4pwfwtj5ghzTh3Y5iqoh6fplehSKgLlSnMcbU
VesbsNrVHNij6U7tTToMGsX3YokNgSjtljbQ76gEkGfP1RFTPEpsHxQTTWZTEh9ZrHlMlt9A6RWo
Vaq4ZscLsk2U9fIOuA50MjyiD9UEbiuNvaXdI07ane3pVKPczrEmkv1IBvsMf4mAEqMYuClOxx+n
+fhc2MOySX2cR1BMe0Fz6YSq+NpttqLJ4XpQdFqEk9+Ifrwd+eIOK5VO4UPzWfEgDBN/tntyvil0
7WFn/4/Jl16s0S3zjS5FOeduSjIrAazMhRi2t1Rr9CqMHpAdxhRiHdecJce+ggRXbWOgiyjXhEUd
R2No9bbSAPofCTnWnPUXul9nONpoCPTAu/7td+8oue9P+CBO+NoO7SVaYD7WDxvqns5v3ANuTGnV
EBsribRrS2ZtvRBBIhjeIgQ6dGjI7fJPP4rrbiAaMaLS7FsZr3l8YSr2yCyBXFgwO4LJiDTnh+Qq
vEhuA23LoVrf5EG4WgmamkG+4GEsYaU7XCgcMAKoZ1sTfL6nDZ6WKGjyen4TTzzMuQitdxpxti/k
BEo6VFcs/2XxHCl200p5Vd3zvvt++fhOAk0b5g4S+mqgw7ithVPYefY6mTE7grPGhEHyeU0k7uC9
CZc6Pi3cmyA3YVQy/2peXsnHZvhgctaDSKVcQYOKC+bIMVyH++9uFBACcKTyavrwljAB5lu0IwWS
mSHhODIpV4v03Vqa8EFr8ZXr2LL8CpGSNow/pJUp3wTNW5Q5P6Z0srgHtXmygzYkBiW6kUlmMHHI
9BonAsgRxUyccCSK3N6wYJlwmcrJIJzGJKKLmvLFFsg8P7DFlqHOmrZax8sj5ngWlSCXo9uYsRPV
PySmmsmTqYQaL5pu6AS7NQRYPi+lfc4l3TeyTGiS27stJrQO+5u3FdAv6KP1IlO8m2vXJyASZsjI
RpGG6lHgsW4CVhr2Ha04YzB2vjnHcFKB2ZRn4TWask1y9oox2S35wWJGCare5ifmAsFmiGhFACa4
v1obfzUHR9/Lc8XA0OcUXhJN6Bc8tZt/hxXKIfjjxkla7QNVXFX28/NIkfCB9UfDgcG+ZbrdZp+2
LXP0T8K//bG1IWZhZc5De0IU2y7QXOtC18E9Aeaoz/ubQDpXWXa+CUUj2IJL9lKyulR54HPlcSXT
7Cs/moE8G30k3ojyf+rVMKtIKs5UGE8zjWMo0fjPfAmLf9X9g5KRoP3gA4KM8zSVHxJcSp4AyXa1
H3q9yQTuNkU5I7DBPNufaxHuSsr0TeTxvEq2bhFwtp/5lgb2UbrZX37fdhw0gcJqTDzmLzDmCtMQ
8ZxBojN6Bpup3oAgFvoR6Y8vY+9DZ0qEvo9iv9bHJXbWlP3x/4W0RLMFfTFCkuWelYu5Nmebt+hX
e+nxAK7qkRG7qwTB4082/ISBU29d9CU35+f5jlSqMp78ZcPnfkAwEcIX699vlUfYC0bzFKeNVPLn
mbEqxKmAMp9rFrN1idyu4kgnCOi9VN1CfTQ5J/CG2bYyyLgCIW8jb9y7KbkeQqlGuh5T17Ja2kKZ
HY0+UqdWaY138uRAaor4lxlQMAMip2NNVrisSM8awB6N8lhNcigopRrYRt4wBI96xCJ/GYsN4MEP
z5qeGBFkC0LdH3qHfI365bgsAtxg9/CHW5Lvybd05RHCqhF6Kr2aKC7j2mgqAesmXoUBkgcUXwGO
D14sqseLduJrdKeYKA1QJS2MzXpS7JS7KvZbVEZqY9aQAnE2e0tZZRO/K8gspfjWiTkBnHrkhfmn
r3nweJoInNbEM1MCU492KsbsXTBeFyNqRCtvRhrPbUPeopR6ogR7YJqGI78PcuK0bIJXyVDzk9xA
LC5bTxCI1loe2mja/XQvoMZv5Q5QgCGwIFjABxS/pnxJ2znNdTOysE0Ip0AF1234aY4hJZvYr2rK
Tb2P9PfqaDfFgtilChuyhlqT53QKJRNR1HIqTnqWHYAQV39hvWgRW5suvuzTE8re5YJ018RcGJxK
7rasmvfyDjbLZQTy+x2URBBwoE+QfjrcKrsCeh834MRwm0X5jMz9l+ZwVpmIxkhTWmFghw5RgLUd
KWPN/C+2obPll7xf51nYyioLwlUb18zkabayU0ZO6QiUY8Q3XkzpRRNDn3H8MziuV3f5a17UEzpz
gFcAqJpl2Y4OBmuXwgfEztog7ljb5LtuAJKlK3LUF2osr9pr1s4QAxnZb7gqJHILIR1bKhNjG47T
63Uk5fEYrLqzZS5HIUY9CGTItk/KN1BKRCSd90M8ZuAQJ673tWHO+B8/sY/aNjVjQ7fbEm/ZtcAO
OWoDMy26MTiHNDc89nrx2A4zzIZVFnAx0JKCpZNbIlPLubwiKHX0SUEIp2gcumBptbWjnuJgR7fY
drpTt3nmxEj7j7E8Qk93c25aEk7p+OItrxjI5tVVAs+/DSDVIJP4+FcRrodi3EG0CcshDYoB5Sop
/QuUb8hiVF8MlrTR4Jkmu/LTHkRfxboSLltAkHmXofAEiBa+VE5iSNM+9qOatcql9yEn+3FzOYmq
qMeX6l6OaGLvjvokh8QDM8FdurKyUDqny9eVHF5K/GjpeH6SbR1BM1yiozOhKQMxvAFxuUV6meuw
AHSPlKYD9pE6yGDL8lCv4N0IaHNEJuPLH1ZHxOjiyehCF82gip5fuF2jRN2CRUlPsUmth0LUDs91
HRzEdze/q4FlIXE/6Um9WbfPVUckQ+yGGekaxp0dOz1WO1yyZ8DVh4YIdzCIorlPwhTchl4AzElg
pG8K76riY/1pPjWDkgKEDKYGxk0eTTq1ZdGlulwvX59mcxuPNtngmARsmILErlOf1kIF66x9Tqim
ka0DiCTPktFYgyribNqOSH0WxKh1RCZIRFOGKinrsesO5hGYVM8B08wUuDBIkdDEDTlJfF3+Pypc
9E/2kEu3JpIIY3I0a/Z4309CTz6L+Q4fvXYLeAV5tdswTNxmv2oRFN3hTEVB8poLfG5u9lcjWBNN
UnfFGZfD/9KNkNjPaggpicDNlX13Lpdxl0W2EtyB7+0KxVR/BiJzC0l6eThRnycWZ+fYElofp54k
yNUIZ+LcJmq5U34Zugfz+CXXOS1UwDfgXBs1a2kbD5ao72jxF5qdjMvAo3C5ZOwEYZpZV0A4pg/m
ZN+9OSwJ/H+E7yGPh8XyB4yUW2Z6WMX/552j5gnbWNL1wbTychHgrA+ZESeR6+g8I0zE7SUQf2Y/
ap4MJzQNOUY62g6KzPup84qK6UGaENyUJRlO4KHbUHB3gK7ydus0ecXsmDeqvY19VVPpqf37oCT3
GsiNZ4SHjxTXJny8VIbxiCSs3ePmzbCk1utQhVq4BzrFOnevLvWBDZmFOi2+aJKBbSCbw6QMquDl
2EO8B/hG35Us3yvV67xkyz9iXaLG7sIHI4Hw/HG8b9PQaKGy2Tsf5JZU5oHDraDnVSVx5KrtqPNL
qw5d59OX8gpN/nxpo3TZ49eJOmgG9SIEIoRn0T3Kl1o+MuFizbdCV5R0CEY2c9lNo8VIeJAuPG9T
xvLv5zjXmWv06ojxE+GJSG9uJCGSD8yqcnJKl1t6an7JmeNNM4ZvsCDqDIMsTRs6oD33IahUuhqo
lXJlz6kQYW168IzqiZcL0sL1eyLaav1CeZa9sX6Ot7kRnu1vE0FiCbu0ywXCe3cRRneN4M285I4x
+Npennu4b6Ux6h2nhv3q8Uf2m+Jy//AbXd4b8V5fpykUh6PjXrmx9C6bZlRDUmL6Gtsj+PuzCppa
5czA5rA67rw5sTI4xFV3/9T8xfsYoXPZxOacEJJn6fqBnU0PAWZG1F2CV1/qMxV65/S1K1jpdG0x
5qzk8Tif5eN2CrWN9ITnOc293G+WvXXdzob059PYJRK10OJ6G7qRq3fWUI7V4R9t/GA4CmV2vy/N
4g27SQIfd0FTR4QsEjCpob0A2VyDHYkD6vaOX3o3iHO6NFjZZo5LC+Yv/PTeUIKLgCUqd0c+BqL+
VVgm2ftGYu9tLA+o6dx+hCya+h5hawHgMk8WeWO3auEqD6SkEbWUfQNeksyggiikj4+kR7JTT/n5
wCpmNcn8b/owTgWXAO4i9GXYx1Gm3Ls8TvI4St+nY6fTxl+J9StBw7KiiweOdK9WNwRauKZU1sio
+yoyO7r2rZqElI51E9T2ruz4COUnto3pLsAp3loJdnKMUllDD7i00O1NJWdPQ/qqgh/ykuxHJIBM
4FEesG6zhiQk7j0D4nPIwEG2wjbtzC0TpECCfW+SttqiphAh8LnQLSE8G+PQWISEjuC28SHFsoAN
HeL97H4tmHzmpJm/720N5mHui2VbWZnzmUn1P00UpUTq7xkUWUbflBttGc8SmR6p39XmKOKppdYw
Zm2922YKHCaMg9mk9qsIr9TEsCYmWLKeZNyQld2yUZk/FJiQEPeQlSQpIhEROjQpmoJqT+wpUFNv
Gqx28zYbyTfPim9zL+jfa8rkssWtVuhgG+Bz6i5rEB+JigO8yxkD+t/DYse3G/s2JlYlkA/v68D7
5gqeG5ZDsDjsIb/29bX2l69TaMmRZVr/decmtjtpfzvhokrQtr/Cu+O+cIvkxY7B7vFZl+BZoB7m
x17Jk8FGWE6ckMZl2sZo07kIxQSy7tbN49j5icjfUZmRjFMG+yzYiiU0nL+VZmJ3ftzhI27WlD/B
ZBr6rzboLdat7vVT41ExhKE8cKpjOEeKl+Wpniom/qXdKBcXlYe0+MLWN6yf3WuDQW38Nw3Oprfa
CjRP/Ss047KEyBtvgKlOOGaQ8XAJ64jwP+kx4PuXGB4SUDgSAuQh2yDNkYjg6fAviQgX68Xbu29S
wu2SOKExv3xqCnnfC7YyOTum1Tz61JD41qk55j+3F6mmr1L0wXMDSOg6Mhru5v5numdOtk1GvN51
u4zQlp4Is+zAny5yvySjeFMrcI+mFtWo/1hKriErLgtEvCdhuwsGr6mwhrEihk8+9D7CFdW/uZ3X
NOf5PM1dssSakPEsLPSt3jpw6cBFnl+5e1uzYHxjNLFOW1kjEcXmyJmn0/89rIvMycduowfdP4pu
VkEKfwlTKAOHboaCTeCzkjkh31ixciH1/K1UFL26P/Lefbrf/Icfi09luMi3zM14qwl0q2knuhTl
IoDHouy58IhDrl6DJL9WrHt7YipItSpIZGTjSeqpzswq2LhvrDvfw9rrLT4HnhB3pwuc4dHABydk
/bdd+qvX3O9YffUrOez0A8Np08UaCZCCKmjH7r9L5XJKr6bJZF2PaLkWrBuhiAU9GCPsm9kLkRHA
XqjQWiwApmvRoNUb0JbfrTThGeCdPkh2Kg3Z0LADQ+186BzWcVvnapoIDnjZyQjJoQ2Y7rLG0mgF
eBxiRKx2Pq4VryVU+ebHzRjl7eyXgxq65fde6QFIpa5XO4x+4TqGZg0bZ07wFjrdNJaSspjMGpOn
zxsPfy7xqgU11gOimj4U8NR8FjIFQT+jgFqXMNwOt/wy7Bia8fvc1KfpXXuq2yPaCota4PzYfLDa
VJKIPAN2rcvu3U2GwgcOQzzJJWivdU0ZBN/2GTuDpB3I06D0UEWEpqiKPsq6OSV+TGeVyTkyB5N7
ZOjIOjl+6e/BF6+8eoPSVjj8RtllTYBPK4oYCWjP8HolA/qiAlDRpPT1qVgzS97Q3mz97xFE02CP
+jeFosuTJ3SCcThofDO+i5l+/RQL6SWyD5UqPbvuWXiBMMu175mxrxJ26+Ab8KfDY2JPPHtUT0CX
3EvrPlf+pumYIVB/iD5tbRrYq1+BhQkyK1i1ko1AgNFdYXgvMgOYXlMW182BAzTgcfea2xulaQBS
1L6XuMuHFMjMstUFmW/qrfDbWgIGIi4WD5EMOsIFboLlh6p54TUrF8l6S0Siw8Ea7ky9N9vy66uY
TaTDh0eWz2ecbA/c3G1M4+R0dY2JJNu9UEeBH/7gXUYmrgJmBiFD36QWyP1YpV/NnYBO1tm0uuNh
BoEgrr+4VIPE+ge4ImqOk99iMlH4at5zi1Ej4+L/hR3J8WuaxuHe2ilkYOfgnDMi5R8wyzAFrm5+
LLcdkUZ2Ro3ZINiJ7C9U6HM0FJe2Zn6MyQM9L5faaO0x+Z4K5VJvG1dxTdpg+NX2QuOeVjv5SUgQ
0kSKOF8Srf6UT0PanuD0yQT48Q0MkIFnTxaEUJ0/kVzgtQ3+TJiW3gq8FIitl3L2v02g0/B8X1jh
jD7nofyaSWrVYZ9jjYUrKcuQ2hSbF5X9rAH4JFGMJ+vZO2LcoN3TL67XTjT04qraJvi912Bt4Yl4
qmjKNsVqxW5pUD7ufjaz5dHTIZ7UFvotjwmX1etL2kqjxD9xgec/pOty7qxzJW5gX4YIT1Uozeah
IyUgr9VLCpiDlOTlxEDVWPrUI/Wn443IE/j/WECnP0MnGLYJzWi9gXdqzfP+tASKaRcYCosXvVCK
tPQXk2hvI8gSVSOO/xNGsg4wkudrBVKjlE32WwvOb0Apu/oFq1OXQVe/PQ3d2DThX5mpvtYYsRTf
m6Egmmzob66WrIeCf9Ptmm3+0lB0/7TitFPVvsogK4mNUC4UW9u9cMGzp2ibj6M9U7ICKr5OXqs2
PzrHuWZgzQr14onmyavoOPC39QvG0y2sGnwNKoKnFnCXJaTq7YEzQ6Kz2/jXW8LHhAgKmBOsqLsW
bBrEH/Cku05PqS69gpc18tnHuegkqddupFW/284ajPlhcrXXJhKQdqR8htfI4cs3sWnKLcjgqdMj
ZpaJdwBuxwxco6qZL/jEwh86VkKsr6Sj/JxytZlLnTmfPUYr14ok64E9nNIEM6t7+ZJUZiLegrDL
JYMRMgh62XzZVXFv06M8C2Ql9T1YNdSh08qH3A2IM91sU8VZwwLInfIUv8bOzqJsBkYic1oKClxe
98ubQj1stSp806OuoaSHwaplA3fZJ+hDU8IIdqmc9VzxIfOfZ/0LvzYkuGo+2XEwOfTvobN9H4Nk
r89l3V4JpfB6O0YfPvtWxmaRatk5HZ0mtwVcGg2Kbulws8cifrPVZwjcm4QioWMRQVSq01p4h0/I
Mj8OpqL/kdWvVnb+Cdm/uVyd2ouceXEOUOb1JN23MFNKONvBZokSpe3TadSWKZlbbwXtrtsuEetx
vBU4NF/yDAV5zo0yot/ngZ3P7EexaR8vA+1cc+Lxux50dD1Ysgzc2qvvjvvtHv+kYxRF06qGVdZ2
ItgWpWq9rkuA3ALGoxoT5jCsFzYYH7QBkT1qMkBQ3twZoOxtxuITS+5DrMTul/gvn/CdZUTOGPnZ
Lq1a5yaANDbB9OSn50L4t6d2HPBEr7zgGwzWRbyTqT293CvQ9PxlUAY/JdsagnkR2RC6xT3uCwo7
GYyd7WdGEIiZv54hOwjLUfne3rse+01L+y0w+9m6Fi4k/ShggETdxZeuRmSigpTs/zQ7Seet5SQL
ZTN5lUnW/44FiAm8g78qK0tGgzwjVaAlPzZNbwqv1lpNJoa5mgpX6l4Mm03hAK/XNFhyYp6M45QE
HjfC+m77PdPA8qZmwhiUYEfkYdpJhyX6+2zYlxv7X9QTFvrrg9Es3DQypCcsJouye2Qnne0Gjwid
YJk+8tnLw+q18HF/qMN81UtvcuNnaGaxMoP8sVf9a7Q3enS/ffSPH+OsyTBPsnypi3loI4uyI6p2
gQkQQZlKS8N5XHyc+jiH5ZYKh7qiUdxoKEy4ZRB3b0XdzS7bUDWn98p0JfSzB5zYI6lya4XrMPj7
U8eUIAbXsEPjwQyzsV5r63uViLwxBgk1MCv2/4dWugDsGpikfppglFFRUlzfHtvSm1ip4js6fcq8
M1nKOcYL7tMbGb+xZyew7CB76U3M+Qo78Olmy2HZmduWJtuw+RBX/Ea7wjZaYAzEA8Quxl+3IiRA
00FRrE2W0d1vk7rsluMkJ9tICTlxkkdEkw+XS0QRMEZQ3pvDtkdiT1rc/hT03tVxY3NFwO3V36Mo
5WOiD98RwQE4ElI+LNED6QKZdCr05Wtly56ZS521KCxFD10971UUyjh8Z4Ywsg0zEnp6BRIEY3GX
bMHi6lf5aKr20XtxmMbr9MxJsY7S7qlZ9PbYjKCWUTGg8RAWCbteWAkmJIfV0h9hfQU21uKgPKQh
7aGjZKAtk3tidsgf5ReogD4nqpyf7BEEFx3oeXgt4zs6KVLEgoW6Nu08P+jK98Bf+xZ83Dl7TA4N
BJtXNmK+metdhbg9/GpNAZI0c3vJOnZWd5Kh0cZRHs35dGlLxO7/gc3Th3xaX0qSg7VX9tuL0Tqf
ApEt4wr/UYiwpU3vmvDa+NgtiaT46bUv0ZoOWkQlaN6CchNMXyZfU7fWzCmhc7UjKQooD0NM5n4l
VlJNogIByLVyX6BqU0mud4Y4uI2zmwj8tnofn7pw43pFwo9x075YS4XvA+YfzjAADjNgd6xFTfzo
v4guDaxOGiOX+XSjr5tICx+X/3VbebNwAZZynLsFlGH7+71YqMdBYpcIq19Ee5pKbUF7U6DYhPKy
oSgFxRG+vBadA/THBi4FNgRlHVyAuBzmEANFTr39fSWti33zNnDhN2j0x0Ke59dWUHPjXmBPEP9g
/NK1YrvS2PTgS2LS0WA76NMQYua44R968Q+O1kZLfR1D2VHbQ8J3KcbUEh2oaClbPpKDlLEeNF50
cpb+49DAHDZW3A+aIlhrQJ9iA6PgyIJ5I3UBLglbjKF1nfRkXhCmvI8Vufqo72rq2aLrkeIW6pn0
4uXdOQd1UHg5+qPCr1pzpjp81gj1YnPKxk88ghIMRazjXlkfoJ4MSGy8tCZWIxi+PCHr2e9DoSjd
qQB4h0FKsximP7F20+Y+wvm/uhvWCJg8IztW7byEY21URV+fYdjh2pBtY8f3FHvnoj8NPZmeftVT
KtDR0z9u1QNQHaAniz3wBzx6/bicmOORfO4ul9m/iBDksmwXP9R9lJPsyqOPHa2z5scE4/RnDjDH
OloGjPQh+7saAFUQC3URELeDipVV9QjW3nMGd49bE2h2EG6WITzl+l9/oPZWcduIO9+uyz3r6Oj6
B6yiffssnBN0M5jAFtl9YjuGMASzaxd1mprhVcTETSB7L08Mb2IwapUfvibLLLfbjT/0VTpIjQ17
BHm6F+IqWLY0nrLZ0dlcB20s2Q6BRLd5usBmSV8iHdaf8d3Gmk37R8yzqIfuuDzV59cztfpMyw1v
jWvKTxPGHvQUZyROuXJrHNd8nmKMQtLk2cbSm9Niw5Q+rVOhluplZkUcXREp2b6CMWSG7TMM2azC
gISC8hf1q/tC2MhtEliLDPb71+vXgFy6d9IAnZz1fisYLBC+Z71NOtr5NOq9qgeYkPQ3RLSf4VB1
sVocHqSvMXcWMT17Tqo2rliKm++bkx/E7LN4hZQEl3bqXirBPzN/k9AcBrYnI063LS/63J/AV/91
BV0p0yv6s9KgtVdKZJ9ftMRz6KPj+wwhPG4QydXY4KZE/6K5YoHmpXFEYTWyZFg75tktcq1t0neJ
bLDUOylZy9RMb5ARhq4kkWwpgTVM3aZGxjIpLpxLDTTLsXpTgdJXcBGQXQt3EjKjaE+ytM+oWQIE
5xOYolM5DPg9H3DJjWP+t9fUOl9eTR35uBLgHvNdv1lKPPRyRyUVSxx7CNeQigo0cbIruFaa117S
eqG8SDy0hjAIa4Nj7l+mSFwjU01De4e6nLuVTP/zmk6Vugkxl35ZW/0QFxJ9uaF4HaKQ3ftubF1U
N+kvj85xNlbe2/S/DXDDZFBLUjlHYGtxBodoedAbCDEQyxwpz7PhYa/4JTl+HiYHO7k2vIIulzEZ
t2hXPA3/Jr8CUqgYih6yUp0RuXPgUfIKoqgFdSUHJgZQL6gvYOPktUsunX19pVg8b6Hd19iNWltS
Vp/TrMm3pF2S4lbSSkkQ4hPJH0c/xltLRaNNGo88Uly+DVAJX2DMhTYm/V6HELyox4Z1cn63U5Ty
e4yJX2jQwcd6G6sN0pq9DFM1wIJpKRVvw088VIz4xRJmbaw5Dj5QpPbqBNdjPafg8u8spI/Sx5fF
sNYTmIHQVL9dT4szUP5EuAxIJvzWXQca0ngobbfdm1XZjl2z/bASB9Dl+v2lVzNi6enSk51xZV55
KgfIqvKP4A83ByBoDZQQy52wje7ihuYK86hPGulmWsAsoc52jEsO6sq6LD253b5P7jv2Zr9j6qaW
Dn/YzwyolpPhW0IVKvqJNYQwUqiE3tkKfgghTfGoqOFEvPTss7ftf000HklalnryMvH3kV6swYAz
wmhWtwfP6ZZ/8URo2hqFS3UVLZKGIbtyhsi5PvLxQXB2QXr+kUxMbWpz0rphmuXfQfgRIJjnl7kY
zJtWsTMXBLB5LW04ek3tD2RJGNYHx94S4osoOPEUJhE8YjLJnxbhCVO8yZr54EtigqcY3PHGDcQf
+J8CzsslV4lQXVuhEl/gWxT7F1hoKZz8rdrgEccWf9gvqcDG9mfGd5/Zo/gTUFzKlCSNlHddg77C
kPUDXgsFgbaJp1Nhvoe6L0GA1XU/SpQ0Dp80+0j4aHEH6/Yrzzu+D0EN5h6U3sQ/1scIyxToCk0X
kqT66tZPUnYatJpBVjX+FhEPbdTsITRBRLMPJxjh4kug0pwDJzaXUo5dAkbIq5LGwxNYomETC28S
1CGOrWC+8YprAk5LtkHORklqct9wdqEGoo9aNfjq9LvIjIgKbU6t6zMWou64vO6JmLhtSZ74TCam
rBQRqowyq5v6DyNVu2tYEQMZvOAyo1cyacQtL6Jh8HcunRULznxQRcNzdZ+bTXzkAdTapR+8aap4
O7n51+nvDkD63P0WZkSE4pmBH/MPJS1lSeZJHpdoWiuPPz8MYamQq3mkWFxF7BrZ8yf5HI/CZ0FJ
hHqlXNYJr8MdOva/qou60+LgQ9L4LYPhmAr+YuetMEc7F+p8UHZ/GWb/2jEhTNItYz/IOhqxiI6W
xWg9qXOhq2kcQ5kKcTDF+ucdS6TkMMeFsA5QjpBQIHdm3j3b2v7C+L+chaVdNa7Q5ZW5zdUVqKGD
ckf7mnN+GkF+ny99teKTtfYbP8w5PQqzNrjnFoUppIY5NoJWqcj54JK2AR55UBsCXv8HM9bKCGEg
LE9dJwl8oREnc4E9NDVImO/AVwYTuP8nlhSVEeA2divTQPhO2sgWnG2LaX37kbX9KDlO1pcKcECX
gPp/NRf3/OTm8YwVs2QHBHq0l/Bu/Wzk/6rVQgoYGoE/evky06giHmhm3oLVOuLFRp5sPKpeqJI/
iPLjp8n37raSsPZ5H3BfOrrYPfBNqjZANFVqh3Qqlzn2ityXAG9Satox8h5zTZ60vAsYV3odOuJN
a/xK0v99ksxdDx2G/x64bYDZ8VGmubs1mcaJFLALtyi+L6MnVTWtwcYsgpwseJDAPja+kcEuUG0r
FxhuhZ8UM2yTufi1WvadNthaDEsEmv9moDtYusjWkv13c28tR+eNr8XG0ndWVnXtoL8QqOjKdTZ/
ybQr5SB0L+CrqDYK21PVW1dg38LW5pfA9BXg9FfqL2CXLbgcSHRn+7gDaTNV6qe9sJeT4Gsfaa6W
d2+ftbNTsb7WIKJ4beis+Z+57KPkq06AuggaNFVfBI55jL/62Ktu4hg26g9oBRYFnV6J6Q3J2g6h
0rHiQNxORcTRclZ9zAzanehfj5P3Cxmap7q8eNpZsGpF736GjtWLAVkBkZzWynjySfS+SjaZYmta
2SkjgVobL31/0nT83Joaq8NxaWlGf/VsNFWPIvoHZBzCt87jPfNZaup32rZBwtqMxkRtyhrih8O7
rdl6IFhtMVmbfsaYPqbce/+17cX6FTb/k5Do1/Pk1bKnOyCqiac+VKBjIZa1hVmtIAJcv29EQzSH
mtQ50BFBKVWembTN144nInulrcl2Fay0yV5DgU9u+fy/P70sVvGTNgCFZp54KO2EkeZUkiDX3yg9
olEpGEIj+u+WC6iO7EH+DymarZKL//gutcZ/hCW2krEvFStqhf3GJSiegsIk3ljR4I+i3QSsuazX
vaNt6OaNeVCNwhARJwpZJlE8QdG+pD83MIYCKqHyVeMpR3mkamH++s6S5vxFrRynbJBRGdwhwRTB
ca4WUk1ohdel1+stu8walYCCOFdIKW3Pp51dfoPMyoEpvXzm2SRL/TRtZeZf4HQ/2Ebb4CMG61rd
EYqMLXEfxGAkqeGnxToUj0mR7vjpIOcqfqxUJn4qG2kv140/wMzfEddRcSaU833uioosFuf3pzHr
HB0783IoO+knuNUhS+SFxLUGwvpCRYnkCC5TItZZxm9lxRy5vi2QPmpO3Bx2HzTBwJlnpGv6k0GX
e9KZbFG7nqyFYX6vUNhJ1otRcybroRzlc+V2vV4yOW6DWAB5fi84rJxyXkxM/rY3jThhlJUaqJKv
8693BE4sARbNIU4V4Za/D+vLbOyI544LNa7gRVBHUF+vgj1laQWcP+OaBJXUxMzGmJBlVEft+4pz
hGID0Jtp9v7sTuLAPq++bEQmzNaN9NN7ri8rSgeR+Pp2n7b6/D0o5yziR1Aw/1YVap2TeVYBCYVM
EQT023Und6DZdK6/b5uplAj2E0F9AfJhq3kFnn4EsuwCgWko5Ou8VP0QtZochPod21nUpaEHLA4b
s9glk7+nuKS0TU724aEa3ykZz9SedpZJBlVZKvOu2jgBfKC7HJrD/BOuIgJU50QBe2JRrr0dcU09
cwZMSIXapJy5aybDUsjKsgRRA5XrPVdEmgbAmXbfKt4HKSSbALbVuw7Wv3ypUvcu/y04JcRmbt8h
Upd6iK65yVoFxlsi/zaXAZzN9FM4aDSi7P3+K1JifUNNOIO2Y6Kak2kp/7VT7se+Nbpv/6cM6iSA
VqGuBCNM1I1iJDVzLXPGoLD+85FeofHLa+vQpm28JYcLDaGC7/FkzhnvXuLGzIys1b9LvlmF3YOU
HKyfzaNq3NOWsdkps5axnp1B34YyWg1bfEptfa3L8Em0eW2DJEpOLYONSbXhfOLnUjjPK4L26GMI
QUln2DuixDOIhL80POuRM+pOCByOU14kq93RFVZ6x13hjJEYaTRt2kbJZuEN1L0HhvP+N8kRJUMU
lOAfGI3iHhlPHpGkbfMAmqDIWQAEc/vohbss9fdpQgyiHa6OoqRyhKcIrpVYvLkAy1vUplo/nTOd
+uKvrXGSsm592F/42rGWBox5vIiuM/hRnhxEnmT7dxv865eriwVjQYMo3p7wD7rXTswLheJqERaa
kPLmdhznqoPl5LHWIKPxWaxKxiBO0g377ROK6fRfL18yMDZ1mZB31YrC0VnMmVIcQ7rwlTft6VED
6/aQhNa0LqDLy+Cziq16sMxzcefLzoRwnP9olr040PJK0iR/pRHibF5byB9c4IaP+NyJY+FJ+Xka
R1jd8fLZBqxQsxRT5wTO/JZQqOOfhJvBdKVXYulQd12yAAhglbIiYX1OWhWvVTYH2Qya9OR1SOAY
XoNH4LPJoc2KOkzhYZ/2LMLR599xBn4haxDJdlKzjhaRLFHjXdWjNSPCo+kD1mJocaT4iByFrVmt
/KMaZDLw2D4gRjgkrEqbWpvhjmporXne5vzeQg6VfVfqCSR9UEzt7Ljn5lai+F3AaAJfOnVpVlUC
fXfj8sL2FcavcsTxC8SnQp1p8mccHDJ5itbTdkC6x/4FXIH0MzibUwVRuxkQ25aozGE7i2bt05+Y
ix4zPM+IYkDeiWnR0qZb9oh1M7HKE8Giz1XwBKxZeS48ifaovq2jl9556v3YEes7J+ZnEoDeNpsw
fYw1I0t1qpn2ZWFgrQQA96XIhLkM3AVX0C4z3fhxoVW2KGTREa8Xcd0aSj28VebV7kN/29mbJJ1B
kAuO1CyDaR1QiZ888lPFEvR3U4rZ7SGutngoM+2XoexOVStWPs5uAaUPHaWRpPV/5SgY6D4ScfNy
iI299QqB3/pujZDbw1f3tOxfO6EJhcUinNATlzbkydg1fcx+uhcYsz5dwQl3roS4f+QKKufDhFGy
qoY7bBCQT+WWotugQL1Ba76BpjDqfgyFvAj49oxwsEbBmH9tP4dvN/3WzRtA72UgtOhxOVuNwTjr
hH8ouXNxsCABsu3S+JKVEcdqnb8EFk/xAvOieFjnAd6tgQySbvGxYkYnljAP81amQ0lZNaC03Xfb
Mivpd5D2PLBA2ctdl4lyr6jU/u9v/aHkU++hNlpxK9eG5hvI5RZfq1DiH/utUpHMkl7JOfvRhGsi
6azCiG68ccsXga4ZEYZedHY+GRYn4Mcujbvk95CoMMTkdzDrHdQUxsKJGY6YmZjrbgKpi8PhWQXo
N9RXKPRJM/7kmK7sYAimrhdD8Nj2V3sWyXLDspbNG0/wstTcifQd+CNU3FK37y3KSwJYksG2gbhv
sflNQLPKauZ2+EZ3vqbMlf8ho5suaErMtdDOVzuKb1j1o3CE9CcWFKiuDSQZwgyUZ4xyM1mA9mOy
cVbvLWpaSzTTmau+OJ5a/mRS7TZqGuf6mayszG2W0QEC7F1lksCfsvdOBlB0EwkF5rPwcNwgyO1y
q1lkewKSUm8/4kE30S6D0XUmiQx3DyJBBN5BEnxbf2jY3JoKxDEi0Wv6YCisCt2KGCZbuhfzxbHT
TME/GMyqPNrqlQYO4/74g1/X3d4WGz2a0qpi35roe1MR37GUwK5cW3SoDiL64oIgjY30TN4BsBGL
ztsBUMcuiBHvTUdR10sIPfahgNyUgIXz2ev2qla4sv1ZWsyCi9dwqceEpE7rAd+1Fprzy1NAlyIW
Yr/yh3QnzuEDKD9V+WRqgn320ZHZor8o58Jb9o08Cc+Dj8k2SMsnrOd1Zfwt1a1bQcklSwr842Bb
bpZZs+wQSHNgA2sxagfYWlgFJSk65Ti2mzJ9S5KikGCay/x9rLVgJMDmnd7luB46ecR4qaQ1A/+P
rqj9NSOS4HqOm+YY41Iz7tcHeJhS6d0NudWFYBAg6kg4Z7DFpy6TgtIsn/s9v0Gw2GKixySQhA5h
qW4F+imohJkjdX6hYxV4J07Z/uyYE3Ix7+3s+iXeFznVpjKlr3pT4BL6dmKVes8s01ZR/auE6dp1
3Llg2R12++3gW4fQ4BlofvCWkqBSFWviQIHJ5GngToLzcdTurEWBm6VyJW3nQlvhhWuOIGQPC6NZ
Y5oj6iP02ni8wgbVhe8OQ3TLkiRu5LMDdPfCDgo2nsO6P2vMGwN9HRINIHv5G8s2b/66fC0D+opl
EKTXKhJd8deUOhU6x0RYbigm/IDBq/AL9lc4/ieWCJmHrv5qrLE1JKRyrRCPD0ZTM0fv3ElkDoia
PDKNlrbJaE0u5IZu9sqzu1vm4lFzg0beEMWJfiGPlhXhrqX5OiGqDvD06va8kvLyOsqO8c34KlX1
oYlZmroruHm4sb6LbOMWRxdAmd8nAkjxB7UlJOJyNm8+wGKR+FkQBxawy6e9lIYDne9NQrshhKMK
qWFelNb9Lt26ZB7Dck5W87fy17UG7vi7k+z+l91b36KDsdu9WVY4H6Sqiyy0tD73aJb3oK89EGSv
/av/dcMjLDzn0S+nTz0bWHxud+6Oj6RdPxHipTx1fpeDHCBgW5NN0WfqvbMD0tVsm0S+diQ+/XtV
TUHkEb+/3z3s+EzE9q3/Lhz+T3y/R9AEolzEzCxRVWTloQx3faVy4Z36IBy+DHs/tq8iRMa0jx2p
a+TRb6efFMJGFiwR+GfIRuVKaV4N12GUEgNYQ3mulryKMvyeRdzqXcDzeaoNlvh95Sf9mAC0cGn7
bq+chC8+4VnULo3NWl6JC4xRO1eUpraBjGbOpdrB/tc0YZS8I+AySu0Z8JsijibZUboN8SdBiHvw
IoQ8HCSzk/enbi1niHG24nlH0J89Lt7mktkkdGB6lExOFs9Pbh3CdD6S7uwBzR+IvZOmG7VFC1+/
gIfDWZa8AVYDW/pSOf7OaVGBxIXT72w+dFNOk/twK04u6DSxzNuBl6xmXMVpbv8iuhR6UbOuuARl
/WAbHEa911xGg2AM/ID/fdAZwYnyVlvcXyr2vfKqKo7yx9DKAoffVWedPAEifocttZQNJNw32qKF
7euGJeC5COGEix/iWRVkuFgRcLXQHR11Nk2+xYTWNlicBoW2KSycUA5B4AdCPKge85ojYtS4lJDi
f8a+C6EohobGRKPjloVpYr2xtR9taEkQ3Pgt7HngrTHUPqtVE1GdlHQ8BRUKmD5Gy4fRPGM5bZm0
8VP2edbQezaCbQ/+eha8Rg88ZwwaA8Dz8L531Hvyd+/mZVP2rsYXpDAdTZ7k8E9F1Y639sqAgZNc
FuU1NG7j42glgwn2ndkQLfxaMPbkP2phZZjZHbBRbvhPMWx8oQj4Z6kRiSuvSPymGP0t9vyBT538
CdKRtqPaeTIv50NWmx5BDSOaavRtTPQ2qfCDvUJMBA6QeN3uYOs7R/HRaNVjzuJlgD+U8oLVKZNb
iTj7M2J7dMPi4E9p+siXih/axC36dHsjRbUKY8n30PP+gJwBPZLec8J13jBjF/uDvpzQKM+bBJOx
aFCnmP9Pr8iU8wQAfLgo5QMNgd62/LLfC5ty9qISWpkX5IU6q6xUslBhQZopvOSlebdjsqtIS+Mx
6GI49sBvtcVlWyT9mwpLOLFGsJfLlhzNgMO5ojBtN2e/Gclpk8IjkrPNFBcpcNUbw3u3ZbnkmZ6s
PPnrBngt6KRS7MKPqx+69gp27TNRvS5CYvWBmsaDvAn/+aAL6Nfyi9dBGIhk+g3/MQVSN/2+eKTV
UWEepTO4SPL8etMY90FP3Ib7cc+RQs64kmfrUCrWbkHZiTK9wB0vyLnMRkCdaTeYFfddwG/AqAj1
uWJgGcJIii3jNviYlXKqrmp6JJfzjxe/TxzvOHV1wxDVEi27zOroWb9XKsozrV76FPTc3UCFgKLd
qRl/sNdfAqQGlNFCy+psDLej5drntKX7PuT8Ouco8jILQAfIxPIrvVWdypwCIWgLDfQatoKc7Edk
7XVEjBdZYtpKAa8RAQ+sT/ghcxnAkkR1xCiDDDpY1MyIbw+BBXp+5hzoh3oIq9JX4TTx0nWYpGvC
W6jmipMeYOwpT6DKT9Xxv0Jv/yBXJArL9Yip2dHXdGWW8zWIyesSo/oArLHdXtzWV+lIcFD8TQ4d
Fxjdqy3M5vwcCVvsRTkvNi45Hcd5s35xl8IEbFhTetI0iA7zSTxDhOP0gvi2ImYEkQaHOtm120oQ
aYFG5hrCsdYrT/H+XfGkuVJaAxwv8tx2xkaX514ocxO1QJxfHIG2XKaYoAllOasv5eLX00VK5SSu
N3j7P4qICOERMf2GNLlyx9V+mbZZ0vzdw6oGqZpv2z2An3l6ZxH9Nngg4QUQbghB5YNuqLVz6R9g
LsbA0oQBA/OAUJ9xUlTJso+ZCLm7fhNnOLgNI58lKOUc0OnGJ/ksdEVuvsGYSXxFV+pIQb413+np
sCWu87YL9hn7FF1vwAxaDpEcxJ5qbv6lO4Me1qi78J9OHCugC8EAzUMxLbdtWjDaA53s/rrkxpGc
GO6aFGH6kfBtBOoHNIxlB2Rl4wpv0f1Nrg/gL+wjMMNy3YHrLMMkefzhbRXe8agQmpFGyuYo/0gi
8jtJUl7/WNHix1OadbKZb6e5HhOCDBmlh9T+F4zPP/ivhGf+8h2bn+k6vENCHzB0LzWg8gR5dl3d
YHWSJ25yW94TK6waRVb4Erd6wvZXtz95h0K6s7b8g+9WfvldZnZOaKRdwXOm0ab5m8vfhKzfTLSW
GghB+8ZGnFh0jjIPhWXYEjdGEHooCBhb9+mUOb17YTSU5dYmQV1Fi52K4ajsWxVs1G9rlS2IiLoD
aCdV/rnSyYWS2eJBQt1UJISOtRloKgPJQoumhx0BLuJyIlyQvawTN/8VO+1Nf9nsWGmfLJWxondw
QtHJVRO62OVZtzPhpr63fd1wmvffpG9lb7aMJTXg8klJzBlr7d8jZJ3qoVeb7sfGrT5k01TJE6p+
kiPlUNFOBVJBKc0T+IpeXq1JnEkKF0OT4YI3TNw1lLPvx1EctJ5BxfgvsLGaGuITmNBJuvD7zXRq
r6mZ44hZ5OzwhOjREH68ED7yRxYBy7wCeUdkOdG/OYXEBDLW628fe1dffpxNgfKs8kY1XLCEbdfY
F8Bhq0PPmJjX7L0GkCqxT7vqjneXJUtqcFSKuYJqSFwBP9/hosQayzlVo8hS9GI2be5ncBlg/Dn/
vLB8h81mDpQpV5kyRhw/xk9SJDNmnW8JRKrWL+uQ+Wl/zR2k2o1ZEPNOQsYicfgQRjG8qKp1rOhp
eGkFUHbHctbMJlJ/a+lkJ4aGvQ2BCdGmh+kCrk/I5bZSpsYl9n1mSP1itj4MwwU/jgT6mDn1GB8I
L5TX+AqhKVRDkVk+M+AW9AhNFuMOq5O4c5QQVJ1zQDD2IEdvRNemci46dMUe3wsDjKE6wmZQy5IU
Q+MmGK/HEUY+yNHBe279VNeMA8Gy7kOBTKiL8mEI7zYzWJE1Vu4Ezn4evzU1X7Vx25G7sS7xYMJR
JiodyJ0+Akhdb2YZlFxEIe6eNrbD0CLna28UZcPdXGoLQyM+4rQXILhzqaEezq4V0US2HBD9OVpe
xO7YvHLU7fUl1vPV/cZsmaLbCucsNSeR7Lghubn33f3B974Q5WBSMDLhQmZ0Foe9lhESS+9bAdwv
QSZFU2jUKuX2eRqbaz4XErUVWeN2kN5BuUAMKmek7Yjsip8q1El9MyIE3uB+rMB5MnmayH5Jvw1Z
6YgWF8fxDrDCb6v5yRfcHRLmzcbMnQv7roLgctVY1A6g9irvf8gEV6c8lCC3OjBjkoGhGCiP31Dc
AzGtjfm6XGrftbQl/N4ixhTNVSubbdS+uNnX78cd5BUMSUvMDZlt0GqPDOFGVsBD8TBLxNch8Ckl
l9I9ycTs2+RjcYl6vwNhj38BnD9rJs2FXK1bpt9+zL6q4wGS0/sN3hLmorUwpkx1tYsD4Ts+sYnX
9YcwUPCEwoeZ4F3PTefYY559zZvMLMxtRwOBnSpCDSFPbNj1iqkB42B6Z/G8Gbr6XX5A6kMvjBq+
ZU62Y7LKXReOuK7M6VQBli+iFAyd/o9nY3VSKMr4mZ0j746Rj+CsLVAajz0I/ImaLbktbGCSJrtc
DS5lL0EwmYhXNKfmMM9AEQ9/DB0ig2jr+rBInrSuQOjfS7Dm2JiYgvt4i0KKIEhrfFMtOvJKsTzV
oWDHJRQbYVVJfea5l4Ma8wLkIhF96rl9pECX/m6FhiMhxf5el48RHr7cRm0tIVhaYXUNF8j3z43v
pIyc532In+eZkNXr2hA53nrDMsOxzqV+tVlQNJHN/oCYIR63TopnE4gyn4bpfocCL/zCelAVw37g
PnA3ntZAOS9cFxfYDoTng5WdRn8VqhJf4lF2z1D1b/sx/orJko92nFISCF8pV/ixeKZATdnR2St/
5uxIO3ol7ZPVOdcDkY7kvewm5n81s0quPbZEouPtaatL+1BCmpO//Ld4hjyAnsb1S9EkGq+paWTU
2FicKyADeTci1SOGs6XbHJFrpIjUb/Iq6i7TR8Hyo/R4OyRhxpUjhVKVWZ5Unwdt1C/wQXNVsqYW
8xiwQclsxi43ux+OxemPcgwzyFVKxdLN/m5eMmTzKupLMXoTnh6pS5yFsFT2dhzIL2OC6KLmanfY
51tK5vBidEXWsHkdz/GPiA9ZK5SqpE4DJzp0v+oDSmImFrBvpvq1HH34Ku//EnkBWbvQ36qgph7E
nsblZro0xpA0iUvaNE8SDu/CHsNA6pgqP4/Nl0Hw7Uwcsf4Q4h/b4Jgp6rldfuUdNsQnnBUyGsGN
eQgaE+VymcljVSoYjvndlSf+5b4XyIfbcXf0l7PTg+BBcZ/WVu1jf/uWnY8I9X9Svf7zUkZCYwYL
tZ0PbM/gIvF1HdREaNKgwKovoNyNyeFQvwACzclM7jsLQh+mlT3tdeyukumX5qPYcYOoP1EHq/va
eMHLOHDdqTfXWnc6fmBFeoF5jN/5Yaa37G8Wbcrvh8PuzEdOtOu7lzdASmAIPdued/Q6cISDEuPI
qj4QkkDVNSvx5OHJJi3eUR9mpTzPwpglGbmEHJd84z0a+UpznajKIpaOg0SZ+g2sT1K7xhp71WXy
+DxDNnNL3wfVxx8TT0xBmdtsWGEFkk4GrpA6Cg2J2zybiwZIGaF/B3YeI7QKfGGetc4R6sHQ+WLZ
QheVPI163ipNQ31gUYOhiCYGgwNUNX0PT8jBN9q9wPL/0vZDnF6n6tJKs3P2s80W7lTQHKEMW8iH
wYoHsIY66z4SFQQhCJHxQ+ZG5coW5ZL1D+ae+r/2TF815y56Jr4kk3F/RG6hpSEWDlZNvJak+WE4
3M6ziMr3I9IYHPb0z4/3k63xdg/YhGZSzYuo85T3MungR08RdAkrerlChdcCF9UYX8ml4fu14d99
i9ZIosGUDbjMQ7mmXezlogPZEaGHS3xhuO5cUsdnhvMQHs5BjyivvMgZqiNPUNjl/ZVBz8jccYhA
3xPpElx8w1zVZN4901opO4eHrQjv3YQ18WjtFLTUUyuKfvidkcLvGPsbr43DfLA3WxiDe/7WrGN5
edayy94iO+zeV3lW5FLRfStSWCj8EU7MW4yUMn7JQ4NxOBWax8PDU1VB+crV/3eNbX1DlM3/zCsj
vK2oo/VEZLv7w2d3Qn+H5q8JHAHRhLtd/jBC7UwINEmKFx5C8CIt/gkEVCm92vREn4nl3dlELVXw
QWzZD5UFE/epd03alrMAj966WIoANsydbqOUMAfH7t/mQeRFQq8dOfuWK5wSCg05KDvScbHr1Uic
CCraR0l5xKpXCuwRXnXlFyPLpXXIO0YxO/pbp0I3sIyj6E1ja54beHENyYX2qwi+S8gQbf1b+bi9
Mt4d/UgP3Qemz1ISeE4Ldi/SQr7yegF5i5ejD7GEA076qivKula7Xz/xmFtYajSfRz9tL21L9khn
cPppuYA605kHatlsa31HzC7tnMYb2cnhsgNvRgoYG0pZ6xltS3AKYNX69xh3pmrc+R1fNvkBBmXW
e3pkvbgOK+piA1dHvV7p92ukFYR6BEK5+H6qR/P3F916ve0JBQm51/XvH8IysSE80qLteG/4xi59
aiZwp4J+ohF7YNqiLf54jEAUmzWl584jwHj1UZnZsdpnY23iYwu1ADPE3POfyX8Owum6faE+cMRK
SK8y8xvrl8hZAX6Vt8lciLIBN4S4OYn7HjiCSeXqy154LZXkZ6LPj+wa6KF1W3PkD+9JhRIqN37D
TY1l2B0F8UudwjMYHJCm9o4g2seczkI1Iph2F8jMApsOKgx/d17ucCC8Hp1dNMU/rLTeuPa5pGg6
Gt77Di0uOuVyqMOdzbhWG+MZs63nZQQ+EeFituqJpIcUSTOdSLBW6leNu7h3OiZggpL7EQpj8JtM
PlBgGbwW1ClgLFraX6lW486t1uYWAMAOfE9QW5ECx/NgYE3t/h43RV6dlIMl/zCsn67UZV6E0yiE
9bGkZtc7LxFXZKGXHlMynNgtA9Cf99dFbm8MtrTHnsCcrmGtSIqCQMfBsDLzrTjyycXUY/6GsJNZ
Fv9TdG7kLyJwgqqoOp7P23BcsBdCKO9GPnL0pB410jeL+hPf8xOxomY54QIX/uLMeFpDzPbZj9he
DQ2RzRcVfrf4IYhKqiGa3m55o7B00FbKEdPWaU8HUBLaiWqoUcXhKDxIB3i3nKn2iMiz72j3BEqi
+vhslICZiiMfV2A4tss2b66HgYMb7C0digxXPjblULKHr7j+uxFa85Je5Qex2ORYMWx8eJ1clebs
83/O8OJg4IYi7rnjjGIVAFgPBoG6bU2k4DN7avFexQ+AkBtUnBdYRhhedZ1WUOnCGWKT1z6z/CEZ
vEt63m60UnF6qp+LXJ/dnc4G4fi1yToxgDIpcZvTU7c+YK7GcCEPNVM/evbgMSAP6G672Z6mqXRD
2yxxdlPia5U1FFJhTeLOe4GOkRul8aysJ5sBz4JhcAv6nQT1v3JlAE8xiFTrSpm0OjBKA7ubqt6v
6D9K1lQHgyC/rQLVxIzZYgxt8D0exnfT+3G1qCll6cMI9Z3b3syWyaJJS6tVN8kPUohiM2qiacaA
sYBZYlWDxcGkkqiN+7eYPBakcv3bCZnq+jmoNRPQhpCXrtVOBSPCYlIGosJtb6gFiyQ4G9XtXFKd
sxedG4a5rr3JUwtSaiP/cIlLnz+wvC8PSuERmIq3D4fv9P/7beqTDJmfv4pdOGOar3h8XOkEjfjd
eNC59Tuhikn5wWjB8ziiZdSi0/fVXQNBrrNDv/4nGGzvqRg83Z1v/ajm1BmWrn1QgBN6oE5GXxDG
Ff2CLJZXOdthPxhjFNTwd9gd65kNmQYrIgusbvp/Y1YZRWRTWpwu8iDQCQqmb3hyCGyLh4/hTumy
2gQ8xc/t/0ZHqtJTl0ibp8ENHkvO67f6PZIyWM9I3RG2msnfjt5+6Es6JouWOYdoFB2lFQPoV6zF
/kMBWMyQAQ2ovaCMdNFiuqUA6Hxfxe3B8o/YidbY4T/nY8u7P/kNSwhSWzOgOD8Pr7CC+Qrq5qIO
AxEhbe60+CIg0pyt3FssCtK2P1NtlQmSfl9o9d+BSIzB6Sqq4OlSGY4M9+wVwEF+IqbzfYAVi65f
IffFoXjh18ZADo2/L8PJu9QTEW4i3zXNzVQ9kKlRUhLtslvvgtZbuu6U+L0VdIWSnyYpy28sOPMs
cX3KzinvL/E7bgMizbxcqnsPdZdbPtxsLvOJ/x1kWhriyd1UxzgmR0iXIjMyv089x1CQB1QpBc9o
XOmQpnITnXLSG6IJm0dp+rFPpcNlSEJcCr18y+k4CkYUbx430YlLQCQ0tsVpEQlKJCcOzfl0ip9o
q0+phRs7M3WlZIb6yQpAVDNEAD8egfYAZRDmfFlQIeuajrjpUBHo+grq4C9t8wUM8488jYD4Ge+C
ffHs8u3VNTZLHGJsWXEuiAJHZW1vkpIvh8ow8Q1u9R9UGAEY6JQS8Nfp+ljmzdbjjv6v4QKynC0a
0brdoAIwOIirTHTA3bk8ee4cgdds5Q43h/NJPNGpV2V1QVKyLl3ubNqKip5Enfmdw8i90ADYnI26
geSf2j7dMfu0Uia4D4dszOFkcVRx5d7nrgn18QXZBFMeoyeQCnQ74PtY6zVTjYD4V6u6ZIDtnKjq
68/tVb2Idy7vZ28U3FhUNpES5HSxIDbt8MGfuXCywgaq1vatFQe1rlIBF6lC+17eZ83D4S+1O4g6
s3FGTBYTEVmee3c0pf7eo5Myqt1nHohWFt5MsOqfTSb5k6E3sVKoXHeKTgl/Kvv8K4NOHrpb62fR
kTGN+tJ2n2P0qTefqzvablYFgeDqRux7DpbZGHm64Jggqs85Qdn2MVGMpitOV7ecbNqp+1seyvVE
chNdO5meySUOg+p9suabpuenCN7Bcxml9mT4Ss0CLCjLmOahcKLdvQMejcopxDb0Fu2Wfs5PFIQl
FMWP7DMZQPY9oAp3PGTLu0iAiT3KNaoqLVW5BokdBeExEAZrwgwKBuGZN+Jg1Qf3LZsy2gTrHZsh
ngBFiVVMjlxBuwI7b20pCqznDJV7haKnPSlgSQiZYb2QGr+mxVgpIFZKplYk4bAQEuLU558fr89G
zjjUGS2o29ZpXQnxbio8RFIhVN2DJoDzes9HoqKC6VI4w/BmXyV1CFBMGv7gbLSYRwuSgAhfrP+p
GsT6WytuNQl07Hdhz5iubCDv/mnrOM4fwyRGgjmK4tjACdSjn2Z3NiM5wvQEYV2OeK4QjjClVmEb
QaLAxkNtd8IHpLcGBR2cL/DaaoI5keDAW1HgOBZAMIdA7o9b3KmZzrRg4RoX6rGbTn7ylOUqtOcp
t2+QkO8+qG6SZa7ZtpUgHLwCDGTNnDogkznH6DLgTpFDytO69fDkb9rOWFgCVZyfiUp1tmp9bbb9
M4h4jCCEGTmlpU16qS7Ujz3RKvWYRuyy/8NYQtqcvkFquRpUMdrD4cBFsfaKazXQdW0S4KC3xpBp
fLnLsjVD9zJ0nG0NIDAQiZKq3Qsw/pu+efSCbeEkiTWoHOh1tvgZtq2zDSQsoV1xI9Ceycdh6l4p
fEEmwFWfxpU8weKZsuRfak7bl3ePkgudH7Z+sbctxfBSi6Xb/NwENp3F+ldrZSry+djCDyz8llbq
4WVxTnFNrXqzTN/R+pIPodtKJYhFd4SFXqrJlWi/1bxXmOyfCyZk4R4Fk+rToXFcVUBpv6r6MhMl
QVBsqHjdhUCfOoI/UOB8tR8LNE1ZT2NsI7nxmIkbhQikDxbyMXoWRycKSBbSDuWLqE2Yf5emHOUP
s7GMMo4ck/dFJFG4oPjhg6skziTet7BcRz7zbbJbxXOqekN/rJjtqhmPPx7qR+bw46N9ra9qC/9r
0YejHoOrUVYnZXWBOvSHpXrDuV0ui7hK4Lfaz/+oZ10560ddRV4tin0AGJ7jxj+yYcZlFmo65nib
Dj5+HhP2FXK//Ci2G4ISzNA81aBF69QlD5XoMtLNRktKk7bZp4OaDsm9nSMWQsOJciUVzz/dF68d
Pqhr3s5Eesz+tG6/kJErnduP85xLZFMvyormVzTyeIj4yhu5aP99P4UIqHq0K5R13rbsbXCHK17x
jJMBdMaKf+3nF0VT1FSyfoXKHaJZdxcVduVYwGlEfZCL4bM6jgpweDNws/dcWXeNBqURHb5xoNiO
/yh36TW+RiKtlMwieUKpLDSZAZR5V5+NNoTY1FFjpMjnKUG98nISjh+YQCpTEobk4I+TiXC6ZAp2
X06To8ijtZpLjILJ0J1zjH4Wp0ybjzVgZh/C2XVR4QbRdfXASYkK8f6p4IgHnU8gZ84Nz2vHb6kb
uYRF30TAmJPHBFzIMTnnunmo+2qUKNPILR7DqdvHi00Okkop8AGf8WlwQfqlGNjZvIr4eGivOaZF
OLP9lrG6V5ottryBfbF/v64LEDTjpbaU0bgWDBlukKWgJGaw5x6g6Z4cfD2sSAV9aXoXisQ2gaQz
uvMqLk4xCYvkoqsW8R81phfuPfJF78WNboCV9wecaPG3XsicQz+XAVBFIzQ7UIGh7ALZw778Vum6
O4P5Bhhnp3E01B+sHHcoSIvpwik17i62yHdnaOYmbBghiRM73HmjM8UbcJBlCXA6c0TFiMY3XEbI
RKsEbpFbKI/y0zF8LMJAYxUSU0lHFIMWjktvUc1SbHp9uivS5qF4DhbR5/4m+JiZNaKARXu7hQt7
NEsxzlWoZ2EIp6AUnmpZJ5nkTuD+E9Fbor+3sXQSbV0GzqHxx+53MM1BmAb/YDlQupXO5sr8LELY
v96PzIwglhI9+HKFeX7WrLcWpLQUz1QqG4ZNz/7oi1vAhX8KUZLXQTWtLzZUzl8VLzrep+HNSquy
lO7R/f3wD+jCNxCVItAyzj0Pa48MTWo3OQ9VUEaNE+m5yYbkj7N/91/5L3EXXq065TZjGNY0L/th
vYAMaSMhT8QZGrF0JtYZt1pr/V2suPr0Rn6U8eJrgBNnhVaHp0iqH3brTxEyMllfrbbRuE1sGOtX
7dxRbFHPNkrVL+whnId9z9cJ571n0eh6t08uWUqYIwaLdxZhpyhhbCcjgDZeWzrSvbx5zyoYPIFk
54Q2n4TiWObLMwQsTkrLYe68aZlPhoQpeDIQ9b1AeZ2rGb/KfKdCiJWQYWmVSEeoHULRfX8wsfMg
EbxOXB3vIhq+BbzGQH/1gFyTeLPP9aT/BrlIGjDQtOqUvHP7CVRNZUt9Whb06hHmpdJNICl+dDEp
083yHP5deY56vRuCUkJMtT1FAckF+lVxenX7VxmcNznfom/ljs3JbWfvrX7zVnLPy7hZW2yFHsMr
wSKByHQEMsJTVKEYkgIrvthngYT2lRQnYOG42sPSuND2gdwuzwVtAL6MVo+4kk9Qlb2/ofpI5VD7
QI4tuhrDT3aZcRn1qcoGkZR+D+SazA0BwIDW1eN2x5Y5SYumZpN6QD6pWBwHkT8nPZLdISzVkcL0
a3AySGJK64rtQrs4002enh7yKhzYXF3slFqYNHzacV6Ir2pWs3jvAVc5XSW46wbTIM29wmaIqdAY
DOtLRLfXgK15qIMjQ+5IJTjQRE6cA8Klz9fj6B3kPVjc+qfFSXOKabkG5ol8WN8Gp/sC8k4ru2J1
4I3g0RzxFm5x68cmCyTiiB1Qhw0eilhcLaeJ/Fk3VzlFMRanE+qh1DDl03+eugbqmvK4apMo94aT
V2ZTSMGNm3YqHi9zkoxDfiudHDfavymnUjn8Oj9TTrAwT1C97XecVGuhvJl2nVJMpb+I5fGq03PC
WpXo+U6wZPJmL8DC3GFA7IhU4qsK/dSLvanA0OdLWGWmsMjS60DFAmNt6kUxs/vmUmyBoWMyW15t
h6T91tblE0Gq/JaSSbvzg34yxYN0190m80Bq0vj4mhofsVa/pNNxnOUp1Yk5e3/1lHZ3IPhnbkJo
uaOqFDQvK+O0QnSiSIWOXKh498iGCGmB3gQSAtXwfaGcec5WsEIUQ1HIdwQlBNWeKij67XzVA5QD
nYxSQGzU4uvOb3bq2nikGfRp//6Ms02jnUoZakTQQn1gDEbCo3pJzXFDSlCbR3X25nmv+KpSE1FG
lcUbyVi9g0CANvIl9+N/gYFjy4381fe46csJmioobf4QkNDgjQ7F8pF22FFPThQUoW1Ar9rdsj5b
joHb9OFaQEWMJFLmrBWIXgYKwhrGdjfCo8V1F07du7YJJ7X1vQ/TpNNQt7GM2msudX7TBMGb4X10
4y16uIzl6iK9YPtFWfYI2E2lB4kuTO1MNQ1YS3V0JjuPiuWslYTOPPEeSLXD6M6YQTo8ScPLPeqN
0cgLX7pr51+xisLPNoUhOR/3/Yu5DnKJj0G6RyHiZi962EFMbf+xcO2enAJPl38wLMmONZVDyuOe
rsouUsUyV7TLsJEawOkiFhKJp9bwG1iGYbSUbtIK24I/YjFHEEqYByW9D5WtEbXGP55zkUEk5IXT
dAm81Dsc4vj7oDyudlndiCv5uNoeyIMz2EtuT9weaCHGfn9UF7Gw3ueoJMzhX/OjdWmDhyBalepA
D5m1Wgl7ABx+LNsfVomBF+v/popgHWfR9HxIRO1r8OaqfYWcyEQbqwBpem5B0igtz0YT7ftry2/c
d+fX/NU64My0zdI97JHibmkniH/H/wmU7Xj+JtoJq65jNo3y/ARuO4dDO3fhesSYTnjC8AFzXDBJ
PAWdyUXKgIIPZ3efGhBCBk+yVnQxbSvWdilBchcLQMfoIj9cJaj48O7bpMTzx/Wk+/0ToynlA+o7
kpWUIaAIUZmhFVK9pv/wX/3xkKtJlhSQLnHYsM/AYIniohCEwM2kgvrqPduGQ359wdZe9BdbZMQG
3oO+sUq9satRVx+q30X3YA6a3lDsZjx0AXZazRp1klCAbY7CKzwMLopV7LPfijXiTCA/F2/x4eyd
nPFGumYGXgP7wb2FZBt8byRFHH4FqjN0okP1hquiEyrR8iF/MIDf7dJ5XAtmEH+ZEKKSq9s6fksy
moT1QsNpNUszQHDenHaiuWMLstPT1mOt6s81gDdU4gWQ8HRDrBvfIsj/7QSqQPKCDlAjJNSYL23O
0zLdTTlGMDxsKp+u7wBhcgcq/XtTW81qnjg9ehhOJKtJuVmAlxTL4XbaDZuqiomYLKQARKoTO7WQ
rJzOO2ucwSjULOlzd+aHIuberrDySZTesL5Hb0YwtkdJ75arl7FeLyPhQp78GHGVJePtGrNSozBt
W+/cBuRp0502MlS+oZrdwS1gAnhGzum/k3KEyNoyzLoItJdSoDvynTd5idkPHFlQ6yEzYJOaAPjA
EfP56AZNU1YFtxZPUWTiwHPVdwRgqiJC0rPZ8hJ6JEWq4k7wEZ5H60ep/2iYljvsnnzuUldOivhz
hLcdgEZ5bbAM6TPVbcAnDugAW2BVnd6JJ8yu8iSdUyZ7zdjv1gcUl28aDe6d1j9S95GnwdDXuJZP
u9veHQ1ZWJCJsykcuh3fvHtI2mBqPed61Yx3KskiRU5ZSi2YH3m4w6LCLfSJKIQqK7TpLbsIEDG0
Lhrv7pyAHKGpmHUzp/zYqTAw/dQxbcYabUTlcQlY6jtgsChoLr3HsyJBXpnl7QWqtk9UGtK+2P3j
EVudjdH/GLun8ujQEdu1jyfjDv4Wjjm3Z+5lJWLLIxeQYkye3dF7PnBw5cL9R/kV//eZxLGdir35
OXiJe98NhHYwDcBh521tfq9e6zeeXXZRJ5XcVa4K+Hc8Kj92+IHBKb4eINSeFVkf4JgvU61Qwwd9
E5Cmb0g7gqqOQq2/H3CQwB5a3BJl9ROlo8S177uoxAdwoj/xl7J6HUAbsx9SpDxDVUWJTUnWR+Fx
W47+iEWqzwvElqudqMoi0tLxHUnM/Z0tqAogokeHic6+8cN3Hb4TKy5gsjJyn2vPbBOug6ehSFkc
LDCGMpxaY3XFUv1CDRQJvM0uqpvWAe9Ay+ObokJOvrLV5zrM+gJI/STIAQt37Hb0iLj/YTideNqp
WAz1w10LMKO0jy19K+IipayUZrmKfgvXWfNe9goI5jtzV2J6Wl6T6+D5Lv5v1ohvDjRUC+xSG3k4
bhQlxFMSL3+t3OoB7GFjKLzJpRaDATz1olu9O/Ir/GiFfXHur5U162rMegHQk294ciW2INQdpr8R
gurGuNemtSwh7PmcHmTQ3EHEB8UwxjmCjxC96qyKx6X/7cnPdO/hrcihylMO1+mrEgqpE9HuzYwS
+j6hNnKP+PLqHAkV2xIccP94geEm4HVU8VSSKBP4Gj2g6ulJhR78yCcydIgcHpblL8IEviH3H70u
9xIU4slNDlDhS8DRNE03TlWn7LC8NVip44B8RxRzrdMWX2tJJHHkBut1CEts1GrlCYijfhdFV7HR
tA1UepgPmNTxygA4UgNUF0xi4b5Su8DxlwPjQZHEDoMVk7Xw1mGkmYbjaBFgHt2lOQFHnNrlX1f+
pNfADiIis8aOXO8dBCee3yWiYuyq8+hLM394ysEqUXfZcfIyCw5gT/5XnhpSCqdMIJ+AcF/w3O6p
yonfd2fkjnFyjixSGoW8fthhQw7IO60gDnjLZmNHqh2JV8456HTfmCzhsDocBlkSdGqURk4SSAyZ
SQl9ImLrBf4zNaPTunWZeG+fXz4punxjIigQwXIfliKy/Zz3Meu8ITw4kmMJs7gGrd0M4CANYFxi
00pxsxoqCVhwPraCyB+g4ZM145B66AvqhXfmKacwFqiGTi9K+3zPVdrEGSztL1kzr8J1SG5fLfIR
pCZs/AtXH7qYPIQOL0BDbZWsFyrjAhvwLvDbvHeKGKKOgBxnxg6+tTB1iFACNJTI7cxbb4pAZ55r
Fgx4LsVYUFT5ESwM7Mdqp/lg+JUa7O48UTHEk1H4wHNMkUA7TLJYoYufhRjG0Zunc8j4ye82NAtO
m013Uy7vW43gEYoIc9qBQ/NeNzPkEa6N/Zn4iaqS1XEJ+X7dQiPU3reeWlAuscoaRBP6Svwaze6B
S5h+cFlOc8gmqlgaFp0mgk8PxwjCZIY4jny9OJg25GczxSd1SSzwGUXEoW0+Tp2cod9FaDGxrMYp
5E2bdWvyS7A7dPBKHCnSEFAoclx6J3t0D2PPR7PZOOS51QS/eTNu9YvuAPvyiFwMRH8U57I6Ovku
ItonK4W4KeypuE1Sywxkb6prkxNhmCEvPtmneVZogIEbywuES885LWWQsFw0RwwH8B42rATGlNEA
hWbxMheNUFXHmT+GuecP8SHIy8ZWtFlZkQugtASG2Tj7SCSg65JA7/T7Tp2A6dwF7YS5ARyouMiw
aZxQibltib+WyUOUcOBoNdE95Dq1S7JgJSBoAHCvO1n2QGF1eXBYGRFNlJeLhaY6oxV1HufauJOz
y+nLvkDGpLFN36C7yEiG5cqSlT08JmtebI4MjX1nmqHZbZgUcGGYjm8Jq5xD0GJ5qnaplnE5VoOw
aeSs4gvBCanOHqgJkV8AQsLupbcvI/6eD2C1NRhLTGtrjy9UdjU3CGGLolJhFXytzOyYUA0z78eg
xvnD1iZu1ZgPMFgDxhsOZrEQ08bpmotJKBvPLNL78ljR7HVLuhav5M5l2xaDSpMkgGsvt5uQoOKg
ORKDf2fUtWH9GvfJu/XZ7TGODoBv86Swx3wUmD0hRzjJhJsjm7TdUr82eonsKasPOk73gA9PZsrh
gTwCDLXDcCFDUqtq3JsTI2WdYhKtwhAcQpHSxDsSo0mUVWJWWdrDW6HUb8PW0Gr2bINNxn3d1WlL
DhLLeKEwVqBwBrsKQT4tNIwS5zi8CGd2Hb1i3R4ouJKFi2YG+6hjF1msCvT5Oaaov6YEqJ3KITqm
DycpI4kDT9JYlYLyro9Lw6G4TE9bE3D6ytxaBsA2lDPg6TaKc8GcXjCdp0Pe2ne+XjygwKMGJQve
kMOmNqVdmxp/4eNFapLzU3vNJcRsxZN0pphgC//hkjuN/sVuXTfyBzZ6EF+pEOjpkLkXG9lkpzTk
0LWTbVY+ssOvtEl1TlMlHBPRCIHLNdcgs7Cfe2lgjoIIcvy25v5N2g6+pmCjJJJsi046QpdvZXdQ
9hPE3MgO93mwoA51bGyHXV5LPhf1KFaYigMJVvoRbH6d5qmWuLKRY0KidpMkRRvMZEIrSZz0YoR8
ounO+bGiOGqYOHZ4phhj0XVLBKQSJkzBCPNrkQcak74QLPG3CsTTOEpZy3yffoRtNEwr7MwcGXgQ
VI6H7q7dm2VKaeW6BmmTEZ8waubSSlMqu9dZMyFiPVmVfrQcQGeX4yt7pb4a6PCR/0P8xTkiFTb1
fmrElZKcPSz6rBwihZHxVGss2zhPOwdaKb1VFqSJyHxpQXe5WWmErocxbUM8NMPtZQSFSHj2cvkk
cWM49gMyIuVYA8DL0dvUNJaVNCgt3s58j55HjLLj9x93JtpKESaHWHr/f9FHpSREIvfLywbv3Z3B
Kba3XTInttTEA/QzpH5WgDYeV55RHp9lb/UFp28NbQtciZKaMvZ/CjO5XtvlrGngI6nsF+oCUJyQ
HgybqV266/1Hvy2Ry2Fm+lGesVn1iaJ2rpNczg8ZzaMu1nzlotOhQplp7aHfBYShTvtqABJhbB6p
l/9gW2JbwaqVhgmtRZHqyTbRpB7W1Yc8fp4Q0ow/JqdYfcnurVq9mpXgQbRnQzFc84xHBXtG2wT/
lKwCHW0UdBvCfRiHJY9fqXdp3JaTNloXEw7XzQyfCaQhiCZ9OXhL5FdlfgaTIblLL+0h5PgWBhlA
l5MJOXQ5FxmLNtgIxMD/sjjame4qL9gwbrbYYDntEJVYJVAqLFO+eH9FxH2C1+CB1zmvf3eb8Cgg
ptgbgisTrT4eyYvfh2qzjUrV42AWZyN1jQ+XSdPvUmcXgoDnNSn8ciw6nTbHfCnFHl27/e9pHn2W
Pi353WyI+eYd4Y20hSDP8BPqgT/rCW6XiCErB5XNo9N9AIgAkUzvKktCuW9YdsE3B/JdZXoMLo0u
WbSbgbN7+flhiIDLjxT5eTProF0YfOXpR1aWm2I0AbJ0QJSgPqyp94F9owHz5EnmCs2nRfiV14Gi
4e6xveJY0GE7Pwfr5mKP3Dy2DRxhJYD3jDOsWgXb7vdZhXV8cg6RzAaM0jdHjA4BpVe4NDBxvvq2
6ZkNuMRNJ1fOE3H2BXnOX20v6Qdi+aDHCgEz2Ck6jUex/bpeEcdduKp1Zx8Xat9U5lcchcgRhrb/
1lX5Xl8Krwsy516Aocfj1EvTLJ3tAdwGysqxNEhXzZX1YeGvfjai5GmMTL++L7ZFSARpoU8qxDgj
gn2baUXXl+Q0pwtR5SX6q71Iw+beInd/+JM643k3/ATOnfcjzdJ76VCUTZFAX7S2q8tnI/Tn2CAJ
gKFTjRTO9bHHM68KRA6eS2EzB3hxXtX+jKQX36/btWZTwWCka4nVs12rcGcSEF+8VY5JDarIJtFm
n6YIvWXbZInheC2GFlO/Az9UvBeBB8zMYmfru4IkPV/NTw+pwAX+fXNlYhDkBrfp6o60C1DeGz1M
nkNcBQ0PUGpsay577xndtcK349VYX8cogkxI8xAmOC153CijQH4XjxvNEiBJi75C5ZXS6Y0hgQJp
IhsSKLdV0N3I6d0OOCuxVjicTf/Yu5C48uT372Ct8FqC2ksuI65taLv1IMAc8ifBj38WPJ4Zk9Gi
ZCoACn26MiEfit20jHN17ImCvDWl41fUUpYUPaFIEwjuqiqXYwZkFVT4oX4SkUzxmcR6O9lW+FLT
IFG3Nz9xHUcrspKH/V4K0SXFpAE3ujVAzSScOTg5jgZQky4vzwnxV8xwqvq3KbUBttEaHsGyHuEo
6kkJNblFrPFhx4Di8jGHkUnaWPR8Xto2Ynco+OpfbHxD1nv5rsNCPQHZhBpa8bWZIT4N+3ZOzGC+
fwsgw5pC0+WOe/XTlJKtaMRggpXCus5dqrltz72p5smEwciiSo+zvWaqCNYnQa8C9zwrwGIufNSJ
0vYKPQFj+0ibdebccD7U3kqJCBMYVa3rNf0TWvmR35WxvRPkWwu2U1kDVtdXjnmjezri/6deKQUj
WURGh4f9mNCB0F9YQTidu/aEGrRtW0aERq80Yuw9bq5tDpdaOeuZPUCXHso/owzAOiAurrmJSbn7
FYiNweow3+ff07ya983/C56jqvX70huSEI0KPpfZxUBHQ1VSF5DVc4ii5mCl98HzpeYHIPkHqijw
9s06DsXVcyPb7nGtYuKJeb0HSQoVUVy5e1x7A1SL36EKGd3FxiXaBm8B6hYeunOr3j38GPlduAol
SMhKpRlasJK7KIq251hHkKeXx8C5ntG7jbnfWtDNvDjRBkDTEo5H/CMgBGj+DnUiIATLIrzzGHLi
Z4R+VeCAz0EqbygyLR9GmQU6UZdkn2K4X3SOfaejoPe6p/jiO/23Mc1UPmltObhNrG6icHgdFVyn
KexJjRauRFTRc0Gx5qwdlHKPFAuFvsauLqy0SWeOQcdOCmgeo81n59e7crp644JbdL6KhHuIYsk/
UfXiUBOaLnikEoGoB5hSJIFj20LGZ3ta4dJesx1bnTbk5PkbTbv0pjGARs4jll2YYDPg0+TI4knH
P/erhXXIB1LYURgpTqo3n64Ug875SI6x3pwqh/h7vXgqN6EL+vRHlrw8a4SJTEbYByGyfqphxWvZ
YyFPBagDGEbbtMWJtZC/+8Tv14Vkr2zVsg9uN92mf72pjyZDjqLAzI2inebdGn24Wd/TsbvHeD+z
TJ/Szu2kjqfJ2sqD2QdOaIToq2AwyZJl24K6nGKYE9G2Pc9/NcG8sbcRL0tcbbbvOqSFkWi9xgwi
7yHg3bsj7HB7dJyHJrYLAYPR6UDPmGjeU9DCOyvEl8qd/XF2y0ElMaJ39U9cmYgCgz2nfb1/MHF4
zUybcFeiWXFtFFR8xFbK45LZBt41OwmE56mCQdHweQbUyTy0DV1AtAS6x95cDcDjU+ISuJpKz78J
7jcCLOAER4B9LrVTu9IObzt4YfnETFjrXTmaAGDnwYMs3J7Prs+TDCUg3jgU9MjzuqGhpDQMlXuh
YwLbRAtZucPMynnfFSTlfRMrDzg82+xx6YPDWOK1cB/GQUpmHMWkehm9Q03fqo1eSc3xJhDWkPGk
vRVuAXu9RBUyD/ZoTnx9BmGACnNedLFfYrke3urbwB9qqNb5w+BEO7CzaQ7zWfzQVjR9eHp9ZXYm
MB5edJj9e5+4xKn08OwppJ8mGckY0v0H72LK7jGmaDIl0oFgY1oB+Q8gL9x+modmzT1ADrRtiILg
Dr3sYHfIq7ZiWDELo0dmY9sHuiSBGE3pGJoSf2X8ed1Nw8uTd3Kv4D0/c+NDCHEIRnX8uVxoWEsA
mq9hZC1VMoT1xhJ7KT/ngpEX+9gj/UfI818cwzDn1OU3+10K1sx+RgjYpkfUUcqLBkpG4VI9TCHs
4J6LT6VGXTuJ4Egoktjk0YH/6peEHXIaLiPd/ycx6OsvCrWRZ3n8efhkmNH8gBFhS6I48zs+IfHi
+jOpL0PBtzYtr8yrat16fdVfkDRl3A54sT0fPsgMxHPKoTAq2ZaNoMlyBUGvS6Mkn2OmarYoeJEa
RB2lm1xX8PVggAKQA+Jpn+6XN0gWZAatI+ncN8o47J4F0R4jveDGmGMf+WsuYYWVD3UwjjaTbKR/
5Rj1zuOQBzIVSBUcTm6QaBHeQFMZMBcP4WqPasEpQNSmf2LE4Is/0pNV+TcKEmtWb8xMAT52eMjT
6uo8y/6zn4FSa4W/LssBnKQqFuHbqkjdN0ji4VHv+I9N7+/TuR+sdfuoL1TLZYqNcaqGCBKUNT50
RBELN398CmcYNz6/zzLBA5xAvXwaT48DTyhb41Iv0Tm8uNFw+bxW8ShBMXqcYmzS3HBSa4ALHjNY
0VjY58dLVJszbwnaTxiQh8zEQUh49MuNk/b2AX7J/z2hHaLq3QT7X2hIT79w+FxR1UDR3+x6P6Rz
xmo/NteFONEI2HJ2tylA6vPiwLQmxrCrp6y2RHh+93j9or/t1lTsJ4pLucL71bsU/v9CJa1gdWn3
z1Kz/gFMrX57IWFvNOYqbeWi46GNnhNzk+3udPT7LGi+W3QjqMat5vVmlZVh3RuIvaWyvIDqxc2o
lCj8mgAfo/32bCaPMA8CwNk2eSWl/JIeTfHOaf0MZh+h2am+jXcdYh3Yh4N3hSEbQi5oiS5L00oN
G2lAhTaxmi0E1pvAfIB1p012ShmPjHoWUbfX8IRkWK9bKiDdUZ6uoHQxw+dLo/DG/Axwh3/d1YMp
F4D244Hmm7vkwShUq03IB9h0FNCKqclmOmjwDxeiR8SKL8f0Dl4XT5Sz14K+6pq/MFnllTsVRtx0
oAWYDRPxPdmqry0wvIy9q9Pcmho+ES9L1Wd1MTfAHwzJcTJ1Rp6/U4rTTRstbGZNMpuVVY/68f8F
ZRXw8pkKq/2vwPDYF8qLNcLWQW+pvTrwnahM77PwSg2RbUzH0kVNtO0WjDcgXCvQ7Q3JAVAfEv1o
cnCjZlKVqbF5RoKlwMrAjb5Yyfl9DX9AYNDAyBch9zHlNfzjVTvmam5OKC2AulBSeFndvK1Lm/0l
nLvfWII4sp848pfJiyA3oSNN909XKH3I2MyvRp944pA2lVqAuCzuwbgB1WixlPsPxSRrC+igNMSw
HP2ak7GmkfNxtq96sVyFy8btM6sE2NIyrwhIZv2JlG1ApVM5C5y9ENVPZIG5WsML/je+d+z6+EJS
lllieVt3sqrbq7Agi3KTzGjJTx7nid2vQAHSU0dMG2OKvXrVIQc9L9lkC8FXEHuYwh4ROn2Jje6+
J6/8eY7R1KjcAFGhgQiI7OMbXsONAdXzCVxbbi14/b2GJZQJlM5l+u52ENZ372+qrhV0XT1DfS8u
MQdEjD9JYMHuqraxe6ETa4Jf+zwvXo6VHeqp3mOU+iHLGw7RyRfy0Al7p7G5R+jAsO61s/D/fNF0
8bXE+RX+4847n5tQLooQ67yWhvo20HS8A4hX/WDnwuwmt3PEiSTx9SY67j/hQxJssb3HQv6mS6aa
k5s/UA+csZt1MTZjKEBVHjJO/mbu+Z+vV14hfqRJdQvRdfDXHqtE4gqRIqtlC0PCtIHcf49drnvA
wb3kXa4oW3V+tJIs4z8l1IhAEi9XYjd9sx/Si1zaDzoGE7YolsTjDlTLFaky43BDYRRix4jrivg1
i4e5jn/UZaglVvA6kzjrBVwCgcOk3d6ggLfBRsGLysl6T/zCGaY8GsbWZHOGKvh87nwg5NM+2ej5
qiztjbxQQGqgk5KnYEmVIZf9jasLLKn6prGpNomDutjr+UBcVPra7b4V+pUIWEYOIXX0UxFjPuJX
zR0A14AzuyI9LtLTi5+PXFeLGx2Pn7EvyOoC5tL1rfuPDbmrJ+TilVpGXrvacZ/7tMhToJlzJ/5V
XIn19k3gc05x6cNkZ8T9klbOpFksTH41lkxSLRQQ2uaMURoGdwlCddz0jQ/isigMPuJGM1++FEIh
8NtOWUQ7i2EPIhBeTl563KLg2R+K8CU6L+ZIenqHukQ67mo7qeliNJ0FYpj09i9ulcedFnVcyZUt
bpraiB8yenAVeJbAowQpqLYlSu0BaK0/3PDAhvJVfsJ9nFnsHh0UvpfAk5eAa7zozPI2DgAPqiVs
DydkMjr5Z5nrigQ25Fl8yf77zxf52u2BTnluJCMqiUWcRx/HrxmWzudy6hzcRio/9abCCwDd4FWR
2JD5+FRU2eVnKIlyYwmwW3a0qCOX/ABJLxjyjRbo/Qaqecg8kL90WKIPuRnjgcvEvfItNzI925/Z
kgPDOu6kiZMpY0NoXT200BBKqj83uOPw/vzB0j8TCzhLiOH9mzDi/KatOqg3TcBcch9dKapLb4qC
qt5wdI3Us8ugQrGZOJZOIt2+EB2wePPH5Cm3T6phhxwnFW4z75lAP23ie85AbqulD1UwFFsphsm8
DHcjLWZOL0D+WzfWwguQvt0eYfQQA9kDS252E8iGnYlvIpEYz5+Wf0buOKuHzB7aL8QlNa9kIIHA
eQlVZkCU0dNv5WhN/ZDTFpzktw/7Whxn+flPB25ViFwVDLgBL+hpZBQPUjjiu0roM9axhjjiiftQ
NCMWpeDlUN8fXRgqswfgIjFfevQ77ySgfE717mBL+u9WYR0toq1HE+lxKWSg6cvwrz5UmMgMBKPV
/rwp3AtG4mbsEeP1VBTl6/IJsrGZv/ncHbIWIZSxKv/lbk/IUe7b+k0C51CV7/QjqslZbJx7Ko2E
/EAt+QUDQpi3hyI8qoDOwxpFniZ3XtQX+r4XT1VpwnS1pF1ScIerKQQASN1+PODf9HiukFk2V4ND
jNAYRDGgEBuW6sVwsT/R4c3z+C26Bdv1h1+cZ73TWvi25XJUUERINUEl1dl0l/fTo8M4q40kIomB
J1a8qAsQzBlitcGBXz/fDqWL1eWzyOG48gpUohmLaFShd506WNWHglwZ4UMbfrOU2krSC5+nVjSG
WwAwWtUJ7IpueqN6rc/maPQcF3wCJuvhq9AiIuA805BEYacf05sDamzDfv6wDc4AUFcZPmyBPhdK
8Jh9f37B6wObhHAuHYE6KZKH9A0nlvIP/OHM2IO7IDL/Brzf2B6DsQzAPY53IGveF76Lbd+7JCQS
NQWHizjUHdh7jPAyS9H3jSHOmT+AALSwI9RPxxD7W6l3/peOJ8kL3tMMONBSfhtdqgSd1SyEe/dc
1xXW1Xvp1H9bShU5/ReeHY2I/K1BDECv+lbFfG3/ZQ98bG4H0IJySXzKpsStR2E0vIjGO9vLo3pR
hpJ6IgnmjP8SO1781QlZ0TX2F85uchErCcJR0rzWXoW6znQ/lVPHhx2qnCU6GAdkpf5JQVLMD+wF
z/jbRC0E2ah1oOcGh5kQKHI+X99IWKhc3MFlvx0htElv8D2aDyQvF/2VayWxsIXkCHCN6duadjkI
bRvmNpLxP8EcpeITyQl3BKm8g+HzxUuYnJ29990jArJXormaS7yTje7a2jZEG9X7uOGBGdFMV5WN
ZGNJggtKwpImZPWEF34mbDNRY0C7ooJu2Zy5K8XmtN9JM4aSYsiIxE6hCtgWLcEnKsNMrGJ0Ij7x
F/iX9rAtvv/iJZe+rVqQengGNjacjjDH5A0spZjfyXL0ja57DhfBiqsTtG6lPEDCJsnyPPRjczQU
jXryL0GRPmQxX89tOcZNmGN7zjR3QxQdN8HOqwjt3y64XHvL19KGKElWaswl15f1mi5DQM+d4Xr0
Q4KUnUl+ShAg863BHwNVkQJOd8XNzQlkrkXFlK4ClnCikqlYILDfNQyvF38NeSnNAD4uU7nteTaP
+uCD6VRubgXvEiO2bwOfuaQQf9lH9sEg/XEDRikWPbMXJfnTaBgQvx27iZjK4mXdqDS5kdNyTaUT
tEKBUx3m5dKEn4YSsh4rVBlVtFOfDg/sAYsMfAIcznJYk0O1vnONnKkp5LE0Vm8iibTrlo8nbvHW
bpU2KTVlKv0SrUNcX162OZaE75ABPGVtuSf3ZMB3g0u/oGlI+akZTDTYG/7HZjbp2MilY8WZ1Nz5
mJ7v8tHlIk14ID78+1Z6moyjUlvaUjxEgj7+CNfCht6YO1sORxtM6JZ+P+M9kbZkzvZWgXyTG6Gu
wcKgj2otV5wHDtWcPQl/86ECGEquLiY92LA1GCwhvPeuKtOBfwU8mQH9tp3dS0GSOnVP0ZQxWK1m
Viv+7K8CPWfehwFowHyhIGHcqoFVMGxmbWsG3HypN5T23QakFU9LktOK9gRvNfBq/d+QgZzCa66m
NrdkF3kltNpvMTZheL7mtVQuWvD2vmema3GJLA9EIhkB6BBZ7NkG46HioOpyXI+EXsdML5Obi1W4
7/gX5LEGGVlKYKMSa6HMVFnZLp+s2ocd5K5wvlKP7uecSJibEKBdjZ+wuqGT4FVYEbnajEUDxiKJ
u614kfh3Tc9kYRA+Om79XP+pJoS0FBSQfw2IY4JfL1f2YfUFQuOdL2lMeXbuojnskpupZG4sVetE
P4YnJmK5669KwxNk605zwrD1Q6zbOSQSO1TkwcV7+6Da6J6wANGaZChYf0RYCRyH7Cp/1ZtMzoFE
kk0cdNa4UiH5c1I+ud/DkNjqgmsFD5XZiltvc3gqvX88bXLJ56C6L6FUdcFPVnlw36Bp5uhs5Org
gKEw3GwPE7cVGeK2r2IqvHYhrPkkbbDtDj8gxuqtw5bjdeJy7D2P4F6h3eM4/Uh/Ln0pLzvTZQAE
B5+2PcGPl2tSR70J1Di0d7Vn3LVWdR/BFt2cSY9O+cNnz64vbrwQn9PJi3TDRzrZlZyGlautsuJE
9DatKr7T2KgRw+pGpvU+EAp0R+Opm5QofNFhxw0EjfXODgx82rkcE1wiGEMzU5f5WzPgfD70rCDS
r/4Igcqr1XaKKSBcGA6gKpbneVc+0cPNQ+QGNHGV/pN58Gf5b5vmFD2/GlXNUQxn2YtrKpwMSeGi
t24RbvLA/5LrHvPmFwm8vPEf/BpHkmwwM8UoDze65oLk5jxTS4rPSc2/M4UAfemu6a8CmA0Sh48V
wWj7ohs5C9ycZWmBFVlhI907CsToeOXa6x9lP76t5UheBe5MbxBHXw5zHf8OopSq29hvxCeuUuM4
GBxRltfM5BCzl8OLDuiaEoMojPYqoAPI6n2kMsyUJ+CtAtNE4/lQ5DdQZdh5luhUB3BVd+Enquw1
klOvFQ8qYSS2UBRINxMNIpSV4ckX93lxYfcjXdYXaYOTt5J360tg+wgLqx5NZHAT3WQ8tANJPsAH
abrxOZzI11uMQRd+WxxmBd3495amUbWFrxWHcf+Wy5PxRI/mVJrGlyF2g+Z/Lb9Jy7F11pmujIRz
21lYPW8atkmaE2hYv5lftsiz8pb8iPEuAvGfDoP7MZG+c6m7vQrK+kmRFGx0QnaG51MZfey04ZOZ
QyNv/yWfPJchwhxrTaKADlunTRRTw1PYVdhePmByG6J/Mcc1j2lYXwfRnih1S5jCxJTTcreHl62i
wfyQe3LiQDddLwbknW38MSZVdQL7hBgw3efuWyorNqkM/oZ1h7cMwGD+YB95M+YDPJ+ESr6rB916
qsrfGN1BV9TtZCZmwyqUcqBqEsBuA/gs+PmtBGmM+tcyT1hCo46yYc2yilP1N/e/j7OU8Q6TVjRH
zl+kTf7o1AdGu7jIweJci42TaDGDnmbqOMZgg8GlEJMxrOhWVb69XFZNXpmkXizDly94ShwKN/E8
43pTkJprMCxjqDI75A3ZOf2p/v1DB1gS4F4o0RKMgrznc90q7vq3skEiYcf0eVkQvCCO382f4RBt
Eg38gFGAbHFxLVC1Y0j3dSORLWgAKv6w+3iaoqMIG5lhDvCT8P1WKi7wHJ+gioPTGyFYmUZ61Kaf
JY6UOskoILthhCyq5wkyo2SWHKP6a1rRxfvdV7YCu9sKWVLqu+onJQZYaAb6vs8G2/gAws0kKLHe
cmBVlUyvNHeSOwmMqq4JDY1BVpRIF9Yrx/63VOL+sU9/bHvyno0yYm2LfeW8O8OwbfvHPgA/+mTF
9pVWSiHaGyD6igVwsWUcjhP7ngL3C2ZjIo76xs9tGbEDMLyie4EiRLrtLqQKGvG/7GZEVxUfJKty
YAQmsaNE3cDuMqU6di4UVPLw4GscOBb2ir4hJOHIKeuk3vd2MES2jqnUJPDRDPiv21wDYlvqtSlG
B9g3iIBvhyDsj5pXKR5eykXP8x4Izo9WZGPf/z258YZkdMS55pmjr+3nzTqAkQA3od0dLBd0637d
W6VDOxKlgkUAmftsy3EAjiAct/jb32SCTlbSHuScMifat44atDutDPzeYowOFg2w87iSNScbAIFn
LE9Z0ICVDDlD9CaDg/48NQK8hGzLb8zxGXVFDoujB9ThWUOhXCr0a5bCm6uJuohSIfQekanMRo0E
Bxun+gWe8jQ3XqnUc7/6Q2+cCZ5PD0ekjiRayOd1Yukyw4eVBI9tFIEGHgDffKv0KEGb7XsX1eF+
UyYfZqJUaP+MHUzMVoT5s6n7dFW4SVf1/xpKZHKFOsMccozkm6JmCAslLsGJAj0Fpdq3L5BUlhOb
DNywtfCVeFsmeA1GHSYwyuxCSfmwAtFmI5qz7PWqP9SPiA1W7K7LgUznW0C2S0kvJZZi0wqGW/nw
HMoVvcFVOuZ67CyHdvNRsOCLCW+D7SIW8NNxJk/ZLuZYg/S0xV17IP/0gaFIyvXBIePsKGxjPDEz
08YrKijy0lb2g784qRgE6TJUorETOcUx5igj4F1oaKzhxHuBSGgY3ZABzYNZSR1kP1+h4O5bKWQW
OPpndMgvxexbUlOwOfwc0o2qeNgiMy2lMMvY20sB45R3c7tAWRhf/VXJ5wE79RwV7QpzeFSkCbf1
sQ4mnYlk3Njy5hq9pkEievrVU9UDZsLs3z8GuncAD8wvt8H29J6qVJVyh8TU6BPt5T/zYwjkvuXP
Bv6+6U2nK1nAJIQT3znzhn/jciFr18gDZJiZRwFKvFGnYGvyK7oyIQm1QgpoaxOKYQPMs0happlP
w/8PZa/2lZBTvavGrnTOPvhBKToL1GeaBzYrnoS5sgfprn2kBgtzXz+jLbKlFMityt4LV5kCQzHE
q8qaacQexUkqHZ88gbxkTzz0yabe8txlbz9F3dgwrbBdAKToyaV89xn33xnteQXyWhHL0WE6FtE3
vM8LSG/LBQrWYPdO3FPiERY4PT+anR5TJu3JOZ1za851R1tYH8gVzS1W8T0P3kCNKTh+/CSqlXXH
3Zmr8tU+uDC1rshs5KNmysJDv4RfToPbx42A0M3JfPHAymi7/4lS2m8+eleOx68TVrv4fvadpU0k
6y5PzggOrZI5PY+g/fKur09JV7U2X4tAL2oyczhe8ItLw8eZHMHg3r/u6ASrtGRON4I4tLHgcHFj
R/9CcdDrqvTyVwr2Y5XRVUZ7gY39nhZJEQedc5zpkv60S6IMtNbEna20OTC1WgLNgjFkm6cBzIF5
hoX6SFPx35YRIdd6HmsOqPh3BYp4pzD2Oi5AHd5ZnDaf/1IleBbKHLFgiFO9yFDRMbp881kv9MaR
mYqzAtPHVLgr56/9shJUFv8gi0OI59WP774UHgxolc8H9KbiWZ81UOfxSQ2Z+KqIhFaR9wnKVTvu
HJtNqO2quflCWldBOHctqLeq/yOtP3UOPgpH2GHEo8MKxf4wx6gyZYxxs3XOt6UuIFMat7pcsKN3
oTlwaLFbess9w3Bp5kaNED3aYDPe/Ba+kPshzKYq7JZ9W2SAisubU0qV9G0IXCIyLA2nuXGj7/LE
/7il//VAIm0bxYQUivuh8M4wCUdbq0rMakjHOTewoF5fpK9gKtEeWXEOTq0NrydrwrFAskG/QA5M
GhCMU3i8n4+cuHNMMy34shRcQ6CTaHgvwZwwCPehuymnFwBmQqQ5bbsNbnOEWvcS1w6sSSBsRwlX
xgUQ2uGu1w71xkz0tLRsYK6KXP8qXi0BLmCIegPRK9NGzaLdNO2eaevZm/KHB+E06yrp6fT3mqJv
RIrNxMGJXQ9OVXsH4K/UY2kxaLOBIC2hxxWgKhCNgY7N6JPIbDGRngMt8qnLk4fIOd4E77H8ZQkO
c3yB95OrZzc8AJ3XEReLv+CmFIzfDBrmVo8HitwxS7XSXJlQ+Hn9xwg5RUSI47PJNVST/FvO6ep9
mMdB32vSt/IgTqgmwKRloNs0g/yu3E+7j9FESOHXRkarrOuiXSjV46ZW+htfvHnZPVOFqdeX1tKW
mpufdEIFg8oH6GfoOdkkanFm9Z2y+LtRE9bMq2jecDa/jGl3oy435mxM892eae0sExtesn0Pz35o
J/O/LHKzuSApn22lNqHClBm9vwRuxLTWoBRUVDpD4kEOGFcPpPGLwGiTScxYAAzv7nfXjsgcxW+P
MWv5jD+GYqtefsRlY2/MWpF6/C6NEhcKVHOhN+UArPCs2ldWUfXeEQlSiwWpv7HSchYaZO8RhS17
IWKgviV3HfxrxxRfV9zvECnyXjRuUTX6kxIYDDRAxakrMc/l3Wnew5beXme15P4l9oQBrc0JQ0Zv
BduA9e2fOuIS4X6Yze076Oyv8z4jjzSehWB8UlmdY9qw4x/nQTP19Boo9fPhphT28UjPnGERSqu1
fmqE/2FC2WKTjy2YwjJ+i3dbmoqrUcpsdS9te1oen77qdz3Z6sbIWBX/JHbf1fNPWOsKHkg7T56k
sZS0l/GnYinBjt+/GSxOSUBgemPqze/bJU4/FeU2+4aGfPeFNqPWEdCDVeJKAzjqHLN+9vzaJ9BN
0+m9n6NDRIH3rT3/BS6WzfFw8PfXSGlsHlVnXbb9ia5mfb/71TnT6OmRgQWxtpWw2KpQyC9FYtYs
55mGC+aPoG4/1g9MfLOCA6UYU4tBuK5gGCPoZfbKP3xn+ZBoc0dlViLTlzSTqaVW7s5kjps/Mraq
idZeFFfD7IqnihixGqRMc0ktiv7x/fDYsueuUfOK+aAccO0VqdxJ7iCABb/8cfSGogWW7oWX9upG
Om5S4W2G9UgnPS+sCL1vzYdWS7G9oLfUhLT8Hm+FUJhy+gSfyyO05lGGLsVnEMUAk8KCgukd9b2J
8poK8+e9/jkXjZSNVR2sb35NEUTPlcr+lQvgVI88vOKgqpAoXZyrdUfMsisV8k7g7ndL8V6lQFm0
TppVC9NhwTL+7PQEiWR40gPh0o51eeMsuyZMvcjRLEktqpuLWaO7cABGzkfWMRHVpMCETmrDYp9x
VwjZUgqalYxC7748ntugkL0sXzP0TIRWZJ6M/j9Ntb6TVXQsN3qwtC8PA3sEvQDxuZfnIH61Yoko
WlGGhj2ji+ltrrUO5y6riGqn7jSJPO+3j8PMtYP+mWGqfTfNx8xrLNGGkWT8A16x3LTSdZfDT754
My+YG7EM0HexCSMb4zNViOkg/2ZJjGQMMImntf+UlNI5+AT7sIhW7O8HEyf1ket+ziHmWvnptja5
6kBPjgDxzT7G4gWM84m+8abM/+tU/8oCTV7q7eckVH9Cj3ox1k87am3zkEkZdc/R16XzmpN0uTOC
tjUDIWqRDxQpLrA4rElBukana9wZlStgOgeTSo1ifQ2LGixGQekKYoPQ7XC7W/9/AG8iESI01rs9
Zodf6vEaBvqSlvx03jNcwDjk+HA/wbO6T72oxtz3bWme8f3nvhHKdjT+/chKukWpXRxmre7WNAKr
w+phg/V/Ah/FuveWmQeeGAOIzajinSTapD+gomzabwoS0/RonV0h4uzRajUGIGPYU1Iq5z+UI5VD
VgsJNMsVK+/sUUPaZLHM03baz/M9TSqwbdtCNsFxv6tTcSXY631CMSJYQgJv36HCFe8chLoUM7J9
98U+NNzVCsYUN5tRg+4FvSRZbvQd2SY+z080NNJ4QOzAfEUgdBNP8HXmJnEBzKCI3Clv31SJYSbQ
lA+bRI+qayAmSinG0PKD09wdjNX750oX17w3Vs5mZkd0lAz4R83hTkCT8CEQwzszPsF0PvpYc5+F
tjxOmhtkVBr+bE6tts7TzSrGpOxgFUEzSXi5Y+u1pWyZeOmJQAYjaiipZe3gPtvAJz8/ofX8vOmQ
rQiH/+OGVaY5a1qmHjVCZ7r31SmR6r9vP3dypFbwN27Axc+JQSrrK0EG2I56Vwpkea8oSCUFOurK
OWrqIrRBODXFlLvryrvK8WQFLEHyJ4Z4VtVYVJGvegeuKv6L1umZVPaZf4jNNkIkbqQi3P7vwTlf
KzDV+6kNT9BiyoGPrA5DbG0qszNRyhSWbqiKweEMz2FLcjaLdT7zRKyoBwM7D/MKt3DtI6VsoikZ
DZvPIoHgGYygOhm0Z9XN9nOeNr81NrzOOtWsLV/bl1k+5DYsi3+fqd8uCN3yRbuGrJKuVk0U6xBq
aFMbxBlA4AAUbtd4ce2v1tN0E7RO0RkJx0O8KIrPCLNa9gMVy1CWDABxRlfpinQWOLNcBER0X9fp
+nPrNtBp7k5b5dWgmqDQpJh+UF+rDJUedytFwQHPQgMLZM3uMJX6svl76OIrCCDNs5T1zziZKIj5
0AsyZBM7UV2UJH/gwSqatCsfXmG6IbVnvVT5JF+cdh2+TiD4ZSgIYx8AUck5vFaZDb5Y2GonA1OJ
6otSQ6ydWcsFRaDWMNpUlKZEBCyS9VQ6vM0Vr/KphzAIvQLbKfCJdpygiqksj7AmQpkM5QxPtCTh
eo0mmYLnTKKZ9MHDdbME/yznfcRjmjT0YZQxZ5zAy3jnM60+oL3gTkVtxNPu6SfYAOdy+tnclpy5
4i7IAzgtyqvyiyFIXHEN3AGdU+mzW33UmXP69wsvQqgywX+hiKUDNdU4A7dDspGRRuTcK0MFumCz
MYKmpHxiDcuar0OsBuHs3CT+P0PpzFwi2tka0RGtL8PXXV+FPyWKoVoeS8CCwDavbbQHNgK2AoN0
vijB8KeidmqtlKgBeZ5dw7X6bG5RVcFaymUDWKZOCMKgaTex/gB1P19hI3TVCBepn1KSsYfISPr+
c+Tk71sCIX/8tDhboznG2OWW0s+6+BepKch7MCa9/4zqt18znwLT7K82Di29qy4RRj4F1fam7KEp
J1nDI+IhZ8Gayyf8FVyD/NwCXY2wsFJjcpcndypF7JeVFG0H/OfJ14h3ydY2p7bCvvdsAT+4chpS
Mm1Igk/kD4ttl/vC5KEkG8JiSSjCWDCPm4vXTUmkmB4pmipg4QMVwe3L7ywrNHchrmd2IWUQ4WWf
UbL6yLgKwKmoBOGuPcFvMKeGi/fOIV0tmvGyFz+ZZL8ukgE8+C2+fZOG5kXHOehAI6ywPKqWDj3T
VISrcQ073ZsTfbVn7xsFmsp0I8IXMSnonVRjRCaQ6Z+0YWHn77Dnw4BqMs6FweyYwBbc4BqzK6fO
gzmp7sNISHdqxSDHi80A9MoZiCKtUsHS3njlYLZpAlZr4+OHHxaQ15mtHMa90li/EursRle+x2ut
i/N+pzCJK54mKygyputOsR7IKs5/ntPP/62mM3cONgMuZ4fvoVo8LNI2X9W/R+c/NgShd4sCcTay
VaOCwGRvcRMGM1rIJM65QhG/YNX9VlNtnV5d1xyfi2USJvHrgr6tCD/Itfb7ZXgZOqVZNwiwckVJ
rVtCo6oOac+G3DlIYndYbzNOVH/pGfFIxcmEhlem3Xfz21yRkvtJKLy5D2c17LkCtwpmehMS2qMG
dLTT9CiDRWR63uhJojwD7nqmEPT3yzshoQmMMe9yZRk/MG/d64UXMgC6EbYpr6NRoskKZT5dAEbZ
C9WhfI/TMOZARmuN/bkLNL5oAyHqM06Op2fTQbA+DimCDYXQeQ+ZG9evGgztt3WwkLJ+suGvrswq
HAtRtTani3WOgXYRKTwigsTUg3mbvXWe/BjeT+o+4P0zCqrQ4J3kCPe+tfjYSUtI/HexDI3qZNW/
KwEarDhv9qabD4NdH59jkkpIF6e4J1pvos21zFXzOxhHVBQ+lwjlmJrolITEdzue5MD8lx687C7I
BP54NCJ/AWpcGYZqFbTLjZDuFNJVUpgu5tyP4ZwULoGYbkbg4f5ECBWob3yKYwYTzFUgeQIu3la/
tGuCAOMu9pnA8cJUC58ZJNoXqizsVGgUD1/cHTLtZ+Bpkx07D+1xcz6dtyZOsHeT0Gl1U4UypxEU
tRkUQ8WWJdXT+nDB4F1d8bcbQqL9FZ4CE4KO4L+a/oQHKSRmGPYjxJW4omYpqVVqSAdpQMY2NHqu
1L1Gd8pB1K7nuOTAY+WmbYIy/o5u0aEn0sNETwjqE4PI+0yV0idH3Oc8v4tpJJWcrRQn/zisciwO
TPMG/bOvSMQRy3qWXJHHTrqyE3Fk/XOXM/thGo/0hwa42rxHcN9T6v105CFJOyH4ihk5B+6cFh0d
wLt/pRH4XdFM/OFNIvCoZA2gEkIQMNBu6nCS/jJZNbNeDdheLBd3Gh2brTnyvFXZ1WY7CthBWkxN
VAPXxcKj/XnLYZ306DCqCgyiBsYGvMyWupBr2Xiht6RPFZhdB/jiZVii9M9weI4hg2ctnyEwEiAD
rWTm4ESmwr9CgS9QeZFegNM2eTTaUdNVyxPCVGABN4A1W1McJ/ia38gzk3S9CbCESS2oGYKMvgJE
UDc326C+6NorrYBtip5XJokTApRAQoaC/M6174nBEk0gFZh3y1I1a0jfeIfMe6zoqUeSwGw0O5a8
ijR0oNns7krY3SQdk0GQ11rT/lDLLhRGNAay4iJlre/c/o91QTdMYCxubHLNwgO+zIjS2pObv6GF
h+bkVx04cg9GIEdt8ZssIwYFOqwhlJPNH9fXd5WM3vqCGey9r7yb9dqko2fE874dZ+eIPFJMTqpF
H6i4Nl8xrNvzvFvp6gICUhi7sUZ3VvUcM47HiyMIXvoR/bbn0flDgkuIVdLBG6+pGEh6KGnvP3Yo
e47Tm4iY5FztL/W5LJVsdfZfAg3ktJ5eBlsFExTZOEGo/gDiPpbxxey+UmoXt+hOf5kZk98jyfBv
FeNsLLG7hX/uTrVSK6Vuwbh6G2/Qt3fKhI2gLQ9d+qxrJs0GKZdv/on0kqRYli2PlUeYdWyhQ1EV
M/Fdou/r5tGZS/avZUR0wgpMqmpdvJ0bvW3p1pchwnsDKp63Y43gYDEvpMeCMqf+Dlrv+jHsc/F6
Qx+GnhlvHGi8ZfZqZOyrCq2h8/SS70ao08IVH7am/ulyU2np2ZkEPUf0L+AJL5K9TNBrIrenMv33
W5yhAB+GwoQZ9J0dyJ5zMOgrj5G45BYddudupBlLqoV3NORMNiNiMrSIgv9fCTIvsnuXqjl/anFC
NUrf+SyDCJRod1KVdQu2r777/jFlEEDw9g1yRwrRhUXXHgZwJf5bSwLBdiIqJgFeYby5khoyT9oT
CPTZCAnN2vERCGUfWP3IRC861yYnNyxSUg5z/QQlT0ogawiUmeX0TL48ei7mCFusjyCoX343tmPi
wGYFMh4e63kMIdXVO2cMxPqUza5tA7u56SknRSSJ2E4o/Akg+p45L7IpaH8tePv0EHrVQId9Bvha
QL+3IP88TOJyAFh+8axP445F9R9u7ua1pISaXFZepCWP2ezj4mctUM488vICi5mh7xumDVORn2PJ
w+l0ELCVBfk708KeaXEQNrFCggbEVUPomOhETYgKMjshbuBxwAliRwVS2CpFMWjXQmdN+8YjhaNX
lrTCXTyNafPZz1wab+S1CqxBJlnjrvD4ip0iAZNjSr8rIjzpG5Aapt7C1zIRbFBNqhWTnJKwD8i6
OZ5RX+C6COAYe/xvNCq4KC9VsNbeybBGPEFGmuRi/KfnGgw2S+CrHjhaa8lUTSUgfXrw4vH4slxF
g+45kPnLDW4CqGx9Ts5Qtz6882TnowHCMWWCL+45J4Doe7EMKNHwQ+1xVE8m151+2ssPd6/sJZiS
WaFMxrQ5Fm19cmDyLFYcgC9p2YJuTwgQKgOEQaQj4dQXMkLrRaxKlWgBPUfcCi1Pyr8z21AQ0leZ
AmOEp7bxjr2jtcGs6FotcxoIITJKz76MYQb+hjuR8UD/KvJnW7YB/pjxhIg1kzlRjb47v5Zgv/KX
/ooGXPmfV/dLIGPEHt5IV5Pa53NBHDK9jl0mIU/wej+h34v9vJqyqzZUtdhcz3rMo8z3yK3+58cJ
2MriuBwrDRjT40MkDCyCv4M+jFupX4J4PJFpPpp0Rv2m+a95Y7AR5tbp1AMFTGWa5sFQTNPnwS5X
5SSJr0i9zdcSPDr7FxedlEqcFXTXCPOVYiq01OFm1fgLFr542+ZcHnhGxr6bPzteZRDs4pfb4CCm
bK0eR3uEp7LO5xOZ2S+FRljm6WDVhl09G33on3w2NJUPvfPXbDI2zwspPJ+M9HRHPUwRHO/9zIn1
Sh9z1uF8HBzH2tJ8whr4Vm6QY/jN+HVcbFSpvh7/Vfjh6VlDWMuOolWOzB61rIDpdXj+KNR4+kmq
N/BGswfvYRUFQ9Wv5+vQowotwcL21xZl9lCwUS72PbMBKnRzycA1doArZnEDfz0ti29eoiPkNvrj
SdAkMjCYQl0R5lQ1aPsMFWHl0MFSLxn4YZHvJh7dzkHY6r+ttgen3QsfWOp2fHPFFWhhpBk5X3q5
KfOZMryj9T0obe3rIgrpsxjUec/RQ4X9+sTNo4xIPeAUlAQ8o+tJqKLpxouofliGyV7HE5ODK2Uu
/jc77yFHL82k7ke/dS7pTFZbZVIZxktcLD8D24umbmvEJ2pIL6X9i2akU0yw+2lH8/4zcA7HCwe7
DEKHuwO+ixOnqocvW0mfDCMLGoPb4wfQ2KkIzNIKVF8bu0qiRzQnpoOlghJgMIMTTpahpNZN+cAI
wkO2hRiMw9VZx950ku+Dzmk0kJMBDIwEhYmS5eclvd47z38Fqvskbq0Jq33dWX6IkR8sX3rE+Ser
8lVkS8Qyy3A0yO7aDrfNvpzgNcJ1vp3wZNTF8hNpAGEOaWQdDV7jhM+pvXufymcWH8R8yv1gEYOT
myXlcGjVToWEwxnlwh+NfXEfgDwAx5KoIah/7dybj4B3oPzgLaqvJCV5X8iynz2iCeJVCCOaQ9PV
A0jLZ20mRGhSg6cQxDzTIALSw5A3PkH8dncsu3OqAasHxoEVZD4JEwD4xG8SZirM/10ODASeQE79
7D+p+Bcgeye4wAX77qGNrB57sOs3/N1lWsjHuNX1Bkyd4Thj9BclyYQ19/tkAfFyAFSSxDDUej2d
uvPQ/YA3/Uae0+N2LFFFfAFJePtxvwXCIVe55N7vFjI1aCDSm8aikoEZxepjKA4jaiBAbaDxRjB9
31w6x7gkWk/sKdskOm+lOTyPJ4D9JemSALTSSifx6VR+HZH+1AOIYA87HF66jx5MyJruBuebfL4x
W2CfdutS1INr7R1NZNXN4IB/grO9pLIb41Ri40l9rMQpgLchjSVz9sc+3teDFpWxirTTfXckosf0
lO548+d0T0OqOls7JMlGvCJso5LeOso3hX6pgc4Zmdt92EI1e/rm7In5DyLwuGm9HllCwvQ5uMt6
DRq8orB+dtiHkioe/uRcBtIe5gAKL7nNbaoN+cgF+dTCSOcUw/gRqAthI7tVfY+i7IHRtlXOnRS4
660UhgjNnIBiYnAxpiFtV3yK11mz+V0HDRXTZbkKZFdAkpl0YAPh8+BzLkGFxcGm5rWdhaMaxNcK
OSnBmoBEEspySupsr1xRAB8XzD1EqOiN5XmMu7IlzbTOZfulWsgBXqCtqCthip4Xd/kk229bMtyz
zxOiRvkwT1YQKQekcoUpvjJS/+sNXrXv+7Ee7/kpfgG92iHLGzJmG22EgYndYeKkSZEgH/noq5Le
X8GsG+VX7QHXT7lU6RbAZXTKh0aOkE5TmnnI/ACaBC+sYqd2bw+9wOEGEGrFYODsRzFltWbiYhL6
d10PXDS4fj6y3Hu/LmgCcSL8NA/5y6GB/pbCEOHJquadQI9B6vXQut0uM43UgOjB18rvVTEc3s6j
mA5x1fM97PszQ9fXvkXyWKWwEPwwrLzlBPS+Vqr7pvny3xtds22lO66nOys6+EjHRM+MyNlGbi36
qhiv14N1UEh54trhD6lML0y0mdhjRFf/0jTls1N/S+Gj5flZp+34hJ7viWjUG1PJgi5IGsX57cgy
i9pfQcEwTCNk2rKk1arbG2Mnq7W/CDYnlIRSTs3ZDcGi8pjIR+ytYKdccQHHrviQKIltku2b75pV
vcG6MS2spayW/jMrK0gcOT9egHcDwtCgW7Bd1hnZgTydxyLAkG8LlljmFf08SgzxU4/EplG5Wh73
+WlpCWwkkk6wKVoWFYSw7VrQmvT8eaW0k9wz/D+OPjIXpxmPC6GiaClTcP6+Vf5BlU+6cxmy7fCV
XUJsnYh9CQLolUb8ms0ZFmIi1rtAbrbe98lhtJM7Q8j8M7XJeUeqa1T9AjNJN3K1DoHzuOKIfm5T
ITGCOUgTaCLdqCC5Pp47WGJG1vZZBdtYfAqvDoys/oEMT1aHzJ1mmCR0pLTWh3L82LDc7sqeDVMC
W3/Lq531ItqqM8MY1K70oawEHbsMYD4F4sD3zYjUvg8++hi64Vo182oePnYOh9dT1r7VQde5ZOfv
LP4d4NbKXYA9nnpMFcK3C2D9cDeMNXBAJy98Z1LmMOB2P8lEKfiu0B5W8PyrzHbWCbYuBHFMRTUN
48wWnJ0Oj1MpCYuiYQBvbDbZItfc7FA+WEDaXk1ckjH2qdqfEtP6lY21gp/VwvM/7NPgvJKL3N3d
SonK6osY7K7fGY8LU8EmTmgW7jYD14AnVa/fUir1avjtW1ESIn5MvWzlZ6DnZvz4IfILeCF0oQN9
8pMMA3uhrgHl+b58RNO8scqMv2GmaxjmSMwo/0FWutufspW4DbowqLG3iiOTDKYq+gFeB9qH+kF/
/OYi4JQXi0Dcl/MHMpm9FZsJ0l3AyN2rrVxKMg2H3tPruAqaAdaGtpXnvnPloEAFqkYlQuuAMXw4
1JZP/c4mdlL8NoncP92g5ss07DRs0axgAh0UNkYkBcF2iw45h0sUAx/3UWmXQKIUWyTx6JNPn/vo
G2N8qeBWWdP4eLHNidnhPTK1XF30UqSoJa7X8uWBTRB+8Kd/JQth1z9C9E1UqEy4aLiAiaEIdlz2
QeMSlSIS/f86YFjpaRjjU9rQu+PeU03XVo0gr9/UEYVM8A6wWN3XoTW93mkShvBjpMBuCoqRH9R0
/Q/7QhhmhQuL5sH0p5+JDls2EF9QMCMhhVbFKehZQWWyd0kMQWDQM0UAvjxPS8DwnHehLY6f6nr2
EPgyt+A36QmkajQWd9vueJxVoyQuzWb99rpCn/nuqap8BqT7lQpuUEhAKhre4jnnJcvsFbo+/ezG
g8uOdYsfVF3rf/Umq/tGKkv/8dNhea1g9VsBatElcS5Zb44GVgWdpSTrt71KOCgOHLEhV7EHC9RC
Gb1HWTx7N0u+uqwBAbJY5A385O1IxLcBfxGW6mabXuNvDJkZp/PFskdaQPUChZ/IpKtlrBMNHzIz
02o8fj2lWWmWSMVbIrJWg52eGeu/+IV0Z04kD0au+d4yVQ6EuERkwO8NvtmDeNKYI4Uxn/lyqLR6
hbTiDL9TBguYhKk4mpCzrqZbTwd+0DCbpeZBz0R0mb5dNBUPs6Ephbud05aum7x8H5h/yPBzwljG
tnaYeA/crudnXDkHLHY1J1LS0V8JszlR0dAPormXGhPg9xCGT6b6RStflI3G8qM94LBe0CbGIEiS
ULX3NaJragJX1EmjeAPlYfySM/jal8C3oYof1ecO4Ze1BseMWO8MMTK6xO1UdC+JaVAupJSVL1cm
JwVR419zgcIeCa4vRyhEf7RpQT9DSiOA1o8EklAHbwfLiq7OAxmO/A/l7OC+wEcOoFH3nojn0AUM
1dwTSfyESme0U2AbXKTqkxxEO8t9UGbZygz2wvi8rtS4k9+kUhTGBIMQRkJGGe4vX9iYsWVd4ul0
boohzJh57m1jjRixjk4rMdNG/+sAXTdJTRSQOL4JrYog74YG85ztcuoomXu80P1LR5RegCZVGsos
dtVYO/1QFwtS0MUR+lUmT5Ei7hXSHvsPNnXI64ar6oCOVAxHh3PpudNQ2O7tDT5ePdKrCa7PfxMq
jPR2bpCuSDA3VFsPPRBrKD35oHKSh4FdPr2xukXUgkTLowIAtf6stenqrCDJRvh6TqW4hL7aaMdq
TuMvbgHxL9ZhJtzXr8rZJ9/UEuPoTWNbSm0aVsUJOnkLD6rdgquu1TUO6P5I1XW6VJMrRqXBzZrJ
c+EQb34zQ6WciNTIM2SIN+B9JCpJ1ZdmvbpfvtQGmpkd0XumAEASPXWOeW6ILL8c2lZQ7cxauG/7
lwfQ3DURzTYVRDjLfbdABSY4wSg2fGgthry1YjFnCmt2itgDydUskgrsklinraUnZSXgRm9MExc7
Ga52EpFyF4/6wxA0KDdvMxlJyKEqsEai9YouIKx+j/WIp0jcUGRt6Uo0poBklKRLGbAHaR5T9v4c
MBKpT0TRRuWn8Q3Ip/Y8N38bHO+eStYOzQ3NLLxHXxlhSasoBODVLmK39Y4Vrsdoi5cWXSjNLjEP
ScyCX0L4W/fO5OxuoXc9PddRl0zt+OGCqjvQcHBI1KdPxx5iaCAfO3kcLh2iT3m1D6bO4DyrsDuR
JKOGLLWwVKH1UMyF0XW82qJjnXYAJj3jrqrLJJmMmFHRIlQFlX/W6YQVNd5zuUWbkizJsoBr6+tB
hh7B8Z8Q+PIW//wRapJNDLD9OjJ4iKyj6CbEC4ga2nf6u7wvS6YnUpWGwmqbvddcVtE7I8vUKVdh
veaVrRdRWjTBWeqTWRxTle9p9uehn/VMy23qthYUmuJ3SIRlxOMPJBF48h8OznMRTrEWY63hQkHc
YHX7/8dybtM+kk+DSzes3B6JMIMGdcqMbrcUwbssMKrrmEQXXuSEvZsRBpTTYjbH6JM0x8Cx3FCl
OLBPi9ePU0tBgrS/DRGpsnpAt5W1RctQUq91fSd4UJsi7jlvbuaOrG0GP9qC2eZNpwnOqDC0z8Ke
OS6RmA/Ah6mw4ySFpCB2hWV4vVWWTT+Zac7z/45mSmI0ew2JGh6LdtW7pwble7sHrVdEW1UwjjqT
2iZ4qMmNIqDbp3Z77l/3ewE9FwH+OsbxRzzK4ZUwexrEid4gPg/R5qt0FLHj8l98Nl7Tpsmzmu1g
RzlIvXAoDgOMu9JID/otW9GJ2BcMUfUH756Gnqq6jUVUaV9w3SLUVH9UyfOiVXb12fr1YvQ4qUyc
Sk8iyayqjjeMIA55B6+dsMn0mbBbOfxlKPmGrG0lQ6VQZqQJX4viPBBr0cFmHpPK+GxawaBq+Brc
U5DPLllKwIUdJiDpGOTdefn82jDiY8D6BrXNPGOcXsahXmXqjt47Y4Z5kQZrBgWA9RtpwZzhddWT
UfqGNF22lJkyD8ozyqxcL3e+/1fGFtm+0qVAewdyhMJ5ZIO//jY2nu9NutBUwDEGJnrBq+M/rDJ7
RlyqBEZwBPE46P8pTNJ8b0D92p8mhvjeoToCAfshX3Yi5jqusE7+VTGu5beoG/MIaVYK54DSncTA
e5t9FqRpnQnLvQGIi5QQTmprZzJKg5Yl7D0WCOQ30gMzhPSolu7WbYfCJvBbK+JjDLhElckfMPHf
QLASu1LK1q+vC1vJsLwmYXl9hduaauQZsxOhA+vUxdVkXy+jyKEGnArBWduS7NS72g+VzAKjDnNZ
d+Z97gJs5jRV/17aqOHNpdYeKkAVKl/4pcpJFD3RyTlhz6JuBYVwlX0szBnBc5LujLEtflkQ0Qez
M5heoyZEAO2bmKKjA8p2u3VwYuSm29Sp+rTc5OCbC1veBUzU0Ti1F659Fss2gzcUI2pPJOJBNhpo
LgBfzwJpTANtjXosvCoOyhgXz6PNiAqvZtsJK8DWQ3x/WEbXIv77FNnHXhu+8aA4YaIvpW8FCemm
xek56uoIYhyk8NrRXat7gHnILW+COiCw5fBm4WkObUSBv1FxFKjGaVqnhYJu/JOpK9U2T5u0+V3u
leiianWkVJ2s/OMd+FmdQePgK7Ail+Mk0fc4qNA4orS6w3M4RjVlnU+5vipPpjE4n2oqY4Y5NyOl
McaY809ooLtXKMtALgj1GmtTq3vNb5F2JhqoSIwVpneWpocJkzpHUp3pyTZEI6PCN/caHjX79Lso
L0SU2WEXBWS8P1cSc0/Hqaa85NXXz5WxTuAQtdWDCl8XzEwTDHq+uKEa00EOHpyxhEBOzqPjqs4F
/wp5aroKrwzOgVJ7O/SeM9SAOYGEuVEGOVT1tB6jb8Aq/Ur3FDwYPJkKvOQHGtzqxL3EQnB447oy
QN+jps7/n+OMZNAaBZNON8hGVgQz6WqQ+Ha0bWpjG6hxxuuUrYgtvaqUxNuAt5lspOSBM1gXozuD
VSZNi1OVFPNIGlS4pwFemf65z+IzPIrq3szZ9e6W4ggnDw4Nq7cHg4eH+UiiOTOzEE+Z07p1yS4x
32QJWYgGX3C4O1LyU9gQJkSZSVcycwHq0/jGp6VuTcjecxXLLZ7KvoCdQHcAuzs7NSmIcG1a83PV
rPZqLW6TL7EEnFC3WGHvwOQ9yzn4adwwyG6AA6UjuVpFHHL6wSMUS0KFMteWunmlge7W53WZWzj5
1x9q04bh6Dxxdqeg25aPrROw3VXaOvGhq60cpVpptQnxlgfHqF9q3TSDww98unjcq8V2AUNldotV
PGNo6AWJ/EBcAeO3MC4bcesxp5T5/x65McqaIWS+IV5Kimg+AqA5JKBOv7DmIo3zcVCw6WLFXil+
TOMyzordc7PMK/8ah/EMu8fazFBeiOsCw8C6LULAci8joiGC8Jd15kj1YQc0RI8EJSgtoEw8ZOJ+
TUHRGA8K3gbgGWY/GcgeVfgwA1HQs63zQ7IAu5JnxA5UvLoBiAn4lfccbnIe7uc9A3bbm2tifIYQ
wKzHH14PESlxbbZlRPLB+J8fbDCQODsjzsDUWHzkqSLdgOu86k9muizisfVzE3MxLtxNgncM/E4V
FYXhkAIdBCnYAmi97FyJHME98VUIEacguWWhQGwBxwVa+XfjP74wGP4OT3I2UKCQVHk9dddXA4yp
otzRsYhRf1UvfmhsLcbD6T7YFpPrdZLkuItpOK4Z22n1VK6GwVIIuXqX8H3shsKXaO4ZKs/J+kyn
oGL87v6qBY9bWaoweBt1q9kE7WXKztKWag/etNRaC5v2oe2snLweI+gLsfwV1T8YdMR7XtlwxyKU
3MX9F3qNKgsMBOJEtThjNFuvH5nCOmhMbiO/73ti5elrBKtx1WYuVwyH27SnXv7IwT/dDDMIwqC0
zOmMBAjK3yGt58WTPcu2NfbZ/+zfpYBkMBwoE5XSXJo0JI7NaE4m5hYPF6WBVD9UrBU4lkSh5Vb5
+4Jk6ULvE5n/EaEcraZTXD9s+gVCytbXSX46z5xFHarVtCLj4dQgLMQ8YVgO1yMHAGPeOWdIIMCs
f+qPXXHsGgKw6Kv4KYmpeEHcjq9IIPkrVVLQJMaFhLMz0J/I+K4iiy9HgH8fw//nIUDor2h0NGBK
RSCtoHje138Uu9th0uxJKriTe4u03IgNdPMRDnAP4uFNv3cIvv4+8qDonxgxFGLdatYdr9XwPm2L
iw/uhaKlh7BxMW7y7KbFhB0ji+zjMpf1uYR0jn/5P2b3e1zGJJ2yKCY7C98z6kw1uhSZiuJokScR
Drxqemf+QeNgnjfHjs3lq2LAmtP1NLF4kuz47NPCtsoKvNpdcMPDfxG9uZThpYoWXtZ1A6IG3E+Q
ezWWlgtygj2/UXFp1/nPSbkbEnRXZs5od+Un3CagBYtsvCl/dKQT3a1ENchYxhZdXMNAdz/l7ICV
eF1boTtHqC/5TwZA97f/NEWqzkbfMr8KFSPljBgBm1IpyLXWR3B3h+3l0VCZDdMrB3ZVkq0xOoN3
hVQD2kVXeZI7X9f5QQ89AgmGTYPK1vXkUlcFeNBngeUi4npMAYkSLutRW6eyP6MHW05z+BZQdpUz
Blbigi+TAkFMWXZNKUoPPfs1z2ks1t1JIpr8K9PKqkDnC3RcnjN1StEqakD8CkR3RpCaSg/Mpp02
DzUvdQ+fPp6Dib9HhMNqY52NsRJvabI1HbJnaTPSXb0w3DxBHCYSibh9PUR/0NyqrWmNxgbw8htz
EYBmgXzgy+xickeF6mVFi1nRA5alD1S7llQm346/7jcGpm1QtQJ3Yro6z4GH7cDRn3BCMREYyqA5
qZGyinlwqis+XllRz0xz4I7/HCziFSKkz+h7AqcaSLMU/ZjPxMJgExb/hB5j2mReeHdsYVVn/Od3
M/6KtnPKanigjTwwjDxAFV5y+wXj+9PyYJyOSop0IX4MEHPQ4HRq1RUQuTznHm/63ToytqHAJ3vZ
6Cb2i/lhbWb22fONBEmhPfuJW9NHVKYsSU7GNDzrFezWKbhA9oKI0bDiqSvAHXWXU1rjYZLpZqZe
hhDopYBVaFo2gJeM2FCI5rfJZUL8xYU/v4TImXqeSkSuJc72yXjooMzLJKCZAHkCFJrgySoRicgI
33yO5U3aZzb38ClEG/vS1oyDedYbcCzUE3RQo1FNSvIVHwCc1QeQ7vgKE12ECahT1E1nvfB+6lZF
5HWnVLMreGHbCvPPx+N2yKdQyEZVHf6CLgEB/XUhcvqvqsGjr05L2MpCeOea6e3BpbhS18Y8O4fo
xcCaJhD6ncS/Y6XGTUimKFrcU4ZznSfslsucOwR8lTYzibyP4npGQ8s8A84XxM9PHfSvUjzVSdZu
lkzMjaF2SpcB6aSE+Hc4VWfpaMS3m0nKqalyLFbmDYXev1tcobf4icBfvavE9wgvpZtdCCEhFmSo
81pEC7ah5GllMzRR5tef2+SjHl9zsmfjAVSmB51juLYFCBevGY3tspygrc9uu6ayG9rQyMrVmghk
Aw1PKzPJF7zdaIBm5Chig8bGzMUqu+ifPI50q3Lfi4ey1JL/E2TpctQIyleAfm49DZQlKfixn0/Z
nW2Aj+uANlgP98FQCeshlLsC4nz0K6pwKTdBmxdd1FZddCxkHMOjibSo4cIYKLPRTip14am10jIo
VT7VHKk0IH7zQM0TPPplWiRwJnFfC3la4c6ysaIcQ0Dn9DTsn0Wj56P+C2yZ1HSn1dE2RqDskfju
hZ7ALjCcof0rnCPheRTNB3s2yWgh4Cyv2g/5F8tE7uuU+4pOEaXAYbQFXrw9S23NtkrSHAU6SxwF
oR6pnKoc3bYTtMZtIjzZSnfEn7nPfBDoAyxHKFuE8f+Ylfe8xytV+70AJTtLt7Bt1ZyH8ECar84L
llpii9DakpqXsBTTxWs85DVlf+Iq9eJc92skc0hsflxqVyCHjGSani8PtFAaDfVcN7CZwOxxMZgn
PJRskh5y08rzb4p7KdKCVOyIdNc139xxFklaz5ZzbmHpMMoPcqIlB1P3fWw0RXNGLcGfmYCcM4h6
tNiiVHB0KPXO0/mi8z+9r86+ikHTTQ1J4Ko4yo6sll3384UV9POLP9e/ffNKXBGpXqZ8y7AtIo/h
0L0lWzioWHsfaWR5w2/ZJ4me5GTZdDmHfEz5nxoJXAJU6Bj7GuGaoYWajfK4ihvPrtf05AROcj7/
6W6NztiSQYMGIvKUfkr+YVhVQP/by8TMAcnT28xin0jsmf0ttF7jCgTDJVc20bZLG+l5TFnanJwp
+UjeGyeO2lSt/mo/FflxUlJ8FCBMtTbcq+LYj8Nl8oURORC+iXk4PPOGEpCHrXiKpIrFE5G81zCJ
r5yss2Bujsm4Y4g2+1FBkyBvj8HNwRX6ImEnrPce29Wz+uyvTwIzLu67YJ+Llly+pta0HGZRvmzu
bjHWbbAphbdFzMCWD37RPT0l7wnPnekAabszo3CgNJukIj+VJxOEctVX5Ltz0EJMCjqJUz5CIHcM
RzdMhv16WBSGjqZccZV7fpPU6SMRsjdZSHobNVwISEHFIP8z80I3RzxaJtI3teT+4CT24+yqFm1+
yExPthMX/YLcVyXu+L82sTs60bWIuNU10Xby5nLiHzhpogACGNqbs7UOMah5ISDO5uwlxWGBc0Rc
PNXPJk5RjuhXPT88B9Rkky5GPoFs7PaFiFQmOBtLNR78trA/WMU5qDIOHhJihzwt2m3LhGpzAOEV
UueNw55aqmN1rWmBqmPvSeDnjt8svZ8AZVo/nt8lGlpKhQvbnkCaBk/If8hRzxlMYzDlURk759VA
fGPnj4a4toKko/NhYxt4h1R2zutYuy7GrfsD8+GcR9yYyrgBZlD14W2ZzgrHCPAQO4u4N6cHBpVs
DQ/zfCA26kMPpDh8cqhdFa5mLWJgkdjvhtdGEep79h8phRdJmyfE6ZHW0GGEtKJcMM0oD8whq8vK
+cX7/0GK6mudVizg3f8WCbmB8U5nWLd2eHiiebESOdsw/u4va8Fvq8M34/A8oRJGfndy86VCZATO
bh8UUUOMVkuLbNTwUrZbp3Xnmy4eHFeXHSmZnZj5nhhKtLKlyTxZ6HTyd0jEqmf7/cfSpX0a8EVN
huTeVfBpoCBgcJxhF9u75Bw/jzgirMQiBXjMR1TOxVz5xzXXT3UBSaZxS/QvI5mNCRtiIPt21LQm
vW0wBMmA6QMz+xuqc0oopMO2nX+KY/J6l/BB5SPQF10GDNxQUzlum6S2qlbnAYSPekdL8Bsyq1kB
ozqg8NmqawZgVgg9cIq5iCoLygZi+Gadjjk8GEtrvcYYFUDcAuyMKBgdPK99Bytl3Iroi2kjrhOo
kGobdGd6IRlHLCDXGc0wtTTGgd8A0WXljBPdqoIefH58KIohA1E2hK0MEOm/x6mjnQpv7UCOzzHC
VogWtXVp8vwuNVYCDVsXiBns5Ytp+Ij5Uv01wWtlP3fPWs4WzVa0gJFb1wLpzYw9eKgqOO1DooP9
W2b2P71U+kGNbVSC4HyV+cIu+NNufw2518JVliHXjBRqQXf4CsLT0V5y4lsfvyDzKmOacvnPjg8S
tTnvJct8aq2WWMbuUqRxIBkq+Vw851MWkePRLgPEv6bpprvoLKVbQC5NLzIid/0gaJBLx7603VyT
Ljod/Q0eKVtlEB8bU4vB82hH+ju8YfUCLmL8wMeYdJ3lYmV6VlRGC1gs/T8IrZbYnk9CThW1dfKA
gaSiybW/9kWBSw39Rfi+W09iEqhq2Bwx8HvnhKz6IaCqfWp7gNjda74G7QnEglWlvKAqtMps2Fq3
G+yKr5PVZqbLzAF3RJ/vN0imYvR9/JrEZ8vK/+KOaRNBENk3vvJ+3wkBFejjJemt4rN6+TrHnO3b
HnuJwJWo6sHP15m37iTxDjEwWD8rO8fLmomho1VTV0ebpKrm6d1CSOySXPcdiNoi+csavboohtKG
ZT4aiyd2iIFfHJZt/t9JP7GxERY2E2dubShIKZtj6AcMBlg27OpbLWghFC8+x4AVUdfTSq1+MsOx
6Rq9X94aTMfoHJXalF5AuE4OGr3LfSXtIBF+IfTtUV8y1ZNxPfAOFdS4YZWnDqsfpYDAlYOc8aky
R4Ilfk26OLhJtIxRDZwmP5TOwGU9TqfWUcHBHjdOxy9/Tp0rv3avRxoLE3LQ9LUGCBJ+bQZFROIf
QROXlHq540Ln8YSrkICosMDwqgLRq03wnUraQpeX9JnReaP7FVKOKd0+ahFW7Yt625h2ES/QCCNq
YABf6r6lXaowDwp4DiMIQHsO/bJOZntcS3IJ57KimWWITRyZuJ5X0nwgGUq3lHj2Ow5ioIzLLvyo
CrvtE0OmpxYh4C6DLSGCKoj8HSX2x71Hn8XLT6NSn1G+NOgg/gqv8esJq1XgQsS2aZP7OCi496D8
ZACG678H85w18qYIosTNVh2QqaFstbO9lpwtp0kEZLMJ+iaA1hAs0qGbbSyNzLLPlC03XKzw3jqe
qMkk+X7KykXYtycmS2knVKe10jVNM3hBqZnu4+E2cuLhIc0BZ0qS49nFBJTI1HBGf+gvbHJKZhcX
cr117/nzRUlsRtS3jfALscFqnJrbbdCZZHJZXfdvMUuB86/t+3f8uxiKMzhG9chPjL234m2Irhlo
8vdsOu9rX5W8hdXSybUiwy+neFVa1zcDsC/O2DclDdA+8VFrUk8N4mzGc5HSsK5bScbr5NLHgmXD
wif/Si4stsnVzdhOJ4TY6KRALbGgapFt6F41enZhNI8sWlf14Ucyydkp83UVImRB1k4ToKRNmPs6
l7EtHpB0qvsHG45qf5IkBPtvn8HrHVbzwmKfhpMp4TQGwfxuhgzbrDp422Ax6LgihDNHu3cyojWu
oWxjSk5ZAI0T7U7Hjvp/akQg/J5CEBkkz6NB8jbP5FpMo5Gs9KNb804Um6qZ9jTz3cSbp+F9Q21i
Gpx/hJGYAHWiftfo5kSauGj9isOhBTTtZkCP44LOPc6qZ/lL2QIERLkYsvIXwWl1FH3IbOfXgsc1
yXT2wFNRszQ31twnrRPT4qGj19TUpm4+HJGH2TG7dwCE3IK4BUCubsrOVcKmE/wN+B01A6vEi8Tx
x4IS/O5w65pSJDUYv9SGsZKIAEU0w6uFSUhEOqQHrNmWJ3zYuTQ1876BfGb3ZxbOMiQC/W4z1XgP
531Ny6rAuJovKU9RvTI3XDUdsq0i7a2S2OrBwe5hMXZ7wcntnh46MkHI1iIq9hNGqIPANwftN0eL
K7ZQLRCB5agswIv5wKZZ32XaaKsT4p05OCgNU0vRQ94Q8hjZKhZbOuhWZTVuoK+8J3ZcnQhWFw/g
48HDIr5I0RAurIYsH1Zp71dH13lBV3H3YEspMrY3letY8SG80O9h0WpoeOT9xB46k+sAi/sx2vCk
1zFUbAPSBK9j9z4jvS3Sz0ePu9HV1F9cKmcBYigYP9NKfW/tMpf+Q5S08Y7QkuCnIH70SKHTWBju
5v4VjEVxFu+wPv3V938zrinOozLY4SnhWExN75gfgOAtU0XIMnLmlSBpt0Nua2wiQQi5U0Rzu4jU
PNRehQiXi1jmy03fKyIBbB+2l0QAr7QGwdgK1aKt7QDqqP7JptiVo/VB8uWmyL73MIuDYUfFFzZr
X1p7ON7aFIbGKXSKKmha5EXlDP4My5NJvdwQNXh0BFYm0xi6BfyIOb3qg0ztcLkIcqx7C2m27IHa
KmfgYH6JmDBwASm9h9XPnRMGKJbuYmUSEJTeJ3GIFW+tTiXELKSaKPd9fEkYJ3+jeUijx2qjjO6H
9EjF/H6HuqyDqs7hK5LrTHa2dHzw/yhRBtuNDVdz1amnRj7rKVZxEAVviO3RPLvpogJk1LES/iG2
vwqnXgDFI8IiTeIQMr9jnphKd4yYGu/148yZkKWi16oIhn06NooR+Rcv0WIoWRM0Ww4MwnEDKIlg
pRtB2lPd9mY/WfeDV6sXNbh0Cg5sEDSkrhX0nW2XPHcYckL1EL+D+w7Z3ynnGgihd1fF5bGMdWd/
Y0O3pW/L+exrmFUz9CBbgHIYCe7osSv9p4Va7sSgnfekQ8VnnYQCPoG/HO+9jvd7W9s8uW3p2Zqt
9dGmhg+gcLTIkgmwVLYAjU6tHTg7hMvwtRieJMYpLuL/Hb9VLJXqzg4QarAyw/WCQKwF+d+F7FBB
jYeIOwTWMOHCZ5z+loc18A5Ksbz3zg3HyXQXB20/dy43JuBDwpHOLvacHaZVBjRbAn2vkfPYsEki
Ax77i+pP8GiBBif9YE0oJ/oBGoBqd+esSfQ1DYSRiPa/5SOIHNIZxAOvc4ipqJliOw5qAsY4hPP+
Qk3SWtFOZ6NljqQ7sumjgu9LhxBMYBUhvIaJlsKQS6WlvQ+QzYfLUpZSagEIlzRmgKip7cJsRfLe
jJqGBbVD/wSSgmXWQN1IVZ/u7hO29C+WC+ELwjGtVmdbuBzCnZuwloRNqYU/2FFV0aqM8th8l2L0
ejbDhiiR1/CE+rUBxW5GIX2CPlv0d8o6+SH1CuSekh1sTrUlZjYmBwDdnzauxcevUmvC/6INgGWe
qDV5YqyMCtYHwMmbdj475liBSDDWjyaa19egY3VfaYfkrwJbIqyGq0liDHYH8RZq6qLkBPTLSn0b
lNsHt8NlsAh3MvicP8HobFDJuBlXglMD9G97i2Yqdpr295SomM+c6vKPStM8syUmHwmrBVgJpBTt
EcSs8oZXz1aafJ+s3S2lBw1QCffGH/931zDSH7tiZfKdb45mXh0qtgwxvhA/jQy/xyFyZ2tU15xl
cLW+6OiFMzz6USJBnmYyE143U9AximsComYr+8AVTtXQzN+BV6si4QE5HZVb81LytkrrDBjoY/Xd
kX0NwSHMVsNLCbgxoZPXhZzgNsqWcZg5TvSz2o7SoKr3DN1oZIjY5GojPj9yKXRnWZDAGj9hi5He
803O3Fyb3Ca6PtPKPctTUI7lxjsxA1AuYvHIQg/iaCm2hystyfG9b0GoEIceB7FZUTDq/ipPZIbD
vYTJ9lfkihVZ5+sn+CS6JyxxJaK4RP4vkdnkmpXQDGAdt31geqoai91ZKE2CGskS+IQjm5vkhcm9
A5Lda2RgBmyWrSus7OQBrdKRmZQoAQWG2ymMeWQvlaKySAoZoMbzwbQHCP8fLbw3Gj6L0tqbhEw4
a5nmF7ZjPY5EJffovBkM584UVJuG9g72vc2Q41jAMQ7llSTedepBE1TOOHrFzdjauyV1GezbkWtC
/GoGkV/55elLCLd4BFYXgo+MSDcEOi0kc1SNcp221QzF8G4ImZH6aHE5x4F0uOY0AGHqGmIEpwNS
3IO9eynBzKRNFa/M2B6Vs0n6N5paw+fB2u4iFvnlNDyik4CMkazALGUpzV+J1BvwBSR8Mk1F4YEv
I1mZpxaaldmu8JO8tdCcsTe0i46+OFBRJcBbArMa21dVERaNCEyVapgGsOFk+26RT4ylcjl2YLHl
Xntj+T2+5DxGZqRAYVIKyaDBhaS3NnjUuKg2VcpTkm5p17id5Q0ywCOipJSMZGojlI/TlVX/KXsb
j6Dy870L8SxO+FVvaofAtQqUIqgzmG373adkNR7NVwJEWl6hJ/J2cFDxrAThvPnqvYvq8D4lErR/
hLiQni3C1BU4TqDwwym4LEkUeOHmqLH6f7dnGcbormTDnlbp7IN4wOdwkmm/dgh1psXdbH6t8O5d
L/RZ8kDGk7C4CboYnVm8urwHosMF5k9XHKEVZWXLDINqHQa9hlMcWMZm/mPSY3xbfb0xZ7W/rnND
9pdkPh3U6npe/sNzT2NOfbPITzidIroxnrCd8B32Fo4wswOAYdlmOj+J0ylfb6Oj5aJoSxOggiH9
jovWesC1XSasvexwucqehxTgt1ytnsuYAhErHl/N8yoE3uZj9zdK7ioZaswc2hfHycccLu1MVj6X
BiXAKx5MQDFiFcfjkjUKbwVk4VR3lpZ4JutJU6KGaeNhEziSwG4t6P6Ys1gCmVmOBdr07jbfLtq8
pge9RlIn2NoAlixmHtzlxhYiMDQo7w7eevc543eHzFLX76VuLw8Ay7xLnCEBdlpbH7aXO7gRfdq4
LGb0B3t/Eul90huRUcwRENuw8AqMD2OzLe5s3wiJD5+BZ6ctRDLY+fbeKCMt6vaweKBmLBz/i/41
xgsCJymskiapxYlMDIaUvX+LWatorjRgLhzvLu7QGtLUdQ5w8PMsXq5TK8pyX1B2B4EEsnFvsRLw
06vVVJLyee/1DPq5p9NtjYClImMUCIMkyk2/GiETJt8IQrmBa2Niuw1m0PXTljaEtnMMQRL+NPbd
Bql1LK7xTlafBb0oFRxxRemjAS/KRGGBXiFrkoDVwoMIqbB9p3xoYSaMIYAWgn2UV6Sz7nXbI+lR
iK9qovPwDgyS57HddLXiyEYVHoNKT8jPkNQLZj1UQseCa52BlRXn5TiWsFHxuPJYYLR7fCUALXPs
JU3o7MOlWadqu8qqrxXmWHlL9LF0PZaLKT0PuNCDl8sJJMCHRZoJNs1ZfBhJTlHWUnr+aSfSDcOU
T/lohAzNNao6AiW6TApbnCX90dvjfY+l4W5g78CtEHI3SgeH4O57MjG7y1gAC2Y159Pg3W2Le5DA
DK5hhnmvyDKutOLmKTi3OphmYyGWhgknETs/R2gC/ukr/GcGMnngz+77M0AOQHgL2scSZjubyvB5
XaesQ/GYYpNHkzsgS91JfXGSWN/DGys4VPCET/P+kgKOg11ZxbdyAa6u3O26qPA9w9sseohSQX/X
DwjBNwFa8rUdVpVvt8fxEJtDw3HVGmEu7ZJnQ0E0Ub1lcvmz30oD9aCDWplfkxktfySZTqwmJu3F
z1Bf5jaG94pqCnLREuzR9YfiLYMmfyl+L2BE9Ii+P6jbnUhMv2yn5o7qQKA2s/XehiAeU5fQAvcP
4Ws6rJyahtk90y9QARX2/0iW+GiMRjf+5eUAHUHMD5TQbADOk9pKlN4dmbP49xXoSbi3F6uyR0SS
HPgYoqG3jKaKvK68Jqq+iu+nC/ExphMa9xxs5fCkjxx00cK1AvG8tha1LvoKZ3hYwXY2UrrGY1RC
ZAicybBtjwO8kvBye4M3FffpTsXC7Hr9BNpRZQi1MZKlBYho2Kgyhe+iOsHA0oG5cn1zKXTd6wcB
s1Z+W8O6kIbkA7WbFUP8qqfbL0tlaZabfUtbwHpXmJYgbtnGKB60Ii7nmD53Lum9ByoIh4/bkcA4
ZW6y53rsfYmCI64Fo1VKVZvk6MbofnTiy8NTZMzFOCLLMlprgx3Z6B2HBFeii6HYdL9BbexTuwp0
aFY3/MxDlKF+iyfO7RrYxHaCBvFv5CTq7n8Yq4M4uQJ3jcHh6tu85Vc3VMZJCpZuf0L1rSEFX5q4
2U3KqbbxpufFZGWbtzHTTZAzz2riMXSmvRv56nkIHVXv2EqEwbE+x97/V1b/27+gzxquYKOoYytz
KKDSIls2g6kFdYI2FDSkRlBOpk15O7bnCR2Ed3I4mZbiLxg1cyDZCMZD/kc9DUukfgCskIIh+8fq
k+vyxOkuRTpoyKq7WX3MLvLnJNAvGb0fw8IXPilJyhHxL6F74rajtIj2qpfnEuevBQHDuuSQ4B9H
0jxkDPoT2oieWH2THwL3UFGI7F61dUKUeZvNwH05eY04L5NARlYU1rQCBO8PPzLGMo+2uzXjG5T8
RAZ1BYeRbhvVwOd5clJMBSraGME0eZuer/+IgHmdISv5GuaOzwg1v2wsa2PO+yI9E9GsIW7QMfiY
ShxwY6KRxiBoj8mGAMmLqEED6tl0d1CCAMa+AnCDNC8La8M8cCSXm8jFZ3kh2pxVgA9vU2Nzy1cN
RU0F77hSH5X+g+g+n1Zz/WDSBwQ0gqb6nca32v8Q0MMGPGCtbHaH78zStEmn0QviEZrCLYwL9Fxn
FLRTFcILuCgskPKj8RO0pXgjitndgeR1hSsXKb0pCyShj/T9rhxOHRwUONNmEUB0yojDc5suBoZS
FHXkLdCITMGnQemdD3MExqm2PDIiarq5AdHn3Vgbw84ULxxbgVTYSJcj0eqbCoH4JkkXna6ZWjpM
McePQP493TS2Dh+FLxG6J08gldkn7jajXdMkZByDejRziL5NiD1ooLSxCt4RXRqRXUmzf153T5Lp
A8corSv0nDvY5y1y+0roWJDZK3lym/RyQbUIZRTf+4LmH+MthTWYLku/IKDzoYRxPZKGHPzteBu1
vzSKH2EzNDpV/UUhrdnU0iA/OIq0UKxBxwMXxtnXwheN3bu6dL9DDq2L+JnKkVJB+YXSUSQSnonJ
7LR3e3i8OBhznXHIjIFsxZhEPVYS4zJszsbTJz+pcwzc0WQRTAw3vbJ40Rg8DTO0x4eQ8p11edL/
q4ZcJ17SLBLZUkCHTMEbyY3dLQnPi6GatRvd/zaBFDJZyeFxr2tpGQb7gIuXLEbT+LXKbtfpRFw5
a0C8DVsiyquWDQc0U/OgqoNHnFjBe0IaPO22ToVeRyogCZZoyxX4wDrM5ex84la70UShUbQaLQPi
gK44d1cnbw6L3O4PMv7Vn/dIdx6BqB2pO20wP19BH/Y5N+wAd5/CBpK2stTEIjW0C9cv7Ljs/mFF
Fg7nTlmrmJcyPUiZCrLicwnDQvQL3SlPZ98JH82Ou0SrPWAWAfY36V/m+N0z0xYIetZ1cMSLs3bg
K1tzuhGHpwcpCFAcGItpTloJ/heJvM28YIzv1Y9XdqYOCuj4JbWmxTRXhaj2YL3GVgsGaht1MUfj
eNhLykjMxdQYfvd1Q4d8z9+wyqfna7LSftV0a06aTE6gaYxU3foivkuPpcGTGBp+4vvTNldbH83E
FpmhPeGLzPGkiaW/JTFoG4nKcs8tIB8ZuCsBOFpAU0zL8kfc0rNFseBXlC1jaGDjp1S3jyIV5CtV
zt+P0ES/9+cwtP/0fc3qUfNX9X0Px2HUgr8EJX1PJVGkq8Wg3s2Ea+/X5f+Zqvywx4CijuV2Bjoe
OFW0LSBB7jbXOEwPetekOe0gV3pN/yXiFxZm01n25IinOn3K6xyD9eeGGvsOQqrSPCDHTS65O736
OyutbZFWgzXuMnNSzFVtOJ76Eq/IMI3UobIhgFvEGbC79v0DL/P5a0kH131pKw+Bn0GXUtFdNwrV
UeZCEuxItGMEDcEuKcEpPCIz4HlCTEUm6REtZgKFrevfhuOFXoz+eWTABK+4CHsSjqcn29Ew/hqN
gYnq3DAEujo9jHkD/LspUEF2/OBW1EPSQBtNA/pd0+6emOK3/icp7JlVZnCYbA2ZtxLGYsasRt0V
0QKcwxKgTqOzvEZjcxKMkQRn4U12AK88eq6jeLMY98ixT09YwZlKgrYyC15gAe2DOaFAfObFNsQp
aJqfJA5/n5olmkdfInBzQl/5EjQEVATyH/tEQYB0OyDiXyUkN+4nc8sDAzhRi5PBsJQOsSRGcNOk
0U9RqJzEkOYy8rx5C7gHmF4KyW4Gotbw9UnXkZp8Y5Xy6dEP5M8Xwl3km4oQ48lc1BadfFSr6PlU
kIxxuMHihAVk8khMULvuNzzMTvOlK5q5d/jmmLD4cpiVf7hcKVeIMYeOeIOy+1um/gzjHVbaGNQy
XQHh/JIIYG++xVyKC1iW+hXi0zUAaIGcYhPUmxf3mcBUAwGi+gqMD8EhAfkef+5jyUUnAZXgb7H4
O7xoyFzlZDRglwzvh/sGWRFPmqVinmqDUhtaAwoVUhNuFOrAxDVjqWu3O5gd66m7s865c0/4ed90
5SJJcH1FBBNTJ9n9yx2DyqrbEesEyVmVw4PfWmpGqz8lJoNWISywtsLk0AJyW3QJeWyFITQ9Jo1E
j++puUJmA/FMw2fexP1Yt2pdTapeIms6i2/xScUV3y2siBM/CH+sXa0OHYML+7g3ly+5t/yFfZ9L
oE9Z0xf+z58RVmUp+1kJrm5m9D8/8ZY0a0Qu7PIjG8jM5a/IubvaGO2tZArWwcajhAsXKQgiDiSt
+VAzaN3nmd+Qdkkd6cRIN1vAGmVEyMWVZz1I0tCvNtb1MK5cwG4aYa+4EqUaQYEPKO9yWI31lCjK
CadEv6Ns8Z+jhyqfujlSz3XpZqoCA+1TS0TFzhMVYXB084veALJhqXtHjQeLPjN4CRy8BsDJW8+L
K/SeqV0CBkgAyiUAlwLeW53rSwWfxXKY9r6+/hMtwlvLKO42dgWQyk9O1CYGyAPebb0vn+m9vFKL
8bs+0kyTYRY5BYV/yCvbVcBvS/QP6hkubaK5XVUk9L32S1MgC915LWVY8S63NKVjNJxBs3hZLC5Q
EtL64AIiR0aUT8/JrtTYbmfA2QeqlXooYMoBOKqdbvSIg+6k2z3BCInUL1l6mKKYFjnIxhq+hxGc
OPCVhuhXKDS3O2Jyzcv9CPQTNrt8V9IfM618GCNC35wjY9iCpf3WgLRllKcuUcxiY2ABrJkIRigE
vJiEll9DwSWF8To8doxJF0GHw3ZEI73LdrSwP7MXxcp3NSHwSy8RVaUncboxiS9mMZFtQRVrzKrv
/f43NToDRVLIlhAoixd8G2UXecb82JDWAS/okg9xo6ugwzknOQYSht6d6YlUBqqKqfC/CHCb6tjQ
+Cn12tUhl4riuxgt7EPm8gCUvO8KjIikULABBs6oDgrInVMjATv6KvE5ASKou6VN4ZYwk/QLU4vI
p4FCKcrUINt82ebdPjjK3SkNhAVdvnwlqMbHd0wmbDD1KxWUGSrf3zAD2qw9wPAML0wu2vTR0wWa
Qg+Uun9BSeNR89kqUT0XWGNTxTIEfwQKFeAw5FzLO7weQrGUOgHKsEuzjhtltPUKIeaBODLrKjHc
Iw36lZDZ8i93oEsrJoLMEK5+gxuKhWVi3miq9u7Ugsl064K6Xj4aH4zHt+Ig75od+hjs4ECA2SeG
l0E9AO9/8+ieFwOgW353C4L/wyK1llIaItEY8zMaGC9gxzpwIC6hrYzvhfRSZjXFIbBYHdnh8+7V
lVFbkDdVsvvlfjZ8XpGzRRauwhcDWBN90q3rt2Kq04X0YGgy4aFhZKyug/QI2xW9PvGjR3NrUZdQ
1fQt0l/cCeFzxfLwIMZQlBKbNwk/WvhV4AUZ5dt/2GZSvFQRmmQaeY7I3fEW7GnkLi2Wg0TJQLxZ
quR6Y2zUlidTxuk0iCN006kvYrLJlFBfFa9sqaDPCOeD3e/CRK4EDqrMOw9KZMc77HpXWaDqGq4D
uwoRoAKEvgRfHAk6av2xL6+KUrR1Bg2BSarsZf2OhhPqMjA98C/9IgXDTMBC0FCgUvi5c7D5YFtg
uB9BD9WmWjclIZOtFcq9bJXqQwWt/2yZYQIS63MTczide/3MZ4LOHF/OV6oJ6HKpWp5Qz+pGN8dq
DGbSL5oMDwZQXypJm48tP1ReWBzZTuYXb8gjYdij4pxL/NOSLLUMb5JALSk8WNt/nWAZlU3zPvrj
WiXvmgq9e6/xGa7mEfEeJNCUp9y954R/8WKqMaZGJpha+7ZWk3W3R4Hy33JaL5K9EO6r/RtpXYp/
EgOZSV6qHASZIjHz3HNCdc5MmANfKK2ME7gmM+vwiMYDnny7ZdsRl+yMzfo/ysJMbZYsBLmQAl77
CGHX1NWWY/QMgN2ZmOngAIEoexOs28JxrUHqKnLC4/VkOZvih3QEjSlMQ+3e2GMBRvhBn0CRrIWV
/ysh78KAsUJZOk5hAv6ljIhg3r0ANd2iSoGFumQx2pIShyScilBlBrpcHVtbwpxN+XAfv6XuccGY
LKLdM1oEWOwhaA5Uu5JBmUhJxfX2zycdu3Cw87PaLNRSCFPoHOjo5U9+RLwO5mhBR9enA9+zGuQS
WmqlGjliBfhaDQl9TF826Alq/EFs216FFlxyPaHwnadjXnLlmcyE3+w+faYMVgzsbT2Tia3Akly4
WhRFOJ/jd9hCegjJcbABg2R40tWZYnv/UWj1FkafKtUsSwNwZoxqhTRUT3rozvqkoLqviknRv9i7
Edw8u0KkE+m6e+cY8fT6pexMCLWV89SK0Bpkb+ffYCBFgyBfFsK/Pt+yhx+qSzIj4BC8+MLVCNbl
XQutZjALggpMtK8dkfYkaN4ZoxckfH5fgJNE1RS8MZDog0pC1U0/bdAy2KAFLhqHFQj2726ncF7Z
A/PXYOLnwV30z+Y0QCZipZeEH/ImYfQOm6yryjPV15S1YNqs0GX8d3+gMBrUTGFV+uELuYdZjqCu
ZHyEhlMv67TyaN6B5Huz4VnTvd2kTaFQsGo6dWZ5lST1QEBX9324H9fV9w2mMvQDdQjLmJb5SisF
NwKqO6X5BtGJtq2lFlkNXJNH6Q6k53VfekG9A6OkVlx1PKmsiUvUTRPWs/F03YA2LdEZy2YW/1I2
O7ifSfTBCemvMLxZAssLwcatppHk2t6rLNDK+csRJWnchFuUbkdT4Clr6Rquc0MvEe+p/HSnp6vl
eoazRErKIt7Znv1jAwGLWMKJpmoj+nr7dckbfBOeCRHLxKkMWqG8AdmBpdmgff+ZkKD0B4FfgoyT
FEydmtlH1Ap5ev6d8i90Bi3xv7uXMdaBUOiooXUgtCFw+JCe7MzinI1c67k6vTo9xbpIxvIbfoLE
5u19xFOYkGcz3Ip7yzif8Cgo6gTrVcloC9NfnUdBH1z76V5wOL0836fp6fUtDheQHSS1/SWh8TGk
I8Nj4u1n9mkmx0cayeNX6FMKUO+FVOVuUD2A83N3sr8ApnxUcKt0v6j20CI+xtCbOdego+IjNFhE
MXnWMaKZeJo33oLqJ9bspMGR5ZpRoP3de3F+Sz3jwDTIWI3m5D9HgwMZxbE2ejrFKWmaZvFm8xU+
bfyiGUVXniR976O2y+m/3f/7I5/+ZxnO1QJO6OprvDwW0Y19Jubp1IWuVQxE/DNFceE/fNqHVmCl
exuCgn3fyvT9wD9BK60nrIJdRhJKkCF3lkP/2zcwO+2on4rqqJuP5Zb/Ek3GVrcY0dVdUpqCeZcv
ykis3z3IQqXijT4Hv0k3FEkAaaNQO3oIgYrT/NErF5hZLBhDfHD3n3a1C1mdU/HZYb4gFrhYFqr+
VCz72wC2rFURLQXNBG93Iebj8puZ6YDmIFs74dpTX44Hc/SmUOs4htG1iuEWXcE5vd2hurdqUVsq
qBrgGFeJMoujJIiH/LuHh2mem/ug5HS3jLCQ2q6nias3ezodXoVwXrR8bZ7ueFck6D7kQk6hckiQ
lvwK5oa8PQ9IDi/1zj8bdaob1rIcrZeKnJ4qHsNBW6lalkd28enOKuTU/HeZb3ItEDTpjFvuAg/R
f7elQjCxVXckuOFd4OzxHZFU39Qq0NLnu8vCWLNPFO0pYyYiuyz1DKO/ZSkW/k8U/aUyHDg9Zg9M
e9A6/qn9mqjNKx3oGdi2E8p4gJp9RrtF4KrLIhmdonxpFGohmgMaH9aQjTlTh2czv0X5O14qs/wR
fbIlfqxws8slAz0fGFW3B4A/J6GAlk6+7O2G3GesUpixLUBe6Vgxas4UVc0IgzHdOqXUqRTWjsci
KzcvGnG0VNWGOMDC++k6ZD4yBuRyNi/6haOOicsQzXp5yP06j6sdBfWDdPtJFj2eHqtQr1Y+KgVd
v44E6WZdzjWXGA14tIb3mceTSVBY7faBEIL6fmjIpq6EWUuPDS6dQUEVhb23Jre37FQvo6kGJrKL
6Czv35MMh3tWaXlZVUSo/emRjtk+EdVrlLMmx62Bpzek4YUFp5rUz08kS9fodDEsX4dsC/9lxpTJ
Pwq13GsRFEtqotA0jvxPveJigpOnn6y4Poy28iW0Xv/Q70xZeIedHjBEhAXOFmI7H2uS4rP0TyGT
L2qILQDRrRgw55c0s7U80vyDna8ayAKcki9AMn+NaESdOQ921qkR+lXbVpW/DHsHLtZCQjeXs+OH
lYfhokR0HjYSypg9PDqXcdAu4LB3ETULfctruYtuiVnE5ngWNHPz8uesZwcd1r8Qw61KPBb+ESIr
rRBgR+w80GyBX4byjO7LE4R0Qkdu9ny/QbpWMmMlJGdG0FeWqu8Ryi8AJ5GOaHdQresqFjy0Z/SM
KmYQNqwysxTvjbSp9mNbE0vC1AYlHKt+u3UcdIqJkND/qEd39c9Vlmnn9Nv1OhHRI5rstvWddRUv
+gkgm4u8GJ2l8Un01RgS1asD3Ygj1li1hH4RyndItTMg/TBlpdV8CR+Vi3ObsIAqj1MdNipedAfq
7WBO5wEfFklNcVUtydmuIo6g9+5FKA1SsNXCJVsJEIt1VrBaArFsT44BiZNa73qhQwAsKD3IE7Pe
LQNHYqGfDLyLD07zE1sWNBB/6ojIAcb6tI7Op9YQpgxfJKg7jlyIxo/iPTKSxNPARTdT9gP9/MGZ
bK7HIr6wBC5VBSIibc+ea5Dm59+ez8XhoSaaYvGKJzVHHdaH4ih5kq4vB0CMcY6xOSAhNiXm6oed
EnxhOx5p0NHLIPokhphr8thgVfbWWvRf5c7GpN/g4i2kQpQdDHXbFBjrdScHS1NCQDayoAi1xWxQ
J3d2uQjzj6jJOTC4/yhs2die9deIhsLhHvPR1336qXLAGQ8LQ0Aiv51Am/BSa7Pv3MbOcxX6+kQF
XWKW5smUFqPy41vR4PxHfGv1H+33YVQnL9sIq+vn9b+KwevSPniFGIM5r4DSVu4rdPI+fvelsF93
0mMvJxnIxrKTWCZaIai7x2zKb5Zstw12vGKsQGewhfgvu3B5BDCNvOzCUD8QC1qSv77HOCDQjMQh
TeBaHVPHM9ToAxcO27u7uSykY2I+AgjuDHTzlD/Ny6HPdKcFzxlrlFXJhqG2x/Oy5CbqhyRY+1Jj
a8C9YaQcdbHAzv8u6oIMmI7A9E42Yy1HcHcYlNbz09obRqLDZ3HbGq8xHEbEV5fcq+N+orVi+k/k
3PgDmfjqdQyGCRxZehrg/Z04zJ9nVkWOI8ssIB5tfJE8+EpPvSiuiVVb+LWS0j2CNmb3KDntlSHz
Fj1Gv5TOnRwpqGa4W0sMTcfzqnMmnfuIqJjxcp1//ETEX90y7PuGMXSOgO3XMtsqrsqOW18Rcj8L
RJsQJ1h9oRRBy6mVIZP+JHFDaB/YnDlhbqnTf/NqsKtq5sp+ysaJ/5DZ5X9RusWTjoBphEcq0g2i
Q1im+BeDJ4HuwyOA+oD7tk44bAoVyYZrvFwdW1vvPeGPmJD9w8XrohMh8DGUUYgv7rWcaLD93KAM
+7+oATRgbSRhryBSgNiMCE1/ZbsrVZuvVGKOg9dmBUWknWo0qg7/lLyeiauB+k6EtrGb/IrVDt4L
nYliSpY/RtYS0SlzeDq4LRCpoQPE3o5m8rTt6gX7lUrKNpH+ahcOpZ7NSKtwOMXEyrZLz5/h0aRF
455XJQwuEotj2foojmB+Iah/etzG4tVzQbu3HXlurkuOO0/mU3UJ0uDciI//nC9UYew8XjImOzTw
nePtycLkBYSOTajsTFlzpOFLSU4UPdTsfICoAQQn5FU/M0ByXRt0wuzJHqpbAGkXX25enPlBw9aV
8D2i739VT1OH5S5coEKN1oCIVRk7im8N5EVxmZfmSLxtdm9E24zOwxkZTVwvNG2NBCzjd11UXvO2
Ga8jf3qxj+drMDpxj0/oZcGzjnIwd6xFqcrL42pcU8sMPIdx8IaJC9sL+UHf1Rpkfny8/zjjaVbY
eu9pZOpLasgv9MM5mWTMiEXf56N3bYnYAcC2IU3FsEl3238OXHUPCcmsEHS2bvGN7YCMflQpfbdi
ewffiDV4nudatvc+dlz2SHjKMzBM26ZHUoTcHzFz+fcd79rD2kAiqlAu8wtsvzaXxw5VOSSzjzBl
qmRXwqrKJRKOtpDxorL+oUM/fBn4Uc7Tvjkta8BlFfiPNezuR3Y6rieWCCqC3sCEW7zE30cneoVR
YAVNI+od0rlyRinsbGwpf3Y0HEOjCUuKw/+scZVXPCAfNe2Ohl4b/rSZGKJ4qqtl3ty/KD7hQC7c
FIPOqdlMVupEseC6hUgn+NxVU97k3S68lJPhAMIcwRDpCH4Sz6zE9GH++RpXMUkjVP8XiN3/800a
IVo8OEHCkkqVX3/p7Ktovi68Odg+9Jl4BH8y8ppWd+62an7amGRXvm7rnu5hedrl5EJ1lUnHDh3S
hYl2fenYw5GgrZXztKZ7A0ttWuDVuK3r3azqTNajkCxusFTVjMvw+A2/F8l+2xLh/CIAbxrsID18
rVwKTJ9LxzJVYannnSvUVm5ShrABCZPN0OOFjKpSJJ7/ddGJ0X06a6baO0mPEjOVTjeJtnoV+sG2
ROrziSPV7LWo1kTEgkidhxJdNhkvA/S4Jz47seXZRy4TwUCtU1olLxJIdADp/okdIS/5q9O3lVX0
4N6p0hEJ28I8J/ZN8YM8Mivy6aFyEYOBZZ3vqD37uQQNLioFNTTZQ6VVZ2/27SzRUNVoqsyzdDUI
JY3AvRcMbFhZ4RI0XBKJ4g0cjRUEmm3VFERHDcOxNJT/CtTHfcAI00ekr2KaQgD+AyvvVrk6s2bz
IXuRTWJxL1uziMVxwK+ll9aV5DfZKhq+i5ZSIK/N0MMlaI5ZNcDR1GEisnHr8j7d5gIFk+Kry4SZ
J/d7ZfRxmN8rouHqGhSPvvbxHgr426KMJ+I1HsslofErmBFRnos/8iYmpo2F/uNej5GwHPP/0q6t
g8znbmXYdJYIpr0MlKMDVZS4Ig2DmfWZhD51qbvoRv8/cgP12syAH7uMWlTfrD8RxdlJ9mYUAKy1
j99KfCK5pRX1Dxf9y/OgEz+Cmb1XyGjGVO1Twwwb8596+y2nmChM2XHoOx4IQzfq2O9XDchie4m6
ir0CcwyNGCQ+3pwI47eCgf+rwxyZvFsma/l7syA4DNaU2GaENHS+2GweBqTN8X6b1w9F2Ed4s0JF
6p4P9X0i9xaBZAaCgein955oLKKOGej2v6ruOBunErUeyzfArm7Q/oNZSxrV7N0wxLEPJXyOC4Dp
NA5+t13rUjLwpBEkZIYhP3oE13PX9XhcGhhDCYq8bBWZ4/Lquff78D0xBMH9K1+C8v7KYUYJSmjv
HpN9z85JUFByY98aDZd9gwIpXvNIlC/v9G0IlqvpoutE70RCIjG4oEp8OmW180coyoYCcQ4sFSQS
cVvgOglnHyE0NAdC+sTiSW94Ou5SBKftRSObCD0snXtbPdyTJvdCy9YGaSN0Mj1f2xa+SQLEHHGI
s6mBnbNkOvJJ8GT6w3dkqYi2eG2hHmSpwMMwiZ+BCeVJ/hJogclwE+9faT8EoWDUDt7lb2EkJoji
yWwQ8UXOj0330ZSzGknKfT4LAjwo6pW8GOwWwZNVqRxtkmY6iKpp55jxvU64W9rPNO/emAS9wcPh
H4CRQqGY9C27WJIaJ313lMubk4Q7TFgrMucum1eEWefK5P/q8ap4WFwxumcZcXUNM0V0U+qxbo24
054lG2rdNJif8jERkRBFoGeIHriOPArgkpm9atovskNVWUlwye0N9xN2fOZuvqRQfbI60IywQ8s7
OX5EHwLRlXzmDhCP6utm5ypuykVOto1i2dtW6/PUeSRvJio/Eg4DeCkBwiQaRNf+D8fB2cWaR4ix
EVZPLwxLAIanm8sLkHRZQMUTpRCEGePOdI5TBc7jGQgaDQ/UUYLGzVsxRbDvVmQBGQUDGHbSxGYa
2v/tVDDijYocb2GwRzgh7acm97bXBPyJZJK6m6qzxTI/+7rpQh/9O6jhZWUTorwobUB0U/0cdb0G
ZDDMjRWVNVAwmuUly4W99pEaHcyZ8+5+6t44T+FTb8Mrs2IWd6locwE3e8FLI9LMYaOSaEStWWOg
NltEMEepGVUEDP2WE7AJAoKkod3jleckWz/irwZhfBIPVnOcapBw4XA/0EoCqh/ry3Cqr+7BDZwj
D6df0bn1PUrWSAS8jftljcUSI/PlBUGY5eGr3ig5xgDOW37qmujO55FkLUJffzFG/TdiGoBH4m/L
551hr62JslSQz5L1pQf3OOfej+XJoITPbynN7f3HUkg24XVCHyhgmUosJrIo9mJtGQAAiWeAt8dT
mDCb92GfJQFJdeDjx4KMjYD/YdppBHfPtn4p4UJD+Znvjf3UwozNg+mBxT5POZJceImHmgSqUhb9
PSxg628tbNjyiDSWicG3/zDZzM4e0UzicbbBbZ+KYeFDEZB2L1DkhaWOdTIzUJBTrLLVe4FKHO8L
fuoZY3TeXRRpN0zn/3C4llnQNi+5mBt+BPQS/9rFsLZfLa9u7WWvJfv/vunoNNVbxhYAsmBCnJgP
ax40FgHIVEwTrQliri60D/JUB6kq0HUjCyAKGyOowNN3pmKAgKdSQ/IPqMPfcr/NGXc8LEGPlG6n
lU6bZGNyredTjSimsBgX9xEXJucYRNdtYlwxyQbK2Qut+5VD2miI9b5QPPLc/kUZOMGdkbWf1hx/
ptyBITxqQIATOyYT40CLvQW5l+PR9U1AE/uo/Jvm/DZqPID8tMM8l4T4cO8lwYFBNwNRY6bKDwwh
HDdt23R8/YwRcrJs+A1TEqXzkos9C3AmteYOlgNoitzfHsvzb1mShJ0hJgbjCXsX7HbHHBDdX5aH
vWFBDMLHwyaWPt8c9AqXfU9l9MRFJRb9+KbzhdwYXGcKCTXCKo3hM+nB17NC+mjM+D1ESsauXj0z
6YBATh/b4gkwVpc3uMk+w4rloZTYtPNlBZDKOcKMJirdjVrGFo+txyKK+y1JlZ6RwlJqvg/RVXQQ
lAO68N9U29SBFV2sRo/se94S5ux4ztimVt+A+yoFL/eU41kub4o/zAyDUSUWCnON2ZZSIZhgUW5a
NLlF/ARtEM+cWoZ030IAd4HrI1xbMwVHWQjx3YQud3AceXAaF+Ab5C6DILgPTn7p7HrHTKORS6DJ
XKJ90tgmNXpeXXMpBq1GZuMWSjfr/XR/UT2jPNTF+QawqmA2MoQTKWOxObBkBQmCjQFRInFw9d1q
amu2kyR2KFt4riTg604i6WjupcCEjWSzXOPj1Hdl+tByI+hQNjCNRqFYHS+FjxexMEjc2BGJCZkC
ZOIOu7w1gAuawHaq2bjCBwNWfpaA7iad7gpgotBXmzfX92RxzyNfq0xQJISsKii22i/hr5nfzp+E
utoeF5XKbkkcXSHTyVHmE0+m3/ZFhM8Z863b5bG2YnSjwTYYAtmEfX6grZPy8Mvm4DtpmYpX9mqC
4jQTFFYcA7bQ9zZPLtisSrWnKh57s9JPOZx+mouCxL2k0ePMW21E1T7TIau4NRlZuKMlEy1h+N/s
TLWIMIiJa0btx5Q6f0r7IoLLbvF0l5QXEDRVzuEBKaLin5HYn/X2LEp2hVYRwJKMXld5Pdmp7Ily
ORkaqhkCSpW6yDjqa+7sFTHhaAmJJg1HvsNc8xpzpCLUa3sFu9EPcjOkmgZmbUTfMhA6ArOXHrzL
LH/7tRItRmUoT6T0CJzV3KO/QSlzGxLvIcIBsh6OwrbfPhh/F4QNOylnDbjGYWtjkVxrhrFdF4yw
Dbffv0+yH1E68PufF3/KiDwfJWVUv/ZwaB4epIZAOczBBz/Gg/h+9pB9uxBG3heXgySUyeW9wlU1
3yIFj0TxSWenmuG7it4t27m6YbcFcXrV9udgJXTZo+hgIk5nfIB/OttSTZcKdOMY7IFvqX2ClNn2
vhG3+HD+OleterpqH6rHFPy5QP06jQP/ENRpz6Nzzb8TC8LAh0q5iruaVyb825j+x0ar/M1OOg1Z
Fm07tsEkrswZMrLJ9qNd+56ETndSWIk5k8YgnNNMjO1eAbCJKkblv9TfFVchwE03v+t53v2dQxlL
WUqt2fVlGH9jHTLyoP8cupbvdopfUKZKIA+geLHa5+Edgizb4Q6tMB62cqInfXqxqSHz33afK0cT
gkxb0RxtCagm34IQHGvVaMm1kimvswFlGbifzBEZLEEDOofyZ4erCkxSA08C/Ov6vvC4YZd4k2JT
A2dGYZZWAlbwcKcngYIa/SJyBIYPP/hg8ZhCD9SQOHVJYmWmmRUP1f2+CM8W3tyRyWjMPgTvvjYZ
vVljapk2ez1nJqSmrYNiLJrNBHZkONu9YyOQ2ZX6NfGJ0YIteqvkOdxjuEMG4lF7UIt7Ze5RLRpc
oj8h4wjVqtDVlbKvcA/ag340WvXuiwSoTmwGWpw6oC3AYwT/dFPu/yj/xmpLIySmponUZ1jB8YLR
XjrET3ka7CWNFbrXOCeJnvGsxcqYtF3q8j2rxK08PGIg8qAJflrfelCDrqR6oyUjYOp4J8H6wzac
SRj8Iuqyho/3MueLXthN304mCAmy6w9flfTXcLGUImyPNDhT1biHJq6bk6sHYLCpQkvIqJiIpIun
pLTrDCNhOqNRz3yYwoTsiqvx+DFPskXpo6NgABCxctHDeif6dlcZI2tR8fjNed+DqlshQBHCslne
Ct1ZfOMgs93sRKfjvFuWbZZrpueXdYq+tHhdPnICflz7gbP32mysRhoWvpzSBBkRkjv8BheJjqaT
vfinZSGDnLZukQrR0UxyqIOdLWP2gXPrdPVXHBdij5u1y9vfv5DRoQZgEkdWh7Yie3jyTwArxcFB
holfJS0cqafpUgEJLu+D6lmQRzHgUE64E9vjhkW4JBATHTq302kJyZI8mS3GOFoQOv7qRJJnGda2
eQb9txLbZinJVN6V3IuNyqmO1j/EsxvNTpLiNpzss/Q5hT4R8OaUeq9NT10qOXbgqVRs39JEXBgS
2CGJ9fmhmRrqltGG/LB6o/8gG9Od5zpxBSYXAdVy8vJLQRZKvR5Gn2IPLYSTOlRKpAkZsBXtBj3k
FN/ey70jj5gJmAzeoEGAMqXurQzNxwxVfBcpMQF9QL0Xp17v8PzGl5n+sfWAnhGlo/ZwTJie2iXH
+L+fSkmp1Z/W6OAQPNssmzPz4PBrr2JAiqQUXsLPyaUOCxlo2qohZwf/u6XVllYONuw2HvMN4m7g
hIJV3+ED5Hh44Io89PzUOOjgTqyzHFXoYjp7o7y2+mZONDBD9bUOJDeQbA6j83cuzNP8ndvKyUKZ
X8gd2f0TmbkYAo19VuYGqd/pcs/3So2NytX1GmaXRGyOgmn92NisJEk1AG/FQY7IbItfI9HmCyl5
+X5KGi76P/Fb5UbNV1FStY7pNIyNdBBxO0GV6+rCA0QdBJrlXv6D3hgNCaiMr5Tl1Sg2KKli4n/D
xI+RaCQOpziR57c18KWq6J6DPpr0SgGob4CRbwEx9z+CNZi+CW6bEEMQzctOzfG2abiVG18KkTiU
/v/Emsir/vn1lkV4HHaRRK2MLip8Uqlz1UUd3fxEDMM4kGGvaIKo5eGCuuKYVZEIiXRBiwI6V2yF
mOpqb/zgCV8kU52j/aFrg4Iq2LJDc0UfiA4nqeBTzEVnEVTtnHJoWinWEtqtoLipNKfu7AW+q1zf
DsEH9MZoVv85OKJoR3/QMYmBnmazdmjcVf9DrX7mJSvUqtlRnshclr1vFnSp35ogwUQ8b0KC1jxr
EXsx7OiheVEa/3l0jMxev5KeO8nFrITlGmsVl4yUNefEE2o709BVm6Lfv06gUVA5wGrXmEoI9G/v
ND/DVoID1y0xXLdAGkkqbRRIrcO/q+6zvm+/WmZlg+gXklT3XGAEd8LT7ErDXhlw2L4UqbSJT3+k
NqOv0JNVJE0dk53E0X9NrQSxOEnEN5eDUYoJF6XDt8XtjApPgzHkEzFn8Gi95750sa9bZem2Xwzz
GKIyIk52q/0OlUal0Cbg5eUENZsD0vulaitO45qRXt/6KABJgbhIc+AjjD8GogCyo3H2bNzm46u6
JeQv37tyL92/+Ip5FqR4L9ClQdf5kwPdg5kmPO2IoLBkG/EwNSTyRJZrBbLl5v/vb6mVJg3roODj
1jIaz/xqRFUq2zCzo/fVzj+uycGPwp9HQQk3zqPwXTzvYqmMFVbgOJL2OwSSYbRAqwhjTXY3IMpc
dXF04C0eB7AphjuREW9XIRyI4XUBOKVvNsZE+wzTmjqT7rFb+IPc/NVly816+8La/+yAUeEBLh04
o4rueuTqRA27a4bHLS+us2LIB6tQUWq9JUyM1vfcrWxdTAgCR3PcWjSgY1LE8X8dSVrD6+8iBeHV
Hox2mNUhPSsi1XDB2oI4JSTNB7lKgu0dNsWmBWa/qeto4ucBBLhBj2UgdGwcf0xG2OcsTqMeRhf3
NfxnHnSE+xR1fXtfQVCPAVa8G/jsxV13hMihz+p0jXP6bKscTlpsjBHA4V3TSOPIMJ3zhPeGM7zl
7gLFEaKXJn9TQmK5endO4mUshm1JTPiaXP4/VSiQXQpwLU27X8kKVX4MYSxao67cZOucX+OZfM12
BP8f3ksIPDsfvwl97FI7ItI210bEpcNyGkj9tSac9OtkEwQtohPRaFE1joxjG6E8/Pub9PY9ank1
5at7PwGwYLB7M+5NOZPfJgjI79PNVFp6Kkw04RgoR6JAcNe1ztygq2FmK7L1AtDweqUB9u5GPeMn
fDnLY53TDP+rq+QD/M+t1t8TxfKHPdd1ViBXbdIJ/gry6ITXvfOTF1VeWVS5FUOG5NkWuRKoTvq9
XOkQ2zggh47jjwui1cKhLbaDxsJA510qz2GTYTNf0qi78A2+DF/1lByTbQ3ZDXZhGqgF9irUf0rl
G+FmcnoX18DT5Utxwr0SehJeUyhdRHocifYnr7wwj4Bi9+6ZD4eDBLsbN44Ow0jI94CyPgRsLUk3
BY9JH01WA7b7BN5PCraDGoi5TISYbZ1xpGo60f9rrU1AvQh7WVfJrLev9f1YwhA1PkGiBWfh2uSz
kbRHeWTqB5x4DhZkgU/N51CXUpvAe9QGnHziI6Gj4gNIVzbKwhdofpM0LrPjQAfTTqzMlLPB/oVa
tmIeqGl4lIhZKFX3JK93X267Yp9CMrvYgU56wGYWjS8KPS2pSLSIzIcQ3uM1KsJz0J1CYV3YKybJ
1t2mAfVrnE9PGZGvaw+Rd5dDSGEy/lwKsWLJ4vjPp/jJBCOQKTga3Q3+/5n2HfdoBanCiwFK/HiE
htB38M8qf2Dqojf0PiSIujFrXfOwxVhPx0JdJbbUcMcN+r0RUWxs+LpGeNionJMhRvZUIDapYOqC
xbHdbDRhEYf2BD6KsuzURA1XuF+aQfLYieOP7q9nsLeGN65VMqPdwnAEs8BsrQz0b635NhOEgzN3
AZI0JgBDu/Yz6SW8FhOLhs0SDcKfZIJ/XuThQ6bz2ZU0TPtXUg5cIj5RsAqlxbV3vh/88N3ddnun
zMMDP4QVi+jPG40DLjL7DmUd8dKTXV9W7klC3RXteyG7APmiL245EhmntS/+rD1Du9mbIhiskSMG
fnTSHKINjrd9Son/vdWDN+r9rBZZrq1qIm9rJmMWXBGYBu5Kz3CM5D1iM9CGi44Bi3zuXih5Aejt
gR+NuvHTBZO0K3ARp1siaPV6nBjdm3mTLKpnX06noK8FyCRO3rzTdg5Q1T/bmJEossHasDHYGbNZ
swb1wsyeJFdI+QqRZ3IoBQhyVtKy1lcaBmmsqYxwmpbHhQCLAs8hyuV9/mVfjJj+37NlQen18IVp
y1bzgH3DUYBCwnt9BJPk0LLn0gDXA2zePLt+e2RP4z/xBfAe5+yrwaoGWi77o24aHWJiysKO1rwz
4mc7accVzFFLdVdCsF3f93soZ0lkUGD6Widr6S0p3CLMGvNeR2LPeoQHIz1XgZxW3lBUmTi5jyTc
IXekY1FPnoHcdHdHJxuIISduOG0aHZXgjacdzkR52SKM6tC2I1iDH5RAQCHfmf+Q3UdE/zT176Uj
yADAXNX6o/JCmigN5qx495stZ7mrazUtqklhxpwxdUQKKSZvAFQQniaHs5fRIYrEUySYmJ62Jo07
U9AS9a2dcHESgzlq0yhMbT++QOKw+FT5nqwSZ/J0GuwSseTNopi4nJkF+qFadFiO0OS+/SIM6t/Y
EwqcLRBPBStQ7S5BkWB+6e602nnZjL/L97+Fe0VecBX5IfiIS6Ruw2lOjP0O95i76mT7I89P47BF
Dg7Wi9IclN1ZZdPPtD5aew2c00/TlptGXPyggArxcWn7mWLChWT+X10tyimbO8ZKGoavg7OGACjl
paxkCsAhbD49Hhwn/5FEYApXT8GjRqy77LkAsg0CsLW2HLjqZkjmbHnaPKENWRteMplLuNtKTSNg
yMkxzmrPDbFyFGplIEejB+FSoHkO0lNay8/PmJq9beepzUYETVfGwWsOMuMk8KeNv4zJol4ZRV9v
u9bYpG/aMvoyemHEYHB3Ia+eRaX+vcbbpowx3xZWmp0/xUvr4ksipIn6oMbohSyJBx5ijpBoxfs/
BFMKO1zZi137NnJQ63MPKGp1DFhJf6dtk/1JaCi1qyBePXJyXom4UANCcuJzwIJd3etoSVR1z+VP
q21mceyjd4IYC3IcT/vuz+9fC6O/gZGRR8U+7AJIWXbPH7yfpmXnI8IwbWNTS4HW0go+O+LCgKeG
3hg4KaYaZxpcyVENIVpgaZxBih6R/q1r5exORrNSeeeN+czvtLLqMhevg/qK0rVasCWCpE7+2G/7
F5S41HhpLsmMBLNwYjqiQOr+CwZregXTxgJkU8tlz7xgVq9hNdZ7o07ImuamSR6EH3eem9XYuaP6
RA3f+mMHqDo9WrYYTXyk437sHmbu96kGiXpmCt6qtvgAWanP2SV/kE4okAp0IOK+frr+USg4Mpua
3mXXPae4kY3LN2lJc2up20aVBipsI0tiamdGq2sFuTlix1Gcj6YXvEO2vOw/osfmsg1l9nGS1m41
Z1vrUxGssh8HH7koK7/a/PMb7M/uIFgFRdghfwAqZuOIjqdIiNzElTY9/H+GjnnTd/vIwSJtfIy4
D0QNE33WpxGxvmF97DGECWM+TmTLlZiLgK7ZXXcnmHniUhTydtzr0Gs8gM8PmChLLpZSkDzXJ06t
XPla9C2t0h4/5cpJf4YJLl5eZnH/PuZIAPPcMOtEYqRnpbGF5DM4MvbrcnPNf1vhRHsG9Zl+6Xe3
zUb2o7An4Ob61SXGZ5yIJx3UzSgJ8BPZWLQqIdSMQKB8TkRZ7X2I/GnRSBWuyaxJl1D8ousN4cLx
xm5kfCCcYas3qclWMSF6t7BR1dj4jBri00ftSJvlvGTDW0fTQUDB+Ha8/37Hxu+w9+QzJNsjNiDu
sNeNlAjBR2gdZQkZuieK9qWmcKbqnVHhs3JNh5Jlckq0DRoBq8CooPMWUOJROmO9Hl1egMlBGUdE
e4HpdB3ivBVSQ8G3Ju2pR5rGFcGS4m76lx71Fb7Gbg7go/UEyvYMmy2ek/OUnMwShDszCqQMjjvc
ZUCfpNrXKSAH7G0MkVoInW+yj7HR64f99bQ2G6/RRr6vkea5YuwstW0hQ/IF45yUr+cGFAyaUns9
e4L7h5OziPxes6OBbt6M7+gr2AP+iI2kD7fTOei2Oae+FfYFpRNV59/T++qae/nGFpk4E/AiA1Ad
ZLvKHHjxK1TbAkDFSaNIMDXvacna5vR8eAxjeKqmcuAIhH3PkJgpWJqnhJh5Ico8Axx8CmoI+Vve
Pf3y51aQcE2M4FJgCo6rOqheIjN+iVgKMHr3sjqJEfruL5TQtlQnWWvVA/WnqHuXpjfJHCVdlzQn
6Dj4JVt5GEgyxt+//SWSx5yYZvyq2SvdSBKrJi+dOaCJrfSwvB2VWLdCZut7hgkkkhDH/ZlD28we
Y/ddpGnspqggqsZAzbsrHNUocdiuj1u4p86ZwFy+EXFUBxmHU1TpGrwo7GeGVXamDPPihnJP4yWv
saXoU58lygnNcZ9Qo+qBg3jI9T3L49qx4SWO1FrAlfs/N2TUJ8WTLZPMlidEQ42t3E2+ZdaAL0JA
ztr0rclHkpiTG/2tu4Hgk0M+CUiygKIll8khJYAVlD3Y9XAWXnYhpbVYkR9JlQEi8ZOkTnfGzydV
mjKvChSgksonvCXwse6BuQkjUSCQMJMmgYONygvg/Cepry+LyK3Qj/VZvlnydw9quj8rKRpC+EL1
7i7RObS5pmHRz5ZT2ZlGZeOWC1abKNOf8bx7ibrJkKVK6Kk9vfm6IeaqXn426WFF5/mDjs+7ClLF
6M3W+kuab8JuYQIYJgfUwv+msFo/V1TwnPUtql/oEYFFt1nzwosevMFor6DUO6Tq86zB+RaCPRbo
F94nOvKJElTShXDSx4vt+Xnghg3cr5OkJktiWR5pjhsbk2DqwhkunUMWXgzVd/HzwSI6Ic4zH534
/bLoL1sxtE4HXUZqoaFz4u3YkCg3HFhKSFy8l3ok+wmtYJjV+uyfvxsjA/p1NOaWwgP7CAHFn73H
0QHftlbsmPM/XNwrh0PspZLhTTpxCg2oUcwQDFfGxlivSV7xb8k/4qBZiKqOryjmelMVn5PSn5Mh
1YAP4THWPiF/K3vApmSmiztAcWSg8wj+7BTWSrRSXfddEoxKQFqurZdBMTHFbsyGjjzey4kIfU+r
3+MjoXMs35zW6q1YyeLwwjpvgiYRUvYQIbu1b/gXM5s7rHKpquzhZXtb1GffD7IwQfpbxV0yzOgL
Rh6B9fMf8YeZEpExvuNumdmCq2b3/LYeqdKhpZPzwnxrvzJ3xQbfoJyveU+f6i86hh/jgqz+I74M
eL5UiI+Bf1xJ1AjvCrbDN+fszCNj31lxW0/C09qoJiBlBCy1vWuLR0M2Fcs9JNWRoW8AeF/npuuu
fxYgeyV9KSetP+gwpxzRc/13lnzQeZ/A10t1l5lLaHBTLmQ8uXvqdHsl+732eyBx4UxV/w9QHwJI
THwOmt+D9j4CYGrONpDX+sXFL2+kQghmCjwwc6//dlB3OS1VH+P1u6ARl9IFTnRdqD/YdHFyNY2w
mXnB/jnJ8p3VSWVelc2FMRTC65jeosTZ8h+niTjruqg3oKbMjlXnmvrs+9UvtpYdgnp7/gvyx3lg
aogSjJ6Y/UJuoZr30TeHlIUHr5Qg74iGuxG0SY7/fuGasTaIB1zjus4iqg4lwIMofI1QXGRsj4ky
jXmeqi8JDBQfUQH8jqhPEiPq2dLlqFbCS+g20y2/2Z1sEI0+SeFT2Yxxnie1u2NJ+pnjyuwKXfw0
WOrnjSrdiXDjq90UMjuqlMt/GWuYXRkrqPjKDb8vc7XtUexN+d/fY4b5UX1RC5E4b666V8BF8HmI
hTpa5886Oby3DJgeZBxGPEhseCQVRMn1b5YpnnMcxpm05DOPGt9sqZMtYmHl72IrOxBD3Cojgwyd
UEM3ZS9BSXZFyN+UEl4iyOXaUZsnMSO4Xwxmtdy2P4T+mDQtflQfdIOimAtvGfG6dO7LHQvgfkz2
rqCAm5NKYm0O5+kdEcjwSjl2j9wjL3LxQ8+9TgoPngCPwN9H6JuNbaWf/a5pf4iOgTazypBLh8et
uZ7uWNAJ4S/mZAgfK4IrR2q8zIPnoa/ZpF57WoQ0JcqkXQrcsADJM/AjkkDJ9EEE4ntMBjYYf6y4
vVEaL0xprenRVTp9YtZXt2h5YTagYsKEHbfiZdUh9zYpKyu8xYb/EE3coyuaTXj8Ok/G1ELtr+iD
u+qaQggAbZnxJpAlL6ss5bVJye08XoNhHTWPOHvl5/kvg9Vci9jKBvVR5+BOELYwdXE+wVQKKWXV
I62NAqzU1a/+Umkeei5UXlGdCFIHOq9c8HbLrHECF9vR2VPvxQFhZm9p5K6mymytXmGTywByjBHv
b8dOme09lh6zrDFgC7QZm8+iNwS0tIn0aPdhQ5SO4TEdjayF3sTngV58i4qGMXF+bS+qk1QwxWmD
ldyvSBAdbTpDcqS6iXz9wiNCb3+AGJe5hoHweQaZ7k5y/TNBuT5dOtyuLPVlEK3etu/ZDmgiVpJA
jOBZgNXfMJOsopoU3Y98soSIw/GdAamP1HIzZomXgp4W+/h+4RiVVCWl0QpOdeP/YeFIuIhRs11t
E245W63/vkBh2geCH4pHdVXWv/KyMIIx3mgb6IFgtRCi0fx1NzRRFZDsp77CCgaEm69n2eXlcSBp
/8Pt/ir++jcz6NrRtOJASYyNIw8EExyg3mrebQ7BbPJzCjL/5CI+eHd6MOh1lORg9YbW9LomLzc0
XZSb3enY3J1hEhO55NVyF7sCnx/Jm5iqIPbKVfJIaUNv/fFAQ1eL0mElSlapPcpFyiGDlUzerTTM
Xwe6R5QSbpPeGjuFRXJmUgF5cpSa5Wh+Rp5ooy4ipJlgFc+/wMt6VqcEs0vTZIFnKgbqE2UaMA6f
28uAc9CYUk1WkNHT6pmOOwfy370HWer+lix9y86uLp/6SG1KsZ1cBBit4BqejfDaOodAqEFRBPIJ
gzkS/KCB6w22hJlymku8GpPKZifkHqnG/nJlSOJagtZiC5Kv+925MQoe9NUD8rrh7pYnIQHUHvb8
FQFnCh5G8XGsAt88K4pXB92tyNB23HS7Rzl2nSVKSkg+fLOw/KQxtxddWc1yK7c5/1O8VPZ/taNl
X6dBNS9pC7Svl7U972X9zdXwynECZNDrCTotQhegbxu4incFv/rXOf32JdW0DHSTjtpJW5Vcf9eA
vSZBIhmQZw4fwQ0vAzC2EytFJ0UEup7VfDM3H7MUbtQ5ghNlEcXwe3VYJW+CY0T0sz07feGNRKpf
3eswVGQn3Y6YytKiOHfZvoQLZdnOVWBCJjrNxYj95TTalz80tlPvNg9wDN8AlDJEao+LAEfzg/MG
eNWepzqQSgWaTdXTRFxDVhhJLvTW+RDRBmJuQpe1+PgjtMkjQfuGg7O0TEgXocJFcOx7yg9FVBOz
T3/envf2Zfhm/rwcwJwUWPJxv2GmedUtbRzMfdunv4cOO4waZY0/f5+a5bnYi497f4CTqs4q7gBG
BIae94UszqiJuuSSKcc9UsPnf/DgSv9edEEJ5EihNaH+SSc7ApNAzbG5AfxZ6zL9wTXix7ZV2+JJ
uJ7HHXDSSCrXq47aEBaHy8fpoFtDwSgQNUuiIcSVwKlWjViXzBhbD4ZWBKU0qGBLlj0b/Gy+mFVA
2hliC9UbdB7Vfp3ZBleKBJeMgQanHe30MnhQ1vStDTcFLav1Xe5usdSesTMBKPgWLfGcNtP1l6jC
/i1ySvj+C92Q08jmErJkTHCudfm9rABZYi9m5Tgqn2HsAJhOlcUYTM5p1Ptco36Oa6CBCxwEqUBt
hvJK9tKLIxCBufpMLIRvgWpKzxNgxN+axAHrMusbDzEEGPlA1C3il5dJYjTqDr4gY2aL+P/BzgdO
Q3jVuSWKQC85FmwBCwXvpHV1o62533F/Ux1ozwvmHMnJuMx140tQBW2plTCffW/WC6LctpEsGS0X
YxTsFqncM4x9n1hs4AyM4XnARdECEFP+gMson3TEzc0YSgMPCoj8y6C0xiv4eeXEsKEazHTm4EaM
VyHkh8WFSZKwX8tG0/OuxQ4j3mNYZUqQ98pJVjuxjRdHbLPp7KUuEzRTG6c2usVoFUINjHO5U+u0
jL/7czOFJuP/PnOhCtXnEfNZYf5so2wKpYtK+U4d9iHTs67Ujoig7EAxIDEs6aYAzw83+QZW7kMk
fOj1Qx+lzp3nLjyGzWnJbn06NYA/lgSq/bRVtOvWdCkYbj9BE2/34TNwPzHlbDc6BnHyAonq2g1n
9bmyRtsZXWI7nw3/2v8UFK+UhT2/JAtQmp5e9mgJk0awlGS6e0LzX+u0OJoaO6BrM3szsvSNmwzQ
3ukQWb4bIRMMFLKyA6NY1JJkVmuvbt+e6Te5qTbH69bpwutD9tlimjJpyq5Ut491R/s4/79hb98h
yhJJRwbo3ZDkFd9svefFl22T2WFf9iXALSGCHtN4uPgM5maUpwh+yTwBD9kLGJfX0Kd2M4+fs/CR
BYPj2MEPCqD/TuaJ7pFpdJAUcAvWT3JTc7aSqqCistURVy3jTK4PjZkJtktTU+fvxXys2h8eoxzs
DlyPpnWsVHsB2VxOsq3TYJ239b+HZs0K3H/oXoTy8bwKh6kwZMQFj+R9HxyL6+MREpBDH/KvFPJy
7A6EVS8ufKx6awdQ9MmQFEpaslvnR0V7Jz3HUlQgr525y4TVdoA5+k4Ybr97H2hLMIIH4zK7AS/j
JSoeUu9OKkDy5CY+2dnP1qq60ycDKuJOQXXDg/2p+d1Dn82ENxigfC+JD1iYo87ohgd7bmq/tB+w
8ydItLPzhrJmMa+W+epc8aB30MepGN41y0hAfwBk7EVgcnc/NfgSX7c11LpgR6qBUZ34mhUyB2sR
w7FOnqzomdFdSSI/0W39l3j9hGNHv04mdbNdcmjMN1xpoH4iwKG/lsmOTeyL4IOa4YXcQbmgzRy7
5KEm1h4QZ6QNTj/s5bheHIXkM7Hy+waNUogJCaMdfh80mAzJYuU6DgQWaqv5c2asZHk6FONmGsnM
zuvoH08eheybksAwFRBOHHfpPQLGlWrlvrOkB8Fj90aNe2R6Kts+QEESbM5zsRLrXEECudhXPSc8
IP3tMHdwNJlB8G1u9vShiY2kfUOo9MMh7hlpkuPM78z1dDKoRRV3jPm0o+UftUdslVlz8Zvsr3H5
JSYyUzp4VL8OYXJQzjKCDMRqPZhmsQiKsK7ZaK3J4dZkIl0evOorKAlovDxDlACus8nn3HVXIlyI
A9XVxx2aA+kjsewsj2nbJHSUWuwf9JKFq4M/C/y1ZUrv8+TuV69bFkHisURE4eBwd6y/vWMuQm3b
sxQSAKtOSWu6WYA71O0OdltDovNys0AbfG7cR0zrKhAw9lhuJ2LWejPrn2s7WphnLAyBW6/TFFSw
GiEJJZneBbbB1SLEAiIIF6D5gt2sc1n06ds/4iHHYNcLk0UqDcEHSaj04BbRiN8q5Q6CTqXnm5hF
e7CVEruv6N736bzglvr3qxazP6hf0qSDzF5CvACWtbFUY1H+fIQr5nqIijBNvnhfLvwfFKXDaHvb
TX3Vl93cykXKlLA+9rpq6+fiHNRJhfTCUNTk9w7vlEJzlu1P5Nld6bFbdM5Td2pORAtIXRhOsQg0
xdSWK6nI8xmzjzSxJutLvYfzdVSTVvZMpAByAz/An5FhJAsbzXP/p5MoxgDv6tmhN61bsj9fE/18
2jghvuY/ukbhyvRgwHRA8EOr+LTiLrhq3iJuoHWbea534MUFuKWs9qJxtXq8T1bAhU/9epOPI08L
cyUFyaMdRGpRgMVFQSf91T77HyAWGti3ZWg9Ftra2BOtgYQ88XxDnBdk1tv7mT59V2xMBp/xix3G
f8TWDtvsltMNvk6HYvtWM0HKR4D5vkUp8mbkCsjaLHbiFshOPeWPVuvWbGCbzV5D/CHKOGmLZrsQ
rQDx7ZNXXUfkf7ZgmVMgMGx5IDN4iW+fpyKD0p5BgiRvOh9o73GlJKg41gQOM8cMdHCp4bF8OCgS
/VFVikdwFiz8fapvrN+SdthqsllG/PcCKkODRkLP+GXm73SMrCQVib+olp0SO8oEzsbPKdsTKVos
jY1yjaf4AKvtZyVkbQUYie6qBMmAV2LOH1PGGcT5vzFoCzV4nJR2ZO8mBlN/y28kfJn+7g727S5z
qpFSF7Q1TExRWOZCQSKcx1AmYN1YLwIDpYoUzRgw8+wCwUVZ5j0EJPknXxknr+kL50swqcgr3rwS
vog9gQdID+rD1Tvr68wi/UBQsC1yNyAUn/DLDjt6otoNUNG8NV4mULUb46u1nUo4Tv+AJxgA4Gu+
JBF7emfm+xl6Fd1vhExQre1WnU3etCdIuJghx+0OqXM44cFtdYtzwDmRCeOlNP4XOvaUF22pTbZP
VrAaG5FPZxk4VRS7D8FqVLYYUMoNx+Zfbrp4TTFB84t6Cr7KANKQrFfPyMN5lfUPNqe2Id/g705D
AY/99tNae2D0A4TV9SdoIqhSNLBtXZZTN8D9svxs5dy50JV9WUtEs6o5XdDfXVVrSp82Fi67GHmR
MvWmSmoKxOFbXo0ZEGahwRIFlbRLz8ZwvD1aeOavyQSb3cKgQKELJ0+3Tm347cO8hfBqL8+T37NF
1z4UpLd6VjmbdOOZn+vN6LcMwJYkkl1gjXdwNY9pSAcA5c8dkGJdiB1PJNgS8Vz/faFJGe7XXJw5
OEPN+91ZyvSQXOjYmBBazxXT2HNhuvcxeCE0QMOmt3Bb+uvAZtd27QwoQcL3VPGUFJGd42/KdqVO
OhNhFz7wtxan4z8XetLOPrac+BHp0hzCLC5z4PZoTREAGeckcVDhgWbmvJX0TO6/LiMjB32yE8ue
rEelKtgCJgu+cgTlPWneA7WgM45kO/Z7Bp1q7LZVFS9jQa1u2VgZvGc7nXZPF4Wt9LCYZEGiwbl+
rjwx+JRL/HVerozFMQfSzsAf4CGpVabQsFYlv5KRy7CfaX/8gD2TAAlIzMMZXGp1DdHSB5crbnjZ
Bk7KBxWN0AMP1faY/yGLldoMu/TjjZlPuOEuUrf+V4mgYlHy6NrGwD6PBUqSskfiRQIuS3oOx4wJ
4Zwu3Pzkn6EzbK0wOfD9bCIbctpuodbReYd2ipesME3FKySrx+tDDy98Kv+fkbNUUzYq8vu/X3zf
xbxVR4EesPmQlD+/lK687VaAWjWhqK5Yfb6DhThdBiR4XpVBz/YPyiVsOS032U7FYTMDcSPDypf2
vYl70bSsGE1PM+4SMabmOwE7Kn1vcdNampLExhUi/WgAawB8oAWqWawqC6Iduai137HGCyqwQ2xF
Yjp49s8hRn5INh5ZFg2gEG89iltAV6ojjZ6X9p5CwoFhzb04bFy19ZbHl0Zs/dPRksc+UfsYHQNC
j1X9mtAjqCMLhTjPv9uDZXa3i+mixYxIC2Kw1yN50P3ppDE5Cg5q8WL9SGZz4qzoTDy06uXjuDao
tbhNbgzD42E+NvEH6lteur3qT43WeQjSuvMdkNJvq+DvzWtitBLHrTgzTEBjVXc0qdbK9VK7ISCS
lF9UkhcOwBU/oZ2zRy4LZiwCTG96pTcX0+28+Pc1g407uiFWLOUASTre9qJD4C98sftyyakIp+lb
2eB+b8E0YBZQzTTC4ZKf+OlEZhusRgZH3OzCbTXv/ZOGn8jvG9KvCQKuT4y5pwfDICTsReWjIzB/
lcKTBPiDIxKfBic+M0pLpAUsAgyD7WaK8G6w9oNP49y0mnd0ePaud5beX2Wx0rndXIXzyrrvjEKq
UM7iDhkVZu/DculPnLoOlBkENL4+F/7elsV/8FcRac4co969x9VoZu3aLCbAYysyqg4OM/6ZJvC2
TlaQ24TTCWI7tPoJzNpXHTS43xiQ/tT9KCVmJsb64R16bOvPfMnCH0pEz6pb4rVM2EhiKZZWyTnt
WlQoRRDR/ScSzYaw3Xx1CKkESFFwTiW3JxfIx55qa4ZQQKUCrCHPFzJIv/jr2mrtxbVrG8gvFhqS
NyY39qvhqXvVWu0jBB+O8eYEuPm4HA/bctyv7p9rWtZnS7C15nj6m1zbhLYSbs3M5Nox6aO0Uv5u
p9k3CUg7xtgE9SrxGgbIFqtTMb4aXXiENi0EGUehRoafi0wcWYRz9HqpX5/cgn+NhS75PCVWvHqo
Zl0BOxxUy7vUGBLoaDIsxy05JV19JRc5VL2LQzeRuoWpL0+YKFKP6LSVzhmiedlNotbusSE3zcCO
T1gJBVZyDjn3RxrW3kIEFFGGh5yjhCxNLsYzhKmLnRi2+4ZjZu1i7DjtirXW9eNiwmHPR9PWIsgJ
TooSXaDpv/+bnHDG9bHl9B0xAR/5QSK/tjghfnhXt0C921/b2z4EZWq5sJDE1ZSbH104/Blf5vt5
7sUlJ6jkTj3UJ2RJCU9FbDyTHfEcOEIvZJ2XupiiXKs6EdxUsTQu0eRfl9Z0cI7FAoR4Kk8l09tC
cdihUgA+JiVYSvDZ6TQxPGV3vGhZt1O/0qaMz/7V0eMZCTB1iaWunef6j7CLx3bFOtVKMllneH1W
BjEknuLLjdw2Ql7dMcbrlEU3gj8P9FdxVFYxtRFxKAUl9lnKWni53maq5a23bM02kSVenNDYDE4s
6e7rtdl1GvfMzfVW83QmJmqY/Usva2X+wvuBfHKUWV/PljXZs+WNpLEnFuWnSPc/zFKJY3SJK6IT
tH+45AhigHiXSI7MPTtu8RK6GwvfFhiW5Xgn5AQVtQYthB8LHWjF9NslOlKb2JS/QvEVGKuwDHLe
uvihvn1xfTy+RZVxNxjZkfUOI3nHLSoKQoYsUhMUhVAwcIdy9eP8WJvYSb0BugrypGp7qdyTUQwC
NOJ40dTkQ5igodfElYPvdUDZ1HYwuZqFiao+KR/JT6zGsaVcyD/o3mKZSzaJi+IcNszfJ0kTHlr3
Z2YY/oreQ9Dx9QlG5kCKQvBeS50oqVUB/Xavh46mR0gWHFNEBJCVNy1OGNpQRLHaL1xDnsKyONaz
Q60tZ9o2n5EwEofKKedApIVZLDzaYFm9RQuhtuSCeKPJzzOusEfNN4kE7JrGGJ58Md7nxvBCg/kc
L/ZRAdHv04gW1Vx7bJEM1rUI3iLY07HCWFZZULuyxURgAVer8mLunFS1aL0A2y8HK+kSSBY+gvgP
yrgz5WHYgPkJVbq5ILlmLxzC6Z0PyPby/DSUmf6q2K27H7SVtmLhYt8OeDPMLHf40wSl7kfzfXPi
xtFnchX8m4ddLUGV3uaOrBzA8SA0dqlDHFelpcmEFFwr8GAtFbU/8yxfU0milvKBSm6Lcx5dplRd
qNOjLu8uKvqhwpdzTQz5uMtKljmRzUQfAV8x9n1V4emdpubmlqUFSvEeNxwx7QgLktjE1eIW9hIY
PLI9OXJc3xJLzEavMj+j/flPtbE0qydMRSpYkwaH8m1Jlpb8+U+JY+jfoO9VlUSngw8IFwCfLWPe
m7rlXlB1LDKTi9xKAdDAwpWHNWHjkvBYhS466yd5s/YTWzNCONBzd+ecrFQ5ke13+n6YPLxz0wIe
ThJJU9PN3c12bz559UI/CUbUyx6yAEZrlkkg9SeyoyAnzCHHyDlawktEH08K2aj3FfytNgehv1Y3
2JR6Z6Z83UW9DKRRErFtRWIv6BvevpDY6KRvciBCjoCwAE4fMcyi3SfaMPWbGJFzX9FqfYGI+ms0
er8mI9rh6TlZNjEXiNw/4k0yNXvF/1UQhpI/ILivmwhvtc3mD1jOu1qP2XPI7bHbvhELST2jkq3q
10go/rDtEgJIxsDD9OCJoJ81sy3dqgrksn3aH7RFSUnlLBqxBYIkxMBApEQfyc03abWso3hw0cjG
kqTCsuMXx6fxbQDYHLmJ7pmJX1lYeGrdtHn7H1j36sBtEK/UXcZMEzXIhME/o6nEVIf2p6VuWiEm
yPAc70O/tOkGJ/QUPmvkTXopSeCk9fcUCMfVCogiNso3hd9Qf0B3oF2/toVAgBrzDPrMq6Bn3YRh
V36PsOjuTbjfG0mA1qT3m1JyeO4zH/mzvSA4hNUsvPnOQ9Bdy4h6AdlGIc1EZvfdhOUbLAjf/ujq
U9pWkSiSJz3TAryOs8pZ95g3tSDPUXh/0pPzZeuc6RXwPK2D/glDHyvyr/HSj0ssyCnTD+BofS4A
vKPy7nswERo/wuLzlXJWAIA1X9QJ8lfDt10wDWt85TqfJ3+/nTxdGvZpEXV2QfVN+9JlMbCyqDEN
+5RxktGcbIlCLDNGEYBBbmTJE7qQTsbFuIIDix/qbNU/ppI34aCilaoqrsByMUCSFOkSuAJ9QDa/
V9vGFk5crbB31N+4knOexyUJZMrrHdbiwe6fP5l0IQuGLm3Pr9tSjNFoGUm7tGB3O+QSPuwIJBQU
c1ofwTenVjakSQZYfFohEEFdX9yu0nbWPuT5Xu9OaTBRvvT11Lk3V810iT5OCYM5DV3/jeNWEhfw
mB2UCMO4VqFZfhCm41ZVBNJe1T3ndrsAqOuwGiw6NMkQf2pj8xXPtZc3fyhqLjoAbxPXwYgC/cGL
I7ibeFTb8XvX1YnnAQ+j+zp07ev9YvYxd3ytaIhADp3M4hTMocn3Ij8LysB5egIlQOILkvFhm+R6
g+/PFgjY3ta+Knd2cxKhD84h2K1G5dg4hf4JlxqOx6He+W818Y4Ml7kl31ai3KR/8+SUZPZ5zVZY
I0TBKKhXywlDEa1iOQluQPjs2OgZcjGIrbrJDz9Q5FYgms28ovLyCyRyw95JqRzKOUn/cfHMAy5z
WL9KgQuxK4bWiFGT2T5oJPLZeUtmTdN+n/9jAV8MX9HGGDQ/tFPmNsgMXaLk72LYxktcZmNf2Dhf
2ZyE04xJniJiFkh2eZnRic0PQB2ZUO/OGp6EB8p1pNjysl6dLCkeP7ZhFwuzC5qoxVz7NmtO3Z0a
8VgNSDInCuXl+k9kCfRxWSS/RKdKvFNDH/FRB8RHieGysQrsUVefCR0594OouN8Wd/cB/6drnVCI
HY3/PN2ym/4AfShron9nFxpoWOkn/aNasANzXqU9nCX95x5XgCXRJuJq0+Ca+WhiTzqbyRvYBDDJ
si0slEho2jEqQ88x84kzoC7fLIDfRUGhMVErb2S3KUC75MgXm2AnoDCnOhzt1qqUj3MNYW0+Yqd0
RgYe7GvPGFsTGhJhNOUHzRm70BSGc4yYV9Z2T8kGgDWxbS/rxWfCQQfOyiUjhhPKHz2rJzBKIp6T
pMsuACaavjkK7VoaM9Epn2A4A9ZG0U1eZhlWNqcukuTrspS9kvNNgTVxApjJL8cFZ3u6KstrOPWm
lO+5S3+3BXSvX6O6nVO9jLFkbkPIZzzKOTcUxc7g1oe0EpSMiNJJcvwnISJU3mjK2eNTtiNcPXKH
HPE1sGmgdc5WCCZSw3POKcrZHfOxCxqKlC4oCbSsPWBUKyzbrSv4IF3AIh/SxmGKMVoebYXSuICK
qIvA9pBb8inw/li5EbLo3aQJNyVYXcMnNnp44q++ByCDMkkDoKAg4iREMJgEFKrSSxgADYDyNMsV
Mzaap7uc6CxSPrKf9TRfwPaJhxlf5AOnuwb5qNb67GaUZrdFnvxxXkmNb2L2IydWT7ZF6EZA6TSi
tUucIFdmsqmYZJuoEgwaZaRjEN5lw09WIvgaT9r/piBoQK3dWpR1NwhLTtH2TcAsQk6a+i5eBJPY
2pM6upqQvXokPFlS4iX6d7YawG+0uk1O9j0XKOpnCxdu9GuNr4m1IarZU8n8MfmnjC0HyXE3Rw+4
A1Ia68yRoyKn46QORJYM+KgiwBoJXmIstfhVJecybPy0uAxzMq8M6baI4Tl/olA/1xVJwxlfp2yI
OuLd17Re0z/e6AuBmQiv85YGWGUoOTOSjfvvZ0IEus6Hg/lffzhHcXoU9j1QPZ1uyXGzcFZeVqfN
gaYmbSV3h91Af5tS6FmKMR8C39Q/NYtlKOb6X3SkjVeNCJEl00JKWTI8NpR2wDKanT5fW9/TV12d
K44DeYr5ziQc+wfZwo6oDOHLQ9xs46Z21bWPx4kKrbsCXWandisXfG1gt//ekXI5FZEh1mrqaiAx
faNHCqVVdMU8DDruvpRxf//G0MJrHoU0zExo4h2w8axI1uBdRMxhooQ1QG4kNV6TyI7BkqiAW9SX
g5NlonDBVAgEL8IXkeTsona6WSADnFRVa24RkUXKb9nYikbYj3To7DxRVeWoEvMQN7idInRzAv5k
CoRdemkO5I24nHi2bd4Mgo+1Wkp2PQdoM98DyTs7xQVBi+1X/JGklU6eRnfelOiTXLG3sSMYjDfP
x/LBKSFk0WvZMUp6d/7ALJgXojrpybGJEDmWZl3nxCSy/Em63eYdzOkZP1NI9yydTJat7KffdTBi
FoIujcOOjjyxVfKrS773ex4Rw2Xb+So3+lH3izqbKuTxiKbcbQjuX6rWvT4k14qH5QBwfHL1pYxE
9UNN8pkVeEk+KhPv9n8xMSeAepOMyIMt+8WGuxIWmDua4INGL5VfzNYWssEjGpI3ZdffXl2gT5B4
T9fnPLBLuQCSMJiy8vSMmZ4DAxTOH8wj3pXUC0XeTfamOeRKwWp5cwuN44mM2CW3dvi/vhMyDIHU
Lghnx9iUqaBv06OB1XFtNoVSz5mjbxjMkGolDBFK/lMyc1Fh49wQHGtrM7FsUJVfahPA9qpshuz2
YUWmyQnEOJAg9E/YFNa8gnQ2D07l6NgMM9l7CU88KMIus1n4BRaguuqCg9mwCAk8GjR5b73F00ge
DN4HJEDtY982qjn52hXc5vXaeimdlqXyC3zhj0khN3GQjWn0i5f7OLw+K99GWcr79XnhwxPEJ2NJ
YvyQX4+vqM/eiwkdCY1vnHI2YieAQgrq/5v1wcYvPIW1aGXMvlDNNNWJATuW/uZXBks/6Fu3ROjZ
jJj2pI/b6CywKnmGYZcSKmEfWuhs+VQsYCGPULAes0kCcGz9CMt1bj3D0AipHSHFTV+9+kH6PZW8
2ZJ9TTf3PEzQVRtv4w3UcuRzTW54qdKqzrfRdb7pnVxKYjvlG2Fge8DHZO1M424DohC96WgQumLz
1UGPa65H62LNsDG0N5S52ZVDciYR9vpqL1i2SH4yBqUPo9hWlz7CUE8vN90fKnhq/Eg+QBZY2eD1
q/eqs/h/QutJJ6AOrwHAEif43drp/+OWDewFMSAx/yTj6cxqdwFBN8lauDJC9708W9fISFNR0Mir
TX6ssOIWzx7h+Ghl4mlJbQVJKovQ0EXDWKD2ZiCd4Iy8nPpTqNUSOTTyvEDVPlsV0BRu3iym6+wR
H5nTvj7d/uSloVMtWfJxk01XrXlJX5hQKG5yMHxGRDYP6OJeMFkVXEdPoH+a7ooJV6t14VAitvZ7
zoD6wtyhXfuznfkMlpV6gmM+k4qSsKGtBAPiuTi9IN9gzQxd0AIcXKcvXOQ7Bv9ORZU5J1ne7nWa
UguNcaSygSKeTPiPv29bF+9jQSYRPT6k/HPycM2Le1eiVjD7XBTFI2PrxgqsGpXmJaM7Yv7wns8w
hWiH4NAe2PdDxzWRAKWs9WnZJZN3ocGYlgrO6gq/TXLdbC7aS5YlA0ANWHAVghwhoraOBMj7mdsv
rmZA/rZvdNi89n1SlF/+1p+tRYrSJE4RFaO4WwW89woQvqW2jiuFPRlmJVeyZpyzpH+bmZwoblWS
t7W2inHU0SSZQjMh21eenlGK87c1RaV47B3gNI6UmxwGueifsUm/Vzlb/JFZnOuQYMrhhwV3QFaZ
FRhza3mVcZDNGzCijwN+HvojLHJm4ZKXxsu297q2nHvSJzDgOM+0Adxwzz3KVxZW/JaSfPdNhRA2
0HcTzFoELiu4BHBn/5UAbDq5qIm8HR+b8VOmZ5GWUPWhQLDtqEnd5XqrgK0sIwAbtgBPFX0M4YmQ
Ne/wLKhs/4gbZJ/eVONUJL7qQoUXUsx/AOwtzGlTyJ33DeHfExwYSu0ri4wSLU6AL1Dg6AX5rGc+
IG++E+QvgcYGRG36v9aalLKfnoh/+IVK/T3+4PHql4OSqryI6bRtMAOgPj/2oS8q6RrzVC2btfC+
yhLLpWoMLh+eTgyuGR8tM5e2w/ANDXZEfKpjP3kc0SAq7DrvPHeNdP2JraYDXMq5vv1IxgE39LxN
ATEuqsN7xRzUErC4fqJAcrAe+gL+F20IYZJ1PzwdS8aJaXkQCIkNITE5ExXpBk50eKTpT6Ne5GWj
xUEyLfIS0+vHt9jDXmat53m5QKNUK4YB42CyxmCraKdd+kUr6UUBW54aVrWoe/C7kyNy463qCaDQ
F7JEZzwgpZHqwmtfsNNCz3LX01z1bHqThLTHcv7FEQxzB933C5zzMe6+FPy3g/11NRKD1uK4HHy4
FcJ6uZdwWPJy6CBfaBFnGOhFHDaXvzm6w44NypotlfQz+ioy0hnoSVJ8mQymJxPEOaR9zDQX93ui
HNe9FBEyN8fTUsJGpCTQ350wr7zIl0cbkThsRtUlFTRpMs91gtt4U9kp7UVtO4uNQI0kFZDCpjce
Zskjim3VfmegktZ6p9Jh2OCzzGd54v4m6zS5+PyolEk+v0yC08z/+jFiPJ/eSh5uj3/+wJEDESNu
Rfx7hGarcD365yFQrszBJrfAarqkQrEhToVIxk2mXzwYrZ/VrwESYlqKZMEHw+F61laC5K+PmXlR
iQJlUNgd81vmpjvTevzs3BItENyddfaSuzdqdGKDhfp536XHQgm/fbvVRUiqNY7q2rCIVB6HntOv
bWIr2RXqNnRb3ro8yrw0Abw+4ZuvWDJ19XI6hpb58LCWaGEkdgSdv/QR9+gcMiHJABgu/OQ/J0a2
Qo4MVRGbc00cBUWp29Cg7w13HZ4Gv+ReBrzTCUwT68vHQvsg67CyYTkEBjF2ROsj6FHo/T1QKTOy
ktaOO8v7JZTIYQDRPC3DaZ/U7IimXAXvXY3kTcKhLuKGuCU5Cu3eMQw5l5kSyuv0CmeBbjlrp9m5
LFV9tEZwH46phSffIpNuQvRT1L+WgWna29f9KXsueo7zwu33ctMR1hTAE2bLRC7SMP9nEybrPMDT
rDUcwOlHReGHCcv69icoP87Jq6DNAMTQvzS2NVBRzLsC1rbdXi4qNZTY+GKCwh+S0YCtSE8/KeeZ
DLzFrXKMrMVDhx/hs1dKzspZ9bhBb3Eik5ET8O7yuPofKozzqOC5bqIB//7XUnhn8XYEmuhlW1Jt
5XESblImHzVfdbsRcW7SMwS2xbZct00qZVMOO2bJlOjmkZSSW5UraWIYgwCNE+b1xzYt9mk1iEoA
+cNMCvKJaio0yEPLljmYxKGrcfa6hcKQzRL9PKj+KqhNy8BMIwYYGonWE20bmJt3wJf/eJ7BOYJd
nTgptCpmuXswIbWUWJELk5P4zSzKQY7zvmASAaWW62L8gzGvUhcFK0pGNnUeo48Am4N10sdMaZ7O
hrwew50vo4V+FHEkCDg8k4v3/EjL5UoTFSpqpyME/t4ALosE07uf3O0DaQuv7QCwY+hgQe35xV3g
jULGHm79qozlNp7dqjHbYU9LRug+4jxAUmanlJQjq2g/ezm1KI+7ig1OirKeXN0ZLi3eLv7C5km5
2zNOiJJn0x1zt/B9hnEEowI85WfjvMha1fuX3NXAXgJ2Pwi1IEc66ugss1NPlmiCEip4y2hCX8dg
2sQTXOrHylWgQZaq/Bv7gMyNFZuALZK+VEfUGMHyKmvmB14VTTboLonEXhv+y/yGdcnKEaUqwfdI
XCwWb5eEPPlTQkRrq43ts3wMUscXMqSs+G+WLg3njwVtLeCXlpWTLTUxuFhjmJqxdlYQ2WB46CAo
gNBjwpt4I3dj89OlcbC0ratfbjImsn5yiAa2YCKQQcG//iZ4KoMfxuJadSzXm64mEejN4mzhp3eU
xiNAQ5Ky38elPEZNZLycr7CsaXNkh6ii+PNwmpOViZOs3Z1vSNOozdRT+sJCWdduwEgreDLEVvhy
ZY5R2jZyAmCR+32FFYKh5HXCa5E3xKCfD4Ubwq6FsGya+lDHCf9a62/ROf23eWdGtI8hk2iJ8go7
Q6wn4bg0+tJApDFNLV5zROTKXlMQ+6ZUP4nw6fxOHQhljqBj9Oe+jZ5dLbrASyP9wvoy6BVOnCvx
ch7LbDrrie5NldJEcsfFWUwdPFMgoKBlbDruH9/CpkURmuQoujNPvTbUGooQeHGZSCKuVIUKBZ9M
qSy8sZPS/dXcjZjmoHnhFdMSxSKLTBqAj7/m2BbgNMn/kqPqpTACrR2KPLSsf4CARc0vD9bDJqAz
KjEc3xRyiWf+0QPa4WjWNjTJLyjXd0CSgMKHRlwxZzx4frQV4B7Tx1Zo3hDPy/7eGISIM3hodskp
45CCxmsNrnq7Zadnw+QKYD4zWtpo+FzLnG1LhtFvVK8Nh4cEysdSIxlXOLednWZZwj8X3Tjxpc2f
bFwQ5PsCk1Fh7OejEdBP6qgyvLDROh+6IzLwN1wKsouyM2hmTxfEQcraat+NgPvt/LGjFfKwR6zF
sccH6Tb7ve17saYqxVCbdaDd2aSpeYVitkaVE+YD3mAs66y1UTWIQZxhZVivrCEnqPZtsi0FyCNS
VhzwpIFuJ8X25e42He+sp0dwOxssO5T4BP84V/xU6YP/BRFOunXcVBuwYk3KzchsI3SQn1srqTrP
NYRaYLpNTBNTH2jro9DQNteiNCmeKD/nTJXNqDCXH5zAW8vwPDGm1fK9toKPjDZvxcsmcCnHuSgw
qu/2OBByr55T5nwRbZ2dGq8edKB+UD+MvBwXy34zRSE6uUhAKvel4qVmhPDdqRFVofEzj1FJi3j0
AZu0hzqXdFw4kejthHLDBVsd7ZYQ8xI4QfiM6naVj0Je4C3vu3sVepoRiieSdA0CdghR8/HcMoch
ZcLlJlGLUkHqfk788C/n3UDHVcDNUFOYSl/KS1OYFf5s0Xcifa0WFs+7rOW94WQRWCdBP7g2wVvg
GQkOEl3X0Li7XGyHuY+Y7CKjl3rLDVQWL0XtvBv3/uLudbeTuOz6hXu7FSKOO2ss5S6TOqihLd4O
xwTvHRQT3YzgLFGi++F/84wdaYcPCiYRuqAmTZHg940gNfWE1W1y/MAkdDa9r+7hARD/WQ165rMS
kC41LOylL+btrapadSFJTW7K9PAbDmT6eXnWK6KUOR5AAbCq2AMiyWltSTvJEeR0PCFx/xrFr3XF
w7wvqepvjpUVpYgCp8lhpwJ+DTERMfMnOYybUALB0iCl4BfshfpsHE6dJ5jhyGeYfybqqUKBGdnK
vcQG6D+fgAtDX7TSLTNEUcepNNP1l8aVUL3Bs1J5Cuu3v17NtaVTk3IE9BLQXrlhbSI3ZLN1+gkC
mGz/63H2GRfCb96vwtOFQc1KxtZSpTLRc0Y31Bk6u8iz1rZQBUPpEM2Stb1QB/NmW3D5yapyl8Ic
Z6XYMpZ8OxT4kHBACKuKpCJO/36a00pgkoZNORT0CkYL5DFjkagq2fJlp1FHt1PpTYyBfxtDC95B
bU7AXwhRgnX/9OiPvseHuR4702lgZ5jfW0KfuOs0dQKwiwVN2tsYn7aOOHxLWYibm35aICxJaid/
BGPayaF/vMU16ptFzPl4vrvwShlz2g07pSWxjoL33gAJXH3QwfKvFLgFfgO/CBwumr5IjLtm6fwP
NjiFAkHPbW+HD0tFvoD3GmIV8Eb4xtsU0gHY0Clo/+xAq+qsRIMZ/Nk294o2Mdgi7Tjur40r26BX
Pq+08LblKaOdyA2IPbOMfaVXcAijb5i2T2P0ZN+J0p0B3Q/dB8zMALSxGIFKmfHMNHavFCmmYiLe
3ZMHynzNibvjqtiweoq1t1Y4xq2XgEKe07RcJQvLh+doyOhliNRsLkcTcNF/JxyQuG6zoyev/LUJ
5g/8MDVOGt6p75ihn1kCeSWhiwlzkYxjbkJ20SUcBmYUcUwnlEQlRqRZDyFUqLi5j7EWj4COE6FN
WVKT1zEPHIWseOE7YsHrkDjZtUzEvHnwIq9S993XOPvC//r+nsvP0+ckyg7nF/eXrx/AaDgrHTp1
j1Wg/FncK5tC76Upt6lmyiwJRMY8tcnEMXw7hfjog8bl6aUIYelv0XL2hZwrJr4kNPVkYkkWBIZC
ndLxZzyVImB2SgihusMyIHHjYIsktrSy9pSuAoTpFsHpKZIykDqU/YFFoseKbCB5JlmuBseofoSD
Mw8P+Qrv7D8SrHqsGAuJK6s5Mlar7hGiaEhqEnjaa5vjrefBfTcdWteELClrmN6Rmk1vsXgO1hHQ
uGfpHjwqYuLNVMwhqBfp8h/mxqAN1dHZdqEgM4nHQxvlmZnpBeTXUADLdDumR0g733O/n6pY0NhD
G3eOY0zE6DffQ/Bgs2eVEeF/j2oaGka2zUOMcyv4U3SwMZ4lbizTUM4YBHpQPzRG1q0meqqNZ9M/
B1Avco/eTH9zOwlbgB1rUW1LNERf8VnPALO4Z+2oSrghYPeJVnqwJmTcrtP1ZitlAAyWrFR7GIL+
bXjygTGEe1yHEBRYY+W0oQ1dAJtuDgY4ubmifBWgSwi6D43vKmsA19gJyXOvOD20525rMRPTvbXy
q3sO62/OR+ljZpUOOiGxRq7HhdHqZyzjlCXyUGgoYx2fM1okHfFAk/Wo9PYiY+BKFD+LCJnacUo2
ic6t6uYNj7cmcVQGpmVLE0R3/wSOGKmLWOcXvJAqKrjJT9+RiojVV34M9+LjyoLX7vVvntOFdhQo
Cc+LhnsegKX/HVUPT2PsGyQt6/DEWLwdQ6/2Bf/peLgfqQI5OvnOcKGPxKAvplUn/kpMOinw1NUC
wC11+fXRU1i/SATjwjVbzGk5gYAYA4zmXbzi+Wz1dGLdFi8U5ck+KJZSy5MaMpF4xtw40tVEd51S
n18pGNBaJGsQbwksc9H3Q4Mzf7XQXRtrrT/945h0T0WcVSTiobR1ctxygkM+6h8KX0wWw53YJU5n
YtYUkaqEUkiNc5ru4Gynaz2g+/ySG1LlqgGOWSiG7a3EkRamxAHNHlP0JKdKam3elHPqtrmyHNLv
jWYH67HURz50+GEtq77XBFWgrn589s8m/3EE5H0sx2/VTqsU9k2J5b90Y42Dg8v+ZGHV9eelnNNd
OwXZtoB6vN0Rc2Y4S+sv2ZarEm69Jtvp8jpDnzEqvoLHwdnWOjsaif7W+oDGrmzGM0zgSGl3BFUK
Iu7/ADIEXdBNHboiYPYQRQ9XLgdBG1oKq5CXaAbHu6pBSTJawRBpUx0+axV9MRuR/rlYbS6oYrwI
oSFMZzbo9jls23m4gjIAilqUqP/VlCMX2EK6QO0ljPqslCYOa5NnxHfno9jlX3YU8nzoun0GTm18
0sc323pZhuB/gGN1DoqVB0pq2hsA53npbMQ57kwxxmhWyM8+1eNFRLhdhztp0OAYB2KG1SZnv6I+
gCf61bLJQanTGnbaC5r21Y3JMULmyYmHGMD9IXAhWt4Aum94Smvgbp8QOmnqv/Zt60pHddxvmJ4c
jSHdF35vWJClxkzBA2RsmfmMwzOK6KjsIyhe0cDnVkFDab0VndklMKZyU0skdon59d03YyZQaJ3x
wksHx2QhNmX5U0gYnMDdJ1a9TzKdIPLczOpvFuWR40KyRT0wvsGeyJAbHZK4t3guBxLTQH/jnRiG
x2y5rt/U1/Fo1X6Xt3JYAjzX48gXunCVcO1I/266KruhaAx32W1E76OpvsM/hf8gLZiYTJ/xUxcY
t/cwfzXZk+xvfOm3/LBAbNStDqROfrBOk+O8u8dcu9Lh0k3H88QDrWLpK+LJbu2BC3OCt1EWrlgz
XByi6uyZfh1K8+TefCgBigwF9ahSTbUM2uJqnoAQdnMce6Th/MSFb3f1/Y45vkSdVSho2iDKIW/Y
Y/LewRMVSY4+XQCk2Cd/GJfwPohIZtGYjPrAkKqyo/n7lBfWZhN1mn/ZBSXjGkhAkWWkwdqI1yP8
swzgudfXYYRjUxhqsdOPtxA0cxAlY3J0MCWdLKMvUYmcBLwBx4r4QVJ8+eVNcayCk3uf0+jvBL/S
wjVMB/lwGXs1YNHTAxm1IlTszpuw00Gl7JmEcufHQznxhT/ZeSBWHHwFnLgFZYUdkhw3Xn0UGKDM
2wo8gdnpqgjBl11l+nl5nBYtfaCmKke8ahtSuuCqX9lCDZ4gF2SBjB0uhhHYOX/8cqr6TDfKeCS9
qzu638K/hbpJ2lS9EJlCUVcPe6mVq9LF/soIw+7T15f5nbU2+Aqd0V23EUfFUXpN7QcguXiywQM8
YJl83oT3MykPtjABh8qV9WAkgq/qUOsJm3GXBKQgfaIlq9jwDWRB7vPK62Tgqvj1/WuLTP2JOYxQ
p3i2LhJG7BbUCTGzmnPXyPUUFOcWNrbbbGbhQ8nhBJloZ5riyJtd9HFQT+BxJ8dd1TU+IXAr1luX
bDLfAqVZ0UA9+q+IbWVtDsVc5AwPYC6NnakskrxsWccIdCgBAoIxfyjiQiM9hdoIzGzfgcDFMb4h
OpQMnmF1RqitW0Z3+cbHP/2J9wF/XwYSx8LBUDQeSRNb7FA7GpgB2r9PCxSZaH2zfZBM3p+hDth4
m4TfHkiiN1dWmAqRKo5PjlJXsxOjzUNDUqShoTk06dqk6pPG4ZQvtZXYqlNmkRdGAOKhBmuGttqU
mfNdVyVW62sVjLATFN+yPnJyl+2zdFFgmOFVTnOnDfA3FuGSz2tprIggFiF5x7r0fPaME9JCO/QM
Z6k8pgLHSPK54tVoSOa5dIrpIyF2h1RamYZ2TADmiYRN+9/Ha1OU21d2gLdAx0i/IgTvtjAj1Qgh
tGFjpgYQ5vmfIIdX77VHKJB7qQs0aGu60hQ88eqEqAuFA8IJJITdIoqigKoT5Am3bauPzmA0RtX6
pM4MwTd5KK1Y/h+fOoerrwDY1lCXKlj+Ra6JmoW/DCMzhyOrAD9F9oOKp1DJ+5mQW1Fw8htFdMu2
UNC1BNAXKj0xhcaCrsvIqsAswkTytDcarg7nwKCrFAPQVfpK2+peAjAr1w+RbEZ5URERBv0vd32K
wjDyMQ3N+sIFdj6G5ti+ycZbT6LZm19IV2RsWb8yU2cB97t+zcE7YdlQoKTVyN/v2DJGWoUBVQyk
T9tcfsZArS3EUivyyf/uuJF7r6WRIHJxKbyMJfLT3BuSN9RVzGNbXgxIg0ELcBCsIRk0zrl7Z0i3
NSNN5vY2u1keca3TvspUjfQdzfSm+B+58jmlwU+FZDA6N4T8UwAksLitPpdzdLCqsYpK8jFn4MN5
Ni+PYRZrb7uXIj2ThX85lvUctb5VI2EFX39m8mJJKIQ1R5enqJ4XqVCfMadK9MzOiCFv5BNUMFJG
r5DYM9PS9sErQ2KJMMmrWOYUPNb6os1JwI+5jACV64WwiFiMXB0G4onQKI1XAMXNOMHewo0Q1EhP
Axl29qnuxvqq8YS8k+vjx1z5615uTSNVmdp6l4WHZEUFJ1i0GONEN3Wnpa5mF+gUdW2QYTXK/TQV
p7gRwQ7QKZQ0u3pVyUNzuzB0R7WZMxctasGJHDYosEPEIqd++p7OYJM3WAu4ksE3og3NJzLE0tth
0bl4zyuCP/+xsARIxKPuvwI1Dky/eYAIJvj8R7WoLCtwdL9IAIMa3+w+rqIAgCaGwOUNEM4gyclA
/K5CytrtDE7moEoLl42PsU1snRnyiIqezoqCNPoEbT6WVAf4kBXyOTKj3oFXi1ZgxhjudvsCJ4d2
ZdJGiT5Pk3+1cGKVj7waAFQmEdB/W+Mm0+LmQmR/OGwNGGTdFUlrXnqUMU6ezxUxaey8Hk0LCBM8
gnKwSyonAZorlRyTSk3VA3J2Zqr33jBzixHPPjTuSIC3SLAXi9qMaNCD2tI1sMrc7kN7GB/jPruc
rQkoF0f0ecyyPRDQ9c/1pd3SxtjcQZz2tyUwnfMnv4V0XsNGPR3zErskr+mxq7P0I0nQWE+ba3LA
9A4qMrJ+93Rp3AZvUUVMTdWmzLP/kcQjQxIbWPdy/W45PIUutnOanOBlML6eYvRMfizeLevKA4uh
E7b1DrP/dOyEvVVocJooNuIyoUf6c64+C7ZEaXtcbb6oqTfbloFHLFN2igRIkA5XU6NFG3nkyyBn
sVM+5ZpHaTBH4ucx3QkSuSyGEGMGcMRzB9MbkFBsmTpxRxrWAJWZOVMir7rpMNjf36GZOy1ewS1P
eRm0StOEcpkVss/Swf6JoMjs6PfRoLZYJRRevmLodzBhFh+Lw2shQD9/rGEej3QpWj1Lmt25M5qQ
l8FajjiJ4CdqDw5NZRj2Wts/aeZeLAH5mby+jx/+oYr6Cg+Vd7WBN1ikQGZjfIujwRYnDOBD/sLd
J+qW7/A7AGaXuFR56FE/P/Cz1byL5vpgEq9Pz1YY82MUoYSWIe0unonQJtm59ViofxVy1aKDNDgz
IKiXdIHx25kOBCyLAJ8mdos2sMPkEDgTCbasMM9GNNTkyrzU+e3Hic8a/qXBG+j2GlE3vZBC9bq+
275Cllx3Q8ugN34asELq1R7Q9GYOedadP9C8StdiDETCObKegnEJeQlooWQaoViMKoPM/KxVioUL
Ri6VPzIBDxS1eGrufpFtdUUkOADg24ahjS2vFAI4mnjjmC3tzuanUjerIZb3VaKisoAnOUDTChX7
VEKKbaIbB9BhYv1zbF9/xkBhbs2phSfXNVnw2pXJOSscHILzdwBC44+d9y5gzB3yDD/+ISJw2hqK
1BayEGNcwGSwvzK5ZQRffowq7dr40umJNQuJ/DJPIXxzIz2NjQl64dDEVrCld4qJ+NSFObohPQGi
VRPt5gFFZhy/SM2cVPQD7k9qVmxbzmmsZpAc0xq+X8HQ9SKzefz4nF607XoAMU6QMdcvCkbHohkX
/Wrn5/BcuocV7NHJqH2hgTXUMJ6Ryk/4OMhY7FTNo90YVGe92MDbgqjc+UymGhdPcnMxFmYlIGmO
fNCj6Kugi0cxpTTpNPsmQWADLdzv9NMN7F8r07t7P4g4LsApuzzusKf+2Z+f09YK133K6VFMKjNd
TA36Fqona7mErDQpQFuJMq7n8i6hfxTktL4A+wrirLnUqokMviyyHmPnsgtBo4vy+wl6qBRS2B4F
SHZg/Mn4v1kcXR+QMVCF/71ZMyyEg9xQkX9nvCeHps9SZyeaw0CdHPgLo8uU+dqTDBsIVy0PLzjR
jpHsF5JCExKw78kKk2MiYEIRVw/jRrtbppw8cK6Ewt8jQplee0kOKJq5oqVpYvOxZ8cfuQGL6GQH
q/QK0g15N418oHLKxlqaPO0EVFQtvMYzGkImSm1O4xGgybDOXw8pjyqhj4Iv2Ls5qtmEJR4VRq0N
+j0GhI9PfTvFigv40CJyt5xr7rH0ORsN+nJXFVQH0DK/bZAVgIRtb920u8Tp+KUflgS9Oyn8TOry
3AvngSorG9D4a3agN+BL21ctRqt2kPVf8Z3DSi/WaWKYhBMCMWjgDwki3kNNfSz2XB5Q5K+Jrk07
38yFjsr0w7GqYVI7afZur+4HJ1LyLEUtKL7nUTPrrIlb4Mr7Pq3/7EU/OCTyk2SbU+fHm5PkV9cy
B0uDCznhzJKsmbXJB4+jtShJFYbxDp2BXWpYTY30SkICpgX43sfJDm9n7eHQ9TNzy3/ApkumCO14
ocyPr0s4mNJi18N+BHIZH2hsYA7tp+6IeTG/3GScAlstnvL+BII7yZebD6lf9uSJaAHBQxGUIulw
9C7seKYANEjphTE6qN7WC07dWDOK58/L/Rq3e+V55G4sNWdh3WUx3tMLXbgwMiDSMeLDJNs9f93t
UyZKkWYBFxrEBxmq1LRIRIu6yhBWzvC124+1SWHMIkd+YNuWwWiopaiUpKypj6lV6VaCgsCDxpmG
8AqH3cCpX2HEdJPtnSojNVwaHtX7c+P2/6kij7RQ7pvaiKvl7gcbRSWx6NqCvg/Wai2TgXc7n2o5
14UiTYzY8YTSRLOiifPXLkfjOTZlsm/aTJcj9Il6/pWceh+/fTf4pn+f/7k4irq/NDCFYsxS8mWR
ZobivBzLFlhDi4psCMp2MbzO4h8Dr1HvjED7dDDrbWWh2LuGEsjRi0RkFCjSGCQ4lwgWliklhXcl
oYrur1KVd56ynn4wRELY0GEh6eHfkTZbNOv8llPFpQ2GZJq2HOTDSBkbLw61pfslL43EP8N1wwmk
uDBBpsFhJmBPcmi/jWUIpOSnvyIVDxjClsRk/hPr6xQwc4Yfat0ibuymFoWko4OeJfTCctZZ3Em/
0StOmUL1P682L5/LKfZsBUF0+sTc9ybysh1OKxmM/wb1VB9yeTld4bEXr/vhz0vhKt3g+x24SPLI
a0t/c2TJnRdb8Pl/oIYcLsR76fSf0wspT5u6llaLdxoTw8AXRge0lS0MSwoTvonpwwsfJXq40RW9
uYnOB3clWz64wZh2icyn+X87O5i/ONmEWBDsvTtx4/sJTJkJupPtVnIED772pHuslzqhicbod5xu
Gm056smoWZlKQ+ZhO6Z0hqxFLAk49gUAS0mOWDsHcICjKOblfWwhaA5HGuGN6Zp7e2rmcl7r84a2
RZjARmbcDxbCAlqLRdzpgxlSTQLdtUsnInTdOV8+M6qHTB/0YofL5enF3si+EZzCd8Ao1zT2drWe
1KWQpUzzwrOG7eADf6eE1DDcfqN4cXwoc5XnhRs5fbGCHZ+SWv8d7RqWeEjFPiwzfZqu5WsNlghK
ae00d5qO1wZnn2+rC8+ks9GSOZI9EQ3X4rskQ/Gn22uqkx+CBIYYPM1LV3HoDEx5i3ZzihdwjBEw
N9Hf2F3nt30Z4Nfgnt9a69/vggGmGIF+rFjkN6oIAHmH4DJKJx1swz3ZWQ+E+BgQr96M8ApH4hle
LFea/TEMjEHZkQyrj+vfD/gvx48g4GZ4zuabxSuc/OR7yqEH2waZzHw350rRRAJLBB8s6tUr+Ydj
o3gXEvYFIhJsFJrcvwdaBZhOzY+a5BsYhcvN5RW6i4iCh9G6eLbINUzaZT5EvKSwUdpzFhS5JjmW
UOhRHpQfNTKu3+jOEXN7SfO0b7CH6640a68Mm+ksvbO6rOVUd3o2TDyVMhTgYNRaX/maEqwuTm//
rzHdVJPdVhMAAyA15QV2Zad4grUaHcBP091i+1kooqXxH7rJujYjIpu09zRCoj3qRdW3Dl4K8X06
F/QOwFWtgwQbMALcZITvwoJhUMsrbycJXcAz1aKl21VLq1w/SC7D/jlzGmLtn907G90qcqMxJZ8J
RIS8Eu9a64HwYqj8coFIKjbS745OJSrpjXnazNy0eliam+aSeedAnQYVbX9TTNUv5EXOxpdCBWAv
eyS1sh/cArez4B7+rZ6RetobpcsZxp/03oJZX4dG22sd7D2xHArj6KFsKPXkasIddAlHK6VVA9yV
h5bIlXzSGd3ZoFR3yAeSuiSdmhZZLEXXPRb4KQ8IkNqAXyiawf1665+O+HQIFiC0PbVS2cvomcMz
Jton4jL+lF4TrVJ9gbmB+o2iTGolBKy9XLWlcvQUKaUGXInN2/qQ2hCDGb9AEJlmFJc78WMiGI9r
UhS9n/leHNkPU83TViYZJG2hgtCIIuRU0X8sQrQIKaiA4XenLbewz/ACDKftBQ3wdYoXpSTR4KZX
/tsuWtI43DucmQ/KJXbzC18OmkxjijIv6/ZN8P90asAMsdZqCuIuVFQqCSLIRZ8ndoqP99fy2lxc
6b6hVxpfTjsVA7YJrx9cA2j4UgsNFAAB/sTURVJMQ7ZELZ3RHZZazOerEJn0aOkalY/ZU8X2f5Ol
lTJy+L38o0tvwyvkOk69y8Hc5pijjfIOE9x5x0Fq1yLdM7JPNs1hbBVUHCullUKFAB4ahlE/dBL/
e3ME/aI/1RArl8Nsrtibo95JyvsOJRwUgQp9VvX142Sk0gLZVijZYXtqUPxrvEJxJM8AAppuHH16
dVIIHp3KW/4fbEDd19ofoxuQdnkmUuTtxtickr/9rrHfW/PlTyGUhMfM1SRxvJeIe2/8bjhL7leD
DBIEpdUvZDv3I2jC5McYPpVF7b8OfJXnZ+hYm1Stgx19MPuzJvistah/+aT+x+qgPY1oR2ejynU8
2TkMg4qoygF3C3qdCtQFN+R1x/ebu6U62VUtLq3Jy9k0eiR6yf4Uhc1hZHKK36lCnCe1sy2V6eMp
Pdy4F20iUvQAg001XszGx08VbM0lJxIFu6Q+0pfWTXX7z69k/mTzP0+5Br/ul66stdYVJTGAzrUh
DC45uRsE9Cu0DOKN7qH2Wj06mlut4tUBUiEfqElDZHfYT4gtuZNY88GsvOemZ+vBKNuQeL53QWxL
z89R2U2wGj5vEtlTPZYS1abVpn/3LF7KHpN4iPkD5oOFyQwRpnps7frsbGQhwG6vPxzKURCM2MuH
aaY8FAooD9cAm2k52mzlb3MPLQUPrq1RtozAnSRehRmLmM7cs9TOBPc4tYLWGeRZSHnBYCSpAvkz
uIP7ll6eMclvHktgRIg+urXOdKi3nK6Uu877iDeA/Ra1HIeZo8ONC1ifQj3nYKrRRwnDYN0LeMDU
maja3q16Su7zzhTnM4fnNRYKxdXcZSnwF5YrjM9KDblASutxXueOS/ukUiZbffgDjzOsXhBu5K9s
0Pn9jaRiP8Y+4kQS940IS14l+3dQirgFvjdTR7cueI0EiOqAtYtqOiCLOBeuOh7Sk1YnoZ+c7Yt+
xLu0mRo6Bp++zj5MAlcRCrYrXbFwFaz1zdri+7K4PAVrgewrCNVWDfe2nyEd2oooKI1P+HtvT4Lo
z3q02ggd0MKwcFYC2S8AoaHDXQzTN7rUiG+QmODE/jwAU2ZfWu+9ZqVlbQvnRaPTzFxuY05uXGXg
DJuhYVQFTMoial9d/45WAe1eSusfTUPtTkqDwJqL5p6+sZHj99T7kdpUe12tr5YQKMQ7Lf8cHC6+
1KDdNlGkgqnI79lTgOZJ9Ab6KR00hm3bzpDnqHrFYlJRTxM+WqkQOwdFQL5GzN7H+zK5GqzOZ4hP
dWczzI1KM+QlEQYcDRwgKNxLcfMMEvcb01mZJH8DYz14SeSXTkP6XtuwgJWaAGng2muMRZ5YaXaH
ffgAdR5AZEBf3cOg4CN9AeFUIsDxaC5kjap0eFFpLYgct2ZJbJSUkJ0w1hXI6RS8A3+ARmHsTuiU
zL0BONLbc9IXwWJIFNShcHV8cnUCyyNJSHqg/E12Ww7hvYwr4QD3/dnEnq21i44BHtihs//Ga574
UQjlAY9oX9mV0nqdONgEUhTyKGOJZXYEOkDqir4PwAOw/NUvVu7ED64eZjbsM4+zND0QE5RsA+Qh
oeX4dLjqhSjcKe5noVUvDwMs5UH6wq5gdObAtJaljjZoHtWLIDFCdrJvxDoFFEElOAHTse3oKg+9
zslpkRxs0K5ufs8OvuetvBdWeL8DGJGq5OL51HDJgiZ+XjBE9R6ugWGhSmlqsLIim4TJD98/+20m
DWHXgLMkey6/EOZhMZI/I8goRWxaKI9VBiieTEj/QmrrmOapZDbg94Pxos7oO83XAjEuPRBImzG9
oumg79BhkWHn7o5R26aOjB22Xd3uYbV6Zq/TZNNS93w0FZ7GKychTSuJiZUx0Cph7RpqyGdhLHQA
wM1UVJb725FWmotbJG1ewlnFfgKEEcqEcZVXjuZwly2+Bnn1lNXWjktVQld8HUF/sxBlfnzhETWQ
+RDnEySI6eAvS5uVgMzhQgJFc5+z9LBBMDnXSCK8JjNWdHO+j5GSyuisSNOmqUg3+KHiQgkPGDuk
+KAkzbN0nv2DbetNAkNREqwyoN162XdKLkW2aJdPnW0QqDy960usiyr5/LcO1yp4CcjZ2KxTnpUJ
H7qkOgZq2ln582Oz08Roe9MkNL5NNuvKCo1rQYn6XUHaE/gKFRQ9b4g6a++n4LP/aWUF8yWRSDYB
eRtpXc0voplKJCb7OCWG0l44UH4GDSdsOlLAzTT+4ktkx9pzEIgcLahIafDNgggFUWhAgy8VEgsF
DgswufDLlTsi3sZBi3gFL0TzxOUVA37QfoHJmombfFbw28CAA3Ihq9wjKqoqGjeN+COTMP0XA78I
3HH3P/49zcWy6BQA0fd/A2rmjRCe5u26vlkm5i01rGfvvVOL0IoEiato7EL080CKu27szfGSPJNF
NSZrIO0+lZIZmc6lEW+H+jLR9/Slin41DXodAtZutwv/SoN534lxNB1200dqTKefeuziqEp/nPAx
vutDIwe1BnXGhyeOopNsL3eiVGLCUuCrplC824bsHnRqgvqMV6m8QAjrmZLhHWIAXr7M3c3ezsFG
8Rdhxnwjn0fIo/B3+S4zsWRLhcyLUxdlOR+hCTtgzyoVZXz1dx6yrhj/zLXz3kz0Y3V/nrIt8n/j
sIn69Js7NiXfZ1AdNKMPDuZ0+FnwHmqebShVaLY7s9VB4pes3qdgr7+JKB+oQ31uD71ET+LJW8W1
myO5YHStxf5vCi8tWzw9IFgnRkKKo9cajSNuFeNdpUhhR7QS9JE2+nguRWXuy8hv8d1VXCnju/9S
9WzrSGaFkFzB9yuBF95+OnHq0UKB2xyBN6UhGpCSyfmD6EAJW9PG6GT9cYbMTLqg8gvQe3e3KroK
mTCIGe3ZE+yGg29CObRRdxFR/YXRz3kF3b1AhfBkXMLhTJkgEsjptNno1yLAj1a1qxLNsyoAk0G/
iXTLSeqly2w95Dm0eFv40kXOsSvZNfNI6t605rlsDJP7YoXjAB2YCS2Kw7GqincjUdrdmgtFAZJj
vYWEiD16M+gfrEYOHOs1txCPI3QaHmvow6DuVN8yqb7cZhkhDue9P2iC1TCGtH34oQ+LJywPd3Gf
CKnClCTbQ475sfPQZfWGf+KOJRuVL3IwIBFOIgvlcOEyUgNud4fTk0OZufoKY4HVo8GwCqUpITm8
gZwittmFNb54tdFhiKZgETmXQp6Cls//spr21rK1h6F8HTbc+wDO6R5S7UacMnG/vvGWcOZg+c0l
fhiL9cNnOsFVEZYHE8UTYASnAFr9sxA99JnDDh22YhiMcSCLGdi3xL8W0oBCO7hOmCVZwhHTvqZW
ao2sSx8VORAVsor4bL1P7kZ9R1phiylwgY+7s9FcuR6z7PWV6zfHFmOJoKO8aX71L+5hZrcqquxS
ZEQ6oVjmrd3LPT4LiQdBEruHYvgkAqowuxlU3OngrgegWtsUBsxACp2bEhDdcY8pmhMlBaf9VgA0
3tXjf65b6xqMVGp3urrtg0Ir3K1dzty+ABidWFNlvmW9dlUWFW/Bi7LQcQAnPGttnksJERiIMFM+
CEk701cUF7qL18xiRMwJNBloHzX/uTNMxiStDdGrk7oMr60pg7yuA8vMVcl5i3OVECaU8Mzh8e3I
iysTmHHAjPMXOHQUK1wP0dUBg6MbbtGZsNH4Ae0wawty8UN/KZZ55kHgo34Li7huiw1ZwYH9kdPC
DVSeTh/SLeMD/3v0f9Tt0TESA+CXtYDc2+vU/bxTe+QoZuwOP/QuN3N4CWCbvxg3peVXRMy6fQAg
zi2NBXQYTioA4Feyse5e+3kdSwkY5y6kHAZTWyWLbNBgS76sZNRDCFOkemiOYnRdtEHnfmsWEaCM
ioTR2xGDYgNy74+Q66ZnooGc8qEDVFcUc5DiimBSLFw90466SEe3zvZTYjXh6XkxiuNd1phvX2vU
54qIEIAy3f/AjV8T+W/gFYraK50ovpnq8KEOU9aHVlatHHV0MNy3bKofQ6fvBQuiskgi+T4jhgUU
s2cBji9U+8cSlQLX6Aq4JaJSfw+PagREYm25zXbqno2sBuO+GO+ZK3/GoilNDekH7amkGilkbBU2
iZT4mt7yuJeR0wyX9Plw3YXkCMqnybAKwqYn22JUR8H2jleLurczZe40OmUJvRBcbzQD1aiAWuIQ
sQdE3TGm/geliZpIocFQbS3ioJOr+Nz93q2/9xzM8oPDB2SLT/yfk2x1gP0Z288FN4x25g3/YQmE
opQ3V82jV0DCJbqwAXcTjMK10XDArxf2lnFb3KWPxT9hdrPY35wmTDi4i0YZYP+L1xrQOd2v2h6h
1Yifa0ZO+bYifitc3P+rsFsrrYskK3tpxvXMiEOf32MVMfDNOdUgiWwkDAPqvg4gGi/lyE4kVOQr
DnumCCJjHMYXTzdUethH2j99sI7Qht4pfE6fnJS++O1oAESW9YVNR4/WhTEqvnDgCnFXj7wODHUI
/Wwe6/ajqvGH+BoSQ4irHUcidF2XnroyxsKfO8DsFWYagoYU8xa4HQ1zpjgJOWqnirEspDOieN1Q
flimSJDL3riWDPaS4DkcS/psyS15nDwz5qpzLLXe4uw8LOprxaYP3gdyfMvjc5qkzfGD0/+AiScQ
VqMQtp2A9RODAsCHT1H0dFwqzn3iYoW8whQaDvPKdRs0KlrxKaLDQelcpjNBL65DIS1wfFT1s+a3
C5y6kowOBA4PAvETczoBRJhqnReNunwK+r+7gcJWUfDUAMwK4H8pAldHIeDmIl5mdyfiA2aRaO1/
fy3U/ezIG33HV+SYn/1ra4zLI5ahUCOf698KgifHGIp0MOPYaUGJcu3QDbFiQt3+UHs45VmyCM90
lbiJgcCc+T4l0lIv9c1pVkOpwHodRfEFDMp71PriNwVoKAtTkPYFRqnfyt36bH1if5o6Dt2jLL3W
SeZIK/bSdFECjR705qxrx/p6x8k2Jjg1Qjw2E/+29beUqS3LgQuaWBVqBL3b5/2K8AcX05NhX3pV
Fpo/76PFFAdDwkGd852JgVYeCxu2RijdtRzQzUfbXvqTH8laR8UfsUnnIC9XxevpHe40EGr2NgXO
nj2uaTi0TiMWd6UjIsTrJ0kpCXh8poxXE9TY/uELpkyyTUq1sBzuyqNmNdGVlj754Wj2COzRzFqP
QhdbpOO9AZhX8QBxrE/+55W3wgN6yr18wswcrZqDpq1U5DS2M+5uzUYwetAeBcI9MCKrebhTDA22
PBgiMjj8PSlegcOAx3y3FZbLrphPuP+JIju5+xtrEUZFJ4g9IgYa0f3BiHnpsUWePCzmw72dP4pq
t47TKhX+nv2IQl/PPf/0o98JLGVl1GMfhVaM7EV0VUglqYhoDLIvKHoub9yOkBjrwzuKMKgaREPQ
Q5V8nv9kK7GBKL9gMIjhPkDYrwiHjwU6QG7tgMwxOKvin3xLNgf71XKyrQy3hFTaxHIBGIjsNzsT
gtx1j5WGwCKDyxE4JcNx7OxbvjZICCAQyAkwsED1XK2GtuIyr/gfUisJtJ9XGw2Bwo0xGAAMa+2I
cdsP4DgyNW+/zFDIAg8ilVCjCri06ncuV7lQaQ+nV0bouUYb6dij0C2kLMiRpX2uo+m2OCR/lBEG
DmXeUt8vGBrNNlqtatXKBTdXsFw+422cIJcXMzcQB1Q1QvquqW3BWCNXeI67e5VwJ9LBwo/35Eoh
WG+2XyWQIgP4om2ZeCvvBKSknXa9/bEReTiBYSdHFzzBx58BbGzbVbYM/LkYozQfuPAqki1/SJUY
pemObDUmA9023ja75GQXN3puQvCCwnoUx2Mhh1ObT/+fKfXoaSKLQBF9IHSiXVPkea1smKw2OoJl
0DVpVXy5T6NdDYug0uo9PRk6iIHAH28oBAT1HDcst2C7hvL835a5CQcfHWiUj6GGWwAVCG0ZE69U
czrFXVgpKfgk818e3t5C9/ecxioJ3ks0o1iqkw54vQ2DqdV8Q/ZplX3cQ8VGmdq+mNfnoP7GQqis
1/YUGVBgKGMJbTjpOcDcbML2IUUNsSeG5uYkIo1ja+hSrVcDliG4jCB1AfsUqXN/R8wNz1zI52c+
yhZ/VAHXVGBSzXtVhN457WeEfoijckuiS5xxIzPrHuBZv9cbYu30UlqO6o+dkjKfNqS5SxfyRq29
PWBdy4lkmud44LS1jf74DDYyopMV3BNUsB9Jd/xJq+iQPdsQ2lGrwaaw6duihTdmlX4MsW+jdn4S
pcqHBouLfMSnM2tsEUXL5mibWjtRn2OWgxF2h/z1j97vJ3I2c3c75KJJgB68cMW9vm15LMcvz6CN
kOOTAmSAmxlQEQbiiPxBUb1U7Fo4HdmOT4I9acLwX/rwRAfokcNMFHpmseZL5iXM0kfvoAfozoBX
hwh5nxPMrG1l2dNQmvQG2VXNLFKVlqashZa+jtzpqRxTo7UU71nr+Wf9NqO6oX17P7ODVEkK+IVi
6XbbzK7NeUmtuItHw473NC+1cwFIybi34xEPMyru08Daavbg85oQwDr80NSyw+hYGnqv+DPgurPC
S2hQ4NjbM80YUCbDiU1UtspgO2LEmwfZOjcOOWnlq8NPcE5ZvaFuJQPllnX7ofMuT4puFr3GWPWj
hLcP6RRmQvWZ1gSRloKHVQhAsBfekD23ZfYD2X3wgeGZKXpa3YL0tFuWAaPsJvVrz4IKSKnDcjIM
y4vdu3WW7p+HericKDiBFY3X6F8K3hsKrMMYByzNZKTC+et1CeBkkAee39eOhjnxti1HNCEFDmA5
ZWSIiI6G0VJZBNZ24gp2XNwIwpKUevrjNGcKX/8BVTARP+rG0Sz1ijUETJfY2Nn1yMC4JYumWB/Z
jvRF4G7szh6DprTLL/THQNreKPigoDZjzAszpD7WwnnV48fe8HTqu6ku4Jyj4HRvTYiJv2ZBsUOb
cRSV70a3z0SgpCxVX6S12SB/VRcdfVtYBiKTQc17aGOG+gWuKgdv2k0M/iQ/kTkWpzY91GDa7RZ0
VDBHHMIAvHUwa3mvxHrQ/OlFshMC5BEkRQuVD3bDiyDv/sptBui7IguvxL6BwRKp/peboPjpJRrF
Tg60GjutZqdU0ZskUmnkZXZbgInTfl0RECDX7g68Qd9+Glke4om3hqdwxlvkpfnr/yL5WXPONZ7h
1ym2PjFzj0f+2GDstt3vGeoz0RHzW3jxKbCTKT2yIzHlQYkj2FUEsjw7yojduD6LpZk91qO00SnI
Eh5qzzvVfPvyJqJQKkCeTd52ce/P99cum5CHt6OXTZyluQUKiMmlPp9yZETyXldlJqR0Lc4PkewF
lO0L7Djao4G03ubldAPRv/NYS0wQHsFqXRL64Vo+17npqMTeUnZHu7PRT3/jHP9CJ5XWBo1u84Lm
O99SiXUyiAGKjbxFus6ZznvpNLso9GQB9I2d98tS9VOL9VSjsyIC6cgsZRDHAWcfqSr39PKfOyxQ
AZaWogKmZ9kr6DEkkC2eu8LS8l/Up1hlYsk6kJz1dAzStmGYZ5snG70+9kHZ++M9bW9inXXNjmg9
4zRFalNeBP3CabRO7OGq5OD82QwseUGDOAYK7Jmw05ulcd+aDWpqrjaWI2WPwuwn6dzkRVX0Q5vY
5Gsx8Dv0KShnH3Kp5cfb8lLfGnfmGVFJBEWrYc91XKELRn6/Zt2buNFNxQlEtW9d2Dnp3/BBzH7D
diQVd5TZcMhazakYcq5QaU9oH9dbNra623Lhbg3CQSvv5jXoPoGOokIx1eGHci+V+3GG67jKFYIX
YxjkGpYNJgce0jF1YURVq/1UUSN75D0P23e/xTdjgqj9SH5uMyh+q6UsOBJKD5bggM0Yl36XZFOo
yPFnFzVWUbUZ9G8/Q7IM8zji32EelvQvKuF4F3hbhcR/bFC6opjiYxn4ARSf8JW6LEwDXm1Gi7qp
1N70CsxwSU4vzGX+JYBoRg/As44xVD7VOQLBFiNxPXfjgwnLMflz/ayUYHWH+H+D/HMqp0cUobTR
79OAqIBJTNcheIx04N8OudKvT+iyPzZI73tpyiUR0q7JlATRiM0nxvtPUfvweTuoslh1G4TlP1fV
a1GO5+5dja6zY8TD+QYZN8p08lSDd1bHoIhNmpfcYrU1I1fM4UG+JThdeYvuRNfe8qh2Svq4QldQ
KRhSnTiSHxX3eyJPwYqEiTt243ORv//LzIx27ZbiWtH+4JJBrYHVKPM7fckqSNToUn1af2rUY06I
CdPIqg5puaS9fsvLMWL1Blv1cxq2hgAkASbwcqIdOSLFfiQKLPSu1jlAIY6ZxrB/TmIkUcGFp9NW
edvHVeznaPWZH9H3DvnBn9nE3Sxs0THQPSCVPmTY1CScp6c7Pkm4k731r+9fkk6GLM+4KrUwWBCs
XCzh0UKGm4/K6tVxruI39bsX7t4cWqAy1dfDEEpNJsKLM46T5MJcMVUHwHDfc7RuOfhyJbib+q3G
dqyOmfekP+uxQZWUlTWoFQAV8tVIrKlinXWKnbGnag2kMMdzunK2bxPpQvMFs+N9T7nhsFaH0j7w
lR06yLTwxxklkfwzFlkQSqFKLT6kDAHsZfonBkM3acUgOjQTluOHJ37U3au7R5e0K80zne+2mTgY
x5aEjmNVqYCQKlNOOeSM5rhU5jsyGQkwLo6gA7oGwYi/rHegimU8yAj4x6uZ++qi7h9bK6ftk2JP
6vg017YH8wOeGCs8cA4qSvE89qrRmWDgL0V4XfiGTT58l14sDt9dfn+QlZkyoKfSbiQ2jCanerxJ
2Imd05yiPX9tOyjwStpQbCT1DqHxeXHvtpasfDGHtgjjwvNEJUIbas9JJ5342f31OxOhRGxW7rzP
4EfqnKDpHoJJs/bMjXbRJRGfo0ykMayT702tHcXzItjz9iUUjMVPS+OsAgQTLLiplZr6JFlXFLH8
OZHR2PJKeyuq4rukWc8+n9fKHTZRk9inmmWoYd3M43b5kuGsfERa1k/f/q+HheuH5nqAZdGr4HXx
/wnZMBVJbcjtmoeOXWm4GXmYrcwagiIODioMRo0lhLWcRyOFZJeQDsdrx/oK33thmgiLDPVG58sK
2XxwgBsEPGs/K6+F6IBRe7Nti24tBetQXp6EgpyUPPG0G8H0DceynoeTRyazl7a4B0xuDdaM2vTm
UbBFthrlik5AjMOzVQRlsPUulZl6zoeLsWAUz0fyST1WVToTxUyimVLWzsSTjWjRctRlE091dkPj
wts2cnJMDn/hXTmYRgNyD07CPsoJ4Et6GUwP2GBG2q8lExl3xNvF30+TQT1bAVhMUj7E2hZwaxrs
so991KhYK0X6yjPlZQqEMzfc+4PDfI4M/nQkginKx/+I3JrxwRXsssNyqKNj+Dtj9uzc7rjkA3y3
olPnsfhbAO1XOdegFN7q6hTbzQ/0M8RrbTZiJn9ZZxrAKCq74gNjRG5lRosFwNS9eoZxa6NhCvKT
s6UJT7eP2ImvgG19xFYM3jziSTkNJ7g6+cX2WiAbWo8qiaKbrodrKDiBuPp6hmtu2X03fbe5+6vm
tVLx4WNyA57HMLRS8xcmat7vA8TwUBdtkEnjp5NA00wl9O0pk18m7rg2U+JMXlNzgJt+jBg5toUD
+dOZ30t6gqnW6H484nBXJbOkDxLRp4cemU/eLlhAI7BYQHoWYK8DYl8zpC0Y1D1hc5sl0lhhRGxY
bOi77VrQ3eVM8NtRze3n/T2nGNovSNnYHdU6Pkd1ppOYydkJiC/ivr8B0PRUAoSvH+M2t2fepTea
2+xB/Zwd/3b+rMMbhITvRR+aFwMTKJeGWaH1dKDQWCb7IFgIytlGmAk3pF1qHCEI0Qrq2UBFs4yZ
lesMDSVqS15jOQgh6cXzdX9Mou27uc5JZpmwTqkKj8wxl1Fpc2Wj8QO0wUBdA4LcsduRXBdi9049
tmc60/fEXZBjwcDhJdUtdeXjcPSibJ1l4JHIUlyuRQGqXnUsEwOgmK2NrSouZfTtpAIZI33ckhae
O11BmZZOqzRsxnftGwG/VxNtJkXpj7rJ0YZRCo3C6vmKeLiRToXme5J7DSkD9CgWzDXz4fv6LXIp
EpmUTZdDj3J/k4gp04dya490qsHTBoAk02pzg/IpBjVEduMmmy7aAoXuRARDEW7odc6m5ZeKOvH3
blPj7dtGYB3E40ZWj18lWKzrIp2UlW5i5GBChd54vh3gYNr4nIlWurS5L74vzKCqZs0WO7MH6E+U
EOhDlNOGQfamxybUabTJh0VskfTabr8Fee/X7ShyndB14JjVbfT4IPlzbI19hkpMykJGA0ff0ukI
Jh6uxod/zPhoGDILidw0ezoivwbKW3EOxB/uDAgtogQ7Ml04XQOeRYKSf7+Keez4ZKWdzjFGea1z
SeaIaAMHGr0p7kaqx+K5xVo+ScIQ3otlES6S3QkyWED/YLLa3iY4HkqZ/VmfJA5yyXA+EpLCefhd
oZtWL2Sgo5Sbxq6/dxC01cnkw5rnCxZsAEywfLx3XA/F9vNR3B/CjCIYxjO4OYRY0WivmSQaXR9I
JezfNkU/fM3n8FYqcvfT4YD2h017BA4ctqAi1QkQO8W9dHuRO5ONEapY96PucT+7IPlAbdr7MFsx
UborJFRTKww29Cjvo9z9Ngo+6BgQErZtWQkJEVRRsfFW1Kuf+MkecCWnRcdAZLn77Jw2EVPi67rJ
/Mma5Zf9fQyDNonAK9HZf2CdlZ+O/viWNzYR9rEsvWWawIKlThNVohAB9B3lGV8fdKftaR74Jn7v
7s93iHC5+katOHWycjcg5hFjIZ9erO+ssAQh8lwjxYSGxu+Nm1vwma93MsNVq6GA70Xs5QGglgT9
dYUMz3yFLDmeA7jzqK+cPcmb6ywog4As8w7k2dwZUTJIa4F/739KG3zMLQ45PzrD9Ure9mh4Ex6J
5nfo9JTAvC4b5B6xDG4FJMkooal9Z+wFfbXdpxGokgKFpaEvSYqoT7qAs7SXu0KXxkfdHFm/jy/s
htlaM6arQ4JUP05FYJZna7zPfl2vEf6VI3zYhvh4a2N1KBqAiPs1xVFNkk+w4/n0nTTLFYS3Me5o
MqKaiL30Zb82ruZUZnMB51+LICK0MlJeFwtkr8yzOU8NxEanVlXfIX10sRmbM6FMmxsFlW7pnzRl
O/00jMZIfmAHNDPQon2GMp4FdxXFr5sSMseknG4QDtM+Izpz52vi3O/se8Pvt1DjRVjK52f6ceOP
no+wO/UwjS43D8m98BTpVKEbDWbECjFyDxuemjLFtz+vnMVBVj72eUxNmYVvodSyYMfJF6fb1x5X
2UgeAYdE7mjR+PUTKMXCVyagVHonJxU+eQUnxTxM+kyHxtQXEh1QxaI3RYuOEMJCA/fQ/UHvQ8MW
4BnHYbbHaQcwfTwvCAP41KEzxs5kZcoUD9lo2A2SmZta/Tb2ShlMo6kS9t42poQhm0eYge5wb3gd
SJOjmlA9yjTiSzZw6b923m1GbvQwtAthDgQ4MB4Psd6U1dcb6x6N9hoqBh+XaVtV0Q7BwTnEFTS2
gF36saobZemfYAXY+bEE2DUN2iaScNReG6kWqqwUtew4zDrGa0sAzH1XaY80PacqG/0XL1Wb5vlo
WNfKeWbOkZ2K05NZFceEXx08jXWsiE+KXyEIyvieKYUBNEyeSMs6ZTN417GQq9njh4IGkgxzxIL0
sYdBFH3wo6CFcKwz3kly5XD+UGKEu3sgL/M5riQsxE/jfdejgheGrVnzDfX9qEN3rbWWFDGnUK4a
LW27AX9JLL/3caxwZqMUOlyLay11yXcLJP8FUNmIlLVt4bSiNKxnSAJ1iB9SZp328cMUPP0AUnu3
Nv/gfdKYDpcDOWauhJ/LRqZ8iOFqMcQCY4RSbuTBa0IZnPywKrG2Xk28VqRPT4Mqb34GQ6du0kcf
MnsiHWMVCQLfu8jFQgXZrtavs0vXx3u8f0pYMWrb9sBUBd6Cw/vs5vdZgemO6XuWZt5yCNC2K7zo
8o/U4wzaW3F+ZHVr3hC7zk18hQRMyIf0yChyO0/8bxMHZTx6dvAkHYZCW3qfnxJpWCPbR2c/k46q
wt2ppheVwmp5P9r3kVYYnNX48YS0HRrdOSUBc3HKrSJjSqbAqM6rN+wKzuZbf48WKI8KpHMSn9fP
LssTsZhvFWpzBQq1/RGwTZOH+iVfVoQpEee320EQog7SJu82DBpZ/Ufidt6wMA2R9LuaQRMc3UTY
8VuyJblkBPUR75oFedh3Lmrt7TJLxZ06ppDdioYwy6YbwFNcg2DPUEq7x0vaQf5nTgLNxtf1szKP
HE9cZlat76FsIzsdMRhgaINAmpYfo7edNRWVmtmfZJh675alJpFHOLSKPeeBKLmi22azomXlEa0Q
gyFj/sXDx3kkv98tvZm9r8WKgEMylqhu7zqffsBaHUaIAekEDn8QbhOFobgWYiJI+CpgzqVSDVaz
QbM5szeet5evfSfpvpq2HnQ5jlsy8r09EMYhxvFpCJJ6NYpWl6wjbedD4xDmO2HE7cKbqWli1uX7
d7yquMFMLdh7M/PMj4FUphHbXC3X4I7YqK0pwJP53kjcR3DDHvp7eqmXr4Vkz6Zjcl3HtHe6F1Tp
J8F7VgmvnRFLdQEcnSK0uFsMTO1wezuOV0nkJwqQsTDAFPqVoAgGFAd7Bq4s0DaVTNZ8ftKWJbE0
79I/V499H7KAw7qxpB0vINGsrg/OpGJXa46FL8eoBiEEaEuL2XJmHl4PBZVooviO9393gCFGzKSf
c0vdnPh4DSz2DAYE9jmHDRqvmEyuy73D7Vx25Ge7IZ6JX9IpIvMo8OLHfQziqdmLZJBF4SyJSjhg
5znTb44+SDbU7C2kOjtPrCrpCQvdHZPVqbbHsKaTsbdRZn1dvU4bCF3OhYCtmyC2Rw7E6lnAjO+D
MqrA/T2/wDUeRprA9slUuqBmwWIBf9r3bq4V+i+6uKaOUonW6e+SitlWfLCjzPi5dYUS2D2IWOS3
4Oh93WCxWyxsfsgzr7TA1trVvnBT1ytrveGaWEiMUgQ7/uXIioTdbia4IyssAYt4djmdm5w108O6
aBcbb6EfFaCGAxyzmS45vbosfS6t34aTBkdp9ln2IAQOJyigtJvSE+wtLDjGEA1pommbVC0XQQNQ
JtM/eQk8RerEdGPMIMMVFD6HCLHoYrEouPfecGZJU6pnBMvMvRMNzQY+NiAcmGDjojwQDbMkFK0b
GH3gKaB2VcNbfIH+8aP5pBH6YIPXnt5+X3qJvE4azhgzRuMvf6wMKfIiE20NJgyRtMoFP4zm75mM
1mR0LHTKmbokuTZH+2IF2uWYXpwDicbs1wWa83tSisaWpbwdNPMOCr27uX+bV0aiij4EJnJWS7EN
cKCHn4XD1RzfzChwujkWEaAsa8eAVXbvT2YZGdkMEBJTN6JLyzuZHgWjYOAht/BbjTSuESfnE9yM
PQVS6oGs8FBQ+14pPK42j4Ha5/dI1PLuFqQ94t3BntG7NMYJ+DLLSE0Buf/l05hyYGUVtMr6sVGl
AE8OWEXjJS7D3+/FRhvwiIbdww014tc+Ebv4cHb9sHfsf4ypOjIVgWzDWoe01oFGQaSxCK/+Kof5
UBJiILz94BGmqXzlGrOyunIEr0vV4NCChUT8IMIxz8TRFpR0bCroACxQwil/wnVlqDhFMD7SO7Xi
Bebb0OLT2BgrXMYhJ18GtQZaGxtrA5vCD0FRCn5O7SM4vlh05gG37AYWRr1ezKlANTTtlLwEJ833
E4Y4IJ4h1uaYojY0aeZiy8lyDVPOyuhF8MAzkAEqztEaYNGwh0r+6jn0Hq2F0N1LlZ+GaP0/T4f8
Op+5PZNuxzGxIBJQrM4zeYjSx5g/pMM8iNETSjADJWrzIW6EvTeXhwO82wagq4yUryUBG9q+61V+
PySJwY6INhPtoGsI75k2bwdZ4riAIbp615bsVU6zXQpoWIOjEgD5o+6JZeKcN9F6z/RvwJsk2KMT
cevHKI5g4BrytlQMzV4DUOWnJ0TESn9hLjC+oorEqTLQoab5Xn9Rt6O1BXV3mRwBfJLnzbprZ92v
zLNaky8UMk+DscFIHY4cTP7v0O1hLin2lPQI+I197WlrXtpkvzPFDRjVgE9SIq5sCesZgQLFrHKK
K3j6rn29rJVVBQmbzZf1gGFeMUcNOgx8bWpXZNX3RBek7U5i6Diml2LznkZE0yD1lTodARpQaL1W
lW/bFB1M5Nb5u5igju19ogs5UMEPxnHiObFifyvNsongXcTDpAOVSLc/ZII/CL1ez7NdXBVkOTBi
4et8BK+kVJxGoBr171S5bkAcf8vFbnLzgbUQ6er2nGVZqucAFTyR2XIzfCi/GV03YQHXhuDvoCXo
9nc7Pf5mEvEYtPRVBLbGB1soUE1ZeE8NXNpYjLGMUMktoEIvlDz0NzsSsNaq2NArHJQIJDsRlaVL
tIDCq0nYyVP3UZX7JHZf1W3qFQ0kDcM/+7TLiXzmGvpatW38hFDo9hdpVtMzU8BMjsRacNQRVNPB
zwhmmm66VvuJkbs9fETivPgTJSg9w8sHFjnAvORbT5FEIKo2uF2N6+UJA3Bttgzeu1QtYGMaZS1p
lZLi7VqsHNBXj5oTXsSbJufLe+/TE2FKTjvcU1nNuOfqugv5hBWGZWULhPIFRUxiRISgbJSE7K1Z
xr6jjI8KL0LK/VHK/TJwJlpUOyH7EdrFxQ8r36TDJtYJvS7kfy1ZBPYNvjYIyoDON8l1koHZaPWG
rHvDUgGXsoErVQ5R7z4jbL3G75wMmqyFkQ8fVNPaBY3Rw7Xz5a9hrzM9v965q9uZ/wTLpyO26+7q
sjnqf0B2LmEiI5GzNk1+kQqHqQ2+IZ9p5nKQQMhsQgjqL9VxQCFET4bkRquU353L5mhs4wZ3lNdB
G9AxtZLdpnPEJi3slmTxZ76zvgLDle9gseu8We+uPdzbqaghtym4/3pJ7Iy7j46zzFTLNY5FIaro
aWb9VaP8bEUXxq9A0h47eVXoLNIq4NgeXRMzJvXMvDGVUoizYWjLVEso+2F1TrDyDRk+P0uHabY0
Ya1hyLEiVos36kXBSAa7k95hoLci8Vq48hUXd2nrWACaDQonfjD/DEgvSrchody6lIk97+Cyxiud
clWmoYUPHK3ll68DbQOYyiXQgXFAKEgKP4n+bPNCaHUOQNiTgc7xbdZ9chPUWUlPovN8uqVk7oTr
Nx0OKRU06gFG7BUxBkr+Ux6okqhRDGVzDh4SmVWWBr78Fh8Vlh1T/CyrvO4SQLoibQ0w2YhTw/iI
1Cw6VXaQSXkxP6AE/9liiRjJh1zCw9Wjk8eS4nLfrncX1AqIpcZpnyd7lfnghSj0tva8sxtuP9kk
nky2so+I5VQuwXAj0AFUkYIkz/fVW/v+rKTX9po5sONWuaVulXQ7dQ9xlVQ8yZU6MQVN4NRovApo
fXeDhfG/rgsq9FsAG6zux8c8yOH9cekV3+6cZFR0K5oKUIAkgX0+yLy1e+RuwkUEOy1qQz/28SlU
nVhDIwuqDAsrOaWVkg8+lT9ds0fbKPx9qjRlHKsjgdRsoIeUOWeRGeHbL/Rc6xDj7A0y0565X82d
yodgTZEWnsuLeNgsztWWrh2+deKV3DMaq/jwXHiDzCszGSyuWgG8T1T23QVRoLFBkHX5040AIefs
ltK6mjc/2QaP0k0iBcikRpoXFauMvbWjEhwhJpg8CmrBGEX7rjHzzFWaU103c/io59cBgq8sszhm
bwKcfsZHGkexO9NgDmkcYiB6jxQKdHdemcGkOVTmTj/kCzWvPut8XVQEBThF0tnyVyxGCv0vSzt7
pYtsviJIpxx/p69gy8rShw3fP0fGtd08bwb33mR3xsffI3U3T7eXHG+j+EkwIHv2c/sMJExGfQQ2
UNW7lGY6aDn9foYDFLexE38AFd1FR7a5ozlGJ6MgcWAzYSeOl/UN+BcUE+GU45g8z+q1C/ez55bc
YTqLXmh5+7pGah0+wZ8aG45uoQQ3pwiDwM3RTZlXYk7jXMXu9PB6uY4r7S7uVS0N1Wwyd44qFSij
gl3HLo3/mCQRZuzVw3+8knDsUqPzmd+z0msAqbKkIDk8T/xDjrU6YnKTSMmAFwe788q8Vqw0MDHr
0g5Lf7/Jfs+Q5aa+ZFVe0vIaugHeVSW3F8ICTzkiMZUPu4Qf/6cUKdruHGOXpHXOgDYMdTnG9hpj
SdkU58eDM2wlPePm/uRnulQoZyp+a5fOLJyE7fQJg9dnWq8Td7NS1fW5WGZvM09Rt9meV7Igifcj
u5CmWRHcY88H0SfDrj0c3Tfj8bHXLq9vu+2jwPfBKxWZzTBPInZCeTNWu7WRTa1Y5yCfHlqtypD9
s9pMqmt7j2KLvvmmoyYDSZozHAkRRev8lo+CeBxYjBWEZ/WgdMtNQbUI5CcRu5kbkZWuG1iIaIdd
m2G5XvClcmvCEwdBV/0vMHqjbL4CAav/D1LATUlSL8XQph68yQdzdKA7RCTUpPtNZfgyr+uiMySo
7s3D+k8w8FEv8spD63Xp3symATaYrm9qD0ARhr5kv3nmd938hCLCcjmtJXn00XaBME+lfXcxwwdg
CGsYwUnpnesp4zySETj4q2JUCZ9q0+tbnIU46HUtN16QAh+jEWOsH5j3KyB4SEbFPbqzgDh5cETV
6Qr6GdirIB+jFOIvI/kjCapxpVmZgzKnv1G8/5wtRiuc1bQSJofFYtLXva7+jUWW8gLzYqzZnUWm
mlc3HI9eV5iF46bEudHxzpLdf5NlMgTMVoHUZsLYtRclyQXJ3rFPhRp91zAdahCYGc9MTXDkRkk9
QlEgY+ArZn8RlMeOj3Tow6XI5nTo3KAJQLvwqgyOhZ23xMxQMEu/w9soNNGnjmrApBVY9tVz9+KU
/5S0yZCzp8oc3y/lTBAhQ/h8kY9SI1DLSZB2t7Bcr8CPD9C1JsQEi3jkaUuKnlVJfiELoeNB0ZeB
/960XV9y0xNiTt5V4D5D6Fjf4WxVSg0qfCzfe6xZzKe/oIfRkgRtGy249JKrdTeNDVIov8n0XWmG
82wnC6uHqveOA4SxRt8m4iuhegHdRy7rZ4bB9AqUqd5EechIwQdw6SyUklDgPo6YXDVeEiDX+0uP
lS+Z31Nno5VK2hOdcB89xQUWtYv2K1exd0PZW9OahST09+Wl+ZsM86tdg74X6Vwu5+bdKsicwfqj
JfAAnNx0PKpMMpc3pi1XhoFeSoK7t+9K22T4mieIU5O6e8T9vVFOaLQLboQTynpQlw7bXO6C+CCv
lk9fHPLZGW464M1kKVRLsZTCxWYkTW1BnXhyUYyvR6eYvS9mSKbwnTd2CAMzFI1+iufsHLZM6HrJ
TssNk71DGBf7Gs7a5hQujQx6enL/HpFiDiHv1+Qi6QRqgUzoXaB3/sYG7htV0yRgr5lFSEmzgscn
qPcmGZVj3Z5ExToFUHKSpABJwE/AaxtDKcU2xcQxzTBFCOvI04vEEvMD7qp02gt51F/HmI0DE6rQ
lpDhCIyJ/w2Uie1TEIZoS/LaqOEYlUXHumd0rVaY2jJ+FXfeUUC89gHdSp1Esdek2CS1Yeoi4mU+
eXLwvJS27utIG0ZVpCSp9s+hJ9i67w5QiG0Hg2EGF+2Dl1SLSSCybWMWMvXZ429FZCmHTa+wvOn1
xzftQB9pVjYUNzk2MAEbZ8VksKEA716wLSxMMET6auaZUBbAFR4yVtqPppVfVd18UabtGl2DY/qd
Ay13x3DnogA8VES4EziV5sZskE0O68sBenzxS1iEUU9Ct0DYg0xH1+hxRh+aFH43IGsT6yONc/JP
mJRdryHlGoVh955HyWs8EgJ59BPLbgyenT7RkhtOtMbMRH2Zq1vPIKESG+CVxmZ9XD1HBdGdK+69
hTT6YbPqQ1rfDoVapY9OPtaLA4YxmDnfpkgKovMY+iDmEl2Hh0l/VW0T35918JBR/GIC5mdutJnM
leItk/K1T2tUqL1PmKH/c+YBPF+C9hXuWStpBaaFMtK6p9Wa5Bim4ALKUS1QFYLpHO9PmWc0m3D2
4iSyH/SOYUDtmy31gQLUm2AiGSWKZ8DjgqCrAqul2oXLsH30JckFwcGPIgSMXkHz4/29Byv3V9mg
Evbg6mi2jV9j+DJ7APxlaggcxAHS6TXwPArjFGe/vuL4g5vp+p2UU6E/IjpI3zDBvWkNKrl3KMIb
Sq5Iy2E0jxWQutwqpzPxbuBUD9VCHtm5KR02KJ8Q9SNv5ygwZLZJebWR7hEmGJYEnPlUNsCN4BJB
VQBqjLj/mEihPYOfpyFEVPesTqFQiNenHPqdbyeYiXfIix9JzIby9WzsEcKLeTCgrl0YN7rWx76V
KZ/UtexUKrhaYtSXUOOpFyxeEP2XlTBfmT92cXqQjlnc7RKh6DuTFPeFWhK+Qj5pPryZDhRpEb7R
9rlI0GamowhM/q4+D1SnZd00kV3PuzbFTDs2z5ONRCJ+hwkafsMz4RQCwCULV8dwjnjnyS0+gEBQ
RY9ewNxhU8TtWOCEC0i67NPLa3bsG+9h/bVwvARUAaUDMnqLQEe3kE5r9OX+ySEPKr3Ad0G32ZYf
W5ccvgEW5pPdNULGpTrnlEGRTHz/BTEqB25fHhC7bK5ptxMkdiJklVDWN9jAR0KcqPt+KTo8vqmX
5ExwH/lRKLAytrri/QD0KoATWuf94W6Guco6Ejf8HXsw1s6cTmTHuOwM9SDmiFDuMawQi+I5naDq
cV1c2dm0nmM/G8/+lOWV74NbV2hkMcURAjwi5MwNHjDnAEkag+dyydT4d5T3bgrx0bRDRmWvmMhi
OL8ttpb5YTwLwAYXHIMarl1xAgbvQyPg+Mpb2bIkUXoCHG5Aj8bI0MtbcUkckqNYB4d33Pvn+fIm
aBjmTyYG6QTQq36xJ67Hv2asB2FpOIdre6NOM2lfoI2x1DX6cjNDJ59HlMT59G9C6kAkaqJ2RQTg
ra0CbQAf7pnHEoedJ6Q8WM2oUUuqkCxB9abX/IntckL43UVinh+tWP6BBwxYA75ALCFYpfA9Ig46
nJHezodFggTQ0DVn3DVHMACrGU4u5n4K5FRo3ES+ZQPh5fEEElHjf/RscZ2gEV9mEDT3Hj28l9Q/
gqp7rda50eOreKNYfcr2/d+s04vW+8XIPxYnSno1fwc4jAkgvy/BJT4fnZRbSVsyfqMWGWswWcgy
1f5FFsfmtyUFuPDF6ImNhSIkhqJ7NyiQJSRQL4VHwTq7bVbFFS4s3r7nZBW3DOct2OVXwvx2UM/x
PKOVIbFhtEJOgR9m+rpW9IbWHuCxQzJznQ85C6A4lAAAHf4Ui0ZsTGiqgZBcMabbJ0l+GEa+LCbU
yE07IxfTNN01jPTAbORfvbEnOobSOmoJJyPx3YVROT4RHzXnhYXk0juQq78QXiAD2GHOLDCyYCJd
VObLmnbuy35K8idIdNtUfnrOCRQ+18aRPVMQl1uGgvCnQNoPbYVTuYmWPktxtBlGyoKb//ur3MhT
OQVRCmam/mowzAo+tL64YjQoED5uYWJVAuwIUV1d4HACXaO82on/5kjygoK1IZe3r8QT9SN9FOAo
iLPV9rCG7plYOJbvgP4Jv67mV2Io/2ZK4mFS1E+wryOf5WnOi2HlB3g5PHEBe1Is31nTVCKNINdp
v1geb/Pg14T2+5Zq8H77BpdmpGwNqxfKX6eB8fLNQsKF2giiht2Ce1+eh2tROFzN0Z4G6RGbfJoH
Er9jL5pk4e0IbJ045h7UB5EPLM1GpcyUsbIRc30OK8c9wPGe09PT2h0J+q+H3yiXgIijW8VRT2n/
wU0nUd0x1+nSv10lcfn45MK1SnnCFpepxuCzj1DH+/+sRoyqi+34G2WDsNVhQbuvhsmxBvYWq36u
KtiM3nM4sM9LIZVEIIdZcaznYHktblG7yaDxgXp895nK34kotALL1OMmzvcztPym/7S92cRKhWLF
z03td67A4Ky4tup/8lI/4oVKJ6ZWiS77UNjBpJHiI7wHH1CuAkId2q2mLr8WjqzZn8A2x0FhkChN
kt73WTQqnZu29db2foZX2Na/DjZwzyoy1KLMknc8j8nZRGmJQn2NY9hAogfIzV2o1P/GT35YLcZ+
r0B5sRZYqdaLMzF2L1MkhIuJ8R8OCX4TZ0wRkLcamiSRrZLOwY3jixuk5dlX6irXQmk5T2TJ+ELL
iuM+XnbTOedBSXLIm5a0eAwDXsUo/aVh3Odr5gC7l4D8c6N7jre0I4k2M3UjHVI9jsR+so4LrskD
cJUZX9BGRr130kTO4GH2j7rqDBxVdctoOEAFRY1N0/XQXc6apxJ43ORuEACP3THS3exll9+NrKjA
mdbiV7isTUTE2EmRBteC8SLD/ipYrMY/K88MnjYwVMqrelIkzUVrKWyTVmHiN6zP+FVt3MkIa8FC
Vm6Jl6v156qP3XfBMfMJ/pWOvoxgi9aRBa0cNbdBK9WEsNvM7xabIrfSyJVIqkZVhlva8SmW1qh9
RQinc7PwdP8/TUhug8jQbHnMaXIQ1zmMK1NnqQrGDRJzn+BlxTOzpRzdjblXkpxS3hneR/fdXlRr
PQlmhadh+vXjZlDGbI3hpOpwJki8pSF11QSkYXcdunJuUbLdAI+tgDd+9YdTY+Yqfl/FdaM0Oxfn
U3YOysthbbb2zkkKj9U/ZXSC5Msv1O4q9n5FdH+tpuSvjEgpeuAhJe9DLWBoNQ6F0wE59nB/XSTZ
sKAIYMwrZ9kWzpAeENRSmeCsRIQo9EWlSnZ/fMt7rxKjq4hjdrqQpUtqQfhcHnLTviwJQawpYcgj
BX1LMmRTYaQtZkWtFtoWXTCbjvf+G7zanC7DJG9P4B4W7RjSISmbTCmzechjQJGotkZoScRoeUoh
wfjtlREOG1i51netEmI3K34pl5MhTcIK/oKcTSxmH6H9BF19rnZYaiEAHUrH43sUtL744cDmtqFk
8cufPhlbA8MBAh6qp9ENxX+36uE9a4+/Jbk2KQC08HI54u6jB5f1uzlZqZRuOyLcUA0VM02izF1f
kv0yoox7DetOUl0B5zmoPbGn5fYuhwDI/KZ3H8MTSuQUCzOCSkDZrElcHpzr9CRBs7qyk7DKIfa8
gu7pm3qsa8garA7X0VJ1GQIhTxWmEUDwlFRGSXse0QbZ3ybCsIETbdWhBvWi/Sc4AO5A5s+1+9Kx
QqJ120ZW/U0iVRd4GsqI4ubQMt4C+Jmi0KeaRICKEAWZ11bYUfiJ1cdZtWqT+98pVjbrVFzPP3Nr
Apt2g+E3uHAxb27pkUWTTz1YJCy0C/8C4sJIT6v3I/HJDPThkqw8QNO2SbzKZpAs3c+TsnUllrus
VnJPaKgcnBDC9CC9cydWpITYK+/LqwcYSQD+V7AfhfseRCxmLS/OsQ97+EEBER4DVpi6HhPLQ7hT
mkSvy4PAkXjtwPO24aC3J51uUwdpCuJ/fn5V9rfhrB2Ppil6s/OjFB8TztIYvO9nBgIbB3aIeNKt
jxKQXVwMf59a8IsvJ5ut5uyvm1oxpWOouBT1DaSvD6+Aq1FjiATJuqCBanlGDNfsiv7q3l+UQP08
anxxee24tEFAT366h5u+icQctWKP8YFoVz7Bd+PrUSxA0bcFJHOypXhqhsFax3fjo/rQja844L8Z
dRF+sSOdqflntpHf6SRCyGRN/1QU3QwcAr6xR+wit9ZoQolxiGoxoO2bPtkVC1w13jzAdCN0giDw
xQUHyncjIgUHWxzG4K7Rww7pcIbfU5asqGWudmbDE8Uc6JR5OWiXOCRc4D/b1NijdLqyzQNnWJ97
wui48h1mlDTN6vQ2AC+LdBTSglhsJMnCJOZx7i6FhbFvvSctN0HP8/LtLyWV6a4v9bwvy8QOHOP4
RY0+RRHDLY25eDBHwF402AofrSCrn/FkfuVyQw9mhbnmaXusg5P2Vip7OFOJk9DaMUZbN5vfYVoh
j5Ke/3Utj5ajEkWuV64D5rIChMtjyqnqzYdTpC/ZDeN22aPJbrHJtg5IhYPlWMuCvPdywkm3xWJc
NlyH5B48x19cZkeUGYzDAFiEdA5bg0EQmsqK2yqkiHx81CrTPg2rDITQeLgZ9If4UgxcM8+7L1fY
g13+aKx76S72dsNrC3C9O7nEN9PUtH90gS5WXWt2etqqjMfoSXpqSpqVnKmm33kDx5ErCpK83VtN
cVo2Ss0FbTCX3vdeIMevHjd3yklVc9f8t/cw9epaOos4uT6+FVHKtN+cq//KkSt8i166pjQd4UkQ
pty7yx0h5yDNeavV+YjpuB1ZeUi46rdHJaEr4y/1nZaoiqG+N3VuD5Iow6Up++Tr9p7w4FTcD3Jm
7EuAAPCZj80mgJdIREU4F/qe/C/zIW4D2xn6ybehMloyxIU76gaVzXRnwACwLMx3chYSXlaKwaIt
ySAL4ACmYTZ/62nRNpB73mimlfM5eeeKrvZ1kHxMHe4gjr/9h0YvjL0zv+8oLOkMUUKJIqtEHRdt
opZXxXxxv2MqtbOHwFPhUFmVVWXqn82qGQlfvIxcHBFvPxRu6zC5kE/Vxgy7GPX4MUsgvj+F8/7E
44TtRCYDdt+EzB4vcqgDBLuQr1UO4//6TY6ANWfiyQ1r7cGRzeVyOaQHkRqaBLKhgAPvLl8gZJa5
gQclx0XJrTjTQN3py7s8z1R40Rs/PrhiV0GcXBF7o4vQk+ihz5kWm40HSjMo+WjzLvAWlZc2SKRH
dUPOSzSEF343eXN08Nx9mN5DirwkZQt7iZ4gwy+jr+33EGsFgxkr7QFauJgab7nHk8K48JwVLM9T
RtdAOmEcnf8luu3m+wr0d7UXNiCaSJ46k9sDNaO2BpvR8zCHdmGt2OxlczuuMCuLkHvCaClgbeis
IUkRMFB/uxL1BlJCVQKjfs+sKEzmwKvk0tRtlY6YnCkbnDCtnCP6CNOKpNI1TTP9CEi/UzA1nf7A
o3vmpzABlMSGqglpNZiupQNSU8k7J5LAEBIbFS2DFZgJ6Tt/qMxsFh41czz2m6Rsf/6Kr0QHiAl5
tUu8OyZlJKVQlhMnF/vZECIxO6BrYqm4u4eLCDO2H24B4f3czFDN/4Hsit4Qh5mJs65nWrGP2BN+
Jf1NyiRD56CG7a8CKjSTfQsFbD6e13k0M6ZqshejKL1qrNpKM+PALSsMx6DpJ5eR2QqVtHBNj8cc
yNDDR0Jf3yF/XlqQHgLyjtm5wwUcrC3geW45KOpFTwVZClYTCtIEalrAvBN4Gtf1YUR7sP4m2uAo
KyGtYTjdzqBV8+h/XGVjFphKAx1vl2J2IG0hZ7BA97czzYH3mhQP1/mjEFZscSNSdtJy0212Rl3e
FhaIeW1xw5ORjROQSHIfciiFweRmtadLWfYHf6YzUOU3XjPI5sviRxG0BXHk0AQ12qqZFrkR7yzI
v0+Wg6nySNg+zE+39uLpHsDCPxNgfK0yEWTWgLRU9YkdgCCAO8wvqMkQWGbsZSw2w9maYzYfV3+a
BL388WS1OnHvHUsLxAzU0JJ1pt4tMhwn49i8Er95H4OsMxcjhDIjahz9nomXd3NtZ6DS3fNdQc79
ctpn+Z15zBGG/3xaDIvdq36giYaCmguUKDnxPXlJDNeu+dDvqx4uX3ZuvX9OqDfKkHMDyVKtCsnF
JzmWgjyOCRRzOwPubPeg8Y3WC18TRTo138xo/vcRoic+s20vbpztmT+uZP//st+LA7nYMOwZkH3o
3m13BbbDBR2riPhPnXnEazhmCZJ2wybbG8ytqeFi1ZflT8vXS3Tp5Tuqebepq1PL6Cxxk02pinsJ
XxztGOyMCr8KQG9FUBws1ne2eDGczuu4Jn8VxKVsYJsAp2Zm92RA6RCPoUQdtjlWCUs4ccY+HsRC
0Zy4t8p3NVwFgGRaJFB5cbEgDvUdXA6fQH2wOf5nc1eH2EqS9oP+JLk67i7EISAo775l0Ym6RLSw
F55aHo6AAVHVzaW7dmlmKKvK61bHsPjBt4MxBD2z5Wze2trAlmb+SdCAG8ZGe89sAc4W80DNWTMU
PKuRBTqVqFOY2GGAbkXeLhn+jkXriU5XaAUlg3BXXeC4O+c+vrk/ENqHW6Ag6asAtdpIIRqbuXUF
fnpYUFNSfFDyxZMw2Pc37pa5snzsDCjY9HV0UOPK9qiXqDCyt3DG60bOEA5ik+raM8uAAzIEotxl
CyZ8JxguDR8gLqtIZNiXsi4wO3DZMWueIVTCaHz8HTxZ6s+vPYKoKo8vcenOjYjmlQ1m2gf7B0T/
aLyR0+jTu60TvRl5Gn05RCb6iDrElWmM3SAcbZpBkvtNGCPm9NLFQBtdrVZh7/VwnBkZ59QOvZ+k
okeGD87lwyJpHGu+xhDbaN3po764HaH16voYp3lcpViTokkIEPPVvu2p3nW7Kvi+2+gmaThO7bn2
96Tx4vLb9JdxfegJfknBIJtA88PexrlmkTQ6s/vpyuw3lIZC8E1zTPFkrzwTmTOYoqFetdge0EfP
cyOouRYIMQiRnLuUz2jD7gTma3JC5UL8L5LiZolAFIXacSLpZAuV5TP8XGZ97/m45XjOQT9DoLW6
OzqafekOhFMImBbo1yYPAAYEZJB4mnS3Tu7zcDw9ah3Z8Fa2bP/fAGMppGrldg0ThyXU4EblO/k1
MPw3Ape9toZFBr1Aukuywfbi+YIK0DjKGqiosXGV7LXytqR3f2kryUdpaHOK9GUkMVG78v1TILnO
zLc3h72j8yO8WXN2nyZHfSy6e5Y3whB5CZ9drFjZP7KzKxszO59MqR8N1oCVYt7o2T9O+ofZcxNN
awfnupbyiqeANa5B7VGc4CqsDHderFgeGtYx61hfUoYwv7Cm06LTIfm0tO+vWygJJWN6WUyi7vKG
ESKb8PNW1TXMhUttGNo+wu/5MVo1STa1JQEHw1FbpGoj8WJJr0OkCBsjG8BRi9kNUZIjXuiRm1BY
ZD3zA+WMzwOAn2XVEmxF0us1fNBomb9ZGs3Ot+Dx3V++kubDFC0kSeFIZw91I1Lm9+zOxiH3FscX
+ENqu2uqm04FSPWeCZrfvwz3SdGNNEwTuV3g2gbeG/uEmuW4W1uHA79NHV8ErIjnEijZJ2yFLk6S
15TzYF2m15ZZa4rxCk5FbEA0HfuigYesZiUWKJyN6LL5CKYtGW3+zqYtxmwUR7GbWUrUCCiBjdg/
9qxG2oHG7wnS8+mDZ4UNMv4Tmm+KNYk/dNF4E9ynAv2qYLzR5lZlefeClQMI6maBIeWYoOtht8B9
6LorhHUFKBQT4uwsHk7uKBf7wrXHAkB4hSjXOI4pSUVJw04TD3dDSlm0FHhQyLJ7ppr3hGdbckV6
UAoYw6VSCR/VXoxcn6cu5RU8fSX6Ttf+kEVn6Xx9BlgshJGlTOWWC5d0JaKvjCcs8RNT+BVET1Ek
y5gLKMBkJccNqdAfJGPjQvMBItjyRF3R4rQg5tl32EG6LkGEPCnPU/5wGcywKCMtEcVmIkOQr3is
Q4pCVf6mTrTS98dznbgvI9w6ETjLebOLDiv6XywXT1RTCJlXphlbWBIbE1e6HwxRDDg3n0QZ42Us
PhQRjTxA0oSgwIaNJZglyhvQ/BQQSiLdvM10RMBD+6n6kYOuMQFCgiyuiIF/ylaAQTC60MfOOEk9
TqVHbbpwuZxAVRs7sJp6mHPynDX5/FBSdtkNt5e2VzJtFArPpyjsQ+QWJ+82HeiQYPNGG/GFq/Q1
B1F8Ff3BvmKKIZ46lq4FHhfUG2BjHi9DXIkgqbaPzgOj1At9DPzSubwwQpVvRpM1IkRzuCH79H3e
vtB5lzq9H48v7HdPwPeNu68eZDfR3epUtyRw+RhHyX619nB9/3z4rceH1/SbvBOeFh/LKZ+ZvxrM
XcCqIBlliV2LqnAS41rcRWsQihxrKIFlAeW8+lA+RGLWA3p1TBQmfWt8QLDH1nJq5YLk/NitDO7T
5UzG/FDwxxvyfzihiV3lonyZCIOvydb2LERvU/P47Qmz/tWo2t3uGomVdpA0vwBXR9SdyydxWnX2
o0zLfL7if7+XAdmlqFoNOetAmrb0NG0NPaEPVTPHm/JAb6guUaNMs7/fBVNMzzGfd0fSxvCG+vWJ
SyhAhJxqNEb5u8PXQz3sYxlGQ+LSmo+YxnHkAKVJja9+45w03qVrqi/wquWRJXPIRvE5yLWLxmQf
yauhALoZax/7ro25G6nXR0k2MJG2DJ1PRHcWwK13Xr46M4tfI5GIhsvNaVKMPtsFJOfyU5VQ1pli
OeRpCceNzgYP6gBvaJqTqiSrUkyhjkE3rA7BHbhYmhwHrZOj7mdcyCR8F55FTgZb7N5It0qQW8wm
MWU2mkSLcXQrRe5EvgOWqEXgRRdTKpZW7W9c5yH7UZydHlK7KZuEzZEtGp2tUB7ib2nRqWAH5lhz
JY/M+z+nLjO71DRd4XmGLDaLOqdaUcSKKw8m44yvjbbaEafFam9lAdBYuK09QqjTzoAFDoJhyzyq
x5bY84P2+QPv616ITXp1sokOj1NrnuQ4/NXuWvxxkDAjog5Rc9o1jReu7inHphOFGo1lrMrJKEGn
IRYtNVtwxifEoDiH4+Xy4oOVtPjbjRUIUErUT1QKWTfByCzZPMy6nzQ73+39ipo1P2P7kbFjb004
g32oSTC/9kYzyxzwfCxJj359ejogwtUxKdnnXIzg6BRjSOteGznEFrQu+OoHMVlBpbwbzuNFKweO
09TE3LAF04mV3VrOXSGywcmEb34turrHm2B0IgCU7wRIKw+pL4itrWrNSMlL/Jrz2UgZABYBu1iS
VIPHkA0GNkGbFp9X4NdHDlukIH18P7AkrXVKWY1APKS1OAnuPr3TKrLBgUati8WcFZGi3ZY+6O0R
OF5nfbvpP87nDOEa1ZJI5WTIjdT6mCpvUadVEPKejsWXgKTx8pKO+Kt+5kDK2KUa5P0ZKG3UXoRq
cpk3hgrSJRLHRedgbHK0IkWp9grHqaCYAk+o8tv1vh9YDNKfjYYppqfsjEMQ9N2JS21bw9n5+uTa
A7Dmgqdv1SMG9BR4lF8eseuIQrA1ScIsk6MmYR9FHHDySbXxxgBVXnSvPLxWh8b8xhtxd1EHYMh4
eTw0I0MxUGwPSDbNLyK+x6e6B4ECgAQBCmIzimoewSDwM92j8dISkjCyndF5CpUyjq7GcTg4750+
Rw094v3lS/tOm5NOSpoTmNICU/fbffdPH3MouoLwYWSsQ7MOgvdTr2z4B146OHDi9lDruGRWDLSX
64WgRFm5i0ALRuGPRpUWNIAi/vssJC7EjpsyEZjTTmUZzYlXxMvrnKeZL/h+EXzPLnHBwut1dm76
qt+Nk6s3eykqub7Eatib+H7aDQZzfPvgLLo20+WsgQ8UWaUyX8WMzyPTVua6yjHpNnI0vuGMEVKG
1d0H8Ij8MysHeU14E5LRfzeP6uoHLB6vBkB9ajlKjFSMXy3Ox29M8pS1KzD8Qefm6jKcgdPxNXVA
yra8E+e8R4XlpXLeC3TNTgzSqGgx7vvqFwc42fdWLKfWmG+TQiitsk8axX6uilLD9ovavUU8tquY
2rg6Ex894ySafBVjkrjLftUs4AYJ6d+QC9p3c2EjNHLhMpYjD2LC17A0Ivz/RElHUGBj+Cra3eDB
kEQe4IaKQb+IrfqExM5tvKfwNrDv26YnPxFiZlWw7Q+DwNf08groQOqmruK0fyx2Fx58JsU6eSze
K55dCd7S/TmRwWfAspDjdLkDlbY1qcxqjnCE+pXwIDi+aTdNfvJm7H7y7QpCTP5stVv7ZH4P/yaW
WnkM/M3fQbZ82eDwz6CGb+BLK/siS2qXvPEDw5ec3rdHbxux2SCXLuRMN6hs2V/0C+6OYmGGfTOI
vGVJeFmuoU8o8mYLtfbbAy9yfAglpUbUsSzTfx5aFgK4HxOQ19AdfOl/YWNaWTetepBvweN0pnWb
FrPLkFYGtiUMfiRLmaYYsq7e/MkW8S1/0QbQvURM99NwjWKDmvShmIkJnOT2c/Qhe/IX6s0v9OHU
wHU1TyWmsbO3Ht4HqW4AIk+2EMquvxldpNQbtJpTAzaqZwYltDiL5nU0d8vqKASOVehASXDEyauI
OYPdAZ2vHARqNE0wg6xvcmrBPPI0D4niDLAWB0xMC6PTTXuZOuJnJsX3R9jI4ortWzUhVhv/Lb+S
JCvrkAZaJYmg298T3K6HGMD2usdNBDq1wLMDj3jAfVhP8tOU44IsntwuOSAKFOvgLAK5xCke+5V7
jKpxGr3Sk3eabhKYrr+4QnXNrzV0rcy9gkCGcqSR91K9dkeiCZ6k/WtwRphx+pB/e5pU6n4CPTyI
eAJN1hPAu5w+Kl4+CbpDKDJN6HZyNpggTtF7LxNzMjKihGLSBoDEcKzQoqNUagKDpX9nrgGQc33c
qELWxVGKR+7oZ5KwZUm912F330mio2ajREVTee9UFlm+CTCry+VhG1frGPX0dOhA+obNY7aXIyF7
qMgU1csTMKSaO/A/z74ru7n0FxHoDOQ75LK1NZjv3VWICHimkTYYa17/rRI/GN/at/3dIds0hflG
8ih1wIwS9fmqEJNGokn4hTd/RLSoxWjrZj93jaWcScTuHPOdfLcoeJb5iKG9H7W7ycBal3Ww9Qy5
gESrfZ1+8lpf1VAfo6hW/3zKhBnhjFSKOJSSLBNLSDXB5bjLQ/uRL+KXfe/BH1iTPeYOHG2gqRfM
AvZgL1CMmm5BB45+FVWQB+h9FqK5wIwN+oER98EyBwGfwCfYNK8nAVooYYxmerH9exOl2MwcXXot
dkPGON6SVu2DCKQ/VfMjU3ULraur9FBe21pXYX9H5kwE/QjLupiEI6FX2QVcYA0qnfigt9c5RFK0
y6obk4nMtw5bMG7F1E2E7UwiTTVLDpVMIWC8FF7jZV35CXJ1mv3gh7edIPC4I0OCK0y2jHfEWJD/
fyjEg/aL2cCVrNtkQ0dG8KA4yxlrhmadcUysvVdHzG3Ed+RGmwV/R5H7T7YJtOL0AXFacjo2wQgg
NuF4JiuoHPDBZ/rO6zesxwsdLUxxwauII28gsNqQKcpRG15ty6IqnNLQYmrJWClUvQRCi3HQ1NPY
AiA6lQjZSSPUvzOEuhgS+nxa7SFlGhrOM+dN7vVzLlHmVLIKV2/IzsTOU0fnkWuOKa1XrNFmBfmS
tp5+1/xvCMErhe1H4h2zbax8YDUbcGtXUB7zEUwc0CKVzJ4uz0x2aWHMjaVsqlczFsCSbYnQsPA/
1gJazuG7eljecqC/Wdq0HRWqaFxHbNpbQ7ZfRaU7dsWGq4HThvkybdMKN1nh+o/w6NNJ/TiAYsCW
flIGY6Q+SPaSkzIXE4T3aNCgvX5bebgQpfrWy7vV6Y2NwZROvIhqIs5Fhljt6gbukxIJYvQmCflM
8oKtOErg9CS2UtygzuZEVjXoq371HFLTgKUZ9TMdfS70A6C/R6DkV/p1OQIkmX0o2sATh7w8550J
4r0NI+WWg0lEgboQ+zDYAuN019HtKHJLNqUH5FMt7HtSrHdOkXRFNZu5i2R92E8DJC2WavvG0EkZ
wEXtJ+F1TeCxfX3unyiW/ya0yDVkGlp/pcPyX5iiJvgllJujPYVpNI2A/YCuFeh+QsxjVuEBguFf
p+3p68umf7fE3QLkD/JglKRBJZWb/vgApkL61mobmjMccQGBsmOYsJRsFPTt1HWPk1qchuau7W6V
OQKDnle8uyxYewrwW8KvulbTfBGuzIzVWmSgvKXKeSNrt51dcJ+U/VmhNMelxI9pDspCM8SDEb1e
WP9Ro5FtRu6GenBMNGKPNvkWesiK0uhDHvle47jPB7o9hVdepTRPwr0vtb3I7RiMuweqZjDP3Tqz
lLb850eLYhJoQll6O0dDSOP3IMPOOQeHAU8nUNGV6uGmBuZyeT5VaOklf4TRIjW8KxZJttXbl9El
xmTVyVomkX1aIcm47l+2I/jNKoikH49s+NdZ/5fDcq6ehwA3thSM7xFwl/lDtRX+4geFFbPLX4Us
KChiD6Bu1ACDz1yJekO/RO7ch8NTY9OYpuEK2zjvrt5umebgjWXEI0jC4fLAINCFKOUV9k5Rdi8L
xH9kSqCh/lF680rH2BEzpPRdNhuwqUnn9Cblv/ACP8eq90nKg8HIgugMlS/4AxP6+ckdGuxWbJva
t7TkZ9PT6Dl32IG33aKF66int3VnJ5wTx2FXWZ6VcR/Ln6oUZiOSlH2lX0SWQOEJeXfeMka136Gg
1JNsVjMtdpJS02ripr7RDLPVRmbkcwIN7ER/R/BRjyrzIW4CCEpV4zISz6D1bfDz8iFrxz2N+C0i
4JGx2RS/+XvRvE/lFc1n1d1WgUZF1u8Sr6O7pMIRGncgxz8NSiKEKKrjYyRNnabnHuucn6yDg/jp
ZM6dYd0xo+c+1C0Il0/e1vaJW49nuFETEqbyX1st7b7jBHhkwK/EncDApNwF2/xfMlx9/eoXH/JW
VD9WpXvvSrkKlS1fZWBg3sJT/y0jJFw3mzxsNaO8FahvGCfJ5J0CzbJkKvUMa3YwoUIWTXtc4aTS
PgmrA4cCKnHRcPTqyRLwx1xbKejT54pzZDq0NofF6J4zAutzqMuwC1PGjJhBeFNS6Z8rQ9sXSwLj
XuHKgpYYF/iq7FsssA6VP3nNejAfI0pV1XQSAgiDGKfZU6GC5FA+FdXcWnfuAVbVMN5pXUjU0hkB
wViTJJ7xGvVeyV+bKKwNSE8tZ991hEKSfduvK9j443gb/52ZdtvbgYQ9VuPM7s7x60OHyhzqDJG9
V5Js0RLWWZCcwbQZK3spym1mz99frVULdqzH8N8XatZDhGVwc6Xmj5fRcR8ISBmoTx1aLwaPz5iF
2jo4H8Eg5n6od8UOXRzyXNtgTUexJ+jDBOx5YvT5OX4WmfskQbX4ovi0rOLWFTZo2mqRRIpvjVfA
JykYi0JO/S4Lkv9e9vmGV/lA2tmS4kyEOC9fLmHG7C9ew+hrgHLHSCU9IfFaJFfHdxlUMzE+Tmjh
+Wzsw5L8GaPC383sVfPByeCUYtEcerVD8l1sywWb6iOH+0ZTzdBt1OSZdsOvjFlKWECk0/Dny8C2
JsxsZ+qGBghmZuDvr4bvTUftxr5dV5feIPWIo0qoQuHLhv1MfpJhdAtpgIPuU3rk57YlnMynhsnj
JYsuNiaubr7HXEZy1SnJZLJcXgn6UovtlXaJis8R+uAWQ6YEGypedHYc9Gazc5SBbrD1vL+kyem7
EUiW+IL9NiFl3NoPjvD33EJpNm3Xek98E08CCI+N8SwTo7FjP8Z6aoqL/lL54vBrBcX4Q0y238sp
mNdl27vtSz6gKVDtdcxcX4WBYmuzmOC5KwvSxo2Lf59TmccXGQ479ynId3Awcw2wZ7q0ZhMmldr0
56oQU9IAErMYWF8GuFDUFYgDEDKZAtvbL2tfF9U2OzryfIU2tBEewWgsr3z1ZBxCRLSzG6QUmMoX
e5QX10cKuUfIBvLhbGLA4GwDdnGYaxxt3X45YOINGIAkt1XDplVXzgjj+rHy8/4n5n1aUWywtORE
/vCU3Gf9/9C6CjcTdHQzuZvMvDEwn0ESrhu7Rq2Hw+7ADdhUbdLKnrZ+XjmnvrWCtlaVo61hzlE4
hB5tveRwCQG23eDXuIUsTggC+Bq3XvDqxGuv9ux/CccPbP1pkWwWls+cls33OGvJqb/QS0dB0JBE
uvrA6YNo5bGJUsfnW7i2SmzFUguU/7ZsZI5KsSXwkW102t4Dw/rRz6ZdBT9VTW6Kg9iJE7uCVJEK
PDgb1YxLKjMQC40WmjECfxZqmppRbvVtHGl/Xk2GlxruY7uixZK0JyskNZTDZ+HfOpSn5WljXyVw
toiPe0YThdAsLMtr+RsnYZ/1qEzPvqUxZsmAJ0awBrPNuCyL2sdbK0diWV0hBZQ6/l078K9Nl0Ys
F38ve+cpWRzali1MCz4nB/oaLW2sn68DQRIb+GUBxm9Xvpuy7xsVsml37qY0HVvdIfs0pvygRRnQ
a+KL+EhIaUvFBHhtgkMOUTptLvXrHwvSSVKJPBi1jSh8cZJIuhY+miuHtum2nGH0Ok6xN0sAJFB9
zX8w7+L+QVvxkssOHMU9w1BXCfYW3o5sbai5puMZoRePTEKa2lH2lxY4BJOcFuMed2DQvCGz8Xrg
2/3nUJBGCrJESROwg/tWQn0dnOlLK5pAaql5ogMsjvlJEkvv6nk0zq9V6CqbY+aH3+DBUuzkMOfB
nG43sXE+lZ2znkTZvco5bkrWmEQmpFUJtlDtXxDdj5jmz/67+q4Kf4/QxzUGb38oamN8ocESQOHa
Ki+1l8a+uop8F4LYd/Ac4lXmxv1+SczZKQGqiZ43XI40Xj/ipVDI42uXqvbbFVa0Z7PEoQZG66CQ
eMhjcpFXUMf6gg52s8xjhsgD0IS1HfVl2gIFrHHkSFti87hfzSZpJVi5GfnuFi8aWVdcc90R1K93
04EGUBzDbPaGkDyejlZU5loQK1RTn5P6eNzFsUyDoEuWLCddIEToVUcg6W2LcVDCsTJSbDwhNm0+
Sb3iNHc55Ms+eSx6Wainj3DPXJdKDOjpIvZ6C1+fZFTNoIheOQmHt57f69LimXSHWmBr6BZ0CYEL
Y/G24OHspcOjyfP8uAo+dYqD0KHVzGTokb0VCCDEcjPr19SOgyIK9Ba2x5guKc9L9ohCCRNWNEPA
2TIYbUThLKc7g1xv6oVSPQPhw/T1JvOARquWVUyDyWj2YiKeTQoSRvf0cgqTeyL4PQgu+cRdLK9m
F8U8I7PbKSMc5CMqeRnj65bkyu7U9p8bbyxXydHSOK66fumAoZa83KT7zzEvIKb3pq3eoAWBRZsa
ODAuyjqho/3JbRvYv/DrLADH6cQ1vM0Eb160c2tZJOeEKEPIXfwWLn9leJp+PnARpzNwJPQhl+iW
b07cWuHzI8SjD++KQ2P3zwXSP2kcCLDDdGTCNkLnQdQDV4w6a5cjWacDjuoltI9jYWvLoC6goSGk
WoxWWlcvY8lf5R17cjZ2rXsQp7K7CpxSHQzjH5NT3LXkgrMeHHGfGBO6E66DAWuDMoZvt7jkeRh/
g2R7AXyDXFihC4sSYQwegxe9/A696eCK7EPb/lx2rERAFuZU8iUjdQcONQ2suuqgV/eGFN2q+WmM
vb/Q1eKj/yODUlyRA0LhW0en9BCPpVcoGuUmUnfpakJProinuEEcgOaRGDFFUGv8AKa/Ogd0H9qr
SEvz1Gol80uB5mYKHnlXvlRtIB43QISJNnLIU1PAWiQrblffHOTKwejrKXDNwfbwF6jiCWOm4+Tc
+FQYSVItOCfXOF3pm4vvU4K1aUTi1GsngQT96T18t5E3gLzfTWLpkAqVSraZ3bzrC415UXwFnPeh
gW0d+CQFdf3Klw12fQ8fuFocPp5gRcts60MX+gtM9KRO8TeTMH/gcA052YzY2sMCZnyldkIeaMzv
DvcrelKpkGt0ilNYYg6FRaCYbSVWVnzsJH3crQm6JiMOVzUCY9/Fe5aM5njA9RTru7wEqKbg4sto
jDCEqLEYQwzJFIOqqTLbZ26v/0pgnRS1SgpI3hDfesvVb0OL8ghVIXGqyiYneoC7bBAcKax6TJba
bC5q18MudEXcL28dPPNxxHewgsF4T+D8p/nHc9saYxTFw3i26X5I+WblsSQFt6kWaz6ex8gGaSGu
sGZ2S/4UOdddeNwE2IHDglESmM+xnSPHImDFn89VUSmm57K2OgskTUC0uYbJ0SX4YgkwGVp0pYnb
DtsX6jeNS0O5AJBor3uQhcwfz8cL8j8PbN173/zKVagtITtwc7LnpeJjTOjcw6LcnZRIrTZ08iDS
kWtq8OIE2YonisCiGl3lcW8FVpQgFkPJ+7euyVQONJIJuWJAdsWtVD/ULGRw0D0UJvQzabqESZuu
aenrE373AFiWYMyw+au7WfJb/BAXJ6WF++PyWE/AH9i66Ee8lSMtLk2lfLZmfiZAzzhjXnhjwpXd
V1m2qpbFfx8PA7aM0Z+shnDKouFT2+i+03qx3TIsEVn6uA5YWOVetp2/4Xn50puIZyrAQFV8YyVK
Q3iQqhWzkOb3qWUjGRPD+9iS8MiNHMZu8MTQKWc4M6fIicWTweOJEV2qWpVSgRnClfPtH6KaR43K
qEZw5hNOM9f4s9G0VmuI8qiRkRwgLsi1uwFjNO/xzQlYDjOvdPS4EE7dzereD/l+l3fKYupDfLTc
Ih9zzXcPaOg/tum9A8ak8y/XFDOIageewNZ4heEJedWQRSjkF5lOyneBNw0mX7/OmjDAxJWqKK8U
8+Yz14/iLJdTJnR21BulJQgYIVDrQ9a8nRYrVQB5CKFydr65xQ/F5XrIB0g9yQibqinGbLexrm3f
CpqpHxRyOHPvWhrugSgJA853crZ/+dAn/0neXN7nm2qg/pljusbldPKK/pB2wNfMb3tsTu3XI6TK
Klz+PaBSQtLLecTkSmP2ZVXLhQU6qrGdSCMboe58/Np0CXk7g7Pqr/YZir9ZEijt3hEWXfhmG0gp
790sYG0FvVn+NFGLi/LcXK/vWd+FStVWNZ8lpjV6FzpRD9doUp7A3KoyfxMOGnzrtNTmkoRnBs+m
Ixs5gem0vRIiWW2okwEMxqX1Sk9EjXFP5apbvEJnv9Ytv+/di6O4POHr76L62/q4nU3I+lVZPwbH
L3CXQg47H7G9xirrJm5Z+CuMvgCC5GqlMNIh2d2r1Jk+PXlBdD4kHig9+IaXdIBoNj6rdvrC9QeG
t9iBH7hXvmodfvrK47b/pQxW2vnNqI/LCxMLqWAXVhO8T9oD3Dn2qZeQ2xc2O5re/ZZP7eOzx84X
nxrVfDH22G827iWWqA26uSts3UYbuU0Dn4q9zuQq1cH82Wazh7SQ9nJP5ZCmdYKJWLCQG0yKesVD
H3S5P4b9GA4UgZHkX398gbmP3XFseigt1yNA/o9+CMMyBKNjnEz5k0GAKc4/NxfKB+2fG6qkIU6f
J4YDdNDbAMZcxLZs31secoKUKyvSVAQZUQZNnLrDmxQ54abJ7+61xmhCQAU+m5Zw+nDekYRNLLkR
epPwnhypB24zqIe/Xh1Ff7NFYu6HBgYKe/4x5aUg+Qzc5yF17zLZchV4DIbO7mntTmH1BoSaOpTx
wPJnhWmNgsNzFHkA1yxan9cwJ1mggBrACYAqy01ggmZ+20NDTG2dlHis250QkTotG67PnUTpeNxv
UkCOZ5WokCnEx7MWuIx4zWeoOqu7s7IxkqdNhyHowwYcwZLbObYIlnoB5IdEX1Tmvt/2nJg8vKw3
wIffHhdUOn5tT4qMXeyVF2A6U/TNgWIv+CHiWJm6NWWgiWRfYU67Vf6+yshkok8KXuCr7kJBvvVT
pF6ktmBvpcr21jRW/6uS1Y3WsJNDmL1jScsI4udREDoR65VO4o8Wfc4692l2kuq6SYY6Q31ibhKK
2a752TOEwhabqogTmUqeFgtvLbBnw9jjjnfnyZQVxQ40VBGVFH9+vusz6ZL5X4SJMy4l56eQlCgm
drn+FQpS3jwHhp+rvoMnfwE+ufReDK/e99STskFjQw87/+ErFWY2mFm27YCRjPpJXyU/3ZgQP/U+
cbC2GsQH/BQR0mYChBf+vB/GpMWl84SKzyFbbTYkRjtM0eUUobz3jTXY8sPCaEJyoaUV3Z2O99d5
SOX2vM+ucbVDSxlkNDV3fn6WPG5SEXdhOrvG3pjXu0H4WLG8NODLTui9Nneia3pBWbaW7yAPyWqR
E8+SdaVUGCkswNXFuMf3XCpCvwQM2Kl61EKrzBsV6zdqUxl+gG+SxymP4oBRK9hBzVa6FQFraZzV
F0YzBLJphWQn7a9wUx2JnyZCRgQH/PGqKkkjVpuxv+2cChtRhJh/foFid1FT6RKcQfrA0UYL5Ql0
KXGAWjXKtSAAN5wVLFKLfQdzmex3Tq20QUBCCmvM8rYPTYW6Q6lstKShWdEuyU/TM6DKQYl+XvyZ
wf6aut//tid1bzjVeI3qSJy3teuG8v6z9rOf8of1/TkmHjj/bSFZBHslJ+R6UkSlPG5TsljzPiCL
idwWBYcK1bKdwq/U/JNqRqmfVFjVtvqO9bnomtrzdwequcSlACF/fI8YApf5rKhGtcyQp9QXeog3
bU7XIs0OUH/5oCzo4rZ4YCKN7XXH3wg8XqJX1B9QZBviPIFSjXwffxXXQrAIS6J0t3Iupw5OiRk4
h4BDSGuLQxp/ZGvMYHGEpgu3QtWR6H/OAWnYJwOM6U4zp3s9WVsQgXp/btIBWgMVSMZd8WLlZFI7
9FYvzd03lGX6MDXAUhN0wjWJCxijNkieZqnvbkO6Qv8Mb8LVOA24JEqQdi/sYcGxXu8K9ssOUZnV
CGYM0JLxEEjMexllWPTL30yi4UuBKoLHoR31yzumit+vrH4LuH8kCZJw3BwDzf075N+I1nlM4GDj
Na51aDIlQAQF3sZ3o/8ZqqjnvK5AHaqX9oG60XTGGjs5kh4Ey1JG7NkXuvWDyiqQMDtn7bmzlPMF
s/jVD63LCUuEAPigf7aBZT3ByB6B4ALoH2y+PjnIiJ+eNZMsP2j1iUxbOBsiQQ1hGrbqW1d6MHhK
ONg/sF/AcKg1W9d7uC5UkmICo5oiqROsCrrfkG+fRAjvOhOvqjuvSmCXeStnOuU3tf08NHp00c6u
48y6vQ9uuZlKs8/LLsvDFZkQasoRKUx7jCfNV+s8IhAranWLZPBM7jjMwcjtOzAmc8f37jaHainM
Vxji9O2XGWySforM78dp7D7uFAbQGIYZ1431blF1eSbPNOcfPDKzmprn40LM5TpPuQi8tMUXGKUN
z5Xnvx8V1B9FpIsGhq+5B+7y4T+93R8hg9zmCBXMjfA9zrkwYdSCkN7r726IiLufZ/FE5j0EElLb
31RB4kyypKYME8e+31S46q3Fp+kI/RrAuTGsDp0L8T5qU5oXrLngbdOQ07jR/19Lutic4B/FTNxF
icYXHoQBYMY1DPTRYDohhZkKQj4pSrBK29fwA3f54/og8/ns4Ko0AkZ/bgUp2NbfpTuJMnlKo0gB
VbgljkeU8rDgbBjQZGSqCsvU9Lgz2fp3ckRJzEORBlm+Vagew2UM3zTOEegAuPCVmEmFVgJvxD9w
YDhP40TPrIi+C5LX43iNrtqUgWQi8OuqSUg6oH/qSG74WmSjSxaUg9BsUQp6jgqjOOtVci7YI6BX
T0oF1zLg05OCstwILLXgAILIcUGD6KuVY60ZGEt1MhDhSF2TexoRGiNFuTzRUA2D1GG2JJiWiseR
BkAoTaRcAVSgFEoXJK2rFK8pt6Lw+GREy8xnGjlUUj15QPd2BUODxfk7EbNmhYOoE5v7vfFKEnjB
CphCYOy2ghrESCuFybomWOSFw0B2X7IgoWQuOrcLQ30WjJ2jI/Rt88tkac3sFvv3cvleLP/wThVG
vFsqbhXKakUu8qg6SxmmHjTndmcM8RhAo3nCZdfvVPLxX/H1H9wOVfQaf8HyJigfOhkehDqZ3KSs
9TPMsMGo9N+Nr67zeh+V0IwJM7WYbveipTChqCteeTvLu54DEv8gZ+vusvgXe8oFo2sNchCRN6CW
yJgao+nlKJnUz4uCe5TbIaf4uePzx9hEaTeiUXaAdXQxrYRj7AKRxGpPs2T4vcsMRjguBGRj69in
sFfa+7s+pa5CBq2uuJm2c/lf2vQkhjgdsTQJCvd/pl9z8hXt6YhnyU2iUySinpQPWOIQsFWnokKE
kvnzGZH7v6ghDw9l18sHhiNv2wKfHQTO1DBqVfA84k6W0SclN1nCPYu1W1hz9fidlaMAgzDDfp0y
BjrDHuD4NPAXoPTFfeVwXgfWlCbv5pgOTD8vJvSVTMRMoR/MAj4mnBNg65lVpoy/XnWoco9LHb9f
RI0+REbvWuY8+Pj0tivigvteNSwQvrQJf8hQdqjwJh93wbimAEjlMIFsOQjDiMZ5iC9IFvLHSsHn
jzX3XcRicihb0W96LAHPizaxgESoy8RzjU6aAVxqt3qyeURc0prpxaEHNIQ5jXLyzpGgY9RU7o0g
3TvPsuimbyVofSjsBLaDf1SdealHG8cJAcuMWpp5zJIzLgVkWC6Mz1Ruw5GfBm/twqTEN0bmWg+b
ILjr8HEEfBM/bjMI8wriwHG4MuZ0hN3y8IzR6aj8zZ1FNXoAlLe4CFWOaOhibyAgz/r1G512jBNF
/701XQzaaZxICQk/LWeZQ1WyGbzp1VEkTbP3/X0Mbtg7bqNCy0UBXw2lpIVmVUwhWc0I1QdOSglp
O3+sV2QL+Cxilurb7imKEnz6NYwcXwP8FGHVnCsRdCCk9UX1bPDoN/VjRjCEsWJ5iSUu9SCmIx/3
Os6+xl2N5BdZ2Q7mPH/3O3Sw2zqzu3hJOhVPeBqvmbdZHONUCCRFxbnvfr3kAxTYFdCktEDnRZVK
dFXqzffq3EigLhn2FVhm5g1PlHjhbNl7DmL3L4Eq4PsZZddDjmzfGduFRi+yNesSOhl0W7Stf77S
wDiTH7Vbj3MhMnkU2yuKXEcK6UQX9F/7fLM6520uSNk008yJO73K53dxqf/vb8MkuLBKnyEZRUuY
CGbD+UZObIxZXWljSNUH3H9kaNyEUSbcergZe8aPgtN1gCKaIlutwaiCIFhX8pIfxt7xIte6r/3g
vPgD9YuFGPuqmyoszqfd4mPDaiFunJRZnGpSnroiRC1nhkuen7+FUA5bIaqR+J9HuALH+3Vh3iK5
24zs+i21rXDDgFcmfBZsHdqXjLTbDNDqtspOaY83akBo3rGDtxJJNDQBXEz6PaWpovo8/MMgsBPm
3HPCqD8IZSJ/aR7qEbuZw2kGN62DRqW9uMfYM90+ewRze4+iFpLYasfAbp4FAMNRVMGfVd9PdV/3
qJRLi9IQPZ24zU0HeTCkY4jNIt14aYMrrew1cu1JxNYEjH9RtXC57Kk1HcfIySaveKyjV+fN879r
L3hYXJFuR+KXMj0345p189lGMDtMugwzeBmIQzjzgm06+ik4K/VtEQEOFXCFSse/PRDJKz+KV6jV
9OUXjsI87dHketdJ/8VUxWajpr9Kijf5DpGk+1bzpQLb+2O85I3OhlQGldTNWh/IUVn5OSTwRql4
kFCzJ9uv4OH8EbqxxyMWsWdlW1K39HZvG5QPeHSRcNEg8C6KtSMqfYWSRzPmigJ+RYAIciNPPddA
ff5LZDvXqnqe/CxmuRPChwS9FuLJoI3/8II5gVuyYHUmgw3T4S8519KLf1cUvEGH8L8baf1Pnes+
QZwL6i0rdM0hG/OLOAu6qfaXvJ5T0XClryUyxCvuKQTNTOxr/6o/5XMjDjORgYQbVEVTVClCooIj
6yGhJxaVZdqTpbOPoERtEv94vXSMjUv7h78re6a8VH5Dc4dnQR9uzrSC1EnUOlfcd0qA590SqCx4
Vr0Hd8FIF4hV/LTLAATg6chlBr5lOV2U74qp87eq9TncHmQMI4SCFf7q6dMqdtlBAz/GotDi8uWx
0imbRvhrLb8z/z8mHd7EVptwPPSKq4wkhszjX0XYydl1KjYINzP+RIRsbByWuvMsOhan2pT5kD8N
edpwuQW0p3O3tvsIDxdNF5LCdJfcLw7vLmB5bLG6l9JQ9Kc64F8JYAmB0dZCX/Iqty5I41uNKMSF
4u7BwRr5mEDf9MYtZo3W2s6w37d8G8nPiRcV4nFK+lvxoZ+DxPiOwzrnt2buBD9F1E+zRgApQ6QH
V0T+WhWVhuvW7p1RxsGACFPMunNtmPHKgpRF4t41EtBQwBkYOrrKU8I0w6q3kTwgQgDCcMnrFLWx
vVDEyjeyzteHlqOrx0qlQLPFRiYlTZh8Kw9obYJXbkpY+jGqQHXjokNI3ch9M6eiRWytAPnGAPbt
QIIVu9X0sxdpHOoVIcIyuBzlySvq8rUD2uylHvZQCPyc0dJr+hQ9U6E/uCPV7WuTv+iEbscGyG+z
X6lGgk1uFqSziGK2nAUYAnULMeOXmKd8pqFSVCppQjE2ZHoms3y7YDrc3hosFvRh91fxouErejwa
wkThWCvQ2UEbt9RgH4kPyFlyY0lO/P1rtsdPr7Co/McTzsutvdB5qNyCBFYjQ6q+Ncu4mNhxCZc/
LKh0LOgWZzq2Nu4nTfu2Z9jQfD5dzxwSsKrb5k/Uo4GWOrNwR571SrIFgqfatYkNZD+KBUODj5iu
FhOL5k9/9WMvkdGs4E5iJ7IMo6+H4NWsndHazCaxD9isbbyuKwsptmREc+J6YQAWntPN6DtvhxnW
IJ+2oyVPR4DUsL1XL6yaUCaIRf1OMswZ0b6RMhVhD/A6uxuUnzNJe1Vox4syGfQ4Y1aWJTWyRS3K
t8KsKGz5yMf8NFuR7OitD2rnEL3cSL9OKJkoVXtVw0Kmq93BmK2EV2zmW8/G5VfEDZYX45HePLg9
CLAbsFaFK7egU6GbdPg3S3iwABb/P1np6+83UwVgO6roO4HM9dU+eOPkpGxr0YtTszOfs6s353QO
ruz79ABliB+soq5RS4g3zUHPFdC4qp3L3XO4BNTEQtvqE+jA6wHCRrugOkbgWyH3MKpfmMdWT0ij
0FL5yZOCrrmtqXrkRE8v/x03QapS+pQnvuGGxzFxaN+2ai9Th5HZHRbHufI8ynoJnqmwtStiEnst
VZPLdf5ncolZTuKEEFl9FhDiGfzghNTgKt5GWQIcVnzMOQWXCQDiYRzy95yl4jQcYY8uoLcQqlOK
glFANGV6ZhbRXzjnOelf61FFpY35R3+rumT2IWLAkN8EoN2zn8NadSWeyf9quNe9fiFj9CIk3s/9
4t4IUKKpCTI+c4/r8hPIW5OzwrEdoRxvWYFbqPm0m2rynsfytbOb4SIv8n9U1DQKpiJoanks/h5c
NYCEZXFrhvg4ugm2OyxBmPR/B8AuI9PILeIwppb3++oMgmbDOYyIzWxrfnvQoNlWXtzVAzlDz7dh
wgITc6KANG9LdhLC1rMxmcDhWVEbfE1nRRq+FQMoL+tbMRc32FAdsmrKljtLdlZ7MOj0kWks+nhg
ET5TOU8glbEHixyh8Ke4quj+ze43FjWohEILbHweEU3MJStkxgIdA4J1kTgYN7UuJL1PdyFq4Tqy
mX8qf/WdyotzOk90oysJPEDFpsF8HC40Yuh0EZPYGm48FUyctOEd7ykSwHtYfGMFds/orjfLCBCV
kwW9sU83UvmFZntYnmtpMMOja2B8CAthKV8d55jAS0HuaLNz/ev5AKGntRwCrFwCBVs4lHyT78JQ
N2bvgUx2ukSs6sbs8+QmNBGdWCIrw22qcB5gqqvjFRvybe9t7RYiMLCdbXux0fCpb02jVXtwCQ3Q
v1j6jxTXcoeS1yj1jAzj9hvQjSWHthSMDs3RVga5qXaqQCxuHUQAIwnYAcceiN+pF+hYf8qAS9Iq
WSM4qDIKZb8ZlJa6h1ABzErBGfxInpDQ5cP9ol3SjrzDi/fYaLMiPKJECq60U44hLsaQdN1lWDip
XbxfDXc9aW3nn5/uipjugMCbm9LBL8NvrtHCZnUerjBEnH0ZASCI6bW1ylWp8e3D8Byo1OSMeNbM
rgcceiesdGZhw3mW/fQRHWDWBseZsbauzXQBwwE1sBU47m++ioybZuCsDYY0T3o4Ai7ljszGkUJy
PlgqEn3EYoGzTzRx/VeZ1ux+xmo2jJNRMpQebFjmMLCICtFdrIQiPaAXs1wdFZZ9d0agUXjv8at8
oKA7TIsdL6kiazPedwbyVb3bniTgoN/lAfVsP5ypTc+YANkl3riqu3/eXp4p0IeMCEsF+TX/iXge
r2VOtbgcY1XhSFds6BO+2QkdAzMhQWyJgS7T0OTA34QWARds5pmFGfS/R+E2UC8dHdpFkFeMXtj/
55hypajAnwdazkGgDI9NY9VgaIw1bFRotmLuD1je6ugNGKFVVVYrHseBwUaT3O+M6C974BscjAaT
wRb7TqnxQQGqsjTzcrGrLO+Yawhn7Vr0CdQJ97t42jT6mSIMTEEUEOuXxRywseqbGa7h4nZCUaGw
pf1yf32QIRK64vsR7/OhwaxuTxzdK3WeX/i24mBh5NIQC3YfmDk3h8qmU5HzTX8FtPIXdktQ+tLs
nv7Ho5xis41AFYE9qOJ1Y8LtbXg1FPLttt7LVS6/7sk7q6Z0csjbiUV8bhzOoL9LzuX3UHAIBl87
ohQJPR9hxrazEVZEB1r6VVPvf9cCknk/nz8Xsj9zo3jz6rPxbVoDXqIFeGkMuP2Rn79xWkBTqBm+
Rtpzn3DY6/+GPiUEUByl1qDFAY321prS3pp8sN8p6R76b8+w8BNemb04kFuQUEyCn3CdEJVXfMTY
H05uvPoDmrNb8RLVqR42WbvMhjAGHUFcHff/MEMxCRAqCh+zToikk6EN1m2d0fLtGFtJ9l/dvLGL
k+zUiiHrQmDwSJeJJWUgmZRISnG0vgrw6PZXI84xyqaFB853qr8h7fYOmg9Ob0pECQ8w248rwVrh
sClbGhE7MHuQiPSZW1NuKaTvqCg+um9KrtmzUDzxqg+vZY5JIsSdoXHdTTQJnXVEPZFDMcIOy5O4
RWFokmz3WvATsVka0TWQMHorC3CrHDT5SzZJXXLC5/ly8w6CkYAFTb1kH0ovPM3nh3/b+02khFJU
OIcQygbGv9AZOKAW6ZrOJTAnnKJG4jRwW+c8bF7c8w9rHWwxoMeAdEY9enBtdpJbotzKsbtBRZIf
e3YBufW0uEYi1FzuDDu6jspOZrXqu6DPUOMzvhPdeza5AelYSwtmypOfgjhvnvDrHJu50fPDr2+2
Ck5WAB6wt0W48mdx7MSX2vee0Gu+U+gMaNe+oeoxGBsXK3xrbNuyAPf/eXe5Ek87884JzxBdvhXY
EWWtlHx2a63+Ne02LHqhChs4tkzPfpd60ty4JRDEoVlS+X1O3LJzy0RVCobnYzpQrey5lsxIvyvN
ey6C2GUjpV4DvSSbU9HgEUzScuPJ+unNCWMCMh1/3Hhp+ysM9eXL7/LV+MHZwa7jBtTNxGRbTSc/
D8c8Zfw884ctTSwJiQZqE+IfRIOVt2P+7DouedAUkUvC1qlmqFe4od+0k/APgp55cdh8QhITOl+D
cKt2JiF1W6UCSGaBfxzXaNAYnbxhDWnQ2CqSm+FA5Ekb1Y1diQEP6XU7vH03FXpw/yuUrBAzgiOM
qSOFZ6S/hw9mgsN5QDh8kmmJvQU08UsSjiSVd7F+iVC9QXMieOx3fLNjsNFEyWX3q87yWI7PL57x
MlKoHUNpuiF37wZPqKyIjBxAjGUoRZZfjamfWLXgLTPj7rIJ+rf7W2RV9rRGDpF10HahmAN416CS
YsbxKN1oNly2ZOlAWbGBRiAeLFzbTsag2pX/+mEZOF9kszVNXi3YHG0yzrKaQNSgZe8lD7McqyDg
qW2IWN56W035CBKkmCusD2C8/yqsmlSa2ve3kDV/pCxRPog42XOuiLFjMSW0MfeYQlNgIOesf5pI
lwc04DCvl9JqHhxfGLkbdS7jmRErd2jFqGcSnA0/Z53r7SMizXqe/pEVtyx3TmCnvnfUQk2V0wZX
gXAZzIEr+4vs2oBYD+FtlluVI434xhQUBRkRocmr/B4O/sz54pJWKIV4huebNvqMHALz419GSouK
b/YFIHF1V4+LJFYyU6oI/ACNc2vvLZcCjJlDWXofEclfhBbg9CXGeM672pocBefQg4Dbz/stXa9E
R1EL9mBvc2/fYTFd8aj8AfoTnxHnJsi+Ukca9ULyXudQ8zFUDTAT7rpZth5kIbrQoYGWDqkw288H
k0BDEmSh5RNtuotxVUu83sBvIpcN+ZsDzyE9nGG8HjviR2nxQfMU/ncXHBpmXHttxER+0oq0+mqK
IcjAUou9nW2P0/dE5mSPrtRtAay4GHQajEh1uGdRPl7VBgzMWfHHS6Gl+pOp8rt2dSahVEMR5MTJ
PXMTQC7Pf00jpSdm7C/7LBYDyOTW9EAjXZQTR0CfPhAqUgVKYXTsi4bcATIb4f+m4mhgfWWttuOr
jpK7udVnt80UgvednYh5GwbQ+8wAjxtqOBdie2wn3UObZR5J83OfEX8naCBpc+EclDfouYXaPTAS
YAaLto9PCQnOGCtklXhtDvkGaaqmuSJcvR1wtK2CMVu96kncsfpAVSY5H10zT2a7gAgnZNQOjOS6
9lANSpVTnQ3bbwq4f+GozBpH6mSx6llxxXsti4iwpzXzjvUpyX8mYkDHl0kd86SmDYj/i2sOSJe+
juqTttcMcLK+HFvPPISOmGqqXGPwu4DNqgUWje4GcWXLCpcnqSFXtcGcbPq3urj8ZcIIqUUqRx0D
f+zNXF4i+Tusw2Jk/2HexLem40PSLkgBYcLqXb0unBu5dYTJFN6ViwK7+EwLXqnPxsN5+V7DTCIU
UruCDP2zxwepyXkILYA3kXn/AASGRfTtfsK4FfNyc/eqkGKrds+pGHIP/CaZb95ftc3QNjQ0E+fY
XfhPTObiyBVwGhCLxkAIjyESc5SFz/jJ5qycbqDmObar01XlMOR0laDFUPZjsBWmugxvrFL0uceR
wQ/0mEFSXKiboSnn/zL7veKYuIqD9GyvEA8E792Xh6fful/Y7GvFLgSEwtbURmLPdEnMewl+5bgW
9aubcl1SKyCqwcxPqgEwju9FvaXFo+Xto6RBDQmzrJUiC6bRtPigsQjy9bFCIKPbM9+UZRozIWGL
p+/C00ubYJ1l+LPiZIVq+sGdceasmlwcGfEZ24qc45MWcOPEpQxjtcen8TONHyE458zXisaIuptS
dPEpnYdtUVDm9P8pkeRqSP+jM8ZCYnWMbVZ5pq3bM+rLWNqtqJ4BbjCmKT6ujFT2RwAzecb5bKJI
pizslpw0LpEKFugBbOlb139zaMu6EWIiEryfsnrenSjBkL1prwlAp45bD4c4LcLCGaFl4Sty0OBN
1+7pwgtGAGAlNO1EtB41Jit3J8hBE2L8xY5fMyb09zNcmlctM6MTQgzLwGM1wdZn+ymWVp7yhyWW
Xp9J+q+9DBUnH8PCnF3uSFfFBOh5QQIrS+ZnrfCApOI4zj0scI5BReRBXGifXxnbKTQa6qiaEIyA
GfkY0tXe7nQNwMj7kOfVBcHL6P/9Lbi9q2awOg+N5qgQoDitsJdRYiVIBbeBH//CgvF1Ai7PMqt2
KLuFNUjOwmKqTIs1vLz+ztU2yWikWngGKyD79PB1Gfc4/iT/k3wDgP4VjUq6MBL/n4juxW1YH6dU
bq1bE9WBbUmzb6j+lFRPNhjfOJi2hGebb2fd9sDEqs8f19yMRD70Bml8i10U2Ie4oX39CoJiUSeg
vcsS4ymkhj1iyL370l6EXIMud6qoAM9AoQuRvNCU+0kBJSdf10WIV3I+jMuWOy4uPhRF6hwb2Ks1
hXxk9fvT5tftnoJS+Sc3DVScqU6SW6B+QJBrK/zA/XNUjH5jl3w19zOUy+nI+t+Po/MFzic7CVkW
BjlU/Jbtf2OQxFC6fCR3SQSzoqa7fSr4Vo/v8s9LcR+vOeeCejxJjcivfShvZEwtmSZ4Nkpu+xF4
gE5e2ixtUF6zly3t48rDTfFTIC8Ln22Cx+WxpQYO5pg8+Hj4YDhRx1tNQ042py3Ml1kO8Go54H3M
gW0ag7smMJysqiCwD20VBNqQoJfNyqrdEOWRsOTub7p6NWm/ky7hYSUTXAFE6wrmZM7V7ZYFrR53
wJpLSeoD/89XN85bhgpYrcjLPiaGhv93bWLDl6X6TzDt/DoA1fAy8zij1eMK+HidxtNV9y1JZUU1
Ahp5LT6VUDCIapur/nbE7Iu+HxtUIGFhm/pkPtcLQyrEVAEtAdzaa74nrEgOqgCH4pJbzUd7o50k
eS9OfmYtsNVEL5nz9nfvr1aXW2ekTaKPXIzGbsPd5Z9UoEpA/mupPGH/t1otYzFVR6jLGWgn5kgz
Nyi5TxR9vC45+8BOY8sDSmrYf4Jo+2U12lYX+iqlY280580nbGp24zrMDRTNA229KqlsqZLqkjWa
XwRSfoRjE/hVa6Cnvq1QcoohIFH8KFNIv+TsNkzx/MeOkIhphpW9+LVk0vTCD3WkmuNYjKXZxcAY
XOLC+SimpAHvDCtJLeSo3HisCtLXha21pVxklxQHyLXO44rn3scsnw6fXhx2zKUaNpUs2xIAK9PO
qkt+7sqP0QFmGz2mnXc0RI5L8GetlNcV2+CVlwQC4oMGBUEjJMitPbUo49tS2X12ps9tsDPYqrJK
ipZBSQZM8SlYcJ8j0klC9aJZTWvr03fzUw9U9SnhQQ3lZy9LneXEhpBrTPibfGbpr1/j1Q8LuG65
oyBjGEDHlrjszvanQM2s0cAc6q2wbu0PhXOletm/r4gx/5yF54KwR9JEmasi6/87AWkW0kNW66kl
Ou6sXfX+Nn6ucQv+fShCdFrrFGLjyZ1XqKMeiVI8ERtZds8VQUzSHZbIhGgW0xcP4nzzyzd2F2Af
S6fGoLevH0bY/Wjks4JYKWL6RUJWF8zNkbsyIVb+Nd3oEDT1iYKeJ/k5qaQzAU8tzmRv+hE26nub
9K6ApvyJ4BzVmup/aT6PfK6SK4HafH2Qlmm6Tnh4GNdoMPDsBrVDYD6jQTuoe5lTbO7hwmfBdLVm
2GJm5nv486vbarfbCYyJbA5dJoMCz6GngL9gsgArBIFPuyZ6HJIAlAJYM2C35UVmi3e5bleKKzmX
Zrojnr/kUznmlLrFquO1EjtIw74qMD5oBRo8M3GgPHKyW8MPebQEKGMpIUPu9P+txM+08LTqT4Ci
VcBbOpazMpSzn2YfyErdP9mDDKns15CtwdgXcsFeE3oCoHFCqPI5hdt4FhaiCPZft2HVp8MTCwqm
4vRbmElXGIOlr3jcY6fvmvG4wFtm4va9cIPr67hxTfJNW5nCJZCQO+lG9u0HxdJVGuGwOQy/OAYK
UQDTaO6IVQqEaYnhXMIMP6PCSOjjCrZHgFLznG/rZBN0Ab7iEBsvwrsxQlt5p8GZP9Roms7QaHYp
k0Pnei73GGcNkLPYhvPIluxy6nrzRa4iB2mJ4vN3V9WNB4CHnGtNmwrP0y5k3u1V0GLSI0fY0PJG
gYkMRUpIQ680ww4zWxIaiT+9fG4g1hsqD60z6M9hfnc8i36LTdw9yMHT5/hwtVv0vxueD7m3bkAu
I/jABjgDBcn9zdSShsHaIt7tL7bxszAl90m+Zp+gleSqTyAndFfdhrhS8UQc2GGBKNPjklYTwB/u
QjySbV/2q3CZZcd4khP2atdKQPizDjuUGEdY89eWT9rk8C9mrAIzyzP+L0izhDYqLM7vMw+Ef+cE
UhxUjzBYncYFvEtADP7HsKQri9kNbGVONVCnKgCaSgNEL+2eV4uWj5pf7DLqnL9HDalKAjx2J92o
gq53hrSL0rcw94CeK35GpRbNx6IrBQGgwhA2h+uJho0fMkt01CoylGkkVrp/kmK8weC+YnCPR6FB
ecn5ICJAW2LfnG8x3bAFx/rQgwFuwbmj9FfshmcddZ0zqjZpWY529KHqVdkbErCoXzASS9vSQ0kv
WvvcPb3QH0a1xI+/F25YFiYuTzUz+5PlAp2N4RWCB1xXQXnKdL+2GxTNBfu0oo1IeP9REMACfcm8
1FdenwNgTyNmrLluDylVq2dhxX8Ne9BUrwE0joQQY+jXqoUNJC9yXBWvZJIoeQVpWdyUo+pVjTwK
YLR8kmi66yYm2KZTnlLov4aLNQCvzX9PMkydkIvWilHh6mo75dCoJVsbVgGfKOFoHdQenkpDhWsk
23nFRKWVeYFoYN8TJca0f2Ezz89RFwMmJjsQC+iFJRYX+znjhVUWnWxGsRkb1HNPPv8DAPNotvTp
XTvuG9g3Qm7pp7ViNzkBkVamHcc77TjueyAXblk2LJGkyONNOmRuVCUXgj1zGkS3ZbgBPXYnUSp7
79+TJOCGppfbFyffaGV5gI+lumHt6XuSCnbmvmxy6wpy03FRvF779jRqLa418ZkL4FC7mqEzDKPW
cqpDldil95661UumERCw1kTOrB3llA5Cd0lbk1BWK2b4sfbJQGImaGsuPXfzIHB8C+Tf3OJyKdJY
DGrCET5GJIBmLi7L6TCBblqSR0PkTsZYNQzho6NeY7l8Z7nvKaNA9LbNawbe9cD9YRgnW6KMcdr1
Fgf8lLWg+JKLYUd1PyLAtJw+cqnYvGYCvn+tsFudESn0li77pYo1YilKIeJAEf5sFzj8k7NL65MD
RYKxnvGIslBbiu0i1PC6apqx2qy3y/LBLtBl0cgmfxN9yVA2pz2LaUQQ+CvKYQdZeAq6YHQUXF+F
ba9mB5oIZOhUNl65RkJqrcl9gXJn7kwKfhEKh9fniIfKimHOqSLDGNi9MS4I+ESvctr1CF/K/Av3
vt4ddgD6MC1FdoF8hxha4P0fpTH4bUV7c09Vin9gH5ZCAQCEzpff5Q7Y39bLURMu4Hxti5OvOkw4
twWAhwNa8Yun5XRiSw0jvuBcYdJIu0oXjGdFb/ZCmEOu9RHtZedItU8H/LxPsbZkOIxHiKJRbS7h
5Y1CIQY72yyQFKEmkaKJDPr1wLitKfmY5O7Y2HVHIt3rCfHnYyKVvzWwGq1sDuK3xuE8wbGttVtR
ITYz6Oaaap2JPkQtyMwzvaJ/+G7dDHD9GLBFe0NYwzNR/SN26MSyQ4JEY/Zyyo9PA60mu37XaMtk
P8UM3QY17U2xiDteNJmHBaMacdF1pjIV6ZRq81LIVPs0v5BIVvfFLzOBChOc65o+i41Ql8N5L0UJ
iFlqYKPF0O9dBbk/Oz2o2bRMiGHHBooZKnyW5wUXcl4mlqlea1QONvTQr/Hu5Au89E3Q9nguycGz
PyYprE4FdzyEQUxSUmr5F8vxH+5qqQ7LMrvTR8FLa49OXGFcQhEh6fKoLGKXuHJv2AW3tOQk/+JE
7FRsksnt25ps7STQbNbUQNFeaRPj0E34MIQ+MyBeZs8rneu7nja1NELZD4BCU5BOCaddfL+3PTVa
Akn1g24V1j2Ltl+ijQhR6YUWzM5XZQ1OXZkddgbGnOs/KQXO8kYX0lGVKgCD6Nc7Dqu7IJhcCaos
w1d4opUd+1TABw1t1VurEL/b6o7F5ItqmWhZQsa6qibaYFF0gfwmElZ6SUdRQuaKdQuVLyMrzIh7
crVCbnpzQt4Bx00ie8+pw9d5i2ctarmgV63TrpUInaC1PQEF+vLDGGT95gPMZRyfZUt/aFJwJg4T
k0fZTfgsKi9F5MkErvFtvYApjgxx6yN3L66JksKNZwPa2cZhaFMyrKmODR7pv9tgzvXkM0hbT0yQ
wVEr79Ldl51Jar/Z5YECi0bdbRA/kP6ECsUcsxvqR6GPmvX3hXxgBRi+xU7X5r3a/S3VS8naAk+M
AARJ74ZoLWSdH4gX2EgKDQ6fR9rCXhBKV8C0rWfiiwtMThJT2QlM/iKSFYHJ/r9VoZk8dPLkqE7W
YZyNrRr535/3+kh7XArDYYyD9aurW8RDjnpboouyQmRE37f7tmpwD+3smfNsBd3fa0Esr69HJ2Ve
FQN7PhSy6ymmed8JsQE8WJ5a6yc5mS6NZ/yU0fXRX6eacB0qg7yA2VE/vsVTRNLzuOrQw4tQ+VcU
a+FOzHUACyAxxeWEsFjlrr9IzEcrPEHq1L4ua12h92RGrBdHFZWpltfWmKxufqq20baOcgdyOzBK
X6CczGZDvk+uO0DYZZXHFKFhxfqf0CVzRP/qKcPa8PLWnfzMV12rdqhG3/TFyyfIXJMSz442YT5/
yHKAUW5hdewACm8rjMQQdN4hUReuBhRp6PBrkDUDqQp26Ps6X1LpSbdIQLeS6c7J4j6JYS0hv8BS
bnRryg9cBbqTjzRGXtbpRBRcQ6zIoc7ZKYJsnV85FGXbAhy4fvdFTXoul20wV1knWlacOBu2+h3f
vOHChWW8EavTpsP1TZ6ZEQ4v6cER17jj011B0pkeYjhwTWDeFaF6orkoPq6pqenLARkxeQZWSM1v
CRBWOz1GPamy9Tgdu9F++o9bwjrLh9vS9uTyCjDPvgQl3cSVnzO7iGAXjw9UMP8VNTqNxI+KDBq2
I74h9Mnqk0a6du2CmWEfRsECSnzJt7mSc26xeT5UfDhyjtSkChEDPFQNYzGiRMVGlKoWxO9wMstc
QcuscJmwP9EB1WbPj0Ahlad9x3LKPA2GjphqCSeRjT0G00yIUR947jWDPM5vJZuo+2m2SAnte+jq
cKX9aLhXu2Sb3Fbe1gD1NZP+FyJZoMnB4sia0uYZPLm6/OtcJQMEjTXkI6cSykvKnWHskNgPdazc
/ZrQMuirP0xoqn1DaakT+z4DZM2LFrlMruQW/Z0hEQfMdSBR7xjmFMsCvde4RN9R+E3pl+I2nnOG
yi4kX8W0FEI31kWSTxoFlDxkhYupm+rdOTOvfwZ8732qPd1w60iBMd7JgGZ6LUOLCmePrndsLkaj
0oJQt+KOfRx4EdgdC7XmPWd4Lgst2lXmOgy20SJkYJNpWywykHIGshvL1gfM0cf6hC1tCNc73q1X
jtlB0uz1++EaFP6KWpc2qvnnrQkMDx81CVy0/Sa/ySmsv3+Arn5ioN1LLwm+tuwCCL3GQEVqZXqa
Ge5VYtIWSkuvBZCAKXUFROJH6S9MnHO+66bS7jlBNR7T5jA7WJ74H0ebj4QM3htA6tBR1YcX4skf
DdMZ2oM69O9mxxbyw00qwqg0yCBp53PC9R02MME2eDShQav2+FvIzVYDRUuffjGUgSLJ9/v88GjN
/qqELECnNxG1tofwMISHGXXqlCWZyoRSCG1nVVy61ZJQgygmld6IOJfNZnMFSRonKVjsc+F7nElF
/YfjLee8UWbRzzBL8tfrso9blwgMkOFQQjcvBHghXJ2FVR4j8GZ0XGAF+utJ1IlCbqCH37UbFN1A
sI7kRvDxPiFam/YaEb19tehZk0IqZ+pwztQRBQdx1rwRQZ0MiOKLYRxAnuBfm/4hTWSKfkeSCfiu
MXmTTgRJjJOlHBf+aZuLh6L6/c9SJxACagXlZxHSPMExEPkl4LTppv96gyP22bFdCDOhKstGSl0u
brEHD8Z8ibKwOCbIbsTwdDh34ebroSDjgCVePOHG6vPk5MSsizsJVrhP2ZL95rNB4+cUgMktSXts
AVGdtYdNGYDZeTIxmo4aSqdfDUdCaaJgMJepHrJG/6Ov+tqNUuFL/uQ65QID96RzlybvFzDE5OVx
EM9A6KSSeQqVNSgzQvTqP0P9EP2+YNp6skzpjvCT2D+yKf6a8BOgSi3yfKt43rdkZdwVSnGg/EDz
Pkz36id3H+iCKhqoGVe68cmN31MiRO+EdSeNFh1jVwVzTqlHLxMmTSiqpExxN1jnjyVfdLzoqrD1
ad8w2U9x97h/rSOhIWI9dNZDge3Bw5rXLdWZrtOF4jGhF+xGd/xLlS0PGXydKSQqU0XMBAqEucYN
hYi9hFHjVKiiZy1Sn5H9nHNAtmhjN/90bB4dzBLhOw2NltWIEYp/6cxm30NUL6XxFTnwfIvmLKwL
6ivTsSBqesEf8gmfHzW8F5V3A/x8BlK2e9EdfRyal6D1JhqTZW/+o5kX1YEQB4rk2/4UzWBH7p4r
hYqv9cNyC/5UEgvAm9UtsCxNUbTEVXUebtykBCY3StKvILLM+EvqKc3rnJZOQhiKZGYS0Job7YRm
uM2sJTE+gAI3wSsG9c0OTPCZk0csd/W4ahwKdWX9LFrJ0XJG7WdSOV5I+3q2Jwh+dabwRRFzQrHj
OXpImWIeGrmeKbAtI4E5vLjxpPLuu+eVjo0FFByCJseeLyRxr5aCBjC5x25k2wplxP2SN0tXJFQW
jEjW9SwbH8fByAXyP3GsOcE6peW7ELxG4fxf71V6IjJ8yrwzaukoInD9Vo6rCIo8r1H7Tmrt0VWk
VMYrgY9uw7bRoUQ95vKEL3IsyTF0Xyy6FB3gGX7smdW0dD9XA80ajw/jZmmxaIWDQicUWnzaW6Ii
scYK9aQWlqLVHQma+UxNW4zW/Fmq4gbFOyCLbHKbhj4PwlxTX6BjqgzF9EUC0i8ys/USmqr2gf/r
wG4h5Q1kZnkE1V4IZtZN71nSAi7n9wiLYq2mNSGa4rchWw2xpJdDPkQy2gt9Ibv2KF0kWI+Q52lt
nW07/eCNQTYYs2YffP/CfNB06G3Xr6QEzegXun1EXpwyT0962xPnHO4rJNCR1ETx8YY87aNKwAfY
QoV1/4JT9g33bf7cN8gCxYeUrilOfFgDkd+CcktLbjcRowrHWu0G3UZQ8NPKZo00aaiITZBKolnE
27lc7GoUacfyaTO3QXUIQOMp+mn9QKbtOLu0yzrYRcqBZDCuGm2W85maKxXpXm+DcRUjkFks3xNC
RmJcNySs2ycP2wSAEEWzYVJcjh9Bq2Cxa2uXAQh2zYIi+t5oPHKKlAldv2gniB9TK9NuzjDezVUx
PWwHk4y6RakzPGhLVPvrECCFc3CDC3cIwzYZ+QG6KBxAngaMXhQZptTIWpfwD+53T1zLyWXp4egJ
+04Il8Pr6ZJjN8rozXXL3pnRp5zmHyv+JnsX4uDRMjlWl03ZD6gjX4mkp9f1CWI07jp1JpZ9s6vI
xK/RApeF5Rh3Btr1j7zJg+Hjt7JLOQe9YUARrMwCUeASPakRb8xAi5/eQDIAHLwV1WqQjM9pUHqN
CKXfoeoIr3evY7OWXaUNTvy7tU522vXSynptzqkzf4kiPGwXpRCXaNZrG0JUf4FPrbzXBqfTZDTh
xm5iJMlYM2fNrSWq+IR0JGfYabtR3U8vgkWRFL26s9QAOFQb9LceY0Sd+Yj5nKIyGmu/gCpNWJ5D
ZzXAPjV6OE/wPTBn4bCO49Tf0KjQCcIrhqBzqQvcSxFw1aN6kJYfkPWwGmSXURvkyBMsSxxcva4w
jRNHxKA3etwpxRtwgCELayFnONJU/sler7g9G4C5G1/2wYrfoC2z2oCEbj8MU5gDAy9OoFpwuMg7
LrJ35hGgQlXWsf+Bz6npq4CNEDuJtya9VOdfbkeETc8AMD/AsxPsRnkCkYOR1rn6KriKbxGR5xb3
ZZmVUqQfbD1M1c/XYxkwkxm42RMlOHeVOdEW+y1b2GWblD9OB1hqk4qMmDagYXfaYWxgZZwtdS0k
pcbRwsnFunvDbZYBswn5pmdVtiHbY/LGEkXdDCy3qYQySO4QRJDczAj3TOZTONIFnJhIqYbtfAhR
C6GzWKgUUXCjEN/Rrf5F0vV3foWZzbSg/d6U5Mu+IbPMNl0dfI5cTkstCa7mBYwKArTpKfiwz6Av
Y+xswuuk8ssYDNmotWnqde8B88nefFfZ66TeqydFlseK+4pFvsAJOuxLOgtzidgdH08DW720IBWu
JaQmuOSaycvpFCxS4zKMhJ+lqJeasoN99/fK28evs+h7KjhcBo9ylDaSjELRIQIXv63pHAP/62AY
yn0KJEVVM3psou6SXuF0O3QZywOEAPQWCrX/JxvIR5XYPR3/ZPXp8ejq6fQhsv52Mp291OTvfaEg
FMASC3WKmdvqI9Rw5pmdOdkVDkN3g9dMDd2lsTUWBteEn2j2NXS2NwKuDwbaUa5f9li/ZUXmOllH
i698FR6Oyovgj5qH/XA7zrZhrCJDGnYNd/BGwDNQ3aa29sQOz8oojYNXh4gBXnFYRTGu/lwaiJ40
5S0B+TClXPh5GtacYq5g48vx/LqMDytAH8XlmEvdGdZyDM8TVyjNo2+VNP/5Ze+NY94iuROQs7oo
d57BzbN/00E2Rk05P2C0/LgV0/7fDTj4CotoaqcbDUqFxJbnzoIj0rimIiKOsEmyE5xF41aaTR/d
Ulo50pW3Ka0eEB0JvkODPH5fQRN6SMOVNPDimRR2xM3EqIghv/96eFYbnXCSHNJTE8o546OxZJgX
RR/djs5A4Us2QrXgmD9kEQewZg1rPaLwIB0kZ0dUZAenHRsQdmX4AWAlSCKOlEUNanvD15Je4dq+
vVz6EaYYTC+XUuLxDTvJwloLfIOs4vSTXsLlD6wD3HVUgugm3TcE43vAg6S/3SfTUnoDLycj7Ix8
kQ8VnIW7rGPrPCLgrVDwPgz8VqR8YqwPY4HmWAlFFGwpyjkMsLcZeZ3rX2kS+IQrTF2eW6h2+eDK
oW+twuIUuzg45PKqkPUAuFwV3F3FEmhcmO3B2aXSkOpT8CKx/T8/NRRCXFkTTtJAesjgAsZMFfR7
Uo7a75B+2sZkbdVadp9BKmMqeSDUnePlL7Nu4HCRAOp8hE8rnZfjkTLq5RTSKcRpT9z79AmIgm2b
ImMemX2tvSujeaNIe4mUPI9abu6BnRu86PAG+whWGbGG4O1THMzmLia9HmJ7QwqpEKGgco1o/B1B
4xpewnOORTKusVNksSa8AYdJkzWPdNJxa8A3bVBBxd4AQ+pcmAs+UhuawuueatGwBkcWHuXsHI+4
hBfmNgrMTLfhtlkrAmRtIGv90iQcbRA9f6/DqWc/mPbuV+TCM/OUWGQUBv0SrHUxnC1a4IzbrboS
Elogc99bd1hJucZD8dcpotFhgrFWJw16a5AxZhBid/klzZfpzcSQC0Vp0iQE/fOAdixTXglmI26F
A17mkw+vBH8p2TUkdDv73WknKan9qRqziQjI3SSXd5WCDltp/ALpoCkBtlR4g1iqgulGXhvYWzEj
fnGtndYiS1LF6aYdW6g66b6cekA1B8nbbQE6nMZ6tmPC3Qq6+afShauYgz2mLLyYLt3KSd3Mx4O3
KvgFvvGng+dBsS01MUDSF33zJu6Od/uAkZjLRQxbvmDXwBD8PttU2USKK6xLP+opZe7BhQUskN9B
i3cx+1hjRvO79tVe7AaJINtW8kpzcsMyUdZiyW8lNm0eXqg6Y6RMwkyrfGQeHZwZnPG406IiVFAH
I6Jf5VIWGHubix6fCjPFJ8OQ6rY7eDICrer8bq1i06a5WTHVywm9BWVxA96V+rlc4gDXXLqKVcTr
uaRZC9mtWOAkSkreU+14ckyAixwYjUc0Qm+rvWnGnKsV8+sRU6fsLBYTts77y1ZqEaKC844nj8ps
mh8hXuREtkYGF4E7en6IY9wnEuygdSD7PM+NPijFfY0wUgJU+P7jX72dW4Ic89QnXcj6nBmRYv83
O0zdXdonDsEtYAyh/CDEmmq0MIP6lmSrTW3tFwkZDfg2QF8l/X6enN0T5zfUrE/j+PJMfCAdc3w8
fBxYdKEh+D7sxXQNsxhE/0GEfcgFxyPIw7BmUZeDxfMuFZsCWY7NUnk76o5X9QczXDNt+SkB7hG3
1V1OsGlpzu66cnFt/M0a/bvg3XaRA2MtaUGFYD+ID0CeFC6SGWgePRTmmLrNmxOfM9RC3/cyotBz
xfFseq9AysFlf/XCr3ZyM7igkUW1NrIG9trGoFalPNKfG6XQFLnzASPjrHSmYgu5qvubwG8957Ws
u2RiFMOmVDTGRMn4GhXmMiUQ80ioO2DRHXTg6PzPS3R48wPTxTy9jhdTAdinD0fpbUz8o6O5zutz
WzmBOHa1qn6V0zr6MJZxv+C95Fkc2Z/RvmvGCR2BXBFyHBjsC1Jgk+vzikraujF3zokdpXeuv64Z
LWpFKt1k5V+dI+QmeVPHP12je9E5FFxiO3p7koGF6bx06yAw0Y0GbmWd26N6qQSTw8SQlzyiwrec
RF6tLNxUUCSkJaBXpKDMMigKR0Z3/0T2f9RZSd6l+8kM7YwqffCZjAkuCLfD8YRp0C1vf8wq+Yzm
0MXFYhF0IOZnO5MFyOr2nmWEGGUiCdrtm6gjC8RshI8TyC/C1qkDj3+fswWNjSbFX395kU4te9VV
YO6yC7oyQxwFfu4HQ4apJKFiEeeiCSme7QPM+SP/cVBdKO+2YqmUcFGGi+hLdKIZvgpCQRRk3QAe
hMqk3qtqGFcThftzR8pY26XnEjH+e8QuOV8/vdY+CgP8vXGpxQHTdBaieejrmsj95VAEcPXVDYQM
MmQvgRgG9M43sWPdYHWJP8r287NtjvhH1DnUEj5E3khblxOgzHIoUIuZ/JCxGWpVmkrIw7J/1hRG
sLi60qF+hoi9mt0KBYmpeoIptVw3Lf2N/rjqz8LC9GIGxHvlwhhqLNrtzcgx8tBBGCiJMjhhNfl4
zk02S+C2ht6UVrRI+kSPwXhJvWCWziD8TWmSbwdry5PgyCTPTPCJhvHm8QEqRFfme9FiJpbdrbqP
iJpR0Dy37kEXK5V+GNBmF8l6wZ4tPWo3TcZy8GGmcbOZEVsYwBzJSE6q5Wun8FmeTWSXJgITBUc3
iKAKhFdBN7TqPPaRUA+5Qt31029eGVVmZAtAzY4LAcE59pGbaSXcZW422BK9XZWL+rB+6rrKa3i3
HoS4iKk/btF5FgLDLGWyFLDMamOXPwaBpck4Ic7D2/XxysrFnDht8rpvHVDLrkbQ5rtF7ZZYZ9Z0
IB5g1oLI384xgiOkT+SNlyXE6yg4ytRJ/GXNAp0RXhhXA4CFfQevBTxJ9tETHR8O3F0bCB3Stceq
1xoA5uu981TbPEWGKWilD97I6DFIR5OcPZtpgXitLbrUeaeOR8IoqT49TxvLQ4gqNI6CD/GPNiRg
xl9i9VGfjmXYbQs0ZkTY8CnoUpGuDzXdkYeAvK235zhQtXiGaFoiDdL4LW5Y1zpztp9Ual+IX/hC
iQHYN2/BfdaEu4uLLE8r7diFDoLmW39/Hnhf705zL7aFpWafD4NnkwCofjz0ya7WolnOJfCOb+EW
Up2Bttx+smbUyB0cSIr8ce3rTGWyQY3j3PZpLoZP9tCc4o6iInXI7hPcPF9+0c9Qm7Zy7FCoAVo8
WzHaRsG+z0wiowCS384l25N2kGYn6QJhCOq6yT2f1qG7sUFc8yhyMPXLeQpF1PPlaD4pidiECXXz
keOejzFa8TgH8hwkdJzEnA++ua+q6lKfep2OzQVfnaTIiNCsTAu3nvVYnb428pqaxm7xKmktz1rH
sjQPbfJ3ByHT1CFTSr6oY7aVaPxLK97QbX1ZeNWFOW40UNfLTgwztrcSy5H9M2eFNTtO6PPrB3IS
CHs0BkKNq5mB+IEyhiERURlno5SkEg1ScbOAn9JwZ2uQqBi6W0ZpT5ZUlMtGVOGl1myKcvXmnXhb
l0xOY5kETVgb0W1MYGpHLJDE3iiG6ZEvwOs5TSZyi7GkjNeyqynhIX+ydvIXaKfhSO8VcK6V0kq+
PTZfar+Oayes50tlx+88NovB0JscxDYnCu4VeixKjKCncPJjziL49RXEY1EFNOjFuhA+PXzu4bHz
LATu3JlabFK8KEEjwQGA3c4EAdqtLz05LT18D/ArPHdGTxXcUuaPRLCuFYfE8hIzkBoy+sOcMcrR
4xmkdcjVAvPjNEeroWrjt6ampz0Ob00g4THdWRmXsOx/lbng4d5LNhIvPzLEPD39ZvVpyKNizCFe
oqPdmdz17JA/DUwKAEH/g8baQ/gzCTOi6HuEhGCM1lekl2dSvJBzU6KomaqC45QziRkNdT55tHDi
wztuB8U/QxIhBeRwA9bD6VHg9EkASeo6VpZ87NlPffeGO7P/YVDJLbVZbLvlmNCE4GQAwl94ZxDw
ARTpIuHVgs/2Jk7ZfHuMTSd7Fo7nvtectMCupa6ipfCy053FXxGN8nSUkLDaHhnH1AIpBv6iutK+
ubrPAMAN2dtvFoXedMMDafs6m/rFyiGXVghgYMrpN8RRFkm/nmBiVIUcs0ITxNxrwmSiORvxxmg1
zcyg5h1h35oRSYokbs7ms4LZqVrmOHfIZSZpuPBk8VJ0Ebm9v1AcWGv6Fovh0LVrS3JeZ6lF4s1d
jKNQbABc24KFVf6fl8f8vMdk5lEBZy8hDwghk53/f3sdiw3SXiKjJqiLrc2yLwU2tS93ir8wGMzQ
nUVoe4kE8nuOjlLdKgEfuWmhXbOPdyF0U79o02oPRxC7E79r8RJKU1oY70/2DNRLtgtkPIYO+T/n
5cRpcxQZIDCNptUodmigUpFoPZtc9kaoU/5r4b0f2lZyAM6fCdBtjFGZ2lRkQrwjtzHzrSi/AZ6L
Sw6WK8HS/g4lAtp9gqdKNgDfAIR+FQk61TiVjgFIordvuW71643UiV+EtKSbimzkKSx0z6kBEa31
u9CLNJbXCbgco9SadoDuzCB4p4xLjQ7LcuyxnK5xbZkg7LuTwzYm1u2jeDIBRaKCruAfB3mrNYto
57Wzyt4PvaG7t4wdocNMYJp1Ujul38acHqhLWpsFh2WGoPMuVTC2+im5h3dRaNQJElFo/MzWeceo
yl47qeaQlAg/jxbgG0NVCt0uYZn3FpeTWGp221UnoEycbT5s/yB4LqPCLpQqV43eQzZl7DjF/0ze
8mV5MvcdviCvvoHKOo3woSpETMpI+S+67Bhg6AjjfUe1h0nnkPKB0MYkBey2VCeECioaNeD1Tasx
l2WxoDRLzTSn0HKWPjT5pMebuhB70NHVkfLmu0dI+R9TyJxpiFRbCgCoo59oakFrloQ/akt95gol
WWixYhu0HQzqLsF7zI9weMCjK4IdEkbSogXLSgN3dnjSZ2jJdPMZM24Igum8+4h4ky+1QzkPMW4C
18jDAM9l0krbKbiUcQU1A7+aJ1O7L0p6/upEkrfqHnH/9FkABmnyHMJZUYkqQsa3z9EebBQ3uVvR
N0+rI/SBQb/KhALr7ehRlMjjuGyx6oNd/IdGw1LpqxZqgpCymjOrg8/kwCDhpcKO3HsGTqjdrHSp
zsC4mKnZ+V639GfDu/xiDk7vY+74oA1K6gSLtD+C/r2UB91KSh1omGJj75euk7ieZHHbvr94ASUx
9n08w/qToLmR5Lbdz2+rTKiQM5X98hBCmL/q1H8JBijFJVtgq7n+wAHrsXoLNRSh6IzJ78It4Azg
DoDZuInbCChoKGEg+3mqdmPrK6otR7N7HAmNhcATikn3ki3598Qt44frw1h4bCWit6eG0Jnp9ck9
12okilOXfXm1KQvVXpkCJcHtZrQeMYE9bVmpJS3G1gY4pNT1AayfjX7tWJtEfyvNFrNnLcRjcisP
x7uqYUrf+7M+CKjAst8YpYvVBLdVmkuom7SbD7XGOF1Duca+CUw6wFj4wA5JemkaAoR0uFjhGA7t
Eo/V0SogqhGOaxO1hGgQTE+Olv0Ylj+mH+8CPYR31NfeZKpZBBvAGP0vOmq5K/MSlj41J+c3XHNk
xeQAGrNIlb5F5CAjW1EThsuRrT5oQBYXW6df2WyvrxLL087VTRy+ua5IndK/aH0kcQctHyzYr6NA
2uocbFIywSKEehDhCEmZFwXmo0PDcvVuVhqEUd7/q1W4B4sKkhB+9ceIzQV0z/MH6e40h4p0N+sF
ZcwRCShaRIXdQZl1BiHFJizLSANWNjIdSeZikiazKwgI0pAhg2TC3FmF1bbirAq/1JWPZFysZ8Zn
ZUBvTS67EnSjoeEUspUBge+IQ9acQQfwfFaDUKVxfEDT6pYOgBTTYsZ2yzQ1IM+NWI5gbmYpRkhd
LLzTXoUH/8wXKkhpN3kQRQjRGgwmJjyvkW58hZoYOzGF1P3jZ7wNSMf9XgCKx3kBbYU9XwbAO8kk
/DCFmMZdplCqlZD/3ujFgFVfLDQ+f5rqHu1IMeJYwYZ+fygur2r3KvMLZ/gsqxwD84yKG+rcIyzF
0lHPDfUM27Rh3YxM1deVK9cXx2KFv9Xgdlun3Qs1lKa4B1RlOZ27XFpyi/ETnksZLLaUcEtGunkz
9BNg2Q6rCUSbxpMBtQu/ogPVFmJ39UEZFChc7MOumPM1fgNNqsBGuMiyyQhxevTG7o2ZWeMaxEwH
MNfATjMcUDzsWeJGNGDPIM2RaDr+wqS/yCx5P3xeU+mCoVZMOKAq3ZAy139mhB3EEH3PmEehXSRu
CBCKrLngVZ4t5UcyWN3bJVU7ZBR35fgBBxcrBxuSY6apHvpcFjpIJxg02VCZBK665W3YFSgSeQ+w
Zezdtk5AEQ3uAL5qXbTauin7YGdqaBzdRM2l1F3ncm3kOD76MJE9tEOrFg5I01xL6iPKRwFhNFue
Q+XdR8I8u8N9/8Fr2mRstogi4Uu37dKeKiEQ7VDanMcEQYSOM5ixHNPlRWGrPqLXOCnNz7J+LyRO
VVdh0SXFeEzrLWX5hda2QdyGYkziuRTDa639HRJJm8MO31exp+y8eRoRl4MiAS2U1tOvam22vcXU
tfVJLxo7bpP5Vro6BkYHjfStxBEjT48Tic/QmWgNp23RBCvMNpH9gYgyD3Ue9TeTBhCzqUy5cve0
PuhYKVicsYNogtLKcEuDLn2K4OzLBdmrOVhOnvxhvWRPzg/ADd9oVV+vMiZPF0gObkaGt7KnnC3+
9K/ZgqG3yOV3/yIQmdE0thTJHKISFL2XE7kcrHCIiBLhc4aECwa+xZvlwnZ6edxvhkzyDHvqiqbF
R3V4dn1h2q4Ysgi3mfkqJCTBchXHTXMeYUXvFwiDswdlagEVsRBnrRt3XHqeYmem/prFOS1HBJUh
iuCA9kx2y/9xHC6TMk+GFsX97RSaC0vDwJ3Zdn5At+iQuU70et6AWxBPC85CosWksbtVLrsj82Fr
KaS2pMAAhCYU86NnJOBtHJKkfjSGB4zCbfT/tHaC1yLKj5VhW7USNqqPO4lss4jiVyWEGXn7Rm8X
o4QrfhwHRjwchalNfm0w+veABaS3HHBtcPPbE7x4fOeJ//8RGuW94B5FEI7hCQd8JaPdMAjnJ76x
cvZtrAyGUsHOfXdBJ513srzSM4CKo0FLV6po80sl+BA9HNlNNMbGwGJrnJ1cYfsf3xtX9gQefAQy
SqzvWooz61NR1cx4fUfWA6yaWpJfCsXmOe2zMG5A+KzY1jwr7D/qFwa0jRPCyQh/+MMKR2lY7GV6
r9MORTkb+LCv2wfPMXFNDZ5vyfyycVh1gdrnfU+G4N6PIg0Gn/936IiZ/oaEe34mdcAdLb/1Z+A3
mzKsilCuBzYE/HsqolKMMrowxD6pnbLnLb4xs5Ytr0uy0w2+4p+/ndpU61xCCqAxWNoDWWqINaya
hXadJJAOOq3sgh8y74QP2070tBzfh2hXQxqskpb2qK+6iQCm7OxCUskxXJ58BXPi6rCErqsvB62Q
0YT4J9euwC/dbA7NWV3BYnXUbykNHC/JMnEaBiBiC20OBhslZslr+nlsx3MV3U0wgPMxxx8BgD0I
ul3rg7SEUUoLI0OYxKrMwYrZMnjIO9lfTj5APB/4JHsFBlNUJJo8dzBfn8gfbnDuhjXN10BC1Xcx
HsGOkY1qD6IyoYbFTLWwRCz1KeqOfvqtCRF4gKY2G9K4NfbnTrNNrIC0RN+qz11GmGts+mR6m8zS
oNX2bY1TWS1doY8ZSWcdIHxi+p83jmRD43fT7ULP6FWi/tEEyFOdfJk/oVA1UIOMs20rsOiJQwVr
fGPIii3Z12Oz8dVNcn11LTikokCh4qTREHkTwHGY7Hcweo6pybIEw7STWhcftz0Il226EJ9Alcxm
eCtEApbrTjuhpnUUHfPqTsTWYS6lQwtdUNTtdofyRBFf9s9JXs7RScpj1AaQrgqBcAWUdABpUhLg
3l4qwwdLftgD+da4eQwB3KP+PTawnRoAGEXvQ/gZIsifZ0nJnQKU9+6E70/QvOYGNrfh++KsjS/6
JjCEz2DsKwaMeTOiQD5nJOzZHfQucbd1VqTaaPoS6MvuD5PFbDx2jjtiXNnk14Ki+qMABwOOZ7K2
+BvFhz0NNA0HtDdLrzD43HpCi468lBtvrPisHhxG1Fexv6PmrHxMr9laUbrobeR26ZYSs+j/fDvP
YkaBug/wYZ6Ablfjq5uUfc3VzV48QmmYqU8P1WWzOraxirKH8LNPBN7XocI13d23bxS3vPI3twOE
YuaXGk8CxmNLgyBsuu/+URU3iDwl028RhzuzLE35jBfvquB2ImZmTANHy5L6xNqPfHwp4SSjx1Rq
1XUcgH8t61aF9JEA/x+msBdZnHwtxdQzYdha9x1jRjQNpjzzqilN0UPrX5GqMj0ppitOubJRVFnw
nEWZMXME8mYYMfKNk5k7vJrmsDMCO2bUfl7NqVMZ2OA88gcjuEitWfDDgWnQyk8gmH915lDBCkGL
eKiwgEDkH3hs+XZ2X+DG6HjUd6BwDno1xpETB3ryU9RsOY2EAwq0l4wqWH3ok7d9Q0aAV2lhvgu6
tNEcBTorwcP2YbwRxMmoGrnTtqnoMjgkv5Kqzpv01QkTSdl9XASHT/6OSCgmiCPig4OsbvqRY/xs
lz5BkVzL5emI/8XiCrEcirm68oNocD7vWEwAKksxs7Pw4W+ifKZCRaMGPZeLICeq91ac2akZB2T6
T4LfrkvdY2tbAMxjgmYrIL4ukzTpVnKjemue1N/yKh4E5lQllEB/DCH8u1EWRcOBMMIzvGsyGWiZ
XRVOPixcMgBHqcW3w8ZHBqGh+FxG9afXtWCEPiKPBXt4LzkXO8himjqutBOC8tmc9xAQ6EgczWeO
BZqAGmcZa1seO4KbL76QzuSwGaPyMuM4VGgwgiQ6ARg2uxRQT7E/E8uQSEHTj9l2N9IX7dABfYON
PKTtJfRgUORh/IL7A2tHIcj2uZ6SogMy3PqoDfmKYzdf/2H/R7+ftXH8JfvOefpOF09gIfNnV/Jk
0NEa/a37quS5DCPZI9uE+2TS+tCBk2Hxh0d560jW+SQq6C4YIQrn9w3ZBbgQttXlGZy8ty2Ht2IB
yJQzAq5bH2cRAcsaCxOvK02mKiNXtDpjLE7JW7iOwvIdV8AAYPBBkVcNiXKDzfqI0nGGL4v/rET+
k6fSLa5PWN3rMCLm/c/Z0GvQ34xIzrjm2Xy38US4BdPdjULZz+U2GZgfmbZMbd1lnOWy1cbwImnD
s1s/kcrcYGXUX1coGzIipTuC91pm8ksMgUSAD8M2MUqh1DEYnjOvW6dMxjaGuW+fyJ441x6l0nfK
XFpX7OX3HpAvi8wTpJPwuYI+bUZAFpq+qCkPnVCWBXmkK17k9idVBhtTigz2sXE4zgQrTUXzO2xz
2hoGRb6xsS0UVtLruwBZoeynYUNTLG+EqgSBPH6dQueELP/WiAjkeEg9PvH01BhMkVZJWdzh6Jbt
BQ3wDhIbGDsjvdw66tnnlqToYkoCIrTu0XsQ4Gl133RTOoEFWo2e0mOPFFwvrCoLDuKTG/TCvJva
cgRvDSdiYqXaJ8xzv/I+PQEiVbI7N3hvi1qNeOasrFgiZ5hTwKVjnzMOni31LBQumd3FgiHYuHXN
rZuPGd6OwjKRwMalE2pIQvFEoRrMrDvCKWC8668Zy3FpWYl5XxFPyYMFxI/hkqRqtc/YnplqSo3y
4g2ibJYmMzfHQNuEkexZUgWCavTHEvYFdSlF26aRjNpBoi6Q3KN0LPRQc5h/L5075VtkOBv3xxop
LUDXAwbbz4GaQSQ6u2SOGconDSNkQVrSSwBHpZf+h7qMVrOgRMldLb3PgC3pKq1Elxe+1/KWQI7w
3nEmjZuf1EHwQr77M3awHdlmjXaD8rwXSojT4bAuHM5anA+zKYCZlwORjo1T84Uw9qoRFrZ2ufAN
6mFc0d4ZagtqguFpve91tA7yNZ+KG1oUieHdem3Aa3cX1Ibzmi+6knqJlXH3hgaSEMNfWUOJzWRu
41ljSCPA0gwbU3PdYUFO9rDQrEoicZfwW6ZC4i9tGrcOC5g7ZtYHO/Z4uwUX/g15ReZ3TAZZe1re
T0wDETUO1VSsa/qNPcMYMd+gii9OCbeEZ+5HVkMIBlhJcHDkcawYb+rhnyiIVu9guBTXQrW7A9cp
wTz9ehslGqfXyCLSjnmSc86w5t9voA/x+G77OKamTYuZVb5iRy3281IG96JMfiDkA73cDz7DTh+6
DqMpvovbFh6ho1DBVEDn84GzX3TawIlCRAHtbMYesW0IMSqM32ZxZzCZlFP0SOK0Sg2fRJ219j9B
63d649/zn6hOSdWynzQtKGxhQ1JrX482cOOf3jfKfgFBkvHOxZuTKDvyoLp7u1dxqwbouTOtsQdE
yIDHxhZXnhFtmctkRDkjVAF2Wmz9KLUE9yiAJ4MQdqmWONexosyMCWAr2Ghj4TDkUqQj9LzT0VOb
u4aht1gMPAghemh7Cf7lXFcFJRLMjZwrwQFTmyJdUwAQfVj5qUxpcA3vCedrI45EPDw3Sb4f2msk
ZclYO4h5TEfJM1+eOEe3lYYbPxDYpysWTNfCKiCoKlQ/51tDwDMYTZOD1oRMNXwKovz8jterd1Zj
2JlYNzHej2kJTwyfUdqxGtyJP9uIQsrtpxJDskeJ/FqXJHZ8PGTPHKGD3NWEiXY/6lLaqbFmURx0
TBnUkJetLzAIKEnH+pm4Gf3zUEg4J8o2JTCV3LB6GHfEtbiXs1sKwAc+DbuDcTNKPpSpPqRskWJE
kgyKed5ma87CBBPNW+NS+yviPENxlBiriAn43Zagaf+W9OuQVS6reCnvOp/24oC65cYYQAdSAx+o
MQahhXyrpFTlRtlF4ktLLqeOVqeAPwANZnoCSd2DMDWSqmB7DjwJbjckTK73jKRH6GFT3iOUVc9U
0IHWpmaPNhxO7U09A8yWvUNP/+D7NQMIRyIOsiTUJzkgkd2Lhrx8QLILK9HgMz7kIyuQ9irXVsCk
DaRz4b7X9CEozs+egDyhlCwZpRbmZUW6xiZATIghW9b2ahAEdxgfaBGJU7r/M5y2CzKSdF7lQszo
peYnzGGtbBUrg0vji0rWVlcZoTnq09mJcLyprEQTTzP3tAWXd3MpjAOwNv/Wbzk7qUVaDb08qb0A
I5L/TUlCLv9xNxx3sChOnrt1fV79FeERgwYselvJvFiHioxdzmC0xIZdeXy/szVxh1r8c4rOFYrH
4jHlVr/iMhMl9oND6UdBqYlJmad1hPdGNZgXgbt9epm6kQmPXh5tN5EC2qrGaezJbG2r565cArrT
cYvXUaeiHALmmxmaDn5y32WuiiJBwnax/xnUXMe9r6Qa/CAuhqnsiDdc3I+DNCX7yeaV3xqP4agM
fsZ8Z3fwzvKJ2hiX0QF5jg5elj2KQ6TkcQbG+iN63j2rzqQV69Q0FtL3vZFjSM3+KI6VM2/Y+Nu4
6WfzNA+jVH33ZYEoQjLl7Rgc5hA5GKO3w4RLltQpbx/aAdhgITkxOWFUg97KipsXw61I7P+9JJoC
8z2SrHHngnViuUVWGW5U2J94mLWZzvI0Uh5DGaDSgQmVzzBq43GE4kyMYsG8PSqQbe4iinESACPk
QmcfCBDvBHM6KLdValxAWp/TNZa/qupzB8rvDCJqTOkSIxRLTKd5k2Qinhn7k9JpI23Pn2y6nVCv
diJUZbZR3dzNtMNAoJWmgiI7X4SoThn2vJgKPmDVTF0obaku3HWTVC+BF6vgaJzK/miGzXu8tpTZ
yQQhk2VxRqXtvF2Z+uyVIJxlJGwO4YQbAcjy5HmyGYP1DecAe3rUVmbp7vONNkWHPOezY5SD6efM
XUMSbija4K9bQOTNcDxRzuOL59/XuP7civ83wG3LMyXOH3tz42BJNUDrtstPculx66x3toebfWk0
XQFu/jbjk92J1AUeulrMaS74rougxI2mgNucIm3dSWlwruOXgST4E4xk/BXQQQCNfwDLNa2Yz1GJ
3a5yN5/XCfB/RPvPoAUkPwyPBwWlxAV8KmaKgbaATRDIOKE+6ADit289t0941X5Amq7uB8a0bzHu
DylLO4SFdyukIKTluZNjpsdXzZnZMhK0Yq4kaQPOHRak8eMNbqSnqeHE2yZCVR0KfPPGvi1cD7WG
dUe2Mi8raXrPW47NXBF21SroXjyoxOgO+2EoiUcsDSx+6iFWl8ED4JQ9jx4/yCKkgJQc0pwPg1+O
IBwPwQyN2QmX/1tLuoVhn/IjFx+pD021TGSsWFcHgGVlb84rvTi0VkBmPcWtxMUTSg755KnUSEB+
V8pPO4m6EnJGjZYTcB9S2mXqaocvUu0T56ptWCeJFD67RJTATvLSkxaFlezVHBAAT5+IA1G30njB
ItAWybfNtOx7FTSrc3L/XH+PU/VgQOvhXFUIc6DE9FNJ+cPNaYMAnq9CbvLIbIQIlAxJfyqi9bUr
/AW/V70BNq833k7JPWNKGByWLxEH8zJtKhzd0bOp577kQ6Mc9UyYG5vs2SIBcqSnNjiXjgxb+ZVB
5y0TjQMnWjMakxCCnTVyua7MqVdvFu9G9oyZfyzFiuaI6OzJuUJtJQfERe1V4ZR+XnxR88b6ygwq
ca1JXCH4SXt9Mj7UGkLMp3D8MVawVtaYlaCRXqj5hFfB3kLmOr+bdtqpA2sDFoVez8dZwooidQca
mrRcKy9/BzbofNkeLfcGW6F9gUfMcZZYvlHtxg/w3DntAqrKYJRWEReA+ArO5wnj6N327sAgKPfa
OeWF0/9JMyHbAuPoAv+rcD3Hshq+hAQTgYCC2NVrvHk5xUgVyFiNJ/zAvYxe7T4guDY5w4JvJr33
Y+ytD78vt8aDi9L9bTZsWO5P4+Qmnjrx1k7aK8pFc7rDTJdhRR+4avQPs/yzrlxa32U77Q+rNGyw
oSSDltXgBTSeXeNe4y6M0gNB+THVQ8LdT3hGvARgFnaEkphrEZDL/FYQuzduIcGVr0zawK7qq4bt
pKOPWAyr8OKJBQluRP3ENRrg7JovDIVOmHTN70QL1knJRHPhErTYFk5iUCYNR77AzWk4M2h8u1Lp
Pdx1pwv8rGoXg9UqePyOcFvi75Ig8o0pYt5gTuRaB0t9oruJ9XrAyoglbeLhO50oIcwaK2lSkCRf
lZRTw2aV3AG6ZOLPUyye+adbTPnyxsjtXzjIY52taVX7H/WI4rbSwRzya17qNyLtsXEa/uIetjRw
qj4JRV7XRuQAr8ODQpZ8w4kkUOH7eCxktDJ0OP1JkbD7azCSYeSrgBXerWxTIuEWNcfV4uDjGEUX
rfBcw8cHBsO+3OlQ1bvY8ovQwqDapBpzsQMI0lG3xciqDkk9/ZGZWAAhTPWwOK+dEszs2iCWGnON
6zohUXaw/4YdmSYy4ybBA88b1Qt7Eurpbt1XPEw46wv2U5uonbtfx2l5lE3VLSDYKeDN79peYx0U
omzlF/tg6jHe/421GCVE7hwNZfBLkCG9HDvIpb8CsH4hZ/Oq0ppmK6BSg1sdFYgdBfNfE3zSVust
T+9vb7wvb0lxTHJW4gDwFcjbjaFjKVzpbBoIw4Wsk3gnU3k57HJj8BuEYjwWMF0Q4jkaZKxCQkGx
SU4bz9BU1sNvMRP5X5+HlZSF0gmz2ld8h0AmEJJGIgZsnzo+mgoTtzSnnlJyMWy+r1gjvd8QSLUG
3XzKjiVQahOBHgr/oS7mJBc3KF2VuL05s7sxq2gBa+ftelaSnQHniaZF/HkCkkPI3g+ApGPgiWvz
Kjx/drH/r8MBhkdRBRTE7Em4O0c8411uRqpxhP33sDrZQkYf6g9ueq+zcZd3i/5X9KJZ+8sdpYWW
bh9iqIeLD4R3VOfgxC2uo/v/UiYlKoklEvZAaOlgYHDW2QEANHkoLgJQzBsRI2zD8SkljY1buASf
/8fSi9tsJf6xh2FQT48w3V1ORVxQYrGk+bbp+yavY857mH6xjNhOe2ZTin4PrWxa5pebAxRHoj1f
JwFqG/Dqy3kuSgg7y/2GV6U4davB9kFnY0ImFS/I9nDi71MsAvk01I+7s/RvGdZTNX3fcgyIUlrs
UEhn5L0qang5Q1/+IDy/D55Lg+F/v8FBuv1BdvHFCXkSybOL9PymTt1+E1avq1a/NoHChehtgRYa
GFX57BN7d9tnc2Ducov43Kk1f1LRJOzKr1MqJ1TbVyCsla6yu1eMQj+k3SYgLOIVXe6+JEcL3UeX
eg6elm7STTcS7AGgHVw2uo0se/1LXS+ws7nMxTnGPUMuNDXY0MwgGVVS5CRwVCUUZWJWIxQ8POdV
dCAoHID9D8XIuIIMi8WvB3A9wtRjWHJSUMErfIbNGD4gAqrXkpLQNgJZjuB7PjzK8zaOHm/e+DIe
Siwf4kpDgNK3FtUqdOFBK1Tzm8t1F5+fvOTiGU+JEcnP2CVBXpvjr1W3OrB/xT8W6bWl/ZXW4hHZ
At7PXMDP6DDWbWbO+qQMnqZAuzHUw+Ca8XWfQozaRfV4vDfkKGn225cedsOwMSaNjgDxs52bpixF
g5txnMZsS3w/5vF0M9Yo5adeca+ksIDFgcucEUFx/YEMOow3uOGYAZDAv69zjVp84TmOF6eqJAFd
5R/nePdemSgUq9w0G7rOJM6zBBN9T8zJ0fdAid37FNy84mhM9xlyV7S6x4lXo+zaAGVjVnjmW58r
mgVNV77luLaBayzJkHpFe6nXFN8APnyE1KD0mv834MSEiJfoOSHF/YdIyLisvGrW6w9y35duDcEw
LtwhTqYu+nDliN7+IXQ80e2/ifV487ul/GWCWjE9bpUHGUrrnpbUJ2YT2Ib+utih/mO/NxrKxLb3
jH0JcFV6XirWnjjwDmsuN4z592D9bAhiezTw+wcRIBE709mdYroC2JTN5oHo61cN4DguKnHqX0yB
OnvJX9BJCa/YIDT7M1MslepWihL7wtrAAbNChhfo3/xsvgwuzF/qHnjWWa6TByj8ireeP6czAD6d
z+E2uH50D/gqd12xeoVSST/vWDzAlMhZSY3M/4Gzwe601SxRNKH8Mk7AD5U2tuuE+EJbJ1alckSy
xZV/CblU5EziJzHaCwIK3XJ0REgOHRFBZpZkkc5Eim6Gku48toec6OEBtdfNd4Mtpzq9/9cII45x
HDn3Qn9KfnW1gsjPemvtdjHKXckeho62gBj1z/oxuieL3oSO7qZP+D8Pd4KrpOqFmGkbK2zkJTd3
TQHL5ziQGVJCAUJhSN+e0U+oGJGPJZHK67KyMiZxrbbczeYR2Oeb690DnaY/kSI+sdmOFBiiv8wC
V+Syxtl21ZsDVv3vdHMRezyvbcILODXsA5F5BmKfj0Q0phrKqrQCqbMYvNeGjQmafHTBubLWrDza
lcykbpWLo1dS0YUaoF5EmehH4Ga5mwYk2JxAV+pUsURSOoTdsR7vurR3e9vZiKk4xerK3fCHhyjv
fPF1s7GlYBb3k3XXqGBxTWB1UGpquQLksbt8MVWEvcT4VvBP11gaA9GmCfBkkOCfT1J2VhvOqfOP
hVtWOYD2KvENnnaXTfEboo4+WySeRTiQHXhGFfJBPW9nnPgYzEhlYA5oZsK1BERnUycjlD08W9DM
AnkdASotUH1n4uf7Xqp3GlL7nWNyFTz8WzGfs7CAWQxq8yivlZIqKBllkUwRtPwvttMDcQt4ftXA
QbeE7biPrSCFlFxMLDLlgiL60BJVt3o6aEo4S/sYwzpf4PxIUjD3V2M9Ueiw7B29AJGDOMMd3HUO
8IsDvhY5zm46jIvP/XK9xH6IHGxDNI1guMu2sVAMRXihGu6D0N6GSz5Asj/5WuTCwQz80XkUHuIc
WinK/82M5JlPXnJaZo+SPAnp3XoaC3raWSGC/VrTtHmDfUkRdC2tRkJDMvjmEhJTBhPbfp9TnPgy
ZVcjbYMV/qd7M2xinE7yTJ1tCUeUiIGa38x5dZTKX9bFshnzRxxC90Vuqvvzk9fXpR1GjkLgG8Jo
cfM7hi/PkEc4v02mUdt7OPH6A6eMZ7o92y0J5lZsnNfXsTkY/uQ/6j+qdsMWSMKTetPsuAT4i7zh
beu0TyXKAVr1MucJj47FK2FG24zLto2DYF7OBAB3iAA31ivgctUUXw5SMGPrqo8fm4/V+fyxHubb
87cNrYjwwLwP8N/uc/ChjYq+AhZF5ajUPyvFsH3lgMACANXJfn/M5U86/xIs325+6Dq1ORZL+a1l
QSV3mLS7t0zXkzXMjLLB7zc9WLEZUZz19SwINYCsuM0RKsSH7tB75I9s4CYTJnwClo+AOcRvlTut
oGKx8TvQA7p1CGt5WzEpR2eBxJAb5+/tVolwtpgwoipLbwb97iPFZorapoTeSEP+XIVD5rlCm13H
ZSOwNrwIop2bL+NjXs5QnTeVA+e9dv9ZOVDHa1bLGzKdE+tJSLodLB3Y/gzUUlytCd2d7B/qB9Hx
tF4HKwbV8yVynUiHuVvZoc/8gbDwS5A+kuz9PfV9jyAxR/i7ifrH/MPB0+7EVrHFimP2ozU5nGQZ
Yo92Lq6t62dd7rSY/tZtPqys7mkvBNrjj4tQny/Jjl8KllZCuww/8tOGXZ5Ip0RtvAfmXnpqTbxo
0f8WYIBjkdGSCSBdo/yCqrvpvW7uhpBTa8YAUlv6AZXFRJjhWm1QicqfZ2LLoV1MMWZREs6uVmTZ
nG3IyCJcStzbCyz1YYp9uNTKbVwIzBjF6gxMw4SqykllkuB1V019u1krV9ciR8mcXY9bAzvOfYPl
3vcoopbbeSAiZYwOMQaeEIy8EjEQyglrsNZS5S8/OFO4LrSLm+6KhfPul/hU6jkFgiBTxetzZIOX
OUKOvWhPGo7pPFhKzmiNXMkgik6uoQvHL5oQjMbjs02bUkNLcnKGgJdtFirI1DfRJY9zeNlMIll4
mycZE1ITCCuvx7t2PMZ820Wq1sk3gYR4Mu5yqY0WjoO/NkosQNic4pTjm5H29SGW1hjDkeUvzL6N
6WbGRTA5a8NQKwtpuW4N7kkjmmWAt5tyUhIr6D/Obz9PUS95PUP+jR9cryucbKQz7muuYOQjmpOa
aF9L083RUBVXgC/mVIuV45WbCaKJUiGyRSLyZIP8F76iL0MRYMgULDivjufCz/d5KGdjG3KqwLAP
HYGRvQksICVkOh2iITnJKDc3z7XzeoopuDNlnG1TCU+t1URB1CZNNsEHkZf06XFseNk33BpwKCXz
0wjhPyBjzCqTv8SM3vEDcGxb9p3QurGH3aPYAyExWrpuQS5S1YKFFmQGvmUsSWnNG7YcgNlI0jme
Owe9N0iaMfY8nk3VYfMzktxopKUEBOGS8VYXtQcAuUN2LunLyg+znyAxe5dg7682AY/w4d74viHe
+yPC80lp40fTM265BXTATBDaXuU9hMr/d2ETxeCIgJHLfErvaa4/BaWq66F6f5BT53wRS0Hzv3zw
gPQCrUunUxSKaxXUwIGrajGE0GHy2rPx3LEr0VMhd8t8iWTGiBafmscUPUt4//vH5WJS/4rhjWLn
gM8ramWZ+odjgvD9swdYXb0k+nyrBQzpMrIm9vGXt7qgOIQvO1bq6hQ7VwKNjH5fiPT0K8RGYzRi
0FrLvEm/50QeK634JjTPv4gCnKrZzG8gfm2VSAfpKuMu17s7cXhMr0kAGI04/wSgcbG8IiZkQ/B0
3d0SZx7HwhiiWCG+FUbgPeB13kAStsV49PeJDW+/sRGx3GTa3yxxZSD9wDJ2CGYTB91/wZc8sw2P
hiSXN/SazfbFAto+nwOzOkrzLsbHUkcvU3GFIE64y+B3qHvpQ0jRmHyCJUCPAi7eA07Pm8FRhKLY
Jmopc89duHJBOMfGRg3d3hV4t0SuBGRtsOSTmTma8GiuLOCs6r2q2ZidiQtVUoVa4Z3E3mb2FanX
OortLLDLSe+WZDSwbD+I9gXvVHPHx8hHHcOFg8cAdJyyUey4ujqUIxBRnhPg8bv2SLV0LGYkQXY2
U/Wv+ozJw8VMdig3NNXGD10IeqXptRh+JOVykTfHRdt1bOc23eq68GZZT0NTPHizt2/FvNH5Jj5a
0lKL6RFY+BRjgxiDxy6A2sFAfJCvHPwXjOI9yd4/EOcBZlr8Yt0rXlx/IGu7R9v/Mwu9Z0srfIZg
j51xFDKfZNJurphl4cah5BID4L5y7gdM2Y8fLe2U6pWSMp7eKAOGPZF7n/rGEiOjeGLBfyP8irkc
/ImcmKfRGmJPp+wglZeVD1UXMmFMcKQqOhpnD+bS8xEzseCZKf0CBz4MpRpivdG2E8zY9lxvzT6X
X8Sy9x3TxQBmL2SZt8QOlFIuxTAb+s1BgAQNYegyel+ETNNRoR0W11kIBKCwDO4D/YyBBViDf19e
M577sZBOm4e32i+1NAYEq8kbT8lUbIlisLZL5xM0MFsj9oCAcqF17FvFj7YdTdTbZYFTUxq8ZeeF
RqbmpEhmk7CgpZ3SUMCTeSVGXrrGhVowTVknl1vF1GHtdpIU6BUPzcjlhYTR1Gz6+DN1XCN+M6NT
jL2levtYKSOjVeTbavfHXTiWCrFndHmK+RLNsZPd+ckH1UEQYFoBOXqoPImn1lXgYYjh8LQrNrW4
9j1Y2XMDMg+fqRhENRAXGa20izHUPJjnKGcvaheFUYyYBihR+OYqI4fTqnyegeK+CxbwncB0leiS
wS8dM7OS/RImOZfiHbTTCZSViMjESwck/ViaV1Um6eVN8qus/PN0F3VF1yf3bJBzEKJpbHZeKwsW
8tOpYKk9UaPYbm4E7mLp++MEfW7j4mNgO5BlhgINoadkTgbCyQWNtEXSM0IpFJCD2FgqdUP1YInA
MIG6Db/hKJdPfox4CBEUqPTg8C48ulyw8Iz4dC2uvoXXcnVyuegRz7KR9+Gkmg/c0pfdxd8jKXav
Vha+VEQPmcw7cLfcmt7q9VOkpt8bSaxZxlqV55TxRqjBx5LgFMjnakAUc1KzALfzHJwx4XXxnnsX
JP3pGgdFcVe0qpqReAEG1+PsysdeZyy1IloASo+SlwkGN+lrkdX25tmtSAhWtsEzspvmRZK56wCu
xLIGSjUxgM1+KjSL+FBBTk62aqx7Xwbp1Z0dzPQS2wTsC8XFyJ7rLEJhipa/MnmsnvSn6zYhfR4f
HVbTVwaXQKRxWxIjebPQMbhHBezyPtqYwc6QxWUfY71CXqjLdpTVorhLSj6ATIp/cEWk8Fslfl2z
+sdsPpyFXwXYPkAxfiBC1nB8eL2Iyve3xO+AzrM7r/mXHdNZ9PfNRn1bXvXBNIuqkpCbNGAzes0u
rUx8qZuYmTOqTDrWM0+NOsSGxgMQ4bFBDgvxEeu+3PUGJ0EjfM2ndMA9dUWlYdKK5QHWobunn18R
rcqOOoTYbk2DHILZ4jP4kn8pAVTwcJQt53JH06RnJnrMVv6zmCK9ppjM7b6UR0Gx9QO0hq7HCjSS
ENxWjJlFFrKY7Is8nRcOCcVX/wEgMy+vrrF8x6J4z2W3vix7fUXfxeU3hXFnm3MkPuVTTMLJ2bcz
52DGVvhsvRk5n2KfNLndIghADcbER3CvqFpP7/+ZacwTu+uKFaTDjjc82TXDlMY/grE6yPCjjHTZ
d0a2ygsdLCk6Ou4exadUimRmwNflKI4kBfd/RhIkEebdtUmnsxHAb5fE0UWXYR5vgl5LFBlO+Lrh
3HZRqc3FXCc97tnTFV73XNHj8qjgPAmXWoPjB/dKXTFGpcYeFf4TdB/T6YXBugZw72VtIVU77OPQ
kfaOcy1gWeqAC96Lg3trZMYOB6ED4AoWCFxzNwqwVM/GzIktPX7TVJhZPrctYM7YE0fv7ebXZvQR
9Wg8yUZ1mGe/KBCAKL61jOUQa/CAQfsrtJoRkakX2fi6c4sQi3VY59X30jydVfS1umpTRPwgmfuL
4ToGizSVrobzPoqc/k6BxdiE5Kc+F3q50yQWpE5KfhPWcwrUfI0+x3UxtXeuRsI/mR4EcmesnSDf
eSUuvYnFp67r/g6MIbQTh/FQtXtpSc9dnqwutQPlc9q+VEmdAABjjRoJlhMQcvNqiPNZfk8MR9Xa
/PhC59P20+UMJyB03yb0oXuVGcAIXKoFJhWqq3NpkjIdch9ae2gzZSdTAXNlqMKdA9WR3ONkcAsc
VGLUF6QmALj5x5qGqOmMthwI3jL0upz62R7BXR7mHv4/5zUshGtnV0dKuQFPFoMNZ8P8h7pclzc/
escxDu8YCMknlP8WDNXuCkeqdhZyWkrSPPoYS2LOdfGEcqMMdhNq8Hd8NwUAcOxhL0kvOrmPyiqr
x8xiEr2ZPqODBV8ndEU46Ao1qEJnhAW+WaGl+GrsI1gt89zXLJpOCIJmnkiD0+RHeT3GpcOSg5sA
fVLI/ke1lxAo9lV4sgllHCA9jJpgRvComVjcOpymyS1Qm2ZwWoTqPGHsmtaMVPW4Ynea588P8uve
kFkQ+yAoBcBpP486paWSH1zUFOXRM2tx6e68sDGHxXgifBvrVv7BkpQA8B8ArMGkcaj6Nznydix8
ZIesQ+yPcPlGQi3WRpCZ5K+hAA1NlirhZHwXn6EH8dI4q/PfF2Zvr1ffE0n7OiENmrNiXD7JhCwd
xRxinW+64taiTLj0aICVBdgKsseVH//XDsROXGwGBaYfLQQWug/4eBkbAdrUaniIXdKqmGs8WrYK
QI26a5avGmdw+yOwXX/8M48wFyeZLBFYYDS0Hobe8bogf3gMH0cN818SHE0CytQbqBSCVwcSB+yb
90Hw7HWni9gepgFEB0hwf/CYL7RSYRpH958QXkkDilxxQZis9u16pyuTuT37ZBBT5KVKJkZPQ3j5
XpmNTn4BglQsiLPF5JwgKT2dR7A3T0LdEOgDhH/6bcjuRD8T2CZurokdBK461xigNrWHa/Dss7fy
awAnD58cgBy2i0Za4E0yUux8YQMU2eSDHEC2x5WyIC/xyqcDB0Ld39yZnWC6jYbDiA1lbB+jPVMj
gAF2EiHnIOPLojl4AXkwkD3E6U95OnSJuKpHOHEl0ZJ1k4n33wcKNbjWMs3joSrT0CjcLeQ6TOh+
9yrLnWQk8uR7P4z2LtjYofshk7lXQa4F+giqljHNxGYaBCXSXSsMWDQ3w+itUVSzu1tmWJuUzlJK
URCillkERygK1HDSsfb/fsR1iiJUstAOp0eQk2eTNomO2fef8f1CPDTljrP8bnXdDUAbfOQiWFpD
6TLWUlX11lRg2u9Ln7WjUQth2DeevQOfyGJ4rsFMV8DX9l4WWAt6E/IpHb5L6hfaxYfeYVcePuZ0
a0OXtpTGrUemFdGPdS2b8Fnm8MIQZdxbgDNB8ZBT/L/jNziCF49FjWj8MbpDkk4wOWPshWEFObvO
cbQculTHgmqW0ZsnK1t6NyRjqiSuLLjkXg4wTJ+jkozYVYXUbBahadNhOGqzZ+XjKH7ib/+F9bm8
s8AgC+K7VgFpjSouTt0zH12o+TYTxt8MgkjW5HJG0IcsjKL3kQmd6GAJWJuDcF6/RZJZ+qMZUnJ5
3a7JzYTUca65LHJkdhxpbSt+sgOQq/v6qougosuVGm1aiIYWjHlRAUZgNf51iT+ctPUML6/Wtx71
Wne218s4XEgA9V71rc16VNQOB9amYRQR58ZNzhDQxPZo9lmPBBSAzzoru5u14NQ5nRvOHdcWLIuZ
zSlnCU23JXTZI2vSPFp9rMJ9KXvFEx0yjjlzzRf18/Wun/MMtZBI9FAhmaMXs1ahrsagUiKXNoHS
+7cbs2iOs4Nq3nKp5d+qoDpF48VnAFsg1l7f9y6kMLgGHj1l/T9r9vvrvxwaX2PKM1QiUsc0zfko
tEdheM9Hh9eIPR5FW8E+ZG9DQmOyttjU5yUyyjcpWk+zU6OKbslgkMKn4yVsVlV/S8+1yFI7lakK
jT/yFcWNa1Vq9EyRbQ0pXe9bpb+1j6izml24LOCovfHVXAWlwP/Eqi3HO/S38G8hiR/wo0wxru5f
C2EqIOcziFCi6dE3kRTSHA7O3qb/P2iItlMfb2qg3FnrpbLetoafe56xaC3/Yp5BzsIlyl7SDjzK
3lxuzTFQvL+yDbw195celwTSJ5IQrfq4vXp/9I9pL72aemnutVwuVxJEZ25qxwv8zuHDtwixvfae
q23tiU2klbi+JeEo9+SjqrZ/e7kUush5bFc8n/564L/mZU1LuaobGSGusJcr1lhAF8+/oshcPlCD
2Xt8geWgI1myha1KaVZ/b/r6MJAUEe0Sd9N8HkaZU8172lz3gLlCBhMhX4UWeIBSW6GiHGK+0rHL
fSMz0MPt7Hog6Fb0OY9o4wjadkdEjBdFaIXu/8s2sUDoygBmB0peeqtqBukcbUaAEZJZP3+gGMiR
S63UBLFX9J7g5h6usrM6Q0StLfWG6uPgm7tvK/s9nRyrFzt6zTGCrTvxOxpiB/pqGqpDZ/8zV5JJ
S64VR97L93MErGN+nmyLLXbHx73kmLn8Ld02zKo3X90OYoshsgBoUylifzqBZ/CFxQa36I3C/JSK
zUKq0WxpEjj8kAA7zlZcqzW5la0wMexwwlYA2CI7WUW/cu++zBbxs8RAReatK2SHSRtFnYscHKau
Oo8sRqhsahYrYXxKJNclOKz+J7BCxDC8HntR7Burr3EEzOxm5FTy0EpmmjLGC4OIuxJVatb5T7uX
vJQHn+mxsF1k21yXwsUfZkKnIgb2ibRpa4ubet6bajKqBLD08ty5kDT94JXhRia8v/JmQ5PEgY+X
DX8RO6lE7G6ExsNwDd5iz6OKgs8Z9AnT5oOqj+b6pFBlX3ErXR7PHZeWVmw9D+oHhcp/OGU4zW7C
J+jQBRr6NNozoetEfzFDC+hqTLbxxb+EA+wKtolYhqZZCg5YAydmRmijkDW7xCMSvqopYu8QI4sA
w6ZJbEkulnDg7DICcWSYa6L5B7gwr0coV2nB4PUzZViZOgDexn/wG754UXgQDJ+Sf3iG5c+Mzacz
XFV+HdPRZb6X4KEvB/aE5UbI6wQAbpAy4HjKJGAKDfJWxZAYef6kV+9BesmZcmmgYXrsDZxMjLB4
mz5urweFhmoQLes1Z2XMuPl4D7njfzBQ9C7ky2EMF7WCIrBXwfhWDFQU9EgHCQwzVfR91S3mv63n
kiTlNqCJZc1bp206ThLTY48UBR0cFBfZ/b+cp+U7BTTWw0KE0KsuEupZ6xbQCwfUVlJdTIKjWyqo
e4fZdUakw2dNOp4mlei0muuP5mgW/VEqrqKEi8+2RJ1xauMhukOk7/LWb1H+CrQbXR/YvjllVbx7
NRLr6CDTOdDBPPWNIrYwnJwvUOYpmMDA5CsuGsm6XNTmadCsRN1pMQG/A5OPuajX5esxxq/vn4PV
XloEoxuuwYrP4E4OP6VWG8rEcOh7kKUBsfAf4Bsd7tsAZoeIEULmEZh4G0UDBtVRqwIMrPGlmtc9
kMsvk3w/NaBgdQulh8uXC60bqQA3aqQorMPsu1DprTsPT9M1dZJdicB8hGF+c8CoK96sbCgd92V1
HKvzCGeqZUIpVX1/V+z5wU0pbZ9iV05x5clh8azl5lhzI6S/C5XmQhbOD+lU+oc9psSujyiaULt6
GP+mM921BUwS8LoDUHP3cqJroPLF5cNnOorNHz1rdCfUt7fixWn2Xk2Mk+Aku8uo262TIkHY9AoT
kqWk7WS30s8YXohGX5pwMY6IBfwqt5tHW5Q7XOLwFhQLTBrv/h+PpDaKaNZ6E89h7SuaRFWwzg24
ep98fiwIakg/pgWZtnKsehWoUXTVVCyoEJp7yCJkVqlfQhqgp97x9g1/8u4fi8AVOopRbtFPK58g
X+7osd8MBFU3TfTclUVPxnbQi5XbDhA9ZT67ZuLuKeBBIc3CsbFSex1CrnCzRI114GSf6dVuYvTu
vme+13JRGcNnoO4SjvKdCo7XmwfJH6z6WrFkLPPyQYWk6S9kBSX0oHD/OD7ffTxJTmOsgfSU8MXS
l8mKD5Cs3CIpmd5b7k3Yu4Vppz5OqKvPrlUzoFmwi4dQ0hMWuGHGFpW+PFH3JIHrUILQqeVfir5I
yWze0do1RU7ZKTzg+872YEJswygAf+DGCbbF6w+55ZXcC99h+60wsueJfhGTrTIyfX9vfKHCQ2Ts
8W8plTF2jhCxT6U4YZc1OdUYvkuGVvk5fYMcIWCtyDe4HqkI6zvVr5Vl8mnuPbpaFAZN0Ez6pkTl
mM2qb+6wweG2LIXM0PFBa07sNdivjLWkb1CRhHYBb2gQ28gx/D0WRHm9F5B+EM0ZaRUWBJpeIBsT
JeYRprFKcP3GZknb1ORG8XJbzClmuHYG3FcUt2uiQDDA+vVWPtI5zZ8pYjhMRxZOdLZu0Hw7uYdx
kg8PUiDfHxcaohQI+so9YhiMWeORiPABoVxxfM5VjI6/ziRHD+cOaYNTuxDUV30Zn45dYWA+OrW6
p0ogofztXJRhSYnAObNy7PukCsonWQj6WMuJYT5Ss3BZqyL5Sq62XPuqANIkAylywm42AW99wKFa
dvmJGD3Gl9S+psST7bv1GcHhl/ruKf3Tux3fXGvtDj+ATzMvQkQQ+iQ9mEPKP/8v/Xd3eeNI4Vyq
PMSnvgLzNCUF6bOIoaJj/J+r/3sKOcCfrncnb9G8wiiu0okcpZMNuv+VJTzKZh8VJ751lYWxkS6B
2MD/nc8zHW7MNoW04YxJ/qx87GzEvO61o00591H5QuXv2SWEd8kViHqm2aIue7W/nS3bbi1u/YG0
s0bQHbl7aFO8mda30zy0RvwLTFgDZaeaopPtwZI5GMWv4xvs8WuqAngkMQvfh5mlKeGjZnBV/Kdi
d90hqeqyUMZRNzSKLxnTdNt7J6zeGOEb1LjhedGtRo8x9L6D8nxF0K8M9RtW4V8Sgg05QvC1WxpF
1xhXmvCTPkycA3YyFC/9tRQwPEktWhMBaTJyxFGlCeDMowFM01DcxdZ97V03AurHkpz6jeVIC6+9
63LwkJ1Hes4N1M3U0cPCd1teiXVt8x4Qn/3Yj0lONROY3JzIRoJKef/VlrW/60e34U1PfD+oo21S
tdJOToR69oGVJIZOxhhqGzZnDqOjXiiMHj9eqwGQZugD6+iYDuIocAl0i0JJ/C8GF0hVnlb7u714
ylUZqXfyT5fgm8qirwqrE2qdwml/4vR9SzGTF9MHjhI3x7bitgubApnIottWgaGMPqKtXdlOXa7N
IbK6vOkEP6H4Om/XbcNx+kDFXJaSXuJvtpi80OUAJI3cQfHtTQ2Jr2uLbpaPbZ9zGowyvE3xVxfn
uYGpuFMPNfJxvqfmNT/lmHDrrdjYVTMfHoFLy7ILVyC8Nr6lNSSZaKthcIx+iV7jbvi2mP+br1XA
5KBnj/tZbKdhwzzqCF+b6fRSNjAkS/B4wIUb9t42F+8wM1g5xT6JkEkOdZuxt1ERvkvjtIHnap6e
fS7YZ4Om1MxS8Ad1/AxJvCmEYFpJsT+mgfe6/thsGNnmA7Moa5PpgWEQkHAkncZmWL0+0WDHx/ve
TwWX1hiw72YGj2LibaAbb9Y0F91hnmyY8IyC/IZYANoV0yEuugn0AE1vJiL210inaSSnPtZyXDt6
0pMTVLwDDO+rYqPR1rnpMY8Qx13tsWUvcZKnpOpW56dWQqVAVUV1OxRbvupQ2fHyjbjuTiDWzWXs
C/O8S1AlSDOqfP2Ox2LEwwp1KtF52JBdfyOz2aQbt3PQ7q20RW9rgP1nwEmat0JVmmL9tql0cmKm
LFGjW8sb+pfhZyUq3QMM+2RXHoHyA5JUwVQoYJPO9BjbF35BglaQ43S27YwSTNhPkBjpfZSUTwLJ
w9hHUyOcI4bnXf9QGK4CzqyVQgY60h2G4WfDyG+qY2hocH1KjbQyzSU8k2x+X2Dogc2P8X6yvyF8
B3wNhy9q+Aq+rfICCnGuoHWyxFmo+GsEFWFE4AfPuj/XJoXbKfTg95+gDgHFCkN99et8Pj+l2jX8
TMp2CugcZia4SBC8a/IldP1gvlmOx+2p0rpG/phIet0oVQLxxs/AqhSEhzU9IIGymzvG1pebX/LT
hSTBsBRZ1lHadhmj7IjPnR3B8zlA6lTqmnFmh+arKsfYGhnLze4qu35ZGyxJFHBjy6+EkFbPVBiI
IKf+6QuY9KQ7jA5odULGVnT+uTsGbu0mjCaJcYSmtC8utqhLEDelq+igNPji68vBncRB+Z4yNdPG
KB2yz0uV/OLlZg2QUIfMp+1dArUwJ/+ovTjcWnh6kKDERx2o/Z+2s916Y8Zd3KvDkWrIe7FLjE0x
H1cANb8HXJqan9std/oC8e6udi8AdcZdocnRyHBFy2kY3nhJAbpWUFTx5dgtQQwiVhaFenX47v7N
yvFPqUqpG4I+dqBOsLeKNlLttIHWFd4WAnKBWW8tAqsm/ZchMdAsyH5lbIB1ksnG5kQSIrsBqiS7
6nUl72OCW/q7gu+Gc6njeTmSWSpIqK/sHPcUKyA8BrQ76qSKzqJgLgnpcd/pyH4EwSogxpMi9wtH
ucYMsd0wCrFu2UTisAbW2PQCBokMdRpvQ1so3/ioyLMOCgCNh5hcfXIbaHR4CktDJGSx9+pkfW3u
g+9RXmt9HWEobEKZsAiL/xDvsYC3j2i3A/feKych/rYgLGJrKvLCr+AySxBLwTtZdYX76QjO7jj+
K/hYFWRANeKjAzpsdw1JtRhClP8+5RTTQyXtSsjrM84COBAJZkrqY6d+5M28K8KurGGnIRhSmCJs
/qCLwpJXeRmVsvYLhbdTD923di9468m9KLWWvRDH046WwMk7+uc9mYgjnhU+VQX97irl9fDz43eP
5EdKEC3kPNtdp98WtfuAp9I5SFlDlbSp+pPuB1nwB5PO2RxWtZV5JauTOHgeMsD+wkL2vUc2FBUk
AhSqAiAnesoLKHPFx8GS7MkqrjBGazkl0SDpWYFql1CzWwet4OD2p7aexFJeyYmGJ2e+9DAo2zg1
eoPB7i7YetUmhvI6sDRmhYGqGoEWKmWMjlYSWQVwsSGA0G//b+o71Sdt2AKMdUGtOPRqmLzb/geO
rwI/PSNurMXh5qxYitEiB0xWnuclM7DxT7N/qFUR9eYqA4rmc1OZWiAU4sAFUSCa3+uOFBkM02d6
Pxys6fK300LmZhx1rBfFm1PwyZ5bItenq/KFAhWOOUt5omQcOw8SK2SygAnm9tMDRdRpfAH074tF
Nsjp6YvLOVJJN17wpOGTekc03FSMF0m6qZxMvSbFislYhJn630A+geHUAOG7iRTx2XS/f/KAhmU7
tKzTYSckQuw6IrkiBiz2u0HMScv/jkBMCDreqjMAlEh1eqjiaRI4yvnuLcLb9ASruPSqOGM0H+wL
r/k8uOkVUnl3A6YyylXMWAxvuBCiQs1Gj2/wujzqsYK+XHSsDfOqFUJMAAAYeko6HFhLSKr1/d+N
Js/G1Xyw3O+KcBjBAPSjjSjc0Yr9DjWtBhsZ2ESvyuWIR9T2OqbFcCFCM/SCrsv6JpU+TYojKSSe
S4PHwXiN+iIDTlmdhUV0uJci6RL3IdgOZXPBRp8s3BwjfZCqYA3CPEoOcgtOL3nSCzpl33ItvweQ
PcCn4MYR2MkTb3dsSYJ4fgTUXANpEChm/6ja5CbXgOtXXxvnkDM0vkfTI8+PC+Bh88kr4PgHImUC
kIdWqjD1PVOqNWt/25ByFN65l9p83EEUI/F1OrG0i/2v9TbxhJzq0FamsuM2kapYA70liccyzhWD
n9H5ysJvLbO8UuS8ikOsQNQrOfjcYVI60j2nJRHcmcuiWAeuVEcKtxpU56zYgaruE58MWagHgS6r
QQ/5Zl4TXO7KAn5Phm5zJ2g2GDk+k5XButgCDMMdqcLgydM5OJZ4pzMaejHydwPaaCezUu2n9A4H
VK+ElszsadsgxhoLZR8qbcyjRB3+bMwzBtWIe6/mPUWR3iPee9zlAHGZIApPOoPTtRl3JyxVGq/E
IUvwC7cRICEoFuN785q8R660dWNxah2Je/5eWJX5zMSYWx3lnKfG5P0Vy47DRHZTCl/Yty5i4vd4
D74itc7pENhjr4NG2lw7ouq2IOQMQ1L2R6cBjb3LVKT4W4uHkyjhcbuyRaqVIahAa1k++HpWDrVs
N/8T+Cho1HESih4wK9jT6M+fVl8Mqp2mDhFqOoOnjNbA39OxWIS9FvbNXb0zPa/d5jOqEWk+OfPS
I38IQ/IfE6mC8S0dIkvf0U5murqOnE5+xwK0dEX25Ddpk3ZvOqr2EoVpvx7koA471o6Pt+hf00CK
0KwXXCZRBk/81U/V7KpVXQpcDF54maUGWrLDCy48vQMX1es6bjglAjkP1udCiEWLskWtohp1+1+e
RH4aL0w1U1BesmHP1A0DExx12xoVCRnGNMP+fI9miHcXoz5q40jnyimKpW6WFCc1M+wpfrJi9R1F
zLUrHo/E+Tsoe1WiA+QohrpJtKSR7z4rgC3XuzbiZOpWVFbuMmA2wU9Qi4/4ZIkf9P7XcTpgiRCV
Rh/alNZcgbw3ZZQ2SCCtq6miQZpvsuvTpoffPhCY3LKIuKobk5m3xE+oFUR6YBWpAD5dRVbfIOnA
MzkwUbgXeG01l1JJkkFLzlR/j4JLHLL6yM0IU8Tedrt6SVsr2vq3/G3rtmvLzSv+RUxy/XDt8kAc
gV8VJlMfhZ3gyI1dROjygzhwxriclsI3PMawejwowxOiXpRALlgJpxQvgUDSRi/FAtgVahZ3NSrs
b0wyvP+meRLiYcTSiZh8lS4C5l/F7j3b2WwaGS/rt4Qbg/Va4fIbeiZduHtwNj4MDHsHSLZZeacM
FvQon9M4ZdHPPstKQy/zU0nW9kuEKuNNKYqYJHAnKG1BFnC6UeQ6RLIwfPxWlj8QLcYzei6IYAts
FZycj6DMNsAGX3JVDVul/f2MlZSMPnKth9YanhWU9rvwXrTvsMvVguLXATL3RO3QqOgygWhUWHRx
jXZInba/GP+XBSPnDXXoASEwEbL6PnhX0qkTfzGcVZxWUIka7Vp6PnrtZJnEC7Cq13/teD2qiIUw
aY6+xwvrrX5hwvdv8i+vpfQFyFzWa1/2X0B+zRikQW8cPThUeYufzgbijsarlBitbxSj3N0STv9M
pVhDpwPSCSqCsTdcClQq/s4OMdD+Ig+1qNC2lMOLOrATNFOG9gvZFPU/sSXjZ2PeiPRrS9QWom8n
BT2lezprHXFyrG2DkGKiheovrN8DfZHS18e9fpwW+us5rdbAA8qocjzPPiqYAaUkv6+HaVHjNJDc
oZCKXF5VM/1dF0kmXYSOkJAJz13CeNJl1RYN5TXWEpFg3zJBnjGeTURxrIKPGphtmlzIMOqU1By/
FyM4RF5YxkT85Z3a+yLQ/1IDy2PbTTOY3MXzuEeaAQhicJ8NngbBjBg8dfEj/CB2Ejhx8idSIsTO
cn0gf/4LBIjdo7UGCt3qSrTE/t8e89fONyFYf86fPL52nQp9y6CZ2Jjy0Nccdgo09JC5WrAe7gaQ
qrsycZHOugjRV/GDs6XrSaAIaF7+FaFNVOaqTgTSuhPbk8sKOb8PDSHJL85zzDeEhvdgMjFU0bXS
UzQrvoZwxpvAOIEF92DR5hsbT93A38toSPh05PVcSmWyiPTWFblkAFLmFxrQ4Dj1Sxqf60t8AfK4
ESnyQFT+QqW+VXv5vtLQ4T2d7+YyFd78j7c3GYb3SblhDilnsura3uZcL0+Niop7KAC4CO8fbqQF
cM9eOCriPThLLBvBXm9Qzs2Cd7TbhW5nhDG4uHJHsaXP+RVx+3uzq8XFowDrklqX8nlOVBKaxdR3
VJ8me1ho85ma6pngruuKG7hxpjCDFedhfqiLCs4RNLUcdKHh0YyriwvhJMOzRzpXS/OIVQJUTQcg
zVG/0a7duYLsfQ83neELNF3lb4yaeKS5Wsm6oQHAL+RUyvCjVpJLHw6WiYKJZ1nnZq94N+GHcCH4
aOH3eor/al3nSFOjVtcamW4rvl1qHnDlq9j/u5V+sEeEhr1lc8m0cKGWyvaHpWrGRiOXuJV5d9JM
V4uBDPa+Vxzg3mt3lJXh5b1zgYzU1iWxty19mQvbzuskGF0ew00FBS0scWn2ex6w+hvoLZvys6NJ
90119lU+tNHOEuxzA8yrMbHgokoYOP/XGeETKwi3rFGFrmHFUIVPMmt2ZiKK7Gn5ZxYphOE2EmCI
2B9y2YlQO0u0FdJvPlhJRvB4C114f7AXJW3pZ9oRUA6Cw7DAP8ec3wdWhP53mwiWK3bQiIp80+eu
cU/meuEC7sAxMmTF1lUleJELT+hS9zxNOrrsMKx1We4RF1bx31EoyqLehjDcYN+0oQHS77bbQqze
+uYX8cCqasQG00DDqp1CvYQiHOQSxj3gbZtoNyMTQJnPs5Faxmmx9begGAm2jqkg/EQwxQrSaYE0
YORxRN8w+DtsoVmVzmKLfaLFGdWD5x0jlZW9fKo4y56uF4SN+kfha32Ta3taS1hy17ib9MuZGf4L
Bu6WgCnT6xCdPgr1Qlx9BBs7SbbjV6kYEhwaBU+T1GtCONHV6hC9T7xBmuDmg1RMXUOlDaS/39N8
sCaQICOtMkOk8vGzJFQ4+GOML8zg1DsYR/taiadN7SyQ2zhHhuZlVqyZs+6QvlovuHF0FHnUcu16
yg+nFVNJXiZnij7L8PzVTEormC5l7SbRGQdaLgh7xMksE91eVWFM/HmEg5AsvkaSrdmDdDdv6p9f
4WMZnk3sflhbqH1FRrxoquEIcQxqYNololQlzDrF56p6d02hUhFhHCvNOatYeAx6oDDGjYYeAeTT
xJAKNM3wHClDNlAMj7iFQ4nrYsP7os9x8FMOo1SMDzPnJlqFH45KYLgK4DMdrO98PVSuP1dUS3J6
SwokOcu+Yqw979Z1LDVve7bcmppdGvP1yPGPMoLUcdzc3CrrDrfJ4mlShMETjY4/SLtCKf1tRGbG
mTuZxZLkLhodizPfiTRpAAucvD+KUGpPpI65J5/3LOT5S9AVD39E8BP1d09oiSN/DidJl8l5Ua1U
eSHaXyrBxQw5GqmLBbDMdFX/9W1vtMJZc8pgkX8gyLBXLMlTfM5LC9QB+hI8xTDMVgY2+bMt+SQX
TThHBBj5+u6ULWK070QqDTTSdsIgrUuRRDXd+030q2mY21ZbndQMQgBile4gcYexdIDvINbljtSt
lHBoakN1cJxCoJVonOjCMGRALuD6aTVtmYMMgCX0r5gE5PdoOPY3GBsWRq7R8gag3l5kg+kl+8sN
cUCUuRQjk9/F56B6LDI7r+ZPDrPS0vc+BF4KlKiI7Rcp/MRR1eOVdgTchZUASpzmc1sHGm5pmDvD
EKB+RtTpC7zdwewKT9/VVTveICZQc7G0UQa75GjzFWc0d7p6XcEWFgvFF6ZYSxwcAyckwndfSZQG
Bysj0uQElzB9tf1dge828Wzu6MdgGXP2qUyMw4jPRLu+vkFDKQJLx3AL4giZ69IiGmLmPWUQa3uW
yAEBZTMsEAaF/2XGJDRGTnLzL7/Q/g7aUUT5DSBm9BDMuptbJELyNP6n6ij239+SDxFwK7xIVrfx
zZrPKLYkKq5TrAA9zKU8EfDX6nbMZX6k73CEdTdgSRmmI/iloD5uQwtAOIcyp0GjQT9DgyUDR2jL
merm/LxL7e1rTKytXLOhod3AM5BzPP/5A+jg4VnWIdIN248aZMr2nowvjQRNPyK8n3gemka3ehSK
r+rA0dHof+JlpeAaW3UQT3SjnNGMYitDfyTFOqiEG/iZewH2+RDsQET60gWZkj/CP8d6m0VP1Wh3
B6WyLhbSkuFv5S5IpEeyZr0y2PRRIc3TnEL2mpSTa9cXrLeh4lG/fe7BTcohiAW69q0tXUOC1Li6
+ReEQ9AWscWn1UEdwfszTnALUGok5imjte3vOgAL4EZgUgCLmul8XyMWREHG3w2zRSU0yj2eEMNa
591rOiaiJlY6rzkMV+wnUJacx70053zoydaBOAczq8xlbhf+I5vwP6GcZ3zzXZe0Aq5qRryKwf3h
NBmNT2k8EeRNCSmE6T7wf4/qaupArPEUbRsZKxHwCL3P67ampm6N5TWuhzuRVshcoF6IWyBZ4PAN
I8RLziwc4HF45z2YxqCVko93GeiZM3mHNFqej8hnmGVEMRvyceE1BFeJzkbHCPwckjutKV0KJh+n
y8y5yEzycUV4yyMaXSRd6FJp/jOc5s7uV2f4XIjMltqXoY8mApZtmpyMZrFmjqNtL9WPbKmwR98j
QdqpkbDLhE8Fj1AkAkAU2ilPIZlqKEA2JfP9wJQ75UoFZ6A77WbLV0khfCfGFNmU8oV30hP4h4Ds
ZbJX/bga9frPnr7cwttAoXnLEAvzlg4UObZSWdEtdLNL4UGDO0m/P/N6Fr12GY5wbton3mYd3aQQ
NbACjUDAqmEB0EaqK40XKPOuNIeQxAisJHiuGLOq2PGAnHAWwGC26x7mKIMSctJOc2ftQdNbYI3M
QdDDNgPRbk+47TN61bowtBfKKtHdgQlwNothCMmYt9/yRc/dsQVMFhsYaMv+g5RDLQi87hDYMHu/
fzjgsgDosFBRX3TBWGyTYXIqno1Akg6Foo8oED/mp2zfgHlxZDNyIqIAFVWgCvlN2MTlpM8FHCr5
9FF8nyOwSoB7AGISaYgZos5r3PygynFc8PJvYTs+Z8NYgTFTtv/0Qsfc56KEY+TzJdh44P3cAWiJ
47eBxRhYGZZmX62Sg102djlUXbHFJ8CIFgnvt2184lruDxwf6rnxJksWGuLDFXuxZ3CecO2AFXHF
vre07hMRZjw1aLeQVu8tMvAbSXykLtV+kfQqCGN3rzLUUiFt61B/EZea+kGfGs/BT3JXZC5gjat4
w20dyGE7NVrKp5bxK3jdpwFGgF5GXH5qvrmQ/nJGcMoFRmbX90aePKI11myoQ0ZQWoeKudkqqEOS
cTmIcCHKbcgPr8ocn8daBESnsNH/N2xtmg1ZepeKnpWcwHMaS19bzkwpa9qjj0Vcncx6lqxNRef7
kC8tVKUvvIOmTkQBm3vnieIVK00W5VG7ci4+2ya6BSYAmDey0hi98zYWJQP+AWAhg8hMRIh/EGXi
tTi8BG3WBuHvqVSYsH6+iY955zcm2dOgatNb6o5XsSV4/Ip2OJ7/sI7N90eGHndM8TYC7BoxxMgy
B/q7JjgPZevx6riZSa086p1OThgY9g26ouq44c2Zi0Pk+LBRz8V4qGJhYDC6vQsKjY9/qYuTjRJ2
Wll5COkfMiFs6RjeF8E4sdQS/qq30kuzntrBPYGN4scuLmaIKnto6SEdC3otnQ37ukDw6LIzcUHf
YvW4GnnZneijOVCSn2c3UMzSHRghFjaWKgYTT0f6Terl5dQJlnu05i7Wle0wVV8hiGj9qkMXxwnV
RkDXbbJSYgCVAYFtT9+97KwuFo2YidkGWgPHE1St3oFE/RHC7IW/xa9Ob/9w3YPePWxSMQ3CIpU+
IUv5zIGXMgAh8shS/n32mlLELW7s1DGU3a+5T6+yB3ZoPXjcDYMG2dcS4GYcBY9/ZAfPkxZmn6QK
3Tf3QbzfqNAXd/2IsNnzMTis+xqLD2CrKuUURHML2zkMV2ncGcktdN9/9DdcbuJ1lE+JNSgNGZCV
+cgTpbOwa2ygShNFqoet013ZXVa9mAaitzRapSYPaV377zN129t3xSzaerb7tKl3nW1qPW0KSp2X
OV8D7RiAHrM0UYWhk0hfmRrUMmdWgE9MdxjiG0u+ECafNIfcyaOUgI8k1XghLRoTbM5RiBxcMRKK
kQkY/ulhnlIrEUZ+89mOdYqhPsDfqpBusEBiGeQJfZAAetmN/XZSKfIQ0APOGDbUAn885YTCVZ4d
2okohRsduiQSSFFuT62Z/1ufet0dsmcL5+9YC0bkcXlZnPW+9A3xwVvMhEW1/smpURcBGPAy8vjH
lLZsKXm6XKICGpTJV9o6oPP4fF2WLnHSnrk5epSz3JF1a9dpqg+zVsgFygVyef1eEj1b6AH+a3k7
m4DsckyBWMqDCsFxRlYM+qSB6tXBan8p0Wax7SZ8SISP6FmOHO+w+RipLbYnXxduKtGiea45k+AO
411dH1Q1E+Nsfl46SRsTyF4m8MGgIGhChCNlUITylY5xvvJdRu2od7TAUfOb8oxVCJGYnB3Dw1wk
3867QrY+33niggaZpGJPip3UDGWANt/31VEvi5q3Itv+CXh/i+PhKm7wBjrl/2ljzCmjI44uJ9ug
Yr9hnUxov79zVmgej1UjUxGqrNnxGHG9/ueR/ITMkNbQBXqDv3uuJ41FwxtHpQ4nfZn5kRlmo0PB
MENrmT0i5v1nOV8X4dtpkrU6AVuGr2NSu0iUbyJjTXvCle4fw/yyEIo5G4Pot8n1/rkImxWDrFJT
bIWAHsutO+2Vj9J+ucPzxdowLOBg9Le1baMKroASItdTawMRFxYRPuvdyqZZ+H3DJFQme8qDyqU9
4ynqlI9zBMUBbYjqm/MIfuzCmP7rB3Ef22oXQa8b0sZajqVtXZGNTMTrYmybW2q/ITACJos3nO90
HwThMVVQ/x4raROG5KxzJDJqDw1R3cFkwLqdWjKFC76AiHleSHoJOp9siRUhBkigSTSPsJ9HckvS
WiuLp5LL/6tHr3rgvjBPi5i7L7L3FL0ZYkt3/tQE56h02EPDRzdiaOhEsAoE54Ob3by+DiDaYGce
3Mn9+Y62yaQBXWZAhqKok4zy+/M0nGCz1P5c1UOXzIL5HpjF9kiiOli5KSZuczrifEENHVmpZ3aR
41Kv+1orD8hrOMgXAoVFtPOT7ki07euKrxLc2eQvX1kobHeKy2ScbomGt+n33GpO2gbmH7C7VIH0
p2IoPwOMHI1F+LA34cK0zejThxpBa0OqiLn9sr8GAlN1Pg6+uPjxjHnCiYyopRrLrj9Bq5lmIOmq
vKOZPvgJTqUHUz5HJ5Y/ZduCaqKs6K666cFUFYrYPF3y6Py27rxuOg43LjvJmycCLqIlYZjswWiu
ZHlshaBiAFiRCpKFi3+1qiaCpEaBJFzhs6oDmPx/0shtMk1Gd8522VAu+uqj77nwS7EVYbmbDrzh
7ijyXphNEVcZRnNLY8SKAg8/5ewjIvLUb/kHP802+etfJCylc9NHiCIY1JKa4+jYn0S0v1G0rFTl
Hg641nl+aonIw/Cnbie9g1r9BPgSYgykH05pEyRdTs0Ynzw9FVE6HqLIvefm3QbYXS/OLvPwLUb9
WAg5v2RsS9AVdmV5/hpU6GSYbx6FmsGA1YToP9OF2Eo+hM3BXlWvF2a2zOXN9FEq++koJM87KE/U
k/cRTCJlajz5VQ6Jhn38PFzjRtvnmNemZ0t1iWwNRbst+eQ2p6ZOLaWZaOSXMZPXv+duCPfFuW18
knsPliFvNqJb/OzQhAOpBpZ0v+XkqvS4oemK2itfvH6SJPPfIEqd+lyXQCvINMvMLSc7o5Aj6tG6
6MYyrl1Wzdnuvkbz/4LzLwGejr1zDJYI0u+i3Jg/7qCiHmh1P9rpvSbrjJz7Bb01lJPjwkyqu5FK
LkK8cg1M0U4Pvw0/iv4eVY/h4RlbUiMjek/tLHAdVEjkeZIW7KEyAZYekV6xDzk9yd1ERpOefHDM
ztSGZ8U1qPQa5Nd+uW5AyJ726U1ES3QwuiWhFN7wjKlQS3e4BPCwXU3T6DMk3Gd0sNzwa3SNUm4o
Dq19OkAdMHopTxUqW5TazH7/GEg8g+2UNK6OzBpNseaWVaDjWyW7xscXuM3IdfdjnyvHIHbvwZ//
yUy71sIhhiMq/J5KsaMDuRn8+OYGDM6Bz82Sn/JgiMsVtMFNBfu/h9tAelmS/YKfrRfSx5sEQ9fF
ytYLJni2pVyr4UMQB1nJ1NE8ty9hp3uPWm/GoEECPq77WR6eGd2/JsRW83SFTEqhwj8eJDaPWVSl
Qz8c8Reev+b+xJccc5ndvQBL2QaBVKpb045IpgoyJKkPPnfKg6HNdCCck0qwxnSeXMF3bLHhe+58
79QnSI6JJ7eFyl3M2heP0QEtvuLmPmu5ZBasnZy0Dd3y12Rh+uV86lfMeobo19/rf3/PWlqi+5bl
9nbYfrVzNnxa/efDah50RWG3vlEwttTELZKLD5B/0/zzz9pUUfrOOPvtYL2hlBQBZU5Ltzgi+c9K
a6iRGFixm+Z0h2qTsrBK1p6j3Gh5O/8Fn8+vLnR4LUWvMky8a6rvBWCXXinrg/EpKewjDlGpxLOe
DxaCw3e+uLYs0AkJ11U9Bf16b5wcsHAS16+vdgqNgk9dvWtssZQlsNMo/MiNIt8mMAkFTcwPqsM0
NZvTiyG1SjmEDvyBbUik85jmJqw2oy/Q6pbPDsHXvxfo6pdNYsJqdyMcNTy84kg6oBZPGGYAt+G5
LWMewM3Kf1dYkO6bGAFaErjGy1OCOu/AtsjXTb+kuhS5YdcUHu6/VX8+inflaXBsofUBW/5+pNaT
9q7EZAQaQkMHTIvkfIvj9BqTW7S8W3w7nTr6t6w4AXYBj4f3A1rsArX1gvgrD5U5hfjK4JHPfZhQ
WTMEz1EKNDdppz79UqNxtbBpff5dS2SiYZsUo4WbFxk5Z9RwHWwYrvKgdcO7Xk7irJv7XqEGA5RJ
MOlS7m8mAUYSi1VzZNjDrJTQR74aSum6kWXmYF8OQw6Fo/6ZpOOsGtA0Q30EVL9Z091Ym4jBsjxq
p2ohhwYFKxaVzBMP5WanIUWAz4MaoZ2u/Un9w9RdKbHJVWUtIHDq8zFEDxTYExYqoQ5HOAyJUU3A
jy1Z4leqrKDVC2d2XJAyuy6Tm+EZ3JpvlRq1zvu09Ubq1mFlMKZ8apbzM+/YjH22jgE3QKM2gfxU
AKYvq6MR8+lgecMtyIUT07qvDWCR4/lqXmVwNpExHRMKQ2Iv3XZPhHR+lMtN64xc0KvmFHRHCS/g
gaBq/d3cdVnwRQQ0ZtfkKquO/u5OYXNoA8WDbEP7KshOG2QLMYZ1s8Otpex5Y8mRYbBsGnpH/7sM
iZSLz28uvsT++Uqe6PkFWce+9eAww71U5sQK1KMJJXiitPHbiceNUf7Wbi7A2c4OnDMItQpnk2y5
Vn5BFali8AZ2Bpa9MH1+tNukkY4vRb+Ks1PKX1ntU6pcndMAT5EEpVKLxJB8/KfKu20zoyXv9av9
srl7u0p3joDAcqhy1aL+PQUyPvSfLe1QraUSRChjYr/ND3vGDFO8BcfMLG1z545svLBJqD0tvx2T
ZovKE5sAoFFwVc5pAQmSdy7tangJo1th5aH9sDdNCuUWNp1sc/ZHQb9Rgp1g+tD6WCAcU5BvABYk
86XtYH2pQwL+iojL1GDaW+5mNVenCHhXju1Rt6tRCAQnen6DID2KzHIcO+MBSew6ZlDZtfehc8jI
f9PxUi2P7EMmY6aee9DoNsCegKyuwckLx/g/qwIGfDLUfHzPvFihEalKYQKnTZ8uckddMQoHurke
ipAQEspiNrVZ++hm4x8cQOX6fEGEB87eGP6sNQ/v5tJaJEI2Tg1LP4zQxsKR4yla209pk7aybRW7
mM8MOFY9r4NiyoWOmoopE0S6fQ0qryT9DT1gfyaVkvk1oLL3JF/Y2IHA8wjV1SB4qAEFweaIUks2
BHl+xX9ToYnxcQZlHwZO3Ts9QSuar6HhPDS2Tod4rtpplatvtP3pkGJB84h5o6pCPhMaIBviSJyZ
uNMeOCB8BNpjkHGhns+RKP8B/puF/UQ9PEbDaaV34uRSXVcG4e66R2gOY6pL1B5xpg+qv/W5rSUt
XWeqDuIo8mhAefzUvdkRMkcC0neBr2b5bFFMxGW2A0Br7Kxhg3hPVkbAwAptSLHaYWwod15PhVQV
SWOSDsKo9hpMVZtfzgsWYgQxRQKMUFbyCF4laAdcHRaneIQIgoVLtEYLm0YORCCtCZFQKutB34vv
QrFLNGGuZC2bqomXZ6k5CTsAviniIJoLzxGqFZnImt/IGMhS19DrfLhxvnnDiB9m3TMg9zUKAsaz
7v0T0lB9NuMYhhs374XwkedBHRjOe+KmqBwL4MMtkkczy18X/rsqLUHNAsUGvH/IhozkYNXj6YcC
HVQxaZIE1gp3L14bEShyJgqr6CWl2BlTFe/fr98OR0e6CwdG3UR/wSGGGKgYrExCC1ybmoebpd/2
C5eDfdwmoLivRMpPscIxDzIXQKX22IOt198eQqzAaU3DyYSVJFSFuXDUwA/zYEYprtv5f2Rv5DrU
FHHOL0F02o9YQ7qmkKw8YoYF0uT7GkeIe5SDgKvmRtK88ryQKAfi2baIVxzddZVlC7w7NYYLQPqn
riHmg5TpCYilSPnQphpI5rxEsWhJ2XOK/EqWHOjJyIfzV47N54NDnM6Eg6seFi5lqibAhqqrWGXn
E83V+WsB75I+oUi5uwE8CZhTMHu+f/E+BPHQsFBzeAQgAd6n3oFY+m5pFKle9LoFp6OSSl5x2l9z
2HsCkZ/2nTqB0X45ZpXKNF4oSIHM/bFDMK0LUvLINtcsKRoty+h3b6km+hopAbdlRJD2LGN4EaL6
XYLwDXoRNk6gsdONlOdhH35Dd1OIpH81OHUkfhHxJ/uoDsovRwDUcgeQjHulwKIa09Uu0y6ryBcy
EJACiJLjlbcdO9RMiDBhm8kdkrbGcnNR7kEjcyHzXK8uCnB7BiWnk7NX8qO4WEvHvGVklb5wkqsB
aWyVdgKZ1Kix3g0cUOHuwDGmOxltPVf4plei55erNAKsj6gXbBE6N6BgajoGPtZ/jCusLX6Tr1ip
c6WR5HlqxYiKV6GWjBQmUAS7K674AdNeCdhnZ0wD1gVXJYf7/8G/PCIGY3qhuD0Fe0XT7n+f+utN
gbyh37bRDF4myyuGTUd1zDdarXBnjDyd/Asv7EKdjiBqB59E4yixE7HDCn0/UNzPc0PczE050j62
TzKe0EVwRnHokOKPimYjBH+OF7KyBKU8Yt1fn7qyjDJttGQm4qwymmVgbLmn2tlGaN3/UNulOR4p
3dbUyxKCK/qhQQd0QD/S7D9AV47iMFcLLtfxSnVxXEuOK9+/2vd/xwr+bdsxymnpJKf2vO/33rBH
HMtg+u8FruP0z0Rg1U7lTa/Cf190c8pvFU/s2Lnz3oQFtG+GkrYWc5Iud58l2GlZnwWbcPRTVEIJ
45ekw+EtpivUs3z8g9YwaSDBBxoKjq8bRnb3Wfp6XIVXndEhk7YVWdpbF0QaWcjSMICN3BnV3P96
OEeHn/APQ2cOcPGQjBKiMaqx9aUTJR//Kdh5vjdLTiZfU6En4bVJecdprybTSU9HzHs2bweHfem+
aPhFqdBlkyFvZS/g/ZRxio6CICD6SvoSWmqH8OSlJ7rUf9yz4acipyhLFpUzIQNLGH7E9bB0kt9P
MHk3PIj6rCDu4J2aY0UeW9mbx2vtZHX6nuCYDBZtyqwRzgOA1Xm26Hp54SvcN6jOlEwtoTIpX7w2
utk2CjNQYDFXRUPweC/GMIlJk9HD9B/n+1cjq1hBfqgCon38tMG4mVt8nYTlk0D3oXPMKEKrPitE
+WPr0NArepfM4l/BWGsg2ULymoZE3FXJkf4tYxLHFJ9MDpiu9CkPDY0vKJURxLCcNBiyPePsB/Yy
EK5/J9JHxP78iZGnSjPcNYnuA0JhAd2i+an0SzDpjuSW4dNpqW64sDGVwDChFl8N00YmTMBU44ND
elqKbaqkv21l5nFEKEQAGwvkFSsPBk9GlqjBj72eqM3y87fUquKn953TdfTRDkU6yQ3T6F4hV5Ic
mXNFW3qDner4WQlvG1XQol4SMyU9HjLtptkWjXjRjVjEHJjm6EGsIXsLrKUMer2e6kzfFu0AV72O
pts+x4fGoFcLP0ioY+d+b0iT76xI7PEDk0uHb7oe/+IQeoIa4q13oErVPglmtx+URCN6TT8wfmZ+
UoxbrGet50kd5G/5J80p2cNyXfdaAXCWd9MlnNDcB2J8jpRfwRedAnYuZ5Tumc+VIp7Jr2QDziNc
VgReKnxbuQWfrEiDsKYZZmEgXybWAbEkH8e0U81aYu0GLiU4JKaJkqOagB/QJL3P4zh9zwm7z+2m
8EXOdOWwYk2Sf8x1oWQjp947xj2UeKBuHca/ziKgfJGN5XtBHvAW4O7f4BwGKz8p5DPlKwRBFq4j
JHTiU5M9pjPj7244BMrdydU+k3DOvYr/VdOxfKeTpVuDL9nxvJ39h8Am6xkdtCU5WVIV/ZaFk36g
J5IKmId5lV1QdSKqbUjwweB9YpFc8Prh0/7mAvlwPYXbHo5OqoBzJqaD83lyplZWKvgIxFovImYF
jCSN6YmlvnliskOILv53yT0n3Nizi1DSfEu+Vhfo39nkSHRwiID6mh8f7jqQAFvY1MpFPAVyrISL
W22UrhTUzMj0N9KI7mpqtfHTMMbeHLRQ1wTJMUw00rguaIMr790u4j2ZUdAusV+XzMDR87bQXo8F
AxwMqIyez+MV4FrrrSeL43kOZTVUy3wZWliOSKz4DuPuXP7xeId/Ry1Etwo19QjbuzQo+hGqRiqY
h4sG3K8lrS/ZiU3pNkphXpJebTiLuSVKq/WTy+MayFTySj2tcfBnGx6CieUM8SA+6TAFWVXQuK3Y
7NhlUPLFcXmM7I5veTCjsPCgyuSK3pqPXvx5P46Fy35SCkTsrb4lielyDWjWnQ42TggolpxhHijy
OTdeibPSg9uLlU4SB2ATPF94VGZUyd6bdxFmL2ZNhz20gmCEWcEWWvxf8QPQ91jGQyoZQtPq3DfV
Kz3VnpYjGVGvhfGBll2cH9TRREsNzseGulu30uWy6IQereWKFICA7A2l8Oir3CSAQQrJouV+vm32
ZV9jDbfHW6C3xaGhue1Rn2I7dBUzG0wq6UjCBpSUQAiYOeI0sCcoYO03YjxjJwrauPou7fVTyhKi
htefrB0vCootq51I1EfItbbcczWD5cw2YQs+p9QyEVca6xoe3CKyH/2yrSh5w75txCm8ng0CI00k
RVrB23/Fxa2AGBgsbZC+vu+naKTrD9zlloddNvElWpcBvo+6FUSpmiynMNuoQswKsnuC0ajVQ0tA
EV5laKPWzDddWuqb9JPKuN6BsJu5pih4J/wHYdSgknGxtdxAbzKSJ7SwEDtgrndtw8HMb9pcCuow
7DerT6dQGHOGbho7IMNn3nQQ1kN4RTzVJ4aw5nESaxEP4BofHT8lAvaI/+JS4Sj6UxWe4CP+9ovy
lJd/1nts+v7Aj7Atw8ZpZBZ1OrXn+AtyISGvhBV2f18pwIQLj0MA+3aaupZ3TMQUGzTqNWyEpoVE
415mDle7IRTjRrSulnJnM/XLnkriuV6jNlQ9DlW+gYswuSUop9K2sZEbblhg2P4JtLIMQbAD19kc
kPfOm6jnNih0qSxdqJnsgu0hBox93sTiWhYJpusi8Fssofce9FHTf8XVmo0aiYrT99e2VyxRb/BL
4QHXzHb8kpSdqnh/svI+QQO/5IFpRS+ZhnKcEGk8WRjswGlA2U1DRc/SvIV8BCVi6gwXsjP9fHRa
fsV7ZsMZBLFPLuOC8Pjb9hyQQGt/l7ukBpSLTeA9qogsffFk1ZKq4NCMZEm1Z4wZiBiFGFb2ytL4
8cTLy1dcyLyIaG2GQ5YcXa9JOMzJANGim4v3fuGO60AJC9L3Z3mEoUiXcbtK2DA6nG/2tS4eYlID
jJRzxgdThiWjlQ3zkFbL9gDhV9dzuotOjBFjJqWf3kSj3z3LUn6R1RMhR/UfrvwGVGpEY+XpZXv3
4QjBXUxWiWcYlV0mcgPa/tJPmnFQansHqXq/SJ3IUYHKvbLdoU3/LgzHTkHSdRMQC7DWIap7esU7
kXwE5t8t8eliAQWl4+5I/qsz+9bhKg+4moLJJl+NzTCXp/Kpfq2END/ZuUvd2ONX9vFvP+RBEuQf
qE4rv4RnXUJIY4s7hywlyXdg1ovZyKXtnNsH1m5vstfcMcKgILKNcypeqsE5fMleGB7sPbXrKFLo
hYkDGVEnKJZ2Qqg2i97xGdFG3yi9EA+qAYzm3SwcEd08lOQVxgOh6XTkctIDW9WHyCSgX1RYg6q7
laMq40Tz/ic7ksFAnTp/6Vx7Rh8wLfG2Mzh1IZtEvgEUqkNkXVUmAE5DXMAQnOsEQEnwX9/e8Df/
a0+SudDJVXh5XtJuBHvCA/6iQWZ4LnW6Lu9agV51rxSpqBcnz0mrkPSRqsr4MqJxL0PHE7JuUqEL
K6Y9ug7CxOiU8CPO9EYxAF/cB3kgx84MxcgARDdne7WYKGlU59tggb+ChdXVmINFS7/C8zIqX/zY
ik9Xo2eKweyGF1iI+2/vx0lmpb+YZw7MwsINYcUGspnVYqVfcQoOS1AKLRxFJds5xsoFluTc69rr
opuRa4ZeuG6Ig/FlLyTUr/IDrD58DP+N++X70FTsAScfhX2QjcXvceX2mltTeY00CeGw92dgzmfM
aM+LV/0PFD6p8zEGjDvGVefzvcxK8FA4IA97V7Z2qU/kjjR1ZinqD89PzGop2I4h4gVSglxk93bd
9qPzVPth8wIEpI2oG8RSpE1boKoZs3U2YQNuooVhiWopd6SeXbdK9k0hG+xDwA/cWrxql1ypi7Ff
ntPt5a0RKxzPTIFWteL+qGAe/UudaZfcarB0EjOqNeJ9Z7+2OA5m4CrsfZ3xPkgSQ05myCxtkzmi
3ya0oLWNr5L3YIga5BvVNbwML7Shpyr9gR2DkPlxI824GXGmAG5BFcPtsxROq+YOC4CoC01BkgIM
LC7XRXR4eXd3VWAro2VQ1EBR8lG5oSD1FcaNasz1WhhiD5jjkWPMRr3f5eNsWCnAHAnvicu+p/xV
QpjDj/6HS5ISm/msCtJSXFIzcj1Pa8NnhHksasStlc9LnDEUPUCEQUVkkieP2rFmJMKSYfMCQ17M
1qbt0KMWIFeunC4E2jnFyetnuVzlSdEL195CaswkuD0X5yrGd7tAiISxQFYTgKAvLKqOWMAufmiz
llRnMHDo3QrDvikI3wLh1kp51yMDeH7uQjAJWPL5OJZ0oVwBt91vSoIDk5Ztsv9pYVQ025jcQHZ7
chE893m9GE4bAXAfm8Vf49WJfzOL4Hi3OK4PuqLp+sBV1fFeVvLnGe2tgiY9xtetgh226j6ToPPg
fmL0Ch1kvEQlkO36Ijs6TDcEwgjEHI4dGq0kZkxKHpiBPjhntALOilCc5Cv6Zbh2IV5QcGGykye6
yeorEmE9mFPRoc88Fa/xVwtDOrQEa6AB89Ah9jV73+Sal1GskzquB75cg3QNKqFmJ3vWNOfwqCEd
ezj00NW8g0QVx2SLlwH5IKvqFWG0vn8YHMAnRHo20/NAyUZtOddDP2r+Nuvvngvk4DI9+rWmLk1u
eiVm5Y2tVNz+B/15bUDyPZ7YylDIN3YZXvY0Pri+MSW8MDNF0WfRkm/AmaJqZ0YshxCW/7qliN0Y
VwmMNpxfFfFFJsdaJucha1qfLE2ebbqtm6JSLX1ahN66rTLKzuG8o/3BrlHvobAKIFA1VT3Lc910
QdiIo6ELOaIr99LYvtJI7mNZ7KZIw0D1euQCGmnYMO+rjUnQkZkTeQNTl8No6JdmqQeM3Z3AQqur
pnpZd6v9z05QaMEjoN3YBvk5g59QU/gOHnVMAHXQ2z22KiptCTBpwC32P4eQnHvKemVdY3JaS+dM
FKGhSMQgfKPWQ8olTPQERGAKrv2t0rJlALoFi+Li23FOb1XcwumtDj8SVxcuZL1O4MjntXANoTCH
WiTTO1c7pPEzmPTal1EmYsNZeyiw/R8fD2EN3B39hNzqUGVosL77FXhuf4FBG1l4hI60fMY5jDLH
i/vYUMD4QXXo8gFk5QoAGyb65SvIzfdzAg6tn9vBJWWvlP3CwiDhUTl4zfZs6xlfnJVeyVsJ8Zz/
HwP8pPYycXSXFPRJFt0AseQnyL0W9sA6zQ71MnLtcaDytVwty3ZjrBtEGVuELzNMCeu9mhXHBRTQ
VQxtlYf8BJ9TZqkQLjgb8N0AejFUo+pikKndrbVaWy8lHdcfzRXlsqEtLydVvvJZKVXm41BSGEh5
++379Pe+dIEFx6XOdEIEfvY8mZnE/vjurg1GcSJ9a3g8F6Jb27khcw/l+Zu/l2rLYUFubTnylQXb
KAwPrO56itLHFi81qAfC8mgaKS8K5q/OLFSJPQK20WuBEdpZnjnSt/I74w3414/dfZi9Lz4Lpx28
VFekvYPA1lYh7wjxzM8Trto59ySoc0ZBP0ooGe/PXhgraukewH39KrJ09u0ylCjb4m/ZSdtNpU9W
hue3xwzNhjK6LoHZYdQph6l04l8/6ugjSOPzVFOVzliMYh6qGvOD+5EmLnhud+BJl23QavZVumfn
VvpwvpVQLUcP9w6VNLm0QmbfKiYJdFXtnKxDV4UScsGD/WoJgqMebJYIbkeVQqKzpA4/BOqzPxWi
LFSpE95BfGtiUcPRoi6l1j04rVZ7aeq28uKyud70QS7dCeIZLk6Za1e630OHI12pr6nfNo1maOcb
beIJFZyitWDvxs9N1r53yxkgAYQdv15qQ4ZiYHH5L4xSZQXbZ8Ub/3FnIEtZVqnJJrz0zh0ANjYs
Cd2ngFNDjtE/Xd1xw8JtRRWFLAPTRopDZZfnlgFnC3IIrr8M00r5mNhrqHKhwDWn0dSlkWHt/Jy3
giZGuqBTfEg4wBr3/xbkGXTYcaqsWIalMucJFz4jNNcrb3iTFpLRNyGkZ1QBRMAkH3qoXNkrz+CV
DWDJcbFHLhRjAIN6JnlC0fJ6VKctLSGIO8jgQlU6AKBRPokqpeTBr9RHQtgXfzY8CZ6OD5WCimTv
8RFf5PCKMO+Vamo58lg60S4Uy3iNh5X13JTHCp9Kbm53QIwpzxKZxUG/nWX4hY7zwVdcd2WauXzI
B4jwLayoW0luCgnUK+m2vMDi+0voNQwf9Fd0G89mdlMEXQqP83IJxk/t0YvkZwwiXQ8M2ZnX85k+
+iLLX3w6FJAce+dGgS+Kj2z9h+J8teIHCwFUnP/xlFTXFMfexq8sytSM44WHdAMnaDHW+l9GeAQR
EimDWy7T8VsIIYHzfaTiWb9yyNygLwk5N+n/FOqX72wiQRzUTiAEQ8w2ZiQG0ijoptkyPPdFga7o
Yk4NSBNAYLo6euEFEP0l+MvkrjqNBavnmp6SqyRYYFbSTh33o98DVbjao4NwXBQXr84syn0pNT6J
9KyE14CBW39acb+gR9KplvPvkIiHgFQVlzQn1YsbqwWR9mfd9Hf3rZ0sPRAffLnKoEJiJ3nczBG9
z3BhkSnoHDWVYNYm6k/w+7IfNR72lylP8cDk36MOeWwPTBWc1RTVRbhW9GVdtdxLXWIhSPS8O9iw
N49pME6jSnfpi0X2MVHzZHmeipS/1h+xTJfOiFqcOoRNZ1SsOv73gyLSL09gR2uOLY1Itf+Xu+wj
wD+Lr5NN/7BIoOz5sVpR6IrR0peTDf6M6AJLmMQw9yitCgkHOKNCfqL9tfcZf7gC395bC+ItDeyO
KzhXXrTwa7PzQi8GpJSebzbLAeE8fHbFNL0VTPN2GesWYMY94H70UL3u4bevgjNkpI+3JrqfKHde
Z2CkJG+NwZb0VtkRxTeOgTfIUsx0nHejPu/wiljWgDktf0qwMyqJZnVKchW10flFp6Zz+URLb/1V
zMHOh9OqFozSozJzm690zgKr1ijPpaXaTHj/XMu2fZuydn21p2izIovJlGE8y10/7Tm+RKYWADUT
oaR/pWpJXCeNTe1tb5d1hBW11e1e8ckqP+0HcoN+rdXS9b/SZpOfRXHs8MLjiBGoSz7VubZFmKPx
dq32qNHtR4wb3T1KWvGmcHNWjEaPZe55RSXeE8r3MBoql0dVYsvnYHUNZrBuvr0kikJJ7sGz0TN0
44qfjTNeDhI4G0S0Wm5jpp/1ikwnuzFydvyQcKgb2QiSVMVmQQPWGoMpcM/85d6H8n9Oluf4lp0x
ZA0Eg4YRzFe1DNCYALVD1ytLc1kwTfpVXEh3oeKBaN0xD6dpHrdF6BVaJulEHd/AJpmB6FU3H7fI
8mgp0PQ4aZJ666ctsSo/zpxd8vfs6FP50KzCp9sBKdkzPz00chBsTc6pE6TMMbN5UaqXblG0FwdT
lq6oH73jIA4s33ISJDzlFSnaaIiGoW2Eiu3s27WAUzikbGf4sVayD0HPW2Ifiesk3TKfufM5vnvs
S5uef9vs7gzZ2+kvUfnZyejTFA5Y4pxsbtETpjrdoxrEn/yEudOwdiDnU+hQfgNZS5RiqmRZUInt
kX8jYQA7JvGC/3vehGD1ZDAZujbQjSvF6Oy+Iefcb0+Yjd/4r/rfTBEqsLWVZFUGVz1AQq/Y266z
vF/P0BBgOur8chhoosXIfKYcZegyyJfU1PFNq8HOYd40/bLJauD/j8+KXbo57n5mcvCjAdWKPxeE
pnDpXj8uAnjST/08ThkSbzsoZvbySOgxMXOivywBCq0H3ptgJpsf0U+zmWlN+3z9q3WOx/zdxG9U
hhfjzNM+0H/OV0JqJpBoL1FzR8LztoHo5gTc7HP+dlVhFH4sVaOReBXgVklcBcRSrzDJZB8kJKVK
iA+qYYgKpSNpiSbrJ5BaxPmMWcyle/kQ6YEHeOxw4LM+Qi88woGmtGdxLH5Nr33CI9C3ouDjW95w
6Q/mLahRTjoK5vqMrhWHPpt28pVqU41/Fp2sC0uQqF6qKh7OdURB/St/31b9MgWP48VdlRDugjzY
P2xCLZdCThe08yaceR6+Da69RVVhNDjDkFMmooOJsHYEHvukCrSHZrVY8iu1kA2nAqbFDTsFJEfs
IRvLOX+IzCBxJci19Icne9WJ9Gbz7lr88rxJ2/4eNcRethk/4PWdpxazdcos53MPYOfjzxJGWY/s
Y66dVa39pIPHBBRT/MXNQxcm2SPsmD+2KkwWojdjaYiytDwOPBCOXCkVoRHUVMdsu7JELAr5V9dx
ZTrFEpXj5ozu+NMjJlTmEX77FJDSCwKabzFlyMru+uTbsaehR6RSA6oV3LnY5r/z8iXFWAUXD6VN
42ahYefkTscjzDp94Vejl3osoY6TrISi/dWyshz5SXrW2IxH49+dCorkk6nJaSSM4Nq8l/JKk6cn
hho3bAKdvy5MXHd9ngwmcJWEPkLDNFDu3MufDMkheBrm1Da2UFEqPyLApLx6/rase/AdJFMA4Vb3
IKRAMDjgvYjhXhi2z4clE1I8NiyCyWGneJpRiIAZP0Dnqfo0r6nqYfT/OXZt3R7PdVYCXlENcKGR
dhVfsgIWBlYlOCSHsZOcg7zSaH3ylG4hssn6Jl6oH3E8Vor/mWvZnxKxWQgY5lGUa9ituRc4Jg+o
FMbf9uPNbOpW2phco38pZbaFWTUCOXDMkL62HNJi775GY8+QIpahFpDFbBkvKrjvGRTcCFZmNgAo
gGxOrUqJ6ali5EwS1+cirJjfKUnE8yiWDtVElxS5sG3qekpgJPV+JVRLVfdgmni115EgjHBRZql9
UX/Yv8A8Ig1GYNjGzb81WWL0tyAUxAYfmtFMJfhkd9+17tKWcnppzmKMye7nshFTr/6f3aqV3Nz8
tjSXj8+nxmj4dmnyPBoj+BMlwO7AVZQwTLCusRZmYoVNryouQxhvAbQK8nRozbJhKT4tFUQfAYC3
5vIsWPBw4HCgjmXj45LC00g+nIpY1/blnLg27+hu28X3ZiN3j1bJhXbs3U4nnmJiNTRtG8Qtnnmo
uM/uroNGi9ip+//nLo1V1MgGT0q00XUnLDYVvZEJF1XntOZ2mMHz1ilm54qjhAVIPt5El1Rflbzn
zRF06LD0ETz9uwQxtPQnJmEjNrWC19wZA1BULaawjWGk+PAPkw/Tn+0vYD+XLmw503U+LXEjm0cE
dyU3VWyIwR84dYT05+HrM4cx7BlKZEWAKpHEjzdyDK4FrF4kSNCK92oKaP9wJze3YtS16bAayXVF
4ETZgfI9kKe2UTsqXd4S84/jgKaff0XYMm6z2DKURiIB/NPwMeMIzXMK7xHgwYBRkNaQOuSNkBbe
aVh0H10py6/86K2eZy/U989eOir94uxUomZRLBG/7MzVuGbZxvkKJ38Jv2R1+ItlomRCLiUv6BT5
+jsI/isKFNS/PKhFt6WwoB8NlwR0XF/OurWeGsAkbvYEwZmsp8KqWtoByJlkGckJzjqV11qKjy3k
bOk+pZ7NgeE/D61IACfRJ/I6Pv1lHjoK7YsQWWSKrosQ1HDuMI+mFT30P2skXC40q7+sBa1hmDBW
nifKa5ruuYUVUqxVyNX/M8ioq1T2NBNmVY+43Su1DAdtk+0q+K80h6YtBfLTOHY9n/WdlysxhLnt
cWrhbhEWyN6ETvDMgF1FL4iJAV9cuwB/aVQ7bgPhyrF5JpDZZzwYRm8/8ExXUw03ihiDBqU2xgCy
D7avA0bHNh4VRKj/U2CXGT+EyoREXUh2o92RAVXQzBYgmEHTJoRDYGMJF6j3LnvtbvHR3o24p3Ow
OWrqtp2DwxqcWjGK/3JAS3aWwaNjm1h8Y+0tMEVoUxI/6WepFry3a9LO9Twr+8rQLWFic3gieEK3
sGfGVyP+wQVwbTZFmhRws58fpvGYjkhw2jb81VQSJ9au0hMgQR8tODJu+rMLvCFjBYJuOAFU6WLY
dqRvZK4Amlh3jVG3B3n1vWgZTsSEY2/f+btDWnI/0z+liB+6rZNK6llsZH6abwpNlJOIw63AY36j
bI6RPzqOnIjMZZ2UjePLVhmdXm2ZX8W/ZkdAWV2CI+NUZ3gZqLPn+q9IIk+XQ4jETAhfq0M8jVo8
ZMlecUlgYBJ6pjAfJpaiHr3c8MhPM/DY/JTsHofy3yJa+VriBgov2bf1TQJd2ZbP9qL8VlBQnwtV
SLz/oT5Orq1GuNyGWNqvbYbVerOHgLl6fulkMplMmGjjpVXxwkJH2L4UEhRry3tHKYAVlQJESBek
MxK5rMp3warminCKgPqoyg4fhWcUFmzlsc1ZSYS3D6mfhgVMl9wWmE5pbRSxoW2VpiFuqtxbKBir
12eE73rUVdPjOhCtx/B8f7JkbWSkTMwSHipnEIG37W8mhdEnpLbZBg96Eglac5O1PUmNTEcaIpS4
tedk4Wy5yOUGXCQr2zg7geTx4NFoSkbbNQX7oKS2zbQMacAbajSAKQaphxxFw05lgSiVLqyTFJNP
aptnTsXtpRtCGfFNxAQ+yK4hnV8/2Kxt+k90nFn0ZzfZQsXgevHMjKbAcSppjqjlYEn8GWCUQ+F1
ttzw/3NVgZ+IYTWQIqutt+Po04nywbA0nytJQbGXiNF6ObxYOK5gfHUT6tbEG+vXcRZXUT6zeZgY
ZP1Cxs+dWFloJJ7LQc9ebr8SXahUrMtvL7ydgdfjDCGWD51qjterVy5oXtw0HcEomZxTClOILNsF
qXeKsiP4xwyPechaB+ybOXZwrtvvJwvrAQOYROh0BJAxLaXdCr0eylsU5j6w+XRvbUNFyuCV6K1q
YLytHKzY4h5/oNrPIJJPaluKYP/UVh6rly+osF31YSpyc3gPwIOgReJCObE3Cdvu93SLOMy5TAqB
1bmb7osF+jXKZVd8Ok/RwDmd1eIgOwBl0u+4c8d8FDRUL/hoE6Of3dW79AtEPB+Y7h19jJXUfJH9
KtgwcT9L/2+utIOk6mJV8BclOz76qNl00HqoZWz3QiypBCE5GmuYvuDxUQbL5DRrZpXasYbDI7/9
9vnGUvtCPdzfBvVlfkK3YPLku9Da4fmVEbNvM4M4JDpxsGtN6EmIHCAGKwuoNYqkCAbrs/pvCmpe
ctW6xo4ySWCPYKwLRi+W1DH7rp86g478YJCdWxF9ZT0eLa8Zr5GVni4ZGyESvAdUWUCnE6BrX1yT
TQR7am94aLVrUC7RRJJVxg+X+iQ0KgbZCFz72YNtyZnxYPHgnXEDaYhnn+4w+eSsp07oTvMDYu0n
DCU/WGF1VCeLjSUSjcjhdLjjgDkD/iO4G7Xe3CFVioVwL0eDDW8bKQiMEeSNpR/7c20dTR2qWDOL
04vnZQbiTENcZB6sCwXkB/cF384bFYoU6vdmvsCsyMLVvL91YrDEJHkGct8sMKZ3Of97bk+XXOR6
o2j5nlOkNjfMB1r4U0GnH1QIpKm8zYkbBwhltsHU5166wTSnAztRueKbqG921JjE9TDOJpy0go4M
dXST/m9zK110SOKNLzQA4ztCprV6ETTtiYYr9zBrp+teuc8CdM9ylVlnBVI28bk6bMEHXV4ayNvO
phE0C5kZMKHlG3e22oazeIaE7VeHXIkL5pQ9isvkkPH8dZsEyrvSkkK+6xxyqKXFsfBTBAGNV+4P
H8N44HB9+lRuKsHktmxBQ9sOJ384Vo5PLdM/dLWrL6hIrBxPI7p/nsYRxlQnCdOJ8hnbWCmA4u3I
2xQrHASciFt1XKdxPo1NtJH0ZCBCdfAk927k5b1yFyucgPSJdr54Qk4JdkampI+obDINALsJoo04
wlpxR35cKOSRnIJQ0uB0hjd323GFgDjj8NrTVULVKWSPbJgWe3K9YA9ySwL7FIDG0EiEMgo1VvZx
3BW/xHcj466+XkGPhZLlarpHYH3f7jc5dwIXelAZwVBUJj59+B3IrSMFNxGVXZM+O9kTeByLkmn4
/JiIX3LYXRkugTWvWp7sO7EDeCHvzeLOlYSyOhc/ld6ehUlKbZ84Hsp6MLUf1uHwDFQ14SRzJUDf
3XNSqqP/LEsXkl3kFlCQYS/idRJqKRW2gcbqaBgaIxLeplxVnPzDNjVv3ZC8jK2Yvx5kKp4cFBuG
uhRscAurPxNNf5uFXQCc5iVgPfJqRuUyyH+IkoKnHc+brcYayH1lIaTM/B+4x4KEXpC0P/a0cx8d
gcl+1t0nGqnTAlYreCQKbCZC2GxoU9GunM3joLU0Vm85T3odGj0cUwyvHO5sKH2t8cFLjtvq4e4H
47x5eEmHULYvlouy/tgZ/vNtaRFtV2aMysbNR9e3SN6EAo9QFyI/t1ssAZo2OeSP/c/Xhyji8Q9p
aZX5ODrDABHzZUiVaBCnFcLLePeI6YYJ8pmfPQe3QtLLRiZ6dEVVWP+XvCWOb+xZa31ux461qwbk
vkf6qe62N+Ib4X+Ph6RhhNhwaAfKBLofX1uXRXZQoBO4YhIE8hdIdF/xNl2RWe1+l2AebF9FT1F/
pyImhi/MfBAA2oT/B1hU0hnsjZ8kA+l/hFw3io8UU3gomyeeU1tAddKrKfdTEbCicU9AqRQIhkAb
NXPTMwSNfqJBxLCpcvgfUaOMaPwggbTeApmMLD+XeTK4eoWDkNdOfi6fzOZ2AnDf+LaFh/bCvpKY
ZKXBz+LQUQo80AiZVcvJEKbX0rQnfJTKot/GdXG2P2M/81jJ3b/iHR6cm33TmCYv4eSgW/p3rDs9
33/NxUQGXYiCAxBTiTWC+jtuMOul3zDCx49NEHBmlydy7tw7/huGAOWkDttGJ3RfGodkjiPQOJ65
YZS4hT9fP3eUcuH2ShUvI4SC6CUamUw1AvXOfbJ1392Bcke0FVxzvK0jz1m3LWAlCTx5XrD8bsbF
aEBj/PSLfRvF2r3rfXnrX3oYHS13y2OUxsd23xU4nADZ2m2cNuGxaN4mTvkNEplPxVvXZGy9sX25
xhGD1GqICBC5yx/pYM7/mKb7kqxKXmeZeNEb+UoMYlB4NnVO4mHMM/MloqCA2NFW5fbVHbBJpPkB
MxypUwx1hYqp7PGdnrePW7cdhDTz4uXFVp64dOBj9aRkvsV+abHpYzh2h9OE8uVEFq2uk0A4cqPT
FTerXPmxKoYk2RUDiQNmmXFGdgFclAQ1Xfsh95u4dE6s/u+xqba3kJ0G5CUnxVxRv7szeAILj/Rg
wzGb9sIxuvzASQT8I55zqgXi0mHvjxkf43xQWwB5i93Kp8Qp6BRjHzRxA02yKd9TO8+kghBqCGf1
THrnEF2puQcS3oKZXeDCqSNWXQbtS6W4Jo4YT71IE3szXLnEb9zNkocUgHr8uXvbixUfXoO75GQe
VeRhdPOmqLxn9ZHXsa11n7oUajaTrq4kAR35YxEGzo91vlrCkg2moIQTui8OhtQ+j6eOLe4iHHD2
5PWA9crSDjxgdcM2RliQ431pPxTJ+4fJOkpzsJqq8NeYAMYkPJdsQggtgXKx/2YQcLTnhWz/Qjqu
Q17Tlg5jg7qxtqMi1UpuEk6OYE66c1NyjnWlGF2roF3NlsihdHdW9k/Ekz99tUQE2dcufxsJwu8V
lDTHpvrwAMykgikPJ0L9BLuVSF8Lk0M75TtLoCN570ychkv9hmQPHc8pnwamxoqOCSqnVqwWhytE
AMSduzxxZZMqDARrSQgVf9zc4ZeRf+IEJXJ0NFASTgr9a48keki9LA+9QSaa/RT07N4027ihgfZo
7h7I0BCv0XktGl7x1NATsTK8FzZCyd8ZnJngwR861dDE5ytgHvxpIzucPpjrXUSc3G9lg7liCzQI
oaLLnnt+qyZMK0tdbzdvw2rG4UfUbWnrTZu2J1LPh73CSwPzfuwszuNbtkMc0sNK5plMXarABqPT
HLx/DH12pHCj+XS5B5FUC1O6IhLwkse6hKnF2v37U+1iZFF6z2TLnBykHCiuaVD2JUZbDwJMmE0l
+HPKbOdf0mn++X/IsV5dCczhp6ZumG5QOR8SuFeXq0oyINhtZ+hjSMqCZg9Ws859FVdjyf2uLyiH
D96bH/caP4t/TAjvQEGxRIBDSDZ7/l0D97ml5rxvKFr1CZc004Ue1WbteWFCDhn6Z6nA7NC3v4OA
/vrpWQrANP1dkjVbhT55tEeW1CmpUtk/8t988TYBxsMCrG1JvrZEjq1le/QRGYx9JfArVmMIgkoi
4rHpaHNoyLVZBZxYhpJpdiW/MBcSIRilAbdlv9WQPrL56N2PrxzISiVsWBSFvrQPaCXP6X0M9CKx
JnfmFqtuUTCc2rfQxMclFoL+a1wTraleVRydr0P2uB/nlw+tKxIKwMfX5lYnuBpFWdCfJrfGnDxG
wjYCA2b6p4fwELS1NVSlSUADYK3Wwi8wnzemrE3cSIiJZ+BIemozG+mBgmy7qbX6d+pWWaOITQPv
9uWSP8o5NGKs4CdzzAucsGkwVeGPQc/ilKnWK7mpDM4gxzDi5nf+7POeDutAHNsCjLj8Q9HjZeld
UOdPBUXG7EXz+N44SCZ/yQTdEKJYUftFPBhKYBB1p4pnf35izyExEAwLBGZZoTGW4FQvLXETdPiV
8ZVW6AbsjtlkgpsuROcirNXs5MU1Ox8YTbcWj1+6FnvlxShIyY+W4WgkH7+kA9eVEwgt+zA2e7VF
WzFQbOfxFCXZUVfLMGP5TJr6YIyjMPrkhBviok0WKTL+DkIGd5sl5fMmBPZQYgb2cvB7zecZVYMg
qpTNX712bIQV3IXo/+S3JZZ7OVL8l4KMcjEc1T/naiUDX30zfcpQCsXEr9aMbdEq+uGpdxISA/Zd
qgfkIINkKLi3BMgi5dcGMgPWDxA+nAQAMjyq050JygAdcrw4wQVtaZEh6ykSPBoeESnqc9ND034i
uN/rW0Uot46HUyphElzdnBMyCynLXR3lubbDISGZsZU2VpQe78sM9kSe+UgaJj7cn7XegaygTwHc
HWLOU2JK1yIBPXZxzJ9cWaZFp+WbwimuTBY8SW2MgOjXJRVOjlREtpq+bEIKSBt/fdXQhPLTLT0h
+fhcz5EcMkBuwnB3kIjDVtpgZa8ENdypAAMfwI4JhmU3MJWByhoeua9hBVnyGSOSXYm3PQrzYWxd
PWUJPtZyuoy09MXrf5LYtUqlClACJKi4V/vtkvdB2R8nWywJUiisASA1kF88jCVgtTGPjo427l/z
2WdY11OtjhUjK39gKqpH3+w2TPfNT6PGMDLiGUWh/AJ+zM7R8s0AUnq0kGbrAw/AkBU/GLWX+cdT
jo5bYZxmOUq3/BV2pyqvvbJyW5GoV2ieh+gyMhc65uvc7eWg9S2YvLCaFY8SNUxKtX+IsH433vbf
D1GqtOQDe+YFxGz7azaXZVnzhaZ0Bk1FJDx93kuGF9PPU4siNoynBjWRAntPa/PeoZPjMhR80Jjx
cybXgYsW7VuDmeffjNq/BDkbBXsBbVoaMpF/KCn7Iekmbnd7sgrl5MkvLIjtxdAWu70h5PUxCMel
MPRwBoPKqjtfQBqxwgpVUIn4vemH8X8s7tsapk8Sm4zyEWWiJhMjfOf1G/zkvtrHh8AAZECLNTIG
ABlgn7nL2okRA2eEV13QsUNdh6WZgkfOGxeh817YQE6hl0mcoiOEIn+XPUhUT2t3sKAeErpG1ps9
jUTaGIF+WtQg4Uegjazx62qJ2rCVAm9W+pU1OzLy/YdZY94qe4g0+iCaR9AHArE78JduwgogL53q
3C4E/cMQuoNTspB2WBVN+7aE6SB59qoKVypVwD1g9nblswr+n+9Cky56RVtPweA9M08K3wcyrsUm
1pl4uuzHmsoQm7u5qinS/sFSToITDFuJr2t0tNoQ2XKHdjrVpd6rlQdT8RmNii8iK4wMZHfHJ46c
orV3lmA0Sl0bhqrFc3+GX0jo79joAiCUSURLi18CFr04cLnHZ4RZw8jcU1BvFn1Lgt5tCdyQjOSr
3fOHDtJPjl3HoGtHlvK+TtdJY76LPWFZ7tB+Mj8kdQ/zpHm9sp/XttVe7iX4mZjNXct9G3jgJ6b/
l2PbRyspFQjdewI8YvfE2OpzscqS6oKYOOao9DHFigiSP1OHqnRg0zkYmDurOcS56TW2AOYDci7v
eVWrQBVBQHipvZVrpeMxxdvpJfoZUH7REr/T6eNmEujj6yuCGYENYjnA+dxsD8LgM0D+GwAOhZiu
LF9P4VvTyiqf/dx0F8Cjgro293D4BzTuEkZNDyqFfgaOCnSLFBRbBRazPyHJ2KlxRP46mjZvNI4g
m9hlh8VnhNhywRZn8bl+LHzLLpje4Jejr31dCwyWLOTRSI2sGMklDBvaFveA6Tbe9JNoctPDAJaR
Ddkk4rCANeN8KZ5i0prmpwM8sN7ZCguMdri0dHciQdVPdSPYjeKeO4JZbkYZU2dX7smmgTsoaJNH
jRmIHajsQGYpA6adLsbgvVzB32eZL6YoHa3d6H/5mhjLt5bmthaN+VyaxHf7svxBkWBOf1EHiVru
wGABbULaL57gQfJm1G7aS6zf3NlHLOUURv4yGlqoh9huSZJRB9Gy2S3G4Svt+EKUtz6C+SCPjo4P
JnZCfEX7KopGqLW8pu90QoQHcdhz8qlC3WMdT7xOsE0r9DHOIQPuUsF4MEicej1M6XNvnbigMGLB
IL/CB3CMI0aWESM2Fqt74RfCthoi9mOceU9/F8pKTzvW1g2N2HOFHLnMfIFp7Eq2UxVMrkDXSXxV
rw4D7y+12iC1R4zmPwROv75LO+Ox1uziufFmqvfEy6IqFBrWYpQtfu1HRgiiw5JA2kJoqyEPxF9p
C/mRaWD7/IZONtqaspLhvF21ID5CiBPPincQXiHLxtFwNJaw1+EPGagdel3rXysAMMbwF5CpDVLp
IJOPfMIcDpemWZrAsHu4runK8qAptHa4U2km0zMvu57oiRJ60eVYol1YDkHkCu45G1nXLH6psrKY
VBs1C2oEJmbbDnhilHgzlcaHxrr0jxENtI2Gr1OKyXRMCQiKXqj+4eoNi8HJpTuq0w0fjJgj7eSp
egTiXx6nzywLg8MKtSJGS2hq3YVV6/OkAsdfESBsBvjglomgyYOMhwCfUBqnk6yjlAYMuWDmztkt
wVhqK9xrlfRycM64SJtjSEtesl0zo7ozllcJC2A0EOuMQtNGnPUFqBaZuxYs3+ehu1IJoULNM6Ur
HhdCu59NsuqMEz24L/8EYuR2R1p8uv5iGvcqGtcKiS79Hxxhq/5o4wtmugwFXig4xLurhMmhv6j1
kydSfhzyhhTXWSCxTgYCZHJC6kIvB46sUk0JDaoQLhS5n9SHISx14REMcvc+SZEj/nNf9O3b83yH
K+MEXOk8H9bu6PdwgsLdXJMiCRn/e5fvu/MGsgV08sLsX0AVU5zXH6IQ6Ha09dW5sVfYOXM2HP2e
3OHtjQoKo6pOgC6/ZRSZfobd6tyb5pKTF42WNTrhel/oyCzVq7Oz9YZodJ9hjblbEO2IntbOPKzn
GXd5Np1ZAP0yj30h0pfqOwY2UCnjCCkjjU2HV0fSG8fGFcR2nTf27ZHwt5GrYn25ROQOeozYEOYM
jIDKsux9OYt82XWVnzDb6YGekFZo7zFhsygmAdAek1aH51qiPDFfbSDWQCJ73YoaVDzv+Sa1cKDd
f6p3uGAEz0CtQlLr9Ngq+oUvXZqKZitTmjMkmdJ+8Du7WZM8N14a850JLKA8Ubjv1jQpRNSN1RM+
CG5hpVDX9OBZhPDAb0pFg/gf3mddo2Qa/vIKjH3+so+6/iRgqN4AH5IJwNIf9Y9HIf7bvmeH++ir
ouwZrJXh0uxeVFMD5kZ9rtFovezWLx0cpgfOMVBzddQAggZmJzWOGPVmGF5kCGqYuzv4vCmq7xIF
W4i4cfwkUoZ3AQC8lCyUZg40PcA2KPcXianfMb722q+HSraootCSNsUOpiuvzwR3c3WUy5pdz2QW
IhjcyaOrUrz2+rmlECIz7RMs0r+ylg2ZSSRQizCIO+xd32/23qHdlk8883c6i4A7XJt968ZgKBhv
YXXz1PbOfjLDJIZXuFZ9V3GdPCh49Sy+pbblZgTZdTRCjHFUhYJK+MibdFi7dbjmz20jDiWk65YN
cgLMAU4RyOu6JpmXT/0MQ6AYXfJejbADA4RX9vuoUoimcFCbeAT0Pk2Oxue9k3Ra32ZD+E+4jz8C
iF8Jv5ttBx86ItoKVKdIrwd4JTHR2SkpCoGq4ym0Ur+tyaqy0p607Yj3iu8KpMzBlpV0UaCTrxhO
BYL173FcIlIU2AnngYdCv7EFDArKk3v0M6NvHJWF7HLNyb/ds5LDzhvAyk6NhfdsrxUL8kaHLpRT
rYHfcsQdwM4GjssEmhcYWf0n1KWd6MTMJj5qVPMyW83Bk2ci35EVUmPyFJsYfsVu2qqEqB/hytDb
ar93NS3ajtHjcYQqyoZvBkNwD916cAxn6AXySRIgQx+3A9K3ig69mLwx+BQtPQWSf+6ANU5GBCvU
MXsXZ10zfBkyWwfpSNbeJSpna6dWqSZDblMOcfmCnsKHhREyWTK15OQXpQS6sC2vpnJpgze2Z3vm
vtK2yVuSeCq5ccztFQsYdfs+p0+GZ2dNgQzD0K3Qu8tztkIGVKvQ+/FQV8Pn5ff31k15BNjqJRjd
YLcbIrv9VszHe9JHVJGJECbX7AdPz24BnRvTq4+GZ5FWcifcq0JCwJ83ZbKX1u5gDabrZpqSUnMN
rjkjV5yGt/18lfJEiyvF5i6LPVJMD2ipNL7HrnF9yd5lYbx8cRdkeoBrSkX/1DKtVYTADqq2t9eK
gzmoW79OSEpIL56OA1ZbHvyMkY+wQ0D+mKoJG2VwzsrM4SQwxwxTP+zbygJ/lZggYuwQrtIxvcEG
nqjhdQycUzazNjMlfqq/ZhvgnlgBNqMVvIXwkP+qluWMxfdr9meMPMiwB9Z7TawgMLDQRcoM1ItD
r4afi9pAtpbamDo8ST18txi6qXRpeWnKcyawzf0HSHfQd+cAKENOKTDqtyBfr8ayRvro4A7VvqFj
L2U428qO9p62Y8PzwJm/b5oGS01ZxbGJMxEYvy/wb/zRQCPVyLye4u5/D+E66wDiXprFRwWNVB9S
GNUlyYcLvP44vtSe8yMI9DTy8vEXUV5JP+tb8sa6KwwMJ6AaYJHqgsLbq58flrPgcmuxclUAgt70
qmsrWg2BR9t95UbqVlJaptce9wKTX5WcDAuJlOf6kSXO0wWY1W1rkLgbqvS9x5SQbKpQzDr1FnYb
N4lqks+U18TKRkCeheWsIAvbfp99qpRuoAvKX74rw9fqUlA9pSAGnbzbjXLvxgH5WsZzvuQsmnH6
ZlrAj5CUo5inSSB6Jwct9u5vgBAmRMNPwSJLPjcU6P8UumgB3w1KdRFFmw717hSm+xvXzM/TOjZ3
pYdfzJGfn9b42+h/i3pbEQ7/a6fktAwGgdMJ4wfy4zpj9wwg5Baurf6R+KcBZl/tjRZJI2XOk31/
AfhYHhQoNbbnZOACOIYzglkHMKt24Vhyk1XxxKbFWe3GHiAxvg1DJmVd7kvUffcl/vvSxl3gTZbg
rHxHlFWI3t2wC4SiS+gwbT6J07ezOTcnVDw+YmJ18ajs9EI/iCxisVQ6cxvq5bXkM90c+VDNNCq+
kR8h/Mp/X3WYieOMHICPgLtTJd1geheBpZH1xyVkrN0PX7SL7HIsQW5Qx7DKS57659+tjCWaCx5g
+vV2V9zdlOUPgzMmt7DdO+QkLClAJxxmw9Y17lONwxQaE7GVgwq1zDj4OnCR/33LCaEz+kVm4U34
GiK4sq9tEhmMhJ3dnAdCYiO90BPpaiRO49Ox//KAcbBaF0QlN43bayGVTomBbIowvNzn00WGT++d
7M4IRGcliDE3i/LSYVRuSJZX7CEwDWnsN/63bhNmfysNsCkL5CmkVD5/vHdg/2Dru0XyB6IOxqSj
5UBpAbEnNTr6iBDCTuKuAZaB6CW7aJVYNopzQo8/xmi9q5PKpq7xu7pi47EcODOaW9s6iGYFAJdk
XnEIgHDUi2SEH2ma/x0iTAD1UaeFcQkwEuMjrg0PZurnBzZh+TVf31OgcVPKy6bESIoh3fBDoWjv
I76xPJmx1ENHymoWg7HCAnphbRC1JmcN3PQY9u8v3p2WCtThqdAhXL8HpMy/OoGTnZyizLZWMM3v
V/MX2GLFOGU2MwHf1/y7nZetr6yRL8oMn0+LG4O/PQCHyR+GxAJgPfe8rhM5xRTTqJXYuE+XHqbe
HKFAawSnamZXn4xOYNkb/4YmxqKQDLKpLF8P6L/14f+k43ryQhRCYyZpGjT6Wz9ZhUCKsScdXZLv
6dT8C64ho2VuR1SsGK+Him+pYJbmzSSFC6yhN1oTtmoB2qt/+lVZvhXxUpqnRS19j650GP1mna3g
AEALSDgyOzy95ZC75t5THm143Ywr2Gohddq1Sk2WqhOwISgjGSpYqzPDNApGx/Bp92qttEHyW8gl
fh8tlp5PJrVIJry8/blZnaUI9nBaKE8iv1zmEpf3JIXG/sp56vwY1PMlhdBk1eqL8omFGLW4Fwyd
4b2N+lCrbX5QMiUhLS1Fdkq2AVmT7C9m4I3U4R7orR52ieF5vDKk9RndGddtKCu97CsMQo5iyynI
f/Kas9+Vuyt8utfHgkQCdfz8t2ATFDFWOaQ3ZSJ4tNBnF80LMOP322cBHI6Vctd3hDavbbKJa2wH
XYmW3bLTLbG9vmhalFgxQXvaM0pkFU094y8GztjmT9B3WXOvvzRMyo5/+3rcvYgSMJJorWG/ifGh
eJ2ixtY3O2jDqDDKR+P6CKAflgldp35T3z5VKOthPnvHB32SZFuoX4VMkFHRl4uDSGxoU3vihFKx
YabKY7WF7prqpK9ryAZsVzeyMlGhs4nNOdyUbDhZSfEcPpKXzQ04HYV+UeBEP+1amU1Rjpz5n82L
psZLjc5S13YBROOLdSd7i1roYHmzPhT3YwEUc/bzueeXD0p8Q3B3bM3C1CCK5kDCCzhGux1kWaLK
QGdzQ+raHNaTSTJhAg1p2+xsPrrGmRV7KKEbKxyOvoyzGcfNY6/r00q75h0Rd/iV0MBmo4189G/T
9MWgRvabNQgxVk9VA3DJ/CnphXojwWDJdHCDLovv0zn/JSCCIMl9tcmzdY1rL8pqZNVGjOCMtWgL
AheGv0TI+VObyHohi8OaR70meRWLFP4WeakPr2XcUJAtPjKi10FSG4MU5oxxLpf9/oqJZxgG4afy
eDPosutIUyctg+phDIrvmMfPhVfhyPAPDrlGsWeSlDlVNDwdUaqRqP/g5kTsM+bKSYpgma1d/u4c
O8fqW6erfT96yO66PzzjXSuwLvuOE+ADRAemv9CeagIYsaZeFTJHY11qv2WB5i5bzNB6BG6ZwWrF
m+vUKcyAaWXleIsEFojU5SFIQ48y7DRSEGzecSBs/f9ZqSNASXaLKLhC2dGaLNv6QIcUDZ4pymMG
k5o07OfrfyeKo9fV1ORRJsIv3NiLLEXP80rALt5LYDjhA0b1jPeaNM938/dv7wleI8fZxTZ4AWlJ
4qJevsNx9NIixVplhp6ELPpjtAU1cfuVO940IRcFLtUKsp6Qg70pzGh3pGNAYRXbvxjmCn9qUuA3
VzUe5XBstIKatnJn1D3C8gwIJeQkYsT/QTAlTk9j1Mz9x8MqqfEptYqwYcX0vxuKW9FoLztHcMgo
cPm0Uv0IzsdHAFmOPf86DnPEjrFTO+R2hPI864Oh6kLK5nPgJoJO8c0mfZOky+hRVYQ2KyyL6A05
jQbV91qkO1llzINd/uUM6icKJVLsNqKucVIRZ76zN8I83c4yi45+qGum4VEniu+9KQ8OJhmgfIK8
Ifm1ScqXxIl9tsmln9uxMYKeGmLuIvwuVCeyslEOEnDvLXa8+6nC8Z4AD9wNq5LIgRoF8Lprdq9O
yIWS4jJYBWo3om+dZzLv/VZ3TydRtjBatSRuIDu4inRgrXAnXQR7asEbn4pIhWCC/uDHGf/SPqHm
ESqPwBKZ8AaRM282NmukvRWSTYm3ZXe7EZpQWA1ZFicbjrlpeXRkc2linooCu+cQeKSR+VKGIJGX
PTzrzlS5afoLRyrUPOz8cfRtFBe8gZfkysRog3MNuzkbwdY8W+wHnWOJTgY1bOzqoOFWYncOhnoN
Ktw1KHY0Ot/2Bl31mDiZnp1//Bo4ORu1M3H4Mmbc5naFNVqd27xiNdY06Tj1LGl6akq+0JluKzTj
P6u9pMyPENEhAJdSznTw33Ru1L9EKLi6kfJZzS+/2DDrH9fq7D7nvpdjpQb09FlFm/tOkmzHltXS
GzyDaYcb5/zYCjH5fvsnYE6wB88aFdte9Y+TzYTrtUT0VMWK0Ijx+kGsZWaTid6Wv2IwS6Wa9PfC
IwEOn+E69Di5gGrljG8YWyLSJS2VN4TwSnTJX4tM9VA33s80gRwbsgfuDLZ2M2ZOzWPYAXm2NYr3
QG3X9OFYylLPx6BFPMpskT10HY4kiTAwtDerjduzFfghGRFE0xbjv7Ud1B9CYzMFjc2lgl+9bycy
frFVyzcde1QoBVu8FNE3BeVvYzsv0kgtKGq5a4xyQkxcJ/pFv1oG2Gor/bmYS84doxQGWE/OxnZt
2H5M5WRtIBvefWLAl4WY02+PU9PmzyGdJROEuD7XkmMxg2Mozj8VhSwQtLz/JW/Flm9w9kJpQ5Qw
u3swyFx77q4jwYMkjaV9y3XQCNhD8VgBo8qGMe+9I0Ll04PPujWkB14ei5pDhOx88kIqZVldtkGY
YsMPW8hoDH5PsRqtsoY0qtHXROnullobwdPlz/8JkiMX/eHytX5/md34mo+TGPKDbawIeX5LfhbV
iKA963TpFDD9Cu3V1jFjUNwgJxSMtgNPs4wfgTcbTMgK/vN0snYspqI8Jhq35QI0NrljMpNg1xdH
vGXcQFHA1mKCX4zUOaNzLAdqVStB0SlC/kxrOMzpNATJ3+6g1GOfFxmxxg2tftXSKbXbYsFZjYzc
WkPAhNvXWq4VmPmuUP3i0V5JAUR5ekxeiLeimf6xwqHg6qoEkO01W+u+fDfIGKBs70MFakx9SGYE
FtS4kmRa1nvHqqYo2stK6oJ+wDaFRndYTRQzPDevr+5HSI6uOOM3XZOUhsMNexX/CEkrsebG5jlh
4F/3ifx8XiRGavDBYfPXyan/RiGQuzP7zWEY64u7BAh6cgVoPNinptIWoyQ1TsiPJt/fxoYDOxeP
35YDcVhG+epOaD2ViAZ4nf0QnUgg//YVtK6fiGqxwy6PquuKv2/QbhIw0Okd6zNJ5TpdlNZmiStt
Wgg0/ZVqBsRp1buP4OYL8gebRyPJGDcwy4ripvj2qCcpkxV3XoWeW5vsiV5Jt0B3g/AWWMc/qHBY
bK7QUo4EwUISEuxsxL54E6RakT8c/htL3R///cby1n6hj//RnLBrDyNb9T5/zZB8p+9wk0AB6XZR
aZiUrch9dJ2xXDTavONtCqnihaIt1neJQx4R1I6G8Lnj219iOrZUGAw7WNmekjGgCjpQGsiWl7uS
9B8Yirmb3hbxPkjH34WIBzSFVb/T+Iac4GXWpXDC7sfzxKUewTWi21AkgCfEeOHh1DtvSDkRXyIr
3Af2iBwZKUMh56LF67uZw/3Ih73Gbr9K+58xQR2oz+Mmuf1RxZRlKDVpWGX15upLIy5T1lOPLFrh
rLLSTz/AFWomzWnqkH8zJ3ZfJFL5n7N9vkBqPncT5FF8enpxwUjEc+bpAxFphsEpa409tNEDDAd2
kvDALEuT4yBNNFW9a1r3uRV0POC1nOlZQowTkGsfm4bXj3BNKcOuOgLsxpjdakrOKovahZYUURBr
5ROoMhysStuVxn6U30ssMzsTqtwgLV8J9162MjhCzof5GkqMm8eap2Taji+uNCFBvWgXev5MAEjS
raIE6S0SRXygXr02WT1CjGJ8+g3v6Os/yC/gqG8V2HwF7H8zBoG1SI0J9NelbnlU8utES8dVewl/
vfe2X+H2TzLM4kfOSO9ZXarrdox64lO4OTYkeJ4fBfag25bR1tN5J+t2cd8h+B//OD+z4N+vX2Yx
aKnPd1OASWB0mCtvqubSNXpp0LI6bIazEb/0Lc3Xp536IXax1Y3ibIpgixxhYpYLyMrFboxAOpF0
0id2FBmaI8E3U00vaNDhD4IHFbCdcSdQNmJF3adzodXVPM+AuisztlQjJNwuN7UCl/gmwMvwYvax
ITLwGYZAJoFaYLQlwJqpHhevTIdoKLxib9LpSYeEzreDkNL8nTgho1DXg73fqta6JyvtBfHageqS
MLjoPuCnxR8d82fkF6148/HTJlTnk3BKw9qwwETGXDobo4GmOaX7DN82MOBCurFxdfv1uNh8Ep/z
uu7EAtmv5MYIbNCbVQfndJca01nwkVmDu82gsd2wLoG1jHsBlKLyWC/ICnIeP95qryni9rhqm360
W+Onr+pWt0jOMzHecpqJlvH69Rnxh9Qp2OFmYpoF6GdVAdrkcTxYO+VO+I5MizHZiyq+MJOnQx8Y
u6LxHV0XJ+dn0YOpwVRGQAwgkSp6dUGyOZDqo4oQsFXzPIamkF3xVgs/zd3JGjLZxU961ROAxWIk
juaDzhsgoEfjra4Ech5p4bUeuCs5jCvzth1eN0FvmVsnuD8cbaLWFDQGbdJk8Qn8/sGXof+RjLlI
dKumNjLv0B9mVsq8YMhunuq1lYRAIQUs/219G1mC7nwQsrOpEtVcvjQB0DAX4+jayzKlYZ8cxgMo
1SJwPT9Y0T9NTpBIOzRH/U2tO4GLXk+rPKg+a4LgPtnPJ+ku/Knu/CG4+AknxR4aPh9bn7M5RA+B
FLd1ndZMk3C0bnqeByzcTO3qLtzo/wWauYTSZ4Kag5lUIkobU162ruu1msniFW/SIl88mvIKs+5/
ANeCdnDcd1sF8VIoc5KCfuOzCIhBKjecJQYSShneyA71QyWOxvsSC6sMd/7ER5QFWuA/OoFUKV88
PwwC/oqjBxV/kLnmnFU18UukqsZO8QyLLBqs0cw84cKoPYHO73CtmRWZhOPR028otnuLEiy7KCYV
5RONiC0pRCCYYYfgFvuy+kbOpTCE8vXlPwhk9Jq1Qkf1/e0hur3hl00LzqtOqc+kwMcnfdd/3XT7
039MtQhfeFn6+z2Exm7SkFEuLhI8lWESVeZ93AnhEX6dpuNP1l1aXdMmZNEC2A6MhUagdNjEXsQv
NCMvW7TkjQtuvQSa/TBRkNJTui2z1YbhjEea9eCkAqfaAKK+PoWMhKZgVy+/1GVpQLVKtJ4cKu2f
ECDZ+GYIKbNKF4zmhSLeDrLGJkKeb7orb0aJW35r/dGf2PW6wuOodceJVNmclWOfuJe70c06lv9i
mK/p0c1Ft3rOM/XBMNz7+8By2aN+IF6Yby7kez2J+kQrzKWzkuX8LCDvOsLwGHzyPHizkUxoh3fD
QMgROKG0/faabAQ3oBx1MGmUewoMslTC93HAyJ/6AV8G20C8PoRRbYNNJwUXQI1jH7Rx6SHPqJd3
FwX05JtMEJyzx5nzDOUZnGJwpZQtsgDiubL/1VI0bjRT5pFtuQhQUDziGkQW2RDvn/cho4MA4ytc
Syyoai7qRkIW8T7REFoSGqEHNEPs8dWk94iXubdVIstLk6RrPxpmx4tYieq1VG0ZGg1kmfXAI1Em
0cDem6ClzFXdZW/6FmVdmruirjhXYMSzW3TclrEQhAvVD1W/z6hMsLMKfNgqEWt+gbTQF1ImayqU
HQgcIaOXUuUAMX0ueGIvIk2LQrrgzKW1o5yBu5faD1em0k0NHLIolHklVeerLmw9KVwsdtpuIB8v
liWwA528mFpgTRGj53AQkFd5IsWWgOOrwLsuu2RCHzCxONxz6tdB2Bska+XvXVFURKKGf2FOOIVe
rElwyqZt5NhpeushZAJ4V9eRAV5KWTnw1Co/FAVSlOJGKsEUX9U1BxBRRZ8bgW79bQ/A6oFIToBj
IFKvYMLhUNkVMYAydNEF/Z6c8tru5Qn6YhLU003XINsqHCYL2aO+wFNJ2Xcj2NRuikRCfOZrBIlv
SpayFCclkb6nzsIXUtXvn5D8Ry0+u/WG3AACL94GcVrdhXoAvL6VOBhyOQfSzT3sRwK0lzOGUbgt
fenfwjIKWqAP1OR64dLpmUMQSk18DwMz+4IH/mZq7cgPd8n2qHSebcw8su7eeZVJDPuUp4jjBT5A
hrdmjil35NqU5BBU/0IHvY5njkwrsv5QPSOBRsFoZR7O3HW2cUaSvPiaZ7+D7GzwbkDqxu3u9SCE
ZEnDa3WJhSJdsBvBMbQTeughZwmWipQfLhGuPiIFzl3dmCtjGTwWtoGqMAbjWglTu8Kc+oAx2eNA
8u6EYnAo+FycguLCenAA7knj+UBkbmyoDnBRr0k83ZPvNdSMoguOQJxvhbME+bkxldKpQaO1xyyX
UglrCdXBiM16nU3M1JleFVb4iI88Gi8yHg4PxU3RLwFza2j2SaREgaqkyumWUc02MX8n7o/8S4V7
MZSfOy+mwD1cSDdKqpM06KYtTZupY9RTY64A7dOQkV9ndKJsUsNflRPbhYHV1bQQGDb6AoBZkWbC
OwR0EuxEZM8m+Yhz+//X27xT/6M5If6MaTphFlKG9SISuclbOwNun5mASfu0rm58ycIFjrJN25PW
lZ7/U+hGJrOjY0qeNVy+dd+/i8/Wb/ttOAOZlNn6EMNO4tccAddDfklbMqttemX+pKe9T9wBMpII
wJzAXSxgnsNF2MtHNm6LSvTvRlxkIWaYpe0pEhvMx/rCgI8YKyZVIqb48wrV5NjLcWV5GsD3DLKP
8GPJDUlRWymAN7M8aZ+9b2T6EC+yDkr/sDAOECuYQxMl/JXIqiy+M4OiY7xq0OzmXhf3QVXD6mZ3
FOsIxyGRPtIxyQYJtuQ0rqm6kJrfSo3iYUTCFDlJX1/nj74KTshbi1rhA4LgIuqx3g16NqmNz5Qb
bycnyxo7ZU1blJ0YvXulxXsbVUJ/0xUJWLD/ewvzcZOVsfDEYs/dvdUYJglkvjKEwki7+ArgLrN/
bB6ESoWQTSMqtwGMBbBYbWau3Nu4E7ddSEBwah7CDg1SwUq+F3yNBlDpnlqJOiGt2cW694eH6d1w
J4jKYZCWi89fULEa4g++2LNfz9oN2vYvGOVEL9zP5wpdgWE72EQcDAI0Rrby8Mb6X0VvVHsAcLd7
i1I6gJoYefVu7y0SWwNWHklX/dLba2i688kvBEWek2xs0HQWUtTi3f/OdNYA3O0KbR/cFOt49xGZ
Q5cI8q/OPmyqVX5VH6Ci+kR8pioSmHkHiGX+/DhFFMmk9cxUxWKJp7Qhz+nMQTF84/LbXOHUr7Ca
K0aOy440TaNX/U7vFX+1NfLFR5OeUuxlwkW87qBASvhreWOYftlFLbbYM/qk1nWiTXXlMQ1HuPPc
yqey0G9H3gXsqb+EUJKRbBInQDQBiDy6GQcQlojoFtzxF3r2ToXOHZ4jzbB7y4vOLTTdqPawb9D8
BzTZ/gMN+Xhm3sWVSd30f6rzZ0pC8i/vzI3Mq9FzCOSssz9of/95ikozFPK48pr9pOggbkXhyV3V
+XENh5e7223go5k7wkATdmDBx95chgL/zGpDdbWsPeP4WKMT4Yj7kAtmc4p+Pk/hf5CElXnEVpsC
G0zWU7ukzsWdCvGQIxQIexkeA0jeH2U+zeV0T9+HK75STo0I6mgf9uAU4LMim/uVAkeoFXBOap/A
ntr4rSn+o8qwkmC9+8HvfYCTikXuJpE+dmzVY4UAEX9QvkzQ2rOgHIVAykp7SXUsR7a32fJ5hnna
o7XOKGv4wfH7unadJocYwvbhLk7iXqAYCJPZq5ckxkUiVjUGNGDG+ezheWTKW4rCdSKtcGucCjyj
TMm9i8e1Ec/LTrs0h8uLhuuyBEiLT3lMG5eYYkAR1aVAPSMEy1OoDPvPKiDsd/sl2BL8rw/SHE9v
GRccdhrKOPvfK5kn9bXTmTPDqrDfopMnvdYH8uI5Y5WGExNWvqXeVRAUoWWdk/m/KrYZ/kEoOUMX
dNHwNyLZF0hXm34zAZQ3p9nQlRgJsyA/6Xu1/CjXY/0NXnkZkA9PY94oNsc3BZ3Zlj2xB2+NSOMo
FfrT4ZJxjmmjiDelWpZmOeynRL1cIke/PaVYXFMEC+aA0zBNhhOuBaA+QCKEIzijIqwxPRmtj7rU
21F3cmbtFbFZ2M/Sjy1KaoWmMD1ffiJ7SIWHpwT7EpKXSiledGl4q9E47d5kNC4pUZgO2718oT7l
NdNP59e8CQDlSvjXcg+A8Gao+L4sevU2mKVr/GZGl3+iAd/h4XCyilpVQvO1tPgUbOa16aWHRkiL
2uUCZpn1fX0khuWGW+p0KanpS34XIuelgqyqUupmBbdiynSSGndRz/S4T2hAcfanbzF5iWZyyQNs
S9+dnljIJi4uii/7IYbF27vcYFwDU3Y4PYE3rSe4Kr9Ary4MuF3GGN7Z30XXsL5JCPSRF85wC6b6
/JPQWQkumhcLk82mA4MUMN4dLTF1Zsp+2hoR+DdjNZqOKPu4y8M94ojL8B8z3yIgD4wxp6XV5H0h
MbVMuBUdtERI5rUWMIzcwnOX1F5xBKzRImKDpuvPACELzZWa3GTjYdm7iPcgyle0J7Pjn5DScYy6
ynE7uA97aeUKApF/w4QEvkAyLPOGwJJ2qacCihmWDHPFJ9sWBN20zWUmYRfp/4Tw/LJo0OENa2pg
tMrbQ67yqpylX3PQEMDzIYiqw2wFqogKguFUZLOnTum4TnOi/fDZDf2hLaXmpraE7VVOvbQ8SEwh
aTftCU5IpUTRicwk8XVdE2b9N/Pj7YzDHnthwEUPIny/2J5MQfjeDFv68dBxrPdQf4qg++g4z+sF
KXLY1vFxU/5Pkyh1smUAFHW/7HhX5y3noF1fWvRJVrXdbDLEkB/Y5EaXWIFybqzdOaVbMI9WaY8P
YoVCMml2FZk03G6+pLQiLGtbQPYo8oO0HXnXRWU9BdA8Q8EP96SB8zHfrevDgUKZFVfazc/mKYt+
F2ETG+kgUThLURSAx/SWNMyehnPdS5HFvBD5moNITX66VUab+Y0/2bZ6Pu5GSztNJjDFyOBCZyJ0
eR5hloyXNafP3EEA5kXqmUtnnjJgldCNsLBRm6tiByn1Hs8Ni4ziMDzIVOK/sO4bDJBv+zwTXD4G
xorFOd6LwyK36Iwpz3nfdbklsN+JP0TXlgyo56cNiewkp3YaLFwHnooMTcGkCW0lE8o/BEQjjAI7
Gl8ViMRaVEy1lsWieq+lkmDdMCOVd56FF7dr5zJ7YXJZtFp9j0APGKdp8QQm0UKvaYaENCFk1AcA
hOiZru+jInhR2dx71hvXkOyGyJujqZBSHmD8Sk/aiAw9TpkEnEekh1SYxA96DSKYaQP7UkgMLAxm
QHtM76/JzeW9V/afaLzl8Purkdk1VNB7LteaFJQiWiVyoAeWqCtvhM1XqynJ1os6nvynneCipsbF
KtTvh7ATbi1jb2UujQizgR4cblMrRE1VZDh6gruf3naFz5UysvrtaFml+8L9c0VMMtS49a7TbkI/
7RNdcLTqkUms3CT9Jm4QP0WTjuuDH1vc4SEKUPaoVIooRlFy0TFrqrskEt3vh31HY0R1WxHlqdjL
1L2sYPs+cnX6XihWicHjWmS4MJe+Xb7YTGJRu0yG1q9iF1TessBzXozh8wLUu6ozxOfWp3L7d4A+
2BGe4Jiq/kMzk24jXl2snYZPrZrma52Z6/dkTCd2zs8tFnhBcIunAhvFlH52eDk/7HAlHOE1GHrj
TDHXWparqwJW8eS2lJ7QIbBn3TjTyb5oGcYfy6gZPdDw84+TGq6SdMISTeToEmtHuKDHCn+20+2h
npYK2U5C2DToqTLNlGuX9mvKgcxpGoOO0IEUySwHlhINOCLFFsI/vJG7IiTHZJc3bApaQjEtqmcF
5qKDY6nK814V1qLZIg1RZQchBMAnFPvpjGlUSvFWMWVf+CMq/fK4Vixfkah/xpoNa8jw6lCWVKjI
kIUJqfTt9Mf7bqDjaexvYmtwcrJTa5R8aNyxJtAvahWROo7ypqMqbxaYkwqcRM6lSmQUmGc94Znf
MObRzsc0smsmgeiHl9JNJaVurbtMfUt4VjIVz/Tf9qG51Hx2v2KbPGbEVNNbHid9D9yPfrdfV6KL
lHIO8pO8DOHpl55ZBn+h0z5+UR5salD05d+/qfv0trFxIbSnbeJ3jk2HILvAt5KQCWjliZqrX7qH
buTuEJ1aZS9XbcUyAfIk5kXrnNJHCwjNTQUKNikhKstcKfnA7ffhg+2JN69sEr01NBvt8kdfLpPj
Cgg5li1L7iSHtqz1pZ2mkmynCXkNLEB79Xkm8/rYYCNawqrRBBEqCAUien/jEhAsttSsh3wmeBg0
AKtRyZDVA1r3jb8MiwHwFWdbXc4eChvqR3oDpIvWRjFtJCJVFn4yr87iEUBKPjHWCNBh1yHf9w6P
8m6bnRM5WAoiA1lqbL7x7boIQYhLmrNhTwpL/Opi/cBqKxrM4GrRtx9hNATkHPfL29EYteLQQhWR
Uox2yMetqSagP7Lp89ijXGGtUniZPzNVWM0ZhyL1H86ppXsCjVFwhejEEc9ET4PUczAUzRaOUvkL
/TY6djFrfkRug085sPAx9CcprNx1nOJH2AE4U7/jkLWokdV5hPzeJbPSYhbLAH/Vqj2BHva1Hov/
8/28iaRlqYzL/K2DBp537OA2REpwasjEBCJScP6r0SpS3238SOrelIfEAV3gqa3+Z7sEdalXoZRy
Goku7za/PBu5ezXW3fmNMt2EBMK1WxXy0lIaiRO4TeaQLl2EO8rj5jnx+AAbfzfBYvGWzSU28Ju/
VC/Z4EB3enMIsJzPveJip5pMppklOolqsvkMB5z+r4VZkBX/q1YxC3ngg8tA6HcGHhAfH2+jeGKl
qxT9KIXykvu/4QsXrqbqG3WUEaHZvOsilAuvz5OiF/9OmLSgUySSyKyp2qWvHttnZXVVtM+z0fSu
5VSYmXgd+IzZ+IAottkRpkN0LiSrN1TVtIc3E6IbXgTn4KiXQPBc5NzBFFl/SS2MsjQx0IVrk8GQ
SWY+t3okijJ70dfvXZf4T/9sWUeNhpPVrirH+p2zAzts1/gGVNG7hlb14w9hC+xo9f3WIPXEYz93
ze6L44Z2svE+JEiZf7TXNW/PT9S/GseDLTZM8RLvFPvw0uzcCPoAjwUYb4bYUM0gHZZePC9JPryA
iPq7Cngc0mLEN6P1hJtwvzrUq/YV+gY6/ZGTfrmuXJnqvA5LYy4fBqlYFjbIYQy/Yo1WYF9exbYN
DF15nx1eh837JvQDEq2dMQbOKsXnjnPcdudX+lOWGu03a6BS9ctrg5AQsJBa084hPoI2VZiJE3j3
CCi5dVN8RtCZu20BampwM7/ZUfxGBlp0JkZw/0DsSDab4dFUqLE/y+nczRS/cfLHw83ikwzIm6bA
7a8zN0lrOtF6YOWscN8c94Qg9WW62OY34biSF7bvwGNGvqQXIsYBYqAWUXGUgIhqbzqQ+zJZI54N
Fa2DXSFvnnW0aa2hwotmXnzeSx2kNNRM0kfQmYXHAPcoFSkS+VPpo4prv0triEQ6eFHqAaCtG6J5
CvmSZFok7quXqys4I5roHO+Tc89QdjWuB71ltkDQht3PODGC5FH1RbSSHlBY0VIHPUvDkNv/znTY
pIHKjhd+huZITME+nQHTgzeBJ265Zoey5ErSRTDITUpF7R7M77seuQOINVNX52n5LTYqNCW961YF
5vrIj1vwfLbSn9ta2KEy+NVKSVLAj+T5QliiWG+UjjSqiIoMBw7hTiTpDyTyclY7xVEPET4hB3TH
srON48i7GONLzmFC9ziEYSjXCxfdGOJ18BGHKu2eRhF811o2hlqv+9JnNBkX0x07Ez2879VifQUV
2+2G1oNnZ7z5n6WzX5tqlgHbkbc4rQNu7lTm7aQ1M+tEH7FiDZ8yco6e/IJ/507ECYqHbzuiJxZv
+1zTuH4fk/oTW097P5eGcpOFiiurjFQrZosVPP7iZEgJHew2PIXCw9lnV3eY0pAHCVFgoeUQqXgc
nHgj2o9/11QfHJioJaIw3cnOpfxoWpB2xjK1JD7Mnb75WOQlW2/ovDqbXjxpqDjVFGQF3yEfk/0j
nQb7EK6a8PevJgZJ+I03PpK5jKzyHMePAiMOOMKfyVOwmURMPLBY9gF3SOibvTitw4q8mrLE5hBA
R1qcfHZ+OAkm/hTrDrowelVpXazA3mJEH/1q/pJqbdQC+nyQabo7njD0IL8t1fboTOhYO7BwMyZ0
bCtj2eAmxuHD9ohdZEI8tgAAAMW/KYwo8QRF1seNa0VVfGoybWMdN3uK6nIfeOPcy6JD+FcS1SZD
B/j49nvJOqPFFX86BhQs0naGjD4UDBOSCppB5wTvWVIX/NVlpvAxBfCW7lrIx/tRDJ9OHlvjGNHD
6NptIMdFBrWbaXVeGyDQYyq7cYA4b7+b6j6iEjVtlIao9oEUy+PFiDTCNlEOXU3WXXBHhoz3zG25
r0+IMhNJomulu2cvMgV/kmdkZnV85vYo3bwbx8wfGZxNp0MmvxhO3O7mJoWu3uM1t1ljFrrfsJ3G
141+wWgJ8khBUZbTaxWKXdwnzYwCndQ/NTfAWpcWLs9dVcL+Xlc85n2UjuSSjKa6O9esp+Za3C8Z
VK+YFa7NjZ5+WbpfmoI8rqUmmvyWZfMKPp8oJGXeg3fCnSGNl8eggIv19mf79NgqZzgqM9Us3D23
w/g7igc0NvPrDkHFLro7qtyiVp5DkARCuhxsrY+GfuhHi42HhyUpqJ7KBzCOP/IbUnWfTwYxU/FX
fUx+ITVQ0Ru4QINNenISiWCQ0HsAOTXQKS51DaSJaGjChNz/ilTyeJp0ApjX0UOr3blFk9FMR74C
WF0+G4KOe2nWBjI3QTtB72KhD7f9uGajm6tvPTnIFjGlX/bfhf3KydRnQWYJ+qqlQ4ASZ5jqqmiA
M6WbSe3QihZFoiBNIKxh9PGlq+kjlv0u2FEeUIgO8+sOBah2uJRBusWn5ukVp8yNDg0ybEtqcEsS
SbExvS9Agnhu+kOa+fJAgGtkzVQMy9Zwfi2XrkPh2/FPmJ4XukuqM2wJR/erZ80+Y0RlBs5veYep
aBS4jfwe1JXDwZf5FYbC0Svq5b49/SAwL1inOlnDX3tHpYKutM8VvhVm+gBzii7mE5dgXgiPKOg8
+Un8b2uoPepb5kZ+K1G5nRQGxx7Pfwag1p4v5yrZ2zodhmyJHBcNm/FanL+oDgTb+OLNtplzlF26
x1Y5KicmYocZ1GSKKxjDFBz5fmCOJ3XWApsk9A1/8lBGpH4HcQMPDZrps80B0mExQ+jvqbJgiFcB
oilLcdW7m5/HPpoyOnJA4A3J+WB/fgSvLf37hIswMBa68GjTLLoAbmN/aiTfKCYTNTm4eQJunB/P
Z458zPe2mIVzmdm6GMajBgSQ2pIqX9FF/NyBMzQi46vt8/UbsVlfWf3MmeNgZQmxoZa3ZzImcsDD
RNgl4eYQqheUxjSYsEfBmbiTMe9z9Zo9BhBpt3kPzQ8xyyVsjSwPojGR0awe/6JXRlXW5IKaftDF
PaN2mcqQtRmVZ47LqvH8DwMYlKwJnMQ8jSIgc7Oey5wQIjrraiQkiE253OjKWQCAHarisEVb9VBY
81eU7dC+mL54YieHx3OhKz2a+BE20xNUiGNOsj13biNbjmfAdg5Fup8u336qK/3zJ58hyH2ua317
KjsQMlZdEhor9/gTmWEljIHhKfizk2FldKBcfS+sycmxacX4O8A8CfCpMlXYcFOZYj0o6TPzIN2z
Vtqe1/6tt63LmwuVNRJ1Zwzrs/7BOfXreWUEXo6dkAuTGQFQ+YzFrJCGRt8NLtsr+7SGeyPcVnrc
ElDpDMKEL225o5ooZBwLBqDkfWEPKPtuG0uZz03TE3vhL6Vz2PUDQ+24jh5LmYUFisLmxO5k/iQr
jgkwG5UMS9dxLjIq29LNiNjSZM9VALSiyKoj9onqw1neGoNpLznoTvFyfkjV4XeYU6Ye55GQwCt2
t7BtUnfKzzuiJUsjbx0mfqnXJ7OZ0MEJJb3dzHX7u18C7G40LyElYL/R7XanV8BtHTyBnM6wLaJV
Cook/AWdyGlV6TIf2VTb5qm3S3i76uJCjFTkl9+FruXphDMdJL5lkZjVFkm5QYWrTYBY0sOtQ1wh
E62VNLBcyAOEVfK/JOa7hxD2A3afUeVvc+5BX5mXkJvQjyUS2kuVT1UG3iPgqEagJjVpAalTGaQM
5LMlAzrXwUflJ9X4uXEgJcqnxDaUsCJOkFGywQzoEG/Q31EK2hFyRsgap6wnSVmYBYaNxVU1AHRo
jtsKxT/DZlNNCRl9hz2xH6fKshl5KHWnd3VEtd+uFMLtssAmhVw0zmI0LxGH6O9XE0YefZO+78/u
LRuLmMeLraETM56QSpkUVsSC9vE7EMzwtobd/t/eflbvg9XT3Z4VLiVnsVRK8c5XH5+clSBZHrO4
ZP21tj4nnpRfYiIoyOnhaSRg1cWplM46xLG6RfyaIpFH6f9MxvB+UFVB7buBr6I2DRepn1L4jDJz
RwO+R0mqgWnK5IttNEjU/L3aADmBWMkq4SOq24XKnNq6oHyDGGeqe2gljLvKFdA0NNRncFxrMxo4
CX+JUyRHmpYJa2B6U0xjJZrHCD3G/B+iBRVC8hhhB6g+l4dfKu6+0Oy2THzXNQJo2KWHKWmLu7eg
vMKczLoXOq/KdkbqfeAcg395LyeEAaRc8usE4V6Nx08cNeBYhYdnrnBgsaXCd/aDkUpvcgIm+ibS
iVzHGvHP7kfZ6ybGr49akFmoM+GzPLTNHMzR7qzYtES/n2j1CcvmOVXJ/66/WM4TdLx5Z7Cfw50g
RuyJslo63pHn65bx3UR6LWgp2rmCKabXV176Wo0gPTDcDdtTkYNefy5J6jbU7dny9ia6xnEp1l2P
VPe6E1PC7GJlfZ9so+NadGpLCih3UYSdTiQXR/SFeyk03fM5RX7CjuIPxRcOFKREE+uM7GkWG9aU
1fDBVD1OFuwrjImEnIczIHiA8RH3QBPiyRBv8IPwNlMOlIHdVzb6gEZKLeI2dtxk0pkJ/bgpd9Lh
ohXrghTO1RFx/d1b9pugFzKegoPklcsWWgdX+ebm9b0d6kmLJcHYQ8fD2GdvJiMF0Eb5tSnGG8WO
vsyLlUMhkyNJ76MEstcmWYs7zIYd137K8i7oRBtIHRoo9igGKGXG+UE03NQNtE0zHIrNOLeqDqxc
Nwl/0uEShR5pDLDtZyWCCUuchC2XZT2p+ClDKDPO0rQXJFyU1ZqMjcYgzFlI2NwI9GTsBbI6cH2+
mrY0EFFSKv+UZMwUzpkjpXPwl/mAXrbxqZ0qTgSHIvLCm/7SGqbfhQHt0gSAaKsY+lJRUOzgac6n
hyjUDTTvsOz084HAacSlGDsWxz7LQLUz5qnvekCgy9TIYpj4WImoIFpG9K92Bahr18tQWqo7UsdG
idmZFe4dIJX1mcayF/wBs/YttqQKvcuD+W7Vy3RE0slrl9aa37LMX8prKxh2iLTufre46lSEiyne
UWf050VZifl4URfikjFPvieU4ry+eWOTEPmj9x+ole7aaLhNtDec5riIiip8HSzwQPPzjQIv7eHm
KjSYkd/R8zP+hotGGZvXlGguqyl+/+tIWPMxNX5fmwIBaU5TVm+pM8TKPn+kkKIUK9+3ARfdpehW
NChwKqXsdk0asckHWCp+dXINvwY/Kj6yddRVwoNLPhVLrBnly55IwMWJPTR87V6lsw6kUVpYe4R3
OmlYj960qKZ/qvOR6PGeyBVd7/9y1S4D53Qj/ZpsXmcT2JE4wnOHFp1eE+I9s9J9WcXj3umYQcq+
18gRX4Jf9AfRiF53idLCkmWti2hN7Ws2Vo+z2R+/pFFetqs76+/U+G8YoM7SZSkV3yDJdHwN1pv6
bAXfJ0vcMWE0Vye+dWUnvJYWRNRLERV59DPUPAx0PInOq86zW2du39HYPv7Kr8douRMhlQYOYL/5
Mw0JasSs0jfJsMApCKEqo24gY15oX2sApnmc5yu6XgHeh0hRBO5325FXC5c0Qck7ni2o32stfjj1
PU2frTejIifXcuKFMHZzHZP8JVrsuNLCoHBiHp4+wzpkHKAejgW2NoG0gbhzKZ9K5UGjiOB6G3Wl
/XB3JjtV7ZALfEGeofQ4VUv2hNaiawqI8LIHifVnm5sz4+QJlhHIWSRwBA+nm+KnX1latY/tfqsw
oPwIqIfGBeNcOzc/kzFeyli4ZEWsDZi1rLVKGMTL4q8pjzMHrXishhix6dkjebZ78OMZWzbjfIk5
kTr4vN43uZzW0cQsE9Oju3TwHjjCM7/4JyQnuYfnw2VKiqyjDfiOdeu4Xps9Z1Qx9QJdGhOOuhv5
mW+9rbh9CDJEk9qzxX7qFcs09sxo8ERopUGa7w15U6fVtkY6/VCo8RbCvR9dCwd7v6vgrDjW0xMi
Cu42npb1ztanCMlnskJZzHE/iwHnwz7Oj8rNCFKNzMEcjpmbA2vg+h5OaPXGl77jhcSs9gIb6tsm
Da0+YGZRLifHl0W+kQUoU/YeWD300G/cExkIu0DsI4a00jRGhW7sqlgpWgDDtnoG8EUva4vVzP0O
NBcCfp1Gsogm1r59kEWH3+wvOcs+iS42DmZQHUNykBzXtRX8+naZ83HAoLiS3IoVbMdiQ56ah48l
Tv5uXHi4uz2KS+F1NsriU3evoOZy5Z7irKMrt4vX4VQGcTJWbDEoQn5NPq82C4rSuob2tCrde3lZ
PIPBPzxF06kDie0reGS3fHFkHDBixli7Ys/19ZTaqn5I7fnWnJ670CoTCfEnkMRBS3XQoTsNYREA
5zVg7k/UxwHFHOZF8QvgPdqHBlQ/UC+qS8+MDYjbE911EQGuGToivImxxyG7GbPE8MsC0+MtyFkf
iuS61ktKOgvB/rEd2aGLMVsdqE2PLi27p7j1oodt36yatcVO3CdzDlFWTDBSzr+dH68iXLOCWwvo
4gyQV5JP7ftelbep4Lx6c2mHodpahSLStTbbm8pSfzd/TPh0HSDyT6LqdJcuRHBGXIIvkxuqLdvZ
hdSDBLZFDc2FV/KkrwtN9cbbfwWfOlQoQygRNnfMNWVR4feOYlORKZX90sOj7qI5JcuuqAaYqPVh
/uSArrCQohxXixIeAcIEJ5KOpYv5vobAY4aw1eiIh54VbWgpMjtOjBMorkQXG1HHCMiqPbIbBoBq
mr01C0ZCIci+lLBEUZ6MPSHCnLSXVV53/lA7gjJF/M1DVXWzbGcItUNRtSVvkJY+GBWxogO5BM+Y
SxXP3ShSlWLKVFtR7T50/7Nv8UuBYtaPlCMbmq/+hVXYhXKbnLPhBHiABgpOHcja58jt2XpY3VSE
1qo/epffkfn7D5C4VAjSh+n0adG4hKepSQM9fnrcRkRV9VhpNqRZN9f6r2k43R81s8Q4nT2/frBf
q4/WGq3BBGHmE22FRWb2+6nRDSd7rff7T/tIjl1TNYPwtRTwKCPCb7YXEEt7GWLF5efLihEzTX6i
kC6ZdwbmAPdIa7jDA7eYQ5LNXhQzh1watp//ndr+LIB2f29i1p/K3+iWXZo7U+fQ7KBZheFl/cdT
WFYCa+6Qlj3fbwS+r2kzTA3Pl0MoUtow39Ap7VCCUK1EBxN35y73nJjHQaPDBSY/2WPMGoDAV8IE
4itSZuNUA295hbz282VRgPQNQL5nImlZslDWee2eN7RIgzrdFEX6mbKNcD7PBpSsuqEo17RoC2tp
6NAd9mGeiJQmZ8y6nv4zHW67RRBgYs9J0agiaXnD/day6MW88XA9u6PJVPSoXCiUG5NRdtN0GFoI
bKU+mQgTra6bZ2eX0Y+pIaL/S6pXBA09pWTszdbaTzJsP0/e4x8q5nC9FsQMiakkkn4DWgaodQMo
lpLiJEfCYIkkCwdg3Ze36rOe/oWyDjPzrdSnEvaLKXeGAUTI1AcrDvBO01SiNnMEiwWwZVykDJVz
Oi2KUMkJgJibPEAb0j1LeTXXeugEUTSTxpvhLiDfbTbWV8OWzMR3TJk6dcRYkkFRD0SVvLGfNJuS
ngnFKC5JaVp9gkLFZ9itYDfzXV9LYnGRymtmAjCwK7xsBlH+k/0+lr+ylSYBcgeDMkDkGMku2/D2
ZSOrK5WS8dS6NI9oWAjf9uVfbvqK23hSdpMBPcEF4f5lIWmP2C8EVrHKOxG596sudLakIAwNgbAr
kxqUA2HwwIeMr/G4XvviiCt9f83ONNNxulYOK3qEGP+ta0TdRpd34c6WfUXKpkT5NkRYopW6+mtE
cDVJM7Pd0mIxCtOysrf7HlEDY6r+bKg1Uh14TKTbvwBBXGdCe+3jFeK+y6/fYU+ABA7sYd5FB6zN
KYp9t1S1q8JbKmF7LAYA3P6NGaRI9TZXXKGTGXZXnANUQVNXjHlu6QJL5R1jf40+sRSuinHMws1w
EZ+IPxry/GTRpoBsSj2IJDbMh4A5u7Z2MjJoAqOgNCyFofMuxSjJ4a7Tt4OQiLP5yDgu+rNpmmfl
KVKvqin+qcMdZx4nMZx+GGrpUW7ABIE1sNaWptAiCgitoHiYIoDt7nresErdzBs7gaLe7uc6hUkv
P+nXDS2oI6mnXpXqglpZcKbgOgzYyR0Gis1ZdbMQoB+tFRT1i/sgodhcNNyBd2a9n9ZPlVzCG3AK
3oN7vpxIgkD+dnDfvDqaIno7duRLWfU5sBBVYGr3JyivgRhQjLRqZzUCf2eWW2MNzWsqfl3Wo/9m
k1nOGfvJzaMkzMnEado+5zUtRN7B/guvYiwsRV+t27BUQIuBt+zme1m6MPlopy5dOrJn/OXVIBQU
E4yYtmg+QBlbRzho5XPeMdrpL3wSHzFuEBsekOyeolaB8rbnBvGDsYKetJUDQXwK5OiJuXpFv001
2Q8o5xno6jPnIQgfbk/dbX8+auY15fkcfIAokpZaKfBCc2/pZqIsHDgDYUuFeZ74gIbj89H35ErI
7Fy4RmnUYj2oLC+s9Z9D3J6kiQMQ+qDjd9qE5wKOyH6nFB/Kpuame8uLHNQiH/I3NcXBcK/Tck2C
0Lez6QeJPUPvQHvuJbGyToTV7PneAvY5nrqXcBDZ5P5r4X7IwtK+QZ0ne8aQQhnrP+HhU+QCO0f2
ML+1cOFYfjn1F4Qhryt4Yr/I0K70ReEgoFIr68Q6Oz8ow4ykIBITIYB5ySC/LKyoWnEwooxRyorS
omm/dT4qoSyh3gH5JPrQKVBgeHE52+nPEMfstiucL0UrOyaMZ9TUj9ekOnjeMcfoNCyrHk8GGiyc
FaqmeB6/Nrgz2gLXXottGViUJBDPQw1nE9uqcWYUUejUrWP+KPUzQ6x/dEMuSVJohz4qMLqziSB8
v4xcPQIy0jv7sA+NqMfyYHxPMY3Wi2YISk8KYOYvN9xo9nHSt65yMxPKbavPY4k8TjEVfYrn0ecW
FYqGWqjLIvJFl1CnBlNWrPoALo9/jhqXbn87KMjygLoIWLZ9Y0qWP1wf8M2YZeaMj4ncEgDB+p4S
y0C+CLQhf6xpfk2lfEMN5w2rltA/YR9sdA/YQHjDs4f6IE02BPp3naTAGXa0eL02gMmuE3j35AMs
whetBVsxo3urOkQcgSUyXutnn0SdeaYRgxs0IXbrJHIsiEpvaKmhy0+Pqei/mvy5CKxObIuYHT0D
l3Gw2lTDEznTQC+OWhs99vhoE2XZEMKaMdMsWGapk8Idkc7TjEZDJEeK98wZ5OAYAyKux4UiY4bX
ESEqwhdX1mF0OO/ijb1lZkless2xe65eLT4/syakX3QMqpXOqZiGwlsdlw4C2so8R85CdupZwj3X
G5/XAejHH/kmrBClGcWKjPv5NRqU0TF2OFZV1wKkykFta/0Bp5RbbYXxyFxg/8Rz1ed246RU1Znf
nscYsI52C5Y7NN2M7v0s+1B+1JPKte1P6MQbHFYvcAH81J5lNsGhBPdeQpwXCYGS/3wEA4JjwxPo
R5KDmawXnTw8uxU5dv7ypdXLveKnS7JDsBPwWSG+KPccGtO4rKGMq8j3OYnGHmXDQa9JBcb5Yt+k
/MbOz2q/fDYKwgn5AftBZ+q8rXVMSiSJRT4br9tq48d5YiSeRGUJBmSVGkpWY7eept6lSEhIKBIT
VJ5Uavoiy1FXbyiXOEpmYpcPd1aifLPv6v9YNaGRjKwfgHfHxzSUnTuJddEVogRzTCZyNQlEL4A+
ivXmHeL2JCpkMfTAZ1xFnC0bxd2ePOJhfrygE2c9iIHAbLXbY/9DarTMATNPqjVCms5RLvtSrHZn
wBUvXnz7wLYnmXfHU8CRezlBK29awgeEAi+MRiZLb7Sf6coDLo5hWjDwwc/ZWP6t4zykVNnIQ9I6
qviiyISy3mYaN9iV60kdxg5gXUVHYJnyBHeVw3eSoIJ7Xhbrm8JaulQDRZ8ArP3FbP4AGp7TKTYi
d/Paz9i6i6C1A2xf9e2cnW5dm1hcrQBBqcmJl/3gp2NZ43/ThvhcO3Qh/W7BMzKiyErpPT1an80R
LFQ0BYdi3tXrG2QYYDiQ9fYzkwOQNdENn0Xlp/6ApRDfWZK3XFcJRxD860AZ/x1dEK3g3m67v9S3
9+2QA4Fa7MKTR0qrh+cN+KckRSsp11wjno/ITxtkHm2zWoJNw78vb8nivQEdr808hijG3ViyaR2r
8AZbBhlYbI+Jf0M/UP8IgDOFW3Bb8ThNqnLSlZqJ0BZhXLsnsTFut12z6KH9GkOEbjSa0nUarYb0
pYPbkyinUqKYXB7UX3WrBZLQ719QwK3QofT+k1gDghDDSA3W2SuenabpIK0GakxtohK2jSj+u0ce
VIJVTMk6km90gF7tr6aszTvBicYVVc4dZJiunUqz502g1cTFByCXcbUTqGNHXPAYKwjO/5I1j00Z
FRjVH5r0i4yFo+xf9x3V4dV5dvklnBBGzyctK4pEF99tlglOIvK20bgJEp677pPhmhF1l6CD9jeC
IX2YW5tcZxg82VTGCCzvRXstT8qxW+yuKvkb9iRTYjlgeUHl/La3ta0GYLeuLMQAEqWuxWVhx+p7
cU+/D9QQdyUEezqWccb5qTvnu5hk5E2wb4Ha9kIsiaGS6kIoiUSnRV5me+XdfF/mnJINXrtkPiQy
579mG7jWTGwPU4LTtn8MUqVdFIFroE1NeL+4jcVhWLcwvw8ScITDayTSra1LDdSpV9jDSAP5rSCV
7XezM0ex4K1tGdaaQEjK20i42zr4iZA2HeqZYI51akDSCpYzkrQ2zXGC01Y3ewrwDMaixPBzdPLO
67yuxT7rWL36sBPn7UGZUNgVmLLPwi/F73QeqNXSa8bpjQ6TvVMnVEz3scJbDCodF/TxCQLH3MIN
powNQGWSur59W3p2km1OzJfamDAsxuGezEnd7TaQ6rwM6i8kPloTXA5jTWSdIosGd+ffDey5+7Xn
YhihPUnIISy+eZl8lFGbtnI51tlUjf+dY9u+vl9dj+ZZK9kxgXWW+UxcgGDwE85TAxju+CTXRzwM
00L8nYn3F4I6Exm5lLY86cJAkDd1WguYR2poYZTxWHBW/TeDpBMIBGcTNReOb4/JC3Adffbco2Hu
H8MsLCB0DO1jlJvWQ2kQwZGXduciamReWbw1U9E3HLrSBcuVN74H5+0dfToY7kLikpHiTrXrQlXO
nDwezCzOIeWXLxTTYgqTJh08kGTseVjDbMrpi5G7H8NAb0yELV1RbhYeZ5P0AbsuvAC0Lx+CZVyw
gd9MLmeXHv629xUqOMTjLtrioyEMjXwnpNtQ8b6KArwG2hcL5Ibscd+MW/eEVdT7rMQI0Ojg3xyc
GE12ABBRImDwr+pTR2u7xS2lH4VU3pdQYxdSoN/rBm61M5MLwgrO7ak6GiK3Gs9rxrm2i5LO6nxO
KuUbrfztVjqLKGJZlcyzHV1o917+o7aOxV8tsTIDeToJQsciqwbIr0fVQxpY4tom/Yi70VL4Pabg
YNoj20thPJy9dA2qtPk1jFqyXF6qICyT5fxdYxGAVGxfuP0jSpyqa5JYgFGDVXCOwXBTnRWNbYZV
uEpXLc1OyqStB2DzzS26+l6qTxgmoBKOjnjWfb353E/eprvjjBy1+IMIZDTpDI4ySYhlsMJj2e4n
KOBw/tmMnKsRPi/HnZLr/EQKZDkI1MxWFallyKjCpqAtJxzVXzW5QJryrcGVn5BTeBKnadUVbqYB
4lZibfbioG6g0HSS8UTuauEUwgiO0dBEpKNT2W0fqMuZBulotAkGiRSSU9isXpr2cjGOzehbJMIX
1OZ8HjefIlsJXG6IvO1GbgD/vawc7gVzHPSdG772dhlTyfm4ksfOMxD9STnHl9O1l5VdxctNYjeq
U0Y28XlwitCa34aqa0gnCbcSQUF+drTG/6y8juC9K0UHpM139b6ApVSYSwrQQtGsC+JM8wWMD7Eu
+YkbJWiXALmVNMBZ2v2dqz60l7hUD+An47gwo063sektGht1Nl4lac5kShx5YDHZqQQMnVHygXCz
Kva+nICzJR7Ef1dS4yEnIHCsa2mfCqloWW8twjxsjdDgimg8o12OfV/16U+k95qqHhoarzjVSv29
v3TGDQZq9tK/Rv6iKmG1TFovublEGx2g0Nu4VA+NuaAdVLCh/CnSBNbTNY5UcdctxBlpjs+JgFur
YiFbRp3XfalBPBNaCxK2MXyvwhpyvRwhJG9aiHa0459t5DMRZKcW+bNTIhFDYsdVTve92mqK0cGX
kyNGyOXfuzx5QDHIhlyRFEbSTJFxPMfnjOXUY53WptAfDs8tiuJsicqqSYE2qXAhSV/a9eaorLjz
lKxgb9RlIV/bpNwqoJ8ju7i6k+5wPYiFwmrq3tFayLS6uu9k0H/tYdvCyEYDm6Fo0YcWlC+wIAkq
OI8ymnawzha6vNdLxyhhs8p2wf4TFXHpnoNuNnZSK35nWWzJNLtttlb91vuE3rYc+4yZBNO21euk
OQ7XCp6IfYfaT6PtZa711cqPdMZyWO6Qa8iHsuJ0f3HQXFnHlI6ioArwgUCa9PrmtVU47YOYJUuE
saLWLFMlrjKb5ASjB/eeJ4p3P3lRw0sfDqI8Gb5JZn9AyT+digJpYegKAo58qp6eBYCwVpoqBSUb
SkV5qyB9Kko5nnhs0ypmvuIXRluzQVxvsqSoE6XU4ixtP/h/zS9CK7sjcVeEJXzabwKN4b9Au5VN
ZEP0tglGMYQYb1p+vKgzzPCRiiAp8geI1lAhu0u3JmVDMtg7YsF8k7DV3/xAsRRTcor/GUUd2uj5
PyPY8LStOGo2FvKKpsrVceVftAVKNpoZl9/pRQIAOEcqOzYeS8LeWJH8bpEXEIi9bj1IyjSZgWvD
7elj9A01CJuv8sxRzAFVpMKVz4CjYUQDtG6Y5I1aQMFYlMwzB0CpOHCQqSQgenPu0srR+jIcJDOg
bEtBYZ8kbTylYepXB7xKZcBBCXJveKdn4ofEGOZCGRZyGcvq54aA61C/E/Ch4N4UKRsb0n+vIEfg
SLiltjzueAhgO99PyJDUQU/AqIz36q6M+U5ZA+YPa7sL3zMWaHBMQLc8nUj2lfgxQqUI6PyHUGpI
p2FREr0IvbGbdZCti0SqNRcbSbPjOlsaPrSGb8a4l9qbYErOG5bAqtIJ+P+UoD04rg2MT5SNn/QT
FfHkbU4uGUGManx2KJ9RTnBDx4gVl2YQPm/7ZKHzuT2Fxk1HUb6npZyxoy8teguDzC2d6ufxTV6M
ZP/5Yt8bdzX26fXHv6I3UDldbLJjnRbh0BTEP4mikZgTLKaZ+foN4AmLYoqYCiu9TRkJi+zUoK7T
nkwHF71vi5JKEEzMv7yVLSeH5b97qUM/jSNdyKM/BjYaX2fh9HquQ5GTKtwR03OcdxW4AC3wjXvk
b3iRZl6kbVthTh/dIiZpizVa/55OFAMsAUJOJV8rBAw7EwwMkbQkYvxvwybXYy2JsSEDNx2Dy4OH
1aKDNhh0vcgP314J3NLE49yK3znmgNClVOkihGZc+DE9EUL9MjUGHcJOKYOraHIfC4XNJh32+udt
GvFguVGIBetwgd8kGl0M1sZFAN3Af9QoR80+4Wx36ql/uyk8p2e2+SKD3BOGivoLROc5tOUWN7Qk
8IrgNE9GSt1EwzQEmhPPL5n+StoCOa0ixLJLrzumQz087zkryabmX0/jVAoapKgAFg9iuxfeNLqI
gbyWktK7v9zYH+i3Ae4D/VBYffy4QJi1Nxfl7Wekw/wK/5UD7ic/gb9HHs3BFNaW1R2R57QZMhI+
bZpo6qHP3GGC4NMg+W7XBbA7tHKmRF9F/5r+0kxGGxCJBin383AysA0RU0loTqDQzuZy8r3ZKdTC
lfNNpyKeCuez8VX0kTgtMmlsDNFc+UT19W3j3kjagAZuJhPi00xSqJrlB2TuvTxDCWgPeOH0HLuT
GoBtI2gKn5tXg+y5HJoOUeIvCg1TsRzxhCHKouQPrDrxySDV++M+GvU/FVVOL2Yd4KE97Kzil7Hq
f/IAVc8gbebme6sFkZuSwoaKw1Uw/w+2RY2brODzuQ2NFuhYI7StJ3bXRpiWEyN3H9Hl6+yzgJkx
D29/RObf6TO1LA+5I4SR/BbjbueF1u8JljHgH4tMTE8qpU3HKV0qF0+YiTxVGNr1n9a52eFMD70E
CF7/7NYvJ7RM6aMUlQqQ1ja54YMfQ+chhRTSC1TL04FrJ7PDhLvMpSkdTRDoy2RZM9naWvSkGzhs
E5x4V6UqKuN6YjoRXKqYrMFNQLIn93G7oWoedoiYGBn7+X0Sn1y+euMuvvZ1DEnG5hBejRCCiGNV
p02tPpB0dKtTVU+bjIZNqTGF7R+KY/P7XStza0WQ0mYyWglsS7GrmYVgr/XxiNwKBlpiiewuJeLm
/PCLZyDcvz0WcucRgD5zmIL1wRADTKeeJ3sFy30pA4uR2Bef85itNGlLKmC6xhuX4E/P/kUs6F0l
7weJgeTSLwSGfPCZz9Fb8tAWR4CMN8UEqooi4Ue2E6ly80xQplWScUEwWGvt+H/La4k9kHSKhxuO
ft5xuGfnTf/7I0POcN0PIl49IQQy5oAFs2sk10Izs7HMtuwu7Rxr33efO3yTYEGnFXX0nhsjqnVm
aRJWH/rSQYgu+fZq8swGczxGFGxaI2GInCoXh5B5TyA3E7aVXgaoD/K36CjryUtKiuBJilpbbbhJ
rtcFl4FB+SVozXLbxaRKOTMgkAILQ/PSTat+lHgm6sXJ2qcc/GM5C04LdoOKn+xfZnPpi28cHA/R
jFdsXX4P/8qyY79s9EBFRGCjIMfdtqnCkYMOTLy/VWQaPVMqsTH76gx/FsIf3puuKzsDYz0ytQsL
0zF5Ny9wnQ6WlIl3CNbrgyryR780jGeK5WKs2HO7n5Ja59If4vXF/npuZ1V0NDC7yzQ+Qd48H5mH
qN6kMXDe82GwcrPtBQTGm1E0UV0TGASEoFAVdsMj+JXM7TlyMZr0Q7nL1VV1M6NfoSM/TceZ3pPN
2yFQBdvyiyn8P7cIqjk/6cHVBJmNRLWNkb+JAoaJEcagA8BfClu/YV7mxYzmFoK2kRucyhCqR+jU
HQSdnTYVSjBP3dNtQz+pSg1CvP6bfaDS5XH8aLK5fe7v5NaxYqPvTaTN8NnlXV0Kd5oYDg7THgRV
zOJd1IWFFrE+b0MdWUn3ZmaF5WVPaTg0KLKhVFOcDKzGonZ3DC3fXxrJ7FSue0eYXuFDJAlPSDCj
+kmU8Uwwa91JDmdxx8TE4S+D04CAkyOYtcbRhODZwaOlP7bk/wDYAuu47MuT45tesWUnLAjJf+bx
5+EmkYLOSiAj9LmfDZ+40Y1FjZSCuyDf5Xcd2FC7ou853VxApqEDZL8y6O9Sbbh7NBJfkpEjmSnV
4ev4j4bJ3MgjJk3CDDVkQyzQE4Iu7kiDW/2pzR8HT1eIEIfqrasDv9JlMKrLKIpntPLCBMXYDEoM
Q78uzoO2AmrlilFBYJCduX6lByaMSRNWsUnGK6wOMzyPEYjkIbvkalcF2xxZDvxK9JbMLPZoQomv
q3h7d7p1rqGy3PwXCqONCKZxbryq1xAm4vbfjoaHFYrSU07k9YGCRDJSUL6NO/GKLtdWXHBWtd03
vGz05aQjhiA3YKVbu319ZKrlbd4vpm+g66I86hg+qaF8Ob5pMOBSpfxiVwey2g8INmA9GUVr1E7i
T0IEU/hbQgyTqiLciNgLYkERHcM7qjmpi+DxJsGlEs//xUtuujHOVoqBQRf0Penn96Qh5yYPG3pJ
H2IkfKM9jjabtr3InngEHrjeVLwuiFuwwP+x3RaGi/RWXiMVFl9vYjdQntmhlyOv74rr0r3aruQc
bjTRoSImkha+VD+64hMv0p5jmCl/vm88xsuultU2WyaOaSiAW+UmvJfea7FjysQNdHAQeUm8FE4S
enygHyKeEfty3olWvNP1/zUi8Fi+L7RnlJyGU8gRYr2OkpwuFjqkuPn0ACHYIbCN0kGvIYBsgGse
udwxIF4F8jZlow9PgHiQqL9F+hNm7ZR2GYW3GxNaAJAJy0hgVri5nOg8CQxj0wuzwWTk1gpVK5vo
w30PI5AnexYfrzMOS7vrbS6pmnFU6/kZ+ESztCx/ayNDjTzIDoi8QbXDkdjwUaAWFt6b/hv2d9yd
l0heTd4gJdUfFk9mHkDH7hC3jcvzNucT/2PGPgv5hzZKkN0BQCENP+dbzVKL1tQgEBO7GfHOONu7
NkTzFotkqIJwyJ6o7J55pOHsZdJc0AWcksVR+rA1Mh8U53B5BU4a51nufmop1NfWMu77HjTz6xNK
0NUDxZ/kXNNfMp44owIG794JQGoAU09YKtXHC+myt2wJyzVCHoohLU87xbojc3hEmmKfKTCEtzVB
7Ocagt/CBkKS7aP4MAiq6ibku9gIgXuz3QP86ruU5t65H3fZ6L5dkv3Yk0JzeFL4zy2RhvACpagR
DFqQQC4042ocSDEJOEVaiSwcZqPCBuJsRTxlmLTkR/xsiVyCe+UvR3HSn9RUMWQNaKiwuiPCxDGI
iPCdsMyTL9Xp3CNvUK3kRDo3XSmPrafp7jwM+tkJOkZd1RCVdVjH0Kyj2OmPIDL0ASLIrgMhlDa1
gMTMjQTFEvhcXF7Oc93XLjps6wv1OE7E+5yXQnh5GBqOAlmsGbi/ANwnuR+N5ABGU8I8Jg+HlB8t
hU2blL8/PvfUv57NbnDsKaHSh058UMYuntMp5f4X/1CBoFMSYsAJHSfvGJHY0L/6ILPifmQfpfAl
DXz8YfCWNwDEcoFFo9iyH1cX+AuFgkqVATNyFGvZAuShUnX8mRh1RUQUMMLMIcyeXxWhkGSZJ1yQ
Z/ss3Ro+Pc1CT1yf4pyS9/PRkgfG8povioOhv6MLXW0HQiKwO/h8NJwCBQyOHKVdKoF2r9NIBNqN
j11E8pjUB0vvzXozDi1N2iaSgEQxhIDmvKwC1fFfgbaupB9/QCzGOf2DzX2qAs3KpVgxkc0oyTVl
VilInqFS9Whwz4eT1xWOIWuskAE2EWELcf6WsjhmFCYLTYduJf8R7uhHSU55ykfXsNPfoqJR5v81
l80E/FMn0sgWQ2wBZ1TbB4eHzINPxg5By2JIY16uzbDmJGgF9GZF7v4w9JGZig0hEEfL2qJ4NhdU
b98ow497CYQksO6Dr/ZEYpdMlSywlhUdR0VaEhxQ47JpnrhrCM8xg7S61spzke/gsT4jGZdylvOa
StbkhTu4kC2sssO644LZKSjaU0NEf20n3Jeh5iyOYTci6dYB4rlnKez3hzLBkJcd4AfIlz3G2fwV
0EDpX1dRHZMSH9xB3IZF4vZ0LNJVkdOZER4rMT6jgXwZ2vSktOH9/iz8CJbfERhVHXqhrE3K7CIs
KL835U5PeyF1VCSX0Z8FJjZoah/c3gcJTOASq11Ucgxx+84AmgWcVzyZ6ZKDpASjF1fMRKwuATI8
2gdLMJAVDHqMFDwWTziaGzjtQyVWRJ3uuMSAb7G88j5NwkNKBbvcHb6Mo1kghndc9EKjKlLZoimR
f2fP4pwGyXtCkUhxGPx0ulD3f/1xIqzkfYaizhnAXKEhp6ZgVnzGacXPsKuoPlF8UbCL7c2emeQB
dax2rscXgQ1hRPcksx5+gL6cuVWUZPA8NE4teCN7bPbCLp7D1NJF7QnVJ2mjFs9zWRouGDZYGF7r
bP48XD3ks/7/cgFWzoe17wx+dlHc24PZ4ijdjJGe47vduu0VwfthDQzsyECr/bslWEEUw10NjlRh
wuiME6jRYl6YBLc9ykZPSO5VG048MJQhMrKcdMa2yO2YetMsq7ZYe9PiGnqJOGCU60WYGiO2xH/c
U9q+UyP/XmG6yQCtQ0chhWHo8Q5Bfzqgpd8BsQEQMWtiEQcHyklzkPT0/sZJNIgAaQSd8gAIiKJ2
sGInuAHo+cVIkKktgfD1MiCvjJpYedT2tuAJN0znBOtiRDytIK4rsQlQvrhmv7B2hLK1nhgak30V
gBm58ijyWPBGIS3QoMUttI6m73xFrviuBZv4IR6iPxQjjq2a9xJdpx9A3nvz0Qhr74BqpnzVLkze
K+ME0WqIflDO0jTmduHC/SKuDzT9gEmBnFJIifMJHVNxlxJkl0vxgcl0Sal7inFk4p/kA/vGgv8/
OcgKvtaKKgOjp9sGfaGxKJJP+RbCwVF9hhxMmm4v8OXuoA4Pv/5saO2NOV03QIT5Y2MIH7M654X6
SqNi3Vpy4ghsbLp9ECbWh5s3zzz0ODWVZO//7QsCuV4kpnRwZrzNejAV7EyUx4pPyyF7rx5vjhUH
6c+SjPqJ8cq2eSQfOP1FQDPVQW/Vxhb4zFjLDXxYgYH24J5J2YtpN14XvVbdC5AnMNMGoOOkspgI
2UojJR4L1gWGyjsbDbmJ3FyE5HMtV8JDab4IpCpmTNUayPqv0Lwu/azKqDhCA4efnVNzi2Q127F0
lh4+XMVosDjh9xPHESqOmVHbJIeEZ6wkvEpbHOM7ATkv56TyhkYnrVi+zE/WWOoDQS2JckTkV176
5YfZ0R1wAiUcnpAZrDZ6VldndFuf3aGajyeW0J8gNCaaGTjTiKGEJeH1linVcS8ODgNxub+QmrsJ
awtYJoP099VBxjAx3vJo5B8wOy3utY5esykwsZ397WHi+UZ+/Pg7bafPMK7H8qh0yM+CFMIOZZ9L
9bkGQDO1sca34Ay2/c67PxZQgSJKru+H34ISgkwaq0txyIZus/ygRAzUFoYRXfRIVKN/dJ/YRNMf
JAD/+U/a5W6rdVYaN4F6AecaTokyHczU5jTWO/BX36gBefcVXrPaVn7EcVWO5t/Fdcda4bCfbDYr
8O4/TnQHZIQ8UJkIPIwYF49tUzs4dPJGafOqcEuWwZnm+3wwf8d9tvsQkC5wYBCq0Jwo/zjNWvpt
tgM7WosPdWwSEzGHzto1wea9A6I65YN8Mbz8Jv/4NMMRGhP0Z5RlYdyHuWV62t2f/ZMJSbWKMnTN
cM98af+AGgBaRHHVE234vdPdCykkE+olE6sVqU4PiotCbiuSLmUdcu49qoN+hzuIc4yc6ZUqmoMA
ys/BdcDeFnEgP+4XfNwWsJCufieiha9iFZkJbybbAKTGonBp559odNLgB9YWhW6dQpG9+GVzZyJ2
IgiSqxcFsf/fqEjxqUD5Onl9RbJVKIZOwtSA2JX4JENofKLNjYbIz3QxKRiyBIrivzmbGk6IO7dC
Jy2zCbChr4BPC3AloxLrGBOXqcfMDPbgSGTmeqlQCqXRoeYJhCPansSCGD46codIl/np0B6NTmjo
+hUHpZAXIXLp9A3HO6gfhpq2fMl/2OlIFrjnxPsUcXCPb9jP4VCtmpIxtPaK/Q5FpuFJPLH1PcHp
eaifpOw4YUANhzIzYHJibmlOxntqrtA29gdVmzB5mPZ9Lc89VCc3QHVedZOnI8HD/zpKxvPpiERr
YAurL5tV2hWlwAxWcl7Jr6DuROAhLMJsE+rwWXdKjzPgtdQjmvFxs/8nWk+09K1g3s2VHokEox8J
Wla3krcR9mQbiYY4MHXYAPNnlpLHO2hrf23B6hpFlB//2HcapQdqw4CSgBSpSmewFsQAPqfoNBQ6
OpXCgNDgdjtKz1t8Z+J3Ujq5TrdVLLszvXeuKi41LfV9TdZl1wBoljjfgCHKdFez0OxewFjGoQcN
78nhfbMqSUYw1wRVFpfnl6rk3OpHiph0XU/5I1lYQQyS4g9lATRtDcPwDYgPQIxruQfP1LDAfERW
L9Rcnva4DshQ0FVAtJcvba3cZ06rI2dkEIMJsTaCfpkmaQBsbgbI203N4osgwwuGdQRqR0SibbXw
DH49twmDgEYVCoSTd/S2usJoTSbcZvmTBKD5pVRKHjTnEn/FIBeGJHtIl19xjdSOXKxWtImfJn9l
UNa8oG/fQeevJF3fWjXNxONHsrmUeeJOnHRCnkC7Dzjzjn6I456Gy/XAJNiCQ76F17EQjhUoMlb8
V2z40xIUbDnzgUbEdYG0qI9yYzrI2k65vAKzsNOj5iMN71vT281UvEv7CRzCXBs15V37u41vxbvm
41dTEyRPhsqKHjuHiPnBLaLaWQFsD+OynN9iF5TLlaYGlrPIoHO9SYOA0bu3e315ffKLqo3L8DNx
P1X6S/sC1PUE5byfWoYvgPRGhez8Ah7QT4JK6clfYsmtuYuRaXiAsN8Rc/PjCYtnhXsbbRuJwNmv
Og2CBbVeBwhM/978jNkXFrTlqhSVEVvX8EFlH6V1fBry2BM2dvMZ7n2WF9BNWbVXKOUAtsKOXUXF
Tx3lzPeQY9reBrAnlKwk9/XtY197Ao9lcDskS8zB3RDWs3ZvVyjqcpvElj44KifeHuRvnd9HRA6H
FzkHiMLkRzNRMWiJBDJLovtWpMcgNBJR0ctpMRwFqZioDQuRtLQ2kFuZ4xN/Sh+7GM9ZMDHCN84a
p1+Bbo9aM5bi5l9YOhppffNDwoTimi178z96JNO4RLj6uWt7uuZ9fZ3GYCkqeAGRvNBtG+K1dbeF
E4XeDG2TPnuLTaQFr/1LhlIx4X7WcZjOUUYoG4kLlvxzuoWTCbuzJ7ICOuNXNtX6YARtuJNbEpBq
7lWCeKS5NeqD4/rAsoAMkPe7ccuDwZQpjkyAc8E4F9+nDkIrzEZoUdBU6Yfnk8NtBBSpb2BXsniI
B++bdG8WoOZO6GjA7gJhY9HOQiBgAx9XpuHywrYdqYtbYLnsXmbq9zD8zGiWuGOGm2B9AeYboLHs
1J0HGsB3r8FQiAl211/0P7TjO/OGNKbOJFrTCpE+vnulnGHUGn48hKNQ7hWgHxiqT6VKDhYY0pQZ
GBd7GD3oVobNNyUW7/c2RlrcxWK8YxO+47kNZZkvgM2EFI+R/MC6/T1KZpPwGrRI61kQ2rQydo9E
GqPb5oHljbJaev0iGidcz+d9cMDD7yvBimbVYQR1PIhzmSM6VDhKwgiUwNHNFHO3gev0ElptlUgx
8dpvRYelmItw2k2kBvCwd5c2jxAaXpzesTDMQoG1ix+5HzjcikNO06urw29rYTFE+ro69OMjFQOx
xU8pqfOGGgo33EvXqRpXaCuTBiWOzJ1RnEQs298jSGBMNDzqmJamtdybD43GEujiJy+CSdF3/U0S
sMTEqI0lR2St7EHhm4+2VH8QvgntkpezuFYRaybjf+WLFVul9bgWV6aUUZjB3b4uALH5EtEVpJn1
qxr58iqOqRGvr3ZjovEcwlHE5OwbOEmFTit5e1ZMD30rrJBmLlhOaQqO4xeuo9/ZBfc4Wi6nV2i3
/C1RNnRRQoFeFCaCzT1PATBIcNbbhuHkJTsPUgQ33QI4pgNrRa80aPPLb+Qahm/ws9Xhuf25IPdJ
wn6huosPLf0iulp4uekPJBYSLD69DXpfW6CgPKkPLrn6LkfK39ebKC5u4SFHYyUhE8e7u4T8B+97
9yKTaj+e/uNQKNuGeOvcSgk/avCSb0tE7wcB2nLYmblY0Nkgjat1fHirPNnH6dXK2E+WTk1ViG/X
i6tkEAXFYpn1Dc06edq43vqePmIaVXEICE6bPywkezBZY819wbzcGUXl9LsyWwJh7blsQkym2pa1
AWheOZR7ddyKx3FaEeYa7WGGEDBHvOfNOBfDNQhlx84GQvbaYUzS6n0W6ejJ7J9nuqB8KrIH/pJq
FUQHdZnxs04UFUh/HHoXzN4I5Z+vggElZ3L6aRwF+z2WaW7JAF0R9T5byQLeZoTfw2q3JxTQdWWh
bxauP1A6waQE5VQT+eGSrjfjLhmIzvZrmmnrmrbzcOTtTb4NiKdN/08bqrr6zBWAxr1MRXiYTut0
E+6E0Mtvwsq9HUAb/UvOTkpceol34ib5UUIw3U3ruM5C6Bv5v5P2ZxQAEj2jEyilfBYM1bimXL1S
j8A9e4YVTMiu6da9w5/cc23n/2nm/H1eRzslAeCwzKPmxpcu0A2nlV3oe+xjZsewx3Z6oMQ8PxUR
EHb6I31wuoshVP6zquX+W62WyHj2CNgH3FrdqyHyYWRjrMkW2+AhFgrBlBZiY5BkusLPGM2i3JkN
Jpgma1+a95cBr8cephUv5JhYBUNI8y7elOb/pDKBFXjzpx9xRRVKCV95SGxEYNmofdQwj6GEy5Ug
6EpNV13NU0DD2sAPYM6dVYR0WYM29tKTiIiZn82NnEhEs2LOiB5qYZ1wc9GYVRDKeaIVSMbPgco7
+g2PvNIqTPMRKqYRDZmsNXr42QF2JSvxRDI6Bj/qKpZZh45yLRX3eItlQ0QiiAJGJcJAKR/6R4Rq
WCI/EiEUuSocvKkTuYm8L9kPcRE0QCJdwm3pn8zKmiJIlJSDiuKKvnE4J8ckV078YXDBigF58xFn
m+nM56zlhs70BoXBYsphry0QBPv8fwKOHDb1rxGeNwbG+hQHPFbjPsByqJnBT1F0cJBRSbCp1VfB
zy/vjaWXM317Q8u6eETJZx+h97014NWlMmOhNQpiXjZXlTIO/94dj2bjl+bD1CdIFr92mSO/Px8y
a6nnxjhjPgwKIDKHEPhHNrpvROVB+fy1ao5QCbYnoEnqLTkmdQCLMCFY4th7M43n1KK6jSNCO5nB
j0EnyoTa0LPi0HEiRuWF/3d6yDypmOSwQ91itRpqBeDtO+Zgv8mm19O7EWo+cSPo5DlRZLKPv7Hm
lg7pOCStO4EGI9LV6GzvcpL5HmcQpJVweisNZK3Y833/o4PME0RjF2Q56WaiQ5ti31N65O3l6axv
Ht72wP4faNlMLHqTkPMywURGY+VYUm5R3PZkv+hdM7RMvi4LA8R5H/i+6AvU3bbSXBUCMxagr3Aq
3a5ZvYU5Zmy0ofB7dT5B8VbtLzkueOAQqfO49Wo+KwVwgQziCiktr96mekyqKwANBNxE6W4ZAs86
JdzlWIvnnLrc7OOSrMd8h27xzB93MP8kb/nYDRRob9GLSpZ0bUNI5oqc8sfkfBr1nkRBeArJi2g0
f6zHbuhJlmbmhl6/4bIZSsF65s8W6PwuLv6W8JklGsU/Tt+tiqtaMTcvqBxNj1SrSstqJdphd6Bl
VIiCMy1ke0LjdnLx+CiBCkz1YMBn/dka/dU6k1NigN6XIch5d1HBa0tPg56m6YlkI1TaauD8TGa4
0/S8DWw6X2YuYaNvEdmQnzV/6iJhyZmK2l33wUFOdkHGYJMeDZjOnND/Ajex/NJNBjrh2ySQd/8m
mmZsoUgQXtSHpd/VrhWUyxTV86IgtUgcWASpRkgNp8AUxx4qPg66PjQrSVAaCuxhwYUZaw4jOcya
Ly5/xSwtcKx2Y6X68oXJFJv+KcgiLuS8XSXkA4zHd//bVNKxxCw8IqHgXW/MaQhTJ0LBwStDbwm2
+YZdP7+9qD2s7W1LElloQKnGesstOb07nStw9Suk0zu5QcGdMzLbvSWYa2/F1p4g7Nm1rwYqe8E9
tHwxb6wnuOC56Gc9MZZpOshqfYHZPaP/9TdNd6WTCglJ4kwvxnOMP18TZqZNPSPV+LIVaDkQ6m8m
o5ZimQmiLqurdRRHdMdpl+cBc9SY/EgBzFAZYbbNLS6+PONizitjVg2e+/yTKfEiQjH907KZmqtQ
cw44txCPQSDeLGJUIHXvEBluwA5bEaZwnRrv5/s78DD7Bkv6ZJdUfPtsCPZSDYliXucH2lNxH0LD
1RD7uSuDA9/8T9tbSXBUjKE1zkAJErfKKqThlUWKd+UGNNGIrWX5bsy7GUBm8PvNYLnO5bk8Cvk4
a6MkhLNhq4VgC+9Rw84C30w2OiBAgG+7RpKM/pJCm8VzgHjTInihAomXSwyIsd4gkhMtwjgoKn7Y
ARf7irEls2kB446g1s7fKu9J8Bw3DeKWsxFpnolM4HqVIdId2mdsfFEItVyYNhglzYhZKM2MfKph
cTKMIJp6FRPfN1qLcrgPcbcp9gOKbL1hNiSGj9mWSSXQp/1/5ERhaGPV645xclGodCk8vMYxzbVa
0MIptXX9xv8os6arsi3UD8mT/jO52IvdD10dONdmiog/Z0Mn4r5wUm2T/ORseZ+t/6yT7tFE+II5
uWTKUfLoV2UeGI8ErLFjW0heA14irjNpClCHg8kzW40Ny3RlHyTmTWCO/yi+xs7Lg/ot8+h/FBt4
MaIvv/Xvd1FHfHK7HQJ+CAcbq5YVdu0iV1VDV2iPFXN1o4SbrOgQvTTpspt+d+5rtzND9J5lYZ9X
GnKHp/uosf8niZVKxVpFoXwCAVMrC8trd4NRWfeppiXpaCGMuC4K6yUbiQSXLLzV9xSTbnkVStjm
dgBhek+8n5dUrMIkObjUNyKwI6WvaOKMlD3TpUcebeLfvogPOFt3WZQ6ys9O0SdxTdannabC2VpZ
xR1gFE7rcPGaRde5jnkwiwifhKVvwyK4eK6u20Ba8CNps6PMMtvo7Ym7c5NeqcaTEk3Io7fQFmEC
YQQFli3eY+RKSSU3kRVthXv3hk8M1mW5dQMxD7l61OP8HrdHUzptg+wjmQ3vKCIfTMf6Es9W/QBc
U1RKvdZby8Wz2OyQP3uQbsQNcJa11bi3BC/1vQXpE/1PBRYLxEutaMQ2weCw4jjWSf0GLRQOCBto
1lC5VqHYJ+SvXDYMISAe2320jJFHpWVHyqBd/bScmbGk6orsMNJr8VTKVmciW1H3ctXiYoHtrma0
sJ3RyvnF3f+K6FarWmXk9LrTC64cCxARR3NVyNl6BQhqDWOoFGgcQ9nYA9EREE8Dg2vMPNaXoUAa
i6R6VDNn48q7uhYoTNKILVaNpEbYFKHNz1d9tOWDpboqUXe6TcvpXMm16ZqUfI9zW/Z14Tx7V+L4
mgG1PSPVL2gqdjYMosdGa6s9syyKUQ8g+vmxxF1d2T3WbIVyxzUqmrnmgfyhMNHI0tR45oJ9fjFN
qUw8V28+JQ2OmIRk2obpbiJwSoHpEO94jZT6KUfnsgB61JmrddAI5wbDdGP/D9prkJzLxwxbO8F1
U9+lN97SHvSlgE94+BHnVENUUqSJP0dimamqmq1187Zl5Jrah6Vp8Lal4rQ8WAgmcsFBeH4jUOxT
3WHouCJ5soRoKg3EScCXYeOF/G7cxkkMddVTkdNbHexQVhnnHyyAtZcyNuxmzOY3K6affRKL9YlE
bwo7jsb1pOOQi8k86wzGfOGsv+VIYGJm2WZo2Z48mioH5M/BH/pn1rBvnqDoq/VCNP2zhVyCLmQb
Sx2tgCdyRGABAEAPtJf2teU1xIBNglUTuj3K4AUkVZvNxFC+4l7WMuNpoX/6Oz1DaNf/Km8mnS+M
ibyn2Bxa8INcrtfefDwleBdf9fJBjzqaOyMRiG7vslEh55/Lk5zDUmZRi2/IAoXEuyY9JB/ZwXhl
EntPUWJ//PdfpmFX8jbaf2XKINRn9/RxznwftBfJRpZiM+U+jB584OUtisIkmquZhmFF3RehUehn
gX8YTrxSK8Fu1PmB+9eyJ2nr1uix0EN0zihC47QeQ3jryG1j1kercX3NajSIIX/VfizsQ9j5lrNk
LndaWBOqZ0m3fxnsCKbQp1uwuIR31Df4Mqbss4JEAInlCHboPudRQzrPmAX9ilx0ndBZz7E7nDVt
ImoVty6uvz+mCg2HHXmqErC6ilxE5dLc16DRO0SJiOpdegIMYRyvidwsjyNd2eq913L8PIWVOHrS
lmN9DAxcX6cHBenuSzUv2BLIkB15Gy1gQMKCOIUfbEmsYNSJrnv/tLgkFrQXIKdW4rtZPR3vkBWa
Cc9v/fV9KaMxbHqGR0RyjeLqceslN1Jb1Al7MYWtI3QFoRS3Q/iDToPOX6ZyvFooJ4PKdyVJ/69m
fvH6YmicSSqwqrYAO3GKL1SHbb4WWKHq9BwO15Wfo/3RmpIoH4CG28HV9KNEV3gdz/SuqL6AVeS2
Vt7gEgaudd3aI97Torp9gohIX7oJKXmx2V78rjXq40b9B/OD8o68MI3RlEW/P7JSvOl3a+Uo//WX
XwchYwZHtM4ED8Vopj/pAu2zBrFm3Dult1eVQ8RoNIm2AcUFNucPfyed1LMJkTHUwRLBqEpMF/Ia
MrChOEMVDIVeUaoXJOPcXCwTh5S+GKNj86aFLGv+KYPP5li8LgvM98Kau11yazZlbdMMDijUH9di
DWpyIm2n0+85R03gr7KKd1/ijCadQyhzo2sk9xgDD6mhMWtNof8vKDWuYnMTYFiHl75uA/bqXw1U
i/+1XuPfs4+hb+nOwboFIMKvhI9ZSu3iqSsCm66aYvDBBAxc5huOe756g9AlWtn3dLwtp8ltbCEH
RxVEuGEkppZ7vS2Bzu6TejvEMVe61Q1qsnOUbVRqn+CpgCsVbI5OPNuSpUkBS4b3p87RlfoOGiZ7
zsXVD+nCJ/ch7JXgR2ZH5RG4YI9obh0Qg3sRRgkAGpa7k5fAznO6ZlcLT/3cPLGfO/1Nb1zgE2Pv
ak2WeodOvDTQh1t9DDLAgPJy7dAxECVXoh7607r+wzOWiwhKuF5DOU7g0IowXi1gg4XsHn90ogut
TFh+nu8Pyb27H9cby5sFWNo0JYS6UiT7WlA9cZUBG6dy9Jbx+Fb+dkj83giFFgt/HZexe/eIkigI
TNW9KhiVBMdX+sgUxCdA7cunU0B+fYqYwe0Skl//FPhcFFkjGV6mZ+vVPEbbcjjEpmpuHRg+wrVu
p7v6WFzo/V/BV6STWpQfUwTXHtvIMYoD8ekwO1P8rcoHqSvfX9Nu5WPWaF7ylagQyjdHzUNQicne
KIMgiYVXUsKX9a9TQwgyUEMuOBL+0FfgK3bcdbHj+8FzJhgksJvlbchIJUcq7KZCnsWDJ97xqtD0
ukNGYeJEwoYOVBBDbPuhiWWVIJTPMQfXwX2VFGRB1W/zOs2vGdiBVgMbgCecv/cX9lnI2vTCG2x2
UfhNcxvHz5aH4V9814hjuU3YAsnstMn1lRkohz4KLv6AbT3GlGkp6nwpQDzfX6UBnCWw51AN7k4H
NvvnNkihIq6HVImviYO0SkWkzt31yj2SiVrEP6vAaBjpSHmiHTvkcp2jWEdGuGS4f2rhYtuATccu
fCdrN7y2PcjbeSQPGVIS0Sy5JnOWmiNTaAzw5U9ZRqk6ykXkJy2UxTqQlHQ5A2nt5G1fOeCdT0uh
tkzsba9In9dG5n44AYvbv++7kRcrnfuDjZXVdBXDezSUF2Mw/ZNCf1V12f3ICD+Xphgkj+5Lu2Sb
iFeu9QNAwPkSDl6T4rUUs6nv1sMINQ74nBZZDSCUcExunoWHqLcKHy6xzzjnzM1XS+YYdwjQdycB
n2f4x+elsCPd9JXyLyjVjWp9eAzM4GjR6ISq7qPGMKgvMyS/TaNDidaXv7+bhIkXrArMsu7/tLYs
0lAjkiknjiQ5eTEGh4AcMFbgu2yIzLP6iK31efWEnBqGeJV3fWQclU/KkpsxxgjUe06HzuAwsvj+
KUVPOng82flk/ScWlPrMbPPmPPN9BB6yLrFnMY6yd1ZjUYKaxXaw9JiCyWrH5pXTrTc7pYO7SV1A
0M0ANYC2Y9nzbcBxVaEmink3cqvx+oK5UFhAGuaG6HiP2ME9uyHO5DBxWWBv/L4qmtEGope51Eow
aQ9/JkMfS7lqIH0b2u/Nv4amipNudiFxt2lKVCz+bin5flsHfVPs18ZXAfINgAZZDKJxZb3FmiKj
q6yhIiJkMQTfXKxLd73oQlFrtATJgG7jcuvvLG6PpzS1IdjEriEK64WDTcjEfON0Urm9wgAjLAsD
mEzU3a1cs7Oqr7HMltlvdcF7cM4cGkq/bJ0/6U7KxHthnV/MJ4R5isSmY5V6/3ykbFNSdP+aQjlD
Cqbi6DPTvPQRkIgx2IPyDupMuwiMLg+D+FRj97x+DM+cKSd/uNNSU8Ao7QKX01Eut1pkVXCLKBRb
oxG96VRIUc/WCDnagYl540UblhmZUj0yQfS3DVEUnvTRHEBfqSgPooiL3FZfeD8apQml9VynLpBO
QJuh1sry1UeR4Uzo+FAm1GCQeXAm5rby7xCEEogJEpMKS8gTEdnN6+gYwFEKyXmpWFfFSIN8OJ22
ELRJvE357DtgQELtc/nZX+tD2lN7gF72m2vdj4y7j85aC9tiRqmV5228z7Qa107r/3ggRnzVWAJR
txPWclRtIoCb+p4/4sog+c07K+L6wWx0BhJg3xCh/sPhHbfWSsCC31m+y8iIO72K1kBkTemcovnZ
kudkmXDn84Fzc7Y9ARSJXsSQokB848UI6qJ1RJ1YcT/Q+aPV7Vq2Q3tI3L+qex7vm+zw1HyhMiP3
lmeL2RYI7GG/8J8M2/S0P3eXjsPfRf6iiOyJPeFFcHT9CiFO7UTVItY7OTy74HIunPkYJw8qNTnA
m+h6VKa7vjRdFxqQuktbRt8WteIMUpseWsQ7Xfo6aSlMVnqsUJmYJCIuHY07qaJ4ufFb3VWfASHZ
nBvkYnkBdDA+twiOci3FcIqvG7BRN2WYhVy82ONYxcwmxRyYYdfUFhGUEGjsEMTZK1EDOIVLzBDL
YezgXy8c4Fr2ccnnGaVfQVUGfHXdEc8Xxou+liH7zFH4aDzfp3btkgQk0ikNAGcqm0ipD/DyH4wu
4P/BgJohwDz9SnKM8+wp7fAZCeTgQ5w1O9JGkzh0ArRgTcbLDIZPRF07RhyTXStmBxkU2iJ7jYtx
kc5/pA0RO2oQt7dAEGsaE6EiUeyAGc3I/BVTky8VXtkmZdZPYapjfJLzzKa6diXHaQjGHVmk5la8
AkNPs5enO+vAfXPZjcpfFn/jgpWKk01xvFESc9q8tNmEZXByVKwRYOiFDckbcd/GyLA4QmZcAVoy
EZEXd9x9V0EMJTM1uD7M/nfZbWJj0iJOFeMOFkkgf9jZnRjxQsyPuB7y/uSunKeYczQn5Xi2cpnC
LAaHC5OuqkQOMNCpc7tIzmt6OnwYTo9InONbgxy4+v547Vhvpuu7CyWLF+16NP+2RzDR+PMS0xfq
bZ4jCr04DikxPL2/HE8omxz73OlUQ0/9OVkYcMBf/lDxPLdxRwvLoVAyF315jRwKeNQ57gCvjo4i
wxZHqxC8pEC3WBJKnFCisoBw48l+5yDMMQ2gN4tk79UaJ+h6xZCiQ7AhOQvOqf5pM6gJJ1vOQI0Q
E5bHSqdd5k1sQLt+qskgWbJ4sJJQeGtgUWnGTkCPXIyrpVAY2mzSFSTt/nlhVJ2DFJDupDxV2Nd0
QgqbbEt1YvAwrwSZ7uJNrwooE72N2i88S66BNIr/wWcmFsbFCYoqajr5w9qvKJGIf3qwJQN/OfbU
hJDqLM55HxJATSWsJLk0DFj28YEqTPZ/6GFXF3cUp2R/Hsx7beR0tMMSmTF8j+jf3XdVLom7ROvp
9mfAKmT9spI1N3NJDbOukEXGGw1N1cxrQOVzSQMFYe+0OY1/2SKnLAtqGxc77FLll6zEHPSFQ5MV
J0gkgmNVn+oZdXs1UACJSVvmW+E4lEPkjFWw+Bcxjy5mit40w1ZTfUDc5unqO+fZTadGxXWlikvg
mxC+1F1CW0whSHdWTINPKkddcurck/0nOi9kmCMC9r+sGN/pk3zUBXbs7r1vdGBltI9yMbYx8bTK
w14aAZyR4+bdkPwCVfwesufZmCF2rbiUJRaKVYx0WyFbm5asBHfWwooyi1Nl0dk3tot1UMaz7iHo
/rchnSbUQjxqt+9YyaBbYcwnYPWqWym5Vp5Wwd+JWoo713Fo3TxPFydrt094flwmEUsh3Feh/q7C
Ss558pHMOVYILzOG0iNYMChPZgpEcFo6ZlEXnUea8teLzCHS9GRnVE69H15kFvgSje7l+zONJaVb
1Ng/TkFQ4dgQKbyWKMoXZuWiJ0pSzmDVOYBbls3leIqncpNntDgbI/iUl8htz89EhAfQJOXqQO0X
oFmiWEUZ4WZuxyln7fU4ve4rp3fCEVzlGgIN2gzpt7UyyU15HsSXt4UN1j3pl+DePnyi2piO9R5N
GLjMbV/QnXmkKl9Jdof2CfFsZgP6wSpcKqyYsc/4wZTR3hKiF9L5N70obBOAhWzMsWLs/fMWwq8J
xRCElS+7+HYn2Zm7jYPvGZldPWvXRPcUgvayOEmCwzDF4zjYchPI1pjclFVbhUJ/0QhOUgR9QbfH
WqzbCUjRzY2BEFavi5kM+zbMDhI30M1gOXBRvKy/reKf9UixAZwOLWxcU2YAyQlqb0pHAa0r+SX8
/r0INPjRTWawRC+FzdfsQ2LYIUQhbIMN4Sf7bg7VI31br09AUtwZhtAf763ypMHM3HankDhO+9aU
4wJV/xkfWBYErB/CVKkMQc4kV6Y5j56db3glkKU+HKZKzeyOZ4JBhpfCG/wapkeSh23sUD5YH289
Lk7f+aDkSXr1nznVW6D/dOPaNMgo1aPFSn7NbIhOTbYTCV9j0Cx6SSW1x/Jm5q0+f9cgLMh6r058
KZTaZ/ytpTAGtMKbPFXtAWF47+yCeAmPDxljqcox0ANfzOzyvG6BdkYgRzXZyXdpHcry/Of3mTVK
GvIClTjnn5+xYkzEN5H5gdsAJKtx2DtnB6AZeT2nWkN9EF/+AJ1Kw2fVO1yWsfGshbZKuocjeEUY
HUW11Qe1gckKN7pmVu2MBIN3vsMpzja+PMWK/M38KciuLFnTD+JppcLV2UdmjvOjw8zd4MT0gNCp
BPLsoycK15Wtf/CICfieuGbiDJhdiw8z3p5iSmtcFoYEvmGzU7i4j9+CAT+Rehwj9D1xPlaHkSMV
FHzITVwCe3OG2jWCqqzHHBCC/b58QNcKeAXMUimj2BSq+iMbKHBjSz1si5Rsc0KnsR344wVBXLBX
IjlSEQ8wogzRU16yaxf4lEtZKGrxSTbFiXFe+LKb0dbsOmUd3Ij4OqogGyy71UG35LQRZ/lkZ5/i
Msn0IOXDn9Et/DjiObLcLYooy7jzMYZj2VX/QvfoosrAI48VYP7C1tKi5SygpE2t6g3BAPj/NFD7
wNGYYJRE69MndOdyk6ONPjlQr4P+othtiwMqP9aYLr1EoHTiMNEGesCYbis4G5RuwyF7+5w69z+E
5/kQ2y2rVpanFlK72ov6Emc/5Y/uj9SrBZNWQW/FLEsAFh867m3gvUnywSuvrNt9BcJavi3Y0tMO
HOXTsZJvhUTkNvuv9+mNGB88aibh/2W2MWzwm2qEi1mpBedQWPy1INvWiFJbELzIf1dT2k9Aq3PT
cF2tB5smQ1DUjuughOM4TIrBy6wiYD9QsiUWLartir8HNS/z9U+0zEJG4s2KKayVYtlbYNglSUC+
a8ao2BV2AZTVFEOLHFkIffpJXm28CgESOK0gwqW9GWBuhgUnUARhkDQ2i1UFykw540Wudc2S6CUH
H5BRab/hxCQKBMXiYBhyBNvMwNA/IbT1rhi7YzOp/v///1EkJG0qFyEB6HOsAnhL/wCfKOBDaUAH
iGi8GdAUKcFSwX/Dx4baC0JDh25gTjcIbU0OkJ/hvXJ014AAkrfgIGDlqY/e+AwpPX/eiDQtercd
DkKYR2QpOXebhdAIH7iyW8BvVw9f7Ac9Xaa9KdaGa3QXepexnv+g9vdtuNN+QkbaQ2hnDzsh2WSn
4hLZAkXxs8BKTt8K720QfymgoW0GicAbtd6bwhNgGNhvIFsFU0Eeyn+htB7M85JItZl+fOOP9TCZ
4CFLJ0S+Ud0lmkQRA6smZCAONcyIBvHWfuCebSRKsffWO471mn81mv+VY7NdlqCADCWOLDXkIXGd
cmlmEUCgTj6qcQt24db9760oxnOZ1LvW/Wv8Z/U1z1PMIMdj3dVs0fo03OUuJ7xgVXmhESVJ2F0S
GTrflBa8O4Iubh43CvANDe0obFs+yX3M4xziNtr6pFaRehErIqFYsp5ufRWbGRSBXIUAWdx38H4X
vTh1lKnATFwE85p6WPmH1gpg0O8KsilxokewPbeOKvhmJ5oi6l0DasLABxS2GtB22T3TjyibjK4j
qHDteDFyAp+U2ftOmff3NS0aSXIJHM/uYoEHYCnCfCCnOhr0jCD9lhOUgU66SOhKXpA6k4rzpXMY
qZ7Vweqv9Es+cTxuwiVCbew1VYEHDTbsW54+Mm2FWqxm/4a1PtjqlasuVdCj97xpqr3FQqPTXJlQ
oewTvcq8LTNlx5F9/PaK8W4s77enThZ9+EnCelb/Zge/sRidzyMSRlF9wMupIcAcaw4HnT4cdumk
oiORBCizQuh0QJ3JTzqE38fNLLyAsmfObBMw/nMGWHIxiLbyEdFtQNCK0PlDGRp854cipdTRUmZk
IcDS9anjRTleMpy9YryCv+RhOgYoXW3c8bMgsJT5Rn6SUjpGCj55c7cVoIbTI/atXwtl11dWXmVM
SWt4epf8dlZw9dKrDQnRxRKR7PK98J4YA3H/I8u80eHndYMmEgNn6/nJvtDXFADFdYWOhfKuyEoS
sOS72F0PrE0nWsNmycqQl4hqJ5WybignqdCW4jeAspCz76anTjXmG9ZnIB9tPdhS5IIJeOEyr7Fc
X7hAp0LtVq67Xlw7mFw4Z9URaDClTFnH95Jd+3+WwYssqVVsg9rS3LYX1H1zJbfVsotQu7qBG43P
TIPci7F+mJoxPyTcLQAnzrKE1XQuzemmlf1YFEvzvZyBJusmVZ2XFDcSJc4tPLppL96xtRxCmmwd
Xwld8AJOiAKF/SsRMTXr3SwdLsXTk0LHV07yLBD0Riwsx0jLbEvwVGjZqyF5BWCg2FzZoAY3SNvV
IXUnQQCJAUfeAGWo56yZTgvI5trv4EWDEIbIWuyR9WeyYadq5UEj0kxocdQh/TbGOM43UXzMHCjq
qY7z/JHsrs/7tc/i8oM041YLxRAkUfYr2nf6/JNpM3bnw0pQwkWuz6Abqme5O1Yka5F1R/mT1X3m
U+HdkuOuuyiP/uHYB1hKDE/dbwvr5nHeKlCpJiPpXKjkqcrxrR5tnQ3FltVITafbojHzxwftzZfN
3FJ3B/nKkQPIk/jJXlt9CbWZmyGDxA+FGnQmUSL8vDt9ATZIj60vmAqJTC+Jjny8NDKcyxzYEE1q
zfyPvxlhcrqbem7JS5tnDZEhZpDNOmCeYZ6C90uBuU83Pnj5Hnxx2ubQqRALEc9wt47t8SzEm8fX
zRRUDL5VFBQzkEFoHvCMCSR0c77Gch7NOUThQ9UHLEAV3VHVBTieFrcID84v/3Gaoz639h+8nYRA
A5Ux/HQSNSDREg98IxtyBzQLXGW9fi6vClT6o84kNGKGvLMbYP3wf5gwE5Kb3hHgkQV4aDyRa18D
P3kE2sFzKr8aKKc3D8YKtOneNLT3/sVo2GYLdcPSvMnIMMK9oBPr9yioCE5QJcxu3dYT+i5uf1xW
8INDX1xDKeQR00HXtOeAHhsu8L0ArIwVS9H6HJpmdD6KgGBH+D4T/wXpHM4tqQJJjDXctHNU1rCS
9TZwyzCUW4ojLt/sRxhEhfOKglcNxWw2bmlo12g6ZnwuTCRvZAAMwtSYWpBCD1i/pOo4MOYdiCs5
Jg6A8Aw75a/8OnczKdfBPN26vr4YOvyS9N8SPvFBYFwXZXLHwXg9A76m9cvo8aNkv0bOZEzFXebe
WqfVYSe79ufS9JR4rRlQqoyglWRR678cjG8PgthKCVX4z4EYZdne5VscETM8jmxhotLf0sBRES5n
v+CkC3OJPfYIJAGXzii3iM9ablp9oN3KaNQOhdxU1+N1QuaUdf3T0M/HqDQEUm9ASdEMHyhztS7n
yKGLqal6jnYhneDPKuZTtnnqrTlOOW0A7on5lbxUJxwKmPuEQesI9k8+MKIaYxHxjOpF24On7HH2
6AZZC9tdxfBjNWNBU1KKVe1LRx3BZr69T28dadcn5TjuqKojQl2IwhhjOPpQMBqvmOr+enBNH+wv
+bhzaejzFlQWrjPO0FSAw8iYNTqo/iEDvZs8NtZBJshUHQL1dDUbPyCpPDPKv25rlVNToiNIl2YQ
TP3Fl0SDCZTQE39PgcU6MJbov/efiUIFmuoS7jLOgflAYW9hoEB/Co8K8UXbYTG1EmVM8rck5VtX
AdVpnLPDGf0KSRCVKetQjqgFDoIznVp4knlq4sczTChScCMTffDWC6AjZ61rzDvSQKdeD6OPDkNB
GilB7x7hQe4TiNwwRhUjk9fwy+0L7WXZHqk14iHs6LsDlRGjltw3dwG3t5/ZWy7s2Ih6DneQ/GW5
1g4qy+1v+8kNdD1Xgfm0RhZ1PT1AcmzsQTNYFKEx5B2IcW7GF/hsBFkuhJchZ0ZkWZZVcALslr7z
e7FVZRaxYNArVr12iTrGxIq3/QAwz958F8UEXvn5WbkumRqffwjoL2By38/GB47R73fa1fZszN2T
0q/iEouAPgKFVg5ZRGtXSvMEKC0+Yd1rKGE1xqYYTe6f0ZdtVgFwAzvMM+x50bE/tjjPSFYsfOZr
tA6u78odjt5LPvOlxcZ90+0BLUSmU/GmLs8Wx9uKIiCoARKDatG20+pu7aTLnCrXYpU83jJO3pkq
/1n+iTV1vNaBzeq4ShJki1cmvPruDO5TBYLAJkFBDZK4fqRC2AWDXkuyXAVGzlZEXx91ptG9jeGx
23PSlgfPJ2GJ33jENPLDZsC1lK77rU5QsgWsK27MoC72yzxtkngT8AjIHEtIGevUARLY3ohc2/YA
pJq93yPaKzs7m1w1DTV6/ouctg6E2VVcdo39vGAEurc29zChzzFukcjkEPx58BJytIbd+MbXMUeU
9pY/fXkLoALkdpJPvF52mJlkoE5gjXU678HPFnPbM3EN8F4LIaKFfI5D22byhbmPVhKy7CjnFKcO
nJYr1A4cfNmlqe2PffzlEIKud9LcOYDnGWnXObcfKuqVs6i9adStX7Ro6cZclAIfcM1+GXZlOhSq
cj8sGdEDzSLDmOvSQKRiWz2sS/ub9P2evnY74o557x0MQnspVcB6KUdISZNRYo+DTqgB/OV/+Wka
ShBdGUshgugw+ywXwuL/sHllHtdoho0MNKwWXUjlBOR3APjvY7BqOcvGwVId3/0cgnPZ1NIkQphE
9AF04kQAXQUo1p9/Q8Zf50o/raY5D/cSx66DqyNuwwS/nV4J7lJtDLhlHzUjgzJX/f3QChE/iNCX
Ca5KLbwzGfyXQhClldrgctKnxUhrgfOpfwQq2XPExSY9S9xksik7pOOaNj//p45HYec4N85nO6nI
ku9aUb3Nm9RvtnbOSTLXCcdR2nCSArtoJdR0ZYpsS+ell8M1JfOFXu2qBEFW3A4AvXlRHtqwVFDv
Nyu/YcSd10l0Wzm6/PHxonZI//mJPDjkc4mQnKkcvgwlB1DlRGdkvyH2tnMYGs/90NxLG04o5y85
8IL+Ybu2aKN9lXzWA57/VXoPS2Xzw0zhetgRbzUZpgrWF7+zQviCwjF0ZBw/Os82PDB2vEF+rVUC
67CjOWNDgWkYAVARFhPQ25FTzwNjlnrGMqfu7wv++t6ol+xuxxpHzvtsyFhOfEmTj8OHJrGQ7NBu
NkL+hper0XXk/on8W0eEJI6OCIcI0P1YVWMh0O/sAf9uVy4KZtz3AcxmaStpeAXJ6wn3w/K65Su8
hPlPt/WdISQOSHpf8ubBPDmETjYi6lCafFpxsYtwFDVs1MYRK1FvVHuwNesvQ+yk8H7gZUn0slVh
3Qu8C4vOrXMk9mVqNg6LvcT/kAkGy/JV8jqKmkrOuhKDlGBL2hL22KAuE13WWyLO8RxTnkTCi8+3
HC3chuQ2Mz7Dt2b/M6NTaJTq26+SZLpODmd8zBgO0xl3hJaS7pK0xH204k1EsnS9djQhnqhU/HGs
+sWTzFvBP8jUt6BYU9x6ZH+Svsfwc9WT4tmUtDRo2JIkfWv9vZOlCOKqmP44TbxmiWyvSHo6C4r5
K4o9XLBnGsM1R3knpNP/9xz9WHQeIHNgOm0uT9mz2dYdLXl/UHOzlkkFe5ziJORUy2nbsbaBKLyG
kE+GZp1lj0XOdQE5n4VeGRRbD+qQrWHMRmAlsXpBQ/BU7joVqIN5qJN1l9OAnvxpRohDYUrhHqqm
XZE8gxIaeqIKjCyPZxKR/Xhjxe96uF5YtYhmm3/Bj4nD+NKbsIYhbxutuK1LoFyh1XEXMwX9kSfO
sWvdACJcCAIVf+F3F6zPoolDdxH1zS+ELuLnAwYDtChHlZso5C65tcR9hy44u6rBUNWF5FVl2b/Y
mNfth9c2uqPrPRpHGt+6f0IRWd2El73KP27ytCIU8pmJ24G5RuayAIEwZuthz+jN3pen/2J+HZ8V
CMMRPIueKYuAeBREVU/E0db9taRnHxQLQJugpzlR3+kdAFO3AgO8BdqA2I69fzb0dJNLEXtIbXKn
NmjJMqmMd0K8JeVpIdfbalvkel2BZngAcCJd0IyoSfQzqDkEEBPH1t7YVCGAZ2pSF4HenodzU2Fz
oE+HDHS8l6xCRTIv8prb4Lbsc5keBLbFRGFUPgrkfyU7KtWSacuX5nXMOOdqrV5gULOb3zgthpvd
gw+9qr6Xp+UeXmmqEa1Zj9BtbQ9+EOwXb7LEzSQ7eHzchH2bOoyCQpPx5qiC27XS7LDiO3pIDMbs
9Tgc43+vm4F4C0BIpxpZrhsxCJle0kZP+NBlDANY9RhVAomi+gfaDyKWyXpoyQy8pLGP0Q3/BuN1
cOVEdlAwIEUDQo33sw0CLVnVb7l/45gTMlkrgVRYkEiIqdahbI29gyWfqVRETxaVkNUEAckc04yX
7wzMOailJ6c988Kx6F6HUyswNOaDB2Y5fy7co69YIW6ROHHdeJjbCCy3zIGcrlh26HaKM/HYbsVJ
gCTftAyyrM8IUhCzpdP6gtLUZto7CGu6N54Fph100DZA22Eoc4tOty3DWA5fp+NJR0gzUkKnAHVs
z62sAvV1u6Smwa9lLlCgDFmDgb9FoUBhHSHvBPva66/eoxNNbrmPpCETqkO0undetJNx/RUidxVo
5hYoyVbEkWRlPo107snV5V4KLWQxFOOtZcCxbUpT1R7cT/erZm0X9T4Jy0J1zaZHP3bGoHoCn+pR
2OlAK3JZ0om9PMlr1hlLKYu4PelmhzjR17pYYlkYVE0NbnscW7JLQGZZ7jPHFiRrIrqknNERc27g
fdo57Ll7VGJ6nrrv+eC74zLam7v7CtT5ydb3xKw5g4LByU30ju/jtO9mAA6+f1/6uz9vSxRrDIy6
IYDkYhkCipfNFaHagW6deTfhuJLmcUC/OsCJrwZF4fUviHRMrZyYA7xt+plC9cG4c9ow9xFWdy/d
aExLJYfSpzZ0wdhbu0yQTLKc7SRTv7z0+xT+KhFqAJtGTIPb52P5QT9IfyLyl32/FCG8c81isEbZ
TPiT9ZMKshUy2fujA4+kKIJsSq3Ha5atHc1h1rUpduMxRg/SKB7sJTLWKGnmrD2CxiGHd+ZYvkbl
2xODcnuUS6Mxxhh8WaZQ625xVMXsQYVQxdqAKQFh8COl/z1/SZiWpqF3VEpmlaG2EbF5Te8ohDI8
FrAE+zYV+ZrxnM0FTQptyF4bWXvrKdIXf5rt8kSHdFxe/QLwMybq6Gm99P8kK/L6oc7zXssdfHJw
cgtDMCF9HMlXnvLPv7+wLoW4Y28ea0u4uFBGh5+xfU6yAXtbfFN+svsA/uhE3dsyb3ttezVl5H3b
tLcjwuxANtHu7fqQKXw4PJX4GB6IRd/5Pe6caCR/J+MZUN0uHVfUQstdj1J+x4qSR4l8UxurBVX8
w7YEpcjTnUYVohpJAHbnEW0Ec2yOHT4T2I2gR0+ZnfwJZA9mEfPF+oi2yaJ54RplgCW7RBM0qPQL
sieYYCILZuUNKKj68zykLXTE8BSmgXoK+BBt3z0f2uTshdkC8B2vXPh/tLkOGDo6iW5lv58kgK4f
26Aldi7+BABQutFSfRKaP2cOP7idOVTqqRkOi6VhB9aavmMV24rP8R2NwPjMUofDMGSe7uKWzYnq
5z43XcnPB0p5zTi9KVlBOd7WoIQVni32vfsGqT9BQc970ZwUuo/rBFltZiKE/OWpZvt9+olq+Lr8
1YrDbhPGHnyI+iXkwGFas8ykjpIjHNmDFZqQ4AWZfamTlqjELI2x24o3H8HMmntqtmyIuLQFDJ4e
19aYSz2+2vkklF7AuOLgExZBacEnhNX5KpDL+muzQAs1KMfjh3+bcFtd4AsGorFnvKgjHTwJ7Z5m
4EswrMmOmDTS1FIopN6mhMYQr3gVkWLkUkml+qvGYIr03TYQ8HrofChSgn7xz70A7cKLqYk7tkU1
Np7K8Qwpvw+C/sGtf3+kOzbbrDPdUSq0luFjS0D/FZqNh2yYExqyzuQ1I9GVThlD/nlQ7lJSBum1
NodF+xVFjrcN7tHGyIfOIDubafdF8xSKxruoUXEBZY7Pge17l7XhxuJltxWnqdbh0yJFGrcMoXUb
uPOTpvSPg+1+vJxWxl0acsPb/cefYOm5sjcmB4U1jVN3wUT1c69o2XW+MyRYx2PsdqJpu9wOTmNE
BNXIxb/Vgr604XjMPxsT/tp55T9kyjrCuujf8FHhuHC+w3cNYmNQtKK3sVxPUjybQ+lrC5x9Dn+G
clPakJodjUdwoXcvaZG+2+MZ7IcY/M1WabG6r98/BA7knqLY2YLS+Gk7ADUBgYeQY8l2U4pSyNvC
gTgSSCZZNginwzbK+RlkzC4N417DIv872ByG1s+q1ooWUg5Z+loTLX8JqX4KJUx6MPAGHRaKO1eX
AMhJhD+9zBAxNK4mGTCflX1GjNeR+4qxpH32Yjqefr9WAWcpm2dJv/IWBdIn3nCPeEsYn91BLP0W
r+l8WYqcA/Uau+fIbbeJSSbszA1pX6OHrLrJSKWQWsJZjFmKMBo6uls946oD1TAgimgrXl73Pcsu
okjWyBEwx7ggwpNUetO9C20HRZz0GJV6wRqP53ubsQP4Ik2UNkCrkXc3T2IeIOJ2EOK3zaxfSK3x
+uJ1zV6ChHSiISyZ9aS8on7d4Rsgh2v7UMOb7mGFLURVq6Y3oF/JyCWHL7giAz861FQMhuTUeZd2
vyuTeVbv5GG90KqKGcqJPS3eo8fkXEWkJgTXYTky4Gu4U+JmD91ixlaJUybRTcVYSN+YVfgvVsWX
aP//8TxQU5ZUKod50eVYSheC/P8obmrO/EAnAiMM70slkc/ShCCs6N56M0tTDthp7grRM2WyQQH0
Q6lyybUuwGHMBUEaVxLuUIDcrrtLN6+8qjnBRl4j5VqL4rbl1OHUalB2tEZnjDDXg8/PgHD5d5MT
x0Ll/ny5B7ddZZvVnv/YgicFIWIA8ym0yNXf8qqJ+PBctMPYg7ma7mbs+F/8Z6A5YkBImj1GHS5Y
oMom49vex87dMhc2ypBOUURkSrR1waUAFFRF90TCFEcoHruJ7hVcd1MiV4hONy2cKP5sqVdPq/WV
o5XHOhfEQ8gRSSycRqxItOaEuCkkv7MQUrctrAXv6/Jj3igqnPBae0yrUDXDCv/Nzl9+H/0AwOW+
FjtPSRt1XL/f9A4qhfZqcLIkteLV+YvW0rrhreoT40GysHLyhiGNutuOYe2IVu7G3kYQVoKOYWSY
yCjydgiWvzrZn8grlFAoqP4Y+lBGU6Omo9+inZg0GKCrTyzsDEfqM62R2KwtFiE+Pb0m743q7vGN
16NZopBTs1pahhNNzSjVTPxsCrtoJaTZwdL7b+71uMbyLeI9jnLbcQeUxY1VS7hNeQkCTVnBibP1
EcwOGDKr660Zl8rePElnLswJY191cvToG+IMO7sQZ12Pe27G8RaFDgXpSaKghMjLk6yz7SgJnW1H
rILwqpXXH29ULII0+/6novqMj0JHWHEa+eD4TOk0CU0tVOdpiDcxW/Oc24S+602AXPA3oKlyZkiF
C5E8wP1K0txZGq1jBeVw64D8cuifYu1KlrD/DJ3fcw9ezVKF441SsPgcDSawWQRqmncz1WvBKYaH
JKhWP0NQNxr8URBQWNynAwgkIEHEVAJ3Vv0DLltzOOYSg4z4WwVBXYwjJSSFY9sRlVfwUKw0GEPl
jNeFemrq6w2Cfx9UXRPbdlxHQsIs55geVAl/wCIRZxDApUuirPdXUXJlMVulKsAdybxPknzIEc4d
VdFVhKF46ufSmOKgRywzYEMn8p2AsrceQUSJqthA6HuxJzK/Sd2TJsgBmTQhDWJwcBQYLRdMLYoN
gdVZY0hfcQgsSO2bi2GFf3AXZzjVYULDoMYIYIDMCiY+1S834aRR/xKubKxP64jLgCmevbuo86eb
C9JT6UMruz0ZbD/wuSoTHfGspfL/nFHQAvF6F6169n8cgKUpSSuZAPiA9SPOx+0geQipSE6AQk52
GSDfXmPWoit8CJft0JiTP6BarA0JqbgWGTuU4pgmZk3gg4wu9z33rwosVVB32mb6JDvp+5DmaohO
XSxWbByL1/4A7r+BVaxzBEmxe/UGn9JUxD+Q/NVJgtGsfuL/2aaIRLNpJaaTH7L4buLsrSd0E0Z6
84GdsgFFtSsS64X4rXiYvZtz+5rtJpyk4MdyB8qBQe4fo6RDRKZJHW7ZOW07HLekyLo4wlxnUUUx
Rjeyr6J/7654t3jrAQqcrqcEgghadhdGkwG9Tc9t72NK9q55FFnlN75BmIUiowo3a5zBfjx9UcPG
b0+Iujmy3qtnr4xg99bm/X9v3I0XolMmB5XqdPHDN6QgSU44sPdkFYphe8HZDsjpJW5xwx3hWnrz
ZCvGWo4tnCRbPWQpmYHX1aG8CoAyVEVd/zEuEtGJKyYapbCG68LHjUi8c2hXCrlQBhyw09LqDHQJ
KLWTqWYGpOg0oFF0IqPddp0UyeTmnH3+EDO+vDzaCyHMMcuocUWgbXKV2kpIdd6sEv7qhxvUiaUG
xSED49xLSHQFkY+rE0WQOFlME1pp0Khsw6+8I0MUODnHRMTAwWgb/q/Z+az5r9nTuJsoRW/6DX8x
41zK8/AMP4P/0yayCZiAe+eK2RgV5FRannh5GVi4kTSzkBkEmBlr9b6Ak84QMpj97UlIJVb1YW9A
6Z1rt2rAS1nLdpMPAFxYhBFDlXoGUXL7RX0wqnyChPHb3WbrRAgbL9PlnQRzV63XOX2eOoX9Rovg
Jv2C7PvLYqMhAf09ObALCTmO27FH/SAK0a7wp6mVdwEk7SWd6iWcbngLJljYgMuT3KY1hjCUrYsA
vibVkuu/0PrpezLjE9RjTmCyHS+5PVswyXdpSNGPrWKkz13E8spd+ilzQEriZtDSPjuLXoPFLsZx
XJSb7KS22B330YdQVT1J4wRxjAft3uv7qlMOv8xPD2ldlQ6r/KzpBwjQQWk7t8LvqNmb2oUdcpZd
DT7xaviBQk5Ci2XF6P5u1lJvGHGSL7DM4dqP8ewwe18/mMEjCXL+THT7s1Uox20bWbe32bXg5WtN
KThLxNuit2u6zeg0XuE8Ab8eBYvcaBi8W414naCphG/4lk6hWMh8L56Vqs25cmP6bMPwPxC2JAQS
hL/BofLmO7oTelYNlXHkeU9Z4V8OxXOMDB0NjiGRHpqUKE4Ccq+3ccgGPdEYNlTb8Z/JTzMhKTXm
8Anq7uw4IeTL9f8J/h3TgW2uwgyqJaXfFwG1JzIBj/04JOg8ciaumSesbehN5wGM5NAHC1Peg1bV
VON4BHmTS4cjkYUrQui5hJr6wXYqVw2bcu3g+dddWD4Zp9x1AApqBTaMkgjluGlp6nyaci/gbS+g
BYSqOCHUM/iMQTCfSVL3LH55N8TtUQ3G7Dfk83EyvAe+tCrZZY/AbXFD9j1FnkMShlKm66lcirR8
xIvxBtMC21KyMPEWdckHCc0UMAYNiK+eoEeMmZGInoLz0wJjlZdW91uvGdaGPvhvNZABiIhW3JR7
bFlC5kRcGG3b3QYx1QctfloJ0kcw9cbiQtKlQUmrvAeyiLsoyjs3axAguA75wVqA1FEYNurYzJ+9
FLPvqaoT70yhOdFq2kP9CEQ3hipNpdYJSytbuCIA3s8Gnkixnxhci2M7mxbjVlmyVQ4t3rfjuGaF
L9oMHdxUvzQHgfnNch6EcfegXjFtEZAZCMYOn/CndSlHXtXUt9Lv7uob7G696iWp2xDr+INYm98y
6RvEnEfTWpP4dCTY2ZvQYxaBvsK/X+KnLGJtdN3d7tkZneOhivb31obtFR2LY3kK0Wxl9iROKks0
YKusI8cGqGle3BX+L/J5ej6KlZw8AA7P//Hb6uYWRMkYn5JHySYiGklo58krcjxmjTMcE1oa4mjT
/xDUH/VJgyH6butUirkOAS9WMnoLEoAnxEp3ThUm3vVKN6MZIiRtvr6dUtk9w3j8ts7T8YRbkv74
hj9OXQGPoAZnoDOVl36YQmTBS+T6xeUsQWDXRrSGwBfoW8a7+bCOQ2C4jc8EqhicioOmaIxl+uSo
AVJT/gG6/UVhpBB02iX4cD5emnCIGIkip1nwpIyYEoh2dsrVX1cCBd9o8FaAgJATXP8FYJvwkmSt
4jkpwAzETB10wqF9w8HzsakEkTY1/U5GbucPVVOsAbPNLtSHw4QRGxQrfwSWkrqOxj8ZWheDBUH7
NOE7jS61EaZ74xG4vAuPp2kgvdOV6Nngcwb5tDVo/wbXWRfASGOlE4kD5I5h4JOJd9JRDEJvMwqh
b/QuykQ0Tf4ctPfgiWg+eTlAfmPWoWwqSlii+HJuuANX6aoidiZ5sY0+XvgrEqxyJl2TrjnLAiZ0
klLvVrZFwGDLtiBQcxaoLmog4Xq68XO02MmnWiRPQ17Us1hRJ3B6HTPEsxbrKgOB1V5rlLJytdDS
ha8pGtf8IaPsMyeJpJlDOWE1NwJR+H0ZsjiEOj5OWKSK6bgOJi9+i+OoIgfPwWRznbLdwOsrT4VX
tS43BF/1EYb9N3xvtYqTUNxqgnhFYN0oZILMpWSt1KbVmrqwN7Zv4FAH+gPenGLa80ou2FL40bis
26K8VRwqBbMahSY/tNn4To2RebM2rv0wPMnZwaWaJXJEjl1I/DHNIW4iqpZkt99lBKLa7jZqUhT6
Zf2YjMETaEOoTZOl/Ggftcf6ro5jmvdenCLQWnKAUqijXDDQAOYr/KEg1zVgJpGKu4gx+4PGIHX7
yjtmWfR5NgZi5BQ9MZzJfbo4AJsPd7WeXslZuxh7A1DFmg8bQJRDFJZJh72sMwLhxNINVRixaqeZ
48XuwYhwUwBD+M10wRJgqp8uu7MuTV5559QQ5c38WUcXC+6O30ULTUFuZxQzhJhnTztlN38wPJkq
bOuxmuz6Is7ycNUYtRZAtXYbqqJhjXG1kV6HUu0ZG9lez/UtJn/t4CGEV6TcsNuolOK9seIl9ydP
Pwwu0IisDHspQZqpNayzpbB0xh7az5EglHrNpP/FvX5y2O9xAVzxKgAbtVZJGm8Th1Pk+hJvMiXK
25Sv/qZrJKoBl4/0s1eVDL9DoQ/tY/1RTvgV7EEtMwyK0qXMbsIVOYLwUUTbo7YyT2b9VE5WRvIs
cj+WFKPzF2cwUAtNvLH8lG4vDtBhpTquwU3APnzr/jDsFEUrAd1otkTgkO+2Sz7u/5vLQmGXRMpy
Cp13q/kjOiJ81vtkJdRtyvIRVqOf+hKLfCAMIU5SeI3H37kllAPb0wzI3TAPm9SEDIBRnQdA/1k+
HTe1tvc4AOaNTxxHpmHcHvMf9okOZW5Qsh33oAeifqhXztUA9QdmFAwls+vXMFOq3wTwNeRXYH+F
kkFP1dkfD0GhVdf4QaQ3x4PbWLfGiGWW1FpUZ5KRw/bwjxGZLAXokNzp49KH+O50eryOEPfpKGhZ
1vQUeTbr24lQm9dm/5GxF6lNxJS+Gw0ax9zbOqjYlWgubCde6g3cjgwkLkrLe5PqhlxmeQrUmwQM
SgdIWOP0a0NfyV0M9HkNV3CPzY7gy3tJWTk/tka/eCo8Nt35KfQL33r8Ne2rP2BkZP327W7zAWSy
TS5XYSvB/JZwLWoZ5MKDF59Bpyw4UVM60xSEtiFKE0tlzNTnqfAiibZqfmy+piTd8Kwy3hGsNjZf
rvWmgeis2YlaIbyKEPr4/1EicI/L00WbsBcJslZtrYanyRtYsuO0IH+9PGQzjxOp1ZZYjbROs3eh
YF+GOKlIuEtV8PEu39U3IY05PGYumIHA7F6vIGuWZDYPtQgAKM+z6b+L9eAQ16w8eRhF89X1hOV3
Yv/24+fQIoWSiQS8QTu3a/7Arj0TJrKBpBnQLIluaXbnGHFi1WvWgUns7plZ9e1atCCtvf2EN+fJ
CbU6jApRu3xAIHij2b1pKc9LRqG0jwFhbT244pnw4Uax4U9s/t1jWoT44BisvlgyRUOr9nBDVxIc
Z65PfAhCJtAn7pxKmaayw1nsn6ww/D2tmF0mPxhQ7XvidhdJ2x9yICFjpn4yD2T7/1F2BxgSkgpw
nw88r6HXpy0bPRVgw2USlmfediarVVtebusEbbtzWnTwuz4CH6krOK3E5SrMZaQ5yZ65qHkTlSf2
2rq/kdDSNu26/wDAPlfZB1ljQjq8BkdoiabDuUIka1YKdtvReaXOyVTIgPBcjhVw3T3mor/PtHju
5ySW1kIz+FXSPP+l/PQx42/Qqv2YwhUjCrsBTRac1I+6QuQLEAjS44Doqpy2O+lTskgibZQvrEut
vC8IiMinUiwq1qaKmVDab5xNA5vLzP23ye+0Ee94iGNHBovWzpO1ZpDNlr3ht2aHnLjFYy4ddyVu
fn2uWComQNhcWUiTvqWqpsID7inXQSXMEC9Td4UlIHMVCAM/C5ZI4J/bfidMCIlOFfwI1N/TRgXg
PWrkZ7g70PP8jlH78fbhYp4exxKSWynyd6wFEgNNzRqc3VR7blwNInmHqVaA7+GxTGSE2ocuuO8K
4z/u8Y0CzdrCjV4ZUnxWjpN4ve+cwGGlr3ylivXOrnpVZh8DpodAQ099+LvkXavX6Bx5e9iyhQjC
VihY8pWl7ZRtMsFtEMuHdTqPhHPSVbx7kyRrJQArUrZPW6ZQdJzmFyy2tTxSjglrFpfjYrVIVtMK
hdKOO1auMmKjeU/Hq72RXBMY4s3QnNYuS+iPPnot1NGdayEzM6ob05WcMf/ZQazgMIIi9Mr7cq4x
fULlYa8iThjevFWzjv49RjXIPxjautjjdGE0Maae910xghbvFWEWty0tU4Y5xFr2fJySbzoPBOGk
zJxTYBgPno7S0XLk2RtegflH2maDanyomoWAhjlG8J3sC5G0Krnw4pbE59eCRclACboieaZzYaVn
ex6s+mc4mEnw2ZigLtPgwBBDmYhUiukSIBwqmfGsLuTZ168ikT2VszfFr7jpynX5clvKBG+MyDQ8
6bJVmy3CM0I454D5LMmtkejyMI8iTDPDJXC4Ec6JyQw3LsdWquFBDaii5lLmj0GxoLqea+tqND5V
c3CyuEQ0ouILHjp3g2uchieYfJCgJfpwueu3LUPpoQM868PGEgMgmwmhpWlzjBf5pSd23M+S7weU
TWqAS6154OkVf5yEaVi1cQYdijLUjry3+SLvykmbDQ3ocpJ1s+OQYWoEx7QWzWY1x9PQMVTxal8+
ZPCh9ZazykQNoVCg0mWt2W3+nhx80+1ua9dThaZTfWjkuJzv19r4kezcPwZ8/yZCCzExAUhy2yID
J7jkcT6JCpKl6Csdt53O1VbqrbswFzlHxvVyRO1MNulc07LAPOaRcJh+yACeqfzIJBppfQTX1lqS
dZS6BPXhdPYl1syEFCq922oHnKvguXbEH//BlKTKPtm8B+DfLrBlJ9CZqn/Fos9l2EuH8BfXmZE2
pNg5Ohul/t7OSYRjYceZ3HDKR0eWVNZgaKGozHurpfdXGLZdnCC5N0F4RZGif39NbcZdlrCH82KM
eWsI70b697dmndGOd7JfInJLN6sheLD/pfV1Zhd6sF0r9xo4R0MEfa4l/87PVpppSUekBTYljzej
wFJG0j4KIbAQBb1gZ7G1UD/nEWyW+I59s3P3NnXi47NKZ/EqUdZ83nZ8Ylp42Wr9KUY8y5N4uaHX
VolwCpoTWyIRsaRalrV+Sp45W8GIM228YIBFwtMWZ0nevHZAa29u1lvLjIkOsbBNgvJ67k+sIE23
VsBpwlvSOtgO//3rYgY5C8dArTIu5durE/x8DA34fRSowlEwWh5EKlg/cWHb0BcIFVoBqLbuyOJo
GZU5ogwgRLE6DHaU5xG1SqN1PguAs4+CxAR10J6Dbjskju5GFQsltNUZUPZDyWoytFkgflBldODK
X4RBw/UTdv4/10DciYq00mxGn8w4T8w8PjCoNFwsYKLn+8CqyhmQRHmLVz196eeiHZXGMEAzVC3V
oSX3yid5ewKwOP1gSAdrb54qi3b/hNL7hD9pmU5HyiYKK13K9AuT7pqyOy1djKB8svQp8LZyocyD
PSeWxkdgDCRrQCVo1exnCIljiJ4Us9mktUn5+prlyqHkPumlaNEIjH9Bw2by14NijNLxBEuMy0Gu
h9T5CKbwOVxUD1h+ZWeY7GKwoNAB4SKEctWoKxLkmd5Wt/es5hIt9oWibqLIh0s7t+gywFnBHgTd
WCVCxM+Kx38mRNz9VKSbKrdfQjTwevP4VbvAXkYEchQ4yl9hdRBer0TtHglcyrTgeZEe7C3NZdjl
TXehC8nGHpDGxJ+WQjpY4A/5ZXoQur0wZV+4nabjmS+7ismdVDLJYqFdqVNN5InAdQDCdhEHLdCr
cwXyYPkLzceG65Jgs15ukqTc4u5ze7NYrLXsvTrXl5t8FfHOoNrZ9iCw4thFsnOSAVEScCw43Dbt
s0zL93W4JNzF75VRShpW92MI0tfXTxzPEYWlHctjzvE9jwiSX+OMas7y3gkbLV1Hz3Rt81AdW+d7
UXZBdTNGTCw5jT0TKNcqS8VmJewLIJOlbttpoYySbdCvR+yHtwV4hGZDzBf7I3QL807tfozZl1WH
GHoe6hPgiEMrYRRrziktoLB42YxPr5tsdS3HsLM8QA8K91D2MH3ndqAwn+6Jb0h8KjqUCKxuQwsd
fAa35z8Hj1fwDZjJs3X448BGtylMlwPuNEyUm7jRaupZKW8+L4nop1DF4RBxYcxqla5/PUtsWub3
86hxVIWV3uADSSE7WHru0YRbexyKh2FrCiSqYTioixoIMyqgUcz9HeAtNDA/dqGyG/UJCNx9cz/D
53/7P6t2EPi0UacelzZVmy56oLCAXBPrUxBrKPMzerJWYzyLbt+xbhh7zOTv9kxSSnCgWag/qcT8
VPb+UCWa6scUssZ6zTeyTx8LUOTjJeKwS3sTcTUDQCY281ltcJDouS4ciktpWXeiPwpAxu4/QjyS
afLcdzpiwL2DNUQQ4nhLHJu+OgbRJhp+/UD5GVYwwgsZVBofvrMD4CXhT6BJpSAnVDc9cARn8R/h
qunXh/BBRoQPBqqsid8YZReZgGY4K8s/g5dqxF5y+bOvp6bru/y1nl6aKiGaTRCZ36b8gsqnLUTy
+ZdrOe9vUGKKbOUWilevNRHlaj1LHlWCpqqvdekr9uiMLOscuMiL3shJJdBZ+pT8D8lDZjHXuVxP
kDKpv7fVpOStUKoCLchrkXBfTL9OX3G+k35N0A1CdcGeybjU1BeWkMlBeCTYSLyflAeoWsiSxfsk
3Ge39O50LWg5xpVg0LohHyZFVBisHDiK+W36Es8pwEVl7FKuFKzy1FgXpgAG/olr7oSEZ2/MCDDj
dIq2p6ZDErIEfNVv8kDnIZNGGcF/v7o+ezms3GehdYWjdEa/gZZliL5vj8U0lIZMKy2W1KGtz8oz
Y4Uw9mzccjSESWNF2JkDNS6bO7BQlPYis5x7g71DqZyQm/ruUt9O15tdO0yBO8EAQPlg/tkaPsww
HflJ3vkrhfpbp5DQVVKp67+8LQ01Bl4zG51eKjTPULIRp2eUi/UCbWymox/yy5m8vMYLt9H5Ss9o
GOpICaX4XZgCL0sD+fy+5/QnfQFJUQHsY7FSS02BqnCnomh4/Hh06/iNv/RaPpWSo1H3+Sjgd9Ah
G3lIVoDGj+1fYC3f/NtHnLj5CEZZ97XM53/pWRYb49tChmy1MXm5W/xGxpcuLaDEgrOk5eDgRkUA
a1AVzgYGknJKKyJUbQAhcrNcNucFd6z1+9WZpXXKiy21ysXIRqOeDBtNewHe4GEC7kL+LCepxNOL
uyD3aDllzBfFiQDINCBNNAw/FNOQP+h4I5QE/2XFo7xz+UBURtgRWE884LgT8oKf0zIqF5etH8dR
isoL+0HDIxS1gdiir2vcQopCLqQg0Au+z+BLncyQI7ON93C7hVHvq4CtC39MqRY1M+WRq1PMhVtY
U+4SI6lwzO290OavC8CqU7WD2Kv8N0FcK8mvRv4+694AhKnq5qAGwXlWVJ8OJfyCBK+TmRAETVVo
ZNjieXUfJgQk/hn9lWv8JTybNoo/Iyj0zdHApJdm/YdHFCuTeYETpxSYJr816JSttPp0UQNcc07s
5TssysCuSND/fgAxOzi70fed1cW0UhxXnyhBtPgni9ASL6+nULM9FlRvPgiVJeOhGLEeyb8v5BWq
I3qs6eJDknPXkrSx9KZ1ihTvnbNozsfKgCnbfuwcNjMc3Fy8GMuae5oFJ6Us3Hl9GSDBGWWywWua
zWLVKUXxwnsMybxCuM0iT4/VOuRGgWVMLYgniqMW8jhdxz2mqvMuuMtrtMVS55EkZ28wkRZ+OYOo
j2u0BRN18yY9UJq7WdvVVC2VdpUy0djDkpIP9fpE/Z+D9t0NViXFP3bWHyolECuu81lAQYTMZYaQ
qp3J50csrcK9mIV5NnJPib+4N2EoXDOaawwEyL6eaHUOAoBCrlCQqZMCV5heXLwjDPV9cBSaHRgt
58D+Y4mB8FvQHM3w9NdLg/6ETTIJ7jGSPcItIXBrvLHmtBDmYe/UlEnNhrWD50HsH1/6eqbODXaC
M5BbyW93G4X80AcVUylg9iMB5zDCYiiM5q4uHB1hho+7BpU6FFNmXVCHEONcLd3UdDec5CBut9Ac
3WCG+GACYZ8B85LATMAtXabNp7wefV/rjNHwWK/O4tc1xU0f17HGD3fI9kEYSCa4zUQC7ufUbPsJ
kgbX7ySSz6cF6s5tg0dYVlk0CL4lOVRsLgG2ThIpIAL5cmUXPKnJm43Vt1b/DKgPr0/JAHvOAxXc
LXTbYrwPearEqodZ6NDrQwC8xLlsSfSS5mqD7Cj9oZfmbNu0pPz3VtvbYM1mdpNV5qHtjSLsmmqB
zsZzpt3xgVA9DBkxKr+bcsHgicDbQUAPUvvAyNvySa/nMeJYnVx2z/ekcBI8ZaqQ1TtaRvDNv3hJ
xbKaTYrbB/bX3InRbL6VIj8FHINcqk/VhSTKDe/sKfsPVAnrrqnxVc4TlZgCsD5xEEjIHeZk/lUj
dJg+RHrtIeZurt4FSI5J9khsJC2Coh57fc5zkh2nz0Ew2CzbItkzi7qy5/8n1gFRSW0ymEcYJgeb
S8JKP2aEpXhurG3485xQd1W4fn+VyeVSjQLoHmzrcKCVthEYwv74PLqMBeZ+/zvvoa7xL+vWQ3+k
iW/YWx8yW+UULLmNqH5+7JhiVxWmEVhpdvzA4XUt88qnig5BPY1s7ResQ1KGpOmZwFPyjocGEIU0
DxP1J6MWZFvTNWHXIFNxLvZsaDEsW+/WSPEyGOkKyaOGslq51bpzwKfZA06syp0XLFvNuc7+TJ9b
mP/2Yedq8NfyGaCBmDWkhlVnhoknbROdD1921v1bSGZouRFDP7JuKf//EWIJlXBCZqGFNnCuBSAX
+jhSh3DEEnIN8qeBJ7132A6ycfeLeCrqOcaNl+j5o2q39cmNaziBZ7m0bsvjbTW4/WUIpOwv+yLS
SR22b7du2S16Py81WIfdF/n4FMpg2Wr6vyl+JPQuhRUBCBFr7bKgEhGPJ+MaEscZqM141u/ViEA7
GBJ2qkvViO+e/iz9gZDWbdJO/OT19diBcv4Kr8ZrMMlM8Hoj+GMq5GXA0jVfOzBUDpi+sWkTfsTQ
+x0Cnps0ncTyad7kBEMmoygX9i71o9X4T6j9NLz4qvh8agGtRDxxuQ/DBc29/QIIT6V9N5T7eYsP
1YyWLRhPDsZxM50r1qgaLGd087Rj4rHHDNGhd4SelJvghmt4jp72nqBVpC7a2KjcoEQiKRsbeqdY
cm4oq/1D3PEF9wsAxzFyuxyFMVNeF4jiLyTBxEwnT92vXOE6QX72TcCusib0dzYYPAPc0qvF+7sW
5BOF5fkDdoEc3mEu/vodc4mYfCBhdBlChjvbH1huP0us1oqV5uh22LkTP0EoH1wRUv9p7NSoMu/X
T3d5OsWsUuOKY+8obnUQ8zbsUmGgtbyCugYjuVpWiJI5jzu/pRXyUj+OtEIUTLoXzHXLwKxe39iP
/WHBcM71C50L4Ci0OaBXX4oO/4VDsVJeEqxcvq0z6ShEM5dpp6fnCvS7e+IMncnz1CZ3cG2qr2ri
hyQ1PIJn4/LAmPi8M+dFxrSsZq5yn2yXqetAgnyJytWEl+x7zJpFuqIYnpn/1jZHosWB7skCltTu
oUocp518eUv1j4YT8UC9F9JAgAQ65/XpbFYrXC0BB4cH/1gFgxD9QX4KPfh9IqqhpFCr0DYp0NIJ
OxmNd5i6TMSguVKUlLy/Z1YF0N0FjjPGyFBg6kflcbA0ISIC9vqVbB75gm+nCwyukXCmzz1ORD6f
cESL6ISiyPon9Chg8eY4Ah6ezldByy6kiw82Rviln/B9gJ2Ov2BoLAQCJ6ARzX9Xe5ilLOEkAcrd
kYT8jtvraw2lGbi0kwAdtO72wHjNbHRdjfsvdOa2wXdYGy0xYQ/NZ7lYzkbpN6ghuWI1OswsLimE
o6vxB/iXhKT6PZBeXOb296jlKCmcVFpYDmp00vLbBv0oFaoK7g7yQgq9FtnmIyaptKFbEHqQG1Vu
GTiL2fUO+CYvSX1VervykKjT2qDAqniYulxImP1JmromI3IuiNxNG14RufA5/Xd1I/Yqrw9ztgBU
CpsOvt4kWWg4ZqfPq4fuF0fInpy7ThbuJtYuVa2uFU5C3O9j/bdTBtzrnu0zo8bxLMvaI4Ml6T0R
Aro9Lj8GUQOJKJ3RCnrXBl/l8EDlB/4gVBUqksm24h0Kr9gkrKnA9/Ah3lRUGKbVSZzWgpdNCo1l
W/kh0geSMr1hQ17c+ZTu5oH01j194PiyH9CC9GjYztMRS0cporaZ3Cb0vUbpYKdntxi1MATGpZOZ
IilemMJVZR5Spa6AeVtDP/jjAoY/vGA6lUVUG9Hh34i4PEWVn1ZMgleegbdBW3F4mqdc5vcQKkE8
iuLc49bkG6f5i0uw87GwKA9XnrSRJVphJThKJK3If2Q2BxIs5mAvcSyIbCwYYmQ64ylS1uUeCjRE
9C8y6cdPYru7C0IXqjVA4nMpHZ316gLn57gKLvtu1KI3eg2DcDseJQ1ZtomJQJpnigv1H9OPYBHy
Y/L2+0cNMmWk4ZZsNZbCxIXMZAJCT+uJwrmalJquiM+lQ+QHVH7LZoGFND0fgvf8XxCrV7v1nY9C
v1jgdzNBcsXpEywLg+Od2E/bxIE/a/rhQuuYNExcIJObjPYOBnM08x4vfkM0jnJ322PXawf8nrSG
/AYWC4LQnkCIipWGEOMPCWxrewpd9/yXY/zKEuqZzDVgxyj0JxXpos2142CJrbUsXve4ygw6iaD4
VrheC/Nq02gEjpI4c9sAuYSlBQqGZKgXOxpuS8RrrNUysOLx57zL494/BtADPop6gumYW7bDt1gG
QSr8oFa+lwG6tiTTqD3F5ygHHvs/o1T/ZPtX6c4isUt46flKZUWYmlsqmakz9pDkYVnInXlK0az2
bHk2Ch131d2/Bh+Z4HydFG+LA38hZlSMViIzAcEZQdHDu6QYIA+M+SkXQZCxgF3dXjE8Sx4JR5Oj
K7IK96hUjM1IxH/UJ8kJc4cim7UalOif7E9r+27HF+0HGJ4GubuXObx2cseKFVKnf3VpsIF95bO9
X/4kL84zRNuZEcDQthOghMnwBl83+C6WcM+4yRJH7rDgCWWqCR5sO5W3ForpuIGrFfzCTyuA8HRC
iISuUCfLl9P5+RbNQ8Wsj3Xl4lZ9XlGvNFHpz7IWFP5UFGQDOU8/wERtGxngy0VWqnsjqPiZrOlB
9Z8BlcI3xQ7SoIkYBdqVr4nk6WTbTQsokw7dBq378oOTmOh2jxFIYgzmgMM0MR0tPPJyYIlS6tD7
Wvd+kjbD1+OtcKBo0s+i8KrAit7qKe0iK8E9TJvc2+da96ztnmgEj2ff5FQQunqVJ2dwV1UPMFwC
wm9Bl94SeG0Y8VGn84hxEOdNuyifUIJUBChc+Bln3hkyRwYniGJDAKWhlaU5EVQr3xxkWNb7wmVl
lZcC6+MQIeeE7zgDqjTO0C/PVsZlsBW5zYXClXRVstzrH+BhqlqCPRRO3o65zbISbi1V17khsN0r
rBE+2qXjLxTu1EKzSX8jK38z74aaFwHrIXrv81qHo+ttK6wCmS1V6EHwTgHzpTdMyS6h/HRxaiLE
tHTtGufy7Vtxdr8gMt75MDUfGCXmCapdFe29TtiAzIhmcTL2pQ/feE/psVvBHmJPEuc4oZhPj1NZ
RWaqT1zZMVGzU0FBx6skzRMz8dM3EX2sgjuWJvp2mQqKkaXnXcH5Sq6TYtwW8C2tPqUUMCY/Zf5W
oYgm0dNu8OolFi6BM4kFC3w6CCfRxLM/F77suZ7cM04/h3kSCF74y3I6MIYHcX5eNjFgQKokI6UX
OoBMWnnpbQAt03LmNrVLnRIVEHek6IE+CAnzXXvz5m7F/c26d2ryumgdiUov2qkHugRx2ogIwSl5
k6T6sNbp0PuJNre+s/YFUGL/3gb5ul4bqqo0o4lUrcqE8clcd1c00rX/MmY8gAkwAGzahsh6urfz
5nkzv8EJv4+S4lFwZjNsSRka0fzDZMas4zx4vFB2Peb2ePUMrtP/V7IKvi63rx9imkXvuC3LVDY0
GAufwpTnAbHgvZAHzHSbtP9T2d4Djs4dcnr3sIB9wFFOuKJ9dYNu2uzGdKIh/3i8t1/z6qy7DaIO
tMs/y0fpQSGJpdErekBQIfLtWRull3cmFE0f4DR6xFoWU6HghVmNIf9Av7N3mbAp21Y4hGln/U3M
sPVcOMhMN1uRZzEYLjPFONua2KE3PaduG/fSv6lzdY9fbKXYVt704aSM1zDVueWvJQC2oG4q9fKQ
xM/3Fo/RHm884ntrHGW7qGtN3U+41IiWV9bvViP9d6uQIAHJbbTQEfr17o7lj+nzfZdS/lZcsOub
Nj5/FYMJKY0XO9hfBHHSVOHNdpTU2WQTCKgraSgzZRC+9mdD2aZtUOzMftmnmkJ8+1OZy/TnRDRW
df6UydQ/vukDZLoDPT8/XpfrtL9gFxpiJ9XyqMHh/jpnr/CNklDI+AdsULtWjnY2oWGzGGdMNXu3
19Z8Le1cldUK88WjECpqTK+VXld4lT6E5ij5e9pUJHUk8ipdO2lK810o3aslH9bbMvy/dV6yNH+5
XkH6C9D9Xu0U7+BrPkNN76cokggfMy0tnglNmtugF222M4tB456sj9cRsihi+orwE2Qbw2J7L5W7
5PK9cgM0gGc6yJaW7/XJVa3QyWXlaO5wWa4Jz60L5BPpkNaeLx9CjDG/gwY1/8GFmbJw8WFLm/UP
4cF5CXv7A025BsGGKH58gLc4zgRRmSNrzw7zdNaH3ko/Y1BvXpmqTdl/q8Ckj0bNPuPOSgGjeQS9
OpXJLZ5kVzMs4HFJhx8JI/GFp6RT3LPzzVnQ8wLqCfXmijTAiZjykGZ2HNK6Er0W6OdaJBLWMn7E
eAABSc4rEhDlUB6M6kd/ji8eu9zWsno0oTQisJCJM4rxhGU6egsxm4jPwWe7YJ4jIa8/wf3woFaw
+t6B4hgy0u3+26U2DcJEJ/gi0lkCw1RugAoZfAMcpnpI1BYfUnJpEQf1KprTRsmt/pKy9qYEOONn
XiDRRrL2wt2lrvRFx2fuEcmWnar73SbTKgsFTKR2Gz4MmFhL0J9SApvAabCivlIjuTEvae6mrBQH
bPgPdEMCd+TVWQiJYyHNz1DLn4aJ27WL+PrUshla8H7qw9c7dnGAIA+gCxKA8ipDRNOFfAF7yWC/
wWfj4G53+nHI2nIVea+c31hErw3t1J2QxH15EJd6l983cta2j7Ek6BItY3hXtpgQEA6OvsEyc7gU
VZF5VXBdVDJLZAWZwI0LOwfyXcyQ7v/pNwVIf7dVYWx+H6x9/O1sOQhREaliw5Sy2Y2wHsqmjy3S
wXItTWULt7LCQAISc6IDyRkVp2eaH8uoJf1wlFpbOm5ALiQyNw7Zu8hA9d3OHSZmzY5omPjZui03
NOH5w9b9z0UQLrf7YZeJ+1dOJFfAD1gw4WDS3hsfei195ycWU+6Gg436xRvMCEUjM7tt9NiCz3X6
EhKRmX0GeQh0+/pRZ6S9HdG1q9HIjCH+ivtCCWOSGKNbBJLW0DFviYLHdTgIYLoedq+X0T2jT4gl
IuuS7DZePtsH+8yNvmx4ksjajFvWc5xXbPoRqS2WnYal4d+1nmKXgQsZT8sQ/OVLmyut7mNmtqAT
+sEXiWxJNyGzWmwZN3u+YFmjy12ea/oN/83qarc+E9CnNJ0YLuq8GKOkuQCz34sWc1qKztkC8NVR
iIci8+bShKbEj1TfWhApJtBj3ylrT85cAsBNwugz7Lk413OlxMcNAiCJuTalHGNsX+3wmiBvpggp
778nBr0E81zhrzf5FKxmEp30sBodBTEdcnmeVNmH6QAqWYq4Bt0kLpg3OcWjxKDe0+9zgVa4dWg6
y2P51YW7LM/hzGj5au5kZKZ8kjX08JRHhqvr/YYLk9MN4OUISRj2jEj6D5PXKYIlO4gntaltFsHi
XIoxGoBok0GjAP8u1TPgsF4fjMManzQJXuR4cGnEFv+hBsfRIMKUdxsMCRHku1HgdtJuulG1hSUz
jiDN8i0QCpcrP2SdrbeK5bYwCPJS96QGF61bp4m9M/Y+ozxSQYosT1AH0c2Jg5beZClQcQqZxeED
G3ED9GD1BmXYsJCVIptgV32FPqRpY3oKaBGx6gPV7MMduXolDskezZolpevs098X/s1waVwYgRLe
gleIcwXPnQ5vKwyD1MkCfwYzPkkQj0TiQUZRyGGCzGdp52aMkncjdf5lEeTrhw/l9nHsG7Bfl53p
SwOOOS92JGXM1xNw/rizBWHjmuvBa/3HNuIuss+x5kr7K8VyYPAeZafJXjOyYQruGZB+balvlYHX
Tq/oLfcYhN+7DGlWLb//v4lmjV4hBMXosL/AjENzqI1MIxtXEQOGQQerMqe4E69VPXn7gsyV2Ide
OrIxgc4sMrk4L78h5nAqDa6rGshA/NrwKRrw2MpB88x5pzIy6hOUfBlVAh9qd56p+QQlGIVDDUJY
QfftC59haAq9Xw+ILUpH3fknNREomg2yY20qY5+4OF1EHDpV1aqjNlWiUkXZPTL1zEdHhEy95D2n
477Ymqh/GIMQPwvAepstVaMA09C5xAL2Q9W6JXXy6Jq+2UeHQwCn7g/fb/Yub9em+xpt90yHpINZ
rGZWLApvUTy1SCqZN+VlyRbjy572X5SzI8Qqh7TkuTAeEl57loo+iQyx8rvmQJHVvMOXMp9X6lRx
w2YHQTDOLrNXiN5MLJOnnU68aEPWZcjbR4DEw62eg0rXhadxziWuuLhOaHAofwnNIcGlK4kcXaQE
ce8E/TNLiSq1PdRwYLe+ycvUZFPeK3zFtfvTNctOc1IwoXgyyx6zf4FlbuoNvXg8mH0HiaR1xSIg
i9G6vNNsTqS4oS7Gb/R7p/CFVLbs770l6HeRBEy3C2mdMKZ9PgCntejLiFwB7bp2dUhXItnOAYCs
CuFzzQSZWbqtFA2qG+pMtrJ6hoP0xe3tvUrX5o5mAOUzP/U3DezFMqhCxkU7d4/8g860lzI0wTPR
ojwZM+IXrEE14LEQf25pD/z84PVXATlb0a3hIdh8WdeKpS3NrGFcOiN/wdJ43qkFnFl9J+Sy5Xb+
SS5maVnmV3Fv1mUlO1ZX22Ov5Hpeppl++zNOuZjPFJOO7mmMy6FISXAuzEuPd3pxgCcN9awkzcxZ
B/8SDsQZ5MFqcWQltw/jZ9E/SEzvyYybWI5ZrNjmVSRhzhwA79X6iBeGpeTQMXQsDh+iPa4os3kF
3M37jDn2CraFNP9uu1eFtDatgrthSvkColCFwmsucXQhQx8iWvqS4VxNR5InlW6kLJ4DtFD+a57H
XOZuO2DJFRYLhue/2/5U2f/MS4Hwo+rwONrpdY8iqajMuM2ezhFekI/RlI6nBQz3klbm+S0SGwsP
YW+y4G7YNvy+Nq0J5wDEsBrnoZP/Jr8yhyMB/WmchaoeCi74+su8d5kpr+b++5KU2Yk9SP8+WxrJ
CiSx2Tan0gykMBlGQOXsR3XezaM9s8lJJva/rqU9QcXeDtaptulVCSO/6BhuTbb9BPfplnkf4/Us
j4oGmClaMxd/ycwzhPvtx4a2yjuwo8ACU8CSxiwitoOL8kY5qZKxDinM3GXduuZKZLlHmlYEz31p
u1pC2sOpTt0WtAr2tXWRFrmXcFSILJXJwvDoic6SAL2VJ7NXwZNFXjVDAoeCflMl4jrHYcGXuvLn
wfJW4B9U9uXWqBmo1HrnPYDpAcpHuR8peCsZb9M9A902TJj6ABI1q/z6GQQTB/2VrJRHt8I5SHx8
R75m2Rd5IvwTFHmIXGXESgI7GjQyEi533KyO5y8I+GNEV4XxwdNH6rbPi4DnBuhAtFF5FgAzhqE1
i17ZtEgr7a/PlDu5H/YXRCAxBbVemp7tDMiNYJmV+tgyvtCqTcz6CjyMM4zXvjAkPtVSJ98XPmzF
YM8L4ExS8NfXSJAC+H9nLz1kylwapI4DtTig2GR56lGxq9f0+AcF7YWh/q+EY3oCELH22d0T/JGT
XXKINzbxUpxBmpuPt566N/Mtd1yomrHgf5uZMywMzt6TLbPcoSJ0Fx09RG9rRYtcaVzPLx9sgGaQ
X8SdfJyiuda+vLilrudRJIPTfRbyKdKV83txrIKvUNqE7PUgAnonhL2vEXN75PfaXO7LOnm7MRv5
pHBUvKqO7Ue7TbCsZny3qWKrmXeIjvLEEzkikujLSuypbjWElqdbj7YvzhcgGQ/U7h5f5db/z1En
FKAVZYLlZhsw8r4OJpZoXWZ+98FXkwf6cVy22GTQLftt+yH3B4dXRMYsP7Lwbk3hD4tsYYUn8Scg
n/XbN+QNtW9L8bsEvxqo+iCx6l9VLJdPN7WwQRKfHLv8hZZ+NIJyVQMbYvfRspvu4IpvAHTgCMZV
qXSgQ/aUYwUkEoIz4ow4svGmQXjUdIVRrvHNkIVG1jhmlExsWNyGEnCXDlaEdTWP+CGzF2GeCX/0
BVF+w7H2vFJ6qOh2WSQNZD+6yDAMwBp7WCfEOLc3RIGbtW3gqWkN29eNzLzfXObfgfZIarQuJCUT
+FNLV8b078CTBhAtY4uf1pEU7uO2vXHaX/KjmKOGr99VmiTsYlaFpL3Yzrv1YfPpZXFn9wUtyOai
IaVx8xbddAjBCtuPpfrKRo2Dt2WQPFjPYoKvBOxl1stDxiTwvxmYLY1l6wFI/3aLOrULP7Hp79T4
TKXlOjm2cdRei4mei98kRcL0O8jdiH3MJaeGWU/9yI8hdHEEVp/XW6nEwx2uT97P025ZqfTHpHhm
V6OTcMFOXsdY3VkfQHBlDGglno1lcfSAGE/6PcUfr0NkZ0ZJzSFSpFr/GKKtuzZ3ctp4kNUUGkPL
7/Ulc95OnXmBTE8ynvCzUbGQRBEeVgsoNZn4SPuKqlceoq2RQOgGiutvLMmRoH2zZ4/ulDOyCgOE
j9x098moW2rBHRewbXe3GiZzm10ytAW2Jc2ahnjnRUKJhoz7As78zO+6UaRyiwA1YW+cPMHlUiyw
kk/AWcs39amfmPmPyDRSiX7ldGz9cyfmCRi66Hiz6WIaBGY6Pb3caa3GZUlOPk0UlsROV719R3Rr
9f7gPLklT1TCIZcOnggXqVs2F4BkwcD58oWGEIGgD/LQout1QIiteKEuERBfRU35fg4VeVwny99K
hGcnF+Ws4s4rxF46RejmS2ClenLdOgdrSUkS1V8kc0chSeqRIiYyCO7ZDI4evpTpr7NUV6vNX8bB
OyD9gFEhmQ2y4uihcsOTbvj8ZGyHyJfhJdYpP+U/4JUKtgJyYdOu6BybtyBYnWFnVbtvuaiVzucJ
h46NZ4ACGSNrXWeqm1kPJ+qqVT8nUQQ/m4OhAtn1X9LKhmUIX90rNRaWLn8txi1em1mVAPfGaNF1
6XniHlBgq4EEhOiK+DoSrDapxgkO6K4kjzrqp+YjYa8tG7aE5pmWLhwsUqOlPFoDs/AVa1fq9Unv
insfAgr1WvoyobkGHg8U7O9xvm0cxiO8bZSGGacnkhLxJcNRMoPCydqplHjY7+5KqJitdmx1kI+b
vPuT1nnOy21ecTwfpW0prIzGq8s8ogXyQa6EhmLkD5GrfDw1xcicYSKXEWA5tHRB+9nm+4lNWKOj
kLHWydOFBffk2oLhTgW1SSNkTAYiw0rzbyACRcy+CFJJNqksEv2tAtWQP58GW4KA4cEyDd+J354r
JD6raUvj/Ud7inQL+64R3eIuuaHnQwvVxkYRCafpxPKG1j6JYQa2MuEbLYjwuTGq8aBOjHFueiKG
HUmIGwJZwfzXB522dbFa6FbaJ8gNqePH0r2h6QmCfMyj9xxerevBD3oqZdbKf1Atx1BJUrwjb8rk
kgnXcL5kalHYARD4JtmSOxNfxxaiHbkMXbR6Y0cNHba59fnnHpI98vdI1wXb2Ac/bSLechKcguKO
1nbgyWYiNI5de/2CMWAmdH/U4UuvgO4SRNhSSuJBIzwDeZpLD2bMpuvVnuduvLoJEwKpASs7BJY2
QdniPA5KHqNJ8NRJb/7OimFBOYy0wg35ZCoyHgOh8r5ZhS6mmE8DYtDo+aanBbmUX+9oMXya43fL
yXcySJfjINl08oYzNMXIHq67mGsH4FDZzcRjIQ7IXS3VJ7rSTR4wiqJjqXBb0Bj8uqDg2Ygyg3bc
ZmMEzHwvBS1VpIUgZ+eY4zcj68Eg2ZDYGJPgk7qV8ZIFFQ7P06hI7HkjHMhC7LNs/JawDGyj/x4j
Qk3QK7CqQNg487SIfwiF1xwsqTZ1eNf1BC1LG5AmGnzuPu0VoYTpb3ckUBT+hLpi8C7udgS2rukc
3e+6j/tNyLVIPoipAJxZB7CM+t7ep9kQPwB1kI/qW1BvKd4kDYX8e4J+h57oeMfEV+cxrGG37Ehb
0YfI+shIL0lreChvrlRHwZlkrwble5rK1GLVmpbvobqwmN8/TXjktxRQPdvPWBzknF6jlvnoJshP
FYvB79QYo398eK535AkkzFFwkHkXn+nhlxn922josVcabttstmY+TPYurNXwjmRda972zqMD6Bjs
02rnyWt0XfhQbpW8Vy9oHukxJx/qa8bPOs3zzDM2SxOqaHd2eJrpPcZD7Fj2sOxQI3PkgZ1Z5l1Y
m8kyoEW6sENezvLmueiYdbPhTSUZS/CKq7UhgnnUzq2gttbNkdrl0XhFUrnA3oXgxylsO9o04SxN
v8a8Ol2Zhx8ijtTh+tyxskE59/HCSKLRhHlkpQXfzVGVso5QYt/x2FJcPMWGYtJKQ5s7IWl8jUXw
x/hSElsJaaBKb8tFJan24r5TAwzrw+8rBKR2z3IcBt/y52fU2PU89qsdxN2pv55q0McFOI/pnEeB
85VPIgx5Gqu/BY3e9sDIjKM8i5wUygLz/Dm5ezpXvx+9kUDECUqpHsFk90UHxYAEiovl964fKK/A
Cg2LekHezwXmwDduVGH2+wogsH+sRcflkMkn6cH7wOHEV2K25HwU41AE0J8MN3/Yqkjnt/RcLirZ
drGzONVR3DBLYO1n6LKpTsmNDcF2B8vDxZgcOKZqfwAFdc/upiC5cnJCjNCNoG001gfQnRC46h0U
i5zDCH16viPv9fZzhApuH/TUHYYV+LnVxmqtyTSzWIk6+eMg5i0jrIWEUSPG8oxV73IjaGAm7Qx3
ovBjwR9kYK9yduguIbBbo3ELutd6+NGKMY1LcKHGVVKu4R68fzzWVYb74xSr25zX6Qpee2OpEnBK
xQ8JVxZJBzUDREuNRjzRjjbSknmo9IzemRT0q2wEM9jbkxelh8q8LB8FE6ZlWHvYJFVwg+cw8K/m
TYENrmFTqMxMDFJ2IMHbKZtVuMgvjadPq0YOGSYHxUF36NRc61aJrSdlHvAs8cGSPRXzextc5vaP
MGAofjBrppfiNRnZ9KFE9H/pxUmj/DL3oWhR7ij+7p6qa94mpb6Sglj8D9ugGyZsf62Em/fsu4fn
gMFjWyPBSkrwBCjWtrTxX6HB/24Lw6soLjMrJQA0HWaBaAmWl4o6miS4kERXdC+IoFSWH9W6cqIm
8rovrpJU1iFx2KZdEOFGNuVP3myOoGzrn7S86l39DHwLm+vxdC0EmalHfPBGW7T+78/W/sFDukSx
bzcvtisSGZwZH0zEnBlvBkrDVsNigdqOA2iPRVGlh6dLHUBWzIV5DtaSGzMkt2E9MjfcIVzVBZOu
Kc6LE2RWRoPWA8f8UdHRr4rQdQezEX+HwPgMBO5L/L1nP9fNWByjChVfH64ypKF6tVLfDpPtmgRU
V4vZOlY+cCcfMWjAo45d8Bz43piU0mgaLzRbvsu0AJb1zeS5bOuG+4UHifVhjPDpQ6DtQyyXP4Gx
4uNXp0hoIDNkK49H5EkuZ5AFoV/3dFjiiReWXrI68PA+aTVfSHLmqPTrtUizsMLNRPw1mIBH8Tgc
oB5PK+lu5/hZn5txaT7w3zRibRw3aontL9OY6/V9yB1HVS9zvAJQ2GU1oj0/uowyOMK5kNN8YVFi
QA4iP7Ps03pUMAL/DWmYXIxFu7qC29UhdnPOKgggUqROQLHR4gvBA7DojXni4UMd3HL9kfTj+Q8m
ExwaInmGRgQqIk5hk4ps2MeNDfJ9j79FAXRVnGkaD2YugzXfnZswCTNzPkV5xJVOSWOJjWEBwPe/
MchHzsWJr80ZceMzypchC7cyMUAPESDIVmE4kwvi+oiFerGR9Ph/oKVSKlsSoLxTlegd/UMVNvym
bnqlhiWjBLv1C6KCz6B3mo91/HEdo4g5sySlAuU2LSNM18k2fZFCGAiULOFg+Yb6or9Hhsim1wpQ
X7ZVXYu1Rv4TwkezI+0YIGvSc3TH54F65sImxenX3OzD/txUdFnl3LdyDByxjXWUWRiY4ija7eC8
3/rX64nxIDvPlEGlp/7T6qF52+s58DP9nV1gslVm2MZCpTLZSDHAMM/P9SxaiZFnUti0OoS0XQQ8
1XTa5CnsxpZ4GzO20xj7DiHnBMKBt7vf7l6kGivVyOy6CQM7gFjJ6p5XWEPiWXxypDvK1ybpRG0R
GhS1oktNXSbkG8gVFshoqKowSUr1O/+RMoXuE8hQcfXrFwciH/ilC0sMBmkBqqrDqC5NOBW0HM0i
c/Du+wDwuhFLLae5znS4m8OXcLUhPKt4IyS29KxVBPngSlmGI1Kbjhu253wXiYUQGYFA20DDP5GO
T973IMVjjO8hVCfuywdO8BSdNS4q1/0oNzhxktcCLJTUlh7PGpFWbzCEpQ6/YZ8CgZ5qXll+nmKq
7sMWluwM50a0smf0M0wVnyQ4pfL5wLrS+XEQLHlLWYqrtIGoWK4Gzjc54Iqc+NZ1RXBhsqnTO70T
yMRCnVp6AXs2vfDzrKFDAHdeHvW0P51pNRgHVCSi+37fRfE2R7Rzo4EojXHEbrjsN+qzHjtcNchm
XS5Ew7NVjnjusL4kRiY/p4Os+ECpI3H9GImAjdHx6p9DbKr76bCC4juGgo7z2N+xZGqF4qui2agD
rxnTurtj1mKr6jwsaOzSuiX7hgOs55uaBwdvF4Pnj71DbVkJ77t9L8THn9nOreULfQi8JJeUvFNM
FK2wJDyeqRe5cppzsC8g1/7hmxSqLWrOtiD/xaoOBJNNVIO54G+nDeFmSNYgEwldK1RicRN/mAd3
vkLBZO0RMOkrDMzv5cugowYHI+EBSJ/uYgIcer9s7VkUnAHd0xxZTRQmuleWfqkadrzX+lAjIue6
O4qiplBxKYXwplzG+eWCZXPqVI9zssS1xonrNrCDkkbToxYbrf6k1UZAlYZifjupCLh/KMeKhGFI
Uj1X2Uc0cpjWEOt0DMevOrItp/J6Z5kAwu2lHTGjEyxXCtNfT1VHuT2nc5TJ2RqnTuDkmCcXK5/z
hRsKEmkLsoRdTcHrvzRL2kJBln+eEi2Bob6RVfvKFhUfIT94b9yccHJevVfG9wF4MXAZAsATOfKj
7uCykuPZmOcAz+sB2Mh+rjKCSkqZh8n5rwBT8npFRRIrnPgRdm8HgymaRZSy6KsV3cj7V8QJUvdU
eg813M4Sppue/hb1dvam7H7r7vKsOeR+I2Rv44czIzYiifDZ5s1Zopl5m35nQi5LK2uUL9mlXM2A
3P5UMR3GO/j2W6j3U0Dwq6l5dDOuoJB0yvqBdlizeGypvJBwEgLsF3e3gCMR8eS5BAuvW13bHqSl
rETux61PdgJ+vnABUooNK7qb02XqwzR/EiBaFL3s/ykDh9CPWEyORJHgP/CN2rPLOPKdXE3mCPc9
Fmjk+K08g3QJYzeH8ilpD19wWPCeKOij5nEGzgehZOUR3oYknjupRT1zD2tWOu1A0exotm3VcQEe
u4iP6eMRkxvaA0bJGLcaegkgMce+nrWKPVp1YOTjlSQLHU75jdrSHQiNSOZEm8ud7lTyOOv3tsS0
1wbDPC9TEO751YvETGMefVZIUr0DMLc5h9kGE7GdC1Z1Vif+FcDEoz4BZAkh6NchQBpVWVP5N3xz
XnodGzA0ZVAaORjABJ4o9hHGyx5Hj/b3aXSeoFlfYGngm+s/BX0ZwoK8Aev7k9+0laLwtQz8BqPG
pnq9dntNoExinEM0rDt9SCeIJ0ozQNpc2xiZqqhJHgPdJ9kscKYCHiJ6E0oVZRzaDYXwdW9XBXpn
0buguA0Ci0NgDQYBvqIOWmnNoOc6kCnlyWhJ4EgUXGMJ8RYLaj6kqhAdGL2kkws0MheOSXZcfn24
xxGgxlpoNbMzUBhsfy6bgkSGytsDs2wYcFSRxA3whte0USO2L98noH0pWqBLb1FY6yiYm6hJNIMj
AJJU2zsd5zKrzu9MtpuOhD3ta1Fk/8WsXR5mITbbdUbGgHOXGsnY9X2pJJGQplXx+/+OOotQE2rL
mo4Fc5gZcFr9FLWd/b41IXe3oNt1WywxMHEUQHDYEGdPXzJ+X2FZljSK6p4jjphHqd7hmccKOZ9W
LNPKPWMZUQ+X7s6NYeku4PL+5N1shl+YBJ4MEUA5tmb/P0Ela5KlZUEq4IIEBBawWEDIAiyMcMog
kAAx4C05upgC1rj77c1YS66RQkWqMnCAgKue5bcpMucFNprubIbDvm1OziHAHdFlWSZI/rGa3WSi
tAmPPIeK5gYmyRjnBos4YwQWT5rZmTn4LvrphyYjaBjD74L52ubqCmkuURBfPRLG54+xRYkRuXLV
KkKk9q7vAYMCM5J8VTcPHm7eKhCFdHu62geajvN4UbkZIvAZK2chcPzd98gfWPWojDSEkNnVLajv
fvnOKsYSwTaJvnz84rEeYf1ppNu+nbk48W7I4I8m/jPZk3v5hMtRTKEHW4Di31oxI32COw2tJ1iF
QwIKdNbEvoWtKLIVD89WfFUkMkz9fEMAyL1H1iCZLmByxt09zQGAx/fbKqK/XpOOEX1D9j9abiA5
QphK96ttWdaVy1nnmF+fuLeFJVUVBeViZMmg7vdNo6k2wgRDoBCxw2cNvarcdXhfDaQT5kNFxQ8w
9i2ZPJiVwezfqusQYjPOjz6jIBaqhfhYIoFGfN+TTM7yVPaOO8ZqxsLwmvxNPI2ULY4aamzqMWFM
PuV3y2SWjkEtynjA7IH3M4QUEI8BKMjIaVKs4HFcSa5Pmcz05fkV77IOplU6t7VlY3xlJvLuBpJ6
gW0BFXLyUuNqcvuQdBLzzsyUe1/QPVIf7G+NgaPUm58RZ61bTPVyPybwLjF3MEuq1RB1T66xBoXN
3VyspBzuZRglXKGZn8rsz8/JO/RsZm7sLOXWHMg7lvVSX9s3meTrTtJ62cw8tv7dDm8PPhABPiYM
/tUwPWCNZEDASwQjmwXrS9V5v2jHtw+ZOvupUZKXbYwWVWlITRRFUktO9/5SxLG/k6zssPqoMxal
qSwxql2gondzAEZrJ8Eqm39dVYc8dK05RefBnT8wqk3JWV+B9Om3VlGHmHVXrE2fRbxDtYceL6yM
oNTPRUByUXMk0dDmr76sF4cG2tjG+wkOzm2xD6k5aVyxezgSgpo9GpHd2Axk7EQrQy2ecqeh8Cle
upolhtsZRPnM5/OEYnAiDqu6xvnkGtArQJtVCXpUpJI5rybd54RChRiGZ7gDmQjE+iirLdW2mJ+u
O7AN3SVLUpgYoHLATqTGuOP/gd4scHbL66fD3qsaN+GjmjHLiubnX1s8prhX8VKYOVVu/b5P6KjK
9GveR4M1uvWqzmqJwtnPf2rPBt/CAZaSwfJOD3eCcC0+asmHDn19fnCvb5sL0p/q+c09Zjrb6jxt
qVPVGsPbdmgIw1O9Q/oVbVJ+tiQjaKh8kEKX44Vuq34G/E53W/YWWZFo21SUY5sWktxe/IYPI988
kxGbeE23PCwEbIhqxQL0ym2FKIWnJ1hMbF8E4neEBa4B1rEbNmGJbwbVj5RMCVjMMLSVQHQhIc2h
E4ET3fBx191kupeKZQwY9hqTe5NP2WR8foy8kf6OYjL/P7f3ES9wD2OIrWzxA0xASDJLpVNeWS88
FIlGDFIrldTw2gGgEVlb4AGOyxUWOSqpGGs7DsMko7V9Sy0TVf/krVJ2+2Gd2Y/Di+NxHFm+FYXl
FbCNHRxJGD15c3XnIPt7oMSDn7yTwPZMoxwGAIgcAJfTi+E74LnZVd/GHLob6T73VwVJfvezZobi
PDwn0MyiUcJsSBFq14ZnUhdkH//grPG3qRSnZl8I/kNclkKBbT2QwLZtcHDKn+sS+6LD1ce9a3qp
1B7UYHtWTiNibaoOga+xvI5T9ZL4rPdDzitsx34x8NAN4BNcNQJE/b038Xzgt/JnpoF828BvwEcY
Ip2qeIFS4lV0sqmeaTg4uAVpWhrh5sb/EVxSbDmRL3AhMXtwA5GkcuqpifAhdURoSr/VJ6W61aqP
Y+Hqo+INogQz+aCGg2YgXav5tXQw6bhOycQhdnxvU5hXk5FPFCe/jqJP+SKQqiyp1iBZYLxpUFG6
kR8jhUYC+ihg0EhuSVOElhFJhNm++k/B45f906G8HBDhfJuHDrQiynyCvQ1+ZIZegk58MiaT9aCB
UdfE1byMlmji0q31XXM+RSmRuK4kIC8wx/VgZftrxOVLt+RauMCpUb2XPcdD9O2W+5NlEJOChQMh
RBIcUmBa1kuzVbecu1N0+eJWbBNIvTUODHET8/bp1P6U8VlfQsKz/5VTBtJMFxmM9hjgbeOJQhVD
3zW6JiHYgIyXQ4wjKaWQihWEzexofQWbRD4xPC2352U4GHFRbfIPPYW/ehUZ9x8WKaV5Y3VdJVkE
r2hqomlX6yD14vmW8zjhTiKnIFXP1Re3zj6JyYO1hhYS0Z+6jq2DtYzy6RcZkOdbL4PdpU9+q5xE
wu+VHxYHy+fXpykprxXmPV7Y/bVE7F2TrxapFK4YMrFBmQK2Hbnnj7uaQ+iDhpjYFY88iLRgvi/y
l1K7SlHqT6DKEc3slSJAdc+79iLWqaH43le345kO9hh2ftl1Ry2nNsBHoBFWyAw6OLq4zlGx3LH1
BKXbgaEGQ9kDaq2td9i9PtJGzr3VA2/qoQLMqyuaawLB9WhAtd8Q/vYxNEGu5fB5D0zs8LxpETfq
ch8CUVYctEPFdLgZO0cTlcMjJW4kb+V/i3mCwTDwr//yKo7sP57/m7DPbJ3ydNvK7Fixlc95DCJN
xoAmsf6sC+qn9w9o0NKpXzLCOR1lUhVbyq+tswmKE3A6KDAyzPyYJ8Au/XY6EX0m6ZUcOxuGfE0o
mdI7828djAzhjcVEoWlAefDuwK5ORDdbCyJlXfhSbGElWN0W6kixKrlQkYCJOFxF3kLqojh2o0St
CCHSa9XgWuclG2lmpErfnJSgH/NBuWW+un3jGEflKJJKVsk9Lf/8UYqhWG8zqyWemmzxAoM3t4O3
3J/kNKaT4043yXO9kDlw4jgtsn8OENg9YTBAfOsms093j01ogAKbaz6zuv9eryHb9AJq0HVsEQJx
1xpHlGSVE6EbjHRH65S3q4CZbIm/nxv7GpUQ4V+FdglIPOSon8OWjMjjBND/E0nty0VncGt2Z6WN
MISZRKY4CBCf/KdPFJTH4Pgfrx2hefiJmOcMOphTe34xtiuOFe1WibtCo0XqcQZCpWb7WvPrKL70
9Wy1yxLOI6ZD6PcpRxwT0f91eDR/LU4BJlLOVgiuQpblc1279NwFvr+R8CTh11rUSIt8+Nany9cE
MdQ1hEC+3VWoUN5N/kysLuj2rJPJtwk9W6l0qaUb1hZDjlDdvAUUxtKMfsa/r4srLEPOPtqrrW+N
VUP+h7z+WBYDAUvcUvNrbQWw1kngDNei9Os45nVdWWez5jYda3e3cOj5XQCxBQ4Ihsv/AR+MTs3y
VM8naAGDxzlqf2EVaadlxiT/Sp7h0cAGjWDasZvNpX0ml9txlLrUDhyC9DepEMhzzoun7WZwLZZE
PIF+tGDjM6eLT3bVsdbAkEyY4qZNBm5I/EtossUjR0zZKDLBnBdp+4cCUPj7BSv7nlCOFupuMOgR
AcYgBajV56Gp+4c3Nzs4tyQamKfTUbhWu6OanO6JYzguEm9F2Q+lfO5jH4t7QbbOKgCuHIIy6LrW
2WZ/njrYm/tCCy+nAIHUR3fTdF8s4xcY5TREUEqX2mtRtCGqPlH14xJhUK9vsNRbwsI498bRH+L0
3Rp/78qBb8iaBAkwOECJNvbIh4kneqwBPkepi3SJikstD/koFI/a4vfrHHR0NpEIsfeSP9SYh2lX
qoSKFZc++4TVc+4NAUxBZt9GlzLcaF77sA80EOaFFtyU4Lq8lXPCO0Ffo37VzrofYWvs1gL+6KwF
tBCa442ZFbe2Ru/+37SG0rFGL1v7oDGk7nDzrNsYFYs3tPP816jeTRLwHt7wL4mB+kdVUSpQSBm2
9j9+vpC9tMRpr2xGfzMjDnV2RAIEfxq5bpkTnB7/rxyiMj1geRGqLQlNNTucMdmxzlgOYWYDWrbT
ERB0r8xyq0uRJJ4pIfUhl10bRgkZdy33Jd9NZ8M96i83N7nD+A9iZVTw3ewC3hluPDiWSYjWcSHS
QgKAx3gdFje8xQbibjRaUnAW+dexTtrtFoPUAm/CRqom+0tK+0xDHLrWMDvQi30kBrmIshy09xiL
ApNY28Y3dYY6OpBzpISH88C/3CQGhXNPscFc6jYHcjhYhsd/kBbUTvVycTRloNqC3wSId+lRLN5C
PqD4rAAYLdTKIa26qK9q9nuugpeEWZTEsRA+VR6zNL9xcJ4Ig9PDo/YAIihTA80DcZQLzCMBURDg
AQ3JLKovkwO/40d+NEoPb5zibXoXAbRYMJ8VuE/SCeksnlyHvTgKILfixk21vikmdZuRfF37JOMy
K/PZi4NhJD9buH7+WQwDwFzM+JB4lUNjLLsiQ4+6RuZ+taRLVcQlbj6UcfFVgizVoarFGiRtJwTx
8Abwy/hI0ycxJHVrZi3FTNBKZ6dBmWSuO5O/egWg3W582tDpuK+ApOD4awJ6VoOXjkmbbP/xwnwA
Fegz6xYiHBsix4wKFigAnljN04rnsCB8qfyS/QohAl+Ftjd+q0XqbFOBWYe+5Jmxc6xisJ+YmjoH
WVRzzAiogCogNnfbN7sAx06W6d565r6sSAbVuCqlp6GjmP5fjvuwf162kVrVdg5Nf6S9BRvjtTRT
HaxAvJYqnfQPxENS9BKhD9T38TlVOnGG7559EDG5xHDxp0jNu3zHMLSRHeCeV0+qiWKu4xzKfBVR
UsALSmCbLtpka1JjKIAyrOziqwEg1AN4YZMznbHtNJ2nxYwcicE9Wz44TvJusRWCq0xDqISORAOc
JQx3/XxYhcTHbxFpKBMjuLF1s1TzlIqVgDLaAENhl8gdwRBiFVRsEZgbIHhWFCFDL6FZe0CoaqXP
86NJaSKVn7LlyDLBYau9Q8pGyqb37UlYfwnQIsUk4t5UIZqlijJ1oRrx0SLp4clfIGJijq9SiRI6
rSGrtx26w4aEerC1RgxkzO4w8Y/TJ/Bc2yDjJk7cus2O8XC0ExGLOjFhZp7nVXX6DvxOZ8+EJ0Jy
kuG8T68ODqCe+TcNlqKltZ59HwEUTIQT2wZt5zJ0/w4Z0TEI9D5rxVMM8OwScNLqfy2wlMW8qbHp
gSQ/KU+SEsiLjKULCstrRBUtl6jP0Guimoa22FI0wg6ph58Leq8yPKPPlUArroM2PtOEERLnej/Z
DoeO9c7FAwCukxufwSp0OrhbtPboeGY2n9kVkTcYpGTaIT2XEiwGGZID8yvSsJjKA7x22UaVs8vM
lzCp4oLkfD57uhngLQfFDmOkk+t+29ltpsfGLaw+BwnYbfCI2sGQD3/bPmu6d5SASI+t3mwS1D2m
sQ0Hq5on5G2rMUYb160yF0s4x3GibFtqeDN/KPZfmZaKjNzSeKXwxOqDEkpd+gh7zCnxvwHiX+fz
k2vgi0L9DgLpbEGvNibNogg4GZCV90veHTZIj9XzCgXziCnP+yVPXRAAIIPBNCmMBD5+6FR0dRdX
6c0pnVRWehBmRTOa3hfOpje9OsNmc0gzGnrbsl6AYLJAxr6E42Sj1s7zfSy4MmdHobSGHOH/xYVr
J+vNHNN5ZfvrfUkL/VABNnDe85RNsxigqe7oQqSjUHR5wGumat4sw/+pdqDfFOGtumtlHYpjDM7B
2Kydt99ZvnYpAR16kR0Kca3iMfsyRfi9TOrUm/DKDsb4P9ruwPjGmkxgEkXVQwHyMOMxir3MkyXg
D+r5VtDTsfAn28nzGY7ca3RyFrGIbGH4F9UGnp6RloJIUbr8Inm/QvFAE6o8HyTyUJ2pOzJe0J+Z
7B/JSpuPFPrnVdnCFSa/USZidDMIKTnpVOWrhbodtFjJ27LaN2r770AqIH/YQFfC3L/xs0Pjb4oI
igkAje9SOJ0TU++ZZRHh5eGUQi5ikABpEZbiJKY2r0l63HJ1umHaQFLjTGIedmH1EAyrrBnlROAA
jC6yEs8PTSOin2zk4ZYHe0L5gwpy4sGLZL78TPco7gnXTSRQ5IJcD5IMoo2A37YPYdR5pWFpq39K
bLynOOwCV3BFbqJAUxEnDCKgal3W5l20YLTxj/Y1BudHHsvGUB1JU7/JBLwtxS3VKrph26WyzaBe
ktquN5lX0iRXsmTrp1lUwRPiqklFv8JlXVucZZ6+GVnL9G4E0bFQWtwBV22S+blZ6gaoOMwsVcwT
mEHV8eJoh4uZ4FkN2xE5vvd3W/aA6e4l1IE4Uvp+iY+gv9KKcGtdrxDE7aOfmN9/ON8BC3tB3izw
0aq/gXbBGabuNuUTZquzKrfLkqP9T+DfFyTYBL099GQb9vdi6eddcPUfBPORhNIig8R3Z7uFid6G
QNlw+KlqxvLJR7DZWjjevJaqXuUtRRN2LCUr5xHc76pJGqWl/RX5Vtt/mvvqsk7Must2c4Hc1Fmh
2QEtqhvudm1XSClX57nANHnVOe/kDKXDvBY3R4aeQ/lEoCFGkD4UrSuFj7BQ3jFD+jUyQGqXKHsT
zNjmahzTn57Y4/bgDsI6kl1lIBc6Qlakb6lNMntS0euTW8gIhsJiVJemWBUqD0idRLWfMPci81PQ
VKqCvVIkLZBi8MrrdWz0KFwFYuvZ+S1M+ArtOzH8S8Mli2/G2Rhd3oeq3sthXNIbX2DD7IHYDpNr
dMbUpGrLktVuvS8cvDwIXJNfvLMM7TQkCAqsihCEwp6XEWShNkfFSHQnLLWxgoa7N46ZmhKGgqO4
z+W1d0IhlS/GHRRihXMopztkq18sToXaq7k2/9aIe22lWHS0phfr7UZ6dUeYbWGvNJX+7zKGhkpB
QHDRg7c1T7UjxIhJd2pkQarHnU50qgHafUzqoHEXmwr89GlzuNk6NB3I9nqiJcu7qT2Hghzq+7T0
KeXFGq/47z5P2PFa7XFI3lpdh/2fiTWRro5cDebX5hFfJoBkR2Zh7KdVfLiiEwZyPSlZNPSCEAMF
UxzWlKGW0suBRF91lf//G4D/ZBJMK3adFz5Hq3mRWd5mnz3/6vC1oEWEJveQkUpK2hZphtMnzBqX
LkWRoULNwyPHB6x1Fq5r16pUKckmFub3MnjeLpDRFUscwFg1FVzgTFiCyLbTbbzpj0htRKj8x5mI
V0In3G3VAuAVysA6JpQXuSHlfJLLxtOUp42ngfNdEs/xhbfNWAfl8vDHhZTuXYjRFYWD+rumOx6y
OH4yW2eDfC0QmLPRZxapc9aTND7+VDQfmNrW5z/l5KPu28FLD9bnS4Td6BNgfBwXxHIwAmI5jq3w
QV/mFHSm+UmG7trF7kXeqmrtqSCPNs8Aukbc8DATCEkHk3d3KMSHFfWC1WUp0IGF47Tf4jojYB7+
TFc+u3OKnwKMZrxSX/4WHs7HJOuNg7axFtFCI4V2ehHc1ndD8kaaUeTcmeCe5vVNkvIsN3uCj6h/
Af4AI+ZQfda+9zojEnO2G5bIKelLhKjWBnwxsAOumJhkuSlIiq5lHLvBbsN2OlCV+6ILwYtzxFgc
eaFC4Skxjco8vQGgMvrKYHQ/uDw6Uxl2Hc4WprNsuEUFfz7jPQBxiRDJ88bFeeFkZpFVLl43qIya
6mn8SQKw2ZuiJYYTNdfEX+3o0W8tcvdP8JYl83IOOkQz7WSLlNzvBddvloNbLhlo/Il0KyIyMbE4
8bfMsQBUg+YyxNmxrSqdek7Ihw+BPzNmqyzHuKeqqLgm82bjdNPd6JOXEb2c0s8VozuuL2xsIuJ2
dtfkdulf8mFMwvwoQIvlVV1YqxGpNeol/cBQHt59giqGgJoaU8SNArErYQD7Yxv1bWmHN9q3JaIj
Wugnf6qkp/pWZ7VP85SSsG+K1zIJB0TVjlTPhIybGouhjODrJFEPK+0Nwi4DiEfKp83ja6wcbBkh
eiE+NXUXXMYGP31z30bB7J1McgJSXxzhb5Dr45gEzltqEV7lvODyvZcXe0d+epGbY75uVCvqiWwg
SDK7A/HlRDxgGhyYhxKWoYGqEwoBLirqeH1Ig3s9113VeoJ5acXjT9mWK8/yStJr4qeKUmrD2VJU
pE5RwLjFHMiv1Zt5VKbz6gXhJBlR2Dln+XKH4Z0K5H1mvUe1D3AiiREjjIOued2yhnKitKmwBSSR
t+pCzFN6OdZZ1l2KsTxSz98msDmnCScgqSE6daJiByoiNGPa6Pl10cuWyTUnzAbiU5YSR37fAWjL
V089ABcb0PNAX3GO+W5JIHaFp3d4D449rh313Rfr5zE2voYv2V5ZTv3vIs5yUGK0SugSUbaoOoft
ioYohUJhgE/C79AZnW+k0jRNp0sSZqycwAdAymEvWQLCqMAd+al7l/8VR+87fcToU6jC5x+qpqcQ
hzPnRg7ufoad/YOzzn9Qj5Kj9mwdcBNMO4SJ943YqyC5o/sjfoiJWttlqZ+vyzGOx9rEx6wkLCkg
+USWFG09zvkywI55na2Pd3pBnWhA6m08RzlmobMrlULedhgZ9SLS1tM16JzE8O55jtxgnAKNsuQP
kbs8cwZ1BMCTVQaR2W+enMZaXbfp2WE3QW++6QRpv2Sr9BR+EIDscjTeQbQ4zGHJCZMAq58SxTmx
uKfNxrV8nsmevFIKP9CIy7gVnpHEOVkU6cvmE4d862ROCPI6BX9eBCqRrtAJvvkMxUsO9CSLN0l8
fwX/ZrmpzbkXRZTUWVAuBXMCzvKyzOhWDYVUDrPsFFX2uzCaND9f+8bXqcZm0OTxp5GI0qZKJv+w
pUl5BMd75R6aqCstu1MOO+oYAJ1/7tqz8gI1s3KU+ZQ6xzbZ8vnf+ViJ8tXKvrEu531ERnRWx5pG
QuiaM73aLMv/9jOzNwiYrscHWrQ1yYvDOYAtFjGzXzMKl/VBEH+FVuJbqWWJglFC6/qwZLkxvV+n
bIDRaiUGyj7+GU3jYKKcxAi13b2KRZYiTRkafDcHb8CNRchFvqcx5zy/ZVosHfUc4TMBW/OS/K9u
n7HlmCvXAjFXezSKmQTVJHDPz2cpykNwFlBQAq63qEIq0syxBtC+OEFTO8YbdyoCWkPzQv47bvK3
4w4wMUUUkWBWn3kaL0EfWvwkJECQj0iJVhFH6BKY45ORIW7X41fGhssRHHRE7LhRXOSXtBuVE1JR
3MeTmCOEv335JZWMW3zEkxVw43t6nxoid7U7HTIXbInnS91wTI7bbm9q3x+vxc7RnsRutaq26ajq
Do5jNAoofYywRoVJ5fF+vH8dhgpteFzdmEQTXOOw+QrG1aBxwCyvNGXjuOffkfQsvqw0PS284inL
5fV35cjXOi8ILiT4yNyEt3SKAYytXXg/5losrVuTU3bLnlsP3UVOXZvKJ8YOdN8qx6JHDmes60+0
RjSKDrlaiaXC8o6iBsHi7or/jOJOsjr2JaZR0RMkMMRGXUWalUDtGqlEBGKU0sw941Byoa/J/GBQ
hKI3RmPDXiDmc2ns+3UbeSEEcY5b/jJZnePvg8H6YajQ5tMFwEOEWoG9tt2PMLiFrb8bqsSSs8ZY
ZIOj9dl/p++zpuXJIwETby8ZMA2MPGyOSjYsaO5YzSlU0+N8rd4DZmTmgOxEN6BX0Qr0AhbOCXJM
sx7l+o7TQPAPuUqBuD3i+auCtAYi//recbBNIgs5i5p1YX7wjiUTXGmjJT17dfCgVrfOm+FP3ZyX
c491inJS/JCMBeCHTro59W3l+yLsUpLMywCZCOZi7JmlI7XKyqJ6p5chwQULlMj1oeIQ/IXnM+xb
ZoDjnNk4x2mDhUf2KgGnFFsIBylivPa0qR2t4tC1rbF/JxTgO2JbwIba7Q/ioxouEx0pe0IaLwWH
uFdXkjqsKBhE8SS2pIEHGGMYv/BAKlNqonwxP66GwXf3YRulcxJ9NPJM8TyLIhD1v20wF5vRUDhD
JrbHYMLqIgas4tV/bbk9hvgxuBBGjkAc69zcU8p9COftCa+07JYGiXO4Jw55U3IoHLKdHgl1FY1b
VTyZ2Xe7ljeSBnLPIQFrGR4cJOJ1Le4sI6+BiIqTVd8X4ybgToyPL8W3HXg2ShXg5c6HqIWtAPJK
0DsjRZZ7mfzLYy+XPcDFvixk9Qcm7PlGUeyGCc6rNmmyTRB/Kb7fyXROTH4iaEG4cNO+Q4MRxKr2
YmwLt1xQ3jJTNYlhxyWySRSjRa8lx5bKC+Xkkfww3WWFhydlCenq2tPK2iYfAxohd9loQmWNR8FX
Lrp1n9k7Gspld6heWe9JSp3AjdRrxb50JoLZ18oT5tQTfGjIw2eYm/naflx6Q4oSORrUzLp9prGP
BV8xv4bJ8wtjCeN8tsCZQ4BGXckMnnqicYL6GGM3wfG71oEO/SDdZf1GDNTV10AuAac1cEzjOyzc
zbvjHpQbNwyzvy02uBIYifsqx2ITmdfVW3QmSrY45Kuegi95zQqXNpBF7PZcxoQz4D2N2FFszU82
l7o1uggnyyttW0Ik9rh2MKhOcMjXfHQu0qNHkc+YIKatsCPbhFGWJraYv850g7QsCI1x8Gha9NJd
/HpW7jbF3tVC2d9TfdV6X0kvCJQW3XzCFA+vxyP7FHDBZ60QbjssC1a5aTU86bT0YT3akA8PK8L1
gI8uQT8WlydaY2YB84ZvmMb8dyuFuqvo3+2x5EVOGWM2c2Df7G+5XWUCjz8wOke+Uo3tQ5qLJgUQ
kQKiT7rzI78Uf4gcNfJuH30JN9nhfmG8paFMnzODT2gMyrYlXlEO/06NDYTu1itShTAbiWlX4Swd
yQjRDLJQzoDmQwyGe7HKIlTz7MjgpnqOzEU5SttMp5qdt2Kcm4qwCy3Bs04I3laTANWwnk1CMBxj
vHJC5GWnvKvoi52YlhJlD7bWK/xARNp7d4vFYfvXDf9kq8lTdIIpU3Ok+bZugdbmK9OmU0pbHiY4
3YrL2qL0ESaoLGVMbgtSyxPu/MjpFp9YMsdaso82NSviZ2Px5i0RjlsaKOhf2+VE0XCqx4w89ytP
4vNpyxEZxrMrmN6j5eCJpQ4h3tJasaajz7kJJ319sRGqODHTce9LkWyiUhfTywyuXfKZFQ/NgEJZ
cU7YyNCWEkXy4KvcUY8sU1REMz01On4ots/jWsmzpPjdkkTKSK+7ilVxLC2qt/gHgOZy1Cjx3d7I
RK7V3b4tZQuvjvfzGI9xul6x3XTv2QYFfbDfTOpOLN27CZjfutQE0t1bXcgnp7kKMNARA40TSYZ0
QWcRlyRdJX8ovvG1l5MDllpzCE5JxorA9WSf4COSRTdie8g+peMCGr7W8bYVSLCKkzKT8Ftm/NdV
6ytPBNaxdA0teANXqWxn19c6Cuhx29/PyD5kWz6WrKfcfeBNB94VcDrUwCw3tYb4raSRC9WNraFS
fIce+O4P3cnfP7i/ezHkMn9RjovONRapvHQOGxWVuK0PIvXPAfRZ7c2wn4xJ0w57iRj8WckdBskL
3+FAKptfXMxjrT3IfDGjDREL7y038W0Izr7XviOcfNuc0teY26TWmtcfWuNAMhKX0dxCOOoAkD7l
AuGOgRzjWFd5DEW3lcz3U6If5D+OXsjW/ssdR38Jtb1NWroKqWW1dKsUEyp0ezj2f6F0+u2khsok
ZGNEPXZpzwjQ7uI2ROkOyw9KirybExIZEBaag+lFWDvf+75bkC5NtXobdLGuvGi7PwjVdTHzc9XZ
eC5P6epjkSmvfhPDdUQWprD0cpWf5rl76Q9HLs5+wxaAYDbdxwxXtOhPxsrymhQD+U4bHH/JUfDX
ETx60eaO+dCQtN0uRU6INj1jjXkkd+yMG0isOieNWtOmrPcxonv4XofKvqcvuqEAALbhQLcZxR6m
Qs8vY008VJX9UHVD6zjKiTwJgF4d9+9ALSusxfuS1M6nn64j3z0GtffDT8nWEgMjoQF+z7pgj8Dz
ePql6Z8wJjOtXlFBzkyHrDCEbTSMr8T86jlJW57/dGv2StFDN7QQ+NXddYuYBiEWO/lJIAoExon/
HcBQXjor7HF02yIE0Wio8mQ/BYAD9SUwgzIAJcTdEEDC9GN7Ddjmj4G1RRdWMqLV9p+q+H6H7KAO
FYRQHOLCKPNmIcBEuFvAw9q2PSMw/lTqEz49es9WW922u+ct/uJh7+ffrG2Kjk6ZIdd2QjzbDpy4
AQO6EfuuZhNDkSj2vsJeUvaBV6HqQweIFWyoDAKs+hezMvr3iTuAQlVx8crfN3bEcgFEOTmvBUsk
dtQ7BNRgbuff2WyYj++R6kPWM5f1eAiHxL8LlhEhJT1uA2zlayK/u96N02/ps3tNEaRHhMwvNjXG
4jVQanTA8n37xZCW17/XG6VU9bP+tmSg26+nWGsqLeebJRAS+XSW1tdcRupSdrYb7LODkbAg7eX2
QRjcl7evjZZ3nAlZj8pp0yxnI2XaxJN29R4759qjHKPjLPE7qft5ErLlO4h1tExD5gP1INMWtFsj
zosizMjBKNhoTTVza0IzuRXWrYf77qTQLuLEpLxbFO2JYSeRYxq41dy7wIYcH7iQy2pU/QG6rxZ1
YfKJ2q8nSnGTR/jMwgSAvRjfxIeCG/5qGZwWz3aAq1tjSMAkeNrwFjniexHs/SRsGwbC9QgAfSyq
gqILQnd3cBCdsCf1HCBmoOoO4Jz6dYGaXf5drrkPD40BdH6lv8UkUqldHBr8FXEU5cJ3+L2A5qfl
QSW+p8ALt9ssw3Xo/MkLIFfmvErRJJFc75eeOITp25le1AZzLAQNVF4HlS37LiWAsvkVDQdh5Rkf
Q7R/+lPqAwEtF9eaUmBKvsFZv8HnzK9iEcQ/IZohTHGEW0ZJfU0wtTG3OGS1HBS3eiSMrvXtlqUH
bH9aIDwo2spW9j3YcnsyGmCyrD0Kc1pQM/q+S2cQi1JNiTMGQD1XqDsNx7B1ipjBpeBrB8i0bzaJ
RTVJaaB06gHZw85Fd/AobUHQkumT0eCyANyquv+YdyNM8HIUSDsNUxqsmR9YL8oSY5E9KUcbTM6W
sKCjLGp+P2bN1pPhYqyxNFfi6AmjrOo1A6lm9wk2FISmMP39i71mp2XIJUggfXBqHOwQCJ62EgCk
LSyu0jB9Iy0xZ7K4CvhjagfOd0kWOzYpxhhrhbUjrUN5XKsG/6fg5mvcTRNT6QwMz5KODLgygE6d
5nrLTbtYTgIHyaP5pCbLIvrIBT6eUEbMsdEy8Ilivgiu8VMlgufo0Z/dmcMskm5vf2uXimA4EWII
IixwFa0skfl6mSUfCibLJSZO0LkLX2YA/m2GrEj+upn7jZ90CSnMirLLOn37bAsNZvEfiN/J5hes
nnxDhTuG5zChIqyGvXej6tcrw7bkbfUf8rhLQBWvjL02osoiCQOvkgeKAIsiNaS9Bfv+StmX4OOb
GK02k2NSYSDmn8QheImPPaU80EI7hrQxE/42lwa+qro4CEKZfsRFusZsmRIYtjR3vAvfWt6nQ5VC
33xZK2gstcJsB+MzIiLR8sbQiOVe0n2bspYxfL2pfdiGDvm2cICsZnat6EyX4TttIuHRcIsEt1kh
tBF5g3Vw5FGccfSKAtZ/xwdx1yFMDWa/LaOwcvOsxDs710etrdNLr1xd2brO+tVSs6WiLt4vobZp
WCFkb4UTuwH1RO4qsS/A+fqwiJdT7uXHZmHp/ZEs4iQWx0kUgyqbV2ygug15bv0uu0ln4t3W0rdi
tsCsRgvFD2sgWbj6i6XmRz6S48a/+EwVLVenaidxx+BOb2MVMSQkn3aZL2uesc3ndNBkgaCdo106
zL/BqnpMW9ux+LI09enHm0HRYqcWpzk5cz+7zRC6C2m8xf00bgtmXr/QurnvqmFGZcrmncxvhlXX
ER8O94MI+MFvYIUliA17VisjC+G92w1qXfZZpexLBfajw3qBrzTwi8tYkkMyPeUBTpYiXRJrOQKc
3mYioVnxK2Lvjv3B26OnqOONFPCYwsSCIgoQtvRtmkhAQT8xPLAxx+jsT7NqSBIFoX8JtIQEi/Kf
05ZSY+NvtU4UgnxY3CB7ngLxGi/OKiOmOd0yK9esC7CSACi4Cd39ZfnsmRKo/LoHn4MaeWm0zNzT
70O12MKECR36pyiFrvrwHMwDHfDfSA2OyaDzjjSPI6l5nF0irveUlc/7en3jNuaNv4pxJsqbAQ9g
UhETUMjAAfiTcSG5Hj3w+H3Vu6rkSTTFJr86huQG5t+76YJbpCFgVqcm65M0Xma+uwh+JfeXbV4e
a2GIbWEfXY+QQl1TkedU0QvM6pg7rDhjZ/PPjACY52BKgSGFWmefc5Midpzk7/jDsZEYLxM/ui/R
N2I8n02R8hmsXO4/NE6JmSuxfOalhlogEs7EOpx0U3m9EfebNceb3ljnooaqjnNXInR3LP7J/rd+
upfAhr2EZJolybqwAkv6rmLZUkKG9soZ1BOs8TkeLoyUVfeEyUatqM50II3zzs1RWGBuMSooGQfw
J0k31VllE07acdzgFb+AKvsPjwjsFf5LrUnA8Omdxn3RZSCHh/uOYcRQNBDHeNivihBohucZHbwI
rM027yKVr39ZBENshwB3gujcTp0jqAjYAIAazS6RO/FNeVFqAG8KROn8CXR2RZ8OJQe+0tTC9u/N
xdhlnNRNayuncZ4f/P9eTA4Y2YNFn/carf8jMoDqA9pOdNOQfPCy1ce5Ty7v6N0n9STxkeOT2Kx7
I4RIyDTkr1Lr+qgrol4oh/LIKjeIUGp+/TCR6CXpr40XRqRq8IvWhNeaucGyg/3UdA75qUhLPCVp
YaeUcyvnXzYd8vH7/lnL102i8o+pDBml8pPJyTn9uKN6A40mkjUivqWnfbYsZaZaHUUdQtYZ4It3
q5QPZtPQFmUWVhjgMOxsZwqz9ao1qaf1x6hvlSlBsstV2PeHseetnBmWLbrefO2JL8nK74YwkxE6
z9JVv4XOYs4Sk2U8caDlsr2Hhc7Ypr8Zo/4Jo1wXAvLeqQajEc4Gf2Ay2Z+Klt4mDCyBPT3ezSzM
t9gG8m/NPYwuwL4eXo7BwYY5yXTbXNlHl9W9BkzDhCrpHGDG4QbA6mmuN426P5nMzewEAv7G8tHo
5zVhnjkMKeIUM1rEcfABfuPGV9WoQfuamFq6TzNzTl9tTnO6ogmVZuneMM0VAEhMu3zcWEC0ZR64
DvblQskj3RjPTeI36EDS/hDiReFbw3p/XI/L8asi6qd5RGzweX/ZL7/qUxpZ+Oy+cvR6OEQ7NPIA
SzXXAN+tiPXWfqfQkreU39xZPJcQZR+vNtzCd3TLTnXkZALFQLeeFn+1PopZe/Kff/s1J7O/W+ox
Igfdv4Dmb2QmRSyAZWMgjSxTm8JMfe57Dlv/Lv3dc16V4aFOVVh7uzPGJ/Y70Dk0D0OKtGUHMbUE
/cmY3MAS7B8hAO0ZsUF8zrgUNHAvtraHBk0MdDr4fLkkrHyyGEag3Xqp7drJ7bp63XzIRIHfTUgX
m1afZb3mDNQJW/JnRF3T5jy3VW0s3GqGcDlWbL/UJBsCEvkNYoB5nlpGowU8FG18L50EnSmvCBWM
WJQxhEJtMoVB5KNzQAGbtW2NE8DvVKbh937aYnfVBQ9Gd8Kr6KQbMoVFrWN64CNCzrVNqggFaF0p
VAdwsELMaqUsSiabWHmENd6NHnpg0ihtwqDA7gG7joa/li3xc9Feujwu7Ch2rq0goYwMDODnDxNx
dE4wbxnJe75gPC3BrYeB5cYVYlAaW+lcPKs8EiWwLVddqHZJ0pKt9XDdAMe10QHJHDKPUMTjipNv
t1cfwtfB2KwSpZFA9jta2Sko+Fw9Rq0HAodQLkwy+8jUMSK4ovrQ3M9TNtACa6Rq64GtmYei6G2e
cK0ZzBQFG/SD38XZBqAuoLRQI1ETCXtKzahI05RVGHQ2/f9ypoNUJyV6rauUx7LKd5jLzRvkeaSh
6dP8T74ecCiibo6o0VGmk6HC/2usXhGKwT1/5Rh70cZM9D8mJ1or5xKIVa1mS/AHpMdVoiju+IIC
vdZF1/YsVKUVSd9BSXTkB8fB8Y7+feuqB+IyD4pUj7DCm+aw4IVEDlyPCpvmaTYuZdp6fKR66rK9
GtIzusjcGl6mWDW4v/aIw6gBIusml44AYq6fKSk7RC1quyZ0ibPAJm8dH4hO1JKkyQevJlK7E1aZ
TtBGRIrMlrFuTWn4oBJ/bX6oLggHozrauDANTiVros5WjpdL9X+RXMt7qkTGXjD4Q8hZJNcD/xrD
RKlm88ryUzDDwBZMFXzbHxkJsXPuDY/v2S3nsd8wuZPCHF5vnQ7PqBOVIqbGXFml5jLuCQKXwTqz
t8NfFQM22r6LkcPg9TcupMQlmerV6y4GaTlzeBboLIyXYFANzAFN8oa8IYrbi4fPiOg22TfFAZ+Y
zkgIKNZVl32nlXGWAleESLgtyJ+kLevzeN0ImqCea1JGjdrK2gkViFTB8ekPsOsFyUS7kkQAft5a
rq2dkPEn33ovfUF2rUzFSfPY6QaSPum6iJc79cXJlZ3xlDiqT76sy4BSgKA3ya7eS4m9Iy/JyVSj
3W5ZIDUXmtWoennikkSO8pvRimc01qaI2zMt/LXpRiIIa5ByAb+P9WqGjTnRu/xCO3jt7eGJIZg0
64UpogxCwsj0joUhtr4SAlZG5+zsoDg/Klnu7KXBsNZ+JtPXa6EwFPWfx2JThmpiV8aMjRY/+tJc
st8iRkxt/TQuNDH1fddpFkP3gYtI8F+Cawe8tCzyNlx+W6iWmcbTH7IQzjvj5m3qlvn4E6a4F3iG
2nWbmN0XDjPM+Pcj/YasUtH4qvSqZdDA0/MOmUTxKGMHrHKBhyqdjyrnBI6iV4+VBDs3e4onD2X5
PhWz+Y/bHDIsDzaRsl6xQWY65iJwdvXDx1JWV73WZcdunvot8uiQejN/rErd9T0DmYIae8JiPf2L
+1euEoNuKE4iboEtDobI/CxiV+Bz4fZNdgZtpVZiM9RPiuoSijTwHIir7rwQabd/A4ZMcaNWoZfn
fEXi9Dhoxh0v3ykiqClzXRdQKHaMIVfkPvIq9yukriYlKk3GSZvb2njcRG0mMU6Mb08uX8AxYObc
0NnIQ3v9uQw7Al0dXs6gOwdhZ5Gg1mXEHdn+hugj4U2lwqH4cH3VahgdMnqx/RN1QUcqGM6ML+Nr
ArfZ1qDqPXpefLbneAtffESMpfbkZHcIp/Vu/l45wuchN8ldvDJjMDtTxgkCj7AB70fUUBXYoblX
RV1A1bLPmjksX5Z67gyPfJRHIx5gq/u7axOe/uKy9T7mxxe4ZASnS6/jBNT/UCAVE3gfeVWarqzy
PAAkaUoNhr4auD5oSB9Ye0cmwvK+dl30XpHgvh0SIA5sZX7igfDkNGgoIOFcz2vFDkn+qC8EVR3f
Z9v8l+eZ9RSxDnpzm/UeOtfYy9chT0QiGGELcX6z9ZKbtRSd2MImLIIgCwboEEhN5ejIPMjKYoMt
rt72C5osTdTQ5uzqiyhAA1Zc7IFI2ewS9+1R0l9grV8mXbs5O7KhxSPLIVhqFtVdkhE1UPHtqvKz
OQpVtYo4+IXzN2MMoWyn1MWff3MKIoUSwgqz7p6O38CvXG3w0KU0Y8fHzpHfl2ofA+0qofX2rsTl
Mz45LxDuJwW3Wqao4mbJdcyQyqxThl92AQp9acTtubCwxWL24k7cNuaUibQvWCBALUVt7+KcmEbI
wpg1FU/TDa+gedeGQAbb4BV68ZN8oipxZJTkKx4xN3vpGXEvMZMQBKmxz95Zny88uwJikNKkbGxC
iNBhIh9u3x/rxLlIFf+DiNy6oAO9RE/JiRqqH7p+9fMRDUdjISW85ATmFRi5hdRG84yOBFNl9PyZ
IPPd3sEuGs/NhTHKdfLS3QMH18B1GjWrGYtPDjjWhjUA+QykjS/mepxGrIYmfyJjH+R/80FV7hmd
NOIabcruZwg+u0Z6eqoMYigmC6bob3A00VZgF1ed97VMj37/zQuy8ZKczV4iWs5SxN7pbKFhUUZE
L6AwhLp4q32A/9xliN7XFyGXDxHZ4hfBhNyJYsoiRC7S0rnmK0VPKWcwhtYT/qEbDJdE0jod7GVd
lZ7R6dGzwP3wcWyZy26N3ruV2x1tbobws4zGUj0TKUqHzkRmDfIxPCYUb0EteQO6ozCETzLuwjY9
Hrcm0pmbxeDlLTh7CA9WJNkJuO+KtYi3UoOQiZYrGoi+I9uSpaKIA0rlZA4W5q8Xe2j1Mcp5OUcf
202KbFx0bQ13e4ZbxQ3SHffWjFmB7ctVbvCUV+a2kJNUArywgoFDyEhV4I2rwaj8z2IRlXgJQzyr
WfnenGcvmqobVf6a0Rz+g+wpEuFgyrcot5oxNo7hJZanRoA/QSjS/1qxNMDwBJbh1mtXWZEahOav
IWLN9ueUpYRZ+E6qr2w5ZewKj9UoO9sjtl+2iBqoEQZDHpBHbPjWAJ3uPCFMNrBwJ+TBuK3HfgZU
/mHXAzRGeVsPCOhCfzSG5uMjuTNjqLA0ndqJI3S974ALXXrjoT1ZpYGSCjDrDJCvXGfSnnTgFmXl
/mkYd7o1/wbfYGgdhGxKgaqDhULF2Iy+zCLmxy7w2WNKCYE9HJFX8FyG8j+HPRv8fq0rfxuCZJGW
xHYUJ+QJZrObRsy/4raUeFm+HszrXrIeiFIUR/7BNCgFVm1fk9de42QKeI5N/lTYl0v9viWbBIjy
S0B2gGXI6TXWI8kALbFgOLE0CKGkzJHjfd3LtKJRvpNbK+c9JyELRJxONvwH1KPyOO04xe/yIflA
qo/vQ5IW6jfbBnTOxhJbSz5ZgL2/OOj/D0dXwvlrtto3ahKbL0w0U0+Ulv0nDdHEg2npCWD0vuVe
OY/GsiFZ2b1sPROsODuTlDBsk8TSvEx1l2eI3PUVJo9LXmosUUoUMnO6R12jqKaNsb/9cpbThj3n
3OUmN90fdZh5nJAUQ6I+I3vv6Xn5OjA9l6uHLaru1TpdPPrH1Ln5U20lNrsFpa1NOOAoLqQmojI3
2mgry/WmUSAH8Ty9l/IXH6R8oEwioE4DmktGeU4cOnNpxlQw3PLzz2mGI/k2WFlASGp1M0Bt2gvj
PbVFpNXbjO4zsjR2xmSntEjMkcUN2LtG++uFj9FEXGqDCkREw8RwrFGCsF254zk9atIUBzgT8RKK
QNPDWoByta1A793loXmbTTP57LbZtkE4cH83TDi3WX3GQV+RXTmn2IPBdAKSRCPzpB74XoNz8Qg3
X1sUVLVCiDVkUlv3o/FYZtPfqGoLk96dudkjD1IhREG2MLmA5j843h1hoMyi2ayb5jn1zvRrT+5n
rA0NOtIfIL7TXbOFa2+EX2NdJDzDwbKmzOcvrBCCNzFEaX9GmBluLhLkf1D1+EPcjSBDrxvLlDWL
Oxse4/bjdllYjc8Zl8m2uasrmACYEWLW1JKJcyafcdEZrAtsEIy7KJhQUOt4GTvl+gN77t7tiewd
v2T10IYGrTCEkT5Y+l7YZEVgvIrcJAmBmzxpBYofw+fgvizfq5arRzsgUEIM0aiHoYwsc80v0/Gv
OLzRM5hRAbThnHU/MN196HK0W4GtZ5aMKZN15+m3p0HBH4S4dtlYdmmTI+iZYIw5EFrBjldWaimO
37yMJuWULzm5TjWr6a2k1uLrTRoisF25ZRV+NyHAXzhUucnXhe/I5Z/ccAwCG1t/GiUY8UFViIAB
XkmuTzddr0sf4JxZKUT4XWP6U+wQMRHhPEDQ6u6yYrRmq4li9wSff7z3+I98DeeYX/uK87NBKIuw
6cKBGl3Lmr/vDYVMzGHr63ugMmT1f9ytzTezWP1UcudGm22AlE2BN6gM5nAnCN/+96nFb+OAx9DP
ALdYou+J48eyDjrgwWgZeE7kGnZOnM/CE9f1V6PEaYNQIqMgiBqQHhV/uAoSVDPsLUf1YmG/zB7K
vjJSFiXjjXcmrh4G/mw6Y8f8YKIzt2JB/OJI5NHkAl2AzHpANlfvjYU3uXhE0jtOR0FQDUHcLt8N
fE0iOo8hfp7zDbuYVD21FOip+FxD7gYpVa5P675+cBvswTY45EWIQGjHG8wo8hCqaLjifK6up6C1
UaThqcmyvGGuWiXZoGLtuQj/eQSCGniUFiyJGptvbrGZXPLWxJdyoWwEnjGuad5HMefPchYNPJ8c
vKeOFkdmw96Xg6BX/1SF1SmiwCbvT8T5ZDPM+BNeTWYrAOj8dpRUhEFH8b4RmIxUE+KmgS4Q4/7i
xbcKmJPsxXa4P7h0Dhu6QuTQOFlViPHnJdEsxUJ9Gl8b557bO+tr0rFYywYXO1JalUFCsdmAkmwq
bZ3FuspXKO4psYrvBAmRta1U5FfHJAv3IKveXtq5MLwADb225i09NSgLEaHLe9PYolPvnMlxpPwr
5V7rS+9NiKFqmFQ0GqrwCuawyepsDNK9Caq/b5DoinBeR3g+lWY+AmsqzikVKK0uWcUuSCXVCHW5
1acUkcd3RCGjjpeyJGhhdsJwB4vACv8xxnyUXOvQEOZieWQ13wBfxWM8MtvTjxBFxUsq7OFP2lu4
00VCfVP49pU3xZObLbkL8E1t+NkCnnRD7ZQHiW4+gBXQRomTy3v186UW+J88oSH/F2luyQJ+SOMR
+QSzRbH0NuGrYaBai5INbb+YU5HIjhv1AnlGNFAvfLh7TCB0TORCqdCvMWtTJ70q83dpIZamZCZn
kmsh507v9ok4GIGvql6qygF/RO3sU0CzbrzbtEbOE5JN6huOQnIyq4OwTt2RPIn4uzPZbTg43ipb
kzPoPklKq7NcXb2NNpOmE+5yA7UuHFlnATlQMqp/VrVcYD55xxcb1IT2zTXO4WM02i2As+7MKehP
fhzqiIf7KvtpQsQh7ZTJxyncBP/sOFskffIbzbreJDeH09LYni+LSnC/xCmKFhwJeYW+ZSlj/Cc6
X4NMTMR1BVJFXbh2RWvmJk1eyN8wMZD1exBZUhnGofoEwLZE3g+XhHOor3TKrFOI68iZZl5u+5xJ
rQQhHT9lanOIzxWpDtYV78zaYDO8KzoIMuGdLT30QHBS8COjYDibk/M8eMq89Ldtjouxv/yBE/kV
0XnzUsAK4V8mcbXAqbvX+tkVUreRsEMjp+0RaXIZ7UtIDzDmM6iEkFjwGR8CCERZzKVSwv4iDDsz
8X2VdE4/jXxZIi29rM2IGmUnM7afMkEe20ipYLzeg/cpMTlp6didSmd7OzuIdwDXULAOdrEDBYog
xFUX+METFHOqBA2++99vLrhkHQE5fqe8ZM9Wr+Pf8SqUFK4OUw1k7dJBuf/qyjamQJaNtuSSZi8R
O5qZjZkcVtmBRNqT0boniIlBPZ0rEd6yhnE+xUZhwueJYv+FZYvS54ha+28OvcOkdAjomY0DibdR
vDJDbXuS9zGva+JDEG6kdvBur99GOgs8RdNBdn815h5GrwRLnRuZ+OmAMtd3aUuy1vWFxWzQRPZg
9eQhEDmp7Lh41emyyFZahMOhBZ/aKiY4QXYFTcce6LIFh8AU61yNzlm+OTsF9kukeCI5xhMdGtcc
IOqX4Wh1EViANtx2VlE+6lPwxLxkQqPOaN1J5/uYYQdVN1VfnFRMG955qioByKJiKZ+ghj68DL1z
z03LVo9H35DGEPJBfW+hwfyFTVbuDdKzuERXEiNTPDpvm1JyZ/D9VU/nKv8Ca666bB4LeYgnlrmD
dqWwNR9Onl7Rhxftl3T46qEWUbs5sKyruaJkt85sV8mbNcgP6CYc/uo33uchm2FFeXCGAJ5eTG+t
A76gyudfk8PDc/CA0zwrh5/zd/+6N41C/nDa/kcP/yhVQtQlSdy75RMKkvE6S0uJIwL7nkg5Ic5N
Fi2azqPh1JBhdoysIgWk6A1I4r7CCvWgxk+P8xBNFh7vA8CvR+d5V2VNjM9QP9TWm8lh8k1X5a/x
OM8wdFkiu6xcadGrAqiGnyO5k/kLqcu+aO3LDg3EGz2GwFcaEUaucnOq60xAV8WoWVk3fX4ms5rP
r+5yiip1SjSLiVOPLM8+UR8bV5N22dk84Xvj8GtaafVZyj2E3MjccypV+gKMdM1uYwoDaFO5dVaf
WkeCTMLiSCn6R4PWlXBTcNnEQF1Ztji7rQmnZwBjfIsHujETgfiZphAfCtW3ScVqK3VwYqsJEBN1
WxN8PhZHmwiZqzDX/52SldDuz5CtB2oEombooYeRWZkL5TkkJd2tDBo7M1+XmGk3O/V8VQfwfykw
xE/pOfzSmbDKGntZFgiohOxd2KoEfSV5xV4duyKiqDX7Xp0oydOhFiSsikcXbs8qz0eXm/nANrTX
cBcXFSrTex7sPq/NW4hdrqK5P+XneoQSbOwWiEEcirLVb7m1betXzbs9vQ9IKwEwNfotnXQfwCVH
g3xGjTnHtaEQx6+U9cS4sw0fssVi4jaOoSxlqOBYEd74xcfuhzv1hZYBRCi95Z99uh6HoATsTWlz
k+EQ+hMajnyyfTalrmRBWq+IuZpPELVT7RpFrOsy26WdOvC2VqmewIjzCB7ZQR11OPEuotdoGNzN
IJh6CfMGlOfHDrtdt7i5bJk+M2f0bEpObzwN00+Sh6F4OfMHRaM5dPiY9KjlZVdg5NVfkKtDP6Zl
WUMnPCn2d/PHbJFTi4ZN6IbFAV/KB/MT38DtIkxZvSLYVrODKlAt7cyHqv+ViPrVvMpTxOsxe0V/
5DOMSPEP0FTQ5zNXFyfqslUhm83kHFUgldxFFsiE+2oQFVjvnrUXGZ4hnQyiQX/duZ5uaIPoXo40
nElDcLT1WRHm19qbTumD+IyMLzQM5c7/lUzqBUKsFMMC+19RT/Ve+3sli/Pk9XAafhB0GhvoiDcG
4vFXgaPD/G9BskqacVMADAXflzLqTVVlBWjdCtQd5HGdc4xc7ydHP/3tcGRMalZU+I/adjU06keK
3HlDfXSoc+HXADYIwDYK/JvPuDzql32r0oyEQ0YpY4+4Q54cDFUW0Bi7rduINx/g0vLReWvztcTF
OO39AJHmEGcdwWGJrpbDS8ZvK+LF+nV2PBc+nKFq6DuW1Jm6tzgRW8xCFdxpM1bB6PNlSTRneSmS
WBRM5nsraA21N3jLdXOInwolUarDtML/mqnkZqG9rC/46hduo9yGRUkgNYacp3gDbRc+0SoH/Amx
oU/4TWd1Yp31v52XYuNMIBo/MDxLn2SOG22/Ry94bE29JoYDpEOp/IrmbpO+XZuGMhL1C5j8Zn+x
Fy7ijFtQN4amcNdDYdDS+JgEEiMq4JWwyqP04I/DlWVNk2WFCr/bzxALp4z6N2YhvDLaICKxMfS6
6ifhG0eNFnwkKqBIUIv7hhJsSYK81WK3x1ayKROU6u5AZGsdfdMko/VTFS6C1D7zbRZSVMUdKOnI
fQmtreumag1QCXUQ7PT/q5Hr99L5c3JfztD2Fy88FIxxBv2Zz8W8/zUuSd7NdHcx5InPgxz6KzZq
7nwVbX7heoBsxJzU7WJId2WmJT9bk0j1D+C2OvYYXxr40sZizLp3lDVCXYjPcJ0O+U0zCeFHMx+f
lstFPBgykXwhhv7UQ5hPeYY5gWwcjDZsD8oQXIORKn67oTSLvWr6O4IpgjdIxJXqW3RpvJbNHqRt
pPeVGNoyc5XjGSPbkMeDmg0vHVZDB+kn0RZc2aLo+I2FDkZDJOiF82aAilpy6ME6Z0rFK46efC4N
ApMGkZfk3FwjtYLmSV96ut+ATs45rAXJeCjVsdimcYFs/WBFgrEPUdr8iflgV8UqD07FXw5v/zKf
HImwpQIQL9muMpjxB0l7eAK+yYEkzMX36iGb9f9XIDlaOFnjX2gfq9k3svnkbW/bEbZ9LWZbk5Tn
kz0qIOZv0jEw4efLibQIK8wa7POA4D/P1PHutJLghSB6waoa4qct7Ww+clgJrtMJIVZIazTA1SzR
sVnUDqZDIfgzr0CdXaB0Jc0Jy1n9T5uknxEVEzn0nF7dId//JTHa9WtELQKnr+osKWGAbmHI3wu0
rqIH6OM+Wz+9XCaQ9M35lUWsXPywE3kwKJj2C3ErsXPpp2fglKQBXI9l64ebR+REm4ajDZSCzhBl
2YDAq+jPHnnhrnvURwzVG5Xwel9ZcRDiKsMjwHbh/K2t3Y36pNQW3Vj+c1AG7xSC8kLLo9y7lB8O
F6/mA+dCdz48Rg8lvA7EU+rphnIB4Ptw+Ns3BBTDU9BbvcExz9Rs+Dfnz3NXwocSmXQW5f3LRx2B
Rf/Mdl6uiBlv7ZkveJhH81uEJ3e/8owyDDjY3IMgFhfO91EmB02ozaKaFTTPvUinqdpJOvZvjxdA
X3c49hls8xJMtsPYHCWd8g+jl71ieIKG9Fk1rvxpmhEbEWL+oUXTD4Dze9y98mJ1TRv7APOi5+Qy
R8LCDAzwt4oksL0Mv3NFKVfoR1CBsLfzk6SQSNalyd/beKMpIXcyFi+2WVmyNHJlUnDR9xCeUmui
FPU1C7gK0/9rKYiXyIS4JkQivRE8k0h/9vlffcj1yISq4I7QZ3FYfnvPjbs9NGuCr2kx33YYlPKh
mLwgZBOwiEx+vUIDuzElHgA1qM7vXeSc2tukYIBkqyx2aHBsDqDRE8+d82mAGVAeQ61vvFfJdCBH
lt1QDj/vSmxB94mkwQ+TPXPCw0MP2O+NxQ1NuHzQVybkTSweypfWzeJGJ5EovfiYYkorjcHWDl+a
+s5gMnOQWvIQL87Edk9MfVOulZM437n5Gijn1ErjzT1XNTQGO0CQwBM/DPhnH5X2XUi0lDKXTMue
ixMg3AAZmxzQGDMax065w6a7QPGCnNHMNlbF9le8dqyJWRUqfBZZD9LCb/Vr9xvbHexsFhb6cQ+R
UFR2sIrCCjOaPrm8bQG4JJXFlg1tSdJYH5Kj/Mx8kB8g5dlO+6/jF48+NrPZFwK7Ycd0WAPiglvO
rHQ4goSgwEkJk8gvQzC9NBIMWI7CNmJT8IljCAR9vLENTG18K5viBk4VnbRp+tTBT70DXoF21mCO
S6FfS9v98RZgcFzHSYO9T8pcw7TWPngfiTHjA9C1i6C17WYCUAWRWH8Qkob6qBoglfRsRpBVH6Cr
xv7Tbf1WyfFIwOAw1xXJPamGPllTGmUzBU9wYNztGVE5XcWW2hAI0UzdjzKhePPpRkznJZIfU6Mi
oW1rTKjoQ3xxh3oSDO6k0xjUOfHTFh9prYrVeETXAXEYU8XgSRYdq5D6xSXzIP8fqCnnKptbOECQ
75IOhHmrkdTcVfGZv96UnWxMEB/7JP++fvY77PVlbj4Cz50aTlG5seM2bcnoUIj1TrAObpEMpiOe
XZwp++6OWv+kYyCD+lEAo1mkpudk+NpjPvwigUEKZSf8i0c97US5B6n0pQflTUWxO+dZV8nFaezM
vFzzddMX5GKthH+9NUQ5QCRgpSBCn1RxEmq+/3MrHjN7PeK0Ft9xRR8wAavi+WRiPQItE9JA6VNf
GLFnoOWgccrCln9AC5i6XDdbSH6V1yD/At4UHvonhDZB0oxFZYFv1DZu0r82wSTOP4G85kO1v+7M
A6LJ39bH9U5Jnnwwe0oq7NLhET1JFsYvqGGRh2EiQ0akvxcs+Oh25192JoJXIEGNbKC/k+DfdG52
AV3dklE+ER7o49jL8+4dP6N0qKDMhYfEhBVmdsu9hyk/F3GRc2J3fICyZjssXDEOvz7MdT7qE5f2
w8xppkfps1bGfhJDjyZRrfJE8RS60SkQMUzKf79a275Y8xA25g7cVwI1GqLHeJdQ5p7GnIdkhF3n
zWc0uJazuzsVl7VBtix8uJMJFm2aZHXGwQraHgQSdb0u0+deDnJv23Qu6J/MuxMcD5pEX5ZX/zaY
1/2IwZwOqqr72BYtHrEI8M/5Lgy0XUEpJeRGCD/LUh5liT78tHacLew0CAdeOOon4VZdVsmKSiSV
vKJGNWTRkZ17NxTcn6ndPtYGYQafG0KvSj9pzeNWUGGawJbalB2Nx460K+UUvANnRJ5IJM0WTKlA
cRfvga2K7+tnhw8i+V0BJYcZl5VW2Skse60+XkOxQoaER6oPHK7ukD90vXuSXAU1ndcnSRcGg87V
7kmD+IikoJXMt2m5pXvRX1ccR5+WmiWhVJ0BYzUbDLdWITM4G3ysJ5ANs9TgvHMYCrCZe0xeqgt3
LFaous7l73WktyTjxbT32Rr7C1P+7w2nHz4bdEnFldysgbuZPNPww7SKb5G062kHy3f0zyT/uCCI
kSjc4fvjHXUYVhAI2wu8LktVcJwN7nnp32eBHhnGnoSJQDWXCmUMbznCoT03FtAstpM/GmiXiYBp
lUGmC88HE4WjqEPjg7b4E9LAYZ8NqyNv/gsPq+j+CHyZd1KciAfP6mGbHC+I0EycLvgZG+oyajMQ
Qk+fEMr/yDTgM5EBuYTMTBhfB616dS626j7dOiPel+g3jNEgX8vXR8I1hsoYkE4Z3gTTKdJJdkoj
BvZnFgWuyIHcsNq9fytJCTY0LdN3hlZflE0F4CFliPwBgzrjPkVGkKsxno1sq9WKZfxtO0t6d+UG
CChjtDNu/2DFR9z0Utpyu3HjTm/dybyBmBh3zd1MG7CRCP0QXhGsv9xQsV4WjIb1DgAQyj26u/wo
y+TJpYH1olA2wXn50l7Nrfeo3gmXHhV3K3pVXpsO3iTILm+lmhR0d5u61STc4+16O678DXByvY6S
AhY6e+TMnbgY958EVRVsf62x3IW9wtrX5MbODqeaBqyY1/xtE2EYOlhYJb2Lkf8mBBVuglWpEvFX
nesibUKNWFy7NZbx9rU1iM2MeN1jmoKPORopJRSXrlxGuaoPk9dp1knMnVf4AKzhtV0DyIc/qQ46
aZLA79zp0XkIDZAcG6yK4DLG/ajzGROiOipI8CoWDhjY4v3MOcg8WxOKIH3vRzG2DSjKAGAJHkkv
2M4ph0u32KsdMAZanwcfA97vxwDF3DdMbeT2J+iVPmgq6WroPk+mPVAij7P8eQbtkuNJaeXNSErQ
9s1apCOJkTrDhQ1/vxgEReVtSeVxXzEyuiDFGI1k3YGcNxRnqdBrr/WEHcIltxfytMPH5GzHld6c
FBP03culP+SJEZBtXAibsabncoNqQ9Rtjn12Ar8oQ60RsaWvkZIfSFCXbsnBxyOv7vqlfzUOMT2x
n12Le0RUB4P4EMxs6nsgAOXRqv3hdIg2maOB6ceekOycerFjVIdgtrrl6AxfZF99vB1DDFn2v/CZ
gUmxYXvUsl+gNbEsMfXfkok+8xttyCSrsEpfJ1RgvNzNZ67juBF6X1vkiiSYDh0Eur8rXOqEHwuS
KYFl+aqSpXTUyJ7SzoSnnPjLl3bV8cKSgO3PEAbVFCb2i1SZZ7dNNMGp/7qYH1oph9ZCkIFLSGIj
4hnNqZaG0eccMLhBB8g3voCbCoVHleyo61X40kg94ZhsLeenGogXwhAhbk59RCurcPYrc85zyxgZ
F9AOI7IbJ1GldhzyhMYm9ozTDtZyV8cKn22MEeS1EQNYMgIvyOg21d+1+bjRkG3IKbjZjxqQKiZ0
MTNiUIkPvl5asgGJCQh1w+j2MXipDm3t+Gbp1Z4mSFSiHKG3GlPeEwuV72D/3JtEgfl8nCQdY/MX
Fg9yeOFO4nyyPxhgCJiANcausJxgztYCwCHgM7N+ImkI0URlyUrhgksiMBoLfv1h+U1Xcj3XC0TG
U+oI5jgY4zDx2BZjiHaXP8VjZUEp7nC2gzDijv5pXHzDeoKAd7FBql3lXHhIzj6ItJhgSl4DN5UV
xwJAIx5sKFpfmGl6pQrJQQB7Yo5ZeR30HNG5KvyTbhZJyIw4OV7Dw17NUqYNCq+Cqo7JWB4zr5pE
EGO/+wqy5yGU7UNQoSXiXtJUlHubskp9itscv2IAG7Fr6+YYgqONwXJFuXjrEHdysj+QppsHPZkQ
+QGJKKvDQxwHNIHGjr3bcmoGqJnWlOGT6PN/EuI9Q4KB7rntJkUGSKcwrN8SJd77hw9K/iUQxAvD
oIYK308EYEASxk2J/mhqgIFBoIF/PQPKBOQnGEPSOoNqEA1Qm/17eqKBVZwEJIAzibSb4cXUV/dl
CSi4coz94gRBr1AqANTfwCfsu9EiPVM/yff1shnW6e3/yC5zWbNiEnFPQhG1ZXypsmJwSpJy+BlS
WxAbxKpeHXVYpxSHhICIT+t7h5xSLuzLwy3vsp/w/zLKy2H0s0LODRcywRpDaDvhS1NhU/DCpckr
WJFuwx+RB9OvvGmU8fchBkR92d0TT2HvX3YtuhVMzQFN/L9Vqh9n2BrBTT2e3y0skIFX5RPWjjQ3
dy9Sq43B1TkosDE8xR06yZlaVktkQIJcEL31RRUJIV6OMARF2tAjX1wIODhW8+6qVW2s+mitS0jI
kLo437AlsXOFdmciPO9Q+Rh06Z4CqcL/ZBCe4RFEasjmsuLeqfrHzUa5oi1lGurW38uj0vHBZymz
YfgAQw+p7RclleEUVRsQ5rwRfBbMXRO6kErGadxv7GbMghNfM1ArVxyuc8zTDQrp5mzSjUne1lTE
pbX51leEELufM82AAT9k2ZlZra1u061xjDM4temkc6QvFdRlFHgOz5rJTXjLF/QXaQgy4TnY5LK4
8wW5/El1p+Wfm7wIfEXnDk6BkVumJ/yiE1qZXSh6o/zeWMvB7X8vp3COxP/Z3x1uiOo7g5AZOqjp
uCc79iUvIKSrMwwkYW7QRGIZ0E5ZuLr103O9x+lcK3r1dJlyC5jRvTg3B6s+cTXLhZtL3s9fbPBM
iLwMFPFWSfu+RMjvlsPu5Wd4XS2lnWggdf5zAEMEDBDSgrwvbI2I6MXbV8qps+S+PURhVmFJsvZq
vgyUhosDyDyf8XfgR3HMSyH3BnH/z9HMCjBFDtEo/h4aiUayZOGynFlghg0li196woRIF0t7sGqw
odponBwpy2q1jJnqFKH9y4VzyqJkvov53/Xyd7pBkr5Dnr5FMMBduYt9tLbbbE2fDdbKH3fEXYQO
I4eQo2sDD02L/PUI+xOoaMqbBLtckkVGUGTyK6l01GXRMgDLuYFF4FtbpKAjazt+8qBgWPXxq+aI
HLdqKoXQ0xE27x3rno404SBqnaKF0etFYVpsolNuXxmLTHClivxS2+plyRjyANgTgYbAbyoDrzFT
V4NCrxpB0BUxKPKWhNkaF+vWeMXYZi24TooVN5DzYKjGxP8NI3MTS5R7S9zVudReq3d+nT69XC7M
6JbQlbvYlQZy6IEm2OwqOed9nChYQiarW9CvX3vX/dvbKosL5bHNC7V70LZrbdIvz3QXkLS909Cl
PlL9G3ZHZ9BETvjoEbiUzqkdzt8b7cNDtheRF9XOvQVgnU90la2r6q52QGwvBVYJ8jVCm7KlrfOF
5vDSsFEOyKE7XUV0Lz1HedTA0aQjNh9A4th2JrjRxYSPpGh92R/HAqFsedrY8WHWbuAgyzU+arSE
Ud9veff5b3CjX9FRMCAfa6aQQmaQ6ALKyMuY/BJH8dtGRngCK4Heft9gvD9T0m/PD7t0UbZ2tz7k
bz/P1vdyqPV7GSrnyxvYAFFM5ONtECbwHHugpLu8YZy+MIRLtMB17l8orT44BlcnP6yONLWVqGR8
I6nJrq4s1Ga/TVXtA0Bta5KDY/ZWtYoST9mbDuIss5xiUQAqfcmWF5FmHvih9ZdwpHxtyfYSQwmt
aCc0BQnrho25HuxqnogLQyb1pl3YniTZryqW3l/6c1Nu5gtHDx8K4GbIDbxO0zTKIs1TcwKVeTdu
oPQQfbm0g8vex2WOTmPdhOZkc/1vUCIGJ7ioPMvOndECcJE3Rqam/zv8RkSY58QTjgq4546p4rjp
lAxgD/i2t8kN+NbtNMKPo54YA/owA+iB7/F/Rc5wqSJB6882MkkTM+koLWmcokiTsFEosiKe96Lc
I2TMKcx1LMTZGqA+vmPIG7EIstKhLZnD/zh+im3UEQRRjjEN2qdVdInHvLIYUzEIHvx/mPMlKDcU
9DIapzrmobWruyLjIIqUaVq6jsyr90o2rz0t1O9yKIk+cMlVz47hzcON9Kar3mB8UDNhmEOCdIYp
waiUPmN+6Sq8jSOqE2AsQnfFvwYx4eecNrZWy5PhCVahT6PR+ZEv1BF2qzCGHI+PDkr9oGkrwpvG
65X0PmFoJoC2lFeuKnVg17ELA5gEvu9HhGg71g7kUqYEaPycCwZwRGGCP4udPG878FqcbBfoNean
vfHsZrTz0VVUJvmT5Znyly22LOiefVuFXjGJrh2SJLKutJFN41bMNkPywF/vWYgCq611GeFCcBaQ
7aVaI1SWdBBoIHR+i/oYCcBByul6zQp52ALxAXa/7KPs9HDA8N77ImmQ0F4n33AZK1PiiNcyhq1S
idjZDgXChjfIEG2Xo3WkO/3e6hi8DMb7+nRkpgQb+CnRARa/7KNbyelgV4udENGy98ckqXel6DpI
ix9VIjP+iBDyt93Bg2ISN/gnIsa33dj5iJpGqvWDH3+G2Px98V41TBK5ou1Z9TYb2S/L0y65PPHU
2TByjC9boLJr0c+KdX1MqVgw6Df65HB9LTeO3kkGYAEQCZQC7A2hqtD+vEEqMWMkB2I31h89Ag9o
qF6qgueLM7pY3TAfbuuof0cS0hzGb6BPgH4snKvsL52nQCZUerIqStXip2TWBzhgGuqajtmrn1SR
jz4aMSPvuhchtM5g4Yju8i9n81OHGmbjC3L7A+e9KH1UUS6Cc+dpV1+FyvFVc+da+XlYjB35j+Qf
FPXq90OeVzf0Oiok1M31q+1M55ZPhKxcl3CueaGXurqP5QPsXr5eBT3AVRCaJSfEWYpU8rj3JubB
55sQEoiHs7YWFC5zKqtVetP3EJKbwIr7I3JXM/zDNQuAQDb3rI+vv9clBJ6ATL9NZ95D8RiA9/ud
TI3X/aGwkBa3mb6zninmqzdLvqyUoaPYllUhARVv/4AxnFR8MYEawxEL9H3Rig+2e5GsrXS1XzPG
Ggu9WvJ75fZeOZHTgH7JlSXlVwq41zewU4aoRMCyuboL8Ym4/XvYoFtc/EhWAKDqPPtswvV+eJoj
VeCZQ3aKlyDHlm/v6UJ/xaxE/xX7ag9jtEqEGYjGIaPYkFk9Qa2C0iGoS4QFL/Je6chjbb+T2ovg
ks1veclih8elUaCMJbEX2rDb5tCWg7M3yhqcHY86Fxt+a0DW6qkCX8v642EbL6rvimDNG6Otr6mM
G6vznQvpJm0PYRUR+A5ZAEgqoKUZYKs6GLUK4Z6naLSJyLIbPeRzouwV7FI5QtBlV3xTCMujhiOR
cwshr+nqtCWNTE0LJKNPa+n4GOa05QasKFYNWexzXkneN2jPT7zJMuhsynXFmRS4zG/8YoVQO8ze
YmK4Q6pq/ZmctRb7s8e/5LIcH7B+QQ1OOodNPRe6JpUQ2LaBYCJY6Qx2dPMu7pEYfr+o012vT3h+
nY/sfgQqPfTlfgTPn1eqig2KCIlD8szYuPhrc4TvYkwe1nSl64+EEs/x0kiVmeAA4k62mSSEa2WP
G5gR/X5IMDsxweNRInM6AvaBDlehdP1vmm5qH95AUaCaj7x+unH2ZizUp7BHbeIMK3lSmsqKsokG
TZE/FBIVQCbS45jENX1J/pqsmv4OGuapz3wj08NDsTJbv7A4V8icLCYCizXtJJrTWdmjO76Tu/yh
NJYafJhi/vsC0TEzzw02YCIpw57C2GrNNW/HQgePR/zp4trIphEpUfmKmk5nY5IF0SS8qCBQj7fN
VorpzEShY4Bzx+GXBelfljjMxjHGOCM/je3g7tx3xdyJQG6KFPon4JcJDWf9hHLcIbFS+4cStb9a
Zf+axQD9IEMTAS11ZM2HNm9/fREgSx3YgC1xrl7WVc9syktGHsrRCRRUMqqdlBEZhr7pUK/G9n1t
7cjzD2TEygqT5KfMJCZkz1nk0INDuTKv97/MAxEiEAgAleXZjzXwVy+CTRuZy8OKGcusOrGrLrJR
MIoGgoH0BT+QMg6rcJxIVN0dccGzn+KNF+sfrtcuhThAr9YALjsZahi5dSpESWCiHR8qwGI0I4Q4
rAiAK6SNXpGqao1MD6lTk6fIYYte+6o6J++/qR3Ur/l6FwbXAs/aKRpajbiDu8uk/smpXgrD0sx2
LGirFUcZ25oHETmyHx8Ji30NoDtU1O+/xAT8LmMNI+OPZRngjPFTAWIV/oDoSlxHgtANtK7F+mMY
FKKrECpb7DcY3L8Qm4RDZk2BbzKVeopYTWCionX8Gt5v4ladFOuLv5arawT3OOqzGHfYbiMmvn0N
XvVPDlgwU5WH13z41TKOX98D3ZWhNZDSKnROYv/NRJfpfETfzrJXqOupCJF5a5GL0jZyUIErxbVZ
I+UANJGCFJeMJI/FZpaze2ITnQ03FxD5uPsOgxKRSglLAcmSRO5cnW7SJ8WRrNoLXocM7qnqRYJb
wMIPEbsKoPsqFsb00hOCWTByL7aHsMaJ77x3ot0WQbOo09VKq0tqO75AKo9Hqw+y25AvNjFdmsPc
24mCoUpUsHvhzA6VgZP5OuuIZ1+LSHthC+CDGIidyulAiftGOdPQT/bTOHMBVj+wkgChWzWClxhs
uFzDuyr28rCxY6P95MdbLaGnXLGtWclCN1mqK11awOXlT2HkNObSNRgcPbbHfepbt+Ih9fFWcF8W
0U/TT+s0OGZYEqp1d7Jf/emNy4fxmOGBmoBSficuZI//JuzVtYKte/GbV0qzJS3uX7jtayYdRzcZ
f1VmokLeiOXTpbAiriKhB6J4JVmTS0xZcfqcg8QzvFsSrOQGIOxyyqyHx9qeVg0AMJF3XfAERyob
iUfkcS9T38bJJWSH0sqU83Ih34tUUuUTKWhjj0feWvf19kD9BiB/27QWA5RPEnBedZRLjEnTVaEg
jWPgaMn54534bsizpOtWUGvLKLdRtFeI+xGBZJG18kmY0tJnyQaR1W6hZJ/tOc7fw9K0l9Zf2PlJ
DAfsugKoKNPmjbNL/MSSrRRHD/YcRHXHsWYHAmTb3OT/jBHpyR1Nkt+GroY8us73ypG6iubn6jRl
lHwLUhom+PmxwlLaWAMffenW3x97s93TijuSWQEFBdDBQALps2Jw7gCJlwsPOBf6/gtpOpdsU/UB
hZApb3+GG/57Hl1+qbF2yI9HcfUBd9uFLVBKjDcW1Wg1QJgUKu4vu6Vg8PQI3hSbH2/XS5j2k8c6
G6D+ybTB+okhLaw9gw+2nUtZVZ9LUaOpXoCxVipI74ZbDnyr4AVE6Z0vHnuoBdKCsO2ySLOQXpSP
Ksqcb4kk22X2oF0kQyHum22t6BZZVHkg5xoatYPAR7/9IxN2rXE3UEezNvtw+1KNEaQApmu8snGA
A/7qTc+mtzuAK7P7mVNOYNTHshUEwINqo7ssjfJ61Hhh+x6OBHoV7v+5gkWERPJc9Va5igTnKo/j
Uh4uc5AA8zeUMG+UJNywN/XL+5Mr8w/S6U/ZqQ6VoNwBPhR7eZL77MC0tqoBE2nrhYqe2qlniU9o
jjhGPEz+KLtGpgtBwPkxAHJzbhT8SaGqd2Mzy+ud3nMzno36KiASpkHvW9Gf2iQ6HTC1/Y0ASTAA
8SfrNDntig0ne7yxtnWU6+zQZsqpPXWRfUNWne0Xhzvwexui0hgzQZDbltb1FU0SCI6FtafPvxfU
TrUIr2d009pJZa6O0aS5DWJn5C0L5vVyURf8m9jIUitPtpkCRt9iHjKofp09I+pMubyEj6ADkT+5
x9m2qIISEIfjkazkTIv6a9ZfLcnRGoiKHEU3KnBbGDpzEY/HbWecsHmu3g1ORQDuGtu5kQPk/naH
WPaszTm/1rI49mMSsLAjFd/0hhaTKtVRbBFAN9vs2CUlZA5h31IfUPv4fK0UAgx24de9OZyltQtc
TK5Uf6OS/Nv3sLv/jftLcgabpNKeEWkUtvyXIXjSWco0NJ6Zlf6QcwWQe1ONgUGIOAe/jxdFO1mB
qUgEy9bkvGr+ilgbL35OopzBrPUcfviLvF9d2CkvOiqXW708zeh8SxiwWOLQos5uSTshqEDJjPR+
tI/HX+DkD/1pATRCxWWw4WzRJ175WBAsjAW2Z7eMzBSdRGkPyUpILJ2DUq4mt1UdEljrbCiURj/m
wtTv+Bmzj9Q6S1ew4OA6HPn4vRRDJ8eAmV2VKxMR4lHhm4lzQpdYPCMyz6d2qY5g0H/Phb+BIXFo
36fJPFNPaC5abi4KMx1WQ2gtA2gV04ZU/hh582Y+PbNR7e55FnR5vDIYBxDpja3jqIkLyGKM32Ip
ycbFmQApbefOF++cOUwtNDTjyN3GIJQzdk+dri4jUbpaYsGTDsDrd1Q/sAAwbZBa/fgC2UHnfBx0
PL14upVH2gUu4KfW3c0hnoyEypjfi4jUQ8cNrGdKuGBttvvLFwrmyntSgHOPyZFdV2usn2kgiOpH
HzMs8TlTyCsCQklt3Wi/aLonyiLdp9LPhqvU+lD4xYXKfRJc/kjrwQkMM6ZAYjLw7A5vKWDTkZXA
kPNV1bgEBxIUxZn/yCYk9b9gTWzTivR7j1WcCAUKpeKOHHqktb8Js3y9lVEVYHHhONAx5clQS/No
cEBiD5ULjQPhhlypb4gOvI+1imOSKm78d8nrcjr5V31OLrp3nNPoWKpajri+n6g/OePK3Eew9ORN
Yrl147dRS1s7bXtSY4JPHoxYlmTeR8qkOE+GKWeFylKgLwznHrRKT6087bG+tu06EVo0R4+AlFPz
2NU+NjQk+pPfVtM6+h42g+PPHvMcRhpXzHEx2wHBsMF/eErPiXfKXnYLF3xa97hU9gIDQAeuoltD
qS7CbXLr0APYzKwMMriWT46awAdkt2m/mabpZlCIeYp6NNVm5WIa2uf31UbFVVAu1nH+/HqiRgyu
x17Jxa9mzUdckm31yXBaANsVbu2BiQsnoMQAh7LNktluby75PS2wqhDB+cPtxfuFZ4ZfmEy4zFYP
EV5RyhITXl42Hz6W3KNW66hu0j4uc9rgXIwyPbyzDDktVVNTOXT4ZU/VJKSsTfBY1EsL5LxtaCRj
HzO007NfgheoVtCOICoDJegR3OI31/MCSz9roHAR3jZT6YRG3D3GgQ4sm0siA7vkRe+NaUKzdDg0
QrFHz9J/9JM+L2BxVTeKafwEIQx/odLy3Gdw6DOwx8SLTufwYcWHUX+h6WPAJkTp4nLxwNb64Pn9
aKcrj4DlSD+XruJU1817XehvVN2yJUv9yj24hgghegx7Y3DoH3vmfy3dJH2PW1WJuoo752muW8wU
sA0JGJ5O6sn+gH954UzvRDAtGpJIIwLAfz9Vo7f46EXRR6G1AV4oJygtOO1VYZQVRM+FRszfItw/
tuy9lMdENyJVYSWQq/yJU/lsQhH8oxispQBmBHInLhc/fHQMBd+0hmT8vCSyiDy8lywuHHA6/bws
Bw/z8ju1xT5+Vny35oFMVVqHkNQiytY5mMOw+5q2JiXh9j3HxqmH5vI/i/lPiCfPyehBFjIugmKu
bpIK7iwzQuDThKcgEANn7RyZBVs9xwtQ2KVVKKohthu8oG+4te4klyQY3n5Xfe3DQT7q5ZCCZtSJ
eXpGhs9WHWwarRw21ylb8PrAMJ/2RbE7jJcYHaYerAlgk6uQAkOoPwC638DSZKbDiSEYyJe0KxWT
R3qd1ZrEjuGt8IicI9pmTMfH5dmh40Y//EQjh8dbo3p8Xah6RNBIdPjm8lY3AY2XEGOkfJH70AcN
sk6v9mROFcGebqlRysXDqm0GpmddljMrYrQvYU0ldA0Ctflmcb3sSS5NDZozxj5JTbBoTHrum7dl
WVGIYTnm0ZhyhJzisBE8OJsnpWjDo1+Ka/3MIhsZhNasaUC5a3rYpmPl5MT6iRXsbhZ4Zypoh909
Q8KOpOJb5RDmnVUzgncJnuloxsBNn0fP9vHT19zDQuNnpMYTmmq1eE3cqbYf2/RlSihJ8stnU8OD
2BNfeCSPqTrVi+u1/Pz4YZQ4WJsAjDNa59I432xt9cLu7NxGsViX8FHvWr0x0wMsP+UhA0w4NFnQ
GyHAiDmPwH+9BT+Pt4cwKHq8NWpvxhEbRphtbMf2HrDQq6UyXqIbvTp+daNQQBb8ZVx4tESBkjq6
VFqrhYmjUvx5P18WSshT80tvVDTkwOdKL7Wl/GN+HfKTPAzoTKdHTSyOB06rwqqHuL6dhD2VC0g7
uEaHIfGfPQza4lV1R6oMRyigHM07C83AlIdIa8LXMc2WOb+8t2zv6/wLV9bPFOjnh2Gr0OKpjcEN
NjjlI8L2XCotyh+0vI6cfLoPP/VwVZ6vxcucWY9rz1bYnQVqfaIQ0a/G0mbqHIcEi0uO6rXEke4b
RtvkEkKNduttb4HDkajRwhzlCli3wKawtSTdjjqF49ZPGDnmX8RAYypYyeC+or5PCZMFwSctDJ/a
IEAfHV4cxxzGuUA0FEXx3K9PljPhVRp+gw2ETIyYTwCGcJTnclEnGBf7++qq3XDG7+y5jU8JwVmm
U/h5vZhZbVC4tQrUUZlb2zuGI5aHnxTRQqWkIJ4eKxehGXWrz6dgPWMdPzeHbGAq3fqi23z7dNwK
yY47Dk3491dVMDC2H75Da7wj7xkC4QcguJJk68gQxR3QzPKZJv4au2CUPWhpNt2IVmal0ePU3O9u
3WyVOCCxZZ9+3CKj7XSGsPa76u2nWy2ePAboFpoCia0Q6ocZEtxkqx2gk+HxxYqv4CD57cfr51Pt
0cy3fTd4Y2YjXNi63QBR1QJAu+L6c6kgE74VFWd0aj4NREyk5cpgmgrivvPtS2Yf000OkUxdtNo+
/i0TJsD/h7bAWq/P1gZ37kXYe0M4EZxi+0Bxg3wKLy3QwY+cykopyl4RO1pxE1TXP0rukt+3EQ+3
0yt1kQ+swFYofHwnYn14yWuKtZ9J3cvmererGal8djRsx2p3hgDIjnoTVJpgB2o9ZPuElR/se7n1
Hzbq5qk546zjTFUFMLSnC4hNzGw+IW4OXmYx+An0z2ZOoWhxwuNGdfwCgYg4oLlQQhgHs3degIaO
r8XlHJeifmLR8dYJARjax2Sa1FOB7ahMFysiGk67ZMKXksB5hpn35S+Mfgpin1PSpAUuGH80gOJD
3T2kOVDJtdXCfnJvRW+VYjCh+AlU1oNoTdXeZfqpyqUE7Mu37C/w+Zr+OgK7q6Yy0ET12HV/6rFi
IVXRiWQLwflZft2TcdorE7fxQQzo2YNrp0YbUsWXuFAwmBAj/6JkJlDdMXiybzjXBGgNG6jgVfQs
EjMMbDbOPQKOSOZ7wdJl231dSvhZ5A+HIASI/QBfcdig6Ph56pEYm5cWoibGuftjOM/ckmhwqGUk
JMI6XPkaecqGkijhDjMTgnBQLoVjEKEUb/yXRNziYMWbLUHPKerUZeIPF8O1GY+4FNjYb+XL1z3J
E1QFE/FQPEUiw420dX2+/mmrIlh5MdID22QmdiDKwngoRIjItTUPI2wrMefq1DQOvwcQb+Ma6U5I
uTn1VVTvpA144dXcefEvVpUANgSQ0HllLeKxBZEyjV9dS2KFNlIISY0MP2lcNx+Yfp+G+HqXlQem
qocuJXIxEAHlhI3J5USJiufFfC5IBGOCVlHn5lx+58zF75Lq8gelfRsuIICoSYalJVw2fPRauqCo
wKyhAglS2oBVhWN6KToZFTdRM5nU389ztWTabFdjyH4ycOHHmJqwRH956c3z+h0Rz09DGPmm6Oa6
p/h+pzmOnXF2Pvy5DZLReSS1ZeT1W49XZiIyyfPo4N2MSFbqTs/LjqX9V5Xfcjd0tqCCpU5MnXMa
xqYwSUXmAq0SBHf2nYY+p/LhzXCV3QHExAhr7z2cxZEqprjrN0AaW6QL7TKTEPmc5tXuzra/wLe4
i5wlAplPF7JmShNULHGilJPInDOdVuws5MeiuxQ6NzduD2f9Dk6nng+GIhsDrVC0TUqVYQC/utmw
iDYxVzH3Z+gJAK13Um4EG6PLYGgpVPcjtZbFQBfQsbDuL1clLKaSgR++Otzu7O4P4wxYxSzkkT7S
ohV7RNZa9WRtJHjBfvkqSU2iMApop7a9b871aN+LO/RH1lB9D6iXZHzVF+pTbxzQ8VdNMdcDb50B
ugAJ776HwonnPj3wGfGeDmIheVPxvF63GIf2mzuIbq/iUlUvpL29wlausLMDh4RiqyZHNu+umUS9
t21qc4GMpnhUBA/qoxNCRkhy/uD1HkXMvGbKPrKTJvuRp4EK8/2bTK22TEeeQIjIK90Dy97WZIP7
USXJHVoyc9XyWQA9I7dn9kiEFUFSNMaJt13xgdXEvMHf+ax0Wrt72RODD4hRRn5wyuZhPk1aboxl
ocq5wY2ROjmTTHkmF1JS+wcEgXlJ+SNjkqdyt19QFAJVaSElCZW1NN7aliN5+/UbvNTCXsh6XVG2
M4gQe5C90p0IECX8TvpUS/5pnR1+2Td/qGb/2zMt3m7QbbBROwMJwIafttABvdozSICGwAUUWabl
lHME0wuMngK2nmiTWtFe20jLIkW+3QWVRRdY27qW+/fTCJxmiH/2Y+awTt0wwLeoHFRiWu2k4jdN
r2X6wmQpJG1ys8SHrqalSwcY4X8b2tEiGF9bK4ZvArPuJp7pG4sY/pGP8S/4kkqkB0nLwBqdZnC2
oJCw68ZM6uDDRuYkAbBzK31IcKMnbocig4Yl7ZQ5Fg/FqGG0TlitmFXkqWY561+Eamx1ion9I9B8
EkBeLI5V5OgpjZffDZjl/KOarMw220XTLYDYCb0NRIN0Kq7qHHDMSKVOcpODOpTEXv4ottt1+vO2
ptcmwLxlm8sCVeDHjKlaZOvEJ1XluaeTdKcT5LVRm9JAvnsnYdhLaw6Kabnnoe7qDgFHAJ3B2+hc
zaWdtHhTIGRJGuJyuermpidjErNDO5Hfl9m5RSb8cXq/W6B0GLs1Vqsa1/sl61oX3o9Oo3E6aFjS
sR9uIvy+WOGeKBRRmsWr/s9d4/b3QAWagOuC1/Q0P+gOoKACuRJuyFbIubHR3gxlGWNOIzLWFiza
2l+OKkfjVWanhHkv5J3kEUCngjrulVMucQo+LhFZ9XZVNddm7uA1S58gjlUnl7Jg8vRDgiKHkOaf
fm99dSaLTn/iOgyfAcB5vk2RlW+N6vZvEvWFFxTabfcdF122rn6rJesUERto/hH+oSRYz8INd1ce
gCydE9KnTFJ7uepErkYpsOoHQpp7HkKRhmoS+M7F8YFeC6/rjAcbUSIPYipFRoEl+cXvnau+3Fd2
0cV0iDpBLzs8yeFwb9wHJl3sKimt6zD0jm76YjpDtTSOq2yGnn/a8ebISSuxHZvTJ2k210VqH6sa
mDbajaFWGWLBZSlACpGIgBuGUD00K0ye2yuIu7mnBFjHHp3nyVVc8xKN0qKdFeZiCt5pKIRajzB/
rRHZP6CFPyGoll8p5CtMcMAOyPqUSqhtrCw5JcmcXBNvIRmjVC7Fnifnv2xAIU3kE9XLJavKyJ+0
w0nYxi3O5vDZoUlu9yWXA9xt5wBkHlxAVOpZVSiEncx94wRp+UQKz2acgKeX7gEaFHO8bTZ3nJxK
LmazadNXYsP7F3AU6LH64hx1y+/Aj0wVUfO66ScImj7niTQ6XNlqxH0me+rlWLi4Jk/iEX/2q1H1
GUjLMGEiaugjyKmzuN0kshQlXmttaI4YzOteZd13Su6wrmKX56WRkuHRpubT2MlGClgY2SL8k6i1
b55lFq4qWaYa2TNwnr1yMRsmZetlZ6vUu4EDylxOZtY/sQNDkQNC3IEi/hetv3xUmvSEYXer64e3
EuJYyzG/1fN2gpZFcPzH0UbkavI37zmxP+HIq+x29Vg+y9ZFndTk8N3swJg2RZmpmw6br4cZgKW3
RjmW8LMEp6l+FLCEKW30wxRF+avPzSjiM/GlKtTYvxtkTZCxZiAYfh4wx2HggjdatCYqYGOIFD0t
jueXzixEanckMclnc9qmh3z786SoKcVawHwDkhquo82PQwwzoKjEpvy76EKFB4Ub/MEKlk2Fnlgn
INBRvHSgLniGWnIu+zXgGc10a8RB4ll9oQc9f0gPOgbUIPRLcY71/i4CraoChbQDuf/cQYvvtVzC
IburaCxzUTveqyx/tIInWEvIP9QovAbVnfbJuRt3SHGmBsWho6Aypc6xjG7wlh0lkDZZhykKcahd
PO/53ygDkWj0FbtV0XDZlKvD8xrW6muYnlaRsy18wlHldZu+86wOmyC2d5PcP0NtKnjyFeza5gy2
VusaDJ1AzEItVVbs9cVE8kaSxDYIpio7te8bU0Cw1zlgeMaG6T/fyI4knYAZD8d0UYY6iRpZDlDR
+kwBYWTGdiz904HaKFmLj4hYl5nmnlLxu+5vNd+s86c5ZAXJoLtwm/Nc1CkYXnoHkal2wiHAaPNa
FxnCW0Qmwc115iPp8+LkuJJt71GRkH/XIxNpiwq5gbrSaD6h6ta5vKg9qCClqwPQQq2vGsSYF+yS
HMqa2ipAZwdAQnOXBf02hzdkLdtKQbrpVFQ5ytnzfdHfmNtjAS7hRMQMixsNxKofVQmVrNvCRmee
gemI9DopEmqovOG9AjusUfgEh4tgDxjv9y7Nbfy5OlrEYAbfuesR5ttT6UU4PYqMtQo712EMQpG0
Gar4crvGojdDrSDj8XcFRR24sD+wdMftgS6eF1aaAkVuYRlw3zwBdt4/6j9EHZMugX2HItCYizWn
AVBoDAarpS8n9lQmFx4nv5Eng2noZ8j6Egn67PFjeQioA8YxsePEl8ltqjwbL7eEdNTXqMsaSqrZ
Dp7qsNdLtwiVXAGdX0QiV2FWYVyZX8A3iaySNahshw9hiiiaKXGlVJQBJJ5EBHbF7VFLF2avZFIt
k2aUK+fv1Fvz1ohI2W0DYh4KG5l0Y9oHZeoroMhwqZf2n8bzRjSfhdaDmGRBYO0MFh3T4ygSiLFR
IufEhoyrJoBMpBNCrgfNvFNXAwn7OmhYptWbsdyvp3prKeFoTYLosAHLdLvsdvYw+qtWUlWEv89Y
dFu2H0UxY9fWjcTWncxhLZFl+hqJ/imonktD3Z4LjiwZMY+Ix8NLF1XM/4hjbRG8/DS1+K3dVlvv
ym+Jb3R/ZzoC8ich82bR/gt3UJFkYiigwMyz2Og/7h8uV8ajrD9McWbNCEmNxazYdLOJ0cHpKIO0
CeHSRbzwN8wASVRpHktihVNWEXJikmPjHYSdChy1WIwq7EjOPHRP9xIQOqOPCMP2A3WEUCPnQpnZ
HGqgK6IX133He3UB4NApa7R4UtyJqA/a/51osOUGC4HDl+yqpgqBC3EeD+hBOPPsDz+DbJy5moI6
BKu7krkYiJ/muSwNd2q2k1ix7Azra4860VvRbqnatbbfgbCBIEz4XZggc839pTCfqcfDEm4yL4p3
iFBEPERgGGetl42tUrg5I6OSbQHlp/0GJTjjz5JD4pv8L/T2LqbCIB9lV4wszRYbkSZorM8ThEnP
DOc2FBKbVQ5ja/u8H+Zt5JmpEsTDFvye9fqriMRAqR52XsxwBwFOcAogjqikZ5p5d/DujTYwBrtO
kN88oVokVrCmzxpOOORUETefMfYjRq4kRVlQZSAGNZ2eqOE7fEcNL/yq10YsFv+IT9+aQ3Oc8bLz
/EYgfLFGHecaebffb4nV0ICfMosl7bEQs8Gj7hV/Pfp1XjRr0mBWU0yYmfcEz6ibojErCScEim8x
27YieSfICV46r6urZGitK6dmOM5g4309bSjKcMWvsYlzWkGPkamBZmhHMHUAw/r6b5HcwmN5Dpz8
5p31PLaUdW2gr8EfU9V3JNFgcUt6zT+ohwYni9tXPsHeEYuP0R2irqmf48qpidrrfPnDh85SO4N2
QuVzXRg2JkAzN8BcM9gG23r51Mx5UBdkPV/F1jlu/syBPDXQ9oJyzPzVCeqz5TlfOdCM/K14zNf1
2X2XAAbjzhpoYOaZtkyVFREOyj20ISTdl74kKHSOs3j/YTm+L0ZCApSHdqiH/gyrsFsYnoPVEHcX
hTKKPEonP5z2nyKzkBJE4YmDLqh+Ye7iqqIhwTZk3+cv03XynbNgUoT5i4Fq/gZ89RSp5LDSk1PH
nj+dkWaL+vkSQfCkK+P2/TQYpM06k1pSqqSsdv1/qKS30yY428X1rQt8LpnTDzop2pHLZ3gJJMUB
7ObHekDDrmg13k8rpkrVcw8fBpzpetC57P+cexu8xjWtTWcDP7GvM5nAYnjFW9YMQFBcmetWCnBU
RzslMO2hFhuF10SnBULnRqOR7xF0ZWky8CZD0801p3VWZdeshJbJPl6NgBaIslCdu+ryqUxBQs2D
j4MHcjJZpSlOS48JDSLDz71A+Bsd5o5C/LpgmKEQ2E+w16hr6qAJPDbEAcWPRX7vKHwAmagzbyEY
27Ghm42jnPAnF5w75KjetFtjfgNgz+Z0Rvm3/oQnTJ/CinK2iiiyJis1NhyHmElbygFuG6aiTS9N
eORBNv3J46XpHOWV+++otqHhlEA2JKfmdUCXoymKPVSIvaR+T4p3MdmLsZ4gBkCccsLGfDm3aZPU
6aHnK+FOBB22oVJn4fXdrZlP01bwHsGWOV6B3Uyrc/t7KQs+mOG6pnyt0NolDkoU8UfdjVnZsN+h
AJiDzgG5n15umv8sq970O+wVy79PMWWNxNQBI/w7sJ1yud8qqec2+nbssocDnDQ2nPqP4kxPUv7+
bAUI6EsL4cTfcrPTSPdAZWheZyKoNeF+JpITYjbzQ/WXwVY2zmfm/egcb95S61S2E+3EP2Hk6boO
pNNeTx4QQppC5sArWoQvggGRz/6/2OFEYSDsacvX2OnICUQbGeJv++XGmVCl3DOe6wTo3G3h2vrA
pC385EkOmuG+BqfM7xdHdrgPjDmpXotExJRSv4Lxf2GxJXtjYO8pXSml0DYhX9vBWlN+Wbx7wenA
J9ynKpAW+Kd9jdJIe6eX/u55FBK50SncFeK7mNWAV3hfJP+DHgwmUaY8GQanCBb6+x8eJ0gtdO5r
CYwludON9ABYrH6/r6BIMTvtQ9qKTAjhp0sykXwBlwQwk/ncXtOkJ2JF/Oqzx0aWk4srvWxy6kBQ
CG8+8NVyEA2mjpFoikrwaDZqg03RdIApC3ndLc5FsypDkRpm/+JbACAuQQ3n8a7DaVQtz5bwVb7q
yprNR4TVu+xohOA+BsfkSvMaGJfF9HuVMbEO67MkqRWXPIQFv0vyHkkkVJ4GM9hYpfUECbQa+6vN
l8Le/tArFaGNvBVziBfvN9Lfo7ebh7AHdbex3L8SlWBamBMe9wcDnQocc/dQ+Lls7t3M6jc5Enxj
xcUDxBMDOlsLuO9Ja9dRDPzK0dzTSHfmHDmZDWYLaJlZpgr6mMfzJoLtO2e8eENvUzW4zGw+l32+
x0FZt06zi3yCpE1JCo62tDnJKhRSLxgnFcgOrdrr/Y8SnWhytho+eNycXw5O7CLHIb7cn2H+H6IK
F6T0nYE6U4WVDOgUyAbOv9zFE+QS6eq/OVZHFJJcDXvasPwXlHZEs9rCfQ+A2vGVKJu0D+CMps2U
BZS4OT9k4VLl4GtE/0oXLQfukGDB132oLvrVnI40qQaReRsZ5I72czMMqeyA5oa1PsFasEnEECpD
6g25R//RnMiBF2Oof8F/OQ6xtmxRwwd3di563DSWMA3Ix3GhALsnT1HAYt7k412LHuFv+DxX9vXi
o0iBCaCl+Pph8AAwh2XPapM1h0qj4YQSx6pJtdwIUdWiTMxxuPWNuzYDA9r1jkrxnS3SqfE52kef
YN5WHtA0Co6ZYCb37JIG2yIW8PL+ps+EGaOPLLdV2AhrQHFec1t3j6jtDxtDqaThnE8yJhX286oL
PrkII4SAxVdj0hzbdNA/38jCsJoI5OmJ5eE2JlL/iM50qHMVgOkpTCMVUGm0BQ5txu1S1elN21hx
fTo3khCuSjD2Ibjsa5up4B/78tR24UocYXpBMCTW0f1dgGRdAt3Opm2SSBbdI9AgcCW5YwAWeA5z
fn8yio2EKXmXBvJ9IvbLm5zGW25UOykhkWzfBEXi1s8+UNC6GCBJh8LqpUGCuY+mnP2tcLyljFb+
TzsTluCLriulWJHL2RiZD9zYLi17iQ0yp5/dCpJzujVSR7O8eo80ClUGNyVtqGii+Fa/5npvvg8I
KJ9cwAbxP/Oim+6c252pK56KKhOzi8lw/knrsJTWWdfSIwUdsOstbwhe+WDZEA0jdeqXe3pNHP4t
UNBm2RmVTktaFMay5Ioi/MHWVOy3lOXM1nUDQpkRKD3tV0i8dFTB3FxvAvLKqOMKwxL6vvqnkXkY
zxs4ZSdROBId/gUmUJMT6w6/qY2jYHdNaA4vFkNJ9xN3HEHhqb8ZFOOvIEcDugBaiOAIugEoD/zd
KZrdJyLPilzBl56pP1KJJ48SEHQHiyvCTgpjnhARsgJnMIxZ4cnR956H5nA6fLvvk/komjrjLuPF
G0kxfSrzunX6uTv+VRXppIIPReLqDJqcbcKjvv0SF71f9zenxhH6OspU1QKjKAgNteG+PyHnkbtf
e114kpEWk8y2ZqHvaxtGCtK6XgJokd+AJ23/QzXj/031ZqhJ59jGDUNkNr0yfNvSTZPBnYYqhqIc
KJ65FT6Yg+xwaSHWOKF8vZx7dh4UW0ix1SL4Gt8nzmUVL4AiN33gAY1NF1hdvqygYqT4NISFJIrd
AGmR1GSSfJQPxA/xYXBQtxw8fEIdVt2n9qM2tWKfuc2HWLBPCz0jMJtyL3516SjeDK+T+YM2k5pb
ojW/ak9myzA6h/1dcjDWP8Ra066JVj6tPninyAQTd30mNcoRDz2Kl1/rtfF5JuvIZe4pvxxNSaCW
ewmkKp/4TFNU+fLTqkZ1nfWVBR0RbJcxH4caueT3tHSdTLh+QCacJJyhjxsEWL6wiNmKdcZB8yKm
b189fceXEUIc3M3OSWEeg7/M/3cLx+1wf7Qp2H6zIV3jCmliThCg6R6icDfxaAj4PBMJ+qvCkGWA
1s1kALGeE1E46nwTWDfsyEs0BHJV/w47wau886Pw3qroFI9cfRsU3xg3HJgBE0F/I6etw73SH27E
ek+kNpb6j22StXXABznhxDpMHP1aMlGbNwBMSNbqOmxNdpvVlz7FZQZRzg95547XXz0v4B+IfPvN
nBzGOzVWDvjByCG7qgu/VO5inQYx3QgQ3roTSfECD89mGgcohx2WMiZHj6wzPpUQIl0tI5tSoeQV
hgg9/Da+b/tgh69aN50+nx54oUcwAnScMO1DfVTKcrwJ6OGOY9kmd2q3CTiyZcKE44TFmL503ukf
ObSBj4Vden2D/+6Gnv7VVj3Z+IWdZ8dSTnQGhpbgHsX07qbxvsbSsRZJYYHOI33SddhCrBNLqinB
dXg96Z+mJqAtrx1n5o42VDH2X15nWcHGwDRuV3xG5FfEXz/Lq2KaLzhCm4weKx1DpaBhR1AZQwVd
htrq3BbazD3MPMLOnUSV8QAWmINSkXbdkzbajZDV4q5hjn5sI7ARkSmTpW8L3Edz+uwcemuyMbRv
mGUNPyrzlXrDqJ5KHWkPHnuPD+z+VdOnHMG87JdsXDYfIvgmTUoo/1SZa1fZiR+8LqmpIblPpCJF
i8YRmPJf7HQ3RNz+lrlDo4JYfcN6kDmBbR+Qijlc1uPqJcwRgW8HhH60dhQ8K56tQxgYDNbUvH1F
Vs/sAvvS1gi1jT7XCB9LdXo9AI2VwWDYGYRYPurLWy0tzmr3rE8izLqiIb9dm2xRMeotZfY1OPmy
EfZhkn+ui6A+/iMtUQoxEA+Mps2Ls14AH0hCfYW9oC+BlWyfryn+KjjRP1WN2SinyL6okWB4wnAZ
9GGj3vLe8EC+LsLapM11JbKq47jhstzk3sgen8XgxbLZgsUYgrMYUeqJFh4yNFapKVCvq1gBqqlZ
a8+ioWtPQsWYYtnnJdzNMq6LPjuC3q0AaaRRfzSSoMx1y6zvDYatB7i69GzKQNY5E6Of3tUGoBd+
H77BciX+wN5P8zcfw78JlkOHkJFR21OBdDdshIYYZis6g9mQ1fvVWTFQVReQM4OWGWYOASoujp/V
A/aXjkU674LL+LDdwn0lH0HetlDB0ZK28raxMOcE6yc27TOTzeQGgGr9JgIiIumGAS9E2THYFEUU
rKH/Z/TC0ooqvAqoJeIvn7EvY9M+z2Np+3Uh7Wf+yX9LqQwmvxBPg0pG7xBBMDqITJNnQKJCRksq
aecQLfzVsnCp9XcQSzz9ZUSvxk40JvlsembfWI47MgSbIQVWMRW3fjNHKCrbBEH1sO/qkvIAROd9
Gc1dzFI2yOu0tedubzK1Y6DM0VUCdg7pC/Dx4TQcDkxv/7KMTmCiXc9RI/xF76nw8FAlTurWXMjH
ty0LNxYW2psS0jcVwbbgXbiNRFZX0kw8Nup5J2e8MdewYjVIUw9OBkHPy11zw73TrJNRAADyeUC/
WgMQMUDs7aRASCeC7DL9f+6JKsDHED4gQwVGJNreRO88PU3gFVERXD/ECnYKsDwCyts8xP+JWpbp
gQhEkr92dndYW1/fDTaF7uKv0oVla4Oh7/gJv1bUNQGP4ztRNRiawUYE8fstCovSBQl8XK6HJFvc
toZvUDfr99UsjDNihmY8QDPoRJQAHNGd7zk8rSGs55iXCwLQgf3FI3wG4j0dcGv3rRLd2qNq7+Eg
Yl04MohFUPFgkfV0goTeD4GwgdyxEEPsPrSZ2bv1T8RGo2zDRtWYsqtEVhnbdUEgSCJVqn2naII7
/V/2f6n9M37BrZDZNq8H2mXNBUDZGOBmiX83lFmLVYBlkm+1azMqKUIhS6PymO6LPANqkambTi96
4FD2O+Rsj9s50KaAx4C5q48smx4sz/7LQr5ZnXFyfKSyHEEj1tj9e+kJUZt4P0hH49wb5d2jcl+p
wIbsRPcS2bI8T9x/MSsPusMpgpBJ0P8mQYqBk1aw4nM+NGw6tS/AneMh1QfuXIj/2rTjWAEpwPkp
GWz40MBwolkbZB/su30+SZxQLF26hYQN6erysIW/7amppfWxnAoVRxWAZ62dsCaf/EqKCRXF6oOg
rCLUpUbR3DS8gL59C7GycEmMsOQwSAYEvCMq/9iiaT8DOERg506hJQ6m3nOg6T/yNIDILD4EhmZe
EbZZNDDkMj08t/61njjyHz528Mzzptjm/eDSuxJ17NOtfiz3PjPA8unFOom07mAUYFvkclDVg1/U
lt8a6UHKmxBsosCV801HiievcsL86IG6vrq/ccZevkUCN4pBQCQy431Q8jm+jjFdMSbdPSDJivNp
E4vmHo4T7KE5baNgWWKpey3hNm7emZQT36Kf8NPumDKcxO48dLYqFY0xJAnOjTgiZiQmhRbWJQaf
3mIho2qSPSCTT3GyL8jzwmhdxwwasyH2n9Q6iiCKMVBgkIW9uq1SZB/bQEiyORaJLkmdNfAh7tqZ
x9kaGDuIOcK2jmQD0M8ppuDY4fAuFOeyXQ5VtU+2ARtX7JProZHAGo0FGX/VQs402mynEis4ft4S
EB16v5dMM7nln5/IHp8F84k0pnLn5heQVM+GxEPuOsSoo3VKY5hWfyyNoGYZ8ne4E/jy6GRLt4kx
GoxKw5RtZ54it/ZcKPoEh7jLnA5eXIpSu7ApsMs0vmL+mbZ9O6jWuLgJg0Ik06GfdOPLd5vs2JFl
JUJVlFwi02pp1HcPWXD9A1Gs0lXn1GDkbWBmlTaf2gZ3FHsFfRBVKANrEgWCKuMqY5e2VBw1ms/6
eMrvyyrSJUrcCeYcaMfKjAYr7XOVFvheINMlIepFTFKI9SFkmKKWNNMO7KBsIOgZ/HSlz8GKxSwB
8OG7kghh/hRjOiBzpmDmGhDzTlHIWNF/2uKW0aky0/BtaaJdxXzTtqirw2kuYtFZm7yG9BgeakLu
gEWPkZSsq8hHjGGouoYHYXjE16ZSsYC35mkLiHXoI8dFaBq/qrKye9KU0D2loK33A6SbWIT+xH0y
Q59kdWKBpVkWtkBrY0iV0+p8kM4/m7Zv3ogQo7qC/ZaD0V71oQlgdwWStHTANyBmJT+LjSC9qU4m
hA5/JoxTVd/hCHXz8KvQDAned6rnhrk+PctCVqeLSMBOayyhRKMkYEBjIx6GROgHr1SAyz32r7/p
fiqKux5zXsrJjHpxDXsfEx4XkTCbkTuXei2YdbUwUQrihHgCqboraC4a0G6xs9/X1eGsbuj8ySZ5
Fwi2sVT/XuKPLYAi8vdbRgPLVYd4v3IJIE9uuaoqdbKduQT3wMJsFlnsaqTUoHQXKlkk1RaLXBm2
/sJwAY5WXjOq2SfzG4hLs+Vb4uG4+OqsA30/QUlvxkr3RHyQDdYPE2GUJ6vr732dbbpDfIAZsCHC
cZvasWwTmVmoBaziZ2ajJST+baNaEpJFnsNZoJd8bt65FzhamqsYUPSHqKC0BiyakwIagrCvPh5f
5zOMT4GXf3M52SYoG/+tNDpi4FXVDmlF9SXhfg4TXAL7CjL0uxYqHaXSE3+iD9uLHiJ+Hk90uLTM
Tmf4SQQ3znsUCWEkeRKsCIEaN1lm4/F9NLrGfnI/iH0WL11opr/RhVZovFeKOvYT0zp3HVAJhywe
0xUB8ux5s5Yo4xLk2Y04slQ9Fq0ADqjHlNT1Y8NoM5I3QiCXxHFEIj2dxwwWHzv7pg3956fi/GD7
0sUWQZB/oZI9SudRtxvaXLr11wlEDxsjSh6u7xLCSvvBdS0PXX38gYP6aquw1zOr1sEdOXnnsktN
pGa+zgSxax5fg8JD3WmUUlpUwC5n1CFmkPP5vGRo8rHTfOXIYne//9yf2QIL2j6o63baGAiJ719R
HOwTJ0W5TtRuEeOYkN6C+5Q0HbRMOg6nh543J+DDgLwhWprlMIiLwcYO3jVHbDarlzA28OQtsqKD
Hvxfukps3864+eVIu6GouUMccmeDGFg+Vt+csnD3MWXTPNzZMQQHvkQFh6SADoI4EXBhl399LB8p
x2wZ9bcaAB0ELyjMhzW+nsBTKwnyi9kuUZe3kP7CnyjOhIXAjjP6Dwx6B55pZIdDTmF5v1Nf5C9q
kBT5uujaCCPv93apauVTl2H9ZCYa2IUdyLBn00NqDUasTJ9mEJILTRmHTp8bB8acXtNVEAvQQ3cg
kJaHxrZQSIR3rUGLjGXV2CrdMWzjv2XMu1NqJcgeW3JKGpJxMa+08Ycqrua+ApX4CQj9UK6hO7Br
A5Qs8Isr6rvAaMkvhnodQQDjC/Lut1Dltv0ccFXB/TI6IDhxJr1l0+QXTAJSpilseSDEy1OwpO1V
FXpY5WOMVX/VCwNjmZKAm/IoTE+Eu63W2I8q4L8p0kCV2k40IpRV8s8ooleVT5WKXWtxsr3B+a6Y
NIVmOKavYkbhLFTOiYRqMG6cCillkMT543Grr/30ojJsMV31DUHSa3YQoEgszIZYRuAQ7V2hMbjq
smnRuBN7E/HNw3mBK5cqokP3owLdXv9GbxT2OGO+Fe8qD5I3xApIeYLRZJv7MVytpjcYhL1ZjIsH
SDkhfvT2ETo/NFpFnXa0FvQvImbT+jlzVtb+2ulkXXMEqTZG4u+ozrmuhO1hKpfCev/hKJSe/VLk
RYrXdCW18j6GqSwqMD9P46BEDJp5X2HBkGnzxS/j0T2jL7AyZvV2LsrRMMHRuuLFsAxmTqsvjSxj
b2zbw941yeQCz9JiucH/pJpfD4kK0GTYTACDkR3rozGi+GFjpkPt9AsYuUvAlb40DUD4RHkiLP3I
Nwtg7546X0B02Hz+eCI42zSm4tkeZCqZx+he8Pd4XvtsV2UOxoPGpkDDuo5rMLWUdchv+4TzzJQK
b1fMR46V2TtaAM0Qw2/CpZt6RT0JtToGW1ceARnRNvzXUyY5bqP3hli3MflBE90st+kf4pUcUJWz
9U8F6RSmyW641nxjwWCPSNTshEawtuETWGSNvGxT1WBPu/cZcsqepcfUPfznNCzYCObeUE+eFc9u
P7ddCplEJNxcY00dJoes0XmAOR8luLTVQqvMoBBqo9dWPN+b8YFpj8t/Ejw1CRgUjus6YrcBRGNP
0ldBfNs63kibBbt9pgAOQ86cxFMjbqkWRrE1TFIN37EYIGZjhRLFX7szhHBZFGlMSjKNHYyL5eWt
Ti7FMvDqnQjUcfhUy1ZCELyjCmq9CbYxbJ06QU0po2fO2Q0G5Rdfs4S8QpiFWGGK7Az+jZ38So6R
VssZUb2F3XZKmXBMYKsi805aliqVaGjMsMsgSkw8vZi7mOZcLSw7JAbPbJEGdAlfeHBGerFNw19D
h3pmBwVI++lrp/FZSACYNvPgKw9rTK/fT05X4ysZgMm66FSn+KX8KOjCNCZ9EeoxvnlviSxcM7mu
N2JC0jadMqMR4W5AfUfvkEXzsgdOcviMADczHknyqYazf/qQ1hMNpJdg3NLI4FjdNvdmn4V7xqOT
pUeb9bcG83GE3BXN1BlXhbHdHvJ0QgAM+vX3l3JWno4OLX45uvP2w7OiEw7fljmH7A9RWEUtv4fI
vxHsJOVJWIzKyyIyuH87ng/1ut1v/iL/qe0SvPdv0p4cfwWc+SzVQNvLj3CznBWrTasF7b750W+w
b6i7Fa4wLGfUPtmk2lm5hf9NeyUh2xwo0E2PEGjSLTw9gdy1qsN+6WbOC6x6wRkHXXIHW4p6mV+d
BPqPZSev5j5SM1anpl0LQETSAVS8fCquL3Awth+V0ql5Q/ELQQh4olyInbkIomRIrwAAIqBF6FGw
jpQSxYBEWV6qMfioWa9kbE7DeW+hFe8/2GuKygPZkgHSH98Rm77xlUWr1gXwp83d0ZEUidM57S8l
R2VKiJyz+PHPpFuaHcKhJQeH8ls+KKWZObAzy+KbmoeUvxSaww8QJ63Vp7W+FDFyrEQgIzLf5sXC
NBf+ZKDLI7+ImfyjLqhG1Pm9ZbpC7GqIPH0+4H4FVFXeK0zagQ01dwadai4AdAtNaJIED2Pyk0MK
avoh1jOfogdMwtRmqAoCSt/wGZ6pneXP4KMhl58hJLuaapF/R61ll4qgW7sJktbdRZdHiMEJZUcB
cPDb23MLrxg/MKMWaep2dVZk8D9ZSjGfJpRbHvUmL5dcdxaDir2523dWI50I08uFEu1vthFQP79y
HdqI4VKfegmJVoBGCJcbg1AJnR+u12tYISRLWX1jP+ff8r3lX7/KD/5Oju1dHfH5qrcUPp0pTkuN
VG1EQ793hwtUBye2v9nbD6STzkV+9h3RdBM4XBVOIzDKgcYuz9ptFSVtMnUGZUQ9Kx8RXQZ10BZ9
z9a2TEQCnDYknctM/lUIsnGH+eP7I7w2AqON/NwtgSQT9sr0rxjK6/Ti+koxmdD4GSnp3tHRY0UY
/eIUs8o/HqLLVpO3qzqdUSip25HkdvjlTX+hwnspxjfxnjcG68/I+8/sdZXSBHMwVBWuWMIEW+3o
ebiCrlLBXK65VWfFZ7csZHytelfCv+qoWyC2ui9gK3QKBh4YahhhYkWwbDRAl+4ei0AVJCV3f+y6
LTmIfqp+MMXpMTMkT8lBajgPeS9Js6xxJ9fwi0GSW6S9zLfe4n89C6oF73XCS+offg98dfpHRizm
PqwqeTjrOX4oY3AgWVGgmp994amb0W+JnHbm67mN8KFpY9nZyS/b1thDlqcb17CjFj1YpxsFxP51
7eR+ffVMCTctejL/GhqWjCb+vx1sglHBQxNyCGV+VSGVXUBxnql/C6af4rQkO2KEfa8LTOW39Gyh
ULLbDvAx1Cs576SL2Q5He7slOFucMxJfISYMONeGxhNZVqP9zZrHPX3DtFwSmJuCNVYW6LQjVzgE
zUvpbUgnc9INzD0HTj0XYyG7L/OmVE8sP0GGfQpWoO7SkWNa9ZwiuEx7bBWbYIr2yBtYbhCaxcTi
UCxXNFw9kV2xUXaq32vUfv6UT7H7qCHvQX78WRY2uegA278dDWJ8IOgP8ECsTRxEw/lJhgZxEi4+
3wr6R7iQ0te/6csWuL0pS4EuvPGr9hRbFeEkCyA6krTrmuL9AYKvGqE7jLfsWgB9+hmhre51e1d9
p9orXX2rlaPTOnGeX/ljpKkVXcv//cYObm4rVSOq6gCD+nRtUWUnL1A9Q/b0f6ku5oQUuQewcjXn
lrR+ch5UCYddj7Tgrmx62H0wE9gPMvW2nJmudo10fw+U4tHrrHb3BEcrtppG8W7o84JjcSs/NRLp
hwauFP6pZqxTtt/nGwJtlD92aEXJnGgbWLvf1KZ0IYcJAhvfFYmqpWu8R2mCj+VaOgpCqCvfUrTg
QY4px+yQcxgLpmHOKm5fSYZVaLhCxZ91lZ4vg3jSPFxnP6bbpUVY5JD8fqhLjuFezGyeDZC92pLG
OUP5aUazQczPqWbgw19hWxJrEfsdhQo5CJzcttgVCNf2USBqXCJGqDgjfxSMgrwmw+1DhMq8Sk7K
nplH+/WDGftB93pIXSoQ0kuYl3X6xH0FGY6lKMGN0f65A8PFeLkQZULmERO84Q+WkYYyDI/wnCIu
JTymPwoRC+SqsSusVZW0DK0h7YIccH7EU+ScO9f7Aiv/JdmnERBMBeMC5QzqoOrLuKB7iAK9pd/D
hbTepX83/pC1jl1B+oK6ZmSqHd3t0J9yROqqMMLmiovh3CtIUA4oTQZIwXGe7HG3ZKiqGpXmYxlO
gyt//cBo9BvFRXpJF9L/LyWX1+SjW7oc1F+dwMQzRX6RNZS9Pq+tqwcuH7P/48d9yGfqbtlS/L/g
YNMLOvzme+2G/hmKrYCeaPSIm5fyDni4/j8KG9DqA5TsN0acAKisZmsaWbwHk0uyqGSiYqTgtntA
JxeZ06YYkTIKdIMidwx586YRWEcMiOc1tOXwGdvZUgVtUEWxAZv8IdC+r707uE9Q1GZShwtbMaPY
SR2W0cgC67c30fmOAiMge7el8jHSleMebMkDNLoSlNe9poc+nXFWImQIkfudb6fKF71uJUfd1jLI
5+1Chy/5MS4eKb4NPzMFb7Mtz9QMV1rnSqpEC63R3PnuYxT+oxZztfValIYJsScF4iCvzIgT5RFt
Q6P1yt8NtfqhR+7duMsISe9Fq1L83+ors3/ZB7vk32YS9nUhCcAIYZsF0UZoqIC6UXqxMpt8v8gX
haASEmIoI/gEPyFNdOZfxIsFTZ8j4zOQx7uKU7c8X/SxZNzE6Zftz1+KOL8IgfndQ0t/E869kdy3
kE7Pw5uaIkPjAYVjGiuKW1u9vS1N6P3+vTqrS2q3nuXbcYSGM3aT0On+goYQ0T53B8Xw3FWjtcJh
t4AFqUWzrexp46oKfwgLkseWfjDEyFtIEZbavCh3UtLQ4zfKAcZ2NYGmH587IyD2wBd+pAUeiyDY
AjoWcN2KNpP+Ea+pghsp94yOV8PA80XoqS/B8KvYu+bqEZ3vaQLcc9eQFn9VW8EXpKfYfHtIg281
wyF71+6wssR13PAKeebrmng/HHjOblpUKxns9a2b9MeH0c2O2GME1Im5ocg64kc7gN5dHrgAWa+l
UI9LTNxo4zArjIrejuqU0MnXv4xUJ+t+1bq4TkRvCku13oWl7yCBWylFaOOOR2kdiVgXAInrsODT
cOfI86XPmCm/5qg5VnrIsnsI11jcA8qp89ho7k4uXl+Ncl/ta3hDz3CjG3sP4vymoOXEu8WSon4j
y2o/DDYqiPZkUisq4v7h8r9we2pBeOzyWcB00huO+X7gT8+516XIggPPmzEeqY5iwhjzWXgMtJLl
5MRtGLZLcbEbstoZ/kcBiWrqnkG8H9p9SqSldM9KmN4wnGm93tLZXByfK9C1AUAGTSsEuR1Y1sV6
MkAiMALnT8WgRp3DR6JbeUQxZTNW0TFo/dAK7JC9jD/dz5cwx12d/NqBLxtFTOYBmTUGLTVQkjgI
YExt/Vock23TKaDuc2d9pqYHLwh8HJ7efVJeCTqYnSLhT3P0qTIRjlQ0yWm6ayg24hxtRdhahZhJ
SlyyNvY1D9Wosi/f2UOLj9MgZbaqQlHNEwgW+yglBCIdhOtrZTX8jiGkVWEKB8Bg/rN8OjZUwq95
LKQZAjPTqZfKcv1NcVAleerpzizjDasYcNMyRu+KVKeML5Ws+AT3Qcwt29dDu2wLjENtQsMkOOa0
3SHVAihCXHSPLZsXb4n8k80ZMpxpKOl4ORotOEYfYytPhTvnESbn9MZeFBoLvP2yXJRIpSm7D/bn
QpkItRgLROu40c4n0zttHZPVgjcdCeje+GdIWwZxtYkW5jfibRmaMO/Xdu7lW85Qbn/5rFXU49eB
UR2nUtkk4zIwI5W+ki3GsDyckrxKbIwHdLeJS94SQY3LjVHoIRSy0dFekhH0Hxs4g2VXYe0yrG7f
vXLHsORGePMqxToWffonAcMk2QvYxPJar8nS1f3X5SYUOxcQISJcY/mb4yh5mRdDOrOvJp+e9D3w
zhDiwTG96tHf2X+txM0uDXtIqYiwCVb43hjr19yECQb/apGwfTZinHSiTQWP0q2TAgSlxP4rEk7n
yAOrxMmXREbDXDm0OThqe6xAPiSXqY9hdT3nm+RoGV+GqEZbjcK8fGZWZdXDJoKwFEP3a0pEHM8N
Ob/ZfTxoC/8i89zM54Bk+EqAovVOdZjIkazdLXi/ysDKzARaeKKbo+nRx8xR0IHY/bum1NKu7/Pq
GXFTytQSVLLf09D/lhPG0vTLkw8DcOlIQAstMCIe03QW/2nWNzDNJc50khp6AJk+UYtiZ9IBKHwq
Yha7Gdr24uvmeTH7nDifA8HwZ8ruZQGh9xlzSsISPkPaYpMVhuvPU2+3qipdJVlAM+cOk1asxdmi
6szj1/XQtCctIMUqqIF7+Xw6XUJLrm9PK350AhrELYizBopQoz/aQhwpfWTx5vT0fjJWOapenN2Z
6KdSmj/DGBG4fx3VOyYuKH6DPPW28KK5z/8y0lNK64xzGasksEJb6OGVSLIqGdl/+n9Wfjf+gfJG
yIq8zkfNDJ/zUlKdxN9pkDTzQFDm39Y3MGlafCTsUjRV/S2p3Xj7oeFsWuqA12tW61eLChavj1pJ
kl/3blnk8yph7zY+d6/uOmfjXfbIxAfuw0QgZXiDevYocbWTB+GHVI/02SgF3+XEKW3yhw5Hqq8V
0UoUntP9IGj3ylbaHIwo145IYy+SgLbbKo5IXObaMnXy9KdU2UdwQpEPb314TJwo8cGd5eyqg5iv
KaAISWhD2x5AR/dQgjbtDwBm8Dq7eB48p3jiENHyZ6ziDfsW6jmlNlgU0rX4Ws/ppIGdLIFmwWRw
7NMoyWV8YTpgqp3k5b4H5/P7ths0zwGTJRw1F6/k1E3vlDdM+dqGkK8V2pRLTsl7n20ji7okOUwk
rHqi0rXtR/rD/7SSBOIAWYpYqWgPbZitjH0XkmjF1mM2XNawZZpVws47Uv8C0Mwpy+ZytTWOEJYc
045Vnanid2ed1RFGORS/2JX1lXXzE8gjaY/J+gMDyDDFXc5kmM8u7qyjFO7rrRnAaBXgA0QsxMNJ
dMhbxnaNdRTexrZLAzzM1gBDUjyYoAGS9ob5pYkivO5oOWUI/0CdVmrDmRF15Qvv+0roTmYiyxZR
NYUxvmdTE2Sy5ysLMDsgKyr3kwPUYi3i6Uf6dUgKLp2Gs7j2FeMVsFQ2b0RTjmEaINRW5Y2v7GuP
tetzXaRH8gdpH6Ic6cKEKoOPOvx18Ld2Z3hhXqhStRFPK8RKBAJubSsrjFP1Bca5BDD5DrlnPY3x
rqBumG1+D9DWFOYZu031UNGKIPFkzVvF/OWWBANg7welUSdkz2sNDaxmyhX+A8u20SRHRp6qxDxa
lCe6RgcM/UsE2lw0Dkj4LYe4xwGRsTirH9dZSp4yGaD0icaDwhN/NWhb0fptO2mnckxT7r7rSzWT
MW8FT2+p4SsYiDToOy0ZhozuggAA1brjdlfS5ytNuA3FpvP7gZUVSwc9OIOuuM8/2pcHEtNWtBhg
q9Lzu2/29bv0J4l1+MoYYs3xtecAzl+ZIHfzCgmUBwCKDhHkLYe4HPNUAnzFz+F7OAp3cS8CJ2jx
pyi5KY8IeZwx9u+7JcpBrMzRH8oWp9affIiXsuZOFCNMiu9RhCCAfArpDCKM3l69I7MFXI+sEgjw
x5t1uBIY7N5o8XVo1ligI4IOPlmeNyHLyTIU9OfGPHhKzLALZzzrviIUjovkTlzklRxtcZrGQ8di
Tnegs32NM7Y8uGHO1X5+CnZ3EheDLz2LCG4i/lyBOB3tRuzlE0iizyzeli2+T81CRl5ezcx+zxib
H9QX5FHc27DQXXn8oTXG/3n6LdRELFO3Xwfui+g+1zrm805eMDKHzBcQDHz5S+ABc8rPovcGGiln
JYmUBMTuR52pV8w2121pBRMiP11Y8tywo29H/jIYHSTy3m/rsL5Vdt15kuXc0cDB55ucV7MY8sLU
irQCciBm7aobbv1B+J7ZJDbB5sdC+xSQGuKlNzCdd/RgAqRNm+VHrUL3RocclPalGZBnWI1Hclzm
jfoa/D7Q1QlotK7r6XDsncRIRHIoI6sJOhPf2HGxM98SIRRdZ/NA2Nv+s3oBtV48NwW3SPHP2snq
KIEOID2Wa/KT4mTv7Qc9GzkQIV8+O/shuAGOpZE3KYOmZkdMmZ18gE5YwEr4jYOhG+CCK8qNLjoy
ZLZyz8P0CQky3DoQ1a7bxFAX8mVzMJeinRMitEAVErbhOvU4R1IHox2YZmAEBhMy4u6yp5Jpd3G9
+pNQ4p2VZT3nboYKtSvR7nxv/+X11zjXOIIlxhSWiQwwes7zq9h9Z9s+x/mb0VcGxhNVl+u3Z7yJ
KabffN4fuPmn3sgbj6sj/t+2dWeiNcPl0gXCd8k3J2JMoDOzCYzOCCIzPCo3QEFuymDQeuYO+Z1r
ASywXFMXpLcmZl/ilCebmWTx2T82QxHFcCx6XbZ17JcCQ0txl1Kf+bEOgQC1tMqoJwbgmbgb5g5+
INAj0+edxN/jJ0lLIWlpG+hJAABL4Mfi0uYdk65i1QhbEKbitH6Yep/P0JbW8Y7b7HBi32jED6yT
htM8gpHK452XYGHWghhIe3pgHKGcjav+4ByOT44aMKDQQf+VBlenDNf+g6qO0nkVr/AnCfj8oz7y
iCJrhyQ1g7/O5fGPbhJTyGQhtXWzXUSJcgGpd4F+0hkVP7SqOxWOR/loFUDLyPW519I6iwNEu1Mf
Lv1r5Yx7zddyXJtgykv1LZ/Ox5SVVrW9BykXKKdKEosQKyRO4rpKHyjlJdZAmURP78P5PW6G9cuC
0AZfisWHYiKnlGNpbyyMz8dEecTx3DQ6NIU9BfQBZbySznotKAWQYGyw9aSQM1pvYpE1jcHHTaN1
24JkDY1iDogXXTqYo/KPrfy1LGYVs22x7NxytPv0P2Ab4dbgVvlkvDkld2jVsjIIQJWqtVNVi4En
IBa8Nzi0+oJHH+0HLtv+q9HzyBd6+9XDvMsx+xJTedDUzd+66LpqnZuzm8DsZVJ+WkZrS1qv83eu
0rQltvZ45LR63So14sohkxEdOBPaP46rJdA3hgEiIRHx3VNUd96jQs5mC7pHxUntrn8t0FPjdbh3
ZYZd4lYwK0hwkJrtOw9r1YZUy5NZv/X1ggf0QTYVyoGzC3HH/TFf7NHn6eAy5OhTHthvARSsx+Hv
JktTKv5ySxy5kScHsscYuW5wF7NQeodbmzJkIUCuB3upwhxg6Bnq9Hui8zLG2wDyq6TfSfmi+3uH
NuhebYcb8fGdIxdYwL+41KlyIRBD7nBSRGTkSYT9zwVWtr+xsxuylLYpCGnoHsxqgsM+irRzoJ+/
J/phOmScX3lNf5E9Jro+6rDFi2ceOVuUsyZ7paQJLmLzxc1jamoWIx4qKF9ZrGfJE7nSWl/Re3w+
zOhgRUJrV/OYgezqhTE/i0wNyHgugxMQA5MfAL3St1tqS7P36/wJheuhzYehNMJdYyAQGQ967F05
3DYVfA9sX33U9pNYIk1GfEBnx7QTuyz9HZIPK7rFu+9YQ6tq0mVTuD6yX4+Sx/nRGDlo0GMbj0Ct
Tmfdk9gILT6UrZu5IWzLBJUgaMqrgJU4FIrpmhYDwcL0OFQaoYtM9WLHAFvhsqlAmS9IDEQORBnC
Rgyi357BLlQKrqtWPnmM5RB9mGe52PC+rkWNLfT/5Btu22I+YizNB9qwBwg1MNJpH93ChAYvOSJR
AnPAJoC3j2imQk3v9Rg5YJ58vYiQ6eQd/WKIHNx5SUErWiSJeb9FsDOr7NPdg8gwubUem/LA17HG
Wa257Xe0jlcSjeRT1B7LIDCbtnXUP8khVxwm71HnMeD/nfs0pW4KI/Q7wETZI2D8hOw4kVUt9LSJ
YVQXhmsWCZ7+Z2DWK0TL/AXkrPvkg9c/sg40jg+tVy70uJnFU3hgn79ESmtR43ejOxv/vt0AR10e
uY34UpgTNQqSZjy4g0ewjrYwkQO57QQ0LPfv2Ajz5P7x7zgHcUTL8k7ntNzQ8BQE9X4//QukD1yQ
okOHSl7EpIWlu12z1uOT0V9clpUvKC5qjSm0NPvdzTZ9lf5/A5d2EPAgD1r4l1+dk/SY9kOiXFCD
oRUQ5ul+sHrAygkzyg9W0dotSZc7w8ZUs4ZpkYp4KQF7B1mNGN9OSz2mPehfDIU4ncKcQ7g+7DSN
y4kP+GxgIVuWVQAKUtKTCC3QdxMehP9yl+m6OKO9649sNVyc3p2pK8Rnhi9OV4Qotp7Rbx+SXBEq
QIOND9WapkDo0Rh0E6cNq+GZE0GbdoMB3xvhALRmYnlXGXlta58Z03BjtVkp/QmPss8Kls+f6eaM
53N5c8YcJLTNi/sWj45+polIdL/DpATF/26bB2ppMzxEiJ3x4B5nmpsmkwKBvn2eJ2FzkZ293xIn
sQcuFPjWKi9ePJ6uAc7it8FrmoDNbeTAK7VQcncT4+2R4996hsf6MouC8QJMxMC/d9tLP3O4IGr7
Qrb4v7OZ4Rvrjrxj2ddYhU+JDTwexL/CKUtwrxT0BqhPKTQqxiP6zvf+2WZbt79heuL1sjocIWAL
RdQUqIt02E531KJjamv2KloG6MdYnM6VoNMOalUN9E7qCxcy2bkRbiUsVUuFrnTQ9x/fyNQNYHia
zXZuDGQz94CzwvSVXK9wjZyJwZ2WN9jT1lTeKND31QIvNUpJ8Ft3f0H+nOg8fNxqyfet75PE8zKt
FabHF0cayRb+CF1e1TqO0IZwzZj72sKmdfPsLKxtCRb1tuOBDCRI9Su19ENS68iNkRr6B/oFEvxG
mxqeFu1JnBHXwrFVcilzj5fKLjq4nYogGHyVMVDXq8HxZABy38ZF2X2ZeA3xMGHuQXtbADAIOARB
DilGXVzJ2oXHUDqlb8Ob8RsDIS2Vq59VWABeZeF/eC90QHhcoB7oG1OxWgjNuDI2nbxV3qMF6RbZ
WLuEzKgAfhBMO6NA5WBxBnvVzeArsfzuvlVi3yDz2jOnhvQyKXRm+waoGty7hGhXKI9zXA18YHx2
UtomFJ5J3xDxyJwqIqi9tRvA+AlVAA3cZ31/ry2FidPfUIFrxZm4QMP4oXI/zUWrEkm+yEIW83d0
OHf04IjsXiHhSws558i0OT84F2G8UCGqBtmkw+Zm1yc2qVDQ6M/+8vKEmeGGNiJEI9I6nbNb945f
v2BW3BuJ0Ekw871cBXp8ybrmSohFEAf5mMXYIy5opx+eh2ojOrPEo4r3x3KtvnH+nqoRK5kM7Nts
oTwE8iaLgxOjIq2QiM3pXlx5LD3yufH9ToZKqI9WttBwbu8zC7UkSNtvZuEy2P+tK4ihHQaAAwgL
2mLo5yVSn/4YQVaWoTysP5Wo850YIdO4ZPd5j5Cp9ETRHQal34PaIp2IB6X+YGxa90D0UIe9ClWG
F4QgmuvW/856AV5X7BtgFL0IcoOWt60JSInPXVCYmJL1NXkXKQModcPmwJ/tAqNswr0zw4/svuWe
WT8JPkquBoR85oAIFyrRP+jzS7ch2iDh+JGQwqBGo3v0GMM/HQ1MuW9YX3JEPVVCz5NR3+lGrXgj
dvMMBA5WVYZAAFYKwtq2RZd5uZ2Zapu/WKdtx5oHFdJk9MQFMy8EWz0CNSKHbRWq/qYw0/h8FsOn
9r4ea1L0A3LWnTKfOIs7cK5TaN4i8w6lKMwJiMeWXQqBVG//fiv1zntq19N0/J3AxfAywZka7cgL
jFqmMPb1uUxslpA/Wownm8VkqzppBNUlLyY+5LHByh0+8SzFOV7OEsRzx9GDkijt2foMKRL9z4Q+
gQVLXbBVRz/UBL33v8RPmDew/O8ogd4RAJ7sn3HTL0l8QwYF4Emsrx0Q+GOyUCC4udatuFAvBgOg
M5ajANuyyyP3S0u/2/ax14hEUCzr176wOho/wRr8fu82VEK6v85fuyv7EebDPDQzYhjlhnRAlVPF
HchjnQ/3nIqIVss8oZbQRTgIS1G/N9+dY2fae4JFGJOrDIa2M0i18r9YL9QtO524TkKcruXSXNFN
CFu7hCz26fnP4rJGuPqMysq3MZX5FfhpyVMcODCr4vBVTbUBpdOh1XE7hfcUDVf+LlroQFNNb1vk
xPcoGp2Koo1ZB6NAQ1rpgXvLvKBhfJFxv3/YL1XHOIK1/vErg1LkD7pIhQVnljFpXDeWRbWjCtDL
A+cAmTAwt0CCPBWM4AE6qQkpm7v/UV6Ua6DnGi+XrCTorIzlqx2RGgHurrRmESXs/IFHsCaDdE1W
udoH6btriX7ywx2WMzKMKNlaukhQFsf6HuzSjrdLN+bI1CJTHEZDL9FOCEUpbjB8vQwKYnjMPeYp
cPWKEkH+qyttpMKFaOiCXRko/VRdv2xYyuiGuo3FrpNygw7qxzIHpXYMAOBdf5o2dky3YIP1ZRK/
q2uGIugBzg71nR0PL2lhgVqTJeICD7r3DH9wsiLLO6URvV0ktUPm1ufbRvatZl82CRPL62UIZkjg
IdSt7b2RP8UGhqbhiHz1uYLLaaYDMtRiSJdFjHOo9qcQmzPmD4lhMgrrWqgxemx+bxWdZe088UE2
ng1hmM1/yDG6HHcnRWBsop4BViObRMlOAHLfYEOn/fdnbj23DqyV4gzWV+TUUp6M9KpPw2j+eo36
nXE1TD1x3rvsSxn6LWNlV4dNot2XnIyRwD1NsuXy7g15SGxpYvswKmRN/GE2DFiZukcEVlgEtSCI
q3eDUBjTvJ449tM2VIC1YAI5+zglwED7rBddg4/2EdOeW699iowmYSItksmIHy7hiVdjylGa5qK6
A9vy4RWZRxHatq9NCDjhiWkJZERvzK9mLPoGIQ5TqLE+3TOR5C9i6BiAacMBJ60iWbYvxmeflIv/
9638UeRrgFljTWefbhKfUFEOwbm86ZCG5t/5z/V/mT951w/IHNvFnAuhMs81OxyGMpevFMpvIXoG
UpaoQRc7kPAcuTFb1r1cECXKj+vAhB+nPJnAmbhirOMMBAKLA4Urn4w9syyeHbWNz0ZWWoXe/0ca
O4BIQRlwY+krH/ET8RhUfQLphA53qvGxaNwGPHfPs3xJZ1ibzYaAFO5ZgeRlbVaD/uKMA/YiGgcu
3lshoM5Irzu8kc2+BuwliJu/mpU84XWS6r1xX1jQOrWo3CIXoBWU6MoMR6axobNQyuHXCpI2SF9S
KIl8vvs+o79tKKhY0WZj/1cf+fyHLRo17I6/wmUyYCbC5wR+WHuQoVS4VRjCqOgWDibIsJhV3Wm7
wqoDaON+nKwVN8OK3yvTo7EiSliVyxJQUFfSWyXyF3ywyNbjwmTyKs516EC9nDQoRoKzWzgKut+q
Hvymi0EzNzLKHM8GYQpn+pENwvsHZy3Wr10eKLUIFS/JSwk7iU+OmwVZYZ4VgwEDCeQAzUkvp0cE
JSdQFBHHdyUIZW/HCx4PHzJBeg/IWn7aehebfoZaOZIuVNuILph7p3/OFMHvw+symS57PYW2MT2A
DDHj3ESrcGHuBdk7/pcQziT5Xe48Kez02kUrp6s3KhBKRU2x0yOnPRfK0LW7LGea5MfkdWRTkovz
LrHc7E+iyQhWPepnxidUAehxPfXTq8SqItmDxt5C2w7gSxGyhThSJNQKrL9Qz328lRN6q0I5bVm3
lruwnt2OWNMOaPaikMZvIeOctENo0Lxk9inMEM54X0Sf6Vbkv+reJSXad9oldj3Q+Fo1SOrwypWY
URtYW+J2+Gy4HrB6iMY08aM48XWoaA1rOZgOxswbssa82U2/ZRXkcsPha697SPgv8ZDJ6bZ1W2Xr
EfAx+e1n9rouvLHIFl0p1PJavTAqwNBSLT6qjR3uYj5s2riIA7NMwStq51PfA5tJPss7F/fynD6Q
MprS3wGYExCKWZf7g6ILsRCwpJXmjV4zGf9Kr0EN+21ViS7ncYJr4FSDIPiU/05DMGrOzTOUAr7s
gE3W65xKg3oPvfsKNrwxc7bPTpwh3MIlfwWot4CItLtzrJ1+XhOAkLN1ASjixb8zQ+RTktsOKSOX
Bggc03O+xox5ipSZ+HJIco9GNlpUl3Pdq1Y3/N8tiC5hAEgCViVavez1tM7TCFZEJFA2SDuSUhe7
79MVVmrnpm0vlmgphVkULJkytD+lIvIE5wXceszD4HX6WtX+vgUdv3OZm0h62l12HbfdH8NLFv0C
e5YVUpoZOWVYSwArbbohMB7TrGo3NwBXjK0T3v44yWdRjgvzV1ka8jNxJS4cEVg+qM9B9KBwW4U6
zctz6PTLKm8SkO9MQVRLL4Z00myXjtlj7aJB2TRCOdnn0ZUjUItnakcnh4AWXGQFwL6ZVtnc38zC
u3bVlC10dmEoUdQ4IJdb7RDiXtxlsDJFc/O2y+icDroUMLfxqTQFz2qhbAGzYzrR/W5TWXHYI2Dg
QmBLL+n+Cj0reVQ8rpcLvBZQLyPU/4BkIbEq0zl48W0K6rPgijBWz390RyW5f0gfOrnpjn/UfcMz
KKJaR/Hog1FNyYcDeGXDpNjM9g8RVaQBpUG0zWEi5gfrhQDp0+OglM5mTU1Vi0pLhWrTtodgPskH
cj4RQcM/0GZ/uBUXaWp9xjzbdXcxoNVuWkbZXlNKUCijouGSMFcHH9ufAS5sYU0+eSIavnPpRBbG
5E5g10STvWim5fZRExUXrfL6Mly1UjYS0E9NTQjki+DnVhmfkPYtVebzbHqYWbvhoOyJ3D3f3MhM
7ruPo2+bTOXy2pgvSyDxwNXtjBWD9+nIX/GVahdRLOVmR2sfRjy99o8i8e0F4QdPLUUeM7Ck6XfN
zKPTyX5telGOGPVJAl8s9qRKDtgPn7WxzY1lKhHQNoPGV7LKgSmsDXUCHyOKe/8TvjV5LO2aRupF
vlwvLUvsjO87iL+xXrBuvcR5R3UdSNBlwtwAo++gVtOne3J/2xlo5aksD2snGUYzT56PRzoAGL2z
SxVsBYaOwjif5Bsu5mDRiHFXAf4xbID0mr+YRB0N5H7uZHbfDBu+wdqZfbDgFbQGqLIDR8172Za1
075Vzqdy7jRLdfxNob0Kyjxbu8mbZ+rO92JmVjvCBc60g6DbCIyYuspltYYYzIxLxCs3HUjRAK+d
Z/lEehIGbamaw/3Zg6HK7/uylAEUfcMu/HaG6jkjNtaJHr92hha6jR6BqUurG2ULuM6ozmenQVd3
pe+ZQiMPtV45gVNRI5gNbby3VivNO64y8Nj1j+QLV6YtxNlHYBf8oTQ2EYG+CU+A/V8SbKYFmiCA
0WS2ikRBO94fsjFvXrWGS6HNsbqJTuEn8zp3CLooEAbad9+AaMStJ7HUvGW2skWbOL3B88dlEcKy
v1PnxfCt6nMyltYSQsKkHtV5642CdaVHK1BLdDOXjHYeCYm7e/6wUG9VxuNoVZrkUKH2Rz6sMzbg
Jkk3mR6Jvk6h4Vb9Rg0Wtc3N9msiMudBNoyJR+erPvNpmPysMqLIhrnHInEzu7QXzlZ2XdN7P/Rc
3sOrnU0nVDOGRkjnAgJgQUl0ri5p8cd6bVbXSkv18eZaxOLChipOyn0ST8GJA5AakOkEdVaIQBLl
QTH/sXwT6qXCohd2s3bj87Wuu2i+NwCz027dvE/hTMnF9nGMbgKvKPHmw10h94VJUfbv5OGxkSkR
HrQSLqzIKQLMWyo3vW1SEQpEJdAl1CWFCyg8eKeh8cfAAn7ingqTv48kS4lONd+oxiUQfKisGZqc
aZARD3xRbAjSdxiJEKrrW7MdSzfCxgPJXO5dL1cKv8KVLJLsDU7eddEnpx/SW0cqWs5Vd1+x0D+t
XmhZQLcdF3FlszKpeoPwatGj5V4qMKsFd8iHMldMUxexZwgjVjhDMNTBjjFR14bT0ZdDRZ1rm1sz
64O5HfZ6TLnzkGy2yL57z7IgdC2mB2hJCoQYFlV/jyu107ln/gxAsR/JIlIcVJrTWAktcXg2L2QJ
sIUz2W3zS5P3X4Xj4Mr81cILM4oHbJUkOvPHtjn/gMVBvFHzYlR/hG6K4eAEccJ5hJeSqRUhR9vX
gh6BetJz0FlwKkNc+K5JpXezTJiYwUTqWq9Q2yDoXXtHHGeiFXAYCynk/A9M/E53ssbgE/iT747G
cBH+WmBnwocTQ69VA6ZkZQ/QbaulAAGj/Dsblujg5E628f/c7zBK+s2xRsuJDMHUSeeHdgmOwbVu
nQdOnHfhSfhzLughlsY+7NPpoAM6OCsnR3/hZIpc3G54BGASWk9Um8DIs3B7gd+4dPaTH0b0Nh9l
034GTSb4YEJjSYYpE8lrjqo8LhHE7zqDrGhWlr8GNftl0UeCaursF4/OysRc1807dV+bdqvOIFjI
8RYVa3po8gLMAB/1ccH5STS5il9TYk3hFjHyKT5yUQHys82S3+ykFMo0+2NeHt1Xnjs4ictS2NZJ
VuHyRpYmSdHSE4ZdNemhOgeJckzCJcxo1Fd7L/vy+HDbYZ02oRlmNwxskrrmCaqZPmfq/Pn297H1
qXXc5kWUgjHO1YzqIBHgfde5NpbgJ2i1hAgRxgAMxbOK97NdHgxjsIX7G+BtjOV8MSchJsDIfW+s
CylsflKVUn4UuadzuhF13m1/wOU8D8qiuE4JScfxq8gxg0WXUKbKSeiW74bsP7yYQEBsyediFpKi
1hgM3toLIJB1NZI2AvdYY34F57gT1CCIsdLELqHxztRRF4YmMsb6UpaQxemYeWBplggJ1Y5/zdTC
IJ0blza/4KBi9aL4EAP/lyhCqthNdj0v5z7fhvo/iAQjHp76WD/t5XAvjE5si7M4zRIx5gaU6Z9R
xUzkCuMestH+gcqW/cNaAd0swmh8cWfqgtM484oupV2LIywhE2yq37QlLA3ZjBLGYrRkM7WgeYLx
umI11j5EqJAwii8S/i2gOnbMlBaROLAgA7+JKm1Wjzaq7oIO+olwaKrSv27D4kbfdnnnnkEag7/R
mjHYo5txfb4ORbJ8xMJbX0pHnZ5BS+RnCJTDTeRFQGFSYif7M8rK0UCaHF4RdrsFU1AlkwHQQ878
7iT2Vuh9kcSPR6NPlAPK1JlOeJ8enZ+K/ug6Dvt3o/QdHeXWM3sXUvX0pYbNhpNIIo/SluX8m0uT
7VFqCoTV/FAJVpP0iqdNEsV7ceFm6FQ7p1xs7TN6PH82gpI8uaEoW1XCnH1HXxI5Ucq17TR3QXgD
kzCEKS7ncYdmbXkfklydljAiFNPyCQMxNEu9mvzfYU5UgVJ/rSN2I1IInmaz4HtFhpdxlfzGQ1Dq
aK4pc69dn0qdmAGS8++/ysBJu0FuphcxR+3YeQ7CJTwXmrUcSbwUeu0m8TxD7Wzx5D8NBSZ4GZH1
Y/iF6YXoV6J29eN/W2babqr9HRTfjLVw5CKxBgYrQxjm4DGFWQTFd2d7HtAK2sk9+KeGtF1xCnhh
qaqee/ctGtDqAo16g/0fbl0fdivTQ6L+D6Sf74CfGHFP4IZ8du51jYtIYNm7P8UIoUeV6OnFQvoq
R7QjdaxC7lEf/x5nSeYWCopfDkhTR0piSaEQyKKe4X3HEK+ohofRLEiwxPZAyuKGdGiPqAybqfjy
R32LIvrfa1mnCJ39Rvg/FiGaGT2fg25PI48j5/Mv3wy2uJGkUZJT3gdNKJd9/mT/xHcVup1M2/Gj
oQ/NPmuuvyRvVT76BnImT2faDd/LjzrMQ37/6+vv3OTTBv6tNsX7R6O4f3oVaZ7FrjCl6XBW/0MW
MK/1hJDh1xSPooDboEp8mLbIZQeYQDU5igjxCXDFFYEfkVo9cRT3cE5EW4xGQTmO3mzwnY1cj1Cm
jAH01to/0EwYslXjHiC0oSvSTcEXgKVu5M00AxEGixfpk5w8K9cr7wnJ0Zkj5eoBHK4HS3s+jKDK
HyCXVYm7GxuNOWjtVPAGXeVmxinQfHTgB/TGB0mKcFqK9PGt19Wpp0c/+hPIr0ucJfVknmi2l7WO
1FYT+EE998mGy1uiBuyB+KM0PcTJVZGDMtyoMmF6gblq2i/+y7EgFy8X8YDCpwj3tFczDzmbfBgz
aXP/9j0yOOwkntE3aBspI5UvCEXGtcPIC9pJND09hCsDjQe2DeXroEp0orsZ7DzRS5O+kgTU2eO4
Qq9j72EiWK6DCmWIp+txREm3Y+R++IXzub/5FG/FCmzJB126Oobu4c8IVLtTUQpXGkOuBJh653Kz
tIt2prNTAjByqffeI8sFyGAQPBaa2+QBqffG8aYFrJ/h/yEL/4YZOOqOuTki9g54kcM7r7xRcbRN
oiTXPvDpjaMhqY37rR/Mxv6Or5et9C304ZTe8ixp1li2AuSu3Vs8hQtGt8AJixfZYEqJUA+ojKIm
J36OhDrcmydophhjaL35TBr5KR1z3Zip/pPuKZhozEBEafVxARKJHsEj2GVZ+7+kTYstTtmbE/Ol
jG+x15B3jM50Xdi5GZ3EyLAim1g4rJJpPM5xPfsRs2++/f51wO2WFLI7kRxHbHXtFA62TTqm2vmA
ikqgfDzwGYOrpX5ET5zVRzqnMUj823sWgU3uxbvyUo/YTDrHO3XwElC/K6F9Ri0kFn/UnMonXATH
UsRrjKuXA1gsQhX5BXv2CaT9sWbDV1wM4OJvBpPobh6GQKVSNl66KRAJzQoxwvXeEUBMU89wqzz5
etIIHv4hkETXe0JZYZsYy7aETuf/eLmtqTDOCWOsYa9PpHVEto4MD34XwACqU0r1oKNZdkiJWUTw
7zJvvNQ8jR+rcT6rhrG8jfJynrNJne23xLpg6x6m9gP0cwwHhfXkbj/b4n0aXEPny45DrFTin+Ql
V6xIbpJRwYJldPKT5/YI/06GMGxzTml9clRinC4CfICakhKbmAH1vw9EXSvWQic1DIZKnukRPlOC
7ZA/fd3oQPYTmrZ/+3hg4tzsrNt7aaOVo7Ik1LKWAqv9jlVZVr3rwWhq224KGHPKecFKs+Rj+ZV+
2u/68qFSZb+rD90yLC0F7lhP8GlNOqG3XrcfvKyoVCPAY6iEqzd3odZMM1z3SZkhCL0/8fDPb0Jv
KzR9UojKW2eo50EwZCBLFcwDD83NmV0PJLe/jA2KhyUhm/hq37LXCO3HEM1ckJT0OcF+hFuXWSxY
60OLpKEYyqe5pPvRflsDCdilMxczzF4EDvHYyOn1lmqVACXRNVnxcETC0JNycBqoNqdc0fO1F4AR
2zL259PmZQ5ulhDkUxRM3EbBNKvv5BINcXjMnBEmNcfEWnHxWrK7i5Nmw18epIrJMaTHpJodAe6B
C5CU33QluE/7yd4CMUdWPu5/JtOvJOdwcXiu58ylXKaA+86HLgOb+XRNA9W4jqOc/3Fb9SQ6OC91
MauzW/mT29gOrgK22iwue4nWOFuS33X7vVbZo7NuCQqL6T1bhhpLvOBRxDYKrEhxa0lM/szjaCUe
Hd0XSOJrCu9cVVTyD71zccITgBSWEq05X1ytzIbPuG5HGd287I1b2T/uDLQP6ctGnIAcuN9q592l
ciyKZ6PO8gHNIvt+ddt6pLGRAvkXt9x9TO75p5BFkMX20wnakk33IbInRPrAYF8vvIF6I1ugf7T+
uaYxoZe4sPNudSIQk0o8LKFkITkA8n7b4wIESPgLAmBh0aT7JJYMysZ1UE3nsSqdvCWG7d2F63oe
4j28JgOnQuZ0j7Pks5p3ztDO7CtZtQZQ7wPszjyVtqVEivpA56Cf1GdWnWcoA73l4npKkTLCZCpY
x83bNuQIqPRWwFaDBOXLWJ6J13SKMxG44CqOngJuddcdyL2DSYqG5sKtUUxvLS++uxBBz2MKl19H
dUApcFTprex723p/GJJBEoaS1tkT8KaMlGX5nm3BqZf1D3iLMRs6/V7v+0yWINUJj62xZglAFipQ
sasERdjmmm2TH/nwNjK8F0KyTxXUMaR3hgEmcU8gd2LeWsr2+O2Eh8cBAEW9NRMinDu5Uth6YEP5
oAEYX06L1MOKcr1G3d40b3W1CWi0nPWnZkFpbI6cwCMYcD42AwLVX5VXB7woKHhu3QSLXAaT6WXS
R4rmkRy1fjvW7v3t+2clPioTrpClkdsPz7PjoQqrCxuY8iw5MF5WAnu8iV2fDfiiqyXxUTlU6JDB
qpVYjG9CD8EJmZY0m+IIXU5IY/gVNJJkzu0O0FNWJrkKxYrZH3VWVaGY6qpbkmvj0i3gUwI4lVtC
cH23vNz5JcB/DKsX0JM96b9igkAwRJwT/SazwEdyqZwU1aP4hFDhsGHL4N7zs2EZVw8Hbsw3P3TG
woQMOaRZYHzSi/2pIJnSKDIoM2GWbue6IgAxE+mHVlQ1pPPkJGQDJYZp/ifTchjfZbXZ/m8YUXEo
MkeFhISRyRFYbF9qcmqu6gq1huYLIEmt1o7kh30qq1AjS95upqiRU17E/ctTLsJ4KlfC2VLgYYFg
L/rS0EvK40X1NUhaw8Rn/A/giRlqfbtnxoQb1DNIuAL8PXPbh2wedrDQJ8cduJmqgOGGd2DfOpl2
mc3Jx1ndvmX/s0ouC1ZDWi5zimvBRh5ziD5ge0l7KEQUz3Sa3ptJwgsM/11Wy8hcDYDLgJiP1svy
jh9ev02nu2Z9EWSQzdEj2rUag7MLUpmj7HohxEEnPUs88ghjjR9S9zK4gyQ125E4ffWvpywV5GKz
kVvAKPcsITdIiNoj0IXy89NOi+Vqy4v4UMqIk2sTHOyG5PEqPGjQdX8glU2YdUuZvZEpSN2Ivfj4
0Y7Ym8fWbB66xE8lvNyDMf6y/EUXVGVj8ul3CzUIKpigJxrRiopl57PdvH9Bo3shWSmdNzWtIcod
3mj5053RuIOD9IzsgAKMVNGBqwaQqZgBP1gAYoSHKKZAkL/iq1moDIkm1d23/fli1NZUZikPQQdJ
CI/RZ6g8+KdrNsafxoN5pOfaa2d8CDMFPXU5kAf4qLn52j2zWmS2iEIVC5Rx7w1rARPKodFr90NM
eJ7UHgcPdnPwS8NediVSVwDDv+VXtKuv7f+yHTak5+0/Z0jwV+ikFw7TzYCsc5l7nRKR1M3KbmUH
es8aHqkfFHnyoAdaV+OcD64sK3ozJ21/s78rWsubLWw+g9MomTHTcH2y4EcpsxnhZKSyEhKzdXZt
QzKH7aUoCIXPYSanf/oOckYYa/ysP0XWq1lmKz0MUVxYKn3mcbNkfoAMGOcLnvLgapYPnqzf7eFj
OAfdINV1eGVrpLOnwAeuI24kuakFc/oU2P63wlwPd8AQPGGMQpptWkvkccGWHx3euSHwVuJ7H/kl
p6A0Fyw72vYGby9K2+rKmnjSs7LSSqJ0fBM0sOb+Vj9MtbwB5wwYQuxXdviqa3z+2jAeS/CnEQOP
SVs6LrDXgXWKJ5q+rzZWNQl5wRFjcFKc00Y0jjvhi6Qrt/pNO1OoiVKMk9EC/z2uBCQt3D2isy8/
3wi7G5ch1gQD6kI5wytbS8l62Wxd7zibZPccg0z6bowP/QBNz696TfPc5U8iSjbhfAGgRIt8Obwi
tBDJakwDE3R1Zgk7NAbJYe/UEHX424sQiKcfEiB20B8oIGpA58O6KxW1hPTnltoZgVZ9BR4xhukl
GCD3vw9jyjHawRAKBwFksAKx1pQqe0VP+BO7eol+pxk/LpkxzrMqs4VhJ4d9Yscw+6dsgEkOVUKK
wwIrdytohpj8YHCt6n1bayZ7cW2/aWbyyikcONtn+AwG9WR5COUuvfF8iVfBmU/gcMr+Ny+Z38v2
Sz+OgPOHKyvKQoH1eLark0cAMJIs7/b9CJHIRtQe9167EDf6XyiRo2KOOErIksv24gMyGw+gdG5/
cgt/OEv5/gco3Q0q1sDGrnmEfzU8qYg4nxYAmvVLDNqr41WnpPnP4n8QHSIQ+ntfYr3LTOlUBKFY
TY86QAe+LBp5e/Z078qRl+/MGYyxDC78lyLxnE2QrkgnsqqA4JhbtyaJY9LE6A2AnuriIK6AbDBt
C/LSv8DiZhVYT8WWauHekuirWdFbEvuJwPyAcZlumaC/WMJq4whVi7UUhN1XlOBg7QOo3tle019c
l3kdzar3zCnsayhCYYqemhurLuRf5IBXpS/Qcfk96wzgoiYHFXkiTfckUUgArqrApMz8AfWrx1ep
MQM7YDeDVNZHknF7bd3gFKqdfKt7jjNHBTiNCQxXQVz6rmrUuGtnWkEG9XtzJEzGSkTV9EiPx+RO
op7isN2sg7M1Uiwrbl4x7fuk9PxEmuYJv8LSONslVEXrS0o+lWuC+ngYOOLs6Y1BdcK+qm3RZgTt
KIpF8C2Vl9fhsq1sMnmrSWGLCbLrPIk3f6TndjfKUmeCxWkm8GkhQFd0fNyRa9NOZZjOqX0kLER8
cuUXfCRe7ZrEA8mM1Au41/uHN4YgfYVhi5Ne/7cD2nh136x/olW/w0pJvlJilJzHQ/UFE9oDDNq6
F0NYJ4BfDkohGwZ2uNUhkXfuYCEydniPIEjAxWfWle+zApfVwxN7FOzXA560c/MvqqJHaz3ZD0ss
dmMo597v0UIlzNBX4Y7IQkl+RWvWOz4v+6GpAP6g9rcFi83tRnyVWBdetmJEzj+v0pyRiJhC7eoM
dfU8XkwJd4A4AlgjKScc0aOGcP4OJ6urTe0LKshuSJZyMa2zxC8wDtgtOdyEj99cPDw098a14p8C
N6JjYaEgUv3i5RtJhIZ40o4ZDcoQSMtm79XJ+oWTpAIkzCKxQ3GwaGhoCnT3KE3HE985hhhUjHX7
2gRYxyPCTge19hQ1C2DpJpbbJlufmJT4FDyTPippKuzm+LPpFw5uLsf02ex1Mkz4K3RYzUDwSN78
Ml1dxo3JqqBHBWEq7F4IXzfmq2P59jvVZPfRoDDSF7LW9oZ/qpE0WxUpqD3Z7Eo3AyqGjEafSXHY
CVC/w3voL2e8fbXsc7zkJiKGgKdvdgq+5DQnKGa2RlDIXrfCXf0WfY/wWovMRhd1pJ34iPqbGp1I
Wl5ejvtWvvDNZT8mkSMpRUdnpF1aoZZNbhg2lHt8f20uXCWdqHTfn8BAHh6BaEJ94VU+NpO1LYix
ZUx9Q5Q7Hko1cnF7DDQTT1f5tWt5ewE9w8ShsZaqW+cWlXQPIqQaFuZY8Dj46IdMDvKUKPZ19AVk
dq2cRbXGiSFgA0yRWgpfa6Rc1HrOq7supxqGuikOykdFM/vYnpagfoxpcZGeh9nS6lJTISxi8DMW
fIudnMTdjr/fI4Ty1WSSlP4I+iXeTU87179tW/LdX4coVIZUB3w+lAl/Zs05roJVRg7fJ7HmXuM6
8aG9Bq0VRzh2p4K/rlzvATGz3MEgW2gei9zM38zfBsFQRAk9q8mz7E6vHKN8ndVRu/dwas0KbUjX
jhcGroaY4Pz/94lB9056RJxHjoEVF7kqRo9FV2YUmijFnpD4n1+PMho5GOS97IGZ87EMSZk42+92
Fy5U8MI6PNzbh7VR+Rql6KzlIj9hdorW4u8dSLWjP1nh+1bFAL/2QyEv35m5bgiKAatmq3sll1wU
M8VyZ9ybinxnhedIqrT6kMV5L+Mb/wUuFJChF9GQVNuWGiPDJpVD9/CpUyn6tiG833Ja7CN/+PYB
/zDtkRllfvjONzZoRCsbOYuo9jD/w+Rce8bo73bC13jDHOk6s/UyS3zuGBs5kHFHAezzm4UdcmuT
wzbOWKnHYEZOKWowesoqOu7OdnJJ/CnLD1OEDgRvG+TpUzqdwdAqdWDX2/UjxR6412VAZMnuVcDo
YJA80meWsZzTMvQzRC2iveMrXEuz4ohkt0HCSR2vhLfpUEQwTmgyMHj5ucAiHqTSLL3GWh4W3bOg
VpFhBjgT7BBtp+K2tPfe601BmenhHM/CjRyZkX+jOkT6ssTCYOZzW2RzyN6+CnARVfRXnoqzDQzF
xWlEwkDEUPNzyMrQWOfjMID+8VFq25h/96ZzaGIfEKafv3bDIl6bF+hSYixLJLGs+9sWSGVr+HZf
D0BbgX+To4fJRWg3NoaAwrTwJazz7+Sy4Z6twR6XhjRK/RJI1WF6GG+r6sFrNjEQBdPyGTkOy9ft
zeTiR2yT/7mv15meq60+/hy2l0IzR3HF6y/gxFTUobg2/mX17X4OzNdF6+FZbcuo4/IKIEaUhUV6
i4kBof2IgwdAUpBNhyG4bM0PNheQl6JLCYDlDItJFZNck5AR/vHKvBtnxfKLIlK+xT8xBFHbT2da
CjrpPgKywmnAl+j26A6Yy5pq8DVO9tNnSjFQJ/rdfvTaMAiTrBT6cxVojJF8C0Q9iNnkxvrFEJ2t
8e06sytwW/a9ly2KUpIj5ZkGLTffGEMm0/XcAkC3bHf2F7pz078uFzN8NHZVUQnBZyRvx5cYaaPV
9zakgke7S+rbTeKZiZpzRA48Vx3xjP2c9ubixnI61/W81vBah1KoUUD0g2T/dXLKugBY60Dze6hi
6FA83OK/1ADrbqhPF68iXYX192R1Zsc4ljDcluxjWlO1W6viNUNb5mb9bLwOaa1sBxzNT9PXKHgt
6tf5mjUyrFO8kCUjFHTxmQWoTq1YFPdz4uVCPv4qM1qSMq9agDUYr0Iq7gAqVoDjEjDwFtav8o7l
bhPPwAEeOVR4UnDubVLWyY9teNgZldNwHwx74FT6mjBM01qeiACpewr4gD0KxEFuuFpqcJedL7QB
P30M2ZnKKj/xC+F9eS8U7Hm9O9DuLEqxWQjvfislKCtye0D7hwv93O8Uz+HH7E2Rh0O9Bf5R8AWs
NWgiSVDwTIGp0S9KZ+gq6z+R4k2by27lOPDniwNoqCAAEz43hWi041XFeECn30HRgcicarxq+Dr6
x8wln3txb9osZh5DfZdSUEiyBalAFiiJR73Sik8mZfNL41ihaVptKCXjBatOodAy5aflxMa54je1
uP8Gvjn8vhfxcKtFsdpR8qGeTyHxRJUihEvG+KRF7hfp6xnVlw06Kk9YoUjkhYMqFI24EVtj3MRH
z3Ayhsu1Fq2/vCukDM9BUmT0nBtkMGT3cs5pxEbGskavJfjUZipE8cCc26oBfXZomGcxu/yJxWKC
frAVBPKMhzdDZhjOSFBFWa4If/ws7STyDoO6OM7jQG3DIitBKmC7csLiyqCyUrjXuLMmj9TRJ6iX
LXrjFbTfp0lWdmq7RGimOogO4qruzQgStB48hRulfA+N/6pBMziWmIJ1boBrZ9yZ2jiOV52l8QmY
AIt4yR1NBIy5v7JXfCSuB/rQ7WCY9A5UX0smR8TC5CdlDzRUsTiWlHrUfuY+NRtMEFfEjlCCwSAk
2vyrunv7cfiK4K/ze0Go2epZV5TsJhvjmZWtzSR+xE/470ySproJOmEJHqE/wkJ0cRjLrojduYAx
6G5PVzoX369YhP+9SgaPpBdmu+1yD1C4N5tpxqOnyR4EfHrAGN5B64uGlQaF1cuk4z7ugjffK9Cx
qlIyefCKQZO+NExANmOu+yu4INo2VFFplmjZocvUHGEnvDB4SFfFXOzAL6/U6MtdiAqO/5ZXmB9H
CTTbpfrMeW2RYuIdtbccLoa0tzXyW3ewpA/mWhC8mBdPWP2b9HzrQin5+mnn5GusjSmSbXT8koPf
ax/dq3iSNafPBRg0jUXceF2yy/P/e3/76rLEzoW+fiIUjxQKMk2qMwLaYF0Fb4Abbdk7HthTW20k
xhRMEKQgehDYs7XPQBVIRaQ91gj/4lPrdzFq1EfMx2WuNZ6G2w4JD9E1BRaP/Cx+qGAofdkR4Fgx
+alY2VMkeZoAoFVmoDmMb8yiv6dmDZ8+fghisYhaBPdnmap0vWq1iKNh4JVX/DMnH767s7eW6nG5
3UqgZPiRedTjNhXZO3gKsDDtkncBw99KQi7LBgugVCuhkk4aIY8BLE2narpygoXpMlnQx8xqg3DL
DREEx3fP6NWQwLGO3JhzKs7rVHJQZVcwflZHv4Kaz6KAQPslBBGFyW3KiOAy6vz6wi9EI2YSSRFL
xRzDmPV4B6VnrF6INhg97lVy+hLLeJ8t5EHE8CfXMZWENc3dWBAKjR6HppZe1cYHUTKQ1iCQyQAN
y54WrRD7U+pq3q5UvDQl9Kdi8D9dFM6WoFOAfj3OtZxOgGKH/kSPmrT9hCKbjfkOj1Ey8yUawa99
Ll6B9xe/bXToPfMfiuRaAjv8i88BJ7T3erUMz5MDHZs0QV68MJn7jNCr4G7rttNexMwS6yA8RVXb
M6JV1yn94cZRHCIbmuO0kAURrJKryUuCqT0MUCtQLmivwackTEDjz2MmIiU62i1vDy3S+/dEZSaU
05aAyNIZ+/yX8Jd8IXQlkD6Un71qlfSlZIT/GgLBH98QZ7WtNnycKQt9VI8amzULqsLltRSHwS52
1RPy0E5nrkkm4F9z6Iptfp1/Xb9gp3hQqKBZYlw1pzIa349RA/GzJdLr21JxBQ86yAT58f6fVAju
hYCBWATHwfCPMcOY1mIkhVGfh5O4t89N2t8o3U2+7XWfLL8B/cWHaKZMh1g2ZM65yOZOy6JKEitE
9gDDB9rEBHaWUXszlFTr6SG8CV1P/3fV43nug4os8tEa6OBueNy2n5yOoGZ+NDK5FV5uQ8nuB0is
tDr4Dr9fWXwwsDyShaqUZsUtzhoi7wXHGB+G4Mk2grsNF/zn9ZMyWC1Kd7aLlmlQurILbvzplPT8
XspQ6okNDAN393vVA3hEIKO0VzJXIptT76gEVwCwsoURsIwaRcuJpwXOW1T0g6wC6bU/cFYyD1tQ
kV0KZrBX+iIxzAE/98e36gIeOpHpFZG2JGN7UmmJCdREB90fl42oR4cE5JL60GhqEx61FLi+QBIE
VNzUghxCTWuhDLhmER13q0CskiiOK2fytaqvweT/ZsE9ckWvikYaLch3GsQx1IygAB8Kg6KNmHp5
CaZkgJVeye471xFKSwrLD6dfxNb+TN05FBCTevV6APxZ/CFapJBl3CIqzn/tAfTrdynUKzt9lYWF
3cF/EXNRkuubmGRmkOqG7stt6sUgtNPw3CbJwiMc3HmoRfQTgN44XCMGzeEggmQ2dc+z7U/7urqE
2GeFF8RXvt0iHC8ToqSF48Z4kHxRlh51nxCr42l6qwFf/vQX9PCX0wNbktWR1Cqpz7yhPdVtndKM
NBFG6QjrKPXcRI1W7juTzu49R/YW7QAVDGLJdrgubgddTjZZRMx/EJr2EQg7hn14dluuHhAiqEZN
ULu290iCPlhHj1V5tN45wuYlhKdNKRGqXczsnxPxnAlky8kG128TbLQDBPwAwPXCK4hmHVjZyQO0
R4kaMrWSLyXIwno5PaMDZC/W8pj75sdSFFXs8q93QuV+4XvcgN5CGRI47bpoFLIqO3Hlx5vDfHzH
sHrj7nRovxMiWMpEvIZay+fPWCB6qWNt+zIhS1lxF3XzC5U4raxjnLWeIqaRdxwQNLvCh2n0nASD
LPMyeVgwj5Wf3psEPa8f7koxst7j1vv5FOZLuQPnzw4h6Ehsis1Wlix69i/QtSLtrjgM9N3H2gAJ
KHHF2ExQhmtc/zga/HaQSwMUWbYWLwRY3NkoqhklRmaWksBrmYzY3fbA/EwlXpzJt0AkL+kbeCBa
+LN+sCg8hIFgREnwx5Hf1uNjVI8OoCuny/GG+XjPGWpogIUU2RXaNHKUgzo0uESTnKv7GO+xpwjf
jimPQuWzAeclkuovlVeJmtWdaj45aSqdttw1tmFgK2IG/fXvxv74KrkFqb3KTsRJseVFNp+7zf7k
HQdX1lyLSAyDCfj2i+MvC0wVifFfpNqiDCdQh1Y6R9pN345McT0kIX2CCGnEiAqz97ayxbh17B4j
q0HAG5nva2Xfw/rKRISPiJ817FXQiDGZXu4me9/J6YPGaqeV1aEfd7YifCYROCl4FYhLIjcU5cG3
vu3PGMV/LfgOPoZGYVW9MUZaURSMOBjh1hBKnk1oDMA4+xKo3j7rXav+UZfjaD2sLvEQvEjZ9tL/
nwTR3SuPQSnkRSChwddqNwfO9sZrxarnC1pUXiPP0IfLLwWCfQlK0SQQNRJfU0gN+Z79M/PhWKom
iR/R1fFk2P290SdowFBYtHSQ4oo39vjLLeDuLv/1IFCbYk/H0YCYLA8z1mZM2hLSw6SdQZ7FfJkQ
0LLShInvy3+4ValbGG0YHOZmnhYrj+kLX78KXgVErPG9iui+UOIjdO2uNUA2HhENRicfKsV0MK89
svLAEDnKCGy+1MMHN95EtTJG23RB70IH6yYVuxqRsvZoxu+Boo7vUs4KZ+znTr4dTY3EtPex445y
ARXyEiSqBwZbZybg2DpV2kpSyyx5YAipuNX+t3qYmWUl81QQPoyRBZBJ5cdF7xHXCOOHZ7NYqxmn
iTRYKJQ/ohms07XU4uYvoOVX0/oP1beTIIg7/Fysb1ms8L/MybqOPm3QozVH7Jl0rdbmYhIDkCMR
QV8VPmBYuk27HvFnLBH+8C2l6x7lvg4Brapc4fp5RR+Ml6dijNP2zSjyGc2/tZOmNA8m14TCPE0r
4aUQ7bezISGZ/yMTsPeMwAt1CLWRZ4IslgDI+OVU7fS+VfLUX7g8bvX21cj+Z6vniAx7uxuziPpV
IdEffQXg8b7GQ6t5NzAChPf/pKEoWM9JUlFM1XZ7pVurw25K8e7yWQ3n8zf2+TusjoueSF6NzwZZ
spwXcFL+w8+L2afrTlt9E6HqULTIh65MXHBxWD0Opj+ByzQS1tpxPiRKh+ykLWdtvqzT7BlcdBdI
il7vRPzlmYpN3YEi7U8kihvXW7Vw/TQLVG1SWdV5w9Rd4LfD2da6YUf1kibNOnt/4aLxrPu5eGtJ
0yBKg1suj5ZamHuDCjJHpUOEVchseoUxXkgTpp7M4RMyUOTtYrgRZfNgwcbWcRXTO2LbJJz7DyPc
GlzxIeF53S0zm+0gUl3XeQTfFRFIZFwP+mVl5GzH9r6kDQ6AYe5LGI/tioaZiwhPJLCHBCm2gTuM
OwzOoUPpdSvyqkIux9eWzUNtOAAU/SWsEpdDa9mqkaMxTexlUOGWDKC2+wsSxh6nafcw4AN3A54i
l2beVVHqnri6PlPIObRCzke3fmQvUjVNqMOjnkHieWqEoFYSjut9I04EEsNO2ZG6NAUjGjnahEP5
eSJMi0Qz3XpIEk9QLGSFuAzusK9J9asBk9VV2DkGwal+ybh01LgehgBDEI69DFE+sKJ/uMinGf8l
Gn07jl399E2ZfMH9wgoTAbxSVZR2bsmUMaEdMKB28RAI1e7tPJrYQbQmgoOkIgpGPCiLS7Hfm+KS
pOFkoWJx5HpNOZZVBk8dWP1wf/6PRj2p4W0q1eX18lBWQx4WtF9pcu9NCQIRkh6njnbTztgNksUr
d/J00UsWmO/PMhKnnxs2g6MruhbL38zA89SPQCI+du+HRsBxmfpPxZ12Beo4MJy3Q/TRcduD6tbS
v2UJUtPrI2/4mi7o+m/q93R7D9XylUujws/EY6m3bQ8sXloZLnW2DNaxK6fDYwFclzDndILbOcvh
nZYoOkl8ncgmIq8bMOQwepccTdRQ64ir1lUIxe5DjqAqSLkVBNmWg0axg59wCKfn+9YW28FHZ+ov
+FnnRvBzi1Dcyw+e5yAcjF8cmQ+IQoomfTZwGMYU3onrVn8FzqyWua7+QEDqMCqKUa5hxKGGayvt
bEeJSHadOkj1F5xEtHuxLlkSxy4WHRKFz5bCqD502QPPX6wbAfWs0sx+dB0t7bb3K7ztW0ihP50I
c0/Zx7C9vGK6n3T5TG0p+rfXRISscO0rgf897KGerdQU4J51jXsYHVeCRC9DPrTnuVv532AmTxq8
1rlO+FSDL9K1TmgSNUu55D8r+a2mFDqktaBsceEM7mb71w7qpHQmGj9WDNJxJVpejxfm4IN+U6CH
k2zwXRPnTc/LxAuMiP1xlqjIa6uTS53RBjTAaff8BBSfdir5lEPVL9VsS+XamhJN5pPIRZb3lcS6
VBjej7NYDCGOkubNsgP0co0SkUA+ptg3cK/Z8A+bj5YHyoM9y4pNafHA3hkt8c/meervb6x+wdMg
3jvRTJb3L5wDHq+z8ocsYNXulHW+OLY103PtZJ6hAlg3uWBepsYdxLPiOqGkB42CR/TW+TSpaRWM
qxP4bhBkx+EuLd03z93oIdCDpRuLGObuIOWgPpQqZRJ0rkRzQyDO74cT0YxssZ7owQ/+t9/QPnCs
yjCoHzL088RLhqoQlhNaHN26B47iUmRpVA/ZbE6Sb1pH43ivDLlen7W3v6R6DNEs9VvSx2jDY4fJ
48Mdgr5wqjwtmmX/91lp+Cd26BBt6+dYtr33O17GHxmWHlzMTq8dgx1xzOSIWM3dZAIjL1QB72uI
yp/zikM3ChV0TjfoNSkDLxp/w1ieSPiH+SLxMpR5zcnXV5wI2xXUwfUDZfAbCZQyEIDJoMm14yDt
LZbKH6YwSIgCjZwnjFbYphV5yZpyBwCeBqHh83M61u6zdxlsSJvrZJspIZdntf2+ize8sVFCjXDe
zAMpI0jyF9omnHReGnTHu7aPuZaLp5HZb42/KbstelvOJKviiVqecqknVRXe8ag380QLAHib7wf2
Nd8DPz07+8duJNEXtk5MRngNJ5h+b036NMmP0VcDYc25jkD21qYTHSDcWIzCqlVU9qUnmJvF0GNV
1Bw5PN8JmAaoMDbSZ9d6O47hiGdYmiusK6mRAVugCHzRBhe5fR8lb2UitIflnM6kvzCiD2ucwn/A
SHY2dfMw/og2J9rLVbI+1Sj1pe/pC6OwF1HyU7lG4GZtcys8BUgPkeBHtjJJkovotIPzW4Kegm3r
AzkBhNf/kN8iJnLoJNar+jGNpWai6AwLRyHkcAFk1AJ0dtGdIdkkEx8ZMenbBJTFTJeco2fWVq+6
zs0BTB0TpoYwBQ76A4XHAOQnQ7cPdyDxIK0GFdEpcv/P+Yv7oBGFXPxbICtzf7evTci94SSpfMa9
BetgcTCYC4ImwfYqE1QwN1sQiP9NJzUcPKCK24L17HCxsL2a3hUKU+/ymz9H+QqfnAW+dDp6fYsa
ERjiXbCnwNN0UxLw4/IEMwhMROm1EsUEYFEnVW0cNzFndLZI4V/OjubRY5RXli638x4m2sz+n7b5
kwm2KksvEEljy7IVoMUVfRcFC1eTDz08rkPB2vW/2DEe/N8v2ZnDhcE/qv0EeiUAD9fhkD5XQBum
hjWeQaATiTNEBzMqLojygHPBGPOr7kf2NrJ5zzfoWvd7L1GAwavoo6mcFeEWYfHORh/TnZ7Fggpp
FBWbixBC6XNnEb/z8C35sK6SXB6S3c0sQpmF4HgOStoyr4XYydTrF42QdSNUx6sHawKVMv8zPFD8
ughqOo5jO5g2SBGA8YXXdP8pNiGc28iddKxVwW8/Y156lMHbkAYbwKj6fyuOwmLhDhMwuTAOnn23
iPxFy90bv7VEOUagU6TTzdJrKt1vXPW+aGeShbnHZ989Tp7mOep1mtJ/PpvQNboAj3rYJUpRmCOc
zPy6a44YZm8PLomrtrpGcVZKG7/iKQr+Z7cg+54WzY9npNS8PgQVd2GOmWeNjeNpfQi+p0luezH/
uqP1TV+wUb31mUe1Z8wXva/WR78EbpYrbWQCvlP7EQzNIAvkOWII3NFHba/adJhF/3l+hQvHvhG6
JFxnl4po9Gf7jjKJ0Vioivuxe6YmXsBVpI/7RqrrU3L0P4/HfOhXc50XESACnzwoVWQANmQzQJTn
HmriV7ve0H7SdccpoP83Pq483zPCf2zpEiSqdsZR892dyKCSLo5RhAfjcV+G7ox8vIIoZ6mO4YBw
M77d6U1SnxZ0/KzzpiMjqlnZHn9rOzyNNxq9n3iDmnoPapxGOcGdTnE0l11iIMDwb2qrkvTfuA8H
lqYV/BFiXaRsuOiepafUt7igZAbdm7r2Q3Uv64AikKX5Cq6o35X9v47mH5QcTPKrciavoAq58jZ7
i2h6oORmS+LETSkTXpd1EvPXknFzurFXblkbZaQ3JHUc3G42Lud3i0Xcrn5qXXO5FO6MTCFtfNzL
04y7tWewcaqwSmVkI0/v+ElYIjkXX2BRwOEzS2mDQsZRFc5WRVhUXgHHGS3Skp5PTUg8+PWSkREN
2kqWUVncuIsbBNJzula5W8E02uJoT1JWWjcTkfni5SDJKlMf3+UAbVlOJk3bqvF9MqLAWcpHI/r1
RQ2sbh1sGnFqO4ha3Fm9oHq/ennKNPJRuZNDGCZ9h0SvVclxXi3xca1kOrhiZkRD+3UpxEeocAJ/
JF7y/0OSyq+/R7forfuF6y4PjOPnUrzjrz1VHO1gq8ktn1TMgpH7WrzQbC9ojKFB/vbCb68qDi2V
W31QzPAG9y2Jo1On65OHjglAHe744j4OMYumRQ3XAT5lo7ta+GgRDTU8067C6AKyLsSvVAXCHomB
hSDg+oBIP/h1egop2wbKoTlovvWX6UQJkBoHlNaiCKldCNc2GZIWvoolGh79B6V0lPQMyzIWTjaL
eBVEpOdIqflrujegugjCdvH0YnVFEUy86iPnVUhKrG6Nh4OZhbCVdvRkiaLZcyuuSxToFNv6qSx2
5ZSxH5d9WUaQSOEa5wW3+SY3rihPn2rtnwZDfOX7YKelhfGusRaT7mXYIyG/gfX7XUnSO2zIyRdu
UBZdjV4JvBrHG+HHyxcEEwlLrViu6uXG7JkjN+WK1K5Lb6th+bOfiGckztCbD/LTADeVNcIByAo/
hNyfXWFQkR5QGmefwe3kqZ13hoVVaPMD3dS4QnUI/F30rEyw1hmH0U/BSO3z++tr/t1MlnL7zYZN
vf5kQ6l5AaLXbgCxdS/nZOO9kqtPhseM3PPZmXR3OVgbon7FUGrp4hUVlF5JPIBNE516/UnJY+f6
E8N+3yL7Q/dJsjCCUw780QLpnyAHfAGVsXAZtvgpY+p9ui/0GDr/RtNbETK6N4U5pDPoFJn6w3Bd
yox036D6Ve68X5DsrnHwN0T82gCcc01F3ZcJ4lxKPWcdk5C1xWsMhzJpgyIbNP1eYpTvVCu+eg2k
UwsI/oN5+G7+USj6I3oXRi6q3IVLKjCoT6q6uC9oTXoLzsjOgF/IhRQ9DcAII5U6c3m1rFMTL+gm
9If5fGpp6Jnf7lTN1dY42PMPWjm/pxMct5Lp0YIrt4DhtIO5rudUWLKnnE83ik656AWI5RNmrjVk
gnOjPv1ZqqF3fsoV2rxfTwtTjXa5hlMbk51Tzr10bO3Oa9Q9ssmz038seg79Tm4PLB4vKjC5Kqmz
vN//YswazDkoCK4JgqzfzVE8ScCbrCYMh9ojwdI3R5CqJg3saJCIcBr3f9u5ga19gmyhYMy0XeSg
6GyyDiQAOYuJieMRSug9tNjM3oPOK4Yhhdq/qmJxLvQUJvUXYn542yzJA24/ZqoNwUe5OHS1fQ9U
DmmE9I3zAqCVJc8SDGibgDu1BKDqII5Sm3AvrlmExlrCcbM2HdQBRMfrXCtxYOGGBYA8WFcMvRTL
1ab6vMfSfsXFuLE2eorMkkkIke+5umiCGwjoQwhVl2so0vqcm9B0lamdGBfhFPhAwwU9WiBoJpeF
e/7kA1lF3JEmvfGHF0fIm0gr14vhQuaXcH+MEXhvgqHqbcZE6VzrWyf1FEt9K+TEGL7biZi58x1L
bChKt2INYzk72UFZwTMs41af+B+FJtYLg//NS21YAslD64xk9g6EFswyaT6HN5Jb5SLYZeV+GBW1
pRaf4UWtDSb20j16KIBiog7L9cyEywcNbGlFSDHXPnQ9LD1pO9ENLP2DoLcB7CZs9MK7kg39hDxG
tkUPmdqQ5qY+LCruOmTiFK82AkZ/yWXflZTtwOk32hA7xJNTaF2U8zFlrmZODahUiESkaJ3CQVuf
4JX8apc9m8tU5QNoDSh0TzuXT/ecqyrF1qWsJ+tJirhKMhFMLMlFgW9gtiX13icvD4HLS3EpXva7
o6wr2ZrZgZWmWHHqiWeXe/INCHOnazJIxQl8rVLY3lCpJQeFJkEmDMlnHuaCD41iGXw91lSV9LwM
T/p9T0sShl9PVbClZjvQ59kbKFBiBQz8TRSv9C/+KdQWBKmn+OIpUkM7XVBkg/qZ05E3gsZTEzLp
W7vr7RAWi88owG/BGYyxKrcX4lZe0KeAs4tqt+tl0jr3frDAOiikC5qx/6n+C5hSB8JxmxUYEbto
4d/6Yp397YzU6Oim4ioBlCR1pKdGrkjL15Hz3xqIKeFmq0Sh/Ed1c1w3a803eQzNglzVxbult3LD
gnFIJywI36ZYUNdvNd6toVc2huq85wUDMxzzZf4Zwxb1nAaV1kIHF07ovjsnZ3J5pycXGSdDGy+8
/LqX5ZmrrnT9ch/awS/PNiL7YmtdM4XKZ53n+ffRF1WBQTEtrr7ppFKZFGGYaVQhHXdyiuGAnCjG
Qxm7LBIjZYzR4CKaUlAgLpmdV1TF8kyTyQHBq3HcybqwU5XYKsRkG+G+EuGh7djDTUI9mXmZvpt5
s3tXZFU3eI5/0LZsoocrq4Fa7ecpr8v3bVLmtMl+3lf4CgWxRzfQOcU2u5ySSZEA/bP8V7wQ5PT6
nDwdAJExUgC1quZXMltciSC6HTchE+y/Kw2DDE2xDdLx+X7T2ltVZhrIiXBeTDSyUS7+9f6mcOxB
pT0EDfl0ezVSetj+BrhZkYm0F3KmEOFwD9g/iVIBqaHNvVQn0f4F4NQsDD237MidV6dQK5NxRu9r
GM/FbISXYADfBlBmFn93ZXKd8sOWPEw0M7CsfnfCFkbnKVv2ZDkuk8XplQem7+3SIsM2Tr/xSt5Q
FMGecS0rQT1GBL7JVawdSNoqO0TAAvVV+MZzdjSfDncg05MK+/o9zjuezaN4q4iNyT3V6pq577hb
Y4d9tE4KCMDnOL18FJwmeCpSOWJR1nhi2ZeVAdOpQuoprOWjAk/c2ZmdBV2q+Z756InTt5/Lyt0X
66+bM/SxVZJ7t7itFiVrEvinXL2lTivLFZUvfiS3lqpVgggJr+Nxt1JHjwMU4fnEuwGk0CYK9l1w
3S5sqIAAqdhwigdmzOTPc5cHwaZZWTtesJ4Sr/javEKPilBKno/hkP6esyVuRErQm0J5jDrsMm5T
EjYoJ4CmEP1AIPBtg6sDPoCgfnXOg/j6Cqr72063t515RCDLBjS6lfL/KjCiSdWS0tVJOEWgZG4T
B2yweR53GtgyW0aNlN/qda/Lf6gBBmqoKHTxtF9b1ixygKXKVgoAyzj50iihrb2CwrFSUoNsTA1j
a844mtnzaEy2/64s6QVSsBlTGsYkn+wTQFI3391j/ft/ar2JIrZf+MSQG8Ow1iWMlAV3Xhn8tiYj
wmapdwGVBylkQOXbvmAH8CmqcxglU4GfMMY7vNzYfOywhAKbar80XfiqhJufW4nSjbi9P82xyoE7
9mxAkeX+LEboRlbiQX5tEPr+/V5QSicJBicihBrSA1OfPUw3xWS6O66lFmC7rmRPtQfF3wAveyAx
97ENDZnjFhAmixdRxLE30+YglOsEeHol68Tucm2x9iq0/+YU9zRTVq2Yq9+g0WR9NnQvvCfUAGuL
u2XHPrvHwE3MDCiVc0pqQToH0lh7S5A9nkHBf+zCVeoWIejME8cgFH0lnCb2z3jUWSqVuNlwELb+
1HlD+nRE6lAeJOrqOtWVkDvTLKjIfym7qE7fyxTSuokganCMP+T3+DyvamuIT9cWPFSkyMutZQVi
ICynwPWTSN1guEnCa15waJ/5jZl0LYn/1368nqeaBS0wBmNV6xECXNKxb9oPSG1Cq8K8Ity41K8q
U/xJtXyvbWKcsf/uUJ8NJIUOrkGJPqKkbqMfaVcthS9/p6louaOzLAC9U/3hg5MLs98ZkrDFYWvM
FcCgCYBt+BzJ5eH02ARoEMvZhxLDcFHBGSJGbV0CSarfUtIklf1qVRIKLkgb/2DzuYftdkaVEeKA
mvKnBwvK1cnEo2Q28wScTUNHN8vpFpZzZUEzgYsLBbllb9+8eTTVv8VrnnpzLeQ5eVfRn2CyLWHy
P1GPexPrya4RPKEtDPUm54Eqmuvxh4PZtmygL21z8msJIavqdjI/UmhrXAeCZOFxSjR+6UfcV3py
/vlKP7D9nRlGC8pVPpg667rcnYqcI9qt4zrWa4SSGeTLlTZOsP3phqMa+QGtm/f+h46jfzptGT4/
wujv+7eOLJg59BDbGfJX+ep0/PYrPNMLdi7d456VzO3fOVXzpDOwCemIOnhPnvKx7SApn9wm+Jsk
A3uKuUnjrTu7u9N3N5ddFKajGQnl+T6SzgTtLXJvYbFSZ6iQYCmyC//Gvqhncz+A7nTTQv/+579O
AQXPPmxa43EoxYVMe0uEIA00rWFG5hPdZuNzNft6/EpF97lMf2jqlnadjpSlQhXFxamu1QY4KMV+
NJ6gt+8q5kaVht8wK4hRUR+U8Xjxz4J5t6jkgDcihsvwez54v1fGMsBJQedMouvgN24IJN1XO8B7
HE0XSO/43v4c4VwCcFpXH3YSV9WZ6KUgIiguE+NeAUHdPGv3wM5gfNAwjh7FYf034msGgx0XCsJW
uuUkpiI4zaHqjmgXW+IIJebLFW8GmG3GrRtrh3wBiOxHuXm9TUOF3oKSS2WMxu9d6s/js5a07dSp
KILmjB5RYPL4+fyz+6SKHcbCAnZPMDOBmIXKwRbnhBMdpRFPRjO2InCEWcdALw1rgQsOs56vG6AJ
5cI53nPAJPXMnAvZ6Yerup/R/x3/thqZJLwGYCtHKNj5BQ5fyeKZHuSOEJEIPtz8e4u62Mj8Rrbo
AsZwA0JY/lrtgfvizF5/QOBCDxnQr+HVyDQzJVh/VIBayYgtqDuQfQF3iGgCj4tizE57mVmf8VTb
s0OqIcxjbvy/zH669GvGAuZZjf/RK/SewvGSfFvARRnhpLzWh9JBotb3FGAmSQ088EIbMt3+33xM
ZKjuttbeIW4OFE9LzX27EjsUO/LqVwKdP5GcMNlT9LzFLG101tKTa+46ws1BF0X81QbjRKiafxX5
QYbZlNIaxJwdsAOVSvMSbWgQQRgm3uK1BTqxUteqSrNCS7u3rkmmo4XRA/YvpqN43LO/1M5S0mIB
jnHGsEt9MaclW319K0GfWh8gtD94LCqVzWYZjPMLq9oSb58KWEYBL8iHWUZWlVJAuke/8kevQi0+
jH7NTic5mrJxRN5UYRaqq4qR5OPyV46/MykDKh48XMYuWJ4pUODID+cwQhI8EAG2tMW1KUhbCJ5s
QpItv41xjDr01mldwq+1+iFscO/FOvuRxjc0gLNxet/lhDFqYZ5ry1xP6h9WT8Qf69oCJJMeZyDW
FTIgLzCnIDung2UiXlqeeehm2ZZGVuynen11ZomBwXHskXj4D0n6yJSVRu41HYoe94eDkDbP/np6
LAN3l/AbvgAdB0+Aqk86oi8ja1XXAePLaD+QvGwimO05mXPtsBw+z1rghwwtZRzjTeAbno0wvaV4
bGFZ0CJKj7d8IoAsFLYieh6nh8BWZ5ZtWE2+D4GUbxmlW97RD8ElWrM4ArigKmt31YnqiMlO+oOO
IQjRGxJriCgdSreK/gmMqkW5u+T6VSA8vMMxQj80wcPX81jAR4R4pZdi4YRqJw+aoYnyOQSkFTo+
I+fcdugcoYJPixehysXHYG3yxxwgcizrpfrRgSt5mvmfIZS3SvC1YkDzx/cuh0iGLk3tjXPTlcUJ
Xt2q0jrx7K9TeoQgwd/9Pli4swbua4xjIbT4U3vHzVABV78YPzl+cxTyGbJG26OF2l33qPEypf/Y
ue5c6H3rEOtMPRU/7tuFKASsxkuujdCG9xY+JbujePAabTuvkzDpww+IZ3KQ0i1Zk8F/MsztQvZc
nwsQSMZ/n5AiQad6XLsds5yxlGGLYKwXy7QP/ZM26Z+VfExaLNAjd0q2VWkBeKPSmEnUuhkFFZzs
Q8EI08pbrl/9kl5vcAL0pEgukYDOaETbp19Y16ddh+rGySWchkukHPZF7W6i3AuVWtWNOEgiSNPv
jMHwVtNuZmR5WI9eXZep+I1ZcfX0M8O7gmFT7oI1tYBD3/GaHGp5NbhDlGHCpWrlGsVY8iHmjjy1
jRKYeYD5iF8boOSY1AKZfCO4AdFif66C/YZi+DzocQlaxlpQYJw+Bm7/Qxo3JWfFq7dPeWgUh0ID
vgwcLDMU+UGyxFYrix1YyfbWo0nhasooCxzdIo2vlCG008h0I0B9Br+gb6hhBo206dFWOn8UoqAu
mygJdN/9T2lokh+hSipDNOeoovU2Pge/y/ykEDY3MjSN2mJ3yWCrXnRzU5JyWGvu1CmpDD2Tu0yu
Tnqt7hGpbfhnR7LVwJ7enwSTSh1xqG8XC9ec36aQmG2b75ks8mwcrTYDefrIKdWqAhu+DNOmSNpr
rluvrGNUtEPc7WlCulioXiXf5cAQC9oczQ825HCUZpC5/iWuqrSvqHmEYTgZT53z91yttkeERZ1V
K+1vlYQAxjULUJdwXrbl8JE9wjU4ZDv7gO3hbNkJhiDeaAqkOVi45lOwAIEdnIilFlw5am6tiYfn
dWOS3tJxCG1ZQ2tkwDy+qhlsXURvb+ecEBRbbCwQJxd/vZsuTniFPEikBzwta9KUsXGtBuZYZTtC
rwXBNI8Wsqnu4lEmu7Lcjcno8qGxobGvn4Uz3oNNLZX1WTKcMY10JMQ9DpREPWSU5iev9FYXl0HB
54Ff9eJ+LAl7NQBNJUhN47U9lIVDONIcgZUFi1c0zH2K5drXGnJ957p1aKoFImHNZ1/yQft/1QYB
dYCZbVqlqQicdlbWkCjVmH/jQjMvc0L+ButVjngysZa+BSakYTHiYjG5+ELZrsGWuo3KxztSVxrB
oyvemG9vvEwICgWiUhJVY+RaAK8HtSD4JnNNRipT+Fe7viiDMA617TG2jjno3AajXsQAGxb4zx2M
4QdxRMA9BToFSbtUe6k4FRbBsGHO9c+Ly0PPNCN3REFnV9faIcvlg5zefEEKh+bGg/4DnVBoduH7
4kTblTxSCdYDkCCpnWqCebe8Pto41zKiEb9mspuqgl5Qy33DVyE9gRDW1+u3EjcPd5Ep42fOhsjU
4zie30lf1lFfISCg4hmpw8pVk8uqjntvgwNasP9ezHYKLiwwTO9LLjV8Uu6M0TLU8Oo5xuZJD/SX
ym5G2tf1W5C3kJ5t0qDlrPvX8PxBpLXLpNSpII6nr1BFJieWueSNXC3Q1iLZIipMtquZsyiWJ0ru
SUkObZ92gZSc5wVDL6qHE+UhFeWb4zn4teELRmWOq0bK+gTGt7X0RdifVy6LA9d4qsjLXz/WNBk+
0rarCrTdsZxiIYFguCjoXwPpSxCpY0QZLofrgo+F4uhbpGl9HOX8qB+S7oeD5SpGLqI/NO+94wXB
gPZsaHrfQF922jqV5/y+bplrD4PFBMd0dO6EY6TXiAgU79pDs2ne/BLymx3FVZDAQS766TvUYzKG
hpLcLNyGgsctP67jTij00Hjw1jApAUqH6aQA4h1G5v9Sc5Lx7nX9w0oi4LSXP0Li5wDCXyashJDd
9qKQUcpJAKfvO7qdSnVn7O7tg5n3SS70WnV6ihG3CPgw5ArSTdYkGexWjyrzp53txzwdEuDCx51b
Tou93RZVc5H1JZO3NFlZ1QeSlfWZr/l2vAYZQRheOmUSiSEOLjfSYAw99QND4JyEG8FyVUqQqQVs
RZPuWD9oBdPi+/GFyn5eMCH2rlx2yS2plmO+IadHrYJcNOQilzTYqNUvNNkwH+6eTLSsu8vDE2QE
NMjk4rdfyO8mclMQ86TZ1uHLnVdqxCdc9ucV1anybzHP5O8SVtk6ugZ38ebZmuKcxSdT3Xuwubni
JojC0aeXO/n9HNOPaPIoaz/0yAwLQiNe+88G9lOyy/el4ZmusQ10Mq1CppUbCk7pqvA1gccF6kbo
7CJrBvrAv58rGLsHw0HrOxebXDKQDy4c++nqUYpaMxWChomxtomD+7GdebDseNRjr618kZcjCvRf
V+nfYZps7uPCg4/LMrJd6wXsoka38oeO2AIdMLEoNYMvWznvY0Aojxu7q8RtuvSZmKLM+KyjGfaK
SuocqCz9vBa+G3eX0ny6J3hoXrlE/HQxHo8MZEPyNWtySy52Nw1ob0mFkjXcC5FbiIQ6azCtEmlx
OIVZ6s18q6YLaBIaaKl2Vs+6WO+x8VB9nocfnCcKNJknK226CyR5WSbBgjhkieyTYvr7I/lphTyj
zu4vORFSYx2Zj454FuRuOwMDgkMVvWqhO+lXKOFeVfgXLzoL+9SPiv5MoczWRtshKZsw46jkapKA
uJh976ZLUeVLpHTVfHGzjf7EADanZSAiVSlVukhEk7hjtZyLLmz+sT/Dxs6clK2JfuHNIOuXJ8r0
vo+9UcqFfeFAeiKWturu0SGdrBzfVupnpiNazvU69vhE4Gr79h7KzS6LU2+lFGSs/JfyV+aIUvmh
3DldLSmhBVcQsoyxf9I/BRVhnA5lNCgxYfpm0EHyjmEMhoEJkGQBJkioUE/8Wcdd4Hh3oNw/Os65
FI4POP/vcWUIucIAQ+oczVt+OhQcTPlivQqJKu/HkR6E826PWQg9aUStWd/RaoWtjMYv+D3QhBeH
8WMcWiYgPPM08Ov0qDRVlFJhqUmXpfO6JrxI3TGnfJBZM/M2gBWXuAQPD1xkzs8GibuoelgphBff
hhzHiwrhl35GJ0mTpTCkcA5BclGwUhIKSBjMCoYPReKryf7RC+ppojmQDSqBDg8j4nIfIN1B0Q7e
TVgqBLQbJ7weLOm1TT8VhqnhAloXKRAKaL+UPOUk7kx0wt3C7BvGWA7UHYo7wASvpMQK6dxFz5Ry
QzNK3GMbmExmVmabgQF/phuxSEM+8XZYdJkrUaK8dP3Y5Kiajxv+rte+Q44Bs20Dqt1LKZimJsey
dsNQPtLI0nuK6Xa2G8cgQ+MzhZc6JwOyCN4VuJwLsTYMYCBjtEOoS3s5LHs3etEFHB3XOBL4FqZG
wbbCXRXBcqMO/w+WTmaxrGlYEgVBNgxaGg1wGPOXQwmeayZZJRFcgv8O709Ja3d/RLy27I/bCH9B
UDWBOFL67rnS4Y00qOX/67at0OCpqVPMvhk7gNCSd9wrNe56yGd2TZ56dY96uQyOWb/N7zV2iB6S
rFjgWkKHIJ/Fzi201GCP9JBeEDjH9H6SGVU0bCSH3hSi5UDCQ+6OyRsOTSlZWd9fAhdntv76r928
GQhLOnArloN9nudR/PfKcdYsChV51oKsMe6MBBaOr01s94nxk2D5bX4h9YoUG4Vb5iiwt0gIlkMe
RV02vaR1dOBd/ktM2qhdHxbs03fSuXtb8WYHpU/ZcPWtnw5qYIqzh5bWGZLJVi3PZ3yyBi+HZWDE
Oo/3y9C2F8nl51lZeSMj9541h5jsL8Cuqzr+5peYOSsqPdxbPOxu9tT3kyPS8DGX1Cs1KbhPPSN7
CjtYSanoXozLWeMio+obcGQtdBVrkJ8PPDnSGYdU038hy9FL1QatAzatzDtxDMZ9jSVTwn2/f3Xm
79p0eRYlDDqjNFD8f8WBvKstGs2zASit3cpjb0GMYjgAd5MRci/oA0G3PoYuA19NPa8qKUl0vB4E
9KGh7p3jeMb4l3ElQqENbq5JUSi9/4eSoAaRm0YeQxUOOd0AyPHqydDCy9c1UxR3Npi6LirXY6qA
KBCOjD17rnrqnFY1FLmW3HK3SQA4g2KUWV07bENsahQdrWvlrtTnduKCFj7RpvZBfoY0R+PXkZCT
WlF0roKJyjXZEaxJRyURKrqKxXrKwkHCiVavTSADwdwGivNN1g2cYvNXpa3J1wpdqFjfU7LOuZ7i
ZYptNn/h6UamUEtmvHB7t/Cvg35lzNLHErwPFlA/eYhweLE0RPNT8UIph2f6DEpmaR06QX3AWoiv
tXBVxLR6kucm/ppEj/bSW2jR7lWPzFzv3p08g9llDYdIL9VMjQJ9FtmMk+uuIzaa5OL2ULayMCu2
Jd+1dox5jePSrmaiqehX81PqbqfpuJslXsT3efnGKbGAg4cgaBVkqUBmd0BGydBRFLuoBfRV2trz
VDHDARkLJ0KTvf6C+xWzutk9Hy/wM/gHCBXSLrF7cLpofgHfN3KW+xy9eOOdKgb3NSmJ0aM7a5SV
ukUNMYQDCRFyDz7mrZxOx8IkzP5YcTGDuD0FIEyLmdU5tVz+jYM+J7zmLWg9BSNO1Bi0/h6Powew
GtfswV2LrgK943rLSl0KsFreC1m6XPYS29z+InhUeQ+3RSJUtHyyxgwr6I0rVOhkCZIcomqk8Daq
6JzOumTAK2ePmwZv60WW0pBAXhmC4xpbqatwobm1qUWRpGTnX5ODWfEZvJn1089pjWvSemGIGKCw
HSpcAy4DPFbzd9g8Leps6Gwi31IYbuZZ9e1HnTYq0nbp4Dvu8aoRBEQdBbOvGaJ8PrQr0nx5NChc
VHRM7DX88ey36V3EP/goYigW+sql+TnjCskhiMoQLRlytGvbeZPiCHshw5S7kbroYtE52qrcnm7c
4KzZ5PfoBfITOPaSkdhpbx2AgT+SOZmYJWlHk/0JJ/ieq0rv43K6c1ksQmHEqjjSzCljcxRWGk0f
61IGnL+cLC+maIh+CBeURDFegfFsRZrxSJHXYdT4P89iEaR/cP+dUapOY5/kibbhk/H5B5pp1JNK
139t8n2WhngjFaBxO0HbQvE05bNA1t7QDdAVy3fBRqWxGw/QUA6w7o1IAewZRq2ZZwgt2E6U15Pq
+DBNqSRTbjsm98qumQBEInnbbNtvhsdDD471ZHAKE/mMb+Ad2Q8JR7oZ62T/H/1O1m8HcyzZ/9w7
B6X9LqaSg4PexTpMUh6hUSkuDEU23ONlgvPBBpd8DOleHc9YxY0eh8hWssw3YxLLJRrEjymiQXc9
Qkaqv3k2cQgC/kKbiKD0Ey1szXBRg4JI2vUlBoEZe3ac3Tu268SKeG/8nX4WaMCU8r48T1tXcl4+
Mb2GHYJC2LvWSabFH2vFx3OBc7EKrNT/bNAMxiYGuH+cvegks9XPin+77yej3gq2ixaPUE0dg+4d
cw8ZMsJGXwGw+C4gukmTjVc3JbpGCUxyWtu1FKYDGYv1b/qqqqUj8lKE61hoMmQI5/+Ccw0IHbTh
Q0r/6Bvg6KAo7b/FrR4uXwuTCFxTUMx5c6xjEmWXJhrNrYFdkEIiRjUY9svp7nvfBtncKG7bVtuq
BGAUYu2MeI0RDjmxnqTw0q1ahlqmfn2zZv22F0CZndlZkU8fx/v5WKoyhalhf9DvfwA+sm3J4xhN
jmZSW+2GqXdDlcn584IScyIx5Ea95jQlicoiQ1KH1CaYMRA0g4SGzfHx4qyGM3BiEHk19S8qrGnN
xS/XxePgf3NUIZnZuHMAU4KBSM5QrZfOXUJOnz9VCdG8UtSRew+mLWWmFgs17IRhA0/kR4IkHe3T
syRoMomtpWGxvsngc96NSoltE7wueSmE8lLrQQWqZbmWfcBBCvE1PyhWgeBkJgBxbgIMLGqvqLIR
zzFjyjC05k959jnoWRMVnBFSzOxFIAlJrFUszRD83JnXk853Ne7wk1/miRqwfImDF93fUYf6ESLx
0nGMLHMWhEoJELXex857qY24gsbC8x6yxZKv2GhGhVOjtE9CZgK/QvxKvG2QoR6mLxGnoPt9uQAr
r/AX3opKDkiDhRGmZBVqB7og7e+os9avc6Mg0ByY656jRdWKKdAPfNiETFJe4KfcGeEBctgyc3OE
RfPmEu/3jErDNSmDZVYQbsHXU/edGSMGD+BRX9pDl+CHCC4WZCNqy2MdZihN8ILGGb31SPsQN3Ic
5i454iYvGzLyK0zGgcyobj/jZH7X5eIWnbNxGMI54r9mFDS2QDP7uDrYnKkzUOOcsI3KQ+IaefVa
AITRkVgG9AmGg+amAjwSTMsXZo++fnPDOckDDl5opPP4/j0AF6yV5MU7Ir11sLgyxhnN4urfkDq2
2wpJsTQ4UuO3ALJv0mvB30EX6eAzPoW+wwoyo9gQgYsn/P5gyDPDlL2XBM0ZoE+pVcc99qfro2cH
FniXBFdR/paI4w4rDKL5U8bsyZDTVeFmTjWPaIORog18nF9g9WVtWxKJ8TEtL9Cv/njowouTBgrO
JBUYvioELMSe+GgraDB7RsRUcmP032kGqctG1c4e8MoYA9R8bUtqGH7T6jEYgxqICENNIfIzq/ou
AiJbJ5vqgo6jgWH57qZxHGkVno0UqDxqlyytA+JO/DfOTqx6feT1SCKrg3J4+Vv12jzAobGeNPDF
AIYxzwBHnAEBI/WMzM+ju5YzldVE/CtJiBB74Cgllwi8xv3csmIIDzeqNsBByZ+Kbv484GwEi7Qv
Tw/mej8syvZGxPERVU/Nxt2AP6RCyxinAnW3nzuYEvQpogZmwn7ygr4HeNSUdgkgm2iHqw/IjaSO
oUfWwDLtOCS5hfHLAYoVxJa1xB4Qs3krRViIIS2OHoCTSq3+w7fEisvD2vKX4HrXkSY9vFqOrwuc
U3h8uSOjov+V7ZPifDzksKTwdS9JfdRkSEgtwk6f8V4OV1gHXo/CUhu7zheMI+EE/AavZwkxzQI4
xM5Z4rv6qgWuZ5otI5yYHx8s93eqPKXJ9xyl6xEoG5uM6HBQ+6hRi3dClRhuyJajosrEXqd5Ucxq
2Ar9TDnWkRCLqcmStcvmR9JQQB9Xfgrn84AiNpuHcwHUBH0t5CNjxbOHwJuT/UGCsEmboFUmFmIN
Fkm1hkSax2os2T2kP9YPDbKbOPJisMUcLl7ysg6HDrnJMRAUXpwtMoMNaOLvqAhJk97OHLUpaZb7
o0uTv8Qu+5GlIFdO7I/1w4CQnl8d0yG0eeETAC+px71HD4CFiuQTCBN5PrKUh7uZTcuBKSwgDwqE
GeYY1TlS/kRjRxMTQzgIHRXCe1bAmeCXvmohXE3ndoGLyhjQ1A/Al8IgBqvobOmH6HHtRlXc+HMZ
c2I4d6rigWq2rj47w77AcOl/fybXZ9sbOFCYkpZFjVovVafnASIIwi3xDpJfvlQZlMLOZSJp9rY7
8/dPyIIq+LA4dMQeT0EbMmRKywTEL7bfsbokNTKP/GdXTQaki5d6bK3fC74sECikFr9aUlXtfkK5
ghR4S3SE4EufTUFRh3ftKSvuLGwgIYeBqRlduDb5SoTPPl1XV78xhSrMt0wNEompUg5cNAiUjVvy
OlKmAsQJBhoaBWef4p1MKJanm1cUCcMDCFghcRtThZFxsWrMiT2lccitKOfILqOhKXaICURt0eYe
uFia5k8aElJtjEvPZCvPj3p8C2T+5JLSLpM+6Zt77MMKnL2D+OYJY0681JImPZ5ac6waD4uQhi4p
bnmJ9GBh6KidihLnS40dBUi2VhNyJnEtlYFVQ4icKEjSNkfKYtKI+0XbikaNTzWHQp1BvjpNDOtU
nzbEnwhsqqlhjIsecpOn9qPrjyN8Xb1Nu/9Bmj3nJ2+MtssCUzxsD88kmwu8g+9zydhiFzIrO/M2
MG0bgeSyQ5hD2pSlt0Q4OqwKWsmuF74/EqaZMecxvm65TTo4Y6qUJkEaGYVPuthTa8eRyoFQh2d+
nLuN53inE+wl2LU/j8ejgPB/VSe1B7I9l24jJrVjTOSpNcLT6V+yQ28HxoRTIhWb5+A24rQlHprn
qys0qse26fla6WDaXh3fsm4/ig9JI54oyy7APPmcN1Rs1DD9aLC07GhpXoaLfiLuMKSb1vpfRbWC
PwAs/Gg7muJXEfqXvvDnrE5OzGQJ/4GoLuZWUDFM7jIiQI9DQDtCEGuNS4aGoT4Jz6iq0dlpoIWq
LdFjqIiiBvGVwmyQV7H3fxoKIfQEH8GsjtaLSo/zwj9bMGUs7MAdsBuyp14wJRMV/C8o/+iN7fdJ
SPALh2gKx/8HvjfwvTEofcnKz/WXGLFtUgjCqqCjj+Do6G76hP+auy/XyvLZMIhoR7nYjG6n46ps
JPMibLYuuxXBz5ZNBStdozlZfzNUASaU/dZ74POFMgVbGCWU+bD5yN+GQHRftcIN61hlyPbV6no9
DkFb6oVfkxXD0KV9nvPRO7JqIKV5grbIAahRIVCKlxYIMIrL3MfAu1AjWfrpgGwXbaYHGQunR8J0
RvtD4P8iii1pRsO8gW6TPTOwm3uAxt/YH+tki6ogWPiMCuLre0b6eH+nyM3hzb7ZB/V5R7WLbbGa
Hy3IXMrNyF2xtP7mJ6MxsQ7c08lBmntb2y9+HNmXgPV0mwol31tIdiFF1/3Uv+EHkWIjrvyROLtw
3+hx/Yd32jIEhllo+Zbxn6c67unzRFq/Lyab+eZKa89wyKI1qMUYf+it9fXaKloFXk0VdEM/p7PZ
NCb3oRihUNilbF5UJ3vH3FRgiNXSa8VMfmvry4nz/pnE2NEK2d9MPBkJP8JcnyAeUlF6+3xzV7l/
rWKpb70muZblCZoZKvMjQjg0n6DtLGq1ehpSRnGhJMgpl5eN25iNdiUV7EqrkqHGw3LwEqoBDArB
HZlrpbTzrpfSNDx9yBors9K3i8Z3mv+LmXeoXUW+NPipd5fpSkXg6rtYaxhPShvHmLJrox4kTVfn
go8IF8ZniaQLuDXtEBXbzyb135etqDkRASGqVwkKRqGGWPWQMO30C2Z+IvbyvnShmD91YYF1UbRv
A7GhBhOlCMWxAGWEN8atI0eaurbgK+NNNUvoCjZKTahS2YU9cJqHh0txQLnC/a4vekZ4jQVzLjh3
bpNupLvfJW/ZQYWv+BgJLhFLIeRz8gihYdOI3YziFk40ev9JSzSXuBkgclUmafPc/LIW/kOtSjGL
yk7eOGC/zNWEfPkibSyEA+C0rBiKhWkbZ6bS+QCAINktEj+XS1RYSRDHESMN4VDJcBM3NknzSvM+
YrphQnQCmCSKh7FlgX+39EMPRSjoP14C/Pj6/bNlyY+NATMzm9EATiKL0/bOK2GMlG/BvHBlEPqc
u/nkyotTpQkkP3En2iS2cGGZ7BwYsOvTA2X4pfDhEXtVkBSlZrtReaD+GVEa/R+VWJ3PvK1VO9BD
sr5OzDe+j7/b6/JFADBSUpb+i3HmHsTqTzHo7awdfiTPEIUgeHfeEI/VehA47KJMBRCrJM525OjB
Xaf0FrPdrGlXgGMi0q+QghQ1oAnCr8hdzW8j+VSYLwbTeRlhSOhrIhR5t0p0MfzAoTHvXeYv8upE
aj7DhnOJW7f1ATfoSXKsJV9s5Ans3MqzeLe4nu6fS+XSNv/djWoVlTfv/CVXN0KBceyryY5kI6ax
2MTFGPt4F5DeA+hVDfBAnNqcNDnoIyROCrSOgn2b8vcTJY/BgGIDZVWrpJcv457Eyuit/iqszbo2
CHICsmO0R8QA0D8JEuSPzyJz0fEQ0uN94za8g9R6TT5mRjTgc48UKiRKCwm1w46J8XAxT9FYA/Pw
8XhysTg83MxToIR2EOSiPNzKNxXvjFaJP4UR2QRqk0qtNPQwyMl038cGh8LMAoLoFuU/3f1QswxP
5oCAYQW2CyIW17cGtO+136Z1EEP0ageNY+okIwcz8Jdk97KYAjKO07Dd/XvqGgvgK7CpLFryn5pa
pKMvksNKQaaOCcs5RAO8frf+VQ1pbnhpQ6YNKNaqvxIjR1cZDP977wwdwah7TZ6b4PkhkYCiIrVv
46gDs8h6DgLlEk0ndSxS7hVL01RFI/e7mVHWx1EuLU1+V/WZ+MG6+DMRjZA06u2Jb3iqiTY93ryE
mu3YRni4Yh8en3gH8ZThJA0Rk3jpv6aiXfSSPQ8aJNbV+klC0dC25jnsMjO5b9PeqxJWfdiZvH0V
brZD8F7GajYX/9yg4gPQrYAJqtVdtJMJiycpZCnAGtk0HSepfDOu/s/1kMNfMXJ0GvxzyLFk8B4F
c4M/rHdcGXy0zLGMjWJDs0w/+wUA36QEPFT4hibbe19Nw/cehikf0RORbMsovJkduaILMSfgH+BI
YG2UCQN+Rr9xY86PwRnbVE/lB/mmt8zmrlQjTZUN2JSm5UBaywbv2O4JwTNjZrQ0Ya9Le+e+dQGy
oBMyj+3Eem1YQx8nMbQKWZ8r8hCta+1K/rpVmAg2JtWCavsDHCyFTXdBGjmK733n4UtJIkUbbRQR
2cd0o3Z0Qeyuv9OWhQCUI3BhGeBkBGj2Snzxpfh0CdB9tnCzNLziB+jUNvVXYiDzGHtvzh270vTp
SCOZ95CQOHeNm2gk1M87gX4u7uZ7G8q87CKogcLlAuCzK47HQbT0cC0yZfRyUYbtNp0WHMXFdX2+
RVH7wqD9twKayS8DpA2yMoZmL6jmHWsVwiu9BQiQzsp1EVGTzWloRV5eJL+rGz6SJCnQw/ibiD1Q
4n0S3AcvMNWmbpDJuPpsgkLjsXlnjwjgw+EsSM7d48gRaN0n+M1xnLcWqBGEdomq1hB2uQfoz7o0
kLy5ysDqypq/SX7PzxRwFhhLcZFTM0budtLzeBLkr89Hti510QAlSVheMlxgipmokkD1DoHDmrax
U60BSc2GWKWk9wN2Jou+pfNc25eaTO/NZ997BWBWVg8kopwsDhgBlGY3h+6oHL5M7nMVzR2pi69T
R7JWhbv6nPAM0CQXYr5SkrhzPbKscbpn+VTOta3E6TtljEP0Cy+NJqw8/nT01I6p8XD0yNN+bpP1
6UVXOcDoSmGcoPn02Uv88/0FkmXOKw+X2bns8EFLqQh8E3D6YuhLYkvsDGdKXYxSvYVQGbfcQkqf
6UJT8a4f7oIIV3hIUCpEolE0I9q4emegyodljvbIhLH2SFZbCZWklA0KvXa9K93x1qQ9td3NSf35
6y0slsNHKuYGNpIXHlw6UEYeyU5dR2CWHBZ7d7J9rasQJFw6hqy3NGtcTMAcoJoJRtLBm+cTcslx
uZR/WkpmpXWcuUottLnSGkcVveS4JpC6ugiRrfnB+6OlIflB5UPj+DLOAK1TA3tu0MxIGd1qEUDr
ehUzMJsVcy0PLRmPL4xzf9I8GlDWrHcC0daG27jaYatbTg7VS+F51D0ReqxxipNda1sNpykXRJN0
69mUURuEUKrYDHJtFY69ABz9U9CThzTxgNYwGtvybopXifq8+LghMQvEjku4GMswqSSxMk0qEPu+
a00we5w+uCmMtx7sH0uHmMAIem8pzxeLchXQgs7JSjZE9fG21xX7YsgOvxA0uw7YaoKtdFehx4sb
qcxZcqFyiY0uR4Mp/f+FBh/5qSpywTfEFWKxKjXh2XwFFBB2msAEuGZEE4KXiEJmqQyUTpcgxBQt
a7Tm86BOaT/2BD6lWcoB4lSHljcFBoiVIimPHfwCPl2Ljq5TiGhY/l7G6vuYDVPjkosVvdq+xYBo
mRYQGyS/ykdqypRnyaTQdbrM//xLPDPYC3rihj+vc0dTdaec1tFS+KWi8ChA/5HIwm9l4EXKuENz
KnqfS1W7oC8dAKTlcPqYC1OHNA2dcjIQUBK69Mv83L9Su/YtFWpTdChKJuJRxIOcE8RH7sVAaaLu
j4SJ0BStHnQclmJ6fIsv1WtLnH1jq2QQmfI1Cr+eLdQweQO4vyjIHuDrdW45OA0A78M30+jPfYQM
BhtYJtqmUKPL/MkzZDfec3Xt1vJW3adAkn5z1dNSHWljCo1BEgWBnGPuLfuq6Z8YNbFjSgdoKTLo
W6PUzwDDvOdm4i7FPuvBa5QmxrzbP31czphKQZosq+HXnj8/03ZHysbD+jsaj8tRH1YZu3ZVNsUF
axasAiwe977cq2a0EI+oWPkJ550oDw/J88UTZ48G7Hq2eO2BpHWsy6DO7YhHY8yePIwDa+KxBo6i
bzyoeckCNsOV8N3FgWwSbMaoJXdGJcMhGWOEd96cGA/P7Q+hsi2iytooIsTbehSTWIH5ymLPmoCe
PS47OR5wb17BfIEZCHYdt5/6DGjJfWfBOU2xpEBGaEM9l/pGlwa6pC+2MuX2+xox1dGJ2iG+V3pO
aQGG9opqzJvaoaWQd6fksf67Nqi+iOv1aG+IlQ62P4yJQs8diDEZaqLxe2p40Tjwtm1QA1HZki8b
91G6eKSP4IWynJeYlH3xWnUVq3dMdeT7FDdWsvl6JjsfzsFmEQLPar5DzCEIgPAwBwHnEZSUWvaF
Wmqus7qQ4ws1XtSJG+Vjs/73Zm/MMhNCAvvh0z1+JycHglNM35QKWn+hCP0pFYHpJcSpGB43LA6I
faZ8reMNPR/s8dGS/rdRwn9f8f9Vd7oD0zjqkl4iC57NaEcxD3mBb8qaP6cy3BgafmfthUiNtqna
/621epzK1XrYapLjl7POgjqrUkdK9Ax0Aa1F5V3kPmHWrtKSCARBra6QuDadg0e9iHneZdjoECw/
3IcQf3asPLAXS8tDnSdlKFe4awnolX/uXG47vPFO/oimWvgFH17e68FUEm2v6xT8e5lD2HM84rSo
W/6drXilLc3wUngXcdd1fC7bUw9vzeXGhPATDwx3yH8Ahi0OL2gEdgxy3myBcHCAwE9qgg3edqel
+CByB38CnTA+tjbcxv3jdrnJmncz9rq5IEacR5w5tbU2XS+5ZMC16ZfIUWZHSDiUYnHN1a5jGzQz
XGPRC8nOTZZ1iqwEPLwDKlFO4aQJMMzeWfOwl9AbqWSHVtpooTImnjToiqRvfSWZJpwutqSTxn4s
qdBZHnNwYvvfnEQzvHqUK0X7MRqIBRYfQEyqeDDhWwXcVcYMShkbuXJiAa1tIGD8QHR9ls5z74l0
vyH02eKVUrHKeyLM6enJH4PRv9Mj1l2FI2TyM0pvLL1hMyPQjPL/KYbwmQqoKybZgyCyYRi5u3uP
J7yorFn/L8jtfnkpiyOKbZzCrhxY2scmfUHj6n1/MKKUsrY40hJ/X4S7sbVHketP5/+O9HBl/fp9
/xeR8HPKXUn74Z175d9ZKrtRbh81MwQ0FMnHocXeveMepO27dvFQIb/3msG+SR82nW4Bl4up6mjG
TCCcHvIyHvvbrVxNgsdweK8c7oTCPHf/uuD75OgKjPWTPsgfDOs3//ujhWw4bKZG75ssKy7rIBnN
AXGKWF6bk3wm4pM+mRGrIc4f4MNAO4VcayMnJ5gI0NDkvopw8UbF5C9jF+UfZnfrM4ca4VkV4x+4
KOj5F8D3qJnCT3rf709e2VvPfja0yp08j7OuERUOEe44Fr56SXR28rgv2xqUmuAo/B2wQDC9dA5J
TqQ4wtLYe7Hp3ZqrbYYkQ9tXiX1USqdqWdhbXZDvzm2ANt9mKlU2UUdgjWxwytxoWYRDnU2YJM57
3rCHjNXmZiat+w62QJgQAX8y0uQUNf6tPNb1RiyAtEhgqWLxtwV88ceckobaTrW6itigQueDwUeH
RVICzLmqkXMgbaP4isn6PsMQxqlt9JvagCTWTeqbfxgdHEylFIsAdLBl0TWEI3kuHq7YTQxAY4Jw
4IePNAz17iGFnom0cLhOZEx1bkOWEClA1cLuK+dlQTmiwB9ULmX5gHo27Qf5BgJ4RaUJwZK7gRx8
qXYgnql60TZZuWNnHIOpB2WSylYyZL1rnmLvOgYJwQcJHNdwtOpoQqQbqSFjYZW0Byo4DEGWZma8
qLFnJDarKKswiNUyYvn+/Fc/xFP0uRNN9CVj4yoOyUNZreVlBI+KcropCLQ/xsQkEjoKcjzWVZk3
8YKdBPPKmUETPQQxcyl99Bt2zFc8Q3VkttG18n8spYuoF8rBvCoJsZUZEe0pZ4xbS4xXcEB8zOTO
8+NL8ULdvSZuAdpU3lSdyposkem5rjbOAS/e1TJZPhPuqQeqAkna4G+c4sSscu2erLw8RCYmt0YD
8GZmonpohqpbQN276DTY7B/zNg1nJvkcw5bdqD6v5KxvfXMrNq+DkhlQvD1Curfopou/yIMF42GO
DWk2Qb6CdyVwhIAQb8lcnHM6gnkUGQYHb5WK0OqP0TCAJjj280iuTAC8k1u21ajdfvier/W8J1xQ
JCL66r7eQJPR4IPxHid5z96AAC2r/ULbFG6Lw1FyhjbknalIcQ2MbVHBD1bNPQP9kP//DheQ5+NE
ckm5+R1fy8hn7NumF5lwEm+2piZI06gD237SIz+1V5yOAvVv2JXII053BNr8qXPozPHs48IB65Mn
CG26+uWmQE2txLWJ2peMyqRUq22FfkdwMF0kdIHZyFTlnZOG7U6pDFAnZGR0t7iRC/Q0ZZc09bUS
fBAksD2lc1NLv/yEVkQHbgcrC66K1euYxDPcG18IPD1Vj0IzcVf6URY4jLBfDGptiRA7Y/50Xnfz
R/SPfNU4Dku4cWGTtw9UjbZ8K6oZvwUi5aEyEbZGdwEwEeQDj98GxdoMM/rFUCCqnuWQxHBw46Cg
Cjx5c4dlBZhHkWVBxB53M2IBLEeWXaL6CGGA51aXkTrapO01nuM1ptigjCk9QMmBw+Ik5BJCSRkP
IHjXURHZVczHGECrScw5kuAgTICFlIbyAXPQ8YmEwJctLtkyqLUCH1Zl4OqRxfXLErpAgYMU8qCF
+cHgKkYx8S/L52m605lfr5sbq1pnJN2EKCxW7RXcZOMpNqcu998T0jO6I+eSGRIZzTGJ3WzopsUV
Jb6xFdgry6HsMO49oWe+g7csgZhBGvcuNL5CifosNBU99xIWhAxxX2pqEhAqyq094U9nfozl0TwK
ZI8EwFA2xkBAxAvRZ91TPS/lcvJ9N4zUGzJQMNPPL10/gr83/nJ+mz2Wc5gIEDhkQ460Gzs4aWGM
Eym2Dpp6VJ/km3ZmjEMb4HQAGMntWJe1QgqJ0pLq2pCqE+cGAhyPik1njj2hBkzoj4YXWiWQcvI+
QbfxWF5ZPfkbT7RwtLFUtso/mk2WtE6bYl9sbTWSBBT4lLO2slWVSnk2WYs43wZ0BCh/BZgIewSJ
exeVU+YoBOj43ulQ9okjm40v3qQBQrkGceYQWRCk/vvkQD9A7o5EIXaSikj+MBHit47/WBFWMuRO
1a2lQCi5xUgK8+It+RPWkct1Hd5EiMsRZFOl6C4Rf2xAd7c/eCkRD8nk4uW5w+fXbXT1dMvuAzzo
efu6ePj5pUvNNdYOF8Zy0fAz5mxGtBwy6EFcy4UgiSngAC/RSWvMXkzBotewE2RsSaXv1ApHUlqE
QZqN/Q5MGbMo4QbnlLgu+CYSmCUiKEangos3KMBNBIy64lO7ZvywvpLI+d6hucp3JY+xor9EZs4U
qofoa+wLDJGxLENyWguotVIwGgih43Y9AvarGacU6tLPlrx/hIvgbstltrEg1WIzkWVbHSeiBkky
8hm9OsnRblLUjHnzrMTj35KozwQ59M2iWhWJAxtxTM79zvbTqBpp6GM/bpqNETQ3ObIoF+ga6MHf
S9S+WlUlFzjckQPJtCINmE3DQ70Xt8+1oY0i1Z7h5PJyPDqFUFFj4jeuQp949jQ4IF0ewTUicbXs
X55ulMUHOWavsMFh7amEraes254DZd2G3ssHuQ6Na5m/m7gOgJ4173EJ1owf5cx/mWL9APmJJll/
A3tqUNbyHC/55NTpdH9F55YjYz41w6h3zur6dVfo5Bgzt84llcHFQ45URIymWgZNyL7F0XwpVRAL
DbNkKlIt1xQnTtCd4lYxjwsWtbbEsM9eWzohrayB0zme+1oTFI/cj8ceXJsJmZR/QiyKs0RCaMeU
3tC/P6vKZ25LkX5GC7jVO3LZ2L4VbbxdhhaGXW2loRIpQuzpte686bvyuPG8Zh/kboMGIrCUAWZT
KaSUFje/+IkwFm4jFMLO8HuWhpK8v3gDYizNjNr7P3EaCJAiXXFi8y6vfwjKebrpRwTvPgzTjZpB
whUb4fIxAd80k8E61wKGxiO/FNwaPKJP+lcOjDwjQmcVXfNOy811cQ5fPFIuXOXpV9GU2T5YJXRI
5mDCdY55gB2OVT3mDxiqT0W/sSdru7oHNyld5DR++KfRBVLaqOTaQihzCo8ElVkAYWH8W7Pj8reu
6tUIyIkJCJ/3ARg6oFO5gWavK8wh8XMxogkGA90j1wjiPUtFjzHpDs+v1OtDmEitGoO8Mry/4xRm
yRsM7vD/oKIQuv8oW/bK1YZCILjc/pXcsQHAFnkN0Dwm2KHMsWLldKhOereCSZvKIXzg85u/q1Af
mF4J7cPF0MyyQZxruzxDKM8QBQRmtipxBDK45tD3F+LOxJZUbvEue3akrae9YbVEYTBtilbrTyRJ
ZvbPywcxtft4ntHxh/XasO9no7Uz9oXXlucU/0Ybka5m+5jSx/6Ne5RNC38FnZ5j3N4MSXqIObjL
qrJtdTdpBh7o3hIU7eTrl2vWBB4hQ+cg9HQ4plYGNhSQLin2NGBUz5Fa9B+dmecEDM6giVSZyiCM
sbF9OQ29O2VqV/LqWXot8ii2vGrRGcoGV2Pyg1WJIWK0xfaOU94n3PQsCDL5Pv6B65mrlqi9S30F
vJmIIzAe3+Wm7TnDp2wQVmkZxJcimHd1pUPn3ptH/TTPxvjQKhJXEX78zCjLQGXHWi0K4OM7VN1P
TPfhMDMnHYl4+kPY7fGZWUMjaQJPLX0nOkfdcamfn5zoBdu4bAJnOQj/Pp6XzMH/duPhPbM89pDT
rOce1djJySISFGwniilDhM4driTuedO6wmmCLYX4lZpD9Vv7b+SQXeXUlFBhnBy2ey9fWtDLCzGo
mFZBq+W7IjNJuN+c/j3lOlcY9xnb0EilMiy3pN5X2pJOyIgkIPVtB6e3nZmP8G9j2YVZwRNS8nQ5
Kz2NnnPZBJr9IXxqjJCAU3pTaUXDnPpn7uh+90ZO0ekhgu1t6Oe+OrrZc7Iq+nVEC6gOS49w5FVE
6UYZpsNEI+MZxw0E//jDq+L8k6B+kX2raG+qfdaity7BxNuaPJxh2Jq9jDVfAULtk6427HbC05br
Ulm91bGo7vc2ApV9JXLKGsMly5pj7m8cCT6d+xvCCHz5W6K4aJeLRNJ2FeHIuRoGyidP8g54Pk9K
iIAR5FHzDPyp6TIsEB+/NVLnl7QyxgRBniqnoNFwLJkzpDAjBkxDdQt8BIm6YVfAAzGoDdJ0z5fr
LGC3GHkIYcXAUyV/9I7k7bpzX2GslKZXAbY2TJggcL8x4iceCEiKVSCqsXvI2ZG0s4TRRFLyluIp
1FrWzh2Lxua8PljwOj2owe27RuUEmEhHkIETgfup+LJ+rvSl1dQmq3ZYhuVqAlwmzriPPJYYksW6
dGGZ3rVeWsg9WUuFv6cVuUnSjW8/R+sWeiO53z14/aGBPLZEgxnJQUSEIF1MYSt+gXVeRnzk7SDE
RwfwSVcxmzSfRI/iAFTeOsSgzokvKvifYwqswuBmrWNipy0CEN2XrVjUZ0u9+wH6Lm/Ylxvjxdet
F9wNZggTM3LSN7Ax6lvq8LIW0HKz4tfDOr8riZVvHM01w7zOoRdQ1uKrXGJx9MF2A3kcwEboS1RZ
8UUgIbuGdgCHZXfNUYo0mdrZXGzVICCFiz7WtKcLGsOAVoEKHSLcilo+bQCH0IrT0Pr4ilm4drkB
lmsqW+dNiJX8wk9HLt2FdURIPWB5IZftq28E2p6T5Vk1hm7KdWNDYE2JZPvkDTg1UQJQZzmylRR3
0Ldk+U302LGptaojDYsi+LGkEZszs/3oQ+fCcP5GRyvYJ6T5YF8R3s/gT8u8eIyBje8HgWMgsqhp
sh/LYX5sXdEbiZyEkNDCBMKOeuwKFItF9ANw42gHP4EkwPc2woXMStQaYuEAuksD6zO6xNE8Obqb
Tr19bTNx6KKNP+wKc5TlpXDkdFQ4N4IZgBFTCJi6TzjkH6PVwnv7l2C4PrXoRpkhDM0pb4Swe/7c
iU/wMh/XufcMeO7EOJegk4ZBeUb0qEf9CqrhHZT744IeNoNQWQFCqFiKQKRtOHwkFza9ZmFwyEcK
qx6bGYJtu6SvLY+aXfBsk4n+X4rbI54JcEYUx3dk228ise6y4BBG3I3Qen5AtcURjgybsdJAFqbN
rKYhQXbDppEkddgwpnLAVu53X9d9wsvnquXeB352EVMSrKawX41icU8Wf2p1s83eGlS55QOcUlIf
VCAZIjzSBMz0KIHsU+vNt6Z8pscuvx0eL+j/kVYNQcRAkQDbhzwRJBXm3ARYXZwuPG9/qexFJYj2
w10aJNpwufu/nA4a12jB7bC+7GwFG1l6GZhuoIWLh9KUGnyaO5TWtO9kfROUvicA3vAjxbLOmJkH
WbKYkO1O5s9JTeStYQuUJYwMNwbtQPov0zu61bK87nx89yjkMcBNPUeDEj/8EWJPczwj+e3bhMH3
0LSW8C/aR/gXYz0r+gbA9Zk/EciUB8sZj40neyT8YoAAQK5MSYrsFNlKqeBB2oMX1SE2uhnpXx1U
3HIXONDsvu2DknbPEhmsXhVY5JGiYMb2iG8GAhjezgWh9vNPBIQt/S7p7ofw+6u6gY7d8OMyxTHA
Nv5zrHC73WTdubb5I45rGunbJuq8iGp2lmJ2lQ5vr73gWi4MlsvXHwIgHGLmdzPJ4W72lslrK1U/
e14GuXeM+8yAb8i/3q8XZuseKcftODSt4fhlvW9YB6qKqDiNV9ZX07+Gfz0kf1ouF+JvFOZZYMjf
tPqpjC1XEuO3ge1XmIWMbbLkOloB2K18lsicbbWz1CGTrM5H0CmJ4eWPgHwrgWA4m1EYeI9ZNqpN
cpcJ2tjoy6b/UZGA+fwwuuZ0UbsQQdNzGBzbOfOhN1XUoz2rRHcEo9wOzkvYyOM8Bt5O7PdrNGFQ
L+vZCSAg+dxsYpmRvL1SUqu6IKi94Ra0otOD+s5m5S3bHFDQsFukbXs55gG2RZ9p1K3G3wtxNDVw
6zMGTezPr9pioZaj1jhV6BfW1zCInEbVFm7JEUS9K22ntU8bDFeVfHRw9CMlR05D84b9Jzz5eTp4
fb8CEjBwh5XuhJ6JkXHybWMbN9MQXviGz5AuyNYEYlxm7XhzdKmdh8Rv9uVqGhXWC1RNus8AMBmG
T69aJT5/DZsOr9WLVdUM9ArZlVu48O7NZWb1nvNKvxzpRVjLJ1onLpfrCksLqLFFnOBVRI8VescF
SYjKc44uouwVj5vkhd+BZCLOrmUSPPc+auAV9jwzRCjQfTT90HwRKvEYmvhVpEoUwZCdAmbwu3QU
gih2FlWjUYoMY4wSQsuvIt0do/+b6ZjndU1zx6KygCcs4TKdGASvU/Zgh0TGB6wpzULkLurW5r6L
yszFHCfCeqwRLsCdcQOQZhnfECBzopJuwwHuJS7c6EOIdTGA9DwEb7Yy3Zi5N/u5/Qh1AEgIQL9s
cKIX0JY7sWIUNNSe4qrfbpSKDXQqED4w0uEb4xlkrwAbEm7LnskTUrvnuWXV/v38ZIiwu2CsbNjg
N9VvB0TKlaT1sy7XXeV9My/knxmg0ppo7Tno3/YY0+e5Dx/br+Ot+wZG1yuYuITEwRLVgt2tk0bS
Mqdd0jEl/Q+AvnyxO2uZkTk6EWLICXSJe2exIAIv9LNPCzyIcHbmLMjBynbqZeyP5qTnAHJoPYxo
gZ8Z80iMhvemVbkH2NBbRf714kCKuwvYg5RWOQlns4ro4wsOvEjKmFl/+l4ye137VOGv4z32uqEk
I0xKqMv7npvv6TVyQvhD4StRB+tpGPMpctyYodfv34dVNFJBF2RpESH1ucbSJtgSOdiHWNLStxv8
MAtlr75KKHwi6hcPuBbu1v34QAz1y0i13m+kgjZhqGQLOuA6OArLjgi+iTmCnssKlU2AE39HvGNr
5bxgGWJLqXSD1Qw4GNgMJpR4GeioysFvQHoYchvtRB7Re8zyCYdPHGbMsH03aYVIZouhI6ayDKVa
e6x+r4i0FTpuwB/LqEyN8Nr/n8bD9O9DMVkKyDF+28y0Ta90U82+a6ILKKX9QwfAsQHepG1zuxlW
+FmgSkl8q9r+oMBLYwWFu0EpuTKHn5/bHFbgJIxzKMT0prYWwQUWhga8WRR74rraGd00Zlrdmn3+
MqSwqIPyK/Z096qfckySZIW/BTXnpz19wRf5ghEtM9PifZM2sAWkTCcWirkp8+1NqdUMn3WET4U1
uojojp36ffY88X28vzd/653IC33niFusKucjUyz3C0cxJix0wAb3Dz4pRpfZHavtDwAWMo7fWPA2
xiwlx09a0K2EjFLjHJqy2cojXEZfHqvDmndPe7kpWHVOkZ5Sbq70LNUjfKRsDfbN6uN4qr+/DQJ/
ISF9A99kqut7etmmUkJVXjnjL9b1EysfY5BWCRX8wVpcI+6G6iKpZi95Z5c+SOMnZXNB4RGxDGX/
bKrcqINcGEm27MfbXegwP7b/th2Jp9w0LsrMRCt6aMMY6L42l7bhplwJHoeY1qLscy3pnRGYWaJX
mAL8VkkrcEVP/LCeQEXGXrYaK94yRh8qlT2NRjAHVM3tnTIwHDrFcbsy/9Iz4nf+VSagA96vyB87
ijpU/muRLveJYUUnXiIeYmFKAarT1C62NSXwWjVIqeVwSD1/licFheCIxFwP+38VvCsy3RiGZxv7
KyXjrn8U+7AjkfD4byCY0BI3du01K1jvG7uDrmt2grgP1YXX6Pq99C2ljwkr4aCc6kvnyvoDdApv
HEgIIP+1N4ApX3PYX9tQzRuH/n9J2kB3TrFw+smEnz3pPFl796ik6Pt83+ySzBn+G1EhqZrR52pe
n5Mn7U7uLgCsVdrDWNkwjyiX+8DwheV5Y6nisNC4BqDLxRu9GbUmi6ZwVVCPQ6mkIgCxGsbi3Wrg
/CnR1bPmK1ToCB6Qdca8fsriINYXmkqs3xfZjFRtZReQ/qK3+O7ZDSNxXitjjhZO32awRUAkKoxj
soHzyYtqYK6zP3+L3Ga3NcuEBX8LZ3pIHB0B8K14Y2l2vZ1dionl7rh7sKij2+m7riOFJNTyP43o
xr2vGwHozeneqbuilj1NgWmst1eAYN4WfDyFItIeCiAEaKLYYLdV+ZDUAg6SAGT4lAh9N4OlKl38
0ES3zbR6877E/Pyf/SsFmEjXXWCj0V9QyDR3LBYHcC21J1P2xlxuiGREVGavUQgX49EPqKITPj8R
AEasgYkf0csBxIZw3DppDpJ8Wob+IO6kjSXa14J9LPrafculCLwbqB3uVr6mwKESTzNXFPc9ePH1
QzxdAHFivN1IKOaGEfkvWmJCmSWqTd4dJxS56cv8vXBIXoCqO18cW6KSmdgc/dBCwHMX8Z4rh/hF
3qmt1Ap93P0Vx11X6yd4r0VCePXMZPCbkBEaOGROM22tU3DPni6XCv2In/AqL04bX3HfbmmfXfLl
pZSLa7Yznl2kGIkPUi+NkL2vARID3AHyAaFi4/nEHVM7HPa+PYiojXtfWW0dppjcjn9Gl9Q2cj17
qBayZPzMqfBD+MAtzXYuPDXrNBpSNv7I+6LSNLeQnsm/I1HiQAhIvDy2EslmkLFDhtVKkuIDhseo
a6z7icTul7mZM3VV8LODIAZIesvySlqIZxKIa3b6wLpNbAuWS+tAXm6Q55BMUs7FP2CvQ+9mplSk
fxq31UM73wBue9nepBy2S/8XynXudI6sOmGbl+csCtO8hpPHAWspOOVSSidmMDYeQ0YELisfWmI1
G/mykXTVGULmnoQ8F63j8zkrveWoRoXDZMM2SxyBRPhAKkSPYDhTdW0SZc9w1D9LeY7OiDgNITiF
wRVWKT2MH9oair8p6Nt8IXCmFATuqlcz5JuIJx8RhtV+UckltrFFl+JINUMrL4O7M/IfYg+OdhrB
6juUdIySKrMcsKmH9J174FruRU+UZ/POwIVBLc5URkoJEIUzA520nyzYKqWJvKqixYor5BleXmnw
6Ca4hTg6xzisMIOkkSBK3sCJUUVhFVnGLw/EMLBx7BC7DA1Y6RAP9T0kA8STxCGUpp1LxgmNZoxN
pOfJ8C5lNmMP5Z65dZOkS95rxaq0A+YtIinvYeCqQUQAsXBxuBQYOWvi4upknZcdNF2RBQd7rjle
ECGlcACLa50/rVdkAgPpXQl+BaNjBAOGA9Yp4vV/Txqa31nkLZCYksFMCH18LcL6w8nxAgr/Pwoq
Y8uul5yNdWdEROd/DaXE90g8WVON0lCEcV4w9hIIUxzP8iW0Bw8LR70owjICmso3YM9V5A0YCP1e
iWVGL5kluigx3iivsUtyDmQD1pFADaSPGMOeJeXfxOilyO9YnIikHPZG+srVP2yZkjmxuuSczU6M
Zhh387TruuxzBJklCQE1/Tm09OSUNS7tHLe4eguHUh4iSuDM+oA0kgKkxZkcuXeI75uQrUcNcqtI
EPaN/p5vAyyUmJfmh3Injyr7YD8y0KcvZ5CQclab98liwxCzD4FfdAKr/jCEjQz38YG+t/LUYEzQ
L3hYd6pA+e75xhok0zjd8VexEmfiI3zlTHvyAyEWm65+29+Ot/IBmCTD+hJV3zJwZntveivBpfVo
n5lB5mNmr7dvOYhSzw5WazDZJLMWM3VyY6tODsVKQHtF8EOAXY9edQu99UVRSPmwx+j0HhnN2+nB
Z/T3A729twBWkNdGQCbNKEJvlqaHUVdMl6qBzBDuMCF1f1fzwbrGkCgiYhjppKHaYRHBrdiqjKlN
Jb6GAn7uFapud7eCWl3HIjNbCSFnBTX54BUAMuV15h2mq8tq0SEwvk6HNTA/mYxwsPqTLDHbsoIs
ws7wBZ2nDO2ySMXBjSKPTroq9NQbjSKJM3b0e08TCV/UKBZqD0emUTGWg18gUSQjQnwbY+a3TLlG
UdCpGdDOWHOwAG32DGANhQsYuCQoz2eFISO0klvieEq4qY/4HTLFjnsjVOjN/cgldJhRybuYpeAI
ocHHv8Cl8Eljwe/nYY02Uciz66TiuV4h/f7ZhCCTO+sQ7HYxZC5d44RXhRsazPmPoXERm6KVdUVF
xI7bQMTJf6a6h/IB/lLQpjsezPuXTtrm1jtyT72BGJTomJbTmLrl/ipYthtXbXGOnIz0JLesKV6w
Oob0DjGV4qkYJhIeJO68WBH/hT0dgmCTENYxunnPEAnbtyuI+cReDKDc74uAudAP9fWdsAFlgogT
lziqmPFqns7CzWkUjm9SCIZ+hsJC/WU1+q4W/8WmwroaFHqY5z81+ybnkZyw3stbIE1qC5tSuIWt
vzBxDJUE9J3dvlMUckjwUlL60KGKP9p4FhnZdagzKFaPdI0ktHhZFTQqI5p9SkWtUKrPUH1pO0xI
NlNSPvX6M+9zfWLoMd1/T4stEo56ApqssuJ6Yepcy9GyYAPLnZOMU5QANFS2Qmzp5mHfow8M4gzu
PuVDIbrZpUpqBETg9YGaY++a9iYjO0mRGsBrzaz7Nho/PRm3bKJcn6LlvYaHboFNRRzc1ePbkHj8
mDtgbaUC3kGLhm7KrOmPnm4umfpseQTYEb0Ki68C++SQddjefJrVU51vsxz7wQFV6oBahJf54kdL
jypoVSa9BezIJNAagiGYv2nqWc7kDbFaee1BDuJazeU6OQhjvWXTLCjm9sZzLyClQtsUrleWXedy
+QY2D/FWC4bB7OuWoqOrDsOXiVReUrNBEwIVY+BWwe9ZVFsLBZHKwhtI72cc8f97/RB3+xNa6obl
YmC7D+wj2PlTxUcLDhjdhdBk1CyPJHdy8EONUlPso7vbxLch1j3MJT0I2MVN/+qU65yrIatUJzeb
1LYyU3YxIU0SmgaxsB9BX6ZxV0TsLCwxUKxnOB29lHu+13slb8gBR5gzxvASsoR3szrBkH9UTyLm
4L470Wnc4/QxIHut55gzhcnWXGj4cN0qn5yCvxWTNChdGt4yl5DoEMjp7+pU8KOTqcakzNGQx4Ym
NrHi1QrobTrTKLYqjXvmfCJfnKxVYiRTep6A4QVQlMo6oz/WS1mVdp0QmvNhexRtx7ZA8kN3R7y6
VACoX9SFJCMwM1tiyicAqWLdbqxX+uCNeV9Jx0a9+uyABbIGno6Ii7zEFjtNfUVIabhnHfKWlTtY
AishJ99NAB7UFQ9dtx2ccSliwamDNiGz0lh5OAeZosq6/2ba5bZTUw+/suYgysr23f6mi/ExyMfR
RIToJa8t0J8WKd1Gk+9B06YbYOc8Dmp+b861zBlxzSMnqHys5jZIcL52IwBhQA/qw/ydyVBxW4Zg
KsVK93fhiOPqoLe1N856pfaQqzvwYu/0LCjKo89LRQJGm16qCAjtAXvH+DbGaUNzn2QScixRqV/h
XvTWdVNFovnxDlkxQTQgqq4qphO+4V3nOiXlUcI8SoFyqSTXb4xS1IRZxy+lw7Gh4J2z01xnAwG0
g3yA01mQrK2+Z8fSotvLbPYILTtX4LHjy9A3KykWOJnsKVlYe/k+MIEuS/QabY7ydTx2LS2KYqEB
QzZPFKV9iFDLDkZoQ6Ts+OfpZ6jcyz590QP75Bpx2EeFgUSGG4mEIhwa0YZwgQEeGQerw+W3FIMd
Ak9d7ZJ7YUxI7/2qZplxezyieYGRdX7Jll+wU1UGC5rMNZu/7Ny93FNPi9y3gt9c8kSWgv9tdd7K
/P+/weYX0CXX/s+t9zIldbeHfJoaV48DRtt/HHxBoIvNDhtyGRgeXSE+pQ/FZNO+muq4siqL/m6c
QFQ4HR76ntbtgHbWziwbEuWqe43heYxBijWaDmBqdBkpDg0mJh8OGpD72+0n0ktFH0uP1Hpi7dnd
mhu2peKrkdGZwMtuebEnvBLtqVVXrZefZLPjsT4c+LSuSHR1lTVOkIxhFP2uEET5eOhYqlpxWN/Y
iGzRv7gWjZHV9/NWNevH6GS2ZVcCpvqbAKWF9QA+UDPooEio02B2fw3CY8AY8LqlPztdCgZs95JO
Bh+X8oo+NoHWNeySVocZPa5Gdg/l9c4rcMD5WnITt95lk5QV40LdZ/dPUJMtRtxVWFUwMGkIMxpZ
oLCPqgkZXQfAwDmUixig/Ahy6FTCvWBbq+pAsGdcyxfRpoVh3HbsT3B4x8R1Djx0/rSbYldfQPTV
TuVhQaJtvOEh7Rz5bNkf6pqWB3UBy2U6wL8DJqkC7Gx7fUNZXBVsFjHmy7MkO1G4lbLd0opATDSM
SMNWT7bxzlaaGwNYf/HezFOz1xn8qShjEd9pSH2ktKbzHcNZBC2Xtepj9UL7NvFg+c8eDK0dn5D1
f3rCBxG1EjCfYmzlHmq1SwPgMEvvpUh4OiuzDxD+05QzNn3q0aoMS6PBS/ijiVFFOrRTlhBIMv2s
MFV23VPomE3HXKwbTFy+9+dG1OSoC/wQnrYWe+69uXCWABA8il6tFrcednH1XIxxXjIXg1Kou0B8
B3EqDMNst7UHg32K6ltpoRhNi0cgeQW52RZSLsUslsaccx67izohpO52miaIDvm8HlIgHs3EHxYk
ZTfjASQmCTNwLihwC2YZLTTf0FRbrII+4yg3L6DbPecvz1kprMCcgRzVda7HpXcpdoxIcBl7ELWb
sjVPQC9fSHeMk98mhqnAYDyRRvUbpfzaNhIzJTkWbHbI1qSPhzwt6WIa60VVP3TKLVc8Dt4I+S9N
oij9NUNzaD3uh6MnFpOttTQ9jQpXoO0rq/Boy62xgxkKylbEz1eofO5RSUte8cJLKvHkfCOGdUxf
2hLZX5MosSVZVEHdnjURGGrp/fsfOVB3ltM37OcAcxKbd/Dgz+EaUWT5jO0R527hpcUrakZKhYPv
DgmnkfLYvGEnuER0WLxb7ttZx8BYLpLvdbw0nvktXAVwXb8+f0si0cx0TX4HoAhHcX10xSsgi7iw
jqxu0VSIT2Mh0nDmzYCR723bRcrvjgnsYMkPi1co7nijGKp/NgS+t4saYqzDK9RKORXJTZgsGbof
/E+f4AHCDMrBcJgUnTRt9zprsHV9ydlVrhHR/iTgi1jBTuHkDXlTfQNAiLEgwH116EteDZokbhAN
eZxVeDR9rPOunJ1coVSZGiq3EuqmUJ/kT+dSy+0q0adFT9PtPOv02gUY9VFOgIWpNAD29z1gmOjK
G2uRsB2Qk+yAOmkismb5OrnNoxJKmEV3/KDcviPZmApiDP/m8jloUN2m8jth6Er9x5/pWeJDWVTt
o/pNjD26vDrAKUIYAlb97DP+7KJG7tbhRIDT2iDW460ggvSguVh0vF+MNet44hfu2HXlZaNq6ew9
ta3CbqFRvLKE8paGvZHL0LoGDAFpIz92UFGdB01Wwv1GmnvDuQVCo4oW2Fl0p8ZFzlwnnfGKauIs
RkIxozJm3blEc9dj7nqzpFHaFz4u2+DI1f5mJNK7BtUqcMAmQVc2L8FgPAlhuUrsu7gl0CBx23KD
RJmqfzRKHXlMnECCgTyd0aBp2zC9eZ1D7g/yyrcU3wL3OQ+W666d+gF2+BweX1yDAX+2f+o0OiO1
/Pwu+mhDOgC4/KtC1ZA4WklaGa0Ecv4IEJQtJi+hOHM8OBir7EdMO4/lbVdfyasZVxLVJHE1Yczi
BmV5Vpu1RnVav8r9/b4cYcYhMQ7jDR8pZ2tg9jkYV3c/SCTTUxFnVgKFyQ3KqUfvfwlI2RyPUgk/
aJqVbk5IKfCZ2mCZzKHejYwh42NjGnRTlBFhTUGcS6YiXlBbleQeCkMyDlOodBBC1gEnjbEWekG3
Zh85ooAr3/11NS1A7gQphd47ONKS2wdpgz/eIAoBXQilC0MPKywkZhXOhrUczYep/SuF9iT0l07b
hO5iMty5pT6f8R8eRWP+wdFGrHqC/cEy2G1w+NRwD0Ry6Bizt+kAV9ASq4Mr2GSHPTZrlfjkuviH
P6jd9BI1od54/ZbMg51hBAjgjrL+YiJ67AXSLpvKdrBr8mPivWSY6s+suQB3pWQEyhl4l/2CdG+b
yUwLEy42uOsbOkANt20vtAIyRcnwy4UU5/jSuBhXT02i4G/uWLjPMRjSaVSQ3m4SvHpO/efRox9o
qnYIbk5rQiuKF6gysShDj3PmXadp3lDesp9NeZ7ekMWqsRymtAOdR5OTG4q2U6EK0KpVaK/4Ja4Q
7LTp27YiLjCQT15kySsFwgRrTVMdTEwgSRRu1JPCO6t6vSetmaMYLVtzVx2fwmg2e3/J5Bf25UvQ
Z7CR2t9UEXV0unXK5zEv4UIG5JvD+w8L8JpEa+XzDfIfKHoJddS309onUcHEYNjQx4GmbMeoqaso
uOhbYm76LQ7avl4GQHY2HUenO3beL8gh/NqNcuu6c/qhinfSzMhv0OctnSnFhSSViHB163HzR3ss
hEDOfG0wHCyzSh4JOlkXskhX7ujucxLS2y3VjpapO4DTkchAQx0XU3x2APwliVhrh+tM0PI3eh5w
ug5BwogNh3RjOLEEPN7z9KPeHH+SOu7pJsTZsqeQ9/RAPyReY9mWrsOmPvTdvQdWM/ToWbdeklhA
kZuhivAKU2y3kbSiDOikd7TzqmhHoJbIfMJRGrok19USoA5CbSIvn3PHFyWREI/oLlnXYZBGfVMT
OlbmExPe7GVRKRyNpz1U8WWNAKQxfN9gIqWIKixlqP66TdM9IlfdI0iDizZJPfzHHuI2KP5mGdgy
vEkeJljMP+NveHqnWWcLr3f9958QLwJMUJYmMdqKsPquEGelO+nC1nIPIYBIEXrE3m8e13V4rZYz
5BgZwCs8KaaNTvuGyDVf6jy9sDtrCbI6GOpNhCFBbCKDkA518maxcJnFml/Qz1KdpifjS4ConHiV
aL2oVRWR6i0pY4IbXq3tOe1rR9ESTjRPJugVLrCLqVIgT0Yvp0kw4M/4I2sTIv321YIJWT152LvB
QA6SLls30bfsSO7EuQqzXGotv3bZRdz5Brt9zonk0dTimIC08eL2WF2p4M/jUnl1sk6W0aoRbziy
fXPmOaJTNUtgeugacsqrRPIlST/itEzG4glyy5clwT46Ix2fayEulwDrqCjFghwcoIia9wbP7778
H4UaoOHufkIgdvn0hyzTPGseQ6LWtGT57FSEEp4stDUs2yQ5UsU0qB99tOCFrzNXcrv1RiPL/Fxn
w5Hzr2kGK68CFmBHxFhYe2t8EO22hhsPjcfsxjse52G0VS3rnfDUDfr0aMSA7o8axvsV9HpTwqyC
gn30cq7fvfgSnnVvRd6piiLFHrUiVYsbLxshvGwRIsqXFgVI3eL+Xm7OaPRAJTbnWqa2+7abfZVD
h80zZBHtIQ6Hbo25mvOkOe/3MBoD5NAEUWS6+um9E+QodbKIeTY8ntXsu0rTUiIUMHqNGnfrwFdo
A0vnmHnNYKbYmBzCzzUZcJOmc5Dz/SXX94pKAPBjdrW+M1As1WM/15lggsK0C1nLaKs4mkcdfv70
KvFsASVwKMoNHB/+oCpm4ge6kATsgQaJlh5X7MMmKtNL+1xMSd3/lx2cyUhME+zZmuYuTiEyQ8+9
b4QFqcBO8A9uqZHOOhcMYnHRQgpQr4jploexZOt23gtNrD0SEhcUEZZOVpHHQX3KE4DYv3anzjBl
ol8HbWOZn0TLM7p75IHVlgFQM4vsevCjNlSAbhQOTGPEDHmd3xhot9wVYVmBr/yYaTOEKiSXuCTA
kwLuT2sCyvjaPI2AMOKF5kXRaS/TrHLuT0YcagHPLAxoJAm4XaAVGrR4jzXgjGTmHk8HLElPe2h5
JmZGYLI3B8tJ5VbX+CGKFlrIiZw1++lLoNL37e0vwnQZ8SgExb5zYKqckHmSp6RilwdRscwLSxNC
GfFr3HHPqKGvBIJPDhgFZp2MK2tUTjq2Bgqu54ov5YnSOiNKBpdnMPXlh8sMzPPtc1jBLiXoKkQi
mASVsi9pJIGsvTPPAaXQLkMlVHP31OixazESzladwY+RxuqKL44xr5/Hg6DCiqoI0M5TkwdW/0is
jwGvRA0p1iu5G8DGIr8xaG/Ke8oHjPX/3voqKG9q8UtTv9bxyBqw6elqUS3PuUsw5jZ/3GHjOQ3w
3fzh1leClN/Y4GY9YVcMm+k0lThlQXHe2MQcmD7umQz6zZUW7t5j80ilNFDunGDLBBZvnPCwQ8Ku
TmgOTnfudF1G3NfdCwdWDof/T+GuFEY/etOWXq4cfIcM8tVVpwhE8PeTJQmTlHOvJbuUHNhFBRl8
CkwLwDviXbLwzBU8vKCC2CeIzYgIwhI1PxhJsD1UF4MQ8usXhUdudHhnfHdZADCxO5kSENYf+rvj
LJxO7pMLRtsChFcvyE7kkNI8aRppWMYVY2pW3oQGIsjv43+s7BwX6/zOPbyYrSzbpKsnAAup6Vp+
nVxG/5kRreWHkYKz+p6J3v8oh7cNTXhWgo2MDcpPEC2FbD9930GqIip0CL5cHUCZTQBKOgNkJCS8
flj9gu7ohxi6cbBvkLW6T3qSe2i2IMTAgYYmBM9IqzDykvLfcRk5SeHIuKIGw1Eq5wETlPysggwj
XVhsr8Sl8609MMG+R+3DpcpSNX6xTuAglG1BJl/kh3wMnPs3pvOiBJvZUOy0oHALC0v2pCgfqNcS
tyPw8pdpgJoP2Ovmbm2dJ1ZO0Yabw+OWHHuZdw/UMU5FpiDiMmM5gRrakPwhbMVsIrXAMKAbFl62
Z/SEqTFkT6H3iW3K0qu1xWIL+0tbW8tozYEtWPEuIH4ha/+2VKg7c8WR22MGSR5+TYgST7pX9eOn
q4ZkCfUj0oDteR/ExMapUrHP5I6Pw/iC0ptnag45tAyYf8kXSP2qjSCLbg81j8u9s2qEbwlYin9e
6kwH1soidqA5BCJZt80JVE2zLwAMRsjqavKhudZgeaj4LQHYI0HsO+2UUN1mWbj30UlbChwbKJzh
hs262cr5DOA2i099Apd08QC75B4xxe0CtOSjm3IG0gOS48eZXliQjOdjBCOxtNdNLYWJ990SrQYU
l+BVga/PuU60L0esodzHGblQ5l1smkgU1FZwcXb9MVQvO7DDUX0Iq+KjHuZMILtGK7hbNhit/3/x
9JfJe4wz+DxyR8XFq6YUQhN8FlXH+/s8BpFdz5qWdlwVkwYckyfVeT0PFauimbPtrzM3xkGAFWyU
p5USYUKaXplDmEEHjEZ/CxPX6RdqcIsZ2ac62BQgiwlKGT/JZAypKoerWSpBBk8oSPpZgt97A1jx
gprxeEREWt0GMz/FPTzT3ucSr7/R6qWUMarVL3hdNSvDJMV43tPA4A7oB9TRcFkNQBZT/MBJ1Bzd
hCjbiG4wd41hnkxc1bIG22G6SdokaSrB+ATQjc/GpE/zEdwWvC06lSJ8XvtjOqEfM4gh023kSHGc
bWbFkCmrrkBzHhTpvaDR2HqLaOhjYRgkT9iJuRzH/G5b4EHkiQwP3O/S9QrmBE0YHc3pOxpXkytM
opXy1kSCoOCiRfkd31AhdEwzr0o6LQYwWpdgntkYLpXmXPw2gZfmME+1YbT5wBFwsV779/YiI851
cd9xqIoP3fckX3heLQ3t/04YdfOGn5wKB4TwDCZPkvd2haTQxnszRNM7g/kk4ggWxJQ78KUCTxnX
CRBDyC6wuve60LO9hiSFqV1ReSjdvBKpc3b/iKPsCkwiN5jgZqV74TgwY2GXhawfAKr+IcgYOCZR
izTH9JTkJex9RKgFGCbenpPeAIXpY2eZ54z2ajqRPQ5OSmEM90kpfXb+eS/+tBQX25VgWk+d+O4o
48xPRfi84CK0yzYTruV4v+bv8DHv7LuirTeMg+hXBnrCyKkN+pyJkd+tHW851cmof6WqLZRFrxZj
eXeNUbhKTR64llYyS6espUuo7gmt3olnZMWySjycUxhp5myKD3CJa3s3nmzM+juAbMCqe8Qd8wab
oI528319SfFiAPQEHstxoEo2TQvKEBPnqIkCtLet86zAB0cZknqRha8QtSBoGZw4/PX5GVjAGG2h
zRK6XPc3mcV2Pgys+1jiANagaKDiccIiSMJrpLndy6/gVcwkLMKampIzoOF+xIu4sMH1pigfeAQe
Tc4e2oJX5NYilmoJpmv89fa/0Ficgmgo1kqxdYS0vQbrNOqB8FmZCUMW7kHO1+/UZP13ic/Ux+QX
S4P0yPSN8y2DjdO+h8IoD+S1BZmPMKwYNh81Ftjz+EPTezR3YJdMWsnboJFYyQxptnR6SAjvRGqW
dMK/TmcEg0lpOC78mVwVc4qBCDvMIpy6PS52vILoZQ4MtKGHnrC8CiZLODfbCPzYw/8VWuCAKeVE
cCcvtybRr3NlaxuY+GxlgQ9dGoyLH9fnE3QiWqIK1wqPa7stLTcZuK+MEb524L0sJ5nZL/QQy1kx
UYslJq9kSgUsxmd2sVFsZAGy/dMt65j+NtazErJKaBk8IId1fTJYejzmk0+xYI4FNFpfhJ+ry54v
upRh0mQI1tQBLnk8jwF+9/b11e4LsuzJjchEESqCUBA09ePAdbpB6c89hFMml3gyZ4PDn3ZnVrdD
yQqcbcjtcqUslbRtUlPHtYPm/Aggbna1j4G7Crr+NJoB+OQuPlDypx28PugQlON5GVRkgmUwjxa5
MvvfEV13LGJHaJTnMlYlIrPi3djvf6EmLzI8PqOM5hdQ/4ykTrl3OBGc1oqzh/PBK2iM4e73mGrL
HPMOcqVk2B3WjVTnxrlGVsIOxJT2hfTt/4bV14NmFGrGO00uCCiBUsuFtAZeqcuhPgkFe6Cqsk3g
VfBQ7I8Hq2s8VsBCpMjdkvxV/iw8TX1dGFjJpu9B7bLk+4BDMAMBP8wpIf/HYDAZhcqLAClZ3Y1p
yeUVXgRaVRT9KF0Lcek/gjH/OnVNVbTUJ1URtk6vTZADqrqJg8zVI6NpMmhd6B6UZiErTO55WLyG
TVoD+RZqqEf+Xl2LcYQtQGzUaEX4ilja6c8WljN1NNghpmon4HdCmJVAYj0x2Ga++g45xK8TPDsR
DSwERf4DqwGUdPv3FYZhMrKQqkTGBc37JFQtcdgA59OGWmzSZdit39lzBOd5ZJ6HvWuvvaPn8q/c
ejjK+pSSZ3I/wstIct7/cHGF4rWKW467OQh/5ot2DxhaRLYe/+5ve/5CGLbB69rTr3UHb+PAcIic
lXbD5Z8LQgYeQ5X1Y1SI29Un98hQdkpG5i+zavcjgP16mLx/flQRmk4Rp6J+2nzRUODSYQv1w7Xk
uU3r2ITy39Sd+28BCz00xpmk1Vnjx+zVpBXgsF4c6EwRwJ/NR2TEk++5d/IpUm3+msKhiKasRgPj
/qqF+Pay+GLhgDxS1/g/hnLvStHoMqaqD6s5duJWR/zLxo7rHdqki0Btcvbg8fhIpvurYdTzKrx0
+TUI/ZW1OJAZFenL0iMjqneW78ROboNCT2ogcwatTzjdOXPZxucRc3kxSB+4k/pEqrknoFaYlSVz
HVE3liEQ6uyCmb8vW0KSOdaa4nxKoBiMWTBImVSMHbTSEhIATe+3onJLk/i9j3J3Ibq9vxZbmmue
UNOTl9iJBZlInI+aCGqHCv1lsKoxeX+okzsNbcUZlayPbPqQ5hjVvexCnVpXOBFyugKV0agJ4BM1
ifroew6CsTeR2KWQC2zUvXaEduMjYFzKL2Q+a8Vy14gJfVczQJCQeuHLYi7fdB1WgqRMhm2ZHexd
VBvrZ3TRZxsdZFvInc6H0mb3T6f+370Mlt4s3Rh6EeAZhB076lSZewUgJ+hJCSgC+j+mWWXYNG1I
JcoLKiEw+NqnLz3esrQYa/018NdpiY/WvmyHXIFckeA845msOXu3Gl6HLuAESWGbqymLwb5YIWV/
xX9VKGAWHhxccZLhf3PlRrUT1KzK6GJvKW6BXL+zkUMMUmyaxSi7vTmQDde9BD0h6uotXBEJvFJ/
klscuXd3vDqvC4bxJh/MQzmDOb8jozL1y1mVGwuxvTrfTBY9TLcD6QW+t7eL9JjdhOPqBYSPkifQ
NNHoCfOZjVrVlXrS1r41fWiNdRmqFCyhrdT16lOvcmq88zkgKfHXwqLRYC+l5XaZ5Gxo1lLC/AF7
saHP54RVeZMWJtTkDosGKiP7AWQe3MJCbB2k48sFc3cH4wpYUcT4mqoWqQ4XusJPHzc3p1oTe2em
lMlFtcY5OEcneqLSFNi3NLn5SjyPRJV9ENmumX//uSomhXFljgy6cEUDXyZ2dztZJrJQARI5YGLS
P2dIyvgc+0QYx3/ytjpFs9KvN2WMwDCZVjkTWcoUz+wjSkUxi5jNfwmLwQGWujIeEbl5KuFog/vZ
Bc8Jw87IOxqUI6bkIFVNiiX5m9lbR/hsCh8sxnPTdA/3f//egUgjIzYLvMUw14PnztZ0E1Yp6iq8
I3U1aYZkHH8K+LCDqXoLrsVgwIeHhI/jch7kVfI1oZm/ON6Zs5uHa6cL19pF1lp/gqYjSM7P6f54
V1kM2ezCthg9TJmFLc0Vuk6zDdDjXXnhvMog73egjFIhGVHeFAPlJXYEidps2+b5Vj0Y8mAgUm7+
bdjGA2j1HZO+d66UJzakM8GUw91qOOPsgC1JYWwLdfCQaBRH0LoXL9A2BaslofSLHWy8Vdz9a9Bh
TAsTeUZKrdtd9d7EZeyjFaqj+9ezjY3vTkEWZz8FAFlz40BNPj3MvlyB+JZBdXc4Z3KyWzpqMokm
eAaCGOnsR4Per9FdoD97AggHeqOswNzmlAJVI1eUuKU4/S9y5jpcxtkj7pUcMeSP/fClsx1Deytt
Fgk3GVVmgMDAtOrFfRb5p/DWj4fYxT6d9q1s7OXh2DvgVDfb0Sqc4kcSqGPbnAYD69FSc5eG5rTE
iuxErsD47xlegLn5Ls3Awy5Jsu3sGMSdD45NzlWzwK7eTMasnS+skpvTLXxMfxM54eIA29cg5oPK
Eu6d0v+vqqW//145099H/o4tD/izHvBNoBYdp3GnZNiSfbCRjW1F7gxIV9023LZvBA7qFTbFo36q
uwXxU2smSxdojDGpNytfxezFYyzl5xCihi75Y/NSoj9oliVJl4lzGvtYWRU3ZASgU5angZ9EDI2u
C02zfDM+sEZBnU04QR6N+cJJkRW3nGCPote09isiExMebV1B7JUqwk472RyIOc8EDGdeCz5MP1DD
OtWcOhX+DwdPN3seHmfxqKG9R6UdWVe3x5EWjpsBoPPB7G4IzV9XtO6Ah1aiX40YeTAqs4JMkEJ3
0s/FWUUdz9bY+IyISfIoznAPRoD5w4Jvz6EOMQjCTtjkYuV+Kxsk1q7jWmoSmvgHrEHUuVGkrZ/i
QmyrhaIMnVku6oGWUlrUyywsEg5JjvXYNoS0uTbPbTXMzl4EZPcbCmeWqUCh5d8hsqnoS9WFdpPN
x+3J+O9cjFk/g5+UA9r6iS6j6fDEhQpH0oDG7ECcOFsd68fdijK3Hi5cy8xX89GdFhuVyZZgnX2t
k0fuqOkxUtTmfX4YV5Y+8eZR7Tad9GB7BqhEhnMGmjXZPeUSgNV5xIytovJomhwS1PZsB5+MVLtG
R2415NrDhpAb8tvqSu9L5cAslLilgHFxGI2yNZZPvX3OX8hpPQguVFxqiVTBV8yPkIJCio59n/N8
dSqFP9+ZiPiw2PhcmIqo/MoVQ/Iv8dv0YuAXE17OUmxG4/AIkEx5Si3SR/ziNlicZeRHfazSLNfG
eRT/TFB2EZ7K4Ub2Nxu8CtX742kPpoKX9wEVTIoz7mXWfSxk41y2T6JO9gc/zx6wVEePuWwJCkeK
ndU0yPdrFWUZxujyFlP45xZI5P47F+GSaETFAgD+cloF12JcsSZa+zONf2TCHALoqH2twLeG6gLs
nYHS0izZICrKK1DQYAlXksj2E1WNAl5OhbOG8KPATUZRpshwBB+xbBDUbIPD1Rg1BPbJU0U9QTcj
elv/FV4y+2m4kaPtWUAzJ0PyVzwtEy29/bJqy79NsTvyn3UrCbBwqC+TWBX1p7V8HtiuxqM5npmJ
6sRJ2694o+H3uVk7AweVuN6SFCLy2pxXv57OQwUh3STDrJWKTLpqXDd+tjfUs2PEVnFmy0qMD7sG
aWvIqx1rpuVdQoRkPNUBAPiHWXffSRUkxgmC5IkcRUkCPB+KX0rS/FU0HXewlcXkg0+7IuFlMby0
U/TI4aE/sCBARkEDAHuwkcjUazHiF5f02QsyWhfpyjSuu5NTtHPlltAOEIu82BzZtPISYPEgDP7Z
vp4eXIEOBFN5/eXJr4tOpqNG8nX9oaZz0YCf9He9+3J48+wjbArIORlluzhu+9tfWCfuwt2icYYg
DWpbK62U1cxkQPSGJoSTWPintQ/o9y17Micbt2Z14NOC18KKDVpUrvmcJzGF5JQWtGisjDUgbHj+
1pCRYmKUKRzQLznvrqMl3KWzTcUZiBDCTtNsG7bxxPwtqcpbsRjI0XuVFcXKYeLgZBRi5kZOShHu
hZhL4tjB1cs0uB2LhcGTBmBzXvgy56kPkL4dtelmxhOJ7O4Nm8aI51/TmkLl079H2WojicIYaI6Z
C4+H9eogQO0A1ma+zKIEjZgkdVp2YTz7CIAcba7qRRI5/1cXuwmlP0WLmGrjtR+WaOZ7w+tEen8K
Yopyag3dkumT+EgVyTiezP/lEorlf/vJrxeX5At7NoLdvNZxyuxAvKVpXhE9EBOQT/hdmxJ6VyuA
okCA3LZKbVz9nGVFEgkCqEP9Mc2jhk61ikf+BHyCNNHZ4vuZCnraQ+hnQDpDctYkTYqeoit44EnP
PHlG6OTUbaj6vIoESeDnz8iZ79MgeYnkOZFcVRi/zokzJYgmEL8OCfJrEl6A5WPx5vcMXc1jwPIm
DBC6r0t5ELEaIdEsd+ZjJKWTVNlGovqGWqtC3kjh8H8PcZyUs4qKna4wOcfpGCl2HGnnQznKeij8
4WRxqa+RJ5wKjGy32FQn73UTkq2iCovVW6KfBvG7pHOYYVIWzKre+OS/aJPpUdRbnaTlG1j0R94r
QDiwtA9dXWf7AwN2TL+2/mD/3YVQH4ztSExmGzDNJ9t1Tq+ca6hq//tLZOc0cFX97YRgXbjsLs0M
RVx+nNdE+GzhEBR9WSV4jXhPW8AoVV1FiphMo/E5UrvCuChcH0o2XH5Yplj/7YzovYJeQ5psQ8zR
of+Hg3VghXgWb8FlIPUMcstjNl+aOxfGd+kFMaFSU6G9QH/Ri3F/cE03iCBxX2XH1s6gZdGwWk4Z
ir0IEQ8CbP6RdJbUIB5Nvf7ux179dtwja1XbNHfHRwtVAj6VXKLKR9Wd4hBanW2R5eC4JMviYzSo
OcPYqktgYXBgU7Q0+IrFL+Qfwax0TCPAN6wQaGT2ICGU0V9n8p5anysgDo+xQ4ECLYj/NcT7gJII
fmrdu5IJBhntWuw9uBlJFWVIc0bXVWB1fP+v+NVGxhm2kK57lnCpqD3NYlG8EZyLuA1KUAZJgm0C
WIUVA1iIierOs31MWkX8ys7FFkVLGrVwaASIRNClf8xykEKEXMddYOptu9uN3psF5CrtMWNdXNBQ
xlWvAPBmlrBTusQVOWLwLONcQls1ReDsYuieLMm2iYmdhwCn5LnGA+dzlMZM0jkPVp1ddXuK37Yn
2+uFgNRHYTlQEefnfb8+8Dq/SA1HVZ5xd+mVnwA6yg4HoIrXNJtdSHcqh1vF5KgiLG1MBudWXRBw
QbZvAxHYsvj98SB6ht8Zvn9W1kw8ToZJ3c1lCI0MeyMroLsoCLmzKqMwsBBeR+avyuq2cuzPIO26
tS+tcs2PHMuyDwCuWB2KgmNfehEKW95LZiC0SWTkoEI/yy2/XEI51eh0DqSFl8356HAeAfhin0On
aN5V8Vswc1qXE9X3hkoMmPpaf8UylBo5oNeG2K77MfF/Q76Vjsk/pcHh0DKhNvc+WJwuPImW4wJO
O2HJDSuwkW60FCvnQ+TT0zT8LeX06+IzsSIDA+cImSMRyZx/sKc6Lg/lG168zikkJ6rg1B5lPr55
7RnIrhmrzXCk7BgSfmtHZS0wcOAVaagMW9wZvyFQueVg3u6ozRVXoMITgfrhLSKEbZl/FabA23aT
HwiPWgLuF2+5i0O19ibpXnCjarFkMMAPZ13fIaSuEYJS2dO26IlTQo0u/xe8sQ2DuLFfU0JrhLd3
BXRfqfP5OAKOLm/GJuxFyqrp2sfTx1Lj/R55i+406P6iQKd22+UkjE9PFaOARSX9XxqLUmArRTB3
iZGe3GzgKvLmT/fHt7Z6re0lHOqnrEFvrAaZO29OwMEMSZODAOcXEWcgRbvFTQXZCt0EKPZapUzA
PamMmAkeYPBS+RR8g3lHLgmmkDOsU40KA+g7Zm1mDlxjBNvqdJGe/p05/edlWxepWyGskES3uvef
F2aQL23+n/xWkhHvLApkR/q6JTl7a/GC8ZfTRrE+NkC9NjgMBbN/dNEel46eCcViOD8m9d1PD4OX
FuJbSDRy739b3qhqe66/zPAGn3Ho7BKdRPRhg3RjcqLEizw9l7m2zKhySnns3JnIdvsrpIg9w0uG
drTIx4OE83IT96HeRYVJ0Rw+GnF1pPBfzcI9r+3z0PDzkNcQBxc6XzDMVufAX3ddvedGf3ky81j8
1BxjCIoQeTDUG32eOgy6cpUxbPT+b+mx1DXdiTSSRF3nrt6L6PHArJI6XVfok+iI4uGhmEr7Nh6F
lTEp3aV+WqNWL+vhuHbnsa9tUlXexBDkODP2YR2HVGGTu5IPftZjJ3nx55PBqWtf+QfwHxSLWTUe
IqMNXoDdj5aTCNi9lAwobRPmyHmipVtKBx8xwSfueO5jc7+nledhtCO3Nb4CBCJ4j1/oYoOD8pCQ
8eWUe05y3BrNV2bfHcv1KPS9hxWLRIYfCH8WCDwFAaBJC0cMGkb+0OHUzOoe646agCA7BZ5rmkmy
Yen5eDi7nlHA8JLcimh8chqpY8BjDSx0dUL57blKjuGqUpwsYiMssXo7f5bohlOazqhboLv60P7F
pT7r853gVqmt6kgEQMvCLNdhFWCYBxdHLtspsmsBeRHdrFu63lJk+KZ+JV7HcxsZhkDpLdcd1FkX
vUL+BJIxQbIH1aZntrBzGFE83MeRwzpCpvCyevNekH0FrkRcyCHM1xNQSDmj6Vdd1PpIPiBgseQo
jV0vtj1h+fwOr+ZnyNE6vi10N5HdJPjDicGxmYsEj/781maaXZjEoqV/IGRbTDLF6JVsXcm9Jv6C
C9t5khxXyqEAy/JMGievTjSFWyIb8pmJ27mXh+jeCRzF5lZnJ90x00PlrLsginK3ESpcpHNL9zSk
4929ccfDOVMsaiKuHYFKL52X7EcbINxZHOSjFhuRE9E9m3CYVmioM/ueJ6SmRbhCMJUTpTouJxHh
4vk9RiJBgpGmvytbFJoPT89SQ0weCcRMDSazqFzpXgjl1gl3V4XrNX6sqy9mOpR/3n1ICP/xZ1tX
hb8H2mmdHygjtcRHamkxAS7HCNhCFNFQvvEPq4JgMLFkC/dRPS+BFpwFFGH4/3OkwRZ4rwhoA1Fa
DZAif80mnBLAv+QfJpnsAwrrjsSrUqbUpJFPUn32N0l1LRCYrPNZ0R50FGM0osjS2yFm1DxpGnmO
DKM6Svhn/Z+T678GmF0z+x+RSAnGcNKGq884OMvAGzsJHVijJXKhPQ2uE0kVzkkAuJ+d16mou659
mTYj6kJfR3GkwiSKgF9thhX8wLbhN9IJgo/UvYK+u5bQPDH0XU8+eQy2UC64u9rVU0HrlAIJ3KGp
Au/efQ0wl+gucR0bRg3KBEq0b914cRQqfD604zPGNnkatX8a1qDmiPOrEZxxyEotvsS0ezfT0qE7
OKZJtK1/PI52mIf9d0/Ho5dMJy3uMgPBhWE2hgpRvxv5o2W3550gvvhu9Ng6ug1WLGmaThLgSUL5
du5awjQX6Bsbja+LfDXNROuUdswk4t65h2KiUh7Oe3cOjFSGnr/CIXf8CIm1b0zwDBZUqpK6CyWV
YOHYTdgnH97BK/2BFtzzJc18KWcsrmbCOGrm7eeIzoLTDBjvVYm/tQukhotqrcOfXymAkgjIqlUt
Ti2dn/cS1LOlx3CkUOIKckEYSIGVSgXu4/zn5wncqTQ3+WZIpYWTYOVNznN2L8RD0RNamAole8l0
XYCEXwcj/pKHdn09jMjCXUuxoWSLt/zBheW3lhr60T+IvNgwyXuk6sjFEg9e4BRrOG21rDzsq7JD
cjoWz253q0iH9FK+VqVsd91q0y7QYqF2F6NfPZnvIEczAjV0WqOTPpEyjzS0IrYcPJHC8MLTFk57
SdPER1oaf7nj3Ipimnuhmn2ICfGkFoeBODYUYCue9lT6L1+ZCGB4JO2OjMSSm46OriBLlIJOsXxz
kYJXWMNcx4qg8CRvgMf3MHj+yzIswy5ZQl2BL3hyWU6f1CueGmWU2nG2GLMpMRIjHWcMpjfmFSP6
5zlGcFgwORMM8u5kxfy6KgO+mUlNxeHQuAJ7V7cL8E8m3/eYs992/d4BsHjtjBmEHYxlnxLvIIgp
+GFNsovziKgwSqSGlBSoSC2mF1FnZDHYEXiE/i3ecsImvaMgGBXV+1HYPrUcR2X/5R2TlrkMl8HI
h5Tg4S6whV6k+vHdM4Znhsoa7S3qCl1W2mbUxLHZmASDSk4AkcuNyu7ZP3EADORJsmh7QDG/1/ur
RP1RePnrMXHDcMF4bfVkDCEZl8+ljMaU01/CTHrlsChNqQeanpKw6L1Qdtx/HCWFUZmvGVT6QpTJ
OYytaRYTPRvp2eSK9zKmqke56vdsxynCu8iBmY9kbkPEVZ7NI62xF+DduZmd6QpMypRlhDwgxQ/P
rOxkfEtj83r2HgiPeOMVWfV+BiXAA0VZhqH1wcdW3X9XcRc69Nj/PC4c2LKiGQ3zXHyQmkZ9VD5X
6VWdWlsBt/WHIF6tv+JvRlu9AR3+602g/txOVYQ58vMQtZdFsVAxz23jqscNj7O6BAAtw9Kdri0R
nl1U0RawWAKjuHIsKG5X1zOAdGZ9wbw5F0Q+mYkXH6acn5K/5CJ+AF+nK6YZ7QY8Z7PX2pMx5INE
gfrYu/MYP8dBJiUKi/C4wNriApiaHSDQZn2Uno7dwjKnVSkQGTTaOe0DFx25iBbA8w/bVVbTwP7w
CJEl4UOYuIFxC7I/5jKVkgxtUlusDoYDpr9tKp37x19kJxPUfe/QJ3f99fNpGcCudLvp6WJlvjcU
8Hj+efmhyYkLKcXk+VbMlGK7nKubY/2S93z6C4iPvA2CSyZWrjWqRplj24R6olJ5ua0K1dhVLFhS
lD9ZZreM0VxtV1N0C/Nhc2x/D9HlnjBMuvyGCRQS7iaMskMrrJZgxiphPJw+Mx2u5rgPr1cyT8+Z
gYfqnDGdmZgCPzKHNVLOJik0uxwBxc7INIxJyOFClC6Tq9aAKxj7N/6UeukwJBNB92iV+WWvW0qN
8W+g/ZZLRnqITgfuKUYdi65OkWuxIHx0qoUTS6RxiOJwZP4ikfpknYXm8l2Ucs7ajh02Xmr+WugC
bbFBVvgRzg8qH9aLABRVEo6Tv0eEgIh2GUnz7+QuQxF9X0n9ssGSsQeF+F5xXrTXJ7my6m+BBW3R
u/syz+lomMjRYxbE2R10w7HVvpfJxq9IW+WDg0KCnvfNjcbvx+duKuREw1dIu8QAcgWK2erH+wLV
i13/mj1+949QWIsCzlAbCWKS7Th3BLk4yFl0X2rOgaa3snZp/66+m2GndT00xqUIk7+A4EOQ31q+
M3jSo9qEEan6V8KlbucHJLZgPRNMc8BE30IJtWJt/bw5BWrgf/YlFvCQIJcQPQUu8VvqQLt+egZ3
Jun3Sn1EfV0FZbgKtQHnJy+5mR91UVJ8nOAC0AqfD71wkgWvWpgvJSMvPZW1BMgHD2cSkIvQIQMh
yhD78H6QErV2VDTR4rMHSmrxujsE0M164DrhhfTtJf+kvixcvGXHzAYfUfDYuQKQiwPAbY7XRfjR
tiKYmGvTZblSRizX2Ief5On7kMxODJY/EWwwPxQ2RPGpDqEhj7ztT5ITbaSO8uUdKRGr/czsvMkS
uM1SB9DTF8Hh2LTbvZdocJB9re8NJc0+F7+HHngjai48Z7AXhbIxYNy4E9ofuP3SCWfmq8Fo+0xu
bjK1Ubpu1eRAD+2HeonwuwRNbKDi+8ViAwCh9UZrHlAtVMryj7fmD5rlU6TRVy8KJ3j0lHglp4WB
5BH3ZGbK9He8xxEjzybXTh3XfSI9uZ+5f+zRqkhJ8kawrJkGTJD5jf2e6hws/6QzdBnTEzqDQPnz
kGB0/HDfFspr2EKhqEBtpOUmLiwV2y/GUXRvCtJYZ9uA1+HdW5FdRHMSyppn04UOqPbbSOvD+Qxz
5IAnBgR3m2YjzqWmMeqKdh/Z1Bb3d+YRFOuHsqCGh6wRfvmF6iNBs65zqwNHmsOxoNwY+/8H6cZI
G+4ZkJmWbUmvNKX9pVRwQCby3zyxBo5mWO3ROUTjK0wAttruSWIsEC3IwKQAdmjlPxqPP/mYFi1e
c906EKFlnPMQRI8/XwUX4HVtRXHp8meg32fH/yPeO3bnHOb4cMCx30DO3KTRK2seZyvsPjQ1l/FM
QXkDYlT7355G7zJmEzScVjWqdIuTHHdIbpZqgocmMAwxNwSzzr8AMTrm3U+MEMv89JhSi5WNOZAy
AEaB9cnLS9plTeMDybscAPODYgnreIdMYCIdAli6THdGhKZG2Q1cMwHGsynUSHiP3jFX+F/Vo9Vv
8SpXlxONyoC1/X3mnoAK1kFm1HgVpIOJPA3ZZX45DDpoKZHjPmCZEMMQJcIN7Xo4o1edqW9ixrNF
zGeOUIpDOWCqtFOj770LqIt0R0bJK0Af8j/7zzqGpaNAM2sUQ46zaikq+kEOu5yfYDISndgQFufr
bj6OeQmrzI+wmu1G08tP7uUPKL0Tg0vrB8o2USZ53Xifv+WrMwDQ+qqb59XAVsHaNAd6ddCJZt+f
16O47dPtkHRwduR2dokD7gECirVC8V9ksV9jNX6rDDbd7hTyL8olqTnj3RkVO8m3phNiW+DbcaKH
wLdt2uUAr7Je1WnoxskV6IQYu9WF5LVlmgIE06ic/tQZud9Wuv8o5UMHK2ENos5xaRXota5QwKuL
Q3z2WiWNVHepSQKL8uowQV3nbuJKJG/rznIct2KcqzYk2TdfarQ1r7/RyqlnX18BNH4wPT9sb5wo
3vtue7OC/RA4ZeJFYT75yDb2SnukxALHlrl2zb8D200y968LXNQHobCbyDgUgUVE78SAuRXaVos6
kxeGq+uemirsaNOYbuT/PTuQ886nDj1JCeiuPm5QDuyJu8N3NzzIjxbPS4TjqYwORDaVhQOqY5qs
kLxxbKxJWIJN5RXR1f5CDIXnmujd8RvM240OSuDMzdc6uJgKjquzQDF3BKZZFdSyRl1Recj8Yjjc
o2FG+KCJVfLTB9OSlBPcAi1WZ8gZQYnoSGbBmxrZVLR8q9k+i2vlb0nNzGTPUM4QP2cUJIfNRnqn
lPCALpDnmtxjv9p8hZeuVqsvRVYsd8Z902nrivD4fh/IN3TeY8PlCH4cf6JSq9YxnO+ggIBakwPz
ck89I2DOBWeqy8pUjHsseDaneEWzppQPOe0ra/bQY9wadQ5C3BMItoaTLpXhrHByEmAcY9Ady1Se
9xp2yBYhStc29qJnph0uCwKWiV0kpjhLCsl48W+1eug3PPzV9CodRhAgj8L0mjzppWXup8L3KMIX
rCeqS13+PAkN2Zjg1EGRRFM++WEpiTFbJ6cfWx53nw/nsEGZgaq1/3ZjuEFsVt1ggsrBZbLrxWho
0r+2Mf7CZhNyaFMFXL1ckBSsndSVDZH8NVOQk7P6ntktjp2SdbADOPPoE1iMFVNdEakSGzTeOkry
cnTmWRcCQiwIQCQTy04XBnfTatuZEmcU3+kp+JiQPy5gq0jhBoigI1enJ2IF6bP7kvN361MXdoRM
Lvev9LIEOF8MMlY2wTvwgaE8JzLHgJ1AFRhXkXwUQrMN/gFZdaxvl4Q7KucdIrBeBFOlgvZMSgV3
8jwen6KVHzZeT8cGMS4G3LwAU5VDqCjM/5qjO0XPPsyZUGkr6VioEs+xD4P8mYmb0MTEI4owiNAq
DLKNgHMjTjRW2LaiCI5cUFcGwm/Ohg91b8RXyBDyQ46RDgFu4JPU3VFkW8x8mkgv/BT6hu5zp2yp
QcPN+WwL02o5Hq/4zLFQVvbz15LUOj/xeXyXSS6hamWAwAaivQRf4lbvn1mnJ8CSwlDGQbz9b0Gb
EZNJ9hQUx9bQO91R3gLQIEY3v9XDNfqB56sVxHGgtjOyoA98VqmjnhgVeVKKSvTP5Huu1lqJPhr6
UuLyQfrRYhF/yJ0J/wCJ5bUX/tkbVUsn+nopF8s1I0PEApwSmZMnzbcL5Si+udWtI9MMBYd1rA+W
tQUp/dkWa3o/7HOQKwax1oSg/6JbDaEl3L/32zwQs2hZR+po6jDtZ/XDEUkionfZrPLmI598xjVL
cCNdIijhtAjEljGG3uZwJYvom80J1XV0XGtNialZNZhE28I1J/48amst8Kyhso1bqlEBWediwxwp
ySeOPccDGN7KtnWu/Oge4V2ppstYg/cpgq6oZDTzSRiSW+mMYCYJk4qFZW126nvRGrwvrvmw2Zy2
5K1IcTsm1lf3eranWnmyXSMdkG9Ueo7QHIDBuKtu9D4VfBCKF7VC9Vy9egGC+zJQoZiPFw2ycmvH
3gYVlRk7qw87QiDIOfkCXZZ3+r8ihf3zsF9sLHz/OoMr8u7K7mcOh+dHjedqlaJYmBqKntmX+3wO
vnVoauwaQ5W+Dc4KLqIL4zI2KO93ZbAMFbtqt1tk7GHUZXaaR21FRa8zJpPJuXII9zjc3F4USG41
ZCe1eqynWS9OFtwpx83MlVTFQzWnNkDUONrZ/96/gJeuFGZhcapQ58JiWoPbTl/Y8qR2GYZyGxjL
nSvEvkcTe9o54klxsUbyM+BypAWKi9GXD2XDLVvmPw/cwBgnqBtCBofCg8dfB91dEpP8isslZ8UY
VU6dxAx2fKjoTM1DzbfkeT4M+piva2boEgclL25ErnZyqRpur0bUXXHoRYNbIUeb4qIgiJD0e+dR
hKWYSTjD/EkDoag3o1dX29uLPWNfJzp7dayRY8v0s5xgDeBB3vqrLaT73dnAJj4Bvthr06y47fFq
oHgshP1/ki7jEn1P54BAICNG60wJkDrSX4QqM8thtpgYQiU8S5vv9QMEBAcuRXvEyP6XEWMArqSF
CNzvmqzuYzyAQqn1Whp22p7mOXGyGXXSM01tjzodgvdX+ae5zjnlYiC2z5WwpSlpZE3h9R9vTVU1
OLa+6UgXG45a2Ys+QsPHwx2Nw2ItqmGGgME4BEW/W30gj1vUeEe6SsGcQjAt54RCtl9LiIsfOn55
oOp9d9rYJAbIQHjGyc/ka5e9YqEDax9ERZjoEniZXNW3wDAeI9+rcCISh7j2BYDA8QEb9+ZRF+mL
VeGtTaKL0YDRoFSKX1qP4dfXFyrCN+h6Gph71Tdd8zjeEIKcEPiiInIEHGvx7irivNmzPTuyp/MM
qRK8PxkEdLbFdeq+FX+x7Bhm2Q3fSq10wtmuxTKTOWbXd2HgkCtScP3n2YG02adIDUOGp4cG3r1f
smnlrSb0NzKs+aiOqN/isSS/uZaszijSJK0rJtwURtX2+bPXgdW46ceTNp2OL60UCBdBE4yH2Fkh
oyv+KqSzmsFotI2IOt19H6Xja2QzK//Fg0sAyqfFk/XzfPWFL6FuY9JGR2kehjr+dEbiyZxpBhsY
dPExo6Hn7SkGX2+0KejqCeX+79aZpYInVCPAPpYzH9j3NUyykpaoW2cFCPaO07BOW+Xg4nO9uHc2
zqYke1fllNQ9MfhP0sPbnYztreaxEaUlNoKEWcE/4LQ+ckMLvnEohiDk2Thp5SYuglImaba4zC0X
6yzJZ/hfkVRIWSOQKItLn/efzr9GJck3vZir9NfAEKte8A3s5Us+OwLyk4hHUp4rluB1DVTIfU30
2PzMP4kILpiXQNnF+Nyw8MoBaU7Ow6owV9jvDaIo6FPOm7JjT4b1z1pfY0yeaYFnqDxrP23HkgH+
U8XBP+riG/1srMVIXhbCacdnd5vS33fj8O/e7nRrp3xa74EP+tNtGLBqn34WdytqgJ5wnwupggba
IYGiyyTZLqj2TcLZU02xRR8hQVICvj4An1b9vT/0rEvrlqVv6E0GFUFhEJw65SZTVv0/PgZzgfKC
A0JZwJdz+cJU3vbIpZvd6aHGtylj+L9iw+/yKr8g7rNYimETDS1NqU6XfeoZjPC2rx/8yAs0mBVl
DWmDBPoBGlHRvVE9MJ1xWv0+n3h8UqSdsUXdEPfKHzhp3VnCAHAehnLfGH+/xlirgnXkpIh6Y1TJ
Vlf5NQHrExyOgXSxw0EjRL9wfAI8PJ2YiuCOZ2Een+G5p1UXN83DI+NR5g9UwvEtM1g1A0qCC+eb
5qalCWArC+oscDwdJm9yUyRe0Y0tevEyh61NYLckluUIQVefeFEEAqhvpzqZCy7myZBLm2x1Hijj
d393UsgSrRYdffg3Ewfj8cpCu8Zney5MEpJ8wI76ibpFvDVWxrqsmKM6fRqoDQ2DM3PTLMKEtxyx
VXYJrEs2tI+ftJwDjQqVWvqBWxzs55jSh1pilBEwV6fg/AWVPuGVmwtGcKGfCKDq4FXM+7TLiIzx
DYK+XsntHFucvAq4/aCUSDkLG8S1MbAAEAyU3Q/6LES5sMkEXXpB0+CdxUoS0RiZYVP77Bj1LRDi
aE/R8WF58qVI3cMk7b6AN05MN3/O+qBz1Pd7VFhWWNbJzdFuS9HZJ3tDCIxr3SfPeibi7yj4cROw
GCvky/nX+Sqb3pPNbl4NpQIyYWRG8EJtYombDa2IxA7Cs0thcLv9iiGiMWDv5HBmocojoebaCsus
D275NUg+vLOMTSFOZyC2+x8UUhKF1DQ/A3IGIHDOUuh1qEq1XU5U5V9G92Ue+wQZXQSZ9xiKdtsS
cjy0bbywc2KPUr2+d+xcxkVAHt2RITxmE613jDF9j1lIJn1Cc7guJTG2EDNzl7hrhzJZwDx/qMdh
eSZNUp8vhTAmAepLE6aygEcfUqJgHpV1JAp0KpNxBJ5lVowoYt0zVTClaoF0P/Oj+R63EYXUevOL
NtU41/+SXRJ08R77KJepoZzL9uV4s9vn3W0bdvRYKSIXq6FxlkSoS5VsZ0ZJ8JkNNsPhtqcgIDOA
64bc1nowJ7FzMjxx83KKfa07oQt+RsLo1GKh2LZMwyZ/OsDUjxbSjq7C5IQbBUJ5yr5cuupklWd6
m1P13VusVOe/klAeCtp74T+CY8WJSlkQaMQTZDFLpfHlg7aZTbPHBhPTp222VBdU3So6Jr7CLEtS
LbO3OxEiW9bShBK8Ndl6GmWqhIapp/lc1NLZGbCukjkLeuPRbtc143qWm5eukcCdwzK7nJ9TuGQx
pHKQdVeW/ssGPauWftzWAOlY4WadIQoCIpXZ0DcaptxYfyENKqiLlwkB/BSVj23FauEG1BRF2nU0
y/amDkYo349piOLt0j9ZgdXUaYx4D8UqfPsHOhj06anTxd5i7twsfj3cl3GH8thNTaQZg8ppyETi
HeNUM2fdoDurONLuCttWLAmQ3YznxrxvUkjgYYq8jYnprs81qfdrqURLANakzqVTy4bMFl8TF4X3
wV0RpUSYvQkg911eRr4bO0/nq6O76deSpgWFYfLcOENtcx8AXvCPCt0gqQio6jBDeDp3Tm2JjM4y
GxlPkIjyUTshQQOcfAc1Z9fud1/MaAFoZhfINt8NWBiP5evn/OhCIXM/0t6zIjaDonG6ej/ZFiWq
+N5rx0hbaPo6vSkmNZflJToCpndSrqaoE91D1txBuQjOtYqHI7zf3DL5NkzY21eNcGEo8agtnQ2J
24+xn1wABDm/+hrF7JfHh4uMrU7TcHlQbLk1bHfj2R79c19M5FS5f+mFt7qgqT1yXx6XQ0D4D7Zd
jptHBNS3p8U03u5a5Z2pOKrabglDFYyFlYpc2QkAo/BRUo6x7EcJdHS7CZnoDRxks7bf4unj3k0w
DGRe0Xd5lX/bnngoj/ZzGRPsG1dCJFVgwYRbJdz+2P6/hBtiVD+nHB2pV/aQvJIQUOKgQL+KNXis
cI29iK+G3CdZT8l0JhTSFktraMBFcOibrOfDStjevWk9zjE0HoJ/WEWYvV3uFkYNluaF6I/1nq3q
gAwUHD9KzK4aOtsocvqbNl+jz3CbCJQiq7VDagdK57XflqldyctKzsZObnXEhNSCxmhp7PX8MZfm
B2phGCfHDZuFQSWPVhkLusvJYRIjXynJ5xZEbIlZ8mC+OQmutHDB5S5QQzcnpm4OU1vl1x9gfTaS
obqkArIe5f248wcUblyZKuTXGUZAYERMiBGOGTacV3ERQT9gJUlewakILXTwa2Z+ypsV5XRnCXkw
mK+AS2obMA8b9g9JqId0GJJYwuwMUbSVcKbfewmFMNFNOSg2y2Ne7SbD6rlG3TNKpElywKPs+bug
DTJEK1yNuPtXPePFIe+u22MNr+v3czvBN+20FVNapi6VES2enmzYvv8IhPc3PHihz3dZQx5pPmIX
yHz4stWqW6oWQ1o/6oHo2yH7sHl4qccVCXOWKkmkiLs/KDqmXBqEOv0StRbvL01bGr7W7yWuweXm
/4iVSPM4jWdVrFl8VcjEEQM6tJkN8mQN/jVJs8eTFcnW11ogrEYovKp3Ks1wm0TK7kl/temB8h/X
VdNZSoG5kVCw/NDl5jU4pP/l2oP4P6VBsLX7MuTI6ocXvpZdfs/24x7qiiet2zsAzsjWTG3rizLO
t7dSg7XwVzq7p28GofPAW91Esi5CDLuEMM0kRERY8psgsvfkIolYfWv5MmnKMXO9kzChCpFQdzI1
818RS9gUwHA7odVGluNC0l0rjdwLPHOvwE7w4mpe3jtaxBiMlFLKOFCfHRXupPtCMuV37j/MQXLv
59E6KiKKgZzCtBbB9qRfl/gL2IzadCt9H7SAB7BLBowj9rjGolhQUO28bXw8xAEa2LsSluQ5Bf8R
6ghI4kPPCwNTPpOvU0XlJPUkXBUfrQqGgN+pcHCILYTQmqZDHkldRN+5JJ6bHTLgh1ni0CwbkpNl
luRb9exWL95PC8//83I9Ral9y+pDaQyjH+B+HCFQT9S6OXV0CwwwirzAb1WBSDYbHvTIfwMWEQM8
KRhR2RKXDt1NFpRn/D9sg/BdKDA4wocHcv28WZhfzsfv/spamI8qoSYuq9u+c3eftZ6E5aL7PR71
55nrAopifwOqi4VPVOS+PF1W6re0FvezM2JpcmhqL5B1bDTpHwTm/5J5DH0w2sDLqe99EK53Is0Q
Ij6ZIuDRJ/F6pOll8VoYE9Zjctg88wqLcE4NgEXt2NcWRMGVmYwC5CY7KM5jhW8Z9KR/DwVpjWN9
+PgFgAjBE9d/HQ8BngQRPf4Z5Bj11JTzFP17uTR9kAwGYvqUTsR9Ajlto7nhK2WIbqJE2SnRzpS3
8PpYxsNOLTJ3vG4Cu8TwrqJAjfEf7YYB4d5GU8kMKXKxDNOJfkWTRe1uQ8sVDl3fTkkmRvW6xkfq
ZJHPbEHhAwTHeycd2NnRNCyph2MaAsy4pF+GVXHRzbnx74UhRvZ5/uz7QrII/TFTwQbi6hDgc96F
sbdUZII5MsDZNZLIBl1CIL1ght2MzQ5+5xyrTrHTkZWLfIZFK5bFpJsYzKehBLCyWfmBR8Jv21go
h9I7IJSowzyukuiuhc0L0amaLVI95jbYaj9bSB4RM3cD9kUyJp+x97fs61h4N24rBJf1GUQcLDBS
0vGokSPfNkWPIoolp4Gl9vNBRaRVYfWPUrLxn0In8ILLBWV9A2PZ+Lz3HXe22HKMojIzzUue6lrG
7eAo8GmPgVQxXDgl5aSNQqnL/dh5w6KMrCPtMDopVTO9pwLrHl2eWDEUJqkLjyUzucT+ElMQfUCH
wKWH8asGD9ijcuewslqri1wN4jGoMgnJHSNv9Qy+b46x/NIrvQuewzdtCDDx0Ie1DhB8oK4QUnzq
iy7hFmmC9th36yyVO80+d9uRmLnjnYzBL2RC3tVkGxOKTeeALAIa1QSEyht9BkHzV5cKvDgBWghs
NuzunLYTwbrA7mpKxYCiye5sqs3TQilHF8H+b6+ytzbfkTYKtYZhHcDHbX9yAoimqpwBxcQb5I0V
bcLhpd0hpzaEpUnrIQ/M8Wvtw6ssPZ2p3c9wK/iT173dqazK2BWr/MCAEpeYIztkDhYNZTRD18B4
p07qFC902A4OjyabCunzImq6+WG61wKKqeNZu9NYAWfIyzxuGdVYC5PairXJt1ByFmy/2HdwMdsm
IoEzOB+sB5SD8Qm4PRWhIo5E7msgSL9fCImlwPCVgvPFZBW6T8c1LNsrXpAO3O5or4M+1CnhTEdT
ClWHEDxrXG0LacBQNf1sXSIbt3AO+BhgOvx6SCYTa1B80LbbrQgqsBryuAUoIzMQUrT5Mp3087ST
CV6xVm/ABUXesE6DZNRaxMKCi2rQfyBN5DAXgJoM6ayRXiI6xTh37/fFrwmm37xqYKq7DA2uw/tK
WHlcWPqRvDf9RxI9pfZFuSSvYRmXi1YaiaLmF3eIEeAODEugoFH+K6BOhoSt3WU7PWuccAtvAx/k
UERoRMCax83E6jxMLB4aSSdWyC0qYKtFHekguEt1gfY3sBNGOoq7qsgdVD/i4oTlXEJx6D/0FBI4
id6AReqoZqa3UUCNr2/Cn16j3DqpgTIN0BemsDztaHBRtNT+x8MUMqslSCqbk3eM1vZVhuRHv9Y9
rK+9asBkReoCPCXIqLyZGAEO7FSnM+gFpNS0ipNXoWFmmSvDtCvoT8ZIGJbozIyXJAKADEJhnfR4
ymH77OuVTpACy3bKY3fN3NVcHXJNLw31oELSJNN5MntnwfHOdYFKd3IEEVleEHzPmVMAhW+bQ+bP
iXrOJ2TLbO/Z7fWL+a3w26ZLr72llY6iGN/AsQoNxtYQzwGcZeafuMPg4g9tSYzrMUiohPj67ZGj
UG5zV2x8x5vwtRHfDNybh7vGMz5q6PGnECN2c0tIYJFijiEFSoWTTimyP+YszDMhMKz637hUiQsz
SECnxSF35zwNok+PghAnlljSl1zi3q3UKPz5h8cRrlYZIhgE6g8/glSGcJsEL3IK0uc/OrmmvD9s
k/xXoibIk34sIsjwE7wewxuZ+kbG9NJjpN4tX17EyVkNv+cNuXUtG6XHZ90ffqCFCN5uxdQOousd
u2FxyQguQthqFB2NhMrq8/UABNZHKVSy5zgM7NPL/vi4hC101SXXLoaDaoXTlogG85iwPPIWy1Bl
wDwvIlH1qjE8Yib/FfBx3PKWSpT80K8aGiudVyItT2plVSqBh2cdXBic1As/vSPkSU4/3ZmbqD4s
rjKC26StG6MJ527+lVFPk2ybmrJHmEhiVGymUPklXO7Xy0UEQHoSJjcS9TXh5p/P2ZgNLSfzGUlm
qEPJRNbxe6fRJym+GOR5Bf7CUesHpe0d1XkKSZNPr7Wb+YyDAFd712zS8RubYrNXfG1Clfd7ko7I
bssQh+PZ+k0qG28RT5pyoEBfAgVlrt6k99kjtzmazmbCeXgxZUtNa6z+JPP4hfmZDkPV2Jx7oxPj
qJ7TpM3EHihFF+Z8+mU1FTRGcyp/UJklyhV+5y1PfdTBEJOe8Eqa7o6Aq2UGJRsqeuAobAvQOzb5
mA58sCoi2LXr0uGK/N3q3yXcuCJPDYnIwgNWdB3L0DrOXHRqyYGyH1yauRLPs92zGHEQN99QVg3O
TcDWidb1SGRlaFjpchH27phALN+ZadNx59BNC8Bg9ImVmmRmRDEwpIw52vr2j5+EDnUB35QJ9y5X
CVfMSaKFsz8ISAYYr+ervoyscb7mfh1oUmKpwTG0NjnrBFYk9Fo0UZvG5OZozl8AyVpt9noLfg30
MhFmhIIeN44fc10UshF2T0HLF912hZpZg5PSN1cPhGBMOFbIlVuxDDKIgLYA44P+Gvf4PMnk9XYT
PlXnmZk1R9VPGfAUVuVLZnf30mXeCUPjrv19KXiQXHtIoVV9qB9Qm3K8NFKNwUnEa2cRZ2UCDMHv
8bua+K06n+P3lbFSMK5cjI7gA+1WixyFBB6tVtcvJWj3i1RgU+SIuKUxD4E4qaraQlV8bHXp9EEN
VbHVl6xk/P9oPavdJh1B9ekZEKexQxr2wDcDxP/b0PIhPFtpZG2Gzme36uTbKAxVwXZlgairwdWb
Ib3eFENgpfapHF2fz+Un55VpNvmkjrLGRiNv675+ya+s93lSrdqEF/OTaCCky2QkyK8Vd8JIpJ6k
JZefyOpIQyfvmyME9pV+71aCX58yhRYemMjtNED3evnM0D0qXNa+bL8EIDhHsDxIP9+lforoB4he
jBn61E87vLroeMXpqMh5AqTwk+z3dnHJh9yk2TJrdUuIK7xcGpgTMVxYKxpZ61iBDvcrrV5uhMFa
v9IMucZscwnC4jS3MIm6KDSMYdnrDXNDZkJb5VyHAUqkt0YjRSdeN9DBs99w81ll4BAl9Uot8l4k
3el0jcrLis6S6i3Nyrke6P6s7cABVCBvMcildqh+TEcV9YzuZnUyNJo+eRGMflGFaUP4jG/dw8+9
cSC2Eqhh5qNOCoOuqC9+Rvdzg5Dzane8sX4+Cs9Qi1mVRWA1bKPyoCLyvSs0/nK9Cc/7WKFN0S9s
Y8jMMxPOemp2bdaCTgLKrmj8f5/64rXt6jLNRXxhI6TZlHPvQ6b8uo3AwR0u1yagQwQKbqEE0BkJ
fsydnFVvN72Y2p6YT1v8ac5naS5t+0ZjEq8e5O2XmV/YQljUuHUPZgVP5N0K8ISH2KBJ2G+Q4DoN
uWBWqgSXDmGrvIlMsqTjG0LqBKf0PgwQW83IBPvwX9UelRbxTFepl2Vlqsp/nGtX/ci+aetnhBJT
2NG4gZWAol8qynq954voRmswpxm9Th+F5qIKoVPoy5+qKe45JgM/78aTfdnXO4aEuq7Jc3ACiQCp
t8lQoeGYaiMJAAYY2rFLo6hCOZ8atldB3mSHH9aRBeZbpTeq92gVblpvmiyfsZIU7WQZgibVqUy8
NbA5tSLFPCjiESfqwRa3NeC1iVOt0WB6i15FDLUF+HqCfScrc1edIHiKCM6AtCDhCGZ9JASUrH6W
faKb3yZspKgu6iE5kI0ldpurq+Wan+1xTLhVY55tp138wAh8qs45arAHY1QiE1UM9L9AuXHJA5W/
2FulCVBRsaDNFLc2PLNuPUa3HeTJivByTA4rrSZK9auaAh2LZoys54fA8DfDWdQik+WvwuWyoopl
u6FhTCTGsd64d8blXD3DILwL4kt4msCebsSFcVKiiVe+QZWolVnt0t3dUmrPg5Ys0tASqIKbUvz6
u7XWjMACNR83eDcblPW3EcxTZ0gtvXxe/gWrKsRXgKi4LcPFQKUz3x9MuTE1rbyiv0/SkiGgqfCp
2lC6CnR29Um2hcfcUUJ+Lzv9DLz3PwHqR9Tcez3GncJ4HaX/sErML2IxbK3Xzap3pfDRmnqSXR/E
al8IblDasaJ9byDlEaV4c9bYCkUYAs2T70ggISXn6OjTSyyLo5q7VyiJ6Pf5Q5F90ojx7yMqj2Nn
z/CRZMuNaDSY7uFeTRIjxnILVMhkraDEFyfitlwOZqS2rDnN+0pJqbTXuqKmhdp9eXQiMGjfpGMM
VAPGeEe4Fy8d4OkOXuLuhhds5nnVMeyyoFMaGX6xzEYcaGt1QV1olDh3ljYwt3G6jTC3sKcDkFsO
IoQUOSdE9QBdRk2OSNZaKjniVr36dIql4WT/5XTLiIv7zCAGgMoB/ZTlzRvBV7BQERAeLRkHCiv2
By0b0K34bWCHrTJZ4O78IPB/KwHWgFhJv6y+8gZFHZZk+x+K8nettKB6PpIFmT0LbGAst0Mx52ZF
MSZC2ixmdQa/YjZE5lIY4oG699g9MqzVmigdwy9cq2N01yI8qHX9qp2w26E/kCz6CtF/LmH5k6pu
lR+al5pUXxTC0pzXikuiuWNPPzHsxierZPW7cQ9tBjvtVfEGFCPJecLtr5jP9M34JkRvERY+chim
DTuR06jcaHavtz15QHVxMqszyK6ksKYArI4A33PlExPmwzbMHkbuugM8FB1MbVSBxxsLGewTRvsE
70jdZ4EV/cutvr2rXc4vMkxKmmdQt4tA3HqrppIdhxon1LasbDf45PNI7x9/neibPiZwEi/wZMRs
c+AY5R8bUWT6caXruZDRxDjPsB8wnBpdWkcJjACJR3vrbZhygV1RzIrg75E4rTwOE5H25COaHUkm
MDIoZSoJJ6eEjxu0H61ney8V65SKBVMXq+QbfBm7WIOLzfNry0K/LP0ThtDOZpqVniP4SoqAqQGV
sjKTdw+cLtT5NhMI4NrjeDQNcYv1zYE0n3F/8XfJrCgwbnuPSclKfAC1zdqkWCYcqybfQH93jPWK
jQMRV2l5zJ49ef+f68O5Hb4MxtjaPyD+Z2M7w4kT5vaarpZbkLDePkNEt6oxP3Mcgod3YMhlBH/R
wDG/I0ug5rGUyLRhuw7rDWUqI403nmS1+5M5n7aUmMb9WrzN4LOWm/mNDhLaCx5RBCKhBHn0EOVF
8QrOqefDthnYBt9ADLXQLqB+LNiU+Se0wcw5BdqrpS5uu0rqr4ymnkpsps2BpD2aIJYNTNNJXrMK
i6C2AcNENnDSkbkYS0FgnVZPnNN1Ux1oiAzeS9RG1oataYhTeRIaDn6i85lN4CK6+cD+MyIWO12a
wKO+va5wckqn5PUEjiEItz2v94ki/SemVF/cXpotAtC1utTlOo0eMGdWlnxtnZOYVzFcNSUAthDp
JIBFUiBEOsFDLVgtfsAgGJGv7RQ8wnPmcARHBV1Vgz13SdxVMyzzmQsMgwKiE5CBsrVy2Bgep1Hf
LxeIpANf9kepw72cBwK5J2FxFUmFVXnuR6M/aw5Khn8atpCSePrMn8qU1CACRLqoYVBLpOKfMw1/
HP9wtuhzT4+GcFL0Q1kLbJJC5ZP5fUkjiC35fontrA46HoGsfDI3LCcjSvdBnSi1XQJ93tMVhigH
Nqgp5OTGgLRixHnv4T/Quic7aI5pXHF8CTSWzLuCwAqJd0N0S9tCAP6X59p6bjAcIZ0CjtUBcVWG
if+7sXDIUrq8Qp9QC2VAqKhvRkZLa0GXNxJFmkZihUqtuMZL4GgDlRYJQxcT0VS0eY3y7fy8Jzt2
HcStTlCw6hbMvYdifEEVPm1qXT2NTZkRYvM2xUEzqePDc8UZKGtEmCMJa3l9fAeDeM4X2CzwF6TI
Hb8HcYGfsdOJRWr2lJpN8E8XJkPvwD7+60qbyQJMfbJoiztagixe1XlRffCE0OPD7cHMVtj3+zDO
nIQBGBofOa050XyYk2ze0VWF9ikLeaT3HecwarWpjW9NbdUn1Q3A7Eez7W9qa0hipVlHBtuIBLAA
diFoI3d1kntHKerpQleWakB0iKoc/P3cX7n5aEMUaPl5MbeYwIh9w8UseQ+Quyv3h0fdW4MKB7Zy
44C0odAtQG20UX732I3hxxh5JuNPogkq0Rjdsrkmt8Rj/yF1IK4zUL7BkzCuzoc+HOWyi4GQNvCo
kER6IXeYZdbe9wgLuXODwsyklw3dByaD9VTmIv1GtFKW444b5100arPOzlWtCnQHStfSHE37neMK
5S8IoE4U6A7H9/qN2WWQGgVYVeMKMGqGE/KjPz6XdqUNJzQsUjXRd/52Nnd0rlCQwG7bIGcxnWYh
kV/ilhdSkyk2CO+s+q2gvQfBD9+zfEb+vStiCOQGEnrhLVfi/+zp/3ARtp97BSUSM0foCsS/Cixq
w5dvTXW1xLJ/EMlmXmWb1qKkNMwKUM2nxcLaUTU7O76L9LZojLzXTef7WxCXaBpYqp42Tt53tiQn
pv5LEYs/9NYSGXCsMQN94594KjSqsRcCNciUYfJLVZeUrmrBilLNqZVfK8zFOscsCRtJ6ABwIhRd
EsOjA7OVyGr44Wscpe1l0EA+FeGcgaF6Helxh/2sTTjIxiKmuVB8CuI+0OcVn8aD/171QNnQC+sp
Muuw5wqlaZIpbZ8u62dyQHdLA33Y4E+Zyd14uxYGMeITiBH2om+5JO4/RP8L29WhjCjWzEQm/nXB
F00Gqx7zjcCgjLCrBev0V4K8VFBkE9wTSla3IQTM9d4JeCg7/ihUDusGJ2abzFveUn9xNxWPspj/
KsI8xGhgySJdv24IRKrZE40ciHE1P6yLxUdm1yhUIzwx0FAMAeIA4+MWL0+VBauG8HlC5zmNNpTL
C2rY5eFSXggLIARgGnIQopG8uAHiD3JBhfhLcfVDMarL8WDgB3eT1baY3nYwQbn6hzlfkvmpjMS6
4E8lGcwCwrpjEvr8y4cRPtvkrmv3z1dnKpLEUPkF7S7oYWOC5aer4/z+onedk7XhNz9uMrVZjWk2
nBAu592UPMI3PLH4v6WZ7HpAVgGMrnpsfDX1ayoqbuU4E9NXMjMKeikpzWjQLJiXqWpzZUhwILka
S8h14igkNLmBaeaGKHhBassj7HTLuhfh2oUwdQIJEZzjZ15Ls5VZ0S4ezOf9+SzAwanDjjYOlW1t
zbPU95Y2hrvEPYaEyyN+MlETlMG3ROkW2yXlPE2yGn+wWh4hOwGV807Lj91R9940xUFfidBIxi3B
2tqrq3E/Iabytg1/0AU9VUDvf5kDPamJfAJJq8c+Uasdpo3zRrgD85MaI7yrW4KfSmthalIVzQM/
2voZe2yfF2Z2lYVK2So63hsJUTdsgPeQXcyohAuSQV0aRec3c9CceRBqziO8uHZpSD4Ck0IPxdh0
04Ex1NRb9yF3fw9vF0yjbHRfbicS7VdBY2YGhSb7LgY/gtIxANM4xu6dlpmvr4VgTkmwFITdTJRn
LLt52jZl/blYf5jcL+hqQ5TOqUGrFj7kAhVsPLVtwXbRLEJETXlCHGjOmVmfEVpT+EkSv+R//vC+
mGkSDNDMX0em03wMxq51QWG0suCFs8qRt3FgVoz3d2ZhhlOaVws0oSWRf0qQRd5HjFVe/y3I2/D6
2eD4eIaqJWjqw5GJFEkvT5vMI0QRgmVViKJ+j/RWl5fd8j4SaPIYDCfG7Y5DFfQ/whoQSMB1xQ17
t+/VHZNSjnmaosrMMZJLhUhwx+ASkdWs8Ag/Z/zcXq9RTyd++2qAPL2XmZVZZHsjD3UeGVfctFb2
8/gYunwyPUkYaQIF9OmKssiXNVqt0Oz3poMmUbyDzYe2Tn2ARPYCpTkmZSZasXES7K0J+xt59Shn
24nsyoTmKPxQhrxKLAnpj57Ad2WVcV/59LP7OnSf5LhM/HwcikF5riOzHbno5U/TGxpeNokzrUAs
W5UuDf8G+b43EC96yxBt/fO8KbvFNH1Xev8DsiECofezigJXtBoavKvISSwYjIS6+jjkq26KXgW7
/8AOXytwGz28AgmF32GhNJFBPX0UnRI/0CrWAPL9ziApRrrqj6ZR7vUY5x+cBlGvKos348xbtHAz
IC4qf1SJwFEz0Z83S7hQhZpT77Jq91gEySSVe4OTOAk9wCtgOnO9Ir/V3d5TKaomWcdV9FwNeBxo
2/ZrbNQkkHLBc6FVpN7Oj0JfSjGc635pz3TiCxB9urm4Q9IgULFl40W6BJM+BYTpzIs8hCwIElFk
5bWtY09zLhBMe0SmeangGMrMIvvHE9KYuJaU/jxtEiArhr7hT2W8AGSzFll32ckM2CDvP/ppTexr
1AAT+AZWvZWYW5B5Ylq5nReTv+MIXYmAM/Yh5gZRcpAeb6bre8vM8eRhcFiERFF7ie5bO8CALFzw
9AVLhEB6II6S8ReJf3ky73j6n9ucGAJMidEgOZ5WQNTiGlpt43r33rhakGB696LrB2SYyT2cYfcz
/Lz4bnIw7NMn2MD1yEQY5zDZLL/0TACkwh3mvS7Jwf7zSTBULxHEZU/VyYqTqdvO8cbP4L44sKtd
rhTjJ78cW2jo6Tqqz8Lk0HO0RDMU0YkP5j41Im0zliooqhhvEA2FQpDMDBfpnE4VxiXx+6CCuuTO
zj2ouuVhCCerQEfe96MmsIdGQh1rpQ4RbXNVgOByDdrZqnIED5A+7uTvphSoROPZ3DvTehOPBUhY
M7sghFR2QcKRzNV0g7QbGhXlmAiNLgSTpuuE5ToKINR2+FuaE5Ob/sMRv0B6eqMEEIfSHvKX6AOq
8HkKJGna37TvhiCZ89jwsQ1vpp6E5E6yh6Ekir4nqd3iWg2AAT4ir1Lj/sN1PQuLVYEG3FG0EWul
Po2iPMW5RBc43TXZMFTgoadOP2QwEZfegepTvuYPWYuKvQGfFShnT2cyOBOlyrZeX3eIiOxQ6zqm
VosIqnKLQ3lqstw5+dVQqtyyQQdTB5kz0Jd6ebIqn46eA3YbSZ8dBaFVhk5nZ1iGme56/KjhIgfe
XC0XSNYr1d+jR40SVBvGTKPMQFlx10U5glMFPmZ2bUlrTN06cDmt27p9iJwVkjNf/3YYxfvn58fz
aqbJZNdSKi8uCpFZY1kEV1ydXbzJKtE8c0Q7nyKmDEqRRJ6Ro6ERV+dIuaNdQ0d1/lr/uVv2mXrw
MWw3sX68cYeoSwu6tw7SbUzKbW+76Ff3glcg7SgVUFM9hgJFnVOoA6me67vNXpG0ao8J4GuNyO1P
dl7/VZdqpzEVUO0wo7agVl8aBMyAma6SLXtbUoo4xKSX911HcOeS7kAhDT9hk9aPOcZBtF1W+XdG
IguQIhEg0FXisvv6CHUqLi9GPu6ENakWKe2qs4BDGtbO0J6pIuEwR6KwYRCuyo0MsTCLaLLYgRlS
O0Vrpu3GGKzzNlzYLN7RlBC1IB0SQm1mHKfTxde5YW+kg0ftIOxwAdc8z3Tu7tu/gJBOiY0GAHyV
GyQ41CIcBiCzkQOOSbJngmbflvbKJnCvfwYZ8wGyGUz7uMpgi1XztlFomaEeCw1zrL+3W1eiiq3z
rq4PfPPQl7TK9VCaDmnb5iq0R3/wQvJd7HWKHcRwQSDt1o8bUnaoMFnmmVXrmDdeThrVHfY7jUJR
D0I+iov9Ords83LxjdzLBQgyART0zwdX4/S6v3I1eViVCfBI58l0x2lGfivNatS/TTDAdl3VMQpE
gm0sc763QO4crskphHjT2pKqoI3jZdG++yieDwXkEJIbJsVA4atBJgps77sWgppEBXLxt/VTQvcw
Fu+n4iSFi70i/CcBLhjN5Rw2D6NW2koQwHZ31XizkdHCiUQj1ctstxJ3MYTsn1P2gdI63yugHeBq
jd636EIC1mI/c/Yr1TOc6FlpSZpTgMJxhnjyr8EIGYtlG4pzM9jTeUfskZ/8PPv8EGB5+0BOOnMI
DM4elGSuqeKwAye15KB7GVwiQP77F8TEIq5nYTFyVabul3PsS+IfDBsedZaS4pvZSuBFcdDU1nWW
DdfhQ4mOKwwOBzoyS7jZuxy040BCqF/b2pvVuHf3YE4gXHpAv/KQfQh8Rw67KsLoBEzhdRFUIMkP
sDIkUbPP12YCxSVjo6wXcCJMO7bI0vRKDT5G+a49Ny/kY1R78IokC/4dIWO+KxEguEAq3RDiZIqj
hhJf6xdZtZINbi6Cd9SlZy4Z0Qgrm3HvlnnbVG62kRGCj71JUu1ZXes7Qi3+WL2r+sAPQoIWDADr
GTu/5CIWVa+wVbqpkB75o8KdCVpOQzNmVp3v7T0pa6CJHUECjUW045trAS3G9E+MwR8aHX5nqf7d
wjoB3P+W5ZUF8TtvjNFdsGWlwzgGCHPKRPAlp6Cqx/gl3CygmIh32zFpoRN3RvHt2diszBp+VDuS
J5RmmarAlmvHt/haQpNtdQECbFBRPHIrdxF0IRRdV9NeMKmydo03mDIjknIMsWDXSw0SfD//N+e6
tMHJ0dyB3Ocrxr9Fca5WtyRSrdLgSvcULtgB80+XQCnbndthwHQfj8Quy/lcf6ZvS903rSPGROZp
JlDVN0/SSVY9M9ggqjsn/MQeNx97e0Myc9u8CqsdjoaQtD/ABGW4muCeLRQXuLJPi+0nPj8wfbpv
QxSnaahosSTU3jaKEbhybKIxz2mXfWnaRHDEvyizGBa3WUBdkCyrckiH27a3qAeKzhVIs2dJTpWc
TOjeTw3ySJ7MJ5zATJxaf7AH67k64Efz1B0bWrxNyaoMh6sj6rpnIGlRGFVj0GlbXZDls5xT0ykR
rvrb0cCGx0V+WB5YyXHSOTS2mnWCG7cveTpUhnQF9/BQqMw+yTFB8FQXpZkbK1IrWW0NBD4ugFJc
hBWzrL7I6XQJbd2dkAVX9RHHq2iuYZX6LzGlVgd0WfXpMUpPZiT93LAmU7K4MGQb/4CwigvHlqMK
vOomPhCn2LsK3JBEB7FYGahe8JXA+s31jiO11LSix2PbsphuHYVLdH58ZCRQJB4bgdLH56GWf9aj
LP9YbCMOeFFqvVWphpISl2pzgn4UKhbCVgnOdnuQNG/XkVHaklmymxmgIpqz7A6TFpBaglx/ifqg
X57tsgo6OL+Pq+3TqHwpXzN1Jj9z8zzpB2kci3FwJrMtCqLvIiXzt2IxFOefPwsOy2tEL05MY5w7
d4Fj+15Ol2dnEUs88esF0FEmcieA3o4deKR7OsV6ukpbM9QGl45W6ktttMZLIwlOqjkLtCOTo0bR
4q7Gv6Wyvo11XB2JoMQzY/F6jcnDIaJiGYho5EypJMwtrfIKYUhX8Vyb63sE1Zmvkyqis69N4LBO
TunoWVZmsgZcRSXpumop2M7qi30S1nvP+r6/+Cj0BCsoj54RQ7L2LGyo3MnJnt892c+yBazqm8tM
JXjrdbWj4SlRTZKtCGJSUJikhoOXt4cPYQuMQkJtTt6/4+NnQvn1usVFqeuF4EgopCvJmNN6I92j
PlzUK+owmQ6LmHWzYiEMcu/v9EuIfpLrVUKpZyNxM6W7PLbXq4GMjsfR5LucxbVLv9szEFhLqdoU
0esiq+dLoiLRBJ+mkZpkj5RT44WvyW/msTcLOr1Rt7qVcdNnGZPiQMMS/9TkVap1MT8UPU97FZ3w
0gkv02RIQ6cWqUZyHYid0X7YGbYvwqQUgGIR9+Vtuu/7SxvxPAkwwvF0QlzPL+xgsXRCGHQKfM06
f2RlmatLYsF/ADVFG/sNGBFRFbNM/l+hye4PBsIab54j6ifWdPwwB3li9TkccIhv6W3D94tkbtW2
GEwbt3Ym4ksyyd7K2l6yzfi5ytG7ZuIfHt8vaTYdJFvgQenBw/LDdeQ3apSIeo6m6uN7ZAuXJKbJ
GYtnpvzeNEhjsRyngn+T7WEOnoSFyf9mdKPGRXkxEbq2YZzZEeWMaSQJtfb+1VmXsvV9EjpLDhCI
svKfsqEY+vJx7dOAeicqACdxus//dMV7teS9cob3WMHYDYVGa+amoaH/5L+PbYXt1b/Qs5tGkGKm
ydHQDxHzmV+OmYXR7eO4qGj5j2hrLbKayiM2WlLPh3iaNOqr2OJZ0AOu/blNGDJH42rNROGea3Fo
lr9eCGIGj85O1BFj+WObddATzaKWCvyKcjKUexRwpjmRbJZCsBUfwlMxCFiWQv00zQyfb3oJPkaz
mYeGGXgve47u7eMRYhadfE0yLqIVA4r/BhklYjve8qdB6lvjozm2jtmEPaf55sl+GEXJOn+0GA0F
L5h4VUNIfdTGdvht+eHYnvGKao3Zl/99e61fd6gPgtyeHh0aMtsC2AG5ugoJ9bBx29N5qtXi3qYN
vZbAuAsi37oOS3okvzhJyZVptyWLsJYv/oq9qurSvBeX4mfkTPhAXtUB+SxmJV/tM+dlHNUCjF1V
mbzEPCUhy/iwNgih9jT+ociXap8QetVuUhAeVHDsRwYja7pEB6QKGa6pPmelSrodfX+rL4jq80aQ
F/dy5Kl7NDBUNNfGdM5GGztY6RVcavKv0MSlDrJ2QHJCb0KRX2FVs9tyE3eUVlAbOU0O7x8CmrC/
sMENloHnZnD1q2fzZvHaHj8j2VVJdlHVFAHGmEnn1v2WhCUqyGY8VoQm7D5j8Mu4/oWHvdJ+nDJw
iEUlemCWnR3bXe6vxtJOI3CoZK9ZiULZyyz1o1CQ7N2bBNNyr5gH/nmEB7zs3HNCkiyt0b1eD60f
LWwEyfM+TDThcDWdy6zGVwQVZO+cfuz0dBNKKfpyHFteohRhQm+yUtavHEBkKGgSwTUAeykn9yrz
GJGJWq24XAT8NsRBKcJA2KNEUUyBNY9fwwB8IEv6PeehJ1R9P/Xoume/Gys2E7+BUVLBoCmGP7NW
bBukDwjI9TYQZvLe+I3wv4BhEl4sIjeqdliGNG9LA4mZTBei5nR9jr0BfGb3bq5H84bgR3rjwkeJ
zK5QRpt0FVpmSg9lUMR6Gn+7xi9H2aF7upeZiAAhNvHQlxq5jCCJf17BQNx9bTZ451iZ9jUBgMUm
MNgP9Fu3I2yrH1NbwJ34Cd0UH8PP/TVPj9PMWdTlJ3ahEs5/ZsG9MG3fTTkPjwpguqwUvTx7H4GP
KsmZPVveUOoMMWZjVipjv0W3nKIJPdmJRxKIgceAUx2XhK3oU6fL58wV3/NLSklzdwdZmbC/gts0
sqIk20IZzWTXVXP0up7ObseGJjxQUtKa1nqDnyzBzKEu0wl7mFzjH7s/vVdP9NwwYBiD35Hbv88D
HBKubUJZ7jP1uCTb+Ic+v/3Y2cgS+t10PaLyg2PL/VZa1DuAJ1ojFyhcWAyfNB2NE9SHd2mKnECm
43syVUSIqLzOpzOWkpJULpXbGkircQo0SW0V0aSxcCu1b72d1xM0YAryZ4wwvT9YGDNu6t6T+864
f3+UrbfSqRg+3YZ+dh0ykNWsYfxDP6AkTYi5aDOoPZQqYiMjLUtK9HfbzT3r+UesPDy3cm4KFfGY
NofQq8mCHibJwOimlwecyco+qTl1iPxccDgQy+JmQEOoiZ2X09jC9M6TDLKssUoJGzbnjWLfO1jL
9JxhsX72DPUPROJycpNt1hQdHjcln5j6tKLOfgHB4yju4M2Ncj9YJxsUbQ8vpBSP18y3vSOpQm78
5RYDLmyF1m1xFeNd3tUCOmzFnUYl3zykoTFoDYJDIYyjC0QxUKg25mQ7dtJJ7V4dQH4y/QYNcsPg
dqKMeGz4AZ4cdgcdMQUvXbem+R2hhZKkBg8bx0K9gaxJmtBTozGkUYvF/FBFNSwyeWMHWn2Jh3hb
3WR+X1gXJdYBGcCID5XIVXmbMMCeM79JKenT1nJ5jERvHNTocqdnh9VyVYiD/g0NMc3mDGr7QkaP
uFcOpXeK2/IVR/UPlKRMmjW02UUtZKb4Ha6NwN5PlpSLKufrslk/sWerwllD+84l9jM9KsfOKAKj
3LQighjQOSo3bDqmcIdtqNH8+/JWVaBMU3n1t9knSH+XTfyNFIMY8wOD5W6bUgMCqwuXV9w6dv+O
r0Bho5if+g5FVNXiA9ql/taUKjhvZ8djumA+6daM2CkVDqnw2fOm+9ZSn8klm7xFFV5u6yKxAC0t
PTZBR+dy0jMGXqSYTazabvLwWYERKfd99Isu1mU0JY+Fh7bt902FP8NSD83D2dUH4lUksjMGbK2E
L3HTU3AUDJO/Ov3Id+sjgXFeoKKDbl1svTLKE2Zk9G0wLCxR1QEfs2E2WGZsKHskdXfye3xGvVbW
3/zJmUPL+DUDbHXexd/FjPbkE6aaLskTCPz8J6OeCiaJOZSMR1kWgGwPTkQSt9SoBdtSE6XrzW40
8UvbLm4AB0faHCeWwFHkywzXEp/CDlUGLK/FsvsSBZViN0dDDkwDSirfx6b5a16bbBn9EJphPxy7
eFqvNg7VXIZtSSM5hyhmgiJJufIArZ8Y+QxjmWhfMHQ+o4GzhYN+vGPdyhK7O3bn6Tv1PMzAowUb
CtU2nErNCen0x19VWLkEEJ2SKG1ho3+kBaHHvX0dXFgsFyC7rTjOuK0zAuxvYG7XCluwQVj+E/cE
MHK14ws8FN3Lj/ovJOqhWx3tYH6xdAaI39E0VweHcqAw1b7bBm5n7KoZdJlR/w67eUKoe4arg923
Ba7OQUE4xE4Eslkz8HZwHtPZEw/QWX7g+gQKOUHwiO3sWWfycJTxYEtcRZtkg3J53fdI2mq9gyUI
4xQw8b5ivUFHMSvgOTSrwDToj/zytywfzzQl8zNUAsC37zXRwQ8lLHXeiL30dwMXxrU/KCWnKjpC
kg7N85Pa/fCbc1wRrRIjX+7e21mQ+Xdr0xYZcvjV2LV1FNVZNnnV4wb4eeTWJD/bK13y7d/1OuNo
IbPxxeAdhGcVlyhZ7JDRfc1Rxb5xkIh+eEZhfJPZfyxHND6Fq7m8P2loKWLHfMvqNyCmAyS2CMze
As9w4dePjV98rK24cI0A+Bv/QThtLgOx6siSLHzOwWF6LB/jIZCNF6Q3NQDW1AVYtyIgeUh+5AB9
vQPtoOUEzpniM4up4Xs4eUsZvSFmvptqT+Y+4uvFBYoEIv+J6Xyh84L+6ohUxOGAKKCwfD93zc2B
IdD6oEJsxv+5gl+QZiVH9Hv6rUJE3BFc7YtMk8BFTkRVMJ8izUxwNxTJ9u1+5VOMG6DgiPvTxBy0
Zu5yLaWwokGRkvQtkBFdQvk94QGLsQFqpsAKBxCDkFu6OkLU87dGNHmHm4CMyCH6Yq+ou+NG3omU
o6W4K3nDkI+fGtotl3096TfwN9y1M49Ths2TeAJuGAyU2DbUrP/68W6YX9LQAtbweyjpbfQJGbDm
/poTAIiKt2OcA8762fKHsokcoL756Ij0wqghzvEKlOrxP5yIGd879EoPf2qaNzjp75mQNqY9ueTN
NQ8GbVD10Gd9izWGX8jVukt9SZBO81gomwgXu3yrqetbQYgXoL7FD5ye4UoXuTT1bDTx+f46Cn/a
9hYy/6qmA//wIn4qEzQS28SSq9hdbaOuxBitJN2BX3IcO100PYsU4u4ezLwrztK+iEWR3ipXZ172
1Q9pZMaGKVjOJFBWd6yWH7Ruz5xohFWQ01JIA9FRKQnXTU39Lw55uAm1RBVBZHZNHETQ/zOyUz3M
88d3dDOewHXfRh0d+xXW25YDkJQ5DgIaIfXMa0ns9Jm1Fj3EO4/34as5JOasIkewd2TPqWDTIEBp
l8kWJ5BOrLYkkT+RT96r6lTYE5G2TIzyRM18WkRKtK/m1oI0P9DjX1936iBnQczpDmTw+l9LNyZb
3WwzALW6Ii2k4hROQ4VxMGO+N4CFeubbn+1eMo6E8BERHt7vw5jaKuyhCgPqy/LTKDWzOauirKwm
owfZ0bfE3puzVBeX7YAI2oPxEbNLQGZMCG3uF4l8SbGaJJEGtoM5Bvdf6d9gv2zDwoePU2kwN5bN
ee60QpasxG8FOJUkMJwLEbpOJyzDRE+m0iY5/1Wh6/2OwAsozfSxjaU8jRL5eRM4dAPjKZaHGT7O
EpeW5Q5UEOFX+o42zpSoPfA9PptPTpjkAeWFrbCJgMLKRgtewcTbYHsvBBk9AdjmXLWd38wWgkHz
tUcTr9nKQcUNYk7Lb/VqjAyPAfqQSVwADCQBJuadSfBwN0bmEfqb1hBvoL3SWfDZvAO1JQ7BCr6d
oG1DdbO4NM3Ka0Z5dJ2NI/wDj58yO7RYVUoato5F5ZVFF8TBJmAIbklKYNN0q3DdhZTgJkYFHl9R
CW6ZP9Tuqq6rT7utvT0qLInYkQSQBvWmnofPPoWURKtheJZixBPExivpANrmE5iDOFSq/9wiit0B
aHMHMBAi7oj0AsDJHRDAiziIz1hDq96kHfe8nIKN5zP74S03UDkmN+rHQxniHui4/2ILnrsdz477
kKDy+9Qto+1S2tTvSTSQjwhZxI+KIKW5GrcPaulUvxqVbro5aNTPvUnxBrIOSW3fXjkbB7O7wzHD
Y7t/hLBL+ibOgGWMWUt0YBgHJHDc9Hj4JCm8HY0d3sScY6Icqcb9Pxr7nCMAqCVL6F+2aNVE+UqR
W33v0zGWy7h/SQ+MkkRhUofaD0RHYGye4T9Qrcqppuf8k4dUJVaieK5/J+KYbCaD42JjnAie91TC
1FFM+6pannBSUDS6MbhlXZ21Jp8ub8pe9oUcUxFb7wJVOZJpSh0Vpe+VnmknJD3kWRcyZeoNUO0Z
B9yiEARKdBAXfGreSyIw6cMenXFZfkNapqi4n4a0CbExDDoYag5GaBjvaBZzru+FPj05DOM8XibP
u/YqVjx3aC776mAbikd4vY3DgLdPS9U5OVM0Awfq7O0afrxcI8KkUArDZGpwez5YVyfa6xs4q/aF
x2khiz5f3eWvOmiIb4MXCU7NKmNOGA4IyA4T+ZjGjGTCy2i0acjRCFiy09TezTdT32xVdIzV9r3J
SM2H8tlVqmh0qyaQP8TV6X74jbhYkAensiCI+tf6PmMYW4YQUg7nwFIxPJRCzHok3BzBowRT8+DY
rMDhhHL43fkp4NqROSk+SPKBQQIOdObTkpKIXwfFeDaiq9pmF89uayvmo1OsfQSRvlFn10nd2V+E
i+cIUGSoUHf4uIxThs5z1T58hlZVtaVNhrf3VUzYmZjOazqWBeJlvd+PUuHnTweqW+riJbQTTz5g
HK5oXfTrE4flNaL9VLRzVIf70WoHp4ewrGQWa/fsFsXcpOODxw4s/QJGECvIs/eqTrvZEWrN5Hhr
gVsROugfsSvka0bT5ICWuFw7JRl0mgmuFj5tqPvrZLa4w1K2nq56QwsbDSdAKzFgqoVfmgYHBoJ0
bUWyrSxFdQwDnsaGp7Aj+kdLpjwFxeIulxHLDFwIiZqAR5xHvlYVH/Xgxo8BPdqn2rKhmokA3A9y
A4xqRA34738SNZhenGviKW61v5vnkBYNlV/vkxf32+vcRfApHiaaRPphhNF8LZ0ZRjnvZb2pDHd0
R7Y5Vw38M/cnqS8vISPHI6yLLsvIMSksAjSbTGd5ItM8OpkFpJzVURzDHsvGJBDO+dvBB81EiWxn
elkxpw1dt0/wbnmUw+L4dYQuVTWnjYqe7Gxi97da5NTcJ+kRDAIXtILn5kNxaPL2JyovCU8+JNYz
aqyx5m+DiJN94QLbbZpUvffR+3iKX+vhg/HOskgnBgLTKhnofMjrMvk14ne6TI2KFwPZwsPs2LUG
VRlDh0zJSUCaWgjArXp+dZHq1L5eowAUjwzOBzkD0QN60wYW1kGQMlxKHAWLwYXlAccuh9G5PtqT
MQhDVkdGfuviaPOzufxOrTMJvm+plLk3XX9GDYtvPB6AQdEMDkGoFpBrQXOHmIRhYbkLd2hg5ilw
9o9j3KFxOoen6s9DI5fGbnc48EUAv/PgLZljZrBJnkDj+S3bpzCmt01MN6RL9+kc0guPYOtfFA7w
YPaAmZoGh1o4EzjT68eubF+z21wNMhdUoavslUuYKSTGJyqAzaBEIk4HDSGvojkAsyqGF94oQwY5
sucRtxYmlC134Hfg84LddqeU3oMDZXJr/cSYY7nsbsPya0SSI74PTedNF6oPe+cXN53HBHGdc6dP
EcAKbwQIde8UZP9be5qOoqa8HWUM8p/r2HqBY4yodxCFuJWQyJ8V64kPeULNHBg0ZMK5DWggdiQz
ITgjVcVReynRInH9CSOfTZPieqPTM0iKvv3/ffPmUii4gtq67cu3hjPjwwTFthpRJ01+amHAwNNJ
ylTw1YYwGh/QRHGmD8ZQ/ykof8UqB+EYTvti+jna/0p5PtTNB021pUzAaCU+pz7TJZVQ9MYwFINN
Vb4Xq/3O0YoTvyOJpDVq4ZEZpCrqkeNxaXTObi6B0tr6Ycv4OBJ+HGM5OJURH3DS8cghku/YS0fu
V1NY+ZQaXLiCuc0BIBORqcyetMYHogn4UAe/8P/G5YDPvEZ5PscIF2+CQMRrseOfq2+U3EuYWw05
yxh3IENoS3D3eczrGBKIODVi64edobu1oY8TjgwgNpMt2oW30zBy2kP/bZc7bRf2UFOGXk45BYcp
Mbrf+DUWSq3KcsXIUI7CaSi2fNhvXhhFi9Z/ynXLffMCb9FMpXVOSJMkDAo/p4ZfaZngyYG3ugMY
7YiTHKutlGIHoPKDv7TmcAKeU8yMwKlhz9Dobvsl3pI27afeKTZZa7pMmvj3+8FAiCuq05LZhv4I
hkHwkKXdAbtx5V3B/ITS/v3gUrUxf/ZHVg0Wc7+jLVodlFtzo0tpk7CekcruzwlxnzfPGe1z94IZ
/QtTkXfUdFz8rg3u7j+HmaM2UOFx4cOLqIfaadlTNalPImZAblA0vm4QqmjtUREibJOraBFIT/cH
Udtt9tk72pFAsmYuIuhgwLiN4CqZMvAG22/ADCe3qp+6rvAkag1P9yZd8z6seG6V90zAHmIj7yND
HF321Zjb5z/S/yzIvk3sNi0fESweuFoUaNcl+cgJwskewdjQuUTTsfl1g48cH/byDwtS7s8ZWwaG
PBGmwDfwyS6JeUjb96sKMflKFf/KQCrfc4CDHfNaM+AoOi7vOWHWcbfZ4B4rzF1WBfziePD8IWEX
FI60zQncCfWEmI93liKHWFL7wnnZYs+ohlIRVHVJiGniy9NJHmlQdDI8rmHV1VZW0ozplOFO4Ch1
67kRODte619mJDr36qk2yj7JmboSPvQk2SBzoaG/v/PVLxeiuwQIUkAB/fjejkI9lO9ux6nOS3ij
mLXXggDnGjJOYTdInoHhbTWNrRMQmfKXXMupKxJd6rMcTSLf3/XP3r+NVwzFL2LpnPFR1i52pN7Z
CImuKe+a58QfB13ZVEPQJ+/mzQI5TZokAJke80LNptI/r5jPXwo/2KDiYY6cb1p/AKBT8dJ0STnE
BehGtezc6Rka4rfc+iebFTLu0ixra8keMEWyqLOJOErdR1iWq8vjzGTwbHOERkj922rBeHX2oiYe
DvSDWVX0PFHdJzRf6ucXKJ/9nQhnFPMclj+mdxJ9dKglJAlrLi+pIChc0UJCkhWVOXULZ22wY3iX
xc2PW1HkpK5C3RzDEO9vvfjUjIVr9FbPYRJEb3yAN6RCDMiTycjis0p/Rj9mD1GEtyhORzGTGBw2
CAZRH1BF62W32A8gmVJIqf/Hp39iaT/Qicg9ADOUJvDTvzSE/jiroLTUDo3z3jL3YFloWtwyJXba
FlvSdtN0Gbj7p6sLz7PdQks+YyeJ3bfJCcLWGl3T78GGJ6e9oPc1TVC4x8hHl4zn0dOKLfgdaIgA
j84SArIvT6/LkwoxdZbgk4CZHDiUzOxh2Vbo0e6+OH2oChi4T4ldhro/0ZUgxP5AOOE8GbJ5JZM+
jOEkaXx9AScTB1sBfW+O5ZNQDaHllWZCDCm49ENB/x+A99W/qD/jL0zro3nlKhekSzgZ+2qDnsVa
e+dJn4MhtYC+7IaWWBivp8AincUpOriKcDyefq9Z+Dy0In4r3p+xzWQ/7vx+K+BXttXNQr/t7YK5
Tc/YLrweYLIpJiR9I3h160c7XLncU7ETl3XggTNuyYtQfGImmZBcwByN4eOqgjJOhFIlFkrMtNTX
aIRQR+rHf1PNkhpZTJqwDSbJ4I768AnLt+SztSP7nrGKq8L9qvqMcO36n+lLTshTxz6P36H4LXex
pZoWwBk8N24WI4B3V2W2e5LtAfQypwtIMIkLMD/NU8UG61I1KydE+cfsrrgBDPLVcmBtEzzc2d/u
DFYYAJiBo3SDyLVHEyzmhgKMkZzrbn8tt4TGzecc9T4tMR5709/SuikiWPaZz9362N8Mdpk6VLXJ
8v6ekANh8CkWYmpIy3rG8390aRNO4etl0FLiAsGlH/eQ2RDyiE9h4IaV1895SPgMzUFaN28OJ/xw
Fs3gr4I2YsjHc80lidHkn0F6nqRSMHfSpiq8DS7i0Ds8SLNTWR2ylajIycIp3VQBipDm0pdv8S/2
pcsw7di96MUttX3t8F7AI3II92NxlO44NDPJHj5iUxE+GnPMSdVzeJFfcvAAEUbeNOxY1FZ3Wtbz
2GN623xN3Kc+HjH5v6SKtn3WkBwXB2Dza2sdAYjoSK2I9fvq8yPDwCK22bWyn2gv5t/UrFVJWsW5
RR6o3gPJkIM87V9vIFMwqeG2R+IIk5YFs+glgVy0L4KA3DoI2IpVX7ZnyDKU4gXPyOSx3c3nS5mQ
do4oiRHM11UkmZXS/JMY8s8KCOIXpx7yXezQZac3L1LPHSg3Z09DrvHSWR8EpMuG1Fk3H9CWeZ/b
ugUzSSWCIm3YP6tP4Gl5Icr8arley7VC6KVVcln31/OyyTyLsnzHgO2IJUFo3IY8i8ykZXs25to1
iBFajVk7QIV8QHh7CXhAiVLCwIqm4m5rjF7xrICwt/5o4sglBoul0zXBO0In3XYhOrVbiSrnpnSn
KycNBhhCxqxdf8sfz9GQlgH7UpdkcQZsW+O5rNk4k7dpViLbj2QDQYImzASCI8VXFqphQwvbLto1
80zbK8fk3lG/Xvw3G3PObCsXtdFuZLClqsJ4fHoIhYmd+qAt0eavK/s1sJwXCyLaaT3+t6Id2Sts
lGOJGv+ZsIjF+ybLdwSPE8p/+FtS9kSEW8UBUDdM9x+hamMjI02TMFKEApHAGN0D40IBkyjO1mqW
bSJzJRoRnqZBw8DaQs5Z1JRUG4jdhBt3bLRy4Ilc8Jh2ER7bCIvNs7zEDDJWkQ+xW+cs1CnlhkoZ
bM8pBYmVRL2d+8Su+lAABGnPQypItQtg9yjVU4ILmCGmr59zxTkVywJPd2rr4Ghzcce80/zwwYfe
STldwRxzEAvtNnSKutd0yAyJlo8MYjyUyc+w5Rp//Ud2vLeWomAOTaVQd+Eb3qoH9d9dr+m5F+02
cw3WBJVPaFU0IJMpG8/+5foVsne2d79AXk51sCHk+UKh2CaWPRnLnOGn+vfhk0FebAenQBUpLn25
u1UodNE0qBKBScstLCx5vlD82o3rj/DqlnhoZ61k791J3kto29JezbzQu2DL03R8RXj8agaDKisA
Uf3AGHHv+5ypZOgc+0VZVEFcfNnWHgniQZswRRBpRPDN6l+kpwqsAkTHVgw7BJFq3lsPfcMO+9Bv
U/VMnuXNksAlGNGPgon7W3bFBPBgINJLXdDXXQH7XPY7xN6NZy+BGutm84LTHXbM3O0JD47NGppj
PGsfEMgRwX5demIGj4NQ726us04CtG0cxCFyLnaitpn2lLFZJ0JgGEhwZemUtD4fNJku31Mip/b3
xUeWJF1ScngUycOgQQEWaJEuVQ7sEpy4lZg3iWJ7VJ6dytpZgMgCRFXsFEsSlzoiWqu349SDFwkv
Wz22csF5r4QeO2w7i4J/BTS5wZ8xcON1KY4C/UlDcLxTcBVg70AhytOMXyZs4unYJZ81vraIPEh3
Ubt4zfz1dEblLcDFmIqkgxihNcVTumMvbRjpIEhuoyEz1/TrXrb4CfbOqgTf/rl+Uh1L1o6iEm0P
J6Fft9lm4cN35nRFU+R6e4TTfYyEzMjXZ9dJa1lyM7GMQ8cIdLkhyud3jeEe9AqU2+xZqBrm6Pnj
dS0JZbQJkm0pf1KF07SpvEFGNPmwmV8QYB2WRr6Enoau1eVuEUtzMtyos9bIUZ+Xd24O+qiaJeuJ
LtjAKOZ61fRX6cv8gdj1bvCgxzpWFfixX1FMJancLU7h3Tlc0v8IxGp0GwY+oGLhT8/SGiyzzb0i
MTNxQ6pXNBaI8AhViJxCK+dGEBjRrUtAySpSAL20oeC0pxTK/mSLxAXARKjG58jXz8AIPz0LQvRy
+lR5Eqowdq4TF6Y9o7jIs5zR+namE76BJrd+k10ckn/UsSIr1gYQZjsV2Ni/9eqb0hhPEB+FqxvC
9ZRnOfyS9hzhxwKPnri3k/m1kVDZDD/EnG9a/8hYhzySEw/FChvp9pmOl9lFmIC6vTXVPHz3Sen4
4LY7jFcB+0EqVjLfdQk5WrRp1FrqJA/uSo2xmYY8l8ZmzTZCt2A33yUJHsKYQJsJnZgWTBXHNgvE
fslefyBWHXecnTv5kJlcYytROR7pktIsJCUqA10ofDYfiO/E9IdMzCWu4D8SkATdcJbNGrKfo1+c
HM0f+OvvLw+J9la2/N46s8DaKW0nFfGjPD00cXJeTH2grTizICpYUqhnMMh+wC+R21QdJSrWBy/V
13iYFo+YLvRXmgSVAJDbUU48T6LpQ2U4gDBXpsj0tvdtXSw3dN5jxzTmI3K2gilcBUFRjY10lrZM
CARTfz0uzJ4T28jBk/Nr4JYTXvVbDKFCGC0U31bShnp34ucLwvqEQFsCqB/qidtJS1sciGeq+rvX
NIzrHCaM5LIEL/IQ1+M+lsBNukMU5uD3h+j8sJi9fkfNVvTuiOznFtoS4aS2gSQ1cuXoXc+yO2On
pVFgWZtPFaHQW3oH8RhBRf3HjZq/TjzXarogiyauRcD7SF36Bo3Nx7l8YtMonpC3ND9UekFPYsKS
EJlvqAibaSJID01HapYWlQA6I26k7/I1iWNkgsiXJt+aozxwYgU9ClcdtX1QHFd4Q+fau2+YjCIE
ToxdYzFtuXgmxqDyF3obK1Uv4UqbbPuebQazbJH1K3UKJIwNVYwKM6F8Hidcij5rmQOHZoJCDnBV
I4L6BqWlRtgoyZUMb4PCsAKXbuWIDfFYJxGKtXRtGlOYAmOWsFJD3LjenRdBj7a2f4lp/GlR+Yd6
0grZ8ARbW0k+Lihfr5QA/SgjGxgSy9kGeHIeZT073te0B2a8vJZk9tWz9fLe3XcOJpNW1jESsNDl
TdEvaRELuT/sjzBW+yBhOBvAJ+oSAuIU4iNfzqhpghSdmueNFtEll0R2nRaaYGuOhThzvNDwoYqw
UdBTNB+mBRnNZa3BTd1jJ0U0QIk0IVDjWHwUudjzqEhy792Rbf4VHlA4GPs9+nb6FVe8UsvwBGfS
7nfooBwHpXmXdxbmp1+m3h9Am68gEodqNLTgGwkUgXkPgXx4b1JF0ATDMZJ+caTFJDjPLf3/eKXM
R2Gz96FB5IIiNN0Dd7eaVvcwBv/caOx31kJgV1cqzMv0mel/V7VBsV3U+z70gHw+9Wbe40xk/Lyw
iY8jX+PDWLu5AEfgcLsk5mOMAaW4hxJkW3bFOujrXiBh2et/KQuLuxLsBhGvMdJfg7zIe5i0XRK+
9qis8QqrCZWPLM3vOw8KM4XcK+1aVTALd0mKEIwWQ1Xsov4eSywj+OT9YQlSRuINh4QkdY9ytXme
FIxJ+kT5qqki8k7f9nk7eFl9jZtkyS5lDRYLt5D8mCqqOv5aQY7FU85PfCqbrhB2oYkHFHvf/ERB
X4DYFv1U6sseMfuUX+FOe+Ix6hrs9M6AIwkdxA/e05RaX87RSV/qjf7UvdCoc91ms3Nw4lD96hfe
Etw2afhhWr3FCS2Bti6p8sJZQnzUEZLof9AbozEZGxGSlShybqcBpSaglDcURl2Wq6GQT8QXaoQQ
eLTtQbMi2KtAKefBPNnXHcVUhlF6MYBTUgtirQucmN9c/Mut3oYEsYQjrSTYkHkMtYwQIRcBx7SK
48TboEOIQiwnxmWKgasxSuIgNFWh6Agfrr7shdVmhZddX0XS/16B6rbi5EMMCHdmIqLRIqc/rPkR
ch8+vx4zu+CXU9dqICSEImfI4kJUgqIf5+xjZjnshp8QHlv9le4bnh/YoKpfR7ROS2V8qsJFvS74
PCAZ7aKYAEBLIuSnj7l1ZbsfyqrpklX87+YXBCVAl3MTWAtU6vj15EStEKGSm8PGTCPGRn9qEn13
pZbDkZXB7DzyYyIVZpbwE3Ryi2Qa0uO4LCNr94/fW5fUJg0voyCS3a7gM/i5yqARjtpRbv0gQFN9
OBWVWTmaSuCIT3cmLtMwCPGj6LnjlRNr33j9Dsh2T1MnaFNhllwvywrqhzp7LUavzu4uZCPWfk/x
OgMcXpNAMOfpBmdqYV9tdBkpJ8iamMQn2Jzb0EpQ1iT5sK690XLZaw/YRR59xTjFaAFAyyrwwlUg
7qtHeQE3DNa0I1wwJ9sGIRwI42hLazqYve1lZOUFekCDf+1lcTHx6EQXXNZSJKuQG8u+tDTTu5do
w71jfPcACb0FadMRjxLjpui86I5DBgCk+dQC15DxUNI9hasnmX+adDNSy1IY6MqIOnp2nssGZjSq
HqxhhXfY6+P1DlKSKPjvpwf2JQ4J/RlXzmAFXl624XF+wPGMXMZIziqO4R+2HFPuAZsuuone/+vK
U/4PGJ3o+RaeicgwX/rMmDpEdJrbv4OUc7uPDYbIax1IYSkvvLtdf14R+d8N99WOtj+e5wraMRmr
xlCGS1tSX693IdpVBwy38KGC5QYvu//JSTZIcxj8eIB4fKd1q8WzcomWh/y1thyhL4JuJgIxf2mq
xjPBdbx11gVW6HD8aw1/eF68+7HXdzrMUtpoDgnbtye5JRZRni62aK5DFBmuiUdxDmxg0m5kRQwT
VQurKN7iOjjknOLlWXsoRwORWS7EoCe/lmiioY8v7tQtk1NuIW3rvUhaZ9T/Yx7RHUVw/ELoXjnO
y3ymtQTIN0pTTYdCO1sSZjScmXKFtS6uZAMpdVBtZZEUnboqQQrifbFI79IvkAEWyWiqsQNYvDXT
+zXc1BC3gkpnbNUxwwvm2zJdQSuHDMBbus4gSRtvL936k/5GzCE1KHZMYaMTUvIR/YdN/BGv/5UY
WO9fH1Wtl411lu4HlahbEn6hmsFxRSGJMgGmg09uW3/je26TCrY9MvPyLavXsKCkyOvHX5RI9+b2
KqWhaRwutbdkyrS/Y6CQVrMvyb1Hrj6x7ddd9pS/g4PRKTeEjCD/yiFcovTLV73O9NypRGASTqey
Q4ShLxeiJlavoRoa7c/kd826e14y48IEXgWlzpsQKFHrjoTjinXrkVYT6rKWkUSIq6FKbykJDh8x
ErWXddCW2I/0kSvWYHInXwGUjXw/Kw68mkZY2/IGwB1elmNqZVm9fMZjOwmFKtwqXN9xLY0i729R
VOmkPBcwoc5QCwT5gSrKemb6wcIZhSj/Juqbxmto8bhJu96a52U7pCsx3xy34spbi9K2gnteke8s
IFnlbR3gEx2e9z4/dNIC2zdUv1AxWamphHvMORMsH935ruLKORmgqERbtVyu26GzFUfC//Gc5sod
f3rdbApH1/cOy9R1W8bbF2Wyqnz1XMQqThPgPX+QZbKTQLUKyX/KzwSzNwuEyJbpoDxTCkbcgNIc
Yrs7Qt4WvtKIAHVPGBuuwErDwF5fi9JdiCqL6tlbBryo2BIaJu4oe5l3FDItmzHGXl0AL7n5wQDX
C7hzZgK8ZS2G8m7lXaf2WjkdypuQQ51/0oFViHcc7h8X7IXmO53Au/yS4fdEpDToYbjDZUI5fhKO
vgXN4Kk3wcOwblC/Nz8yRWX8KIUex4fjObmpdADZSZbDpXWOWB0U7G089NzS+TTHDETDmeIkt25w
tBiMI/Mex3988odc2H3IWLjEZYxCuPfvJ01UkdO+4q7PPMz5+st5mMCQme6n+4mDAxeE/Lw/JOJU
4jK50CUPPgwOkntB5gPCqipeL3tEETkKRaytOdmISaaz4te490+mZuR2yBqeQWQO/lfbEkle9rXt
WwwfIX7C61H72daxj+KfrdICG08Xwn2mEIL+oHOKaL6Ay8eW35qBRh+EIbivsdbdZJYDRzmWCz9M
Vs7OvBSN6eFxe61m0mqLBXG91Onvfe9zGBKEZyVS5fmGxEeaJL4z1Fjj8gccSoNYRgyj81FoQjJJ
+MRtTOXWRtaMa5Js0SvTu46Ag2FsYTV+HCIKEa/ikOq7JiOlRXwq2NFG6qHK1lFQOEdpVYCoykWA
qExqJLM7tFwjuhmlrXB15sDOChLUZdZ1zN4Kv7K9P3fuSTPdClv3jwZp4XhMV5rAIAHP/g3m+g+5
J1XaEBI62CyZrIIQj7Q0+inVtc2POQDlsOVWmbpTfin/cZeuY3N9slDNqT0rmEnzAUISkYA9F5VY
HKcFxXHeCtqexxeiA2QBklcifZXvGQ4EVgvuTq6Bt4qjBahUWrsKVWfwc5J7gH2cgoprgtoIQRf5
owZA6xycZBJcSB6zgayGuA3hMgscqvmOUrmWsfsyPr1PnAuJGOEX+Cvzf3ehWuLlb9UwbDxCYwDl
rnmQgGEjUx7LbTNY83Bz8K4bbXQIyTGL0Eb5WRQNPFYGQK/X7RIffTBQyvr7xe6DXIDTegIm4Gxv
wkRY09JYSSVZHeB+DLEiD9IYYpOGaUNGFQS5eKslaknQeoEvPQMxT8BmHqFLxTZquYNaGDGtp9f2
8kxuyCh+6V2eAWrEMNmlfKRWdaP3A6Ev9d806UNXN4Ezw7yM8AqBSrhWxsSoVEFrbQUJCCXd1tVf
yvB2HoIZrDB1Z+qYUVOL/O0V/pgU1PnTHFYNdBqgYSqgFI55mZPCi3QeeVglCNx2BSQ++knjXRI5
PZ+EU7JYORmvd9njzfYhQ8y3ZjEx11gt83LqYdM0MhHbAzuH7G2CCaQ+bk5745TRgzJfpERMWyLr
ROQsucXT+AJ3O5XG74ArissEWs+e/Zd0PJGJnfGyVEtKuK6DKf6Z2bQg9fFfSSpdmXEiTENyGwD4
RZh5s4VN73qFNDfU+rAn7qTFi7fabVBANk+A3p1zCWb713le5K1G8X3/mHR+tnoqtd3RLJnnK3Mx
afGyeMgOvUQDo/khe2zpo69/ek0dnAaTCQVKtd5Br6Xczb0+wL3eVI/CsykneNCCsxvBfT4XPt0L
O9cDQRqjBCl169IpAT/kv6iWv28RwqyUPvsn1HA/PcfgDzdi0JC3GM7oNYwg/PSFPmhoUjXM5nw4
RhtMnmyG2YZQqk5GmIjpitV6nwD3xCK9+Xb09NIRVuao5gmShXhaxulBVsC8VUDJUlkp2wwmSxKw
zDP8Y4NErsxBtdvQy/gb9mzvqTeOUBAhTaTSWm/JtDssIDYhYZKH8ijs1xbdnuXHUi2dYJxffwVA
xHM8GRe4/HfsWZRvJmVSPQzROnwlgustNSBzRJJ/UyiT3ZeAkgdpUa45vfPmYfT4pLrxPJDdP5os
3H7Vh2Hib3PPnyHX0H8TbkByZzL/3tIGOIGe+vShCMEYDck5Q5QgtomO8wRq6faG0qE8Me1WIPhb
9i1Rs2qPvf7vhypcRXKZET/+1fBv45EOwk80sL+HSWu2xQVugB5PU/jf7bE/Rh1rNn/lhCShOnWT
9mOq/pi8mf63TfOEgD6KaV7u8vaguOBdx9kMODSZQRkpvJZTDPriQq/fUYzenlXKw/U2iwMMYsZp
Zx6omqOOWLeymk7uDg9Akk0WsHomOsIOEIW5rWXlz3tzks+LznTYAdMf1fv42lIipMpOuOFp21YZ
T3Yqi4GIQp7EPYoc7+L6aNHCYfgVoccup4GEtw+sstEzDPhqHZ3I+ubpACU8jxxaQ1jCCXCumq1a
dDiajPEKEmrg38IDLMfD9bsJk0928EKfM15q1wcDIMzIvEuLBxl7xew9wI77GwDXSjChLm6pntM5
dFrYBjxTlHOMPWQl8oR0StDwrUJpGZoYiesD0Z+T77wxjztFqC9+9a3ntcFQrna3m+udDKCs3mwV
vnGSqWc9kQ5+5UK8gOJLpTcbJwwZqJEGkLjEtiYgWXSmgwYvaLV8QrwyyxV7Vz2xf/2tPtWLUKST
c9lC2pLZZzqwcO/U3j87xZhXBmYkoaN6ES+qfNY8wecyeBauQHWvx8GE1nYpbB1ivFYfPsDLImd6
dlMfTiA7znSD9W9OAHGf2vyEXl5IaLSzh/ulij3GGwtN4IyTmtEvdCne3HUbAuk7IZ9euFDIgzZA
72r8/I3LswEt88kzVbmKJFKbopOiISUSPcZQQMDfg04KsjhfupDQuP1p443M46Bb4Okb2MsjxSV6
L45crPJFppw7ln8RJUpFzWmZ/70s7j7bCB4ZV2e6UcRXkpwSl1WjpwyXLVT5kxedEZYuNIHT0j5U
dzJL3XloVOVuRqsn4liRmseym+hUSHWJ9buSpELP7XAzr54jhInjnzShDzeYZvE1RnMmu8UNu2bq
3T2off9gng7YEwHKnNH62xTUyKAi5SkVQuI7JwdlGih3kxOfwdMZ16mSIn3Gjjrzy/1ErVxc/CYK
oqT8qg/5praZh6F8386RDF0VhcMlnLBo4tD6/bR95+8RCHJJu/uEaT4D1wG+lSdV1rA8KRBJ/vsy
zluntyXCyi3EFnHo/a52EI26hc2FQFsYE7d2B1DV8U090AJ8kfdOR8p4fgIKtrYZjypZPnvhHffV
vCtCGLgeRkGwpGtRSc3lPjvKA+ZyKvxI8R7G7/pZRGQwWd/fYKtonebWSNYYRO/MJ84YMR2izH8s
bsHDXsBhz6tXoGAttT642Mk4MzUep8veqL4lmeLzNw3Txb9kIObPma1nJ4HlVhJojHO+7QjWH7Z+
NrjApUQMMf4A/Zx84QsUtdeud0SGUgKOF+J0vfn/7QwDDMYoQZiOLTGwfixBU8LZPlRccIWJ2/0E
KKyJ2AKu22SdJ633KymB3AVW/VL37vZuH9XgQqGIHDwxs7cWAyEBCGqaxhJhaJ6TLBZU2i9VCzVZ
s3NZcZEa18pgjxpWOEjUotcPL6sYsnyO15k80T3oougljNOiSshvKsbG+Sf8Zve0p4RFs5JtXsYD
rChvvOdmyHNE2tNZZSgTVDhcl6dFOlt8XoCz7hQ6jHjHXDrsheIcYvvC0/Nv8MTDLRar3O6uD60W
i2SuJXiJ97sla9lXwBlruxyxQh/lWOwqk3iopFnawMBnnADBXmEgXFgrLRrqb9wCDER2oRzoS1d8
ZeQN+wc4hPj0iw0V7W4o6IFVw699pmhkGxnecKqbGY9rfOHne/HcS65DJE7vZlKck6tFerk+2BUf
eHohtzukaIiH8WVm5lCu2h2F+3xRIRH/8cY5mqqQ5HM9K6ClILkshfsCj3y4ZtnVlLZyVtBBwUWA
+Svvm40ONZjMX15zhF1GK+qXASN3Zy24i9QE5UDwB1laPs+uGTmdqhKCCRjTqRiwt74tzlhmymdy
6yVTnj3WezfS8Biv3U/FawTpZQzrGexW71er69m2j2qRXPc2BO3Nr0yTalY9AkS7T7zV4oosWwP7
OlDSOKT41+sFLOkR0Pziul11RBrKHuw2P728obmECdmX1T7Qbt8P77gyF75/wgJrbzmU7/7Y0L11
s6rKuUZNXmkXeLPYYfwaZyzF9jJe0868kXcC/vRqseNB3mn+BxeUokZ8Xw0dWCY6tNSWzsZRaRZM
Y6rCHxswU/QiHP1bUJBRsr8kF46X3R/2HIS/YxyLu9tCHu65LsbpTh+A0cd+MoRxWSs96z7l7NjY
+urDfXdi6rz/MOq20L6h6icniPD5Zc9l6AAd9si8hYIINLFi0MI810uQqMkBEE3mQQ6Jr4DqEDtP
bpReUfvMszJVRaauFviOucwem+D6Ps5KthFMPu1tyZBmwrrnhRQV2OwZ9vk+nrXr/79UGWMIJwBc
+pNwiSbJHAGpBkyJShHfnvVlbD4ZMMifWuOVno6XOjFteCHuQWpLL3MulkAGHDC9K93MNOLO5VAV
tf5jhZUk0lGq0rhEDn8eTYVMO9bM/q4wUBxlguFACanrpN/jyKAjhKowdqPRp0B5/A5pG8DuV4Yj
SO/KP+w7gNSn3GeWVpMV/34Fk69kvIdJUmOX0SGP7V9SvInKFPIqrjgJGl3v4ZNIfY9Rh1qEpHWl
jU0ePh4gWK9WY1wmZ5qkYUIlnSSUWddzQ0AWpu3kh/grAVzWqkTOlbicj6XYHS9iLXwDnHcOkm6Y
x+IFPzwTEK0Z5JqhmNck/Tc1EfgjASRSkahfAV6h2FsLz6pHMFrcvDvQWn3iLBZsaDq648KIF0TJ
1N/poKH4ZKE4+rxFiyrBMSlA9fN5nHmhTjCHZgQNMyw9G+sltbHp2C//ixwnfX5GbZKlB1RRz1hX
iupRxNLgM65VHcjma90mFs5XjBhPmyk12qK80LaDgGM66I78hjOhkRM811kSiXumAECposIeWkrN
aHVaOBfW4GE4jkpfI/p+Xtc+cCV0/hVcuAcf+KfrTA2EPPpqr4A5PJXl5cOAqAGkR+n5cFFLxN7M
RayJBFiK+08sdqPu1755QYvOuJxXFvsOBH3W4qXcKU/+4f2/E3DyLvHw6ilrANvcFa2vU/Pe3BEG
jUPMDVZeQr5FtjT5zVx3NcNANjW9B8rng25AOLn7yVrbz69D9s5+7ZEftJOPc2mEo8YZwwbwo3RP
qlwLSAhuAs4Fto2y8U+8CZ9eAatrcguH0Vl/cd8g4nwbs1iTBNVEfvfedSQG2PaWk4GznkeBJIfp
ZTKjfEPYLem1mTPMzu4C4Rb4/b4z24eAXOHOZb6u6R3Bishzph5MuhB68uJga0wb2mec84ybz+pI
zUxvrX3IfhEhN+oxtKs81/Iy7EPzHRTyZ8M3TIyE5ZfbxtQECvy20JeCOFqd4psZlAa+bmM7aDmh
8ME14YchcnggaD3A0WutMYYvnvzlLv4mGuhX4nizpawbI+Ypjp+lXsBIrjB7eMgPJcN7lnjzbDYi
Kljn73lbF4mOY+61QcqwquEdRaRqCSrSfZIcTpk6bpJak9oZfmHlL1U3BnRVUyKzLiUqXw4oAeaO
Bm3mmksPOXLqriQN/furbAn4g0DIhgwEngl2cJiyvclANb2kicg4TdSLtpypIreicjFbl1nbz0CH
F95RdCuTw84zsMDKVZesA+ksnbSLaSWqU9YfKKXirrCKX0cyfuo7p+8P4Iip2u50uZaghPqzp8Cy
eSNP7JtFLB90AUwRELPVvbtSJbTPskKy1PlWlEiSDmRrYPJ6udTmupyJj6cuy8MLF3yDImpj0K/1
Y/b8zZIoyZ05+Br4JGuNCegwhWU2Slzf01rav59e0GYtm2WapRiw2JItimzuESoaF73fR4oCOobH
b2sOl5izlNvgoIomfUkDaUkgrkdfoqSpoJgcwDNt1JGBbxd4c6m6TfivLgpacVESSBFDIAYRcgXH
7gmQijtszdDTzy4pdUMHGnlevwh0ulTfmypoznMwkllsMlC8KIPvLlygifC6ksmlX70/5Mz1DfCS
t3JiNzyqExbrMIo3Y6BerBsk6DRBrNus4uswM1nYutnT7IDYpqpbsAUde7TfSIV0Ll3qk0iIusoz
LPck4r7tL3ZT2DKPo3yEr5wR7J+YB0xHbYQCpAEUHMEVAho3hyS3pj9jLn6M6qNRk5dbLTlDzW8x
zE3JzFqeWGrUq3oAaPkUmK0VqWgEtekSYNXNSHyPsBzXSepWzzJAcPiW4o/+FBSv8b41O7SoYHHF
VK6MZwi87MpSYhmB5SRyuHvwfOI/grVZj0/3QEJNC53qi2Q+CC6NY0+x5a1ROtt04gg90sh0t9PD
3q5XaxITTl4gjdHib3vi9ueywtU7h785tDFSFecj/qN9V5YKZT52oqltmUZkxsMTOxjvmA04MPuP
2Gq6s8aCT8pHPggh54ZJs1Hc6Cxsd6QeQ1B9Bf2urZbDHTbivVZg+u9/T8sXNPE30kTt1+8HnRka
+0i+XH1jkj4whDRfWFGZEckl2oCAHhktWjjNZhgXSypOmxjUUx/N078SK8ywPC2f16D9AN6g7f+R
L766kX2OAZM97cBJJBb5EfZek20MWhAwh+5+ResA50g0NZYVYx1hZC0qFTrOAUR0Tvrhwzf/84So
XIzO7EKbmGRLPwDXiTjiQdAw+HBb7yaE69WDmtiUp69QmKvy5GAwfWzKEslQcdu5pHNhij3xlES4
t92fwwDqgyzUV0bW3V479c3hXpjBu70/qQolAUUpsqdCLSGJSj4O35wHtrrTqgQgZdnn4EeloyHC
gzW3rrhESuAspfHkzcSJF7qEhilzctUIJFSu1ztXukdpjIL0MsYOPoSS/EdKfw6wOCMBiskCNn+K
F442PMyUWCKiYuzd83vieysbCrC2PY8ICnKUeZHmKxE3Wf3S6og8RtrfSddqC87zNEDCvQF3irO+
bgrGO7dIw8/cNIJWPVTb3ho/bCP9StJCF65SKqA+Dktc4E55XoQABfXCONArVBYwr2rfqaHdGLDt
lu2qN53I44/J1Jjk1yr+0AxotU5XRDaRyt4Pg3RUsirF8wcfMs7v4Ak116VvIKh5jCdkWJayovIr
DqO8QPwb0ptK7tIK0rY89yUlgjCk6UkQU3JMwT2yHJv3S03jE7BsI7oRErUOFRkIIS1PrLIpNtlF
fwfJEwZYa+pUy+cZtf+9GXKZx+tb1KvW45Xw6dppzYbIlBw2E2A8tOeZXIGlTT7rxgYrbD/IoWEw
pSUeW/Nnep17Kpmqqdmn7Z5truYjvWuVFiz8cxT6OO4R75ju4Wlw5Wwh/OtgI0BGcXuIYyK6bmvD
iLO2UENCZaDvvH7hOz5HCW/eWSjI5GYRlk+NbGfNZz//0xqF29u3YMmO/nnvSyF7L3wDwb5K7jZO
Y2BmYevFC+JLAfgCgLKphdvcvwfhWDmpzWwL5yrzHxyRqj2TPNDc4G5j3tA923XyFAwKxy95OAOP
EUl3HrAdcufY6Q3JMlfLuKbRhjq5QzxJ4eXXkcDuCz20GoLa0R38MlU+B7p85NnIMm5y0XdhE68Q
gMpZ5M4yD3a0yx3yI1kO6sPb7lGa2pAYLpfqs73999JGn96L3HInBfQ6WhoNhOYmLo4FG9zsIHRX
SA4URGtMqC4Yj47yBQCvkX+igdULIFHggS+2VkUiTaAnjqckBUiSv+CALfEkZt5uyEAzKVmIN6nS
9xVVL3WC74PQVnjj/JTBcgj8TuCJ1A/BIc5V8tAl8JiMF+JAGEmN0PqsYLsOrw/93J7plNp8Mny7
H/JZbRrQf43inYE1OpRuqaGDGuscCjz+PNrWVkM38f9ntWjPTpA2QfW1oy6KU9amHTIZeS9LNRYz
7X9zKXrcYOW1PcytcdHXOs40cbZ0RX3QLidfp+sw1R/YRropF02r12kqKGhewZaW0kdmdcGYyBRG
LA3y759eVDi5g08sFV6+OFhQfktRCIKFG2AcdxkBy0WmDZ/5cBeT1521riL6akGH4RTObCidlsfS
6+DQSEK1Cvos7cO+c+ffjdBxE6pbkHgVMJQc5PSUAu0ZFSMYCaK/eAK9+uQyIw6uTlSmsca3qKrn
pKEenfxJTMisQZzqzKk6Ej5h5UGxE0IFyrTe4qHFZwHUcTLAiMyzoSRSupGmGtoLgCpYv/YzjGdK
6FNfllYjdBBPCsgdv+NEkGSX+roAPoxZ9mlClplCG0HGNaE+kQCkkO3a3eGkURjerNfn0ZUIkJJT
Pt/1rQxba1+/iRENHBH3SjQE1n0AKrhW1rUW0QVgjUCBhVn0AImaHp6MI+YdVKLU3tSK1Wib4x+D
WqpASFkYBibUCXR6ZQkZVLtrguxggwyXPH2efciEqbBMUeByT0G5Z3nq3qvxF1fB+9OR9gyte7hg
6PqCjGVa1VYKVu6KsTYFkWo0ScaqFTwBWbM9g034vigdb6ZBbOqQVW8P35e1/+2A+s1cx01yRCXY
sA+/2JQtWJ/QgC8FaWWq/YwOpC/zTP0SmIrIEbgwxdx4/gvRXUa72vRt2VUpdQb6pfy1jOFF18ya
KSx17HzD/N1IJP0Uir7KwopYSel/BCM6Qi7jRqBQIM/uzrabgbQ7jtHqlc2L0of6vNOfYUA522Cg
Eg7HBEP32jqsqkJ/QcRlg+VwJgNgXsZoUOgKG7hyXqikfy7PhpdLMoR95wh4ckFyO8YffvpzP4LZ
3LbS2G0v/GlZM9oCiPN0wyyZagAtAoCDaKMxYXkSDXJZYoimcMH2rUrlypqFGcRL7b4oI/wbMylo
5vxqJxX6+5mxI0U8pEWjGS7Vt0tqQ9Hs5EF4/xblI5o2t+x3Kz/vsXK3xchd8iN2KLoILTx1Ws+G
ArH/2IFbDzkIoeCUgjXSeU80tROjDbemGR+bhWr0kYjSA6F11LflbG2wLvAkhva8QwI69vzrgNjR
pqMuhL4BCiyMMYhpVk5gR5LbrXzadZY0tIk/wi8a5TXkdvXrEDPjLoGf/F8g1/NW5THN4w4H+qKQ
c7WNsqaXvAI7vdnlZjAgCamLlBC596WVV7Dgg9w9tVYTzJAZi6X1EW4PdcZcjo64bRuWbaAW09yO
+nzjcDXZMB52DWcuEYm25QgWw9lMF2PcKcOyzUkMPZqRumOidlKrA6N8NyygMGdOUjAsaHHYPuAl
h+r987abA4EFXhiqBIX7oCZK5Qpqm9smPE7e19Xa0SgA8aO7DGv8fhIyDLstmtm1/6Ckvk1+2QXS
E7aVscsA886JUufr+UhjepbGkeX9OZn0UXOLpp0xhOco5wjlgV8mcWjL6zKpWUQv7aKVZwwb1294
ZLvNp7SEOOSadL2bl1nXpBs6d/2pWJQB0RYIehpBqpvh5/QBWxPUMwedsAW1ftLB1m0cmRS1aUTz
OE+g7L/vg5B30+FLpQdlcQxtsAe7OzF/OHzArdMyQAT3bEk77N/F7BA9TJXALyEwQK5t+S3xIBtg
+Pl1cDAz7TFv4ZcxAWnWBhCorhuj8JrhBXmrS8CmwtJz1FGcfzkKq097rdFVGTynGkMjr+8BRyIE
EtOKnCxURrP9Irj6ztq4ivHE1/8efNtPj8gqH9s72RT4JEwbNkvB2xTsTm2iPUYutYA7fu5Pdxpw
IACl3z5CNPMfuGmtqsIRidLxcbmd4lPelmuiD6KGkGQQiZTZx+QG4DcRECpXC799rkzUuPN2xA6q
sUJwXjrmU+x5dcRD9dUDFLKJKjXclB5hSsYqG/ITAHGduRy6Escq86+s7/iwyc1HXcSbEWZVMzTp
PvKrS/TTQlBozx5BeCnaZmCJ/pccHEy8r5QxYSuSV9vMPSCBlWoMMeXSDnPkqTWB/v1fsRLJEzSq
EFa1hV5/2yvS5iQ0TDdS2PbvcNRbrf0PoHZFkUkqMhtQLuurvyb49eSW/suFprbZrfq4qiHAWny2
Ipm4f2/oPt7y8S4g3WA9mW96L/+HFW2EiTgsHpcLfIQRJynqSYPKuVuo72CR6EHb7W0fYGkkEZIE
v1gBTa5KDIcTXk6tfsaVAeLAds0m4/d1yQAQhcoxmnKc4+3VdRiW7iyyVe4JC7Ao0Fj8+kHuot2C
DAcejBaKSSnqdiJcAPmPi70PCUt6fY9KdoyYwnFNMnEP/8CN8XgGbO2c/FfB3uBAXriYcLA1t2rE
/BjLIAUyieZtCT0mTlmdCdCh14UeWTRVGir+xfQgXhVu9m4aIsnuWPLCsA25Gm1pcbfCztR7j8ER
MVzTljRTE1BxRKoRtH1MjuHwsxCORMDLqLBD39ec+sNU1qVR+BDHvsS5F13z1srEj5zPicf2W6qh
gCc94mEOBmzjRtgKqRtHCxI4nsARVpqO2ignYzWwRrBh4SpUlm6h4UyR4a1XZm0VSlKMvMkS2DJ2
2M35C7sgdvGaOkTgSUAda2qmb6TaZMURjzB8umyIqwAJGy1gBS2Ao888IRY7K8H26vwC8TX47vhm
avf1zZMjsGzmiAdpRBSYxbvcOctw7PTUl68oJEbtXZZ43GGmBvVNokoIT9hoTb4D5V8cg3a9xlG9
Wk79QEyv6Q8xcfn4Aq3F8RMrq9XYtdDfZd+DBGnww5PcKmPArfeFCcBNJDAtax/fWqHNAJXJY46V
fDQgN95AEurcXz19V3dzXlCYmWPMAupfGO7tcqc4KtGS7cElrkN+LtJKYX6P46/PEWA+Bkd3aaBD
jzr+ofr29BaARmcs5395sjPmC74vnjL0blQdJhzlZkKJLzDoGn6AAT5hsCtijlj6TS7HN3HQcS/9
8biXUFnrGKMOG5UAE0gUOlpNO2//7dSkiVNztsNYOeGLmeL9hJPMpPEsDn7zTwJF0MlciYW874wk
Lyx1dN8+8QZzRd2b4cwIF5bRe9mDNBtNX1qCo+QhnpoVi+8CP77noyYZVTCzQpL8uD3lFXuOl4TS
QDk3mIC8ATtVbKg9+hJ515Tr655ABmU0BULQ54ncXB2V6MaBy379Nwzo+0YOg8/U/OnoiS4bDJUC
lSn+tF5Rig2pPPdkuzTYBUT6QqrbS2Py7rIVDwE2pkBkiHQrCy0AcGjts4WAQfqDMP9Lrb0dLy70
q2dImWWjylx3Edce3vzULCWdRQOTIoN2O9pcP53OF0Zir73m9y37jAD2yk+MRbA3gtR32bEFm45j
AbHyg727XZDHDE4vZQ92hqfCnxXYEV68AdJJZVBeio/KLFpw6jNz3jbYqTcWF8hXbI0dZNBL6OEP
SSuGI0xZeoP8F6O47Kt38hYmbWWoBBit9w1rH0wxk5FnYGKV95TAtWY5fFxZ9kgR+oQ+VsDrLXEh
vjDCf/RlkcoZ4TlECmP1hU59WuocDN9LOp59Ssb0R0sw87I6IxwhZkEF+BCSf8WXncoDym/euzdt
5qjoJwdXqNjFtVoo2Mkc4K8tKyYJWxsDTbPGpQEO9Jyb5Mit37UUcNdbb1HECzTR2C15cY6V/UQ9
jP/VMdlKzVtGdK3h2GYk1sZv8Oz1o0zBNlCexN5HtjK9OSwvtgPZCmh47akP6VFsULF40blQ/Bt6
AhH0KqMgbkgk+asKbNsL9+ghKeRIKEUse+POeycs2eOU7CG9ZL9SDW7/q0zXutp+X+1JIaO4kqCj
zfYz64RCVo87WBX457ffeR6kvtC3yXokB4ytZJjVfgT+VPjw2w7h1PEEa2Q2ePkUOB5Qvk7C884a
P1vupmUsLkFNNxr6SEir4XI088qUE2GJbiVA2j0Fu3DcWjf7na2gDD79FnYf7XMs1Xk/ilPTc5/i
X+giQk5cS6kEUV+LV0AAcS80WlEi/xe4BBrm4T8v+HSJFBUGmQ/n+Xo48xENMbCaDoyotpqjt2cB
LCirc+JIwT/nfLZRoAJS2buPVeMtrBBR1+NqEs23aPmyNbBWLl/oXRGbACR1v7595CzGf5HCoq8U
/oMKY4I3J4ZpXqSCuA8vi1jJqBXDEjdPCt2q6qZM4DqPZZ2Ht5bCcOrM1yVfNOew330RowKlQHHz
7fWobvVJfzLP4pqYhdwWy+u7LcaxuBrCcghc2dk7ABhKN4pIZmNmSD7T8D5NpD6i0qsORmAdBlMK
fTfjfLpOoGn12WH4UuA9yxDCXdO/KkYQkEmYrtFkHpxR4FZoHc6RnaF6NeQkA6b1ef/78M9Hvdk8
5+6oYDvE/ON61nmSvuBTdczny1Lp2SM8YVhq448BwTPEMC/Vb/bIXZSEh12ngOdEf86jiRxsWYJK
nnnCqmd9pa5f6QrzAxEIZUp4gNwQf0/rtArNGRDBGDyemm1B41QWGDc6REG+GLBqynWyrVjEsMPe
pkDT3DB/+N3yLoOQkVFLmDnk6gLIeI8DHb36G7fzUTJH3+BXSHiVqxX4Cn5zEgwUMGikJI0fWiMu
rsGjk9WRi4Qz7OnzN1vKinKIpbaw4nuKkouoAppn9HrKUb18xQnY+bFEicjJQd3SmkGWh6wT/DlM
aRPbsJGZL2W5ehdZUwrY9rvPvc43e+O1VkATsTfks42lu7EVJhsxgMt2snADnhuJMP6a1XVVp+zx
7HAxhNF/hwn0HimgAUoNGIkEkLfj6Pqfm75PQkacXnIi5x8x4cgrMQJuT3UmhAXxF0tn9OpdWjPC
Cp1P6sVeYNtul7BNqfcP6sNYsz8stN8EEwpcGRJ2a0SAAzFfJeMrJN3ubMARNk+9a6DXneChkz2a
QELhreLHpZDCMsMc2ZkKYMCjhazv+Rc7k8cpKLhlncHjAQNznajfuRm1SfTjOeFaf3GJmpcmtU26
IHPawJtbOn28KIYNQCFYNDDT1a8ztFZV8oYE3/3VkQ5zLf8zCKrcrXgdstFyjfUB8bqjSDgHwl6o
rzDUo2aH9l8q8j0JrITLML93MvgEjyfriW4PSGFBvXpK3QINt4CPCe5iZ43CYYWMDEzUxB0zuBMh
Et1eWTWT9jiQGUcwV9TgtWHH2nGVVQWHjJT3yEgxAXClt57p4+fEAGFu8UOxMWF0R41hc+RTY0/K
5eq+KGRZ4OoJBwPHy3Arhe/GB1heV7qO7iMORcKI11qEWLMAb0MeEHGLQiOMP7eCSkyiSH88Tdzb
/CbYsUlnZUIz3AUnTign4qIXNrIujlwVUQ6gTtz1CgkBPsrSkCqJJ5DSpzQgJTDH5z3J4QzemyJr
0/7ltxRVTANcfvZhSsKsnGdh+0JPwDC72jP6CyzjeV744x53ODAK8VQ+laOJ1R+vozLi9P/6SSUm
faU6WRKCNezS5/7stTCcvGUTAjGLUnIp/2p0XvEKPRX/FIS/h2eDycRGGCZipHu1EkWH4A5UhYe3
MB6wF4ed+zHdChLYFuj0NjA8sZxCJaIau3bw9Y8jQOkS2ZVcrjx8VomfvtlHvxM6azGUZXYJmPpa
6D0hP/M7SvnN+RETJ3HpA7AO31SFTRRuu+VqXMTMEVK6TIeMvPA36TirkFQXavwRqGok+uqmzKGU
6M4SibQsZj+AkCpoifydUufvKzZmNWxLow9g973uKxnAiBF3wJonGhRfQq5OSyUSgbu7aB9xHO3O
v5lqHoOyC6vQMqih8KUVDEIIq2QeF9X6zUBvdbD20LwdBNXzreKkMfqmf7NjuT/cO+IJFgoyfGl1
8svSPvEZJn3bMU4BEnUp43yjjt40vnMYUnpbBKX6RSKsqisam1JQmV7yJATTPiLHhl4ZNatiKf/6
cIWNZSZuETY67hxliYloNNpFHjEnLRcpLmY8+YHZp/5OTBFjxj20qrIcy9Hz3xdttYEM7lGu6QQM
XS3HrDGiJbCTtBA0EKQQCq2M4tp/AktSqUWLn6VNumbShBTPiuD3BPZHbq5TupPpsPpLeM9pC/hI
0fUtvmqtT+1PHolkQqAf4p8gH/+/p681jE5xEf5TNezLyy9YWS0PrOAOgBo+CATwyhHxTFh4/1QP
r+1C+dKVojtMyP1xZ5s3u4ZCllD3ifDSqRWWpZeV3axxqWcX2tGX9k27h0+G/Ukny8ZE6L29sNkN
pG7QUgYcfRd3fVUl7/SAVnnld8ipHYd4ExhQG9+kjt/5cqEnv0yHOzi1Gf0Eflh3hwMUduH6SSH9
aYGsA37u4Humi66Rs4lr0BJC/9NOPnvv9PrSQARszArjSinRaZ1Us2aiRjIV82pt4KFKoyMSImW0
CfOTJqfRFK7dr7Q5qZdqrVEk3kTpGM8j7+0Y8qyiJ9CQj+WNn8XLfMSv58FpSXdXCGIuEU7TkpOr
s91/Usx2SXYLzc88ObN0plV2EpvRFkMCV2V5+KF22yVkwTG3gEJoDwdHRYbkXSlq34UaCiWchPk6
zcTfY55oc2Iod75JYXme89OPapFjnJH3wHUZ1RL7jvI98A6jn3scEkAWRHWJz5GxxrIkbP52K3YF
0maKaJfQUz8CaTQMP8IkVulD1gN4Yduy3P6lZQLlpnO//bxol9pqtacTiEGgfxtEU+U+ePZyGPlv
tkXRqjECKM55biOxkmwD6jCauqGNlR+rHJRZLCkkHtUViS7H7CFpeUjJTeFnZXBIh5aPgjqOqKd4
7w8S1+KiW4Y4nfWw4mL90qW/PxgFoelsCEDrVIThRvtjStll4BH+Sv2Qi/4grI1QgcHVDZ52iIYp
/8xFOJDN1RqCgjtLsp+CdCQ86OhXNRzHhauI2n8QxbxrTJCqxsbFIimBvvr9r6I98NApV2qRlpUa
5+XIkBPCjlxPuMasQoaEkWH6rdEquhE1IBLuCJ0GQ6t8iMzFhhZ52nuicm2QHrQkuBKlmC5z3fCF
kkYA9YvTiyjgW0QvYe+VWjyZnzBHOzw+/eCSjCKvB2gW2wuXkXZG8G0FXsDnoqBkF8O0LFV3f8WA
C0y5/owevp8RRDLYk0+v+gkZX+sJnM37UAJWaJDFOjAMWTY4GgWAG20nkcbbn2XggNvMKIEFwVZG
aWj4SDPr+YTCe81d0wGR2zfJji1+BN7L8t4qZ06Ckpf9VAXKixSCDUy2QyJG6mCcax/ftukyFvHj
HBowjsum/PJCJpEN3nBiU101fMNkFaPEeKRlJ1/4Cv9wGMxP9Go0IdLNYIDQ2S4rIC8k/C5cj24c
ha3rGgy6DyCK78C2rsxZfAPildSzwjgnpg0me7CW9ZWKFkCRxzmpVCQEH0Ij0F04OnGY1Oe1hgoS
Lu3T+Ln9BOIeq4mNpeHQJJyaSM4p6E3X9UIb9JzymnOefrfm0wDzNd1h22mzGeuYkWVv2AF5iLZ4
WXFlnvcdOurgiigPvzTJtelUtoso+C0fq4qSVESSw/bAhs22KpnVU2vPa2kukH2ZMvzQro8lHsP0
0GtlQNuVu4D+4EiFlEzEaslG65lSnHvpeTVFeIdyMCebpEyou0fqlQPHnLDL1IVYqxGiSHjBfEqu
24Hxr9RCO7cLquERQvpBxuYLu2sHxQjoRz7BSbtdyM2M81ELX2ZaGbggmMbVnAucuXtkXF/bbGbn
JztgPHGSv4hHmu/lLhPPQBg40/wpPCGfJB/A4eEsfWLv5UxA8VogOWyUrRad9/vXJC2nqwjaOwiU
DXes4gzZwIYZch5hyeFRjyfnxAZnFp2ZaMqEQKrRGw7dFgM9uyX89ig9Zih85EqDS0QVQKqnNM/Z
fRTXcvUuBTxsiH43d+CvZNT4nKAxWmJlRDBQMTeCetuf9BDgq3bIdSBjLEV+qgybbfuGUW5atzzr
cn0AN+hkNphT7VDu814cLE1uHb3nf/KLnEqs0ie2KWKqdPnUG5M86Wu12l6/24gFdsIs94kfP6UY
7Itm/AHAYrl4zX8rVx1WXA4qGqmGYs5xwjemlAx9TKPyIrhqiR4PE0m6DJPxV8pyfXq1yIMA/XGD
S14x3VDmpYtSKhnXTP31G5G9yuqpGc/oBxy1JpMKuwp+B/WK8++8BG15B/Hb3YVg0R7kakzcKXE9
CMAJWHg/EqH9ZOBvrQLIOfyEC+YICVx7SF4x3PlVMLVT5Ff1/Ui56OHbny3FE95Khui4S7uFGyL8
yuMntpga0UnE6QCIiTh7NrKThBGepnqlOCuuM+ihfsB1lHk6AcZPLW3iCDI2X2doJSwQcSlB5czy
fFLFxfhetHBzjSfbYROGQPE9XF3psmuycJcx37+KKJnj4ea6QEAxo6tjhh7zdQW/rthpvuheyIxC
eEAL2It0U69U/5GfqhDdN01Ea4lxD7QOETtjAWahuLhJ5+bkf3sn0Bzp3N0MRheCosrFbxiyHDI0
sjmkNN5bUyajGeT8RlUwcAPxNUZeIU68rFRReX0H69R23xsC4292b6BbVTVSsKve8MtGKzs5x9k2
Udq5iLeqy0MceGnCoSlTzu0bkhIB3H+2MJsnEkJS6i+Q8ReE7LF5gkpbLapC9r2mmZ4ibWuHJdG3
7lax78RsrxnobKxAEs/zKT4r54n1/nZNRZM8AyWcdZsf24g5+VjhWQ9iPSV9Rgey6j86ruIuszE+
bk8zqiPW3mF2oyeCJ1Elk5CtbmNEi7jO0/Wssx9rFCH0TtN8CDWt13ELwHns7jFodzCmkdecpmpZ
uIkSqj92uS1rxdWTCgPg/6mKvWZ0aUh25atG4Iv3wdHIx2UFSZZXNMimsbjtO6a3XvxEtEVm2BRU
YT7yUOwKat+QdAAEgd35IK5MnEtNzSPD2CS/Ekee/v/ukAERc3zATKzVX8a7bkEbJcHUijK6pzCS
SY9eTKkNJYfRXq2V3GrkfVc6NR1m2fWSV9pn0KbcM/S31fBZuNvtMaFPx+9GYuWEViKFBniHAaOI
Y96IBA7vXb7H9qRQe8znaTY8nNlZnl34t03yi3wBtHfYcTXb3fz7KFmi6Q9voAEpSBjZfsYv5AH6
BDBcRUMumalItuuzv1wr/4UTTjX99sr1U1l/esEWCm9cJT5X+bz/mSwP8PlYGfi/P5BDv4JXfYgz
0XD2ZJLr3Lmo4mqDx4mMy/nv9ms2+VE3nPZFWd7BHA5YbBXU3nSDO9NA82XkTF7sktbu7hhJo0wI
YKlVbrC1sGy6RGWfAtPdF5fDc9e2dktUAsGkyb0hVt83vfLGY0BssGqW7PANo4coJMM04hjxMe92
LqZ96cL1huf9KAm8/33rX6fKnlToun2ISIDFZo47Yj87xUs86D5d8cyCJskdNVkzhE4YtXLyE8HE
+lZ1vL4z5slZGa0ZN1Q9XAaQNVMaErpRfkBq/BFuSWxtILLwNaXgyB78/6qDjX9Jow7KTA92UPy4
i0ihByBAMmt0dwyFSGgH7rU++E7UCMY5uADfAvuDCpHRL0tN3e/aFV2avEidfBCNVeJRvJGulhgR
KszbHIY6sez/tKDv60fI8DrQyC4UfKGddC6/WvD9O1X75MfW2K5OCUZTJK7mdU6ZUNS9abKjgA22
JtWwv0c8X/4SA3zohemfyVApi8BTYdeaZtdNHdIEA8PTRTJjAG2pClDj3sCDrmUFxz1AY5lOiZaM
JYC4J6R61JvoNMGk6n6NmI1XLEjV4m/1DNMQWZ9dGXNF43Xz37/RhKskuvttaVbpbGvJ060D4BEE
GGvoYKvpC49OCvNY33PiLJSJEeai8V3NxDMgJKYv2fkhPQamrpGOv6mt7Xs1N/eRv+tNGAJFbaBl
GaNQQkO/79o8vqoOGp91iEsMq3weBVUlv7zSVyc8veQIAI1CFFAq1pMm6r2Su2k4wtBCuwMHDN8s
wscpi5saPAWMSoyWqebGx4jr5QPLOXZEgVl59rbHlA493oCJoUV/27ao9tGMTL9mVdffUSMn/UK2
TEJOSFAXey+807LlgvDTchfF1NQ+GFtmjXIV15pfY5Bd5NuULnAmQmZTe8SbzdDpgTrKqj9YiGZj
cPorzg7ii+DNxmpl2DIalZYBqv1f1ZAHBcz3JC2ml85zcgnldYpvUyuN25AXZRHwULvrH74IZrNZ
2LSUWYe+OJi2cEE97XIel9tGd+kLtlzQ5uVMMY6YWKp3Urp0wrTwxXi1v8mFtpA6HFKfUajXiMBj
buy1/NwbmiwutVdWOfkbBCeO30S0ZjGaZc4I1aM+cLAYhdmfK1nYSZsouTSo4XadzWfof4L4Lm1i
9SwC5Bk2nfLQtD8cZhxR8rutOnCYQi+YyZTX9lJ6ZiP82N0zpx0M3Uh+XLA/0QQyBXvpMQkxqPcS
SPOi5vNO9ZgrxUDK3IsczISkC1lGY9DiL6tu0FRY34TVOeVlLVYjHWH29dG4M6KlJVGXN0FxcDe2
9Nvv8UOkVSM1yUp0BlnMlRUVWkNJJcGwqJzqsaryhnPaGy6OYdEGLV0aXPm0SA4hXxT/paU9P6HK
rTauDKgO7lzCXj135gTEtuoneCjQ0eEFBvdG3N11CfBtXRVia8YweOy3wq/SojXNnr4gyqVkCrfs
WQ4VX+wlKL2Hj/+g7AwxEAme2iZgACz9KxlRNMoCwfREZREcuLMn0AXu8/m05mMpEf6HXBfe7sIO
zdCkSClPLgAjzJzZuewWadXBFI7Cx3XOZgE5BtTjx6jJKOgPZyxmyEVyevsZU5tBfilxv/nc9aPS
SJxvkvMU/pAjONCf1gPDsH51g6woCpnN3YRWsScHK1TcCP5dJmSEmZculTiXy5L8e3hJY247ZHre
+M3Gx5SEyqPWU0ZCZOkWfD5Rk1FfmeIqlMbDnpM5mTkEukjbcWzAsuzW0g7RyIwLwxyYcMZzXMve
lWGCVv8P8+lReT+kqLEps+B8MGz9PWAqgveC+72VtqV21OVrL+SJmgmuKwpTod7RLhgdYLBxha1o
R5Flqa1OJ1KKnaWVlpponP3YYKwLUYKby52sAw87aoMjoDS1/lVj3V7G+jS10lpPnwrj3b+HBTee
+3jTDshMrIxyDsanrVCWbilnLuH9zq6nWysnNUz19nNVSoV9DMD9bbbSLIEsPyRGFEQBLQTB/9MA
LL/OT/bs+wkbZk+SXYQOnLZKouMqxH0Ij0xVr1nqtSZQ+oPi1rTseKFXtY2e7XmY3xyRac8Eqyic
+Nwm5lQjlSwwosC6oghxgq/h+VmFZ/0evNllgpYJYgbn3Y+7Pef7Pz5gASx0Wc3SDu0lNIq4lmIC
K8rc8d4aOTV1wErFk52Ef35A8+NhF0E+UIqhJ1atlPHbl10ubi7qNwHi4F5sa5RT3gTU8ZG97SYx
Ddl/ksARhNxqjW56Q2Xf6LnC9HIMA7wyLOlh7PU4y7Oj87uMtSgwfdw8An7+1/3zq+PZnfba+f++
Ax4rTpk6XojBoDC7FqhCyFWjlDOvFCaGy06lZDIpT/0QQ3527Rv4LSMoatkOBDuH+86msbbFFFk0
HSrlUStHWPGy5oz25fqLpeaQXO1x4iits/vRD5rKKa6yR4q4BAva9pxhX9ce/s/q6aN605kkyBH2
igfRBMV57cOLWLkZqYajTw3I47wA/2yueOSwCiOfnBvzv988f3B9pbXQ6BWU4Mc27RZMersac0oe
Q6f3zTovFoFW7Iuu8bqK8ip41dpar3roVsgiKdBkfHRYSdiAcLtn8HhgLVS35znGga1CVacKEN3f
o1GhFA+Fc485QzY+/v16jRXwUdVd0WCXMpPk+rdYYF3LwnmmQNsU7xcFgGJoVj7pEf8iddnyEGiM
mNCbWZ/c0JQAkbskwKeuBK2bynT0vBgdcGGu6uwq0WebP/66b9CzdrDO2NryUFmjLygJEWqx+dXF
9bTggc9upgebAzzQ/9y0iMGPE0WAziMiYrpxzDwFP+ausMI71uY2bPOU8deiSTqvLmBikx3iGuV1
mjUruyLCVKp5ADCgiMqRCjbpj3h2G3ymtLpr0VxZmQeIFUvL/Dfv2LUycuO9wZo23W2n6N9QXx0a
w2T7DKBHCsZGvNZqFMbdaEul6ugQ5Va6hqon7OAGQuA+FN0b1fi54tjVSg1pUrmIvjF2NAOCF3jK
HbRG82+RDgTJJGRXC0iT4IYT9Xs3/E4DiSf63AqYn8T3ybX//AoezzYwyRENdFnnXhg1SPmG2sSt
j/peQoQejYYq0Q40JNWMz9aBz+xNAlIDj/ClXjcmG3Lf5vsSYwqKHTcyx3spmGOOyMcDw02ScxPM
HtydtjDglTLWb+QTL7iQedbnLaIZnA9muHRTkjBT9IkdKaJDusgQVpFMmACaicg/buuXzj8ZetgK
PkyxKIPpgv2+AGiPrI0SPg1G4ZRJzKdBxiIZ/xhF9q6eSU8S+EpKbbzB/Y6tb1ev1QAjGCMq7IVf
9+OfLxgNj0QQuTzDF20VJ6tkb92B/AMF7yhGxTADOwGdlIUgMIroAJY+BHQ3iRFYWqR3R8oUtxtQ
qfjNatgJfvcl2NN5YBoI8o1b3Ta8GIcCiJv9Lg3mLcS23TyikW+8zsYSwbCFqwK+nrZ8Aw7rLDZG
bLTbyCpLxp4aBtwCLTKNGm1YKoaUhulFR+JwN8PjjsGWJl0KSyqsobV6Mt5We1BkT9cj92ZgIYAN
g7vyWzCjsalRQdbUj6Ag6q1i2g3AltuP3M5hcG6dR+zZCoil9JZFoe/fXFlHaJRst4Tnbp+34wOB
R085rAinIn5A1dq+MQUbCdbFdZIGm9gjlyVfpFPRU+6+7AI1C4OLWQ/yq601QIEv0+7opQfbso5d
0kZdLnsQdIGkMTitMsWyF0W4zrbhouYjYwAwSFCc/L3gSZ5iJ3D/aTPm9d1e3uiZjHhGbMdZZKw5
3XsrzgL9A46k3wk9qv3RqtrWq/vvAk5KTjuYCY+SdXygNI/2j0KwnkpZxFCVbLOU2GtOARDDhZts
QPMjxDkWEhXGqpVBiO7ZGLDHcKpLZmTSULmv0sQAJ2OLzwaQUizUdYX4wm0c1qaucMCeYULblk+B
DGTNB7k0QEO0Ul5lDF+kJbZa+UtExaJV22ZMrUVoa8FBI5EaU9Fx/0MQmR8WuBJsdXIBwfb+MHTg
eQeu+COn4Qy+1uBf4+iFonOyjbKFGCHdP8fAFiBYOsAct0ujJh7rFFVHU2l/krCj0HTlvjCJS9Hy
4YZo1eOz6Rlc1oXsLd4n1+54efMdqdx5SXP/LWO0alsBfY3y+LQn1xog4mvVDQPeCzQhnIXiTla4
/otbcY7w4Lw2b2UoUq5n5BA58PPrzRf6tLHkWyRQ2kqMws+x1q3oHwRYJ61RkibzYhHe1VDDbH1Y
+0MVI74D3MWn48RCqg5M/JWlbXnfr83owa8/HEY6u8DVrm8aJxRyXdcPltFzsJlKiy5sRWF75/xu
Gdz4Kw0GXXUf3puU7QwP2+ZHYnfNscP1x0ROKcLc3T2gU9F7K9Pdniryk0jfMTX/pS8XLuLs+1KK
WEoD7BqciQATPJE5bvgrww739Ek7UElIiNRjlHQba7r/BhsJhssXFLixHw3itM2fSWkjU9K0uq/V
WvdSTd0RI1Q+vdOnD5HULzCHFwkBChvYrN+kBhwDP7/1DMlvflBllOF6pDVVElBhqTwaAJozG6ul
HY6R8LHpbs5yZB8FK9ZB3wsQO314ux9zePvwGgsY1lAl5LLihKrAePf8Wysz8AO8rRav2Q4+hwCp
bXzXGNcsy8nHjGtNW3KX3LB8U+aq5qaC93UF+YzU0UcOcHVAaS73M5vlt/mndqr14cIRwYjJNSge
gvik7I+01a9Cfg05ASvGWzJClIWaKwJXl4hj419Kjfok4MOBsXMBoBQveTzbIOL9DQ3t0gW8zSel
ixirVg8t+gMF6qClq6ahBo6c0NKTRj1j6HWHM3Gz0tQZmAWCOEywy5awm+C6p+EZuAza+oQ10cVB
eD7iO2tlFMoBLQagTgf1oLJbYaQj1bHuzP33QP/5ZqqeYsM8syoV73/tHPu9L1ouq79Ka1eKAcr8
e3a5SUHKgqRgntdgXWgcZHy217kw96IIb2g05ThYM3HThjjKD1ZjgyLxsLUsF+BM77Acid4t3J/X
LapG9QdRXysjJdUceXppIp3Bol1ZPNdMVf+hzjX4THOBEJhrdSjeTou9BSIJVDX+Id5Q2OgZWTn4
jX7tCmzKDHfH1G6QYTugbRlJkuPxHJ+2BfskgNVYhPJDzHR0L7zkxAXjJ7FDRXELeVwKdWNR6qEo
ealZ2/6XRRqMv5FMs5ovVv9jDfP39KxXbHk2eZPMPdZNkw6pMXDDCGa4gYWIFPJ0ynFJHIxZzLs4
/sHjkys8uD3BGN85DLXSnwbia2+0mWQHLngeQrRE9HKjOCfShM1qQf/fZ66ONw4Le0vP8iZzQCuU
uxTBRzRVPk7HgRj1jONanA7K0aR3K/ovbC07J2eThSdPQFia8LNSc5ccySXEAvcPBznhTtrkjBIm
E3NfBc4E6z+4aZNhlPG971Jr14Njww/WS/eoe/5BeHEa3ncn6e7eYz7wFQA/N1TBWmw8ZtOmqETw
uSkTHF0EHUBMCVPnyKA7LKCxpm0p0iK/aCPEjKn4sp2I+rEEW8oRDt4jR4iHb86rWqO/bxKiE3FQ
z3Ijd+VIKu+rHmEP1U1SMzlqmYuO5DfVsxcA82EhDh/iDlkR1X3jmUVf6iejOsfwbWZRgpSAta4c
A4FieMSBGikX1UceKxmcdtKnPlJAQwE0MmQjNRssrYtR3YMNKxh+0/cP89YJIatUBUOJzsIfny6x
VqNx6MgAVwVGAxxT7MyjM1bbACR+agVUq0B5iyH+7TjqKIWzXnOJPEwz33KJrtRBYsfYehCqTG6W
Kat4hZfXcKnxXToSNLZ40YcNUJE2BxfOSZWM7SKwkfmquBCSYhLqXbkvx3vxBBbmVKTFkaSAqfjI
TQjW5mdyO/jzF3oHNcBdfqLzMPBj3Ch3yRMhVlkvUk9BTF19m73g6s4ojzDNAbQ3/UtPC4nGTpn2
Om2Q68AbSKJy2NHyDdV7trbILFTnAjuW/Uf8bCcM/IVl8EABkhp4TyJfunAsu3H0jA4PPRIYxsNW
5w6D5VfA7WcUr1peolUqdywqmznLYokMDWtu3c8spDt5pBrN+rdJyygNgJEnqzXM2xgmyf14cDmV
T4IHqm0kmejCFlYXPNkpQhqSspjzJs+sbWDPZQEawXyVroMj7virE+lWTgCXK3BsRJ7j1HklDWIh
uhZcXgojnLiee6S6EDlZi+iBYCS2PPdWdRTtlj+26HaEFuPlqyqvLcdw+ySpJgBzwXktIBOwMHSr
1KoQiwC1Xay8U3+/U4F7yHjOIvZOheF7RSWkfi0xwe6oQTS74v0JWhOTjI2nv2OsTAsUv4SpmL6L
8Kv/1uiEQEfhQBNY/gsbLjGyyDLFLvu3deB12lFEg6sKtPQsaP5HDxVoBzhPYeaY+E310FOfSAly
dK8FeV++79MqX4oiId5/7fse7Vr6vDVMUUUnGBLrR0CjrvTND9fhbJ9buKf8BvixCKUjnlw7sh89
zxeRK/kA3ufJlzTSauw4uqRT5PgAEIrOXmM3a5L3V+5lzNig7G6UBPQlLVxNQKQNLC0Nir3XanOM
G0CjdVu7NzIANkfUaDQBIiS0ggmDEQ6bqVxoPBiXRGbtRMSVVNU0nzPSfnR6v4ND1OKmg1XNgq96
qHO2N2hQgmgKdoA5pN6rdEkw1uYlhECTZEdrcjPiOdIlhccWVKNjRxgo89HcR6a/YSsXxzKWCQRO
OwpzLmn4JF6wl1WiSorl9o9H7yc/E3UitThkTYi3Tpml/qeym80tytXGVZqIS9v9AjIIB1H5QH+Z
fLHx1cS9no6aGfbq9srxfSdPcSkILR1IN3ppzCM2nuUgYyMJs9VfEvM/K1Hc2jIEeFBajL4HG7Tb
5eC2Q4inhSgGOd7T86bk9iB0BVU2WS7g5yuyi23agdEhvhnT4KTDqbEfG0kKldT+IeoY5dMbhP6I
XLxCvEm8vKQJ4z8ezVjofREjez7M9lfYH90uuDtJbMKR7+s/SjKyCPZGvUDneCBstMZouuLifE/X
QvRotD7oIRCjjhTUBrjHOrC5i9WcPeQNsdTCdBr1yiUG02kBK+re/aubfzv+6OGPRwRMBQht/Lhu
1+VXLNPShkm+x+GfNKBrDur8cWkpKa4rWjNFyoECoRMdxHBq2uJnFnbcU4USVDXfksAH97BsrrrD
Nui7Z8NrGlrU5vtzaJVLslMTo6FIPBcuYueDSs4OWutI4RnNQ/G8RNiXUTT/RPdrct7usnvY5U4P
+UcQH8j1yD85PWykuLLYJz0TvyejjB2OFApT4V+Od40tJ4DoqTfZbD1+LMkwPfjtceV/IZFIVYLH
JZ860KsKFokJohDp9i/wH8pIiyVL8KvwKg3FYad6t2o0y1HSjJvPR/gTafQdESYVlWKigG22LPLm
su9DbzOmqM6DSMgihBiHh+RLwDirhPwCkQFVYp6UGN8tG0eQw3qgyd4uRtTflpveXE9jRB5RvgCL
WOlGZDEXs6wdgxPQ+Tuyp4P/JdPnFz8/z8HT1p00IXeKOogsQWvBbjeYjYAGmaaURctVuw2G06WQ
ZY2HogXrRhSBGGJIWBdmmE4/yA3RwjWzZAHM9GUDJQsztqCJozE+Rf8IJ4ZPYd/DmV9pKqgbXY3D
DlTRGWBP6TJHgQamYVzhLUxFYSsTzksjiQ9IHtvmZoS/gYrpXEc30UERHiS2lYf8ibvX3Dq2lh1q
ddfivIzD6gZsHDf0/w3C/Ppfz4H5svNijRA7rVZYUCoNvVg5GiDQ8qvG3DIA99xZgyhpOo5bFT1T
mEYvZK42ZoVPnZJZigi1iJqOEhTXvhwi8A8LAISuUGZqddDtoQUJX5CoADwXI87KAfQtg0IxlUxG
8sagKL7bZTxH0JXjASHsv9qU7YtJOb7b04elDD54mQb8qcIFCPa88lEsRQtFDzOKiAbWRjmOom4m
Pt1212PeTevmdQFhsSagThMAxktjGznpGdwkqqTrWjTGgvPNpp2iAAMPuJkfLrmsuJjjfN2igDxu
P1V+DzyG5VcwRyhKS80VxZnc3zFdAOQK/qpbnU+gGdObZpqHNJURzRhjX68FUpPnOPH50YVsKCpw
xZWg+8uZhdgPFsho/qM/kjR72FOkXzRAtVU8MvYw6EzexDDDVWvAGzgOcEuiI/dCPed3RaJahfKe
H9d9x4cTvo4Pd9dwvgce+p0/gVY3WP81jnEEzaPWdmfPFncC6znMfo7QRXKYT8Fv5k0ZLrF04Obz
OdYbFNmbh5nH6budJAAAsSuRLfJ+TykE531RePgiH4XfTLLpjpdtR5D/Id2s1uRg/9wsQkegCm7o
Ovf4eDgbnjIJl4jLsxPWDYGwvakLfTrkhobea+EnLczzDXlsqIwaOgTCasEX81VTTh95CUuxNLbz
tnPRa/7vqpo/mHve7eHsWJmKyy6J+Gy7OoxrIkEY0QPQdd0o1Y+QS3SeUTmFfFL3VXY+ZoxEiqlC
UMxaQPtvXl3UJQA0lqeCUK1xMTuhokjidMixB5XeKl1Z/LFWvGf0Bq4y+DjBrB3KahyooV/q/PTA
M88p8CmzOdF+zxNnNj9KoeA6kYNlEOZBg7UrwJAIaV7eBXIxAyfqKEcIEjCIFFKTSyaAUnHkqjW8
HX+vQM2v6CWWA23PIl321c5lbNyB5Z7sIYt+PUeZAJr7YqXAimy9mIjHE1nnqqPzuiovBINEcCeI
B2l88aixT4Swq6VIlSAm3/LTF9ra6Kw79THC6suy4dvHHLgtKJHlvuxcaIQLx/XVhCnpgArC6m0o
LP5ZDWaSAF7H8uoTRV+I52+lDBfeLP7HkTPzaA6QsFmUed2wVHeOSPyRPTWRFpM+Dlc+EDzzHC34
dxJURGpOMBHoEyAlNLNZjITqP2wrr2pcOrpWd6j/L0HHP2Q/eSvZ1sGrd3FFjZCCf6TcWzEqopHF
YhIlNsnV5boIjhJ9KEu5Awl88FQoy4MzmpxLfWrRLgVs9zwbVlaxeXQYGrApxJe4oECeAzp9OTz3
eji8HcsbpGfvacNygXLK/gB4lU8rFWaldfejF4A1hs6vOwDQRXjl+0z96O2E0l1DmK4UUpMOcDUZ
7XObjGFvVOAaYUJtpzEFYtbKE2OaejJn6cDgV0WWq6X4P7eU0Vmv+6iJk3I6AGigw6UEDF7JrKio
cnxCcKLf/MGQSdn9oKNZt5LaHcMxpptOwxt2QtQKsIbi1YsLVBvsiV/uSl1b1sWEvpXbSX7ZSR6c
RhxShIkEicCF+C2g4KyQPynln/k1N/vbeyL46qQaOZZzzxaINII5czAL9HMc5twK+/DNNkpoXwAa
t7IrE8+15NSIK49lRAHibWjm/reKzwPGUfj04eg/8/K4eWSTK/FH0zI69PPwAsx9Q1u2+mFCEvyx
8hExLjtf1UshrTregM7ZtqRsvGGBjTtdwc3T+DUTYzLN97zFip6PhEyiWF0f6r+EQ14GB5n+SEbH
IEEmKUN/5MwyvW/Bo9ZqEQmm4Ij+t4V++zdVa7TAUi7B2V6Fa/6FBiNz8nWL+kPPPpEiql6wHoP3
mtfoXy3/ZkDoaVrb5kCZVTXnLD9LDPYMBiYOUk2JermvykUvhBwwkM5TGcCgyMBX+8aErRUj4Wfd
imLDcz7fTc2zKIq5Ln/dsolan5xMiNOLDqCM/+1Cdo9Gx30lqjwYVvVgHb98O1seCxuOrGVJeze9
rZsg5PaKT3+F6k6bab2iAyqWoTiB1pU8dnA2fMGNbBzN4SHUF+s+7EWztCgdc8JfEPz9pXDdjzKF
qwf2ywSnAX5XvQ/j0w+WG1O8q/RoBwe3V4E5Z17qOGHyuvR0MJpJqUdpnGI35XlLr3FKY1f/dk4Y
/3TvIAhZprYb6lsyPEBt/sGQe1bUJryEr4kFBWynMK1sGsdxdRdHsaoXW6MCbPJ310gY4BmI9gmJ
MCZlvJJJMJ2kFULQ3TjQwBo6eoDkAJLNHAFdW2vXeZT/3z0dEJCcpGBWzU7Nf79XW43hH+hJ19jS
utBzRz7BgcQqM6FpBMn3+RNeieFP0jrg5Th/vMSmA3VZnwhCbMPFQLmq0WmNI2m5CpIQw+3gme8I
MLFYLg2AqtZ2PXLAm59ekyPFz5olgRqKDaClmhV67Migau4GO5DaaoLDPyV9ngQZVblv+9t3bS+b
FTyRIsxXforLdN5YPkVo/YWRH8TOVOakuMrm4xpPqBPdg2BPoCRPwo9m+5+uixao4PL05/TLinFJ
RB30tZ9/xz8BTQYXZE+AnO4j9YEEE16hi7nz7sJUu7OYD/pVBg/2Mg/2OFlNWiI7mkGn5xe8kZeU
ygVSS7lGw4Py76t9FkoxxhHgojHRCynu3Gs924n1Xa2oXpLSAypg6haHwcg5RGAadI4KPcWGPyxG
dJCK3/i1XtrvvaelhMBqtza1M9G93aFPjZauLutC6O/szX9uEB3EizC4yZSGpqW0Bxih/2NkwYWZ
EuF8dHW1/1nzYG4nKkSinZW8Dni99YQFP+UcROphx3PW1blSMOx1VPh8LNl/yoojRc8GQEYx+IIf
zanB5v2weQAHxZda27cvH+1y0jhQ0UE/Z3TYH2O+sfMYaJSWW19IWJBpn6eRE3FbkIfx+5i1fpf0
SSU6AvfFq5jpaMyghg7AarpzAoNq31J/x46h7tIxm1Uf4Z3L24bSAGTiLGUemBPvEY935wQoiq1I
0wJEgVKBds+8ZUUI+ix3g/nYtpclkT9z6k+WE4v3p1dVEAeg4vjXRSo7QouA+Yi7nd6F95CsXNGl
CWtRVnsiILMwGLDFyBzkoZIVgFyHZZDZpqqF8PgJ8XfbCPPBaI9QbzTvYuISbDa0T5Xv4kdH74jh
yx9e7JTi2sOr7T2/v0QxtxMmqM9HCtJSeWv2cFzCY6piW+kFKOab1owuHpvsUf0LG+okphx674ze
H2niXKF/mwE0DgehNKqesCN0QGdjjUmOQ1lbjpnZQapErnc5UEUT9qKracZ8cFMiT25HJg97L1k4
PyO388lXft3WBmLdmU5+KDHS/nyaC1HkEBAFIGUMghlygYGswQgewHhfiYT1Qg/mmvTwuE2J2a5f
CBggTFVHFR/++WC+7VDZzIR66BjnikDWlRUBRWjjpq2CSLWgfSWNuZzcFCK828c7RpNoX60vTxz5
CzVGuzo1MAPru+Yu2CXADe1yqyOBdmpwxGUe/nrNbxfbjuUYQM2ckEHktRjGXXCTN06A9AkH+NE7
lg/kCnN7b83YzZG1NbzTti918+rdv1KoffMbiaz0MyTHBzoUif/I5mVYxXreGj7WCZ+J+cgqBJxu
ZlLTBLPRcibe0C7UupQ2nOXmp5XmFsVzSxeaZ4bk7zXsJmfSi8Xp4rMUhrAkMPFogqxEwNunFU5/
VBP64pl2IVTPPnp65HpU7vVMhMsG7T8D9cyFtJlu5339QRn6q/ALsIXg+GG6GiF6833sQG2xq8or
1B0vS+ez32lzdDeyYWpzJ4sslnL6Smc74RusQGVz6DJO1oDNm6HaUiKDeqct2lzOoO0kaNsHTW8q
UG2Zwi55WT1vcXtH+WvbdvV96Ja9YzVuyC4/ZEwTPpxhkxzCl6tmB/iE0Wg6lCOi0aLviubHy7YK
f/JggLSMoJydvD2mUGVTfSA0/C6WOkt3yppjSxEf8nPt9hGdtx4ZVU+oEPcJAuh06bFRUeREdjFd
qPwMexj7zytb1SI+k1LzHf0zQ6Mg3c96wOnakbP3mi5K3kUOrGl5wZhiepif3chY8Eqfk85rrxvH
09467ef165caDwltP+OPMU6mTtg85rhEcGsmtTV27DP1MtKzLodsnIwCT3Z02JX1DmbgJTqprqyt
fuXyyWceAfN4y1EKRZq78ZytComDjdT1HAQY79X03/Cz/R1Dl05TjeCNLLfOaFpiic670GjC+wVB
DJIxCWmbW4K3G04ltB8hpt+0iL5Axu5bOL+9y3GgXCn4n7nlDqtHiMaGBHgiY1QGXLPbVNeQN5e2
9/4zrMw6dP7jq6LVWhuukhzkLqCf99yVpB6aUbrBAA3yhlbVOl9L/zKNMkA4JFO3DU27N1aCmRYS
iYB+hPWTyQCn0CzaMaQ3Q3i+k9NGJobkQektpCjbAlb1T7kjn+csRtA46t68LvPJmF5hOE9MnsNg
7BCed/v2GLW7CxfjmJ/qxtP/UDoO5RYOOys/0FmsSDH+EoOBf/0xa7XEW8hGhZEMg7ObDvC5jYbC
GRXpNeDxvwdI59/RoycsXusCP9pmcw/O9FfncQcOLAovB9wVEOcJ+W8Bo6KkAb5Xzu6MrOcRFZRa
JDcv+96NyXub5scf3CvhEDrw7se2jEFzARIUfkF0FllBZXBfBKj2SK1IVD8rt30TyEHw8te8VP8x
CuduJOYFiB+ykXveDEUj+/dY0ERkFu9XJLe5CqUi1rN0XkO3Mb4sPOKx7GhtWLyfVAyMUaVgoC1E
bu/sj2rWGu7E4LXdYNyEjbkiIGQJYHEqRS6jRUpJuwNrPiMlB7tmVMPpFjrDvzKNDWt0s+OsrG9K
Ksiaa7/ppBhLHBxvYFWwvukcZJ3yFSM0HhV8IAV2ogi5tboqR+o1d+eKvX7jhpgsA/FG7hu02n2V
s/DXxVIX2A6F/uzbfX7uQmL1RK+Q/lrfst4oEQnokGZHvOlAzfAR+gONkPYnN0plbFCgN6kb/ohG
jiwRzPSv0yLi2fvLeay2NqzxBm2hneHsr03VLWIhIwsCgplyot7wrX7zKt0mmMxUuSfi0HnEI0Du
zjVMt5KQ9+JK/NLulx0q44tFmAGpoehpHyr9pxbtnQDHvfBSMWjaNx4CZfEm8pdrsseVibxIkU+f
PtEGd3/4jC6t7+Xvb2tIxdUCR1TsEu3MLMCwxW5BhkwmsvsoBJHyWCzU4FxTiEqlMbsh0oU1oIVv
C23McIuv9vu5v2ipckuE3+u8B5+6K1d80EVzq2hyO9UvKW4AvzPjeRWTx1/JlxF5dmHM/BJoC11m
yobH4ALuL+qbk56ahU/plfTuBW2Tiw6fjfDGBEdUWAvc23y4vYzHWWKCbsLUYmwJANMNLDVchbKm
/1I/nOC7hDRcuyY7tKRFl4rQ70gGjZlFXWhoLICb7BshFeIs5epu2jaAbcVRghoaoW7JY2/om9V+
KnPxJ+wwRFCqps6OdmPge+CCUDbTgrwUyLOCnJ6HkHD3EjckMfIJ2TT4NxS3FVtqDgbE9BLS8Npu
Z/4ucVPn6qJfx0VyjOXvykIC6YueICPY2o7zO056KW6T35P4T+harsN0Q42gR0vbE2G+33lIJchI
ol7cNX+7qOBpcH3rWIp/lOeIXO/wGEzVgBXxvlJGkG/jcZ5V+lBCxFaCr2cPbrLM1v3qHhlQJU/C
Oct3e0zo3xHB2SmHdSuF58gvloRoCBSoqv7n+qIym5PAtYZ5MgzNCVSCkc/qXtcOwKnvNmuGc3KU
6TQCs+E4HWXqov+h5k2TSx+o1vkGX4fY024ZEc3loZI/t6SdOi1a/KgAyL7FZRy2N+j04ZhGnPus
Ttf/17qVF26W4BC+gxFweb4BfvucUfz4+HJBT5+pJeMqEuDP/8xMH8yWWBuzMoA8rndecVNpknTi
hPiQ7vg+12hY6C19e3q/8jUq7KJixL0pqcCHRg+T+BHy0zLylV2TDd6d3+daQbdP93ZWENfn1YIM
OfupLnGagblyO6N4u6Elbjpfwlc6I2eYTsWTfPtZCQkiXYgeL+9BCe7CWY2PjBFEOX6UYbs26vHS
R8WfCE04LbEpq9GF6oCygV9X4eY+0C54uJzpyNxd5HK/IFUasl3zUMuJHD6maM0KWoFDmRAuqAsP
x/uwPuwCfgt2zkcSIp0vAItCUkoeLcrEf3pUgjks3waOaeiobJlH7hEvaeN502z0N+M3KnZv+fv0
NYchu8+WpYnFlMhnWvzRW0TLI00a/z+rzn4mt66Sp/HtVcSpBTff9MPQnfk+ylQ+pMCfWzRFsy+F
cP64mSoAEeuwZ2egoDmr/XvKBPwMIt+iW8V6AfkQu6ABu2LCpaPofV6mrX41x/1slLT49nTWUp7l
BeEv+N4H75B/gUxwAoDIqAcLPnUtpyZzVivQegZEiinaeiZdOpECRCWkrTeJ9rapJnAogXzzZUEK
TgZ73HGEDkU8l9rVPXMd1cL/dajDQhb0XyTEDh5qL+E71OBQkzlZRRBhz59TrqK3S6mlRZcLXV86
2R2GVNywUfMfnMkWKovJcdRC7OcO7t1yxdzwBWXVwt4Ssw6RIMG2+kL7rxY0MP2BOn4A6INvR1E7
KgS7DxKroGc1zFiicFxxuKRwO43fCqTnt6djFMMmD22g7WQSBkuSXg5En48d85hVaSk1r3Y6shRh
Us8j/yP0yQAOZbCugE66O1YxWu3QjKR9MMZgvkQk3CVkokQGh/hc4FXAwe3S8VxW/Air2N5+5Edt
0Q8h1s6xfaU86egjILJHZY9XJLH8K2J4OpHofkWyTQ+O1FHQjyuS+fZpoDPwOORMgQngAW9sqVSx
4eH+Wpu/C02AKvtZcTHtGvz8/BNVYjS+U6JtAXmqI86SFkG5Lc+sq473OpF1idBiwatr8RUauI24
0RoK67989cKgjDolVyXeUky8fuLowbKI6JNLwKSfC+oVHcmxiIrc1YhTSeCmRO08bjx7nUGsSoNq
HRbqh/aIn47B8s2b6UqiB2A4Fo6htIOX69uDnZHlAknMW2lQiSkXouhtnm/QNs0Z8/iWxxlugF3c
Is3fW9vjrQGonOss+9dgJLluWkHzs7RX3S5ZdFwr5kd3r97HE9OR+VODIBOyzRbCnrBpBG5D3V+p
N9sPbaKshf/53QCKD0fFObWj8vBQBbtz/Y4SYQMj3FuYlQ6Q881VkHxorxHB46jc0Ds7RrydXya9
kTq/orB8QwQZRwlo+Xg55oeMD1HFfAI3z8MUGOrmy0GOykdXEQkl8UJsQ+40/pRy/PUw97v3yFbq
SsYkd6/FvS6utjUplBQ/Z1pN2sTeXF8r8LirI9sK8JBYS9ndffFKDtL26FWGjTNKjk2nPGo4C5AS
XqjMcuicMr5qsAVd6HGk1adk3cGbgyh/JaddT3KCdT0ACzgRRBhayIHRMX1Y6Yq+tWPpsMOfmIcy
Cdk+tXjRTlh5SjShcTi12KjjzL34j0GUFmNC9lUaIjk8yDTEY3I9vLxRr7Bwzq1sZZ7erk0hfjkf
bEieesBAv1r+kE1y0Mu4IRdKydvZDPMsimF3PxSOTFGVwrZkZn9TODLCPmTqirr9GBaY3KPActiO
IBcn+KSIBAYNtBp6HCQGLP51JXSUowPwLWY97Aw+KMo2McYDQbQKgX/6acMNTzqN7kEOZLHjqzKs
sYiQ4lUEGVnV7GjmxDrYOxPvvaQ+jmcSGUeficzyoWyuzfqAvOs7hWOccgSsiXaP6bh4Wj5xbnKE
YpqVRcVpnuri9QBUxRz4lOESdWGcjcJqkwsEN5o4vt0rbjQf6uDE9X7fYYYWYbJ0wSnsRUZqeuE+
/MThiBTT5oYKXDb+0zExigecW4gZnBQ3hLkYZrz0impiGC+/orPXa82IlOEJqMaQsCEZ30jfLQiN
nshAzzxGcZWXqqHK35ySkN/hhjaciRrg+rTp6+9Ccl+TYPXuN25fU4wRFyvRpTfpty3rcco2bmYI
b3pI/nkXdfNuAWrRG/Q7kDIc58JnYp4OBNju++YPFB6PSEjLr41wObYg+JHWfMPAbAg4uhcH3Vy1
cSEy3xRRdPJaGDKQMxjbQJZVOz3KoiizeNsyhUM90BZ7LtkFmoOWrhEZ/vE9Ye1hx9mlDW/OH7/e
Bg+kf77aGOzRUX18nM4iCaEVjj5LT/XqY2nF3O6CH1wb6bzjFHOOcBnntQn76fnSCeFl3F+ZK8l7
sAIsLnnK3HBWpGrcC6xGWg+uZ4e8Qj8gDUW2VSZtEn06ALF+VsHtSbssiElvbi+8DdIv6DZFRhn/
svk/KCPlGSc8T8pckH/sX4HzDfgH7eeb18nUQaPpt8Ce2v2O+MUbQBM0dql2G72Sm+GaDz7COYI5
GXwHLGc7dRoD/wG9cuJ4IPzigsOcn4hDZIQETx0VdaEnWp7zpqMcaGfkdZCMVBd37+R24ptd9ESW
zGXr+OQYtehYAHn8vRLUyMC4TmzapE+V9ijvt/zzmX2WdENosiKcDL8/YZTtEKDkwfJ+CdnaMHpw
RfOsYjLuzRwHMrIlzV175xkggvAuZxU3HT+RX1zLGQ3oz81YSZiiCoaG/SMUnLUhONtwXf4xqcl2
lbmhAUvy20Ol047SPzgnWHEqrtREG5JvMPsWUgcGgFvKLTex8dGqC5Hw/Y4bekfhiZyQ7Ofv0wgf
FmHprxjO/2gRbKupvX3qiXV1S6aNB0CVHnDj62klUdKhk9k0HT8pr5WwZoil5LWDYmy2jCfsG3Au
El7pwmwlAPEJJAz6alQaoQgFjCuNUagM5my7EK6W7jd8PWQK77ElWcGT7dQuT7h2ZmQ11k4Yuxkj
wc3Daz5dFdxmzWsyUqjmRJC7uZzCM5p0v84W/+aBOZL6H3Rw/lvXquRoLaG8hh+5kGDVerRho9NM
uPqLinOlpV6rAnAGVRyS+mvs8H8oRRGCz13DRResYv943+rzh+RQe/JoumHB6VnMOdrLWYnzI1jb
Pt9kEEtGHb8Ys7aS8qpfupk1/yFGS2YUE9elcpv2r7Z9OqKYy+n8AD4T6Zg72TVHyC9CGfvMdNwm
JjgZmhIYW8cumwxeF7FsqYGroC/kbVak/mpay3sSh/ZhQL/3MhyFuVcxwDzctfrv5q8XR9jg3DzZ
Vn8n4s/gaEt7WMfJYrIyyXvqnb9NhGxfdRu4dZ4wgoiXM/uvbRq2qKNHEKWL5QJZRmMnmijQ0Pmf
qfqZzTnSzREbp8T/Ph/iINrmMzoh378uZqvJpN1b/QV3xGTTseQtIc/EiFP1BZroztbzzb2OMRXX
W7mWySTNb8kxpTxFAs0AOJHxibnZvBnlH8Eb1H66Nyv0U6p0/usppwAHoIB3skn0dmKE783hjj3E
qDZ0xLpMaNdAqVRDXvOa+PmhIMEGfQiaLdlR6wZ0546g9DJCZJ/JJD56btFV55rnDq/UEmrDnmNm
9E+WMaQagfr0g2Gw9Wndw64cOrJqvCj+IAYlAoWY7WtSOO4KYxhL6zobVTK22Bsqdq+PNDKPDXoQ
b/y3X2hlwK8JOLSJX2g7c7DysuRtjYF1aCpokW/yfWAiAtSYzOLqntUsoMGFeVn6ohF+pl0rVbvE
LnUZdSGjfLks2td4uGC+J3ryqj8cg7KvRbrrwXhL140byT33rXSvk06tXo9+exHgVsBW0OQ0n66u
84SRYwiZX+uBwSpJ5r1m+bjtE7FCLOjp1DXUojwMRvFPQeal49QHs3TYOcLGJg3btTsZo9rYzSpd
rm28B+VuSvBThgcNJjAKQCPZxl0WK8SDeuytgL5gP3JOdmbpCbU+o429Sbiqhcq4ovEOB0XE0S3U
r3YJI0Xp/pTkJPiraWtCGq1KhXGYfieUIHab8aYxf9aOdV1fXcNVI6qL9fEp09DREKdztzDBQCbE
ay/MA3FYF12sGIsTyO29DLa4y6TYRbYfG0B3Z/fNrfGhZBfL0AIks4RW3tbOFPNXQ6OtPB0QvC/J
E76rs/xVB3TuLrGwb61VNP8nty3lwc5d9moTIlaWrwumcEUi9DWAWF9SJBbdWVRoR/gI/FrosGe3
ETbyxmCNwA3JjTpPaDjAoqcrJjnFr6I1ucC5zBv127uB0oyQSVmPqft7Qcbodfrvc7GGnTD/eoq1
9dXuXk3DP/XYe7qOpS9oJY4AI2rSlw36uMx3Rx3WZH+41b3NcIqABjEU1hHYkvgi+Tk/WjVOgkHX
jWWqQhu6gGY1JsyotZB2sySHGe18ZzofcOOX1v3M5p1Kam6UWYy0qkghShQJNf4YlHYBdVC5pkPp
zUZwvnmsnrMZFsbCclYDX7Bgmqh36c0cKB8HUsgCXzQ5XmrMPJzA5A1k1TSA6DKkzXJpPQO4uKpG
SaA8A6J/WYHNAI80exFXDo+eaCwYCJVmpzYjeo2DAnZ9XcJqg7VPSKhiBYHTlSrmK0xVEi5fU1uI
SeTP2O0267ucr5dwJ2te/Jlw2ZqUyUj543yKVDq/vW3rfHgFTquRONS8XJ/IcNL2C6mhJEfTfS/0
uv0Z33FihCu1+h0AayrCMcvrE4sdNv/sO9g44SauCBoGnuNlW+3hUJcYLZyqL4vlufGE9jTjezZ2
W/ngF20qiP3log6Pu+MJzOO/W9QkNd3Af6R2ivfV48PXIUcHOA7//QAEHvuJ53E66XXNIkZP8hJg
4Y4N6Tgq7DM8N7nMllwp1J+Q5ZMDWZl3rec3/BaEP5ByWbeN/WKw6J+6g/UVHysaikvjNqZ06eeS
4oz5rqaWH8ai+ZOmNzzBqRGNSqYGS8mfI7QrlPiLROqM6mBdzrkP/QxKCqu2znu0n8156TT1zQjd
IBmaQvttDMDrtd8kZBZW89HHz5eJB6Vs8mJfnygr8N3B2pwjCjJ9+ospYZjSBPXazDzc4KUOW0Ov
QtxBG2ryhOdmi/eSwBF7LdNYupRtM1xiy8yEQrcbbjaKRjzz17bjVbYzRD9UjqTtVq2w8DHxoT2M
2bsAOb0f4xKjo9fJkLDMGiGp/YHnTomY2p5AT2xPABucFCsBNVzLSViEgP7GFperoBQJ+9eg+oMc
PY+kdOeYN5OvH4kuZZMzsOJrb/azo352SMPO05hcmaQLS0OEB3eSXfaEx8dxHkFnXdCaxsDekXQe
rH8ofmjzjEXqkeXoypIDRnX8s7LxjVzG4HdDlgpJft9cLBCnXuSyhWT+0d3R+9BgzY2+2HpRvTto
SKnwQP0eLiNCwRhfPOFPLLb5ad9O33nReBvKVv+vQtjRpcGLKJeombOxX95EFojAH+DWjE/30HRW
efy6tf68wY3n6X8G5XFWBzeM0qC7xvB16dyKjnPT0QvBF+O+IR9pXRDoFS+Ze4Ncq4e581IlSyNF
0/emz5VeRi0Vb5/rhfG7nmdbXV0PfFBG5Qn22DCYoEXn7/DOLNXEG/300zFvPUl8orno8ql8JA2j
Q8sT0BqDh3HYubaviHJE2LNEdVa28h/ZsiGG2VXcPH+SweBax1BboaqVJ9ZEm/wKrvsVEL215h6z
n4uo86Z+44JdgTJZAe2adf+pza6vnae9j7dKhrtGazP4H1mJ2CT54/VDQ4/JAq1kwfQrx624KX0J
MukgpdRemE6tekE4tqvZTG9nDokuRflXYucHlgHsmXI6EAi7LbFxsoYZsEI6aDvtptLUpDFDqSJn
a7cWV3jD3S2y59jEVQ7DQ3N1KdwHPi9CGdAfjUWKULBqcERxjQ+bDJg8/e/cXddyQ8Zki4Gt/HYK
M9w27ZQBaHQTo+n4HnzZPq3izyIUyrJl+mZYSaPM0PaSViMjawQZ0zxPcU7yp59jD//I1oH8z/sh
a/fqBYyt4E4tHE/sXlQAaotaVVNZ4vpcHGIwoZFcq+ULLISVLqzdkpROXQfx4gqKa3501EtNG0a1
o2cUWAtPthAOKccy5mSU0MeEReOudZyScz0lEfeYLo5qaTIvId7DJShqFrmjXVXxAtRBuW2aVOHI
/xD7cFzaaHXk3SLSOxTR7k6HXwfWH51QOou4L52yWKn2Kj4deyU3/+pLiM+WN3b0wTy3r+C5hBGQ
R0X6+p60hHUuuI3Kn3MsrXbAOi4A3bYYtOjNTNrr7O2CCSoH8Zp7DcMQ63yfI1u+RI95OzPothCT
ybSxMFoo2VOkfYGqFV6FH+LaVTm99tDfSoWt4sYux/hHSuou8JSQim7CcyIxynJPQwAqXuApQ2ti
YmxRE4nl0DQFUZmTEYb+2pnS4caP7v0EB/arnzKbCtc3N/IPpuFwJVHXzpZs0GnfC3EuHbJqQ17T
dxofrD1Y/cnLL6bbA/eB6LbNw3g19eBZLwA4LLd77SbFDYAreaTohIOmcJdZvexju2kiUSITkjpl
0l/SdeUIg7W8rixaPbdo6dqc9eMkNFBoTP9RKgnCxynN8PX6OQeX1gNBs44+8b6MDVEG+DgOZgSo
kBeNBNOwOuEW3rWNU3712wrxayJmlI+V3XvCfj/nqm6hwGjroh07oEeSus49wGmbh3y9ISsQRlD+
2YzGIVMXDI4IIO2fb21OB0hqu+8tYx8H3+MaINNLwcMEeMJMUEk94owCRdrpWwsJW96gP847aIn7
wxQd1Z35QnxV6ZzaHTD823MZ6/lBe8AF6EaWhgt7g5UYUXfdV0pQdO5Q7BSj85cOn1DkcAqBS3CT
mTgIHGi/wZnafv4n+OqP//rAe0aB7nn8ocioOBoWooe6tzEtoGq65AuI1IglEe2wNyyVKDUBWPXk
XqPp4z9eihyVyCzyjGQn1y2Jzx3na7FrcVp8u+yIWz1F0s7rhQW8Ng4iBs+CUSNUBwoEcWkRM1ej
jjszm9yp7i9f0fsGY3E3uubASGS4tv4bDKxW5XVJTXhXmQpB3TDBGsdANLyY0jAMGA79HXI9H7HE
QxjrMudToYUbegrCga+3orEza99j2CgEE4yod6gqiNvzJfEBw7ptfcjiipk5CmckiKsZTaeWFpil
EkeZsJd+6DDn0yuP2KZMc7Z9VbIzOWDijFSYGS9Z5pmDNJ1esPxngtbj3Ko/Q0qAA7jef2ojSbbG
1p/s+V/x6q+SCVFppaz1/jkOcyUJw4JWU3b6TtDCmvc9lBWc+aeXfUxCS/h9PJ0lUkOq/JyFWoJ6
oxYPowj6zeZ+Np5uwHi/npyqfLKEdIukiUsg2hjaDTPTT026r3gYWxiVUH8wvtJEoFmJmb1eNTU5
2mBNp+kI1ibkogiIrggMcsc6cafIJWVtxi+eYqpF+2JGTHX1j/sjV263Nxea2VLD+LJCCHm09FXj
Xn02xVph+B4vEz+npItlg+YDc5po4KiBfQyA5uTnLynpt3FdsvX3w732rDEcwuKQ/LVhsOVnuZus
o+dag3GtSpW1/zBrfe4YfV4nnVWr5eyRXPojJpL5PYdvgqwk4cqQUgfntafAOQbg9vX+svwlRVGI
V+Wxjx9cnzZIon1zrhfoZ6oRmp6/c6CVeZ0bqbl6WxJRmFHgLIwawkdJV8DZcF0lcQ6xaLrZVsaK
vnzTVUH98zgEDWh6XqDiotajdQce/om6c0EyVcsLVtGXOwMiWzApejpq1Tjm8j1k0fjmfzH7v2sD
XUBeXpFoTI2NGei5f81SIkho13/N3ZjyOeEjczNiLWUC38Uwe9OfhS2YFI+2C69jJOAPHJ3euQdV
m7Yw5cTJD36XQuWDNoy9aVcpeCbEuKiLLqRqwEBEa9N36vXjUax0cTdoyHej94S5hFxPsM1GxAP1
kAVyqSKsITEsn7k/wD8GzwC090ufYZnOdMAxOFXdVsY37psElwNAP0OB0oqGqVl8GRoBfT3TGVya
7Ic+ByI2VCxuj5tdjCUM//YqlP1nxrwbbH3hHKs8wJJtfvYkdghuy2ns8uFPUwfgxa4F+Yzufivk
oUb2YBZ2BCbFJDajH5WQMs0Q06jw/rsqHwugTKb9IxS4OBmmknzQNwADtoHy2Z98XjBVcXupq/EQ
FYpg5T5OzzYfCgEljCacyl6q9M8sydg+puBUKgv4ykCoWske4/UpDxABwuBgvARbiqnCKCkh8hra
ayx05YO59anOJDLJAtSqVa89CzxQJ0hhSKCnFXBK36YLCJhD67XNHWzCqhjvzGMO/k00GQwIzfwp
kbNAZhOzAcmbspFUv2QTTSb6J+c+4ucqm2BIwMT8K/xHZYAVoD5ZZnyLIBvr2TA1U6y3lNSYnucy
jw+Em/SYXqelG8MahUex0N1BADlDKl6IK5GTnRA64sjz/dgoKE9eMPpL4wsk5jLJOWMjT0LD+AuH
Eq3rwjzwZU5rfv+gRl7JCITCrKILSCkUZxKWCJqzFRi46wPyPwUTDSX1nv9TIzEGgfxbgVwUdlqg
vbqof5vDHtkVOT1tIA3Sv5K8RW+MjoIvVuuDInwOR9cmfagn5G1I1tBKZNUHDJdn7sBwHXOI3Zol
tR5SN4pcH7O6uosjobKKFaYVw6c77KpomcQxRxVC5bGr1rtjm3DtMXvH5wEmKS95S0tAYL0N5TQk
ApPza5czGyCKjT6iWZnOlN7vARMcwocnwjPIojxaLibTYnWt395muRX4SZXHHuM6HDbccOWP2aD0
qk5AxCQ9I435W91e6LP7OvFElu2M1PoXKW/YtzEvcXz4c4Rvcir5kFilnxEROHMQUx/imCJWghIJ
ha8nVg69mn8IkdjMr1UnvglV/GsdrIRL3VZzUdVSjWd8RYdKIrLrOhvr7n5RnX+WOX+ciZh6Yp4z
FmDTExt9qCOAYARPmZCJs+eiToY9aDXma866GKGU3C87EQs+Btlzjhco7+qeXAqjqFG+xARyZVIK
SkaTaUCZkkEw1f8Tn+uKXqwJI7ASxPHdPZuVqSsmqSkoFphm9lJQWlhNe/0RRueZ0tWl7hSM02VD
rIJkv5WOI8yMr0PdejU0ezR073plYOksdIy6hq5ryCLNz4h1TvzN0YkRRQopeUFdNVr1ujZN4nE/
/LX98jDLPE0z0iA8EgN0qWXViSRU/NCEgkP6FLz2Q1UiOZHjUkCi2MYvYCiC0KgiC6xFCIOnzIv+
sR3oNeKBatVKeu2nvIUjSZSUm3Xn9FnPYCDKAMPc5WFs19+TavBzp22jmph2bkrsZhOCaO5+tDjm
EiVu4sygO8UDf0PIEOf9WxebJIoi/41OfC6wS0RwKh/pI3l+cxQ1FHGml/AA3bdGhaLNhPiJYHs0
0ppOhFCN99BjExG7xDFuP1M32cA6bF+04CXXgRIOYQ0OgZgJua+8qjPPZLjWOfXkVxE7SrhN0EjG
NZyyfpymGq0rtCg4ll7PP49VK27K46Dk5dPzgxu9Ewt7dItSGWa5RByU+IRYq6IjcEHlpi9aXGFf
pbH/Qpro/t1i+p5wTt7/FzBye81WO2Xr7lqgDi7fF4S51z9fyJXGfgXCsvqdfMc+j6GhIBtPATTo
6SoEnHduZlpGuDatE4IUxafhbMccssdo2dme2B/424GW3fkOiKImsCXen56O/MHaQv8OzK7AY+zC
W4WDjPQj9CfrlIWeV2ZZtdJ6iZ9ASXZDVU8DJtr3vJ5hvJVzOGiV/gv9y2JSJyULgYyDTzDJsDDf
CirutkyDcm6txY+b3srYDRiWF3APYnvKJo7FAnw/4W7sxV/dQnWmjxfmibr/s07+z7DgxWeJIfpF
Orab0tI/wTaTc5WtqB2zHNKrFr8JisjauIE9DChWhpsZ4eLG+nljX3GS2bzjIt8nNJQtiXd0rnot
9LCZjHSzw8oDRP38UPklLcY3uBu8HudSQBqhzChSIDAUv3NnpuM3Jw0k5JDRJZpHZbKsJXox9HOj
mO1nIpI7w5qEMxZewcOEVwt4SeoV5ek7uYycc0gQYuW4tQV1S3LX713wN1NZXhQ+1QukI8wHQb5J
21t2Ma2JaS88nKxy7S9oRHc9y0de0yHV4m87wPI7wJzuchw8P1HyY0CslZColSOid5um0Q3ewXqw
4P/kq9ey782xRH/PfGm5J9M4xbLj+02a7gqtOqpRo+srnROMn2msV6UxvyBXq6wO31CY/N7C6mY4
7gNsNtfyjvsYi4QwUul9p51jbWyjTyiyVRL4EfM6tltL9LbrGtV0Y71BlvfjmoL/Uc5kTYuLncTe
0Z6aSEovYsGO3YJP6ZGe0TcNSok6aNYZrEQM+m0dXhDf91vJMdho83UGezc9Y9KO3Zt0xpNYF5KT
/9Xy7YEIPtCphtTUMz1EptWKB9pjqwMU2EUw8UCg4ZGVLg/QWpCHDbx4+Ei264vm8Yvk7r8vAA9V
zz8L4qvWg19YMz7YF2uE3+VkyUlEc6ywI8oU6BQnFSD7OPKb4AChurpxXc6j3buDS7HFUU0mPYRb
ZERBYzomJFS5k/pMPM2gAzrUDZ3E/6VG9TyAbJSSdYNJRnsKGR4GRo8pJn/mzBblEqDB0gbnyOPH
WwNzKp+uZ10q4MoYDi4jmvUKH4Fof9VKr8A+yvczlM3C+VL5h+qoqTnZFkInd+FmPfqPpchL6tTO
w5+L8kFYCiOhk6Nv/bOXEsHA41NVQnuIrgNS+Id9YAGpv31LU8/a0zZ142aW1bZnZ9gg3G5j2jUR
0UejXGIKSsl/IAFVolLip186FzOMNp943pIxjcXTf5SylGrA6B+kK+eO3NCqpcvNtKE9G8K4OYbE
B9wFwe+9A7L8sZ3if3EiLa79E/vE3Ka9g3afDG9KxUcbSo45gXMdcjo4Halr7ODgkPMYpyH70zp2
OEQYpfE7qyJq0IpxFNtikwmR7UUoCSibdIGxHfqXBBAxDqTX8RNxvqd3kz2tz0w0IAn2ho5Bgen9
XiMcGjiHvKbSoXCniXQ9N9+DTz8wTduFImpct4tJqd+bn7cSojonfDB9MssnHJuU4MxdT97qLdo/
dmlmM3JZgy60W6G4ky5/F58dtWWRh8aCYFFn1dY/S3n6f2KZnN5H1dqCwKy+EmmFcmLXWPzMP4Hb
S4+1d7Ai/+dHA99xgY7bos0RTRDeVU66UiMaTE6TXs0qybmGTktS/dd7IcU5facpcXo9tCCfWoym
z54AKr2FgNLxIuk0b0q08dNzOkDPyYb8129BkrDkr3EkQmZ3Uc9lWP819B+ZJQVrmlcoSYeLbFoU
I6OINgCThxCme3xxlRHxrS82zCpsmPx+EhoR3FjTYfrcRKfU8Qb+yz8OCAgpGKNXr0YADDPF09iI
+6wnmoxrLAq0UeDDSYXKHGbElrUT5PmPYI+Lli4J1P+OS+ZaxeUK7Aq5htmH6eK78ilnHDaYUTCN
6QXszBtucxlujsjgq2EZAqchqkCxphzmZ8Pm4l2vsGOQr3Mk9zxpYcK7J+Z/VRP+iTHY0n2z4T4f
SdNcLauZ3myXAkatu0m7zJbTkvPoaaUebEFN1dww2XgNskDGsjAbnFa3GWR12/ghlRZHRqoht6DK
yqYfHuE6Ve+GSpWLfeNHfBfMJwDxorIArf+B72t2ZkaK17KXHixJqMFKp4EC2ghNulroMc1ZKIAg
OtEhfqYKAfCK3AgqGFRVstKoFe3a17Q444deth3e+jYwRd9RjgKPkuKXolHHjNzveryKlz5avGjX
nUffV2YdC0qhiSKcK7mDtIhCf6cMKUY+wbLN2Yii08n5NL7t47Te0amDgWK8fnIb0hGPVkx7+M3y
r3XquaegMiK4NVyUB1LKPRuUvV8GdVDdlbUTOHZ/eFhk467jpU3K3J6Ijg2naIDAtPd5YDqE19v1
dx9pcm9JSmFLqBLOfk0HwtMe8zzT/lQZK4TkIYrt7nRGC3HvOehvTepLnUeDZP3ilPV6EupKuzsR
Bx3AzD6+Mag51rbq6RXzNM26zuWMCRBrdpMZi0zY6QIGbH/0UheLosyvPBW57m9wBO3rAG26yQU4
guVBtTqyf3edJxYD1DL/T4VkYTAC/e3kWtUD+uOFWk7ZpvW8qdFzfZ+8qoznkHGF34z+z7O97xAl
1QHFv+fWROEyZYIEtdX/ZK2FDY1+9f0YATB7hyHpgCXHvsFdLdAkk3S/wjBzAx4zVZPX6TQyJROq
wK+RVrP0VqeDtXnlDt2eoY9z/h1oD5Cs/Jt/vyRN7/cHUkfU85r40dDDCb0a5ujMDBTECb2PRy87
1XVQ58YrKIkQcUGwPmZiWV5HtDCjZp6H/23hukPu/7JF7yeFX9f3qkcKtKD+yqjmh9JEcdRlmuR9
l+6ygvdFeWWUjot7pkbPR9u/Dvpy64rkycfACTYMFOen30oWRrVezzUHaQfkdu+xrwL7mvyWXAUQ
S37mxrlENYs+/VoKf9BbGA5HCKzdz4rY6cVVRlbSLsfjvM04LcNJjH7IRTRxzaqzLVUp4ltBfp4F
rl8EI0/rYZIU3vq69EOq82Kc3J4AgBOocBDfLYNKMDHOKrXlN1dzF2EJIiSJG8AabSLDpO1hp5C4
esvHdv1yzh4qcUHNW0fi+aHxt/JlfFPBoPYeTIIk31ToCgMGAeVTZ51dldZ3Man86jjTD1Kk6k/e
iqRnLSHSrQkcC+u8LLNVOpeFqUWkPM56zakgn7g/Z1unQF0jOWiyQvfn8EvNwxt9aIVdULzAifPI
OhKhitbLp5k9SnXBKdkKG9GHpsGOuR6yF54+z9f5wxaDmxVz+3R+yB282UeR84Sf94opwfxjZaRF
s1HcnhZnlnGkjcZQsh3QhejbJScxa52lVE/PYAkEPLdiPfJeKOvPV4xaiYR6WDgR1wuKCsUtl1CK
AmCUqyq33qyxj6YDIoMLYMxaJwE2BZOU+Pr4dL5dGemcu5Nl/MI3IxKkLLwxDDZiIT9nGOrgzk3q
V20oy7Unm0oQ26gxbWfoIkhqsEVUgVKJS+cEfiTEyO9TSmN+/mOFQ4UEt8meQdRk4X+tFSgmssm3
Bd1EFyb1ICEwietxfetfswlIapy6UyYn5nlvl+sB2Xlum/NR10w5CiVST8tQgu/M6RQ3JZVTqbp9
7Leab1GZoHgCEz0H4LUGYbGkUjihJdr3HfB4mCkmLmuA7YGiwQn8SZMKIARF6P6/IHCKVtJKmioC
GusoAQug9LVSWAq6RI9mfHc06m017k3Tg9UK2dTWzXaYucqkWBgQRrPNmLj09l1t9LtnR9/Mn9JH
UgwyqNMcQBDI1CiF1XvVdMlGhZmzG5De7vP+WKQPfGAxvz3uH8/E+0gQLUkZZi4+GojfR8rMMGEr
BncZUydfC/uuQ//NEmxE4sJOHbBmopuNex5+UbcoCxJplNhuLhkAO4yTfOddsnk3T7XUw4Xaft+s
EroCVeNzDwWaNPQKyob6t1kTxVdcJTQNZKMixAhgNbxtKCPjVQUcP2O2p9NY5t9vskx6RnXVUMRv
ZhKkbLebxW7brGkLTh8FQsSJfO4rxGyB980LCUBeOU89GCFG1IlwOGIJGpjyTTkxS8icyp2Edb9Y
IlqcdBd49ABAKP9YVEXeqnv/hONuagUzBl+VNMq33ZsV53PeVms8ju5XCbOepM4naU/SnwWT2C7e
QmKHP0p2k96T4v7duzSOPUoeaUoAyfF6cm85R6wFi5HgTT0+5It+KKyZLOPki19AFyXNSVOP+6X1
s0Xa/N/b1NeRJuYRKlK0qvX4Zitb57g7kY6H0HkQjMntwOdStXF+59GiODY09MmbEN8XAhbTlI9Q
PS3hfPbsCsjt+VZ8CjiFV0SpubvAkVzWuxWxWqFDM9Fy3SijwvJT9t0xptNtadDEqSGmajCm1ufM
urFTTqLfXrIer0AUWsY/Wicv/Ouxttpn5USW5tKzFX6ysogIZEGy+abvugliVULcqIC85h5M0S1G
wzVyLUsmlzpRAuJycuy0ZMTG7UYFkKXGPoUky4j+b8C7u5500z1SG1ed3HvFHAx/tHCcBYbsGurm
L1chG1W+DHAKdNlOIMAkxlsvMX4zeFEtR+EWGyyQFKzb0jQWdDooQITfX95OV1QWRNrLZO9flihv
us4e1VwgbfohnNRXvyAbDNSRrYRggIz87l4gR6dvYWlW9uMDOXAqCKO5YTKZBeRYM+DnibIjqz/w
Jyhghw4LtkpiMlH/8foAx/J3+dhoac509dUqxnOikWOgDf3IS8c6icqIF91rYQejr1f4YJ3iuvO3
1RdFRzcHSVEnuxeL2CstbUtYq6vBZlhPiqmV62chWwYIrPURwtz0Vn3oudN+NwstHBfqhzPmqQqD
6UsWgx29b0aOqklH/d0Pn20nFiFvWd9eogSRGZgBp1CPCUr9eFEsux3HZIRPGrmP+I9CYiSw6MpT
dlqXHwTZh/uz7Wzt3APjbhI3ATq/Uorc0bBwg/M/259sVGqrfjGOTL2Eo5jTj00YdlUq5NrnbnxY
6iKIULFeKtGtW+EAlkBGp1e9R8rvpSI4xEnm7U8ltt4Td2SXhsfVf/1gyHzMFlkypnV/QNRaAvf5
jnM0V/AMDymLji8mAoGOKhfzEtfK2slSAmFmLxp2vN6WZg9QZBrWQK5eNaZeBFqgk8xfFCP4DzS5
NEic7b3V2byR8JAhEg+nnCF18j8Q0MeEormW04Hrv8sZM3200Rao+X0WlexxBt8/N8mEoefjRZDU
nFdNPpFQ3IfIMkjqDSQfV+M1fGc6ffDJDyXX5FZbIbDzCqVWE3VzjFf8WkgwCHIjj+tlnD3LN3cm
HBbbW6RY6x6OHwhNK+6ARIlRabJuU00Cn2BMT8s0HwNckPDjt+VD5A07v/G6Wc6CSvyS2bdu5Pbm
1j4ONVpbED/KDAvmO+zb/jol//dYrRUyaC9VDqLcbmfD0hLdWHCH2HDKYPt3zZFmGWWcpkdd1MhP
olENBk2c1pj9tcFSUanl7wn0wIahsjZWCzBIWq+IrMvc1bSmodDpH7/8z1dBE7YtQ2hjsea0wujL
8BEodpL5vypU1uVnB/QPLBWQv+jvwqBxF3jW/tAOWS5/ff4XBNfVXsHpNzFeQMItummwawjnRnva
4dKfNUKZivuBvvxrgZ8kI+YO+B0UYOSLq9ozHvVsk6O6Se3AtEECJWhrh0z32gOLKSjxLase7NvJ
kvWOy9uBZR9ijshlLddZm0fLe3WNNcZxVPIKASocZzJFX1KWIIVDujITE0ypNKDbY5ME6zfCXp4E
RGly8opCkMAlvJ6jwP6qZb5WlZ3XY7joWJNQMP9rzlWQa3dLX0YQJWGN7i7TZGCwwVkLmkbzMsCV
bYPfZHwPFc6D3KaYN6eEerlzEaklFfZnr/j30uHWQwxXXAMKY7oBCTF0+K6p/iMZ08bWsGSFtHkv
BvmSqGH9cXQ4T7W0yOMEIBU1hQgHsS46VXE21gkc46M62DytGWj1LN8c7Fr+2YeQ575T426dnDDp
/m6JWzjnAXxttkKO8cgPrq1UaVP+anGk2dDiCvfcMeL8u2yqkYhmqodCzafP/m9zYRvX7od1LRHa
4lVA2xvH95d5DO3KorN+z8ebzyKeCaFooHwxU2ZD/WaHnxCV7XcAGROPC/BPUAy1zwiv/jSZKxf2
3JWOBe2aknia8UrmZ0qF3wCpHXTFErr3TdDdqsJ24ASEVn9sM+WMr53mOq1F3P0GESuIOZVR+8T4
AKgWB+2aMJxxdBhN/7sG9jw6+un5UyEFYjAd1TNU7JDRBQTAwgb5LNRQV67HBX9W1wcs3UwDNVzG
PavXdp+vHQTHUZxZhByt+l9nK3Iel6mcMxGWiTulPEpqlj3D/lhXIMmjCEZ/ZqyOblIu13fS+o6H
eHunjgU7CKGwUBkcTxvuzuC6deb2cr6H8FAFynU6GmwlNyAdeYTJ44WZ+1TPqUKQHOMP1b7XI9Sz
sm/m/mYxkgcwekZ7AsC+ffdZnqf8aJn+RHLrZqoSQaNO8qVTMz9S6d0XQCiSYn1qj0JXifpGhHYK
/2r4G07mOY2ZDaZ5Z+is5gzgHApQrar3qNr2z9HyNrWxwRx582O2lUNyEnZkfGJoKVGpYOIK4sxH
2J5Y2AdEeOEnsQkKXmjXqnZeklnAnipXj08aebR0+ErKEQrQW8M93h/BrXIbFsVmRhTWktaApSiw
jwP1p5AJiWLH25SbyCTPn1HQfGGolr4j9qSs7M9VVDbkYAvYcZxOLov0KfC4/cl1iOkGvBQzGOQE
I/CbbjhGY8pwktPqMXCyhExFy+kscMshmleTPb/fdrQF3JGz7TMK1wzKQUtsrxQwNcAt/2Rb2is1
q3w6F/YC56Y6ulpvP4B7oJ46Yfu2f8ZmsFCGtfWUF2t/H7TO6M/lZCAJw2SxjvNh+NdRt9L6yQHr
87iH1RLAmLbkEZR1unrr7WZ39sPrFNODjCUTvr5qlkqRrzuZvhEPC8kL5HJxqdrlbMSIVzw+2Zk5
ephlz8eID8hSkvH0H2o5cAbjNbyhaxMg0HRYNN9x2a8mBPRpKwJKtced0jkmSqeqSjAiaa2TDMNu
X4Z/iibPOwCaho/fYGVkgCBVNOvczaB0Y04D+/tZVwVf0mvi0paoDjA5q/ohyRMpI1ZW0nR9yXhF
Gxkq7Fk+o4pGtF3gXmi10Ix/hYEd9czO4qwFppW5DBZuTzkv+rgZs995FoFGEK3qPBC5+hPkM7I1
5qYkBSjS4T409DZ71+W/bFzxF2+GRyg0ZJy2QDtdLKL5tj1j9umi3PrFHhi8IfOD8SpMAoVyiOK0
B+sIgqgRIrj56sRcnl/xyKa2RfkCviDYTiFsb465iojHo4TC2wjIxzg5+qqNYPVxgoHhNQzktsf1
AmYArJud2A1MhDCUHFnsbAl45IQbbLKJSu7S52m1NzLJN84matIsf3WD80jZIZONvHazEHxnln5f
uvpH3schkkRkxt4I6YekGNxZMX8A7cjoEgFdmuT1Kbn3Sg1ZV2mKTRuMWwwG61knl2ddKDwmKAHa
SZQiueRUykp0PQvcd8tPgUtozZy2p1+QmzHmkdVglscqv9RMmq1nhcA5lm0IGGi5R1z+DQcVjEX8
6aO+mPuPZu6cEetFobYOz6mADBbiLVJBz4107VBz5QmwLhHPON/BmyTCP73NbibqOPY0NyvBpMvH
7iOL/nAQiw/D67LebJeubyt1hJ5suGS7GjYDcMS2L6Vxu+rn8HjXnY0rvpWp/EMbKxiZKxf2cEBH
Di5oMr2E0/s7pxGl9cML/dwhqnOKOXxkOMNGO7QxbwE8Ixg9KFKVyRZo83kusOD7DKGFOeUEvHlr
IK1eTuNhwA6F93XZGV1BPvKKE7Ds+zMFhangpdP3ChidlbaDnGxvhgyHXb1LwFVQqmWqLK7OWgUk
VZXxkjDvudR8JY4OAPOpTMpuy1Bhqkb3t1We0aHMXt+WlqaKtGCwZBEZ8KhLpCXvmQKBC2lAkiic
xk8JWMVU4Mh++oHh1GlPxDXeMC7Vp8l84bWKsbU4DRS56y1ymiRp1JPfSHKo83aXPiqGOomYcp+L
p76p7jefhHidBDpm5DAQZ16IMXt3J/ZZRc1GCT14KXEqmFEeODVZIMme3ZdmZ4J727fPeDL66TLD
k8ywPHWuWGJ2Kj9aQ7wI8eIoHG2wwcbWmaRnEYfHD78yhC3nF9mLS4eywWoVks79paan863fAHqZ
t6ZU6mgcvHU1C1aHWxg4aT1f72ZQL9n4oz3nlBUeRuzCIDpsj+P/6QaQE6z9Wy7Cg/n2gVM1smwe
qII+fh22okxUjER4NYHW3Y83551dBZn61Erl903nlU2sgjENQZI0TSsUiANHIvHa7ytw7B+ztSKd
tqoMTgRC6ShgbCuQQ9AGq9fWiAaoj/vWJNo5h+yRoG5u0Tn+Tz4Et+ph7bRs2QLORl8jyGcJG5VO
XE7Qrd9Al4EVHbYnk9EoJvLUE/GuBWsya1MgSdoLdykzICKNQ1urx+9Y+ywuZfHX1XCTdg8iq1lh
SX3XKZ1zEkBnyBhCZmSA1O8d2+nbVNP+WaSkbzWun7pYhgqQnTh4MsVXnDJXPs6TDQhEA4Som31R
OR7KRfzgv/c/H0BEMKbC+Eb5+1E0uOq6lOGO8R+/cjndJCq96GYFCHXH9vytTTFDB45h7lbJl/gR
efhlooao51fQZR70t+vjsVQtr3YJT7+lct8IRm4JyfCVKBaBSuxbY4H1B3H3MJiBfXhTdU9Pefxp
CmrU2ubx0Rxoq35a1lPBD675yNTZzy9XlE3f19zTUshD1srnsvozNQ3oXOlx4bEgyEqoVQ+fGGKO
CGXqCepP3cJsHdOG4Dw5rCoEzxj6LrYJOzezFEsvPCHb9YtdqZp49yKTpJP6zn1I33HtNfkEDXa+
B2SoPnT36MCaP6ydrjzD6bhL6mKEtJEa8G10jgGs6afDdrdmkq/eHcsjtDeTVi1h+hbGTnYFeY6O
wwzLWfLOiCTRK0j4Rs9C4J9d7BjPzAHshhV1dVCZmFqn7lYUx3zTLJDCtx3LESPM31LG7ZpyblyP
wA5VhrR5hkxFFCS1K34Oqd7NBqYJT2l+NXBnzeay2/CpL73FXkjc3H+xjOuerJadQ5wxbOBYZx7I
9GOno+fy4OMJUueoRXaoH9YoIzwDeS2CKX+3QTfeWrbaoIbL6n3nMKwJ2x1trj5V1ZbJCC0t4TTt
pPQd+a+D3XO/5x/XugkFe3XE5/Ed1gc/1qK9FKapWqtNgTzPELM6O/uFuxTbQK9tfohNp8BG8/kj
kqS1kE5HWZb5MKdXw/foQdzLNj5+jMFPcRS0xr1sl4aSkfC4l7KRWSP36kxZ1mUV8wTU2AeWHxTY
w3LzIQLgtxrFgIFE3wbY/m8yINwdiKQUG+YWj0p19OK+SNbogQCJTXo/Ay/u3qgBv+DbV20jUHxM
6acbEaCBDHlQBCNs6mpPZ5p6I8wdAtQpAVzZAZMHYzvhqJd9dCtyn2vOh4DgM6uVb0LmYQdh2T1u
6GRyY6Gwgqah0lI5T/G6VtvvpLqPqILoZKgGRaAKKPZDfnhna7mvq7eJ/mhVHr4V0OeZ6XaQ9W51
X2vIbZ9y5MMAHHCH33zJXfRZAO+0Humgfeoj7wMh0jkbdXR6y/datlqonxgCEaHYlklfm5meb/2T
2MU5hgMA0+KraVA+x426KeevaaABY6Y0FMAxO690pUQGeLvXuM8SjhJt0WkIPJiTHzPm5SHvsc4a
s9FBiwyhPYHTpc72Q5wqb95wpdSk1RMGnmIxgZmUlWVoc1XIjTHmD5DOM6lv1Bqhvhl+4Gqvkxi+
YqhWZ9iphX4SFew2YnHmQIN4gIGd6nT6JjaGfOd184FII3CrYnLEMQ+o8s0InRMqPMB7PRGEsDi/
RZLmVA9nxFQvXWKS5CWDjWx+YiJrc7aFz693IQISbNh4m/Dq7FPiP23GwyD5Je+tO8rQ6MghAcyF
2QU+rWMVrOMDTS04HIWKN4SdEMS+bGoCufx4te6jIYsHofadvMmkhZhx6UXuVr+B6wb25q1xN2f9
gOHTi+TymqrQzBcXdrkQ6pCy1jkBT8Ng9qF+nqbWhNWabEeABEFdciqU8uLKoqzGGTTB64POft3U
8ReS1uIdW2CGNIF5w1swKxsbG1fXscM1VQ3qSBGfxG09G3TfSeLPZSzqFwqU73gQhpsTdrl4p6U7
E1Ra+P1ZPLhb0aI6qy8i+kZSxPebSIa+5ehwhhQ/hGHKVnHfS2FNa05uxN90aFlDwq3Glg9texVC
r7bS3wPaC8Cz9hHQwDwuGBlCHl21e7xFKJijnFt7RCe+YCh18JS82rhknlYl6vZsC52a24AfDkvu
DrrofZcc/93GWGVniHGdFz0uAkxwzVqtAIW/QcBiHI37slVAoR6I29pywL65fXfigTHf3X+t3lEJ
XbaGZoRqLsK3YbwHuziVSMFBq261ojXU+u8cagQAt/yql/DYBjZ4gL49lXedhnMBgiLm1k2/5/Bf
bmzHIlG+Oov5yw9edAvkkWw70W9tPpHkoo0ZfurJsuPbCLD22CXTxoOnQPf3Jr+Gw9P8qJkouMML
IJQNy+10cCqyBir37Tb2dtZ0MaFDqcF/1TGurQJtKmAEVS/N+osFLmD2qwdlKk/jkLHwcaEtsWBS
jPeE8ZaN0rWHZFQ3nW21FQ3Fj/rsfUY914x5wbmoG7sofLdtYafXbif6cdzvMCCNyO4YjQ3ngWDV
9GPQIM3jI4rN2s7NQOBnTcblCEhc3JdKsmtBUroFa+KE4RxIOMgFy+SBe5qETTU0NYlUChRZHfmd
v7Wp9MZyWVZjOKxeEqqAfpzUcSRQhgsgYCNBRgR9VCMFBEo91pxV4kt1fKwpDhz1+WCwbeUHzyuv
ZdXP4wgwk+UK52Ja1czGQYBNWoEIx7dIp15Nz6prJjTnswHL3AWTRjQPoiqzbzVx7Xg8dPaqYirs
+7riviy8EPV6HDSQpD72h2ZqsueH12wK0a/MIP0cHPDVUq2YdSeYLPOJJY2lSNvjaNHUL+l/OlRV
A0MKFIJNN/kB4HTVFAdEhWa5+ct/x+Ll9qfBdD5TjspF+McBemnqZKLqNyBjmOf7v4kJqnVKM4rQ
2k5dBj36kz/hgpU+EMQEfanxsCPUwU6i0d0pNtktU7gwaKhiaO8rOKr11pghzEc6DmvXKcwVHs1b
tVL7LhIBfcJ4KZLtV/jtzQe6FQ+c1lf5RriTXguL7ggY8IWZ3B5XV7dHtOOk/DsBXzFBPoEKk97b
a1Jr5rvGbfWCqc3jcrO8a3dAUZlGat/jZDsMnTpwiwN9YZUrHbm3z5nhkQ/RTFNqh8WURT2FxuxR
Jhg0WxjSUSnclPtiW7Vd9WZhZjO7KoKxSeNd7p9Zv5vQuIOJwUwTnCyTXYMED7Z69E4E95qWP9j2
Wu4gZ4Mx+uf9V1fFTD669/BYfPbYbF+OzG0DIHiusQU+NT55sHOs4tiPDdecmlzGZTpN9JOy8it9
vIAOJvIHukaemHbDvzRhA5HzkJeUVtd7iN8oJDGl6F8y4HlNcm+eTtlHAjanh1O2qoIOhyY4H/qm
qhbapwudRjKpUct/tFe+L4YJqtaiq4IuGtq1vkWF7FVkn1aNLKsopHQNUU78RY3H8p1w5jjWRq7q
T8mbWLAL16FiTGhye0YkdDQWKy1rZum4BSjMQLyCDj5IEx6JO5PLpg+R1m4hLHafJ2wKWCUcHdAK
W0glZ6UXHHBttHp+4kZ/tYNM+aOgOLJu3MSzgcyM7zttLJmNWDAH63/zKNxuk+hDsM6l8f0dNhs/
noTYQrxTTIKumbxb06daSyrRmzutbcST5jhhB4ZN2MndJZADwb2FAdlHg1P7dMAY4/dNJ3QojtgX
KU34OFufCtG+EAEb6lE393iq8myUH3GAwS3D8hpfiQdHSAQABzf8t+mZE3XlTEMM2Ll1atH3dDT+
oWqqCWsazkrh0zuiRtajL14cEbFvxj6MEgc/7ucIx6U40Mq+Bf2mO+5X23o6VnZC+taYOy4SCD4u
JIka3I7Poljlm6JvRjoTxFTf+p4ctnqBXCH+0fFKy7KT2ipHBHN2ARp9Exr69cLJESl+SE0YhrDL
xdhnp5omqyyv8KZZN0zPZv9hMN4V/RXdMlMpFfw6yodLG7fHr2fVB2O4HQzM6vjNZLLZTEkklKUr
GGrF4ScBY1+Hj0Dru0rLvP7BUDs0xf49wiu4+9hIWihCfEXiGZDzUeLOdO6MCJTYXNPo42ayZoBp
w/Nwx0kuKv7f0WGNpoc/CMAIalCZQfX6wL3zN+MeW64DOPEQ4wHAS1kAO5THyNoeCBiflhOKnbx5
qi2ElLjJPq/9m9pjVGbJUIAkTEmNTBpT/eY8KVqXFl+3VdOaoNtfnKBlNnz2hRZ/YrNFarbhDL1e
EizS+Ha02GoxzAZYJ6g2rCBUFTsyUYObN6qx/MU/mEFtwZeSivQ1kTCYU1epaXptqHDUQmQrPeQH
C5gI6K90VTleFy/BVLZSXa5f6gXSLp3TXcmqSvHHy9ZQ+0ctobExDYIXHXjVjQTP9EYwlt7FQ7fT
xkq6OKR/i/I3AvQwDsm92SscHsMo5tAfhwY4JrmaQQMx/4Qy8+ABA0UGzKYikltMWbAp2kv/3ZkT
c4CE1xRN97dtfxHm8X1CImnGuKgtEHSd4ZhFG46OiM0m0acRL0VRF72gSnvq1RpHveAAXjZhAUIL
+3CO6d/kAUN22znqlMqcnKT7+ATgTf+O3fBwmUItu1uMnI8U0xOxRbD3O/aUnELOyfwUKp60ydaJ
8xYKZPeesX/z0W1H4l9vPWBzu3Cbo9A5EtS/k4EwJgYR8C7U/dZ9Z872xZYmenfbVxBjQgbB7zmQ
aH5zxURWlty4pksFyibTFCtqNJCT+/n0mI26JzNzW/CFyPUECGGnAIOtnoRoQKavByLvEl1G7+0l
eaB+MytdC7g3yAi5oH0pG5/Y5awyEMjiWjzatYsToose2xYisTjRrYpxx0d7X9n4U8znGA+l+2H0
IFU+pfgJY4cep/WDlh0vA+xHHsZ23UpgrBOo11Zrb9kJQ45GBFFCZnPoEu43fy+sUsyf5Ekc3kU7
W4Pq8INfxD+VNlK9uwhfzpUMVYUDeCsNQzMIyw1i2Y8Msvqo9o0PMR7iiv3LcTQeG28CTov0X7Tm
Fyo8QQ19D5GsVqltp8YisyXs+8RTMlu+xFhn+04ZrTQF/x5FagZTZwvQPrk610NAmS4MTvgUpiuM
756NvO3b516tlVhldk9jlbCV1cPdGcKwpJaVZWfSxVSBbrL7eiT0IoRqkTzxYoJbv6QiCebD4u6d
OhRmw8mIITyteHR2wUNIiYBNmtCrIZSZqdfCrdwqiUxhJzd7AAla7ToVDXbPwElBf79KkTtomyN5
q+gcDpmTmByZoif3m4V5Sac5usPHGSMEypuNwr+5PqV5m2q3IPEuvrljztC0H+QlyuL2u0Vmf60h
XFjvlSJx5rnM/Usq+XnsPxVvSQDXxBTOxuDdgJ5vPRJqa0jMdImFGqdNmptljmPSHf1BhvW7NSv4
9yjFshp3yN0KJLqbAMX9+oKLwyknv3nEmEw/W4+SZ3X5X7LeJVtoeble1BnyArOmHs13YGcOtPtf
3oJpxMvwXdCKbXQ+zyN3djRq/R6DOHZ/pQoQfGuHcwpDUygnkCyZjWW69rPYMyEThjyyFSMHYU94
W8zSGA3AqVxwBNrZtogW/DWiHkup2FP3DLEL4D4hlpyc1fH0FZhyjy4e/mBZUGEhZioKgw1TILfA
0T1Y5kTJ34Bk579xH6RLtQ0l9S+PvUoNv+CtdongGUNpOV2DnPy7tYa3wL43gB/qwFyxsjEsfvYQ
OLryHYJFboPsMoFzaqRqTGNGh2kqdaHwX1DLr7/20TqKTnGAj9pnejnmQVYd4XLZzRq1Un9KdCva
Wvpd4H2SOT8LvOiou4HpBsVaoOmh7DXFXAGgqyCbTwNznE1ybByZirolqXhJQ7oyj52dvaox+Ja1
WdewNhAnV2DSYHyiIC+s5QKcRixKjxmujufnyIzWC7RREFOS0tgMgM1LTgC3s/jQN/LkT9g5CQHK
SmsAFxVhbHOIkrAHlSicH60UJwczZVbRsy/EmEqbwEs7VLuktJVznnNso396SZTmd035PgYPJXan
2p4actpAxclfX4h5kRX+S5YTbFHfz0W7yyBwSPc4s25dMiwRkFdMVaB27xbGcAX5eoc9zGixuMjB
G9glAJQgohL1zK4cBHkKykilmLdxih1rdJbFn7rtlkDYisYIONJPq/tD4x1iUgVE8Cjqfv2ljcF+
q6m1j6ZhxtC66rQnKa9FTesn/Z8K26uexPE+droe8YKw48eCFZcwhF1BEgreHES86vAJsmlVZVdA
LYbq7gWCyKMleT3vN9hcqENfRS1aEqGGWWtssMQLmcHLoO5uauaF+P094m/z5t4TVK8imHR/Ds4P
TbQoNYWFeUDirW76mP9E3XYsWgfZWsloW2TzaGsbWETdR4ugfKX/kEb2KLG+T3SDwofEHm6sEx82
c4jS9Rdds2sDuv94FSy4soLJvO+Pp284vCdKH98uPQIMURIdL1jjNv6Vu7kjQNqvAmISL2MqZHSM
E3OyZ/Ji2GRg11+akM0FOJCn76amTNl8xtaFoigd/iAYLwiwpCsCBxW44URYSlP0KjmbdpRnWXOO
Gt/urmShnVDb8IOVQNM5o0Xiujvu50ojcXLIpg6IZldNJDmCxx99eeBCaUcjV6Vi5wfviXOYEc7X
PIHFnsdG/fkvAWQkcZWYj5woJEnB0B1Vj8LaiuRJD5r0Kw6YdiQn1nf9cvJRCMPE890y4Lyu/wKO
8njbv+2pZ1Q2O5g3QTQKZzuPn3xtr9rDZciWvHB+eI6kxZreim9ZofjWs2GRONP4flmFDw1sl0Gc
mGK5YB7JlRaokZ9iHxnulQKvmerFHvVPUMf7ljxWJfNxLdLq/n4NpNt4bX1jalm4ExTC0bQkJUmj
Nmugj/se4eC2wjmnzUDANWmsQeHnKQK5YohhBFAYzHbaUsIEAgvHakwIfp7P3/fs+z+IQ9k3MN2L
Hiq27ePsHOk7hFxcIw+1EPtMxD6b6dcPMQryY6RFbQKUXxoANVhtdQrMnQyPZ2slwMSI4WnpdfS5
p0BVEZCHsBYzmixkyoK77csOgO3wABDtnzggAty4JEH18a9obVPRSHHKQCjdPnYnRM5B06xGrOLg
8T+4UeuQ2T5UjINi+GicDMiNlF2e6wf/VyUULs+HuxDPF7h9ph9sdQD/TNsLRvEcw/LE5LxQ1EUS
XGKUAmNNyZR5eyGfbtWEAY12K9ahkVCFQmYyDV7lBcHU2u/hcGmqdqVLcUldJU9gOuxDvmxwav6v
L705mJlQKcddoCm0YvZ8kXQgE9p8R40USB/chF/5BRUzwUCQFp/vp9FAFXJm2Yv095rEp7B4ZA2/
7Lp4rjVIHuAhXFJ7eni/bZVkiZbEWWcj5vnL316a0l7VTO3HyTzzmEdx+VJuEf6iNF6pxWdiPEzu
UcLlRDx2igdNFm9XlGLzNdES2wircpHfDEOPvgWciThuvJVjHMF0Pndi7vW3wFHxlZ0WaKsbG6ZQ
H2Lng6d0RqzUr5c+8XDQeOpteo5reE49psQlnf6kZ1qk9YXLKASKDzEe7JHl8qnUqM9l3iH6C2Ln
z+D3cNQ/hYLl3YkftxYGepDXLS5OYS0fmcOsB9yRsLGYHaWC2KNlb8la9GWJ8BK8YuKoaYXcTJaH
GOuouddJB9DJQ4Wdw8rvZ2Fnlu9ugDZy54kD+CuZuFQs2To52PPi7tiUvJspnsS3H55XSQumIITt
x6lkfHUwGUI+PWN/lkOriMeLL5jKSeHYbsYBGArULBNNdJaqXoMql35DpP55rqq/crbAkBw7mK8q
1FxvFOEpOahWhG+Yinwy4ASyUP5VdoMH4KbWu70SmloSJfyTOJWnlCIApvn0FybYP/gIjPSUznKJ
blKntXo3uCyDP7ysfaW4AnzeZA3bb34BSrfEpZrbwyyCU+joX6TqmRyx48q7FzyhqfLWoCnDCZp3
0brhlk9FEsFMQ42a7FAdQEqJYhNcKlOjWOCOcbWGwJHwQbAFS8mcdoOql2jhDVJZPIv0dPR+CU2r
kkZKyBaREmb4VKAu9kYt/fMO6z25uuje1jCZx/YWN7q3nHkegRcuPcUIE1JdRwMED/fH9tkrZzph
uy1zlxLa4FEXcjPIJDeb9yC7F5etzMEwo2My+ZQW8j+wvXAxPAPDIM8wjc04UR7KN57jm5LK8P58
Y1rPR2uMpY0y4dbUaUb8SPnvKpy/ciX4oKRRdUceIracLO+iVkuCt7FbY32bq3vlUTme6fJT4bmO
mvp9t+x26z5vO+72dJS9iXhoYsHhyDme/PWCZHh4iY1Ke7iqbXqDO76gp75JdUvxiPplj77rvnka
RTSB0vJhdqiMzFrAb7Ki9syUG+X2wo/6ke1LTIaKGYAO/E+y9yZN55mWny5gnE2S1oX7YRJasyOA
wAM2vO0DTZlFtABsM6nKkVlAQVPjwJWM0dLIvq9AxfQejAVYoSuV5SYIev/GEC8Wn7WHEW8alw5k
wRuMv77sSrpeCnT4rI960ph5if4jrwskVyGDDraXhZ/1/44C1ig3rCYdYumKU+XCj/ZoLKGcYNg3
m0G0umcbGsmNQDEoF/e0mu75uC4QFziuafx6kN2VKh329hf2Wu51fCEIb9Xdn00nG4tYC66gF8FO
F8pTkWsMrVnV60DqWQxMpan9IbIvUatcnkb9WgjzEZ/AW77TmE+oJQOGrxE0MmUxBglzeI4dt/es
pNEqogVV1ZjQq7pbDmobGLJBJgPSSFVmOrBo15NXSawoB2JjKKq0VHpRunYbpuaJ9LpGTshs8xes
uhTO2u2ofxQS2Pip48qUuIvShwfXZ9DGUBMtsxQu0BHH9sGyx5M4sdRDwybJ0ov0iu8VFnjH7oYB
Ogdu3Yj9hr9fePYt9Rs6Sw/nsITDXHuGA5qCBRtF2jy6L93UlXbJX3WT4VitLQwfKHkJ1bXvQs2P
O8WaLIth/MGQu+a1KkUL06Sg4v/DJxEVM3DfUR0ESBA5MbemCsR3mfS3+wt+e702t2HGbyQ5j93W
dm68b45Zkxczq5nMpVfeXIk4VY8Qm0il+juzJNZqpScIWjh+f8xcaO2OYg93t9nEctwHK3b6IJ4X
1mcKKTiVqBgGeUfMH81bylb8Hs4I9hDJ/A/ELZwLqJsVxx/yMEDYTUI4/Gh2o2dgy5P+IxqCdVZ7
ILsbfzDp74GbellYYxG49RdTEEeUqnrxVAEQ539VD9TILkdc7wY5PONnfjAmrbN4/h9KYeWlmLd8
RhXkM8uXTLeBmumRXRvng7l4CdtJi/8zX8mNqk3EzrmGeT8v3QcjzrVYklxZeYJtlOQpkAq2Hb/q
HImR7OQuCpUVOUBZ9HDTJzJn0qc1uj1jALPAe40KtMU5ccgcyFofqo7ABiKD8b+VD1LEWRnXaVdg
qD4X+w25WANt1vgKmLK0JQDF/FtI2pGQlvmsYd5lcOHLHIbaK+IEIzQLdBeQAiUt4FGGSBTK/GXq
tRsDRow09pSN1+DjOMSnTGQRGq97kvHHV6B5JDEY3Jz1U9/4NHbkZA+9t4okgt9pOYt1XFSpGZf6
CHZ80eMhC6A9jq06cpx12ETJgIddlaVmE8uO/F2+X6RTGVz+9TzoiluN6kA/mFlVYgyBOAMjOzJo
KB+aqJhPClBYZ0yXCbbaPbuIBC/GorwDnFnVnVWbtG98RVsrE/QakJfc5ekOC6w2v+loTK418ubb
/I4eSZ6lHndjDlV4GCDYiYuRTgdnLgy8l3jz1DWimzQtJeW1gX2Ys8UbLH2P+O9AaewbNJohNIuG
LW3r17thnCrhBDV1in0L4qagZm/WIDHj9NU5p0pUi0iAdUUAloRk9gPk/VhSdt2NPQn6QeNesLoP
t9cmg6JNsJhBKe0Dqr7taS9eFG/6deRsF/9vj3B7l2Owe2GN8nX8FZz8FtQNQSpo254SURpsGrZA
eH7QeRV1ys12qHy4WAm5cm8v6inPP+RCGnVUL0bGEbzmFptDvkTLYiqKRcfJ71GnKfkd2CJHPkB0
ZIRJQUauLndGOXd/AeGVjAT3bikPVkSJCfEJ8h2rKGpLM2UF3LGmq2VmxSBfbRL33Fu6MS7phxqP
twKyPdzTizCndlfVvlKTQBLWPT9wmaFIa9OgLVKiZNsGVejfaiY0H/T7b9IggOE64dvRpkxkaGOq
wUdLoSx+s/f6MUcw74xHZ7XRl1dIzRFtjq9+U7m69MTzFYw7usc5q4gJmbIHRUXesJyf88S1ufqI
otEDE9e4KrlHf4tg+2uPR9tNulJL3vSbV1HHLs/sptKOsagVJFzgUvFSU/6gZn+9iEQx2MEW4eE3
vMgIpVtFr3e7jgIylI5SAUeuF59wcEj7wcW5YTRY3dU2Oi4fl4FP9dUa2Ya0NPfiDWQdDvwofsHG
RLkAlmdNI98X8SDXNelEVZ/exP4w8Ewlov/o+LKAhWtrEBB+/DGmU8T76pgwG/dAl/u8K7fjAr29
pieq1gJf2RFWXT++9rik7dhITT/+pZsQ361OvXfVguovqd0sirFsKSlpT2lWppeiNRL/xlroajzD
h6SQu0JIuEcGN8Kdw6JJvC4ODuElBhUxBZJ1tdveEL/OdLbAWuH1bOwdtyKyRqk7T60t2xUSSZd6
MGZl3uNSZoFkC/mmoF02fO6HcgFAOJWBlHUBLlhOiBWRPyu9hkwnqD9gp54gzIy8bvGbRhk+7uTt
Yg7PwsRttpDXZMFsF4AtvasPfl2vfYswv+GDhPQkQjk/SoJyvPdSRf3joqAKtaUe1DzRwVrS04/W
KwkaN7EHyTD3SrTs/uVr3DFVHjzjsnjy4RxEWebD++DR8z9cEXyDuegoatlDOspoRhUSdh58MKkX
dr2NIU4dwc7fW+zqdMhTw2R+YCsJ7IO84ZJ5DX+PnWTp4X8dKWTwDrD5eVtxcr2KenpEjcQGbmJg
r2JCQ4XUsgtRWqp7aTepBLLtRzbC5NlXFCN0EBCyXEOHl29QWgmMMzCCQf4Kt6lNtVJvo9ygq7Gt
33s9tSxS0WNIOHiNLFyYp9s2B8VP9YCtqW5vbRLsjlmqEWbSJf6paluorr+yz2enO8qI9ne/Am7t
/wPywsd87rKOAXocbaDWFlO6wd9tuSKTDtObe5AWAlAMBP5ol5baf3Ke8lrC/Z7dK+yEbuE13YvY
kHIsRY6W1GskGnJ6eGkLxYSOfZJIH+bZiRFSaD+6ml8ToPdBy6zP7QnV1lkuAjIR0LhutrR08ocA
6bxHRjYRlDWZqw55Vg1F1zzqncKUX0iFExGk0HSEbgtaSBtXR+pegSSP/id4z9dDzClwihHMCuvo
I376LzutMoIJ24/i1n/VZgp75kLXnjNIGH74NxKwDTN0DCBoKV+QoJOs+7rFjZaYNOc9v2KIe1Xy
fzmUoJEGhweR+5KPVgRt1AgEg/hrHl+/Fhhrxea2izUwRHRgaQd98/zxGEKumvomYB96j5JbJqTY
rNKSqZUmiwwv4OgvZIHIGoHIX1Blb9hMkSCe0D6IX2+Ppgpx2Rto8BoY8s/+3q41PME/coWlUI6K
zgCd0W5kd3ZKDW2jZGGb96iCizCgmsWGfQDDLl0GLj1KO3CEGvO4IsjW+DqrAOlWtNF+mDJkR6N0
cO9eD6EkbwqTkNn5K/a9WuO6Qza2gBcURHtNXsMS//AGAt42TzzC9cZQa8Oi9ooDFyV54i1veyQ6
NO28O4kcK9/Zq1qBPcEzeu8WTVedOblIzatby29NmwKAd/dXUy6PEQpjyQ2B6eYwACNYx+87O4Zf
upGOAVhgmkFbFZ/Z2p/KDZtFffk2TZgSmu9hL+bj0vzK4Yt4wn1HuMwsEBgKGEBZ2mdskpVoaeVP
ovufi1CJN9Y1kZXagslMy3QenhWbxs8qZBClcSTR+YABflPfmqnENx1i2hayexqZrQ+C43FfYj/b
82sfAgQxnquC0BVesgmZy5/zSNzEfpyiDbfVSzQfLCRosEdVmF5/2Ez+muZqNsppWQozz0Od9k3U
y7DJstbPUns+yKF1A3u5UBMh/5vZMxyweKFIH6+HbJ3zsgJj68ETHrRlMJenHCxo/IMOEHcj1h7t
fM0ClqRRiu8Qfusb1jH9ee5+EOxmPS8eOkutsm2PCAwp+oFudj2fsQxLwN0SmyC1E9JBOm0Coj3d
ze1hsexEGkJGSFfbrmYI/LQl3BS/MrPmBZE+whbNkPwGjo9e82M8kerWVGG4LdzALJlemDvRtT0y
ylnJSAtFcNZYJS48JcsaFoSKYyvER0N5R49FAQm5Bvyrpbv8qurjASV6udHHVcJXyQ9vbkeQiYdr
E9n2Wz25pFHpDdcEk9VZny8lcso24+1hn0jBZbYngU+rfbJ06JwfE5dgaDmHXuWg4aFgpIMFTdxu
s7u8oXjy7agxjbKGTbHbb5uo9kcoqaFg1KM7134uj746/arbFdiCFBHW0BtkEzahKSeE63LZwjiE
wr8gbw6+IvKehSb9U25w4AXP1Yd3MYiA8IrFWIZ4My/tM+s3XZ/WHMyvINqc5qvyQFYJii7sfPlQ
E8td7Wvb8yvT2OnHj4fiDddLgxok8ITOCjx8aSfVqysocWuYHy+vXUXa/+r6dUfDiQ74PLKegMN+
DBAjHTudlBgMpc7LHqg2xSQD/tJca/dXv1pCmddBf/56c0r0Y9hdOVeYDpU6sbe90gRcGUmu2cI6
PzDXQLgW3FyI1TIqc2HTh4SirwkL0rVw6Kr1GAhYWv8W/gjj++ogLnuXdWRNLDjm16ji0xDajKhO
Yt7H2RXbz3Qq0qvsGJZZzfJ0dLBJcUwkQ4zKV/NA+vMKNEOtftirfXSh+T7ZtesQ6yebx30kLKjm
5dG+J1XI0AEtLvKQrTbRPlZuknjbVbf3u1hMGkEQpXhYcLT3wNlAK40tSNYwetzGvw/zTLEApGvi
+aqENyVCywLZj8jDLQeQESCODXl150OWMZ8o8yZS5fsNIFrx39b2e++togrmHyZJRV5neGPdFBkC
DIm1l3XGTueynHV2mTG9MaA1o3giZrYYvTkhTecOLeoVDp9OADm9z90Fxfeu/+HunjdTV+K/3ZXV
2fARszlzvw22jyWE5dbhDBNoIS5ZfbyM7UT6Fiz5i1paR9WBTSahgYyX5BhxuPq+Iwd5pdgnDg75
g0y/KNADaN6UCgr2QNHiSo5/rFYD43RnPcSapVCbohs6j+MLdW5qyvjjQ/xOCzzqefdMDN+Txcd+
QQ3JVg3stxRTd5xmAlPAYdhupE/+Wc6x9b4qg6mC2ezSzRuCKasgGysikXAoZPOvptYgeO5q240m
1QfmWFok1biJBULy9vmUdEX6sRzk+6+Fa5iPlCUzg1uLpo3Ib+nZRKZzBO+7csVE8SP96rptgWOe
SpQGxEd4t3FQXG26HXy/z7ZqArOMjr6yuG+P1okVmnQnrgqJLQy0Z20sfdc4ztC3jl7Bk9Xh9NCT
mImqKPf/X+CCp79kIHyCNONnwH6KzJ5wUdwZzKh8jRpjtyNOXZLZhZ7xhHF5hU2GdwWkxllAU101
rzcfgJaIRab9X72B9pTZuEWYHmSfDKEGYZvn7P45MEtv0XwA1kNbmA6YU7u7inwAK3cAkWzhVG+F
+TCdY0Pgn50LCw+uhz07tdJKutwVmuQfYTPmYz3hZFrXCiWOSpbbDE5FhgnWtjiacOZj4Zov89i/
WbD71ai5Z0ZXsBjlxNU0trAA/siCyIaUxh5nH6h5jVZuscCQBwHgvzWkyX91lXrRTfUTgzqa1c2d
vLwujEQcAOGHgltqMYTclXsrGrapeBWPRlNhmYC5w/TDZfrFhjrrZw3dK7pIBKnICgwatxqKZ2ob
4BiWRC0MPaTWJ1P956V7ZKGB5ADbLMbruBUuHes4oPKV9wf1R2xbAJmUDKQGdHfxbAXRTGtkoB16
04ci7VPWZY3uMm+KkkfwXWeEl8FkAjoPaCVpoAqTIumwLe0isL/KDI0jnduRZwcTdem3eJVFf4al
6koMbv5DvQg+Qb6/8cfz6/LGq9/C2p3wooLPNR7yfc3IiTUBSq4oGysi7eAUVk0GxULkl23sref8
aDOZQk1hGewQAhldAq+j5tVyawP0ajfCzJdzHna0Zl9OcWz0eT8cJlgBQpCoIJZFaokqoU5XqkHt
NnAKcCHIKDLiGaow10jvpMXeHmzMGTONrGYgqeSG35ERkwK3UyAR+MGlF53XeA1Njho4ddPC53xJ
XFpkBg4L4ArB1mxfAhBGpO+SUBmuij4hJATbkcuG8Ge1SWmYvslXybqZTFR9ZrmKwuW11+ULeTb1
KjwfJZPU607ENkrNAtj4JrpeugZwRjLg8Pgzh4nMgtGD70VS4BAdQDRM6im4S+XxhiFd0PhOquO1
KmlcJge82a+PEdu0xlzAsx1g8FeT32Sx6jl/ZjqDpb37mP3Yzk3Nv5qWcKpjJ9gJwAtauV6HmZy/
4SV6bJp9uLQr6jRG+I9nKq6bv5D9qD+4kkZAqEUIwPUGFUaAkoRzkuc9+3VnMaPXUYIHQNzLdpwP
UgZAT/B31LhIwBjJztBhSu7zE6FS3B50O7SmMqoEOmoz72TMRybCiYqGbMWYfAuPf3XCWUPSGlu3
fdhkd4p9IRpQaId5MMZJ+RCZ36/Tz5m+VGMdOM/ZgNZ6IjAEyPS+FGYea2Ql+gjbYKyNeCgpBjqv
Eu1fyNdlKbAHtLYETjr+p8gDIyVy+rDpMgWdyekBqcVul2d6q8GGzK2u/13tLM46oxnKORJyShTQ
uh++Dq9Neae9Kbo/FbKo1Ez7G1EIo/wnoGOvt87ttZSfbKZUqdCtVWCTbBoVBcgHxSB/yrS9dW7q
vwKYyH9fPE6prIZWJgwyv1rPHH4/DtE6UYzDNO6gbrTUxqEcuj3i1v3RHoot3EwPslJ4r55RSg0A
aqDOdetUhqrOIeGxzZo/sb55pISL3vBQhCOJarIzK2+UBRnhVY5dTFS3KAXL8pXlTmIOgNjNL8Sg
jXMzq4lK4bLHnz+CBu57G3RDjxlxuecUprfXjkM+TiKX/EIikHr54gqdygp7cPV9u8rMaBfgIaUc
dpNpwxprzTvmi1MSdkPgenffrPcl4j2l7rNAgcuk3XIQ9ZpueF13JHsyCYnX8AlfkgJ9nlor3cGw
aWqvsR9LrSvcCnRqNryy+vxd1vct0yyq/mohYw4wZI370bdiqx12kH3BGV+ed2khfC5NPoz9sEM+
EDdH22fS2wcGFuMy6UMkkV203nwNG05OrhyryUBftBRa1gMJl8C+GstR70EKY4nQ+G9rrAPCvztv
lMvoFtNlgReTuh/VhPDktZn0NwNv43sFuc29QHYwFf8xweDKT9CQIlsatb2vGR4zrilJMq8uH0bE
6jKL8KBpslA5ZYnjEIwUJjgjZdUgQdlCDonlxIC+fb+pWUhSbMBJlRe4+QzhYd38fStWCiB6L9WW
eoex/gCMWM5G3aczWuna0tLIh/4VEnBFoGlgKk43zvJxtQj8BddbWwL1DV1leUcARnB9Ro+mid4x
IxmSsUgMkYnSFS/usYsoduADbPgO0BWR2S1TnXpb2pXeA+7u1CbHffqaofNEOqp6XY5WDh/RfpB7
SOgzys8G9pVwiiHUdhb1NnAXifAcG+xSkKhSc4Sn0psqC2DP+g1LfaeWO/bB4YMG+rTPQWDmjvH6
vXdnyLWslUSkobSwn6NzZOb4xkdW0lnbsxlidyfxjDODgwheRexQqq9KznXsHg8x21deEhfhwv7/
SFDeftoEJzRmujNmTdm87aMxLJO75YCwsLadhsbs6CYfranXUVK94aGTUThxB9uaXZQBQD784WW7
i5+l3unDLe8BpXkdjrdPZrhkbtvF8Ln8nlUCWOC2HjiI3i5MG64QJtKdEMxT7As9yVkmL5NChnRC
znpdWKRAYhoJGBth47KjiXxNmOIEdkWJmepKZudVuAP4efjU46lwFWHHwWhMpivWDCIhtJb7REXb
6PSp/palY/v+Z//cOdgeTkN/yYkcBCiHMmh9qj9ii57CbiQ4kuBdDVOK+JS4HO6kFTT+KV8xzdUZ
ejmjte0Oq+4sJ9K/KVA96KVxowTuJsX5Bxfgr4fGSTddT1SDcQz7oZcd117UDtqqvxTuwEYqQCPW
ziVmMl4IGZb4usfcdTRhKzOeSEDKoGo6td05IgnR/wBRnR2x9u5lxv8FsCt6QhpYdD7csPpJ3Ju/
vlh7Lh6pUSBdNX/xVycWpKPZqUgvbqXVd3X3Vd79/c1D5r6yKUsEh/zHZiZt11bYkhJlDzWvo9vJ
B2CYpn0bZTDuMy5ubPqCWeyEW+fc5fG8/+JTpYbKx8XUX9PthDhFJCce6sHyucpPeD1QePdV5R7i
nSNwt0oPv2ke2c/S3mmsuuJE9FCGyfXJXn7YzAlT03sTANNtmHOD9z9JofNBFNYh7XZtg/UKx0V2
Po+rfGbt8ER8Rs81PRLDv++ksW1x0LlkZaCXgybFCjBgPLCt6Q14iMO4VNME0ca6royVSb9DNfI0
PptBDWqwe8a+uazaNJTchd9IVEy4MWeNUotPM6s+ZtU8HICuRjOaUtDE24UhfJJMAtUMh6alTK75
C61p0ELDhsOQDMder0Oz38Bqx4L5nNsPJB+b3KjsO+WliRlN/GC8reex1+wVHoYdIELXj1USwfah
9Kf7ZBybhvcdLZ7dlGK78+6jRdXHq9zyF1QuStjskR1quiYUtmjoSC1rUEX61XGZKn1Hw4wOrHGW
PPPKMF48Z8MX/5kOAzn47vg7FwegjJSg5bTM1LcsfqZfgjW6V0MV33iZryt3rtZ8trSC6RWCorDT
AHX5z0f2ymhrGuFrxYVy/9jKWhFjnJybFv7ltPxYCvCXM1ln9o1cN6iiF1YwY6Kc4TTAa1hzV8Jt
ukcIT/gef3MWblc+uPeYJTMiWrAElgNnwsaXAH6egKwBKgOHwE0GJO05UKGu6zrciUfwuJroGmjG
E96W+lkaP1uAnfYlyXDmudNzrmQ7RK1dQrRChKF7gHmZ/XtG4YyuMLaOeQ0ZzI4l5O817fXiB+2l
L/YeHJbk0BaDcy6vpDrtK35iScOvlp3PBFQt7wx6iPFDz8DMXJn+xBJ5+D0DSz8r7qNG0VrB7dfH
28fN9HJIcQSDsKU4svSd8/bZ65BdhIxnThejX1uIihq3kZYaD5zQlsQ1xmRmxPsM+J++F9Pgvq5P
GJNoPkA6MzMSeMQUu7dG2cgl01FQqVB5lvYYT07zqUI5O9nvCksl3B8BJz2lren7A86fpz/w8kOz
4sY84HnoRC3YBMk/KL3q4eWxsmiNf/AQfrz6kU7VA7Xl3VCi1J3L+BnSzxivAJ6/XNQ6coFj1uv2
j+4bug53avWUa9gw+0JwV1t8ElsomEGCXRhnfFMlJyRdejyRfk7Rlj2F6/4xvPLBgzqYr8QlJ4mF
mPy7UjJ2pIShX1sQDaCSQ7Bgu0cpcQHv31yJKGFr2j5SJtLUjNJSeONJp2vDzEf+YwqqbRjIhcFO
G1hXzDWDrndLtsaVf+GpmBDQaWZku5J4D2EoTOTQh671eXE9AGoWjlkq7GAfvysL+cdweWL3vQG4
dqjmuo7QSrc+JfFvkXmCcSEg/uoND5iYdiqEBdTmqmaXgvcV62s04GhHa98PuzQjL9h5D3ugtMEz
2Ky5ncYxxQkRz5vZtX6UZtfIRTZ5+23S7pp9vqw4UBsWkNLuZ7xRNtDMwkjVutxGeFpZfWoq7bnr
33WjRmY33Wnq+h23ZPmoeGZNgDYbuQ2qjQlWThuCkQ0Clt1b/Sa1BExUL3CPHor3xvBQf9gOwpae
aEn5lla10Tk+qXyjYurfpjsfHv4w2mtO6KrcALHTXkiwyRjlaTZeVQJB34OpN1QfCTUG2A8mS2kH
zsa5JegCpuhNo9IEtTq7l2vnZzgCaQ+H03fIZZsTdQUb5gUWbJgutY8hknLqh7TiR6SQsSP9T6gL
1fGoT4y676JCx+3KF5rceR9FJOLmK7B51qphYlfZ8sxYdGe+3DI3IejJz5k/4gSuuEfUqkETQdD8
f36FZZHIieTBJYeUM27/qYZXd8sGTphlk5hLoEK9sNLoJcYHr6vqyNhgYWYDa0vrCi5PHnAHBfeg
CsrmcMYPtizNpIn3gX9LsCQoQxoo3QD8akrVF5TXsUgLpBt0sqWyh6PpVvvcy6CERE+LXi+KLVYs
3nB7gHCpnJ85KQBHL5xjobL6SuyUhPmxEYQWxQqAZQxxkhx/C6xvsoyChS+FNwot9fpueNFbP9Ya
yksL282EUfqKjlU3OpFFEo87SdpVCF19hz+S1oBCDtJLY10PdQC35LVrK8u2b20ie7Ymh9/CAFl1
jczYinVN5YuQQ+z+u5cWn7+QPfGllg8wW/dEbpNbP5KKa52bFPNbR5S4XFhHdCxkq9aWomN4ofJS
Aa3EgU3SmzPZ+Vp9VALKy2h6mRAr1LsoOPpIWKmdhunVA2x9LOpvsbOcIhTXKr2ugmlTTJvoMEOP
+wDMUrbgR0TUyA301kEevskpJL7C+qcnUwlJPRO5wdhVgftlyBnIFMA5CnVVOFtN+FHEUAX6VTSQ
EGwk7KBt120VctlYioK8WtWPcF+SVoYXVpDqNaW+LWGqAW+d2s6AkBhstVKbRRri3S6OuJDjdL55
BRC+JviShXGF3IJDeCoSIdNTdm18AiHT+IHPAwI7FlsqXEFh5AfKM51v2cV/8lAkr5Kpr5vcSxhi
CmvTlHQ6PbFxf4K935Db5Z7BAM5bPzbyGswPdCIBykGUn5a6juPWFlqsLCYRQb0Kzop1dNre5+uR
rdgE4MU/ChBc/Tu4ZLndCLyE59AAq9I/1MgT1pdZnrVovJ7Z+gyOV//jxz/n0MErduTtN1lR3yEV
8Hkc7lHervPQAszeRNkPFeDYKpKp3jgNiKTVArjDeAZ1rpTG4WFFPqPH2hqMtnayvj/2nK4yP6f+
634I0Km44E9eyuCXUMmR8DC4zuBtxaaYbTJY9oxJd8WJvOs82t3D7qcXPKZ+9kA07DQU/QYSFnQV
ft/zT/BvLqRPaWseLRVuZWduL9os+/7vLJANNIOAWIFvVL0kNRf2sjhfkyLL3v776PLf7oj+os/G
T0A2wP0CwUC6kKvh4jTlN+yclzgg0OtO78d+lNHrzRv3Kxp7qY+XDrn/gD/RKgTWBGdq2W5+ThSa
Hr4r3QM7juej7snYLKkKjzMICbjqeiU99fBw+sIScokIfTaYIBtCvHqEb/uERuKNeOxXmZefuZuv
mCrnqzfHz9X8aJ7AiYfUgB2SMYNGOxbx5hkgr5oPp+hvRL6G3aRCUh22yU+EjRe7JVUq4yPbtulw
JnZVfpC6Ec70A08ysis7kStd4IDw5b8zkYmDwLftMYG9+vGePNlUxfHHJB77A/F7DZEm1yS73G8B
iTtynCD5WmZcfyQN9NNfOtmZmJrAmIoHad+J+OS8w42KHYg1ckGapYr9cmAwCjwIsNrbcFOv0ARm
TtrGJDvK4IeEWwTQrJviixAzZ9bDG0WrIbdc3e5zZ54ZpiCRVRU4Ant52bv8gYD0bs8uzlOrIqbX
/Rvg2xuyMsBZRF2s8YRpZcnXaF+4sw2zfZ3QSbwe43AjoPdQfRuU/+xSZ70QyxxN0zwRx9JSb81h
+NeSlighmmjNsLBBQV3Heh/MCSdD7hY8HyIUaQ/9vSDf4Ke19DIW8nJmrdIKZVeReDtJ479Xfy5a
+pGANtoTlqlCJIBoq60rnQN7QUP5ixCzE+739CQr0akaw9z0DU8i8JqdgZwqDy5Kb93lzZPmzrKG
SWg2y9Ejz0dzoxyX61gh3SS3aP4lwoz4JLqm1O0cml56IcHTHLKd9dm1aawhznT9J5nUxT1eLAXs
lcvTZs5lLCxN5d5K6V1778ZCGULMNvmoAcOeZb9TXcW1kDPQcn9MX7D8X8vGbFYbVVyxXkE0bkSg
iaE0PHmpXw/9mcbs8moBcv8ARVPqd3N0gQtuWaIj+chmsjiIwNllyYDWZkEZ1XqhQpi8TOZplHMe
YaeeeOd6S4E1ISzyGU+aeR6iRClutUAYp17e15eN3aaSer1uKN7xdykKe9BjANaopE/3yaAE9TQd
A/u/3TaRAl5mbF73RQyZAoVQ9UhmaUKJ6LAv/rvZS63FNhuLDjx1Uf+pvfq9THQLSUR7lLtjGTec
J1e3ptDgifLlcZZSmD6IXq85MyQr0PoPYxADmy63cXF5N1uhlqZiq7ntmtvJEpyE7PZ6MBKBK0Ot
ot8eoNyxngl2qpLvwyhTt705vhVigNjdEaMWo/ROr+beyf8kcZI4vPKCCAgMPzqr1Bv7Bb0AUSMP
V8LM2PBDogoTV9XjaKI5BjnF/WEsffw9mPw7ukgfgQhMDs1bUzBj14qAmLwAE/A+xePlVq9NwZir
9Vys0lwFkzkHbOczUC9XTiw267wbre6i64LLAWEJUGCNPeGDqfk9CEgebtPzQKi+Tk8F0UZpCcNL
X7Nm/OAmSvDXfbERjYAViuJBOYf4tiMdTwXYxlatNhCLtUztKBpDITjaeK88Kxh59yAh72OhvnX5
ABj2ybRJFZ7FcAeVqGhTGzaxw/47VmvDxbgUUf7hPg6PGe9mwYex7pFlPXK+PHy14OJcvKl5xsp2
Su6qbxBq+6wHsy0M8bubal4Nb6YLrkA+jW2XH/XLcoabrGRjfSgZE4MYYSomM9L94BmbDeJYG9rH
KBcJMkhMouHOlyoz49jjZUwPWgeBy6xukqj7kiqvVkOOSzQ7vqruvEHRBGXsSh0sxRxTgkr6CAFx
2vKrAQVQXFPigKQD9j3Igu4dLbEOCx8ptN88eydABMsgeNy++BYGZoTgFTsIdSv9sClpQR6/nrlL
VPtOG91r/6+x+1FWvAuG5CPJSOJRZC6ED0FNLmGzPJujEA0si1DaL7UmnhCFq8t2aKb4MKHAuynb
zsDHa9TWYH6fE8PvSidAS1xscdKCOZDZ/jchZ7sTItEczA3dfw+rFO5afWnbWVUqoLx9UOwTM3dY
5GPRhD6TyakUZjOGwXmuJ4VW/ErgWPtNqlouMd+fR459asnXJSaoTC5gmYSxaZW5wZa/cRf8m9C9
42/qsL+0/7aya1/9DvC1n49zLSk3TVb0UzCqhR308IU53/bVTXRXN0ugLk9elqdzwqXbKcG8uPVM
GkmAgyhXOX9483ouUwkojrdFzAuCjPPljOn//0YmWZUKBs3fDjpnFwhkVa2+yZHAwTJqQD7BUBpZ
oLwAA4wahIo80syhdMb7+LuTT2A7ZGsl7jf9ibLgWUY2UM1TBeQNFxqqweSrwlXR9LJqfjsNqX58
/hQreDDnJBRH5qr3TEwTAfMijntJojU8E1i3DITEiYDAEDPIl4dTOtF8GNhAdMG3I7vnp2izV4t6
fagQWG7q65c1KxxLHVButphhw6i/cPYopxPQJUheXguS5vO67PSu5jKHLbXBiQbuK1M9nrNEtcRZ
GifFjkCq5a/2WXP8y/U9xQTHJ8YbAxJO9cKa3Lv6ueCpIecKQtwFR1qdUIt9TAu7l98yydl29M1d
KXxL2Vl/cUsKVvQXMiHTsE9c/tStPZDXZR5sTL7LwGkz/5Q1oyQVAtzpQId6Fg1X/CvC5rDmLAly
Ymj2XUjif5L0LK72X+uoUNLNmlf+Fh59XyLwQAx3U0XE6pwIWyMFPY+KuxVbZt6AuDqRjkSTEG68
7l0BNIZDJecu8Zhw98Tbpy4qJY7j+m+em1ufIn07IxtrfvEjAMEhk8jRjvJBQLy0dXZ+SiyF+FUU
rWprBix571HON5VgDX3+XAFbjss21B1RJ4rYiKLA7QXuH/6YCwiQMUiF0exWxs8GUkvJmM6UkIop
8e+v4nVNdzrJBsgnLLD4FZEPWvjn/QoCJg5IOFYrr/0psTMaPH4bhnf/3yHq8+o01Y0s8ZbhNHR+
MGEXVg/pV7FigbebG/5SIIOh28kJIcZeTzd4f71FVefFjn7lzp1as4zAr6v/vbtxIi9YbHx2EvJ3
OGtlM2TGFBo6Dgb/LOwS2oh3ifY4IQHmvbe2Vyblwv0PaCyWGzqv5nvQWJw7Y3rwgZuzbYPxzwRR
iBrAoYOdPGR4jhO59iPidth3zyHQzFCUk/Edj8D4O2h+ONWNtPToWNUxEwFdTpg6fMMdBDiAp9yZ
hsmrQxV1LRLktQjyPHckeozzyW6EGhQfnw2bT3xigEmp+cnOwY8VqkRzZP4yRG7KNuT+8eTOqwHb
fFzyqtUxPZhHDSQkKJZSiUtZe86xxD40MBEZw8tylE9dS84obiLnLZAn/TBaARMhY2As47gpxrJl
+kt2idrUQp57p5lYvRxCx/XG03tX2J6a1LD7norZr7sopQBZINGl9ynQXGoYySg3fwtNwaz8DcU6
eJkCPVvc4GKMGzPIz5F9QQKc6XvYsI297//iJ4tIhg8HSlkMkca3VZaU6f1aJV5US38GBpG1ZOTx
GU8wNnicT9KGLra92uh5y3amDg+YKGlXmzWlYlZXwV5+ssitz6NzT0loGWxt4ei/YmCaq91Qh86L
Ka6FQc6zOwDnm8CmsxcEM1XjpGlG+Wt8nNtAvUeFdc7Gz4gqrY1/Fa8lovjhbDx8u/b0StUQO1A7
2hYFp5z6nSLKLm++ee6jbYXNe+982fEJhil5CeRSJwTtDvAvGTS7EE1YD0bnTPn2+E69e9Otr8UL
V3SX9OdtBwmPlB+uDpdgPWZJgTrqNpNdlJyX7PkrqYgNHjgE2UQc7qch8XIShf7CHIWiYf2N3PKc
+HoMOn8dooerk+kF5jBE5Kj67D95p5w7gSOQktEUSuQVydFtlTijvhLRctjat8UL6Y2b6k1hySWI
d88WGq1HElzMkX+W1dxC/DQmniV1aa3gMdQ548KRBDMJn8DmTsds0M6p7SwFF60rVNf6uNxTikAc
Fle7g2NJuGvAnh05PWAoGqUqXqsLvFyhaWENN+xyRXDdnak/EHJaE9I9FeMtTR9HXejzuGajOKIS
qUGTi+8XyMU4jgvBOGo04d/6yIPz91xpm14UnBzY4Ngrw2csuoDzr8+t/EkGfxKHi9+HpM0Yt1dl
mXFQDFNqgiVv9y+9k0yzJtljcUw5JQSy1SbJ0jo9SvDOzml7amhPFbw63BZWAfxSgrv5OZRGO1XN
ruPET/x7DWD6xPGexPoaIYj3LAvZxhMLPrX9ABNtn8ql/b+/RjMSw4J2sxnewR5jss10LT0+T5vu
1tmP8WDjuYtOAmPDxJrTbSZaWSlRcXLe5VxEY51nfez/o8E/Of8nsq7KQaTPXVpDPg1/3TNyTRQP
ixO9d9TKJ0/PKS76Y05EyYllStDuxOStK1skz0AgSmr5q/KEDOsK7bUYR+nO/zDRsqGs8wP7V+ms
a7OkwV0Ye4wpZD2rCXMpvHw2trFWqql1l2dPXLnHZutkpEnBs/RxTsUdvVtWiAADFQfx9bN6x35J
gCXknr9AIY0yGSzSfR6R/JzKVkvfQvu/2lhonxZdA5kNk98t25Qr51ZJsGSGCxEAprRuLMEshodK
kBCtegWF02f/pMoCBftPhsJvZkUSXkPmV3qkgS5XNMb75e827QwDq8w4ilQPkxUcK9eCVGSmSHCC
sy/1SKbdu5TYFUNjKJ5y4X+TklwMAyQH/dGxLNk9/i7grBnHcYhj/VCjOTdj5uJRpjnLfMvcBiTd
BrytTJjA77EBbz4GYwt0ISmMWjaHQaDZsYeFj+IX4oMkerlAS2ZsHwCMrv7zC4iXq7TtLCfGSNL2
RRr9jIsUiF1u16mQRqx6G/UIclge7VsPphvV+a55HwpnxVvJdif9nkG6UuZzgMBS3oReXzcqoGRJ
NTxMovH0ZHqjfNRdV+sKo8xwfDAfiWF3RIha7pOLE9qKbAShFYrLjj9v2LIDl/eO/nJWgcLUQm5l
Y15a5QZu60Q5kvSC4KSiIVNqaLJ4BifkdPdONi6TMEgSFUPIgC86UvMzvqAZxa0XiXXfpj+SXibu
Abwa3sC94ppa2ntsiCDjqmq3dk5d+DaJDmzGkF09CCOTcotZJDxZdJ2tmJQuZ6msjFgu45Mc/+Ya
HoVB/ah98l5eBzpLmCraA5dgLrfqRlQefEykjyydIDfBN3Z//2/3lSKU9FU1h6nKL+y6xnzuW/IF
GxQdzccmiZ0bKCJQlGCUKX00OSDM+VfpcsdFC5X0svvUZWuWFu+ehvF1M9EgzMp+vG/7stK5ctXk
SY6coZEQFNuSFOczC8Mxj1VRLVkx6qyj/ti5EMTOtZMUsfMgPB55i52DkgHmarbSsO7UtikSG38e
Obp3eA/fpp+hniGz/bYGANGj/3A8JuaLz7KRjZVRtLXjsKsQtJFx9vmG1nLtrbFPR/K4/6jNoQuw
80kvug+HVkVYiMwH0qNIXeUsY2mL2B2a5uZo3jRgz5EUwm7T4+YD+67gljr+T5SqX/0Y7a8OfHCN
K26QvWANFjVGC+btfYNn7rBQ4d2RzLHNnHxc2VOxLnMO4Z5qPDun2mdKc3FH4Qq4Iv3t9jIgrpIZ
KldN9zUpQv1eq8oWxfNlGeXrNNySAKoC5sW+arhN51afH/UOTVoPbGrjlxD/3akB9am7QdAPat97
w0/FbWjdrvE0mnnHScgmzp8XCb8EtI6Hm8NYHmctmYdI7ysjX1DpMxFEXQrbse3D7ggB13+GXXqW
g1sbJrEPcD1SsjMf3gFS/a7V+GgmhYvjh9woVdTa2K6vSf7k8cT9/z0HmCrysMPYnwLq7ukmbbZi
Go3zBvU4pMPpm+uaLs9Q9EbAVJ8o9zAy27Qb0P/teoZF/Qj0HSuUMvtLn0iVqR1aJc1JS+v8VXax
6EHXDE0hXwCTp3Jji9GzrwvXnaF8VgONwIhTdfoQZlUFR86ZNYCndb9G1xNSn42Q4TifzGyS9zVm
0q7wnRwO8b2Z8yGF/LNm3CD+Eu9eitonNT3Ng3E7CoA3ETx6DY4cnZKDhJgfwG/z34U4x1IP8d2W
BaU5OR4GhKEFraBCQo+cK8lL06dmjxmEqTlAZ4e5XuFY5/E6oINrjDIo8ysyKw98slb1qwKOBQoG
FyxUipSwlnZQlQsepPrlmhBhphLqn6TGqi9JiIyaOyWvoemNtp2Qsc1ANXywzcpVre8QvK+00Pli
ewAh8EaHyEico7aiw+lQVmWvZiJCJSzq9P+0Xxq+uOcqpKiOn++PCS8/yFULpPrGjQQ7uEtb3hbS
fDvghFpSmRLVPMXB0iBVDj84vif5j1UZwrIWnYpzxMDUOsYwyF6OtlHWlStdoP+4PLZNeH8jKO75
ycg7Y4QWwAtqamb15y55UV74uqtYXkgajfXEy69L5lxiaOr1m8VU1P6Rvvu4CrisYkUKHPE5/EJL
J0BE8zP+T9/01rqFGR6zIhu7waLo4Mj519NKe3mwLYs53dYQT8BDY8qntXbP9Rjnf4WGEPCO/Jzm
gPfx7c9qaulT86UQZz+25a8T5MNZTiIRERa8oK5WVtmPqjH4THbjDKN6uwJmyu98OzFbi9263zRR
BB3AtXLe9es/kvExeZcXg6Q1EsR8EqsNpzpIuyZURnErkzK1QF/An+SM7p7gUkDpv495j03V7mdi
mOg6tyM38xWu8JFc0h0i+Qtmk/2FfUQOCpJ8Kf6yGj7qhFY+fTBGNvlJfZwmXT76hkTbG3mWCVJu
L3bz+zQSQBK7/lJDJ5LjERtQOJ6dzbRJPu5VX1blhyVbYBi6Q1Mam+VoL+RglLwuPLsR8i7L+YjG
DzF7Xlb9JZxV+OOBYzt0EdAFPidROqVPeZeVFoV2yl3mNUtu4nNHC8rWCngMkwMVvPnjxI9pu5D1
qj1VZK5FSJhdKOlskIZu5t+GpMWqR0cMC2Jra1UIaBBakdBUlNPI/3eC0pvxEy/yHOWYJyRqEEcw
WsCC5D7iHnnslHHyVtUgIGCC33fnlY0gNWklCcQCErJ2yYIkwDKpWwwNJeYMF0qDJ0wf9W/EaLwj
SEcpd+dTr42JshiVKAD67s+KCdjimH6lRY1VG3l8BnLFNnbX/0wAKmhIXQF9PEVNv5eYNqVY3Jlr
srOMekKmfCA3vt4DurVYrKdRRU+uB996/9MYjI/ldd/5S6WdayD0t+ZZrJXQeFU0TcPLhad/xcCB
8FWOArmozsP3MVAuMpSCzYy9DMr5MZYvs916zOKoWRKpbuiDuqy54P8cFwTk0MDCO7EK2dmpNJS+
d+xASKE3r8O0wtpwKkFPQNBlyoJENroVWNMW/hFGtbsGzZlB0YzZsxxWR41QZFkFzCW9zCIYqgSd
2qM04hjZ0Bo9MkXOcFku6Pi3/ZY+NJPkiRf4vH+ADOJYNUMZmmd605SO2UcU//IoikABxTEDJyTb
nvMm37MyaafCvU/w2G7obBDDWoFfji8fRp9ZgKozmcphE8Aq67hQ1KaR2UQkdxvePh6LTPHDbtdq
7ZMPVki+tACm1k1N2bqwQCJrLovkjMWmPawSJgER5O9Kf7PHe3umzJQ10lx985YZF5HqW11c7t7y
0vn76RvRojkv1mU3g0abLn/XWiFEJ4HnMu2Rs6Dbdrh/zdv1FAB/ArlMh92cAHWx199eJpjW44C1
hwIv4rSMrnJ0KuAx1YcZnKR97jRddRnr5baqAyilQzt2DczR7f+d9cFkVi33cT+9LUSZvFGsEKZJ
18eaq697xzzSUY3hOY9MD7UwK4XM0j5+lGnYefdG3s5FtpNrNtgfWVUPTr5jlfpMjgLem91JpaAF
7HZnE6SvEbYMiSB0MtKHE2cJfzX3Ga6DJ34I/w0sQFopTPWjjM7r6yzU2zaMZoTBqPac8D/lTPf7
HIIa1YlgEXG2CdR/ukyUTiIMpA7hPExoVHNJNDnSa2tfoe3PEr3kY/vfWSG35hQ6tZFhWjg6qhVb
Q4y9A/CWaUx9BYD1UhApVN/Ud14dJ7j7+txjb7ZJfVMG4lPLK37uHNzho2zFFUKS+FAxRLUks9vP
sIwZiBzEiNn7xnlRGcL6hYrf+X5aAYkOq6xxOIXMHGseKZ1XPBsQoxlN1/CnsPrKMmw57pNko1cj
O2hhvOcM6+ngVu0CH/bYBW3pbF968kfvVuTXniznl5mazw1Lx5cyUf+qRdy3ySZdlrO6+uet0kar
89js+tvEyqbnEF3a5dscKWk+swOs5LztDXcTQAvzj3EmtMXhkmERWNTW8U9E9h/2atpDFtp5LWUS
txER//JPYeFgkeXUskVn0xMLiUM0le/iDrJcyBQfFZ6AzxMdp4Jh77bWwAw28xB7D8+Ghf3DIHFD
1gIRb4gghEhGPpWaJ5GYRpM50brAwWUSxeVHs+SsojhHaW66+laRoq+ereiNgDRyXlrRYo2GB5JY
b8+lUEM5Ub4fJ6tjQ7Y57g3V+pbZzCJ7TksXmMOtUfchj/aZWMg1gjtFTDM/HSVnDoA5B4FLgQ88
EfKc8Vil3ngISwDv9W0UnKbPgBSO6Y4ezIJaEIHVzcSdB++JToIqklLou4yxQnc6kN2vCo+EKVI7
nIGKZxjJ6z8Q0g7cf7qedyP6oAUNz/NI9Qs/TPhAZdqKe2qHTHKJUQcT8uJ2StgqJD+NN6z4ac3F
VMdPHmSppziCCJrIz+Kwur97/b1ugG+SPU4bn5GhGYqzVqBu6Pcvb8cCFCYrJus7om/xLo0lfbYP
XIPHD+afNps8Iy7Fe+SX+Up9XsgjvZFqlyvSOx4VifK5otozs8aFL0w9a8JTA5KvVq5HJgH6kjiJ
2UwKyeXst+NIWo+XFpGg02xboxfZNRVadK1Vb8Z1eUdWEZcL35iAaJI5+2kv61tkPlp46+y05ed8
8/qKcDjL4CfpLd9ljvBNw+lni/fJcZ4MtNHEHHB68KrBpzaSMwxFVi8W0wuZxRciD1KvgyXAEYEc
j1Vgo95/2Pva4wsjoSq9vc5c7rYrBkJp8O33Y/QwuTPFdTKdxwuIS1mAn3DJbng/t99Tu5cqAdC5
zUNUmZpI0NT8/gMtz1XFdf2K++k8DBQZsJXB04PmLQSf3YQvMx1GBZbh0bv4t8REgVDCQ58IeX1m
hND+mJ5l5cCFfkyz7WG/6Es7kbowkp/k/tY7rpcfZdfUKakv8N5Hohh6GwE5gN3GX22Mgvv+fDgI
ICH+40QtV/TqvQPvzNVdqtx7vAGlDCspodNn/fBnBvUCXmME8j8WQ5451I+W+VLOZ0BNJXhM6tQD
+K43am4xXiUscVmBisCIxCr+0XU2MwxSBbahigiar0j4VLDY5ULFwDVVlZJE03zPKmhVTQi6iRla
hIeYeh37fS/32kjT5DQATAO44YEpxB2c7V+B6PSpDdpgCXh4E2PlrHuHwcKq3kijRSifvk0zo9lc
d5S23Q++B08D32gEYtLA4A+C2K8IPgLzbIa2a0w3EGHsPP6OznCtFTyntB3/NOz72D3o82uXGTeb
nmrAq9onBtMkjvwRI/M3VgsiATEQs/m0dqAfNfZXIjm/Q1NqB91kHTE2iKVmFi8jjzNcGtUTXaQN
weAscEXW0zexH1O/g/yMnOGHreEmzTRBPpmqwNiPhLTVahgu/j4wEoWB61B07ynlCyS/CHAkUDi+
YQupkfucand+yf8317VRnPVTs2v2vHmpzymfYWXNCqRqOVJGcMvB8hmgZMq+cwOZBkqRVoKxkCoo
XrWTXoEZj52gKMI9gb2EYQWLktL0pv8EYmDieMn1toqEmirpAzOXEZrxiJgCJM64QPEHojMrPEki
ot7Vksmp4TcyiJcRGKiBG0zbd7BOkuL5EvkJeinOmICoMddPNuNON0mBFboSJAjeUXOPjmgqczgw
xj3QIPlVDV5pWhHHIOpY0Rj0BP+qK/lP2ZpPaDynwT07PDZM4vObs9DFBwKZdvNlE8oBkq6KR8jP
EwuF1GcUxHoX/y0DHKikWCFr3SToZaODXboZqy2VD5uKK9kMFb7zX3HFEOrYjhANZptbY5YUTUcO
M+63fkusBLUQYJ3KKzolbfd0siYtnmz3cOX83KH6PRYUw2yhNjZIHo5H6fqPTNLeQ+m83WZVOfKG
TpHSRTRWtR6GXcEC3f1Llyhn+tz2VATRnXCEdAmoANROb+HIj4Q5gojNDzgbU2bvfWHeGRp4NQDq
v4+7ofGhV5O2tvEQFTQf1x8wvGgakYzKVL+x2emnJqmV/IFLlTGrJUzhlmbnrFWn+knwf2VR8JC6
li9ANadZwkbAYaRgYVJ0isG/foLJ1ZfdpJy+qdu4AAlS1KUV3OXhr9xqFKhb5/e+01KG04D77eGx
+OLmiJpKihL4wGSnqkGrNhGHzMrdGg+WRFjH/UWFBJfDEgJsCIfCdPfEtx94TGqPiUrmngITYlBc
Dm5MI3KKDZPjLC8Mqld5qGa4Ek9sBKxPi8bVziiC2QRTPDIiFZeWfgw0K5irgsaMCBDx6KkHuynD
EdMKlWxW52rsVpLRW1vJL60SGgfN+9McXIukI31I2p32ktmAGz+JAjivPCIfXk/9rfqcprlsLpqC
z3BOHFbcqYBPQ4fy8KkORKUnknm3QWwlfMhWb515R65l+T0C8ioc8sRyvWYYBP4FEpVspHz19TBM
f4UDQrALwtf9FHXkeMfqFFhYPBzR/eKzECDzbgycYy4eeIEk31EYMi9RW84REvk2zRkc+w9jcjEz
+T21p5TXndHthl9avtL54On0nIkp1vTcp8nX7LWcfS0rawwnabdLpFhpA2CVuULkHT3+LuWAqKiA
2mUADJgtKshK+eH6mH9UgZqy1GqYUGaI6YD2jUD0eZENvsPDafj4G1kK+ncG7k+3CAqplf3WW8TD
3rIQe4PCtm8auEdIaGpB0qc6FiMl8on6H9bFNf26SKtiNhksfNDBAmMfYnJHVftRyXp8+ltgRLip
k+PftDNejjx40+/qCO5v1bcU8Psd+bLFabtSli9G3G258VIJFWIAEtX3t0U74AI2PP04vJIzG57G
oL7ZX/x4ArOMlDFjQY1qMh7CPEA9y7dBsY6zKAWb+PGRohY+qfv6fR+1mqYWY/7/y1+7awcRWYev
DRgqHqdJw9SpD0NrYKPOU5YbhMr1Ilp8fJqJrVV+kjLvaQh5qLMe+zqncbWfFSVe2s2bOyBiUgpD
Cod6spCenVsF6LONKd6qU6yxKiQ6LoABix5rE0UfETWcfnuBDPjswrxVakmQa3+ozOw1DQrRLwwt
343MUDl5RMXyUfLrpiVF1DGwK0liSQ2vqR4CSu4aHlDEaaCf/8wj/jogEwYMuG4zMVdGo9DGcUQw
srvcTD4/re1EjQ3LpLuL7Hk/Vt/U9f/CfuviwufN9QcRxx4H7TujmSildrSf2GHBXcokuHk7kTiW
PWTPAYLHmguOhOdh+4oQjueb4qumCHg8VDPwbFvimTn19vf9ZQFtV4U/YlayMS0eQSIVB4JrA8Pl
m+agfKoxvGBJqhVaI5xKtfE9rAe7HEy4Nro/wyfiayqq+iD26XLmSanWUbyXSiF5huSl1P5fNhfd
mtEvgZe19DQTHWdlLJm7QJXqTQ3bgPvvYBEW0u/Ug2qD3nAo5soii3GQnwcSR1zJsLivwsiq1i/m
neZLnhOPs6IVWmnXc3ToytePXjPqELwOzaiyQDDDJ9/iFL9uduwrmntM4dSR0Gfh88wD5lZmB2DI
vgcTtgHA/CqYjvm1WAOaQtM2Y8gptQBlLWFhyaRlOYGQ132gjNR2Kdj6vKXFN73L2m2D5JF37KZL
qoAGdFNnLmBVGoi9ql3Azhuv2Car2p71A6HbxMuufYPCNvyC+meM9ipzNH8Oz+F6iH1i8aYCsGUm
Zjkd8bw0DaRLv/0Fvqe80tVvJfuH1Ny+uRyXF3R/SeaD+L06dWd3OKPVd3jCkH4l3d/1Kguqf4sb
nOKtzUwI6vTlBalqINJrA2SBgQcAd/9osO3jlR+JGEtozGK1pNXQdGTgfUchzWfx09Q40gpFdxas
UdCo3Us2/aNgWRKvvqgNKUNcOOna37phjWo1saFfxFc85A3OzRRiC0WRBaYXKaskFRBSoq5BZY4n
uPdaWiaDaTX7KhMlHEcIl0s7h1PmPgh+hwKe/LtN0DDdHZByAjQITPXuifnE51cvVul3HLvaeStC
D8pVrcPQS6a18gs5PiE/JNzPFRvVgD+dtFq5JpKiaLBgD3F6n51vvmmkvB/q3kebCXflNHzVuKzl
jFF9mQRLd8W0atI43V4zb0KzJZYNxP3S7Cf8uwVq4fNQ5kzOcJ9Uw6d43CrkJNnOnXR+iBaN9nIr
iwoOVBpwiizRI2mbSj9HMVY9VXwIMlI58ZwYPsPIY7dhHqAa7Jk7ft0+P76/uIJsZ+HetC1+0eih
8s2+GyEUOcMW9G2ZLE4B5R9dYkcUAsBy8U3Y3qJGbGQX5F9LeO2iK74vbf1fTa3XvHSHKacxHQPW
jdxKmicB1M5xVNVMQdsx2jZOXQvYuRoU1tMtMvCbNRx5LMqZN+qQTl7PZYXqEr2+M7bja+Y/mZ1D
NLCINN31sEzfW0if+70UKBNFdtni6JIn2ZZEZmOcyvY1YlSsp2UmnShA9bYBFdobAajmNID31mni
0RjgjC11BuKzTD0fIPGvix3HdFLQHa8KZrAN5BKIPzNHwLbNK3C1ITVkt9JaCBLl1IMA3YzQInDE
xhfnaUwpemzF2T6pKDYW/4Yx9cTpNpnCMyC6zZGOf5L6AgvYjInwFIed4pLyRd6QHtXefQRWFH0m
nivqV/DDz2lRtZZC+FNuj7/Z9MAeQf+yxcqR/IyuRPQYPL8DrymmIROogcj/cl+Q3UiQLIiGpI3m
lsO/yEu/AlBHYD1uAmwO0Ha3OyYFJt9p2AnrJhzbv85mHllrprlsOH0zfQKhSm+7tbyosmmViyTd
jsVtMRwMrA7HgkYRcsPARXzvzibAQ7yUI/I88Wlci4BLWSTjUVcUoHNZpvnI7xPjz9V6sDP2Q/J4
6Sbah4bScRuR5bqLTahJh8NEJaIf0xw7Mr22M6d2lyTq2Hqy3nFhC4Tq1yYf4O6dtFbyqyc4hn9Y
oBEF3qeIUbEBWfYpu+PpSF44L2/p1HJk+kqDckOcwJCz+cDcoJBYq5XZy2Hcpj92KqM1FX9sFb4p
FhV0UVD+3KVjzTJb7WII0uWtpfi/SJyodIlqS4A44IQcHErybU358wCdS35UpO548WbBEJk9BU44
kYxVmCh4i5rQxA+v1MZBp4MWe3wf9j1fk6G1EFPI1YM3sMll/Z4TFcxM5XWtfb0u6fPiUfSvfFz+
O1YnkInijofCafQTgM25Z5KUCNlcfPmInCeEqTqUuI2Du24kgBnPfEFYOuIOktiSFHAvkrAAYSqG
DJ/j1j933TW7jR2grn/+2G8fUF/DuZcCIUB9S/HRuGfZDDluJfKZjaGqosDwKPFNsyvhPGn+R/v6
GPvr3nmyagD/PsB1u0pV1MqDjxTcuKcCm9FM+agrMhdXBFEVSr/CFTppDh8oEtAs/bM6KyosHaAB
Yz+1rLni2x3R40Hle3zCN+QkioD7Ym66S7V3udOaQcvw7YOz644BZnAW9suYX1MD9uPndJJbDoy3
j90R3d+8LbNaLCtKGvjmXQJXmC5x7aHiplRnqwdakkezh310ftvWEHhL2lKr5S9pjti7S4ZO7Fyp
DmRuA/7cFYg1QAORn+NKDl7MYZoPO/l7T+VUxrM6fdAbOubTHxA+cjUfmluvrKz8fmJI3u+ypsrN
NxEMbhTp3geAqJZgfIzVDq0GyQHsU8mMH8Un6kCG6aNgBUFai47DhBU7vR1rFMBSkirHmefR5S6f
FXKANc2lMZidnhkSAjFArsnFNTfHOkzO6+wqnFT1k/E1MxgguDCPgmzY+neqLyP94uSG71rxV2U/
v/jYG0MYxtTfpJWnIVsS+P4I86QLTMAE1gr/2ARWaFqkc0xkEyX9qv11hIEZ5sed1fSpcg72kgeT
gF6FfTT85ezy/UJE32eyW4ECJVXfpTNR0G1yZnDs3Mb2oWVvA0j1Py+wEscJfsop0Wl9GG9liPPm
9cAu7UDxP/nW4R9KmgsrrWUhRNxRoxx9RMps9tFxtEErOu3ISEfeb9sfaqSHRzu+M8VzMEP1SF+9
XeGTjBWjgC28T3TYe73uobcYEKFifN82R9T/yR9lEp31mjWbANakyPkRbn52aOtgiQw4s5BhaRxN
nrlxGBPV1kzkgELN8jHeUNAG1pRoT0OVAQbKkHHYaObXVWfai3jvEJ4Br1FR1SfT4gQ365THzc1g
lbUuq5TRrWYmOjaCk6za5zuhLGOhuQrH6Y2Q66OkqlRLRVyfNOOtRhTX34SiqaUtlZd8OUcZUYBl
HDxyx22vn7gOZrVQT48XV+icWI0/kf1vJKcz2OMfvwubuVB0kPIqPxNfhhtAuUIDDKRoVwbG02yE
tAwRjvXfncsv9ZfPDgcokQ9Ll6GzPOsPFfxicZreoVFxqYqF2nWjZlZwwnBUFeM3nPHX8P0hSsnZ
kGRfZv43CXkqyZBI7zoLflZYksLI7P12nuq6Uaj3QCHCFUr/6nZi2RIZ2Eh8wuVLP3x/SiSrEG9e
Pwfn9hXNYQrwwmiiB28BAsK1e71LQGWD0+nM2j+/2bjDxdWwuTUIZtxQTP5hawFoejBCpmmfVoyT
ThlbIKNQRaufZfSOV+ZqaLB1HKYldAZ0nReSqfdO6HhztfheofymbGlR9nnKvNlf1dVHn9EwtsDR
K9iQt/HHOmi2QaSGKlqrXYFp/Q3o06pOsGoT+Ml7+q2s9IAIQRSWG3m8ED3zj0cJ9s6LSs2oFIrX
tnHMeHt7ysza27Ft+jHxvNgtddCNMg25I5z+Ib13OVuJinXsh0qwq3Hae2SjXSvSfL/ohZ+fXUdg
21H4xtQomjm4u+LGMlSVh11/S5NmvgI3NcgGRcWNMIullzOKd+6BGefPjSv+o55xjeT4Aa+hcM+z
vL7YL1mBSRvfmkuRpPc9by0g5fduQH7ClUYCgMw/pRVCFxdmmNGW8p9vEs7df9yDdLbbERMwbxOq
bq8ZbCOMmJSlT81aXlF39SwwKM5nF6icgzpZsAh2MQkVg9C7DaeOil99lrW7iSEYIw7ATJSVpVoT
+72ddhMysucJtcKYaz7fUlJMHe/RN9EMfd/Z2gDgi4LVzgyHN37FbebgABMg+a/aSqJSQoj+yoDz
df17502lM3FQ74ToA5gyggbilhXHGFH6U5UaCQggaTiQy7G0ATuvpM9fCSsfzmU8xS8WcQsw+8pv
WIOpq+KGOl8XflWXVQqvN+WGA5mpjvGJMlOy1zNA1olqBzTeuiEu/10BtMmHXi+ZvTuOvweR2Riq
Kh0UjOZ7ueS2zgakLChE9aBlmL9O9fA/xiQNOSeWwBRwv10A2e0pTMw3h21lDusBp1eu78j5Ic3g
7ID1VIAZhICK6FykEPzcFgoeaPBVq0KI94awohHbdI1W/5n+DuJjogsHJtROLa4YsA3ZEDbBJaMC
lazgn+YCKwFkrMYmaqa6bDZBtxuAPGs4gElF2OPQGTT7Q4LI+oR0QOy+mkbAg/PdneQTZhk+qqVU
pQLBC1swXrFue0S8JMfnUqt90rFWwjEJLAR1ojaxBynSf3BlHv8sqTu567gc/IMLyp+KkbUfa7Km
wvHLVG3QDMz/2zspXElJgfUaET+x8NWgvOiN6N+VlpLu6Oh4yK0eBeKTQ6uo+Lr2KQSTELzGmuQH
AxBEB9nm/iwy9WCxwTGgf1CiF83DG5IVBZq6aQ1aIrnhoISQ5Z0GcQvf0oXu8YYAERkJMvHSBx8o
zqwBTrAkEBFn0C0pLEeph0qtksBoJ1deoKqYjLGdtxumD7i1xSixI8Fm2fHRa7/SiJDDLp0w5Vln
nem2JVjFLeDKlp+ZtyIvMMig1wK1/Faa/wc7qeyKvkF/crj+WGPAHXaVHXAfqedsrFD1rwgfuVLr
dZRyJUCZROoXbdhkwmsbZ3qoHkMKzcqjuJs3ykb40ySEZQRjGBt1pvFhMVzZy+jsCONFmtdfM+SD
LDQNTlcOQKFr+fH1aoCU3I1UPnJJkWB5kmd1bsa6iB8HfVB0cnqAaLROWYqMutmdm6gLmlnbHDYY
89b3q5NXHX+VqMM0/vyfYhx7S0V1Zm8z8LwusQhC/UHC8zYs7sL8rmva3Y13akGyOXjKGJlwEU+A
fHeNHs7mXWAs+yDaA3ZbBA4DEoeL/dUkINaU3QWsqO2Ln889GjAY+f9XIstr+aJ1KweDRPbhu30N
zDh8zXg38QNxfbwu0cKGRLjCPBR12AioKFFVzstBJQsfJqv1VWIg1S45oNrS7ClgerKf/DU/CyMB
UWwduXryrQCvajhOVyJm2MXsw+MhYFclPd1yumbufHe/ykIyfp2RCcVTWqEVsbHt9nNQq4vWrcyI
drnHecw5BpJtLlLLX4pBfinbHb659qVjjePxgP299cUwCbFoAiNCs+CAHWy3ntW51HqEAY87nAbG
TO3dS16+N5Y0ZsGjL9yRO7lv3g4XXdKsrhrdpk0dPF8epO4Ujy0ZFlU0AQQbsy1plYD4kdIF7GzL
9ryAgL5LXh3xUIL8whX6sRX/M3ay8fv/gieqcKGOBQmQjN5oU0ZRbhn8O13jZo1J3vOBrExr52iz
XYstgz6UhWA5ReB9UfNaqnq7GVGh57JMNerUDdqj/Bi2TQXsPUiatVYcD5FN8pkE1fNTeB89ERfA
q5tHlIMFhTf6Fws6gHsi6RHVEvtOl2gxg2iqNGwES8yubt2LX68XQZVA/qRqA1xZ6Ev0Oj7m6Whf
gONfLoDncwTAU4txvTgJI14kVwbaV4KvTqN6bV75sQjDfMs2cXOLpHx06/5XMltOh4txkHf10i5i
9uS+GdVXS6HOBEO7fS7f+un/i7arOw9VpddcFUILkLDwjJLAIFUX7SMoDKTi4LOZCQDjI7HXWshO
kUxBOvK+I0Bvy1T9Oc0HNgGQvCjIIchenl54UJYAN7b0mJDzcW4BsId7NM8z0nHFnqjIv3NCHCYk
mhI5PCL0Is/MbBrqxav2+J9rgQ8ZrMZc8LgSi4+bGcwdghZvObulPDIyi+/uLOW+vXBestPkn+oo
PLgxid6MHi9dU+ZK5SB9wh3zHLlXg0vmBmMGWNPs9j8NYfTvWLtCFHRGfsgcm3ButZw7wt5s2Ja/
oE6ItdctizVUFGLhVafGQKLoOd2KRIo62ltKEUGNZm/yJjnM/BKqY0MlBLQQakosgN1bcDBaiBS7
aXjtGzzDW+XCTEgHOpBMVCx6SCXidsi5xYZTijZ78QZsKWoRn+FjD1hJLVl9x3yN13n9WJG4MCoW
9q+W/R4a7jBdREOXdR8Y4u/vSPnjovZiY1G1E/MIr+UEmxvmligMhMVuT2HCN20wxGhOIBD/bqpz
TZ0K5UxsOraMu/Wt8KqHxQPxUj/mrOU8nvUpzOowq6nuJttlhi4rJbo20FSAVSFzF5SPh6N8LrvI
gH5E7PCsYjcGLAS76JvRKvJFfEM6a6ncckm4N/hbhnE3RVGRbl5PKIhZlpexpEojRWez1fOB9ZHk
Z+uPxW7Y8/EBUF0/wnndzr35QA/B8SKjdRudCWcbcxkNb46MnI56vCONkHNLqz5v8Y3Fk/y+Aksy
JABAbEgdGePdZZaxTU7bB9LyeiKUOOU01qeuqDKibDGL8q3Wbuu0L/z0jZdGLAUdTnCjoRAmkcAG
vWVd8LeLi6K9PiJBcni94Qc0Inb1J8znJoi4q9QJ2xoDvDNRYk5X6VYxs1xUJQDZLNqClCrz42IH
sToTaDlcQYOW9WY0GfDO/YhnIHhspPEKgO20e00kaET5Zl8Ij03gs+1B4o9NPipLakQcnBontlWZ
j8L/mHm+Vd60x5kbmssSn+9qQZl/0gaEwHUbsRM4Eo0TDlkswb4KPd1u6YYox02aYgMARkPf13LT
NjSmdAlcJY4thQKI+Fpo7GmQ8145Kz/KW9TTVaH7L/6R/wxL91QX/j08pBeSh/lHKoKz4LReIesU
Ih2N+bUwwJRG8rJDl8BTQoxFk/OFhXHb6RcRsR6sRvDanRE70pp2UoInu7ZjDNVrd1CsECo77djY
LHgUsS0IgU7NQ3du03LnZK8JQiTf6syrxfRLftiSu1Cy/IkhjcBbKo4y+EXeWxSJVa6QjCtPYLfL
nW5LRWFxuMQLFuQyyXmTKhhb0T4IUOg9Kt6z8NkTVjip5mI8PVtA+Qk9TwnkHK7EmHNLrlX0wyor
YtvFQPykZVp3VMOEiK1/tAAPeoLSKbQTR5gN9DY3H/xjT+ZBPyWc99NIkQoH0xVnOscj0Kv922+0
NXetoZV/GXaMIMk2JyydooZiI/f2VeUddDWxRTEUU3w4N431wBI7HSehrf7S4fn+kWtoy+maLRsL
M9vnZjM1u4kgEOtmZRDwnEHPyEErBHttPotkiDNxQzp+LirHeyM2iKp8Cp9aDX45VwwOFjIrgONB
UMWwdWhGedbjjBz64gTux+dbCD96lT4nQrDpXuzVeQQ33i8SZAWelmt5EAWObeHMBsy/P9m6rEBi
5T6BdQk81maPZBYYF8+geN1LlEJZ5lIO3Y+w2AOY3+DUA+V59ZdOSqHYbN700ms95MHIYDv0EyYo
fjWWIEX20x420JIVDz0Y7cZvDxPR54RmbM8PcJ17y9Cz1nL7FUdlVxj96vn7UotNVnpa08xzWJYN
cQt1O3ZaJPdko/l9GHBrwuw3VFyhr1RmtBndHFcA8/sQMjIIsLkq19P0ZaFyYN3jCmv8+WWuSLlo
AllCVIDxVucT84IV7xCb0WdjrkwddI5JPkEYLD2EWXteZEzeH3jOG5bxGG7Ltz5UtqsrOMSUj7Yj
AeWNrjxBmmdyi92sCl16m5UYVlsGwnVpGiisZYUbowPgcL55TXzuaTn8LndhPitLhqHzbnhC2f4A
WrJMgUuO2fg1LYxEmJh+9L0h6tN1GQA+qdgrPrL9OnDadvhE8nh0Kin7uT84QvWqIN5W/f0jojJr
OfzfNDj+rwogesGguVQ1rFMT/xpGtiFObR87eub3wLlHwS1/ie05hTgbRgROVFv3p8uNVBQKKOkq
s+Lu+FU0AQ9xrQpErjJ6x1RjroIgPZXNsrK9Cl4mQCkBBXzdmnostpfooyp2Of8cz53HhesmDQHC
Evpg96SUCcF88Az/Us2iKw+BVCrbtiOGUVGE4N5MN/pkYZf2pVyew0Sju2bdOCnwGcs6JHlcL1rB
42+87al5XTwtljckI+rgCrCfTLr0IfnkxN+Kc1nt/WdG9G02B+vjD/m4tiY0wa8uEMxwoJ7YpNYL
Nu1kKOWBVb3mzBsZuwbfbRyjTKfQQKnOLsMuBZhaugO97ccFsMtzb8+WbQK+Clcf2HgKStB4k7bl
X2jECAfbpSowbY8T18REY2bwb6Jubd5HuYaxVUGhFtEhDhC2Scp9uAEz9REJV3PUZBAY5GFhALH+
5sw3tdP51vICtZTYibkVoHlni0SKOxBQ1IMn6glg7bjSaFYSzfZFSq6iMfep0BohbZlnmQtWHwxY
Lct4a2vSiNdjg5vXRw9AbTWDPp1/PGjz7lkeLcOvxL81cT2Sh06ikfl4I3YUZHKS5+AlXW4Pn/B/
Wz7zCvXjeKKTSZ2zvj2AsT/raH6Y8SAuKBNJXSOgxoA9KfsP8oLxOjuEBUxkyoRAXzAcjJF1gP4A
j/6NU/M+UscqQ7zpgYkCrhcbrtt0Tu/enCDA1XOF9UwyUc3mg9Z0NtbExE/UXG6jUVF7e1QvDKmC
WXwQN7AMwQKHQQfa04iOPDboMH7qTMjCCcPj3gdgg70akpAOAFkVI/4adjPap/K55Ia4ph2Wq/si
Gzz1nIXj4uOlsP8Gp/ABOC51rGBPo4vqaxeeADqGxMmT6e6s5uc9he72vcdryjy2bx5cuKRr5EPm
Kvft2z1tK/uufIhK21xjFN1e4UIck08XR/8QfcoK+ZXI+OQyGgiZAOeL8W2pmCsqzbHzwGzsdjAs
d6Q19iPpYv5ohR2BmG27dyhhyGzA4MZSW8J4WaLpLLVAmqBvfhGmQGxqi9GZNu/LoxKsQtushNcX
7JbigOdp1giEZrY9x8JDxQdkIfMCj8gokMCOlX7Y8PofM7yGL1byrxXvqN8c6H5o5VGW8T9625je
moPaPocX7phADTMZefPbEEG1xHoImX6JSLVVlcD683G0iVMS3oogPYjCogKGfYlCu0RWLbbht1Yx
Yw8AkNARKHdYcA+gu+pgLy8nwQX8/dDw/zeaZI5yrHjRbrC7QK8KoThh6/F9gRhbD3F4BaURWDRa
ZHKpIIbflooTdJ1FACFtbYIz3rBCeRf+46Y6wD1D05CX12Kz0O2+DphbRwFO6w8hSrgl5+jMEosY
6l2JC/6rQWWKOgVCDYycoOvvbeHAkXMa3ynFTfcuw9zqhTFlg0aQQJL/GtsSvNWJyoZFgstfL6uu
JK4w9U7jIoP6rkIZncmhwSw4u2BQzkXQZlNU69Wk/tqbK9GXObRC2T/5p06B8f2j2FB9yF7xHrIk
V25xExJvPhLUnYMtTtKV4rK/4QMVmuF5dOFiCZ9y8VsQ4RaV00j0ffFktcrRPNs5tadkbMqSow6y
Mw2ErAd75iWUbNBGx+07xayGud/kapp6G7dN0G9USJ/kbZrVFhIM9ZMttgg1RFPSRGfZwh3xEWii
PKNg9zoiACS7AfC0yiHGdfNlvIVFpyt3EeSFhFZ99kW/auqxgMxQr6uOZSiydxcna23wnm66Dtf+
FFkz48GOI/8BJrLHGzMbJQKNfQcXlt0pgJFoBs9dXrek0DzUYw5NjSoETfDjqw/X0oy8EM2RfPDA
jBAGx8L9WscPsLaqgclx2uKv+bbLsbYklYuKArY4gYRuwEcxf0gH1+rwjYjITua7AloQrPOvi9L0
gb1V05U6wjKYjtlxTO1j2VciRic+n+g54glxsgF1n8glTJUwVjioDtUkGmn3tU/DjVtuC9b/4iTz
m6vuCtEqRNXXUYD/YUZnTs1wsnIZPQljs3alonxRCc1P+qi3UQEsCGuAiEtxFRp6TXr6vBXIp/L3
+zOvcTJZpcwqjfKYt8tMjIdEE+LygsKMEK6oIxzv60YqMIUrYy2W7SzdvIudD3NgoEYppmZbxC+k
5qg1zH60v1dLW7JdSePuEVUXT9UWMdYMZC3GtVUIy4KxMj6Oxc2Ji0wYMrdFoqNjChEj5nC3P/HM
MAX0NBO/FTFaldVFLY5ssBljqcx7i/tjBKho+16n7ojI93t+H3UpD/gWkq4I9jFFVHen4oeC7Y4B
MDo6fAcZX79zmgwUeQDswP6G4j2/VajOLf5rAV0aOpQoNuaWhBRbB9X0m06PfcV8OO1qCJ1ndLik
Lrikr6JxjvfKdukyAP5P7eCbkZrVWp7iDxD8Te5qQKlY6bTQ4ze7PYiz3z6HjMFx7wVzpPbPVtNI
O4t1o78EzOMaWcRoxqWc0CVcQMHx+cn6WWEp5Dh+ExjwdcG8WGXliWgpMlG+YXWzbEcNzeM5ZMBr
IyOYtygIl5VIxiC4TOBG7dXQf3ve/0BMeEbmd1tL8YFyIpdDPskiTLq9d76vTWSeSTazW0lqvrVm
XEUL3qlNuvFRhyzINVCq8jRK3TA2HmwhRX6tNCsm65um4Xoa1lrFDfCy0CgeRKQRaUjmZ8JebZEs
6umfdV0OwXVSZm9ovpuUO5hlw/G2VtDOo+q1zFGE47BU23DrmqQK+z4ceRHSq0zIOSb4TWoLulIG
bgbEO0WnHEFqngHB31IymhzTHXr8FkSX9iQUbIdNdCbSixpqSMQ0xzaN6GhRyoomAGBOLRYNCF7J
PeNQjz4bz8NgFevBtAi1JaGBDFgIKGZiLGQX0PLxVNOOoNoJi5BsijuE7M/O99+th/PC4SUGkhd9
dUxorYQ+NepJWb1LsiZzcSpTEZNkUtqZaa8l3jcrVLzmJdY27s4UvzUmVPsubAmDcDmeD7PcBDXA
ZtKLribbTowvGU0qrMaQ+8AenJ9u7/J1y6wX71Aau4PGY9+/PYYk8HlSkxzsB5R718MiwsA02M5+
43Vuo/Hv4TNUv52CfgClwSc8Bv+uxg+uNmTzz5W+mnQuZPwWmxxWHspiWHZIMHyA6V8zX/cO/b3E
5/5mSA75RVTS0Eju1Gt9Qzj4Oo3bXx5+4iiUEVw2dDgE6B0ld4y59ANqeexX7zqQ5mlhM0RuPpHi
tzsrtaFJxu57VfNi4b5FjZZOVAghABsjn1UMF0CaZy/Ocabtz1m64VH4DGDyeuwxtg0zGQKg9zko
h/tSkK1IMZMwqg5Rvb2dfu03HT7FTegqWiEnkZCwSZoiCbGynBSkn+AflfwbZ4lJIBny8i/O2ojh
s51A3Y6PBsL7hN/VJRd4yNtBODhQo3SWcWIK2EeQjcGVUmHSgC3ogVrkscC8NOodK30sQ6sdB29d
a3vmVNWtgkDUMs7ZIiQZmC/p4YkEwukdu5jn8qZFHTRUsKHlWJDuV4TcMegeGUZz5pj3iNaYI5IV
Qb4oyVM2zKU9XGlOxqQlj5VDAaHcDALjACq6OElKzqgFG5+eSrfp8cO9KP8YcADcpy2g/CHiZxHw
WL0UozBfdUMgOkL2jfuUqmSqSzvsfM3qoyjEWZsIwMjy73JqwmNFxKjfbzDpKkHWIC1OnAIBTmMv
HfuyZovYJ4itU2XC7u425/NeXVn1w3tPFP/Js23nGW8IhYeeh5iTvCxY8EGY5pIMjPzensznBm1r
z4MmHsM6TT8jcbwJqE6hE9y8yA36NIp4beJPWI2G0MKMjh+RYRvmRZvUlo15LprjRMux8lQyFXRc
jpWJ/izj+vLtlUimGHTq2imStG4NEIbnXzqhJMaO/Vc1q+buuDVEcWPOEZM9blPbchhXtlpIzOKo
FfhE/KEFZRyaVvlZRAY2O0KgLb3ze4lKkP/TTVcSQtLZXz4Vv3DU6hO/7edgfMwt9ChpHKX3J3qG
TZy5CS/jFPY6UulePu+ipn5kQBnCbSZwplVefl1PRI4McK+YDO0/pE29yuUngOYg5IbWROIw53Bh
jZ0YpZEG8i5F76HPslJX7tr7XIYI6n1kER7GHUOZwSgrbMZZafu3lE4elbX91lbC28QH1HKDwv//
fBw9qo/d7qqN7I99wNPYY/Rov1QKvAVMB1l0VMq2iytYqJ/R5yxye/0uUFkxP8TjVda8L4dSYeYu
8E2qAqW4t7QXfT3LI8zyIRKxrTuqTvvu0DZw8PxFhTxT2EanwTb2QR+Sn5ley0NPY4P7ZaT9EPoj
YmgUJkcj0st9eXSjGA+FTbue9ZZCR9260RgAJ2/Egx3uflQbLiL17sreZLxuMaUvY9sg5IJqTXWh
TEZUiO0e2fOQfYuWEEkFIFIb10E1q1t7CKrkOod9JIqACUXT647Ddcd5mvH2Ghqq+rTBfOwqQGOc
oaciE4f031OOCOL3I9f8O/NJ/XKQVAYiTQKrdVhn/IrHXAxXP8sE5L9QZaTfDPolHUO1oBF6QOO1
GWi9Kt35HH65K7PXdczLhmPxgGt1pfWG0cVC/vtDhlgOHC7w0cubstoar93ajYfELECMi4vkgKhZ
Gdo8+6r7zdkBho47/9awU+Hn6cCdaAOFM3hZzgZnN6SYpULWuDpD+eFHH2j27HtcJe2nlEQODdN7
Xt6VRBIJtx7dQRiN6cbt5gWx+rk2anPtMCL9+tm+TCR/A+M7tpgtwnOc2sN3wM+5AkrAuN4LLtQl
Fc1PCke4ywa2ex9jFbINUXT5bVjjfWNmh4ALNJ/s6qhmLlJlvFPkZUDI4k1YE33dA5oUpGDb7I6K
b67aSiw7IGRjcRQdsAv/2T5d6wSOCY//MetG99qPH8hQdh5dKpIYjm8IO90MGEIpq5OF0DGcISbS
Otct+Pkcr71s16U+HuBRLxAzg3laZXlPHGgaSyuD2MM1kyfM16Scrxa/U0o/AUypmYizbO6QUrcX
LwV/dO4bWL8Wu+5qWf/5AkUwR/VKrJcyhR1XqOyy92p8dKQNQXHAneVQ0WWbBzzve9KHIFJeA5VW
icCbCnQtPXJizYj7W0NeHsuJJFWm0UVN1dUOZsAuEP5H8aNz3SrpM4ByX4/nq/e5NXch6MMUie9E
+hSA1dsbHXn7dBpbkN7RL/RJsfQqK8rPUYTOaLgkJtp6nvQUpzYuq3c4Kv4qIFSHZytwgElvnx40
OpOsQFE4+5PPItmFEdpoxd6V0snXqnGYGTNfsWrv8fTrtP7ZHJDwplcB9w4H3YgI7zlTs2dpbIP9
TwaTLCK+yW/fiuvwXn0RflGHselcdLJbOB4aYKS4lpLVxspl6lavXLCTLFZYJwIIcOmME+HJ5VGR
pwFHUEiRRe+rSSwAG4wgc3W8hHIBxYrmHyGJv/B1DByIJf5Ad8zCiWUBvZinjRpwSRJEgv+VBWU0
n4Lzq9hs4U5KujjwIOsgNU6EX133AerJFkL5wKr8EgZBSIYgIshQNixZjIvzL54LtBRj+GjEL9TK
iQsEqfmoEDdQJ8S07x5i51PmlUM1CX3n+dt8W1sMNoTpvtYTFK64h4d4EmIg2bujlHLj92JcX753
3dfJPipBcgqVcqRCup4yjqXFaVepXOofN0WSMNXrCJS1nDAQj58Cug1Q2enwjVZQSkwLQGeJoH6y
2xUllBWG/R0dfGGBQw50Xnr37sZopeWo33I0jgRDJZ7Za97c1plKiI6oSVsuwT+Xg9nPMD6UJ5n0
xAx64hH8PZRSn03SY3+zy3eD2Z4TcMXaIxsI+NCavya9ioxINR5VLE+qDVIK5smYpLnAzksXHfd0
BM8CbKTCzNz89UbnTB7mtYZS7YY5dL6w9b8tS+EbO4JrpzRq3V6GPbOVNwfXDUwfZmSqq6oxzuG5
1puHma+G1wiMVWtoZBzstmQRtn9NuW4BDXlE3lWQKy2tLOiLsghH3Sc/j/99lDS92GKwP6dok0Sk
YCtrNSL93nD2RIx3Zam+MwhIHZHwNlKsNbvu69xPQtNavvGs7dkcuc17nJDvPXIWoS8c9at21Oej
BFAGQzGdqyWgQie4lBI8XBthp035qfLQpzn5UN529iZLrRTNd5f85iSNSipTplrXTKxlAdG6Rx/K
p+v5EOfcd6Rp/2b3TzEdJ6uocPPqMkmEQjXyUhVe7ywjSYOnbc0SxF5CfcG//QrDkCtTBJbv/9cH
i19CrjvEu5jrXTau1MC/mOWsqkEE1GtxfnKCQSXdSIk/wrwasNS2x/Pv/Z5Q3okcH63Xt2pdqx2l
McYf3wiKxWrei3j6qWcXQPSDUkf/GiFQ8YfgPA3DEz/firnqx4vmVCFNjl60t57zOnkZyhEOcghq
DR+EWbdzX7p8zRKbnHlER1yVn81EO/BuNMwkZwhf2lYVbuU67eH8+Bk9h4cjj9ipNVbDbD5OYYsk
+4RDa2drFO9KjLz4LBNh3rmdHwzAcJO35EHpZUPVKSOzqT3pmNJeMi20/ClIeEo+ANEf0WHo56fg
6Gvi8S334VicMC4nr06rHUcHf9+DlP2nKWqNJ2u2gjYpO9haenUfgEFYH5LIHuxJ881UYTR6+kLA
zA8zbyXPwR8qtINnR3vx8HjvqEYlvALE/BtUvFYbijrWz+2beW1lSrE7TboykkmDdkzOXsDVJOXp
ZpF6Atz2zxZzadlX76CQoV3e5TeBLkCnebLe15hJi4CXTMVW6iL7EpfCxXNoQ9RkQ4pFoDlTv54S
QBN4VoBqvcagyJV6+JeOamDXt1P1uzg9TmCgrCs06w4imPoEGyduazpdfCr+nA2mUM4bzbn/xxJY
GTVOpIw9yzrZEY4ShOotxuOMNqRO1c2O7j47FnccBtrxgEYXTE/m81SGYt5+fG2UoaMCmvD5czQ+
wGoOBnfWMf7wsRGUlzi82fnBuzrSTY/JtzfwyWKF/yyv/rKfizw2gWIf9exAxlCZvmQ5OBPsSowi
oOPXB5eQcNF00BwatdZQwzgv/2RPkfwgqxsE/zZZ5XarpsiFu+O8taHV6uj9mhu3I6MLOUbgZX8R
99s5rO/EjLucd7FlC7gHoQOjbr8Q2S3urSMzw10xoBppcNm8onF4Vi249LlKdZEOQAKCQHAZ7CfZ
vukgj+e/jkoaz+oBCSLhGdsJwdE8JNF5lIMiI+NW5Qx2mLgiEfrXXSq1+LIJvDY+41nyBs70Ss5U
lhZmaLjEbmlLDU4mXlA/rN5txaA7KAXv//Z5uXezXiGeftHoktcLxVGH6PO+Df4bM5nzPi+sa9CW
nK9ZNfa5hpvXEVXmGsRpGaO9RnEl6NZqgTXsDpYWIbZBfjKv7VledpMG8QXqTlje0W4P5pzy6Ksy
/be5xwiTkAGxob3yZORS5xZAfwoROaTl/DUGpYve+DsYIZRYhCipnr15x6IEdB5TM3U+JGi/me3Y
ucjDGpS6BXHkZidqVhcVqt2yd+zsAUWL/asxAV4K33f1f4DSlwkD9n1or0/O0/kxbWaXP0Hg+c1p
tdMkYRLHxwI+QtvCWPIo1qTHiVwTARqiSLv1xkwkZ3KHmcSUis0xDo5RaYtCeO58uW25Pvx/c78D
XQsbHXKw/6YdLxTUM88nfXPIlKYjQFJvNdTQCbjZCHro0aHrITpvX3hZlAf4Y81uzTIyVmAh+F/6
QVAKAI4a+74mtQaKGlQBX9dWeAGik8Nc7668EFtvNTx1pMw+7Id0AVwFoxz9HO7Z9d/vrYuLtY7t
vXpQz+aCt+OSRsmi+CffFVkjHp4H62Zk8VFTIceczI3WEuUuaf7fDlIBXIrXAaFWWbWQv8989qMY
bQD1UYH2/dZkMxUJZlOei4yKdqt1ApjEzjv6zJYg687os+4wQgR6CzUMXiPb7Va70FTY1aPZn0MP
ext3v9/RZiEzegc7ZkmYXqeg+stD1qv+BH048DKk4kEQep/SbE/4jLC5cXkZaoHr3P+A8lGcm1Jn
pjdwqu4Qusis8vkakk3q4HzI0kz+YXeteKUxL4iOr5Q48dTQR44F/PE8dZeooe/cd1YcQ5GWZ5DE
tHDoOxpctJqNxHmEi2CYXQ9Siuf80EyBcTOG0su9A781scTmJHr4ye5S7krjbiHnlnxx1OSk6AEa
C+AuChv7GWKl34AZ09sqb7f+RkfQss6PiF7glEFnI/IynSh5fvgom2zvxbeclPJFZeyUUeDjjf6V
l4tFo5u22K2C79rnuPYCYNQ4dME6pq/Of69QNxJjJbUUFKIvmHyU94RVUuGGF2/s+jT1fV8uEpIf
hQEJcrRPsqLSgNuLzL5vRL/mu3mrMOzo98nmwKQ3+yAe36pICNv1EDpsCylSYLsBovnAECK2vAio
7iSGdSLkDvLZUoj+/zkc5p4R6gyD70h6jalZPX9rqVfLKnjCFGySNmRk81MBneW7+iU1ywyyO0D4
RsZ1EaGd7D0Kor/h5CKHD8UMJpoZEkq9/VsiSJ/PDdPSeDtImD3KboPSGdqB9BBuXL5gh1RwRaPH
NgPusEkwhaUzCYBygvyYyxjMdf0ypNgY3Ev78/YQVllZ/BLx+oGkDjAfrZtWdAwnnbH4688OOfDf
ZTGvvnSTen6F2j9zed+fAce10qvFnAafMOCFWRyDvYqkWBFu0YoeM+n367nrcQqLMvzGya+N/1ty
gdyPma/iiSj2UCTY27Wy3zDkLNd7XfXiZmGz9TDcz5LaumtpcBKmyrGRcFP9JMIIMnHsklUD4HCo
scujrm3kYd3/oPD0yi5VBzkz9oU6SArNUaXTGmXY/6jwNpab2GDxAO1FqDlrBFKif5UiJJbceifL
II5xP9kKmZK65qhYf+BrRpZok0VU81fygkxsDqrWpaxp4WMmfM0oSF+3HOORjn315D1YnyRb+DF8
8L7PEzD5j3YWhwuFoaFcKYLmsqNCGGUYRnVat3U/9UDgcTJ9ZemIz3xdtbJrL/ylfYGxzvZD0Mx+
srK24ElO5lYHXZzmFWxv/EKVj7Gv97IuqwYB3fEHgjmvH7jtex5SZwGiFkNK80U2wwKCZTgDOCy7
1O/MqcnsVa3VPiesEZhkIk60YgDRbYDVaJ6k8M2Xy1OnDpRbJiZbBCrUCWULMa6RGKTuNsuThlH/
vAsp3ednHf2KBG7XfX8tbr2ShjoZ2olR/vv5F1jlt6lnhwJE55O+l98WD7PuvLq2eOx8giLzj5u2
O7mFB+/+ycAdKcgrjoxRL3t4SA7GZzy49XNnLe8r8rI3DJWvjkHMoCASOJH0Ptw7bUQsRfAis93O
18D294LUOU+cCwYQm+RdpKiqDhlvSsrzAQoupAuaafyC+9CUBcpUdOiup4MRz4cnNmxBrUSRMAar
yAgSI57uWpkBLtrG6+YemYZ8mo8fQvpofAK2VxYADpnIgdBmBOa3rxI6Iyiay/2rJLdrRcpJ9WXH
8Eux5C2CVaR/ygyxoTIG+eR0qkHz1iJ1648tNpX+DU46kJ0VNJ4GXln3Y7NxdQ7IlCJp6z/0rhjQ
2zcqHSpwNQTGP/btMkpjnYQpMiZ4MOMDxij5DI0kIOhrXzn5VugONEMg2SvNe8hAqUHoz0pT0ZXa
XMeMTm0XYMPsSbLXcApfO5XtiUgYysc8kaHf0Ln045veUUPnJCitmrLiCgimCCyYcnbtWTCCC+5j
POerH29qXIWghpPzOTE9C4ZUBs0Xyms6MbxmncYhI8sqPikZji0JmanrRT7yZsm/rnv2e+yysesp
/UkLLywmvalvc+XJIKVQajKjxDjGzMpuvth9aAJnOt6qE8aSHBi7m5O/wZ6N9hVmnEZAgjmNf/MX
vhirNwidJFVw047mOoCXFbFDUDH72rT3Gf5uglD+2kNDDIQ3Fdrgw/W5ezuXWLbfOe6W0ao2wOJ/
n3VeGKbm/DeDpHojGjsvZbVObVfaQYvjbx1b9FI6JY8yPtmkEJXtbK9Ys2ILtl1evHJaVHGW2siy
FsNOXmcNn5rD3yzTvL5opdJfYVzk4NbPbsrp/uxhwjjIUkQ1aSuQB5ifI6zD+J3Zy0y1KysT2eq9
VpjF4IUWmetKmcv+Ya6P9OvjEzuQ99Otkpc65pIv1ul/hrUSZT9ydr/zh6UiBOQ2fIHyRjRyX4O6
4IChL+6GsHe3HRvJB+ZZcF2H9bxPLCeHzLJ/+OYL/OvAJnLUrECzuJTO6bHlY44fDZ5XuLV57G1z
rTzhj6e3Y83l6Wt6JU+htD4rKD6hazLFVQi4oq2qPG1Ad934MqDovXr4XUpFDzB982y8OfF74znX
Kf0dNQNeOgLc4LXH2U+RV6LxddkLCaH2/CohZ2BdQCtGIdFYnJ5YFwgmlOmRBZU/2eugDhtaI4Ue
J0UZuwciJOW+cPs5e0Fs5/nGB6p7GXFGbFrchFwJx0LCfc3K/ifWGU+u1vaqhj26P7UgI6bJ/n/D
gEnxCzfpfRXe9tDLECtDglBpWDGPcY6/Ycr0UVO+aVhFA9BaDoDALTzWegkgMKr5tJfoM95aeOq1
GQtdm+GRp3mxjv6P/Vu7ThlPcnQpB44laei71aErdbuqUoHXhA+qdipWyBgM3VnI3aLJjvOcI0iv
MwGMV8IO+0RtSOCdxsmGY+c8MHhkOa2nY0JiJwlZIEYccPcTk4KcOXJYAtOnuHAKeY26lJ7RIygI
D/4wjHVCHbY/Oz254emZi4up5Ssldcy8FHRifpM+lca1iwZiOrggF4Hwb5DnKn+0+O8C0uZNI39q
Snu1k9mg2lu1N1VgdIhp+ABr6+fKDRo5SYIYGiO2yUbwz8f8qfNbNapJPvi0qZwwT+5d4l1Rw/Ws
oXtSnF1knYM0p15V7SyUUOffGCfaT8ngmpoGdxd3uLfAmQOCwW5ZIMyZnO+2iv/MxZwtThJSh9bP
SNiDsV2LDMJBgoy2dDYL3B4n3zjUshktlq4mn68EOr+egZAsSGqjk6MjgmAc4tW+mVXgYqXdfg3d
fAfN/ZPICcgjdPXn8HKpLw7ZZ0NOS/sr79fkFtRmuoJh990dYPiUKYIlz224bk33MJlMyV2ptkI5
TZc3SS3cr0JVJDjafiIIXPmcao9QkrHVu5Y1IyV7/nFJPMTroDBkUBPt+8VfGuCgMlIy/0afn8/4
ZRijjYWMm991IxpYN14yD8d4OdmG09bz6iA/eh5YhWXntiU+F15R0l/PQIj4C+lRj58KVT2iZchd
dWJe2uU4ViQ7A/lyN/8Vx1K44BBm+QCyE5vbIL6SfgM0VGNmqh6IeJIN0dipWpRJeHF3YdB1CBv1
ZNqHutvfaUETJJE+U94WqfgI+OwcWj4NXChBYHPt1FAEtPNLCNbzfufO/xqszWgKGfnt+v6NgOIl
pcmMDqu+NyClWinmuqnF0XKS8TV0jwyP6EwjSFYuLEc1M7kKILeVeinEIz9dpeHfIGpdWQyNaRd+
/yS3dbcW32kuhgkuCPIXuwlep64LURrYw2btjTQE+lBim/rPOrYtEqGpRo6kxoik2HU9joAhU5Uh
PQ8+EqaJQXNvFgUOH1mdQQUkQJG8lPl6zLijwPsW2IJY9JWpA1O3/nvWEbVYcTu5zOx/Myw2GUD7
CVUPdHUmsdm9HFkkvJYDGVeuR3CWA4Y58pUW+HxvJ5RAbmZykn/UdYk58if/vIEQ9gOobUcvKfuE
xbvVgMF+qG6o/qRW8Dn37EsZC5kk/7pH8gXGNX5sPligO8+fxULinoioj5IDJR1wkDJtP7+tTq19
XIlhGkIZYCSWTdqLsbxewFvexOKqlbIVCdQwaSEbBC3pueAbSgvijWsLQfsGrBDKk4LrAF7wsZkC
zAeS6KNp2kYWkUeLLuX+49audvdB2T8vqx/LwxpRO79MZp7dyWDn/h+5oPoBZvvp9iiK3THSvgmM
xsDbyEJYgJqUnxCUCCZDJGh7yPT71uOKVmN7JIPLBuH2UEebuITu0A5cLk2aa6OE9RrSZ116uf72
txZADIxhgnLlf/hN8hCvzU92MOK9oKNq7+tkQET9E8L96kxwxFG5MhooLU+Ud3KI1+m2u3EedZnl
QiuxkBbLwcOqhjyfz3GwlwZZlw2QrAlaUzUMrAJCPAIFDr/nqhFiHDIxPfBnSpo18Rt5xtTfaZ2P
yHO6h455WOH5qzRYYed1ggyAsWXct2an0MPHRdr/txO/8YXg9QwYpBmqOjdaWS232gIX2Lu9P4ID
52ZGzUDLZdo/YvDvXXejBfCEoB27FiHbCt/ZgWXqof88nJt0t0A6LwckgGMDcX6tl9kS4DlWd8Gx
bQOJONg3PgiU0Ym/k1K58Z4sIhvGJYzCZEVqpDKL0IYD41jtEQXIVy1GvH1dRje+5DYVn+Vv+FfL
OhITRra0Qxdo5qWn6yKv8bVWIz1dl+APVDGiU0HRAn+6CRdCmH1l66BWz4WpTsNjYRVmBnnu3ZPo
ll2t8eeTA2VX9+nD9UdZh8pgGaSNcmyYBSmVlPW/njxZnzJFXefo9KN9MNzHtFugEspd3/RMnTxG
8PsByfCGbFVMuhHkjzBhc0wSQ79NG2Y8xF9aXiNbZOy1pBkyxJxivcrhr4Qc4avHcCkpCbo+6m0x
ZVjUvFpH6DZdIZrZcSzAXR4evYNaI0WGghdAOEIa9ab3Bz1Y8bawP885pAN4rAni5jEiwNBsxNCr
KcvHCUJY+VE35lPP7Wq2ZjuZAe95HZlUAyIaLv0pqgDmadcSMLFfJkWbEngFt9CYeWbmTDeQe50z
vuj5k38i/lMmUspzZOVSLvqCs5kg80kMWLYoppuqIeCoCkO5YJm5ZrDzbjioQWmYsFv0dRzgn9s9
mu9SbOeO3l0p8IxzwxWqqwsQJVzc/2syvDABD1hPHknt67FL2WU6PdgRzjlfOlGsBVwo0LMQkPaD
BBxp6kwT2qpW4u+zcaUbfPzVtJxknEHSbcedmOWxkOjBX7mljsM3sHx24LBDNT9N9OceK9JLRJnm
Y1xICSu2rfuZrzfeBpg5Jto+2G3zWNhel1kWoYFGUWHse2yfopxWAgu7W4zOAnmd2e4zNcOkHMkz
WGX/BoW4slcAVf3gECMF/XYtyKfkPpV5AfZifSnsg6f4WC5qw0Q8WuEjw1gQi0LE9h8fzP1eC8wX
nPK/6ONhFxZz/BBdg7tMaGKOkDkN3p3dwpUAbe6KMSeGtAl2jIyh8Bg0d1gIkTyTBu+PwTbYR+w0
WbYug5zvmBOuNhA6EmzIpz/MYJT4mvNcLF+ERIlineh+ZNucBkTDCNj9XygLTj7VQu14cdAtZn1l
gHqEgpTuWvdU2rHLX63HduJBEAU1T8uk4MIqmw0toDYPi1BBueUKHoSWV7McRD/A0JLWD+MZFuaC
TR5xfUd4WJZeCxaCSmlUwMKG8QVidnXqpz8Wk/6U5dfXew2uI46NJokM0S2iTGql9coSJDUuY4Cf
5eJHOt63W21hwiafXKi9DKvNpbnzd9LAGIuzgWZ9gCKRlpmGXGotff+gOoWLCx3PaDdcuaeC0SUQ
SwMbgQjc7aAes+I0Bi+evldkN4HVZOQFAoFw13/HLZUqEamzg9v/0m4a6zRdh4SBIPDj+GBSyqjH
MOMBglXSZ8qyJahoCPTeoOWyJR/jMBdx+N+xf7jE6TH9l2TttkWs5ocMvudV1XqH2V0mRX6GCV1o
ULJGnSCGy2fZZQH1FMxmzF0zb0XoCLbdo+INURE1EGXLCHa4AsVF/dA8ca4w1lIQxyIjhHcM2lCI
fWE5/1ueli6DOasTc4Oc16BQ4lqIVMTwyIVs0z/VOJa35icJ6uXOcRqBSOcFercbBLz2KjMoDxMd
9ACn/zBSPde4zLzE34prcaOJsEu1cBdR8mCaUuMuzOkhnSEjijtWBROPhVlzPy2N9Da1x/HpBWwz
wgsEn8q8GpQtJ+hFZk3tgt85G38LcMeBvt6zgeLsq96rho2dShaHK/glAb9bktylzzB0A/he9RMf
ts971/VJuXAHd7wfwR/sv53V/OZI67TZArUYAfgeorl9pS5Rry2xtgEix9LoFUyNeLDwxYmq1DqP
Bqvinr/rpoIpyRoUm6995TVtMWqxrNQK7CydPbA9K7T8JefZtW4iEp4lBS6NaAsbXG/yucQMMHPN
FZ2EvMsy0auq2+aiJkwMewsogl0tpMoWQ4IQ/oCtcn2+awGGYlnaupZMiKmC2hFyacDsh9r2YiU/
xfuemyfS8ucCeCj1DqGfxwvI9XrqNkmjXw5ax6oNnpQpY3MJ+x/qmdY9lhsWihZC2TOtrVGmhQgT
FQv9YA+jkhmyD+VuugMRlhU5K3gLEWU53802op+3CtRufH4zG29KSJfOFutpEN5UK+SEZGx2baeo
BRyIYCq0Qn5wOkLxDPVuao9YjI1rOwX2q/nLnaWTzaX7ysK5iIpBRTOOstwJdBe4mGZw0EhVgwWe
PPMDBa7hrKYlT7qFcYbkAR6x8GcheR2AP990O1Fj9KigUsqC6O/7V3qfFB9moP2V7E2EdGLFSMo2
y5MCB62RcE76ypZqX+vN4MxCyJN5P6EpeDezn6hJ8gloLkf2MdhQOzCjOaoHfQBXeFxa/mr6skFU
li6/JJR113z4pWzV5uEE/433gQvYLJtPdZlXF6UHX8x4gAGenzg4tMXCYyRAjkOEymF3KPbKBWvw
AuktLw6oWw067oZo5wqEuiDT20LZ3IiD/Xtm3hzeeHZ9a4kTqlaRmdKDNgcdWtMaBdMQvPOiQ5Zn
bbxPTMEyL+SuqHoopvxT7h4DT+V89GLoxsllOjo53Q/HyHuIlTvdgnukDQ+N0m7OSW/t23PQQ1Jm
ZJVzUdqnZwHiQ5QnGU4gbnQ2W+pLn9LeommPSet+qvPN4zYYHQDv4puJWazKQyppbaoFqmPFrrqj
7m6E2RO6VY/WJLg9Q3wa63Hz3hkuyj+Q+2g0R6Nu7witSWE60AlKumBfGuMMkgXrL827yonB8pSn
PAyOZTapKF6M/Hw1VqKJ1aB3Kxjp8/SwS9EYCDUtQ6SIQSVSYmVpXO7WJM6eL2llGYJhyC5Rzx6i
bE6e7JP2zVDM8XwgB5s/S+zRuVLf2ayYGjBuoP61YTpiS7BOms8uWOUb8Wv8cM2jcM4nsHDC4sch
RdwUypRK9RVPYaCReODb60cozNHRUGoh+wftcJc5FqC4Hhzd1o6TRi62un9/1nQXnotuchsNHd6o
cynyskzpcoTR7GTb63aVBs4CZp49i/D2TH1q17X1cEgBCbzZQVSOhVbmKj7Ct2uN4iZ1mcncdz5j
A9QXYDZQNvPprIXUr2+RRvyE1bN8b+tSREJRWNg65x0EMZMnvcn5mlwkFCkeOL7QkbRF+gwIO48u
+PD+A+U2ml1RTjTOpKZTHDTx7v+patU0t+2zpXcwwEh6PBgWbAe31yYJVh4jSr+noZkwH1oYeuam
XyecoO4w6dRdets06S/7/2lBq/QH5FPGaF6B92kUxKC4fzcSphHkmvfcofK392IP1P+mWuxBPzsB
Ebn33MkiVr6+557z7VtAkInjaqC4pMAhHrmiXO3cpY3bpMO3uMfqPN+6FA4v7H1n09+UC0SEst2s
wlVEq3+GlMzi++XMICLSRQ71dzvlJuhrA/9QmM37nlP8z7oQ/NWXr48sKXh0srC+Ng37lwH6KJJB
l9EBbTTbf+sTrfFZ+jstgtzmIpl0TE9g4XwhmNAUtZPRAjf4SkiKJ5mkpu7GAdCxLX7Mp1HMKBCK
2o3Cz+jIUig+qmecnkW+W1JAOsmFRvKUAxwyJL/8JzgZs1kaghxTXJ4aEzyU+p4ZRI46xVEdFD1c
r4YmAs/BAhSKcywlNOAPV5+Di6C+qWZARcVgKPxmPXTYs5exOCHfhrMWi+ManLiSTGI8pqeMvOyJ
F4zP5gTX7Kn9rHySX9BDYWEbMHh6Ey4Z1c58hsWZgo01WVLJieWFhaOGc1AS1w/a2SqtMGaU2ZPY
+RPcPPcQ5CGHwqGiWMLCQi+2TYmWe6qmNa1syoNQFlsEtV7P9J6Xly0PIXDlj4VtrKdeIZJMni7n
h0nt+TfmJyKfQJoKE2yS+qli5kWo2gz3siiOWdByKCVeSJlKmk5SXFGCtCuEfQgWudKqjrt5xZ3h
61/Jmi+BI8JZoQwo/dZ4ItPvcfyo4Yk4ePl3gw+j+iEcWPQSEv/YszVinjGhN9VGuW/Ypvb/N4Bb
cv3Lj9sWayLyHSMv+TauCCiZ3Mm31ommcHC/9343ZOGSp1yyUYT4Jcqf0x92YsvFOUjFcbaw0nVs
rL1lTy8iDWIxXsRNFC3Z5euTr6Iff3O/spq6IoNwOjgkJucC89AeT1/k551AXau7YKp9ltPGJXYF
sIpUVIlAmWfKCDvJa6rJjYfZ2nacV3hQEHHZPbl0Q+34vGRngBDzWMcTdTa4Hu/IPEREFSjwDUbv
7/+QWXoTWIF318vi3GAOKkwkXYzvsRosaZPSAlDEBxwmxkdyCFZAF2updRHWukJkk+d8VwAmIeG7
ebrVgJ8a2eDcFGPPbAOAFv1RfhAcSoOupLGgFWP6u5MUzgih1XK2CqIOBE45zuMRE2zjfJeAe9o3
L+ooA7UV4tHQwOn2+XLQcTq9Ry5VumLFNujxfFyxJ3ljo2bx4ewJY6c6eknMTkCbeBEUDuN57g/r
z98xL305ceazWAswvtqJxvIURU7X5/tFdtHWoCbHqN0DKLOPzEuYlm57AyOXQ2SmhP/mp9pmmUr5
Hwp/P56ZWoz7b4Ox6tw6ATJ9AM0nrsG6fYUx1kmfZcHWukRVXyj+4pbf2k0rdp7snKVSE/J27qKv
lfvGI37fk/C1ZNc2p7zzpJbrglAuSailH8x9pJqpRL4li1zaL6BdB/xYeTfTIfDqlXgXqTuRiUsC
mfGJQ42H7bIjqRp08otHHbF06ukBDbKn+XpNhxTB0cOr33YZy08KrubxBAzTPhLmc9MqH2XR+Gm2
N8apIWa8eC7wYT+x+Ie8ben6fHNTKZMkSiOUMpBQ7Ojwpye2yeohxsxzsdnzT6hGl+J03RRjzMpz
gD9zDD68Vj7UHYgsdFOIeritgPImHAY1n276HpepjPkpB/DLhMZ9BTUF9J05PhuTymVXbc62H3Bd
kqe9/PJMUFLwed63E8PyLLWJNAmD4IkhjImYfNpazFAeS3ueMstzDtJKiv2ePjroF91/GggaWeCF
SlvfSchmjOBOt+cF3Npv4wIp0SlXjQs5psTakK8WALJ8QtUyHUscumLGForQN/dCpPOGbHtNdNEX
9wKzrrZ1C/s68qhwMyPwcDUo/em8slkXQAxEX0LpG8Ts08yY4wp43dRqS5DRyX8QRy/nkXK9Vfgw
9e8aHPi/1e4qISQCbfU3eRt/x0l6XKvXHWkWPqek+iO6QsbF4OyK8drB64vdeWIHb1dOdkJa2BqM
MWNn2S2DVNoG+iv6UcAZMzGpv8Q6OrT0E7KsCFTF7RT18BKWOY+0v7JmtMxZ2AbAd9Cyr1sGURs3
3H8y8PeV0rJDDDQQlDDAjCSso48VPQhIUHTsJsTtWoRaIVNo6o0f5PTKLtRtpvRhJWbafzd6Wyck
eJkA9vEgQY5mk8K89GMbn271ULSQiQVqd2EUWjnmD/JscXrpwKEySyWVZPu7oAUQ8NQcaO380Y2p
C1uWMMGad5313SrEJvoPn2Zo6D5GzdHuro83lodphhN8xE+W25qRG6zrNkzcs1+xWOOyFbK86Wv0
G1Go8qZHfKR89BZNVTRWbR7UsXD7250Y34byujqVg98CnMrGa0/7nzz9mNe5RBXC+f/yBUkjzPgV
aos5aeDcZTQp7KDyFhyC1U5xusA+PF0xNhOrXVHg2IzttSz1TTq8WsMehBllm7pE7h4oqYCLqM/P
Y92cHFVVc3/MynjPUTNRh5dKZBvF1yPXPh4YE5jjA1IrF/cFfVDaJFawOEtaPrB0vLw3cpl4s+WH
3mTuCLhTJ98mZPuWCUyal+RG+O7a0hI2ckouqHBINXUo5x6dlEjqh+4xDQBMK6HR//BDc29Pbm+x
WNrwNgxrNUHpNm9hSnrxF+cZ4pygHyg/8ANzoL6Mqa1K6DAOG/gnHT+JJqQuzuBjH+JufUF0erk9
OmvBW6tEj1ysOEI8fPdVfnYtvsgWmNnORGt0faFlySr3Z9twGPJfRmNaYMajDGN9FwRbMtxx6XQe
jJ2kYdYte8u6tZnIk4j98i6qtIMLGHZVhorKB3nfc9N0wufbfeACFcydr17K/9AW+saYHWVlgKS5
Mzai2d8JTpzh1mkhhP3+r4IrfAnKeY1DLzddVPcY0E+TPKgjITn9mk83wV0B+TWfhkxrvrz8/HnH
1trlTm4nySF2IUZrqh7g1S8EQAYxWTROYrUmicKLx/+Y/4kdVBOdpgqbN2dIFPyRvTxS+JiL231e
tfY8vd9lPSrMVOzhqOKBaIQVwjEU6onBncO7Q1EZSzydi1JwL73Mifu5u2edmidajApZl4hSZ1MO
/ILuXVjLVVeCKh+HNDzEA4/Q2ukGfR42PQPxRJKyDs6ehLFzMvTfCC2VMbYVkFN5X+NzIZI/W234
/S0DnlvQCOFPBDQ72jEV1WSFAvkhFoTp62Gv5hjVbrIc2SGVDDM6jV8L9vWX7KlpwTP8OIpk36wE
bO+hTI+OWx88/S5Ifcz7RG27u2vNzzjFYS8FZZ41VYgSkPjb/s2d9hSkS4F6jx7xEutwopPoUCKO
1wRDmunzIUBchyX+qvj85/IcOHPv+rqiVai+FXXH+eg9B/GovPB4Lbkfkkfmq/5AWr/KRhOxsvt6
ZYHP1aoOgsXGBXwa2S9VjrOCHXeFD00aykVoySXZ9ZBaaGMIjfdD1hXFlHmSowg1fcRramEvpFUP
bYDYdWcF9FcPKNbf3xQXUKVfLHxYQWFWZ1IcgtPkxCGb/BnYNfLXJQnmK/AetBVrVQITJgbAHXbd
m43zkwrGIhDrGEGylUp/hsGYBB7TTK81J5qk8OVdDg/8oBUPgWAw1i1Tnk4zhTGHGHzjXM91J7OW
81va4FTvM3H+YLApF56cmnLr/apm2MFGDC01piy9DVbIw2IbuUQWLPrUqkD9I0YXKmPCPwYSxkiG
9C88z/Y180GFIYLpFqW7AS90Ggz9MjnBQ6i2KfpvFt4ND4aE/CyvFWM08WPP/0f48kzofSuow/rg
2IGHfqOVgxYsbxVmxcMLOyON6AsRJcXXZnYX60Js5HXhT/+LCpG99r4etlTnk8s4L/rV1jSGxGeH
ufzwak1nVnor2SLvwiNMevvB814NRjeQIiwD+a9HUMyGYqwtfkbHKoPbXdpqmmbCkb6h2+7rtBSO
Ui8xA6x68bbCE6iN/5UZQMMrgcA5kGLoaweK5XHYqjvvJf9186bOpNheP0yQhI9jUhNI9Cjfl10q
AVhSAYf81oicXHPuzPAy+gUIuLpIAoV3VycgkePKKPfF+srPBlVBBVqmoOd+6XdjgtYV/yy60kaj
538RFWBCHlETb+N8TFDlj4oPECP+HuT+va9eqm5mR3x3G2nRwZCucLx/cWVNm/ftSk7jK0Hxl3Jo
Wf204DrKwVpF0bGcwLwSwsSWzW41JlUyQjlijjlY6F5IMZ7lZ7KRxQNu9L+gdcRj0Td2iINEzELU
EEjtc52ZaGxdXIIOMDCBghYnMIBp4Dnez32BYGfPwpH9RGt3hF086mGPXTCIEvLqmukNVjjZul0y
bQvNiECtqcmtfe7XfE5DUe0OlLzysxKP2r8SkyqZKmmx+w5IS6VO0+YHLDfnfgxm/9XVS09nJ2mt
agZRX4HXefl+AxztqL8qfxQ0aCPkMLuy3GUdtPSbe8TilI9wTx1F00Zfaqcpmfmyxb3ZPoo5ACUt
KeQn7GI5Lgw6mVrgha3YwVYerA3Lgh+q2eVueY2KDtmrxEZ+f5kvCqPiF+8VG352znOQ8gjJXF1w
/OWm9LCTF5YF8TLPsnIC6llZ4l3jWDQpP8q17r2jml76IpV8ZnuTTKQIXbmSIkrx/1ry6OQRgapD
hdr7WRs7Bv0Fb54uV6/8GI602f3nkV9H0mNAYp7OmZItaSXbFXO5CkThh6yFV9WCS3ugSjpl+ZCW
6aPx0VPxf5xF1vP+d1pRJRuAzcW7PLFLfn749oExKNZ63aaOXafLSOLk0gF3apAZo4SEICBlLSwU
0hk9foKuHVfbMYyc0Jtiq1Lc5QWLwvypEfI68FQVNgY8Y5/4xF4PFB3PJr5HtdggmX7AwSZdYi6b
inUs0fMZD4h1pLxMIoOMwSuyhE8YUW0TAd6DdPnhq9rTE7xSbLLTom8xKwisCQrMz1eKNOybZjM7
J4sEab3yf/a4SCFsdalS7wsPV+BfVFrdx2b2aR0YMDL7PxQ1UMpm5ULLtvZfcyduCj72+T/T+blY
X036eoQrWIP+on6jmMne+TiwE319tGO7IWJQVWucj39qtU1YfJEMpuBteNIyrI6z3l9jBKHq9+CP
GhowsS5MB13MvbgBBJtxjoaG1nSoP8QM7hTvjpUTuOSHKSrub6MKdu5KzBrths3WgJuGpNbfoq0s
PrHY5DrImxZvPyzhYWoQQMvIlOX7cPLb2UBR304lJQLfzob6s3QVubKTzrjd/ziZzdbbjEo23sO6
RQH3tVfNUZvhEVIwxz2a5J6cqJCje2gUwYfsMXffhu8feQDZIvFzmcZHkyAH2qQzfEuOL9zSLq/j
vBdMttAGInkJEr9hjbtQrHlFjtxucoE3mT5oqQHDOKQk9dNFif5VuEQ2WaGl99y0U6PkU7mlHQ+I
VFXnKBH0Dl9B7xORVdz26vU75vHHFAXpkD2ztvKpWIiQa/YW3W2KIq6YO4WZbu7qa7wMLifeBKJN
hxpB2iZ9hAJXLGh5e5P1FGKQHtX5E1rvFshpf05vWg0hGDBxFNbltwQYSh4geg5uEDTszBUPv9QT
HQq2vDvFhqO5yph7IcWKQjRPc2y7nKWO4aZue6T7frNOUTSB/xcUgb+kLiz6Dwt5zBksQ2px7t2A
EIgCopxEx1zzj65CkISVZItpc1U83qzBgk7l2O/8d6JrQ2XeGmNcQUDGwhhH8xk5WJ83csFSt789
Pr+BbF6toK7kqBWcmfjIOcBtUqw50Gj+QIC8FbSiJGpFoEuFQGggWK8rr3h7w6OVlWv43TUJoERj
85aCi1Y9O88moBFBiHLTsUUoNz+5oJROSV9ECaUR/0Ua2/UUs+E2+8pfxrIQoSMdSNl/6XPzNOhj
HbKnMQE1tfcxVtWgLTZl0JpwtZ9ciNbfzIGynEYvxuMgfl5vGiOjO2bGX1hDx9b2/EQprg0/ZArA
ZomMceh3IhZuUHOKZF4MXh/SXH/Ap8duQsUbXIIOPg55t+pahevuAPXKSFTXbKlX4wpG0WGoDRvE
s4gGuoLPEp3gsheWPcvuwSqbK7lpD53V7FhOMKXKPVTGAc8yhTx/2TqCe7Mn8maPpUWWDGW0TRpu
PFVQKickaymJUoS5GOufIJFhKX+/UDPzJukhn98YyY7/Flr3A42yAONAIJPNAzl2vOJ+f4xX0tpA
yl9AJaIeSWSBqUa50fuiaiMdEwQlhSd5woMYTRT+l+xBpGxL1eBzYEGJVp4PLNbTArBgpZupGwF6
X0kWN7ilUBR08QziW6BubIreuwMw7jCWJ+DdGc6DAtI0ZDCyFisQyWDIcM2q9JNAB46LfMt07Wtv
1kn1YvAbxI3+N0SfbEibK50gDC5aDzW4N5Yt2lfjfww57W+Orc6K990oMHmtQ44rOdwaqcbBcXpw
dtZB7DevR0S2kn8ePnPimVJB5ELmAhwrj4V4i51mQmNt/r5+xsOGRjVfekgH7MoeCbj9xdB1zb7Q
4/+qK4AwMJc6nikWYkGBk5ryi0S+2/iWP+LMJo0fXGQ7Zi89GNCHo/inQ6j58gc8c/oc5bs1g32Y
rMTU0Tg+DqtMw2s9FkwtEIzowrb3Q4BJjDFxNCvwemDm/vtM0yf90H9Qbk1pnrb906LeottWCRad
8ptP3eKgmYV15iqvEF5z5soUm/rT+rMEYthY4dAKdC1PpyDLaJW+OOKAzd6ilajqpxi+yDLEDEYA
bAIrrvsQDvcxkzx1EIxK+DGAWa34S1/Js1r9I9MOhe6xdQbIoOTAyc5Q7Y3goUETh4Jwy/BghOEp
W7SSIb6Ms1ziVSuIP2rCHebN5M+WN/NUVvRYM4XaiipYD7H0QaYv9kIoNMsbS7LWmtZRavJxozzH
u4cVdlknBlFZRYSDLKNq3v18deVxi8M6Z0vYLzeh/y3R2gktC85lk+u2ZZ6cI79CIc7JFKG/rDIs
+gWt0sw9TwbznqI46jo9gvtzgt4dbEySfV4Me8AoRnVolwSkKF135wuYKPZArJPkzcMFO+yUP3sS
83IE10FjZaroYP0Nk5fC/sb1HJQ3WHGvOjZuHtyZ0C5SCFcxR6WTvv1uLJZNLQxir0G/utUJUOAf
7yR5dVasg5zZT358rWqr2g3ikCcSlMkZTVRnC6NR8j8rNrRiqFYrJeo8WNTuLfFq+l+CJRSXLJPk
8aQsrahhKRbrRL7VGYe+P2htsubYYOlAYzqDzIPW7kDHB4dhvYMtC0KfXjFg8BTNtXDcckyl9TQR
7GWvvzaPi3jURkW7V+oNcINa3l86HlCj1Kzy6LpSMn/lmEb2TolC0LVbxLuM29L74Lu1k7R6Btnu
3R0TPObd9HTogc3i0IuNq1NIsVy8kBeU9tuGJiaPg3KAeBz5ORSA23inLcIpNKjP3ql4pCq274BE
1acf2cxlnVymDjkeS3BDLg2/pvp1eKtIKHNDMCv+ejiIr82KRb+MW4OBFrM58B+ba24BS7TBYzQ9
Vm9B1yOlVMmuyoxsKlDkNQFTEx+zlkxGpyc1OJzlHd736Phizwf4bcYFHDf07WC3X6EM/xgM24mt
7ZU1VtxSf++5pSkYNoIdvjoqCONWJ1466bw3/ksUmHfuczwEiZMrbwJcctyCiZ8j1Phfhj0fQaUy
oTty+6sTGXvCfy8lms2WBPRGPX1jvJMeLtq5PXuzHv/dv9qGKMQSbxVASmXvC8Koxd/rOHEeK7HY
P1LsHdvr752VmtO1R60MpgUpJOhQ0dWtdLwYuyA50NdExsZpTRyZ3roe23XviC7wD4cwiQgmujL8
ee6mWIohadB1sBMUYhcsVzkMcjn+tW/RuvT8WqeiCDtMymwXB49gEZEL/igsDbQly+CbmYK+63Z8
2pK17+CcBTfb4D8korZR51PiHpEp7b4S/AbX6y71GTNhBpq5bUlYwVpdGEH1Og7Ig4tVLstc1W9q
ACQh2oX2J2UGTuOD0ASTGusc8NX4wTFtI+XkPWvz1UwlLPyq2NF6UEE4RpDg/ZsgEajt9OzfsuqP
tR/tq7cb52agTR+alOrhaefFvuywUNqhk86njdoyLtOIhsJfy3VkY5bMb8Xinl+XEiimQ9wnPI9U
oVmS+DTMbxR0aZeDxlYFyemVH4u6Clm7J6/hWRoFh8LSgvzCp94lB0AtPQjLnGgCailOygvY7Fk1
Ra6Ebchlswq9UQqG6AT7b08A4Yw3Lx7u9sLB8aH1E2qYebk7jbSN7QaKkAD3ohpeJLcmgNSZVr+A
TWWxOCCunGfXS1pSSERjz8M+ryNmn7OGc8ao0iN9zphI1l3C/e/fQgkffYqK77hwSNp4bDpdArd2
2aF4XqJBx6QQkU35c9usT8LwMA1ynGU6YrQQE3dz5jwxMmy3NlTNxFPf0sjzQZQTFwJiDKKu6xzl
0mDvktbtHxva/ACev5R646838JYF69fJpxyhrKb+5b50ze07PJyDKu5J5lUii48DUsTbErg3wJ5F
R3Rm5NKW+Aw86p5NMf2RfdrITvAmvucfTzQj8lw57WZFtjAYEI96fvbdxrFUehhr9bivuWg+oGvI
ZWESnqQuyloQlrrxWp/p6J8Iti77yV9xdMqk9y8UZRWm1YXMASSIa2IT5cmiWXSUbfXTGv0bqWFF
13kmIa35BrDBaZMFwrF7pMtJhQXG4mX6OWQqMUnwgfihx9DlzdjdFfccbroD0SOftT0U0YUu++gF
86GbTC+93N1kj+okquB96pXnawTQc9laA0pswD6zjKLImDc4Jw9WnPCQl+zE9PIb/SDRQhmqI4Xl
aaLPFZlTjEZl9Q130WSsW3EIt18GnzmEROqzgahtU/3OC+6E5zx6RVGMbZQy7NWoLR6au8dHKvqQ
zBroF/vdT7CUFmBMWbPN4XAlJc6BFsN+9P0I1AKJDEfNSmeXKwCAcD3iW/K8z23JBmzGBQdus3X+
w3lbWgSyef9m0SeZ4SCXvhkbhTqIahXtBznGIBYF1CYzGVJuCRTUDX4QW28j8gbMZ2gYmAwrW/q2
8nc+0VCKGWjs+eljVZpXZbiPwwx7vdjpdhZk3Pe+J+YMFfnT7epaVFxQyml/GmwXSflu5ywjrNSK
trvJaVafAf8WThlrhZuW1ayEWR4PVCqd1Ijk2l4Cc4ybRW/dRFCsZWsBAz2rpmmHx6AE2nXbbQOF
50IehyeuR58fk3qAmT5mPWnIN7NEOb2lfyfc85gkozf0+JUNdjvQWJlONwCtc+qWKDA0AC9owzVR
eUmI40t4v53kxLo6k72vvnJv+Wojx3bHA545hrGi0E+G9tS5+6+vEQHKzXxe84YUZoEawVD4w24G
gne0bNyVgjOsigYOSrRBqty/JjJ3DZtB2hOypOJAXtCqC6G4iA7GJGmD9fXb5bjciwMHA/2X4mk8
fN6LVIDuyvZNqaR+qo4kNSaPl8SqnNojgWs26LE1YVGmCUmdtBQLHJo5PC0Uq9pH05cCXMzBjFts
gFhqhhEFeEMuiLV+Ka3be7UYMsJwZqaTx662SXYgbQM4zj0afktezEdSHOA9XI7otq0SVWyPL9jD
OiQplbS/H2MxrF9OXVsh9gCy7204T7rBimV1iHsrUKrwJiT0Myya4qv/CglhIf/tJ9pAM/SNpFzK
ggYHxRuNbuFBnlNSwu5WzAb2MjJd+So52+YuMt4G4KiIX1+LOTZYyloRpp+8l7FS1fGG8hy9Rm4n
i04LnCk5rPdj4pP6RzdWf4zkFidkv+0PppOdy+H2rscVMcjKr9lWwTJkCkteghyn5jAwaHxfLIXL
6T2DzDBTjjUByvXFvP7yGoQnf/uF7rvQZmRS87aFaTqlo8fwAzgIGBVbdQjsDt0dGXg74Ss8YQ88
1wYnDcqthktRtfomGMU2YK8ST/XNmilEcKERvrxl+/m5Own/Dt1sfwtKICFeTNq14sS+6zGF0OOl
nx0F2YbZ8c6K5Y3BVbLa//OyV5TBBnOD8+FtktWRbBCoH0asCRwO1pTYfiAoLLCw+upR0CvuWtB0
vqcvL/LJcA+/RgHJaly7nBEux8FxC6AdT9k03k4RGepwvIen3gILj7RO9MlhO7uB58ZC934hdLzt
kBuFJuGoMjM0roL10W4JK4UYyIW5M3chiJoCKNVqDFUeVEodpOUtWViyKQEOU31EXDXUvtifgvR7
aRHZ9DGqiarkef5ctLe2wta09x5qGpBUnYIZDyZlvwH2awWX57lTPcKK7BAtD9aAC0ngFJnD+BQh
uSz1OMysLC8zlUBVSdS53OGT0wjeL1uCJjrKtzOpu7JTZ3wvDo2HRAaEQU3duRAxDVBAYGlG+nch
3Q3tnit1WcorlgwUZOM0/N+Mxa82M9Ekr8yRn/n+Em9hFJOSlyySu+A7+badHwjDiQVYD6ePeO+x
YrYTSi3qeo2h2N3EfBTVj5EWuge41sTT/QhAHD21DYIFz+isvwIQ93GqysHC6CG1AyDCCgwcDvuM
2nuv9Od5EOvEW3CkmZ7Cx5mHIlBLgxLZ79v7VoCkc/ALTSwXMyFcuSOhoTdRKen4o/6F+4VmWZiU
hK1JfVgFiLxnIweXl5mD/NVqnQy9hsPK+BZ1/MOuS2ZxzK9Nsy9KiOsqUOy6xeW/vrg9M+waNC+T
bjE+q4NF0xMW9mb3hTOBfhqyeGZZIaEfBUGX88tJWW+dxZWx6qzi25aYuGihTlGBlWtsmLyzAT1F
bUV0hChu2pczvsMNA7O46pZ0VRlIWhURfOevysoLlydfGzZMYUZQ9UANcX+5AT+OW0LiP5TgYxge
8RlxrB3mxSK+YUD+FuHEsY4kEZu4bjADFr3I53bJQNScAei8CqJ/m0//xKHnrS8d+XkQvdbKpY08
7Q/bMnJVWWw0V3orTYbfwzNQiM2c7CzR9NjZ8Yimf0FE8fTO7T9TYRQmzDtAdHG3+jmUaM2OiTIC
4KIrlE053DUJ+6qewz7pWJzhRtSxZreHiov5SHtcSzCHjZu2y8n5EaGJu5vSnDqQJcSE/BAhEaUF
SzmfdXPbYAKEgSpgjZXx5Nh0/AAHxY1Hd4+huU5a61Ght1wlSFtC96KMZkAEoQHlXvxHThBy42zT
LU7HX115+MaLeYkU3TgL72HbVAr9X9X5lr3ZWGEO5oK9XIsXvIpufY2sHiz5OuXJpJI44XvSVPEl
4wrUIpCfsVkbBlp5maa5ngl+KO1p1+z8hNAOEUz61XTQ4XWJXCCp1I0cxj5JhM6yFkfynrP1CDwp
bMFZhJYpnJEcJr9owoxQtb5sJBUZeZOM9n2dByCxs2v1gg6Gc2359h/So3OVuDCUvsLAWx8TOCfj
cG0NR87td90Sw8dQ2Js7vzCoo0+ZIDv54pfyABf3OhJlt3fbW6Ojsz1jqXsuhWpjxDkMe4tq4S9d
9AsOXAyhY8tki0IOgpxbr1/To1XytQKpXhsFL694NgeBzbcG9PpLpSpGPkd0iKyjxpxQNrTnqrLW
hEkoylOhgMJQvgcI7VHDcAHQBCGcXlaX+6nZt96tgm8jAN3FPDCNgq8vIZZ/yAfsLrKD6Ch+wHW8
tTLAztA30JhHB1OAS5ay7+uZlb21jpkdcvfOOioHWznItPtzv+i2+fTJtjBmPak+srlksG6xI5Wt
BNVQHN02Gn0Ua48KS+l8iGMaO6174JPg6PsJdKi6xEn4nH0rQNWGcoW0PUuUu07PcziU/KAxas+s
BP95aknac/P00fBxAcYq80hIBE5TvHSMZRp+Aer0Vy2ZzzkAvY8Ze71F0o3qMyS4knwCOcDMKssG
cy5AucX8piSMBEi1mtCjs1AswzdAlP3jNabIPKMEC2jE9d/pWmnvOm2tTQq3/sPw1UNkpgtWY0bL
RMjes6sFsj+1RQkpiXK5Qe+KZRbDWuscjfyo2gWAw3WgbHGIBJgqYA/fK1vgibXK68Yn1lx025hO
cKgsC6XFfu/kYw+vJs8mdkcJo+Syo1OIBNrcOhcMFq/sunB/VXgfDAFq9dyE3cWiAOC9XQ2OYJJr
Coap0yPwJTkhOxspaOOQwzgLk5bmt6krY9qxE8gOJjhbzFGPBcxGptM7teMuLOTMtyvOzU4kZYdL
CPpKF3WnLXU7QPmRVoBx0QMS3P2BpC3T4TyVATL0lrmAd/cp6tHsfHxBLoglZlrqG0uG/1e3T8Ua
1VGttT2Gcnajbug7GLFYvB+yIWG023qsm5+sqqxo+1wrZFsX5HvcdN7z+lHWiPFDTKTdHqauZIg7
tr/gcNWr5oz+niVOPSLXZv5m4utmyDBpsH/L8+jkyi1u2smE0E2oQUOVYJb4PD/mE+AQDqC+VO65
2jm3zEXo9kVzvVbEcy/nDh4/SxJenAKDWnOx6BzxTfzc0jMyKb87nn2lHZ32I+ENLPsDGOIymbA1
DI8lZ41WbyOu3Ga4Wi2mmABhDt3mAJBweRQu0gW/SLAUm38JionFxzMVW3EJQpwb77aaufTvX4o1
6H1pht0aFJwWNZG/2n7KMxGfk/ith3iqglGNI5r05DbkiwGLFrhun13DPSEvxkPDDgYpSRJ7/bjV
EaPHR2+9foG5tKpUFWRtDawFLV3yqAr8zA7hyU7TxAkEHmAY52GR97b57QcMxEJdbdf6ueR/kz1n
lRmrU6fsPLKst9sKuuLVUPHla6txM7T4ZLXPf2Wnean5rXoUQSGIk3sL0yDSbH4LJDSJ21bAwXXj
8K18bvG6oqHfMs9JxUmgGUfNdPdW0yKHvpvVJHbUorgU63hR2KkmPdZdVFGLJhKX10ZhldT1clNt
azsSPnmL7M3XmKrgPZyZ5OLUGPOxy8ehSlyW1d/gJND2gPVSjuUTnrXtc08zxiHzdRya/v2yWST3
yf1eVT/jEatHfts+9vL45RBqQ9p9fItcysJcdywFEDgNXPPjymPwFWP1u7PDb1qVv46Nrb1GUQ2B
E4TZg4Pd1P4ManXGqV4gQ/4lZDrVwHe4JChiG8Xw728mVr5LVhgnmsAMFcIfG5wKrZ2h4Ib1cc8t
pVzjXlTmdKaOzes5Pcfs9Q1YNzVPt4PLL3Y/YmFlauIu7ry5COY5OIVb0/n+/uwL037M1aJPs85W
7Ilw05bY8hxJQcLz0PZ7XvN9d3mAOfSJMIZ6l9+kHZJxOWW54sGyF6/OVtyjtB/Q/Vr8BQRTtwuB
QZHa4G9WZ1UahNtqUpPc5Rv/Fkr0u4YIZRKCrcfoG/oH7losI8DOUx3x0EDU2RmX56qdvdrrLJC/
zHyi2uTW1Dhf/j9zblSPaCdFCK24BPIu+pDzZOq5hnYL0XpSI8qrj46eBmaHrRxQIJLrBgY7II0F
0JWnmhNkWcHMH3SDOARz0ym3wkhhf5nDZVKZ4VG8U7TBTM7FcAcUionZkZU+mNfexa2QVt79Au9O
OrWx4NPhGSkTl2pHlA7He8iMwXMoiCHbaVZVzQMevrOGN+N0lZ25J6eamlvqGrlaSFQy+LKDKcuO
8qfqFnrJPRefGmKDWS2wVx4o44QhNVI6kpalJ1XnoWLtzXzFqU7C/lAen/osODjQcZu8LJ+CgwI3
Ao8VWpQ/DFypMkI76qAMoGJlNxZVA7yyYugZhrdsOU0QaV4pwsmMR8genhSQJOt7c7hoWS5oFSOp
Py2w2tuFMqjKzCgm5CoU8UHm6z/z+K2mCufa2jAW2MDrYHr3fNxZUdPzefVOMp948bJSUKyj78y6
k+p5hkHg85YXdDOF53zJNJurYmlr0A0ccXaZ20tPyu5lmjuc1+08cQ2sOX4ji2EYIQVA7SWtT3Kd
+jnjYdfhchMT/jLJS1l7lJQWoQ6+WxVkYRCqKET9F0tz6fjtzVVzV6YwnXzhUv4vPR2HaxRGaWmv
jl1s0Qmivs0xwdgHuJLTtI70WAzCPZ4OT/lPLK/dQCvoDjWTIhgV6XDpTLztCW2kRplcpQXFIG2W
0lWvZWShepeWP196sM5JWawsAgr1kVaJ65fMKC7QFcW4CUlV/SJd++xYR+aXwokzY3qiNFLeu9Fo
tL1q7E9U1OKnfSHOxYCdYcUjx0LX0NrvxACTgl9TMnaMeA2Rsqk2/26KBscLg1GhG5qMpkQ3LEoH
vzj33nodkiv2rr2kjmxc66N2DyGA783bFlSzzV+QCJoDmdinqm3AmkVi5MPCErZEMMwRtNLyfmzE
hfddq/yo9EtNReMjnCa34t0wE24wdFGpLQ94J87Gh9QhLAWddepno8qFz/YDocgg+bVvQraqlZsW
JxB7+r1dE3m11ZAAxxP/4aYPeq7xV/guEShxgqGJbIKXmxjf4vRA+Cag+KjwEhp3QCBcRIAvOl6B
0rklELyfvkvqMglAWOuawEusXZlDwfTilJMbSqljlXd9yUHZjDouZmBNbt4yyn4/TgVkBMpzKdx+
MLdMNCkHRWpED8zYQOw4NxdlAB9P4CP1s52YvH1/5RMk908wIHd4/KNZSe0EdKXX7Tqv3yglMiSC
3xXqBJKie75qw7nq4fzSuwA+6RdLvq0PVt1/Rpy6yl5f5o+7aNZciq0+Fj3DSxbA6+9mS/RD8zR4
ExFVROetuahPVoFMDW/FwYeLIBkk3mKgZa/cDlW2PW5Bf0pNvwpEgHUcWU34BhuwbBmZdyBEoBSM
OrMsjujYHDJE+Jweyc3Os1E8CZxEGSndg+91ec6PNQ9RirrFappA4pb5XKFm2MBjlmeNSLkr/fVJ
pmI8C9VLfvhzV2Br6zDfloVv/tdz78iDFKSVxkeEvxYYNoMTHkO18/I7uIQvO3pTMiOdLkvfGfc9
Dgf+7i5m5OPc0LVn4zY0A3oA1GpkxK3YULalZ7UV6wutFVegFAZaNyQCbdMKczBHPnWM2Ej7nf0w
Ml6oDSwHk4Y5zKYfG85o0Wmt/M0Lv+R0PRatsFhUPaK9fFXZjBtPzmP+rQcQj9BGcCTpeqaF6u8I
ijVncyqv95aj9NYEx+NHc4E2JTg7dN52Jv2aAHlh4AahFbDVBYxbQNkbBzdXWiieHMiPLkHNMlK5
TdwwAGam24uoATIfuN55z7Ml1byQ9HNSlFeU+Ymmui1VKSjlcswOg4p7n3s0m0xL+N+QT/bRCXpz
5EB9A/haAWwYwe/Cnd8V33GgR3AqE8FufJsPwfYZeFffPKZ7EoOvEJMRGECaNOV6SLfIWj2cl19d
Cbcp0wAatVyitOO3kYuEXtPNsgmv2cLkK8izifhYKP5W6CKpgmWqpSnWxWlTcaKjW6yRtZmk6Ik3
K+SBe72PcrDPgSUuNEjT1wfQfs2HmOUVp3wIR6dyDTOkMu7jqWBKixPepUG/bp0wA7B6D/g989/y
A6NziQZ7NjSx8Aw+tkJ7ThH36IHm6x/+ZkaH8Ve8WM9aJZdXGFIW5ZOXjJM56CW2yPEVa9jSi3TN
TPAMKgpCuT6N0Xcv8Nq+H7yr2vnh/+/YOqXO6n1L5Qj1b7WhGqlLo6rJv1E+fvSkkNbiBHXSC2ih
ylg4j5oCaWIasCAXpG1I1/tt9VbzsGhDS8XPv4D/sCRIULkyK9bAhnuxa5WBDx4COeBYCgYN7s/1
JLZgpVz91xNGURehULQOOoEWpFC09zxEq1WFchD4Vfu2hHVybFrfy/XLye3EG5Hd1PWqbV1dKUud
XQRIhpwrM0djnCxLbiLy72+gx8wvQHIqLyoT3zE5m5K/FnQN6f/ymSPPHBX+OFElwpEjgDENOTAb
f2E8znQr3J58NCNV/ddPmQo73kAS5xL9ZHFu0Cd6gb2L+crzOzTjYUdDm6q9ybrb7SjGxJYFsfqe
2FW8ThidznHlCMVrwYJ/Zq8VzVTCaDZEm+lkD2Usau3fHaUtq4zJOA/KwSCbzlizxULySMiwoL2U
5BuH9/mHV5LWkLPD5LzsENbfKpn+1EaFRWdwFLgKs1axPc9hmwkZlb0X/G8JFWZztlnkaXPg/p4O
WpTZJoIimRYldNcCQDs3EdPVOxxiiJMrb35kGF63OfAef7l/m9U8o1VcLcdx1M9UIMirz/zpQ2Jn
fmyBrFwpBgkaZiniqkF9+JvzfBEM/LLsDJvutWIZ8OX5JqXXRGvHxudQVemutwmf+jLsJoD0U6iV
x5F7a4wPvpvjVVfaRujh5/SAw4CJ13tjyNBdI5bPbEuhIoQB8Bpl1+QCU3jaeXLvvaYfa+W3eoUu
vqKOkgrHnCsKU2upYe6ps8EiWOWFa2Zq5dk5PgJspyfxUnIAzU+9jJQFWjagogBeWSXG4RWyi9tP
MjASJ50Vin1BOKo4zVmVL2dpePplbpID6AUp+yvaja48dAetUkiqC4Tmm258yLWVhFVpBTacfN4J
ZwJWAF7sz5rcwcESrX8GzEWf5f7gauW1JsC3EAnKvAsgCNu76L9HO3ge5cEuzSL/p/y6VJHrfgA5
4tmtQxLPNek0lL22/3SCCL9q5UqniQ3Ur1W4fGUR4Z1Y9UMgBRNRsXQS0txmW5cURof84KAyifyH
iMQ8lM8OpSUFhQ0OmYcFY1jmEpkiv9jlFhCb8lKkfjJznL5uoeebBJnvyrw2uTtm5RVzsg9FqGct
tAAHSZALk6GvsA/LxAaYTxG4zH1dgEcKGzICtc5sw3FdDNW/1xKxw1KflRZLZPwY8ckptVmQt/HS
apiEqjjnPQ5kKSIuQCjmlZKorPkvAxJDoRQGmEasFCiHAqD+X6Ijy+NKWljTxKibv8mAsPiyUww+
sALB9dXqTSsXpcmsoo6bz6SENeQ39qZqgdAop4d9BCJ7HSxzpAQP7XCNh5LEdGH+aV+eIN2ogRDe
KpEFQOSzxbQ8TmlJoOxzG6PM82M9mjpM1G+keG1SSK+jyOlS8Tf0792EnLy7nZ5j/KyQiZ231cW8
XW4PozAvBz/OKm3o70oJU7Y9l557333WyV4ngJJJaWqnEtAwv/ezByHEpcHcbAtAQn0lYoSs8Lq+
TlpzTpAN9Kg+j+bjBEmIUXZLNWgwDL/jH4rZ0eYTuv8VLXkUPKspEg2KKukM3dl2Qn1ehMN3qeSo
jis0OEqXkMKfv+WSNZb3eHF7F30Pdw6iNuHqjxZ+p8HnjsIRdQpexwbRPHEdxhOTG68hTgdV58+S
X9uenGyBcw0uU4o1EgszRy2FiXuh1RXQv91BdO0IdsNIExb9Rigdd1n1RauPUKxpVbQJZSbBxdI8
Kuo0urSqQNahQgLsrp+dWkhTTYRhZqtWMkmAhpTiSiP46JHWiy3c0AVGVFMBX4rF5S22QUNp248z
YpcU03bq4tFAn/Ji9nsnQ7tJKqKIltt0ovVEl0A6Vr8+ZYj3kfI13j6Uv1ti2Yb1bPQqIwVP6d2a
uEudZqe1cbxKIGBRVl6oio7aMISAc9B6wIo70gVQJqMNNUup22VmPmQojI2EjGQjvDb9UMfkegB7
2YKvqVi5GDgkqLBXLIJxp1TNbn3fVVOpcVzQ0DfuXMBYFlWvuSvL4sxaccVm0MMoQkmhvgxStaKa
x9aL9JNmsqVtcqy60uxpm3Q4MS9HO14aFzXN4hztER4ufkI4T2xDbUOkV9m3lgYqCD2dtVNDf0+w
ifMwAskfZB5O5axlTWrVF0djIRGSG3/U6A27m7siOdbhJY0bgVvda2XkhdK0FhfllpdMOzQ8XWS/
WGNs83b5boFeqDnyKgg0Z1vxoiU78x5D9nf9Fne9dj6lIJncziwV7hsH+f/1fpTcNu10QWJ5rn6u
KmLo/t8HHqAGun75H3jr0YKfOemGy8jDpi1YPTiRUo+o3+Mefniekt1a9B4nbr4LvyJlkWuRMKy+
zQVIRKXg/CxwBDD+o50+f7YzaSs/YP5h0ToT0xb6KWoojgyhd3i19LIOg4rE8rv6a95d86kq3SlR
GvRQNct8KVYJc4+O6PBfjBaoeTPB3MIQZ4IkSuPQUm88xM6cZ/yusyhnhUOdCEKhqydly+zUI8yd
TVrTGCLBYbUm0dP+X33sFDaElbjhpD5QJItLfoEr9BDVHhr21mXrWNlz8WhkzlNAxmIwPKpIPrRm
wm0AJVo3nf0Txv/VqqUlOMVmb2F24bSddncwEgMQYQUF6r6MwRh9KnTggLaQMfGIPtiEMUOmL83O
aRLXRgedG/Ndj59OZg/tZ/5xFsX7/DY0pRL34xa4G1yh9HZFiFFZfIc3oS+vTOwaimbw9l4x25il
eCVHa+V7lPGX+1/O7VpR+aTqnBidsh9diEhZgjkh6EI7Z76NqIn0QLzlrBQQlsWp4XuEdPaa06Z6
KuAEtiZ4g0kN9cYAvM4cUNbIa79r7AmtWXoV3XYok88z099NLyOyINlZx08QymO8/l9ZuVxLeO9Z
JSgx5Qw/arJRg/lulGOj8VV+xf7j35iDCxr88a8D1kaFCGOvCWKHJcI0KjGluM3bDnISXws4Z2Tl
ZGsv4NIputX946KWuUg+2L+82BPMc06GWWXC+QkoII9rdAwrsq9+bzul9UHwiGg7ffYNjaVrc9kz
RcNGtCmGTqGRx33fJxRRkGDK+qqJx96m3zJl5bFfUZx4fXaPH717rBiaXpJVyV5/tmNJFbsQqoma
1RLtKnLjnbC5OauW5RIJa5EiQYOobQM+i6NGfwcgAGHEZfu/wGlf/kNzs9/32DPQaf+GTSE8P5od
ATVLpZJA8pbmCaRTKwUIbJOxn4XuGOM7NR3VoMWp1cp+plpRQi+URZpjydQvps976Ypa1eWm2VcZ
iapZr4S1cXiAWVdBM4h0m18NAvbK4TNYP8SQUmwnzE7I5ezeRr7p+s/OemxqglGJ+Sxc8NG025YA
Y5+gPIo42M9+IsT/2XEq2Er3XNSi9Fzd9hlBDObCT03ABFQzikrtB95x1RmfvjBnORS3lTi0yQB9
rvtvDQLfmGjnaYGV8MPD9bqO1pi1m4SE95krCw9dOHq+dZSsrQmeNthBd/SkDDVy70kPgIRizTpO
li7UXvQq+UvH5YcGGkNFPxRtD8ZJVEBgoY+1PCkFaN63WBUzgTrc83xXuMXymoDM0l7YCTleR8Bq
0aVpw7MX+IgOkszuTO+ijW4enOLGyTSzlRK12od3PbXiBVmWETYFG/HRmkedwg2kgTfJPt8AOm3A
/S9SIUgi9tXYGJFN5acjIjjD8Wm6HGya+nyk3OlA1a5n4/8ZiTJOElEX9iGM4MLtruq+OI8mIAqf
h7W97UdzXq9xBGUiA92RB97FqQtnmknlTgioYmQhBFgVyRWP5Sn6TvDMZb6Oahd143/fDYH9t4Hb
saoZg7UG8+tLUl5Nw+ahZz4muBaS/uZr4tFf4taDSjpIVKSEeOkgBptRfTHpbk4r/qIrzzObCAJq
SIZeHX6WMx3W0wjFHOdqFfWXy+BBVuLyaN2KXybHn7iWHn/B2boHdGVYN2C9dqEbyYthmW1VxXrZ
cZnwKTS2HaTZjvop0FjgrNd25iLu8aHsT98C/idgESU39sjlhO7EOu7YbSOv/9M7tG0+WLL+vu7m
vc8A3AyS68sc4OKMes4PmQRqXn/Q869Xi0voCOV7yqBE3L98oaEml0DrTty1/zKj7rF7QWNq77/E
Eqc5XiQBXTxznCIS/AUEMAb/gr2AUqZxYs5+6hdM2U25rMDwr+cacb1CukH0FraHcBCtZW4WWj0e
TE81uKrqAxZnWqYB7+XILZQTyOcl6B0ODM9IggG3B4txiJPyJuxO6PtdIiITPn3Ka+LNEO4lEGQN
EPf2E90EpynhZ4bCFICR+Ti7GbcJmWCwpORDOSBCdfd6zNtNsV1FO7v0yfEZcuT+DUE1jGYhaBrq
WMK+9N9FWFjpEUGxcvl7nMZ0k0CSlX97yfG8glm1K7D3gOE8lOc736+VP1AsrcmLk72kcunyr9/k
U+OXF7SE14WBYAs+Gj4Yt76FMidi+z8RsFSrgxBwgpRnW3KBuQhVUg4TPdyZMciv4yOzxMwn+AXY
B50u/sDsjp1KNW8wa75aDH0sMaOplF6jCvGEIq+vFkGTdjALi7Y7zWcVYpuml1RQ8t1LNNf0RG7t
n65ouD74cuTY6RO1R3qnmRZJVBRrJcmMNHdxTgWY6sMkYoVcT3YxKg8yZxRwMYdy2bM40/fLPrdA
UuiUAkZPooCfyQbtQqWHb2zsnKp2MrQH3EhddyF2nhTgF5ZNSfQ+ydPARn9lg9cp27fDBwnY/9h5
812YFxuSSuurPb2QiGWqwQtKobPs91qRjw7m84vtnJcowP/xnzkS3U2Wh7fKT33Fmj3zPg/LPGFx
uYRpbGwvRnnrnLLgZAJQYL0fdZ0QLuXUZN8I6GuG5hGGCO3uXfglkYY5WLP7E1jdwlK5eu1ykVh6
/+5RvnFxB5L1+rvxVk6O8aARQQTR/HgPnipwGVKlnyzWvdphbDtXNH1uJlO0hRtiDHgNJRVtTiXi
27vX6ibiPKk8ROyIDKeH9taH6UMvp8qovDLFR+F1+j43ijsweJitw4fuwy15oVnZCEgv1oxFfNBF
/uKmhRhtb3KH/qn5TIQfOk+5aRNc/flPFaallqFBtpKAXDHwzL73DOjgFIIctQkiLGZTi4+oLR7b
cHG+s7Ki6TjyzRiJCZipHpaaZEBgteiWPI9iamKnbrX0/Oe7i7tifJuq7HkldlIdEb1DNTi9z9cl
0OwKKiOZ3IQe0iv0Rt4IbRQ0MAYSTY1Hl/weDwkhxMFevG1TLIsSsXDkgsFj910pOfcU9hDMdtYm
ZWpg7qU7oYNNhwJq6y4F9lTcoKyyKOlt/Bsq50QAIqxfAOoa80SmGTZyPEoyMGz1irllSTXz6++y
qGK3nO0lTzWDvlJeiMwdA5ZLQAJB7TaSudr5LyySJOVSuPvO8d3ujAfuFva001epL4ui9bCv6gwN
LXeQsPDZDza6KZF0mMWaYgxWeHh6qX/kgPdwOJIkJsB72U8HvkeDDT7ns7VewHSNn3a79jJ04VVX
AyDrDnmZwWn/eWEoDSHbJzwAptBIWMeL7OMgKLA7KYCmGVxMYtZmKtzFhLiJtdsA7P+fPYNSwERe
60wQYCrCyi3+DPUxFPNzS1TsSdgoT3OUv6X1vMMNn5FSZKLjJe7BPPGj9mbjU6wEK3V2K+UqCUP+
eTtiYB82cf/oVgGycb75Rgjn9v0IIjqE2xvfMMECYwMOWdCVSK2d9kz5S8Y3H+n/hTjPuiV43cgV
nmMlwq7/28ida8AZO2ARiZfZlKX0mvbilfGezx038eqnALzN5DJjg1WlkscWrvADK1DzegKIAttz
VX8j1J7xcrB4Fqcjr2ou8qVL2MeuWcHqNLKDQrqgCvXbALRwj80lQAFNzU4lKqdZ9L/X9kwcnwpF
YWbyj+cJ4JBIcXUcHnCMj9pXwQgYyomEvWex/STtTKLmtk7Gne6xkaYP7iv/LocswDX0EFpJ/8VT
So10DW51tPlFEnfQ9p6+tVFKqPYxNDq35wOH/34Twx5pN2hSfqyc8QrseJn6MODHifMBhZfOn/sb
6FAaVGTkNfG6zlwBrllSHZiNa6LFoKqqkl0ynvarXqDY8udcmeX0h27kA9/op+SNk8tYLXO9Ft7h
50Ytt4UAZXow540VnzLUnpk1+2RMC5eitoyUFfqgjDZeh2ca0rb4ULL/W8yl8vEXNypMIpLIvpGA
wYl5NWsTv6dvRrItkib7j5yGb64KYPtJGJDQJOLDasl7s8dVZOO+DFKQcDsYz3KwDW4oNJrIv6XX
Ra7pi4dCtu0jaNLA4laUAhFK49+D4oh1G654FOB+9weQlIEz8HaQKVtonwRBhhVfNzcsLWVER23Q
cG7yZIwCnRE0Nr0CNe/kxs3P0fHQXQBJL4LBcNzNX5xsTYqPohu/Lpf1ewzEt/krGnbVw75kFM2d
Azs8D/FWlJsxTNJr5ZVetZrKBZDi5uEGkEdvlIFyrv8JMR/6uQlA4Zd5B3aX6XXqk0OwZK9GXoqz
2qN9ESvxTue60Aojl8Lbrk8ciQxsTCsCpHgoZzDB0S7sC0NSJTcPvY9+WXsC5Wk5qW923J3Q5iuC
7ks2CWuaxxff8eBx0xUfnrhYxCYj3agYjm228M9enTIkWZUUb39SONHolPCmNJHaCA5nMH2rw0C8
XjWBuAMPh5c1n3X4W5/KelU6zoBuJ+u8OkqrEk5FxE0h1e9LV4jOBVsrcFGyfYnpXMzgk4HufcU7
nr/3bAVoOIesqeAYlRDQGa8wbcADa4HQPb277uKW61+OtGyShPndqwhebcrEHEBj4G0BLcCxk8wx
/nezyUPLMIRwEUsUVDVI0sFQvPh7p2WRFIxnX6PPWj11VR/DnWkITCzgNSV731hMNIUubbtnYKq/
MUTB2SJcna0aSNFELF3k27QPHVlabomV7hJ1XRTEQcFF/4ial3UdrMq/JuNs/GsubZfrN9N1p/gu
daHOXK6WShF0svFbafAcTeP0gUIpeuGkxU4kCAw1GEI+I45kKNAZxZ+IPSJqS42/jLyOJENlGXx2
HmaoZ0+CmzUP30Pc18Lq4JtASeaxCk+F0ec5PReLafLjk+c/IzzpACClSo5dfP82905bPPH708LA
P+QDXzknRUG320Nb0e+QXxTI/xAzpiTIabLjAdXghyYwjV1r+pLAJElG0yzn+OI10HQv4eXbV9Ul
sBOUmzLCzDMn2RZq4L68lcu0rbUbs3IXjYJXXQS5ur64mCwi39yVqAzutJIPGNWaE4PuYryGyOVp
Ubq5VUMP4fL+YCdW6aJ+J60ktgCDocIq12hmlRAJLkL2V4bPxLTIaERsiFvFDtW0nij5DsU7IOI1
YtugMfDr8+yMDmO0llRWMvrnltUxTtKXLISXGhzpmZFNFe4oVJ4UB9SecLjTqh1kwOPkl+D6E5De
ZRkF/bfIuxBrvto4p3H9eU7mEkooMD5bXuk6dP+rBXxy4oo9WF1J74UupnGnRA1OHn2iSA4pmp8e
SBejM3LYEaWhpbldKzH1mFDPKzsw5zwmRCqguWAK4TZG81FFHdhg3xfRB7gpuha9zMyTo+G6CzkS
2lF++AG1Fe+VdF+vMmuCa/9g3ZTT332TxBl4kw5QwclJA6bMfG1iNtgDLeX1E3wD3Zl78X4caq77
1W5+i7FWvYM7QRrTUIKkvQo2X0jYBd/87xAqJxoBGgHQnceJOfVPJQ68LMCNOQd3PupYspf3xNYU
zR1W13QpJJBI7wt+aErxRyWiKg5QdAFAubEuVQQTfDrHezOejYMoBLHp3ZBC8rAhFERj9cLODyWO
ZEcxRsoN5jrWo0OQQ7BxPK9Hs3N2gXNE3sVnFrWeYJmsZmYjv6kswr1eHpiYFkKqsageIW5TxFo+
NwlvvhakZoYPpS329Et7OeXekYc5QZoJrXUf6mRXr5sZHdQIfm+ngMtmvmLRoqUPMSUvFlFVri7Q
deNgyGjd3oMAukrYP9Lyz55z3faJBwDO0a27HoNkJbrLCa7seQSLRM7McLGK167PX3vp6cLxxkYA
OUp6BuZ9BBDAukWYcxl/YjBpjJMoybSTL7EQwTMMaWN3+CMTo0MD3Tb0ounPJ7JgFdRfnpS9gxdF
V/9PFBUqDiGGCyywTm7U7HT7zmAuFPOS5LdGUA53XhbBNEWc6jbbtDeDuPeWMQwALj9ixlcho1gW
1dFttj6BZFb9+6fq332f89i1ZhG2hrYvD9eOxhoOoH9BIjrGD85EjOlb9mhQnVneBHBpW81MxsvU
RzwUf+ROXCNZ8QisaHcZCHgNO2YaYJRXrUcULqMRMBueA89i9BLr+kjp+j75MTgj7oQXvMuZUbOh
zCaj27vc9FOqKKozbfHX/GykHCBnzlG5F79M7HbFHwU6ke2z3mtjCaTRlitzLsEhVM9COuNTkviE
Sgmx1I/VtC7gOetVYxyk1HcZG+ag89Zu7JW/IwIAaXoqdkgf4On2LTZwa9tFN+My9lfV8ynQocDT
1wSwwBD+fYrX4jS0u7RaqyTgVTwuDsyuYv9S904bLAcWU3hNyE3gGjPHeiEoEyn61HTpFlw9KZXZ
vKhvHyevsq12ElM1uhmOLgPyl66zjCFo3MDzM8UoIqQ33G+prUbV0Ieg3DzTex3OUlBGuvh4HrP7
wK0j670lN/5tCnB1SX9naSuJctibRLXrz/PirrHuxretYngNcY2va1xfwONQ0c0+qFYyGpN6e4XR
bIxR3hMauQOP3tJXA2Tnl6ptup6BfT0cKm34iZCuLYn41T6OxhzgKBWgpLAgM1DjvfM14iiwxJtq
eAjQR0UXXvOx71DnCiXcaYjdtJzxVpRZDSfiF9VlT66OwAybeK1dwOy9tAepylKbnu0/Yfnlo/wo
I6wII8w/j9Tz2LLJB/FyEIwhdy7EJlgpusot4xe5nuu2tXf7/hVHf6WK7aMK1Kd+5JUiNUUwhVhg
ShfdJ0kcgo2WeSgWomnUV+ulE/hmMttwbZFcIZla9J+opuZTXEygUMvLAWzHFgfTIi8WEcS+C5If
wfj+KQDdEGC9Dcn5RL1RK5bfZ3yUgc3Q2ljeI7npxQfgPb2dCXS4C8W3m4Lnlad4IUY3Haokz4lh
3sOLE2u9nUOC62sk6zwD7Je7NC5tbu7/4NCbKROO5zeyZxFe/nKkR2ByNTJC1bJqQ42CcT8VspBS
nqh1qQb/WuR3G+CDDepSVFAbHCZYio0LOSqDCiKlzNnVMy8gN4OVmV87+C7+LGTezUADD67egrhf
3qDWD9FTux/qg98zjK1dGNYMyRs0n5THz+hKWOfB9zV45Lobc2uuNESm1SuXTl0lizkFdmkRXPJY
Qq4eqsEVfY3V+W1zmvUlrPJxyHjX8YibxkZphqEQOiEPrFSVOLR0Hzpt1P8TdXO6FMR27MaOTLrJ
xicS3pCfdmapxKFWjFD+LcfM4M6vlXtW9qwLeikWNVaGbETx7ZYpiyE/nDGvw6ksPiBewvTJDJfQ
U88iFd8p67+i/KsDa6Pd1DWalHTY9rNw4JauXT/uHrL/XY9wsPAOblvCaaF+Ll9s+4fNo5MDgE2n
EKUIFAPJEr32V3Mue7+xTzwylsvRnyG04lhGJ6CDt8ZxEIz5uBzK+pdFxPOFO8AoXp/7VEVh4sKJ
R5yJJ/Vfc6/Uyu2YmCU3y6TWZ0X9eiunuSddr1aHv+liKRanmlj41ZPxqJigTWk/gB26IUaCxo7B
c59WFaayXXDGzG7qNgcHaA632fdFmhRewWl56QGGUc0gSYrgTsH9cIvSWNSK0GTd2nhuRBdw8tft
S87XrKs6H1phpV0IKJarKXTanhhsV7LgK38REgNDePXHO42FcOXa7YM+A4e4bdo29VBAqruB+uGm
QQRfLq8O1tHsruP3j7tZY0kGWIQG81aHosIeHVjpW4o0bgDHJlOFOrZZcvbGeUFebnl2J/WdxkXo
35gTCjGUuERXnp/7CqOW8O7Ii/F2Sw7tfEqU4F3iwpBe1hp+V3ppiJ5Qcq3Sf+RMyFPIAC2n47YW
JuWjSZDZ6XVwKRdhngJaHfPwPHTXUduvluHwJ9HJNNKUBsxwSx0rpoPqDKFRqtkOiMjI96k1YOOL
XhG8iZWws286ixkEwTjhclxAgzr8V4VcKwp3tEhjXE8R2zUOvdAmoqlftO/U1LLE8KwcgYmQqqzN
lDp4vyVbuErQxmFvIQ8n2bw880IX0yMP8V7WkgEomntepTUoqzXab1qlWOyWvM7+3Y/owkhxAUyS
R3Ed+aCsN3aSa5KdyCzrM1zaGWKjpm7Ky6+50DjIBefyxIhxGVjecYJzKsINQqbkLcuHmvr9908g
sYfKoBmJIP/TG2bMKHXvdt3u2zLwU7XCVvjxNdcL854zmAV37/4+iVDldOJ93LEbFwtAwhf3bIUe
wpYa26h5HbgVVF0XYYylkZ92sCwCEX8gFPtG+ifyFn6KxX662jVxGUfsUnDCuee7nMfw+GCmAVVH
IZNgLciXQkbrq+08UjlYAHTrkqpQBw6IyVMT2TfDbutpbIUkpvkxG0C7W+sbbvBGPBn1W26jcqC1
ggHu4iyiV9a5yWoWj5mq/XCdPuyW6KuQohoF0SFMJVB6qHNS1kC672Lu3B4eBapnFERaf0OV4dzk
ShJPDeWGAm1kRkQW9qxhJONc5ZRfiKjUobwr8lQ4Q8/MU3jQ+W7rjiP5FN3ofl53pW4X+ddoVO7e
NQQ9AUdZ0iqXEmOFmIQczAmlZy4yJK3vWpnPzZrjtsYDLYV98Cay5kCIOKpkO+zLjsv7/qgW8UJg
9p88Y8+/chlA6Gf7DUIjhxqsFe/TsfvCD7Fkif8NK7zjTj9qwMBM4EN4BkOoO9RtpeVJvJXp6Qma
Tb4lCrzsv7Ac8SKcFSU6kTx2UQGZeCNxLvv+jFsF0nCrPuYvdwqlv+VIGn78HuCCQKeKpZbhGJJk
6KqR02KdGGkOsOLhiCDR3H0ThMa8xNmpw9lUiXyUvL48a78qDa249OEmTPrutMuz+BbaGg3ObsL/
8u6bLQc1OEDVnrUsJrBNyJ+0zopsbjJvqlyfgBY1Sy+n0JUrQmD3FWX19o84O9yz0WTQfeiYtRh3
Q+NwX8C8BcJBp8WvUWpO0uJF4Naw7NdAzaT6LAdJaFw2Bkw2Ml79AVU6qYl7SMcaQ1c2+PIZn49n
1p5sF0goydfvJUwtK0LEivJxtFxBZo/xi077z5aY9xoc2Kze+YNzVDnOxfSNvUqZ+Vt3LnMGQMio
GWIUYZI6AGeM9vDLMkMXRt1EYcsPxkBiQqbjlMXBSWQJn1CPGCLd3Wep04AHwAVHBFRyic+aUY++
QzFE7hoRUdk/hSGUVko1D0I3kA5jHZGAXneMVbSe7gd5J6rgWjBqWcxFoUQJOkaf1klGDbPd6j88
InG4XR+XXcVPHG/5xBOsUPaXapj/uwxQvPHcDdphYHpwWfisNUdXSjzgxd+FMpirZo7VXvHaXL1t
YMv1tK2MWSed0IHt0dTfOcIL58U5OZBmcXZvTR8dlCKAb9CSHGv+det58fJUBLcDJvBE+6nKmwDK
DQTFmGcb9B7tI++JhRFS+zTu1wEq9VtM5ajGVz2XQzxvvtIlhUiqI5pWG1h+3kvRDFxfcIaMTg08
lIK+eix8m1zJMhxvD/CakB8ccjUEJ2qzgHjgy852Orb/0K9h4tJjUQf1QXy0Mw0b+VYeA8Bpl5pI
R9YNkEHtIfv19sVkeVgWCFG+QQN/c1BVEsrTeQvV8L4uHPAvj9rja5W9L6kdxCOkYWROB3KhznmY
78mTgOXXm7UodJkIoeUxgMnsjPM3YW5RPZoJWpUD/tTiOcvmvE7tziwuzloqzDnJnAvfW80rXQ8s
3dxnOU3gZdRpg2B8KUwt71+FqFkECZAraIs82u/pEGC9ou2ngxG2yaHE/HQoJHbZLtspT1QCxk3u
2GMlCpluWwwf56S5OD2mlhrhJJo9qofdwkXuvDh44qoCbHcm7coMARvUM/YBwm8lAWQr0uXe5vko
r+99XOL1C0D0gHfaj01808QCpWFXJ5EjVYZcvFsr8QOP7x0yZBbeYg3SX0f02l7EMq4bROScJ2Lx
Ozkj3mOLD76PvNBsHbFvsMgmSPUCWkFHCJ0mJ1EaNfWX4yGoSPwwa/6OynrRm9rHI2Hq5cR4eWV5
ulnsb8keM5OQP1BsOusPt4lpQSagGUYn6yHDiKe62CNx7+J9J1paoteZ2vwvH2V1PXQDde9MD/mJ
Wuciu3FoLvfPf9ySKzbaqJGSIzICG+2MpLICKB/NM5shcMENQLdzT4vYgDBuH10dJM4BZ6abz0IT
UgF80MARCT4v/O/mUbVqBgP0Eck42k8VdKzt7yiAWr8tub4R5CBIhyDwj4BTP8FX3EqB8Y+RLq4W
ROx51EAT2ssFJeJ7EZGPSs7A+rtfq8rBbUwjj0bRKIE1LR0+WkIXU3eZl0AepGf1e1fbyADAfdFr
Xvja8rsiilTc+ARa2cZNHTt+oexp4j3NqsWR+c/prFrcLcuZe9b1JaC87HCEMhgiLKxnocJuVss3
6wXX4KMd8UDT72mxYqDjg33keQqoRWRL8MahferRZ/ACWWjVInYYcS/Tor6/AUkTYdZRha6Fmf87
qAkQ/vbtMKzzhQ6XmtgsJZhxQp35F6AO5MwtdKUDHli2jwZYVWlGqXadJlHmxH+kL7Av+X9q+Yot
qKFjOeWYDUc67RbKCfmkoPxjBMKtskLFIM1iGBbtLeRnv9A7YHVcPv/rTOVTwmynuE2v1ejhG7on
qgkwnHR6APCo2t9hmREgivu0mm1uC4m4UVZ8J8ZLdJnx/37DcSHqFtIoxxCmt/t7iy+WVKe9wYZf
24jXsIXq9kPeWzfNhX1EbcjrXFrnVA81z1w6nyGf26ZSF4V2tlR6lDgLVp8UqrtCbxbZkCUHQBpJ
C7iFJW/VkjBErvmZTxh5lVf+/0hLMsV0TgBbE/KUv5SjQA2uDpReqOuyloZWZAZT/dSr2TT/Ffz+
RR2IpDGE2ljdYEYfxhLrRqv2yycT9iKTfTmm6goQySrHoazzUF5ZMlImdOxrOkRz0T0/tAkFDSmt
78/mVikzyLFrMUSlIf61WYgOwMS2+JnxHJmfhnp0l83+FkaIQPbQKMx/yWExh418NmgaqWPjour8
bvhiHzNyQXJyGLK9jbvt+ZQ+IQPMjA7L76f6VDD80korWDb2FwnxviN6gM8pVriEXB7Y3cEkrQ3L
h8lIABAxSHp6aE9yYXrHyUCl6OGcNKbUNkvsQqFxun8azXEOFXp8uMHbA4sA29WY+sDxzY1s9zRa
IOcqzap59synDr9s1fFRd6zr1Ymnagl5o66idl49h7PEtmd47qhSMrvP5vVfs59norAFmGOUSBI7
LJSPK7pRxyMRzK4HscpJmODs1+2mdUGrkbC4g4tdjlGnpAiy6f/lrz7TO2BSQN7vpFbqttsWWek7
3qLS1fLn4kqPTrjgfC65eFkV6AMb4Foj4RjwGGPHSmg3d4gLpNVmJO3pRFaBxx79nH1uPvZYo9Sn
6CBGGBY31ozMB/xCNvsaK5auUklAGta2HttOZ7ck3vI0VzSM5zyawaVp8aiIyAWZTwRXv8VBA2vm
WZ+7pQeGw8bViBiDGwE93UoW8VquHntTJZnTiFPmkwX9MTeoRALsxed+/EiEJqTq6zxYQ+FBn7L+
s0KcrhnmFrsBTDQFu2y+WMVOAr7dMG/tLfUeL4gDYZmkcOtBgAjWxBV3jMIxCmRkLbCffOepv9tA
PabXbArkH0yDfZV/t4WYGFqUlxoRacmZFz8MFmTB8aMIT4eMbl+z46krO9bUBWRHG0O43UBYGq22
59EFfqn0C7EW92Kp2ahGZ+fRwB2gRg2HdeZo9OIbvFzPpARi8W+FF7E8WcFvDLLgV0QGpXxmDQAM
UR0IkqEjYRr62cknozpyBnvRQfiQFDwzS20JD5oS5fyEDya8fcXI/Od+pMMeURhpYw8KDWMfa/Tz
UihFQNLrgjqLjj7Se4PRbVDFmHgApQOwJQCS+QENrBROntEWUXBkVgFYYFZVekxdDaeMgmW6mL13
0iDSGEfZ1EWGwvyWxiSNwwQZ+TGm4LbCfs+8lgE8HFzbzNuQzr23qkh/eMJErPZyL8SF5lK3cTk2
SxLePPXpcygOICw12B0Ryyqv2/6wVrW2O9DftxqIyKRd9TzN63gVM3/wcAeMBP4UV+zboM6DrxVz
HMsVIPBIgWK3B95Fiv1JyC0RCVO6J1azslK2GW9BE4qBouBq/BcrLzR2tCsTG7xNNoSup0QrOJJ3
WEj2Dl730TNtaSskaLWjqU/9BLU05f4JLexw+AXUxgOPFoP4ndHh0mIBgirFeY9K3xetOQ8ZjF4h
3vG3kKCOIcqWNf52QKZS2aa2+AW6gKKax9frVkN4GSX2uhx0CH5iMfvLKYiisZYsk4YgHRMrXoum
5qRoabDeswJHCJnjoyPbyyX4tsOeWURYRkYsIs8d+0MjnGZYa54fyuAO+LRVmjW5T8Jaokkp0gse
o3gAfBp6djKhrgGrds1oGq1CxqRdsU4tLH+Nz/RVZ8r3LaB8Dibizl1iyZCYOVMqF4iZ07WvdIbW
5y3SjPGz4ePXFnUOZEG4UjEzDRBXQFUlRjL3p566HJ4EjWawMUxazP5mTrp7Z+7OGB2KnM+i4oGN
pEyt2g3KulExAIWelvROSMlxIoFFgU1KbHnw58tp01ZQuRHzaJitIghsOsHBlgH6IWf4jcigP59o
o42a3l9mY4RQ4hVekH0ngmEq/0OHvafa7tzLuxA/CXov7zCbfHL0/cUwvGm9BYHM3N5KSnxLgC9O
KhYTQ4mhlLitUcetCE+XtqfP6amtk8PmkTxJIFHUoLVT3Q030mVvrPr1Oc/yePpLExbRQKzhqxR/
pCAuRyULi7KCNpdOZLfORj55mJzVGC0RsLJn3S4aiPaogvVVN6/S++F8QrSIBvEvNDgPl1PDs6Dd
csp5VZkH66Nt2L/jXGZdWB0UwgPBx5r+aPPbaNseBYHFgXiVqijRjaNgl9EzEfPu72uKDa8MC6Ps
U4VYimSVE2ivwevXERvx0WRp6iXoQaxJDjOD8ngUAz+qmm2fnvtB0OY6cn9yBNjEyqIjr4c+3lrq
NdeL1oMpp1wosNLTUTKSqftK17fUdKbI7yHTwhczhAE7BV7Fp7QptdypbK0k71FUnYwi4/5i/Gdj
UngkAQTS+rCDtCLKzA/Sw/YBFVXS0iSJq2FG1zR1XjvCZ38MHSnTPnH56vYE6dBb7F4rAm0eJwxq
RYZgsx9cCmcydn0yrj4g7488gzyxgnZk7mU41mjdkJB//uc2vphZrtziBee2sZ0b65+RN8ewF1oa
fg8HDF5PJ2lDYYnux56yy6RFgm+/JdEISN6u7GNAZoe2dOL4hiWHBTds0OFwZwpVWZeu+nTuwHUf
Phje2wFvvhNkaIZ3Qr61kDPE22BI8ae3ENbHoE00o7ZrjbuBRHxnzhWc7UFRzRZhOGMeEvspbYi6
4jQNvDFZJ7wond7Cz+FdYDbu/V4SIVrHH8jrI72AkHVB881s0dzeBQReuyleazLex3d+yLfHzhwy
Xgylj0adObLWM7MKPO1XcVU2ydUovEGTzsr4g+2pbvuKzTQtYz5l5M3j+JQmEMsKcYd21Hc/o2Ye
+WF8KYo/615NBVQ0au5SNnYD/9uJZreCow9OK74Nys1WyNBBbNoSwoW5ILtMfDznhr4ZjZOIbOqj
tEH4+21qAeQ4dVjBfk1Zdpu/48xk1Z7Gj2yUBTNpbaRtdQUlXqnb/h4P7uB0DiFftiQtww1cGTOz
+mHlF68K7Owr1qAX02Yr4YyBxH1OExxnNM/OUNC8+bA6Le6n/oIovw5FXuMA5i8x+p3qdeBElqay
wlhIWZ79CFbjhQnIRnVDoa/cZFR2jEVDrk4kkH3JAsMhkw2kxjKditFPthLu+5L1zrKIz4amBGsN
9/g+ORBWf6uN9OpQ9vo83MFx9sBImDh+z/HHTi+LgK471C24ugZO87kZylLxAfTAuq8JuwPmObZn
7MhZpRW753ERLZFFJ/FE6WVE5W0hcUQO618N2z2+SknpZKlwPsgkd5UFWTx89bwto5+3fYn0Ryxz
ufb+G8mXRJffSZkdr7+hSPmNcf8kxIJhl6qj+Sfh76VAozRaC/u03BZhGzPpsoyODkfKGTvm4Z73
/hGkyYEwk7r3jZWC5rpkN5AwyylRaknkZxG6aIJ44dEmTHeOURV2Ug6eY+V/ef1VRGk9pt/QM48W
IG8ie/QwUJcvv7i/aDEBFR/k3qSWANG0JMX3k3Vw7f+KAMATKMjOymslu8XNzR3ArCaP/BO7Duvg
LfhVPB00D5IXt74mhxJBesWkv38jRobagiwFeh+2heDIXdgEs+kDvd0PquDxIh+m5B9hDxtKTSju
aU1Ki0FpCl1tRSG4bjwGa6NPzb7tGvSBjTjQxVdJkhWMcoD0Hs1jio1GaE2iu+os2fyYpA1zbjne
/IxnCinfWiBbwD7J3zPHq4UgrpGnCW/+33wDQWZdtvaSIuy479tqNARJewc2v/GV0MGzkhHDF5QO
hE173KGWXFfwFCdCsuBBlc/Zy0QwFsaPviyHRN00ISWjMfAVEGCq3oiVnSQEmOeqdXVHh9dDrDZs
O00RdH0Xhzp2nePlrtDVC+6hN92Xt52f8cSRaYJ3agX/cWWm9VDGDSTwwaZT8f9bDb+bR694K5iy
x3eUB3HPUIzPXAgKFwRWCD2f207AYSBTv3OImsKNhZL2HdiXewQTfYdySXmFHWECxbkRbBzO/+It
EFVJO5EJbymzHzLJcV2yV2VF92Ms3e1IS7UkA19IEu908Rkb8ZEUmPeunBlMi9t+1SNyP7C5wyiH
QFcMpIbLgBycuck3IsWQcLPIDRstmfFkBepY8KSl2PVTZk9pt03bg/meMyuHPVERGN3ZHUTOpKqU
/tJtcADc4MAuHKVHt6/sxOI3fJqEG2kxuwIRNKsQSx72o/utdsi1hm8rPkAZiVLZKdMRpdMJcGRp
jrfj/quakv/o1yTZBcGQS0DgNbrztUCouwjWatNm25tpA8dPFL9Xc/MDLdBfW793H5u7qODS8yKb
XLOr8qnJbOaayJLRR7xny9/4pgMWDm6Jwo5FgLHOeIynqy8iRMdnszrBiql9157pBrrM2Czu5LCl
rXQMETXinpKjWtfdiJZpBL/8xpFQabXTcc9YOsexx0DK+V6ilVL6QSJHgKjLUcHKsIN+MQ4Sj+gF
SkLhQDYBHTfBakRgnw25zqnd8lXk7cYoqMAK7W9keB+oulJ3FJiruFdOAdAGLvoUctn/wZyGrh1d
rHjDOms624WFfVTGeoci+5c9+ZaGaQ68KfW44VYBveMSK8HPhaHnNcOf3r5iqbYC57LqWt3AJoZl
h3WtLpxMKn86UYiCnBlTav3kgLAfvhDmKGHWZ1G/QOQG+XqzMBJFs28MZBKX1m2bjcP4hn063QaB
bnTwrCQ1RfYh3GQL1zy6natB/JlGVhdQIxBd0E/ikTK9q3GZY4/285fa+uwaw6kfiiLuhh71LMJo
gcvXftyV9LL1wkpOK4QHGh20/kCRzjHls3wYwAgjsJQfu9+71+RvrE0mV051b0GcBBgT+9JWJItn
ux+yvgMG8YBwqf95YtyTqkeLBCFVYrqcVheBYMDyBAl9YqTRDNu9wd4JF1DWxZOJTIH0aA1fJb1H
Od44U173R2eDp1jC90AuGarJcfjtZC6XD0aapwXl9423r6KWd2BswZrSf60MPowKMh4m61DRmtoZ
JZ52S1t9S1hByv8WLxYxvGqAbOGY+q1d1Ny42LnBAaK6TrUyotDosJbmBj8TV76VikpaR2ZbD1sN
Z5Rt+9+mI7YYhykCUEQRZsDPjX1FLuxI+6DRHnTbx058QZ5XIfdpLxYjIw0k1jKcPH6zvGRYGoaR
z/tGqO6q6t625FW3AvdJ2uauEFNFiruCnMk3R2CulI75bMKsc153YfAPAY6YK6Dtj+5NuuooJ//8
LLFCtQ3Gqiyp0MX9MkkuimwAS9ql6Ps68h1tbfESGlfH4WHX+65xGovHd2FwINZNqd3NUMtxNJoS
d3sbhNwtbdzSLlm1kLhdZTOLimo8oSmojZxf7WCQyOa1mb+9YrkF1yrv9xDgBc8uQKAIyrhW7T5i
o+nSInSxCIL4BExj+nNgbatR3DrbCqzO15/1i8AQfYWlTGVNyksLZvCBSARUIBECOinR7v7R4Zka
paHT0m1ZeFIHb8pgZO9pvHae8Fd7E4wPPYmt5eGeKPS883BpzA+Am2L9EGufRWLK2ylPpKLRK9hB
CzyV2Rc0tstOAbGm7EBTPk/N7XSZDzTY3NDw+NbzfiLpO+GT+WkXLWggSq/Ht49nN+HnEqx/5ieq
f/R9ircz+dCQ7V7QmoizzOqvnZLi8B+KljJmgtobwFsZcerRMK0vYQvjBsY6DiLtTPoTnd1FF0/W
hWXVgfv299b9Z86AcoaXXHx0nZzi/IY43QsEbcYPjI8cLjmKScofFtH1uh/K0Y3GEjaSWHJlBIZA
6D/jnN6V3sbgWfcN15mU3n2SarZZBEQWjHTApryEjrxQHeObvnQByhkuhuMMzNTIZTj7k5P1wtwD
Ri6iu05G+RMZzUA6klmX/aHeGzJbzccGtRu/7KHGylDa4vNWi4ImLihGbnnuJiJetzUb5nB5cH8O
lX+UpBd9uWNbnAZaUmbtW/VyGcrtPZoVgVP2gwbTgMeGXINXV0mfUkrKGarHpXFSuTmX9fr8Raix
/NTGzEDhv4P8Qmkye2/0QSpv6OP8QFwSt5e6NbCE3HGZTaBKoM84hMm9OX17z/K7acqTDwxuhjfV
dxaqRY/HcRX/eNEsmmcQ8KtwfN3sQf4zvMc+cbmGZSvbfvWh5SE0sV3GVH/J6nbK9V5U7yoMrdjW
4K/GTr+AsKciQ8EAOeWLv7vPW2wUJnmqaEe4eWY/Wrgai1XbEZoMvJUVf5uKo1p1Tyn01t9Ub+aN
mj/MPlTT/a+Es4mmlygohUejJn5otpaCmgHdQvlyQpK7TOUQan8haCCvLFnW9f0pZj/mSE/OjT5F
uD3eNKshbBCy5c9ZKmWVxqZpx6QfaOrcbYDyjFEpdrLEgdXeChZp65OaVvVYWJF61sCg1wZGUcLR
4z6Qfq96skdkyhmGszXM/JsTyud7oRzgA8Im0dJ7ioZKsAnRErLDG0zPXYvdeBMEOvenxrciC+ke
rR9HmwjNY7w/8nub2DDGMfaihvo4fCLkeI50izG+4cZKQe9U7q1kaFFRxVFGEvQY0KR5MJLEBcbv
1P1KrqLghn/+pCDlNtMSMSuR/PQvtpUZC9FLdlGadDhxrsYhE5ji6A/ymHarsrJPLDT/B2h9FRP5
lN84Egn2QhOtwdnEjS0OHH0pml9Rm+hQxq6NWU9pyoXOxlLXLzcEwyV4jfWXdUUKEkuWOJag3VRH
tQqMTXsrmrkjDZJpZRkuwgspVHRN5ZL57JDvre1/3cZfE5ivjbcZh4soXQ8vTu+wGNXvGgefjD33
aOLf3mBETyv4eO+OKo75EKSSb1KpIUELDEiA8y867uJPuvI8G85GPO/2J+sVIzsxs+rj+FG0l8dJ
y/U2+m/CupLduQJvl3W6Hd+IlCu7xdy1sm1zPIjxz+Iuyq0dJ1cC96G2iVGS2XJp9e3X2+ASKzBm
MLyu8ZSsPbRQazDVfIXUvpHaGs/vzLMZG0Q20Q4y5QnnBFgz6zwlSaRQXncnbMG1pKSPM8nSsNz7
fKi/TyGldTXRN9lxa/l5Lc6jFbBvXX6f0oTd9CBzJrZixE2AkIwbfTRHep2jcN3HchJgY94PBLcP
qnkXQT8QH1c86qOijHj2e0VabChi4MobGXwzIwhCZa/JhC4hRjqrTcDiewKk9r11QX/DYWTSS8IA
uglLB6yJD6WgONGPYGxOLwEX5o66cy+gkTCFCgKnMaKGQNY5BR1+SXJKQlfWvdhxPCy/Fmc10uwv
h5Me3Xa7/yb5x2Q/bVyohLg4/UvdDOLkPpENslqmlbWsi81PUnV8vDNobtcoHI4DSQ1GnSgYQedH
ZZZA3dljmcHcvi40heYEhkXq2nrET3dnS638FcQbgkAv+k97AGX94+pUE116V5FGq0fDbV+efEF5
3Mz5AqYAu9KCUVLg5oqg9828tCRn7lI2Cg3oulNw9n5OiUpB37yHpULoKjVpNvDyn9mvgRMsyP/k
Rx3a1A5piCfwxM2TNi2TTJkzPhtKD6j1QEkGv61byxrARSDSpA9RfwQvTdz74HYfjy4XNT86/7dO
bdSwJoT70e4Ji0z7P+qevOKb/G4nSMdO7FA3+rhmQlXGuG2hqbd81W0RtRtuiH3rjCA0R9K4qlU6
nRM8Xl/HiNFGJyofaaGoak2i5ApXzDvsVO6vvNQ3E8yVnvl1WqPg5SLUwho8LozUX2aooclQslWT
ciOnOJ8UtDGWlLgMKT4WT4JXz6tGzwwnZxPuOaHJR4z3d/RGOAvCuymuFmtMDoRYXqu6ZMcIueYs
urS9Emovf9R8OuqK6l2mSncxACscDhMNMoitXnZpFnrRCe/adL9V0xexFwgYm8ValPNlWw6n1evd
xM+3swDwFnY2m5+1KAxUXwKzFrzoG7Da4xzW++C3oHUedF+Jiom1IOU5eqCp0oL8+daax3D8eCtU
HB7J1G8g5jZjSkTgXZSaDQf7ih0B5ZfkNs60JmZ61QVGBDFTlyVTNPpUJKeufEUho/+ivBwGLWiM
bExoeugs7UtKxrLwvWK6JmIZkkmfP7j3xX4ghOOmydAoOMKQrDOb4ZRR5r2kHErFKt7CHkeEB3H3
Fg4+jKLhhBa3PfMoUQ/3I1W6iljdBh08LkBYL40VLr5QiMp7mtVyOSAh3V7ao57KjAYsOnVEBrB6
pfzod2PJNrxbBhbV3V8ysBdC0cIYL6GuRmR1qd7CgFt+Hhv4f2H5UfNu+sA5rJ1572DVCgUHujxL
gj0AMZiCxzMdp3SWhP9D8svBnoSMptP4r723z15khE4F420+cD96xDJ91cPl4aT0FCxFPkKoGDWO
Wiww7QVCzXNSGSrpTOgkF5O0CsJz/164OaMQGN5MCQtqWxJ1mMxgp1qAl68L0rSEGXLzdVw8reuy
KwKitW896P0NDjsBFpCEzrGbO2Jm/MLW/9uLTXFOemwk9O9B9L/sC0UVm8hxGYBmu6FVo1TsCOv3
f9JEYEkOdupX1cEYVcjwrHl0BDF+t99eDJOyHR6KVphtIJMWkD0HN4+oFzREfnMpAD7cHhPInlYX
E9y+0jRfWSAwxaZUjEOsdYrtrguM9Io0Siw2DvrRPHcDPijTWsU547wVHMngsR2CZih3SHqtMwik
C4RFjN9RYqrvuoAJT+SZEUwLdsuK+eRoKNqWbO/f4709aFPyz89hhVyKHdJEc+eL1jJ2UchdJlqb
Cdoirj6JQemhW/SJQ/aq1CXo6cVejKcVRayIo/2o7toejRWtDsVMwn2rKHKz77sTDEW5o2njq2wm
OnMAb99P7LOc8AqydbDFasG1hmxx/9SCX52wZ/Bt4G3Laj+gg5vB/19zGouUnjOhKqO/8Qgh/yvb
smTAY++TNCeTlkCBU6vIDZjk5pqB9LhbPzFjm3AqCO9n2FZ1fj+A+j4yEw5aGHTyc9Himhmwh1+l
5Ir4tPuBmPC2fuqWWYUoDzLELTn2fTZSO8DgaoOApStNj+S+OHprmLf6dDCyd4FswJ9dGPe2CfFE
yQO+Luvhv4/wxfe77QStSv73m2HLQ9NqdeVhija3ISZtByCbPEExO5+1wZBkRsymaUsfz3CCsN0s
rQw03ZQW2nlbSLudW002WSgBJUnGbxX2jv3IOqEfFlwRLqn4odUrM440OuzLII9VOi4S7LlftEhi
HzD37qnUPE8PxUFOHXprYSaWGJKiiR9V3PxZyfFIpX/hlRFuv7ZSdclf9YGGE3koz4s1wrqWeVRY
GY5UmVWyvRI7Ejc2kEaFALJ7G/+y0OGfhZjskoZS/YGl1jc1Dx0fwNTP06W+i6moGXlCce4k/oYp
vP7I+4u8CKITUVaoaJFQTc1bAvu72vpU8SdoJyqjFVQrFXKRmImI28Iq8VgI7iRqCEgebtjvaziR
4BuqQXatyewYUEvqiA+GvRQGijHFLLhKTuwAzSotXm9243Pux2+Vwm+w2JsAtpYy9OHIqT1zBkWa
nuEqqbD+DOoPD7skqGt/tOq2PTGFNa9Mfek2lPTs4Ih5Q2Y4OYlNddFMCU8Ec9Y2bX9qky8vfljM
94wScmUnSA7l4foi6zUs6HtiT72VRUI8p4Gqv4gfjLXx46hxuXDOjOs4S2/nrm69MtOSj5OuwQVf
qBhCiPjQfjDNBWNCuBGs2H87wq+ceUvjA6qHBWGQUUWdtcpH2INWW97nV9wOh4XW2lIbVi1JKuP5
Ww+Jj127HB07Nd/sZob7o/dP4kpuP8OqIuC9DOgNmKPIfLH08l9HEigfYlSWz7rCWqdcl118+HLV
rR8IFYk5bsVAyKNUD7K6OWxpwLD4apqd+X/iMbQy3KOFsLFuCEIE8KeXUrlh9cAwdLd63f9q+/eH
R67kGZZZLUg+nTz75429RPZxii1dTC83fk76sJRirFTqjGDV6dU8wo5MAWerobYKKLL3YLaDjtag
nUzckBCuCgnD1/cpJq9dAz9hRyapmMvz5u6pH82jbIWLiQnRN8a8nZ+yUgQP5kTlbNKdYTwgmgzZ
RxWyWSUFgp10X3grLqKwtbfD6mzSFJ9msKgwswlL1nCp9Vk+wsaV7wlFhp6nWlrjTQB5meJKNpH5
1RwayNTae03QUIusnE6SmZS4FipTSFn6kFcB8GHd4M0agAvGOTN9Ii+lnITXH99MILa7Qjh7dxor
SKMNCwHz8Dh3IzaR3YaneeRic2eg9k8DSi4njGCE7PjdC4Q94H83x/eQZU1YjNhfho06wiQFc6RJ
KaDh6gLgsATo4mYXUEcOGaAPXACc1f0E3oaYmucFVDGVL3ODyaTVZwWqMvkWOr1eh9X+6UrDQ8pE
Gp4cHa95qZKh5HiWXlhmGkTndiu0FrroVUgoLt1B39C4w1c4ODUzq+GV7mkh9gsAfsgrP5q9Fdv3
2vY26qvedJ+O6fyc/UPR9P7GiD/k7DwSgP5eTo1dCS/MiRkYfUAGON6oBU9WDaK8lg6c23CSGYB1
+5h5qgGZYzfOVYo+oOGi5nN1qTalMARKJCl3vqMAfMAIqPyQ8aj74424RODBP78p+TzlasqQpS6b
bxjvesBpKZrYRxO5IrGl608SEwO4SooYh0NujDuneQGxpslcfDi6wprfUSvbqMgpL6AVf45Fr02m
sV1XcmTQVHFC7YSvVJWV2NM6qh1nK+SgltENDRlA9bnXfZsR65e/G4T5tImfJA4M28iAAUDfETbM
j96/1TkcZamtCAWMWiLF+uKx9Sf9QUy0lDNilzII4evcNE0gtcKR+YuHKTIOhgOiDA+bAuLWPbOu
lhjj9FJjCss9puIsk/ydInVmRH3tJiNmcgdovJwRj+MdQ2QN/uOi4W3RdbEFTuWTfDhx0yeN2X0n
JWS1+SY9L19BCer0rHzOtqbHeiSsjYWnNEizzDs2zu1BEQX8lw4kW1tnVQVSd9Tm0KNzpUHYhkHQ
mJpo/0LW0SXmKx0ocswuZq59mu71wP/fCo9taUIGEU9z+RKypiuLrJvQVQcORWAoOjwbZyfyliK6
fNHuMA8dLSmExCiE1nnYwYrMpzPkcPvaqAx43DFOi340Gb3qLjZU4B+V+mbFWn0nOZD3fSoUlRAH
DdXLkXOYKQQ9ZdmERa8jGTrcQ6VzJ06/OvsdwJqYysk3Pu9yoYKArKq01fB/rHpcYs3YSEHQZr2D
JuGAMOgO05+2+uatCMtpigX/rUjH6U2JK96FIlgMkL6P5nMmfwchR5frdysrpHw5VOspKejRR2qu
E/tZmyQXYeFLcGsUe/pkc5/f6EGZrsvOx+DOhFdoSOWqm/eaqZB7D/TSSM8ZmzTuuqQE4ibAyDa3
97i7IsoSaLvvYr1O5tA1zU6l+Vm/4Qdt69b/5yW9Coaf3XRvgxVhbbQNFN2WLxPRJNeZaHnqLg4e
JMTI+8PdYvFUMKf/GV3RqlFRk8i45buGtVnotg7RcEAsRfbzkwHLHcSwIB6xCcxoTtrqpryelYkj
SRPX/BqbTrl+P1wSsrlDCHg3XuMeIVwZLSIyfM3eC3dZeM0GLJLOTp+vC6yTws+UrQB8TCY4Z5FG
Pi55556Hp03tLSScsgrnQjugc5ozHg5bKDt+lAzxr5P+bxUY+7pUD8Bwr1UNLLDEUoSWj7/sRfT3
3frKH4e3N3/bQwYuW5LZShwD8X1qemB9VfRTRKjnLBTHG/Mwb6UVu0aRgjsLkpHNFnfPkhYuH2gw
IQO+k5PdHgNU5kdCZMix85rLk6CRXYDoyuyo7qDvgIgkaJ8ACmxEproO4BJmFDkDHYUY7poG7uZ4
/7SApjlyeCFjwBUPBkOMrlae8l3ef9aiQrDC5yJku0ryNNcVVZXT5qcoETG+ZSxcNomc3YIijrV2
rw6mOuyRguXsmPQKDvPUtsl12j3OrZwk+8LfZdR+ia77FudyjpWKmkV8c81FFFcqCIDo7650i7Di
Rbe9JzKb+IwVaVcjO5h0m8tKpYzHKYqZ5DXDC70kO9b9wJ9OoftjqhWM4c/EYX42M3IDvLgK3K3E
gxGHvd4dsgd9ncWi92EIZ3w0ezjoJoznKw9KCmWf8fg3ZLJDwGG3c+pU+s4mjOjSbeE26ijOrbAd
EEW83S3gR5rH0VkU8ED5Jts01NYGreDnokNcXHk0C3gZdMl6OT0xCvNy6KXiCTAT6jf0rXNTjUoI
leQY3LdZuKRg009yJXjftGRSjznel30yr+Crh03/Oqeb0OczES2o+XsWeF9jeQHjEnjIliJRLJK0
0k9KiU8Y61Mq+WJUGP7LCggaeupEWoJezuOilXhczWMswcqvNt7GAiqTWDfM7J6b1Aq2obVH74PR
CjVOjqdGVdrvWBdZPCJ1x2DR7/e2SiyFspdmCd0E0Dt0/GxgqIQF9zlHfdFssxzNScLlZmcuKvOk
mncawQcQAXnmjMuh0cKLZIFFByQ6DJIvtbeAGD/MNiYtIjdAfJ7pA5B2Ta9AAWNSk7uNZWLrhszK
gQid1d0aUwFkN7jgsAM6LUwxgbmBLi7v0MxNb3TURc62Lh2rLPAe/rIKNc6c3rMUo6SWxnwrqAsE
N5WmPK85G4waQnEgNTzXN5Iv5UrKhgT+QESuWDC2gcKBPTsl0eqST8V/EmcvsSYlIxZsy+L3DLTs
IWWuAMZbgotVk4lXXC5ITV/EHbJFYR+SIV2TfT3D/465XTx5LjSQ+fT9hNgvSvF1mCzauMHlzLjO
YuZGmmGhv0DCbR/zZur96A0JlrvFarhmYbMc7FhTR/k58MHeSFXAfQ5Ifww4DpkkhQMIg3yQBd4y
p2WmP3LhiOWLimPRsmDOZl/Gjj3hpkitFpNZCUMV6tJShTG7uftp7f6DMlmQuEdZzNRaAMMJ/plc
xG7sIOu1YYfKNVAHDleL1N5m3CANbEgFVSruvp96krv3NLyshRI14p2FNe7mEzIWIqEroUfKtAb5
FKk16WPNQXcSn2Y7m0/xIiuzdLPCEIVOWf7BrjQbSazSrWWAOi3xNjqLmtCM5XlrYglKt/i07x45
qLUwT4R6Mkise46Frt3hjiWbq+KhABCgeS23riShdXMBWBxUrSUmOvxLXUXkbRLu7HIlNxWW889I
HLSP/UBWCBPaaK6Vo/VsV6wtTkUSbuV8RF4NCOxzLoH+6w/VjreK6l5vPj7YmJzCTnIKWjsTk7E3
MZrNAzXVXj+nounn+Rmv2YtPDEpcDHaL905hS5fHM620ZyAKCxsZZ8PAjutbQLOr1CsQxcF5DJQ/
gxhhR4Gd+IzUSjDSH7CAmgaEaYNQYvCMNegUo21xoY4i1fJHWl7h7hKyBuwSG9CvY7dK4oPa45pz
AHj8QtQvKhDnjbZsrVr1cbNVlKnSgCFE7PqNMoycdu85yOreYp/a1LT4104HvaaHp7zb7CBABfMH
exnKkoy0VdNnKpCoSImpaC49u7ulJMnJ4E4IrBUGJC67M5gYdYz008EYbOtdfJte4mJjrPaCUbzq
aBpiNIqwJngOl2O9hr8pd62Nr+CVQXlrcGQB1s8g0fMULLvfLRtwCCtdfsevPrE3KnmZedng7Os8
a0dyTwPn0derOp8bxyQLd2rmq7B59o76fCV0HIAGyZaCvK4gI3Rj3AsbOGj3PFeJBxREEM2TgSVU
k1hMj1D/958HpA65ZGxhwcmxSZmBkSmM76YubPytuM6YohsDqIlKKQiMQF31CacViRG26l0KWRo3
LzdlaXGnRApIjZivJbXvxdg0Z1x2eXh7PVEKcwBh1p53euNnri8jhvpvG+97Zvq70owk945ZKZ1b
d6AxtAiuQCJKnB/LmK+grtAYFXGyzrNIcQASW3RWmjRN8uhLwmk03aXLxGVL1WqL9wc9NKLRy+5g
5CMZNNcfymIlXzGSsbusbxFStsLlEYyujWsLdsnYnLQ42XTQR7w6HNPZ7hvaMcvy+I9DcADOJAIO
mrbh1EBlb1rDJ9VHgqc00KYj8VvtcM2vhzRVbL+lIxkHdM8SgeJRr/pBvsoeRsxrqY4gOt04D79O
Hg1UhsRptJCpKQf7GiepIwCHJlj+XXO91cufg/1cRn2qcQygOUtuFarxkUrwZyK0qhN9vaQ+TPBh
RXIVzQ+uRHWSQQYVeih+tNkbQncs23DkcTSe4DTKSysM7fyKM7KNDN8mYZFmvKxi8P7AhvbCqptu
zbisgPqhRm0QWJUY1yBzLPzO3wmgn2Dj2XrUq0uLr8xbS4cVeJ8DdcFMXAdPKGKe/qP1C1bDrQ4u
thTWvQdZbEWC/0Ufq5F+/5ZBl4dp4aVxqzYT7Ga8kGTmXn+spAcjeIGHq+80yQhLgJ5MaFQCM7ZS
XlUz+PVpd6nkxL+GesT0qElrE9i4d+Md4yIdt8cpxpzVJXfBj3cGn4DFeU+O6tGxlUX+WRKGLzsJ
yoLtfVDQmPIKw4b/rXOdffu4SjNgmWA2qkJBOiEXB2QauezFGkqFrWqPo5GtQze7jyi4lrU8Tb9q
4w9Zmtq/jEIdDf+JTZTmM5dA0evM0yBBCobP+9P6KO8HA8azak7zIebw00aqQ/t0E7B4+dfdUo+u
0B3UP95tYRIxAMCcZftYco7+cZnYP6PhD98kBPb4M8Lil9H6tOjMZgmQq2jwztrqOszvizCdRL8I
1XEX28Yzi2b6t/D6UldPAdGKcjg9F8XTbJOGapoHl7bTTyUDHP/KzopP7WNyY/0N2kZyFptnVif+
sVHY2LDIzQx6XH9+tXXbqKTXBQaMouQ5e6sZ6wV2XP+cPYWDtpLW8Jn1d3Y/8eX/QVR0E3lHQuzO
G5B9IvggMpX1lEcqqw4A7QfWOZNkhBfXiMb3nNI3XSzqhxVBxjv1gwia1BxfR3bBarpRqKFbfZ0m
NbUHgX9F3J5g+yZKRaG3dL241g59PM4QCArBVgnrHJPfNlL5xDN7q/auMQzWSb/dtOBLj8LHa67F
v8mNHLsYMHhQ8rWzqqWS0yf8aFglQcSTWTSM2ug8Lwxv8V6zn0tGJZQbFdHw8VCiI9bYl0j0KzOM
1v91im+XbrMlaeSBXGFuRrYw07a6fYKsKnZdaPQF+akNZ7fPs5b9A4tIRyoPfFyfTx5ytDVz90z+
XxG4646KQA4cdW6xWofaKNFf35p5G5EtUyvtUokSnAjERZWKVdkj1+9GhMr6KYkb7oq5dOezzZc9
tGMEBQe8Vfxjuhhu7G+WLp6wwdcpTSRpiCVpVoMBiw6Wn1dfbLzD014qalqMgIfwWN9jQX/fP412
vTaSpScLKVRLmjY2L466biRL0EjBz8SrrY+As46WIMdtAIkp3+vSdUrrUm2VQGzrbP/HGJGk7yGI
w0tLaWOmKtUKUmLeioCrl0T1oNCQUXfFO481jgB1c4hp1YfFWq7/6zD5Wpm89kkFeo58h4wO/H2j
3HlVVG4tLj7HPNpBW0KxJoQ1cOukhJHKb4g3DhJg5APqbH9nEnfBeVYJHFQsNvGpe7wT7d48mH8f
wrQNnwu9UmdN5UDgzA70H8qjKy5Y6kuEGavY7Frig+SeJ5LPCmm/MCxSWWOp7iwUm7H6bC8Us6Ph
C2U49v05AeCgLX5smbZ6F5L6r5ZoM1nrEVMl0c83eXUNlPbEot4gabDrccCji8UeJsIoGVxZhNTr
KY4CLBpAUYPmG4o1I6sbNUuZAGLeUWk1X6K3FjeY6nB42kAhu6dmLeAxyxlBQtPi6/sR2bbGCwuR
St0IqYrisHy/XtjCCT6PYZTucuvVXhgAf6Bg/ep6Ma/hFGwsgmij9IJi7wMy6OAMyT4fbXKAUT1L
dofMYNDCStL4MNvIlAYKEEapvwMoo/qK+D+vqLw9gOYl8hjfYPydKvfkJ7aLxT2tZvcbvrmHGPgH
SjBTJELH8cPQ3xl15+Hsb4l8oKc8fPAryPZw89ZuVJ75NxZfVswvFQRusAuvU+Qua7AeDrHMcZXd
GSDl0L45DoD8UUIBN44MXL1hvovzz73+ufF/6I7fRFB77oH+7OVty8njYAT1jWvvCCeqBPNbG7d3
mi5Z5WIdrNesZTWepMY8tOCQwuvEKczOdCCbPdV4uBzFC+++5kDdFa0M3UzfS/Nj2NQ8JOEHU1gC
u9cUtkvEx/8Px6IVphaGalbTq/j5jgWewh+FbQAIc7j7ClhaoLUI4eOZaILYw73ql+oAZkpqLg6q
LQUvhqYMk5XRrLpq8hVKHK4EdiDj43HhjzzBru3XJD6o4pVzwJA1JkSy4PpXfAxEQE1l+QCMIHH3
WxRE1IUUxqRPUCfUV/NX0JYYL7rMyqy8zL6gSQH9vQCT7l3FDKwcVQvAp47e5AqimYUm5thjgW5k
qWd0ULFbaSrYaK+gG1YkMDDVO4G/78UmNpWZv4bJtsZsBzc1Ha+gbCC2AsljoCEV+tOHYBm8Qf95
7mgdzHmvjFlfjWF93LgsaBcxWtdff32CUEC6tvr3pfx6PFnxsCmp9MZV3liTwh8Jz6HO7cO6Tpba
CWdGVPboddBbjiS/yK6ecwIPqkDOI782ffJxWNEkLDFNffLPivFU0jSQbDmolITmfn4U92YyzdAR
gHeBMhMAIhFOSJ4UVhNytY+PjZgN0QVoivRLxYBuhnxkyOCXdA/DDACO20CrnnfSP0jyTbjkCwZK
ITG435QqGn9ofSJbFWxFwYtpeCikZamepRn2B8GDVHsfXHPoQDN6/YBIMie/q50KbQnHy8O4YvRc
WZqoamOMcLa11pPrquLWaZhw2xMZiWFlLhYWWYw8qA9aFvaIViSSyZiqWpWI376Anre4aSD8X+Wh
aqad/AUYC4k9/cQ2zWOztf9tZtf9HWd1mbkVG8+MN8idgCN9lDeS+uCUUCEFymQiKrvG29BcOVvQ
WT5KzVrQ0Mf3YyOu3e2x7EZrFf6BOXfNg0p6J+3O2UP5dgSaH/MUJBPbv3kZC7JuGNA815adOfct
VnO8vtlEkD6oJB9E03Q8kObZyuWmZz1jcozGuCjOainzYMGi8pbUS8XGLsv08IiMyidG6WarkMHe
LzY1/1mwN+it8FkFw6KvghrCu9MEDDWsd3kxjl+kwfp8L6bTeR+2oH5ddPTk2cY87xlsr7Koh3Ox
izqVdiXAjvdlg29tYOgQPdImxk3IZM5+gxkA7bYVYd7oYRsLHXD6UsVJIM+11PnqgSKyWFobZiNk
mBRTpPW18uzzTx9KH9YE/JHSEh28rm2tvx4w4rT4rH4U0TpLDFUiIQAEzqP4mTDmbMIGO9WctUzZ
wJ+dgwZVxGWXCJG2UWTPWogk9YWkz1ClH7JrOqH9n/K9bSqUPZSAndJSSUgktYiESXYdO/BLaNnS
uqYKd4iz7YFB3FaLCw19Ya0EVW4kFrei4Lg1Vc7bQoOWKvY3u/QWNYQLA4Bym+jSe8FYZy27jIpb
r0KWQ5I0WSeEXsrltIoAQvxyuTuM4WyF5gXBCY1P+TrYvFKIjwnCpuP3a292JaJUN1DZyCzYjCSH
PPQcknyFpRq89I0pYAAtresZ31crqsjQ45ll4kryVLAu6KLTvE+sBHccUFPTwg9n6QT1PjTr3y/f
/TRb0PV7vYZLK6qnGnI0LbX4M4ZRcuIFfo/xnBIhD2HeqxacVR5y/ofhUFOLX1yvSHcRtTQpWVhp
ycx+heh7H5s7weSEyUBaUvNmLRnjmXO/tBxcbE9tlmyD4//pe59//aUkDUuTx8VOcC7EOetn58of
UWUBCqI8F41QzIaOXqFAy6hdfClEBLh/UbPSVnn9PG1AUW5jDpN0OZIdpl4lEIdlzpNqhLUepjt0
V4p9X4jdLc1uetYlzxdpgbvmBqR3mBAHVOu0nplWMSlbb0cnmLadjAyWClSlIUFT4O6otDqAVc1L
1vYRNl0o2PnDBXrT8ImmUIusxjpbWmsIS6HSsmdvFTXfknFBpTvA//iH1o7JKtvF1O0KIF11kld1
xxQwqSwolZmWS/yBwi8R22onAYWV7sOXo3uXTvQ0kU8+pHeISnyIIjesI5VOay7rxnx9L9Dh2lsL
WLhrUte+050N3fAaZCymlYnqXViruStWw+FgwKabNs52+HmQt13MX5a9FFr0WXrl77IdIBLeNoFU
BfqAsF5LrytTIzCoIShYnvKYPY40N9GepLKRDxbXp9y2s2SAf6ZmJmI7Vh+GGWtkYtxGd/Fl2gvH
7sk/huh51avFTG2gpfpBeVfRL6ZOXEzfMXG1ZOhd8kKxjN8bspcZCTAIpx2dtK0EWNOLd7Mpg7O4
Pra5ZdUWrQ0mjWgp0SW/U/fxQiqzaX1/IPbeALNOlie3Oc2mToTOPDF85z6mEJ2W6v0L/4ooADCJ
A5OmFVE4kApY1GjgZuKnqCfi1MDjxLVmAyE70HVhBPagWgRViRP6PFjG6Ow+en/VfHvdyaXekGWB
aEfjlu2IEpf7cBa+Q3AVBm00S/BDsiY1dy251xIIeYBIUWo/fc9x8bzPHXSB/1MeUR3KyQH5mFkT
f1wFcsUQZIk1aSkaaY80ttvmV/qBbwZVBQtMVM5uXSnGkTzWrVzBIQAcsMKcduE7y/4nCiIVustM
0JIEByxEFFE4v7joQAvaGLF7K9UJkbmQSF8e+5sLzpWCVlzfn3pP3JlKtPXshTHBkztBht/j/QJq
flpXskcQIiaoLcYXfHLB9VoutABZofvscHBiMWfRpPv4DJfNfbIAHO8T8tH9yNt2CyA+7W71x00N
naGAD6cD+VWSZXvuxX9CE/YtCDi80PJOLsrxDjjPDbk9jgeRE5zW/J+Ziwv2nQCTnw0ZAoOLlnJZ
W4o1ykdMBE81vWKnU+ID9zBAS/ol+5irxSBj6zYwb+T++ppAhuLJtPRUVk85vA+/B9MPtWBfP2HY
S1HNMVL5uPSeeEMCiBnpOv6OKHXzQFlhSN6AKD+50fbn3QfrqIl7sDGx/QCEe0KCfHsWVMtaREcx
33VRSOdscjLSXpq6fKFQQmDBvlJ1GIa8fX2qfhbgbH89eUuaaNUSpz/Cze1/VJERAGgqoDqBDuUq
CSVyTtq1TTLqZvlHtgT6Ms9JLupzxg5/T9Q3U7/RI64b5KyF3hBmOusHvkd6MsONGk25RqboOLuV
xDgJ/LAvuH4nb4TXQb7zEeOik18R7KunKCzucykW7eSfafml20R5ZJc0qIzyniaLXYgFMybLw+3C
8eW4H+O42L4FCaBPkce4mlM3I2RCLRtTwgx9NI205Yj5QnQELQs3tqEYorE7Dyr8gE+J3P7v9c8U
XbxVcrv2vWVMd6jqI0d9JHjW7IXPn8OGRhmmCNL17TRi+FAeQ2PzurfFnBGTAB9m4Z5YQIYhSx8U
WGCz54+8KpAhuZhBQejhnHX+x3zhj2iLB3Fm5llqjsRDGGtE6ae+GZ89vFPFUfDRTqSKH/BksuU9
xa8FB1r3FdtIM0kRIT94hdcvUCadAPEk3tCWDfNCVQnoE9T5dM87u7B7VcQ36YGVDFX3QFErTuB3
IKdnJJrWpufHMLXjVfU52pJYwTz1sFwpNcMMXsmUrSHhOvJu9yttLuZwdjdqbvSfCGuF59t8FyP2
4h2veXjBZ5TlUO04F2Z7ILNeZiOhf1vsTAyM7f8qPPGGoWm8zBJnjs1ekTZjtq1VmikKof4gHfDe
jkkk0rM2cfKSl6mEvCZRf3mzNmsfgAEaA2XWZMBs2mgxEkolE40nJpaj0HdbuwPSlIV5SwEJDn7i
zZPtVjWj9/8ji+10rnRSNrNOrdt7OU4LaKuxIAmnL8iCfBSobp0JDWoysjZMXps2DM31fdNJFNlc
6tNSHsE2PYs+CEp9Eku9HZat4Zd++CBKTGBF7Rvonwe/VRW4WKSKl8GgG0jtJg9WddfAYamOGMqh
xyo95d1mhrLyce3zfeFzkEGnQzIj1M0CmgJqAsGQ/ygM0BF2IxqASAAtIrsthM6pOfbfspp2yMW6
FGPnsApsQO6dVoHy/yN8hJJxLKnvacb4js5vSIB1XIR/8xWHl0dcMnUZnKDycY5Kt0puvLO0wkdD
hj27T+elBaG2LodSzBNbvUz5+A97PoieVlBpR1Hsuy9A+DlEcsCGTRHzikQm9lP7HmudZrkzqydJ
aSZCWzc+BNRPWygMiSHJ7mKmXM60X0JCyY/xueauNzI8diXDXFKPjtRhYdGYnilFvcfVFesxlT/3
COtb/QfQtCnlHNtPr+UgYYu5NCeNuDpfh9V0bip9aAJlpnNOHois2fJqBjKxLHvLF5S9MD6acEkc
DXVJnVEui3X9RvGNy8E8DFEycjnus4Jj/+tFq7wHZ93MPSifEsYW9+SyBW1V6RTvFAJtXkzws+Db
CjXZzAZMAlAcCPN/Vl7Zt6fJFrPRLgIPIL+u88ZWJeyw8IMe7jod9TQ6UrmbvyfhvWRZw3RqUbgV
RrkmAdz7uqMr4BtaMP1FqSmu/2QgcYcK3HXQcKJkyUTIM251ob4Cka04ybueMFCF//yTKD65A//7
okZkBI23T9g6AUz2BiwjNWBF6itJcB65f7HflsWl3gLZZ7ayAgc859CZ2qvD+lM4tWLbYvldUNSy
JWJI4HQpNwYCKCiQwVn+NdGQiAQmc8clD8IZzuGdza8L4YTz29cs050C7CYh4+Cp62zF5y7uzWeY
xXaxvGwsuLyjMGUQRcB/DYQdC9I38BWAX0UcBSFX+RlutpmyTbKs7CYDpXl0/Rzt5X2YGKe+3lJt
LEfSu9CysJCS1V8153suOK4h1tJj3W5p5WsMKupmhis8JIzkN1Vd92zHEBiJC0Eb5+v6RKnsNIMU
mz68ELveYhshrE9iYnD+7OH+TF2mnq35cmdfWr2hMKEtuHvdprj9VURSYY6MJjzv+yuqOnCVXzf0
p3LeQagUUds//p8J8EvZRtVGY86sNafDd/4cyA9o9iTG/AL46bav6MUe6Jf9c16fYKEFPxl6lD39
2r3SR4O4NWG8SJaH8OpHkIwIxKYLqUGoA3+V9kRZGenECLwOaNLllIBN4RbIyEwd2+V/UwEB8unM
5DB/DxfrSVGC4fJ1UPwithjuhcber5/UiHYgaCkIuJiuUk3FlhI11IWE+RGZsn9upWH4ft4UALwp
oI48YqpLWj3apRJUsNIhccd0U+mi3hB7pL1UXH3DBv9EhreKqNzrRwHGaJMoyiBL3WlegwUdyYIt
QNvNX8o8ArXzvIpREbLQPsl4b2mnGmDn8NOxK6ACwtL9XHFfS6GUFypdgpsRGDxZV8wmdHYTShGh
S3h2s++0/PhvvvnOIPnQQHrinT6QoD0sNumQLlEEBgs6/2OgovuQ9JiFXmHO1R+FMVAA8VbyytmF
wawiVF6Cjlq/FErWNxeRduAOjvaZAhi1+KCwNc5+2grQ5XnnJVcVKwnmpWTxw84zhprhwj59PBq2
5WNKFkpSyVkYzpasmXNK+3hDCtNSB0tPgzTWrF4fgZ7xBwgCKmy29hVRseZZYTQC7PIZZhWDn0Yx
/OVKUjNu5Nl8PvYygXUuQAYD2xuUNDi86wqpTepG8NTPTxDvJtjWJ0jCKHMIYdgwDbzVcegQ4E6g
ziB362dPU6L32xtrg5Ke8oGwZHwEteGvf2zusqP7VGMgiU6ZK9IBCDCLYxkvbuqxcuEfTpncKcXn
Ia6uHZom7USKGaiep+How1J4L14vcKb2mRkYT35irf3HZysIY2k0aHsmiCULE8bRRn5zjgYOdjFL
rAzcKxCSNdFes3xXBrYzzMMxWD22HMghUk5C492rBz3IPlchDZioou9JrbfHTIOG6uH12FkMv3Y1
paZAKtnlqESOkhx06Au1+w5leW9YM8+CVaILsVVbljwv+wAd13mAHPIwi9YcjTbOznegPcPdZcXq
yYD+YwxY7RmkujkJKxk9uTowcn9PN4SVWRLSf4owBbs4luhzH+eyMgeAO78Xmw70Rua5/ydB6o3N
DqM1Yq8+DzBMOqPQZNLyJKJ+vXD+Toc4gJ3PN5hsIiOZvphc+uRaDY91DUwBPLVF8tibISPkdXXP
wMZjmkmDLh/XMOsr3hio5TGZ0KkhMRJZ6YwCjhwXcS9IxNaC/Tku6+ARxOJpTmzCTIiUQQu/+lsR
yoN+7Ka2nYhaCn5nAO/kdAI0Tl+OnuOl9ujh6J1DTzqhS9IvgPKllGOm94NDJKLlOsyQFt7jUsFK
wWAaCD42YXM2mpIi/rnf72hsDNPqvJxJXG8NWQuaBR9GkW1HzGkAQIi0ALkAoVAIp7fZTV3yDl53
dBGOHEeXdWqIgC57ctY5sLaWusorg1jB9NS66xeBnFG5oNJIQGFI8V42t6KlVA1sbgJ6C0caIQKe
nb85FJi/SWK97Q/F7a4cnTOYLlS4CbMAj+Oo1hP3fNEkU7uiNEljYlcw7R1vqWAuFBThf/P8aKz3
vPVoYU0qsvaNun2oU20NUEuMMSrEAewVWAxBPDXD7n2e/O87COaMsn9o99Qdvkj+r2EClLoqxTnq
AS1BrO6nxDWdQH6SzGAWW0Oem7ORSrPbZWlb89z4NtmADX0QN5Sli6d/BfoXxadAdTtsWN5AZgDz
PxVYDyWU/YbyAABx6O8Bvq60rRfz0FkqG5yEcOf2ZC2WnS2NnMIgNGm59kFWPFCvx5bMujFTanw6
CCxBQT7UIJLJAgwC/BZ1IrfSsDCBajnmK/2DCxzURUw+sHOLRSq5w0eHYYMPCuEj57Aw6HaD8hKB
GY06tH8cyHljagA86RoPu6LlSDNw//sU/o2fQDFZpj3zjmoG1g9jXRTDmq6TOoQZ4+AvEQCAEm+j
GH+ql3UT6q7UQyP6ztnBbjZflc/P436Okc71kuWIxTM79+qiP2B7nzbO1/HVqvr3PG0xvJtYhJKB
LLneBg2MJ+lMSIq+Fc0Kn7aLsRgXQJICCcEyWZ2TGCK6wwSUu8jGrPuW9AJnYlASkElUr7ekyjxx
2k9YjA/x0IQuqOrtrZ4gcia/gtbd6MqeIUeflEY/8zFCvb3ocDnpbPwg9bX3RsK4cmPg2AreVGMZ
TH5V2znVdwmqwfDwCVv5xp767lsjQNozw7jmW1GcT7+1GOOGCAn1roqpng0MB1hw2BZJbRVCEUGl
i/DVOveEfy9/1ein87Q/WQ3a1ZRY38RZbKOhKboc1MoP27ir9jnu3q5XP/6yXYLeEQsZGTZnY450
LoSGBiyY8rXC/Fl7Y+/rEo002c7XQ2AWny1EEKqP6ufVeSkUWqFnqL14Z7pDcIxVrd0Lx+MqGV0+
TFsFWDWxHxJKdH0yAOYrWS0xzvNPAYx+Sts/gbrkWzmoKuNo4ehZkWC1KtD73XEYGYHyQOPF+2g5
oHrmVmKmaKz+PVjLZJSsYNSCdMY7bAoujDYHnehpuS1CswqW0TIeBMJmxtTZ5ATfCWBlTTsFOr12
Ox/5FNlvxiTzNCoXE5KmJu0XPtuyUwanoHcjls7HUvkhRmZLvDUXfddroXua7VLotoTh059huMda
7cDvZnDmaEHd5RAgrJ6YhSHHsCcD2tyuhE9a4FmRb6hRg2bOHyioIud4OP/NbLoVyw1nfslo3lRS
AuMgqrw+AptJFpWMeXEXubcnEzFwwurKd2YsMM+R7kB7BH+DSqkFezOVZp1BhQkEC4qtuuWhVBbn
+8n3Mf5qQ8VLNF763oJnJ1DV4+E+oksR8Sp/fFnruoqXIfo9/r+qCwVlevKrJcSDEuqpc9rFQohN
gnVetfPAWs3HUByx2HT6zzHQbfviipe07pKRZKiUrtKaCPEAYWV/KvdUDJURSe/37MibNJxMP1Ja
Y9OibqvTmaDCcBjVpNy0LTPs8LeWe2AM/6w7sK4Kb5SgJxR58RJoRypPUgJM04xHX2RFr7/G/cNc
mFCBxnHg6xS1ed/w41UbpjiNOT0Xz48U0qdyI4wpPvuAVJo64DjYX5YTgalPvglUtSfmWgeEprbv
NaikbrBk8+3NMjZxkbmpxs08K7X+doCvuE2otOHv/Fmq5WNv59JWi/5fnsdFodA6Rc4hwwIpqEl8
86iJ40ANhIJhE8YezGvbedHKL1yvPB85tN0O3DvdKeKpI19qnlzGmQcgp9tHwVPGzNVcsX766yKm
FXuMhgeLSn1/YBE6pGaLrCmlN+s5aYqWYhLXKjWvWilzs3Zvtd+u5NITvkPGBI58g2zFM+sg9yqX
0sTrMYRMX9lDR4OEFiIM7Arq9eICkVZuOIHikT/8e6mQY6vgKc5DdmkbXQuBZwh/gx6hF55BCs0S
+zh9gRyxg7zFEF1wIpuTvMqxzRTKm4xauXUprU68gR2Ftg62A1lPo6qsVxYX5WHtgYZJSeBXZ0xc
/td2TtvFf9BCYP9pXwpPwtLRgurScM14PujmSAoTuFyksh7rcPe69Mwap6YtEytL7Ci+mZJc8Etb
/AvstayTRn+5sPMHesMymX836hKNSwJYDgXRmxbmaKBGCY5m0X2fjJs0Qu3CcnGzRM7o/evX1Ar/
B9rwtgrT6nECvNdmYNCmuEfR6zGSBWHmRFxaAY2FdQeGmkn3+x0/hZH7S+n0Om3oL+mFuWY2CLNw
sBlwOnKYAl30RA7Z+nxeERoQfHqlifc3hdjAet1YvCceoE5RzyPG0h4haqwAqvdwU2D/Itz/iiOh
Pqdlk3CiM9J12j7s/IXZzcoyuckG2txRVIGK8w/VafK2ApGzlVC+k6/Nrgw4jSNYDsMEKjhw8GnP
JOeYTlufNvq9ehmhJSnW19S7C+qOHd4gQmybGBs//bVeP0YTF+o1q1WdujFlbJeIZw0JDyJDJ/+l
C3hQI564lqHNL3EsDJtf/6HtrMfbHlK//nFmGjpg7MZxAey6y8l/kj9ooB70A6m3Bz3E5r4l/FtW
SV5X9axViIP+KeYuaNbCZ07DPQTcyIg1am+AmkLh8NyzRKquWHGZt1amjT9zdMaYCeBxdqc3PrBI
5aSJczuhaxkWif9zjTLLxqIaj/mNx/K6+p7vxTRq60AbRk3mGKCAu3WD89nUXxoV6eQ++kDTFla7
9wRLkqrB38ezgqsYstsklKnSWfKSgwdGyPkG90xQnGlXyEzQcdoVCbzqzJQ7a6A2ZaAPFmeBtENq
jPTNVSUcYfGlhffis5lPgAUmtC2/HySqKu3CaJ8wV/u96MY9LoAFHU7SHTk0LzcH+HZsbP+LYfRv
yH7f//zlKmYN+NMCaA2O2AH2L+tO7CgBSPXoVVxhXp6vvICoMOU/LWvMbaJ9wFrcwu1MPwRmSu6z
Du+WicXu6ZbWZ7YczK0YGxEceOh1QrVokSctkgT8mVXospmFYmYmDsgBbHjvWszaCKtzDKowCQWa
PQ76eaKhxEkIa58Tk5kRbT/IofNGDQgl3e0+45Dg9xj+VcA7eM4rdPe4w/MPSTMQGsKVgHIhA1RZ
p0oJZMPUs3Qe5R1s7WRskzvm+dkdaKk2MQ6difXL+gbGIT/51NCHMhLy3Kzbp9R56WpWhAyQzQMh
YavPobIGhws0nNVurw5c+NhPA8tkB/PggC7lfTATHyYTYdao3pWP6HFoV//y9n10PbQ6A1NELuyb
Mq3cd/IOb4yIlER6nlzonQwgKwgkfOupiwRumiA/3lPZdLTIqM9KjcATyO+jsRPZonSAt5K0TxNJ
WDMMo3HpIj2DrO28jVc99wL674yM2Lg+dPoVf/2P9j9N4azCKeABJX53Hpq5o5SfpELlPs8MDyIQ
BGqEbPKHBYkkEoK/8H/Tgm8JKGXzG+vbau6DPnZD4mvjRKSIsEk7QSnDGAiCR28UuPiJIgON6BHv
XIwrySGt8TbUf1lgGh0JqMDvlLNeERtWTGRgEfRjT41q6CNoSDl2SWpdij3GtxdqNP9RdQdPgwU4
q6cNTetXwNYcaSBw0Of1sO1SW3N0fqyfuqqVb9idrRbBwVVV000Nuw6lmnoPNO4rm0bhs8XAz2Nd
SrWntQ9hRXe3faIRfyPWO2TMcHzC5PXQuaLgCc8Jx3H2Tw3lXMU4GVUn77D6+cHTVAKjjF3orGhY
sxbjgcPpq9Xjds3BWzNbVK4TJ7WsiBujjPeyeG5TBvW+T/myswKzpQ5rtDuTc25+hvOVHo1n+dUP
PDqE/rBwl1yRwGG0VFBJuqESmGlf4yfY9Mu+EFO/gtVUgGX3PrRgalt5XY1AG9ak9QRi+3HIiqBB
PbqQFidUmBaCwof82Z0+gk8TUOaqjhGyHWK+wV1FdXc2j8kdI0/hA1ezrWJTpWw5zFC6aUvUuL2S
gLI/+7TANy3gByjt1TEGDe0mPFYB4qMMs0S5QiMoX3pH7qEQ/fJkEKYSX0Yjfa9f4KPGZPHJD8g9
jf6ikchJ08XAXUxJg5O0F+dAUfYG/3Q/tZEJ2WIvceZda0/gQYDS42+1UYZkzqn/1qPZ525cRWBQ
SY2JRx2U35KoUdg2mbjLlpBqlKTu7ntjvavn1TdciuI0NWib5zAlIe+dUeKqC+uHM/pksGRLPtfs
vBc9uHzE8sHzFUW71mNU2QwLutZK2tFTb5m3+cyHlaQGEH0cFE4j4JXtHzKPzo9LmAZKRVKFA8jX
KzrqiDq64IZ3i2TOoeu99YImLS/YyIzwU2lgeep6FkFsGObInef7BsYH6WYoQmyPQ0PUH7UbB42e
UPD7l0TAFdiw7pOhSUf6h2urD+p+kE1WJTAiDQKS1jdIT9hplVzkN1pP5Rk9D1YiPnjayp41BAhu
pJIIoEJZB9UJN7X02nuZyS+v9wO5cO2WIfFku/gp8vpJGZWri1Tm34rRhGuxtDxWOWdy5kVyO23d
jrPI6FoxB3htEElbFDubtI8sgX8dRFboQjff3ZQa2rLb3iQSXIwVK7leN/UXd+BFmY0jXGoqfYxP
hw8HSB5MZTRQsJVy1x5PecAM9JDEVUhza7o17Ad12SoaGJiod6o50xeM+RvdzBQNC1Mfapauf5F9
ADAHuQZboEGUsNO/xxsS2vxbUyGxkJafJjtJOKm6sbM+IjNGwDl3/KL5Jxid40/V75C90BJcYQen
8A0wqMZbA6TdRncgfM0JxkZZNl2hu+ikw9gHUwOZ9g/UsOtqmRQ2XYkr1OUR8bTr4NbSSLI5GScz
yOFpKrT8dcVs0SD/hCkAUGXI8nEaT4YiTvnH/lp0K/MbguEy0MeX6r0wsugP/zyFqy5tvJcNlQW5
oCXUBNWKcpl9pMDcrBMQo6YTw5VXUKkazojXkpi3eh0Dv/3MQutBrwY/yuqa4dahBnDAbcc69Jot
YUCirqdsErE5Q6S6ZKcdk9BRd0KYC4swzwVtaFi0yV9f+84fIEI6yQUytq7aqxWTcooM/Hi4Qb+L
F4bBk0U98t9J5+2AZr4vh9gwL3YW4dE0yrmUubrkNspXcY/6sh9jBOHUFm6/MQ9AX846i/5n47dU
dnK0JYfvsPzmk61eLzl+r2vXhzVfi8J4t+57jXghkmZaFqlsKLeb/At9LGfNLzTQ4PPSLnyWFQGA
iqxwVEE1gymSVXKci2kZfHYjvrFPN4axw1oszXaBpKi9BZ1Ug4DBcUa+ZRVxZc3jHIEcLiJ1VQRO
GcLRC5txIlM60NLfFC3l2V8xUmJpzojeHSBpfEfDs+hKKvBQKvgdrTmQsYND1KCDwQ3xv2JtSIt1
0lxoqQp+fPpafpFVO5O7rzz4UMLUDCtfp+BJkivbAw26lKh61giwool730CXcQBIPURDReYVc55z
8A73VflkfQS89HhZdzC7tmiNsgNqZMq/yCfwj0dtnQY3NfUPB7PzRgzdxLd6HibuzIhXGmRhNE6Q
ifHmV/RoizWYHbO87T2A2ebnddusYJIa2oeb/kzj+JglOs1eyI4mxK0HLvgihXWLptH/hE7HSKIS
byr17N4wk4N+vmT8cIwspHZZ2CAfY6lCZbfKplPGyuJj6CjeDvcKR94uo7lx2Qt7HczgTRytNI/m
3eAZmuqLO7+RvVjYksAVarnWCje0JoNO+o3BBPgJXb0m3ZAKGw2gfBu6U/hX58/c/8ZYcZRsPqfl
Ma5TnUpkXlIgl3Di+RQP2t/eOaDVWbupJNcVjEV7wFXh6O/fT0K+XXlk9JZxizonLo3VQTZ/KAX9
Thm5jnt77fvppXFEB5ME2jlbVqL21BlNC8oo3TnD1R9qSmBVtwQCyavreKllfpDBi2M6wBLSIdnW
hO5aHgUs1cSbPEyeqhJCnNzpwVf4dJjyUgekvqmdWW+g+/rjZ/SacqvtmlT5Jj6SoPG748m2DoCT
670vlzRDaTz0v+HpwpSEf/2/k/jXKtsFPKDwcSW0E83nrNrMIUEsTrqsk95QAevexOsh15UGp4Fn
u0Ktnw3JsAow3leQLMW6RCjTd4TBjHn5NFlYOFI3kvJb0B+mJEhMR3HcrK0dp7Trnhie5YDxRFFn
HrROh7KcLebUmr82OfLN9RJ+GfoO17lImTQbZrLHRDzQgZ+UxwpyPFVLb1H80qCEPfandZW/eDPu
xn/7zvyxDu5yGdxF2U1TrnpHk3RILw0rSD9ksv2SOopdVkfrKYbiTDSJ6fqlR7RaakYwBMnbsS92
FoantB94LfH7DUN2rNRfDSbceVmedLEnxRAkvSGVTNFcWRGUspOVIPrHpMh8Z5/u6kwF6XklJdRF
CMymE+93kE/CdpvZ82Lt5n798zLcre5g70B3OOZFmZ5Jym/+sWzOBHnOTwe9/Yxe/8xi6a0ix90j
ZNrhEY8OqO5E4v7HBFO5uN72/W04Jqo17sdncNVSxIvzxC4OTvzyX0+Up4iR843shf3qse57PXa6
DJFwg+HziKNgEMhmICR3F5MHzUowKIJE7qaLFliL7gf8lyYdWb3oc66PSTJJBWaPWDVunn/J/WhP
d9N5YvLl/UZbhU0jtQMKQOKVD3VaC7rFCL30ir4CpKYOhXgtN836qM0vRM3OQqDQ/rtklGvnRm8g
hfjwPtzXGKOMlIEu4ktpGVQea6HHeC1Pxk338W71Qnj3lVYTqyTpbatagmilWwJP/OKuZXYYEuja
k1NSG6qPy/5ruZVDjp0qlEpxYmpcVLGH7434sTBq2VNx+WS5NgFGhTFOHdaqzGVjKTb5QiQZt+zD
EqhLWKy+yy7K73z74A1mHpNkOJplUFvbsrB6XuBSksG6BaM3RDUCkxgJ1QymVAakUg1SreGDNz7A
NM4DT9AwJL9XyVhifehPMxPjknZ5nJ0uTdVBViMvaya44Or1SID2b8SgnxQWbDpuNW9WuOL+n6bH
SikJTQ3arLzKoYuYgDP/JNDNO34BujuFE4dfwOOThaDRk0XVoMO7C1Lte+8OW4tWGt/4QGKMGOzb
+mWw7HxJ7Zg5ChcksFmQuvFNkqdgYffSDXXkNHfkPStyjuazFfZ9kw6YmgF+uKuy22h4keADT3aN
SB1VNJSewSsUiKGILKnAwrLhGM/By18GXGjbS+u1AOCmyUxt8r3WCudnO79MjPTb/iCO4EzCrr+a
EJYjYoKxDUBJ4jOgGwBo8MmDMsdjBvDMbpZ1LdmnNd9qyQEC1eZPyLw1xnRpBYkGAFF334R/BP6Z
0+JV+7jX4VEZNUmQ4ddhrUuuDcsDz+rAREIQCSOHw/IvENfl4xDK7EHYo/5awmMT0V+mPs2lGLSw
9x6kzI3Z/I4NMWPe5JRCslahmlpKD6G3A8XdoL3+P/6c5LNL+H87t65dTOjFaZkMGxPQaSU9Rrwi
2yBu/WOHvJmdk4nytZqjCC7Rvpk/+zqdrG6CRc61F+hNeyZKqb5wv9f3tc80jTpNEDpc6KptbO15
UfH2GJVxBNFAM7KmJPkXthdtq4jugMIrza6HcQtpi80HUoyV2ByUAQqv+7Q9+U8N2BLzCAt/DHXu
VIlM2ua1mPH4i3NDAAdiDhsGLfLlhOS7c8n1J8kISkubK+6gP5P1+cVs1FQ0oP0AaIUIaJV4FJhr
sSa7fWWfD41RKaLrhkAmK5Q+DjXwFll4nOHbqn/WVngJEyNsDnVQQ5GqFP8zhtqqOkuB2Acg2wvg
E3crTq+4MhTb74EQ7AL9zXeVtTEmdNYHu2SGUbkws0bBa4ywl7YVqfkpUrA8TFGvGB8U4vyjpPzG
ubbYuNG677VqI255/4M+CfzLjqpOk3F01/ol3A+BHTE2zoZgkz4AhX7/CcPv8Bgi10AsyrPHpPuo
nbLBDfjgqVvNM3ExVWJeoqrlFsQQU+oD/lSJu7zFsY0n8SpMkyfBIJGHwNnmscrkM6eU7EB5hKFU
Hl5Q2Pw2RUT/QzUqwypF5LzTW2+y6CoaZsNkKhubC8iq+I8Lk1N6tDJTl8fWDgT5f+vKI/cnItRV
ob4tHElVvbJYNYVBJsHuXTi0SLEWr8FTR7iBJYX41cZTKjU9eBPq2lnqdsMpwGrPoekCzohm7Bpi
fhnYpk37XnAPWSvns1x8Qi0Z3Z+IRgb228fbov4qPWEy+hDcCarG7vpigk63xUziqXYmYzf2v3c7
jnWcmkAWMrO6MHgiZAMGHHeJEfqNzQN6Rz84GdYlX27wnBoahUcrUauXnOVJBgm5O3uJuRnQfnMt
SEAMutNUCyzWQKZlWJSmuMUoIFIyTiveSs7UaMejoK1oADgRJy2JXPZUnwI0wsyFgowP2dP9yKZK
jJSy+wkMqbI6BtF1aMgajQSKpGSizySgDIsWDDRCmUgKdgicxq49rgFPRjKuf/lPybThg4YYCY8f
vHg3qvG5AjdFNSHPM94t0KkraqPH6bMKDjMBpQGE2ysNaHc5UTlCX3AghMro2XD56+/X/zZGQrPy
9Pv+xxJn0DYM1/Kkr5sxBD64WFe/318gLUW1k6oC0YXGX8erAMRACDnApwCs0zzcUiSFjOnSrjBs
3sqZ4MFXOCzspWP9Ihvr73UhSb9vurastexEskOwE2WmPKPtz8NZMtp+L6febLjln4cmlRV2LeyP
Uxajwd7qfIpf03W5E/JsoNr/AHnKVNMs1ovUJro+ewgRk36gNzS1GAEZRXHefScL0teBEe4G6aAm
RxNKG3Wolv7RBaUpte3ggNuMoc+at5Sr05jvmpcXAKe75DmFjvAbRBEgG2hw4XTyDy4l1Av7YT0k
HYrMy1BVuh2AbEDePmy5y1+Tjg9yp8kn3E1fnkR6sOt0ZlIqj8Y338jFVXLCLgjWEiEcyL06EO3C
Hq8zBOVvH6WFchD0GECQebzkySSllQW8Jhz0m1LRm03x8HxOBZt/JwLKN0csriHaW85l4K1SYoO6
Z4kMrHF160TLu62RQjGfLdOnfcytceKamRbiN4AsUJAG1zJSrY74QC/IXunobDRw5rrO2zp8vB7V
s+DyxqJNM6p9U2NUI1w7y8n5xkXD1pJ8/D7x2/MUvUJhUAfe8xs0BC+NyZWSywqaB+ezXvtsbJmp
LdZM3fVD85RGFWlN6ae642iiXeVp/EBva+VzGL4MJSu6meoLGV56gV8PO0TktZXMBb9vqY115+lc
H4geOiebySFLOaKYPo3VuqsBO1zd66GRSk9uMZnjal98kpHOQt8zGoB5d28DTDWBIjL0DLij9CHA
9/EdLXLqKXmBo/sMsG7QrgW0y78t/fnUO/oeSHQq2STKgegvFNqGvibhUYuZl3XB4xsNhN6xNMtx
/qb05aQ8DEN3BWVzZVj+R6Deg22o3f5Bnp448v26djfAB9sKWbKYfXIT+R+8AxLc5wBZRlVgM4RB
ivxoerSBnZF/6scbAyRQhBlPauNIr30B2XLb60g3ih7ZJJiPHHQ8s8tEm+pbHwSgpdqODnLuwYKp
GqWeJqJYTMIF23ZG3ciFEDlF/oe4mjg10zO1k5WTyUY7JpxihbNlgaDUcet3zHjKnYJt36Gt9CH9
1AeXqDsnPU8DNes2XtN9OJ44PS5VY6rf8OL914rSQy8W24XB057nyeOmhKXCMnZyVZu8hnqjvt2m
E6OK71veR7g8xECKJWsuSnQIcBN/kLq1Gpx3+uIA4ee2k8FUvyaavcjC4Hmxvi8+idNrg4S83LW+
jGWd6+ZG41k2RsJA+i8aQ4xNabwwjBqdm1ECkG1r7vAUxPQdp2dRakbOneBC24EdYFJBjxDus5eD
gzVIcYuf+qIcpR/1bsHUZP4OauY1oWYpyCbq86oei1FxDuAxayBN9atWAw3nQdQMsvSdZAiBQ1vj
UH6iGUnV7mLfOmhFr18QREoU4QWzgBD02jcrj5ER0SiAs39GLRIIp9+uajyQETWT/1SBuHi/T9Kc
B2EJBjvLpTlXcO7upMIH5yuAjx/jx3ikLW94iP+G4/GQBzD2sZqh1kPnmPxwC1HnEBiZNyvbg43g
zJ44Uxo1cIHER6UBRlvs1q7ltXMynHQhr9t5+0fClkXwrQfz0jDFY+YYeFpMdAAjQICdkDCs8kiG
bn0W98q9UWam33Jsf6Rh0b2GJN4ev85Y3q5CxhF3afa+XaYQQuCLAK8Ai8Fv+50dTOWvBqSg439N
+Qr4I+stP4qSLquJBFvLNV2LOkpLcHCwWYImbFklsvLttPfLyNHQPelIampX5cCSiawsMmT04pOe
GRSeE28X9upVGqLaRMglEEZPqNRGFcEv2u56TOP9PyhJ7fgl4QvzDeS5uk8NbEX/AtJH/kZze9E9
3kSE2VaE0h+fd+1MrHy/mqpk/oqu4RaOmlFCYRDq/X/rY8QrAKDsDxAYDIb0QTWpOp8Go22OuVZc
tCvWK1jCFXcHajOnvShRaHK12i1ITlI+68yV6gV6XLzg6lCEm84lvVdtc1OMlpH3eLroBxxdF5Xc
TejkcjG0IU4LOJpiZ6xddmYDu5X/jn4+QjkScVBA1ToAbodTZmlNjDMkpwQiPdabohYaIPIna35q
bf5iqHxti/DrESz07akJl1AKVqvB4iteze3CukVgRG5jhJW896XyXq6FrJHfIiCKXdlfVl/VYoP9
1m0xwaUPuc7bp7rvMo05ointAyO8cWPjut3WUn3OorobfEWayBCWChdLtm9oU0L3q93cNM7yXglz
GlQ5fu73dAa6jO60vvjBBVHD5WJkM4MOaXk3uV32vPq4dY1Fhd4JGg81TboYFIj1GuqFyucWOcxC
NyeajK8MyBGHXgBqd8fODoSp+xI4hfDbjoEKgEx0BsvKKkzICQ8EiyVv3ktWKUre4kAAb6pvilsi
u2Pd+jM1hJJ5GOse605U9AqpkQFrfsGXP7qFKyVzr/0l/lzlweRylEk0z/UA9MxSUTpbLeG5pHms
mL/U3jkNoV2knNC5aPjOwNRY0uYIS14qhcHwYQyMGzTbCaHwYdzzOmRwsFlFlX6J0CxsHvU2myDr
k4C3EeGguPHPY8b0ClKeP6bQmzccHDegIsWYcmw3QOqdxWP5hhlcHVRz5pPeIXarI0U2kmJ9VJXO
PYecoRFW4PKblwLxY9LkyEqjMbFCJEMrFrJJrcjRAdVI1Vyrwou0aJAybqk6XD6+N3rwj2/U4ORc
kUEk4VlcBib8vzNq8VLrHvAmSFp5dVZTOErM00+hElnTgqUm+fb/ypWvhRFpGR52G4kMWqh3Sb0c
fIp/F5AwEjUDgDWh2R2vA0WM4JYk+AeS7rXSon26ZszvgZtVJFrQU8+mqTzdK7TTzrL6hIBcFS17
+RQIWennDSG8ARAgOIAKVzBLe54ZdLR4Z8mNZBqj8i/pPX7cWOnK6OaQPXWs3bzbYjL4SurQo9Gj
7uHkrdH3sjK4R/iMZAlZ7Fps6q3ESryXb19sIGxAtYAMK0vjLR+ycKoQCE95EqnIJ4VB0Z+fZfkG
zkvr09aFLNgRhxFEv+ynKyJ8Sg21WswtxgQ2OAlvOvqJEZQp1UVT8HN7wBveK3lpzTyL5J5sM29L
cWZiRzZwN1LhYIjrzwveLpY+YjQCpQPZFGISdUtnXohA3o0di7Y2ET7v6+FfLcZxbnoRKLvMwlDB
lUTMSw4KVdFOKw52qyHSuAdxo3j3aelObReXJ4JzJZ7gkooihLZpTDuVbOprkmGq8K37LczI2AxK
NEBw+eiHXPFO+JR+eLB40+aJDquwd2le0QGNFBheoSNzyrafAgOaJTfN/2ZDHo6Y0R9l9FstDEPK
KawraVav234z40/8T+BVFwq1BQXOwLcKzRM33KPaxfG2ZVZzJexxTz469/dxjR9lmysC07mI+pYu
dklWv6C6OB8FFj//qFlMVu4Cp4xSgstgc1L2qSYjCg+kIOuqTIJmKIcMWbm6leBe8FhZeeIdntC7
8RUX6K/3MgGd80GTRtrIA21kt/6Gc2kyREWdDK2bzgqrwPtJSyK1wYiudKx40HpepcH5THyRnrNj
pqzjEGXk86pmBW3ROIPlbpmtZYggAOHECsojds3QdlYsTv/PZHE9gy7JAzQ1wh+ptWSwsy6KQEJA
RXRvC5t9wJEBJbk1aEo5/8l+CATZV1bIEiMs2yWrjB/G5anSI6khRwmfgZxRDXPTULlECFkO7WoE
cdom5gtIfJvN+AdscFz2+dKx/OQdSOeXpSEAVl5GxXkiHvmYERwypeX50lXWrRYm/FnbIgQ1J2vC
VN7J7JlBwtOYtU8Ds6AXIvmOMOckrUZXmelgj4EHPKO7SOemmee84ID8S29ivHZt+EPonvGOyvDi
3njzhjI3djB5EAPRc6kcqk8EeJJESLZdg1UtxEKkqRvhsj59lG30FvARBlj7qtEp305Ribxlgwmy
lDoDv8Y0U4/IUDud3jyDBafH98TYeqN7UFOHyWqcNRyU418oP6YL5QFdZvVQOQc8Es82zF/d43g7
W1NXZinMOtGVm+BmXkwCgov7NwVD2EuRosEhgApEu5CXyrfn3+vZafR5mNOBczp34cJovdC2hpJi
gj0CesNGm3FUtnx56h71drVqppc5bT8HYRb1sz+jL1loYt2GHQr1npLADZFY8jNZZlG9k1Z1LAgf
sd0knM6l2rIebbXkMewV4KudRcnuqnz8ywVr7MB5GjxnYwcXcL6NraeZbtpnHFFtCPjiom/Q0F7x
g7ywR+b3qUxeaTWpIy7ITG0iChPs+Dq4LSMk93PcU60BBMiQXbg3me/gS+MXFWCbPCy7tCQ2ZEEM
7kfIds1Ya6RTF4f/S5A+0Y1lYdU/zP3se2nvHvMgB4rN6+wc8rypnpyQLPo40fv4QuElLFQMhpQf
xSsF7KUyAwwpM2fARgRSTn7+KVYzvfK99tWWj4G5e/sKC3vSp8zb+Ye6ta1XIpWbHzxsfJe8pSG0
StKHnQvOl1vEz1s6F6z05kITE+GXulTHVZnxZos33EACxsAm6rkdV6Rum5c+ZTCn4PjkIyVOkHQR
UnjHEYfcAGb7/kIlKo9gcgHHPqaFOC3yYBHHEP4B5TfEB6V84sWKm5mgYbrCs/BU81asz+ji5B4x
tCOeCjgCntuPdmGcB5mr48gtEcAEsrlLDmI6tJRqFm+0jek981M3/4xCc2VfCzPDGjIIG+6UVDA8
SD2Tjl1RzxhhlBe7IgtXuC+Dn4V9so9CKAjuv92rr6Mo0fXj2S3fVitDsyyCtQVQbx2t5IjjkIyV
53XMg6EsM8P6YYWRxtEsMR7BJ/USyyjPivs9VYqfHka/zyyGxq2gmTFXiwtVBLQ72acNrZ8NSMEN
0pQp7RHAT4kzrw59NMhXXPDB8/fXxP9wxm8EybyoBFyiYU79vHKJzvlBn0XAZ2mTYKerSQhlH2fH
5WV85qIKNq7gZk7+PLik8kTNyIYlbV2pULUWM3Z3Mo0TvMmlI3AV2RYrDjLezpJ1X9prpUTLEGj7
uxFUG2rNlkN7ey4N6uB+IeNgyGfAI3U8jH8+mq+06FG2HU4ZWOKrI/erVNHaJV+UG4MioCK/qV+X
l2WhgpuWKPL4KvYkRvLCjPdvkFkfsjL2yWn/AyDWgOuc7zGIk3/aSImyfQ3Nh2QHCCe1o0iADkJ5
rQD7ZTuyHJ+B3naMX8GUJz7KjArRIXAlyTSHGPtOYrIJVEADzab0hB3rF4RyPcnm8E5y0QFrUX5g
qx6uK6Db2X1oyirPAbLzDYsLIJ3W/xn1IcINe710HXFRqYb9615yizlN1ZE7PDzo0KefcHjmomQk
x+UQUySWMCSIK/BgXPRV8VtTGz+nWT2Hsdq+TKlUDwn1A0qxgyBQJDAU5ZVMHgZtCe8Gb0HqKaDS
VWkhqelbepAiU722130u86WQ9Wy68RzPz+nJPvPqZD2OygHtSDQXrSpJye3nhIAqjA31y6S6iPyq
fE6pommgYUeD1Zvy7ubpJLXkp5KBKig2Nt2XQ9+hoBst1OIa0Ri7OfheMp7bKOuKjGXt6+RMIVJC
GlGngLZEN+W+eF2KnDCtR80ybX+nCYLmdW9+hBY1G53O7A26mQTt/1OpUcvWnhYLcaJzttyj7Fh8
x12gvo22fdM9kJpS1E7mvsBT93C+Q6nxkftKvh6eD1PL2K8QurzgE4njYweVdKEIwV8Vn5cahJXv
SnRxqBJQun2K1M2AKqVqQfDOK8TvPR1Ul18bxBif3KCYe0iJyUl2k5thXCnaiCWmpuL98o0Rlsze
o8SdX+10puBn2vFJ0oWljdVpj2EQzLUxJytJREbTCqT9v5MTdPiTMTlWRZ4hRWPamyue2m9AX8cB
cmltfBUNbccfjvIaX8haqp4f/Pz4ifQSD13rOiX926B4SzIxERcQJDJx9JpiHfJ2NQoGtTkU/S2A
dOgc8JXIzBeiGsb3RDuggrcG0k+wVcJ0kiOgkDSpJi3gPl2sVdBURGju8fdRUIfG6L6Y7ajrJmp6
iwZelLP5pNy38InOJlugGUP28PJwWS0e2iBZowMGzwZdVBeDNjMZfmgJXKE5N0VaucADe3bilI5Z
UbvhH0CZVqJFFTqiJGte+HpTVg81f+9COgw40DU7N30QE3i23IDpnTtu2GPl6k4MRC9ktOIiFpKC
b3j73GiMEtWQXe2h3n2yJzfUsXxkXqzvriyJFTE/pHgc9lhT7yKMnI6Vx3zIeTR36x6HLXOGxlRn
MjZ1ENyjxfPs1n0DNNciDslenBP4hRIb7Njpkd7qnK8UvAoRIpErp418ygl0WC70Mp19xxB8acJW
DgAOz4JSOt68noOwGuWp/L7shNcoFVjSyDzLzanDXqZHn/c6LQWoO/m2g1o11PDZ+AhLePSC1N7g
JHItaNh+719HYhVKkrzd53aU5JvteA+lCK2pAUAHqgfYbk43JUiQl9/7idj3YSRKamSVs5PYnY0n
EFrgJfvBbMDc5NTjvCr2hHkYEyvdS02Q4mLEV+c9CtTWn6R0XntodJKDh5mc+HOuy5ZPHTBpQ5Qx
Fk+bGXqSYoDtsNMQ3JrokNj3XkQJN5REB1tkQLUdTibJJBVcfo3EXorpEoK1ZMPOHXKPiAoLwDj+
DfNUwesA7G29S3fk3bgRBDZYnOovRvcy4h1+1QcX2MWj+8tdoX1Qd93YugpY0MmFVngHv317q9Uk
5qy6bHmNRbefcmlhmusN1vsu/SNL+Is/sWnOtiO074xAxCA2Zv1OvtVu1ltV8fiiw+w3VWzEHCab
ZdEsJJznZ08c5KxKhpOmaIicmjfL1V/0XI8As1jnLkKWEHJ2hjcDed21IdT0FIlXZhSwtfG+ipOt
7r+KLo/t/ahqmaJhRBFzSpADSLBj50hbTZku2Rm0pRv9DwCKDL04o47eDOZG3h2to69sz1/Ki2Dr
hiFr8QGHvUahd0oxvALYlEKUsgUm2SEoU8hYR7cpoFb7bVL40t1Gzz7Bqnv9BVHBYxe/U4MEY7oT
SqX6tyh9tnO1nzWG43+hLdAd6h4j+k/M6N7KcuvB0YInzMzpa1cD6Bmt9dt0wNZv4p4sIlqp7n3b
F0T9/li7XqEFaGOmJar23fbbM/KdSvf4p2DjpoyKF6EnQwDP70ca3unRoiP1Br+GV9fSkA+3+agy
D7s7Ro4M33n7Sod0RTWq7cCP+GuxlRYkP8z94AvUI2tdgYYhKQwbWvjOPsKBY1VxzRqJoSfEEjo/
e2p8vHTzySXmOHKCFLAb18z1c/US3YDBmrhtpykldWaOkaOYm1dp5FQ2Og0uiD80iNdQbE46xU0k
9fRLQqOoCL2rpwwJeMwXdG2MddBmlvSa4bh6neIiR/oZsI1+WJSQT9ebYDoAS/Kb/JOtYUmlnB/W
2Z/qA3qwvKuw50h9EIBdkG7qeAI1gm2r7SImwOpZ8ryfjQLZ9Fl6PUAGIdlXDxmcq/SB6QoZjRn+
ZghCPiybqbb2hoZbTDkf+4ZlqakzgTpRxzJvUbFfY78eMqCJ66slqgZxFcnnSN7zzYwOQWwfXkyn
NaCC/H70wEk8qDW5ypHb78aYoNHH/lY5kiQYj8rP57i+g1ump0rNqO+0+UtyrBZOhSajOLVOE/5n
mAabTIhzmX2R21a9hxCcfKxs4sQbRJT6TJ3ipU3exbrV8dPxYVdSBLlKmWqGQd5K79hbull9Xkf1
hk1hCrBAxU/WtfVzJI1/k1kMYBh7h++hRKOHoRFRnKxth5ZQDP1sc3+XX5QOCM3ai1JA3csu5lE9
layqaPa9XV9APYjlNxZDBmZp/QStVZ5trRyD0+u9MgA/S/oT5sMOrnjxcC/Ce6zew2CqPXIJJzH4
uTAI5XtuZWWGE2cawKhhmcLAYe+iiRBEjGHoG4fDWmJ5oAlhzH3buu8T1r4Vd2/R0B2CGU+nz9uH
fGHYcmdgGDZqkP6jCl7bhNJKGjjeUJJ9qGuH5GWzC6JEK8wXQruFD7V1vDnpUCBFVzycidBV5CHW
q2pLMH85UeO0qKfg1yfyRO5h2vGflcq5PkbVUbglgKh+ixL5mTlIs3aUew/K3Ltd5JO4E2u+tdRf
pxXVylBJmbkYi1rniLx9evxFfvDx+dxLnHwRqIQ4nPcT7V1CuE9Ik8PcV1LfHoHnstLME9Js1Z6G
mVMCtm7PjylF37EY42/n09bVNjyHeJ2d/XVBXD0cSWWR0MleXWLeL5VQw3FkVwDZwwrcvcbW/OGu
nDbNsqpsWZS4OAOJ+1vyPT7hkpnu2M01mpW+qLtvBFk1jYPNRCSuX2lIEYsAhFcxhZgDCtb0YYT9
lsTvbnmNfORtGfPQP0VfS+sDdjI0EF0lJ5HofrdTPNQ7GeHfaJ/7lOQMh3cKYMZ2QDtcJF5DBiUO
2cagRbUqQolKWGzZ9OAHLUgo34OqtNo0bbo7vylEBzCIMgENypMGuo8oge2ljPls4mJbFy7G5HG7
imYrOCiteT9LjhHMSiOSJckpfnZUrF/e+mgkEHgvLh79rnLMwYADNJu9/T7Ehwu80ZVwPbK8kt1Q
9lX9qrz6IEdnsAKDmUTu+vIXv60jDAh7byzWaoH4f9DvcMEmVzASJ6wF2o+WoaMLJLonfA9AYink
Cd7G31B3jq1lH3lGx6KEXkyiLgeggad4sg56Vze8/eu/sE3hCxizbNyjU+9x72Ksmv3qqnBj10rn
SEicbSTFrwD1kdi4xzom8DESfoyvQIhe5KNoVblK4VzbvAzJ8GdgN7mS2ZsNnYWwa3WLSxkVZmjO
SWjWa5FxhEx7hb7RxWwOeqIWAdsHvTEQHSoll3ZYZ1mTrjbt3kDc9ZQesznUvPbwPAsrsZ12bw0g
AprjNLHv5t08cOtO3iwTB4wiXsfihHlt3mAhNP5I4hV8A1KfK6zp1kZfAQ4ZslwUDygO49SMFPMp
vomJxFQCq5VyOj57SDX3q+wHSECDxrzz6VuVT1ctqxEDdGg+41iNvtUUXfniVYa+oIULI4A/v9Ao
6kyyyuEuZNWvPIVfTQrPLkOjV9AMQ4MizXwMp7sW1wchh+6Q52BoWIuK8IiWVVYaX0fOGEWazd3F
UYeK9FuBsenTRXlWhnKIU3/2bcK+P4b3yVwD/BICF/tCvmhvkBhuEcxKbD26wM+YvrVmop3Qw7AJ
OvxjbmfR2ar6tJv6Puwe6aKcJ2qiXFiEDOqpkpOXG8aJNCBp69qwLy+BEDadCrnsuvuRerFmQe5W
YdKASTxRZ5mGt3KmssY7JVQrbz51HzXr+3QrgzvLxfv/YEXApPQmUiRDEo+sKxK0EUjvQzyIJ0iu
E+jS9QrGi5aB0Hr5EAOUlK3mhhYz9EQ2oClwGKVXe9ipZU8UppjaD7BDEZ/cAIPsd67Kc4D6JqlY
OcEhbJwOSKqiS3WIckxNyocCoxlPsMfTGXxXSoVr7IXafEliy1Tb0I9bZxWHpDZSUv59CxcEbxwy
F7v5o4c/mM1i+tcVnnlbNpYztHgwzpeeipf5xMEVuyn29/7H+TY4Axuca5fT2UBpVjlBTc37yEDz
DWO3mghWdKmmACfgNMkQiYJfcEBVPINCH9aR7PeWHQhI3xF6BCetLVz7clxuJR1uNWsV2u1IwBFU
9t6mRKsgEf+T+3nePE+plgCriUsgBuiW7TvwULXJowT1YauiKRVbxjCGHSzWV8EtisUxKgsWuSrP
2gpf2dXtvLLb+SOED5cls1hqjCM+1Ng9h7BZ3FlvG0R5pRw/WfTJz1k942CgElkpi2PTV++EfcCC
7LBq4htS5/LlGVYaOkl5aoodqJ62oLGK3svyTik4buDSEm0vlhJVpaPAuUHfIolGkWbNZiSwc13k
8qTVHRm08z3qtqC8B8uG6vBd7hCdyzLp/xiCz56PURROCplGGUloGs027cWNW4YurVrvZbDrhBET
2zSBSxB/ULkCAlBmah2xBarsG2kSCti9bCT4GkykKcHrz8bY/9czpbYvxskzlLPTvbopbKsejcnr
Zh8eHEFhvojQzpkQL+pB8cbeayKozSwuYev0f+7ujlXJABaX7TITR9CELQCLtx4B2zN9btu47Kyd
msE0+BcBVmVGUv5hnOsBywvFFtgYUntWgWp36sDrOY2L/oRJhW22Vq5trxvzJRhKAJeOSHLMMLMc
KchZ0vcnFShf7JPmiXMAiQRPcW/IoIAwtMH2eKTjflGTDx00ZL8EloKQIv4vxmPbLP+hEgkYSlig
2PavUNw8v69AnzEo7wqpRUxWQL7XZ+Ca/Y/Lhob8FN74/1HTlv0uzUUiYJgoGpWmQIBA5CNuUWsA
8PRLdB6Gz+g7U23Lt1VZmpi7n+20l7GIJE3URVoJdyUAnUW1sEaWQJWf5qskWQ5gtQAzN6s/zmMC
/xmnMiJiHwYefbLtWev4POhfWqBljplkwZAtP5MV9mScyG9XFe9My4i5L99M3D8/2APomIgWRtjc
fRj19R6SrhDC5fmWeT6Low27weZmsMGT6GRyYtMedhoxDh0JKXpMpwSZx6eCCu30OsIz76OucEfI
3iECY3jFlW7eFtr1BaKrNL2bT6HMN4amMs4K9kZngczY870uoNPP4LefUbG/+MMVunIr290FHDVD
pEZHbw8RFFPr2U0lycsx3n0R0PtmYO5CNYQ1+muzOI/CnG1areX1IdJh3heB83+TDhubKtsJP1gC
7DhdyhFVXiayVgvP9pGRJRQ6TUHBS+g57TBhywOUwcnIPBlKqDN4JjQcIJWgSYZ9iJ4zD6eFTJQu
/Akkf0DdumPgrOHbWyR8Nk/QM/rpAnhuX83FmEpxw0UCSdS4vCdOWL0XjCTt9AzhM3cabRs4IT/a
G8lN206GmR3rwQ/PV0FWOg1vieksmTyM661agAveigvvpvdZ9f/CiSNm5VcOyZEap+yPwz077TCf
w3yPCOlrhRTpKMijfI48j4YHJGn3NADoR5TBjEan7BnZAvf7NJvGXhsvlkmC5CmJYLrwll1O0spz
vBaaCRA8gPDv39KRAiolYvZ0E9jqCyD9Xci1IVwDgS3BbX/X4rHIOvDxz6/5IEgwGuFcCZU1elRJ
ywD26LkiIYk+OuX9t28taYo7mLO/EkNcj/vCcv6QxONA7oA3Zh2lfRQh0YPaKjBdoH6cgyAQYDL0
73GPmVqZwHNeVwlPi4LUBnybMdp39o7AcVJ8l1fyl7SxjBLHrtunQX1v6RxYrS6WWucd0C4hjZ0I
Po8KIsNM6cEJJLq4lHHwfYSaTiaFKYMbi4vEsxIYI9eZEJTHTHucZjD9HGURF+RtGN1vlwnIa3t3
zgvB97tYmL3ttDnzmgFGLRBmJBj0J8icURd/ZtzmACkLciyUSs7qIthYTS9kGzw4/U9Z2X+EVAu3
L0cHbh6vtjnrSNJmZiML7CbEpyKecv+ZrEHjbSc2RdXghmaWrPbIQ7hhILnkmkVK6pCedJMOW3br
XMPNJ29+slkbyMAT9H/y1M4v4ii0JkqFAQMHLNKgYi5ILG+4dGIqXjhXG6f3781T+fBYaIZG3/IO
m2HXZI1C0pTxtc+/sqhwrylABTN4KdUfUpIsXZ/yUO91NmQsfL9+ZjmyNIumugCt/nqJhvJ/NyUn
rF7yf8HEnqR+zIXN8MXEMm+XuRljQPByg1ongJs8eRtMxk61AcAVCbVDWc6j2Fo31aTJbpwL3Obf
yP0FHoQL1ZgKvh4e3EjehDk17uDpkV9DJ0jfW5zmKdnKrAMFJiUCmvd32DGUK/p4NlQGOvSrkUrR
YV+LznKfZDr5CWAiQOmxpt8ACeyBdHPRg0x2hd+BsNLXzz59+x0J+STk4FwUTztwH5W12XUt5rKH
NJwLy8ozWY6pRt3zEBCa/SdjIm8e88Rwj3ZNRHtxMGbkVjbZg6V9hENzgCJ0g4qx1oICa6y/QRTA
RXGeE+o600U9Vbzwybu3WgXzAptRkTE8iE7GgDp1TwA4+p4RLUDGY7Fi2mWiDLEAhc/Mokwl8Spw
HF793XX4N7HZchAeUslLjYtjZABImLb/tNySRZM3qS0VW04VBYg8d0G5PORU5LvaKNDTwYhAAtZs
EG8YfmO818GBPHE3SOStKAEm+JkNh9YcXqz+OCopW7rk2ILo/P13SwD/I5f6G0+188VBjrO4PsBx
1LIlHanIpysmHHZ+ThwtvD8oce5uPmYIPukTqK7o0QfnEqNF2YjHc1cfOiSFdNGQpVh5JEJBOzya
3Pf3xngF4tFLKoSO4sR++cgbU5DRHhJmfYBy1gWIOZ3JBfndfg8Q9gv2URdEkYIKI+Yrv8anGC73
6lnkMwuaKVvw1x/gVHNgEtQq4HcgcKJkcK4NQm9ci5BDnawHiHONwPlldPOLQH5FdiSNFV/dm5uu
tn+IgEA13h+8TK2Y2AF9i+w4RDRW6vqPCrUjIoodrIi31buMbVd5Q1wWBFmyWxZeiN3OwcjOLLXG
m+/1u95amOeQ6A3aSnEZr+KTJb/+8wHz09xia6jS7PSpIHxDDHy/1y2AIctQPMviqgOjFwKEBb60
/QKS/Ox3SLBQFF6nL1nd6WylXQ8ZgBM7p079Kr0eCvCVfFu/UDIgzCzWG9Xbli03RCPW4Dk/llZ2
ko/dpvFLvGDsDw3Apq3wkCqCwFHEgl3kBEqDpXIr8TdMGwVrZd0oGmxhla/LniFZLZe2fZiluSfn
ic2stY72WVygUPJHX6wNMaBT7vGfER3VB7yWHQzqeZlA+T7GcL6ACM/H9enZ6P543fIMBYdxle8Z
v/UH8hByGQ6UV9BmBwfcwUzW2ZvHP4hpqymTYvTcIhscbHYqzsytT2Ppg7AWlCRe9viSVuNNbdPp
LAQmbBNEiUi9dU5Yk9GmaDrPwSPX8xVLTe0Mmas1VRS9Bvz/BTB+GxcoVY+WkBbY+hZWgudiyDZa
DSPtTjTpc+HmhE1S0lEbLBcNWgp6A9efvP9J8CuHXgrTy7c1iGVTauG8iCVIyS2S6a7FR3Red4x1
lQJG28gnd95F+Kl3A0oqiIQ4l1AZdw0utX09QZA4qTEzCVh9UwmPC+mXUxA83CRg/WmB0o2QpV+U
8hwobeghOAgu85zHjgPwXl7CMx5YdjQxQfUZ4ju+0IvFIW1TETwqsxOvCRhDiKd9yxjvrEWbmQep
XzVS7iHZV951SJeVnxGdFbhhMuII1mRWV/44wlq/MrgA4pfpRNk3EPXbPPJabAdjgn7M9vJ1EBks
4XF53naKAISTE/7/r7PjtKa/MpdT87keKnD8oQEjcJCU23btS+0tvZRueil11dMKCUKbC3ptiL13
19AETZcZUW7nHbF4TzWTGQPk99QCfQElBMtKfFPI22O4PpOup1p6vCccueyQVff3UDBRJZJIpaTK
IsO/UlrahtFWWtyyaMyiDXQmB/IGJxLjjO0RM3/ByCQeS3SQMM9L5lJn7TdpUfJcfS2CwtnQXsDA
D/jOOiOVXXlNKl+dCMAT4ylLXqEvT/dx2Vif4xI4tj+SFyT2mkMbH2Gguz9JPwuYIc7WV5ChttDx
4paqKSGi7R20/MLj0zhi7nBh5MXzMGsPK4m8OltvOj/lujV7AvIV5HmuMe2ePv81ORuzr+NJpIPt
b+jkGBnvx6JeJRe0e/rXoDwq0eO/BE1Q/QcckhEl3oGYX4t0hwC93+nI2CRN18W+0pBE045WZrGr
iNTv/DWQuxcWS1/3tBXbGIPZIuIDjTrR18Jj0SuoxmiqN6qIvKa0dQZjiReJT74rH5M3eyj85dzn
pk9joOYuONmbPN3f5lx5BLq9ixi3OJ1j3LrqQw40ptQooWIVQoq4RHgh7egX7zVXztHCR5tqV1kj
NBhtsYljBYnmRZrkp8DBDxpMi2+lnUwiO3a1Hu+qU5n/cPY/Vi8UovMnymyn6DQtiQNaFuewAvXg
gWTAObniOWQF6dO42n0f4+aL4pIJWoJlTWiWXH71J6HsxK5rbiRjhByGoBLXFrIvkO3oJ4LkYBd/
R3iqslpRxJgJEHGB6ZLxzEL7rZKZC24M74F/8uJeAJXO8g10RuQkywLJJLb9Bu+5gTNHCmzMeIxp
WD9268y65M4DET884+43S4sn5xQHTMcYSYDxFR9DUIdnjoDVCiLP5T2xiRvKN9BLaAgLuQSi0ANS
dSaGLvwXMpVjcYH2oKLuogxeqyj2ysDtcI7XjnCizzFUAq1nVpbNf/YqlrfTNwS3WklLTFTGkV47
fYxgZLp31nCySKfN5PoD0lyXmZn7AepoVqh5r0GjtLsFu1RoSaRC155PBMkdDZuMS29y5ARKvbFO
ljEgP5lwx6ZCevL0/z/NwBCpTy7aypju1XQ/6P2njPFqeouXTsTQBp2Orjv84AoW6+MJFT6R0kA8
fjGRQ7qA3pAqpyB0tLlgLl38TmldA2jo+T75nEZSGhvY8Jdo4OHwOspClzzGjKJw/aOVCuSbJoj0
IDLGYzlm35mPWBYtpgzVIr/0anFS6UhtSIyp/23DMevKqcuCcnw/rpDoDeWYuzpz7tSiqE1/K8Tw
1TFbcHa3yWuLNlt2jyce3nrCkpslnIH/Ivz0S+fiuUxTAhKw1WC5uCm2D0eL2OterKZx7PuYWQs0
ioGD2EHNGct4TSKAayKK9yjKrHQAMDpZar3Z2kviYM/JWHuIbcZ9bqIHO6x6GLgJQnzuyfJw35Zc
KL1KTSew0KRK/qg/NJCNU7rGQZ6GnunraCdr30Orr0AdX3v0NocT0GLdutDTXso7EY3Y4Qs1p0t6
MYpf2Q3YHis67WsS8cT6BqYaaKMkv38V3B7amMJVsRQMbVPU8fYoI2GSsstg6H1n8iOuV0gpH34N
5xvc8LVXANdQw34/iRcdIbBJkrk8i8evDSSdkzwv0Do1vH9UhWgb9FFMDvsaYz95bC9SaqQqexwW
XzNH/7Ox+h8zL4jpk+rgiYOAXhoKI3Fb50G5tsZTFTpyAfurgEWQbthDQ7cQMUYOI7kbh44IprBC
n0n5eK5xQ0Mdw7RhyMIjwIFVwY1Y2sA+08LUFjWsiLnp0xVw2u8XfUXtxOSImfy8++Yl+Ixqvxa7
BdIuoZFkvWiOK1EuDlr5LW9rdeEJ5bgs5waE7rlfISecv9RI0czjVpTLVuQ/z6tZOhF4Jpqs7TnJ
FUkzPFMIC3Hjs19AGLS/xJT98dk9CKqcmvs+qZqExJLhylSOkQQzkHTYpm6HDzJeoDqjp66F2rpX
zNsPPoB5wkCBkVnGrIk/7nv8lM9rb0yFM4r88g7T6Z7L80ETHoNgJG5H25upztyLBJlI54BmoFcu
5BfatCFCnTgFXC+46IC0/IpBR7E5pDd/63OH7G6zyWqEudDsYObI/UFHDCXKZIPDPybiMhQ2RarN
j8bGE8fp+/WMz4366togBqHoQ4RKlU56olsnPyrq08UxHOzqfxVFozeRv2dYQX2AP4Hu37RionNo
IsDrz+3SoTnrpsPfHYhTmuP7I1CosGI104tx3gtYehPCt774XDjxJzH76BuB2NSf6SKBaTrKXVdO
wjBPQIR4lT2sLJmkZl7JekTdG0MhuswwOZpXOyiiW228ozYpFkGQtsckj+D7QEODV9JRUltyofxm
X5dfco3TFb32+p8ycCO1BvfjJ0BQX6yDxo6hHBo59+KnlVcsakNSHheb6kBel4vaFn9JYYouh9+2
FOn6gpi/UbRurbFqUQ9019ciyFefdePWu4csMqFKe6J85IzCivlpXkQsdZwJT3S/wKjW1mXanhsr
ZBjXLBw289ZxH81E46Qciigy35Brw0xhKYROoGq42WP7ijxrPWsKWeOpBoqzGiJCcKg5GLX1DLSJ
8bYRkqnzan/g+6IJJEUGMw+QnWIf7duZUk4LuBAEl4xRhtXFXrgYaVFJzzm0+53ueCghDdFcPDDX
HQRvL8tPmgwcDB3bnC0dWhJTVfjDe9wiJchwm3sZS6YJ+HNOlpwlizd7katEQ3JliM9icLcRrNtK
fl2Wqh/KC5M57J8qT8l7sWH7j7cGmogVMjEPaei0jGvR0F+hn7wwZs3uoPaGWzKn6Z/td+l6PhRd
IOj1DU8uSTI8B84kLrHh9feBeDRi7oYWcfe31b9BjMERrfAYKCyhuA41TfiVB4v8ZWvIclHiPUl4
QYxUjPGKmhBrP/oWGS0WMi0YzvA36wu5BJjnnfHUdDNMG6koIc/dpp3ev3xgzb2wPqGTLA+3USP2
DDrGfgMVawCaUGjK2DxFanLEYUfpEt2OnrYSRqJbI4Lg7Mafjqi4or9nFAXDq8/Dkm+lp1CbNEiD
tqkL0y0X3cu7NaWgrBamp14T0uYX6CeBXOFOGBBdQh8Btyd60arAuC5LmvLXqRrjT/iELz8qLWFi
zRmwgPcfOOFc8L4u0RrngiGzTxKR+A2nCKAhe6A7h8iT8KQMnFi6XxJnDytnpF6fEAQaGc4JSt4G
rV7qUT+FduwToTyJG580latxb3b2YrZQoxMfOuOJYv5pw4SMwab8Gq1+trXLbEa82QNftVDLCmTZ
LhjfMqlm329kADkIewRzJQTgCQoi2N1PkcnT8DdrVZd32y3YmWV5OFIBeSybV7YB/UylCFU9ZEJR
Vj7vRprr9T7LejoKPD3+rXPR9kde/mCNB6PLeMKB15QANplleHWBt6YiyGJdv25FjdLkWy1PfJCz
1AFaPzOXz84exkBVOBlcTcMgQDL8anShv7MBOpMp1rTg5UH8PsBhEI1XrXjPxvS6R9TtPqDMLwv/
9o5jagXKzPC9cpmgoPQv9ipWBsqSA20y3Tw+Te46Y2c/WZIV9xNsevLPRXdti3dcOhodEUHpDQWD
VKbZpMHXaqczRE8DK5b3XTq/wOr0V/YandAkFn6u0zhRvQAYbcVfOd+QJHhlMU3kj5+XGBWgES+4
GtczICIAcfc15uxsWj6GFWNmbTRPmsSAAiwE3xc8dJyqLHhP8Aj0gQwjx7KrzO9IJLeokRtDk8IW
BW+PEHs4Dr8EAyAZZX75VmIaSBt3uSBAXHR8ueIq0095Qmrft50pTGEbD+CGY6JuStl3eVc5Nfos
vCOg9CGPIacYxoQPVwBW1Z16GTV2RypolQA1ZGXW3a0OD86NPDrrG6qSMjPEV1xUFVA8ewNGfkHp
qOPG4czdLa+FkhO/NmeVvuEuuenp4VB+6z8e/Mm/5qmbtZYPj+lXWLfkJirazHKxWkf3v2N8ufDx
akwPjhQaGptPbjjJvrH6RquTRkR6ExoQ3v4jE9xYWXERNZvOwLGf/25cE6p/fhKIWPGLnFL+5gBk
8hpTUYU00SSI8JuG+ZV6pZ7Jb3ovitAdwxUP0xXkmvN0baW18BbaANAC8VyDFhDAdRA1StR3p2Rs
zxmy/CEjGqlcVNYG4tDQ8WoSNsjZPhG41EGrPZpdKdImYqNG/EmO+sJxjOxXwIi92PtM07oWg80c
ctPc1HtRyxyFtgrcVAyx54WIHk0keOI93qSOFwnvcvZcUG5PeVCzWuFgleSRP5s2l6t4wv8L+UuV
Kp4pW1BXbRs5vhIKSQ9zfNQ4cGMRBfs27IFOlzx5lMTrdpJl/xTvJWQCZWuzxx2aWF2bw0EU+WgK
aRsUXm7uimq53q8tBAxhRNWKeUAi/+qHPmzK6noY8P0Bwo5oR1Kghr8XDqgLPGDJ5C/v5VRAOhU1
8iETUhs4BY2H7HVxfXCKUtwnlbKJNpGjl+u9zeBbGuzwmKvWnfMGzthtXzZaBL5Zr0KOGDBICMF5
hIZT6txh3lOqG0zPPgC8LsCxDt6Hvp6AP3vXgMr5jLxN2nVYDRtyoKn/Od8ye5Sa1eckJ4EtUkEx
fbhMpbF7rP1rQX87BQDoJAdmykAk9ihGtra7P9dcxe0LG43mq8jyJElvkG+4UXwTNl7g3XwzFU0E
0+Yyxk9xt7KgBsiUIzzLNwqeZiZ6l0vZlvm4w2eiTDRwHQoQbVrisPAFEx2N/qh29QgGBNbvsFGU
TcBMQgWPOgU29XHhrYYzVBF7uQ9aJbemdHxJx3Qw0A5YxXcGfxIdh07GZ9g62yYchvy+Br0GA6Eu
utWVjDe6lRBpGKipwgMsD8G5mz1tJ1i6L7FKHwJTkDD0Z8KqBKQY4CWLR4BUJWbj4wH9qbQi7+fD
yrIOO//rLZn6vsU70/HZytHXItS7iYcM8VL4R12NE4scbP00nMuO/m63j5N6IRol7yGpcrVqajBX
mQvIZg2mNc8NbtxX3GP9N0RchUcxLD/RddpOeA5qZX09BdhVCV18DhZNSvq/Cfp3za8JJS4Cuyis
FCld18nrFPn9iM7dhdv8MUU4YBtFTmN/1B7Q63gxiQYirYCWysqCtj1oH/pz1ZAb2iBDMgXZioVD
p0y9+8efI7bmPw7VeeP1fxwWxhP8fCtAcXKOCEVjVpVrvA43lUEoBAd/C2461xPUbe4+gJr8NEbt
mSU9AYkkWFh3REs3u5k7yrJ+5Rrd/gEClYmhU9StOZipdCZYkdRUkF33N4MOVFzzIW3G6ElPFBhn
zMLRffVVPupXhYFYGdB8IycZtVP38FwNHvCEzh77iNivPQrt1maIGDAYgvn+gFo12dQ2aZh6K3Eu
R0J6jVjEuSKQ0wKqRJMGjjLbTHfed3iKMS/t8wHFcVLaoUa99HU8PfeNOkHivRmDNGUX7oZc5+4F
gCjSp32JEFuGP02pZBjxMNkE2pC6H48Ag2e2+jaQG3lXQuSbEd8v4SI4t5yHc6AGw7ungMYdveO6
foCUbrZ2HFACcBT6hily1qkE5qcrLNmum4mkB0Rs5S/WX1tJ+37q1w7HgVwU3OhKhpAAIdZwI7rm
32bdD5w4j8Lz51o9ECytlUZ/vEfX/wN4uhXZZUkxWf2d5OLEp9zlB8ZI6/P7gXYY9lfM43x5WyC/
5ZFUyzDQ96BqBbydcHv9xWoHor2GJ16W4j9jWFVY51yIyGubM8w2QJhJmzaG+FN60an/GZoRdsV1
M2MieeLu2Waf9ydTrJQutWNnq+F9D5RT66ChnI/vz+3OSTTvSHkz4dASk+Xney3/qCV9VMFEQ/c0
u9fUIGr9CMg/BuVxhLZcfdC68X4+2BFzDsxUo+tWsv+NHBzaC0eog14BcMa3VrmXIbua9O5qaBiN
yVSxMtii3eHEjaC39G30c/32Rs6jP9AfPlEcO7L5rYSOw7I4JqMziNCFOtKPhomJlM145UlTtH65
MAQFgsq9YdeRSy0PzYAfUqBS6SrXRYiZwHT3vl0QFskwvrj1F58On49UhdUdJ4evuuWLaxj+qUfc
TfhwIDP8T/kVfP0sYAfOW4KM7w0hmxNLCfg33Vf47MGR0pbQqnuW4D85peuKYVWn22GjJ0iphKMP
d2GBTOgucw4p6t7PLmigVHKuO3YU712JR5YBNwGst4bzWU5XNc0AAIbVnzTW38OyuZEa/Ak6kgCQ
MTKAqo0NtV0OSff03zfUHzTKbFMMOkIfk9zOqvNsozFBgeY9aHcGtP/6sRj8Pk3pm/m/gQVy0hK4
Kiwvih2cLsskf37tofF1QZ3MrMNULNp6Q1V7CGmqjtJMUF7K/E5GVivCyYEgFt1xYNciHALQb0TG
pWfbF7XBPwwGRXB7cYawktgz6N/Y7D9J8+OS2XbtaigRQB68/4J5g/97v/oDvZIZW4lpeqlA6oeC
8s5M9JkK2YFPvnZv+zkGYzFls1CrryazsiGefTqXsOD9fgzNpxwhAmFG2KFFk4pvWLO6GcfaHF7X
8cLCE+gUmpDNw9yaaDQJJLJoIkoiproET/M5BK9flLFPaesDTXMdv0U0m2Ms06NfwxtKHAUo5hZo
GsD5VbdFSN97RMDGCYEXAzZLlIxqJueoqYJRpkX7fCgFfOU2bg2wsmQ5B8lWSFWHGMcEn/QlKduu
gxK7nWF3mDK6QJIeZ2vUqrukvj858BkAL3qORS4OY8UqdEv7ttw3yr5RTzMtybd2m9UfaFDd5Tu6
31+rsLLfJkhDIffmc2Cbk99fIzBkFDdkMHqxGPHhQe6iw3M06A4B4h0+LUwO1s6VBqxDzGYjBd9T
J9hnNtAmdv5UwULWdR/nHOPZflT7ERddsleP9e4YQta5qz6vERBJ38ioHT0J1zsyMn6hydWFu246
Gogr7Cg2mnwTAZapOgUD4+8TlJITfH7pQlSz3sG/5xDf+pFkKV58eEj3bJTYe0ZB3pT9lcHY7WhL
BL8I8hkg3NWQDFsNE5s00HTPhWg6VGaxXsjRQVOlAZpdpH/ooKHyMw2RWuuKyweT8OHoImzjvfP6
bR/lHF4Z5iyxFQifdWci0miQ+XsFnrQGEw8DB4LMCd18+VA6f8MHbTN41MkwWslF9ONFH9IXPqUP
WRa6/fFlMfBDiPJQcZuiGYgoGI2QqXgDOC1K1zLH4ouWcURq/VHuSQZZzV0j0WBs/73ntjXGE4N4
FJTRfQiouHicU+gy+xMlS3oBn22XIMT2+PRVJrlgY/qdDWuiKro58kRg0q6+/ZdGIlgvgC3Ri0yD
IKu1FIFn+r7ikgXK70Eh1qxXblbn3xe167Jf0znQwtuDdQgeZhg/TlFPRzqNGLC8ckxrq7Ljp6Q5
Nk+mYvuLkWaYIYWO6qxTr+S4j98FinKTDTIqRT+UthZhWy63ammibLlvddZgDfy1Ge4JxiuVa0Jv
imNk051k+WqwdZexbuSbjQn+dOLtrH2Nvi2ZKFWywAxZvqT9ExOu1a4GF1C1wm1HKF22iLhgvOZ8
6KHK57+Bo1F4h2QUp5LuSqukR72duq6hy0p9JtmrRpskTcWtYJcqOUMhLwXlATSt9F+RyLHvIx2f
oA1nsN2Z7KG8BPsS3vecs7bK/VQhWsjV/HhsaRYi2nZNdwjKLMXvTAH8bviet41GJUx+is9ePOV/
GRXIQJscsLN8qo1rBwAFCm0UHPIoda60Up5ngcyzPAQpBhsO2fBwOKVMKdLQJDWH3edjJknnhhwx
UMLIIOcKeO5MQp1au+rwV439ejyLcXbKtqktRtc5JGfP8OhGpUJ9todZd5C0Aa11hVgXtY0kXL20
ngWn5YkHnvPTWKcmPTSTqI7nN6r+U7AYeUfzv+TMwQcaD+NypT67n6w3Mgsq+XwRvHLwQOoM7dYC
fYpDRM0RW2XMRiG9vDo9QiJFICD6VcGiVLVybhABL5r/8aaDk2SQ6eOHD/pJLu5h6zuLljeg92A8
e1yPN+wUrVQVUrxoZ1UJ0NxLeAOVPoxJaIm8dfvKT5Lv/Szzrh30tiHlNrXbARxZsm0f27x5zNov
tALWd4f2fpUJP2uV1vvk+j37s4UnNEPIzTFad/zV8wWOZw8UQxnfbwd/6f9jugl+viGGasVKBmc+
kTrdbcCEyoRO2yE8FmokJIsQm2/7mafE9sHqLxwI8s6D00IigzPRoLXSJw+HwT0F7EdPTUDHd4fO
nlIR2rLV0a8AspDI0NTh58QdLOZYFyEUoV0rlA0z1SwwNRc+hJM5/MVWBVeFqoedxvfyrRxmvj8m
/EO7/X2XwPYDABGGGnnSgQcVE5I3d61cHNFDUksqx4XXElHvZlivo9b57xX4b18N1iSWRExGZo4O
U3XGGKBDzGbMxEoNX4nXxYQ3eI0VajCwOsBT4z8v1oBO51r9G1uSPV1ZEsfTeFizGh0OZnCH3yqP
awSbrvuW6D7hCYkKjVfM40nyGscmTgOJGoioKW2Znuy0a9dxcbEY3qmnEzeFSk8ka8XtYUEDEEFD
FPZ+NbBprZntwGCagwpBgwetkBPAp3/pzaDxLnX4oSvli//NCD0LwN+/ayZYsCUJIwbRKe+58xzq
Z0IJKCTXQ6KybSAhDXv78mF4WF/vkgvygDr9wZn6EAJjcLHUEwEgxDFkt8G1za2N8nYmcS3Crsfi
+F9kOb3QO7pZr9KWoy5JjLnVl3rVs7/8gJmLYQgotNVwNoF31mAC5Tx73JPA9shWCIAmsmNsLPdP
RQd6ZKWAeY+QKKYvsWaEPJCcapgUtr0n8x53Z8IxcKlvNNBm1VGT2Eh+PMCRyJdFgdetb/U24ZeY
iqOIDk6KJ2KOcMNn8DBuDiai0QZsmmj7oTaRRXszErLr83DDIc4VvbIdx/WA7/znReHIOITq47nB
iAq1M4p4bA7ofFeg2Y2iBQHkT+Z2vTgLftHMdQIUOdCdJ/TW+P9ufgx2alH2bHkoY6bIRXFye5fm
49NcJ0qkxxDIhobV1XfhbIYPoQOe7+YjDwtNAh0btuS2x/NTTW7xtJtMM38YF6of6q5SirAmPTOJ
+ssyenMQEAKGhQWbAeT+lY/zLExrDZbIbcnvlPsp0nvtKrkEzHtscLkxQLHun0TO6TgygdaFmeJm
d4481OFM1kgn/I4PGMJB3wZDl7ei5cJv2Dyjtri2vtt+vBsLHkPbTQ2QP9r1QrHF/RdseXk2zqgV
cdd622EZ7TpmVgrxJhGyHdavlOZ3d7AzvFMKGsp9jDusd2KLShYzj3RQAH5dOW6JZw1w4anvQEmh
sH/ffH7UviQAXNio8+jFLKi8sX/t6s/+Fzqsfe8cAnwozOCigONbacvxhnDq3PAeN4V50+w3pane
ncIWVduyxcCFipqb0LQOMHDjGF3+60CZPQmsBk9yaRfmtqxofB5UGWIbRE5Iajhs7X2Zu/HOcAKD
HkcGERjZyPHNoRo/EqBV5O91yiMWG7prIBt3lhZhs10ihk5UPpBqevmqGMqmRGcheV7b+p8aFlBt
xzDRkl0DQX9wSofU2ntekUizQhXqFrgxj+kef5wTVZBACTvJ7pmrjXzT26+s+1qfn7fk9RHjvdjr
2k/Mm8ZY5e/YZFD1sCBfe7loC+JsNZ8xylTBPAjy2UCvbE7XDb6WFMg5dWPTO9a6AjOHBhByzC0G
o3OAz9t/K223OnjwOcvBN+fnb2QUveAgDdbT2O/P7XnC9TR2ZZXJyBrstZ6xBDqayR5F4NjVHbJw
ThlwzPps4wsrxvbnMpIkX9mBhDDkNhQS6yN1j8HTEaIjI/mKncJqoUHAvE3DKrS56V6fiDnDHujP
Ud3HQ6pkw8dk8TX9tk933rQvv+rH/zi3Ys3yGG8Z2oIJc7TEu7+9epGLls9Gca/k1cmvoPBdiWzk
iWglyXX0cbPraE71v8o/+stdDPZqqIOwrAQqtxa/a3ezUecaiwSRB5f5TeSdRADieOrHtzy9C9co
Y8zPB1cBfuj2K/8b/jnWjp6IbGuS3Od8MYjTcxw2vPGvfJ7gf+IiNyr/iMJxTw7JHON7NlkjdjtP
9OplZvFkx6MNLEJ+vy5QBTf/aYZJU9BBOQ9dF4JUov67od/l/r68nYnVRU2t6Q8nOAaDRGCRVnOk
ixRHHh5gcSbcUqnBOmR5Y8VsxdEMJyaiy2P2nYW0XmvoT7CbIUBZr0jm5qW/9iRsMW8EDRnu+Fov
SyE1/48cwY4SSUvNU4BVlISBR9kfNPaoUp45IA4nmpILBNVsB23zx7P1t61Nr+X4iFs6/hyCF0Ge
fL75jBRobWJd/zcJXPdbVJkkv0NbX9ntJTUg5e9zAFQH/aCoK117k9CM0PN/n8B0RSb0pz479GTv
M6GuHy4gOU1o+tzaQqmsEgBfPqzKYJCSO+4SRRNXlniXkzs0kbssVB/A1hI0b/Q2BxdtLg0ljKg+
LWWrf3u49T+CPAslYvaUmxm1PXYo+Zx3OJs7meHWQ4DSL1rNJH1+TIT72tvU3FHiVTAnSN4i2Mov
kisIBQOMe7m/ViYV5uXKbi/M1bQkXbIgLBn8iwOxIq9/9koHJkm8StcyKVBkNOeJXwIRuNaDoKMX
/PurZ8R7JEAtdpmzOjHuQkWHBa2TXo/Uzaf1kxrKzVCA0cnDu46r2Br9/cEUZV5BsK9qPmBJJoYO
1ddW5ld2o61gHmNg+dT/uKKJD2DcNbbiOY0ldz05gTtUO7nrg8/tQJQLcb6zRuKQs0udGSEGDBDu
wtlcmE9pq2W1AZdww2+llNUN2VgcDYKXGkDt+8M8uZb28PgmP/LDphy1/k5DXIK57lrzAvbUYMXz
JU6Wo1QP66mOZS+ZuA8mr65AWd5ao+teVQMbn6l8SMFZucSEiCqi9gHGvAtGUzPNd49Bs/xakMGu
nRlA3WJJ1i5EH7X57fUAY8BXO8OfR1WYy3r9LjDsO7IWur4/EoNC4T3WAJgjVliig/PDoLBLuKjs
FB1RvTLUd6IWymVptgiA9xO4h0bmmoT+fibMmpCGyCaXbAoH2J+YE7qa3YXzViwMXYjzy8Ln/r/z
0Glbdh/Mz/po/UO4n+cGNLC4IBEUHkC4bKNAnqKW4VwEc7snV0flNw4htV8o3Y5DVxrD44AptAa5
dpHBjvXekkWkiyussKJ3DVLn5sxz1QHEbuGm1amgyR+RfQa0tUNkSPIbC4xQ+UsQqxIX6HWyOvkO
1VUVBCJpE2njaDmtx+OHed4OH0pIb16oL7XTzLXDzki5Nk1guwKY8YeIYGCnLR/EeqGCVEq2iU9v
qa2u4kVybJPOxuliZucSshbZIJvHrxKGhzY5yNyNRMVrYXlJtnV3TahUYZ+qV4dvav6b2hE4Gmrh
CK4Tvlwty4r25BvgoCv3pxhX0qGEhHfYAl08eyy5VhiORcN5ka6Mlo6Ur2IIEXbuzptZPWFa8hPW
sjSKneTexlxaAG0SU1by5JpPcWpTUP8kSDnDRXmV6qxpWctnHOrNuHermgeuHBPfBiiPF7g5gVhC
Yk1CNhA01MmzJZ8zptsHNO3xeY1vnnBsHdeLpLrzHfFrcmamUIaxR4P7rAk9hbA1t+NPt6hRDJxt
HiKD2MgJmtrowPseNBAqznIdENs9M17fkzA+RkTAAPWk0RTu2WEJ2VRTTtXlhXLLuTqzSg0Ai7Iu
sklFsiaXjUODPco73kPwxikGvrJwQZ+HXc0b9X6V4HgskjOyNuTwRBgC5s4w1ZwGf+H6wTGVA6EF
y7E/3PzNR3aczEhcuNhVrFO5xKBpi8ieW/bDG7oBonukFv/nROy8qFGW1MlAlO9LAkwlYFkwTscQ
2pBm7JzOZgqJbfxeqzavAFCC/TKFiSzZb21It/GLn9d8BNKEssPZZdOpub6A932yziYxGm3izkUx
p+EWeP4khH6GP7Xt4fkc62YKLYsS671z/n4X2LCtLSJzgBnbjYqfTk4oAJ0j5wKS9b6KAdXr9Ynk
n0Knha3kRjddWRaRUj7oL7JaEY5aq0pszZA8/EatjC2Di2sDHF9BfT/kdmFzrMO8aUGDxRsDv6GW
NBBfvWCXu3diDK1+RxGpJdMTLQn/oCVhHuzv92/PXzLDBvRRCj1EAK7vDlmWQrjt5qpBY76t1XqF
ekemiCnJJmRmtla3zG8IilSvnb4FOEbXC+PZg93RW63dRxVgF1YsHE4sqHkNbGtPl+9ar+V4gDqb
9K2EDWGAyMMf9jFWBhYrKriYARXxBJgtjQ6zta7rHJp5hmloJk26kHWk/QLSThcipek3vxaiUHD7
tNiNmuXIRCb39XQgIBr7DqgUAK6nGtzzzeRR+mIj8d+iS6QKJsygD0OQrCxh9sppeerljLkYxFgO
JfgoLmQ6oH+VapCN7XTGuRJe5167+1O/IMttBZXZM8A1Dbz5Q0NXUA56vg1KNUosXHBF6Q1JjVjg
plbmzCh0qjIGQYJhyNJEFRphlmt3EcsYkNL5o17vT6dHOTYjAS6ptQq2o7PURlLAWEDBQBjL2U+Q
C6gVq731GdZgRIX/vQ/NhdvnZvhB307Xk3bIr1dwdbnAeVG/FfyUSU0DmBfDo5TzMuP53Zrfuw+1
RYorACssXMV0AKgNMlRSbB7Vb4VT+ot+id+aRVskxZ7OvIW7xrmrKHMoaqRk3RPmyjgYKsSRe0Ly
rLdPWffIctNwdaxW8zeLepxkjYl3o0BYvlbPIbLkUiR2QDMfppvG8QtbxuSAO5xIFFA2J6q5txq5
PcnuoVZ+NbHrmIRUTSeMw5moPUs2rPSHcBpu5ni2UdL9lKkEbQBCP3DobaXBLdp6FuK1g0dvRy/O
stLOjci0yN3WAkkxywcwuowijPdxFPxEqB8TUURWaSi9CZRgTs5iblvqTEkXUpibkdYwXJ0aUCPi
dtah/eXn55JgKBJdv05ZXl6PwL6zf5uKKEx9iJr9dNdkDkfqlPm3A10afxFjaX5cDgCKngwTXIEz
aF5XoanHDbspzpHrpNcM89A0nyjFN2u8t05JF3mkvmxgj8t0D8bxGj2ETE6iQt56moDr7ByR3gL6
+Q+1633/5KGdrfVytxaaG0JaoUqtZE8qpb2t4kYb4JuRRPbwCsNkXdv4dIY7zJsI+vBHPQjlvbSS
ERlofP3j4VB/QZTh4ZMohZw2doHeNh6SuV/oLqD7MdGnsRcncvzlH2SPtARitEn0xL7TiZhAFhWW
9V0VjF8uA4vLHFM7saIhMoAOIwIwUCoZRtxLSUfTe/hc4UlW3zFyYkM9vfs7JhH7Y6daI9dRVv1m
PZVyStMVNVXkbqKxJNuw35jZYfuU2/g+irMiEZO7M6GLXx/Ja4quzDsJl2EgfUIffxVmVQw9l9Za
I4xj92S+RUjFQLh9z9CXk4+XzrmNO+KaaUv64oASeHicualCWhz0eE4qtNoxMvCkg2HPt5UT25fQ
iVxbN3Dnaaz4fQ61HnZ+4QII1Z7ZxVyLh6AtQOE3vL2CJZcJ0m+u3iI8/wETN48BRbJIZ1ObRXom
ZhYwRH83IzUvzdcTwcMckfNYHMy5u4xaL+lbHNIo6PgcTLisBiIV0ohOOrcJx2pwP4ay9e8EZgJr
BPe5fhGyYLsz2Eehegot8JqWbo7u1xl3oMOr4TwpudnyPrDztwnZe6hbWJ2zmziY4hwnVqYZ0RKp
wrrqkqwk8/jebRB4mBJq2AsgNVysG0qrjfSnDwb6/5era3bUczizToqdylo66HjAh1OuebDleynh
tOWYN21DaxwfiHm2Re4K1XFlqF/2TYi//2tSWl88bVKbIow3lFPY0stTNXjO6n+dklS3WSGmHboz
/yVPgYf4iRrIYhnwEdRlIb2pBCSsnBKtMDHNH6X9zPFcAonXYKwxJUwaT7LWDHUzfZPJd07iEfdm
hx7NSk4W0W9sMcUrEDCwtIV/adypwN5llDsEF1Tn49IKG2/XP3s5MDhtoKPa3Itd5zXaBDCfQO5y
kUXs6QCEu1N0R687LIQG0O9XPw/HjK7o+NKy64m6o+XZa93HenRFxXr0od/LO6paRBz2BxKmKfom
TfiJBTvJVDz0X4S7k8lBV99Pfx1dfMB7R171+BUKYDKQ0UyJOF+f4yqxKRCnvy+k2K7HiuRMGyyt
S7cKlStkzvnBrAp+tHNPcPw6tCooTlyd7RSC8KQ4uiQfsol/r5p4JSE3AK9sI5YyOxBrM7GtLWBE
kCdkJeHvpiTeNTRJ5ILLFgI5FBnVEo5zkj6yTCChY0CYZIawgod+fVLVxz/dN/2SEHdcAdIkwmFx
z09vYlluCJKualDOurDQPYmXMX+ZIRyNHTgqfoc741qOWcD9DpPl5IwrfAlqRDAuEP/0erGH8kOO
pjh0LWBzW2fZoxXseXlhjGGiTC3jP92+GDmzBuq2STJbT+pBEJK/6HEKZ/Z1Q7S2f93fpfecnJDL
XEG0ZITYBbqdrM2O0H9/OF2AlJhf5CLHPZNPAbSl7mT03DrgMKfG0sX1tR8WZAO162fgh908ZvFC
hhxvvIxiMbKMxmvjxWfphiRWipalOVIIM+MoJwR2rMYD2WWrTVLOjme/TiJqaoldpB2SWtxmqfoC
4/BbqLT3Q6iy/scVoUtk7j2OD63NfrS8BLNA+oZRmcyHUSOSR8f0Xq8+32mfunbNniRbGaGn4H8V
MU10yi5EfCTmnBk5s7wp74Tp+PNlv6mJZrhu89rjZeLMHtzbWU6qJBou3c5tD0fpbSaTOUD7GZRv
ewTiNeq1IP+GM5qRHnssEclqve3gEZh1fER5ohaTjtvKLEJyHMVh6VfIyy0On/Z9qye5Vq6kAEu4
mHUbQWiUJmYFdMqRmHVZzLH/11tRqD8/naLZHqH3r3CuMrOQxRamKczC71VCxXH+o5u3+HSMr2jn
b6ZBVnOB8RY63sumoWEnAwct4ZF32YFevR5tAlcH3snZUpHPjIi8MBZ/ipqt/kw+kYqxU458lH+G
29SF85eEJ36poZnE8qF2p+txcvBN4+MY7fjVRSIEoRTNc1SrZCJQ4rrD6zFn4T9RthjqxAwS0TpK
1nP7Ts4RD/glVAODgYF0IKF9Wj6FnxiHu1Lul66Ioc6rSfcGfGMKp2rWJTiGYRCkZFh3pcD1rTMT
4x5wiICpkIkBifEMay32K+BGIMWVMLkXuXJWQsStsAQiogZVwI0kd7/1GF+Yn/lMRf6N/o0kMyH4
BCAm/nA8GMb/Y5G+jGFGKUgK4y94PUHBgRxbqH4WB3yczBEIu63TpT3d/WYkpZBYKkDC/B2U8mvj
i8bVUACK1QvpIQ9cbBtE86UsnPtsJy0lME0FBZU1Oth9TJzhaRPSNvMNbgrz9Dy7aHcbA1I0fvVw
AlM+rIt3zxLKK9ksQJhkQgvRomlKLDMmxFFFynKp4KJ7wiSyzVjnNanuuBXo7lI3I0L5Vtz5c5t7
j0cGX6fPSxMGX/nudB2yDsy34JiU95/ltEWyXyBwIrxVqX5xBSuCahtiJDkFXhqJa4j01CldvnpV
TN+nBrASU5O3XeEytuYsme2ziOf0YmrQCoMR0UVldG3Mh0sRlFqGPpCj52aG17o4/HTKLKXi/PNN
97B6NBpWJDOYG50Cc/24LUmlJb/8Sgo9EqwRQ0dANvmy2DIXzoM3ebUIv7WwWfZdqc4qLemidhxH
Egy74Qx0xd7OUyg3kLolY8TelUpXy1LjYT3qgPobwkPJWByycKklBinZDBvgTQ6f+WAeHOzX9oyN
6Ay3J6bosMjhd9HmYAuo1vVFYkxG4rlF6xzQTK7eRqBhUmPjY3B8LcEfs85ntboleU9eU33a9f2L
/quGR6mefHoJEDUzOWJyDT9nQGSfhRJiTYZbhNHX+Rw3NEYHGJwvAMEITELwb7fZzG6TYVnvVvXJ
NmaDFpzLaWYSCT5nL/a5t1U/iWq5Kb1ZIipmnMNyv3hExBo/T8qAD33PJ2EyL1B6R9M7JG0t4wSC
GnTOrm8CLbjktuZQskBhrb57xHIKxnu5B01og+uVRVPxOqtNvv1pYEDUEc6z/38YuUWhXExAoIP1
RjokqjorgaUEwZD5stmk/DHzH1RsJp2cOpxYHvWd0lZQOsoEZf8Zar6FNOS8lLxdNBjYbVKy7JOV
4OEq2JjZRUqdkaHi6gd7U3OO4s5mhIoueSGyZMWTP5/0HXumbtyBagqPs7EasQjHD+G6tCFjqiF7
qxIsu90ZX09MfcKRPUZKiFlyhS3D3S591czf04Fug6QaoqdZVG27LF8hMjKE+c5a1B2tRvZaZ4bp
XHh0dCO7QQitrG1smEnbU50kng69guDVADVkWKoD5qYZeb4vApz2ipeoFDjWxQdgT8Wd/EGqtszq
+o32QH3u/eVTdmvEiM2lW2bDfWlUHeJcE+zneQ8TSQfPLuaoCm27P86XVdL9d9pDYJZuVvpdPo//
f29YH8j2KhG5mwQuVeOUZqpIFST4M5ZIldhBS6K1/Ra5bLgQbN7UXJmVzwD1ZpmwBigw/W8+p9jT
uK/6J47bhv+itinQs6gnKuY+NU7PAhZrVlz4S3RdQMs36HOc8lJ9yf1XklcE1sZM7qt+baZcpNnp
vctMZ4Uvctsq0bEURUdglsjNsu8PmHzteQV3bb5tyRbWDI7sj99hNrrjOXKhUuvWXcO+pca5YxnA
TshWFCHeu12jGqtvCIOoaC6/Hc4ts7zNodxK7j8jqRzuVeJSSZa8P+r5M1IvxAJhzKhpPX5XmHCp
I4cS4mgudy3rU7xjr2IxAlCgSPba3l0vWcb50p4AhohTBGS1eV2GqsvuYtSJQ8wvOqF0Nj6NGjbS
seQrcoO+myu9QOBNj76e5ZqFwRXB/U2l4vUwLEtwQymt/jhvHQS+KEODn1mmztxBKKRN/qHyD5G3
8gaadGBv/LCu4ZZWfoWXKc5Xq5MDDcnwU6JZ8HMCBGlfW5k9m0ph66G2s6WI/IIinO735fRxZ6cb
kQSg51HctP1ufTUmhIM0ZrQ5Nr+tKMKe22zc8XyH4bSiL1z1QQdOh06yLDJK8o8oHNj386dmxRvR
3/PpDI/RH4oEEoyTa++qe8Swtvsxo1MotHsl0Sk/u80WtBaTXjF59qegm5xO1SZNroew7N2pNKE+
GBhe0K2XVvq22aRbmshyUOqv8HZr+oYM+eqIO1J6BU6Sat8Tkqk9a/3a8BPmx0WRTSjLqZV6uy89
q9i12fLA/tiHb3rbCz+CTWmsp9MX4GBXCtcS1hJZE4mCXmUzZhjXSLd/ux3mupKGIgWqq8RSgFCB
VssmlD6/QGQyyIxozv+Vt6tI5LyZz3bc2xWL2h4vbcVSTkzNN53U6k5DJ1iKX0ofz4iqgcTo0Y9a
YS6Fv0+DhxAmS/6wAPvmPzlSRURcDVdGqP7ad8gsU5J8IG9Y16VKi70X2fbReDnA/UkZJPFYh+J6
+eN6CbiXrvtRDaQHaI4Yr9ANbQY9S4awjjQT0i0OuIz9eB+aESTgucTYlbn5MFmaki7s62v7T3ix
Y7vIIn16cnVq9kZb3a6DDP6QpyRKUUocv1j3fxfSRkwy06P5cgnw8RcSexTzFLZrG2S1uFRYOPrh
Zn3cWiFZ1ZqjoDII7hoDIv0lvsMYPyfvmvHLRlMJ4rHtygpotsR1CWqzXhJSU1jYXwc3KoDws2yC
a7SSL0rVhE3RR49yyjI6zQqzmtyu6WggUbaUzhI+JaDIuI7PkZznaOrfTJ4JpD5yV1h6kedXXmkU
8958OcV/3nwA6NJJBwviSm0xdmz7+VKxq0Ys16zmUo9nHRjm2zE90atM+wE36RYYS4dl9ZkD/g81
iuXVHNAixLqMyUyT/TIjQ6r7sV1IITxmYDwNJ6wacO4zxfgRofTmx5GLockkk1bt3i89a2IsrUng
LfazpMPz53oWF07sOjzENndBYdWpKkNICLoBDjHXPLkMgnVbRfqdam49yFZeveMETXiy/9jtHhJO
yPbR9jgLdUAGnmXUhnP8VUn8lmH9Z/ntteX9fbqpBtDD9Y8Sgi4OgHD5masQpbV4dBCguSp2De4S
LoFXKYp1UY9CsR32Kn/E5hBjJpPlDegpJgfrpt/IIIQvnKsx91H+cpT4CaM8zVQiBb9i/SIvf58c
LbwoeUEZn0L/wHxZn7cvnXuuUPb5wfJLLd1VffovTweCV9rydpqBpNGbV6fy84PdrZc/jWXgWzC4
HgT02ZgcQeYPjLIH/lciWSfZnGol9mLJvJvJtmnTEHjKF8cSHEnPozYBtZv5ATiAstpPApRknSl4
U+LwtNgunpjuGi7/5S8pvCMCeSoDxOO4O9giX8HDaq8UDZf19X6kdB+BEOBRUi8j0VTH5LaFGodM
bASJmvesxi6M6JbdTGp4xFpnOJFEGaIRgUyHzSgUuYhp4K9xuPeXmBviw/zpuRPIlRhyXw5dNeAU
Ht2z3uerUlG/3xmT0PDs1/EaqnLMsM6fR3RDCI88B6hE4nZ9rSmtRRx+MJ5QYQFePpyUNi39kWWN
IhmKoyOdjoIFTPa4ytXEt1TcReuQVcmKSJNNeIajB36lXt4lp1ZyvrehY0TcHwte/ZOa4lxpflSw
yEEGYNKpRi0OZl36uuvxwGA4kWZeL9N15dBa7c6l4touwmISUZF73tJ5wYwik4vCdmBSiMFX0C+D
VGZ8/js26s0W78M/DKs6nswt3VFds866htzyQQsvrCgRVJU3DvRz00NmlOyeM/Eqe+CnOZyEblc+
8hcGtw0ot6aEU3RxeczSCbxzV+hRSRpshq9o028JG/KRh+35F0Lpmkwt+YVXSyj4707Tr2R+oq/Q
UmsmEyGWCVoWF31oUYHqwF3fF1Uypk5EFO1dknBnEhZTDcZH4Jxhe7ubxsObtZHY8Wt0Tjx1ynSd
Fpx8OSRkyxcXaITD2iQlPIiDTaj5D2NICp7srtxYvSx/y2gPIQ07P+yxKXTNi30+aEdrKOqIHPtT
Wuggg4TxGlkB7bOEQHY4BeWHpLYgvf55KNOtH6vDap/qqUvznUjX9tQw1S3vCzMlxzbDc/SAanUA
Viw486Hk6s/yKkjhqqdMhsL4CHGhoJD8VV3R9fdT9utBngpAfgdSkEaWuStHNAETg6xmrRM7A2/v
SN+EF6f4utksYcHa+UycLETdOy0+UYmF5UGN7fixGeHyhHek/AvhHJ4bO9QPkgQAUoj4nBcwbl4i
OQzS5AP1MkGp/yVXp/TQc37IxvGWb2B3RTOvWtYXIoTq30YmbJyS2QxjvqYRReYPgPRAvWzKjTY2
gLLrhwkXq9jwG+Rr9wR1ZEmaZw6GZM39zHmWPsKuQUcYuG8WYeKHrlpveUi0H4t09QTTxiqESUD9
yup8ibUHQv5NV/Y5CuOjSOQR//c11avkpuTz2bP0Y1foTqvvsfRjNA8GE51Zd//RwcJVShd71TvL
fH0j7Xci9Hldr5q9wJGqScisOy2yTV4toU1HM4ifgSU9a6JtmS1dN65Cw/XhEerMdNW52ZroC6f4
3PazyzziBJHnxj+vmJneKXEJ9tEVjoazezbyd+LWg9CvB7EkU+pTiU63Ym/fTRcpZkOmKReP3qD8
l2rwKONC71DhOYjBDF+AB4eRu1dHbcIym12Kd6clsokhmQiKxKabhJSO3bYjBBT2zJK5JUTgkDIT
I0KxgpVCxCo20ZbSXOGEQIoFgHm4ueFJLudc1/St2+0J9GWss91J2duQ5/P2gSOAEbGo6Xq7czQq
KpHcZqI51vU1ToE6FWh3p7ClscuvCfRI6Wrsd7BexIF8oCQ/FHJ/ivDbo56VRIYhcNG5K7l7jsRs
G5S3UbWLY/zxe0/ljzgUOHHJl2utQcyM27NHWH8dwRuSarSVpSiE1Ey1SnBvpLosASXg3vcyq8ZY
k0xBv8C7jcJwslVe39bZkvIQAtsRUgED+3tVC+ScUgWq3Ub3I7n7qOqgdNgX/dNBh7fctS7hX8A4
1J8ukibyABuDu0bhmtfV5QdNd8zjPI4exF906mgXNpqACCEIsHyXYdtTHDyTuywlDCI7BFNfbR5M
YMG3m+xzMVKbUKidgJapSeU8YNkVYe6GjjENWktMQmn7Vr14M4/gxgE2UpktRTEIzsYw5QdU187w
+zhCiS2L99b2lgJnH5nfe4mAXWjpSr60+brgDGq2zYCuccbNMMcen9ra9yf5vUPbdX1UtkRYBSOs
RJJ1p2kG0na8vE7prRH7VD6g1FNebisznCKkTU1ORiePCk8M9WI8Rb8xtM9p4000VgDgk3rO3gFX
J87f5VyRPpk74OWRo+UnQ1NrzsjTemB5Ggwb/ueu0jW8DljKLvS7cEwEN+KmU7R8xscfDkMU60WN
EiDEEjhGy8BZu1rXkhGya2s6kPvsIWjA3fnJGupbhWKT1KZwU/q77OT6TeBP64BO/gVkBmWtoJuq
3JuuSpiEKflhNS3uKuwqmr4UeRavhilaFDqIldpX5hlws65P8Uc4WR+W8fq3MCCIPGo/cXQew0CJ
PJKLStbiXhRAsbzIlJCRQc0s7OZqQITsni/HwFI+f/JEhTXIyZvABCj5eMX9WI3w2o7nNxENbcCb
p55kL/Cq1cd9HT9vKNx1tz7BJ57/9rU/TSy6a7fkW+0NU7/63OtO+KUtqQN4Z9bddtC7Z6pgd+0F
WA01Rz/S76wum47thXbB/3404IlGjVHbrLdAEIu5mb7rq2LTvt3ol9M3ryCVXjSo458M+UVJsIvY
015CWLjgFdsMTEY1dync0kVh29ryBJrP8fSyM2vZmWuI7GK1+dbkheRIgUlaByN7A8+gFMpeA7dN
N5eRbz7ntoF/kgGkZJY+1XfD+A8dVI3xqNeiugqiJ4Xw3cRf35AX+sWTnkbI1etxx1cs6ydhlBpC
4O3hZMVcApVrfKZpfySbXsSQ2V2JQMl/n6y/7RP+ENZtT3GlNRIBUCoYR3u84RPqQGx++WCLAA1Y
ZuMzGu5RTR7Se+LwevG4oL6CiILaY5eH5Tsc0RKcYnH5YzHXJ6aXHYs7RgIwgX46/LaoW0eylep3
OnuwvAW7JFIK60WvRl0rkf4tYo5nnHiLiDyke5sAiHsTsGvELNkk9zwzx/E0rdxJJm7yJtSzUj5Y
RBHMFosc/YGSyTYzupKvVTbCqGnlf7cghVG45SE6btNV2LwZ2SuQbfRD44gIaUyQTTEvyK1W2tvF
fypKsKEYkxJmOT75XScqACq+FwWxyvG4eB3kJWWmJIF4lvhAHBZ05QphgqFcP/Q2d0un2wwuOlzW
4s5LMABB6lgO08ryCN58JsM5ikfXa+ON3Hnx6uGMGVHBkExIdwNCQyg/oaoPbbGgKfxm6fb+nfhM
6oTcT06ydWYED2ENL9mTcZbNcBbCqT9hfNBrPdmEx/kUnQV/9VtkummJr3stgQRPnRVEkOvLg3D/
Sb+xxhhFJ4MLIPnRsqjjnDBevS7ATagupRubVYvvoNOsdur5qOa//ilD5K1RKfbchozOrRgohkkE
qYK0JFyG8aCt7rZzKF3zrUq1HgghXXitZyYEV7QWUBrXnbWB/kM8UCYvvIWqF/YKTJGfyySmUr5H
+WS7glKi+wX1UUHa0hS6wY0l/Les9t+tG17K/JRZ0+vvNgzUrHNM0aCcxTD59eZX5O66qaauVlUW
4WABja2tBjffv2p9XoDQc4T/t7OQvGNn/LSsWOVi7mhNgjydCnW5NulZEV/FseBqKsK7BTZKo6nQ
yrapGU01SQbBBCCKqzA1I+/L0IGtm/nzxor0hAK03TiFNfX4fP5OS72hTzpeIRwHlXWS5wIlenAx
jdnQH9+SJRwqXuuMqCs5HKpXx0UzC+XbAYtC7Klj6FJbAFlrSyjcHj1LnLfo/260aUScW21ElmZ7
SLOUdDxIS+fwe27+NLNSgEdMHPUN3r1BR0nC2l/kgIg/cUqeBX7DTwJBCUh7IpqCABbU7PzL7OBy
2olTy/Whd+Crhoud8WYZQWED0Vua42TsB5ieZ3j9QNlOz7YDk9HJ7Bz+Ifq9O+z/3oGdopa/CMOn
b/P0JDDcQ4rzKRzmUpQVvSoGxXXK+zKtyhGUqIWVJA/JhJuwEdbRm3lt9qXm96qBbBw2nCZVqV8l
qOwLwB6aIX/T2TDv4qDEDU7XEJAV9K4fl/RGJkSwLVuR0Uq1bJ0Z4P7kv/FeB+UfIdycNUL9Srzo
8NPBjS02KF3KhY35XuVzEodFIwT0L8gq2m3JFCZD2z9bRXpS5ZdwwbLI0bV2jzQjksUanAKABsSI
/2/fpp9xcH5M9I/p0ADHTGiFOUV9Fc5jyhFA6W7KC6WUKYPMyssROH4Bu6FeiK+SCzlGgejXi2KV
IGeVdebK57k9U57+cRLmKPuKL6RXDjoJCpAjlRXfez9tq8oFbltYuNlPe4qcrPjEMu48wXu4PEto
W+C+RIxc3RhQHt7SEic1gT1VRasAayNGd7rwnZKtxQqtDiX7gR8WjaZSBwfObbU7mHBNRBGMOSzc
KJxMyLZ/Xn16P67xAiwKEI6YnELlDIHuf4kLRCl8u7l5lntup1x6IfI5TVcN4LhxaU9cZQL0jiAp
glrDUI8p3tINWpLsA57aaObYzS0MF+EywjM3jIkBE/3f5X5g7UQW5GMIFN0YIQGsX+6UCyRmhNkE
gChhurU6ruqPQ2yiK3KC6Wjz8wgXu3GJeiWKBw0SBLPfN96dFwpmDjaQoW9Ajotl+O988Edbl0bP
Cdo4zG3kcyGsSPW9BpNezEO9Tjy2wBJEUQsEvG7/huLQuUwcahW3bo52UWnn86+Rh/Mn+MsnwZoc
uUbyf6n+Y4yyFxmCAblSPeBmtVuqn/wDT4Fy5VAz4QJlfQ/ACSTXL5LaGimxGRsYcJ6uQUatLcVf
dj6bcoTi6gfx/e3wy+/hNoTd8FFR8f+Jn7ov3GSWluLl8uppoIYKN4u0guV4z+aeNOtegGZCczt+
ESdSmLSrcgQsa25+phVeckzHHRsn3GjJukXuQSAOPFJk8D2reMQgskW8MWhiEE9kkoK3YVQikRUq
QXnYUPE3W6jnxGIc6ZXsWP8ixNXfBGibOfFs5Bo+g3yu14mefbd5kCYeXAfDZ6jFXvBlQMkhPrG5
C6L8KVvxZMP33gQAgb3+ybvcfReXQPNLWwFMc+RKxX9o4MfE9LFEAvT8GVQRkry9XVyhapiPEoT1
tBgyTnq7c1uarjrIzFrQ9Y0TPdI4gNUyZZ6v6TAM57XKfwgYayQL+DcGTGVucZZ99X34HPEDvP8n
FJyyjtOmc9KoytwF1Gx0xsCq8quBu9OshD9vrLYkp1xbNT5R0KFWMaKygtWL4b+/qqbg9hui7/FZ
yvE2igz4o1WJeCeIN1pDbUYVGP1Ff+u7vN73ZQHWbkOn9fjkuszxmqK9Nw/8fMV4UxKvdhFtBFRq
C/FTBqRiZnY/kckTN3ipjfaf4ny7IryUOPxEZNkIkThq3Dp+y3x5QLF/jrxFSumDTDEpenYxjIpY
7YaYxxjkQkFaAEoDLuTc7DT/tlSVuaIXDGcliunVroopg2q4CGHL4BFm020RBUKdQjqSF4jQ5FOx
x9K1/KFwMdzGeRBwThLUzQSYLblX7Z/G/vioFgcXBpUDkihEM1391yXsXQTV1JBk+gkeg35PBtRK
Z85nb2p42KMMkBq4Iel8eiYYlO6GR2KO5G3ORIsshHjQjw1kwuAjob+XPT6Drzihr1wQIlJsgwpR
GMsyRDiBHkY6DAWyfOXFLbTg2+Vo0b4a4GF972SGp9ZV5kKO6BlnL3MkMFp2eFZGKAgCUddNAXcx
3aVOWwY68hKfRq2BzO2ehILAY2KMcyUOU1ZIoQG9WdzLOyjkOcGzDE9oEHOhVe7suFKH4m3KD5wt
LE/7uOnNJkdJXmF6hgHg/XQjsk216kGVCc87pn2wIjYUCFn7npisRZYXHaElHHT7SBOmWpoU4kdw
ny2mK5L82JgjtmYUv856UPIFc3E3YklfLAbcxxxsYzfg0ewTbnT4yiuLUe2Xla2WDhcmv+wci+Nk
zaC9RAulyOCt7ZCu1Fm9HDKtW9M1z3lSNpeiaPJM604aH2/D5QBLe8xNZQF0RX0XH9r/e/eJjRro
7AJ3QiwClwnBuk2rF2yhM53qKXdZpOv2TfMSO1S6EfwrSiDknWQJJ4VsBxXzH2sjx27GT1w+uEG1
oJ4KUf/PryLhTe6qIWU68QenyZAaQ+6PItP+innsyJP334e/0npakxgx5CXfPtbAJO632mSDi1uf
QOWFADwc58bDzGXxjIRr9qH+u4addRRmqjtuk/QQkDB7Kb2Q7CBQDG36ZPUssswMHFVSGJU9GNCl
wYetSi0p7VYec/Ts/TNItP9rT7E6cyQ3Ojzfm8IMlmRdEXbUxAYNC/gBLQLghVo8Oki9nKtxJbfD
o8Bn3D0K9v41Rc/C75/iJK2dmUJZV6wquyrXN9GRn7zRiA58+Cg8vdeJD82o0N4OCKYamp8Ja+/P
920OMaDRgObazf5AzvdY0HCVJMhDVpphZz8ZoD3Z/CATVUbcCIxpsbCBy65naQLlBkMqQAcuw8n5
Iw3wBeN0+FoXqWv+lAUdzoA7YeA527EW/tYnDkVexOhnTR8NXm1JxAnoLyKQsuxNPotEe7nmumaE
pI1jG2/jpB1fikyX08D6CFDVH5/TKi9Os4ED4yWgttEMR22VjN/dXOqHM8iIU4+sZbN3/NtKE3OF
2PUFvF3IJp8QD1C5lOcP390ljcAiSWXCeRAv5mEwBWdhykUymsrSbyigei91cxhpls32HKpTQA42
sjDpQYoHG+WtwX93Nym2VO5JzAT/0B0COQLxVZxvb3etuGODFLHYxzPGc/0Em0P5l4TMFQz6ph18
wMTxbElAAOmG14uLgf75pKewNJq77NyBsaEBZb1reMmMOs0QYDVJij0fm/eNdh8kDTvEOiS3e1O+
6aYH4+R5O6wyaR2+ROEcvqD/FUFYQBDIZ0Nz75uRT/Rmtq3hQUzCv13wiqn7ZDSWx7lnLiSTNUcH
J/ZrKhQhVi1/zFNXQZNnT0mTRNnHSZJc2JzCKphN6ut4MlpmIR8NyMpRhXaJTTPxm+rWzkdATXWM
wgQrhIFBDGg3mXWyJeKqLZSij5Q59R+IWwoAL+9tmrA53RL54Pz5MNBBb1cmRjlpqFm4dRSaRPZg
9jIu12kR8HCigUTUBTH+guPVOHa98I06yFDgzVhvDO+HqfApos95loLquMpibDjnvNywJMB2g30h
WGFewC38JNWqrdJLZXOQun8kqXBaaswqKs84ph/ut0xX2lW9seRLMxk2PXFbtqQsgR9jKCeqDLRT
3X1Pbjzn5MGouMqnFLtLagC3a+SRipJSLDKKKtTtrmHfS7GCUJSiYPyoYu5G3KsCdv1KTeFf7yUx
zHOCqclB2v8w2SZlN8vpB0UuJrovFbWwFH4/wOPkyKA0x6QEMthE1wIKMGECh5vJllKHH9aRxjj6
QAEmMNcjgDoXktxwTG3G7Aiq7Lr3PJNjL0upfXnAQp7wS1Q0ZydxdoE/43S7DnL1qVoBKpxix5ay
CAGWTw1HlSDosIeoyBu2cB3rrXJ59/EdlmleghhNS7NkIy0wmaBIErxO99ABV2hnXi/aQvkY0xD6
CjKt0hYwN/yQtEQ/mh+CYp5ewRbEunOdZGSl2MvBtBz3KxIW6eNC/HT2kX92pHyGG9pPrRK60cfJ
Utap5Ye0ZGCQnJK/HIK9qv3NWac6D7nXKESGK1r8dVVlS89SfZ3TeTxvPN+djxHw8S/cPnxn5P/B
iA7kgrPKU29Xn0kV5n/Ch2C3dRrH1QHhc5JDnlerb0MWunlBl6wWPcvqxY9ru0FXpuIpPH8NJ0ht
SnPvFBSwbNcUvFs00vL5kVq+muoi3gwr/xLgM5Vb3ZLVcJJ862zuliP0Cxbh5oLq33806Afx30w7
81yZl8QDdPt+oWenM6Eo1Gu48v/LDHlgL6W0w3/E0QCqGd+Z7L16FsYneuQYcFvp1pc6Nip8JO+W
K/UBItf3OgI7vKUYWEzRGpWksBvej8hOLPSvaTylcSN7QLPxRnuRPQxyv9hJgOtPSjd/pG5Miarf
x7FON6To2UGXVJxWqjuxM5PxPlsdWyctk1Mot36lS47Ym++mVvj2UILPvEE8ZCfO7vE8ui+rO0aa
254BC7MwOyz5YIr5EeTKazkVdDZGYOovtePx1KSxI1weVcJ7mZL/o4WFM4J0NjXjm2iBsBVCTU5J
YFWuO3HQEex92yI3UG1wy8r1hqqGdAGmLkCx+dAsbUAC+6LF7DFn3dK3xmcsiu1vYLHcQbgNkYcK
4ltUhc7r5OoPpT+hQT+ZtJQUn3XckdaeJHOy9mip+gW/okN2HmM4SGBcSddIVoTaVrv+BLPxFuqN
k1iaIs5Y8UI/DisGXQXe3yAAuhb3vU8dwmoFetEPmsfhuKu0fO6QyOqRwwc9Fm8qGlS4zyIpuwTK
dErrZbl1mEio5uoWSBmL+JGAXmWiCigYiv9voohF/J0RQlx78mPNmRcjKKTCXm6VkqCASexKI2t1
LEYAU4IQEeQrdESf/SzKRH4Mtc12j/Wrjf2BRFScFRyqSyjgLEIZCeEAfwnsAC357RRAvWUuqyfa
hQJ5jsjmFMNpRcKmVkmWInQKp/YLLp6L1zCqbSDSkhbHdwTo6Mk4Tn/NtJGs9wTFAtcpXhc9nfwB
zpCXDYjbD0bxd2wmCZIo4qcP/6ajnx5xmZ2OCqhDHn4kgh9Cs+oBNtoAEvCX18pEYe9IIyKxM/S9
x+epeVPuzykl4Jn7mXbLmQLsgsbn5iMC0Qcaizlomhz7OQzbSRZq+JcPPCvSzehuAYUUlmtv9Rvp
vnDy7QtTPwEdOBmV//UhfyA/iWwFce4e9a1knpc//r1+yDtPh88a+g9TvyNJanfgvDF3Ew/xSpdK
MdttnsWCZLZ3FdDIRXNfahjDlCqihBuDEnEZJJvkECiWzZKdpv+vvueVSr3iaaMOGJxMhqNUojXM
2UuId3rmOVmONRVSovZGOmcppEB+0v2sIcN4TrY6IFyB3JtvPusKVrUM14s7y2cMRYPEQysMIsKa
GKfjsv9a9V59qzYFI+3DFevkULjzYaGbCqeZ87E+mTdikTUti/pna/fdVmWMktRhEJB0mLtD9ToU
LZxJjFd1OzQuUla6huGW01v8fbIvFcpB1+XGdOmeqQmMZwGaC1fcmPEUFN2FFnsmPSztGjg/6oAY
uEdNzzgjvp4475kE1gWtA4zG73fw6SugWFrvtD/HLjb5ZCsbAye1j1t+v1g3b5lLgrmkpFuHi+c9
RmwBKTJnR8MVfcpguVsiPRcNaduFxcHvFFtr7f+B2YhFqutmVxN/YzpK2aiJtD+uzKDzj1+1CRIf
to8s5HApYPEwMVlPQIrrRX1IKoTSiDoPH70CSsZf+T3fHHGklpqkS/YyhVuK1CHK8BaHjYvrOTx2
potVkK1N08Sx3lZC5yBXrIXhWlAihjRDYyutfsDgNnVpL/PLpRKCg+KFx0gaQTXJrCH//fofqUjf
Ek4xIMVtW3qprZtfVtOJybZ9NdtxywAc6DPr+mp2P7PLBZPLEXWlIZ++sdakQsT/vZd8IBs4/fya
WRK0MMZ9Xl57LRo3K46i0i9r+C1HcI8oV0zsk4O0L+2HB6Hrwim5L9b0EThL0ga1vcMECCdaCPzr
KFJKNWG4Vea1WrZmhMXG/OwIE1clpx8UC7tft92/od3jMAJMZGj4RWDxssx2Rx+NIaQewuTtPxIO
pV5A6xffdR2Xm6GeTFIbXTU2KaXDGlIZVw2sAbR4SE5m8ogSNZNLuCdlyLjviuL4wj/5iDc2Xtxi
OLGOCpHmU3JieQ6cXCtK8MLZTSog9ZJgdAUzcnnZTXNna4znwXKWDTsdLm+EHMWVIxpi6Vx+qsmy
KkY9fY1K3rO/HXnUUBTbcGUeaj+SMRfb4ONdRJydTPRO1wHXB8Mxwz+aDhUSKI+GrnSpowSzvcbd
DTnuHwRWWMr220j1utlGwdvoLeGKQIZzyuafUAKw3jJHDyZrXT5gABFtSsMDbc0PEPEOe1QGAFG3
XMbwkjudmlcsGJ3o/QxjSFigC/WrqXiO4wtLQ0OSJ0ecj/5BUUuhgBaCjN1pvx+4Fw8d2OH9OYA3
4DnXpus/bOPQzSrxOIrvZBV/YIyWb6kpnWKaaCdYGqc/8DvAkjO12j8qVDRezow3S+bgIku8yF/B
1zw0YaFzhi0auGbmPydAKNK/4kar7RSLodmMBTBvwi8MoCSLlCaEzc58n5Oz2mYNJju+UmFtRkZW
uNYGhs5PxBhfzCnNMqqJL0lJ5JmmVsAjNgNr5e3ARthHHjdAEDYFIcojg68oh7L1htB3nIF5B5vZ
KLuKv6YcaYgQ0JPN8hUoXvMJp8to+ZpQbBBwTv0MI4XjBW6Y2ZX1cMdPiALb4AsX4qQStAzJSJ5x
WRBEshU389HqLXFMQOWYFbrlk8u1EObgLBzfcikCLfFF6xb7jC/Mthlwty6PsHUfWWiArIsmntSo
Upe9Ck8UeaeeFpCcP9M1safm5D0F8fTFqrPcEKHfElWv714giIJ6AM8QwZe+yBvnd5okCuMHa/Nk
kNi6EdPMzKsUftDcPKbRWAIaaRB6CaLkB5SQycvrjN1iP2Xo7z0FPCnx1GiCA3WgGYq6FsaCIPuP
fqGkuxNiQIswOFYKemakIvM8kNE+hMloEybQNQqWSU1jjSKDWc5Cv5grSlqhHLupOyLwsJiGxpYK
gHHR2c2vQIA7cyjP8WiC+0o//d2shKz2d2qK/hgQFzboGV6QULpiiG4dKmQZIeN7TTKluyh0xryz
KmV7kRdHYnVUJxnsDaZDLTBh19WWh9aU3WhvBlOUZ40+IQ4THa9gu4zivGuaPrUMnW8GkTue8p5i
KdcFTuVRo7cmJIrAJXoUNmW+PekiX89MbFUNKtgPN8aGXF3ffh2LnLd4sAjApE4DVCDI/2Mpz9x5
hNh/hSR6dlTllnvVBHbfnvxRINDWWcEg/v5eLFQpPSPjq6XO5IKRGra2wxtVLidSwm7ploVWhf6H
CDdvHOKkEWbBkpNVK7n93YBGPcwmuozgWqcsEVEAe1wJCOWIQ9e/Yf8NwYZB1GXuQAw1VzOEH6pq
C5ptKe0MMEyk4gPqe/WJWbv/dTrlzIOkHy/2+kni3y2zn9tUsojFsEKMt1n9xBXvjCIRYxfwKhcW
NoewElRX21sIbe7D8FY3uSVcjyw3UXdaHThnDy5wL7wM8Xfl/2BmFxAv1ECY+aUA0kXkiUkdYabS
25IElF/0SFkxaTjws07Hm/y2qSuC59QZ7OAxhJ1zfxBVKKyR3VhKibKkwVX/6pjn2eCTotVFBjOi
TqVdjbeOuipWHHugkdXe1bvr6LzhasnEoHhCZrH+LRR+L/Cxfogz4ZwgSptq4qCUrqEeShLsJWhd
PZ6o+uO/hq56W1YO94MTIpoAurYcHiLiwfRGCAqIkp3JBHpXOcorwLt1rS5kIUo0uJMcsP77t5Ep
ZH1dcfP1V6RG+eob2FCVJ95/6C2lOWwH153OVR88nrxkV7NBqib/aE9piqiXNX3HsMJ0AQqz/Hh6
65a7KdQslQsgIBxKK1gp7YB11PvEHRy953N6/JBlgQ7ZK8B3n/w5lns7sVl1Pg6cmDAyFo13lkTM
TXpGQDtk5BlP3sQw9LeM4jqJNWlqlj0EXSRa/3xLXv6F/yUByJJrITdu0gwl7KxkEKsiu8X0QOXg
eU8KWWzeowq47EW4VgSAZySbXcaOXDBf1OU6t86g0KndveRFD83p08672TcdaIit/zHhGn9yy6Km
W8FjfkRG/MppMTQskStdJA5VPeE4UL+TdR4/boUam/drjbMtfiasl3qVJkzkWRveI/MUOeskYK5A
LwtKC5ojRrAwNuN9G3+MPVboEZ/qyNNGfMDzfFDVDarg/8twKWZ5tQ7anKAawTW9bRdNdYIvYTb7
sCh4/AHAeegj0dEsCX5zEYVrgjX36F2wDHeuNFddx/uukwMeRz9xnjoOOgnaKfoHWu6Cp2zf90N9
TCRovyiLk1zBpqXicu6Swwn57Wk87SsA/sezT1xw/XOolvn5VhBz2CGqFJccHhaSO/fCoaleFtXT
e4C4eqTHD6dWCnSuqE6FHEaVHYIe53g1Z4SnT2/ac6BuNYdzDCQcSNlAMIN/fVMZIH7sA9JNjlUj
0T9n5waU6Zklk0QaXrwLEkviTT61w8ua3ageWTFQD5zUEm5ULU4zDcmbdbeDpgcLJ/zLQaDy0X8+
GAGK3c9LqYjbLIbU4k1CPlmiGA5kDhG0LwE7J+oJSfjdO8tav8YmjHlwo26VCqW9nSA2QS5gyNS2
wuwY3mxvIk6clT/m/j6V95PAF12DuyYX8n/3kJLFjLkCdiUMHfOEUGjXpo5NJDRZTxl7P+9GTDX2
5iGzpAycMLSYYFGssqstP9NqrL8aBHSiZAXBLfpuKk8Gr9liuhHaWwKSw3KqOTvOLldWa7+fOKVh
QPix0pc8vssbhIakUz+c9vqpFO2gDxpaFK/E6j5jjnvUaUlztxoaXE/QCoyqOuJ06gaTzc3JaxcU
371217ljbssEwwOdwWiVaXmECWdJutZBC26W5GHrGLL8kxkIZpTx4wy2j2R9L0Hj2X4RooXCbNmC
QzL6KL7zx/p+kQtPHN677IqbzJGd4itG37KMNKaJZsGsMK98EbF7/A9sdG2Z/UUpu+mi6VsmSorl
S17T91gPfxnYIU1BLxI2NHZClw0AYcG5oZ0Qwe23R1mbhbwNsOo0iopdGEN6ECtnSZqjvCbGMPFT
xyd8z42spxSoBcMxGYdEas3xBR3NTVBbtCGkBBjSquVms3z7q4nYAAlTQ3AAYrRh2m9eMaeVfJsF
wn0y3uEX8Hyd1kXKhWTtqnJrjigDgGNAKOmW33hX5Jvy2T19Tl68KJzHzZTZIu30xfrzuphfqWHr
rYiLk0pumeXuK/e2D2aBnqQZhNli2KeMuz7TkUX5PDhuCCYDDB9altZnJ9VMSgo5jZ17wztoc8NK
UsN+3IDiCCfwA9Z+rd3pF7NWiSFGbueImfhdM6JlyyaWo/ghFeyaP0+QXKeVQ0CcvrndeZwHioBi
/ak2636fk7lK1BO708SkRtCWRswwMPyNSfgEnrTBztfhsStPYcLTcsTc/ruMpZyvR5JLWa5h5vdo
5GsCLtRZXK5+7sKhnBfYa5fOQnEy2B/1VebF6Yz1wL6u2MqlrJViUkPShcQHfmbu+C8juV1jdOZg
DewDRMRz6zvFRo2SayrIpeic3Vu8g92msQfIIJG4CkrARrinkSaSTVidBMchO4oCYRRo42jVG+1A
6tSMlXFPRmfvgxFzml3T7c7R3HlBoXT+vkpvIACqUTH43K/0uuT/2ESZkgxmcWiNCDJu/uIXvEAs
tFMYTytUUZrdsKoLoSnOX3affCKaciaSLlIHqBpA0/bvUdXCFH+1W+J15FmBKCvJ/TV8dc0YwZfh
EIcO6Ct1KED1tX7gKQaQb8EdBLnxBcfHm+ETuhDzENpKuaTxLYs+Zjm4VzPuTi31gP73TNL6JQYd
iv+k4xakBXsbAi6mM4vl0Vt86yEkGA7ToQQoah9u87sYjVbG8RUWY3xIYIY1xWmTuJiMgEQAxoYk
/kalFMZDxhvH0KUC0UKQvoU5VOD0L4378gnNLdcZ4e2v/pevUoVNMIS2DPMI6w4eVZJCRA6QwI6H
JeVqPxrpLhbd9B4tuYbK7/f6gzwAe6ZDSEFQuy1nEswE7g7XS2/nyy3tX4jvTuD6NGKNKlcI8qqE
X34t/vMSsH/zGX40BLZqMLi6Ay4fqRN07+Fpfbzaxk5htskGR5b42xEd/wwaOMMWxD9mdH5MIw/E
DKC+dpLCbzd16opVlWuq+7lwpct/vUQz3HsC19U19Mp2PgVgPbIPnHbkBhheTuGS3eBEXsMYM+Sc
DLSsqIgwSsd1ZCW3GAAKzWPZcjvVAFWAtBNR3yxZGsNNLRwzHxaYqpYD4H4TGcsXSORWxcsXYJQ5
SDloqnAWxTZIay9a/6OoKgvnammHeICsZBQ8qBG4oDoGEsuRMZ6vTT4vEXFuvT4hY+8T+2DsTf7V
c0JkqLLJf74p1l5ivPeTHn+pL8bA+lWYLAmkgzB8bjcNGkjHHSIaAzHcArKxH6+rq3NiKG5cdoVq
Cf3bbcu81s7Sejpunbc7ciF0tqO5oLKkiOYLMh+n4c6x1RsEjqTYdB25q+iKrpmqSENVIymxiqSD
rtPN1VQ4AK4KHOCG4ZBFbSLH7LR/N7/VFd6Qc1zw7Uo/SB97l2YYdt9yNCanpxf3GBdL7/zmzZuH
ZwYJahWyhjPVW/D6GMrTuGkh/zaGi5BCAI92FoWKHyoD8OOyIMt/ImeMDFHprvAy1B5jPHPT4fc1
NMhAycgW8TePIWdX3eezJTyYl7hPvVByKx377M9UeJzudaBuD1MBM3J1tBYspBZCIatHoFUsWjkO
wob2V3jwsxMofjKBGbRAkyr4+kA+v+ryn26AEWexynHiqfFJphmnhp3iiD+2dSuGH5kzGu2ZqWhb
Cm23MbTTpsN92T4oN+XD3txCTQQJWpyl8GkKFSsynZZnp7MKVGDJwNGnrBA5WTHOjaEi+4LaouRy
syHb6j2eoaN1/TwL7kULsSW0AEwAyCql5Of3lpBzrqGEns2y/twFfWAkVAftwR6GWx0yC4RsoyCr
duHWJBZruasQv0MVQfXfGf7ZKfVVKGPMhtZWfaCYOWd3hj9uCKkk0btLT6biyYksu4foCWf6WX4z
DXa6q7yw8Atm7H133amBYHAYkn6fAqYYi766rKHH/Ijri1jbCmI+RujQboL2W/3Qg/5evxC2/bHk
UU86LBUyCIUZM0N/7Cvft1CpWijnkcDpKHHm8sZqGb/HWALAcparNRlEI8M6X/8kAaiwyXTCbCKX
+hoQAYiWKFQuiOnt4e94by9boXu5IM/LrufFWefYUSzX3QaUMhCK+L2oPT1LpyrySCzlXpjHJsAb
WpPJwPE6oi93gWT9G/DyHgM/6BoQ2o0auCBdA9UbAOZfC+kehOtqpaveRElkKEkod2GZDXo3lYcA
uyQ8l6E/yN4xZrCoyLyp9tcLsRTpC+wNvnt+y8zBmvlMYUra3JSKSuvCXVNP1WEnA8DaT7A9U8EP
lxhHNpgdXkHACvZqeQA3v8PNPZhZ8OtOJP2hY47Hiw4UbsA3mdS8Db3afGoOQAgklOn2QsCtKnhL
29P5+hJFyzyOWviIQg/AAm8R7PxpHWUQdoR1bMWdRMpxyMsOQw1VZ28rSfo0/jQaTEAKjuRSN8Df
3oa8mgo9rB4/6H0SAnqP8FGY/50LkouvC83eBMWZxrIM62rC6AxoysbEjk0yYw/ENSNgfcs37X1U
E+dtfGVYw7JZM1998ikdWcaewaXIq/PUT91xqIDyJ5B3Qpl4K4RWafGGaeid+M88cI1G/mTyAXb7
d5zJgL/oVj9KR8xNPxCQ5DVnH+Ob0KrxWgS9lxPKYopHV8rvpDCv4JIxUHi2cxDC0DY6D0iYFDcX
o1jhiyNJIF2AG0nlDPUX482f+RzZ9+NkXGeVWRcxFyAkdNNB4DrtLzriq5ZfBdKMZ656RfPVhU2g
u6I1zfnz47upVqu+KSFXjxkWEtB0PG92g2PZdiciEd7FNF3DAXYN8JHmtU9ZJT4dY5KN0/4e59RH
Hq/Jk3Bo5scpFp4XRAJ5ElM+0lGgE3WJ+vX/L9vis92ZjkK4yQG0tvU7r+9Rq/pa5GhjRrAXdhi4
yLUOLTv2Vvh6H3CSPIFKctxOdpAk8jkfbXbgDlnJx9rZCz7tPLeg1d9j5xajYgnHeGL2yd3NAgOs
5os59DnvqGUsEHkuepdV4PnCtRZej5oCn8W4KUb5EQXdON71QwBKdrbfQP53LB2CYWNszLt9odXz
HFaPuqXCzOF52r0bp4yCMYt2kw8NQEF6RiVTAtI8Vu42coFscoP/0sQglHaCykuRP+AG+1zRmhn6
5t9aAhWs9u6A7gEhr+LaAkyLOMYXg+IFCGZ9Wnjiyt+p0C4bpMwB1vekEgSIZUEHiJ/Or1dLPBC2
abMxnOZHAFGNf12CmzdJr7rBLoLMH3DH7o59l80/ZFNkNWU07PwR6xWXctRjDEdYVwsxp0wT4fYs
5KVdEQDJtEEDrIPsK3DApBsCaOOPreIVb/ebwA3M84Xext9JLWrb9A7SbGxa3mqlr/Saa3yfomTb
1RQyhYU/qZb4G2wBrUud/jAKg5c7UaD+uspS2oLnDCXX+brPuqaxGXRpbNGYpuGYOQdNFXaCWg0G
hOOjZeP/3ym7sCdu/NEKCJbbHJXhIsRQT8y3WH/Ipq3XEU0lnXWW63sF0X6EBaj/uXEw1xp83m9k
HESb0KQYZonyIfwQ16Rg3cE1mpEJMV1Indfo+8sBdd5I4GFkVW58du+cvJLNTiHzRmJ7p7ctlyNr
GePxjWTWfU25SkCngIIkZcmL1ZyBTkkqiB4CesMXJfGnm1tokktMQoQZUFn6DffAkS5u6VHUUhQO
AX/20UFWOiw2HOWpKmNc+zXMxFLPf9UsF3Lz4ELm/q/xfvKFW/E683GsOofZOyjZBxYvZ5elDx3k
RF7H0e3kdOaY0TlDcJf+78Hu2hZYWN8f4E33VSlLWiKR/bprpXFj6vWseqQLH3bwzaQlyx1mygJo
gavuO1mlwi/Hd1QQUtOq6qw7tsBIzNcjxJe63lDEev/snprwbAJAwSYJyrZ9wD4AiO3hVGLVRt/a
ihhg96D39VRF4BoXQVRuLrpR59VVZTQWsUamxYxqlgt0B9BdQGGT5zVJiYdySrjn8zzoQ03Ckhoy
KuZrPXR4V7Z1bDOPf+Ni9WXoLw/Uqe+oCOW8GApyv0LNotwU9Uih/pIbankHAPTSwk8dN1kcy2eC
Nv3CuZe/aVsU/AaEd9a3w9UqDbNMbhhk8WNdg0Xw37qSYIbmfs7VkvuHRJLEIrqtlACLBjgYnrA/
T2i6DRRSwhsAtiFQxctWec51hRIQlm17Bq1StD8ZHqaezQFar6T8XLbPqzMAybc5JIk7r4/ISW0N
kz5DBIKDlx0uLDMsy9xUcadqcWt+LQcNH6tAzUbvXVqqtfNlXcJGfaPxJ8n9VHV2qCOxYVW7HdT2
JAuoq9Z/F4hLHFch4laBR2ckOKs03Up6suL+gjMrrxP6Z0rdLJYmomRbAWCTEeGTuSvltsoK0F8g
1TrfpbfvenkaanWiz4EPsfvkNAbykLCdvlwaAoK7PEmfIMpbbVQYcbUtpc62M8BQnvpD9tHoZcC8
VmN2/83XG0Y9VwZkWlheJ/ax9mHycs9zfw7+5foH5LZM1nAbikdRPTumtt+NjkALg14EG0z2Oge0
MlkNh6IhSBpKXglz7TWnJA5IH+qFbEkg8TzxaIfqgQeZajnms/Vo3wu/F/ZqjRJhYGwmcVm2Z0Ap
7/afUmo7+2E1FdBcnvBI63eJ+dkuUkNIaU0h56E8Gut8OBIxFDQbLfrR9g+BWMiLdQcZtVYsiD4e
j6+gpGCWugrg6i83YRa35Qoj3Ojg7r7r3AZYdnxbXluiwV3peZe97ARCxVkZmiJ5rYPGV6uwR3gv
UmJrnIZqyJs9yMzc7UCfBfTsW8NhD2vr9rzV+bWvCRbiflszeAYejoHKj1FM9egH7eysOsThHA3P
sKr5DFuwIefAkDnz3TkNNrnqtk3mX/kfWTYrZ87ONRiJZlXkRvRQyYWpbnp8MR2agzH7QPPXbyAt
H5Qn8kXVo6sFSWSPxndnwfDN3w6z7Bdre7HQCc46Ay1yGWMpVBt40PBq5qFUKQLzQw4spAs2giQz
P4+x9WHJzWkWVOyTbIrbVBiwFdyDaQA+py0CJicDsMQDF8ObT41e90KWZtnDUG97+OP0yG+YwYUQ
IzAxNLTmi4lsFuMtiukLCR+mSM9dL+OVvKtlPcw23bfH9fkbN0e8qaHLXY5IvNjafw5zoZMA/dgL
rQSXa/U3c1NNHqyRrKFae8/GdmBmdOewoYQqu2hA4xj/PBtpcDwSadQ3RQz5rtjNKv8WeFq0/hz8
rVxGIYEWMD9IXoOpaROKU5iWY8sQArTYf8zrbW8/l5ne80WYOAWeTBMeXzMaBPpU8n3eVb3xo+4N
waMCOGN8R+FuuUBQonrMhPPh/6ADrZdk+bGmUqQpLdptE8AgJxXPucFp9b5jU62DMB+6RfUvt8xl
eRxRfaHanT9rSdyyvJc6RUPSTYC4Z8WLjI7xxFsfxau2MN8mNtwTe82IcIQYZ8+q5k34I+zBXXlo
1mgIk5dgLdD1bfG0T6Hm6R0lrjQ4z92CKBxm2IUNAAF+6RVx5BsgIY7qeYEUNlswwNr5DU0O4/lN
eaEw8k9AtxDTCnjweDgni8BWs6a/U4Po7a1DOOXEeCCbn7ZPX6S5eRAa8tujLYZukhSuf/81IURO
PiaaLCnpwXYQ7wmPW2EgG3Rm5PmSG+EelW+JXPSEwvBEhvtxvO5gp7WIFNPGxGDNmU8hUZuE4peB
YCDYxfVdfJB9dxjBpGHLRTr9ZSJK7craICAIqk0qzpIfaV/qAuOe6R5AuF5790BJaDSsosacUqFG
7ahazDBj4glJmAACKsQ0YVbUaVO7DHwhGmr080tKWNwznOcXscOWy6dhQ1immk8eIFMa8IUqWlWq
JtKIdURCq9cvqB7jJHc3RPq9cs98liPWqWIzh4wO8zFcJy2xNKF0LBVKNNcqvDnZT55Xy7mAQKhk
8QmhON3hfV13Ej9uf4j43DtmaXtHxyRrsqntTnJ/0DTS4MERXaPLj/SpRgT8AietF3U1wSKffFPP
mXgj/GMd5NgpCFMF31WyCFiFfNpyMqFgQShVz+m8rvaub7vP6kGijq2X4vwiezZFzyOL/l9CgBH5
PqHeR9IedmZicrPDEn2p6QlfNYS0YjpvwXQsDojCkbL38Y46RuChsOCEh6NI6vEbX++h63St05NP
ZFoxz9P4FvTcvBoV2zxnVZxrs8/bpHY5Rd6JBTzEg8cm7pnogQwmpekb/CSlkPfU5x7VgY4GZ4M0
+TLw0LRl7IWGB6V8Uy6NMb0zhl90nQZmvjdYMON3qWtTcqu1BXsF83SqsPUD5fW5WcJZT0IETdbT
IVRvdSW4IGQVVDqbxk9BnxQRbIu4Vy2oHwqMGDz71IJ0KvfHxE7HY03C2JqnnHmhOSzASf/K8Dy6
2mI0ST5fCRv9J9LEDRr5c10iowVlZ+AjWdkmEtS3kFOAnW5WQxpElTogF4qCI1WJuovXsXAP6RSg
pRTaDH5AcwgQWPbA+og4FqSs38PUWqw4Ht3W1scLbKQLGP2uvW+LHVFYOM5/yyASDFjsNct6Jwz5
U/JqmwzfD+z39g2JDI8LslLvZSAUC1kGkmnGCqivsxNlBAs6+CqKh4cg938WXDk+0BVY4mUvRKvn
GFslF75i/A0CeDpsY56Phwkt37LApYEUSVdc0zfT4Ywk9p2yt6E60U/q5mHQnFSlphsiOvwREarP
BpJ5+QAfcyWGawojjhwiicl6MJYjuc+6RJIWjWBp7id+cChZhJYEgqfyipzf+0c8hq29DmtH1Z+Y
vVc/nQfml/41IkdNuJOY0Mr5wsM6mJj3U/Rcfot1oA9Zy/tGmWj8CJ7KZGZeiarLC73I9uJY5WXl
WSZlkDYXhetnahAv1YjJYCPdTjQjc6zJ32smzwvAwtQe2JvhCOBa067OhjltDzaLGfdx7bP7fZqH
U5feLaLT3eVWX2wkEVWQH3dzbyzqDGF0V3s/xKXfQUdlx2snxbuT+EE2IEV97tNZ1qHYv3RIBbXK
v7n3OQQEkeeK5cflzNPpgNCanVRnu6prNJ56wIpG0OD4g7yOdlBD3d/noT6NBY7kUQ9yha4ym0An
Q8vz8UUr3Q8UQpApN3WXPZ6k2xrzrI+GTlOuj4nSyKy+jTU4FanGA2o0b9S620yt+XV3uia9V+xC
sk0NfmxO3VYszB6JkohQ2Nw/oFpcxmYEIMAf5wwnMOxPcsZza3AtszPXJY4ZMH8rnHJEmVjypBLl
fSpbE2ohi9hZT6voeJFr2Di6EBhlp7Jy7yNedQUa68Yh/1TUkr2e9CcEqODkBda4VkoB0+YXKCdG
OJ4UIvMuukFBMfWvTO/hHTQMaMc2QPhxwQUKC7X6oGKXIFM9EXHcZhuzixbRoRsguZNoOq7+8pXs
XPxLnaXv9MUxwxHLJmV5dBvFXljYI4GRbU4UV9p7I9jf9zxi9+uutNT3qJlvD8v26y+rGiapG0KE
WEWE5Yp4hj5ZzAbogLIRFJ0OCyCD3K0JJTIaC+rxzFqEgL6Fr1NXEPgOxyhDyzBgnEwcI3f9E0Pp
WAYyvyP9LkW9t2IecaIGNBY5lZZh2WMl1/OOuRxvsXfis4aBQrk9fFS9RItCvq0AemwQg8qqWT7F
++qCB9H2sRUCYPb2gpVG3rWUM1Km763Zeuuh9YEiF/Eutzj3ZslfzIcFC4qOOfLnmZVx+SUeDcPd
lgRVsokXpKhTHdHpSgbiIJWoIKIkG51iddYIwRuSqrtF628jG8OK1fptAH/qPauo6kW0mHewKU4N
gwM2SlEAM9xphkQzseha/9P6012F9yROoBgicJE1tKm7hIpnuvh5OHXiClvYPLCe4h9xWWKtTUse
r6cL8Ns7XkaDNDk5sMK8EUyS/zcT7NNaU8OfGOVlh6Kj9CEs93CrmnO02nPoPXcchNo2S7VULVUf
7nkK7F50xx4FuS/8G007C+UueWaZ0pUZmHXsR+k0SGtETybvvH8aeG1R/d2UuJkEYBDJIWnbYP+X
9KTQPFvpgERR3qrvQgWFhO1xOwum4RCAgs0GPObllfvx0FM+WTGgM/5HYEtFssiBmcvPiu8IAvrv
h9nJrKNlJRQJ3mZJKI728frJyTpNmU/MmpOe2FRnFrwTBuPojB2TOKrnraSgXFeR30NWgj4Azox8
/dcT1gNTqQlR48DwPkd/LUDRDMV1QVph6VqbjJ6mrtnxLxcYOiZ+rmpZhNKuB0EtyrnMAb1m/BPv
FLjcxKhw9SnoY1RUW/SZmFEu0OY74TgQ+wzPevU7E2s62EVve19q4GlNDYM+rw98GI7jUgD025b9
yIeEwCkivrLwGsacExuXV1SYiSI0s5CztP2dCSYJVG87QqZuh8L561OpSy0tp1tmxz3gCkk/5x1C
atJgyzhUFH3v31dVzoAIrVqe6pOtVLEvDN+rT3VXmul8ju7UJjvjtanVYSvxHtb63mOQ8AIVTYYj
I7HwJs+Rs6Zy8rlEajBqOpIMp5t61tkFEWh7HOs/wUS595g3oOcUKrrP6DmdPBoVOyoF/ccwbpXU
k3TQwjEjBaZ0j/7FMMtB6zPPP9nrrQqgtW9N7h6m8/2yO0HqCWye4vDm+zWnCf+eh7CnJtEDvaqb
q+NLOYvf8NG6dzrb6DDdGRNOsareC+z8ZFKImFkFMgmoM7mUFD6pMgeA07SPoSOPu2kmDUZ+sRC8
vZBdPNL8LCY+tNOIU71HAVcIGv/80kp3rm2gyZucZThzXL7uaDiKZcVWc/yQns4M8fAsQ7rbD2AV
o2927O8KjEhiW+PrxpD51YXZ4StpeKiXZkx+a1GWBd5emvX16tSPq+YJPHny0CwoQ+19Shnqsfun
EPSH87zqxikCEhkNWNbUZxfDnLNvtTfUTcLMqLdtiK6ht0glQ8S8gY/C+jCg58pr3SsrcMyQukwX
BhzGMAglq7h+Qxw9kPucQ+xgEFcx5DepLz+7Saxk1x1SqShZFFgK9tSqRa7LefDw95c74PO0JVGC
0FGgCzhlCRaWc9pYFWnpbO10jk3+/VdI+SsWn5fzqgeNuHmdITuZURWzi70Nr5r20ix+zqbjmzip
YbTkOCUiLmzFwaz8PN+VJtJ4Cm970SBa2rp9RQ1jI7RivnFHRY+cwUACEoaRBscENQ5hbw3O9fG/
iE4l9ZikYbrUYnGQH2wlC20B6FnSU6yoF75nynL4MQa6PPg0LN/RTEi8o5ieoJlvwMtPWplt0tob
nBbo3QfxuyGptVnCCHHEydAbSuBRtaiRlJffMcVUVK5S+Exhn2fTPzNMYn0YlLrhc+QUhBP6XzI+
XJ1bj8rOmruREepjfh4IxyBxxc0e3D9+akVWA5Rg41/6yPUrXUXxF/z+2OIFEUN3DGbWqj6c3Xfy
6uv774+I9BlZbvgCBiSIJZFrdh4TRn+YnNFzpgipeWgDqrWuhDHA9ZtAYAlsZoyjUhf921ewg+rF
KpcVJiK5iDBk92dgy4q/n48epgOE6H2+1oeOYJI168WLN2rd+N8z8fYVaaolJzCZ/S1dvNfAoPHR
i/Bg7J8BaN9POZ79YMGblvq1cpUq0l9NwvbsSXq1XBPAalbUbOIBaPtMY0rWO3WUk5gbwq4hCyBC
ZbdjLUIUoTt9KQDJcKdDqkTgdTRV6lL2cX+NYcjvzjx/cbTVi1cRVAK93My5PnnSPAdVA7b0JLw3
GMjQrucdDNuHEmfP5y8N35x3GNlqPn6eMs2PAUpD+OYwHqFnLyf/oG0C3nBNpzScAi6ScoozpNQQ
EkP/5aZzOJ1Z941A4zqBVdPyL2oqm/r7zgkQlwQzWymXLO0FvXEo/BuNiukcX613HqiXS7zJmE9x
76sZGPrvoTpR8jaLKyu4UI/wANunWnV5pgV2j/ivyk9jSuVtOBPxUSOxyApdNcEgIixGDi05o2Xt
IeP3WujfCubFfajf429X6dOmXp2yzfrEis/qWlKhbnh4gSSqjEF/6E7CNefHDFojW/gul1dFr/9r
4j0/57tAtfaLf6jxf9ANk/bY5GmnDQ9BmEdR+PW4GnI3ZrATcZU0v5y9HqhLF79T+V+p8bKK25Ig
g7vWrEIQMOEZieRX6eirTGfFEPzMyjC7kH6RT1c/j7KrtXJxUUeytQ3eDuRkYFvSdewKkZrMaHKZ
YBDjWBBGuEWhHPeM7MAuxpoY1XnJYBHFvj7We11rFeLeYTiGi9DHELLzjbVS5evueQVWeOq9twml
F/dJM3HIvW6YPmyZaeMI9ynFSennzM8GdXE9/DKUJIqbOngza4NgG1Q8yCWTlfoNbb9cIPU9r82d
b54foYSJNVDzXCEqKgdjQvZElkXP3vLwg7QvEBPeF+6yf0fzo5dDA+YVAdKOZeBZpqktGA1+AAxe
gf1ejvL/iBlb2qLXQ9LKshcCBZdRhizeojZIKUuGVZTgIkfwni+uhNeUsBPaIpc2nB68+/zLaEtB
8knEvir7q/LxuGQz4VsYw8WLtmtwaP2hPmtRQaIXimb5ntX6FFm/ZSAcFJjGL5WuCPtqWoNNBw12
iV7yitTp40hqXVd1ykcpVuEG3DR8KXIaXAp4iY3q9avlaG8GED2UppEobmD9Fl5Pgv7V1GCWqh3S
1Q6e1uLZltq5G4EmTlAZxETfkrLW7z29bZ9+VAgzbCAEcU1FZnMniyWBMkg4DZV89bhMU8XJ73fD
KB2JsJNfipgzL0ds6oh7mEtnCpSk1oGN2QOyKVxTTnpTrrqEjp8wwHWxHYmW8zrPibW46KriL4u7
oRocp6YoU//D+VFxje+oM8J2oiCXiIu0+SKPsWzcqygzsrclZe0zHndVjzcZtMqj4udBNwMhru5L
BCznSj91nsqA0kV250iC2EZVQ5aRpYOHA1P79yjE+WDV5NTwP08tLtcROSUstuKDA7wCHmNCJED1
xLS+fKSGs1+4w2GEfFFZcjMxFcPtv8UESvQCf7f76OgqrimElIALd4DNwmT3bL6o5lsIfY2a3CVD
z2DoNAd2VZ0cwKKplaNnTCaXkAVAMFRlw1lU1/Vu81Mq2l4wSMxHvC5RsoO+3F1AjQT17Eh9CpMk
S7hkkPE26k0egcaUgwpyOwHOmPw1PX9MrJLDD+76QXqVYSUCsXvyd+h78GqbTmAccm3QFDndO/ry
cMKH3PMVl+Ds/8a+9IhQ0kC/dK3DzY4UywiJ1Hj6FVRAwuzmb5X69uL9m/TSDL5WouJj4QpKVmfU
MYVteLdxOm6s1BNZt4TTkoQYYOo2sIPgFGgnFJQhCPzVMBL92RWCpo69kINgeBHot7xakE0CkRdZ
LWGimPfTtwmsSbmBYgLMjZ8Lm3R9CXJKcmKENQIOlVkl35PMILNgvFvqeG3AH3Fa5bOogKXXd77F
ZSZic4My+SBDfX1xqDRmuulthk+fVJWMOSOlEzUOTKn8XNDFdEP8JACWCNaZYCF/hcR9YI/CgvKI
dxfrYGeHv5+/z4UC1DCE4NKEc8T4kVoNwuGBjyTW4gy4NKYCer+5HaC6oWCEBYKZtTILTmCkjU0M
dC+bkIYw+0NWfv8ZQrp78xgoDJuuHGrdAr4/OdH6IHT+krlfd09XLNvRvbJ/c8/uZeBnAHXX2HxI
fQcsdGoaTnzrM4BZq8CLZEymoQ3rBbheYXpJU4MR4GHYo0hD/TbQuD1VTcpD/rknX+yRh0MLek2T
R2oDHQfQa5yEm2Yl/3hTtL4GcVuDRJECc5Fs3ZBD2ZK89yf0BIA3FZPdh/DcwDXoq4utkZTu0Hlr
puWIl4GAs4QrB4Wsab1V/R0E4JPq6p6wTN2PT9FvbGrVBnOM52rLkurGYh2NFCreKCH3i4F598gF
ILUQPz/bgy5oWNezT1WLrZfz97C3qFK6WJNKY3rJhKGEFO3XVRTQX6U6QXtv82eLuZctESDRgnCv
Hk22c0LIKlWB9eAxQeYL50Eqmpl4zQuHUdilktMbuvpjYx3qQ1GY7cC4d63F4tDqcgEGPpxQmimr
lyAnibmvYCX9ZqwvVMAxKY+oCnR1tKu2XGxfaQaiMFFT3MyZU1snX+okMhF9B0hCpbyx0YhSpj7s
JFsmCE75zhXJrmh/r51inIC9bYj1BtuaIfxEvmeGWPYlWXPrULWtV3YCkEd6b7cW80Ry8hqSWsOc
6foP3Hc6QMRJcsEtQlhaa0dNFGp+Cj9N+mMe7UVVXboQ99A7fBDdA9GweDZB+JFLLxvNjUi0jws+
AzScwyH7k4El8sJ3EP3k7yTnd9PiXIxwv9S5KHN/+P5LD51QzQkTQFq5RqHj1zCf0DZVdn4Qv27N
LNj0HF2SPQuvTA7XXEi7Rqi9uMiwfLjOTTOodoHED3djHBzxPQFe2oxLwsk+xtMLCXc6SF50kl2p
KflVxN5G9bdjhXgEvaHdHUj4Dm0hQbXAzjxnlxpBoyknUfjaDIpHJ01/0EVCzsoXKY7fCgFrYomq
oxPvbufNFWm+OqsOhXKULRynSzUPeFtC3ZKvTio+F6I9+NXZWlxRZ2BWTVs72XzhdYfCbGSAzm5t
Zs2XoRNSF/FBLa0+ik9h7Vs8Rjx+a+433zr/VsGl2eMOc5icohCd8JobfrTNunzmL9ukY9KQfIZT
lqWWyDrY/5u8DpN/dpwVX0uEHV+/tXa56lXWbnz70g9ZwhIEXEXTvVjDb8wM4ZyXGuy4qQKIqANG
HqBaYU3hfs/6N9121IGlC7UXA3lPJE8ezmirVS/JD72VzPwFQY16GOq4zoseClQ4nterZ2B96Vyd
bnJEeIWyMdZljxOrDDrl3zzEcmEPhr1m6WVL4wGg48UDl/jq66raLy8Q9Yo+nzoIwsE+7cTmC4m8
/QXYgfbR7OnGC0Dwdqo1nn0jhPJkrKxj+evnByNfRX1K2g9nOh86xgz0KLtEaOjbJSiv8QL3WZ3a
oaLT1pnzRjD1xdGnG93gagj58XyHOvcD+2Gf8OoNiX+XCJ4f8Ghc0bwxS/sAWqFInU9iqJYNqHe0
B02loc5lQEXTJ0tmO3nquZexpzPNlO8YiNQgE7V2bpicpd4IvaSSUU3zonHgTm2iYCRTDiSlFvDn
u/QPme0eyQqlUORJixIhGQuohffVfeFaphkUJ+DhLYYi8isKcJ0kUMFre6FX+UNDPmOBJz4j6bYk
uAH44eFQq0Nz0futROoj8fsNJfufs1qd6X/1ubnhMd7WG1h5W3Qw57zx80Ozgx+3ukiqVxNQDopC
2gVQWiYVw1nI5Ok8o9lsBsgFWpHvWTWKC4dyRQE8FDIZshGOUy3lN+u7NI76cXlAiTiC6fsLCtkv
ZPWw8WKPPgEfGHyZ8BA1j9gnYBCfg9Bv+xMjHec8+HkimwTqub9OFAV2+E/fmh9MngVSw53Ry6O+
wiHPBif+xLahjJoq2M7OyonGgItRsRyiT1s+u7QZFR9EF9Gry92Zn0ba+Spj1MA/lc0q+08ZoJEj
3daatxNXdsqNvDoeBu1nxPcQg1fp4Is2wx7sW0M8qZ7C0MT4dZ3D6UcOSfOTZzSS80OHDCmWteCF
Oq1BmJcOstZuCQg+9B1Ht8G/FqSte3u0uOkPm8NJH03umNpv0FBywLAH76jrrQILnnKHytRRGim9
3c/h3rP9GJgo+GSFW2F9sHsPvbiGzxFqF66KFm0PN63o0YePRJWjnyffV40F2CXw7eeCWzLaRot/
/ZCBjL9FpogORzk+DHL4uw8FJwuNb6+aEX0nPIycgXzKgx1buyv7fWa/vvJM5mBEvGTMvORIveeC
HjVB4fHgklU7pq4mJsrMBXq3F7fknSIuwpTYvb+Ze+vjSCPipxH1xc8tCJcoFyftCSCIE1wKFkBw
lpCxjSrbd++N2j4NoYz7R2vixTyZPSwlxdeTpORPiTlXbyJW5Y3vX2ckZtSsxGfHPa7/JXOBDD4Q
F6uF04W8RSBZLoARQI5fE6afsbP8CQs8vt1Li3h61xi0oR5tfqGBFflC8HlvbqVVi9LnzUTA1gRM
DBWLWmN/WMyCcDs13bvkx6a+xfJb64Cj6MIbEObnF+1CTgI0f76nwQ5jYS1B+aR+vw8kC+UVCdXJ
+ofmHloQB+lR4Vabo3I//qB1Jm+ca5x182w4z1B6nc5+QD2r4lDi0uIqdBmnnBHc22/pA+fiSS0H
oK4+ANqsSiUCX45dAFtVHR8Yc1SQqj1TwvKuJncdyWc2c2SdKtmqIZ3jxcmLG9XmSbrTgLZBUbKO
XKbUGho9mPSmhQkGOZObRx8gk3ALiC0d31uP+fnV2e5zXQERUe0UWmLfs18Dhwpu7NrP1xRPCorl
OvM1Y4+Qo2GGsN5fn/FVx6IcjsfhxeuDDBPJB95WjoSCxGV9oPWUhMWvs2UiSnn/mSS4A6c35Lho
ipZZ8c0n5GHxbMpuqHtUa6sjVKUM8jpW5DMGM0VRaVziaC7tOS33rBylXJcWYnqhOTHJALZxEKF+
ERxrDgdLxHomBzllnbW6JId0wINcqYA5YrQc8BPxK2cTi7cINmjPYoy34T3r2ky3fzwfvSLKDs9l
OAhk9VGg36oEiAJW3HP8JBlPr9xO6aE9/5IDYmeNlcHSRbPVcTa7WgyshCWELM/AEXj1FEMyUTqX
seFkFGF3tVRvQzkkX3VhpjTLy0EMmO8dX1NeqIt5nwHmSI8joF+dXWbkRyxn+bCwaLASUuWz8Gyl
IzObPcKqpLhbNNWByCMNr/rRhb9UMt+unHkHFRI2RSKfkxuSATSM9e9nrg6bFFGNrCBODo5izohW
CjekxUA2Ds93BixceXD8G9JBoHr1iOrNSXVkbqPab74AMw/oVvDVxWQNFL3NC32G8TlkIcgoXg5I
iwtbRcGAdCIh7Tx5wDasEF7gjE5suKde+gio//KVp3V9oIm9UHXFhaHoe6COy+wAprX0QB99OpEr
xfx0bPJixE5ZsVsdpmYImrz7HVq/1Hgce6ksflx0Uiq7kGuC3u89QvbSysX/cErRZEeK4Irqq2J0
/w5bx6PTUzHpCvErvxEREz9PFeeewyC6KofPbFxv0FpJZpI4lYENoC5yk8y2ZlQ5rpkgaG+X3ig9
nGUZQWu0QYBpLGhEGyUSiZDk2YygB5oErsF9tFeoXwTRlZ72XvB5FEEifJ9xcUrm2hAnoo44QEt6
qnBtsbwS2CS1TSpbPEq7ah/OwaNhr9TPfiM1LK50Cw73DfNHzdfPmuPKUSJ6jpD/Kn7+U5rXT5D4
tGyeZxoAduu2908ybEBOJ+XqfyYwhyq8L1ttuZ25a744VPrjXQ9zfff1vkynu4E4UwqQHjMbOkmo
LMYG1XUkUtpcETpMxuEZoTgBLa62U45iqQ6osLTm1oCKsFcqbNzOLdxIMKBsHPwsKrl4KFrxXLww
cfhfSGfrbeFxugcUyVmhkPtbPQyk6MAx5g0zY6BAJIFra2gIH5gjG5oiSx8MoHVt6T8CpzT2noui
MjFklAJ2T2N3qhOfeslN2cGBrejUFFuJZq6xauVnfp8+Gth8xALcEw57UvitmQsJOvWKIObJ4Z+Q
pMbcJPOd4uu647AeGhfuHfMG82ke+4bxThxjjW1koM8XxoxIaL0gKgPazKNA6m4baxbqcMKZ2UxZ
5YqhESdt5KJ1MpbnSnYRCzjQNdL1ZgitIs8rLYXKbfd4PhOXTSBYF4faKRFPDQccsPfa9R8bg2Vd
1au7s8+wS9WCkqBE41nepDwUs7fX9din/b813jhtjh8qcLVZdxxRV78zYBJWHh5NsYo2UX3Ul/kP
2FU4jbo4nPpA64fa3deI9MbaKml7V1ECIiBSUoo1Sqt5P6GMJlmA5eNgQ8OGmSa7J3KpgZMVyYlg
seYvyPA8xirenBoWS/LJpMVkoIzEzVF4nz7f89uV6ewX2EoYHGy68y+IgmW/KeGR3s49uLhN6mSW
i6ElUHbu964ZWNHQyDE1PSxTEw77leviavk0px/4mc7g4DF625ShG2HDWXE2qPOWeH3WCi+cW4/8
q1O4oT/pnn6ec8tz41+coi9ZLakI1wJEbuwx2BBYXKEzg4SCJk7cyEWSeQDFviFh3QSpGmMgfPwH
pblSkMHiY6UZDGZyh13SqyXL39llWpN28TdPwkjJfW2FZpnUg8JVYMO4I6lJuWzLD94mtBvalgL4
PxMb9XqbMal0Mgz9MyqR2S5tzPlP3IN2VO5TkqsjDXI/tMHxHrp0bbYKKFXtzd1I8TCX+xBep6nZ
vF+LG0bPGo4KM9kZ6wLal3XDmdvHwYqjBzx2itG3KxYhE5cFQgQglh5WQdV13ED3y8gbd+o9hVnT
ykOZuBZvDKhyMqeJB7d3uDGLuVp46IONctfpI8tr8HT2uF+k9YozJmzp9qRNHzC8egjtb2D3VNUC
kuhKR0IFY3EqP4nbjw/QWSac5/xN8K1Wz+Dgyv3LroJOodzT14SVxexiScLsnAZNuHOZ0EUJjUgW
N5TWsXmPoiD1RDTmTxsoWsxKM4igt3MBfvcIS/BifJbAufGRNaOP5A/NLba460MVdULGPQRaNm8a
Ss/aL0tz5krDYky3jUuM0/HBMPhxqrO99jDpKrR3eiJOvt2/aKDBjwPzVOM+hBTzDHb6wLLepGsI
VY8DzInJd+i09agbJwpwI2TXwzN0hLgbBbK29cSHR0c4sjb6OwOoG4YrQGfo2hoNoz2lQAR9/1BA
J63ZixVSY+DGGJUpXTeKS/GSdt+0U1r0VYCov9eLlYSlc3rRKkQRbeUb0f4UCCyZAdV4Dsjvwm2i
xy8u9/NSusYCEqjzg3uIeYKbiAF+aZ09Tar3JxRczETybO7ViZXGhHMAEhv7BZJbnoHrxrSt/+s9
Jr4h9pCOX4MjjHrowgL+844+AEtf2Ftl2hESqjFly5uExcI8Cun+NPtF510EwF6JXePimhv4aT/j
sdaKS2vgwvHTTBW5pSev07RxsKCwNcnru93dm+17KHa6YWTUHzIgB0Mn30PvKXh2n3Ps07KcEnz8
AqoUjvsfSIbIp8TTzrJk5MAY07JlK/6Yd3m7TkIm6Tk2mpf7o/GfD1atomkc0C+VKRiTHZ7zGtJb
fVaiV+50z098P+m+/oraM9lNx/Mn1H+yBLaiyrcH581V2vtZIZVWmlKs429mjQZchxnX0dbTdsSq
RaKRMocX+vgbwjXCkZMweap1vCI6Njod7fHfNqLW62205jpFGMcz9eZrH2CC7d9lrKliSksOP1ou
tWaYgk2Ujo6YxtciLI1FD/h1CX+i58dpwUChVEC0/i1ttpg8QtPnYA2gvqS2BKWljQDm9LwXeWBT
+q/xOmMbtvetsW+lyT1SRKj74gb/wEFbx6bL6knllhi9kihXbbVxtikKRGqI6vF4u2WZv3hafLTZ
TwXqJxFj4W1GijlsZg/xZHpjBi99amQcgaxd4luCbo0TtbPO2vB7gUiLtuAC4yI6aNN57Zfya0Th
STvDXv8Xq05KGKO0mu7NzwEwdtlOM2sKj7K7RyWEqpV38n3s19oB85W1T8Vko9VYLR0b7O/upjGH
JVHfOdV/CQJ2RJkkQPQmd5F4u1Q7txy0QpzXIKi8YwiRX4W0Bm8yTVzzoEKUZSMlUzpea7jknI65
+rUm8Wo1g8zj5+M9CtBJtoEGFAl0Aksg7GgMmHzUGDtHcUv7q1cDpHwb7uslcuux9Vv++iT7ulp6
ZaShjs0RhBnlMKz8F9dFAaF9SjijbbI+hb4bMyGd5B5fLDVSkgIKoKmW8DrsI2TLvwHWegBJpxnG
6j00BYbwuZayxQBtd5xI9ZJkzI/xuozkkFJzOfQdpAyYwwidMAJbD55z8eOmjjeFB89Z5KuhaNk/
TpUXP+G9pYlQ179y+Qrq3NXf5Tlv6V1L38rYDTz5RJEAMfQCozjxK0WsISSdhTnUaGv9t+typ8zu
tXW4E3e6uBv6WNDY5B4zfOhMf33kjrPmB6xYYGTDMzGGyJmuNInvR7Ezs4XM1kmz4eRoeMCHLIJH
I2hTR84ni+hdndcplbxbE9QuPvDeVPVt8TfBjgQv5FVOI9LF7wcX+F0szhySVcemWBPoMs2LwfoS
4f719k7d+O9PqLQRzbJ5r4w+xoRMUJp78KO2sogcuDmbnbPlts5phiqENbWnEvWUUnNhIqWl67QF
njq+1lNezjatux0IBq/RuOl6MrOvXMfBnLbf7s52Yxbb7fojJmAsQpl4nT7799ccHgq4tCLD7w85
31F1f9B5q5XxAZlwActC9fMAVnhl2ybEql+w6JLBWdFxznX/xrRqUWTHpjLu082bVSrsI0TU5SYE
yIobN5lkSbMepf89Fy//Zo632aMfS67kYi4a1ZATRbAZGQTU6TYJxdGsWmAn27nlgRaDCR/dshTq
NYEsLPYrDE8IbouAUINC24guSLIq+bZmDU+N/R1mPbZcBbWxb+dMwsrYAqjTNUvcAbpj+b/ab51A
DjNF1yBf89D+o/8aXfL9L378d/DX9KMjWNDsaBffDDXauF0LQhaFKAO76oQz361QxqaKO6Gwu2u7
rLPQCjpTk0uL4tL/7pX88Tx7phVtRL1UnyOSEFPJYgY9BVIVGO9q40DWEhNVfLHRwDn8Bd5MhDyS
+sSeuR6+EwSacDGa0AG4pyPMtjGRGgbR2NE/XMOxdF/hngLyV9me5c5JoVdJSkJqiHSu6qtEoeYK
LCgD+z2497LZorIL+qhu4Uzem9sSBGCwKq57s7n9NEbzK9os+KOaTW5CQsusUfjId6J+7BpSZsv5
xx+mdwQUKadnP3YPxRJdDSVyJjCKhgLG9RRhsUIOEplDgwlzpZMMv5wIcLacTxvc2g/qPrs/wh4Z
RkA1t+OsJwDcEK35wC8/9JgyYU7dFaAGbYBBoY3insm5CYPotpujrHJbX6ABCsekxFRGCKqSqR9n
5S7pSDb9lcaciuKybRB7QVqoGbfrMunHnJpdokRSp22mQAYTg3KgIffbrg5Ho0NkOA0n7hHokByR
SUqC2afT0ZUAUTumc+N8DDCon8b2mq8zBq8TZFTvnYWlG5ADCXsjdXaOlPydmj0/gaxUIurEopTo
dICR2p0vvgpcB4EwrK4mFAlAgqU5193lGCC//3C47/J7OiUTgFerXOtYYth0I/Pk/AIzhhV3vwt/
FWNwVtXJ4w5n8S5pf3Dy6wAVAm3Rqg+w2YoveDM+OP2ty2xhyDqFaMtc6fL0UPYGJ+lulxt529Of
hWpiD49GIa8T1YJOHi7nSiZlt4jWRESP7QQuCTuMiD1iQHOxWIKBb2ule/1hTtLA3BuIES1mcXfg
iwoxi+F1AoyFQOioy+oCZMkpXUud7SrkZkgU+HFTtXdugrzSkZpMjpUDbScyeAudLJSitTAmgmhz
24zNlfQc0JgKAuYgjqyJwcgVw6WfnucZ5Y+LV1sYONSVX3s2VMi8raFlWdIUkubjXFminQ8LwOIB
lXF+VuX6aYhlj5ePUm+J4Lq/CYkhfjTvmhJkpW9yqoLIa0kD4RZiJlqZF6L7ZkvQrAgT3r9Co0OS
S0/2PNln1/qyLCKUHAbtLIWmAHfs9r+KPRsnwuybpQjem1KRsLkdPXKszmLlX84uNDyG98GD/jNQ
iqOYM7EYGp9HZ+czMMOjAuXR3d6dSBdbtfDEOQhL+LthbYvT564zemHl+cHruMkTq44xImcpdAZy
98gRYhPjkZZr3zNgMXxiML6jaMA5JPYhIPkw+leNG9rszwTVSMxlmjpMQeFPbti5zJKOQFrsDq16
JqMM6EJCIFCcHwWgCUMcJC79fUNuZrXa+v298Wj9w1Gk7M5fXYDU4Lm6Bvlu+dVUnta4Y58tGJIx
V4fSz130TxEMMN2Apt2992sESGJEaCaGEb3bQaAkX3WoV536shM/khZispFvWgCgle0V3gZ6hCzz
l3JJAPMgbyYc0VipsjTPnbYve+TO/L//K9t5B9WzUI+HCImIksOQyUIvOhJ+7DiCjI8E7zdHRiZK
wgNREUm8uQ9GdY/r8AxQSpwnEDTYyZ2+HULB++cAPyNGEtScvZJHq50ywMRe7oAb4cY6p069122B
3HMYs7mCPPlt8s6tM6yDWFu5ycRcnPZtncti7CJ5LYYRtGH6AjGmjNF2JjQ2hQ7w3lnJU10GbsU3
oDnaxBE6iVs0PFq+xW6tFuZ0diyy4IlgYya942E6tfl6WRLDWBfdVsKg1Qbim3JB32D+wc6GXhlg
eAHYOfBJ3MrhR3U67m3oQSGoj1CqRBK8xf73Tt7yC+Xq7beIAUkTOZjHygnj+Epyd5mVZzOwo/vW
J0eYPA/GY3N5qNMcQPLbjdE3WKv5fvRaiYNQutKC7XPfS+04tQ20BF7P07vuDBvUkoZFaFjQSY0Q
DfxCxhnNgUvhBvM9SFF9r7qOr0Eh4Csl9zFZJBTw19ltNGrUJwL1XlWv5pBRqEeZ7DMMi0uCVZMK
dL843V3p+aNXKLMxtMmEGObueYnWzA1f01GSvcy1Gh90jRl5FZc3JerPHNI58+/c5p9nA53Ndl/r
yqUU11s3QXXbmYK0NYVel7qYjoAc8QVooms2VWio6Rw2DgyEVZ/Vyd9Ev7ezCuUiVzoh6y0B8U+K
Lv8b7hAmm4Wr2OnJfSBFvqukfozg8QcbYvMaQhQ5ZBLZ/OrfJSlqdJAVwpAYU76Ha85OTg4KwKmv
nvOEjsJchWelEZlBRgII2hUy8m2uvklULw/6Rj9I0WCo9swlAKzWsBappdQm9FWUrFb2ii9XWY1N
42L1GUSdtPJNGUx++qqHLaRYxjXML61+peQLVeSBtI+QBulNhMP09OSJuncZlg61qU6sgrV+Sl6l
5OeV2U0Rgk7HqcNrcT07/vRjyaQ7PZguUGwQnm/a1s1YFirq79VFh3T7pMIVriHj6/HqxGX3YzEO
0E95ZHX4CkPCUyI2ht+gdmniGrthaOKqs9YjVC6PR/afOJD4+Lr79u1EoaQWzQiK2T4OJyvLLA7Y
UvTxwnS4EjrnL5Iv/iKRGRxHRZf4TnFFQ1O3Rx5QOGJeuNT//aTMBDCICOHPZgtl/KdMMqCCVTju
/oHtC9DbNo9P41FBrz7FKu5o/yelSGGSymDki6/bH2rJlWo4bvSZeQble8xyvt32eE+WoO+NuyVS
hD6Tm7g91daG/OpMSD1jKwpWdr+O5RtDxCWtcIy80TKtnHaCqsAX1dSpI40CLiqagA+0ujiFUPqZ
NXIxf8l39KTu8GVDW2tjzf3a9l7SK95NxS1bX9S9InnH+hBRMFJRHo8xYQE3mG9nKxun3/pN16lG
4ezApU5LV78rwufFLg6Icet+sCZUpl9LlJ/xCDMOG7PvtlFfn+Q/E66lVUqaZSktwzdK+8pCnZz3
9KscozN+ndwD9nYkme+sSmoNS+lR0nh9Y0ajVGKfS88QHmBWcEv1wNpjRUInkJEZfx738NUsyIr1
CYP6MY/mvP9iD0kzPmmYYtRP43Cy9FREvoa1TAJl7HaVbjwA9RiM/8WQwhi1LyDIiRdQyIyDNaFG
JM/xwSBRjJwNQ61+O+r+XcRic+VOykXD5iyvN80kfLDqXDjyDsPctnI2UGIvogFkbLvwm1jIPe/+
i+TZz1OokguomBuvTcAo1XykElace5dYORShTCY8ZFaMzInIu94I5RCSRyeL9cT2iEb5NnVBWq/8
EmzTRHK+7RMlIo7v0YwTPERM9szBhKMPx/38rSwhqi1fBWFmhk1oqtk85wUCiGF5Df2cld6UGkMU
Q464Rh5L392XuDIKzFsC9nxpRgeUJjFMEL8NuvGDlXjAege9Hf4kQnE/pL4ILPZP47IDvnDM1H9F
PALmZ8GU2mRooJRLG58uYd2iCpA7fbZFgk8cfMjDp0R7qse9TU+qfrlAhnXsKcBy+4U1rIHrOXKD
p/rOcdj2A9878zIaFZRkkGjmv3YsZQ6RJkMdG0ieg+Fg+YHbioL7kiMm72hjT7XApkA0cEt1IR3A
kUSheN1EXy1oXa/5ALaYnbi3cduQtINzukia8dojOROeVncVHWmnwLpRD2ekss/P26QSKIs3fusr
AyCRW/B/mk1dB8aTtyndz9plpfKyvvPByTPyAuiqNKzLhXzRN6u44JfJzc/rZPYl2bAcNa5beh+9
IHf4+RNWB3siS1NC+FTYEG2QIvkoufEX4KoMabObe7HjZWnsqM4JVw0bzoimqypbwHi1uZKvMJ+7
A8OnJtbfKvvUsBS+jv1+RXpYdIP21qIhEUt/zfb0up4vjrNzt6l+YCWsLDus/+1f/XKyJ8DzLb+l
MRhhIMHhgxvKvja4h3jV8SNrQhi1wKhN3PGXsyEWE04BVRZy7B0tUPaoD11+KAoaz8Xgr+6jFkOC
AT8+FhSuSXZFUGQXn4qZKgI6G1YEeqq5oTMtx/33eCGzUZIFgGZg1fjFLXTEdsT4NrMCktyhjsqn
V1IPNb1J39YLM9jOsqpU1ZX6BrogJEqI68lWtWP8tRjXP1d07/5uzhM/7tt8wYpr2p3oPWMnj07S
dujt+hQkhd6xdKCx0MMJCmkFIRIufs9mWvbxESSJjB1J3FQw8KwkQrgOSSpD677gzVV1s3RzEHXT
K64zGV6mue/5ISa4fM+k0egKvxzYezpReJoR2J4Gg5ewVbNbCs0Y7cfxgcZhdlF7ZmysUrzA33qv
rLKnLZiZWdnCWaa+gSrPSw67XljkTW4yHZkUbdJUYAlgj+uzulImxhGnXWGauPYu3VtdxuseCAgm
ge6+IdBle/cGDWVE8h76y62I3HTWoKLQ6eHsz8Wgvp2ErytH6l01epLpLLEO5p/sJilUYLWql9B+
p2S2hMA5XYMWnTAewB06hZiZyOyA0AUn7Ju/zcllmwH07W4Rabur+woa7TcWDUpjzEJR27R5ZtPT
r3RUsVjqKMBRShuZR3MROfB/jwASe6MR+EftfmJhekzOSvP2oWBtRwg92bWP0CwFeGPYKBTzwUsg
4EBncvSMmsOxdrDwjzFPV7IIwzAtHziA6whRVf9iOprZ7cRP+xs/QUVakKwOoKEKKM3LlsP5P7kD
IF1WOkSolbt1JroxHM8py1nnAbWykcWwoCX/8Q2cnVrwcaraio9nWBvHF2rxzyk5cLR82zOesfUP
wOZpYKzggImNbwr9TAZdFFTX1aREYOs0yyfKQQW5qJbcGWePKd9SGTjYWNbFTcnOF2n6ausWc5Rs
1nPZNcPD7Tat/DgTJRpMwwcg2c2Pe/x7lyDIqPBHQb6hplfWpS3lfmpK1Qdu80sFF7KdG3Wy5sk+
M0E4d1+m1UtjBgwFLMm1QN+pu6eIjjju7i8CpoEDLzlQmLGZbFkMvHi7rN4x59qh4PCPZuYTY2zx
TZJaH5WsHDrNd+7m+QAReojdlAzYOcAn68CNIE1/riuKRrnMUVkaJWfxMq6CGEDaYZlmwAS/gLk0
kIbot5ETox2x2FpiakrnAVG1frNsmnRUksRaeV10NMcU4vTPh2gR+F3J5xPYNDdYxSkY1BbmL/14
vo3y6Wp4SRD91a8T7myb/LZxC7Nuzt4/x7+PmoNnkqeyF5uQG+QuvEXfDcJdd1El8jWK54ZliCZh
FUafU1sALk9rMSg/duAqDiJX4r6L38foPgAzWP4NrRyMAND5HPVdMHnfWFOHpC2tkDORQL5t/78e
rWT1DoKleZa1BnF20kF3nQNlhtTqzvaVFSKrcUqSZrKIob8zcnS0f3BK2xnhc35EbJ+4EqRsZJDG
aH1g06NPGA2wCJSYgpfbDWPHAvAW/NoBJYHkobxIyFsBdtA+onW3wjhkrw0yTTyqDyKULpUFHBGz
+OF7HQXeWB69K3TE5R/eW7UNNxUuqfE4cYEpx7/5aWIrx2ewbf1dzJz5NRNGnTgok1HjrN3+Sp8n
B2v6aV2snrCNfxatee8cez75fDKAwU5zDAXZkJsTA7pCfkLu4JW6c3I2kMlfzlgUPtyvf2umy9d0
YBIXq3nCJbwvWNntx7LFGrZf3FrcvycNJQaX0evpTRvPliZWSfPn0cvvqK+aEG+WAWlwesHgg6N0
0+RpEImHQuWYpUFnTLLrJUb+1UpKQDSiAza+b5rWyH5+srFaXOKD1LSlQKwH0vVg+5MRImnoBl56
sGZOZDD4y3ZUfOFLarAIwxOg2YKFm05NsdDTNOqYCitqquNaiVkoM6yBWTF4xQpOo2JLCNkxhlSS
27TllHoOAK6Ks8he61tKhYBVFsG+z8vc7gTscTko9VGH4Jr+uIGmv8ePVSl+fQljZVJE1q8W0Ff2
zwi6pIYekpMg7bAVnxae3lXnGUXR4O7OOvtvzpRW+kbsm8/r7hhqjBOUa02OIWtExazVWuHzM+M0
BUmlyGdr+1nRWqvpGcDiDa55RBZdBLjNW4/SENSsHykJCGyaJl2ZmqGBqnQrDYjMC+UKqOVT84DT
6xPHPYbgW/+ibjaaPVoZF1B1NbTHInlvpaBXs1XIeCxKmIqUACVlMxu/DpsmRE2/kz85ZSJrkq50
UFJhs6RyAfnCpUcoJ28is3Z3WSiqB9JL1LnNDbzOU/N1rYvsIJgfBNWmI92g8TPIN25K5B4ch2gf
AAgQLwBO6q8izT+PnbS4jI6beGdC/jPdUcaWlprlMOK0aee4PzavzXHyQvwAb9v2pRQ/ZziS7KvY
Oine6aNYYVqm1KprU5w3ztULSNul5qtwBMwGt3lnY/E6jJIyyKQU7x/thSzFYUVdg2iNp1xRAyKW
x0Irv+Z6POZExK6zceFn1bOZts9zixklYuNSDIo7dmcKjxPEvUPNPSzkAa/wtIIvZx8sf9iVMwaa
7r6mVnBRVj5OLa36B2qEkYTsioefqU4RxmRcHk1NoJHV4V7EcggsCQHn7mbcEzWYiPDSc9DDO1yl
mJv7UdNBSNOWtpce0AjvN3koBTIdKmKO2TRc3QVhdYcoQkJgNBckS9wiY3rJJZJ4kSmGSf7zjfc2
uxM8R4SyqG0DfuNoJ6C19tyiQCAU2kJw23dvL+VBaZOFB8pot8dqcxha2pNIF3D7o73QTonrx+gW
jRgVCXhB5mSnP9nW1KKHct2Z8d51WI6Pqmj+PGPc3ZQHHDNZiDRfryAzXXxXK7+zBu8KuMiHD2u5
3blNBTjNMqJecpULKBF2Jc/BcHAtGuScvo4sTXE701uCKivq3IyYaAQW+3pZNqe4sqYt7d57M6tg
MfhE+pG2XUZUDd54bA7pHJCv4T/2coN6CM+cFswsYa1uREM995zzO1mkSU0vYbTb+IeA0v2NkeiJ
0oqCONFsjh4hNHZfuf1zTL4eQesjZJswwC9Lj2f3jABLw+z0lgIWkt3ShgTjVtK/ozwVGLXKYBjP
LD5SWjEG5Hq6t+vEX6nyxqT9ZsVlIyjsgTONE3tphxOpd1MYbaGPMdRmfJiwLVwnlbEu5joS4WLB
NvBmnWCmGeBmMDiG5hJgHqqlH5BoC/2yyuJ2DLF766PnRrnjyrtc7szX23LGwG8DFRp6mXv1PVqa
McI2YLxGfSN9cgW9mFkf5KjtswNo+0Jwl5WGhoUq6JEHTWl4XSZffeu2CSwMhsqEkacD85JjKSxl
VmU58/8F5lb6b79gzzo3XnGRcvgyzCfa518ALM7v2E5HWiILp2QSq9Zu0DfVn9r3whjBwh2bU3Yz
GkYeDBmzi4MTRccbZfoFQQbM1h3asALZG0ZRzMjtwCV3kWQDx8VtF1kB6AeLngi9u80MWXyxhiUC
uy4wTpyf0Z5nSD4ENcWzqT5f5Ur6oCy3ohgMYhtHHKvK7OHmVUJYtnSX+qvDBzhqQiZcHEfgOOmm
+N27SkI3Z1Gq4QUqv4SjkdDnfiAl3lkHi9n81L9zG4kyi2OdVcTbUU2GHsBGluryPRWo76TvjFT6
iV6rwBmih5B2sqd4ACbY33X1C/We0iDi1umhoHhOdNyNX3SWXpNeen2EOAShr0H6Dfv3J7HVLeuv
c82HxSwXjwLBsShAfru19d4XmHRV4WfhtZZG+89L6BQZu43bZXfZZNXUORZaUN9jx2hgmeqAcqOs
mPmhqmIINCHiynxmvn0F08HW6WFUOEgJjz2/5acAeeVI/Rh95AyHeID+wCjl4VLjkKgmnnHK/4rr
ts2aJ/vLII9Q3rw7V24s1pSJRkHZhFaqw9l49fKweRNES9ENWNPuQ17G5zzm3Tl7GU0g0RIDBjL9
OKQx0xvyjCz6Ot08mxcAAL8Wsyph3ClGIddEANVY8KIz8uhE28jPiayBijmkZ5h0l5SgtODnei6m
Lwq7sBmicZ9Qq6QH2IOhknE/BsKXo6zP1xv9JWzV9ajuruErI3YjMMlfqPdZAYOj2+GQ6w8Dv7va
dKeQOcK5tlsagSAUIbqQqdGh4Aq5vEnqomKzyaRZz7tfItQaV35ey4hAU3hI2DyErB/ZPeI/WOjt
G/M/XYPe4QDJZCyy3RoLzqpaiAQxM6077vscHCYQ1QUNYzFADAF+ZVupx2wCuSCT00RbcOwk9jK+
loC8PYRjCWwnQZnPgKbGU4EpFITUb/WsluN69UVW7IHq5i8cCAwTw5VWmMsHDmJRHuTcLitKs5au
ZLwtRqs/ui56KB+LRObvuOgliXkGjwCcPMm6jSaK81AMimuyDX8NTD8NHGmFiNtysSUlhbllyc2X
Oud08tHzucnYYWjH9aoo3rW7jkAG383rIXjrvlIAO2bWZ8HEw/9KoNOcl4HOARGi2lp+Ncd9S2I0
zfzdnwLCcA24vmqs5evtfwhJIYKq3lHQrvOdmN5PG0wodQ6pr1rqYgNiGZjz53mhjheDbSHeT72/
AA6Ny3kMx2bE7nH1aPiixit6E3iaGPXq/HKeYNIGoz25uXpEJDxout/ov+EI7VVW8IBhpPuDCfKt
SRfhOloTAx8UEmaooLzcXIpviPVU5nKW/ArKirbMN9NPibisfWvvgzJY4trpLJDVY+59AUb5+QC5
yl1JKtqb1Y22ML8IP+PX5Z+vgzTncnerddhInSryWiFq4Aj2xy+W+nYkC4Ls3y0VoUJhOYE424Cd
zbm+Uc8FwPrQkW6NfV6vLofoHqL+9/gFUTfOCcB+0FZHf1ieFvnwDK2i2sdDdPwMaljIwes6sbzy
n3oGloa7uxU97KknqtlGmVlg688+oSFy8ScVFKgQZtmRV66pliFwHWSLmnRYCzr5pVnpidcD2EE+
O7Dr6a+TjgdflGx8aQuRaS0GZT3kdSGB7nD6lwUD1Ozg2VYZGkqw5guIemUmmy5O2V12L82SBu30
7Qa48SEuNDf1PSfn1Wu57uH1UjLnRRlTyUJNBsjHmppgC/3+QRf7iDGNzOvL3q1HD23KVRYDgOdN
DstWPl3UiBTTWIcTOD8kM74uhFeq5RGe8df63PeYJwcGnhSrliNe0lHr+pdRSiUIIc7wozIxyZwt
lB9zy+H3OW6v7QYZf5qJAhKoakVILzCZT3R2xBKQbAwowncfm6+2TGUs6ntAFL+1slsDHNF4J3WN
oC0YPIXh1QehyAvbJrxS4Fo7mzouNRWJt3QT31SCG6mGyGzXtqDegT8HBqE1zVeWa6anWT3YV05D
bL3K5xJB/O4oqT3Y8edZtZ7Rsn4juy8Wa4En7PylG1AwBeLNN2SnWK6BxcggEtvv5Kr2UPnyxrB7
EE+fnvK415rE/HP8TTkhdxnpPjb0fgZr+uIRGZwMyJJXpvb5Q8gkXS4tPAw4hH+O+pdXMKVhmIti
eZ3nlOXRCvNSFU7rkQCJvtsQBMsgcN12SVY3Et1aXvs49nxN5AVdJQO4qDkApyxZ6tHsvThMrJ7b
YREq1IMGTlKdD5gCc5AJlpSrSi+iznkYfwb3WYCe8HG/uGEd2DKEys1TWRdT+WR+NQ9iQTN83snN
c9ZqCAKAGmxYlvFD/BZfzZKg2IOFIsKl4M3pFwCDFQe3IPGAjtZuEurRTLxNAVYN9EGix0wKcqRp
ZDWEi3tfkvwEpz0VGE5hQNS6AUKeTxXJxQVcjELEqO863SJl5L8R9VXlkYPh9tomGTsAu3T0duza
1hrcSs5ZXZRLj2JXCzWBLRM4NSr5HA5n+FC3DtLZfe1QJq1uguXc44KX1ZZuFzQtTuj/NbL74HrF
SjxOeHQLWJ3vinbIAgqGmXMSwmtrVP3G1W7j6qmwm3LboZUZQxeEmABwvl/kY0CPW2HWLsmR0Vf+
WHn2agJc40qg6qeXCuyW5e8PqtYveE4e6avubKQlIiQAFh4JBcSFcaakXGkapzMnJ0NDfZCeMt7A
oByRYn4bMkYawcI5Yy49vAr2zQ/vMvoEdNV5QMzJllD7LYk5pImRlrbsEjxyilP53dfFmscR8tS6
aj+NClvChiaAU6pn0JL3Ozl6l7dOhId0q2Xp429smhYasOk5SwfFeyvvw0JGfWq1N3my5sUJu6uS
HOpNabTLw9RYF8fL87YKZztu3uyvxggu8pEx/FaDyIJJZFciNotkJzO5hQnhILb9glZZ1gtg2fSw
qJ9G76omMZgIPFX+3WYtUqDmoi7n6xR2ZOJSQLSV+t02kQSPXySK41kAIsD9UkV3yV5+EGtBTi5q
OpwYioocbL2si1cn8QRqKDPMVGA+xfqYbFcbJZIkSFkE+WKqqYGRE6GkMuFteb5twBfrzbh1R/f6
cObwBIs1f8PWd8+jTO0Dhyi2AM+5vXj7+NBeTMxF5Sm2U9X9sSZf8L0EiXoyCkz11d4/5+UELTW/
bBT3B3fR2g2+/GIBTbmF2OcuvXxeYok7IAI9TfaEwz0GFeYdkSRwrUkZXpX+qB/8wbKSYHjSTjDT
ywwVOOWCNeTh+bQVV0+w3cEJPlLGQ+Ri+SxOECeRNyXRY0nwo68TnS7vjWGieqHBaEt38Dqz7qFg
Tlj8r+MOmwzDziXo7uQ5z5a9tdbBhId94M0VQ57WUYdJAwtMp6gU7hbhDgVFEN0ST+aMYV2dXmfG
gzqYjfX966aDFU8NuX0NZRxfiGCp6tik3FBsBl5XdD4jRiot0wtoAZ3YLXEnDe9QBozBLCBwGwSU
g9cpKqec2APxsUFvuNNDNpR5hJ3jAjYUtXkPhKsgblZ6hxAp22AqllTFuZySeIuI/XJtkFAnK6W6
+VYAgsV6RSHKuL5qu3xy6jqCq8g+sQBbtgdfvX7uDMzwK4RqRaX+COcyMx7XhqUcOQ++o3k6NON1
/4ktuHyqi+gGIJOcQYtiiCcZt0CbOMNX86OpEOIkzTT0oVgfdjxk5sFKmJrS7CEnE2oxp3KrAwqG
n7SCjw70pa6PdO0vPZdFabGvBCkp4t8DEt5F2mEcjQsr6Gys76EHEWYUT1h9HWUjF7pB52K/snxe
yDDepe7XCVkEcLAlAL18txuVEsL6z4EQnpo2C4Qjo7k+2jHR8n5ZPW9U1aP5l/UHgccwHTspl0Zg
XbE6/eusRyxD7FRAuHCQadzVFAsUaIUyhqr6UGOsHkJ4xk8rQX7PIQQ+0sGqP+G6pOz7wml8BTJ/
G5N1f/kD6q74UVaaAMbPrlI6wThfniX3q0ZcRc0N/HckQjDFXLtpLUpRXrfAVoaRLp5CQ6ic9XWE
CV08g2yubIEj7U519gQHBmdtzoCsqCk45/OZ6QpIc/8l4GzbSFyUZ6WXoUh+MMlRoMBhP4C8YvB2
e+x2qxz8dH0yebtxMlYV5Behou/enUZHt1z7Us0xIFfEMuNLeRqK5rTzvZjb08vDe3RS+U1EpQaa
GNi6bRp0LXnNCcUTi/HqWpMrtS6CjiBTeE4xqBDDYTZBwM8zdQ4LQtavTmEwQy6Qrdo8NcOs/+zA
Xt/Kh5VizfORMHw+WRYVntMvYXYnLVUKoMGZ9NMy9RCIGzN7dLftVQvtAOGr89t/rP57ERxbUdFO
Vxt9L5qp77woTGkS7suNdBiUu451Z8riww9dxqMkrwrC4u89lBA8w2SNGgWqdhn982itRDjCF970
dAMeHC9s/LsSLqVR70mJACwgXv1ANlU45uYwNyaPID0ocUGDMhVr49LKZY2ytlNT8tCnRvmlouGh
mTV/eG4GRv0U0Ae7USt5pMBGCtLkTU+xKF1qygB0LVa1G7FEkjTS+4PDErMKampf6Qupsr8LwpL4
CGj2Xqq0TdE2Qvnn+kBn/m7Eb1A2BY1aLdmQaxao5fNmTBCcebnpqHpOqtahAoZ0LjC4QoRfyh5k
Qgs8uRyaF5ngh/abKV7Bl59kePLgonm1vHt+C8hrGPyfWgDdt1dOl0tHtMZviA97R5iVaOET5mum
msbHmtyUpCLNhLBb4tccNNv6nk9wCymUz28KJ4A7TxEdwq/siKv77lrTWWZ4LUoeKv8jsqsSntGM
W3rl+k/8KoMrDcWFBTz5mBlEq5BDB5u9vlNechc0Un0Q5DYH2ExJozzih/WHBnNt6+FOtLTParcB
LqNLo+WuqIt71JsWeurNC6Qv6Qwxnkraqs4uVQMJEimAzaBKa9phzO7C/Qt9mDVqV3p2x/mEAeLT
tqhJawOM0So7K7kt5yT0UX20xIRwT7wq33Bb+FtBskIqVnbH7iwRcJQnj2bNL9g2eKQlq5Mtgh7q
5caPbyba2znLieUmnnHrv3CEgMWmYDRtfjB0NY40sdBlrBnwy6crbBW89Zeddpk1Al2xoDCQMvkJ
0f7vYrd10Ui40uHkrQtqQ4qKpgPRs8Vaoz9kfi7BGrITcDCpHaY7ImPjBtKX7Bw6hLps2s66wCLK
3cJ6yd2GKoGKjieyAsieuYGInzgduS2uaEVc+ELdLTQf6gwf111mYnMgeIssbh4TIG+f0tVnbjHC
IWlnGXvv5aLEgRk9OMeSTvmFPojumIrBpUbixHStMpP2Ye1xKuvaVxdq1p29mjB8Bi49ysgs1Kdf
5yx5h4SuRZdNlU5XHFf94y9KiuVvRvw6iqvZY281nGDwVJ88w0BlMRllpL1pSKUtvEXIXNEzPsJb
TykzajeMc+vDqlU7GG87AYS+NczuG9VuVt2YRhcFIk3gzzQ7t2oERmhEyhFB9SMG8CbFU8X0WOCz
YwhdAUiMdidkVRUhQREBwffQ8Y0gfAYzpRO9B63Wd0jVFJIxLHisdd2VY9IMNfTHrYlTfBfDPszf
QBnXO1Tlu2AnylmHciM7qroVZiC5LFZhf5lySCVOzqWf9TXC4Ns3HLiajBznAun/ZtlrEBOZvBwM
RT0qlnTbK/sxSW7VPOIKSju09MRcTmknDSB8kHmlSeZuZvLQn2dzuI3JDon1zJZZUFOrVKP5E7YM
KWgrdbS19Vgzhr3CwRyQoc2bvRUa7zT9zHyrFdIJk/48AkLsKtPDi5tH4IMW9bVMoS0jg5tIUgS4
xWMjnrmzysTU9szwHrXwS2EXalm2DTLsvXa1IHPsi9EfAjWda6EgjiA0O7i1jWm74FaXvazsW+V3
uMc9oSId1HEmU6k7pLckYVqp/Auy9lE6HUNMCpje7mXghsM0GH5+PRCu0btmqxYTRZrFQ1PpakMt
NATC5eRWhLkMq/rQVzuxOCqwlK3kwzvJRCadUCEgYTOzX4LS8Hj3hD9tjwa1XXbcxnB0i9+KxB/6
R4L2/LHOv54XYeOZSHmCuTIzWhcg6Kq3+hfLLIUVZ1kjy3YA3xIGEa2JfD/105Pqz2iJkjjdkNaZ
F90XIo4Oiwb64fVjqe2ceW8AqAsJm898N9sqTr/0KX81wheXFCxmq15+s1FroNeg1LPhxAqGCJ/R
AE4UywNODahh4Q2GJVuZo6aOSeuCKEucWwnf0z2IeuXZjfImlFbNAXxrGukWtEiLNqu9E7tVSRuv
TZDkT2ZSquCJs4mhaDbrHsFMrsZTkDuVMcwwNGsHRykETqcTSJJTjfJzYEwqbtSl2egHWgfRmqgH
Hbt95gHobX2XBMSoAntta/FnjKol3VNEtUHGNm45Xr+CUVt74wY1VNEOBIDDkZNAC4484K2Wu8te
2T1NhAXMaDA8z0AZnFTBIj9s4shTpvADDLTlPGT5DcxJcgMM09cvlML4qx2MsWRd4utn+ScNvQSW
EDkCvLfC0TLQRdsjKovP9fOqE9Vy3OMsTb/puahw7fU3wl4RrDdkFK0KgC2P/WyzaM3WuAlgWOHO
AL+R9e4e3b6CtVJRfuPXlnx/cbUNjENAly3nw2rH1pFDAY8cOcXQJ7+pTd/lUxoyo3f7ZavpNYWI
fGg3ipzOmPHQ8FOYXWqGiswYopQ1jfIVfpatIYbQdDdPOP1wxKvbF0eYbT0DIi7r5ohx90f4IbfS
21sZs+3GKlThjFq4/5jNSuDFHsiyqj2eujcUabBqOE7wkWk6pz1JWin5ck4ZSHRop/xysBKDRArk
GMy+baFyMXFzcInfqsuDV/cXU6FvcGjXwjAZqy8PoRjgYA5beRs3gdeCrraWTC7AyzP5EyNYnkaC
f2VuIR9huoC7o++FYIqBe9D6RdHq3TKDzl7UtOqAmT1/y1rSYjQonucHWeZdBxnFqli7G8v8Le+F
SmZCCPpaCxPld2PHv6+CaWLuzFWCP+4nSg+J+s6crfvgJ7xTbmCpkC7J5eSk4aZlKvcDqyGTGUwi
tiMqaetZZM79I38NZ9yXqc9cIIaw96WZkv5qAvYmLKTJbz+90+J+6OVZF32Q7BBw/AZoYuTTRdIW
9tkynGWfId8baXpBvqZZVkb0cwXKNqAhdQWGUFybrs98LsMD5TMIMg1VpxCpqyC797m15TYghQnx
gf+xPD0//jpG1mPTog8et8HH8218jxhts4Sq+FB+Q4VAX4Os2/1KJNprka7ht5f+3tmp4Y7ostf8
ePzbDeTIcaeiwJCQigX5bIUlzzbHnf4QUQJ3Nmvyvbjv+DMKjjKvJUp0Av14HgaoStmrOur1lIC8
oGouaybm6wvVLw8LdYIBD7Eds/OXt+hcG6ZwJ6BQ5geC68e+yXCPacTWBuni8bI6iicfe4XnvsFT
awzppzjODQ4WAW2RJWh/IdZGgoyruaydUKFIm8gEFzSldHWWC6cPaJTuKOAJmZHHnRyEgf0jjOf3
8IcVBYcTYxiMpiZu5zHzboepLDffBf6uYWXHtZIrqKBumFHq52xE4E22kKulRe2fN6Xz98sWvCqy
1JF6mxeFXYL8mRCx3PYV/dstkqkd609KT9a5H4IVktwCjIhXtZcJzvPwzeBgU7NYIv/+JY4/YdAX
OpOU6Bg08rScsKm4oejRnIP/d3JZuMhm5Z2Euy3HE0RMr4M3ZERbzHaquI0wc3PnBD6Zwkcjnz8Y
tsHa9mx3VUuOwj5Zpw1a+IUtGf5+SATCghZrmKIdgobFxjWzPllIbpF6nnuy8vhZH5BNs80r1nJX
fS+0MHYP/1ok/SVMESdJg/B+7nMrlia0W3Lgbr9g8hAhNSEC3ohyggewCfvy2bKJE0NKm0XMwBLw
MSnKFf1THl6j0UgzetaKFoGNaJslyNfmPEKndkaSC8xfapj6yRFM358Q+z5vVMbGLJi38P7bDDAN
LczhROMa+LOuEpcr3ZYxNjZwMGkxeuBmZ+09rhS2Y6eMK6jzcExVYbmg/Y+R1UR1J8PXFB9+iHMS
hX22FBJKzgJ+8hQVUJOgHjkR2I6G+qUDHnNanyGkdrAP+jCpzZUNEphynrsDzkTYx6es3pZlw45b
vzod+uKSIX5AttyR3S9koZYwFoord3KmYtB+gcuGm0NU0hNhddWFVimVilE2MBqXYOSt/CN4jQ9a
sLYv8vJwZ7nYI+h1XjtKKBT4oAFdA+HF/jCojg5K6nz/EU9ywa+cGN+9Y2cxVTQwkkPaNbeC1RFy
1GFmO81PURbEEB4EiaoXTc5xgd+qh1H/b4XXoHqW5nolAe3bDVQP7mE/vd719GrjpySKj7vFDgdj
qMvhyLgM8HVrMzCEo6zbni3NLtnCLMNnRubjt5dyqsQRTiX9y7V4+V0zOjQizkk256P4nJ2yaFvO
hYxTLRTNYv0n9Gm6lCEJGeeX3z2xMB4gWh6Ejg2tQAMubJmZlLrjZzECQK30TFK1gGrHydVJWuug
S/CT/6ZbK0DfeJGWs/+HExK2cf6QOSwxtKHn0ZM84zn/g6KIBYsYp3QzkvqsrdMRK6kVHuNcIr9Z
kwfHqeTIQ+RECMD/9oIid20WX34wpVLVjOrYpguS54ZdW9pnHF7Zj3FWBq92cJQ6XT+JRDka4276
r20QjwSWE/zFm+YWbJiozDEefxiprIpQHMLwab+dkgEms1B35xLj+9nhacWVwC6lHZkAsn4LIR+B
FmXpVjxq823MylgY7qcRmlCq27duMzxOIkapdcgOyqFJkZ4AB7PGBqZeliUeD8yQPWkQuxnEUeFa
zl8cg7IQUZ4+3woyM27oegazkpw88zr6Qr+5HhrG/xnFTZPZIO82lQwuCvj787peLzjz1+ewmAIs
xNBKuYwxMgqwKDTJ19XLJy7Sp6ALo2dg45H9ZUrE0uvKe2bBnXvv6tp7vMCBiOplm2DOtjs0bU/+
eLqHlID29CaPvCQ3N6EhCFi+/dgF8tRlPcPM99MLgC1diNxaUdCCFxJHOcl07MPnBtp+3wS3mo1R
c2uTgbXJQXHqCuBd7Wlf0Sae+BTbhnrf7oiOQalFXHsnyILSbVQE2p0uXW5IuypcqMEmL6EbPonE
l7/AtL9YlFU1vXHJYMha9SsW2vJcirlgNJau4iqyIPHzwX5nRYpK+kYC6BWGJkRTy5D2ZGfkV3TC
icxOltbYa2GmB1j+e8YTfH7QOKIGr1q2e24M+M1/M6cUnA3qce4Mgb3U5WhxtHgnyYw28ATu3/Ce
dROkqE7u5fNY8vezfudrpwuQXW5hSNv0iME4a8g1M7wecnJU+J/ydtFiq87m0kCJcos9WuUEOKXr
7Ec0q/ZLsN1X1la0hKrsA1LUhgv0NXs0upJ+83n7N2jfIMckOEgBxrMJsbtyk7oM0GNEL+gCKVwC
S2+9rIHm/gLyfuebARz2D1eKY0ebrmd/TA7NsXdDzNFwviXlr0v6qr9K0WR6ZmKQCuvzLvkKsof4
zR0Htpdu50tsJvFpQ/JfhsYW08otRQCnW7wdIQjGb/sZ8H7/6OABblfEZlO6ja+YHpAwkxg39PHo
kL0yM/LkPLkg0RG9/9/yr++6COentveWKexfJezy/vXqd9NXYcAfqbcStWBBWl6vVpFdqcvz5HpG
Omutmx+Qrs9dnB9692chZSGjUxDkDVZrFTQeRU25NYsXuO5NX6qfdxBoWRY2PKZc+Ar8bm8zj61W
bQiTgSFgfWLIAAoGZAp17bU7Lu6MemHfr8Yo3a1CXtqCZhYETiF+DWjSLTPqxwEVMYzmGKlnef86
3HvJZBV0uxJBppjeQaTGa7cAeWyogTyVuocHDMJJEkRvYh/EBmlGzbmMp0TDaNIlaPmsGgTbWUAV
d3KCTyrDKSENcOJNN3xmkyf1nqn7WTOH7NPaq3GS1+1aba1vYV1Kma0A7rNLOhDBIHV4z+MvgM34
I/qMlSLZ9/hi3Lgjj7QN0kLToiMaLzG0krBegzgQIh9UcGvrlmWYmFib5WJsdRAQ2qZL364v+Bjw
QL/TyTZDefcIqVrIs2NrM35HsYbhddKNb+yYp2MfsbJGSmFpr+l6YCRiRnuI7Y5ldfllZJoEOOdK
B5u8UtzJVoRedn1N5UFut5GMR9fJQn/cScD22ZUADu8zgHmtNTSuVIEXQMrDHWJEg0Gpu0NcSZN6
epaWaKhNZu9JZbB7J0oTWs/gCooVcf7+nGboh4+G5HMi2Gm5Ss1iR+OcZR4kXxTT4trqeS4IO7y0
fDIEbEfuk2uKkG0UYXLbBGxn/vM2HC4MqroDJFq/rh3lOIWzz+6ouqXXsmPDVDR0iQjhDm0RPvz5
KMq96NVbA9SFVekCvoJdzNmyn7dq4Qqa+TKcMAuI1JwivIb2VwYC6IfCiNy+97omeboSdsFoNClk
3dOjirHdnCv/h2RRXZYnbmGaTuuQ2KU+tfjAH0HITCcbBxFjzlAhaDBvOq5qifskER/JS07T7JLj
1nMEnVsIudHJ96JjW9YKy2YGiVGXC071jgmo82DdXSwkayLTR+kFX/C7cwy1If6Lxj/G2zEoQhaj
MGlpi66ciSs5ljGot/XyM4nHSv2ngaVpSwhmMgzIgu+lA2fghcTVgAlkcYSrI5pZxF69YgrK6gc+
p8n8/b0gSVSu1D+ETdG6BK6HjpwJzqC4eKtI096mQm8LYQMGN1kRmqYAYQgxBeSlAZH01mLiDGNu
VJehoTu398rc/ynPO+EQ1kER/vysdbx/tPpOmghDd6ZrCEZJGpOXpqvVw+i7EZi27CXyMJi1mqdh
+TUX3Occ//djakBD8h/WzArNKEMl+hhCTA752OAe0al/kBtg4KdSyILXK1QKzvhi9futQ/oex7sr
Fv4rHA5j39tJUaaULyavZEvsr3mFrrb83s8NSMyjAGvnpAD/CK8WWE8bz73siJjJa3f93uRIRrpq
r8VJMw9qeY1NAVjMxRd2lqVOKSqG/xsnSPr/mGWZ/0jLB1mBVn8+8pWyGu2iaKTCarv6JpGWDEfx
kREFzY8cqyHXbKeGBfT03Afc/PGpLk2BCUkYd68hcykcV3UBJG5WOFrrTcjelCOpxY5afXetu5In
fJHPX181FFoaNwug0+xZQW9pMw4c9/JISfa9p7VOO0u44ssSktauSrXtlA2Ig+36H59IALs0KDcT
BLTTSBs6Z6nKWNGOnVk48+u1jNVlx4sFWvak2D+mNOx6a7TUH6rxKgbeIf7AggX9OIGpriZbIYKO
mGVMrgVZ+G/Tif8nvft73EpiNyC2XGTl8Mzxfh+YGhH9w/HtfdW25wuf9tqxIM9SyfGGgwJqk5du
NCJFk69bbqoQw2U7rh7S6DgX8eJbkiPceKSE02BFQdabTubFJw6ppqd/Q7ED1/y8zq41c9cfvHUz
5YoTaNmDDk7unj/DGIi6+i047ffZkGv01tCpOuJ3pQZIRaFo4vqFjcD4CwzfX5aEP3Zm1Bmv7Kxa
Ghu3tS3dCKzQxHimJzb9jJrnCIaDZSQzgfEnT490GIyqzdRBbc2lKqCHWcLsfMghA0L0pOY3/+S1
slnlAMlWNjnaf/Ra4ES0PEUqvXcFPXie4KnuM3LMmkWJapCCVRi3V8qfi9sFlAi9at4KnP7fD2Uo
Tzj/DmcyaKSuPWg914ZcZGdmcl9wuLQ5K1WFZXqUnYmImEOF+QrdCzDsvN3amEpxnSMA37cNruXh
VwJgO1IMRL+RdWMWiY23FaIsRvVHr9c9t/vznmljY+/kpC1oL5D77k8Vyoogfur/ms8EPlmtdRWM
1NoaTytyJgHpyrWwwfHeo63vXmQMoofTHZHgzzIebBqY1jmuHq+YSSZGp31+yITEjKEf/SCW8r8T
lHpDz+OJrmNRKr52Bt/5H/CRGLM/2q+CvnjaSyHZvs+UaVUMaQ8dL6qsw1ws2SR6Ew8XPD1x+5t3
utO3EnBCMzWXa20B5n7jsGHNl/XWrAUbrnPWbXeiOqV/mG2JDaez6lMDmrOe/K0Sopsxf9hrvCr+
zSRFVtMZh4AwZr3l6ooJ27YZ1IocOptJA4M4Yj/RCGFX33lHP7Wmhqm7s95jDcR8QRrU4C7RJmES
aAFFmdIMI+ouZYnIcaCJfVAeJrFQ5vNbI1BWUqrxjEiY0xILmv3OnMIyyDIXxe6SSEbVmwhEvXGy
+4mSf96sZzs9MryDQ/U8i6o6Kk0uSepTD0eNT3+ZkqNWKbjHesmH9pqczUcQ6wMbkl0eWzuCA9GT
CJ4hYppxIMhvf+lMVZFCKgdlmjmNcsy7Ja1yhTtnWbDhlWW5kBoiYqypBvjjo8kTGp9qtOffyexm
yMa/mdjk3NPEycYRk1trJ4b3K2psB45Qepy64r1FTDaU4eE2lB67SSZXM5bGQL9J3g5XYH4dCiOq
xyh4kHs1fgXQ+1lPJujVRJNUnjlbSbQSeWCtm4i2LkOvNDYrfZLLzL02s9PPgdNwP+boauB9vgZZ
FetORBbH9cr1vDDSe0rVtzKOFl8hLkLUvakggof6w/Dyr2tOdR0Pl4tuK1Pn/wJDASmGVaJLOgjq
7ERzVnVRk9s+RGLjKxAy1oPKtx9RO8M8XNxwZe+9q2J05TPJ5iKZJvJN74xMS6/aeWnjB2iHMixa
wx26WIBoNCymIohls6uaTdGSLOwbN87+qHbW42SywK6aqBCzPlFXG8JAtPtsKIGqyEatXYObQOcE
5xAelkXlFBKkjqnk8/MpDyJsYwCgMzE1bTzAhI2bmmpQdT1mRbERZ+b0XDgKtd6DnoqnmJcCYhPM
VctM09Hxhj6by+61vNqonEUMA4NFPqSQhuwpcwgs3dXh2i9zt+BDD+HohtrhClaklDRg0XnSpi1A
FrsghsPUQLMsf2er888VRIXCQOjON68Esm+3Bk59YtkNSurXicE1+se52QD2Q2RTVfutHz0gLVaV
kzupznkD53HIOEhbGjy3NOLn4U8Q2UWH+73qLEOwVOBm/zH3obITy8yhl89FJ3gjvlvoLXr+vt1N
1dWj9XZfjdpIFmTzIoB3wGaYX/MVsg0I+Hk+57mSW2k4gpWrGIhpYFgbIdervKlrfQLY3URv4Ebk
W3OerszYaqvmxXZqO8YsHpyunyZJco8SAt6KtjZ++Y3mzJfMolLNL5Rggws5x/do4y8TirdFhlcE
fjjtUAiE7TDoG7ZBmWdtSb0Q2zFULOo0aB5TAyo7Z8F1TiPyRU9ywVTwcLRAOBABxaD0IcSzSns3
qAKYiXGFOgemuxqMJZF5iOeIL5v495in5BSAAjvdbnzHInchY9RIBpdZbPidrPk6MSA2zJ9hxSSe
kOJ4UjM8oYPKV1C1peNdHV5FeHtqkx/ibhA1SdefBLK59Lb0D07SwovZ6MUkw+5vWZXSL0EQXlUY
XN8e215XznsCyDUAgmJrP3yU6K4pI0+R4FdDIFeaL04wBXHGWCPxiWe+oSZdd5gr1/YwuJWmF9m7
TvPZ57nS3ThBq6rwutuwVV7e0iIFH0qjUukgAyJ7ZiXiA5RTMnl97EvbzOYXUSk03RJNQguBNaIL
+FWtVzcmFhuPCHaP5424ivShyHgTBr11BAwBa5DuBbujttiUwrWyNOxnXx7uLe5VYNWHRQ+fmjNd
amJ6DCrpbA3tfhkFVeM/VsEdkFmTds+hUq9siE4oy0Yt9HtW7tFKQ/byuRlTv+DCHQ/Q6RG/fGzC
+APF62Hqx7MBV9jc1vTzzjFalkr8/Nvr96gC26ugpTh90X+XslFA+s8q3X/Vjm8t//MFgn48St4h
kaKS5SFk9g3ZCaJsnrmGb4CpuIBq4+r77oVPvXr6veWvj7udoHMVU0Ej/ieHspu3hjH3tLCk+PNj
CI33F6ZdPdra+PeZQhAo8jtJeNvtgMPfCYLoMNpKsyu575Y/t07QbqnlHRGA11jrWWIxbRLDmOx4
MJHyAfvD0i4jc6H/p/l7eUj73wS4+sg0ty8WZ5r5gXBSMFH2ViwvbSjTzwYcCNGgmo5fzhrC95eZ
Y/kwpksOrdB0hTO0b6DDhTFQlbTbI7iATXYmSLo/ZXddU7OqUgZDeOSeXfkJffWUN2J3lHg/T2qU
JWjIIUwM81MuAbEtyuTz99aR4iUFFqWZ/wunSEJRTnvxEaKMo7szqQ/1xTFCd1Zgt4Rlc3Yx0m68
kec77Q+gbKiAgMWheIKufPXfasmJX9VQwKczjiDrMFkXNKxqdIi/lTW858rRJ5VY1hY3rsOJSFWw
sIG+mLp0Mubhs3tqDPMXvhmwnRcqEIqthE6BtChNX8a5Pu1yTfRq3r5rbkQSrV0WOK28GN5zCo2w
XzJr76PK14o3Vk+nwr393ksaUKcdXJUScnq3M724Eg5RKr1FqzdhOVgyiMjGNT1FR7vQz09vPY/M
2iJKikNEBt/SS82nxqv/wcVHAjP/C4R20e8zZab06kRZM+BwmbwYP0/ThkrhsjWqeeKcSKD4fzJK
mVqij4oPkmftPcIFReaPMtw4xy8cPar8Gov3Sm7kspzo1ZPtFMvRhZxuZhxzFd0sR3B9VbTwanCs
m+a+nsjmnDmpX4etsIqWDhm6qk0eAQreabre/hmYgwCyHNQHe7NpEl0IMtJjFzG1q38thECFklyV
f6SFFAmnY2s/34QDKOi5pmVswfwE3h8R5d7y1Wj8h6+vD2C4LBTRp5SfipQ6JpC4Abj8EgCI9v25
IOIzoHdkJ9tGaPgL7gNN39IkxhiDkRmEXAEccWvkxGS4E4hTD5WAP99PsO1a22WwKxQr5KuVZTBR
rqOtu0kH5HmRa3s4JtBd3fgE9R7wHZwTl3/xQ9qaMqXu/LwVr2XIm7ZvWsTcUf3GrLst3+iAGlAO
46Gkf0lfbjM4p1Nr9mw4JIrO3UMNsZZwnH3xkePlKmyQEv5FGKnerq5K+sW3jFmQN+Alnrf9PS65
GJtWUgaMTcYzpIIsi+zGpk3sY/xqhayZkkDNDGdiT1MpPIl+mxpYX4rtjXul1cmMqLj7TtTLSHPQ
HX8X2hMYGv0RpGto1nHmiNn4m3h20f10NUzd6J6n6dJIa+mkbltt9QvBvt+OM2A+vC+VX7mvGTV8
c1/vrGm5RyoFOpSJwfq0lgab8dBeVcp0n44KrFMLuZP0tYAg0ca7NYRUka+ghflQenAoiSut+npu
6r83BWktC6rUFt23uTBu5+Zh5PSiD6vYriDnK3PG60P6iAFw0EyHgk6uEC57Aq9X2YgjM+JDq5XQ
aphAeeJ0FS9GvtI5UX30pFcd24fnsgNeuGB0GEx75G8YdahlqcxPQxMJdoIgkNuFCsPov5+cLZke
e4LRS7Zckmt006NVFmXCcLyGU7FRkxEzyf63LqENOZi62SAig+iqkZ7p5Q2zMH9v/c0W2LEml1L+
aiipg29ylesDTcNgkRjK3oMMJDFK0og+xFiUE21GSIcoNpMdeNDjQx7t9ve1JbeFr43dIEwjKO7Q
KOxpGcbgUOGVoxEl3AfhDE51hQi6c1AzCkW8gb/JuQdMrgVuGpa4c3Mp+5mcLZIK9iypU3ZnYDUb
7EJtWSEUBYd7J5yULvkVFLebEKqcqCfSJ24mxZhQfIUtPlqNq2MFcHKGtuRbgFezRHvA23KpJ9Nh
/D7juH4SHqwZw4sXTHzhrJR/oHu4Qpc+Hj14umhWuB9LPcDtwSfY4jDYbGNgTrtg6W5STnj8F7+D
Qf0khzou8nr9qJGCjk+W7oIglszBu/s9OqBhMb9I2FS31BDrM2Dobp1C3Fmp78nU3zsdwuZPy/eY
XgE489HRaZitB5ecvJgR2gCVexLRTecxfHPY4Uav1GP6ihLqfkhVXeHAfIosXy8uL9ghCFl/UB+B
rIpny/ddpYjI8mRS4lZIoMRnisJ3pI1D1aTVjT7+vzlwCVXqXUFlITggsvced8j45XTHCqa+UY9f
cxA72btdlcXp6tOAskmMH09zx6NcGMwEE3Hou+28zd1WDGchRnLBk6rJeNt9+EuUXNhN7VqxaAeE
FtaHZD9SOBJ5Mhol8H7CXXFqf9rypfxDGnZFTO/TLW92En30VqTHqicFUJ28uKjyu0KksFiLdopd
T5lsinGGKaGl6RIJVuzc+3eTU+2RBKUssgl6o4PFfIKbVPpJAORKBQbKDDFhE5EgkDui5QV2ROvE
1cT8wcfNu6uyjWaHOiS1MRaSyTSFFM+NuplO7H+0gaE074fzP5hYAMuaZH3SjrEo444fQrHc46SG
gsmMJUIUz8XdWHCTdEa209/Uw2D+qohOm3f8KuZDE8lPFUK3XG5iZIar1pp507Zcd6bfCovJDhyV
Oq/hrxC39esE3kFY7YLxUxt4vjSgxkMEtTc+hdr/oLAbrtCfVm14yW3oaFmqMBbW7Auosq8Pebtu
R9cqAOM2C1KJPEiQkJo5/l4gVRW9thtGvdxMp52pauyyzWt+63470H79RA+yiSHui25CC1xbczuf
yKoC43j2b3NlYmL2qB1enKH4CVX95jSIMBFNPvbJGVg+rgN33bkQ5i0QH+cZM7KtG478P41vEARk
jccc1olTfJC7g0flB+g2/ma1Em+D+/aGwCl3T7Pqb7nNG6bfpy83RVc20y46THG9D7Fi+ce2CXPm
us89WbJ+EWDID0Rq4V10zSy3bJrPprIOUImdxstGm5RIq0Z4E4j4BwSfbcHDxrHY+XNrR4n7U6wD
KKPDv+qhWSHxnz6OWkOfZhoounUUUDOg0c014Ai2TX+qzHgS36/PhXQnK/oadHkjRHVKZdMgzUcX
MsqIYM4wCG5PFEUQKQmYfH3GmbmSYeO5qcH6FYGxbg1XZ62lSI6Ed5+uWk4RXLvlKkRM+mK00qUZ
bkKIukHITPTFOpSYsq/wYcCGqSojDVPjJrktfaI2uQ0KaFi5mJBGCdOLpw9kyGJIBG8twJ0brs96
oOdKfg8EQe8u175KyQkUzdAd5igCc7Q4Ipq30xTPcdkogjTRGPlgFK6JlyxQsFxhTQRaDq1NSPEd
husU/4tuavAL7B6GoHdAVT1JD1tAIBvuC/wuJkzFmxv/9bl08E7n0nrFuGlfeL2vA/zfh4GBrugR
wnzTlSjEvmWWVyk+dLYjwByCyANU+3FrVHCGLhMRwx1bYFfQgjJGqdRunH2I0jeJpqJuJaJmZmK/
xuYwCd6AEP8yhwCLwgyMsHxYfYrwfOCyfNzCw3bm8jSH/hxCNvU6EA9K2EcD5c8jW2AyQOpjuEtq
IY7Pt7HCWlHuwx5ExyzBmWcVTzIBegvolqhG6j8ib/1zfi7uearA6dUhXQiiuPZtgE0K7UIqsO59
vu78NNL2a8lBrl8giOewEleF+9R9jn2RD9JL/pHVNjGm/44LHQ+oFfym1u7U+Rq/BBaZILr/ip7f
cjqi1mdHR9pbp0Yok4I4rjWLcMD4h3yEjRF7pT+1f51pR8PTczYpn2lC9e0eUWGc3/IBN4BTc8+2
E4tmtsup6DCf06APXy1x/8s98EHgYgABVKjGOCmiMIbngt8o7Kxm35y/J6chuOWnqxtfeEb1wu1L
EUholLzuGaJOhIN0617LnjoIP90irnNS9CHUGOPDalVVcRfjlwEb0l9TSYymhAStoyTnJRhyA3pb
G/K/WWB1Y9/LwjtS6fHB76qja/TbtcwFbIqJeicfqGGIXAYccSjJtdpHAZPy09uqQfMIeOnHrfzS
doREvAJ+9KzOs/RBjxaQgjmcDOK18rg3N15IOP8zPcZ9d1cYlgajrs/tvVAz4l5JDzOd28HHjECo
i9S9qG9HLz0UFgUQqkQ1Eiyh3fixEZNmMWmZX+HkIetjM2wgm3+CAnDICLwEwpFxDJgW+h8uxvgE
2s7MDnCtRz9HCtPATXZ661QdRJUJAJAVgO0+mbqagNwa18SWmn0JajZFARixLCAOKvrE/QJFol4W
9eyu38KJ7yuWm9kEtN57LXRTyXOp1sBl5jW1YZmMAJKE9PQu/P1iKawTdK6e3aD9EtRbX+zHMNwO
Kp/V5QIHxN1cA/jm9NzkI1WjgQdyO4PUiVrtzOE1DugJRp40Abs96msUr4buvux5bRcdCts5idj6
AheJ/2XAEwd+oGUlhVraM+Vq/NUDPXUCzsfAZiAbgytPepG17hBDOJvBo6IC1g+TWcGN1dU3UCmB
Rsr9wBDto1HufgcMZnFuBXxIRvh8GaD1SLzV2xDVd9YI65MAMIiiAN56oipm8VuN3eaLLC0gQkLL
yGqvd/kcazOOJ2SwUVRytPpRGVYFR0kldGZ7AhMxwCTl7lashOspHzvi+uEj2Lmf8oOg0TkhZOzL
PkLK6GNPDN+eIs+sEUZwauY1Oqn41/0ndv7NC8nLpSpvSlHlQHPOyo1pNCk/BC4x5eOMb9N1mmoy
dPgs6MBj3F3DuHUwEcdyGxTjC2+fjht+yhpRX/7oOghvDwvftLVJlM2kMICIMqCtWIDuYDbNIARV
okvHjPCP/BrC4GTw/OCuybYjMgyJMMejuxoEh2rVZGK5Jg7Kh5Q8J8Rw2CbdKm8OXt5x9nU/6zJh
87IbHmIrU6+9FnJa6sQaKMMufctdcrL/anTLjb33b7ZXn6p3c9oFGR8MfiopdTbpzWKAsdvr8Gsd
FnlvfTKU9EWpPLVt9a4oA7GY7OEEg/Jz7Bh2rFyMbNaMCYHyP670mcgfxhgB0GzZbKLmY7tojcGA
h9SYcaKeLSKvplWjKHnbuXkpCnSC9aeiOEpbqFmGhy208zxQHXz3nD2bT8uTy6/Yec1qKS0Q/n9q
AzZbES0K+ttzWaCoD5UQ0KYQblb8el973ZvxM+CO22m0AKdMpNeppIolqzPcqNmL4HNJ1V+utDYR
88v8Mr+20zneSUSbayY4DfPoZVgybPbUJE0CTl+apY+A7jVjm5Iod2LIZuxFM5DIsTIcZd+38ewf
Z3tky6GNhlXrrC3zke54EVCXcOx51pTjwj8UlbdIw7Aa9EyPTg3aa3AHnd4rS7NX8TJuHnGYNkFC
HspX0l5FGuQBF8WqMURM8okyzZ0c96Qsjv1DnwEFbTYue967X4AiFb1AX+pNhQnZrM/E7oOx9h0e
o3SWM0c3NNUj9bdmPSAhQFjg2PIQcQjIwojw20YabOHNgeLNpzNXSvT3ILMgXIhriVDuJqQwOqzr
Sy8iLwR7bEKDSzDTFNbxyCJSrfGfjqtIhghML+qWJNPdR3xCpUP9j3o98FrccgiE9nKSWjRJIhVc
VaJIp4mCGohrPXIN+FV5STvsSIqnR2wncxXfak4yUN6kML7nPrFZy5geP6QT30am/t2P5ER/zn/U
/M/HbEADRejZoEMc8fo/iKnqt/kZ/VFq6J+og5Hat3IdcQNIPj8ya+hV9PLLtvP1VCV2sxiJC9EX
rtfYlzLaqaYxYZr18FH58exjQzQ90rSp/6pMO5FU4iwmuLkyueD+nDI2WTk9i3bdM1UC0kEXgtO0
30ElNnYzlToynYSwpvw5XWcAPbLYmXtx4H0TR+1wz48h5fPqwad/KNHkwLL2iLuvLeCUfyE4IE6d
Tey1OK9hOz/i/8NO3RQ2CAGnSmJJKSsY4PHwHCvXU0bfgj97DfW6Fec3u11ljxN+78tA+ggEadNp
egszP8MvRBEDcFfBcO+bhWvqFcHWp4Vf7P3B/8UFYFiAzPDxoiXnqura4RNrAcoGd4JF/UuxAH3s
dCOq2p4JBNorePaRNRkKnopcqTkiygWDkQqDGPStMWWX5OPvUe2Eht/ft9By95G7x4Ei9hmeyNSv
itKox0tq7ZsCL52ZortwQtvluI/mlFqmKGCAGn/NGP1xWZKyu5UeFhjAM50P11dAYk67tWylPked
MOHBrxSdmCviNFAFd1XUNM8jDESAplKRa7v9tAZ0aTFuY5njYXDPqEacfCdQZKy2qfUkvl+ll7J5
HhXXgdcA3XI6PakkF3yE9Ee3f3cxph5i6kayDvXsr+9aPcJKndOPmvruIUjxVDKhS6bRWaKZwYYy
gEcRvmGV0BljqnmTTioy4DtRWPCopq2QktoLpRHXEACre786skgQjcyx7bTUk/UBQAvUMDi5/DKu
2HAvobCFsO3KAGpLnVNFpzMkLI0V1gk+KHwqtGnWFfam0r+yzWJK8tHPJiSSXeQ45zue/ghk15//
mYm/OaAXPfd1HguQj0ku3PEkTBuwh3pEMDT7mip7iIhu52lSuxaTBzXVMOPB9iEj9hpoc64HVMDD
+jwtOH6DTWRKgIApEFaKn57SbWhFVRookeqRPm9+07RJs56WdO5qjF04Y0TBkr+trk8Kry4r3LRM
BOMDHtWESjiTNwLrMBVrY3FUni4eDJ9kA2ACNT6KDSDvExvYx53leTkJlrt7PkGAWIMPT359B2NJ
GnZZEr817F9gZy8TNKD4jd6HQpv1h4aH2A6Ip6hw2JZ5KBXu50Tit0dK0NFl69cbYDk+sPQWgsTB
sSyfXL6dJe1P5BOBSofcpOJ7CR3yd91Q+RhenjVyfoEhXYTQdupCSW4mnRTAYOxx9MU/Ne0nSvRW
0Ds2gP2Aphslz0MqU+o8O7EhV4HCZ4KLuYTNHGyX3VGOVgGGyvsg+T0laAFXTdB+zFanQDHoRAq5
6cNC60mzHTCRzJRak+BLGOlAK5SRGEoTIclPQKq5b9ivNtoPfbj17f03xSiXcHe3tnN/dcyVToQI
T74cJZ65kPUz891sOnwnXxiqhOXURiw7KZZYKUgjQcrv6024Oi6evq1bK3e/a4VTyla6eYlkkQB/
naenbZDi9p1VuZYrMlA4Et+XHqLX+vBe93CJEaB0rwfeRtkvUckbDjPOmADw5EJ2bZbrKoTYDIVO
hkArXsD00tiD9QIwjT/hPHZ7zd9Nhe/tAsusIJaDnwA86KdFd3Fg1UiPnKATxM12SqBuJijCaXmj
kM5qiqhnL6rQwuWcFgIWHnHDqdr/KT+86sBxc2JhG1TW7K0xYvRtNCvdKg71yTqozAwOjJHObGCr
ZPjFfCvW94DDGT5n9EPD2rV0grfSGbvDmr04nR1kR/FtoweFHV03QGG8F/Lb5xo3KSaV1e8IFWEp
HAnaY7b48F8ilGEDxmb2KVYX8iewBGCo1g+50IDUIKT87ukTwhe81RLX36Z2GgkYchgV+qlS5dvt
ijmR71QApm8UJO+BDQbUshq23kpgZkumFfTVFSHpdloysI7VAjen56BBC1XTXWr2kVkYCgdRqhzP
OzQyHab8M2GPnboLEqZpn9zZ8DTiwRAawePF9AO8kyZLtE+dnSKw66o0SU2er17o1O3IcjP+0KsH
XfcEunNOFXDsJz/mAAjp7b9B3UXFxmJD8Om5WI6dPHu33cGRaED0cHzpieTqyO35QVYHuMOkRxgN
olgHb0ISZpFRHSF0+nK6NqOb046L4xrUFslmLR6xhv6VtbwTbjLTNKGqSrqH6s6L3B9JYgOoztAh
OLwND9fxn5d/bYCa2ir22rFjnShTajWcULl40AhCrxN2nRJ1JSmjllBNR7N+8+oRUqZt3sxrOu94
90zeSxYIvQNVuF2Ay+s0sXT7pZDfZmktOyOJbgWvJmpxHj+x92nVI2KfjJJWdic2kVepwbjGpguN
iwfNOyNjH5YbSir6i8ZPL1sNCJJN+xPqerB2KYJtdEV7s8QPLr/ufIWmbHM9EO7QYaFkGJ/g0S4T
No3qh42Swu0cuHC8RTXapq3QJZVD65K710HveLQr6Yu7M/4CTJc0Wf1VObsjsrPB9mDoJNOtRzwP
hhZmqipf9ZjLUKDoZKKs8C0NtWMf9Bppy6fX945xLnEnwWg0haXuF7Y83uHUUopITfBsdUHKEyR5
BzoI03Pot9UgQDiGpdbBAYHjPzG/hdi3OD4ksK5oHJhDu1LtK0cXd1khzwCahbAczdNkWn6fk2QB
wh7O8xIgQN0ubj5H+F//9S6oQZMqNl27D1ae1g7lPbeBVb4zqxBZf6G1aGdvKolPcxugUYFNmM6L
14cUDjAk9gqZUt6ua9EWbPLBobhLbRYNKd2/bY4bdxreQXESxQyWeyioT8R0HpSp/uCj9g87oJnz
vWNqLcjrS6KHIDRbmy6yMUVwcBPgQPz9hHA9+YGhXw+p2e0+LNkZntmw1jMLmsi5nUkvHSMlI4MV
VmbSS8pskb9yyV+1zF04eFV6d08XbEhe2iToh+uwAEMXPPLRMbw7HA/y6Ez2MUQlWBSdo4VqBPkK
ND3OzCr9R5xb6Lwp0EE62VW7e9Q/LfqvMYbIyaJLpD+BGOZopp4o5Stc5S31UHeIYDz3Ccu15wb2
Z6ajkjFeZfvGSlx+ogu17JAekek2wJwqF5SG4VTpDJwmF7jzVRx97VUY6HJ8nXKsM3w49N4w+2Y7
QdVK1rMs8iEFt0oMXx/gtL16mqqAgAo+7yiI/2c5GvTd882EJGQAnOfRFIcdwg85UshbL6N4c8LO
W01Ob+bAWX+tJH08ZYSzpDl/LCMC+WJBdT5FiyB6DGCcxM94R5Nuhvhskwfem9jCYKovFP2Xa6o7
b5xQorZp54HO/0RSlY43zri+mNvArp4Agws/+kutVf3U2C3DIevtJPnLqy1vegoJPJm68VNElN0l
PqL6DYnI42v4enhWowZFwEomaOW7HjvarJ/wD50mDZ8e0oVX7oUESEnPIMCCoobJjzAKOcKSBkGY
dKerGuVw0B/tCulYJWO6vBmVN43SsPswj2Hx2ixGGez7XYiPaGtPMRv8LPo4zVov7bifZduwA2Oy
oqWsm8I9ch24UfZ9OiEj6WTtZ2FjANk3fTK+oxjwqTZfzlG01+wh+szv8ZKgnTQViSoF7CE3nA0n
rWs+17Ak6qDDt566arki3IbJcA2tPWIPnHr3tIbQZ0xzisIPeilVyEeJh58M7En5kjTMNnoUlew6
MmosIfmqzqx0t6t/g/UKSi4ZJeH3tjabUEvNWlfi5Qv1PVYJlVtp1LEwxjYjmj4SeRbzkNcAtQhK
CKJC3GwQTZJh9djVasGVapqZHPnOtth6RIWZNYdbYEgP6nqS2jT+byzaN63s75xQhMxFJZu0yW4L
42QclImq3hquIvPCzoInGDeaYArO1m2mPg/ii/h/vy+l2/yKEo0eL7bLV3WvABgpMTgpyox8+Res
uG2OxXkpPft87h/SxLwBBpV97DnVg4IMqQk8Tbav5vhallDUrR26blEF/8a8NYc0gSxl9gMX5/or
+H7+JUCDeh3LPIBGHVHYXnwumEkp4eFdXW4qZismiD0l77lC8ZPwP/0jGp6l76eC3UJwkDIxUzJL
vHRyKpNhXWn107L3UI5XtobFqKrLiWy0Nkng6GqPZONSF9v3UenPRh1VEAAVkcWMgG2TW+daKAJW
a7Z9U3VHsY+WDH47KkHYn8hw/wTlWXUmwpj7DHFYwISQrpYNzc131lvR7Xp/696q4F7H7wTtPbi4
B+ghNHSoNW5XrR5F+HaOEnGFrdP7DTgXck4xXZ8ayR6XPLxvY1ELWuDuNI3EF5DJSUjs43GmXM1e
3hvaQOv2PuleAjbFD6kZA0F4f78oMmFL67vf64oUQcCwB10yBfU0mUdOh8iBDZ6yqmQ9o0/95UdK
8s52AFQ8r4JtkF02j3fvRKLA9DFZzwgWcQcfI/FiiWVOc1HymDYFWpXmszzTQyidW1nnzl80pWAu
kJio9WUkViqkXYCpQRKYBwxSeOane+a/TCrCDPWLVsSPDZL4RFW944pto9BDrFO2cKV9f+W+MVs0
hoV34HpSHWPBl/b4FFWbrU2X2FN98tLX6da7OWRyoLuTrQzFDtp5/04vwV26lr77jVpkBGwQXe7g
C40K0G2O07eIMEiojCUmPSXRUufBVZIUGBUJrsZaHq/2r0lFyOiAExc5VGIEzxaFSWGwXBHatRqM
K6HgkbHwLgd7alCr5h88rV2iNaBXS4TQiQiQ79wIUR8uHWGkl7jDzvxi1vRKmYQEuu/ol12meURb
dOBET5TT3PsZMcvlyy2DjD+3LxDakgRyq9zXYexoDw55eIfuiCxjvxTeg2rHp6P35ERpc3bkbyt3
txf5nh6L1yRZQzUYj48HDYuNsT9UBKncAr7tb9TsM8cg6ykVo3u7TCeXn2n/+QEhlU2vxNhP5jj+
0VXkqS/6t7fRYFMeWda1uCl4VVoovLiqAyNuv/6gx/MlNbViT+hk+kVDD+oJTNR9PHOYAqfv6tLC
t4QHMc9X6Y7ng17ja3DUNc+EItRSHCiHjLnwKwDGCcgPHI8P24KyKDIFUrEoz82LZ2d4LImAyGRX
t6EvDbHGc9RBv3iqSXCWNzLlwxm7GGkjGgyfuR6JhMF5wTx3UR28L+/Gun9QajgZSyRjUkc58rek
Q+YFJgFDRmOGcjS7/BSnOyuVaEvJjQbqoobj2XzmPXDHFNEi5Si/WTtTJAaBu/KONWeC9utyuBNw
pWB5IgapGTBA/PcJSzwZSI0BDl7xLUJD6Tu9pni5T0R56a7y/LF67jxLQH0zoztbrq39i5eU//Gy
b015OuKD9Vn9VzvKrMkC7wDU0epBIXTSF3hDO27ouTfQk0eT8ljURgeXfiS5WrbPrjZJmxXAWGiD
3omD2k0C0kq6xZ6ItNQX0+4FBhtlY6ykZwv9PwoK9XSv8JU2y6H+UOYTLpg6hj93dSloz0RCz9UC
4QkM268Pp9s7X1iPm3Aep3F0PXyuxitv4E0netkeUbdCPM0FeykXeT9HtFYTsSuwBL3wL31vWHqU
1T6ooD8TFEtdd5BBP1WdcHm9PlKbnDvipEfA4nu4UHj/rf91o+lwtyugquPJEthJZ0SQeoUc1cHu
cQBJVbv6/rHey+vEX+j4nz2E1gs1bi2rkgV2JCPx0yFpk1XYcVot+HVRkrEomc6K+12ZO15s/nCA
CpnpQhtZlpyT9TkOc5r5NNzrN7yFx159L9EDGG1I9xryjQgcTZME4VGQK/Y9dMN71PjOUqdLdZxw
tqR9XKe8nVEo+nyGZdGb1mi4e/+oQ8xnOjFkFsRp1RJkkyi7dkMs96eDB73/zbSY0ns3KlR4tmfq
d7m51uUtSA4qZgJUigPsfVOpzxnKOYOLvu1a+tW97+mMxTVHlw5t1FGcbxV25Qs3LBVt1LkBcBPT
Dc3V/4+bzfKXhfs6vxuoDfVZj70zT7t9ck0mDP8htUxYjbcYIP/VE755q1N8sFiEuXDVjl+qkhfA
IXwz0o1gkJD9sxn9dj+6vNcZz/3DtnN1IX6b6qgqk7d3cDkQE6rFvYYKFhFPQ30IOi4lgCn+7wXV
lvUg15kuvAhRkGl7jsdlvZTG2flHUHtl4GzhvnhO5JOpwy1o6CXzZOpN6Uta1PvNNealzZ7u152e
52sKy1xYJn+fKzTUbBvfLbmT4kduwcCKyXESi3e9enejg+2oQ5aQDF2kNgueKOLN8syc0EfGSZ/2
r4LupJOvwzHCsf+t+6f1tsNNNGEo9/ZnO9Gz5rLO99H1onS3EMhBE2H1FuO8giWjG6fuvWWAc7Pg
pu03h9YrR0sKDwAvbJVig71W+RT3ZchtKNuwSNbpWhftysMURkm65r9rSrpqiO3BmclFdcosZfA+
7VOJbk7DYCMj/tmIIZL/4UObEoREqMcwcCpgvRnmTW6vvzpRMF0T8xQxi6EktMyBPyZV4EVHZjAF
A393j30xbLJU8+VgbnPL/rWkN2eUCL2LRgWHRV9F0G/V4Vw0eQSqvrSaVHs+PXPmZqRFA5Ittey9
4wlUy0yV+aMu3VGjmdjgDcpnyzl1ONWE4ypjOFvOlh5uMqqslNOG68lUk9UP/g1EpCB6NZDCFSOo
qc7roMcuUDj2APBo1GjmnEVOGuhfW3CeZwshgnfSoDL7e8R5gCASrz0z0NhqPFqSKLXKISBC1M9G
sRaTADWi9QttdHr0yfVP2U7R/3VVEmugKOPXrYuB3qw4dZeDxFoetSf+GVp3wJYH68FyxsdFZVPe
ldnHYDh6uyQsqWvFSLCw9LDMqAJ26CYxb+H3oNPTHrexpMICUDqSrl5hPpBJzXCNaavAdRuoHQfU
98hCO6L8XIo/Fv/CtXNU5PoeTYBUnfM20MgsAFuILyJm7+gXOgLgiy3NX/AE2t+ggrteujLJOjpn
L/rIOXPkJoedl2c8A6zVGymHVAMvPMbAZAd+QdxkIrZKdgsASLVs7lby9CWLhH6+hnGBDIQUnds8
ZCRj/0W6DUqqlTq8kJggQpcYDSq0hrjSyqOQhWEpLNeCx6GMwpWACihEkGS2ZTNJJdowgv6LuEMv
96YFvBUIvaJVHHdjUDqST33Tt7aPn7vOMmokflzF7yZaLWnxSj4trtiwY7DlwvwM/sPKXXl+xr1q
/9HbhLK8hcd7XZYpaxtCtLnK2lrzxW/wxF4jt60X/mRHkpEbCjheexfFiQVVB5ct/exE391fX7hT
lpgqf/LpDQUT3/oPt+1b4me/MmwBt4YSDzkQfQm/IIxJRS8ncHe3qhB+a4O7Njc5+nS7nnGmmsvS
YYOK5dRPmYgV6epJ9fGXIjLgtglyVLBZPbV6a7XR+CRxuCrpWpr2/vjJhgzxpFu5q8pTCZCJTRPB
NCe1K/ADZM3Tzdl8MVqU2+PdnYZSule199KF8+KepYWEYw28Asb0OidYvxgwITwz6IqYATG7ymsY
ZKyvxz/xM0RDsw16PEi0jB2JytYc7v1FmlWd4XSsF8g/Nf70wPzhGarhiPtIphP5GdnJinqaH6Ay
cQDuASrlSTtwEJ3yR46/jBw12FPhI+Y6wWBTM2ljMrt9sYjLJdC/NIisW4J0tgQYm+r+eUscs0nO
xzO891yQMn80Q8mNAuxTjZDud5b2Lto9QcBa5QoQ+EL75s+7zPe1jSBR1MBVBH9+Kv7/MugXyl0U
jnBLpgXNt/kPrsEdI/24phl5tiH2eKKufb4ThmanD6JZ57UC+lO7R+LQBosHZWO0hbq4zQG2O19+
Rqpl8R9IBZhx5QDV7HQ+6gaUwpiJzgU/Cqc9/vcY1THOY3GHpw3bFRaBbEZKUtwtpbqIu0U7VXY8
2Dv+TGKXi0G+e8a6GbVJkeBEWEK9bPk9aze8sk+mbBrPl9jlsaAejWyj9RaklBe99oR3R7HKn7L4
QUxl40rPSpooEHTR38TReC/Ex+6y5aoXOZ/zEUGsA1vD4OUlidXwYyU7Ph6ujVg7liqjEpJMIJCh
U+T6ydL6ef7yZ+S/6Q8GvV96+QqzAwcdFi8FJB7JRK2Q0rUyHlLfRl2Uq5ahwxekYz38zZOXcEbH
0X8TUMqHkIK8R627QZF+pc6u4NKjS3vBuflESlLzJDeggROgRXVQtjgH6yctBd5MApyTeMBl+UkO
NJXgrJLq2zfDc2FxANAc/Qjv3b8e8cqmtJSuZEmnqO1sFeIZMPZAbFcX7ljFLDSdbylVODqQdKOr
MlKQF8hBMfgiyCAmtU/8CynyTry7hbu/eW0c7G3UxgpPGFH1TIoRqpwKMYuH8HdEVBHsfz1CUh1R
/oSJbFikBQ0FIpj/3Cg1LMFh33JOfvwUDeCLAvWfmTmVghzMcEvri1EDh1b5y55z5BP5hMR3k00j
TUr1nkNh4wxfOqGZ0+Kt7ah88GTQfwodU/Lfc9Owj4ag6Od8kJTAHAA/aOxIHVnfzv0YlhE5LYyq
8ErfdUEhdfBfqA5BTLASFTzyMcOoGeTiEw40P5DeXMOrKFnJ9alVDHfgz6K7um3SjjoM5HR6sqJ5
/4L76hNkOzgz3C4q/UjxoQ0aBC2tyT+6yI8Pyt1o8lcCJZllouaYq7nWQ+6UkNAW7QdPoHQCCoDa
RWXOCQ00HQFdeKwR4cM6q0/P0tNmku3MGILUn+FpiblALepzLdmF0fa/Bc12nNpWHjyroWe8fLhu
kta571Lx3d3C8iaAcK9xHM3IRy6yrc0C1yYsDS9pYrazwzDbXDAtV4oZG+WZFRNnl4vx647t/NTE
1pScrxfBi/Fy5sNm9YHQb6/WBjRmDJxxNtbtrAoXpeOs0ywcqpPTCCosQts7NNZ6dPagvI1HM+Lk
igcQhfZyDrnmm0FMn1GidkOzcf1565k76MA8L5IFoYTw3g36ZY0OYHhu7OluLLFaFN6jW1ST+qae
z/oC1HbC7iTLn4V6leYsZfmOAlbIP0RUvTIvtyaJNwnRbDxYWpH8NMkVqwCfte38JJF76j2FBOOq
o1d3UL+9fSYbwTNqyd/aame9GxdfeuCIJJDuRFp+zb3vTvffduSvR1aHNyu4T2PEeEGSGMY0NgJb
6xeaewxSWoh7WNjQTRcyaEz8cJOzrrE8c2BBQQSPacISU69qSY7vtLNcUCm1toTWhj6Bg2t3CbfP
ymrTFNJACCa1tcN2zMeb2iaPwLnJIOWyPX4Yh1WIbdtMQdGMKdKLH7jdFLw+luYTirJA2ymDV1H2
Xdjq7HxKmTi2z7UT+jXRxKsLaKHF+BKEHtZlGSQI9Lnp9p9EHR4LF9CJIECJzIoxRylea4dQHmW4
4rjLX3hJWBoX5nzKpk84sv2qk815QplDyTWQK8YHyEfRWFI+CWzl3Qhrh0sRWj6Zdwh1Nhi6ukvs
Tn8clj1agRljLskEF1IgNTVmXzvvT6TohghN6xwMvyxwOc9JpJjg/kwGvwTFxT3r8AYlwZSB2CMw
RkS3DA1BSQLFk4shWytEj4FsDn02G5JPz3cC+/HKvO0isPjilO3EJfC6Y3sVsYQ8f1+tlqGXGUNN
o2oqsWPyBkDlHYUCAVnO3A85lXVlERf7KyRhS7M/7x29iVRKfnD+FQy3PdCOT3SVukvYtmaOMVKQ
nHqQ7sssNVeWF9QBcHyfzykJky2TMwNtxOrCikWkvUA8W61p9q4ngxHEiPX2lLTBPpjZpPdSlvqg
GJAfwszthgplIUgeadbcJ0B58fYEmnAn5SvvWATWVV7N/OfZQl0TacXFSiCNLma1L4M+b2QfiQU1
g3oF79wBWtT7vvLJDiXeyLUfFxg20Q0vHvk8n8xClyJ7PfodTmKQnKzCBvKHHOPKEC29JpCJhUH9
R6txZVBTg7erKne6cAPnvo0PgOccmMMW2zhxPimmzU4QS2jGlhpDbycjv0qgYdSsTTGvdQvr5fSu
y5onWmvGiGz4xwk5bGafCwS6A9IZAxkqI7F1FLC/5m0uvpQFfAmQ50SBhvfJ2yIfn2lk7M/niLy2
2wbR6OcSrO9UaO5HJ306kGh98VlWPQjtMPU/vvVhucBCdxbGjt3Jasz6WrFP2pMzUtoFgR7sKq9E
pt/RRQzjT/BiqLTmnE3MZE0RYhbjHTA4nbXCf3efYYkYl/22EYHqKmHD89AlV4uqGG4ZCSHsXG4M
SZzAAhNBlge8wguj3G5eGzlqU61SQYV/recQ8LSwxuAAX5KI4+JSlqDB3rdnlVxwU1E0OZvxorcy
AbQl9yd14jpYDrbaxoiHVk0I+SPAFuF9J5eo80DFWn0pw3kRtILpOPzGr5dLdsLCTn4izI8/1I3Z
Y0f3JyNBn92qoHeODZ74gKTK54GT1hLpRBGZidvfu3L/+O96W/9QAuAe1Jv2dqtg3ifkgwU3ec8z
ns/ztIbzG2NsfWqstVDk8eAV53WGoveC9BbkVbMG28jLjeDmPs/+pVPctnOTTDv5nvYh420mcu1m
ejmkceeX8iLGSOgn2P62pBgdDvXZK4vGxiLGTMNaK3F/KDC5P43SZaF+Gfs1wNw9qf+tTeJksIk+
2fgx6NwPnWNDb9nGJiYh/t54YCsqIAhgZloEK2jPzAKwV5cQAEXdW1BCtgX71f9Jxo0cHr2uaUx9
fPhg7cSYNJt2hsE+F19ocGjecRWAjpLbm52MFm1pV7ZyoAJ3IIdc0DB+f4JSZHVtr0kvtBl54WjY
BhrGZlpshOqiUEyBQKNjWVUabe5WnfngS9DoEH8MT+GNqAlbRn0ZMM/eL/ezKIK8oTx8mt0kfTM5
Hk7e8Hm+tILmkANdps/15G/GWjEG68eaf98jUqyXW0jX7AKvhANnWXKihQ6FaOAwl6yI1JSfUJDQ
5IiiH2bTckHe5sLBwu6Im4PTmUOM56foi3EGl1J+Af7e9QOHma7K9N390soVqZGmIFKuxV0lsu4/
AFKwMgm7wcsYaWX+PtCve5s//9QEI6b2ychbIhYDfW01HGllvyOx3nQJtlVfjKgGZdS42FjRn3Xj
ObeB9tRlDaV2RBCMvzx1isqhb9I4EXss0zOIIteMGpFnVPhLoUa0njN26t2AqxCb8XoV5Lj6FP4E
YMf8rkdOIgYuiE14kMKbKBIB3m4OSohxtBR6ZQixxhZvTv1ZXVapgutcJmurNN05WVaLuHIb0gZu
KMZKdvRjzo3DSQ16doEi0tM3bkeATdpzM3obfAj/4VvepbeBLQQyYv1WBG8+sPIbWSXP48jinpDJ
lnpv05ztsGErss7C1N15bFwbgpWQGzsZPm0chxSnV6pTsyU/ipT/0oQHs1SGVgKPuPdNhYe0NGEx
hDrNDdpuIqGBW+7UfL7+S/EwOq1JY42zDfEIbUcMtcRLzutAapbDdDRNIwDVTEDFtXfDSDciapEr
RSEca1NIXpSPQect+JEJHwqKYbtrymlVQSwtK3zj9ez206vSFsbbsl9dK+c0aDSu4/vZaoF7iGLQ
PeDK/4W1pInMlk0Uw7t4KG0JLCpsG6BDpMqIOfPKB7GQ3reaJMYoYw8v8r1Y++GqJs6uB2D2aq6N
fJ5LbEaWD/P/tZd84tGEcRwnsrUj5YdwDgcLeMPIgH41TK7TCAOmfRUYxyaaYIOsWg3Ds13Eova+
CDsixxjjPljGR3iuAMzKpB+aefkQG8SAskmmeAAxCwBn8zCgI7bT518ZmzVyT5iLdGeIrwwM4h1c
mX0CaqPqxkACdX7O0VPgBqCnn/q0QlynlXe4bq40fl67sB+iOJ1PDkQPnQNFvRBNQzbIKDjmiC+m
P0YIWpPiKBItP+32qm0KaGjJXwy2hAjLme0CTcPZJ2tsX2rFYWZOKsMXzeEbaV3xoVGONTQkpNdh
axYEAHS0wFF1nem1UX8bLVmOcuFjTZtfVpEJCQa/szbZJ7Z+iQNClLlsiCdQZdlZK9OejzKDaSBu
yUAZGKwFx/2QTlZV3aMwOPougaHXZwwVqEVPrgMPQ1pRUdq4TE3NFel7z416y9uPlXhpOVo1V3I5
sJUTw7UOZkJoskH/se9637Ikx897rdSxaKoZMCoSvftAdKH2EQWo+nLX5R3sPOI0UIgwpABpZvsV
jeZPN6k2FTxfL6sLaYe7qyzZ4diyLSeCv4cOhmJArB+hr6+H4jV2KZiV362H1PY6Bwt2rxS5RpA2
/SI82MjC7cEzrAPC/WE06IpiZEcMlPwJdh/xgzEVngwl0Yo5eDbxFCs7M8fTpqgb81fuhexmuDmS
FE86t0WVoYO1QYMYn7slUa6h6ObREfxfjsEyMpaWhHVKtQAgzLp/kwx7WAZWpMwtWldNh+RhmgK4
AufgiF9vBZK/N0SQP3UXUes5gyH9BrwnXmg9gx36jeHbTkN55wUShjDBsfz4MCTHIuYg0Aj9Ncvl
ZofiIkRA9jwNoJxgM54UqVWF1JHSymHiyoCer8k4HtF0Jc65u6xUDUgrEB7RU0NcYvy4PmEbOkTG
Nuud7JE4oqGl/zZaNECDLMfnhSwCJHrF+TaUH9r+Vc6FXo9sdUdXCgobYgjwO64OC+oP05L0fG0+
a5uFCUFgxv36QmlFbHE5riTsWBD8D2bKSYN9Na8sZMkG3mHXa0hxk7irx6sVFCz6hb+UAzhz7P/7
MH5Abv0ls9DZ6XPJD4PG9eDQ34nB9dUpWJ7tIbmd+YUsxJ3WIjSZRf0zg8E3GamEzZgZbYXoEP9C
LOFItjLy8BB5EFDkSHFbemk81dhlXCudKreKsz1qmBvfc+P28hlp4LOjqjYEttas9kp+mfKf2EzH
29U5cTrdssGf6pRFiXB+IvC6PPjMjYZ0rM2tmDwWTrEWoHJ1S5i41/sWJ02I5XDB136ZYl/0K0CH
XklizpOHC5cz8SvymlrtMm4UKBYIuBF4YJ17Bl00iKBnoDUrWoUlOUTfntkPQotsvdCQe3i5Op8j
SEdj0SfdwVq3f0eaUZuAe4asexq6NDLIdF7VgcBqayvqD5eMjXXJa//JYnN28bLV/9Xh6k9YONZz
/oGH5Csx/OWxQnME+9JrcbaMRP9HcZwgzb8RrUW1RdB88ldVNTBbw8ZS9zcTc/73JlptOgzfrPgw
QG+H/ku5wUkdKrNhxg7Ar/aJuNWXwEL45jz+jW7q4tuohiHJjoPDTRwlggn4gi2jT8N8OO5jYWvg
iFFFPjs1WktW8mt4hZBATRPBejuJ3f9833+RKgxF3/L5ZjOowNi/B/NQwH1fF5IIiQTHgbaO2InF
rKsHXZ39ji7Voe4DCd2xNJQVytOM0NR80zquYqSFnAE6Uutfw+NL1u0BoFbmRhXZ7ETlmIJmVdNv
NgLV6aWptP0ZcKlgAS1DhTlSJvwiKrMuCYLYbc6NN09xiraJeJqJ7lMZOvs8n9/6hoZDhfY1zSTo
PcAYVRpLeVZpk2Oe1xgfQFf6Gey+N2jO34ir6IhLrPEJ8bm2pDyu/VnTQC1bLkH0xwAldKmaTY1e
nJduDI0swK/y5zmF2cHNnsn5L03eHzjYw5BgfMkZ4kNXHs8DI3kpOy6dCk3cMR1lBOS1GyIMFtEh
xHSB3pGyVTrHerucRH0Xp4sIU97cPkRyx7suKiXjbpA9lFKA9Qklxbv960JPOh4JavA+zr952c+h
oqd6iGEVTIvgvv4Yz5FFXGhWV27gvL7Y89BC0ydMtgUE3/4Z/TGL+wLIGHyWG8MB2Xvfawkhf16O
D57QkolujN5njMDdn1ep9++uHhwQ7RonEISnOmRHtavsQQiX/2/GzU/rvVGX5oSLZCun4BwL5aye
2N5QdIfyWq13+cbgUJEn1++CgnSHwhC6FUzhT8rmdgDWcCi4x+377+cewX2ZnH+JshYtj5X55eT9
O4iOxiLWoIsJ52uAecIYX/ZN8CXiWJGrllP91ojZLQ9oFFIklvCH/Iv/N20Yb764dqT1Mmz5beKB
qpQG/FpVQYnK0QsWYm89aHjT5NZ/ubuM/I2lY2fm40igqByKSwagM4qn9Ye7r6O/tbVv0+gDHrKf
SKPAayw0X9UTM+dWXn9T0IvtnKmQ3ZGwZygzURSM+PX66ID70/ELNV2mt7HoB9JCbHqjpZOAT3Py
IkfUGGc/WmRtsvqMvGuokXIOQdnLsKxfZVsyf8pm0RvLvqupFUYvl/CwfD/tMc7L+HrQi1PFwM+5
XArtfJ4+C8gSo2gG7NNUPvBjqCZ8Jt/jevfW+5MKGG25V54FZ4e5qiCoqBY4qHYWWxpeKQ58552D
AXcrgKjV+in8XmyY0ia8c1g6PIicLVaTwcU3w8EwQS17+my/Q6xfMTkxGXB2PkKikIwOvq0RKnuo
IzmGIBgcjGYLnPOZgpIAuufuyjRqK99wXnCGmDzXEDmEhRC5jCyplouCLTZcliYOaF9mlHx8bX8x
+Tj0Cq7M1yhISA8+mCx3VNBhtr3q4ySwTB3YIT3pI6gLH+K2NJpaRH45fxfeEhyrGVuxJYl9UAva
gX8j0UepCcaSWI5Kubx5T5NgVL24XpovZkHRNXsYwXKKqcztDICIlVUjDEBt5HJsh5XoXCE9AGOw
kPlun1yndwPmsp/Y6MuRyBVozgkQMaIZ8A84giB6bXzK+zlSXyAaDvEESaH1EGGFIs4GQqfLF9DR
7vAsQdXTB2czjX2ZeFf/DZrNXQLqTdOzmlSqcYdfM4LNHRIxTwe0KjrCgQQyPUpPFTWWnoMTMdVV
FQUPalNsfzcmpgtLu7ZihP6aiybKWG+lKUu7i6twnqXDhMbRt1H06A5r4mC+z7OIlTCbt10r9PJz
LWCUQvcl2qfIbGjStRA1V1WmEcYvCcX0bYlJDtIoLJ+nheiqj4gGlag13Vx9O2Wt4hIa8YAkmDVT
+WgLgXshl0zJHGLdy2xRVtAV0r2nqq1CDZtSMzVezCc5q/V/aura8LXzH3IkXSSZZTtqh27702F8
bzgNr7BUokar/31KlBj0EDSkSGp45IgNmfyBt6mdW5PrHpthjrxu9kYAGGk2gjsgSnDmJ3jhcWI9
yfbkrQ9YIBK38edOEivXMBcYKUixlYqWL8ObFqdMvnNGbpzvu288HZV2V9QyLj06sGyUR/dfvb8P
YysZ7n8YjG/nVJrV74Ny3rw0Qy7jflDUlvBeyZl2l7BLMe1d5j/mtcPH+1o382MiC8950PK3+q8K
qMaFXTXZYRFtrzHjNceIrFSnN/RsoD3duyYhWEynk+CGMIS/VkZwFQO3pPA3FMmJYaLL+nt8S+5B
oeomOBdzqHTXMefzQYWE+DKWMcBrg3pCFOU2IDsXvqZX8Z52gOM9xJIdZxWEAs4+jQHpr5P/4zct
gDlTjBUeQaj8Q/tAzCRgGT8gQmLRTc1NwoePKHRsAPUM60Hm6vtcZFJ5AC278IejvwI1fkz0qhZR
Pmrs+gRiZSTZNvQQDNs3v7qBvIMLd+cEujIBWhbQaTzW5HBXn5jAsn4sjPd7g5YTj3pYadJxSZGI
ryPVihvc+QBatOw3+kTFQvHSn33oaaAF9Aniw8xDc32jz1mhhTkQI9QDzqBxGkLO9aeNqgMv2B0Z
doacqhE0y+KEmgpWbZEmEb4y9khzZreibFIID6/Xe3TjFtpLTlUe8W0bxcYRnklaGp5HC9ezriew
5pu/7qrlwBCt59RLfpG3/sdyHRHUfySFXKuqQZYdrm1NRIfv8nf1kK0tz8+JSTdxt5Dqp6SVNHse
QWd8sIqVIO79DHFbD0YmoMYFYDSYbdejysx53kpnq5x8O3ePluti9TkCJ9Gp9/yyNrR4VoIW4xzX
rRIHKwP9CC/zBSbR7ZTq3Zbk5KXpNk7KLQsKmAJV0M3n/U5OHMO8O4pviaYv1XiM9Ebv/XaUXNa7
tXWjre8oeBr8I7PsONRgI1ZsfSsoq/PVDoZRQeES+bRKFO+vzdj/ceu2841fk49gjCvweE4n6o/S
etIAxNKBxQpMwqBe8T1EI3/2l5h4vK4j5LM8EXzVPMI/nvFUXpGyqtGhH8mGfK1hsk8xXmMQHjo0
Y+0UmeGasfiZaGDAxMUlSsRMmtAmqUlsrmvEwy76s51Xh+i/lIUPS5AsEORgHbGKek/2x33tZb/d
68QJiLnp9sSJdMZw2mEEGmA8xxs54HA0lDTVPnuvIDl0hHSORBW9Ku3gJLGO5Pna49Cvgt9EWaNZ
No0axPIa6YEFAog778C3TYWgHBog5pAgZLU/trjw9FMa0vUvEJP/ORwFZKcZPPb45slwkOS3pE4B
PZ+t85hwO2ROMKL9pt+jtYmIYWwHbRNOVhqM/cltfufVj9e4Naaf/ONZxTWXn1b/2KJbrrgv7D98
6fAL5o70YDdmhIvB++/p/tWRVyCTkca4M53wGThb3RtgXE/8Ae/xotepdh+0mQFQiTFIlUI3bm+V
PFRtDO3khNGnQxZnUpF29d+et0+tQXvTWzjwL/PUKZUmMssIbPOpq0i7jNWEeBJ+BogE7Ye5CU/t
lkFaEEL+89blXfkzOe7CnEch4z/hS8mW0PjFsFOoeLxnynJX3N+DeFN2patdbivUrzyZ57W0Lgm2
K1o5GlFXphXvxDsl5rnTu+hLnZoiQEm+xJQC95ePXnzhPTo0yRGQLhSZOiWRsGsKusdMbQBnuqdm
9gKcDUsiKdwNRtyWQDO2tmUZdsYf7XOby/ImnM9CTFkoORmmmaoI7owUG+EYoY+yEvxdz0of4n/S
v8QmZaY0/pBSzLGSkEsNKU21EmhbBQGrsBp76A5hs7gYRQl/hJRgnexB0/yWLS4Xt1RCgtb2j9Y2
VqXuqc2fG7TZlCp8jNrt1IndKrmMQ1q/ZxT4mKm8hmr4PvoYkwYdXua6pnWVmGWLgLKjz4LC8XR8
jmeHTs9wecIHwYn4rZABxT3jWNFXl82LJAWO6Ujp8unbVztREwgioP+c5QMlZgrJ/d9FTvqgNvlJ
cqi19i09L+ZVkViw3hQA0JyVLfirwbzz7rtaT+KiEh1mpHkhVk4AOABbCi3gush990gmI0WN9eOL
Z4CpVfmsygN/e+TAzgmmoCndy0NngKX38AJVW5qTjyEa8aReWgk24FuZwNw/XdF/v6k1G3FsIOBY
SkG/6XNbTBBePBe4MLCUbWfpOj4EQsB4clkSTBYzXy30bh+scbEQjwUT/nV5MEOznTSkGlW7Ghnb
IhDlw/Ae0cCL0POPL9hl1kkfQ3q2PNrbGATG5IOFyxA4AAcNEgOufcavIuyyrWkjSfaXi1lgs9z3
hzsp2qVK+wCt8EZA1rnN1Er3HvO0b6VGOIEQ86JyuVA8ZsrB0BlRJ6oDrEH2Hee/5kKMlhQwPHWC
fnQODA2G4o7QobGnHLkj6/WEQ/nXBIHmiVLwQh/27utD10bahFOLbN2yXKJzzBwjeTDigdxhkYw7
NVIR4JzYg17qrUuD030zJ6ZiRMFfzbZ7G9BcSKTXEDdABYTZnmafd2DBUI4mZ+ksUgD4/OH9ZZ0g
oXBE47H26C8GxIHPe17e9FvUZb7xz+zKzJmc+HycBVdHW2leFHNQ2bD15fXumNT6WbC1lQkI7viX
k4WWUeqADVPmnYw5+byLl8oKUClqvXb5OijWGB1TpCgXapF0VuhDn3H99CPc8yIQv5U9zR7hi8Ni
kP0L9/Kf7Pvw94MSXniA1lkBzOrBAdGWWI8U583o6/mfJK2/UPpwY0Sq0V9pR1ZlR/BcAXb9E9An
spAU9zAPXaSpvCyKjkkQxChNTgVct53CZ1gJDnnyL2Ruxftt9p2Wpn9hjUwtPIhe+d9ga1nkBVDg
ygHEJBVJsVt2GVqmOaATfsB0XsUlByCUKPqrWa3e3BFx3XimZZuaPHzRgrEHoInrrQnsOATiLoGQ
u7NK/+v5126rEvjPb3ShI1ALAQxyxOrfRZFcx+8RT2uReOaqk2TpszSbNUyzF3g7DVht7eYupheh
gCoLzVgu7YLTEc+5WqUmd4V3Lc6F5TsieqY5aN/M7CXJXlwPSAtF5JwsmlKaYp7xcHXH796FOJWo
rM0ZqRCp+G8dU76bnxb93hRqT+oLMXWKwVex1j2tkfBNq/hqP/om39g8azP2QeU5xRweIk1wXAMD
tXHczf4ELrBlKRmoza0cGzhcc1aO8t8HYVFDmmPmaGDpPxEBEHB0W1gAdN61WwTTrhsVMLICw4+Q
QrBnEiBmSHSMFnHt9hSjaVAAxkW8Pq4lZ17nnVGfbpaEJLXIdaJJ6Dz2JWZ0RAnStJI7Rn+1sT1u
1Lv/r46uGD/yvCyjoNWWseyiZJvIdsfmODNWhTjrl8SakYR8tilL5QMpVgnKh32AzZFg1pFsWakv
0UyKG0ISrZNvM2n0vJVNkhaYbB8dfPpGKb9p2RunNxpmJIydbthc0O20C1hUDBeAqrjh1G9gEKIO
kjNskpsumVxIGDeNRasR1rhngtv9ros2ygjFYdHQLA6txkXsDtJPYY2aGISKmqfUCkNq+mOk0rRu
nBUYHc+tP5ggE6fAIVf91mAOz5NDWsEMuQB8+JtjEwTz5vvt7yQPXkJUkdAo0Myay0NdjUIBMJkJ
MkB+itSflbm5UW5wAZt+ClJgBpX0bAoVAOMo5bOU7mjeu6nYj/pxIPcnjOCmRPcHksgkkMntFlFl
px5hKTVq+cqXFBgEtuJXo7IZF7bb4X6mFn/g9etTUP3OQwlIDJbJfps6PeUs9QO/cdyx9omcwO9y
OA35Y62WDKlGsNjo1KWDpS1VXen0MNmYqefFI69mdYOccJoDKfYPjhFno07G4+/MpVMFXjtNkCsd
QgABqtAC+Q37o5YqXRkHT24qxFThK4qqeJ9T/Wjad7RrHHpAh014VvNjrw40CPhsB9CqSi+nGsNn
IT9zYhedPAUu4yP8TV9kJWdKgGU5SksSCN2KE6BdM/Y99TN2dqG2XnlrF07o0BQq79iI4CXZjyac
w7MLSDkKbE7CfpG5bppgRH4w0cVM6CwZPnPOyB9hDWv3jUFfuMqx7MaeCokQTbgu7+FZoYIX6pDM
Zn4NugeRk4RIUMDOuT75GZ7Hyw6EF6GGSkydeBWturfcnFTIToMoK6fDce/+uh+erAHEXfu1+2ds
pBtsALZKvCAJ5xS1zvYyur6PnmlOQ+KlfaPEwPf4ZlprN3mhzps9jPAxwSm8fN8IyE51cVvZM811
vvwI7DxDLm8dIwmn7QUmmkmiP68um6Oia1W9nWuJjXhwEGtuBj1pZQpkUhdOU7uROTq21XtrQi5d
n8qwrgp8JTMSEQdYC7KQexVsRpKP7mDcyZ2dDVcQoM6TjOKP2gjCnBVsQAFmqeimVigffw61R/nU
qNSRjFFiHP2iGEny1Guv5zass1QJREC0xefRsqjLPq5RogyrISWj3wb3B1SrqUAHK2nDcTyJt1mO
T+njTi0BUqk+gT+qkxi57iqjKyvqOA9xssf7nV1mKwu/lV8kV9U5mJNBj7E1CA3JvPe0MZojeDIj
WOf10zvY/1o9Hf9DB1OvJPvpNVoqvs2wyd+k/H6ez92RFrik58t1HWU37c1vM7O2D7+w++/bSm8W
hyO4FGSJ008vTa2ZJyGc9GVevsKWF66llwTQgb258n65cB77Y946EMrEfERgCKviD9/DnvOS0nrs
/mScjsM8dgcxxJjV3wplyvU9ILmtp80yadbLRVotS2ZZV4zAgnXWsSljDdfkmCj3wpJhY9EcR4CC
51KhnSBYa31AOcJNl30M2sQk9/7oilyCNGNgvnHpDaQAgOz98xaBvwKPOPM9K9RUvVGW11PrQoZR
9XOF0ifqc2tgaMwOngeiRjO8GnpoAzibpGK6lrSMNuuieI+aj93z8SfiDViYwRXobaAFo/W9Tknn
az9PU2u2WLpLZTsjXFir4nkN3/dEWrL2iYjNEIk9EY6RnX+Fu+y+TSx0nT1my+2634VZleSD7Jx1
eV8aIJgW+hKNOfENM01DLLVPnjIgqUuRH2bzNkgnxvLW7xfCk38+1dkovCjVlBe2FLndKzB1j9l8
0xUbY9f1xUMq05K4lbyZ2niuj7lIppQ1bWkPkZQJDQFBJG1ikQEtjkUvWw8EI+QgIJSAgu8GTddu
rUi724nepwHrgeslxViyP6ZQg3DO1JSxRiABwvuehhZTGjJkblD6pVjJh954G3o0hPV8WTIIaxZm
7KFwSGu+RiyaLVsKBz7XUG/8IhOlKVPD8pgqwTLmRnmCqQSjivJB5K15UowASBk6oFGrdjBdOpJ5
w8ulyqgFgJyAcSns0lZQpYUMgXoUwr2NpawXCz4XRtLkNvF+/2uSunFoTeybRzsvn0xDV1RhacHX
Ur5Jetijch5+Z7/+18pXRj7bgKAznAnucoNR3cHOoYGUWbW1AZtNlAPcB1n+9ML0g/VnpjZ95wXh
J2i/k7PdHHcQXqMvehTxoxso9+X0ZUqsfX/It5IlET59OuLjlUAwXureyxGkGLaYbmOKp4v6v5AF
BCpaSlwoOrcM+u0kSY8rT8wqdQ64SIksrdbfpOFaB677h4lAR3jHYrdqrrAeTAWn4gGEdKLs9liS
ldugpeLZavkIGjfJFcvh+zIZvVsYg1wFJvzLscm8pKVoONZEbS5xypfEjLwxOMJvyRQqaMoByHXN
TZm/OrJDb3VSa5T9EO/SfoTKo3A2ncT7BdrTpYkEZ22lC1NqJC0slfsqy7wiDYgIaGgJ2AalBFx9
PRjTriiNelWK2oGMQ6kPxhcAF7CnnYJpv5rnlwB919mvoxCB1GPXQKHOU6D2TGI8ggOOCN9iXA96
ZQ9VJsUo++ns3i8zqlCGZEG5oScmJSVDcAr3kvPHCyS4qwcxqwTQVC90eOE0xmlQqIU5gpTeoXL5
jgqqy4df514sNe+YTVpJB/v40iUXnbQ8S/xXgYo/HfdHONP8ap8NtubzdK/hOIk4mZHtCJrQHMg5
cSb2z/aEKhHJWwknSBCU5aXEzEkxeWVPhxxVWKvfwU/rie7J3W4jFpEMa3WHL6Oc77aXfkoAVehb
VoAkfbe4y9mlgDjwAOhKPvzP+DS40k1pNIbXSPhy0y6WfgFtYUtTUZev7FaHP1ibTb7reg8OBV99
GA228+YPhMc2fR3di7KGouLkPiPn/ROKmOzcisVRPouHoRnBAzucK/RsjJG8W7KZx3ma16cskMrW
WkhPuEmLbbeIxfVFT93ClTcEkeR7rlGQ3ip3Rcti4SFviKspDjespYrvhHeEClynGQxV9ij0QTfn
1lhVtHLImIT3cqCkvzlmZrqsCJSxJswp7vJ4tNyEgLbZcSlZmdz5Hi963RwDp/RHN2cPwigtdjDy
L9PMcCxEhBr1RbsANIbP2gevOJ7fIzch86D1ZhhMysx/dUITDuu7hkHN8cZnIRMTVEW3LAPWFtU/
lmjjHbz5607pWSteXyJL0nO7IOYYhBSnCB54KkYKrNtfy0LEZ8AP/1wdBcwKmGyAL+W2ObZtRnEr
PzLwt/57V7xAe4nb05YNjv/ogEY0S4IDvCHi/4jdK1F9bGfM9fTkmaS69GOOtcay/WctSXBJufs0
fEqgkMft2T06lilL8yujR5jAiIejkMe53+KYLoV0XR0qh7QBDscHbWsUKJZDpHbtZZj8/dA/xr4W
+LOxNBdpkdHrgNh7NUod1wwjNLYk/YR75pkeNSxw7eeOT3cuHZ8oC0P4Dqc2knqwSSx4oRoRQKsu
g1ULi8DdiU7mxxwwRZJccrnr2P9qsgbHqNs82JV5p8mCZpiGEXkVAL0dzDm+t4X66qbsoDxidVSk
2Sb42/wg0xfJwIFRsAwt9KyjLi9uyXVAqXucWUGTKL/E5gguOrLjCg5tFE6hdO2QmLjiulv2Bcui
UkjuPFz9vCO8J2botvMcV9c8o3Vu5Vw+Lo0sDquNgzTDO3nfNMqUwrhyHulsQMFWWCDtA+21hZbR
KLKH9ki24jcQXye6POsMpnNwakT2amO8eer7N0X533kk0RbhZIEEhAvljDd9yQ+lacd59UnQCM4K
j+UoWioLDFNRbxGM+5O449OYKNQXpfMjTfF471vvPk/UpYn6S27R8HAV+jsYCueu0EX+b8NNhSOU
aXIZzjSTOPOgXOHg1Ks9VUMFECxODI6cOM1tHsmi5VFEBj2qBzHdFi7nhcZMNmbKD/7SMNkoRWsJ
X9A8RzbfBxIF7zd3kLScjhAuOpRWauoLBUR4m3hQl6jvrVw+p1T/10T8rfiBtoMStLrVzjSsj3z8
NwpUgCJN5V17b0qBD5oU2eCi8+8ytYKOiDKDc1udpxv2YZw4hb07UUbAHsFQkWbNICUiFGYonCq2
i0RsIMMKZ+k5v6ddnyBZDtUFJeOCmRrOf8AMrnPGZcUyg5X2+fHs3UkJJtfGuvAnI9ce1vj2cfTi
QqV4h+OYlxyNlnB5aeHU2UL9Whj2BpJmPisf33dtDBXiMZAbVgyH2KSY7ibFF9UfPPWElciAsMt7
onOsbKWOahGj3AGzzZppMHYoOoCG5WESZMvSWknZVjWyJsLiRsFJI7NFrAL4ykhmtp99w+2B+eye
gG7htnUPs/wsDkTj2xAiGUxAa+uC1QMZDn/GfW6VmHFi1WQ/ZW3d7N+Ouh2RppxyMbBQsiXp6+Ko
uw+quZ8mh4bcBSiv3B/mygZBFL7/vBrBVVl5WmCd+GGFsuDVBNHh7Jzew66/gxuvAZUKmD3DqyVc
hcGS+hjTtgHN6RsZftMf0v8oWmRBOE58sfKTBo3PXJV9kTldkMMZx77Gx1NOYmkq1JX/1ifPlOVE
ubhISPu7UPbrhsy/KYqAL2F6oXFbqRMBXCtM26NXExTL1n5AbeaZg5wgG+h5GpvMgUonJ7t90S1w
wOslomspd/mClrBvBdL/cLWO3L51Gv4xGdh1OwIxlmBVpMMkDduoZk5fo2rnXM7wKm1AK4PTrcH9
X/qoLuZnGC9E8ZXD/yL8RoYLjNx0WjcxMO7TFnmoRj9/b7PMng4w28cGVL/F/4BS5f3JJ+mxmAnW
ljZvro4RsgmFu3dzDMFo/mZrYcb1E8UCiUEmZos62EZ7CM2rbPcbkWx+j4aqud6C15IcmL6NKauU
kYpCKXxqzT0jDF+7BeUZCz/LaQzZCZ7LnJIPX+Y8+j4oKFDkWpDW0PXB54kBD0hGUJBG+uWGz9P+
w3n/xqxhuY5oPozFuobKgkq2aHfRaTXx/VCV5L+EJRy0nq8kVhbM6yPeqLhXb6XfQbn1ayw3BJ2h
+idS+E031YxBRrIitsl8TIyewXi5pX9qtI+XBAKysprAhSc9Xc7yP/HawZs7F8++uCQOHCed1fw7
8Fw1Sy4yov1WtTt9CnLB8jfJeVNp0vUWvnEDAgWQdeNJISqQ+JAGSvcisrNs6HYFrIB2mSp+QNqA
JzfBvWj3YXUtNL4zZEf9K7fFLPEC35G1BvUQF5aNu2cXCnWb3ePVgjIheF7P/UsoM/GcnnGDEl1v
m2IHOUule1+NhwRgLjU2CV+/ymDLnFhoAwcOTj8s91Jr5TEun9r+rTekY6Bmgqe6M4oyJybKVt0w
yG433TNalQJ1IrKpC+D943qcpKjPG/yhf0cVDAaOHBDkfJRjy+cV4x6SyHUEBYVmNJyTZ4Jt0ZRY
37/V9LD9G+xWD69FkQNa1LQ855PjiQ/kWRyLoEuQfCKZjH0YhE3JIfvPus3m0GlAV0CcyReI2fJ8
zl31JeKb04Xaj3UGZBP+QJIKKQ64iqediCIFYbiRzJe2FyV/o+w/0pKksjFR+HhYjAvK5UhpdTiT
tPBezvldWAl1Ou/LzkC02iSAlj0VnpON96AYXQmrK5XccJ7eRGCEpg+iCrApxNMgC0wCv5LHxOvq
CHwgKxQAFWyyPsHGQi7MOKDpOjyuKIqEEhjBKwXrtl3Z5H9SwQwTb3tYXh4C8klsSX1xRW1OnLtj
PIa5XAtTBKSx9eZ26k62bJodr1fnX1i70U+s8Gkrhg7RjiZNo7FqMSFdbqGr+sKOG0hMt6xC9jUa
Hc1qU9E5YkfjKvd9jFz1U4JNPojEEeU8RBtfpjYh/i4xnDQYT7QNzYmW0xlYVOXowGU+XQRwtC0X
+Ez3p30FF3oyMjXgMFEYvyJqHPJQNm9gYf4i/HdUO3hXUm1Si5Id143CfaJwjmGaFpH9sc6Ypy6Y
0PSwLfbXThdVrbX6enyWipTv7fyn+np1XawRYUDpYepRrTSpgj3HJvdgeaNmPUEKPRHWaka+U5dd
VN6KSdqaFDOeu128k/fxiRKD3E1ISIFQTWos+k7QGf11IhEO0IPkBSkNGLgEYqaM8xjO0mqjYJWI
y+Wo0bHc6hlRTvAzeUkUp8WKhgcAxXhSijahjssF9GUJW9ctTcfrMLdZGOuGgvWUftgi4FQX1I2R
DiLUiKG8OzLxeeIHsEKmcXEEWz1GpGnJwNSFwEa/v/bYS3C3Ug+WDIky+h+pIoxJYMjgZK+0xOB0
DF+cyi0GO38G0Eo8xFCqEUP4tYG4uGpwvIMTvX1IJBPz5rAg5yDAKFX6jHAVyvHHROTXS6nR+KzQ
20h5bB4TPNcrOddbSbJAdmHNlYXUK4n/LynI1vE1Cg4uCiGoeh3qSs/WFfuWR4csblBBVvC/uYCw
DuTbFswH9qbIaaSrwvgjN3TPcHiea6/GWJnvuxxB2EA46mpg4KYAynDtKjJremcAB9sVUNwVPtbB
9q2hSUXGIVqZOWAr/6ELiBe7Ma3NHBfMPSw1GIFozI7a7AXYWNOunKUVT+iC46XMaKUeEbS35k9F
N0YxVlc+kn18ddkXr1ccNM5pM/8nucL75rPalsGfYvTYlKh/RUD1YFN0wDGJeqmIaJSMzlLAq8wI
RYxiDZrvSAm2qf9gXlMGyQMdx2pdT6SQUFMmvrUsOz84XIBbqbZh3+vqUdEe+W/8eF3x6MUevp9f
urlIIjvr5dXUamqEE/hMoenyr+oUW1BCyVhrnroLCyrBfsVGnBsNBs37I5hiT+fq3OA2n1Ed+Khw
c6E0DBRsMkszk6CZYG1Pk1stWq19vxBVwYcG58IaTIF0gGPedn0q4bcG534HbLqogP8hfUIpNWUY
6AT3VGsCEoy2IAgIG8W2W1fdTNeYKP4r7Hi8FzXLArDBH6GQzfv/Rs/9+8BPAe40Qps1D7/KDPKi
C7yL9Ef7HJHGuRX/ONM+sfUoQJCpeg2GldoMRwQe3VpDUDtB1jz2J/DLfQVxe1aYAi0XVdCA4ugn
ptfE5C9oP+qKuMuhxvrY1mhORbyOIToV7jMtj9P0uEylVFFKCi0mNVDrYP0a+QpJOwXtn/kjxIpM
3DioJf+hZqDP7LpXEpisceL8XSjCmYFp4QbveNODgG2XqMHddsLSiMsUwaJhhLLZVu2EX6FnymJu
eK57Tifjz6YhH33QEYnxb3NXnr135sBdKNAoOaaECPuPSVtySE4qNaNv2OIVK70VOfGPK7hA/taS
TJ0T/aoevxfYj7MBYX8BDTWlx8g5dr1fmWZA3KYUVC3QvfsJaFSK8Ig8gfqaWyOhCezTOAIBwmi7
MpFRJV8S16FDLSTa2YKDjn4e7fCOJ1xo6juMEYsTFgvB8FmfE9Mia1l0SPCyji0YkuMr2mRuealr
yKQGIohjxSrOAx/ctMAMbTFWWaitxa+mSVBYQ3XFsHJrvwCCMAmE0EAw60FzZe21l96ky/hcJhX7
FtwXJT+ZRDJI9VcDhRoVlOeLoVH3kVjEUfJR+KPHjykuTx4BjRgoUAeMn64KrKMaFTlq6bEjuxRO
50cg8bBqWJakXBQceSlZ8B2GJfhSAVG3CGLGq01yZFxvum9i5sfHR9QU35L8mI/QhcW62sEexTzB
LUAe5Szi8WEQOiTT2nCzB3Sq6BSQQW/KuOvva+OTp/68Hr+4wJa+qs9h/Ja1HT+QaY4Fi/UMO5tj
skbXG1SF7QOyHBfn/0qV5+IFJrKBV84jIPy6H/HVoe81EQzwIxLYCCddMc0acqRQwOxvkmRUq6LS
wF/7bSWzySkPIywyY3WqS4oJJmgKekgypjYLX+rV8pVUydd4uNc+I/lAUOJZvS0/1ZUyBsvXkiiI
D7irxUrA6W05WYeXZQxyG854AQyJIXsuDPFjZ8BovnlO7ZPZwgfsLQ6YeP1ozBK0phWAJEnaLHmK
OuoSrSclfZ+gH8S2x0OCm7cH949W8ex4N/k9KelNxPh84KXsifLBcTH6622UH7H6ytWXWTV/4HvQ
5IFIZnSNB3EFyrjBcg410IAqHWgh3yBvFYb3ibHi9S3Gi5qRIHfvDrkjBKlbibJS/0o7ipNMaRqc
Bz9ripaHDFTNsrog1v0XlzJc1pGPjo7OHBGEVF7ejGMebInlGg4S8xGP8uDXlyN4nL0uvQcoJ4QZ
GmQ2V8CFqZpudbPaLeRpvR5f3VchGm1yXP/ljkjkscA/fCjjKQhrQ3Kz2lFG0nRY3GZ2RO4gxFne
POwf+lgYZib0dCHw64yVfbX5lc8SwP6+11g9aZQPqFkkBfVxjPRycL24dtrJrfMKPXALmeWNPNYZ
Xn6sg5LzbpFUufC5Tgeac0PtYQWIdZVr3lZdOLFUpWtR1aNatpTtOOsZxniW5LPHjZjUpj1B8cb0
uySHVlLrJylMQ+LtaenPhmcpBnZn+dPbzBzexPVbB3slMhs9bb5WhRRlD6ebZb/dMV2wEpCpJJwv
nc4AYfJowy9tVzZ9mvJxit2gww8p7nN3pRPVGqeo4gVvfHrSApu2mT5v24+QUX43wWnBbSATHxuf
4dtwe3yIOyLAnsCFO1Bxitge/GNqGEYjMdJy6jBQFFA505kMLaZHUbRfDRfsCT7wSpN1X/AbBnGy
UqHO+CtDcS8jCF9Ww7nrBFE8WthmImFUeozb9mbF3HO/sHgMDZesqAZMVxtAPCHpDL5gOfFtOYzm
nlCuW2Lk0LxMphcr0X2JxKSYSCOe79a0GFLRKKutQGRH0N8ywz9tyOU5DewOixJQFIFinh1tbZ8/
uthf7dRy9SUVAEOHopLG31LVBvqrWmZuRjTVz+e+65E9VvyLjjiyfJ+DWI/2m8i4Uxc12EjdSgt3
SUhJF5kHDOSorLTKg/jVdLkjWV1bQcdRFL7SJzUqup5rZlUdf+5EeXw/0rFntE3ie/Y77fdNio9S
Uhyfig2r5pcCS/DWjur+HeQSG5JP+NcUrKdEIUwvdYuSiVxxUHz7tn0jyXzB1XqWz9S/A6N5pQUN
Eb8SGareWHnhGvmmzXT0T2kR7MGr63QOFY3deGpH3v1Dn8xVMMWegMFNMaokm+FC4gUdl8ovNnEZ
DGyWosadWZJT1wCYIkz6R6YJwO4b7eDlGDp2La99wwFG9Wuk/10vQkn3qmd14mxBO/DKwc9J/JnP
XTrkV7nOZYcIHgiBqQwz7/C6XJKE/hYsBl64XI/gm80DRWJrgESm6xtC34apAve3WLJJEbqaVDl6
/61sil5juIR3qcJNzFsq5jMAnvJ3aFUiPwjfI8LF+O2KYByldKYTMwT2N3hy3sQ6dOyPqiW7Yp7j
aVxJGI+ab17KFG6OuuoXClp9RtP1DOJUqnJVtbC+ZB0cTP56AhlQBJv33HAxvn4cW/51IDD7/d1E
QDznl7n+T2JQoxPYeaYYbYX2rscbulfSGu8R7Hl1arnF2blRLdOEevu5PIEFwPO+NKt8xEKFxzqq
rVmqx/5+wHaDBMaauHL8SUX/Wh88LZFlUKEniEoVATFLM3VF8+WDfKbSeAjLBOcD3Hcsl9Tqw16/
zgQNO5YVvv5GjIs+FOoqsrU6AhByHiCZRAWwD2ystntJIz1tnXBoUletYwTjdFNlzWCgNKTXQY1Y
3p2KeY3lIfCtFgwOWmnNR35Ni/n2v3d1ItNEglY3qrkpt23C4aoCJCB/TnEzFTAtEn/Sc/defIHF
sylRaAwwjrgvyOmR9c0PYmntqeLwt6hArsChQ/s6Ia39jecLhKnq6S2V19VK5x+t4yprmcLWLC6T
5vVtEFi5cwv97t8j2dd0AFvKWyna3vK4bRK8q+rAH5PSyyaR80MK4l0Y4/ICSVbR4QdykvHjZkhu
Tw8yFZ3bXmIuUfaScDMHBDsT9dJedVlKh0d1sm+JDNlmODUy5ZaSLNbpb0cL9IKxatb7yDS9uQeX
wQl+f4ej9MZhGuOsw6OmuxBUYbRtrDPCIeN3+0hkUMj9eN5bNs9FC9llbg65ASX86v9zdTjHJ4Pr
L7Y/kAxatcMXOty2TIZ3QxKzpR8eL86eKGpSVqhKUamwig/JRPJtSyALPg41Xb7I6RgZYRPbECfR
u6oF2s3x9NY0OWRVF25btr3ejRUzMi4HgW7ZefHMTSfnT3DN11aYSmAaq8KzeWkJqLX4yz57pSeJ
xSwIStQgYENiAh8SLy3DTQLGC7/n0hQzNcVihNNJ6II+CWw5v8tP8U2Y8UKUzKbDydQbwWuMgX/u
hHHEbXNkEqazQ3JpM6EyjVqWb/Bw9yldImcQSCZHCpG/eEC2JKEI12WMdRSd2YhE7KYNYjAnBSc/
cGe5ASKpnx7TMpPJU/QcVO2GpkV6jryrI8jajUZeCgkgfpBBiuOsoPqKcYI/3qhUJxZpX2OFETVB
h0YZVKQCsMRCoA8mVmt6Y5KXQ8gP8g1kooU4iFD1o9g61q5N+F7d+UXHPm5JjGwXCD71jnroiNmA
WCtzcj8Svtveolx/pF7CzIwgAswAlFqGt26ig6ywI07uYYJcxXOz6B0NuG0qN+3PrWbxxcbU9q25
aL7B7zK2xHV8np5Vn63WwfMXOA15ZtJJ3HIrxNSdQEeP2wZfeaSpnLL5PVLRmDKySFnXHxyA7fY7
mJwsZ8VgXNzz54kK7GfU2npt5lIF2v/7uxG2AJmTRUelT0gJqbT55QFR67z1/ybf2rTd3R6McDqt
VzLSBHLdsjrlsPhp4bbPtbBLndZWByt4Ejdb4XyHVSNhezEddQdmpikWEN8WhaGlgUu5GtGgRAra
Lby6we7GrHpWApdbQQ37pN98Q+3G1LlUyJBrTzYJK69NPti73iAHpEsbFZ7lCva7nDUHEKx6LFUn
OMbrx2EOILlBpcCqj9y71d8WtPGkcncMT0KCjSuF/HFc7Yg1d3bxy63cy0pm4GMn5M3Qj2kgtFcP
kS1NXBQs2PMvw4MCHHdvQX2qQz9Ym098G3sPhzwqSirf80GVtaVuMMXrOMUM2CzDpgwjbWSZmaJV
eB5ukLan1FALuRT2MNpL/iErkqwnoIAZdC9hCT1AgH82tS2SBnHEWYUFaJB+Qe5XTlXCIzp6kcf5
YMa9cCD0ShVNIuMKEr+FcU/wmatQSTmlWTQRTEGaxIdorcVFOAD4MAa+YwU+CR3qANl9358FSJ3D
6t5MXvbpMHeSGAZO+SKu1Ku6GSWFMcHPk0c3Y81BbHPGaxMROphLysswXhxJ2no53WickZh/Whdm
BXZNWtrDkxR5/yPMZkPWa80VBVEiCDQ3zsaTjrPBWU0X28NqiwFBNKtwtx155zsbFI9aw9BmnYMg
5s2rrRrMy4ciGVu5rwTJ4b267jIR3UZS+v4lLD17CEWsloljkKFuNxUsQ5HbZjzHVB6YvSD/w88W
obyld7fq2aGercyzxi9CkuJEC5+PLmYRThkD/fXActKoYmmjBLj8mSEpnBkU3oZiSX7YwPWoWHGn
FHwqKx3c8iCDqS98wzfXrakmPS1xrIVQdsYothDoKRGJsNSV/teYjERoHhOe8JfeTS8lNLhdi5ZY
lZPjB82Sa19dDNjqpR62RmcUj4B8fs3qYPzvZAvsMkMnfdvx/HBVeOEPVpdmWI71+3QTO6Gl5LjK
h9QIAWSrNblu69Piv8Xs69nR18tw2UTRmeVpPt5j5/2tBLQWM5+/3drhBicnVxOi6A8vIJfbQdz3
ndMgtg6gkmaCH7MWCWZKaFxcxh2SGtg7c3gZie8T756AGplTUWPFs1qVeHc0d4E8nlfIgFJYd0/7
3NjjSzF0kyHx0kr0/jOoDrb61Y2Zq9mw0oueg9KE9RR2Gq8yINIxMMoeN7PwQE4JWX36e/dbgSsr
WvL+z4kv9xHind376Q/emJcDGKUAIorMEBwxIi+QDh5l3l10oQO/dEV8bF7q+y3YV18EXY6A//aR
0ZiAcUS1lMjHhE0ej2ORcTCQ2JItgKATTQxopqczIiA8dukIk0oKxcFI7w59XPrpr80qNdoN1TDn
syt1SbsyqqVtnEXiWX3idlQm7jM5/6id48ZLR17ZWVfRJEHUasg95OK7nt07N/sNkA4PAnXSpUca
qj8BRh4TBvzYd0i39QbVO4/PornP/QS1S1/f8hGv3qTadbD85zLC6S6i0qj7UirhpXtBYuqTjjrr
NPUgah1U77qYiZeSGEFZ9jlEyI51IVwB8tDUKkXdEg9Psjllzm9vNfmI4muFhWKLJTVu0t1ugTZt
rmGDpp+4wL5aLytFsPcQunTwdo+auaMFoCMxdsNclCVFlZpvgth8A6NWy2KRYJ5s3usszBLoso7v
s/YgrjsDdryb6O1RUZGbiJ+vRJCFO/4ZktNMVM3dOfs8kgrvuCuM+w1QyOV6ZX/LZLL0920V6hFu
OT65Xq0Z1FW0Glc5ULz75FvE0xdZeMQ4S5rSJX+vzJPEr8Jymh+vQTcHFb9ZfTC0r4OhtzD3pces
WzJvUAnhDoxT4WPunG0It+lPYB7jFW66zSFGdaoSIQJXcRlL5GwrDXmAKCS6/Tz53k2Gb/M1u3vG
szsqfiI/yU5TZuXqGqx+lm90mL4RZe1ZEKAr7Zi8EF0TjQMcJI5TRLmAPbj28QHxFVvkm09CIGZ7
Eri0AfDpS+LejiNFWXbp1VjjAzydJdLg8ce4n6cqF2sdMS2Lr1dd2LhaUcgslD/6mtUh4JnBK/8v
k6d+jmzF8fcbsRGij1sjfKSQYT+QGrpjg1ZEKe8j5o1TrxtpSZ6DtWR5NBiZYG+wpNeF45xdgru/
sny7+2mmiAG+OAyTg/nR+O0UqTrpKhPMMBtm3qyZIJL2nbJnC3MGutW2lxd9FgmxaFIbK2sAvNzF
kLsZMZdvQVyO4kj6CBuEqMK/XvjpweDBfrNmUsbWCSFcSMR10tK5wwZfYqcG95IQ2b70tfRWpCqd
2QMxOPRWd0rMWRCoxf6HKBjLX9cb+j1w3UDmdkp77MSyXdt26dVoKP9vLn/+vnoz253QBngs1Yh5
tRn7sFK3KRKfyZZyTqo5ZerDNgH1bKmdYZQB5qdyP+C9Rc0cIBGnjURibMJlZCnDRhX0s/U6OaWK
qhWgn/BzJjOXPyLMR4J4qDohSyXKH5Pp3J0rnvIkzmgvc9KDvjUlxAdNIw7dIgUqWK4QdSoy2fkF
STHKt2nMvIATZQ0SmJpeOWCn1L9w56k9SI1gfo68Xhq9I8nflaiKRupAnVahInCj4IZFyA/kq8u/
Tdo/TmlYWHk+sRIWKgS760YF7hsDg+PCLpI7BGUQ4XdAevKlmdnPmhcbSGikc0H0MIkTZIWJ3V1W
NNg3MzsggZG04CPCLjDFbrb23BSPK36OohIBc72i3dNz5c4ja9qsxRTtCn/ZxI5tiQ5oHuyZtZX+
xtwVAWDKvKen+A6LaX4NHmghbWsxVr9S3BNI9HKJW6muC2CCsSrbR6d19N6+0YuBQmOSa4bK8hNz
PSGgr4131UqLrFjb+2WTVbkQCrE1W07c1fMR/VEE9xb/lDtz7DQhfEvwNsBQbeuQREDsTwhpMaJZ
zCEfxUP+SnMXxEYjZu5Dllx9iXtgwXQpjaXFbRAREfMyeYrmlSyqb4zwkVUUY0e0qgHKeAnMJy/f
5IarNl+Nq8ygkv7jcioFzgGZ/wNy+11H2rYu6G7GfFs2CiTv9jzmEW41RztdvEBJRBJsu55t1udo
rWdwxO7cAfLIoySy4YhQoNK3zhZWYb0NPOKWkeBZZsQhgtcDCFJaIE7RblOV2w5jp6CekbWtTZ2B
xctq0mE1NsODIXdG+dO34WLUoXpwgVfl2A013c4Jh9Z0hhkUW19HxCpbwSm3yDixQmT+MvHme1q6
RD8qZppfM1cQ6UaP0/GvDdOO145PAJwecRZIEMn47JzitHy1puqn5v2sqlLeIZIJJ+tXCGbzVmxS
RFRxTklkMxmG/sIGFDM63gTrk4SQRyzfVyiiEiP7IecS7/RUUEAmQg5A3aVT/pAhmPRNIy+DkD9/
6e05alnxPGPdywz/mncJPZhmLHdd85anryVfTOLd9M+I1NyXIyXnV6FqLJXCk/Cl8mH4hvssl6IJ
bnzGy/PhBMxsUpbw7RND4GGn4TRGd8+54dHKvn8O2zwiH6GgSRgQfKLrD1PJNLU54CuXOJrfAPrG
VewtLuoNFyjaUBatK/5PIrFHD2g40WZOQksEelux72s90eztwnk2deHkVqdQ6yfAJFiSGX2AEhhl
bVMIwGe0H+ICbtea8nkTHlhf6GuMOtQxPxszgWOrWXYONeUsZ7TrYAZDeViGWOfBwrO76WZtryLt
OVIs3oBnFpKuK2pz0rYT2KLUxo3ctIwmcQNR9ULu8rTIq+iPqakOUVfr4Erbr7Sj6Ji9HnqlcxNV
+B27JrgKPjevpxo01r4TiUgqWJAZzGnRy7CNUO6MWwKuJKvjuvDaeoUUAwyIaV5cwic1L9IMtdQ9
DmeI7sWDljvoDbDAzA/dS8mb+fqXRzD4ORJ62D6VNvVWJXqvE4pHl182MdJuE8JbAger4klKbEiw
HOKhQ/I32Xk/SKqB77MxyRvNr3KQqOi+AKi8JLPBEnQRCyUehLA5GSZ+s/tfdua0+CmEfzgynZR9
p31xPrzwc5SNBWJfE5sfFwb+kaj0Sa+5LER9RHyJJWItIm2Nsj15jyVTPlfji6d6xi20Q5cxZg2M
CSehRWQm/+n6x4CwPp0je60HlXiwOOIqL9IVRfzPkveokefOWXCWnyL50cAV7YSK7Lzl8BDAHgaF
MIB8bItxibiACEwKlo25QD6Oo4Y3fOiAi/7lztxLnKcQ2lvvL+yuDq4T9e9++VpyhyXikPADQN0A
agxBmUdRcEp3kbHeXg1235pE7QHRUPcd9Pwr53lP5otWKCByc8h9soCQstPeNUjoFdNP948T/d+2
E3YWlA4Mh90zdGIrZ66vD6kYCaTFn+85M32cvwtO5eEsPVXLoBAKCNzEvRXeXRKBPmt8AYuJz0yT
Xvr2EtRCvZmV88lQ0aEi4hARyHlMWACSJQk5jr1PSVbzylYwj8mFtZrAvDWoTkrmv7F8pABT9SX9
7UFES5WoZg6CnYQB9JgtMST2xgieBt75PFyAO0zpp3lv4KWG3hM1jBD/pzqEm7+wdv6arUGKasHB
u3vOkZ6OpiG7a4XnBcKigr1VNj2tpR5nhAdVH0NbtoJs3QIGWTvhUH7D00pJYT+79CTAYSDQ9pRg
gr0YzCz0hMLdyu+0oRZ3H/9Gcm4fn8dvXnqG6QBifHucXAQA4NSOxLbhAHvxDIOSThfyGdZ0FvmU
wdIQWBuEWwRMxM5vM2EYYuqwxrawQj4TwOv57OrnyOXlSSLZGG5UvgWOFxb6TNLGSd1TzzNjD1lA
FsEvBZCh9jCBSQyAekrlAuJY7AAn/4MikZQqcfgn4FRtcKIfSSFbK0DBG2q4LJOij+0YujJtnAw1
yzfPg3k2z7bE/rFxLll8nvLAgFRdy1f1Vv247PmUP0Uxd2+T6wmBVnUv4gVlBdCHWCx2BcGKJqvM
SomVwE4Ow8uf6K4dM50UpFolhLw5W/eUu1h3yWDB7cD691Jx4mWxT9hiz0y8Z67ZdA5jSuDjI0id
HvgTbO02WzZHos/021oELzdelhN3k3u1QVc6WakOQAQg5GfYMCHMPNaCtr6Pk8+mWVTD3puZGKnC
gDU+8LSOIqA0mPq1tB/sobFXlFxZrcsk3p0KZZMgls5AHQv98BqVN+SaxNI1oH/MyvAll0MQQGKb
JsRNEbujnaOEXHGSpFrZmtYSWMiOJabiLTE4x2y+7XOfs1qUnUvlS6T5ljgK/901zXdSPCb/o/Yc
mDITnp2UHoHr/W9WBYUyDFL4AFIy+GLlqd6z1sFdkXPdjojCwHPL1EreRsJAos8Un3FtqfjIWUhM
7ixw6pVyhXzynx4fGfLggNMSmbhwKQ838oEUf27OcAskWQlp4zg9shcgp/q/EU4KlyRSmaNHz2/J
tpAbcWPdJTYZnzkBS1TnMH5nD0hkUDh+Qg04g0UyIqnRqVuPpiLCbL1Atnppv22s3hT1bq12TPi1
fO3Fpf8/j8vMkdm1COMiAat2Kk+uidJd+wMn6FwdYzthIlqITa2KwPcuHhfGBDMmGzSTvRoGGokN
F8ldHYNR7l2vu8DmdLLfjDy5i79Yha94tEUrtha3I9ou0TAXCMBPno5hseoCaiPbE+VFwneoIkDX
nsgE80utAGOmBqr/T2d/VHSyHj8azJ7yWbwXPr9A5YlNfK+GybJ0yr8tM3zQ39W7p+2xe5tgkcIY
IJZxv0iuNoDe5Gfb6ae8VxpljqL5CGOBtcP4tejfcCv72D58+ApdSNFwdfttcNX77g4vTTbKgSvq
LPnnUOX3dvShRRAPoa2EcfnYkP2iDZAy1qxpxZI3f4tWJuTYu270fvh/EBPi6Osor+H85N/zPGYG
IoWOaxyLWyWB2IgWa5aG1ucvaepTfCAb8kAHXSKvBi+nSbDPefhUxk9deEpxhoBuJ/WcV2AnYtJ8
nEaG6oEyet0Xzx3tQ0P0lKJnc9N2HrVqo96e5rsplwiIajgdYe3+vIGMIKLMmYB4u/9+7I+aUPbp
STjHZH5PKFJrXmBE7zM8t3VodJSWpYBZmGGUJnQF08gvieE4QTgOg+jNPA8f31/vsvGkm8aBI3/H
++hBiumYxIrg3wvoZhpeVssABlNNJVCkNEw5usrCSkZsgln3ONa8uuulJi5zQg60S5pPy91sjG0J
hJc9ZfPwkt1Bu/KrKnyAtRbeINlQIfDARNeLzGJULdt5jUu2XoNG+jD5zyHlNY2jwQX8+oh9x3Gv
ibTmePZhq2HB500LyXCvUFqqJjsXNOYoMLrjSyut7CcHZnlb5ACgXW/njHNcXGNvFbIxy8PrdYos
/CTBo2vVQHtsQ1JVlo7W5YN65wdnfWG2SOhBtH3RpZesXeBc0Kb3MXQIN79pEbiPDWLAY2SwUwEx
xEFn6/QsY1+NRNIZzYsJTfNAXjJ5fLkwQkvlO0LxXItG3Ik5ytZYceZXl7YATQX4PYcnAfx6kAb3
eEgst+SScJmuNUjqQEhp5u7192ylPIRTlFLateEgbCvBbseEmgTPmYPbQP9e7Iz0u/NCSlXx81BI
c3pXH21coQoeYd5HFoAYv+sDlcz2UZyCKlXg8hcXr7TU0beFetCbvt/2X9dFxqLuMMF7fzae/1gH
dEBC3ZWsUsOfjd0U08BNSRA2EIjGxaEJ1S7jy6HJTfOyEIaGneNx3+6nkz+7nNPtE2PU4Yr1KmXn
0x6s0OYp68mF0TLHaKgzn5+89fBCxqTs+4u7pOYM41VLqSQKWDgHlVxtXYQu2hssu7cMw1nKS/ML
Snb+C+u239+Eyc69DIMjc7H10hltmS6RBEGOKwNq3hZmtKrLB1LTOAhtn59L++ciSrGDquyH2Q5F
4R8b9VsnGi3PWzMDhUXNZumsCrOBeMEQfIBVenNr2oHf/9lTEI5GKO1tuz6/jP/tVu4gjwDNoT0w
jDL93G6jkhzjc/ykkrk/SyTYOVoh62Xw3Mxtse+AEeALq+dKy79QRK+OvYhSvgH0nYgp3blmOvnn
bzuIOxqy9ZUxaug7UK+JBm23PkhzEIIp4e9/KU90mugATECAactsNExrGV9aFgCzucqvGLsfkGtm
g7crCXSkp0BfJEcbqiYCdoMEtASDgcrEB1rO6NJP6XVDGyyEVEconuP/s0Es/gxhKUXFfXujf5rv
XlMMg65dR/6ulpsVSRtk+Wy05pxlgcc9n7eILQ3hVYyIHL3gdyHHlp1AL1TY2Q1ffO3w/x4E4J8F
0tPaWUDsrHKuGjE+HxyColHHfr60uFhEnVQ5cSuHPn78yTS6j53NSCggAKkdRLWM2M4yekygP82X
RlZUKZRyPQw25dkVweY7HTZHDJzo5/6HYcS5L6mWoh1lG498vU/jtRX+lOp2l8Bf/8jRF00EB9X4
9yjVWS8hhBe437uJbpkhZ3rygypSFf+rSnDICUsj2UbkBORd9DUQ31mRoRwN88HAdtIfQw1jeB+x
+JvSrbRpvvCcwUZOCj/jNat0YppULPswWoqyTMitNuF8cPPb9SA/Kgtkrj5q+LMY6l8V2Mw3Gj/4
RUYg7O46GZTgEDFEg5de2eFL9M/zPTAOJiLvP13RBYGh/KXqPlXoQngRL5EKNK1vWiGW0SDvNPJB
LNBKOjxlGSEs5/wZyYNXO5OKtYHa+FUTo5YIFN87zN+6JUiJf3jhkS4iDJeRX3D2M8Af4vpXHLTC
Vx0XRO79PbbUXP49XiK92JOcFn89rkFD/9a3tmTau/Uw3gagl4Twy5rNg1pBvDrz0arLM0fNGDPX
1TcJxFquODi/41qWxbW4atqSuMBEQd1gJRrKJ4RrS56Im0uL7peAeztlRrLnup3LjfotDxc3JYaA
w5dUU2fPrp22zVaapAZQwJPmn/5ETukWJ24KqGjlcUHMn6AcS1/D17jcf/Wa4SPzjuZZONr/LJj2
ACw6IMUarXdCrsUYDF/8ghzEGSoL7gXk+9srUVAWc4Xj0o8+0ELlyYmiFV3BqE5rkc9rp0fCJeY/
8093d+c3BLI9iEQtDIuVJE/9lvR924TU3OVyatnDXSCofj5dgWgqphJE9ImxIsZFbnTyL97JRxAc
jqrZxFPA7+eEMIRqe6X55hd/sCr9lL/OzcCjdZPJuz8DnMIGFb20uwhOWR8EzoVpnhaHZwmgwa7V
esnKToJUq17PLGc7ozCz96v18+fsoAvxqIw+EvBONjD0QoLmxP8fY3sGk4a1s3+HkzPMRQKW6cl6
KirFvsBRS2qB5PE5tfV4Roa9f6AwYIehM0eQGFmWeCSVo5aFZYXQHvzO5hy31hs+arsTQaUwN4J8
+dV+ngx4y8MzBao03jC7CQwR3Qxe3BhngKIFYFTtzlH1GtaDl90kalwQFcu+YOOxCa7smAendd6y
mNBUB4Et4MqCBGmzS23soY6HHUzo9CbZJNh9KOpJm2663KVBYIEqr2izVzjFMFmKvsbDZzh8ipE+
hwJif4ukQ5vpauEMIPnVz/AeakrACqO6NyVyeGKEm+f1yH7SlU9qHW4Dg12D9v9nWEs/ES+wVhOC
MoBuyOF0s0BqVuXvnL5hp/Lvf7xKcECfKsUY0iS/Je8tRPX1+T9TAB2LszL0t50c4ysjwJHgVnap
qUHA7sqRallivNtonuxwSh4Df9ecnpZCrh49Ij8cv7or5SV9v7SgfYp77tLyE+jSb5TSKTpZIesc
chnVLtOHMpZ261NoLl8hUlg/xABAh9TsIa1FwiZUyFJneOhtt6G4X60LaSYkVOFi6lovFnzYA0oj
JyPCZxKmYiHaNMjUdLtkHHhYWkxnnpxQ2CAW/pOVGXG7mdr/H6BkCzA1359IdT/NUrJppzf8g/PT
h9PGdnZtkMa+MbML/WSu5Aybq7hJgtTx/DwadDKqqj3msHb92EgoeJEj4ZW5ceFB4dzN3JCEPhsD
kVht/MfNJLTUIxOmYh9mxO2od3+EBakOCrmMErzszh8WNs1xI25ItOGnwc5AbKb38XKGFMzz1Eug
eHsDPTH3k8t0EuCwm87B7zc/8iD/UH1N8b153A4JOlfQFv7slkUhyufKZyJ/Ai7AO7Bz/ZwNnJ12
lWT9LYBs6Ph26HRh27OOEG6bplM/nIjcLUSlILPPQweUH6M8EGXpULlPhNN27u+c5i2MYWoPmX1G
3xxBcF2N2bGyfZtUV/vzjh2V/E4wi6noXoDPxGf9pe1AvRntenKJeFNrTVFCot/xWf3/PElr1oqd
neQuTeChEwAijdClbn3vP7KLw11uJNFc4/sMB/EEi43bUWxPlNPRexgSpmykXXSX/Ay2dIuZg0Rf
g67pQu1ZDBRjrobLqyNLz3RS3fHN/+WXXn24kz+hTMbGrKCk6kLGePg2ZYv+SNcWOGRLYPj3DfPm
e36BvbdqhTc6LqHVa6JeNI8tKbbC80k1TZOTkytfpVa7GCsW28QweX3eIRAykEkLfHGpXlGl0Q+a
lurpMLPqzh0kfX9R5dcYjwOIWtSlwwVpDzR3f5c7eTcuJnu39fLzzTcVtaVo0Xm9UxCbhatVTPX5
5YJKIMBaeURHQIJ4hf+36iB4gta1lQk6bgoySjEGqPqof+oJqueMJWpcIUVd+oEQmFeQecDFIvHL
5ZhVfJqqwSbzessqSia4lNMF4J70tOz2Qj6wyujy24cIxeEKWSAQNqBFuT9fAlcsT9cGrE5plL1M
k6pwo5DLdr9JBT3waJmQMWv2ComFOwhbqfqUSnkt7f9UKgG/RxXy8zW2I4soKCfoT3tmR2dpzSim
lwLsnWhpFq8U+RCVtFtzMwT9nxuO7DEMp9ZxOkEC/8Sk39AfzrvoCbCtwdUSvxcrCMFm016sppd5
qv0+Q/nti0GjXI1c+3CMMy/I4oeCXqO6tsnChCizIBKEJq8UIUiwDHNPvVmjmcswvnTCHWYruFm1
rVimbm/h0F/mObQ//k8LaTwvwOFOve8E9cyB6F2bVL2v3fHdlJLg7jj1UHCR+lDZNVdQMC+uWhBK
5FV2GggGHhslurUtfJSqSn7i2F8OQzaxVzij3iMb7C/e72nCkMkkBi2NkLmtwxbm/kovrpIV0kSG
TnrO26CryGJa2qLFe7dC/u2PgC3WOC+8Pkt4O+fpyIgm380gpL1kPn4dQReRYFLFrCjlVvWGzksX
VjrPaC/tNd+YT8twwvwwv1gmQzNSjUINksgaU+dsFK53txl7jlzFn7q724hjylvtfxqHK3ubQwha
HLVrtjOu9ctaij/Yjb18Oo+v0ha/t7WJymdx6OrHUOddOwoTQbsnostSDVY9/9BWhlOwQHvSzOem
bkmOUH3nM+j7gv0AakCqhaHv/5zCbx9PCO/mpxgt1wyEMV25+ksrayoX6Xm8UZ/UvSwYpqGuNJ/R
NgEO6mWtZia95pNkQhchSIA1wEA97gHESpXVKLcJZAY919M/3HfNH12JCbElJjGmn9bQkCsP8OjR
hpgTDUZ8GjGvfNLQfOrUTf/i4oA5qyD4aGdt1bibiQy1YdiVnBY/9ee6JQLBtlyEVRF1xOkG36W3
UBDFevb2gtesRhj1z13FWSwotX/e0rnFYjjdOw+DkMlU53TUsvJHZyCuxjQSvSAFReHqFX5L7APe
qIGmzhxlu//6+n51hkMmrK0GM7dq1hZeLBhCYbrGrM4ukFFwCFE7jBy5ylUn5xNKTFt+ZxyBnXb7
PmB5FdmMLtAEWAKnJ7bcK2PIUL2vuLwqf4hHOqzvdy5e24gz+LAFFYGyVWH7zbW3fs7FROXPf4Bt
6Z+9R7ImgulphvvVZUnJoTUzSERsSbzejjjDeUj60u/I7CHLbySn4d/yIGXEdBUXJ3p8mKQ6KrNs
8deUFhbql+gg66SHpijrlHHxM4KbGUz18N7GdBCztaOzY8HLXf0nc23qYWCioMRLxgRpJYw01l1D
m2qW2pak97u0j78o3Vvgl2RvBy5+3pODOeSHnFO/wZZQ5ZJJlknrvV8ElvTqBcmavSRYbDMn3rDP
wcHfxcfnCDv5rTuEpPUO5tcfECeK/PaG4wKMQH2s7jMjmn0r2JCHr/4Vl9pa6wwooUQ9vIcGq0PU
R9X5FcxrmEoZasBlgYXCaKVtx0AW04N0+w2Fajx6GuEYcfmsmxJ4zFfLmYUa7clnikNoseIjgHgh
hbnB5DST0YewH4CyhVGHc5MDPyVlwwGyL1MwfyM/Oqj459dpI827hf0AjYuwCe5KcxzVcnkuGj8X
Xms60oxMfWEj99g0mzOIdU9P1uTh5INRGJJy3KGel2ir8JBWGrYgVsewObEfFlK73u9/CXVMrTN9
8qcOuU8iorIgJVkzraeUrpP9WU2IS7lXyimYK+TBmdQcvDIRrOlcZ/bjA9W/1waoIjEfLRVdG5k+
RXo0XNEv6dPIBdz8Q/eOLlYzz/UtIPv1ixbAUF9Y00dCbMZvoDaC+Vqce9+2SOsqHj1Dg2hI0i5m
bPQDuYan4JtXQu5ucO28TslM4pyyUOyEdqXGaQDDFHlq4n1lYH9Fe4wmkw5Z9xmOTAQ1TlpbfCEb
/8DX+abuFKOWjciqdHLxd6qfFJCvAzoaIDpb8lFCT5AsVWWPxKoE6jFERUxyzo86cG6AvMiHq49l
lgCcowoR0OfMlrIjUhS5IBknilO6d4tFI7HpcGS43/6REi95uEoJf1uYeb2sQit0bxMaUC2ff7OU
K9OmTtP+zPucPm3yfw4q60XSIZycJQtSmoo3Ntl1ngY5HPa4C12YZStpTzaJ59IHnIvnxG9Ymf+C
kO+2IbLafM7SCnY73AnwvOcTRNP8CBVKzcgJqwfwY2ywQ84mTN0eF/0DZeItUtuQg+eR5BF3rb5j
rLtO0XGg93Om2hY20M0TGpY629hexJS7fKpgUEHbNj/zkt4GhjOxVHmTimkG6/xA3pSmMHrYX7bT
xeUQ9CJic0psZeMDjuXQvwZ95bPharAhorujrZe4MqxeW5KG4YSsFaWAbDoJD2N/5nGcyWpiiSoO
KzUY9GlFR3N5P86EiZsOz+Nqp58j0cDq5rVV4dSiH6IRAJU6IsLUP2WrKy++xEhc510zs14cviQ+
L59NyxEeqLpA2G7vPPgPr6zMx+piKVeurjeU6p7BBdqM/417q6u1dzJu5F2SIbzj++552eA4Lbb4
QvMHGceQVGnM3VoD0VXfwyJJrNvVycf48z/ggSgPUtJvuyQ5qHBLRUroVhPK6UkC9hdvTvuNNh7J
RSbXK0izhnKaIDmnNFoJKaUuigsyHUUgBc3iI02PZx6NEAT6pW41G4p+tjgyE6JZLQT2zbWxnExh
glXFxEUP9hWLS3cawYxjIDdiYJnSRHzdSPxSCgF0fxorcHS9gfq/oIi7WASVCv+KegJIPKTdd537
RRSWrfNe93ncmyenLwYw7B8Xx/jkzVYa8/PMyKuWS/eumeuI5oZL9gZFZQa2I/RC3S9JjEazS0tY
/8psJiLN5hYFkIZ+MgVxCKuKZUCuJ/NzGsrblKbWNWjDSiBoKScr7cDaNAL6wjGtEXIkdZ7mTCSZ
OeIJFOu6GKYo4Sq6gkLQEsX1ysKoDHnjnAvEI4e0nURdQqlm7O9CRAoTReJM4Jxpo/Vp5XuqX7l1
WmTuEow/R/+6AmOUWq3Rwl/L5VGJG0a9HO//+HSynJLJPUhmCepo5SKeyJOW5go5MQ4JfMEr4s+Y
AcMnJV1Gm7WxIjsLH9r0A3l0zBcze+P+Q890FAXSrrR5FnkWIiKNFcE0PaHKNPIBCBVwpNbsEavJ
m9N9jE1SN2F2QVA6QJYLCwdLjShGzMN/4aqBk388DZ6tYBQn5Dh3Tcz6mjT2nm9LMW51Qcg+TG1h
OvFzgmMmzxTj3m+JLNGqxefPc0blWjTFTiZHphxMYrh0ECjatfWaBOnwI9VECdqtXxUCMeGJiTua
pAoebEYInoszuHtU8NyKEOewlhdWRv02EClu+LyAVgJz4GSujddRVulwCPv2u5TbSpxTX8H/2B1p
YmqhQaCg/wjzQo5GWbbC1TxWMdIne7YlTYH3LObS/BQaOoloIkiLE731RCeAximWY919eJFC1CJ0
L0wr42LZCbyRN1q6mKJcQ6d+GgtXo88sqtJpyPeXvprIyOL/fRKGyBQvpQzUmTb3LVycURIXn7KQ
2TmHT7IJL8CWDSuw7H0Ea2xigqwd6krdM5N0DlkTb4dvr58V6gsikjRyFzNDME4pbwuXaPyOK5mz
2Nx2L8kXfXxlAi1e+ilsJNzIEzarer6TxVXP7E9HiWwTD/0871UAfSSuEfpwO1MAV4JF4frWFw2W
F+xPHRmTw3zZrq5AocY230/7PIVkFG7zUpMYBdkrElrdQGtnmWpuZKNuA7LeiB0nBCqRBkDtou6e
BIm++pjnQz2Nyk9d4fDBbL+WKIdZX7sMISUjzy+5J+HcZ74YH8U9BlCjB9Iq9IRnF2+n87UWUx0H
A7U4COd3N2tubM0aCI/k/AvLoBO2kmfpdKYyxEl2CyRwmrhQm6137MGd/1j5oxbjHKkjBmw2/UJh
yNeJzlDbct7x3L1pjvWDM2MSvO5QyiOGp1fYXkz3PRy5baITdGdGCpUBJvvyVkV3e463zXYEHtsX
FfOgQ60c7AO72vixkhdK1OBwgTAa16OW43xGjc/eSr8oaqCh9wf2zVSj3zyKy8DVYgr/zLBH06wr
8sfv5GxfT4O5TEX5u8s/UGBMUwUHlw4otGDjZk1uiwpcJvaB9Y8ipi2miMYwAcZU0KuKD10Klcqb
RVnox3NR/Hvm6OkdnP3HdUBeti4/WtMbbGcgQqxzQV14NztPXCWWlWwknmR+FEqDVbO9Q7rJH/KQ
FG5+JoOL3hKC2AxqPC7+bukpxEip2rvVSPgoh+P69acFJxO8wJgArpX4KFVi3PHDvRwvKsNVvKaR
tI+IMdX5Oba00QpqaQEPv3Os/Tsmdfr+gCDaJ/10VqAH0dY0jXjVhW4oqUW+Vgr5MhXvpNZDUned
tQfvIRr4L/9ppwY1qL6iH5W/KLLpMBMXT2lvyuGo+q9cE5KmKamHTRbvrHgrZ4NP0pv4SKBEbDAG
Bznsk45+/swymJ9Wny9o1rcu/O6dRRZ9V3rkGEQn6/Eu9hbzHB6Q1/wM9RqOuKGmXZx4hqR0E+bY
Lh1IidN8db/rF2h4K7DEypBKsZ5v+0E9iF/B/KV/izGBObRTGfeF0Aa+T2q80Pwnksg0kLMZyxuh
s+F167fPZgSGtjYcogfGDf+sDJiL/39HMo2IXzZ8djGU2j1gP+VhUONMAQf6sZUCRyaYMpmyV0pr
oDHPnME3mSCVgE2wKgpoMVMDuCZMaGyobwGMYKVe5g4ziPLE8iuzhCMNULwS4UXh0kRyziaVONhi
9s22ErElW88xaHp3ELnU3TIzOe4mPa/Hh3HaS72/IXMAmGsxR3ZhVO68ZCm6wGN8BrLc+XP/gQFE
F2J0ulFrnHicxlExRr3gTU+YnbDFmDggRUZCgVoH5MnmKotvuo4ahbRjaCp5XuwcsHa9k/wDKE8I
WRqbFrBWOe1QqDglM9w+J3ynYfOKdUEQMZ7P3N8X9ImcWxyCnOO11Vxc0/gVahLZ02ru6uFDYC0o
+hcVbSEja9MloSH1Nvb2hhV2WHrtWwxwj/PUsVHgQDuSgemGYds3GWGR8e0fyYi9Rr6tB9WH3AWf
5/RiVRSvRcuVbCXZVM+FOQbldf+CTEgud/SJdg4YlA/PmWDT/TuIYRQ1bbARy9Br5424ena/POTZ
AioBN2Pimu2Wyn1RbA0lexqBL6Ph8yU57o4gwgIDkG69Tty+NuBUvv8fYOTWmDTJDPF2PbbPtLDw
uHMsyeGewczxoklJ6kU6OeKUvTUb0zLQIdULBnj+DdK5+DHfhxfn8awiHeRSqs+otPn61Xf5BW3C
tMO4S1nCrNTuij19YneALQ11gn9lEiCKFsdlayCVdIqazukfWtHiFZiPPotnCPxL+bMB5Nv5mDHD
9uhXMCVMA2adKi6iLZGACQQ8ej17oszjzfap0Z2cQ/X8Px0Cj4VCo1dRGwCjtedYIp8VTdBKsuI0
F6s8jblagZRy4qYcYW46OeuavRYONZ27JWWh9u02XYxHDB8fz0hDepStby7qShTyBX9tHyzGtD+w
kYzXhE8eklLbSWinmh+kNUJYu2R/FRs9Tb+3zf5Tchl4pKoNFOsZN+e+ECWQTX7eDiaTs1TWjWxt
76a9J47mYl3DMtlDy0Lc+B5NA07jNZCACqXCdbDEh0AqaBuIGkKHV4+NOZHKzYT6fhHgKZTX245l
80f06OTEmqJLilOCTbSHhCIXMa24t5fGgUUQDUFom90p7vjL3F0m8XP6wHvYaMvB0Kpzgl2nHqa3
+6pS7sK5SSEf94OZvXkwHxcGzwu0AB11z7MlJs3igz0zx3fFMznjS2j8yXCkFv8AcDnR/+giqFdP
0wdDCK8HlTSRXO3o1IrbDUDxmAFqvVmbiTfNx8sZO7tH6OtqW3k8C3u+hgc3v22S67av7iQeHuxS
Z1S4BVauy3WrIeLrs7jJ6cxP2V3IOMBv0VwPMlTl1whPjx1SvJNMxNEzyBTJYC2BZqFwcgjt9/Ro
khZv3iLdyn1GxGnXssa5uGIVBMYeSMRdXhChCEfk5SVFCnVkZFna82jatCqCW+KilwZ27T244AOy
6mvkLHFgQc0cG4OrZRErNd0wc1/C7WWRTjAqm7i/F9MnxmZTkpZo93NhwpunhRaB50+42Tn9KmjG
0qFgWPJ9xjv54SNXWzdD482GeEyMc5NU3smYl6UmYs11G336tsLGIMTHoIHTbJlvrefuuskXtWB2
qt+X/NK1DAYthESpIDI08mlAaV9kxLGBYoK6yJopHDusawZO6Nj6Yo5vSmSoCFWWnV3ybSClQ9qy
QNMrherMLsDu9vm1/KpFzpz6M8HesgsHOAwXeWQV2HR6jS9SyqW2PHa6TumOJudGqc4rxxxHuyyS
8nJ8boJkwGExENuH/zmEUX4HHtoXywykKbU22skg5pisKpXft2nHvxUXrrbcJQ5WLlLHRqe0HVvS
z6vpHTnW7FD+qJCcF0QJFq+qr9OzVfmZ58SRZCpXa9UgMD0EhTvciMr8x31lGxPiVMsaNqTy3IQ2
ucDpr48NX6CzfiJm4L7o27HYCg4sqnCH05gztkhsEX6gfeBe9Zknw3tXuMbu5zQwg/rPMPXjvaey
i0/bgZBEPkYCPmU1AbM3S0HvigYs+AzRToua9FS7d+2PPbhXKo41/NuS+kU5wHW2faf/LSO8ZW4O
orJHJAfASlvVPRaJ5Y/pB+GSqiDQZSz6HC4BFfnH0rXxondRymY/K1OOSvbwF/CaIH5VS9ZPzASM
CR2IyTd/hgctLtHEUcZS4xSNd9pEJjW4OqhXdJb484dbs3nGyUJ4hx34AjLVmKsT5cmaBuT1o7bn
/XsUNjc9F/MqP/6YjLkY1YLGZIabGRHu4XP64sQlWPmwH35vFHK6R4mVBZwiLq7NoPDAUMSh7fBm
+22m08CZyw0nq2mjhT+B/1RleQnUMB9h7gpfP5gFSKLVslttk400Dhk/rpsUVVSabItPuUpC3CTK
XQrnWL4/snv5GZNfbtnMT4kVtjcbn9tWMZLBEqf+C1+R/cJaiBXF3Nhd9CurbmdbJQzbEwjsZaOI
0at0IqgMFD9A3zrPZDiQ+TPbuTFk7BWeEbawbujoehE5cJ2w64IqSy9yG3PN2J4SkdYciyhXGuik
LlojH3rR2cEJuO9OT3OX0g/H3IL3XVX9XtcQugGMl4EsWSNphZYFH4mxn2qkqqcY/IqzWIReeMo6
zO6crKYLQES8YaQS/JeyQdAQmb/Qm46h2nEop6OTUJG6SEizgNiWVSA0AWRP52ZfK9Qp7uAbgbED
Idytk60Q6TAmYcHYH+XgVRXdd+nu7TyzJsqMq66VG+O1BnZKZ7w12CAm52Vt4uJnYPsXR/3sPP/F
tO/FvEXqTQf4TPY8Sm9Fc1eg0bxbcNP2Y0UlUdljB3H2aWP53uQiNQOd/47LKZT6AtOPtJBe02aX
530esNtoqZFbQgbj2/Elx7FsINW/PXrYk+5S0BP6LDTAwcKs2zhdRJxrMpYKeP3KzNVsGGxvRJNA
HlC/WLXUCWwlhQIkJd1RM2mDuoC4+HkSE/oG6DLVtFeJK3qCx/NtcMMhokttklXBR+X7E7jQLAUP
K2MzwiI1op6PP/P/W96kQW+r9lX0Eb9pSRJKbhCSht2p/fX63RRrCZcK5mwH9JzLd89j8YCEGhXR
RKuPk6Frc/jqqJUgkhPN6Z1cR2QW4Ez7RlPPtfmE1YsXx2J5VGqzFMWCBn+9Tgua0m9QGH+svBXz
CQ7IB0yTt7vjF8p7raHBfm/ZHb/BhnLXWdV1+AXwqQtYnnynD2J+MjZ80scqy8xqCCub+s++Wzv6
F7E4BGTuLEYY0Q1SJ7v6gZYZ41xStG0cUl1n1gMekkW1A0zxhvLtUhqGharLF/FFemvgdjr9fo43
Alup6kLU7O2CrtaO+jMPVgWdL2i1K0AcUJPQr9na78Ck75nWctOsZ8o8pIHAJHLJtM4/4Y54ILL/
dECnmT7kG9JwTLZqJnT0c0E5Xy0ydflkYYCbFXMO7oWjuhC+rFsbpGcw/FmvOKH3X9uMADiSV12j
5Q/x+0x+e932HxK/2J8toFPPDhoHNeDwO6Qy6MPTRO/zo82PmZjPF4ov14WNsScM1hPGKx0opIo2
WLzSKHgt+koXQYHCWWX+Bxx4Ws3XXsv0RXzGilMIYKxF98a/GTkhpO5on/qJK8tgPlItnARSFHBz
n08Wi9h5NRYMVZdi8G780e6whZlerqCJxcPpZFpUrGaIvUCMB0mpkVDc5B8Tdiiv+6yEnTlN3NTv
GV2kBREHWyB2vRdSvPlxu/WXmRXrwyaCiwpcjvGMsXvKEAzCRQsfHeIUdOQp5ipTP/+ch8XD+foR
mdbaeeUt1tnLXuHsNpnoeOkUuqupfqmTN3jrflNsc9OqnOYPhwBUiwYYBy69e3YgBICF0PU7suAW
AfTuAGSFCwKzAgfjFMUJTh5AFyl4gw2VhCITaQStbTX4IvtE+3Mo0DRMfI1do+RlpExi17waxA0I
TiP0V2jFA7i1rBtru8pbA/Q8/X/y7HZFe/AsZJF9fhdKNQLnimz76NCPjd+6zs/01o6VR7oLQncJ
zM+UcXQlM2FIp1DFTAShgQ4uADtxkLchxLGO4ZmKP00nnkVHaf0swaaBKDnkaOazp7LMNa8HixSl
kfxPNFMPwygfSnJmc0en+P2QNehgEo7lEN1H7mFWoNCzdGY3Iqn6AZfHSKyDc1YtkaIPNc3CFcUq
Ntal7grf6Y6spVvGifKG5hHFJHhu2FRLpQxUpxOXG/KBROGl/9tOPFnJ3CXyx5bW9f0CdcfYk+FY
2XijgXmIFPPH3xOoAHgo/viiF8g0DbCvbFFwAnp6fzSg24BPo1pLtHgsJoD8M1PYP64quWqPhHj1
Vqwv6UwxZDhfiupAf6c6ytXOp3OeiiKwDVdK/fBILtjKD0LRbAOOcQAqCGXWFL5uWB6dtb0Ry6gS
qRerq209O0snwHww4DLFWcbp7kUCEeNB7U1E+50rW/mCaFWoieAAQ0OApl0jPpZ4rLn8O765/2hs
w6YTftEGHnYbZX0DtYQSvFOSOXYud/aCZBizFeNl1u6vmzsz64Y2iX38RSF2HZIs/hpuOqSi8wSC
TFRgJi6LuFtwjmwXh9fR6BzQ3S5u5ly0EdeDHkcsj2rJo0NnMwDiiQAMbQ/7ZBGoYL61Bwr7yy8o
DJo0Phnv+LyXdnuXm9Vg7I1NBViCT6ryQjcoQMcll404hMv8bFaLMuT3zPZkEc5TB2ehXM3pvAsw
X8U8fwL9PbDdfbbFoPw4R4aL+E9UhvIyprtqumqiGBAOcnP8DjAxHkt++6YAgBDZ9bCq03kG5W0G
vSpO5mhoErITS9Fh6EMx3l/z3cenX3/0kFZLR+OyAAO2y82i/rbDBsJooSoz+5S2PHecwRuFQCRW
vumNaHpUeLc4I1RJlnMN8iD2wGk5v6tJpxlgnWVACfGVGb5/ZxQsT3i4tXLI9El+G1a0Mndb6NfU
IGPW5AddrQe/hU+nue1IqWmGM/7e+bXdwAtX2mOHECLlzpbCNM/LZyacrxiJkfA4DXwBtg7qt1f7
eVa7RKgN0dIegrAfVbyejwFirjCarKZV6NWwXpoP07zILiquKYN7b7/vwwCnt4OXr41IaHCdJet/
QhikHoXdoxeSSd/groOQhpissoHDpupDgo8Jo/VITCDxMdQRgpRzCS7mtTv/MZ570pnG7QwsAL70
RDxCfnNSwvwJDDIaL1obBG8JwBQFthP63aaC07SlenNQlXloMYQjBrXYhfCWwMZb4lNtgDqmoz2N
cPjs8YPN6n25HF2ahvylUS108eWH0pmSvLpn9ncxoUTIcHS5oRK/eSQNAEVHAgnWLqGSSsqywI45
glAn3X1+6b1SMMyqMn3MgIWpshsIE52jFJxdmmFPwBFVEpN9TpSM/Meeu8vRbTE7PKzDV3Pkyd/d
bivcPm3b5HCv47jkzKJLjCPcdy7ARLl1wL6P84HmtdX3j99KoFejgKxbmr1c/ItYXly9NGtkdNEX
mKWsUCzf9WY5OvwK65779GH9mZhCwCuoo9F6tAJWnrdkhMgeGbrGX7Ddvtq7y9LCrUEOMQMHmzVn
ElZN4OILY3PgzCbDuogU33ekCOVywfbC+LNswEN3S/m82dsIz0KGtnxNmWIC936bPfE8dTEs0CR1
2ty/DOvBz9XlM21Y8XOgFnCrgTQkI0cUNifA4dSFdXMT6MpH1uvhJaPFcTE4szDf2QI1dsYibiLh
YN3zQ04ZZ/S7GfE7TtoM/k98YvIs4DtXTKLDG4U6gTsNfP1+Ygaj1/zyOXE4svNK0oUb7GUSVeUg
v+Jek9M5Dgcqzg7w5FDOtHpe8DYugBM9+9A6vnWPlJ2gKudWDav/Ri1TCKI18TP40OGjvy1BLROH
5r9pvc5FtMbOv9k/X/hKRbulYFPqqeXcRF0LXiw1rbwi6OfUOWQ30K+2741La0oqDoN21NDag6mS
JIuVeSfhcUgf4Q5O1PiecHBFbQGnDPnt+nI68+r7i/aMOFV/o0Gx1NFyCO9ewYD5b7vnphNnP/tl
twupsS4LkqXdyeAsXO0jgrBR2pT8cyp2yi8Nd17oaf5pM9iCbdqeBR84LgNJDgXgTf1kynvyj4hm
9Xo6vj4LBUi+hm/LCizd3+rMrlKF9OtMH3FtlIrtQFLPRstmEKN1uLOkP6/d9F/fbkwD0AS/MHT/
uJzAeF1dldK9+VvuOol28Ncd+6kBDcnwjZGjg5jpXa2PkYBACOj8UrjQAhU1wHa3QZgOqwIOEOYN
7NQk6xtriSKWyrzXZhLXJOikUpDH92cLthQj9mL1gn+RNSjkLumYUb2r8lLN4vpfTOqhxM6cfQvA
qYBFeLD2Nk7N2cREANusQ6pNyoS2bQ14GF1CirE89FuT4oITQf5AIMcQyy35ArhvB8Qk+9apt8bt
KuIhGS76Zx5Qcv4JBHaNVkwUMMKpJMRAJ71MAnVCSs5yHYTNtxw68/g3iPbQ31YtaVZRIOBFz/I5
GON8FkyQ+N5G2Gr4wjEgw8D9TQ+Heh6NUj62IKzrzQ4xLIhGI9vav2byoVOrI4h3C1pAxC4zGf82
Siqm2Ku7jOORLwcECET2KjGBTI7+1Yz3k3m+WvC5M+EUjqAWyv1c3D0ZBg/qIKX0rVLlexla5jfN
N2TiQ+sQS4xyZNok3KeU0hfuUo9rs4EZQISKkZvWM2tiV/dJTMN7iDjADB7wdbL3sbPoBw2TUdzf
u6dJIgFv06FVaRzczK+DEfswMFBb/8VClUtjfvcU2Vz4tj/NPv0Yzz4QleYQpUX+8i/YfGyicn3q
JSV27/qpsarkLvGN52aFDCSctd+QBUm1VgzZf4sSpKcQN0uKAKwj5607d9qHl7+WVuvkBaZDHvIF
FcEwOrX+nQLmE+MwBQtDLSX5EciCCCy6BuUfh38P3BbyB8dcE1Htda2IZGEpGLqkkW7wDx9qV49T
DYgUTMl0iv9ATcZRvrP8H4nXYkZpX31pskAa1yczSmueXHRyR3OqTpEWASGgQA8gYxhyWxzspCyq
YLexgQQWJc4WXphc+7M7ihNRwsfiuQSVsYYGcwKizv3xpg5QSI5V+9jy476o4R9z432KSk52Wudm
du0SENbKyGa7yhPgKXAYr2bZW3L+CK2sF6M0CnXGfuXx2g0gfOUJ0TmF34yoanimXEszbHF7dCeO
T6qJfGW97RCBR+EABvB6d/gsH9LldXJHNOIJsd5TWQZyXdH+zXD+TkjMSRuM2R5mA6LwGcOHBg8R
pD4awqpF8XYL+3OEGY67Utmtqou2fdckOB6MrdEwlAXbt7sgQRhKo407SpYUqL298VPJFYyRlmgW
Q1gF7HBo52hCgmnP/ZO8X7fI0GHkAIkHEQOCgLLrrupzK4KdBuZjON1AtK7XKnfRoZ9p1/cnFaFh
PuS1P7n6L2rSv+NUsBOw9dNh2+IwFmtMjX+YNquQ5odwHqisx2khURKbZoBTRtc5RdgzW29DLt+4
PmAoxHhceZLAjR9EZc287XERNsFh2HoozoeIJ2nAo5bVsBf1hn99fikcgF42Ma5LL6BuYJ+Ak7PO
IiXPj2i7jMBPFoB1/c9TklrprxcwAgcc23arQeJ0a16uIMUbqwTc4XKG4IFd4Lb8CoLOv2lYyXhm
QatqNSwhKKgaVyDsqBWllSsQtk2lxtUHHNl4lLUAfJH16RyezdkyfBeuUjQlj6wVnhEJVRtLlbXd
lS439JQ1dHcs6m7UaaHcYFv/s76avBbhLZUI6su2mEy5GqWXENfKtgQn6nU1PlrIln+ZDuM/yvyt
cLk+CKPvYo1Aozk3HTGiiu2GOsGrc0Ees6q3iRaYyOPM0Hri0/B/30ZUdDvKpCBCw5T5hXzyVU6s
oCpAo0GhH6JuvndnCbiFEQJpW4/SUz6rlYPzrXPGt86CHguTAIgN04OmJ82ro/8RQGPuepbzhkzk
0Tilep2kKaN7XiSRhcGIuM3WbrJhj/N6wvX8fgZmtXdnlarG8SB4v2j4XZKtBZNL8ReWFQ6oHq+p
KZS5sKc0+HuZSr/Hwy8eQLrfG2hRVMg/mJdGFUaLXdrC5GdMmaRB4GIzMhME2vc4A49a/bMslPO+
LFuMgEK5dHkjAlnD0X53qRc9+rWTZjUrZ22ozIn7cjszaqHpz/ohvhuWj6dMsEn/Yk7AahEAAHcH
W7bq0NShTCHs13ALr5uR5too/BMBx59Y89gq81ZQe1kCmn7JOOBJ5Ot1I7fO8fWZWHf4+cgJ9HOk
nejBdpvSlibH0+pvZirbO4F4g5LaiF/XDVNq+O61AcjQTGNKQrJk9zCnhO/LNvifkojoCJHlYPc6
D5BrMe848r+c3ju88WziWKICWpGOO2EsQ36+4Crm2JwhplxGdEPQia88wkazqNGQx8pkGnR0euWC
dgYkgXo3rlaZNu4bf1YxOtPmqf5v9PDALTAeq1R63o4DitgRrfdiq/lHRJua/pE2xOvtnMsS7/jR
WDSoTHOJlIbEQFVlyScQqMSEX5ljiMZ1rJj+payQFvo9zvMTu5p/mYtEnwwft/12eAwizhQS0aYG
kzQc66gRqjwndgY77MXeRuK1JflL0ne1FM4bU48XkC5xgGDVAWqzSVE2IwaQRRMG2GqaA/aE1lfk
ohWenKjB4Q2iQYcilQ8jmlIHKKiBCxEhfUhG7a3pc5r7AOVBMRkn2yiP1BEYvCmgLw86NcBBWSRm
VBCb12gCHG0VYRHfDV6idGixvNY4vWl5I7KAONfd4LmHAvocNHtByOL+9sSEMBgzurIU2Us8mE23
I/I/alIYQAtWxbwfw1N37RDlCfq6xcs5DUg98/bRmgOVhlKG/A8lVA96sBo+oBlWGOruIBDAvKLN
PRH1rQCKiS+TcWxWDKoI5N0pIy+oIANCjsUrqmmybPBxZKIIjPJJmGPcGCkRReVbiRBNv6OryuDJ
bdjL7BRPDFtZddlrfC66++VtW9DQyGdvUfASw7vkly2fiWJmYgOy2wJk7KeVJAJpqKYSvfbWlTMb
N9SKeZzSQUgwK7OnmoPI00tMrUsHYqgFmJJwNgB1aJy97jrDw/brezijvhVTied4nkmfDC6Mb25U
d/oxg3HqFTmmiF7Z8n4310khGRKaEpjVCbFbCP/u5Syr4ajyMRQbWiOUyqs5kBJjMy3aAWWSAWCB
FmbXUTIGWydVsvgZQ79uRtti1ITKHwWBkKx36nt2Xq+ITFrBViJmNhFm+ItZt6lUPkWwUvmBhWTY
2yhle2oZ1V0LQ99xuXvFiRQ21ZBbSy5hoKhP8nVIhYCYGi1llMis1miJ+jpmVfhqUxMKCkhsmTi6
R1T9Sceg+kk0mCb0jXePhVu4Y0iJtJlgVMk5QNxTj5Nb1alZpJO7OoSx9D7A3El9nzBzUdrrxfTT
w5fLtWsX3GyuvbzPudEpCoboZ3ErJkJdrsogmULAtCU4ATsVyOJWHJohi3fsseKTfsxo0hkpGmlJ
+gH9ayWwFjLKadFHIQbOySoAzGiiZtDYYLzu1AtNWYKLgvCtS+/FNuLwdWBA/OzOiuwcs6oNWziv
vuQcIyocmeY5R+32QgK2LfsyxIVQ/HPF8dEyxwuX9oHf3vo0NbbK/61LWuo12HaFOE4k8O78te3R
NbaRT7CM/z22Dnalg9sIqLUQbgnMSig5C9Gyvo67a4RdQj6ttULttJjNAS98bm+WmBBMk4OB2iRo
t9GQOvrOb45jcO2sn7Os1ombAKd0nnJkfiEdEGpnA9Vx7FZ2Gb5YT5XIwLPXo6g0Cd4hbxSD+Oot
N0M3TkGg/5v1NaDjfCj9Pv/cu6C3rC+pSSQi3yg0HBVZb8G2gXl/EM+X6uJpmvSr0jt1mB3whBrD
g2nEd57k+LD1+BqsYqtTrPEBU0dntictmZSWInAyaMiS9FBXmLOIHFt56KtjGgGwvu2hcypIvOnZ
yEAm0vvkTm0ej3yhSci1OpX76ffp0NXtN1HNg5Vb2W+rM7x4GyXmjs/mUOdOY+RE90wH4tkRfhb2
b5DgZd+XK09cHPI9rjFaBWxQUIv8cXhiVXxtIhkBa9d09smDUJYo0BGRd+DT8jwUKUaIqIbYSmcw
OpXjh/gI/yGavRlUoKxsC24wcsPc5sqXMIksJNf+u5zr1PaljbB8NqYu1QMA80urCl9EeprjKYdl
BBkkSEk8EpgxeWab08EM1p8/cEWHgFTYkjuYXK81yX7gLEKgQCLyqmbRRLvBi3pozzQTgghJNQpf
5FOt18R+Sh7OqzGiA0neYx2A7ZkSiD4XI8zgn0vOP/DnoVSeKpkjzEKEBHZaFDJEY33LpakO5tVs
J63bT5XiW9piQyzZyyMPDOpEdgQC4oR9OU7xO/ejXZWWcBJkY1/rDmzZRkitiik824AbpEMrL3cC
Wg9I+XL76wZwHS0dEW3284sAvbdjQMkAz7pVEcob/3yw2NSWQaZLs4jQtWa5ltztUoxwRlG9xENR
ZuY4Oqrcdmd9QW0mhf0uu3V9zpAQkh/VNz/VTb0b8YcszK3Nj8CKF8wV7mtW4cei1ja/aYNdQZOU
cJAXHGRGa3U1p7AsgAi16tHMke4ZSsb4kiZ6rb2HZcIhJfEcWj4e6x/x6nKSBT/rQ/j+W9JcYQCK
OZXAxedb7MOc1CXh2ymgMS2DNF45Knkwv+C1qoVHvrWiFzzQH3F5L5qlSyQHUquraE41bGePA5uT
kt2FIT8qo7JaKVMZL0fxUValfJaKfyZbYUfvneRmo7wHveDtwa8PC6FciodCd16Zk4Z8D4RWTdO5
lexpv5eddvB8Hr/zUS9fkBjd/EOKxOV6AKZEguXNUf4aTN4g4gucgNvlZBhR8AnXZVwrMWeWiYyk
o4mXLpVnxqvLyTUJT6OeIPAFtDv0CLqu5dOIty4VUQpUQPYC+L5UMGU6QK0pV49GHADZPq9FF3zf
OmieER0MIWb0iv5ekvj8qL0sqinSWA/pDh94qcIsqzZnFjrvSg0ryS+G54VlABMNxZMkm4LeTpXQ
xSOs5gvHU0HZq4adZ4ovqNhbyxwV6BbLg9UYM0+hVOoH9UW2zXOovz6eTgraDUNT9SX9i8tQA69H
6l63X7N9C02dmszrckDxiOz8MZlYZqmYg64p7stN9lHZRoYLiz9SJz8gYf6bF/SvazS45aKXhO5L
CaxpvhEEHCpwiZr4VIwC5i4UCF4A2ZCIxbcs+6oIR09+gopLzo6e4+9DUNwqFpU+mdW2bF6Ym6Pi
T3fFqfmLYfz2VVk7czFCVKBprUaQJoVeh+k7LtZ3QCCd5KYPfc10Vnb1wjjCj3evvWMmY5T41MEn
aGWNz2QirfXmLa0/u1tO/8sWJIIEGRYiVwQCK1wo8sU9jjFBmuJ0kZT0cLcF3TlU470ppJvkoBhX
AJ+UVbLBoAP3z20Y6DCDbuPGN/PDbrseUsbB5UzP/lGW5UZBMMb8FgIveVrtwS492P42YjGMZfZz
nGglq3UNuOn5PmfDI4fPyYZe0VbOWH/bAQWxiWRZ8+4OqMvNE+Ajr6sGQaXk+rzJq1RCXV3F8v3M
SUvkEosapkRqvNMZeFwI1XHaCYIHr+dW/fD9viwNWKf+izZas69hQ5ssqcTaDiMnRPJElFUuNJ4p
zNLFVipcdls/7eZzFhT/UksxU6kX2W51A+Ti01Xvl+lcfMsIx/2xEuA83AGsyA9ZK33E9xB6zr8M
yt5Wh8m+pZ2bucV/ddoEzjlGzLhce6xehPifYIs7seUHRccxrMiIu8DKM1/+e8UmZ8ikNSyG6PeW
/gWrhckd26lh3tFwxdvOHjdrWnMzFfKq6LHpaQXQDVZFjDegaN4PTCzxIrpHunTDFYA9iQ8HWh6J
s6dRhRvmnXwmqadjjeXDi4Hw2+SEkSMeQaTcj6EtcnCQO4HtujP/Hw6e3ZvkJhVebKsujy8D21ks
LvPiYuu+PQi4LtIWvp7ljZ//3PZttNopfCb/GlxmLeLwklnKiCgs/bi83DnMh1ZBrnHud4nJKKSD
PHYOq9Rc5p3tky/4W8YRzTnust0ZGXjuue2BdTUgLzw968n3u4+iHzH3s3AfKdW5S8daT4Sy3IYj
+WsVG3NduywVfFk8f2dW0lpw6eDsZ7ubSTuP0NPI6GiK2KP7tUNniSH5ja9IfmF88yn/4CbND4dy
ENg14a2BasdOMEAp/h3IkpOsqlANEKglfIKmun0u7q9GCKZve2K74NqNlv2fjR+B0J7rrwxoRK6T
qMg0pGFUwMTKqbn8OKgkAjsl1RiJKhgPbJHYZNei3djE96rcHQm1WQLsieUYkTnbhZn99XaxEc9v
YEyvun3wF74GPNd6mhPnB4X6tlLFd+5Ol6NpdebJUDR0tLrbdAAeVD3vtv52/8+pQg3SIa3muQrk
clpS1rKxDw53jr35MqcajKbvW6PzrZJgyo5WcMWwl9QhJzBJBnSxxLd6g38RXwYpwchLbw7QTFmU
vxEvq4S6N1/Pcb6i/QAlp6TGPxArQbAkX4D7T9dfXSjmvkBuJ+NilfG97qzQfKTPGhyT3gKNW5FO
rJga8x0LM6XfjeQN2n/4qgKj9EYkqNvoykz/JTB+FK1YwVj6NzlOsVYOVX/z/v9utDRqE2qGtvPT
haotr4rzuGb//O+AffzRqnikhFbFH4AG4TdHCUXq9xmKkFOf0d2N4f+/ikAtk/+v2oPz7lDWpzaU
Kw4AxQBSY7rjoeA6uA+sVG9AQx1FEY72lwPu/t1o0t5r9DzZDggVNPbNekn9y6740AkwZmul2aEM
k6WYjuYumh3YCQj21Jct1u3+KDWk2jHjJNo1miobL1Qrfdfzp8cxUNSZ64U6ilmicRT25jSOf34e
dgBEJnTmul36+InwYvlfsHYhNS4YSTiqotkrqEap6ejNLmY0LOUNtyWCLaBR8taILsnXEoypYRbe
d9YjPnIree+8Xf5TN22bRncnm5fVtGoUNME9iQGRvQGxtMcBQBqUzT8rJ4+9ShVnptNgRmY4O+oC
gpTUnBb5R+pnpZ8JGgr6brdI+u6IDPfJwMq+yfO8UAgSePDJbAO7XXslPIEJ0JzFDHn8diIAHi/e
/CZDxjUDLG9CHqVY69FB4Z/9hHixmTAvn1sd1FFeM5S3MqISaSXsTr+GNoqUH0BdCgZyYDpQCcE8
jd7wiDW3Irlq8X3BzFT6F2lYFnat0dqlkxoXIAEO0vODwTer7RDHm9FlZO01yPXriuBl4MlpITVX
5tVQbBE1VZvwz1qx+bGe7rrCxtTR6oDUmjklE1YqJLZ3GcfkbJwKiqy4Iq3Z2iGT67O0iF14sQWi
w4HMCGCpiH+sog1TWTyWGpV+f0Mi860k4I6J26FnGNr3ybhJ/aznP2tIWb60CHEXwzlI7TKULGgw
FIrBgxMr/95QB+Zr1dDt4nrjodjz465Y4F83r3EQfOiWFyG/mimo6Os2/QE2mwRW96ChZPhSP1Ui
5BCfCqQXhIu/8pM9kJ2bwoMpFfECdsJmNKSl4j9lS40muCv5sojoyndvyjT79ylVxrSBL6o4rnOv
vnZjqMBVRcN6OsTk6kOPE0jHdKFaaD5LxAcUkoQsei8qmZKfAOD7BoKpNtPRK6wFVAOipvd41y+j
rjVyVuXxG/LDnY07H0biKjFR91L6vi/uX5p6U3/mjHnYNMjKjIarXMFy/Kh1SIbYg8xcngps322g
VbMVgCXg+m6jelxxMl7pQ3sHoHXJcoCGPtVfrI9FSNeuIFXd4KAsgPxLBVYBwLUruIxL2y7CaveW
iT+PCzJANEpKsPpBo2zEVopvZlz7M3HrmCFMpyTFBJPEeaJqk/lcJ8PTfWqcR6W5Es2p+iVM6Fp+
GdM275WCalr1UkJj9Lck1RNm1UJh7OWXr+Asy9CCuUv/Szr+/CxqNuwRH8/puo8jyJbESPFVxZwP
u3+0elFytZcJ4oNWlu4bzkXbHS8Cz84C/ATsnkcs5jKsAcvdMiAPFJZkD7NThPryTsKwgLUzZGNH
6q8bn6yb3/xMvergy1r37ZFrFJkP1xMliJ/CWxfjIMId6A0BAy8c3weoX6+NXWvtOgUskZ1M/uXO
hWqaVCBFICvWqjqcVIr4Edm1mFoqrmLC8cNEkSOKVhouasKRxJ3mICGHIXhDVhxYYq5QNWBauVC0
6B2/IUkxQEU3KT4yaW/NacJqv4PCb+bQypojIer7ynhLdxipqHxscWMS84zW4nxG5R598Dfw9JgL
WEpNlP/EE2KLqPFFez8JukjfYG20LgdhBssmPKIQuSLFadHtk7EEv+rUjH8AMIuVryrQg0MxGnov
umzwsTocgE455BQAtNKmPbFKtLI5C2nnfF0AUF+qbN3IHPLGJbDZP+xu0GtPV4hjqvx/zcxodr4E
SFnKGkVgQ0P+kMr5ndt/r7aGhjiDn13frZIJW+FhEolwIN3ykXFRMO6sPmLd9xkcaAnLV2r8XOtj
dFxinFtPNVQB0Xy3wEcBHLMB16LLqwIPPJCOAHRLCs22sQL0hJJY9VR/jlZyEjju4eCOz4k5ycf7
ZGkqqL1VwgixNs8vVd2Po0/75ndFSokzDT6sebrnYIJVW7p1YLBIIehJvm9CkysMP4og93QidToA
AeoYqx6eHu08s0F1G4KSyLbXD/8xPGk73eLnHmtSPWFmTxfsntKJfBqWf0W32jnOXG8YWJdyND5L
60TT3DHl8uW6Op0ChcpjjJlnmUWYfTUrbVKo/Vm/8dneO5hOiTRXovlQj2DFPOfgm+7Aj/ZskPXT
8C/uaOIO3S7tHiWrCKwoyPl5Hifv6U3SJprB9W4eCDbVZ3FgUt/7vBA+lLYJb3BmMIOWIN/C2QKP
5O/L2Rq9/XjcBWxQTzYD5fbXCTwg01YmDYL8Er1IP0M6VYNizGnM4oDJVHxNLbTbm9G6nIhTTkbg
K/OajPZ/Z7U+PvIWpStc21D2yp4H+fvS4Pc+JUxWDhW0tuyxDG99Qtx3UqzZ3u8x363QVnyOTpCM
N4Ll3pKUqRsoXx/9H0Hy1stQzoC5AJgKxzrvKL+OKRC9WSItyYHNCVsfT0zbZccAtyxXYKhA0cYa
YwT/oLiyISdA0tBH2O9yj8utGGFLECnwZCdAfpwr4kmFCJVMkuTyHCaqBJeOpYOFAIgk2e3jHm0+
SVMiqUHE6jqyr2bo8LKC3QVU5oVv8CdUAu3+NLcmdzrmd4uUywplJvfz8N7sB1LKr275j5QedvN4
Ldx+myshe9DMWGhQ284eHlpgib8oHlMuLhlVhOjTmsTAMG6VCnIqWOKRZ23tK7291bxbPCmwzYTf
axenfpq2edszWXsOTD/q3yAoDBh5ya3R/PCHKIIxu5GVy65qpuvjPiai7uk+wil5rW5sPOHZGhaa
heOJzd2dmrvO+mLxO1r/cR+b09WPmqhzJjmXecIONTBRUKmeb6x67BSkVLzKdHzyvMs2sZBtW8+P
vDrLH6zix+CiEUMRW9Q63JhRKuCeeeiTeGvGPmODDOki3jYRhgteCkEflPJGZ+jSjGhVtehb2/pe
b83JjKmvegX6Y8DpT4VFYpVFqalNUheOJ/QMS7dS6vphFBviyb6psN4vesmO5uNVHOt8b40mDHdW
hy3x8Sq3TQTyb/dpmVrJNY9x85iAfiNRQh3NMfw59CFzOMYtUzZ50lXsSOUL/NyUvLgBnlj0sAI0
Dd0wme2X159ZW0LkdYOXPZZN+xuuxrbrMSGjMYbGwDYoZrybStNWyYWamH+Yaiq1rnPxPr7PYlMI
mDDMQ0efUf7BA6+3muJ3VCdCUIJsCIjw0IESIDeRH7jVK0SbceLl8huQjzgdkXjvAw2fkJH8sZ76
UnOJ8v5L2e9ZYAjvoV+/9Gy3SRK5sbs5R3ge2A+iQFbp7GXIw2aQIk0lI2MFiNWlitFN/pYwPvg0
YCH+u7IRve0sQHtGDcaexs6kOGgG/qRmGxvajejqDfrvQ5bq9aJDmucgEKBgZcSPpsKvazl9LQnR
GmMt/lLkA6AcsExqTTA2sLV4+XnxY0bMW2MjoW3CNR2HiTsywgCCTxXlsGfZyupUnv9zCvSPTKP3
oKzOSb1wtOCoVgKNXGm4C6Sa2LmxlfHS1WMw/SjED5yTHeRBcitBkwhOrKHBCIz4HzgKonqn9jpb
HzDpV64lnj0Rc1B3s7RscwWwYipB8VbzqmBa19uZCfQyT7cqh2vTdwjAa6JsNKntCukhl+rz/+qN
90LBwobr40xLAzDBbAh/PRAPmT4jfTnp5mlyfHJgtUcOFTds4lELOxEkygpJFFqiPaCud7o58466
z8VeVNRa2LAuCH36TYLdrnU2jcafGDoKPcFPrV+4M1m8A8oZfckxOfapUr+AldKRE5Pz0SyplVK7
8jsu28qHW2mBHq84RqVifz+trfUhRpAUfpNeGcGNlai4AA2ZnwtqqVKNB1WVEKDfQ5a8cXT80SH8
47+NtVE6IGkjmnELV67P8sBLap1SyisJAawG3OpEaasCpb0nA8LV1oj1A4AUdty8Hb3yv1iPLtZ/
+npn/PL22sFNEwXN2P2Et5QveO6GuBEUhv7eWuAaQSYpjdpCXn5euvDMF8BoASHFQ+8htZiXS/vc
b0mkAr5YnVGLSzB6OremKLYK+4A/AxSWG33ceskuUXEHvaWEvvD37Sp2TRIdPCavsz4sU06Swq7j
G7/g16yvx1YvL7OF7Pk9dPIjrrhYs5eupmuRF7ZhwA/SwPLKIu8SklsezaVBQkfglSYiR6GBikMO
YVj2lLFPtRWZI7SQ+5mLPCdOzdK1L6oPmnNc80f9ONTtowAxRif+5tjI+SEB8sh/CAecxiVGm9gS
eHPfmX2iTd+RP20FQgKwYIuqxEOUiUktR5AqPbbhpSU9cr4Q4LEwQrsmJAv3F0ZfUs1S1oqIlkN8
lTY73kLBpck6EPKGGWkcllEAM5skMLL/7YoM7aikn6V5yLxUHGN2ljXV5f3NvS3BGvmw3/4Z1kvy
7tsp5L+mCAIOIkVVhj86H79E2UogoqkSG1hXdheMYgFNo4uFO1KSWptSTSikt+ej0Vip/850T6rx
CI8svhNYYAR9+S2ECTMbozVa3iDsE9YfzmHEStHjVpaZQVBmFvJXlGoJ2ieBU3xdVLjhv4BzJbqN
qBo3od73d/k1FxGK2FI39UhAPkS//t40n8GxXS2xV0U17dMJYRoGPOTebkIImJB9O05YL5k3HeKh
loGwgm769gNL+W4EOFZLwdXuku2KYN6BkQ+T0mxWg8/kNhdTL0m8euDmmoplMpTvb5qj01BKR12s
HUqFVX48DZf3ZxmIhN6TFmHKj2nfJR9z5iXG8VTAqiOUfN4FyQR+TN4UrvOQFe+wtBdBhlg9C0mD
xhiLIf0o6lr91PDF0ZKKp79Pcq309K80icCgsgzP6RQFl6Vub9188A7xyRB4L+mOuhsElEfsrtiq
kW+erTlxwdHmZTj0hloOtiTOyvOSNY7U0ile7QF8sAd6UptPCMqGq+o5asUw1fCrAWRd22PoR1at
0Llrf3CGu6IH1AZCUdm+DKq3v1crFlGVcVpjSSdfQuajMWKYuocLpyz/rj2Z6Xg4XnWB74S0CO1M
Px9qbcDhqN6E6CYMK2sRC4JcCLLW13b/XTjxw8/l+NCNHxYRJxckNBgRNYPsDexUt3JaLOhKv7PS
swmGoms1xHPywjYPr59rU2STdivBlBybyPeRDPnWV2kd37mJ6Mm2Pl4VTGA9+bncZqmT46I6AFtQ
GllWKFUomnwQ1YPUCR9xY3gb2TyhRos+y7S1hTmCnMmGbTW+/pMamLl8C8Fm/3YL2VepKz+JwV7M
bllBnutT4EXiYltD56GxFPznPNMsmSC1BvtodCRWXAG0Is/YmLxPPfF9lso2kHbFvtTgqQTQPRK0
if6LFf7C7f0TlVnfXwhDwhq2W1E7HZzr3q7ywci5NK5k0Guc1K+9eq7BKRv9OGTXoQ+IRMcdtukk
OLT00yDES6u3SYpWu0kVp+meRySk8t3qRAPHllmRcyM+JZmoLkOIEeS5zjGHZroKyOj92iCHMWYZ
kZx759jXpS4mp2PL3WurMuhDFPYfFXHI+knqQLht+9iocC8oILcCedVJuF7JQMFP3S5J3hChEHjU
kG+1Ck/uyMZkolVKXdJLGBKmjPJ4gOCZ9KoUVZM9jg+S900wsIswclLTCxCI3JPgTj79ukEE82Rv
tircKq5W4+TxxYQIG2/s4394YapDgpcM1uKjIznX+WvSrX7tR636cVAOh11o96kaKy0pkRskgHnq
sYUSg8idDQ034UJqiu6/j2mw9brPtEx/m0ir9HWMCAYkNfZT1C/SmLxdulWMXpSN60GvVAiMdctT
5Jcn+avwG7RExmZ6AYdN2uGa2Cuq9GrgGc9edjwOTVs41buQNuU4kihv8nuHYebU/JqzIKffxNIf
IrY6PaPTutNeg1bXXkwVbQ1JJqyxpTh5nh2+nAiD7FpOe1P6mXwN54RBlrfj/33GYsdktEDsvfjJ
nApH/u4dEgmmRVgqhSLchkCA460FsmIQ21QavUZrwJXUXF1Wt9eiJFNCtvMq4n8tUzsNgxWz14+Z
QlOL5lUZJi0r/KHGfkKWsnvpb9SxI5vGl50GbGPS+ZyLqalCQ3EdxhnQ3hEQ1UVKZeTQCKmHjqNF
f7sc2o8QJEB5XIso6gy6Ist0qfRoGcJII9AT8XMsY4okoGZ1jiE6VHwdKKczD5Dibo821nsjVHM3
I9DXxSYkg0MeiSiMSZF+q3P46ZOlq3jXsRcV+xhblN6KOqrW2wozhyejAYXzYgMu8JeOKOCZ0z9l
VNEqZIN7QMuLt2NmP0fvXbLASmAg7a+xH12biw3NWFFEqi8zzixXNUCubtMWZrLUT1VtmymxMUDt
AqAJDXZxTM8+xu5auIXBbTQmu6An8UIusba5NrohJiXKXbm7SGwWuxsWI+i1WiO1IN+A8qCv7k8e
osumRBVA1oeuGp8HvesyT46MkWrqVn63aXTPdzL6wV8Ol0X/3NnCYoOhlbpR0zy/vBpT7DVqJ9mM
/ZDi/VPED5Ps7ZUxAZAdkCWFYSKSCWsTdbN2HjiMBGlj5hPoMQ+Zn9rkxB7lCy0E7C8NAFjeMSS8
Mk2zX/zyLpY7eKEdh7JiF2P77FLox95aUfCNFjZgg+FXPM9ZMxAp96lwztSJCBIBQuFVv+19zT0w
YK07hIXjaJoExBicJ7q6N26IJ5a4tcBiTmxH/igw4KPyeyrKD2cUVN72xGNAaEdr6LLHP/YApHub
O4ZoGWcuQ7BgaY895rmvWJxq0iuEuqOXHSJDdQaOcfqOFpYaix9cHW3E+2oj50ezpEbMSDla2FB1
J/uaaEbGp5Bma5zwGFeLK+Xf4I9+ZbZTsZqjp0yB3iU5UzCXTqLFO3LU3qsnIaVSAfcPKOq5Laeg
9gYa0nOyH1SKI3MnnCKJ5vfvJSdRlRdSd6Pd0XxQDGUErfcVR6vEwfSsvOYo5Fk4yjdaNoepsFSc
yaGiziC8S+ZnsSBDhOHcB3YyUuCV6/8/pbU3sNFVmnyM3GJlGwEbJ9DkOZx6PTWvDMHKv/FtOwz9
JxDzjB+c4cmAmG08y+xIJ4sEpfC7eWT9iJxkZfOBX/X86QlJfQRwhrZavw4AHcZ4wBdqleV+pRCH
8o7SfeOqrWrma+RuSQbgwyYB5O4uNPVx+kwQbEtuFgX0JdkjPtRBOpEiuF050cftftNpm0EGMEhQ
pABYzWgb/txarCf+v41JEhG/UxEMamuTtryOaqbBsgIcXApmeA0Ge920AvAVpICCMzPoGkb/Qf1f
GX49wANnL7yls9huAwopmW1d6zZBf9sYz9+2TmcfwsDHNvLF0enBNnquJQ5PU7kBp/N4yP/HF0T5
cu0T+kTMRv4Gxo1Mtm+xNbFhJq7zaws4ThZTOeiClg9rWfRwWriR9Nj5W0dssOP1icPcy8uLgFDF
skIkYRXtNcULPTf9hToV2flojHc5PTg0XngBrOT/w1pMechPYo5gL9O89NGLqp1JiG0uPrh7krP1
bqj/o7DFLPlvITYaH5XakYV3lQ75QBw2ckix5HWrlf8vDypzf8m7sPvf1D1lyHstL9SWqCQM2LM0
jrD/BehgSWL0+OQJXeDG5bhlOILh8l5Smh7bQiuMV8uDEg16HfW6ZbDzA5kCx79kdGBK2CQTO8FB
AiAOMmsYtfWbU0dU5lmJxjxRSpiJ3hKu7iMAFLwCpY+F2F+cac3WQnF/k3ifVWSZtFDbBBG1YY6p
rVjQFO5KGMMupMten7dOkDCiWj6mDnJII2kyVxOfDl9aJBT7iyzevyzF8imxvMysbCTTEFL6Xk7D
/6cudl7jEitTUhF/DRg9fQlieb6IJy9LygWzTI4T2HByPCEa5xAv8JF7nKLBvfwVGIQO6Cpp1bmU
EKwXSZeqBADS5fLHc/ie18aa7MaG90gWN5iUMZ95fAJG6nby8XzhYNP+4bSnwF374yaj7bhIHxJJ
skbUHjiZuqEX4VS5jLgbXy61Q2jE74JJwuiiU0AATOVZTC/NWRA5jLzkHiKo/+gXDlqFO/60O73B
F9ne3qdE4NOIKjo/eEKcflAjd15mlTpjhw4B8DYHSP2+LNmBLNdFdkCCEMstNGwmF+op59j3wupY
mRELSigC5nvdUFPXvPAB+J19mK/XtMz+rDTQJlV1UXY7lNQ+i8ydRsV2OUyBG8ZlZ8ivxibAmiXt
w7/0b+KFQoKqY0xF8oSDsUEC0Du9XH2Q5VbIXQcP29u2fzCCeAL4prRg5BfSFqJLk6NFaEGk+lHm
kSvj0rSG3SdwXvUdAkP3mOKRdzHLLeDHbCuLnujB5p96WALQ50sNJpqiQZp8124m/0qwTQ78VtQb
Ic8yyD6gVL33+6tVE9dM33+z1hF+Iku9Pz6HgUEvsASWIpLIJZuQj0O14MEUw2k2Ekp1slUjqszA
S3yGWLiLpcYiJvvMtML7nI1M9mHAWexhBaYgkxbU5SxIPuSp8MC0VX5/Mls44DNvpSu5mfAApWr/
PxCgsHbz6jdpx/KDJLyfGYl4NanryD3rane4OwtYc4Q2UdgnvXThCIVCZxCNxgl2qrRTSb2pGgxu
DHA333OjrqpJLQjClNSM9TkktDeno1EpGr4AtapKct03dDNI4Q+j7F2YbBOICWUcbRG9NuLixIXm
rK4NAw9GbPmy33OJwda5SKmh9FlBlpKfze85TmMMpVU0BF/+u+hIvDTH81kIUQWorqZPrlet+v0H
l5NAFegk/PcFo4cCqdyqnzacq0+daBS5MMdN4/eqVQcD3zdy0ge+5uksygHZEzaIo72kGnUX1FPg
F4vVTKwn7YoeD8verdgLIogxANbzW2bNPkdNM/6AmHC2/ugIuWijGfEWWZUAf3dh9IczHWq8vTUm
sOwDWaKGRglTS/jJwIgl4gUgMW/TvJLHtUqDgG/xE0fEwvB3aQYylvc8u0KzHDKQWqvpl4OYBsl/
8/K3cqRhIBMfi/cPM3gXQgYkcw4UdZfdkPyUh2N9E+abE+W8ALM5VE43PBhSUKQJeKU5QCGosFxM
E3DTaaM8nGSv36mNdcNfuT2q6OrHrOaHR6Qw9iTABiSvP9u5mmdBnQlF9D+0UVGtJtt9JfgkxihA
j5E9ms9taiQKLCMasI47Exbdc2kjYDAfVj5Br9RaNzCXCGL03GIKnGj006YuS4fJCSUvmtVy3/OL
h6I5eecR5aBnz3y1YSA/9J3xUS0HU4xwpqDIIaKfcBGLgvJGL7dzbSsxQsDD4aG7hFoW9BJlbtY8
aw6NPNS6fHSIfGcdwDlKOKJt1HTGHXsLS9rGuyyhsxjxAjmfNQ6GkB+CdnfHV4Dq49JP3AQh1aFX
ZYlJ77c9gGyt/dUUcQu90FF2KVJRWfW+I3xnpj7moDPhudYgqYJqbhsx9EM9YKMH28pc3ICjNZRE
Yago5r06VCwJ6xxHx/TwlJw9gliprhExW33RvAUi7IBnnGVVLzSD5WlYnYF72wd1V/3ZqtyMSXht
CzOPeTSXfLoE2YZGsaJrtatzOThR18M5MAHQW4EQAbjujdowlb38NWaETI/Dmy2eBxptbb5pe3Kq
Xta/05oAGP0Nn7YFD3VITqXFJTidcbVSPijFElv0WYzqg1VKgJLQOdV9lTTVGnlhmVdD0TUeP9jT
VPAD5PGPJB8KbJPBDt6qDgFRI2YySHVnUiUxm+A/2KD2+TMAFk5gNGB99MhG+IBsd1wj4tMLk7aI
vybtmxg8zeZfOf7bLrJQLp5hcZalMEbjfW13e7BpP/HcdqwMf0v1ei3seyjzNN790SHn7Eq8SQjm
BapZ9GX/JaOzOz5BtKsJsutsRHhSQpMRGU7UQRe6GmxC3bBvzUXsrxKu5oPI0+EjZXEYxg23+3ao
Y/vtV67GSJupbZuJuUYURcdvaGYXcpWAf2OassUHq3VNhNk4CuhP00B3JjFnUQ7hKBwA/tahaQKy
CrLvNUMQfrvmRbZjoj34smXs1xdNkX460iQ//J0JSmPwBJ7jsjR31aQn/Y0bxUr7O7SVLb2fGYMg
R227LZ0cWpvstNBfqocd0yeUnR5BlzFCXFx/UFsQcUM1AQ/OpJrsaGwr3xxXzugzoxT5M5oPWK40
KphGClKnZYayJrYSr+knOYZhTVngt6hpNxwyAwOcu4lkKro/b995SAzzzg0uyIy46vVs1GBRecNU
jJq/VbzBuTP0P8KxpF8nNwcNO2pAIdUirU3J6pBZuFjVVszM3hk2sGbeVy2R7JZqow5MxCg4akiz
PNN4s2bpJ1kaGoRmVBYjQp3Oe98OoeQWLnVYR0QqGnpf5AfcZwSHtzAV9nCzseAjdV9lahKUPOsc
vSYoTbpBbxWJXXp8nEBeYiwYhXzLq+Tb5bnpzH/re7Q3g2oCn9eOdORTNH3FRY7fjM1cCyzjuNi0
8x+EHfj4qVjwGFyRsR46OZkW6Oer3sSLhvKcRI93CBPNtBQxcA1ATjdBSS5BzD/FA3eGcpPqBI+v
uB5edXIof+nzho8F85sX/btqygiJjJ8kwlHWc8C+AfgnXzoPFLdRzT3rTITMRdqD7kxQoMnDcVF+
kD6rnvN0mEyiYyrg9yFuk/bLe61rL2Vt1q1x2ognVAw0QXTl0+YTB5hqfO/jLKZtqDSw9D8JjyJZ
Y5ymRTkgo1zA/3satLeUkB3UuiwKUO+w5FJsc/iDkvc5R6zmU3fYN4J87aHA8SqvKRb0T63ewkxO
MrKgJuC/lFbwAlu9yWYSgBhz9CwbO3ClMb5iGlPy8DZAyI4vQ9CnapMyzfzPOKQjtcOaacklJcGc
bbiOqqEGy8mHDU7m5tWuNLl3RPqkxhX7B7SEqAatAIOfoTVJa16b2tdBw8qDbXfcHyj5VfHyNxRc
yPkVn8yndIecmzL0gULYAYWGkhgxZVO6Wg+ToB+nde9IG0SfA1CobV6lrRx+wmlK4dDJqiySv8Gb
/34vAnIGjKjLeqNHQ5cewJVAGRW5d5KxQpT4xgRnyuVbNOYSJTaV89LxyiPd836Mdj9UzsPTQYTP
6bf5JUogNppy6a00+cq8DP4eXLV+8smpHf1HpQlb7vFPjB9RFVytA3Shna1RLx3MaA83HyPpNu8h
iwn9MHoAuB+X/koCKczmnQO5p0YQme2thaTpELfTtmFDtcX+Vw7Is3MZjLHFSe6EWjf62XGT9q67
5R+wuOHUPDAn39cTBFPMzeOw5fI05HoIVR+KETvkPfg9VnauNZrqfnif9VurneqXIvA8EMBYsMRe
xJncXYl0/pl5kEVaiYKPjlyr3joNTasGVuougRpBqxkiThR4u77YaQWRbSoE7/idDsZmoDWOC1Tj
wZY767xMccESPRwmHlWG3z5swVjDaXMLrp8/y6E0VLzHy+o7UG70gdaL9Z4+p0pBB7nKjJwbURpV
eFFhrWUo6LnsfANtJG49NgNBztNR2trJ2hnKl78UGoPiFt1CbO/UBX4Df6dCDIa5IoWAfRfEgWSa
aWZTvJnppRw3jzSki/9cF32SKhJj75PRsqdSEZDFJtZkdvtzAjTU88cPzcjPUokbwD4OKBFfZcJj
722NzjEsv8rYrN7GAWS+jhPVUOlpEYzMvACAnx9WeGM56OMkQuzJ3gSh7gt15y/6cDojieibiuQH
YD3D4r+hg5322QACs+uL5O+dPXs5FJ/xidl0zgUqisIJ7A3BP3L1tYQ7JQQoHbZzQnsnJvWIB2WT
OubFqV6KBcFLgedQcT8hB0mwsGbQ6r1DsZR0I8sd0r9FC6oHXjiz0wKceosbZ/fHcfkpp4ev5Wrt
3QESZbSa90/bSrGp/oftTrxJ7rOusOYMv1tm2S71YVginQZnssEI28RUIUD6C+Rsxik2p2KgDHVq
D1AIjR97wUX85hDMh9UGX6SI82XOsofIKdqPo3JpVwoYsEs6E6ONAmS8BFEkqIJMwQwMLVKQbUiU
ogaPZ3+u2VSuIeftcXoyZBUpGX4StwohYMgW7wJ/ntGIU9e42pn0qymH8B+1JX2tcZ+B7GQYieAa
Hx5CRlLSAcDjszBkmUVRH/Ztj9HBQgW5ckWjxZ9BnEencgtNfVlQVkyGFegGM5idaivAjY7j58E3
eQEsGT34shweWYCWZ0v2Q45wQBtZX4erx79hYrIKfKMTPDXZT3uMnzDCuhR7lVFGgNtmxPir5B3s
n6aERIlhVdVOz8ItxnpGAR1AlxS9JhlNtBj4bMNUiNOZiQBNycjItPCj61r2RdxSTt+WM+C60jpV
SA8t7DpMqKj4PsPfg8V1AZPGnsn0AArlHO8HYmjFfVCVxmrlyvCURRi1+6rwLJenkk6VYz15FNF/
9QMEmbxdDn/lVwcu6IbDQen7ohx1VS6EOGWta0oAFgCXRW7SKYYxETTHapxZ04oP1OLmdRHG5m76
nycXhzCRBuxQeeHJgfBNPL2NPwOLOMWR+56oAIyBlFAiQ+YkChuUdMmD0noAbsvy/bj/72YxMgWh
YfyytD+3/oKC2XpgAIWSQDDwbHGaEpfVnFGJRzGcMWlwv7+S7frjuenQiWO/jTROj05iLNfLtifl
SvpbILSpXJaqlIZCcGlzEFJvMDIEhkRemUGNFw3FQVhB8mnyyfNiSMnxlcZYA4wa0XIyrkpMjLHy
DyAXyA22kpwnUK/0+9aFhd/yq53Th0OQkrTVnHe+YobI/SI+hcPlxT/EmVEL8bjboL2FSJhJBNj9
75qhqmK1QFi93smz9nLtY1e3is0YQqMxb5aSpA+MZ/VrxTVNu9p7eCfXdq63GFcZ0hl0JOryZrA3
EN6xk8wWkArPbXgjgAjaCVuAJpnUbxT1pU8P9xx+PsUUOUACdyUpVElUGTd7a4zSN68VD/ZmL3wE
Vkel8EEf24CInxmmue3skhla2G51yDSbs1C5hqN5aC3kK1QXm2IE9rh0TmAlOLNCFKYPTRNQR6Ky
Yfa621YXnLnNlpKbLeGVOGiDsWIAmBU0SiG3+VyRPVFjo0OAK4eOiAew6GW1Em4apEg9T/20hW57
MkaBzPUpaWxRcAFY+SxUcrO+5dTvy+6BX9OorKOOp55kAYD2/IxZSTbbqoodLWXrvDD1dNnubGuF
Jpbgz6/G2yIrXKrWl43738XrFpxr/WBI9dS8ocYOoCx1m8DLk8a69QRzPuWXhg1ux/qaPjB3JegN
NgpKVG97An96wx/yr686FctZwlO/tS/90anSxxwQaMVy2YPlarEjAQtogxOREVidO/iV7Ww1ySgl
cZbSRYegmN6M7mXfGDPX0NQL/7qDU0G1lQc7Nwaz3mkp8TanIiLbWk7zzJgNZ5mqFVBpJdO0ec3g
xCkA6h1G/GPZ0BOqkqj6pNc7y5ZWe7e9YjMA5KLk2V7syeUjyx78gWRHOPbhI59ugEL9HA2VkRaG
tYPxkNdEvF4SBlipG3pz/OVfExva7unE85w5s73kWnFuwFknCXn3DNeXF8mZJwLZrpqnWpF1OrZ0
+0N/zEQmshxl630oBV5pTAF5klX2U8f70aw2Vxjl3MTdnIJN6OcRMO5xhPfmd2581okuHkR32vp2
zL3znRNlcolW+ily+p2p2KXl/2ABdlpUdqbB8yLSRgtaVzIlVCLkTDpp1TGfvsw2eWOw2ipeebAf
l4zRS5CQmcQGfKjjfdsH3hzIKkxJNSzZzechcdjGIRSgJPWyhDw06RgswtjiwP72bvItC+lJmmNO
sXsouHbDsvnxOlbnlNXeOu34VByrrBqdh40hrjTTuW3+P+OV8z6jntNCyuSmAy/g+8w+HBSwDLWU
k6/iNA4fd2DZJ6GUQlmNyDDbdVpUsd/pAoSM3kIw66E2bwWPwoDWE5qBDIeWhxurK1J4/lgvP4eO
oUZRNGz5wVPKLWpAOdJ4SeVLn8oEmql9dclzpT9HQOg6kWjHn39nZPuT2CTQYeARP0ki2ha+f+7c
0YX2mSceMhu22ZhAL7X/c7nIMWjWRximO2fRaIIL3SctMoRAaVKkOh5Fgi3P+upDFTq5p/S6IJ/t
BKjzHjLzI3YDXzNt4046WlenZReu3MuGHYl2emMBSOq/pUJR047hcHyYenWfuW6P547IfSSXWPf7
VUs55gAPC2gA3M7B8Wy/VaV0/r208DMpe2/2dRi1YjRstJQQkvqmrtokKAiFRK5X2S+loz6ptpeF
0RmVZJfucslj1Nn8LSIDCRoCOS+CF23AKqG5Oh1UjLw35o5BUFVTG3UTEGgCRU1aKQQsdDCDMnn1
6aVDuVe604AbECqoO6JTeqQCMgWg7RAh2TP9+TTzBp5D4r4R3U3u/pmw5xKYqLgvMj0gdQLNKCio
3zZ6jV3weyCwvhYhokYuK4iUK56kOycTLFwquDfs4mCv/MLiDRiORc0bw0w4ScZPzmLFulxElYYA
Q/tKJ2+CTtmoWh9senUOSjjJR578fxPVfzDIA309i1nlqbaw/NDMCcAsp1yXIHWBWyI8mHrbHynI
zpS57tPyNAKEgGHMkAcLKa7xsFEgNiPkMCxSzoKj50hCY3zQKASfl8b3VDqrGAX6Pi25kb5krGFm
jBGWtXpN1LD7XC+Rx8yN1bGmXHkf6C+ZPRHLtv4BOEyBL5y2fvS64lrKDvIm1bthGbXQF+zj8m2q
vj9BIBhCunUcVtJid//taBjcXDGu3s6K/inI3DPm3vqqj51o0UNbAxkD5iEOdNV/NwPQnhE7QEfN
4Y7IsO1fIiyNkG4CXnBgn6D2C6mhOTbx56QmUw/oJhW8BkWjro/HsSG5pguL9HdlBPv27e3V0GjP
teB0+aNGgSBurUgG4WEym0wxh5S1Dl5c4eEuOs0FZ4nTcPTgREQLqykXajxFaOjrlaAOm1avA+9c
c0hzGBMqa/lZbHLE2a9M83CJD91mqFiJztI32sr+cUDQghJio/vxDUTWzc21rdv2KxQJ6pXhYfcv
qliOERitd8uQswp+nj1uiYVZDS3HSfKI4XsO1NHrk9bpybBrAC4rYAFrwP3cWlp+gKeFyz5RkIkI
wOrryME0oVk7wP6WhIqWOjY5By8hswHn14caeqHLZs9Fh+fiHW8ApiPRF2iXwzjQ8cHZX96XRva8
zn1fE9a1qW0NpOhAy23zXUL12zWZELNCXGNIxCCIlQwvNPJB0EefffeySYkBzhe3LGJKWRvkKTcy
kJ/+vOxBgglhXRJftXjgvsx2AVLByCC/IHe26TpIi1p2LdvsFdqcJG3ZbOyG/Mp9nnKXuxo4DpMF
5nVxaP4OVXr9eJSIMAu841SucS/d3gMQ8FQpeldeP8PR2ttRLH8ZCZSxZNKuwEaRZ1Hc+dfRsdBD
zTNHQPNrJkBiktwnzxatZqEAesBLJpu3kuxxvMoPIyt30qgkA6ZbKV2ziggjL75E14dbF/noH1aF
wQ67XZyRVsgRdqV61mrsH2GcKSdGUGiRYYgduRpV0tJeaFgs9JYIWVFl58pfgsLW62SJKYj/ruM9
eeURpmSwz5NY9qA6qjW8YQfF2L7UD8Ou6BpnAeOlDL5kwK9iB2Xp2VQeqMp421uoNE3Txq8LtozC
XCrWQIITU8dula71eymb8oCU3pOtVZiiyLmXVJMRTRy9HLM1EaB75lx7Izk5KJ4kan09Q3RY7PxF
o7I2Etm6B/JHtfbtG9DPadl1Q8XoYLlzGtBs7skS4jTHjKTrslCIEUnGajkLLhjoGe9lyIY0MAu3
Pi2khUNTmAKZJmXENOAssAq1LNYYFlkBQtlmcw834Raydi3OEckKfbCM6GLpdAVCp/gTHz1TUdqn
q7nk7ZFvmkWmg/OjoHaCgW39dzQzvIvByA0rQyYo9raD2dWIg/ek3YrazDTyn6fscsgxHuDRWak+
1ktZsZbK4Nle0qaNqi5/4ZkUOWyrw8M+zO7XKMUNK79F4dy/Eb2GJinkiT8gD1hYeCpCFUWi1dtk
wXniaYY5tcuraipREttH2gvmSvAuqnBFCMsoOQA5nxnLzgs6Rux01CLa1NUM2j1b43fr+wcQC+59
AYHAxmGTlzO8cV+juYR09poa95OrpND+INxQ51N6EBFWSMlUC842+KgwvKdUKWe1YDONg7B7JxeV
vhIw6oY92ABqlcii8sqZyYl5ypK8ymb9YB+HWjw1nmZcH92RVhI4mOZ3cGMKsJNY/slAy7MOBYym
Ktq56QN8++PUIUjP0MlV5ITv4Wldl5QW1wD/r+XZDcZp0VnBEkWXJ/lKvaWddSPKGACEYIEuFpS7
hEQfIDDTtCiSsROULz2eZPRp/RHLIOEogc8EHaELQG6U/uqFvgjm4WncB6os/3D9tPZysUFneebU
qphe0T5GKs6jVGtQu/lGv4e6q9E9YB9YTYJ/P+Ti8bZ4ll1PoEQjIykf3cXjJSuHf2YRUScsnpvS
Q1HI3v+QsRXqnAeBissyoguBnEmrYLynrb1ur/3N0RUCrxTjtrR6gmjcDEdteB+zaQdL1NHI9Mjw
cV5sEwaKKN1Nh1e1BHRtge+lLLN2NizSpZ+ruC/9WAFH9fIhkpHeREu5iQAd2w6DpuDGLVay+9Kq
AHAGzU4n/sNZJ/7HPnyTQ+9wi2vYxBOkWX01WyM9DYcrAal5yLJsGBa9Df7jjowL7l3nPOkPXAz/
AEkO+d3D3JilR8uzhsfUx6Aq5L0iQymjCGu2y5rqfB7vdYH3Aqx2rb+iGrUi2wfriO9fCn1+/vTQ
ZXgMAaYRIlzi+PpxD8xmZdS/jzNMGhDDzr856lpD0vxjNZuWClSO/MeePQBDv8PH9QXdhoCHciid
hrpxCsZua/mFJHCmM+RsnlDCd0wMZADGNH/7QntsYopmsuymJoOX3wApig4qb/XO9J8kHM+XjG+E
pfLHWW4rz9Jlcjn/HGxGyMZ8bsM+lSzbd/zGg9lGtuvE3XLCuKZ+r2XV0APeXOuZec6afLgkGBYA
2QK1Z96bw9AbYX/yZTSGMraywCr6xRa8V4Gzh5VLxxWM0NWSkgi+cmH2AneUJCvxjaOckGFuCTbI
AXxQZODT7s/Uw+H7S30npSHSZv39x6uvuTeesMpkw4am4RCHvDCkw086MJ3ZsuMG9g2gScQm5yJU
5rafyU56XBtFtFiL6+qHlMtB0rBhBOkrdLXKISOh0ZmXVHPaqv5nPXnBk6cC5wgpN3id6v2SzO8b
T5PccEWypKcx/R3alXvBMMTngWPfUghPGDI88evWdQA6H8jWyDG6j2z9jcirtnL4wrGmsYwG0qgl
keKZTef6ynIq5qN12V1gMoBJLFbfPuk7FGB83fUU6ULHBc6N/e+mMs0pyyarR30Sfq6oyH/zyix3
qaF6Wo1MCgMsUgg8XR7Ndkx7eh+p3r/3dojRa00xkxpujbLi+Uu9xNg586rXsJ/LNamC6uJ16LzX
7uUVwNIAh50VC+3h1ekQuyEk3/R4yOOOM6MvDcTl0eFCAh6eRd0VpYX3kauWHyv6w+Lp3s2aQTmh
4gmn5W7lgsGwAXi8r3nahj8gSpME0UpmODyDp5lsujr8ynCOdcH3/E466gcxYW64X74a3tqW1HTa
ZfwfFjydzojqwTdnuABWsTWSsrJY7a7tYIc7F2HSm/4wFDcAVqWDTC8HbR0Drl31WzWioeW5dIa3
E+7TPwSCjzJfFVxpOkGU+y8uXgJEdgHro4go4t5MiINW5KuQG+8Fdp3JWHRcE3wBbFBWR43c7qKi
SrBeISPYPmdzCNGwsEGdrVVzJEZVIPHmXY0+EsFl9QOscIkOtHyj2OUK9B5WhDkCcqTd5CNJTS5E
gTwxBD7UkuGI5N664n9FWZPyJkVpTzQiQXWUVLiy8Th3shl/pg3NZFUED+GBTXua6noUj5wsb2kR
IBGT0H+aVYtq1pbDIepKz12beZXN8Ym8wOp7Gzr3hhPaZK21P1BcpdqO+aG0zuJb/LAQmOlyGnzC
8q3cgTv6rQewsk4i8Ble3wCWHUxZdB6If2geMwfW7WemJdhtF3XYujA/Yur7xE/vp/yenEisnhwY
AVnWgxLbtMXhLm+z7HCGSccuMOcsQ8Htl5/wvAIDEV9fgkVf8zBiKvutQEpj2GQGIRTT1iUqfiIb
XyJCH5TUJ8v2jJAimSj4ouedyfvTn5qDMLdzApB3kOJIBOFTMZZJ3YP3mNTvr73/dRxj2OCYzhCd
7c8WWuMTtjQUIs+LtkwGTcu+Zwq0fTDDBGFisep6aDs92ucyKP0HrCOr6huu25YEsyuLpLKOniDH
v0EV1hMslv9hHsP6scgsWtUuDlu6cLTY+PXZjMbQiGu8s6HO/LH7LovkOpCTv5hALLqNMO66AR50
JlTLTFmdayuj+qIyVxtd3KJAzepKOlo2DSWLhxhEirwhZohRGg/2FmJnAOdDZM+0jZn3EEsZ8VEc
jqIwQjcOKFRCIc0whoyw/L9rphcNaiMb/OhBJRNmtAnghQkm+ylB8Tv/7BBk1O7D4ZJGyCXGn6TA
ukzhpp7WVSUBAUcxoAG9nIJYPbyK+hGfuDZz44ewMeukz62m2u6ow2Ofq0+1z2x4pmhyQS8W6BTK
p8oHpB60Nw8gYF9eBbLXNIsAIPdDZ8VixgKaQItbkcieZqJS6XGODN6NxW4xnzvIcgonohl9yAQP
GKRixyKYUzBC/Y3dV+rMe9oLd+pXWLFncR1fhj0iRbGZDfuutXO8pAGuHEi8+EzQtpMX3dWKCNXS
TG5b+PSpkxQhSjRTNHaYIituMQCJqLcXScpKW0IeWO3YrIUAtOWHZLFwyYZxGJ0DtsYCGGbqT+bE
qJl8FZc1opIhmaaIQfX/m8DuWxw3JFyGGdPxOvT7GVnv665ZoqbcjKEtcEQTmjIHdUEq2mzWHOUO
pEIWXkUf8m2Xm2YqLtXwiV9ZDUEjaXSf7yzwF8GddLx3J7VXY2SN5TXQ9o7ROdGT9nR1T+Yzp9BT
WSGcrSwVl5eCemg7phUzZZjdmXbJ/fxEd7Kt8x+4gUuBAFBXM3Lk2i1RVHEEQ9Om6lJrVFGXcc5q
aYRIhmwgYq183pGGSBL/H2FhqqoN8uf7gGysJlwhm+2lUEpD9m6Ps7TA7bLwF6kgZw9m1Cj/9Agc
rOt1PMbDJ0FQuEDnDyn4gaOt/Ih0VQGpov787z5lPWjFZb1cjdM+SU7KCO0NWdtXxP91s3fe6cKr
nhPI+qUC5gkNeNxU0btXjv6aA4Z+sL/K+cP1hAlyxT3rhcmbtBFOec/umYhfCVRwGfeTaAvPS+gW
SgodwNg/PJLVPebAXFsJHcM0UKM0yi5zwMKVScfXxWn8kfBgWIye33aai66GSd75RttpFYTzifNy
1LQgmyWSb3SVPewkX2CI+L+ZNIS1CqqFi9ebVKRSW60P9YnLdFaoouYT1uFZ2aWOySIZn/CQhdpn
hGyw4Eh1CBkCVXx3tuUP4HXV8dywzddTBuPvjTyHIAb+UOhiK9WF+Qe+dNQDtkGR0ga696XeUXQd
w+SneeH1gqnjzDMuAabDIY50Kpi1pRhls8sR/qgqRTWBDzfRVADZ4YA7mF7fXFSOu+YgrQvGl/e9
dXvsLyv0/RP0rXF6KV5wIYkdMyiF4XNP5Wt/f4yidOfgAd/0W6KBQXsiYEXGV5uY19WzazLqX3H8
3amfRWZOhhPu4bVHBfFllm7lNfVFoD/Lpn/cAugMj4ztC66lkOdtcCV6+gxxexnh4fH44hT5U4xQ
NpXTWku2azEg/yPGIQIvtiPIK/WCZauyPWRSQ7jevjbSZ2RqkUoUo9YQMCBiWnvIiZ7novfudHzs
eCPfDd8pAKImxDOY0aYt/mO3yQkNXTsA5wF1cVESq61eIYvIDldpjCQ4C/3ucaEJBms1j7WJvorX
baMzEv1ZHls3jM0dmrwpyZnmnm6/3eORhqg7XQNTIg8+YogkfwoLa8dnQn+i6g3OGPeNu0+tGifp
ZGca2GCqKNs5Idnfe5q+RDJfVQB2b9LZjzoYPKcuA9g0cmdjdZEhfkGThJPH/KxQdoMHSpH9idEN
tNmDkhdQ8oN929gFaBjuHCMx/LKhm+zZAe2GMYkAxtmgeT+gP5DNH2WM4Eqna14ene5iPKTB9qQR
/0pnDS6kjQWB59t1B0gdxBVerrKzzOGXcogfYI3vwVWxAM+2YQpW0/tSUfCJ8o9HF1WD8UjXEkjM
MoT7uA809m2nRxzgndRjt39N85VznnSQGCq9kMROawZUDblten0e8edb7Pq1ltLzpyLQcdih90HA
WaK0C5Xrjl+gVkFrxhXbePyJYKh8PV9roRMia2Lk+4A1gJ6aJB/3/i/fEEwhyG620HmPpOPvahHI
jfS1B5psiPOimWE511t2No9TrBvcKWoH60T6aXCMYMVHJHvYqMigGl+q4TnAQMTaiygutj0Grz8j
u7Zi3wk4LxWmWsVNa5o2700+7ItScVPTKB4RQ5OAILzH1JcYpPpuJh4fPmfWW00PGOh2XkSkc2Jr
n69NPVcTaxF3V4fcj1vfZFF1DHUOXHELDaY7KF3Of5RX5+IgAjWWIO3iDpAjFn+RnHqNj2oxK5/6
7fi/PtV1Qzf+dvJclltjo3DnnTcFDnJQEg45znxhlNI4OUWGOzrkWLblOPE0auwqdYU5C2lhtLeW
GKGT2PiAvBRXXXQzicQtCZATGsa0d6WCGUDwI0l0vPP4NjenIuokSAd2mVsEhb/VR3Lb/KpQGtwJ
nDQ3GDG1tBapzTdzmSoQ0KURN4Q8OktHFZijFywqzLYEurfXrN0HyXoXHcn+DuujSP8tkl4iK7pD
XDC1mRaGDubuIp3nQlVaOejH+3uPVD/fMLWC+vSjDnbC154sCfL26ogxWI1fxJBxPj8JCbYD6Nl2
RX8QVGS3XnVgTPu5EcmLpR0R3EheZ1c5SHRInHqRdxi3mLaorg3Nsq9HsLBiRIXcgIOby+WfM6ue
pJHTVvFydaTbAspUrDlYDWtrqEs5zVrLwZpEDf2k7MTZyYW2mvFrG9cfRKCp707r+e+px6Td27KB
v01ifMqATOuz4rE7vK9uBmtw48JGEZe2Xr6yTw7veY4vGIL5JCUoFY/emcUXGiXm7NVL/U1Wxs00
eBgKoreYCKudbnJsSX2z9HL3Ur5hGWEuH+lBnfBxUYHQiv2T2jGwggHPi7RdCpCYXf2hZgIenXKq
9RMI2UCZ7svYUu9O4tSG6mFV4JqhY/T7QmR2FGaE6WRRKEJrI07FIhrKI6kdf0GtBmtmWIBdUblS
pJIeySBVyV3URJKDImFwopxn7J/J24mGD1dH2H28xoJUTkiuCEAgB8oDg3YndDfgGZanjc4tgWJV
8EPzlIpNQgDblTypG9yRlaUm4ioxq83NwM+oVW3IbhWhNDLtcTlmNjntTZzNbjPUVQlnuYguZQWv
obScrNTx+4k9IMIgy9k4ACuzDHWUuIEwqEfxHlB7ro7GeLb1SK0easriubyx3cKwfE5LrxEleLJr
GB7squxS1xmOvKFJVAZMiayIv/lanRpUdl/XWe/jn/gY3zmNSvV7/+iS1lNLXu3qdDrrbtee4odD
RP+v0gJsuo3f+brDOO0C5bVACfbwO3QIHEeonzMXuaAxbI8FXmylbRtImJxCI37njU7ur1mDUIwu
WQbu9kQVlUC6kLuNMscOxsSWzFKDhQfqEc8KAUR6I8mJvruS2vP5NU9o5hlfsaT5ePTZ8OInfV5v
S9If8LGBZh4zmIPiHQVedfurb7ee1pgcGNDSs21Y2pbtr8Sd/iyK8aNwtAtF84bdAzZ+R6PZIjMo
zeEYmzldL8vEf0AeeWKzU+R+dM7jfLFdwTIqCElh1imI1MOERllBSKnCqUSaZENp2Md/EWU3AlAU
dL1Oecxkz403cxD+79ZgLb71AdrQJcUo1EV/ZUagFNRWLjFNDuB9UAqUDwBG2I4OV2oHqA2QOO+B
uMXNoBcDEFCmqAxaFy8Iwyz0YisR7jANTSvmjz2WlfOFvWXCKPqrnP93hCZoQ59HrvF5aPpmFNOF
63mviD1OTSzo9cKy8I0WJgSTZcZ3bPwFb/Qt17N5QmSqt2t6r01B1vxhhu+0d7hT9rTczQQwO+h1
Twh0vGZbOo4jtxjQcx/the1Q9xY8yYYqDaliYcJJMiRIK6EN7MqY0y8Ty3pb/WdZFDaZYBtO5F8u
B4LInM2KLYuweNfjwfQ8vLSoIFet8A81sFX3F0fOhqFTRQuQEJJs5V9O4bGVAbEgB3kENPj7+T4y
vG2OEUmQppknKdF+MLO+sVRm/dOLJZZu2VVtlJfSpOE7RQ6bet3Fo83CGQKlh99T3O2tN5mGAxgJ
SL49lDb2Hf8cE80VCdr3ClwdFh4zAapKtcMoGfWiAKzjYBj3JQFneQ//0eSh5Vnfj8t7f+vq2a+3
zDzBmHTLQCWJ8ulOsuvmEg+9kd/h7HIPI/fvo+glzyM11Hil+y4TUc6QkHlt9wuw96yx3B0UeLfZ
GcZ1w/A950WztEAarxl7kLeKjy3sbMvrrHa7QIVhAAGMTy3Y4jpEtv+lndv/eNcIkdKb11seaFIr
J1dz0SC6S2SCgMNZgjAo3mYnwnJ0Vou1+EiQnZxRvGUtlkB2Ndq4UERv7ZbY3heIoa8wO1CiKJTs
Rq9Cc8ojeFE4dgEP8+koUYcqjFkqo97DXkIbzFWhcV6V4SsgsoSyXpZWZnj+RBvVgwqdzkGsb2zJ
Cqn6Koade2UhJGEXbDBaSRG7IPqYOCcurOM9NQ652bZCxvewx6pEHbHP0t0ybqNNhLP0r6isrszr
29Msa3xseismTTzDBkBPvkhwDRKAsbIZIHUb3SATOxsqzPhhV5/hqZ5RmdsKJZ21AEMTnbhwV7El
YjvofDNxVFB5cE88e0P/a1Kz59G2uuFmQA27wkr2j6e2yeyWkMZjZoEzjcLL855OcNsb7xueA47l
ymOefjqruVX2kfMaOsd3+9+ykVcpnAgM67WxJJ96MLcnC+Yql+wkWS7XOKU2OXDmZRTB6kxZNXAg
DeS6e/4Uy1Ox4fVKCseYcxxYFzsLeGnpcULds05lhW3y+NAMZkut5mliEKDy9uLESJDDuCLqBTtI
wHkOz4RHBW8Hs0rlijCxKl3nKbV7kY/q9MiIMOMqlyzUi/dmbcLvAApl7I9BLvcIKnSDWRa3D4wk
+9dDMXY4ipJKyN9warEQwjB49ugOMZC+PEjRBWAQJvvljuIs+Zyl+up8tUCMQqVcqVN/D+U39q2j
0AWUCGxq/JgIxRmqnA3fw3NIah4rwllcaX6cm4sdfvsg6h8sHZ1DquznOt0IcIAjVENETbPc4t/+
IL6DwEGyFuDmGD6Ih92EUuNAWGH3KPogaTEnF5TTIp6j1419vHSmEIegWVuFJeT+Iud6aWBNhmYm
hLTQmFVxNQtXF07s+PBYm1wlzxfP2UH50Zil01G0pgAxtQBqq17ebet+z8oIPifxAeH7/wK/jIPA
GPTQcFipIMgwOac1vPE/XYNGmZuIg5NSYm1MxQOVRE9OEU/aBNcSQQ5B6f6r/7bTgknTaSpjzI6P
F9oidHzyvtALxLcCD2IvGOybEtjX6R0kz/CO1F5S8A+5Jztbanzc15ez8vjuTSv48jKumRm0H5Hi
aklKDTB+I1n7VlYWKxrmak/X8178Y5Vangq9rzqYiqoGQKSLRDtOHJatpkCGPjFj8zqZhfYLoYFL
5eXrZquEUEyFSQz1TFwJD7khmqENDVSGg1YlRBq1/fFEk6jguhvL4ibYLoP99ZtE+lh8KR1/XzDe
ypDw43wARU5qPNExEO/LKLnqYpuhKMABR3vOiAk9lKio7QMwX8irAudgMH13QwTtLfJ3uQ1KUseC
flSrDqVxFAb/9WUNKR9zFY7C3mfbV6kXoY5vwlPVPRWkjLGedxWNGfEKs+gbPFsswnlZdyitluHQ
mKa7GyDvBa/y1/tuUjwaUuqkKi5GQRjcJdS2M6Ay6ojw2mFiGLCohSpD2he7V/KtYFa8MoyKojzG
lBnRK0tgFQfurPc1UTZAUR3thk5nx/7JUfi9/6rkYYEGGupMf+hfTdYSwXY0YEjgoKAyQA7kLRi3
fnqJZdD9yMLVsDjv4Q7nEcGyqEe2y9DLMSmMvHicEVEXNI8UoU95blWEcbEkvJTUHDRYhumVlDTC
n/clGoVjlLASvikPPXLYShK/ohnR5PdbAf7+gnorCru9KdEurbThTKu1+MIMf4g2b8QQsoclBcAN
9n7x8xkeko3j3ZMej5NIPBZOv9A93foZL1W5pre5zltBsNh6UMceteFssRxoMa5AFehs0lsLMtJy
NoHO0XoowE6G47V525zuxF0Jh1aaxf60gpoR9DYbbti6cKgvRsCjSxuViN7q1Xvq6nh4oKgXXTnE
5f/9X5sVkP6sWYuArN4c8pY2pNhuV2yDBcvMYY+2NkV+omWRVRcZw8QjluF5gEvRG9F+TsCxR2f1
2p840IneYX0seq2C+pqMabhkzM3Va6n7opcl3Yb8xyARaZkZNATz1o/EirVakfIKvAgEKXGcLMis
yFE++UAbxp0ApdGMUl/iXGfGJkotA6FZkpzmh4owSoxfzfDsaAvYSKErAYKQDoyW/5d5MJPGhk29
vfhI6IQVaLoPGsqvGrhFlo90s0rxNLRlgFGblpLqRwzWQ6fw2GxMjKyqSxh/yd3pgpkDMTxYnMPR
542LFSl6RTRrB/DSNOBOgiUvtW/7NhtHJ1Q/F0YygJAaa8oxNi2yoV7wDOiIT4wEIbNreQedORrm
ebUfMLaFwX0OB2TWzUJRBNWdBvtaehGxzU2fwO7ShDtyCKsNvxOuVa2CGkEEOBA3VZvm9xucZe20
aoRkjmvAub0ezt7gHjTjHdArJvJNy59/k8Xi2gkTGBxPkIoqsVIx5aAbGVXR1pcNLitw3IKfPBNO
QAQGRt3WzbmsnvpQ5QuXO3ylNEXlS1J7bi3DduTc+Omsb7ZoUtujaDS+AUc6DohbYNAZVnuVGWhn
GczYdLUkctty04ruNGDAdz/w7syOVVXrC6tP1Q4Xn2F3H9jD8eWtuWLXz4xf2ZVfy3auLL7ptcFR
YGeflwb8KzLRQ7FshtzNVMsMdlPXFJ28CZTU4TYowVmQfNfQWG+jAeR0P17sFjyte2MHI0CpclCv
p+09VFm2UCTralZYpzWI6FCIni2+1/s9gQ0zoeepwquxRWLMhJez2p+3DYCWtXOZsB+DYQN/fNkZ
XVResVYnM2kiiShFDTwUHsYRkpA0tefz3iEdmCB8BTdgoL0zssxTrDBevLppnC8c3RpVICmTaCDv
1ackw/BTBMYYUSuJ4JTqZVvfGcha/xbwDAbEWDe3Spx62QcfUARmImEJ8ghJt6jX1TbXOy2HVM5C
6EphZy/kBxzhjLsg8jUYWUFiOxjPJFiOcE1Q3pZGhFTtxrAET6MgsXCotQBG11SWO8r8oxo2WK2r
cghdm2UZaOzqZAsZMaKxF8JdfzthD9dJoRm0prFgMmryzERpngNqJ+IOzAKTrWFeBm87Tw8zJ8a0
nLFaE5JiZbX5goeUqz0nZGnEcbCMenJunoPxYxumu4plixFG4JbYRd5IlRc/jnzulnU85/GlB7r3
3mvohxN2llxYmSaw2e4j0zQGSvQfKeYA9dhVlhKTUhBO4MOtT3sWFTQpdrVrG9MJym52DHBOnPfb
JIpRnIGITNDFtrZ7uYtSBwk/2qi1T/DJJTkPIITR2RoG3QPqeMN2qUwZSptnriHz5GUQE32XJIiF
0DqNaga74F8ihNMSrzUMmj/9D0fjyzWdfjYpIrIhhdqKFAVHpcFizrDf/rhbwtMGb3vylS9bBtdL
54gIxdVo89eZcRKGRLuVh9cgPWY5gXnwpHqNTAE2DqrvQOGA7UtFtU8pCpzZ/85wGH9nG6UWBhsj
khCbBqME2NDVMGDwRKL7xuaS3ccgqQLd7w3+rGvnbwJK1qRmYf198YhOLzdIH3CQupKYULMItUEw
I8gH8buytfY5UjNrR0RyE/zA9xo7fL9wR5EoKydjkjePpDRk5lQSU120sPRBiRXen6N/DFCFnaSE
+HSCR91KLyOLzEQK9ceI1WJ0IOFo8eVkyBXyQFnUqMWJG155ZhjYpdGnytGyC7o3f+iQ6EElPbl4
KMtOPjVYmfdyfiy9x3NyqneJgDwBD4XsWmSXo+8Ao2kJvYwKMg/baKkKHXAL9Ck2O5Tt/L3WE1kk
lGNdSuEy92iepuWKqL/pbQVCZSigjW/yRozhoXasD1qoFgPXrqxDlMTwH5Xn3qU3EPL2Tp3GxPAb
yRHk8LRZC5BsDOWqqNvZ/AxfqOEBwwqJBXi13n/82Y4TR4hvjPTXX1aglmq1BE3/EIZCEY6Ljsiw
2c3k21P7IXMwiNmLscbLgqXy84A7c2CWhS0nTb9BiRf4sIvvdbtm9xMqDqhuZSMnM9b4ZL9OTb0Z
a63FOLb7Swg9aSKT4Ymvv1YV2mUlt7z8Zw6GT4Yn/O2CNU9+n9/KQ5gQsxVQ2d2Vdyp7pjRsvyEF
jhiOFM8vReysvoBnA64DSf4OvYvpuvw4iHWhqSmPPPQfjYAiVMvdzZjQKatE0rLT6OGT/dUew9ea
E7LIDFyPRTqG6jrQx37L3X9HpfYIz8pTYFN+1WCisgJBTqxiUa1sYBYR7ZH8JCDCp0ux2GvUUTWI
EPByw+tmNYsQfDhpc18UPo95q1bd12mRHOkRBUr7FKq0dMwgh1Yzl/ti8lgp3Os2I3/fmyUhzb22
P1dfDYTdTdstrM/x/cZYuJNazkmUgXD2KsrcemHLicOc+KFpz64sHy36J8a5p0k5Tb33LbI1cSNM
wc3snzC1HtBYyAhF7o0eX5z2VydfKt4ThWvHP/W943BdgxECsv2crcp0YXOi8MYUrTXLnwGhRhdC
D5U9y64KtBu0quC0RrZMON+2e6WsHFAwAXALeukTZYOgF0sAuT2v9pGAUIqhu3t8RhylX9At8ItW
19dagio7F4hidbYAmumLRJ4mVD/qrealMHHuBcDouiRjPHrWFTb3nK934KvkK3rOAttKXb/hON7Y
MdZjzn9ZJwmfDhz1h+EIKZ01ZgjKeWiWThfobgJOSgnzD1HkKfs8EZWlFVh2lXkgCQAjRH75EUq+
fU9iL9rvzDrFG8pINwLJl99YaXqEU0M9qUCMCErKXFPXoyTOrTqWf6ASc9LS5J06IuiIrC3MTIJC
XHoBccFHTKMW351T786vkIiGl3pwiF0OxZ/g2/7OAs9K0qV2GZxG4sm73z1DoXD2aSL00WvZkl8l
rODQ5u80HTx7rOpAgagKN4ZQgc5AnLs9Ln2eoZSIZVe1iYTCw0M4/Q683wPLvKXRkWrTGcfWzhTP
b/bE4DpAANfa2a4wytKR6qDe0DqLIrlpyvz0RcSvvgSzrmU9QC6/IqryvwbDiS/2KCle2ZY3DG/O
ujcFAKrYyUEPoiGchzfEnvfcCk5d5vDuW1pPiiA9GweBIZXUmf/HsjCmdX3M2WRkx+cVy059RmK8
y4qm+gP7JUPqRi+qZ40BrC/SNVhAWgEXd3c+WpKdtvuAWP7MnwrWG5buaqi2xuqscIS18B/pG+Xl
VArARwiMur/5q9OiobXqnNRKdUGTa+QUjKyRdVSQ1YigtysMApkNmmtp/Ob9ncpq9uYkSMh1Qqe1
prtHS4zr7uLHpGehPXglNPnGFHqRmWeXXXbOl49HQLnJKh0XUKeTLuxD2gpTX7kcR5ZV41/qaRoc
kfbPIbzhsiwG2qhDd/Dwnl/7jb+siISzdGzHhSQQh/VeYXWfXkPt7Tte64XZm6H4UOyMgAPptMnJ
ccAp37FQtvCfb0h/5M5BG+MgeUmwBXVXIWuXa+YbxZmcXf0w+H30VbgH2tGj7x1wmnb3h23fMJGM
MlQ7mKBCXKMD2ANxgmP6ZI92ES/gHz3/zQHXa+2cEU3J1DEW5zMwFb9Ibl75UupJqVIMNzscPLKR
j5+FxEByW8/8epaJNoIvlKtcBk6loWYMHKps8v8XyUsWG6+JAyhECkwLuc24W4beRdCxVF9FKb+g
HpPgSYgn8z6l8ogbCVEzJ9c2JQVKbiqqvC3elHLZuAIJsa5CDIb/c1P9oOvt8WtK1351M6yNz/mO
MtyKOF/t+w4mvkAeqkiK8rqdyC66jd3Zq0wox16mnJq1UPeF7geAPWgKaQfi8XW0Dl/jXy7iwR1w
0dF1zSWopijOf3Ogw+g2ZkyCEuzltsFYSm0kyL3GDEWi1xux9+msZcUXS12WPQ/gv8Al5Mkbcjt2
SrZ0JoUhEDUUftPnIdGfSb1R/uD+TGS8lTv/5ksTgjTXf8W5vMSrA5EECGq7uCIf12UKguHNFQrO
9PA2v6PCcZMManIE/c56jcnoQTZASCa4lv7b+omEFWDWdnv/0hKMll13WLIVAw2quqwkRQMUWkYW
JQ0vz4N/P/ysjccLDoGVv47hW0zylMEfRtR4Py3nfkrBziM+uqZ7uMrufs1lyKx+LnlD//Ozl751
B1P9s6RFX3K2Jf8Q90h0yeO2D9XBw8vxjffbnOlM2Wb0+weWns4uuAMp0a+3ITStA9ChHwmPwrEv
kr/8bfViJBWXcRGUtt6rLo3gNkCpLqZyg/yd1I0sCw7esn1wTAp4DO7Eol/yk6e/h3D5TS5ZEipB
dKg1xlE2gEOSn8TW6FcATY4Eiu+po4C4J/lI7b9XezhMaJ43scidvzqS91ArnKwskUvLi7ZB8Wha
oklDP7jSkCtHBsIG+PbFPlvTEyaiJ2U1H5zqJRs3gtU5ED1JYxL/pt6ac3m6FlSnmDoGsVPX8FDf
r+itzKEWCnjKm2PN9p0l7K+WrutJ5HNUMVcHj93NAwgP7GeHbUswXZp8YbVSkKEQqj6Ksc8USVfO
kjcfTFt7BlBjaJLXaCNpXjRL3hkzR/LV9QaimAfkNyu7nq+r2whXW3f9mb5UhKx1bwzWvB5pxt8z
XWr7/VTylvFfaXycpExHaCsNpeH4nkVnN+SziVd1L1XdzLBskSQ9FQIX5DfbhC5VwzsuiSCjed7z
kqsjOAwjdnB9hALORa5XYUwaoj1lmrTJ+ym+2ffTazIbx1UjcB6zL3NFBdZTvi7EAmlo6AFEMyTJ
xntwHJrpEgMBh2R8g807yXgrLYPEoDLD2JIfl5NLuIO2Iq0W0Qcwb3N9xAm5tdINJZ1iqpzhiDr7
u/8fqGTAXOGDN2BtJxHc4u03E1D7yi+ZdYdkrTYMojowlNHTUJh51UfkTUfKbsNKaDaq6uhyMFfj
ak2G5reATASqi7eC63REhjSmZtD+kGJwDJVmWK2TXX+d6E6U+Us74BPdY20FXr4hHYl0Xdz6sOzj
6cwpCXymsjjx/a2DvooOMCLi9vKXvZsorzAnwOCTPa0A36+frcXAsE2xcciBQy6ZFzuQcdir809u
TL9yGPcTdrfAgncSbwxnyIQVjMC4ivIvuN9zrCE/pl32wVtqVFgySUqzAS5vbL/NWr6oTgxsKnWT
06ADGIKQyqMzMYhbz6Cg51TqZKwu7AV2+nKJEjLOsxAPg5yUHIZw3xttNxog6cTz339gIh1AmjHL
Lnn5AjRDVuNY2KFFYYGcKTVis6rvdm0SLZS2m+eHq0rs4JKBPA1md2Ypa9ptmdKO4RyX3WEwFK5l
8z1Xk2smmbOMzOo0hc29gn2GFXnsmu0QSr0bOo3q9vORxO8463p6pycWgB7k3tSnxyC2zIMv1Us7
kbyjXMtf0RJ3/Zws37ODujEr6u5ONJQ/R7QujNHchkBQXzpB6bnfR68nGKPAA5VNPfqkv1ZSK5Qx
Tv4+D+GcJn7xUybDRZvqqiAaiPZFibkWsWQIPDSbcFA3IDhXssfNzo+NRuJPVTEnH9+JxcjDtvkh
rd/YYw1PRlFpA54TVdCY0sad46iEbqCv63P86FxyOldK/aol5w5oWMvqsdGcloJVrOEqcLFMf///
peOn11oQBjN5fvN/cJzETqUO0SAslmAL89aGyuXIaQYt1tjK2GNTMIFRrwyoHxaG9qYh4HFvWHBN
R6byZO7ZyY9FQAbrnuHoZsgpQY/1XLVQNV1kDxkT94OBeTX3Nlj8EYD4PSY697BbHn3xb0k5qFxP
8Y8Ua48tHO+ZPxvJJhmjwpUwZksNDmlgTnvMNureUYI1TWQhBlbN2J5l0Ujcy+OJn4h4st2GbbRJ
BEqCYf47Ob9LaY8r01bq3Gme14jVmA8Y8O/7Ugd35er3yWKd3tS8wC8eEhmWcaaPhz70ayT6qODp
j29BHDBnKd5NYdR7xrK36iE2W87WsJqQHsMj/gjpatE/yw4Dy1r2OU7w19gBAY3x5ZlM2HsG5PQO
dCBmw3Wm8k3O3iXLbiHWVnTwNcHO7o97Ai73ercpDiMdSPy8Yjk8TmydedT7v58uufKdczEbxdhD
oND2ptz6YVo1Xo894BxyB2uvGxDKM1Ywojr5LuQjX/SywgTAYMc3n9jqK9DM4uaRlhmO6IicKRQN
mvrLnNNuSUvLlN1IkG6Sf67iRvVWl+KzmekatgzN/jczQE0qO+KL1My92oqEsieY9kah4Dr69cnf
lMjk+mCZ2XcFaVNCijoaCmB/qOc1qqeHIQEmT4S7jYKa/+8DUtYztbezRvdVG35AnhxKuquYSUwW
UADhAYWLJny0uovR2NHD82QGPujQgYuMDfg4MUkMRNeP7/4PnsI6PQ/Q+fI/38UP28M3WzCx1A3Y
v/v+Aeek2NF0yyhtH5aL1oh1ZFW4kvHEtXDcjpQkwAVlGPUkKjGvfAndKsjDhkeNG5INFSuG7ohX
tUomEgkPJNBVx/o10tVkIQRr3xUgaYIUbxqvy+isBk+kSTHqsTazz1PaBWTEZ0I8O09mQjzi4c+i
itqybq9zc88Nfe1ql6TtB/uclo7l6GQ/AwioD/YH67vOtoWZRZNr9Wl8qfC9XGUzhnolXEHSdKWY
/wdHYUIl6UKwyKKIxe5P0G4mX/Fehf113HmVBFnFpyEamlCPZWcL5Sens8PkbPLy7D162zdnASnj
QvULdxTs1D/68bWiQHACbCw39gRmEaz3od3s6glNILVbCQSeTH73LhIh7I7zn7GK2/N+aBIvXOir
6Kz2A9ZeEU2Yog2WlZj+kzOXKMAs54oVOC+wnQ6cQ/U94FWKTc6guDTzY0mn08Cv9PS4cZMTFbr4
mWMEtneI1FZy2Lycw8Gw2rtnfFmrBxyzCbgFXlwXdYy4otRT9a4zllS9oWzb9DpehDmGhzbobWJm
7Xbs/Ff7OWEKTH1f5PJBjWlD80zfyJeMCAppbMa+TVHKa52nLVxg2trCemKtkSApI1jocNGu1m25
Hq11bIGju2WZChZdscXQfRohKy1Cn7DCPb+y2nB5ChE48Nn7Tm+nUj8kaXc12evEgcYy5qu8L4dW
8bN/UD+DDh+YDLqlA6gXlmuGFK5XHeMWTAxiv+AW9q68GKsPibQkKP923vfW5krALfcMc7rCEVMi
SDnBcMR9/SwSrVKCwfZOZclp+eBw/K38NUFZlgTiHBfvzlsHUT695XN1AYJsxubjvdPynModecFP
R5KE1MoOsRiGc7CEaPNLJnSljXf9xD4AqEFXZqvVAFEGd8zeLD2rl5k78oTH8YFZbBkPwy+1EPzi
6r4EqtFteRGdzFurmnuhJ8Zt56zbQg9AMK7Z70YHpHeoX5IuS432hJO6Z7ZpGoLUTCeIE/8Dwu9P
HS4+kY+Nj97H7xsfzAboOXK7/0gKK3byRCEqBIp9TFlCd7ZsY65Uzghtcr7JSM4MY5HNEdfNbQmn
XWUBACMY1bfborGfvMjxATerm3ZURkT0DjwygRSe8sgnFVmusOiBTV30ggSmP3npcX6pTlDEDE/e
gdkWSwqb93XQK+5d0BhSz5pYUHl7WBDk169vNkMZXhhEyCDLH18BdSNjWAIqQunUdPXtnYjcEVJ8
oAe6z2IGnkyf/gr+DS05ZpUHXOiaQ5Qyg9LidzMFVIIhuffoYYeXTYzhsJctTvnY+ubMs8aNQERT
pyPCowuDZzvxuRkMMbpFfmcNtUig04Y5F2rGzMdhN45bV8McpcMiZFglz32YYBxKDbDkzZzixn4+
YOD5qit0nQzpVd+GfLirOgoQ/LU5g5GKH+6teOKTLdCm1XjJj1a+/SMCoWJShTma/0KEE8i6JspZ
fELz2vokCqmlDkoLYrqTy3bELGl1uv2ravldo5IswYhbHgQ/8SthcKrDd9h9Dmr3vp1VNl4sVomq
E5NQ05xb9ZVm7Df9eab6sP4kMLVcwZKJ+Ijq2qlfWMERVR75CrCzYKUUzpkwXTiiTG+406hpazCn
NFphY7cvLEvijFdKtPqA4kWnXJ4O3J3jYVtcYtFfLARIRq1LIac506PC/GBKXAVfHy6i7upjhVT/
S39LTJQuW6kwonXu+pnsr320d53rdddXySG/ukErN/lPBiSY4lMBvl4cAu92KorFMnAcl4zLR2BY
DbFRPwgaGRAV6THHvtMGuXpbD/TYy0ZW2UeMrENmSqo01Plw8V6RIs5iMazzZBsGQiCuTt60JcBy
cj+7Gw5Yz9BvtX0V+pdkiRlDLP6DabeHY0ZXefhY3Li5He5I3oj2Rp8tuZAboAWutf5b6wuYhQ6a
TJsTx0yzj4RdKkNe9islNErtKp2Lr0hpVPdwuPoAhPt3oe9YpZW3xokc9jluTO18ximGXSStrsyg
1OnXxfy7xKkTxo0n6h4pfmVhbw+rh57KjV5LMyfAucRN96oNVtLw+cl2m46KfNgg3i8c1QspczkP
Tgs+ty6IWVXbH9wOTj/qpwc2wPAJWeaaDzW78IM5sA75c9TjQyjwAsXYI94te9GQoAoD8PFhIn64
zVFEuatjV615kIXGcBXJhYVcchWzl6dOguW1tIh/mHPbsTjlkUOQFIuY9xj2YO4AYCjyRz8yHPcP
EVq9pXKeeKZHFkggfKvodHjMmdeByAItKB8QZBHziJwDJRMcLhHoZfsMnGpZMInRmg4ACtxrPggq
U+oSov9Q9zCwFcMqt7LIYN2jniiUoVDjcFWgf0QnMF3DZyt+6ZXrskRKu+ayjmLhFpMYjPluMkpc
dAp+5SJbrs/f4KK0L1j+EoRXib3CAzMAP4shuCJryoO7fqDTuuDB0eteN2h2Eo3GWmLwY/Y9YdNG
E6en78km6Spo6hd/P0K9h+4Ex+wqx1J+eZfUYaxhuLrgo9BtzHtJKwah+Pn3NKu1qW23rsHpEINC
c2S5YWMLo2dj+en7M3wyv+CDQ07Nf7L70IFPnfCq8I+kVGxxFVFnKjQh7CV0/qaZQKdeSnVQxLfT
/0IPUHxVU6adCqv2HCNTmk52niSX+NRrrmm4M0tP0Bj30fXND86ciuAC2zqHhcGV7L8DQO6vzds9
lbvRj+MBqcKIesLwamian0hw57Nnk8kRCCOqZdZ02ZMHt3G0hoFmWuwWEMGzTX3+gONN3F4R6iQA
aNm30SXJ8iAf7CzD0DcMsUbaT2VS+fqTwk1zI507iPaIIn1d4dgDKXLZTjMI4pDkt/azk3GhzuKv
DMjdVvRC+ELBBBnOUMgZjS1+AtB6rmVnjnVt0Nde1TPSveyXKXgRvjOcJmPvqw2b9ZhtQQM4EIdu
DNDyR6heDm+OBoaXQ+PqMeIEBm9lA6BDHbHL2LvC+vaQB3HW+u+j8U1BcrU+Nv0EMssrvQQQj8RX
sW319WBKu/A9+K3RYOQNRFrutbxC/VuLPT350f5LwR9X4D2XRXpfkeJ7Iik+HKC05LVJcdo8B5LE
paJBa0g7JNNlvoil7a5KgyDeT7vIUW9NJhgjA339F+GY+WXfl7NgRPU7KvkrzuldHh+BaFtNwKH5
FojkDgx+/aLLyQsrJcSCw8nMUzCZAL2P/m8vCazWVwLfpdjmDzUTo1xejUj58wmhZ/SbmwqqhmsO
D//1krgS8tAeEQ4ALG3ctmjU1BBrGxxHq8Gq2XZOHQP8eppfBroskdDGNx5w4YWxmyeoE4T0o4dq
TIVCFjd8VaMSxM5EPob/mWCSa/lGMCU7Bs+0P2BpLY/iCJ/XdU+WcezoQhuaBk6TchwghlEeOVCI
ywTBJzgQgHiJnRz1E70hSSHaUCJZCjUdpYCjb6z2T3B3KdJUME3iD3o9PIzXS9j6QpRHD4RxI6QA
W9uYu1s+/sGimcwUGIZV28xqpsKVQyi21U8ykxWqk0mx/yvj2/DKNRIbDSMU60NyA+WmVYi7Dod2
hxD70E0fboe49m2Ir4DuqecxpWnKrN2VVIEWTK06SyHge+a/o8x17XjgvqbS45LnbuX3B5XQgD/n
iMAN9pAy2ShTIkmmMPKprRVaygon0UQzvctz8Y8nXrKELpLG5TKh5KI4VUSobU8y0vncyxc5RCmj
BfYX4Ai8zWbrXjmBUJ63PdhzW8Ns4DwvsQBL0ZuM1Kvfcyt8kW93OHVz36F24JnZN5w7j2nebZby
7aH2zdN/l0lR44RuYuDB9cyCfK3Q/sIBNmg3Lbz4MO/wPN2LpfJSvGBpVNa548Ofd2+jZcmLCqgH
WkyZxc2KdxCV7ztRb3+fabc27UpuZMh52kQzzU3LpAat2lav0Jh0NdQ7/slPssi1us/N2/XIu0VW
DcJvdHEMwTcSS39mi13iLFGPpwanNnvBt6pMc5hQA7KCn4q2pTbkyQMPooxQbtf05r/4f1Su1K53
dEiEZHhVqLgomYjO78ItxrGwzRpmekZ9ly2AQboqwIY6H4R0Ddo5pOHXK1HyF6Vf7W2CB4ZcLNoa
nkpsVzCsUwvTVebSq1p7YevibrzjGRjkH3MUXlIXDTpSXXfdJ9HQ2w2VEvF7vcqaFsFxGVwvpu1I
DwyFDxNBgHqgxes+RwUT8RnAYfj5poC4mpZzHaYWG51dZYcj+gBu0UxRzamYarb+NHYuOq5MnCN0
kDGLjA5Rp91bC1A80pTCChn/lt+3APEkGcfAZQ6Gm3Yrt/yy6GxRYhH7miLs9JIBFiTwmG8MEKCM
6wi+SpkxqYx7i5jRP1Ck/RpY50c3K2aM22uZE+xMCc8WwdAlWR3xW4Ft+fqWMGTTUsNbcadSbOHf
Lta6skIHcx+oW1W1et70nC08GNm56V1pi3j2LZchTRpYEy/FR0CE4O7ANVdztuTwA8oWy3aUznPy
eWcDLRFndu/r9Qr2QAZAe0doZEGEZQ6/aLylRBEm4Be/eh6BvZyYESzD1i0NyuzvPKZ3zl1A90aF
4pKSS82N+SXNuqd99KnckTEYUbIREe7YFDK0RVIUjKJa0Tf+xP3oJuUfV3n3ZVG7PHYh2TKJzmsn
Lxw9uKNbHqmy8DOwrUKN4TjJNJXPmAZgUTmN7c0rnFH6KicF4Av6qMTUKlmh1DLg94Ijcen+88Uc
GciRBwafbxhZQkYMbP7/UoeQHw4SFQlPzDY/+kaZ56L9UBE5NJ9qlWevKV6Eju1leFZkiKOfVZsZ
dtYuioE1JvGdovhv43ghd007tT/hibBfYSzSvhLBnLUaG0lkRWlEc9b2AioSo++fEjLrhA+w7nHE
m/AB2HeRXJ1W3OXkz3Fo1Lh+hrnNVKSE0M84BlLONcx9/uuLoZ6pNf6L4s4mz3WsoQqWqaAxlXmJ
b+kKKq5OMCAKQgYXyRSONtS2FaQFggYvqYMcAzrl9+iZMRREyvze0slM79A4yrWTtdzAnYjaV2mA
kdCIo8Xd1RAd1BQLd1FFYP9LnUt2ALKD5HAEeR7BnX0QGLJeM5SwXbsiMw96vRj9ILCz+zhbT8M4
47+D9Y7UKzdm8AmzjQ8BQwYpOHIGgDwdBNz0Lq36lcvK9xPGQ9W2vIIfD/61siLHFAFzNWtRTz3n
nacam5dZgMcf/RDmYwkGab7SKsp+owiIvSCmpIId1MH4R7lgTg2k3PreULXOrAWzUfEd+QT+kiYA
BtK8dtbW2hvkOmusvmBcBCM9E8uH3KonQuXQ9nVf45JC3X2YJywIxVnK8Ts/eoQYl5Irb6zg0XNG
7wPb46/yhzrTfavlmqR/nG0uiPz0cFbGj53UANGW12g5mu+ixios5KQwOx3V3mcrwWurs8BJR/RC
y5iu9y9qXuK5zR3nXyv+imAfWpMzygLMm71oEoz5rxgdefLS/cAKisb6KvSheJ4hpF/vU7dWFnra
A8qZhWqmGvYjseDg0PMfEk7c5dshQll/bP9cAOJxOD/aK3up7HDY/L7p4d2BPClG4AubNxpuZGQc
imNLIycMWQDNC9m9UCWh4kTrNNj6TPfwrGTZOEkokQmB3DKyi5Co+s20SrjxvVakXIy7Bf6GEzdc
z9wYl3qB550pBotcV1kDpokqrhGZWT9k9BNIZNroggf6tDbFxJEzaKmUUO/6KhoDuzE6VL1pytr/
7+awx5anRGqT4z2qfCjE5Gtn5EMWmyEkpBZVFnraLeKm40+eI/oT/57TSxbJtQ3NjhtPpKo0xdBS
wdiDRAYZu8kMYCVhtNqGCbfqFWYrJ/ade8V38r9NH7xpYbYtzZzvgGp6G45n3ZAoW6L7bYOegJdQ
geX0ByoUWHU34bDDW+m6tDHkF2H6IfjRANK45HDyVWoju8BIdiUJYbovAEqldJmyplu2kqsoEz+G
U6zEWpHOEs689qkANxBqYAePRQUJHUyRUJ+6z38gXfzsm0UBYZ+nfBpHcZiN7rbOOdiFcvxIZKci
HU3mbHB/LVXbRnLByMPnz6mXC7siofGKSXBcAkgLN1eas03cY7+J3zq/3XuFwtlQdLUaJNIcQuQC
HQWe1NGPFXPD4SY1qL+Sr4s/H2zo2bf93XwvNS6nUwrBHp3dFr1l6QCElHe0HhQwtzZ+ItoSCyca
X4O4n5j+EpmoT54S8AK9ZPfWkKGpRQjIjwaHn+IRnBSDakJq3WshIX5WqDWMNXLuxiFtZaDC+jXR
mFlI5c7cEza6qto8Cef76KkNWnq1WgQdvOqZ81MIGI91R0lM0xQ1SMKziLVyYcKySp5aHeRMH6zF
LqLGuOXVXDPaa1erg8QI5nXC8gjQJQe9YjMYa1inTt/zkONdCTWEmuuOtJeb8fERvhhEFcSOsSW+
/wq24sOpMo/Yq06kMa4HGk2etQQS8cj/uOCkJTiuogmL51WKh4M8YKUIrprY4MK/2F7IOb3sdEvu
sSvH7hVzRaHttViaXBJrhuncldV/ybZN2I74vU2EY9HNHMyYcQr4kNFzmZMqDO8BiL4dHhisJOr6
FFmqE2GEfXxifF8p551PXM6idJEY7yzUG1Qk+T2u8XQHtgzUlQ2vGXtGO83+LZp7v+nvZ66ewCW4
OrC7PCtoNOe0eU7w9Ik9kA6Z/AfhCuM9XzA7BkLbOtEj/W8uCCyiPpWR8mOnqAMe9b8JmVF2qGW7
pIwXF3XjNR8w5uKQP3U+z1SVHXwopb/Is6dSfovRQ/5O8RC1sUL8wrYnPObdNHIzjwy2f+gHs0bz
Za9hP2Nbzdf7ULvXZJud+r8D3VNYuIfTCPb77AZHByDfCPmGCTY5LEr1Tl95a9IRtNqbFtoJdhOz
JoNKmTm8MiOewVz2lVL6jrEpkbb3Ry9f6367qFAsRRL0wzCcHbRcPkEZ44l/5VkOEyw7P/fyJPJt
cDGuB5gsP3aRrCxbzmYm6laaxd2TMrJ/5O9qN2/mG+XkayQzCk4BQ08ZCIiRhjHvJsGUkNBrZKoD
JhwzftwcXcsb9Hx/MXvtj75Jrs5RE6Ri1Fsm1dMdn0H6x4J/+JptApROv54cQKyyLKWuXC+u+mSY
BPyO2quh8x0sSsMf17HBoRhISCvu9u/EnTHb1OfSw4npv5EBfOUThlE45pf+VIWNeaIUESjxcV1a
yLvW8IqhGhyaea4cPKRdlMVyHBoYBZO8irhczRKnb38EDm11wY/++t83bgp9HaFAe7mzturQLKiI
SFFC264FRPD6SwR5K8TeFp6ZiItDHJyjzLeJp4iuCqZtkH5a+ArW/gTT5c0VY/xJyYUbz16ibYFN
KoR1mMD8dXavF1EJCQgh7GXOcZBkqVulCvMsLFejn7+808dikKt5GxAy7PPWMGw9DO4l43I2nDMU
3BpFqC9vIHRSMOOYgDT/CdY6L5GQfnwuVdVKcaR/X0TwHgduBvPuXnXAtTpFjfohancgTaJ5bbrf
hfMZr+QkgG7Mf79GK7NJVucBeEA+h5opFxkT11VK7FQGG8Uha1IPsDGb+hZex5kW9j7q9mMVu7YJ
YMfep4NoslWJ9y1zwPnJtplUKniAjUqXQIshnbcQcSigZPr27Dw7GTySfkynPSHRMY+oOpDqIq+g
3h98CBgDo0PdCIHVUE0lgqyBwW7/gV23YUXTkvu7dAmxeRwe03PFTuu6bzmsab+sOgrZPbwY5jAY
yePMB+dXLdr1w0D9fMcen62Ck2MW/B2c9z6ZYuzUn6cUZbYPiV8IaCbBX5syrExGHb2+xZO1QoPb
4oO7nD6lKVUuhSYHWBdFaxP74kzZa44G2mVEQ4FXhZQMK6VhqRVcADf6ciUAeMCAai9IgHNnz5sL
BNKkB8ILE1yZKw6caR5tfmxcq+Y+1do6wLlQkdOAkXxkyaBW9h4vnKCTVG48HPEwvPFuOUlOKl6h
55PpKqf3qwm0mNr70RgJziy4qLXz6zEaScUxiHT24UiiKXhkE/kpeSoKrvb08DOVb6dkC/VE6/6H
C2ltjLez4laGw5w/eqVHv52yzDuDKtEaExDf4QvdzT4buMFLpOiTpuZC3HOYBAKAjIcPX02IM4TL
wVlKR8Eg7DNTbvVg1ginQOULDIC1LzCGOdQywK28m6LMSBmRBEBjtiUxuAF00YpgWwxIMmN4Q+xY
7ktvCn2gCAwf74euZqV/CiVSpnUMzj9u7GrUdjNoxVDgPwBye3JFUXCFbCSP+5iSY7WXWFOXW/3E
gokolR/MXRt7nbFm3MiXgjrjddDDP7zLYnMTkFJYxGarzgpnD3EL/qkVDl4VEmwNjOV4lZjDuEte
PzEMEHx22Q1HE56l1Bh/fjBV8eE0ABd1II/63IEYUpqx70wnopxPdwtdjnJYUwKZiN/NVW6yKSib
HGPlnBYNMqUFh1Hfy3PMhYeADFOVnlZu3lOo4BGwZKOwh3isZvVEnK+jKjR6eC1138T/FkzOIg5G
Ra2m+ZZFTlPpjJNZ+bZnzMCrNuWGjgzX1r4uXcq4xor+YPval6gEPIySHHbJBOunH7l0WC8PXSrA
LIsd0gnb9Ia+lAtw7Yqs8mxLSj8RruO/MT2cRqJ8gpM7iW/VnnoeKh7bYIG6kIAPgKiKLRI4eDuq
z0yaP0TAluRp2X/KpP6JrflwwuAzk0MGEXllpZDiiinGMF8riHKlDvG4rsarqsmAE9lRenbAFTgD
g4td5mE27yAohf/pBOxqyYW8am2ZVmQl1GyDWX1vZbm4u0umI4oPnhJQsuY1Xm3W4ezPVcSrvSqN
1oJi+b4wb5cQ3k79xbZtUC9rNU9jvKVsl/6Lmv4DzK1MJO8b1VeoLoxHBMrX1LE58L1GSn8T9ZTU
qzpKMtgmez2+jWk1kgGyrG4x0QQtEUD6JiSy5JXuVhcnCR9t/cYM10vljiMO13ADTCYkiRDpwbFk
NaWhjPOvsFMc8oOVW2BRC9NEuzcTm62B4cDFomHIrvtHzlRTCdPra4aVhHK3a40l+NHxXpKq4i1U
oGKyd8TQlGFeRM/b7P4MiRUME18dWmOgw2WcPSY23kOx+UXL89c72Ko13bCcGrbJRhUO/Ynvc/Yx
4iiRZwjheaJsQ7mniZIkErqNBQDI+9I533FigwmSapO+3qNZO97fG8cDOFslbpOATCKoc6skmFJ9
XdkzdRkEA8BLXyfECM5iB1Cv4dmlfqGjVEs6JQYucKfhfeAOABKmYtxsYMvCCGtePPRtSQXm/tKg
jUCAbMXWmEXmsqNZ8HX4XPMmpU52PBf+0TcE0NzztTtaKJV/IUClhHQ9cp6vMr3yQWqS2kKZvj9k
/Qin/Ozfpnsn/5Tlqwd1RBDsXkFy516irf3o3dbvJOL/TyHlB0hdmauxMAVJRAR8Nwu7Ob6yNRVo
8ecQ3S5nM43ZECZRRHc+HRJ+K7IlisBfYI3nuI/6/k49kb0a7Q6hjX8qnBvSAdgHN+wrSZcPTdf9
01Mc4NbpIHa5hRUEucNxpHVOLYS3/cKpcCBLAQinQWfaGhcNWaZoHPqWoyBErdw4VSoQ56szd/U3
77baXpHFIfs/5ruN3XH4SYZ+bX+cSvVtfZ4h2Mvk/jHxanGQhOqXRGFjpZisoJ5XNo5TPhdidXrz
qu9R4d0QTiVbAGxMXVU/Cwg3dmyEk8mstjoHmT88dtF8R92PUP3eIzQ1R7+ekxhlFjZgkfcE/bpJ
gOJ1HgTO4bdmfNPyuKztoToDNhANnpf9ePe5eyTjNX8tmjUixm+LUEKQ0+3YgDnQQx0yGU/1Bslo
SPe7fSGBFW1Qt7DWSsDx04Tq9Df1dK7jb62jBc75DTbykaqE9gfIY8t9yuxAPx6kvFtvlarE3yEr
oFxy48kAtRdAcxtMhjYMzU3sJFrsIvN62ezkb50BfLodZCwCDg3+9OW2EWdI6qvQSc1dgJL1N7vJ
r5y6Q5Bipr5et6jyfUaan2sBOoGtRuHch8SboWTDVxDnAUmlarz8bTuZE/x8BvL47NzZbqMTd0zt
qPOCSKmXRnGai44ElTfabK49V5D2JtEJur/CRdGuEXHJW1P/RNJkH7NqqggwK0RnnXrlrltYeLQ0
fHihkt+oxXy/Hwln7NYno0FpIjwNPhxOee1pKQlrrpHqyrAwue/qDQclK6NUR1C44IddRi31PcSo
l7RM/JmRZCW6gSpHvJRugTT0EO8QAjOtriKMsxk/ORao9+pibN6siWwYzqdvxA7m3A76u5IcG/HW
oBzb/ttB7MPVdPMi7LveoCM/EMBez6er5+H5CqYFIp7yH4OKo5+Y7pyYCfi9cKgryu0LvHTjSGtJ
E8MT0YTBxFHOV0L2zqlhO7zZg8PERMvZRzwf22LHIWOmwqqmMCu5+baEM5H89H8EaIl0hUTaeZ8O
mjMWbqVEkSv/46PSaBSHO8aHRAFlC363c1FvIM/iFVTYqqIluJHP/iF1sw7ex2sVjInJQcYyjv9f
kjFNKhJBgq577CErW+ULyzlr2+JZ4ADpKZQu901Sf9m74uanqKQd+7EaYQyRmif4oZYoTaUnW/I6
UWbrUsqG8k7MdNm7k12sf80UzZQsvQuLG4Pi0ly/ZdQnyj8V4Y+uSI4/TJvKfCeJ0YSGbtsXkPVh
58E/YGe9hoZawp1mB3JV5de74DiMQDJo10AWmRkgM7rWl7nAOzAgDleaSot5kXQqrN23wGd+1GL7
3fSYvPaAiD2UmMPsAWK6a0YeJiS7gUKikRqE7Ihn7hdLbzLIuHLneCsWJPQXvLPuEB1pKGnAcf7q
N8vBZFVCzWVgUKqrmigHU4LgwtoM5aarBuuRBUGgBAUWeLjAzfGz1VWUv/txZX3NcLocfkWgfMNm
0IEAjQ5QRT9laTA1iQO//LWouXmKwRVgZ+qHyljAzowxtalXLXMSTIB4Y6a0B+VW70r0L25sMQn3
pXjKa3dXiHC6aV1umwkTx3NfdkD9/BUBznTJFahLM0IA00p1F5H5NtPpS6QXngzclEsuHaT3sWEX
Uy6egbcXwt8V2siIXk1/Z4sL9SFuQhPBrTTfYZVzxMOzgY0ca648NrusN6Q6YT0PQVbP1CuoFQrO
EjV93utl9n9KH69gn7eQbyd+7YUyEkMoPpebUyULpmewPjsb2mN4Q8wW9bgMVUFzq6wy8plz+Bov
7h9O82iHENvSLSNp+FwlLJXkNBuAYqQHDSqo5GY038F2gids5CT5P2LugoQma649v/xKGqpGwbDZ
hOB+yW9urTWQfm2if0ShVnJT3dWI37v74bMaVKcwPi0C6LSUdPtDL+sgLJ7kFvISruXcOQJtMiVu
LshS29T6a8bxm9NdnlHETd9C5S/F8VXbjR+bUUrgBhlqz2Vixqk/8tt5E57QNiuKKuCDTwIBmm16
qNkLNBnX/SB+QQz8sVSDNVp+sK0JQ4s1ele/HoduBhcCQAkD6JPtK6oPZoIPmB2IggwOxT/A+Qij
2mgL7Rb501YB84SG0Zr3MgQPLOo71jdsdSZ2CexQBbVhmIOOUl6WptWzoNy174xOTWLAi4DDVOZl
9SYb8inTFCbA8TOgli/ti+/3V9+WFz8Mo7gU68wNeNoUYaqjyKUQZ7h/UjJOCLlZHr7fFw/ex/Ec
HlxhgSY3jXITKBPnl+syKTNFRcW3MqOoSSLZh3euQ1j0fYaHEBP2gS2hsmDF/V1X9BMl0bjDlXvU
YAJvd5Q0NFJojkGHGKIIzKMcZIfWI/gGa0w7jJXy1nppuig7w5XcDSIVRO9UDS88FY+ScEkG/5Ri
wkEXDrorN3aoDQD4oWWgSTXucLTGw5jty92/43ZXOmBvGQlU0IRLqDZ4O74FAHQFSanFa4L2M+yD
QPjNePoddCvq/9cO+jUsQMuTaBo5XbRwCFeH+ycpQV8ohEW8N8iLLxBvT22iLT7N2bWQgBRIHgz9
LQNAkT7EUItU/Ut+SRz6IMCiCF5le6Vg5z3Md5lCwOvDaqbTWlo6oOGfmkxmYBgQyUwHpVxpAmF3
GHu3YtaiWcjv4mdzpEwuV1x4bWxICzKnbx8+MhdZooOkGZCZZL8tkcZcopRF55IH/OX4H6gK3oBv
o94SBCaeLEbMLRsd8fIhz2kl9AKr3Gho5+rKT3KfFK8A8BVl6MoQ4oiFPAWxf0wJxroORJHHLojJ
xRG2rqkhtCgNEDSgyihwHa6+V4AzWdbb0PVWPnqbBSCgN/7H7szszm2eNgwsH2pS22MPrYF7TJZM
donW6q+IrXqiwCGzikjDY84y2o8G2dgfXKa5nC/FnHS48KxeVxoQFZIp+A4q7VkUbvucmTp4978p
Gd/3CoFBp5L320mXiJnSz1zA0NOxJaLCgTOGEDmIjYsL8iPkoyc3Wqh2qEzVdPJHWDlrMspM//Bi
wl6Xh5dWqxFMjfxzJFemOR17hNsnP1ei3HfN8pz8qDGwD/KEdOhjT3Go/p07MW0I5i0DnMTwfgSG
j720F2am/QukLjHoC9DTQFCnwR1ByUptOtdIiiFlos0KRA12aFUjGjJRa2trK0QeDaNIsLokmY1U
qcn9RAsgYK5KTYOD8ZuMZhe2LFibUElkzzGvkWXroP9JLCDiN3lyKMjCc2zcubqq7UiJS+ms2ykY
enITV1GhIqYLwFHWpLbirxHiP5UUZT926Kb2u27Nxj6t+ssvKGcwU/nBDfh/2F70XOAcDC2bA9KP
TcFBzu1gbYZxWxfAcQL49DFPgRz/ML4IqVRW5i0ONaGu3ldVxDin8qrk3mKu2qclQqM1nndQ5E3O
s92jsSZFPunODhIb6NdEUlMWK0y1knV4wRXwFvmQ8VX+lW2n8U+lHLSxvJPxlwu4nrfVD4kdU8Iy
cCo7Z1D0y9RXtBlsOZDNJ/KwH0ZpSV2H8y+aiuc7UfB35oocRTMi7QSivwNLuXszZF3E7KWFSTwo
tPz+II08bB2xnRhBQdOLgpkvvLyWAtdJbP0xlJMMD3XgQ9DSbo9nRi5y+oEmoAk3ijloXM2SvDuP
aM1/CniswXxfozy77/YL7XQa3BPyoKc9HRCg6/DItmbRB6+q8oK8zPOfKCkkfcsAkY51DVLf0QzV
xbw4fktnVUWcQQUpH06kkCvJWdf0ga4i3bT4FzibIp9mfvKHv9N2RIS9N25TbADZzuqA+HdymUJE
3UnOyxJP1j0VH+CwUKCqtKoqXMSIj/yJhpQ0MRLoUwwlgtGrCyDd2p61dlys7wwRFfsyjYwLtMpT
dnMdfCOXCinJFl5LBafesOfZIujGeye+M9vWUHbxuDMM2WGfai1r15gHSOZ0N9qXItb1ox2mDnEV
x54SxOksoHC2x0covOfyU7/4Tu0vMDYjubaypFObTcdbE5Xe59xp215F0BwVxn9DFzJCM+NU6J0f
OEU08F2PW8S5LvELQ3BYRKMV28licwy8vwGrJgeNHDP8U08OdA2rdPLBnPfB3Zy4Oieb8YuNRESx
g3OIm0o+3q8rFnM6nONkWYpIH8IrWap1xJaUOWzDOoOAgT3KOLFEFyZfpBhdx+Iqv81+EOmOClz2
tRUjBz+FFJcssthnurH7SE03+Ke0/IS8SrjzU9qn3tYHF+ShfgMVT+WrC/nDJJctDqYLq5R/4AVt
CoIYdTyYxNZGZHHOqXRxI15UYl4FUVbrXuDaBEi6OBy71bzQHWUVCdfBFIAxhr0BM9k2Kt+4HPix
bAihpM5i2kgTsjk4tp3lcrX+hTCQe5ID3NduGayLLMP3SUET5Dr4TaB/W6HznUTM2qQc9IwnIfu6
0bnrpYFwnJsSwb6duO0kpYl3qjcRRAcXdPv5FjnO10X6RAj38RAWRX8eyxxXV2u6SUILFl1eWnJr
GadYSRvtQqHO0nJZalTsrvcSWy5gTA+qZWZbwrrFT1IYYisnHZe70G8vAnO26UreMDgwVaJgD2GD
Y32UvH98NfnChPffRthwCKhaaAki9LS2L86Mm3jwfMxfxmXJ0WukMwt1v8V0hpQe9OIvyDPeV/go
9vIvWMfkhIG/8enrbWwfEbK1TnprNK1NIiwaAP0OC5HBujXFtIBk/uqKpmmGsrUYJ6LvOsM0K5NJ
nro0OCyDBGoUR/wnKKFKb2GOSDAhmwnPTp4h3LcrXeioexVZsDl7I+YLJ1BebNbrHftzWZ0tUmf7
0ux49wqH3Jn/OG0DTJ3HL0S+rdEJ9bAfO7FaRMdiVjoOfoWQFBUVnDZmXEQQ81P3NnzEN6plPx2I
H2Hdt50WTqrPhJkNsIa2qM8h8Y6+nAQx0LHCsjOr3Gqtwh9c3msydxYywR5e9NuKkFN5iZSqgz9E
qG6mGNcMalqbS+xvTuF32WSimW3GpBXIkXAQErGmw8vmP3wH1fH46/fRU6bZbl4gI8qwU1VvPH1H
2am6Nlu8LmIPLnuqkqVXQqnRJthCFEke1UvzX6Unxupahkuj1d0rNtyMdx2Duw8qNeOOTqg7NYFo
PcG4UWZv3WTHnb6ivcjmCfJReb0xjQ2CMHR3Olei/OsxrlYquwdqQTU/CKDZuIM5AszGFCVLMqLb
qyo40jRapvjn0O6NCdgYOufBrkq4xMWVYMznpwvqbElmrglRbvE1FH6l2hMtXEB7PdX4PkjKpWLs
r8AV1leNzYvoKfnIxFbRBWOCsRy76TNG7b3gyqZIcRgnzvuUM3PNPdFYhDrn54ZJzYo99iWTZYRS
puIhPTJVd6Yc2M1FxdKd+UZx5K+TsjmwXBpa3cjllK+hxLNc4wMX4OMrPoCDMwDiFzoV+SPgUKKj
uZ4UICGOfdhHblnrs3ZhcpVy2f5K5URif5wzhyk4NVHaTZIbxxKx8IxyFeWblQRxS25BQcQLPDRc
K1kHddhW6Z3L5yhrhiufDPbJ0xr0E37hhqXvPHyDfZMd23OMwKoLElTLZCZAAghtEZZeJ+zbo4mS
YN/Qe0AKI0ThHCq5RxaNqf8rDz+UMr9xmyndhOtLwJHydJzQpPEpvHs4eMCCqa0+CgHsclzB/YvP
u3Oxdop9VBv7Fi12gcZRCVb1Q6563euRAveHoYum1lcNt+SdpvbYFGFTMvZ/9eytM0t3n2Voh93Y
hkRbw9Nw17OwyCACWI35X0GA0D2ngViOrUrTRqdH5SmOf1+vJtGYLTJaKCZsAIRTTXUUlbcRNi5K
NbvPlL/gyGaOcQn0uF8IayzK83OMVw45MjDARHnsdvhi5DQXK6oa/3K7fMy/Ga0mJK642qj8+Mic
3+9pR83WwVhFV1WFDuJLll6+T+JEEFvPMgwVlzHFtTK+vaCG0SX4y1JDDl6jhsxhLcO9YEb6p3o7
ve5auM24M+Qqq/cYGFe9Ugv73Swq2pw9LtB1r9HVz+j4l5fwf1zwI+6csEM5L7DQ9zRTBwJW/Ou4
UyVlEasY77RRr/XS6iR7zVIH9CQiVFf2v2L3yOiHTNake/K+W6p7Vh6nN6LQWZr/BCavSzczwNXJ
YioEn7DNZgtxy3GkLnupLMfywws8G4wsggU+xxZCs6V2h28U96uvFzgaCBocmszsZLGOwP10YWH/
VM0La3pDCjJymZ3PTzzWEzPaN3dMoyYxYlU9V9XjPSgn5LunmTcbTVRiA91kiNuxRTntIudRvVRF
q2n5seuxDYz7d2KbjIELdiDtvaV7t1PCO0PWIj1epHT3MnYZtWZftjSKpzePAk1ULS/euranAxQp
oB6GCgJBKI68vxjvK8bRenghGArGLb7AHJ6ejvZJWi30lJX0H6ULT0+4jP94rTPCOIFBsN43+yAi
DjU+d58UNY3xxHYe+r96L1OMYqVflo7DvkYZEWhkVyNfQU5WXMG7s32Lko4UeiTSG/T3PEhAcXO7
VrkysmDIu1iGSbkPYpcKU+1SwcJJoaIEsaRHu4azSLombg/9DUzmgem7sMx7OwVaAscCqrxhfgRd
CovZDjQQv+I+5b82OHiEg5MPUUnP7hIsA0vp6jtfIKp8RXbWE8OCQCgmwIDlp3eEi3NHVV75wG1G
v9Tqi6ZCMt4owg1Qw/+Q+AEsa1/qRXKxMgXu6YTPkEp//cBniai9W/5lrJlPy8uJczdbyOzuXeTN
bzcZ5e6o5T4T1TFoTTdgNyUNEpBCVXBpdyUF5C7cy0tBa8HkpjOL1YAAdoK5pU1OnD5e22Je9beL
Uonr7TO4meyxc4o5RdyrC7QA3t6fg31ayMErujD/Cp4xQrNJDTAHdUj9us8ogtaOJ960L8b9Qn1L
gg/17SeRk9FVMlpy/iW5AMFCri1SGD1gHljlCNhSLMLjlbVKshGJkzagmd7BwA0kwRnqGYjV51hL
Y2dXdfxfml3CioQ+E1MpfCc8RpXtXjmq3F880u0r1GIMBJMu+tLB2z4zcsOO4tXhxTgdQEaZ0w82
OEGuGc6EbYX2SGHLSqNe0cmM3fo7ZSN7pbPdt0LYCcACmNq7ET9rENs4wFrI6FrNtGfrPoxXo8Bm
Dm8JKqn9YznoYQPva8hsJrDNkAxlZfYs5zmhtjZN4/EWlzJaqzUKiiu2KmeZ7GBj0a790t9sz/xs
0Ni1LscWMMnCREIFGuf+m7cZt8FLY749WXc+od4Pp88KpHblrw90dtpI7wMhFX5vW3CSLLv89cfL
eF74YddnerBLQcf2zWVAU1QI8xzgunF0uuT0bd5VFfWHz8+cMV1Fky1B33gWcRpvvb6MxI8v3t6n
63wj+IBPAicBniJ6YdGjyytJKv+0pmqrrxh93ECM7Ge8Di7Zy56kc7w3I+oqrV4eSfDhv3jX0A+v
N2JtiucCrzuygV0wQ4ReJsUNAPWtN9hO7iwIDSjUtYDhc3ktSn2nuU1PO4Jw/zmQZ2i4rDt7VoMv
/eLjccXbOi7AseOOgSjZzMJRrg/mOpNAUoL4gmWkdB1oR3tFDeWvFkIyJjB9hZRo4PzdQCw/N2Ay
QP0vr3MOwG+FK+anPsmNZXLLwN78W6taLsDGUmMWGiPV0CplQYVGIdoV1nXw9XQ25PAbz6MkD74i
3M4QxFwCsOVumvKuLPflxNw8NtdMGFDiZ7f6aobcGv1yvRb6U9hFgLe7tRvTgg0rVVZeVs/X26HA
G9IqhIwaMOLZpJaJLfHYIHXrgnv/jtGoXD6teQz0vn+BAZBJI6U4v7fHWFXpusQ5VD3IjeApmWGW
lKC9bdSZ/B1BMj4X7MLurcolu0RmFyfgHtIGg3G7lbkZXsv90iihqHI8+lsKS0N3djTDICTtVMUD
Ki3HNAELynl6p1SQVlAnqUmrDkmCU3MCh7+tnmlqXa780BgcTnyPkvWW3EJEySmNxPGwt15L8Oe+
nrTxf4b+M7H3anzjb7qzYy2zMqD9BSFtZFc1dqucxf9XstZSceKdt0goBin6qlNI64l3gg5vRJel
w/yy6cdTXRHWhQQYkrWvPYAHdInvlVxzTFTyHgCSuP+V65Z3fR0z9JJMj7FYbVrd0ZeqcqoytgQz
HfuCmtLkNGGgHapTU2VcQkUH8J2u6Ec8WSF2+vO8I7M1NN5rbHDspivClk3f2pk5lKXvYFo6QkV4
PlB+0g4WB61iCpmQ5cLSyjXaSUTYOIHU99BiEyQnjHJlYrP49e84hbkl4ciyd3a6LEeeGrZ9fOM+
r0oLGRupcRNgsGNFgU1x+WG6fpZd+8R7/4n13BLdcDULTpyTs6KqZwl70dx6yPp7z6I/gcVxq9zm
2UX3n32R6lTBzxNTJL4Ylu7upC5AWwmt5DY2XsQS4iLIuA1QzJIoYg7LA/sq8SqObuzqF0J3SHJ6
OcOm5XduHpViiEv4w/giIqL0s6ZiBumleJFeybaJE1X+wV1UNclaXl2kSGZ0+wYT0lH4t/bcYV2f
74Qj0y0hTJTBzPzkwVjihob2OUkjUcagbH2H6aNHVDgh0K78G9oQjE4IthjG8TdJlbm3YO0vt6Gc
QQiCKcZ/Db/nr1GoeIdhvNzN/qtnDOkp8Sw4cNtc+h/q0MIhNpvVBdkhevishtN3hvoPrKqsaSgw
UeVYc6OOpibQ7BaKagsHyPtmVtH6TuPJSABHdlsrKfBsboQMWajstszfV0k7trqz+s30V6AzC4VX
Vx5hRgcsQD0RzAMRcptekrdxg9mCS7giErGTZg1DLUdhmsfXCqrsjJt5ylU6+L+SPdw9nGjJwch4
JZURvaI1b0c7PWpTZ7GTZEiu4VrJtFw5FXie0VLBPsd0j9cKIcn9x3XBgWbAfk9u381mki9aOGLT
nLYWPgCGCKbct0v6zOymjECHbI9fgboKrAt51YE3sIToY+dSAgxDKHWwNvikfyGic1bgUoB+VPcR
I0GN6qGAu2nGNffQE/xJhwzhxuAvj6Qm/BjvdlYXtuklRMgMviQpCBGKd6tmPGOu6GZDXIxLKkvJ
BMqusniHy94mvDCstFsrieNZLOelk47SckKO6pjnlIy2PIBRrleWMjXOsAI883DnBvc8oPm9cZ9w
aG9gFhoZFlHNvk4cG9qhkoQsZrGuhNx9vO79aoFnL9j2Tm0ldoWKNAWbaa01A0IPjRTFldYeQVx0
lo1VHlnmJn5aer0XQ5o0T4MEPpFrb7Zg+3xx2P/Ngc1Gk0IysYy/F4Mw9zlsntGGdWq0Yh/lRH5l
tfjgzc9D5jkouApQUZJqSZNTVb5c6VfZA/SJ0cJvgcvLpzeonVH02PPMuR8BoLYf9sssoaQJ6vWW
SnSyVs9GSVssu5fC/9WjiXF8Mm9/ucpXNTe0R8biyJCRTh68DZh8C6uJt6xviKxh3qyNuDuyOe5g
Qf1A76EyAQRidA1x9IS0pBhynR7yyFimnx9wxOzxKcok+SaONEMNCv48K5aZvk1lSBB9x7Q/XM3C
4QRxOzuFX8SKuURUUcYK5LOlHAKglfFGsBQ2Lo2mRUprDzBeuide2+NdirxwC7MaDE85kalOZP3L
gHE3vh5ICbmLKhWlX0IouiThpuiUX+PDwe4dRl1ih4j8GbTfZYS3qdVHV3e1zbF3rX6FgoXGIj5B
2OC9Sv8s8CM0xOC+eck5Jx2AdW51RzYCYYDHt84YlbVE84+WB/SAJ+E4z3KwS7ibcE+9WhJ2htzY
Mp2GHI3NrKv+B/+TSHSo+Zpteevlu4RxQMVMd/F4m9+bEGd11qggLvULh6ZUKJRIEX3Sab9N7qOC
GdLX77na233v2x4A4aarcgH8F96ZjpmzpLkbGZALFBjT/+7jmDUxJJXoQmfFcpozc+ZQ63d1tjQS
jiPAdHwODsU9OeLqOU6gtNyZ+h5il6LDzC3VsJD/D0PUpbqiPHb+hx43IYnPn0XhqZYBSJBLKT3O
SY37KJIXyy/d8OCM9ivXIzpCJo/yYuIsZ5LCs2CkkPjDM6wG+KGNrxgsOaGucCYlkuPfjWdP113G
pyllmYahSJxFPnZb+qwPEudUHdz9m/DyPuyGxCWpJsAzOQE4MZB7cIrQh6BlSeHhr1sy/O+gEGK2
NXVZl5phQ4Ga8oI8yHRvo1Tmjkmx544QduOXdgodpzRDEAuieafsndSbywyKJ8u+BmZzkgoskpNV
mQrBBwZKofw9GrJTRmVYd2X1uCQNJVbmviX0F9sAcmQMFSqy+7BEvFd/1KgjgIoknHw+WUf0psbd
16CQNhJViu8/Vh1XKeN9amxRvWBX6BzOTEsi4gjOlh5YBmynQQyOlRLnl9yZ8vpKVcyE4Q0veMSe
2/bjziBfDGWAKuFTImbd+J8qXYl5NnI3NF7Z5srizKNLq/Wyrc8wua/+s9PwaE1ZzA6K9mLj9vXI
9MwkkcZ0XyBVAHA/P7tck5mFuKNSfVDLDd4H/Jk46a1G8yOI9skIxRcps1oxVtplAyjVltO5+So4
0Zn80KoQTNBVw88FxabfYqyZa8kssA02CzquLR8c8nwPAdXiEMgUP9/e/4mxRs40qXoi8cRNNF0H
x6mkiv4rHN+YjHy06KShLutq0aQkvGabjtZLAWec95Pf4inzz8+6kdS0ObMBoNl9HB4RF/rrUdtH
gk3sHy2LRPtDnYhoUoz++2RmNCKbyT3uGukFCd++yyg0LHQnBknXUCPkyG9k9Rg8aZynbbbzu2wq
oHzJzg7K4tbkWuslmQnv46pKBhl3v+slMcq/O20+6lVoK8MGgmI6Cy0grhwXkht3y8KCQ+Gr1OMf
g2eJYgkkHed/j7Wyb3bGlqGNqHqRFT7ZYDPHG+msmlAiFntP/5ubiFrEqLn3rrpOWazVr05NSawk
DF6ZW9rgn12W7M048j5ASsyIf5aL2vY+4tK3ACTVsaXiBmbTlt46jbfozWwIgGacaEUFbbI99o/I
Fa8qVVyZY3scNbmU+GJINb5hU50AZeyzudjDE4UGYbn3E1+5OQ4pnJJ5SQItlNUO3sPabH5Vxf52
s9lB4ihFkuq9g9qVyHm40kGWIZcNjdr0duY03XnG691dXD5eROJZn7IMSbzuHJ/akCMp0Z7ROYzZ
otwUSPUSP2i39X9XsVwJtCUzBXz9GqNmGbMYP/ALppfvDNOq8CVvMt0jWUdKVta26g2xSLDGwsHm
D8fWzKgkdJ+Jb8s6ENKTC8JAfr9ANYZt4baimO86CQIDMVmSkPavUDRwSHh7LCa+tZUH1tAJXG0e
lETenFcAQVAnaGIQvcV//JUDgWMFXF28oOMvByMJ+XLY0LiKjlYYFeXkOJkDJC2E9voR7GwobGqP
qNPkvWbB+ES+b+75UktfAQHLJKI18UqqZgHPeU3Oe+n6di8T78rokSV2KU+rTMc6K9a3gcuwKN0I
khhoE7iaskqD6mLLRjeAsr33ekbstz+hpJ8MJIadusUC4EQHAKrX2itCju592Z+nrifhg/dQLYVC
YsE7a+fANo7RJWVsBXkmTnkWvcrtLWMJF20DdziBnPOwfONskGnKlBG2wL0J74W4rO/RKfiZPvG7
FkK1Zm2XS2KFDi9EfPZDrYMHl5M8s02uvtzjK1aPMizI1FmVzLQxREyJ/WCz2+ObmtpH/01p8pdO
mRlIynB0YFZvGb9bn+qGqbO54G4eHVAU8TUHPr7SQpy+SGNkBbQxldm8McHpso9z5JTqqm3Ny1pA
B9UMfv0xuf76FWmG8gUPQFluy6W7x2VohoPPWKpyh9fUK/7Ucu5kdnvQYTEduQpjGbIZRchRln6s
fwcSR2CFzFs8V5Z+LoxW9z2kKO5Z1eImiGpiR5j4fh5eyFeSm19ikL6ipTQbWtuz6KISaEi4b6FR
/BxMCzbHLAR2AC0phq4w+sNZxkiwcPtg0KgzXh/Z6iESiWkYkzK5JtvOa3zFO7taSR43jeMOSZkC
6xDrtur4tTqstC8k9bcpEOylIRvhM8Cy+sH0UYsiZ3cxXaJ2xT5dkPh2fEXk7V9Nqfihhw6StO3v
mShsLuBrcWver+N7bHsWcwFAS7BLzvZkM4b5VmXmyJqjLAtAvusfXKrtXUK3pnUR7ZGRdGcy8ldR
aWrCfExQADdxcqmpPISNwnFM/9l4ZEmx1vO7ALn9wPXoN6yDwnHvDX03OWIiBIGMudOLAtZXJptb
UDk3SasjhXMYNkKXlffNPJbV/GDE5ufKMe7WCOYFfXM8NLtiemWIqAeVA/aeG1YZrWxfw+ItLR9u
skY75rVj5/almlfaggLdcgL6eL5aPB+g5FQ6AB5H+zIoV9VxnmCrADWt5+ewW8olyv0j+00kCP9E
xKXJmskvIcOpTmvX007UIu8CnbxwMebc5hKOKgR47JYNX2alfm8kmk5J2OgP4tT1Edd8OH8o3KbN
NPlE4KnXsZDhk3wDA4q17qZ8NuIfkQEEHqp6XNcUjD6CtC2A2NJ+ejVSXooX7QFDKcsPTIASkwue
U7YsLz9Mq4S9MkpPJEHCvFNkMYo0LNwZhGgH6bqEJmUSu/r8+HpMe1+ELeuTEbF4rT5cJfQskhzY
4dYx7UE5CYKMq7vkFcOhzAkKf45pVB1LbDXF/2GNndGCZTkzxpW7pokezyN9AF44mPVbstzz8xwc
T8+Rlm8fg3yEDQKykxB9yRz5GKFwrJGJ3TSajMHAr694zx4ntGheVzUd2jqevGJWv3SgPVrs0UOV
xwzhViEb8RWYtvEhye0+jn2zAl1dr6uzT4jK5hvB35qxIHGKYoE71Pm0y0KOrTfsGiYkBTR4LRB6
u7rA/detjy+ylyuDP84Ajtu+WmBypRPD0AfVarFSBwtu9iIzygRXUQu3bNKG/q6PldGCMj1qiewy
KJcTsz0ZLN4SOzr+WPMJVyRqLkI8/Uv8i8TClQC3ZFihA4ZhAC04q/uFqdHmHYwNrWuculS3dU6O
SZTCsGtti1wWs1md3NBwHShGr1Mdke8MStw5+TjQ7410ItPN5BwtSSQiiN12y/6m+RT9cZ4pOjZQ
9DxCEYvo0ryPQ/J51odO8jwivurIiO2WFmZJsqGojfJ+SuYjs/lnkT8xOewf8N88Vs+sfEYz2p1Z
T5dXm8eHGGcydpUCfTTufJOFDRvLRY+yhcW7d4oypV6QZR157Qtul7dbkMGbtT2VfPHlBNJzF4T6
S2ofrIehQDcBusZyaEjQHUwz4h84wf0vhM8UsNjPgp2K99+VfxnXlB486S1b2U4IidhikH5tVkIk
j3FG4Aqj5vUr+6wf8Wp+L6Q2tTdbnpgELAf3YxHi/EcvA7jDTEkNyd8e6kUQ24QFN3Z/1bl3wE5o
MyTfC0AUpw6+1HZ/IRh9HEiAslqWk4s5prz4lVrUEf+yiuYG0IyY1teo6EsWTU3AYK+xZLSjB3Gx
hRiS/SR4hp0vLs633wLpIi9DuOrugO62/+HUbgPEPP2BeS9OEEmfxBtJI6nF1HmxAvz09LhXfQKy
879SqQ76jFZo5r7Phuty+VLU3PsQfIW+3JumuqJPwGjn/vJY/eOgYMFdbxcvfxLEbZRSNqvAJYVg
idBUDNpnkKXURIPwL1HgCuXwAuhs2jo0PjZf5imOLhbextVajbJIyjhynN1K+cv5eMFXZf1bXKNt
ryoZD2WurguaPHRNHD5szCH5tMPCX/YG8lmlIB0I8dUAud1bmawsQXJPgC65wWfa5K+ZsiHJLHCp
dMrH0gaMiFWYyUmSRHxaMQ79rHazTQanQWh+VJYp0Vi67vkLJs7mU1qOHKELnnvPs6JrNqZI8a7X
jyCvkY71GK5YeAI1yA+UL/julWmbLacZqUkTdNr+iRrKP7+m9sfkEpQqj1WsgkO4Gg+ndx/dFTzh
9hOih93GOR2a0R08eHvB6BKbifS/1rAhLjy69p32FAVb/TkHpsSktADeH2WlDE/YrunxBsX020mI
cJKnq/DBeRMizfiunfYk0JEkW5rdsdgFyAAHoKpe/usSpDg/Pa/Xp8a7JFeBoqjUSsFytt1bGhuJ
lUG3aVUkVFMXtHsOH+ffInxYBgyt0Blprlb8YYhY71jqy7IPcG1XxVNRNNuWi9WOOW8tDRlsp6rZ
Q9H7Dw0O+4lijZDh1w1gD6pkOr1AjJ6MDmjpsdXMAUUL6Q/npGI3v0iLSvFRr2fFhmpqdvKXz3/x
pqasQFWWmk/T8NhcbiS9EBxIny0TmFa3ms2YLN1weFuU2qvg+ONTg5UuDS02sK974uXOMlJ2q+mo
ZOfWGZ0fPhdjq13Mh0mYYRXq24b0V9tjBRhf+ETuvjN/b0scNFXsG9UeOHj7WByqTMszYNslkr+L
s+zLlNkcAE1XWCz5EdnWFnPeS1rasISY+8txyDqgdH6DRyMbfg2sa8bXEqu6x2vJ42JgJoJUvZ7P
05mQ/UOSwsAu9tOk7zFf7VdkXpF1a6tnyRRSV5KnB5dIye3zuaYiKfO0rWYX20K9Rt6nWKyFfBw9
wq36P38aKdh6HPSBt+sa+4KkHtHzIKabRZBLLecP9Jf9AUm3/UEO7ZIyotaxAVGhPCY3+fYjX3FA
Amn8BDG6GCgoXI4y1tJOAgE6CmD3ZohMF5gdrPK9+UxqRUCJRXXDxbK7iH6ak+4tKDXONAEJmjNB
EAW87tKoJ1YgHwgqgQe007zE1R04h/nJmdt0itgqK+VzTRgUnyG8/wG48ESNe6pjRU7XnRjZhC4n
zKIjt5n9sm+5mg+lIMDZy1VuR0q6vXXPD8MTq5CMiykbnOBGyjpAbRwB+2lN1BvJxw/IfObW8gwO
s7EaWIQpEzg6BwDWxV2v2yzn9EojYfzbfqlety+v3039YqjBv43FCHUOh3jA3GThIWx9WMu2AeQ/
eTrsUWUst+rnl8tMu9pkxtnl2rDiTGVvs8d1WIcHEiI5OD1llH0XWZUQQgNXuthEwNg8RXXI6xoU
GDbuBvBDgSyUSOos37DHBcwbUWDtgIGSpDDIkR7qFBNcU8NuTYrLkNsGinW1iq9QvKvJGOJoF/Xi
RNR/+We7eTVdkP3chPI/YmaExHcCesCs/Hg+lLXCBWyU3h0HzqgR6hK0xpfbDM21HN/aFajwhVgJ
RPt8blZ8ZFYpzFf7KjWTD6ds74JqphcU3H+k8sUad3uicIkqA642DS65oI7gtz9iMZR1QyDAPFWI
RBqdZ4EXqRcaP5Co3PiC3n+xzhOteR5Pvl3GhuBGq27MSrb6b2YnkCSnL4eeQ4Xxu2bOp/KrOSik
0eSsx+Fh9kfV18oCRRh3X9Y+5B9Z9x8YqbtlmHk0nuEtDyBgYUddYYqJo8SIGcNKRZVXJB+OJBYD
n3bu9Ea021oKbfMUfRjp5G+AUCUpkMs7VFhIONcUbxvicWdJfG+qo9YUJfNbmzMePfrcG8hF7z/r
mys8U3O0ac5K168LfMmT9xVh+9weOnWHafWco43P19clqis+pe1Sw95pOj3K3kqj5eiS3+3sJWnn
jisQNXecGNBvvnXUVvChuhfSYup0186WPnu7x8OkXJh8YYixoPgqi0SJMzoGVFts2B9G9/eSFwqV
XXax4P8qmHBrPTYuRgHrIoYSOnh9K7WnwCb81LpWXA2Fd4R4GijkuK2TOcT0cx5KnI9/Ntv0SKrf
YOKUuTn86X8HNDGlHUQGlrpR2JXUx16k5sxsMDcB6fF9pe+o+o+s132iRszrFLS1+gnBoFT5rzwr
gnHspH2tSrXCHfX7Ny1CM4fPvZmH8vOFYHgjwob42X6Vdky6I6TdQHkCRm3/u1ahl2aj9DG75+m0
wyNBSJ29XJRRivjGgHiah6204GfUgVm7brzCKdQfFOjR02p6sm/OaJA/TX4DmcMM5fLSuM2R4IHD
mz+BuoqvB1FIK+rwQs81hVOuDY+dLvPChFiyUi2FniqHCOUEQzYPA1XgZhTjYH+MHxf9NQjYAbaP
YiyOuHjLk6+C/8JT8jn74IK395Z3SjKdSHd/3lHlujhPBwJ3dYaQR5ZXeboeSSrVYXwPW41xvMvD
dEg4VmYsvbg+1oIgk3dvmxy6KYFkLhrJMMV0EL3Zxst7rwpqvUK7kfBZmCRu5HK6YbuBEX8dzgSN
Nl6/W1woPvelF1pzUnu06npyREbEqQlTUE88TK1uGj+OAWT4m7U1BGAXm1cA60dI/S+mFa2PWQyH
S1RD3S5syuzgrMJtXK2C72dc4WYASBxbQl33HohZ/JUZnqp4kUWIcTJlR4XIB0jqul+3wO1fNRhp
dHRuK3XZl+BYXnwi+Mz3k+lIylKShanrHOPmTo2SkC6vSRf33mOOMJwrbxxliYFWcg0gIwmnvJH1
TxwvKEzgRVMVbiQAev1PtvyOFNSqUFkXV/PGhhxJ3Ab9acpArV1KexzcCAU1MTgSGe/lvy8ggqt9
omjcLLs2QQJ7jpRFmyle+tmxpKqy5El2/A2Fs/OiFFhPCMHaVsnnyRuoaHzhj00vv4p8mM9hvuDe
LTn4CnY72NXRApBw7g9tbsKYu11ZqyU4fwknFqlqCSNp/JjpHytkaYaEcUAPMzWe2MoA5ilWxOlj
QIdltfOccqTEKhWtbq4XXDL8nx6aNiRm54QqMS/PHXy16d/Ghv3rJNi10kgFV7h4pBw3H9jgVS3x
373f6md0a4hYnUhpUbsFOl802UW2FPmcZuMITitfDSSz8bDrBdvyrT8Fk0rKGgr86d/vghtyZ+Fs
3KCqZxV/CCYe+K6pMofLwbu7aCSEPDwHV0uLyUKeLVLmKeZ5L99ctxtK2VXd9Pau2R7Bty+sjxec
m3IESu2zaHJVnbL1aV4EWkioB4+1ORD1MoZh7/dBxYC6arYBbkUGpbBMxF4dlex+xULZVwwbn45R
2g0A1jTPdyccc0i/dTGUGTQUDFTSPECCc6kRkHludDDBtljdQXc9kVTFbLRO8H1Pmb/WinJO64xL
0B0+pTD/8DZQpPvzWcn+UtW2q2E5CniNpJhe21HI5ngfRypc+M6ms8BNktlrOYooGYVRl2L3/RAb
aIWTwSyDt7MmpVoslZAEA8MqjE7A/UXnpBcv2N+d8KC8o+QwL+e47PbOmLrgkRCAhWLaIPQU51Q6
gxgn4fKDRMJw3ASpgLxkZSuRMvaS2wtseEDtubWvQkBZUlGhKqBEX35b3nbmFUsFGsxrnxyAVfV3
44L9JR/t4gufUwxWmeK4ojBp5N3IC0AhKIJUJYHnzS8u/VCj6utXw1ZkMsaF5lmmv06mK0VpY/c9
Xe0FMjXGhKKycxmcsqa4oyE5IP/ENkqa708SCtTLOZJrmINnxX/Ak4rKnylIBpiJDb5NRVHBtBWK
sc7fYw7VfoaIush20G4B9BmGKX9qrxkFSbPG6smuUAGbVPyQBJynLtIBj6myxDfm7Pewt0xuaYIz
SawNw6C+2/CTSv+rc9q5EFjetwJyeJP1k+/1ThBQZPMki+jpQoCjU4MeH6YSIR+yM+7TwNcxgNjn
v2lY8cgJrg3YowzD3nDB0Rs2D6tjbHoiwIvH6PNsz1Ou9+g5PRWQGKWgIvxbczCmYIWlgV/LlP7j
1XZs5Qv5+A0D5OH2dLDWJjto5yrQ44GEqbMhz/zcZ3uTJRJqC4XCcGwDDx2M+mm5+zPE+2nfIVdA
/o1qA0xp0/ijVSrNsqMrjl7sRIh2/OgiLOaBN+mrYMv40yZ1Q/hGGbdh/qbTff8lAhrlSFg9ZDCT
YcAups5g//tEKhSDsmwnizsbNMIIc3vvdt1PUB9yb7r/+cL3L0CgnpBGme8OEOfbSPV1HY+ciC4c
/GmooxN1/aaHUu/VsqzFNV99/B6t/hPxytgN6MaPmDUoIzunFE0IHHLwA9KKXUxFc2sCLryhnMuO
cDQtKdlzCxfr/+24gsTVvjSzSSShcjW2BaNEs9m3iJm7sW+/cYCvb9mYhYCXPsGMUUkCrGS8yiWw
SxG2pJwnB4/jkb5J9LFtPfi6FuaUYZQaTxcM0pH0oemCO1Oe+PEAAkuHHwymRkfRdo5Jr+DOfyo4
SOMAAhsfx+21Umc2tAzHgbpnR49RArAkYXY8lliKmwP4kAUXhnDMBoVjx3yyCTpNdbnduytYvfSI
CgGnJSh+TTDMXNWr4aRgIcYmtmEQ5ysqWNVJ4z3NQY8aG+acZPAibaHD9wsaVfpeOuwMJgOjmz39
Go9KC4Mff43BvsygMbAxdVP5FrzmOM9Fp8fjU95PyH2Ay/rQmUZ/E9fd1+LW4FaS9KCeRi3YioYm
G13WzhgZEpZo7W9Dm1OK7Y7rxr71ET3rw5Y7ATkzZAgRXAugmr+dW/oEuEzZ69gQvft722AY1JQJ
glhf9e9rXJMSsQ4I6YWvjEWXJzsya6LorrtxOOVuByR2Nca35Gl79PeN2q6oocTRtE7Xml/l0FBU
cHXhPbNnfLK0F3Y+hWTihHX+PNkyW3boRCBZvzVdja9tYCg4mmvi2Fg6zTQHD84UUKiT2dxJNheP
H/MazAN6/SfM7rDNlNw7gGLqukYfZWn2DN/MYYMb0EaMMYK8sgJlcAHNhzxljElpd0vEM9Ggugal
EEgsYJgEn0GM9dMzeG/n2l2IalXxK7tTqwJe+d6nlyQCQ+pnBgW+MQZknU0rBlp+6IBkfQD7qpLg
pBFsF2mLJBjReDfF1SzqYdQ540fjeJDjUhqTQnM44wZz0sm9hzbiUI7aQnHoihQH/Pa7JSgjloa2
MYSbvtBPmyZ0h1a/hyXXrXGoIJNkQvk1tlxWD0c5Mzc/m2CaeGuAArJVAw7/w0jlJs5WAjM2R+Od
CAffWtAwQ+IZcai7ggAnPnOSfzSszDN37nk2f98lB7k2knQJrs8pKprRRGA5aE3pxkKxHwDwX8i3
TT96Cl3dLRfIZZVpbXfjm8pzjd+K5Owdz7Qok6BZNyh4x9NcZmDU/SABOBGL4hQcgOd01VyKIFIM
pmlQPtae0rHovlm4SKA3aZw7ioAyxmR5b/UQ3rP0RC2K+TM2pD600A+4hxPuUQt9/r1+Jclo/TnI
paCp1wR1nZrSB7uBMwHni6MAiHUdC51x2jnSvYUAWm6MjnrXLEtoGYDzz0AXNaQoqEQ+xk+losGB
wTiVgLzouEaJXFdmLvGtqybQucdGrCwFFGcWp6xC2ECd/KPhAgfUDPcUVb8qBAvakpSi8fCQn331
ohS6lzgDPe9X3IaMga95c21dP5yar8UErVqwsu6pu48yK9PKeT4V1ASVcYNCVhJeADNq1r7GRzCB
CcK969BphR49AA7rARJfxlYgZHnqwDf2HohWx099VOAXUGUYln7HXdA19/+iUwNc1j9h9mqiY0+/
M2FonmB8xHibWURzx7jz7Us3Zpi3DN10QUf0fbm1go/10SG6hvAmNYSSRQNfryClfkW0o8yUwgar
bauvkq4s9qfMBtwTTZF4Q+Hht+kjH50xJBkobMBKLAYwLMjdIjqKyg5lFa6KHSJOsK/qVsmfMtyA
niFMd14tF5sbxSvjrUCAWoqwR8ntP/SggEl4fN45caIxtg+CtO/l0LhBhyRFBrViym5/NS/xwUMX
26bptoi1UA1ZNbH0DmtbTWRRq+b/If8ej+mjJ0VuEclqQNDRww/L81JIY0uBDCvEcfHFieeLjoV9
wPQt2vzHc0xZpMnghArlWuCJjrB9aY0wobp8d9U9giWqnseQk+oKT9dVXPh1HJ3vR4ZEhWcv3QMw
mXs775PzCAtlArcLh3MBWJIuO/sMWg3utPCwZgjxlSNw1i1B/vmjpDs7SpSgf1XwpfAqCLWaoZ4V
tfqcBPmAibnrYKXzaQIprRp1DWlxlABoyORVTjck95wQUJ0QTWdxWUqyYL/GrHF2KT7QJ584QvRM
GYFTw5/zyqktw5lheUIVzx/3K6pIBgP1ugd0NlcPvvO9FeqvXo9/E4R1BHy4L4B2jzfgL0HudL/5
riqjKP+gTGn3vwUhAo6GqsiF5sVVnrLWq74naMt3cmR4PiG9aM0i7Wrhl4iEZ8bvNJojbcMGcdcY
89DLUI0WlEgW94oDxGnxcdvp0Nr2Ol3pTunZZjkY83sKAl31sN7o5IhJCgqaRsaEwH4uqvUM5H/F
uEoJfud55q34zZuAJXaMO15oTFoDVRUe5sQA7FzqScMapsYlud4r1Z3/56ERB0EjRp6Q/VuirxXW
4Hfm/TQk+wsXCnO9l0gnBBWEFUBVf0X89j5JVDIZOQu6Hurpqb3qKpajIlFofeHAp3THggpU5n6F
2S8VnWPx2VX2g08UHrXitYLHv8bZNIJtbaiJI2E4VI5vnBIRe0tpRE5ht44n8+hOMtTxVCzLwMWE
ZZykdRJfYsL49TJgMM0aUeAoDb3CCfWvXv1yPx/m1dAyhtc7UGglgrisMgauR03Q9/gU11Sdbikw
Q223tQXGGhI01LFmvi9DqxAy9RmSy3qjMQLwYlQuJSvyFKiU41d3bJeuFkY4lNSQspZmyFNjbfLA
0jnJywCAnCO35QO9SrX8vLGcBPgw57zZBewwBRmVFqsqfPPG6Yg4Y96OqPSRyOIHcZNnKk33qWxl
z07q3smDvsnzLlR3Lgth+3MRPWhMmz1k/bwyQlTVYwd9UHVa04hUStE5aulJboEIlFsFOthgWQqx
jCS3RhEN9++m2ZJZ5u/lkGiB7jr/eEz9nZTErzIgvmynmWBjOXYwyS4++F474x5u1en31W5Qay+a
mxsOuyD/QSfqOKUBI4yiuYPuFI57kZrRknEWbrfi7Ewbz2fdGxu51EQ220caXNdCsx0EcLyX3DEC
TruIEWzO4gmVz0P5LPMTtxpbHF5nvurY24R2/sHvQsXxhnPmNv/gbzT/zCX2BkHoppleWkY53TyL
KU1skQWEC8yUI/tkybJdVGTZBBFVfawYcBNS5sQgvWgacVe8ZyXthJFWoBH2/auIuKPWHoP+ldDY
gppyA/TFpSD7HVqISmbA/TY6DQsveVJBArOIug4TTzJHj4Xt7iaDSUPR7iPpZH0mCB0GV+mmyV+7
/qoa619yxZr6uGyOgMUT7AliomMxnVyotRuEU5npq/cBnPlzPllNFYHlM+rmaBbDz/iCQcgx7YPj
dGp2TJnDKgKe+vkTL4+Z4xshciZAOnxElZFBWBIhOjDOGWLwo52E63kdtBQWaP+/mMl9bZQZQzUJ
9oq+qRlUTye3T9+TjO1Wn6gR9Sr1a+VC8nWhRGj0tcNMfn7x9HTJnSXoIfGb+BFoJQ2a7cRI6uIl
s8vIGUgvw7Y+L/33UJ4K2oM0WRvRT5FurDCtZdTq5NB14op658JzaRzFajZqWxEzLHX3IE3+RAEW
JRls0diYvd3ih5kYCeA59uhGw9204Nyr7g3xQFrCwN2sP6ZP58QivDnlLBC+9fxPSor3g/fSUj0E
U2nufftjz4m5qv4zn6FoWmhE0Y9zbCuyY4BEdlfq8q7xMta31w2Yl/FZLZa6LMixeo/fXti055Ka
gR3l7eyOdhatTPTGRP2g5awVibs/XF/pau2u08hheupuPYML99jDvWZzBm/v4cImvwQgmQDBJSFQ
yQh+EovIbv0G1GjqVybLg3/HAxFPVrdOJ0NL6rveth1HbcbGV8gJ3nQnix9SltEtIXNP/Q24TZJV
sPQuoHwsIsslfpfuBTwUMnKW9xkgHL/kAR+6wMLlZXxt6w8AtoNqgvvWZPTRl7DP8X/YQUZtQBp8
6SXhXSwxiDgnOspMoP84yetcs7+wv32IkFdKcompsTwsNMFPZT+7y8PrAQTRDIAtRQ+l7SwcuSjf
1tl94F+KriFOWgoYe2qBiOXS/P3WSr2pvuPke0TGJlJa041jz98cTbgA0p7kmqbfSu4oB4YV/32e
zJZFacsSu2hEoIw+M6xVF1AwJUdt3hZwUhLZ7v2E3uqk6glDRCvmnXxvou4nEnlDdPsgzwSa3J6s
Cj2EIrEIWXW65L2NJazbUUmxirUWY1UNYxv/JQdGZi3CIMNAKajyqIysaCldGCacXzUbnOpbag5d
MK0UQodFFIHAq+8vqR/891O0TzJmbUWdU6aj50t99LOx/TdnOY2vo3slXP6e3QgsDXY0qskqjYzt
rhYSmagh4El1BUhCAlU192JM5gjCByjHozHHwLDtKxWPRVg8xGeWOjyrj6XY/vKDsWCb1FBHAABV
MxjudiiM7bZt6FmAz4y0pIrXnFJgceiFbcOMoQYO1HoiJtSrWpN7p3ZbEi53CJFO0aEPazGs1ElQ
KdeTIIz4nbtg6wEjwcLnf7ZB1WC0O4RDfIK0xlzIOrHc6gZfWyJs2tVWMias4Flb4kUvCYbyIkDX
kh0mtoPxMejLBwVxhF1GiFodc/Iawu8zcBhwXjyuKdU5Y+61e8ypeVdZ4abrgs/3962qH4G+Zs70
QiMRF+RDpihOtd2jUvuyO5k+5x3gumQ8ffUN11PEIRbs+xgzrL+lj0r1wsej7/rFxySB2nWeOyUH
aZPl3XN/yGQqQYGzTpBnfw+ODtAi+snZRu8rTl2nzVmhs8vjkARXvpj3NYAkaZ8Qf5AyKWSSKN1+
j6Ev+42TR3h2MnMXFY3H7vt1BlLveiZFwFlKHp6ucJDBtidAh9+vLL+zEqUYxbVnZTFDuFv2LwNo
QrcSHCKR4bMk8NDCOnrpWLw4NoMXk6dYgF2r/m6uKetVaSTjk0UKbqPpFR86rjacgAUDjcdBJlqV
QveFpLfxTPEwr40J9BUJAqeXqujzzvhvb0MKmiDRoV+ZzwRrqJXKXON4Ou2BfbzebHjnrPoT5MAf
R6LowJN9Inj95jvNQBSL6UlQLPH6Xxb0Z8KZoR1PxT8f2qGJp0pgNwcaPZMIneuItRd4Cn+JfCs9
4rDVjaNNjkY0JbX7DLxzjV90AglxJYlngn0fHmsDYAWh+sReJ1EsDZgdLS8U1TegV4AyjBrGDCKl
YFe6AfqOPiRi/48ssMb1T+iFTa8YFK4XQ+k70y5BkM4dTyXbVBLpPIWzUz4aEdXRM/POyKwvkx3H
13izm2b+0CZXcc9s0w9Kvx7QtH6dUx5cjQTM/Sm0VV87NIWorRo+JHLo2Ol+S/s8trrDmMWkTC2Z
QcX23k/NKve5CPzco98nx/UmTB7rFBD9Hf91mtWUkWEcWBxmB0zVYSpYnoH6lKKOHKLnKym+qK2n
cPZhLn9l/nf1sYvOfRvOKDr29aIdRhB1Ryzz6P67UTOzWcqczRu8t8ib4QT3mAxa6YhS95jxZgr6
RGrZg4Q9oDhlNzvdTFkJpMhbVQlEkL3TLk0xwwCwKCu+Gi/FEAvzPo0+bVoQtkLgNppKg+jgnkwq
ihffxX+0KjEnshcE3aN4C5/oe4kwLt0JRD8/EO2HnFj1yj9aCIfgpzxDQzkqx7mj+R5mbSKQ9A5d
HhBUFcniMBbNW2lXiq6b7OR6/wYT8M80tNIuYlZaiAHNRmqaFtDjM93ky4W7aZLF4m7OE0Aq4UTr
FnvLe+1iQfmdO5Z9inc7T0KRj3kgZMv+cY/OzLuUv1lkj62rZRjoiPJ6frqIM3h6Orq/hpNX1aOm
+2PnGmyLAW83VrC35xZYuN/y81RwQYPhLNrsIVV2bdW+8ud+0PnBm09cUkqzFaVoQQmktim4noDy
+GQmLT8SWfcWGmOkx3dluNCi24WFG6zggcWVj2TnAA8YRREd7afyozCgAw+4Auy4ofTMRLkLIERl
PHc4qjYPtD7xBY7h7eYLVKbxBORJXn7u6uZoKhaL3NqN9ssXMfUKhfHOTrZCUb6dY96CefW06Lzt
clegNiwVQjfo/UXbniWDn98mftz8vHO2ogC4xy7BzKRsIHslx0DvqwcdWq8u831d8QtebS+CnGNP
w9j5dVg2zM33d7Q+vX45u2XEmho4djbsWrBvaLt9ZGZuqNFWG8xjLMVRSZ3qNTA9EBbjx5TieoED
vAjqxdBgbXOJ23s6AsPhPnBgCEWX/tcIC29KIm1NWyibDm2UQeWXrBvJq0WPpQqBYJnwMhRNB5cX
zdaACzubnH6wXBcUM7Ih9DMZkaPEG4A6Qm6/4ypZrrdMix/ooXghq74hlpYoVYCZ8ilcjWRznebW
1WwXW+Ynzn1BhUjf534ApVD+yYscS+BaDMeFtfxULLcmio4iX1x+e9f7P5S77dSP6A5W8atrxqwx
SZnZ7/BHMAyH1qznzP2+fiqkHyfAXrBkp6SqbR1AJbYlHEakvQEQeFnPun/5Z7BpVob4rOhq6xxm
WM1g/m/Q0iKbLgL6RJI5+z5V6pbtO25cyRb3EMtZQCdMDqvrFvo3lyg36zV2BMs3J7eUOfGVrSm3
93tiTIbzHSiFRbSGhfC/k1XBE6SHesSdqbJTITGBAfUuv/n2YOeTUOyOFOHsniaVPcGXnRF7kAHR
3OzSOnu39X0+0APyPzNzdVYhbp28u3bz4X/7lT9bQ1gRwprm5LmdFKC4sWTZQf34ERSmw26kxKbK
V115MZXHpkWNJrS+mob+0gzzCi5tO1FK46IWQ3lLqRtqC2H90aNxDmRyC03WRAI6Wf0mKDPCrMmr
h6e8sQgbfl0Z+A4g0xJXU87TME5IQ2vu5T8grhk1kc+6j9DuJdT/e1zmU2pt0Fpc/oVkDCUXsW4g
qbCU5smG38rQDTNziZ7eUaThGTcy+bZwsdxTcKB5MHsfC0uIxXbNSZVwbCX5s/0LBvMYWMp0A3yo
J/UyPKKl3mSVVKuYcnLrL6Il9ZJO9Hr/GTAimT+UM2qA3FWQE6UYH/ThRyrwO43RJS948s+KuqLI
WMl6rFJFdpr+uhcdeHrXtwybs/x88K7XPnpwNnuZt+aJbSejUs1MlpkmwWl68+X7F7zeOPoyIqOt
3h9T2QKtll80tGcczVTaqgSwhFKLcwpsFeyTBgZitXbDajlLOj22SKqjE5mv66pRy47w5Dj+Hg7n
IxaMUHKHJwJnmXEhwAcHsWWpPvv81UzxS4PQ/6/b1M/4vsq1NFrN/a/GumlaJDUxWCCK8CkzM8I+
IgToi6xh0IZEdCXC4JnmFlWFH2nMcYPaunYWJ0GekzBbPsNYMZH6zNkV/SHWD0kaOCXhU0Sl56E9
TLYjb1ggnbIUlW72vTUNHCSuHk2GRLFa4Qq7PjWoBZOLQZME9xtt1sYvieV2NEyiM3BaTL4SnD0/
7wcsr0SNxVKA0RjsxdZqrPXI+boRew6BASiNSqXNZSExY6KZgUKrO9LuyFyRd5OjwCQA+cZV3/Oy
Fvskt5+Cryovn+CKDFXODMwZsPHVj03iQ8MVUuvbeg1gvDFbT5dQw4m8PwxZqDb0Al/49pDHst8Z
5GFH8y1+hbQFpH0ShFVqiYfVSIOx0p8puFHKYwVOseSVUyjr6EylHioyLsgfAz7kc1BbN5CMNQo+
ktbRGbSDABt9EZP2zgXtM5MrdPCUK7QSyU38hRHul++/TX/0RB/r3HIz2EXBUpDDKgTmLBOSlRvs
sPI2Bfb5T7ttCGzLXSLP8pqldf83zGsOV9NTjfYtZEinWDj0xt/6JaePnhGal0XMTX3oOAINDDBv
CmUWmT3ZeXa1qK0mer2iYydDI2D0VUxtsESsc2Sl6DsQ0/M6S0q6kVi73mNgMIbcwgo17svqi5Ly
cW/8a9AiXT2AklgvbbW4utLqmU8rfkKbPuiIk7aP6OBGG8FWk21igwu8PlJqhuo0R/HyhqgAFz7F
BC/wOGf8uIUG8kW/Yjqmi7FFFdR+WIuRbK4pJG6fPaTDJIdsnHFPd0tuOPoEAh6nfHE6F5r9SVdn
zRGr8gG03lmXVS83lNF93hLdPLnO6uZE6IZHkBfAF9LQKuarMkinDUszRNC4isRnO3yAGgMQZn6u
nvfzzrwDTleIXQi4789sU1SBp8Gl2Sh5DnAA6LNcR8kYW2FECXSuUQdV9fQdYFiJ+FmyyG3MTG1e
S6rth1AKebSTUpf27QoG2DgI7N7qw/6u+HVL9TOhM7DqkKWxYR4R/blENki+aoGf405kgJkqIX6L
a6/ydvHdpY8QMcKcy1aqnklwpwFDOMKmo5fYiIEvv/U08i+TD9GMFk1nY65t78r0cRL0QDnbWb07
45z/ivKq1djgFn6z/dO2fWthTXafXF//SMWwJ52z3Mxo47EvDUr6wTOYG/FbG2Nlt5L4KRTHMZEO
4o1oJ7vGQnVada8vS2sYJI1cofioc1rtIGt7MmxuSA6X/segKuWChcEqz39uy1lcPO5pTijeXAgo
dBrqJXCdr9tdLxUVFTpMDx3NLy6nGTMNLRudycRCoiqjQieW8C4rWjQnkOYJ2IHmi71S9/E4WjKf
iMiY9HtJpVT+6XGlyYDuahKZgng3mEVu5IwKVipyFW6XhzaJwMUIwW+VQMh5x6/4+R3BizEjz6pt
PYiAP7T6V8W+PFfpyCV49xD/IxuOSXgvudXfhaCeFn3eUOuzQdOf2faMKjl3vOrSpAC5t/vdTHDc
T7npKOcbiylFG4VB0hLBow4OK+R9r8pallNVh7UZH1JeGnUX5cp9pDtnH3q8gh2bh4Au3B/VhT6S
Cwm5LMHPyNDEojfWw4iyqQBNGF5TNqv6Xq0J0nDMcxaPg9QYpz2DA7Vf2Jh+hnvTu3x1X0/mO+5d
IqyST21kMiLKza0HzgMGOubKwWEwfI0WDu31rNdW6XFCm91fNnR9oUwj+TZZfM+u7uq+esix1wyr
EcFBPIhEEDZk3mPmP8//0+qp/luuCPb7diUDiGjtmecN1t+Xww0P3JAxvHhZihLa2breF1oxcB8d
iWjqYQ015ZwWpLUa4TkJaIAs7LZzLvdFztOiHtKSqVm2RoPijAf1dawAmIZCchRl+knmU+xIkes0
5gOU+wT3ufzUpyMzMUod5lWAotf2d0/rAN/XmzGVDbLc5pCOjsNHd0P9Wrb9q9op94oO95EmuaJQ
EKIhrR9fS61bWEskBGTKdfEaKRT/erQzXDh9yS+e+ssXHjXsRVNy4AIwqP5/n6T3r2/T+t2oxHB+
2R82icugYTFd8z30kLXkhT1b3bY8sLcwlvTKiH9u2Y1WYV7J4L+wS8bzbotGPqc6fYVd3suAwcQ+
YfhrBi+o08FI3Q4lj/xMGArIxlPBfWfCUP/ZaC6xhPLNUQU449PHFrzMVihb7hl+6VpP5XdDDvz2
7h7XB1jheDXdxmI/tI60izti57zUkZShaTi7rku8oUUAJSh68ffdLk22sBSgdIOb6UBUn5bh6p0+
NAyyH08Qw7bbr93cog5cvRIaiJbjynEfBqYEi55eAEsmHgTs4xSMl0Hq8VS0Gynm5604txj5qJ9u
kTXeyGtQxYCVJOkrowkKUZsK5LifM/SLP3n3NRiB1WifMqzZm6yfAXVf6YbcSZxcqI5LMG/OtHLk
nWSOlvogNJ11OMw6DDQX4WRVVF7EpFcaGzREK5KwQ3+boNPQVc8kL1cxDbauQ+V2srGgVgpYnfE5
3KYgw/TuYAWWnC7/o2wRE0JEDHYLUJShhdqElQaTgE736VNQw85UdmJHHshfe4nAodkrM/3ETXtS
uPQSMRQS2GXrxSyw28jbHzSEZsEJ7cTcZJeYQwqKUgYGAnl8PYCqnLQrURkqvd7Xk/hgG31nMoQy
FyvyKCFKqJlEa8m7JvDscZDIKK7tBM91h8Tj3AWd9hylG4HgrpU59LxzVZ/7Cj44aeTCGAt2PIaT
F5efAWhgwcP9ivjWNRLtHFhFu5LU0gfQ3X1tsi2jVceGEZ/wr+tjufEjaf/Jkq+q3q5w9m4KWiRQ
dqSInmZzJPKomnUtsbO1NFNoNVxqj391RPfUBHNnyC+jx+KE6Du98Nj1YwfwfhsNqowCZV9/aY4u
G3db4c3UkhlYgCbXQlZ9dM/mZZYp7OmSjOEQYaXPF5qERyXcfkbOLseqaKIkPKzpA/so5kw5mHIr
QUFmrT5jPFmKKyFs7re51YXduLqY817ay+OFY4oHUcmiVOFYGm6DBHYr4n+wDo0Pq3sScZAA/Rto
CIqPsZZ0GJkJn9blVptGNTEAU0Yf3laPwJnP4cIHppTqbtjA9gubADWs0BJEwC6ltludLLGTPp7w
nvAwWUpcLvrHNRyR9ym8kAOovvkMckizKMJxvV7M0aFZX2Ys8s+9dSto+Qz4rozC6DTsxlgCrMw3
opSi6upyZCRc/JCtg1TVkCyLqKvhyFHKu95n5mRcrsbWuFdINRJJ5yZ1qNank4Ae7gauQZKEQ3qa
/yveIGt6c/M7nWE4eBy7kCjsxe6Y62HIqs+Pg+ItB5Ta3phM0qFfzXGX8YL5ogbTmRekk3BObshD
rDHbL/iruMLhgcal/75zNxeQWOMSxPl9KcourbvXuUEci+5wX4e0pJeUxNXb4CL9MG/4aMsVU+6L
VUZlzN0ChpM0e9eid6xobE7PnGeAji2qaMUO3muO/r78fFXLdUeAs7bxFj3vP0N0HFCcPemMbcAn
YJYVZHc+nnI03gUUEksLX0e+oY9a/MB9Bu+CKMFKH56ergUmFLj9Vh0SE419i1mVi8TviSLJ4Cvl
3TVVZyiodQAm+fEIhCqImka+jehcATU2u61H5wc8OXKeHnw8DF4xqMTbbkW9EZmd3cdEK/6zXG7b
xRC2jfpqnsNpcvs0jT+Kce77sTLKdCjh6vl/fx95yxT0gIGzGOc63sWC5SZiLmqLChQ3GgwWx1AM
Q6SF0gXNfRWk6EiXq+Axqe3iQeq1WNzpP4wBktezcnY0wcFGRMQsWJyDm7DXaLPowDj5QURYz2V0
SiifDsoR3BGLmfENfBqrDbXXwLpgpJXprW29SmKgmBuluQUzJtwqwYe4LIS4cCKTzaDfFD9gsgyo
dIWIwpTGLQTBNQHjaAHCBE/2WtnN9Uaul2+Aa/AI9e7zJfjwQI/YbAc7ShDYdNR5eUuzamZONQuA
EeyxUBVO1eOSEYNKhngxtlknGwz5xzV9xlcNE8MEj4oep2d5Gk2xYt8pOvoRoCNrDyVcSHsk2if5
FWhN3EkG4tSTrQfpW86V53K/1lp4+80XFHnUOJEmvpHD6Jad02Mw3GIAEaKGmM2RdTSaqpGJb6w7
HIwbSYe9O+W4ikN9Cp6IONqdYNTyz/ZB6kA7nmudO7noQ4zNB/RBJ3PTVfkl9MZF5xiHkRF0xGUp
GsQPNiP53+7zN16GlrM6WIehvpqWS4psntaC78VIfp9lSXAFZfLTqATB6d8lDy5HzilnR4IP4Dr4
wuN6Huh7FgYYhvxJl6RiXJ0jKq8X53H1E97BZ0GTSH9ChXBxUz9PfCiFH3gV67WRp1mqgLxdqhUG
lbhFR/8ODfyfZIgMFCRBY3Kv44k25Z50AJROBCyAm/S7dLD2eH2p2nMbzA3N3kv+zi5eycPFEFRV
VN62ERothRN3MdXmNZ2X6LB9qkMjZDZzfTNgBnwy8K53jP3QcIwIql6yrjwHN6qSJEBO8l6Vujm7
sg4F1JULjPJgkAvOCSWePB5KDQjatoXoymQboK/a0ap0eCFyBPUO+rLh/b7q1id8GkE69M28+73Q
ZgPAzoIfKkZ7tOkwwcrNASH5AIOqWdLPRxt0jeNobtbJfqr1uE1FUe1raTOv8Vb6c0Axt46lysNY
ij0M9DeyTooxcWUdFziVtH1ZOrItOECTO5qNk1UNvMWU2Fe4POR5PVmG8uYTYny3nyGMqDanLJIX
dISMVDk6QgXYa4V7HwsE3ywbyyK46roH5HLYogzXEe3MwDCWvW8Vqm8vzyd9tY73RI0M+XZRJTeR
Vb4+5oJ9On49dpnKVffay5E03dG/VvMnWNP5rWlvTtSlQbovVq4mZiDt5N2q7oV6yquOtioYgbtl
tidjEuaUAKqZkBqyb6ysrPSV+TvhyJssvKdZQCHlaD2IjfwmphoAXvtuySuDZYQxivbt8u2lNmCd
7dr5gxx6I2Lq09Tmr8/ds+K7RZ/74ZS52hxAmOUPGmrN7MHSu5js1KwDypyJ1exMIrDX2ppvpAm/
jXs6GvNwO91e8BARIQx/XAsenknzEdW1AeRXickGUwn+AOdLYqk450pn7AxZvnNWdtwLfr4RmGvF
837HoebtwOxM7uHkNoTq8rBlTm6+fh67k/p3hVYwQ4uZO7rn8NCZk6vE7cy7sWxGQS5DsYkCiynK
zSqbyYrPJ5wUZyC1R4rlIiy88ZZElsqd1zTfmGTv1HflPE13UfP2wLOCfgwq/51seZ5AusOxhHuh
5QDW5jUWy4+ki/s2vfcn9xS9n64tqlBLfbK4/sFe5bxpG12YJ7+esdkYYGlM3mEWN64DqKi5B5Fs
Qm1i5tSVJfmVg28A1EEnRsM/XzbxOZjep6T3fypN/6fB8qMoARhWoFFaYvQPkcn+wo4gP0mmegvI
mPKvKP4AOFFl22LGcUi9Sy/e37L5B60tDw9aTzEgYwI+FLz4cO1uLOHY+zA65sqDVc8aJs9CIQ/Q
3W4emqS0awbxi52o7WeS9vtza+L6w/KFWRfMRdfwkuzcZ27Wc9/a1CF5cCrmO1/+fJ84BnXpiUfw
6gQvBuUDCzDUgd5ddtvFbEJgEr/BgIG56p2eGa1T1bIF3wo/lxii0oedliuGowiTrlsPfxphSm4L
oRO3YIdK+luIi4Q5SyC2TcEkA7pdbQrqrFbJv2/ALI03kNHmWC9tQd/AbDA+/obCIO4A57ySmm+v
K28NrXWIxBj9jKnCwNZEngXzEDW6DlbFV7MqCQBQPX4b1SMEiZMvJzAvp9ASeObqzhseEN2JyxwL
zIZnBqXij9jMmaUmAyNha1pj8QAsrd1DDOnTVSVuqBhnsIgzGJEpQc0wmrab4Cwk0AtA7dvsSTfD
wNl/wpCMkoFpenvRaaM5vgGgo+H42fAIXbqWShjJBLxXZiqU6BtAxhJO5D4eSNQp6kzbK5szp5Hp
Sw5XwZ/FsEhkGq2ciFVjwkW3ZhvzHjYQ8mQfjQdEx9j1H+mwYFKab60Do2nhmN0JfvV9W1GHPDur
wjJI49Y8dI03uT7QDW8wU3tEbPWVx2X2ETRlKtkXiUxDUdeA0JHPvXqq6iOkc7lNchBHsxPkvL98
Xyg7Kbx5yXvX+D+ygosxAUyP0qoJaIX/XsSOeQDSJTEwMBzT1LK0UAR+l/A3bZnfVBlM59o60jp5
MSlI7qSk1y2In+IjHXjP8SdPqMKE1hpJun0bfeyOx1oiQl2YnFhWlriAvgxwWsHmCxzSNmxSHbY1
Wf6fmG5CdOWjYVc6BDnEiKpCsZpYxd/8VhcndgLd2OECc1tSJCXGXDOr7Pp2LiRZsH5PAvONv9v3
7fS1RZyQFlCV4bfQifWRp1Fb6A7Tjzxcsu2I11c5PqCh3AUexSIUVyZ9xYCzPsQH4jkUrJ6QBKJ2
nsitTGANwGqgPA0GalVgIa6AwRzUFcE+4avuly+cgJZr333QX6buu4js5GpTnRHly84HH0zlpaG4
dz2lRM5r/d19Em0/ab5b2xBtDZSP3HGtpzPtan+jkbOMGBZfme7KZM8hU+dE7iaYksqTAmU7buLr
8FTet1BdCJ0OdioLTQb0pdc3jiFZQtxdX7DOx7pUtG4WtVS7Us5vZgKnpMlSbwt+GczcMt5K3Ai6
r0TKJxNW+XK2G1qX75FRdvwuXHTr42ykEqq/CbQjwkyvbmVj53D/ppWQivaCLyy4XLvOrcpuLvtJ
nSFvhF4i/vzvm/EWnTkR2CoUBsMQyJAHy0C1apYL2y5KtHermBtwsvgKW6SXJFbOw3bKGI3H0oc7
sSwYt2YZkgU8GYgNjSLZsbfWh6Y8xAkEGzAF0oAOyELF3e04vxERIaNj6s700n54g/mR3E3NhZLZ
SigaHcmtCFM73sTKK/qK2b83/nfTHrKBIVNXawI/Up3Zuj1TawE8VXej/gESGU7em9ZKWkOnzthx
igsY5/rfqcvmxnpuV2Y1EfHYda+R+pldNBYUEDmnlGkaFYXcYna6j4ghUr5qnRLr0WA+DS1q4S40
XdQijr+fArIXxzHhoNKXZLWcDTbolxajqlnWI+22xwGGWZwhh+P9YThsabDCuyjYnZ6IJaJfef4x
BMOUmUJuQ4vSwsyt7jG2k6R6mYDothzY6/jsYDAleBzJ7ouGJ9kCm6SUQST6O9D1KbbK32s0NFEl
NcW2JUGEXs4Pow57GuokYmp0HrbnfVNMHMBV3GEhOnWvu4IckU0aPNjJzpC3qRpbzDyvLgSwf1v3
rst0iDQPmo+QChCHatKOwKJJzDE4mCrZnu6S+RgYnZnHy2E6KS6KZeX5EBQ6FcWUQkz4Qq5A4hkm
Ccp4k1sz/JlrnGKLv28ivdoFutHDyeUaxqJIEwxa3Fe7WO4wb6dZEZn0KUFNkkLd2fNEmY142U1k
2B3g4M8d32wOFkqoKC5hBJcp1QEJ4HAlOFilgvpkLPN6fuZUzU+8GWw7i5vI3bXzOr0Oc/g5RL8A
lgbkWPU9sI28Eo+N6SiO8GdMe44vsaKU5zNzv5LLWjimalyYfIt8rzcwO0qfANRwhKjMeS3GVXom
D1oOGHg7l1IGpDRwnnd/CWpx0bNoYLHqSe5cIaZKZg4NK9/vFLf80rkaGVAB4Dg2ssrWsMp/yuIf
CT8wRnzToD3yHjG0o+IhFN65tdzTrpFkb/qd351Q2ngxExUR+YzqkDohln/6M6Z/kN2qobsf4+mn
cXu9wj8GzhcSkap4rfuWf7XIuunPX5byH58kwu33J6IQdxG8jcxqHzJyw3ZILxaHMkn4DrtRpZIK
FQ5NtelB9NP+2XPELV9ESxcNGRI7TQAYXA54VOHc2dDqP2hMPJsH7Sc27oW9cUV6uMYxdEVBFFwg
pCiSM15j9XC/Xti4ivQt95RGT/2tP1T+Fpc7j6kWCmV3kW7mvmFP5yjam4EmKK1wBnsvR6QJI6oM
5AhSNRfmdiKuuDpew70RCux/A/mBQcnBTkRrOKZHuhD2enSX7jYFvgHWuJRs/uT/Dj/f7mQUH2rH
zeJ+uHEaq1D7QJZzP5yxeUB2UuEelZR36eQXTtqKZkWpVZjcyZgXZpYYza78aX/1FE1X8HwyKVGe
zEu9A+Vc7wK1qRJWnRPkwJfXBNPLFzHVaSZfLRgKVaiDJ0c2piN1JFo3qFriy+0YNFO/e8LBUMHM
8gF7xqPxPGCdbTqILICwscGLQXhrizGA7eHoH9yStmZa7tKzu6u/p+h0LGnWxRX9sEtPZsqmOOur
Mi9nupovTQV5ZZNmDSFjPAGuyP9v3rJowQZNIEJFhTidZ16fT7DfqsyXoR9DK69rs3wSuUYotCD/
pkd34XQBo+dWwknUao/fa3q0u6rAwZ6TONin37CFrtWIR+6PAiMfq0XKuUOyEqoGqpF8inCAm0Vv
gclyyhknMJ2DrflAvtZuIwYQZWSQm9dCNAYSEm+CNEJoJuZl59OK12KNXH54jIW9Qd/t9z2YTtQc
uf29HsocnUixE+jTHWjn9KzyF+8qbx2Jlg6jkyvmRxoojd+ZzUfVcl/FcAA0g3HHAOYmgJmmGr6W
O3cxzC3D5P98r20FxPR8O42Y/JkedJb2dYrmacX/KcMY6+hCCSJv8eooX+bb46dhIx23h7ScCUGY
RxCB0aYSG0yVDd+sviLf8z1iMOMNz4NDjFLkITnGKcElMlcU7vMjHL7f5DO7F5ZKOV7v8Uob69zF
UeVVz90w+4sQTFetaQGGtEcmg1D5nngL3NQQ5JkYY7VmxFswtImV85Ya2WKK2PYUIHEgYjy4mIlg
tYoCxgayDChvf2dn4555UBPdTojsrl5Q6MBx6FxOuwdnH7pvPQmpCbDHFPtiEKc4vHA0Yc/VJesF
fC8UCmj0I4t9kUNZp9oG8L1vxF+2P5JgPeVWSNGTAIOWZa4jsMKHQLmeaRdhi0BLd7ouQptsZt/1
aGtj74uDxqBfcktEMeK+rOH+JT7ay/AaXa1ym2vKehL7EAzuQLDX+/MeYPAJNvqY39rZUoSw8bI0
VnpANFu1K0YygoTf2Jz+YtBmrPCdilPprmJOBKDlcch7CzPzhrsMRNZQ9W3o7qXJtKgiBu8JDxWQ
tlQE9mIGTwrhKcr8g9CctVESAF11Rl7CMFO9inuJM9YY6kfcbfGJ1TXFIEilUNt7x1E4p+sUalmY
NOZSTrovJJMaoq3QmN30EyJGJz2GDPcaikpQaEfxMUIk0e3+0/cUQjB0Y/HYWPyayMGbHh4M0SdR
wOE3nNtlwpHI0rFPwKEhI8iZmamJuwpohhxRXTQXhcoSlDxtAE5/wUG79U0PDASFpIP20WaU4+JC
V6fqxZhNSwzes9f/AgauPzWWWwACEGL34JWj9eV/dzMKtUoNFE9C6oDuNrlkgwxjeA2ytzeVnuGa
pc+gOtMiYBAWLGhfViDsB9VqwfXrf1iahU0Ose+o2oQQpYnNmda01Uy2S8zsf32z2N5pJuZcy0gq
NT9veW2ripfcIThhQtqdj/YtoWvtdX4VKs0wFNeh8skJqhRGL/Pw70DyoeAZSF6C6b4Q92yInq+j
R3hKFpBlkQESyjhl9E3lCoPsOk4GIiZZjm6aLzROY4ONHH+Gfy3ct5RnwnglHbkbFMV0eczE8buK
3vlc73pYNfV3A+G6OyRfV1br5327r54Q9+dsqq6ijE/IY7HMekeNWauWjP8ZbPquO74bAQYH3gVK
vhr5Fd72IhbHOzcJRQR/XHZqkydhhWnqrCPvE64teupCWUSjCCMHiLPzBz3XZEwK9RkfoVU9+ndw
inQkfiibfWB59z3btrkTfPu3ppK29kE0e1BsG18Ecw8mr/oxF0VL9Twh9umtR7D5osoDA8lmPCZ0
RTqZknvYtF1FjfoiY9u5ge5tQ6WAga5PyOoUVAnZIniFWsv/EixlXzQ+YkmTZmztF1wT0p22Wi7/
8E/IiBmSjqW6eXMdZ0Ffr5WaI/nxb+6THdZkl5PCBMEoc9sia8K1yoKLYpHV4waro1USo7TH1Woy
cwcNLV0lmv203lMqKqJc/4uyBmzw2gSpLWbNKNBMywD8gfUp17P6iy5gua5ihlG1w8WdkVkYPxAQ
2i4Qsgw2Sun+415UFJsbCQEm7W81C3wONRYxcfxl9EaFzsNsDXiWX4tf10VKtIQtw6kqKfMNoG3N
y/kT+zPh/zMilGeImjssd7HIw08iL+dZFGwCylJ3KcplOATVsq2qTgvO1LkbHT1XVxsb16IkZY1c
cHSIViwKEQyHbPgYTu6p/b6VKdRvCz60CWWyZkKRF/UbSbDaDOlD4rhbI5J/qney9jRYdwnc+Gak
RbVaoFGtmtpz076nBctHxdIoQ0X6ZUM6ji83VQOFGVFrKF/a3TUHGlDtPs0wzicExRRzlMAa0fO8
+TlubypDODjBm50jV9CKqKhXkp4+lIZVFw7OQHBEXHeQAl5ScThfDzBqSV/h5rjQ6P5453TuZAAB
eSp63cJyEnYrVxGSLuwMLJ/EhWclGlR6zJ3VLAyOFJ1aOaaNrD1eXL0ujk3+RVNQum6XGeW/BGoD
MRdGrtnXqZY9KUvSbniBqd59LLwrKsUDGlIAvqXW9+KvJ3sdZ0tMWWFPxSHN6CPF4gALuh7E8S3C
3nv/0C2MGREjw5B9us7Pg0XVT6JLok/Ljb30USKdBYTjohdEUIzaJYARiuvvQmVz/T3ZD9rP6hoZ
hgmRpv7nq0ObGp8OthhZ4tDUdgv1OnmefQ6wYIiqtISXYTGrhPDPWZNMGC/P2JVVCc975hS7yEIG
fIXkkmiD/AnjK2jKlT6JYSvwlUvD2489sVWh/QaNbH9fqzoRE2xJC1IhC4AKCIELFoSXDwGJ7wc/
3NvfxP5P9KovSuFMGfiWQ2X0QSOVK2Y+mn4NG6inTbGtQrWuMWS6dfHghvZD+4OKQzmP8mMTSZoW
eJGNF6dyIvffxkrUVNdvF+P2EC1gdegCZZJpZGAspC8/CvVCbu2M3jiv5K/KLynZuvwiaX32xfot
0ACjt5vLFHKHbJpK6QjnWMalWLraJh1OcVrhJvtjn+oqK07xPBylI/ky2H6iXg1r+Zlcs44gubh3
iDcyXmjGfA7nx6QGSVkkPDHfeGCbmgNdzHkUDL88EsY8ydidEiSZDiivmbgUth1zuQYBOZa7hfxe
nMjUrpbNGTvprpexyUMfG8HeiUacm5MoA+lRhj9kCfzkqUi4ORVjmYh8xuJCKp4wovMBUtkspeLg
MOQkKN1zU0gD6ma4CK5gQeP3jTGBCgTUA3sbVb71FkthyMaVruzffIwuIhxpjvN7UgJdurla/SEX
OmOg+wD76FKnGaIbEZ2eM0mRbXnNSSv5E+DkTQNrlR/inHE+U4hkDoDzBPh3MgbOSnQnLyTnBNCx
7aMEMX0oEyHYUJbztgVYsh0SaNeEk/5wAns2mdpb9MAG7dCXkfpPapV1eTdelEP+twmcMDi8tnpZ
LaYSgRnsg4Qb48YHowX3fPp0rQdXHuVca+5SWc0/192TxHLEzEV8ESH9IzEwZtxgsPJx0fBNLd52
7yLy80Im8Qv1BMUVNgVrglZroccPY7w0J4ebmYp3xPhV6/wW59VtOSedrwIGhKtvZzaCC8tIv8kH
sYAPeRtuDn43cdDZ0ZBQ+i7KcQqVWdPHXO1+k+tRWWo3WGB/kxIyAfUUdZKRMG/TgNOCBhp4lijY
CFgMH84tVRm5WM9tQWrKueJpwDFYYPjGxHRzIeKedGAePxqkR3iA7Irt9eHEiqWcPl7TfxC3tbuc
irHERTqEEtcDuIvQH1Ucqtj00GW0880cuDIYQ7vS3/waLge3dxb30T9Nfy8tgkCnHhlgvdHgzit6
sQkAViRhNWMPvpbo3QkldGGdRiAxMl3BNg/dMEXn39CXJi9OjzNMgilm57VXmznARSX4/BaVGCiA
0j5mzKoS/sNl3ITdTnX8mcdvlSguaLBPzoNU7Ot+WABYCbHWJBqb3VG0MO1B/TBAv9lEEw1mLhWs
6Q3WSOGGmDvOADGnmeG2uPhlhdFserINg/wtT3hLOQO72AIOdYytrkhrEdklCCla8Es6lL7/W3MY
4cnBMV3HkMr7MFVd/TbMS2l3mtCjRhTCEtr/1iq2PBVHyCXNTLcKj1fjr8+Cb+fCTQ5a5pSmHERi
OAk9sOABSbyANh1JzwmGsq96OwmqEEbdex7IvViiEokZib55XfdBKB/IyCXR4gx/GtvKxbnLp8yE
TIWulpUeO9fL50Byyu0M6atAoqQxwPCb9o/HpEmBC/XWaT9/DytR9uBdRduahzepqnXlvYarqabZ
IP//EaeucBGJ9MpEAtuKfi+42jhiWgKs0zIrPZ/m0+vHNWV3xa2qtMoKtvU6ISbF2JlVrTp5OnUl
QxequGaodXeZJ+SlpA/xjmpnVE9IUKYbUI6Qo7hjw03y0VvXeJ9lcp6KL0/qMq1UVUNECrzcaYKK
5NR97qzzwGL/97ipcLoS8GByMZQtRlXivyk//mXRtMO5dZpLnYxeksYYBwUGvuVspFX04gDqpWWX
QoTr6/OJDmWTuOyDrrEon0QTlSXzoaf/KD2a7LcFU/opkzVbiiRKFFf97zWXvgEwX2CWj5peQpn6
CF8HO8j9tzfHC9mN1XZBaS3jAJkNeZsl+eSZx7A3CUgMdfxQhPCynKUFi2i+TI5C+JxslhKje3ZE
grmORPrvKXDrJ4m2BgHCVgrzfO7P36MeICWaPurG0Tc1U0A2nOkB3hZFom6ZlREZCAETrvtbqWma
C1mCMovNTS9PoPfki2xif17qRbt8kwOiSqZY8TH8p4MziC4mBEIIpwJNMqDRsNaYuJnbYAgKNPBD
N3DWN1EopHT4r+EWxj/kjTdFs5oEmkMUwWvaZJm3yIBKLsU/RnY+PRgeJ/JQiFMBQiKKzERy/gmu
h9ziDz3AWgNhZEWgDUyPw36QlGJr6lK3tVElV33J+JKI54h1dBaoQWcei+KyOXoFQJjS+66IksGY
1FpfVFLavNf4QVa3Y8U2g34ttv+uSiq95vOSy4AjrMR5Q+FtiDnfXjWdaJA7TXA5YuopuY6mnblv
qBXP6yIwYLiguu+LOYeRFO8uNmilxgZ89pModvxk12QbZoI5tJDpbP50Upvrvm8RseTyWxbuaTc+
SsvsvQo1rZv1tiZ0gtIt1kuLkCqKfG5pl16/EnwE/tQm4d4G0zUJNUgF0NBKXGHovmAH/eRqTahC
22/xUmMCTPvEqyr67OCw2FbXwWODgK66yojp7YKHpDEg70kHaf50qek8PQ5/vuZd/HVqz0hu6pry
q8wevrps+TPpNP3Wpi2hbmwEyOJEFheQlv3UDgnpMdXIE4mpay3ia1965/m/PZCCGOJ09blATsID
PmTnZbiKukPcayL3P38cMvOZIqO+XBn4NL8YSRRBu9Zh3Z0meUp80cYJIO9SiihegV/E55499BOQ
/n5dy0oYkMaIjI50IZMDCfSu4V/0fqRf+UdrGk5iWvEPal11QTCVDixV+aY3hIFwQJRx5RvPVu+n
VN03b5bYvFA3PPqAJk3/Fd9CTK+o75LMHgZIOVSn6WDtrdohaG7KXq74qlSz9iNrWtVkpfF82Xsf
9GQrNXarL9fEAPbEss9Jr9j5s33U2I0ixPuH3Es/9DJZu6IfVEZU16ji8ZUdz4aDNo34OafHX/CI
KMoPdSGMA6o1NTRFntZVBnMT4R+Q1s9TK2CJjNyEgwxjqhIoCvoM0kGQ/8iV2wKrSVSwOCwkeKSZ
FVg3J1/pKABQiZx8EeVwwPwFuO+zEnD8thxiB7as1WnceV/xQ+BVf57O/xZCX0Rhzu5r6YnBLSO9
zMq1ZUjBlS7432+T1+SE4v/8/JbgTO0nPNERsV1XY3dsccpNFXU6vKx+mIkZ0Qv3vmiDThlnIM/B
IofYxaOo6oAo84BiLMj+iGRIgfgaoHaVvvKChKkDWSTceT9ApqV7sJR+Zekrp7t9GO0DNkDwQyaN
a+z1kU5kwOz0xqMG1WVxdoM6wF/UHhIV0tELsZRa1n3eyqGHtnj9OU1tJFThc3n3/g2mRZXkoQ1V
kNJ3LZ5IJn3jTSsbSeU7V9x6rJl+0RPcTsU7qEvBofoUqnyNaR4deERrTC8QlrdZEA8x9YT6DFc2
UJZOSWkkeYABM6TpVj3Z77sLqSDBFduVX7D5Vb9OkjZ6zj7mEM8XWWuvDT5zmuZm8SI8E+iuuJlT
/NcS7B7PoWa8iTM0SbiQe2ATtM8id7m9bPB4TCTJ7VrvL3cgBgEeBFdP5FB2lXY2kM7uLMNdh3HN
GUtad9V6KS2cKSo1M03NJHjLcZhddEzegeROn8jYdVvlrvmWjAkTdpoOaip3a9RgiEDb3qera23L
eQdA/WPGOlmG65e3NXBkhRrzURpgxS7eb7cJMJC5y4LNZ9PSr/L8MQkvS2VgLpA6EycTyGJfFDX5
naOqNEs5MxLsn8A3jjU5OlOQ5ajAZSB7zckeASoPKOSnyTMqJwmk+T/+Ux5+ylzTt41zAqalV+Vl
0uWeTfMT35DdQQWxYXEduBz+3469xDgkymVUxISfXDsEWbzhMPMQWTSpopsQjvUlM9rh5doniMf/
nBMdx/IZv0cfZvYBBriZa9PTYqD4w9AoIMlG+sZV6ilMOjdFXutjJHk5NmhU5bbv64KwiBPOfqqz
3nJMLjSG3CSgw3okKSmPK/IrLY5zD548TqVJFxoJ7UfQl4mfx4dvkPJiE8t5bO+NNVNaYwkVcrN+
RFgz8koQfD43TrMtFJI1wBU1B1E82ys5TkTInQonafTdPvgG1jEKO428duu0rAhXTBqdycHrRuVe
4iNlrq7ScJ3Ek6WYxEDd8522BzgIUkuyCJf3lbxrdaLMMzfmlOB8N51ns5zp5kRMZLw3n/A0l9KP
o4cxPfweKMx8PEK60idFxX5DzvAEpyXWOImP6pq2iEo7jWIXiZlFno2t9lL8we3SA/8p8+ipFjzO
KWbxOdyYaG/y4X1tvod8r0iAM/0SHPGc6mWgLrWGg7Cxf4RyfT95TrdsAfx6AU6GK+eI02uXGhNx
SDdLP2yzazABXd/2UNpDK4t1bi+CfKph/ADaKl2R2Hg1dgOAne6QzGTHFsD6y5EupCcjBpx0Gsay
TBVuT7ffdOtLpPScB1pH0qtMrqNGT18xXqgOqZdY1ANJ4IDwR+x7kYa+859/CiUKowy/QUOkdAjA
qkaQG/ctytAoJ9NKrXNVtEjMq7YnTk8G9kSx2+z9x+HwypYYoIxRtplufv6y/VYGY1nKhoHp1HuU
xbP94Ki23h7xDc+TZFOKw3NdaOWwBbZrOoK2Dxm3h8qDdSNWimLMIq7CRRHar7SAgTZ4rsPocaml
wRaAcRzP23x2Q1PftLgAsPEKzrBILH2CxT9eFNp8QltP7y/F0l7HjGH5+jigfJGxCZRZs5yE0tCZ
pApU2WGuNdEEpWKZWZa1R4Z9mrrSZkfo8JBqsPpihWA11uc8a8ThVwDN3r+sp21ucgZv9NGiVraS
lhYpc465VXz3tAtuVJzLo9HmLR8j/koSNBg7f65FqyvUYb5MK+JLMyr6nfsnFHBRw/hwCDtDNYiv
hw+dI8jJDvQvjCQkwDdGHs6qu0rd5H3rSE3M0u/snjv6/wlgUvJN+1++jZHg0FKGM8WVqtRlwUX2
NTISu74vyYJERRjgNRrFfKxccmvgXZ0P8RBIPHGLEzwSNgMgnvAo++hdfqkMwZ3wpdo2F+20DDrq
XGmabARVu8lyvCwdZD2AofJN0cuS2lgVe3Ilo5NSKR6fa6iE+xB14IsY/fVSjqYHbMKmzS82SIps
7fhSBpwwU85Www97Nb8BIRrsjaobizLCzUq/PTuohRYRuEd3Z5uCwFG0LNMXgYsl52V1DNue348a
CxYhM5kMM51AVInTxiY2IYut2T5ixBcIR0JpONM30MMnZl20jGQOcgrtMpNCM5jleHHS0Y0qEC3Q
mwVC9fJF+qsDBuEP5DfII697Fcg35W2IeG1gpj+38W27L4ZcOcIlJeqAezPpDRfPDtJmRM6x7zu0
7OwiORiuvKirX9/Uh0h1CUCngse7GJcpIj+Lh3guagqQHLTq84CYnUIPqVGkwPh6sRj/8y2szWco
yENJ8Nooedeg0t5B8u8voZovItq8EQJfwtvUnDL43rXoS1nQS191DFbLCb8c+m3pl4kSa1ws52Y3
VvI084CqrjmeKYRjMkkbjxIbYdaD7Edhr/tmyLpnJKPmmb2YBVfoiZsW1HxHGuS5PvR0Ec+bvlpb
cvjjbPEvHFGj+GZTtHhqjudHZD/LuPpzvx54cvjJJH45D2BuyiFVWCSAWeQCvEoTlyg/ARvPl427
Q0aVOMzDZ903ku/OkGdLYJVjpBBGVrxAcS5cbH6ybplLUVnqH2Hdqat4EgG+y7L09WdyJjI9c9rS
k4J++UVSgzVQBY32mGHE9Eu3xXNPwzUVwQynhTxnxOZHj9GubIm3n8ch179DKe3iVUMeb4iDGEzN
rbapoW+/TDCfZHgpsDeXOFNY8GIwbAlwKm+Pq8S5V56ylR0zJ0F6UOT1JslSvpX0xnrImrHP69on
4OABkHA9ry/ykVdbdoyDqI/EUx84bhc5M4/ozZ3HCwOcZTZrIEVCmZ0rocZsRcyBEH2jAW8WRSxr
xFNfLNLxJ0RINzuYewtoEZoD+gfgKWNPoAOtWzTuQX+LOraiaybf6l0deM+TjuTnEhMStf2IEf0v
KIYXXkA3kaW2wXJiiC6Q1zowPSuw73hk9Jzv0t8pTqCpYC6h7qFYvsnD+1XhlrGy15H23esrjjyn
gZPOnyc1ydvyI3vIwINEbSYV5a3pbARXvNJeCi5V90DSjax4yccZR1eY9NZczcp/Rq/huCcHLD8n
MwFX78SOJfNxPK0Z375UcJ92VNgbP8fEUl1kL3gAqjIPilF2nKQOnsEpfB5K9drSN59UGGHr2b+1
uBgOtJwUpndLYV3aPM+LvbX/QN8RFhfphHTG/U8um4SrzMRk9DvLouLQgOcSr7NMLNDGo0hWzkmt
UXVx8F/u3m268IMkA9+Ln3iSRFaetBlveY8e5BQeGAqbzNOcveInAYvnbj0klxru9sqzn1b1/Pur
eyhXMQPZw+qFTpxBROMVj0SwzECOmymFTbvURmZTHWS8t0khtZfcEp5ZVIDf/O7ykRVOt4AlrIgB
wxkl/DfUq0lorwTbtHNnvQ9LpPJmiwm5K1z0e/WBSleLiB8CpiYbrYLbXUvWoWe80O60XHPn749v
PDjAqjl7L/4i6ILEbh7UJzpJ7rMsAVfiIKHZ5BWlLEKEvEQhhhlpSm+5xnyDWB8mDmwpW0hutVUC
G6t1aIzIfJ2TMO2Ga0YDorwM2OGsNBofTLPUH+U7WoMibDJ0zySAVGA+AO4ugceIHBlDLq7hac9g
JNjWyQPRbZXdM+Fc+y6PfwztztcgFdY5Q27XgKHINrFdxtp0/WYUMFMv0BRJmuoldTPLHJUPpJVi
IVyydO8Bqn2HlRn8x4maalY4XjO+sY7yJLqCWuvQ6e7ZLEL0S29+uu/8Oix68LtarBxiWgPYqSBR
/M0zne18+a2x+PS2hAnJhSx2mfFI1QJupqBRa5cdnBiaA4UH6O3FBculPnAD4R1j0XNo9folVg7h
tgHFSQ6FbRfBmVlakiKZKG+YmC7SenhJrN7mChdBYD2Smhyh38SMHokl+D+i1uzAVkZ5PiZwt5/E
RW3dnZ5ozAQDuiZd+1JoG+XsDOeqFtH75cBPgovx8a3VRUEXXeeQf/B2ZqBSX7A5QFDHPGB5ljwn
PEvLPt/Sc2LWGAkx4VfQ3n2ZU//fb3OPMiGMfnTmyUbRUvKPkHZB3I9i7hUIL1R9ICu+p5SqKXAU
51zjuCBIEC5k6UOAXmO3+ebtofBEQ6Y9gGl3CT7/nYq5nE++1y82NuiW5brL/+trbMdESC+id8bZ
aoZT7Zs14s0iNQ+rh3zjf6ZPoqKpdsbcm3lwv4HN9Bg+N7kJpU3Pe7h6L5y5CdYK7RIV2pD0XkGe
SSTk6NNqAPDpnpV8/o1x32TAw+U/IORxZBEBmvLSRgyUkT0Jkx3xOp/JzmZ/l5f9EiJaetgqeZkH
ANpJHCMMKMWUczAf6LZKATeQeLCtfI8Ef4qs524fHz2iwcIVTc5CfcPFycdGD6ufEZ2F+J8dAC+3
JSudQr57pU+/iXFwH6bzq5KpaKB6PwjJZpMQ1he8JcuJ+ghHN+LXAMqv+tfRHEdyFa77DMRbx7XE
4ilOVIdnbgR7hCTAvuOevUsBEzNfgoZrEFmz4hVUgFH+rJ32lW55WZV5g/GD7BBW5FM6eNhGq3fY
PoI9GYjm/E+cBvZcSDO5bMFxKB8dwxGqAHUdWJczTCCvNMkgNmSsEw754qJaD3jPxiLD0B/pgajN
7Iil04xKxpY2A1QK9agx7KfYQHp8uZ4SQiB8u3HcvfJrjFIefpCTRsNB0rRrWyHMKDXr2JiswRdl
KbtEVZodyXID++fNRPh3gMdC/01z3YqmT/UUXVWooh3uurmq9TdUlB6oEfvRxB4JOdB2gZ+ChBcz
Wf+f/5pbwKf3on7VjHy6fZV01aV/Nat6y3r8CehRHDwIqYEwaRJjqvT1fZcD3dwFrWTfhg71vOTJ
DgfUp17WZgoY70OKyAtTvaysIqbnpmVaxt9N/6Y2zrJvZVKAmDxJcr5nNnWIfvsoNQpnQEMghVNh
6PNfu5AyEQSreIJ5O7wmNAnzoT7Ya17NpDNXPgMpvWmnvX2la+3XgZlB8qDQkmYz4vayAMtNNem8
W7sxT7stC8T8xDC7zSAh0lTeL34Prh1E+jUMB8KTTbEKj94Z5Ub9Rg6LZsvFe8IMzvK0z/CTXpTX
RO73ufVjmLadioj44AasVhPP7XRJ6nZScrzB03QqF6yCx6f9Dq5vsEgvq/kaokaP/Pf0F/umPI02
A2i8wQeJCVLCT2TF8+wkFMjUpj/oGPuyOofV1Jj5d+IOr+cfBnWrrrj4P2IeBQLp0XFN6lj7lrET
1rIQ1ncuhVkz99oO91E0KMqDJQWGbHYDfZrJfdZkKzx3Llwxrn23LA4l+2J4Kk2O59il9M23RA0A
bNSCf9bqBjqErCAKkQez/704SyCAjEGUamAp22YqwxaZCbB7XNsa3ByjtCPjbDgk2mXsKyT3iR8+
hYkpCZjzMxtiR9w7hgd5FHYBTS1vEVxh3Q7a/cBmC611Z3Sveq6ZiLBHz1XhZH20GNH0g/fZCTGl
KdIXa+M7kV8dVnKf/ICpX2wwoViupzxjgodkUoVKKI5JY5qUeBfcxfSgkSvp+BscRbWNu99Zb1DJ
4OIpWPN/wAg6FMPfcgCPDyaxC8cF4ghT8tuDzYNo+YupJ8eifsfh4zl6dx0pReprcvMyh4qBOoY7
Bi9WSpK09rJV4sVrTONzRNnEqon9NHQkM24WS9thDqT2YzFRfc2F2V++ALOh6UxWCkS0dY801tjd
3IY361NQ8vv9RKAlSSPXvhGm8RDybRy9jeuIpHGtm3189e/wHuRaTWcrEo+egIIHvTY+Ud9Jw9Jh
pN1eRauQTHZhQHNP7qz4jI78eyCmSTT290rhGogpF0nMj/O/Tn0h2Megfn5W6EKsIEH3rbQUbPF0
DS0gM4LO2bERMk9Wiw8j4XodGz1Qc4vjOugGtT/dpHK0McNnPSa7tYmqJdx/CEIiz3l8aYXszaKG
gC09g92VdW6eOuS4TqvCGxKHOUFOO8uHdMfYpI0f41QPHWpHX5yax24eKFkAfAMuv5u1zsKC55HJ
sC/WqDatGhx7HmgTBdzWBZ+DESLJ0z4569HX/NUDH/7V0E2sNhAkr6tkD9kEYtfjuZ7jIMEbdfFw
pDUCZiYGQbGEMsje4Vv+YnKz8hdSBsNuNGj2fLS95xTtNyTgaBLjxSQ3CjRLP7a/MYVewPSpeVQ+
JsYGMreSN5SUEzfUL++krXVWSlwoUGFJfQRAB3O/egxJUVMRx/Qe4DMvL08rmseFTrFTMWIvjXKY
cpsmZO6mCvW/36Kha/sJ0WC8cibdSxirYbdXKeGVKKaOikrI16lbV0vZVcYI9ie8L708dB/kbvez
monc1l2vaRfXAArZ5mipdJDqlme7xzqE0F1R0ZFiQwbqITWlx7wKndE3evSjbabdYMuFT13MGk3i
55da+dU5US56W4EzhkLgnS6B790cZ3R53bv10ShA3L1q7WqPiyK9pN0xaHcMEgAqrKIS+DySp72S
xYIYpx4p7Hl0LPKSQa3RCDoYCInJAZrcnxXQuy1B04NfL3qE+2f68YOHqsljTBjyFArIFWWcGVjP
nKvjW6YJJ0xNMKfRVcxm+TcndZXyFzic1QxMVZxkv0ahTR0kJgmBZnvOgsyN+/4GleyjNLilmB3R
jpCYPx/JzIIAlTwI3H0oSJO15OpYBVhez2RTVnZnQJksuouSqL4d7KhV9ORjJ/+FRbqjJiFym/pA
65fb7Ah1f2tebkzyfXyFit76r72QJzebr1P3wTilLplkFdb4ZTFwjD4TgaFHKloBmkvLHu0YN2Q7
2dc3h1Fw5KTEWTUJtGeFRIO5sFb+ii7r3MROzauelKRPepDX4B/AYD3lCCc92sbqk/xOOxVyDWTt
KvjjpaAgFfTGVYq5AuzoxZRvJQ8DGkXasiu+o8JuIuo8rD4jxx7xm24Scuf+GwA7eq0qdMuKqdka
eQ6d9leRvcYLBOXYbGmpG7yQGagisJA/abz4MMSHa6/LvRA06bLrqonDoRlBblCsJfbK4/7o2eQB
OH5t1ZZ9rnPclzX1G6yHW+yO+p6vM1WBsJaDkX3xjmW3pdza9C/AiF/3bYBvHHQBOo7EJPXFozqh
2KCZMGrC3EaSUbtsDuyIoGSDohswxcgiYQbknCGxRGzUgTrjeTLm11zPulU0BnpB7ugV/xH4/V0G
G3r7kJ0MAqfLQ5tEqJ7B9NXcxXjQE/x6m42IimGN4dofnfy4KV6utvHN9xRkG0JOHlOAewdyetfL
EA0eyWacfn7znrGYMkUeN298u3O//50FkW6m3v9l0Z5+52JlNCExbCo4qj7y76E1CIPU88SGAqkE
RUERW1aH6qu4k8gdV5C9d/+o3yMn8CYmjaR8+R17/XUO8NKPbaUhwCmrZHOSsEoV9dN8K+qHeMtI
Kc//ap6JJ9LozeMey1Nz12mpdnR3d2mDJxYamQXRcts61L9fnkYb52jWFyl6ETg+NjVx0peOKKmY
/v2KDbtX02Z4GBV/G0jgkZQ1sejDHeFmLjjKJinWxI3LVPkyOyZVpy1uKbukorLoFlTqZAQ3LR52
6PEIk7ms9T5t1By/ImdS5wxZqq1w/VwBjh0j1i+Cf3vbU7+DWYx0xe1MsQMtVG7HC/VqcscdkApf
6ToaZ3QKsUgb3NFkUlXqtiXYAzJ/ClvrrSRzlHn7F8F+9tdaHfhlYcm3FUd+7K593QcMZ3oUGFS+
I2kafORb8J9xKXwMIxio2cBIxZWQxVfdI6YRuGKpLV+S/Y6fSez9qe1kM/1s1lrHRvqlvSP/qqF6
OrK7CmOWJ0SoCkMaCTHGQzYjozzcrTQlc/gnMLO5dQimHr+m3BwDDSvyQ0zLwC6X4sE5453PDUbR
iyRz/zKTcnmqeYTadLZQv2a71Prh2fU8Cen7iXmlvvEHIW7h8RD+66JHkQDGJY9HI0jtS005h2Hs
OliFNksqtGjTzJN/v3GgjU/q9Dfp6d7SW0WaMN8QlftW3RSBm/j6ymBa3kJEHgP234GsM8FvsmII
KJr1f91wZs8OgE+qt2dCmARxNYG2JSZPLBastp0yRVGubYHDat7fxR3VJvJO/rd+BOUesK/CgZiv
t8thn4oKlNyztD/SM0ahXWpSoLrsaPGpY89wyZ5V+PTIirrZ2hMmprpzyBG64v3eohRs4LNhMtZ4
yeyOb19T70sW0pWftUK2EOf2UDYkzAwxcba47CN7v+B/s4BV18liOWi8J4qQBd9UxANH+Aemnrmd
2uVqviLupPMzFY9D5iNpaLLcBhQT9cJiuFMLZQlT8I1jhdOlMNg68LodpmEFeSEX1wzrlcxbFuVA
O4+t1sp7Tu7FBGDuzefHLr1hYFXp1mn20D2hfZrakM7t3WDxjCGdhnrndyEosLn2mtsw+h8DcI0d
6hLitAhxaE7fFGujDnDalz9ES4Ui+wcE+rWpyRZ0sjvts97U7XdrMTopp82QPGZmIOTLI6opNtrv
mmumM3y+FF5C5lMuUqqFSBUTfYkte81NuSsgqjtpmOuEDGPW4tQ9PnegzZuuApPLBGKlQUdQxFP8
mdzzu1UJPOHbd7L3oh8iAdk0cqBQE7wyO+HdiYLdKWwaDJqKinxXzF+Ik3PdhDH/Unzb1nv3oehk
RunebJmUP6REV4mlbCZcGNQ+bFSPdUDL0gL6JNh+50pcCRb1HoUF6W12L+K4M5j9YAycgjq3v7eZ
OhmGmppLvRS7bMx+n2WrMoAeLPyIkydL2Vo/lkNTqk5S3DPsK1pt/2X9kD1dOm0vjfzjRTaZlKSp
ap1Y8cSHDMmFzOI/+0zWZmX3p0aojhSvGp1W8+QJLMGCkvak3plD0BvxqnqBY5jaOcVvYlFkaRpB
nNcMiJ1YqrFIwbNCnBNzxHbpsl/AjxeGIKMksFSTMGVtOWmPxljIKRdm0a5DKv1OUL3cd1XDrA5I
V0UZbrn3M3Ct01cYu33yotU6bl0b+wjdczuxagA4JQGZ1qRMcZXorcniNqFhOovY0f7Ar7+32nUo
E/8W2wfuY7BYfDLm++ZbAdePBzieSC2xbY3tBvyn8EKB8ZOD9p6kQoyjeYHEd2nMh+ZINgrJbQVc
Hz8J98E/gtjCMCC+A5osdFTrhKj+tdL9q+A1/qFfdzg1J5M9QGV+YnLq0bffkIheWOh2dC+13Qoc
fOtMx8bNujSxiJ2oKcZKIlpd+xKcD64RcVTOt9skcTOcHrV/kUJWh56cxyAqcAauMGFiW125EPmd
4v4Pb+drOVKYTENeU0boS63sA1c1jbB2jjsTvaQ5b3om4c/5N4aXqJd5i8FVFmLeVVnkEQtHyLIi
uz732vFJUmVp4qdvsSK0Nmxty02tRxwM4BDd1rwpS4AEYWPiNsiyxtM8V2BLLX97Vwp33feK4GJ7
MMH8A5ty6yCmXP8Adt71v9WpW/uiWSf+o5xDzaJwgt+phj5SOZTI/TRNM0C/q/qYxymPHTTr3g+O
4+ScoDyTpcN7cAj0smzSe2w1ZzcF6EeabqxHbRUvk7/y+QuYyBcOiEw67DPdnMMaWY/BzahAU4eq
TgnRsBUOB47JGYhQVk9hY99DK3FcxPzJcrLSwMUtaPOq5g3viV/r0fCW9wbSYLcVBdVuIRPNW4Ay
H4rFYpmf+OaXHF5Llnna6QFqUHoR+NPFWcY/HrgIUSUyFe0xNpi2dWo+woeeK9cOm1ZNklNjrSqu
9NELihSautCSTMbp1ShHDQ8c7Qk9NgpieDG8g9XK559v4oYwl6eIDq/Icp1rxSB6Urm4icUeaaz7
+72TNjq9ComN9H/4thh9wsIXd4qO/f1jh3lGSFpA17laXX3sRLHkzSkLqH/44Sdw/H1EJNs9re+f
K1PrsVVgkFMV2KLkj0WnV0bAcmcPURHnzSj2d9TSN6dmAivpL/bdVE8G7VmlBQdCDnkRsRNlwgvg
/XpTHdBeWSd72b4z7duRn5Mo2X69Bzo0hgSHJS0Mj5GEyBQcXO3I8DVyrxBnd/R8l3UHxzE5YsKk
FJc+qNWIDPVu0qm+V2WfOrJShSw5jv9+lGrI1tzsKR6rdNDa/J4cU794wLME7r+m/3wRbp8EYV/C
wHYrBPWuqbChMhMzBvoDFffSYUu+KJM/YZlmUAhjGWtuEnwZ4pyClQ823B7z/JCAHSsTfQX6MBAQ
WgXP7BVEEWMUouyVEN9N6lZoma2TDh0wurvQpJJXpAdFtjKld3/wjJmx3hQnHwQY8bPAhG04HVTE
s8Z5pi1PVMcpA53n7qjDQQZh36AlMXKrqbu1Q/XQ8Mzrat7ldSC/iw7m9pQKlZc3aF4vcaYDFEfw
L5d3MKYYceYux0H4rqj8xbwR9m5alneDmEXjh+oyamQx1uSBWroNJBrEqUlm5utE1/aT65j/UfRR
oB4AYoY7DFZu561FF5B/3uiQTORL0FUyyg/hxAg5Y3bzJiMiij3spXWEHmxUt/tKhAQ13Yo7h/EE
UOQr8IkEHHuVRutO7/mmkZWZhXEepicDzcUWw2Cn2uSm9mTq7HzZsrtYvFBbN/1Z9PUSY7X6+jCX
aYnosf/CZaah5213u7xxelA2McY0x9GELjm2lScMImmwrSswj5fOHzSSJJKmobHqYegqWeMPyl6b
FI/O6F/ED5dpWQcgX5LWvQfZ+hIwz/cDpgo3xah/p7Dw1LY8q9MikhoyYazTxU4wM11tEHYfhwXf
qTNMEAyQGNeFGodWQ0e4IjFvKdejluTadv2zaoOj5DUYaXCrhds3uC22Ffr2T1LdOj6QeY3PRJWo
sxqzqOm7i5YA6x2O2MgH40NF7+q61Z5EfNkHwhqVXA2l0Y65LnkTZNXxnEKhuizBUjl4KgZ29aa6
sqPbn1aZO18pyo2JxBD8eA+MKiozuRBoOGYo4Q1I4ddxBkTXaQonoUFqr90yyOVnGUKGhuRb6yqm
/Cnpwxoptvzf8LZNTD6OwMyZtl5gT1U4drhEW8KFudmZM9QZVDpNYbOd2uqfl1E12Mu4lz6wiYVM
y+X6rJo8X1XUVoqR8MeM4BH9UgesS28y5WW2Hsst+EeeReZdG3hqL5q/47DB91GFonGKd7RtgW3e
fW0XNJM8s2ZbshQKvbQMRqGCPjNvT5qgUn66Elr2tSQIpejpFhqoevrdSma1cEpYFIrvqZFm1V5z
DMXLWbOSy5sF8M+G8z78IY6bw26h6uutvcvn2NXlqsVwHrLQImgbxazh+F42e2VmU0o6qivgVBBq
BDqVpXXsGxeRODyvgXvz6xt/x9Rbioqt/vLoRfnSFTyb8AI2jgQYS9OQ8V/sbSgPP122VWoKFjiW
PygwjUec7qOGnehKxyrRJOtB/4bwlofZDh/qbvS0BRVdyuF7QtEHaGhGC91jbZlX0CZW3mi0l/aR
jITY3jAw3xXJy4Kzo2C0k5yO36E4abH4NMJNhxf6CZPNEMKZSLZb18+YMBUX7KRhjytfUaSxPfpH
Te7W7RYV8MHJaXqkpJU0TiSXInPGcdt46wrLfXvb4xchHml+kA8xhMqELBfRNY1/CvyMn1vmnwqp
2UwEuoU8yW6h7AGGiDAhQahodHKZU7/tFZ9a9VqLEiqUfCyxUYFvXvRNgVx8vIS+LJMbuNYhbEa2
vITt4c9yRc8bcu7qa/2xelIvGh1hq6iUVoPukJPcd8mLmLYgrAiPs5wWYLbtA0h5T8XQ9PynRYzA
x7wUoc/0rJwf0A8ChVvcbaAf0fGbHEd7/iM4h5XegtUFRyyMcvMFv1SBlvr+dMNpErXenMn3zmOH
s8bXej+1aZ9H5i1xNykSWAHBTNE2dR2Oo9yxRJUdItqO0LxkbCH1JF9LAzmTWmegV0RGIyjZDXTf
F/RqAFSJ+lllltVDdC9Qevz5S/X6YqQ70v5GE4SzJnnem6HecSvzxHfUSM1T+tnQ50mXi0lYelpW
u5wFA3tRFVOZ7dOeXn/rllUG0HM3MAwBLOlcO+Ea59MmtXpqjyDyLXTWoIRDsVS+mS/YG0cwNB2L
VM8w+jKZQwNynAYeR+yW0KHuJyvf26KeT9ozeAP1N31/l5QsBUxJO/1H2L1Mog+Y8dL9flrN90+/
CmoI06HRjn056pzxGUn8TCGUd6+o+W3hR6TljPJu08Z300h4EwdH4sPGDFsuiPQ3sMEgZPKYnvIb
YvX0L9wW3V+4OL+PWhDGxz2HVb89AcisIWpqUypKRMUr+qH8V6U5QZQlnR4/8E89fLFm7gwn+QOi
vxESS9bM95pIHLsw1Di/i0BfDMAqa6q/I5LG+Wpf+6dZNljasiUZHzac7BsbcXoxlqfJziV3o+4v
PqI4/6g5dqlRlj+E4y+uEHK12B7Vbd3oomr4LDbEmQkbDlTH/hjAKRbxpK6x+SSB7eUVqJVpzvyn
PEX/Ysico7vrTti8tIVOzMVAr8ouCffiz6zrOB9qivuxr0rpXpCDvWJ7tRsnBDuzGYpTuNE8RoCl
kV4OIPF+hCUPAi1IPB4Hhb4U8HY/QEJtW89XMksInIClFzM9y8V5KC8EHZ0J0UyW9pOHDLf8vvpQ
dg9Nods3DqdMyu97Wr/ZgsyMvLUvSxEYBbNoq+pNlrlGHUTQ63nMSLAAg1M+MuIb55efrsKRIbKM
NU7051MqJnLpVxRepS+2S2LD3tEPERzYUbJTPGrWGZ31c+54cnMbT2zkHBHPWTKLEJ9YcUNoaSiM
rRvgJgiiMHRMvOB66KeTvC5l4JQXKG4ozaHn86X/9fNQsb/HYEx4KtAptK+EKE8sR6VnKzr2tPnP
qFb/Y5egsUrB+V7TQ0Skjxt8sH2aZSkQMwAdaoStG2i2Xrn/Y8DupwjDA31tZHUagiRQOKNRAQrs
ciBqAZ51FcFjtp9Q2pYWK4UpAeg9SSE2Y4zwIiowXO9UQUCFwFXcY4B16fAxDxGrDmZZsFg8yEJv
aHP2Rh0yW4M86wswxmt/AbPW3WQBgwG7EhkgBG103RiG4U3aSc6ORxELaDLuRMmAtrLUrH3q0K1Q
JukiLtKhXBbQMltXTIm0OwDU6iYInQbnfuqKKr1Du3qXWErDE99drL/i3EWt9lxJ3yFdMpzKUiHP
Ke7B4Z7J84HBOumvnmqzC3Cr1mJvkdLbTJJydvPrGhUUPRot0pyVoKp7BKUucHpDFUhlBr7yys5U
DMeNMkPG6HUFZGRnGlcjhLuA/LZAmPEyAH1i+2NJ0h9nnn82pIinGMQH29a+S6jSJnjNX68ysjMN
DNoRTCXErE4P+tHwXHL8ns0C2GXPOqOe7z1JCRcvwEH2RlD0691f9hSWl4IcBmFP7sFGlLeqmOnx
QieEKQ3RujcVRjKviatvw3VBUfCnXBQRbyKXy511iax54fup34nHKvyMjPkSlJULmro8WEsf2C8Q
77Of3zcJuJq6sU2TLvg0+0BOpFh3SwfyQ/QMUnapvz5DR18X/xIWPVZkpdh2wScrwjbAYBLeEImb
26TuyAC2nTttQ4UtAuRJD/kbiCFHM6EMnQepk/G6ya4mQ+ELvogkqYTUP+aXouP3t/XNo8+s63MY
f8zGZtFsupWZwIARtRTj6LCDDh8rJIfTGOVy28u+69FBeoHNGXDGX/UVzCNff3sT1VfGTmh1Gh8U
NQ27vE4Hj+KQH4qFbXwr7j6GQ+3WZ09ahfP3uVylhC9EkvmklJGYBPIZQ+JVFl5KDq4u8cuSAjl6
0Pc2dkQDqGmtFUtTWIaijLDYUViLq+iHX4DsMVKYFblCPZbZ8e9wkcR4JrmsDRSOVcHXEvbfrzhU
ItUQSaAQEACgi/p/8HiffOro3ZgpzchI46MHjj/5XqjQLsdZkxQ8pM7ca3NLbqiLwDsVyHcNPG03
YX3feuiGKtg7cuu4ENLefIPz4MALUcKdBhSuPXPjOIO53Bm2A8Finfi1tamhf4nZkJkAvrrcMOkO
MUQpDx3ZC+6OK4N43vw2oCdZuQQmuL0H/hnVlVij0EOQmf/vjU0E3YDnR9aPOvlvpbUZPBGSt+Hs
/TY9rkcmiuwaJ9/GWtb3uCNBNVK8LCnFUoLfCGupJt/we+eE2+0q6bQTFF/0PGHbEuVQeUX1BenT
c339Iwa9yqaxxn65XMcWBGmLOaFWZiv5SP0JTbswnASYpT/NPZsOQ7i/ywagB/LU32oGXSBXMe/N
B0bV0JJXgPJU2/pzYH9duzY2Oqw/jxBlwIxTBdDpx/V7+DfQwLFNYE3i1pN64vJj1qo/27P9Inm5
UDvQJfh15zLZXjFY39OBI+fjScvj3prqVythm4S3uCsniqCtFQIDhMwbvfFtfM/c1IOP5tIjF1g9
eykzR3rVyjJEmnWpV5HmE/wfJNefcJxBWcnyTBIEo42f3MBmFI9qoecAo6Dyd8tMuW/5nh31O4Qx
5F+WE6Y9nK47qlp/FoMNLkRzrO3LI44xyWVKempEoqLwwRibRGqyN4feuCTocy7Wpv+P964gG6/f
tqdDaTcBgceUL+hjzabnNHoann3cW2COr602Ejb1qMeNCeu6Gkg5qwdSz1UY5KyJpGLY4dvRsSQO
TThJhvnwR6+31u8Z4I96kvdGccOr19UJHjpcCkDX7RuUgAek46Rikv2TrdojxqCguwTCp9Lr6MZj
L4bTyMw2tq8RbcgoC+bG2X2EmS1nlBZasHJZhjRTiURhzGJmeV+xi4VqKQovO/Bf4ROo1plFSNnA
xICjok7K5xghtg7uRQytPHZtUC7WrSCyBOmX5HHle6cyqOFXa+i70mBTKaIZ/n6pCXDz/zyYbhHx
njBw4xQz5elVPKm9EvJWQBCDuOZMbwaUP+BAeDHaZRFR3CFR1zlZo+BmLvpwJJVj407rUAp2ohp9
9E7EcVN84F39wJYEcRWcpz40bWywyUpyTrZIPSP8CnwScCnDTUlooXytky1wgJI0uK2Yy1uF506e
SUrFXHHPvwd59Tz/ERxy2LxFJV7ODs0pKLXx2m3BnWC+rvFwsZpIEmqehZtmXTD5S/rlbCg7kp0G
JNHCKd2yXtmVO38zagVDXxx2BiWWFrmFBoJeneiCb5L3P7Q6WOMhU4ZaYcNzzYKUfw5XrMPWe+l7
Ie9xJ2lqrBUO7Fe3teDWbCwF1k7V3J/a2/vBq1KZ7m4s49jMS2a02e6QwUk80+8fZ1ezlZp4aXHY
vhyPPgUxuirUfGyijvMPATtC0MOcWzrCo+hvVp7mhpEKaN5TecK5ewYWZe5XQMsO8KBswJd7Hmx7
6trDhjtdm/l6e7TxIiVJ+2MSw8no2nLDVmolmyvS7s2EBUS3NHKmkTyTR+3+YXVxDPmO5+VZPRGP
DGZnRpXQrqhDilFLDY5HRr2LcvoCkXROdpWMp/lnjFz5iP2HiXqB5Te/lJv9YlRqB1gcYMBTySsk
y1NPHDc1PzuMJ496U+IDAwGjTIzUBoI0IJkMkxXyxINlxm4jIv+tcdSujA1Ztg/IewUhb2b1j/im
K/yfOsbDMzMzXkt22vYeQJjvE6HkyCxd4OoHiJBVTnEZgh8Hq3D6WgHhmrjVbWg+KnTPDxay26uP
2XSfUbpD01P2HNksw3M99jcFbPGK+jWBdSTl4LTT62RO/y2wI4Lo1T+XrCXexDmunJ4jY0Ouhfv0
EC53Dor0QI4u8c3iFl8CxgNwna0LaxDa0yJQu6Z4kOMC4OPZC6Hvl5x9ESxzBsbjLgj4CV15XnMl
IXAXV8WxB2DySuYOPgVBdVJmfVfwuFmVJewfPedy4q1FICS7qTV98QSzoQgDOW6sQuy3XPf8yTcC
ufTcHuBmeWVnC6cC6PmK2LcJwyAGlX4m+tX3LANXGe/llQh06uKmyB8f3ugMqoXuguByw9rJtY0r
SFDVttJxWQ8DSn4twFbRhczTejNponK24XSj/Q1fVsbGNjTiWFvB0OOt2UUTohGe854jpTnVXF1w
OillPPB6/f90zWvzNJMEQPUSj3SMARNXIOvHxeBaN/boREluT/EgZkY92/Q2Z8C/JdusmAKWYXn6
WuoNcdLLb+4PZB3xlDKB0knDD+m6rME/HoG/Zm56HdywtgWuWQZieGHEs/pEFL4wMS7u+pF4vFu9
ZQDU4pPlWbTr2z0Wp5Zt32utHgmIMzxAfWLWljS5F9QFI7rvwQLrAtyHN8EDrpzPBE2ENLCUMnmz
GIDtckVnE1k/bzKKs5mqMZl3g15p8ta4/hRulyw061egk7YjhP368anWxbQHPbDcSKhoF/RYXy9z
IzMSsfyTppR3OB3VgPpioyvQC4npfmYgcbBNXYJdDjsTGLHA1XEVD1JcmUsFdjrGzDJhXllBbOJX
a7679f+SB7U0gZLfaa2b/K8HFzdz2zXCBCT4h0vYwhCWcIbs9pvHo896nAdFBQ3xETxeU9aeCPaS
IdS/F9SjL/+hHtAuYO/HSNtbWpkcgGIsKyxpx4HAnsicY/RSKWgwE7QmHWWvUwLwlRWlTI3KLv/F
RA3QdWlsQ1OMRYPO8Hb7XpMeM3EoMPoqciGn5XnUhKwjPrOKgSLmI8IhEt4Umb0bd70/2+FTMWni
yT7Dom0zY58o4+AGLWoLb48Sl3QtlFEigmIWj4FnnAYO9NiGvVhLYXP2szCqF68nmhcGUGi3FeEj
ajKs8rKXWoMmhXrcTzfPjGPbvfC1IMwKgwec4Rp9ejFNLF2OOye9oLKk5/iVBbsMk8vKxHzg/PDU
ABUgPpcqPSv8M7HjZ540hmvEdcfSyGi0GVVWcrlUU8lm3mzWLnZ2hDs5FuWnIfDHqgYd9zNWmOJS
YXDDZx8qf1/L9ync+5ng6CHdFMBD+XkcaNihIqVx1eHkU3gnVBDuodtDCqQhcTr1PxDgM48IN3ca
9h2xhncFebSHh96X6nl7bm9iwshdDKVpXst2qbbmSjub53fZc2wJC7XVS+MuB5DMn8RMB9V0nDAO
Mkr+VdfnAWqVlVZU5Spv3VVExcNtHnVADuLYi0dDzBL3dfS2/GK/jTYs+cUQDOFDRvJMpjr9TZWi
7uv8d/n9nLc7vyuj/AnA/6VuZc/k4DdU3LbQneOKBrZxSR6gA72Rt1MyCGt6XkxfwGV92aQQCOzQ
HJ1wYi9WjiyB+qktJ1jVQjUyBEpgLn7keexrqsvEb9vY8G8YJbxXeJ0U9rc/k846brIYOij7J5o0
t/P9STy+ieTUQSwMEYVUEOJ29CNqI8vrhpdVbalaPpVoXQIIjk6Cvv/K+WFNwqszdKQHMNOWzAoY
WboM9E9nogHSpyYn4wSOD0t9vEebMDhvlpwo8R8PI3GmG568nLnABeW9Qyblnz+HZbBp2hUXmfev
JvmTAv4b0+7ZEN3wn0nAlX5kRIwKna2c57cZzefpiUMV6BMjZEEV5LfqIXYrkdewrEjgaYlOUvO1
B4eweDsyyONOU8KtYt4wBBdxl8csBshbtrx2NzfMh7hbRjs451dD8xaTuJ8Vdi9aTSu2l724wrjz
48rRDLWCUL990nH6MixDLHvQw/bfGrFk2XDr9p3Ow/3S9BWtT3vCbRu5I1e3/24/GyNCR7/inJ9d
knz9RcOq4Df9HXBYMxi+dcPyvA84JxY01coKUZ3FclxDfPoIcRGJU99iirgAD2kOoEs4sRnga4b4
OjG++sJFuJtXc6tdnmjP2n1cOd8xgACDCo8rx3enqb1ZHyI7KetP362Mz+qLNM9AQ2FohtVUu5Sj
QiA76x915w6Ogxixd8QeqVUYf17fZrx0osyXA/8okCrb4colaO7H6/GJgwSzl7s/enVu7nanxL8t
nHlVPsg6sgE2jBmE2FxUXtKQ/8uwvcqUJ4oEvjjxa6sEsdcgYdv8k1l2qJ4yiyG24AozkMYFIxWu
OJQeIcddShn5DOifSm0fV57Msi1OAirI0W69jVQNzwJtNOlwoRTvChPiJB3RcViOIyGY1gnhlf1G
P/7aM9Bsuh8T7mKZw/uedf/PNiJN6M960OP7DuuVtX40kmv2X4wGDZzU20oR0nSR7woAjFxHf5o8
OU0FVFnvPO/Z5DRrkSwNwHSG1O5xTHiGVNf67VlCQTdS8PYB7vchByYRcIVpOg5+SGsNWhttANs5
SZmZdjC0x4YIQvFhtoKvNEPFSGngqoKg8p8zldTo/JiIUsU6ZsWlcV6VQaXXyQGVyDtaMnGZ2kWF
IxoEeKzn3CYHC/X5DeSlBSYUZD06z54L72F66QX1D942atTg+Yti+PwzFZPsxLnTgJjmd8ZKeISq
xaGN6QImGNTqEQBiNUZeFSEOm8yPt6Qx5WxumQlqkFmPT+uYinPV8ZM2HWF6mFToKervlwjV4C4d
8/0yJM0TUuE/XTSU4M+GyY21nmtXc5u8Voh6qEbCpPxeu5DTMsM7cRMty5RpEi/hm9wWeLwwtH6k
JHbF2prouVDSAkwQIMZ4ZDf0Y/2y3he5zFaTlCRuw20VLXYN6RQvuIUsN6IAW7Dxy3OVEZmNLOny
jeLjF4JerQDNw+p+sAesyHe5F9pCHv3iybKPdArxbRd1arYH7c0i5d10D0kWYouUr0LNU+t2CQIB
WENwbrjXyoEqHSrXtSVy93/qZl+OSrs0yqoihEsYAThpZeYBsW62qRPASFa8JRhkju6VkN5/wMVx
Ka8n1nHEm7puCY+h7OIOsYqup+PmTP2dIe4LpsuOea1N3RimmKpgTbNlKb/uJCJtblLtQ4gbWnj9
eWDIzSlAsR8IOqx7VKVlQFCcB4FTFcN6xhJMkD73/B5Fjo23t5LfhapCUP3DgkeAbU+1Nvs7o64R
0Mt5j0VFYkZJnWNNZ8g5lM7vebc+pfRGUZwqM5FQyGMakGtz15nvn88mkZwLesZ3Bc8FLyXpJL3I
z4S+Yv4iZV0F5wWPZmYFWONA4Ixxn+jgQmRUXt7hfEmeY72maxEb/ibJI7IZmIQJFZN9NZlT4ng6
YDTbHJZHrfeXElhcus+lEZtIrVLkBYFLql5XGwROtFPSIAxtjR5kbLq5jZwEtQ4E5K3z1//KA4T+
WgpLozlsZrmBxBuKAsSz1mYs5MEuPIHkKs/BnObGKC3bb+weDqaSov2KnQADbV/SefgRlDLATzTV
LBDJ6avv1Tvn+Ilo+qSulP3SrbcYYWiL1N/ZOPxOhNMa1nDLnBYmdRi8LdRScAJIOrl0cGE3uk1y
CW6HWRckKkgWTW+7JX0IPQSHBQlt/opxvVqcd9h2hrErCL7xW7Vlfdc7/ZGvOkr/jfOy5ZRiAej2
YWa5HcSgAvvqFE+JBoLZO+3fEps4xnTIN1RA0YpQXiDXiMr6tjYgWcE4Z1PCa2Tb8mlV28uzC5SC
K/KZKlFWO1EtB5PQLqQmOSotMeDm5gHe0FbHmow/s2nUbdbDylIqavwBnuxe55cyQnCpHz2EyWeL
1nD9346JuZSavbIETUExlUa7E/Rv7tnjc6wWGfdQzlPWxTYqqWaBRdBP9/LJ8r0LV+BFChchNenN
jTE7MM1EY/Jtu3iE3InL3B/2IUrUSscEcvTDb+4qb5l6WMHfN62aeaxGIwoiUXVcxKShd/qmGI3Q
Ipgxb8nssP73h+gniisc7PZhUi/QmSUgnmk7quLuF50ER9TFwBV2kOACpzLnWnBnKAUQMnZ9oB5g
Gvn02sM4qUzcqg1REsSDAHUXaSHuCqOD3OI71fxz1BDBiekSPQbBQb5P61btdLbXu+E0HBcl+pJ9
tMxArMwhNGVOlyyls/2acv4Mzs4Xu30eGp83iEYIYqxpOk7IlmG0az4l+tgEIkp/Loe+/Zl5+oep
0lO04F/1x8rl03bfp9sg5RsxWUi5xifRON26zI17yS63c4kXIzYPI0X8hjz1nQHw5pAJQPxpxXiQ
HBy65wE2IQoGIubdWcivDKA1qP/vpO4FH2TbilIomMKk0ktmgupYkKSdJNDn0pSh1fhbxGCX8kuz
hU0mP0sYlwo97X7LG9kyYwa9zokGoQjitcrfx9pC58Gxil7WSLjvcrB+F2hcH4wnpuZL+460YsNs
mMgWo8ibrz9ICiqTC1VxCT2uWcfq3GInk1E7xOTGVTKnevGT6D1XBXTzRz5JUrhCMkhvHwlWjuN5
ULiaMdIzk9DKPTasBdn530hL8LsC+CYtJxY2+ZFN4kOLyvwKCAhIQppvnO1Oif0TPWICFyf18oYW
8ZCl8VCUXaJGOngkmIQEjvrn5uTmCWG2PGLzHuGXT9Le3G1VFqs9Dur2n//viDPmLSUGQshxTjky
/HTgt+wA03InsQ3s512TtdDB97reRNg1aPhBchyvyONbY2SxxXM8j51GIIn9+Q1p6Xf/C3kBAbIU
MD04iOaHTT3QCQsE/706ctVmL1xmVl2ZYejBHFy6WvPzExa6F+VBrlidmiO779iuymLE6PjA2oyW
XBl5CNJbARExMnX6HSzSvM9em1gaVU0/jogm+M+kyte/77jGN0qhklFnKnP3QMsYYak5onT/HuR+
NA0kpxcyGtWBMcwk7JOTM1o9e3Hzuo/Bf1HYqQp9yNQUW63WvaK7CPkuEPYWKVWHk5V207TjgmdU
l1yDFQuQj1FrjGFZ56nMhnwFstfGGOUYDuBj1UUJtjocbdM8b+tGCRuf1eDiXXWUiZI/XMobGWia
ZpHC03DwFrEMRAOF8vcYrWZWXt0FxVcfbQojmaBRVF7CoxG8tVCvsg03028LWsSLjmXoUxtYwTHG
Qr0zub6DhAs0U0N65oFuSTQEzQO3Pthmu0nATt0KROHVEp+CFEaGDccpnEy/jI9/0Qb+595CwveQ
PttOrp4isT1sozpRXrPgNlVfgsFWZWWYp+dgv5hj9gWWe1BzvOsc3ZxriqXldJ/REnkrTEoEBXzG
R721zxPCFejG8PitPNQcLq9MKmg02rryCI4kjrhjBG9kDkmHYNdyeshPXRy3NH9993cP5dPHf6uy
PLY1a8yh/IkMssGBdWnoYLf0+ai1XVzyDP54SoyXA2LUobhuabxC2TyW2OBydqYYEYQxxSzzNtDo
OeWjuNKVJYj5zOvKmx9IJCAndrvztd1t0WAwbFWomL+5imV04CggsynIvM+4mg8cus/IW6rvGXgq
HYqnCN5XsaJ3jLXPQyP9uWOt6pTduJVdL/+LX87Pu+9PUXS1iRgPvxgBmDX5APsEDts+YPbGPZWR
XuhZpbncTh7RPvvIDj8zoJk2Vo+2iKuf4mwUuNz600Ue2wDQbJRBVXh6/sWcUe/iZXZOgSXiZ7fY
lFOFczPNv3zz1p71mkjlaYhHmOHzAe2NmIqbhNhxsBzu4D+gHKq5z/5CNHihAEPiRgF7VfmXEWJG
JhbWpIwCC26rQQC1J8iDmYt9z24J42uVRaK2LFVY6hUpPbadaDTyJJYcDQWq7mapuDwC/3BLYCuG
pIFZurPQcBO94qQUu68Kmj0C4fJCJ7OuG/CQycHna2tlkHysJDJTU9gEzD2ESfMWYHRkg7sV68Ep
i3U1kLyaRI2vmTfNDv20FRuTJByBlvGZEM6S7Tlq6A/RLmRrY6XG6Ul/Q6nxRxTKTzp+T6Eirmbg
NKO3KWCbImZGbHC28zEGHgU+LsqRDYGnqW4q0ij8Bk/gQzUC2ptdTJSr8ES+znXiMjqWEKmvKair
Uk/hsWVNuGzfnc9K5hOnoUfeG9ExnVT2Qyx+y0LQ7yPas76A657HrO2bfPNhjX5MmafdUlz9y+JY
9AFXybHmyEju1EF449yRsvyY9lFXG+3GERiwSS/gSVgm0qztq9x4nKZwiKCmE8OPCk5PPpz1xLIh
nvKRLypb9NweQtvVwSfW4LK5pGjoLggs/nQdIaWw+JRFkz9nLhFrqFrkgwCZf2is3VV3bwIFZdjv
Gy8Htc/DtbhH9LMbe9AytLz1iOKjAMGING3SCq99jTldaO19fVrDczY8fhB77S4ydH9CJOfdzgsf
dMgVqtUz9WmQdwZZ/Hso6QNQa5JXVAEUl/I2rXD4dy/GtpanX0mSPx9aZn62gRIVfX5mngu3m0+E
s0LaQ+LWZnTcI+HdedmL/oZ+w3s59Il6oq8CHWad/h/GzzL5CDimXJpkXwbEM/QO/c/hZin92TM0
wk38V6zXguLyhdHwEGo+KtCsG6AzmKdmbAp/U3Q/USDoGXDDSq8lFnImVw3hKsZLidTR7Nl97n4E
Q9XYjglARWWpAjjqqhttfnk5399IQ7FVVP7cb/z5aAHLfZiEcGvLzkjnpByJ/RgMqK3/cIaOBbwR
JFIJNXXsNoiqIWj1if11Gl/wxMuBenl2PrtnEARYt3EENZ1+scTVTUOyujR/jfkdUO/oHycm0yXJ
reQL+T3h3V67/CkQRPXXPvgjmpQNaYhi2oX5jOcZgQ1n05TPwoJs+R+JOHIQWbNHk9Zbie23kSEw
Lijw7/17SuSp4m3VZ9t1MbY8mbApC1c3YuEupb8HMiZ5AnFSvIR8j9Wms71CqD56MG90k4UROFKM
mdrfooWoSNg6ievgEZAiR0SiidNrPmr3+OFOMC9Zg0czmD6ck8g0ZmqfHF3wHueTNl7jlV4/ntIu
+1WtrzisJRMKZBMGNy4D7UoJ7+dMv9UazzOp0QV1mLcC77fXnwzN3sIiAb//9lXu0es+227hwPRp
yvUW5FnDv39N6t3Fdfc/sn9rCcp9SoU3LmhUN8kkdnFduEP8UrX/qZ4biEqLiZw+QNU7bHTUJk19
5//sQS9W+4SGpIKDKbhQrrAzep/YlsocBPcztp5vYYG+iwI68naCVXdTRAGSIJqIwC5PjPhqSYgb
VMSTmWty6N+gSZRSmgVjD+A1tOV3j8wfH6fbe0hwRdlxskAEPqCXjG9rve50QimvfRFiuOCoNZtj
q2tI+TjBwYhd3hrEp5oPb4m+UtYdE++f+uykyA5bfvkuIkHCy5uhIe2OVSYFwFZb8TV1gjsMTiqh
aj8YuekdOgNjEm3wmg3+lIOJ5UYaW8Rp49arDMK/DKPPtGaDdFSj7cnGj8Oe5n1Kfsvt4t5mFSlO
kd210NM7aB/d+NuL70Y2OqoBbdPx8WS8K+PXqASOzS/faUn6SrYdskUACucluMZ+YVpx+V1IVI5x
CbBSTBQgJZ8OqEs+nWRsf6tU0OS+n/3Czr0PtH4epagRDBEnjhSK7BdCK9uup1DAo/7GXTfbq9AN
XpEWmGd1HKjWE0ZEH8S6IzrCQawCS8bVp95vbyKXoRgOs8oeLcRJF3jr8xacqQkt1rdfAwSxrHs2
mGUsACjtyBwRJMq0/gj/PP1uCPcQy78RleM+MNqV2Lo5xK7oiZCeglLQCWyCR6RnZ6Q4IqtbPzST
NUZNfdB1qdOCsOkSQAEX2ikRgf8fTXUhzXHurtCOk348HIpKHsY71ABQs57YKtx1qZfQU9+RnC8p
aHfswzPtOCDQ/ATeqGzApBtT7JXruYulpS+EPoh5mJUhBa1zIwgGaQ7x25Czfyes7D4um/W5TbOb
dcEQu3NQK2secx4EjA87LdYJSUFkZxrKH+0nMagjwVHyjSEBUKQvcJi77jtJitLxjUUpG0Q7TzBP
+alxaeG+BKe83EKMo/OHC9z0wtYe3s5lARYM5sEu+wtmZ43F9QgVrjttZ9dE9sSflweuSrKUca7z
n3pNBSE7qpvqkZEqWcmmWTbh/qUtEcDtRcSXFFktSENQQvNsGYNyT8+ilW4hjLPuaNDnWEiLNXPv
U9+qGY7Ego3/fe0r/yqzTZOrgBz9hXs07Vb3y8pXu5oqIbIqh/qwdRa6s5fQzwx9B/Tit8hNguR6
Zxd3XaWJngmUa6dH2CjSfIjOEDlX/YMARJdELCwuySLD7HbVlTlchb3g5xsmAia1vFkSLesBvvLU
5ETqWY9p/2c3XI/VF2SCinITLOVutFPl1keY10pyrdcNHbzn+zKhygKkdCtXkKGCbfad4cZ7XFrx
sp3NTmCjjPP34y7XuS/4gSEdMoMb+dVYzzBkkmYr0tApjpUcirjCVyHwGx7HiK2KipmcqOGiZUr5
6tfeD4k6T/VGuWSC5XjmLC4b73/gnc1JRBUhgwmpFrcaeGt3DMdOR5940JE1sbZTb6A8OUBeK4xg
sUf05IwsAnhwRyTIQOIb7NUZFWi3BktEuvIFTaWkbIvMl3hNh4i8ZTaFfABzlGyXYmi+INAaeTR5
aSiFREGH4+DjjI5SYdxq9OIEnT3CrpGN2d8DpMTRx29ADhTiMccCVF9cCNM4LEGJEHomxSDoqd1F
zGLQp+jLrx69OVGDUWc/HXkJ2dC5nu18gs/cSILsu5yJAz7+H6tOAA0UQ5gvhG69yVKfRGbMRdWg
EPXJ/Fjel2dsW66p6bgrN71OKn+M+45qdnEpwkPfxQvReeF8sfEGqOVwUhx0N5iXZywzYWE1qE1E
CjGdmg2Z/+ug9bh3IfslIQC/+RsQWnfcjDTW7rnlFQgd/+dph2hbQ3kAqY1CVJlx1Nyf3SjoYgbC
nNhjuuHU5a8/4cGtaGJ+D4/c4k71lBArQEdRxa35XeqAO9zeHlAJUOC4erxwo37ZpZ0cZ+NKbPV7
iKog1nwnsgAOD2CrmCl0dE+88/TwqvOK4jeNte0QwOETdAWcz8hXhQyQ/rAE3h/Kpkv/AizE1T3i
YfHFG89YoQFume7QnU12VOyuhFCSvC3fECbWTmxZaz6x/pQQ6AZB/ix8OenGTEyq935FIuK7WQs5
SHA9SOVfOWbgPHEb5vvZg2G2MSsBykR2nyRkJBATERKVHFq0N9zoPRb8CKM4F4H56WGMpKqUWtes
Ea7VMKGNem+qc5Vpj8fFsyaL5PdwMLGovp6uIJrfsjD4YrelhK0YkDqcoJthlBqgKrBSwY7RK7Sy
/yX6RPa4W+qA8aeHoP7v9wHYQHj7NTwoht2VCM4wI5+OXvcCn8USXZ6q08vCBH1k404wBILlovFX
/BHtmFFyoFrxXZxfcTE1a1wlfxIIdI1N6lYYndtbOrVbF4jWksAy8k1xpG/Z4I32AjPocKrNLvuF
K9CB+npGTrXeSnysQmZZYPnm/TWdQWHmPI+tdIa3Vm7CJNAXLn+Wy+jnZQvrhcUFqXH/dIxAsukq
0x/eHQuJnrJ6p2uP9XEXEKFM0nlCEPKfUzWbOQQnXfkKj9SwB8kJlgokMasUlmUWEXDiUiNZPtZb
xMfbVC3ile9fDaHZLA5xjZj/ypNUF/OfdCy+gMJQlyb9BKeSsydMNZm06cqplhgqIyxZC16Nsg6a
oIH+aXUd9cTEc3hSHomErEccYGkmaQuTk8FIo+/OvRYPEvrZLDuKLw+7irR/JdKTdf/VlPjyLb42
3yiZ/f0rgo9W5ugIbDbkhZ0tljI3+MZu1SyFx1OrH1v3g0IxrKeYV+HFN8TSb4mnucMVmgIq6kgq
Qn1g7foViPjM913HXANqgcxweMwqPXUpj7s0lrnU1qmynUq04m+P9sW8P1uU6c3A2Sd24tf2bjNM
JzK7ysDYHfTg3BV9+OT1rs7ePSBS6aGS60Tujen9muoxNA0jq0mpMF+uCzCHu7lR8+hJJr8Hdllg
2S3XoZMEl3xzg20cr79oIQCMPHyqVJLzectTAPVA1PzTwAq5+rr9wvC3IlmksIHMn31C46L83J3V
tqKs0WkyXbLNZsmup/fumIu7JbHynHrVz3JcDEsyyEWb44o8jclIn4hPzzbMV9q1iuwk85Sjpbuf
slLXOm4vxdNzaARRoVN3OAZMDdFxcsPgcE2qZrIBdddkqtrbTklry0znIa5M1tJxBqHNbl+pdoyl
uAx8Vt4fxchxEkYa/ATEIY3vaBsuk/y1dX/R/MSLmwPoQioi1qFAlaJii2VZiZtv7cNIh8cxPQtf
K0XbTZRhyvdC+o6ySOKjeNOplI74k7YZGAbBlAqSg+tB7lIEdGnoplz2GbzUe6LU7Evwcxnht8rB
EBLnGSUCsFtLHSmCH4OAyWEgKKKmhQP6WBRy6MRY74rWSoajrX3zY4C0vOQxvB81FQ+mWfdkw6pa
GGuHzegKGPpGHwr7lx0Zb8iZCxxiypfinr7fDKyYN3+cGfFQu/2Pm5v62AHzFsHcbv1Ue/FSAjaU
aASjemgWChLZLx3Dk87pgP5aqY4n5r4w2ELNynLrS/04aeQMBY92RXXEfd5dK443ZxMFMT6u/SRM
yEfPTdGPp2zLhnlJTr/b5f1JyXK1Ld1qq7HS2onr76nKWIgDrgVBZW3sgEIRl2vNpj2l+gcfNcl5
FcVjy9hawYoGlPVNDU+Q/cfcbfImJzfqSORZuPbyYz06HIbJLzd1pfX1WIjy2ndqcttpO6+1+yDZ
4cZRrT1hvi/QpPSRlSddaeaFjTUmxPyhfX7Ylc/k7DwBgPONq06vB3JHH/RxrClFbsKzHUt0nHKl
BglKTZFFfq6o/gIPes8shOdQkBoG8590ED03LVYSnzFdTbw81ZL6WcLa2MEZEHrx3gqz/EBdUiKn
iTEa+lq/1+boSIrjW69eopJC+FBDqFtjLUJ0AwDk6aS5t1WUpt8ta05vd0Tr+FcUO/1kXPniOrnF
lIXpIpYh0vWVbHiGs+lmYgGLwvOjEZec2+O0R3sI9ArA9SEAdFnVkQ8UDTgtpHP/YH+v1blSCo2y
pSLNftXTZCuWNjDGoiwEmKrgDe6UqNw86v7SNnVgOJXDJos3pGYsN7+sF1n3gt5fnMIkE+88ucLa
yEJUI2qFi8URu9d1Y9R1UT5WlOAE+g4tKmd450odqK6gpwwX3osYwx78WW5MMMnkQQLKQovytv/5
uNjwch6bWNnHlib/AttELtRT+dcoIEGru1R4Uvg94zyJxca4L3PDuY28Rmj+xMLfYzfWxiDB6JLw
UH+WseC5jeEyTmxRHJ308wri1kkwcnuuzMnOnWFtRUYe4ZaVm01g6kRXT8H+kNCsoiO6qvepur4l
ItehnY8Ci/1E5oZF6S3YSTPQVCGFcMn3+GVTTvP6pXLXxqx0O8Bl4nmgdPJIiagqhDqDtDVMiK78
ElctmMAFNi/subOxtNTlzjms7mtG8Vm/CsgOecgYrIS8B8UdaFtkAxkdgmrt8A32MP+99thCfXgR
W5fyafGgKd8rAPlujpxSFoyFeYYmThqKyHklPPLNdiVTH+z//dfE4AtYy3zUZarKGZdRwsrOZAMw
yO2vieboiNlMsZd9HUguuhRfjjIwYCRPad4Ym9YvgfbBlPcMozMVTX5rLTlSOu+CwLtFREptr29j
PRCXJwid42OOkHrgVvVErYO5MoxLRMyY8yU1s+nqm66YjThT4vrQdySYc5Ztc/eOvVkOkJ+V92yv
LC7hpdWiyz7eJ5LH3I7yaNv2Wsg4ugCkzne3dH8fu0wPHRDn0QGZvRE1exdd/7/LcfKdegFK2avH
ublsxiXnZ//VShGbm9wAyMdydrDiT7g2umalLizklna1K65gpHdm1K2C556O1kEM4nTLhq0mqEUn
oBz6Qnuf2NIQQ4RBBzZP9ihQbl5Gi749l+ukFydlZ5I1+7t6j5xaRDZ2dg8o4zWd7Ts/IK6iFIBo
4Zw+XQxcBVsnpYTyh8FcrSrykxb/1agDoqqmJqu/MnJoYbrm9Z7nqC258sFZSABV5HGYmGi5ma23
gKr8A904btRPDsJycLe+r8OvlS1dYNnpAHI/tD+iMHJA/kCoTHy3oUCyDWwvO+XC4OPR/IqJ4Zi8
ynJchCebJzyGAGuUfH5HL17wii5Oq/kiyB/jM7FnJn+dkVgeayyfx20Eyn+iTfydouFDET61LjQJ
QNzH7yS7lO4R3GDYGV4SEDBuUoTtXJyP9YdC3RBdNWkbr3ScrCM4YJdczOhe+3qzh4bsWKBVIfFc
CRnSXNMlNDWuQ4sOLDJEfXKBBSUlp9gnog9jQ7dZtIjw9Q647APkNoi9w9XwpXI0mo1rTiE4SZg+
uiTlP9t6qFrelUoxkVbTEJeoCebtEMX/veuvujitunDWqg4QST8udoVO2Xdh0iyEGjBRn77+ng5z
JUhWcKWC30BJS9vgxGJrAodyj6xvLL1juyESYSfqAHgmgF3SbDuohR1ev6yw58brUS64o36LUDhJ
TuY2MQNXrFhoVv1g9JkCR5nonAE+6EUJMcOXbCoNMYYw5On9mJK1P14f+dTMyouQHcC0ZH4P8X9Q
0RIZd3cfFbZiC3XimctmUh7gXN6/px8jzzwq3SLqEY76r4qpmqulxL6zZePseAH+OdXLhPrA3kNj
l3NfJQPMMRcLOfxledtdPFinSJms9VqlDh+Tc3yyDo4uSqHQFY9Hvg7w2jF/T2N7N6BBVmbIhFng
4LPg3YwC7WZKmMj80AGj6zAKxDvVyCm1WsG6sBhIZG9DGL2vjbQAGV/xg6IPsjiW7GNu+e/nVHFf
bYxWWnB6Z37HPixjcx2v4WS7BE5p8N35eEaPDmPJB1IPP+0/9bWyVIl7DZlCr5EAaZAzqiyUnwW7
I/iTQddmLzgJTP7oFLGv3VSAcF8EvzvkSYeeoNXqio8VYlpA9LWMeZZTpxosjyINIkxE+ORO5pnK
QsPv6ZHBJpfdCI6CriW+tOFdRs68Ym8r1a6YLKzuILtotDrM9bZ8Ef22n37ZJSc7+VYazZKqcrHs
rn4YT5w8PsO8u38lSp92mpPmIUBgoE7BMlQdzVwdpInLpV9pduRhkrqD4D2dYmyKfIJkGs3BKHko
zuDMndJXS1bLZm5HTklucf0XeK1wtQk0GQsZxyBExZKH/iE8uvXjROOdSyBn+CCB2wvEbMGHCX+5
4VXNg8YdzARbu3hfIIoPbPyFkgMyBVRkCL5yvUi2aA9E/pS7JqNf2pNsnAEn0804SAEw8z0uDmbC
uREiGQsegPGs6YtQWffXnieWc4saDfLffuZ4UGXQOXeIAT9xGSH7kDoy0zeBoVlnmBf9fNKlwp43
NnSKDf85Wie+wADyUi6f9dxL5L3fJ8mRVN/XbURmMyeuxB4Pz9QxG1NWMF4dJ8lqz0XlgawxbjxP
o+bSMlAFhq9jDahflb9/YzTX7vSDND3mHmO7ZxicC6OdNBWFMOF1JKVvieUaA/kElEBVO5v4KrsF
UDvFjiVQNTzBzO2QrDU5xQWxJ7PplWUQlDmUEkdvy+xCOgRcbfWd+EzJSCbBQAVf8fsRUXI0FP6t
sKIC/xt3zxORGpJIzLennbMJ+GA2peS8zEugs/CKzYk9OiFFUIzxjbascC417SGHfAHhD+i+j2CT
WzGX+Oj20moAF9IUgH1z16+lMAR7Lych2+BRYMSy0uNq9raV2chZd+PEDLU+Kh+B2bpSCV+sPKqf
K5aFbRA+lnc218HDE4qgl4k00DuTKZgySx5QKs2+CDtUHdEXAmwpeHo2USPkvRt5XcYvaYppQ0jg
AjokG4HMWSiW+dpCx1xruHxzRlX/9gxGW8FUqWnKSzl4f0TKKJP+Sl+EU2PTHGn+mLhG7NFqPGsZ
eSSUFAOswvnR2SYS/+XDrsPEvQ7tMe94Vw+W6QSjOI2NLcTUcPZr8Oyhvs2diviiX1THxsLlPU5b
yO0yEng1Ymq7mQxdDXom4B2u9JiYlw1gOnXzMLWxoq89JYKNFL8IuEsMHWRtTnXxpSHVM0U4G55H
8BGe603AJm7thesn7pnre61Nu6VO4X3F+n/Qn5tmROE8vVJubi9TzffNq3uDoyhS/++3B2bRLsqT
QrAXSJU7VTMyQ0notAAprggunWkfQyXGqj72QHwIj/iwe5DSgUB6pPV7RsJ8WFRQAJ3P+akYwQhQ
4c1z6kR+h/AfYQXzXEpzT1W+phlly3eik4KCignqMOzK+KOgDhB78IsChtFeKrkL5dIKynaI8zbJ
n1tgwzHfqOwL1A2ecpVu1UqpKqZ/5OMDwmQPqb+oyUxuA67oqMGt8Ir9lUzsAqhIMg53b44HQtGU
oHEJ7kqKLrCzS/FadOc19b/xaKparXik1eGuOBF1MxkEdG/BfRNLcNMV01QnOResfOIvUC/wzYe/
VObIMBpoC0uQy2t/Dvgi8EVsObmeHbzaD1hJ89X3+bUBwDpQD5avDYxGw2EbwAfOxm5fBvUB6FLq
q6AF5yqJgdPxqVNTIYyo7KbXZCuCMHU1kCkitdeUbXlAsGKZ+Hd/NcVsetm3x8whoTsolTePTm7E
7wIPdYMeh9irS4u3BJz22mmz0JF4bISmS7PLx0G8mOmw6oBJdqJlmM2y9Fhx7y8Br0IUXtVUGa2s
t3oAUSXi3gavg+iezoLkI/ir4GqxORlHjC0bRp2I0uqCUsOad8AsY/N/zAqtShQg6Xdw29FCIQEq
poTL4nvVXMznScJdhllsIgw6R8JSnIEvr3zxie7DackDTyW5Ub4hmVT4FfM8+bS8mtOLNaIldlO9
5VdzlQRcJxDQhNtorSuw2lF3vSUQCtJZn5h1CzfkC230x242PRj78cg1HkKCgZRQTkYnmPHsm9FH
trTwuzeN/anjTxb1jCN22aF/KlifQIOmDJ/CVu5QqnNgHALp50xXt0auZrym8312rdHOH64cy3V6
oGVp4s8gXeycXhZOXjk96D4z2+pj1xOmc44YJBzc4LLi7H9eHK0vuxjrWv+jHhaGVpoDyFCkzGNA
C9LSTEETLpH0F1OdbCqy3mAH7F+FlACR8/hk03xhhf/XDsj8xCOu6rL2goCntoeo9DKvEn6hcGBD
8O/FtbJt6Xlu82TwAbNC63uamfbQaCIAbR34FilrKbPPc2J18YUQHp+P4SJF6LAVA//A0SLOtmfw
0TjX2lagaNHPu60zw+IZSKuv+/FQJHYeWu22L1gzAjx18ca5csXksYtVZes3bmsOket/fTcNQsK6
66nWekJAUVU1oPk744+PbUbt5p2OWjPznopWIkofP70BUAbY2pjsDx7nhtPzVF6bGCY3m5yP6kKJ
TNT1U1Hd+u7KcstrMyWS94xK7GLxdnByV80md/eorOXjZhaNYeJrGnGawU1eyWC2rUYNcE3bhMCE
rfa3MuU31ZmHQ0qdAGc0vWLd/cOCos8UmLxmPSneZDn26ibcuWo+snCkX8hJfG6eHPmT3fLSr2Xh
5oaKVZRlXu1vCh++6h61k7BIdTVRdmUYkv+cPAkimSmNt9u0/xCKI2uc2WVKbGmUn3t7UoWnNiV4
jmuiYU1HU9te4P4x9chURIV1dVLMiivxlPB30TjQmD871tBWfIDL4yA3rwcEfPTQPgjiyqrTg0A6
VjD+4aGspjMRJpL7OZpRbEZKqntPwVkCri7uANUA041d5ZGVnW1eNrhZsIKaqVSR283jn/2Z+/Sc
IYmw67uqzJhr1lHPV03XvztR3kj5OT4+KXOOoUaLuFPmM6FD2l+vReL3oFxG7dyo88y55wiHWMlp
nMrnokbRhm81iJLMAkiDv1K488maw7IbHewA+q5lGLep8zMXMW2qWnK5uGEImcoqD3yOWeNB5Acg
o8d3vozpxNu+nd9u2VB49wVC4HWYhsu0xtKYHzVYVKhrUOqf+lQ54bUvctqfx467G2CW/BXNOU5s
oKjNgcuN3fakU4uq8Wxd8GHbT3pCre9WfJRQe+GuAQlCKYQ05TWdgLy4tazD9yogJvahRvFVpB5C
vD23vX+oVx5UUj3t7nwvUp30QTWfaDnPvqFosgWaXfXFKV3PFGa3Psk2rWzaerkjQ5tfCrw8v1iL
JXRGtzT/Fgk5B77OJequ4Uv/O12120Puup9DLCO3NPv/Sgbp9nFKl29Z06SoeZ6QyHKpVxQRDuAu
fSGGn6aYFjWANfCBK/FjZiEzMy3cph92SWrwx23hD3R0DFgihrwm4HSg1qT3zJjHtL40rHcqTJTU
0R+QigP2AVSMAwZ151QROrchZVd8Wi/bn8EKhWcC8k9UVAQ73LoXHvcPXo3m9zcgKTo9ZgQ2PQfo
zCYU3D3tlJVfMeUCwV8xvr2h+51Mpym0LNVadbJkSWk7tAGxk6O2+UFu0nvCth2gPQr6Qrqak0BS
Q3qRngH9Vt4UHtrjOS8bzJm08p4HInd+BgUNRQQ/8GFcN8h6NcxxKixDoOaCHqnvllzMqkECAJTU
bQdteqcGsIeA2OhQayQWEmqTvLatnbi7KxcwaFk0ZGjq0bFW5lJP9MgpvFWQcPb6tuE5Yc3tyrId
v5xZoLyPSwWzxXOpeecH+XGFaASR2m/N26enE0GQChK1UYQB6gmxwIlpqBjxwGadIzpjKFzalgCR
/piB/k7RIIaANxdDLn0WyeFApzALSTeyF3dMEmOg7RZ1wD/xz1yCANLUzV+R85Huz2pvEchGZies
DGADrlNuShtKXzFEEf9ytPbLIRHK/5lpbalxSN0eO/E5QTiBaZJAyIJdk9veswtf60W1B4wy75b6
nArGQ29IP7kEQkSY77yj+7f9PvGcXd1WYHWiDz+dK/dPC/arMGQG1TKXYv97/kYEiWnAEsJq4zIM
xVtPLZVTkfJNQubd+bbhQbWiReDX4g1fnJSV37tlu7XebAK92CvyOrtXN9Bi7eduMg1Ah0dHLoNJ
B6M48wIOx+eCp2j0cYQ+v1zxMye3QWCaOa+RyMwf+QMcjA5XeZL7AhRySVNrFs/FK2YVnsLtoKBo
5ku1uIsyJLaJDmpPXeyNIkzqCNEwN1+kQcA+WYxqLWF6FkSUFiKn9x+MmroGMWtgiAZETqm9qayr
9luMdc1Qnuav4Kn5sziE6yZAdZZlALdMXVMDWhwq0BS5rpPnSQH9jyHoOQriD2+xOqepYmRAkde8
vPxrTpnd99bX81dBxp+BkiY+eRt5IcWDbmMZGcFBb4QdbVAcs7uZ1W2YnwFUtwLPlX4GeSLk9ICC
JcbXI6zXWeIQ1EUaFu+WDZEO2djbiLgxTBNPaF7AlZSFmdKAtJoafo06FhXq4JmbWWIS3PBc62zJ
un0ShpWovbGQi56WdDOvzr48q2kbEdVO4zFNhgsETD0Jsp2Z+XuvkFMgXSd4gwzQboxCCLbW6CpT
UIPbCcDs7UXqH/AQ1wIkJzDcxsz8kejLYqqmb2UG2MDiRsu6kHtI4EggWpd3upb6vomnteWCJAwE
BknZ7n9gzrpNCKVKG+eOGcj+kJKg4XpC5rWmX3tbklNROD+yVKmTThjQRdumha5nadGJrn5Pc7IG
JgWWPA7L1efij6W/3tnf8Y2XKAej00YsDbiQKckdtmo0uC9a4/RhCh7FXTth8aV6Jec823Rb+1E1
FX1OuICVWFk0uF7r4Sm58z8X5ZWpl1jsWdkhP145W/oZm1t+nx38vUSWf9lY+D1fFvLqWEpO5bL/
IBeuSz6/qT5DnBO7xgwfwK5tpMXpwnJIgRmPLTovnR1LVmgP6HmsZqxbif+cHxxwEaj4Dyo9lymC
MvSaSsnMci9e42ih3/Ic4hCQqV9EIPLPKeGsgtZT9iNsywAj9jtWtNVHK2FYIbA+UNmFakfF0kKN
CFkt0TbarvjSnrvWFnyL09u0+UBcr2ypvWOnx3FFOZ8QCxCUyVpuTcBCFrk1rWKaygCuj2hoi59p
0JdytvrK5hSi+uCBFWkOsvhFaResfLaAqljLbTPHEvOFcBCqPP4huqBvGOQPlLxsh26/foAb7oqN
53uVgxOoVUb+EdNVtgxa8oFXHFY5ts9CbOqwpQnuKHICKcAU2nsbmLeSGgjTMBJpe/bEkh7kW5qY
5DOsb1pKuYdgB6z80aR1V+ODeLIR8Ol3GEmddgO4zBgOC39curVzx5PdyB2MSYGXXhdnGpF+Cu3W
VsHEgJZpah8yoVLWu2Vx7zJTMfGxpUk/PLQ34YjQMZaHMF6t++F2H0mrTUMjD1L51vUltW8EPs64
mw0frm8PDDUiTj2mKC+M/3+rPBGems/64ZpjDrujMpIYnftRd5scfFrDP3u6ClAx1S3uVquk36u6
2M+ywemwNea30fq03rUl8/MUZCsVB+AGW4QqTyWMhue8BdWCr7lTEo4YTrPvvmilAdIfSEJDAYMj
mEBP5lCSc8JwFkgYeJuGfDwIgwRSqkaOBl6cxrDofZPv5B2tS/255ACjYZE1xmKGpfmngh81F5OG
swGk1NFUxY/ZWmquNlNnNa894pDY/0f/1wXULl1AtfDNw6skHFXzBO00QssEwnPcmMnCZLlyz6d7
o3LMLQxcRjs0wEnYig7TOEXgOVFzXN0q990xxisWcZTnUsXdP4Ft1gXlu3Ztc2+nayCHVz9lfOO6
otJSPq4uXZCmEC504JAwSS2u1aq9bdfIhLK8HO4vYsFUzJWjQwQx5y1H4+FxYyOpLBf97xwFJG0F
bEQcwwdDv1nhxS9986gO/QRPy9RE6BD/nouUPY8Z9Qqe2tKfrMxtMzh72WakXjX72XWasATPSzPj
+4x/IvoLG5f3g/4I5J6EYYyoefg5OduU0J+TplRwVqJMoelpwmK2JMA4LdttJltNIr/Qrhg/P+po
KyMSqRgMVJAce1cUiXLwwWAF1FdUaHqgzKhu65Kf5CTu2Olf3g2BAY0zCW6AZFan1PXgPAOmCwkC
oiVw/FNBmNR41Ctjl4G3U91lnvJyLmQqxBvSMiln3yGszC9cObfM7abj45OUoS+qx3rKhKCKd9tK
xAPnSt2g+U1svCYDYTasEHxSbRbxv4ZhadZzCvC/qNZM3/8HZwHe3/pD+p00UxwXzIRBiecENi6Q
+s/wyzl4wiBtAC8yGgl0nK9rzGX6gRtTgNDHXCgDzPpJxn6dGMiv+YYRpWLK8btU76LXWjcFkkpy
FwkLjUwoo58d8wyIndj+jb3scQCplTsuAAG8OtKYi8NIX4OyLFgzDrGlOe6U2+ateIgI4AO0P1Bb
It48l4UH0aaqbWRnjSrNU8RYxHKq830zWbYskFu8dIuJFaVIxYoFu0v0hvlO47dN2Fp/pGh6a67E
TPwlbm725Sd50sBLkJ7LECuD0TmlygNdt/mnPWFRCNQTPiGfK6D+uh7NU+3zoT8CYKrg/IAwbkUT
NAhPUxfxk3+tLx+AefVri8F2nlFB3HRqVgYBicn15AdJh2WfJBPsFj1foiB1slu8dMn1a+YKh8xp
GIlbu4i1DaL6SA6qVqAutKQggAG9ouMdCHsc/dPEO+5sVHdfT0RZSkAXvkYTJyF1RjPm3yx203qA
1j7quo1JLt/MUulxvdHClaRZUCHf/SZTbfbb43S30Gq0saGX0RTJAMd9/tndfFJ/2oh32gxk3vqL
48bt8OJk906ezHZSb/TmC5TjoIISqMysDUbO2xmunp+LbrgjCCpp8gFjnt1zMYc+YY+tCTm7hz+H
leP4r364khKbQTLGNgiiut3uuM5bxO9rEyOv5nbY/7XV6ZdDnerhmzv8uXMF1E95ejTdnKRpZZxb
/OFjtqkEk6fDeav4wHKAlVmOCzVfoG2HAclexJDm2Tz6dhIpD4qkfSlJrWBAtpH9b6+EzOW8AfAw
H4boWNeebMHTEfbIOV1Eeiwa2RlDuwTZf1re2jfwPquUbgl6JMAGZRXTmW8E2etJTxNEBk5M5w/n
DIxVGIEVoHSq6mN+Kxh+i6iHE2o+VqlOpDJzZ55OgFY54WPobKc9+XsabQaPGovvVG+nctnMCa+p
HqHayaK6e6C/yjXXL45wc+Zl899jc1ossGgRbHR5llSN6c5DZ7eFPFXyS0VQMccFONuQlVEQd0Db
tVEOlMbsmeEhze9CrJWr4BEafBNE/kmU3YaLBiw4UJFICylCiAh1q5ZtyqsrIN7Tk2Aq0WumcXZ0
y/yjNMFbd6tcV3rP9SMMH5ix19gvDeVIF34B9omWIPGR5Eb8aMNj0qlDT7I2aF7E9FxQQR3hBj+J
hmZBjQwHdkRyQcvqLHvf2KfQWGWybzp2ZNyvL9sfNh72R5REWZcc1GUXS+35wENyosDOnIKLYE5p
T8fEGM9bGhg9iSddoOgfsvRfgxNwseSB7Hkt134jQp90+Oh2RuCPSpK84e1klWa5RR/eMtiaVX9H
yYygILHAmrtn9XQ311jio4aj8/7iFcuQVS2Cr8O09VMkw8SxhQno74S5yLTXOS2YXic5JH7q689e
J87+pxyccbjON25W07oh5+Nr/onMICxIkA3DW6cewxhUczWkLXxNtg36MxGak1rBm8e28Vy3qxwA
fQC3lCLySUwxp4t3HQZLJE0jC3hx+03AMejWpGFKRgseGcAhzoJmodoC3BpYX+InzNg6vHb/eIyk
D6I4xGhniiyXgmSgmt5oUKlrpJf1+n14Jc7Bzorc/4/HRpRM93k3ylMNlCgfmCF7kAmveUddHZBs
dLRtL+OW88Ctt4UsbY3lEF7mnX9LR3b8UlWXpF6/UyWiReJHbyz0f3AvgeEBrG/D7EJrZomXHNoW
dHoRKtdWU9Ky9o3N+PwWMZkDURwSGRVEkdR7dfEkHzXWBghmkipslsxL3+r8Lzlubk7Lm4A92/al
dPidiMuGeq9wpRABqf5AINfft9imbrO5flbMDGEo7Kzc4OYuscPlkGFqlvzfM0okD++7b7XpJHUY
USKsYK4KmTxm8xILGIbpzMuTyeT5cgE0DzsKMTFnD7XT/Rbqwv8BBXuf/cyIVh2tOVNFtddYqp/x
0R9wQQAd/CgFdlsCqDlxl4t29Sj4d7wraUoYIHXmc7wV9hd2DwCY4dobIdNs/A8kWfnHqffM9/k+
D2/4OoEO3g/BNvYFbeOGrcqWzjQaulPa4CUmnOvkKhnG9YuTSuzTqUGKZm5aw3JosB1lnkhv/Q0R
mjc3ngRJLUjfZkxXIdvZJBOTsj7N1uWEhlZ4JYbiGDdxCtC5PXsPuNVCkANT7v7iaUbe3VFGEMHV
9O3+fNm3xXRaizkkLz8L+xKYAINeyQdMjK/2D5GgZtpodvgOPHKi9aADRq7ldPKxt3ez0lygavWZ
djD42XDCmEE30+HRncU9A1ZbxzBDkoyuwC4wQDWy4aNMB3Qt2jAZgob4dMHZzuIsbRYJf0l/bx0k
VZNgBMKA5zFGQcyPuP5GGtwOVw6V4BMLHnNYT8EiNI5qZaJWOVG8BTS3xSMlNZVuhNibeSb0ww1O
YNVaMjLg4MH1fkSDZ6sfaOqjJW6fsdluQhujRbt9AWXUP9jwq/d4UDZHEIucrbEcBj9R8/NC/SOI
bN2f87xNefCJmbPB0zAGQvEuH4BMrPHYxoZUVBH1DqNavxH8SKtl1oF1BHNmBZCFsB2BwzwpUIRV
rJurBqWPx99IBsU1m38OQNLkLkE/RojAkav8Yst9lthpbrmp5WJ0It27htQvKAKWS7hwfoZKBslL
2II1+f8B60aXE6aGab7hNRqFIxF3O60hvwrOMMQpITkV7uggkYKbqHS6AuOMDf94cAR0XAbckaZR
VBVi/rMcLX3k7SqFbCKS5gOyjW8Wm4mnkg9f8E9Ppigp3Kq7WbEZ32nQxanbE2VzdeGpTVj+FOaz
pgrBzjkQzClYbHznn/n6bhYlPHs6FQ9KVSmlkrGHjUv0mL7GPuFul+D7To6iGhUBgty98JgnD4fv
TySihR8Un1Uhx+0vRbT8Bbumnhy25yNzJ1oNGXwWu6p1VkBDjwvfqfWHjDxCP37FhDwTX0ZZLNqS
mb1M8qgbvot5n4NAiPPgV+9TTjOOv+QEu23mKB8fEIEjzs4fDvI0v/WeEubjpbZ6WoXvXK1uVG5f
a/l5S7N53tfRAAtnLTw7+FyWwyGTXt3dub4tt2Hq3oDYdA6EPPTJRBt8OgI1n6y1pt8Dn1vn1+0h
CnOcDBHciKDKoB8+Khte0jdC2el+Kwry6Jlvk2XC+N+bvPfuuw/O7sX6P5zJC3Vl8TZs8cjcDxmy
Um+TjmHQUy2qzBudbgKfr9d19qhTP2rRfzfDrlnebwRypshNWXDcPmIg+mQzG6xClmVKaqcNzq4o
1SK0qw896jn1RgPZL6RXxKa0VNywM/3z3AcfumIVrDgpONc8vX4f7Z+vLy7xaFCOAmrpInX+hnXB
YhTzUG/oMc7TKpiniSyGhttfi6wUA5hY8y+K6iyJ+DL/CcxSw223kw50zMPJxxD+R4hGIxXSGg/w
2en0qFdhwbo3v+QdGE0XtLgiy/Btks64dZ0z7CXzbGlHxcdjj/rkDS/ilyg0weAL1VyLB8ZWy5hi
FJbfWtLFX+cf4Wq200ZJgRjzSUHHwdsmG/bjo/kJgnvXJKIz3UHG7rB/FgUI6BGqvwQVZfrMagLM
4DVmW1JTyWtHDVrQWz+xH/ppChMvWFY8D8cylbEypxwE2/GbIts09IHXPtVgZJIJnZDXdbUuz5/Y
OW7WfFognkMs6oAyh55y9W8vKOX3ZYVfeyFisjQUZ93CPZfB0c+QUVdNp8SSKH+M9swBWwTXSBQj
X01taTk2srCymoLGImxy/9vbTuhy020NTncgxOKz/AFDUasJC0l41Qh9fJFmosUIEfHkaRD4Ey6h
gDztF7ksGPHyL3pDwkx2nJ5tjpHN4Ncg824Kf8LXmonbq+D9rl+U4zw15yET8BBmyIXyVm7s1pEf
TG0CYEQBiAnMQNzCEfnWB3m4ALfZrDWGCGhvH54UVFRH3KcLHMDxKBNbobb6Ka74yAvouju9EUJ0
InmccSRgysRgcKit/BZxouorbBCR+3XuQ/JKStk6MZszApdX+duZVaR1pMA+rByu2xl+haaKrght
1VoCuDKpuV6pMGJFqkl1qqjEdWwIN+0Sw+WFqGkn4HrGEzbY2ZUx8QvhFykYMwb3aUxlbY3nWI68
GIbNPAniXIBI4EITyYVec2Ol2k0oalnnnJaLtC4u36PYhqUwupGK//sL9uDRR0pI/3Ee6Cj6h1+C
F/YM90nE+Rh+PQ+jihVx2AQ+sH0RRwIIV4xQ1XDFY43hlIaUNo26XRsqJLFNeMV4eW6GjSavGM9g
Hx3DT4qw/k08lhYnJGx7Jwb5jiqLPpzaKSG5Qi4d+k4KQK8fVxc7OIuiwrmRZcfez8xrkT/gxQ7b
ZfURdMfES95LJtDMlXJJmKk7kIr5xHxPTcnqa8DwT2e72FUFfGYSwxL4VLulKIuYivceEhKHSu4J
XrRGSh7wMv2IYqHGUFYvJ9xCeC1qzw3oCbRKZJFhrR4dGQmWycD4csaJM3gKKXbzCuhkALRmdnum
GZrKhotI/VmC2FEhRVGZ0LQDIQxRNZ0RCeaiZ1WleHcNuAZQAHsrdPC9TZMyEuWOIdNAstia2jVx
+ut/o3BWYEQ739O6TqAuJS7hyMQ27wWwcst27/I0/TX/kCVSe//Df07s2c/iOX/evST6FyBxnZhW
rCf6fQ08Aq7gznayFc1ckgu+aK4gCdYE9QKqL7e703jY4DC1Zw17fbzmpA6rMdkDnRdk8szwJT7v
KyqpPc8KygdgdkmU5qqbikpE1hHI7YaYrK1NLNFw6sBEClFIzQ8iqa7m5YnPuEp6gWlLRCXwK4R1
WnjEI5bCuaWMlBO9fHZ6sIw+bxBhudrIyQT9nLdjFNSwNko2w1/aSGkGeN2wfsaX544DmPtLpgZn
0mfzIMzPOgS5Fx7AXJJvGBFe9PteDatwxKISfSDKGKPWi4CkHL4nkPvEVI/x6lPrrVwuDqf5Dssp
H+BZAR5/aEsFZ8i9ca9sr2Qz1frpRJcxn33cdDFDMchBLJEEauMihACei0R0cWS4AipLaNggZTIm
g4ok70L7LKGYBnt+KMazAJizOPjArmBBS134trdTujcibV4AiMA8WqAf/CSzaaWWB1fGMqpDiwMD
9MAr6k0YhoPErCz8yE5A/lI+VFyjiKA8WB9SzrtestHFiXEPOW719FZ0PpY2lsk9EGBtCdfhtPmQ
1TNRAzh8yaEw40YhSFH55gAH7a2YT+fOzlg+EEG80kFz3I3Zr6KUHcp865Vw+6y+EBKjJa04vCY2
SWn7UuVuG41FeQUhckwpuFgoWjnYCYUhatzv1TjpB9G9u5DnYSqobKL1sMJCunJzbvsqyRHsXD12
m8RKngNNn+yMq2j1F226+B0PZ7nKlGavIDZB3IKjIp0K00RdDR/yiSo/y00xCcb5XIQmcI3YdFxl
qObsLAJ7ESlGR4OTAe4RhnFzY40CXrUrLYyPxPznRz2DXzBEPl4+nMNzNx3Yynljbj4dbs+fQ9ny
2FQWpv4BEdPyx0K1BsR8Qy+1vBLfVC8NV1YrduBaDyIz604YrnwRDIm+jbOY6wdT2C22fl9YrfJa
EoUcnCxSqs9MC77s9aoVITjwoZe3dFbpjqJ4i+mxP9kWfN5MRwZ0Gi0ga2MY+ueFiymT8HF/hknC
BGCcJjj1r0BhjmqVVwf7mdrIvmXTWFYvD3JJxLu2p4iyBkZgRlX4sO29d18VgZ3f+ZqzPRBMpCEc
O86jKh0S3c3Iw8nP0dVQriHqqEkqRJ23/LtWWUXTBpVpjizSasjryW6RL7TZUUz0iDFVw9gLqsGf
ApUFGxygmmcv4t7XMBXvy89jCFKQb22VMyHn/B0wp3xl0jh+7n78pBIFBHeQahX3r9aAriNpUxRu
ts8uIBvkOiOimOQT49DVnrm5pMSB3kLU8Z5mCIKrvVbgiZwGuo5OqgkFm0w4kTRYLiNDlyVr2wY6
OE5bP8is4AO0p5Q+HGSMlWrddED97bmsVwx+EszgfJ0RVGL2acN/tAu1r/hlebmWEUn9PZXK9atR
VWmwkpnP6or9gCvOHUfWmojPtvlU/H8Y6Bf8mxS/H7lyekhoQYJJLqFDwc3Yux4Rn0mPRFgjsa72
yTnFJQNrlXM5OpZvmXJOYkW8cDbNPuNpg0ZxKSHkKLtkfCRwnl/xcW+Cew16kN2T+KQGgye90wzE
wfndp9SodhhGsC1bsaVqhFXivdn0Ji4NH0JKkzfwM6e7YLPOyAdMZ56jOavsGXwJvnlte+8amH/e
xSm7W3hhfCNRFpmO4NCYYzUY9LSiFwBzyNJeqHDbfjgyglQ7N9YqE/NbCxfQFDdCSTWjIk3+8XQG
L2zb1z0vmn/BCsC7O3jzJYfsIK22MyshJcxbghzigaB+QQG5jJecRp7vvJ2hAymeSSVbNqxi81Ux
tkrOzu412/DWTJtidCSD+2bGACpifo+VKBTPfy5LuRCMRpIl1yWxsTZPjGRY2RiO0/YVSWV0+fV2
7Kx9kIUVr7DUoh2Y/yBkKsy/ew7Xd8rOJwH6q43C/abdhz3Vum7yuy4nG+VAEiKDxgUIJQX1JzWn
ekCyJUaBlvxKWlsuWsB0KzbVhWkheu15i5effNOoxru9wrPYfJz7t6iqS8LgdpiWgcWqd50GkUSe
wrnFuuZ7U/LVu0HCUuDz0aORPVbFtDg3oRDTUaNfmIJ90ORshJr7nGCOJzT8c6bDkht9mar8Dgdr
PKSD7v4KqPB35b+3kOhbFVkbASwdt/sux0fKsH+sz0L8t7aXj40fUsuwWo0RqqfxHOH/7sl+k8TZ
+/DYKH4ikcfqrY6lgD7kSHDzGOFqd3og8it23JEs0SOUsTSBShi49ru3ADPRjRHdL0TV7vmV10Hx
4QIpegshT4Nyx5FAi6qQmSsezXhqmwb8QJSE2oGutxc2HW7eMXUdUQlF7hEkZTwO3kJP92DurDqy
sKqALNJmrFErDtWkW3Of51gem3xl67/CR+ZYDwSneMBVT3ET4RK2SaAWoRIoV3LSIk62MNK7Vmfi
soNULDLvpcfMYq9NTH1zjhzC+PK59x75AY1sF2R4Pn4TCN8hLy3OLIJd+rWIg4bKwNtxqW/s2AOa
S6GZO4b2ICuLV5fmxaES1GF6TyoApEPcAam+U3tuTzPGJdnFD5DJ97PJ6WlqnOuNbb/ZwzlTwxc7
n0T/Ww/vPRzVZms+P6oiFNwFtF0E+sRSDK/kt1tVh8cTfeinTeyfWHcIN6JfQAYeSHiozAuQwAmh
erp2dW+yEx3kvj1YUJ9a5eiGTYEqVKq0j6VfS7sM8qFawxQ/YwyYj9W0jGywoFgNrckZMTUjIFiI
2m+wZggwZG/7K+S/Wd+oTj6m6loWrznv7ZQECjS0zOoZkGsQ69qNXjO/8tInf9RxiMby2qJVzc1u
ZTFS/lHHNqoR15FsbHRCErx5wqdk6btL8nAfVTjx97xYKfB6Q7QQLTVaySih4BkCgNWZlYiMIt0d
/2Q42x7V7e23O9BVJjYDPemdZGF5wjMJ2iZgECLIpTZYEqYE6Z0nKYFFbofPSd+5lZ5whuaGUQ7w
NZHquunX6HGNRfBH/vj8lUcfYIOSVW0Ya5P/9pxIMb6kYJd6VwBkoyWNSCd+BZuhj/QDGztNFMm4
pZ+OEijigea5gOVMtNpCVObIJKgCZxNClDOqApNKdoKPOMrOIQPltg0T5p4+/hmWIB547ghLDXx+
OWloB5MDISIeZvJ6tbcXclCs6DxQ5lMLQom5OruyML6RoJ9oxGgOIRj7on6885QKSOcsinOxRnRI
r1GtOtL7+3q0VjfmS4HQHXDt10YcXD3ARprIYI3s8z0mbGiHGTDiFAqRb6DOmE+KUq+tuPjjjY8r
mtwYFS9OCsfpF7qFcfuAdd3Mtm66CpP2mgh7QTl/z8GGo1cZlNQmUGEiq/YrFsGbQ97aIZz615Rj
8DfAsN/mwomxjwZtrVyZpidY0AOMNbpunOBqZ8rBHv5Mljj/s0ri0B9w4lUFJjsWSkjHdbG4BLsx
VjdI/Lw3eNjgep+kGNBbXAyoWAm2kNwcJWsNWWLdhglPnGNvpsOP8JdMTI9aPiWpfVq2sL/z6Bk1
eMiZZK6cx+LS+clgGjOy1bLZ/uXXYTThiKqilmvTANDc7U//m6V2KrmoNnmQ0qw2wepeO7JD/wof
pUKeqQPIasQSbf6k0EyRn+uwfWHPk40feju0lT30UBFjJrYBAwDRQH16QJzTFC9jOK1e1B9mI8d0
qw9dt6/re3ZA4SCTLqRmnb/gF+okRxPgPXY2N2QhDZcYA30KHC/kFe+v0cMJEfxchaM9Bv6E8DdM
QhwkT0rcYnQ2sP9YTPhHBE1dnXpAqvrs01RkDV1POalma5jV4c59SCnhNnGGGQA77HRZN/B4ZfDR
RihB5WaHsrDezNNK6fw+yLqm1u7GTfKvQerOryl5dM+AkyyzUe+3qiN5XNzxRBmOQT/NaJxQc/jL
4u7MY6vr771Z8Jm8eLLr9+ub5Fd4mDtIxw2ykyO6ATr5sr2ASePsyQKIoXZw4hBo6xd01lQG8kmA
jeBvS8ifFxw/saNZnec6OJy7o9Y+7Y6cZ52xkrZkNZ/EGWMFc4qRHs9+whm3jfrNfabqpUI/yT1o
sn18eTMkuIatf8uTW4XFxq/ZynSpwjNrXTBL1HVIIw9Z+Ox2v7yaZSwfr/uMbUxWUXKGwgshxsK/
DkqFMqK3cZO1G3OOKwcoTswI5Cd4iZdgTczTPWYpS2rA33sKuUaGdt31RVnAsfoLy4exqe8xreKr
Q13cTAFPrlOhlsapSoeXeWYwzPRVtzgzKUuwUCBslnMfelh/F09fc9xu3RC1lYRRb85afoErUgEn
QByXPU+YW5E+ZxDUnqJYyN+uY95bahiYLMy+dMHJa1oP6j+5GrZn1P3EUBjFGPWOe1HU3xFi76CF
aLj3Sx4jRT3k/FFAXt7Y/2udDUW8y4dLXl0ufVl6MlC1i0sSW5JhbZ/X8ePLiW8G+AOw5rSc2+Ly
BMSTpbofZuySOrku6X73O4BzCIEsvGwBmzRuOT17DKkFyqDodn/btDPtB+EMmQKvxlP1OqyYVTWT
ccCtpTu304vMvRH/4RxRnoygnvUAoPfda3y3GHJG+/YAoBa6yuBMhXx9LrF1x3CqSPFnQU+r92Wi
VL4HGuuhJdxRPIQQvpWOyE2Ou+SJpX3oh7F9jymr99q5Lq28zXrFL++ctXfXciWX7qVllTsp+OqL
0splMVKHBU0CEQMwfncp9sImDK/J2JEXNjObeFM1Knrm55poBvPv8uQJ3DeDAnLvWxFmsfdmDWIo
NrDspVl8eeZixBI8N7ZbrfEaki2qLZlr+f+ihuBtBcIeXonmA8qqyBBklysI47JvSoc2qfpY4j1l
KEG7fGb/HImlp8tTv5MLfY3Re3vh2vFOr5agjgllYpgiluLB7Pz9W7fVXbbIqGo3KhGjigpgd3t0
lcIhsnorU9mIg+0bSI+GcnCkAPhdj6im1BapEBGDqHAmLbzegS91nTAFIscfxEiPXLKu6YlNqi6Q
ukffZelT9tlky+uz+3LjFFoYHUXI3IwZld7vyFvYlKe1JQC3lkCjU3h8Y19nDsCoaqKbhIjXuaqJ
6tBJSDa3ZSI5dly/qduf5OMMFO4K59hlw+G6/5ProhX4zsWquN38Hen4UyIhAcPJmm1RJ8KUtJIj
P12a9crT4Fo49poyIO0MKHsis/c1w+Yo0zHBWXwzx1/np1E0AwQos8Afji9XEA4eL3phq+MOnLb2
6nnDAmiaDPAKS1dsKplyk1Gl/6tN+1gqQpWX4Dv0J1vGGkmIGDjliFZv17B9T0Of6ZLQxi/SR17S
GfbGFuneEMwMLxaAeNIeTsi3/m7e9Rz76NAcHL/PxblM21NfVOJChFFk6+hAozsv4v6dZB+/OTPI
WffaPHcDPYz79gB/m/P1COM70Z7V3SKx3BZ6qhfd4cpQFjMZb5IpDzlpUnPgjYAdt4iEDsTnlhlt
TWE5XQlSuw92EEfIoXfhPCXxr/BZMH0UYDGxtcLXZQk7AO4Ovt9DknmmcQdyPkVMi5iudOv6I7ys
FuabdXgXxpy/fvWTA/jyAOrYTyuNR88BcpKWTC/7MEZ5xbiCoknHaINd/2RdCPmscTCKh0t0I99u
O3hlsKmEEmn9Xb9J3Mz2hDxeP1SQAedg4rS8JZrHP7F//CEGnw3USUsbPfUBHaMz0NHrBcGaYQlJ
GNG+knT5eYP5qug2Oh7XnSd15T9kgUD0nlkdeY20/UKboUGdyeQaUl8Aah7NuePZTtGJ67m0ucoh
oqXZsCLNWvBbg5pHTmq1RyldugepgaGSwHJwbOJyVYM9Ag/LXULHm+7GfHtGuUqjHP//Mu5O/dwG
u3ahAXMq23gnBJOzEEaIBswtAiEEgQFu+6a9xIoBVolu8h7CfXVDoN7GJg3qNA9HzP8MIWH3/UPz
zuCU5+6FvPKD7HDJcqKii4rKuWL7/MTLz2mpBPqVleSft8Eq/NMv7W+zx/s4wWEoC63XuCP9FyV4
kADt88oVRGV/XLzLMm4V4vzKhJT2sOYQ5XCKR+Y5vQJpHAYCdUZuBLMJXG4pXbiiWdR/XgL01IU9
IMED2TUHWx2MaTDbz+a3sOWAT6NCsHTTbC/mbDpBgMZw21BpAg6uJuCx12rZGiDxX3daCwd+akCH
2cYDcrFnO//UiPdHMvrGMeNm6IwWYaa1b0teg+ETmRP5LMzYIX+046EigFc8VxLBMUbnGeV3AbVF
RaIbvTzNn7y820Rq9t1zRk+ruCqn3I49qF2x3tInVe0dqB6rL0LtmjT6x6y6ROfXEz9o/YKMKSUN
C9MgPyOU9074Q6q0aTPTO6eYCz3NuKS3tjs9aAVwMvG8B0FyX1jApxEo0W2bgtNLqPg3Tp7DQNSz
jI5+cPsw880n831SukhdAf+CoQvYQZ/ta4r4ecpoDmE/Brf3HB+3uFnoHLpCHqy2IxCsykrRHGAx
98YG22/pExet1efD5eTQ/fktEMf02TW7OFIKJD/BU9qKrbGNXFq5EC4b/s9KmUtIJw0m2ijJ1yh6
k4+86Gz5gPrAh9lv7hJeSpniShmm2vYuS+EQHtzC8O/XMwcvB600QlWYeEO7VcgqUn483FafrgU3
5gh+yIWviMqu3bwhYVaJ1wDsEajrJWMo3grJLrzJRxTJX9lZF90OLHZpwIar9dQ2QE0MUdo5Tfd3
tjq/dZvPRp/xyNpK0r1/P/+pmPtR4gA4vo4O120vKtbFCYKjTiVRCituSWemrO05f0OggCKTtggO
E1WkIZZWs7GvDP9m8xYy7pPtEhdIquh5OG2KknB09lWzDY/xQ1z/K03NDDs35Y6egGB26YQE1TBO
yR+YT5kyz2f/zIxWNxPwgNrFa6Ec32KoIMFR45o7RHAc8oQ4E4RHKEufyMvjR8rS50YCAG3w2ACS
cxNVNl69vmLNtiZrxK2SDz4t8c8s/yQKLiVzjRI7WuG8JHZRwsfW0PgYnhiEnLUYlvsxks2NuQId
xWHsnEZSLuUeYheJcZzib+fwS19/G0lBlA+2n6yzN7OGUl6BoqtdXQJsQAB7KTr1cPcmRl2YOV8u
GGEvWmQNj05kwG7SxiyT31MmCGCBU9j7Rowb8UZKNhPXyYxg6+2/eZHcpEym9hlr/DR3d4NreYz4
9iD//iVE9qHZl9WHeyavw0lo+CXOp2tzS9XCqLIcjg4Ithudj4JHhsvnBNEAQEa3uC1uyYefPMJN
pI+ArdLHUO7BgZoUbNzs9L91gslJRaE4LYj29K/l5hG7ans5sJ+cz+0lFmlpa1mZnlUmKmiOM3Z3
AvmDj1MJ5fe5dY73htTcxIFbEdSmTfrnZros94l5FJPikyLs9KUYLIHlIwDhwWLUCf6x4fNiZavE
wSYNesz8GkH8fd7tgR+bML9rofKELF8Kn1RyeBD/90iwFem39WOJ21/vIh4ijU9jt8hQ2UlcpjKr
hCe8f1R+bt70oesqGlqrT/vqfxr1aeuqTIh3Dni27Ezl0O5hNM74oZ6QeCggyA7jgIzYhkYqyVPn
CKuoJ0DBHeCoth7UDJr18kGqlTEi0WkTG4vFH9PNv+pnGbMKKOY0nmlSFhjEQ+fWkFcHaF422J0v
WSYVNMF43dGHfLJgMEwNMuzUAyYlDeqLpGH3WkvW/N0BTbOe9DsKpuSzgvrtJMlp5BH5qaVBN3Th
VG5WE6COXmiv8yiv9j3sqZ3qa/h7wdNwp6VJ6o0qEmr+ZZ4CypDhI6a4Ix3Tj3LLas2iBLPt3+YD
eNk0ysPSoy4xp6si3Kb2+HyAE+w0VPngW0v2pZ/KyCaDP2EctoTuvPu2MNAiZFmAZ9kCNj7doP9e
gGwvMEkaF1iOAQlG8zk8R5wCiQ2Y8vyA9gH4E3fONHr5CniXbe/N6qhFGn/LccTVgOQGBYDWRU1g
7BMM4r2TLJFjhAkSp0osmDvJM98FF2CAudwl3p+6JH/eiKT9DH0mWDG9QQkmzwU7ZIP9Ithu8t37
AzaUSBfU7mVed5yv+mIatORs0wTtRoIsuRRpUWIa8BrsXl9gxke3atZYL14bAhfjhsZykDUEugCR
/G4xxtQI0Bawgtf8I8yo5kn2FKGGl9pCDL48RHUf1KX6u+Q+3UOc7ZqHKY4TAhMwcmmeiZ0eJr+R
3P8ddPY27joDoVJbOx16GfDJRa4GXd9p43F1YHst+kHsgCuaJ1QjtbyLD+Wjc/ebcGhFwM+QdPon
ElRTzSTt77OuxIHJnKH3MV3SpSoqtw92g7FykVQaeeVqTvP90y4ux+TxCpDLpp5l8XaEoeTMMi5g
xLK0keJ63YUXWscg4QnldBlvmFl5cocp2Sb/fBcoz/9RmO4jWRC8pZQg6c6eb1meMGeKecBcTddT
D954lkCGDHKomyxavr+Z3XcyBdForJ1Y/cYh8V5G7DkWqyw2FMF3Jz7mjj4Zf6pGd+oiiYIpx1DO
RnxqYbe+orDZXQbZA1+RqMy5yUJP/LklTvxxlKS/zxM1cOMjQJhX0EMmEQZhrLZp5jkwMWngXXtE
6a/iv1ZGtA6SZR6FVrv88YGuZ4pc6i7blLVafctpl87aIvuh17SXWwPo1n7ONicYxrFS9vg6FVpX
CyL6KayYmvb1cPIPxvpTq1f6PTFIIKn0n1r99gUlQLE2yo6G2xlFWA8cYy0UYe1C3ID/qRkTMwmS
XIU5NP8oXRLxRqSMMuBpe6lQEtg2hy7OaxCpKCjY2qV4s2sScR5S4HbFNhtVk3ccTvXDLiwnTuHM
QuEaYRxexvSu72tzB0l2J/k38UpOr7UrgHLgw6cJIyuIWRPbH4/pEC8zA7le6FPU2eYeK0F/R9Yp
zwqsMTIu8f10gtZQFDGjUF2PL9GxuNhogY/NYX2gvWrKcGFkSE1xgFikGeMAh5qBfdRc2ynPUzVG
Gna3MwyyAe40dY3s8Kl3e6IApXEKxwzjn+97SW1Qx0ibd/4OZpPSheGynkiwTsqNcctg+NM2WWIt
IUg92gDra0XMyqwQHr3YuabGC3gJwiqn6HdxxYiL++SwQbMSdHlvsNFE3caZ4PKtXUcinh6vAa2E
FldyDYS1HXgUFBJnEhPIKxBKkodI8FIi/fuVQqWArWw6fLUjQ85GOkIn53tgQS+TG7dTNheDHN5C
9Z1W2v3RkI2feYXP6Uc1JjgbNGoM7AMcIfQQVa79PuM0THnxDESDY3AuC0W9VWvBEAsiaYx5yHOI
kKJHBqnypQwpepzJPL7JX4NYDyccSP5Q7o1sTCZCy1x6PRF5oACRbZYCycDW/Yen5wQulp3l2AOW
sIptrZjNyN0GGupSmB0/3ENWIN+CYUH+C1Hp7xhkzqMX4jWsJR5NFofek/1KtqiPegOv4vpF0l3I
my1jkSB52U1kbF+G2Ykr12ZI7qLbJw3//hyMkrbXKeGLmX6O/R5Q/z0Wm2qZx9FKJD6MtyCEeSNT
cbrA1yVqhhI/duUHgT5YaUBkoBmhqqk5Uti3R+fB5U2fb6WgmczIawmYDgjNI6gPUwBWRwzWoo03
jAfhuvt3vby7nskJHB3/+sz8kZ90yHrJLHkaoRB7+Spi+f+FB2wWXPbOWbWKx5PDx9WDD/fZdqYh
DSQvupDtgxejt+erjsBQRhz+FPSpGzT5Pi6/fxP/vHtIcu2cy760NEgEkdJYGtBEIWKyhaIXPoWt
O87/oQ4m309/rhYytTHvvnVRwtbwpeiqWaoo8eqt9+hcFY3SbZLw4+5YG1eDbeK2e/UsjwAwzzxJ
KUlFvAdmkJdOVz9nvUo6A9ukEXVdLWSDPKC0QwCXchCAdyu6cGbzfdTt5MqxaL8aoNzK4NT+/m/9
6AmbRp9YYBSNcVhiFo8nYL+/e+yUOcLhzKpAuA9Wq8Ru1IwLzO0/nS4dUyydRTO6CddyEEAugT0/
XbhzsWkP4JNnCzBSsmRQXh+UKC7VyPF3kqoNg4ZfdYlsGKnGta5TrifeL35jBErk4SyUt8S1oYM8
njzkwH2a/NPfENcMq5Zon9Dv4YLsG3Z2NEr4OJW2ZfVjY3yAkF3pqJo8rEVtzt2P0f3Fb4fdWIsv
BMqUxxEkpWMv+XWudAqGYzcLoh3hA072USmthPVLgAW/hEXR/2jLute2RgUhfa3vFh4HFK4Fw0kd
MqhCGOhyAvNzIqfThhYVDuAbNvm+tuQQGK8CRE2v2TQ8bGLEnG82CpD/ZWJhkIh26zjzy37CmuMo
VNcF3dK9fhjf4R7HaOUlwACLFiECSbQXEjdCRTzzQk7NTZWvDgqUQglHHv2d9EC+q9cd29NFNeux
cgug68tTCPxaYap3fCfDuVTQrNZrJeb7Qwt3Y4Q/ZLoza9WqDvUBauJ0cazca5ofWCk3SomUEDCh
RpjbXa9VvhNJcmXJRvNaVMth7InAexVRo9F5R3tTSVETQjntNALLWy6V/sMCuiCZJPvTcTl+SSCP
I0sU+FTmYNaZ56ksfHrHslWNUz8kfBjLMybHF/RXkgrzkPCf6cjlTSbMjmjPhqNwSq1gDzv+L5/J
P/ejOINlbGxKdMlHG9EPa1m5r5rTzW5XaH6YkGQjUWFsQVuBEHd5uxbZSe9eyFov1YVmu4IwXI4B
QecETV8aA5kvSFmukRTgelB/eZu3y2DI0KJ57cUh09L0WtbvhRm8TuzpiW+GpPvcpEL0EQO3LiRP
aPm+YhBdX5eCtGunhGui9Ko9oU4fmEfybmdN/EAfQIJY0EG3Nfa5Cigy73J6+M06ze/dt6EnTOXJ
52qgTWK9iO2uV8uFp2XnW3A30/nb80DJXa9xXu3M+qbkwmleK96jsZPX4hjNByHCvVvHtU4fuw2T
clvH+p6McsNhBpavJ1CDVsC5wXtU/FP+tzwhLAoxwKuNxzVv6peY6I7F5smWe18ksT2D8XYG/gJX
mEm/SrZG/xXw2w4kMSCDMpC1MHMJVTzuXK0px7S6Yfzq26yMGC58A9gMcSh8r+AtYQ0yS6hmn9ey
bLZSFB0W73EslVL5RX6sL8bpifk+2gey2FM8xo82Vf++llZePZkIrJVrSFGEGxP+r5rqqKkC/5Db
jQAW1hVqO9Nxr77CNCB32epwuyKiTALG0RmEZ3ej7ph1Q5++SqNxPyO6jEKujXSupcPwU+hrbgZV
AZMWZ/yvoRNgCUdRRlivN6qR732lBdp2ixzSSbLJm2f9MZQPNSf3F38fJYPbmQ4BaALE1K/dhGFR
BxBViNG1YDmicg3TbQdafSNQKKUYn2esHlVzfSStWd1kewu0GUgT2ccBKzEzfxEurjdjTCf5vUJo
rlbs3euoDME7xARk96dmqyLlz12c9fnZHk1iYYXWctxxpWTuHAAWD3eL0ZPn8cNQYYDWYByufvVo
1zgNwplAXMjo45WwQeek106o/cBC4Bd2LNM/3yLK0ODxLjzBF8mBLyCnPRjhwShkd6di5TnYx1Sw
T0iq37HAafGm3ZI3XTMiPtU9wbP2Jt6hnsbw+Hebz00swxmg2bmpNpvjQBp3B4NYntblJYNOmp+2
mS6WZhiy+fRbd8nvSG2c5D0sixI+hOPKpFh+jO4+krOcff/95FceH6PaV/JN9C2xbJN9EjaiyWz5
nSi3l19H/n6oNdW3qxmkh/mtYCSHg7bUwZRlt4FQosfe1YZLJDatag8+Ip7qeKwmhCCe9IKEjdbH
jLkenUKI0GNb+HXO4iwuZgKZqEDXBOVzZ5KbSGIf8ki1H88n0eV+rgntH20hx9l0XOq9zQ/ZyHfh
AXuutQbPj3YMgSK52viZSjaO9rZEtfSxEHsoKkT3i+FCOerx7QTHP35hvcj5t9YKzIjEaqhGM0Q6
8AltOVWcdGbRDMFsfRDGMRYQr3ywZvhAwYzy+nD7pMlVaCsFYgv1AtmZie6Cwe/3NDMxkw0Uaqld
cx9gle/ULi8g1nTEMSRCtDK1gvHDO2pBGy8uCMdfUioRDXcQWhqUghf15QuDBjMBZW5rLE1ixUz8
h8j8GKjYD1BL95UkIjmaQZ+XnpucPwhjBX7FO9aQOtjG/d2rTLqzt2OrCPLN8E1+hCCorcZ1QWXP
YM8iT/iboYUPLl49tt7mTRB6JeC7t3Ceu4224m+KQKVw5IrApPLbZVjzBbfnIPF1+Cr7GOLNIQIt
wSHwdtlb6OtKwQgfZLScHUoJ4+R359oD47AHN6moZKojPucRGbLmlTLE4IK6UsphpkSogkjWUHEh
VndaEsZozdIme0+ItJkQVQYKX3fVlo4MWaUtrLbtAdAk5zxam2r3EL73F0w8cqVjkfM0q5UavjLL
rWlMUI5mJQBaLks0K8T+vcgp9vQxecYCNA7fV7thqiA2KCTxRn9fcyssks8/ciZqtHSairyQlvli
keWuDoaTuIFAgw3dxt2BmD44xsUS7TQrCAieKvZVaL0jPiJRElMOxT4P1CYKnQcZ4TjVX1bjRSRo
lIzTkxH24Vd35+pjjR6X7rJdoPrun4/MrG/tLXhfb2Z4v4V+8n8d67rtVULcjm0GOfCXuicc53D3
G04eYRVS72gvut6JwIW3f3Bvb3JMENfSoAj2g4zjrp4hMJvmzayOspXyue+s8b1aT5E81b3lH72h
QzaJmACh+Nkw+plGkgLyAU9lfi19BDpTN6pNqcx/u8p4/72ZGOI274tAX3/Jq4fvOWNQsxNMI4Oi
UYszfpknKBYK5OsPt7L+UPx/8Ht0IHXooyd4ciNpT35gyw72/Ez1DePNTrg5PrZUW9nPsx3U4FVt
gUxuocjD1O/l+8I29zmZ2Zwo61UqT/AW7VWVWoB4T36JXm7UNIdK/TM8DGNQCv9VgNrj0jLN8Q3c
RBM7ZTdPVC9drTk408lLE6BYR9SPbLnohkt2inNGxmiCIrxyhvggrx39AgmAmpBwaj0PEu+twp6j
88Xq7Kuf75yqJOW3v6Ufg3zl7iffGPkGoFYr9uTY8oYAUX1etN1bGkcVSJycel5BS7tioZ8oTVXe
zjKAjn6kNYIMsniBWF1kSeW1fFHSMVQrae3iE7i0cVrvChn3sfdvEceq+sX1ri0unsok5zlnN4Gh
8+uN7DrG1Rw9v+q/HonnjFSHeq52ATN1SPdDqcU4BUOZDObpIfLE9Okz/HSIKiAmaHw0YfZd+7DJ
BHJk5/Em7/ynfBjDV/8iz3g9EyM2T+ywWEyLFL7VMaEbmOLZF6WWH1H24XlVgoATpQ7MHHzBrYHc
ZD40GgGxyfic7biiSvMZbAtBkIl+K+eHeL9kVjDRmvnQGkFMBIVEQQZrlkNf1E5HmiAWXSTdw/MG
axa9WFpw4u+CRQK3c1sg30i4REgqUmAPfiP4RzmzxOZMQiea/EjnpKY4bYqcxt4aenL37mJK2DQQ
akb6BXGjmUCgiKAR/516mVV/zrR80mK3i37fN/BBgfEObw0JP+E465ex+Ojd+4ymcI/brGNoJ71d
M7Wctp21JP2zyVVXIWglpUyvm59YVAoMOS/AEvF8R6JUtnyovWE9UzSM4aoflQ/Vco6uOph40QYF
g0zGETdWG/p6laa5kqB5EIOvUBxfrMc1e6YISnqjdk7o/X2vvmtmzPpTe082Xg6N5/su6aug/rnn
tqKUk0KpQIIjGdqe8AuLKzw3gxp8tTjSNggYmSubLlrA5iGlKINHA7ZHMtezbDo12+QvlRI9uEST
cA+yOrlAvBbUD8Ewjpy0Uhp/eSQvI+8YarOfn2U+qeI7QOdhLpO9u/KQ2W64+ke6VVUT4coU9yAR
7SEq2dimfLzHmoELQF7OtseNgY8dYDpifUg84hRtl3k8rDg5Rgu+q2dQ1f9nV/PgpYmKrVZqFlcF
1yJboUQXwsYtM1mkr+5zXQGSp8yv+WHRgxKx4MVezaOLQf+foPViXpPWbFZKL7fyoxMYeEqldt7E
AwL7foXRn8tqCoFtsdQnXwji1vavKGp98NQLp3KSVD+QDz0a2Ym7Tk7RQjSV9hg3K8OkIjTQOCM2
ZqQ7YXxEWTJxmUyl9KvfhKMwNxk/5rgpWSvdrxBzdzO/W67tiDZdQJrdqCl/BFnJoyJ39EjFoKsv
4Q3tW5L6fr0psUIKeDdaqLDrxkycRdQ2Ld7xLj3HP1PplQrHOzLbVAiIeoD+XH90IWYl5C8Ab64x
IjRjK4+BOfSXsO6czP57ZOEJIozNjlK0Vp2N+2eJEDbYoQO3wO/BYKw3AAv8h9D85vhssg6/3SP2
1MAwzqOOXmFdkJ+Q4e31x6acN2MYyDLwymgBLcMQGAn3G2nHPXTRF6Ib/ZdlJmwroVkzrvQyXcOD
BsMJ7mVYFxlIWJLsVs5VzWwkswC+vDKmpZ9ZGu3Wjx9a+xc/5ROs8Vm+fN80+PxOspxj4h12FN0F
ppEBKNWjkIf1MwZx5+cBTUQl/eSvzsa2jV8koiBLtHhcmJ1VY9qqtflTWugS6Iba+qeDHezrTmg4
NRc116z9KjX/4JgUoewXtXDWJ/6Jon4nWONYiBMtjfV/0C1eGwPPxWISgb0MB75DGYtkCQuHV+sp
sKBCZ+Qwdpp9K6mPUrFke5ZLuhgm9eNWSXyimzeJF/6dbSaXrhg8kRcn933KM3Tw2xX1DrT64Be8
Fnp5Z/M8SP5IRLP5/IXcINaiTg9jvhLhrGG1eiL2s0n2LmYENjHNfj6l3I166JEh5mngwq6O/mEO
XrlDoJRaYFzLi1cHo5/9EM3goQoZpfUzLDuiWSpV4LmJSClL5Md+flnXWyqx/SanFnvRC4arLw15
xOqpRmploGPRum/AOuXSV4fSujLFst7HPvzeYo8wdsfWdW+MLFt/pyMuY7d1z/u7XicnX3hOdPzq
NvBG4I/+1UgVR/9hfb/IOn4yie+aSgzCxjot8RLLFnMrzR7Xf0oQH1vfN42J5trkv24i1FSllPxQ
olOlrC7UvNjZcJTuX2Efap+6gqC/FSrKmGENYiGEuLVUPukb+gxjtQDZoN8ThM0NvILIpU1GuwP8
akH0LdGhHS8jKf7zA3MqeHginLQSP/ZNj1Pqo5uflGuT0Eq9b6EKloC4/vYnuRZFq6oXuUD5ckwG
H15gt7QsjKccrJ2+0jYlRVa37y+eQR85zUMsT+2orjm9eW64ftoFlEkBkzG09S90LYVuPjKZcXa5
j2cCunuAFdLWb6Lm+bvI3O3Z/AuwnDgDWV2Ky/95CE4zomPBrWe7k0ZdCCeS7MuD2UyTLNY63N8U
GGZQ7gSFnF4xXOpMDt7TExT99i48S9AtQY6OHiwwfOTF56MoQ8xSFEj7gusHv94QFi5BQYQPuVuo
xdlH35EH1wvRdWhHUdO4TGTanCwBKDXJAO3SmngfuaH6l6grpNnsYoPkUb8Fjl2pGnK2wr1CBHqt
qCu1zB/FbSb+kUS8MiVfITyqHavKwr/Xwq1Gtz633U/wJiQzqXB4h7qM1hKgCevvDbt7zNbPubAB
QnSYL8YT1m+Bsyt+a0AbvFki18OLai70PV54JMoj63MtMc/AAskod2cZ1ljiQ7XErLX3ZnyjcGdY
heoTcsEjQYfSFsh7X3hNlu/I08Xt1f8CnIqZycx3ol4C81mfZBYeEJwHpP9Nm/MXCiYeMOEZZSz4
iTB6h2qOkqyRuTmHV5KT5rqtLvHFHCF5DPD+xML6pd0TLR4y3O0tgu1jimFsaaAqMdtw2JlAb8IC
MluGkPAy6q5Hdf3DJtv62p+1aXs8cvfyWjiosnhia3PQSKChWFRyb68aB86bVUTxJUl2Ks9iP1LY
3r9WAawxsYrPaA80cd0ulSmKmh+2240Sq9DeFUwBTPan3D4rSC5rkudWbM8+Q9xzAsiXeYRn+hlm
rzoWmdnYrLShkeIPZ91i0EYV258MUkYN9JTVz0ZAtiiT6Bf5di3Bsb519i+QDfQiIn5YkRdFlGlD
5cQ/MPQvfenA8VKyidZQ2R2OC64Wia0yHX6gD6v+KaCSYC1qJEVt66VibevuDx5QjqVaFSkb5/sa
dqoVMjj+6OBXroHyn39S8qnGF9J0XL1/3y8sCYEbwl4ueRpzVzReMHRotCZS5HPpzF9IU3u9D6Qw
nvG9kfJ1C4lBRKOR2RmLKN325Rk0sW6O1pf/L37+FoeQhM1OHEkR4qT1NV1CrPDtuc/880TVjLG8
2TFTqk/7HODZh0yKeJ9bFrN+Se7VF9QJYBnABdYSQIW+kSoMIREChUn4n+54XiHAUIzI3uJRI4Oh
LsJDDz8Jei4wj20/Pn/UV831Xmclu5Fp90ebZVy8r/3kMqIvhkZUw1e3J7DOmfkQDt8t5VcdpFiX
yXkw2RRX5sjji9CQ9ZqKY6FHlL4y/uk5zV2hdrS+Z3Eo1hSwhB7tHrbpSUPDmIsVtbZNsn3Tw9Gl
wC/LWMswQqA9ybnKUcnOiz8c9K3nfoJ8NMK70nuMRVYfSu1JO4Ksp11Vz44E/maUy2Fe/wQGPvQ5
Dsha8J8YaQQB9zzTvZyQzdD6B6D4iKnaa+oXFWnP+JV1rHQUlo7V8G7xf9EkeRK7L+sRJQijNCfS
JpKojJsGwc7fQnqyvcpaaBxP6m6kX0TPJ5kax6knbnFy3wM1mHFQVItYLVHf8Y5KA/vgqoIiRQ3J
t4NKi0A69SnZUlbm+lhv+Ko6SXYPBPfueZtlSHLfiYVwhx5T6UaozzT1aI8G2c9+xFfB7opc5zhi
3LAXSNZ3wsqfsEC/Mmpz+JbitUbTqUSPYT3WI+mNOhTh6/RSXzc1Mk39CXtAMTgQSpQ2yLb9Oy8K
BGC+PDVeSCg5T7A0+z6728XPE4axs/VCgRQt7fRAaaCTUNWQd+t5Ho0NNwtMRnWIVkCm2BfUNdzR
WBxGE+IFzGsAhMm9jQ302h+CTVw+yIulP1/+HViLhnszOxxoG+f+TAFFlVE4ZzwvXfSk69ZR1B42
kclvzKNwoGYFRj6qcSQcnrXvzbyj1nqmRtcb0LStrZxV3jhpE8WWpxSb+LUJ6SOQJPaIizsrU7eQ
tU+9xjYgkmfS1uLzr9ItXo1WEgJbiCfiIgRN0idrTGoL/MEYG0kmGdS0Ut4SwS+amUopELlqQEn5
BDuB4DJC5PgFw0YPBFhM4iRnJwgy+izeur+nkjKBc0agf/LMrjIREvXsfUFl5r47oDFldWbdFMHS
EOVpXjlg1f9GJwZQ5CSzGy/Cu01VdKZuW0nNURVzyDk5wsaqETV4xIK7Qwo1grz6iLAXtih9WGtr
qKdHyB9ULM6PE3BlkPWPuwdSIPi1W9acKkyMvaKvGIFh8qiTVGfx+2TURCb7+BK+oo8N842112uS
ZORQdaHNSdaJsRfCDb8HxmPkl+Ovl8+izLjVQlrtvKhz8jYxWbyJRr8Xbxny+VOqx5wTd0fcENTJ
Kmjp1F6/jeTC/6lwEaMzjmdgqvqSQkWriqlMVDdtT6NGho8SbTJGzoqYsj6+Dri+JqVw/EDg4Xyg
ui2eNpA1bbZJ9u5di77Deky2ifpVp+DJv6tafVkwXFPM54p6vof6IU0XCjHoK/myWobmy+J0kpHy
crGlVrd9v/wcI/6bM1QclHXpycPTdqYHG38711qc8tzE2xrc33bm1X8RpQH+xnup4jZmxs83MtY8
27fGRSJzrc4nOOIE1MVgGjHOw6Pq1XYJ/PToQXfPHxSMPSOLvHqB83xTZur8Y+DoknZevc7kX98+
5gS/tvWrnL3OmBP37NTUVvZC3e1Dxki4gHtYBVvHtou81tAXIK+Yt8Mg9HHPtkHLQ7NqEFp2uRqH
ryDRLYSVpVoCEMhJg32S3EdCUZyPNBwxrsY86XBW+8carzhzGFiZTvv+tpMnkWuK8ViD11NIk8zL
J2JEOYLQEfMrdt8KnUkP4oxGVxrdmrk7MxE10M1h3fcGu49NniyDws6BQEbLUBAP4cPhTvh7RRbv
lM/N+64iV0PjytSUu4mC9t5+/QN/Q+wNACS9EXgNdDdAu6vrwkC0QpFHu/ULSMMNQxhrGfhx7t8c
eexxoB3JLL3nDh5LfZLJMSG/ke4nhh2JXlf3xDhRvk6EIrZd0pUSUjcMF5yzxW6euF5yF3Dj8VUl
2iWRYW9wbKWLpUyki3jt4/7gy0uSjK48wpthwHFN3YT8L0K2KVvBcMgLQIjoGGMWwmY7ud6SfsYq
wx8+fzihuQqQvk2sGk9A1sVDXRjQk9Stt1f6MFNdH8HWg+bD0+ZZvAahV4PhP0Jwt8hVWBzsdQoS
1mWM9ZEkQ79ljYPpBIsdCUGABKCuJUm0Szv0fZtH9cZ+6SAVujGhIjOdRUj+iBI2vfvx1pTI4kB1
+usif0keuGGILQYy7zZeivIp9s7WaHDY/VhgD+UexHNyfWOSy9uEtgGY0ChN3uNI0Ccj05zCP3gf
9mHvID+K1eyNDrOyiDa4QJQ9aQ4/L9fw+v6dOtCZA3t3eYZjoRJUutzE+OgDbwCZhovXGa5aXhef
w/8G0kCnffHTrJkugtNYLLg5PHjUajAsCIyiGh4FRAneKJXmY9Pf0521O8eCV2OTbyjFa6WZ/gDK
o3sKoIKerVL42RM+b8bJD9VX1dzgEek5iDAapRyh5OAL5cT8dkaPYe+fBPtGHccfNE5lmffr6fwE
CUSYaS5DiGCh1KyF6Px5cWrv3x7JWJvfyGKSP7JFPD7V3m3ZqjkYglqXAh+GJwSPFqG71XsNqqMo
buU+a8S0v3V//m8oalHJosL0bHle2djak5aSYDeGQZTePIwVVmxltDA79lD2Eyh+kcbrFbxe1fmf
oSfQaIb98TWmVrD/bdTRuhXKoai1xKNH9EVcvR5I6/qPD06vfBLwZF9YtCXfIdOGqstMQn3/mNBq
Np8Z2H6RJW2AscJUDdgH8dLb5dNp1C7GWt8qaSsQomzqe+e8h58Xd4vgmBBLeX5jc7mkp+2BQ80p
79dv9Yox81I6IADT3dZtERLKVoMgnL+2nS0ZUOXsHAkpc8sQ8w1kAHGyiYtqK/9RkBjCpkNtcEz0
fqrY6jvFqSc+GplhMUpBPgR29nZAtTDatBznFxG1F+U8phy6bCQjsIPdNS3btS1csAd8X3NiGRV2
UIvD/87GWgqYetxjJwG7N8y9kF+AuXQs+7/2rLftmpQd4nJCh05idGd8AZnmT2cJzUyqO8YCzoS/
5kqt9N9PQK6LtSSHTlbgXC8RkyQ2jjC2uGZaYveVrDuECUw8klqn2tPUC8fY5RPrgbi8iaHYdzpf
udMyqq13q+dURIJe4KE6HHySgbDJswvyXGdah+2p6bX/pZi0ZngVzMc5KipipQYnyhN9BAMzOT2j
GgrWB6Rptyn2ttXwpc+8JaeI0cFJnXa9346nPjKMm5n9TZjidyHymF7+6eDi1jEYNZ16Q5EnecEd
CpEmLGxIS68CTp6Lu7WPSZFi4uQU9bRvOx0mpnSzoPjuQPMWaFrl37fMC4FMYS0NADNiJ7luvIui
IFiad1GtHoAuqngqHiZ0fAGQ30R9x46H8W6dFCglNT8aYwEhUfHtFFUhv43+f4ghSDn9zC6CzOC7
Gm/R+Nv4FGZ2q7KCUaHtGsGG2Q8s8t3gV/VJ5QxjU+jmVLzKwbp3ObXN4DL+u5mrvKl7MY9rJ+nc
Pfm0edfRnmFaUBvCWQFZa9Oau5SbnK8AMon12ex97oz38ew2/NsFrFXTJikgD7itodnERFow22KO
t38wvNBf+yySuW6S7+Zf512oJx1tqRiVzh4SxmU4DTzp90HKEtc/KGF3Kcsr2WdEjfc4tsEaLIla
deV5hDo3wzOrIIIxMkJ5LPmpJJvbV/GIYkFrmvGv69mcGm6wQAk+QgqnW//VZXD8UNuDgjYun5RD
DA2VIi48wsrjeBvoia3adPqJuEMio/Ixz/Lf351pUkiXNzApU3h+hXrC6No8FrxKd1zpLa1ElGPD
rf6K6BpVsSDPDpUJpRhANt2L6/UhfTP2bqBKNBbq6BUF4lEEeGiSB9MMxK2m5x3yvuVitLM5JUCU
b/pDrEqffffrxNWXwP6rz76qjLvtDRYFijqy8KT77pdq59dGGkKhmdeYKdz+oUvnSA0ldVRiMFu1
0es3ufeVGqmoiFkO/utSskEvNkoTYlH165scYQIY5H0LGHtNjV8TEOgeefcivnN7EOLubgcIs3Gt
KuM5hqxcyhgHs6SRb28DuwYXGftYlyqizxfCWYgeww71LMC2s7EOYFTBf7CAXXgVSOX7rgQVdL0j
P0E23uQlMSo8G9zK0WwNwMocgnp/Iep1tCKS/vL5mYm3DML3e12pI9zxFo5loEaMAlDgnXKEu4p0
L5SyDTVL5Sm8s10wEd5JnumSWaS2qwI8rCo4I3qfp8OM7OrVd4kSRL3PwNn550ZR0HhhTvQuK+mv
Kh5kLtZSoCDIbRsVDg+PlreRThghTd8hRco2+K6LscJdT8pMHWVU4xNV9cmybnEDUbKtGXqAMfn3
UF1oNU0rxMCzFJ+/YB07kPfK7/hi1DSXKxx8oDmFkBmI9xvFKggL5WPXsm/+JzELt3V91uezGokO
1aPFvScfkVcoNhUJoZwLE2LHOEqT09JqztjyjGTyz5imfKR/7W+0MbA41j0Naju9PaU19VZShTiw
Hc0JP8gUvySu19QA804ZKVrYb+JvaIInbqSR3mlGCkWtuVVVV9Q98E5RaMscSttBu+W5Dkz1D5PT
/oCzvmjwXwsF/xwsfuKxlsCL7iQZ6/A57FDLgyfq8OvLra6Y/l5g0VOA8p86xyrRZpF4/n14m8ef
3DQLhuYr8ODR7+Y5TS5/SN1eJxM6BVfNfxzPUGHz6rhM6dXpHhr+a+FGzuMlSXB+/7O1CmB8hOfQ
HKDmrDN09mt0zEdiPcGnfVJUxC7AsPnt9MRwhdMS4Yp/MQ3pbRFJKDxu77pK/73nRrJXC2RiOBvD
HnXNDjFUPWLLEMwFhGqT+ifrCRQzWVeIgrGEtmFCnS6bFHUU+TMJP/MI6omuUzzLHoVoNGchT8Wa
4JGlT2L1MjtDj8aNaVR0F7JH7OMYxMWExolRs/4MmqKNhwCQLJpCion30JEczvFB6d0ga2STw//A
4RECpZjvAy+JUgSsBS8KjjvsotRR0xC194NOchX4dunYRjQ3n45FDGTCETjgxuKJ57kbetr/Xmcg
xpF5Lo/zWlDwIyJabreR9+42bnLV7Uk6FL3vww97TCfT8eBF+Y9ic3uqpSCd22dDDvm5gNEv+vHM
Cs8ersMayjURdd+454yi2a1dEiS52DpzoaPBqOQ8MPS/J2WiwkEbpcpvHAqK5vs8SD71BA18MLTi
b6aW64nXImCUeI8OsRWxKEFMzixmmYthWJuqa7+PGLI1hYhzHOqnG/Dh79lUMmbKsmLRtXtwfxvo
RfTUrCIXWKB1fZlLCM3zqL8xAFdRtaSRTME5Ix1AFsK1hl0EM9VDQyGFYD5B5jFxKfWK7boQn7NU
+jif1F70Zlw+Kc7r6bmK/RNO1mezGeeU0MykVI2Cw84S/WSMBcg6I2hyMUSOFgePZ6OPJmIsKRwO
u33LSOQBaa2rtvHH5y1pIQgyZrjNUNhJ6SohrI9vcrpACK8ZAojsY+pT6ORjrCo80f2yt/hotM31
91BTcHf0Sjmihezf4pne3J1p3IO+L0o8lB0+QX7eoBXj5lUHJPmj2KWFBGZ/yNCum0FWpSW4bf5v
o1iKKiGii4LkIID8pmP0LQUB8gGboqaUD1MXpfVA2h7KIgwFtf5pd0/7OGJtEb+1W/lJrxqstFdZ
5MgKlQ71MYybF1M7Y51pKKYfpvKdM9yqIOapRFkKX9kgI96bl5dfHuJPgXIcwpfaQcOhhXDKuyZk
ddn8QBlKARrw+URZgLzE903Lv3zNw7bhzhskVWtlGWP5VSiRc88JLCp1uUk8LvayX65XnxWNG+/n
0TWNubwbUeil1g8JIZk0V3uNtRljIKd6K5qlb+yd+YNYZtR0H+NX8818GwsLbZZ4Q4v37a0DOMJH
edy667Lunr+jjGyIzkwiPN41bNZScXsPm65GITyAGEfrVh6A4lTu2UNlEhAMdzj/1MQ6ldd/dD/Z
Q9NrFuhrN+A0siBfqpUhh29Z5ygeEMZFVIUlPDbf7s6/9h97DjnxkVafxzR0v0g0cegHEErfVSfa
/rQafQr7BSE9O0PLvYloIRgFj4TRmw9fIhvRfxvuQSYHpfxi9Kq8yD9RSslG5nvYLQXzC1++wzx1
sK7KlAoWO/F7GUvzobYp3wP4DqKSeDY7RKBIq2tuJ4xV3k+F1RIJDPSO5D0wlBsbttyTQqHFx2te
o7so5zyDaQWMoRmjrzV8MO/8YDj46Qh0I4mJOmoTQ5N3fX77EFUo7PSrlCvZhlfUfO0+I+VJKEU3
FiaCLls4EXowXvDoNmAx0y62v2cWtxXuacDvGbbY5PD7M0+3WNLhJ02EPueFMxN2Cfk6HjpmHxoU
IDltlgrHxanuJf/yjJSVtQHjc+gy5gXZDKNLLUBOfS1+6bK5Kdlaq0POgE3e+pG8kHDE4gdryef0
RO4GtCg6AGzbJb+7eUoBWZthQlPyQSVTNnZhDYynUK8ykhAxk0oJ9/F0h3WVoUs2I0ZRFHTk9aGd
W4fQK+NBIScebDOIKAjTAwor4u8YjK9UuLbqzO9CyccJh2oP8Dr7XfU4Qk/K3s8+lgLDP6oEqsfC
alsWSIAEmDOewKlY7bcBMnsySILpjPXw/j725XUagxmmrUoTxCVxdnCrkyIhAbV3dnj9zekFk6hs
gi/vkZg9+2vbAnuzinGfrRP7RJylhFeYSo1Xwku384REAbXNyo+WmxG8uoJUt9NmfFTO1urVQA3m
c0BHWEVMwLW0rQO8y+pqR61wnfw9wmHPND0aGb/aDZ8LiJ0b7vs/FEAaMxP41QubleV4OXz9kNNJ
JkpDVN48IiNuzo2oajTk+caGRLnfV4pNEk7fXSfkhFN3wLY947ohfguk0eqYTKRK2Q2NVmJloJEC
5uEgHd/nTGmWH6ZvFM10hdWCCgzh+XtCwN7Yuw9NwX1K2V75OnBrl1Hw4f0H8ZASYlm3Nutyvk8G
5U4uvnRLkOo6IBNuNIkHsdD3t0sQF4piNZxHv1oiBSVjBsIAS9FjC02BlBeJ6e/3eDvuFVqHvnTi
bRwPfM+blHqEdLIPtffIPiXEbETEyIMH/3qwIwyh3W22zez80KD0lhFGLULL3tZF2VihhMJ2sz6w
shufJcAY1z2+5qIWoBhSjaTwpGCz3t3mFs2r/7TixV5euiDiUtdz+hrWRZHjrrnPyXOawAEp+uP5
Ra7VfTkWR/MnQbz4hPDEECtAlkIIZ910c0R1MHXDzXkhRwFGbMja40YJnkriLCpPD5huQdc/ymDk
p2b/lt1VNV8gYVfBWd5oz/JKVC8aDHyhtw9TNRq3WK4OzCLKHMLykWW4H5eo0GKqHvbIIrmGEpk/
2iX2SGrrVTUKcDqsTBm/sSwChqz5isKkVQFf/jQuaaKtBrv0782BRoTXiJouiQhcj/ufPGQVS1Oc
Zl0MNMwMuM5YRX3/M+uuXvdTqsm64j05pZO24ndOwMEmGX4iA5pUcVSaNwKhel+u5zlJVWv11+po
Goc02NAi19HuFGFxZxjcn2JItRHtwsv34umDkPKKXz51MfBX0aRFS4znQtKdqh91PUkgNBsJkRSf
bRDLm1m7F8vWUCS33SiC1KYJbzubbwdoM6lK0r+u7raLg7omx5/W16e5TRw3cbY4+WX+UjgYkEoQ
1kpoetHXcgc6iMvPlfv20LUN3xY5juQNtU8owVYmLNsXOWlgzkbCJdiPEr830IYXtJinZoWmZZLF
3gRFVOrRYq37HlnjiPC7/TpHFew7LeRSPMibe0rVHul41vN9q+33/wkm4u1sPksqYTzlPa7ELazB
JKWkHtxwpipZUVAfCEc722psEKfuzi1ilC48Echk4JmpCqxTsRWscKaQ+V23V9bQSqEZ4Oid+e8f
ldDYESEVf8onsDqQRWYlqA7EMqRfy8NMe5SwXhBxuxi+UC0rc/a6tOSEDbFPArB/6YiesSU2mk9S
3ruHY+GBYFyi2LAiZEbybjupKfWc57eXEpmfz5Otq/fOjd/OJFTgmOGuiO0a6lEAdV+7wiyMdozw
dhPtA8WLQQPs5BIrzL1mJctqsmVqEEflWjmqQkWo3x8K/L7EGCgFPi1Sp1/9gCdsasaLilrL9mc2
o4UuIkGTxS5V4fclfaE8EhKDuj3IanmTCM3yE2WCv6lVga9r0C1SCpKTeqHmjpvb8JLXl7DjyUfK
T9+opZhsIUA1/5uIaflSnkdKqhsrrliAJeJHrP0prIxoJzt+AP6rgW+XmwBoXK+9I7N9sPuH18fZ
jwlIMoFjH+H8eMAfXV040tjP7h77dGTVJAwTn0a2/smVMbR3MMJAqHjidzB8NPT/T7efEH7OGXUQ
nGUkhqkwkqpK7xmlOjttMn9wZ7fofG+qoHNArLjB0D59cWXlGgMYI8qg7VdK7G7u8lYCeg8Z7JQf
Eb936CZOnHWbZwsEuvUpNdElsi/mKUVfngYMcsNf4qRVvStd9J3mRrYisY8B+YWOyXCmbocW5uyO
/Ea/Wg65IiPWjI7X+jINT4HMja7lPMXou7eDpqiQTxaZCN5yazaA+8PjIvIhblCEh+a8VYcKj8TX
MJ2lxHjzOyJgjKaEk4W53Oj38i5hXaidwZexeRFotTblaP2DthSp/B6soLREXG3KmGFRmTMY+FLa
f7pcAygdu3kFRY1EuvLLaK4tS6gWqfqYm6NJx4MRx2L86ZsL/XLn3lUSZnHzkpiMbQ1BcwtFPn6v
IiEkyewEq69qIEBjsh7z+yLfFvACvCP3Z7h/9iu7kiGq6YC6m91bBmYyzNHnkbM5/F+73s9hUQDg
Ebq1mx7QiMAORZWp+0zMSodylfwfyylGIrltg5anSFssy5MIcT+FArdrEUj2CORmjHX1ZND5qSvk
qgFgfEUoQMAmJ4jEfbXEHcYIcg7eC/qhJzIs+7l4V0vIvZn2TDFAI1WLXL3/eCKTEtCyXAPyaawc
ee+Z9wLUrcJfLa3ZY0cqurv/1jalFDZCQIbZPWJXbs9N9g9zkRUwQgYVRDO6uFA1oY9PTIgTXIUE
sVsrCiIp166S054hiSCew17pzFPCu+OhK7EXmd0uuBTxwW5xLqjIMHjSb0iT8gEq1MQmzUVuXf2d
UHLQJo/vNdyVrmeUTKQUeteCnS1Hn8R3IiabaYHmTgVezwf2jd9TvbVfXUKjlgjeCveUZwbszaUq
cj1sSaCVwllLNmtArCkTygKcDyaUVoYu1Hy+sIniX3dP0+zSvML9PuDdk2p5Jk+1vR9o3RwdFSmZ
dpwMnUjdvUHi2lA83djroI9CLarVJH77OZSWT1MznE3kHeNO+Bv3SSJ9NwIJKluGOghibuU2PLui
e0nspclzDAfMlOKpQkZi1kPe4d7KOYUjEAh3Xfaf5k4h93cldquZD32bg5GpDPNCieHys+pzdcbY
1msJuzAVhJo+VRQcJJoBxzoM8kvEZiwjtRb+QrOKZXWLsJFiuvWGh66/jlgJbo/EiPp9BorgOTmp
JOVtXOckD0FtADpa6HqColx8jjsNc/F8Rj/V3Oq0gjYVT5bctQb3gXM4IbTqy0VdXO+DkQzk07qL
VsxjRmvhnFcy+l/baWfbfQYO4S8NtfUKM2FjGI/MrVVy8C/1iWiGKeSDiKgCXymyjLlBmgt0PmKT
H0DyJKxezeBC/PCffEJVBBh0/Q9IfMcJngszpdxtRJB2desch+SdugvnazoCprXav0bmCe6ntRTn
j/s3esXBMLLelQjSweNKK6S8/tNtqvwiQGlvKi6mmLJeCI0/nQyIg3VpTrM9sU+rHfZ02rYn+AK8
3OVc6WWfD66d9MgiKDZIXNQHEI7DCdZTNz1/5BQM68ccL4egaqw3OIe2cIgBCv73HEktMQgmntSP
YUNc6jubwdaWfSyaq4yT3MuUauQ53/kZY1Xl8ZT8g5kqqtVeT5hj7/jPFbbQBKGwtQVThC0PWqiS
WCvL+hIfb5kUT6l5WNIxXbP1nSykUlkCqXFIn1bzPh6FOBLtn9pPhpAxueqWoe7g1xzAi2MB1pvw
soCBPjr+C0l3RQc5cn+TXSTnPig57JaEJYn1LJQ9CH87RUca9XBO3kMPgycvHQdShHQvUYBuGXyM
8c3BKNFX8T/vhF8L5g+ScJUUxf58Z+pR5xr5bFudm9Bm9rBWzjalpmgcfRKpmHjv7oOIPWyoXhuM
S5tJn4ovlvkIudSOfykV10KC8Ig54YtEoYWn4jUrktRxKkM5PTx67hBqT+QHgrZ26cGRAT+lhN+K
pZWJxmVEQQJY2v/SGQUIKsjfZwCKZxCpdRuuu4X8jYY091CDQlfENpHtoywzLZQ3icQYNFnzwofS
xkkJlOkoARwLQ96EB2wmiaQUOGJmzrb2jy+FoCQcp1vquVe/xstE8VtI+78drlQV1w2XlplIh/2g
AirWLE92EX8NsYqdLWhEvSMqFB74DtjAb+C39MsWr3/BpIt/xhhC3YcnOoys1QBJFi2YN6XIMXQ0
uB2HgfmDXxoztqr3nwR8KvVAS6yFNyIMc54ri1YT4niYcXY3d0MitfKyuy1Rvkwel4/0vRjb6WBz
ntYDaItiYNSWz3O2CtbAdpVBP5OERvfOagayGKQ8vAA9TAH2WSLmGmH57G+2tIG3DLpN2Qas1tgZ
Q4phP5pKhQhWPLsFbZC0TEV90jm7UrFDUumpf3KrZQpvDyuASy/+0iqPpOXC+jE0ZGRGoxSud6i1
/0fgRb/5RYdzN2xErVBWkLQscnECRGf7U0moTuDVCv3aeEyUgFGhgOXQ80lwZNiL4KPG6VKPjyUp
OLrZaKHs/+4if82LQ8w/VFRYsiXrtUn100XwGjsvtKMPvDPGcU2JNFkY1VC+a9iTFRks6zKsmyCx
MGvq9yXZBcIFqT+q+XDk+/smjeaPeKPOc/vj7oMRHQ0/8ZQ44NhH1+5EVwbyetvW0iPYLYrL+Xzg
UXrtqvNSYyZwVuG2NVx+TffJW9bN8WX9gUl2zABON4wQc1FZhJkM0g56TOlJ8DVtHrUQsRMWsJl8
p9fXIU1ujnMJRCjpBhEhlVWhF/8b3v4rShS5q5pU2N6hTtycwbZr9Z19QH/oGhPbBj5uhJtW5AjX
jAdAmq0uPCrptB6qi1NeHmeoCKKBngNL0dUA+Dk2awr4ufTvYazje+KlFbZRNUsocRx3PUhmSZjc
25xPs8mXRRdGFIEDbmR18InV4rwXI8QDkoXEd2bJUfXBgQJJpWfewZtZ0R4z+QrvB+VjdJ7tiEon
e5SoZivw2pSvKHkZV8hFeLF7k7XZ9u9n4va+sIFPaavOZE2jXyzj9rU2lEWtU5c2T7/SWc0858BM
P3Osi2PxWPFy271vd6Ln+V1FMRBCrvzAqdQhUgDfF21FUNdvYyRs5Bqm6bxqwIkBVatBh9bjFmMq
gvZheQVfUHFRm4Orv+MHHgvBsha4IJA4RLgclQQ5LppYzzyt3DDhIpwBJ2601iHXvKryN8DOf6pf
Hl5b8e4KgeWKEDnpX4efD57ry7mNKQ+A5WsrkMI+U0196ZQBsPFFI0NuLwb/Ix04Ral1A2cOm0Tq
9bcthCY9tkTpWC2Y9Eqh8Yz2dQIt0RvHaUX2nYitVtaPl06/6mONphE/gmhQZeokNSgt9+BlG/7L
Q/OSV+Bx9bf1lsS+FEjPcRVJCA6JDxbk6Oz06M9rPrdCPmTNGWuuVnBXGMDkYzoyeCsfpBSLWcfw
uAjlvg3+ZgmPG4RsVNqG+Bs2FTcfIJph+LDwKuPttRx1RuWUICoXWtT7l21bmu3qqInk8A5ix06Y
FPKj/If9CwRvNe92HIHVbhFM2jTQe3utCKXZhZsqC9xcY0lx9NgYBX8GZriWeYBBZkVmQdjA7I7o
JOFpvimkbSpDCnqwDa7N4c+FD45jOCMuKsGI1Lx38ZsOkbndZpwv185Zf2wtWXGbezhDBFoj16Yt
VtWs3R2DErgySfgUTpRUrU7sUsbDYe7Am/rL7h4FFcwFDRXkFm+szy1Fv09oOv+K+euQARYVo9LK
++LotlnbMcjHIzWNWtW1E3yJczVv8dGczE/PrkBdsDwoyFP/pJR4T1Gl7CspuE+m2ObRozX1m/Dw
rqT+RwzAzT3/1IrWjRAI5wU7um9V4Qk3MVe16HIH55BH7jNzRNrWVsEnUjz+ZDfQoCTPH1fYeL5x
9NvQObzb261Z+lY5EbvVXko0cJ44qOGAinwyk/pf/eDKvM8d00Cntuza1vzRtY/g2De8j+h2yPKX
ZeYnq/Eknq27BqNwU1bR9wJp5aU0+sDSscqVcx2PUf/LR3xLI20RA7wxOCsf4qK/3yvMc+/p4uY7
OXpkhkanADHDMbGYOJqgbFe3/KDp1gSmQGfkVg3N2grVHMAuAaD5y2FlvvsT8XN7A52Iff+62/Dh
x3m3Rl0QtIKXAnyBgTt7I8w6KYDN9pp9os1rY/1PmnYTY/5dB2q7HorXOIKGGoBPtyaizYC1/ZHk
OGC4ogjHk9CsuphF3pKZ+NSKb+2FdZHklHMOLhH7EuUC2WnKELfzDbWzgewJlTlVn/P5DOP0ppXR
PMNCfrC3HR7LvQPdhor7/1BrMcrEIYXdPqMM/jAvLyDI+keog2WltDiLOcs2/Pvrhga/9HI+3nRG
RnVhN33MyHkxl5W/0/i81NLja/pIAmmM8lE/hTHcLIDg8eY/1GJEgYt/tyFIhmuok4P8iTc+qvPW
lluV8SYFnjVqQX+V1TjIwZRsmRun68Z2nc1nS++HNZDfJt08IYHCq1WtLJYYbET/NT1e2Mbo2Jyj
rB7YrKePAZ3oEM2CWJt26NmyKJpbM8IDPUK6NzI3lDleTtHzcD/VeENtEtcS4TuneudvG+hR/m8I
Mm4AsNYQC6rTyppAyqTIRlFYOSKNZ2BwwzXSlflgq2kcdrZroQ4xFkYVGThSk8UeZd5/h8HTsiaM
SLf6Fe0K0Zx80PtqWTRiFjaCzWNFkYKTjxJC5YC8u3qfZOMwJiNQg3sMAUOQlN5OELALlEecoM5b
3zs+T3q+4vlZ/BNGx2SP2CeIgR9Sk8hvMPNlNgKej+2KBQSJgUEae1FNGk5vuV2iIJGCBkgOQ8/A
RI7XpzMH9Z60sfj3R3D4fzPJpo+Dhlb2i8XLp5+iprBAr9lBdmUO48Icj8qVir4uwzY8Fdq1pmAL
TFRVhGtYIcY/Fh9Yk/CvZ0t7EqZgQxX4xY3sigV6KgCrtDpIbEnsTnhm2CvLbvQvn0KT3BA/47+H
yPiq0Vj0JFkmoMXClcKJAEpPr6R1/KkFULNPVhg9kmLSkJdpOPNt0uJebBTWOxQ0CxVUD3s3DF9L
TBbf9TwFvB9BI3LBV2PWaMSRVoKI2jKBFC9Zqf6aYSe6Z1teenJSOxj8TR7ajSog8mV0Sg7e2tXW
5GuWCYQwUKG35RNcCyrFS5K33RPbpM18nlV6Zr5SwEZXfju79Hqpin1pvMepKwPWQxwo9BDZpUTH
rUkYmvmLo664wxZItOA2ht66NFoeHUc6vm9Ymm9YrVwqMGN7h6sakzzYLIECbUUrOyA4n7ENFZWY
/NweA/SBnPXhe1/qZXhCtEDuAUz2/EDjD/u7rRADm3fsGg1+6hw8xPdCuy5OAQ1bmpIx6fk9bKOl
EAqYXb2hV61MugxAiQW1R+onRh7Nq6A4mpkE4w7mLd1J1kuW62R1v6sDPoVbFjAkjQGtbk4+RNY7
MCkDAxSM56KyrzcxYyCHOfJyayYn6zi2q/GAO2aReD1szlhx0SxX1/2CA8SdA4d11/8v66IMdF03
gelk874XHoxCweUPpqtJ8hglxX2531FSMsKQRYI3TTpNSVw0sYWB1Mg2L7dgt0NCWg1siJPEI2Mt
XiMGbNwnrEbus86tgQcKBCpgwutGLqWZubych1SXy9qNFCQe00zLDiAgnPLpxX6NQcBpZO492nFF
8GcVdD0Cd0Ali0P9jEdLsmO4bfLkF6bYNN2uIhkU35qmwmuBygausBCMgQUOeeUleHrsl2GALHBj
ujk+v3BaGwJysOMWRlUhseDn/RqQbDnBlUKyLc0SmYAQDdRCi44r2wfgWCJl3r6oQuTGbarx8qOG
eV8WoVzTw7dEfQFtUngDvQZkFENmMncdjZ26ceO278dbzsiC94Q6Y42yIh7Pvr1MNri/Wx8GZpzu
YzOXhsWy+u+tFLjwkriSwfB5ZKLm4/bk8Jxtucbuqe6KqqXsfEBNCmq3AI0c7luNFaQoEPArTPse
NrFlkIMEeoCjoWoKUyA0v/jErHOQdlh++XP3pA6ZIZ2BmetBWyUuX1ODWLCOf4WU/Ch1GNg3gDTB
5qWse3yPSukYPuauiY03aeT45S1yLBDzHiPjrRCx9X8C23mExp3AkKBVVUX/jo6l/Q8qZM6WQQUT
uue6///MImjNIF4FHARKdocn1+DXYNfsTBSnjdq9qeBM2sP3TGIUbHLgqljd6SorpMFxtJss0tol
JzN1xpPXPB4FzT7bMU2x2Le1KN0S2YsWZ4B5UBsbLspgF6gpaYnrsv9u4X04+iD4u30G0sNNZm2Z
pS1Y3SmoxKttECJSdYdOBWlkf5v3r+X0n0Z3QeGoZga3RQxJqtTdUlKq5o20ZvkVNLjl3s+ggPKE
yY50JMNaNwCd/x1hLdAnEnVe7Nd5pGAHKvhTjTPbBFRGx5U0PxGk/MXakmOpCacPpzNR6CChDZFU
W/gEhFe67+fAAV3tK/VogoUbC/uOWl4J0xPW9QGQTBmF/ASFmXJpGG3wTGx+vVITHGS3l4Otf6Lj
hwD5R8KUxiz/9ZrWm01tP9QERhwFJQG//St6IupykbJ/a0Sy0hTzcVIpJoFJaEojAm303r5nBukR
rn7sIv1/LPoX4OOy/i01rvcRnrnmnFvUBnli7nni1n9Clix9ln6bqyG+SJjsJ86UD5mHV0cjEc0h
bUlRh+5gF24FEhTUOA1PWBAIiKRBhlM6MTlnsAhoablYEr1VaD+J1PrfKw9CTVs5oWxdOU26f+fl
Ms/aY6F2LHFdQ450uX2Ri3BSJZIa6JYqwDi5rgjsPR8ZCzdNIMZtVYKOyO999CLiX0q+vuHhQC1X
yYdnUIcQNgbSLHqfnWrgXxQQ7TuOO+umldhUm09DaE9pewX5RdO3t7edJsxCoGuc/xzEqeRJ6hdg
mU6C+/ACvPK6eDjmn1Qoe6KUWPvWiV8uaMe8I6zI8bJLVqon9qBw8EBvT3gSErelPxVbc1cU108y
6CUoIB5VT64tzKYW/koRidsIfVBW8O4Elc52R6TD6d7V2+uEesEVBy1kNDLQVYb8ylH+EGP+h5Ja
DM5E6k0INc/LjsX1ED0ubOARPlsek411c9dc9+gjViy1qB5y3w7GiDlV+QJM9IncR6LwecUiDM4M
ROEZv4185bgTwB/g2jcYslc0Mg/rk4+WuhCqzZE7Kn5tsT285Yp+5nmkzcM47ffistMnoFtqKCm1
s47m91rE3l7NjsW/FkATljeEUYA3OdkoM4F4yw/+ywpsfCX1cXoUMLu+67eCxwUJUcWwL1Gfveuy
VXndYq0tMrF3fXA7NJek55ruA7moCVpVV+lK0b76zTUFg/KsL2cHOaHYlBq7sAcFKtVdsEof2MTc
ZN9kES2pUR8JQ//RxKfUMfQToWjxOLng+qltMDL6fXjcCqP3L4ZkzBXB7MhVA2actD6W1fFPzpnR
DYtkNSY+qABduKMadmpDzm0h88oL4c3r6Q8FDMjS4P0BuKJtDb1xKUWGImnUrIOQzd1p0zuG7hRB
sAm13oW99YzSiYPvaq9+X3fnzjgQRmrkEj4SkIHAMSVnN15ZOdMnGn6R+mn3rCbR2RaLuBydY5hE
4A6/QqEV+GygsM9v82VN13Ok88iPpaF26muP8AlbTknSMDqF2ibMdkob18fHnWxtPKtJ/Yl0q/tB
rv+62e288WAGz1AGbsTHOF1W/aX+5XeDJDN54B+uXv76kBZJDdAQET4UtA58nsQzThxMjlfCluUs
VNfLLpN4hruvosSHX2NuEFrwXRFJR7lKAY1ziYQpIoUqa80cJSim+BUTOTzTQZU71sNrPyHmV81v
/tEKxYpX4QrVi6Maf7mtS846fb1K+OUGYZnz52awgFu560yN7nwGc/mTKtC5MPPMZ58o4SvQfeQn
fvMasxW5ddw0+b0ujLZmm9VUS7mMeVmVD+bsCaf94yMypBL3PgK+pmowvPrA47Y5lNN7U0Rw4/lg
7tcwRoOrxEKmK3wh79Jw77PrPLoUz5GYR/K+/KTlrdihDCCGuJbLWPyo3r7wAkUagKxlYX03iYti
KPKDk+/hqG8ySMGgsB+jic+/pwdcxaEUu5DU4SLc6+dRWrMoAvT1qmyRK+4m9urbGPRx8P8i7Y6m
vw0EzLbEhsc9cQ4+1NFCocxhGa9bdFCm2PcN8oux5/2QNda3xLczQhycBMcgk0EKJ7Rk1QLeigkV
NZIZAzKCLTNaG7DKXqE2GQZIeILXFHSitbZZLWAJ+BHODqNOyf5XyGrP2Ry4B8uyUzjFaF3NeUfE
C2cIzLNl/cXhqiIIGulAV8qKlvslH9DxodU/nZLNOEOAhVgGwUWyEfk79rr5QRq4sA5DamvuUn0U
JrWXHUTZXzCYV8oNzgKkVNDkHN7FSIN6s+41M/LarByLoEKorr1Ads5UtABA9CuE5JoQHoPwYa+E
nphERffx5nEYv/h5Ag/asPD8D9yw/+l7aRA4uhIjLO6sRoBowQwYboiWIGP7EbixUPz0iJQkFijL
272pUXSZeu69H9I25k4mkbVz7rGtBiEVgca+siEAuhRJ6iGno0lau/0IxqdXIYexBRNHUNRoQGXv
P0n20zivyDCFDTtc3hvV4ECEyiSkcbeW94avyRsATr/3Oi+fGpDesQMtBdCuB00ikLRupnYnnMIm
eA0nhIhdbu91HISpiXlob7oieEv2aTwbyCXPVSoSptVWXvLbeBxnjtmaAeJqRRrrraiLA89cnpd4
n1g6gA5INDj6OAcVnJ4hqH5SMENea3rPspF0Ld0j8a44XngbVUzw7A5rNB8n5QFp95Uz02VqcCrq
qn3C6F07uQ8VGcKqpjn/0IMvtVPTmbZTXM0OtJCX6wZxmIEDA3uByMOu422bVdut2ZdWsjfv7dNI
awX8rYyhzGBfOO7q678BNhoz/zUm1Yd69roH8Ti9DL4chclTCnVzAnNDKo6nsFeQR8tP0OHL8O5d
igfMrXD01SN3PWXYcCF2YkiI5WAYtwv0A79Q8u7yhjbQKO8B9Es8IAy2npI4fYa6WUPprtm6H4k8
7q2uqFOoeuPBwuALZME/N5fEQYBROSHbEUBpvwDEOvS/8rkl7pWKc/nDWiWh6h/YIZ6zIhodZK/c
EtxO/66LkoR65QQbPbTmEbH1Rzo7H9/iA3tiupAA+14u8D652muacMu1xG7F3ySEkTc6QSPaCEsx
gBzFD5wvuM1RkTY1wMefxDT/xUxZKll75WZo4EUsgrLp0RkoOUoOip7WxOTXD3r5IPGpFaHTgyKj
oNC10QqHDqi8JPAXWP5spLqEqyCeeLQxleYrhSBys6uRQlSKwG8q0VqN+EGVFgaHhS8TpcLBi+lT
XeVLhHcblWAScXwD8da22X2ZBx0flS+lKvqx1z56VVL1trCXkYMUs3AvXFSBJj+YmoqI1D9mIccB
ay3aW66A5IESuZzDDw7nJkS0nVrOzCp+oJnxdUZYTdJK/wAmYQFPTCnEZnEkzBd30sTInt0hrPvq
IW1MaOsgidapDReZ+TY2Bf5YjeKKUyZ2tU6eGnIkscJ33CN3Grj2714a1IvYweO2nXqDhVmvF119
aKtTPnI7HKLTkqzrWO2SXIB8fHjS1PBHiqE6kGp63Y6w0dS5jFhgHRdVxb82h48twYeSU6UU3MGz
dqRp+btY55RlQlo7Bwpmv5z4ywgJjD8MVy8JX6WQNVaGJyvvs9uBHgGlGN3GrjLnrmQqNqUzxNCK
Ep1OPHTjAL827BFuAaj5VEiLbVedCSl+++VWepkL+AMgNcbM5OdEpueOWrb4vvSucNOWMt6HzsF7
U06QevjUrTUDHGK86RlAqFolcWr1dvh2dfE0Jpj2eIbUTX6MIupJ4Ck7TEfirKCtPnvoobJlzlZw
bZH6Z7wlS0D/HCb733MUnqIrcQ0f5H6kjLUtoCNyb9X6twfBgVQJqORaQ+oJfAYcvJeuFSOgs/fR
ox0aegcxz3a/HXD0fZabhOYbCIROiKaKcneREqy1LxH+RC3wcfMlqggRTlSWhJibZVBsdMZ6t1id
fTGap/IHEeBjFfbko85jjjSLmVCqjiGa50yHBNvTjbYW6lPH/8Y/xEWw76sc7W84C6N9LmI/lVJ2
TSBNIw2u1LqnmYJ96Op8ek7c8RQ3UtYfguvwzVV/KXUc+D3UjYeEHW7hM8rF8OBZuniPHeiik2M+
vv/lsZPmNh8Nq/l8gQaWpWJ4QuKtXCZ6uqvJZlHbYv/vUp7gNonzkoRonTnCvbJ6DuvahSkNwzxJ
xdq6LbRCIg4nCJ7wy87/GRYTqjeaB0uIZ/8vZUcJEAyvEc1lP4QGyPXzuY05RLyiLIwyq15ECvSv
ZAoaSUmmjKn+VxhRTGo1GqTD7vbID8MiePHRKv48mq7ccTChQPe3VrpKbb3h+B7g1cp4PFX5GsjT
SY8RKt4liPpPBg4tDtcdxAXDUCDrN07xGjYG5rD0xuTI4371WnZPbqMQ1H6D+mxSzJnfcSQwgA52
rIQ+t0uFAs6PH3Vg6gBm2dGMMeaCC+IFu8+yrkdonA4xFiT4WASWP00CIhWuUFwJGxPwdCxgvfMH
KNQc5YrSo06obkjDFS/4jrh1/23LHlfnQoWg+SLeXvU+Hm1KrXODA5QUnZDJVkxy5XuT+orfmWPQ
bJJg1A4GGLPFx16yk9j6z8t8Bq5sfHmPc5iUyIi/vomqiLwGQV6f03JmoVjP96OZKvAx9lxEo+JI
yGdZ2zNGGk55XbBITGKrUroQkkfnvf6Z66fL2V8WAy801Q9xDODreK6cc9BBuHGdMJxTrYPB4VlR
DyIZk+Y0wSUzLXwXN/fG1l9Z+0i79Ck6gISAK8m3wOzuX3J8MqhGFc0ujOe4Rt/1YJSGzHm1Kr6C
SnmlU/6JbYarozafPEnViUCxueCoFxFPpWrb3wzdT2Dxud7AZ47PZNMyGq3R6NaVzQn8pLXwqFUE
1wUNAnC53AqckKxf3b2BmmQovZog40E3KkxpYzSqhNWdCWS6aj+s45vudN//QwTy7GR3IAu5mv6d
gL3qvwjUcmdsBSqMrBfdRRxmz2Ux1Z9wExidjXl89Vos7CFXo9T/ExQKz75xFZiPbFWYJRLB35co
XZ/6f0/COSbaWiBB7vopfcSCuggo6F7Lj0VtU9kpMeMZVfqh9gTGlMrF6wn+5/eQWzwfUYmce8WU
RjE2Ombr7XfKEr2m8kBxKce1M5d6z5ZlZTJXr3jD8g1q0BWIIpgcq0IihURVcGLJ2WBBgOMTxW/D
6BsMuj2WkRZH9eXO81eF62Tj2QxgYSf59sJMWHMWYc9oeWalpeknj9wCpTV2oiuDw1/3eKRtUlej
T99CJ3U8me/5lzyWhvNRkKkbOoewy1MF3e8uhDvAx6PDlGFP+Agg900QKxKxd33Nggx54zw50YgN
Q7A5JKMYZPxzwrQGCHz7GS+iA3LRRaKBVzJDQeBkeeGWNWiXIV4vfo7ETk8/I5FYF8B5fP+yXtzc
r8mjx6S5D5CvlrCcFa/6ITwkAxtY+nNOkVYT2QEouqiqHE7ZXeoNHMxUVGwp26MW7Ol2EMqqtNaq
+6MlmpK0dyGNpbRVHsBdsgRl8zVi2uvROZ7Sc5aPRm+gOyNtSOQKRBipfOfKHwYmGcJ1eYVtly//
csa9QN/6hf0n0ltGNQGfn2G0CuzD272ng0qQwcBAXMJZZhA+5r6bAn7ZUolonHVp3aiJ/lQR2Of+
N5VuAog/vdiZ3gzUC2rx2uJjB4vqXbKHlZMiSZ++mrz3AOmJnS3qFvosTTxM3IzZMcU3reUxvTmK
XfzzKQx2mEzB0TGmrH0mn8mw1s4b9b0PY/vCV/0zHRUmCtj2XnC8b3lpRYuoYRsXHiM7JEhruV5A
r2RJWD4Hz/PmZkgrC9pIgSfXUPFKbNxIq2dECEZULcoTRVYKZlHfk5i81ouDjbgMDsXWz0A4nJxE
cDc/xhusQSuCrODkZ9AHnx59+NLhXP/Koacg3sLL/O2tDLX8sppDJUk1guszhCSsYsrc9otTpDcS
f0YS/RbAXSYxqgLuVnHwpsdaNvczEPopMH6CiY4qiuCNS/NrqT4GQYknEyZrBg0RuiwPLKzCaVZo
AWxh41l9QTXEMIJszFwPv3PTS/JNv9X2VSFOWhKsjUJkTQp1P9pU9XTXf4rkBq/5btflN6B2ggHX
eyVQz0qHeYq5pMAJFxUbOsKls2LitjxebD9Xrjs/8kehqclToUbwvebZlPCccjqlzePiDCSUuOm4
mH94T6A5N4JvfK0Pmv6mNHSSMb5uz3kb2IA3DXF/9TLofmF6MJAPg4lRS4SeN3AjUA/pgctI5wGN
c7l5Vgvr8dgS8LYG8CTQ9sFkTBwkmrgunuYKu4nBG/kMj8R9AT87Dy+TynMtbNIxjn9pQj8AlOdj
hsUbKxudLyKo/gZjWgLvtzoTsat2pLF7MmXc2vpd+sxTCTPJJgyzCfUZ5hIX57iB2eaOsgluZtMw
y43yCv+csd58aTgDqIKAdX5/g9dg4rAkefaEfdp94gFOBFIzXtDsQoMay/Hq8FaB8AZee/Fc97Dp
zk8ID7zTE3225u1esYL55oww70E2kf/xPCxQzM1ZPyoSQhQh4n9Prk8+MRwq1YR8ftea74Fwr2bh
vKaV3EDUZJD/haL4Zy6SrfAiA+wr/VixbMjamKqzPdWIveyYRc9ItDyIBqqB6WDZVx88gJsglxly
vBpQlzIelnbXY2AfrsLm2FNb49OhwHuYn/4baxPuRcrxEDkEfdQe8u6JUDV92GofpJh5VxlIDy/G
u76N9MwM0gSNZjuAYP2Go/VrC+TCFtnC4KRtdSPq1HQnQALO/ooBBWIuhzvcMt2RujJOWgAVCahE
aOcalZmN5SjmhpD6q51BG/zi6rSEZAHttvx4cFF6hveOVW7QMCZEZ9QMv6OdanDoz7JfM8+3izaV
bTRaMk+70cwB718weEVO6yJdax2cWoRbKHxzlJK1W0BYt5qaMJd2AX5wY3gIUC7lbW2Jv73yAhEk
phNR8GT4LAj65XB7chauZnSQ9zso8WJwXagjmWBSDhGiMUb7c+y9RPheoqiJHQeBhhhgPtllNDsT
+7WiDSNr8zgMQOyhufhFfbZQBh18c6nD9FcltF8NrvjNQ8ZM5mDDTo28u9C/xO8VJWZMb1zkLdVq
pzB9s4RQrAIKKDCx1fgd9sKMBsfXRvFJqXSC085Zoyq4gsAVLTn+rZIXWy+aTETsOHgpOmYEc0it
kB1kqduCCnhwDYsJ5hvvRv1BXLCjh39rHvBvJwNMvt+Tqvd1MJWtR4G5T7jSy1Vg4mYH2Xe6NnPC
Ca6tacXZ/ZeXjIP+rwdfYI6Wc47dilapRWJNgSbgFjGXT4YaIwbEyrrDAtpDUKAp10NXIrmaJyM2
ivnXGVQpLQZs5P+Aw6Ah3vEyIFj35bdFbIOmGu+KOcMOWy1xsGojJZVjSNPMnJgtXzjQ8zXH8+RC
b/TrxE5nGkyWQ1+8WFsheSgfxN2BNpavTdvElUpZcJ5YoLTL8o4KOOmmTxZaTsmZaex4kQ7V5bKs
S9HmMxUuz1rlQHxIN8QmPge82rFTOQMLQhKELG+IbFOajwstF+sqVnvh6okXsaok4SWXOzTBB4+F
3n85LWv/ah2eciMSMlsQhnwuaLmUhg4Ztxtdw78koLbMwBzrv0Boh6E3fDRCADh2ntvbvT5BC7Gc
K8RjiMDy1KOh+FTlSKsFC/PmRrs/WyF25aEGDSJGGPzYsyn8wF1g7LPK9eU1tTi74Uj+pLEuG4Eh
KMXzKLxaWXz+XvR+F8svJ6WmSBZUIUYzN3dT0jzQ1oMEIcMMFu4flqRxaXSYDX/i9yWyAP+qCck/
k5pPgkX/T4z+o4mrgowV+LsjNbqjyPxE/cdmOIdHZblX6VzXJBMYsnCqDMDw58nswVOwzn0ZZUq6
Xy9ZPVcAP78PJrdDtGu8vGq41pk/S2plmYPwUpLNsLL3eG0D5X7mt420PaSkmqdR/g2USK0OhQ/t
yZbO/hbQ6sa7264emp8OAle7uL9acME3gMSCSlObeHozBl1NY2lTXI61+eZrc+N2/GOvmlAUj2tC
UmHFTeFq+VFnvPjBCxi7PrNt7lndTrsJcgyzyg8Mt88QxFB9ZJn/FDdyN/XWjVvAZqabjET5i96x
qjNXgIbFQghwwY/ZxfsbNseAITti+elmBwyh1EX5SsEFjWYjx4eEDSUaHLTiJCnHGcF2NE8ss4gs
CRp0ilJEuMRlYBWB10qDyo1YBDTgLkZYvlhwzh5POR40syLp+kaqOCGjfwU1Rpj6Vb7vlgiH4uZo
zN2so/aTxEfb8MjMzhgLCIK2jam1g8vt/zP0czZRSF4QiaIIPHtDYOrClte1ze1p35kzdsXBsu3L
hpPsF9wJSXIjMbdYgdxfOA0wvvcO+wqASpByKgmxp9A8ujQ0lxEoX8JeD7U6956dgTp+IWr6rxwC
1d17a6sTX/H+SxFXQL32+ch5wi8CxlZfXEvjVkvDxVSntaunzX9vyHZ4T9Ry+53Yo5XK+vLD8tvc
mCRWfbySsnI8bt5ZlsG/xji+WW4DrshWL6dAL53royiuSJonqWTLhDu2T5TpPtV0OT4Nhkiubefz
MojxDs8yFGyLaTojtmvm5zjC7KymbRxYMgkqnmKlUXl97K13kiiaFjaS81GvkA+hfefNOXUKdwoL
onKHTylKQyPsnrwOt6JrE9MCho5tXhCqBH2sHe3ke5V8jitblrIXE/fNIc+ICNywjrVRoZrGPBDi
N7yzCbnZnCqLDhXS+t2WJHo5yxScpaUA8ojFgHhW9q0iEUJcz+gcRyjwez1hFTgQ7RpY08+yv/Rx
cFjm/gA5diFjCepwve4lheGmIGommwJcD0X3aq6i2EUQZ/cO8QTbLpx6DGoWf8D+P03TZh1FSf0X
LifQqnC27t1dDYtTp0AGy5LuWsp/oZNb1tl9jl1nbBVsvn0DfcivpbkCi2xbVuqKuZuhDZZomg5V
9Ubz2IpNeuWk+X2pXNPNQXlYWy1zdDV/UXcrGmJD4HHT6rq+S9V/RSZv8kHxdOmtUxL1fDVoWxnB
5B19N3kjyYSeGH804NkluHAHgnjbKRstyxGm7FZ2aRORCTgIBxXRyrhfi6p0qsCgoOWs9bskU4we
jW54bpqgNDaKduSB171BHQ1HTF9FGXfEj7SgaE2T7lucvCoInZ28rzxMlKb+0eb55t+STrkWh2fj
rdjxGWXn4oR6wuG3RATIbouSpHYi1i3vP+RoYLZE396PyzEb7LLtGQw7ONxfSt4cauMo/RIhmuZ6
ecqP36wZC7z4+sWUnsKJb705DI3IL1O3SXsVBUxMT3F5SqIOdx9F5M+gMnY8+163oXoF/0wfK9Lh
fslbcYpz+3wdoKNSnSD6LFg/2s9q8g8bLTvGwC3Z0p+AFfITF2nhd1MwuPzc6tQiCNgkIk5MtiNZ
D4s1lBTn5JFA7OKF03xY46pW6h1uC7yLOGigY+H1Wg8QvqdsF9LqiE2SV1ARca9lkoq3aow2Hlil
dthuejsQ1FRr5Clp7GIv+ytOaXrY+leSSFFxY8oW4TrA7tXlvzpuXD0GEubHHhBO8E4UnjjoUQkm
sgrgTZK+8fruC9MQTvNfu+1vqMAUrtC2yQekrbNJZymgsMceCydbQ/ohwQtPeTMsFAjbo+XHBxYh
ctUedNhueN4vn7+tJkxt4lVQa+hcY+4CQe1wIFm41jRUb4hpmeWsEq6YJ2jKFmADQcrpqbdDPdHW
32xeHTqfRRvH1ZFXUgPpUVm05ARAemVvxDcNpVUWUcilT7SHc1WE3HPfw9/dMkzVOHP5v9Nqxm5c
HySfdTDo3GF5o4SF/TwkZ7RYmnTnb71QRhIn8AyEcpiO3CKy6AbGKmnLmjmvfLO44PAqqIicI9m0
Zd/ui3c82bwg7zAfLnEWF6MUrELhU6QwhUfPrXOTyTDkj3VQaVNFjNeRkNtW5GW0ZVOfOgYXjIln
Q4g54IT5ykVJCzy1FgI8Vug+6cwyiCOyz+ZyKgjbihcqy8Z79XuXZFg1ha3u0hw0OHHlB2rkIEbl
qFZ6X1q/pofXCsppSx7/KyeECnEY18ITCBWHzupj+WZo0BUl1u0FfNU+eHGJH8hIDi6h10Pfkg9e
g15eARrNC4Ee6UBQCu7YqiTFe8PFsSp4Tfaeh0jZDwf0eQV3spuvE9FA0pzqMT26mpulPu1F9Gmq
eG/Z03iw3nRxNR+fiZvfmmsflbvOyOl6HfykZ7+7uX3LEAbcfWNGDXDWjRMw1LfJ4a/wxyQXr17H
Qwi2qNIBJeqKpKW3XOyVGesUDl7+38PbVyR0bMwT7XV8hiDfyvO/F2bEYKAX5uD6h8uHfTMx4aeJ
Mp4ZVkjBFbLHeVEb9Ipqt4gQ0B235SyqmNIKVtEpDtzE6Ujv9xGb+KwOWBeoDd13JnQ6KiUfh5fj
3TTOrlsCzQuO0z/Ddg3MGblFD1RF4MUFt86EoU0ZW7NzlpW1kfE/hleF+mMcpGcbFupi1zkBkiJO
Be1tWFy274blnDP14Lxa/DZTSH8kppgGvw71Leatc3kWRsHIrHzcg66O3PmpFTRk8JSXsOvkKDJZ
fG4/au+WUWVQ6U2ofr/cAKyyP/VNWe5awpJgomDR624SOaBJ9oAnlh095XAeAAJXstFcC4ioWKWY
RsMsA5efNIk69FLv9NVdpXa8M6FU4T31tHziLgawMyYhNNsCGZiKJKkUz5Zuy+MhTnloaCUgZ5Dz
3XSEV4qDocQ7h3vnWsezzQ5ycedJJYR0BGHR4HJcAbC2VUnGqYEu3qAoCDLaUg1yHmFn1H5jpJzy
W+TK7EmhajKaLd9KUjXghT2irbA7dy5cJl6F5HNsD3s4ud6pv/0swdZDNF/gVZWGv6i1hy6DL8he
zoRZJs5GuUJQWrcvB4KDTGGkH0ElL5AQtD3XtIFb2+XYKmXezRNlYpj+hW2GVLzEH/8vpNQ+KzPY
xISlv9x5z484St5BD3Pe6Q7eTb0wxGuyPqHuYxUMumzz4yrfmqo1Ip2BDxRnlLq6g/ZcHuVk+jbI
Cp4itBlb3KM7qIinmJpkVW1BHE28L6pL2w8jYvPAKC8Ikosh5WMN8+Dz9yvlCmiuZuzovUnwoCb5
oCMOJNwUbVbdmLWMeEiuTfvOuy94qhv08dkTN/NHzxMFCjDlnR6cUqF1k3gRJo+BQszjDTSJJEoT
hE7T8GV15ix2dzueQ1ffdXcBRB5SNpp4hwmK8D9Y3fjvoO8Lgg8teQL6ShvejnhIpB0l/nAkyvyd
Dl7Ay7eW3PxzGfsHgP8rtxS2trutPCg9UUmGaDIJiHQgFn8Hiv6UO4XgRt6O0M/3jh834KBy3gzg
KT1icQj4N1dfqUjEc51WRBvcLoFyff+p3fYCj5xWC9Ru5GYSXPlc+7LRtFzBkBdYP/3wgYwbgav3
+Kuf7zKf34s6Trah/+3bpRFlX+t+CujZO1ChX9C9FsYHoKzNY2smY24yBKJfn1qHU5NAgTVbJXUa
khMTlzQTLwmH1Zo7JwuBull9ttDZdYY7yd6jO+nCxnSznmnPjyG/r8Fh597vEPN67zpWoA3Txfqv
Vw0mHNKKimib4Fzh8A54Xc5hNmCp4ZKjRgMRTGLwNzjr0IBaQX44gLasf34zww4Z/EqBXDT7nBMM
OpuDyug0Htnvj+QlX//gSNEc9ti5r7drXWC0ft8n+IXWtA9JYw2CDWYPuOSeemRxDGIQnCerbOvQ
zifAtueuduZ7xaLzxcY5awpB7ndWECMA1oUV0TVMG+T+DdzpgxblPlEZLYeQll5hDeoiQ3g+ZpvU
/TUg+MG/1lScaKnq/0afGv1Ac4GZvTsE2DnUJ2H9CHn3gJ905uNGacyLXJVxOdjf8MbdRw9mchSu
yWyLaMVnAyjyVcQDMJe48RB8BsK6Zk1piZWAOhAT7/R9BrwEmjjtBcxQU4uWH+OaH2LCjbKqelsO
+55XC0hw/oLhvoHOJ5lC6ccPA2FoKHQWqFPEEzV2UhVl3pw3YSj8xEZQsSt/DjrOm7/iXfaCvvEN
Vx4xb8v0UVhWmxYpl5HPXBProK7f3rVDgkBxHx/SlofXdJb21nojXwPNGL4THur3/kt4BMWTRtD/
iAZ6FdkFFeFtdJbODgulwpLp4HhFoYchXuyxhh8Kcn0F+Fsx5UuAsZWQ2DmKO2s3tE7O0zb3t4Ht
di338ZOIqd2ZdgK8QIwUBGsmWnjPBt9H7kjNpY7CSnRLNq2bBn5131a+t6EQoPw9TdO08s5s0XuQ
gLZ3BZ63ICG2mmz+VnI1FKGuSvU2xDuBRrohksqNUP+ypU9G/MwgtPKQX+VzCgrUt9LkyFcwTO/p
raSin8zd1jXMuwrQPIXtTqqWtX4T8i4adEYS7A6/yV/FZSblRLO34dg+obqN5hHY1d78rPdK7hrV
vQYF5Kg1b0Hu+0nx8e12zWJQvlLR9artCof5WfF/Aqg0nkp1CpTjrhm29gtOLmKHVszRTG8J+A4A
wtYbD6aIr7boTc4yR5JJY7wOKzYT0FNjxzJmyXRxeiGUuOOQ6SOWQVzQkpgTAw9P9PXn2M43XOjU
J54sRzejIzbd97JMTUvA0oX/T6MHJ5pziALDbvqMsAyIioQmX0Y8kBRrvajCG1JCr6xdF8xCGG4B
omKl1hb1l2gDdM8ay04UG4Occ+coWMnoRG8oHxrgsc3T38DBY16j8rj8lMarcm7PCQLVSDzWvOgi
ys7g5pxC10DxFfiu3kevYptB4YIoJ9l4UFFx8PbLzXDw95JbOOVqroazO8b8hViQ9+oW1zxuaWOU
oFfJAzjKjFLYsh/L30HaRmPvgExX6FnCD0AzuVNg9upj8o7N9S09EvfYmPkxHEsrDqfPe7VFPM47
7j1h4Pzu3acOR1x9BGemb+Me9EdJA/5ugLhn8MD7mWJFX2/cBoygvC0GMMVCTIkXYqihiEuLOZ+a
MELE9GbVrqnhFev/Tv3oXjm9k0zmCKd7wI3danTaTOrRVtYZ0RvwYL546urZogFCoY0VHZCHLDYu
3vw5t8Xi4/ILh+m1jXuZ8ouhom5fR+wAAiaPA1oPYsbWDUdcR+seRY/QBt5lGCiUr9iRMtEF8ngp
jIVRYzdT2l6H+jgOUEN3HYhAbkO+LKRYs8nImIbPEYLonJDJWZ9E755ltPm9iRSVlRWu7de3KkdM
XfZmwcW1b29X/S425DFCkWKjhFTkL1s5d3cm7Rep1PbcYAsjWCOcrDxvPIqjh7W4scrI96a7VZL5
x+MVMFagbV5HoxDaayK6PqFmiDNanMEujqvEfJtlYTwIZwF3WgZXsA84S3tVRpRNDgc14qdKlWLc
P/CCWtY2XTnAx8X0U9fyumR42yycnq/l7OUIowXMbKE7l/i6cG4edz8BWx5gzOgWrngPH/xkCZAb
tyT6VpOR67bR2c0kichlP+m5YelWjjp1hBia63El/7Xq8Se6A4yIIm4rYsirFwFWN8yNiaX0T8E5
FgQVbBBNhPwD/Lyi1B2+/QqRRruR03Y6A4vJxg/mGoLUG5IbMsZXJDOFBnmjpmD03EPtJnqg2Gud
hA7mpwz722zJFf6jxg5duMRcEbFKBtJF9Tb26P76qELxHK9lspnL9rlm5f0UjLSpJtXmK7ZiHv+G
y4KulA9swgMkJZAqxafv86p6NKEV8RxtUPoWjbe8dRERFhCIqjsVWAz34wjikke4Id7nqmaG+OOz
4vCCtswkrZVxJm9mf0KTzPe9qHp96epNSB0/QURbwnpsJNqWJ1G3ar0LKFt60SsO1hYsEqXIbd92
WtE2q5dRosEO9cQ2fbXfi1dmz0df+qBDVHIus5LEfq7O++TtmXcot4+37lo6htKo7X7ue6hZZsJo
SbJNSaPVQGGlNS/zvvNrWnEdEVYo30Vit6oAzZJvFj8dZ8x5RYju6zM/wQ4fMtOza1ZbZoZ09czc
CuVQl2LL27QierGaim10N63wFqgcSxjBUm4H1829fQSl10KDYlh+ShNy/Jv4TAZp4Cj5c89XjuF4
4YFoMN0R6+UxTKJydyzWKFs+W/JsxNqI2Xy1RpH+PK1fpQygr6jX0dCQLRhkd9XVnKpWGgaWlout
5R9GzjcsFWusADHmdSNAtk13Vr5JjByCIrvemr1HViTQlgbYVXDNj7RMo9Ib/ePlNyI+7TXTb2fx
W7rjbBFL0slxCGYv2fyVwftlqzjKwXDB97bvgzCpix3KqmmSzZojh84Cj7+wdq/FGspmt5OR0OMa
sAkpliNV0D6FGUmbKN4Jcl+idMFmeb/DFnV6LH4v0TuXGE87JDHr2I+xmzJ6BPdmqS818HKRqLCx
WIl0gGWKwXzUIRXaDoFfZsBuO8ODJRa0Z38GBXQESBgXv+khrmYslg+0zOyZCbZp89LAvI9q47uv
EssQ0Mr+DxmXCJXtgk26yP5sSRrwuiimCtbk0uVooT2pFDX00/f96QJBozlMj034cn6VsqVbIDo6
alxNARPYUn9NkuPvvEkrtu+/GPfZbc6uvj9BoBjtKTkSNBayKG7si9CDY839DjTKEZGLQzz5Kce/
nd/he5756Umwx8RmUhLIZY6O1g1L9WzP4J17VwmXZ3hr8YdTi76Y8u+hBgKjIQko1NSMNBE1UH5I
yIrWUECFzCeFK/VQrLSpFR2ByWK9Vo9RUc9Kx4J94JLXKIhkWgAkqBXXkhXUmlNn9ar+pkdTbULN
j1hTnnCibkN51Za1jFeFmXor7V/RHd6K015O4YUfLpABzLeobDzMTM/hJ95cMA5c4SDbjpk75jDX
FNHMUZIcCq5VlJRWjD+ZDP7q6a9wZ5zUzUAtfoZFcvX+RL0Od2KUIhTqLAqpk4HMF1Rfm2UnopO7
r7CIReVFKVr56PHegUpeiDzvk8uJ+oOaRHgd9dDIGmOXEd/6Z9ghITMi3lY9y3XhxGapdbgwT5E1
KsCauPrSjHvuKhh7s5EpLAQgJSpsbKiWICuCp6hAqkkz8DbfVycpL5Af9FfaxOTb9TJ20LkeTTGw
AhsnX8AMDdjmidbZmq7YcOedmMjBqh/opldhYOzuwSU0uHxJFUzxw9VloDE5nyxq9n4ZwewSGRD7
7KYUFlG9VdeKxokxRxvxrmt2n5qazCRvZERj25vxrLDjDj7x/jfh4PDxBNN9Nm+Z6x04i4VXt4cx
NiyxbC/ol4xf1dyHK0cybRWCg/VCP15rFFwun+N1M9GSvCqALCUULng4q4TmgTJ++pH+qs1nitcI
IMlwXeu3Ka/NtdFHFTtPVMFehD7r32ZMp/PRy0vRx2FxM+dVmKU0KfposCoPPGAMmHpv3ijigerN
rvqHbgnIOUcpaYEoqxc3SuLUTPZ59YXVaggMCmUikLB7F1Qi+zGUsyOnimBNklPLbZlF6/WOhQwu
T+RTiexbxQ4G8YGM1I3dbLY8nXcZtd8H2s9wY2otipFZvkI/mzECEHPgH9UM4C7XXk2CJd0pfxEU
qYNB24pTdBPvbY9FfX40QInos08Ha13ZFPhdFY7qqRZqk+xHBsV96UFeohf0UvEao2mpAc/SAxhW
uusoEenEbrQ0fkGDFiABLr88k2ylvKYGpfX1WU4FPSQnpy4u5IpdZE5SMTIPFpJUyc99U0nAFdoe
IxDlDBRGdJfO4XoNJEf4TQfF7QgvMqBQEwVa0XdlA1FTGuxh4IgpR9Ns32qwXHKSgUfmPckmbxkg
cvMN4PeQa0aCYUgs6tdEqUJ9rOU90I1jpOCnrTR1zUhPbdJ6K/Pl49JEwWTR2RIcFVbgdZmYzMZL
dkeAkHnCjDfU7D7L0MSM2159OmxSzd9f3Spt/ruhrKGywJR9s+RV5RXesjHyFzNn0JaIADePcygK
sCMfvCpjVXlOOMmi+3Cc7r6v/vLLFGwSIierNhBhQbqWguBbZhcEl6X2Ymn5b9HEvGtjMieWP5Iw
KXNoSVkCY4ZKEDUyiG9r4t0wiq9qdja66Zf6ysBVqpCNk3icbcSFqIRarsc8zIAxTAVV1V1yBFV+
/NqL5zMcnwx7I3zHyrLj6R+zhaO1EkcskxayIk52Dqu9yu1wMLfKYf31z44P7rTdAe65R3GcydgD
x4Fc0xo11w+/koBFCgICkjJoVycko44V/54px7drUOetqVi2eU+PNFfEQTxuTw0zwLFQdA6kpoRI
jahvT/ffnIyKuDa4LgJY/BSXOS7Szucg7FeDS8HeHySFiPTBW5jQ+ecCSWFZfg2PGQQAUuLf5gLw
cSeXuf8OW8JYh1eimx6sma2b0WceL48VibLTgPhAC2bx3WzpKuJSSEFtMy52HJ4omwZR9hJ27rfz
rBsaBuNjq79ajTtl/vH6eASboZT8u7qt3Rjkn3mhektcA/f/nkT9iW5poi0GJwTewahKyOvpsnib
g2hMsC8tttlrdhaa/sKKerGEGDvvLxzy8pBuDGXt6fT8ln9MkgrJvTKRUqQF5ImK3G82p6l99Gg5
UyReaQuuqHr3c6Yjbej98akxxoJASk5PQbiz4rtEO7gRyoh1aK6SBFNNrCfgqguC29PgJRfMbDBw
4X1ATYsV2HBQP+2K/UsYc4wscOoTwSrfmWxcuN6gnKFBDzm7TzxAoAb8Rvazx6FU4XSJp8CN3+96
Yr/AbgK1S4PD6jEqbU0KdgB7YvTtWarl7qHxCjyBxwZiPCm2JPlG7O3v5r7sfzPz3LSa5sdbWBwn
eHFMgIx/h0H8XEzFYUuL4SH3fYwAkYf8lBfLmeXX9ywaoizC2y9I1+A4lu33LeLLWz/BE/NYidat
tRW11JqFVbjfnLlbjzlTktU6cnnlcKHbx16jcWWd0HcwHoUwVgx5SOa/fPm3xnkBwNak+PGG0UNv
80igEVStOTz0zdfChQbuYFoTPP6aNzOLCR0W6dyvNdWLWI9y9fb6OKe0rwtg+ccQi5ALUrmYHXp5
jDkq/wpaFozvX3SGBZLu6XcTTPp7B4OOsCx/epUqtOKFIAacGnLU2hFogb4lEp9wrtxo3lKXo/6b
Y+1t85u882rH5Qu8RqDTFRAq+ByeWzdPPD3u44lLFnxdCT9d8WfBe0L9/xHnXrYq/LLYOl6xuz8V
wM1+S5HYLmjzhZHL+aCWXy0xRzkKNF67WqJvcHu4ymRhDQj2QXU0q0/yfhuEexezUQqUwAcDYcdj
mHp2GJ8OIrWy6ogJpX1+mX/Y/B4CY4KHRfJkLczP3y/hlysQISASHG3zs2v+pssVxT8BdI7ESFov
PIXRUG/EYTkiTZ/oPtUyBQAb/B8SPQbJ3WLMNBX2ZkccKC/OFtSyObQDDqV/45SLX39mp3K3igwz
yZWDiriis/PNNbD7tPSzizpDoiXd5ZuhJWPi+FjSHcpamYt/G54Zq/kj9IqImFUjLdLn63VKRRMN
AxB6HoypEBFV5W8/hBwUrtGEJZWZfaEqm69AJHtl0fTcBGz+2ASG/I84udz1kXTWgmo0FmNI5TyD
tCdkYhvK9Y3ollgzJlLiyH5x2RpDGERqmx7h2MgPE6quXZMRfoqP6PVnEALR+YUfIbUGdSMivhc1
sXIhclbQqCBkenk5cRu3wJKcwYuMCcIXqmX2FbEtg9VRkft6OPvjXmqfrwCX2IbLrYG4D289zYd/
s6Heja04ibI/3WShxlk+xTMJwQP5YReD2uKBvqZLcsbnrA2VZmpQUyXsTOsIkesYOZJ16YFBv7wi
yQdB25fcvE/I0n9OkJVGSeo84uNrLEhebTYb+o5frLPZYb3iTgXESmDy4aMVMIArPKUd9h82nLnB
14L93hEiPxkHulm4wCzZHaaocrRjcn/NUBh8xaMQuR3M+lIYLDDmEuEytG8L13TpeFuMgw2cuxNH
i4hIf2BrqbJdpKtxnuSwtti9gmj+MlHtdeW28Unl8107PRE/AJ/ssNccV5C0lQNBfLhUuhThZOL/
ySDTF5VJONo525QimJH41ZXWH9vsFfScltJgIPc34sEgucep0x+LjIAB3H1TZyb/WTxOjLnkhLSh
BbNiuqgSnz9a5bHUb0v7mg+ojTMjxPvB1iWp/nW4AhOHmqFauxF+vE8zQMWvcQHPbRSPUp1rdDjd
oT2bmMtBzOSO9EhHqRppL9lmzty4d35P+zhtNLdGQ/NN6iURLHSJV5XA7ni3lKvW0iI8aWlUWuV4
4X2R8Yd5q65SC52BBJuvGsN06+IAqhdZGQEw/Dyd+ytrU5WwUn5Ntf7B/0GdBHOruzbIgkq4j0Xi
tB2zpwlF17Ld8Eoh83V0adPC8w/wZf9YKBx+V0uBV8f63b4lGMrBX7R95FwPcIMOlD3uFkMJPc+/
7TCujf/e/wiXAQIzdpUFJXFk/AMx8hopQXry/hUIvreVGp9rZQj9O/nuyqEAB0z4W7F/hBKDH7tX
eWqQB9cog0z1OjA3YNl4Hw4kof4hD3nOOkGfdQlVHgF+MzDipqMx4TwZZV7XyJHfFAgqsXdHtHk+
603RJCdr3LUN9Ub0vXbk7cX1gOhyj8+iEHxXVoKzkOEVIVuCYyWcWkkC1u4cxss6/UvdfMBcieRZ
blmH42pzgZeZX+eyxs650xRvp+21FqrOvd+0gTfW0tRmNT37TkJ+2G/FWm+VJ2RwDobr0oyoUDPo
9O5s3HNS7QzSkaJlKe+wraKCULlYy+wVF03Ae47tai/nEceGZ9Om/zhxFyVGo9grviYog+sBWyz4
sOdEErywFvhFlzqocf7LAFjFnzUkcOX7dAnymFiQt7iHwSXCnsrhrnuEBcsShKIvnxrHN4dTGH6C
QNuocimY8CX+LfA9579hwcNPD8loC96DFytjla+jdEjvTOueDrkHcab6sGWtLjiJ2OFlecc8ygNo
XODSHOq8jgQP9xbIKbO9qpmZuqAt9CMHY4zVLftNiibb1EX1Jy6NgySUqHe1zooRB9ini15MyLcF
KyU9gOf1kVcAxFcBSPvtn1DS0Idk8toMSRALPgkV6TdXhaL6LUdyRwYaIiTSg1cQhrZq85F/R/53
LhTtUce2faTSkw9ubxee/x2QoOK6U9d26iRhsvq0uqbhBu71S3BBS71oQ5O5PRG6y8YKF/XBZKyS
ovR6lObGv108ppTPUJcKgPsxsfnQzjH8IXIppkbbQdi4aD/y3BQbky0CkWzBltnpqMBslBClZjdT
TpN0AneSAvxINpaWgB85KH5LtBtQQxDl46dWcNeNNQ5gS+K4D0rkhfsPJ88gPHE7WpwfC6DA/M8Q
E0/ESWg48TJop7megWJ1VaHcLyRIcQLSONxYGrQYgpK9emLjxJPnqYzTRyjD62DDuAFyl0FGn8Jf
PVi0DYPFv1ikjnUmlEBpozLOdpOXGkQ5Wg75sCuLgXvmmgkQeinbyV8wgSptkYbVZkQqPzKVpBLx
hXT21D1ZGwvWMkVJKJyBR0F5+oFJfYgaJ3IZvEt9Q9sr4p1wud5Fl63yB+7ozoKg/Ox862MJNx0n
u9DO/3Eq4v0e/oOqoErziTVqATeBGsgTGBk4Jbd4bxGFCjsltkU1SlyA2nFyQiQ4Ii9cTgiyyF7T
zbb67ncPMChSkAWfViJAwQVidvMPTuAauefOtuam0DsQGOJuswTHahLaNQeY/UpcsNbZ/AtecrQH
nrpvbgzEbUsf0oQVkFQnWevCaqlihYdMyKCUg4KbkWhxPz0UCCAq1pYSDTpozOHBEKVi58FAS8O5
DEor029FSOFD3EW2IPQtHBYcycskQaQUUH1SW4PTXYFhlVBWbclk1tSGbClqPxhRR+jYaKeE5sfg
YmkMPhYVJTTdoE9kY5CwB1mrRn8gsaDL0l2HEAiqWbZs2UD7ENdr9e1G99i6KSjgTjqQII136Lpn
kmP1tukTtkXM7WW/q6ZVFRmA5kZ5PosJLMkaeCRthHkCeveKwWhfEAl3fgkdo8ZXUCTw2QpRDcIY
2dl7mfhQ7u1KutsGXB56+cRLuSgSvEXkMHKZAlDZRENq3cAZx3zi7X4bCmDJn/Kpg1b1HFkyQIjH
RAFmmNmHfDhA2WV/d7ZnUqOQkesbswp7GIIC/t+UTzE2jmrijtK3hJL3ovKtLnyPBW0+J5JwZAUc
Yo8owVcC98XmzKEY6XWPRN58MJmVsaxrOFMYp4Qgw20NWK/7XuWf40ldmcoe2S7S+qlDxg7VfleT
cJN7YuW4wGDk4vMYKb40ROl1GWAOuUIVnWZyq8Em9LjrYwMG4IgECKMmnR/musnYDfPtmUxhU+Jx
Fw3EgMfeGJttb56Pxyg6vJiEBNnoyCSCmx4QLY4cWZsvsziOxN2wmwjmu3OwQBXMxymFequdt7Iy
kUyEfLfJzLZ+47CXMV4pdDSI5j32lRbO5DVnlKSVu+Vuqi8FYUv2KTioivl/mArWvlytLYVNxD8v
VpYUYAD3Lfc1Dxu6TLe3zZkRYT1Zo34JecZa4vgIOkEIXRtrhQ1pbpjoBfGQ4Lw9oaIuhg4X1sgo
G1YxzbyNvoWvE/A91e3XOeitwe5YUksQwRu3mhHpN1AkC8s2xrlhU1AvI8vi4S2IVStXKjHsjRDY
jtufoa9qXbZL8XaF7WkWP+lI5t6z9lsSLOxFmLCICFBwpWFlsy+y2LZVljjnQQNPYmfzRBRQcl1I
0u7zmAxYoEvmRKzKhL8rQ0TJOein7CQdHRJvCH64vtfgaOQ4299C/+ehMeb1iz1rSl7A3aToxkP3
QFmniY1EhWCBEw/B1N+Vvd3QRgq+4vK2Z/XSWgGoV8cfIdVVDXNolImmOgiKhPx91fae0ykSElgH
lHAAf8g4AEOkOwAgZNRQ2w+XCWY6iTwT6ClKYzGUOZJvcOAd9t3IZzFiBZvjJWeYVawucWLt5OU8
Yi5bpq6d4aiviOpZjX9ddGS5f1yHizSJiEUbbH5MVesPceSXEGlbAn9JKeD4vps2u8UXXrmXU27J
Qozz9+Zd6E8izFy0vsUbgZlLvXfy2GlOcCtsGUtFXr3VFJRH9+sLFgHpzdQnGB2TNsLRgb9LlRt3
jamcDWzzMmBfOYLW02b+pgaX0kHrsEkKAL1/3hMnE8Fh3qotYcGrJrfXuefC604VTYoiN0jyqxSA
QzbK3FT19vffoONhEIiwHOZIUqKY5uI0MSo+d83vqeGPvTEV5TCmv1hXmhJK5iWLF8EyXFmcD97B
+zSnXOuV16U7itobRb5NR4zwKJ3ta1IwgTFKsVpICXmgvxqzbnyOD2qJ7EiMlkE5hEpArSATh0g7
N3IDhNu2L6yusSza5fuNyY7Srud9pKjipJRbUMi2V/MG/TSxmIcqG2IHBElH5AIbpYqpOq6l7v7c
226ga7v6bjlTBIKYHfTEZZ7Cn6n9GsFsr1Mi7/cyEEKRAt+RlM3RpWIGTwHL6ISg/1i6K036vQZZ
IFAUaxznpsnvdbSMWs8FBSFZbIEsgOt+fEa60bjyvCRfj/fRrDezKHgzZSayMRT0JBfntf74gvom
7/bvfD1mIPZJRZ2XiNgi8Pl3pPCOt23lGPfW/i6qeDTF8KFxjACRCD+UByi0l6Oa3KeNSrz5Y1Q3
QBtQD9tX20jTbTDfZg9TqJlnHJFZKA3TH6Futy9ut13TAOWrrQ+YS60KLEaTnDlPWpSr9IyLYBye
tBbTMsRlRbdVblr2vgPIw0abId5aHXm4O68Wl7Q7lmwZ33BSvDnri5Mzzm7g/ein26Kns9K6E2Xq
RBdduCwVIlOokmGrRYGc03QY/xhSIPS45yknwmQKzzKHTv/mp9Fg3lEX1hTgtW3CxjB0GZ7sPxDV
68wzVgqb8iPvrzHNUPcESok3shpoM5/XVwQrD/FSIYv3As8D7xlxP41Ov8CrbFSFsR3WfG8RPkKM
sYnDoiIaVxTdl7oa8EgDcQ+iEsizhkaLZvxQt0C6R7bbADZMEVdKGs/0kNt6zpSGY3xdkJHAW101
bSYQCrorsk06lZF/nT8CHCM7FAOuik80oh8ldUj8nkvYvzd8mmujFOiOzGfwsTFJz7AL5UejZvvo
3CUFZmhH4iNBLFHamD5P8oT+kP/4iA9Fj32fY3hfvhPlEqS2mOfRz/D027BOu0VyDiNqdKPqzs99
Rf1XOwyjjfSW4JP2brWHq78iON2ValZijHI6mdCRJiq9qDkoJOEpexvdMffoznWVOh8pmoQNIY9a
mUyIKZQW7CRW+GOqvsq+bN7AgOLOWZs9pVd0II47lWXHuvEz+uFbNxasBj+yRironZdi3gpCsAiB
UXbtlRiLeFAxe53gLW/R8Y0LpO5KcaFsOhNl4CLHs/RkPNzYA1rXSTtg12UhsnRZDIUCnTEixtgb
4wZaFnggW8BdkpcQ+roQ5JLqXX36RtNPy0I6882OAySWu4SMh/iMTqY9l0PdAEos7ZfSjYDmar/R
5mL/dixaDm7wTsdpgv0cszFt3gRpSiL0NIn/wsN3WwParIG5R/46YWjg67FWZ2o6vM0hyzxvnY37
lGK670QA5c5H3zRG4Nv2NiZ8SWQbAgs5GgNlE7wGsfKIrGq6TgI4HJMdY6EAHf24kQ7SlL/UKlnC
yFXuUPHQd/pNMSpsbi8xc1TeeWUMugg7SZTrIIYtzIxpcoRY8txDzUrpudtinBUhagHs8wpN6+ow
zLbsiZqeBSdxA87xqAibTxjkr2fPfgw8L39A5mQjY3Ka2wpewnnt6hT10dR4i5eALq2YL8ILRggE
GeHu96G29E6rT1KZObrq0ftHvG4rdvc0d+j2Rj/YkjwSOoTkgpxWH8KF0jBP6oeKWL+3vXxAkup4
7PHIX25YJc8zVLlp+/eYEdgut9pJMUKS+X45U6Nn7O2idK9c/IFfMxfjOrGufn+DlRImc1Yq5dOV
Vt/1NQWEITauwzw04suOoCloR7wuSrgiYwkeM8UpL95OJTiSVHCosxHtgU66Tq94DO1ZfPSBnBOV
jy226sxjibUYoSJuwsYwOlyvCYttdbc0PlAYLh38I8nbEOa0AXTNxMkoFI8jLkKzT+df7pv9uJJf
VwuEan10bZIIaw6FaodOQqcNQQ8o9vD7FbIK+r2AOzJZ1fc0+CsorJK0om/F//SYcYUuzi6ae3zI
19nKB5664NGeN0oORTzVmR6kcnvV1F06nFyO2zcVYIxHpnkioIK2GfCDPZA86BlPdHjH8mUsiAVK
urYseN4OvEJmO3rh1D5NH1M8yhXkWRARl9CBM8JquRWznxfopdQ2u2I3HJ2vI9WjnhbOiHG6MHAA
7a2D1SfTiC0Mq4/Ndq/6gaAa7WhxiWCX7LdgaY9G85EtvCvl1Snj3LURtpB5QxJ85SrV9ynOqWBF
WXJVg4r4P/DlRMqyTJ2W5ixVkyRNuYLdcSYvqoO+fgmC2dOi+TzOc1OQmndKmEwZ6+mRD00pfp+t
+TaaDkj/afKvNytnu3wrrS90Ga42yLd9hVTB9CmXBGc2oTS2EIGBfo5zvFpUvyejvmfYyl8jhaR5
yRNV6j5GK4zFY5GSS1b8l+78HxXYVxrjnkZ0OCah5RPCMaSAQQz8EiHKiKTjPJ3lb+Hzie19sjCb
AF0gzWQKokAy1DaRW8tv4bKX0a0kI9EvTTx3pks4+UCc3mqiiVBI/bMHFQBHBBVCGRbrccqNZOgK
N46YxaEOFMoGnQ/u4losdNxY4icb785ckLlBisEpNA8RSLH3sn2zqrtcF0v+TJX0RjcAvinIJfY3
I/95UpgLXAlHS6QlCheLamnLSAOPQ3R3HEZukppNoFDpLyyp1Y/S3fXW8k8KTosMSbycq7djVkKu
I9JEnPCo3+r9lnRRI/efWi6QQvpeQbwPi7ObGzf0ec/8cgm2TXasduufyUTcc1lZpnVWg1izKXh1
3vd3oaTb0C9WuXNMk/Bbb/FJeJcIiZ/hR8Q/2I4yT6r6NwaL1qCSXLyN2GrXuQv5a5w6OuixMTCD
J3QnKAtPpRMP2BNIAOysiPgDqLeE1StXeDFiir+VpDMlIbSfxo453tTP56tJD6v8wmTU8wXzQ/Bz
6qEgaoI6+eh/ugKdP2T1LLc8tb9+1G/A50N42LMraO6LuEn/ggc5GNFPhsIQJZaUrV0ElNd+DAM+
IXkStGm99ujYJWRIt/VL8gDLeYZps1aVcUpkukvbI7/dLuq0qzAhT6vej3ihgLoOYO+vYW0FaQpl
DAVrpHyLyNPl+kJslF9hAh64uWaRfIW6pF7PFAygJv3lO7W6TPJWeoWeioDUhhY/OuicVToXbbvQ
5oMfUz18ubo4ST/StSNiIFTpXk6Z9H2PVGs5VXztomx8sOxi741fWWSpO3QAbgJ19rNF19bjt/kZ
oG4ajJlYBMICp8d3NeIB4NNQmva37tRqDvUEWwb/6arBMKVbkTNN1p1KMbs0aoWWJjpOk3YUrblG
ypcdKBREZYhQEbJij67shCDkRrc7fauCNOG5C28nI63hVBv0fJRctU0hcaGN6OyErQrDt8n2Chuh
3Hiu8RDnIge9jfgtHZAlUBbKWDMavW1rLhqNmUMhqHaaFtEHnMboIv+PnnCCGtPxN5VdDspJt9Ds
V3WTmkzn3NiDWkw8Mci6EzjS10rLlGcumagbQATiaUrg05Ut5Z0CqFBLw80s8CIJdV+XARfPX3wV
eyGk87ATVPYb8IzIlGZ4j4uwVEHdHBa/2F/1qRDXmUN6Ez/Fqy5StrmA9UL5Xqu4EQLKfAsQUaYM
6Kc3AJd1fOcGFkFOR+dYUAjoJXrt140+ljH6lDVDAVvomO/bvrBesmm+RN7W3+Rh1UcbIShXaAoa
azjJqKIxeH0+RzSNoP7TIEZWlqSH2yBqL6oo2DTKpJkuYVj23+h/pkkmSF2yRU31o3h9TMRs6roB
1nY959ofXXoYNF/9gTRl5WSTrfvCoAD61w+PhRgf8OlQF2nZS9RylpObiB+lwBqoEOg4cU2MkeDQ
JkfIfbVTSxB0kC2CBvLx9QoB7NGS3H6Qsb309ajZpRJ6OhUsbYae3CvO7JPRXT4QSuk/N0ycz8pX
yRezV4vUuBA+h3o4vSkIjZ6UJQ7f+XH0EjIMsbEA/NAjgsJVEtD1jf8xheKeBsanbzxgl+cmI9NH
Ke6f9C6CGV3NJRt94IxGRqCuLw7qv8CeZc8MQikCShiH4oVG7b2c92QNWWWS8go09BsbKKl6kSQl
jX0DaAqGbr6tl6Ft3wDDw8hsc6K4oiGeeedtnqIu5R/aMNq/1K5qxVKb+e7kMR0olYnMXpmWlFVc
mDR/80DTVScxGmtxFJn6OLtO/ShYR0IZVN1zgCoSIXzu+HUzCvN/7sFdqimUlULZw0uI/w4hH1ZG
x6eIu/XH88HFcGrxRw/5oyJF6Zu+Z4OxFvNmGzUlfemjfb5SHQ73xW1oSyjvg3WcmRn/FrCWRYN+
ZIUf7+pIqPWvYNz4QNXWgN4CcWYdy9EnwTbRTenVCetVeaPPUv90SjGrCaIRhLgOklm0Sd4H+bzI
rkfLo95RoYNt53+KrOdQ33tO59nCneHYKqcofnyJuupprZlhXTyMbVwoUMAO3nsD4q0i7cziAVdS
rqbnqu6lQ8Gm8VAzKqi3mKjN2ONrWkjo3w9Zdb+ZCI90M5Q7pok/SW5fFygrP+/6TfoZd4d1KgQ9
BA2acU1++nAZYDdpbh2j74T90l70U2fj8+7TQysgQPn+bnCwHOWHRCxUDFjka7Ji4qDsswHbzvhn
L9XxDg6V2aht0bXby2/w7lWNsR+QdUqWPWaqqqWRHRCqaxnxJ1DMq+5zs7c6lauFEMvkpWzygnqN
vhq2b3tGqQWNxZqZQQJuAAimLWt7DXdtJSBIKQbGWBVKkx/x0EkzFOrARLEfTQK8k321MhYecRm3
eUgAXQNiZytfnvJVjgUUyUmZRbZNVfgcRDP5+zZqLg/QTOIfD7Pobgrl6tELXV32xYeFMFviPOz4
4rDB0U2SVL+DaaThk3dyPhkMbWARnDs+mvjK3XxiPNK5yAMEEYyQs4xPK9+jUggGatPEE8CUGTlX
4Lx4iQZ32qZGPBX8WhJu7ZwW7AAWfSXHL5l9BSxfLKeCHOabsV7d6A68Zu2RnLWWtp/K7KecF5LI
J/Q6f1AYqP4Qk63cPKw5PSAGYtuWobhCjqMkFw1vRuynLfb02MYztq6TSELRhRtshgXU/GnNRTYv
Gl+18Xtc0KtZbsUbvtD8P3SlwqoUCfqH9aJZlZHFRiA54jgq6+pK+3vylLnSSsHobYeWDkg2L9qw
fAyUIg78inTBrIBgRYbMSfGyaBFn0JVSY7TyXpJBWqVTOM3Fxfe6URjrqkaxIJbt+BMAGcll1+yB
0DBN8vZ64tInWu8WLovYO9KPpHGPUF/UGgmF58jKOb3q6hZTm/D3OjrVrN9tE7JnBNYiERNVI2cb
vgtGU4/SoThbnGGS3clZRqO8bTT1MVcA9syOQ2sB9+lw6YlylRMli8p2vRMloXk4OZy7pEytvTLr
It+ALQC3qYge3ZBdj/mkZrqbR4zK0g9Xb1lgX9ik58/0bpRSBGVv1EdjF+kjkLHDc9OaC2MwtYZN
mH9aHcFLi4MBmtotQ6E/nDoKDv8Eq9TodYVAx8/6f/pyJXBMP6GrVSlatPF4tCNkh3zKM46wM38/
SGOmM0067acOzxqvEK9UFJcMlVQAKv0gUGi9+a/NUx4gffaNMkpy6dJ4AFzWYC/k1tsmmjD8Dmrl
pXFYWJm5EVVTj7xVkqTnN4VcpYBr94ema1/TFHesQYdKb9WapCxUn0XMEp9SqY5/Yxn2Ebm3tyFa
oZofsGY0uw1Hb3WUUArrOcHhAfDjHr5pR5M7zLhRBm/KG0K9zuzN77fM+5dgPT6lP6h4NaENpo1m
5YVf+CXiFL1e51heq+/A3NtGPr2FIOi8PZShjY+nXkrwjV/RutCH9DCw4xACTXjNyzIzYiusr0OE
uH8f8KPb/kzJ3vTiPGjjwXbsH/ryySc24RBwiF2SRLlV9wpYoJEZ7z8cVdseIeBOWmXnyJ+g5ZuF
VAWWqPDDNXkllZuJfafPSdcPTSsIONgAV+3EDhnF9f5DxoH4PznoFtfoEREG2HQIWIo9cADZWoXP
BZ24Z003neLDL24wIKSccZ7uyAzwDxwRWI1zfN8EUiWoPj8LhTcikzHjvwmGCQGv7rqTjjnt/Mrl
O8V58IILAM2beVHUeoIsf+Px0u4COcJz1Ob8jNYIALv2K1Q0S7n4k3K4rumSvZ+Mqyat4SV9Bvef
fDxXAQFGltXQllW7BlKm5YnKsT6pIB+wHJzvwt5nRRY2mhemCnA59nnqg5mTX2NayUzJ6sU6t1aO
zSljVWOXxQalIoSoEQ1T/ivLLm/n3F6K9MUaoOhvNS4NrhYePXlpGtyJMgWgPwF8o/KUK7VNK0QO
SSKVumSNE1pkmmLuiD8Z5TY0tn9xpLCPgO0l0v20yNqn/NMoJUKxHOBGm4H0q1y+UCHr3DhV7Rjd
f4MhBMeu4ehxHiH2L0mApsn18oQNmqYRth7XR6mae7aIGXDDuWHvWZbpRjG9MgKa7F7zx24VOjJb
fOfV3OTFQ2C1qZ41iuvUx1ybyonlgKdDo7TCOUAkTKGsVdA7lw8/UqdlLLEFZfMKlBQln+o+xijP
SQEltiMGnBG1oM+t2RbxUk42VmwUxlLlmF51nax6qubqy0f6Yh0jWXcNj8X8OUaw775Jy+jt0Emm
ZQZQfmjN923iva+EvOgijtZRBnMxL69g/XGs4zSgJP/fh0ODdpP2LwdNFxgtZol2lAXRd6iHd15v
mZpFG4l1h0DTn2VLMgzgLGFtJ1ksyldnj7hPOU+S3GQOPZUlJr65kVzBmmWTL8wvggEsHKorSowa
2EArf3j6OOy860JutpStppeHgPWDTnkqMurEBBUL4O8w3aKgQS8C2vniHW5UrABAh03woAA7Krpx
bUOc0ZU568U4W/d0DKm9c0ff7U+59MyRItO0kYkRod1lvyG0ie4+0iMssINYv8pThwUMBdZm3RpV
4eem7SFSav0fvQwnn5Y8h5KODZ+/8twXTK5ufvj16ceL/xvd0Yn5F8JREgwxNROM/HtuEtlg1ovP
edIY6ne33amMqd87EZJ3fZgqSfr4itB4/8ur50vOfUqWJ6hXHAS4+so1O3akI/jZNyBq2MEVwwDK
HtrXrRTkGF0+eYtvaXTFsHXjWmJmTKL8fDNmWjzNF7GljtSww8RAnR06175wlxCeiG2zO9XbKS1s
IG+YDL35rkubpyGryibxDOd2PtHgXdaMl0545RZU/7divqSfnei4zPCPmX/270bCHXn+eNZHVPNX
cwkyTd8cZjTiM/mLUs97/8eiIwffJlztebHIT98fgynDwIeUKv4N6OiGPnP/aKFnwYxnyyZG6MHG
WDQgJB8Sqc7Es9bQLheSDle5n7xsSm6+sjssNwhKLGF+mpwlhV+SIxFac1+JUCaq0dIutaEMm54w
tJcxvsQhDtQkyrCj6Z4rRMJx2sTXzVViSLSa9korl1HEIaQ7nJTo84+JmhxLx5gWsUfZTi2vLnKC
mdkbei2yz+w+4PJJPSDYpoYF/AFkIuoSf7mz4VfX7hU0a6rLxozGpRVGiGZobFYdryg0l+o4QTPV
uYgGKpCkf1Ah+8/GEya7H/Pq0YFx1Kxs+q4PqihYd8mDLsJFt3ltp+C6Wx/S1E+MDVkru2HfdlCv
W3dKF6YoOHXf9DRQYEAdRDu0aReqWxkwJWlRPSQ17De56CqyaZ3/k73vI4FiclZ/vVMOtkr8tdbJ
xhQRClT/SuPkeUAH4eHnUOMFxto8reiY/OX6gw124A9FYM6TrLifQgR8sN6FX+SvKqLWbHxLM9/l
IGUTBnrz9KBCEnAQWQ9RyDCz54s34TF48BxFx7c51LkeJ2e1WPvMxToB0fmP/3NOKdtf6i4MYvSZ
HsXangJ7SoiR4A4yN0vD6vwca5kIpZnTKWqPf2lCIHiVGIr/BWs+m/sF9lyKbpUT3/IrfmAeK1zM
3ILOWoVBVf4KYYQ/1FcWCR39zv5Uz/Udg5cSBpPzi+EDDOlF/7mu/FdkrzSH7g34AP82/CExYUHu
vP71TSf+Elx2+pF0N9fjGu5GLkxR0IzqBPKnJN4DsTMu+IlS5E/TAZwGB15+rRHoV8q6kKbl2Eab
vG05RoJaKSG7tw/c9yjHFh3EB7J5QJ4EgfmxOb23tczExFtSoh1drDczrFB+MexwBuB2PLlBGGa3
56xWAMBzlb+J8rP2q8XuvHf/CiVNv3AWqqyc7KbvMcdi/3TgaNZBNzjq5ciC1GUkV2f+Lf1Tuw5+
Fh6Lw9uKU2IERq/tQPTpgkubuMpkV0IvPHG0lM7050Uz1Gr+oiVuAF0m4va6y9rCkXRm2mNSQQxg
kKvc+4PI6YCkEFJuTD4633SjXbKd4gfY3VoV9df3oJZdRH4mEBf5qINKutLqjY0vpkPUxSfB/gSp
+oc7tfEod/1uFu/xADl9ATDpAAHTYhOntTczPI242Xm6MFQSyYQ0WBRTKpuL1kEkGdr+6EgQxZOm
Io4rYCF0/rGr/eWHiSBxwGnR5Y+rThkaQuhbGFlilZ9CqMKFtKwhS2kXjZp+S/fw3y/27cEv9iqx
rNwWaFXQwcDG3Ab53PkoAT12JyAJIDoCnzl26SaaACRdO1+qDUsjSeTUrAs4kNYZF1nlnwAPA68p
X1CVeQs2Y3CoSDV+4U71ec+JVXDNK43jxG1cXVbaEKQrUvLr6G2QixDZJxF9oQ2igUIBr3QEB//y
KbKtENlwyHJV7DwFGiYCArrM6q3MWpSLTN8SPt4QvzKaF1APdUE1jx6BpNKvq8uFnoqcY7gExViB
qx9y0mTHGyY9RtKVtMZpGj1bcw+EAhMRrbJGw6WLcLpfeBym+V/CjJD6rNk4AkAslWqylUwnStLR
eAdvxTCNou6jR8qS+68i5ZsvDN7GIN5KviCl3EvuzM956iXlI1zpI2e+lc3S4S6ydB3+GZ14p3eC
hvdGCCSnGvclsYqBRZ1Z9C6oscDO8oHfATGnv+yUgVK4STkOfYO7U/MSCrmIAH4ezdb1iFBekCuV
245q5Q+/6KxyQbPUrRCtRDRi994qyVgDOFuE8pMfcZPC3IfPBYbtfgR3kNCHH8cLRC7V6nBDluic
POjCokDpRv2pTo6v+cbaYm7LgYVCyOgoicdMhuXWIldwtCe4mvsek72G9eTZcTPYgeWvW0NZiKDX
mCJpQCeU0IEHntyDkvep4LZxpMCVZVNvJbmR70lCylSFS/6lFwxQOvJ6G7zHq1o2hl3oQYdlHoVx
JHHh7F+XXb325tEhexAEegw7mM7uumLaYaAG3sJdA7v0fUqKeMWftCmzT4SZUyaHbTQvD7xau5fD
PeN4n8dRDfGE4N66l25pL/PAZwgqIUoixs8eFyDSdPDZGreRE/qOsnKL4Z7XV+I9f5Gy1qHFD283
j77JpkEPIX+M+dsZmxCSCV9SQPoFF/ffZdmAET4q/SMB/Ro4u/9aeZfEtVHYgMgBVjEn6n5Su56B
nV6Dtf34RYNGd0m83mM8VK/jDVryuzelEycx7BLQaieqMguCi4MSkeFpTWyPgn56AUJkCcYadGPG
BwIXEM5XCl+w/YIkyo1JM6Ul94Lxbk71yJqDNwasE/KXwbTYagAqTZvwYo/wcuXwuAnaH2LKEAoP
gRAmkO3b+/+RTUL5PqOdBCShNp80+SYG/YhmFa2FlSNvDrm4e1UhAVijlFZlZZIicsI9BxSZgq/e
Lwj52c3a40bXhDNQrh8LBLdWZzJL069OxexrZaMk40a/fZSh+HIUOFzb6Go6/+dEdF3YnoVsrbSQ
amjyshS7csEhvt8afHrSt7tGjaWn87EWk4ZLVhidznrmJk2ye3JA/w7Fw5cNa9sQl5EvCakGC6M5
OLeEhpOU7NVOJ9tw4OBkCXj37TEUZku9rEyQqpy1QJTkemMdDgPgx/bUkcN9zYZVL3zuwaukhBFP
seynvd8yG6G4TuRix8/CET5O6mob4Zsrsv/V3uXbG6EZMyoDMrQ8gthTi3tdGpkuA4yq7rme4VBZ
q+L8fAZEqv0nN/Gpm49aFIFJWFpv94p8SQi12/NeGtbsKOn/7Yk2YuoL1rMW4l6leT1uV16XhWaD
3NC0TpiO6k4r6Sr8w2FAq4RdpmfahfyRjGG5d7MiuNecZ3pWD10Ycx1Um/TBmHGWhuAd3SvcBDA1
3X3aXwrUMeBH9bvpK5opO8f1bImW+gWkcsN6WnO7ilCpibpMZ/biKOnWv2B+lhkAtZyoSnUO8tk6
WvdmTwnEySqkBjjxfi+27he5AQ46l7KHfp/zg4fx0CfPPyYsnePPCpFjCw2JiJ7oQnOlXi1E69BB
6plmWLxKBUsY5jpSCuV1rc95DADj0Cf7NahPA41iE+w3OPknYWintu6fTeg6n/UQ5VMa4bHruuR3
JzsjCCsVSuaGvAxJIaHg2ZAUfL7fHJ12m1/JjmrDmA+rlWrr4yzaiy/15RK4xiH+8KJqWuVuQc3L
ZF4Tz6Tq+gAbFGY6jZJW3YgW924kpDtOA7g0vgLyATk03aBfa9artqtAi5Lm7PhVSK48ZSMykQTa
NqVUCV2/WEmg5+jPtpV0cEgnacOapfz65hDW4pt9ZirTyUMwOFbnDoredSpMJGGHcrOig6L7LzUj
T/Hb1bETJuKVNscq1ArwYcU4NODu8cJEgc4K20UA9X/krI//7KU1X+KLzB+y6MNPlkdS450D40yT
1yTlG39ywBHc46UXMe3LG//WEV/k641/K98Gg4WRcisaiACINBqYLO9wyFTUaHFhSz7Ltp5P/F50
yfkYjb2e1evbxvzLPafr6JQe4rZyPuk9sneIYqGgaB88VnpufMLihx5TbnK96IhN96ucyfqe3Zym
93yqBKHviUltsCZpE04WpVUJI2eldrpp039a3hbqIBR1dkJaIvTotV8vZasrd0uSzL49NmIpzTn5
rXLz0QjxtfqENjkJpi/7cmVdLLEdHkecTuhIrYlF0T45EsuILIhVKaw/w3cN5BqlDGav/njMoIFF
HVUUC3UuejPS+zu2Mqcf+wy4//HsF5FQlPOoDu+dK/vdTmI9efKocb6BATDHl5SNLUbpUPpdDKkc
sv+IVV722tEIykHyZT5snMnGzzVYWe6X7PB/t1lGBOvbWWLTor/1r78T20CAs++rcvaf11o1ROeS
pag0jshg7Mc56rq+xG9ssKE9lOF6oKalGlCgcnDMYf2jF2XSqHHhYibF+Lk8Z8Ifd7BjI37GE13M
7zYF1TfGXvxPMPgz2OMZNMihWeMZaIzCoCrE96o/B+ZBkuV7zz8C276K0tGTQewFtfnDUR61HgxQ
CNrPsRlRRbTBs1ptr7VwR/fCf/LkSaP4N8CCIgPijtDEmgnlPbneROEILocVtOFgUCNokhVZNlNC
M1+ZPHWVjFq6ZVrOfU8YURsVnWhh6CQSNAcFBzdDX1MSP/Fa8U3C6S5GsAjyWrMZ/lZgCrFgFVaa
UjCnEx0SJqPPQ1W1AYD3MiwWLo+mvEGLmJClvBd/AdQvGXt3NkIlaTeVMgVUvWtHsgm2NlLTbhMn
zZd0jFmUZJ8lYUUWULN5onbR+Pd6u80XDxIzFoc79mIs0eIWSapEEGFoEQKnMLhV1TzUJvrByZjZ
GLtfRNpVwr4Kfr6lcrK9Yl60L4EizWRSnKa6V9P0ybqsmPP6uFuZ3cTDi6tvidI8FVwNsiGIu1hT
XZ1MBEmbEyLF72uGkEYIKwHEYyIgD+eq2Hdb2OcCMVVQjF7EZhLugNCayaWHC6z8R6vcmhJveR9U
QzatZ6EGbWZMekjnZAZ2FjtY5tEzVF3SpPKkDLiMSNXd4xmwBSgfICv+ISN2sAslwlUjYfjW6Mml
meZbvggC/tkNkHmWB/N35Negufg4+gAiaokYhRPTHFIPKRngE2ac6wBn8B0fW7gr2og2K9e8UJnS
UhGzYaWLNHdiy6nAwamsDd49V2Dm/vIol5bU5JBERmiGq0NIRWnygTpCsxlhsipkgKbbEjvKS/YS
rSw+ymc+ofpkbAPlLiDwe4gsKzscH3cwNaOzHRoJp4c8cEs2AGeCAQhB7UDMg9HUfCe3vDrvmdFt
hRjueJ7EgNkgWQCeUONtjrdeuDv30fZDdHtH7IKD25hV36JyGLU0eaw5J4jLzlH4mGvdEPPQ+lPr
B1h4eb47u+Cg+tAZL/lqyQQecSzQwdnq7k1LEDLs13+IUZYl7njSHJZj4t195Bu5uenGscr+bzbV
APguXk52S9XizRmjLCsUJ2n1OTUhud0IC6A/AQqGJu+uBtoIhGjEzWu6MHD7NfLmXGMf31AIgH3/
3cDdetBouwqgHUD2I4/bH91mRjUOcoB5xqkOBu8pBif15M8HlTEFdQAm6Rsq9JTFHcdesP1oXOax
EviaXWkc4xaaRFKye83jcoUIO9QJ4ST1ftS/RUdl6uiHPwkvvt+O8kVO849vWM3jh0iwH3/weIqM
kxLdRR51ZcaoevunnjNRNwkUFUarlOX//7bSq2WhINNaKa+osnjBNXXi6vUiDA1rzPpFfU3dS6Fs
tdv5LJanvCy5C33nR1wsiCDFqPOxi13ZK1E3KgUMmSl5ryZ3Dz4GmYuSS0+rukArk7rb4OewidIe
kuPtP4UAj473r3NkBFFN4bIDq5/mUom+An+CldoNr0JwyTWayhYpzB5zGHEb9Oq2X34j1mtFpScv
yQvfqLzECKT6RIOffWQTOXtCD+LLBcWyb1z9IGR1YOSxAggd8nqg/PyMQKgqNiw7ISzhcWRO7n8X
zcZ8X9Tlw++6bf2BYMvtimfTglEdWPd903FviqbEm8TSfAeJKgkeg1xJDRkvC3Wt+y/i30a+guoK
xRSvmoIWR5Ct/KPP2b7hhkf/4n8RtoA5bUiYf70S6u36fYGdRjzo3awZShJ5UYs17jM6QQryTTtU
9j0UaYNwaE6bvQkjWfDWrHj0JNFl/+EsBV0bd9sfF/1GiPMSxM7WpbeCMG05e3XFCF9Z/hbYl1jN
azry0pyPwaGG3ZYpqKNpFSRy+GNpktJgu7RyjY8ZD68a9JH2WFxxfjN58WneYEesevegldGfFo/8
1MgeIwg7twd6xTw7Byb7pAiAWTU15Aip4xebMe6QvJziFfwEcDiEm57p/McKprxdK+0Z/9gn/RaA
8ji1XdUVGNEbBR5buLjM5JDXI/WNQDFCv5Rsq2w2fwuT/c5xSZhe07E+i5DC5XUHVKYBT95VKvmK
lO54YMwND/hULwgB5EtX5EWZUR51I+O/Tq7YQGETIjEz0Ks0qrTa6Jn6pDL1OXtY75M8Zsk3wSTc
7K9U0qHURPvOMzjvLdMQ/XF4XYMljZ98oK7nZFXLBatG0HKwARnfurTlLE0Gy6RYz01Qm2o49HWE
vRhfrJczo7Xjkt3LRrZXJ8XsqsyR7c0HHsxwPUu7qEEZA8HL4u++/crchfyda9xdXUe+QwHiVGyA
P3tav4hTQcArxMywvjNzdvqBnHwFCf9I7HDcNsonT1GqISnwveQShhWv51bzrWuT09+9nfZXOC+P
l6NHq2qQkTd5Sm+WT3HKHKHjWVbR5AYsiWzd72X4bjuOnoVvkVgUdbMmmgd4DfeyGYvebvW2Pjs9
OloeSK4lxqz6HyOWpc0RjPsKjfpi8IVk36KIVlHKTEPSsZlhQYq7gv5tf7u5LMT7JXOl1kkdTzbY
cFXilaNeYkvxTUxHjrvzuu5vJ5paN87FVcdERHrxsCH3Ogjh7Mg65RaCw1JVIv9vWWYkBnbG1WD3
cTVyubgImgMWa7UOLfc6ZgiublDbUng+xk9ISBXnhoqBydUUDn2h7h0R4ZYXK8WsJZZ2YvySNzM/
VdCrWejyaS+lOzdiBBgxNmFcGDCwjHqgt99FcFecat5sR+3pQ9z6m+J5tUHDdRFmMJCdv7+eDzJc
q30CWOf5cigU0hDzWntWWOJN/WLMRuQ86sFsyi/slpfZ5qGLYTd00J5lVFD2x34JgBemuLVFR32a
viICWqozzsQFD/GGmkPfvdB1aJ8HVkCiGS19RshL3xeHG1VqwXOm6GcnmGPnzriEH03uSL37QEHn
oM59Cd+9liqFFaAVrqlzBRObtzk84zrjvOmzBMPan4bL3Fd2CuJx6Mdy3aN/A8WJ+NPUx97r6NDH
trlB/jP/iEWaRE06qCsJoUtyTO3nmMWCeyC+ZT7PJdiH5GP9OfXjWzZZ7qC47W6YZKejfPlEl52q
FWopkHl6l3NQV/ZOFr1JsrKhvT7RIygfeOdgtlBb92Jfx1y4oz5LlE458+fWkS3rJD/cgFEWHMx4
/sKveK1ttS9RN5u+azugBs2AUnmF58+oKP7p+VZa1tzZ3DYCooVIKqCyZfYICpIMQ1vBpS6GGOrk
83jFXs/tw/9+a3of8n8Gqac++BXgvPTgYMPri3gmMW19dcQAwB5I3zI/W3aZcb3AFxY3cT2fvxdo
ZvlFEpnrMak1jobplTOH3jui7H38hp2jcQKSAil4F6kWKWHh0aFU3F5jSC0SYKDSMfVZAvWm+yg4
eXnkBlLGRdYoFD10UHA5YL17liQSBBCVlY8vSLtxoSrbvZ+jBuF7OSjstdQBgsR14rJqlmVz56jZ
MjbwIzhw65XjfAjEksgtiBpOuO0ceqHFA87kDrHlkadZWfJEcRTlV5AzTR2KG3KAShxdJLxrjBPU
H30Di+sSdq3l9FW3Cq3daqShUHd7z4QSXuxw9u6yTnvdiVU+WnIdRCzdGec1kDORcuoe3BCU6wuD
4RtTiRaR4ZGdupP6i9qfxfZQaKjBQJDkVGFVWAutjOOFxo1xaxUb/VO052AqhG4DnCX+4a/JIvCV
eQXnvSIePTaz5usygWgztvoKv+nQEFbQZxA/L+EjM5Iffz3v6SNewTAGVgt+YEEYATv6G5ZpOIoT
zH/b5Zm++yhlec6vyu+ax1zCr9aGAOTTM0PwyMIYE2nNVlHJpoGsHlMDDDt3UUJDMgsYjeGppHCx
S07M1zJb2tHN9+hbUFapLe9+FkJYJRAuvAibTk6U0vKwtJ4YkqXtKS1RdMJffZ703SUUoJVYKh+p
m0rimwQZ0FCtXHFf+b/et0hTV9Fnm2oO/j1T4JsthSquD4/FooX3Q7RVLTFTZCZSLILAoknc+Uol
ZAHlF7wu431ICPpwbGdaH8ab+RVOQJEkiYIvNr2TZoodFOQ7RS4Dn6yn0rDS8LwPtv0Y4OKHWa2F
jOUkxRCydzlSjptttUcLeWHqgfmPDiYtNkIAD74HVyPV2xk7BpHO6C8m7yaVOnmkowbqLHBvG1AQ
YezUE1lzYTH9vFGKruDXWEBgloAvljCwORYPwUAAJxDNaTFGPDwc/0pGWARy47srG1aTBK2FiL9b
6Qy5pMUl0DBji7e3Tky49DKVBFMTyj1Gs9VwLZ1AcylvtPA3h+GviHyEZrwPGUPi/XeKrg2yeALA
Wwn21pdZ7F9Jfw+2DEGVq+VhYDZymX8Mu+uThAAXvBGbZylVunxwXMdc+LPDVHrODE/DU9onC790
/3l7QHEg4Vl43YMq+2X/k0g0xfc6LPXDwtPsShflQLi7k1K9CtcdAsD1mZ3QdgWXIEG49oyD5KWd
wL0iq/I8KFTvu6a4W/P2k5J228g/tuxkgQvGls/tKrVIG/8vACfowhh8mg26x4AjeKl2wvy79XqL
DNKT2oJRJOFnhLoUhdsJ3uLszFoGffWsWozaXXJaIhEfy8KnXgTEI03u1d6VspAXMlBoHZyZ/SQC
dMpZj1CGOgtgNjTPKaWo5L04Ula2/0D/DgDcuKnLnI2w+6pJDIJlg3yhfxC5XRahcH8t0RGS7NiT
/32CgqMz1naJovx+/2hBJ57jqOQowz1VCGLRP9jL7kJpYSkls8ofa2eAmtP8Q/531nKYC4sE/1ib
5GC2wbhFatuKn1Z7I8gSbiaSMMWDfCDMhKrTgyDGYVWfh25oRBc1G9BcaxbeoLFzOexfqcF1pJ09
fiQ98WWeQcJ9C7RlG45Qy100aPEoxammePikQ6PjA7dNk+5kYladJsyvvA0jeD4/BVGVKcHYZkIN
5mdYAywRTFTsIQyDnSlk2/QHgnJUCqTMc+xZlaE0B9lk0ZNVLKOytl4VWA25fXcw2tJuzHD+vBjf
WGs1UMCT8QVB5uhEjo8D+Nxy64kIpvnHiuIq74ar9jFuxs0NwSoPKOr9UxfRbVg9DUejanJ0+yXB
T+HDXe/vRL0QBclTEtnkhU+vn7LgsFt2AHA/S8LYEZbF6+dpxSbX4rq2gVff+sXxzzPhx534hN5H
7vhGvEvBRaJofLqeaDvjQ8ApeJrONP9TiHMFJFtlPoyD9YrfNyYj/PUrtYEYsNTezdLOTLy5Mmc0
kkv6l2y6txGEHPScDnJQPTy6+pF34CxfNAtEb3dFXyNARyIDNZWqxcedgaU38bkVtB6NBLXZpDZz
9WPtJ39NluhPLZXS+73YJgXRgVjJv4wsxVdahXioyA/RW70mKVN7muZfMTGYs3BrT3eGl388luH9
VgzudaWLHIP8VSgeSl2a1zZnogj3q3EAK5vhlqcnvLzOeBhQ8YU/54KG411jnh58j/TkxGMFGBLX
+leEXpoF5kszsGccwzZgChfqbLOlhwEKtVWSOZAg5pg5kw9skAYe0yH7Dz3undDcCx/pNi3KlrHm
jw85RwTUbZDEB15CcM9xhCMGNTl92NsZqFwidmZw1bNZW1ntj0hUd3V3eawGp3zjnvPfiAEnS1AR
Udus1OLbR3ryy8lz5rIYN9izfp+VW8mDhGAXD4jAgkiFAsI7Q8x5zWPYKuxrOg2b7BSiMCNHbICb
YIFFlXyaN1fdZBDVZDLNibuv6rTufjMguud5+WeyZNL8cglw+J2Oh5p89c6amE2H4dmBdKA1u3qt
I5iX0Q0FNUfF919G+WFFtar6oKBk+0v/2a40idu1jq88Ph+E/Y0Z14in0D9ipUC1tDpqxC9KZWGj
dVyizDwdlHJPLqqgmMFzWOrxPeoSclSTS7yOL2AOcH9ifYjU+2kkoaxlmGLnd3YFYmE/OXICRA48
rDdsyRy3XEJut/Uw6TYwUqQa6Hf/9Hpr9Ht3CV7xY5wzm+THteDqNnB12Eqvnptlo8rLIBtTV2OV
S36cFcySegDYAVY2XV7/hEyoPdmeSBL7/aAPQxXplVKBY4MIaKcQMWgt/mv3CmqZUvcQykgNgXBX
XsXLZLQTFN7/R8VHfQw0AE1iLRdiX5HPActN1YunGUX9uI9QBk99iWy1ZmxlocU0wc5VVY+ammk/
FW/LRPcCmTmKx8m63ZFxS0r9MP87szW5zBp+goPOyXd8Rg/LNzKYIp9qYndhXn4zOp7DwXy0gu1d
QF6Rl02hyhYH/aV57/xjKIeTaoIfJldXIZ3HV0pXjVFzBUeE1NxRl7OqBu7QTByHy+dFEEEeCVz4
NqC+ZhNNq9llp+Uz6mcBrbN3HsoHT8nhQ/hDbawbqMMKZRe1y6NjHKjoIlxkYCZU4gh4zAR82HMZ
hHuOKBu/PjCUMkSYgJe01vLqcPrYdvRtjHcLK05eYOEEectMq5jXQT7x+d5h8FZr5Vom6ot6UJ3q
z8qqOWgRTcSTf7w7veh5kFvJXF2clWnAfVGTpo8BvgmbRDdZYewON1Rx/1fWcYlrAM2+fcA3/u4S
fLj4RpW17ud2L+3ZTjwjASrt+hKlJJY7ZKgUDHD+qCICE8sZI5yLKQ28/nBsDcrXZatDuE+Nyv3t
hQ58If28HwLCit7qQUmWkpBgtZYOTGdy9RAQTfIUnsT/0+9v3IVPK+4H3szvPYsJhoXIc6kB9aOT
NqKDTv58cXGiviO+uq2DeLHP69ebvnT3+QVqtH+gyyJ1TLDmGUJM25Uh7uYOFWKioUkBhIXhtmfa
M10SRAB3zko2wlhnKRoxC+TwLoyjxLTDjCZb47XVxbqiEwb7ZKbAPLLiSwhALa0rE5KMHgUK5EeB
8F1uV7SXaComtkOIQu/0PhvuzWPLcHN2+qEh8zPspcd9oiwC8o5QpfKnAbZNvgqGf001L4BOwexg
rhAkUc8b6h4U3WEL2o6QaNcdm6Z4UgGq/AENX+gTB+HkiIIMlu59P+JO7yaFI2aIXec+eZh4Dq3F
6CQsHj/uNKHR2lvAogvApbqznMTJM5V3AFrARH/Gw/jQD6FLizt74SdUp9NhGVnmkC7sw5X37ufW
2wW8ImdMTViPDXnQwLbJEeCCLW5oEBg/RmcnaLf4N5+LBkt0XQB0ldgq34duZJVqz6v76rmMsSQX
sx2DUn/ASlyfpWYlWamD0LQaL9ThpuP1145ZR439aEMwPN+uLzuLQ4gMvmy/RK102OA2qT/hzBOv
kOSw8iF4ZpN4tAdyR6k+w2k463ZnHqXtjs+fRRZa5Cqh7ZVWD1v2Dgt3Jfy9BV62FUuI4770vJIo
k05+7UpMcCUbH1+007OGcAM00SP8zgOYGYrgSjkia5275qEOjhCp8TAlccvCYTnLJ3+8I6gw/ud1
rqhPU0H2HgpbQYCFlXL8KycxDiQSCN87pIIlYvuhN9e+ZKWIFkkTFdfSsePQtlQ0fd2MZVyYI+Ld
uy9DLJSjFncxdzkvQiPgVuEFaXn9a3xP8ZN3H7Iql/KO2CPJJJrFZ2Jn1R/Zxhm72iO7Ah6BRrc5
swNE6OyeGeSWfagdASIT/7YZfq2iGZl21I8tQ4en1Q0Aqzw7krPD1KFzOu7FtVLGaYMeQn8Asypf
hF4Y2lCt7Yw8C/ZYADUa7hGXGneCAkVxEMOwtd1ZIGI8OTRekNgCbs//4J3EyS/x79Yjz8/Y/BwK
JcoZL/fQbZEUtPB43vOELTjC0OYqYoaLUU7jJgDGUUcxlKOvcDheFBRc8kLdQWkRROFoPSlv8FXV
dpSj3BEN7Wc8b1hkjAdeNPSgkJ8fznMnBSr87OURJOv+IzL9JJPdKMtc3opyFuWww6f/osQ+5jg9
A+9CDqLFSEs3DsgEBSRdqnIDX8U6P37gcxvF2Mv+LWxQDIu/eAgrrcBBE7HQBgEEUAnnhsjTNswc
GS6iX+imn6RqdqqdrybBxVVL0ClPfMeo5FmEgFj4bDPQkqbh0X4kgb4sQNqyNmcApgwD5iF5i7L8
lmF4Pxas0dASNKsETOTDBA5mMoieAI+pXu5qu9/k2O/6O766gXqooqA7IoQZn5vGySmzRZsUnhlm
pC5v9XApvbIsrhRB15TCnT6oRzsipU4rSiE5ZLtnvYemYPnS/UUeYJbWwDjgzRRBqCBduvKbvyky
6DO/G3zdONrEYCCXw33Ww3dHj6mHw3GTIcLojdArKY+bHvelnES3KWef3KSYn2K2W8QUxPm6ZgJu
tmMSp1t0n3N1hIupDvqEQilF849v04WTH/Z6UXHGmP9X4xo4AUGAoQ+jfj0/P8M6tpg5I7jAHDWH
IC62pyhu/d1GlzkEcrgKHnN2sTID2Ufohmh/J77Lu6iIXbB2IKZ24jQuylCrJviw2F7ozAW6miyt
XuvqqIecezYq/yW6/vr9/dZTgkpGAnxrFQkxAg/3Uzcmo3PnmwdI/qiwhW2fxRaBttSmWGz7yMmx
gdb0VkX4vO6KQTIW/KtypL8aIkk6FBDBV3axsGAHY94CXKytNF9PF0LIOYqKApF7uN2F44xXag/N
1W4kOj9pY/Pim/voLH8GXNYhAojpyl1W76SqvZt75SaWzG0XjQjT+IYAITdNl/9jeQfh4UZSpGy4
fW5iy/gXhzpw90HkhE1OjJpcKuI2um16+YZ6FVigaynTTmVxf/8EX49TkNOua8EtgpJD8icqNHoe
gWWW+AsFdWtz0B247kB2e1xvzZEUK6QsG1F6IjkUlE+8jt4QucEGXGPd081V1RIIiHYk71hNb4j+
WmRiM6aV2MelXI+BvfgR91VKwSrLbrT72JTJdEEwQ7SJ4QEk9MwnJO/Xx4OL7GLwO+Be9zEV+Pog
I44QX4DBx2n/14mx7elGriThaSr1U8vzSuXCf+z6kzo51pOASx3k21W0NFzwgzBAwoQfAuEsThLJ
0V6vwOacbFJcKGXERpDunWWXLyL5HnwA9kUxvnwwNX+vtGp8CLjmkFUlbUrWwaCMFZtYqKaBsWwQ
RdyoKGHSQ1Opt9qAVM6XnYa/H1vrWKHoqbcg8zBVDAZY4//G2vUjzEG6nRb/IHh5kQIvk634Llzj
R1K43QIr2tDRrhSdohYGv6ZylgFnofNUveLcmItZo7VCeF4Bikmkospi7hOw4BvNox1+BfmQg+jl
VftACagDLci33e1/+xB+Jfc71AHdibysnfND5MeIspnFPzVpSv/+PrYS5oVUEM4492NHUwslerRf
Xrg0XUX6AM5k8o4fHL563DED4IYqPf7GIV+aTAb+kBtP+FigDz8I32w+SnYZQni6OLUl+rD2UesF
pNayZh1OAo48v1hlF5in9E+LBAvYfKULaY/hZYBIgc09hWxFxRTpwS9UgEErmF3CNBwfVNPKxrCa
eNDgEkr0cYDtUDYj8ByAzLIL2aOXsLLaSBbBjOUqoXYPqd/4wyzuFieagT5xb5yAcJfeB/OOHK1Y
TMmnvy/WL32RnCmlJXCkh5wAYo8qwcNJbQ04mRgf7h+7bSvBhuOdIm6K03nXeCrR2qfivIFwyYrk
GEtcvGRCNOB+6Lx6Zsa3enYg+OniH9kGjNtqRDgASv6zzGSZHOBriAsVAyYieeYWxrC+RNlJLIS9
zS2n66KZn9K9iotId6X0/cTL1vs2CMfZB0MVkrAuSUcRnTQUJRPjkcELMtyJOQpg+DwfUW8HKA/B
f7tMr9mOFI33zWBai961iPtU6/0ycSF+SRIEhlcgzCpm2n6yAg6OQz96t2VtnbkJPtNsRzRerRIt
Bl64XEcqkx1vQJYo72gs1BmDvZayDYxTTqVDD/hppuKv45Y4ASzOx6n4XSv4fW27p+E2uoNkq04g
Ekh8jlhNEfi9PRwZpkeLX47nFDrRP4X3UzeNdhGoX7Pf/CuwiGwsRqAoitWsUqZbsMgL+lUl7GR/
ftADxct2yby+jMERJ4SePbmXjfdS+gZPdYWVxg+W1ZJ8hVEqvyb/indbFRCdeNYLPwuowip9XF9I
kgVl7yrFDkPU3rM05fMkHROf0aUz+xonpa0jdAHknKf+M5zopTuhgk09shksScemYDjuNIDQg7SE
w9Chp0PXieN2CXu8vXpsmihIHhlksny+O7NpvX2Wl/PYkzRO6bgPR8quu96XAL0rzygPSz+1dWjm
WqtCP9AgSI9f6hXUrgFIbJTFlHNII3fOwHm2VYUaVWpkiwsbuHmGhPurNwlmOhjEj/aodZNEYYda
cEa1NO/Nv1rXHlmupf1ZHq7+g1vFODRIq9IAutPUeQai1MopWPFJ7KIrufLZzSSfgc+jrpEuiODO
Q25u1LDGG6whfLOAotPg2S9B5VRA2/UYnjEPNmaaPxM3T9fXOKw6lPEmR/wkMsze+YoYUogRe4Mx
tKHDVCyckD3ZkJYJQqhlRzpDcix/b43z1kH1sPr0sPbtwlOInI6zL/F/QPZxcq/ogyvVNXwkaGa6
nXTam/2pCqyXxVgGwEqTY80rwja2ePkYnBXbYfetvXvivPGAqByTkJIrGr6WX6KwrHJFFpnJ9Jyc
4OpaZ4t0H2boJk2CnTzIaAjlNY4beVw2eQGDrxmZKke1ALTSzPG5CvQ1BuXGDIpcm1sGrRb3P21W
C9QhdGe6lO4sbFdO8bzLFgMYPwifWfNxrCGenJcmI/jqtKXkgRq3n3dZa0LL6jyF47uqTuuf9hC2
49MhE7BW0MRY2VTLppidsuxYFprYyMxlG7d12A4hdmChaa298XeiPyz7Ttsaz5rNvVB6eZnP7zly
ZTyelicYgthV5oCwOaBB89SQeJJq+jM8MfdyC+a52a5KlfsTezTXf6RiaFkWD930TDAfMmuNH+pK
y7hv5zmEmLelIrtL+ucggbsx4tK0UacuBXrdavZf4fRzydwAyKUXLuDtKtMj5td98u60x4c8o6y8
zdIlmZAbfsv/S3OrZYyDFMzdLY5R4LscI3gTEWZ1Ef+k1Atgh44HFHah5C/sATUxGBUT75mhMCf6
vO1qfIiLvt0nU2UVCP/+yvxLoWiL+PdtNKteOQUEKOOgjU2f6t9HwQFtaOUACzd8eYm23BN1nYlQ
lnngVG4+abny/vHJ66b79PTEIB3k+y3d68J+ipiPi66+ziRCilZe3tMHtpX41kf4lqMM/6WdM9Hs
riz9o56ojwHJDwQXorIinv7/LjiIqYUoq3Fe7wxgRGvKP5ztAnEFvJMUySJUco/4M7HvnXRdiF2D
c00v099/5JjMV2GBYifHPaKCYqKiBW4ORBa8iHOiiaX/28NJbsfgRfxQQeF2W2q3aP8/Dj3PSm5H
NeJsVrtWqX+iKe5xgB3kTt1vyQ4SJMLH2Rrzf7tchc0c9b+7M99ei0rhJJyEsAv2dgGGniUXAybB
LCaQhy+1YSuw2GhiejtEey0SViFrvryZ4tYNt16CUKOjMElvlDrb67JEeWyheiBVpemArDVyWpga
pinDn0dRjCH2if59bQITd+XiqjsBoTOpIa725Z/ZtZ//cn5c0cdg3UTZ2ipKJ5lmEwpw41HCfSK3
BVVy5lc0mXeB0M78sjyC18dHf4LmjtDRwRNz1CkBL9uXVt8ZzGtYSm2lRlQN00aIA8UI3b8KqsRF
e/gtOeNnqr9vqardSJT8LQ4WFqRxLTpwjdoHFJKxbYHpqlAUzlVoERC8vnIKqmdSunNRX5q/EjUV
rvmr6HioXIp2R3uofgEinmbQWrpPu/yn1uZvFKHrHpNVg8jENGgNXgo1KtE63WbI9plKc5dDFHjM
+Y5hNb1m28SSDO1fVuhoc7waRAuz/prk4SAmbVb+GZoSekc4VnDK0ULoIHcO3dzga8su2GbXSLr0
m11Pimrahpw0Hlz9akN1nRH8TT1euIV9lLCvfOk6faKVkHU7vAb7RcI5gKzV10vhZS9CXuUwLc+G
hcMNSDbyYHeYwCXLyUAn0ub78+wcUImsm4IQTBsRl3l/sELLDoPl+TkvQOqrRvVUDHbVA8QsAlD+
i5E+QWXAeIM/gx8kYOmhVaWXVEtyxBzjj7zqlB5B4AdCIFHWEI0D079UMdTx0X8bQW3YfG0f+zMC
irWtWLjBiqBvIos/lhQyiHkVZsv/bNUgqV+I7h/uF7F5mYowldvM/cdQDUySG683BljIjrW+PzcU
na/MyyrrEkmhB/KcCMj5V77NPWz99Fs45iPrxUN6hkZwYAIrdJY/9GCg12deMps85OtR+vYMj18L
VEbaqXxnM09Xw5Gvn+bakczSWvhF9AelJlyrneu2c+YiFseOeVkS5xqvMUThA4yANyfyIv/F1f/L
v2ksVSz5+EpbaTkMmUO8ZZfAMD6lrUqgsNLT1g2zeTK3cTgqbq/aoTo4mn7cQvM9bAqeSL4WzHPv
amndnkTwBOt9ZD1NRvbyBer657ZZSdRIfRFXFG1vGpPgIIXh8VbVFRvGVvBO2JfO28lu8dBQLDyV
bvKqVJRuN8nlwPS8bW409e20HVLFiPxhv8oDDziknRvBqZ2hxFWKesmxB5K3b9IWgbUHZ/irtt6u
XesSa6sBucoqEXGgX3TmS1Yn048+HYIh37SCFXu5/Kz1dUrUpFDzq89ntSofRd5rNuagBhav0bds
+67dZbWfya8BtTWhCndjat09CcPf1E7tSP76xw59MQGTAoMZradVRgqLg4F3uNd9t7rTcdCeYz2A
wig28GKWfCWM8Zn+NhqAOonDYtJ3U8y8+jmSL6C8oMY8fHWnkPV0vU1SUJm9N6UBKKgTSwjrTxQf
BzDcjfon0qWpKJufGqi7C5zx+2U8mxZ/SUYCo+Kjtusro0bFqIxs3yJnXOb+uLkTodUWWhOnErrr
Mfk/TcXmuL66d4VemjQ5QSd5JApWSxCVYvmvFQGEN4fzEhvZ3hbOa0Wjp+auCC3ZSNn00nNJa8Bl
U975bVGXco3h+7uv0yyUXAFhc/BDK9k6oy8IiKiXhJOy5KPzhPjhNwtxatBhX5myNTSY1+q9G1cM
yKx9g7Q4SFnAZrjJ6LszgK/+A37xxPgBAEkzjnlWcTrqcue7+rhM9YZN9W0GfVUfjG8dJ2CF1TEm
qTyRLusetBpoWOndE2STmvKNSLFxHQT+c5O3fudzmjnsFFZ36coDyg4RkYUfA7KSudW3Z1h2Mniq
ZHRVwVd2q6uzfCZpayIqT3Ys8cI+BBs1U3TlhRLZnHiBzA2CqOBGsC6mLPWEUN38RYNvb623Ofmf
lVKKffMm493kDTPPhi9FDLrI7o+fi7Kw9yMM6Lfjf5jaJZEDnlmI3PI5tGUziIJd/5BXquuYcUZk
EQUpBwqLVXHrYCnwjB44XjIClMO1lK6/ojxXyVEgCem4GKUb/OTxpxKB9HyHwU883f8Peoy/oC/+
PpSb32H1KkkcLTHs9cnWRXUc283fUnDXh5TYd37qdk//tSb39Z/JXc++A2AyrePFD/Ax9EE7Kq3h
+FGyQdwrs8TygUepDm7qG2AtANz9RHoXyFTq8jD+N4z3O+b6sC9so+FiqZ7C7cNYtygdS7f5Y8Ln
RJk5tYwbFak+0Gtx7wEaWUz3qp9AW6e+W/GU6xlE9olQAtQmxUrqS5miMj+rsT2vMKZIlQXOPou4
o5Z3saSCZ2EnW09bdRmditkX6a1tMdR2ErlNOjki6lZMI5HHyiQCumMCxai+D+Urnf+0XB9/b2ba
q3x8GhAoeR1UlgUPL7m6CdqPQUprY6a+7j4Z0t1r6aJoF3sSUE0vNvt+QWpyEqwfYf7trDNWLIeH
9/FWWFwzji2ph2ayZrndIdpU3bdRxFxp7Hk9mg6XOw7y3gH12cvXTkinPmi/LaextKW36YKaG6Z5
sJch9bl/RMBzuJxGCfSw35Ps4QvycOLEjNtrOSE+gspeQoyCefZcBe2fnaDqVySbSpxxzdJSg9lZ
GoR+GT2GIoF4adSQnH55MY/O5zoEIODatuD2vq0wI3bI4XAEgK9SIFTBOj1/Wh+deUmK1syCggRs
v3nQufb2/xGKga3RYSJQlrgMrZmMzDWo7csGRTW3rsM+t7VTozwtJ6PKI7Qp7VrCXUTEUb7sy5+E
gphPA7NfFsa/a7edFmU5TRl7bVevva5kqKEj7QVrlo8gfbl78VcKMy4UJ9VUxjTnxYzqN2cwGF/F
xS3/iefX8HS8IB4Dvr0pAiPX/XZQ4zRZge0ZpnjyxSJ8O2hrjI4hG50PzrbI03fRZG49IUuRjWTf
SH4rQjcGNhe4X1l3XiLa+TomxljSXwSg3vaBBU+Qpa28gHMIbD9hXVlSExm69KNY6JrHfd4FRFIa
w6j7aMuN6RirEBsf6DdIjCgfYtWNIvjnP3L4M8pVcVQZ8ofzT8tgmXvWyhHJoxxYFfXeC6QW1bNE
xG0woPCQemwlJpwGZQVp7+mxkSlCDz/QW7bCvl6JmUA4YCgyp41RpgLuITkwZc9D1QnihqdkZUYH
lL9qE75EImhdNY7+YZBaMUcXMIZwOb81A0Nnfan94oEcXdGdBgQjzvC0Viir0Sk0+/887d/N5i8c
fa27mSEnaWnszayz7UFpOk8mZg0wfoGzPBMs0BQMG+Fmjm4eFOBvaHouDL/xjpxh2+RzTwo1GUyq
fHV2f/g4GXTEtN/VeZ4ggKWMMSDs5AWWRiFBlj+3Cd003x/TtN7uGHY3Y1sqAiFaw+Di8V7WySFu
r1LMa1IGerZLvVuMz1MJT2Lb77aKscGzmfAEE3uf6VJpW7EhmJUGggLfRfNC8WYSJhJYYLFqNtt8
eO1Qb+6L963XM9jbkFZnXk5dmK5Zw2N7NucpC4Uhtt9SHmidgGXw6td9id9qpzkSf8TFdf8Zjur1
WWGLIffRFTs/0eEVKVOHfI6L/bjqkS78GdJpttovh6+3PuLuS22Bm6a+eXmqc2Q4ZzsZ9p7O2owB
P+U7x6ClzIRu3aCMrxiIeJCzON67NmY9V9T7ne5HFxyRap5jQKXNspiARyAGjf86qYUJCfspsreF
ZZ3qx/SCM/MsraqpIkW5iCK7SkviEsTDLXb/yFSJxrDnnTeMpVdn4Y2nM6O0fqnJnG1skGNyJKhQ
PWhcNB5VPWmPrcSFNmoxfpReTHvHJhqJj2H4prEN0TJCk4/pAI1KdCmNVOAANCZ5NnuBwvvSDibl
eP7UBztc3W2vsujuMdep65wMrjpapRgwM2mN0uyc+pZS4NcCXce7HWWOBzZGvE1h0qPijVM2ChOi
43plJ8UvGYcI6T7oGWhHTrf/MWrjHcpj81kfMngJdEAJulv06S5CBP0OolJUst4UxwMzGNGtf6Ok
eHwZp2kPXfXWtDQiS7UsiKuDP0JqdpoXgla2nGqJXXkrCyV4GZ+CFn53rS5Lao4AOC3Mla5+XluT
9E7VJaIPtrE/06fPsHQdUhbUlnLct/FPFraX5I5T1c5EavpHRH35vSEuRwnZuekk3ef+gkOxQLLo
lYxME4ROINbjAbm+ibgde9qq18SVD0Sy9ORY8cuCmS+SFqXynbwGjJ5pn8QmEN7RmwEY17j/KOM2
+OitIKIrqSlngFq6yyc/yybbHMaZ/5nncH+D/GLtjee40v7K5f0Frtl9zR+hvXc7I6RFF6nnsJAT
ybweFnKHHnj2c1RtiuaeLhikUrudrHUJu+xrmKy4it5iornhfJAuYcIZsGdIfeclVH/EwEZ4fO8N
RSf7LxiSbXXej9OFQme0reCrllgqml+CJbiclNj3xeT9OLDVFWnJAtgrvKjyBGRoonTO18aNhPKO
sJZCowGtEczku/jfu5bICvpZ+Ewk5MiyeyCFEMlsvowHiUoQOZl19O6sRmPIe2RiQrIN5IZ7z538
zesPY51InFvtwZQ9QvEIDa7UCHYJjFE5YUaUXRhILAB4UAtkFDNsmF/NpvLlGnwvfNEXgy42i64w
wSU47fxmq86E2HVSE945hNFAfuv4tPjEfytf4ysuG3anyi2vr8HNqjSMhLM4avVkUBi8E03UoJFp
Kb8Rj8s/Te3E/h60mfNBzUU9+ZNDefVFc0jrfs8D6jd83qri/A/YlNds0D+JTwxmBr5vqVnyJO/1
PIpGcFwjdwnIReCvhtkLL7xF6ltWkB5tYaBIIRXvzswfnIxFsrSkkX/991KyJ9JTQrRTVSYuV+0F
PEOHct3J/fxiNgItoGdtPQ3qYz8oDugHsQG74gZitsF6ybtV9VdUj+vLIf9NPrPN7XfChgGeZf8p
KpSTVqqRpoCQDVwkTFTNn7BYrdNQvhSHns5TyGpA+KcHJg1NaEnk4l3hy2qjE8RLj3iNrjqeVXm1
hUZVTWjWQlVYwgpyD6eHtcm4GQ+KJjmOLq2/mYHVp5owjQ5RMsjQCCRNNwdV1vQM38O8atGYRrNr
mQJZP/dG6QJJRUS/TGxm307TvMG14iq4y2f0PtGs56JbnBwTR11nSJtwNVBDnCvabMYyohLJn9vD
Ut3ozt70v426JJogfTbgVCvVNobbekKmV4sUphsbn+1l+6VcBUULKAwksRrtMKxzzRIEscL824zk
mj3bbo8ul/wQ79gHAKyRxZAQoGM/GeO8VgoPsH9PP1gEnlQVYzu0QYjWeQYpUpJv5g7je2LbAvHP
3EomRVre69fgNllQFf+mosYzKc5xroTbI7ts7SFNhEr1yjYbEAHkrp46PiWJS4RS5CtsKaI/IKEB
YP5oD5IX6t45P0FEVNV97hjKjtVzP60LxWP5/QW8Y/INjmA3rAF/g/KDTFUwB4q3UIZRzhIXXnLt
ClTBOt/MkeX9N0K7Ykt9bFXYD8mW9T1Ol8hDNCJ9WfG6zS/a2XMfwIjT96d5Whk7BY/F1iTXkd1i
4U3z3E8EFjV+9U9sbyHhdUVS6cHzJ8A/ZyPmFcENdFGkfPlLhQh8RxH6fnLT0L4TPmPRrfoVlc6s
yyS0zaCm8bvXVU3O2Q7E6e4TAwLSSH6HouncK5GDKmFAgJjP+dXPup8eMH6lbWTMyyEQts3kbGH5
xvfhYU05zxkRk8s3zAkcyrNRsHaZDirzHcoPPzGOJ8+oTpP/VA6zQia/slItZO3BOCstv1g+vbQY
goNy1PiRWtooXcZAeZ5FxrChx0/OnsY5/qFtMuvh6jII4leX4RxQ/rIG0Xy/aTLcfJfgMtDHY26Y
5mDiV2oOyQEdhNm3GHNPYgQd8RGD0Lk+CbDMpDl/EDhuTfbDzSFzM5qIoNUwSsE5F5SFgGFUv+jn
d1QgPxcPHC9fvG9bCnSNr6SAulZJNqdiR0tni5HPxivSk8E7IJNHa9tFtkbkEGdpYcTs1qd/BwUh
Q1RhIPQc8VnIGPw1E3a8/kOYSWK3l5zkH5hAd1KJ4BLhGSEhT9+WO8D6isArUixiFDKsWNTeRvFl
VUx8Cvp0c+xWwR4mLV+WGuEJGF6CE6wvM4loQ6a/Xj5g22q2bWTSnOJopJbfy6Sq3t4kEjYpsk0g
DeT8FkzpJuaMRjJq9TDu1hwvAvQtSB8raWv3iytpjuCKGsPksp68fTaBNmbKwCCS/+d0s6sOHuJm
tQqfg4LhKOupKwZE/1TnSHoJFXhyc61iomQRbjhrbgP5S8BLPXMmG5CspLhWC+jOqtT/DAsqklOs
5U6iD6u0qump0mLVFgofkkL2PA0ktDAWg2M3sYp5T3ot7T01TXiAKfkQJJah5hhRx5kN/m2FkO8N
N4LGecmxB2M3IoSZRcgNfWSoXJgI5+PVbr62PpQ8MVkBCd9szW3WnGQB0h9ZKE9elsc0HgCyWyEC
KwcS1T4eKDgQIIRgywSPQ9Gl9djgd4RCDNuO04JsxLF7nlpfPIDjE/rDohHdbAujVDFLQ4g5azkF
5DhOEsflmpiU3/O3lUbLbUcT0WeGT8ji/IjQl4q/amEW2xKWpn59tiUkZp7Sd8csTVA+KruafF2r
P3SPGgdhvQbPzHri0DWU98qqNSohuhCRY1KgYGf5QOM4R7gpRkm7NrDG6T3QmQKYw8KdjhH4qNlS
fb+Hx2uydixHELYfm3gIkNCK0g6up3uxf/WmQg7jHx2rZR950yn8lrh0GEftJo8G14kCA3OhbyQq
TfOsERYPuXkr3dB5BaN7YO0UFcIMHB/3/3ud1PoC65+G1oltEnrNY+D6zfTR/CWNBVqJNV3aavzw
yDy629dUyRbwvsvT8ayCZSRDlZ2h1+SXvXsk1sc3vZvrYZCAjCrG9+xXuNmhWu5ISk5Da34vXJg3
o3SvWfXgDYTkWcp5/uYZzpOfkvNPUhnlPvEgVrttWf4u36Fq6ljZeCiI0pLj0lCstsZI4ux16lEt
3uQ4utZZS/yYujbU6Hm3p/69GOr2Ga11WJn44/rNz37WlU1M5LwqX7tmGtZvtejYZuJIUEdTRu2J
+XCzVpualTsTKNp1lQrFSOe5lhJYkfC9rNUYmLeGyaNcHhSRDESjkhCJI/C/IkQ2qfbEYxk6v2Fc
xYSReVJrQCJx+0k7jijw7ng/pzxGn/9DfUaJgkhym26eRs2scpG3FVRW6TpwCnBXo6PBAk8I9GQR
/hOOrz/tLSTKrKaWV87rIemHQDBVUuKThMcaksNooG9/KJ28UUfV5zNwgHv8S5/XMJszF71GSeKo
uYpJFKWgACg9LHGPlx3zIHIx5aHlR7MUGS8e7OAkIfkhq18f8ARjPVgzuXf54KKw8p5BsOgZeNiX
7FqxfQ4c7q3+jf1hvw04ya9O65Ylc/aCxOH8HRO0sfvCKpKdoCz7q+DgCam9y7NDSzeIoUeKVM7o
AnR7UPWS9d6kQ/IjErk9L4d6Y4Musl/HfuG0zNNKYY0omEyk8uCYwpbmfaqG6EGdSIwoNe6DLWuS
keHVLESaUMvDrsaf16MwbJ3iFgwWCs2xqwNoKGKi95U7dovIBso+iI730sBAJMearMZrSlXt4kx4
J8340ESctjaQzKy2x/eMnduyJcFa+dhTlZ5TVe5FX1Fd17koSmPNPaAxLdxwsrQvYVbGfEFoJ24q
Q2RY3QvhmlvfmGj4nccqBfy4ca3lJd0ZG1NwePebY86nvCLtlKXqcPPS5NJDQi1bxajItKe7/H/2
l08+mWxqwO3mfArezfcx2nqXiOBIdVNr+KNicdZ23aaJbr9Bl43E15vVq+CFZpG90tHouKJtfyFx
rCdvrWixNXz0hmIQXSGpBE+rgJaiRZDYiT+VNPbEKQZmWL2/M/BF8jpEn4YWjKPLutFcUaEDPWVH
swyd9MBNMWLEzgd4VHCYluzPzGwdoUuvxcUlihSLHCa+pwpuFjcheo0tgslrU8dSU2M7hlzALFt8
EdvQuv0jlkt6uoI913PM3b0NtQyuA8Gu1uunni7K60xbvftEXFpRtpJx+p3cwCljVZEpLijf6V8C
YICT6JH4gcjh22o8+ZlwWhmTvhTwvZqgyIpQIvoaV1cY0Kjj1Qgamtbkj3FamE67BDUD9YVsq3Ra
j/HkK4FHYGHvJ3kTt71CcUSYbWYpIbqRZIAwKCOYdJ2rRd9yJIeo3QerNKEMYODpNUMFnK86r1d2
XPRSkBNcbI9+IOg92L2KQbL1CQnCeO8K9p1tNfuDy/2MsXuYvOIjzipbOoZQa0fgGttkMchcXboJ
EkL3zj+87TPeh1BkKl1LmAN4OzzuJQL7RklKk8IISwQzTZRckipsStCCbJkRjkq1IOBoa7sNDOdU
rtJVIOoV1niWI0i6WKRCAOYgY+VamDKsBTbSc+FAjGEPPtQaubkxjCUOCSKhlNTXugHNAvxwN4vr
PLuUA89WnUeUKCcpEx088VsBmtIgV7X5ABaxEiGs+wx0h8uFpMFuKJ8BC1jDXFKxuO9Ac43X+sjd
7+tjWiUy5HLhy8jrtm/k5P+51yv2+ikzESzIcTNCaadNrGbgSFtqXxSQBkixtMsRU3pKbSOMtdvc
mSl0o8e5KkHT5njbQymIpoqIRcK4xcdBa6MN1vQcwXB99u8bipIDzvNBJeFmtNv/2QcspXnXPFV9
bezCwt5oR4K4UYU4gb7Qu3OwdzMe5ERyq3q2+UEqf3JTqjQex8xnW//ichhD+n+Ia5w8HwWzgofc
pwoiZTnGZmOhPcnGLXHC5rl7KzjhGABmuFRsHLFQAqmj+LTTO1fZqxBQJAypYjbOhg4Kv4JVinaq
uSgta3kqMR5Zwur7Julquxc4W1qZA5yF63bfl32Q7xxUfGcTwOKkCs0QDcQV+bdd6m/rn9X3WtNh
bVJoU3YqNABOH1QtYfha25+sluEiv0gDSK+rfMjUySWtnihiUUlgVGbtrv3cHMN9xgflIT/+Yla8
7UUvc/74cpfBWWQ00qdCjfhTLOFhI5Ad9zHfquCWPMYKb363M4FYoHJOVRPglmuE9pgRngj82Jba
73F6AzZSPFB1dzxWAmug0WuMWNfFRyg9xbIZJabiExgjp47Io0A3HCs9lgVYKf+l38rqeCYUaFpf
h7Yk6ng1PwiRcpzU4kRq7YiBOghv7BXuVCW8aUaipyioKebFJSJ4V3txSPAiyBnSlztAQJR/We3I
5JVfKRdqAytr4R/dSZIgHuEGZYOb6cRI0iFB2+bxSgniyHkyiRP2xHF+Ulx9QP1mnI+LXK+oyH+p
eUqksT3TBWBp8qX8Z9QJGd9bNIN2q6Er10wuPDTdv4KGBE1KBAhr6ZkQGEliyChjwlgkEesjxQr/
vSvh64j7PHzoW7elvTHnsLS3+ceu0A2T7fE2zzj/p7qN6zSIsvxmiHsBBfL2tvOsqsZ4gB4EIgzf
myHeLbMFI4ULU1fS63iDyuuwsHVOnqv+pcg3ehy4Yy2jgDME2cfTup34OpKWuwN7j8MbArUmxC4w
eKcna86cm9GX7bdnSMlItL0qdcCrYK18yyXEsBJRw3VWchaHmePVFx7dMcibWPPNv13ZW+6vZJD+
raWFfneP2TwJBth/VwmchpOuzTeu8P8ARtkfEx9yPa9t0ktXyPOjuY+eVEwjEuRNpkWiGYOR23HQ
cqc9QET47iB+2B/tStQschvSbV8qg0YN0Y5iEoGamKgbOeqIvsaIKDdbuIrFXaNFPvk6gsVsYSeb
kP8AkH8f4UrhgbglhopXpixnbzSHL+kAOFV7rdWSRo7xJlbrPrA1y13bVoUKKO1zEWiFDEHlPpmv
h/94PvwhO9pFFQ1tqJ3qJ1muRJksnlSnNx5EsZBywVE8GkXIGvj9Mt7o1cTnEaHFFi0WM3jWtYBx
M/9MJoiWX5maNIePwKCDG3Rkxw+ql5Iay0OeatLVq+hkmM+7Tz2VT7/dZ6nhyQ7VY6Sp+rjwTY3h
LNd2WAOVZIiUTfNC3+FHmfSQIuz4/kVjv9S986y4goCEgsA/audIal6JOZDgbmv0h1OfN+++pV5x
CcUx3UEmM7TMbugHWsE2jywvtJAlG7cI7/8dio8t4tcQjQsfsTxMUFdoXJXWwSgN2SFUcocdxzHf
rtK/VsiizqOa68MeSwrMkscCanlEijpn2atEE1XuKATIBUxSgT/N6794NDhbLDGYu8FRvT609ebs
evgo5QhpZ7pZpHvceMMqISkw+cEj9TfpMSe0i6TZ9CEAA4ie12+JPi+4YGARp5nJhTMwjQQy8K8D
CQ1gxlliYuM1QraEU0tVhKotlGz+Jz08sazMVzOaYsvHAh4+dUIBeMIKNaeAiSs8V+tFJomsHa2X
jrjQC4nZVdLq3F4C0PQLhTu8Jecn0yKvZpz8CYfFYCWFCT/StEcJNmtStmuBmCzVGRXPYoY+bXaU
8ZlPL7e/ViSSnp8i8yS0dkqrWk5ei2y1DcJYc4Jf5sEyaIplGYRkDVanVoGu2snezPs8rdqmdU/2
OphSnwEVlnTfHltx6kX5GazTsvYOZunjqzsI+uOonZvYay9MYWAcb8yiaJnrKFTZsRn/gXf2S9qE
TxTkJVhsVzlYya2P0bpwiLHLXEytVvYMEUYpHJ5TVwNgON3gG5pF+lP0D/EHJpb3K8WH8Ce7OuIb
Fv1ywdrkBQeNxZzLPdMNW2yz1JaFuG2j+eVDQbtFwIqXunjPZ1FG32AGXifIz621vOs/Z21xK9yi
GBwe02tHhNg5Gx1krtCv8ctbsTflIzU7tYA4WZeYFasQOqHCbWGBemTs6OxElsgmXNYx2/3JsfW0
gwMqHgLIMrmjVCAOd/j4c5eUqUDRZLytMWXAss2NJ4SqYhxDQrEKvjtv325/PoRk2JO2A2aJjHV/
eckSxxpzQIWgy+cBtj7reK8DYllsjYUgFbd9+1aqeB7i2qOmIHdb88L36olO/sD4N9mEIp4/f4cr
HKkrwWJ0yCXhpM7/Sf5mPMsnr7XSoaZ6UYJpUoeObHL+mJ6pSWY7o+dXU6G9qfGdV/5hHBR4pdFL
AQolBBxIj+4r/QmEhWpiwysu3M3alXtIlSSbBnk+xbWM53fYu79n769NsrDwofheX7vF0fQpx3gw
mLN/Z00kUOcmRcvb+otdx6XsjoMoJVL2+BzWZrr33LNwG7ZjHnK545K7jP+rPUO5pKVxefDUX+xt
CCV5u31U6KuUZBMT7XGnFdow7fvbe9wtANJSWvtOMLmCfHhwU0rB1EULDv3V5bnw7RUUSO5zg/tv
SxlyZ8cSm7l8aycNCFrBCunupSID3tLazhFXhfZHbCoDSt8QLiXSI0524pX2VJ+hEbPfhkTFIfng
CNBLivtz96lw8B6777P51mIXqOjazRiCYkJD/AG3HqIc52JiBQBqDjItrhbPtdA8YMQk8RJzo1gR
HT1fnJFIEpO7DuPhnLIaF759F6rcngPe7NRkvVE9wATI4dGcmq88rL/EYfPgZQbGzBTbqx0VeEa9
zEbR6Ld/bGAiKRt0LVf8qxZFmTfbR0Sx/vYkhxW4Yo0OlWToVxi0NEr8+Py8MaHgdvN2Ww+0GyhK
PO4hqmEUeSNXawXf8ws08fvR1Md098SksU8mJXN2bx8VOfSdAoQmZyk5omMDo3b8650CmnbCT4lm
MwZjFPjdIp9CX14LPKWrIdNz15sj0w9+RCF1KjyYe99r7P6xLa0VRw4bPRpDyfinQshuHi7gzwaz
6aCfMNfK4UlftwdLZqEvfpV/FRCpuqZMAz8At5yxmm6Y+VcYzxSjq2wgsvfN4IWyCOiCLWf2zEG3
t+NAu9VTxn1QEhLjlSDdJVW5KJF0dNzf3Lt6ywCivF3dL83Ghsuiddn/4a7+CHpv3FW0EQvahDpF
fvKcjLaTMycmL75P6dnhZF5JYHgg5wJ/s/WBkQatmXkxEsRNiLWR/stJ7W+xWgrmjUpUupX2oILw
SZIBHJU0lfC4XtdyRBUROiMELGaoQn6vGygoGQLzMHfiw8cba4HRuof+WdyXZzdLTNMYgx1BwzI6
I73T1IW7yCO9/nAtgoNdmdx3s8ylUwFwIksVgXVvtTkexnB/w9TIFaVwdHEZqUEmpOS0yulVXLdc
p64NbwXKI2b9tZ4SdtJO00H5AEB0A0Z8HglFHU23gYS+pT/e/p//EHaBJLA6KeimB+fU8LOCnFYY
g9iFUjZffi5Jpss606cO30V0LaYYfRtvFF3PQxoWbcIdoyE0y1uyYx/UF+KwLolGtkyud0tt9sYq
Qfz1RpE+aBYnpgg2zgSAnaeja+Vpw8lm7RCngwVXr+J3nf/I1cm229pckeTA6KEvcHOLGy7V3isl
bN1AARt7pWzx3pFtgmwZswUcpLxj2/2bTxXxaccJCAwBxOs6QlDsfIjvt0FYtdcVQ0QSXatJa3TW
qKkYPPh66xjzyhv0l3AOONRRuPcy+lKCRyDbWInH24TN20YSZZN4yR8XzEpkk8phhNWRu4b0nBMk
bZ4lRNdhlGVlxz5+Py08ZSQgLKEBtaV4DtqNhkE//T5VcXwTeApVIfJPLNJxDpWEJ212NFCo3mNo
Khc3DbBBeUmugCnrPigM8KoPV3P77abKOXwpHmnJ0jqsNDVs4c8wAnuqHmoMCJNCW2aw7d5Madjj
xC9TvaZvt7hDvTe2UXZYhefLOH3QuQLSOKs0yM1/Zo2eC4J7zDvW5H+hFQk84/ujfrSjxC4IHW8z
ncxA5lQiLyYhNl5rRj0iIHeylNEA+wSdZkIOfri3xGxMILvm3VO6WmZNw2ngFmxeTxaIk/W50J2n
AYl2bgA5Mb0ruJ7ERNeYriWHN7XBhYw9tA1JOlItgxk49f2m+wqfPQ/xS7zPrzIFV0KLrEhqBTAE
B8qPtNAu6+eouqcAlREQYivixc8/vwxgJoI1UtW765cP8Wk6OI2se+YEIJGD3lfu6CRn394qRKTo
96bkmQHukWkQ6WtC/K/TMrCJqZYrE7ZrLJcY569xxbbrCH1MpR4pIW6rv8Nx/2FEUXYjuY/2y66N
TSqE8tkUpJnLb+rLJFKHnk0Zi0hjN52VEBiCxLPNccRhyQ2unPsITjOittAaId85Dqp/ppc5rRO+
GVkeL4gfEz6xFQdh8tovmD+ZFaqPxUCO29nN35bKBpJYIeW8Oz/YeB/3r99VXsXajtHbKgRrUfFR
pc09tTrHvqkfEjfzLkXjmsZ3Un+zllRsBiTsRs4bp69sCIr0EQ19FtCrb78HeiSvIakhXQgQmp75
NYyCdYuB/K1okAxv5coEsEmMvig7JBpfDdDV6+payi8iIA79zqaAZxK+rNWTxlNA5p7Xa9cpVZXb
FTcLjOStOD74nDd4EtiRBDlCGWHCI/TzymF9xLyX8/oijfl+QhZ0AdaTFR1dmqfN7EbvJCHS6kTt
S8Iy1x12DF+7vTyftQ20RvjsARwQfDKMO4a6lrHWPobBOwfcSFNmf+Qp7ZDaqbk1ectwFf7J2Zxf
UrcIIHYRRiGQUWQUvkI01fYo8r51YEnbJ2mHNcCA0RIqIN6UIw4PY/DIVOKmKFNwUPFfcZxi9y69
QjwwzToO/hsy25Td1Wg1IbcwzOjBZ2mXGHx8X8ZqeZtQQQVEuFtfMtRK1A/8VZWoFQUH65As8Z3r
sc4/INJSiKyz0S1//AYnQakvbJ1k+nSylQoJGPKvSiIUaHktOS29fqWzavScFndcrSugOshyP8Fy
C4R5MQywlUBT51JLdWZX0mt0uRrVPPCjbE974t4bNZfu0gniwGdkLlTIa4kl2DnG6BIi6ujpcclt
lzaxaok6Pz5nqj8Nq4QwFwGc8t7M6gnqG5o4uXF4dCWjABFpVRKS5YvGaZTqSaENDOAk8vwTpbeN
naVXla0GRARK4NlXuvgFk1koB+CwpsSIHumz7eP/O4uamkk3HzEh9fdNZlLtBkFwfYu8uxDr4Prt
s0D9+DLHPQoPT2GaSnL7mKxkVFClpRdOsUucrRFpf25c6xuaDJj9eDZd20r4CStxqf2llrpAQAf8
J9llysq9T4iti1kRLsZKr518CPxEPUpDNwH5i26k5aNSchE9GIZmzm6gmS2asK6M/lbcRXqMesCv
PmIXl6Pjq3IlV4kbecW7DL8ExF63uBIw+F86EA5r9xd6szXPX4A8cDyQPc+WNZAl9u8GGH7Qf+Or
n3zEsuii5rvtr1kdvSQKH+c1yIT83srZg3Qm2+pTgOekuJc/DFet2VKDd/BQf3cddlWVvMf+gkKx
UWPCoIsidm5BvQi/tiola0iaEX3GEOVd2q+9f7HLMHSxzPX/+J6FtidoCJXahvJhlspyyihQPcPl
w3EgJHe6KTM+VAt1cGGEYEu7no2aAzSFniuoFE2jFa0+tcVG+OcvzFayGFFU9EGL0IOC9mP2ulRa
YvUl7fIBfTUpnpc4lOglHlaOMvT7zUDqHojZuQQSUvuX2two9IIftsYXAVbcBKjTRtOD7MzP9K/z
OZ36LPiyDS98xmauvXS8QtZFRlaG2i8oYlF3PRIIG3xYIX7TNRl0eXwdmOoEUaPxSVlPia4MWvwB
jDIXPYjhrhhzRn0nGgWiyjMIlhA3fDEpa90FaGQ5AsG3j5dxnT0VW1wXayiqiZiNmapzEqenOhCS
2LxjrF0HRYCEr8hfb3Ztj3i2uKlN+PFjCOj9Jq4N70piEmHjj3ewR9NpnLniNHXe0FYWogOCqgXb
GaqxUevTFpwVxkwRse8GAdOrBTYqkCmPKkri6Zd4vFpdOclciVZPAFXmCGJVledqgdLn6QrfV57U
HA1yrxfra1nWxOpoXBbj1vh2C3oR0B5U1jPqusg7pfAPFO1dPuvfl7J7YG8n0XzJ4qbcoBrJUXQH
+KopTqbzv/vukByP6XJ21DmK4J5ctzFeIF/I+06pP4wsN+sYpxakxA8ykXuJABk/yoI9OwoQu51L
dUgmk2kVIlUVCkBSSFFPgDN1/yNomQY7XwUChabKcP1y5GNWiCOqQ5XblSwSYVS6vCgNbZIYwxUi
Ix/fbg2OaR/mZKrCg+P9KiQpoTrRuFVok9G2Z/ts8X/Sl1WqKNocSENHnkXTv64Co9NU/SeLAAJL
UrtcmxRSgvsiVb3ADg8uvx7USkcWdVyvPAqKz62JHZBw9t2p0Yi5QTnr5papTFT/6pbhuLjcihWA
Xye0kguwzUbbyBan1mVGdrXJwzAIpOMWBz+FLDhx5WWPRJ4t8QZDJpfZyEsUxDKBEVZBqpE0hmlP
eHr0w8Pi4FyprsEoa8X0typQXiL3fnvtI94APGCcwWzl4E5/ctcKb5R18VKYz6J71l5kMqq8mjqC
mJgesKQW0ZH5Nkr0F+ZECVGgEYXjTA8bu9AGM3GUcswSshw9C3NFNaa0eF0ycvhIx3r0o2lPflGU
vSVd3ROzNXZxnhu0/uAayodQrFloISVM7pLI8tZZlOcb0nlJclKAoJo/RwsGzNjjf7NhEiraoJzg
OqBsI2oBF9qTfzpYN9nnjMsdtkvyLumRLc2jtaUQaGsxULUs+LF/4NXIpS032mcXWZDDPELd/FHJ
c6yCWzh5nC7Noy4d97C6RB4is39FpmHNjckPG7hLvq0/4tkzg3B8yXtzFI99x2klR47PQHzM4oMp
SbS2oKJcjpjuc2VhL32vovUbMacAOPLJtCypj6IDfEcGaoFZUYhAkwGl5HKZEhXmFLYUiMHprVAx
uy3YH33Tv3cBWFU1zfJKFRlrX+cnd/KRiSjfofDCRbeIxOj0WfRORADqjgh6qJtvAszt1x7283ck
CP8MQSV3NqysebCVVV5ZQ8TF9O3oKiRteOINAsSeTZd+mN9pSUnIlQkZaTR4rmcf5MQMsnELmUTL
IqPknbjdDpZwYJXRiAxt7YNVDJDDZ7ha5UsQUcdtt7VC1ovdEK7sMdElbBbOFu+X0GeAAAl2jqtP
euNnRDCrq9+8ofmrlNlZdtRGtelIl13f5xcUQiqo9WVtkc7/j11eVmabshQ7IJ5NGYUofVP9wAZT
WILWnMTKbgmMTC0rSGDEToNDypwQFTSc9vUTHBV8A7vfZxGEilwmJ03Tq/TUw8BCCrWN+qkt4mVN
mLBhQwUosaV2miX2sxMAKFVIgGr1IO0fqHBk7KvHAOQy+OffEgL0wiHiUZS8JazCDNBxm3gelVZv
su2mU7QFVFdfpDsGSFLYPZr8Cd5LWEfHsrPwVdGCDueMlUaTC8a7CHircppRTHL3i0n1c6OmDFry
Ewtj0U0m9WqrgQBnbf1WgJKXpGehfNah5E8y0qBOQZw1QNkRy2hA7QMQVHJe7S3M581IG30F6Wh3
zLPZSvRm3iDSw35f0awhILUNqNIvL3FbK9q1rS73pABOfTUAnP5QvDNLSKJwdAkgZeZOVDqGofFV
ZLsXcVbvX+1V5wYVDHbldEYMHjyGS13R6oGHyGURH6lUTaJsG/vkW9ehckCC7hsjWpqcizkqhZq3
3gfL2ufFvgXPW4if3WRD/mxHTTxUxvZrJJD6jdA9ER6Jw8qewZZDPeECqazWU8pBwDpBvymAj+hh
XcXRu+YCdyqy0Pyz2vjBAm3WWWKsrMOpI+3G/vKvWmB6woil7KIhYo/w/eDKjjRHyub67AWk+NCo
kO+K5Xgdf+SqEJNRdfvtdRAV/GRc0ynhrsDiK0i/N27vLnjEWOJiCIqs5SZSUBabmL9KzUkEs1AS
+2GNfMV/8D2AJLR+3LBeuDvXP7tc6FQ/N5/hQ/NSayYxJ0pTX3t3Ex84pwFT8nBnyxDnA/6AhxSM
LJOEP23Cm26CTzp23Hz3Rjx66gfsVAan7dFJHcYPoq2QjxlZl1JhGIKDuvLqk1YAWNzB/EV4tv0Z
xZVjsPeeagWIipm2k7K4R08hbPz5VnYnvjnxD3z2ct0Ns37yk4/xm8Gyy0EOZealjePr/VtQwHaq
3mRpEcJQbqPttNHejp5S/tUuKLs66zq3c0dKqws/4336gaAIvjuUb+fdwMcmLsP8EtBMLKAwBal3
GA39xr3O/buMUsDNWe0YFgbOM/6nvnUtXhQ4VGjC1sNP2eF6dX3QMH7TAddFJu8hVCkHIKgCHZ7a
6z72+4PEU6saeH4IMq3lM5iCOEh7OW6FUDt197rWt6aSe6xuoO8cgjwchzjfaqApu6LqcWqLeGwN
QEPwtuhbU2edwSR1cQTKCStujhgZvx9yMb83SH8l55Oj+dsSQEptSZie8DDME5YsYPgKEKXZ2iez
q4RKUNayhGDaGFhSZJjHQO6u4O8Ffqq5ssxRPWGcGo9RgFjAVWWseBqqtofi+tjND7LeA+Z9bMBh
eVWHFbuQmky8A2It4t/8w0Ub8m07A51why82FYAgTS8Gf5D0TP/1rY0gvlrVUOiUoIq9z0wPeiHc
Ee/7I4e+je0Y3pbb+zgvxDOWBr71hxKZua3J8EaqOU7ZWHiuqu/zy53639KDLMqghcTdOd4vRrp3
Eg3sDucdyXbGyASmTZpJVhiMKvhI0+3qgd4f9TJ0vaO0jwCUJYouN6+H2jSqdWDvFRsaueoc5h95
vVY3Ugf4Bw9SjLoE7nZ+WPLsG3cM9gPl7vqNiBo/cPD7j5bjfsgNm2eL9eBvdIehenBMQ8VLvtzN
qRgggzHy3C+JHTng6cS70nkXQu99rkaPQ78mrs6HvvGiIDQj2XuoM9lroyQVe0gtvNZYbA6CKuHm
ysylKSAaIIEgwtQI92EOoLbibZSa2n6U87ixoMNPiU94R9R/2FhU+nqMMfj4r2cnd2BiuZmX0HFY
TbyeY7mRL0wZT3V95UKnebSfASHUVJbNjNFbEtBdCCmbfErPtDWnlbA7/BYFbVdgxfJw4019v4aP
XFLUGRd6f3KMZF9WLgOLONmYB2Bmcv5vhujPuqG4i187l3n5vg+KI9TrHjhROsmDvF81JIbFGdPK
Ijasce2KJfcfXrvgxjSIzyQMNSaFQ3Kov4GvSQVcA9IwYRsZdTGKR4ph0D/JQpYRDhEGIGKcz6kk
X/wuauIcmmH9kG3/PxarmrR6yx/28gP6kx/JVgJ4U+cIYWIi3OM8NdMAF71DLjtNb1MhrFDiazCi
0c7tIFIuryh9BUQHvvDJ5nYYuFUo1iVrQKwrfzo8Jv/4BqKczMZEESre+cqO6gMbmrtmtHaEii4t
LxXAaQ9jO9K0p6QtqCZVMFPMHfXv4GavyOxFFNuxb2juuF9GNmYgNyMZhmOkDztPU2kbJmpGVNtW
VcuCC4y4nwrbBkIQJS7Qn8s/Diy6fhytCnqp9WZoIggBQH5R5hb9sVITZrBG9HpD5IX5NOIePBZs
baiCWQVm/AI0pjhCq50hTM+yBi6TxrgdtXtvXcgjKg3lGBVgq5qwJvtGauoArP/0IimJj2obw0Hn
873H+5cnTlrXe/fdjBaCfPGGuEP5j7jmP3wwlRP1kZ+hPnW2MjAChEyic26EpGTlVT78EGzbjVd+
A/z47nyhRnFib8hZuShEiZm7i1uIr3beCnFckDrjGX/dVN3yB2UuWotRNMbByfjoxgHvTBw4zuoH
dcn5PJvk2YpfDdI191cn4u39MQp0lat6+LFASo/I4DAjgk1rgtfgH+TlxyFn1SVM06y0R9Uv67ph
Km2esVrGRnaAnaSh9dkFK338J/S1uGdVQAPOkTqSMgw+DuLCckXuYSAY1e0IQZ0O8u6a1GpXNuHy
7prRcEo7LtcOAa1FLLfJHN9gHqQ9+/718VRs/hzw9msUN1M7QSqmJoJ6vL37XqavvLIZHiLs3obo
xuLuRtJ3Qxkrf59nQW+Wu5NtqbDKHXyKPSJaeliIUJM0HUSh4Dn8M8hqiBhn0ud4Wp7s0m1kMxw+
YZU02xInE/3cYw7YNKkRpvhVq/jQKV/xb7cospm+wGu/qtK25CHqkcoKtOGjhOLqJOkQJ77gFcci
ITOqDEeQnFaqDcboXzQ5dxAor0NzjgrCa0NHHQ8qgRanl8mmDfnGv88IVw1wZpSJIoyaMnQII+uF
yvMrLq6oKThTpU9xAUayd06bV2/JG4Qt/ZPfwP4yMZi+UXCJ9vF/SwR+fEYPyJ1UBhpxZYLye6KN
iEYVg4t78HXSrLD8VtFVtpba11qp0RnGhZOFKrqXi5kdEmzkxH3sJZHgoLXhVKNWcMa6zDGcOWi2
vndgtvZolhduj/MIcoKxJl5iE7ZzagDflBCsg3Km3t760k0GsxPadgh6PjgWHMCWaHKJKf9Y8X9i
h1Zizhfl0rmN2l54IgqFYoWbYt16MK3gZMy1QqmxU6eD9BPs0wGOxMkUcOG2piDGE8G/cNG3BTwf
QqADAYYGXmatRpDwMxVH++3DTUxvVwnyQYo7/9iC0bcJj1nD3FvjlWX0ZkBCChWk96eJzcA8bJy1
ApjiMU16agi+HvwghJOZzbxQGYK5TJFo4pf8LKmzLegs0DfMFPFepZCzwiY24xdGkjapZBivbU56
rKLKBE/ZHuQ2RR56gkoDJmdEhPGVOLraAe5TdDg5hU8LML6dtxc6tRj2JXFAeM33LX5AGHUZkTli
VFdBBVAV1HzME8gfoH/SmcdUppeqGur28R694x9wUYOqbDHFOtSrx8aTaW1jD8MHk1oElrDiisLp
iccNXTukg8jR7zJKCTzGLaztV2ZaBJjyAmGo1AVkBGhzIzW9Bv0BY35TTVAFrJrnxtXQt4ZZBcmA
jS+1478rJ4d3lyr3JGNRHndEUoaTUc3IVtWg03k6a62TNUWD0SnUbsBJQuDLwJMJ2gW7hb3QKj4A
gs9d6KXbYFuk/LoCGvTO8yTfOuBNQZEXOu9z+9J4yaduEzaFCY1RzmhhUkkPBigP8NoLFRqnQ1+g
Am+HOhV2wOY/L+mZP7JJ8DjtS2V0KTfipfB5lFG33DJIWt1QbHw9kEiY+NsnoT9wpv1fMVJUXerq
aVbjHjV9D7nQ+T7YiDDdD8+CD1wUcx3U52WECYY+7HunR7Vldv2rlMU1piYplnidX4SQLALaNTUX
YqR+sPc2qn61+nVtuqLtPG2Sj1j2KUGce5mDHEIBlbeVDWLe+pLLkTuj28hkI2FivGZWjEqWVCA3
LHbK7Js2kovHVIYEKsq2MC1smVLZjedaP8LPLU9NzdEn5RejOI2/FpeUuU+yuT3bcE91YZMd14XC
RJWsnIRZG5F1hMw8AY80pAYhSsKmnlnZxoMZv07bDbb59R75IVhqIfd0A1wsQgUEwSAe8l1otkAb
mop11fPJRY/0+l/t+nDmnRI486+df6apABgJhxBQIM9Her39Zw7benb6odxKs5HL2wNWoxF7/9VN
bnEBkz8H2LIouosBWbWDQyNcqp++SfzLHaO+TgX2cnnMrUDI+KotWJZWqpDKnvCHENTatR8FXvZT
3N+hdr3aJsLJ5c6GiaCrg5sSIe62rgwhVigOXVk+iTSjxREDQ429knTCsYzDZ2ykZjGZK1KC6W64
7/KeKKvb23uN5o6wEmqgiVCaBX2uI9ArRk514k6W90Cotw/Tj2kZY0+GDXGxAyFRf69lzbTVEiFw
8yTFEBtLAqFF8VBjMrKhkxCXXVe/ScOIK2LArqXVr8x1h7IXXrcCluo3NHxI8RM9pFTS1dV5C5wA
T1mefCQCWOOBDEpYyxtwqIx9U4g5Z77qBfiYUdDRg9LWpqdNJUzcSwbCBDBNbMbF86ZF6ytb0ARw
GV2APRWrg9fEZvW2Ikzu8NjK5tFtOrC1w3+jMWMR3aLeG5A7uy1cdnekk3diwi2xxLF/rLd1o1gg
sUHviBqf+802OZLq5HPlXEdBMW3u7Hsa9XrmSEKwH3guuoosJTCeu6N55Jpy4dKHfGR9WXt9EISn
Ykt48oN1U+BeNnpNVd7au7oeJWnEcKNhAmpiHi9HkKGDchB1dKlpRhFG5sLCTiYF9XtXGXHu2DhO
auf/Y2GI+L2hjRaGyTS7WS9x5XdTtBtdxxDw56/e5I2SWwUqCf8JfoPCfO6RsXPDfoNSlfrdOb9T
QZyaUmtGcbwXbdNkVlcBt+n0rGc6/kKzYYaLiszws1uvl/GQhEossXAfigQjZKQc3j21mKLAVjt+
odnv7Yd4gSGwq5wIoGbYSKiA+b7sMk9tfDuSkN1muufSZcF3CuvbKI7YOBMaxNmaYhClTMadl+xM
yZZx9dPQXNCmKyWpGCBzAAfoSvIiuFQduKaZ7wWNEvDYLXSxSDePn7dRbXjoTXx09b5OCj2IsTHy
KByQ1A9wzkkikDtpsb6TkLUoZZLgPFyOqb9BWVHQoGCu6cwpyh0hHmrCVa3UOuFi3K3bD0CRUSUu
ei2k1dWMzkxbeIoAJWh5hP5JaIW94wBongUdTH4aDgxGyK91eA0KuOxLiTDG0AISD/KCjEL15jyl
rKMYpDooMH9w+GQBcrWVal/b+ydwN4leiaAM/4Dv7A0Tckfvj7QFKf4/aeZgQ+sYwAEFp18YrnRk
r9fw3T4T7yKHgdQ6zw7rHJ8IBetcgOZAqbIIhVRIdPO/iuRwF75yQ1erhXyWJIIJXBwWMfWt9WUR
zq99xJC6Uu7FgUxO83g10xvzxqimG1Zkv6bwRLZewh+dzntky5Rm+288wHqzRbNBcu6i2YsdBYE8
owLNT/41AHk2HdT9mk7WMdYMHPulaE8BCdR62126+1NtjGVAGEuThBNLgUsXHEDr+Fk9Aazwe+GH
ppNmd80ktXpdx457c+dgzicUDITzkSkFkXr+gbsqQIfmnNZoBXC95v2pKLkSkozDwz9XS21XRJBw
qxRM0croX9bvo+gG1DHfanJkdJH/bANjeK+ZJYMt6xDkyvhpErF8bOM0YrktpPJSs5QSlG02GsbW
LQ1WCRYQVmG4rL/fVXedSsbUXJBCi0ENVBlA45f8JAoNnQskH0+V4Xktd9gmyEEj5LoWJx63mU88
vgKKBt8FN+OBBPJH/V+gs7/Z538scORSH0KiR6yG1AgrxU5xPO6Y0yi81WPegiuEbknOcc9h6aQj
kRvfMRbzTlSVFjLY7545aZcVohsyTWcKRCTyO+EKwg9DrrlvW0DHqV0PWZxwOO/hkSmO0KIEIbsz
BrjBJuTvKICHgazQEYYlmW2+uukGBV2CLagr0HAi5HHBuAhEF2u12TjJgS0ghWUaaLwXbDgE3FXK
7XgzceXvXcCPY9IUMSBbyjQBfUxqI+TtuiM4rWiHaNZojm9Z/W2OZZX9PTEr0UdYYo4pQ99bJm4N
MPWge1p83RQYBMoA5tVWVdIao1ahPzpSGS4KuDzTRpfMyDAZ2Yi7XS/bFmZAACR76nPXhdzz0umj
Ak7jwUBrbbg3XSMDBXtE2M0P/Rg1JB3lGAyKnCHS5YcHL86zRYMxqQKdBkgUx4y8f5tB0GO4ZcWN
dgLXXnq1vJXRIc5RYCLPzxr2IuJZEwr9gqSFcWvHmgXCywnK+HdFlKHYrmWQ+BbWorvd79n+oh3a
j1gNB6mLFLgKjYAxC268UWM5qM6122dZ4bVlaxF6cRC43XzCy6npq1d7Avn8+mXguyBCQsLlvQ/b
Pr3YikBgalfpRTx+NFtKltl68G9yp3kRc5tMRUPAZ/fxlKQbQqFsQwhNuvYeL/9t6jp1PWxcSe3u
CRET5n8lecSQYtgGj6Y+o8iBwDOr+TN6KGjfJk/yyrkDVAw1NvvvTC8WP0buR1vZxrYEjDznMGZb
3LAAlQvyvQtDAzgyjwNl63F6WZu3VIB9fr57EYMk00pIbNkZZl3FZ6o3qjc43zZRQDOdM4MFUqjr
PJ3AQX5xjR3rOqTPAuWb6+WY/9a8Gc42iARor5i4cQ3t+1EjH/+6M0LwqYkoGFD9Ikf6xAXGlqR0
Fm5QkRKIrXEmxfbq2TihpK2jGTupizCozUnkCvl0ApbAxpSir71FBjuKJWJLxk2on+N6ChzdKVEU
0YA4n0JRlaLA0qa85M33SbYcbcp28QLM3l9ltgCT4QrELKQMLogSU0jWS/+LF4T0nbuE3Tt0dGJl
V24WOCLsmIf/feUb84w/PPIEG2WyKluW7X8ntrC2PPwUofLgzt5N2iqejj5c4vev7dIcx2/J1Q7s
jqsH6OWQ7+7toSHIm41d2XN+Nh+0/ikN4Bo1c+0+MWp/Db/KK+rawjI6rrXVdi2XKdp2u1bUIAPO
4PXPIk7wM16MYIZyO0NX1BRGNm6KmxJeJSrA7wKUWiteYDGZnKnxWa/iui8teJKw+mjKbyLQ4Vu/
0N0NhSwzBFmBDnJHJO83F04DxsKHQeIaK5KinEtBI49q5HXvHrGOTazM6S505orXqxx/DbKE1Amu
Te8GoE/+ZstfzYiSaLJOR88g76c7NGr3dN4pPfNkuZZIdhhu9EfgplSjnptTY+TF9/mFFsXwTChV
pI12rCK2BGP7Ta8C93yXtS7Lvzu4uGrSSS5exG3lrifcL+Fh1hRHCWuUgTQ/dGxgt378U+mnix7P
Shpraxzv150bMYYw5RZPkk0Mw0gJdxCu0deM4JarGiL5wEmBESTLjqLB7Rz36scQjlaFo70cWsJu
a8UhUan3VHLTGD6X9Irk4vKfl9r1IYjmHXy5o5sTbAhiFAhLpeGB9wgrorWFUueJuMvARQnG8LS+
uSap/1bNitU3BVshvcWr7VsHOV9AJIX2X2JA3xSieiEXWPtIArFWEmx7lqI1PVNPsV6zyDM0b+HO
osUs3JF2wGLQeeEPJB8e2yK41F1cSM/LH/+cUzWWuMETGbhfAIGtu4ZTUkXBu68uXofqxPQaoe/n
ZqUJC0SCD1H4sns82Z4WP/woUu8eUZpIVaRXHgbk3JuG86mMiMnVztrjIPT3xKwiTfwmrVZaXXr/
ZQMP6GtVNbpgLyguBl/3CRp9FJn7G+tXNXcAm0MRzMmlSTm1FuCefZAFTatYf4L0Z2bGRQTA3BqI
fcN0HftoTeFhYftKS7mCf7GgppNFMQ5lkoHbVFAFLcMsMDONA0kRXpJRxvEUooIVzSqL6Fp3Pxt3
3Xz9Y0OTxXY7FEAd0HjHMiNJvu4BzTLg6Nk+97FvoUnhd3N3T2GAq7BlgBgKYSjPKH3hiHpCxwZj
xWyWyyjS869Yfycsd8cQIT0ITpAswXuxtC8hY4a/NU6T240f5bUPY5ITXfct9PrNVKaB1UwaH51Q
7ZrPfHOvqIjf18ugZD9b91shybIjxfy1Wk3IPPrGF3YtKRrl+6xbhz3IjcgM02Od7pxdkFdkYu1G
uDNATiCX/E1pDz42fNJx7nP+7vfN56ICqdAWwXyfLcOCveaJRVUoQAMRewQVYUR3I8LmoS0NhFGM
lnBKQuVSdYKwg2O06gKK4pNRUeRagGnNpaPTlBC99L4leUHy/bsH2qzsW4x10uM6ES3HTnxIucro
XnT4OhIwNS2wkgn1g0449VkkvfO6B44Hmvzj1zGXlHOh7oIjgVteTPBTF8ZM3w5BisUoySPY6sc4
xB9ssXag2RzastNj9ieFX7u7cgPkhkiZmqKptMuYzldQSEqO5fh3pR8wAJd/hs/jzp+LAluac2Ko
/yVmR3V5oh3oeTFkBzMz3EARnwzFRQAWoBc6Tbh21Ttd4hbCt+FFUqVKnDpDX1xniUCY9eR5VzAD
GSpFcNRBZ0HIiyKzxmVUOv6tagzVxO4HY2DpHvLpbDTA8AG/pqQrg/55/NgisIJV1xf7u+AD/z+r
XUuZfJ2UQQpdJUSHqu9CZNUHeyy37yhrs0ePglrqo0hQOrRPHNjJg7nET9dm9PkVEENRuZ+s8Vtq
w7jSsRA2RtAKbQeYyeRsdG2n4phEbtA1Z0cHqf1RaI1K/BKJu+50M/Ow8jZIjjHhg5dgni8M1J97
GYywnNDEKcPt4h0kH/l4MXC9VfODQJh3NKS+HOCHWa6a4uKi0TqNpthcRVvAYReiR3DBtaK3QSS6
pJLKyWfSHA/v18qkn10QaGfIizxZfXEQ/2NL6ZeV4TqaBsJY8G2suMVJAv9ZllSdcUIb+VX8U0XX
ofwbQsUAjANl1xMD3FHRdNQz1pwLMh7bZXexMZuK7fJRZ7AOrrdUbn6Ht3pPfqD4IO+sH/9ZHkOX
pVjMxM7p7bPDb5l2smQB7epm/iQTPADVx+DzBTqm9XKIjzH2YOlYI28xtGy0MeKAAHGQsi1KJHBP
cP8P4sFrl+iTEvJLRdalDNGmgLsjAVuNYZzsJQrSAnlehVHk04JpM4tEfJiW27d85MY2DlfBtxtd
JWiCBnne4xl+UjxvBm8gyVV9wgHR5NGKQa4IX0FhITMTkTQZrUr4xG/YX9JTq8E7IakSauNdVYZp
HFTdBiJoXfYhs8rwhDeujdY3i1kq+gTC5oKZKwQMGPnxlGMHhjnfxZYwFQA7v3HDD/eV2BQlEvVC
cFjkIW3W7JkTRTbul3CKUUhxL25ERZVvUtHJbWk4ituEO1J7Ry18hBeMXy2alHpNtEvi/1VxaAt4
0dKBH/EpG1LSwp0yXPCE5VCdg6tFM2s/7W5GfXwcpxvrPBg9tbPlq0exw6Qf3MqKmjbGpRgAj4Lj
GVnu4oF8A4/72+PSJVGDLdWKdDBPueNUWWXCfGFFWpbZ6SLC1Q8n7XAIO4vaAlSjCGx15sHZVHeW
GIra4hCj/2nTE0oqAo/5ih9/GfuTBJdfbcLPQNzR6474O42FQ0AKKRK7u9IcUzOi37PmyYQEst2V
53z2M8Nt60tMQ6Y7noCbB5nxB0HOBcuP1h1JlYLOFoCoJFJa9+pfQKi9dkFauBKHFF5fUypx63nK
YRU5CviKNAzpo0kWe56ShyR3mSjjwcK7gf8oBz9kBdqKireIRURI+UG5LIwPYuNgwOKC3lRt4/EA
86eYxym4kSc6WUA1ulCCN6VwLwn6UuhJshaeB92kfS2qCZyskO6bTUGt6xQHb/2rSWHEB0tH9TCE
d5GAd8pKX+WV7ZmAHGNLbLtE92DUTc+w8qA0GYi5Kw3VfHyoqv9Qgzop6kSwUoeRO0cOjBG90XTN
k3QBQtM8rCfBDEEeFiTCIguRdAeqUsWBxoe1hJg3TbHd5NkqTacPZ+JhvAcPn9ocQbl/7a/fNP3w
Ww8UD9DgpE1YzjunOfcdBdxEvZU1YoDGRKQaPQUXEBCTaiAgLu3ux8ZATR62FLJsC9Uxj1PVUfLO
qSeTsjsJDOYK7prQq82el3eR4JjYEM+6ddJW+AOdPoKwrX3cMnLK4kwdEKovu/JHtPIGY3c9YzcU
HyAXhmRxeLKV8QwAlUL95/Jt/qqqMtSlBMvYI+144VoZLxaiVW1r2Ktil/TMmOznG0ulep47z12k
5OHJpCZadDILky4wNtx14BN/C60I5E1rGmjcgs1WmkkTPDrut2si8ZmwprZDUfG/i3AT2noXjf5/
N7rsrn7BUCCy1OyjRUcISFmgp0enggf4NoeY7vFlw3NJ0T5Q9BZKr7z/LLqE8Kqdtp90whaHfMKG
8IOqxg+LW6BccXuYTrtVGmZUWfeqy3ZRMH7BiEZnHHA5Zm6c2aKeH89auiR4vEjT4dSkRYvs/OEb
zNF1p4Z2WXb7GLOHBzKvVkSkVD5GM8LUMVQ2n0+fEYR7omuGOvsLR7jUaomYuxdfGMmhGBuLilz+
5zkNdURPsD/cHG7C896HsD306lvvu4DtPOFo9jTJNU//qpfE5TXQwMqo8CaM+p/eaH+FnLXl8a/c
yEO97EhuTPFuO5gVG5xWnUi/4N97MZFcGDmdCH7l/00p5nQwEWqyjnQcuJPmgXNj0I5zALBBj6nE
uxtxgeseNqvTDdLG51dVgdtA9t1s+BHsx83xy9/OglaH7isMRdl9rti0qKhjEJUo0Docu7qlXD7/
b3YHuu0VFf72+/ptKVW9Bj+RAFRD30HhzOrHX5R9ZctDOfM6IhsrOa6LrBpBnBfUvkU5yVkght8P
7FgrYFXNBTUixVHCt3CbS5RdBi/5+IuN9dNYOyWWrJwxVVkKyYAt51R+lBH7YUnCB3onsNVqmoqy
0/BmIE5Cdvz2gYt1thkqKNlIqsu2fzMefmMqTlliZwMwX8OVNHWg9RoxTvgBW7tlO0NbBe9h1kUJ
jghTIcyTSUkyvvrI0BxVgIXaM6eE8QndtOcpkR22e90rLDFkKivxzMm3r14mSenhitNVMNoxDJ+n
0wkYW6OUD/H6+DjN5ZZilI3tehtqbM8wyMbTIpm4g9+Ca60Tbas/zKIsOyxq+SBTYWOG8utX5aSS
q0iSLMVi+JmSVNLm+ULnCG09JZi68M6hNMtQ8m6SfiCZ7QV4ZQQ/ec3lfEZbM3bx2ty1e+AYKTeJ
9wpwqLzWoitp7eyi1lW/KEGY3guFt9yFR2bMRrrPSasdl21I12mTRARP8fo7yD0K/9n6JMoZ2NIy
sHmRB2PQm+yVTglz0lUyjU2RHBA1qxN1jjAA9qPzsdFtos+aeO1iSjla0RtJ66NH5rkgOPHleUeL
En13VuKunc+8K3ii7QbGo+d83TNTQjC46xiWL1c8XZf/JX8mTzW9r8eBmDxSa4k8fZs6CJ+1anAZ
9pHJZmenWfmngAf+JFUSezmdcvhMIMenDvtWVCxqblBrjkyYPHg5F852U0JV0aV72X4zF6QCL7Hu
KQ3UxHLQlaE5pn0RQ+RcGeIi1yuAfkSe0SY0fpu1dOfktIIjRPPedBnGiEfejdQG2sBAOmOxz1UB
xWz0LML75HRUPaa7743a4pFnuMDEeIw4gfaDBGpOcYItg3IAnMyrwYr92PxD+smdch27lRgE/xV7
kB6Ed2lZdSm8QkYpqU+t9T+8oRQ6hfdBnZuACSmUrxOU4y1WlMpy/LqWAqeKgDLV9pd//fR6Wk4h
s3xok7nuWU4tbd+tEgsFKlcK/+0YukLAQUbHePwQpPFKTFAG/7Fpp47beRQB7q12Ea9K8JGkOD13
2pucG0YG6kkL7lmwoYXyrvyL9nrTIU12v5sZmlFzlnFe1c1i0SGBhfK1s23VN6CV2Yz/E+kYKtdb
esa5PRl49S0+2+Mm+il5NcdZ24E1kl4TzaWc+/r4IYSC8kPJAJHKFTu6R7YN2F3u25VOe9YTduo3
tKMsj4zji4Hw9MEjtXQbZ9N7MZHOEQc5/r71qmLMwbjC1IZdLGR1Ol91HPOfLGRDZ4pp68itTX6S
jLnWkWZAPSOLw7bO5vhmt3+39zeqtzHWjieelXJ5FV2IBa+BvogaqptjXO/9QOz5fEScJC2L9gzb
bqTkc+HsKaXO6f2mRmIpCIm7eASUniiHO4YGGyTX+Ij9lsFeAb6OmB5HlMXUnK6HsF2DAdf0f4s1
HKVyIkk0kDDD/TDc5U03/8y0T90LdpRDLLt+Ooy0gMMuf8eubsA3jHPjeWhUz0ZkcX0aJr+vqoMC
ZYQwnvDFWoyzOBMUmhKn5loi0EZIojv0XKgJUStRMLeMQLHh6kOPfVHUKn50Ns5MKMZIQO1+lAO6
kwNAWE1/ejzyRiWztYZcW1UbJtlhUZJzZ/hT+cOG+jRUeo1TPmZ8jL1UlYokRTXeLu2csrwN0YcE
iJPcIMYqAul9ld9FKUXD9YBtThuNVTeyGnzbPsYB3BBqAr4ykUmmGFWKUenLj7WTIOUhQjS90N0z
BcExui267cIOjaAIiUTb4CH9OnEGWNcxZESi5cJZg9UdOy0MVlGK7n+sTjliFepZ+Mz7F6hI+Rz+
EFBT5qrgxVFPRi/h+W8OBmYZt1XIhBpDiqzsFOX2yoIU34hw3WMY0faPy4i+Km9OGq8M0sveaSfg
pL2vD7q0Gou8oJMIION4dSTs0/whv4R22Nkjt7lNfqM78h5WfgmzepoVwZCLyotdCX6bq+puE4uf
GUF0DbpuJeGBTtdcsZw48R5j+kMqmA3p8b3QgzfwPOltvPKIGEH/WpMsX61/zRmIOBql4CvIYCc2
9kyMkNjYQWK+JpEOBL1Pn+amImtSXQZ28aeOiDHsRwmAlfMSameSWjng0DjicEF8XNFEbC0xf/QU
Cj5PSNDN45IO0nFWEwlhLPBOq6hvT3W27wyKvPIhkUfYjl2ATKSTet7TqiVrX+uYSVoYqzCYZa18
pJ+GNH3wDsPpmMeD7MylKNFkt5h22oojkcHeQ2pC/JukRoKVW2Nw6xyPsNMduaEaHnWTS2mzjzB2
6Fqm7B4UaMcXE+iz555snvwd132Ie/S1HxEVz0l9XsXUZsE6oWBi62YW4eq5TppRlsWYcwpSEaHL
Qax/E6OJ+RCzKVmglpMmPIQ9ndk+8BDnnjSR3c3edQKxovYgVUUpnSDEDG4DioU6oIgtqby6Z1MV
TW2OwQXN+0zY0wI2Zytu3xuZ5ejfVBVlS2NyXSQk2OBXoihG5XUURQTZcWBlE4kYeCl+JGmh7EsR
SBnZHA22ngqLKQf9KTjZbqGEYJq9B8elynA0zaf0PCXxB6WX6yjXzZQ44vZmywqKIyNy5ktZiA9x
GUtbwIyN0iH/blmKZAEmLjOusIKMf6G8mnOnXY1HeNdce844T0j3IJTlJG/YmohuJL8YFCQVTD78
TCRoNjKKfRcDwjlcE7kWnb8a4a1/v6R1zBQwNgy9uxp/d8HAvVklraKbYZMv7+jbyzPtjnRVb3UK
tLVGrV+w9ExEV2mgnANZZmPb6BEH3EPfQThqxyCJrqUxHHAfKDvWB+e5QkFVcTvvTMRsPcyGa9Vw
3ISOUvJnjQQOX+hxOGMWTzGHn+rUd+/1qn4DzJG+pYbRb/uu0SsjkCF26H9FZxWclHB9mFbWR/yr
GOummzYBpJoW3Q1yFQdU8uVnVfs+NljOIWTHchYS0cDktmSnOdUg21SICEGjQwE+nB/CQwpt/vwF
pNhxJjc+534F406y/0DyO6ISRv/ZIC5qapo/oXOThdV25bXY4ei5zSeR2cn2ze/HY5suk1Lnhsgh
oKvIq3yJLOlkWSe/2ZhXG5AnaRmw9vQxaciAzeuE0CHBtaXKtCGL5t/VRKbC4yYu8blQB16gU1Ek
5giH3l7kgvrjHwEPUKcAQHR4mJJA+Wx/iu9BS1+clia3Q/Se7a9crIgPF7jc4wnV+JU4A3upFwUs
hs0776CHjzQ08YHsa9rWNsmZgfIDqpoVQ86lGD2M+Q6fmzTUu+tWR7lZ6DpVUJaCEpGJXWMMsH7z
bIf1CXEAcRQz8G+0Z7G0GjMyLPnAH3lafftNya8S+gbVwC2QwuXUfiOHjZ4MXCGk8z6HFLxxlZ3Y
alVttIia6oYLXII2y7HvqXer9R69kB5IpnId+kKyH1t8axKNkUG0MTyKR3aO0oXGh37PET1BySre
KFI47wDeexbNZ/dwwplIv7JwKa43SxuoAp0fqxkUuOGd6RPDCqcWUjGpb5pTNRAujmqZb4fbYbbQ
IwmK3aG3zYDO2o7/PtA11ilxBaZ+Bv0EI8tbjQ9+LZqzm9NHPFT4QWXL6QIv0C6jyiaDE+VuuRrD
fMpxDaQNknSmt1yRWg7aoHgBm+qUC5r2YuA/ZOnoJkQpJ6rK7iKfayrFypL4Yc2EbKKBA+fwFU2j
qKg27Q1UsXOfmD0BC8VncrO3fpYPNO4pcQasRc11yho/vaUiw94dFqZkPy408bmtlBPsOxxihlr8
9r41w3LRuNPK1rPSaD7LZI4QccgZhx/ayoF+qU/cs0VroeAGv3nPk/0JsysALeENqBCt/MJXGMx6
QXKEv7ZFE4OKJoePT03tV34vzTg/n8UbyAYpZW6p2C+QmaiaEtsmQIO809Cfv31AoxLK9/f/V3Nj
gMPilqDVDhyc0YKMzh6VtuLk4eiWoHYD1GbCaj6IA/jwPGNMqxkGmKwsINmSQyxqvW7i4hrw/WIa
u4Y/UfHsG3jbBNOYuvX61jp69RwKlebsZBna1kCT97uzB+Z3zj7kwqfJoHbZxy+9tDwwcHFZbV4I
f4+841nW5nLPK2z61HGOkKZ95Jpzp2fAqLcvxc0B5TYTB57TQHNSJGicIRMwgW1vwC0ot4gz0EIk
LY9lCt3/B5z0sYJI/xEXsom20M86Ok0jREHfMA+x0AZbJnz7YkmwhgKNsRNDeTJgQAeFtIEUs95x
4I5eMINLYzFBWcw70Ye/YSDUAdwphb3l1FKUJlPHV4cBklLoUDxkd5hS/UfDKAQv8U71ecHUocXd
+hXeQGXjps8IvRNSFqJi/I3dk/mZZpSadX9hMUp0wiFuqNl52xoPf7JnrJQ6qsC6okAvC1DIKhK8
c8kg68rLrpVzyFQ9OhHt01a+v3621SG3erK5j6WOyQh6go1KwJV8dM60Mo3cm8VviT0cverxgBTk
Au7lR6jtcvr7x6M9GJ6OGbT2FWaiVfapItzbWLB4XapeSsSOJBE/vCvfaF5qfi90H+J8cB5QzUHo
e6O3OxxTRhlwyDEJwYGBp39IHn0nu02/8Ztab+VHHanj2MOUGHpyyghxdiQxMrKDwPGHtd+Uzhcc
GjYm+07NwJqVVYZgHedu+s3+jwcbX8qecu5YmCW15qhTIVg8m7yyItUeeUD6R/KCE2pt7mVEfFGX
e75BEBEwlbH5e4wTsQ16XVrCvJ0thkz4yZwqdGU++QOoSOGG1lOXRRIux7qJGiTQtoQvKtQdvT/w
dcHdQ7yd1LZ47TdqcNlXrQmXbynn+CDS/wEoAEDSmo16BOVUkMPt5gRK4gTPzR61mcH6Ai3TCPEl
NISHC/b7+LulU1GH1bfa6Ur2tKs1VFJLHtsSyx8I72wLINJnr2P6s8XKCLWqSrfzu+FPIzMWvE/D
tilhgPwMKkYEAERoeU1vsyEQUBdqIg41SL/XS6gRNh96f99+fvNmnAsOmbRmwwLe8hDn+wrGIyaM
azwnDJR17SBgxuNu48VeHakiqaWZ6WpBaHKy1+CfD3yt+TIURgt7fprlBtvUgX4H9NKo8ZpgTJjY
sABRGxKbtLn4fPnj1byulMusePG/mBHrVBza3PLMiudxLriyRw974SuM+dxIII9Uok2Ihb+DNqKN
N005TqrD9ZD1x4BIrNTdJnNzHYlu39Q8FuvZQzZiS2JpGpyOzv6BQI4PtOdH+eWogRyMr/Ur0IR/
QT+Zen2UQfffRODlEPQWqzI2TWYNZI1AIjpfIkapAd2kpZFzzX2USiKN0YQSd2YhHF4S1KrQbDc5
vKAdn2mIdrGry3jUrW6/W59xT7kSsftzZgsTuYr4+EjqTCLkmtjEiHCph8gtwTPJGLLCC7QRXIQq
NhdC7X585iJ9wkzeCl2ySXNHxv4Vb34SSyVYmXeBfoziH3DZvBygA0lQsIErm75DQXaxiEP6jM83
YXJFCjLzPypUAJsMZLtTKON0PHe3WSnTcTW07t4gh3t4WYd2uzr2DUHBGJA9IZOjTG6bxHgDviXV
U4ceaQ57ZcozhL4i1Fx3F3yjhKMf97/ys2HR9BxyD+nP1MMyZesLYHLIgalD1VBYUjtXF10lztVb
/AeRs2tw1ShEzAr7afwfdqYINpPvQSKmmhxPQXMtydnR4sI0k0bZ7A3sMv1jXUWkoxHemZZnUGLo
L2rho5TI/T1UylPF3Lwx8q/4zHDkC+eq4CbEZjU9ZVeLlIuNg8XvwZy1lxbmBemBnZhqVd/F7Lgg
XvQtCtGqoT5u+c0mi6jWJSglUH1SLTN4gYpHMCh4/9/k7qjettBPu5XoVLh7kV72hud6X1u42Kt5
+GEGmmusgvCWm9wBiY5V2O+yjXJnsWmuU6/yOAdbrfh8Pz5pWjwXjJnG65ksJdqMs+rXXifyteAs
EDs6JyFHf1Msd2jXbKCVEx3UXCyPH6RR1g9qCaGgo9mMpcS+JGDHKanENPV8dVLaAD/WfdbHny0J
EYf+9P1ZROLDz36dr/kE49XeENPFpBY7R9fg2uXrkn5q78TY3fDTbl64h/LUIxNgpuIAeKwzIN5X
640lg+4z670eYkU+A8MIKeMVRwDr73V8CimlCv+RSPDR68v6i0UXkIephZJI1NYbLkblYHY30M0T
j5Fguq0zm1d9IZCyc/kB07/XGW5zrqbZdgw9zcT6rAGhCvGye1sZgznv2gWWPflVfzT/rvTG1/5a
GW3uNUvg/hsxlxajMtFecAW2QTUhfE2uf9brqi5eMtBusJHmEGRDHVNgiW8dtejJFu9caJvYrvAW
BRfOcMx4me4bvy6U34LUB09oBEc+lRA3U+NVfIvy1ORcXn38Lv3GBO3wzUDSHZR6B4PoUvTu5GsY
GA1FQkWL/9JeaRfeP1ByoFlwvicdv4GHV5TNkD2BXnPd9nfHJ658AddJlS+Erm6hUZswhd3NulbN
5dr6VvdK/Jeb6KIkIzBRce7rxSTY3WTui537vxArumpCefmjMSuglbHJAjll2rQ07oenDNPQ/MMI
cTFg2a20Je90KBS8BN4SY9/IQfKqqqlpjJrLE7JBICKLcLBKocNVVSJm08+9aB5GSpaTKoG1tSkT
yaayJ8fBmqKa46Jc5C4PhrT2eFVj0yxm590UtYxSWoJMR5AzK2wJ+1BRWNsUb1V5d4XG8lSUYyR3
E8OId/yfz9zoSKiOSSXZPHyht8DrcfI+bcHqLX2m8sPoU7oNVQo7pGY9du9eOdGFSEsE0qcaHcxU
KrumT6MJbslubRwvNENkJzb5QoHaTglEmE8RKS5VZr/85g5lnaAxfG0ksoXSr02SQGLPj+Kyefqq
3rQtWvTyKkLZMdr+gtCkKMvGQYbFINA2fvY42mQqoV/Iy02+PWW0YU0Dry2Vo3OKf1mSX957SiCP
0cFLKvo2QCpNyNp+lTWp/+MAWVspfPlc5ov2aTf3UVQdQVnJ0wT3sfVnngvZcj43xtjqA3Nb6uFx
8yMdyOoLA5nxO+ss7y5kwN+C+TgG42yxbtz42IBhj+AmU7F13tNdvQs4xwvqLkzMUDieVpWb0VCG
eXd5dFnu5GNqY7l5sMVZUojLuGwJAojJH0p15TjsF6xLmgX8G49cJ8PRvdrP+09DnoTfRzYRj1fk
Tf5k0Q7zOdv3v4gcxkIAsji0Mel8MGjVryHMqXz+Sb4wK6c4qnvsCPIgmvqs7IMhxN/NGaGTzPuY
/yQ1MhDL3ydkg9RCr0pr26Fk1RhDoVkASRLv9yP2mNM2fuXpqHrPEHmDQ+kbY0o9O5fet9HD7+XY
13j2pIc+1gyrBODBMBT76X4KfF6c9RklI8kOEKbLKhMBWob7CMHA+pNKBnrj/kqBcHqwE+oEU4ZC
ABUzTvveg/ZH83rohU/3u/2tBhfy2DdG4pcjEBJXucA/NbX7ukSvR9HItpWq3AxOQmLNa/f2Xiq4
z7F3mOSQYMuARKShsyCtPk8zR5DxJvzt0ANClyS/X2dkOGpnpdHwb2pPq4BX7e2BVXMEHoBJ3cQC
gLsURAZqkYfej3iBHnyqs7ikOtjaslrdTsGZ8z4MsqUZPhRdzSirfzQHlpYZ3WLlJMJMXVMAcRqT
IQ8e/gCXJB0C5w6V/gdS92S9E8QLja75qvMz25KZLFCjb86c/eumNamap2ki8QsI6axiLsS37on4
JX3n84BfVS0TDOdiwWd7VJ2DwUT1pTYWD40K1UPE1uvQMZ8hvWi2Pg6bGZ9d1j+cMO6L4LQGSGBh
75DuCE0smwa7rw4Mnal7ZBxIgv0qUtSBb/AGGZag8j0IBatkVMFe324LWFoF8rzR3VZ2b9bADBo3
bpYCh45PMCm4ASfq3EQDOwpTnTv/dcsaXMSdheuI66AxnviVdmWuuTwUPNQ6R1IqJJjJ+wbiErxF
aKzdWrIOcXxu0TynuRterccGFnOR38o0acYo6jI6/9lVqdDROTqcFBbjNjrL+LMxl6zJBO+NT52s
1kfZyVrYHgr/8PaxjKXihC1u1NC/0SkwIMaZ+f+VOqZcCJQkjC0X6gNfCRxHihd80/g1CIYIdjU/
Rl3DsexXLnxw6BCHGChLsllS+VrpqLW9ptLuaZL+motFs+g/Z3Zv3t/NF8l07S3PyhYegYJSckdU
gmzhzQde/bamc16ivwk9Xr9bzkLhIIuUSdLsDIEsM79HIU3z2pNqEvxAwbGrQzOIl/ZYWIR3jULe
BYJd4HkDzmhZ/P+WbyyVlEU6X+dyoJs1eDGaYj2oRMnTsCSLALXbvfCVQze6uRqb79mO9aUPbpsM
jwxWe3eOoNk6YAl7KguOVrmKYP4TVOY+ThN8IN6LxpTeGlDFKLVRjR5h07WJSDkG1YE5I6yqmRR8
LGVl6yKlxYQZJDWIypC2VL2iHRpK5vRU2VU9ir8zq/7FtqDg4i07BhkYOrSC+s6oBsjZP+TClX6t
WEjXlUOALoCKWACI8WHbV01ja0eAGwyWjRpnGKLpp4HYwjQ6BHxrqGzm56eS2U3Hs1imrwvam22N
ucy4fGkTosGIZ7ntKKO9C6n6ne3EzwVxL594bOufx0CE23puTvU7bs2kSuZbTZI3uVAWRYiMkxAh
E2whYmn1j4Vb+DFUj/R8Hl0Q1TBfTRu0/blw3DF/LKvvJlY5L7wPUZHBXRMEsTBBUWX4abdmlcdo
ft58GGamlIIP0NpZWCsrLfCYaaJUNKAdvcYSOvq4W395192Gv19ntvQWMVur11LpW2vX862182il
Z+HcNEboNtlpnVTCLyZTarBuSnJDoUnh3vYau+5su7ucWTNbyH89mVZYWk/irAf/GC6ZGmHP6s8E
pqb3Nlak6TaUqEFkI4j0QnKosy/dHla2VhGkZYJ8eaiT9FrWKvRxWUjnrFmM43IcAWg7ff8z0oYr
YrfEzhcwyV4ScYq/i5L60YiFlTvGHtXHQgRX5NrsiGarWTR/p+FDCwZZer+EOQWgGYDW0Aq4LKZL
4umyuX67ZEovuCP5c+/VVY+4Z2um2/BZXBSzcRTPaD6Jx6XlDoXOdb2FM5IxLOR+/pFYqAhgpdZU
d0grn1h2Yl3PKn7LMZiV4F++CaJmjmArsflvs3MOvS6OPl3W4iQMO/z+e3vbrpFHx1YsI4O8q3eI
MqDGjMBsb+cFGbQw2cVj+b0Q8w1em8+dWKRYlntvs5OcwFJQ5D5FG9sr4pDIpEn6WkKzv4rsgSRM
hIXxaPErF1oupFdFslvddAqwaWSr9lontWLZydiDcrmzwp52Vckj8+bmjVCBL7dmzVbXSY3bIaAB
kpLPZJIONlK/uUL6UHbotr0EEWg7vX2V1nEPXThEVyATMoDBb1k35vj+WUh3Sw/KKwxX+A7S6GZ3
zkDGrCLEjaGuqpHCQruJnh1JoRm0QkjLF1xL/j2b6SOYeON5aNNtH9ihcJj471aUcEmi/wbkzi5s
yR10UTShudZJ7FNRgJyKIdp75mzHkBuWUUy5SZoMS6mujW8UvP0pjqV8qpSS6bNu+gSvMCIzK3va
79akyRXFFLcIlusYCTkjKeGITZi/SHMSihI1d8rvwR1JG3a7sdnuLDEZ2zjg6wcMoBvpoV5rPisq
wcQ+qkxDOe2AGtEtRfRZbFLN6oKGJ2t7DhLhXOKenKnfDlWxJQy1q9w5ofLO3BId66D1KR5NEbIt
TTDYvp5OLH4sw5xjHQRnA1nS+jww76PD4O1cw1sa6tFL7ZCZZwzS5DKwQUd6CEUrFlCt5L/oyaB6
MZvErx34wRteGXMFiPPF2IHzKMJPioHPo0CPKy4lbSQWDsVvPqSdcLNZiixW4EDaYY6M5Sqi1MB3
j3bY3TPkcaDajMDQn0cl2lkrTKqrGnMW+C3TcWD78SkuAYPSUuUFz8mKSNwPLQzxVui1D2FYj7mt
ldmt35ESHlEg1XB0o3ECgod4Su2A9cpKjYWCMFUCr9bs6twYLC39/cMaFCg+P9nV0f8gUCbNCmv6
bR9qX+8FZmUAJlb3fNLGGndTDd0GF6vpxFvngZMfsqJJeeduhn8xNnVivw7Dpwarh/7+gNTgeppV
EE8MXMj9EbLDYfolWZe3D8R2359qNjMMnGKLvof63nhQO/kgeu3fqMsaC0DaOxtxC60mXgD6SCa4
mlZ4izke5sypRhgzmbxURSBClIC3D0wCiRVOd0NtOnhxo4CTvA9Kb1Xx6mGEMdnjFVRuuRE7c5RB
CRXxiGoEeUNKHJc3xBvNtJFKbSZ9pqR9JQEpqKuZcQ+WVpDeJUbPtTfPchduvPEP9Ka/P6TkTs6M
yJNzvFjQf+PpGO1m7pQ3u0SF4GOy2dXrn/ujiQqWv20nRAKCnD/9Dts/Be+Uq+D+JxtefkquY7Wb
sYXU1ItSSi5h2OmXQpHBII+OBfJ2zRa5+mTtzn/Btrkttf3qrEPGkxJH4aNF/SUVpbyEYSxqNsNW
LUDzmq1REjE/og2lBHeI+wl2Ntn+pzrJoXzq+m1xTfmUd05ngLke8USbqoKgf/d82HUqGf6UjHd0
PUKziBe9YaTmiW3n3Uq1hCFsTJ6MayvdxHZpFhr9biEbd5V6q7xwPM4SwLoV+FdPos2cyORUbXDM
VRQGG6pBWk6A9dtS/oAnnRDHjXtsU4kYtvwGptm06aMOjmREOgpI13XS1fEMKcYZewyo0zsfeoP9
zd4hZVPYjEapREkGbC5FyNvzL5pX5EL66nqx+lRfuvNnn1p3lKkcioKN9IBdzsCtEdOFLtUhbJEj
xr3OlSBPqX24d7YWGV36HvZO9sKnGkDppGXe1WCujdB2eiWOzRzu8xxrX6t4I7C7xNNhFnbl/NpZ
XFm2PizvHeP4rUCsJDuMbohOe923/TO1Stpnj2geR4nz+7Qx9woLiKHjHUKclKkIL5rR5Ica7BuI
0rmHrPrqx97k9/bVylTRYVnd+lEMTRj6ffir/PxsWOENEmMCwMRWlN1tc6fP5iG5gvC6k9awvv7p
B78leSCwb2M7ydItAouhOC2viX9jiM4p85T+TnUsQgIZgT9TAFi6bl5jKRAyGiAn1tV/YKwb5ZRR
bTu4MwkHgxJsK8YnoRVrrJ0WmGZIjqqpiYqb+kx71pWYd2b2fdKTOmHaq7xyzmJRarELwG0Kt88g
ZGgdjFNLS1BTvPnGbJI3l9dNeT9N/+SNO5BD3LH3eZQ0exaaLzxwBM0zNp30CYiqaaKEFcr3HRKg
mPIMtIShDi3xvevkFp1HU1wURb6KkQNa4oJD6ULvcAsxt83lvuL/jeauszULP48eYGRexJMVCG7P
r9loxWlJycW6uJQtLqD87pMXdVNf73mXgdZCJ/TIG7PJf1vgZq1kQqQolHC1mOvXPvj9i5wqC3y9
OVzQq1VotaDU00XdNzM/f0qc5JFPf0O/Z7Rm6eEzRo5BhwV1o09bwBKaoR7gp5Q9YfplJwuBsNg/
IwlnZ8YG/zD/Mq/7lYe1w835CjS7gASugyX0fpFIpC9bvRzmulSEvpOvFbSdMohHus8ltofcmfrT
HIPhZsz3xifZBlMmsjeDnpD++Ey3ZGuovqpbPUq7eH4cYD2D+lrDxWE0li0gDASPVHRhGkl51KPo
ffZIHu7rGYJuDoqwg/2hMKP5+f/NOhvqdW5ioCAgzc34ynNNGuRrB9VsEO3ZXZNwbJKalZxrmp9h
JqJUQeIMkCiJIH3Pf8iPCA5LsBVXwcy1ARcJTbfVqml+ysiNB0uuOfnMLGl6EbtfAxINLrwHDGcA
jxchktV8qZDeSBQJC58QRe5X/rof4feyita8a4mKzvfUlK0AX3IO7umXC7H5VssqdDEWCMlZlFaY
lYKrEk49KZ9cpWwVgQ+Cn1dk8IdaAvXLJbm3NfO7PFzpaD73p3RpFwm/bO2UAUsckwv8+pnhNECD
O5KMci4nJgthQq9PajdRBsmJKnxz2k+nFrWZo3SUXBu6PEg+SqfRhN3VDhi9LT9age+klWg9w3eF
WxnUMCtGG5eYdNvMhNPTUbY+fHnjqE0SLl6Zdk/rNqCQNoF075lBBRY+hpFGIWEeLuqWHPFGSJxj
29UberFxATdq6Uy32563povWHT6nsinLcytiGa0DDgW+euzJrPCvEUZachhmIEee9TFllKDj51m3
V1kRKkVB85mGmQ66iU9o1zX/pfY+hneoqRImdCPXQpNNIkUkgbxYbwnkzUM5tXI4Qy3j4ibrxgJX
p7O0q9b40JxCcNqwgEeonAJk2xFrVWcdaR83DPeHPhGZjVKlFWkaN7s5yTrEKQSg5Vtfm6Ypt3z3
oGSS+yf0jx+l6obnX59rC+T/aNwAWKW4kjD7cqJernIQnk6buXO9+rYa6uI9DGFyo0nVTW2ksEcI
/EkywAcQnqtlAjkeD2wVro8qNUU240BGOt+C/pbd4k9/Gx2XOc0Be7LJDLHq6/xZwKG3Z0kIUZfi
MJUpA2JXeeSUe5S3K/Otha80Uyg64/KXjzB03VvQSJNqsO5eEZBLcPb0vp6bHyvamwbBAM+pZFwV
VN1JglbhKsbTxbM7PFgbTFIGzuSOcdOudzOpyTrAScYAkY+GhwgMyuL2UY2ZTQQZUjmHkIfVZ0iR
USRuIf2fZwBPq0+gHIC73o/c1WkRPAK6/sAvXDBqlTREXC7K3vYiM1oQSTWEvT70skCiZTdfRL6k
IHNMxfKsJWCsIia7cUemADChzb7qwHkMRy17VyXQGeVUJ5Qy0fI1eu8Sv8tnOdm0M1OY15GW8YQ9
C95/G+CCb0Gk1jy2B4Wb1T/XYJMuP81rUhxl40MsmM/JccXMtZovDYSSe4/8zGbVV7V2VCGmoOMo
1gFQYESXHA+x0vdq98b5a+XAekLT1x6k36rzQefQpwT0jDlSDma920Nf0YGJcZT44rl4aQk497C+
+ZTEhpR3xV6nMuAx3/QBwNDcJTTa/VxFA2gCMQQHxiKluCxZbFza7ZtfvFMA+SFGa/wcxVc36eTk
TbWx522jAWRkTtgMnLL/HzGaFbwNky2++iXPkYch87bpZ7Y3YFBlKP266zkkkOMLoVQ4pgu7G17j
7/1jTTBmPrnMxDZ1dMjKWoeClUKqF1Oqnx7BhCbhvz3184n5tE9k2daJ3wJmQVcABRYJYSQprn13
JkW3uH8hS4XNFQq4/q3o+K/G9NKOLjKtrjduaqY+JpG5WP4+bYZDGMDAW+xLu0zKNjqw/yNswv4y
hdhzKXhUaj+Kj5irgDmpP++pgPGgSL7Ty3X5WhqZ+UzN6ud4dsGF72hWTCKtyo5ymQzuX+n1SWRs
bk8MDGT3VT8nQ8YLz/au5AG2y8hQKOIzFrmR7UNv2CjTNKNSOu4+yAk3VMoDsJMP5ekwa4ZCwyaB
YrqsXWU8+gg6M6AggsWNm81rC4vDnm/0faMILTh0uBUPv/h0oLhPEe3+IGu42J+icN9SInmezXTS
Swt+eI7vogKY7Y3q9xmBTC4XlphVo9oySZrSA0lQoI7+MFbWuIbHkvBLRdyAyxZM8+KgL5Pw5inc
iWCTt4RhTDyb2alq8r6CQM/S8Ykji498BBHASCw+rsW6+X/H3x2o02gxgbZ1F9JDJkcI67khE3GS
aOU0xbFhNwxtse3IuuUlqIL8MOOzouVP4P9JlN47FfAbRFxr596sfhNa08aPiiHZCBm9UkcpghHF
anWGafoI5FEWLCrr3viZ8D3bZRLe4tJBpoc8FTekwicnq6WRlAiH9T3Tc+S8UNYRCN5W9cKiwSxf
cWDYwzren4jhXwGnUAZcETM7ViGGssp8AnSviGQlgjBLAxTJthfm6nIJknrQ0RS7doI5MLqfiuNZ
Xj4oQY1wWfgbkvDgk/ep+II31YMRqIKRzYYMChAbleu/iI/u8cSD6adtbXIi5j4YGnvuLYQUxL25
x6Jbk4ozrETpAzOax2fpe+IucJbQPF6JWix4EM7YPaFWhQuDnhlfwZRTW9utq/WpgReC+SeFb/iX
23GsQUrv50g2s/DQHdACs49AHPZw11AAVDIXCFIOo7UCI8dLygdVd/KEBNviLCOOdHZzEA0wpFSd
9mEj4EXmMRrfRdvLC7HNLiCsXMmyx76+p0tJGiFWcYZBS0ig7dVlLn9H5YqXozMNm2DwMmle5a3P
5M6EYfXsc3TpxMz8D9foz3TEa9grYjIspOEzHMG4eZs4gqTptoswG85IFL2PPSWqAaLWZQ7Z548M
r4n/QXXr1zW/t+qNsEI/ieEzv/M2+ma1weoELfwxeuOHGbcUvsJnFHoAsk17Jj42VSgdHoY2kWtF
8ihMrFOtDE+RpI+PuD3Igan3s76dpHEjol3jlF5ye3+NRHMx2iICMTkYOWHHiusHrajzXXlLGVh9
bHeGeIa9f4Nxw68R+uv0YeNtGBJMB9w57i072AK+UfV19nMFvQCLZpjnojnBMBcNaSVOaoNkwh8W
ltBf8hRE01FZxBg3BVKF9QiVc8L8nT9ro6vAYk56ssse5B/1qgF2mjtxIs2nEYMLxPniX6tmSsuG
yra7Z+wRl87t6fYhxOTEg/umBNvcyjjzxAUuKTM2YAt1cGXWuQ8P1QVWKpFfjUj0E1k3k0r5+gTi
BwqYbl1lgotB3ycxDCTQCQ45CW2KnkIBzVoIr4TvUnNtll46rBGOya0s5Vp6NmBG6Pg7Qvk6Q+AX
e8504LVyyqwviMhVbv03AR7PUmNV1lEaJy9WjulAfSnqTrK+dqODT5qqqkra72VGspaiBzHc+qjG
/sobH7SlXcKo6oEaAiycv5d1TuSNnjtw3OLJiXJ1JOxdeFj+3XaPrhMB1DIt6aAK03OjohYTG37W
4/mIsJ/dm9lbT8xGvmlBKqWyGqMvzX/ZQl9lP8CzuTZeVOm9GLy1f1gfZWMnsy61E5DwrW/hEZWr
TqcJcdvKeGvggHXzRKttTGmcmqijryb5KwUxnsBSI8Wd7/PSSkGm40UlV3lB9FmGAGReR3BrVm4/
9rvugAHcB+qnNGTt3MJJNeXMrC3OC0aMK65o4nk01uxI9jjbc0e6RSJWaYuFRnN0NmjUvie8kA8S
+vWlWABap7VujKWuGwJI19+DnnDsuFz3LS6S7+vip3tdd/4twM8QOw1i0VG6rh2iDA4Vg3VuT/f1
Og5glMFBge6z4apk4Seueg9845R5WQtCeWGd0agkuwLVCbKW54SdG5mR+NKYBpuFCTvhB2cx5o3f
LF0UKSAALBfDjnHEOeIpWJnunX5EIh4wP1OPwO7VYXm74njJ6XJ1p7TaTiyHgRBs2683yM+73pxd
u0bfpOucchq83Oz/3pkcYSjMTzGoEL1zMByvSd3Zv1eEW0s/1OjhQQ/Bkx8zp/x0mkzsvRaFSd6g
JQkSOQxVk3wT2iTFu7+OWU/zUV1+5kpJPWE4SWdVptLgosTCEqvYvVaFcM6MHkef9nD2bknd2YVr
e8rAJ+cHti9QvmKe2ZzG/iBcCmZ+cpn3G1zU4f1jZH83AV79C9FWdqi+q6vpLANoXLzEO3xO+prY
x98FEUUKgMCcfaEkQIlq9nJ+CMmBsRyGoxc2b+Cg77asHhSX2tvZM/Kr/T6IoRDtZItQF4FLPIMz
hk/C0cGD7Ix0diIV54E6h3QQW12uM2iwb73lkDE9R/5c3b5ni1fDoqBq5w0Gfwbxz8xUxCQDanOh
bIsVFwdxXZTv6+p0evodfponGGe1RNMcn10r5RS2pPlpNLgmTcDEoNjTpKmN8f9gqrVuXiwEKasq
/u/XV3oTDSHru6Xnf+tlq0eiMrcY17bOxuKHM2tTUGCt31MMSqNpzv2m4dmvmRSvSc+3HStRmG38
1k1nVpZX9hF1Bd8wKTxPL5NP59hZd9CbbeCDxBb2ZHNS0M6fdBX3UFG4EtTW0PFCae4Br9NbH5ny
0u70P/w1neK+qnqkWgiejEHyE4+yJvX9SQ7tEnv5xYFLoZ4PYcaLvGwRgk7Ij58g09oFqyRLL4dj
3hNQ5qe8y8QvsLgH2Nlz8Nw1wZUwU8NJhqyU53WpFwZG1diw4KYZ+koqB3BOeZAzqLGr7VKR9lXI
bnZp1ZgvLLc1dyQKhWY9GOR37xeOvBFzfmKjieDdaEbiJ/W5+wX4u8H7dzYB3bhkDgt2ekB3XJtF
EYteRhslgZgoJljo/gorbI9eTXNXi3Kz/RaMSNIU6MkU2f/h++fpKteNYSocf9/wPrA15HA76crz
S2NQlhibXzL1QoHDvl2z5ADqMk1TAXvzv72pg6BiLgZ/mO6DJ/F4QYettjJBl+9bjeArmHNhzgvH
1yU8TwqVhY8AmK8Hupu1+UX17zidX68IoglSc3bdoF9nBBaoYmEZNKYiBJHkt1Y+51kOmqhFzEbf
uwsGTwJXc0grskGsjSIEGg/W0iTRkQdR2jIK9DsC3XDwG4WRNsypjt7LnetfsSY+n/AcBFLAjyHC
zjr26F6WWUiBLxnhMS1AfYHP0xNzOm6JX9LCcmT4oBuNqlrpr+bn2l5xn8VRQKOg8Rukm7kp/4jU
UTDEp5x/jBgYQq5XwSODrNGDKmky9MBE4etdPmkvvU1hPFwrm+jExQigyJIBZkK8T2Nr2xoYwxV5
nw2NYVy1onU71KpaO5/ObP7aAzqXWPnParm54CgTM9ut+XwzV1Ej89Kjd0O0Og8KoH9vcT9m4EbG
hmozZEHZdNHmQ8Yi4OKE1WWDU76cTMWoSRJcd9RSg4ZGG+XkIXziW/RgldcV4K6ysQx9gOgcK76V
/mBfYBKiQC1RQYD1C0GTmr6yEU21MH5/dIUyKhqf4xopeKH/EW1eeShCsv5w+ClqKhZGURycdLfv
ACnLsYyBUE6nBqYaxwtLANWeMugtbRNKjflv/loY3om8didudpCkHO/1JyhHuI4jVZv+6SEhuZ+p
qUnDH+PdYINz3YQjk25OyZmvSV1m5uiFrAtIQ9eTOk4W2n1ABBHT61X1K6eHuQ7BgxKWh72bPGbh
6fxHcvrd9AOGIoxbaAS17o0SLaRXJA4dMX16Cm8l8pviHtynXUFYynrLw/aLyYHrql3BIsT9MxaA
OTUoBnaN5wQr3sEfq/nuMm1678/XEqz5wSPoDF2AF28Af3Ng/etEdBkCvGra5Wd5zhJkFjtFJRzf
dzCmdudUHEn/irbPBORRCcYXdEtTAfUZB4pVHy2ZT0d4zNK3gNGFb7YLqCaQUx9lWHaKYWqQWU0A
oeqe5N5UiNlsy9N5H44zDskksHbJ20jTqU1u29KVWApUmmqj28GMEYKHcjr6GtUH64UwyzwGyTDg
sUCviE9rMv11zbFhHKzQV1R9E3BnnO89ze2N4UjTrnnyirldonAF+ouTd/7bMSghsLSr4JlM39L1
zPCgy7CYK4XMguIPgoKBLHuVx9J5FlP5yDYdekSmVVqtzDmDXF0zGeJq+RUgyL6P5wH86e1ai8K5
ZOWHrIy6RohPYdkFrjAJ5wwa5/oLl//nV3VtN2pR9xfh78V66qPwTk/oVZRwitnCVSBzqgBVk0MK
5Jnt4svuhpdVjWEHLDChrs+8YLpRKk49d3uElVayXIktcqrM0EMKcVKNXEsjeNVjiKHsMPiTIDlm
pTD7cMogYKSzlhxgMbA2JaddpAcxGWO3ibSp8OFsQLKWiQSHz0v2PmimQ2caN9BKaW7FuvZqCJEf
hk4RgH2D1mZJgFh02S7lT/3UhbNNwzunkV06TIaKxecUEL70JCN49r+JygzemCEw+xHOxLKe+HoG
cjths/erD+pvT4Vj3PcKqE3j3QBgu7S0TjytOvnmXJJTdSsodTnK+GM67xpIp/WYEZFHr2nvqVgJ
tyZWHZo0QPLVvxNKNqwK5WBmtsAPhwQEb77CnSCBWno0180WyGrMMZogEzkmKLGDaIqY5sjfEbPm
7SpCKc1N7D4uxbX1W6ufNYeecNj82NVOnP5ef5MbVPcWUGyGNfhmekVTOVEcwYAidgH8+Mx0zY3v
WZnegE+4uwWuYw1m6WWBQwJ1+NOnnbmkwua8/j7XggcgTH3hm5AGNHr0cNugq/BYguwSFIhfTHmt
lSv03PJgncETC6l9CADw0wfTqCDWYp3Rs3CLeMuDC+z2qciInOdroSXnSOA8xypmrUt3dlPssuPD
vNS5+8L7QbQzq/ZOKRNM6/evkSSBy/Ewb0eCMdkPrRABxc9qhkUQT7Ih0JxnpstqG22F5Oy0OytA
QjCNB2T+CARceaacEx9MmwWmXqio09kHlsknGOVe0jL7nwpwAFCYFFDKS0+oT2mTO4k8ytITiKkS
y9T62459iE/5aJdx2ExhVjZE70SF6EYBVupSENE5kFWijIXLKhqlE+ACsk74bKGwvHYqYao+JtFk
NFotXqodBqgsQJ0x5i+daQNJhEB2CKHSr1dOF5NZvX5uRY3dO+PRYEw+gVTMH9xGvH0w0Had6uK9
wEpcoHaSQ9wy/ABM5UBRf9gKJswvrOZuNNyo8RZ0ey52LiSRnJePPrvbPVZXVjNyHUd9Y3fuq4L8
oiNHBvAGoDeLqv6TDAwj6CjfgDkYHe2HxApBK6S7SOTesZDMi6EsKJ+YFtZx2/8z66uOIOZIjQJW
FKltJm2KalzpxAoQPt9st8kRBL5XieH40NmC0XKe0Wm/gaeqwXqQ+KrXBPsxRt6f6dSHMknltihk
A8xpschpX+qIGFdV38Gyp52T/AgUEwrAHpKlDuWren9lZp6FAsHmrOWGmSJZVFpfJ+NKCI/2jeMg
vNLvOIGbdzCK+zF728Yoxn/W35Fh0pSkOktrYaCxf4By5Lqlj7mC4gdJT+1ODQlFNHawV60DxPm9
07uDkEiuTb21iDmTAZRRBfb27URSRp9KMJW9tm2N8Lcc890nEai/NGKmzn+jS1ag8Rv+aEtx9dE9
/fTn4KeouiqeajwJ9E2CbIJyur190tIxSyaArJGXB9SSJwIqvLd46EfcgRGCB0u4Q4pAToJIEo/L
5dleHiaOYTCabU7EQgMPao040WiR73n2A71nFEb9uKDdmpMATlTz6uU1Uxiz9NdsYE3L+C3+ihix
i3r6WxWzzF1pHp9WkH4LzuMNMz3Ay2SIkMarGhYUwlvSCq9WGv/ut6luxBeh5u3LNElIzKOS5ufM
c0DOF6AGyGlIHxVDf4muKIHCVU6SAR3b2UacnlqcDXZzYUdkx9VBBKKk0fBDoFaHI+jDCGJeFkxY
xf9m2qPyH6FZ5cqpmeZicyzCsXo+aTGkZwmPB098TjxD7/eKz051Q5X5F04z9HL58f5yqT3fD7kb
jxt63/Umd5aBach0W/aaMw09+XwIES3+ORLvFLJmAGQUDIlv/cn9Cns8uE4oVj5otAAypF28P6ll
XgXMHeSew672EKNTvzYkwe42E5ATh6JqBZ3fzBxc064ysbIDMxKmOerrFkivKYiClWlz4ychAUjQ
zCIgid0sXpBRDU5YBk4du3RS0pg++bKbwm7JXmIDPEVVYdAukOlat3VStD+4VLkF2smbSppUDiah
M3IqgvM2IKl4IimDSH7RgOM6yPVDwZcQsoypMsao4togdotsP1wbnNT7Qk+4oU3ytVI3jR0sZWjK
kaH9nAuVvEwpbo/vl0/yelo4dLS6HdRdkbJ1kxVZsm/F633jQkeVANOgikQcAnX8L0MvS70wj8c+
9Nlf//pznmwaTsrtMc/7e/tdMWSinClVnIT0SBpvIUMIkaTMYJVV33ufTi0EHdFI03QqGLa1zOnY
hxEU+2G+E6E0sOp3Nu3Bd69vmyCkX71xUuFrpIAG/c9aTxXFOFXzl1Bmmg7tnjY/p8z2hXLmZZJ7
ZSTJbBKzYuNchWnRJXkqb8vJJBT2m1si2Yya7aj2ZdIe0/pViTefyP79A1wyZfSzNnedvLwqqYwO
Jvuk6KZUSsdB0hkyd0H1fGFWa+dCNBeDgm4LKoH4eNYjG4W6A7kft2Lu4t2nNBKETRFyTBcedrt3
HZhBA6+gsnMVqXQt7THiUrpA40oK7EAZN0vOjUfw23M+pe+kF6ZQ3CTRdyews20aKwgIHlxAtMqL
PTrV706qqwtpBEm0aFJOApQyaqGFM100m0o4eyiyFeila/lNc0cWHe0lmtBk4hHb+hmJG+v0QjBD
lMxj3Gy6GkFqSqf/AfWJCpUPk4VgIEqn7ls5PqG27J0rf5EpNwQkMVqp7bT8hCd3P4CVjKc1OvHl
Clyza+vfpG2aATEcZKdNjsJdV0bauGNZzQlOQl6TnVINd3NuJno4f4PcgQohXbI8f3AbSjvm1DyO
nTHn56ahXSY5r4Yf2sgybiET3gHvwqDaUR4N86Ejr0GETe9rk6TXb8GfiyqJ44eZajoswxdPfYce
c4ny2+ulYp6Z3PMv3hJsLgXw8oDaaIkfpIVnrP0m5Nhn4HfVzsRvob3mNQkkhM/BGw8+SuKRK3yV
tpXpsr08eNcJv/4vlOBFT2stcc5qKW/PNWeLc75s9tYR3ARZ7Rqeln/m/YZIR69BFiLDOJWs8Ekp
jqjTNsKXSFpCrgIMIXubYfRDQZzL8UKLCb283ivi4jNKuGMiPne0HpE0lLhF6I0sIk/Djn3SgYhz
ZMFHrjvGRzbkJINE7dVHabpx/sLVm9RbHneUW4vmompOp8RS7kS4vgqdIrXrCxOTDCUcSmU7G5d8
lhAyy4JGy0qzncXTZ1UYIjt1R7S/gt8ION/vfLMegUGdqI2bMhKaRQ1uekisiM+tJCgP/OOJga99
ttSOiEXmya1q7CMLQ40evYVO/sPjORoHgRfYUBhZuwgtlw1iCSOVOAdWRb3YXilFc8xkyg1ElgK2
vA6/hOsc/ZW4TQ5/7FHbvvVUTKNXEr/A+ZDe6O6B4oMZtRDIEaVzvBAp4lieb8GCVfXt7blE2pPn
E4nwfxVqOz7fHGf2ytYNntBHm1fmLcjarCjFrJ5QA0r/CSiHjvEm82CqA2ZYKUgFm4i3RfKztACV
49nIPsP9hevNBvK2B2JFXCIata6zYCE+XTrS38EZCVRgAFqp3jkVUrZas03tFc3m/vvwpr+h7tmE
uPtEE/o6GZOt+FIbDO0lpdanZC8OPGHHcW7M+hn4/j3EZ8vENwFVa9rLB8HO9XqkmHcpGP7+33F7
QwNuQBH9ZiaZUbmcgFDuNY3tpW3SKAnJSiUgiqgQmSNvjZy8NAltZTD1/m5xEAlq0mE64Omr80Cj
W5Y4C7KP0HXNxp1FPQajj6f0eYNLOFzt9yufcLgq9B/ufaxkxcKKVptvLHK/A5Rb7+cIMNGrLdu1
3OOHIL5dbMCUXsMWZrf7FPGpaJPr3R8fu0umSpEpXob3bV3niBJOjsoxwX4D8kES7GCs9vgQLakY
jyb3HnKCIoskW/tQuF8SMVzRPN6tFvGSOg8ubY9xbFqR2OC1Yr/phErQXbnv03JqMlD8G3pWy4sO
0y2DOpgywBZhItJS4jD0cwSnabvEaatyseQyaHqNmDvn6cGwnh9DhbuM4wKwCbrOjzt2BhmdIrrM
BuGcay1//d0oLDKjvwZEcpLUSJAPzRWo6R89lrr56WiTLwfn2X7tJfrYf3JkHfXJXO6Ep6TQNDJ8
SaJuqbIUNVo7uU+tBHjN56qWNsuG/+scfyRmfUrIyerVjD9sAueQ4MQHrWME0Vbrmqpxl1H3j4Th
SmVe8CkAlxa1dbn2/0P0u7VqntVi51XrB7I2gmlFOMPEKq6rITq/Ll2UMI89xzSK4AmWWMxo79P4
0rkJSz/5k8oM/5OjUlUAjfOAayIlXQHQAewrHqi13hTLg6NyCIDyVPGC6HJDE52hkluQMPOeUp+r
XVsgd9RDGMLTyCq/N46Ih5eG2A+LLfHJDkl83uR6MpQqOsR28ioUJ5P4Infk55AaeyempSeYh/qR
ZXBo/0M52e/mRnq4KxuJyFYNG+SPCx3GWD7jK/o7NDpqMHJQJL7q1FkhW2Nne7TEepmDNGY1h0Qb
9T4m9Be2yXfKrKJ9PMcFtCPPV227cqc5OS9Zow6rxUwwaGrutiTuKn7j1Miki1U7D8cDh4feWJ+H
ztRj+7RCa1OEirockFCB4NkDNY3SrYEkQm8wSV/LDXNVE9Q4+HhXWcEFbtGr8eKiFzazGDJS02b/
hZAce8BNqmlNiVldFmFRQwuNd62wvS0v+lE0S14oR/D3EY6l9N2H/hKrh5bjzdApgQEq3STB36bp
mXPWylsShlr/F5OAdQr/KH5C6M2LNrsam4EI5nTSIKGG+vBUEMhWPtMTO6KnphXo8ZQxs5tNbvqp
DpksTcRV3sqcNomCNfEcWRifnF6n2ImmUkoxhnD8P7ysWDLr8AHMDmVUoEPrJeN0VBIDuykEL31B
86MLFrdFRPk39fFS2VUo0EZGR5TbVdyA9OpoqZCYxNHnPO01mEPyY3hRgAPGLtGRiPfTmD3YvUk4
+UvTxOGMPbUUhH6Fr8gpMSz17fBGETzdpe2p9bbQcGTiwAHU5zIKJU7VvuwZ7SJkt//zVWwZsQvC
WAwnTwPJHCTtg+NdWcyEVLL4UGu0n4b2DC+XXhr0TTD3zlK/yF33Oi9BFVW2/mZI2CazImIrS3j5
ZifsBdBTmxhR0Xt76+4aD3rECnvBtA+spNY6dHXSCFck8fcpxLJp539EyeT8M6e8zKG8XUe9ypjw
VoPY/UIl4M93RxUf5ILwKoRHB8RVvSOwnIuu+JfgmXrx7jeuLXYtmf4OQtWVjVqLZiePCaaBudSN
qKf6wfZszXPm7TTbY4GduWNw21I9X/ybWl/Smz7mpGOeQddJ6qaqur9hkGrNHKZQ30fTUbyv02DE
pBaS062+hbsJHiuzAIXol7D/ZxvHr0docPkQdXH4UYSjD0Dyc9obFf/AdZSv1wk3k+cTuXUOvk8H
zMGVM/WfTVoMWVELiZjpBPvH71WhyGPrLERO3zKhxUxdN6eaGf/Y063w+bBAyRCT2JV0pLMbDpsw
ECjKHLepWY39pqC5is3k5TNPeGkOzABzGX9lnfr6dB/uzk5yQOdfEtLaGK9h9Y6D9k6EbUZ+I39+
IDdut/HwCQkuTzDLddQsPrtvVafGPOpxLO8iWChDPZydrRrQmrz2SrFqOJdH7gPJSAB9oVgilYjK
vBBrisTJpuCZUGYwFZIYDxG2b0TzIRAvpp+zACnpGM+2QQVCNI4H7Rhz4n05ncOy4ZKtb40ADakC
PJ2YL63Zu4Y9hJMUQOpXwh5ZQEi+IPO71wzIOlmgrQB+XnUky1O+9fOuOJEd3ReKKCGRovU3gPz1
N2kIerPtikrVtm38jTx9a33XM0VxBVgKz9U6v5+O1toc3D1ttP0g61bC11NTXYxkxLEkoqmKr0DJ
YaZbIwMKcc2zrtsI5FCj9khezsCw7q4XNbd0V9u686Gn2gOjrwufErHXE6qd8XS51HTwtogAbBB2
MxczwKzNJT/gfhOCb2FnLdk7K8DCc4LYSYVDlijmqOW+Opq0gn7latlARWlwthuOCUBhFd4X1bh8
ZKbV5ijogIgExkf/DkHnSWPii6SU7YMOQcYnGMk8LuKmBOCWeLX0xCJJ1VVfyTU7yjmwTNMS629U
QTrwVd9juBk5gYq08UId6qRnuMtlM/9c51kfEUgY/u2OfIaoOpLCNzaUFFL0sQDZZBaKlJQF/CYp
Rw2eF9Ca19FB69SYmDcfacyDGRBsNgI+CwXd5EuJWX03KgnNlt1aLtPXzPSNWkAoC8IGxtGGjIvT
emkkeEV3K8lWdFjRgHoOnsEn/BfSQsi8GHQRCr3gLyxoBaMSSTYCyGluI2WYyhxbUQhY7TFitgtG
pi8/k0hwTMLMVS4XjidCHTLFeJ2YY/qZUkX2Vi7jdtpwlFk6S0/9Rb3nempE+jQyVc0fzDyaOOQv
CGk62XDxDacgfJ5MDidh8ZSPbSG4a1QATbT7codsu4Bw4c/8ycGFjInNAQZLtt4U/dm768SFmQXn
LuPCgVAjBqs1AcQ6Iqk2erWzY2+nGhzcTiSBR//dBk0+IfbGjBGRIunWJPqQzSLGB3zQ5jcH2jVU
0snXX4ujvtAy/Y0H77QhFytO6sgMOChj7jn4zN2KKY62eMoIe9Uh4ko71GsViHb47QsT4Ltd/xyM
ecToMCfeExADqVRrO6xZYzZAihHo60OfVhOR03D8KMppwBh9mSJZAXb8/qDZfrWdYDzNV0Ye5lQn
/H6J/7ucwAq/QTx3oKTHGZB4QGY6HWG/FG0qlDsXB211CXq26ZZ/S112BLgIA+5lJn+HZhZLE71t
5kjrlsETxcmc2MaiWTRBPUu5R4d/n2NBP4LWA/bfGtXiGxrTgIAGPplXgoo/y+DLdTIDFQAelOOO
Vrfxg+K70vcDpakjZeB5a5QM10gRAKwfH7NkiDRaxAY9tGCcx89jLlxhxzN7u7NgYQqPzMZfRgDq
PSRAUzKoW+iLRbn05kV2KqemBvmMxflkpCq7us0JVJJq2l0Fta9txJvUHmAs+BazmfHXZwpiftTz
K+q7AguZ+Y3Y8LT/3SL7BD5ZTMKmFln0w4J+0wagOEsiqe+Jp7/DjNGe8XberK87TiL8ifgzVXyT
/WDxk0BiO0eNF8nO01foOtAIqFfzi+qvngH7mkcsH+xaeMAvXR4Ge4p+V3zMQOQ+7+IMyxUQR+DS
SWaZXlkoDM4YQHiulFwFbFqitvP44jzRFV4lvyWoehkXjXzBT1ejSJsUWtWnnoNwFVerp6PRBDUM
DAhJZRZmpj9VHAt2bo3bYE3e01jXTMbzU3szrNKqqgh8CUepsVHLxAMSRoKdESTb0SPbQhVNOdbo
dxuOwLstu9rs8Id8xRba4Qkg3SNrmiotP7cNianGYFtua3L3acmTehmz08TkpilyCQmyUVSK97hG
4lykPWYY5SYUXztRhi1qAk3J2Sk7XeaA41RWOBstexrbYag14Zl+PsWbh126RUWjC7nIiFs0Ewsd
2Lv+Hz0wWXtbDsqqQXb79s5RsTWLGI/20VoXQ/fKz/CCeqL2yjmZFy11YlQKr7sn8Zlds5bN8BFD
C0/UDjQo3vpAV4+6ZZdM0HIcJtGufZYu1x7KeiZXCqDpWIZ46X+iAq78cbJeWl8dLKdcceOsB4t1
6aadLgIvH2AlOXL/poPy52wAYWoZUX8SNez+pjUoXoNtgdP5u1YSkF0Le6vDspK8Pj9NnpfMqpPW
Fj89eIezHR6BXg+MTE1kgTEuwW4zeEGpcMW/zU+pdCpdDGmajYnalwZcHg0+Q4xAqp0HM4zhZwrF
7eVntP85hCYVdQjarocUTn6hPf8hKRI0dW99SniXl8s5ZvKPbcPvNwzKOQGdL2vX9ZAufc3KT5MY
UdqvSmiQSanWZusy1GH/sCRNLltcxLQUYkGso7/0reXKo3tCsWIiT150dStt7bZp4PTSOWkoqOLS
ldM8wlciddgZQFFQwr0LY0rPNXCFJga+boiN4DoM5S2k7z6gJW6tVndzef49/wMMRFHEnbxaYsQT
yBkjK0J7uZE0eQXhGVHXUE4cUZDvm37QMn2H8HunUW6Y1gTPQ14DpoVDrR+t0e5cxUNyR9pA6iD9
Jg9J6uIJJ6DEr2uzd/eLzPQRqfSKXErA9myEYvK7r8JMisILAyxAoirQyajUpdj49gWwdD6fqL9/
m/FE9xofwQVhcb2h4+eskaRZj65fLeZQwTcBkTmM751ibR9w4gNRiuGVrKsmzF5qC/3Mz66ZdP51
tPwyiDRxuOWjwVyaDQttZcXEQvts2tdL+WMcyK+AzLB9JgSkfAyc/z7K/uuE2BNw2FCwJA6ucg8s
MebUAkEABFm2PUsszeHbnY+/BVUaW4X7X1dvW1OeLPB3mkZBXYNFMNm79IbgFp959qBOTSzufP2j
qVLj0QjEa9Td5SC/cC60R0mi9m7dnitELhWmXefRI5FUhh0YKBX4VANzqXkzULBEf7oqyOQ4GX/l
6h33S0IllAwY+1Dy0JUDvHaYS59kfCIgiuJCSHfukXK3XN1klfhAH+Y5u+NolXiOuKDhO7ZIVMQ+
+xbMQAu1LTCyXggeqaVzzGqdSu6K9Fwap621S5+8HvgQz4jH5pGefCjVF5O8vqf//4gQtpKhgHMm
SFp8mMu7pmJuCYQ5hmS8Q8lauJ1EbHy3rpUdT4oKOdRxmIAnb7ieQxm677rcxq89+oDYqLZmjVq0
F9ptX2U0w3O4fSqEuqu7pMuqAtE7pufky96CAaZbE3SdYcdcsGAfSJdqSwwKH14Un9TZcWdPyZNv
sBB3IV8x3UUWJGzVL+RKDHhSnrmwzDvaln10PNbw2/Xz2mMPSN4uelNxMZP5tpdtE77PJJPKN89O
Lbc4/1urTVnQhpxUHpwG6GlFavm34X7oL7l2RyGAUb+kB0mB8P5mRxPNnLoTqxPdeEaQeynJk0am
jWGd+yd8nWrvrgH1WW3cVN4aAW4dw2zGmdEsQ5Rxjlge0tDM7ABvV7gDTfMUcs+tSW+TLIP7Dxye
45tytrfDzYH9cVG0j1Cn7pthyfaGAB0QxvQmTzvMk4yWsIItt0aJ7Q8yWB5KCt4pBFAjPrAu0bMZ
hmNM6vdt+mqlxjYGh1HJppWon4XKJ41yphLOlDoKZkWn924AIWX3M2jDeDMFkTLznQbZha2h+ke/
7mZ5KKDUdGtC0DX0qNTV5yQLDdqu4uxijSqEEohq8cvud5P8eKM/uIo+fRjJSihu5Dp6MIBkUTlT
XSLuWZSNW7Rvo4xeaZ31TBCniGKS4Oac2brKoj4bRqiQ7mXMsnAXrcix7KTmdy93oVFOP1vlrfsF
D+yW/0eBCRF46wO5jKnY3Vah3e3kX90k711bJGcT7Ut+6a9w7ZyUUKENb5DFT4rsUZR/Ib8Kw9sT
O6IzRoN7ahqpsYoFv/cYAS59Ub9zbXCJVBdRaQLfNv77f2/RT9Ng9RNcsD/R/wIaKPOJYCyiKSw7
DWT1oA55hr5+717i/awpL8L8qOAR6M1iywl2MUiiLM3OaIcEK9vEfbMjA5L6LgUYHcp07CX3itKw
xW9NGPj8quRRuXUHa+70zCStTjC8Iy8cGxkkOUN9yJSn1sAODzJz39ubDDj9/7lI6FP3iZTtStD+
wNhOL39XDKve4T1dauzBYn0hexQr9hCSjdscKuEE2bYPm05/qBRe7q8E4nn1MY+mATK/CS8OOcRq
HF6oEkj7d6mTEXxWPcpjFPfeur5jlxX1X7MedSsJ/EBuXtoyzTYQteMzYuLMA1r74/k3OA1s7v4Y
Hp3MN2EbfIISz3ji/oojIXF+Az3LoeUkEecQ31NVNINQJCv0wO2Qa5+qoNL0jYdMH+AS6GfFm0+w
AaCexe7300tmwI60AAM1gIFhNenRQf8jwx9huQzry4ttWKOsupJPKj72Fav/LinuqLICsDvedYN3
q7vn9+VsidfLOlGx5F13YOE75eQCqe7ebyf7h8n4bN93JXRpXoyI5DxIs4qDvn5pBNIqFzQyahR2
CjIfos/DRhV1gs09B0wqhY7HPEi/mD3Xf7iK/p4xaLz4yaUy6plCxGSliTFChLdCcla9h5lw6Isy
wAnyGiWTLiaLxTELsPTDMbF17JIiPB2OSu2th0cqqk817H5w+LBt8UkmRAPMDy70YAnFjdGThisv
+lwltpir73lWUKsDcIVUQu4dSxfmhlpwsJIpEEjkX1yGjbzRyRcc+YRaGKA4dJo4NSK/ZzosWNvW
t/YSVy++C/5IJra61xzRlXPf2KkqA021zXAIi0DcLSa8HlI7UQAAeBL2VqAhh70jyD1cxGXaGseD
xQC+ukndaJZNKazOjLddIgX73yr7DjJ29EeBQlaOp5laRh6kpKy700A835bgh99ETMRl63Dtu80L
BqAUVtxPKQvjxf7ShmlBfmo1QK2uMKA7+V5E9vr8pVZBQ7qdI/ysCIL3Tnx6QdNJh7lbSM/XMzqF
jPsq95ZXZcb993/wHT7+zBJxP0P19VnHedwgEwLouVFkejssfrb5I0v0hTAQuqthZ2x5PZBebyYp
wTCBJpfZ5hNzG92vf/TFm/9AnqQN9OjSI3QitCovyrW9vitKGRYak1hQL36Myba/T4gsp1SkPxo9
cz3M4ZlEqG+Y4EGR+xmiy6frP8uBCs+LJD/Z16k73/YyxPUhuUHpour9grmpxPV4gOoVK3PQMIM2
Oqg1qaGFuFsM6M6avXNDdJdv8hbsriOlJLI+66/6+SXzIGlp/HOSeF+EBAq1/XBo+3NFMYrdl/D6
eDW7taVF8vF7d1qDrbcxMIVrzKaQDkv/x3SZ030B0NeHch4uDoMlfjxYGWKstW+L8wVlmbJEvV0e
1SVYx2cYKtA+peH1fmQdSqCp+kS2/jEJvyR7ZyZlcYRvOUixH52wAXZHxf2XqX8oFFYiwvMmPyqq
K7RzlFCjSDKdQSaap/+V5dvtifA3UWeEITfHP2jUYa8rr2DhZjQlXzUwqNWdzrfXt+qWmoEGb5sX
8IwKNG0QnrKcNWiLYwzc7DONDqsLAa7qnmODCCBU5us/hksphdIbkOCbk1r86F37tWsWKDdz0aOD
MiMEBUW4HfBxDenIfLyRbyoIlASzcbyEtOAtSZFI/1KbuWM5zFCroy8H0qeQQMYoapFHrtZWGZ0J
5Y7z0eFOnObgDixsNq5quF9nA0AU3q29tlVba3kBqlLApYJ9pHyU91SjUhIRFsvyxsgc5OIGyQG9
zE/sgxWivtbsV8rbN7qvLuCW/LCpgo1dcvsw6mMAtZM9b6Sc67cx++pkwBBOfRn9m0wxDH+zRhfb
JllwT9lBoIex7tLpJ+YAz/Uyd8mb0RACKBTCNmRFNiVcaaRZFiyjdEFIr4z7VSXmWagbfMQtHugF
UInKYqubNn3Z3xYcY2KEX3hd+/Mb9798O90a+KtiFYMBmPQJcTg6E8SIOYU42K2V1NA1cEM7sQLi
OHzBNH6IK7dC6KZOH94QZOK61U3UsR4fgWc4eNajHO1uPTAVJ3h+y0oLm7WJ2bV1hDDLCPUSjDoe
qt8F4edq0U1DvQzhhym1SQSO0iLsqRwEv2rU3SRHBEHnl43DaP/DbFHdMLzvNg3FhfstCKrhFOYv
4TAD4EXXecBp7F+6D0jSUGDawhwMSBgeZwlEIySHgehizV18XR1XFigbZaU2SFI0u079mdiy14ZY
o97jAlXrCG5MW/3RZ1FdWgBqHPF2iDvRShMwZQqcnKlozs3x2c49SnDlrKhlYmQx+uVohD2/Taiq
Ae+cHs1WqmIk5rzmb8kH9Cf2B3JsMDInzDNRKDrOatnsFe+Dbhb68QtBADE+TihhU9QOHF0O/DV2
7zgWgZz/b4+6CGaejHAQ3JuweouaPorbEDjhMj7yI1QjEt9Csom7fvtD0p4i0oCqQ6aF7HTR9kf2
QcFXZwFeymnV6QiFi5/EkDTu4vzB7GAo/sGKXyxznB1DfOQGOIobvftmlKk09XWEzJGiHCZ7dFln
rbx1z84y6cmJVmVk5joo3jcJwi10bnrJu3GRQKrLqojTQWetUlSdGUpU+ZBrpGVoUpYKEZLrV0xC
Rp1gbnl6mOson7lXRkP/KfxzRZht8c2JexBqqSjiFkgDAh0K9qLuGJlXdVq9Q0UocG1jl9HVmlmz
xTYCe6JMl4JbfrISC7cvG+QUy2BbYFqYFrBkDSmulXLL6tfRNc203k2/Snnw0JeDboCZmtmdNwct
EpOeRMdGimy/G6KJw9XoA/ZsnXmmsCddvIlPPQH2hMWXb+v9n57OaEQHfrxtIQ9ytnndUkepAuDp
02c7UGwhJfmKQVUTGyeraw+2HVEGnU0aXo1yFYYzJ75aQ0RrZxVeNcWVVc6m5KcXt+BoajPmkDOr
Hs5Yi+rIp4HI0iZVwoFKuCLkIS0LBZcMZHdzHD+68vG8ZxHXXidpmzOAKVNXWDpmMNtnbHO3ZyMl
R+P3kLtF/M+hf+ZBb2A8TGtGSzsAS/TOekGbY5zYfr65F3l4i+QCJ5rCAZvxGF7wRWPveQ3LuOib
vbmnA7LoiM1YlqiJH1vFDbss5daaMb079XuVt1yleN7mxtz9cE/74fsFWFYSP4yWhwGLypLv8grz
9RgQhyJaTyhRxRI/zvEHqLVv7Ik/xAyd1CX/dRIWMoWCrYUGtJqNdblPkfBtcT3eGABooXS2Qoql
N+7iWY+SAJqd9xrSERBlzlkn9wTZp2PyaSWN+zi+DjXihmZdCggT+bORkMa86QWE74c/FN/Ucntn
2jyjlRM4kAF8uPE6c00s2H7zwNo4M2VWdld6NJaDD5HIkB+embBOxyn3RLTmMiiaJNBGrtSbkZFZ
+TIed4I5Of3ZBA/h/F1VDy+uQ33T9A4iOlk2DpA3uZmCn/AL3PgmoKVhTuRkd0qemc1IXVNtWzHX
4HlNTpKMJFg2KjRVvaL1Ol0Ci0TNXDhq9Q1s5MlITi9CPvo+PFFMXm5A+EnBiytvYD559Fdwx130
QWkEHgdYaW8KadfJTw3+tfjCUn25Ck1XXUKX9FFsJ73WdYvfVOMHsRXAwEpnYCShA1iaGcaYRQm6
yxBEXeXXo9zDWbMChWnsXjNh60JRvWkVg4jJHnss7ZU/ZbfUrjAfqmrpGXnwFoe3ahdGV1NMOcqk
H15nUW8TQ4BOG1dZ3T0PwJOVl6XHXrQNBiOh6Kw110eniF6cq45uWHxXObQm07bbZLhu3+hZh56W
FSO4EkdwqZHskeJDxAKxsDjiQxBvYy78nrmSMyvUOtQ/wXL7AaDVs5pmggsll4qMrWOXesoSKux8
NnqEPbFkxX8HupcuKMto101UM4BuYrAVNT++TqxPzE/OHjlBEtDQQyojdWS5425qna0hfMN6g0Ez
0H7CTinDvhDd8VaVpGzT2DMq3jRDfIqrmmrxzcVPwbUt2f8EVZsu4Zy3bg2gHa3qXvSyfNs0OKYC
epCHEuMTqjPFI6rIcblj/cI1hI4PkU/iVg6712LVoJ9GbpDFpVwaoaMUrVvwlEX4nzTvLpThPlL5
lMuk95dXmCRiNPDbqGpy+17cswZY6K9nIT7+t+1YE9t7Ls6xC026+ffWsZCmbO/Ihd8z5F3pOXNj
U5hMQzVzozdk0pp+xwsQGWffU6S5ZMXYPRczfBQS8pJudxdJEYFGfuxjunSmT5t8IlE53U6QEJVT
OizUTFV/wGtYixW+Pw55mp1Aei1E0qc94FfFgUkmVPdT/dXQqOuzJqm7c4aJqt/nB9s3UuZKxU0C
HGDwSZVV9vxVWKgLU/2B4a2CHm6PY4VccZrgu9LLURSHgY7zyJ0yVPAT7oO1zxHdrUGKUIqfaYQv
y31VMXOLaDtIbr8XRq3ckdFurx/MiDEU+T1s0w+SpaNmje6gafRGHS5wQ1olc5QkZh+9Xf9XlLsr
5bkMPiX0ib8YqACZCqd/Tn2NVRBVPHTzN81aYMPfCIceGjg+UQT+hxVq705CvtCDzhwraeqOSHVD
NngIiwxVvHshdLdAqCiarOQGnj3rqUiB8nZYSfECr7cmPngELkEfUREmqzN6acUTWjALOh4XsBZt
kudYWe6skE+Zw6mKawO7BLLACHYI1+iQFZhWzRgPEvUPZTfoXZeQVRgpCErl0OKRht+6srCIqoQ1
8MI7UYbzZUh1tKcleoNTYGggyb7mVB0WN19B/8sarjQ0GALJztAzm8/A9nYOx3GKkdgSgdiF9WfD
bsgYbRd4jPj4jUGxDH000uRFUBcN8BAgntUBJoXpKSU6b71DuZrOT8i8On+CAI2yvB2ikUhiIb+p
JsuecgWFcvz32Tr38KSGGfFH+BDFp5iNcDdJD9EVea0Q6GPgSX7gWikjhEf0Lced1A+dtWr6f0Wi
FZSZyx+CJqTHqAHspr8Lr2WHYh8kB0mHDLbsxIxZyF2Vm5DequM6AyUBzvy4N7T2yl/qssSVzeWb
a1oMIBAsjYeDfiAH2CL6c4p04Bm5eeSEEvXXaBzkKKpsif72pd6w+rhlPhZdUgmQ72/gRfcqF/hZ
r03Hds0DHzOKmtFUmk1dWXs//Qyh2UxPfEPOf0qSC+CrZGkzR0gdPforBAxiLmuIGu5gjNIRaiZp
HqMnLhjnNBFpH3EJQWMf7SmRFVvybRUYOMPIq7oNpCNNAeiywzVB+rIKyyjYgcYnLdwQxoDtmSsB
ClJYLYhhD6WpqyulTGyjLBlylap3Wia0se4X9bLyIFswbVFwDlpHJPXShbeIt+JuoIak/DKKJC+3
ES4XRv7Kt2M7aGeYNRUPo5t5EiOW1vK+CFZoXGnqjX7sUm2DEqfxGT1q0qHbXW/xkiEDEW5l1pPR
md11bJRcrQZe60grzyfnfDtyRK1n5P4g523Pw1IEBEJOvkp7ujOQMmiZ33lUZkAM7JbD/OlVCzTj
lCK+LMCe+pqOQ+dyiJC+gyYDR7ZOTgTa1kh9IBP9gR7vcJwP1Ruv90WPM8e4mNFShb02QaG+yorE
LqSWSdWSvbhd3L7hcGwNsyz3XsK94YJILUIN96XbQic2UI8vpgscD/PykkFBioSIrs0jG1Mxv1Gx
ZUzxKoUnwxts4zUgbFtbnWTrDUtXRBLHMnOqqV2X0Avls27n4XJxAQDi3y2dUXu5oHpGt6uaHlgZ
++HwCC+rhbe4LFoIQ4+xwRCPHbL1R/TFck6AUceTTklbZTKu4GCleOs1Hvj7a5VjWyl7Nu/P4hem
oOe6iEcNV3IMC1U+TXbxccxH9+r9xfbkSkeb1ir/XuvbhCbA0Fql1U0HDlaB7PyDCgdYF9ZgnjMH
CLfpCTlyatoS6lYQqD3FKVCA6hR7ZsgFpEPc2G6/lOovIURQuxF6hgMwF6qTEwCd/Jt9pFS907e7
JftV7uqVChcH9PnIKdnamlm1a35hoHS7UfUnLyhZyTTDlZ7NzHym/cyeWJmOSn0WkelXPAxe6W7m
bK52ClfbvzBaR/JUPYRffzyPv/Fi6T5fW814+AQVzspeII9UYwp31RvgEzzCfF6x2JNiPwbyyZpn
jMOTpD6MrIS2gZLRNCsJ0cInpOHscB675JxvsVowXSj981sJwYYlHF8jO6XehLk8EHZE+6ldYlbl
VCT7DjtMJahA92UldQ6wfa2ra0W4vZYuH++qPZDwJEZ49Ta+qDkxA59e+fmQ/MDUzsSsjZih1jVG
ePYzHxub8QvKthJgeSdv2Q37fu2eheiYKtQc3zSOktKLdgJv3DsamLReoGkJYyU1B3jVj1rolDLh
uZg/PiXjo+/Nggn8GKU2B1s5TZOl7dT8oGv5pIa1uf1IDQYfARc+xqzkPBtfEPmRpxoGjOTSY1ge
DBXgsN9Mtup5SKf4X0NJqjn8Qp/3uKvtQiEKVdOp0cT0O7arSWjKCavADX1URK7vGueVsBH2TwXc
8/VfPu4BUTlYxPHRkqDpPEs43PMcRoqqoYIGiyibUDXJTX5j0GoHHDlnWEgnmMqdPcD5zQqc0tzp
HuBdP41/d1qS2TBF/eTSQG7/SF5N5jjyk7MvS8Q7ezVuuEXxdlU/xqTfY8tH9qQrobs+s+qzN7ve
B135T78zpHWUR5dSrXx19anJRURyboqOppgdYk9QdsH6z5aeiB9pF1/nNWEDXpsobHGNpBx61cJ5
mf+Nic1zyWhc1rc6zL6DsIWUzGKX2RbXMHo7qgzMhh7wVdar2X7drOYY65AG7xCPb0RCnum1Rwo5
QonMBjiab62Y+wWZmz255ryTyNET3vVDd1uLOZLUV81elQ3aK+rr74KMKdAb9JRSaG5LTXCU3aqc
sTyeKABxb7p0fFv7YB5es+Xw3Zd5vQ7zEXE25qsis0wlJhWA4HJoApd5WWdI4Qa80Df89z4zwHeZ
Bi6Epe5IlbNKhCfceYQv1FqDbNkrRjPSErNcJIHZZYE+H514qIVodBVXfIj6fdHI7+CxvqFhRDXB
Br5G4ulE8fC5fS9PTjBs8fUAmm0uB9Hrye7EpBRG+Cszc6sWQAbZZSy9diV9YzaZecSjQ9PB4yKj
ow+DTrveiZzsZWYm/zPWuwChibWCONy3G/CmzqZiZPu8+qMLijbK5VvJ/x4Bf5F5M0JfIzZ+VWGi
mUEcoW9CTI/Q3PNmaGeFdFTOvJwBYcD+V7gJniplz0XzEIBC+ou6bzoJta0ZxsjUJBl9aSHPseoh
Z7dj3pqyu2O/V+Fj7e4Hk3gW7U2uYPdN4K0OwbvpkXG/mcyuP/ykJGsz4CW3myG7r92cb9HcPFIi
grZQE25mnW1LbyQa2dwJw3CQbhtRLThY5b8l/uIRzm1iJ3KgokzcfruyqH5ugODF2zVnJGrTXMC9
VR+Nv9+FpZhmRrxdH/REPtRqc6iMwmahmB5Nf95+8GntLYeErL+AQAkNPJAFM06+WLBKs4QlAKBS
/I4mA8M0sGUUa6WnjUq+1kbhXmj8beUQtfMWBVLh1pUeGhhK/FAeuouJMw3YaGtalsvHU2D4EG96
+SE2gmwaSmW1OwLg2uGWD6Ok0e8gpMllWeG5rky1kuqpVBuqPKdFEoW5u22d3TUHtleFoL/hlhz2
0B0eAPKidit29oBuJx7xwimQ+Cqdy43L0Lu5mlADGZXUt/oYIzg79TGS7baE9xSeGDPcZ97kUP/K
FU+KLmw93+Z8lSGbuO2Of6ZbAiIot6UaFPWHex+5SLgA26ZIh5Md9jIaxy/NUrwxye+EOcXeohKx
yv2NGr06uL+swPYLCrSzo/2xNAhKLX/IxOvszSYFl3NuHid0aueQWyXmhxjlk6wr2xV01cXpPB4S
koOqqYOE1OZniWGB9otffz205NwInTu6uB2J8zErkmDUZV7wy8kiY0bzDqklBzgx2A3TIPsuUQjy
VFWePUnkRAkmDXegL0z7OtAMvA6OjcAZ4j5htn4843C+2VnxYkuzJfRMDgClghqdHoIw9XjOf6k9
CNtEoyfBhaStUCTuZoPLmXnRjQt7wDZH97pR+sz86ebfMKnLRFe1EkfMUs27lkkMs8aU76v7M8dJ
Vu/FSZ0QFqiiJN+1RUb2AXXP6oO0+1ZOL0TUk5wx8rCk+jPylKG7iDxiUnOmlE0S41De2JBFEIjl
S8+sTFAKWwcDAqbV/eSeGLd3BmtOScngfRlPIPGi9PLyYDO0Ic0eDxKsWzp/n2xBi2tml9Z8LPFs
ZmXfXFhVTpPTzArHJ8kICAl9s9f15c9wdWyypjWNFUrKj27QggIHC0W2CB4KDh2yDLANt5O3yG3A
RTdMh84SkQM24tggTjpA2UcFNyLnBeTXNPiy/PD9Dotf7dmGMv/Ah8PEBAc4JyLjVB6z3P070h5K
F1cv87EAHrLbXNXWviDDI6Ra52/LzwKlYRBxczQziwOMO4p8jiMuGIW4K4irpBywxhl3OoybVMyE
xzMNWaZ5/2yY9+yHdgE27qyhumjWnGfNkW8hj1Zu/XjBXd5F5lO9dEQqNN9TnGeWggFgJIbwHegw
tP9I4rZh//A0ysJSCc6cms+I+DqSYYfjXvgJhpmyaFLvWhxdPEaU8SzZqWL5aIg340uPYn60Iiu1
DO088BYtSTRQCUFDcIQxe1M88si/dQJmBREOsCOve7iGZylMk37qsIPmTa7/E3VwVNHOZcMvJusA
jDX8eZ8hM2+brnhnhd9xE25hLXt/dHN/7LGKGqyYLNrGN228FGyznzTAkxDKyMG/Htn14mDC4czs
PZEuq6xlfwO1lTR0n8UlvW0Muxv/S4rVTSoTJllYTazbISNf/Z3bdPDxAyz0HP7O+anfkIhVs2+j
c5uH9FwMKPhskcAWe3SvSj383vU35LZz2lUy7xOlFse59KGYs6bytrxW2ieflQmbKmhXnW4SAluL
lvOAAgEk9g6ri56awb/b83p0ZPdDIVDm2dbmm4jH5hSetmmoRTY48nswxRgIwi54lUi5Qwry0X/C
8h/IMlDKmp7Ek8EgLOweMKx5+xNVL22D9hL7yMqxUq81xfbbHhm7vQl6SH5mTMI1Pm0GYl24GLSA
dD/Wa4/L9Na/l4xJgYGyQVQ2GemBolj6wFawnkwpp3DbsDaB+uoRsb4Ip40vyDGu1ednxTe7qt9Y
KmYNkdJHg8DzT2nsdoKfkwDM4RillFVIi9qy7ErKeUZuyr1Pd6cRYx/vClDs3zKMNMW3zf+3MEwo
1NLzWmeK3hVlx3mYJ7L3nEaWnNN1AAwihtJlmIDjjIg39Tx/vEniG8xFaCoY6cgfob1icliQ1xIO
Zc7RzhT5B1GBDbB4KA1ip3bgciE0tyMtqTpmgIXlHmBMx9K3/hoKgQSJeDplDiLJiE1WTKTD3RKH
M9T0UcyjOynGRDpaHJ6vIeDsvtFwP0ucy0RJHQtDHbgwt/5Zirb/WVVEksq/8iZNmu71du283LR6
Ylw9a3RV7BufNJIOYeghMIvZ3MK+7EcHTBFjX7JIXPpklHw6t6vPLpfgIwu/pQ9vxPy8f3rZbiOR
hq8cDr+5CDzbvpGUFLRoHlc4FaLXmF99sTOQO3PtCC4XlZeF1QW4dxdyud9mZMUy95H1Fr8pXi/v
kwSFoRCaRTub6lbgTc/j85fImZgvH9OdfExVHsgvYaeEXXWRsh0Zq2sU3xziU0ylEWmvUP6AnmPx
Vor0707oxfWVMzD/XGNkEPEjcLEDK00vZaMZ6iJGH0TEzleKb+rrSFIbTbQ70deIDNerXVwA0wP0
ZMJotnaPXEVDT2Oqc+eOfDymoah/oXYkuhebSKupxmcL3QWDDCSw9Raxo9zhXZNOrBEBBsn0AUCu
saVNzz3wbNQFCPVjfNeXjpIvDnZdcgxO3st76ry1VaPULYmaoye0h/CSOvwa/+s5bqIE6nVmZIqR
T/QD4whE4Gz9KH66bUmvnUNJgGKPznU2GUcifMP7nFYHfTkcUI0HZfGNrCrEKYw6Ng7sCSjlKWVG
f6xJnq9miQEVyfGfCPqupPestemSQJnlcHqru+IMXGbpcI6fcl2epaFozG1h+4gbmUt7eTEvVpS+
j27IglUIGXO/u/D5nwp1YR95/nzFw8LtyEO1ZlDi8lv6PwNRPsGsavyIK0PA/1y9ONZ20DRY+heI
966PVSAWxoA1uZYTixUHLsh6Woj9bnxC8ybbO+4l8qxgPLh7fX8glBLjAD5ZdrxLaWRU9qXXxk/F
2u7aVMeYn5QN1Jdnr7epWTCyI98d70TANbPGsDFbEJV1x/WVrR10mu9Fz3jzkqADWwO1ii78ynz5
U9Ms3VTCOC2lVCInQSS1v/dqAfo2S0Scjn4Do9fdA8G+H9JhSWKZd1fmnR8N8KVt2GLGkZ9Mv8VG
XxdsGikE8SgoV7UiPIv+JPZ/aux/MJXV9xDMVojYvbDaYK8KQRaoH93O0cQx2nu/MU51fkQsnyU8
tsJ//fhD0+7qzNsrCjyHHjS1gxA2+WfHhGOH+2PpixjilUjxBrH3E2Oifau5hXFc4TRJrVPwJ8Ee
HlTv8dwhxKlHRofvgNIw26Cskiz2zl3lqq+DOnZEMwlRf7RU7KAdW39hWPIk4KvwbQGkHpexO3ys
Ej6RwfnTHAFG008T846cVOd2i8ez8p4w06GLnPSSyI180EVa3p08S4EN7FgtC0BSXDzEfaJ4+a82
+ZvYXwEHXfD3RKdyGVLI09KYtJ4rdNDSWxP0nCkQGPvtI2tj8zkETgl3KwESebw3A16BK8EM/6U6
xinFaXWfFZsq5QcK5Ez8a35EysVNV2AoAoeBs87zI4U5VtlBDn1nGLgUj7qftBSlObyLQGDSjQGR
OUfDGDJtT82wQwBjV0AZaRnsfkSOVqw6iHwqTFWcFvvInHZV24rU3HMGosw2i3krKg6Kw2zYov74
sQAsof72E9DcCnKVLsOrgPJYg7JJxNVqj+G5JG+bWcqsLL43qVBeGidd5V/fM9NHGUPCV3hszJme
x3MEuQjDfSDWB283b6dsDkGn6TB/jrWlGLOJ9Rx0WDe36pH02G+L0SyYpnHrawCGEVsuRgILqLLv
l9xRIquok0LQH4IXySfqeFesLZLU43y4MAxn+WmOzVmaw7HvdqcBOxkF2yPWGD+QU5W+mxvpMfpY
3WPuTQTnDa7uoqdXFZK2RLWKRt4Z3jcfPMcAP69pV6iqGPEINE7Nrdd4ujXStGqF7fwnMKOtnKQJ
PBHY2kcjUceuH6urYABsabb2Ytj+gQOQ89WVa5VYtUb+FsIZtRjOdHFzTuyTFfP0hghfn83BWjXi
YwZlUyme85pDaEr5U7Q6a7Ovz9ACs7L0CncwnxhUPWx6i1+UpS1aFstB02iw7TpRO0Bshlg1mW/P
BPE3QHhTxQKdJgMvzVGCuxuViovAzaj7srLeASXgG1ltvNddLKRmdM6GK/Tu7n26ilNJY1r8Ybed
/GvJzx9jZaPA6c8+ekBuGADLaZbuPbVZSM62lClzRXNDEuCr81Gwbc9u4eNPgF87ECKhIuFo/rjy
SSNzhum9+LvaUFSirN8ExjjAsAdDedBdbr7nixGTlQtbSy4GaeAyNMEKOBBztKztT68um5c9S369
KOHnEwCFym8diia9/ne8CmErFQ4rj+DdWiKP65keAGWwXHsBlt6SZWDGSASMNL7MDRG4DEgQ2mX9
FCBi74G7ZVDawmofwBvYr40vaUIkRiyfc2cE+2XryZSYONgq7uNGGWRHaE93CAthdN6fJKcaJ6pl
JjXu51FQHUHglfyK81hcMcRYNp1BGVEEkONtaR3wqZq2ghMU6pnjAVn+T54657fqcdC90I3HOvCH
jRVap5mg1gPfLdelUJuYAUIX+UgvaTgsiyKFPHSWR5f/pCo45P2wPbyzLWUSuzzTlrdBCn6TyEA/
635wnIH680AKQHe7IM+Akz7lWVjR3T8k/xXwylgYokfATwJaerh0RcdfIeZeFAhO03ggGcFXp1k1
n7yzBV3JxrhwK8pPT9Z0w0jgsN5am8NU7cc6Ufq5Kf8s4LmaUwtSKdNn4K7QidXut6bqCVcfQ7q5
tpx3ooF02PufMIjHWS6LrEfXBvtdLCsQBv5r/F8Kghy+X538di1kc51cPP7MnDJ+actizHRQ5IHQ
tZPOcdNeFckx8Ruh98AP2koY2+L4F7H6qFt2xEvBKSW6sSN8lvgfiNlqTrtjAu7s4ABvaCZWquxN
6aJZnTztxPGkFl3D7cCIMSl+nC0hJaY3BJIQpu7rozHjJ/ArFQVnEd1R662KkU4wUXFF4aV+vAcP
QMk4lWDQ4FfkTV/51C9hGE4k639aICOU8waZVzMn5p7yhLM1EM3cpEUm8b055OnHegcXEHHkpeEq
FHtiYW3v6NKxxM7POICcqBzHwXJAxKso5k4jZYqtnTYImiCUeWxU30mC9PSEIk6eSH+TOap+LeNS
4pHJm9A/kOsmPbiyGax070jvyEYTm+ppP/WJj1elxjxWSdPfarXB2A82OoTlFbj7z3SKddmC2uyG
P6BwvCA9mpZoJcbdIzed58UYQ22sP5id/tWtCI04pkHr5DQ0AMEBHXGov793B1EnThpa4MDeushN
1/JTBN0OBkscotB4jz+PVh2fh0ELVtARNe2wJSYavAg9ig/1ENe2yDRU9wOowXXQ10yKGc4xBaRT
k22hWMqmKW7B7aoZpbuvOYskr8aVIc6unEsAKyCAEiHGVSziJgNUgsNbpvw+xOEFo47y40j8w5UF
JPlQBfrA0E1gk0XfqhP6yxI4GDhU0Hlg0o5V8jp6kfxdRtszq3YKQ6MryFivNrDov6QJuUcRjhD8
wZxUTgEl0+HNXuj87m8IU6MYQkcSsfRxoYbFON+AUfLXY8po2IflORvJCYVhG+AA0jZwhW+r3gxK
hO81hpO990UuhGZJR9vpSBsUNqywp/wxVoCdOr5iSlgPaqc2uvKzIWCWo+W1mjYfG3L2LKBnrwms
pW0r8YatYIj5EFJObcHW3+0c4JKRLuBjY85UeTqXotnV4/WefrtNyntPWdfPFLTKLO/KCDHSU3X6
qNr0FeQ2oUXVZaw+pfYiZYXJ2LVOwuUkHIItEPSoeCRMNjV9z7Y0UpEUtQvis8FtIanOlWsFqNrR
jfhUudvJSug9is+sAc3+epkV0CfyuuGbnMgjSAQjq59xs287jFBPMvR2fxn3ASW1e0hbmOtvNQWg
pvFaIcZuCshlXjJhZtFGHr1G4EqQ4IzNWCgkhVYN70PWvivLD0GwbFkjCTfvW0RopNlZh4FlWYNa
G4s9psmvkXvVaQsLjZpqS3A4S+mLBbQzvaH6blprqw8nZOzfOT2X9Y4hzNsfE3POG0m90A0CShut
OTxQOR36cdJ/2H+2QdTYUuX+Muh3T31jvyXDuNm13FqAHX0aYT1xuBrPz22oDobVkCD3deT/24xj
tOVaEgbVUrTcG8cU5lroBtY4fq16wffgfMnNGKik7vX1tqFno+TTR8GLN5T+cGwhPyDcyhThg17D
vJT0fjiUXV9YU+56jXr+vkF8ISZZbgiU8UdkqyfjHxEea4jrTqaG3KIkRCxwko2iSERuDhlSrO9b
D2LrmK7NZGitWIy8JNWnqILNGVQEw8hVI2m/UT13N+zWJrkfZScxiyHXGppxp60tIKiX+gi/Dg4m
CPnRBCjJT/O2sfbuSHSkuNoFL95CC8Gs2iFqB7Y0XIwoDOzrjO2csGJPT71kxRWGkRDwD2/Nkx1R
nY9mJxfcIVuiTrC9QEXXLDNoCfsQZM9OGRABbZu541v4I2EegFJplKM7Q8P96ridmL+OQLrLt7dX
Sttyb2pcjdSLNnLwSSp/S5R20+X6wN9EyzKTXdAAH0vT8WaiAE7lCddSiuQsyqQ2bkseuF2gs43T
pV0X+1/xoAv2cN9HOQG+eFpGbx7qixkVROAUQyyxypIKSKfFiNBwNcsYqgstf+acUjOqxyjOclOF
SDIMYntjxH9aTMfuh6ZanuUkYjeGflEdkyi2btLmZsexsQz6/8+RI4rhFLbCfitkMVlzdifDUcxD
h8/TWFvVvBSqoq1lQ+Bd4HItXjXgAkGF0rCO/xhhDyarg6wEotI6qeOYr5eO+zQ12LovAwhVV4BV
vu3wOamEJJEyhEOyax74G6il4AKW5Bq+KwEFOoGgg8Fj24i+gYMg11DY0cB319dsEDTEg9Szo9yu
xPZ+5ZR/BohrPv4pUOxvx6G2vPIV7iCWoC3ucFni307K1D3QIebxXtfNacbSyTZup6O/pvSW1faV
QP/3uKo08ltlnHjkNLdrCFHkNkHkyt7sHyscgjT5RVFr1EHt/K5r1PUa08z9QaLtFoRvB9bCE5T8
o5ZOqcQIEVqcP8fSsC2mE/dVQeUn1n/cSgQ+sb0zoIoG4ECohzs1l1iAxz7D99Cp7wNT8XyaK8G0
ygvrAJWo9kl49Is1l0i/+Ub/hotyZRID9YWEhPCWXfEAIJck1CPn/gLsyzENbN6zUUYgNXV3bLVx
RFnnmz3peOdWtFpOTUWDvSddMCCpj1413LtV+zpxG60vMWtLSJBzZ/A5+dGQzSRNninfqZAcCAzV
V6GvCEd5gz+KlAZtkFGtWMbNF61F8SdjicE6b8BqdphNqHQX+TbceNugkuM5H9btC4HGMAqj2fEL
Evnb2bB2VJCz68c8LuPYFXZbSbIHRaekDMVL+LCZ4SyrLEebo17vTdE6tEBY3GWafsdS192h1uES
nVOL3VAIRaIGC42FK35j1kORFSnhiVczq7PzUAfqyDE+7qR7jnWOxe47gn86KkTtpo4fPu7oOHcY
STc3r66+eg3oEB1qo79ujEvfxU3slveYpLRczJ+DqF7G68vEYfh1uAQSMZc42ZweFDRM1E2G8QXQ
Q3ggbjTyaRFlpr81KWE6cqf+sF5OjEoZWrmOJYBslPLeOLLFPm0O4WJiUC20vNq04nlKG4AOrn+c
fHdjFMQEQG5a1WuANsh2Cn/Z8wNIG9NurOsoApGZ+gi93OZRns6FXVEklNhB2R4hWmywv5LPwqQD
w5NUXy/9I0J3jTNIvYWJNBGVDj6qB26wdAgvbYUJzRf40/+ztrFeFrGz/QpNyScIGTbMUDtGYDoa
34kt+uhh+4ruq99uJojI2lVGkgymHoytxI0iM+nnKw9VXK80ObI8/15jspeoX3QMju4y1mbEItNi
WQxvDx9H5h9nvQ4GdefrnhAG+yf3vAQ/nU00TlCwjs3BqDJPM8yLtH4O9W+PDT3sZVMBAX2SDQyP
SpW9dlHsjLFLompXUhxN67xuuf6Ew0ud4l9nrggaVxMVZlHAtC28GVGOkYbyc2vbKroGiOQDBKIp
K2AgZsiGS042whGDMvfDbWIDMJpM2rP44xDlQI4bPlTapjQT02Ny4wbfLHFtkzZzH6Co8kce009+
prvVszUSRtJESUmHr7bA897ucaBiRdCfK95mc1X3pjJPJ4gmmR3VUPgGTcqJlJ8+qHL3SlII4XWm
NMfNAh9mN8Q0/hSWfnnHqykdHhlpf4qwYfFM6wnmX5K/FHpbjQn3NXYygfvH1tUIg5YB7nCagIct
A9ZwUb9uWVkNhB7s0MQyW9LbU8bT2ibT94hzJ9PuPPlind6X/J4Omp3w8OQdVdYTK2OJclkQ2CVX
D0p2UNp3lFaaNEkO9WoNt8DF4Ld6wyGdO+jo+PfrnStDDwCVHhn4hzvIfX4txBSPnBbrCWLUWp/3
LP8qC0+ND89EH8tK4c9kMh0EQv09FauAfcvdHV23orDphvHapohp3oBmE/FyreDmRZohBSBw/DBk
vLzSKuQnPZJuk2jAVXMkPiTilR7kGHDSh2Z3tc2FNol9MBhXqhCMUUbYd9IBJ94zlbHgm8/GK7XX
gOEThFMGlsS6jr43BaMH/0FNSEczkg3siv8ZXvMEgiOVQTFFkUXtZiLh4uJcyOH1y9DIlvlF90RD
aH8ACenT0I+CpMXKdcYvfskwzOqTrdplhk0+gyOWh4KpQfRRqMO5c70xWyxsxFX0+g37wYEA3sWC
58+bmOaN12/MWFsZDNUt4UWnkrI4zF4MBQqhU3VYeM7xqfDSlzmqP7bl1n1ahk3CR5OQ+M4dso2s
wtlzuyCF4HRDep2+vmcozpheahe0dWUB23x6qo1kH62eFZ0D884X3eSqDQq4yjDBXzsFSEQEWcCp
rWQNKrWvPq73apk8in2nmApJxoSuulhKLZdH3guS5zTAAVT+dI+ZBkt5GS4DonET9cwpEFEt0U5F
3+LWNQzmLGmiQ9TT5mtQHKukCyEVC69QESrXgXrOEeav+kLzPcntcPOj6ZcsP8nDa9dn61a4H7N+
yQhwGZAcDI9ZrO2iIJCiLi5/+QkThUayDVC+kXIUWBh19ABhE8C3B9Ue6RBbwPraMAttycSyrzGt
GR37zBblbqhl4d0Ejix/qgjmUYpAkeQqYqbzx9e5n9dLVzojjd2WguaePE1N28/+P+e/FFkMX9+E
Qb9NIsiIVbvNyrK6QeAe2DY06GqSGx13NEYtNBOeyNFKeMZIILbQkydyKVd4MujyNyOpHYuV/4Kx
Qz7sD06JFz4bqqEpwNgOl63Rvoi2T7DSiaeGoM9cVDcW9+oY7uDmq+ihee3czTz+1imNcbs4sKYw
nL37uGGpU7OYNNj1nKiUYFxTlLhwf4735FU5lIoRaFpoKxjIczXegE6I+9l1KVI9Sv37WF3scos1
LUqB+yG0lSWZ3Hsne3Kr/0UNzeXVyHKFdXQPq0O8tpo4pihunD6OSI+FZuJDvW1fpsc+7Lb956O1
/H3uSqvYONcVMN3BFgAaE+HaB/Q6bNMTV7N1SGiZ+0+rN+j+ZcucpmPJFQVNApPPJWM1IXQPATpk
W3QzRc8r3RIJdTiOyQ0OjTNsXJog+gUr5gL+bkVZgVyNKg6rFrPP64FttrMuBAol+VexFT/NDY1D
uZlXkiYt0iwC1lV7aywbX7HFFIPzRKbDRBodwXtAhlw6uGzCJ/67p0QRKE7ze6LPRGrz73XOPlqc
vsgzRLf3yRKzfk6PkfcruTpyFAMrycNRmVUGWvPvt/7mXNs6nHa1O2aohyA0MgDg/ZNSghrKexq5
XpmwPbzydaNkIxc8dvKDkrISRUx5f2wfWMYh+ZRWYGXrUyVGS7vaxE5m1UDRsmY+YOkO6ZWk4xVj
UqiVr/xt1I+eRbybAf4J039j80gfUmXiNTrXoBSlR7Z9mGkFgD6+apZA9lamPXFl1+t11TZtyiwy
Z9Nq4U81XITsvSh4ugyeDeQX5Ham2KXbgmDhUwHPGlvwQrCVE+SOVneKpSsdl2To+CnR+uIcr02/
HcE/SFFNJjVonAbK0+x04/1APn3OhrT0zWtm4V6rN5835e2OMrw9QQvIw9EIHa/IfJCT9Qk0KXl4
XLClJUYRS2umRYEeDHq8R8Xs8oe+cvs4dNKCKird8QDbpa5ApCet7lqXFmm1+O2yc9vq5SZ5MbdW
hLfHrTiL6fpUHdAqiFYX75hqHPoJhh/Mn9scQVRLrB7zhFDH7BAUcxl2bn42Ckr+qAaE1N60it2x
MxPftS6Av6TiUo37xPFc86ds53P3UNniVo5RZd5/madrQrz/fdyDcX0Z/wDtrOrwDYWjXnVyTSoq
6OtDqXn5ib/XwS6dOoce0wtb/Snad8120qvcglJv/9UMYKZwi4sywPWAbIyxalxTkAMmFa4WxL34
I9ZT2FpcoPmmndQZ+At/WvW32h26gbw5KUPkj1Go4HUHRktQbgY4ysignZXQXaTTzH17ki4pN6W/
v/ZyrfzHOJXIDYbO2WdfSrwI6ScaXxGXQqqligDACYHy6NA236cLqe6X6772RojIPfWxNyinkAHw
sShpwRXOFeFhr+oTT3KCjqdV2kuLf58d46LJlbsylgSmaPumPal9T2vNRIeKSw3dP/9GWSjy9ihE
fEQp92o3ORI2jBRheCeurbrwZyGD4SJVKq/PUNu9u0Io+Qt6NAqGv56Gn0TC3pprPn/TYP8G6TqG
KKbUQ6D4f3SLrFmlw07YZkFxbQfWyS2xCcx0zNvPze84jnFQCXPxnd27gprjAtxX/J26kyXrq7wr
9VEjTS/snCqs1uIuYmM9Q2HG4KLB4gLLu6P1ix/ECvFo3fM71xuSWZNxiyGXAvSVr4yrnoRPhdgp
XP+a7x86ExnbeeHIUno2NyqVF17ANx1zVq5YFNDyutmbbHOP+JZAgVBJpHUC9175zG+SGDILVGOd
5sFSEiYFVr8uPrYfVKKqkOy/NFWQYQbZR2QWr39Eo2OplDxopaLuupKyk9vn70XMxvWDxGsDtfOr
Mx3E34CFT57Ih7vuzQoDtCMC+ocLxP/PeNdIIusfbBmaM0QhN14STZNTLnFKyTjD5gAmQHvBmyYR
as3tZpBUS/GHFxDMCsllIyifletWvURU5sj3zV/S50HOf1GDF4EDCjScJfOyBrp2JEPMt4cMbKfr
pA9I8U9Eit3uFVIZ/ewbBBHGFxoCcmbdiZ+EuNGVuiYpSjkx/l4OMY+G/H7MS6qyBoe9XwJ4mpPM
6bVeVGwFKTQSJ8X4iTLQB1MDWus+HVwMRkyY/pK7JrKeqzZmz5t8z9072PjvEoXdTR0xu13vM5Yz
hL+vD2gS4+q2S8RkQFfeMCKRvfVqKCyfiRXh6udSBIOKLlqJyedmUj1u1+aWCKbKcgmQ9i3SUsKi
1v9M6aFL/3qXFPgGWEX8QgN79tE133be3NV2T7dp1BOb1WyS30LeI0BF7/iq6HMYbGHZQEB46qOH
gQW5WyHAmjf45FO9FmlYAvBhcjxesVa7fTtX7yGrHSx0t9HwcWXp6TVZT1AgKq8t307qLRRJNmDi
8IZbn5tXJjJ8hRVeQi3zPNl9GtQtppekf26gCoeQADkztbmGH6SOO+CYcCBS+OP3c4yMVh+INMI3
Zg+qRtx2+KrHXcvUFVnYUtRT225QRT3OPn8CcFZ+zqKtCrrG3QNA3VExqzzgaztgTZUk3UBjw7lA
S3bkpq7yM+56MXOr5b4i34yko0BcumzhuaetnPqkoVuazl7qMSQpZcNA8TshtoISO+ZraFqMJqCt
XFvTGhoDK75jMBxJCAaXxmW7pg7yvygl7UEZsGItvktEfIpYdLki/t6SlyFlV8KI377IBgtRQ4Ml
7/clJe46ruGnNIQI0eoED5QvaJoKMEAPKCDese9rvT4QaroMet5zSDNmm7h1QCPXGkh4bNPItk5U
kQwHZKgtZ6ujUqZIsQg89q9TlraqN9l1JCi+XWFuWKSNaYMM5B2wmiGhG6WTXvwS8DWQ6SwEfCZb
tEvD1jQLzIyzWcunzM+3WMYJc4EzhhPbqP4fzUUVHyIkHpcxrzXuBKQZwpskb8GQpy+/DooKyOXm
k4lMtO1eOVi2/nEYiO6jQjuJRZTsNsJnL/2CNz0p9b2i176x8rwO+P+q65PmW1nc4xAu8ssouCQz
X2dwSgMDCfX/MUY4HO6+6HEJJWovJCaacvIXOU2M6WYbuH0l0vp2roHJG66CDD9Fd8ISLtkcDwus
MtRhXWP69k7O8v1YFjwnEI+QHVGDjuZHuje+OkIWt8GSUU+ccNqu90HOBbowKrM0SuOWLguztPdx
ZXCTX58Sfbdlbj6QYl0XNJfUA3qgVUrMWZLXeY92m7eZw9oXVKhYuK0mmbiEhhNFxURmd8qdU+2D
gqhnf+irvjnzh0uZIEEfrg3M8rK2cdciQvmQgDuV0nkn3NtwFKAAE34ZHEz9XKAjGrpuhmlas43S
HZz7BYewr+pVp7eCK8vvefdxSyP+mfZuZZPoNSFqdtkI9N21kBRKW0Y1k2cvPX6oqRRzswdStq55
msc2+Fg8yepNI2k/IDQcet2c7oDhz/33hp5GhUzT9Lebd0eiB3+baUqws8nP+LwXnrGoX6pTK64y
1zlCYqKzS9addwU7eOCQ9zeKzPuvTtRQI7om+mFOorxjf2pNS8DcS5f8/YGDcxoZEdQo8MjGfq/2
8orPrqt41EHqwaBm610E6rrIgjo6B7DYdtDyM5QY1sGucRYe0r356rFXmQPBRI5GnUy191V3vI8K
0UhpvE5FPMf13s+jbsNbqqKp7UzZUvpKjm0cgsIfobtoN0KBTM78gtVbjHLGOorNVSfxZv6RvdfI
c8T0qn1/YsiN6J7D68iLv04QT7r3soJCvo6lNd9Pfj2/MUnGBVt7yAZNCebtea5A8HmORGKVNK5E
V7xIOwTzjU5M//gs9D1Z+jFMirDwaMB6yF15+u5bz5/UEZXxGCQvsrEpt1O7fd8IDUIcmH76wiJZ
CaGI+DLYso0XE5eRBY+KSBIpPv9o2iJf6uhXF5IDh5f91J4l7vi1OGQKSF82tGQlepcBuCrYH87v
1Z0mtWCyHR2dr/S/aunJ5Tt+ENIN5bDbDANmzUIoReymOKnnhxMRqHd4UTGIxMJIdmH5rrxF23IL
CCEfxwIXqLY9e+zdCDAUeQAb43hxmluhO+pxwNHRwlYoG0sIZQEO0jWKGFB6gzADdAKdj4y4Guud
GwSbINGfNjTmdOiT8VBNtRSlBDxO3v4QaxfWcjMMPZK+EwWe0fTYhiSwl+wifsDqF2UzK6E1goD7
Wa5JZG3CcU6+VqEjXWaFOBm6w8mUtT4hKy/yfT7Gl6kDxzNAkRZLbiQIBv42zDycweTyJNlxVrgk
GXVYVD8P9rOW65ay3PGYP/DwF4TEAHgHTQzezBnCJB/KLhkVZiPGKK1UIs726qvYJBguLUtEdhcM
qADqS1E8il9u7s7faUoftLuMEsyXuoSqiW5m5UOCRHo/f/yHyd8amdhrMLA413SCHMAJgG8PmwAB
P/XGU2hn9jBwEPQdEmtPYkcS4Be9biSMabJM0h5IBDqve/Ik7jI+KZvTsV5Seby3Z+2lCt5tpsV4
H1Z59boUF643iQuwyG/ceRbbKrmRE4/KndTKL8F5grselhLSjci2BXXcQSQBk/6T/p/zj/Q2cNcs
HtT8TJ4lBMCCEzgBtHwTOJRFebq5SNbVX9w79dvqkBYXmDAdSGhpVhpvi1BJj5VFmrla7Mh+YnZy
lPr8PhYNa5yGrw+3/V3h4e5CObPZnLeLFgh46yTdR0YyMDQ26pnCSBZRulpJN7WGDOccee88uwXH
/F2Irr8hjusKmYBFHuqWkZ3KAUV/paTKGU5jlGhtUrYKTl6ApIHaDHUWZuPVo+bssZKpkh0vyh4W
ilYyClZzY/8MkQbJcb9WQuoxHai7dAVyU7K9AJioXzD+ajfVEhcBl5GfY0q5SDzKKDGQKg0jkCf3
K9i/5IRpV+bx6DJGSbhpFPu0WEbflpYwRmYaerAQjTq5OKu8Gr8wsTFE8SZxKHRMmnS84GzcLY1b
PVNig4NuJBpIyzTqL6GCMUgtWHbI+wjBnC9Ar14aHArGEF6evvpclZADLJo2qdkrdZhjIriVXFK6
M+CD+VbWS3nISXlIZBl6Nh6sjCGRtAPhIos1XfNl+cS3x5vDxZRaXWdODqD1rM02h0NMga+2XUuC
DxycU8zY4+Ifd99QBMXnGo6eQH1pz0zrUO8Pn79GYMei3f4ISYWvHbA2a1AHiaQG0aLyIwYbPEfZ
M/Xt5756dENWsy1a2sA9nlLjh8sbi1j/o9rhJ6pfh3oADogrZ2EokDDZSPxiB5ycUNE3TWQBG0Uy
v/QBLQuIstQxi3gNV7FIey9tonyhstmgcyjknYUVeF0czWYA+jvQY8JlzlGdngK3eG7W7EPzFsF6
mKI/4+2QhPLwLfQTw/ZqFc9VSc3TxvmGzVKM6FLxUnw61IAsXMc2laQ2/m0fVIIywVzcbdT93Etv
LGNS+VpRVmQrTdzNfNEqhtaIVVXNaDgBctY24XnyTk6d4HZLhS+Xq7I/6hcXXGpHPT1Icknh6Qia
C9UB2Wli/YrCaZudS0jNorXg0t2O/F9euKoR+R0nqnVQCOOJScu5iwPDEL1n/+jVXKxm8BP2I0hd
E6DNjJqAv0Zigj6zA/T06Tlt10BE21P5RH3bP5GpiIipVSDOOVi9WJrOb0z6bfswL4zRg2nz1vW1
F2qQ2A4U+SBigNIgDSfPyeXhy91x4uxvjnwbpVC1OjZA1pAMDJCMNsrdSVv0v6nl92Glopih29Pj
d+eZ90GoLflXI7IDScelMuxrf8N08aNKJMi/nRQjVvYpCTXnSMwtjRfyZZDDJRB4utp3hcfJX4Ih
LIQVigfl/ZERj6gQh9W+yz3TSwNw+EuTfKYL3R/mMJF92pEtishWIItojqf249ce6Ygy4Lu2rh3s
IAb7rGd6Y6emEcdfEt8kzhHq1MT8PjWsUlJIkOzi8dOA/PlAjiRQcqItbVXfQ4AwHJX9F1tIqB8c
FImrRvm+QZ2OK62gUEyy+m/cIvb74DrzM+nVqc5nOMrpXmgDdozrUZ6RxRnsDP/rbtj5QQ+2WkVK
BXJvGEcUxHVAQWQeMPCGY/NicpsaVM82DckFeXn0AqWqLG8fM4ewNJQWiatNYlB+pN8ngS2Qx64q
aSyaVadEyznF5ki2lwyE/aG7P7vxNTt11WDB9lCc7+Ljd2pvgmPWZzBHXzEOAOB0uZRtx5AYOBxs
HST/KwP1AdcFGJfeX0pYDeK89dClaZytUgVR86wsUdBJtovUGzoBgeRwGRIJ+llpRHJRhtluK6a2
YCUJLiFlBdGXaLpv5qcpDmoHHjbFeFd5PWckAj8y0vkZUGkT3df6rpBQN9apoGh1CzHVQ9/bG8aU
dpWshQvh889L7fYcotZ2vrMkxWPLm4vyJ4KZW8vBMnRhpYHMRHM20VkwmZi2BkwcLDrWNHfxFCr/
cPwZzDmaucqJDh7zEm8m/npJqnkODFoLpREnxOO14MR5TtJrr77EfgKL2YbVYVateZp/akf3fmwu
X03TO+WOAQ6tl7zPmnlFCctvmolD96I5YigmC9WdKO0Anr4BWk1YI39SrAaU7k+90yNEEQMXDqnd
HhLZZYpw1Bax5U5Zu7nRmqaY74YRE4+PuLboDkbopJraKNaf/o1CuZXApsiTXAtrYdRO7Nu5eX6o
tL4o+E94yCNXW7j0xEXRjQLLXYjQ8F9ZrcZ7b92o0iGUD/VLi7l5KdmIdEqwf70IdG5cGormehrk
iUlbdh7/flTQrbfgnd5f6KctzGnLwqBd23+Z2X2GpCNgxHeRvtOHOk8LNA30h3/nAd8Evnq+FYYz
TaKpoaNfJF830jXhoNnwHROR9PupfbwTQVXF2xnxeMbbvHRcvqdcrrS/pZgtnv0hHklrdsCohp8I
9PCLN0mFRSG+B7otEC2eXRozuTArSBg2e20KYLppcrH62PfNlKvp8Y7mWqovTm99wcV+05/YpJP6
cdWWW1oY+dWpCpBF//Oy98t8EE6H8hMfghdrwa6kgSWO2qcMbGKB9WoaoRqzllThI63vhWhl0I6T
BwHnO+hp9xbq9wAgryuobdVBhUxDpJp6r6wg10S4CMumRJVPAGDJ/2pADTa0ScH7B+hniBuz6nTU
eDc4Nq/VBbpH7Kw+NFLF5PsIcyNj3yM9J7p1Yo0Gy3ybUwUPN2KfcZL5elpo7Mgsr+lG0EeRHC4K
sMP+W7qQuVPoVuM9NB3c8F8xid4cal9eGvwUMw3UiB+XWS01uuQ3I0GIVKLOde2rIuCY5vkiz5bA
avpuim3PjgU3l0BV8rE9FCGPWlTP90OSYFbQPIXEkYC4aThO8K9jHvK2ncc907Lr/RcAL8oJz8HY
eWxPINp0xOIntwcoyX7NzWxeb67byosB4YhwKy5+YYA0fQ6EToacQUhGwPkprSKcM/nhZZoTPsBx
pEnPiHy+iBXDmB/jsZukS3rGIu83J6BfibQysqD4fj2/mEVeotXBEriYbXb0EAbnoXpRTXCgF2dm
AltmMODASGFumVDvafFBHeCjPozBWyaW5scs7mY1XD0TCOY363leYDhB9pUMZSRz/L4aoCGDhK6O
nose7HaM7Xvpizs/kEsAP8u8hmvRhVPOOoKZ/KjTmhwQwhj6vRv3hJ09Covt6VYajy+fkfFPNSOK
CX0qnwNp7bQ8xlGF66S2bi9x0lGt3wV1nGyZNZFQ03twefGHezZq2a6OjiNnF2JuBeOz3B+LCaZH
CNdp7VnlBj7MKgPx0wKeduEAuJ9YKSecaEOnZgncxz6ONyjTycdpfC1A0b+IBdLjetWB22OYM9Bz
iF7VBdODyEGM5sv6u2YeCzuxTTu0/9c3meRXJRrBIdyV9e3HtgWRu3h4yqCFF3M587pKBVEewl9q
Fs1vyqkByWYHIfT9HG+J+jx6qr8RNM1sFFnTp9Ux8Ynekg1rvYP0wmnb5TsmvhH/ZLu5CGcwo6t3
1GYc+2QSkUlnRudd7WXjKb5xaxnkKyKFVOwSeiPwz+p3GxdXS0M9BRqjcM0K6XNzHCCFOJ8xlQDg
fgwHgILoQYdOSgWZNC/yQtSn5RUkYAqyyZG1p6Tv7KBqwb3heY87tedgmJ2hEtW7eRL9gciEx7lW
dNazlhcPtIawXBEO3eSO6GzURkSL9vMps4VtmwtVGZYpBfba3NH5kKdxJHkemEEYifNzqoZaC0RS
M/F++TiJvBrya7BRDp/AL0N6JXAxMXQrBESBglt/Gyo3NodvodCkQm+hmfVkImWd5nhOlWGUiiU+
XNkdynLQGVSrphNvtuqcL41CHu+ilJlHXcPvqxR8urbK26l0Qk6e4khGZNMEIQ69hJ9NewL1X/Hd
FIPE3EaxiCxXYZTcsK9QQImV7R19vVIJBumi8SePpHb/Jxkgc84WorUl1SzJTD2qvdcqsybOPh7D
dVpQcFxDdM+y6PkfE9K7RsE7n5gLIqUC9gI/m0Lsp2v2knoL6dsB+hrKe/lXBsDPnE3Ou4V40kL3
RGYzRe/iy8Ve2bMPIMOJQtOTIaem8eQqNwn9ZVvdjVS6e1Al9hefgqVaEfngMhMddIbrktBAsCH4
bbL1QC6oF3WHqpHdTlQaHB2qD6b941hwpqfPg9JI0jEZ+/yYgzpUco43Hi2rHZGFSc3X/bHaOKIt
3JjgOBYoO7R18hgiAV1OvRVOoHfVybSPF3u0FzcGXSyJm1KvIt7zPsnwsxOlA6rUaZGA9snpP/fE
kBNHsDUBwquHFOCzqUDuESqkB+T8kGUqnoTeTiMjH8hYidqYEq7n9UDw2ZcbPT/gfk40OjAUuZEn
1UmaJec0PA1Ya5qtRDT/meDEdIJJK8dttVqfq+9WtaPWPougt3AnwblYRwvWBvP+/N7XRXq71mYf
WNTu9oqg5ULQFQxbqWyGrVU2rPnX0BHWa5CBGIqKWUNzbNBJEC84TNOFa/FueAWsdUrZoFT+1TLm
v2X22JxfKTKLrvt+wBx476oKFzLb3KmBLKMv0h9vPxIZV0KDejn58tx4tH1B7YKagxf+0TGIicd/
Lraiiyi7O/cFaCHzkifd5Q4xXBQgecKRqI+OvBn75JjxAg6Z81gn8N7D2jhXaMn4E6ID7hMeN95A
MDDouX1rmsUqEYO+iZaklyUCKEBTmSzSy3eVmQPNgpmoqi1FoVhCyOzFj6pQ73w0FP9VoCZxP8MC
VvLAgDZEIE0NWwk5LzKC9m4nShLgwOdsBiH2m/ijv1nJWKJvB/mBGPMbs/WzZ8m+PYewE9OLOW7r
/627rn6Y4eY+R0L89EKXlFRG9FjTdFLW4k1C8vkLL1XjDzfAKOIxDjfovezeK+YkY/C4nrPc4riJ
J8hfR40zUl8hA1GHI4IH7G3g0a/tyVxKANtTQKLWIp4hm6GoW00JQP3qfYMlOuvnbBFjFzFi9cr6
LFXPiFFbwxtGrmmsplPbagd5Zp032ezUms7wIb5lXHAGc2wlUnCkVGa7nrSW3l6mvbkC3FRPI7Ma
EUqsyBYGS+oRC/qwpNgMSrcHN/hGLodLwETt6UI0ZNbvz8yyKwdnWh1iO+3u1jOpIv19IR1yW26s
ieTzONa4UbIH55B5Lkq8SBnQtvQ53sWoIocFTC59pa4GXCvYg5PBKkLfg4L07dab2WjBNFhEI+V7
5yQ2ZAKnvY1cvPM8GE52/Pnfyi4srZM7JoENofDXiVkIhT3hcCe53N/7UN3yqyh8CBrXY6PU8yeM
QssTmEUH+I5BbHcu0YTaznQMqf2cLsntzyNS8M2qvh/MUGKnoej0i2m2PPVV63ubQoc8Cyfj70ov
FFRTjC6pjS5gy4lCh/CHsl9R1qUuRycCVsu2CEuLhPWYzz1m/LnUyTqGREPujIN0h5Z7yXqLSijl
QHSOf6fTeCjhA8hOXL9BQEXHMAUvFIo+LRkv4CsPPD+cgUgA/54Px0eoNbjSOasmML0ExDmsmEY+
JvCe0NJCjd3gOyIBhpEJXsaysbXC2xg8Ggii4AbScAd6duJ0YroI/KmaugZMX25RtQv9T3GLTKMN
4GI65lslMtfoEJKfqmIrBJmN525FrQAVohp48jFgbwkXAoGyOl0XgbBTg7WnCWL1drNGdTW2QnBP
u/Oxhlb0C8zJbL9MHi1fl6R/2XQJfUFu7/PeHodtM3/iiyPEiNmeA5MvjMv+pqywSY6sClAennwT
IN/gBjvOyICK1YLLyEnXQkm88QuG07loRTFlFsPHjC1NTN4B6iete9SGbsYgabtoaBph+H7L+Exf
KFkZIM9WxdVmWEsCL8BNLPI9HWqNElcLbcIGGCXUOkV1jizjCC5DHi6kcF9/4svRnIeamh5htbbV
wpBRAAmEDbrV1M611ubN7eKoju8m7Z7rmlqUGNFeicvhy3EoSyzFwz59rFr3YKgA6SsyqoClXTPu
XJ76pd9XkRNjOexPqamiTTfSpEJgpVJenY/q8LaI43dftvP62itBzuwH/PEB2JbM2u7bKuToZf3k
/uMLuN1KrkjlwKHxdFIRPCf8OQHiAZZzlE1Sk8iuL9/zwzZhQxwfeiVeMHZ5QHWFCAjuf4RzhjeF
hmdq5JKgv95b1dWTGwY5uRlvdDvVvTEIAwOItGS4d9yvxmDHzsR9o0Bq9em0lJnQenOkY6ZIiTJd
T+9T3gCFApAgjjgG/nChg0Jy6sjdM/fLWoWcVu/injfOL//o4OW1jKekW/TiihnNSrakVJVJ1fJB
lO4+Fau8/BovHXmjzrgOuFSwVU+6/VcfWoXY5ptsBppSkTj0KmltXtCpzIYuJeLS03cQTydg6MpE
wLfSHIUH8rXDV3I4JDyOaX/A9Vd8c0dxscG/0Yh4fruVLLXaBdbUpzBpL/MFYFnJQjlu5wBqtOOt
6NfGWHP34w9Gvdn1DFSyPsL4Dfa9tupUIUiuYLDHVT2y/A2GS1Do//wDqn8aion/69uQ+343vy+m
dLboKbSlxLmTpkAdGOuWS4sm8c3zMImVqGTPhJfWVl6B5YdiRQsRXKFfVMVx/lW9oCFd59474q0B
XxDnxxS+dfLLN+IUgYH90WrHMLd4Yl1ij+Z7cz17mb/Bi+2r7tr6s/wjhs43PMao/r3EDyhLMYKW
yVvv1vPtAN1O3xHwvZHqPwGX7Cqi5r+i7BPn7JFd/rV76XGXwss4FkVOUkCLgQbJeYLdHhYt9cnR
JL2EuFwiJBegvqZkGOCA6dw66aR8iVy0maO0KAp1n59kkah3smlE0v88VLvnU6Mj3+myReMVBq7g
gjCcOicGMW86lO6K1pe3bk2W8VcPAKGKx1hjcRtC6HZcDHJPnSSD6FeUcmn630vlhLBVdNiHpN/2
8RBusgMKttDfWmq/+Hwf/MtS1UQvbFHeqIOsY6Nywbn4OOXsD3pIVQCAxGcsZb5Wjs6bnXQDmK80
/TACg0VNjIpN+g1rWHgiA3eUC4RI1NAd0RE1wTwrDN2AAKN4Trq2Sp9enyl0vgHR8Pnf5D3D1Adr
Adnm72Jw0ETUcl+AkICf5dBO93JqDsS7zGSTBb8HZ4Nyrcj/SoalDyYICBOeApWjpf29HIMUg4Em
BQT/7hWlCYOR55LkRmvSzlumkzfsDT3psrrIvuzc+RHH2q/9nQQowM+kFEqzdVy1dJV9LMZAM0pM
MSkhoqT2VidLimY1DL3N/0sH8rf9gMmUPc2N0IQ99JQ3u0XxHwg5W5j4GvxP/mX+p8uRItqOoefz
QJKPeUdYJzbwT5SQleQZ3l189jw+0jhA0QSgprFZzQ+LT4jgfbkzYqi337QIiCz1Yxi+1yJs5b7H
zcO2P9fzO/eONGK6gpqT1dSK4DFpjEPpGohyG3zwTOfbaKNSMFgmQuOLuYn5yEbRCxtXRh8VEVS6
xjh7I6TxWYzD0m/SnKm0k3wV8CuFphBQlDLnuLcExEA/ED3fMKZNuWXAajGYSsbNGe10CQ0VEa/P
AaMt73uUGljcW8QNnSY6oC/4OzcK0OkDfC19hQcncdQY6NEG3XWBRzOyDFRdHVl52nJwLjj/aaID
TCPEYX80STT0E3lNv5OVW7lUH+RzeRopLwBc7ZQOHFb6a05s84w1OwlOIob/SPJkV8MSvlgs+LCd
hvfMj92vMdoFof4cGcZR/LoeQGmSmQYanKmgpi6k+HbEmH5SzDVQ+3CW3MWPCjeW6HGGV7GrKa1p
jOn09tNOQx20X56rz0lRmtqicFJIK7Udbdz6zCRR8BUIJCdDZm5fxuudKm5fdgxxn5lbHAolee1o
JmMGXO4oIN/5gU6VSGCie1HemWvvWQHoAGHg4w1tIIEzHSRGu29QvDgpOyhFxp2F9aS+M7SDTHvE
SoB6dZV8Zsy9L/ETplvHj8aabsa6okPeRxmkl4MSwpB30aehFh+6bULec2AdK15DLrGveKMk83aX
p9jMbQKV5RLFQL554jd85X+wau3LxOVOuyp9dcZnM6uIcHeGb/ce2iT/m627J07ULd9MxOqVnE3o
4ewAMfg30uHxVH2kUlKio8OHU/BYnnm54zk8jwDTWCtaGPwCAk+Ua4g6C6PnjUya5XWDjZlCfMNZ
W8thREnkn3j26UYY9xRXrm5JdWmMXOWYs1O8tWSePs1RVjOWcgdSUGsREeEXyhgZ6DR141FW/M37
imsecTmAMX42KufOYEGUZar2II94+4inL4d0nqgX7wr2DSJEeRlErebO9oWubKuN0/00ShFZ+Esi
gThwTAjh4EmUjGDVIrX3ygtjh28Jw8VzzU5FEIgfnR/s9NcmZyXbJYjo8Yjr4XHThRR/AZZ4pHkU
O2ZIIPW5oArwvMJcUBoIgom5WOQAefS8GtbAZkF9K+BdycZSViwKAomznvPb52g/7DpFIY5P3JuU
x96DB11D0xOpzCLB/ndXhhErfB2k8x5eKHlfKLtu6U/2hMzLWPyYvGhtj/H9AjlmLK/plwqLMoMl
BKNREqfVC1Nnzj93JSiF3KqRRavHsAbdQHbftM0GmCL4qDnrbqP1KJnL6KGnCrwNB5Wxo5xmqeQF
/cSFww1hQ/R+IC9WCoJDN6AlubftGDQgG5inlyQRvXdpfJQUSKZ3hBjZJCsB5EwgSkOrNfROI6g5
hoRr77e6/HYyyEIXAEzo3AYu0OXfnI9UKnhFGYlFK+p1T0DMczd5sBa2hVYsg6tMhl060FwByWeQ
w5FTUXUa92EFZAk5tGIFKfVG6Mj0DU7Qy/j5rwCfOzKHUNPmn8ubPLEiMEsqiiEd3ZB/pUhFw6/l
pjs3LDSJeCP/xiB48SyfYpTC1PLMvewe1bIi95LkJEWpOidNLn2LTTCqn4J7KwpcWFfiKgQRMu8T
g7z3dR4CaaF8satGKhqp4ZOTu0rm7jd86Hxlah7fhDcEzjIZtlajE9yYfFLVcGmM0RQerWnCQWdD
YgM3iKB1TkKJpfmd7VY9nCluquvjRcKiEoGGfWlhgrHcYlj8fuRhgRhDhzhstfg49CETajlNtlZ8
E4vhAVbw4qqtUV10fMoxSCbEuBabQilIJz+UmsgZiQmQWmSyloVkv7745M9TLx8xygrlaZ3j4AtX
CfUA0YMm+E0DGSS/LE1OLGfN8OyDED1gZAiYJyLR/2KzRP8Yfu2TSfv6v3Pz3GqRxTcVPyQQDgme
l/Wq9CEk3pC2OqahrOBJQsq2ZzWIQFcHyYkCpm+To+TKKTxsgjQEwMR1uY/CmkdnfdzjUnwUkxZU
h5j+efkuAh0D4V1BTBR0Iy+VCzrNXtuJBPB5M+9MZRviabOpJ3MXjvDm/MglguZGLXam2/TwMMP7
3axcy/4StraxD2ce+LKQ8lENBLNt4WspROFmyEyfT+Qb7Svh7+z2JeW/UqRXU3vP3VNJtxJlWKG1
WD4Vec5v+V3miT1C1AM882FdNQddmMvqtfRO2jflCBVney3QHo3vqs1mifiogplsz1C72dRwELP1
8imAhmnLRAVprBXYTbLG7cLgedAjIXFN6NtUfn+W0GTL4/q0Gg7qY/vpDSx54rsGtnQ084FVheL5
oyXU/mhR5UqBXQYA+p1ZaqE6159bVwmpu4vq6rnDfBWATI0K3RYlUK9LZG3wCyIGx8LKVdPj+XPk
XN0itzQpHST4laR2vau+kjEFCNq3w9ENFI368pNtsU/z9vJ92CrAN2SrD0wdgjSJ+6UdsYCeIVq7
W6ZADZM7AGINmCMjlZ84OIre1cLT+nvXuY2riQM8BB/XHfMcvNS8GdDsz1k6Sw43aW+ZtiQPDBb3
j3R0geF2UrUcZejJr3x3k+75aXt54zLkFUoCvl+4hN3R4qszwNIiV4M+q/p86e5gA5D6SH25iBU9
9RvDDLz23sxPOacgGpS5Y5MoffeylTGh59VvqJ+s5UdzOO1ZZI696QVDE9eCf9kyP88JOInvdH/0
VD21z1gB2BLxQdfXxNdaD5TtAFQLDz2q9zi7odL5Gnd3hEdNu1vtHGBdvANoqFzEvIIU03YRpnpy
ARvN18DEqYXkShR3PbcRTVxJj0koeb2zfdAdWRM6A93e/WIyPXkWn1GFFXO4SIaYmOgKzUzQSwAL
a6zof//H9T+6offmP6MXP4wi0eesb53ee7VO7G/O8tJe1qvLkljlSTX3HxdLX+8X0QVk64yEs7VH
IFbT5oPnjRA71FtP6VPcm44ZZGbxYFUW771E6pIJqaDfLse3xAN5zN/E3v0gGi6lMve+5vxlom/l
iCKMdOpx6Yax+eO9t2r3i18q7MBBFuv69hzq2O1gGu9zZpROmbJBJ3v8sIzoQu8RZR31nEEgpH8p
2QDXFOyo9prpqP18RYHgF0RoS9VIJyChsz+Em6tTkOdOGCyO+h3c4/tFPE3gixM7T2cKex26IlXQ
Btwjc373cCok6ZbCx0GY49Y9mjsqf+429xqt17H1wExh+aeC9W0IajKFUpcbmXhKs48TCZ/zj5i3
0aqEGT1MNnY3+LK072GlQs4YpS2udNuSerzKZ7vPGNEo6Lex4RR1x6UqPxVhABtGM6trIzPYrrLU
xgJhpBzeuuchcrlo3KXTCeqBGmjG6MSWr4FgYV57osMqhPq2E4UMUgW+mrj2le6OyJwkJvdaw4qt
77b1ykBiVxwWKKP+fLpB0M6HKANT/IUBZXrl2pnP/36hvBqOH3bREEE4Ia7nLzTl4rbc+JKpIjIH
5JxTnSwBfSQ9BPcB84440ijCU+KIPazIQaKwaatIXxE6Q9QxkmFKAe3EYxbUlW2MeP4wfQYEwZy7
P06ZVFuCJHug4MhH3x+iFWyHy5htvnU5dLyeZmqqXGT4KVuojE9Xy40peXiBUnwrRj3CpSq6Vnnv
7/ugJntk0tWxIhr3vCjkFCVG6wDY/Fk+r+iiHSIb9iM+jnamyCsm4WofxFArsifC+DSb4lxu6kER
qXTLV83qf7RiA0ligylrOrUNeF+MJ9Ac16Y504rBU+DeXIFXDsxyWMDTjvd1jPjKorfyvqFyhbYX
FpSoRCrRxdHNKJq8AA5TCb7vWA1BI1/Nybyfmx+QPx4ukikrZ8vx4OWP/U4VSErgcWoJLe4ASlkB
uvqKybQaVZpPoxWp0cMh93g8NsmIfnpFaZ5l9XfX/Us+ty77gFbewoP5LGBeeMxmCSwq/Iitvi30
8yHO39tBRz+ifICQsoPtYSrGvUH76F8Q4ErqkvyMeGE6VNSpzkE3TInkxElokvOjtQzw7SgxzyfV
Ekfc3RgdQZuUWaPwNexAPmTxFfEjciH/mieeSbtEryaYp/h2yvtYKwtfN58N2qtc33BlYkcjCU9v
YPX/trSGAib4Imj56sxBfEHU2+jbnF5zh4TBpoEBfN39cKJpQZUUr3Cb5XNjrW3zB5GU2g0l8ckw
JrvEv9P8BEEoz/4UBSPLsljZsK9FI+ygvFlIrR2gycuGnKZE3YlzPIomSlFbcmp2uNJdbJ2yOfuD
gv+5fy2+wbnPB9OXpThXypVHhyn7Kei4Auw3JdLYYAeFH6b1wH8Wm6g1aL6CVlEwEC7B+FVm3z2M
ZjIWYwrJL6C5Tn8oB1iDtqY+s+olu/bpo3DwbFBsYOuwlv3af9W+ZEgW+pwszNVwPqu1M2cx4Vp/
yuD6wzewQzQisiO9ues1OlTa3MCjmAPNOdZoI6PakGxI7C9T4rLq8j1eh/n+RF9UsY/rltH9C1VT
VpD9010ZSsv9XNbryQEn3+pMDp+EAqGpRK4IcIN0W59RDLH9O5wFwLEEZqEAH4VGfsFRx3OF+lk0
SeQRdtWGMaOCBBHfnbj1xpl11L9BPkmN9kcjXZICPZLPwVKPe28RktcjuF1Ci9eDGNyrEypouirS
RZNeyUaGR5zd86+xx7m6f6KIeHZRevN7fLadJlH5qhWhzVmUcRmz5ZEWDnkseEz2ZDFLwUZ9Jthx
VlLpjoi3QLK7FfpEn8VP/AmW6NT61F6qYd07YoFdQzDZ6qt8cNBFflHRRe29hUmKehpuAjXMkNyA
O93h3efCXguo6WaFNSu6oBgaRt59llK2DFbUzVbYORhJqoynz7FD6/rQb9QiSvgMTQl/0+fEPszL
VdshSzxQis0ILPaOIp/2GriPqbvUtRvRLY17txU56SNhWUNzn+m+KvsOdbFIQVRzH64/clDAG39o
2TzBfSYPMKqbZPY7WisCl95cp3h9a1bzVjCSeW4XY5UveNf//xboMsmD7i9AbS7ov8ZyNt8auJWp
qJq2S+iT+yVmmfHBgJMOAYO5LK0c5PEC3UU5shYFgDinn6zycZgs2YiN0GcoEMRQJmzjyW5JTQ77
49wHG1Ql69d+VarH/esh/eCgKo4KM4aa5qswY5K0VzVUkhvY6u4SBkN+NZtE76MtG7j8ozle/XkH
6rSNfKmGBqhXsF9FBCsCJS4guyca0PR2LidKwVZfHrdB4KVDfvosuWMcuVtezX6AdtA2vOPN7ZHU
ox+0FNN5K3mJ5HQKHUqUbgsuvYzqYSLkojilCAUYvewFPsQYQCWXBLhhKYzrVIwogmT4SpR79eV7
zLDD5CNv/Khkfk24Sez7W2oZe789liitUSjGlnC8ZTPiVM0MPWoF5ZQdcYhSqixeVk8Kas4IhtAL
GHb2mYXG5UiBfA4izBLBfpkPg73jl8X8fSJrWqVE7+FVJ/le1FvVHdLXpZbJ2mHA9jmnQyQeutMy
QFeEdxGXeq1UY919eNjQ+uudP6WeJHD73VErirSUSVDfCnr9g0nMNxQWKlU+Ig0ES6kKmBa05KhJ
LK/8wCO+HbZCzPo8vU3TVwso7SxSPT1xguva/x+cg7MHotbfPkwdmla00M9jMFKXbXOiJKbMXbph
h1sgz8R1WhbxuJM1fC+WEVtFMJyNzPZikQmVUOSFbDbBe+KkXfX6Cw54Tw0oB50x8kJFoiHhnonB
jfjfnwz4/CO6y/Mhj/w8e+KeHNsTvwsXuC5iDb1dwUAHao968D16rQNsRd6fsGnoF1DFSiSYBNor
7jLk4wpGROyBnVlbk8bJBxwHFuaTmMOaPxMHRka7IHZxQIOxguo+CRJJk8gOTjUDzGGXuwRUziDe
AWmn5kRJP7Eb9LRfvfkQwPjdIdFv9ADlx6q3HcxPzA0YZgOfk6EVoJKED3xV01hjvxH0oBy8zDjt
/3kyUIEw8JH449duJjkS1WFhZ8Fri2hxrlAVl+tHRnw1dtv3ijUYQWEC/zUIzjzg2pG4eYW8gFv9
32jNV9TE48e/vsrMHhIm62Qpc5TiuEonntdWFroMnQelZtM7nox+HK5OLnc41gaXIa2bGW59OaBB
OWWh4eFqMd0S3iSzUp+t1vx2llRb90/h02AOkAsCaG6nKXIGhmrNlgoHDIVtS/DV1ozVom9H8CLR
wP+TQluDwbgRqv5x8i6i/2r3UownBQR0StOryp3JVt9sAd4hzYAbQ4ct6m89hhVEV1Ri7Yl38Aaw
Gs+dRfYyiR1t7DYaSjeV/TL2Y28v7fE9dcoyJCWWyg1R1rMWXgLDJApmBfqlcwb7McICqa1l0RVg
PxR+WpI1K7o1MGsQHSR2G1zbrD7XWIga398rS4K1ozSFt3wkEx3yatAId3BX707db7DoV0o4d/WH
3n88CqcPxIquXXEwXgMn7WVcfzNuRZ4/XRIj6Kq5d55/ZOtS+8v7mbP4KKZEePaWUDAOCxf4XwIZ
Wcc6+KpL2dr7SXD6giIMWMQHTif/tfYr//4zPWXgIFJB8YdW9nrieR3nIq0NU492nsFDApKORq9z
4+G3x3/+bMvFEY2i9Jgd2lZF4zmjGKcFPDqrHakLITeMdePZn9GdOwuKDnCxV1cjPcp39PIFIH9T
6JUydDrOfwLGG5ZF1WY2h5dJKQlby2UWxdz1jzErvs7Q1Lz1tAewxIeiGBLd5/m539iO4f22kp9l
dFwd/hAaOpGHO/mvQXTdmg5BvX+E7czt++QseA1nDhSrAVKIOzoLfaIqvzlzD1YHfUjVJPuEiFN0
W0d5X6/JtUse6/iSjIsbLky4Ky2wYKc5WKVkLV6/Jiz9pxpsGLuSzBE4iPy7KZBzapmW8QuvIhkw
rMOM/348jlqctUszjqv40VIBv9eQdIOxQYsxr8HWqvimTb5nN90ep25D8tJ6J5/rbtQUzQtL6IQZ
gdwfKzZcpLpYN4PKgClNxYwESTSXIbqEmAGY4gVQLK2IW0sapNNzjF0K0hl301Ztm0WDdEG23nUF
yvJNy2eHnO5aZU7EuhEsN+rQUUKquloxU1D7l1S0j8jY56iDUdSP+hWPPEVxNiMTjhj7FO4QiBew
lb6sJ15d3JLIbdDbpBTY2BY3fV9Wdyt1qn5vjC2DgAr6Br+9vNlahPGxnB2Ej+nvjMDNbmct4S/q
fMVlkh+n4hRbTodC3KZOKntfq7ao20ojBfZP43fVfUFFPFb/7gqRZk5XZtfRowumOAm2M6zTQFco
PGElc1bT3CqclFlbTpH/d5qHh67w/hpRDyu6g6TY+Wfi0zUedN0v8KsMYHlluLhg5Pfiefh3sXvN
gJzqfDShagmy8X6XoJ31dIYIuIzlJ0iF6kaIB5o6yvScsJeRdq/bDZd0J1Ey5abARI9JH9ZGddSH
oKKwgjmzV+XPSSAk3MXy1SUyrOAODh2Vu/jk8AU1Li0xnkRjxf5anyjwMk318FACyufJ8zJEpUEf
1z3T1biKsnPHClF6mJYxAW7MP0FVIZPtxzv2zwGhXIkn7rl4wG+11VTtsJCcLlMlTlGMVdt77BB4
iBqiD/s7QftKeaFLGs4nSpBIhcFFn+B+R8IEaqAtneZN8p/e0Z75xZMHyXX+5cY96+UTMPwKHXSy
P3FaTMpRfqnokbPyV0Q6RAjn8ALzbybbgXa3v56OCMiqYPbMx/Cwbu9YbbdIfd0oKucTnjW6lOYW
UTK+NfGESk3I/15Rb4i0l719S4IulSqj+QKSGxhTY9kNQ8UtIbC8ozQrJtVEvWOOrC3HGFeXTBy4
bMF4z44qCn8JnaFJbRQDNmxV/E6/A4NoTdZdD82jniqjt87sgTaq86wGWKbWNDI6223yb/Reu+AP
Kerr3OWLhqsiFYOg8SveghA/UeWaoSwL4GUdxETDsDPsoL4NkO6PBTOlWNuGpWygVw6KK6RCLOhh
1VK+fJIRRMRFJdOF63es0OS5PVGP9iPwDVstKrAZdBipnRXSUlfikgbFwfxfZBE5GVqVFFC5Pkng
MKxeFw1uVS0Laib/CUFhTJsFHL5Dc7jseammvEKuR0KgJLuOt+BnS2Torm4HP8Z8P+pSHbxKqPm0
OP2JxsDkE4Oe2ScOYXVBYyCZa2uTcRl1stZAyZv8K3ndFQmTvjS6iFs8N1qE0H0JDw1qMJ3BDZEJ
5KHUskAsIBdX+C6N3Ci/lc0F2UpqGi+3MhaBHCxbFdmW8kvYC5PqKxojXH2QLj+3YyTLmjR3TaNF
4wJVzoNMRTBf9Vbjy8aQbQlf5a/5OPZz1FYROOR2X5JkV/2N1fyzizzXLzVsRZHQgzvo7tI68CwH
iEjE+0uF5r6U68lcjQhOBVD51tE+EPRliE/VSpVIiXdHIU+QiV2XtO1MY+7TdmCu89OktKkQmo7r
7syYsPVih+XCgTf7f1SzK+mgd8U2OXfQ3XjMJzqlOKmB8vRavyK6xxiAsk8HmRqGajgT/Ypcd77w
sB4uFrlHH0unY/yAIqOyJCsL0BRgUUMZHGUcqRIlOjBUjLsF2Uw+5cvuGz0XfwT6AQyOK62hFAGB
t4U0zonqLKMwQ66fJfhiChhG/a7fpfaqQEvjhr0g31gvxSfaoUGeprtvVcqnkvrpAfEU9L0a7iz+
fTpEg18K0gkBYLtluX7GCIMu3yonTmLIxxqnG7ypqK6FyeV9kOAXD9S8Ck0TSGH/fRvWrCHaqwN3
KVichbsTIq4IDeiGNojGtelJm6kktmsL/WMCnmGtnfpZCHqvvcafvK54J4cqVNhx/LMNaklq3gqU
kXOsqEG4KcdSfDYwXSRSnpw4dccPJuQTaGAKTbsFe3IxWBKGoH7tZEXUsSrzP5nhOpEmhs0Qjel4
2/Nyt11GWKp3Vor15FWVReDPLMJQIwh3DK/lsSOAM8HoHguLCbelandlKsfwFmsEgZQyf5XOEh6W
CWhhz+SQuuYzWykcplpw0A5Br1AblrUfdC4KY01ZEaNogfup2/wmWaeV6A9RsPtixsj6o5DlmWpe
/0ybrDht/Mby6bD4LeK/BnYlsqgYKkICbg9R1Qc4wQVC6VyIDqGqLtiEuHrbc25nrNr0I5D9KEy7
+zjL9s8f4Nlw22KOlhpDagoxdbI/SwcjsGZ8njUR09kgbFRtv40iEhMNhfgL3rEE0Dp/fWt6TOj1
80A7pneF1KHX8DtEA+WMWrVX0FU8yyQmuWr0pGVXXQPZcGShM8Wmf1CWEsi2kZIMT0LYFHnmav08
gQ7xGi9cryTz6WMLbZvul6tr0QvbJYe0Jlpg0ns/KmIi0j8vcTxLvV3URKgFUo2H4wjNOnX6iJ3V
hDqx7fqXxyB7oKqGh8JB85ToawtB2TYbgnqZ+qyUH6UcjytYhvPr3M4BrfGpIp+bCjeOV1k66Hdf
drI26HesEypG/8G+9QvjFn6rYR/wOnNFVIyQ0ISdeJFyeAv84whOAp1o54eI+dJaSw43p8oN7EC6
tsRMp1gQaauVJcnmuoxjKx4GastY+w7Ld43cswcfAN+ajdIMXkF+zFQyF+cHg65K5ILt23xtnW3e
34QugLcRxl+mN2DXujQ31Kik4021wxCOTvluf23VRHHyQ7DIjQ0ZlphAo7sSoQdmOFzFQwG+bvKx
fac2HckqmhHMvVDDMepI9gPdEyZz/OrNtJesjW9vu2xF2TbRFX5DL8D6zZlGRgzQ1aU3KJ9AeXZk
BxGXoA6rQNAn7iZ1asfW7Wkz8ofpwJBHQaiJnoMb+EittjNA78WJTW3lHiYtRM1p1/kr73bOOxrR
rY1Vp2wYnVvo2e2oiYOUs+TO8Lm8U36acQLoIO/2j50+TB8jyBQgvIiK4XsoYWxhb4hKqaR18jvD
GfGMFBNJijGEF12jxBF2111G2m6ADRwsYcnMM6MOe9/eHOQgCUjKxXCfhldPOkVRbrmXqxoNYmJE
AvxuPLkjGShI5HTjkuLUIf/D3WiscbhqN86D8fxv+wHi9twCjV7jW807tgtehR6SgENQrwXIGRf2
8Lt04KgcrxHlqaQO+N0ym96QReDNvgeRxUwMTr+JISU90S3NIT15jcaIbgegW7WQURnZHEA3Fjk/
7eUJcAsPPJmH1clujsEGqQAuVcAMuGTYvD7plBQSF+IpKi++OiJmF6EiFRqiOiQ9r350To1WXkiH
sp3ytjF4F6UN3z+KBTNc54dE+TTXu7c5ADXXsbiMo9RpCB+fBHv0KJ3Pu8X52GrcA19z1+JPM4RV
wbBGUqXAprUOFIv5nJ3+OnBsH9RakpEK1r0reRKjEChGLHrtOUIQ5dunWmdwpn2MEAq0TOo2Iply
e3plrqpbEC/3EL93kXmAxVRXz+eM6FWO2n2YOx+P4cAiWLGS2BP2N6GBATwT4v04kjhjD0a1NaeA
iSpDg+5+8u/UkDnS/K2+vB4CTswKFsUY7vl0muZqeju59TBd4x7T+mYfyMig+BZyUleOMEHhBoeY
uPc5wOuRGk+eUMnFGoKCQx0czlGnPaBo/w9VIPqULziJfPkq3XyouekUUSiI/OuKNgcKTT+aCBEN
sSSewVvJEFW5orvbk6h8f2mFq0jYmXdmogQYoVon/CCfDpjqgPg0H5vBwpvrgsnMxKa/wJNc0UKV
2CwE88X/9c+RlCtlKsQnzzhcp4ORG8TlHLBAhVWN2uGe62WFKtfljxraXQ6Dkp7Z8yyiy0uYRggD
KgFfBc3wnoIUg2BfA3ejANoedBFrI99QsJCpTxCBd6rad+pWiy99NmtCzUOg6iEhuIwb40Tc/lPZ
1Mh7318JCdGGJkpswNqZvy31dcJ67OvpBghLEVuhTLnzfPEcDakBarYHZJUkuDUwNMAdeEocIchq
ZIjXO4mF3QkLuK8yr9MiT9bW0LPFZ+Ly0BOhWIIqF/i6knxszXZhHc269qSEN6OSlORwXjV53m43
Kx6r+VA9o1VxXKofETALTmD5karudUASdIvDRevJWtUOnpLd0r8PC5Xvyoh0lM6KrbDU+Onti5m+
X/FhZnJhyklgxGnwJTb5Vc7DgV2ARLFcQ3N6NOlgWtHRUu8t6Arm75ZHujLAXBWBRa+Dj+nJCnZn
LiVqJcVTRX3D6qWP9zusnOfjskPvKApgsjZ5t3lTqB0a5RB3aHfutHvjoh5NeAYHOWyNkY1HyvlZ
DXjejhPF4nxDOrApODO36Mi1eXj9VCGBbbVQCe4Iogjlc6csbVaea5wsI1AzKLxd9dggIw7ryUCv
94iCmw7cq49uTVI0b233yYMqFXLHtHe4Ojppuk+sqv6e4CdO0EPiOQjXpScAIXShoTBfNfek9LRG
r0G3JhtsIhZYd+IpJihuMq5r3cAxlzwjwg+7xgypjcMHiCaZBMy5HR2lujgifToEgkkGsM+TxCnn
02k+tjwT4NNJwJ/qdH83osdPzJi0LymZ0LoeVK9cpBBVtRuqn6/31bLW2za7dkDx4rO12JoHKIuX
dLxs96hXLO3sEfn5RlVqD9GX8gJ2nJ7SJxVNh6mBuH7OCvshAZZB158BR099bijLmKa67+3fTL6Q
vnGcBt9inDLz3RZo/e2vqP9BhllP8pfl/aBMUAZPPgEjFfFIRDAkEcAUj5Z0P6LumulXBgviNNDs
wAurvRr9AXi0OsvzJiPNF6BB50Z5vbHLQhXmRcl2wNw6p2oXCJIcvm3KKikwJ/xNMOphw7Fv11UT
k/iuqNAQcLidHoSde37jrEto6qTZNTzzz/R8ajw8yieK1Dt45qvBFJM+XZquRPwPnXWAXnYFIWR3
96mDSUp8QYPAUymAXuEEggjSf4xAfJkjdIGgvw0ZVNK2CMoYmAQJsok8Erba8boWQfjUIuHzp1hb
SRYxLBitSNJNHxa0Tq0cc0kVb3tBYDWhHqI9jnVctiMXuotIjQVcbUP92Kny2bZp8nVw+dIEmHsy
xvC68bYu2KtyGHWCRCIeyGjDlSfNNPtebI3fiBMNotZTiqD9liJHDDQ4GEpUfcxFqJCZH4z/Pt5n
nX1QzdOE1kZ03yMi7PekD2XsF9Lf3nxxi6hUtH6XtKu3rtscYNM6aF5khynf0J5XUtrhzI9hoK2J
EIqLprlWXsTLEOPmxRSxVXrY1tgIMoGW5PkQP/PIf9hRnp4rfL67LRcs45ZvRRZjWhDE2Jv8708M
44d8pOMoUtx/xBZT2F+3s71C1H3r4TobFPAG84dIQjghvb10aDZYAaurxfGc0WQ3nmXmuyitYeBs
x4A1OePvHmlFaPbzzcYNi4HeztaQyxq+eux+i5CPHZB/nnaGphSyh5uylOKXcU43Woa0bEIiQaKl
axm6tH/GKOwnJXaP9DcEfpRkDdmf/s+PyFgZ21go9Rr+u9hoKMJURWqcxeC/Y5Dj8H02+vKDHP6p
PiPwiywnF0Albb7y8lCkLt3gJ2edfst4kjiZYWYIXZ50yzJZ2n6aMgAhpXFcEE1SIEwxbHyqSx9p
WnvXpDDrAVHkqqDlb9D0aYcE3+4AXY4ay3eFbXsYXztis6T63KPuwwCH/AdhR1STELfPqc9LFew3
stxefXuaqX5w4dSjQ5FtmEJ775uC6RH8YDy5w+QXJ6JnY8RlROrtPYNhKQu2HS6GItJQSbrDr5gi
h67H2G9SPEb/5iSVvzkdEVPN/v2709UPkywg4EtmFZSioNEAji2qsAckxg43kOSQ/OZ6aSB/YGmN
89h2Lx8pyo0vu/FsZ8S1Te+Uhp935gMu5ZOp0BKN7Z7Q94KRFBRHhNj2gfW4K1tHvpGPowUFoICt
jdFGK79ZUNLMvfnk3uVV9i+chfYzLlKfcm+eTGgVF6OGhT5Fc/zxXcEQvZXj+RtrsD/1RZoS+89c
2ZXlLVM7Y5awWq/4OR595LGdvg+ioeAA16S+R4qaxJQZa4VrgcgBuYiX9cGfWxXpcOvFXokXKtxz
B9VozYto9XX/a5MPcIai4kYpCyxlbUzBZx0isqRcXapzuuBAKHEwBsVfD1WDVvCL4BHpnZ/OC62Q
x+ITPskekvl4CH6vcuQTnI6t+21E/9plrLfuNH/9XzFcEOtNFRgEXoVcgUfQt+xVvnKdyItgHMz0
Iq4cQsEwbsONTLizBuBwuLj7e6PzHL+wiYg/RYvNKqHtucugh+zTzBQ8Kud/eV5/YslEeN7nhxVG
DB3gG7C8msoQtvuGD5XkKPD3/6jQ59UyPmnyrUDdyp9iW6AujSoH9ryF2vyMhFwf1ZuJ0ujYBMoL
Sg6RsQkTxA06DBAF/W5AAW2dWYfOsT/FBGtcT/tSM0zCngeHZRene9coUxkET08Bu7XahUC7rkW7
quNmh7MImgJIs08Bcs7oIiK4tEWtuqKyAtxwVFVk2g9XCAO9kO8WXfWMEoZpvTW0chs99RqbLNda
2TVC6CBoaiJtujkITfY4h9iiXSleRs1YXXeW0cZ8a/pd3HI82NNRNpGVWRHN/tV3eeqW7azryrVW
ItBzgUeIh/7knNSkcJ0/wf7ixGmEsJGPMOhaRXsVaSItj36UYa0o+9259xWxGpJysDzIpsDWeraj
4bfYeDPW9WIIkprnDOQ+1Lf3hIOWjmAkOHftroLfXSzZMnTkCbU0dOHFsRgNL/mpHFnT8ILIsCwZ
vIbO05JfZDl8VhtfFDTahNNwPT4m8vM0D0BAtAX2/of68uDr7XN2++i+i8qfLteZsPBA0QOPwqLX
0d8Pfy3a0raK3nQShgdqvDJzwCQbzeT6iwF3txImmtQEH7rwzE8crdDLPwJhbvZ6fQ/PNf3gRZgt
m55rluOvBEnuVI8m+Rb/YlGDsMsD9VrExhx/ZNe9weRkFrUmhs4zZ6/uCBbMPa6+UQDAggJOVimS
MzkSqAFmhX3hQ87wV2VVloj87iJ2YnKJarail3IFPbuaEC5HUO+yQAdnH+mQVN+n2hVbno2KHq2G
GQlgfYoCI0JAqCWwaLZmEVsCkpE1NTtW/cg27AhryxQ8RnvozyMX7PKtp8Zk05WB04L59MeM5F22
KzmLlR9KzQfayLq2qYmzaDZViGR+yg439cxnXNjU5nhC1FQf+umDOX+yVJwVFau4og2BFCFvVm7p
w+O3sHUJpBZAPJI61q5NU1p52IfKE94nK5Atij8Ved9tZ4RRUIZ6J2svQQHA345WxbZ1J6CG8I1R
GRZVb9JSJKNcj4z6R7xERUnWp45Z0befkcz/qkUXREoy81shyH4e9UVGsVuaVKAcTfAs0MjlVaeD
/tCm4tN22oemDITyewQ4tsW/s4ERLKeNE8u9+BZeURaNCtFuokmeQPB0B/AeN3DeIfsgGg5aGYUS
vtE3YjzAwlWzzKZ2P+1bvoT+4ZBSZ3kNSqiQDk4eb6SjInhBCHxdztkVxmsNVeS5GCk5n/nQLlxF
4NkFN1tliy59a+YVKbvM56bFXj5/zY/13LdyfUdQ0/2+wU3NjL9gjtW1vwxL2+G84BV5bbAc0yua
xQ6QHoJfVH4N4XjgToDd0GsQHW2BFrKRQB04qV6jitep3jofMzjtttds1y4LQC6rAxmwvPWcJBTl
DKZB5jssjur4CDBCL9tutQ9CnKum+muKkMjN80KZkFLChc5WOArC3+H28tjBy1PFsL47eVyYTfMW
IHv9tVS31OJloKGvEG2X+NJOxcQFfS8aSehBESe7qduYKrijmdKtIaZSXqFm6JCNPjZGAoB8S46+
absvypC/cp8zlPtgC9l44VNM12vdrE69XlCwD3E4dtXTnIzAAjj5uHPDxFGBo82KoBBh68cEyeEI
3MCouHtzRGPipHTfviDYOQyYCcRxUB/snSUyGe/J8oVuL2F+tEfy1tbwaFZfLjNyqfpoJ1lQeJoU
CqndeD5wZKNlpeMTKROvMf+MwIzsE8u6ShK31XtefjXng92FJYOIyti1x/zfbiMMjq/ckwj8xOpa
7BVJJYJGosbp7pjENvFkZmw/+4IMzpvuJZ9WYoCdua6+zUFD8pGiIAHoUDFG4Q6m4oBFxCLivTWq
cX//2Hs0WwyMxvg8qiUjQef7OkFRYTtLtNcFWlwVdcix/4XtYbIOLq/GFB4yZKpsCFIEacASDT3M
87DmulctK96vjnJseuiq+egCBnxxMIhJzpAeCqxmik7OmFatjn04A4bkoEOa5p49TCGlbU9EzrD5
XIeZ+NxGb5BNQyvzDN3L7DxYVUp11x37VEHCe7FuqTuXxLuYZNAwPorHekZcVLsCEbKEamn3ko15
vv6214RJetE2FIeuQyuaJ7ZPfUatCCppxn+LEU/TXkz6+BaRlTLX1/UebFAdAmnb795Y2YagAKkD
1mRpYDYiE35x87jjjybnEhWIksn7/FWb2cUfBj7X7cN7Yizt+7Dq/6ulnH+s+2vfSGvFvcWsMRG0
NHhvoavsc95+A0KX2tJkxWdkp5DxRikevcChUwAC/Xin8L31b3LKuHRvkTIEktFSmDWt7n0xk0HC
J7RcN3lPZ7DZWi026x+z+YNKRXD91pNPXZrH8pUqreZE5VVZIuy2ktN42/K7QT+Ru50hH2fNAW/7
KXc4LCQM2t3Z0RTwWQHPoLfO2TZ1rizJGnXjN61iMtDIByOL3sQlEokc56nApWfKdjzifFO4QhpT
4sCH9EBN07kxL8T31wnVwA/ogUQbBhh3hVtLXqEoWrmyush8GrrVnDnMZN5wgpq+7lGk5ALFa8YK
UzV6eecenjtOTI14V4mG6NqWVpGMl5ktByFR0UksDMRTRv9u1c+HBsIbOOMSgZlBkpRsG7nC9LvI
x+eNoU0Y0ExbSy+Gdo5GQNLy+F5dpmCC9Ud7uYV+ly4IDx2SqXlcO/XiSSabCbxaJutOIx4WQznf
w4yjK6jBslV8rO99eu0FWPdumzP5g2Wu9wiWsBWZYLvoC2zHvVOmpwyR6fyND7xYWnf6K8F9IFAH
rnlPA2DFR2eIA4V33xQy+UWdDw6eLePEwVyAIxRAJhugyO/9j/fXEvchRZgkGq1CMI6OOicN9qBP
W32Mb9LHRPb/J49cwCcd6A5rldLYVKoUad5oZJzlmaj2UqovkPkGMed70u7lNhplXBUHkL+NWPgd
pbbObqDAiLxMQoj24Vd+nq9j2ZImZjpkN48zldabHR19G4FSrniVdMg5gqCcUBSTmBkoUwxauJbj
v+0HNapgWaN6KIz7pPUURx1w0cmsu+ECDq01HlbQ2A+2PW91W5huItwIZndgynyljXLRCcxbvMyL
rLb9g3r57BnqTcNOShhs8w4GCD+Q4BGRGILVcQQV3m7/MeW2z7whXbvRnvDvEnGf+0dZz0axifgs
J6Mpj2AcxkmvciJeij8PngjEwqe1BmpocjXL11sFzUVBaIWkffRq1W9mxStHUyJBTjJ4s0pFsEzy
0MmLpgyt1UPJfcPU/AWvWZSeY4/HtJa/fSP7Zu3AHNIR+6oQEzhJFWFN04mGDfRqteeCRK3C0GAF
CKThznlQn5suraHQclyI/GoLYmPEO00b06V9tI4nAsamRTyQNRNbgeJFy2/yVCr6s22mahZetdAZ
a0YBX3aNQuexTVB0bBg26t2f9jAs+imZgfUlBywD8d+7QTtwu2wlfTyO047PhgDfRNl/DflQ5cDT
C56RSStk+iJ5xqdKY/3AoVuvTWC18qUCTR4vRFVmyX3aCCTCG4b85UVw1+R9ZuRBIbQtMG+i+SGQ
Tb/fqEaU1hztjbPBKyaTMK2WrGVH7oHmzGXGA5AlKL9zsRRztH2pJBcow3MHsldJ9256MWmWSSb4
pjNTKS0aiiGzSeyOMUyFqpc3ZeS3HkXIII4uijx3ZkAZ9Tha3GhTNkuxXGAQektb91F1zZAIYGpS
me4rZUkW3ASGRnTNMldelZnk3OV3BCAC05Gzq3p6YU8UUjt5qBstl1tobGKCUab6/1F7cUTiKOrP
X59L7RpJ9Qex5sWrPMhrYrrlJFQDBR/Tz1LyGZRnsgPRqk4p4ziLK0DXsWv61xDchyYxspKu0+kK
KS7PISYAiceXUJT1QzvLEWfLoTFm3yNl/3LzslMHwb0X9G3Dg9ZBqrl3KE5zNqM0kI6nZlrzmj/J
H5Y5XtEOkrd1djFYOckIYeIEklMSjYiT5gUB8iO0jPGoe8KV3hqxTYMBAARZ1hnSgtCwtqUG4MN9
yTSWHywW9j7rFNdaq5biWkfyqhlkLvH9klpYcnscPJllEobnWNzO+l/qVTjUd4J6KqL8vqP+7fF6
tCGu+/mtTP72U2htGwybhnH6PCV0Q8fOcgBi0UvReZZShFXazRshxjGO7MvVfQEXnhiZ7OzjZsJR
GH/6ZEDh4Z2RreGe2HKdObKmY58lTfBsk7kkxkPJa31eMAJUCoMxOMNQdT+zJlGHR+dfJuSJRhoJ
fShb1b/bGZsXZaqHWH13r2B2Kue27zabSH6AUb0WQsfp+crrUsi/Zg8ZGIagVMgrC42iP/5+uoAg
FQcFvZggZhuAatQJsAknI+VxMhIVO/mZOBMDQ0EWpHTh0YagbIgU31fwFGKgUPCtu4ReKVbkf70u
wWsjYz03jWAR2PZNcecJrGWTKO+w/6+kmASJIGAQwDi++TyotiTZ/j874kuSoTXP2m8wwQXHebqE
YN2w1yUWa3cjim9f3sBv7rmX2Yil87VP1qjAd7SFNART8lXabXx7olnyvn5jqe4Vg1KUrqv5Ff/2
YmgUB9iIuZaZdYqGvcMDDLkLRQbvhSoG0lc3pM+1EVGb9lqZP9x+4mSBa2bHGYflCELshqDTYKBQ
9FzrCKmT682k2J8qR98TcOMwM7FNSyDNY9C6xFsUFD8lA370X40gaP2cqdPULqM6ER/r1U9WNGIr
BuO1exH9onillnF1lEh0R8L3wJMC78XCs/ZIZezes+NeR7PBg7M3+MK7xNUTfBTr7ztDB1lH4dna
wJ1RiCTlG0FQOjRijzJrAKaLW89PKT8Hht9pd9tB0rI+4NDV15e9xGDefWUz34tzzjyQbmJ9Szcd
4R1JAxyt0b1qQ6kJVU5ooFaudu2XimWvT/wC0Pt+hVIMIYZE1HaiieL7chIPsJtKTWmu58Ws9/ZQ
dlovfKpYD0e7OD2SQm5kSYKWOey+D/1Yd9/jFSSYIbzlJe90DAMqR7yuDIe43CNt8xIz+XyrIY/D
RC+lr2McP593AsBOO6fDW/Da9xFGIpAjcwT3jbPEX0G/FrRSjKaFkPucnsWvaOMTLTM+9xdjHLGd
T2iDehpWYwtzLsUAGaGX39l//Yp5tYtufY3uuyupLUMf4uP0yzDLc5QBr17JDmVUmFeDllaauKuL
sh6iHyzToHMVIq61z69V/KvSv6JWRULlx8Cf4OkS3lggAvwvZ6ih1wyh3X8JU/ciVJeTlORG7yQJ
qmHcHg2Wih0YI6AL2nHWDI2FGFBDjL8t5B4SxcBbmuBBKoG9Bln6Ff3mHy5Wo5QuZV1HjwxeygEH
DjUFvcf3vnTKND22UF0Y1DTDs9WIjl9qZpxXE4imoWCml8obiV0bJMKEa9uqaWV97bNxpTroi68E
rq2jqScs8B/hKAZymFrRlTqOhb9eeycDE7gc61lPu5tuYxBF1YZt8+TGo0mpnqJT0uMRKNlTbU78
gsUtxwVQOcYE77jd2hwkqnlO+j6HdI4yAbXPfHffVMilwg0FykhcomddjwzosxsLrI5yyRkEXF9L
p6rwPtPMkznN70wkGigA3whMG5fQKvAGgtf8OS/hz0GuWV08Fepiv7our1Ar6tv49k1RyFZynfUW
51DnkwQDWI6WPqinOsA97AzwTvwcN39nin3Du3xZgFFLrHNYaXd17YDR74wL9NN1Iz/x+GWGCwjz
4pdTVXl9XU6OjTRqDvAbOPhnqYv3LWnF0YGN2YX6MD0PSKNvPzB6VbMwsCdcioGGH8zbPiTzaWWV
UOWLaoz2gamamVbU/K3HOIWZqg4MjUIXy0UlD/wu0kW09Cz0YwRI873KI7bK/oVkiOLdk0zCpWaE
ORpd0VH31q4+oHAh5FfqMtgDVgpWUMkVzMGU8TrZMgNuKn1ak4cArd3Kf2fRqUrZChlpuSdUR2tm
wLElP5yBQOTOJIrNVomk/cu6mfcyZFTTzebmwG8UytxoDzCLUyfS8S5DXcysb/Fz9/i0t71kGbBw
pDh+dBmiuRjBT4K2b+uc8TxiYiZRxpl4ixy17ZQLzseB4aiUrMGpKfiiuDJArdzdcd3Evx4dexcO
bbRtMDDAJMTgKwmM+j3oz3LF4ic4Td+ju3ecaIAQteyRy7BsVIrO2q2pFiczOq9I8aNpKPCd0KkI
Pvgs3mu9lU5WxTjENzmwXEuWbwQUtQU8UvAIRRAOMUs9FJuXAEl+qXqj73EK7wtr9LeguT/kkSSI
8smOOPmHkvJRnLqHPpsFVIDUSFDOPhOyvcmY2dEEV0MDW1JWJac/EPhO0uQzbcVAi+lNQyd2M2Hu
D/QRw2DQzXAxeBvec1GBYlZe43HX3yGzON88Db06CiPpnB9Z02y8hJiqS9mCs1ZuZgpmtszO2mxU
nKUHLg+JV3TWavnzKGfpvRpkevzVxE3j83gcuZi+1eZizT1qmDAnPEWSLY9BC7l+Y4M3QPhG1i9k
HqwSYoCRCF87qsbVqA+HtphYyWwzQAmsPQg7i54dmGBvjFH/aKUlBgWLGHPMPC1+h67nR3KoB/WS
HZbnJmaVqOWgB1LHJ6xASGVbBCUP8FsBcb6+E3+qaH2YDybrVuF1Pzmw7z8CiBj0i/Q7n8y29ktk
0o2+41gf5rfrwvEkJw6Ochre8yxRbzG9C46SugvACg2p9lf4r+Ek0qaJ7FhR1sZZtXh6UggG915F
LfH2+o8JmmQn3VOow0Se6A1cmVXcc0zoaqaRPJTbCn7Ivvur0ZdPUgLWQ3HcgiPy2DKDcUqZBtsl
X5gxUInQWrLJdM71k5t4BIgvAKyB/HGkGFsgZAlChMEOUWK4mEaYxpRswYLdPZ5onlZeKhUF2zEz
OWuEVfgzDQV6MM7vNerLSIpn+6I6ywhjCXkJlpJYb4GU/W62I5BkQ9c5AMFx2+72hOP/sh7jcLf/
f0OCvcuU756V88N87O7b6qfZZthAiil2lm0A8XFMRAYrFUFDWpFXd+kPG/QIlLZuOMYTP55HBRh5
UfAuN9mzSCc70hG3YLCwfkSdjFF2RB3vUkYbWYWnVRG4F78ANMXOMy/rX4266yiVNyDkBVkUYVdx
WZzXSLHTjUM/f+m3iA263k3Cw25TfctT9+l0d6WgrHAjvnQ3zYyCA0TITNaSwpX73TL7CFygtUMi
fixQC+yLHWmvZ3YkxVdH8bx4RyxWsnpj4GBHHYVZH78/fmx4e4Mb5KB80lELjQGbkT5kx75+RQiK
qExZS/GfbqtG4CPKToTZpsB17HnYBnJ1XVkqOcHTveNMAdXNRz5WVuszFxHwtKMitO+q+NHbqgxF
3xbFK+CMFG/4a9GciZ1uAYaiXtEjGbw019t3zODC6OxjUQIv4HG++uRbZaT6XWhatTQC61lMQIM/
2dz3wAWsBTWtGJpH7Cv78r7DVXP6bE+1s+kEr/HLdGWz3mT+C0rrDov5uR2cdedV7Z+48TV121yP
5OpjBXiHjzRXhteZISq5nlqUFl2fRbxncRZohq+60bVmqNhy1/kzBU+WizVT+g5qvzNRZECvDUe2
Hx2yn69S49hqVizZe5CaosgjnrVDbjy5ZLSLA+gJXZofbul/i01JPVVHpnFQvQ8tgwvlfIF/GjPa
W5/SfSyYHQHGh0/BX83oldzuaawE1AE62YBSvwK7J/vjFHvx7cteLV8WuAXtvWGgY3LRa2jLBCii
AVcgOL/yjY/J/0iBkSpok6t21uRWhb+gkS0OiFSPZ3A22Jkbm3IXCEXlIm9sm+weDw2+QU425xex
XZKUEjCKZQ86NJuKp82aVGReQye93K3LwqH3wuxsOddA+aSTry16qHhMbndUkzm3odqRHiZA1PTd
hieECqd+j//h30Y+Z7ZPhADNiSXhmOdO79smIRbnECAMsje0T+28H/eBBS67QHk5fHe7MOfSkbF1
ldl+Jvme7YyHMhxkeo3mGsjl1xr3cL2JiX1G4kJIi0lpDwRm3EVoqnBa8IR6AIOKsQzBgrR+RnkK
f8yiSAaBQUB6xKRBZo2Rfe0xq8FbKkmQzpUzx+rqsq4k7WCOIWsKwVKDtlsN1LnVzTSVLt/9gIsH
KnLkv5hkVaG4pG3gTU3H4we7ckvfc3o/sqzQXu3m5hLDkz2CagQYcbfQMTGLio0SBA43Cda4Uqmo
Iwv1NRGQHdqXcE92nnOtpqGt3gQhSTw0ouP/ss3fljL0NyHZh4vmMg/6AAmY36sDLahmKcSWrn9Z
rPrysL7SB2dEQ8OxgYNHo6/ffiE3a+shyPz65Och5GQM43pvER5CIfrC9A3Bvj3BggNt0szguOkq
QhjZXWI6UFO4F8K3GsHiCRwdmg6kZWzDtUjDRMLUp6gKyq1AgOgHqoMhqbATmtVkjleQmcgyaXEm
mLbMu+J4sWkl04lG2F9j8pUhznu9ZURyvKsQGZqdgMZZR3JlgT6CiWAmSoGGvv8chWIUtYmrM+ri
4/2Qx7hYIGxskemexBzPr4iTUm2s+lGoOFreoPuzbZHZ7UW/n3EWs47F5FVSOHuZRAXogy7SfD9j
Tjs0djFpC6hfnbqbq/x+kn1Ol88POma5Qv3jwgPXWpFU0sHOGSCaayiSJOhWAlcajzAiPar6fP+G
bLo4iq2GzVgotHESlnVdppmHBNdnFX8HCxHasIzYI+CPuSvqqnO1HQ6Axgx+54zA4TlXBVqXHg5R
NQx7BXTBtrbBkkp8ogcJ/69eIHbfQR0E1ftnnAmr1LWN+YaSINYGTaq0T1ijlNNqI+psU6UhY03b
2nmLU4LrE53Yt7xTUORHtVFqu74PoAuuyXPvTwO3iualKkl6R3xePx5GrgXMioh35Rx7Q1P3f3Ut
LY9jr1MF9pqyXchkyT5MIlGok8phiUqH/7Em3xrMUd4mC0dMKIYyQfDzEb4NbNryxnY25/XyjV5U
RLTGDSyB/vLwyEdaN3MKLCEc3k8cj7K0y0hNkZTXip7X61wB2qmx2QlXZqwTJw/3sS9QFvC11Eod
f+ubRsxV+pVhl2q3dGIURxR0b9r9sjRvCvqL/8MKcOijhaC6KorHgr6tUU5wiau4W3zbIZL2ZEJn
/M3I5C+Q1dDnsxO+KawvixGkPjm51XhahgRYpREDJpFfPzKbHeyzZ/olVEs89lUdh48QStYFgjTp
xqTsvEgQbzXokMgLgb3ZGfhiNjbSEkVQ/TE0jQ70liLGTqC+yG7Cr1TL1ZaoDtg0fZku+t7BqklK
BKe5TXFH+IEJZuz1LYtj1vLjCc1bC3aEPR3sm5mITWyUKg8DK9aMO1NcQFWrwWkWmQyPrJqyPByJ
bSIwQb162pmA1qm6tNLKgzy0DAhvsW4taZ+92l787rTFSI0UimcYOqTe9dTSkzdbtTggmxLdPdGi
jfGihFoOgM3ObhMz/9HJE8XzxrgKVHVR2FcVQHsgRn4YzGFzeeqYemj5A0V/phdcpZLG8RVPTxIN
gZmgbiQv1aL3Yof/dTKReWTFca1dphI5U2EC9lLtT0ffE6ZQ9tdUJPxO6b9HwUMKN2KXntI0Oslj
BnY2lZh8xK4XKWNz7DqnJ3gN0+BFE1At39F4cbTPQgYdqEnc+P07xlnqmR0f8O/MbeYx4GKzflYR
O7aV4ADLf++/H/E7cfpgVazWF1bO40oPdahAFn9BPlGm3isYMPr7ZYOdl/dNfP78h3TXtPeLy6bS
EqxElIvzz4w3cOda9Qn1KzoI5qm0xpX9g2grLhZ3muToUle8Mbrq236iGlHm2d4YtyS3p02COxp1
Fxgad8+js5Abc6m/1VyYM5T5QT/FMQ6gjBjHMrqBrVCmn6m4Ks8YZq2mVcJXhwByZpkiR13HeDr7
iVOOAv6RiQnXySLf+zhloT/I8OoaczBeUWHiX/hGtSxv1X6iVudusG4C+5hdEDVY51ao4v8/cU/k
5jv+UtCJqR7j4mhB9m5lb3sh6+LSDSGqYtrg1b8jJg6k9Ylfds3VXP7+ZV9bmPp4MbDng3n3U/kx
Ljgb0gAjuj0iE5x2WG/bB0DTW6DSLYyls0nfHhiudhetAlFtYbOcJMUorm7DYb7GE4h7jKhXZucF
NsnuiCWNjq3nkPmFn7hk+oQ9gF0O51BBOaeio0In4v4PjS9ODSnnlbEQCcEj7o3heUy2Fkv5q5uH
mSt6m9456xDBKSvOT8R8jRruUbnt7CixiHB8sozBDoFIHJD+LEVkVAEFZTk5DDQugXDpJcbL09BP
lSyOYxwfYxqGa/AZYfQ1gPpNsTQHu/ef9rZ7drpv3YlmBc/QvQHSInPTyXP9VeKY/+/Y1QgR0VWU
kMVz/Kj7KiUCBPcnIMd7DAUPQm7mwP9Esq/mqCJOdzBqGNdBqHWgKJpZL0BY4umEzjhmAjuSCV4R
oNSbw1zSrGZGfwti0E0pzztrmlB12okY7F1rCczeIGxRmwHyuEpfxI3VDBwk3xkVvvpf1xKBaVQc
lgsXsu+y6Aup9L2uMg6uvQVHuuPbPYuXEetUrpsGAj7SP0QMZyNZuiPoAApDtFqTiwNIk/1HCZb0
oYzxdZph03HRXcSsPqXH5j9lv6MQGO6B9Svl56vfEGr+8UH2ic0ZzX0+ZtpyG3HcpZPqltb6HMwF
PFC1H13faWIGdNbsfNdD5cyFGIlDY5ga5sAHAWNMgmonKY+f04NxYtzKRGFH2NfaA5nPHbIiKFfz
HN+iiJrrnoXM3yR/EELBiL2qtskggib3i7B8Sd2OAynb7tgu/oDWxWdZirWUpse+820Wd+/2RVIs
pP5JX+4i1RGmmZsohzX3Zx6rGqMs2kt96YyWyeH5bh+eWXehtx4yfpY0ZrzkdE+MQqaboAcrEkBU
KM+NXKdjtVBOV7H24Z33nAG2CgSRazfeg0sJ/m/6EqT9LouK0lZnpXv5m8V5Dy8CQeMStkDbxn5V
J3N7DuFoLZ2x7mD4rzvoRd03fgqRT869FVSV7kKpSTz5Nk3BLAX1i74hLlNb4Z8qIUZkGYi1dHfs
kdhVLoMzSwz4BHI87zSJJIOJFGoQjZMs8tfuPJXnxwneLGR4mKFFSyTqS2uJWN3Qp26/DbBwMJOs
flD9mRu9tfsrpajwtCOazNJLvCcd2laF5a9esMk4frWPY++ggcLWd94w4fznkfrG2tiq/PrVmA8Z
x5cJye3U5RUe80abjNw2p7eI5OpBtDcYTw/D2M6yHCPaFqMwP7WhbgOlRQFdBqOOp8GjWaTykp4J
/h5X8gN/X4cEG+kOTSl4wRBYbVN9BEdlT2PGCWyEOVUaHuFMKYQ/fhzaDJdlZQMOXPPBiXkEuBRu
qse+iwVHgGwrKqUh1lbog9IzP1d1dygImSFG1zLe+sQj2dE73iQ7QcQ7mUe0a4ulWFISt/iGG16P
MaAlhWzBwDijbVMVZWO6NC4+pVUvJvqZ1LPbg3tl29zUmoOnyGWsrlicRHabndFdXWn/ZWpR8wDv
c7cvUDs+9npw7fEuKhl5cS5p02M3nJOP6b+M+o/h1z7OZ6T9mInMqE32mqTa0Isq+ZiQ8ADJ35ZF
U+5jhjITYi7kVM+Qcv1brcJA2Lr9IOslhZgQstMYPkZg6O0Edbp9iMFTBLwOp5FKlSmGyP8QedgJ
nL/bo4R1LehVgIdPEYOAPifufbf7cOHG3Ij1b6bPuTuZuLAxi+7IRMc38XRZt/CU+1ZTkzzkYaXk
rd5JipPd8VBOkJWMPV7wdIPEB4ICpXPR6kjp7/hmf+xtfKgfeqPVdPbw8ghaMYE5zswkJASN81ZL
YU9Eh+i5bnLs24bRO6orhQiANgp1LuztWscow4y6B77BQ9FAPnJcBCY9UrSslOtmVsWen7bbDGhk
YvFNNk2CdAsns9n8MiFGIAFpE4tLlcYr26UU5veYjU0BV21g32f7qOCIgpg80p79Pd4+0rN7srew
z0Cye5qHdAFarf4+BQIo7GilRRQ8w5vAiiFKrM/YhH/orXbtY3euis9mSM/W5W2CaU9SrX8lCmMD
VRO6ZMN5P9mP3Y2lXgoigYd94Yhe4S626a1a2m3LIVW01HYOsEjdqc5/eegUT9EST7oP9g2DwQNB
6oMf9YlmzIBLlk3g2jf4lmcMYcq3s4rW24+CyQ8W40FkyYbulkKl0/clbXA3XjQlxGqVm+uynsYH
mhHCaaHK3oGMW0udB7ZQe8YIqpbB1PUOYidi6lmr6DQU88KrIJJ1NRsqdQe4cZFqC11JOFHRmx6M
CVrdw8FfmaOk40MNhA2+P57GGJ5je65Ap1vF80oNT+kYpXf1ZDu3AUydbqYVI+hJfaZ4w0kAa+az
kE6UCQWf19bhzp/P6NkbvCGCNWeeNsQSHxZlD0ACwDkndRArLBwmSw7DTEvbA287mzrgsE3rWU5Q
pae0VXXhKkJa8pkmAhSEMFj8j8uR4b98uzHBsze6BS+527E60XWmtqB90gaHAY1jcIIB3uWB1ji3
VarFzVm+E3opRkCz/RC0OhyEWCyVypmFDVqr0mDZjojnv63vy0hTDs/5wAA8sXGvNxE7mBnD2QVv
1msusIcPB/KY323uIVK2bAH90+x1rKkKwUTOnTQiUy/Q3vWs0muUGFZVce7WIg3o/JUGLJa2QOvU
hL4IW4SrRmUuF/+oyAEbQQKc2Pzy6civKBEdqiwSHzEnHXSzby05VNqUCEyH1RHKR1RIJ84Km/JC
E9t3muxP6ROtXSDwLrHuBBFNkuBu3eZJBSUVK2odnkyphY6XcjKSuXikBTPCs99YC+87wwZsZE3W
bT5zFEWRIJ1xrOivOqxiIUMrE6hMv59eK0NUUnlXkN1B5u2Z0DO5qiQgi4iCWvvrGIF8AZ/WySFj
F+hg/EDI+ksxYUsO0qwEjiz53qc41S/kEiOTrBjBMVxXWC9TVc7Hz2yAQwzgUXS5KxUE/zl/Ifek
EW/PlwIka6g1eijDqgCGvj8m+k+2nImDFdvLbMPLt/21+aPCTyQtJKG+h9JX5yB1tOCftY3GoRCY
6DDbO6riaoiSyFbridKTSRu8KQS/Xv8SdlMKlJ9PrTMnFzm/m8TI3MEs0BtDHkA0Vevg/6lARMoi
pm7dHPNE4ubsF8AC1LEWHpagZEu0Naq7+cxRLOAd4acvYPYTfpwktSHhLNn9SHMdPgdmUx4Hxd42
PRyyoQGPsVNrejZzf49VwJUrZ1Dc29syMZCYjZKZA+pFjJiDAVeOra1ScsZR4Q31ZiLNXdkuAgg0
CAQyc43JtdilvbAaagWB3mzM7CnrSy+6hqylVFlT2ILtSnc3vo5J1Bwrrcoi6mlg7bxzqNmsNAIp
wDZ4MLYd30nql19hhCd6Cgj4Q3KdaHt4e13stLU2JFFpkCrZazZbCOjxq7E4EqTUXqHP6AT4SxVD
EXAcuPW373QCtv3Z3iX4rz3N6h5RZSWJsoxVtU18GNAWQ4GJwm76Bk1JvlKFnZMqY1aHWDDs83dV
OSHy0qbvpBdIQaV/bZJAwrENKZT15TLAPOIzrXrjU83XujtasE57qFfm4NCmiL/IkMegXQ5N/Esm
OwEVTUoKfoxfKL+43qwDUFTDqXDjw7tiHyBMYuXHBcUI1+pL9HkLq7sQreYN5Lggo6EOj/pnBue6
vxu37HIgwPKFxktkKp9CloYB12IQf4F+3+mUOpoH2uyO3IH8Y5NNxgYvFZ+svuEjh2GIWwg2fNJY
pyzuN40BWxR7u51TCbTALi+xmeXK4FBsDSK65WdvQ6r06ak6EnwJxq4KcX5zd/bR6STEYyMGnsty
RP1BjHEnctFhBn4dzl/GFV04JyP5U2LLlQFryw8bG/CHjjRPgMvLYNxVLuXJPzM8AyajTXg6LVdL
wJdDn8xrthrtZIhOQbML+LjPXoTusD7cXHLWreo/z96Hq3U3BeIcT9X8nBia8pwyfUr2Q9jl+uKb
OTzOpF2oNvCP8IQqaoaILmGx69fXZs2yUPzH2IQpUh+4/EnQChz0Ms3SyZzb7gksDXOw8Bi1yG9Z
apW9oOlvZ+6Xsa40AjFxT8EwJXqroo7524c6ego/iLkG76DYqAqFZn4Gql/3cC3QzXq4BfjFIheZ
3tFM1u0ICatl7iQ1GweAdIAO+UvTx0EkbkuIN7ouHUPMEhyjSO2EQEnUmp1EobExPiH28nXrBiGe
tWKKhL2l38lANi79/TNOkY13Nc3ZRIr5IwQRiyysOGL2WGrhqzRxiygFGvKWvB7PSqwTntKVVOrw
0MmuXBFHDAL4AQWyVy2MVA335WAWgP8LKZ+KnBzWnQRFdN5AMdnLzIx4KXDE+OlaOLVwKumv0k/X
BVnT9X5OQnIhGYisVl3Ecl0IGA1kJvbp2qBJGN3eZ7Jhjgd9jEk0bkd90vF9yTh0lIV+42eR4Jp+
RN7UZMuvipIwqUeMwIIEvWGP3m0lU/c2BNxdrZ7qDYfYXGq0MzQP0Kzu3/xEgNKQWLJbLKhsGKG5
cmk3ErfSHO0QaAAxvHi5nFsVmdRsjhNDM3lH2qPgRNyZ3ZfKiaXMug9uBMfhHCl4uCDXNd8RZdKL
UH1nlYYpnL09P2geAbqp6H2/CsgPRLRjlpeJz2xZMIwC5Nm2XMBxE3RPwvuLDkaAfoTiO2lv0PXA
p1iOL/voGWw+L/IWWsaRx5gq5J948NejYcbGrHWy8dH3NC/HL7DWt2uZkuXjlI5hi5NoTVdvTLT4
Ss5w6ezVOq5m7GVy5lUmcfXhqXnXBahmJ4cNAnFL6r1f+d6Kq87XtAhOD2QCN/p4TXCJIUTBxVqJ
9I6XQrA2nqR1KNUEZaGc7G4dFz4JSOgY8Dpu1qcoY9ecW3lJc2wXF1zXDcVTLzEktmSmZqYMcGGJ
O3qlOLoTxFnqKjx9xYlXNzpiTmT/iEgj39zj0MJfheCPDhlRg0Jl8wP24TSTgry9cOctiADTbr/P
j+lgx26KnqfeRZUEprTl0yd5DJl8nLyA5Wz/R78L1AzUmA2dMLRI6iSglG34ynDBALP+o6CVvVg6
54pTiXK7aJaM7GpMYfNxpg1iC/7gNNjW8cw3Z/2EpFrorBmn9oXIX7dpPnlZ9nZhbYDlCxaq/fCp
lUgohntYRkspMzW9RttXmJAv1X/OXnfnBtsdZHsABX++tUdwmoQz1LLlhDCpLCBHxnfUDQPQNA5r
Qa3PAeWiN2CqqsbbCK6C0f4Wno2Als4f1flUWCYvl4VjejruwkY5yxwQ+GBGqLZFVuevgjqsKDzs
DxL464zdEw3LW0oONleMHeDTJZzBz/aFOfQTclXZHDYFU8859EC2CyS35qs92wXkclviJ1EK3oal
bqnYweDy17zhZu6nJWGB2eOwvBucnM4btbJl/02bediaY2dsfnu9Me6rAobaorsyg1OyA8b9EsQv
v+AIDIo9p/pJtEiWGmrzEo1NY5q66suwYJdOwt+QEkNO3c9TlCpKidaPLXhJnlhyRt1mlBQ/KMTM
HQOwckttefJe12O/7orcBeAnKuQ0rbpdg3JAwAXcZ2vmWMZ3fnjsiFVOkKhURe1fRZsjWU2jUIxc
9yJFH6Grogy4SiAFszoQiN9PPCSmuxdO94WajtUUgF1KAzUf/kZTrU+ucEJR7+VEJH4mx9QCc60j
04G4z4oAu2JIutPi9KogzamvvamPas2OWFr4Svop9SpuJCFmPKroXE7+N7byA+cb0PxBnj+9IHzL
4DxDxSWDaNSaptTQ7JWMpo1BZk2uOEXj6wtcAYp4+/VTtofJ2epPYyLvIVhzcUBPKiCtYTgBS6RQ
GtkckmVjYVWXiHoCI3gfeOrBAK10Y6kgjRxZ/0qPAe5XCxsoo5AcgKkwIeddLHV3x3rShL48lBfU
l05pLuuhK/uC94IjBm7x6UJ4yVDHp892PH5GOz6XRuIH4u51X9WqMROGnC+Frgt0VxOWoFsGqP/e
nREvN2FNlh5JXM3jviqhr9mM5MfyvPETziYz5O9VqEaSZBbG5xOxCIQDvipeK/kwV58LSq5Hieh1
jLPJoM6XuC6ggOh5TAJpAJre9w23C9+kUDs3TbgWoCeQyAg/if0QGeouwa4tMb+28WhUn59IDbb2
BVJ7nCoItKcDwGMFTHmvbDBJlRsrpkch7TV3tqjz1XPTDMYAvs3VMnQNUKitLvu2pbg3x5FmydVk
MamDC7ozPvfLL1yPXEpH7jVHZfNmdiASkbmN/Ag2Dhs0gv+3LPvEEA4yx6oty3RqWHcJNwV3Pfd7
XuFwcQYeLWzaFb/DffBnTLIqFDWAIOzYzrCca7AG7JU27QXnRv3bXAI4C8jIdy70UIJ9xpfUfZKU
e//WUTtzNBhKJcwpZh5NdzI5bpb1cFJc2AzJ/5jkD3q65UDyNXwHqbX8klGVSeFCF7UJbg6t0vlr
p5xCuumwD2Q/eVVUFPBubJnoMp3hN6G/w9kRFWE7Hhf/K6ZxzH3NJAJY5KQAXGCTi0yy6xyG/TqF
iU0MSuIIV5f3S4V6V5boIf7QGuFSd/Ahd7lokR4chWHnnOl4AUOVI0kimK8bLRqr+3jYw3K5Kqzt
QepRk5b5Ezrki3MUjC93t+c5//83f/45yPKaddxXdU2ls3sZ9d475vDePgqQoRenwNFu5HZ0NniR
VUN4C0aiUgIXoEEkxrMYdsA43MUXn1KNbcd/tsjpGy8heQ0HOEXREz743FpzW/ShbZjMx3fPSd3l
gg3erJHuf6QB7b+DzBO+o1nko4hekbr9GrY+T8MRxa1z8DXCt09ezcC2RsdpxPeaQxKPN1XrPFcA
7ohhzowAb+IxxmzpanNq8cCFIcJcY9QQnZYLCtlMtW1MAimq2r/Z4F3ovl+AQ/ix5Tdksy+E7zEP
uU6y69TiIPeAXTVslvyczJbkYPRyp9lVcoQeWwRMAnI+VsUvKZl7001i+P67+qjwyYH4ZLTE1Lpd
6P+7e0LhJUlJUxS6ouWyiBs5aRSLjdM+rBNMieYq6JyqjbHECGftVNW+q0k+Hw6Rxe+mct3/Jw+r
wLMnlj80oB3lb3wGH1ZbSdc9wkBKpNHAzyZJdD8OnhfcbTMGyG08s7e9sHCQy3NgfClILet2YkOZ
+ym2ba4YC4Ngl6b1zwWLf39N0k1J6Wm8ElXMdo6iNxJcH6clUxeWZFNXt2aRwlvOm4jACoh5IC8j
UgXvkmyfHLPM+29qD+lfmkVX3RIEf1pXoqYFx8CXjkfPkWHk0YNILEgGS/aAq1agVk7O4Mjowpe6
sTQGMd5gWzpAGUqb5hnU5cq7PT7iVVBfFLCG9DgXYVKA5mCvoe44apA1KgMzn36gBGmxc2Yt1grU
qBSKcXuJ5UC5WbvBGT4YXSFS3KhT2Zbilniq5FABHtRcwRD1jYcwu0x+02KO357o5X7R1j/4qoYA
dhpvxZZY1zt7fY0gvTIbbSdeQTTaeByE0CQQV7TULmC2lY/rQcotwubwqjCa8BbgoNhAsQXSlVZl
GQGbm5T6jj1Is/HOIs+z4JA1hlxl3QEOEmeShnY1XuwF/3wM67A1ijSw9YHYN5zHxr3coQhNUnQ4
iZxemCNmPG0EKFjVzqrpibCKD7G6hMTd2fplJyENDI0vCYeeExMnLYetnOpmSTp4jkrxhAvHRETk
vlroGrIQpD2FoAbykCiWOqPyzRBWFPtG9KHBi/1H1jwh8+8rFO5KiBCJDMRXSzg3Ao6LQKDm1MOx
n0G1c+S3ru3HPMXEbot1pQ6E99AEGQrzUuEKVoNr9zSHPWytPRcCZhaH3uMtpMixZ9b5FnLgX/a0
4hhAQ+v/1MTKWq/i5mzA1TGmom7vbBtjVF/reaQYuPQohhwD2s9569KkOMuHnknIKk0E880iODfj
6rOePAFORX0S9eLdgrahgmhiwMKHYz2IJpdpblbr/XrRU4uOH6ydbBqjXvHGdVUof5nx0aiikRGd
J1kGw6/ZCl3SE3U1NAa7VK0wxSUCA9Nj4ed+JtHVdh1+y+O+I9nJz+TI/miPZMj/CE/ZukarNKKH
AJ/4+FCf6+BYe4zsZ9WYfq19kVo/tGU373i6D8wAxiUaNY9w3YDMj7dr/CfuV3QdCW0hpwPWLXRv
V/bBJtJTL3wwNhDawT/Yh/PyQVKtIG3qK7yKVqQrivrUaGrM1auU9uD9pHrwgex8jcLLmTkpTzGJ
g2zu4zBXZ7jY8QCvqgJbfQHmr9HEzjmpQDB7KkHK3kw0bIKBZIoG+nUHFf/bx371XrlOOAGafs/i
m6F3qY/nLkWp6d7au5FtMMCIIi4zPY5nkkejsyvixn5pjrWWQdXJkCJRkhxd7giIZr/MZog5G6Zl
ZcLzWpzYiJnCpZWKeM1JeSzBgvO0EC+lZ9pzEHCZkA/iOHUmMdoSSSjexuB2AYIDaLetISl5uU10
8iaJ6tcif+wUzxZL+dOqKlULHl/teHM2Hoz2EgF3tc3VL4BNF37pZv+LsFXpdEarysn70cPun6j7
POLWtY5jmzRl/9TLRQivnayQGtYKxSOsgOLRKKs53SMBeYOncpIYlsjcf1xiy4frwXELGP0IFn+/
LNqiWSwicibHtTbjiV+94K6pkj4YOfysPp7GWE/LS6LW8UiaLkowNWHYDMqCxlm1zno9yv/WXyLf
sg+xnw+SWN5v3wMjRbp6GKeE58Lw53mZWdFq0w6TqcCEN43nTtWAtOjdEqXDDcZPwnN9F9Zss/Si
JSrUvmgK9eMnIJVg/H6pH7aPT4wrhjr/qn/phDd2lZ1qEphL5HkTOBGFmYtX+hpNqZMRsUVdfku8
cduhCpHpM9HQ7MX7f6NF9/Rgvdo6rbqEhhAjgqh5s6mQa1C11W9OQaYdPYsbQi9uhU6VieOyDRdy
BQPtJBVthOB2+hkEMVUcjOXUwFYLoybmDYpoRo29CGQI8sa6CVe5iGsCZJ76Fe7dCBdNjkjzzZfD
XcvKC4HmyOyl9CFEF+Mi/F/vOIaQovZ/mk4T4/wEGXIqdP0TWpOSxQ4dwr+aI72fFwYmyGwUAcqZ
6AKuH74gp2EB/fFqKNzD/ab9PQwfVX/ImrNELwluvwL+ZAy8H5ZcrmwuQ151Iy/whtaDlXYPc9y+
r6WOA459Vz/U1m90/Qpv587tTvs7fpitLIa1CU/69zp77F6+OOMUWOv5ABewJEBOSZxW8lUZ/sxl
p1fepjOsqWY1YU5zePWfLJ2cJ0SkQRFfW2Aj6AyiyjrCE+3jJACdXB1lEWPkE5MDmMNZR/sDLKgg
NJ6r7Mj5O1oO1br5i17KfS4kU+bmkcoN9/j9rOEK87iuiMrCqh2i4xjSjHubX9TfcWP5a51A78sK
lMF2Yh3XTfcru/iML7WJdAIhdXxXvcxafofD3vOduYt/PEwBLyO+5lA4x85nclcG7iWynLonML/3
9mF+J4kv/6sklVZJVbQ4aaiQp8ce9mzhAY+V28W+7jN1/2cboZIoS2C7EtCzhFunqzUhBXHeZLDB
LLcL5mVLXRYYx0T44nxoPSHDBOxrwdWlNsHqlF6SY69n+HxnG+gr0CMFZW0hFyT5wqx9Fb29H3yc
YkizU47Ph5LU0GHWO3x6+TAOaSNOHkxGSVMqatT41DA5sranTc8wX7/onakE0O7U3q+DC0mYjbdu
kfNeWh7eisfeogUp2glrMpnEOuOLG/RLs15Kct4250jysPGqcerIwn3YBuVl1+di6Kyl7KTCughX
jcSc5EctDCnAE2FaqLp6xs+pzvza6Jret3c6c2t1MdInHsjiYG8w+t94sLvGeDXIcdkMAeIue+X4
2naLDsL6eA5bymltHVSaC1YTBaNcE0XI8xQpY1EukFow6r/bRNFQaGjn1SJ46LUfjHbdOGfS5Me5
HEgjramq6miEhpAtcztw1O8hi8QkcREKPEq9ujJ34HzzVUuN64Nnyu2bWhmgf1VnMOFub28cz++s
g85ZBLQ0XZ4fLJd3n0kDphQteRzgI6QQn4LeZnhL6oa8EmdlVy86+lLIpHcypjui+bHw88KYlOA7
HvgN0inyduNa7cqaWSqfXMrq5mn+CUTOcHppCRhLZc+IpCCzvmCMR5FFfSjNe0FEwRjbVz3F1n6n
XazckFRJQPao8nPiy6KeQOQLBaJp3aSwOs2Z588oENm245m9gnCTAaHbJscZZ7n8Tp94SQxwWioL
QoYLG/+DN8TP61dStp0s/AtXv8aWgwJHCqynL5eeZX6CNPBeYUOXW5GGpIKnicoR2a1jZa6y/+Ow
hYiEjJ/JzkDcZUpMPPxBAZ5XLXithr/E8WPLnXGhfttWPxenOJrQGH8wowPuzVcGX0R8tIkIUahy
+flKoFM/ehStiPBOVUGP1wW4zBCKIZXMdfYUQ7EfsIdiwhFxoMuap3fceBGeaZQPmq4PrQLA8hHd
dE5jCZlIyuMqJkBtZv0XdekRtwntOzC5+cPBE+OwyYDXXCYcT41PNoTOwch7tGnyhHqA1tmuy383
P2+mEToc4f3QpT281AWRZV5C5vucCJr7XwawKhSI3at9+dbekZd27yY7KvsLqkz4UNTF0TniWbEJ
XijZ9OTixUw1mBc7Xb7ChLPkErGmy8ntLLgmO4lVEaD41SRm0Z3WSMERTSjDHSAkgK6C7QT+UW9v
FM+mbAB+eJvsxmNtINawGcoFDODkiaKmDhhqT5rIGwikmXbZcfK534WBH5gxC4fSR9w+AEYHss1w
7qwz4xvcPxNKXiVDYZRjnLlDJLH09j4+kPiCLb489PFpWtxu9sgNG7LPQjeNhD1q5YHS0dQe5dTz
CHtKBtWmZUAsYj3JmIAQFbwKaynPFSWS63fBuvGxNlMkASYUe6k+cSuE8oNMka+r6HXJ9+5sxiMD
mJQHkfSuaBuab9Oq5qrv6PsNjkxXWGXC3VSV5cl78uOyE0nVPwgJKWpJq1I/udya7+J21JHOOCsk
YJHxuVGMRWKYaqlVhp5RJNZtgxwsTDRklM/ze3oY4yQ75ZQbj+eaWLdLfBvNrFGUiR/++YADTmaI
IQv/hTYbYLtuzM5Sd2+hCCnaUWjCK71UcFe1/FgaFtTNfdmmhV86byFsYwhlaXwk73zxad9LlUiy
rPvFC/9VnaoWxBKu2Q5UaM1hQ5TBZXT644EwZvqjK1FmTXhfhui/O+8485cx6IBIB7PGhxzp3gBI
bCPRmRWKo8XkSN4szYovksp7gNqmSByZvtofXjB+9aGKU8nfk0Y4vnrWCc8N+TxkMgWg14B/4RGD
2Ih4z4CEdI1gT5Y3MBMMHgmdWbvsnfeKYo6RMgdrBJvMyyVMhSKPUU6SaB5lw3V7pnusPRJc6f6V
zJOja2KEsazFrlzBuvstfznfRi01xFMzRUBxPAgx42Mpg7nPfpLo/55Urn54FaVpL+VZe/xLlZIN
bJ2T66c5ifs45XalIQul60ciTpgpv307Z6xwCoK4SNayDfn4WPJltTJ/VnYBHPI4G7w3A3QOUAll
ESH4GJZnSFeOi4Af43uFl9G08S77ReJ6rJAzVUqV83Ed7K0r01VxrUb2EwoMIlx4YaKWzZJ8IXm7
aAuKetg/qTwXoN777fbspkkuHfR3qGp9dg85Ej65TwQ8TDUUoNJ2hmtKX6FhQeRQN4ZcG86CUQe9
+LO6sxUPYXbvC5/t+zdZl4Lw1tb5mq3uFZlXt2qSlCTOdBfrTgIzIhFc8YzT0M1QgN4PSaIlHMpo
9tDB2pjzz/e1fJXuBIk72N7QKhq5AAba3D9qw9p4dVMQhiSqnbcNaq0AkbGYAd6JRAwCqAgF09N3
vYYHjA4YF6qKmlylZQQKcTZU+NtyDfHrPQN5K23UTOcc59awYZNGdK/uyZSVVYcMWmk+5zvWcvKk
8j/YoQr9rMZ0MAViPNOPONv4yyKPeCT/IMdEmQn0ZvkQhoVefpB/uByOWXd0eiJyG2Gfflkjumy+
yLkg/aqG1ty73fFves0ZmiuLChtnCYhrv9F/WTQ/FUDW2h7x96lf/jd7fRt3ZdSRlxhZyPxgmjRh
Xs0AxqmaJut8JyqVLqwLclRNy7YqM1UvuEtvHzCJiHZ+KtVgF4TlkzCmZZ1bnmYmxCpc6zbisT6F
zCDtJBrseqzkSmFzdsZRn1V4zceNij//VZqUKupnXN6ZIHs3+TXEytrlR4UR0si/iP4N3yO+hr8N
dTR99L1r+XPyFOhohf+cZ2k4XA2cOkR/0Q0BazjAL1AhbYCdG1pPB/r2d1+bvNRlUc9VDivsd8Wu
CgzVWQlvlKku+Bg59C6LNMhR/A9PBcHDUUyuWrVC43I8fHNeuaZbdw9AQx25VZUaaH8tBp9szkL7
VISsYNeSCVWUrddba09/JJ1L4uZj5Tie1jCGvjRxAdSLCRXgvgy/3kbL6pEi9nnMzMvofHa2laCl
47ptQme0GhmZ1WKhMtzCgNwmjxgIEdZcEGH/QkYCg6Yn4kt0iIdPvp07Z8h18Z+70iIjMqvr6JCa
bro98H+vyLIC4J6epjo2h5hHaOIK07ZlYzXH2jmyUs1H9qUD4htnlFvzmoI/Vv7c0ZWjNIyVbqA7
PX44riO2i5z84yMSie0VIwhq/SJa2iposz95CAc09D62cm421GqWRtW8Ieu+48EMqUnXCKobFCbx
ChnD/6scL1gvTc6vCJrhmn7ddbSkKnDrNqCtFRQIefKcj7w4WZyNfj8lQelDiFY2s6JiMU439cuu
vL3DxPRauadt3oGrGP/O6TjRCRLdWyvo+FpsDGdzFt9bc4HOcm9nrhG5uVtxdxgqqW3YPLSxSmrS
NepsGbYYNYAvY4FxSlmUcmveaDrZHl1k1LgV2EAGvr0Y2SXsBr9rb5ciuUD5gpxM2at9QBfumEyc
cxIOiOQyiVp3IgoaGXx/WzVDMuikrC4CDfKU6LL1WD9wsAIzmbku54MrUjMWJreOqStCjvMOQtK7
7Jl2ZSry4ZVx0+yWBmh2J/eIZvOLs/5pV2s4nhFfCZCMIQ6tF7KsgbtjOuEsaZNe/doxT5MIuW3E
bq8ZkH2e+u9GD10kP4vc0T4cRfwBMvA2hs3drRWcCGl90i8XNtS+i2ew+bYc5C60L1WkBcrRYEzZ
yn54DvBbnCwkf4n6kNgUjEgul+4Srlx3Ag66QZwItq7ucB8/NmGfA/jsrMmTRFKlhvPZ/t4C5fOe
66rZ7EQR6/mUotmY6KN8SJknrGD6aJEvWnOluNQCjEbZJRmg+AZqSIk/MKm6bGc4ipqO0C7kBxsf
TMhj+I/Jac500Tk2ep48FLvG48eUTt6sRlh0f4cW//BHuj+LPYq3eGDF2LdkbgIT37XgJK6KNxRI
64igYg0ijyZ5XMV5Wfwrcn6NpjfkBmQymGAHLccbi1QdMOHxNxUqQ8cF+kza75eqxlb+hWpBhkX/
Vs8v3bkiWeAsQmzHT+X+KM7PHSWezjtk/KcSg4Y2w8PK9GhTeK7+cciT3wTUIjwtGe+tDfJm7rVL
ljn6vGiHxNEKKGl3CH7zToTwwhg1JWrEIDkJ95IYYd1Ux6mDM98ICxLiRsb/SCjT+UFBjUrs6ylK
05ruSq5WOebkqjzVgUNDgK35i1/R7Cx2MFJ/i3OxPzWct8WjrF8Eu6Ihjebw8/TxXr9H3O8pELKb
kjxh0w7v59YHdZZCXHWpb6bqP+LTL0lEGLQtQCJfNjX/tO62GHyjrUzj14Jh/FNME0QXdRPhd+Nv
5ZjULCDEeW+iH3/kk4tTnRzE64DtIkWhEktCAl0NqYLKFwmnpN6CXXwPgAvalwR5jbpEzbeoXv2x
rROHMuUR4S/3hWt5LOb0rK5DGSatXgogb+T1F/6W1y76j1Hv56oK36AnesgFXb3St3WS/GS4rOFR
yLL20G8nwl63tw14BKpy1AQW2nOVuliwShQnCyMRdAkw1y3h8DBwgq10KGb7//F7bc0E8B8ta6PQ
AIE4LScDQm+F/L/peEjraey8L8ly/LvC820Qw/CCVrJ25g2ZLSH2ihKlVpqP0Zi8LULmfEgVL0q9
4SOGfTszmz57seoJZoBt6FmThGdH4m0LBS6hiX6WUN0XbX3xJMlRUguam45+CUQ64LXFP0TuT6xV
h7h4QLRllI4GCBqvThe5dvn/tK1/nDMIoaf43DMD3UHVmEriiu/e71+rE36mqxIHtJ823Kmj81yi
Firx4OCFe9/FGTZfYMOJJyT7M61ssgW9DAR6M11AsGWCCMeoiJf8LxHYDcOWMMga6s2b1H3EGYlO
AhiFTNcbwo1fKJj4aAbz1m9LKW305Rz/5xxO9Xs924aGcr51IJtNsdiS1iaL7W1qfqMrIFcxXapB
Yl9fBNJ6ypbkEsT1++Ix8EiA2ygt8ffn9a9/TWHPPOqWjyoogIoy08fXqt0r/DgZKg753sH4lKx2
1BojR7FE0UnU9e1HCCDqvfcWCq5Tj49rVeNfdgYVXOAm8R1ilRt/zDnBj3fehmOfCsZ/B68ZE/7F
qheFJ3Pb3Bao3tpPrOtyj0k6CAKGk7fYDIkgY+0CG3YBJHgZdmRo19lV6g/g6VtGYZ2J21X6I8vu
IxCKzDumuKYMKWbILbP8hVRrkW0qhztbhLNIJvnBMLiCqoOPCRUcibGqJquE2Yq903bcOjbdhVAP
ic4ByxR3dWikfDx6/YoddLkYEd63ya3xuiABsXhEkLOzwka21drQe90dGhTTGBHG/PeLcOelAHIf
I8r0jIcIV+SnV8Ja643OMWEzilWEFnA1GkdNjRJazgvsGyJsnA9rE4VfuJlWeqgZ8ogtFrsSu8zC
Jnp9GK/CI2+XvWIVETz2+dHVLy786cnrNv5r9cRfgEgSozHwTAsEacp7nPCH8h/hB+AX/Poo0SYp
0Bg2q9S0tznK9Fe/n6XeYp38qJ7lYw4zvFA/YxwPCu+xVN+MGALVQ2t6601Ql365lm1eJGkEcvWg
VPPVvlzx/8dk5HdBeO7dVshTUFiOO3uxMf90ymUiG4ASKgsPhfAQVi736I10Wldw+/ekWMvHGgq5
dXce6WGf9HtRtXY9LRmIBJKRTRoK43UxFOQrZLdZCwuug/tN71UWan8Vuujm3X/oQIfzyTg85KKE
8+dhcXtoewZ5EdUBTV+rgBn5BnAxJYValfa4vZeUipJPHzJopbYHvBWrKBX+AaDdSt03Pd1UBgXt
BILseaMas0PpwaTCIQit+Uxr5okZOVhP1gJ/QRuvx2r5UluqkDS32n5zMqVbdBEqCh21vGPhgXfo
OkUHfTT+d1M2WWxuadhgeAHkHHM+DuzYWTUhdNAH20dJYkV+/x1BxXbbBS9NWVrebC7fb0V++V96
wmCwSYug19VbdhhfDWBE1r+Ew1srBwzVnd3J5Pp1Gu5+R/VwIMYXf1LeVqdhQ6NHaEIbHNPMt9bk
l8ft+OcayWSngrsYQAA6Kx37UNgVH/XSlKipwG5KITeYTj9hwsX6VQvNpURIfyBYhgBIps4B94Rk
HSDfViudN64uS2ze5pqpTVGukxUoKiKZWkl3D9PGuP7bhiq9mq++VmT2wvwiXhlEy3M5IA687+6/
k+k2uohvjcJyas8Qsr3jT90oA2ww4jC18io0RWAanF4yP0muGMXSc6kYiVSGeKZ3oliMXGzmIC/n
ydxpSCya7NPPSl6J+fxSS+b9FGu/CLhqno3DEf5YJg1fqCQsS4kI8wgB9mZw9JKyE+2wvWCtXhAL
1KHID42SzeiJ5hOt9QTc9Pwxi6ckuqM+XMxdwp8NYIWlisBI7HVxIJyIT6Tb7JoEt0CpmWMQfxb/
eP9EirY9No3TwIGElt7qVM+w3Vk0Yy8dPSU2ytkGhsJUcIBOZqhis1z132vmxH3bTmGLJUcqYqlS
SpvqUIw1/l53ylP+vW8qG1pPK3ozqFzx5DUHZTfJWapto4sEoXpdZ4/VkIMaW4ByOmI3Q0hSdKaU
aBg1HmTna6Ob2sWV+PAsTbVpwc1fWdZuWFEG7kRTOZ5U8omO3ZDcTtIx5SJDQ3y8GhrxBjkK0vrR
ccPW0QV4rczH1z02tmunmYUwRRIQfliEKtkYu/g1y+zD4NFSuDSmkDxKmehEuSOmUW034JVBXJ0G
i7zrrEeG0HIDUxEpTCyrs3NJ3b2WhhdzW+kndvzQK/C49/Wb381nbtcTg/FGiKF3yD2oSYMj+61h
r8kJLsVSbVAfVP0Z1eoqnxhIXTeyeg8+z9vDuyIAx1GJXGSPUL5WuBfIwFxV9hFakngOjDziRBda
8Rq9SAXrh8VypzIGOdwgTNJiuCoIQEyeM9SsemvYWBaP8fr5nZHcS2ILroCggTN5tC6FYrcPJvug
y1u2LSHQTTp8SaGKJhUFol4VpzqEyy93BWGgtej/pq8TU+2eBOZof0vnwn0aXl59++KKFCOk1KOi
ENjsCMHll/f+pd2PGEFEAISu/Sj+ry4AM2XowQ7U7kGsmki0S9GrrDo4Fi0fzz6Zinv0nacI79jD
nHJtcsxJgRUygRElKAqivPXupJ7W54iwrKYcguHMrXn3slBZ5phjlah7pVVlqs7ipFW1aceg4OUI
hxnLRlUuJPvQ//ddIB/4gzIy4BY7W1+g5DMRJnp3kw2KpR7Gr3I9hLmS2lupMfe8zzB0J9vgHc4u
MfNHAEfBzGqWhsWWfPQ+3rBheUBaueukuq/mTb4GmCNRjs96ceJxBeadGkj1RdBHQlyq1cdrZ9gC
tBlP4Ba6OU+A0ps8Xl/7jxHdWeBGntKaJh0SILZUtev1i++2eVaJ8mMQhhnUnW6kdsZ3F3z3RpKU
rxg5WnMdzXFAG1qIQDD+BaAnfru/lD0xvnBHQtK3H3CZkImLfXH+y+cEsN7/Hv5nqTpHnPYUZz0r
KdNb7H80YlaaSbYjS8W+ejbT/rqaHJ209VmhccJtXLWFRlmTiUMWqJ7BzaN/umc+HJjzPG0PPE+i
IlA+d2Qd31VEkSqDdQpr9iAU/vz+x68k0dia/7e50b0Rbx3zHCL0XSkArzlQE+rf1XzWN6apyyZQ
OVMBMCBAHb7gnXIpyW5j8u44/v+RyQDVoVaH/cahVFR1HKWWH48/yTXGWORmn+W5w+6myQZVhRbo
jzJUwqC1CiupBwg1cNw/UB96RdjbHHaljH+p/NmwbQY8ee+XBzZe2mxX4B8UGRDmfxv4EcjDSSPj
YXHlfaWCYmRbOkn2LHnoxjGlNDVMOFCoK3uwHOmFUQhg4uUuCOFwrszB+2+z4ep3kwGcSN0KU5A/
WS3oJZy0OQTO/qSwio7BACIZ9LwFKPpGKmoqBLa7EERwDa7GtFA39dk8IUVXQtjkhUI49FFNTGvr
GWfuWvEayiTYsupOittsft0LNDntAEVt4sev1fHtZC0cNJg5iTtkQYarqZtBAmC/Bx0WPYVWJS7d
1NsFYPcU6STEzY8/J+uBlvEnld06yK1mbg51FbxvrN7L+dAlYiHUzZp4mW3ZBQ7bQMQjH+kqoHHx
QtEEnAtKtImKsXGXA89ZcoYnRZL65MUrrWwiaiHwNyjjn5l2y5jeACLHROuUacWna0dvvDA2zE4H
DQbQ3VonhGra43kT4Rxma11sG9eEcdyPQV/2Dg5KTo0PTvcxjdxSkRngxq6LRea4SPZpFE+7XhuI
GHbYuq1B3mLujl2mjewWVriRpJlatmqE2GLcZcmEZs54Kkf3Lrmpf2S4oJkzDJYvjBDkcTqgsm1w
TRWUsEypZaa6hV2O8sBkLlsriyOl3GU8wTpesXsM6riR5lG8l89ODqb+saI6w8AHVm84a4KcsIkQ
Np6R8oZ/WVPiHzZHG64FtYHqZIVxIYyTx0NKC4x5DP/zj/Wyl0bH1Fya7OUSQ1ZgHg/U/NVAk+KT
WUYpvXA0YqYnvDsD0ZjEUDcqZeDTjmanf3mBRsePOYU4RsbKSkgcMTtQZl8enQ3eLLOcF09ms62J
/ur/3AHVRib/B/KHJsIE53t0UAkR8JsebSSiP8U3+kJ99gF1cePt1a1KX8z38cFv7CdZt1Wb/Q96
BKmDMiv2RMyGTrFJ0tJaP5AeR/LkCLlo3qyL3QZ5p9QCP/bQa/LcZBqWtnlFvGsmwPzxA0I6UbYX
JC9iHWj63WwGRNyl9pG7Nw1ba7P1FQ2yvoXOH+LaGmJJZ5stXFo+0XqJaCfJIgUl70nYoc0OqkTI
7fbJTcQVif4j8ahiv1DK2bUUIL7z0VAhzxSWo3ieeTaFmpCHUTgKB5f6JtE0SqOHjXEY9/RkqoDL
xQCUzA6JK9cKLwShsdXKwU8UVaPenWFCA8ugM3YxKWThjlExClfiokT3hY0mHKC0M74YU9e0UpNB
8t78/O+wW/6SboHJidqnYG1euKPDs4hoYIzpYRJiqDfS4IPiUaoJVrUHLF4FqpuGylmBIS/P8fjH
1Qz+sCz+LY6aukE6HJYQFRgvDcuGk79lpsmJ4VC5WdujbHB/8iwK1z65I5KvXP40NoJIccYpMcWE
id/zUYJmnAcAneIJFtt1v+DubEmdz0ONh1+gLb1iWr9nupbsm7nGRBJo3hn6DbXdXpPZ2SVOVAqL
ksHoBU+MZBkab3X3o2XwrAGlCMVYKhWwLhNY2LDR2+9R8HQdpPyVLXwMquSdU6uOzPhXDQEQ4TPs
lij/2OMrTRDdRKu0r+Bihdl8t3vnkyVhEsT4mNNxZTBiqt/ZGpnKyuIATPTBZd8s/RNpp15xVT6Q
64y4a4fNAgFRaBAm7T++veqnsisBbreWaDKDSj/CflhvOxiEalcUoOQ4Jxb83BxGN8AGhsrqvdwE
hQgYixAqcChmAEIrWHs2/HdkWGil7gauiM402V0tzBWG3qUR9Mw8qtorsF3qLf+ov1ToZnzmdyl4
fJsvK/YwTCWYsKMJr+LXDpSqSqUo75zyS0WJUljoMrJJQFd6DSqZq0zXAhvDSsMoxFU5Bdm67IRb
3sCF4/1a5eCSKsw//I1oV49buq9xwejVUsKNjtJfcovVuL5sIzP5Jv+Z81wsxZ6lUisUKPduZAq8
o9lNIy1FSy8ZLzrUY+dhtvwqsUskusdzxrNj0NyYNTOABoznijb4WyytM/Zn4q1cnjGLS+gX++LS
R0D9g4wm1kPCDVEuGdrsy7h2YWSwLugnlYAuwsr3meHVw6pwdTxZwTOanfmRLGIXx5uD62jeoxHR
nqr+8c+EW1HVzqYfadSEmQl24Clkv/rYWsCwgHGTi/j/ELuh/f6g+vvGPOcvN0mk4nvLVAxM1zq0
0Zy2D7aGmfr/BsiA7ik7HLTs1nwJZg/vmkguRsv2SjcqrKaYg9D+26cLxN8m9l/nP0GvBNg2dUx4
iAnBtGeaGFLw+kxXeYA0r94f3G4y5/kfriTk9bgMdUEfDIYytkdnIfH+hWkISQtHmzdGQpABGnM6
mwmUy7G5F7DyiiMDhGcWIRyDfRRLQFr3iDzC9PEsChm1tAsgFnOdaXLJCMOUWocJf/VWpkPPsQnx
dhWVLbobMBpTQVJj8M8IQydo2hKAVkb94TWX2cA33d8qXkUZZ3GFrLodl+pTZo4y+06oq7SPVPlc
S6HaaP/R7jic+QcjmWdJfXT88AWiHiLQDeVIwtBFHOhpRZke6vRSnJ7Eir5x+JMPGuXxrwZUHPyM
qgj1FcyXDEHMU/NNkcKqhqxV0Ta513GDuDoSVMJYWcvx+vCoEi7rZpcqku05jGYdqUO4CckflnD3
WhBXwcVnO0VcdjTA3p9n0tMh6XmFCzmsPUtYvLA7RiiixX191g+ZJZgtbNB15zgMLcxIz3zdgUIO
C9wwuHVdyMoGux3BE3YXoiZoMvuXRntR0ELGMELtjjI9ebng1JstAyUC/faEhy0MTeWMdIkRsHIA
ln31BcceR2hjGYamRSuqCkhoOVo7JM9h4QW5zYcgoel3UnnS578pqbtY6JTg+rGG8DkPK0PztMXP
4rOYGB7G5L/Q/kHcDoZWGIf3tTeyY2uJgJ0545rqPWqo4uqwNbO5EQIPN2b3V66KmOQF6UtpzwiZ
JrLGqeSvhXXT915Gq1TNAeoE0cFjo/bhFCgAy/UTIz+Bcvj60BjlzNsHSr5ATGFKiI+/S10avy2k
UV5xc7neHoO80FhXmiF/Ry9NL2zwNXubJCDC/1367Vay0EhhQjcDdKh0uMMQnPoomUAJ+fUesFm+
5PzkdSnf15MuUAIPldM36nossjAYyx1ioimVVS7pI4WGx5xzXChCGwvRf4NO9tZMa4M1+0blRY8v
Uo4af19WkVyLDmWLLsxiPMWRn7UBy/Is57vMRAmAPc75Aiz1t4yT3bnozxoBAo8d1TWwp2tX76uJ
BJmu/OK2LxZe796dx6x4hBmZQCshE0Ruljhk4hQihcm5UJAhHVqu3rX4EQseWmrIkAxhyXRF816L
OmlflKeV6JnIHkhELbRznJaPIP5tRZLKWqlskKwVZjsfCRiZnvmvDt/F++Imq+dNzus0rjx1MQag
0gHUBzBg+ac5J8mPhHEJQ1PO6oCKkwGK8+Fv10mI/zfUchLAmX0pZZh+9lHShJr2xTkVeaDEKzrV
Tc0pJ+rSMTZzC2VYnKfR0Xoi2Eop+sSFE20fa2iqltaisZcLuy+bbiHdgjWt/cMFs9P2rf1S5fgq
5G6gZM9GJZEhN0zBGbVfQnsX+ni74tPRAhZnBsRsDyEe0r5ONfV2S35fYLX04YQd4hhhHCXVMSI+
dG/KNh9djJfuPJGpcZt9OrdM2de5ypdiK8ADPvtfptWK52sAMpoT25Ul+pPCHNV0rZOI0Ga2CyHh
nuOrEWGj5IeN2e2TCrqvrD0+kRC64g1xI6Aeoyn21UTyG+P68xBra6bP9EdyCZqv1EuFscPXBIG+
z2nP3g+dSwPIQ6F0MZuf9ywe0z7wlvlTj1rl6PJHXNuDJ6/16wYXU1MKQaWl6fQthVKmOLk0GS+s
fY+VJH5gBm+k56jg+lNmK5bUTuihj0kCWsfDg/z+ufKG3HGSBIUftuVRABBJOHm1kFuXW6ebr7mt
aRbmJ/7t46GAWjrqEMtbYvoXvm/xXh8zZxozmsqxxyjhlDeRm8QAztUq8g/+WFijtFthRpw5Uoz5
nJACcAu2CLO0tkgm1e9ru8+1xjpFY++ztXFF+y6k63ND5GVoxG24cb2RX5PFN9A+VJXYvcs/NehE
9Djpn6ocWCPgP+6ssH3wdB47xUFS8fTKf5FBFzFXlzx8REKWYLcSy2SK32/QRgKy+D2AXTx+BMwP
3rTMD0/1eljNk1JYgp/O5OY8qQKFqw6H52ab/hZW4oIB3DS7w0j8sUlZPG6//z9SN09BnUTlP809
feaRrfovhiAwUYAUSZahmd5DwIpIxXjKwn0WcNEMsQqoIl6Iwb5ycO7Sh8+xyRLFaAy8fsnvmhKl
0jylIIrM+8TAAlcKV6sCROWZe8X5FWGzsPCLrUOBrnI0Nq4DQjZpTQplFtBazUPkAhmouvizrx8V
JWIcaO8x+6a8FddvEY9AKCjrTkZmVu7/p7DOslYzSuOwhd16lMZVcIm0oBW3K3ZY3lSquFtindq6
DadDJfRKI6DccDm2ZD5hM7cpGmNnLjH/MDlqXO9C3Isr3YSpSU76Dgu8Xde4lcymdcaTkuTZFPPW
rVdJLzuy9yU2tr918vxfY6qR5rtL7ZD+gAR2JuwHnv8y2rIPuNESiGNyJ/Z1owUw7/mwx45Zffca
9XxUPsIHNzHNecfnfD7RYuB5Emk1G3DHQJ/aGPuroTZyeoZm/UROBG3TnkQcT4F3H9J7yz1d6E6N
27PIssHOnox0pW8H9/9XUCgoVph++6tMdlmVfwFXlgcyRKWnJSAHpY0siGdyQUT6N62H+bqnyHFX
O8pr74IqUaMMXRDqwte7cuHgNhPV/MPo4ZlsnqXwg7DsYQKVizoamOzo8v6oR80SdpJle/yUIKnc
mtUpKLukCzlt8chMuVALgrTT0hOTEecderTlnS9+L+af3QJ/tVGEEdl0kbxhM9SmepNN3iTLTzFf
yyMpSzZhhi8YUSURJ6cDPGwBedC3kSujt/sEMMQnm5PYl0NhwUonfPjqWmhVH986UCTCD854yA3B
8ww/3WQsulnrcw40k4N+UkWD5nUKrDswrOUvuHyVV6ONNnaOp+N53W7SgYGq0hE5N83PcARuNLOg
bkvxlE9srgNGAmI9VIymULwDnrUJryzvdzUQ8fUR+f+p6P7C1mrRl+ZonVuO+B1e/ln9gWmzKGH7
oJc6nnFXhOU1MfxRsA9fC79bPyHhekWbXBtg6eA6CWSfgeAgta2p6RecgO2Yhmgg6IkJsHGYyHCs
c4u3f86BMeURz6Lwa28SZvHrP3DB5H8K+y3CI43+zQLHs1DsXEi5mOzITWMXXUmf24Sg+IMSguE1
L0HxpYVvwnoH3GrnXnDEANs3cqb2IKFVoaPUj2jzGIINBjRYaOZ8B0xoDvECszqHU+yX8O98oVzm
75I0FeH7WwirdwSlPsU84y18hTzaMbrayaE5YKPIeIhVDUQ9cL35punqyEyyKAAV5BL735lD34jA
0KgexrTbU6USZrI0R7+PF/nMnOP11t5QgVu4cWRlkFqL2OOdNEvZ54RsHkgGEVowzDxuCJYW0L0E
5Vye5+cfHcLTPNUsaiFw9V1WqWuL2/rUY7Y3fYZPzT99WDFnnzjCxJ1skgaC8Bli3hBG9RW8UK6c
ESSNjMxceG9KjHdeRAhjjEGi0P+FmP4H6pXHPWnWMAkc0wN5gWRENJxBya6aJE2BOeQZve8plN5Q
Iy0+tGHauWQb0N/1NBQpL1+npHy0C9E4AsOcmtugQ+Fj2flBe0Z9k2u4FBE+qPFayrhsgvnjLpym
2U1Jd7U+2kzNCYx4yIg403aIYD2h3n0TjrFCDsM0qM4sVZDuVdTIwZJzX+s7LDFrfSHiMS4LjyFj
AeM8wakTpd/h/HW6N64RmBmQwxKgMadcEZUnhiKq/G6Xi5dAh7H6j6/aV+LEh0anhE2wmxRouw0D
R1reZUgtIdWKkcHWqR2fZnAHdfZwy/lKn3aYF+/Rc+NLNoj6mpOGHlS47ceRm8bfQHL3GsF8i6n2
QA+4l9yuKKcj2uc6xWJfzKyu63cYhefKZ7xeBvFxtdGIzK6zixjwh7TLa/it0b/EVeAiXfFEI594
qlaj5vHVYDz28BvtnqmcCiYYIOEZK7hD1Qpg5kIEcAPt/Cl2IyaxGwLdKlfopMFY2PwvadliX+8d
4PVNpNL2r06eQnUhRSBFXzp+Hl9NhEOB6eH+ZyFYZ6/P9p55Avblx5XmjDpSUbpycSkIpvOaBpFt
uz0mnHEpKkWUe2B5JMzJpEwEbDG6cXjMML45LqONqTzd13UciBILucvn7KPqryhSnubn/LJ2yOAZ
W+oJ0tTjRNNjNtJLma0SAJzE9fIcPablTIdzrZE0dAzAzvfniKDzKg/S7n1wf74kQmPoQur/tpLd
k8OeuFinDkgdt/c1cmvigVxJwAqQ3cGDWV4KOow/dkvlf9nTyjkjAwtusRdM1XQPUO0vKaTGg+JF
oDjwB6ssJN+4RMBKumQXUAJ9kFBi9qAaEmpxCxAcSAX0HdTJri1JFmyzglJQCBSyc9MDPWZmHLDV
n7Fe8ARhWi7c0HkAmVV1p66vmp/pxb1brWnHz2DrRA2vnIUt5Kd6BVn4sJpGG5f0q9eYOTupv5iT
TqBzcrBrcmkkPspY6BzT1hP5l5gPO2O9Bm7iH68Qt987rN+4L9IlUpKcGigOcMuqi32B+vRCSOOS
Ar2DD7EGbQ2SNbnk7f13aMF0sT3OIAwQI5AtwSWpVhIKPhjsjCxOW0/QS/6/xssJ+yFN3wxbArvX
Pb1Hjufp/0HKctAKQ39UxXWPhhg9s/iyJ6oskdwt3GcWhDO7eTqmbc0VZA5tmsVdI51d0o6pcdRh
Y/FaevriokSWLPGOTG9g65ZePxDRBY7vwyxblZtbapvtkCB1TAUpOPI14b+8i88u6EOvlr8Vda6V
gO41S68PoHFNjAwpMad3Ms6/INHeuSKWx+dnTiCXQFyPYlZg5hrsFBJsIaEI+OQJhyTEdZy2XmOe
O5QMAfEREVtAWsLEmRlLEiBwaHbsyXeaPysRYARPbQXYW15Ju3MbQNEIyVmQUkZe5x8N0ZULCd7o
NdheKZTtkVbShAQ+382aRUoVeW3ufe9co94uku4pBZFxnOiTbWOLZWNN/Zw1+/oH+CZHyFI/+DME
ud2bK6T5BtzFprGPPUwBbHzNm48eEWxdRWvZqBk7hNJD1ntjTLHNskJEXS+idpTl9mWCDgB483xP
33LdbeZsK4XArDu7xXViJc0+sW94xloZCBod7Oh1YyGn4K9C6hxXlp3YdsHuYFWCqS+3zq1TncK3
EQZDlBP7fcMFWXttpFao1uoTn21660bEyObAET5pmjRIN9ETVSHoXFU2OHBc4hlguEXLYeFQbYeF
5me0OsfvteCkFuY/doVTJvL0wv84cc7pxqQlnpDsbag1nyQQHsKYdW5UYBuYFY5x6A2TyuYX+4VS
Gx2H7hrUjzpGFTHwsN7hQNtcxVE7FEjGT90NRNDa3R8Ee+6swMxQA4bG6fNWgPGFF/vrBaBFSk8a
jyw5+gHkwFewVIh2rlu78UkK8ENFM6+vy6Z04dmw+jFohS8xb1SirUqFCWAUnupWg34ZKnTp1GIX
lpDFScSHRIO+iKi622KajmppXuxKIBKnIkaa9eJAXPOxGnzxCxDbYCLU1yM7d7CW+cA6p0R6Gvcv
zAhd6N0CxwIGo7PaahzSJFZsdI1ON79lryvuq0rBo3XjDPSQQrHSo8+kHMopEVvMgO0ZwEMNX8Ft
v5Yf5ckEezdU5V1XajERnB2CmVEhFAvfZXjkHXPMNxUgwArLZO5NIZT0Pzi0tRTaBa0Xbw6dERQu
sWJjjfsr1TJu8KaurylgRwqxm+pj0tawKljUcWIrPuYIk5ddXrI/7Q9OvvYmgwrcfbw1eBCBADFn
J1/uI8E65UB7Z1poejeLWGR8UbwnI7FzL1Xy99vKeIgyB0bcEtfJwPAwl0BVVOqIDEOufCVSBCe4
niIvWBzZF9JYbNuPOZt6fjDYrHjl158nKsfzA6cIyZsqvkTjWzeU3l9QHoR6OpekSFIGlbupZ3qt
w0pb5nr/71pLhPJAxqrzmxjlJD/0gIh7pGMNayA5R06cM6aBVmPk4Tif8CEEljEV+dwPDMB3+gan
bzcsQ3H6MhnoWWAy7Vp22rZFw15ZdETArz+RCdByf5yIdvpT5/86j0mdP1AWgGDRTLO20Hobmgd1
pc8RwIPpQww04p37mkc7zBN1ZWpJApiPvNG9dsMEIalHF4RPeQ4iQqvwx4dceojmwS4MSxtNNNXq
2rAphAyg6+0XL79SqpfSqLI1q2BuCkU42Mwj3FGEgdAsO3Md50/HuxEIKi6zWHmgdl5CH4XfewKI
SSZfattgTLnFQ4NULRDiGUizkCMBltBU6DjHVBBryigLnFYVFa3kC3/+e743cpA3koNwslUN8FDd
vTzMcwgy1FRKK88acncieXUwQTuXG7H3gjnIV+iGBHdReEW6AG2ZHttjU8HPrq6BftKjA+CGwoLE
DHSZA9O1usqZy+R4FgafHWbcbPSrOpTTMnLh1rRWn/xyItUMRLVWVtiOHhUdYKY44F2Y+s7RBBn7
hHU+ml+PuYH+DXmjI5Cpoc+iXzmM1fUALwq5RhM7CoWPPneHEaP58neQCkkovxCaBqRv/I5r+bi1
rRuLCsuJQf+3BRl9iTugyEAdCu8HibyrJOH14RUDlYzI6wl9ps8zQcwd+wBGy22zEWOT5t4JS1ir
RfykWxRf81pcZWHddzSLxx+ySpOOR5CPURsm63zm7A1cStkFrcJpbhfHWR2U7mEz8NCh/zc2zSS9
xC4f5vq4HFXIwidXuKUr4vbi8tWKmTX9geztOr7zY/Xlr8FD/WxjGUHz3OEarvr1uKcxJtECxtBA
F7GxqfFN5hHBVdmRXKvL6HRlpAD4+vDPSMn7Mc8H/W9xyRtYAsf95VxEG6whz6QoetAUTYSHmm80
iFXdB/AMPP3zTYuWi9dVZmJ0Kq+Z4aZXXixINWhAZUhK9zcEOoeFqcXCzoY1KhpyIDOL55cyKkA3
eo8+giNIZ90jOrn7HKi3GqEdV9XtuFxI/dc7c9ytsF3jo20OYA2Eu47AFXoLB+EwuLsmTvl6zlG2
Ns4US+jOQ1Mi3yIM4SqQ7hOuc3CdXNiwIoywrxbCzBYq9POMsApajcBfDW/jc6voEqvPkD6xpqIn
IEFUs/ZCzjDZjHj6exTk+LisoD4TuKCkk/Gsw6WokNtqggw0gXgwMPsXSXuYbGfMhiiCX4C/00RZ
xlZj1CFqw1FFkizmhG5DUxKQc90e/txAgyyyRWYgl6Kq6LNjUajDjujuYI6ggluV+Hpiolybm0ha
TIaivXlIa8AWwtRo+Zv0Vlt2TvRqC9AjQX3V86VlsKgqkJUKNlY5Gbn4VuGCFnQTK2bAdTG8WJrQ
9M1TesT8N7mi4YwlkgyuT5tP3KjYi/X5nXYxtrDxxi4C5amJtqIEZWojNvWzYsze7kb3VsRHRTCM
QrVaEs+NhzDf68GUv0uy9b8UfZuSbp+7x27qDeSp8sQc1MdqOVhNLGnvyV3NHncc7q4RVOzqqxbU
07+M82pYGTW7yZyqEiGULMz+Ng8syNn2adLutOnnEQHKOir0yJldvNyHf/V6lFHEwkO7eSn07oqb
AgXC1+a0LZ+AbV+fy06xGqQqyeVm89rkgnuCEEzv5E8VJuDEccDg21pyoOXVP/I1F32NNw9eBrVW
ZJbTW6iumeR1by5y41HLsSXRtM0TBKngMPCziOmX+SpVLWVYzRncOq13C/mnojwD8M2we0lPp6u/
JuoC11UlB6xXtZX2vXlkM/rxouTTR0mtQ1hfu3pxDbLRiQfg4EvVEZwzZblIeGWjg9FGYclQGCr/
7vyoOlXfM9vFdng/JVEb7qq+g0/jbDYdYi7Bx7vCIutHeNTBiDQzBxjZJsDOj4Lka0SBGwFBEZo6
dnI9v560t9jxBofciaiPp+HT5cdJBtWDHrejfuz6e3rJFIs/P1vDY2pb+L0uB7zDwRnA6t9zE0K0
I5RTftPGmOlqK1vfAku9HFtf4NAeu8UQEWLoFOXKx60ntdZohWSFCOa0YUK6TLU9VGc7ZlK1TU7p
hs9A/dW8vtk/j5fe/C84ru6OzbhAsGWT71KqrNl2SilZuQgdK9k+Gi90TX5/W9OCZog+1lWenQ7T
Wg0mk4Pn9/5mnqeliBhSmO16lqATTskITIDHvpBwCRqbcF0cADegzsHArIxsH1lA7yiK1V7z4nNE
KmyWZNlqq55+rn3TY6WsmNvc6SJhUkLt1GZC3bXKMd6DviFq1FPJmmhwC6yiCbgmgBrUUosJ4Tr6
+9TTGDA5fUcNEg4GAXnqw/r01RpiDBAtayrarZwX9kxc73Jjw3yjXmP5zmKn7frfOaWA8x99Ntjh
BQSSo+tY3iCZVQRYqzBNAixdmDoilda8UvG/5usK5Ul4geSPFyRyP72ZMQo2B9s2BEMd+n9BYOX+
Pgu9YHL9d9J5kkdaY/DVSt07XfnNGXD2pmwQOSvlq9fyOdadBZ+AceeAmpQMJHC75zcRg8vhxK2G
54PNU3+C+HKh7V4JuguSFjoTEljSKP0YgrOUc59aKd2W7HhXNhTFy/9xF5bwysAC2qNeAm10jgNQ
cNiMoBwXr7cN/5Izkw+mK0mnRQ+G3EuxrjUnR7U7e7CUK2Lkxvp3WLytCSdAJ/G8vSf3ORfvN5RA
ahXaPCxWt18DfICoyGs13NmEnJn1smjzGq7voKMRJ75cGT9MnuBKAnrkO/1tMBdchEA6+czvn59N
hZ8UseEMGNI3JTU/gUaS+P0jcHR6JywUsNOPY1OPZDFeAtoFYALkJ9x8rR1+8s3ACBtVCMJPASSh
LhbUUAQJc5O/sOiuM6KsoltARp1fAnlLYdMN2KFK86wgdKynLGMGgkxlfSid5pR0I4rnXBaxBdse
Uhn2qSPeBczKjmp/kc+6JuzY5meDUbsKWOsCyv0vJSbAroXtLzuMSMBW9hPJS9nIwUlWWW/+trp5
dsYHNFK9nLhimcFSl6CIO/SQYnfzJNGY6MDrpWehQI2wOJmaSRoCw+iAv66qKYKFywm4/VlqLu34
i0WpRf++C1cXga04XAKHwVKJGuzyb+mZZgFTgJAXrUogWB6lc1HGYZpTF4AzDhFF7n0kfb8bl003
S/WgeVNUbpjTWqWRI2+FzH56EShBfs+6mLsYIFDMGCbV9s4PnnvbaQ6sfqQZyQypwVv2hkAWPaHo
nR659esv5u2piR55vkNR+6H1sZvFCzM9E0eKoCVFx9Kbpnx4080i2H0kqDWjmoHgqb+LtqY/r7TG
82wcfd6MnrfTSZwwsOe6DHwtMDZvujyLICT+SUY2MmCQoI1iMQ55/vNXQT50SbeGUQzbxpyTU6By
krPsUFBg2400qai7kUPdSoq1EiF9CnPsAVPUOD3ZPyO/7FvzUPLm6xDGjd4opjK95Q3Gqtv+xGge
hLHko2UUPmBMqPlyQ1Fs50PLBhDzeqmaMvbuP+WrfTSsFtpGFThkdb/Gcm0Em3CBjO5T70//4wZM
WO0IZCFHAH0Ljx3lPW9NDbFQwrZ3Ynkh+JgVYC6nKsuHXTOezgbq6HZCxVKSSvj2TuxaqqMwCjT9
CACrmTh8cXgKC7tI5YXYfKug5OUqNclUZidOmlETAbFkoRj1MzXKLUWvOF4lrC9pSZZVeACRatZV
t7TCCr35ZkombPkt07hbJXYYIrwHpmSvUA/sD66CJptkZFQnKywU1Ei1bhBKcJVDZNtMVxZA9iAq
xOY21ipGoX9phGmCnRehzfbxS19TY0gVQ4e6D1WBfkA1oEyKd1ZMAJqRyRxGu7x5iOgrjZVctCiP
M6+ovwr30XnJ7o+xmxfqe1Ww48pyn4syqLEMYp6ZATGS7LNf0I+NvtrJ3WTKM9IX6Mv9SDIcXRij
J0Uh9AIv3eBaLxgL4v+kF/3ShH7UbrN34dTHIe/Pw82Zyu8HPuZ+P5qb1WAAPUP1/W8BQmE+JnE6
61/WxwpxC5iqJlX2hVC51nX/eZTlaZ6xd67kEhAzi+IUdbsywVVRSYpevyUGeQf8hGgO6GIEaO01
7PuOynegkSyN9o6HKOziSifupWmPLvPMrLw6dBb02vGKoXzlUAIwu90/bW5RTNNsWCk8FE4SjKrp
TTJ5fYyztKAc/s2pPglsA9UEVXMmYHA5s4tvNm5yJ4gkRnSnPkN7w8JJyVpHJfFc5lJns4wmJrtG
ymM1dLfa6EzNmGrx130pomuSvLQRkIFJYYNq3hbeyqrhra374jwFHa8Kz+Hj98MCzpXB5VubP2sp
oAJyPdjdgzwn3FACDemkPl2vgauok3NVpw5OIVhNBO7JQyRJ6pOTjIYDSFXlLzTNibIPy8yxmFca
dxq3yh2r/76tNNpe55vnTv4+dyzCmP5mBvsMkej58ZQC7VJUSNrXsFNi+9YwwLEHKEBhcqKedBhW
fL5tfRcmKM/mHupnHUCoQqzs0sgrqqsua02ZXYj5UzJcXMpzUK/PzFiHkHzmKR1EGJRtdk63XybV
/4ZK6LyEQQsoyGcYzlb62ZCziITer6xmjYF0dsF2sDq9ivu8bdYbqcSBfEUl5fDbi4LLHJmIs7xS
EnXoN4eR5tD6Wkykzd87IgmujD/JborMHb5L0pE60PL41azPmv+rQ+FO0qvmU75EwIlYZhMBaLgA
1JFXUY63FCRrSratD9tgn36h2ej3R/N1CGTxSa1D5s4Oh4gXN6P/OJUYYwbWegxYfAcBaLqnrLup
puSwDPicuyOYDjjEoKNpUn7dRHuwkS+8oELQdqjV70iW2OELYarDC4sEpKCor2MAXTe/pepPiVpm
+3cvloOmIdyDo5SNi4xidjV+VeQ/7H7tgIZSq0Pf6z6MIsvpg6kcON0oK+O8Uq+vES1Y+0SqQd6u
VnRrgN4E7WWNeVIL+Cv5NPYzBWZiYYPj7R8zeD5FLoiT6H1d54KaTCh1IPwb9ObahFwZEHHb48xt
tdjnKGYW8lDAU6Xv5KUPaCbUOEw+Mfco+5bPGvylNvLngQdgengWGEGoC96CSyCP81HXohQtgjwc
AJoPLH07SzUZHIyCrNlynypgM9/Mccf84a09dkKK0Ht6wUr7pc+kpyyhjYQcb9bpx3S+J4W8moO4
RcSWRw0eocHX5PKrAV6J1fl5N3Mnd1+4M+sWNiVLpefZNJbKdw9ZGMPfdKs/lORiX7dvhdVQsUYB
zLPO8PTtZ47+6t9Y0rLrQVCeUg8P61i3SNhBoSVsiv0+g0+yiFqNnE7cXWrZabj9MHt2bjOZyGrq
xAqiIsknM5wOvweILgv7hGjuMc6qVcJ3Aw0DTkL531PRq4q6SSo5wroaQgUcqqfGmLiILyKcl10b
IgzQatOcAnr30k+uInLEitSZo35xAWwPpIxAIKdu7XaKbUXzNR8bobQnxFvWl20B1A4KOUa3yENG
3ee/sCXuGlw74Yv1ii+kRnAnRAptC6eOsEOTNHQRc7heVa6J+b6m3SDPjdYjdbUTSXjH+IQQ4rrQ
bjA9X4dMlv/B+dbmmgZ2VG7dzvyogUIkcM2pj7eu1AgTarc2rUKIf59aDXR681JExK6gBmOiyHNE
rnV6rjSoAcfa/OEU6LuJjwFwRRBHkDtJ0BkHZ0K6rR9IM4pUY5ugWohZdv9lhW8cxhXcqDTPo2iT
zX6M5z2r70brJ0Mef3ATu87ZPqvvAKJzOX2qBIvI4OPve1LAiREKtQle4siUJdxR1dfz06cEMNlj
iDIzgEFYb0RwdpqhWB258ucR6/1vGITk8UUzA+krxzxuBn7nyOlOU29jrHfmUJ+BbmkeOiq1/6+Q
akJ75ybwRDDfQhd9q1zqh9cHGK6rIcP+lmYL1CgkIggul7D8mxzlbOXOTpv9xJNy9GI8sCI3ItR0
i18AHOoBHRk7Hl14bydidxFFW9K1nohpm1GcyvaARm3GlW1CYQdBwB8UfRuVpnMxnwniGu2nG01b
hf70yU6hBh4tlbRvamKkE1FoMRxmRv/2hq5yHdiL2EKRzX+YIsGvl8+TnmerFiELJiSeLFOY8m8j
W7PBx1TLeO/8i/F0dbBRSFlPw7ZpHEgx2kBJ+79kUrrc192QuJV4Bg0aU6Wr9P1mc0JTNCw5EUmC
ybSzYW1TVbleZY+r06eAORO0vckbjPaQCs9R3ecUCAC+iZZFW3cRlmUh/NNgqiAJYc8GW1IYDwbp
L6r+TzAgFLURYfrbs4pHEGuo0pdjOX2mdzkHI7WVCB8DFVRpx+iyYs102fW6hF/fhK4ERVcSwbWy
OjmmxU8nsqntY8N9sUEUxVTg4KRmU6IQqaDAKC/0biiXwrQzeMcOe1B5HFqg+lINMcQH6OksiuI2
V0gxv47YM9qaPhI0JFMe2IpqvhbzZpD7cdEfU7ngNGDK9z53R5i1NQXIKPmshbYL7zh1ZgEoBrE0
k4gDImSJogcdhC2hmM+bFlG3D2WVgFn4yJ9cjMyQ+5IUYBVz3sTXD6j1uVCfeHm2vG78Qu9IpYcZ
xHp5+KJCUljjo5Xt5TITjNqWQyd1JCcS/mNKLp0SPBdch1NRlCWj+qWEr3cVNt7MfufHyI2RQBwf
pT2ZQYWDvdmP+R8BK19PateKUR5wb4S7RyMZAB//c37lrg0L7ocLTmMBQLYsxJqyeBcIwUGfG0Wp
gokk4yF8cHP2Bq/otiiJlVDcc9UW4IhGxJN6ajqbiRzPsqKZalWVYWvjtQoi0IIW6f2pw7tD1hL6
CLSrD/SlB94G4eToj6Lg64DwzEU3yCKt4tuIIktDhdRs3Kx7pWG1ZuK0or3o+xq44awgDkyC8QiU
cONYu2ys2dmBWoOukUWzHinpGnrbB1ZK6HOaZj8votReQnR8WAdlHPPARcXm1HDqYIav+y8HuVnr
UWItjffh/SDzvSOjaeP9ZnT+GrWOfV/OhDJ8/jEdvIoMYNDvUUr2KBqgyWk5OGCvJPh5JM9vfiYu
m6g4wG+DsN+54op6+NSTqoC3cMBR/FphM58hrUoM8ajHJjSpUIsTe97I/XnNFaobEOmE96wON41Q
ToZ9uJ73uHHpdfMSdKUQJKwgQRGr4ZBLEzXQe9kIAJrjUeJwDTCJJQe0qnE4GM4+hCEg5xGqRgFa
2d9xLKfqN5awph8SiBEvavEU9y6TDNORqHFgeIzErww+Fk2Ek7KqHfpxTLaI67gcj+Si5tU8fETn
1FEvz40kGDQSk4I261cF+2kY9HlfuD+NuaXr3qXor1XEQCcGn2xRZIcXsW/5A0J3Awiusc2353Nm
D6csVBeIwrZrfvkzzNRiwCZsxZJN6fsjTqZ29G7ED7J8cd9mEkw0c1/yGiqOMwwHobQeKN0Lcisz
hLLGcIuS9X+1H5uSmlJBqMex2fVnlSw0dLMiZYBZD3mCmO8MAG6vRGv0LBbgGtZSoOfCttiXc2uI
NQSdtzZjX0oOlIr222cK8b76X3eJqivweLL0K8Qbbmf1Yk/Z7RmPt/mbZaL/666o50NvsHlGuOl6
EA1N+TbMxbmBu7WFZ2D9LD+fYgh4Umfw7RdLxZ/KNpw/wcBLlnL0SxrmyapV7JuS1DNI2ZxLd2E+
S1h68+on9204yjho1oJOhoFklBF6ix/12dn3VwkEp1aRIEBug72kVUCdeczRMXCDDaNcL/9aBbVv
mE33hLVf10C1cY98bZBtRAgUUlDSST9RHTOJl13kueWB+E+vT+nnr8HCca8Ap0He4v3Pwa4NECRG
gz4zDwuDi3MYaX9PTYjETwoR94xRI7wSWmsFqc8NH7bIgNbZvP2mK0RoMATMqzcwP4xDIszQwKLu
aYrX3JcMzNruT22n31WMpoxyb9m2Qt6Ra+4T2DHY4uXLw7gqNOpiskwvdLFAfARKervQs/9+7UOk
TcKDVcnjvSgzStHLxUXc0O6qF6vbli6D0ifZWxHEoHH4NbgNCaWPlcIcDOIidYQGFTO8ad2kyzWC
9BFgw5nHrnHC6/9WzylC4bGILW9yyREvzrrpnHYwTbjNHE4DMQ6QADna3GNG060m3TpvSQLySUAW
VkRykz7YITNrQUnaGMM529VWb9WIqZlAT1Qa3MCT5PA2+VuiwXiagHaM1XzkzXVq4Hz04JueXtnp
RqSmvwloFOCgZy3ysZzW18XATSOUM6VRQkUs9kW7F4db1g32iqk+oH/HuUbBuy4HVO+MdwIyFXPi
ELGzizdZ6pkMQ0uqNO74UZlT/dMawjTj2rHGoJ1aNke4HATXze6NOpPgK88L4PuyfuUcjSJbaBMi
ofzblwgInOu4OUmaj9sbXwv7CWgfUVpidbwLJB2ioV34oRsnno1jJ6EYv2/s3SdkNF35I+ioH/eC
xeUlhFJ2Phc8ki8hGUeHJHwcbzWvte5EZ53dsS+FGeNa1adxrcqdU9WPEQAI41Z80wXFzebOgBqa
PlwovIxFrSZ+3Bocj8lfypl8MvjOmRNArcP+SrOC6xC7y4ymDQKF/Vl9R7B1QH9T4ZqD0gZXwMsH
jRCqFOGj/SvaPrqtc6uPjbO+4PRUTJ1E8KcBMhmBhOp9PQxyUq37EkHWPXZVry9B4/KhSqzCZHQu
W4H6Vqtubf28tdWwvyj27p3fTtU2/Y8aoSFaWSf8UALzVc4ZMlJOQjzgA8KWW/l80wdi77mln6OA
Qd7eO7NbpI6C+zGdqaZHxCt87mnQSVairjy+RM8ABs67WHB9LEUMJv7NXZ/2fG4G54VjQQ0PuQLa
+m5vD87ab6pgk2Igq8+LVhEjeJCBaqWlLBEeKVjD8PIm4F7wQnvpaZZcWvDE0jDf3MUQOBTJc+au
qK+POjIqvZd1XTReUmEg4JoBO9t3OXWieDLH3tIwKVmDkYHijLSnPV4Zg1Sl174oGyZ8EoqAj4CE
ks/Doa5qBT5pIt1HrxfX2ateI+s8YWUi988TcogJS/1WDpvhV84mVOAKCpTBViOSgj8GVycy8pJE
q5k5vm42XKULwebMs8reAXK2PeScTc82u3a4CVfr4zZdn7mM2PCRPb1MhB3g2a99txXoTM8fbXBu
rqIjrQW6378o/OgDdv2+7ra5wHW39UltX8RuBwTl4EkGovFLMRqCrPld/88AG/N3IWUafU4Rv0jD
ZdRk016mXAGTftrz3nS4RD3Kb3NIWAuCC8cMRQeJThdRb3aqrtvJYgxGxjq3wpQQnmzXBP0qbdjK
0ckXEhdB6oLLX1rYfn+iuTdaXSx80Nb6W6p+GX3zWHwvqihysmmehmCcqk8FuJvGr9elPG1gqsP6
OUKg+F4qsf632sDXt2adm5m+TD5R1+qWv0HUhrWqB/FoIrfy7TdOVLjTLMJ+v8YUR4WdoCw4tons
N8wv1NLs6SbjIWv+ZqMKAjAYjjPuz1NbAWudzxROxBmCu59G6LgZdFZD4tPcGTXJz2C1mawbX2z+
puGrrfkjk8IER1ml5V/6Si6lbJJftrFn2NmGbA1dDoSOOnkL+ZN27XXcPWpZJqmTgIZZ/QX5xhd3
Oe9Y5hrBRwj21tBBHohs0vU/SHjoqvHpO8I+Li5/A1eIXWNkotAjXepsgFZcKeO6160MZMaB3GmB
leIiQMxTuh4VKuOUMlcDZStCcZ2WEFjakGMRZ0WGSr+WiXPtt0bQbPn/fiYqZ+0oaJaq8GGhvn6k
8IknwsRmrHQnaWkNm6tz5UC8pOqbanPAEMEHy5pJJ62DL0H3QdjyyomVzLFU7WmGyE7fEAng6Uss
VmNIOw06/hFyWc4ZHJJFX8ssdwAxFj6xZOZ3JQckeSdzOAA1CuhICXbYQ5TwITOeU+PlntfuAXPN
+3ZTmfvXwxOv6u01rSwJmdvYmzVOhlGIwjIsdy3uLRJGT/8ZpbNtkRG4inwIlyDleGYTY7BefByr
Ir7EqgW+XBUlWbl7sZyC3PA29YQt19jlrLwIpaCqcol5oTwtWPmKIDj5E9myMiaEucIIQ7V0M8Uf
r5V0LsKhmOoRnkON5f/7XESaWAiDewN9ucOfxEtiEBWBeaEPx+pzk+l5To3CI5l75J7L4skWU7vW
UCjGIS8lK5PHC2/q7y6gSrlbl6eV5slU0L5ajE4CTbOrcy2dXA/lbA4zUNUEvTfje6HE+R2POJ4z
8b3WHzTCOpDMqGkwAs0Wu7+3F4W7zLsykz7L/GyK1OJfkBcMbedglGhB7w4rpx2L/JqocTVtllNA
DHXPb5Tzka0bhaWq7dHhTK0Rf8zsRf3KGWcXSvlwPqnzeOQW2CGsTDeNUqoWdDbPMJoNkBJFZYo1
qPAnxEPLBiOa6KQwtpRjndxP7n185WF6hw4oBY7mMwBqMfFsvaegN69EcoNXzvJLBIvvjFDKoaeD
SGyyW8JnGVfmJTQhiP0SmhzOSCgJbFX+Y3nlGwUG26S+ak4AVaB5CGvGRtvwoKUTHDEHmf+tRGNi
s78XzeJ7HTK34SkDWA6PVGdFSXSTsonrn3xdWhnBp307Qqhi5aY1so6lXFGhYe3l4MRK0M8+oEEv
0I9hwuZhmYb3jSuG1IWYbUshMvjqsGOuJDHKXAppsdyklDOnm70ZF3pG5I50w3FqeBvUqQJ01xlT
MnbO5uGZWf3D/irE177fagWtrBwRmGFECjsDSE0+SyWIEdRQPGOMb8AHB1rk6xY+3Y3HbOlvYp++
kePuf2W5dunWweXb6qw3gmtSzT+aDFK8gs8cU+pmKZPZjSrVjOMAzp9bjgkLECs82Av5/ZI12kt6
Fil93BG71dAjEGu8nousceou5y11DEkf+cCkCzEctGT8RolwuKFI16uH9aJCympcOZtWN2g3Pi4M
zgI2wHkkM1EkML34LxLbMNq5g5GYlvqQhqhVI/DkvVmM6pbnGvI62PVyOMYpxWzUnB163k/T7JHZ
A/6zbptcevFFjUEWbGWoIGgXaiIiXCK63ZxXi7DBlPfsZfZe5zTZzmqwQJojcTivEYPqkU6m/v8b
ZCZu4TFzKySBbQIMiEqfN5Yfx8RMVYzZ8nM/Gq2O/bezIYRceNAD6XKT9Ega9hV1TlxUcyqvx0sX
G6KyVVbL1c4MQycSCCaPjUKVF1in1bEmN/AeZlxA3zRbOEGT2L6U3bFJJcqbP9OcCzXYd5lEhk13
Wr6rvMVzZYBmhMcy3zALrTvNDODTDt5IfFz4L/A6ia2tB7pms+4WI27i0GfasJT+9sWfX1FZAYVI
dcmJPfTnMLwMUcmUhO+ttt4Gk66eghzbAUGPom11BknSTM+Vax01DEicuV+Sexxf/q3IjPaCmvna
VWqQGZ7s78kHxyeYH+j6su3/GP3khQpgB/WuAxZcgvugfbyZriQD+aNx4shapkZc/Hzb7pkfIWfW
6RDpr+sh7iCXJrTSVZhUSExq/Low2sDDXpeJ5PylJhAZpkp/sB5yfDJIroO1LPCGrp39ixSEHvGA
J4duBkFYp23mKYnFBt/YGH4THz8LU98LVqKdw7Y+JFnQH2LR11ubQUCCbpracLyWbMkQnSSsHVOq
kZ6++hzP2DKlz4PESUMMmfXInF+Bn+UPSo2RcQsIkmybQJ5cTYu8KIaCqOXuXr76dXFwG4mGm1d1
JrzJluqUMhcI+vBHvxOtqFT7E7HPJ7oBE2GJdWE9azPbKKAxaxU77fJ1bia9z2lYXjW4yFdqeOfq
P5To12f2KacwupIdla58jtYa0e264yYH31x8TdrnTf80FJ9+89DbVUxZN08gM/4evh/yFnwoxLDi
XBKVVXfYDY0OuxFa/rley1OWJfP6xyQUIRQMAT/60NDd9oV51OLMsLlFVWLnXQ5l6e8WXt/d8glJ
NvpSqwNLs5J8sWsv4ndnhA0XcAp9+ZnsYv1smbGWrBSv5CCyoPDPZQFUOEa/MGP4SyTFnhOT4Mu1
9XyInr856l+7WjJC/nK16caNdx8D0Nvh8oIFi+W36+eeyKpqi+twdShSyoMBEXEETPq1Gjk35N9V
g2x4AaepKkTZkiLzrqvYIdsEWwogCdBQDjtA9dSnXJVqpaW1YaOWitWY3eLJhKfXSKyUixMcomAu
Swxy2dpBPX2GlmbDsCpzYZqWyVq0IpPsmmsa9C5BeE0XrDUd0iI1OF/skHjO1Xym3nRWFDAaOHrd
6tU6z2jjRVYlwdVi0H8MVUj8fDoKnzB81670bRrKZFKfdkaxRd3GA3pApV0e8EmeOQcLLBEwwtcE
9Q53t2Tgkk+maDOwp/2GXw05dfdYkZ2WE9pb697kJrjnfu8VnfCslvluCBCg6gTUDnWI5du7MOQi
f+ot67TYRUu9zGlKLvE7ViXQHcA/p3xYA/sj/HJd2Bxp2urCH7DiMFFK0yM58ylwmSnF7Ax3fj1+
JV1jLd+qNpIUQVFW3ZUeULgD5Wvyw55fMJ0XoPtnGygaU6tzK9gXtO120jiHUisZNii6AnP9OnOx
VphZlR7SFs/Uom3Mc5n+R6zcftMQpPAoacPQmysHkOBdYvDPDHftmUfrg6SwquCfbogAobWaJ7q7
3bFNoqcQMb0nOmt/NQgfYghB1ntzEEDFrjB9NCmIzfU+w7/wDDHrs5HjarZYBfmGCQbtAld+ZEdP
JMVpSPb+siiXMvqcAndhqWuTO4S+y08zMIdkxr8rsBrHv3H9v6PSLntqKNO8r6piv6PDTatwFCHX
S7RgleMC1kHtnDPYsFVDedW9+ucOXD/m+2mC3VV5GWr6xNf8IogJnyLXREmX30ouIopBL/1YhN6A
I6UX2umL3Te5y3CJ4I3cclU3jBL4Kg70mpsy1HyeFqvzixXmfsx4Wd6Z0KifNVuDOxOmXNh/lOta
JqcAKdPXSkKEPc21MFuVnlrYGy/hiw2zjN4+J/kj+iYyalrYYqdbZpNOJvjnlHLSBpM0Rnm3daig
kHCfIpGcTnR1m6dHgWcnYVYRYMfNJ50ctXY9ii/I46S7WSxqrT2E/h7/zpI5YVMglL1NghX+gIi4
+f4vn3k4+shVtL5IyPyU7yFGf/w/xv2DLEtogiBeugE2c5b7DeKaXnuVHo01ottnonBTS/DmnCtF
HfIj4QMbM3zTn+7EUbNapfDRwr86xy34wJZjCGXbn2SgdcACHR63FDPiZqwphXQCVdHX6Bsrzqmh
O015kz7kFm75ywN3nlqtGCMbcBaJDj4UAbdwL2JSgfLeoCF05bb+Ud4mq4hKwnOfz/rtRQXVN5EP
UeOmH6NMdNYFN9Mkx8C4ClHM7iw5H6p2pKUomqYuM1CADLJg8mSWXXk0AbGkzRjG63bEovpvCsCa
wBvxZ2cI+t39qRuF8Q9c40Zj9KN/YMrvL303floo6g90d6t4s9E6rWRRGRD9Bv/a3I4+4HsGOdke
wQ0cxjpmjmOediC4zi8+PgvmkBh+YmFnsP5ZBQWfMUon9gelm4u6tcyzhFv4JL0lmpH2gpOwFC9+
eZEsmwgmV0CylyZaBVGjZ0eWcULw/XrxO5P2KR3y+1AE0UApHa7iECJ4vlRGdWSTZrNWwHARY20P
pGaRIzOxqApKh+SVXfXR/ZBSvPwecjKpLlhiddoSm9he78O38C/tQ7zkTMbhx7U5mAcANpXQwb6m
5g3R3WK+4EYYIBbEzZrOOe73ep3yLdLDsLeWXphwlENvilR7ScEYx7MLoif61d087xrDbN/gsZkb
bl547lXQkYMXySlgs2uMkgKDyy/LRjX/OBUjCTr+shFw/nSPY9tDXHlp6cH3hQkwnZEfZ6uaMFYo
wHWL3IcI/cEpuk+7ARRMh0/Zutrdu3TKskngSC0L4RQCv7PtGjCtcogfzEo6L2aiooD/UsAjsV2+
gtzPoo6ZFshwQzsCcexMXoNfnhFsdDhBQlPF8qnqNXgbQCC/qkPKsIEVTH28YQwNSBvLf6OJFsHZ
JV+HfMj6eq1Yl3gcV5YLfiwIiV4Z6dAks+gumNyrhJZYeND2qBdFy9LaGNsuwfpJoTIXxg+eAzYF
nE/AruUM8cHY1Q1f1+ygzzmJWjQnEU1AAPFUfuMoS1dWk9jXbiev0VB/QgPjbI64mfDWd/eu+sge
jqO5dx7ofK3AM+unUKVLjJEZ6lYaR0FVTwWXFF4i8rPcCpglf5Y7jAr29JrlveXt9ZK4+hKD6y7v
zQ+9IN337grj62H4+70zdBVhhI7HarsHFOr6XgkYPwSLcensdHEqtEHn2HVGI3+vyE/zXaYWH4EC
wlwu2UhTPo9dvnbgAU7BdfTNjI3GKCxA8ASYEE7rvYQnUYAHZ5A7jP0/YG2Uq9t2+uGEnWQygiFr
nfdAT0yZybO3LWpHC1lU07kVhFJQYBRpcgMJ1d+BleyVa+wvgT6WbFEKvrBttGtvuBQnprMJiOz8
91NiMzlllQM/tMm77gdf1Jz7/v1Svij7udEQ1z6s6PajkyzlBqI+fTvTjhKCge0REwNU8+/gSpyZ
UGHJGbMnVi+2MtiEkPmRpJGte1TDQ5UmX0nBDpuNgMlswDOpINYCgkYoARry7sAVB11hvG5XsVgK
Vao6TlCjmr+vaUdz7+cdVOuWSfkcwiE8BT2h/LtSL+a6pJYvwq0zTTAr3A4AL3P0FUTgSCUylipj
QRzVD1lIRdrCnBZJ4Gl69ixBK2t/EDFTe4Fvs05tBvYM4VJ2YQn3iTJoEjgJny8pjNdr4qWWXPK4
sNYjXoJsPKKdeNtVVD8+z+VAg6sK4J2bwostEsHqki6mOXsvP/+L/mMSHJpaPCd8FvifeKJwuzRj
Cn+C4C34AKAz5K072Lrd662k7KZlIXedTStZqXVGVShPu+fuiI1XZDpO8ob0JGYjzSd8tY1yiJqW
2NhSgRu11L2w/tOOTo8D3xeuGd/nwA5j7X6dXlAtCWiaqhwbGLngp9kGqbYaB+kUwWeIlEyiDN4U
dwnmXYkq3St2HclT55VfSVpbtPFWHI0Bufjyos2NOI1HHJ+/OZnS0Oq2LXUe+ZC/PV/I5s9eH4sU
OcLLZNsBzcNlrvBTf+cjTDdeA8l2g3ZX6c3sNFwQYoOCjUY7CYcwBgBveb1DTDEc/XIWWuL0LNvl
m1pboCmWCXGprpzbJw7Y+rgg5fmCANq87gNfUwFbljpotzfvieu75cpDdqtbPu5UUiARFC4RRw42
4Ic0t0d3ciyluhmmQArUtSzkHAdhbSDpA2XNZXEl4R1SmjxL5vUcTm8gLtHT8l5vr3HH2sZRjHGx
H8QsFQ4gqIzfKPSORic6jkVt4mbVu4DVe9/JEPv9PvKw8es0+TzJi6anioLselLH3kkdE6A6qqCO
ZNKdWg8qrE1COvpVYDH5aXaFb3/k01CacOYMyNQAT2Bk5dI3qlpZ1aYx8y4ZIQDjXWMnCRnlDR2S
XsV2XeNxqENx+cIrsLySSjCZFvErd7W8eOBJ0Apu4BxIT4aN0EFwQs5PL0LamSqN5BXlqVXEHfhc
n1EjJrFA7Jyw1euk58NHV5lGOmNtltqcswGUS/QP5QFgPGX1Rk/f/9epHPyq5ssYinbMxJXmQ5UZ
9y4Y7CsPqL/gnaOyxe8CZ++wRXEZLS8mh6689unYaOtYc7NKsxpHBMP1xDy0m25h1p4ehDqzeYlK
JcFHoB/kyA0KJp/DPS4LNWuB0NkYA5VefjP30K9WzvrSP7NUvBZijdN7btr9s/UIY1RVDeuL16ac
qIxMy9BBJ+dCs9lFFwi5GhnJl8OsGqXeJBV4TO8MCOkeRpmVrK2ODGcokS7cxcwuQN3WcewlKa+L
VeLyrAouyXEJantyDddBQXq/9dFLtpqJuKC1GoxK1T44R3c+BaNZ+ry0Qxp/fj2F/00LbvYTorZs
Sj4+UvszedUO8a8FRfhvOg2jtohaPH70UPhBN4OuNQGNvsrqbU18krGBL+JRvh4S1USLV+PAKNRi
AWUZIg2mgB6GJTx/O+mPa+t+iiGDLkZjR0dWukHtUEV23NGAQK9xXyuf1hZrUFDAu6OAll/cLZQD
zGeHHt6WeCUwcyAsPtbuXhhG4xlV60DE2J/rjNj0FB4C2ImPdZSb0D8XDKm/0CXTvT4zK/uZsniK
BVkqSmUj0YRHC2mlr8f4Xqd/mwUzXwFiqneM7v+oUr6xmF3zZdy96q+Y0pvZc7DnHHIVAx6BsqoS
X+KsP+d+H9EGYuoUS6ZNDq/SgaWMMvnVS+JW0FBCSAzm+ZqYtHz1MPBo7sCLE5KRz9Ix1oEDubFt
lsIUl7Er1/UyZoORif95aAzHoFSgoKWBvDtOQC8aUwKu2LJExNEGr5n21S/XoaMbUNTXTP7XDwEz
q63FO/NMYvrf2Qe6KfDSedddYWMu21NTQVwkt/NgzIDxWwzNNLlwYW6sjirEgzzXb1DhozRdUcKc
o4RKLdyUbF8QdYH9OE5DgfTXG8abFs49ZTvCXIVDOIiiDtxCCvluS8mi8+AtiCe8hYdGRYWqdftJ
/hpaLKXqrxK8TBU3UEMxmrrprhtOrwwmfxJ7X1yxooRNinoXeXcT54lNcA6Wj1cDL8W3+Urxznj9
EBzr4Z6aKrCHyF7qcggCrQ4rH1u7gigLOOcbazS0q5c1XJbPeHmYFJDLJms5EqnWIFECgDr8qEB6
QLGNKBuwe5IZaT1Rhl+HKQ+o+SM7tZu/oQX/TiCuPrwBDThkVi4l/IjQdLG+MQhPLI8Au3BRG3Lj
iZqCx9U5oletoagACv3X7jWMhGPckZ3jWL8l2x3Y5RphGIKacL4gPPtrVA6M+1HPDzu/AkTtzqsU
vRzi//PwOc4T28i/EQt/kw01ReRkVI47NJKRNS24l8E3OlLvDzB3P9olSgU/EluQQ3DiafB0IWrc
c0USieMl63LrAJGL6TdvOmLXBahL7Rwq39+9NrmoqvK49ThbUP12oGVKxauH9oaMMRJNJBAurMZ6
P22GKq1sR8Rxva48nr8jiDUM3ybxjJO3hq4ug2ZgN3IDNMKbarooQnGXRala6cBY0X6vn1ON79ba
fw7QOqmc33kir5Kv+fISGPSJHseOtAO8FO4/DaEC9qMNEkkniRmBITEG0jMcIDGsqTKKxzp8XB//
3a6EVFhtmg8HciBpIxWqgNHQ4xnPaQF5EqxLxBuuJNvtcee3HZcIXCbpqYsOmC0hQH151xQS+Xms
LKlsLuEsAB/+04Ht22iqVVd0OscVSRbJdsYJOGYvUpU3nWkct0N1NES1jG2LkKrJFN0HIl5yyf1i
smx58WP/IBuzcOMmD3n5DNEOm55PfmhaPW+4Gv6qy9m2hlBN3800vPaGdej8C9MWyohrb/4612JI
duVxOOrJot9IwP+egp53CUp2dDxvabJL70RD9zezt0VsJWO/Yiu/kvVC2j6Q0wZikVaUZ6wYyhwi
84AxwSgMWbwXge1+5ecXMEuMJ5encscGVBjE/ZCa6ZYmNdjf/02YLE0HzAWu9+JNfOC5rmnd7EU6
URNZ28YzDj+OM8KES96oIACmKUQN8BZt0LnT+fRVebZcVlrSFUh6EnOzHBr7/71NkTXkb8rSXN9r
ziyJcKDTiGtxcMMaYCeenAnHfNu7uRe4JeByFturMcNWAp1AKEYweUKjXqb01ghNWOvGzmdF2JGb
aNxuiyDxTzeQD9QSevi5uYokdDzEVmWUWqGi0jp0Gc6kXhZwCh+glSHMKsYAgtFMk//wi0+v4Bqm
OQ8bP45/KP5Zmmm2M0tOlxUyZiDhrGd/8mC0a3S0G/atZuzEkZ2GjO6aNR2OZWjWMw7NEJlalUJW
W9r+OWA0ycTNbmKKo0YeM13S0zqucLQV6GIZg8h6d+EUtIikFQclXdLX692LEO1nl0igrOr6E4aF
YV62uhIE8NIWaAdqrCNPQSsF7iueze6za08cXfkrCrrszLPqyMK+hZDtYi4q6j31Pr7n8bL6fSlb
1Q0hG4zMKCRoxNzXZkl1jLwTT3WjXen/dQv5R8q7TPy6oCsvfOvaeJ8JPsYHdhN6OzKWOBgdGFIl
CAFLKUsRkGX5uWEIXxZRi2LvICw2ToWUN2Af8qoK8JRr30K+J3kcypR7ZR7ZBRzEUwS5p88f1+DU
JlCiw4cIE//QIDmJN/2eAAgHYIbD1Ia7LDoPNdfbhVcTxILnDvaIAZojzZQeSUwUveG8JudaXVWx
hnaHDrl4S8HePth2SwgxdmQTTBIFq36Q8EZ9nTJ7xSphu4FbWJ4dh0YiV+M1z241Hw4z/N0ZyQAf
guGrM4g29rZDdHPmvMntIuAf5fgkMdM2iz4FzDxETCVwj09qZxPEonghuH5BP7zuNxotqKerbWdt
zTeI8Zs8aUCAgn/FJETnH/aBvjlRMWlc051jnEoV3/RXAA4n2EvL6oOSAY9WyHnAm1LNecEbHvWq
6XARJ06GbTQL0GlPH6oV62eKTRDndMnz3ie43BfE0s9hDaNwwRu9quJ/iAxvN08qPuEwwuIXhdu7
9qu2Q9FYDlCVMGHscwmrTVsSNFSLLhtU/Y4elM67dRBWvRuDDFq2Gv+HMHqG7JFzw+nLs7VUpEN/
SKvWbs4a+E/jlXTwgpzwQFIOllEbWaFvFqHhTrFLoZkm83EmlaV2rs+IevPVHOVuqCFWma3dvqHZ
DuDIL5rmuEk5vGj5qL50IOyrpqJZma/qY5bRNcm3qyoCnYNipGarGACBOwUoGVA0/eDxbpLUIAM+
EJcW7NcgD7GPm5CfrRJRQZirpWnJfCNXTyuytMhYk0yNFgnEjeRjqYs2zX5frCqQG7MyJXvANaG+
2j+UIq64xZAmkogO2tuI9clkYBeRKBrusonan8b8p2nS1MXMwnlgH1JDxGOq2w36rKU4Bxq8wjGA
oogkQ52Xj183uGcZSEGuvTgcgHuzuIp8LvFLJGzLk9rsv6JiyxFPkG1TMFnNVEAev2JvPEbaaqnF
LFnWw7c6jGMquHJMHE8KvwDwbsQzc68ys1zmzS/kzjY5YfLTPtbFbIKLN/iQJOfEX72j+ue8/9Ig
ULowUAza4uLbNnpoTvjvwp7Igva34iBm1eKs0D7siepx5HOv5vRYNYK4L3QeB3MMJZUGphkXfbna
CxhUZ9SaNyus31Oa6iiVDgKPRzcMkGDjFDh0GiO2iIbKmaCbOf2iRu2yqOSWusV/x1W0UXuDUmFk
oROCHIJuttS5Sko2HOqf0k3UKWvpm7qoWLEyxqAXpqtgfYXS1s13EOXFyUnQOzNCJ1nxFJBFqCBx
GJhlGOrl/oefvAuKfABbq0/9cLpq5QM6P6XMBltH8AHGu+2dcBNVUrKwWE0fU73Y5MRl00tyPMn8
0hhBDSBolalTJy0MQWinMAre4N1lckPh4duakyeAgcyDo9fbUqdoYaYznhwYXFWNK+2H6h02elhe
OQ8mSLQ8jZMWycYfVJtZ59JhldNpGwaKWAYM9x917ck0rjatEQ8Nb5h5WHDJ5uyKvCPX6lwbyDYt
4oONBbEMkIv8WxUs+dtP/13VunwB0K58WB7ZSkNvVqlxtWRKNa/GGqcS5t3M1EpnXdiV5cCXTqQE
4mG4De5ahJ/HAgjwEWUf/tOaXQIRKTxXCpgiBDOInEZ7P+w8JTNDmFtEHD4yPUOR8vNFtBRHl6N7
3CGnndBRoQup9gGSmYifuFPFSVTsO2Nv4OkLohfbX0RAERyh7YgUEpQZ6X3nzJzXxgmQ1nEGEr29
CRTCyTBE2KBfGIOtU6awxwqqgSyX4A1dYuuX4bF86EcNQwx2SbkL/XVTr+acfjukPkWiQs2uzZ6r
Qo1a3dX2BtnvZKnxKCuo1kSgNnMOPGTcr5SQ5g8IVXCVBEuDG1suHqkfSpg+40AtFkVIAqMSQbOA
Jwog+NyMcPdAMdTx6NnZyTUmgG4gE4VOgj2EO2hbP24W3v20fM5yCXCgmVowZUFV6380fAK7RdQg
KhtgOHV9AorTYZjm4erblLzrs+IaamTjbJDvJosX2aQT1O/M33xwOn+AbxZEe5Jp2PpPSPOgMg/2
FaEaJ2VqlljEeowvoajIqahOb1t8Y8WOYqkKvygDUlpxlVCjFPmvq9w9ZJ6n+AHCn/Bj3PUf8XRP
8dPldJ0q2wj8QHJoitBV5rM4JNYCwuXYCbjolKFQMs2ije24B9iN0N3z6JFxvAnleK77KtIwWki1
JHt+MurxT+L/F17AGuwsFpGtk0HI1G0d04zrJP4MYM4YugWDBKjttm6hR6ts0MQpCAM0Fe6HuUMS
lvQFI9ckaBYelnzCdxbb4pbvv7HniGj6dIHthKilHZHDHZ3qiugCUQHBYIxB/VPtTl8U+KaYqTO9
uvYkvpBTcYz2G6pNxYVaDqkBY/xaRHI3cXkehl7GoI7Lqnwg6y27kwSM9E37bOWfBBJVPDzt9KxM
+tUeEJKqYlQ6i5IE3oCd+pH2hyfbql/UWM/ZV6iRTZXAQ9Z9pHGXWvrcfX9qX6b92f1rq6RyVVsd
poSpj6rFmX6gTcG/bYyhKrAD74ip2lIdz2fXhqJva1j9P5Z4MP1qBHHvytZ64RJ1ymvbzeS72vx9
rLnQkFvN9Uy9vqAPpIwOnVAHCcxivMfFphjYKnenOhqUdeqepG1EUUqKBwhlo5gWpayVFpKvEHSE
xihohtsiIRK3b7T2Y5hcu8ndRuHhV0UKGJw/RQd9k+FSd5o7XLHpWgDehyYC5ocv+KGPTL3SPd+A
o9uWxml9fOoJeOvM7F6ZS5Jjh8f/FV0A7o/ogfWGU+qwVUgrE3Uh7n+sz0hWDTCPn7EQQUkJa5ub
1ahPk8AYBg968hGcYERuqFvVFxxuOfpf59dd7McVTZaK9WqB/975R1mA9RJoEr3xLS3xC4JSmPdR
RbB9Y2qJbWh+dF05ayhAmq6CqmFMmfObK5P6LJ/M7pAlDhQ4Z6n6rVhUOOzmJQk0GfHYhjMXCILT
Qaq/BG10Zl8+TrNMPIvsGaVhkSTlFmHR0goAjDs/STflYQyOe4bAJPk/XWJmPHY9F2MI16cjq9qc
s08fkLXfsNdunxg8vkB4jmHp+1AyXJmhzv9WCJtK0KQjJVB20UFbbroH+G23qKr2RB+fPpNKWYnG
aR2+846EJBjvfZmtQeNPcnN9Qf1w19hOONy8BeRx8Rg3Va/Y0MYdDPPHWB+ct07MEA+vj2a/1QjN
RZhGH8gw6ybWW6YQVBZAd0WvuCfGY07QzLk1eIgcQ94TGTkFpEEKmScOjF5Vsm4yUC4uuLWZDaGZ
wpkRCKfO6NhVDs8pCF6LxitstEneois+0yxV0z2YnaCjiXRAYHXAxyAorZsz4DuK97hVK8ToVpwK
yswZ7l7C4f5UfSIVe0r8m/6tFIpvVPv11/+fuY00AHdGPXW0Xr+9U+H+ML2273CAUu9lzA/YynbP
mePwzf1r1/kCwvpGqID+2sxi7vDhf46Uhj1iJ6xAl75B9MDA+AL39nNL7V89K5BsbvNBLqz/LFXP
GBbkd8RkJMcvlh530yx/QJ/v10ekWeEXM2gneNger/78alI9IMN5nfVv69TzqUsJP1bIS5zGXxOg
ef/AjTQL5TBeRB7ZvYe90B3XuSch8Glo/XZb5efG9cj8dVaFcf7LREEXhxKo9sOhMi3/9Oe2iyC3
3nsGFN1SdCFFEtWLBnV0cBKnV87mpWjHw0zIP31j3YCSr5fZz8wqcGd65S3p29JaUF5V1bdbWewn
pipLtR1LWRs1RFmubaiTfomvvZrlYzQGDtbm7WtDQwQyRA/DO+WuFbUA70d3E0WGxGr22WRX+jPP
3l1omu4KEkorZxyqfo70yB4V7/Wl3xLJs8GoN6NcnmPdIXxmltrQIREDu+wfKWcg3gadkEcCcuX9
mD4mWu/A2ilZYSOESRwtneNs/hNcl4rpSp0sCLdD/FRYCE//gemyhRPS03keCeEwEA4B70EUrvkY
kULIykZAMW1pjzguiKiLHFpxP3Vv/ko6hZR45Gn/B+G3iMslmwTXH9vk6+xyQJ24wmorSYlYAe4c
fg83RR7UQZQabQcTLx4T6y5LklrE1qCOiq8fMQQ04RbxsvsL/CsviHbdvjEEC+1Cx4eIkt42Sqgb
Hdvbqll2I0qBHqNfF9aYJIALewEJzgeKXTX5qzr+QC9jxYlXAPDOo3XkeIMD9orZ0Xd+SAYj9iv+
XtaKtIFjfS6v6kh3cZ0KqOmcYDz8/bRgGbqIMlRD2P7Hcp3EZSFWeyVRVE7GrvNINzCd8GKIQW+J
VycWHI62dRTEIpXqFeZ/oJPbHJQcpluVxJd/YGOTnlb/so9ELTfBoaPwYe24Hq5Ml4uTH/8sxsTQ
L+kdlsLHCYwIPWOSposxooS0lUYHnZmc8jd/4lB567ZvOAnugVrrMyTeSegU9987fzosdqDjPuce
zJXXrJ9bz+yMDhTkKEhOZrej7j3y0IlhL8HewhHcONnXBeZRFyJn53UlIYKq7alGq7mlVQCIvHj4
jekfe2wxim0pN0m0rwEltDFYrhWFFij9H0AzEx0eY2tmst3kJY65eAP1alJmECxH+7H3C6IMWi36
BbtOYExXEYL5lcl9ojY7xSN/pzNMytlsCiRoHNFlUrh7l2o861f65baZQ1UbDdFieE53dGLPMwNf
PXp70bDsOxJXy9+xTIlnII8HvlNNq7teRH0RXyrWhMpl5DZWBuZFYHlNdJNtTMhGAieQnYQyfz8f
so+Q8JaylID3mMr1NQNPY/xBpXMw4q16nvFXdlp1bBk1SEKiTZptADH/s1AM2fFMM2C1/ETpV7gf
gRb8IVpLJf63JXydv4Nk8Z0rp3LVyUoxTI9h9NaGGFhnhYCMEZz98VsEAu+AD21Iq7QBpDlYxCVd
NVjFLq/LIDHgWWp0FlAne4B+bjhkdfjbK2WHk8BJOkbrJYouB3QgtuNCbiuI4VIXZi959nUXRezf
VGPd2y6YtmNHVX9JcTUGgihzL1SsXevWfNey+a5OxlJWCpWakAo/FLPSi8MHIMy2IhQ8DUcEM91O
opeKh6Vbh9BVplePkMxcloj3jVGMU0bpfFvu6Gw+pRmVOkfOUfyVs9xe+9RfiCxiDxrHHhbT/NiT
BIeIkZcyBXMSkR/nNZdmxJWOWfHhUQaO3gTViS1+AtdgxNHRzdzM+RFAJwtTfSWaJow4sAuHjKmr
Ys7PXLsovyy8S3bXvbU4WgekJBVO5wd6X7qRFpXErnRCsH3/LIPTfzS9JIKnNsmzirUDRzkUGSd1
Oqyt1jHqNEJ1/hG+nx2wVHWx4Ze59JR4cACpYdmJs6bxihczuiTUWMxmsK1CLMiRHC6ytgO16BV1
gPPW1AWFN8Tw8A4tasDpnvJxcSRdBASdMb32tx7ywnxRA25JchfrVDuj6KtR1UUgbqz5H9sWtzG/
eY5YJaYrT892MfvxZpZiOQ3AnmSxL8ZOVyQz9t36QuFeWvs5Hg5RXPOxv+WmyNvrPzebEbSlYnE6
fXDETSldAte8ukJc6FJ7Qf0PurTs+1ki/MGKMtkVwg9wQruYl1Ffq91ZwYFY9anFGYTHGtdBzOXN
aFcZefIBmLXPlrWJeUpfti6mTI6R4Yi5zPC8q+/1DTvD8Z/xTAc49xK7XVqf6ENcryj8Hx5u0udj
Rfim00wBNUHLWcmQZcPBUJjAsObSUHlRiQ1JJ7j1z/hThT7KX87CE/PKpjMrBMlrAjO7yQ0alHTb
Pdu3OTD30FTZVOdYNe8v5qBMs+p0uQ6h6/ro/rsSDL028IF59xCT95CefEhI5Yha2ZY1iJ2AHoq4
2d1hHXNmYXg4ZjEF7LnjL1ESwzDeFd2lZVacZmeVS0Eg/U26pr6y4MKjdxr7UFmTWsvAO9gIxth4
oTK+YsMvyG4xY9b8ObDjfNf0uJrKLQ1kQ35Lq01xYXodVMeE7RIeKF72lw0hdN64RguusE2PKE3F
N21WfprEaM0YFe++sfy+5/ySynMwBluHg0jExYsMOYXDh/4O0s5y7h1wsykIwQavoyCunz964J/4
TYZ/S4n4VOijOPFf8oKT/QgM97+5B4dSJ6tWPAFQ/Zow3mFJA+qHeEk2q+Cpk/D1rwihJNl9OcW5
CC+d675jSap1PhEahqGScQFJeL4FR/8R0Fu4+BFZrwR2PUj0C5sWA5y9E+c/gW/dOLWGJE8xFpSh
dqzhSWKpbSEywSBSBXnBQcB+YCY6QyneKaNReFTnkRms1njzbEDQlXXZbp0egq3Umjrk3eOAhp8i
8wL6TgTwr3sZnNNx4Y39gknllieoNEAFLCecrV6PPNI3txsRVW8b1zZO7mda3Jiv4YC4YxZLADb9
mNdBbXLmeioXlFsjDD+JOKbVLy1GDSoZ22zTJLDFBvZOsLafZUzjMDhW6NF8R91VgpiTbrRU6rLY
wbmW+bcLtl3cyshtx08gG52JgMkhj2OiYP9ajY/aDQzl8yhrZFYLch64m2z48iVTLcE2kaFpIza5
LMcOaJRiRGrJyV5Afs7bt5c3scdXLgq9OEwl9z0fzAYt4YJYDXOY0ld3cY1MR3Paa8ysrfFYv0/t
fR7v8zZexsD+1M/RVwigO7aep2hNtczlBz4S5dgSUMFdkzdCwDczipqr4uMGt0iXV7/BUXHWqj2U
bdVr1AYCWRIZXhNo3wEYzUlkItSjQNg5KBydI2CsPa5Vmxl3kHqPT9K+1r5ziFKQrIvBP0vt0nrI
qMgNFS73ZbyUy59BuPSwjdKfoLxUrApOO0BEPvmiUM1FSerwU69FxiHpZe+CRxxJ/p+MXKJtEuDr
MORIci6KJ8DPFGVF9vOKgECLfZterUNRAHwit3oEGhcn5IuXGkxnQdvlJQDdqiFqt/zEOLY4ljKA
lmfxA2R37KB1u2u0Dzj2ajOch9CnlQ7QOmlsF4TBvJirMWRHPeGUgRoLHWWHcRyF+89xBq2MXofC
VVcOa03EYo68SYRf6jkFTTYefCxo7Zf2lbsLaaFoepuugAJ0lOMQspPtJI3YxHYN9VTbJIeRLDEA
WFoss6ajMeiqccLolc8/5ulNS1pB22/k4rg/qFYj36d2pwfPUIAd13ifI0HrlIP8SJjhPwVg77AB
rw13uArjP5c9ZEge1EuFI0VhWn4tNTIVx7NGt6/xO6kuqJnrQHf6aN8rvW8lhGAgZAND3hlGlzAA
k4TI119R1v+pvnh+aNnPDM+vG1QMUbf0/Ih+WnZ3Fd6sgcnJx8OkIiCf9qcm4WdekeaEu0cWFYTC
QHK2hAw1aSBNy/4/HTUsHx7oJ1KR//Vi4DyTP/dWM495J+AfkI76Yv7SdL9KFBw96e8RUizdVO3k
wDIeUZrgvIRMrmLvRMcGJxzB8ECmODGniAABO5wSM/dQXcV2IEsXngS9VfOP7h4YbMuKEM65RYjF
BTwWHnf/2LJ/yZlVseYii/L3ArMK5+cUEIHa0lUfdd8kfIM7ibumQSOhzgG5O+PP7AtQLLQlpMq5
RS8KEBSE3ku2fUtzUAcxSYj73ffUQphY9ZNJ6Rd0I0/zewpdvuCm+ZCbnhE5bB2NiB6E2sb1LZmy
8XX1MBUiwtMizpCRuKEvuiLB9uOrtZz6AajtZxQDRzGrgXOOs1p3Y2axmDmmRKk/tofjtX9v7gSI
ovfoAv2rbYzjCEd+faqizrjtcfnmpZKzXy7c4X5Xuvc2g8WynCG/thN9cEVjA8Wgur6sYCtJojiR
ZMuzz0r5fs5X4ZkJtEEcY4FtCWK8YmskuMBAF7JLvoon7kO9V+sQ3p0yNY6BHPveg40qbiKhrPCE
Ewagw1wVdt7ktNJhIo8HF9tZ5M7YLeLNb9SFTW4RxQyIyR2ixeTpk3xh4QCIrJYOCuyeuLwAn2rI
9t70qrf+faKwiVqHoKF1B3UnbpkYaajyLzuSJcGRi/EdArUh2/NIYLjJLVLRToOb6IttmsN2ntY+
N7doyOqZhWKjacuQXhXnyczjrtlBT3bh9gb23vlWK6U2hnlCNB5z2tno9FWrruwO7sBdkmwokeW/
xULhPYsZ71NK/yDbDIxnRKspoMjzb7UZQY2UMu8XiUu0OfwZayu9ZIhbdHmrOA+ygl+GgaX8rPjC
V3Ayg6dOT4OPVfFenRE8NDYZrB1E/bBTq+7kF+ST2DQRYWnYna5l9RqlA7SPJcGeSbYBalG2FiAR
DlUidtQyYwd3sJpjLqXzKShLw3hUXy4VAHsyxtANU4yQjZMhdsgRphRsrPXVimAXJM0mzpNWzvHE
laEdXw592b7KWsYTlRMHWXMlWtOq+15CU6hfq6C2mB4ihniG4Bf8wA62B2jwdU9MXVq4KlpecN29
55YgSNuXEZXcHof37uFtjI2x2txsWvF2aFygzW1Dt6uNGLVFbpGTGIHFudF+yuqmqqZPe+LRRJBp
sl0tEUublQuuw+E16rndjjTrk0wDq8lw/5I9bzM91Sbed6g0kAU5TPkt9sufBCZD2v6ywcInhEQI
+dcaBTzM5RbHjTVP0YAL4t5kP1lR7KTEAF6P/qlOkkOhXEWKhVSOQGJnvc7wgo5UfO9vriS6KDQT
gDRfa9zI0HvRXfg8wmCI5HTfh3Xqsn+Cs0/2dad74SCHSoCinppFhAiOQrjjwS8VkdHgAqLI/ncB
e3uGsBsL2DW63gtg66e92cS6QFlLYOoWEit2B0xkDWXqeVC5ma+nQgo4NXOdtkGBIceFiu+sxQM1
8NBWLTOvAiX/aR/vB0CEj69mpNLK354L++sOCsafnNnrmiaa+/cQoM72jbDpaVEzzfZT7ik/NAOM
VBNMterIU16kbOJlV7XcwKVva6LVZzJjy9AZanWeA9XVrePVkkIKW7BnKegitmNfInZHdrLJ5yDw
6klOvlRrordNBkuhevXOeGGFzIv0kB4Bt8EBU3hAQ7w7co6afUeZgiVKbTs6rltEu6/29IdLSVQ1
2U7YX0an4mjJodWh3owA535hNilAuKY5NSkvcPrStnnkleNG14N8rHnmu9XSvVeLUtARjg8UYVl7
ahizkTcTosvlqMBjJGr2LcI/qnTrh2LDBOGWR6e/1vfARPvp0ITcs6/yYG2bDRHlB8qXLMGaYbel
KVQ2RnLUFX7yd6/K+82+lp/TArToTNOGVQB8AgxIgAG8Kh0D2X5mBt5smgLJ/ittfeFR2vqSiGAZ
gxrmb816vLeLNaAlTpf4UpN0I7cxW70Q4xV9vNhjN1uhCCI20tF5aTuWc24Uc7rAGSinJGGleYt7
mrHMomvK9tZSnbafBTvOuwOpY5VanMuAxWtWtm3b7jaQgdOoskFoDem6JPVmlSzfi5Vkh2m42LDO
RFGWUVUUqaR2VOfa8H07I5Jwj8NV97Q0u6RfMllopL9GqS40CVdY83DnJK7XWuo4LibJZrJDLckL
RdK90AS4kEZwA8gj0DOCUtGDniu6M93MqvegVokq/nEQRkvedFc3xdEoZzjy+V2Z8UB/Adwl6n19
KwAEPhsgZhATqFYC4xgsYmdtovO3Il2uv5MmVSIB2RABszVhL8KMFfeKMfFT9jb7bcikDJK265w+
yb7xuopdkOYeQK3zbFUqg8dCDJ0J5svLuBvqE/ou64zCyvFvubd4F/CDOquHS5hr+QYuHuqe7uqb
pjkHAQXYfmbxUXDTgOTTU6E2VU0XwoCyFdVYFPbrgVBCisbtu8hOXXcTIS6Q9BtCnNbt7iE/ncE2
+NJXzctbNBzxKD7HSHNiSHhVoiFSMZFROdsNFZQPgC/wMfhOiSSf777RtkRPLN/6r/wvov9mPj/U
V+ARMQktDXe7M9dQ/55D2vCHAi+AYLsdVjf0IGDlU2mrFlKcSDGP7y8BqWED2wlLKCrc3r4p/eZ9
xUumIAhYm8iQ+7tesKaHVDLWr5Gz2io8pCkoB8mGbuKGrqs30HuLnXBd9Be0mdZMNEEbueeXyO41
22lNIfrq4cfid4hVTYDbgPPzFWfkVPRDDecTV0I6X6Rjp4IqS3RI0KEQOGtWGXL24MLZFReAS6KV
rqcv/X1S+AZ6iXtsGZXeP/A0g9df6/Q0/Yuqkzr3/pM/1YTrCeOgMk14+KL/Pd75YreQ05+2mVp5
xssLwteWAkvpECB3uEVJW6WwP89BKoScitOz+Iaddc6u7HW1/Byr1B+orfAYOittPWkiZwcFL7MX
7sVbqTVUbBcEyYsnJpOGbnVZ/gmqtV7TchQRjnGT42Q3ENpj2y6QpHwpp1o3cBBSWniz0SUzjsPs
AS+BHH813uQsPMXozBSAZabn+MQB5g8hVeDsdPSIxQPgS/DRCWw9011J0/hYH3wY71a/cPTYKFgL
mYlpWvQjySV7Q/semQscD0Mzswd5dmEnLEvOQzJTkSpV8DTfBmZxEIlbzyYL1PLvzOBmAl+Abt/m
gIC797Iws/6LAU/+LXO6MHPnQYsQaj7bvk9zu6O/RSygVK6B6RrdEVrPJxjZbRB8VXumS3jCi+sb
BZMXfSyp+LbTWxuKSg4/pvEE/OiGkCreWtsSF3kQqHvqcEWJNi4+e/zbxEUbNlRQ/sAkVU0WjAAj
P+Bs3LeOIunKUwS45kQITxawtzd/44WkdqGfj3R+d+3LXRyqlKPUoJWbObuZf7CgR1KGI/Gi5z9R
jS4JpzcFlJrgIbh64JxLjabVOD8Y4ROUc03T64TF6i0cBNgKzTdjVb/J0EE47osnXm8FwsFfaTEA
B2Y6l9XpsgIayl0MwRD4wuohF9WtpjMrNaZ8iveeH5wC1pcLFJlLnVft+gzvH40S8T1BabpAYDnQ
uBQS/MF0oqXJBXaYeBuHgbm1Lt/DmT9D3Z93usH9hWjuKKe6uQt9C3SImuiymzLNbB3yR1trKrJK
IP79/PJQGSoAzL4OvNCEVjlu9xuSI/FQe81zNNogZU0vwj6MEFisBSPFloq4WsR/rd+ihxtmtdsP
3B8xO/eGwuSRWrNnFEXvdwtN/2cpm+3jN57hlnht+IRMwiVj/TmbrnY5VQB6dBc6/+VOop2J6Xtg
u18AsdaLc4j9/lPxjmzL2LeA58o235vqiUkf/thdPRtFR75TWsAauRzvzlkjZgEjVEm4H/ilX/Ek
cDBhJyVn7bXJj+iigQE95h1farPmY2oAhiYfVzGcxSOGE9yjLGvWGbCZEjhozgbecCDHsOFsvwnP
e6uuAlO3e9qCQw3mBQoV89VkjTKDVetmNKklAYhUpQBgVCVmo3XdH5Ww7aCOQ78apk7J61Tj/CED
S+VQ6+lS1MxWdckpqUGg3UfwspGjpU0wgqVMNbyfvk4QR8Mid29vv05gT8axqswz/UDmyjCA31gG
kEewOiC02UHtQFvkKkiHTwG0F/AUoJ7EfxuoUzchwj9dv41jVHItMK7reoPxgigMSXGn95gugm9E
ar+b1dVgruiXTa2OCr7q/59ZaEXz8cdoblywzXPEOsUX1q1/vNpqEkhXczERVRGs52ArGKU6sszM
rSxXdhv0v7iegUwMOa8wvpIFpWm3TK53RYO4fnJyFKkJKdyLQz0jqV8MqdLCb/JKtOtWEEasHnjH
fCBDKGE0wHk4wq4emuiRpTxyk37bNj4KPVv8J+7oXWYFNN+ofcMp4TWVQeyXDhcTKBT2zfTmaXBF
vvvqdIT4YPTqc9OYvbUCwP6vrGwXCPnOm8SIzoElq9598YXIL1cesmE8IDoua+R79uI2EB2Zw8Xf
/WpYXHda+RxapUL9gq6Th9n2Q+qGvN5p87/RGtcjqcTi3rLM2o5mtobCOWpUVzQ9P0AauJ0+KJj1
sqSU39O3j4QITFzTU9KHRM7zyewxwPGuviPusd3/4vXm15J70EnE+XX4MEHBfCRvwIyg93I6y+c+
N4HUfQEJWaUi7D+Lm06jdmVDkmGS6kgrLy5+t7au0s6yhQzOq3x/RGQq5lCPSCRZtbmK91WGTnGM
OFrU+PC6SzWywhsA3psP+v3ZVPBv1iQ+9vjzNe6zysEuz0Rpd0tALc+6xf8q7pBgxIIx6/13IgZD
iBsObw5uMM4PuktZtWyq56Q/66mKvu73pgU0apDCt2Glwlr+HCxzG92gTYxwNn23Iorqv5DoAXKa
0F799y0IPyQfGQvq9Hq5wANfUToOdFdDf+Ng9XAkmTfMecZRZ0Zq70jh1o7WDubqPIg7ALa6sr0c
be5Hxxnp7FI28TAj0+ZJ0/4dFwISVzu4226HLD6c6e2RGKttlB/88cOK0kmtCOUzVa0DEpxUx3en
dGafVPIOWKbVr0bttHPgP79zQ/SiGS/hsn8qrylgyWYMxEh8U5/CrVSIgTSXnKwO7tOtTXU1KY8J
hbDQbvConw5iKwp3JfqAKQ91Iz8AjX+WRbqA9RIX52HJ99vF7oNIS9QZSqW+eDXXzfrTS4/26Muv
5V6bN5eP3lEvt0xBLF85xY/YfhxIl6t+AHlcoaoM3petIwK8SPHpzxgYprUagDIBOJwmmTYoAXIo
KrjqEzon45WT/1fsHTYhrl51QR9pUiHdzEsXni4QbGpFJvJaGevwFsGTJAitfR94cOpbdX0p6w5T
KfYDM3Wfb026YRVYBu3wi4Ran/mKv/m/7TNddZKOZpluENboVEI8plNNezmF3u1nc9SFfmObJzgn
Z4iwpr8zqlvZ/LVbID5Eq+N+fe+uRIDovaWG3qF4cjC45jJSVWr5eghgFTmknmZyrDeraltd+01K
ctPeizMggjk/bvH+2T4sfVU9mZArBoPxbE6j9SoXWa8OdYnK9D9tW2bUq0kjkhMZy52rM1H9BHw0
3bNPsZDstkIaRA0giKNbcwSmFoPogcblv16mxDy/zYqgp2ElwOgUw0qJis/QHestl/d/ciBxJKqB
NaDGlKGSUwBK+eLrM1Mo7cx4V8WaorHgTcwStn6eGMEFn5qjz+3NMYGay02YlTmLPpxJnVU/MBuk
UPpxIUtpZMDanSqyvmXr7WN9HZDxJnAmBW5rJw0uX1vcrit80pkxRJ6M1/ksE+52fyFbh8oLVjKF
wTXOrJ9DA7Elgl8sOW3SN6Sq9+qdFPmKvl2G6tj4MSNpZB754n+aByh8pP9btAQqMx0ccxXMLPv2
a3BI2C7Uw79TDijhHTpLqS8wglHPXF8UFz1Om7q/Ag73DEfaw/IgEpaQakxogqJDLHPB2mgdXe3x
R69DyNZrFkn5i85Ddcnj2K3RLtFYt2W9pC4Bh52SdpzMl/ICIuul2n/r9+lreAN0oGb/dO7KrUBD
9yJGVb0ZU8tBydW0mV6xxbuonaLAV7u06zEMtj2dnQPHrG89Ol8DYHg3yXyHY3YNOMycRiDKb5Qa
M8nayJjXD5e+dR00K2XIWCvH2pbSiEJVh7N/WDAxsGyYPPMgexnG+rzU6zbOQF/+Q/hfyfbeOll6
GdplSuL2fql18II85ir4rLxom2hZUM46c5j/7lwcs5UktOHBHHBo/S4j8DT5WoUs3n3HpyFwxUfm
sKghtK3ydnxCJQH0+G3buYYoiPHrSGKwVE0um5FJJAM4IKiNqwkCWzDHBKv/vnjA33f7crsb2q1k
eoeQnhSek7zg4gcdvQpfDNtf8vrusklRWeTa1GCrW5zbiaDP8XPUV/ULUD9l7Xtdydb2TW96HRyp
az7lcihNq6cAkTNNmuklUgFw8+x8KpxQaFS1i794q7380nz8P6YAVRmCss5CJA2K16W22cWMBV9Z
2cxh+TSye/7ixkvWyguDHEDE8CgEs/I/GJWeCbXDv9x4IsXlfMY5EaaR8n3u5LYeg0CfH5WAfOUg
Pn0u+1/sY439GxMMMjOGNsdn/2WgZJkifE9H1xMgJO2JjBKwZDZSkUoWlUMe+MrX5d2K10HST7p+
Tap5f1DLvJU9gFKo6rBd3EwR8k7gFVrjVKS3j3rfQ/c6E+AH41SDDhg7scLgSmvbNo0BjGJl0PTb
71AZshgKfHWeIrW9jBNFAgrP9330GW+FIwhO9qa3D59ZgNwNvK3IkoT9Su8tBrBdOAliBuM6+DN9
2XrY/ZlXkPDsQcjqm8uZrDVfKI94v5+KoILpOcs9XhZBeCKJazfzkLqE9XGI20hB/3uueKYvpBGR
8+SBhQTGqSgn0dYSHMnQtW9ydWJgyriyqAgCDJh39Ft/rkqzown80BtVsnTPwVetbrhAj/sGBVIA
e2Toa4nYca2CDSpZy0pfWg4Q4tab6RWeMDRLIZkk4hV7nZG0heQ9ngeoEP/cYcrxsD1UPZzapVCN
+7yyRlHihg1mYg+c7VjzeqZ7ij+gFzdgSEXPtYHlPJCwq9yeaVhECA9tBiHdctk4rJ7RgQ6O75Vr
PDc9NxFOdi+l09ZLZClekjZVQb20BBN3m3LiP5uzihzlQzgYYsa7a06xNeojGua7KBGit/ccgzQN
+8BzyYbyD9Sa0GM4T0X4dE/1MWa3NCbg7qIU2oms2U3B8UcfFQ94iedan2u5fpS7c7jr92s8mL95
+VmyqKlvznC+4ib3Qn2N43JQMvkB+LC9NPTPeP6lGnh+WwUvgA7KEqv/3qWpaAtE92GMQ5d/ZlY7
wdHtisMerROfeEsIhUzzc6MyhRGoTW78E4sw75Paz6/KEIlkZIx9pQkvueV2QuS7l1AAix9x8i+4
PViKbNaSu2j1olv28yIiZsp7k9gsWPtS/STloXUHE5bDd4lr0scIcjzEjB51X3xdrf1DA3CkDnv1
EpY6ppgpPaA8+jGHfo5i55ngW1Lcy0cLScQBxAzzNkmYa8TA7Xf/Asl83wzRNhvGfI4c5tsK9TRj
mfwrRNKukOBMrM7aEtpZqXFlH4mgp9l+5YmfgdrZtPhmAJTz7+brnIxZIFK+XkUX11b4iBEIj3t0
Ob2ng+4fHtlR8gKqxD7/Jvyv+TsHZs5AfaH7Fn5MPb6MOA5q0dOHHtiuvOsi4drFzab3jO+C+N2t
nQCbpAmvD0L/4PJMpQlcelnI5xbEP2862gF1H9ElWwsGmqzfdEsAxMbZKeHTdmGrdZUqabPIK6ec
GCiHBFV8qh+83lzdiA6uOYO4AnO3my+os9wo/Kt7smajhJcFizzEcEWWQcniVf/D/SbfjHz8LDfU
bT/yrSU5qlY7ci48R4iR70rRjLhVHwGZBF/b2NYvi/PUb7mFgLOZHDC/F/maWpWIj1vcmBo7Ms/U
BUfz3hK5Sw4gfKMkG7zTAoHvttfK/w4SG87vvLYRX4nu9JLyEpcdq0DfjUW7NkaLePSCLYZ+hzgl
4naRWvykEQIjegxgoE1LJ73nJxjtc1JqXkC+qxFZyusV+St50MAO5x4IHEUefIurGWcyLpvm23T6
id8X0PLVg65jrNS6KT3HOqWiN4/vCP+WjO7npT0H7kJ8qTrJ79sjx667zb3egQjv2Y8AA1Wt13k5
1GflMdl5msB+4U/PQesv+5YCtyAEUF8DopUBIf7hwhW2R4mEopIxbRKmjO24CswuLdS02fbcS1Am
FDm+Q1Z90gogwIoGM00U+owNh67uLMK8DXvgNS0KxjpXfeC7w6UtqdyYgvMtSsbJDH4QDRJPXGQa
/SP8sm1CL3nK/mvjH2qxx8O7wL5p0X3OEoa9YZUSW2nzUJtV63kQLwkOLpVIu/6fPTufS7uAAey1
PXwQGy/b9k4U0MrSWOKaP5ubNvZ0K1j+hv+YsRi4jgSW0SRReR7WrwGrOyuATkYxkMcmbdqvCFFY
K49PUmZ7aTKmVy3Be8LgI3v7E76wq10jeBM7VHu+p5sAdwOav798xjYGNcR2EnWdonGCWUHVB21t
Ab7FoXaKgIdac0dUGG8quImetb1MEmGwa7DyeuMtuzMk/TREHpYuUVX/M0eMfBhuP8VvzG/P0USp
ExfIpIpoozK0BHlTtgrWB+dei+mvClX+T4CL6VNvQTyPTdQuyZPJnssNnYvFIWSRc+JUEeGab2HR
evQ4+IKOJQlmN59nsszUfwseEFwog8YJ7IwbjGYJL1bgUPjXP4pWodlKuO3AtNDXCnU1NjZWLCVE
/5khEFJNhQs0EdECthSJEIsgzwxhrknohfVpgvg5afmIoHjdwyl0FB6/5M84hacREsyGvLwrGI6N
P+AgL4Sqo//KZ410mmj5EZ7ykwcxwuWAOo5ud/W940scaYmtQshi6kh3jSw1j7yIUxf3SrkzUkfE
cHtZRvFT3FHOplsNBpN01fKmUeck6ZH/ieDJLCTlLB/101s/FgiZT6rXEd/jJ0K3RTpA7uQ7RnHk
JV3dwm/UKebBHpNEWc6e/1twqwrAv0gIiMhEbeEUIdz0FAYOxIFYYIxSPxNeyOBre0r4mDmuy4OG
HugU2zsnTdb/1edV+jcl3Ve6/ukvHeS84v7ldkoV+ie+B3gxw3lrIrNEizu3mk0Zc4h8+JKcpv9w
wrR3qmwi+uN5WAy5JueIGHM2baIx1e6K4mrXq74bV/cEMdbjRdL2BAbE3LEC3RYW/q68ajEBhdOd
1tOZI+qFY6pl2I6dXujaOBDciQqF/qRpd+vHrvITjxjbquEYcCJFhdfWbZVr+kM88nYmhOXaZEIE
XeUdsNfxEqCA8yw8wGSdrf/1CcujBYILypxGGz0dyNiRcj0Lakw8uT4r3oaxUkBYJ4djl5wxjUmm
hGSJH3fZz75Fi55qNeCDycXYU+y5J2dFXa13W8WFA3jpgWuFEOBt/YtLwOhe+3x943ZR0HYsE8aj
6kdBUYXId7kygjF+3N2KDeOYt0/NlRUOfA4RS5IpPgBWfkLTqMyYkOb3ybQOJ1ntbXuMHfjH1xFE
eu+PqJy/vUx1v0xVIE6+SjA2m+OjutRDw/C7600lkxx1Krmb49MvI2C9NPYZElw97SeeBfJ9lpER
3/J8OdUQgpHLucd2G3nKjss13VaboIXricXIJeNcMGPMJiTbeY/zgsT+GpGeAZ6UoOVRMZLgGbkW
qt6hv2lyaZ/Z4iC6T7oLCmeGIy2I8iPjb6LwatcWncDjjdxjGoFbcxstR6RQfhFT9YXbRQb7OuMu
sLl8i7dnfLDKP1Uvwt+DbAk1fzS+1mkswGGykh2wl69oZtUdi0O+7d1D3jXpDd8NUEW+FQ/A6ev1
AAxIpwUxWLxgXOcmjtxpJONOqgtps962XLYlrs99/5acBQJ2he5BlWsDS/ZV2LxkEYn8mN/Z/PGQ
OUt4u67Z84hzz9rGaWc9zUvEzoPOSWy9UhANc1vSlp36a0oPIyLt5lvdzAiPKkfFKZqpLbBSt519
LsarZ//Lg+2Rad09/sUA0k+FGVvJ5ASoLkib4tVxtomrzBHrezd+RKqzRHKhZ1t0hdJgtubVUwku
pMVqN6+/Fcuev4BH70w9O0lKup7Ry3SYr3o2cR6FApGdF6b34K945GxGrw2F+E9HgXYtVHW3wRwh
jqFE2fdKxIo7kBR3HFXMU8HrQ3SnPd4q6RLpK1V/oxADhVwhzOp+IVaxMpyvZA8ru49dwP4TLLnU
Uap1Pq6ovUPVcjndMjAVahX92RLS+SW0ey4E5hLDmhAatxoAEdmT6VnnHAGpmciIs8D5RmboRiSW
lTPeka3dvF+yOojFmB81yb+wret5+RPB3dAqU3YfwHX+ugE0yoi5HRhnEKQdUyeGutISQqtEXxl7
pmATfDqGTXj6Aa9FBXpUoqoKPKHChUrE+BP2sJWj2rMiazGsMdh9WVdbNRxCuVILTld18TFjTulg
0mQQT/vPQDyB505iah0a0V8wkgDiK+kGDxggYrFo0CSd/ncmfJMG4nWq9Xnua4RB6oPDAUsbh3gd
oje/74jfQcgcPG74U/wUfeQiWzv5uDycKlcVczk//Wsmv2TndpRriUeQQHeEPAVRHeZ9JA8/AW8W
cvNokofxnz3dQ4ZDKzetsX1M56MZEe6HSojm1OzjJjiLFv3eJg2uYhazJWpHNchaXcg6frQAj/3/
NFnAh05iKZRahWUod94cjoZGkmcqrLZp50tdvl0wk9EE3B1PxdIuI2XFyxaXuvknv0XJJYvLt5tv
LFBX9n/xRXda5orW/XNc/jON8WdCENgm5A0a7YRk2ltYtFBTc1a+zxScH6/ulvi6cWG3SCtNafUp
LCPkNJGeNjtFuD+DBWVEdDgVmIcb9Be+zDBUPTnAIPO8nXnrrWDH04ke+W2A/c98lAOrLg67mw6q
13FiF8pIyU0MQU2K1vMUmYnBItmRigMWEAhJDS+DqZOVThmtnrsVysy1WVwUvQDlPTElmKsHKlcO
WyQd0UG/rA02mjIMoYA11MYb7F6YEodTvkIcO7HtrPojibfyD9VEri14uax5memYqEZevzu2pHC8
DNi9trNWCV0uNlaF+N6tNNuo7X16ypc+UXTPy/+MmQQtW737A9lMb4FijHdI2mbquPuR8EW1Vgq+
JXPxu5tMzzjJFtc2JMZSjA85nCyVvgWbTZTnI61HYIjTNf0uLnqv+tJZS1gqbv724sSudO1ASccl
63UuQcPTjhrmgRifq09tDJi+otTxO48N4AC+05xJNtZIYXbqTpPQ1tTpHg8J8G5nE49AXEs0ZlK+
EZPBQB9wF3zUDxENYUltN1gqWhGLLEoDDMkBnBTE39RoGyt66t2vogRn3BX1YJTElLzdMFDMifTf
QeAtxoWEYeIgwulS1FDweloyK6nS05jE2VSrOk17LMhHY+0jF1228eDu5XEB0q8V9bYDDy3LECxX
mO8+tobhxAHsq30Yb0M87tMiWCsNKcyg8wOSlf8qN9uztix4FX0yBt261vFB9/kqAo4blPzc1e18
KSUCeGLx3ptEcJ6PQjhGrw66JeVVhfU6fE1JxG+4zFfnK3nuV7T8oSmjdFrqsgdnOo2qN6TVqnQl
XDie/YHR3N4OxJvBpoHfHS1jqsxLEGkmVIn9b1M3pzXZtSfT7HRf1906NATloGHRpm1nOLhSrDB2
STbvZyvuxURmZSD2N90BsokeQjYizZKIHL4jaDwRsKbL551qLjnfMbgu7qIYncQd0x9BVuX9i2AS
sOVP0ItIFEZchuMIo6q7QgwRzPI1N36KqxGAMdPZz9B5suOPCmpMFggmLCXxih2MbWKvoHeeAIlU
Zr1USG9vpsJT/rmOgxx5I7SkKZg2s4snkfwhYcjOFEBSYS1R8MfQmeLrrELwe9VypiyTHqfKi9nA
etycM+7neQXKJuyPkZgyogum/FNqKyaNCqKPrQQMuEA9d/Mx1Ui5U7ZWbAJVXmVaC8M6H00gy50E
tvlOlW2VBJeHVXAhL+4sn/1fJjOSBnRUqo228TOmivdDyjhn6+bklZNUCD/qNGYm1HZPN7SEK3qg
uQuKhJrHt8A4B+26pUKI4c1JxIeB3f80EOfQptNSowojBAl2NeHuHFFmTTY5pBm2Hm6YVv2rc5EH
MqnB4F4S6oCPNLu2e0tWnVdq8CNbVLNjrO2gKnICKfB7J+ua1p9CShtAEsa6So84xwUpDP8/7z2b
L28GsSPOQPCGM48EThSBdusqyqZVVBpTY754aRT732prTHAC6FbpRITTZzKMCJw004YmCfOp0aKr
tOKaQsrTk6s0OqopQqEdPIrrMMVOLrjn82VZ4NhfnAs5R19+Em8KSbLdJGriZTpB36Mjz5umNpwk
QPKF9YUPxKnfmyBDegsjV3K305nXxEp4Lx6I4RvoWOJhbJ5fefc2BqlkbqNlApIm+kvvRuEUJ71B
vufrpBGdGcFgCE54LRmHYmfAVOfoo6K4P2XalSuZvOsrffXFigYjbJHwDi5aUc1Ps5MJAkqieExu
fpr9pV7beWM570MzOh732lEMnAMKsFMGWY8vSyKjwJ+WusOQYGwYe1/XD7Y9D+dIq+UwQNzrvNou
0GkbnqmBX6FQQAiHldkCJ+5GkdJcmun/2R/bT3Y4w6tdA8jWb+z9cX+U5408dLyLxiiOgEqRA92H
D9lJye/E1WAtxbGSJgW9JDwP6O7vRjpf7D06zxmb3g2tRHuDyQ8Y+26cPXPla8ABJktguIOOzdgx
i6YE2jij1XchB7mIR1xcrOWunhkITJO0Wjrt7lO7E7B3s7WTmMlVCOfsOakL850BGhhC+b4l/1Iu
mSdz18ApKF92KMQHS55FR2ciYGfE/0NfH83ROdytPjtiU9T8eY9HoBMEYbEtdeiCIA85GhIguJ7v
ujTOyBr8JUaecHd/gCT7zGHxLmic6OnjkdjeYiMf3rNSJxqtr/AxE0DrCZe+Zjx00nocb1aLPVb0
ATteTFrR20cMeEVSYJtM+1VPh/fws8Shl0tpX1HLW/pQiNonBkxWx/UQ9lfdmTLIYnnw8YhidnT4
MGr3kEtayMuhalN9DKoI+d+O3ycKQeVx9gX26aLPMWbrrYH83rQENfJYnsfBtP+zOak/UFoa1Sfm
/t2fCyUj+9kbP0JlnL0KHcP9F7juJ7be2ShJavldc+tWQG2dN9Cm5lLNl0aDy4vn96PXoqzV0uYk
EgB5LKnqAUoOv3+Vv66ppv/9XNbaNOSOgXKLBQfOTHvZCP5OKNoxtx10ehQcje1T7YsBj0DTG7la
AC39IP/GIGPFmKUueRQhwF42U1/4BVjh4Wvy0ZZlvHFbXKKYMrmWa55uSIrfiwqSIzymRXUTFNS7
5/fMIHTg2Qg37Ml8bkNFO6xqY8LMo2jh22ggvWaTTjKc1EoOPatMG7d58vuRXSeJu49V0q7SE2/O
YkDevaFxNogfQiBo8l2KR9PmKsKxPI1L94iOYujDLl0V/0+KIqn5pwz/JW4IQPl0JoWIF/hf/9xF
P1o88irtLhO3gQZB95a7AslRDnYaAldq0JCtGmuuBxvwF3SDswpcHNdcJ3LCsMF8w1QekRQJ0WxI
b2gRB4Rh2fjmalNh0a1DRkZE7uJW7D3Srkalw96KMsEsg3guVDiwCt1gPxuYWAgJvnbsZ1465iOi
UtcivBoEGUn8mzVVPKMVluaBRcrsCnKHX7rfui7FcVcns6VUrWAXw7YR1lL6VI9eqOx62ucia/wv
mLcetC2fVmxRjb+LhL+WGcTLHjgSpQUyNcQd5ikZeCPLm8PNMGGOyVoqXEv+5pKnnZnOBrP/zDN1
fN3KziMzwjsaqGd0Q5TReHPEmZ4APDewuWKv0LNY/dPv6UyHsX7N8ZWwtAy4aMf+ykzKrSj52/Uh
Ur/C8PTjGMQ4MdMQSB/51P6KHjdcwnBteiv8ZO2H32Z0rujzVhp+i2Rxq89yijZhTDBs6MYTBJ0K
z/2sWKzWHNUjVpJfCMXAIyKpSGNKPbzzwYJQ2nlHj1TxhqHmHy6PVPgVmtTM77jr5PwqYrvQ6b0j
lyBSTMCimOaeQ6G6eYhBzxemzG/mGVfHzWSZK5Xz6AL9tRPiJ9Viw6cWQXLapVFw8vgjow9PN4Bh
9J9Ingk/kaqaPWxXCE9ADrx+IYj7IwxYw9y+pucuVSQ0uPnxX5ZNa4L1GG5otOHWHik3wF6SsLXE
zRDzRcwKz9qgQhiR0i5l+XNHJRSpz2NfXEj2EHNqRYLauyVkIvRB0sKZH6xFYLaKUH9MYTsedZCh
PT09Yl/plFlUKYnuVfLTRv6LHv6jthke9N03bwrE42j6FtqKZpQaZX4Yt5173easUSJnj4ys0lAj
lil9A/vKOXkioOeFuTS3JgwyislwvOOF9MYmWJQdrTmhPQ0HkIcVt03iQiXCK07aT/HHMfZR9gP1
mWX17UiWwJc7K6GaZXCp3Mmm54WXLjuIRWGQCOS7OviYqz5FNy5lFbTz+2drCMBQPS2CshQnQJlF
rz8UpvWKYOEfZ2dT8kM/eH0DyFDjKdo2FnQzlJh4mRzs+47lm+b774DNLQ7B/xvhLVuPRROkqK3F
9LA5fGh2mPzuO2PLbe8RhggDeigvATMjDxAKATOb6RA/LDLlXTdGpYLjdieVCf9UjZIosvJmZ8uB
YSRHb6Xd5GG3Pk012wtuD83kXWe3D8OW7ZzMxuRQgjHlAR4rQb8fvO/cSYcT2CLwYjMKcStHGQfB
w71xRYCiABk3GQ3POlV6PyYgvRVGhmaRp7T7Q5WN0JCoCSVE4zz5mrVkwlvjme1pK9pRTPMGk8Kp
gh6UZfUepZ1M2R6+eAMJG9f/BRtoC+Yb8O/4OLmLBFrrvaFcFFuHCwKVq5Gr4TsDFr0ZHFMZSOTO
PX9T/PNmC/ENj0AIntjBoDwARc1gyhlYd1s/qDh3tFx29w21sZdqEj1ZIPMTna5g72HeO5YWYpyE
srsCnKGiAhGAYHHDb4SpC8i5FYUCtoVbsSQlAOQ4iBZm2OxzJBN2FJsCJD5rK/0mYlPRtxhigqmF
+6pFvkGkmzD09WCdwUMBl8Dm+fznNsZE3cGUDg5p1YL98Zq0Ja2F25zsYDK7/U6ZEdp3sOi0kNW8
hUbh7zX+SIxuxo1dc9KcdSLqPGMqeAIQRxX4h6ZQcGewL6Rn3HG0OR7nXF4xojf6xvn8q8IOr/Lt
k5cWZ5gLLn1LEWU12CIbIVbdcW5Jv2BVr9tRB5mzhxm21B3h2BiemEWsI9Gher4M2LoqOqUM/rs8
npkUVQveFhp0IPCy0jKVcvk4ES8KIXVmBanucBsZjfZ5zRUbN6f6AVhhPnPRPmh6ve9WfLgkgDCH
XNBp4WJj89HCO9Y+lzofmYNjpmp256wOiesUz5OZ4BkFd72Wt+ZZzhJpEaOZtE1IQOa+MCzGacwC
oy8RvCGmDHZw+I+KUup7VjyZ5IgrouMAtdXjwGVZ7LPU2x927XJZ4ooKqD73vn84u2fhdtK7ZGd+
RjUGmCKVNYzdJefg1lxI3Y+Xb4FScBs2Oab5r7p5/Lh1RKPeHEYNQKHmunDefXIXZCN3bD1Q6rhQ
xRlUH2DWh5sG4IaYHovWrkegHLBUBaMyIKRDs0YBTKsdZVx0nGd7iOqU/PBqyU6qaSxnPEhkyvPA
R5Z7J+xkXPvZTWRm5DYcOGrwi5TtmG28BLElRQ3jENvkC6swDE8M9vkqkqm3UPDy+qmZHe1ypYBm
O9RsjCBmfxHTI3L47cTC0fihxEp37/idyJmGkkI3LWV6sKSI1+TrVU4NAJH99URfdDzZ9U1Ci68L
CZh+8vIVnmxxxJ47GbctHMMvVYqLC+60+q6qkbG2FyuTMgIQIwPkC0IdqKlWJi5TTsz6hTpmJ51B
ZZY7DZzEYdm5qRFTT5whBFlVVOWNfpR/r1YBdrV4OQfXPYVAqkWfxzaOlhpDUTdM0BaTgLNghflX
4ttTp6Nl9pr4+bB9kPMu67p4W8ht65tnQy+KDQyItdR/TpzaIhJMjghLAxxPGqZj3Z1bawPm89sR
jUc65jPjUlDIxClmUR0AsQHCQsCC/ln26bsMTFE6w8LZKZ6cLqmyTW3NZ3+apV/4oF35WyKVmePt
vO2vpY+oePlriaUWssGz9/1hha0lsG9uJVu31i4ZdaV47sCKc7Umo+dBXdNM9GHap3wcwOHB0gHi
pC6Qfb32X5opRENPVXexUTNGXjSnyoc692eCBy54o5Pr/Ax8ym6pyrNWwT7p40g6NBaxQCnIbmU5
dqGanURshfwy7bXkKmt85PcqPRmCxZhupx2RyQOWpwFQr2e/YvE37v3l2B8mWigdmnnij2B6GHJj
oo0w3HEprznfQl5zjnVqrne+34cApS7jvSNKPmInO5kdlcZmsCSpcoLIRodqqg1PFTLOqm8mMrVq
Ik8x1QnRsvaOhPCk79PW2Jt9pGOMaT+3LdrPGmHYP34YOKIWWdhFarI3LoLYNCWq7K4UjDCqyaOQ
jB3dTbXb/uPAfeU1Tz4DJqmP7ywuWkp8nxd953L0mPbX78AtLfPOV1mJJRD06iejtNiiXidegl54
/2xEWvL6AfT99fAWsUbCPIqqGiJ/YV6KaacL5uoduD1x00KO6bgFaXl4w+FDPYOE1Vu66xmvu8WI
1qFeZIySiM5vUqFVw5hli8x93ZYvSCGX57dojXKUXN3TyH7Tu90GfSYrJeRTIDxI53rZfbAQYGk5
Kf262OvUl2cdr6aYeSxriMJDLkM3GKXryJ/nszNatr+yxkye2OTyHY7p5k+EDxvx1mQFssRLoaE0
f4k6XVVHZNEDj6stahnh84jHCZvTdFyhnQYwIUoS9rC0IY+Kf/ihcxMYXwHCUaPbhVjVDduuux3C
R1TqdBYO9b4bPTSaLJjdjJ7SfXK7WSKMmYC+8vDztZGHmJ13STy301PzYfe/Ib6P66YLys2qlT14
bducARfSkXPA+1hstW/v7Kh1lKv7qBiGHoOPOXabSR/MbW4Ens8kOP5zf6aETpHcOuGmvCa2wNlc
lrPHgFpPWQ4R/+RmEMM1NTILl2GM/qZRnQNktGgU42vwg9YLUFQ0wGTz+Pu8XH3Zmq9AkujfewLf
8GKHGC4jy456WV1DL2hQNNOY+WnWxom084wEhbqdckQC3nwZNMYpx4ZdGKfT3JonxnaBuZqwnJ3e
o6TaDq/uajpVeyni7lOEXdwlOIj2uGNyQFHvhnpSYuintQa0a9oso+C0mfn+2uQFbEZTkCOUz2Wt
p4OYIS88Orn70S2DppEkX6rNP4J9RIQesxChRtr/ebIlLBTD9YSYsmGdqZmJiVp41XKBImYW9Bm0
lOnlpD9b+Urw+g/9oMCaXaLS7TEEhoWOHJKnqfiDPtu9nPPXRX/PCUzxJIRgllSivrS/P0+zF5ZJ
e+OHAsSdyB1G/UWziRlaPQlTXdiMIktgX2jVykMo0BQUjEgP06N82HE1fBMc9dtVtJUTIKDanmca
jQDVD5wWDSFx8Ck4AeQlBFcZQbmaqV4YyCwt6CRBXhHOekD0l5KvP+4N3Tltj5Xts1sRquyoBj3F
svTUjRrOwwbMnMg6JxSUj1ysPUKsGLO6Bg7BqgexBmSAwetLesCCoqy+BSLOKr55SQMoNd8ZXYCT
8WmLeLyqvbKrFMV2xqK8AS9m1RKsjmq+9Vjx3LE3SKI6w2WvX1bBNy08tab8r3+gwfYsvCkbZm5D
g9fIrqAXWviEUNguCFyzdL/uFI2FfCJlXf3UpTSoXRzfqQbDS4TC2GYPWT6ayRlSoLLXWdoa5hSn
LmWa0vHh13d/de9Jz/mJ8SSSQ1F5yIhVMLyHKxIpI+jtPYVSWq3FjTeJceZ8cG4/6DVK+ZWjCoTo
fgi3ZTMX96P6o+kT5TYwwcaQQ8v6Lknh8bhANE+tmWa1wvdWd5j5+vgB29uCS7tvgIkZEXns/qZV
MwbRN5ytzokSPkiUhYcfQxWbgMoVNYG/LZZgCk3amXmM0xpKdNT4E8e/ngUZcP5LM0sTey/1Jd2Y
X8C7t6ngOK2iYfK0U1lbPvDryPq26ZXbq3tniJI3r3+3im+lob9muuIgST2sdxk/9Is9f8wGZiVT
VTTER0r27A20Mp4itCRr4HmKvy2oMuO0/dM0DyILEJLdYumwHqJLs3pzCbJK9sCIZtfbM7iQ9l1u
OdbxOmtIX3EvkIoL1+metT3E7cFs80FamFh1+ImDRwNKoljbML9lfhaOKfH4SYh+T0XAji0xNawX
ERPZPPQ8fDVHFNFXhEtypV5fTRXuTO9FgWcqshzmHW/g/NFGdczurv/noq6GuooHvR4Hukr1py1B
Iri5nEC08UEGbjjIl9GE0w2PdYwGP5B+Wzetl3ejJNiyMmjNWoeNgALrcYIIp5vuzQBFkX2g5YQp
qXpZCRsRUUW2/WBmP3QatvrkrPUxq9d3bzvBVqMofBmhUmVnaBOusrQ4cmjI4n6T+n+L6dfqDEqc
MIQxOfJEZ7q4VRbquBbUcp25C8C1TA9ZUJPxCt7R+xMPn+kcY1clMBc0Dk8rTCW9lBuuQ40y2O0a
GhAUxFVK59pO0sRyY6k5mjVgzwVpu/onRZyPSQShcttrj0s3jMgZthU5xw/4ZjG9rhbmI11gRwZt
DPJHEnNsIjg3ayGHz3KggXbte6XZT9sLIwyIGhSLaalBSeSkQmIUphhE+SVKh2SRMZByGDvTiqJe
AQP0YXt7n1ke0fBop5Q8Kz9gczJDXrhJV69t5m44RQOOcDsYLlmU7kubLavu6SyA7M2osU8MEXqU
Wj1Z/aBHC7cqiRwEKys0/FRmO0UQ7Ma37jLlbFUteJl15w8W3YME3cve/gOYq37njPPLztVcINrC
SuLEsEdfEq0Jxy1r0RPxco2xrpuKRIueW6bFiAEAmXoCbW7JM4yPG02utzP/X1bUokntIHoFBpbB
OkfrCOPf2m5tJHEF02+uFRUwTzuxA5cRQks1BcIylhunLT2X7rSOOBnOHYPYLgC2UlH0drRY0iBY
eeJC7Z5aBQ5FWtKSMoBRGaHSriMOOLr6rcqsn5phgvlYRFDLenT2TCafvXS4cnYkJhpBGPe5L4oC
fPI0EqYv11rKBM04fCuWJx30sKj4N5qExHZwZuCdyLxXp94Wee61ieNQ8lwNy4NfA3WFKvLcczQO
XnGNzqb18jKjSs2vKQnASMhoTUxeGgdjN0EpCNTQ8xXIfjIUFPrdN8HA3hpNgIfT+WlYnDSCSFjR
rIZELQR4XE+fW8JLEAia0V/OCM62AHMWqYpPEFFsujoFWGblvZwCIe3JAckt/yVl0ytIJiiGbqGg
s8z7DHhLnpi/tbV6GckNziZhnPrtDlJfuONhTxl5FSGKPLDM/0pRuIVVU+GmwPHH3hx/LdrUStK3
lzJXL5pQbjIWJ8kOMfjre7A1XZY4JQOJjQMzbhd28aHX5D1dYhW/8KlqjR5k/8YqN/KIXI+r5PoJ
VzE4olJDdQZcURyBvUqp+WAG8/JFGRuhTk0cgIPBJceA/U1c22kBv7fCU7X6ye7T0dD2f2JTy69q
mihvPQkDO12nNHUyiPFTPsjW9gb03kixvu1HhxYsQq/QGe6cnH+felm32twm7CmOr7Xc9rev/0go
M68MfWzzPd2PSU82reWmyq3r03WRwiwoY8SkQeum2o4lbw22zchqubgEMT/fc9/gxU7c57fIRHaS
JU9HTAXFbrj1mo7ODMH3WkCyFZDJiPYIG5QE1IB58KG3oegrOMYT+W9pPSepJkbWZHj7XsuuYGaR
ToQQREWGxX1Pm9IRlrlCv1oKKa3Xkczo74+GXCXrinEcgZ1XlVDgMx8g1hThh/EUnt3LUGZPm6oo
c+iDwIG4vmrQl5zEwM2EoY/1oH2t/o/Knf1ECiKK/II9biuM/Tb1nJPdVkbfs6OaleyCUYep/IKv
UlX/Td/njc2FuLO5meNL07eMV95bp+h8oQG3ZyKR1fa2dqOxjXgphnrDciZkVZyP2nqFTzXUz3x1
+VvR+coQZS1UfqOVEPaA3dmtw+iV4qOdZjTjKjdsQb+f8SdAS1Iao9N2Sq0hJZUrU0K8BSR5jCRr
puw6IY9Uz6VV+TrQYLGQ0nYVXgwWAc6pbA6LQg4vtqBngb2OMjkCJ5XPtisaGluLKjwV22s29uKA
diWIjyNH7Xv708i2h0CzDZtnKk6lhOU0E8NcL1TUtH/c3QKQ+66Yp6HLQM2I+/AtT/+zpI+7/ji7
OnlKvhQ7V2FXAaTjJ5l9oMk4c9hjo699mA/L4+IOfBqylSHmR3LVXaRjcE33bIJ4EONPflPXnL2h
Ygop/p5/AwqvAZHhQT1pcuzEpN5fMUIi7eVjf1PTbNW9TDmCsD5uezsDvci4ang8cPcFddO8L3rl
0ehnHWkNhbICiKPeYHqd6WrZ/DkAWifnzoI6J/36k+Z/5vEqgbB4aeko04+liTnMC9Qb1DU1zzQl
83T3e09S7Wi3F5+XsKT4Vrwz4lYs6GSXtzjNYx7pAP5xm0RDOZAJCfl2Ju0JSxAjNnFQIEyxakQE
0CyhVD9P7YRxxz7YnNz1zz5+qChfuKhOY0VC+unV5Biy8yaiBHsxj3XPdIFA+hMDwkuBUvLKurXu
/GLYoaXwyXFB8oRWUdOegjEUP36jnqZaCQmlFG9HM7RKO0a0S35ds5P07b0iSJSeKIYqNv9ZcrUG
sN5gtOriP2/J3ye0r2oxrr30YsYk+f2an7Jfkn9o3Vcf2P23xq7/4IydpSrR9G5iVRxXnhaQUhtm
Kq/ZWXK/ZMLbIiA/Nc7SKo0AH7rBynmppdjedkTVGoBfq0wZmJA+5HfyLZMHz19R5ShvedGOMTb/
E3fUsX4kyFn0KEV8eRcK/2BWEPA9T6mzbVi/vDpLglZPHzzLHdurzSBjL6ypYNew/Z+bLHSfzaIi
DrFDVdVBdhx1OjN/UIhPRHGzov39ALylf6IbVCEvKRz8amr01X2utLTcmFs56Gq1nBeI3ZOqFtXG
iylRD7toGS8BHwQIkxWmWvfyDocFx70WshDLRqC4PZZgo8JeeAHWTWHzXU2EwD89QBgG8ApS/BDl
I21mEIcnz6SOi6XWt7jMxpG+CjS0ttgLHcDqxe4g7X8ciWPv7l4lzJ/m8y/Es/h/LmyA2gfEs5Kv
4qVEiX9Bp/LG8acFaZL234jxNuIv8cmOme1M2tHSEKb2FaX/Yq3ulrIzL/aPVdniN4oUOMaek6Q6
w8oVU+iq8ZJyO+44onxW5u+jWBVFqauALQfyrORMyUsns0J77OHvjw514Y6E9waJzFrK5zuCFJzo
HsdSNaD44PM1VCBOn8rtLRIU5TVA1eq2Gdgv2U40YBYxHoJeq3LzLov6y6bd0VNINtqRWBKlS/EJ
q++87yMk4hqPsAv+V20wHiTDAVR1ATfXbJ1yo5ckD3yN1TA8WAh8VYjuVBYev3BIm+xaBk/fttLE
Nm0Utw0OR6PX4jD6FQcPKmUpTT/zjxpph0WCmKZcYvNtKi+JogNzpjpJjzRU/ek2BIPHLSuZzL0R
yK+0Bu9J+1x+ZPY7SqDzguZ2fIGGjxMf8bb973rC6E0QXdVIUBjYnNzneGTKtvQk9z4ne1OiuJ1p
P8GMwMjOpApelcPikygODQDCD+eaf9ZJJvrm7mlkYO7r0RonqsSJhfwXe6E2BhaU/ppgwB3DC6Ar
rf2ifEimhwFJMAtupBjq64RIPKUvVqd0oW3R96dFkTSsgjAmwAb6aSu3hi+fuGRIZHJxrz9MvjzE
0ldGtO2gufGy0B2IN6Tkn2zAmLf/HdZl5jkhiHBlHWToVmHBJdFA5afjbljfucmrUgucfATEeysH
nvwZA3E/ixT4JYd0y8TO4ybvm264x0hyoOCLBpkhAn6dneFZsZPpP6mmurtu6gpGVx0jp6q4lnsZ
DPiBscQPrCC2rAnJrgQq/kJa9YPMdYg/W3ETy+IdWNdHve8X3KJ+jn8RIZWQY3lNHjGY8GFfYmZM
XB58s30RrpAaLBeZH1iWs1HYaIR243AaLT7zZKyjMUKCK+b+HdKqIXHSWdVstIYwKHOK16USFa/F
XX2wr0cgRDlk8A8i45Vhz/ZkG/XxbHyWJ6F2AqePGxifB+OgAoQNHm0QTOf2A9xRbmn0pt8LJf8e
6nDomXycez9giDrgT9Bi3czBH7k9DPwsGOf1kRtbzkPj8Eidq/9NWn1jz2qNopzut6R/gJJR52NN
UZ9Y34bI4JVaqkbJX5TLk5Eeyjl3g41Exi0ex/Rugisgg3MHjQrwqIrC4QJuRFFqeM/hj0Y3Dsov
vtGiA07XLE6fxfTrNC/x0Jsnpik7jKTOv57qkt0kkdcShUyIjZV7O2eKxgX61AZgbApfsl1N/3JY
T1/Dq7wGG9z2HanmALhlxilzrdrf4lsReQ/9KUHbvyjKfAZadQ73Z7smPWKBmp+gorCJ1KBPzL3n
/3u9oqz//bn2YgiRJuqJz7lrytEMOm1BRG/NpkiqxzPqwBUA2H8GHp7Rz/8M3YDnv2wves7VfI2t
SEhsMnf70megKiljGlcx8MPTIZWiJFnZilISmcqMg9I9sNFMNeB3V6teCZx/VJ26+03W500T2EnO
Odwg+t4CY7y5eG/Wt7h6HdCovVtHDyGUThDf3KOMp3FGPxNfPOVgvVikEWgHy9t6GzuVr9G1SZIE
AAjqeFvTXRvjgJyiUQ/iBVb/BPR3I4DTxkv3rbnmToTW1NzbN8HA7EQseMpcIGH3vFJ+KmGXISsr
OeIMUz14EL5GIjq4S+049sXrE7zL0XsiYGNtbq/SIhTyECMOD4tpPkH3K79p8pi+sMPiNzn37QMt
tfGJIOioXpJAzd5z5cz9kHieIJ1IbOqmDBZ6AKf7zAverhVaZZjWonGhRNjy+xY0nAU9QnRilIm0
+TaCMUna3ewT2dxbAmMlKvr55AIm1mOhvGnYkGRVW8ePguCvu75wMkAZAlsajOzbS0F7vkAnLjVB
kt8kNizdoD3jtF2lfaCclNrFNOS2pa/ZB1oc2w7PCYB8auc1RXzRxSB1VSl26epafea0dkZY0eaO
VwVtDA1+s6cJWHeJytjItQit0seWI6iPZrSqdhwY76FZEBWmLruDCWyChKlRbFAzV1R3mjttE16o
ks4JhvShUeIxBQ/gXgdwRFCY4nMtCzaezuPjY+RKI4+ab9bnYe41WLtbGpRISfd6/YAB3wjjYHm6
GcRE88nf/nl9o7dUGJE180EulRegI5CIpzrzTnwB1rH9vk8t23tg+Jo8+pmP9ph0q12pXEk/tUao
q6MNfMRTZBTUf/dc6pJ7UGucIBtnfcwpdeo9Erojo9Dbmzb+GEWJMcKBozap+HxeQQtg2fiACvFm
cyWybG/jVPRXlEDdsbfZVKRRIuf5cit5IOLAaTrWKobJ8YBhiMPTDOyVSyrqOfNUa3VPdPdCKy8v
AW+Nh2+mjcV4lo+0fd0S2go/pSuanR9KwdOnLREM/or6qZLeoi+zzoEUpKXjcFClJQX/m7ZJHrie
bve8mc32gnQLfTAk2hPJbjeyfBp6d0Kf9AgHYXEosnRuJiVd+RHNV0ZwR50wGucsd1HR+8CF4lVs
R/o1EvJGW9Uum0p7V+RO7Zmgh84rJBPADDenRirWp7bR569rARhT065mVDsJB98oO9xTXcsaLqEC
0V0rbY01oh9cZUORxtajN6ZG2gCImsg5cfPFUPyblzedMZCGXWrRqTOQQoRKgEa6xhIk3LKkZbzY
9E3UYSC4x6px7mjBfVcaCxRqVKYXU1UVtYGVT3m8SAtDyU4Ot+C5GR7Xy0tg8RZ4L4LgC4rz7G1A
1NpoQu76mM8UFJy7Lt1Z4sL1M1zKtRXoYSRg4MYBNGzhppH0IYst/XqdwwvLrhHsIlbwOmirZYM5
Y4YDBjKle8FXHLcpfun+YRRQIbv+waxko4K0V5uy5gdecpdbTaSIwRyIOz8VcJJ0VbH7wNRuv+h3
HhBtyuNbaMliZ4g/+Q9+xQfVXPwgkHeYA/61KiwjTDN4HiRCb7vZC6j6DsoMmpebvbxNTy8W7ZAZ
FiwKaIWfOtkwAx4GWmSkZTEv04/+IepCyG5LzMVZspke7ftgDws9wzhClC1kIDIMICWGYA+FYPuG
ijRtsEnXWW6pc5rvfsY1by7HKCF1MuzaR9NzP73XL4QfM+xzjES7haYhVKmGPU09RXV8TZ9s/uL1
pIFWNJFL0SgomzGkXEjJp+sQOkIK1J3IbWMDm1USDiPUvRAbcYlEQfkHzEGkQ3Bht94nymPJA9VZ
IyBbG3sLTNgms7DuEw7dlg+ZymLjCxIDz/S5T5dk6xKjHVRe22peOwCZdlIGG1WMcmmyGxOEX4Yz
i7oGXLPBVfyQiBDtfQDZ5GRum3OuHXkowFdpqR4Y22SRZfXhka4F22W7MwhReh+DmJiHQsYEKu+G
IC4sOAhPUMLt2obuQdjHKAH6pAd79hrTiLzy8tY8wxGl7swu4mAmc1LQu7JGjm93bzI/iKNHdUcX
xQYTewYFedjsiiW/Naba5Uh9rhpbLhyx97djIHb3/D/uKOQKEXAvBoiy5rQbK8NNbqvj36akj8Z6
mQ9Y6aIaCZwFdD8kjknoO5EfqUpa0ci9aL9JBUUsWE4h2iaBOXO7tfYWaE1twTKJ1I5PnEldEgEf
Yjxw86CIEEjQ2o6mtxgkSy9RM4bySS4KF9XHJF9Qu20B6lkItOp9YydyTvOP3IhPYVVRTOQ1ZqRU
XbloaWk1n1krpRkI0M27Ccg/2lKNZlJOdyfN5faipCaMvFBXPzAKiFryb1ywzOnq6VYCNXW+1Ofb
z59bgr+wCJusibdaqX7CyYTGTfs+v4h56Y/t03MLrrTZ2D65oZIqidERrgErlmyEtuba7vD1dFmK
X08gxR+3KZpakFoD0Bp9mMnVwQl/s/+jyjAknQxh6LgUHv2oOBIeWikCyu7xr6F5dl471vVWfYRA
4pXJoVo99x5bqXuthq7yisR3HGl8ErFeFTRFDHvV3Y7ZJi/VyaW80mA525QtCqHvUZ47j2QpRE/7
GrnXj3o6eOCkWGPneUnE7IspBvzWOvp/EXKi0c4obl0T5pJqkAyB3pZizwZ8Ox0ZVuTWnvg1OvGJ
9brzGyGfeEZs0Pg1+S4WfI+VUoVVfVQpu8UOvjDZ7/Lix2b2zUZBzBvuTDHMZzkCN7BWBMubav7l
j19ATjoh3GdI4M6KaR28vDANDW9I8pMVNmVTYS3d53XaxqWcw4+bEvtH4Li0xDRm95QhfMa6X7U/
RhXvi2uuFu/1b5rKUgOJe6RWhkLXdbDo3Gf6itK0c18J8HmN0rKLId/Zb+MdXnU+7oCb9yGHyMKt
ao07ULw2qB8m5wkPhb+JLH1XCWXx6Z5HmRvDGf90v48vcRtrBSnOfSvp8qRwc2xmE+ic8zqo+bYm
bAiabj8OJhGCdFYKGzmHwv1l04/7kViAMwAssl4X/5piSiLgA+p2KTYzonnoXQ1P+NCjj+LgYQJm
7iFwi73PC1lohn8AYAz/yzBuJW40ztkI8L9xI/GCburU9ZXBTl6K4NtXE7FQ28ZZkM+ywlx7EVwO
BwgrZchDmXnrkPNXi7HxLaYE/QpZC4Llr1YK4gSvNQgtUEC2gB9sMGQBpstjG5jYdxNhYkmpXsvn
N8ETyMlcp2e+PrGY2+PgX4SohmNDtrVB7J903T4fxreASi111vK2mPcjpK7WRtT1WMat5E3QRcAs
g2sGT4BKBhouqlU+0RwQ1ZG79b3LxjxnoMnY58aVGPDs8632YTCe1kakxv+FLVGtd+ly1VJ5Si79
Un3bj5MKSl6tO8P0cIslZvIb7LR8ToJntdxhGOuC1ddtrOW4NsyvIFU6eHBpJZDiE+m6jw4UIjV6
v23Diyn6e7S3JAY9B895Ggry52rT+/oTof5EjPgxyo5gbUUf21CC/3Xoo29FyTYqgqd2az17fjL9
LnhWWWYcBNR0PYo2tnzOZo7FCKIi8wCowRF3VjaRrtFQhjr0IY5+Cy6N4XXesBbAiFdXvXKEm51C
dotI0LzPghpcRzUM3z2l1rXdDnU4nPnyQQQKg54it/Z40D36tcZ71Ip4KDehUgEkb+/bRnSCzDIA
RyaioE1rUzSZhASavQoYex5iZDvOswGMvpRAnXmuczgpRF6EwCYZW/ZyEFrHGNEFSpUgdUOLlyaY
crhFAQ173kjQAtFiyDM1xoYMLA6fiBKDd6gjsbtczDgy4tbu0aIEI2fNrxtZv5nbe5ov53Y2u+D6
TfOAqlTEOK/uen3zC3iM7XzPnhyZW6pfrCSKKNJRaWasFDux6T2vYyIpYio2LmbgWlQKlS9YHsGg
N/97qk1089ncE9oqeDw/kTSaYm6NxwSk7U4apgktL6EQlh/1zbgLEHnu23BSSlParyZ55RnV87La
xRYia5lBoPKrwEAkMf98gM4i4rTCMr0eE0mcFGcq+SpfApT0UR/wsbdPkjYw0jZu1yklUOF8RqAu
IofwUlEKQ+Fvsntptb7KwGj7zLtFPlG7CY9D6Mj1BMIg0eNUdp9YUngoBgvAgt27svCfWdJlh44S
kaZ2Rh1Z3W6dPC5PZDlNSTJ9l/PVi4ZUJNEAaDT3pevgcTyB/JPcrHt9MuzF1i62+9fhFWA829rF
UbnfoFSQCfnkrTTtpp5Zwckgsbf0E22fpc42ICBMVXCDLeh0rjFP6FOCzv229ovIvsioe9HlcmNr
z8DXchVR7AS08EgbmgKrkfGZbtGQGMATtGDmSpIzRpb8ODgjs0qgLnkXuQJFdfafvbdmHATF0X1L
Jlnk7cltNJzVKC54UwgBL040LGOd4772SrG7u5mlfmz0gvh9dPXxZ3lDUDcOlzGTeB6r5hkyJZww
6QuOBuY4IQBjiaIFM2vBGnabba5X+HalEeSTHYoJ3rHzvq9J0yCezDyah7pScHBEU5Jq0HVqDhyh
iNeQPRHB1nRDG4Y5cCZF5knIFDZZTteR+cjZEbCblfFz3SdzHyheLxwq2WArXO0du2Um3C9Wxagv
LTUljndysUzmuLoU+oz5tj/LpTj2xkfX2dOk+vkWSqAx1j1Yqw2ksNLtsI1DbKPS9eMR3SS3u0GN
Li7AqF/kIA83YnYu4CaodQilK6nWH4HjOQMIrpqsCPSgONwpCRzySL2ODYazP5+23VemJMwaqDgX
3ScGpz2CNCrvzNXbqhIZ68q3ZSdicCK/a+is5EjzwN10utkzmz7DYbFPuC7FXg7K/oEWopgMJkiN
uBpLId0g0vunmKBCHf9g3cGiUx588LwakTJCiUKv06sH38372s/HfehwkRlEKMr4kMrKhznm5OoQ
5GUcMni97OTBJQT6nldvmRS41W7Z+7bWwD2eePPqHSZ7lDcS8gXCuL26xPFONhFmZfnEh+6A8FfH
OjsXzrln/32SJ9qYM6SHIUn2zlLLzYmiaqb2EtAnF2gByJRmkfzf/vfbg+DlS/q5RjPIDhEhvHja
ID4LontEZTMboPFPjHapeMUGZH9pBhawl/UjZ68xv6z38YoBTeRfrus5+Dar8dxIi6dUl6K+ZACu
kVmh0VLpyhDgV0kGdN8Kkc1mVM9dj5/A0wicR9k0rAjV1Il7KmbHdtrVD1oxCoOgIUM6Nvy8ya+Y
JW5B9svIHz7yVbhoTG2SNEeSl5d4KZHiFVfMlvZ204LzYhu+Jf0JpuKH1cgUkt4X7BMI80FyS2Ez
OEKFofOwC5KpoXqRNn/r3Crgj3LlJO4aDzJFflbNHyMV9ASbfrJPszYUr+PLq6z9RVXvv6A+k1Hi
6ZVoLf4exHSVWD1brxeRFBcAYuOFOXqGq7sJzVk9B8KslA3VJC54GKZdDi2+gxvafUO+slFsfgJp
9pwhOQ89XvabwZjBxWYDEry683EmK0xGU9ULg3E3F1i0MQLBVZvpCm6iHrtuMzGWEZsK9Mwk+K2v
9Y4nyF75Idet4oEfiSz3sCgMXofHYyZu6Txraxs+wBfTvT4oXZJN8909KS+drVRHYBL3CVrh68Ak
rVPsCD845iYTmMmpeJVcrqjWvxTVcpbcvowrfdZYJEsHUMjZGI9dlBuv17fZYebHPrYwqEaVPaPq
VkomD7Or6W4yi1V11m/s6+tEswD8slusZ5tWa6OM/V+eir22KTe9wPQTWxV5Lab+K5fFLGt3F1oj
01Jid9wXLPzMw9WCCKeGMu7yuLRTcgcJjXmsyqxOVNupxHuRogwE1aM7kHs8EMHo1dY63YL4J5Sb
uq2viVdl4t/K5G2knkW0ibI5TK7J3s5E9gQvh0xzanB8oW9objiHgCBn2Xj0nKtBG5XpD8Q2ggfZ
JclmlIwjVvlGxtpum1OSoYIoq5c/qaIHp21RYGxRmqfsY7SPwVbWHpSR3LdxlYGmH5jphEtarF5/
V2j1R2CMCcDBu5eLgllJ8EkLc0BJzCm17C1vvUHbnnYpC8eI//8WysKsjQQymEn+u6fkwVvu0Ciy
kK2OZvxnmpa3dG3mQIGlgsXQiARA3eNj6IWB+IzOWM4w7t8/EGUBhuOskjCqQ2LADQrjoJ6T6wfy
V+ivgT2gM++k5CbgArf3H5XV4XEVDOMOqbKC+SMFNfonToQdZEvmfoVunPrZ4x31cPpKl4N+mSK4
71rS7HuYYytQu70x497XZiqhiF6vMtJX46bY9V5k7/K1oWH1NanV2XTvRl35S/JGBvqsJ00Y1APq
3O+G3f2u9b6f1w0OlTVCc/8hPF+6Qi9SsBc2ZaNb+JMoVvdJ8jRqlbbq9tO/RvziUHGCAX1EXhXl
wqm1qmzpD1EnX1lJTxtWJauwLKfAnOZgP4KKs7XoL4O1pmOYeIdSFYyY9l3fDTBSDJhtpSH3k9Kd
ka0GaD0vja9Ze7hg0nxHXmyCRTs5XBtcr/zQfinJ7Ou1/7L9bQNl3OkGj4v1O8s7q5CbDMkkC6Ek
S8QwCKu0OC1mA57upTLFbGgEIhAN99Ntp90VqGtMReVdJygdOl0Qk2L6/Rcl5C78xTriDi3e5h1D
YFwmORoFoAY9X5nmXGWh2JSuUotoHyv6bxKDQ3baIjYpaCrKI0ukbKka0N5S8i+ZQL1qryYHmDVL
cZVCaIfhD2/KyYIgNNptMP1q39U4OLk0RHmgdZMTDIiWKyZ6kRzx+vH+TWDuhCunax87lHF1S8Mz
5zgCEY3fxAl8L++Cikb7nARXChyb+MhHPNDCRcNHhm+Mb0cXiFehwSn/5GKdPIpTmfMBewm+Iz1O
i4anRNzMPoMz6/PI7D4ffUGh0LjrC89KeCunw0KgQwiOnqe/ic4jFWfa7IcGo4nb0ba8QqrygfRk
NDGbRRpuFUI6S4k0O5roX0OrkC6/jJAJvbgzxKJP0L1/VQKnnHZe6PbyCrk6wyZeGHZp4qovfymt
easZ/r5CtVZFucN9uD0MmpsTWdxo9QDSurefv26jEQIZd4RXD1Xj4OLMvfUBKpHeXh7povt8a/qw
Lb90KPKZVbT2tlvmZMIuSTGdsIDNKiV3izFuUQOzNm/PuN5ZYtjwTZwbS7kUomOpZt/xhv6LV38V
YoJQCxDxO/JtBKm6AMqVkdUdONw2SYzWU86nTAbPw5BcJkcG4aK1Ui2kis0H2UlxlgbsgSzt7FLw
pelIyBhe1T2ULINGdFRT4OxgY2pM8iB162nQhKxishLaEXhQ1hMNcdW+8lBJ8WTlySou7yK8n6OS
rIS9wK4PnJDrX1vWDESF08uCsDNO+4gDhSbEZJUKcCbIYuK8OgJYvriUQzf/8f5KkiFUO+BT0Slf
rOJi586n8WYmlqCS5TrL3C+3I31/UKR+6ZD7atSo3Y1dKuz+Ut1zDaCH5MB5Mv86i0HRBMMla19e
PPoSLwvBfatAP2SUIo0SIXnn/6hlWlP7Q+V1bbkmPqkVfVN9eag88UhpvAp3B9H6zOEN6J+mwupi
0Xh0iZoDtBkgKMTPh9m+hXOuebiPoTxl1/s04Q6zfz7hMNjcX0TCG/nPtSk00RIJfPSqznMb2vCs
ugrTMlvDL6cGn5ffmqasTZFCkhAi4eRt2QTIsLZd1NpBae3Sgu4Sk2ehlCqwsLNd9psZg/DRbLOs
sr0HyYCw4yRWmlJZch8hT4oX6swuSQv9AEAJG5ihJ1Nse2lNik3BRm0ssc4LF3u4wvKF2ZZAOh46
FtmdNsybzF/Q5DL8Y4Zcu3EGIezi+hiUppMG4RAo4fGWQXVdZPFFsRvuYIb/99gRntdmOjXdLBOL
u0WAaW76Y7qkeAvLKs1wU9xfFu2EVRRQaF24damGVOuc8wC+MK8E3Vy5874GiTaSXcxgOsCWSYuZ
r1QJId+FRR43r64ZQBEj4w54GDpSAhqSrqFHGksHQmRfjudyze0Ty2/GNiXgu1CRfcNW4qfB1Cl8
hweDZwNBUBgh5TMHPU+ZY5+LOVb/x2MB0H/GEJSwuOf6W0foHW/MDDCjryarRmwc02Vm1vhFlxzw
GgbxOE4t5c2S3BdFU65wltKE3S28ViNEvbchMHHJ9FCBU6wXEr5A/11MG0+h7zkXDqiFEEd/nhyr
z/BUqyM1SMDfWru/B0+VRx1e15ednestGBF8209W5M5oqaLrP3YjkgCqY5wAtr4v3e80nMGgRA9w
wHi7oIbTht3h+7CGenRqrHrnaOkLZoEHcdq8pgdhlkq4GcGOX/SjXF/1OUgOr6K03ZHOae6v0HH6
3K6WLibq2x2UkxDEaqAPIVEf6VtJ7nHqvg3THhg7F3ZmlMTSCLhJgPUY6vwZBH5RDa56nvrJY7IK
XQU3d8HM4flkGxS4AavvzNoSLAVxAunuue0LCueG0dESf+HjvMjOdARtv69EFGV1ay+bRu6rUM0g
CbrnIi/kHWG0jfbI4p3MxbjgmEHLE22hCYXE2B0uV0pipWFdDTj9BMfGwsuURuOLGSrVeZDPC63T
5H0CexB/MKWrazalm5heYnOiZQrOjG0335A5xmeWWxTPDQskEXYS2CFM/hVOtxcpA6y3I91nE6e9
3BQV36DzLqVmhhe2+Bi3z2sS25wm+yVe/0j9hRBrAmx/K6Abcv99e4+J+WtG1rjeF2nvO8dY+fsQ
qWk9/66TViXVFkFFs6mgKhBktGBgeQd6GEoOSvaCaYjAGiEhxL4NKipxNNt8NDPL3op/OXWtZ1pr
QPIxfXKOeo0sG9H8hoSJUXmpObBQyIviHR0CcoHdwulW2TqsUhI/jhyhPMsIxy3UwSOFlCgWj7hp
6ahYKQbcx4/SJOShrsNoB6fMhwkwPPkVHAlyXZY+RqopyOS6FLfMyH3xqSOAJIhYRT+nOM0IOp/f
GPURo4cDKqjl9oquvRBJAHY6W71tskLZz+t/rL9tIrjGX61Jtb1FO5kmwIll4lsyjrNVgvMWyOsi
2cw5aTP+6eN+nDgXU6SRKSdXJll2UQWwdj0Frr0UgD98+59DUc+WL2blYxecWPR1qXMmfrZXafQe
T7cRKdkXH6VytYNp2FEZtm6oxzj7AlybF9OK2/Tcf6GBQMqRn1sc8XaKzDS+LBmVggXE4pv0tEAP
lRuYBmbUIs9Ed+lQL66qOvVyHkKVd14U9+6ois7yI/+SEczhSFIqfg15ruf9ELOOcoQZWIqeh2aW
/9CSWDdKdY3es/BMeImssL/PNWMJtgjRNU3F9WSoJW8eASIcIUmNuisNc1j0h1+8AcUZj8bGdva7
WT0niJfw1lo/OHaPN13hIheyeBR5w0QHwfqfi6aJIi6njcY/HXXsuflqzwjWMDvJHB2j/FqJMXs9
mK3XG2dusDDOXozyqXPNGVQSHkoqIs/zouS4Vnr0o51UECr/RilXCRVxdkL2G5qgijKWwRneQW0d
3oBkv9vSUPlB4hIOv2aePtYLgIfdSI++zUSTlNEb2pRfY/BeEOYOSle1Ms/m/M/Y4lsgvDmYGTRc
30hDGEJ8162FuAaXfCCOsN1zj1q9njwh6n14JylE+P21F6T9A5uF2XKOBpvgoe9RTBCYhTvs+ZQv
ZYiMKyamzd4l7BaKTZltS8+uXfkqZdL5jc0lVo5X3mNwtzHT3PcavjS5JOqDf3ppMWPEtRrJ4j5f
85IzD6k7BT+InFwq3ipmSgE0ONWK7wGTtE79+5jb0HD+3PZikSmLYs0i9Ic2ZIpAmg5ab7jBdffy
Bcye8v54Hb4spF8iktcL4Wsh2iKgg9X4RVujDqCaXnUdFp8rRH6Gqxd6iRunHY6sLiZptDANO6Su
rUfiNdFMncy6xqEXVgYrLyaHxATAoMSkxmYaxds3JLdyxvBS4uJBSX0oWruRQczsCOhOqmOiDmkg
cjpJMpxr9/xXrt6pVVkafuZM2LuKxmTrHFXWOKbrJ8rP5SAayFJ4QkX04uRgAxPGSXCtjrIDaePA
OffXZYCdBp5GiQ1rFYRHU/13x3GkvBcNapunrCX844R/PqxnesY1jqCWXpAoNN4WOyCu3c9EQxYK
4WIkienb1vFtJxoIy4UfS4y4pqCoo6lMvDO1ELRzwATJZYqAANWyaueRTwPWqy3cg4JItSdW74DK
lLN0ZO4ELIVfn59Qm0c1XFHHTRXU5Nty/7al5s48dqeDKDoIgeJ+kH4RqpAcjZm2oLZR1RvebD06
4jUygVZhWAzNJT4XscwDP/eacW8egjGToYv8loEKDXINzimhIPnwSIKE41K6DCtSCXlUJ0WEQnkW
1I5lCTcg1Rf7u3giUD4xqOYw7h034vVtk21tufP4hzwuNfFx5rwc2jnYcDIu+0tQcTk0ezXUXqrs
PHA713DxYwB8WlEdCOIaxlfkmeSyAeEx80MAtwu7PS6NeWrCP1BIC39166oqzA5XX/Ila3aY7vso
ddrsxZ/XB/0QC7e6sZJ8pZO8Hb4AF0dhrr7yGsc/ZiQXKT6L7G5v5EJI1h810rP5HEEXWRDt8tQL
UKu4oLnuujuTekBWv14oTjyhizL/swlqEfbfETGoQ+clW5OAmIKhulOmt2c5YEHd3ftiJviuD8+J
Lnd+L9ni0Doj3Area8FIVK9iDt431yAzOc12YMoWom8wPDfS75f/cLUbtVGWgz2BRuHmRHfQeq7e
laqTfbRCd+tjnM+2rJIyVHurf4Pp1oq74NGhH4pZGscR2HFO76UdYuF0/v8RuAbty5mN5Tzqli6U
SctBNyEOtyFdTVM6+2B7HmQvI7xLc5h4xw/W57Sqeh1DV3CVzWzWN1ZoNBGbp6SvWNZX/tjVaSBG
6icUj02pBd/rOa8mzDzXqwCPb2ZdJquu8Wqjt1EFtltenIbW1kbcd8c7RFKPy5gshSxshJX4cOIs
44fJiDAH51+ejHhrJiG9OE0HALiKHzPACk2Oq+XzwG9j61sKda/ctSG3iVLkeqv8S1e+6prNenS5
MsTK74blDgoPRo2wSvRqYdVKxZEa6J6+mFCBFKLGeorE5b2TUN3ENaPWxFRl7Id0RDgSOqqmWwom
4M84d/zvyVGCGGqUfHOMJWjiK8HqBiPlw5MaOAgttYkEQ6wMxikwWkZnQgjbVe0L1xqM8Tv3hSSJ
MtRs1Bec6fVXZv6h0x8x7B3toYpzhN8v5ioA18QtSvGFe+A+s8GETfeuU87oG+82GGtBZLE+j4TI
FPWGqV8NIHBh2A0uTcRU+jmjCegVW4DXNXVjUcSsZztyTUPYJnf+vD/XuWy1iNz028OlElGd0bMP
lGS7KawrNKBOaG9oVUdqTuYLSjmluAMSF+WfJEhJENTzTU59pXglwd59C73tEh2Uy7faZSjV7LYV
PSyQedXMOHWoZt9mWVwkFeCVOjxwiVjW/iEGdse1AcByKfLQnlwcXwghCMbSIOck3ZmXCqXDw9KG
0N6XbtlDMYHWe/5v+PMO4hgAEEd2eWJlF0+hyXgYslt+c4qN68eg9x7MWV6xMpm9BU1bTIo4fiNn
niCMb6wzr5FQlJM7FvIdo5soJe4VwLyMvMzfKoz/3xLN/duOs3+NhpjVQiplxbbnZekuJKN1wujv
O+WfWj7sX08JgX0XHPWkU5mwzS9mpCG1XxDQCprfA8QDWqXlxZH4TQFkgjgIJpsurAaoEWHXe37R
U4zIaVhzszS4oCDojMxBLjzfbOIqWQZuAfLMd25foXlToVzPu+TEg+F60eQRb1MYA8l7SF9dcN/T
A5ngMplwzatwhg+m/7iJLZGPVeL+h4eLRQlnM9zCzD5rkUY8F6bh+o3S5UZPeOCE7b4kxcdKHcuU
2GxDclBJWQDk8V1isxUVunZnobT69dMEjJYovErQNMHYG76gUPw87dA1YFVVow9nhngLSC4UhYEj
Dz95CyHkn2J1u7ZzDfibRO112VrBixwbP1HId6XoKjvf+vCbCzkb+NaY5iQX0ZcTPbmU4RbpYUM9
EM6lmNxWOQnkHX9NlZywmyflycZmVSpL70+/qv3I+FnVTesk/MMqi8d2KLyPzOH2+F2o5W5kH1YT
RJvW5BBzJHG7KjjvRblxXBhZE+AkUJQMh04QxLU5LvJSumH7DPLfSwqRKIoyTnzg8A5Kivyi3kIW
vWZYVn2qX3dDoMIY4liihlAtJn0G9U1sGUsCq3vn+ON6P240zAR53uZlsgKTzRvX2bZfgsLo6TUS
lrAG9WmG2fBvAFyNzugMOnmAR6JbKLI+9iMzZZ0uEQ1VzXitEckZKmTepBWnQ76BkXRzB1hM0Qi3
0X74xoYCpzxrvq/a5SzByUnTgyi/jE3lMl5oElbiAeEc9KSXok5/IRfCYo0A63BgnIxkh0obST+l
ObdjWng04qdaiQW1q/SRFpmUpGm48wNZoHPyUVFx62AaTFnQo49iS/Ytxpldy0uU6m5Zsl7JjXZA
LQlb/KYqzT3EXSp6eCRQDOtMcIwDkH+2tsmheCj0hevNjjrx6Woy8nTtniXeTfKfGAGZhruk/NZ7
icp+joA0V50NaO6QK0X2fp+kBGkH4QyliAl/WhUrhCIqziHgkbr7Rwmdnezsy6KylbaNQmAu644Y
IgJoeGM58zfoHh7y6xl0x579XuMq6M3MsyJWlGZiz0j0sn/i8209EsAAb79Bw7uqvYo3zOpGnfn6
fn1RBAX5U8EnqcNAi1yfO1+A6FAYCdj0Px+BhQJ7KMtpvnaxGV0nZb4zDHLb6PbyFBk85kR/JCLU
UXPRzUWhQHDVwHxDX73dlmXDo+l4Dqdeu5mWFp/ecCFWuIcjLvsP11JTUHq23qDwXCie0gSqI/Ml
n3hj994L/9x0jlpgZyVl0WBdAGeOaBlkdvRLrrK5dDdAfI0TAg/yKyg1v+4Yo6rwhKdNaQkaxRY6
GM5zcszY57y/oFDfxU3k8VcBOEea29/Gf2fUYk9iU3hAhpoQ2UBOHiFmTZVdxgjT8st4jA0yh9JQ
c71b/3OIXNyRztUdOr/NEbpJBEoDh5Ee12DPjv1hUvo18cymVAyoCQftYmALl58/v+IuaR5zOzpX
HAOHxWBMz+EFmMlskZ1ObIKuywagNKRohNL5GbxhHH9u6wGJ4d1vJhOje/jdVKbhWqp4q4rv0GEw
zKRUe38KK6/YbuzKU+MGZ6L8J8X2uFJa5HAMeQdQW678zUkEf9GuMT6JkBDDvNVjzGYA1Fqh1Rc0
E+U7/erjltBenNTkcmrjDSmosOEn80LGTCl4wRyFEwqv8NvNcfLzhO8lc6b379csmDBr3hcNvL6D
bPNvFqc9pXQ8U9IWcZtQfdULrvT8q201LYHh4u7/B7AWH62Hqg7qqAPEOGoE3hQz2IU1T2c14cj3
Z6/PsWnwLdNvSKIixINmzsDl4aYgR1swYPgGLYhhxslhL7iVOwGYWPYKJMfz3Ht+ID7LOFT4oF8a
ktVWHYb/q3TYKKeIiWmcDHZS247fuLjQ+YZm7kK2fyOiJneIHapfOlD7uIdZoZZoS9IbsSWWbYNG
8ussbbBRTmuL25bNTwieTkVnHS2lGbSmjFtUd3gykx7+gBWdfz8J2GHSFq2+YfZVjHnCR/cd6S2m
20OMMV9lqCXP8Ods0nQkav+TCyeV0wELV03E9aogPnVeE+QEZEnG5vxfdojl+ik9f5K2Yhk7CJ78
9APWXoH8z57OTw2uP2E1Den98OIIgBJIu/74HcHYbB2GLmEBAC2YVMOVeFD90jNhMz6r6RVV5L/U
QquZVCySmZLOPw2PBQplZiWQpGgrxUCqYahOXOMqSMUlQiZHco+j+960dpzjJkO/PwTb2RoCXDfU
CuQ6JD9b4Xb+WS901/iV5pnFmz4Qg10Y9P+a6cHUzJ6gfhakCNGyfcb2aCzAT58OCRyyIwJ+106G
Xw3yHIzyoMediDXyTZR+G3SeTzIXwZvm0DmKavhrO2p+QPJJDOwb/Q+Z14ElcBfZXv8w0LBckfeM
NhJH4Ut64HDRPRv7S1YuS5iJAR8JaB+Fjamh9bKGs8R3lxh/ueyuJ/OCegcp/Scg13D/w+q89sMO
/6G8V+iK8POnPAMs+/kjpD0yUjwzcDJHTrxI86t4fHSEknRNgLPJ+THspgFxnrUtWmYsyDKiKFOU
0veErpTOxhN+C4Hip554Tv9MePTLNUz3dtLaKpuVpYdz9CMbxPKAlrvbLCaBfgOn44gKTsvP/YJQ
MCQpAh+EBZ9DxnZ+mTnG8oTILtH08noG8adwSBHFSj/Cj+uLXPVqkJB0wzUOFAmZiAyb6S18wYXX
AplFnmBDxWpgSfFKKCU24qRx9/Gs4SfaQGJ8AkQrtOoTZuMKWueqEEt4saOA1a91fwrhhCShT90t
pNx/CNUfNak82ZQupG3g0eLnTBX5LZo4smlVe2t90CXI7UD7aHB5GUx+TZ9fi+5l4BLO1WmuX0vf
nbGCW03Er++jYzccrnUxnZsfXFuSdtIxCxB/8QPm3NwZcUzFIHMXHgfj5wanAi51FVd4rqoEvSKz
oQ0lWdnVjgZUu5R/qI2fcplAKuTjXQ2xFmKREXgh21J1qB/wb3z/1hEBIkrL8Z0QLI9ccUUNxnQ/
tc8EQuPj898W5oynoIG1m+DHmZZEoRHvAI/pT5I5xgITtT6ptquz1x5FMoORZoS+JYkTsAPeYK6d
Jiwukr3374HPOSbR69lBg6qprcZvYsKISRSY0fXDkCnsyOp/E7saNTW0+qlUqCVDTtTeDe5LaAkz
L2YAjulknqNikS7EYiobQGirblNcun4BmNBMfc5JOOStve3JhoVLQmZueErCj3piIlcNS8s6osC6
OMCK8Rto+fXt5fAy0AO8F01H/aAZQrntIxd4JTVkgRFEK/KXPHqseW7WsOOb6OKs/8L0uw/0m+AP
W2y6PKNTTF/9tH8990B9w0JgxM6jFKtXNmHZIT7LvV6y3q+Zz803YxjsSjx83yf8/5ZAIO1/mWKt
y9tnagaAsxC5zMKprgKLPXhJx8c43y1qeKDz62VA326yQqDjPYNxl9GX+qXPCB8gYCCcbxq66+Zv
QPIIextLpedg2PxrApKZDiKbyDetSAy9R0zXWLEjxVhqwJSg0w4PzcLp0bsuKJDBCgi6ywx+GQvY
pyVlQFT8T1FQZ+Xuz9keD/GF2jpXLp5v2+AwbOZalg3OyEymsEauXpHhqfWI1E/H2x57et3v0PAb
ZVCG3Y1HdRWW5p+x6oXjrC09dJ9hX5S6trUPdsYCR+jH4n4rYENEttIlBUBMUWy/EpAsGkFRtA9v
qEIdbQor6KbqgOLa1TTraEZXhEQCIVvjFW/yFDQ6PhxjReVC6O1Z68fSq1H/SvIcZxYS20HJZTmN
eBFppezhhkyikXxbQ/iedDXprbqh2MKQ8C+e1os0cCH/9hB1yCkk2K42QK9PjsWHSnTI438+cREy
dihyEwNlZl4BeBJVmjc3YvZNjvInnDRzxGahgQnK6M1AatDTx53d4csqFenkNl0NHICgyntYcMBv
/AE80sZPjU70or1w9UCI9thLlglJTLPguIThvwb34qqHseKejUErxJNvulkotPJI0rIDQSPH+/0+
nBOyM9qlC0roG33YU1Z13qsjzoFoM8FjQHhYwhnMBB0BdktlA7EmrBteZJxDlh71p9zp1Lnv7vdc
Uxq33zDMs6LxZzoYhRL4QUzvn9af5QeiFUJGO0OBseQBwJlj6Fmc+8dBZ8t1+KfuvVB17H6EGZ1v
WnKMasNQB50y3NEjbS9ZuUI+2V9x4i2IYSzAigesLsdhzLag5iKKlv2zWbnIpj8GHIKTdqc0SDFB
QOWvU/W23yg1IgyEtUEhdFJUwOj3FquV7Q/3G447LRyJ/JTgQ3YS/nFAa1raI8ZYPD7gUGtgNKxP
OgGeU06uf937WvoROzeCE+PRPahi+95/+urDj6GfRJ7PJqEcz3bRL10gw4piySxZo2c0jDNbrg0Y
AgKcXw3C9vaQu+TxIsa2UBj/7+Kx6g7sx1hPqDWG/4xz42f3ZRmCxhkfuSh/bDessEtDmpKtp6Vt
TX9Sq3mDRwY8UThaFhGXvkQsSYR9ZQSM1qTKJJJXubbQMbYoJL3r5jtw4bwZExEoosGZNSaiJrGO
+AoN9IutfSDhDd+qJZDS+f7674MV8ncYpEMCekxCjR13M7sVMI1r1AU3vBojBiG52wiOvvZ6rtwf
CP+KIIw8qb6b6tM6h06/SuIcN7MiczYaAJqjQCvfuJS4q+/eFPVC8hJf8W7kLCnutK1R/TgjXw9A
XrNPM4fYM7OwPGeUndPKTOuLYrd/JMbLC92iCQlV9OCJZeTotEcvwJzHuQes8MXz9vYt2arliFiB
OcQbCh137KHoltQ8QfZFGQ92Jz7T4vE9FTEr+011M5G33eadiFiFxiAtBuV6vTsgXc3ZciO9s0tk
jd8ANbTZix2uVK8icGumsbZCqUqH86nPjlzP8wk77R5k3xYMDl64XaCDJdq/2z+B+R8nyYVK1g/4
2JI0/K94jwB2pgsU8kU/c9aDFUROIOiABlnd40rvxOvnT5mjEY2MAaPsBWS925RKZdn9/Ji6+pDB
PREtfCq1D9MNLaUfRuTrYMp3/Z45OiTPZxb0qOk4+MkE4ZFUZgFBbDoPDrk4sQrsxkyIExsaqLlt
009LXSjrPAOmrzuNnf2JaymB5npTcgfZXQWml2Amn9T65tjlb1DabsiZK9fiEIXBpdnNl53ej/yR
Kue2ITL30Pc7wqfehhB1iWkAkRJIkSulpOCz6hLFKqPF1lmy0o6W36xFaS8evM4KUE3Wen70a/i0
bjBW1J0BS+psdsdN4bq55cK1kf+UFuUSpAkBX0UYlBEhIliCHCFmAzKsfymR0CTmzwVFTM0TTsIK
Z7JB1oHsnSKsd9UBYcSEkPrrrxoiA9EAm1HAUtgvh9Fsg7asm3WTeaUsETDEej6WQVUkM74oEX7g
Us3zwfbuU35TddutebCr654G1RwGbzy5wHqDVdSbewH4pK3ZzcEQkQFHG/mOE/NH9Yne1BEz05fe
aqJIvw93lLyFQkraYV6nmlT/pPCRmKpjoTgvdg/RJwd3HJVlgkEyFObYbONmB2RDq3h/RzOli9mp
t6i3sfwQDK47kgpRMpWiaRin3Tz0vFU+j6EeuZYWDOChEx5qTHRjYyWgN/KpXsNPvQYM0peRKEMa
J0TMQFwUmuQK5e6FSqh+p92D1DFyNiHW8YD8xkmiysP+ygtXuManBP3gi6w3Ey7Lo+ecahrYt3cS
waXqXLMQ5fEzhNY/MmY9Cp6TpDnpFfpi8Ix6CJmIgsD8u0XL6eCproDby90SV9YRV/1e35iFeIeh
L7m3iDN0Nd6JBuf9uFFJu21JF1vX9Mwg8wa9vItw5QpS5gRXH6kbBaUv1l217CmqJxqKxj5TFemo
50YtiDmV9HgNHnGBI/c4ME35oNGM8/E1TMjC6mFh0uZEBdVNheuNX/XiV+qJnUIWyryqqQNKsuPW
VrhO1LPMYFLfm8PSRmKsJWmE+GFgocDttcB6PyhJ34kZl7o1Bz7hXcNbPWihWmOR9f+rGr0duKP8
vfVe5njLgBmbwvAShgajAZmWeYddeaBxAQTJ5TGnlE1GHDxfvQoTRIf8zSvvWYknlHdQwMld4dIe
aQ5ISFKHwsiVLm5bHBbuYOR7jr3Z/jhGpHfEhUBD1+psJs7ArzxXfavjpkLNFhPevmlKSqF0jnll
5WOJ0Z3PxW4NodErOJQZTGoF9Gd8v03U/q2OGFcTrKJ1iYfr1dhbmo/PNXty61GQIs7I4crY6sZK
pZhgU5Hvd7hmxQxtnds4FKmjoACEpgEYGIfEou9+ENt7XUj6OQ1kjyF0Lh0ZHB0wdTJ2tYdaW9jy
7zKAO7od/dmWV6boRaMpmvqJFUUC2h49UpVD2I0Z4NUYHCdIaRJvXA7wLJ9cle2DawTUJiXnNaIZ
HtoPUzPF/KFlAJEHx9mj8BcpH1fOBae18+b1VwxTvPsaRrQZ0YnaipanWrgvz0yfn7FD3NbhhTCo
ICBFUQI01rTDfQe+38sMME9QdmUABewX4bz37uGywQjRSOKc8HNcksyrKjCgjwJV27Mno/zo2YOO
3ac1MwN7OmV+zmE7Hsb1yc6i+2YUwsz1u70RTalhm1OyEC/7Bf/yVxyE9eTnx1duJPrJTVxDc5Do
Vxii+Ycah0JBuGFyaoraKFRaNTbCpwANHPYbxBo4RqQhe7/CM26PRbXn7EdRfXfzul7R/4h1tf2s
RQ2qKJ5VsKJ2xogtfNswDRMarnOL6fzvsn33EAuSb5QD3Vfddx6lyGdUMQwkWGK79Ottx/R2wl8V
8vMpct9hEIjbs2n8PvxTnVtlXDiZej5cSbr8yPFvhRFuIFE4TQkRqEyfD750N/7ewRfhcHpN0FIT
sVVXU0tPL0/i5WRH6pN0kaX6X4IdToOLN2BS8lQdf8SuBrXwTa1XfXJ8g4y/O8WzZz3xaI7fNS3C
zHChA7j27hcAFMTM+lLYMMNtjLJPiRTtVUWsgEnp0jJHbF4TgF8EkgX4GrmOme2yZAyPtbvJr1t/
E60UxxO77fFBX4p015Nuin3tgejpKjgPYdoZXDTvFXOLrK5rpDo/jAFs57QM284/xBbugsFUm6lx
wKEBxcfjnuLKW8syQ0haZOBmwdbUOu4UHlkm0q8mgoFELRmesFTsy3/RBitBPAla80rQGgKnEp31
7oTbdh19b36tf4G88EPHKZQuWmnki3yTkfXwZ1bEilaS87Ike/89RorY3YC1LcW8f701VDipVvAY
WidRdss91agIz2I0yXMqV8CB97yQxmWtdmtDKIseewrsJ4dJ9l1j97HXU3V69p9QFKat0nmJIKxj
p9znex3kDO30nSTn1qTsZlZiCRZ/dl9B4JmmytshP2ZUenSQbBW82RKEUHv+DLszLUQsi/4u1N5G
XVI7q/L3jTybktf7/oj0O+vjOxlvjybSSdAYeNog9XpnfxTYoShQNX3BdHj5bGv+qRfKAw38d/cg
X74HmnUlt6k85EtFl73U2qre471WIH0kWxH6dXiskBO6TyMewd57Z85stcyir4TVDIWII2wyCGCe
DUYCOlSH1nw2ehpF6ifBw3axszHog7NUH9K+IGSt2y3g5hOZdXZJfWv2VEmoIKR0Y3myERUumL1A
2JwiYkO8W5aoQTXunQDQFY0wwomG1FJNj+Sf4JoPRF4DOdhzqK2qoa2GKrmrnACO27XnMERibvIx
dOdcOx28Cm1vD2ACxDvjOBSWRmQ1rr5imiheQ4+fv6lCwrjy44mhZu0nrWbs8RfRRvC/wZjmiBRA
htppHZyFuuxryaAP8Cr2B9QZxoI2Us/8j7iNe/W6nzHsTf1TC+MPOH/2a/O7E8ShnjUNjOMGok8z
k75VaLA+hBu84IsEpU3EILnsO0nDoK8I7H3n8DcgKJ0db6+wrq5bVxMK+R1Xhu2thFD/gD9FKAdz
cpUrR7mdRgT81772ured2Q0irCAaRcAkz12zomiSMEx1b9Rgu54qzCzPRQN2e1skOFuKn7F29pGE
7ICWI1gf3QknUFLs2SklflRFe4gDCjNIkoejB5e+id6bVuDcdqJOc53DwBW31tEFMem5rKz+M1KH
6T69++cb3wbtcMwmbKFdhU5+ueDY8GY7KUh5g92jowjeySNb5mu4jmXolp5ycauzbK8fwMD5AHFE
Ot9H+P/+IpGndjOLUI4yGVSBZL+D8OV51rupOzeVTH/EajpZrRhzdW4pP2Damz/ATryyY4PFmc5I
+NfwlRmQywi8B/VWQGIpn/zSeKVQDMrZeqQ4NWrEBMDZm6JNO81SN3LG/K+63Q0fhxMm5JQRC0Hf
qt4jGz94PvCC5pC17neKzjmo6m3OhIhnGgBabVqygdpdnptvpvIKCKbH1lHMDpfCg3vrWbw3X/Yo
ki4oqDkUvBSRkiq9ziNHH0gdqM9Np3aiuziS69N/eWxRo+0vX4g10Ye/O+mvL7Ap8maq5BRsFoy+
foW+QtPE1TfQnWSxC+KK9EVC1nl9Az6qXXCroY7jNaIZ/o9v55XehtcPihU+tJBspobW6w2T0yf3
DyqlKbZwMUpP2RyzWRVJ830VrtNNvvVoodQCKsR03LoF2+cbmj7yWQ7EO/e1Zc6Y/zo8LmDIRWpI
aQLCdKKZXgKiTmLg2fpXib/FK3YlTd1I8q9LIu5tdaWBYxjQxJ5KIQ/BMdKdDv/NgPjCIv1EgNhS
VK6qqzMe2R1RnkzgTkxYGkbkRIs6GemxWdVCSYA9esdmS2th1p/3Za41V08HT9Ctb+Q6yaSajqfa
3KdOP32/Rp0ca0sSOsAEuJK0xdh1c/1h0JaI5iOZfZhXMLWNPw+kqtklkS98KhSqObuJnJcDjoK1
jzPlgVMpNEYwtjjA4NajMoWT0VQcGgVljRdTe2VOE/YgjjRXj2zeNd75OpX34SFDsXQzKQqPD8ny
vhfGsKCoyojXfPG/1f2DwhuWF0WIvVmBwUNwmgcYpAG/g0rOHmQC1HoDOzpLGP+A9C6e763KRu/f
0j0tKpP6L8MYtxHID7KTPucfY5HC4T4evJa/NMCiRGvZ5hBz6DVsjw8yyFhZzVp8LW5QWjGGBZAH
7GCCHFyyzv2XrqMAdqagbNd4o36L9PlkfcP5h4FTQd6RJ+TNYliFop/vU2AyGxVhXX7Aq3+p38gA
/89O6IdxEz1tWkO/cfuocKQSEfRmnyfdEhBNEcYpDj9NB4Jh0UZVlGUJMCDHePy9QGvBe/uTkM2C
rRo4z+fT80SfQsfAVTP6aeOVmfS4BXNpWWwElxLrJesVoZz4ksA6JmJDrUucrHSYgAkZE59MYPsh
KKG4siQyce1oygnhZ5lHncB9bEId996Sw6MIAZgPyuTEYQRar9lPmKSLW9CuyoQA3+TB3L4G6/1p
hSrss3lc/rsb1moDfvb4CL2qzsv23cxUfopWOqaI/BsS8imvN0IIReNITMHA4MBwcpPOvXcg6sVW
7jyQsXWv7o81jkGdarvoniyYc7+hzqhla2+XI6yOVLpfudlhkaVgBSsakGP0+0Q0K5yQ8Jq2zP+7
86tkUIhpJD/BjaJD89pFKO9Kf4YPK1GtMl6YWN0iq7USAc6Sm86u7VYr3jX7bqEEib0+ZLgsul/o
FPKO2hcuvFRL1edevh4q0JCnhNWT8RBdl/0Xce60aakr9GabdC7Um2AK8yDaGJlBgcW3PRgGaC2F
d94RRySQds6LH9rQ9fnd5HsIJ8GF8sPV/sZ8O1zltNZ7rfLJ+JcLqZ2fasnv7cEd2tHPnJ6243k+
iz4RGRgUI9G0mxfCpcxhGFi9aNMvX56PNT9W1qY0YltoVOZiOG2BeMbijm7taD3ZWJXBv9UwayZ4
pnIjMwHi3nppNZkE+FwsIQaFItsQR74pQng6QgjYyCe9msBu5ucohOZ8U0f//8VR9eu4J+g2LpuA
6Z1qHxO62WbOpTmyG/C72QEAFSZuZs9zdQWYdF5+3JkCrrjCjDzB+nIWMptcu3fkwcJXDmxjHkkp
u+HlDpyOXRZRt9lwDVK0UlV9QkwvDPdhVmdhtlGcAEDyVqtp76ku9pDZENS+AyiKDbyZvlcUv0ST
d8nnQh/tuah8zIIX3ABE7cpn5FHjj+9WUK430KNWgLSn6TGaE5GdN6z1o/GMIO2Lu5c6Zuq7F1TH
2V6YFQrvsrYE/z58ih3Cbd2hQ3ol5yqAR9fBchwVeecN2KseCYvz6FNFDdT9/VfYsySkCVfziURW
wfuokDCWKtHEwwfGByOSTTbexGIcJkx8kT4KY9nnr82I4UrzssEr5z+mlBOI5lhshWjT8Jelsd9f
t7+L3YEwpnQfuSZLaWSuiAv6FEsCL7rXc5b588mAYcsCNVVZbE8c4qyOANEJYMSG1IFiyp74EnUI
OVzzRWWIamMEkRPsb02XkEEmTjmJsZeAZrOssYpwMQ1w574YRI3+vSgi7tblCgyLxC3nBxWHfuoB
y89wUjxqmn5se20myAAYc4ATSdvCjPWFfRuDxxEKea69ChmHEQrQCj6bwweA6lW8QgvrwbmlmerC
EptrcEmlIAWWb9DKTLWEZ9BWjXp5hi3OLS5zVSRLRWo1ITx8q3Sa2u4590mbZsa3Go+ADAWf25s6
pOAiDqou3E0cHbgwfW/fxsgKWlwNJcAD/7+xmkMDyiPbWqFa68aGCzF6S4XgMVor+giSFUi8PdN/
HGEaOUsWXBmXmyy4oeAXEHssGZkIV+RHcFC+z0rCDmdhkRkCOoGumCoHwuwnrovWLgrZTB4s3K7X
Eqm/rUZnNRbMETTXOWkjVweafTothIwhwsWLY660hNPAMBRdFOTKllJY1vQopcgqWzCj5lX400QL
TX1mQna3k8KO03rMwDgDgvldgTMoJ1JmBmGqHTJm83w41jhdCjzpKfookrEz/EtdTeVNX/kANEwk
nASwDztt3bVELyeWK4MYkyWXExBJjVJHZyFHPh6wvRK1fnDZD03UpxKSELUPcoznkPd1LMOe0o0X
/mm43nvvcb4d8sMFq8KHkFgbyqCPHISHKZJ8y9MDRnfWOZgjq79J3gH91CW6q0yFFe3gU/QRlJzj
aNCmFhVT1MSosrhWEVQtP5gcwigy3fmttr5uxmc0hwZALL9WofFx0Bu69uepn/cDhNRuCojuXnKv
XRBYiV6O9x3TAixcJHhReJuSVSz8VcbezIQgQC+SkZWO2BUzqep3Z9QuWfps3MTEl7jD5781LZR8
wJZTtPagwuUsTc+1AqRDod12SN9mUj9A4e3NBBVoBmp6hZ1dP8Ug0TDdURjyvn13W60k1UnPbspG
8yV29K9ctdRJTzMfey5gs5l4YrMOuvtEPOxmsE/7P9QRYmsD7L84x3HyuBBayULH5XvepylVFBey
5Dgsvp0VcHYxr+f3+Y35PLlAeBq+UIFC2vFiLbbUQGYHAbKEmi4I5ZoZ9Oio38XymeepchUWrfAS
lv4jZtE04j+mA+A24XmkObFR8jj4ue5uUn4v9A0HsRFjLTEDTrl66hoLGJE/XJYUvM4jD11zA0w9
43B4IAXibi8tn1/omdZW+lQr/DAFfS/qzi2HdvgCUE3FnpBItt/TDBrG5ajjOnBmzhnVsWKvBg1m
fmMGNHy9WyKG4fMVFDtZJpOsgc3hEjfoo8Ij4fN8wt1U4i3k8mPzHdiT/o9SRwPCHdp91PgIxMor
pSWRltFvbnHDoc1ealKA2RqUhwbgzqwrEveaJQA3HguhbDUu/pAYTmuVy7H+YuM8mLnQYAT3s82J
1wlj3sUYVPqT9tCAdK5C0izMxrYwp5/JdLNaNrqpqAA9WQeQx+vuN3vhcRGE0tS2DP7HVWnukp3T
aWUZXxYhQqv9eUV7FM8Er00xRaxArMeHQk14wG20kH/Zmz0NyxUKYlYq3TU3RP39tRDCWq8/Q9pa
GcFNtfMT8ja4Zzcx28OCyT7FGapenxUEP0rlAAtJGj8U5t8wRyhtbcw58953PmeQbOmb36Jb8Maw
H/HghNObPUNwVkC7D45RtJsVDBBCpwL2IGZ9iDGspvOkRylaHn3nMVToAB/UD+3CcGksGOxQaqlf
klEw7G0b/nIrzbTEaZHwvyEykkpdMIZBhAxz7xXCI0gSpCF/y10E+CpoYE8YlyImlpxPR6G3Aw11
UxZTlp97GoOFlZWy9WBqB+n1aRJWaF5159/NTdB3Q1TcF50/8Qd306OUO2D4MJbyfcKI+atuiB4r
DByNWgCbgnMRQ0mDYF/k2zTibp3pS9fFqfZf34Pn6EFZTTeSa8qe96TuWE83f4ERBkGJ2mJnbB06
YgjJ9TQwY3l1JnK+dvw4qZlRFVIZ7Flrp9SvsZFAgb7IVxy2hlje+a9ODXstYI0oXc6E3VnDMhqF
EfylJ1weQsFfmU2bZYPMVr5nt5EpEAk8IMJ7j2jMoafhHRMSubZyZP/gCFSFb8cZ/nZSDKjqX9t8
69YXvfEDylKPP1CY4y6FGy8N+QRMZLak9XUVi5cWxFdorPpM0FP7k7Ns2cukQIJkYU14/TxeLEXt
74HhikqC1UMRqXqURsYo5h3vh2cphZ3VPqikviTXwOp3UbhW5UxnIfzrwnSaggyE0c3dr650lkju
Yi0b6V+arwRsNV5y+RSR7Gyi8CB/CnbAukSMdiV+9L9GkyBQfusvGDnfEKRmNUhFtT4uq/NYOfno
ji3kA1DqT+sXt/64yuwLYzLJUSRA7YuWqCvMabFi2cWobwOcUyCzbmwV4mOQSpb8ai0arD71ux76
6UFVzvVkivQwfUqsxTsJkW/jtP1sCXdeAwPxxWvR6Bg7b5kBgvbViqI3CR9VomWbn9rlq6/2OlvC
7KgUzd+q20o1Clgo6NPZOHtoLiR9Wc9EtIic5BXvbt7mcqMVe2LrLOJdQYQj2Uvhwo10h/sdtVmL
WX8g26cFxvA1PcPxE/T/W1vIKPgf/DPNv1F12rY/B1w5WwTrOtwIp4UowL0/UxOXl/UmnZXWezcf
gtamZwi+qKD32QcDE8JAk2dn6IY9cTIit8K28OHxEHTZsEYEFiQucVYZ+4t5GXwrx2CWVrQRKyC9
Rb0wMM/xntWjny57WgfTAH2oy2FI7qHgcQx/WWQ1lZlxru9UQGjUYy5NNMPACW5TecjfG7n3+NeT
znG9gGYXOfzqHbrFDp4cEZ8HknPghasUZNRCbxSySSeSpDZLbymjpZ8VNI4S03X/yLF9ok4qf75P
cmx0BFXukI9GZwvsDXkQmP1ttrzJSgWkT5Hy3CFPjsmrY3aXHIv1TeR07/mHXE3O0iO7uWMTeCv0
AE9gxoaOwW0SMRH8At3I+eJH6hzD56mYEhWadROc9q4ZIswkJGIQm07I25uVp9aLbwM0BBqFKD9D
07kywwKyoUN0gHf5xqkvOfxZhaWqbfrFFLaMNBQ8L8RspjFWNdNfBANnAmVV3+da4XEF0I81leuE
QUH3q5ZHfBWhtyipCx1fLxZaiCKvj2Jo++kWuukSq9ynMBltrT5qQM/jVjTc23PyMblF3nDm5Ft5
T6RZgzqAtM16dTv1Gf5aRr6Mw3hSv7AZxljgBDeYq+feXQ+kncXomI8dMERDlFCp3K0did4jIhGk
X1dzKZJslvIXaGUl/jFyKNC+1ilV0Ghqd2Qiq8ykqieCawnJM8NlpnSTqzM2Nat0+kD8/xLCMhV8
1X2i9mVko7lHnot2Ay2+qZd5oh9qwvZlkf6vvjcHP609e1V0zvEUNJOjP1C+J7WMFa8RX2DSdQ1u
TeNgNtsT3fVznfQAqJqmOzxSL5cdo3pZkDbQXeF3mxXZBMJ1uDZXiaAF7cNZxuK2kQuXrLI//kL3
WsxkdG9/laKkX/P7YdskR4mhijNS/yOQOb/wmwUDRdjC5VapT78kKXXh7zNH4C7GOnEJAcaYlaxE
Njfn9SKkEIjvhdG4SGl/AcHsN8sRcVJhXLGuFYHbNxeTmvDqGsvdLdRk6z+wCU9p5iW7q2VeyrrT
6gok03xtlwc8BLmrlcOOfWQHwLgtb3QNVZdwX+Z7591vh295MzCpBRt0ESSdwTiqqhg5FX+5Nfky
xrvDcYjRmxxkmSIrx287yEpf/770cWprlIAvGSPH82+2bRDJbp6B9OTmBk6akhf1FmcVv6d1qB3H
I40JyujylKSj/z5hExscr9ei4GvamnYMOWBfpQfqmNrY7+i6TtqOXmPCx2Jvggsz6h7BUaQw//6W
Hb77b43p8UgzH8ac2a3Dy2vtD5IfEifrJjFMzr8trJfqmpR+LSfKUDvl6VxfFEL5c9zsQhGftWGv
5U5HGciOrXCMgQ23jWIKoycDXAFidUBFBJjNvIGIV2ck/aZVZCBVVhpATJYYWO4MyugphzR0dBd5
iOF6IkfevnFVaNbxe9Es5mPja5AZee2WKZfEMe/hyBSxQkeN4x0v7lgclk1nMU1UTJ93wB7YfFPn
ATZUr2extMxOS/HS/bLYf/cjmkam378IMlvek0IuB4NXifRIt3zjoH/+c/SyMLQ3aoDQrnlkyIUQ
2YT7aV490gH+yN470t04yVuQSklZEm/CD27nxRZ4oLuw7+zvf4rJrcLZTHOjHEAp4y9QbdanH7V0
15iSoGCPPPF0zfOKnkkK29ClyPK4xEOS1koFZtc6P1rExKnuU4M6xv6afN38+tPjHNRYX7LD/rbz
3ISWRgxLd57EWahaeek7CnKy3OpI2BQRcOpgXP2dlas0FanHQQ+Y8SsVqFZmEH7WVqaA0fYwcpsQ
hosHSVYdx6Uio57usbz8+EthP90rN1vycoCmJJcGc2+Yp63c1GdhiUlZbD/PS3DidEw2ltS1hqo3
r0H1ASzXrx7KlrR6eP9q/UCxB20jf4rrJWga0KosBiEljmSKl+VesZBBV0qiQAEDdPoUtSLh/01P
cdcSwCv2gfwza9O0qYwHANS5R7fceX1xQgzrEqvQFHgJZcbJiDzrpw5d6ZI1wnXkNfT/JEtO/u+R
CA60fHWZtE2rNGePVAr0d+kBzlVvFc1FJ8kGcNE1mUUKq2rQifiNUvXRiAGE/f+Qrl1cwlZdhGv0
ILrI7iJXEA6rH2yzAtFPlEfM+xOyPUvF4fDCML1LWMPlXsE6PvMlTrThqxBJ+vSy/gjJopyGMkWr
5fNUwM2tNkO6cer6uIsIaYpw7AG5tFO2wdGCwLkJw5d7vFhDLEoq3k2ZlWXG5UuHpCaovFZVo3Nk
jXW3M6TuILHaPwswGRg3nSYL37zdK8BbkvNHV/vkFJpRh0ImeKZrWsB2ipNgx6ImCN714QOyHVjx
lLG7odYxbVOqpNnJKgcQ2rLC1x1CIbs51CiDArvdGvZkHsnJ1OP5gZBsPBfofXCkh8Z2NozoWIVT
RgNxCeXDuEWn/5+HBVpJJtbtOCbMtJngMtscTC+P4peHq3O+yJ7zhimormuqiLIsAeot2hVR1PIs
sFgCjcdByjfjkVLIrx/1lrp8bK4yBZbynIxTIOgbeNDhNl8CV8wo6KRYJPson1tmz/GNFWnCF0Ts
KOWu91m8U/zGC38NIqVCi1WHRtbVpPqQ7h1kw0r24xoXqtx8+A16/arjdXMVkbM5GUHMO05+0l+X
gV8MQIEDr/oFmSjVPEAnLBIpNty82QIjBtJFD1flC3qPlLiW4MgYLBn+b/18MTkqReEQa1hTbunI
DpDt03EA+DhQ4Gokj7jxmDIObxUALQbrU5I78rRi3HeYY8hcT549pWAU05ZGNBBK84BEhqS1UGiP
IjLQpTwL0T1GwrCEPzUlVL0xNPcZZ/EUyyrjqNOYWrfMNS5asQc5sWvyVeL0v0qBVW2o2fq5/BHj
e8fIUBTE7J/XLcL45UjdxeMQn8BfJ+yi6bOs+B7MJBSfyyTJemx/Ikcps9zEVoIgfm/NvXvPSWAE
Jh23Aed+w7g3Q0QXhHlpmDNDcjbfx2HWqTYIycRm6dzI354RIpn7euhhyeykaldlqGmH9a39K7eo
xWsJbWeebzHKr1FKJfgLA+dc0baIhVbu3UNrsbybMO3EZfACiacv1IzJTtCbxzEqoaFwAhqQa7R1
/CQrhrQVTa/P0Qo8kBZe8VXAEL+p+sfXedx9ZS1S0nX6wxYHjHPmGq3BM2fP8w/P4vQx3tQNYRAo
JusT8Ty1aRhwMDy2O6wC1OifYmwLhYzhBL2AxJpf8ZlSRxaKPkenykvXr0mkrMWDEASOcOqgyX8R
NbclaIfnz1rVn8g6rrniRN8lljnE/TC5dNQ8bkXoeyRkzSV+oOcD/LpP9cxmcQRkGRuqm7OVEptp
4fmNiRM0N+BPY0mnUrw4wn8R6f6Nb4Ze+58vmf4eBYKDqNC4usQ3BtXOz3adYu24+Vcb4h2OJEGa
Uay3SeuXgU0v/0XR6RyqSAd9nssaKKxi39Abr8AjXeE1BtioP64mVMNJei1dWr05iEYophS2WLFO
Mab7QxVCvMto/8LlsBnd0/KHTwpjVDHaShHq8uSD2YORF9Nd9G+ybddfzUCHeGyxg6F8GLwrYlBC
cBrUQAQGG0/cTmNg/lg8Aorop4FovgoouFhIZAl2dEp+JbwHnK5ZVcYOS0DslocGdz/Cf7s7H6Lm
+uvmi9kst+vs9wFIFyVSZAKjQ+AfRN/Ai8T4FVfMeTQhCsotE9mZc8LfxZKh+cLc2bx1db1mxRwK
OokNlPl+kCnwR6gJKFqmDHQAhsTCfPCVBjnAYwNxLSispiS5aMDGuG1d3lRTtnUsBQG3n66LUYlB
QFCWUciJNu4UXtJ9h361fHWGKt1eEpG0s7zcSI+0IZVq1BBXWmVPkyjLt9Ggk7tbZKF1KeqT+9vj
XVrlh62iyOwD1w1uKmF4sjDAtnw+l9JhheBzx/QjES1sMKjOESXepbZZn4jFmCifLGmCTOexuayA
wu1D8XuaWAGyJrecUf+XFonKhzNQ/yJjGB/iKwUtGu2PKPcfq8kstw2Fmo3RPSgmgGe1XGaMw3pB
APhyNZApncGS3QhdoIwiGj3q3Sin44HDOnhoXd551tZK0A6daoQsRx/EgUSk/KbgqK6CHX/OWc3v
wPpA5DMmQ85D7kMyOvguqBJ8Qs3uwLlf3OoGbLXgUjEtOpxQBTUdAnFp6pAUgtUQIG7QdA1VF2Gb
JsCBO5cvjxVSbhCfwjXO6W1IqIGkxBZiP2N22xAao2F462FhxU3E92hhCfeO1j8QLVtvdpDigqKk
hx5HlD6kn0bRKVA/HZEVpCvORbha9T+FpTYolPHDEbY2xxdqi8XJUByda94LbJ/kDIlgIqsBdTLf
2MG9vSu9k2KCGFvCFGQfs911nzB5LAwfMmxp74mNMg5REB1s1OOgZGBEvj2M1LovxSDh6iTg7tqL
S5xd2hZKcgh4N/KWGdMO+/Kh5LkROxIf077L55BNH0Qfm2aWoFnW8H7o4+RHT6S6bOJdpwkyp93N
am8wKGKyRNBjgEOoVSt2z1fkEZV98mLU3+X5+Wl+0tR5uCMDGF4xFstriAy69MQCm2zeEEQ5HWi4
o0TTpQgH9CITvjbi8mGxSTmm2nR8222BPi9VGtgDXyMuiOkBUUHD0tRvHAGgktSVj9wTH2p5g42k
s1h1GP9B6WsxE6RKPN8zHcRgY1qLR4o7CqH9kxmaXp5r1gHzXRSlY6Exjt62tbt4eFF5qOPXpr5D
wCzNZ6U8isXFroKFp7Ntb23DMh/8KHjFGhxDk+cyOuQaQzVYUJqms+VuIcImObWqS3Cw/VZdScTR
4kKtiFUqGaSVyCzZmln36GjGxUy8ye+f6ZDFZYLTyYB1aB3qhj93Yi4+ZkMIyxZGr1gY9uFSX9iJ
VwTuTtTcv34NsrwS81bkE1XwAy1SF2Vd5TAKKN00twGqXLSbbERYDL7hbH7pZh3rm6n2+MtC2/iV
txHbvKkapDYyef5YJloJ8tF7fUbdsYGKXM0dbL2J7wfP4Q3EhMAQhlLGhdIqmiyqiMfnu0Hh8knP
hyQ/wO5pMXHnuv+NYCKxnQ1QtM9LbXE6Nuccywdms3EZe+6APFdRGKCAXYaPh42sRKGFPrEP2YZU
J/ZZAj7aBbJpfNKGzi3wn36L4narOgxDr7ox+mgKmbDe0s3QIbd2Thp245xRiegDDgDC9qql4BJK
aD6Q1n/EuA5ImCm1eafuJBixblot5DsLJZ23UqzX+hFY9zpZqnL5hLErER0p9kAynIeKoHKFAyw+
ybaumqzawJ9UJ6U12Fk9gLTEeGL5qXXtGzoih3zwJxlWK/Dr/yr0EH3ysCiThbBUhj8Fc3a4RD6J
6pYJuTiry71EYwLItkzRhZj6Shm0eySNz0Zf3jVs887yWwTpguCK33q556Hj9Cm7H9Aj0//Glv5U
79HVQsUnisjR/7BoTy0IbUrA2LtRxax0XmUX3/WcBP3s7i3kxCcVliSt7AB8Z5dyb4U/Mjk7i9Qj
JAEwViDglYTjxlnG+DmAs+nrBmlaXJqnUEwP4KbWWYXZhl1XQ9S1SRuUvR00d1TUnskOhdu9/mSG
4SFFlVem+LsjqKP7hojpKdvvMSBdwRr4jgxZJ/ueQ1kc5v+pFCbgCzyvhsvLgiLx+WR7E3qLPLai
yOUZvI20aIlGb7aH92JcYxrGn9YlyEkCqnBNK8nTrowwDQrMcoPCckggN8j06JDAXZLcMUes/Q/C
ggj9OWtPKQWQl9ZjlkBjL2tIy+bdtGQmk2iXhYNxSwV2yYIAqZCCFNrnR/CW6U8bwIipzc547tek
Udr7D0AsbVMxHEN6rSxVKSSnMTq7Nf20LUxf751QHePA24MlfdVNXIHUSvU3yW4gE2fZXHJrZcfB
uHBML7EHMpuool3CSkbC/j++9mqhv1jgJ6S6PDg/IRikNLfJkZtJLL0QSA3LiwcPlZVb+IoRDfAt
3JeZXEki1t5v2SRFaVTq0/mV406bJWJsVF2cQcoU/+/U74igmqkD9NL9MWZRVG4Pgpc3FJJsmVZz
iX+z4N5zhVUzupX5s9U3QJkOEc73EzMr40T5G5Xo4NFgSGVz69bRLsQcCHZ7KoDgL9KtpX35Bvrh
oxbeyKqYup20PI0rVf+eBFH/la3voyPL908gy/Iemsn8FlYnXArqolLU/IVdxqR72duEJsykca2r
y4WNxcXmHLhIdmotJaENWw9VNAOE94nZbCmfeUZC3VOSppRPFegzD3SNBqqccE+HnGBCemXeue0O
rDORSQHk7LKTt7rY4gOHs19NvUcXlBYSOSzyDO9jWRgIye/zp6ibBUdmngYuFvhYOGYUtVrMyL9f
ClXBiA1Wc6p09v2XLX1VF0FHTJks/Qga3zbPCWPILoXdgIkxg/9KJxrW0C3RDiK7ezxxypV/LIG+
F+m53BteDlRNioCVzgPcEUjDlXcpjYGWfIbbXdz3AUWBtHNd9G8vlLoyuxzlXlOw1GRXQjpOZvJH
tlMZCHnw7wobhOP9ym/lwptowVD2FO1vtmoVUMFa6mnCHdR66fU+uByepSKlkJnUhuTFCUaXD6SZ
4a2DBpqa/6K8MF+PcKMBgWpcM3/9uhvLrBPUsQ53Y0GA80DNBPVPlwT7w4rAtWZHSMxbaktRpc9b
wNe3oawFLbyxTiErXym6vs68a+b1q4vw44VZD62a4AJ4tq3bg/paGoMcjhj3hjoBkCdh83Kuj28I
Kg6LSrvYZ0zJlWkqSXYRrfSFiglXWp8VPdQ+ukV0rm+RNmqd7VFzQOTs6nAzpRwlAukO06RR9Epg
jxi7Ur3UDJJsT8pvD7V7XpTeo3niwfzy7JViuJArjpkYwmQT8LEJwb2jlrt9MqNKl0kllEZ/eLir
qEN+oqQvzB6LZkijT6HQLvS7ncRGlsYTOFbFR9j29qjCxmBFG61wh62ymX6jsXZ0S7YCLi8E3JIr
cwJo90d6SkhHyrfGuNGUNFgCYcqEDK2B6w/Pj4MledBp9rJpMjueUUSG4pX5zzfa0aacywzX6idK
0wJa3BxYfMBHtEwddX313keGX33zHBvimWJi2R+KXRZaTbHV3ftnUJkV5C52OCDZ3Lwcr8rYJazz
tR8MFTaf+zDmKI1EkQRKfijYMBD6oNfcJiOJPmnWq3fNDqa2DtuTc3yUm0vCZ9SEKz3y3ABhJVwH
VQ3xZ5qtnFqDjyJA3IWMd/bK/QZzdC7zBdlgyoqFBEmFcs4VJwts6vdGr3vGbQ2SfyA98ERIlHAS
/7iOS8Y6ycY9J+rwiRZ3FEdYO5W1bXym8aXUDa4VdW6FiUXyRhsqphaldrgITK1kDsNKH6R2rqEr
0mO2pzEqvo8clThnW2bvr2bZP4aiEIwNTjXMPE7r8DKPTAhX8aH1IW1Srnp26nLXaVhj18jhcu2K
U4pYAPauCbcqHcA70+F26cdB6r3mEIdYwTBwue92p7hh63kIKKro3ocmFuDElSmrS/fVgU68tbQ2
ALW5dCMIVUk8UOQUDfWbNNSstXzgB30LxXMVfbkG758mZq9sJSbYm0ttXz0hJHKxCf9e9y8lHX0b
KB47SpJFiA+dzdAfq7b/jRJgZZ/E453WFYB47SUFM45lpZley91SCJgxFGlIWzSx5pn+VrVGyBmM
LAB75vO0+ySgEK1izcwbyjCTS+LV7wZbGnDtc4Jxd6Oxp8JtLFUP4j3lfsL2P7KQ4d2UsI+VBGeB
5jQ69keH0MEZcgvVgtpOW1r+CjRJkKVIBABr1iyHXKdoLrUCF+3WHHORoySUIh939evSOVXe9SIG
iqlbGNyr3nPUEKK+qLpcSnmbTiDWGMFhpZamSD+dYSbQ1wV2ZnS3SxbbEM8GbBugPGyaoLnUjrG2
4OPPjwKgQT3VbwA0m2pzmHUW0tTgwIfTwMlm2KDiDOa+5eSrUCzGaePWR66N59bnjU76cXWBdgN3
XSNKcgnF+yjz1u5tbFZdyshgsz/VnibJx21MdhBnznxenaW6nwJQgP88Zw7Lv5Gs6d9Hh/DUz1wQ
60a5tXECGfwnDhYtCqyygop74jLAarpqu4xv5W97RQjugFfsYEKMSUnXweYzrcpOHxZ4ZwoQWVWu
h/K6YJ5Og/fMsxdT5qHM9kayljrP+0zeR0ux7gDiwsuRTDRhwml6IXk1xJ0wXBKrVM5CUF7D2S+7
eK5edPMa4CCc8T+vLfTFn1Rhk6Vj/2WMQ8WMyMMZFHiftf29mq1mA5uudOvQEDlqTbBA1Wvh2OUR
gVEtet0cRnkN5Q2NmmPdnF6wakixfq9qoJpwE2+RQnHusiMFH7APlKGIkh1/hXM+jaIdeIjwOwrf
8DVo/3TA147zXlEV1/7TGX7VX6UTXgoQht6MCpKWn19smzBJEjgizAwgFNa+ZZQAWNHW69h+L7e9
5zuMYFSZYPWsfVh13r98eovsfS61Up/INdktKnDOGEZ4y8YeTUQ8173MAjx0+64t5VR74p4pHMNi
uQNySQPnywInXLwJqcnqFjMh6A7AeHKzjUpQvs2z1hzTZyaWeVB//YTTNftCxbv0C7nYEtgpszc6
Mw5+Z6H8dzp5Gm2nnmyB1UVIDhRIFBlUsk7V4F9yD3b4DCo8sD8nZajcBEDxwRJoWjZ1vJ9lz0Ea
P2iAWizfRNG+X86W2bkRJ9nOlAF7e/ToQZncIWFMl/Tb9Hrkp4RT+iVn25zULvrreFkJe3JZi6lD
NNQsAXSX4TxIH15WwoKROeguLc4hOWsg5rUD2/8S5z2zr+wiDmqyH1S2+9wfJrA0lacUMBJPYn3x
n4sPkPm0+HE1xgRrdyD3sjRn7y6y04hHEERyiMfE56MoNUrrN5aPgdNcYF/7SSgl9WB/IQE6DDjp
cE08HcV2v6CdHXv/hs+Rp/l0p2OdGQRlIpYD3SaZq8vqc06Be9k+lTtrJBKVoy/iAr3m4Chs+czp
92P5vM2wgnzfU4AFmsZLk/AUeYi8iwfKU0DocHr6Ldeo+KNdwrRb53M+p6/C5RwXSGgEjQjtENgZ
DEKFuOqVtxejR4bATUFIGj7lC/XilGWteIfbNSOKOIJ6Zh2KUi98Xr0hIxpBMHziJ4c+zo9FpiDK
FnK6jtnJzHv53zZJqfoZdVarMn8ScJvSLuh2JS0kRVfktCo3HB+yb2DCsQijBdc1phSkTMDCFi6w
RRI5FHlI1FX+8XnbwGhjaHeMCICqke9r85W5X0zenM3/a0MXEl5BIDhtKjbQszrUlDj8wbUU7pzK
bgj3HYv56BoVyumEL5aUAWftyDJOhZgbqQ7utnZzm1Fu0r70UJ1nyh5T26StXQ5ja9kzU/S22zfA
jc/Zm3Hc6y4nHLDyLm+pICHxy18binpGOn833QhOX5lc4kPjythiRTkOuX717doThxTRxY/klTsx
weJI9qJLCmpKk3m4g9g0HJ41lVHHkfXCripJE+KdB6Nn/a2VEnCHCTVXmVyPUHCT2EHYGcLrkja/
1J+yiWF6l0ndzjaouE0Z5zdlm/o/hmMQAeus5ROfhMmrmwOuD+R9tV8R+LXNebyRyOqDf6Ip5x2C
e5JbxxlvlcNQyWfLEAzavyv9nlnsnESvbPTFSTzn/Xf5RIw4FpASSba8D54c59BqHDXSEhWEjhut
0KbELZU9iBf6Al2VtyU99RDtufBWmDAQmI6pTdNEh+hqbYnvO4byMh9nCFF6Iv7xJ79zKqJfs4mh
1wZ9JAuFx/EiSqlC8xj7ROasgH+hufylLSQ9117nlFvASW0D21A4T6tdLw033kyCKNhrBJzxhrPK
2zwPp4+6/gnSLEp13QDuzgwBEA0HYfVWGw0BQM2kWOtLH9nocjfTI6sDVqi68CEG4cFjWaUoy7yV
M7Wme9wK+x6YIu9MAKvCKGSWrdmXkH0YHrz9Ya9OINdw47V/vpCAMyrl+I6fhzYo7L9xItbRsNUK
RVrai468QFRCAbcLnCXOTy9ECJ4YLO16tvGFrxzlvX60bfERbRmviyyiVAfmmf07QSg2aFFSHDMm
Au9t79JnFGELD9PmOPGhjKot8WzJMFPCkB3zCUhthpagt55mNWjDpp+NiINA5ieCxOBZjba9OCRo
h7+wQSHYs29gaph1Jj65kJw/rF5nb5aWAW9IucLXEcyesuamE0aO8mUzOhVP5sNDhwibr9CgGg0w
L5gixCh6DqNFBreTLz5re91JvCoOxDftO+RQ/d2VFPbY+NU3TUjU2rM8UfBJX2W8KIk2Xi6vsYKO
3/RY9h/TB7wBH0GHmjZ25RSTzg4CmhZ5MFpA5TXi9dTmgL02tX8ndGqyLANiSaYshVdXpjqB04uy
R6a9bHOq7TBZaPdKKICLvN0QYYXA5y5EmA2MOeLVNBkNGM9A8lfl0/IaOhN94nGU7zKfsUNNlqqR
zPwHziKoD5yKD07KpIqRdkcMLs6ATjDLH67DmaJuexT9U8DZW4nTJPaNgemJMHjAgV99HP7WyFju
llihCt6MUrn35WK+DJ3wWBEb2EuwPLug+d3mNnbkz6J7yaUrmfEjMWwEaUI6MyyhBLVMhezlo2V/
uDSL7JS/1c9PTgaDtXoRUucAeKwl+DrQ0M4z2zO5V1hxS+IxOBURc60SwY7SkZsCA2zO9EvmfrgN
qgaajFhOOkIhWae63JrEYW3NpmQUwLCcPMH3VDtNMN957dGpxKGcbwBWdOVeE1Dr2GEtuQ2FENpD
vYsKN04b7HpCGbiGiVZNzMX7pp/5KAvZr0fRZu1QSeRDFYI6h3omIVOHoVClYsprOAhYRh1Jo7hH
iIRG26tsmN2OPlqgEYH6Cw3niHnCJHILgXs+A+EYEc4EGdofRDIIXYXMwz2Eey4Rsj5fTRYzsF/u
cSpSMAgoorbXgksMM5QdqhnSsSwlVEmNr9X9XgdWqGkQgQ5CXB7TDXdwslXYHgfcXMmuGptjf34l
q7SBZvsvoNYv9Os4xGhDcKQ/J4JTIeHUQOKVrFjrPQ7WJtizprN6abM3//d1beG3mjjKgb6gBQb1
Y4nuNxFnIbWK8hXGRjpvwOJG8ucvIDcJqodJSOTRpdSQgh0w2lzACG2jDvASI3fO7oiuTtDC5fkd
4CpKVDDs8KHTBpSn0XFBIlU6CR0Ct0meapR9bYO0UTlv/4NPwLPoaF+MjI7G6ttgryJmissvfzpk
GuxD7e/042A8ejKstHqhNbe3FjD1lx5HuGy90GS3eMC2N7pBmFxeEsXHkcTr52oEzi4anDAEPjOU
+DHDJU6kd19j2DTnOFvF0gte01wAap5YbwSPrltlcirlyphNOoWqYwgEIyb8TwgcW80raW9vuM59
aclV/J/4Mv5wOQSA/93MkPH64EGoO+pAMc8Z4iaKBXzfJYUerVPL0W3FN3qCQwlTO4TG2/8qgJ9A
C6WVhKPiVYT3WQ8FCt9jfHBkIpTpK65pjPbw/egOoKXU9PSv2Ny3+iRX0fwo4TUnhfdyJlbdFFR8
F9oqDHVaaFm2Odtx5bGpbz/rIQaYyyzXrix5muPhO3dE28GrpAW7Xzbh59IUiIou6uF/DuXoN7dt
u9V1AuIQMkNhBOheOxYZEnmrS3ySUFes25DbKT5c8wviO9LhSyTFTYLeEX7XWgbzb+Pw2RCl5Bqq
AJhC3LxtXj8wBYwX9+bUdG3J335K2U6rOz/NB9M1vs1JaVvax0puVpQnNEhiyk3lzRg7NlsgM7G6
WJ4bJglQ9APwfDDnc9EfRfW1GIdL6Q5Sxof8/PhM4ZrsAUgOp/zWLqO6RFlTEGZHAZncsqtJdxIh
Wcj9rGEv1mbZDp1a7fri1TiMW8cA9ygThAct56bUDlUb+fypLIjjx2TSJAYhO4fGeHllLC8sotyo
kJNbwBc7unSWrE4DniTedjHZ03zjxZsyD2xzszHSILSxePkFySlRaIv4UFMoUxeNWGKIZSrWwYQN
gwsr6DN+WMtGosa2Pbznlqmexb2EPETzxjaGHJcxQ9axWIt6yu9MxmdcKIcATedIaZapo+sgPsek
5WK8IwXcD7WoL7v5YbgWsZp4Nw30CTVmO1gxE8D7C+gNurZrdTnosiGT+E13iywl0yseyYOflP+X
iUkYT+IJA6/YTSl/Ps2CuQbLQMDUf78OaYHLdnSfBA+Ffd7W6nVETtvWzvDEDVFdyI7gwt/wiEFJ
IKOgKNhHrpyQ7cgsEA3o91T7/PJxGn+N5UFf1AzwcHR8VKxOPhexoSNw/zS5b4+wkVQL6yl203eD
4m0VAuptJYzIg2VnY1ofIDtSg3d6OGjAV2X5CjkNCQpnt21LSBAckUAu8Zjxd42NGinD4WDzqhSZ
8XHsX03vCoE5Tmxv6FBcippnRTB36dvnTWSQo8/uZr5l64q9hSwZ66ID2KAuPI46hA4Y1c0gsuWG
1Rw8qoDvJYoGpfwzBMEqoQtKM9LDNHF4F8FEaCfBWdKQH4IdvlZkcpl8io6mWZvI883QAW7kH9aV
NO58uBUBgLvuV/vfY180JsTmOyHvzVR+vnAMvgWT3NJZUAGjX2ghZo7PZFKQaYT9t+QWjtgsD62v
d90Fu3WDsH2aDp7UVfPBRU7/dR20ZnIfIcpGXP7B2xEpydmeG9DGd2TSboD9EALCbTp5AK3NpS5V
T4fVNmplBccJB+YlhNqompQtOMtxWhrIXDk5Jjbi97h22UZAeAssfv6W8cfJpuHxc4c7cHTVQj7S
ZlOUhanMwG6oij9q2JlkT4vtsg3mYwA8NZSLLaDEb5OFUGVyuooBFruVxG2dhXRVHlMGz3TXi2QD
qvdwXkur0H4xz9q6I1oLH1WfHZ9/Fy7+QyQYyQJ619HuNn2Pn8FufyZtytN8Dev4/5+2LVVYlvFa
P1H0cw1PIDYqzifPpXfrdhIcQpptfzwjr3lFK5f36zzLk2Y6BhFZVJ4VdrBgpxYxRRp4pPhsPggM
lvt/Gw+FAQPUpHu7XkMnJAqUyfqgQzMmrXrJy99maTk6Sc3qhLOkQvkbkXBhQFxm7Rp3o/1aSwvG
RizkX/LxFnCaFbKIyVjtjj23+EsdOG6/0GM2MTYMiDhmf+YpNGP5wu7qglkNqKCdCPyMdmzocN+9
avc3KXvedl70/tR3+/9RgUSusNg7URoXkhqjN3SRpfM2UzXQIHqAPd3VvZQCOWp4ChUe8d5Q2MVF
1gbOL2FfCIawdahUMvNLfsRUPPaWRNumuwg0mIwDlcVGVdHtFBVS5FD5JAI8ap1jTBIz8yWc2P7w
3LUBvyFA9GEJXXBMBR6dNYWBVo8jM8EO0oYBi+IQydeRC1U4PCfxXpHxCFSmcbLh+nyzgqPYJ7XI
d3M5tuYSskDgcd22BKJa2M8rW/R3WPLlI19APpvkvem6ybYb2p+JW6+GX20AViDaoN5loETgJbQH
BqoYOulvq/lTtzf1Dyrv1bXNSNRz1TCxWfbBuDftmt8uaDCwThT9WCHva69NAc17UM4q0qlPLTEN
VBBMFnsvENU+bheGgr8HoD8Lw9xCTnR8CRwoNce5ryLUl+mAIZQvtumXAlIdaWb8N/zqputlmL2X
UGVLgiTGw27BOwpeSNDyxEnRtx8uqnua/HvbXE2W4Qu0KqtP7K9ooq9BalKMEZI+DU2bTUJq9qDL
qJQMHtGOcLDp/1TMHanQbqjlrzeWZqi55GsoecvwpzPYr6hGyaR9v3xoWwqa9I3c9tc7alsLSKRU
pIilxpSFzoLrNAfuCUnPfAg3XJK1A58kHqs0g2PoEdXmnndKQlIY9oEHuLXOcD4A/SCyF/4t9oQE
YKAXLxFmkxaDy6bZaOrJNXlNJt8jSN9h0RPbQadI0aL/SeEGPwEjHY9y8z2fO6e5d9Rp37gBB2M3
Xoyf+9cMvWv7ykBAD6dUSZb4pjXd+iAhOoWonci5H1868atdZuvnSeHISwubkpuEY8oGZHojIJmH
JbqxwDLkLjbYafceaATPb7KtQwW6mXfrF9NWOk3VKnfdwBk2Hqo1DPBfj5gfbFmmZb1YH/liZdfP
udA5I0WqbnzFHi+FdAzSNq1tVsPOEhDr/vJd6Y1mSKU3eScEUrZcEHlUBcF0PYTwmjTyItkIdsRq
G7NvowsEDTBcsIwACMkEMBNG/kAwlsz2/RvHlf9ahAH7sSZTjARs8cdpGW+rxTu2nCR55J2vpb8l
koEoSpOjffOXsXl6Hrq2rL7PsJ2GzB++dnpq6Q1YafRGGKFd6eEAcTPCnD+zZSsPgjVtggcTvUjY
eRusafR9uQGJKNM0RSv9bTv4UVZPhj7AJ54PzMrLtLVHCtrCcPY1fAvN6YTygFedANq1XGjof8Df
+tL8Ne+fSgRX2AvA5sd0ejrGi8bifI5aRc+RP7hUzoMZYpoRYpwi6hr55TovvUi2HLWtTDKXkrKS
GhbWE/WKK+3+WUysTBzNQUulTp7zoTJ94GSBQD0weimfo/vcgvJ3JKQBlAignpKMA6+m5XS+YtIv
3v6yLTjsGO7v8+yhjeuAHtoUNWun3WBcufBJf6bGojMJw7PJbL6YszPR9y9aZhoYtRODUVDHOlUW
vsLW6D2Ho8gJTddORI88eGQcXiOiWf+J6Ce+ZbwqySjpiLYof+aUPVLqHgcaeKjSn/PyphB3b7JW
wCE+ptzCJxxTmPCyxEGsHAgv+/U13xalAx6uKdVGGDtlCdjHF6gtmlw3R7wb301SJYRvFh2iKGFF
WDXSBhxQTN2b13XOO1PAPh6iz91wOGFKCRvai0Wkm3R4qi6lFsvxyuciGA1TyyWAlgaC3+Vtxkbg
zlTNAJAcznPa+FTbYqFPBVohnnAnAaxD45K+qnDyrhk4AFmspWFfsdFx+AX9Rrc4NGMHhQAKrQ+w
Gi/cv9DF0ZomXbyzEZNqIDlkibG33gtL/6sQkDHRivgkF1chB1gjsFTFPZEJY0+GKlgfjJbc1Mkr
lGkKBKrZq1HgfEbneH8cA1OigFwOYeBUxV39oniwSWzFnbQpw3wkzOXgfNNMOZO0jFx2A59ZhdP/
feGdhiuK7+Sehn9j892xF8owFEq4SR8yTwYCtnOS62vDz3Thtsl/01iZjJPDWMX+Es8337Pv1tuQ
QGB7g3fgaQ5bcweHOTfZtn+BqrwgHhz+l4cOyu2WCmGrPy+AvCD1l5TnNrsAOKix2Znr2qM54s//
8g5l6rR9BzTd2W4p0npiM/f4ziVMYT9MzNB0tHfbvtjzAb+NoVLtBuukBL1rMSRTZfeGczeHaTRB
wVZxP/5Dihs/9Y2F3SxB2O5YkPwQNQL2bb8JWAT7bXbPNHCXoetC/G8F1ZKHvNjWgeoqU8xHhN1+
/bJp566vnXx6qXhHcv932M9wXRtfB1Nvi+RdzzOeQTnq+T1531UuliOU+/GbsWoja8sF1Nn+j+s+
T5PAUwheO2Dd10kFuIfkj9ID4o47iSOb+uYrpe9rBohvSYFo0XOpscE+zuJNAvGwsF52O/pex05B
fLhRm+w5UHoM1RXsAYBI84naIyvZqHDz+LRu3u0qYB3dZMOnh9OhAWM96cqZgxtihBK0WB75DP8A
3POyl3oyt1ciuNF/BfyqEPXdTEvsgPcCB4TGFqW0pFwSxIWP4vUp194cb+X8dhJNy521meMFRM4h
cpIo/qX4XW4IC+uTgJ9yNUWWK8MDlhidmw3Vc/nL0dskPhV7Z+CaJ+/EWOXDwry2SsIYn3DddLSO
o4ZMbRYoSKcAmx02GVM5zvW4zKVFEyBphUPx2E230ajdUa7AErsQ3Mx6nEcxH10OCjrOa4Z6LtJq
kx42Scoqi1dil9RCQ5uUWb/eWQE/RFC9KssxrF+eLHSVvDPuiJ+KiHx66ybG12eK9vE2QY4B9uwv
pGSP8P23IhUNGhz2HrWmQo4EsLKrRvQmdvaL0rmKIuPexxzTbblh7oqcuKaVo0GXENv43ettJkJP
aIGC1PFPC0uDVwCXfI1DO7/PKoxvQBTPV+Vy969J2mSSJyxMS28Lrfck/APjTbDAlIt7faLZFVKW
xEq5/NrborWyBQVi8fCnu6lXmVsJprXY8SIDRYw/JsAq4WmzuY23NhATPKEuVu2YsYl4LzZtw8cw
k4Uu01AqBrpNX6aRtapgyRdmp2Ui0kOjpRma1czkFDU+kiK4KtRIF9gtHeI0GkyBxiOC5JXFJufi
5LXJm5IYG+j6FnK8b6Ks2cYtFG3xrUuejM9+YeOCLc5WmrgWYbIsnb7vAGFGeq1cKF9SLImoi6FQ
/+54k1ry6Vi0I5TGEBIl7H6a8ixxCcMR5QoWdGZfsaqmjAeygm1jz9GgWse+e8wFl44zssdRSiAH
2iqa+dE9UTk2lp4Nv9EjenRadfY1h4SWURx1aOmwOlgajpX1eEHqLvmcm0zmvGW4hzQtm+1DSt5q
4egc5Bx9OrFu+KxIY9xMrBxm2SRh/YOn/VkEsGSl1IhYOFGx7tSStlh4vpbtCItqEx3Ct8/prMM7
UQftdqFSDpPR5q3bVDhW68kaFr+oCDQTwCKawn1SamxZAOLEWg/2rbQoqdNO8hdr3XhXwrs0DJ+5
+/pBEkGuFuJVxPuu09Wq3pgHJc8p7ru61Rbg+03RH8TL4j4SItlFqcjJgUAlOJf3vWSue0INrCcV
3rT+ZYX6HVPSxCl1uxqA71Ur8FHDs8xiVlmXhbURCSXam1Dl26v0pwgGPZwHJiL5xYXlmlatrtT/
eUx+Mf549mhegqczxZhgrVtsP6mDGZMGRNS4rkx46T7kQdbArhNMh9wAGj3i0Zvp3Ep1TBU3HwqV
dWJlWAtjJu90gTMosDqWdlRoy/5Zh4Oxjm/ZvvoJt51VTeNGR5TI3fu5MDKiRzRakt2m4I1CnWpF
vVxXVe+NtiJvze6z4CESPQjZrDTVhPCLE9Pfyn9trn76psUhkj94BqYlRPsymKSD0vud0N7wNIhv
tJvVcf/2qITIMvo+qNoQyAWLkLaOzisDXAHU/n0NA2H66rdMszPCTSqCQV2BBUK4rR06sNKIh6xO
Oseqotma3QbI9J68mFddIP7PZHc7S9iu9fpIcj3PJvH5X9uEbngSyotzfR5QpPtIxkHy8jPLozu4
PkaDVYb2O/wIa+BKcu2GwJSau57JbsupM7QTl8GztcKkeTNvxLDRw55lf0agvglkZZG1Yvfj3DF8
dvHOa3lBQYjqDfvsBNbLBWpmdryWL6UU8366TK2YsKR/KVqVwJI8NsesZiWtzA/PkZtaYnbQhq/I
3Lb6KwCN2S++PG0pNNkA1pX6Ey6pdcQRm/acEsbD6ehfyrrf1id8GbJB2MxDYXVeflHhqDQ6JWcl
Lnb+jbZadRnERfCsjmhNAv9AxCAwkh4XIK/9hFiS6PMIrDr/gHg1OetkwoQFLPT8J6SbVxBMpj60
sghQFFqkcXxEul1RA5yQwaitNG24R88939wq3iclkGGicCmjDc9RZBHrZUPO0m7bj/+Hll4x5nXJ
9Ep+UmPlv8cSfEjEDjJLtZyXcVcelqaj3qotMpWlFYPsIYHZOWH/P3Ghscq4hBlihlud/UQuDAt4
eT5arEbIZQ/0JcqF4RGLEV0xjI8HFa+LEGA82LlzEjQsJGEVfNHeY8IX4t1r2GkdGDND6YALHL2n
qN0lUBCHUzridJK6+DczICPsbYiGysoSK2CvPwL4rRYhM9FvZXAWoUgXmvbk3GyIDqNvMauGpXtj
l+Q5WSl7zt+qD6hZGeVLQ+b7S7OTi+mT7pdChQz34daWEuHgqQpPCsSL4EaToc7FpPaesC4hygCD
iac70DnkdAYsTunFLRXfJKbALHvY2Wlvfu6wQM7e8V0oKO/DmGl3549eLocOv9oplkODCHgJzz6p
yUG02YhRXSH1xckcaH17Zozv7AcXO6q9e39j/J4eKqLEbHI8tI+px5tX5qG9bk0utIncGNrTOAbt
kgAMI58TQK572yKrPD5FxhPrWPEVmDth170Aza6F1aJyy0x26rbO466fU6latuBPb3mrxy2J23EB
nw0L3HhA/fl045hVs/jJPHYVZj+zK8qR0i2XaxU+/uD9Pyz2bRFX8sqdgu1Pwd0CM2Np3dRVc8mj
95UegG/m1EDL98oQQnsSTjao1Ym3ff8cKzBfxP2+YcENVBbkM5gTQOFoTh5SWGzPqt8VcQrLVcbE
IJ4fZgNaiXk9qvNOvVymfVHG1RXyEbexfvDwaqJpXLiUt5tNjI5JmdAmwEPLAJ56dRiZDXgLp926
ZTaX3cxOu1VJTu2Nynn1xhHdSh+Yw2H05aalLsbrvsvWIQHo5EYnO1iLIt5IhpBNZUGndDS1HJwG
/7eE3DDz3Bz4TENNbl5m+qMTMS6NgLgoLthQ2Q9RvioCEKIY38wfnX0eS5yQ/AxgyGS5NXo+nI+N
IZg+DnMRIF8XOgiwEjTJbXXEwdJhPxF0qmQX4XLr5oQp44x/fEFK2yY3wUw07U13+nXSJUE5r2zl
j5dh9rvYZ4VHcNQW2/9/K5dH63wQMw0lapY2LZKnvIofU7HVS1fuSbgXNO26Ss1YFyqKT8AFpQvz
O+6uZNMJn9zG40HSenSxC9u8JllRPDXN42kWePL5j7jqbe5Pfji889LeZSNYR2lWw1Dgu48buat3
L0NI9WZpm6EELYZnSPlrPEfjmCOgjaZgH87hDqgFywyy2ezjb2/1QoK5dHNJfQCzT+4xcI9aW+TI
py1wQNm0Re+YY67lYvxAJcpp6dmue1aKUig4oDhbOebebjxidzNXB1p0CUrJePxoorShZ/0syh1j
rMZhTrwZLhseizkvtQNZHT+zxNKegkQCofV2l7l5K3aczCfmEn3l/sgVvv0w8GXVLRxFwnPZLYGX
q0NNygWUK42qJ5YHco+KW88mUXQPfTV4nm9gC3b7k3YX45arN1xns5S7H6HnuvxlLEvVneKskiNw
fkoMDAezkm7lPeYtALzWdL+isTB4m7wLOkg7nXURnVQjvYmM1M3BMSZq6AeOHJFHApeLdC06yhYH
g8dJnIDzhriG4xW5Gso0h1Gh8/9GyZvn4ehAxcFdcO2KBzkZVH5+eG4vQOKc/heDIhMuPzXU6cQb
RLV38jGC7NwDA7QsDLo+k6/Vw3i0jdYgNs3EDoXjzB0H0X2AMrnQosGxmSLGkGgL7Ov7p+ui6I/a
fzuqR0S/xQIaNxHPsE6ay2ejFyF6LF8uxvk8DTrK38qPSsQUXlTf3yRbk4PnErkq5QR8X/f2pFBb
nuS8uPG4w137oBscOj70YNVgWvnHzVd72m586LIt8KvKu/1pBKaWZuYVBZv8Zwj3Mf62E8kSlA8c
b1UVR5sVa+ZWERtiYokD1UR6o8CfJZZrvfDRaazFxOFbbqZnTI9R00Z/ywQiJVafKq1eht9dFdnj
DYnT29u67RSgU37+8V2/prWXmmwhCep4uY2iHTcGBJugfAGmMt7zf53NuXS2s0KUfAD4LJrridBm
Rz6ZxvtA1N/+eBbnF+cuEZdIhSsBGdiEHnguGoRVQtOUhHBcLRODmGNvbelze7oSVbO30GY28KNJ
3HsEyc87Na3ywZgD7QuaiPJpuusW0MMRNI/lS+wD1aoNde6Zec+iJrCTxxh6tILAfapEQZPwRC9a
8Ou4OXliPyPyT7MnRqNal4UhentMW8khPYjJGMQFaZwjCJQastd3Xkx+ELdlYsYDp/yKNEfqEf4P
+JQlBPf6KnXckzgy8ktgUSWSYIomJM4UXPTJwMp/4vrqoZxc5JAgX9Vi3DTppKKsoCgTZUDPAlw7
nF3fESWeeGSb/7sk0Kq+wF8DPhOeLsBF0rdSrKLJvweWwf1wae6MQaoaIHXV1lOuUKVFrLOgKV0K
FiE4IdX0M8LCuutiSMPcn5eo+VrZ4oiJIZWLY0BTQHB7p+AjCFBowTkxtcLxAamIdVkQ1Y9y/aQO
ixqvTjUG71BtoNG35gPMEaGPPuottFBaCg1gZPjjHheO4m5aUnQd24jnJqRUoSLDHMyPY3Ro5i5a
OlASCJyly3xYNyu4aWe65CuDhzYc3HeOoXQmO69YtVGrqP78CD7tW5SviCydNkp7C+JK5rdjZIyu
SsDWguH0l/c6Jba9hLi08WFp1SidmH3Axk4pEnpmCf1mqIySK3HxG8tNdbbLUAnq29x66ERlX+kW
nui7w0+nzJhKLIHn/DJDwtYJsrRHH4smpvl10G6+FrVe80iEuoHqQvpcRvS9PFt88gMSSCMDoTNt
ifFejv6jUAiEAAhSCW7IEGLaq3kO8RrE6MuA2y0jT2RzeMQeiXuYW9HTfzkaTGeTRZXf3YvXATfU
HPxQ1fuBO5E9e0XHkvuD2Ke2y7oynG5JzlNdAGVLuIKpMfAt69o/oh/p2oTH5o+WD8meTfd0dzJ4
BuETOG/Y0wBTIJA2CO7JCAxikMnZedABmZ6Jq5BRVQ6ZgVsQ0fTO1iD3IWR2HYazp9Zi0n3Kq33F
2NwL8ecFplNQ0+Sq1LiScZJUBdN/mE9VmNe638avtSyvWi5vBvBKamd5+5CuIrvvqgJ29gmS9Qj5
XBxIEMkkOPjhUKFeTqY7WmRJ7bU3wNsx4zXr7CzcnQOQ/EhNyIk0l5cY+6xc/9X5JXSmZuzpyFvm
cfYZPfIiYnNEP46tbUJk+R8AYjcqDioamUo0f+/yj0S6jR9g3u6TouOR9S+DDr781CarABj7OGP/
O7K4HDnbI3ZfEHMbIPsG+BatkJdqhmvHE/MqvBh4pcqOI+Iugyp3nNWBftUnKn7K2ovE6NfTDhO0
NP63Zu2MWDpwm4n6POhBOHf3R2JVHfiuYDouPBzxdoUuLnD7anfSm3PIAnIrn7HLVrFdlXgHArEI
QZGhGOME3sZvN849cneSF0Z9ENuGHkTTfyx9b38dlVoBQQ6ly5KMPCJm6hM1yvTYYGN1GR0IDR/0
RQ3tdUQITlztRLkvfLsr2YMuauI5pqGUsWZWDwy7ssXtdKikYgl8JzpgUZQEQvEUQ/N/L5zSrr1x
IXSwckiyOTxQxOUYphre4f1zTp+TNvkKCDrafacRQ9MvlipS9PPfaakdpbjoMtQ7T2/wPXBlH8Tf
SN1K8bkeOjYJdU9YyzHfarE6JfaNuVOJtjvsimk34NnmTCiVWGn8xHyla2aZHQ/8ANKN36d8SqXt
XpVJtRHRC7tzfmmlxXls0osdvUJcLNpn1XRjDu9mgChez7kkoR/4aS6da5znfhMRe2PZnl7Gdum7
oqTDBVcok0TRQcKReElN5VqMso2cUDYRuFfAToi+FxSUq5m+Q9pxTgE7xSsDc8pIV7dwtJUDx5sc
7Qf5Hay8wDSKXGUIE+fSKiGU6OIB/WXl+d1Bd+YuKEwUrObRDwjuBLyMMLgNSe3R1psXeElOhDY6
bzS4XSDzQEvhkUUlv1956rvasNzoyL1oiDVLLjSPEZGsNjfs4Q2eX43mr9Cit8WCuvZEqsR0rSe8
Sm0D8j2fISm7hGWlQZMBDMTjsVmkSRTBnRTpcdOgWGpRLo/pmsuDBzDx67gRtOmGoCyY8o7T8Sj8
Q0TrEU8wFfSCF8ZWisclxRCYk9dpMCQOnZFdGZh6lqI5ehJvdly4C5FZuo9FUBIORN3yHc0zisYK
vhkvAbHNBjGdC/VY0sbPrH2hymHexoufCJrH2OA6X4zmvtb63U68Zv8OyMPRpk89cEBKh1VcyBqd
BBOtpcn/NKk7Jfs605irlBkgjyiQRoD/uj3+rDwK7JBSJmjF0NztFrS9mImkdeOLydaPVPaVCJF1
9aEh0/8EE47SxSwBYUCV2IollH5hXE5tTxtCD5xeiR7naMLmMUy+EhHN7HcsjfJHFI01IU5vR+6q
izrrhj4haDKh9r/mF1nql9Nx5wyQSRLMEWq5fs2A52TspPzECsjLHmItINV6xU8dF8TB7DEBQjQD
NWpiVFmhPpW7gQQsC1VdktvbCbvGOpEI5PETp8zTgMzO6dOqRmc3pP8iueIHfAd2ahRxtq2GXYao
+Dgu+kHuk0t0qwVPhUeOyAUgZ8zZCDHMplsslWxGadScm39Cx6gArVwsxHkN7tuQHdISXuX3RdFc
OQ2E1qb20IMCokEjJJfdoHgVURJFJYmJT6xmfaVwJbksjR8Xq+PE+drRI15FP1ZMNqr123hdGKE6
6NClmPg2Hmw2YqJxWfpgBdexJADI7eDtcP3QCJYpFSFAehpxr0C9HxAZtDZRyq2bwTSJwFXRZMgv
Z3gI7po2JZxV/Uwf+jqKOl5GT+griDDbY4u+7ptE5Jmuv8eYn+zm0BWadqg58Isss7P3X/aeAq64
1XxxlQYJQXs3A/EWptYdNupe4eaRjqKwVY0/Csp3boZNH9P3bdJvrq5VgtsmmUdmdvP0YVXBI1Cr
UEwEASuTnMoIAO/lJNeeD9h11foYg18KQ8efF4mrIRa79oFuxrFpHDThq2kdvQ5ei0LJjlUfv64z
NF9+9tIZhkcOJQwmBgPrR1sMYHB7Oi58b7Hly/dStbul6EwKxGSgkJwPv37yRUUGwxHsxT8rlXAJ
E19X6D5FYAhU+a7qrD0fek7nJkJ84t0K90m5bH+nG3Wy3HOQQYQVSeT3BpN4Lo8D+os9z8rZkC3o
TNDkEEuoK/zhl1KyPBDu0u6MG5oQsQgJcnwQ5Jjnt+VCUnIjej8SE8A9Xf4tdp/eKT3onFgWkn+v
fx7pHGImwEywBAmabu8ChMVCxEfHE84fyLl4TxNGDn4fT/c2NtAhjWG7rL8dUzusCWhjFTKVqyVs
konKak92o8O1rjqr0/Bmn630pxghTJY7Aoacn0UCJLZETBpTQsNTqDzvOrqjm9ZMc4r2K1/9VcyQ
epXvj/0m4sL3bI4vd9BrgsASRIXIASKenJMxSzlyMuzlmDA66LldjlBglxBAL6Ou5i73ZOa3mP42
k38hLXGd2zx2pDilr9U163rsyglRe6UoWGZA6+gg5lJlrH/euSm2BJer0q6Od+O1y48fiQvy8BqG
sE/gIw5vAuZgDNA7HiNgsg2Wum7ytQqLTpRe5YV5KcfFjM2tnpspM+XUJtq7rGUIUdH2pDFs0h4A
x8Qk4i6XbC8IGPd1cvKkdQxe+daUJFKedA0GVo2BaRewRMcNgWN6QkakrEtlliOauiiUEbqlRPJY
kE/5bf/mxilhyMcYx8/9c/DeWWLBTtF5rehc0ifVJdyftaV/Lm/9vFaASntKSoodx3xIVgJHrpm0
HFhr4X5Aqp1hN6rXwbPbfLUcrkWNg2nN5byKxsPi843OJgsL2lp+77iJavlErmquGFsImQM2Vl4A
amk6ehjU7OUA62tHPH/Jp1H8NvnydExrx+Z6PZiAO9m+X+O+M6XLgl6ZC1OqxuJxEOfeEFWoYDdm
qFNJpuS1zpd4bIl91nKYGyHPUPyg4PbfD0cTzRlpvCRY9H4FjwmO2IlAXhaAZ1EnNaPqbGXXSD6r
uCivIka10k4CwX98QpERxE7zKVm7h01FC78pZZQN2plx8V00cxX8+TaMxSAPwhO8CGXRv1ptDqFj
xndejLeIe6l2OmLnoR2Fp5D9noq1QErU/HTKhTGXZASZyHhPuzVqb3KctDeCweUk94w1eo0/UOSj
AwTL0SBh0P1WMZESTA3WOPXGDXNtHYr+YG8+Orz1+SRNMe35V34dVDFVYnnDahIcz+pGur8Lwy1w
yoRNztCHIUuGpI+WsDIU+90KFCzOa76Pu9Zt9pboUK+SUX0K/c1ucj2juIWZqe86FupCh8QZ8kd8
8Vhg52ToVg+cB73V+TOBK5+n4/XJHnGNUzBvWwWYmwTuoIiMElJa4q+70kJXFxR/IQ5d+b6NtK0M
oKNp1X3CWjIW2tn66XmYq7m0K9S/RyE9vpTJSNTSHQrUQwINBN7ATQO2/rcImpRGVWuwozGSrFNd
jr0umc4TVTo+vrrZYEtBzB99co99kzmp90YQ3I78wGQ60UJbtzno6AKlCNmwEP5bcfPhi24ybHI4
lffqHh0vEistvDS1w3g/EfaRq+AeUFzNM0c+hWRjXHIXcO1XBeQKjAYvDxxa2pebhu7T9KWEYC6R
QovIqWC4Ffb9j2HW1FR6p5Guzf60XlvzsWMBXXiayePATB7YYVdmPS8hkd80qhnSoSSTuEaC+ox5
L7pp9TL5dKJfwhALsNeEaCETXz2ly/XLlQZ+3UcEhi9vs9MUzMcltQ7zF1sd4BJuN6PQytleJ/ml
216x8I5hPwgscwfLcLv1QFk9SvxyAiVo89qKkD9CSoM67BbLtO3gRjEvw/qXKYS2ll+vBj8uWSvA
mVvoTvuFSG7/oyho2NOc2m9RaFjDq3n3V5z3OXewfb6MAOT/fDkl3cughYvu8UP4rYEXQCW/ZTQc
MtDlu6u1SYk5/uQofuhsnkMs6oW3eTVzjGejdLi+aq/gWdBm8VNE4bL2TUb5dy9ttZx7oOuIuTwA
Hr7QMom3aAvyw40N2//+i8gCWkipHX5YV8mfks7O6n0iceoL9fjqXMLTRPDGK7XV2ZvSZOIQ2xnQ
z7sKbG6bWHQ0g3NrfoaZWo6bJQIJJB3755trNCjJGbIGEDeu7bNCU860cH9GLcR9fBfljJ89UNpM
afrTTrvIsyTgZXqdSnRdPvGQb2abUUiVSv4/VJJyoIEpGpweVBc6x0sHXVBJbfp0FSKYtMOF9FmY
pGp/gmbGK5lZIDhGNtKGfhaK3Sxa4oFh5tdA4jgXXt7fHPGsTmz1MoQ95R/6tFu5WLmbPQFugjGH
UGUzYS8y7g/YtrwxIlL+wj8r+lDIqzVdijmp95WxqqHPtX/KUp+XIUg2aX0ElmD7Y+UKh91ZeODO
yiqHZ0MLgXcaUlNjP9zhtA5wxx1+VeUhwK49MtiH2SvEzK7sPIO8GG4zdmk+t3+pFvkg8f+Qoh1I
wWISbelPTyP9LV/2AeiQ7GR0tOvD6wqCpupX736/ztKH6NF4SjSC2/y+bqNufkKMJTVapDT+djWh
FqoIv/i6+fz1+SDCrFVqqEf5yXN0LlUPysnsR3v7ECYYJYpSoSwQ3KB/XG/UjkIdY8VdFpaeq3Gv
n7svyusLO7TpTOghSbfTi0LtIjMxV7NiOXNpA2qgjBDE7VzDj8ViqGTqk6oU+ClvHvf4uXyFgT27
LKC4L7Q0VAybDIhGRRwc0x26uWOeYr3eQTB6TRUNwfQmC0jYUyPKu2yKJhe9aob7+GxCpmBIesHZ
l/aPzZ528ZvIb3Ju/OF4AG0c38yl63hfCk0QChIWHjlYpbQCqzx3oED0zhdE5HZugziOxGEjcMwF
o1HmNLnoe8ZA7p7EWWDdYoGke46kTJnbMrL4yMRwTDQWwfenmXfjyMD5TVPVfPV6GSD6TuDZp3mE
ajcxW3Cvh8+ZSsTcU0hc3y9PdV7zKqK+gKGf4nRS1xqrVbQ0jcSUgDtbm3WZlnKQPTUcZ6n3ff02
C1kmIB0KgyVZ5bEjELQkGB/p1PCq0iP4GmpTw9OFYxJx8Zf8lJD0ga0yDIo+jLOdADYJoT5OI8zu
+esIYYwKJ731JWk3v4ebx1lNp0tRRctJdEJnLWPMMldE+eGQfzvd41nWLyXbyDhVFHsa06H458rt
z5MUdBlws5dvwCaD/wRIxVNs5REj2Q0dpVebRZaqZIkDptcQ/x6YMo8aEaGKRAcbi5ArW0RJZe0r
GBYGmiTToPKqieA3lhLGSjqtwCGbZclDsI+rzfXaynbOvxHuZ9lvgQyvX+FYV4IJX2vJCHOkLj/i
mXm5hDiOUcDOz+exejqw5uJVDpH5MZ4RGp4PKWO0aqKnHCO5wSBq431HcIEMJWo0Pk/IyU5wcrBK
HfI4vcwbL/ye2+jqN1zHO4gYym7d7+2+EAUnl+FLd2ueKD04ufnJaCzoRqNpAdhQy2F1rbg2SZE+
xXwdyvVOa6vq4y1cFQ6198079rJyUAln9dw0hRO87n5fNNzeouqHKj3Fm4s/LArj76oCJzZEpbtN
PnjEENs6MDPQBIXTIRxHApwpeoatRvFwLEJWRPUGHsf1XKUU6UAfsZ3PrvbJwb/PcIDFG2hpR4mi
LMHtJ/mjYQzqrot6IaWyK4eC3IlfFNt0gYcypQpgIhQdBVhLALDBmsa6m32BiFkn8wzrFFK+YWSK
Pqb2jEW+EGRIpB24DH4mFqowSWNL0bWqZT7QuCjLTfNsCJDjzagWsBqUKxnwV3q5bakVwhRj0CqT
v2w+Ss8EcTrN9vUvfu6QTl0vI4Ofo3ek1NCF8WBgMa43TRat+2DS2UhfAcztY5SMle3Qxh7WFIhP
jb4WpghNomv14/NFfTCgmf43DkdVtgqDnODC5W8+xuvdf7DMbFWHNSMJ1XIKbwX3KsTphi6fqg3X
zxwqzF2XniTR9Dl5qu3ADLvjY2WCdSWp3h+G04w3JczCKXElmcEQ2K5024bbY0hSqgP+wFMD6rE2
amNcs4133Jcl858zxVgNl8SbHRmfdx96gXZNie72dtDWkXwUBob3XjQYGOi9CHJItyEXsL3tVjUz
EGEh+EwEOXSaM/ZKUof/0i9YylRItelp2/m4anbmQMCVxWVw2y/htoq3X0l9XMsAouibTnhTzKdC
tUEn+UH07/W+p43sunvy0E1VynBgE5tpAGk6Y6UrOnkNiz/IXwcFNbjK/4fNXb5BEecUuKwfxuNb
qxZ83/w9MaJ7tS+sYshsJNkWP4K/noS5R85uZzOd/3hvECSM/54YmECAWIehEEw0gSh0Cpsmj0n5
Y5pO4AhzLrFidYTGDuQtzqmCuG3sTW8BG2R/P+iM63lH9LdQqNYUqr0PX91tqSm/gwqhrlkuSbcV
yUveBi6Lna0kewkzCJUlgGxgYovLDWgqNXcvVfAC+8Dn6sjVr3hBXZotLXdAj7W6JappLl4W3mIS
xI+MYR10wgKa1Glyy7Nz15iqURwux5O+ZhFZ5OObFzzd0X9faCf7N9/c/njS6yuuDWtoGlSK4a0v
rPrSTce++PXu7hDvuvS5auGaneknXUa9PcXIj/g5p8jnzCHtOjuxMzc4kifMw1Jx3gyUzzUNOEIt
Amuz2w2+27T0Ggb0SUuRDWR6YePVgwaJFsejtg0ZVfyLpDKaQd4V4ohZ8+yQczH1O9rUyLai1nuy
gZwvmQbkejxZdLJNqBbZeR9ao/4ILSnbm/Y3BFs/fMTmrA4oRn1prdlYpwIRCvlavXGMKB6NpLJj
vEt3ZjsoTo3ntDBRzTSMkhMS8E83ZFEPUf1PVmm3MZIWW6CAg7TCn4jxpkJfU+oJWXrH1xC8qyVm
n3+sJ6lJ4yYRl5dMJ9BHuujO47LiZjmQyQ8v5IMDyGMzh5cYdcC6s1AkwKKklbq8Odqa5lBK5tRv
/WgzwX/G+P+j24CwYMMooRLdROY+1gSC/zzSIAd+76XKhg4yAcdtLHKM9VMwcuPaHyDoUyLkvLc/
CAwfBNBPIhEQhoRqEQ128++m5kLgztYv3L9U5+He1cpNxGmXmuyG3j1GcKTJdU4zuygAn52KYODA
A14UzbAQpeDoJtkG9g6v+s1zoeUWk1CyyaRHPeRvnTc4Pbpc4W2I+118gYMmkhpMXbti6IPxPpRY
PsWR4+rxOkjhdwYW6AZTAk9tt1bIfLmCoXcvT2aOmRKtBQBD1WIsaTeqF0UnzJScT/EVXgpLjxGS
/65l+aaJKqNYAifaEmYylZ29Mr3DFltcn8iiX2lw7+kCxoBNJWQ6thkoqjaQZ1zvYn38ZHuFO9ef
+aL60GlEYaz0eMlTvsq5na9g9MLNDKDIyzW444PpRZS8DL5tPxQX0LGqmTm8JCwEyEf4aM4fPzix
rUDTQdiKBpmY96amyOv1W1oc1zkUXVTWT/XA698lThstpctQjGR7tCCspDel2AjkE1Ve8KQbsA3u
q731hufMlSpVfzV+8encQ1ytHAmelMjx6GZcHlELfptG3LNzmBP8P+dfPWnRIZAkkdkZbhaCR0/l
bMhIrh3mOTf5JxPxBDJFrXLHo6DuS9eCMxtRlu0wE1KTMdBKvoKK0mwINlNV4ewFKCLQ7tX3EhYJ
CedvqCDi4mHHlOFdCbE8MFG1qn7pM7kthb2moK6mOfYmoVQFhhvA6g8Tx4vSeTGMU507Kld2Ab1x
qUXTx7sBWLkK4963Rv0RXmy/U1MIzULLrvZGES36Ihzx6t8NXVH/hatehUGPWyhK7RtFcmkcnpZI
85zsv6Jx2MRjO4UwQ0Edt0bHkj1pWH82u44HoA+w6f/66tPmuWK76Ls0xr0G8FJ63Y15kjz7p7E8
i+3rvjTxtgAvLgWTn/nm3Mi5rriLYExYo+r9kf4N/HQQR6NTbEh6x6uG81KFIpIqhar5C/qXzwCp
nsalNTRZcsnDpk62snVh4H8DrMjcr/xsfR20J6YR9TtmlexFBBV9TcLa1OlYBeQrmN5tqxURpcee
g/k30WwBNnAYFU2DsT9tXcM0DShTZMtJsFiwnOzWZI1Pe2qXmxRsdZ80+7S2LVaWhTQVF25aezf0
v+1foRbbRfA/IVcALRQODMJTXLxOK6/C3xx64BwwUAe+GCm7hYdDR9CNJxRPT4AarqZcvGZ59S0m
LnYDd63jXtzAfl3+8hk42pzbbb9WJ9UdfDHyBclHgc8t4h5ntuFOi0NiOFIcWoc5ubAfswbop/hI
QZqXLNuza1YmNAXYxfn18cD1tAJVItdl8ahxEhKtS7+8sJ95/UThYEGxHz+oEfR91UKm4zL69Ci1
gvOXS1zdGOpLF+8JSanubENMGL4sbvEkfQ9eCpmntE6+zgvQyzIfY3mONbjkMiGgebrcERO2O++1
iEZ5zPeVC+YBJjDIinxWVI3dD2wzJRhBwJ31Gb+2LxVN35dF/tnYkPaXNVz0jhrH6XHHPX89QAn/
8Ytc0jc8KXaEWILZWEvbVIER3nNnynsy/FGUV8gCa7ruETDNRqYCYJ1lGRuw2BR5cC9QHq0bhCfO
UdY4RR7LeJZg7gUOmtMUyR+VKHn77MhAV84W5lo9KBHutxTU5iKs2fFabfjf5Qhet/vcdtHT1FIF
Ljju6I84Srm2mlkrGQZXDweZq2ICdQr5KWDCGrnq2KV7xjicM2wTda9B7Ta6UZTc4gSYqtlXbQr1
1fV0l63T7MQkKf9CY58yP/0sE3R6KNywXOPc98QYyLaZXFEIcGt9CF8uiy8e20TYYfwwhqTD9XAk
fz2+8lW4zvTPRXfn9z4R7sfqplYYBfvFtYYTBX2omP3eARXQEphOhdC8BAEq4XN2A0bMss5SEPha
JRk9mttTiworEqTAiDo/IEJyLUQ2EWBWG9ADMjvWsXSZXxkg1jQL3aHKtkVZCG17e2kpbroCq+jH
2BWoHUPWleYb0TiWSN+6IQs+AfLDY1VkyU4Rr8KS+tB0ug5tredd+y3sLDGeXyNGI4H67y9sAFhT
Muw0HDXMgzK8XsSeCqtKc5JCJsEUq7+GzkUDl5sX7RZ760EakJN36ynprJMossh25E+7UTSRklXJ
YB9mu1OLlaqA6P44DmC1nPJEkNyCVZPmVgAzxAeHb/NkWq1gsdFRd/LcFoLE0MmUlOrkfEeocB/Q
mymKLN/EHsFh1lLnTgDG5DVg2dKvPbKvtQsQvDwQGXjnl9eKb/IgLwNf5WFRDqLmtOMRbWr1B6dD
Psdk/g2v2yYIZKP6Ezd3t0y46ZYlVOR/I25wUQtsnFJtBPfJ00J+XQuxiOHF8zNjlmJvUotVAmCw
Lr0xtjwvlIyduHVDVNkmACEsuPWqCs9fs1Kte9HUIx3YZ9YXZiIRR0sbPA+JrYwrdhvAumXLgySX
lrmKx4QQfGIJ9bdYONU97sZC3rF56k5gb9ejqhrtZbTBLWFpofWbkkYJbSdjwGW9kNJqd6+13Wk5
vFAoIhD2R04j7WVQHM3ENiYehL4WcvGm+ZFdnfUpkV5iRSLXI9buDIdyFrTobLw5G1AmeWDBGJxw
FVMONDcghdRtLmq8QwDFXViKqww6l3uLjNhoB0RdnWqzvk2viY6Tg97+ETAdI/WtyCVt6VoXo5Xh
sjAZIXQTn3EvtK3LiGDHK9F1Hw8d5RHsvV3nmsqYKDBsr+dWktcC4uQ9tazcOJP93757Wf2Efc/r
ZPyBlrhTg3v2JxzvIsdxmZg+l5fD8faXTOQAE5ykXUXR8mxwRVz0kpvjdOWEG9fk3EeHDKABPile
FRG+SZjM8Iwclo8IjiE626tppO/P9s2vYKhN2zVaP+jMATWL5Vnc86rcwnFbo35xBf1rp8ISKsuE
+FdkeGXKPx6a4neJ5stq28gWn749xibsJFO8bPtHA2+ogSVmpHCColHOQ2vHgCYgQxozAXtVn8mH
Ty/SpLoRdu9aXYAI9McAZ8sPVjsbe962O931nU0EnqZdAygrkDJ6Jn5JdMmATBLTezCuy8sHxCid
+Rv5BHmJCqWCG6TXYptjxDaTVIlRyQNFvgosKzibVdnQvHps255xCCLG9tdc5UMGMyQ4R6yg3HwA
2mucr2560N4mXzPzsBLsgZ2BvTpkkHLJ7v+Rx3uSisk899cjNNFf8pJJYnN6m2rrA7qKFkYsqbQ8
zd18y9tDHntE+f95EGV1WyPRb/fCofa89nlchs9GFm4jIVN9FIZoZ/Iz+JZzDPWs6/q1O/32WItR
45yxbDjUZtPIiA+kRudYHjG2tbt05OKWUrEG4McNCVpX3brCK6/Mr3Z7UdO+luL8oiLdlknvfbvL
LwzPHmj5I81t06J+/OhXsxsP5lS5xjhB3g5djNy9ySS5OI1wSv2+AnSP7Ps0VM9JrPtZsuFh+5sc
ovzEaSTJcWPujCFohLLTg/1QuqdPDEHUH41L0MC+q/lZ7I0JkIH9y8P7yCb6CFvUrsuMNNEOt9+e
RUPOj8zIYIV9eNojDJYE3U9JMFeli7qFoKACIKzUhslbjW79Sc8/bVd8bG2zdqhuFX8rrZmW7Bla
C/3FD6whHEuSS1DaAmDZLU4leng0PMk+PgIGKgVfrevJZG1kvRZ+74gvbM0WuOR7hJnAkBdhwiyR
fyZVYZibc6JlZx4KyOpHGKpEcMdWwFeOWCc6usY4PDMAqBGuP6lM55Bh3/xO/Yb2c9cTqp9IXjw0
AwECGnFGte7egpmBVH/tI5/Aeocxr19HC79ntmKUQCKZwdiS2njSXRpr3ltYbXiu+OvMKX4Cwmd1
71R25t8hYdRoaDMRooJpXSb8Iz9exEPA/ty98D4H1jCH4tw4rQoi2ozUnLRGbD7iwcP2AiYEllpU
3mAa+YibLkEfTzhV+bWbo30toZQD94+neCtkE7QEyABm26wqIRxdcLjztn1luN+ccQ5GZRojSAyr
LFy8ff/gNJgDpeY6etXi8I7WrLp71KlX8pyPktcO8HCFwTBQCeLpZiQgeQXstmrQz95+0gvjUXQ2
veMHmrWzzaOVtEB4mxC2Rs+UFKZNaPxTIvFFgv1UfrkWAsMGrtMtVS815pHMWQvdoqgY/5IEePA5
Zf4bL1fnWX/3JQN1Q9IcLsvKF1RXKlWOZ2YIjXRaSQ+J/55ShN19R/yRocCYi82TnoWRdktQadyQ
cK5eL+o3rhrImcBJT+NUFagOQQrQTjWse4PMUrYeJkzT6ZwJHzyfw8AcOsUst6voaJBnGjyTis3m
gzAEjQ/5kU9OHXL/tLPqE2oirdTHA30MqkPFy0i3b4TCkKiiYB8wMiAasJvnZenHjb18VrOqT8nf
sTV3MET8T2gy89mAwvGmwwAg5dYi29QqakyNXUfhiUDcYThv4T2J2TdUsKDBZ+Mi4pHuRsHo+8/b
8NPQC6H7Livif5RYpAJnZRpQr2Q0WswaD10oFN/ppgXYlwdKI2sDE50RLhiAGqFTZhcjLeHDHBC8
dQ0SDdtjnJ4wh0pgl6fQ7io/2NXDWUQq8FxFTlXqfZXn/L+3nL8Wfs/Wy9kICxpjdDRlAohGvoqY
GsUJABiqgFR5kpmXjtTLZWuo863gdA/+VSgNmeQjrEViSYs9p82LriDeGSs8SgvHg/TeY8nUnjoK
qwlt8XNpsnjv3uSMaaTl1J1ybiW0LTgV0F2gH3Mm4cDJTP39zrjcvBsvd6or+VPfmkuT/8Wum6Cj
wEH/6/hiJurRwFyu9ab95E823xWTPnz4Gkdw8z1qE3w5SX94iIsowea/S88KkDasZq1HIEEpj/Qa
sepalbKw6FTMTUXawBmeyGbKlDfR4RskC14EitcswXdhr+8V8ShdWrwYvpdeC8PVhVkfVIYFic1A
h1u0q93awF6FHP7eKdQmakfXXMkhcYEW24agMyWxbp+5OsnxqC1FVhZ/c6SoDSF8i9UaazJIW4mY
JtHkI1cV0kiVMOC96daJDN599h1aHZhpY7jEcA6sUelWnDb2N/a6mRdgCvzrbXa/dhKxjuxYCEF8
vjTn4SYJ9DR0OY8irBJZy+YbHQf60nu3rQ0UAMdEmIjubrTBmOU1d09RWaBs+n148lmRe7jLvsCv
nVEZgqPrEak3CKBhW4jTIjdiTNmEeIm0seIE4uKKZiT1mvK7CRabi09LVVdv9B+xhBe8TT4Wd+R1
3eTWYvfQy+of7iB/ZzcNShYAt0alaEqEBoLop4EM5LDM0li8EHwLJZNcGAj74pX+dm4ZTMXIAGHX
yqoU2fASuc737EL16GMH2NILJDiVldr/0dHJOcyrMAqu5IdweNyn+GUddTWHfLb13937WGKnI83T
VjRf2NPcF8/udhq9bilErPEABM4QFKP/V/8YSe365y0F3Ftq3N1HNHgMs/oBgxyb9Jjnf9FRGQRq
GISwqiMk8sfU3pQD/cUzaTplEKdY37DHnRLHCGqXjat6nVm4LSTb5YgKJmP8/J9UIZ5JP9kpNesS
tEtsV8uLgWtSyjn0QfA8xV5VizwsdL4vXg6p6i6EPY5KoBGHkJkER/g485inioP0amtzE8ma9TBh
OIlv3RH/BeemzNtn0cfP8D8gGjjMK8U2qlpSx52j2X72GVQr/VipUgnp6p811PtoAMDvLee7qod6
xSX2Pjad45W1XdInu42TnFmw5veUk9AqgWV+WHznrO13vI1jKh6/iHmJA2urLxSR17JIWU2QnqWx
nb+XR+JqCwSfZx8eSXZmrOJsNSsiTJjoWxdD3TaVznJmIOPrAT8J8V4kTvNboYYaZmSjgCvKPWGs
FociWfPR2NL/qxn6QJoqU/3m3hIOjuucDXPIMp3mNm/ls0n4x+45zuQVhJpunh/Gq37nIEHyH7UO
+mPfYJyt8OA7W0gfEKU7pUPS1AtcsxlwVA76BaYcVWwApA6Qh8MA9dC3SWnC/rB94gPETJzipLbt
9VUj6XRA4vhpzyU1tbK9r28+Yop9yO+n8zc+/P0Uegq2xvBf9TeadhVYVk4YsGVwVTXzmT+ErUSi
qgJIKzerrpavaHhRDd32m2JlgChecG4q8kCqIwNVoZOMR+E/GvY0u9m+CTmFrkwf6EP5lH3zDYiV
lYNe2OfrJl/0wgnX3RHoaMrNme1/LRlMkxZ8iOe4+gAlhEpzAwaXpIXv6TLE3Z6KjCEPLXwdFbh/
xrROkUUd2AjItusYqN4tED/munTPWpAgEtqcr9W1XpUChdZjRU1vApgFK48JZGQWi43TYtiykYwn
y1NNCgfdQFt1rdaum8tOSvmeNrOBn6kr91mU+pespR/xbKxShoaei5VnccU+aPkm8Hv2yCjmJxHq
mylkkOl8qwoBg1/QP5dOCfbVqYou6nYy0HSUQXtd2iKZX6uol5pqoMHC41IVuMCX8w+TU4m3qNJa
PwWri4RUSOuR31QkWv2O6g6GG5lJbzVuUQAdVTjORXqke71fzsrmo2VjQ0sa2tDZTBBywajvLoLq
FQKkeoQ8q0r6UuNw963k0ChhTif13p9LENyiCb5H6WPOf4pYA0WTYyaHVoLLAOV4E5qE93aV1JOs
9TOg0z6Z7v+gcEq/uNMEhi55egQtlvESAGek2Qmaxa7UsdQFoFXltgWh/HufansC6DrpufgvqhRJ
/v25l6HuXPsexSoKnIy0JrLoDWrk9XutHJtM4Amx/uDcNck8LBXFgNjXWwSfnSNS8WiAXpB9t9tC
MqIDccbq/2bwpbmvh7OYtxhc18nQ2mg7VriIAIAu1pHTUBw88UvV5XlyaiACwxDODXsSC3MJNzFZ
fH6fdmKTZYqE2JzN8XnwNkZopP+fdKEweh2T67G6zZF0S/s9JVAo4a+RA1Kzusj07dLe3SsO09Ag
exbs50QKRai/w4/1978+IKfIMf++N3rAB1NT1X9fEuSu10alXciCKs1xVZenuaGaXOdmAsULGbZw
mH8mN4z/pvKFSaqGMcsOl01AqcjgeLyaghNKvA6lFAqIUNR8zbkb4sflFAwXPgOB8QASC6ImfAj3
/oTNQHwPeSmMyQ2hkR7UoQEY9wHB3BLaQFUdh+e5GDdAoEwzhdtU67RS2cldujIuU0z9C0RmI6xF
84xdCiy+VrPoAUE1odEwzw5X2KzeX9EiBmoi79fxY7dTjpNcGlCcDJdCtE/G+78JFl3O4NES/4/f
m6fIbB6Oiit27xsj7+S7k4KS9Fzx7JinZb8mej7h5V9sZVwJUJZQhy1zeApMPgcswWtCLilEt4YL
Z8jfR9HetoIJeFjD7nNbcJTXpvicLCf/gwbXtk1pPN3bEx9FB5G3zG1wd6aJQxMWrji7JYlPKmd4
G72Qmdo+5BPa/CUJram+8hzGQJDiqsHQ5lw2/2VROmPpaiox3SJTFkFfLRv7UibG76YCIqY18Wkb
UnUlsQqsiEWwRVv2VJumPPeZogyLKn+khyvz3O1xrrwyLq+cQkzmAZv7V117v68Hx86gcIl1+lT6
FeT7dbLrZxapJ32XK9fka+rIIUPLPWngDlN1e6KH+OUzTral+PSCzGHiUQDBIY5bDH2IucfEJtqX
cGGTyPq8kE+1bwVJGF+TaWMbm7ot0vXN+JIhdKUtymZCIu8iPI+SdRuymFU0FnyhvENT49bmg1Pc
kpaYLfz2m1VV0YM0dUifEpP2A1l2g0Bl9hwPl3Pm4ai8hJ7OeTC+I099tIVT95LfqOtOV+FasynA
YHFZT2sxgmV1F8Jfza4gZmHJIgA/M37PjZk83wYgHFdKsVDRmEs8BlvzjDloFw01YsQ7FeLNKXTA
9rNejrS0LoToEHDzoHw9a6bQROWv5JX9wCEMzdF8n8nk73mC1jMGoqbvjMk+6WUieX8sQ+pyANlx
OipcKt4OJ1yJW+Uxj58hEKcsVji8msIfgV5lLXgCSuAQp18xJoGaHitU4vIDV+FV8n7iBY/aAFNA
Jr3wTXDjX+J4JMbSp4hJMGms0J5gnonjjTLtybxV/tyBIArsVWTAftXOdAzquXCknXCKLATcCJS6
z3fzh9cFpPfVOvf7hGcoQuXmP0Fd+Msstlg79kbPFiOYTzB9YvrB6P1f49BBBsvYIeV7cAcb1lTO
Cj9I7WUtNDAeOOXbTemE3nz3Xlsa8e5ZaEje2ZOyRav4uzK8PTxvPV9ZTFRFZcFCku4AS/qSewku
oQwaCEEjalhVu37xRSwGPsv1/WXd8eb+g3huRwdWtRALEa7Gs2AjltRBWzSRETZ6z8bL+F/r5vFI
hRFtznwUVRJm4p1aZjt2y6lGqctgeEaSke5iVrHZXKa7zT3UMVfVWRBAogL05+tRs/UD3imnIvnl
18UyA8o9hU68+h1IwoeA3ELzoRgafBQP7pG3lFN71+tsjpMCYUcZUpcsxvON5eXQRsK4udaGlkNB
+q6n8d0XrYAb33Klncr5ARcChegoGpzm/iy9E84mL76XBYGFaK9Ew9xtZTjnABO9p+Hfeed7UgAq
yKhazBnkU3PzF7m/om7e1umouMG4DqfOPPw8IdKlimCvf/12ZxyeJ+Rfu9bTpIFywr2BOx2rfMuQ
SzONjzYPQgi+/fpOikkJ9ZgOwU33hZgNLio50FAVyNq57O1MfXVfFQqAMPKxo9kS3NYNjzjYqfG7
21TEdlDa2UpmCNNq1gfatZJpVynljrJIAs1If2r171+kNErrhNVYZfHT4CjUDCmRH9hBmYnekwHQ
qOCciWQAVwhPu2+6iyMZIzYPsPgDSxc3uLLTCigg6gRaCElz5AZ0pgBiFKaawCGdnBBdbAPGdKgi
LB3cWM7iml9LXvdqcI4YlKz+uYSl8LPTAAWs7eJM2GavoBzHvXuDSk6oRAycy7RBZD8VIpkBJdv1
CWQSYsMBTZXBvZrsUEQ2/kOqPMhMFcWksSlWRiHLSc18cYQsx9lTGFFP2zvXyqQtVVT0nSZEDcQg
L4aeJhJSojKqcK5Au1qC8jxCUSGOETA8nyDaOu0XVFOAKIPWSxSJ3bdIT91YC+ENZqZ/0AsD58eo
wpAiu+Sl4+j20obs/4jQ8ax8ZE0Ps9SHUuH742hQ9fe4uLkCGzGVU2fQojIFqUzn4Yq0R2ysPHgj
KPhMQGNjTSogn8e9gISO052MHeuwJUgKJCgXCl0/ofLn2pJs2jHVDtfSoQwqEObMdUC964O0PDYR
U9IrdhHy5k7IGsBGR+ey2wk7pbEjOB6Jq0zcTB6DmNPQYrwG5y/1X8EdG86X1P56QYNk12Q/BML6
RLP9Tn0ZeNqbdZyRuIUOWJ+HqE7pdT+8m5f9cT19YAKNm/AkKFqQnHsrYKaqyVHCXBCqRP4xm5Ti
fH8OaLFIFAaTBlIVoImuLwdWNdHJ+KcgfRdO+41pkYsDC/v8WLAWpGIZKE0nIR1GW4QiWaVYjRUQ
WNLjj2hzG1nVBO/qnuMEcyI4NZKm5XAxD+XBhRr4hKBy8r7eK5nnz3nhEwfwHg4ZVlamiKtXA0Ue
aDZtzImzx6wj5af5x0PTbHJQN8PKiazA3rb4U4p2ljCHLqow2AtIVXUmmwyq2mNvdnYXgYvB2VLr
Lem3wiWPjWDSLEc1PaTXRPaynKG4ccU3rWvfjA05NwhmldYz5/AF0VOa+RfgBJoQiH+4ZvRQwBFk
btk9N/KInXrSWWJw93kd3jSfZBOTRhtg7VecO9xcbcOJELbMn2CeJ6PDSeORksfeYgI+4FlPWrZo
UXbnvNTmqpRrdnp0BvzPQJSDG5U4HMzSkuOmTN/ZYvLIMYRnE8uZ3c0D8X57Vwt0MGH1eIA3tcsp
SMdlNUSoYYxCqsiRfP8eRELfxdQ5mt6RW3Yw0ZPJ8bKYzJsGj0Nh5wvHD5vgcIQNCyUnzqoWecrR
OpQxkoHBoWv6oLvFxpguqijpWvYt/rNNDlhYCFO29OmNF8sjGNwayaumN0PkcmpeEfP36xFiJpqe
a7GMA9/bGJzQ0nPFLyAS7eUm3WG2x37aP5omZvYijUQRF5fuOicT/PjbGu1hnZ2kndC7jVGcDLxf
7bysi5+tJV/9DvJbgNX0j3QcQiB9apLN/XNGs33rPDvJwhIxKKOK+19ccrxm9IDzRm0TDTD7dyVI
B3rTV3Mwxuw2fHTxD4Wvldq4jyJJOULxs4nJt96/IzNiywKQKroikQX1ehjE35HNW6/6CfgROCdD
3VsxS5ZNg9fS58Fa5VirOb6Y/6y7sJTPytRD400wErb0orie+1CVq3m37WM7wohVw2wjqA4TKvq5
DYkHi61zt31JRosXikuwiDrRs+1QVBDFRjRK7j7JvIYvbth4lpSB8Xiq/ZgwLIjXyEFp/VLxskuN
K0DVyZHyIt1UDRZVLFURz9mFq3CyLY3Dy3XK0uiGaGSzgrFXsFlkJqqayijtZKVtj9a7oihq0ggt
t9f9QB90FmrfhXq8EOnv7BlBfgcVZPdsrWZ757ERbgU54HbgNb3P9CutZkNryRdllPa17tg7El2h
5JNh70WLyxjGUm3gbFu77k4z5jVqo1gBEtVBvhvHXFUVsvAsOv4G0JmsLeJcGChh01fSpOuy5NF1
a2KlSYfzthycwbkynxqrd3F1VAkZOEyVhvmUkDAugaGAZ6jilMlpVPR7xGjXrQaapaSQC8AAQbXk
dbco7pSZZXkHycuLop4df3rYwskwO+j+5FlrohPN/ZL6D5bk4EQ7k14sksnPZM3NYpEWxg42x5r2
rRJpjAQLlyq8ZfDBM9efEYbVRMTmpHhU3Q4epAa7OiDr83PnT70pQBA2t7JP8adNRnJpr1DXETZA
1F8MiVtPza2++eDF19EioKrgLCH+aHOQvygAyDtCg+tbLsepClPps87nfUpel6tf7qTZw8V12un5
GDFo53C1LK3HxPdY262U4ghhO5Qflq1qx6IRUZ32NokswoMYBbWRPjza8EPcK9YdWUplBRA7M/4G
/ao4n0kDWcXUTxMtR02IgCEesyCfVLDYy1ut/n4tv5HhBpD4T6BAQdV4arKpeRM18Us/Ol9ce9Jd
wEdUKFANGG+6COP8oha3UNj/b31MlfBviAqSILZzGAeGhykyWm2cchdWK6UaGQGU9iePb9n+GUYh
yHDPnY+EjMNfrrGeyy1ZicKEcypzfyWKD/1mpUP79GiiEJJ/G59BICEwidEkNJ+/nfGsB+gU7sQ8
TJZZVEeIE18wwXCcxXh+tZRlphdBct85+BBxXWxu/tdDIyvBtNwuwlVYAcQuIfJx+JZa0zute+nX
QhNn/GvS91xhFIt13qTInFz7V0Ltz5kgj88orDs6gPeh6YflZusLP4T40znCfTt832G9LCRb5pJX
2ZgOFHTbF9f+1WSAjDRzWIPhGB4HwAPjDJC0tKe2leLDPj7wAAQddhA5CSMR8/O2fDBEKQklrqfE
owphnDWKTBajzvi+dUKsT/zFQ5KO20hdrRLrdojeJ/+nk+bQYwxe4b/k1SdkUPse2tkQEqFiqogV
E8oKJYps/gUA1lJ930kBstjUj1FUH2/iKAwf7CX7lWBmZOUhtS9QFvpRgET6/CfWfYqHuMF6hf06
Ln3YoUwHChDlDvNyONCiSNUMlqDBjEi+al345HIEdFNnZW39tUUXdeRNCeJyTWfgPSBPjsEiOxzm
G3PROLy2Sui2qAQOqBUNPjM4GCZKyr3smML88bRr6ZQ6xVKnrAgaDT2pD0rgLIeJezg8hYhyJ30y
dXoCXxWi64tZGqrHwzufpK35UH3azUK8VcFsd2XZFNticPdrfFz2iAHO1IEzFphA5xfnDPU7RZoq
i7AkQ1BzFjT9ggYzhwVyfChkGN5YyYccCm9hvz5uEcW+7nnmg6GoWVK6tlu23Sx+e62LBm/+8RyE
5c3aitELKBpD7w2LE0eDamA1OLBuFKDOJl39oG0APiuSF0bYtzOS6C8mU6JJlYfvJXR5f/tdOZEz
cGPXMFhBAwYr1ewr44+Tz8dfZrmYWp2s7R58W89wikEKzlnDZ7xo1leryvKKmhpVg5xsbQrQ4jW7
i7Rh6kQevGLHRf/1k7dtmFV4mBckxfJDrCFCZ330nKyrE2S8mDLDT4dagXGiR1Y0gYhKEa6F1YXy
yvtS3SR5sr3fTEhDlF+gAoVnBCM/qSoWEhlW9gcJ+7cxn+ARRVh5JX7lvaNaqPoL6lvZKjhakUeM
/RZZeHNkvUDdz6F54u0JGTAUj5B+S6IGBKh6vbarEIsbrRbpeXZGcsdise41EAQMZ0X4Z9F1pJyt
+yj4J8PCRboHCUAZD8Wv+wYt8tYxfbQteLAFTeqVNGGFljOrnymTPdYoYgbypH4lIB3724oD8qwf
/WSpWst1oirdlUtugMy5paYo99x1IomNydQV7YuR7UdAh7pYPF5Pr3KTba3ld+RH++uH+9OHhirK
rxOhK0i1Qr56nYkNDI4DPYBv7qvNmLrVsEUz5DvWRG8BPULITe3qlT/mP75gQXCfLg0GjKwAm0b6
ZTW22B0mQqOqyBkUi8gsjYfZTWxHL2G9kBcJgaa5yHdyaHvGvF3B1govCM167byqZfACGQRmOFWx
lZZGJ+os71bPsOJFSr4sDwX2fRoLY2sQlFdLnxDqRvqCiMsqFGVnMi9CQL38p/ivtIHINUppNUz+
m9DsAV9a2VxgTJmsHOLUTIC9l22JpFJZs+FkF2OeaoEMfJFdc5MUseA5JKUXbz8tSTvHpEIwMHLm
NyktfKAGvezdPLSle+5RY7XbjfV9JpYK8VvL2ltb4DmfJJDnnbPQtaNEP5lMPD5A8WmCbKM969MG
pPgmy5hW5bh00LY7P7AZRunczyXKJlQorLgyJp/ewD5oKzynTxqhuhQlk5/r8vLN47OCtvHA9SgI
uJuQ2bQgZKuHvctyx6w/KzdzXyUbs8kYAz3TFic2CU2DQ4Aon+Qdq+myPmOqq07xtJQs3dNpwxpO
HNMjnATOgMHQG8NpR+9pzFKaI0yStgFykm+5RDiWKeQ2IDURRSWjz99Cx/AFSlUlWF6D2ZEim3fq
cXz7Ywuf3eomrZNPwvHAb+hCaWGl9ukxNyp0pR5AZxLFPlTCq+JT+ZfoCcChfZO0AO/CTHM5NC46
nFkSUacxtGSxu4zVPd3PKXxRGT/QIWqKOEU4p5z8CuJ8xpSAHsUbci0w2njtcmXuDYkeuPWuSyuM
h6SpC0WFibnQqVSkZDpaUS8/mhwbQgHY0KvQv7CYZUxuqu+BI25aVgUH+qiWY/ollwbtLDIl7Ka4
wTsaCHV5Pp1+OAprMgJjE7qCSpzlqW6YgbXFVp+6aKNMzfybGbJJyjg4N7+M20K16Q+jmIvJwdDv
m0LRaEYkphHzI+20AXhYGcHhA/uYz5OAj0EVotk3E504Ox5Eaz4neFfg8uMw0a6dL1bJuBee4h5j
qji8ap37UnMbzbGTQmhZW9WrF+DRng3cDnCskck8OGJ8+7Ah/tf+efbE10GEpNiIUtTKL2F77lUE
gat5Pxqq/+qyQs91jXtDkv0DkNk2CsNWFJJA9zjSNEjj13ckEh7gnNdFLy3uGYbWhcdiIKgkJeQ6
PCPZt4gCKGBY/B+A2GMEu6CzHxkQx+htfOeZ2IRl/xzS0xw7bgkwVdWHzInzYSDLF+8k8hMOxOvt
7vBiERAVgIU4Ea0ztSgP43xcs4KP40Bu8d3APfjkmiwrMHfnVPVT5mISH1sqZJd4eN5Ir94BFxYX
orn+je6SzoYhVpofYHYDG0d4fL30COK2hofBaEuL/nzak636oyM61DiL0kHhxBjQoERP9bQHxNxR
iSa6QxjH4+ez9BOKHt5aYZEvbUcXZbev0d5V8zmFiRauHeuBQHVQtZC5AcSmmVAIoBlefUKn+SqV
xd3nBDclyn102GXxp1hcEOmUeCgiXyF64ldQ66omGTtPhCbbRxqXgKra83RzIxIcCw4uwi3WL0M2
3q3xRMidCIR0Gn6cnUoJlRGzHPBp75dKjELDfZd7kLuBm/dW850dsjSoGicl2tieZ/vHerMZpIwF
FqK39Ff+ztK7s8ohOOgajD5WPlw7jijzJo80kP832c+VY872Yg87etXdpA/BKmDsXdb6IJ9J2Myn
upZxuqtoaEkqwcRjur9MPy41heKslfSHr6nGPBNf0wa+r+sBkCfYGMN5owBHpX6HIDulQRnSxUU0
D/4T4MXL7gsfTqelzbEFxJvo+N7pZivQHBFd7bUsZXervs2XGfOGmUauStB+wGms+dD2+37W2A0E
+8aRVMl3Zj2F9MifGsjK463HrRZ9rXlG2DXd2+bZhHRb648Oq7dgtQZ9TZ5mkVZPX1CCXmIL5YrW
CJWD6sfQ/7OJLb2x2ReMmlq1i1G+IVN6e/BLxUHdTVBeAn+8HsE8u2nCwwYtyObmtnPJSqgp/mY4
EgqM/cOBxiJO1ycAUyOWmHha3tUCr2YRf9xYBOZH5fln6c8u48yU25PdmHN2f1Wq51hmdK0OMTdb
P/nkyirs69qdlNsfMWXyKcIfN1NGT2HzQnh51g6CM/8ZJTKlKGiELd33L1ZeM1LNdkjwg6/h6Zqg
X7QEwB1d1e93Lh9akxBzQGX7ou8Ygc10IcMGChLIzajd+uDiIIuMu5e+lCb7TMJvwiDBDywmHNVS
POH6/QMwSbKfDqNi0E4gscT/RpDU2nsumNHo7Cra4Hdl0wHyixcS90HN1jE+gQ1E5tBxgPSWtrpG
JYhuUdfiw7WwFq2jFIUgp9pQx3lnjuO7o3P/Tvy57VDFjixlpigFMKtqIE3yiyTjrFnK484bYYuj
PgYmK5O4qmv8pOh17+IU25hK/1E00vaUuVX+zmeIgT1zphty+BN5DIsxrpLWBf9UBqsWMjVoTpZ3
0yEPNSp8qbbCV2wHWHptM7jesb8qdWkPUgzgqrsm6gpxGA6qvSt1mlO8B1qWcCezOY8TUR/r0Pl/
TdOuZOwXvy+/cBswwT0s37XHi5nqmlDJnsIqeVkFrum6DXQpiVyBwojbDAcf15+NZtzcRY8aTPKp
hrKcLPwCqYJ3yHZftm8S1w75yaVFOKPxlB0wXFpZe+Dtp4qrSqaePaAoNVXLv94x1mA9Wff+vsy7
kBNuAZdlWu8ubT5NWRVlSuoh0HOJbZND+qsct16orfcKFSw9DF8GLRsi81H4JggANAl5y8tdFqwY
rYuWz+89H+6FMxVRVu9zwmseIPNpOqVkxFYG0I5zVPjX8LQigXxNF4e5mxOeO6YF6Y/erLlCXyfy
kewFeJBUV79us+32o1v9Ukn29kMlmC1obKsYIsJe6CnhsIyzBbZ+B9W2tnbFhqtgr43CO5nqk+Gj
+XPDVHrPaQUjx9AhNmgOdh2SOhl1zAfYYGRoJyZ+fwkhW+f/rbvuAHGLPTygpTQ3ZsT0BrjPLHT4
O4cA6sJEhRpUbh2YcGcl2pyTgtl9Ej1ZI7cYZpsioPKrbJkjYjoLZJnh1YBODZrc5jh6isxbgwS9
v+N5wJPJtzWbP8Z09qwcpJZhnb/TBbK8DN11XmJwS0TwrTatLPMSzNk+Qsg3i3qU9WUogQM/KEVP
5PkaM8RBJWZ61v/UQmYe9gVADMWj8EDblmbIRS9Vjs+J39I/qEuQxf37QcDuTgLp8Bkunm1eUV9u
a1TMQk6pVtxZ4FrpO6eLoN7/f8e3q7P+MZ+4BSniy+GU+oHkIDPoPnhvqonBsIMcvNMMJ4vN10BM
Ki4cerP/z54ksWAdP7Xq9xSSL0Zv/qIxVkuEsi+XutmveAgQTe4Zqg6G79BEZpbYiK3G7J3RIh49
Br303/quCNi04RJiHMFnlZsnkKzitMgt+RpNYvGxVL63kWEgjnXqKWyeLOhRSg2oPsNdt1AJ+BTi
qpwatRn5x6csz5vN+HV/+Rvm6npK9JqtNxkcFDGTlvdBbqS+xEyOJq8u1WC9XOnHQhmW/qf22bzl
dlsVUKONaSa8ep69zA5oxkTQ9zzlFZpYz26Yk+fsQaKGarhvB7dS4odXQ1WUVuTAlIRJxh+5PctG
Nn9kZDQ285c4IDmI2FMYsTuDoRBWy2vGeAj8U99C0RK/LihjAdp3HnLRB0HhFv6rHcuP4Cv32jru
hqArKG0cWwsfHm8+Qa4n3ebDfH+8PVuoypPJLrtA+feSOTggzGGRHhpwx7L5X1K5gd7wm+P92OAL
UCZy6WO5Oa/ws4GWTWwTwNYc6v+9OKmlxs/eCAqffYDwk/bWG4VGv04muTGOqNbeqk8C/44Jqm+E
+Uv4foDh31keOvwUVKhO6NGuuLBX+MZdlT1yr+maIGycC5emgnhgSlZDXaMgT0OdQZFPJc3ghhuX
2jL2phdpA/0n1YidClUtBAC95yt13C5vUIVQYXken3t2Vjam6S3BKLfqVRQC4HpeGb5v9XEGtxNp
+64nikOgbPz/uXiMsqZvL26d0UtsmFNeDPbv5kexhjgOy92oWduBhGGaOVYd1DiwkyypgBAT0s4u
iAABdhMc5tooENXqXc8uFCY53XJoo78w3YoUwdBPeeEFrzwKbvfVD4e3aHkMew+oBuysaSYLcVGu
WzncjTxNPgF2PUhU8nuXz/gc7qUCF4+UabfS4zjyPg+goy/+PAO+srL7+CXP2Ll9d+T2rx6KKwDD
jGBd07f/hiU81BZAGpY/8Adx8aan9GdoaPTzhyHLdQ8fVv8n27YnBPTQjQqs6DpGJPlZvYUXkAdJ
7o462DY5/BS8Hde9TZFb5CXY8jvbyeEk6tNCk9E+SCYjmC5rbvwnJDnCGmPU6tuJ8R88jbobZDxe
MILJq9Ij7tUDWTvtPm2C6bw2cb7j6vX7LHbiBleWKtvWt5u6LlS9WBCe8CiB0tNliEGU7f3hL7v1
vEHuWhcF9l1LWNgHNhJCIVE1jrSiTw5QqjUlbGm4W2rVBSfg+1rReLpLE9jI/h3ZyHZNdXk6CLI3
0ZbmDPyRzFJgVrHmNh5TdajD7271OKEQFezZzAlA4RCJ48wRi7DPNVNMVjfTuUpU0WtZl67IoUPO
erzm7zGdJxeBU0MDGZmdkrQ/riLVaqXOWuv8OKIqaL8GCF/t4wux27B2X09XUmxMlLJsLAPVuJv0
MLc8YCu3JCvTndTDDiySaBHwXMGnKNDVbN+368sucSG3Vd6UQ00tKYi44MwxXPinpZx401NlOB1R
h0hEdlWn12obAaHQc+mlXTLaPqLhUp2zgnfWWSeOZk1o7YeMEJTseUiIrexLes2XjeFv3Yycu8SL
R01AJluGZWevTpeJOLRc2TxO7ZPovfMHCwtnXZYfOoXqt6WJQLM3vpjk7gsMRFnzLLjY3lrQ3exn
2aH29NzBNfUIjb2EHJh+2r23IoCtasLKFqwAJ8N4hbBhGI/mb7Zg+I6MHE3RIjmKSIpiVUhjDFMq
tgKotCK4ijSzRdFLbrEHp2e2thT4zorzPz5DdCVkbcc+JIygz63hhAVnMAYTtsyltJ9ruLNPxmpO
1/bc897gRbk2if4hNfGkKnAZNJKEdHaH3z5eTkUoWKlgJZIPfMaUkzwJejahJBg76oMRN7I0PUKv
5ExwA5b2hqMq9KhsJN7mQGk5t8Avz37rdiw1/RBnUcpGji4mFdljbLhsXRRMMupcNFMYSLspJFmu
a7FfLyChedPmpZ/DZ6OxebANT2oUrETZIxQcj4UO1YTqoBRbtOaHS9wS6dcRtk8wgvB1I6r9sTZA
C/is/5PizifzTPBHbGyn1xg1L8luCbOXs8JWFe8s5a8cjOv/Ov/LXUSCW/iNfSiHxwNiXsdbL1Gd
iOD9CoKMceX8s768Qp2FT9gn9a92/vlLgKeWc1YPR/AZGQJcnGyQ4rjjcnOM9zpEJG2eqlzOXWMk
UJZmySDnz04Ke3FzSlUNrw2G3sEKvz+v1xoil4dqSt/WIsTpoCT69GyJe084URZa1X8FaM83ne1n
kM3Wt1g43eLHKLYITuNwc37kinTnyKJhwhGcKe3GsnYRuXLVVmQ0RP/ve3wwBnX1aAxOjEFwpJX/
olcxeDBwJe44DtRxaLQ3IaHJrribzkuFwLl/gMu4Iw3jQgPQcOYUT8bxPmBAc/qiUJ43sZh6Jr1s
GYfQO+AO1qSmZA+emaLJHVVz+qy0Rdt+9ZZQVCj4DO2y8vSprak+bahtDhpl4tqouMM/1JJ0PtRG
U53clN1QOY0Oy4ks+SsjQ7xi2X8Lje7wQGdGxR2eCk3642K0fNcJgehefQRH0ZUdbM71TnbxGT/v
xTwqZbmgNHW1y4GrHrwncF1jctem/uxeWeaZZVN1obv4mh+K8Nnb5NELsOA5LICv7O+5VQemngRs
vV5v/PueRiwYyb+ZMAGn6O7ji2s88Y4Bz6JWcBi1OE0n61dekZZ+pX1EdgM4M5pBKo8VO9VpA9f7
kvNuDY9Bpzz81P97IvH1vKUau1OW/UI2u3virj46RD6LD/v9UL2wnalQJjQvbjy/q6pfZjLxe9iY
bpAtQTtVrH3OWOU+hlzK0YSwiI3YaVaBo2/6g+qbAYXLMbcf2NLiUCmWafCY4nrYRU4qW/CrswGt
x/SkquY3U66MF5rkSraLuSFrqo5XiMotK9Yp6IG7gz7i7XrBRYA8qvbM2yGju5LoC/eCYWcG/4l+
Vtu1PFsxFsiEiVqE8bDPTIEha0Ns9pYS8aOBIAAxzs5hTm7acZ63B99n9jh4vgFMuvx7zNCKmOn9
HBQ267fSCRQN2mhAx8bOQ/Egxh2HvJ0c6kAjjdhzO1ryMttBXHglmqPIR8Z7PdTJb+fSfMmE1AGW
Erp9W6Y8svGMzPU52tmRkV7W+LZA2KaHrQjvv4jeZ6g37WnwetzSqGtwmtdFinVCCInEc6Vwz1fB
2r32oDAJmA9vDWt52FQ8SBigFgpG80ksUeSD+DSnzCjmebeR29/7fKm9p3aNvzB8qE22zUsDaM4E
DILJSJN3GnIQLqQUVVMBng0Z4mBeICeBZEzGTty5GNQi6BvKrFBnSz99Vj0j/uWhGCIe5Dp1nbxy
bdB7DeJBP8JANfP8l3N02feYFVRyzjhgUVkU4rnRwbbRKc3kzdeCebz9ASJuur6NpqBszBczNCOS
yad/ByQpiGOPHCTrWVMg1cwT2tv2vxE3YPRN22LEHVnAFWMTUvAtAxDc0OCoNwNbokwlHx46dPen
VB8tfx10Z4j13gno1qBZoFr0GmkWnf1rboEdW+czQa3aExX1WMmKQWbJZg1RJwQa5hmq6kB2Tazm
GBHQnOQ5cfzadeU+stSQJdu4m/NOQhIVIVEcojMgCDQB+XsxVaWt2jYl7PTP1IrtzIljl7pQ2cen
f5fSiJwtby04YdBGDDZLb4YZq+fneWFJapp3GU4giWvH9o4Xa+44x82JQ2g8V7u9dq0DdsfDo6Uk
QXOTBDKrEUS9Zgul1BoY2ZRDD2MR1GH5ZxOA2uePNOS7dcMBUSYxn3wH8lxLK4bi8ERl8ZnL0Rn9
8xHcsfIZW4JHAo2jY8xj4VW3AFbfZAGiMzi2IvlsTR+bJY4yS4EA/zl5TdMRxpvCZUnfb/bIfru6
mCVpZPMPv5sc+qrDAqlIRBlPMHl2QORXaqnwbwgEGW827dOeFB02hqwA4woA5KKlo4NBAQq9QdLE
5GjyZvs9j1UDK94co/UyL1yngkriuLaspC4djiiRYMYJskm7GRxxkT38eK/ZOjswqRS1oA7Rz9Q+
PdIeW3E1N3SBSJZ0Vpi+rJBBIEIPEgHXSQKdnL1otXa2AkNo+poCFMDzr51Tv6lpa61nOpPd72dh
Z7wrAj2L7GDMlsXTl9ZKDTPC+4+izjKFYJoJT1JpNhKVTNKeZvK0AkNzIuh6baATJLaBHX8KSgeh
FXh4KUDd43kim2QI5QXhNnif297fNsj+qGYOPcDzhs1CM5Ow7cTgl8P7xumwiGZhQXm0K/y7KcTX
CIh3IYZhmuaU0c2qjKdtS9E+ehrIKp/lPUNrxfJ56WGE1/QrFKGeFFoEGVlb7yeKi+Kb13ufkMUZ
+9SI8aCu+sgYIWZ7pCMqgeIjEsk3xBidghSx99VmVP/4DVU4EZN1Lttrqmlk/ON+kmdgI3obsQJX
i4KSggyg7gLeIV+D12Rydf4RGdRla5BYNZyHE+4G4iBg8GqcjPhz26kmPRDI/onYatpnNSQ8+kuN
vtRX/+U/jRMFMTaENeI70dw2iUQJ1CjptAzNzP/B5CHAiJDeuWiGPPc+OzsNNj9XCXLyEPrn+/uS
0Q6JSyl9uH2awuxU4Td1Lqh2mq7brlyn/BgPoByuoJ0PooZirNN65bY8MdcIF3n4uuW8jBmDqP9q
2EQh2vQr99LCnkG+hrPbu2fe/ZkPk8SC6RGcJnT2vwUqrmsVceotMQ1CrLjDS/NnB52QK9hjrwRV
wwIs7prEXz7xRA4Mk3WNzh5MkXOm/zBz8X/wJFNtknATqR6rzFkZ2UZ9s4+zY4m8OXYvXl5AR2X+
DWMdowsPVAFQfb+08coAHcH3XeY+It1IZi/jFMGJby96ppLk9z+0hjmYEcB0FvA6zaoZt8jRncml
zfzYKsaeWS/G5wOrtYoIOxybN/mE5ZJcyUAaJFouqqMY6zW7IIXGbligxiUZi1N0YQCDLqkXKHcB
Pqj7VadB+76dqMnBxOhzNsbxeqD5fG+4GkdnMk4mDUgXcsb3UEiM4UaHzY7XYFbJooVp9zaZmINy
DRtJhl0sWgyV4AJRqJsZ54TFTDb7TBLVEzYRp9YKJ7EpHocLgF3HRlvmxq24F7XUBkAcXEFfof7W
EoGOBFxcPw1RA1K4yqxN2/FeAWwHmKCgyQVdVcUlaYYclBRiKbO2PpKyIa0s6SlU58CQaNfYrAwu
hkL/0q9t7q5vC4ttZdof+mckzEQZ7PS6cpq2Pkonfv4hgcjIOLGgbVz15fxDsPypV4vUGKPQL8dE
GOA4Sj5wKgffPKGWc0r9RB3GfzqnEb2jLU3SaeIFrn69k2x7rHCZXxFLcZ/P+nrE2U+zQkZ8JQXs
31QqTBbDaAnki74xqqlVvp9fBRWTTZ0OWsnXMpat+ROSNJOYM+u50BQjenEpDxf2mXakSmo5UTpz
4L4QrTJgBU7Le98L1b2/ni3rHSTGuuVIX9283Ufc+rWxh4kPCgGaMFjIa+rWryZ2ethJzCWR7zix
PcQluErk4xNPnCxOM4+LMztRClWRBFGlDOMZ8ZW45oqRzSBRyucjO/X4F84OqWjPotS74HX1H4GU
AM46fJ9Lhb3LDcf/1mo+YT0oXrKctIezTvxoIgi1VfMrtTpy+Sz7bsKEv8OUiEHoctr9Dg45IMis
jEQWebgUYRcZmgD7sz2Cslk59rSiBLAvvXTll+FdlYSBlkb6HQH2RrouaiZMEyydYMzox+Xjx11q
qxjZITgQdtL9ULERPf4VKmnbvORDbr41fDKYMjb5vTizbcTfSyex7zjNAS2fy8dvo81fQ2jY5gww
KXY1i9OYh/lYmMs6ceY3L/XBbq7G0Zgr5I9vd0YDbUyVLJvZ9z++s+uYq7T1JRHJBCSSZM+mXvyq
ocXFy/gs4t2wEtxi3aSnLqPiMWDShRdFbkUmRMfPpsgDw9rwJIG2IB5KjkTD25Owbm6OSug2YK5D
AXSPqqKH1nV2XQ/jn8NdKbKM2Vul/YYFqSHfmTGxr+s/TuN0+foqMWY9AZOrhO40IwMCW1QXG2KJ
pRfN/SlglT7FQvUHDG4S66qF/qFzvlBRXCbkYlQDpsMmLT8DjzeLr/x1F5ulJTASLg346iFzteZW
8pSLslByCxF3oULba+Sd3gaXYY1zKexDnSffr0asYZBWArpmAJTvuzItd+sFbzJvCY8XzYeFgYsj
DrKF6WoQCpnxwYK2JOVaDZK0pUFUwdLMeInzsMhR1z5RBQ5PxFNkIGwc4YtpY6A42MZFZWtV6Trz
E9Yd2T4iPdmBJkbTKN1LNlGRQRoMxbo8SFlcZiVxYuvR79GsPN3+sfDfhevZDzhmy6fiBICsvGpJ
IM19HQKSzCK+/ZZAGISH6juSuAFpJqzz+tY5QB5WjI2FQE1F24W3PMsT7j2cop+TwmgwexDJXL+R
jjxJnFluzKKZ+ipfUG5e0KJBIuFW1xwAlYIE/k9FB6mMsbIhX0CF6D0ySvDwZQktv2yUxL5YTCKB
USHdaZaPz01+V9dWTbvH1YGGoEHZ+i2+rf6Wq7yWor1lnR92IsZnkC7KyDaKNsHZR0uaBETaL9c1
xhkqHQkSYxTIPcmhSncUIqHDMyqh9fLu5JRMVM6JH2zPARV5FKDd9050AsSs9Nypr94UXHYbllBh
Poqbam89b3CvDOVuRfBDUUvcT7DMpXM1xkm4VNogu2e55aMKMxO39cKuMKOYzSwUZbSIqiYxXwrB
hPEzQZwNIkJ/Xteotfjm635goeM+LjThIQepONvS9H/1oNuTNttlP2X8pShrlYUTgEHi7VSqAy7N
sbTFbkoXO/witqec+g8vsMmpZ3MHLA+HFSFsqQSb42jNZevyaAZVFOX3eJ+gaHl6+UgIA2WG6k85
TQZOLVTonN1stAlb3mHaUsojCccgoICETbThkLdK9Yvsn3vzY7WQLLYJvBhpos4hKLP/7ZLAkj3z
oFT0SVKpRNW4E0dTUolsQH93Yz0bq/oOZqQzZhs0cgnVD0F4qo/QtS1S/YoLjcx8HL8nXtDf/lWQ
CCDROyI0JRs3P8MLhuj6AbLdJ1Zor+gTXTwaBoEhubcIHga9yIj/9+jtbpctMBwgdSXpBekls/HH
+12fjB9MAel9n+2MPKDsAQHPBsG2ZRRXWNt/UwUBmjMPqjwug4Wm2nYze5GcUF3ep6IGYQkBfDAF
Z38Xh3Hn37At13oNgM8aw0AHGspRTgEcjuY4Rq1SZgsjTHPCFvD7rhdLRW86y6FBGVj+NY8Gbj1S
RGM47uhxhexGgRAKKbu3OEmIZ3e3bcSCtgMD/2szGFj5Q3juShmCFGR6ftEg229tg/16k6NEfR6k
MMJWVnTpgakP6g/WBnMXjk0avHNoDpawPtb+tTm7A5VLgIScS85VfYuJirTw/LvZqJXAKToDmlpN
NBynwn55f2dWES2iKx/0bvAqs1BUlu8GAfdLd8shY2qZ2ADC4yvehiB5+QJt9wXW/87xhNc6gzWi
dyw4UQTHiZ3A4ziKB85e873ehMsHqLH19MCrlYaTa/gaqXe1u3wW5Ze0tI2Q79lno84rsjjzvXYe
ZQhVM9d8nAvg8YZf5w6wKPnFVQOkVchOG7xELXK0F0Waf61witv8iO9kz89Coukt5foWz3AAZqNH
6qnqR0tcuocvFiPvrRpY1sE1W0umfsYTo3VJOXnxMdkVJEW1ES575FDqmw5l9kdpJoog65g26K6I
XkShqxWV66doPG2VvI0kfZqyMr+8aCsriB80dPWQU49SAt4uiElKYUPwdfjZs/hKnbYXknb+2xdw
7IJbEzdfbSKyG4zF1L8PlDRiAxEiigc0fJyWCAaJqTfk6e9ONXp24NpheffGpX3iyMrSi8tA2SEx
a/+ZNb+It7cHul6TDqkjQ6JXuGr9slO55G/S1qxdBTrRy7LkUApFo9cddzgNDlQkt4CY2h1eJQmS
jOEDkk6qA57jW2zMPxKulYKW7bLwU+VObw7d0iLKHInfXsf0PjprJJxCSbY+z93wm4VKrdItMqaO
lUy5lVI0S7FBKYelnAyeKxiz+RcU+r2HesgtrD/J1n9gDzqlytPr8egUhBaobghmG0XyaarQrbzx
4tTisGr9M+nblhC9QkP7BVUfhMzSruQwcsNn4tcort4AI6e712NDlN/Cr/KCCYEeVFwW6hUfk5gt
k/Y7LM5DaA2CGhIdBn7qJisksDECJaWhxQ3VrIPpuN5pdvG9b4vHxpQ8bKKqN5/9At+Th2UBAB6r
uGq5kDHff3a9mcxsdxHhLNzJN5nSXZ4ru1DLG6KFtJGWvT0xGRJc43uG2kkmjl/POwSeVaSPIqNh
H7A3vC7iDS/o0LXsNkzauQo8L2MeBp3nuzxFKCiZ7/T4hpNDEYr2GpIqgBZxjAMwKiH7ib0/Pm08
u0PjUCPJXKxthwc45W20J2apN4rboG2fx2TjGF1aYLmxi3wqbf2Xk/jMtwI7/I/ry7eCY76mbsh9
2ukk2Ph4O5F8AzXiJx+QyhjVK977FNFOvn+HJA7f0Md+7HZmAaC/xhpm01rN/7uVkda8WZ2UNd/a
lxzH63T3On57h923aPHU54owQVVMWSlFbzSV+ycGsjVZxYDWlh+anxca7X8Qw8nUj4dx6Zo+/IeD
Wazow779AR9JpwSttJDCsHBuopNKJQ9pDBS99w99acTcAdudi3bjWAX4mlOvr7Hmsw0HU+buygkl
xyWuHUqjR2UWccgfFjtIvx8VBaXuTw+Cwe3zsMDWceLdfYn7hmgCmbG2tLtML5u/bBjtGYn9u8Zx
0Z5uZ/6S5ScXGtYrwzGcmJm6SkKDomXxc/5KF7LjWGY+54lWMjPD/BeyjMrOkSm8llIghprUe9fO
PaAwkRwD5O+rOA1VEjzQrUpJ3o45l9wvjsyUENQ+QYVQgajwKZYEllbLlh/XZX8roDk5azKv00Gm
iosJOipB/oUeM5YVceR2f/8qXhE5H2sq4u5cKXrJyfgMKlyUCJV0tois3gnmVb0NTN0SfmFDd3Dl
jr1CUrIvN+ox1DrfZxBn5rZwcs81njDInCyPSZw3hdcPqWOsAqq7Uf1Dn+1NzuUOCcg+i4tLUA7h
RCmM75kAyarI1nCI4vuuyNn3ot4kL4Aht3gdhNLCs4mMtMmey2UqrD/MuLDjhb4tbP10cthzbXp3
pGDmb6NbZNXLXnPJJlTFpXakAt+Qnb6LPDXM7O/VwYHX3yYFSzPDgPV8BPSy82GT+i641q9ye+EQ
qx62kSSM5dNGohXuXz8oW4Vs2CnrGigA32mNyfROPFYNs+ZBb0ZQg9/MOXTWNidZH611LAjwTG/c
eTUoqHjg24hJyuoq4zHJumUe9BjYEmuk9fTWgXK8xSrWAf4mTweWUdDeS+A5EDXebreYyrOJca73
YiCKWvuIMi2K2MsjRnW3hBTle3re0l2oSDyBKA3vqg/7FKbuge3doRv75h/MUQeyv4yc2PnMER5n
5mi97S5Yvf89p5XbGAOLIhYkYu8Y7BPPYNIB5pzlQC1MqKH29pcwoJrRojiGuqhSYnodueQERpgp
Tfj3VHn/lJSWag15gN0MH0XwwDmWXibYNdHYf+fjFuPNO8FZoAQ3cz692/bhB+ghMGyjIJTgmdPB
U2WionJ4cciOkQuoiUa6qkge1V8vn6Bo95J4Dpk+RTGlqY3C56RfbilKVNobP4joPI/ruzF5MdFr
IEQkznNMInlbSdhuMEwZxsNf8Twa3bV5XBXt6SJAUtSUSFXJwZwcS5kjdN/VeZ6dTkFVh4vRQjcp
3ja7/4Q8nHqiDA/ErxTvWGIN2OZQP6gyXwg2Vi/DlOukl95/8ObHlPRwJcLFECeu98iVJZLiI3i7
H92qt2cJHYvui08Ly8A8pCocW83NbAVN519u/BH6r1UfmU/OJBz89YD2ZqR1aUcJBXnX7YjTsxdp
isGhePqbmOodfnXi97xujN4e9LcwJIdJzla13A9OHGgzQ7SWxjlcigmhkYJzqVi1Lh+2cKysQLyu
osPiUXi6jZwAcgQvhR4ySSrasMxT+akhzfEMQepRYOUtvEm1VeK1RC9RJLWOiBKVWEc5A/rJktpD
ZedsmGQ4JQvF9/sGB6OzNWHOdp931bF8+HsiD9U75ZRMHmanfdcdS5jZzY7XVwWHAG+NTZV7An9J
G1yiioJmsdVsYr5FvtSFlkaGmS5VoWzowRGA4od8zkRL+KVlyWopS9xULgghETM8xWO80vuoJcli
6xuht1ofZBAxFTQBnMiQERbUS41JNxLOVFlakhQssBx0skrBq31FXUc83ZCkhc0PdRK01Yj5ykHr
A/bJVypaf84ymmR4CTiIteCZle5p0NEKxroLYxFLiWTmTGEU/qLJjde9rwNWqfsU4hDi0IRQfGKV
tsjard6veOVRl3l2SIQsLk65OwDfJwG5qAQFJUXrBYbj1VOUYysvRBbMgnSXnHoqKFUvtbLSZ2qS
eqXqXacwvMRh0tlgdgt3AJUpVMNeH/UJFOXGxbZS2/sGefVa1rF/RkucBIKTuyJkXmyii1c564E0
jn/2ReKOiWBMmTU5JI7gLH4VWCDR+s8fayI6G1AMaxO1HqGVCFMtQH7k3d/8U8RWU4rJMMQyhDTb
80mWywQeNYqlHnANAKLftK1cadjmn5WcuKrqvhMeeDY/n9FP0hSSiDOcEt/ORuTdZPEY5CyYEv5V
SsxXyYEnjJOZ8zdqLlFdJGJyMszmFDpS56qCwPdtIjwJLAIdT9AAc61cdf7cjxvGbfGQ8RmkEhq2
xFu2XvO3heR61L/fP/RzQEiTw0hyS/QC4fIbQ97fIxYTiEEmot0WgRosr/zmAjZ9kaPh/oefHnrP
xJi5Z+IiCI+mQw3ElSt8NCo6E6CmUFny8zmjPwAD/qqT/+gg5xjD1VHoXJAsUVsvF3DGp2ztojI8
sQhYxXEcByk6HDZokDlitf5igEP3T9eSz1s7teyL4ILTVAfhLgeUi4W7m/B/OrOAjH746qAEHr7Z
Zm5FUAT3xu3Vf/cqo074JBw/oAq3tMOdVaXiLyNcoCbHG0kWApDlkfdcquP+RjyQJCFd1p3FsFR9
GN1YfWxr0Z/+2/MeTFf6YizaElVXime8cRLmQhgQwJrVbG+bxBwL5WJFdvkR9xVzeOyXB+JSDhA/
upUCxKjKJCYUrQzCLFstLuBWhZJyngt/hN8qVb18x/Zf77A+NHnn3q8uVhuXbI41Bjcx9GBycTiG
kU/moUtUWOw7Rz0x1a8umMnHx0Z+T2M3dPKu8mip2usoBHe2717NQUYiQCTLMdYhAwUJ6vxo171P
DEqa06VtGrL5NnZXnqOKxd6iF8DOmUrhTJfvkjV24boCjqOm+pK6bqvKnePOhocTMCh5JisBJRIi
YIcI29V3E3491ksWRCM0PoMp39JfQWdaztjzj/KZZfhUsGuhcGXV8R2XHm5575wwUw9OqMQkeYAT
xqkbyRvtQjmtYAZUxBk5vNBBMGz0QegmFwBgF3GSOfePfDw14f+kvYhRjVpKHlW0gD89z4vstN/s
eSm7ORaKgyLiK9SweyxPcOAJaG7KCIbzp2cKIHJbxWUYgdzQO55hJbXspCKrehLYgpieK6zfi5E1
ltzm1lkz7XjbPSDJlutZZB+NwO8XNWXZaV2M/LTXQBaBSNKS4CDZ1vl49T7tawQqaSNSV1+fdBdv
hQL3SkZ9gTLWHCuOxHkXzGbATQEqndVxAQnccozTxLxo3KKTwAdPKQjcNDBLl5Xl4l8apVIQ3A0i
c38xI3jdfPak4ewEQEsBgWeYLcn72CjFZbQBC8SObCzTck/f7V8OMfrSuj0k3NvZu2RpIkT2LAa5
PaOTQy48J0XhP7ZjHg0GUq5+3UPmkQLPG3HvXccPIWFCD+FJiDQX5XwXnOAK/DpeuZqAj3zVTxHR
c1p0hrU1IJsEBV9m+JRAcGEsUPPnvW862Oc1IQfJw6NXM8B53/ATFJqN0vLM839CytwsK5aK89ol
gy1fvo/POeGcUQLsNs7JM/s/8ZujUhlFb7zUhG+XyJkd1WSzjsB3S615RJK0dl2UB+YUhRoUAFcS
YX8V5anv51HmwCZ2c5tmza/jraO8/wQcbTuYsNyYZOD0ODFPhDKhnSByB1iSzJNfve8YqqQlyBdh
og1HzNlEEC3HCjr7jyvMVJnGZhooshojGSpBoVl5K7ujaH5Nm5If3Y4iKyBlyJAM+q0FYZeFdR7M
bBR/xphltj6z/1mwD1IyRuIHN+XgFoXJ4A3gYpzvPQXkf6bojJqJtfsJSBBtZlu1+/zvYe/pDDDs
F3U5ESoQJFuLfHjmuHXJIBkQoYSVIX3UlQELoyirM4XtiXr8wTdYIx0fbIoIT1TGjVhBKNr6Ycgj
LQXknr55PLDk3Y/gOtZNBR+D1EXNnZFP4SfMzeYUUHlVRJRMp6GWvY91eZV/oBUMxGyfmBDRwRtK
DwY+urZJ+aeoi86pwVMrGSVXugU2f1bApUODwgP7exYYFePI1y/LVenN0UpwtS7e1JQkZaDwedor
P0fJtdyKUOxnJb4bgZrx30mldzg90N5JzhbdA3P9iVAQhJsQ0bqfUW6ORGAcbEGSQUPS++9lVudG
gYo60aB9U5cf+02JGKLzFXTr2lF+7PfMZIWFIThh0QJJskyboKpyCvryB1j+qJ1/iNs/Jle7bYIK
WZHV5OgCbZUJm0sZMrH376nFxctP5n5YryGXADC7vzTXSOaRi7xLBhZTKw7n8xFprtvyY1hja5nS
DAZIa3MFTFoATkFZtAmYfIVORjuUn9uu62WOpYLnYuc75/ASdrcRdQbNdd4MRJ4knPLpcKi/FPx9
QCq4p6HbgqwwlgPbGGFOyuVRfMgm/XymEiCUU+nImPjna6Jcmn705JyyYNPEIVur8wHR8GzJqM8C
QWXc7FhvJBBSTZ5qPHtHR9ocZGbC9NbCSqwo6oxhynCeaQ4ov5KIdALGfOD4cb867piclmCmg5g+
ISbJfFmRJuJ7hMmJY6SeujDhde9AomM+fYaQnLJLRJ2VCkHFFcNSgg7UOh0TOWZmtO+3Ln9WRD9b
0T0TTjsMwNA9PnzFySR6r+Wel7J67NV6wANOMVu6j7oWivWbHgs1YLyU3AXWrcjrXHuBIVaSHEBg
zIGHtFEXpewd++fl8wqFxgLzon/+GWQ5KbjrGRcBohhU54UBDQWKRYWVN8KKl2DhJNK3zx0tCBDI
PCmAYsGCWfhxy6PN27+Z+BtyrCUWEQiRPiknOf0AbaKLTJWH7SiQ3YvuFjJp6a3AdPTKqZdxhci3
m4CwhMSOz00PT6aWUVlIFMXR40bIdL423Ak4X7iA5QXbKatm3QSCLK7rJ4I9LXmdlMC+un/oHh2d
s6RUpL88bI8W8Pew51aKdDXDGo1IdjukNzAg/2UsUSkNO+viknijy7V3vEaElIedQ4xai/udv70T
eONchbNBMsMfvs6ZqsefmS3v1OY+f2zz0I7VkMuMk4O6ctZPArD0xXrEwa74sOjEmMa7IsRca90H
mANOOYzPzOT23xAZEkYQKQ3rNRayA1nDBaFuUyxYg4rFmD9aNWMq38d2fhjnjI9dSOB+52X8Mu5X
VhQYw2KB69gH1IXj/qkathLo2t+V1Q34wUn18wcMgxSrH6NOMI/AxrvDovpQ4L2kRoFUroSwj8GJ
6sJtXXMgRByQK4hysRe6OgpZUzCgkqrDckSAvMFqaunNOGvvl72lleck1C+M0dAlN8AJ0g0CycK5
NJpT96h2P7itMcC3u922ic4Jz4l3FnN6F51/O1GC5kllYM+Q6KIoeEd/nMESPkiRzW0zOw0g066m
VB8GMpTtuBeI0vxt+zCIvnv++OPtAoYU/TiPlm5QIsov/m3lJ06C3W4jt2Nvv33WWzXEF/ZQeN2X
oyGHcT5uyGcXQoKnXnXMKmqiix1w0DRDrd9jZPf7PgkQY88wrRtjQjZs/+lAvtUQyLUZKbY8cfra
KJ1S+d0ri+LEyTbFbitx6+xIMm1KMZPa5U1YaVuLlem8iS+vPxptI172dCjP+fCFAClGedXLFO+c
O9MM0sG2sitSkgRSgqTdldQrRRga97+zlV9SNWWW2r4y9//cwsBiJ56qS4YD613bzoTAHuwTeoOo
gHIK5/+dK+BGdaDxfE7P4uGG7EfWAcnxdMkV5OqgtoPKyCgLCi83bWQI/VHWW1mVUk7xIZ/y8swP
p2XPH3SlPZYogkdZCjHWuF6Myir8SFZkJs/1vayvo1kadwxK4XP0jykChJ9CdQtxQ5bff47RQLzI
+UVslcKdHYJ5Sf2ikeXcIQ7ptE8iSJBnbokCueg/XEEhvpS0U8pgVI+/7wEqAG9ojy+YwWOnd0if
+9SEgJbllOSJfKHJPSLEx1NjXXl1egTLYwLiqK0hwA3YRKH7RJVRbTWrcIO437abdz/YEzrOIXT4
M6xdY0usluzO50LFJ/nVcOoTy0HiUTB3H1UlvN2oQoQL84CCGAGILb7DjsfU3EkAlhyydjIVuMXB
T7iUUTQWgy4Mt4e+wmS7hOdQNV2A1IGgU1g9uoh0NeTdFBEkpprB9OG8FXIbRFjQf5WhNaiOMCPF
kR0Wz7HiWYlMYhv4O5wsXEyp0roEen3ylDrybvH8PgVUG8ANDcsDu0F5e2+9P8UAYDWhZTKe4APx
cBs0OMFhFeAJRhvDq5LbbbHE4Z4K7eudvxUJDLhwTKKFlMEmEkl5U8glnqAOtZNx/dU/MkxFGmgC
vDVMH0jLDtFW0WcsA6pevp7m485ta5oP94T7PVzPSMoTSUZl+SdLSsPp9qu/2bUGXiGsIW/mydnJ
I+DD2e2vsC/yz2QH18TjdnRUKqwBlLYjbEVNqL5g4EIGlby9YgcwV0jcr0Vv3ZrCfH2tXUE5ogDE
rHX8GIaj0iXdXdOX6vf+RYRl5RoqEZ97yzgVxwCegmmF5tcHhSebx5Q7WwTvWvhGf2w4TNtPAT5G
SPTeDoP15AXJyc8E02Gp5/DYHlAJY7O18yeVfP0OwCyeYvwPBxD+595zpEmE/4+JQv/HQ4XP2sHt
DWS1umhv7khsCAAOHyyxwnsjdAZ8OibKYOXVral8ryClzLI8JmNwXHIgF6Fl/OcULbWjykPgXTAK
W6ailSZrMXo/ygOXegSK8y55Hav9OgKdASgz2oN2U7zk7JxlB0f2bHZ9gzvA75dF2M6SMU+hvk53
r6PSdefKWMdrQQT33sWRIHikjCfmqLifILKKTpmERTGzztedpyWwRvRdbhj/50UMBU8uOigv+6of
nuFqRD++qxiuZ6Z/ZgxPedF+NsVchtN1c6mUFdHE/m4SjYMMIFiwzokq4aPD/ECSiOs4ywNqHpLL
6VlGewL1MgioGfSfDcRJIM9k32Y2HsoDE+kQhgJtnH8hBRx9n1IFWVl4AZm9dGyhFI23p5jXeaNL
Wco/MXJ3CcJIbW+GhvareexdvmtryvX8MsmKNVbCfW7Dsq0M+FE1CFoK2mC5Wqm0aKklFjBqRUf8
vRCMkCxC/0V/Q4jtcCyN3kMWVgE+xKz70Iih6ocO1pcNU6GcB0j5PxhRxQd4d7k4eVw4lsd8OAKS
FpuRtDBqyunZHfaH7THQMsUKYFRqhNnivUiukq2126Z1lf1n7Nn3NXzlcekCpKhi5mWdYOqJQhvG
MQjo71qYq+5hEORIlMJQEWsViCLiZ7VZ0kM8s29A5nRgAI2klUsJLyVZtDZRjp0QlTrugZIiA2Qi
HRw8MOX8EJ9i2hHMIdmisvZtXXjyMb95wPU2k+xoyWLvKGp2QDlwFHvaskfPqs0JWHco08iILQgE
tP9Ct7wl8Uj1X4ykobghGklgOPhvxB8TmAEuOs1Gy+yxdAJAth6WnDUCj9okewVhq5VHgaPxCftC
ryjMfYyJZhWARNOi7QGmKkDxEHCdKlxzTfx7oZKba1sHz4KNzk/2BKEkChlFprU7ZfodATguy62Y
dlUc1Vd+L92goyJkBah6N0TMbqbot7qp+m4bZge58QflUTVugDI/waj09W0dIpOji89aayYb22c6
OyFAgMq+E+9YHqh8Ii56CkJ4JI0QzmGJhRdcHUdy+jjVmFd5IlOvhFb+zTozokwRP946sV4MXFfi
xIzl9BsjIMrAaVOqfieMy4CVN/HA/YgbuwQXSz7LLwpml+mwTx7urxBbIuU658VbhbyOWHmHdjrV
C0tcMk9rygIcy/WEts+Y1vvPrOeiYtNGoy+2RtgUuBnwL2z/VIvTzaXsZv+GiMdnHsFhK8I/nTTu
FJCX/7FF18tOEhjG/ZtomYsdI1IbYhOwLEY6r8wAVkxoHMakO+ml4/iMvC2sT1n2wLh4gh3AnheD
SB5l76iv5+tYTSqoIMAe7ir5VvsGQ9iPEbvHE/qMmkPNOYurZEA0Yd55te1wGaD/COz68kJSXuSG
5V5cGc1zvkhv6Bl9I0bdsZ7t9jL0gMn9YojTYPyXrW7SHZkWFhg6doF66haxuA9t50r/TIRQUHLI
G0zfFrBB7XMDADQTruRE82qJ2c/QP7ZsHGPmhj4VFZPjturoF7ouzEccl7Mbs5U5geQoJAYtMYWz
SUkAt9wMGKfVgdEQ9A+QJAsJfsiQb+QKRZPxyzV++aRiCZh0Fqyqys7rT+oDdRjRdMlB7QHRmRPM
4I6J1gwmoKJZFimWk/2iydY5lDJJ1LqFvKJMSEygqt8Rt4OPw/RKlUkcwfRvqROFQ5SHv1kBh650
3RkNn3U0pL6P62LSnAdyPE4Yl9ik+O86YKD0xE4W8LEF9P2OkebR1yFjNMPDi6ZqjhEh71vnQHgI
+LJYYSCRUrSGEMUNn3p+AOHxCWTTjdrZVmoji7vPbl9fPOTUMgBsmMeMgGzOC5yJUggK5UpQu/wS
IZ2+vIeMBBWCYl1M1gODLHeT+qnnaGeCvVb9wzp/fol0Q0ahJbtXl3j1637wak8+tgX2IAAwmFbx
czElEKLIE+H2hiit7cEKq1RRE7Mc0KRFGns2xPI9HmclYfaZMtd+FYpqrd1Lue8Py1l7t3PlbXni
TWwbF8T4LrgG8Sd61A8V5qjvyRQrtY7V5S8OGT3edWkUW90LF0ShNr4HMeFpmoa8eKSuK3QfOu2m
Yye6ysq3QJA9GJNwxRCs5Mp6xmloXB6ED1hVakMk8E2evqCyyjTWxBcdpFJXwHkIJ00bZThcefCM
yll+ktNpNTtpFoxL6ivD7wgpJijzkzcfhDz547zMjGHeCz4hSr+LB9gv8GPyQqBxkFpOg453wmQT
XqPnudSMowCBwiVCiS2oP/3TSacHyfAHXmbs9LeqWNWmEboWUxHT+RSuCGJh8CiJn2//0qER+w9Z
70yZOioJrZEtUD8v8Jb8GnZCasD0OvKOU8UtQNXXg3av5UfgoLMCUyr8UKRcQ6qVhuN2VOKssS1/
jmeLn7kTT66W4d8IrrRsjoA03VlzW1HRrDkw3pi7RGEPUjREgmjQ9ZQzokM/310B1JIIqQhtMhcD
Rfl5cTc9yvVM9Y5nLDhv01YzgQDO9fibnNoCur+EYdetMRz9/Ce+O4FEwdDV9wRyFkY6t3VJN6uC
EuE6BqzO46MWasi8JevvZWbm2AWpcKih9Ln6ZAgptutyHU75b4ZcXMc6JVAGCU/apKIiVWeHQcU4
GYLofMPICCqLR/RMrGQ/lsFi5mOFhttz9FII4Nkjux+oV6do+NEeRiwdtdKTmDIvGKTtTlwe3fm4
xUgxg5nXNyTu7efNjCD+ytXcoPytcnOSh9B76wSuEyR3SkN66/a2TIFy3Q4EBKPLdK3R+Ir4lzoR
NKKudPg4BzzRL80/dtmzGN4c/kv00Oh+Jtj1QT5wfFYAMXU5Jmchs1ZZPm1oBCOv4YvibvWsVUgn
CteTnRGeUKgt9CqFbxsUVX4dtCJnOqPsSR0+XEugCOrb6MUfDJeoO18e67t1XLZDlFVLt20cWHqG
n/dd3EM6KXgAEoskqbUUTTU2ydtrazLZcWwps8q2cZDpyGjesJ/Gd3wDCpg9lvpe9Ghjbn6lRkbz
BrBXuKiTyesFac0//0rsfzvlgbyPENxw6r96d3MwelHWqW9z7Me6D7zMumB8YcDl1pG3GYLftC5s
9f1uh4g7MnyycrrapoyUfmyBhNsUgIHHNGxjf0BKJ6r4YIPBJc6rLnVYzn8amnbgaXHxt05HRt4Q
yQHQeMv+3VYv9qkaxsfSPErfLeGaUQJ7hNZpjBioGGXhPLLzWj8NeUpscbjsYkHGvFuwgYai9t7t
voZ0BsM0uwlQRDSC8MVkcJBB8nlfayw5fnWLTDnTRUyizXfaKMe+r+9moHI61KTC4EJg7+Q4/4TW
jQP5POo512Oq2lYjfiUroLDn8N21r2rYR0fOrLhm+hUhT4nPc9bOYgB2ltf47fhcOaz8RPzYM64r
F419AY8Vr6+l2hXDnykzK1J5PwBJW5BuNQxKiKGifzNh4zENC1OPfo+L+h6D/B1ifWP1Byj9Er+R
uDsfIQtssLGCtmSVDFdzRSvh49blGqUuLk3lDY7zMyS1I587/dmgoiaSjf0qZZM5Uunz+8LDQ6Uw
2CKZpAER61VRWZvhi4EAdQ/ZnPOLhh9zWCpfYvkdxFabtX3J7DPs7VNxQvKpJtMmUQN2jjZD4dJm
4Xw8heIZvhZ4O9J9S+0+QVcchWgZ5NbKBOmUNtgldPHPoxptWaUPOid6obciZ0ITBE/fd2pQ0zK1
wNGzcf/vid77+7VFailX95tcPEIwn3BB/yuo9ivLO0Ddk6Bo3QTrYEmwIIhxFwzXW2OEznPXANfP
wIMe6pUh2JbdwQVW+mbwIPjk7eoSCmA6MQ4eoO5IPV+SCP8944ceQtw2URKRhRwycHX5jpwCn453
jLv2CqeapvqOr5aoQyODPA+YFNJlPzbiTKEYt+pPEnDdYPTv93KyjEEPzUdJhjbnYVOFEUCpct8j
BUlAp7sQ55BLdnf0z97VzSD/Cd2v02vYo81a+ZkZQb0OXv5BgJcj+IAE7BH+2OT069OTSWD3n6mQ
/h3BHugoDNcjrcCIHWtUtnAGfVr0Nu/qEBslOAcci5xWdrUs1j55omRJcOIYz5uCcfS6lWstVTe8
jPiWH0w6vbavubSF9d7NI4e/atn7NbJy++yfkgXTIFcEIW91TgtlZPhhhHBz3g7XEKkRcdfJzM1N
RRE1zAHybwxiVJkbmPWGQpWtZIprqTkhXVxKTKbp+aHruDSDwEVAy4V06AouUf0QZzE3FfjJ8cvF
AqCzZqWv3579DplnxaH5ahNJYLnWfuHx19WlYRGFF0cKox9P2z8rqUBmBmTQ8aOnk69MLMqnOtgJ
rvu4KcXCGNl5QDtjRw6rHpewy9ebTWkxZsIa81w3ZP3ZNLr8iodWGhEFUADqOimRf9jTBb9HMYB5
nvCTIrYBZCCbGmYoIR6/lYLQQJUeShGuMiznosVirjHLbuAnA6fYmcJOIIPTOiAAfpCxFazqMlEW
h80eJ/0GPx6c6irne8hH8qg3AX5d7gp87FCl3LJes6tNfzdx7SDYcktet2b9G02wSwTfUFr2gp3r
cUMAb0RnXm7sbCgD+AALWMOvzHcMpeMw6r9gnQdfDK5aNm4DzcCDDV1NSrXskRsHnJkHKH3Ffdpb
rqT94LnDOlmSZ3sjA0mbwABWtlQghR4//St8/tJLVjt3CTFj9CyDoaAr8/FWUy2VrpfZQtKtmSLo
iwX1M41YrnSg42MQGybyJSOEVsBGhvwXzLpsTa+XNOc4rSMMxLClG+KpWhFU1Mq02OeAYz5S/Ixy
YJfsYAGynwip743+qMsUwIJi7mjFNG++HryBlBZBHuiJEOkh/9+PsUCDt/fWRSu1Al+uI1U7IDqF
jASxIi99zgq3/mY7G/6Iet022/iQluylFYeFpULPNcmgderUv2TOlTStNh0B2o+ilIPhm+ejCYO0
k//Qeaiz3VznsvpSkul377YcCTAdUEXbyoFkpFCTstY3wPT0emfF8E3oSrvw9yqTGMlGbIfunRCH
eTZz/oAI3tiEleH6A9rIxemYJSkiF4WJt8XhM2W4K1Z0XdtWof6I/wVYipUA1Zbn1g7twbdGbixU
Vkl7a1Edn2OO30/xEw7GctlBrufyzLoPyDsAsMHqlDxrig3nYevVCZpH2mK2PzDTjazxoMwoXquQ
wHNYPp/xK6QUJYMVt+QHMOmW/L6S1s8Kiqwtp+vqj0jPEjvAKF6VRIySrYXrazgrivFv9raKK0d4
BSjxhma+c/fWXXkMRz1AmcVUoszxeUIfeJ1ja8cor65kXJsJIRqdiKJZLVGwyWR1WYywwkqGEbcp
DtkFv5iXSkRAf326ijgo2efNfzqVsz2IRzeO8aLtIrgM/fqAQvq+o6pWKB9xqeSRx1nun3Rwmtzb
1r1xpUdiz1hJm7hN8s6BKo73O7QRGnQdDv2KbwuGYMlbOywCGKUW15GQw0uHeYtVTJAbqNih7V5j
WHL0V5DlLMxZmmBpqERfFlOVlVNX9AAJrcB1ruuXAGbQ3RhirjO0GZQ+ywJcImm6wa/1uvtTY4Gd
fOaB24yAKazOkX9xDOJBb0nVIfwMEY3Wdl3Kfxw5c3Rabt0qN1K+hfoiR5KR1myAGaRGN0tmXIe4
gsYTl7ETO4C8kK5+ru+nguvq08QiH12QLvQSsQ7CHEeJKGEWW6ni1vvqjbh9WNVS4IKvG/Gz2Uoq
RGbHNbabLgM5trWdX6M6CDgWTTbDNdtezRk0mqi+EpCfilcqCG8uuQ/8iO9YEyl607kgzD673WC9
Vsq6Zdh2v0ng5JhxtxkTFuo7n8GWqgSmPAwgSvcVqTt0c8WAyL4VeL2jpy2RgdUe9KP49P/felFp
yMo5orUb5CzlTB0ZwtfXGG+YwCgufTTIl64jYfXopVtnJDbm0t76fKoJ6UKRIX6T8sAfroDbL2/b
3qEy7XWioso5LtUFviyCyn7maAhtQZKgQAZ9uUkOH16XgACupw+7lGVkFL6ygOxO+Aa1mROQJwRs
bSN4q7Y4ycU8+Yts2A1gWwe9F/riGpCqHkBT+qEjdSHlZ2z9flwQfmFHWZY9hufCly+Sw9wlKdDH
GQYZjwjD9XEkYPKJha8A0ZdBQWtgYoYVOquRWCI9aoIfDAjCqJdBk5nUnaKNpCSQ3XEUzCQVcZCQ
SnXrA3dEsLpfLwtuE2MW9yR+uN19u9cBlzUfXuqrqLf+RzIwlFP2bkmpM0U4dLl0+69qC1mARoTx
JYg0PFINyVBRiK/i8v6GypiRvU214GeRJo6fL39alYTTtfBXFI01rVPl0S1PFTTIa/h5LPE/+g+H
lV3ZLB9KVjRKhuJwtDP15X71AxKcTxjhAuBHHlrEHb63ImS5BbSMEVXF4tmTyMs4GqQdjXbQX8Ta
eUNhi6H0iiBYnqJsS6MDVbSvvjwr2lMBTKK//R+rXs7ymOfZrGizu5c+1Mx4Gh2KecGuCmm9zLYO
sBjevcS5mVULIWWWJJhkBTFUdPlGCcBbeER+/VrX8HqA3vsemeCcpQWn1dRDnMQMVV1WKPsW9MuN
pJLCPcYG5Zf6d2Y3psXIL/Txos+UgnReqKkpro8Uv7Uj0gZCenObgpQJA4ca3HJ1VQDEZh0tqgyf
0IeCDfmnOxFEYpAQaP1877+cPRU3TlGYKhbA3VFk1jNzwJcyAde9+K/KVRGRsMgejIN84tkFrALB
1PtSlJKVC8VPUQrYH8qPZCozPOnJwicq0NsCLPKcIx+yD+SxXWeL0CuWHQxK0vQRRaimXniTa0JP
EteO3Zj2Jkb4iQdXJsMYRF1yrsHLO5PlDVhvdU1/8NXm2ZfqtrBonyLKW10COaRZVRIKuNssE6FQ
i4a+ooloyF8NXIwQw7X6ZZTytACSSwlEygDA8HjyScFOjxpccYmZt4r9Nq0RvXpDIx+pchbxtgFG
1vsj2cZcPRKXBuJO37Lllw24XGjRyRGSDvtaKL8Xg8mUnC+RN5Wt2OJao45tXOjiyDwoC5Z2qf/s
8vyAaEZP3chkTGcZYKgvuQGyVo9Z8d6PwiUSSTXrwYCr06w2RBSG+Zm1p8ljAYrbVUtQ1yGfbGkg
5cLRkGnR2yGIxvnAkf4WCnwXs25oafc0Qub/tnjfmJrITafT3T7suYU60U8hHuF1mLRxqK/W/uay
sIQvVaXXXR7k7jrdqTFvxffa2bl2541y+VjbOPjMNaWBasdAgMmc0KeeaeYdIbtoM98hi0kwQpq9
Saaf59U1R0n3JgZw0oYp3ZwQS89ZYDHH9X/lWNbQxL4tye4vtgWaGztF+YUk/i1Qxxke/oMYKerA
BimomBd7kN8tZkGU6smyUk2fjBGyXXQwX5ljE1OqmZAqBxsir5PvJIrz2y6KP0Y9nPMFaQwJKXVj
DiUDMWiKijRIO01Z2GdscRs7y0YzFvwnF7pS6VsX2E7u0M5aIZUD+gCJ1l9eDoqR0tdz7HJ4UH16
XqFeuWW0hzbf8gDHKyd0pWsQkYZ2KoHSwyE9qY6Lvn+nZCpD1mowUeuEM/EQUPFfW0H3gVsiX2Ii
J8URiUuTP/UPEJD2iJR579e8DJ1Utl6iyACtjRSxCOVQ43ngHSrzsusmWMyxoJnOhNLLOAFiZwE+
ZobqA3QzTf3jWRjN799vLUcMcJ48RMSTq5ug7Oe3inxwjF69fIo1Ie1y7dJkqwp9xGEziJi08oy2
utojrLo2KuM6QMhXhT9Ii6lyadP9HdNO5gtuWcFNbrOuEtHP2ws91D/IKFRKjq7M2yfU6V1XyqF9
tCRFzhp0TLGbIFs3wOSWA7zKcahhHW92sUc1IPQLbc5ehn/U7CoWY2fOru9JAsOOH/Ww+Ykm/Ibe
dqxxNtjpkyd6klCGVz72vNT1hp4P9qia2iT51Y1aKqU2Bp+kh6f2tPPH2C7BGsLe9z4ZDD7LNa6H
m2J/80olVhAeXzfErGhqR43L+Xt1JUMH3ZvQl8CJ7ORNIV1mlN/8iP9GT8S2B9HhpmFLhB4NRUBL
rAcYCAffsdrXKZdI/g7ii+FQ4EFlL60/50RaJLlng8uRI7vkVGWjuQ35BscfBjJBhBHjegVJNo28
C/VQv/q54nS0pOcaKDOlhjNt7gw6G/5SOs5ZKTded+a8QvAzjycb1kGOWi/w4gUjNOd+3Q1p0oLQ
+CLI8N/v0AGg80g201h1tXSGbXcPWknhWoFeha0kCCX+3Vopzf4biwXUUvexbit7evG6zQFbkyRb
Rls0GDVOkDJwkhoRduDb9hwmPTaTtpYUTP5xDa6w9CzHNR8u0AV155IRuV3gY11ESdcMArCmv5eT
gjNoEOfBBOoZOSpUIEKaemZEyv4qKczuPgA2d6L4SAqlxjl63kO68pBRpVHNOTv/i7/7qBVwJht7
piykyFaPw+ydvNg7JWxX+ct4WqeWk/kNFQoe/6YfcUvD4PhBPxlC2jfoxmdndeUqzu3rxDP16j4m
HNzkOJ1t0SFSAXb6cYhYLAot1xNs4NzoZ6SUnU0axAYELY6atcyvFeFUa9EV8rFGuCB4KVvlWyXK
biiNmOEelhdmocA9qmvFXUwCWulxlSrz3yGntovCsaoB4zKcyfw3p+scTwNg+LGa5fsgjEl4mrYM
46X9zEfsOFG9gYKJT8Spg/oEQ/0Gbm9IzM4+YDXKJcSsFlfe6pDvoYtyFR8LFMGEjOy0rMB99AKc
HPGyj6AQCwzWbMtRGfZxQzQl1/p/JJnyFxxcMiY9H52TeXmbvqCQSi3BiLMGrUHmOhjSUrm9FndP
n/rVo/mHBR/jNgXB37NHgNx5TeVX/gDu4T+c82EfCoLxkV40KlJdezMIRmAY9GZmaSdaID1M9fWl
bFRpqmmwkzyXRGw9d+TuK5e9v7O2y6mCNOm26Ol5kEa9uB0QvagaOI/WmbzB1fIze7S9ezHFtFRm
2H90OUIvNnmH7iSGoB936Po/J77jTujjD2+DlG1i/H6HO5NkZ7vhSr0jvsOw/pGdZsob/6W07Nzc
AbVo4pjO5fcwrVAcGFor8FF4nTG6Wn5q0EfIwiElY3SlpMQBlPwV8+rcnKEb56gm9ruuLDBkBQaG
/r1wWFfXA7Bwd3frH95m8OLhsnzHMnjAlVdB6f2HXDk7rOzBxsdErJJqkTjTevO5ZprwuEGSeSoA
nCUkgPotiS8poxRcOL9gf6rkXz+n5BxFGgSnVJ/MieunF3rAilj+nnsEHqc0Qxa2BCZh527J5WTK
GaVfe9cpRw34m11j/6Lpp7D9uNKmmvzFtB5wuuB7DgzV3iqNcIoS7etAoUusZ6lmsy5tjp1KGbDY
jv7Sbmykmj0B0N9JOqaNeNK+b/UEzR0YOFVOriBIpw3Ub91GJ2jJz18OkjOQQp1EeQN6fMETTThe
GayXY5T89NPagUpbLb4DgbT/CIHpjUpG3N5rosFeKhBzXRyXkNSbDbH2Y3ox2g3hNWIa4TcSw3aj
GVNx9iWkMbnUgsOCU26BbAzWU0yrFuXqD59/fJzWH6RzN1k+YV/2PLNEyLTeM1Fl3PE6z927Bm7/
PHL1AOK93+l9sGBH1TqvERrdC5lgfBR9VIddYAg3eaT4NB8W8hg2hCcfXB8arsOCSp090fHM3N1s
Jl4lA9d3+ZXhIQBV7Gq/xa2W+G5w61E/TBY85RY0yJKUBQs0qKoBph2jFWq2NMhd06tGuOziwSNN
p928Wx5XgSpmxAiXQMgpdw/IMlsH1UsgPLBMtjvkgTqoO1I4bC9KTuiHHLVwJlbzKzfv8QR6r+8U
9cqDHgJXLcFvrUDwLDYZ8GGunombQq680qnDi4iejzzyb3u5o/GeMCYyV5NIA2/OFIrIulzgAH3G
xb14m17KQ4CVroqUvRL+2pQ8Nqwp1NBuWi+JnOkohxsGSNUjtmQRzqZkR0kwk9cUB/zqRuVENsBi
Mi9u4/sU+4TI8tmDUxhFJ72dWa2jtHNt6F5atigimzB9Jl8YnujJicuEH5mhBwNzUnR4lw8i90yu
JdQoLEtZJi8V5tTS/H3t3Ti/QdlpvcGj1DeId03QFjya0omKA+DvbJLnhCBr25aBxOvIQnFMQCfk
g3GhRzmv9vq+r5ygulD1iByKQS83HQY+GRCIDhID1D12tvU80XOqhA7n6jmJV0x0K+QWdzWC+ooY
XmxTYEsAyR6EYq1XdxglhshDlkUgXw9oVz+/qSrCZs4Urm+v3qT8zgSrAgFhIm9WLVA021icaoFe
RNQoTZWmJUP8Vsg160ZGoKWgKz8RDysLclyd+KPZEuprBSsMLfYGhv+sCfqxjySaTv7ROGnwKTxQ
nzSw3GjMHVbEZ/VQtoZEznTZZJf+rQBz7KruMhH4f1AawAJMGf2esNnK2cYVzCTU39PkHdsNFOm4
gKSyuPY27Tjph+PgGIXom4yUfTdXlKLhtsMIP61si6OdfHwgEeMLO3UO10DPGAuNgxm2bccMg/Q8
0AkC5kYW2aSSY/bbfUtEKyH1s2j9gvzO4znEaVtbJM23X+4vf9vZgdwBUgD/7zkSAV5Gtzepnkp2
ssWd+RLfyEPOFd7SUBemcQWNddyXC6zYWCTVbkA5SN15bNnRUgqBJdGY9L0G9DDWVMfrPA2rKqE9
5gX/5NlZVxBLwL8kccwsgM5+AWPzNaDgq94rtezTHSTWx9vohQv7uPxJJPyXn753THfmGtGO25ZB
RUOJKj0fcLwCbfokgVxyUutk1Zl+6ARXtzTUbT+6aqkC7b0ODB7XH3R769oajrWwb+MGIzydCJxS
j4t5wt2CbjlV/sfoZm3F1TE7paTr9U6+DitAhgwkp6yXZtYySfwoCuHA/McBqhgyabgoihYs4C+R
mgpK9IHR98SsVh718JNT9TQL0lEiZNB/uo2X1YU9sK1XxCBjuXkiVmkaucXOk1c5uSqg6eE3T0zZ
F0YrsQHYxqQgWna9EOPn4MWqJ4hBOvHPL751tILZ9Jx9kEKPohqByjSFSqpVklYMliIsMCDDEf6Z
0k92sZUOUufbjfHUOk0k5r1OIkgr/jcyRvU6El9y30DYbIZ1yb8ZCZxNOJpn3kxbCeCWASEqnh4G
zAzey54LcCpxwa199NcQaikjXyLpqENmfyyrwV7EUsccSAlQzwgcz7gCBJOytZ0d8e06TWT9Qb2d
ZOruOvV8MD06TsRWwdl6qPs7ZT1sp7V66BbkvQfBBcmn60O6KH4CUjwmq8Ve4FLKb/kYCf1prHHH
75LiwQugd+tktdiTyxdjDt5yj9QXq5vFxB8cNXAg33qK1YQv4yeVrk0OW6JKFHzBB7Y0+7Tkow+p
5eORyEk03U2o2cKF6RD4vnP3ZGhIirEZrdc2k3kNyrosFteNkIcJr4supiiRjBghHW+pPRiLfKkl
Kow9Awc4T3qDPy1b/1kbYTHKPUJzCpJ7dgwXy09rMS60RV04S+JlKVNNAdQQB6MbUFZ516CnllIf
YoMQ3I/yNeDFDedHMOMEjRw3krtHgKfr5Sf2qgsL6PkxmbJwTKG6FYshvxj9E1qMN9STQfHTecAd
bTsMHS5tARYcRruvB8oJvkn3cmxkry+x8+1aHiaGxLwxQZ+5UQprhtK8MY6oFgMQXfpZtlMdAzgd
3XVztpsHjalqcAj2oxobF2Rnss4Gn7hs75IpXeGmVPeZF2c7V0rUNT7Zi1PtEjtnd/wHzKodbikB
8rJlGpCWT7+PEfWbrn6xfAGmCC8qkS8G2Pr+ZRmOl/sBkM8yS6xQjNBv+Y1KsHjWHa78L1P8uULo
QPQfIGe6CuBxyldByvjFIRR9Ep7fqYmwgObyiKHPIqeZXiEjmZGu0CjUrSI1UqNAx+G44ML7EIXJ
nPK9r3p0wHF1NfdmJMWfG6NaMVrF4qlP1uy365tlrgSOlw9YHeYWC+NeD/ZuU9LGARk9TCxchTJu
zeUn5ubhOLarayjVB9wp5cqSpvPNKFmY+sw47X9QgCspUTqocY2lrfD4x6+JJexziY27XYwV+q4c
LaPTXdNQTRk87/g2za/S7xY7ep4NxNBGUE9yUDWM6OmsKReteksAtEjDpI0AB8Hd+yY+WCersp4i
NTZtq4eJx2xANwNqVf19OGYlDGloalcF2Zf9wmcW9zY6gyFIqigSTvgmK5RCNEffKKQgHoaIKxrG
QgGvVJe+ulhViKZ1F4ZjONZnwMJw1IJLKyfp+Nk3rFEFU5WeSeS4JKnIdkTkNagaqY+NQUiqm10x
tXoP7rhwB3CyGowGO7rNgy6C3zkbTAbJGzL+qNW4fZNZpz6WaDTVsf/+Yezxot7M0MR+++PU1Vgt
uWM94RFl7HlWyNdSv0fSTo/Ri6mTc8ymFVUS0+nXmeb4DOJC0l23E74slB8BdWv1pfRcwlvGD8kt
W+5McHL2/2cuwPEXlX6iO9Xv9JOUjJ1gXD77TVljxXcqj+AIcILx3wxNOctBdACfRIbPAyfYk2cr
iMb23yv4rH6dJVz9a9BM5L7KhiH0q1hOnFSXg32rF74V05xOclo6+KRF6+Vuqw1WYx+D0y0Vw5H+
J0RxXwSP2ztggQG2hk3h3pHukq0dwyNrLiIH28I27n2guFLbaoPhChTENvQyN/TRI7ogv/bHe7Am
Rh7IlIMPPlzm+2aQPj+heW8uTIfJebnZKrCav4NKIR/H8QsfrgqeVuPIF+TAabIvZUvOonvRqRTW
QtTuVKafnIXNFnBlccg6Yum6MRYPnRwI1jKzKVpWbLSz3WEMJn9OGY6PUmHiRWgLLMlyx4ijOheK
2vtheMwmKUNsIrzGxgGgv4yINVxeKxw5259Y57W9rO2xNcRemawvBIAbxMeQQSCXnDFH/yam2Qbu
iXGHSMpP2JgcOR/NmvJD2sLheUej+Hdux45Y2RrQMBOwj0+P2lyFiocmQ9WjvTdmcek0UkYn7ssR
lBxlJ8XCIorp2sOnKaAnaqRRCrar13CSEnW03iP98EZfenqo8GHudW2LXjwCd010HS4G0K1Rfnpl
3hGwOIRPQX3ssdfgK8EhU+CSMDkplhPMzXO2NYlRVBEfCEmA2u2wFktI/Qv/BD+BJ2LK0NETMYQA
K8+h2YbNG56QTVhPhVvzJW1sljYnnkTpGU3cPTjc/Q5Mym8dTIBIgwPijEFIBPWVHt4r7e6yJ0MS
pS/WBMTmHdJ3ZIaIQc5I2GVA12UWTKxD75tGTdQu45dK800DrMtnHfAe1TtEVXQICeFUqRa/XEo6
ELOeth2yQMuATDD+IxftDxN1bJClIEYHdYabh5AcHig83gfmj/c/kGnLE9BtDQYZJHj0Z443kN6J
N0LItQS9OLMmQonG836YXRrBGravKNBxHC90JjC/KpZCilF49rNxSStNXThw2pmKK30KLmygedgL
cE5EQNp2JPzF1nhYs+y4p7A8Jq6u77QdwbXCxFqBbmgnqjdbOm+51jElxE+LX71rwsXIHSLPp1Kr
tWQIxssi4929pAWRGGI/yW4JKrgk0FqUaUSQfuzpyBcqO4UglF0dkKMSt2BCw+DvKJCrUCFJ0ydA
u5dVz26FtVO/nrEMAOKLbfxq3pnKhAUXjcG0FRFYTNfH9V8i9CoWNvVBxLf5y01xWfrHYj7qjEUT
VXzWtB2qG507iqcqj61OsbzuuJTWBSopReTwAAW9U0Mzfvb4vQB2kLZN6IRNfPUdlGtKlwPLMgUx
jzb7ljlisN8jN1W4YwjoGIjE9zZDunix+Co9KBwYYfpjD2Y097VEvX+lOUvhaqKSnA9aQNtx8zgu
7bZgHXsne90r75P9tvbOn2VtOyNY8jexA0mkDNUEjcC1mRrJ/YDJeytQR4Clpr4PgPjkboythaa+
WCI52K/yIFZUe3kSzMcZuS1e/7XzCi4/7GjknjUpbZPOxb3hIbSuL1YiPtUa5oWpmx3IFzdSmMGY
SpGJ9KAq0aRGFBh6bnLZl+BjVB7NkwLY1325hl/KN7WiHDABWOB0zYS8Skr/QvO5zJ+m1EEOezia
4dcitN/l54yIhJjzbc9iy8+b53SRTS/iyLYu+M9R/0EZezPByuU2iu/xJJBtLLpV7PTRNJUv27yN
wfcUcsBGb5d25Wu0F3OKl4ekFSLJ2CHTB2ltZt+UwP/jPNMnJAMOui0mf2JnwQuma300V2slnYr+
FmmAuYijl/dV3VVjC/QtfEHAQckGWxq05W/ZqOiZBMxHDMb8ykbbLpDKt+U1O7ThCsiPi2+j1wnm
emb3wkFko0XYnxehn/IPyIrXvkz069pu2GbRZEH5yferqZQHGILEpZ/zdZRT7rJ9Yxhc4G/O5Tca
zkJuqxF8kKFCnL+YPmfcy+Gb0caxgoX0n6HoJBxNLp5Z48QBYA5lrnu2kJSw9vat1/Q4ZJajdwRN
V45PbPJ0gRnaQUBGLdG89w4Bmq7ePgEeCjuFM81c3bBV3D1qzbu0iuO1rdIgKHGLq9MrF+0+mMF3
3gEKHPBQJ/ijTl3b3xUEgiIKPu4v6KT8VpMnaC8fZdZAMMlrDP5mkCXedPpcoOcOw+67tAOspjIw
kVUz2dzgCzW+RZvXdZngU6fy/crDyHSiwXWcuuJWUTY/s5INhC8tS0AIgxQJo+FP1Jhi3H4fWwNB
HdtnRFkrMx8m3xQsdgj+JLxQluzJTaljsc+jve2Bz9LowGjVjj3QLIU8yVGZJDxvpw3fDZeLEbCo
Jj2YCIfvJKorC5xD5igPIGEK0RqDBGDP0nNnUdXjpXgJo0ggas4d1DviGK6KJg+k60WZVVRIecpI
C1wzhp6tNQwy4t9mcitw/RQSs/fzJuo3z6YVj8kB6qk70SPrhZHEAyLIp3UB0MFkgmTB6o2HMRRj
DbLrKsTmpjJT7qc/L3plO7jNBqIU9PonjorvcxfH+VH+MbfsEfoZLOhIHrlLbqDranF+ycIs/eNf
f9OVuVImz7IDJoc0X/sC4ZMHiWYe4M9vebd6oMXlLLV6fBEhXu+sAOhaG3PpjhxBtGv7Mgk9ZcJJ
Z1pjIor9XfW5snBuHVYhakMebWLInfAj93hopZiQ1+1iJqekWNkNZsQ5zafLmviBRKCh2bArv8Lc
Xxs/LXFw8H5ntgsHCZB1FKzpvRRQL1F3ILmO9KQ6QES1WJallgWNeuSfaRKIA2yP5dsFuR7NycVS
rWqUuD+798VXms0A1XCSZP5gH5IyOIgbgQbZQByeM4rb14PqdnebHEjzG7kXSgseOHhdFu85XWcS
AeKE5ARSu60bTy0vWe0JMbJK2C4WdPHGA8HglRw4nWj217WaQCfRH0NSVn2uDkP3jbaSCf2HTP/P
BWxWl4Gx36JQkL64rX83CrEP5B9sqFfCm88m4xRDKqI4LSMH8TwBkrb0Q/xA2zhQvuP672IUOkzo
gQLOfMiWkD5nFboM5TPkNzeOJTVUozHuM3wj7Pu78uMr+CaUBpPjpSXIJqSaHNoB80HlkscNa5KK
Q1ja49v4gAJkFetFocnCA4+2Tp4z/3f87K7btRuABiYqfxZdcns2EO5eEqqL/qv86oplKxYALJKJ
UeTyvIJBqTNCVvCcuj2gRx6LhRz6ZWjrxM57BNv4MYfODxbOuRz6/mJPO9gXirZOG7aLRhzoek2I
D41/MS6tKHIl56whoPJLJsk1jbbmVgCbkHpl3aC1tqhfVKBMZ6aLZdqR7O2v3OpEULg6S3BXxmD0
/C5X+D6x1GgBjEsRJJGNi2vmYNGwZWgHV0S5oilaKCKL5nk1qeVXw9/f+eOllr2NNbWbDwleuwqc
M1QqSk4F/Y3EE4ij4mUdSET26MrAY6KjT+HKxGzYFocuHhquUnC1JZGfyaD18k3UAcIOoEAldrHK
MgvZDkxc9d3BzgKt05as9i0NMucCEN2uJBbLIqBOGz9+quHLBX4Pfv6itVETcYNoUwhvOmg7Hues
P93LxY9DRUhaQMe/bjdMehj7H8phyNmg4kiMuNxb0/5AwdWEkjTzR/lUkKr/wJI3N3y1Yu0Pwb5V
7rlV38WweZ3G6RmzAB7eiCQihZYvCb18Knk2dKpYqi5UGlSp3pbvvirlUIuT05tn0EOKsJUUJCqx
jC08eIlEE8dCxA5iHy3rxOIRQXLrij7eXYLqx0FTIzLEbHRBOKt5eArNE37Zp0POrh5AzzzxYeG8
deJk8sy6CE6+SSN2h1IU5UZshCO3LlTyHi6YphXj4KEtcWf1aWmXdzF2IAnE2peH4/fFaKqHlypm
jPRO0ymZQ7W25VsOytGwo25+tmz29QcTLThSwJ9zjNeku9tFz4UY2ghjCtrBbGTrthbOEPJi8huk
kkijoUa5dnWWOZE7v5zF9e2WsdJ9Y8BdIOhyBTwL47iiTw6aoEKb48IYdso8+oY6ET8Qj2vaMhsG
88AdYiYZp1PI1M6jZHeYQdk/+dtC0TXTJ5FsyImdqtON6fE+0GM15gdMyk89s/h/OUPhymYgoylR
qMAKoSB0KAXjg5/WgKS8HBtmFGc/B5lcNe15tlwtHzzm0GfViynEM+yBltyNHAw6o3A+ZIq6K3IS
NtSR3jpAJb0voqVrBZ5KVVRl0TGX/jZIeaO/Kyrk366ZvYYEa+z1oWnAPTa4q1Vua+gwhdLa99Qu
dukSWgvvHrBVzdwmf1RIcTFR5Ofg8aJibQxTBmT0aLwwwhJMGA+ZETxq4KPJZYApNYyWDu+65bNX
27dQ7aRPW9mG5s2G9PfYkfwN3+0dl82gm3bustpWKNzfUT0dtLPdGU5H7TbjpMLu5cywtLd61XMU
iOpZFCVx8cEVhi5eo2dytE3am7yNqc+eAJWo0U0GYFTgR7M3F316tj8aVrCGN6g6altNjVmvCH3U
UpLt6EZi3O2fhodZ1sXeHc7Vn+QEJGy4vDcLdExKMeCBmQsMK4sT7xYNrsXC/JKUdA7EqBIZFQK7
mKDQFcLkAHl/GFd5D8PAjmeSNqa7wHwVrC0LVkyC3LHcMB9EhYUMGp/rRtopiF3A3TlgQLW4EP1/
AbdjXXlMAjMHwmRHNfrMNY8wngKClczvI5+N2zu5Ntuqla/66d289ZTzKSyVF8Qh550EP2sUeYIE
dM2NB8XZ04mgEJotf4YAdGtNyXOGyNN0V+E4CUKkIR77B5fiQABsQ8K9w5XtbHXsfYUHKghNx+Lm
x5eCI0uNQL+MNus6HdzPMMQ8NRzVvGn4jqz/mjndMc56V3euZnfsK3A2S8FHZJpcG7L2ioE/0tyX
1WRbnXLfb2XluvF5LR7A4mrVn3U0xLzhVU1ZH9EEuDe0D5FCA9UqKyONY520ZKcvqbqlZYIbhrJI
WMVIND38cuwWu/X/S7Xg50+AcXvJ+98UwdxdRqlh8cgg5SFIaeTF0P2pWj50etvuYqmkFX4MdhYg
pEq647W3HSAgZ4SDXxiQpwODOse+W/p2i2ZbdrmHZGvJWP4iTMlRhy3ZNzqbEKWEMEXw/9i+BhXP
zoie4A//pJBsZ0xuUdZyoimPuxxsireQxRoSm0fYQ+YLSatSpHi4SNCc8Kjt0waCGuOj5BbN1pAC
p/3wtPSCaXIAKoL9WM2jMVLYl6ZtKZ+iY7wOmFz6ZGr++AqvZPU1an6wT1DH57ZadM90mKRKt4ZK
7hk38cvj22U28finQtRdIqqfuB1fTpV/Jj8obhcG9NMnlMVOFAPxVGW9K8ft8FpytN+z7g1EQ90/
Jl6JlP/yyzT6+scCVXf+3AaG8+TZMvUBYVJf1rllOhNPRw04Hn/sfpZftn0DDgsM+AyQdmAl1q8q
jDJbYejP8jc+uhfriwd5vwKsehtX8dEyYVkbBehj3mLowsxPvOvmXm4hPu7VVBPz5hDbWa8YatBC
O4MFursgBanN51SzZTF9lNU9p0TClVNSRmGYC4Q4yTFUuUHtzT2FFXBxS7fj5lPr9oYetNqjFY1Q
aos913hjyEnokjyJitusPqTNxBP0KnQcFyL+OSo5CjbDPaEt07FzMPntYnRVSU+xz+kq5p3gN4XM
57JYFyb1VJclCdboCkyA3RyjPzQaZSWlQODTl+7kIbsc3jYVPwvBX8re+CZSQPRdqiO/0wBP3sVs
O25HWevAfBMHzV15Pu0iVReHhhrHw4mbrBWv9IAnYJ5aNbtBb02azq1h4rAGjIo3tXQSXADCjcom
VRfcP2TOe2M/Xu4x81EG4O5Av/yEeU979zS+XBcpFT/tN1NRiAaxrL37vLlDcl59w6ulMRcnfVNg
ChX85e0hVdi8rRXTAtcBWxWg1VJ6u2BVrrveuL18pHkHEQg6XjPzIEizi8DvxSwD3Y/QTtmqN4db
fvCsaoHxUGrhN7yrb/5hZWhItYGcCxy9GA7LiZV2ut/93a7qIYhzbL9uZfWpIgGmruj+z/8ZhEdB
L7dZmVNBgbF6IxOBB/JgZcb/zyAdX+Ji9dC/Rw1DMmCk4Q37T1JvXiiC6p/5qb7+69vfxfEGsgkn
kTkajYyDhAt57PVHkNqN7sKBDWPFfbeRHHhevKNPlonLOJnjAIDZa3T2rbBWskgMu9fs9Uy5dL/8
75DF7FmZr2S133ROvjyH2oJKY/yXQ4k+TSg/4phjU+VS6muCffhUO52LUkuH6Hq3QJTpHWN+68YC
NRe924dlX2vYjUw8PBjEwWJhb4bjUaj5gv7P04sxfD9HYXq7GSGLpFDlwP7dCxmJuGmD9lHcu6SV
QujItm6ywaZa+KXl1KFpcvywZxFh8pXAjBCBkec2pszFw0cBggqp75uPR1sj13VgTGt01kDu7n47
1M+Koci/2iojcArpAtm6lpevaA1HaFWonEzx9Oi2ta2dnvi3uLntcizP4A+lg1OS3eU2/SV/DUHr
rCgI5+6mwY1WuW6zC0UkLnE6nKVSf9UXFzuxR4rrplFqCUVVXGLsDYH0I4qVrW9WGa8zq1rt2NTr
TSA1mbaMd0jCX7o8lb95TI0c60B4uiUSSpiX0qxJSqbu8Osx0fGyI8O9g1JQUXZ2Ir6v/MKhgf0i
Y23jf85WTiqBQHqOSWy2QQF3xnVsj4Yui2KL/YbRKYaUONteGS0pcSVlaruayDESJ6BPXIxeIlMG
i2IBKZp70TwDTsqD1pisFjZinf73zlk+LChAvydsra9Pcji1m4nzkD5QMfArcCiNlZrNAefxYKlJ
t6OVUkaVfSq2r8dHniz8cFw481Y7PDjljIkXjGRm2qShuBXM2LchrifCnWVWIEO6wb4leNAz3o1O
XclXYRyRxZhUR5cxxq13y2icE6nS4nfAulP7POAIcF9521+GjMc1AUpWbccezyJZzjXTEmZ0O/vL
Go1EoaVwLLPtHLNLAq/+iiNdjLClxy/ug7hPIsZ9GIfv2LdSawuMe4ydZ9nyDig3g11vBTwkM3y9
LdmSbeAoQ1zJcUUbalBKDRBI6hGm081GC0Uki/f9T7RNhFw0LJBg7OnrwG307iXZdA1QYNjcXQ8V
+gWyYBMOVP3Z+gG7dNrgpZBUxhxmwg0EbQqJsJvkkoyA4a+VsDromFE9uZ9SahoPr4uO/u+nLU0r
WK8fHdjvRCRaMxzLVocDKTIR0fh0/3aEew93S+SatoTW8y+VY/M2yf7vtIduyC8yStHlld1OF5Bc
SozbfxwFOmwTAwmu3J4iKpaOpbhWgZaafjI05ok2pTbwuyCrvhxdFbL0OCxbKQ1tjAW5V1MRrHuL
CD6BfbtFz0Qn163//DXBzZKf0qcPI2mePQeMgwjxmxPMZTRVJYDK72WwCSWMY+o1sf9WO6QUwu51
oOU3GFC0A6g2Ms/O7fs9R5Bnhokk8mGXFfFey20LqjHPA3opFEGlh2/OYMtiS1GAyq5i658zDSZa
hszNhYMFa5/J82UdYuk7MrKlt9HrL55z2FUClAG0uVFDEIW7uPe3ByEF3OP1JRE9uUpdZWFAVBVI
Z/6XLIg5VP7/dMpexowSuXpI7L+ztSaDohk3QXX8md4Rh5Wtw9/IxH68RGKaR3Blc3KEA7uvsIpn
1+0cfOe6okm6d+74hExLoeKtxObfah56F6hc/PWOawxPOwvRhSjnn1o5EX/hIKYYp4AiAe1fhAz/
p/ckKpEtdrP5rGvkSKe76EuspbYiSRWlex9Oicy8KUQjaSX41vNaNlq4D2WkC4t540VYOQ31jBzN
L5Nfi7PxK7OF17f6AAlCfiswS46di5VeAV+ZG+o+a2AqPbe+ymtmy/F9OYd1xwhzTgXar9LBKCWo
JaLKCMX8JNWQcNHNPuqU8CdZ+N2mXYzI+U0tFFhACXW4pBVsKdLkVLoNgLxxB2oJBKBntg8DiMom
ZS0q4+sa24Zbj+f/7BSVPWD7hYQaQMSnqS1uO/JmfUunKVxwsswZWhKkY3sKwssVGTBt6w8CihAF
d2uli2ySJVU9zsD6gvEBsxYBYEnEQCU1NO25rf7JTPt/As/BNZ5yZTg+1piKNc2c7oXbSQzwstJG
FWQrYgMRCSyzk9xJ16QIpReytMlGP0b4SvpdqcWcWH2bVwTNu3E71IHaahydJu3gRg7laluK/Pn7
mJB2lpnj3IeN4zJAu2vqCfIu4TSfddnI3nlZO3T5FUj7zAiabs2Qj8oT5lCyP0mHtBdCvzRfmn+v
RV8xGfOyNKIOWMUf4iNBTBT3WTXDlu/S2jM3olHilMezzr5uwJXbndWF20mX67NHiZteqQYuJw05
iQrflseludtDvJ165T/5iW61Jg9396PP/5+rO83XNMKTMqbf41BEqH4hfB9VrBigMWcZ4WQfVtjY
qpCMqAWZK7YldOedEacb8w3+E8DExS6yPYDf2MAKI+J5hf+PMDJBc+YWnmaeIRJ7+V7IbnRzEeu1
PSWnKlxpqFtg7+TCp2koEUf9SPUE/hu0JRzpd3AWg7SpPpZX1RJGq7GkcuN7gRmdiAlGTq/qDqz3
D1CPK6Eb3+y5uSEOGINn8Y6RaaZqk0RDTd9vAr+ZnEzGJ6p2/4VP2qqOOvRhKNm71ixZIcXgW9Jv
TW70NGmmnk79evXc0VdhXwDlWv8IWUrLZSLDLN+xFHIl74AjPXEfTZv+x00UDxgJdPNayUVbVPjH
Gvg9/XIb1Ucg02pKKA442/T6YFypoxynjtZ3diKY+otYfbdiNyXDwkNrOX2JlFAYTzjdXjtBN1V6
XtlXqrSojnfWyuUaM1/2Sxz/TCcHl/dnkrJHZsKz5O8pzr5+cOdnTjs75cFi/QYikBS4G1xbxdvN
AxTpWpN0XxhjbSWsoZm83xUwSHqf6+Od+i8BkEwGA5OpasarsREXiISVNxiOEMbWsOZPkNz1MlbM
r68YB6KbrjknpSg6QR6l+FbD48VvOX61JpI8X0NH8etTfY4FJOiFlXnwzjqTIcob1z6aK4+fDyZV
vJGc+JKPYdRm8BvKbGYILsWP0YGNVAQc0xr/qyywbxIkcfpO1wcmLW8hUmH0Uhy1aw2NzAVxYRDa
bnzjzj387OWhIwshinhb3gZzC3zEK00sPIXQo8TjMVD+G4lf+OxGM8bRJhaF75z48NVKwcZ6vux5
9Q8MHkFR4emvfMV3bP4N1XOzXC+SmZg75n61kU9FFglN/j6SXC35lwGPdOtqab21oV5Zi8PyZNsh
iftk4Or3xsOQgqeEXNMcXj+ite1hMZbduj25rIjaD84FhK3gOH6QU8sljkvfxFCKm8Lg7b2VqPVI
iUGPJxmO+VZlG3EdebBkF479EvdDn2mVCVMw0xzLHEcZ2+IFTrmOSBYlDqv3Qea0myLQzEZZo1cQ
BLJLh3rKF0LkR5p+8ZmQGLHKUx483YSGqlof8p7LG8Qx+lciYpxh2lOItKv9ordZF6KuPK+PE1HG
/dISpFXn+WAbSnDEzYcPSSCJeRmjLBzBiT3FWcgmopZl3GfZiLew1gvlG1tAeUsKoUiZ7oSrjT2H
JOqe9q8lR1kOs/ysgATeNhgsRqWO0dXiwV+KI1oMs/dbGb5mb1eQ4lHFxpkQ+dHfxz4EdzdKG2JG
+6sSdDuDSMq9OYq/WiWQy7iivsCiPeYwRpzx6GLonIZEL4p8m4FWgL6YJnehhwYmvd3puoaXs81l
0sQExWq9Q5wo91OkS/bNsPd7iHYG7pIN1m3gBAMah9bI6yma0e7M4akU/nH7FAtnyMx7Xvoqt96A
0tJNayVYg6GoHpFX2xNl9A9GiYQwpNlqlUvlcnXT8l+HEYX1Z5AV0pku3H1j/FcjvfHF/zyFB+AY
SBlGmmvu219mrJZwCC3SGWz3ZQ8k5mdzvtgGM3byOk4iY3d2W/R28tSWry3UQbsV6uChoILjVVGM
KOFhULLo9hOnrX2VMtvtQIM0Gg0EK/WunIz+xgKaFnQCUy8ZWkFfD0ixgRAEHWXIu+b6XgzCBI1U
uqri3uy0f7EM5FMWDseKDAtZW5r2k0p/0CVdSnwza5v+BayNvYsudBc9Dk0C/T7z5ZIIcm75BNHE
AUEw0nbhqm7/cUauQGuLjYj0lkQXHmuuUc0v7QIRrJNSOUOaZD8IR+yY0ehzncNWkD9RpZbXJ1mI
ZXvJ7cVkMoaN9G6etMeZjnawLV7NEY77PovQXyQ0QA3E7Rmbt8LrFayGztADrGPABwcc7apaQwe2
l0cvWwSS16tkdWFJeVFwNpAlBNLkvSt1At1m+NTt8N9BFHzY0Z9MA/Ybb70/u7FdkwWOuRHz0tcd
DM05daCG3zCue0Zj1COHrv3weKpNBlZVTLgEr99VGPRNAa6yG2HA2L2xtbZxjhGtEw7oaV69PJ+j
vHi5HUup2l7A07XiQO0i3I+rfC1DR5oRXbfeB2itAvQrIN3WYHJTdsHEFT7AupIjRVkg/7Lgu7+b
HA/uc1nmTO29ZmVcpXfBfbLggFeT9E2OYusS457XhEKfk5mrTkLooY7Nsqa4ZF9058DEFXqiUqaB
mwUyjN4Uohef0EF6AbpPfv6hmNsPqjFZzM4WC9DsGwEUrVvOYCXddu21RSVAqSqbBASU0yAt9mHO
wo3tWdU/Vr0pxnbC0mTy5u01BO9et/VCk9PC0hM4dyUtkXYA0EbDjKgBAG+wdJ4KHOIe+6ellyxW
VVLf4HntP4sLkNNWZXxOAQvA8K1l4rGIJuCx2+8BraiY3U1EPigrvwjdeuX/GJwyNgiEsaR1hBXH
g7x1VDcX3RebVAb2ijMaWoG2xpcKEeginujhBg3ecHRAeDwOEVz/dE737AQfuub2nH4o0dM2onxD
BYH5ys6vR2O+whb/VLHLKE9Y+c4PYhg0Sdk0rh3qeKLfFpaypPaNfvjbLlseckoUMUoL1ZXCsjL4
DwQRWIr06L/bgk9cRBxSEurK8BZKpqPxLy2JBe2NL1R3zKFAbkXvI6K4ovrlOS5hQupV6v4pdlA6
P5lh3iLKu7RZXPcUpxPYAyTdYraauM//atNiMg1/NqrzrdsQgEPcRsQP7WVzuI94VuFM2JZGVLgi
QJOL4otIvFsxdpepzWMORXZvUz8FuvXjNSJ0639YHsAIrWdeEbXBc5XnUpqzQ/C117qCwQcP5d74
6wDPM2rGlStrhsrGtI/i/LKh8OyIdRkilE2AsjUKVEaG7Yr7wsMk5jZBB+FsKsMxKBSSBHb8ggc6
wnjHFOl7PZN98kkOBBgthZMhA/L00Exm3hiGfZoUBjnLGQzkb2uWcnQAZAPALLzGy6clA+YMdOc6
xcTS2TcVYvUnzWSGNovgQWp5djMzbO5jOPR/JLYkfMSBn6hf+XaGTjsEqIW7guSf+mrOZJqbzkAR
v3rdh9yZSsuJRQDrGhEXWesJ8JC4EeCHcPZvbBsbb77QFnO1RQ0bb8nbff3WZeMh6CkAPEJLvOD/
I3/0xnSuDoE5s85AXDevwlAxQIn6dKuwz3H28hft4GGEm556GgU8rDM/G3roDKlYalGWOngiIyii
IdRjdhckl5VKqh6jUp1UGaIuiGXDeBb2bE4oK0dno6S4v+0UKavQaUBNa0EfsAMDiALb3XRJeh6G
BLn7PP9DjIweakrBATXV3rgo0cm7TkNLLYrQ0W/+xoY9584Kx4UCRGdfTamNM5zhL4IVTyspOGIA
XS7kampGrA2c96AvLEMDcl5QqxH2JBwXNxvg3RBzL/6kN09ZK4o1jNrvLafsRzumJ3uS6/nU7NlF
eTXxGHosjhSCtta6zY1/PQesQfMRBYsHJRuRm8ReI6kOYRylhL3mclJmwaffVeVTegI6Tya5oFBG
vV6AhyN/MCQoNsCOlLgq+S8O4Q0rUdvJgHlowumg8T5Qbfus8/u1BxfDhvA6jfnJtGZfiZkqm7Nf
/imooemHZ/blyH+aNFR5yGSvMx4CFiZ874Z86f0wp+Q8VdjawAYhBq3hVGzqApjT+RaKvN6mGly1
w2sT8fHiK4pU85YunjN+xvtMEDCrXRZFdTlaeGOp456fS/kD8Ru3YVIhpZ9sJpJT8VPUTEkrCKEB
wcXx15lLOZFGDRNDjX1l0/cYWd8veDg+drZ8RIHDQ+Bus6/TnCr+2FoR6nWOO+CL95gKB8gRh7I7
aKEZtEY/vlbI3Vrb4cJS0c3bS6QyRLLvKmr4zUIutbGtc3kFU7cXC/kQSgnJiva//03gLz0KQQ2e
E5Ry3/uU687ScFFV2mwdXh3CyJ2I/zlytDsaKQvpbw5+9ECpxoSEyBs0GBhwTA+3D+0dX7yps4Vu
nrlK9UZbIg94cqKEshvVQZ+LLlJ7SQLkvE9c2/StSB16fe5ifkqEZBS6FNOrQfUTcPjZUawgKneS
EOlE64fBtBLFK1buiBSOsmJcHTXI55Ev0+kirrE5kFDrosY6ABM57FyFHal4Rair6zEoILLXkcob
QJ5ZYa7DiH/yWFwK/2O0mNUaerXGBxezIjohYJBa20UYl8HFt4rKlsbsTGx4zM+ICkG61h3fHYW7
y7+W6Gak9pDN9aR/d8o50Xn8wAVfazhh4cZWqg9imvSzydJM9ebDdb9OeoGCzFWphmmqFZKI5BDh
38QB4sH7tZzmyoiTj5p7kZ79Sh8kBjLdgkY9Yzp3qc2xe2GSX0HvYTOpaVYudYcLtxPAS0B8UTFE
/sDTYpFbwylkFfZZaqJtxFR88XJtHK4tGtMDcMpfQBMIJ+1dFxppGPgZUzvxvqh5f9lyEctPyM8w
VmDAwbOpXuElQOnCel4rCoSVHbEPAp05W6XWHMtZi2XmJPV98eu+3lphTiTpZBXrmnbOuP/l74iG
QpYKom5hUfdbBO1kJ7bUTovfcsFwj1Yf0IuAeuaCaLqaoZPT065MWgj8TyPR8y+cVV/G41eJ/hzN
xkQiFhT3h2oA0XwRhQvAThOis2M/SxtLqP2TO4OLFxLVkQgoXye2sLkBQ7K5RiFKdW/WkJLQctaE
Y3GwTegU/csf5guUsbEMthaQ1Ku4tbLP+thAShD7AvubZE4p7kD4Q+/5/enaoFIN0ol7d9O/68p1
KbDwpoUobYuEt1r8U6DFXyHEK/LeYwWI0HajzWNS6LQHWEbveuyHKyLfOZBSkA7bxD/erF1RB913
RIJdYwM1xZiIIHroS0jbpRTcITWqLyHmROVmPewPvfTbIMzbRU59M3PlN/RhWC9g3pYoAT8iuGDo
Yvj/8oUV4RQIDHD2W/O2x4fhgmkIgIlJMGxiVuMWdBRaEFhkxAeBojx/TdBuwIduMCXD/hE4NISp
yN78Tq6NOD3OYEqyf1xTNUDj3RmVM7zfA6BHO3lXkynumuWWNvyHwYespLQMg1oley41x/d45GMk
XanKwGlIIwKSkY8Ts23fKZi3fJzymmHCLr4nY20RtBtvU9+6Afn8Dj10m/f92tVVkLJ70ql9QSYu
lIQXKI6pgOH2yCwKOAeWsYjAl+1+WWRGgHX+oy+eqCfUKi6N3ZUXjBKsRlOIMPkyZiD0PlVTpCCg
eTh95rZjOGem01POwNmQlWa0FN2S6r1AENnhBN9Rx5ZMFCv5e+TN0tI8LFeElbu9yipeVmV9BKIk
C1JqL7FkngwPbWKqS8DhXsZ+Ag+ctFmOBvZMvCOmmumhuRTuvKtnFcI3rQPxBUTvOg3NV2yDWA42
i3vJwE1k1D5NkQ6WxYrxbwq2i/xMS8uV3x7sia5KzSWvR4YLUrTNquwAgHDglYjSxZqB3mxRnEgK
/WmfA1xT+dq+0pJe8XKg/IhcqZU2sLJifXQTggeV/AEZwFi9jptHCokuGIAZ4Pkobknu2jGILjQt
/cVDoefmjbJN5JU4yyJHiYPGze6OVCdg41NXZ/2DSojEURCay/eXrtcS37D5WQHZLEUWLP/mifS2
pnjmWggttSh4/yH85gVJwV8x8y6+fCPaFyqDjYaIXfsuuuZQwgryTlTrOkamhP5kk5REIZd2ROpH
pdp64Ik+xZ3VbTU+Z+QNyTDg+gIjAyh1GcI+TnQFhKtvu2RqC1hSKn4MyLgudg2H864FBBokMOpx
vp0FAO0niaGJ27TcUhCbwtf8WI6fwZ2DpXT5TI7wxSKHY/W79Qst5yRDUdxoKGKvRfFwVUL1YadF
BP6giEP4pozG2ulEP0scYD5rvHBkIu5mp+0C7tPiC6y0CC0UVeSJIxTzZMfjVJ9vUC1w5BNXK3fi
TdMbdNUiY9kApMAYOItNhWXyT2+6Tfy+ETBBm8uhTF7gdHrmYwJLHB1WOKGubOOIuNoOWUNbq17s
CvV9koI8nE8vdAXue6ETP5QihKc7bTpu90hVJ6F9yCxUtLC5K+vPgsWo0coO1yVBUSjFzyOQGB6/
l3uF7wKn7vabV8yRlGazks7Rt40QxOwber0duxSdlMq0RagR+z61TiU9vNV3lwk5xW4Pr/eNci9Z
pGtTCPYhVg5gNPw6tzu/gqrrTkrbxfB8GNl3XCjGoqj3nN+zzA4UwGtaUrnxjkJav0BjBSMLmWda
yvmgh3oRE8jaPopcIivldHii5ViTnuvQ4xq6ywpbTKfBrhnI4lvFsqYIQOtFj+/RQzsJdNaeFuo7
OMpBo8+d6GPVjDpc54V+jV012l5pPN3Yd/2CBEhYcx4D6AXEnSRUO+A7E/or7wrfE3YNylWkOXqJ
ZFHZ3gvROS8opgCLoqML0RhisEPc0TGU0Z8iEf8k/5jy+aaFys2vJS6eWrbxKiKbHqmDETtsuG7V
GETMZIg9OV9c25vf8z3Ap8QURr9s2tSD+NkkrH2jfivLGCQVcpjU1UwUCqfyXH96HueDEEY+Ooyw
axV9HuW41SEFz/QWKiINFAdDP/3VHiqXoeVt3QLVHS9s1ZwOkrPGg5OyBZazEflgP0BV6Z6RCk+9
/MtjMFp5yreRYSOXWDOe9Tp1P96gQexdo/yYiUs/X80HpQOiFnM+JurpwxyqbvbocL5S7ejxIR+A
D99+g9ssH40qxCnJRGgwK9qs2BQkZo8rNCJFJoFmB9KBfVpZq1Mc7lNccDFTG72Oxl9DPTgrrRTN
k8yNFdijBMoTEnrMaS7cXmoJek/4UvJkg2Tl6vzM5iWpzhqF+NIzYDkpR2kNT+HUYKinRXTC/2DE
YPGIkw13zAOvv/2K5RChydMmGSi3Pw+cJwo1TpGL9EwtFDMe05wP2dpTrxajjBROJ1APxQVR0LO4
0j00y60rAAN9LglEsIDPIu/pWIxpjTgZBw/F05jZShqRwccQbmmmBmGx+7gkEXQjvCG031EDBYCa
2t5sUzgD0qOO25KDbf9QPukGgKdenfMu0RTd73XNolGEcJjZJqOqVRkdG6g4g8wvDmqK7jWJaCdI
nP5PAW8Nr86C9bEHrjfUjZKhlm9t9Ob/nzSQ1qB4EF17V0z6hf9/Mg1WTdhnDLy8t0sdaXCOnlKR
QyF8/qf8cP6hS2c0ONEzET02cZjHV7+7oEWSzzgdbGxhLLdf5iRwlz2UJaFvwoDpGqxVRPhAp3rz
PWtzYgKo1tylb48cTyoYFkJhoRwTeNj36QrUiWZhMMYjqKvC4pMaqYB3g60R4jMG9mZxbTu2oGii
UfpFjtdrODcjdoYg8fhb8nb4Nrv1JYbQ2Gyjbl8edZ1kjEhZRv+8riEWamFx9+939Xw+OYzX4WXN
ko09Cvokyja3QE3FVsUkdqxPKjofNzHGJZXAGfLPg6pSxsJsnbFqefzniWY2IdG0EBN4N4J/z3ju
34Lexl3JXZfqgmeYoISxh5qo48T1fsUdCK8pjgIU2rQZDUEcdwuvH8CqxSS3OFTLU6QCqiHeFW+j
3t6cZmmPwHTyhray27TnIgSgWwkvIp3qGo8jNY16ivUsJTfjjflIuihPpjUxwAta8hd+accfDnyd
RTt0/TjrO45eUoOOUazllKVcCiwCxA+jq9meEzWp9As8TsxiEJSbwvGzC7nkbtfmDGRb9+eqOrpk
FT+AUqqsKzFcLck8cNEfSu0scA5HgNf8+am1QR5V4qneQ6uO1FT2434FB6S5Ei51in/3CKGW4+i1
X2beKdV/Adc4oPL6SPXXBhO4lRdvUdvWRSeQmnXDYnNZOUnP/8ofLBsDwVwxlYgf+SI9n037aJBt
hzjDQtlTwC+qKSpEzA6b242hplbe0q0jjJI4oW4yQnG8GlxO9ayPLS8gltHBtkC6wry8Y6EWWCRB
c/etmpgneVEA/s1/t2jo7jgTlOoPdwMFp72VMuDTZGyrhdoA2TNZVylgHEgI9ZE0xiBOSKU9LoNi
1GZkBdW8dBh/0Neh9G+8LaWSmkKCb44E8fZe5maXQpMn7AiVMyMlSxU0Q7DSA5K046CIA5LTeHh4
jd93HEYkQtSoGbBjFs4OgMK+UA6rnimdGVuhZrzNud9ZHrthLjHLMAAVkyBK9YT/2OsaLLUkbBTm
dhwizSG77DtbCDcuDGzIz/rr3m/cn7M+vicdQEyvQJJ+iKwCQxHukmu9IY+c70TCVYhhdvOvNr/6
GhSDiRrNdN0ugxAP5EBbLNwJFGm2CPD5sksCd+MtMDIreWiTlFen31qYc09ABfwa0PIpw7ivZZEz
KVxjNbDdkEwIRd5nfXiOcipA7w7wVfGrJmSxZAw5jQOJqL08dgYtCNXw5VlORz/uiiacwrpOg/XS
QWb47kQiQzWQ6me0gAawYoZSpKVV4f0FSPZytNtsU7agohvR+pkrwUeR1QgXauq3QZzqtRsE8ZSb
zuTfOU5OK50FVueJTKBNvgU4iVvoimwsBG23dOBuCi1l/+r6iYU6dVDKa+xSmaRY4d3Wb+QXGJQN
0b2hYsznPXJySL9wOtE9HzfxwdxZNQU/9r3VDPjkvhVvPjTlSvqBT4HndfXW1KnG2ym/hJWm0Ta6
kEroQZvtebw3UjdsC8Fpyb+TKz/hBr8g/LUsTdaw5tSgJP+s0Qizu7+2XiSNdbgO5c5JM2GgCl2Z
W5gbounZtQ6iWZ53Yv7q4xqfVbFndWGFYJ+T77fAl/y35wYbR3hiPycWrzH+Ivc3S+VgAk00LChk
3Y3J0jewCuEVs3ORhLWUNZGG/ICZerZ+KS8gJFxBYT+3cSI8zPPoooO2Fhf/6ZOd6+v7PHnwD7+L
hbuaNt/wgHWLh4yePQ+CUc6ExX15h7HqJzRSRUdYWQV3pbDbhilRz/IB58CBgGPPz4ZVWIwyHaL4
QupNtuIYwXqmzmEWje/rZuLBklW7m5JDs/7cCRPrvxnlg6LOrFcS8RqfZkNzIfP7+rsuiHtNeVG9
zOPHCGBjgJRRjjbVcX4bho86XWGrhY40IZg4e/cq0BwiNu5KvXQ1tSIxumaE4IZV8LY0+xkUx0iO
CqT2srdLSBK5lLancwBxgSVUeFQMdKrbXZ1ij0uu7dAURzlMn8ViPUbwNL7cYgN55SIFixii06Xh
cNSDSc+v/Fsx57boJstLdjNPzvJPXgZvHUfLoudSx17LmY97TRmxDJ/RnptXM+Bm/ee+hxLri5Ot
cJ/RM57bJY5MK5ek48GTHLZlEihcbLVkh+6jQStIxJHFIRJBmygtLf6oSP5/eu60lCq/v2VY63eC
M67+ocRMNGKsTQ7h6OdqKBkQAPGErzotsH9njezL+G4H5CqIKefGFsKrMMtAvShdEPGWQpWbf0/4
6fmh+4FtKs4C2YRvrIFWTDoy/nKhVJKT0ffSScF+NuKR48MFFTu1uumcKfWPkbdCyq7EjT3qROYD
HnIwLvxcYA/NxfeIg3IfzC6FpDB3Ivry1gAnFMB/qeJQwvypglkRFvx2DsrTMscnNjuZYH6BsSEZ
+H0tlKngWijN2VZia2Strldo0rozd8cpEvhZjeg6UMs/eUb4VEsDIiwTm/ESb0BRXt9ZBBupI166
bzL0/p6EsymyAoc0NnP6p4LtR00Wp8/vmARpS/NTllO/2ajjCXsb2mPnZMkiidBTGPYecPA0Z0uQ
GGimFVYbsLWnJCCxCbf5ABXTNsxINMU6h8pjB5mdtajPOZrTm40jxCIDZYfaP0G7HW74UB9mo73W
ooaMix3e87PEhavVP9/L0aBLAPrfxEeWIXIyTNBaSS+JjuIsrDMP+KL6IOMsoLPWmZRKFNe16D/K
/ge+wDD0+wHc+lBdIdL2k66zfiTpQMFdE/iou6lnj7uaSQ2pkq+c2FyJqyth5OKk6LoDU21MtIbA
zqcA58D4e7bkCHcvrjSw7tTRwdFyqGEkLYul69zVMYaLhAHhny6OXgNyHYBxLGR/fRHIziUwzAzT
MGgh009wGL9AoIiK3tLrcQQ70NGrLXN6o1/4BuVqEwpOdO6FC++hKoCn6qJFAroIVjSJtWyoZ3nR
sSOvPDUKouynsdQ1G5DaetTtz+C0aW39SbgSUuPjN9L2KthLZ/+w4AEwslnU/Y3w6NIY1ebtOUgO
eK+faXBbFvTLDpU83dNuhzJAQQof9PILrAuuw3BT0Q0PYimWCKyAVftE5MVgFbPQyKz9XxU0hVjq
zFh00UtVgyDl3sdR16wo8W16aC2sXn5bHTybQvlAGV6TUwKVm6g/HA/UBVoRrJcGcFI+TuLdSMJQ
31qLBbK3IKA/qMX3fhR+dAuP/luVHnDYSS1Pp7pkShBl7nbtOpZXeVLsKG3QQEt8w6amwrcnoUKY
VCE4sfMgkMXdFDZFaDsDNuq1k9oEcR5GHr93ptwxG21BAixQQZlADkI5nFMt0esbn/HxvJZ44YSD
3IFEf2gXj8eKn0UJW677XO2zpQXfdH8FBFARZOaHVp+WAlxAR3iakXLiUMncelwTypYMGW/aYcD9
arrqQb8DBpDlk8UeitrTbhEwfGoLUA7HZ0PCLOyoC9ZS+lV9To8cGquVY4zbP27CvaYaayT+5tBl
Xfe56rTc+45EpoxzgkJNDM39ee3O4JTmN0hLNOIzD8Y13oeg4trIeZqnU53m3C0+RZqo2pDW9U/X
O+V8qqRcDk+yrCmLm/Rb9M2w8qGOadMW/gEBmHZWvLnYFOmJkVXcoTOmjwequmdp0IGwiNCKcpja
mz2QcN54HhkMgSC/RR8fl4KaNVWoc4ABi17D2s+yG07/3TkgS5aNvTc7a7rKnLWxKF77CNdVbf4q
P2t7Ago8FOGhvV+Ttm3hXEu1BqYFbV5ArtIv3m+bJHtiIYQzBLOAGAY/Q5bWRnrMqgqpcJAsp/oS
6qqW9hWXTB370RhneYkWYGaJg2wOh8Q1BwAw8IBPxfFfdfy8OwVh654vVCLWr3F0Ysvpqey/PS/A
ZX+LJbPDp3OGatYQLqsUwRwOzfOWBW2Qbc3E72vBW7Tt6JB4axZpBqOr3LaudQj0qQD1IyyMqhMG
1WbUERfRVycQOSOdhMDUWz8wSA/r2SW0x+V82JwIQjzEa0pYLeXPYypV+DW76CaOeB16znMhOpY/
E5asYFIN986i/4GvQnpFXwau/TCCoQO3u7YZiyILpuZ68X8S0yltNm2g/eY9McbMcBick/JfPcS2
+Uk7WK7HkfVgKyhF0fAQ63IO8c+1jn5cF2xQybgheto71jKiRl2sDzBdhc+aEBaI89ocFiSv6XgT
CFjDIYi6Qw6P2ighx9GsQ8BAMfcXLojC63kR8/zq23WKKj0xOVVCQFxUMmz8guAuhijgJJr/vkM2
NdS8eiFNbdxc4DVgf0TIhKEFvVCb0bFOxBl3P/kfUUPs8PjrLC31OoT1q5NykKwtcXFON4UtSlur
F3npOb4o8FZw8Lw7D8UpZtdOBzgEJ+Kim1rHgZdqasR7GwuEx9mYlTzjXHEyoj1orUHUrR2X1nXo
UmONhcvrH7eBmt+toKqth6oxqX02+dkDUQlNePms3b057KerkH6FIWTWHo8IBPgwQX48qYe1FVHk
y8BMmwmXdowW/yV8yFvLJEE+HF2XASMeqxYWDhEd+nz8yl3f50lVPwiaR2nTs+sFjG9Khk4NK6zk
YWdrxmn16I1I9ouPvDuPGDriqNgQcNEGsSEdlkvoaTGJwoCfKxn6aLzyfyFAyS4wjS9Ea1jWpU0l
DIsFOqFDlgNTQeFSbn6NxEGImAcYjH2txNaGusp0DaMYzyaM9Ff4hF/Vb0W7n26vnk1PgOkvYLRu
N+ZxZG8dxQoGABMGsuna8BR2ts2zWkAGAG+MOexCSSm7RhzYSzBW9uftdRQ5l47ImDh91EkfjNiC
MC1ST3KhwZCeTyJi+2NZopiqa/T88kRHwxHbrxD2vhG8jmTlSajxfjA8U8zcnJY410K+ngDjH96y
rXNkOGjsi7TlEMyluhX2uz1V/tBBS0gAIdlzXAWorqMvGgG8RH1wXEhIwFtE/ti9yqwig6Vvej2U
hdwZLa7cRLHEY24VDkHJwk8l2blhorILDV/l854v28tewo9tha6IqB3eNEQBr0U387iNj+/e+81r
ZjS8tabjl1v3B+UUUlfvTk8/mwbqG8Z+JAUeFugbKoGu5QYHFZMb5cSJSa0M2WlA0cLQZkpsvQXr
BpN37fuqBFE8V+nHaOogFNhRnSKMX6yQ19dTXkU/WAaSwNhlC0g38v4vfUScTQUrEBXmQ6JSRelX
Tj0DnGpdD9W3da7qzRllkM8qUp2VfWGyun5TspsPEbsinpx1+R2JFCODSX+J/Sv5gbb9ihvxOi44
z8HJQ1rEqgBuL+tSAoIUdMlL858Q/taqSfuDz5ngF5BVU7hBw4Ts96xgL7RnamRiGAfVrxuEuaDw
yIcUv6d1VdHlFmcPeLZA3KO1rwh+nPCMZx9MwaneQlAJ1IUVB7QGiDgzbIHiClknllGDpBypd/kI
cfud0QrIxL2+bmTBPsf2TBsWfrxr1UC3MHBqoT55LKrBf5ZrKAhk2Y/9xyIqGGkQNRvvbSYxtIPe
H0KHu7w935Io9x30KEGb5nGSOBzOKr9t4nFJAyf60I6LTd/lJfCjpXooUbeJGrKVgP5LwvGc/otA
OZO1APkz7vs/Lf1070skwc2XV1c2NdQVJ4jTenzgHKobAxNPxpF0fniJ9pAB3Popghv4oDr6xJ6c
2aKuQnu3Nnw2/ilhtKPn9GZXJg6oPnLv/JKD47Vu5hRhIOfly5aIqPpnytsqOuJzWc9F/8MoCFPC
pbnEs5AspQefeGc1yHAbHOTOWHubrZW++hONLNe1LiIdzt2f585b+3b4Zx7U3rzvQlZr6VkyVBE9
YVsN9e2NLJSQkPq5rmgZJsZ4xu+Pyc2b2uYukNzw37Do5P/9XjsvAFOF1g+nEuYb5FRi+kCV3kLL
axzUslVEEvyl2PkK4kp1ZC1KtIEmjqeQUxi5a1Or1Cc8417UdmX4ec0q7XehLldY+O5KVLw4e2hK
ED4YEdOs5ZB5zYcbb0qnykJkoWR8Xvj0G07VqYbxdcWmZp04cm5OQWC9dFfTfGKgIfWZkA7jCKjh
ywzYoXdmKkiejLOSwRG4CiSiLERykzwKrVwY6tzpNxbiqMkhZ9AD7CysOlRNnLND/m03YgAq8wBw
f6lcVDawLazauJr+LgcZSAW5vVDKoN1XxaPYcGMOc4Pp0l5dz60K0EYR0Kol2r4yFugvKVQM+UR3
xuRms5iDaqUTRicJmVNBa6kgjSirzZwvXA074X7M/tTzcFgOhE2nY2v85baBlcS7xa3LIfFqTPgP
FBqqdzHVonWAWhqWJlSMqaAZ65OfxjoocDnsP1R+ui/+cAomKRED5b04WMJUV4NbnbYShTMgg0vs
bDFSarYp4xAs30OgaGTNbjUHMbVNnRMbu0L491C41ucaS8AJcneoQZ9XQ+vXuc5nWpTOuF9Otyhd
332LoTPdrGplAFwARcVWHqpl7ODfh6qc9dB/ig0pxY3Mq5WuyEl+R/1dOHEQwPuFK8BFZRqK8TCD
/JNF9Q1I6sjXAX0YKtXlMaTXdb7GtNSzugXa7xdzNCdPZOEIAatAoqmqUnODTTOw8MEsDqcrPPqq
zOa+USRryufXFfcEgUM+5Hl3fDyeBBQkbjM68I51PD5XgIQyJ5G+MLbasROhMaaRgmsVLfWpvaeI
LzajhXvBZtGihCar0qwbA9OGAABGrAJdE1oJw+ZGk/T6LtTlll+YLaAEmoH7Qx+anvX1EpCM0HlN
0PzpgfrvwI8ETOhej0k0LUIfntsBZ7iTs9n81OsQhYZs2GxTptRdLePmDMAGjIhUp93SstwudUng
W41aBhE49sMRN0SjIq1TPqZK/rjuQlTTOVyaD8WGPyo+ADIRAR9oXqw90mqD5+WDuzwyWaYEcu3G
uhURpwqU2isCNy0nHqCfAbVEvaRgEsto2jNF8vu7c0cij1ngw1uQfPQFZmtFdnCsNH44IZCrwHmC
1+4Xjt+aquMd6fyevQzZTUbZP8UQAC1WDPV1Id0jNssOjhBjfCLmJXSdJzpSBJh+m8xQfplxFTBt
6NCdRLIVdR67ogEFMw0ExrqnvwlVPJapuG14ydDIx8Q6jNQNr4F2Kr9rnWbSpM3d0IiTLDiCHyAw
9P2VhUEghulWccEiVh87ejYMU5vmvJiMNVkYEi27aTvI8diJtf1MmBP7j1uabeq7TX2rQEQ5y2yw
eWDcWemKdm2d4mQby/yV1Aw7KCTmXpYTvvXhMD1nIm+DdKJUFoi46HCLhQLUQHLWFPButI2u87FK
CMUAJnhEDxy4VSTHK7pQp6mKk54S21HjXDPutCWuueGZZ7DA5d66BJGBg87NeJykxSxY+eR8cSdj
f9d4KuNs4XQ+X5SVk4T1CQpItPM0DQUYDZb0JK6Qbb0bogaf/kyVBKoq3Vl42EME3dx2ko5y0/jT
7E/T3s06mMUdkvdUJkRLz7/DcT5bVJsp9LVB5kqaFQJvkE+9ny82ahUFhIfylbxVE65lIjypkFPY
/nm5gWMXUATWK4FN7cD0i9FMdBj6VFi7M//5cJDc7hCUBMw07BuIYxWNFncfiPXu2OXY5MCXNmvO
9bZJw4ae+FmfGqtyZFJAyYcmhiAl+suTh/XdJPfzPylfquLKJxiBxf24VCunmmmG9Hb0Hg+nkHCM
cog2zOwoRTKvszqAXwhA2hqemv0gaOG4HB0eR3IiWbZi6k/EuvKVWQSgNIyDwb+M8fUxrESnypRB
xDwkQagM/hi+DH2jGOmg/fC3AWfeR4uvq8jiq127zs+QFWoyeNUci7hyNipIxIB0xZro0QBauOLj
gmIIUo3zTQCzEEZuWjD8+QICPYT8WJD2wgcWznE8VfZX2Kqta7ZMm6OoRlENXsIfSW9YGpYOh/sS
MizCJG9treYI8o/sD1v4WybTN4DHX82VW1kWHIf9gKK2modedQ5D5ET19doXfkR5nBNEB/KNBpHy
ZxP2lqGv07Fvsqk9Ek5g8BJLk82M2kTnsFBMI4LBo36aojepvZ7MZmKwtNBQTe2MURyiRaEUps31
QWr9iJPTnAlKfe4f/sXrlI/KCnVhqOExQfUXGYh6oJ3x2dA7zTRWmW6wgzHZm6buYSPenBzjqaKq
C51VF4/71wGbN3OSox7rwXkRB9ZLxsLFw7y7vftqluhpCW9JNrsk59oVkPS4NQGrMdNcczDXjRxP
Gv6vEvdAsFvFKmgRJqvqYYFkRMRXyQX5RlI+BY0un8YWw2rFGIPj2rT14oQTIptaq+A9kZVYFR8K
gQDjVNWTCIR/6flhDgeKwV3ExX6D5kqWygKtbJ+ep/Gd232AXyr6RELakwtvg1wQBchgkkH8Q9EC
zGgYMvcQWecCo2YwitwnrJCyjFlYab7WP4a2uDwBjpCAbpXsi7iFpNZf+qpfS5vZxcyfde06yKKR
Wk6KkQGm+HeDgKVEcv2bboi4ryv9BvfAOIBud4xitt51tTwW0QW+ioGpDVP/KMMXYgKuhZBfe626
VSCd6ca+2eYZ4QQPU6JtXt0B2Puyqd11CMyyPCaauEZplWKto1oRJMLeu9jZxaLpuOlgQM8l4TC3
PcJN0YqRDh8wlWLTmqxFyPiRvLvp8ShWSR+m6IsyWtaTu0ck/6mXgi0Re6xw/d0xLVw4VJcxyHbz
Fk9sIW/0HqJKWlPqiH7QtT5rfpJIaWfDpnPOgJPCjp9Sb5JA6SAgNVlgZvnyWACd0kkbdEmOOBi+
csAU0s9zcEPVzDdBD0J79N/qPNQzhQImMQ56t670WkukTHbOGeDdgoDt+LYmFnvAlbJMsInegxcN
KIQqWd5WcToAKlEiCkIWLoS6ZCvxiXEIJb8y/yeeE8Igfy8zc4zwqm3QjjmcjzKk88Yn7o0Gy/1+
D31aVtlHZcKRc/DtQJkOxmmKOCG5+haKytvbgPTtDgJXsi7zbshOXgwTJehIJuHa99g188Lc3udn
SSxoOypBHkk9hYbYvKA0RDVoRkE+NWL7FhNdZ56LkgbcOggZFeFVvA8Nq7n3i3gjwlbdLEzjcmNC
O8OzkCM+vkhdXkwhsO2e9nb+t9dAv/KcfxI4wc7V6HTDaO7BUEndIPZQ2StW+gkPTbZ5OFLiW6dP
SYnpGcpHcroxpItitGE2axKw7oVvikR1bQkz4T38RMk+8C6mHP7jDTysFUN9e8USyUw4XtfcyTD3
mNrd3Guw5KRybaCK8EQvq8vH6Rs8vuC5L9nfjCIjeQkVsV1vVqODR798SjY3NrSfz1Bz1Rgmr6/X
LQVQZ2NaSCEyRK8k+buaZlTkZv+q6oRF9Hq+GgpGBxYfSKTpHyhRVvj4R0sb+gJaLkPLJQZ+NkDN
fM+opsT6XYn0NOqzaen0VkSkFU5qh1JRC3/NNv3ZJHzOfPOh+abtqegJqz6dJx/xzzfm3uly1pLw
CHpd7ihpx3am9czX9bkCn8xKpt733MBqZWxsCMpaVnHlvT/1X9N3QR0vE7tZMm680kXZrslX36pa
X1JbhVyK2iMxg+XkE0vcEemZPZY5IdrtuikF4f4aKjAeTwTI4X3aHQTOcHOfSYkecbMzzAa7rcAS
sywOXwdxOMzFlpaSb7nqaTKqlUoH8jXmzc6Xsq0KreI0ZVVX9mFTYQCBjQ95Nn4yKR2aZyHSFzQg
bNIuQmmuTCWWghkz0X5R6UIi4Khm2MmiQo5WVqf6CcEpwMedK/1FIG+ETYkdv3ldUpXnEBB20P/f
HwZrTs3ZivfAAMFh5vc402pSkQ/y/AqtYKWe7VXXhptIFFyhEI3dnQLIe9H8eW1w2AQYvaMODvKQ
AzzWWCTE54mFz4xXiiAkqDR2ThNrZKuuSBNWNn8Zbmar9KF3jLldRHhv2cICXKim4GOTOF+MvAJ1
ul2aecDQwol60U/ZyedGrjqoS1ycMg71TeME801nLNQ4yiExFf6Pmpb5inYIhTg2/SAVFSkEsQdj
kk7h5mXwsokafKUoo2SAWKs/JgaDNu88IUvWWNUybNtVDCt0J9yR8TqlY5sLhWryEbi18E3RKXiR
VfEMfui0EZTPJ7xWQLZeE7kF7YAnRyehJmZIo0z6M1RlALQPu7e8S0+BmJjR8v5ruNriNTboJJeG
4j4ua3OxQwTF7sSlOE04aVXTVF/xCoYTo6EQb0CNcJGX/Dt5cjhArXt82lMi7NibBnu7muCVY5ui
wyDdcemUrQZ40vx2zx7afRFWUQsXa/p4RXcJgxYwtcg/qVFaj/mZAWipxLTw4of3m6QbX7OKNb82
17Kso5XBEnHDNN60sNJ4sE3ntkgQwLSWhfzqU9zAG9td+0p3UGeZ/zGWhcRBCS1A8rkEYBqxPESR
TdEw7cObsQBTEuriWPzQNm3k0cj4WBwEaHNyJmwWIkYCo4nUDb4kOLvFQOYxcAASIP4TELIczPD+
ZsUhX1S9+xeZTNLNb7vlTdfxDYgYeMukqVwDHnvbEcJu8vKiqT79O1VoD8TlMgEiwXsSzGCxmlPP
WCWnaI5NNfRCBkDcbMukgqaGNgTVO2KguAyH59hnZM5yfuaUotTAXMC2YRS6EQDqzY08HJChtntQ
tGj32etWLxBmiYP29RPpVL2DqFZERjrT/qeU0HnQpCl8FCUooGVVKQOADgntHhaXsUpeWNMyAe7Q
uCZiukk2oLdeauX6fgRbCws/t6L2Y6KXZvKE8Au3XAzIOSzsLwdJfAHmMZDaNZEmD/1mIYtcNzm2
i5cgfRYVSk3Nj2OnYJNAeDwgiYTl67t6BLv4hF4ftMwjyQiL+IyUoWvJXlY+5MOuTI9C8kcUyQt/
oSYyI5TbtopcZVf8zMH6rIw1GkRDg/PcvoMd+FhpjuINGadg/1U3vBfFbeFAttNayW5kj+U2ZDYm
Yt6YQXaRH79OOFa+gH522wM6VRTJ5KJwZR//H4fwJA0GBRjWFiWn38atJ1y1d5LwLZOlC2QWTRCf
l9r1EF7C6FLIX1HWySjZLae9sne05uz96i02A15gK0RwL+AuC7ro9HbjG7QHM6LgfpZ58BmYwXow
tU+hAu6+9t9Tj6p3adfJdPdcEV9gjLvd3pNX0w96ijf+jGJgkCy2so7wn0dIMPtH8h9UN/P3P86s
eHV1KXmwemvxd0MWhC4+kMobU6VoVTonL3WvC5QxGaOsHXq3whILL0Ki/mJVoO2Kas4HTRj48mLz
6MggqZh/6uiZHHmpwj4AmeU/Ev3OrUmzOVCgAAAH8y2/ywBsIIc4wi+HtndWTJ6ffP5igKZAWLZX
FrhU7Eq/B5lrhuqpMO8nYlHhezaDv5/JTha69GDU0xL4K5k79VWHUuovYE2KW0HSAJ1QuW3Jqtpg
JRqLy2FnT7U11eh2OHYvOdXv8m+MIa3KFD5CIEGVldrrr2iUhlub1JEc+a62kBvPoCJEManBnEsI
9/jOC1GLlZIhGGttYkNVxW1r3SAq/fql/3q6AuIkvU9lrbtTTMVmF/PtDjtMv2AsGvJ6lFC0VsdS
htxbNRbbHqLnPs6s7GmloeSvp/FtRVkX5paiYDsgLJ1vLhDqygaG+QqvNp6adwGlU6GKvvO9jmr4
md/WSbWhBdrkC9sI85dn85BZHMbeIZxUdM7lcEpyIhz8r6j3fIhthQOuKrHTlzpL4VyHnp7N5Sm1
AAC/nI7d3ylaLdL1plFSoprZeN1pI6NpWmHxsOO6BTjtX2xJAvlqiBzuV1mbfCB6GI356FkB2V1M
dmjWAI81xwTmsS4lksB6yLQ4LQhAaDvOYJn+fF1X5IJkYGZp5GS1lQn1xkMQWNTqf2Qu3I6Vy5qF
+Ku5L8IdEbMfnZ6hEAPYVusJcTE8hbpYqqxPy1CcoSVDQ4jFJhEwcEjLmzEA6yNxZpartx9Q2AfV
GiLUH1K52UxR+bduY65Mgu/XaH+sbio4gsPgq8ONgPoLKU0X6tuUGjOT7i+w5B2hQDsLZvtC7BDv
kgaiMfk4pWqDs9s1IASvg27d34O0blBsoFjDRDi3Q/LYwPn896of520qKZIGemWH9drkZ5yqa0sF
a/BhEKMu8odOvfxbxbMPkc+XZrkf3vXb7aXUWDyAhlhwsqQazcoGuLPTRjjbSy4d5LiX48fPtgeZ
CFMN/rARHhd3BsGM65Hk9Uwn5KYsFiwb2WmfOk6vq0q7BKHjlsSx19Xf7f5OPFmbh9nV8y3bDjZa
Fc7N1EYmJvHzTNrfYQrPv51eyz7hj7BSGZaoMqSOdwTbBG5y+PKBlmE5RAqOCddOmaDXtGK4TsOB
kYzfxl4t+ERRyt7kSlE8fnyCpHt4CSc4EM9Z5w7kcvn0/GAAiI0xeQwQrFosAA9Km6nsx/bPVoo3
n23WxydQJmUnXgHpOTxugZPT+e9kjYo9oGbOlpZE/2wjNAKb6d0LR/j1AuLkJQ4a5QBDyb1NOgZD
jXZO2txEPLu0dijTeR1m4aX5GJVhnb+jQk5HSvQk+/nXvH9XFgDIe8Gmwe+8+Q7u7Iuhc4Ujhk2w
lc7H/YMzdVSoXQnftger2lFZazEen4IheMmh3WW3n5ztB+wsAdInAWkXidpFLk3spboHH2qP4fGW
zdm1BDc3d4INRe3fpk78QTD1U4J5y3ZnGse1kTdNGuXfCtBEJXYiZykrx2tZ5L5kGBKm1K4lLG66
aAOMWjAGxGiP0YVGGvPHBJIPC/QtKJvab4A1XajKA/MG3jymbT/R8dBr/gyGNviut55FLM9pdcQz
slD3jQHIqTpfTeft65Sd5cQ/XE3p1kyT/qyYuZIcmuup+SqpRBONjtif/2C/MylkpJ5EmwMLeJcw
w0PRH2dRvEVUP+BrcWcy/aHLoQsAblHvwYRlGUgHNPabmbokahnrKhut38Fc7HHmyC0NCm8KP8n9
TUEba+y/1pmiNJw8LXFx6ZKE0bnkdYGWfx8yDsHFiSvr3iFcnS2BTGmVlIueuySisKcs6w50OS6w
Y0mqgfrReW/xmYDkl8nOETcQLBqZCUATyLxBozRsn2+MTi7fYwJHWNu8FnKZzSHCZs2E+WkyCa+t
z2GBaKlMfS1uJphY/Gw+1aZNDhe3t+xVv9krPLn9s/S1rQnKSsCC1sGnO/vJE0SXs4RQq5DWDBLL
WU19YGh8odx6FGclgAblUWkI9IYhDJXLx3n+aDhKHHX0N0fwJm8KXYk7fzoArdFraCmkV4V8RcR5
mnhoEa8U7Ea02wKuDsEA8hJG1rYld28TAF5Fldo7ztJwhdi1iQixNd3Oy2+NVyI+e6X00xSTWe/B
Xl8y+Et9qdavkyc92ZeAHm7hriy8/9BoLExwnKECrsiabPa0OtzDubexaLxAvAjy1k8q3Ur+mJP7
YHhPmoJAILABbw6PslHMh5XT6hBm4ZmcbTY6y9wqmnHpjlMJ8Zgqati6tY/OEB3mc77WwIGjoZtX
hBMnmoKdoO5dgM9vq8ApL1qzRPm5D+P7I/dLPhnPlm8xqaxZ515+DmkY576cMMjWdZkfQ4HLvs8v
yltJzAiDKgQdbL+dtRD4W1Fh57IqPUoE6nb3nQP62llsG2RwPU6odbaBbsl8T146y+cjt3XohqrA
CYjDoIEiQgfNYGE6OKDZYVGQ4ogvHFRBrBcqT68GmOH3ZzbV6Tz3DU1zSmwkTpV/ylHTmaYQpDBN
VNqSFLwE6SPdHda45Z0x+4tgT3DR4mxyc2AgrF8c0XRqszFvSXBYQsSefzUYiZEEWzaLB+3jmxyh
tcewmTFzQPxIff4KtjdDYVCzIsBlQ/ObPyJudfE4pv1b566ntMa8tVU2Xg3WzcUCjkqD1yDDz/eW
Q3XMC/ICw+qTbVJerWFePCtdP31fq8GjCnKp6+v5NIieKVuz5uVkRAMfBAdZg1P5EYVW1RNdFyQo
bo1LZuhGR1q3xW2QJMERS95yjl0Rz6D5nGPsFerJyetzvXaHqm8pDa6Z5RRdOnTKhPujIxKdq8Hw
x1dDGTVJTuVJGMp8e3xC5r8f3k0eTHpWPPW8Ch8KkFXcuE/ubA6M/jSKTB9KZH7GneSy492C3s9r
IQX79VrkrISTgbO+MRvlQdTsjUAUUbq8V2ftIRJ3J+D7dt0zcUulBQz07G6xSqWOdTCFTCjcWeCR
gYBocl3tfy1vN9KZf0rfAg4K3WgZ3cQlGENVWqx2X4FCQmTKeC+urdIY6qxIMn9RnXjMWo/RPo4M
pSM6K29wCoTV2i3vaywnhvvYGx7h8mpHhEpsNpfMIYMAF5+O/e1MdLSRISn3wFUnpPoRZ2DgOJ2J
xq/Ya1nnT4OM/y4VTXqIAutQ+r9p6HnpdXNTfzog2VbvsxUeq29rD8bFgEnM6yoxePYWYaVyDO2d
Z4Tk28rbK3ehreFnoLGvncjsFH9Xg7lqkXCB86myLj7tlcPt6ISjzgsUcnsq70AllNQnKFEdwqIz
rS/uTY4ET0laJAmnHFT8VsOVUkqLen1maexavrwiYBicxOp2dE9hE8C7GozaiE8GM5lBO8JNaTku
k2tZg/Tv1ONbJ40Z6OKh2xXi+ackI+0mVNvmVW8iwles58eBkgPQlQwowLhOelpaXrBNTxDWSpb7
NNVyqOikF/DYxyntJHaWN1nfq9MmoZv/BdSRLr7v4UCd5sD9E3M4P61dILGSiBAi55y0dj7Ihnou
eCtFV14EpB/xeaNlSQf32Hutr/Z2yRKfL8l8KKhbPlvEQhzF7jh+gbVACFsOL2kNcnSU/cgbeh5s
9N02UByUDgqV63TycL45Ndf71u03fbHadjik5NvaAUuydeWJwpsoaTodV0xbdtZBO+I24nCfp1QZ
t3as61GSYZ8RHDTjCKnltDvTMQlrlca6IRgR1VEAGVR0ZnxlKaxMihUR3u6vPHBmxrHwVFzuknvO
SzF3jhxNzY0UYEIdsBP0WiwoKUiV3RGxjFOK0yi6EIkEJ+K2hXd9e3kADFER+sj8fOHppDItzlR0
KRk4SeDjqCldNgWtNHEPJge2nR1ciEno4YBCx4fr0zYwlI0opSfrOTF4j+u97Los3Ee9r0fsWEqB
Ax1p+o6J8NzF9BEUwjgg5Aqii/w+/WofiH6UJadqzDj3kD34qXLpe9d9H3PPf8ymP6kecQdWFeDX
y5N7u/GUVk1tTXelcfQbsMDLqE8D2TPia+j4zgAngAVh5Mpu1n33CN4VS0G6TuQN1Y4j4YG99rqZ
vfJQ09qkU8EiJtusR0/mkP0WficUteXN9CGHkjT5SwW6bxNVxQqbMUdtnMcYJ+KIXheVctSORiqQ
Ig2+0aKCYzRHpS6MY6ucIAILR2D1k1/3a21fzQ3hxd/DXhPiHsTv59O3EQ+sBC7Kz+uytjpy4RXW
uOV0KNeRdigjc/t2VJ9qNZris1CMdsXxTju7ioQ8Puby8jZOCo8aYomHgJKb3QDuZqL0G1jIVDxd
UmKkmqBGdfxrw0xqlzYILS6KE6qUtwewC0THhfgjYfe+gIhC7zF2zn7XS4SYGJQjsD1wJKVwkC4n
yazgg/a3wUwJ/B6E9bveXjRTaJdUqp3eVVJlCwtSxzV75Mz3kVTwN+/umePG9mOvppbVIXuJnPrp
chapknCQ3lkvqqn8+xLgAHBuCIeWRrWCsASL2KdFAhUm84ZQFcvzQiKmWt/0D6S/BxGTZZ8ubgOO
tj871EsVww3GZRrErj7S+EvgxjNWE8C7KXU6lIE6FSLYAMQiqG+dX+FQ411j80ltEFx1paF5y8x4
cSAJxrpaHxnW4vlSiZRIJ5DCFZDVS5MAfA4+Ee6X3NvNbQDzL4A6bh5RTiK5/w5Xqq6loqan9vZJ
d2wxS5ety00DV1ENN79CwwATXMFKb4zlyATlO53AODHsgq//OKZVPQmyiux2w/5/ll3NfWdw0p/s
z6JveulR/0/OT9d4clOGHdWJkKuN4h8BIYG1INjPi8h+2bMgkyg4AR5UAF21mCCIufdWn8qEXrtP
RHV79BWtQ+AoA5MDR5wOBtgnXFBKHOr1a9TB9oa8JjwybdGQ1dwHXBKiEskzi6HBcPeMkfHfUzwx
tYTBUJXEh8rm2P09gRNPnPXOkz8PgSV9cDkMlmw7sNa/GVe/i2YMMi7Kri/tSjegfsDeBkS3e4OS
2lqJSUjcCpCWOgnhPpoCiWwBxEmELJZY5n6acY/Qwb/F0vrUBw47ix+91Srrt6HOYy556FyDi7lx
iKEZiwY68yfsuWbjtXSL3HAAHd+HFPVrD4N5luF4O1mp6QU2p6P8sOusMa4y5p5ZUZ+ytWRWNERS
1KnBazEmS5ZeHPhu3WzGu/jdC4nvPDRneDGr7UfHNe+Fc6ywbVAo0XBS3uQi/iRuYrmo0qRvHrYf
WqH56aSADWk/3tHict1GjErRZNyvLhWg1JP30S8n1Zpdw8jAh3DZKBYkSbZhdbnL2jNOnqXWn/Cv
W64WbdsfmI9HQC9LxsQEhhEbnB7PZcDW2tAw1kD2wHYQvMWK51f8BTI+Oxw0NT4k++oG5nZ2mEp2
XlzB8Z8oVorlHGlQZT7EOd4Yb+TTHveu338DCdoQ2n2ArmZIARwz0h23K9cd9K4sEC+eKYQQKFCu
17qyw1p9VwSX+snaOUAAYmL0mD2sbuuRfYP81i7ElYA85hZMnF0TiBxn8nWnDUJ9vZb7XXkURlWO
Y2qLSFRhZE5YgAckvfB4WDYWQcMC6oD+jpyKR3SneZ/aXxV3tIrDciZ+0enCSjf2Fz2ZkuG/Tyxv
vqPpI+Ws1E0njpjRjcRiPjN+YpN71p9DPdBz1P3/evKHRzmnh/4FA06OLoZNVkCy2ER9sBk7zP/W
udSw/tm0I0YRWoHvu7q9LnYHDiyQSIL9CL3e+F6MM6b+gzeTdFOVhpGS26E7fa7QS8zZ24cdMgDM
kH9iBcA2w6I3/LHPCDsOwOwrYy4k7kPBSzSYRAxVW29D1UlZE1FEH4DwO9im98CtderxL8l0LIuZ
6CRwvbt8nRbsJ7YzaNp5l9qig6CR3h0qfiOSYmKt6BwAElBBeTdU/nl0+an6QRF6KHxPhAQnUAyP
GiD3TySzK0q3T99LeOb9abEi++a7dSSSnvarR+H9m0PE2SpWd4dkrI1w1pBAXdKWSN8Wv8Sz+Frh
sjB5tsvMX3mdQWS41vvhzZ+ZLFJhAyIYUhQzPSFQz+kaVwzb3Mlhi6EgBW4Tzcfa1aNd/ffz7AMB
1vpjhVYgg0EAQzZl/dywTvaPzcPgeqlEw7u/wOg+H+ib3fGcTagfw8T4Scqq1HhcUimBb4nkU66U
+rSctg2lG9bIGtqnZlmskQcZsMkq1bUQbIUBeW/ERUBbQ+TL9/ijUDbwxKcoPj0af92if3VIB5q4
zNSd1vcbxFq4rq/Pbp8+e+Ar2VEvN8Pwf/gSlSleLeJ65nt0tZ2EHQ/4+DdEyUSfx2gSrO/lvrdD
t91eRBteLKaLbAZqN/Ga8Y7iWrEijCN9zvUw0YkOX6dAzlJLF1+Nq+RflRbq/Hnrp+LyUxkOMajO
yFaDhcvBDwoL3+XoR7vWmC+7DEDM0QXLJCdPAyvjCp8a1WLNKAbPkbCQaMZr8cIoykZRFdGVAHor
GUDC1z1axTyrNBRlUnYqhtH0auB3zYj4xSa3Wp5APSbtI92mhgrRz+kXo4Aib0uxZt/sfkuWmvZs
4SHtDpGPZFBa+lOXB/mZASSDNQxs6DKVl5h0k5WEP0W/tGa9PZinq4mm1LUJ7qJJLt3DlVky6vrd
bJ2WrbCWW1VczXXafBZLmlAwv5Q8wa27KGANoRf99c8SDW533Bha/YNiQwh4TkERYjiWZldNQ505
zcXJLdj/SliVqTD0r19lCJ2o9hQlBI8kWgiHXirHRgMgqOd/mEBSfc/pwKdMnYBFABqjnXGEIE9h
8eTww4cSBG03SAuhsdghrt/IJuZ923HOUkvQJfAjH1RAyQNkYj421MwnK8OdWc8uyMqs8B/cbXhH
nv/EhwlhXBc85Y2pf7ZwgGTNb0elsASd7XnZuLOpNnes0so1afuPT2i1jjjAW+u6kfPHwAunemKe
cFy+LVgsR0xWxAsR1kC0jBLXNdVRpMWMOofnu3jzJcLI/oE6JI9C77/dhORPxocb/anLn5rwEqut
VR3rd5qg4iF8nUeootw27VrPp3dPYq1IZhOwh6kHgw1ZxSqy5hLGZbLmT9c6MjBpS3BGdDmMNawm
0Af/MJapqC6CvWiYgxQm164bUjhnJGA4KWfBEXe0g8jcAGXrqeAtVkLZ67RJ8dt0rQnXV33bs6DQ
wtxuEJLF/iYj+2+w6jVIgVBGhFByE0ATdU4qualH+lQBPgMocEvd50Wo8urUbwx8hzFagznCl0ba
B31sXEJwbL7zeOcUtC7m8IRUAOX9nA+Jljcd9y2LGyX+hHOHT2/MUJq+FRXmy3OrY4DdfNZoISNn
IgxnCxBwsvIf+lDh+qgpvXwXot/AAIk++1VITMB5BD9wvpkrcDsRxhuQzZ2Id1dt2VIEF8XOvy/K
zuIkp6KuZ/Tofb9QpdM/G9QVtzW7Eq9ghg8pdnvvlHhnCzHpBG79X3YFQQSG+DBeYZbT+RJ1pjyN
I0n4e5K9/IxgqoorUM+yGxAqyNY5JKTcRPeTzQ/QFZ/TT48ws1WtPUrGKmbGSJmYlkuk1TpHhIJe
OJwo518FjoMCec8J7I2SbQVAUw7C2GEFMDmOvHAJ91jJx8Ju0QDclvp+Y1u5n+UCHXRWvJ9JDeKD
CwnMH7qKMxos8RDxi44mzu61ViaLGjfdI6nQCmT2mBZa6hnUbRCbLxP1Nupmg8sENHsRtTm0FD5H
r6sdjEI6imXOVEXJY0asB+FaorYGy54CJOCTA2PrZOL287EsNmWKFetfnkcLUNl5EhRX+Rod3ev7
tiFMZo1Y0JPlpzQxIoswFco7Ps8b/JdMZDQpl7UXkkqAbXvkB2EwgEkU0iyp/Fg3lcs++5FCznvL
0mZuVNvDmCmi2oO4Km6JqKD8KmTkUp4RsJa03bOilq/WDeD4sOe6nMEiBnMZ4Bn8nw4tEQx9Q6mm
VywPNF5slo4Lhi7YM/dSzetjtNyDyp6ltGap3cLbQxHzeM57fqPo4gn9IUCzkZsLp7dQv61tsRNM
PlukxClHFFMcpE63i/M/gWj+kHoJkQxa94UjZaXksGiBofMiLMMaBJgrXlB+bn1DVcJoNIxg2zQ5
kqeKJnJ9q5gtTFNrnaEw4R5gA0A2SrwVNydEXH1aKfJrDE35EfvMsW+c63R8HUv90zidh9ev+pEt
7GRJ9027VE4RYyIIohS11RI2WNXhuP1qIjAXgpnpAJNPEXrRff3e43nbOQSduYxYpoNHWm+DaUzM
HTa+yQjsRosOnx09WAkKFD6pYxxplQ1AEeohZaC0eVmA3TVs/wq2qq5Zl9r4dh0NKz5WA1GR2o4h
j4tFK3gu9csJTYtb08qvypEWXX1+D1aOiNfvxEOoi6vVQ56zdMOcvZsAjBhn7HZDyFraNkBc5EGP
80DTk/0nDrBj0C9qteZ3dc1IGj5Rwh0AtqxfLDUyo6LBPV0AEoNpWskm31Ljg1ZepE4ImK5yAL8d
x7aRxEGWiBgk90+RYqDkD+EADMS1Ci0Irp40IYN7y0VP2vWtnAvmsVT2sC4CNZJ3d2vAJ80O90zj
3XF9LRae4ZH0kVBz5s+CjkprTCBZZ8WUe9LmKD4snGs4eT3vJtvfAQJ2EsM9AdyEbcIULg9X1odz
t0GirY3sQ0qZiQmaJ3U3BH0yo5OnJNL/5GMjx2XfMwNwyaIDe5OOwp/bDXrXM4V1Nn7KGVZO9wBa
xD8VhESkZowzQr/OGP5gYPnjr8TjFSuQjBW/mnCKme7oz62b7y8BSFAaM/3gqM5mUlNinfFpg3SI
npItS/IxLmEtfIAEg//qfoAGZhJvbpgh5tnLdSuRNzjXoD9Bz83LjCWuZNKidTPOTPs1C4MSoGbh
2I1Sqtt9l9mliqQulfRy6qDvr1uJWwfaRWbGqRpSGTiYJE48SRgkqwtqC3wmjbnfFx6GwHfoVAO3
oth0OpAKj2EENviy9Jh7CpCCbGf1FI+65QYEs2fVpCb/a0/n3XE9mz2FjjLUKuCRV5sTSgd6OPm6
yKfXqZkBNZxY0gG/xug7ahxw19ojEyQwaNp8MLcHta+LsTPMYTCcw8hECe/rVMAlt25bNd+erSDS
e2uDpUYdPI3ScDuQA+UgjwvwNoFev+8t+KUk9ajTb1Ccxf6njbwCzY5qIkk6ScKTt7xW35IeKIyg
vcP1RwjpQQAcniiP+cHoS9cN1aFPUnalfHvAiTyJK5o2VIfNpm1jFhPUbrkdtwxDB4B2jFfm2cCk
gT+gYW+ZClrrHfjcHF/swDWn7Rn+HLxfftklOzVsx++8NakDPbEYlknCeR4FYSaDni7mOeVLnyui
ilUMdzxuN16AxhCkLVddkKP3TcUFevpdjPQu5S4aovy8W6ch3+jc272hBTCCA9DPhbSc2DPrQvzb
ofq2pV50l2hwedtfTeJdxQe3UuhhQBkH6RCyFpg8W5aYi2cL/fbmbvgya7ey+shfBZ08a/joiR0Z
vRAwTMmlRIKiCu7jJA0OYDSqlPwoU+COOwlZ0I1QGRgV5GVDduvcVUb0qwgB3Qxf2+KnULUK175+
ygCo7zifD/kDj3ArayCn5xcOHPUbfUuSlTZP08Bu8CO08GWF76VL9/8ocvYYAm629AWcDL0PKMtO
9ZmJHopSUt0EcJ2F5fD512O0fLOhCMyb98upbZNns84yVDcGOLq5+BHh/bydphC789/lhQJFuQK/
JoYXGNhEKf84Wun+27ex8fs8jpYG+BCDWSdITQWE/4Uq27Pl1zo6qwKmXrcaejKOEZcN8w9Qp5A2
6drM6AHkKXUPr0gC+H/e0w3f35teGteyuZCXmybZ2PB6+HdUV/cgp+Aa5CxLodLLOhOnkxNyFx9l
vVfaJZZhWOVdJ0i93pkbyvM1r/nFVZkMMlMOK13pYd+JQaPqimYSRteOjGbEwd6MIegKtT7QAY76
8lQesjmADylw8chPxhk0nYQYTH/PVKO2c8AE51gjAMzezIFwW8TacyxARDd0k+cyvegyNAeq5x0e
eZQuqPF4a48V4qW0FT7C5cBDv0o2t/zU4w3m5RvgpOVwOz2QlTqdLR2L+tajullUnQHof4/76zey
dNbxJivBwLM68t/2gJn9COhyfLlE94spTzidcelA/wdJ+/hCAhwwYG0zPmEzzrzRX7bhFiCaafjR
KssmN9pd1Hb7kn3Sn1DmCuGKRGIIccLvPSvn8L6TNDOTs9dTUylWGm5ggObsntDTPLR3oK+06zXS
PlmSOxP6sUkwdEyYxETA85Z0+cmAzUcGvlBevdHbG47awEeeT8dufKZjoANDUzrCMd1PXkKhbMSX
6I57UFuFbhIw5mcpuajJQu81KUHZ9q7f4C8fT1QfHrxDrxVwa6ZHn2eVSf7NsGVpxaMrZlpaUopo
pncXM940gz3NkWPDEFfEb2+I2jMcEc2f5OGhGiCWeCoy8u73HYGtetVWbQhvJKCFiY6gg1TxrPoq
Gs7NRyUb7d8Dzb5XhGTKPSFCFurqkr3qZb0QuV82Whrgo6lVwr17FpiIi0vqtQxMls0z8e9bqALO
Q/tiFZx3h8cCLebmWHhL6TlPtZHuSIpYkfzP5UVBIR1OgvqzRFiqaRi5SN8VvGu0E9hS3eOt1aCq
qSnwfX47ONtxWUuxF/EOs1qoK40zGGBwk9EHUc8ZP0qbNYEbth4SfNFP4jJZlc3FKyzK8rxQYktc
/xLkwKvitIwINHmH3A95k4ej7mj4l1iBb3uA1s3o5qBm2WPsPoJCC44lMB5vxLq3+BkFJu0JsHUn
kkpa+4q0thSqrlDPfyPcBDPUCzksUgNh5t+NsORt5chPWPrWwCI/nM1WEH9lpf3/bxhnKIRC1iWA
iQVDEvZGliZKJ6k/hmFtOWo0WeNLFRPjaZilGtnrV6rjzDO49tgcfqcugbx6z+rF4x8IksToM/s5
Lvg5/Uzb9sYiDiWu3BsKVYQmqgMpfegIFkS2K4jEsfkGqeAWmnD1gN3k8GgHJq9mZn+3V420k77W
zXTdTIpN05BgsFJ3qmdUOSfXN3M8zx9uMksF2/eC7C+IGeXvXvt33uukYNRYUy8R5hYZUl4mV+td
C8GnWlPwtzy8ZmNSMmtOKnorWdb775be0hXeLyQENoeMwQJxsT1l2II+6krepPhBlFk5FRtYGIv9
dNpQVbunmbjwMkcGPwWwxN3ujUxtI0GlR4jfQoMNigsYiy+f8EjKe3E2zzLiLm5U+S6SNwZSs824
KxX3akWZG4LVwaDQoBOxzC2rJTM5UTZechsGTOZSZuslpFyAlNZKpdE2qfqO8TrJhfCO6Ih2meWT
w+sQ6ARNXHlS4IcI43PRm31N/wDOfTCrRMjnhA6X/63qtXRj84qwJ7Yw0YnIrnCoi2vhgOpkA21p
yv6A79LXx/oFzACFKNSXMYMgdiZsejFjxcFgjokEBvRy+ye5DxJEQU27qL9qEK6k6y3JdHhQ4WMe
6PQfCI6CSqdx49ATzUKrbEYPh6EluAKUwInAhLDaVwKeBMJ17QjmKAmQSNpGcZAtHp5ZJmoMVlb1
z7z8qPsGfDMA6ZpTJ9mi9ccuSjpwR64kTDe/GFevaP4REYJlf96YqtkuBmsd9dvEOGY0uYNIEvEo
y95VKYEWStwINcgbmKR/nZg5KlfIafI5X+I2mNxYvFI3P9yIigSu9uwFReiPPbQGbZ8WIjEOBO+Q
moX5DSR1p4v9TkRXS6C609BkBJjBvTZJ0GCMlav0jPpVWYdM+sNQEGqxm9Ay4m/TzKG+xs09Yt0I
nuPIOlDP9YGXpC7MwxM3Uf6JXWQd4r5tHRk2lK7sxaGijTALl4qnPZbRLR2/R0asoRTsbWOTBNTC
NLVgiCzhIONpTrWdIi1MtZddiDn0wD4xN8MXVfNvZE5sxNyr0Igk7+8SGf+1l9KA78PYofHX+JMz
t03T2Zu/EZ4KDjawf+iD83PtUppBpZbQyGrTd3n3MRw2GcCnRxj7PDvzmTyBtQH00qtJaKt5M0Wk
NkyVJWBwhBPm8YguaexcQBKN+OPSA2Y3PdEXUxtOnIgCLh+Mzrj1UUGNgY8GFaadnFNpzYKMCAlI
DS8u7QD6Fil80gmASFmjtYItcpGlsmWDjz3tlitXCgIsyZ/OegQ2Zz+kngapXzHdlKhMiwT164pe
cjn/YGbQDmQ2c6X25GWD1D58B5aN8rm6hoGcvLTE+CrTvgQxkxhvCjNOZ5+Lu4Z+FEPJYMY+DlvY
dEys2nzkygkUpStco2kEr4SZCTdEMVeq2EG2zLsrIYjZKX8K/IXy0ADZaIri7bo3aWSNX9Zygdt6
NbDtb8NGCmoAZyyhGx5o2qPu0uAq1re8FGKl3hzQwCqavkltt3ozQrVXGwOkaBUArMcE4Opk7UHU
D9sK+JLE28rnY9ji6lm2TwyEVZ2ejlSbw2zg4CLgsEci8B1dU6qguw+k25L4/7MtJqQdFyZAmtlc
l1RviR0xEd49PmQSHbronochWhdXtDoaYP2P+nBb2l5nnuH8gElVw+bjyGC/LapDpv+pliXWNfXW
GiAFlZFGXo3ClZ5FZhmL+vs/A0ljaTl7n+4ncXasLLiWOcZ85TapIWVCwXYXC7SA17z7OTOOzT8X
6eHUB5v2TnPOGE6d65002fMN07rYGYQFTHmDo7RK/M/lhLn722663DUrCk3fHUl5KqSzphcF6vm9
XI0JNGvfTU5XSgtLXUSr3pqrIFPlcnJECnD0AuLSTJe0Sp+JG6ceXR7XmAw3oveVbZuj2TzcAF+Y
PvExDz0R7os219l5kyasnVzaC35tQEjwROFCyj5GIaDoVDHFyh4GM0M+GzFcnM4kraAnGJO5fhZ/
vRdSrwCUHPIfcpjTgx5xFi5R0N32mOvDi72uFE1SzKvZpNatIrH0l+sddsPysxeJKTXG2ByEo7cL
1TyMgy10T0g7D3OdfvJFtj7exVluzjAh0BoKlSkVDVln0VJqCXNG3xT+INSJ/xFJLbOs1qQlP8Em
DL753kdqTNm0zj6/WWz7XhEaSP+sELCcvKLM2YpRB0BbdEm2TAOpS+oinNC8dUViYDcrBaliVL/E
jsEiD1S/T7XutgZoTrPU3MY6yHq6TjXrGS3L2gidBBCvjZwv95RBkClHuEvkOV2Y7mrCCSzgMjCg
eHHlyiyUdAvxVrJ3AqjFeea3scY9GySbPKLHO7WjbcxfD78hDuIkmRnLJvOBqTjCiT+Lsy+a97Q3
r5CKHui8112eRU9yn6KHETiD/lml/9ZZn/muXEDWqfTiiW0G9+jDJZwWm+5lQ1VV79tLcFmPDRgq
rwgg9PRvEjf3fxI4BoZejxFuMEYM8vGXCaZiB7xsh+cfUg6GHtH6mNy1pOnRP97R6oyZFNT8ljFz
oN48KZGKcd/vKjYQ2WNgh/uOcHQr/0U2zt4W4LbzZfP+cLCvQakgZlvfvKc1mdfDgDEVz4E7n/BW
MyvTTtWIt1DrIvJkWwpff3D52uA6Zo5wJnw87HVb0Dp3HxQCGUxuDgeMOFJkbxhIRS50tW/u3hGh
NBaaXVfwbAEqNmCDGkH707F259VfbcKjauPZFqGQKEygJB6k31Vs6JAxkNPWY6/aZAY9T9DaNzX/
XLQR6C6JIXjCSDQsRVH2x1FpVBWf3RyTXrTTkmW6Zs4afxHVaCToV6yx7xXeEJoHc1MdOjle6RbT
DPMr9Cqr/QLemU+ijMG8Vu4IdPNCxefyF7pi+FmottNJ3bykO5mP2GVW+RYkXiGh/4LmvP89Fvo3
I4jkmKrCyHmKoI68rV92VGpD1t3F5n1ehmWgIPcOE5CfJBNG9O6CVF/X5YOjPcoCk1+Bsu7ll0mm
Xqb1/av7faxCXdBnSGGZohVkqiQQRKgzkae8FP3JR2D+MB6zBw1BmAXfgb25Qae0WMwKopyXoV44
F2NB6FKw2lzm8lnttB+Ml71OIdlhn7SYo6wuiJnMgXFGG/MxIEKe87C9CB09jv2B6JiGr6r4CiqJ
Mih1JhlRHyLqAYnxs7gkAjVBK6k5QM+Aok4b8WmoqMgR/zmXmJvfutIRNjjPK75NBETzGeimSP1p
VJQvk28yXc604TZqACaJqi6kpiopUvT3ZO5z3ebAvuVjMdftBlFTC+M3oIwzh+lE6enS97ytE72q
Y+jJbiXOyjzYGP3kUB6OD6/7ewsStD5v0XAml4RSkihGxAwZvXP6ONsGRxOUuoirM/sHqOBBz/hQ
X+J6cFBpbvZ3lfeNZ2exzceIKn3lepWCnBPHa+IkaInZGcsnWXo68Ij9hPhkmXSFNXDQHIjc5nC7
df4TyIcuXo+gX9d8qIkLlKY4OTY/rdQo80PPH898zAnJYRzd3hZgV0vGvGgRbURkjCfBLJVXZH/E
oGiRlPnO7dZJD0zWAqM43xGxG9W8UgQbZZZSxEcnB1ie7dr2BmLvcHVbAPy+ClnSbSmLyOSyf41M
LtTEsr6pDlRaymUuBfDDKln2vhpljshp5dLIrJk2voSf/SQ0v59cOOiGcO+9yPmgbqoShlnykcty
fkycPU8SmO0eYfHjhvRL6iXKClaIHBghaLPnwo2H4z7DdXYBsZ7mq0i3Egy6PlBEluhXcu4BB0sJ
d+mmnKTDP2HRhzVQsphQl06mxDEnr31IljCA0t4V6UzILd+serh2lFyyHYuu0ncINhmTiWWtIOSS
6KOGEBpjHJMi2JhiEUPRUOk3dj9kLbw2OVfN6oy+BQ6BR8PWw8PDAI6KLiBdEe48TS5sXODIqV0W
LNaaMlvyaJdBnLar4BiWA6xdsmPzUWBHsyzV+dnp2UkMdNH6yUh29HXjfZNnMC4Bl28M+MdBK5CE
6o23AOzA4zSnbybnEOyxM2ZZWaAYUkexD0uDGexn4dHhvvqva55ad51GxxfaDf2FGRv0v9kzhOo9
L/bwP6D8Epwg2Fz4CzW6UToshAb5o7TSpSuO1dX2x0nRy425+MLCr1CgHxYrPzg50g5O/6F2pCvC
kjm4G4Cr8zSlrqoaTV7ubvlgPuJjHOk3moGMrEUGUMobCLo/eB4mtIbpahO4ySwyRY0WRd6mVGMI
lCP/gtTZPt3J4SpQ5oXafO+0SWSWgLLMOMEWt+S8rOvc26wje381qacYS3dAGSZjxcJAagfUhLz0
qR2xZONZpJxeFvUnLboYJ8eCSeTNr6u11aotcspKAAv/ogSfj+ckUDeZQ72pCgGKh7slHwGjaxUr
CH08LZV3bpkZSIvmECkyNfFPvgD9Oe2JFTQ/FOzO8aKp9OEy7PfU5lITg11Y6+5igbe+ZLCGVg7Z
/lgyvQe9q21H1mlEGi92MUrgT29NF4ItO/WODIxvot+QAWnApGH1LLS3gMobg55kGLVLFf1K7YJE
B5Io4OIlGQrqBiHQp80e899t5CF7R2hEP0pnTE8t9YW9JnHGO5LizO6va9oAmgDr6WO+sopHNS45
hb7kg3kNvDMtXMtFQ538jkHoAdoaSBIv1gllQoLZ8cKj1Qq1vAkHlD/Gm3i2ds8/+61sso5xcFr6
jjc6SmLNn/sOZaBUUAg1+3YFyTXO8Zj+LWya2YJSzFtFdI1vsUc5LborXUp8cwrYbzHO/BsiOc9P
y3ut2suP+yRQH7zhZ1i+fq2xmoLfQKqDc66VBZiw1TldeZg37en2NxONE8g3RSGOcPZtjpvPCiQr
px7vo0WbfdwY4gsk4Fq50DLtk8lmz2sgu6qvZLDvOQbElb2ZheByxIkubrH401036Zlj1Dg0czWP
BjLt+qwYNh2nPqVfJ0pD6tCdrBeKoUxeJzjePsUum1Y1NSCVyw1FYFdu9J+4yJdvpgtuFSMajUio
cP43ZVKOsAXDBQ3K8nDNpAv9VhW/rceksCKKBpvnNdeRI8MvMYaFKs2KaqRwN5xzhPw7IjF+CiBK
YwfQgSYdxtCHFA3uAruspNyd71j+dAzYAWxbJ2HSbdQclMv6n4PkRuHxgqghYvJSgBZU09X8SN6p
CYeAAQWiDbQ55u+YTOTrS781AXq0/RwU9lIrfBzm5lAH1jJUFFdaznAlwoTAyWP/JEV4ttn3enyO
Ma9b5EqDgMRW7G88Ar0GBvKmpVt+27YiYDFfhxqvs/lEvHbb1Xw0DOn8rjVzuMZGTX/Iu82YvFYj
2Nm5DgpN0VzlNsKwRi5CWiANKlpHoZ4HWrj/QeoO7gmc/j1h30ELtftqsQW+nv5s4Q11tDMv3UGv
0LTPqX4hwk1Z7KVCHPWnlEj78mY41MqU2F30cLBduq0bV6HAnKqbFzOEPK4HrIQhyTfFYW1wk+B1
PMd+4MBSuF6QlWQftdyvvYPg3roXQfi56zVEJBo0P9Tvtk0cCz1MRrOzSOfuyZHYDgb/ma56GDqr
cyXlYPol+YSW5szxMCNJQ14BdEVkeCRc9iJZP0nLwKM5u1f2BC1TTHTaiO/uIb4eeoycOyUQ5oAd
bzh3RbVHOcNT9IFaqHuDFOJ2clI2uIGHuIZNkfp0cp00ria8TxUDWJXemrR1AZn3YYiMKWa1qkAJ
g7JftyxWnBpML5DdW3ySJd6GRr9svqYLp57cVuDMs3YzVs+S3u4iGRyBwfunfsYfw5s+afqHa+zu
6OrDUVfD3DvONe+vqQsGyCQkPPCvutIDDHBJU/FvCQ+5EhRIS4zHWkKvPW3HR/14l84mbt+ibgh+
58zU6Z0g8Adp//IakfqpUKD3mtwcqXI5F4Ern21zG71lo8X1JCB6BKU7FyXX20mdXuD+KHpWEbfI
9A00d8LwJvYBrNABfp+Y5nTqBUKN5CbyXZT4jbVklslc3XCqVrUrBYoPwqU61g7Q0DkCmw+cWdwH
86+A6gKQsUQtHcfAnHv8IzPTUZ0WlT0nkKx956hFZl1TD/1AyXpgLSwzXyPnkfCzxFvLPzsWynKo
JbDDswY7P8L+6fI90jEXLLHfRf5Xh9J3JrCE7rf3r7M6QAj0g/cJoFZ2BlPPqiPBwqACpyHJWnJp
UfMwexp9H8cU6a/ha+M7Bwsdho8oKC6g6CK8kSi0w2HzdehqxlzoYPWLLSnEHS5ZyxVCd0Zjz57P
+Eum/8rAdHUOGFzQvF76Pj/EG73opFbBgOFvRWB5exon4IpNrTPGgscj4sL3+vO8FbwxICVHjbrL
y+CcZ5YyXJ9m7eBJzaxTo2gREyvydzoLAwUBobPwXLAc379jUjXZ7qM1YaqK7h3oepX0QLurDCcm
YVTNybIu+myE6jTLphQ1uZNJy3jq6Z3l8e8cj4QAC//985RTiGrM8ihdgWIJ+bJNhNh+Ufd9lviZ
Mwx7k/3WXeQ21yshFQ+gIRRe5IMYQO9mOEYgKdCEuw9nQB+RgQggE1M8ZrBduV7CbYwz/Rvj4/Du
QM5fv5kxjYADVvBHw7E3ipZJP7G4ioogcQH6mixDWUpGEDmG5GeXDtLBsw9WyePU+NUuyj4RIMTU
4mdk5lj2a8/Q5qt2fsUv4ZMJ5hgfBmApijcLh38Un4C26ZwkImbdyp/cyhsGkapjUP7HtGLzRDo6
cAH9DNSgn3bXSnoo/imhCBxXpSMEzaHrae9WuiFISNguAS7lumjKFn/cdy0Iv+MJlCAO13rdMNcA
0GNgBvduiTFKjYTmu0yXidqY9cepkbpiOq2t0EKNPjNi07uvRaS3gZD7fYZRSB1ftbOowLkB464u
Ks5nQpJzfouZKm+YFKZaUP0inzi6Z2Dp+L0JTrDoVaidCNLUJ9RlMjuQVGOpPEwM2SO2e2mPe9hj
RiSZbEPWqW5f8YP5WWMHQR6yYPjeCjYDi8YM/wf7+9Wd9smhHPyDIZXyAO9tQwD9ix0DtQrD9d4h
QEb9QBUF5rJwOUM8A5mfPGhcdvXoGGedfFgRSIEHIWrjf4RJn6IQEU7T6fp17HOqUxXNzB9kKIya
9myc70bB8DFaPeEoOoZsIfCbHSaooTBQs1yJ59Mq4rRJkaKzDzuABFgXfVoZ69NI8uwBZd2wR8xZ
fC+uRZkLeZuT1XIyp9I6SI/QJNEi0RKciT1TkbcqCl5u3n43E8bpPMjZ6HI+Uu+RyYbqCuEz6pkm
idk3tDTt1W7WFBv8BBdlfL+8BOUmzqlMFvrJpGlhGNiBwFPADXqJ9OdWYNxtfDNHvRm0YZVbp0R6
Rj73Yqc10LI2qOm10lBsZBTv+qLIY8FcdY2eQuSRFXwgyGiimR0v9SBIBqiiVF0JZ9K8JpYxcPB4
RFrIGmA+y2Dhl2/TZILTMqrkZYDPIhrTZaoEfxvx2dbcYAb1xlsp8YxAZQWqpBirRIy1QlhsOrol
x/v6/RXYjsCtt/vs3OSn7Wj+DWTwZTn5Uk+7jZnYdBr2bK2jIDv+PN5+ZpY6qofBjzfmrihMYF/Q
e7Sw55U2NQofO1treiVN144Tpc78j4c4C5MZiSiTIlQwGwe8YrbVj4sUgs/F0BckxVHRtxLspmHF
4vWPaLSikoLbwzVSdHw0f7dajZDhp65tC3uKGQZyNsbGOOzXPicLLq0nwWtU7jOy6f2UM6OA0O/N
xkxtuFNdjUnmU9t30b5huKLXPP/4KHourYTBGYNyDwJ3HVRFUdWUClxdHy/kYT6PF2qr+nQOgapd
N63WkVYvkOjx9agxoMUC7bBl5wo7w14ENNXdxxmm7KU0hDwTYpG/SJusrLOWewBJ0uTgq87R4Bhk
aMl7J/Tn1aUY4KYRJjQwc8k8K9X4PrceZTKVdz0NgexLy+C7uzh0XTO2vuKh1+Ubgckr2yZ8ZzeR
r2urA6gAxQzjTp95N8acR9kKkoLMiYemVdDe4AtmLJSX4Ccp6bNIY4cBeOUDtOnjs/8URp4z0VNh
D+BQc2WHvjIfYs6cOuVkAq18FDIMi0khHia/d5d1KVPIrvCd+B0rbPqPdymiL5pg2z0IMlhmkp5a
Y4McFx7s7x5PD47RSa6iQvkXGVjd/W5YTy51ZSbj6wh5kl5rv7Nkgr8YUBngCefstT3SMiqdFHn5
25b665jDiS8tS+Bg6dIsxubOL3v1oT5Oqoku51R4ppKNPCDuV1r5TdR50kxPWDoFpmVtd/NxtMhM
Kvr6JLXggRK6eCFBQrApYqTYPIxP1U/htWR4hGCjoa6Viy79ZjLHdYxYntKm2l3HdwX2I7dUoErm
j+gbZAQog0wQ4MQ18g8FZ22YY1fvcXD/3DInZ5xxStf+NZfg+PoJuZzQXomjuaxzh6AL8pOGjTjf
LzkRRGlJMBWxdVaT8KBqpx9GKno6dEQxOWsDOAd/MfMS1gr/N4kdpcO9nXNopawuZcvZll4Xn/P/
5O66YkWRCxTNbn3zhLmKohJyqiUQ6C/C5LdLkL39pXGISP0ks0/bzGuKt9hVe4d8hbNltWTEF7Yr
+nMY6ULqpKcHUh4ec5XT4qdyi0KpaIa0mphatAimOi6n03WON9Fxl7cki2P+/JNui0lqRYv9R5nJ
ccz1AHODmNSPXMjBLBk665qZzn67H1a7LUTYAbrY0EMn6a0eOcfqJR3cl2wvBizb+3XULPic2RaR
CIm3fmWht06ZJlAg2MkSQWK6ZPSSBvvYjKj0CzKUotzrCo857bLRBRZnXiKxe+6mtHEMzeu9pgKx
I8/zAMx1I79nNKLQmbEl+n3YAc7Kw7166xew9ozH0fVujqMcY2oAhBv9qskb0ogJs2XiWUkYy9FO
oaNtbCEIUl+HbbM6fzwUd/y452/GUBIUJJhrZoEpbGDUn0/56kHagQ5yoqGyEs6Zww/LhVoS/SIk
VXxteKK471/u6s0YDMl4rLv6qUzUc9fHqgjWFEmTuWUIPdidujN73zSj3KcF5Hq6Hy9EgMfXFzUy
cbPWSedEQ8aat4Z0+zyXAbnFbDw4iWTxIxHwldLy0md7q92xUnoYcNw3crpYTTCgpEz7au3/mZqu
9P2Op/gW35tG5vUx9Iy0R0uU+nYhBtnLlYpqEVlmN/FxKSNu3oSRwcynbJLivqltfWNo4ikRgjgL
bSrWDxc8xBZz8elTOp4Wthf7C2oS/M1RvkmONFEbsuSxmdS/MMtlByKTw7Z+R+2aTnEot14qXFUs
ihdq9eiulZPnezu36KrKkbV7phzEVDHQh2zjCdYSyLr3j9YAOfKLg/LtM41Wd5Q2ipN2/uLuyfr6
J/kZu/0qYIUcQag3oemu7qxo06vhnCX8gFOoIzbQoKAc+PduWfKR52MyDHyYvJg8XufezRwp2Hzk
jyBaJcTQ/bnSCQzegKAv4mCFLQtRJSPD4W1j6R3Ce7mSjWFiG6rYfkjQ7FCTW6ZkDU8HuhMItq0j
bonjlnJs9P3miGKAezy8TpH75eWvAsN9QiApn+WeMYLOA41eoQjKyqbq5zhCTKGcmwHj39ksNYP4
wDK6Sf+rfTzdCjtpzEklJbLK/CmsXwMZ+q7Rm5Ek7KLyEgugTqtrBgGa6CIzAl3JdNTGKxvDYbWN
vF7upl2lFaxDro+6Qq5rqAclIKPcikITsMuS8IYwdoBnhWXV5Qbkic3H2ulzzR8MVBBBHNROCrJ2
3eRubyh8/VeM0cTl9z61MBLXIJ8kjH/k7H16/KmjfutQrEbPgHM9hj3j75eWLuCoF2Cq+WAQD7JX
2VKkzX1knsAUqFhWlR6Y4RK8I0N8METPnAoNqKVqeX69PNz2HVzALWpE941T/AxBSXHw7fbsVpmF
Or+dxyj8EIqvUpxkLOGlwQSaq63I/cLVXCckLYcjPDx25M2Wvb58vmJBa71hho+jfkLC7sN/tGHM
MHe4kRjICnEWfZaZkap4ddGWYxtHNnyhhHR7IBg3ExPCG6wY3KoeGT+lawXKXtarwTnTTksoBmtV
KhwPUHTVl2AdIefwtdAF2S/bCx4ztqe3c1aXn/tYvdXJtJyNDMLTxc7FcjzH4bDoi37QyyPYvSyq
/EE2B3z6ONj/dQKd4cI1YqN9XAS7AhNG/T7ZDHOSy7kcWtqDkR8hBr+yhE2E5LefiKNDUcFGl1eV
WAL3c7dxdrZxoqY3j1notYIHUkEz1UTK5/ReIx53ygbAt0+H3naT7sURGirxNX4xx4KBW28cMJ/F
2iY5OVb8gbRVSPX5XZP6tsikNh22DpmWqrkN48vwQHQ9XJaZbEfYUt9f6VNzxEtbxDjWMzS5LpgX
MQorH5FHrcx7R2NoICEZekBT6f79KczXN+iBiLdcVx87WoHRzGgYt7x1f0Ne5GGgZmstddiajE3G
GtvrM5hohQq3hmavPVbjTIu6+5uD59kZOfZ2JMmhw0d3I8zIgG8+79pyAYoc63kMVmChXfSl7shh
6WALa7mGnXJrWXBZnole9ZghqYvGuzXSyyMq+pjnYRd6Sye79BaUGhn/r1I0e1KrSgKXJcdGUzW5
t/KJlUU7Ns9GZ00P3Aj3dPkiYOLQbr8BqIbPg9EMS/loPB48TGjrE8kkFo6KUSAIjBlheykfgrvS
piw2yCbolvkxN0qB+nEa6+TlPRU73YGzYtJOjSeDb59a8U4GCK6JenrnLsBiXSt9ns3D6Pq/A+ui
1pQmAWFfJPFwLkYijj+7cj7Oilll6hNLVWpgRI0vcvEkcG4hSe0TLY7PRnAeBi3+wjIWsEz/ccFd
8fAWsO4k8BbgXQthxvj9yDzA5zyO0S0QAFTaEETXMYs91gSUiF30zTPsxW5U23dKf5MM4pSTKzbW
D14dRbhor/AenESv1tTK6d3YVtXFv61WHEspT+waHNxPEuaJh/fge1NN/Vftg7JvxWr2sW1xPuJa
93P1ndRjqdZaMxFCL7znrO5fwl/pe8EhVO0Z3UKoEq4rLsX/8rUlKVJYDhczIFDSAc7OlUDgNuQs
OlhPrAtQiSBR62bGyl1flKaS6WVpLj4O31R8weHg9qTUYrh+dZ9bgOiQ5PNZHZzKJYBtylwmRXP4
a6TnCJdRefh7WEEgQ8tDz2LWOyTN4uJMMxnQ2By6ggu/EzI8qdZgWSasOlfNb/O9oRuxvjm3yz9z
UaPBQqoMwkDQ1jQeznrP7T+nY+xlyFDhvvCopMBk80czztc5P/+c8rQaB0l2hT56rEX9FD5QrB4v
CYOb7KHivVT95TVZiV4+kLNAHBhtdbmIufEZKF693JhlDQgZpdiPZ62VqUfW8mbgRI84vHeuVV/R
IMIYePzJiHaYOb6xjrRHCaJD3Ex4vUYricTeTD6p5nfznwVNTkfw7HW9XswQBrmlhOGZ/d2u8To9
XT3ogGMumu+mRcHxSaee+5Cmos0FHC96ROfWn4J1N/O4L+BlDREJJooXxre9FpS/DCRxzBGDZgsb
CJyw26gb9mN0UqCjy5oUq6FZBh0oM2aiwghfgWXC4gIBXusWRGstvItteU80nhLYVoXrKQVWhrVS
H2dewXoBpmsbLHusNUyX0yNhEN//Ee2rOXInJhwYpmiIhcFt/zYWFrgcTbBrZ9116itBPlDYgwlo
/Kzc+RlaGdhUEalE68DGz8Abkgz5syM+yPqTCUfosgqmZ8wyrZ/MaQUhGlxYzu238TaNL2KKcSde
y7uY89eEC9p2kL40GlJyXP69fuBsLaw2OGS/8/JWrAiQN+DGMptvTZ6JEV06s+JMmPJSoynKkrid
z3gl4uel80Nmt8WfrpsAJp2HGIrpgZv/PSerai/xEIhvazuBt3qZdONAfS3p77noazlb9YzgZFAK
Fq6LUz1FFuGah46FbMHRpncSrtpDzKPMTVtZSOCEglAi2acRayt06f5Sw/LUJ9ZyJfpcQC+d+W6T
P6qLHtmD/5swbaL5XlhQWItEpryYQeY7OJxfcNqirm++ug1/DRzPPoWZUpn7cUmHMJ9uPas9uzDP
duMzpdb12qh05k+JgPiHtjGo0/BFu7IK8fUbq+UFPd2MEG63DG8zYrBQ1fzkAYpboOYxU2eyk7Y1
oyTYhsDJasz1aT3ByU/UMOHCAlRj/SNr5Kml2wZx0zA5orZSA2TgNxe+5sxSObSrTwnGI9hGl6dk
NpSdqijg/2hn1dQDNh9OKUp80z6AK57lEq4L3iAgVVjYNlEdA3xmhJbE+IbB8ae6QhAEwc93kCLE
d44TtkmH+2uikxacfSWmKOAS1vIn1hzyH7c8kwWTJwKkHvyUG8imcsz0w6cP0yzeHBkSCg+3dmiE
X3YaF3z0F0Rd1gYnLLVAZoTe66Xn8hhXmamv99EC2Hz43sa6DMSD6qFELb2zVydRl/0lHfxfhtBC
mphNHofoLal+GSJgJaCvY4EI5ka1+W3Y4yEl2nXDe24n5bs6i7/QZQJ6SnRKY68KNEBG/uLT5r9i
SJxIGmtrw40BHDDQFbd5lLO7lHCVSsrC7yvLm6ZUHEYct5Jt95VILVrddrrOE7Ntvx9kEmrqwwK0
4nWgOhc5tvcStsnBF9wbrnmdZAaRU5vJv2mT/KyZjiA5OVtGyFgjOxBdyjTDkfhb1IUWlwZWbpF9
XRmN1+7H8S2w4kBW/5DERaqYkdFNRQ6iNS5E7eQUErHs9E7e55qNjB8H+Xz1svdDxMrz1ZbW//jE
fBoZACPdulHd+3ExA3CXqoM5s2TjyWDsPbTU+O4kfpA8XEQb37xHVExt1GeaoalQJ1Kq4xLCbzha
tjUFcsUnH4LHtI4sDShC7yhHwc3aVEk6FFcS47K9K67ZC6YKP1YdOhb+b/vjW+UE7KwgdCLp7Eao
ITQIkG9NwWZCsuaPqpYaH5CxQkusX++HY3ubHYl3YdREvKyKi/MEz0+hlw0oXBdUEuen2a1LE688
UZiLBs8VGergK8D2RybaRcqVrkrSuQXTJ44vVe7kTrDDUNggSzhJME1m1WDx1amozsp/b2Ukb5cL
oDubm1UVnmZfo1XUKDHZGpJ/h96GQ65872k3Bj+j6d64GHAhYzIqAQtfM0FHJ4CYcIhgzquTcJkd
0HoJsQ2EvFRMgE7jplZM6qsze/CSsHQNDUIE/yoYeqmAfBeNxp5X3DRUAy6cTQDbii2prOGw/pxg
X6McvYzcKqbjQiSgph+cP88RSE1NuBeWh8gVWKZZIGO1EALtPAtnEyvycHTd/t3vs5X+tghi6Cje
3+Lvv8eKeFLjzj5CwSlPqzTToWRnMQ+hMrGPMI78d77hjor8tTysuPhRXin0vjv5vwevjUxplXHq
yzQcAWu6eHQmg9ah494QDGGT95NdUHYvVd8b4DTxi1/wfQ5dLLnsrrNGlQEUrCif6TeziEWgynXO
mSvIOfO2YGi2g1UKyJRUL8VkavK0oNreuU9oi/BmfgdPptfOVmvriSkrTd4obozlJ0Vvp/1rW4hl
D0Gw6Q0vjf/2bCQyVdgpMofbLhOkvDiadA9bvtXqaYg6/FFnzAA0ouxQB76aTofz4x+iXjuyTdjm
VcLlpVJ9f/XKx1NMmExVBt645WQ8H2Vt9d0Y/u20eGRK+xo+UTqo47ruR73egtk6Udn3crjipwSA
x4/V3x821XWXXX+R1hCi18C05w/IyeGJHX0K88mpeAaKTML59nHzH5JeyyizgtrCrnSfWOmUwfTC
uNkP5UaFxzVCfNW8bZT+ReaJgx6jpFLi8Xlq7Z63KPbcTIgAtuJlDwiLXNBtfzh+XLJM1wChs7El
8opWkuHqUyWNE0SEVCF5s1UQNaa6iK86hR62XlWhucn3ebgWic8wKNXVxzdJrNZ5iinYeUx4qlOD
XS/2nTfdxbtNRkIVkoeB4SaI+ne0P9TFlQYapFoT6nYD17m2YZYW4kaaGpoNc0zaJTjuLv8nhBYT
V8VkBUxg8QIWqWXFvvAE4lvgepsgEZ3u422v1mSE7Y3ICbZ4QO3NDJYsXzptg/qSQvDWk3NcAyvk
dHkNRsHXbia8WJkSLuxLYNm+kNhxxjuIBifK1HJOex4gkYHNU4SxY670eX4fPVU8Y1S4Mf3Uqkda
6vOTsXt9og9fLA2TXiMlpk1yBxw3EHZ2frlj3naGLouxpgen3lQl+5IZ8QNF3cWB4QFdKKF2/Hh6
Y+9rezuK6xrO+nImGyUHCXMQjdiuQLwGvaaIwHEAyls3AFhwva9cLjYDFAEd5kqOsQqfqZPvI9DG
9wkiHHUz+motbNinLsTDbXAZnA8rAOa3XmYPTDwQBp0YUTk1Gvp1UBqqHw4hk6x9gXEcbnW1Q8KP
/YXs7mjx3cr9u014vNZ6fa8chZOrL3/q4etP5PWr5LSwhegZZwhegDyXNJrWbfXM0y/CnxBak2ca
bROiOQ8XvMJVDF06WZEaZuN2KSfEI9Yj5cZFFC1sxC78Bd9JXpiabtQ/MfSqDy8hehoqCrpjzk7F
Ssx9jgF6/aGBzK64BtKwxpDyXhsMNuoeSJ6BJGA6RlqMGdHv6T3ikboqXUJUyXzd3K7ZaZjIdWuK
2SG4P/1QU+CQLcLxfJvpVihjJVlT8Tockx/7zyj3YWtV9Ly/p/NSp1kpskJq1RSHpzlp6CX3m3hn
Gyd4aiDITgk/vji+o0T7lFNCAx9yoS7ouegxXcjYFPArakSed+1CveWIqk+rCS8jYHruntU5IuDE
NuX8Xf8gV7A+eFHsCshCBIL/nNqqzPMZaEiDXAkISZuMUCHWgN5lFq1glJx2Ik1k9HkjcifkfdoB
oSmNJkxdPw/ewlevG1f+duwXlJXL1R77tApC7YAQLRLijVP4o7NmJwq1C34/Haa15Db7vl29Wvx6
ONZQ+e7sMMeSqFKk6XI4qBJuL63m1UAG+AMH6maBH2xh2hDnycWUL+CDINDVGPIrS1unNhNPMCyo
+PJsXx9zk3uXPf2lMkCEkf3J2UP+RX6DWoxDrOsRMuTwTIIKngE5e5dVEvXrBN/+DCSLKN6kLslE
H1SpvQHiHY2K332OlHtOCNU7fKSAd8nGgEd6h5qbjoExMDu0ezQDhjVECJ326s/bqPYlSl0uar55
3IDh6PNrC7vwNn8axSde9pfEvEE0skTbOjUqslo8O14XY7Sxa4uQkclOU80SsUKlpqO482KmMJk2
s5gx8lbq37gCiDSmK/J5iKi2FvhobhwnxBbj0HCOrLiDdAv79PwawGtPb3rTUU9kAKDzUlo9gyWu
zwsqFEOm1oXG+LuDOXZhk9/Yjc33KCXYQ61YQ9SiVZ3uN1AZoCUDwKFcqVo3S6tQ0sP9C7/DVLSD
qt1CMl3DEOwnf63o96E4liktukXq+FRcGnWL8Kv5o52q/Opzt2pNreaxHzQHT6sGMAMSmwg8jBcT
ZpT2mAgCeerSlzHDybwhU5Irs4VHjfGoMliK0H9nI3BdH+0pL+iWM2nmay8qydNdgv5AR0buV2zu
O95+Q9WDJv55p6oRd3p6AaP51iMsn2A5fMa1xyK6GaIx7c64+6Y7ftlHvyK6WVSiOrTvRSvLTWRw
lkFXy+KPqKm3y/XejexhBCIopohAzCn+kENdUD0p51wiIwDrKlNwudDTLiQCNlPrqvfEFCTtIMKk
B3xqoGWZLIBfYyLAW01szpyD44q1yvY8ryhWVenSLbuMBMNgLlIHcCu3kzg5xbc4Tioglu97mZNu
iQAFAC4mQVsIpvftgR2yjkDNAxa37ooCs+0e3kN87Re/HtJwBR+awwTZKyyiR6c2o3wb8Oux/0X9
+KAYXiicwAwCq9UvQnbQ+aoT9aH/NXMPNh2bZwQADoar5OGRscuAGH5vPE2snvtgd5Azm6yC+MpG
Qh4O31Jko+g+kYMj/399K8WSAxhzfLhQOYfSIg6gwLLUoqOE48lmBQ+0j72nX2lZ+jmGx5Fw1Wow
yK0DKT+KNqNR6cyYb1O2x+ucdQ3Vrr2X4624i2mlvJKUQgXXpF0q6PgPeLDg5Eq9WEceo/DQ4dqV
ZfvM6hUkoDw41DRxI31g67FcA8LpyoA8jjYoZsuv25JzYvd411+RnQJtiTNNqDyDy66z/DMZVYPR
/EOq+vZwa8z2VVvzjD0pgOcMEjkyu1/HEV7RItav08ikW8lGQ3x4bjwBeVgb/pa8QmW/gR8O4EZ/
McPZYSGBZO4Cib++scXZprku/VAb6iAq2h4S/mSov12Btneq0NyzyHKA1WcAa4vkkJvQl3ldSIV2
dsKxAv1eqbEM7goX3sSRKOlK7zGnJ4+kQnJRt4eN9Nw7VD1juo7FUWWp1Pyj+wrxx/1BBC+bHx9q
S9kYkUqSknczUH734e42oNlc7yysPvkbTzQB2iRkLEyHvfWRmArk2JhMotzu6e+BIND5RnnfBzk9
TAEDZL8unTAL8apMTHs6c6j7rPGFr7QcKFKSNJZxY8s3N8VGeeNPIusxSsAXwMjC+UG0SXQb8Mxl
NORCehu10wUa2HxGE2yLUT2a5PkOFz9LvFQpUg14zt1qtDTqkgFlMgI+v/N/+cgGYdlJnOevy8R9
e5+P+2CvTZvACkUF0i4p/mC5LVpdsl6yDI2uv2dTN77OOMdP/0gC2GBIHtTzBycljLM/eT2lGHr5
bwQWtm0EjeJrnyH1wnWDNR9ATSasMAVEQnTcLnmVqvhkES2iLjdwMIoEEIQwmS6LvjAcK30a6rLx
u8Ab5zHQxUAuGOp1K7f3qkADxiYqYTtZUQhiWxyXR5s+SpD1ML+p5aap81YjiqSw2cmhvcaFVR+r
v97nemD9HtAn6p808SAC7nQWmGjVpDXhln6lsb03kh2lJ/Keij8qGl8F/pQVAV8YdBZClmutYGc1
XpeClKF1oNhWVAH7ZoU6SpciZAfHUm0OEjvQpttfxzcLncUW0V9OY5BOEtwgsV7yK4n6B1MSybfw
qYJ5DImSTLx+zSxttoscI0ilELjaNFntHBziRe089YnepRGUSZFg5+U8zX/9riW7hvnRvFzrWoD+
JANgpbT4EEYNCiNkGB9w6VUyKfK5co5NY6qEAAcB52WSkE3qMAcXA5evV1fOiyU/PN7Cswgd/i2N
I2yaixF6SKG6eAgABqVOMqwrPdvDEBmp+X20//xDexeCCrAxTYzZoOmwjWafv8GImWqWbHmbQp55
i8JYePZl8iqO2Y3KkZ1yfuxHi1vav6BEmUXPyMM0vR0BVmmYhix/lG0wqIY/DJaN6wT9b6E8ai8b
o9zwHlXdb8wVhmU7rnpZwOjRqoB+QaGdjDFz/xvh9NTHy/6Z/4Wr5PWORDv/byMyjRR6eS6J3frY
GawyleQS9pj5r0Lt+XQCzVmFmwdTxaJs5A2BnizHS8jjwLvDyQeFmOQzq64UxNkxH1U5xUUMdM1C
DXdj0BO+kDCjLKpLBgt+vIMTXzYW1TTxYcWlCkyw/HI3XWgub5Gz0HxmGjR600mrb7NMJ7jhYhIs
gQTOvroWWYxFHcSHrURRaMQxrJGWMcARyXAsfZditTUde9wYMAnJbNFnDYSxOZgOkDrUuj09hLFj
66TF+CDTZXGUp0zcsl2XVqTTwngWEZ2HEs/GntjfJuMCS8QRuzxrtRzqil48em9xHRfcjkyoBkPS
7DTsGTizmdUTxIFWZtxBRBwDABnqah8Kkx15C26WX/Fc47EbLxo8kDhO80oqPcLDgw+7g4lTsN/z
StYPuj8axdP3w8hk+3wSyxBAGIZmclLCW5YGFIqokLG5etqnNeZUoV5Z7IEL+pkiqpqNIh7uZRfZ
lV1V9L3zVNrbZK023iem20wkFf0agxkLvb+jsEtFPCydySBAy7qrAICEFwGPTf8UZBYn1XL7dBTG
rAyl7Otb1vrmO8BE68nC/5Nfoihbnb/xiLcKrqvni05/bxC7WdqTHF4abV7vA1lUWnqpbE6n6PWE
eqlWQIxbf7VPlWdYwpm6sjRx5rnlRmhIpZLJ3s1LpPzKILjbd54dHmlEEG5rz5IgmqcyEDUStgYM
EEKdWXeb2iT+0HZKPsjZisK6jo7PFLgUNNXOShAUwMpIK/t+ahUUY08NaJodzDT97toMfrgKDf5O
2mvzvUXySnkxiu4bv14pRrUNzr/1OEYFx83nHc3U9HnIN+qALv53yxu0IwYfHtsWbW616V6/fvq8
yRW45SfovFRSTskNAsC/Zt+hTY7tNX3I+x03eAAkrxuNudcab8K/R/AV0OjzIlGZ4hTK3fE/yO5c
Es/kIW7R98FUUOPAaHg3PaohhI/6eIF+KHn21zc7fuYBLSkRzLn9RCop9ds2yU6N7aFlSPBm6jdH
YcqqHUKrTE3Lt38R8LjYkNBJxFnI2ikbUZ4xCdU2B6rjGxalW8xRDH1H6s/qCAbhkAsqpzej+G7y
kBjf720cmMD30I2Sgt33k2EEN4ZQx7uoh8EPJdDoRqC6QL/M7upVDp2whhpK+LswOOZH8KXfK+7s
UDm3ScE3abZ9/tvm7oPqurd8JFvCvSg6qB4t6NRUf3BCtA3bOVfcJkc64M3nHpp3D+iyW7d19eGc
C2lWsrF/koGWqCq3qywc/v5rQQiM9E+c6DoWl4aP0IBC5FyuhRLMhluh3MQEV9ky9WE9ll2y6nyb
/JId7eo0V+u+AYMdp5t/5Q/7vd1mj8t7LA/FXuWeQuIF5y3tLSybd7wty7liuMq+0CO9lQ/ZUI20
GkLjyWy3znligtcp49zZZwy/kT6Z2nmvPJbJpiq8KaxixzpTyUDZJ7hjQj5z2zqtwQOYypcsmDdw
ttqvK0/p/wgl0Wm4/fgSbzOqye+GymUfxUQel6it80uKbARSpS3CmZxEXUTnXWlhFVH1UgUl5MKE
3QE30MGekTip9qg8wM/B8ycDHf5XU5N1UD6xGsfN/phsIKBifR9cW6uwsitPDNiOf9RA92CFEr/W
JyQMN8X3vyUwpuES4yNtCFWEXvJ813zUzbVDk3V0iVndFUULAJQb86maIrxYUL8XqB1ui73ZCt2P
PjgqxjJWRPig5FT4uELSnN221xQc1EqoajI4CxMEFC4+S2eXUJ+5zow+x3tWFOzyaItPPXSABDOW
+BjcVoXzXOTqJRndyp3OwLUvKESZOI6xE8r+UbWgmVzmEaT1+6jSptIHPgPpG3B3Qjwg++4uNxzm
UgFjtD/8BBQsECjPrc1njqx1FuUWeJsmMnF7JwX/8sShuepHeQl2jAr8PiIcBTmrycy57EJD4v2u
tG2gTpsuD0J3zIGdp/MtxsvVOtB0srmKO2f8E/HF91xX7i7e7xAUONJ7M0j4+jZnYeULpkRuWTqp
zSEA5QlkxZ57md1tfgK3BLtQGD3J78jVRM6BrsVT8TJE/IgM3TTKJ5HRkjROVF5GaVP4tSaCbvvB
GUT5AWY0Q8KPWYOAmdto/yIr1YxkVs/LN9sAZvON1NDQs7CRRG3B56B6BEj6MoqxeW2pH8FqieKY
fc+DpKErTuxmqDaaOUDc+tVo9cy3IzEbkc+0QQcD4a7ICzKw2xMbhiSLr2+AK+sN/T9o9noKqzU9
GSeyOosoh4W6Cn4ML/1YLb5WbMXMyWcdFhOIQbDQoThVkJUh7t7ay+/0SEtzRS3pqjuSCx74sdVR
BparASIBTc9PPEtD8Lq/rFJolSFeEcyApN7DwJ/2quP5ZCEfAJIIRTKaGLO0dd6O3COCBbKsuErn
1+bccLU52rIFD82b/+hf6N/IYiul0MuQj0tEhFAsg7kbkhW91YTzkNQbOQtuOsbuPJ90h37EgzAa
ow8lAIgjl6S0Mosb/cj4Xh/BFrVsSLRPGR0F1dxSK0x+LOiNBOKkjNDBxbM4kNTUoAWif2idhlwY
WBhPgmvm5ie8/+OBwF/oTRCoJQIc7BCsKZlFsaRFhOk/t+SnQQPIqPE8t+xzeBoyetuc1O0kthdJ
AyKjFsNYjTflzLhYZQiNgZtj67H1y69yU36N1OXBtg1xfsj0QnPwS59IkxzafOv81uDyoXBstGCn
itCBttuRUZn6Cid/5q9y4RuLVtF8/BX1X+s/dX0vFNFk0NJkwE8CBwq1kPCBYc94fXnSAvhnaZvi
v5NNoH2kcUUxjVcJS55ycxhWwhMJ0evwOeHCLUaMvx7ymUiTobW/rxXRpv9SIkdyxZvmX5j6tmA3
aQFg6UEC4q+8cfmjy1yFRCz+74PNOC8ftCxVgkde5hw26umsPpz9euB3JnSqjwek+yIeGy4q8hY4
uMRMvm63HFhm6nWgu/eiXVZVkaUqHVU77e26Xzo/yOuA4RQ5Rj1UKn4RaJapB5+iZFBD5yFlcTYv
OHqvogCSS1ZnmAlJpwtoA0/zoccp8DhTc5PTWb4WEUyeFSY7yDUYediUjWHX9V8V83Nw4FGm7+34
zWG5H2MDAnDG3TchuR3XQLPgdOvQL3VOi72lEwrQhVDf9XlatTYZV5mSuYivIOGhLfHk/NRAADVx
olzWhVDfOtNo2VEOLqSQJABsyyv3N9Tn7iZ2MpID83n77reI9/K0UQzICmZCRlkzgNJvtfKnEU+s
Vb0LCsF/wZ0xN0BDdEatFnO4IB3LmX56lbUzyU6siEUR22lYyBlHh7stMZfkdqCR+C3mCXGI8lUb
U6yB51rylVX8TaLmxdULZdLuWVmaYcv2utTAQnk8murwq7fDd4ZB4JYOT8Rd0Z7405itVUNNoCZj
rN/sIJ0bGJ6fFlBJWC9y+DzxJGT2+2X9797uamlRBxWzg0GifaTwoVe6k+vZEd8KlHtSxlSl+Ntx
vilwWS9QP26u54QxNKY3v+NmP4Ffc7a2GUpb1SvIvYBxsHta/3lOspG/aPc8M2xkndaOyl6DF6UX
0xjvAx8ifAjVSrOFsFDTx8TpdwhVyWl1QIu5FL19WRbocKpWgxqMOggfVKK1tM8uZoDX2yySKNQR
kFC30iyU+3xK7ERJ11syaWqT4lqxA7DRQR4LPhAaKI5aqV7ofmHvRPueT2UlUTibsZ4RDCpjWhtQ
bfAhat2PvIF8QZWIWt9i8kREaXYhHBFqMRI1ny5VLgBocoyZZdNarKybS8dFgfJQZ2/Ywjv+gS0A
ssr5Hcm9cNwcBc4ndhhLjx2/zpKK+8SHowSsF4YwnKYh22ukSlDLvMBxj69E7iqYxxyMOJmo5OKw
M4zTgQuLI+3ecZJ2/e+yHWSCMsFWZaND5KeJCdN8yAKBqc4wG/4hhx/mEAlpZCUkt6hLhwqF6FsE
ObppH2hsmdBd03kvmPxHAgw37tJC9P4pHaIOgkvKN9EeF/tamAZ/OG+fg3ZvJivHXR6rd7jMFcx1
KMWI6Aj2jUBnIpPCbdSVyiIxnPR8rvm478c5AsJgL0GclJ60rvZY3YMuZI94elwNUbvDbcuXyiaQ
ZgCYcGW+zDNGc1H9oh75HthVK6eP6UOdkXbptavLORrmFq5Uab8PkzNeZSw8WMVHMAHWrzKMo3N7
EJKAcG7kJIOo00qlmcpsJOMw4X+2em2fXT9GzgK+DFfLBfMVsZ2Ew6RktszAafbOZ5H2cxxIEl2j
+zyoTY8EP9lG87glnInoiapEfZpxrK4RAQ0wVFRuBmVhZEI2d5Mi15Tru99L3NjfALxlfOi/PIzd
KPEOQ+bRRZSlPRCS7lMDNDMMqGA0j0eME05MBG00NPQZunITQqMHrvawpJKRWxABtKUp3OCvMzE3
aqe5KA8iN7O5b9CmijHaeyABFrAyP9T8A/5KRg+Kw7JGlD0FwgI0ta34XMWRFNAkZdvN9sW5Ec5x
32DzVlkfr6VS+TrjDox9qcAd0PaxliUBcvVL8zCPweyhZsip2UKbTQiF2TPUthv8shcQZxz1B4C9
nwwhK17D6TRiy5u/z8z+U6XJX4PCFK5klgI9/kebCK/avaztvlphVV/yWvOkkkIL65D5gI14Gu65
Qo485HcGKIsHkN1hZBfme0uOwPnUau0hkdTDD76uyepFMI/7+YYDMFaeU8rgW7IQwwapyptGHCgs
FHg4BKaO4w05cfoT5wc5xhCMZCxQAGyBTDrY2Xgx+WEjlh2eJTKl6fqq4Rlr4PMWkv7W129wntja
k98BqjmeZeNSZKVLt+8JcxqQVoq9HaXX+kdzwA/tjdEm3Il/Z/EEkMwEx8LihLs8syw+rzbQvf8E
NdCxNzskxGG/TbCzdJgD/7nXjIFaX8mNsQBGRmmAFo9+O3w+fiG993+ynJNj+Z4I2C7wOA4TLYlC
eBLIUK9LPBsP/Kn5GC+F0voSff96pHvCdksLEvAafF4uR/ZZEhGIb0DxSpoE4flZWCvW+xNTeCiS
Iq/uuIOsDACPjw44lJQSThooA+6uJxc812P1JwmrQ08hVa1LaajssTVTXWHA+ps/kTQLZV4rnsAR
eu9Rc/ZbQiL+B3DtkfBpchBQcQM1lYlAyQ++TdxNQuzx9H4sYz2iNz44gNNVvFbhpsIhcxxgVawf
VbYp4P7BOaxKx15+w22qhl5vYCZBMWJ8JJSOukFxrGYpCg4niCyNOrFfgPYk46bKE47FC5gwjmGT
WJyCMT1DcP6DFpKleRlEVefaDD8F6GNKCJnGTHqM4iy4H1NcIJHndr5TkbCqleEbFWoTbZ2pMZZP
RcXUZr8dykVVbeGWEAPngC2Z8rdz8+3vFGIeoB2ZnzkWBdBhYqFmWAuAGhLuiJAefc7szo2FSIYE
6X2NUXngKymHkPopM9rudtW+DMM2jLu/nM3PW4f4VOv5mY3nGb9xMf8yT9nH56L7Ioan01mMQZXO
aLvVGfyfX4iHfxpwg4gp0MDdzLAM99uJ9bke5TqmP9RF3H/8C2dFeuzjrVZMuVBgtnNMubWNN5KN
L1xEz27oYaElDvCq0qdv2PViH7rJzCHwf27hUMTN1oz4x6shFkwbuSm4IvXbSC11BE8ZgSLmyFz+
wRarGoTZeFMCMxVX7BAsEscVeSHIqNpSv02rofh/5JemSYan00rSLlaoDeRpk61jYIyFGn+tLjhE
g36faT78M3rH1plNZZsR+44w62uLElonEwYIVSpC01jfRxnij4AGhXl7kIlyEkyJYy7vmdoEI9PW
+U+NFAddDNwy/G7Y6HQjSBQ8v2iR4Ypp8m8TM90wobIVKpOif5+EaLpAt672Ea+BJlaavKd6PWZ4
MtyhkTHSdrrH1h9jZVbkpQ2d3h6MwbT0ttLVu8DadiIoJegNo61m/Nb8kV1G/c8GdxRkPrI93VLA
1YDG7V7tnutcUrl3kQR6sd0DXKvfAyPN7rH5xxayYepJksVm9ka+GA+1j3c2fgMxHT+u9H26WQUf
6tzXeGz1MfCxfP7QY7OvqzGvY6X6WKgAnzBk+/Qxh1ArtE+icFdoxUqCO4koWobt53r/se2lu+DX
iVZuC3qGcKAt9xga1PkFb/1W43XJETItKdp+QMX5KZ4+wowpr9FMYOyp3gtxptGJiPyEedjVdfd4
XStfsV0Upm1ad42sy6NqLORR0pWcCe2nB7tOjnTK1xI8RU+2WnUrOAbPsyjPuN8ZY1AIr5ystSuo
om+8oUMgZvYqwSUH4FX3ZJ22NhID9/9luhlbhTdTIFhSkFsA68hVliBLafHSMuRCNKmALRKwATHZ
UFomERrQFfOAm6zco90D5DER/LRIFQz9NZXtNBCo2bE3QnviO5thGFfb11H8VU72UOAuOpd8FkJA
HvGL1hlCRZY2LegKJc5q+f25TX/BQ5ooOIaKAtCc9CrP819GGotyqSYS5fowjnO/kB28qQZXGXRz
rOtVpEifLJG61snKOifhvuAWdAeVDQ0MD/mtclaXvbt/jn7QpLkWjRLrV2a+whingdgzbf3gTR2K
ilwVp0/hu8YbG3pXOMwznlkROrq1Iq23BD7f0YlTsJt1SMokkIms6Mt01xalAbc2gmhEC9q01RSt
c+SrqW3kRosuujL3BbUQGaOnclH9YHrY75+pKgFNsGZUuL8yCoG1oDaDDRJfpg3AYtyfrWvgf1++
RO5isUHcWZKruKIvVUlkVlJmIGNf7q8yFrSqV3nZpjVRSQBeh7X8OMIuQruwVrZ4ho+P6McjC6zH
9JGEG4WHJDim+9kqBm3z5cPBdJqWz3GpRMm8iXPafbLFsCWC7U/kl3Wcan5WdJ636h2dRiMr71dL
AyDxTKv54LwvWdkGAWtxb6G+tEarJChA7IabRMypvsL5CrMO6KhF+7dmxXm6yrl8GaohIoHoYOE1
ts4LUXmLvnxSwJCxR0fQ84gBSYnd3CVGeVkHLlA6nCpJgnob7KOgG8Q0d9RS1RTfqdHlNG+QpslU
2VnFaY5TYn7y5JeiVcYhsp3NO2GOZMByucPVB3cLgHk11Nb606LoPpbL1A5IVhkEdg60cX7X4rqA
iu7FOaDkelQJ6PgWPG6iYodXv/IQ3D0hxRAYCld4Y/sztVvo9i55+fHYkfyI3Ka9usubuHrdDonm
dpmYPrE55rFW9GAiKu6jAVGSO6gwlP/yK5AnZe82w0yQev0182T+calrq9KqAKhKGLYfa+zWsrhj
bc9vedSe5FGdxGgBS0vkXkFl6hiDK+iHuhsca19lGQW/7slvgzNrJ42YXWdoL5O7HM+FWDnmeVY2
216d1rTnOoWv+qkrjlO76zDbImHv2YUmnlGRE8kHFwniTd551RditOBffCGWgBZUMLBb6xuwtxXZ
YX/35byJIHIcaAG8RN18gJIerk0h7vmg65CRhZEbe0XE3NfbeGGkMwxeCAMPrR3KUrK287+8ursN
x4GtX5+7O6LhvXI9+8xXPllRW2puao2yz8b9JycMgtkR6A4FQWrdRYPcyDEHWyiXvQwouRKMUR1M
zKNgJBcq925JqPu2qAE1qvQRWLyUkQOvC3EQ1I7ou7d+IOL9Fpl+ideD2+8+Ei+c99NbwP8eEuEN
6Z3Q/v+QoU1tTfB4Rz4Kmtw0YW8g4lDnA6knr9J36Ulkv9iqWd9HGIFqpqsq0tJRoM0ewWMZcTsI
9VCbPdqJalchw/WHAJeUEeViATDD8Fp+djF47laXYKIT9xGY8GfQx7b/Y+6j60O1HL378nel3NjP
Xp+viFAmCkBge0n32mRsj3HF8gR6uWJtDzmAHopm2UmfJtLsKYZNM+fJxmszzUyb81djVBkAKd2v
Aob9ujBhFn3vh9Too8Wf4jGOIgtjXlr2fI5SE8AZy98VxHzlmzbMYCgo0sCHwsyfr8nd5MwUaGRC
gnPIROr7PTBja0vfpwtcZqpU6nu5mYRGwoQZpVQ90HyTBPclnU1InZPT64J0vjdLqjHe32I/6E3P
rCSFZ3c8owt7Hv/UQ3EKuP1ijVqw+lpV1tdOeeJFcY1f7tH9XvPRiO0tbiwY2UXG978cuqkHUJnt
hZfI5ppYhZ17dyI58uH3SAGyzo2bFDUOp46o7ePivCIw4Ozfd2H6WnIcJ/UwAtMTR7XVn7qzOsO5
VbGFSpPUWzi3hLnA/brfy3t5FJx1ExduSCeDKoLEtLOVnFfm0ZRwKx5SsZcl+iN73ZGU/3UCuf8p
j7xYDVYdXb3LlRRmhM2fPp2VPdA3DTvg3y43VJHOlRYPSPqcPXdVS9qBI9eGj8IToOWOqKWtVEgI
8ZWMnJVyYUYVzYKqACSJmiWk4JGD0it5vg6q4hN1iialdgiyz5oRmXcBvYAwmzZ8t05XSfVvLH+1
oCgyxcBLmOgaNAiKr0UKXzK0V902MGgZx8yougE3I7A98V+yUyiZg5DA75bX7S9T2c09X25I6AAz
CItvio/JodmpC57tolnzY0F5u34+yBPiwTNwW5mpsrpxQSfGgIjRJ7onEIETRVotTPhkz+l58C3p
zs7+lICM3aHhW5WQ02a3RhKgXJxLz4OHN0jZ5ltMRkTDzjqUL+YqGlGCP74tKKK2GHA7/MdXDcf7
Rmr4P5iipZZp9ZE31I/HC1S5oTTgc00x+h4s9LPV+QHL6spdQLi2JBVJ52IsATtUblb/pcSidchv
IYYbLPNmiOIr2xVHg5KQkqJyCBglJDsXQged08lQR1xASi5NdJP4lnVN1p51hQFTQ59Az1IUal5/
F22pUQPlgpYmy8sYC5rAvXaf1yhwWUA8TAl+5O021W9qGKO3DlxMd6Nq+dpNCcSRYz0sRkL3eBUF
jn06JXg9CiuBytibJR9ky/KaMRvq08vNFaKaGLb2lzUDTvhSpRfsIh2Dmb/DckXrpgd5hBVwLSrB
Fjujos3JN6n3yqleC0YC4s7bC7sV329uF0ksPtKGXc7MdCuTSaW0moMSWaFE4px1Xr2srkTScRGM
eJCr4cqNQg4ThjrgvnPG7falOhOG16GIUIjlKzGKocm2SurcDdbMSY7F/MddSVUj15dGN3D16HC0
QW3Jk263O19G6ccN0ysVl3d5y2LD4sNrfU1m1krnXYHIMKL7P4perbnNaugDS/UDH3S5zi7rehyv
2f2vP1+k7aKS8OPMkRRJMdpabWv1n/Z7dZF9yu83MVN7Rwqyd/SpBeoZvJbyu3tuhTDZjrP81+4k
oBvd/Y7iQ+umiv9fanZDW8sHdvSf69oIlk6hWpRVljTSEMgA3bq3I6FgBQgmC7ICr8s7yPihrK24
SCiujV1IlGkkLoeUn6ZNfac2I0Z4C9bBQ81J6+j5fC3B3TcPJsnRBVjiqkDYrxZ7mm525F6Fu2K7
D34ygMhWOic6wa2xaT6/6rzmaMmC807WISrIY8Xgbaaowwwg5AnQ//2/SkxRqD5ZaqJJPeo4dKXa
L4xVR2gn6qyzgJzicDx7KAP0QxBvI1iaD73eXPIvQLBTXJkdeA8UOjo4x9A7wXkk6DxDS8wcynJP
3efp3WKWJKZTiBGJT6HA5t8y1MEkz6U1uqI5KP22toH5LDt7ud2VHW/w2ndS4eCReCE7WlVj2l7v
zlP9f+MgjdSBQA75Tb1OFnZ67ber6O+/yVEFovESLJ9ibwuqssWJ9arahFdZsbeYl8HSV7yxVFvE
gkS9hgjF8h1SmroQx0cSxpPCxMsPqTOMk5ufF/SiMjWBV+j9Pzi5Fa80sFTBQL5syT3W12LvOAR9
xiY1r4i10Y+/6BCbrL7ucBZsXlVfj+wgrFUlgO20NGUYiLEmzgCrT1d9FPh2pOFJk8tt5U+HLk4K
7W/7HQASDdCmjVguUbXi820rPf8BZ57EDCLTudriqsoCA1xMd75T21egrQ2BNVhLEBUH1PQ3/kP3
uqCjxXdMvp2EeXytqhAPuXkwLerM/DW6S36CVL2TrxXMm7fktLHNk4sxB4zOqO5YBvY8whaW3Wzc
wvDeiZaoEEWgtm+2/2aQtdLPXFI4+ktCDhS+NJ3Bizrods2awLOVMEX4YiUxWSfpAo8W5HBEqBXy
1jEb4D2sxNwdc6bfn+W69yqeNrj38jc1HaTBnY/HmhUfimp/M3MP8u+/EXdJ5AHdJOxsXUOKwz/R
ib1ZKlPfshyjU+WQH2cWfXSbR9ksW1gcLRC+AGerfI7rqMTAmev+cZ/6shCkk3jPztSFzeZRxAec
zAJKOrVhJz8nREyyNIEyYVimp7m2rcBnn8xMMUW3wGxQPsS4h1OYaWc6wr3WLFm6jsnzHual7Mp2
4UKeSYr9AIPii7hz4LAHYdqjnxAEp14swnIa1AywF+Oqi/JTBE4Wojst+wG4D/MwCZpiiTiFe8WZ
psTNL5Qg7SJIscyMOynlO+8dxSP4kxh+pyrWIaf1YxnZqzxIb6YrkulcQDipZxeyKeCjSA4gRqX/
bYd9F0/OrkAknJPWlbLL1HmJXP9903umsmuAiX8axd5jM6KtODQ2csvNOf+4VaNMmNEUr0DhsCy8
oQcTJcAoS8nUBv2azRb+LmxdXdPXxjiuRkYSJjeb7vbBKY8KY53qlXaOKVD3GNUBgq9OK8agbfz7
u7Pw37yobIIl2sTo7s0lULye6gPKw8mv3bBWWYSHKoRcE913kbt8I46u0teh7vnK9KozPJIbXk+i
Rpx/XCmeY5KoqTOwbMGQF2j0LM67EZ/zkdyvLOG3JNXMrD3o7BzjLj5TFfbELBiQSRLgdfhuHsRg
rtQgWtqXDRMINn0CBhuwtOal+P5neV7c3/HrsOeNLb3AyIk9AMGkV6chN954RyOgEmPSlGVJIMgd
KbArNYQYdx1PGeaclFmYK1yJWbMGaFMk7z7N24axFcgYFTJQx26g0HH6zvlZHH8F6pB5V7m+dJzl
JdcqMBwTGObntGwcbvgh8eJBZjYZoEUPVSFJEVtIJ5FxZcZjjQYJsjVJ9fX0Jqc+iQnx7Se1nWJd
oIHexpWnmjZ9y96tNxna7j5h7EPA8aeR7y1S0UjXY+DUHAuVXxYDGangtIEUVUwlGjGb77gT7u0R
LxMqIoV+P2KThjDWvoR2y846ctqTiDoR5yadpgR0N2VOdYmyKWccOtI3+ywEqfgC6tjrxCXbjtDk
wqAPSAMNrQiR2RV+ydKhyBiqWs3qW6dYHx1GgtMdaSlzgdHLqV6LBouyBhv5n9+N17+rBO6V+9ro
GaL7pRpsH/66VtKd15XRVaBMASi7m+qd0MiH5Kho0DbICUai3tG70G52inbQPVZXs96naVU6JsXF
eWODqxWwTx2IdDSG/XD/3/QhN4iqQ+BqxqpUAjkaQVwmaejQTseTzpUfnI1DY0WyBfa2nJSqx580
QiJDi26lxYMnRCVip2KEca7Yt88PvsfAgUfDzII+8obkY694Y91FKjCGig+tEkpSji0JZjjyaYbj
6p03WlL7WjwsfuHje1QN94Xuk0bnG5EgNkTKwY9cSlRFnHSoTdx/nH/oBV8MWrCPj79/BnN6lUjv
wX4E+n4ciZvc039jE+n0sCG3JriLI9KyAD24Oi1gki/HWtObIBOy4LnYONKBTXRnpoo2pQFui5qi
Ydd89NK4rhw+ZvDkgUdK7mbirqYSmIvwuC/Vwe2vlYWPchkNUMTMg4+RaS0TyQCwSH+V9rDBnKnz
bpu7Mo7iQHIHaXLMqtDNrwIJSL9PZ4DlerBpW5s6r7h1RL12g1a/G97wwPgmabzN4jB+vDj5810i
cy5G3eXq0JroeP/BKjNqtxPI90wkvE/8o6CZqy1uXLROpySfAWjGn0LYwp/ginSc0W1G+ncjrdTV
1KmX2LvFfKNMlpvjKmwU/9VV3YaTlsQ5e33TxySrWh/Lq05NpKu0GAfhpd72acFSVsPr4LIrGFJO
MTYrCkeMAJm+D/OtXxd4WQqhH2fqVsdtYmq3ixn7JBB9U3EFf5l8QAMIG5QHBNFTnR2ZT5/Vn95k
A+2DviMDddcRqb81dp44xukTGYDWu6erPbKAVf3pLvBDROssOp2U1+O0aFyeTyRPFWbMxvZb38us
KUhuWUA7p0lH3/RUlxsb5G05/lY0UcLAusQT5BUexFxuVRIw1e36LehS6hv4o52mC7qK93xc/nGz
wI+6fKCGoz36tVvFSgd0xbWt1O2kplKRUhaTrPo5n3BwwGljZhe28AYwp9OAqpBtFQXdo3M+CrYe
GWOoc2uX7WtNd+/QkF0+X/Qx7O5ZyyBv+qcmnnIUSgtk4whrlww2dAC7K85l7dq7Mhn0yKKh3aoC
6sav2kRhV8bkSobKNiS7GfHZ5dSKprXtMknmVWfWlldF7ZegvFSKqoyR0D9RLbUi00lilbKtELrO
Inw3U/F6nLfLsy90hsArOpT+Y5zldCJ7MHbsoVlmWuVahglYcqEdc16Ho7475plT/ytmsKP/h4gq
5/YA9+PorWMQl31gtqkXZDe7kE6Pssp2HcC6nDJs2MAHMFQilCtaK34lJZt1N/F1r8GyVuBWLeSP
/wggWf0n7Q1ObOSnQ+ZYtFXLgixsG0EsMomUiyF2dyf0ZkMGNObD+jNa5BBwmA/f2RiA//B5ETH6
xgZEE707LWP5lKKbnX2d7Flu2ehAMUnpZtKyWBOGPppgTsR9O3aYligIblvxcokeRAGSeNaZuazE
3JcHcZYUKSa260g4cecDjW2WqgU3h2OLvfJQXXkbp+jBOKDH3kS0iphDHpkUF8faaryBasRkH8lO
m9DolW1lD33OyCCw1MyL3qhfIZ19WMBKsE8TuUAwRj/S6P3idjDj/taBStQyh3d8Yo1Q/+hrd+r+
f/EhEqcspTYtE9d54i96+Da22PlEv22d+XLPv4EQhmmEgsLqBEGNyL98mlzSLwHhamm1NI9RRpZt
gbOFg168Ybexfqq1sPkS9dRY7vAe0xy3m+MJzwXrkBM4iZc6tiwAbK9qvmPJsrsf1BdJDsZ8UpVi
KMmRl4ZO45YJe8wZ0iG6X0Zq+KxR61qo0n/zYkMRdQJb9j+eF7Y4x76KLvJFmOSDa8TplNGrH1Oh
QVoSMgDJBd4v9JuvJRDr3IN6X77x6z91KNqiLGfl6J5b9q0aUAo94tvr9l8BcUamZVM61KaDb56j
IsGgmsNEfkF09IdYGX9d/6j//rdFF1Ggce9Bm8/0PJjvaorlgpGYmsPahAz+NX6XM9Z1cTJ+jaX8
miUt+plr61TKkwGySdtwU0T2fOMB9uSJSCa6SCYO/KO3ZK+LcWcDPmS/Io7/rwQ0d8t58NkopNF7
eHPZ+jpmvjAU9MVNvf4JMnM6yIuhafU3VntjwSJ9R+m3HjplX6dKHpSynSdK/y92153C563lK5Km
Cfhalg1CYEd1gsOFNmdQl4XsbwKghlJi/dRu8JH+4qaGmoYNO31P84KaMPUu6yXQRq1RoLDzeKDL
9yKyQ2qS9qtNujiamkp2ZmqV/KleAg4geYdYHUajRf5iVY75WJ/5+q+EKv7sr+zd1H6EZsRDKwTr
KoZhzDUEetnQC6V8ZahzeT+AloyNiNh3Axpyya9fhURH2mUz28UWKvDSZ3b1G9wFDjLh4f/a5rxn
SW5peplc/Db8a1jexn/9OX6yyr4n8CdFutA50WkU6BkP+psc55euF9onlXAiPs/zy72Gmd3q8Cfw
90M5LrCYOBveAyWN7xisCx132Aulf6XVtSTSQm7Q0AIZa2qmoQiDsJqPMS6bbOxBIBeB+UUQS25v
kZEKdaQk/xzz5iTaosClgOiTHWmm21oUJAijlcUEv1Tl6649TG1jYAwxmRd0gEyLuPNqpz2ngNDs
Y0HGzk+B4Ogj52z91kZy5Rz7Fu2b7kPyabT5LGR82vc1D0MmDjRcnhvesnFep2vc4EyYZ8gaRjQs
fwo5v00EX10iCb+2/dvaTA3sZ5q+WM/3rGtgqiOXF6QiWa80tcu2SWo65i6XErpqOeK1vimczIlx
74CTWPnz75yMPfVwKwCLQEQ3OsUou+/Y8jL+5w/IkUHmpUOkZfswXqTrKzMD/5Na1BGzUQZC1Gop
aaAHexnk8VLfwELzrdnMHXA6Cpamux3MHxwN/u8pM/DvPf9onEQjP3vy3ZBX/YPVQu47vRMZ262W
cP509+g/HI2ZrBhjz2h4GF8kFYI763GA02fXFXaWd3iPJ8kojntu/4ee7mpIgUFfz75SSKMSZxGY
Md88SSoPanDyTZ8OUH50Zq+QZRWIDRxReVEM251uJCIwSwgN9RlH2yjmN+jcjGrTy2ZUWfC8PSdU
E1XQPmhpova9Ra2lOa5Epwo3pOQFdb8hJY8xuADMmsUAs8rkAnGVPv/RViTEhHXB3D3QeG26wfn9
ajpP/UXkOMTbLvYOUe5EbzIjWZI6uJbISym/7Q/fIhVzlU2q2BV0bGfT67NTptiMwAX2BE1eT/Km
8vEGnzwf1WSACVnVViTv5ZzT3rH1DL/vh+OfK7won2gAXTID8qP8LNBABn2H9WNmBIUdctdEkgra
9PrQ7P9YXMNOxlVW0CyE2OfJ0A/2mbPvwsP67kQLfL2AbFeRh+7WcQoZhEIFXWIYttL20uEhe9Of
AicrJHpWryfBzcOP6WmNBk3M4r2jyhKXoBVPJHM9sIEYyqpV6i3dCkqT5DlyxS8rrd9rWgTnzFf+
8rfCkWsXWaAbfIKh5p6BkI32l1uTnoQKL0X2wg7kk7pPwB/8IHajpGQzGNX2Wo1+Bx0d8Qwaa8O5
Ai3zm2Lbz3JOymeaUMYvKjuoZ8RuE98Cog4UZg8gkqIrD6odGEiNgxiJU9GpmnTvn02askfm8veC
zrGzgs+V0gzonxas19ThtxD0M/XmwXv8KO3TAIt7MC+MH2UvH75VNmX4oMcJyL84njN4hW4XX9AK
PaFSj4mmElAl+VX9azLNLJIPwKsrtvp4KjOGq0rv453YjT4gASR14k5e9WDLKPoQPfpodHstRW1L
ajLWQB43ZYVKc0ALL9EVkqtaN4eMSgAICsqgGXKpVtDdYdy1FtNWvMtuLdf3TsHTaac8Cot0Lt7T
ozOCAs7pAK1kjlAnjeBb7nWe5yl85FPDQrKzZDZakIFLc+YSXyHbXtE8owmMbUBnjNDRLuWnbCZo
/bXh+aL6R/36Dz2H7srYnOozQ2BokBj05SW07srLwmANaI/Jo6QuV9JkciGGDFH6Dc0AvWhVTiSB
1+hvG837YRk9CwiBuuRaSW/NykA9vFnh7/mHN5bl2rEq6Y5KWBW6XLHDdrjeHATV54gw+LmRcGrp
ghbKRR3lxbSDmlqvD39VRd+YoKPypyV43beFJs7jBYO3Aqp8iFjF/t4x7388ZBO1NEIzGkzry1iq
8163Y6f5qz0lZEflYtvszWhOxzoLRXxRC8yHPTeP3V9Y6LO2/fESTvyY27xhCMsxACaKrLuvNBjQ
m7AMS/JFDlYsEasRz8Iq2NmjzvRLmoR1jwuUFJa3jacEfhW2KyBZ6zd1giFvOyYCAGLeY+KF1HGt
CikO7I3ngAUMjtJTtgJBY8qePEkIdRVbd03mRiHk8jYhvqY6Pu2cRerviZ3XMe4S82AX3arAV9cA
Pe3HpeWBGWjacdQAboq4cHcoZAvmXb/IpJFUyTgALGBybpDh6ETikNjk3YvbnX62XHk9RYQXTpX0
L6p+lmtV/AeQsHALjKJlvwRT766GlqbE7uaHCgDjY43NHTLCgj/BS0iEzjl5zZGKWgmLVZP1j37d
0zL//+mICKpYK3zaB7TdTZX3sF1lv+9oKB+gEMsHI9tXNkRqc2BVpaa0y51fMRfwgwQI8u8Pdk1v
N12O2Ir1XUxXpENWy9ClLK7ymJgZQII7yDIVa1RA6fXMvIN2X99SF8tzNo5EkUXrjOqEi28SLRIC
A0vEAEmXLnZ5r3E8CqKNwZjfC0aLDpEqZtBD7E9iNmwJW8z/82ouzjmuIE9pbcq3SgGa45ybfZnK
MSVM7mruqaVW+hBbum0SB6h9uwVPNbAaJ4j2XJAjO8yMFsJxkMA+Vn650wqzi5VdbSFV8NkpjbtT
oHcx7B7cUYmiCnBaP5gJiWnr/KqhGkTfLm2ISI5QMpzLc+6PieGCBDSWqvkaGtQfeU+ohMp0UH6p
qxxeRcTNJ/LInx/3wl8abv3h8R91g3IunWKITJLZtQ6cirpxjg6HWzq0elAIKrlTqLdm1NuvbV5k
KVxVfYotsK1K2af4/SzN9x55ysWjK3MTqjlJJ9bQCY/3Y6Lfpwi3aPwvbl6nD60CYIg0KmjYwBtv
f63NYH3VAzu8Fzbcg8OzTUjfnMPfFKcRfVJ8kHvyWt0pQkx+oB7XZs5xTlh60u5F1zKVuET8ZAaM
gL5iEIjzvbx9befSl3DUpz2ko6Ujw/SorEOEg6dq0Y7Jvmpwo5nmXm5jlviV7NND8LNJOR1kDJu8
jxEZH1fu/devZd90ae+NEf6stzHgK2du3HQRHtTEwVpM+ciyZApP+q23FjFfkDMgE9WP5aA4Styq
QmGtnlsSQlmKoOgm4m2oHc79M9vor+tfuMLzzUVMibgUYFiw9JkhkjzZX1m0XWsFZRiajVBBwhMm
e4pgs63M9SdZQWIsOLUl4RAPdBhjqKK0wXMNDJIhBePCNpy+X/gNeq/MIdeLdIpHFIig4DO1v2Fu
Ki6XdzTGARNvw0YWgaYRoiMyr3N/l01WUFFBw2Gp0GrFKOlDurF0KdA6vGeZGjTXwiwKFlOBVR8+
aSCz+Gnow0sO8PijkCaAzFCEduAjlaZ7qd36dKFYnmWEVPVJtrf63/Gq+OTFeoRRNHY+iv/qcx05
ucsfCY8zo6NiobWP/LneASRoou9ODzywMgK0DsgdkW6tRVxvowJQshkVeYolRKnnyMBWRjPVGtou
0FzS8/gdBjsEx9Pv4mLgXlirxB4bCrQdlxz0d92z0LXgOlcplLxPnv7uER45WibMiLrzQE62ahw5
aARYAWDIQTjKrQHxRym8MO2BhckW5E3PppeoitB9E2k671p+pP0wckItSE7tonz5iDqh2q/2SfYv
GZb6wEzjj6KhKBctZOR+FisS4ydB3C9aiw465DJBy17TwvKYLwYHTiUk/izDlGCufyDtgManxz1F
ptdfNsCxMIvOMlbVxYWZs0FSeKXvWrSUyfiwI79gSPnwxCDf35XYAbl7Aa/RpwucgrRwKKNuOeUH
g04ropSjLIB3CjLZa8Kmbjf+GxrZrYI/blfcokQxA12G9JOnmHrxyd6u1eLec2Eop+aGwEPvPBDJ
qnXo97Ct1W5/qj/BTpPKh8GD3DWmuVVOza+jiPxoRONhNSED4avfxPXEI1YRFm4TjBulkAEqsuNY
44sev5ZJIz+S2FWQuQtsgp9FxF5JOuuGXf4PIvWDSveC/cO1vJTmJO2fYKxfGwey1+p6ZCAtTtn3
C6YId5IKDrEyCtZmnn/2pzX968mMI2oAAMF45xn4J0lhOdUKOP96Man0kVckK7MKjs4bpLePKulU
CWjzM0+iLovZaBMCqBA1MgCIykv0CcsQgxdpmN6mQCQBCagUXz7xG7lv7yCzjB9Wc6ueUQGfTsJB
F1FLuCG9Bm4oVNEpG7RGRUyuqdEDnAXEsJb0fMqTJS1fVrm+tqNDCf2uEgUYilUNtLvXgnatkwFP
LdDpkfDGZvNheuOMhuvtJIibc1bNhmvSfgeU0KPmxGZveq25Hzp0JFDkSCiOBX8sEKYKcX213syy
D+LgLlSP0d9NpFKPj32fVNMxqIyOV4fC9Mc4QIL+vgA1KNPNMxM1eVQzQue22ywhA+d1p2EtlljH
erk7TrkfDNxlTQIeF+e4n88UilGcLlC/hH6bbuldOl7IR4koNzP+9MlvP4RCM5Ok/6rvhCP0uAMs
5kCU19VJ8inzOXO1Q0MMqcSkpW/O4jMfBZQDOZAwaJndhYMX2ZWusz0uWTz3j6RZNr/ihqMJeo3x
xT6agAd71UAkU8nwCklQVfndgZdlU1EfdGiQT830ymlTOvUyAvtbkyWMDk4RzGscQWLFaQGdg7w0
x5Ulzp7cXisUA3Nia31qP7Y1d34s2OMaZhcwrtoLvjbr/gWDrXMTNiYXJguCCpwWr6KG/dlBTmCq
B33VoopICbUXI9+aDSgha5vNlMb2b7HEYAtNXBWTl17DsTG9uSzdogSWLQXMBDwMM6rvHvQSru4c
MX3ez8OoipyIfCdYecAmUgYziQtQMB+pN7tpJ21YwfqgB5WAN7ypXWyKb9pD5blZT+TMR/VtanNz
p6xanz2XXgTrVnudzX4Rp/txg7Ayasawr6BLT0Rm9EKdikPiYbwj5qUXeCq3U0aSmlDjV27gbrgV
D1D4xhhWx4C1IRBgwtIjUOXtidEFQucKk1pTvfH4l65N5HM/+q62OaGFr9CUwz0iCH97l1Z/8oGD
7aMjG/3TCvSza523xLEzjsaVCNWeHxBHtJtUYPJ9bkgv9yTsefPJWAGZeslFqY4H4W+nqszqX8dm
z3+qmzyBBQs8OvmvoRT+kn1vKyMFllQsr+HPGZPzGWjPl6tUKLecd3is1drjx+nWyK4tCC8NJuuH
ofOxtDYy7waCph2tRItCzcIknIEx3ShMdg3HDwEDEUeSr5KR5YlTJQSapHWjjmo+nVadmycSG1Dn
QySPx7aThvbg9zCLdeZrKkWA2ayG+48R71RS7+w9MDMa4434Au3uOQgrASSyDxl01nHN/qAbZdU/
1ZeuV5xpuwnMjk0u7yDUT75fRtwXGGyBgtUaZwCNZyCulinPBYY96bRtSRInhpkew0MzMRoAk3xb
e6rc58Tcqc15zol8K1Iu7Nq6TlL9SbXFQacAVK3wwaK0xfrjIJbW45xt3NFB5MAUE3GEqshYRzf0
qrulhhoK4qxZIoGCHUE12zCUtmNzB7F6QiizEf1uUNngQQl07A0vZLZZXeqLMwxm6jEctWvS77Xi
JStZJ7HQoYsiXSHsKIUj0PHNkr4+Qzbaz/JZiRuUXZLn541V3jG6Du5EleZl9JVfENE1o6B20Mzd
92vSrYB1X66JX/7tWiygODb+h7WXEZKJDMZ/5antCCaM9LfWQuCY5DK8ZDkg8DfT/BNCOU+YjhRW
GxEMjYxtUwOqCqP9OpYzGIwzNRhIYlDURwpGqb06u1Z3X5Fq1JD9/gc1zXplsjmK8/f+4CWzA0pr
6G6x5nAvjxdIN7TnWGZHNFeyXoc73GZ1hlE5Iupx240vZ5pvCNED2PvpOq7kOtbosJ7fBqmFeKZE
nPHKzsw52MEHFuype2pXoqcWRaJfImfkJWIL7p/ApNP/nkXlqQElCZt/xcUKZYxHiHwytNL7DeoB
dmsLTSEkTskpXiIhU42zv11Fz4IRbzqg1WKeIGNba19IzaYlBS7Z1OCc9RqubUOJyO05vgf/V771
HjYglUuj01X0v+L2QkhR6puBmatG5rbmX1IukeZMEj5XaQkwOww7ZTSKmJOwBsJNQWK52/O6rhrL
L1FBlnWCizuWajxjpSQuijMSxJ4BGAmAMLBV2OVrVZ5MLN4jS4eQSmAx48eNQeWexoumaANRmerm
p5kV3gFCZcQlrHvKvARYnZ3dGh2WgTiRmu6IFKcj9SuOi5rMdFbzLdrMef58BDN5gofRJlFJV+Ek
ttwDLkjTCpfdauG0HPkngJu39V49q3gIAdzRl/Z/7Ps0ES1oXFWsiAW8LB8g8ULhaEUM7gIE/Ci6
23YvV8H90LvKVJ591c+Jd2KDSc7be3EK1la9j5Erd17HiYeFueb+iLB+DH4N2tZ4EztXdJe6iBrL
aHUq+/V+X2lvdnUVn//12Z8/a2WxsGqyPjphjgd/RYrNNVxmNc86nPbovENWQlZ+wzn+d6hxm/Kp
TKwW0BG2XTLs9Pp6soYzcbEJuXO+4R5Ujvtaxg342FC1ZU3EybSLbgLuZeEheKpa0AFvmRM74xVN
D+Dr2Zft4x7o6KndJp5y5SfGPk1eZ3sNHZXoHjKXRfT1oBRrkqIh6hc3D3sYFTBiEffjgAAIXJHG
gpY9MVzMpVAQjDOWmLwSCyItCapud+J67B/hyfFJOdJ7I3hOVEA2A7SSRWhgKgVYMwh1C6GRWxNs
xyNR+Z6LyMzeP6VWadzY8gVTLSJLRQ5ABZqjdRQTusgcHG1Vk1NXxYBtbgYnjogXSQD5fBZ9plLU
FAoN2hUaEvkw5Cx06wN+gbD1dDYr60BQCD+VpGARoesoIpw9Cx61npJsZohixY+vDUwTgsRqwEZL
o6FbaASUjDhASBo7TABbpOpllA8rqUyiSqTCQ4nkwVWr4cjnhdFkCNbNXhUWW762IJBNH0X4bdnz
QgbaaDygfUdFeciB7RicDEEx4VKFLwnDEQE+3KT4CEIIAb3J4UNwpLqrTWiyw9dt+nN1P1lERZcc
Yr7btG2dPhyrRrEBuwsuulCLkHMqSHv9Py8zxP/s4IuKnHnmCiquybd2GibITDIKadPJPOMWLuvD
Xg+3YRnBWPe+rVDPgVnO91fw7z8HG1Xs5Lo3Y93FYwWAfjuOph+QvnZpeZxqOfa0ywylJoXsRiUW
BNnd96Va8bHlg6qGeVkukdNvhVLl4+AVOB36YZLd4r08nXEdKMpFS798CsUeUvg1hBE1wMaYLDus
lfhlkQcjMSiwe/gW41F9Rl9EOge+VeRTyqWrY+JijOA72Si9cU2xCUj0zQ7cNVuDrirTAriTU+Jk
WBmJdhAoQErHebMzhd23DAbHu4e79+QEKiM0ZkMc6J4OF+fCMMtdeicTj6FjuUk8A/i3Hi9zS6tN
CrvZo8iclIfySwr5A2BmgYmiDqN+neKv+8EI/pX2AoyfUvxd0lqTyXlW5BFbbhVI7JsGMz/YcBP6
YULYcEfX4a9kOMuoi5psuXLJCbBrGYu/T4xOhcFPrmb/pvFteVk4mr0SIxSI95qlW2e91RVL3X84
2VR81YjbuQ/3shCF333+t6Qkct9bx7Zxyhq3H2Nc/sKWO2qVwLYB/oQhwivULdNIjpF+LSijNzmO
2SEY1Cu5RyLmCQ6niKbBOGaJebWUlySWzStCVChHd2Henk3X45Jv1QF9urzkT+YKNqtjHgsOBqSZ
endimW969kEQY1NqaA72vNTLlBKI0yu1mLI9IbVkRWIWMlUjoMSIuhSE+xzOlLBiAbBwCCjcNbjh
tGH1yWsb1Ag5IkaExNPtfCVxhcIDSx/KDieT3A9g5P+uGQfmgyXAA/xCLTaFO1ah2V1JORIVE5Fq
skj8n//EcmPVh3SGCjpqpRJYsdkDepEJYTZZEc/OKbiQ5bPi/DaeAQXicz5yw3TjSOOiprY15pPU
tOkMzq79wsCyNt3WnSqYcBgKYY7jKgOVmUQcIc+g082rui5lCm2UwiNW7aJIY+RIL33E9zECJu0z
RXhaBqsOj2oCku516RoEy4hxXhclTN5yS2ZBoHfmMdRpLpJhpP6CRq7qLie5RpzIPjlc2lUEH1DH
cQC9AAUzuf+cuWBPe47TgifovumBThPC7Mvmj10D9KqAe67ghw4qWjKWAbE0Gf+g8kW/54LJdbpi
rTlIuQJRILLUhm1QWE9NLIg/n2TX4ZaL6mPhqs2IISu1SnYQQYL5W3bo1Mhsg65IXxAGl4zP/fmp
930os5zKJsDEdRMFQVSRrC5mpiyflMDvJqS1XwwMaIB/absMBqRjSPq9MfBd5fHTb8t0Jlz7/xIT
Z1MsmrDHSA0CyhJIXQ53hghwwZU8TlQybn0BA54Wg/IQDTP+Nll7EZacCyFX42t9aP+/QrbMG3zf
whxd8QgIar8hkwdAeHzRa6sfax4O1/WOaU2JJbMTnmgQaY7BtFwk1pq/N7E75qerzCEprxnzUbvG
fOUEgZ+dn5m6vSy39mHhk6lEo0TjHIb61rYRosQFOBpBjZDW65sGh8N4K4PGqD0yiA8iayc4akM6
TEB5REsYnEwEkVsGENt8yNsoiinwOheyGVj4t7GAdZje7aQb0sA+amZw9E4BkSw64l92/SHufygC
iagbUtLeprXEmHgAltFWKhgUrUliU9e+vldWsnwfUDdFHQy10P++UNWdxhkat/n66mn4rmv3Wr7u
+rRgNc/uxnmcqY9II+0JHMJB4hqnYC7FktaWMfdCg2MCzBjRCgYA378n6r3VjY075eB06BcELCTd
kco3a3TI5kkbHRUor0S+hwkOhl8uOnvMxCV8fwPtYdUEeutd+JkHpBHKmeOorXsf8IQKKGrC+tfr
y0cpxCHdY5N1jjyn8/ZcSp3wGIGJkb2bym9FnG8Tfac6e4zXSzlaA7VsCoWXQaxKnso7QAM/zNGh
lTqeQu1a3KOXxF2/9Obej/gFpe4hWOVIAsjZ4uscuDfWX02o7Cg/LORvm+5hyBKP7s+jmcWGBDI7
bnTVFGeN1Dv0RCvnAvu0oJD2pRkpSt0T9bUFp80V/PRdr4hrXbwn6SW1SFGMTquw2tWgKxjHFRI9
oNBZBy2CdOgrX67RQwO/AR5wwJqQW/yj4gMdU57dLN/y1z+7+jeN1XTmaCdI/l6jO5sCbEVXkF3K
Y56EohZKnOrmwJFS0/Yfzm1AOq1FETB+5RVEspUynFx1+JQonXOMg0KY8hIz7mMh3PPYvpxC2m4V
jj3FnHOW1utCWtf6jC/ot2iPgdPpEAkpEQBFNJfEthpb9fgh1VBDf1JEUTTm2UkB5+Cpf5xY3Jga
gSxua7KOwEGxIRJR6KhOVcj/KkTcAwpU6PeB3O+yz4jZHf3wTN0GDNA4F6HwlT3LfXKqFjNUvM4i
VaUTHf5nDQJe6vIvHX4imKhJJPZAWv0d52Je6se1qwc061yN2nA9c/5QZdpm1pHs7l/NyljRp5go
f5IyFuv6BN9WiERmhWNGgCvPZri2fIKDJaZc1fd5I9DUPGn5EaA09FQTkmRWmp0eEQaeSTbsMUtv
yqOtdZY8VMcRd6GSNeWQQ6CZDOmExvfU6OenGG0Y5Cd+wPsSA9B3Y1UTluhDUZyJwRjzj3jZ22qT
UVf8/jw6nZfswRAzErUa1TAaUL4rIvJBDO/RnSUS23sD6RBlloOSO7ot9L+P1Tkhg4ncpJaAMWkG
78CvuNVnEaft0rUe3Q0qM4gU1E28X1EcPklv1vxup1jG5Xa3WJdBRU1LnW+ajCs/HniaMrBJD2OH
jdJRLO/OTU73r0EdL49LKjMRIn9weogPPmM3+7ilINYofiNVfN6cJE3/yK6kUytzQV5gNGg5DQdS
jqFaufsKz9pw6LxUhz+vld35S9vFxmnw0o76nf8Nez3IuPe0GEj76bZ4ooYuByS0DHrHxoM/0eka
jt9NOTXOmsq8wlzvAEw2nBImA8OrvPQE1xgQ8jQm9U1Mt2zVCiRK4QAGzjBaz3WhdeMxNDgrzdaw
rs1+BgD3PqQZx98r4KWvylzlw3oEjO8mX4u2I8bhzO57Hd7wT9rOCkZjDyaKOhHYfJBHHa6LU9Rh
XkAl/t9vJkiYoAJZIL2n/Sp+cbkTfsb4PgT1TdPix5Bg0b56+9d31SQ+Zp5K9cJdLUnqRPM6KX08
eeQtKxizz+Xbny9DqP8OoSbveQP310ecLsRY41kx5fomDx/huwg0gvPliQ5F3rk14mMJvX+sJz+h
bXrmLllDZzQ/bsgwAMNlZ2WoikLVwgzH23q+AE3mAiaf2OIpqB0ExfqMFXRuGLIUUhvTutZ+UxLm
7zkZDbIwabhcXqBLTV1YrItWRz9b5g7RSawQTFOTdZNSxG/buNZGk4O7WEGOlnrbSswzyScN/m25
oEUAx9xre20bcJFuOnzZzlXLCceOVzD7F4yscRBdO4Y4bwd/IoEGYEeLKKAPAN+J92BOfGU3057Y
BZ7+W4nfwXx4qd52qHqe9ccFtIklWbBBq6xpTL5Q/EP4YtasWamENRt6XrB0TLFgugFwsNm4PB9P
+xtrlxa3r5lhcf5ahaHHUpi3UmC/FXA6XnbImq4MtUEDIU/qTIarSKvxN2voIM/pKZJ0LMGhz2K3
t4ox4Fj1k7+5NVf2SwipU1zjSviKvXBHRrQDy/o0bq20h7FrQCHOiTOUJFdWaHFdMVSoC9B+nEWR
VWnfq/bq3FrHnHlYz4vZoo1kxH0+WcR2TLnw4YYXhLHuunxxqCUja/QQZjNzLX09ldIFWiq+49OD
oWdo1fevBofexZ9ZDZhRhwsPgZsaZoOImR3jmQo8U2J7nOkgHrC8BrcFdLfFq//WeFmJJKd6t1o7
5HQZ9bVY/4wenzRxEx+C2FWBlc4R4jXpx8Ngritke1hhcw/Gl8B0l3P7/vMl7BQw4/Og4d64JS+q
MkMOF+dZu7W1JmZl/AEMxiEkxfKWKqpmbMdLO/XXWc8/+yxpfR3IxLUA2X+MixeoKScjTVGuye1x
dWkXPGyMrwgJ38JvbkY9UGAkuQEvkzFPVTAMHb277OLH8DIaB7rxf/iRUE/2T9mCwfRRWXuThQU3
M2ddB26pzcqtKkK7WJknV6JcSPK9nMAyrux3uwoOS023GwxG3DluAldDqXDSobUnEveiy5wigiHo
0lwAxtQJdFK6OJ9CkDF5GcvTaJ4oeID7BkHPzHjEWyZkK1jlhSYZYWqtFXx7uOSSxVZ8r0GX4M90
Vm1+JgYvXslOMQqTcgOKEBeuRJ4eQReQ81NKoQRHbuDB+zbhQ3cKQhB10z9oUASvFhXHHU/zuuU3
zwSIRehC7M3Vb4u/Nh/o9jGs17jB1NxUL+nhu8braf41BBkI4CFb85lR83H0+6VjuwL1NMn1HtXZ
ecQoiEwQrGGyJzYflKF8nVwEYdnuEwEZ0Q7LyLXcQEUfMS1eOK2yEapU5EXDFZKktAHp/MQIhWxa
2KL53jJ4XQzZn3vugCZUXTCryEFqNg2nT55j8KOjl8mA8sLr2vREcpIlPkQplv/Pv3HM+uSIeHOD
/i1tjtbqJ3RV8HI69UknmN7+5X4/kiZunIj+88EfO3c5hPeaxlKXmCxOfyB6RiHq2qa5nDzZFtg/
N7wBskpEGFhgY9GbZpx1qEdYWCyszazp2Kn2yAwh7Fxk+9fobMmBBUo5vJ1eEOlNyygPk18CIjO8
ZizMmrL4Pb4MQglVNVrojr2UKqeLB/EUkdtaxezMMqQjf13Rcw/so1dH7TNcW1GIe2hBkC3ZIcPO
3LqgjuOwL1qAYOmC+gS4RbidvR6egirM/TCDm1xSIUksLHhg+Hf9EofvAYTwPfF8qlJDq/p9OfGC
YaQqS+er/85fhtPjA/GC7tWJQJnrhszxCzrbCfvz5AxOhnkrdoEr46ml7b9/YclPi1hNcVzHSuvF
SsikD7jI+p+Vws8NV+cNZ9eUqPtHPfEJjFAdbKC5o+6LEwdblMMUpEGQT+kUQcFrHhf5hjZDuCT3
2oHl2NCmNBc4DyLUIHLpG1g4qYMvdZXK79aMqrJEOjDGcJ0p1LBCUnZBaO5fFFigCfuCpyGm82Hj
skuGQ6VryU8NQJ5/iCEskuClhg+GhFO9E7JFdnMaq6bSA82kggi4Irmvcfp208Bzd3vnb8HdyhiR
mDzjpnQ7EPf/jtFPF0jUM76IgYFfWxceezPI2oQCkMLPSv0a6wDjUZINYLmI5YqqlKLsNI3r4lCZ
VuDhhm5ReR8TNVWQMccnxsQG96ANWA7LcOvFqco7wBawrRH2Mx9NVmyny529VrZXh6QvWSAZ7cZa
Vv3xtrK55cCckG/XSgQ11u8QbmdVmiGsE8tMk6Mn5iOPSD9UySiTvfFiMkTkq++6TYiFEWmmcClb
+vIIGQHv6YGVWrqzuazXUigPk2+73a9wa2MrM6S6Wxq49q64RzHqMGcpt84n4CkDpGkf/9FhRtFk
gaiwBbNdvTSEw/x/elgTUzbXnMtn8ab3/AYRoVO3yF/zXJ8xioMBHPp5lYBA3J9SP3rlzWdIkxPz
nbFkqzlbKmECWGgIeqZGJruVV56CRZLq2Ry4vtkFrRYdmp5fpfs+rkUU9fOI5QGy2GdLFdewAOGm
nyA610LJwYv5vy5Uo8h6wWhsSHIHgSEYNUrngouUPwpjRnVBdlVQozyamLeP575jqCNP77sccp3Z
swyefc4kjbeIDMplLWgvbqeVWJiX6ZU3i6l0Tspii72nFK0hMeCkxxkCq6FJXu2TFlHeCEPHf3EO
3rpd8dlhtkOGgB08iQjdynLN9WEgrF56CcX4seSuYfCncjHgUS2jzXOsnuLIx1X9HPcJeCN2XGWj
/r2J1eciZH/h+7bqLNMCOWAFs0uPBgh7OPH93EyBVrf7kE7GKu0pKCSJxv2rs1gc/F2JXk72LG5J
vfFPMFFwaczzrxspOY3nCMndw7zL9eko9bGi2+EHrnNEHPC3vz3T2rex2oSaF500kQowYZ+8ypdt
VnFMq/zN7KRn5xBJwGz0ECLY+mSmzUGLPMCKk2IlkXrbkiNia7Vrb6XpG9AWTPyyiqTKKHMMCLh8
cr/aiUtQ2KVComiPFN6HX1ETiVuSwIn8+EpacLALrhi7g2q5+5tf1hfLsIo7hqWHUTuP9+QYJGG6
rp1b0sA/45cbpOHiKxo/x57NmPrYNK/IvT+CkXNja6HVH9u6cOGaIffczTnhvw9zcqcdKdk9UKGj
fHORkJAUT76BplB9y1IZCkm+izjBnHbt1fvKTw3sxEw5ebVqlTQvqNB2BQDPgSdpPr77kGhSjnwo
Fn3qjvFbaDR2ivzQ+E0iBWl1j5J5KKrRk2t8w0kCe2SN9gWYKCPaIeHmM2j6xqDkp8OuXB00ZRyO
loOfD7eG0ufhJ0O618bXSAXDInD/Ck+orGc6tazpVMV20+0uE454RxE1LnUBTnKuKO7iG+2yqA5L
pQJbndRXUiTwZi5Fuvh8s19micJ616Q9QI4RoDyMlQLpRRH545IUpI0mUnC3idg24t9/ZXoFJYGZ
qZHFa4grEGXDrGP33aPOMLSxUEhre3RSEHzKj7RBojhmS519mAG5faa6033AgmzaoFaiq0sRoTs3
phG79rR+i1n5pADFuRrdHx5jeYl1qVJ0v9yMGUDiMNJMNgcprDxWzpyjU5rT4G+vZrmDPuUyR0IW
JeFj45whLWtlG0UEiW9PYkAcqITqeKREWKc8molvLNkWoPJNPSyh42LSR8/4ysaDbeoA9USuwPE/
SzvZdWaYZHjvbhS7vXlYbR4obgw5SkPRUzgH375UwlRKb5OLvpkElQI3Iocq7N6Ei3+CTVY+H7YQ
CGQx3k5DK5GpzxC88ei4LZymfpg5mCOESFNNn9GNZQh4FqVZlVZcfYPl0m57lvQ/kGoZ7pYNWoqT
Q6ZzFHF80hANbvawWhICGuVJg4By25tdu96Zcqkv8HeAJx4fLCGC5Z6JDKpRTn+2TQdvx9iTnr+S
DlnGqj3J30wkJOEynvrp5pOLgOiCTUVcIWlO7RYKMXYRj5/ncuq9m7HPkOrgFCWkW5BwEvnToTV2
laSerpSpyjL4QmBsaTCIHayHt7uy4CSKDq2JNxCIIanFMQm6zwZKSdIqIZNV4xy4SoDGcslPKLAn
pgf2owEuZiQnFhWYe00Tw+CXyvKT4HZyyFx/A+QOFbuEk2I5eRCen2Y8pXwU8VjoyAAKDfQvMvYU
5n3yXVkI6nr4OQrnS4JfLGxz1eOhfW7fVy1BiS0l5FdhgX5hTTdm4YQd2aYeUvC7+Sepe3uYDdBD
fRGhgIOj/7TG8rFoxkkHiGgfM8WOsgqdziHyjU2fXORg2bvh20SHc8adI5XKdVChIPD6qWmmUccu
JyVKNfVLzLjIQdUA4IEljcEboV5hIc8V1g9lOm20CCBPFAI9gvlJA+K5ugxM5ubDkoYSxrtreaEU
tlTCAxPVBAYQctbrTeo3uXRLfMNP3+1ikD0TcE4NpZLFekC+sLRMf9kDmTwqaQt4B6MDS60zcs7G
gCfWvZFGn/P650g4vB651BDUGB73L7ztlTLp9AMFkTQdh7cvCxJP+RzabaFUOu7J3k1RK9NeG340
kOaCJAeq9QDcfmn1OqB+0cUUlrPJ5GM0/mJtj7xefwKG+iEwbIgE6NFmtXHWVNjqyNlhtRGANmKn
6uKMM+3RiSKov+ys+YGEMKEVo2Sg6lNOL6HatMUZcuirp60mI0+lNuaI599GEhgVSnR56F1yf7IY
f+IN9uQvD8jvNEM1k9uTnGSAivZNZPF9GW16/C9NTNrMrwi6XubS5nzG5WnqjBJJH76FKU7BJdHU
/e39K7jO1ww3rvMFrg5bmHzE6TTJBmR9FTL4rWepB1REwaw3SR0tDP0z8CxrwZgPHS8YvT34i66+
mHuSNEjvkixQiW2gNBEH1kAxvhWRoWfzQPXFXwNsC4tS0lTFN4iCifAUkc/FB6eFEQlV968dpSoN
gxCaZ7/S+IAs+tTlFzJg46PVEhtDqhWoJC6Ph+NaOKpi63xaMGUYoSaq8d0H4p2QJR1aBqTjOtJ2
gmN4kFNSd3h5XPbbT1dPv1zl8pShpmUQ0WlsD++2LG3nqXXb5Ups7+P7cG7w3edBSHB+rDUgjHNK
Yb4nA0Hdcp8srEBzumoH84ZRdKFpzDkj0qZ8FoTdvBvLd+P9OtVJNKUVHl9cIRrHwl3EEspl2XYe
ddCWRHtphk9SXGeQAO1twUNnl+uu5su9TQ3KPGfuPvc/5A9GbPeR5P7M6Ty4PYQ2Y97G3k/nrGaS
JH85Ei82WeM1gDQC5Nr4Lc1vLhYcn9cPvHEYRE1DKa1kHkrFfhxIKI8sI4xNSU20l8+krQEkvdQr
eGmYjHUtKzXSwiYAlFEz6CjJzBDzxsSFUW+8Pxdqe0kz2mKZemox3mCQgmObFbPbLCN073IQ6VX9
U/SLtQ0+gqyNso7wjLRm7G0rNSYeArO1Zkjm69UaXH+32mZOM4U9HY5DtWezd0l+bKnylIU2jAyz
jbrlh9XyZizNG8k4lLas81a9iibXlryHoRvmL0ydsqCG1jPvLAR/6xhz4PNBpEdanL8C6VjTYjXo
NbwU0byVoU6c6lNN1QWGpKrL22nVq5oF26agG4RTcuDNTSTZ9akuSCIkJQo5HgOwE/EdPDx3oR7Q
nLrO0A8jymvwInj0PqTdsuo0pAm7xDSp8BqklifTBYS4ceNr5+7wZ7Byp/pIZO4Y86kjjNgmURuY
esjDA50cI6CJ5cSGmErCeqrRw/LygTW6VeBB3rOlaYMx1WNQrd4gHV9ebgxuP4hC1mNRT4ZQEnr8
w6yGQZ61o6ZOdN4Lpekb6p4VmWegDlw6r7PZDzw+bK148qzzPi5qohxw7BxA0Lb+Y3owLVod7SwQ
xRSF/0/wLiRNu1KObvxes19aA4eKwvVX7u67wmOTx0OS1WOlFy16oMq0VFSaJXZe7lpWuMHdXUtJ
oW6AmqzuI+8BHIj7bvgYNfqOxC0ZJWCFJPo3wknPizoaVLz81XzNb8RDVdhx55S6qRWRIxAKbj5n
DkBneeay7QZTTP95hMXA4vsgZokWh1EB6YrBDpkNg9Jhz1SixrCl59VAjd+n/DPPII2OM1EOTvO3
TqQK19R5hJKY4FLVNts8kwyh9XqFWgI0Xac2RCOuIpignLv4x/CrS2qyjKG7cg3PqEAYwUTXj0FI
6GI6tgexpQ/C4DeCPKVmhBNKKL/O7vG7skEDGs9RBODEHidwvVDztF65JsQTZmA+51iA71gX0t36
fBUTd57jhlMyhs4jRURPvJM72WcOfg+KbqgeDgjnPobfoXAc0mFemc9i2R0QI3Lp20FHoGaCxGG4
ikSRrqcby/AmMzqHXpgwoxevAe81Dj95a8F/CrYPLB3UcezOzt6fPZikcagRIc0D4r9H+ALFhTD3
JpAjIcizO6KX/EgdUmu4HQmTMPdC4jUycuPhcenl7JMVDhy3qXse6QgXOHscxwLZj5FXk0pc83pS
qLRF8jFs4DlSYgxG1B9+aJXAPdk6rVvOjpCMZDGRisvk8HQV0oCmgrgQ2Jg8aCvy3RBNPe7pgwYc
/Yye8ZsBm7NQfRJgbZkaAyFn8TJcyJsnQOKm9dD1bPzcHIv2pRG1CQx/Xm/qatg0hegLMMyW7fld
flH+t/9I3RVKg7CXxcjquO0V15exBXyNiQkkXkjoXzx7QAIOkZVl6+U+Ifk21Jq5Prj0zOmmA46/
E97Eor2s4HN1ep0HrK/yruDrFiyV/tGrUwVTuExgAo5puZJEOI4MCNX6sm7WPcc90l8CSA6tGZMt
kLWoFYGugyRSU3Fv1A9XiUZYhmIUP6IAE2YZKri0N+jX9vBjkQ+zC9QKQ3CgXDscGooDFe8RAicv
MeKBt6SvSdjLo4dOmix7mrfZxWeUSvTEb3k7R0H9hl7fXGN98wUub/9AsQcyRNtWrag7U2UsY/c/
v3YFenyzk55bODzXwcahrfM9ECs0u+E8bkjbBEahSlG80WqYJmInMDOvkMSnIK9RaF89TMq4eMqq
8ImqryWdvs6sTDKPZsI4Zexw2Ub6zppBR+rozquFspm76elNgxhbpB/W/NFUOvlNAVGfVFn2pZp+
U1DSZHYdRxEsq5NGan6A+aEXzIbMFfmL9fNsYIPE+vhu5SUQCv+++p6qLkDZYa4I0X+M3wotcqwD
Wq6DsQfYvFGZMyOfhJbxOT+Xt3tf2V2/t6lURWZviNIui+iWYK1G62Y56lUyoFhhSJwCEXmHubLk
cC04ao+nFyQcmnsuLyluM/ptMWYsKRyoip0n730I/8WEsVQ93Z+8u5or7fH7fVz4lFx1JHl8r+H2
hs42ge7Zwjfdq9ablGV4RRlsEYcyauhtRP9an6Ngw5DBlQg1aWE4zsCsPmKf05m7QRP5KWrq5QX+
coEVmUESKO0D8ruQUK6x/MmS4nnnYFiX6dqEyTUv7sY1wTiTqAuatLkyl/LVCsLdrwXlsXOzvKcs
+y2fr16JCiv8IKM5my1Rnfycxm4QHq4j8/0EmkuBuUNvjO7MlrnNOtoolL5h8TsFk0vVI9zMdekK
G+g7kAX6PhKdJSKu8NOQCqkgrfrSzquFsHfhjV9p83jcydiVLvINXcmPSokO8yRhpTkkb+g34l46
OcMDBwVFvaMcsOYNCp1AvTEfiVkYi3GZjwsKutlCWecOnOE+op0w5OpHLt8JpgJCZXWItTGbcB00
unJYp/UzOpH0BaNY5P6vGJxEf/QUkeRDaNQpXBVoOgqNKdW56+8SiAMcQEZhcre2Xxkx1IiDFNmM
ZSCYw5FYzmApRXJBUL3auSrPcFe8OD+XUuQFfMcK18SJM5vbpsV0jV0tUtyvGYh9VblX6oem4JqU
T3AJY4gUcmsD8Jvu80/0mhvFPDoeWM6m3ZO5Zmoubd6W1jH7Y8/tMiaiDZFTzSxwMtQKBs/Pzs/4
5dh1Q4x7sX9Idf2lTGpiPI2+zQ+WyeVTqhfGJ6+u3DglO+JG8iU8lkQIvMbMZc0W+GAeEF55eVPx
DFss5WaBfqq86cDTHj7FKzJsxL+LQL2pYHEBTyq9L5wNo+RHs/ElmCfUsCMKUIdAF06q5H4s5QMJ
8RM+8UAmpqJn3/oiZrE0Sh4vX7K/Sk6z+ZlBs/MRl7V3LC6GzCtFbz8lLewFTO4WUtZlKdLzqsFp
pPwHwseW5F5Ag+lrRQnLjblqu+50tGOL6yFY24aJ+ezKgTp6rB45x9i6ujZ5BD5BF1zxscS3ENKH
IoSYTG/9pjCieoQj0tu6Ek4LIyTCHRXQQLOG1K0S2jrtSa3HT36g9HTRFDwWhQxYVivJnQtxkoWa
Tfs5Yn3/wQldnuPhBgufvbKDTPQtmcfKqv4SYyBEcU2AiNGie7mh9ZLtfE01aEstuL4wUQ+shtyE
6YZwn5E4HX6MwLNWiMD9kALL0+gzcPvUJtvA0ngbeeLG/GlDIzVTnyl30G7D/OMuSv3Nb/6cvaAs
JqHsDmlVtSNcJEU8SdjLzMDlq/A8392lea+KlcuCPiupGbkASmVtZrE25pVksun6vfhyX+S/5qXw
+hZ437FeyqPt7/QzYVZ0P0JGEJ8kRZ8xMzQm5SMdHv8pnhFLhE7gbmollpoYPC3Nj4loSHGpVVp3
qtyXxI8n2J1hI4ZmI1yGDTH0c3s2gvMSCrKwgRGRqCfFtI4J3xg+h50fos19f8IRmIT07g14UfhO
1G1la2IjNdblRiO6DQ/gOaNVE0gtSM5KAuUt2281+BAaWGWnlWSyNLpT8TzjGsjh23fblzao426K
mwlqQw4MF2xg/WKpNwesfHT5vhGGy50Mp/qR+6hwGPbf0BWjV3CmLqVyd5XLdz8X646bUmbd7ZIX
xCGiCMbmFKSKhrJc6tH6crF007cHkvTYI1r5LPppLNFMViPaeCbJPK5SSkDcjnQsiBBKT2Jc2f+l
SJcqKHB3U1s6U48Cr3NEbxEXHwk+qTctSLkHdKOUQ74lqX9BQWp0d06xfmFtK7AFJK44fFU7tQdF
sjTQbg2kjvs8zf+1URK0yWRsH7s8GI5icaF6ZnASlQiuZQKTshl/ASCdTPgzKKLawDlLCb8GVtJo
WkQdLcTMD5tp5edj8ebVIC/AQ4fFgf+MSzxXWXRTEtm1fJfBpCIbjk2j23UnvuxRSGK8qs36fBuc
9xeLA5UOwWCaDEMAwBD+yme5DlEoOCeOAOjkFSMC/ZAVZiWproMtkbuOpD6DTZ9BYb5olcXF7FyV
ktXOmT8rDYNEYmXLtzmBENk/k1ASGcB5SqMPr5xX9Rjbo22dEpmqhJh7m4aKd4y/U6QZRz9aH5dS
MDYtAlK9U8HQUgw6h8ETnhPSBSHo+GMok6nqzqPwHeTMOfvQ2lST1TE6Y37+XR1+1sLuEHpfAGjq
SuYA51ChGgPCX5hH4k1CiROsI+MbrGK2ZKV1/G5okj5FWT4b+53OAzHDbg4Zb5goniHH+CJBmnRQ
l2GUaRSYZ4vmpfd1WKJylheYXyVRLVSI9jt1kd/dQ6WbNV8LLquP5ZmYHjcj9opVnXZbiGCb6dpD
zchO2kYPfFIcNicJ6UopJ7tcIY0jDEn7J7IgREbr2l70R6nUgsLZlLfmo1MVTegbliAmoBAM19Sw
8x7ltj7uRM8q/tycMNHKk4nhb5BWAO27+sLo7zhMCPxbbSq32vMqRW+JNGTv/Y0UiprihTdZ1b5M
D+RTSExH1SsRxPrbdEajrQ3Ms9Tgl5ReU5QVo9jIsqFq8II7cnD/OWfS/I/ZIv+XVXEfDUXaprap
LI3NOFQPEdTpGCGOLAqHrNOlS3/GlP6mcuhwfA1CmSOHTiUMb8m/Hd2amaAhnbrTsHK3LVfIj1Ng
rdQ2ThWC8JwVCNIggcPzKud8JJWUoZJB0fP4kFumHPlLGOmSAO5jg7fMhVI1ExsjBIYSGPOhpOK6
Hc7bhpwQLtu7P1sWFvJIPUFRaZbmuPtwni1Fg7/6LqxYIJWNcfde1t58Nb9K9RbOH0zgGVXONlF8
F83xrej0YZq1oVAyTPwBkC5gLIZY4iCEMwp/P/awBf7zYk2AUepPMFN2SYKCVMUywHrugcDU4PSF
iBbEHJsl4I3SZEkyZxnm358lseG10oWCaAJVvSh8q+JpK2OBsdA4+Z3pwh6ufPjtG+qRjIhUp8X0
bX5pgE/DLfjoXlgpfR7kbF7ZlLcY2wokiOXtnTL9240qDYomyRHJQpSrvhmlosBz6+XxTLJZpTLv
vmszVUCB/3om9/uiIDv07K7wxkZOBjGwwA7XRgNyM+sd60ps014lumoZvYMnUPKQfMaxjnvzeHj+
LvNB3kBQjvoOO/5sop0mj2BB6gUPkPmOCYpUkCoqYCyl/qkYgVAPFgOCsO99smZL45Bn0XYkAGYf
lW2Wnqq/CgdVjrYraAgiYFRr9PbfWCWXjgmHG8eT5ZdwYFgsb7pMNEf3mX+LlkOrsDKJItEFktcK
Bs+BU5ZRQvNVkv4ltTVnsCN7bAmIZGJj05dbV1jx1MzQ5ZsIsrV4nfZAxXHzT3iyYy3ZCSDw7LTc
xWcaTT966FpmoVppHtvcEKN7tyL1Z3FYGqC49KOL17aXgx8NkY5Su+bSnnGygRRmZW/2AyrTc+Zj
mef01mm1Lun44r7YvxpdIkgKgU2EO7lNahnJKvr7dae73azFC1FQh9iWFAqfE6RVblQqTSoTl5Ja
88/Xx05MVNG6zBWTGexFIsoEHy3n01R5HDNxoajzW77GW+DiOn67M8Grr1s/iXiRQqhnZ3F7zEJ3
xDo9mLckkIWaZ4kpcVEUOp3hvdZiZifY/aZLGbhMv38npJsESx85MxtomD8xXyM80RmmyzDhoQds
vYxgj25cV6+ZkudSsXRZC3Mp+V3Qzq3B3cIfKvFl62MEUZpUI5paFMK1nkS3XJsz9F189UZ1Iu9v
oGd8+RVvN5iYcmJ0uwKQunZQ0aaevfPuRrGTtfBJ5kFtMp4D2DfMcVx5SVRkbAdVCYTdExssOq1i
FYsO3vWYrzf3Dax7cYEvOICjoroCTpxLNnn9Ndw5SWt2ETAVBFK6YdEPz5oFAj7LrhM/tU/P9A35
anIUn7UHnUfdj5CpiYLQC6fuCIdKzh3pyAtlB6esq0TVzw0P3ufo/DMBO6wt/rgNRl5O/xEQ78CP
DYkUYWk438XBAzJtoEmNdBpaaBCLYRm7k6MJ0hY4UzcxmvAa5Rgd6gJj85OjAtQEz1OHpOsKRSkw
Tg3y0yzy8kpkRh6KSGY27acI/K0yLbYHJRBzkwEie1ASFJ6cxEiM8CC+g46Zv/leRg3kZ4aV6InP
N400j3oKHOnpjfz7uytoCKuC7XoUJtInmIrzRGean7tdIx6tioLg/t1yuRYbd8J2oKT/KLuw+Xai
Mp6Vgq5xVQZcsB2F5Q4MH4tAXofdOWkx7i7FmWoM/IRvzw05oNgOLwYSqUESKp3oee5ttpPBJbnG
Vr/YDD2m2WMWGPW9Iq1ramzIZkX+3Yuzwt32N/ZxTcEzVU3y28TkqgbzJFPI07Kbrdl87ALH6wkc
BPEUGjwLKzRhNsRa5G5taXlS3u+FZ8YIXBEcZKNdJ/Dlvqj39RW4j42WieSr9qJ4KplNIX7xzfKy
B0xOOGPuAgNbIqL4zvKAn6U6hvc7IEkNCDGUvt7e8Q//QwiLvvWBGFWjGq48qVFWh/bCvobudus/
OHWaZlUcATjBp5LZp5PeQL6DjS4MtabtSiRT8vEaFFPvUVoDqPQwl5zmkE9WlxFCNQu8KAQCUXWf
J8oYCyV/k3CZ0mgT7bJIU8Ys5D4zL/5RtB+89HSpChOPhhuR5Vh+ct/X5g0fSEg0nHGz8rWHop4p
nu0K/oZsOOiEUmdF00fmCam+GRC5mP4Z+CsSuEhaTCo6Bh4AiYaFRRZ1UiQQu22/kqIft/GOGAYl
tYYlZC2glN0wRu6o4r85sLUebHVn2UnU667sHZMDq+vXPslCJNILwaRcUQkOScUeft1PR8oq13GO
SnUBclQOgs8JBAmEw/BA4p9zXEnBsMRcN0Udbl3DnrHoL2fEzb9EcPp4WnKHpjPFBcy3SVasZQla
R1Cau/5UTWUO0mzPUzkG4ym9Pk5qyyZD5d6nkPAQUNGVUPdv0Z0i4ixPJkpxhbVTM4sW/UYRkvKe
73LgyLa9oVIpYvUiBLvsKwNJLIhUyH+BgEK4q4jYyoeCicL1QGOwkfA/WKOa+YPxpb/mftKshTOS
ZXoYHtSl2q6O7kXYoC8asbU/u6S9FOuRL+v0WGvqssZQbD6ghxQDdwjNQ3jZoNN4q9YCMWtvla/N
1GQh6LXQn+B4WIAcmZugnB+f+KwPu0VLcPPp2z8PSYimAd00FXccwAKogpACyC/p1rciN66QNwgB
SSOhse1gs3AhKF5SE3xtS2TWY6qerAmTcNMjrcSGQ2T/Fb9e28TiMSlE/Haih25eHV0o/z40eUVF
fxI0l7aND6sL9vUGJqRi53s83i9w4SRzsMsPrbAW6TIn3krsSzy0PXk3mZp6RtTR9D0gB/2bK+Ck
ZiRQrDxunO96JtkLUfKIDJevxEYZsALUokDVkYxYIib8dlFypYNhoh6aOA7FlWjPFPHpsTV5rZX+
WkNSbs4Al5eA8LgpSrAIxhJZYZ7Ir4vV1e81h3WeyDET7RMhOrptIdxB/K7SOgCpJXmFUJH3AQvK
U1cjCThz3WLhLKsMOdi5OCzk5y4ahdA+U9xYCDyphn3LOnFdwEUIA5y/s/5+Mhk3toWm29vyIiyr
MvRmC/6tsJOz/fijqBeMTs9dSeXzIbXAyKbuHx6ik0TtkS1V/g1LI/iIpvMB6pHUXbaIbIXd6rwZ
1xkvbSfkZAYjyGaKmYY83jYBGKZi2MwGtUTV/RaTL3U1XPjE+8wMS9eREvhqEOTZsV6NQUJyv84S
Fva6NXRHjB7UwZXb0KVmuP/iI0iBo/KYBDTx5O5pmrMyasQw2l4cV68px3BfO13UryP48/oAodDi
ejPkYGQlsgG7p2m9r0tp9O8UvQ/jpK0Y1xQ4atbV3/VonjTDpnk7iF/zPoRZrJzCMAgRWPGJdS2R
+/PeaYGDm6DyNMuGtSROPxqvFNjmochUBLZXceeHIaUn6cPA08yxvZ5kAV9XUionRyNsWcw9QLqO
usHZFNAVKri0byloT+Vi7ApOVhEtDbWw8SrQvXifpz5lI7dx7KaxF5L8cb6IygaWv1B/byWyvNzy
41kbGansku3pXlOQtrf8PDm2TR3wRxKJcqdrmXLSKibuUs4z2nWzwLEhJbPnVMVuoKX4E2qzXLuO
v/Nfjl1nt2QZcdPzgpeneMVyJCYqFMPYvbfPbZykR59H1uNRoT/QjcgQYNUSqSaJG3rGuehmHZrK
JbdCVTuTUPFc0PsJ1f43t5oAZZ8djeFT0QnvaKenKkMl2w21i6C8iOVc7lVYvXQgrsZmM6E3YLrt
AUOURS9OfVw64mb+8vF3ei5btXdBU6hAmPnoEORPjVk5Ca3/KImtUtXU2KdslQ02U5eoCWXlPT9t
+zyjh6KWL7xdUD4fOdLKDbcqBSdDycCKgPiqBJ/zd0Ksb8vlK6jyIcWrXBxJ00Rjb0NrCq3iDf+6
yxFGa20+fTM24vZ3dIbZxyMp8AOW9FtUjqSGaMPNEeopOw0eITAoFiHnPSRyxD9lDtgh+Er2kgR1
eqYs8Mcp0Cr44lTdSEmuiYCuGQr7/214jcOynGlChs10DWaC6gJK0cJLLmdduS2it26Ri+bJ5Owf
qIAmoRpdorEq1obqRGGlwdu7ifltS3GRAuiZs0NZo2kjyi8Xd6TMe2wI3q7MNsmsVcW1hVq2J2Fc
Tsr9Lvn4Y6miVoTSPZjc0UYMUv2PCdmKtedlLiVfzsrqX3fj6P/IBmz03C1f4NDd6bRiXAnrtv9K
eATfSkfR3ZnxaB8zgUVID66bLalMOegZ0XiG6vLF6wVXCdmt24VxptBNhQ6XalrMKPQ7ngM0WZZY
ENV8OeoDQp2yHUyyrQOpSAZUkxVqGmoIqbOsun5lnnpk+uKEhMaq2ZgT6gs5bV/b73mmCfQOMz5O
HGE06oc+kXsRrgH1XpYmqRzLXvTVtL/3tf3CBtLFJff+hUTdLMjBkabnJEJuFmkCoXm960A6+khz
+ooq2i850+khgyHIS1UihwAJKNSMPdRxNI6z486czaYe840k8y9c6+5EegawY+3QGclY8SCIiWji
EBMmnw4sgwy58jbLT7mUA6R2SOr2Pqt8sntFYNJujrE55+EGKXweT6ZceQpKlvC5dUHBT43RT7ii
UAWxwvxlSAs4u0tj4JUQP0fkQ7bh8OFqeb4ShZBs1yLJaozO7SvfbQ/MYFJczVgJU9jiD/61+/UG
fsVEPRApxi/y38wubGtNuZUKPetjek3eYqc7kqlr2Db7iv58VzRdNh948h5OwHvfVebBh7/I9iVn
4r43WBsk1dQJwHTAiYe+cytuypqZpH1XS8i60rsHDgeqG//5Ckcgtii+99kaZDCrrneSCb/pXkPL
RtVn9hQWlxjQWzlcivYLZx+jQVVTS0smDiv7BdxQ78w5FEA0n0UOsOnx4efq/5CcfwdK7m/grDFM
j9pYO+io5Q8ZBoPTxpB0kHW6U0b9yvzOOHqHEiQZs2JHyNUMrTFlz1DRfDGt967mUvF8aD+zGPEG
HizLb0VglfAqtdfUB4jWyRFXdHILpeJjd2eZix5BFf6PN/seRDF/HPo93WwEiN+k4tpyrPuOKzhk
Ay6izROjvB7r6m06XRCzVtVLuOauA4/Z8HwIgkDY+IJtofp9aptDYMmFlOYx9xMkYLjyxkXTuYSo
4wZi8ntzfJEwlxDzP+y6c4emBbzOXes9yyfH/FKATn6yFqTtf5h8BSOdpmTRssBDkZ/dFyEL0HBQ
oMTdNYi7BPE8/1yiL/Bq3oUfPVSWmK5IKykbRZ+6X5kfmBcv0TKqqb7qDnj8sQgqIN5PXFTOwtfk
OdFI4vNV1GH5MEo0nmMeE2izlGbVTNfhchWuUbvF2XZnS1/oMDoizexLOdU+ildJUq7CscuFMhc4
xuE4MmQiq25e0a2Hxbn9fAKPvzyEAMZPOIMagl731EAc158ayk9aT/ntEgFqyYvOZY8KycPJUn7M
luhGn6RjpwdWTGFCBcrS199TrxRoyNv/jnFgtQ0yS3lCqq2f7Z5xrQocNNgKahxx3WrSXFHWxq7c
688pY/UnuvzbjCAWBPatyHXIm2589tKuQCdYMcUimxQdBdDG/aMx6uZmLMgOFpRUlG/Oq+CXJfPM
SZMEKvodu/L8HxKK9oIwsMogBgqKUM2Gk6h1gzxbzjn14lchxgra9nUwA3Qn61ren35dTU+4ixJ7
G8n9zuLC+IiK7lFCPMUPIwRcavEFAwPY6LD52OFpkTcOC8SAAOBKAI/G54izU/dShhdxBJbqzm+s
yB91fBvMVOV34ZhGZpPwUsxb4Phg9KgyfRuYhKLxcCSj/9qCGavUw7jHE0oiE+dQxfim2KSavTwW
ie1YIsmW4eYw5uVlwI/xfudVQ7G3eqGPNpmYKraNebDVBqsa9SK0ReVB+n2BZugBRS+zPOACCKkz
ZjOaf8jKRzmHQF262bVVsLsXyi5aINiSHb22Vx2kaQoA7ZIinkqn+H4ADesq3a20JE/EBoEW9CiW
oe8oIYYzXMXGk8mSt0zzmK5vqZzqP+FD0pW3odZkzpkMtQGGuIOxN42IiP7eYlPf/rV6/BwD2vrO
kPImC4RUBk7x9AH/6hXMuSm1TmFsdambRdTWk0duhecppimbRF5ipiHEbAdE6s/lDyVkaA0aBZnF
kIHYTasJ6GRSC9gx8Nf5maIqFprhARnXTbGkaKKbBtJM5EttTMR2qVjRsgedhbxNjUvF8T2K/uio
qA2oLCU65KEhoWrfIhgTZzX1cX1uLQsFRYVGAjf0becV8eMmF+4Xw/yXbp84PDZQvYzXiGuOGf70
2EnOvIuwbiSB71nvYUNnBwTxuNZHbmO5mOcK3ZsXhie9BTVXVCbtgsST/R4sHHiymGI0cjB8jn9N
6XdNtv3TEcVNNy0YCSDg4+kyAWXzJwA44aZaZrN6TuuO+yFlkue889FLRkU/9/3yM3ORby3+ZtRR
O/m+FdNCHqgCRm3hIrnk9hauccbdeHZCvxRJM0Yl+7dl+PwdSw1RASVmHFY0s5QNMtjoMOEwlMvk
AYDf6sRbo2hbj7zRZKwLqQ+OzIISqAPOhun5Qjk6S5FyDBnPs8qrs0QqTFHs+/mu94OcidswNk1P
YdqkhoSCoYtmDh88zh6eCoe5Om13JITcYOilUEQZV2ceIKjrT8Te3UxWftfgUNzdkhhL4b2XQB0r
pka7t1S0BUjU4MSej3IACCGH4Qmu7VYlrHO+jYm+ciEuKrHrA+Lk2bwysmLstvMt8d5GVBG/xuuT
5JlBaAZICpWJ8DGt82TvNxpcp1H7dYAga8r8pUgoe3z5v1MaBZW5+hDppCS/Fge5zANQnL6DMKGi
gGYaIsS49UKkv0+4IP6Y3QYddwhKdIjKuUrGEDaG0of35bdc68xKei76ROF8VV1gG2coV65YqzJU
atSNY0ZgvFxrTVWWjqkONefri1wWnEuO81DNWmI++AoISFrUB/klv9cNLDzIvOz16CylaJMc3lhf
O/Ts8xSZM8DbAPBhSty0bEN24HEVPc5uTmclFlKGw5b3yOcz8DZIUXXz6sND53HyqFVtJCVNUkpN
47ResCa99VV9v29Aalga2AzcBRhgJkXR3+qiKTYTYu9ZzMe/vero4/3Ku0NBcwHIvjVC9AvpNOKe
Md7MlmvDPjfJsSByvDTlsLB4Qtq1OMyMaL8HCUkNNL8BX/i2fHbAWSROigPaZIlwQOMMyNH4YgIM
c9lGLtuzrOQ56mNpL6WPeFvcQWeoTA9kgUGZXZlvRtFwS9Sy9yrEVoauPgMbrrmiCItlSQzwY0Xk
TqcSDKfgGrVUQqTb85Eyrsoxak9ChsTb6SrKnpGOTH06/xisV5ZsRhw8scEmb9/mQXjLvAtB3pJs
5k6QM2qjZj+jNdQuKHKBRl8CW9l0VnddeX/kcdU25rbxbOm772pnKs3MeNY8e47UTZ2FcQWamDV/
Biaou8txyxd8wfkubKtJkL59dgk7v0A3LNBp6m/SoHNRSacvnC50x7kM+uZv0pEMNEQAzsn0z5aL
9ySLV9DMbW/tDtFpnkoyWyagsRl1NU0injOkKwHCO6xSzQheanocs3tijOWigr2QCOcxyMpWVQ5C
0Xg581ogl5otxl5Mgn6VWZairF4XqS9IJwvZQzBbdtrm/DRUuZtjE+BAj+aELW1BDyguWSeb3UeI
oH55QxbAkF5NDwx3y9Gc4dMFXqUzvWKFLoxgNNo6Oiu/dxUviE/OcEBeoQ9hDOpRqSFulks9oYfe
d4RVlt/dlqLGWFqYRvrxS/cra3+whLZW11tukQQxLt8aLdcDbA0IzOtYcdNY9FPopz3DGwr+UamT
ZwFj1Noj5tN8SA0E5owstJ7IV/10DFZ1CzTLfIBcMPjPNdAJrHU+Bzv2qE/B/6GPnJO7/nm5ZV95
/aJmybVB5IKEo7viE8/zO3FMP/DQ9orwS8mVJr2pVCUNMuxSnaQEg+gFLRIWSLBlNzB8pYakn1r4
r8CGnrRMOR+kC4phcVKnm01RvFN1p9wonb4hkK76eaVutSPKNNJMllpIvAdTXM76ZSD/XTagJpbn
PHO4NUCC7qf5yAt7k6uyi3C8R/lKT8vKaA2xbnxPkCFHD7FRB/fDPIlljFlgb8a2joc2O7iA1Kba
lpIAbj0l55OHvflyCrdbj3UBd3tBJQT7vwII9NYGCgAKzgjUzkU/WBJBdeIPtVufRLD9TBeWMs0b
OoeQZggg10RJ9liU+/k3p7KmAi05F6RfDr4tgd0lWkk5W7CbEV+RKzLjv0GCCnclax24CoVuqOoJ
27CWfSzoG1ytsvU1Hpo+pm6IxpeFCH2zW17mcjXM8rRsXHfSPeFEuazQI5nfpWXE2L0eBvBInfJE
izXx+66MqSWrQO9CkEwnHv1iG2+VmnUof8YmTXdtiqfsaC3TJhJZzq/iJ0LKE/QvLc76NbtL43mc
Z9AfXn/jqClSF4YstcF5hdLp6REmedhlW48NkMbAPuJDEojTsxDSJZojQzgsqAvBTkbydgrqrCj9
aNPKHTX1Rf0NwkZbEpntnsQA9lMGraAI/U6/HgWgki+85DTrj1KeEbjxJK5tS1VzfsC5Xlei1QWE
mtUetv7cWRbrq56LK6XDDHihTmwP2Tbl87islUpmqhNg3Q3/UfQHmISqYfTKEkxsAhCtdrULbCGk
xtQ+Au79yOoD/T+xeRA1igo/rDGbkPg3bvJnLC9xGMzr+y45sfebH5lvPPVK/o4IH/U1bxxVyOFW
1X/gJBRTtZKk+QoQ9yDQVQ5qX2efpE4ankc0JwVB5vay6MpuoETacJ2p9ZS6bd5pGMaZ6X+Lr4/Y
h4DoNQMIJQ4AySw0SlKpquuhp7hAPtSBFlIrmTr7JZwG/NhsejDLy9x1yYT+aY3YvxVYpvYJggKu
l1WyiKL4fHBZ4MR2R3LFw8IRggjjPvzJVPz/4mYehCvO5vJLRxcdITG5X5wnnfqSvGwGRnABLGPq
9Ju8Lj1pRPzSmuniQMiHjFzoDKy9abVFxjEYls/cxt4d/CnHM7lRFkbdxwqANsa1Is39DPFabuyn
yppQXnvOy9RNP7OP4AFPNZmdgEjKjw95lXK1xgWx3L5ZVpPk+9RM6q0Vx7OFT3Jb2cpAC8BpALAZ
h9EAjpg1fzepE0CswzxrMtQkoDrTrpvxN5JE49SsHkQ5b39lVy7WLnftlAV0rUvs74fuZ+mUnyje
fz+zrAj6IfNl2se14fdMdCGlzRTHt8LHvBr4J5LiPUtshlW1THR51wXFmXhR84y5Asei69WYnat2
eKuOscreYF/uw5bP+BK2lnT4ci0tbrrqZ7fEN6XLvmkG0hJAE0GmWrpRVRhKBnFON8+rR+PzxAju
yuHMXPkGVfaKOYMoNAEP3ReXcn5tfu7chE6WsP5rsYPBxkIcHAo/ebOgsfc+rfEP6oLYv7dEbIez
SqurM0e+NI5U4DU66j0xZbxMdrZB/6fJ6SikRyg7obl4+NoOSl9dZIzlgYHdVpoywUq2wJoses0q
7MVkb4Wb0LYA9kSpennQdfcfUHNH3GjzKChaTVYCJdKYwntzFIvU3fusEd8QIynvPYCyiubeEgsu
b7rwXyevPftj3ACurOAao6ZO5Gq3EV8joJLVdb7JaPM3xYBfMU10WbinwXaarKacXhhE5D45Lwhw
6SR27DWWT4z4f+nl4fUn133iOTc1/s0otMk6pxpUuGuWldmFeXwWeJlF6MMGEIdAM34BhZjSIr/R
3op8crOCSZFxbL0dtcybSeFBru9WxEZWYuLFp44Q7677ZQiqDC6t7Hs1iX1+4Iegycnjhx8/COi1
H/q5MiYRKKkG6T7DrI0AvssDA1QsqbdtxoWFIZQfi49yCKDkXPMgUKiAR6+fsjmVrqPEJ1ARFAns
52m1XF7d4Uo5ctVfdvcKbzNUh01r4BUYc71v6mduYaApa5ldsM85DGSJ/UZwt7BR5kk5o9Y+5Cs+
UGpfwsUXR/PiIn0RT1NzCGuI/UNpau0N/Cg0ozGL6PP4/FPZqAduPZS7MRR9+J8QXAdC/GD+L2Tp
ULdqxfB5sXevIaXKffozoIlWMcXXMHDiL1Rh5728PeRhGYEkh23ztz5CQO82q/GuhrIToDHinNcj
HVqLPFQv1M3/LBJUotHrOTEJWuF6DtlTtoXO4+MJTOZljWrJeVYMJ3j6QKqlQgoNUavVJ4eN8WFk
GD1NDoCJ2Mh5v6HxEGuzjuSEwtGfZyosmNUjObG9hIIASGQ9V+BdyK3hPT6prwGB4Kmn7v0sZmv6
naFrdSJygdIb0ZKLlVDdlgjmZjk6AXmVvOS0ko3ujW9IpeGomdI/YmiKKHQ8q3PVrBcUVTH2alpR
ANzoZcEo40OuwsfcfUHUjQcncjFIMaSBw32UPd3u6BF+IN9pfg7LLQvDTQVdE1BXXGT3a2/13dtu
07d5RQgTYti7xxUg8cLDPvebHp2Uae7wJ4Lt36wZ+oNMcWd+N7msXoEmlFsBscQJxLwgURJc361i
ZLbHDjVdxUlQAul1DLkd1nDkZtRvnG7LZ9/+ru/5278CX0J0VYTWDjjGJgovX2YOY5E2d+SAVK5Z
Wcr5t1ulHGH24fG6r9xzP9Aj119MBp6wliW2Ch/qcC74D3WHUco5k//7GSYAS8lVAAu1bjTAFrcB
5IVI8VlZt4RarY4lheehxgiYNubKzDj5tvReD8jwtZ8WyhEJv7jBJyPPc7AZFnsFt1ZOoIPe8Cn8
RAFTzuwlaVzcFeZ1JUfabrwLqySI7aDJ+vZGaSynWL49CrnK+T74iFG72jNkNHfRIspWRvOLERmt
xvpl5n2qE/dAUtsNvkjoE0lc+JBtUuLg32Qo++PaD4xmpkN6Z607fKl6YAh+3AP2viHhmTx6F1c9
aUuc3zslVU580FSjgCWfUC1rb43DKBjDBvNi/dtRaGU1TeAwNc2H5BvByRk9sAd5U7F4pkyW70+X
9yT7IfHZLAX0w2WbQHDvadV/sGP+ZdtWHzscoZOKkp81osSWFw7f235UwcRtOE71mnClx5H6TQ+/
jh52cnn5hu5jIkU5nfAlW1AuJKS/WOcATuxCog7X90yrvR9eYopat5nk7jw+cX2dw+MmvTkDdBDE
hRj4bOtJ0Si2NSFPTVq3Wdxj0Ipn8S5YTgot8ayLUE0BWJXEJC4ifOKKLchJMXKDepkhmX7ZOobv
2Kk4GJTqkhPSVr64xoBbBMT3cAsf9YH26lpVYoKS9ULCkl5iRC7ABYle5OogLFgmz3sYyd3PpwXr
PPPpRFCwaV2vMfAdetUowBOHY4lfylHF3I/Cwn3YX234qxzx0NnQ783iPzOdDZ2IKBaTdM1GiPFO
Bn8J1BkP7jsXEzCWKzKmjXOUeei3oPdpsJ8QF4VSEqXPm7hcs+XOtiF6P3GhB0ucKTT0HTyblFVD
PKLRj2lDf+vgdzrFuH3bRdUnnNU1Rhie9/Ci+UVuUuAvfLtTJuLSgRSJPko/he5B7OP7lL/r4MN+
iT/gG6VBNOFX8aiQ2ezFEjFaZx/sjXJGG1c3XLxDPxs1ucyqFSb4va/N2FRF47GvQYblNe0Wl736
Y7jsr2PA24MrI1npuBhbIWJvMAVG9yV9/mqEvkbnYegA7IL0/Kvyj5ESjNYnWfDII8lSLntpSYjL
Qu2o6k3tuTFN4YEdhHk/oBGhUPy/Zq0VolTrDv/R0UF+erwpLP2w7fkFykq297gLreTr/fAc/FFF
LCFvEpS7yB5ivpghz31Pw1qXzagDWvzw9xpJTD4vJ42S7FP6A9YZbz9WjDPuUMpOyiOS1DohybRT
fLuaZNrXl/PAY8QkL3gYwO7XZhgfQvIs3EybAJqiuyUWnCtbnxvMWPwaL4X/XUqgm6NVPSwx05xi
JMELeZ0xsCF7or0eGiChonOzNdfdE9V3iRLunzbrwcbfZfF29N5YV0L87iIwiMTM6v0s4JigbB3j
RSsTEJLWT83jo7xDjA13hw2qW0mkvVvhwjU4l+NEdYcAh8gAAkRqaPHFYoOO8wYEDAaaRNzl9ttM
1/RDlOFHIzLzJ7s6qr+U0uQp/sLnOwvC5LOI0hykaYAdmS/ve46R8mmBhJX0gBd77n40vq4zRtTk
5uknxOFm7fXdYISgHazTGDKKjbmF3MwxIpNMAcwm+jyVkCq8PzZqgrPaMdLkqw/TL8dflkiQeu8B
qsSvCrdrcD+kLBVwIbnCWWVA+Bx6+DKQVTteSqPeELmv4igVjUx8hEbgFUvRWVAMPpa//eFsW6p6
fBeC37Zcf3QiA6T42Ain1Yth0D2IkEBrqfhJf+L17+3mfGJQEtcqiddZ8i70lmlT4aHNuzxTOPFz
YnLuO2I6sIZYbjbPv7M5c482lx1xwXE3YT29/9VNSJXkOwB/MDBqqWYD7amF0F7U+xsWf0rvmEjX
Sr811kVUPfVVLKXqJ8zitB0YnaCTrlF6xf+PvJ0Ca9yrAWWRrORW8cn9WX8EvItOdMagDS8VytrA
+FVxew1X9ro6pYczI7GiSPHAu4gMCU6yHsXcPRZkZXwhhednpglDLam+YDtlxg9obyHil67+Anws
9G7ANIpt71gPYgOuvmnRMx7VYiR0SIPDPYONGiuXYepUjvuj7k4YC6F/jCp05ARgw9qxlU95FAXo
C9pG6K2EDKrkc4qDGa0xoJoFRH5WgwBF+24/hYRroaTsyB8/85kyBZXFEiP7SlbnLVhqWgtjqtRC
VpNNZXuJgG4oA+In79m1QvPPCYy2qB4M54uNdSjx0PFPhU3skIqjmf0nFQWblp1aaQ+Sg0AYHOGo
SOb00Yal5wksLNDOiv2OR7Y57+c/8+Pr7uHZrAASJi73+pStmzHmxWYBUYoRcUEF3HIMpYOfcxCO
uV2Lts6iqgSdElZKGXiwgNiYl4h3w3dTFpXUaOvnQ6G23vXTZi7S+kpkfAGNvxg8LUYzmSf8JTZi
a6ZKr1IXeiOjD07Jl/4OPJc+mjC0gUnBylo0j/AkturrRbvFa4tTYutmJ521nbJ6ZUBnt1KW4kpP
lqynqOonH3uNFutRmwNTbHqqzhr8MEqcKEixbZW5qMOWG5QkpGjQ3DDI4v3A+R4OwpXc2U39TbYL
Aq7dDPhPHWS12kC6HrTL6zNBEItl+DcwFS0Fs/DTS38usek7RZH5CPB2+4UpYukFpI0JOfAwIDtx
HVj7j8qOX4wN/ySWDzqk+aAiy9ndcz02yriAChUSPd9Q9dp/tzpgmNekDk4DN8s0GUvsQhMPyXYk
f1hhScW/x3WnvqzW8gN8kU89iRCSamt3wK3bAjOUom+Z1VDy9L0Di3fY/FukYpAMUJTpcVP71DBJ
aU8XsxDi39ITef4JkIF7UbxH/APRXLtKeiEkCZOlAX95Uccn5Lu15ocA9EYqCqLVTVWVt42skBaa
rjXJMtrcoAofhRw9KGcKEEA43n5ezV7s+gktletuQmcExgnhZWgfiRfZuFlR9MbqBIzRo25Pm0Av
KF/cuyngKsxtBJy/U8G8F0seHAT/ImCZezDCq1iHsJp+Zj36U60JXCcOuKyCq1DFlOnIiblm3ECR
M3NyfbDsaAkdAow0/s1KILiucwuSwrjnHjHLTXEOXb3NlfHrqFs+89lxSmq0MCq4LKjhjgu2g/fr
t63L+OunUQxV7lToI7CdagHa/iymFl62zzGGeJ6sVDBTiaVZXbjQOBb5fBqJTqkxDT49W8AD30Wv
C5XI6iRwp8bEHahnTTdUq8WhPKoYE1FbqIK8xlUc95E1be9W95Ao79ghwWkL6Mvg+eFYgNmZ9eqO
596uqcfLLAw4khXvV433ClGc696wOl0fRxL8+SdtVvoKjweoHQPZyXKASqiCvFnv0dMlMlyyU2nN
DzHuB2Wsg4EHQtbOI0rQWpZdAxlzDaqkWwpCKh+TpW+8Tg/T02UXz+kvnhEly2Om+tsUh7/Tvx79
Ha+7uN11ZSHMrb4jdKbtd39xGo9lJtr4+Sm1DRZy5uchWflapwn0299jsLpFUM+6wHZjX3jCzeGb
HOAG0f8+uWXII34wanweJv2+ljbJE6BQqlUWojhnqMZ6xsn23k3Le+QK8VZIfzdsxpOwOwlcnwq6
kuD8y8kNXv5vWtmBqagWf1MJ8tzxQfmvtwABY0V+0c6yxdM+E/GjFJRrynuatBqw1ERF/vZS8s1T
casudekbExlNe4FueFqsfxqj2KuNPsFPMQ3tND87Sb1I57YUQKMkP4bO3cRy9EAfw7yagicqvIRl
JPul3ZYqJDXizspMaBueCi1AJN/u2ZC43tDFEyFL4ynLtvMFpFVhevr7lfQJOivhKsTSmiOcZu0S
kCPUX8kQvt9OXFilEuUC4JNZLRfwA3Efu7kgW4YupNh6GkDVq4zT51jHyqu70pfLRAxDuEqKxu2Z
Vxh+Ji9eIyikc42HI6VNHXuauek+BGpw3rOBg90Ws88qGMDVQDPam31kxgulYP+2JInFb8xVk+ge
FHE9O586Tw07BdVUh3QHtuysmsswpx8xdS5abfgBF//nggIyknp3kidiKlh6qwkQqHLRv9v2x0g5
TWIpuTsPYSU6z6kYVso38kwxmAD6+JZ4aU6vyTszUctvVrB8PQYAAuiDUjA7uuYNkXnQjJ/ME2Yz
1hvzBhghagERzpJAbnBYtyC/vmOQM0Yoo7mM+MhKU4NKweC6k9CCuCI2C2eK/z0bHYBSQTm+ZU3C
ZA8nCsUgKLWzx/rgfiP1bL7srctwmjvpHhEIsyAOUM1lLWRaknYoQIhxqRcc17tW9rRdQHGdoaY0
7KUkZmbMwozWckLxD0Tzy1ZQnkCYUemfxbV2O5fECSxusEuSCa/ASMR8sN9zvk/Z11v/bjyqX2Cf
KxH/UsylLU6yA0Qb33x30QR12cG2NmMoNwf9VctlWCCyy1BS+YMpmRo83z2fwnS6L1F1OcXtMXgY
DaZuRsUjMrbNZ5LlYG0NjYNsuGOtVVRlZ1wAP/RZFCL34zNxqS1gzSOyvfZcm2+G43x1YYBYahm5
DOyaW8FWNyjctnin/8N1aTPvmI3Tc9MAwc4R4nT2AMkiWjZ0JJPP1ZL60Sim+Xl1/J/rQ7NSsbXn
lMuxYCK6aH5MPJSXXWXPhP3Fb6GaO25pn/Zd7KyncYPGgjGbudgcKa37F2lyTyrJLpRpdm85cr/o
dlCjBtfSkcukW3XBw4O6nBcboGTip8Pw3fnvS5JwVxM1zxLhYGR4xxt1Q4JIzGB5B1mPiFQxPLaQ
wp2VFc5N7YiO7/Ru9GJCunKC9VmHX/sZ5OX0u04+yJXWip/csmuYEslWi/F5yP0y7O+SLugq6toG
FpNRWM/VMUXCNwM4gQeICw4nAq+mfSghJKxK+TnYi3ipksLWHvcVz0mq5LcoR+MirSlsYaxGjMyh
EKrOkrZxZ7+14CBCCCFsQDmlIgr3c3zRjBM4AYaF7QJkuoAs1lPJ2j5gAxspJ8JUOC/KVNOTjrIj
YhOh9/jmoabpGlaMAck9nDIOPNGKVxofoT5pOcO9x6Nm5FIQEOCIgld4MJ21DTvDJnlrnmIL+qCP
NJYx8JkX3HQKLWSnp/PF2TIrcK8yj5jJ79atN+4AaU5vj1fcgjkb5U0YxP2QigI6e1LkmEGRKvSN
v4lhemmf3ShFIPQumZJ4d4ufiB7aa7I4FAYAXrAtBqyLZXnfLvFRpq5QScHlRUYkC53PZ2G9AScK
CA+PA/vGCJaUZXS+iT3Ndjia3IwyRwLPw+FiZFJ6BCOyplrn2D4vPIseVmhzeeSF4/iiWE0WNeBn
PUV0Fpk8TAbHhY2ZFkSGrZ11OxGQhF6T22L9EuoHGlqWjgVHmxM8RqwIxEhz8LzCmQRuOlP7hhar
fPPMiPejVLizIZ5Dz6kPke4CFPUM7N3UJVCF9efEX5hyuQzGFSyJ6NP7V4p9huQjRp3ycIO2ojIn
hywo9AKgLSdR8y6fqvvxbujGxkbtwywWIzyWm+9uM5s77Jt1TkWEH+LbsIkKwzVn4iprMvPaIsuA
qvG0NqcP31c7phZY+IIpmKVQXJ+ttz+B16pjEgWEQ0zW3WDFyBeuQbQEML7j4vfTpdvhwzBShuyW
blq+8eHgI7vumXaMNoOdyNSaiFoeSSJPq+JJCbBaUrhZ4X69WiTDWLwLuo4KAvl5n813wiB0xtKm
BCJil1l2T88+8gajoWsq3f7XQbmVjUN3CVqxQV4Ny+OIo9t00KChj5NdfO/t8dj/mNkSWT2CFJ/W
fPBR9qAdj0qblzMeObcwZOKzjYb7GEMsM3yEOIXDX06d9Jkz+m9UKPE2OjXZMSsd29X/S2dZCcbp
kOGygN3bne72cQYHM5DHp/doxirH1XS+aQSMdNP3mD6KcmrOaBhhjAO4E4q7/26OdtooIWZKCTmd
cq13CFTguhd1BjM0CUX6Mn63s/NVoaMge57SVOA1xTynIKssCevs2ECPj4X3npkKvJ5CRLo9PSW4
NhwCuvh0PxFFhkDeBEDu2I8bLhAPl0/xOLXXI0AqF+o578VL6i95qyGXszB8iNkF8Anf19DU3XWO
8x4R/Hw4CaH7WrRnfzmrYy2hrVls9pCNBzMIX+06PzYxvqQDJVTRcgvxjUBzOWoJ2WiuXJ4gaC4o
fnnWBsOn8Y/s/pFelQ+eSobi4OxtBA1kfS4+tGRAVtcj1Jcpj655+FNc7ZtJjMiRxSLYNq0laxZf
uKxI9CqY6jYzMPcaQMhVMd7o1ZL8J1T3qoZML+VKg2VbTa9hVt3wihzxhlPpNlmK0RUZhpLv3Oz9
n/ruBBeR79jSsTfDAkniBTpabLTRntiz6kkVm7MimWx0O9WDJ4G+k1kI+BNkHfvIWaVYSpIxHs5s
44Faj8MzhpjRItSrLqF4nLgPGTuoBTSCaFk0GJKTWVO1SBkeLN/wr9/xN3dvFMdm7UK427YQEYkb
DofvHbI5qKJ1O0h/ODoScfaTeZmFq9uXEI2OtmaMPFl25905cygg4ZE5+Qalz1m70i+xGswyf+l2
1HNOq7vraecTa1Rf6UJ3EKqk7R2kb4UBbjGDGhqDC7b+9MehGmHn+JLCOuGXNtHZHcBTanbWDr5M
i0hgVtltoSAOGs9K1RA++HSxKE2/7nyLb3dwal74HyZ8Lw6CalsW7FoT9uLYiaedVNte67qyS6u9
yXfhqSlsOiV7wohx8IOhRHZ4pKO0gs8bszrtI9zT1xoznP97Udak3BqpgWUSeQMJyUPxhzz/U1u8
F7mjRS95UrJ0O8/2uyGFf8MV1V5D/gFWseNUCA4Y8irq9U/rfAGEyPHlDnvNIKgZOfGvHebyp69k
8TnUZhISVATvklj+uDQUK5B/FYhtQc13E1NVF6QwteMhejERrKZzeYtfhFq4O9KmvBLj8wxXRJ4w
A8xFR05RklPKl5cFoJwdpaZDL9neu6svAR8FyfhN9WewryZGSxvJjdyZV+Y5asdguonayBikLNrE
s/63czabZmuFJQkQSSc5RP1vAUgaiIAJDj3SjtGmL2xprtmmcmDpDwbjvjMtMPD0cM3ayRhpa0ti
rYKCb4T95CAzhWHTUVhobLtj5Z92kSQZ90aJ3VQyfwJUGZz92IcU4jGwIjXm6K2qSHYO9PGFiBx3
5wnHZmwnskO1xiJWtqikG5NQluJEBfovuglSf+IjTgWYXsLHye090SuD6jigq/rL6mED9wMJzT8R
Bayk5mowy1yGTA5KM/06C3pTF5H4VKSwgQRmDY2tpCEAxBfHlpmWM0IoKl+RJh6iJHLXCA146/0Y
k1x7FkwelPb7N7KD12K/dqzOfGZtnuh3XgzTczLsEGT6KUzrAO3RKmpdksosg9a0LkB6znSzRPoV
JZU5suv4D/P+VPGRZit/iYWweg7aUfiZEROnuamU8lfJUq4L1E/I/s9ZnHbzIb5e8dHTP6aQLXxe
ESjKm2ZRBu5nYh1Tfrz+gMroxug0IwO9Ev7Dsj7GC42AmhK0NJ77DwbgJOwL8KyZ/QTD3Ip29kVF
MAOpvG8+yvzIKXAKXErVvyWfgOuwQHmLH5NKZtrGu7lDrqlkUivBHgSkIJfe+eO9SyIxzneSvZMa
s/DKB8VXA0/luLyEk4q8Ok7CvBcsfi17G7y3WoSO/zJSlP8fOmSu2QQoPe3atXNrL6ABEkMAICqJ
kJEwvH3nN1aNGZgHPjxVflKiX7lTZCKgJa4kdLgap5IDXxvVVQqT/VW9SNKfiL5JfSN67DdG8fHt
P6p3e4NihmvZ1CG3kENLA7nTNt8PM0nqcwthZrxEbblXKXpKWyH+ymKtUkq1a13pawKDgGhnogZV
JBMn1H6IXqImGmukACh7GJZvjemnDCnu1zKYSCx3NobXcL4QrYtA+hGtFzA4qCPN7nMvubIssB3b
e8lsIV23sYNTQ83pLg/FqczR3KVROjQuqJbTcXOzFydb57niXa/KXSj5fvT/DtbCsjy/TcuYANum
1SYgg3+Oo/x3FW1YBKc0l6H1SLry5ls+DJTRmain33tN0aqldJ/sv80hA/6AgEY9aiN9BU2yI6mq
Hd937cmwsDkX/4vMQGL+6edBDMJvenQ6iEurqQZOCaEfMsHsH8Si7G9pywrG5C6EECLkhtSgr6Oq
vU+3RAeXDlCyP1qcEihN05+GT/pX/mZPimzl8Tq+SVpx/k29mNZXlh1TVSaEGivgjc8rMfvKuSd6
0XHgyFaKkF1tan7IxUvho1aduSS0ZDbksct8Fv2ZgCmk0mR8zT2ePZuQFpu7kpk/SNjJjXcHkQYo
jqVLa9+a0sf3BKULxWDwbeOVaVlCHVxyXaN+A3ubNxY7tQe7QgiYEahTmZ7okZseS9uderPiaBol
pnXYGj5RpSuve0sTpFZR49/gGtbM0PCilcv8q3lS96ZR4s7QobaYCCH/83RNYACtAOeTSDSUqMMD
p47wuboQ2OHNMmbjL5sBOyUylkLWe+APi1GfL2qX8HWmi9W6ENcn0N7dAoa3DLqoOuS9hEkvZh0c
nOeb66OHFA9PKRwqO16gaprYR61zol3iO7UdLnKfgYIvtOZ8zmNCvLBbPkQZ5hSHjhkJ2cB+Vz+B
4J8KbBngFQik4UCyZsgtf83ZEv113iaaIuFHTl8YIAkEiNSz7mSLM/TOYTy1VrLAWiIN/NUomQpA
YhB7TblR4PbTFIZMksivn1Iwt6cPC0iiFpKNVoGD9D5WE5egte0VPBL5z9Oc3MIW6WENbjpiargc
E3oDSWcREVMvAjM2deJg2kI9UUCMm52gF7Y/TsdkbdKkW1QIy3kHc8WElf/Fzt4uc368yPhsglrl
p6Mb9saj6lNWog3HeUw9AqsdWNs6JLRSKWeLrOcklh9ZOTGAsPIhXPJrPdaLehXAbLupoYhg7pUT
mTplPbtD1unU/SaFqUeXIdzfCi0YCaYfyhlAfooC8oxaEbCxFZwaCHwJoeGeiqhOlLwHRn8yN9OD
vR3g2OT/+pYq8KWjCZ/8OnKw5bAH6tUzqVS/GXrmOTYCl/iGusaTbekteiAbQYiPTQsYaFBQmbHe
ADDNe8hrx15xDns6Djh9oyY0SrZVJ8AEgKWR2/Bkj8YAzBi4d9ygAilNiNl1loh1fquoMJWL/+if
PgF/6THUG7xvnS4CGbOPms/4S37rl+afTYD9e0uco54GsUaMQhtB+QDeQr+28wxXqmOS0F9py4+X
jWe1J50YcBYf3q4FWFgzfmMwgiy6iCe+7eiWIOgKPsjCKzLsZtmzcQJvdUwnf2eIbISxiKbAAa52
/DfGst4/vHJ51HsbzwGUmx/Z3dh9C/KUYckY1e/Ald0sCeYMlynyOOrID/MYTE7/3Q69rcoAa33w
tBIErG4IS1FnZ3yVg8iItDoOoZZX4FY/KA8uVAakTiAfrcN5nwtjNBLy39jw+tg2r9LUUkJBZ2XU
TMTrYJ0t6Si6UkvXutJ/MBzXx4QlDDmfldd7LHsOybDNAPJ9AqAsjZUokB/oOHAesJcIqtQq6cij
NtaII5PEKl5PUSZhHT7qH7XTq7fMAfKhNL3xFBGQsLLDttFcRMspDISkn+XBw0OGFY13qAbsnjwC
JH5TuyK8hgHCTSEEfPdJGpUpTxWFm3oFZGx13EAF8UJCp2hnN+DzrpS3JJzoyIE8xSCgZFifoIeG
2CzmUojieK5DDl23HqmRzpAu3d/O/ZOrB5ehubPxB2FciasMEPxyc5duHwmgE4fOcH1QUgNytPEd
CIFpi3cA7yuNj8Ay6MmlI908HisrI1MMUP4wkPOhpX/hAQvHoRgWx72OG60SNlSDeHZMmhNBpN0t
0PL+//XmBWf/2ObD7vDwEHqXadkZf0yo+AIAlBaaZNtTXvvnffS1D/Rxd/eKXdFfLt8WJwXcfTZj
5WgkRJxJGP01yum410UW9g0Axh3g3dpdseD8cWo9+Df+RU3/DQIqtmPwztwhKwvOKllf2m66hV/r
jhojRiAZwo/g5buCn/NRsSLYsoSMNz+FB6dKY3HuDCYlyqwAKQSKarg8bVHXnFnucOGLJzELF5g/
jYYAKNUdrl+pgpRQI+YroCEBaCmKelxk7zKhx7bENOIJjjJNyzi+HUPS51sOfAtnFtaeh/P7vjlA
RrVO+M362hNqYJJ2Ea7EZoxy2v01FNWluZ3nubBcKpPbKOpzMFR14hxuPTBYBHoCT0m2hGnqVo12
adi13kJqWc+WeiUuKE5biJjRA6rK2widpkoUfeyO7E9kiJp8GiLmiG0w1EXA7v83tKkqshMtdQGH
5DUEFtObRXUQHZnI4IyOAOOcI0xplfDYwQ7NAoZlXGkwDNM844BAovM8O/jsOsocMJKhoBTxC9q7
kXifx39WAjfE0AfpIDfWMiX7nQE1KP/D30b3RzN2DEZfh5BzJ8Ug9DXNoVsjR3tcZh30djygsG3W
BX/RZnXhAMLMIubspGpngsvh56638u/eEfCYXmHpUJHiCxsxDcQhA+yZHKOSXfejvZohgW+QneWD
qY3vzXFqzhBiXQTrIPBEPY0Irk0BcHDU8awADmRM0ITTsSDG4VKXpTwKPPwuRYsYyKudkKCyBzB+
cmj9YfrcXl6ZVizfXXhcYcdf6xl5Xe+LJ4qyLKDht/vrnIUpNoL9CLiLIzSiYlY5CruxnL8x0Ze8
Ac0HM9VJ0/hmiAv/uE/cG6Cy8lnXUukNxetgCekoLJXAXQrXqX7scBJvu4+dIFUzoK9I4wUEr4M3
AQYPgmyjRuJ7UF2J9w+OTEbTX6K5Gx1URmPKHszI3x3tE526eL/4di94LYXSlCBim/Kg72/5Qe+t
SPldjDiClE4kHHrDeV2+Zxi4tnW7uv8Nooc3fr5Cm50estSR01Qsqw/6uj3VTzg/pgalfmgMAcWT
cniY6aalpw6jw48bjD5J+eKY3Pkg+MqjjZi0F0u8QlISES3LLH456HGt/AE9RP1PaeiMSP5lDSGf
mUy3bSRelvpTidVCDG7W7B/jmxYf/jpHVw/D/wPOCrX0IYi7g8qTRR9b6rFSVQcUETNOBsVrfE44
244rbWWr2arPkYF4MvET2zEygy+jMCImRPdz6PwNA+eskmRLpdObSW3bmJxn1P2MKjulYy6ClY5d
Xeeuf+vgJkQjifR7RCLfee6FeoWy5lErWjYc/w9V5L5FXapHSyx+gNpXhqCIqZeRPTl2WAHl5ESB
rSUifRM1JMRFwrnP9/4OcLxKxoGqVaIDl4tyDi1UhHacJSFcNeV2N9k2DCYFpncb3197CEw5egCm
7YOaffRHxTn9BQaBLUrQGUQOJe6mLVe6yYqLA9KKLKESHL/Yc3HKdyefnRTeOpguj38WTU4Og5di
1VQTJ6HonqLmhFeocNccOreq2elMk2FB4qoQJS7HeEaekxe42ZKCvdT8eNNS73mQAXOJcDTiLqDt
1wB7tPbParT2ozvOBsMjRTiq7mM+Vch+1SheetNgZ26eK8c2gxo/f1tgh7YbGORSJdG4/i+W1XyU
+R/PBzGHsfNyeUKcTYcsKZ+JJ8E/sqSERrSYh1qWWhad+FKjxr+CqFisJ52HzNXdGSGydXyC3f2n
a/ZVWl2muLZd8J/6l2cPdbFtvTmWXuB5ryYKc4He5WP965LbXhQCgWjHM+kBTbO7a/qdEvU5gLJ/
0A8RsefOwgfqLoJtLxtjztBtuGIbabmmKAPMzGM8hywD8bfOBkW0vs0J2q7/kCvX2lGGoWlGTBfp
p/irBG2sLPwp+3ZFx27FPuPWbchB1OuRpfcl2/Z1wcTE5mM+nFTFkO//0eXk4xLNfQDHj55ggr0B
0RATeHAOxD8m3JjUhgjhbncNJ1XlW+TwZp42hw/Abb7qlIa3JzBjwIxJDUYc+1qz3bg9ShihSeLb
KFDuYy6VBV7ImdeO2qF9DHGV/DuTiIldP0VSs0z5bqkXevzBbdtoLZwW3PCi3qgF/hiEpZfDjBzm
0BMdE8mF1CXuxHkKer0JyABK7oAwva0MB6rANTPNcJ81eYGYpGVCbK/eAJoTuBQ+Quy7RdGlunSh
gBL2xRGIHakG2nX6XeoSETIlh35NfkIv6d5jdsPXgQqeGwbF5OqeEbIlEcsjNi/wfpALNR7l/VF4
gMD1zlElWNRktj6SkUJy3BwAL4LVzUZx9KtHG8PQzMYAHoYywS33v6zd9heVgWPu+t9w8HkawoHP
/U9+sUinCm+8wa+Stl9b8UIyHicr98YSPXLicgExtmLliZ3bQZKv7Rw2OSzBQEQI9GcW70erclQT
9Hbi1603+t60iuKPsFCnzgsiFnh/ou42NRG8gSla1dgNdIA6DvG0ucacYGLfhqnEFAKzYCw27T7H
+OouAL6I9RfhczNUww9SCmVrjHat8CfyAlFOdxrz0Mi4M2/W3NYQE0owFDPdsCpG5Ywnjdz1E7XI
vQrdMf36k3pZe3Itf3R6+8EQHOSWWDzQWnVxm6aElom6/zDDj6ljK1XfsBPQTwtl4czgjpWVRiVD
BOVAmhXnuBFJqUXB01jmh2rn6OJARYWOzOh6/TyhZbOAvEGCv4ZPBPo30mXFsydNerzVAxaxUBGD
fZC9EzBxcBrreUlWmXtTN/U3/SQ395zKcAOb9txYv6mah9RslynyHFNQJq6YvZ992WNwZFjtuE31
QaGiEBTXgYvjvF2LYDnq+x8BCN5PYw5YtCME7PIwOoKJ20vXCvt4bePwKBGMt3sBAi7BhdSfx8ut
prtFHfhUG9mULBYOW5KNKQrTTLSSI2LIoabE2vtXoA1gbO7n1hCZo0rLHals/WRvKoggV1aumYg0
gkPfhOgCs1y22Yedb74tlso07RBPA7jf1ZhTk3/DAfrCwfdX7sAN9t/0P7MSw3lQWaCiAwJDI0jA
eBPImB8GBJbN7cWXGs6TdQzwRipaXTgrJ1QjZf5loadIv9GovSW1sw12uXcvec4OPiYsBEvxE8Ad
pNqvbsL7EodrYVB7TrRzG2jIDpSX6m7JacHzSR3KFTAwmSr9tS5x5ntWA+nNVaB9/Qd+zoQxdDiq
d1VaYbj57ZYV8W12AOqnvYCdSCAIdHu+I/8b24cL4VjaCaAtjh1QF7gU7Vd5kIWEHsd4L5Ec/2m6
leZccGGSIX25uSVQSHNgwz3fY1PDDvXuaE7RzE2BqHcudRatHjPfDJT4c6TbN62ZvFQdoj9C7ov2
48zjI1QwAJATY7Yh+9aHn3jqi2MdQPX6PTAsFS7XhNMkjSoasWf6fpyy8FNU52g0rgwLVa7Jo+Ps
MEp5gcpcnmuN2/UCucorRpwagIR2pn46l3MXg4ctKFFtL/GJdInKN4mucJtg9zRwsplaY0gCaySX
qU8KSvju8vwe0QImL2jsE1RwFxR0Pqxwea+bdcPQAYG3+CP3EPIPQ7s7r93wSRVc1SBAsptiJoxI
/0ZrERCKTO1JWogYq2AXkJjNMbQ8PMdRT2IqCyMiWXqF3obdHIV/G7pxqllw5mn3mUa5ZUFJj4JC
md99Sq0ullBqRnb04IE6Wg0wbtG5FpgUH9k+WqDkxWY0d/m2UQXTBeO8Ya6HucSDnx5hlTpicTjv
3bGig0VbUFGayFjOa4ZGVOUsdXI4Vx+AxS6/VNQsj9Hgpv6TSlcbjl5X6AbgYXpQzlTYpFZzi8G0
FAQSn34qdBWCzz/KGg/sb6jefLXi8y9mb++Fl0fGJbCm/FIoVTgcgc4Hg33JEDo9VCtsaBzHM5wr
SH0J9eB+Cb3R127ctJjeblmtOWOIjOPbm315YVX2y/Ycjb62Ki8aAPx2rvQOHqmHGUIz3Y8opuHg
6AkdcQsjPc22nBnDsw2b7dMWJJ0F8yz4puwGaXTukReHFwJeI2h3643a+7m8fDvhF8Yk9vo8zMsn
NDVtU5l3RKbjY+uuy7gHFtQPHmR3plT1kg9esz0LwnUOc5ACkMgIfEyWWuU1ss7XMZ9n8yK5Qzc/
PVr3yR/JF7Xv+SBQAFEc+l7+OKAfowMEkGO5PxNLJhFS/85jbUDTp0/0XdCfI/1vcrRtffVZVeFB
yIhRey37QndS184vnV+U9y5Sqjy5McM576bkaqwLW55bgwRa0Gzf4BAudr6hyrz//qlHWP4cCeMw
CE49bO6LB59XIOutgatQq3fz7Y36DlmtGG7N9aKS7Q2WjILdjTz2uI/SEGGezqpT3zaTwY+6APeD
ckF2bYcxoXZTmXnAgEcQw7Dk+8dm/OJbuaiA4XXvktg05xpG66GDzyoVFVTB9OowBDeKUZOz87Rt
AG3uVY8RCk0tsF1+EVGkVxGppsckFThOMT+Sb1iZlnEBccdnVqdRI30ioj32JDoMZeQlY28ofuHn
63ujEys+PCOp0yI7ClBt7OQ0EIGxL8uc4y4yEIs0iqnUVWZKDgsd3tmSDcYzQT34fjxxXIqQpUaE
G4w9AJRKwOSqrKiCGJ/mo63f6diwlhJT9H+aHnaI/Ne6Vl4QzYPtX4z1ADirpsNpjw9ubfbsOXy+
rgEEvXhfFp24ky7AWnLr5OPujC8gc38mQbD7301n7Cp8tqzfHhxbQFSI/bS+K5Rd+F83HAHlaqJv
MWg34lFW+gRP3LzdRuZoTY8EQUQe2lQgBxAVWN0nT7FqzeHJcPhjcSfAapiRR7+spVebNopfh2yd
lyj7OOGCZAgcQm+IfaRvLkDbUJPfQGlgn+XE9yqG4UWDp+Mz2AG7Y6ZvLIurDHMXRcwp6ZWZzSmK
iQ5ayplTsLJ8rdqjQu6NVMn248QsJx8LaWc+uTji9J1T393Go6tMkXWU2rJFi09NkvsCy0CbqCsc
EQOtAQ2WmJAkOfiFTDVT4IFC+mXxKDItPed8w/0tsXgmIis5yVLo5nbn++EgwlEKznhnVMBtsPcT
algNcS9KDIliNrxkSmEKdLiNU1l97ZT5IUWmoixwYDhYDKAkVf51PJaJZTyl4AAwIinu3KY1bf4h
KrQrO+yvteROcsNIBHhP6SRFxjA5PVT2zFnhC4/3Mp+018qmyuvtYBSkyLOQablCyjoqarswtIlH
+KyJnL60byRfkF+hMaxYZR1kj7qeJheR3CcxMooHrevrAeb6knzLK+5ngFwUrvLfZUXnonmijNzy
aBcJV+eItQvUIYb0iblgtpJhT5WF1DxmseUbymESuGeXFrJBnxJcBbBGkVC1Dj5zIHDw7ZTtqza2
SCDLl9CrOJ89LOfcNlBHaaxCKwZeVYYF5gj3tLvTwOfThua0RLWuSXjsr+eSG5Z90J//FhrQzjn0
DCOaN53OC+Ix1tTm7jnzKVzEqlu0q3IoXQJIkvD8XhOcdaIm4Fyjj6cr9ij2EEh3psBUewuVFeyc
/Ivdrt+TFneimOxN4ZCbL9G71IvVEYjBmE4yUnaa/DYJ9FvxXuEIhG4mqG2s3NoWtG1vFCrplT+k
jU1/PNLpz2UkXXvmSgk8zU9EC4ofYvw/FIOfJaslPYw2P8cPFVUrjlKm/CNsvtgBFrGvC8iFIUsV
z9pBuCdkVnk8/t+/iI+dupKEASNWTZLPKlf+L6OaSWpQLMoHrH7/Rxrsi04wyzA9Ap0YlmNLawxT
FdrMEZgHgblgbVqDmeltWWVE4PPBnEBgJV7IKqEWhIv1YN51qVWVX++1Lg6s2vCsO3UFeNm1Vyn8
0Pk4OXfy1TIwoHtV+pHUe0dXh/rEupvYvmAzqVXoHtXT61BkfIDF7LsPjiICjW1fxHdpnXlZJKiJ
+SOSO/vbF4oinRhzZYtxI68SvPdbDLMzFQy6m0HYurvL+pnPQGaEdsnyeKT3TrHRbOou3x1bRs0N
sH6wqdh05CYjPdayaHNWIVNk+RiXnUvp2GuoVTOP+HDM184cNlD7Mx9F4d2N/uMrJAofc/iAsUlW
V47rjxICOZeZ1cuQiA4+HPa+tl0+QBK0n7E65OMaAXz1gB3QJFqUb1e/sAj+YtCf8Ok8S+JQWLNX
L9ladQgNkXiv5mVJ4g1geOXwg24Ng2S0oSP+WdtJ3MlVFy4FtoY2WIky6XOQm6XI6WL4Pq91zCWq
LILSegVTlVDL+0z7WPgV3mUycu9D3/Bk7/rPYGX3tppTfUKpS6fO96DnxtmT/RQtuO97pCQNCMKl
avUvpnguPqmMO6P74Yd1mO7+yRwSbJwCHbIHktC6qvnklNFckmdkifl954BkDaPnrWWLues6rNFe
92TVuT5OESSbsTSwslqSPKGVtYVp4rjbmQMUmyVHhpTP/1xI5GKTV/JD7u3wE1d09TVDuVoC5+ww
wvOJTHsj+HztNWK3+VgD+NDVA2xDu7aGb13FGalUpKfD1X2mYmzl+99KWdYSyseLAmaBhNn4h5KU
1dMshywtNlfUQhEb/0C+7/SH7hQ/Q7GufdcIi+EHARVQtwMb68Zsc5zArEkO4KEoELl+Yd0Hi01q
cUzp1zX9/lN6fP6ZjaHo9IdQOEH+nVDRuAyVzmfe6JtKBGwWT6E54+XkHKMoLJAkeCQJ9z2sXgo+
wKCZYZJq1b8RiF6mCi5YV17RYPTD9TMGOJ7By7rBV1xaa8sepOe1G6BdZRdmNM4uQnoR9uZLvuB4
0/W126a5tBF6HGjKsq88KGgKBplyM9WlGfF1yhOsGSWVOQ5VK/mRtzc5K0wEtmYP8FWicILwBU4K
DX/wUjZ+MvK5Kwu988Ng9S3XvdiieG5FfWLd5WiBqzJDzLmQYRJ3BxedApl26GAtfdRIcu+YifBH
Ppk0t+zMHiM1jnRubstizrsfkPyIZUw3BXqkkAcDE69cfmQD619dEBRUg9RSP3mQtZSAK/9qHGIG
4sHRrxyhzS684vopTRXNifeRTAFGwzeXdIP50qpzzKC5CUl5Pp1jqpXxLTERqBULxDwBLEglreSo
obO8Ib4pk3wUNoLxZT/iQe8+8LUa9FIXPN0EZATqeC630x0dzXOW5VWndyOvwMZUDRfo72Xzmyo9
7Uqt50MdHpd/WspTrI6b/vXlrLiYVuF3oIQAzwTzxPO89if3DprC97Q0EcqCsxdRw4Sd3rSwzS4w
0X5jOyJWXPsWKnVWoq7nfng+HfgF0tSXqMMVQJVzec9Xx+tDQ4V9xbxC9ACVT/9vboAkhJjCzaOy
CoQad1XiLBkQrhCrKpzK+NjA/0sZoZy06zbHioK8tY17wDHoODx2com2DaXwhS+snvxnyFX5sYpk
J95ntlJV5fsVZXL8CWwbnljH5DGUzd/3aoJErcm3tyc80/7aNY66IodUhiPUrzWoZ+9HCubESJd7
DuvEUAQpnmLM15GJjfjP8LRxAX4aRPvB3hHnCLkNFs68BSXYD7nW+QfpzL/yeMVQkGYC4gvcvpcE
8xDz+b8vRlvuajJLTnKG/tyEdZs9v2Oc0F3ygOcGiJ9QQHu/8oarx5XkJexpCCfX0o5RyF5StaEe
3WVXgtM9OHc+EkUOpSTrBm0ByAB3Nln4fKS1HZOGTDjjn9nXgRaplpwJLn9uxrf3k3HYZROs2shn
19m4NOGqW579KIEqC+XE3rPh3VlcjqnLLOKb6cdTT6TMSFTmmKu5rPg/e7fr8iYCKotdAwDtZECt
t01PpP9Ug70bhXPN8feq+eiPKpEe7MmU+8wikGDPf4ZyLpR9rN/Cw10/vHW4QyskoxiOMoslYRgC
5nARdkkSuAmvgsJ+ydEo9U/9DdxVZ94cgVEPkvQuDkzbd+TIAeV7Z+SfaByUF415AvSNCpwt053T
edCemnOU2jqYpkTdkFwCkg0mdQNCJjOzocZrXL4+RxRB0atTs4CoC52h+HSls2lm1No9BBCnudV6
Sd/VoqF0V331XUzhUFSAjtEnbw+NgBFYFzKbv9gQWYc/F9sp9oCmE3clgu3hJv1J92qvlnlhAomO
b1UDtNRDlO5Pj+IJlsYzSAmTvokAZTFDa3ayFnBW78SW8TbHypMEytOextYB1+oGh73FXvUJwxBE
+GpsE57/idC/Zsq7oMSoQvSD2C/msZ87OIbSBW8E9klWi+keVqxA0CpKJBIDcXR+y0k+OCNcnZkd
GybxhCSQq6WsDMpENWf2vYBcjkv7LrUX4Yw9llf9mSmgLsFnacD7yHGX58iFBoYZ8CeuxHC3Qasn
A90oiHuDKhKRlmcvu/6mjr0u6o216sFSOD6xKJGkEcn+uQv/Q/Yl6ns2ghT489r2/QKqrGG4sBTp
RwbA3IDFDPIevdLfMcAlCW+bMp1RePfi25i14zgZvMImggcd10s66xKFOWqbL9iTw6YE+5U+rQCF
XUIdZU4K7ot2yS8/kkWBXEAVnhQjwGWX5Ewi4XHQP7YWj3KFGBXJgcpHP/fdWt0zx9nm5aMd0D9l
qiRtT0MrfQ0vVcRtxVFHZ1FQpl1A9hEwLdOCMIQ+lS7B7KG+oUnrBuOxO/c4qSaDfzMeI/gA5E0o
XHL436gD1DFut8kEm2kEYaQ00zEXRIwgvZFyFxDTcKuwR5RXPBvWXSkB07LsudSHLUBCRMVGmL7W
enRk/bdQOq0Y/7ePme6dPcIAlXdiW8CbS28x+mAgRKygXVlEFuB941RQyOOs4pulwPDm6rzG15IB
rVHIRJh7yA0yv2LxTxYKnPy4WZW6Uzl98/byx9CHy29nb2X+/C7udRrbWgXZU0D26IjskvWagJsN
JiqFG5UwxG7tSXMtJe9qp1vXCZbDlWx0zi//Dx0af7zoje8JB72mDJU5MtkYoa9ihVkRvXeukBXL
8ZrlzhU/4WUtBvG7nEWPFcF11WZ/++E2/2EQ+I2PCiDPtRnYZZUpUawv2FPDsv0QQBBGrUKapN35
vGJnn4fTCuKAOdD2gVgvUd051i5JKwGM/PLjil8VYoyOJS4YLIIeqC7HyfgXNRWqk2yDTq9Cc4Fn
dhGm/2Xe958Mn/4B53df0u07x6yiC8GgPNiq8fY/C4WVAPspAveMOGjko1B+znyDkHjvOjTXVdER
RvEVYrrmAPwtoYiZzWRrg12Ch1qmJdSn41T/Ylc3plxY9KhI+vYU+dj4rq/oxz+ISLeAcqzxxJow
c2wRPK0ucNxNy/AJkobXtDPlnAmBVk7NtsEqEgPDj0FLfzCFbH4BQx1yjzJTBxcKFHXpY1opDpA5
SjDt3it9qBmh0M5SYZSwzYZUcoKfSYuTMCkjuar/B2gsKbFfhwvsMFQ6mL1+chfWCg8s/SZgErdU
JH4cnIBVc8PTXix2y+9sxAfyeH97yhE6WcgEREg7SM8X4WpQrL7LR7ekoZebjb9gbCU+EuYfBaIh
krCUkTkStmax9P2x1vNc5CsmHfXVO+hru9L6J9VAfeAPzxBifnV9MC1hZQISRjBZ9fFhyddlqKEo
jUpuW/1y8uKEyQuXUfHhO3+7ZTRSlgHfoL17z+yrPV4N0butrPEZHHKF2JTvo2vjKkJ/SFenYTUI
p1A1r0wiP2+xbvmwyzkDQEJb67DAkfw37g/eEhp3xgKYEsi1TJPVDNKNNuUCEwMG9bFZPUvI/pP/
UVvWChfMVMF4VyDrqSZTRZsFcxrwB0ZDn7/b6OYlhdp/N94R/+orJ/zUpNUlgFnBOE98dJQxbI3d
KsVD0NLMN2c1/z4PymLkZ/TBxjlkfaTNdKqGs4xGzsHrDVA0CZWdA0dL9jIMnhEbuDyRvijP7ZDd
obNlKef/XlCIcDsr5nplXUO73SlYo5USVZkhVTGqq//MEXGkDX5Ou1QWLE10MtUNLjc7MlyvAHaR
m/2zB+1FFFHRaMBzFXgMe0gK4mC1L5ftcgzTWb4M1x2keboB0T6azOZ/BWD5Pdsd6ZWEw6V7fb+8
ArjetKJjff2moT2rw2NDK9HkAAe10HlgpbNYKlEthm0TWlahteug1I5egpV3kq9X1EESOLZGh6SD
3xUYcOKl7QzgCxaKi/x+BD/ulG0kon/9GV7HO/DPd5N4PLZc0hXCp1F/mWVqxo1RGjmefJeEF7Z+
gBtJPXHkaGGdEOUpdqbaVg8TSg3TJaOxz8m7P7m4B37r6t3u+IHaJwbfpf7kLylmQUB+90v1Fbqa
6n5VulFaYDlTCUEh8Zx/MFrEmXFGCI9C+bG+b3+6kjQ7W3l27aZBYxGZoEzcfT+MUukIlJNC7nCI
ehLhVCsG2Y936DQfADA/mkMlmoTLYEkL8JqotJ5+6l5tX6pjqcPRUJ1Bb1yTtv5XGauTjIvBetBN
4enBX0PM5EOjCbu/iZlpmjggeHwv7gmdXWSu6UbmCExjBqEu+4OkPhS+dShk1dR7TOKyCxURmXQQ
MeyuHTQEFsyDy2jBXDt3TL8SDVCUxi4Ejd9wNyhbujAEFRJs642OKtQ2+94OQ1oMdO/oXWMXCOV3
WvftbeYS8P3e53wwe4c2JGDZcckWFAT+donJWgIKLKqOUbmWnHHmCLj8JVnrf9C4pdyGBAiWgP3C
8IqHYTV8BIVNroSJWVk1mHCwAdLEEFXWyrF1OFUVjUGdrwXz6j3LhtiJtlHX9u3HT+lIDFtnyirq
m5NuYLCRXZGQXh/fHe8wU7D6aPj8t1WROfu0dO6Ij3JlWCsX6yKq6D1uyZjln2Bum/USVoJmwCCz
y5A3bYuiUzPSd5e5jSG6NYn/jqwzdujS2ni347YAl2i2myCbpREx8yaphcIWBfbVYXDfcNXztpcO
AO5NnNn+MvvIFnq5+3bBR1abS68L8f4+Ed4kPjvWqe/NhyBSKKAMNxLBNCeJAlFdwJSwWZq0mM4F
O+ibBrxUE7s+VLvA0pJu8fmQQ8oSEfGXmwHc3YUFKaRABFxVxPQKiUSegn/CT7AfXBv0p2b8LDvx
w0btsuk+jGfaQwPKBhgyG59EXuMWOuK469u2/HQSkH19nfVutFzEj19BagqLXbV9z5apeSPmRKuA
pK1H+Bn3C94kiXADxJxEHlg1NQZmV58SbmsUwmMgvopPgZ7n+/UdKECf7CK+S0NX+uI1mc2qGT4d
AOu6BBudiznlBRR/x/wpeNRRjl803KOKMvezvIOJ41a+pL7Eo/EQeqi7S1UPs5L0AI9Xe8wG91pW
uEJRSphjYCXKt5SN++6uxdDcs+6KQa/7AN8kvompBmgMQlEKcA1gOvvIkdGYQtZ86hdUavTuDcCT
7AowwmbF0meTUrUZ1+z/3dNmHpGyOkZNMKaBj3YOnXqU/SjTjxQ4nRw/UMPpwfLMtN1V0naEM/sD
ltpg+ZW85BvNGzGSGmTySljH9OV02hXpuyrtG3UrsvJcCqnugwEMSUfy8abNkVM8mTTfCJt1p3dB
c99FgFsX16sS6ehqZiIS5DiBGep/1CAx4bgp00gAW2ptTj9WxiXqAnhqfHmeM3f8O5DMseZTbfno
Tdptdc3UGhm6RA65pazuTTnGXkm13XTgIQymNOV5dlGdzhtoIiybFgfZm8djPB6MGPC7mfmSgpwB
q87zA9bSBDBhgl8JZ62XKtuh9clBe/LPzXZtTXppTgT/HzUGIY2AqWOse4gdSHkM3RHmvJ3+8hDC
w24fbi1jjgazVmutLmTvr/GxiVNV3+rgZxkgf/GHyjR1cuR9K3nkdUCzdtE1MyIJP+3KSNuswMhj
6beNpSjGYHUfnAN/JcNDM32N9sLYNAuAzlHFZCNTqXQqHgt2Tx7N19AswU2bGGN8c2I8KmUYkQ1D
D3vHKlQm0VFLgkY4/pBE0Xu7ovhCQ56afEB1kj73P6I70+4DKS1ohUNDq2E3M+Pyo91dJJ0R12wi
ia3+YwATnNRtdXEu1wtWanwgbs15zh4EfV9Nx3uCEHmyVcj1D0ULed7rZBA51n3ZmYYaI0J7yZJT
qHRB6CfjgGtXWzIJlL3L3D8c0viK583SRBbnIyzUNIyNeZnQWNLvYSPYslLEkDCjj7bu4JwH0a2H
EwsWDf+gKq6idDtrhFgYouG1MxqAFvQeMeeJdSFtqNQX9tnMiMl2CuIu5mTQLonojI3luuflZd4v
7jsmiSRBquheHgrUzvkcmhQsZYfAzwxR7LQiptggJroHwKXVMG1GbwEZQEMRdeXeLOOz8gJ+Wsbb
O8HOP4SIWjYq0lfYbsxXgxfPYK1H+8MRYuhT8IN866ew5O15NdQAPpfXSFYs6i3fNh+s3pSSSQ28
BXQ2BThD7q53xi9P3OxjH0i/0avUgNw9af04Xek9k2zC27bViEvaoP4FgNXv8A1iat6BcIBeadtL
EV3G4fAegY8KzBtHbwIq9wACA6JDWl1OZps3sLm3qGcyNwv57d34mZCqB24vzlyXrJrdH+R7gL9W
Em4h4cCiA4bukFnqU/+kXtGSt0teHphl/q/XbzHYGVNZaiwfk1+Q9zUdCm1ApW01GVPkYSROJS+k
nQy7dPfll0gSzV3VbL/hmsnRiR0xG3wus4A1jw05tku7I7XS8FQtmoYv0QJz3Rb564aMQvS4349/
vB683NRRo5UnVL/AGxpamvMf0PoflGlM4fs74uu6QpbVCnGUBQb/05AgE0Wd+ZC93zdvCATGwZWm
abvph98H5I+yrRy2f9y/EY/rnvHA19lUGyMRFuHjwyc1Tvc3jtZn8udOrQQV+iRt0hoLu5qFBGJI
9sWMEzyN0fhvT+0uGA1b+FJATxTTkhBd4S/qBaZmNz82q1ltR2ZJCjXQaPdyqdxAnqYEQo4al+1Z
GkDkF7wPfOzlYxjTfsqpUxdWMVgjcZD9plRsndSlA3FpF1nI0TfKebspyhoEUfIJiBnGJhmJciZp
Eu1P3zyVqvaYfOptk7TnK2/RSZLgtSrUTYO20hGv73cOQ5NlASTjFW1RphthNAvkxEybIjryfUK1
htLq1+omDIgpPFc51PFXrkoALiCq5+Ivq8TkXQeIH5rzOqRpt4jv2A7Ixk6UXeO5rH9H1OI/JdsQ
K5MniD5x51KdAfMR91jMb69RU3TPkap01/uivuD7S2rjjy618zy5yuODSuJcUiJ7NIk/rxL4FvGx
5p7ta49TDgxjzm5P49sB3U/89ltd3LJoHsP7OTApbM/Yi+XdMb9GmQlkLLF/zE56NXCXog863rHF
D7BnqsScZNDb8wPhLqCJT5iek9iiWK1VuG9zv9fzdHrKDDQnWTu6YrAddd2LfiEYkwwxQTbgetSa
S334yqzo2sK5xnnfWTYzNzc2TpZMuMjBmpuTK9lxJJcTLz7/06y3/mLNXHH4CNZRkSzdlj4JLBny
K0YH1amfINud7abChGKz6zv5cZTJWDnJ1bcYogtcx71MkR7Pi+xlyum9KlKUr+lbb/TUaPpXnb29
8UMw723aMd9V9IXHi2zH2lOhko0DIr8ovL+r6/48Gajxzwof8lq8uB6jo0GvryUpUdsQsdU47Mf+
Aw8ouXLR6Pxa+f1vxceeyFOV2za9YZm/hqaDHHk/qs13iMPZHsHVHO/y6zleo57kDAmvX/UMor6P
zOajFgBIasvyp9tEHIGEb2p80i56wpt/o938F5sO7Z9qkMq50c69NWXoKu8H13y+qP+aG3acr2tk
uuhKlLbDysNFCj7FjpecZnIfXSiH55vHF+3LheHqmhGjtASI/oCuMlkuvcUJA4tm7P2Oo9d0JOui
37hPMsc+NefAhexYivcIizJN+/Xeob4q3FDwdL+lF56HPj37xY1NEmV7Lkgmb3A6zPTJmLMx4ZAu
4q/DQpWTip0kIinSU7FDzFQ1LVbWUXL7mwboCfLJf5EIcT0MCoG1Spayo7rP72gaO1GKFss/oYU4
/3VoWzXGmpdtn/RlxTOy0Cd1ryozGQKta9NKhoR6OvZuTbYnXW4UbWbiBWMDWXGGW0OWa7wPjQuW
O7JrUOgWdMzaMEVKYL3w1Rp+O0F4uUG1Zfb72Dz0AjCsYJLrXXBf/7hTFWgK1Tnvaar33w8/9GqN
0klcsbgBj2+j1TH0jY9O2V7qwJ0tIAJwzK1P7pZ52ujSeNEb/DjwuN4unzJHijg5mxG6lMr18/Cs
5dcZkLwtXykojCcQ4bNH9/XXVBA8YPqeFKJEyoipntvAuPEIOsxIXW/xtCQNh9gfoRkvO3N9yjvH
mZJ/Gc0rUmhEPHPDwsGdCXbeE0UlEMwMOmiFLXXB+yyjDYyn5NdV9O9EesZ/V24ic1OgSrBNFH7a
wvBxKqdA59+Se6wLbVq/plihECt740vjJdqFz0fl5BdB6l6/E5mZjVQiARv0iSlojZFo47G6pDXV
cxTJgyeG0aGqvuYh/EKQxY2djzFzVB7olXbTdUVG32Vv8uuSHpa/UYpkFJa1jqqeOuoNm/es3zxl
r1+q0KS8vIUOfokAjKhLIlT11HftqYSTioc8YCraOr2DmPLdhdbICHLFGqU09Dn0oAjO0AWph9kU
RwxZPTQ6dg/+m82cR6SDDhMQrDYcjsy053WEqgxVGc7PZQRT4cj35RRpRqKwI3eT7w1leaRaQyjK
k4FScox48lzb7DZ7oUKVd8hzRbe2E9a4csrrxL/tQcA7L1vrelUVq9RQSX45laQnpZYHfEGkcMxw
tYN39eIYIs78UJcyIm9eINJuZ92oCH2uEiAsmAOx7g2x+KhGrJByAkSUK2c6gKjg9Nf+/OTyJtKb
3Cfu4brfIS3i/PHDNfhQGardUxtW8Q5Kw2M88U3+8Zelzx5I3DNPhO8SO8YrD4ATIQVpQQs4OFvo
kRh/+olbE3KaHcaP0oVjaptMi0n0hOw7uGV6AHaDA1KzEGIjnziA4uarIIMxJ9QO+Yy4au+LhCwk
R2ymOqmC3mpcOPrtt74LkgNeWf9K9lbfoMCh4IaPrSjLfJGQXKtS0CnmnRRTnq3EV9tK0KwhwkqK
VY7RjJGaU5hxMyOMKA6Xu5kO+VAQpXfRyc7jerjOIlK8uhotNWLBobxan7cxgb366Eph+CQh3Q0V
BbAdtekpMvWeJkHAZjPgqVqIKODqYwZ0Po4HNCBR4YClBpPoymEAJdIuhf1trKZTKWKPexxVbiGt
rIYP0tU8ty/k70iYw877Dp4ifwSQP4x+jCkbHgKEi6MFq5GLQCnpNyWCn9pArxIuLFQZnu605kaj
iJ5fKMbufSaPqXeuUyT3WsIxbTD0XjPnXgBkuW1MTMft+wDXMZghqx1SD2vFN37RZG6T/5eyeF1y
JhPWVsPBWvpgjeIzK2CZYUHup9YPQjP7GrVzvARSu/utMSJFFzrYofp5JpzqsBc627YX/R3p9MIO
YCZEtCe+9Ht7MmKwkTRZykhxZjCUfDgbRxPBOaz5HpsL5TdewhquCo6NyMgO9ISdbLxl+j/yMmJr
vnJQkULqae6znIaFtS1OVJNZr0lg1N3rYNC4LEc8Z0pHO3WxTqvOm1cePK+zLxzDcBiK66HYZECU
h06z11blKQ4UGZpROfGRDu+EqEw1cKYnI9lfelzseVypqs9CqDouD0BPJIG48s8zSfQJknoEYSlL
L44Y5QwIX8CDEj9viMVCPV0BmUvGJs1ikVvNAUz3mnG7H4UV9UKvTwdEzR5RrdEHb9IDACwS7lfE
Mch1fYdV0moejtu54do3E1vB2+2DFAxfGyc5NLu//WXHYM4umaHc+yxYD2wzbOR7nnK38XIcfx4U
CpxarwBGVlMfBxJ4+2kNZrRKc+rCcwPLDtaARn9kC6OvRMT69yWR91B3fR776I71fi15SES+awT4
8mZJMAhs+8i0sQXfI1R/cWkTjLYtQ2S9VFvRo+5/tUsg3X5nbX2XBZ8glRbPzmoaeR4ER8SzL61w
jC7m08ok/cTsv9Qhr2SfLNBZMyrhUBEdUNzTki6a9SRmdQfyYFQezsbmyoz/BA1LvDPk9RAKJMtW
5p/Zu4iMSCVCfTFkWO/M+iJNyA3R6tzeiw9Eaklna+OjyyuMw0GLA1wy2IcylAYyyU/pf9dHeIOq
Zujv38JCdYbC7BTX8c2r6OjLKcMujXCpNKKgoRgK5cY/9LK3YCFIhq2ZBVR/Ur7Vk1g5PV7IzTTp
uSbLlDCKcEkHuU1zlxKcCO/WfvItqk+IKu5yPohLkUPhdIfuM6nEg3nIQj1i12mZW1f5JGwtXxOW
OvxlgmOnGVLZyHM66QMCIQsaSIiJNX3U4mbRjZVMCV9OggT0et2jlnYmGoCucXLllobnWLrKU2FA
VmCyQiZWkYaIwXeu8MhMsWPswkNKLFaGKgMjEJueoGeODIEXGexcDLq2ILngq0R6YTR2vjFEbNEn
+0e5L0apM2m0O5uM9LTtsC/LGnxBN24zeBiVbUIhoy7hwJ5s8mWF7YBT/JaNDFRFmNw4+s2tH/A/
oteVyFQmhCLdJ6PH0Sux29uJqLgiygZB2w/v+g0kTF2TdiisvB/5jQqh6+FM87ufY1w9RdIMNEkn
1AYRuMeGCYZt5iJ2TsQhDONbPrwlhGASLgK2Om5vAGnWka01dklFdQ29A2MQK8Qeo4/Zmx1K0l4p
G8jekUS07mRn0W0PZVXm9Vkb9/juUIQqRm6na4WO/IPdzKGHBuP4AHGyD+UttxqrzJtBBwNg513+
PjDHJsdeyCjjwTzBkGk06oSpgSS+1KsUTVRsyV0PCv852v9y0AGad4kuOXSf5dmL/XAlr2zMkEtA
MNylDDxjm7o/KSh0/hgNsXjWTNCowaDcj6hiP/KE/ppUveKWZ+DZTmCOFunQl03wPOABW4t5lPeK
IPyr5gagEPpfKfSF89XgIzrZkXEZ7kyXXPZX+QNlx4E8prcrkFxphzCD7473Ku28C+BhyLGwjk3f
7wzTCAjkq8m8dedNElev8oFI8KgOPsC5iemdA1SrIUpr9iXNY5Jtwg7kMUviQ9orxqR2kRPYOOLS
VZB+2W045nz/nULJPIFEj43u/Y9R1H9E3UiQg/a6QTJ24JI9rZLpJrHfvm/V7F3Ho5SGHYXXszEE
6l1LgeYISHxto7jmlCrPIarjEG1mUXJKsXfL/MKqFxsq5sLHt0Y5MXXgUMQFJ8LXonfa6uTHHAQW
i2bb9UWdqoo2Wo9jcsE5Y7v09WEqlmE7KEkc7Fr8PXs3J54aiUJnChOrPdX4eVbnxe/kUknh9mOw
PI0dyDS/nZ79cpsr1k4EhdAqXK8evP6jBxl+jtKuPgToChafeG1tQoF56l+jN7Fno2/OkkiifGpL
e/rkUk9/ymYXZ3l6Vkbnq+mHy8c0dteQYkGxoK4DbsDoTayZcsKsRivLBMyQBuciWUwV0IYQWiCh
etZcocWG65E7lDInM0vl5lU0Un3LlXHV/LSgsSKd/MU27QVa+Xv10ndyFldoHxK95MA6echOaEc1
UpPXzHgejgaKUShEu0fYCzSgRCsK+zTLIAJJHCLUh68CZ777fmNRSMiN6MY+uTqp3orNcY6WjJLz
pMX/gphNM2YEUl5yNuYewp+hiWXueh08s7Uz9Pix4/XxWf6Bh2cauOw5kIkxaCLOksoDlqNzvhzt
tYl8J8G3EkIwoObe+x023deyrMCKkVxFte2MyVtSUjHYjHRBtmn5Q3fdTQaX+I6wPdIpXEzqXwhH
eoKR1W+PItMqn/iKw2zgtppRA6PpnN3RvLK23GAg4jepogn47DP74z7lgHR+X4kZEO4EXKNou/3n
iF9T/U/jp9TULJwa4kgjSYsrKNWCRDzDKamaar/2VJ50Mix+X6AKtcDN5EZYpOJyBlYR7TwKc45f
ktxA9JJ4qVcNohpvyHxbhx01Vr0e6NTsJYMJ/5kp9S7IQLSAdJqZpPXqaLOd8upiCdjbWk38Fk8K
9x4xN+KHSJ6UZT6HLZdgR5jX//TPGsOrCTBJTxUSUT0I5eH1unw0civzGPPWbDxcqWMJUcgrp4UE
naGcGGVdW7MTxC9YfTCA7C/k0QY/U3WLOFTqMMlnOU4BJb190lUS9b5pu89AFBo5sK7blGs1p5jQ
DKKZAS/KqnqxISY7oVp4B9I+e1uh1aF4Z3NhYE6D0bOD8BxkbBk6hXO9wR/ohKtKPjMzOGTQHPHw
xFKh4vjxngfytw71S5iRM5qYPBKEukTI38udwu863K2yyE+kN2nbcYkIStBRjXw0vEP/Kbhjlt3M
0nO68Hrn1S3Tp/uwtPWOpjXrcIuz7muthE6ZgDyk0t7cCM/IAl1SV4fWJ9dlkWrguEbHkIbmlave
zZB+f//+Qmvgb0x8Bp5MLS+1Kny+kz1iDN7aGYm/C2v31DuVbI4APiS78zfVb2F483m0wWsa3z6x
+9ZUhaE4prxTrG6P01Wew6BdtZrXyUppR4K7e1H5cBjBs6QnexE8XDz4C344HqDG8SPKM7waLLLP
MGwvffCIrL3AmPiCa7/ZjyF3KWn20k1AZ5xCTxFS4qoScG9aPtzavG8alsa8ECIL2oJS8ni63bBp
ynRkZXfI65COSJj+IDtvDXq6IkawC5j2FvCoD7XPf1utsI7FNSQWqgpQ6I2MRVGsHOpowe1n2QC+
XdN8pwSpOodDk927ppYNWsaNOsdg+p7wWY8zn6j8IpuRUvRlCiZu2d0/MbxGPlqUpL5HgORacDU3
paPZweCHEk4tgXTy+v6a5j+4r8FtXebC1Zxd/bwOL/O1Cq8mPiuiCtPUPnuFI5hVsUeggNxvKARe
WKeqDoWRNUplZKva20rGZHuB5kGazBAAYoSnXoZssxCLR6qCLZ32K9zVTDqkj6kEBVz15D2N0KmX
Lx83wBqHnbN0UTZhWiNHxo8W1CXwCHGtvNnafxP5enPvKiPoOiLgWxLqC/2FK/Ji1ty72DSZcs6l
3BdrHYTkqZ4yWt+vHe8pNEJhZZXXrv9cIb2kA6ziK5RB4OHEZsZ5LVy2y+2YKiofStyzQfHUVyL9
NZX3zswQCea5K+Tr49wzuM1fk57SCScqQ3yXuQEBYlAjVjt/9kIT1phASgXhyjki7Ry90q4XOQrk
qTnbI0bsQLdnLEojPMaXrbdXWuRqorqdRHemuduEOY3ibeyqyIHuFlol+xuWq5X/8pTvKtMg2U3V
EIyiXn7YVNJRZuIJ+INFdbM+OH6IMTXTAGY+UVX88vrkKaxa1RDQFqEHx+4y5eBJNcrnSV/2tiOx
uS5pab+HPte5XwtRMCnzmK9RIiAAMTuwgyE4Ad9TxYxgtq4g4nJ6Ynyg7LWBxNJnIqNqYETeSAqe
wywWRBKApe5rnZYAGk84v7cRDi5b4cGI2456BzTjOIXoXv6Jw27ikDxBO+H49N5tuZkpRVXM/I8Y
ddCbvCL2N0SG0LcnDmpNJ9Ma53SPcPjZnQklOiUyouS5zLl9NK/k1yqNA6Lo8wAEu0+YSzSSDojt
mytHF9/N/j0taYHW4LJSzAmDMwa77/f75Slp54G4s8EXjrLoIugqXPDZuH/fiF+YCJEGOiA/zRgT
4lisvjH/lxCqsrhiOLJ3R/MdQ2602Qib0uFHWOSalf5Ld8gHxqx0dGwke9eZ/3KVP2USKZUb0qxW
brB166zE14rhCnprwea5sjWitKqu30Bx0qX8IRqaCSOMKVKsYmCSv8gUqEb5fIkT1MkWbEEr2TDD
uqtypGMh4HMZkpHSfPUGDbBA6smFVbGILR+MRlrIBTI9l0+PX6mpMZIQ3H98sZBwNvK+P1H4dxrx
hcVPuOBIO+GfyIUqPMYmGzK36rBwkNQQjLRwq8/Y+jhL+a1uHueZWwxKpCL/b2PbcEgAA3Kgfmpy
wzpNjix1kBczuA6U2NO+6a7LZEN+j/UnQ+HcA9oR1r7nI7ii8PSlqHdomHUUGYa7tHjXD0gxQKu3
tmA0eVlVoB1fTUD3d3Ay3ghBRQEGaRfCOcIfF1/5kH+hZIAAF4hUv79TKkCUIhV7C6ufRI1tmncf
eqohCoUaiZPGLvayeZifdiXsoShSNojm9uj+Q+5hKM5x6RdiXdeYEsEJwgQIor0WUvE4QkGH/wdr
aCb+j1G/hUHQ9/IueH8e3zHc7zjhMoB2PIygzrB09qFxxkvUd7AVY78XvFairKj/vI0TZQwm/aTS
GtB1jVlogfBpBmZttkfbz0CANihhqZeGc8ZcViHdnb4jwBkyeH5NCf/ljQrgryTHMA3nIuaIGM98
xnJ0AIv756c8tl1pPW8zbdR0VNI/5xrYizC7RK8RlVq/T0RCDibSBHCyTVOzOfirK0oAwQkQEzm6
BErjg0fGap+uLfSvFWE5/DyLafypZYAjV9NjfCRbQQUSHR9kMMzLBsSnHwBVjwusX/Xp2rFFbCBI
K3dRsfa7nB4H9C+g67sXAAttz3Ht/cixvyIVoxCaqQuDph2OexytNlKhHReXW8XUbZ/h2mtZIrDQ
xePLwkc5jpNXZfi2fP+xHQYtaC9IotN31g/uea5ppB8OoEA8Q0XnHUrVlwMwRpM27V5xxxZxRNYV
BsOzfGrLPYlEcrZB2IQw5S1XpJs+INVqvlJGvkY3NuZDtJZicltR3tQZSRCdycVE8dGEePqoXAUA
mXO9GAVwC/aYtaSpuddZj1a1BjyIZ7pSmBws+8V0tfsalx0xOC3MGYFhODHXttOn9Dj7egDopTWi
+8F8iYy507batiA4/zaV37IHsIj8NC0We/2IGzRtEy6xeMr2Hcb0JpNkCAJrVJN2XQKXOMpwd4Sv
xE8gLsQMcjkx6rCDwh3K8Pa5wUnwLY33+UY1Nzh7lqj5UmwZWlldcgoqkQyt/3+LvrxXPqksIrbN
JhDNFvHz8MBozM+C4TWBfPZoJfHqGl2mY9SmnP4pH3yzdUj1Hjvd21Wo98J+oyyEp54w4FJM/kTH
q4R70C2LKCruhfPNPeIdZdFN/5Zhb2FIW0M/fIlbXCfIdneD6GWF0I6aDW3qjjXvFmEtWyYPm58b
lQhU/omZJOAbIe5mk6unDKrt4C/3bOqJp1XcaT2po7tj0c/6RPr+gWA8eNyBsS1wp5Tjn9FTHhze
zGJzTA6e5N0dXSsrE/nTGA4fGha3Z48/9ELd2Ro/eqWAm9Oe2b/9ZV/BxUaLi/EZ5r9XLhMJXDA9
v1cNr/Tezs4578m5hMuEdcAcLw/P/bCNSeTs2zLgcoRGDaHPWAZ6EDXukILBWNtHxJNloq9A2sPN
+WJJ/1jJyXA+oZ0+kZWKzdqTlWqqS8vMiwo3Ce3pBqNBmmNECtX0yQ3gtKd/8n9J4FNlMTob2N+F
l4wuzjpQp2Bp24ByOTyGaWSYBpcYE7aqO9CFtsAcjz5idu0KYzqLRalIXxQpOldT4S9q8IKQ7Tbp
Wkn+/Uwgb69vyrqQTemNsoQX744e8JsGhtgzG9Hskt8xwBbEKpYFywxJVIVfb5vV1m+mkM0+RCx0
Pqyltop5wlMp0XP4cXeXCjfzKHd8qaF5AujWzgjjgYTJbhSGP1agxHPLajqJxlO+Ay0vJU9olj+N
38HnkOQ+WwYPuKDR8nH4SJV/fPDQRa1aaPRqx6kGZOB5e/3nkDiNXjmyXj2MPOLJGOFy9m6qAt/j
R6fZIxgRkCwcHkPRh0L/0aXP1XYplrMEz+9aflezDm2XX3fcd3aSqxDzMdFiuQw4c7r7jc0De/4r
HNlOOQnoSV3BVBtT0ehUczybw3WgNHiJB7zqtkEaQv7MUgBqM/TUABtLD3ZrilaRZZBAALQapJhZ
3UTgyg6lknH111Hngcv5HkDD1vQbIjJaXC1TMYY13OVT/TuIrTlJ36niP5aDnu+Xoj15nEUOJMwh
RfQBLiD9XnDDQ4JXvlyC/rw2sL3vhaGvvfUjVvI4BRbCoUnMDbDxTs6L+Bi0okLRzsmgixuyjAy/
03bkyHy6mKdBQ/7GSUgi11jvFhwkhx4c+/rKedzAkkMblphXWT8BfrmX31w/zOX4KjSoHablmZ1f
HJ5CkIH2cek7atc++zVr4/peNgHAnsZVfb9HHVZw7KxalAba8IUwaWPLIXYK3gzvduCcuBhwJQZ9
OXSKgZKGBH6KdX3ex0Nc7wCFqKCmI5XSXlgYghgaHrbUKASG8BAHG9XplOF/r9UeoZ7x9bSekQAK
UPot0bTFaRAbfTiJ3mXK+Rg5w8LlmafrxtmVXW1CwJqf0g6jRrCKihvub7Nj48bELEFuMUvIzaf7
L7Tvu0p5CMY4Zca2Y5Z8Q6HhLgAC6Xq4Y+vWk6oHsycvr4aTqHxYkqbKhBng/e32e2iD/F7Md9Cu
du2nGYmderu3EUdnrrMXi1c3CsIj8LEvuvHF5zmdwJ6Q/UiFIFFB+0FYWyRlEuDt3CMJ7OQbux1O
9ie3HTyJHvPYcux+j1NCdlAEFDrdCUmk4Xj6jjF+hr0euqgKOSF1doe/bASG707IRKaYMQ5+SLYE
anRdPmXrPDw5+TgcN4L6enl+fmfjwcW7YUXxpbzeZyooymFSk5G0jZZL88ToyxAmIjv61lXw819R
dAFt4IH5oZesVSpKCP40Rg+iCXngI20+1GXNsgU/74nKRZt59qvMw7W1e1aIqEvjUDjeqcImRSOW
mxCnAxaF2xNYKnImp0KPCqDVNPwe6mCEI7TnPcv+3aktNToTLmmbi1bBGL+sOT6HxP9dmXpPrGQX
CISd12Zi/zz9xb3HAztRhekUbJ0Troy5XjO0tvguaPogy+eg4hV60Umpi++tuCIigZPN5JZpA6pf
S7rHVaStpHIJq1roQ8JRJAKgWCBKB7Mfj50dN/8B+vomE/9jqwFEHe/ZukyysoKlXxEHhaX/z1sL
Xzl1zoftNtL/YS+3OYUtQ0Vue/9x/ehUosRB8kXPFqdRkvzo9BEyUH+WFejHP4kJ2lCyOaksrUPc
7f8WdH2RcdRRiJzrocucXKcZydSukJCi69zag9OvEtAeJurfBbWmxGJMQWnoA5M5kxVc0wETBQnr
zmbLz/vJz4gtOxi4Z2tqjGo/7mBMEmxTM63AS5ZWkWbm1knvjhCq6Rh3KNKPWbDfq6rApX7gi0fC
BkPaDzTXfXKr06anjTDzNLaG72FcmO3qnLf48Kf6H3+qbv+MN8ViPp/8selHjiJouIIcX+K2hFZK
Fw1/ZKXELImGskrqYvywgWJKqHNmH7UZO7L263VubAjgqBEba2cDYOKALAkzHnKHRGo/SkGhKMom
LENQoXMrPSaYpVIvPUekIRZIBjbyOKLYvkq1fApb/XLpm7RxkIBSzRdYe1cDAGkWhF1lPGmigReH
3ORzOtrTk0Wdle+cVQi4DWUGA3iKw13ONmiXvk3ghKDg1zpu06yO2TjxY524FS/lkC2wm7Ws8Ecc
J08muGSozs6lNfmi4/kh5NEXjsO73QEE31+A69Vf1psyFwaSZY1sTTFCB0WE2hO0H3zT2Ii7+NJ1
JAc5e4vgaykP2N6zKHIG7rPsBdcnS9L1pBZafH0b3ZcU9+Zg2f/QR0XAPPL5j11aJugwIbx2Joib
c0+A/ioxWO9kPFi/kbd49xVzYvhyxMkaJTxUSY40puMr9Esib3Vi1R8IVJU+u1UJCxglAHwibvng
bq/KpOtp1G3jmflTxdEQdFFeT4NsEt6P+8VojOiibfO1Oo2DcFu0JIVPDb2YxHk2yQ4iGEigugCz
0OOb876KItJkosjj4qbiQmLLHap6PiPDicJqzya5VKPcX07xaG0CPA90ti+YB9oXEgIWLY1+zUgW
h9oR5xDiEKrmIjQj0rtjq4Wp8ju+iG4g5cmv/6FF3m+0xlel9FpK3D9g+xxCkM/xRxBUS7gA6f6e
UO9RsSFhpyEGVKW3dt0h2yyvNRB+ZZcrgpC/d9nUDFfuLYOXgoFhjW+t1zAVhBxzU7jmMeYsXg4e
aEsV/fIBIDTAGMCuUQ16lB4+Z9J2e6vhaTfgkR2q+u1TRKfwiyQav7k2PFOaNpXqfyFFQ9GJh8L6
xRWFM+dfIhCiB5tsS57nG3l60CPhcT8MI3UVVTixMy7cvIqYvjRx0AAXHOSHF1AB6ofkrpLOn4wZ
2gJp+XRn04uTz1WH3z7+tLgxIKFq42ApR2u5ViBreWUwnKWsbrnu1h2x1yFmml1yLMcuUiGFz/UV
EjhcBFzyyyzjkRGI4loFthYS19pJewYYiYv0wTkZEAcb0J3iQ4gD0KkTrBxXWFIW990LY4AsPB0n
mR7bzPgqC1tgbZOtUZTbWZ372OOxAqLKS5hEns95lrxIw3UV4OHgns2CbmE7X/wc6mZsxeIZX7ZC
yfdk8q24N8GKk1Q0Jr0WjvKkjvZonwBlcMBoK9JRthVotLcIC0FQ8F1RjLG0m+fBV9P65ntyrAeZ
oRMZ9/ni+03mxotZqbifPaaRTJE5Op+BFqOVPHVXRFsZWjzx9CL+e/HXJdZVig2iMOydMjXuQdiW
cZBXhAL31lsX3L+LOQVL98Uw1mod+sBpcZgtoCBwua8/YrgioIxVhNGMePmwnerx3PkubhtIhyaP
ncpNngWR25AxD/0ytQrDXgMIjq038qzl8rhs2mDd458SmNvyn4EyCWPMpOMfPuf/fTv7wgSvi3fD
SeQyuvzYmmxZn1BxHkvQHU9LEeEyxwkYpdVUqp54DrePsy69PlQTUzgQlEgO212EMn9Bn9ZyW9JI
YJP4ZT96WdWmYexaIaKZ9VUELwTt1bO0wqXDN4MUn3yxvXGMvk8LzVaGcAP5Q5AwWNU78rSrOTck
lY65tohnLcCxqveZ4zGFnrz8Y3l6HCaTJxgts8iL5ntLvCWkhpIrOAYhsz8ENS4l+/QylkKAqPhc
b/Jy6AWG7NtJGdAWy23dlTxj6JuITXV4oWeP4yTgU1Jp0u4yUTysTHiGfGXTKhnFc+H8Lw+rwdfy
BE8LAih20hFCQCOSgZPqVrm7p/GdCBcsi+SCTtA4yz0wXDBM7cycdWSOFM4Ra1ZKyzCOV1DMeP+o
oSwjVUDZafByMSmaJ9H2tTEOrU7E4+N2kTowYa4VwwCusNPvshio+gNww3Hcyu76RgA50fNgvW2F
5ua0w2s1ZJNTFTKSEEun556E1kUQDoF+nE2VDlwC/KJ2roIR0yHEra6UBpqPPLp1Mqog+a8MBIma
4BVsbZWiq/CiDCZALYW8MEu5JmTw5UUN9tGD3GPhhmKCvC25e5o0toGoPeJUsOFTzO/6QVGWIPHz
4ucTYIsvrdqrUczNs/WVMgopkNxqoRc4HmbnVKYJuBWkQJ6vaSFk7wtrJhfVtnMF8EKUhxLQlY5J
ujmywR/HvuS73Dnq5eNjTg7Ras11MI+AkavhpnyxrhCwN0NCp4fHOYT28LpkLA2cqGtO9joCiRSA
igpO6LrehmyZXLznk4SlfBqR8SOo0Z7fghQ9+C9013u+cqp6e/Re0GBufGuayX3jMJ2Ob1TAWWw2
81478y9puVxsZVWIdLdpohg7tNl+LrV9nClLuBD2ljhWcpC2MN/1EcbTYCLYvlsdVLq8pdV4f3n3
KzIkEc85UQFeC9BGuuZC7LH1rMUVpC6EYD61+Ztb2kQwxQ9QwLhBGUOXOARe49ogZmzYBSDxVZ7u
2ixhLyfH0TUljHMgmzKamp4fDitPOWxehzzcAbKBwag0eYry+GCPrZJJyMU5iFqbesK72QHb/I7m
QTNXQhhRkT+U9KUMTXa6ZgV8+fBFmSaNRK/BG1mL3cVhZHK/2NchneqRoV1Y2T5VWKJLbUHN6EGk
rzYhP6xLz2hTx/nVkP6tga7ag6u5GlVswi8JcXqaMYJGGNIVk+5JRYk4xK3lvEh0mCSeT2/wtB1w
Gr2yTGVbUPI1Cbk2agMl/M/GmsCl+EyoeeXWGwTFhffsheCt0MfiPwgo0j6CSmaHHAgxno3kOD4m
gDg8VLfYQZ/jhkVE1fQpTxXvVRKxqYRDl6FO8MheiKXdZhqrepBJYKp+UC2piE14N6WozYzpU0Dx
JLoho82ty/mYxXT2hOB+e3Li03+Cp4fzNEkVN4/bPCWSpOCSdkhXqX2ZsTh4XgbJiBMbWjqpYYo6
dhO+M7BFNu/7RaY3QdYpev+gA30CSevUMNKOe/cqziyQIB5UgEeJHYFIIkk15gYTxodCeUAIFLrK
D+H/2avvIn12EUsOlaSq0d86lu5vc2qD5odwG8Br0ffE920PCAsCAWKr7RgrCnCdXQ0Bk2qacfC8
j2vXSzrERdqcl41GVLxMBUzhiY0NQyDohvP5jjqjxFxXiqHG7zbs42MQNZah5QvMFm7Re1ogwngI
EI8VaaYKdz0mpknbB91bhapH5ZVavDhE9A2XyGoPerRsrB63vMORDI1wul9v9VAKGQx3P7FPZX2D
pIQAN3qAjT0VxN92SxMVdzYlCr0BIpdTiNbXEYBNlQK2OTeehV96mv/jPyaZKg3Rz68Hsrbb/B2J
UuBwjjHI2o4Pv5UJZph5hmfQTOlLZarnCi0LKh8bxc1s7X1I8BBAxQosraFJtWUzpEaeDZtHgaH2
IaY2p4uCbG1tetNOg5jEM6HrYOfbTrR1Vpo/Dyu7osvUqkAnYu+bKPCLI9RHqJDsIDa1PVdGj131
NixvPLwRa6XWi3xEPGQ48kXx4twOBkD1g+ZKymbP4A9D/OdAC+T1wZrXJ3viXERbgwctIkIvD+Ta
Cqxp8mpiMeifHsgONG3lMMi51FTtV1hXMIGSvRBuHs10MN9ov3/v4JJJh1JfrKXOoFmbV238Kzct
ngkRo3I3f1w+5Er3Pl2l73E9WDTrwdVdn1zJscdACJMt+KAA7NXV6QXyeKQN4RSy2XuuebSqsxRx
a+2didtTOygkMYdl6TKSvmN7bU+YGmniUfHuOfoP8xoUAyWFGobxhWMB6K2YiuqdrOnFUnOV2F1L
FU69yz/BKkHFAomMs1RhEgtaUuIqa5Z8J5nAxrzYqyGfhMomjSba34dtcI5TL26xKdRzAfSrHreI
ylrK8VXMdpsCTXfKECcaTBlEW3l/SRzd0PtBnJ8LAqLhmB2Pj0+uZWi3f/ENd3stHNf8xyKSgXif
lT0PzTq/gwf/Za6X93vuivNYAnMYbm92fj5qvzPHBoyp5k15p+0SGXaqTudjnQQcdae7B7wmFjTZ
EgS8NRdoTY1YfKdU7X9NR+67OyqSkXH5SpzkZFjRCcNmxE4GXMGm8UZXYyRUlb66eeHLsZ0RYNa6
lrLtxlG5zwscGQibUBZd4zhDmuYSQoyY1Ni2FX16OnIN6GUUSRBA49FSjafacO/RZ1MIU0BkONBh
XOVfQ3U076EfX7blqggMpsDVe313n0HbxtKSJj8e3aw0tTTCX/EnuQq1LRQkOT6LsJ6Udh/06DsI
dVDJM6ouu/cxoQvfN3UdtOPa++FPzpyh1wXUJHtWiVuSJKFm3YVzFYoUBEfOdurCa+k84vRBVQ8Q
jCce08E2Zvaz+r6McNIjDMlLQDpM7YZMbPhhbbzObKrbthsL0xfoiBkaycUGVDHKk8olDqIO0RI0
0yoa4z+0y7gOXOmZQ3KqmThwq2G+WgiUlNIvL/RNYF8RMk3wY7o2AKIFEq3uHSrPs5R2yWHK2/db
7wQ5LebWsN2jr4x40tK5BAQE9fDT176Npoo8kF3S7MbhJtAcnmyibvdNdHfGBIgu6uldrdd0+fcj
BwMs57J86vyVsD59vowmZVWQPRTMaYibxXTRN7olVllX0Go2PlBnLDa5wD0UpnD2osMiMZafRi3p
mpzDvCEDkbE2SE+II1buF0TCLnm3JL9d4iJz0TkbLPPgYow5cVQ0LScv1LOWVPlnEvu2aYmW+7rZ
9glk6FPeagJ5lZDHbG4wYpqof2pAA5MY8o+HSPRtUvE5w3+n9hEd82CMOjVnIZ1g0eyRf87Q2N4V
wXGMVRbneAW/YxQ5y1Ie7EojyX1vaJrDgxCoqo27MCgsoryNm/PFJ0PAGHQTju2+K+AkZJuuwnmk
oeGWaMR+F9Fgs7glSf66+1YqUF+8g63D3VSVo9LQXAnUYy1rp0OduvcZH2K5QiS61CtynFg8ayvd
RQVDjk9iEVtuLzgfX0AVWDRBBrcssuxR1Q0KnZsWRwNvAdoYEW2hbiPcz+OKVpR5Je+VKtPKTCkS
jaox79McnTL2JLC8Axc93mQ5SriDjzgiLcssepa5Cg3hzX399oYVPWqDT7a6aGw/MTSsbVWLu3mT
ceutRswotvZ6R1BGxoqSkZJRBVmDQ46SqVNOOD/APDIZohHxUzts2FRqRYdSK9nrrhBjci7EDt7X
FvBKs96iDldmI7IQFNnhiXC+BWm3Z5yk9ZZ1S4uMl91AACz9ayWMMLA5gmeqKy00Uj4i92gAokG7
bawhxsBCdOOym6m3yl68nhmIjH6ht+75hTRwtYhrvmOSJjptOdAgbApzUEnWP6jlWUqm9PLP8fOt
qWNnZ+hKDqdZDzvvNmQ3YkhF9P9gDjIJQVXncESLvxgTBO7Ev59M/DXRNzmP6sG3hhws9y8j2gqk
jzOUz9vlHzg+UscEL5TjcE9NHWajKqhCTAxzcDmU0/Bh5WI+kMbdGCVt4kmXsH/oxVts4UgrEITH
bcC/OFs9tEfl4UQ5gtkk+ivI//pGd0NjXRreDuczi3NiS+nTdygq548cr8Iotzmrtkv2+Us4mKou
TpFybUpZAm2fCVFz2ZvFgAfECWhI+MEakQYzY3dqBn3hVdQzLWkHALpxRbIYtuEA8yFBTdog/K4S
9GH3l5mUokkFY+w58VcycWxShkJtwOeWGo5m8wi9TfuziKeqaug98UV5gTmespKK0wEZohDciDDb
QcWQLiVnCgvbYu1Pnr9AOpezaDU8Qcwj+P1oqkIlSSTfzsv2lH2qvuwmyA7A0mtGj0pVVl/7ty8k
m489bi1dVi+HWPHfettZYf1Oc6P2o70h9EsoLdMX7ztH+xkyxKpsLcfy3IfzvXGqrNdKUOO2CcaY
A0JsxrMXTr7sEu1xTWbxHzlCXloQaKjYeOIA5BU9W4Azb9GwOBygHMm6cYy5NgR4Cjumt3RBDwJN
a1nLitSCPgTq9y3FHpU5MHjI+FIKbvi5RQ67q1AeL+nhh1zSOYeNsIuvof8hg2IE8BLmejsk3r8w
YOGNqghba3wJDF7zp1guNDKbkctKNOILvYu5/J6Huo6thW5GHG3zo+A0AXtmk0jn0PbcTPsD5dTF
OoGGyjQzyswp6URbO7a2a+GeGFf+8B6YFf8OZBLD92fh6tOeJiidHlSf8yOsg22k31qhHSuRx+W+
HoeS/KfqG9/cX7dIDWRgRfppBTF6mq04GYg3tvLtlgFmQciHbilC0alNoJHXTkjq9ZwoSnHGG53D
aubqe7Rs74tazwDyG7fSh+GRk0kaZFhgPcKnQ3hZRQRpsMHavkmRT6Y2ycopS0h+Xv5IPCF5C+Ao
KKOZvQ9J1aE6wpwBE/YObLVHu3mSvLVkmX7wZC2KUFnSscJ4VpfaAngT9KFgqYm4qvmHacoZ3cEp
boMZK9KoHyFsQ/ZE2VJHToQG9npXHx9PZzA5svAnC5gUdPpU0Y33LP/2ZmZ8Q7Qf2OWZANgW/Jdv
gXwyyXRMOg7FL85kTAp89lBTAb+hKCPEZNnAV159W5unu3Y89+jN9TzoCpHALy5e3eyNpC1tohqn
gdRv/b9t9noLP99In7vhhUZwKSA+V7jR+O3fvEOaKUsGhCwglFSMRuI0OhV++vhX9PlUSVBw4jAX
dqVveVrxCWMRSF+yz+5Aj1KHha1B2ke8+fw3uKK8ef9WTPJJxwe2VPyObR5ZSm8BZ8oE8aAhw/q1
+KVsuCmz9ybym+r6t8gUG9MUEn8M66CzJcYUklH8MM191/C1keFN+kpngxqPJO6DICaN+Mghwkwy
2rC1/ZWdEDe/bsSu2FoURu4uiGgq12t73pwKDxa2hOtis+duvEnXSCy7Hakdc4nZvWfPRc4JbO28
9EoEKGGS55TjvvL4JJ7mhtlGfaUSsleOqc3t73nNoVVDObZCOkY518eDAuauB+qFZTy3um6gKjFT
1B4xf+GSkoQtVTTga7c+Mr62LqflmQaXp+zJnYDYB5fySnZI8xbGG9h2kXeqb+RbV9twV1wGi6Yv
bfTEjRMjQ2Rpi1N7e7gqwfHIr2I7pjVQm8lWMJeuwXWCRcZUV+RkfzPZayYi28qM6aA2vO++zvqQ
CA+wEDYHzqXrWedActAtV/suOkpbRpgGreJrJ48Z/3OwgDUxyRQOF0KrY+Zdkqaifaav2pcTt1oP
Eln/FvruLecabTSQpyXuwAOHtG2AQG3eqzcvMB1EVCCjAGpMTbSEjneKcpt+CkESbzm0moRKvunc
m2RKrU2eC6uYpuBz76ekGPswmQjphxcwKBBqXc+4xm9IGaHKFrC03Vq0QixKtaHGgvxSPFCyCSFT
cnmonoTjPGqRjF0FQ3Xvn7T1a+RJstek8mABoNz0FU/LQ3uBBERA+CiUtWXc9UC/HqUVkQxRURb/
A4xO+A85TMy/EKokD4rPnhnp9rX/Ytad0ENEcCUlmVptoPednCNRai69HzAe1dxFv7T7KhmEwePy
quIwnBpq3kwqJjYjbKTqkfeFQeqO4aZefjEpJ0loi2UeMg+34fU6GgyrtYnydUIE6o6LwDPiSA0l
Tj7EkcydNAeLu1Juuddg9QEoaII19iDVehjyW8gbclPv+2Ip986FvJg2I3WsX/kcteY/O4upVE4Y
n77P8+PcZM2kePPp+l4T3lAmLhah2tcBFjkG+rvoTP6/Lc30UBppuPFmgiTYFWRSePaM8Fslfuew
NgsOZhF4ITwKUHRLb2935jFn9+9oiUEw58QHfqj49Mvh9DBkyX7dldRlvkwhBiz7D2qj6T5bYtTC
+y1jg23e4JoAjq9YfviIOtkoHjFsXMEjNjL+ouop5Kv07UKRkfzVOADO8W7Lq6adFbLX5HHdXjR2
xilG/hd3WPLbE2LLE4NwzLoQZ58fvz+uMRsw4UOh3MhBh510ZLN6OLFi5BO1SEHdRVBNRJdzTyfK
5MeT6JxQtcv030kcPWFoQBVX6hrG53LnKo4eWQdwMyb+/k6IQUc2MNcLY+CbvTp6CQtvXzFWEA4f
394JdJRN99Jek5YCmMHBpvq2ivmHHQfgpFHwKE2jtZTwnoEDXyleg07sODdP1HKRVJ1ERvOLXfN9
1i3KnFMnxgoE9y1Dy4eZSTcpbKC2ckVTQRd0vwNUvulZapUNd4JNC+LMRZOolRAD1OzjEZTY4dIN
LMIHYxPnm3ZDP1GOf0j6QzoKQ1dkpLAQb33Per4u7JCeHH/gsBjElzWZGTXFxWmL4X3+Yz8hku5H
pukns7bdLgE4r3J8Q5PPu8TQZAbsHAZN1I6DHJ6TyyHAonXH8yTc1MDcrvJWO0McrXcAXhreR8pY
yKdlkn6gH5yWbHDQJ7fR3WPfpEDwC8PDlvtQl0vEaJ/0AX3/lr//L3TuVBYiblsO1BzjIsHqlfOb
cBUX3OEKEC1dkgrVZPhrPK/fOF4aalV0WLsHybZ7WPEucvf8cnODNhUZYqfxCFyaVKTodrNw3mjk
LW1lRAXfjUkmDn9gHuDjP582Bei7NIg3gIA4F5dsOy4RVRcZA657rhntVijf50pmoYV3HBxK6i0H
Mx+qrlsRZnO5d+lqirTMra5Wr7ARkFqpEcoQGz/N19X0+yZI4PluP2sAD0TbuPzANKJ0iYYsgj4C
L3tkssn9tOnV0tC41Ytb2CU7PSjlTm0rOys7s+yoKRH1QJAt0+ZY/ihRYddcCWlYMWvreFmataPI
gI0zslzcivF70Y045P4Z9FbJV6FTvJApqz8WgxosIY5VPwl+2N2AYSBFrSR8nqpxXCR51/oO/l0C
FsjWjcpGpOHeqOnxgQFf7ApVzg0G36QylY6pNu26MmslQi/sTdosoQVWCePGqzSf80hlebcZ9tYP
1uvFodMddCCV1qPlZDidzuugOM5NDIiX38v6aStk3d1n2yoF0qxu7ZS3m+nOckXeJ46Jw3+wbIcs
Ezfo9SvBv5v4Rz8d/ldDkjA4rTOeAukJvjFLDHMBfm9XXUhu6pPFDNFilIoICXfdTdyA+kcJBx2M
c6rdTpWxEuGC/dYieCr93lQHthP66GATJgBBhhss4ymceUofA75tUYV19iOKnygCesU3x/2SfHWk
n7TJGmEe7HHrOK+J+Rv2mn8BKvGexP2kmifI+OL4dQN/u5B2J+OE3wiCJrUN0vwY9nBYam/t2JYq
eemK469JD9yxRPjE34ZhFDenn1Qk3FY+xYwgxmz+l5YGpAAOwxvJbMytKmEr7b/A0f5b4qDtcdYU
IfCXcXjYivsNVaOM0AL5Yplvsr5hxcTYvGZ0jsw4XC4CdP+JSFOwnJqWHJMjSBB1udq8gO8wR42P
PcGyoDCMWDPaIpLBq15I09Cjy6GfG49ICuLbiiGBmf4WwkaOwHm8F6dxP9CqstjbWsMGEO7xgO2Z
CtEWxYvc7YSok3X5EbqBmnuCLX3rf2KoLOZfOZxuDpIOU7LAROAxCnGV/GD+BmQe0GwG+ZBt7nmt
cK3+lZp8dnZfQUL2N4UBq5kqHL/G7iGzv6azm7A1FlfjkUzhkDy5Mf108pBJ7NEbU5cTJS+3IMd8
wf9aUb9Aj8PQqfjeO1siyoQ/rvtHELqxs8dirYsMkf9Zf+t/LyOCU/mcSmUV7Cbs/Xb+QMzlSgBY
wxkZcsS7Ggoou8PeQqerq6wznKikDbr5mBHiKoFRWgUh3Wbh1xh/uV5bvrd2CSoyxh0FW1lRoa+G
58EUK8HNFtyH2HXnUS1C/xb4Uwpe1EAnNkt4s2WEnmuZLtAkxs7+Ht8NhiPmQBzt5H6RNBpNzd4d
9/DQlxUSUuH+m19kK/KOMPL0xGC/AwKPDUXVWyln+oOcGy8FaAsieVE2Bcggy5tOgPe3u64nTMhC
UFpb1sZgevmiiqRM6zo42w1Yt0hyBbkoX4cjaEwNU84ZNrMyy9rBDnaEHN4anVOer5XI8a1KVQAL
qdKrFj0GPtOSjj/85vZKzTNdCyRlerTWIiKJRJbKbYtLN6S4PFwZuAJSaUtHTXiIcHWLV1Lq+dDB
30TWiZYnulfE2DXrvGkZo4w0nEPf6KCpGRQfZ9Hk8FrFvQnRUYljAvvuXn3V7vV0JcCuaGQbHg9F
qHhPC8naNAJ//iVVhkVaKUy+GVxSzLsi1mjPMb39PNFf0d+93idYWYXypy3UISg/Wtah3IPq+GWm
wtDScrn7+CIn2mRGBI9wAgX33PSDj4jdP+RM2Rd3s34tHrXH1zc8CymquSehjhi5AO9u3lBA/+3h
1aqVvJE8N8Dqm5QVItzZP3mWf4zzmIAkL/Xs0veU0nBKVjxWXnC/2czyteUBY/ka/Meyb5q4xp7j
jKtVwpc7pEjXomivrPbNRshJUDr6YFsWYbjY041ey4dhjBml3+ac1mmupOYrV9Fd+htQucUZB6ZO
xGfUgw82X9M7j5tWkPBvC4xv0fsmaSDSKj9XIjgO/rQAwzWOsK2ONqbHmKxsVXl9T3UuIK4CIGKp
uUx8n3ku0OZhp0NlwM/sAKUqrfL9G1vE82PW5L5wEPMvmFjFBE7HSecH9FyElIG5IWa1HhYCgif3
nOMTAV/H9h/qp2qhNx+d0bKEIuYcj8NCPNxAib1E8JGvtC2d5CUwSzp6RV1lV7/YuzsTZRYiyVh1
tiRBHAVVuxoiGwBTlp3Tf3WFKOUK6sJmqcDG9UmuY2Ve/ZDUqJLwflBTo+SoWNdnGuINK1eOVt4r
E+E3Lk0njlDpG4Wf4BshhEtdyJhZTGLE8FQ+VuhSd3VCFR0j3wiCiZrbUSIEyx4EJKV4ObMk4fdP
bCcmis7DHpKr6Oy8K/tuAN+moDy6dev+0l5MR17BDD/IfzRwLjVpYb9YutqidTV4RiGJdsHsQNeq
9TNaJpZE2uaNgVoPObvSNlczO1kk5fv8z5RBC01aw874IL5aiUz/mTYnsNro2fu8pX7DSBHoV/ME
RbNr+uJ89JEQL6G3GImRow9Ebs8aXyk4064tQh2WQC+awyf8vDMxJC6mdenueV2sT0X/VwUvTKv/
EnU8Z+viFp/KvWLdp/abVolP85qpRZYCjkXJJBHM7sKNPOKewYJ9iBBbV4jHtJIV0fcIJB76Oj/7
ypFld7Td1C3oYZarnetQrbjkUUCyHS84ZBGLNdwG6GAA0BI5MYFiViTxYvPrP9zhzkcE0HXW32Qm
sov6th2zXf8gSB8Tpk/yFPLuFZ6aSE2qNAf9BPXoj6q8sombMhqNEIJjEAboxNPfyweeMTByaDM5
ZJZlYWJo3MjyI12SStgl66VKA6MP02ceuSb4p0ewlKZC3ExOjGzft7udn48zePQlu68oydBKRP0y
+O36qDqcSiHn66xluI/QZpX5GnqF0fg4Z+JG9z2UtnRUKhNFG6C20XuE0Oot3AlaoVYXiK7DLcCi
4F7AeloP1qB2oVjYMFzTUEIet//N8XXLqi9qeiFs5CTuvtFNaDBk6ux0vaTdEiOA+Aoi2KJEVxIO
5oNuabZUb/lWvmXQE9bGLdc285DyBho7H821TJ622HnCY5Dj5rCRb/1AHHVucBATikgStHiaya45
aeqo+EeTrdbHdTK2T3d76Zpf56A99+gw2fAkwD8dxibKA5a+JkQfuHS+yQT25k+oL1sazKDJ5qvi
t77bJ6Jz7CMSbNqk/LTm6ZNC5MF1Y7KDhEcYQXECbMOcOUs/weLN6P99LZ/D97Rio0V5cfyaTKOA
6cOTi2eweoE6nlA0c1JY/jR2x/714LQ00Tebjd4TVPCmA8Ju/mlQBGIdqsKmXzpADvWJaEM6me61
3IXXENTgluYcIL0zGXIj1mVIdSyUcVCXUjatsh5gu9y/Vb1jp3+dYk6eyNAgZrDXC93zE7Clvf8H
vIEAJwMpHj4Z5zxalB72N82J0t+i5oBatY+rmH0028gTd/sIUURXjZayj2E+Ls0xrduWYybHF/vQ
8WpCjLanJW/69+1EE+7jKFuS1yVMZfaaMVwTa8seyazcn55xD+sGorZejWceE+gQH+myYzV4D69Z
S/DLNagASLKftbN+iLvsi5YssKL3L40ZD0RqmGx+BbyfuZPZDCDSCEq96PbvkiTA6hk9l/MDt9BS
C9cUgn4iLce/w11OyHRB6oDcZYyn4+wLtHVv8EgmCtJUonroY26YkAeoyaojScWBCoe1TodQ0W4y
JQ5fXpZz1Ad0EuSOulMAiOazRMl1i/8QpXJndC0/F4SgCjmb1CDschwhfFf93ggpzsPr67tN/iuf
eHyizbIxPwjMTtHYhc+vERCB2XKhiv6WBntwohFZZQOlQkqAMWIEuOJ3AXvF7ZsCDsnCp0LWVyQb
anISAWgUq4HLTG31mUX/BmXI4mlox186VhL3G/f1xytXlFwYkfJHn/77n9erMPoFm7YBuBzP9mhr
AVWFXv+Z8Ol6i3maNSFuC21EsHUR95I+jzwd1wOfVTGiCIcXnQWOStASGe+pHuZU35VgWH4+iD9o
sxZruMzQ1TX0Xh1RZwRbKDLs7WqDX9qCDsiilp8ttlsXXCF29bd6lDXLyaKpPPILAmGxdgbqK8LP
C/KaUr5jkJY8QtWJOAfPq3BM0cSzvDZODIDvSHw7IKxKkE8bpg+uzu5QMBBMH0nW8CHCC6WvsnKC
fQJLz/fLpjlBlBfGq5lqEznarhKQ34d4PnIouBnt/jt3U8J85w9/tNc9sfh5JN5pxiCsRQfVnSAP
Si3D95BWcWqc3w9aclapABldqbtAkMYtmjk5gtZ3QiSEZj3EJSagTSL2BL1CZmGanLsVgN9Nxk+5
4NOQU/PZdTv+SbkzV/F4nAOWd8Tv+nMuIH8+/zqwULacqAvLpeVmEM1jc3mMk0d6nO/xxDE4OEQ4
8+RqZfdVld66XTRKvYh9+aPGgoxcf7DZYEoeLAYF0W+1arM9PaJk6/6jUakYYoAcXSB6R3J7iHzF
mWtgulJ6WpTt9xRSopFJEWnaCFp9/iDzvNqKIibgknaXX+60oyRabTeL2uQwigFXWkQ/542Df46J
j8CKtUPf8XBn2kpKJfuSOXG9EofkviZyoMKssQmZfWsTMpAH+/lkfbG42gF3QFoKAhvYL/Pqw0F0
wNZkFAfwKz6HLUXpScKROfn6YLypsIa+C/cT6JDrCnwckNqyolxCCysTufbtb7b99z2++0Jys5J6
nCUE/RrM+IELWvgMyn6AcRaT7QAav1g0aycnRIAowwl8vreloAbpumdTu1XXwCzgelMZIc9rXSwV
QufA/1pOOyIlS+WF3uosY26QCdTpqyiFgyNtFKwrOTK2GCseGB7S5PLLkvkxbPrOGeUiZ5jPDMIR
1x3J1OBD8WBqv+d4mj2eI8rMkTuW5Z7fSoYShhODVmBOfWVGrjCAEPeE1T2x7oDkflUTTCo8drHL
pFcZPTi8W9Lp/oGGAMUG22I6AeFmk/PaLUaOFzIYPNBwHFg0h+PVXWa9a75McjC69i73jXpRA3j4
sYXm5a7qD4At3qDfvX77iKhr8TfC/06d3e9j67/26RI2PjPTSToAHiEd4cKgHIjpTG9T94Gv+ApD
+ZilkZGQmdsWXlIA1440PB40OSTUjhiifY+NNverEZV+9+n2astyjuL/ID1kxzvHTN/v6qZcX1lH
umV5yH8uZGSixLnfbd00JmuZ5tx3pPgJWT10a1nqpQCUeHJsQKw3mUenUj+ffcBqB9IbpgoeupCc
DTJWcUs/3pR8B9crh1c2XcZT8zA8W1Yd5SabPzAWQGcDfXTLHlCWSnZIWIszTI3VyPzhIARvKAJ+
/pb6TK7tOA99PPdWg1ebnf7X2OBPF7ejZU1XHGyluy2at4wRT93m7QityJsfKe43TQjY41T3fn73
gTszfdKiwLax/yR74i6Q4vTkSkFC7hEZ46NWgTPX60jxkIHgX0KC8rWGqRPzoiky6o5tf1Tz/mhi
8VxnTcYe/IbvXsR08PUzBBXqpUKJH1OtIHS5qXDbi2Zr8WhFCAJo1kVSFsbQrqN2cyo41knUVb4p
vLLU0z/uMHol/EZyDrL/YqCW1FY2G2CVtwKTB9Ln8jevuzqDweq2XyLT159ptMikwuNyutr/rz0s
qzFSva8yAQXiWwtQr0kxW7ufqXqRt3kPS6f8Yy6575n6i5RKGSaTdIbr24sYiQwdTJWSCFY/iiBU
bkpAp5AfrKbHUeSOlMQ7B4UTSP/E1Ql9GH2oI/yE4exjvR7M8NM9vQrta1adCByS4ZCbsMIQ4nWG
W1CL1ytsb99YkmxT6aLfTzfFyt3lSaOv+UuPE8Pm6g0Xc4woHuCD5t52g2tT8z7lbjN5q9qz8atW
UL0wCB7oqPNFgLwM7rzVU8239m7HZ2Oq6YFLVfJsZWhp3RJcectdD1hXf2/ATuIN26nKhznjjWCn
0Qf09f6sjbToh7+iXJVWAEFjb+JnbCTnCZcYhotRhxWwYdNKue26gSB8GwBd9/3LH7WHOcYegHy3
lq3gLm1ipz40vOOLw26qOe2pO0XTaqiy5D98rMopDxUuxsD/Iv5wFDijXlxXlGEdxk+pTNSf5x5n
v7O/wTyeAABHIXzhUGY3xafF/O2HJEODZe1rsFG8qM2pUUhWQoEyCW41DubFXC59LBgBiJOfV9Y8
uETZ5U+2SfHIevvJx1iUvEPyeHXb8SkBE7L8sM8E0lDgi/JMxMhVJi09+DpOk1D9mf+2wLngtlfO
EEVu/Kq3oDwevtlB+0SkHPkIOcmBjQeLi0ui0iagk7AYn5FFn0k5nfblV+7cO/v271zDip6lSzRi
UyTvrk7L/Qio6xY/EmH2bD7MTVBJop4cd4g2W0SC/lokded2Tv52WVXy4OgpZH1Ytosh70zaiJzm
fN6ofuui8SyUuGrglbmWDeOfOyHa5VnpQpz5clAhVCTuSzreEfqeBZBKUvwV5r+EBE52BwQ0KDz3
W1Yym7m6DcxkbP4DUGxZKLxCC1XJ1zfWeubGzD9WllnmE5DRPzvyVgMxNZW9K3FU/d05O68PoEpe
sg0D1zw9qRC4lUb82ik10/0oq27quwINw+QSE3deMKZsYtb9X1Dqk3OzOXBGZ3W18tlAQmGH+E0K
Ix5OE9cUTh7DMCjOONpLVorvLWnmUg0ESeZpdP1KnTGDfbHK1YUaRZOvxcW+2RPejd4IAXMftlwi
FEsq94CEhDrSZT8b2FgGIt73HNSX8eULPGxywvB9HY/4le/S6BoJtECjZFnBDXEKNl/yVhnghlk6
9/+JkVl4mpMr6AzYRAYUCyDIhVDNPwBlRR/qDxRj+uL8INiJ5AuTaf1MpPts9qloKHD65/wSTih7
9rGR3szokS9ItFGRGp6FagClwUqbakSbf/kzFCYcaTwTq/v9jJpuiHUkGfs8cCUjKs5zatg6fhEY
HeF20bDhYyCby6yWmpXami87aG+5jztSH94ug8dEU8oGPP/TGt3O4JxpiXD0XB9Tv71xu76Sb+8+
BjOtBbsXZnhyYY1qJmB+AxhwPXvOJ54nqQyVkSVE3QeE0Gw6tgxIukJKUG19G/a742ka9MOaOj1M
gQdmVzAEGEdAvEnIQP7cctvezB94+c7+GZDi/qb4cK3kSbTq6sep6RjLvexUO/28LkFzk0aSYqs6
bbg0uwvxrYdZ2SXi1il4iCwsvoC3y0tbnFw/AdeRK6B/8f0U8K7DE/6+/KqdaU0Qpms2sBeFS6C3
HRfJvgF6NtZ9uaqrwM/+5h8JqbfrVokD+hE3peqeVBaEnmX6krSFAPLV+6+JeHO02cQDXzL6w9zB
RT467/w4xx/DSSf6S+b+0gvnQkRClL14I0hwwE3jBXKR5CFVbYcSFTaXfZYCVi+LZAWwSc8aflvk
kWsCAaCsodbcbt/SkcTOOn19ANHtsoIOdKtOno16gCXR4yDzF6w/rRWfSKnASE29Ocb84f+bPnIO
1PINTY0EF1GWa/6ej2pLWbUEt9HUnQG/5gAKd3ke4t4sXvO0JePsqe/XZTNifv0ZkanvwoY/l6JQ
y3sZmEzrzOvbkO5lQaHWwTrGv33rWZh/5/BD1VisHsFCQTSM2AgSAbb0EH3YS96WG6OJgbfvLQne
iXXTiRIPeyVEvNn35ACNUMYx6T0RSedbvSkLuUJKduXag94D98sYL3kKzJS/KSPM2PZU0wDlbZDL
KzYaRpe1bEpH3DQsX44bX8F0FSTbQIjNBvRYUO3Bl+H/Gzr9BThdh5R3MOPoG0Z8wN+TLp9LmnME
UYAiAtY2T0Xe7uWNuSMBDMUzt1WtgKpoBPfIKpEU5OAaktHZiEVFkc+M16I/KyP3TEltmC+2jOY6
Btxm45/Cg6D65fFYv62xNVUko9TQOJ3kxTVe9Y3oeggL7/O60OqEhxc0BJmdemOl4x/BIh+nF+E5
BcXzUlD/gfWAjjiuOARhrVIGmnVrzESmZ7s10AqalsytNt/T3fPsvqaPh3sbq+0Zp193SQr6Cg4z
VMXZYhNxWOPri4FK8RoWj2f7ZVrfK8O9Snd6AtyvlkJPb3UpNqyESxzkw2oTOf5hxMR95Zkqv/35
41Y5lhSxjE+2cyHx2MFnH75AfbTS9ACmZzTmR8ljZ0HqgVFooo2ENuV4eI5QerqgoyjngdYD1Ijc
rZQI2R3oZqaChR2SqTeXhRf5mqIZyxQdncwDdFtKpxdpODwEKFBDfQDOlNoPcG7n5nqoMbI/WsKN
ooTx5Q9X0MkDFjk57GRloMKavxOkJ+wO/tRQa1DV/m4k4blvxFTAGu8WT6PYshdTTXcL9Ee/DeEs
Kn1JHXfPyj8zVzFwKJmCUU1+ySiCt0l8/fw5etBJ14WjZgtalTn9nTsMbZjqGeqOXqxvMtc1L1Oi
lrTUMj10g4ZWhXa2jgSCuiFol8D6vLosb4CtLt8ntA62rAOydnFy5/wK9YUY73XxnzuMh/K5IyVc
cvk5uo2dPiqjJXOChr9dnIFlPwVewbrMTDeEnD2FJrmx66E7Pfkka9+Ws+2bSECtNPypuyyHm5dG
1U3K+ZS3Tk/I5Kp6O53bKSt+JUSkvyHjFtBymwhBMgXpmywxaICAwnU4WDTENxs+T55rJ8AWcr+X
mhSd7TPs50p15HG94ZS1EgEWLCO8NTF7cCGX8iBXAhVZrFo8XR+RAYQCWkOQs9QKVRUUi06XmAyx
z5iWjtKiqSJfSVmP+mliip5AkzsTB/i0TBPQ15P1Z3SEDePZGMgd2y16JyUyse2r8Yv0cgBsQBEp
alvQplsIEn78MdaVJ5pS9KsNoF9PZqfAm4fZ2FkKc5GVRiz7viFXzFO3O5wtWTCF2i0SsIz+bw1g
/5fsjCUMjSbrfgIsLgP3ZpqqZb7R5HD2KuKl2liqOQ+/ZSlSx6lx09hM2m5LX9GIzncEKrcIlE47
HLmwffxYpXXHLkxQfY3CGnGL75BaT/+mwFVn1QI1pQXXo2+dm89zz0jzJw8XKcjI6IDlgmUuljqf
mXBulmTRAtNkGxz0X0d4R0BFg19zvgk9ye2whyTQKb/f+wCDPGmcZ86LI0XucMC9Ksv7t8TZW8qS
BsPeavXfaxhbdIt3H4nlAEuz4IcJ0nvcP2S0ue5GWNORq6ZEHr03Dv47NH0vMDUf52XwADQGPFKk
FbW+RVqBNLH3KRllEeGtvgAcP7wGMC8w1IQsosOAq0HjjaV+VZt9v8uO8P39neio3ZlPuMyF8Tsm
yFf4fTMHnUb0l23NeUJ4h0xqIKPleLeky66XWIbWr5XbvRRfYt9WDiY6wVRm+q/gV0JCT40zrnTQ
RXL6toc09udLStN3L6HWwUkp/I5jOGyRPPLqvO0KNGW5QM8arncNqNS5AbnDYL6zneszYyu0PcUJ
20wn46g/c1Q2/SRXw2cJyONxCvLVv5Ls2+SWYr2B9HMVzvNO49u8176LWBc9/K2bkS28c2IIy2IA
wY8v140ot66ZCmw53RQ/rR9/ooc9g2iyHTarJbJI52O+KF83YBH7jnLvPcjH4ZX2nANO3WddFupz
3Q/SOz8uvitsh+0F87OWHDwwNCoKoOoG2OW//F7+u6Pa2bQiMM8jWYoh3fcU9so+XPiWKZqc7xEB
lRWL3DlqYCZgyTsc8knK5xwxXsgAB9VJ4lGjaVfOX7fL4MbmybxOL8dyc6Xc7c8oRQbPTUtZJRVm
1bmqwMLDcSp/R8sXXe2BNk0EAAXbDGOlJkD2W0k0L7fON4TSwNsyky3wnUg99X1qDTFcPlMKj5gN
ARpSw0j9DIcYIHOvOjPh3QxJrW3Z2/6THqiPjIpJqUH/mP0/dcIBGIQm/tUdFSQExzDCfLzy7DYf
MwJ+aoUWjLnoP1Va7hCzHnD6p0AEjNakRyTKTzXVaDEnQL0Z6X8VUurDKSZDBSGpccSpC3KrrRTO
aip4H2SwtDBtzrMikeCGuWVuCSEq8B6GhCUWKLvhpUaNbu+BBJfPvgZAWvpX0jHteQdQekPoEgIF
e8xivm91/g0iJJsFQScnDmjQO4CllkDF2BMv1W7Vijh9izXPbM3TD4j5vSuIYSH6PUuZJ6E+wsqY
97mhwVcjSVRnQyc8xKFLR/R/yHCg2aMYBbz2xfaqRLY9WEmuDstjrPj8FkVIgBgcPqvzt80BFk5F
GJ6/nhE9+whbUZseYT1iKqF/PjxkE6rrq0srPdpOnMepEWjJz/cJT4LQtej96G7QVPcZPasFWFow
oditkshFP5jDt0NTvLcAD9BdlP0OXioVr2l9d/O9SmRdXuf75iyIeDUJ0iNYbvut68tG2zE9ytB1
CCyGzaR0ltD0UN/AvXBYuadW/oa1ciyop/ovnyPu4kJahnhmEZNg8m2FRbwwxzCvBWRex62MjIxd
w1JyTqMuhPi8ddX32Zj51I8OBE8IQ5tieo4AgGzy/64PdJB5nFYwjCqsQs1hJdmxaMpYOLSUQHiI
AgubAwTeDy5wyEzyRrgd8DWw5fbEtW00dV+J/PO4kl1kOW7jo+V4p4YEKCcjmJSdICodte5G4ogZ
EgK0rvzx13Dp9JwiMSYUTX1EmoqiSIFZ0gEApdsE3cntbeQC0JgzpEuyY59rplrI+MRJaDXtKACT
9KGbj5kx3wzuUdNaj5LHDLOCco017joK6Z3EGGfvbi3E/nU5XXhjhSiTnwHh+op2eoJF5gq+eE0G
vCoN+t3mWh5ieTWZSemrDpGXRh8lCe/RBf9XnIPwn0O3dCTGK3zP4VuVxXAZIngBYZYhgcDQJf9M
cDW43sOjcKJts5VrjGIFX6Ly6bbul8h4O1nMAhxvktXNK7UFXkn9HDnETVQHi23wfCJxYHnqayC3
vpdqKAlzJ7/FHgYmZEvdZd7rfBXAWbfzNzVOJNEuy/N8Xy8xcWxSQUNG4MuNHbx55ADqk7xs5EQc
roF0+F/3syHRxf/NSdcMhwIl4DfTx60zhUuneLT+U/J2zMnov75T6+R/lwtbCO+FXRBEvlrSIACB
s/z9Pw1tMV/UwRCSQToxW8LAtrhRDX733elxS+sAlCKV25txNHWlKCEFXYx2ZmOLAVM9LYnyTFZW
OlyHiyrNNN3+WB48wcmH9GUSQ6qaUhgVkpbzro/UP3N//ZfdoD4lEU+IKQmsZ/rUCe6sSiMwrljg
K4pedgwt2b9lGfAGPSO4Iwfps/gAtHCyGNKTfgjXNb6fUyujZj7TAY4YaTgXQih4fPwwOuh0wYzn
zup2qSFWdjoOdmooVHO0kjAkB/Mib963clelNCXTt3ej2SrCf8RU1RsWI5cozg2IDETa7KS/OOKS
bDlXLzdHfEAR4cqiZU6xZL3K3NGaSUuC542yi77Gp30PZshniZ5rytEOx/MSu5etv4ExYppI/fxN
IU1zJwxn6R6ZlBwprp23hrj0FPaFQCCfwYMFbwZ/5cnQ9gBGAF2OgHdhA64RKob7mbHtEsutZ9lc
hdj4pRI3MMk9MeXdjB/oR/KIMuFCF0i9yoIoOIwS2NF5pYILu+I4IrJ0fCk4REHKLGNgcxquHmK1
BL1pxBuDcS8xi8VxUTmyOg4GH6FQTnPksGy8HubMqNnvR/XxccMeighzJ07+PDtMq3EK4Jj+Rv46
FZ7bYlso76ZDNCW3IrOMtih3M5wgI58Ih+mCg+3xwYnsckF8IhCas4vIHgVn6blNRaO4E0psldm0
UlCiJY6Wgw/DcHfLmEJahaIHUqmlGG7nWDAnlpqDFi9XQg7Wj+b/VPzwfGcp1g6GJbFwjM9gR/5s
LDnmEFq9PTRB5h6/lvIoV3KDcc25mJAR+hhiJUPypZi0lxvE/ZIO9hQBWMBdFvGg4Ngp1g2C4kwZ
hKnb352NJ+P2fZ0Y4YEPpRxVUrReyJVQyTmGBTrbhW7WbnkS1hpnfhFPO6rIDkgmlOqvFG2XASXl
osIL9cnyLt0JaOrluQemY1GitPJG14a6lNuNI8Qy3gSbatcQ0Zmrtkqj4Vj3+6yM/l2pf4N++YtP
CgvgS4oiPEvrQo919d33QAH/u/w5cHgVXkR6oW9Kc9fnp2VcARYat/92Y+aMSrpxGTvSKyywmgue
s5COXLJUhmNgIcS+BDYslhq8uIhg6N8Qn5Onrrs7CCrSP/dn1vGbH2pxifAB3nOR3q7g9EPc+HzO
/OcYbLYRHFDHDrQSKmRDZxZPVVKf6XdNdPSiYCuvtdFRztnmGCt6zw4pH67sa1QLxfATriIayav5
Xnz6o51FH1xhnKHwHWQ4S6Aw3yyPDU+ZCwMQa4mfQkE6Az+KvtgWLs6OAjrzB53wUC3cgDroLeeo
ANbNw/U7rYW44mW75lcQvVaR6sVhpUWw8atGryDyBM7g8meG03OGG6iiJ2e4A/h/IWS/L8wfyl15
i04EzbYXaiHZ7+3INzqDezHSYjxBKk2MIFuJdVct0XGUG3TAdRqDYkhvzk5OlupxpynYHLTQZPEQ
+KOloG9bY4oIHv7Ow4tNGRoMTT90nOSoIjuaOC6FJl73W7ZfpgAdOb2B9g4cNP5z6G8XOz2yujuk
vY2bjmrJq/FMBClxJWxEtW0ddi4/to349hEgrlm6xJPWAHRSmP1vs9hB7x9HEeVZEa7lFJga0A2q
3RUR8CPLGEF7XLeLGDyHnHoG5tJix5r8dALDOosd9+2jb0wetb71K+eEvIF+J+M4HxhWCZM8sKgp
JqYfM7zbyq978CRAU7rO8xeNrcLb1cX6l4INs4o9NL/2h/8gHOsKpWBUJ/+2TAXBsDwIB1jD8jaB
k8XcuswzhdRvcSaUM8UDhPsjiUL/RmzWnrYq47MqHGhsJ8eczAqK3QHiyRB2gxTM6N37pvTYU1wb
xltLQc6nbeKHdm+GSMQeIsuOljaBJk23xbJ8u5kwZLKTpfM4iXcdAZn7mVI0ZVTqJq/4Yw4JxWrP
UdxmsccC4oY+2IpM/5xUzhZr5mWxVhLbYoa97Uu4hcK8fLovc11FF55z1sBF4KXAr7hdqjtdIeU6
6nKnRCE0H8gBZVDoUbL7f5wjICiSfzLQmGHZ8QWUhRkqEaWfGz61tJilvGSXiFkU2JoWiFAtRdTl
Np5IKa5k/x7S92eUBhIoSxJ+cR9qtaNIRUiljIPRvYvICoCf3kk/HvxPMNp+zuOGFQE8AAF6rU/2
QTOvCnAnsRc//RZnN90q9UBWk9qXyAb4rSXZHosycfKINYRtwdIjGMhq4EZVBopplA6IyAGeMjG1
lHPKIyuvW4dJhlu5l68y2g2J3nWAp1yec6Bd7CK7iF+MElQoriNn25SBWv5+AOjWgLL4qdmL0dmz
wMu9m0KdqA7QgEH238dYDW8iR04WZHckMO8wqDSQU6TE0q7910LypouWbo+bZu84FBQ97q44dVuG
56eSCsyfOWtxuduzr80i7jnUi4wlbpbz25OctMCDiJ166YG+tEko3Ws0Xvlp73CPKPOjLS48S6kZ
Fvpbw2fcj0tbo/oYNQJIpJShUXpTKi8CIGiVR9yGECd46VTZV1Dc3Q1Z2dTMGVpGPoBKAth/Qhym
4vJUBaj/JDoLz5MzADdULTjiJJldmk677IJLTDe6qQXXDr0gX3g7RBr/6T2n4Qa24mJFS3uWMT7y
faX0KIo1a4aJ/njfTm7EDIqDiGj/Udpr42m3RWwEZ+audHdGwt0QWTFz3FTvo47do9JsenPY38tp
4Kvaq1Z/GBhTLNt2yHd8YqWI7AFR073YjOOkrRL6Iw5gXC1HvHEHrdKdMMsERlBq9MB5Ok3dN7ft
C+h8YEJjVwB2U/L1EdILibm39SuSQEwMIOV6cBhI4jetxFYdKgpxhEE4DZpyHjdRLieY1f0ntWM1
B+q8qZUs6ykhR7hsy/k/4WTNDDEx5QT5xYkVrMPRxM3YU9c/lChgpSL+JWvz0yo5Dn/4t8zrkYng
0HD4ZdsX+HNExmTz1XIifSL/97KrZ4Q+bFydLN6afOGMlyUx8rLQGXnaUBCL2cCvtqpvwvxh2GKy
AdBUvgxjM32JS1k/icPtWZvh2K7zhn4gS6RnTB3eemDvJNIpoNRzRKpaUco4OjPju4hJvAfE7i7L
YvwMrdJPWP5IEKOdoWmfU+Y+fj4kTtmtjeDX10jh0BmHyl+o5c0WDVStnhXslOUJW/glWQDoQXQQ
0BU0Fq2UnDP9fxDJzMuwTqddwZEo2DW/+8xwI0wB4zcByQXnvDNdiWOoBW19D8vf1Zy6dLclCtd3
UTNkOMl5HnoqSOfQXcEQ/5ODoBLS3BbCbx6xH0XLEC4eMmyu7QEn4AQHhqpEqJPyB8dYeGS0bPT1
0jtuP9uId6fYrh4BkIasUngG7IcAj7C5R8gghxGR2lsvcFNKBZ0tN1fMIBVqpvrPGCooUDpw/l7R
jZT62fYKP99MSZuPzlu65/oLLBtbkAhX5MATuHej+ZaRVpHUPAVXkvntGSPrZAprBJQ7MTYTbNea
giyNunQZ6Rci02Ur/ZrQ8TEHb5HFtsCHxgOgGvapTumOILwkAEXr9s63bOobic8W3vBmrwBABsVk
0PIgwX2k0hjzKFry3XIeQxojlEEeB/VB6qxMYx2lOYJbwpyja9Jxq40FQu7ZuxzpT5UJ5jYckOYc
+lF9/3zNdJQ1ZonazJ+waldLIoLJGEESzwmUB7zhjo+d/CxcF1/4sD4v9fB9arl8GATnnpPu4Ekb
KcEe0q3PF7ig099OOao2zlrJiudbtxAMWQCpBgvF6Ol8AelCM9K1/h1YEFqkc28ijRELihHmsoTn
NJUUAU2SaQTmHP2OQq+vJ2AMLFz9Yq9F9EhaVjl7Ej5R6WE2M7J+k3Qn6S0UxKO8XRJ6vWg04Vkb
16Dc45EG7Te29I+bnlO2ApD7qRXkfKG/0tOd2aUwPXvz25+5V5A88P1SEuPqscMaddXr20lF0Lyg
mIWyyZWrlk+zInxu4L2/7H4LLtcusXE7ihU1rHScCh8x+Lc+cCrykzM3AHB9WurZe9wczCOmR5oV
DsqtX5ORDhsFc4i3F0PqYeYl0cghLQRR2oyEfz9kvMRlGFGwOMuTzxbfm0bJWaHp+CMWi+3kifWn
fM/vcX9pMt8FFrO1twtdC2FMDSJvCxwwwo1vOdTT1tu6fJcgeoixchDVvwIZTkvrWU7Ow0lVFP+g
HtAm/Q+fM6MXapEeC/fhCNB8n6V7ndY1UXcfcQw94DNYkH0oTR13SyRIJL6KXuQhy1EXq/mEpp7p
RyDq3UG69LbKwQ427Jb3FEY5PGW/y2lTmoMMbnPmotbnaFtnpbXvLO5Mmn/WE9RtCd1uLKuPolUn
ObH0ylR4ph0yMXjx4XIqMR337ws55EEjI3EDGehnAKWlHhjreNmAR4HMn/pr4M4PLWbMioo0Ku2l
ShPiqKlSpTK9aXNDfBwTJFfVpM3YHsihhKAmeJcgjl+cqtagxbDpwgL5wQFLz/Pl3nlMu8pJYOYz
Ju1Cv9NBUM06BSwvZHB6iew90Xc70afgEKHmNoi86qCwtk6PdVGLD5e2PV2Dntog/+1vTi74h/4n
C/nr3ylW46GxL/JhDPc3Nf4qBH4fAk8MejY51I7sXtvEb60jQfEeMoeypzXlleHiJlYui1Q9eACG
hvt8PogLVDxaN5ZkGrpYWXOfbF2koAt1K6aZYKPuhJrMPqER5ZZjku5vO2rTnXdeMKOqvqdqd+bl
gkf403+IF8t/JnOsqppxrn2KDc4p0CPtKO23qgipqLRofus1A9xIdTJq8BzFn2uB6DhXhArXYBWZ
auQ6Ufhvr5XW3QYWy1nyHG2axhfC8dOmMm5xg5/mMCvpN4AfFsawFcBlaZodukumt1NdHbLJWca7
3AC5afmlxC8Mvl6L0z6kxS8dT7wVfLIlJTX0zRCC/HGEqMD7qepzRQPgY77cCsqjS9aQIakcS4/F
laajlliQdgzPTEr6Zu+Ist+I9YsMlMLoIDzuU2IhtC/ebhBbALFSHMGFMBLKshzhEAGGTLX+/U0Z
qumCCkp5Y8OxaTlLZ4hZN1XPTeSjzkbIkKLpcyQmKuGrmt5TKF2LdTpF9CRNzzjdoDFFfOT/AVLs
Wp0OsvvufQYV060sGxLH9vjJm4ljX9duW6b5GewJJwi8ac0AmT6lVOq4Lfep+nAQ0T8ZUGBaqa1W
bkrSnQS2zyHS3hu76F840SpbL+NlXMwLm6ISL9IssutrOHftwwY4HBEzUsZopbItEQT+K1SPCyon
oqtNSxvAABUpvRsmMQEkiLDP22vBn/lSHau1GWtXvGIbtLh17bejXcvllx+RbuGB8j72MTDQNurS
kL2BafrH6858Duvw4kQv9WtbkvBAgA2dqcTgtvzjkZEG7tnPtSLadQjplZSR+whH+LU83OYfQibc
EVBjIktOnvLNXmy45HrJZ6eiwYPCJTOCiyI9xftqeYO1jvcXSf87yWEd0SEWr8Zjt/3wgYDJ2FBA
0fikqq+hAg7idLEeZ5FQoodnIq+8nDLU9vkzCTDg07ueesq3Aiskg8IL9MFDahXfwq0Pjet5VqF8
h4EE0+KaAM/JZ7kzHS6+muA3MMuwlfysu5UU1UCXpJSToKw+GYlNoBDiw6H3YtiQ2tiaslb2FjtN
8Fqvw0qdV/2cmIygr4SDfwpyKGMonBZsH4VGmmMBVnSrFm96c/JeGCgvNE9jKnwP4Gk6fYv/3HKw
pfHajY5HrBCsReHtFs8ESbsdSKUNvgNPJ9mXmawhgrDmxz4VNdVhILst9axgURp3lr1185cOFQSE
Yqhes3cJ2MVDGz2QXtRKfvIfsJGiKUxyfJkMqQRyDasQ0TlD9yRDd6SKRaaiZW4Mqcc7ogUiuQZ5
t/lOhMKuohpBIL9VFBYjh+/m3sAqlwUUcE3MbgiylHHgd/u5LNX7N5FXrSTYOlhW7IoLnRpP6mck
KEtG7qb4177DgmBlvyEtjqHjgv7ovWsYb/GJaJoiFxspHKx5AObmPxVptzTk/L0UjNNF01MLje+O
hXV/O5eNKB++tK1rIW4M8axQ/nNe4PW7Khp4u8IR+16gYWDCEnqMbU9gPB8LtWGtCXA2Q7syavoX
wLHp4HLPRavyAwXwInxJ4DPmUlW5aWkwIcOq/XzsEtDTh59fUtffodaOZlk8xwGR7VfQRq4RMWwV
7MTRS44yO2JeFJV0ZbUML4WVE9sAXGrfsp6QcMKtvguJ9JH5sANq4dl2GvHKY5VdAhjCJ4TpZEsL
PLdYRMaVgVq/FCjuuLMXfTkdRA/6cmz7mqKx0D7i/8s5if0/q/W8w6x8QZV6bVOhfN9A2z7q5EJB
Dw7bqux4LfU7WOYcKN0BZ5fZoOd1CJ1eLaoH+HSY4jfTPXy7pOW60Jaucim1/hd6yRFR5/nAOSW4
crNtFw/a8vvZ4SZ1mvyrY+NlfxsU9PKFHiLW0qQbYFtguwSg334REdeXwZ9vOcX0pflHI/gaAGZ3
wlv/BZ4rLAkV6Q7EOH22PjL330omfpAoTF8KTkss0k++9u7LNWKKiapIRNCf0nUHwB8XMOGU/rRb
k6ygr7fuzJNm5HbIf1uYeBSqfF2TlHBWHT5HEO2VTxhhFp8vo/9afl+xbok6wT9ljhJdRHZzwW7a
PWCGsBM0loBi9JFAtXgeogCfvbeoUZCzk8tyreLuJ6c5ufkMvMVe4KQ7AWq//iR9Shy3D/su33vE
tV7T33qZSIMrrC0Dm16iCjPxkM0NucEWYYI7WGNabynWD9e2gPC5AgAfqkDg0Ibfd7YoLUw+vwL7
WjZTZrgq1SwZilNW6fC+0rdGWYBG8BJAHONgCGM7Xj3venZnw6WSlhYjNG1XrzieGXHvfBk4KKJh
5hHrJ0d1HWSwjWR9dzB9bmBZYm2ARQOMprLlvqCSS3ylHyn9Dx5WoQK4C6fC2IzTafg7s32EXsmD
Hk707sTsdCA0s3q8cdAX+1sVYqXfLwFAE3WRvIJygMmN3MyX8geAbl9UGJgfoS8b6WWKoN2Zy7p8
tdMoa6abcO8RDZKUbCTvW/KXvM/v9sgPwC3E9vSO2vX6b+2ruaBMOOgk2jtmq68GErAmy7oOT1Vs
Q8ZxDiPcaESdoR5FzOJgl4A1GfenUgkdiIj6nuDirVsQ0+D8k415lQd5FOZ4F6ccoEoOeyFH53MN
l3QQbqI8Fi4SbMB+WG8hed0Q2PoiEB86oIvnCI9/MahwUnxpLPgzcbCMlRMlyf/Z0Zmp3hljVNTR
+Ow6YBB3qS+aBcnkAWkuPxDA2RKonJj5fq/CjXR5Y9YCpCgYSrH/RAyAXJtrazKo6qHknbxxHcTs
u3nEEs9+JMkxhK7bYqCHZu32y8HI5uDN3q5YlRWwidRRSluk4wqKgCnbA1cluDiK58wDNECdQDrj
lv9r19PVPLJRAOOhcxHEq4nU8KTvaqsYDBwD532eyInXSz9F4b5DvfHEKaU3xLI67+pJTZs3aPPD
kWTP/Di0qxB6/rvXVc9HyzZJ1+D0A1owHxilsfOt0ju1LRilc+RsT/w+DViVi8GNzQcl99GoU037
hEEdCY60YbOs31iT9q5nJUZcc32pR8DrxNshR643OhknP7htK1UYe2allioIjEu4xb1SsmbTk4Sy
xiwlDy1ByWtbU79mE2aEybtgReh6FPIaeLNHOho+rFSEmFygYhkLQ+8MbnuQih1HYtqKc4RztMR4
9YleCOzUIgS2QhkmI4LoLOUMnzJ0FqhF0nho78EnG7KmspSFX97AWciub1aarZwuoXEMjDprnvd9
Xvy3x+SaLV48X8LJRyPsn+/NjGkuU+Hoa4ricBXBxZj2NH5lC05TLBHsEEUHB2sSX+3zylYUIoT2
cESdI2Koo85KCK7a1J6Sty32AbGkwk1ZYnWevIYWIYJgjGeHLVGhyNUE+VknwlmrzjD82PNGMX2E
I1HJqkiyYTnw0anRuipbU0p0WsK7az1o+fiTkaZCrcQJ7LqzhZ0rOJzUiZhas7vF/Nk5iiSm4Hsq
awZRx/tMpJbZhU5h9zDLOlmjqiwABuogE1wXHUpqXYljcCuKibpXB3ku0raFiYVs31dYZmhW+JHZ
a71vvLEXV5PSkSliE7C5yCkwxmu+E7Ign+jZpi9LsGU1tpV/NZp2w1E/07EZ8ckUwdmSqQzpTDUo
hghA3QJCdDOCwJwVVkiF5AKETKRAAr187Z6djew29bKX41s5dCvKoB/p/NwIfxxQ0m5gyFTjpcN3
2U07W5yXv9h53kbNYJQGooHm2PtUp3lr9DSZFeAtSIyqYzjmzwkm4sDi2vrSsTGhvunMGZAfEAV5
YyEQlSMa8Xh6M3tzRtQkYXR+xQzStwsEYK6UMk+Tn4/Z0fOtUZ3iMKnXuuuPTuQOz09O+KLswglZ
AnJy5QrEt37PG8mhHhs5KdJJUGnGDzn9wKFG2Z4RKH/xquBuMNJr12xbSImJ3kMfWpQAQ79I93i1
KmGsQjfYxZhv9zrBK0VsyJ7vpeJ9LcaXNvUhbTEAt0kWRWE32v0R3zd1MG5mJqYre1ccKtfZDDNG
jvsMabry297x8o55m/7MC28va/YFu/WykZhIYnx/J8hbHu8r0MZ0Wg0kPaIZtvLMakay6zs9SuVH
Qm2JPkCd0Tk9rKTIL9F5umYo4IvxZXD3EmxnVLKoNS6T+fz1vhs72HNU6/fLqpHzy5p1xCa+6gHv
lsUE0VEu82KLd9b7e0AU517mnQau2nM/EX2HZqKYPCrYYDjNpTaLxhXiweibB2eUdD0lazTW65Ls
cSok9EC8lrFenpL8qQX0myrksQ4aigdOADQ4Tywku9YH4q/g4RCpSQ2H/6fj4c331fsDwcmnznNc
Pnfn0OjZl9u1OW2Fg7q5a3pEP0ykKZurtuuftKLx2hM8hF3aHqSTjiraly6R/1bvezzEkru7U5L8
otXha5VBnjlUCyCgofKZlxaHEvkc5Dumz/Pr1hmBx6DC/k1TQvWWzscMI/x5I+M6uxkJsOBEc7Z7
M3RIqVqQM44Tk2Tdqtc6sNk2kyd9MZhp6nli6/9DMqxoXkCfdL+jsXKDcM8U3ITq+Wgn6CWTRaZ1
QZDgDJ77fI1ujPcW8MqCoMCymFeTMgreMb9zVeiumc8tpDX6L4YYQwTzmniK3wNR8QG/vsGfdQVq
LutdIxVtz+zNOjOX/irY0T9rx9qLiTrjA/Ym9zmrOGZKPb/Ggy0+Iu/mkT+8QKxR+8/cPkLlSPI6
LPznkMTvu0pXPOKSGZNIZLK37WI9/ewHxU1ndb1AzBA84Eo8iUoM7zxNW6REcAJwPpPLJ4QK0I3y
1hD9a24gLYRhJ/AMA8cIdKCjsOH0qxS4/SDPWVt6o8cdILDByKcVTLWGIWjoy78z5ovT0HFc70n2
/72MD+XruRmbXUVKa9/zLx3K1pTAHpxlgkRFUOScMP4H/pzvGcawSP9sr2T0fepbgICHE5/2SMSn
y4rXBIXk0HlTFE4b3g/JOLPF5m993VeNhVQGdcruQCKUdUgUeDq0AHulgjJXSKeRc8ftFLIE3Uk2
U6r7JfijqUq6t42aHF/5xMT9aGDpwdKznxZl4eIvh9vuLGpY7xG8Wf2sZ1J0dhuU9aLfzuuowP8Y
TfDfQEPvU4Psp70S9fFxj8HCR7RQJ6ZoM5jjR9dZ5h/0/Xn7RWxYunqncDaK8a3UHdvdeoK3kTdp
st/hpRb+pJfftKaDwXh/Dd+S/0IghVBaduQKmmqS1iS/A3WWW03+gTO2dYh++ov5YHVjU1n7BFOj
wd/MoQbruGMlQGTGsHBjcaPHVqcmC5iGZqeLf4WX+hSg9dkY8iBLIGPHtthnmipijm6FE/dSeZPh
6TaPPf9Rs/mQlKKz81DhtEnx4eYfxToVARTSXOfD7+UrlDWhQ/I3aIqwr8f9d+ix0YhHrQLErLgr
KinXSMl1spHW6iVq1rdOJWcKjJU5TguSIxmggYTna6ZV0xszDsQgcGEVi4zlqRmPK+Dk0tX/1EFp
m//7ALb1i0fv+34mpFKJjHUAEuNaVqxo4rZp27wNTXZ51YsugdKWGyFbUAKuW4k3HjA9MR0DuZvV
0wAlzDanKu1SRzLbCjSt9Hnuku+K2+dEsQjBGpI+WbxaJQrqJom+vK6H8eToLEIVauncmHJl4BGd
Mpp1UsS42lJk/0EvE+HFXgZRkHV29DOLhKlsED06KNOCy8th6TJ4m8+ipd0yiOJHv9yaXs8jXHZm
X5VLgbBVN5mJigmq9Plwnxt4ci/M/G/BqIguCsbFCFChX/JV3/9DtFpbLxxbbf2ot2hNOxsI3kEx
zg4/GkKC9GfurxSUB0lwnykJBZB/7st9lwTziRrL98yCzG3DeW/YdIs7upw4DZ/ZBCAEGyw49cTt
AH9uGSXvMsbpPjDg52SjNLXi/+WOL1Fd5SC9c7qJ4Y95xoAZbaGPNwJKtFCzExeIDXouRcOIFKIQ
lXZS6lMlr85BTf2OnITj69WMYMblTLPULUrYMPbuzbvBmcmm1vInhrx+kHIBOYv8XMffqNaUaPpk
4r7l9hoD4KfW6P8aP0vAIdkdkHt/NpzS0nM3La3DGrTOFJ47Aff79SYQ2FJvxPjBBMqkjmQR3vSf
NMic/wtzgwCQ1Eyss2KZSIhf5d+KcDTBQuSMZ9o0VX5GEmNH8w4cax4AqlNRJMoSRQu6lzpWxjAL
B/oC0J36xbnGyeCbS+mzQj3TqlvOMw5sna9cvHX75eJtkAMGj6TDre4I9o0Xn3byrs9G/AisecWf
aQbuQIoGvq1K/kIL3rGO4Bo8cp86aJxNFHaFwgjTZq+YgWnl26X2LGvpfTdvGscyFX/uTHCGUReF
4WV1I9pkk9c4mQwxVRa6pS6NfUzb+mnJrxd+V3NledZomO1WIYVwkTr5bbGl6LeHXGrBvrp71z7Y
/zsW2N3v+4/+MC1WiTYHlBmI5rlrV5jzJAnYTlJsCZn2R3/KVt9muibRRbzQI/GQbLwKQIpydi39
IKm/rwJCVImemURmb9fJ4e6820yfaHutOYpBAFs+spd6CaX3mcIO8n+s0VQvAsy3j4qXRmTOiXqZ
kGILnkny1+vUfhpZCnHJQaOZh81yl1nRtMvac/hh+onHhOMFQyPzCMD1mbwUFdaN9r2TaEqzE4IC
NIAC2jeE+HtyKFkEXML2+Q4gDLTsXfQNSPEPS8hLND1vporKRdesEPzDUbAGAB5yy68SUD9rGLRr
vkJWjBOSGIuXOCPTyrPsKkWO70R90cqEo6TmgXILHmpr6T1ABqLaD+/yJKklZnvP9J8m3IhMoZt8
wx2aMX/kEJUIFk5Xv2T0suozCtm0XwczPSxphJi9Is18fsxsfxG2m8AfGDNP5c2lx7Sv1NIq3VBJ
c/00ilohZa13BwpXhMYp/65yDz1TmUsvEHx5V3zdLLKKcZ4pK9U7CJm7j3SrAmDnXTjO+vr9DVHv
XplslPJO/THqws5t4RGGkjywoulld3wFtLzBT9vDZ++iVnEHxSkhRaM1a8hm8Tp/+1Ho17DjjBcV
oIdiiSyX75CDh998+YIz0ZgUbsgP+RCydBuQFiiOUwyUAd5TRkPbVnwVEObAXyni4kXGXBU/FF/W
0fccz2rht56EeS8Vn4ZQ6dHJvUCJ5yuZCn+PXg5vGs17QqbR4x/JHKl3hFIIlIImQRSS4Rr+gRVq
PxUxR4/0ubz4QBcANMpe52dUClYhV1SbM717NdoYmBWKKg1mpRurUFD5nl77G4FpUIQ9ESAgSiCm
2sNEr1z4P2cLe1YKlkSFQunFM003oTwLA3jS0T70CatApPsObENIyQxQQbMX4OScz4LFPBTk4Ww9
Nsu20BejundhQE1VCvcoDkZCAmeXnyO63QohO8sIBkkIzn/HSV5KguR4en6mYX/S0J5d0WSX8/Ig
viy93Nr1g8pTcN3/QqwtDbv/Kjpr5VncwoUq38aMvZfi1UCaHXKRBlRrBHPBXxc4qxjtoHAzcPxc
w1EJx+OTd2B6jHpJs3bHdlYzYYxaqO3J3H5i+2o8lW+3SVUC1lL6hDj2olTSX73eOIDjIBHcUkFI
FzD2416Jgl7ZKZZyHt6OvX+zA3kOdxpe+apHXvbE96/BgSUufpSFXLxE3TD1Rv7dnvho96KVXj/r
GIZVUEKkG2cQrxeaiHon7sfEArdxZ0HqMIenZBOWPmeid6r2iIMGKiFG1z260JCV1W3ehGDtLMlw
w20GKy60RtAKNCuoP7z+ptrB8jLtc8bIQp/n1Do59ESsBjkyUuAErPqPi6lhM3ZAw7R9Ay0KnzZC
ILPZODYJK0w7Gd8dZAg0cXkumxyZPNB8cBZiqrKkCgLQprZLfSJl+dQX841YL4Lb2Z3IFHxbtbts
FpucwqzUhA323P+ZhgsWZKWYAfYxONTZEwJjHfpxIHaKfYvg4GFNLu3+GA5Ob/jz0PT56HTWiF/w
177vpiMz2qYTq2DFFSJZSwVi6Np+b+2yvDJykGHEkyGADA0aqGy/7Y+sNGrw62mFj/Vzvm0vLEJY
W19Nw5usLpspYFj7g5BOCndt1usH7AVqAwKzTwewJmy6ugzED69v0MR3stsPVrvcXRKTFYJaCr6V
WWURk3522W3tesFnpD6GWsmEQskE1/+a2CXVcyW7wdT8ffSa6fxnt1zBB2KoAImfbwwTBbY+RVas
g3ThPF514FIyBqyOpjYwA2Tx5gsxtU77Nv/u6skOYBZKajBV6Kr5OmFUQP/P7O3rTAcKEvuiErHB
xD+Y/W1COtZm7gdI7RUr4H0c5yxdg+T+yJTMylRybngTo+n1X6uLrpvwm6kygTZqmPN0XZt+z6Z6
S7t88yQFyZs2sblzm7+jpwymHnVo//i/tMG8dPy276TDk/J+Ttm5UlXdRibeJaahWTA3OJhN9ak0
g+KGzKKoN9YlEFSZSg5bq6zs565x0NuJC3VuGT+/rNOxNNhylIYHBoSgjp9aQ6UNllGW86aSBHDS
ae567lsaWlj7ZrIjYrJeUc4hqyM/8sQGtkX7ZH0FskVwpbsueEuAtCrbBhsCm1mTU59H6AeIx+jk
7tFQiQxJ6iGlGWSBYHo4+0r1AOBUlv2WRUbYgqPb6tzvsFuGgQmdrtjQgrfmFSA3CSfPqhrIlBt2
Dx9a3ghZFw04Op8m6VpiPJ+mqy29WA0G12H7m9o1nQbjY9R4n72gEiSL7woynS3Xyq3YQKmN2h7r
FJU/6imkZPVikGPv5eIReBCm0EmXTFIrw2QphyMFAyV2iZ8Cd2rHltUnep1eGqyh2IVITKVihhO+
d+M0Qik94e2HYx63ND1w1W//8Y1wAgxoDLmXVOSIYhuta4EuR7ZMA9ln3gMJc9st5+15YDCYxbb5
DJv5N1zl/3SBOO/tMH/ES1mUaXbW8NLplmls9x6REC0EtpCSDGQVbhfDf7uIbq9QE03uolq9VJAB
JM6zlO9o4wfJSpEqnMOz1wS70xwrPKrFANGCbAvhBcx3Ir2vB5ZjIbIJ5H5ZBaXiT0irj/Np2hkH
78RqlFH4y6q6qnZTpkxgsa5qHnSrdRMr1URBYdZdv7PznQUYPoA3AdG+F5imiyCYFoLda8VVkIwZ
3ZZY9liq4DLxMvAsmljhh2HFfqwFYK2TqXHAEvffRb6waye+oGaD/1O+wENV69fT+c5MSaeCnIOE
pAkcSP9oF7UvAMBSqC2ivf2klxQEKnn4fHfrAa4Oie9jAXFvrsHlu4pywdmZEmjBcz8hAxmT1hvT
g345whEzUCennntsK5he8FSQIW+9tMGo45YQAh/JKakBVAjhzJ5l1N0/i/B/pUywaYo9zgOCyerj
IXl34lnjgaFqtE/ygJFsXbOSD0gY5zdrXCSRIAfT7K6b2LAOlcGIJJj3TNh0Zn9nr73oXxC1D6xU
yKjNtKVJmNwz2UMlYorQlJH194dIUsa2vigSizJCLhmOXty27SaoRtdQ8xA17IgWVW5yxLGYM7vz
35H8nPPnBukPHSFoCexxmitqFcbEBOW/n1QTKF4OAnnjKOryuhYZc7bNGLFMXhEyNofeJSKWgoVu
87md7aDn3lQz6MGTsZeYDR31rTA8oVJEEXadzM3U+FlGcEOqJM0KeGCUH05oYvBKDr3ZjzXbLvKd
5Pc/HcG5z957gUhgKpiBIuO5zKBuEeOnCQTrwh9xAbriLET0Ir4JzvjUw63G+Bl/pDsGrow4Xxvx
GswXkGEgmdz1UPKVydBwWrIzagXd6J+5jClKXdyGYEb3XijEomZ1Y3jUAQKcmbbMRVbuqEoKEJ/h
ZdujewNbiYJbzjpJLMDAya/FRBZSZ40Q7K2+NnbSxkRXVHUEDCpdk1O3o8vFOkJZ4DoZYiflcoXQ
p2UqrFq5Nte4FCFZ2MPGi0VPEaixVFZbk5s/Nd/bF6yOsx8edJMa2PVBUpqCRHZpi3PJI1Zj2YtW
yr2MyTvxbj6wOtFCposLBexze7gTsKk/Nif/WFg8963eENcCLg8CKJfStMJjByVqPgaIddOaPQ+w
DLURMCvMkEfVVzsfcpr0GzxB5IR872MU48+PqxfjPWNNBueu55oLcLXKlyNYVfDN3Md2Ggx5e58c
7BgTq/OODXzIBzbQnQJoiC7PFZtv0oiOkedDvZTxrw0w7/ziMMm4KHaENvbR4DJtv7IqHEq2BrdW
ArSdRGD9d3mB7el12niSp5Gw9h4BVXUjxYQhtqIBynoEqb6B1/OzF6Tz3J3bcq7h0d+waMoBm0vy
2ys7P3hrsadGJ+onLu2nuE6mAWPm5sBaCxWu0DRmoVVNmPv3FbPIsFgGRciumpTnmTDXlrO8bDWH
O5AsZZGpSK3miJCkngsR43L8vJsA3D6kdlzobkG4PiixxCZm1+owoHur69Wc41YCf6B298BHSl3q
2zXQZ9nJfMoDem1Fl3wvoFt6qCcQegj6bhhsEdBZxRj9u9vjCQRxZ9CTPxMCbEYhGPWhM5P2YDT0
lf94NtTP50NCy30dHBBUlnBBK2oqmSfIYvVzWNsgQQBBiCBWfcwI2S6i46qHPsl2oM+1kDCpv4XK
+MKjUrU1SCDxCQjB7fNgMQNJLLKYN0crk20Tp2qT/h9d8Xk6QiZy+FZ4yMQk3ogXvaSWUJJuNuJu
IxW3gb3iq6ief5A/LT2ZixmtSmJiq+bVBpUGXtyg3+SUlCaIe/SrYYV0VLhynL8f0yhFhfbZpOBs
h1ieiUnL85uywtEuK8MnLgPLm3SJY0Oy8o/AMnoiYIU9xBot+K1HQiUUxQH89Bfyz5Jf4vqD4OyF
ZO8WnS12FhbEQWMs0C4oP5i9/EpzTmqaQBKjUcFCmT2b89dwCepBG3Pc6pu6575RMLBXx1h8dIYp
adMTRSulEOW+8+fTnlUqghd5rZw90HWxD+UyLQHcoPpkbDaLU2SvXKSJebl5rmBbawDn3mWtdmMd
1CVas86frmuQKd4DLTJRRAKNgi99BQdxa92R8gFp0uix90f4d6C9JcrJuWWiCU4lRmY+U9jC2suh
sjMPl2tdGDROhCWoUHQNrks9kjn4fedv+OTAtFALe0VVSaLluRsk1YoWZ6RpNPixtu63JShw+s75
N5o992kzoyB1VEEw7qMeTFGgEs7cpMmxv5pyvfIXuEBdbl2dqbGic3ezF7FZnMY3ck3nfSPDRLZv
QrrS2h0eM86QT583cn8gxXVy8Y/HXe+vrGvOjtpW9e3GC9IcVgh3tafetwYwh7fMs7VNAPbYUh1L
w8HalfKt5UTuAmVAYARVIv8WtgaLSRd6FX+QOHIEL+qMwI9//2x8+cXVCxW98CxVXzi+1qFJWwdW
wX0l2te1MNT/+uWYBq2jrwRBsHPupOUWdKqbjxscbxxCEbbeIIsXo5NVsNYcd6GHB33C2CQLIwxU
wvYaBlFbABYCelFNyhxWZXWX5suLBMJtRL35qSTq12VUggyyXxqg87MSl39E7Jx3yMcvUg/8RsGu
H0JsFy96Ismk0Kdu8k6IPm6NXgkgrtfsN0sIfy3uG9eWDLvC1ol/CgZ0ixJIyBX2Wzr5rx7UDlC+
AARO2LxrkjqFKkApnZBfP+1eo7Ia93N8RSMahBpMuXB1hfQk/WhnFnsUUdiUl9Npm6Dx/1YeceQR
s53Ktw9uF3dqSOMgLP3iyfPdCoM0Tk7ja7rv6VvKW898fptLoZ39FvwX/342hBaOS1PBRCKeiS/y
rsgTxsZ456H6SqQ0/2T0ESDdk35I07qB+m44JRSKPnAA9ewx1+X7K1uRyBshljhhvOt+qcMxSvPA
Ni0rT6rhJ2r3aguNe73lT9I4i9IpSnhDkEE74+HMlhV0S8XoWFRcOnaOoLWZtP1vWqorKMxuFljT
BpbTDb921iO9pcYHSq4gNzH7SuzRmTqGwPDZN5UzVJjiofMXGk9og2fY0IGftkkMUzzMUZ0xwvUs
e6oBeRQ8OGSxqhoH/TdixY0fR5/uIeI6n/uyFUiyeARjp5mJw6h/W4UvXi3t8EISWsI3SLVEiGv0
NyjeUEmzJV+n/HJcDz5zuiA7DriLIO3FHVFc460NO6ZJ7DrcShTF0VDX6/N/3ORDDo5H9xzuJDOE
GG/8UY8Hx+h9um1aflZg9J25JwK8z/fi9cSfThMkbsFmm6k5GaG2nKfHnRyefcmURtiOWCVj380v
7uMuRrzV9xZ6njSRb7g3+1dp1aFBMVKXiO5qunBCRaNA0ybHsAdrc67Q1RF4DsPepEclmLMQnU/9
bSEc1zPsw7BkW0zLqeC8TQ8bFR5YEPJRjVfefR1M6Amo4THI8e9aSPuEnP2VtBd+6lnVdXxhAfXt
jZUnlUi1JW7yaMCf5/ynfLGTxLiXMYkH4eYvnjmGYalwjXkd8JS+yYKcq3SezYOvau9gL10W3mF/
jA5wFg9a2/Fl5cZRl/ppntptfd5VK9Y4vXp4MZhE5O1381e3QRHj+u5r+wYXhDAedRINJVjeSTIG
HaJAT7hYuL0HCbtpq6i+y8YBRebBWC6g3Fu1NWzD4NGjDzTiVM1fOQBXDGpKPO81KnHdhwxQGXii
dvdM0/rR7Ea1Pzs7f22EyX3SemW3gDPF3cUPvRLtoc80YKcON4/06sYs1aPW5amrC6l6iZMjViUv
DhZTUHNNudRzfiQWm68ZO88HI1nGz5FFU680xH2yorNZ64obhxRAvwCLy/fy3taidoAZ5ip6UR3p
RNgvf9iAXHrIpNHR3mW6A9BK5a0lRg06riHmbvPOTjBEQeN2/BJN/KYUIlReXnM0EmtVfu+sJ80f
g2UWKfW2p2/hz2jgxdEXzr5HiEWWWiXCrg807NkTs4HXihM7YBK6Xx6ys5V2qz15rMTZ7Zr/SXYd
EvV+WZfQTAOYwzAIAAa/5soP55vTMsqPhaxxkKLPlutZyNAT+MyIR2H/YpsyOkCpRLDYUs3jIEPP
tuEWSJ0Hl87tbeApy9HJFWn9qn793oUFqO181Z0YfPk3L2DUnWXDekvxb+sFVIV1GJ7YVhKE2ntd
TNV3JwPYYo5GT8Atugpdbonn+1ntp9X3p/FslWlALy08aiqJDUyNiGUqYiaTO1xxUm8sAyfaii/l
lYc/rrQ97N3fv1c+M/CbHg8c4qkGqLZUTrCGTdY7Zgh6YhYNdstHkBq6C/60Sw9QZCumMj90Kmft
9oE93wT1sAt43GwYh5ADhiGxKtGZtczBRVirBLcLcQRpJ8rDsdH9SLie9upFWxkryEFHHmXQboxi
rYX9JnlIxlbZA+YTPBfbuEV4QESM/wXwYa0VBH5pkiBsefFbriJsC9YDAfqT/9zUB+V0SfNAXe9m
keB06B3T9dhmATnHRX4h9n05vMTrT4t/YLZSuh4b/ePzIgs+7hSiv4f1tQTj4om5KMIJDyE5AyqT
BDurziAi3ZmV3S3Oumk7pbhZq07CMKg/n0rKG4FXazj3buTE+EJ1/cnM8kbBfsrYJmWt78zTCKGm
Cwh4fzn2yW+I0Bwqr2ITylHwlw6AbBNn8y+cS7c8QUWpfhkI7htGAFI+mCxa33MZ2MKBTdOa4qqA
Pk16mCFTEHxesOuqV5dLHDgqdxPpe7cfWT1KqczPuUYBA45Z2zHIt5h3TP9r5LAI26bwWc9j4nJ/
XeNBcPqZJh/fvG/Hr37L3zSx4CKZ9xzcdwuLbOUL6Xm9PDu5HpKm2XIm7gGAlE5yuqVOvO7e1XcZ
CEdwlLPQfq9VIrd2SvNNVKsdUyUKhkduXkc2FvHvB2hXwm3gcWWDP6NDepPWaM9xUnZ57pynCYLB
mNDEFESSGtljZVgzDG9CHwho0Th9Q7oa6cYc5b+6tw5x6OxoAbS3PDe2PbgKebD1NvKXChQ9PN7Q
CpYmg3KeHHHryRPYKPyDw/iHm16jTE9UmHqCR8ecZn5tO9qk0pyoaPyb4xepDXC77YDJJJVpekol
QYJyfClTiebzNQ+mRIm4H6aTh3A/meaowKtHFlyE1eGne3j9kqBweyMToFNWcC7cL0nUMqkmfyBk
z8XBHZlcvdHTV/igqivMH4Paun99qCuBk3uoZI4pA315+tsv4si5kO0cCn+FtiRtHB94KotffSbE
kHibNCKEEe2M1+MdQrhhFSXhNOs8so7GrxEJMxQSwlLXQJ9FbwWtMtRlOuO9/CDZczCkQP2l/q5G
dZzKjdozxuqdY8gX+AMaLggZUhSBxm+gE2Q8RgG3OHeFBoXQ+ej0tamxKxvm8L4Fej9bPnQ/MQZM
CjutodzRUeDc9sP9DmN+6wZ557gPKZgXMV/pq0G2++fkPE37gaPsEgjslZ7UNFkC1rJ0Wo1PmcaU
DVRGow6gTu+HEzL6t9wIM07V9cm6+ek0FfIJpm+y/x755H4YNytUoPg/3J+Nn/EYqgsuQx/qOJyP
veloVTnBrFpKTE7+X6O4AgyMBKZERZZxF482vxBqqs34ycWbKItFzPD4B6JGODKXVvH6DzCsdWuA
Ch0yg+0hFeW2aHkFDpGg3zClDfoxN7wvtXpTVrx5bgEUdRwrL2hd6+gi0UZBLefQ/co8OUrLyFsd
D8atw7rz8en41dlzM53agW6R3x6PE5gkj9Bqog9QusSqp2qC8lOjddL+X8Gc00DO8OhqHqYQHlzH
Byznblf/q8BqhKDIJLVP7t61UWOrkHOdE96+oXZOrYXWMkjMLF2uozl6Ab5uxsST3g6C5aataC3B
GglP85Zho1F8W2uzFU0UlXMkoZSLN3No2gti4Vo/1lxwceQEdpIGm++ZIU92jaHKkHFkAjFurg4j
OHOgnDqFaZaxPvGOy47XpGg0xbuRHAxSCtk52UoI93ns4I259JSar7jxO3K/FJGc2k+9s/2MvXQn
9D50hwOfaZkY8CmN9H5DUh/Xw8tDixhEjzL40FffzJHo/0skADOw9X0Fk852DCoqsoP14v/n437H
QbkG0Dncvrd/UN8fvFtZc4jedUX9e1uCFfaD2iYOM9PYLw8IQlJDFOvD5y9sdVpqi2sdyCSUut+c
gZBSR6KOig3cdXOBN0YGfw9/6kthSIg2MVpfQB8StONs+kyGwbDW5wfhn7xNhhQ85OeE5aRhPiCI
GW7cfqMihzaKR3na7lom70X3pJ5k9KP2wGg1u8Qre+huhvaj4omqDt0wVawWjVJLVZUpG/tDqv66
/xr3W1012SyyYcMTQM/O4NOoxwS3ums3Hg3znXA5yLDH+vcFYsZmESXJb+sn2pBoHjOkJ1/0szRe
nZIxVqLCc/mX6pPxjZemqFfOrYrV9SfcKQot2+y8YCXrIYg9DgYULN91UPOMyu0H4hbLV1JvvP11
5qI35y6O+bCvQMMWOJ949aaSpfiw0HNu5dsGFymrijswmIqzIW2vve45tIfOEXyBTyR/E/6PTPzi
lA/CNbmGStkcFy11qFgDWHbia7Il4vcMW+JCpIyVN4mGgwv9RJcksH4xtSCi6TGpqOvQRpcJS2Eb
l8teI05jVUo+2wBVEIhTyn8qMJ/25Wm7xxds44nXG9vwMZYmrPMt/vFLHlZqadCQwhRodGzK5NO9
8lXkD1YnlzS1xn8E1YmLUwSHKVROCmncb36I95znmCEuT99oPNAfw4dcnmYLdBcx3NTe0kt1blBu
92SZb+X+/yXfchiTEtdFOeK7lsnkWAK5FXGcBSz7b5e3upuNGv7ohx26yAJ5C4+weS+DqbsvEK3u
zYgF1mZ7Q3qxkv4QpQxd2Jiv4EqvI4ANkbZg1U6VlNcsTPz4yXJy8cCWy+texwVbRdIvFFRSbEEc
gF9U/yoXJYFxCedZje52VA/OY9s+rxQDDWGwIVxDQOThSmZEyMzPTrTG3sx1pHJm7151BCwJ/uyl
G1bnyFAbYSJxzw1JTjsjkGfs4tET89TPOV8ecXR5NmbTz8yC+XE2AM2wEAjjZyqBpB7C2k7w6ZHu
nGU1AlvEriH9KAjLogQrQBjaq9/ol+jmPoReZ5lH6X0QftuimwhvTBIOnqn8nQdcwISQMFgDDahY
HeJXVPU7wM1DGm31UhyZJFQIuRiRNrOpc/Nn1XcygEufgsDuxSuI6cNWB6dDT9K5WwQkG/V0MEA0
bhZb017DWQ8v9BOx8Ed3MhHkS8noF3YdGY8R+AxNUbBj8G5aln84zhF25fgZ5Mn/heBojKHkuWB8
zfN0JSIro5x2yL6UEiTvV9k6qBBsv3+fMfH13udbXLO/WLu5Heb9vVj7teZTAasnmpBMJ+Yekg9B
ZHfiyxGOcTWccKy3NW1PMa4K6KkBCGbBbfUwVSD9pPolDjmGKxLxfe4+PrY1Dv1Sc9f8I34mfP86
l2n4aV/U5SEoBFCZKeppisMzA9HkNSrjuX1/JxT8cVAwEYCbmNdIQ/QNBURF8c+e4UUTrEjsQgay
y4vwj1w0wo2LQnLRLUz/tBQ89/5oK3G7lFFCdm2QvI5QcF6mcF91dmfGFxjTuWJOuE/zupNtv0W0
bGcHEdEyBR+ohYO+9kw0GY8Ead9rFZdXjg3goQQjpBJJtvKcpTjjaPO8VYBmUSJm2t+Kp9CJZyaz
Md9sjhnYisI9KAcrxQi6Cn54hVxOUKcDcpcXIxJxSNxOFxjPZ9n5T5cA23v7b16BK+gmAdA+wVbT
OLen8OVS5XsBoLTgWtB2gB1c43rgnjSSKq73NN2LCOSF1CU1A7A5gZzsPv06Y21ZHkDMELgglFKt
2k2ZwE9NstAN9fsY8H4QsjpnBZpDb1jinx0TvXP26/dCbs5vDJ7lsDy4fLqOnRE7tvYMP926bdKF
IO8H009LSbsK4iq7eSKOi+fzw6T04nNF2u12VYOIPjohxvc+fNvDj3jpQVQvzzH8OpxnWOrPBFKA
7ElvsFIR3WipPzbcXinIy8laNM2sivpRRHAfUXEwzh23xRUHSba/kCFuK2Vz+an5/bPk3n1wKWzv
QDp9daCrqE5Gx34Wn4SdjgMttb9ZGM9MUrgydPu4uMvIEY0wYebhqPuRvRluj9t/dEeHwIJwPQJF
E0rJNYaiFOijFf/Cs1lGfXpaebkDqnBouRP7pbav6EyKCZZ78B/ltLpl370kFOpRrJtV06IWOWXm
wXpOJWbnNDfLp5obaFnSz+ZlFQiuuGm/0OBfNVvZflawGp3UdHNf+vW01DBjIfrUR+tf2O73ES0V
1qmjAguahEU4DjLL1R2eDxHsCzn2d65jVM1Gsr8eQia3MyrqKfpVTz1hjMHSBakNcA9haxnLoUAX
kxVAMLhyinn7ZWsBLlojiufClwv9xjCR9mkSejfWOpUx21FiE12HaL8Z1rp0nqo9kXJyAvlXCJ2a
xVor9qW3NmwoXkYJgpGhQJCuPOAkeZLJkIkv6qReMw3Pb6aHld4QrR3EZH6M9DXLWAgCy//Z7TQN
6ELXJd+9oASOihUWXLcZkWhGuLdXnsTwT0Av22FfFTlS0grSjHrxFewuZ5GsvbMSjDgBVSVNCsIN
3UDlBmP6/JChLPCUV04dpKs0+Rw+etxbPzZ/5md3hPL+VTA301wf1H6d2Io8XWTJApFgYSe6Fx53
hoNRVDH81ttG9afq8Hd+MQRpshVnDyRm4wVykKs9HeHSXgs8DVKLDU9BfN99atLfHVLfZMMZgPlG
KgRW4tYBQ6WbWtVhB5QR9XtND444RuaMzqQOGdPXAD98rAjcpIEqAb82nyC+/WcUHUbvDHVMH42X
ML+TZvQAAJCpGebxO1Y/SJ/+40EQ38RQc2Pd3hs6vIkODTKAjHcxped4mekVsWG6+3mFx1N8T7Jy
v4JCDVJ66jaK9iDousoisLCdyVglA3MKU9RS18Wx0l4r4vDGcUQ69i3sjXh8KkIhRTEAk5dxfsF8
ED2gHdkBf3tgWmJ1YBH/QUwnk34h2rZabcqdjMePWeTKKX7fKOAlL2UcqfuC67i3mB2P5vnCtKWj
HbzF9feO3BP23ZiMITZ/t94ZN6bWvBxsMzi+Dsn6rqaDtR/e3NzgNfwB4xx5Y1KU8Uj+BBH2zp4Z
YyEnYvkMI5w0ms4unV/kO44nJFkVLNyeircHDptslUIGbUIqQp62k5c2meAzMexSabYpfDes70Kn
qvYtGhI+WeQ+qyuq602ln9NfzdQ36ybl9ajMs3DgyFRcQfO4NcCst6un7vrmZQ5cYgMu1ZheuNDy
p6LYQaQCiFblZ762rsYfDjU/nMcBctGM023BUqOULqAByUdyJMMKVdHtx1wEoe0A4jlsOLMZlkXu
CUaImtPMV1QWzF1UphYWK0WhfiepC+ghb1oYP5Do3cU29F8NduevoyRHz6db5fh9IuLpcssQx8WG
vb/k6wunAqNNuRYkjyrRWK4kKOvoMTxawOa+IlKAJrdQRelrlM+EXJokaaaNYcRIaY/GZ1PcXCAt
5LMxPv4dk0ysLP+7NpFehaFvelvWLaOKjNOUiB0aXFJzNvCENDp4zLMveJgDaLmEM/bVlQhqydLJ
DUBIYC3IOEg2rk44Djfvdon8cYDatN66ZnIWhVhchhwjLHcxdSkrd7t/RVzdHhbjQCxKkTKSLUWm
GoMaRJn8Sr4aIC2WhybH8VyuMdaIXAealw9zCtfO4y24odQxTTbksESPJKNJjm0MJQpW/wjTSt0p
I+ryaezfODBOkIBSUoSBSjGhtoV1M6a63mTkF8YlwJNVbUByVyN5/9V8UDK+r+IRXoRdxNHRH08q
9c5KuDMjs2KwJTqU8NHlFey37Fk9Df9bH7ytovQu6PL/zQtqFpl0i3HGrkBOnCnW5U5uMlYpTiDA
l2bjuux3g5OzXnD150VdleH1zsOzxZehRn5AKVNFiZeJiVyvg2CgGy6v3fK43enrJn9S1z3bBO0X
vrzsHaxfayzy5b/HEo7oYo//S0jYsZaqa/qu2f8k3EUtE7s8XRlc6BJGG3CNjreYI6Awgrv+1Kqv
/jLe7KM3eooSiU6HCQXeUBK2hB+mULPh9+uji3gHClwwdL3L5VhUHHS/j6ctdqvoG8KIaHjaoIG5
JN07j0rPvmstHoIngRIs65qp17WYf7fgSSB3cYEralimg8VBpBqWLL1HTAYRQ0JIy6FM/KpDL+qo
SKW2/w9ZpeD4F15lqRLsSRcnjn7E8gNPpQ36ZcA9Tpp3rl5Qd7EdnPqJ8BOj0M4AVS7dIf8nkuAk
znROy2Zl4dVOQEUybNOyqd+zbMGe27oJUodv5ag/j2wGSPaMmhQIYMnHxFwUO5tG+Mz4+rhrSshA
EzmeijEbr20VOO6OIJdCuI1zWjivVMxPmceK99CCiKQaON//aioecNExK7ssi35rG/dGldigjam3
n4tVC9aiv8zvztbuK3yfEUyhxwPHhadzMSetNaKIbt51I0CoZOfHtTnTa/fT3n4ITVIvcb5B+DEX
1B3Ywj6QBmt9Fbeq1sRySp6FPEr+cUs05oaYOZy/m5N/MdTKY4N/H+YVLDWX6vsDrf52KKLAkkzB
Zo4I8UFLMAO3OEygdDDNsDxv62pUpocWSLWp1Gid73GvBLEbnL6vFTBvb2rmNnQAc8b8DbCZ73q/
CVzLRqyWvA9CTrKek590GkT3uoaG14grcL2Y467BYZfAvhEscrXv5xJxYMR0b+dmjrPgSxc4GWZx
L57c23nGyucS1OIsrpH9I/j/DgrB223pOe6TVdgqTpB2kQFTIL6r/MtsBKFYHofksDuPiKVve3P+
jG2orXFHg/B41ZTv5sNXcsXzbyRu5TM2+Vj4MzXFjq9ETfG6lOQ6o3F7+80UXegMIDS5DuhTzpD7
6CpXMJM8Vqvp80y8JfpeivrNfY2+H+f/wJjN6E5a4ZwVHg8TvAthzjEb1cJwBzOszvK3mF4FZg04
U/KctmjImCXI1LFC5Bw+QGBPcgh4aN4yxh4AOfSCymXS2rKqGow4eFxOpvNzjki6VNReC1Q1Vynr
RAiZsl0ugkX+YIIz8gcHt8Ja2jXXJT9yf1fZ1wVRveyBROygim/p9DvG5BTQs4zZkyR2yJM34KUu
4ZOU6w3e6/gngRXDM4TORacq34uxyJFEM+6RYJJvjV00ZWD0liwM33QDlwoxxAjlj43UseCdwdHF
ycs+DLONctI+RRyW9bKLhpn9wMa8uqP6K+Euw8tGw015s4rbZi49ISvo0PkhG8Goqpj4XcrXRQJ/
bCR2Nz+rdnT18biDawKq4bXWfsMtrhMYo005jN/+iZ6yrC+fMUHSu5UBwx8FMGAFZbrWX70gJgIn
pGStbu+OCLv9MtRIXuTPu/4qGO7l3AAU9t40apG6gdxsfftMQhoRXwvgUJRn4mAwdU2tZc1wBM0Z
MV9vemgolOG8WaAaqSGPG1/PTsectwkgKm0PRie9w34Hmo4Fr+a6sG7FU7lWrUa+Mg9VpvVvGRe3
v0zXCMvlOlANel4CqsH7edP180YrpRrKIlQs1k8idcz+I5StwsiaKgGPbAKHizX11wXPJ7rijaFA
NShgz2udbxmG1KgKgAkMEG6N0eti2cVvGcjq4HLRNDm/wXITemCxIecaJfnzA+RA9HmrPiCqGxSB
tc3VyOm7fOAHz+zwpDhCdscHWw7kj4FWZlB09ltOxLnngbTQsBgCgQErVVd5mtpWnvdHzZuAbzWl
xfrZ9Yvf+Q92+vGtHUahM/WPP00DHupu0TuxehKmBhUrebBW3yoiMGXGvougB+EYpWQfcYnQ/9+2
j3FyNaq4so4KSvFreGOv0JIPCAF22owFDJsbwoHqpIxaEX+exVBomrK5Onn/Abndic8yO+8brTtc
d961xKhby+7E5BeVDgwZSacBH/4wBzLKeyfL1wiXjtMSdjzdaucKGW23dyk6GnC1EOyxl7v6aSHx
L9CUamH+ZheyN2mQ/yJ1bGIA9lYoyhJN/mdUM2uGnALbvm1nUuN0+MPNPKnhDd/txp6hP2JvXSyL
jRp+S6dtJF0Si96EBkwSYpbsP6t8fNK9RhpNScTZHntni5tZIH0ARIWdfAN3AR9pGGyN5RMYrkgo
RoVUuPcIGn2tdtcX0+Z0CkYo8AGfn1Di6ZMUYh//dugpETPVtilqIlzoDX74ckKY64hVZ8A0Dg/d
VFdCcvfj20qlM1gZca85qXusXDZO6bpBOVLyzytoomA7PHrDUUwRpQloT24AZQTfWPbXcq8xslRA
xe3hDrRli6vJoXUgr3g0gILXnpLAVxYA6NgBIqTCpz1F66szup1PTPmHZIuFYgAFQ32/5Sb7NzyO
67qIsWrgb9C8j2ZVsSTqOHAjfmZNXGcko/0RBRvXH9qYYdgyHaW4Z7rm/Gjh5p02GSpjZi8xFODh
2AV8WPOtC98p8Dv1s8ZOLz9R2ZnTMynhMO2bx65G6/XnEGKkZtpM/TFb657bO98pvkIYMtJZD4cQ
1lwRHO1KSCt33Y3yrn3Te4p+99xn3OvyPzIy8mDp0LQBgbgJyLeKztUdRN8xQddnWjTwf7XAdmPN
DRUMrJkNAt97NGEgXuxGTXjZzCZpua7+2x4KOd4Fj6q6AH7TpWwij+5cBIWVO+ZIEXtVrjRmmOEV
wIpOUC5z9rbPGKTyqYu/5onAvnPqVq7xKhkpGIr6DLYwKJ6wjFlkmKshoJA9TuRsayEuJQNZnwHC
90a5W8L+zn/SF9FmAAbUSqpc5VY59fdB6OWRzXUpZZrpO0o7NigG5wnQ7e/bs8PuWwXYHM4vAjUJ
MYtI8787teWQOj7W4DpzSOaq4meuGFKp8UE/4x/Xl5reFVoBPuTGd80XIdAjwp+rsXnyctae31km
HE/o8cSUOmE+kj8ziarFJ51MCulY3C49Fw+2n1UtKHV3UYr91am3tfwWRonQj4hMAXb5+7kmCdIe
SgYGmnZcpUjNJXRTIzFGewQTE35Ql1yIoBPLtx8MfCPldUne5IFYWEwvK87fln118D4NIjU5qLLa
5tFuSr8uUSvciHHAyrUuPcMiu4/Rge6nbmzxMLfAPm2StmMi2F1UWY/HE01jX6Lx/fVgZ+mnW9hE
RBfANh1sRVbtZi6mV/ZE0tgM1Vg1IBd66Kjakj9Dy2K/WrYQxxHsWkIWgVNXlOCxieiWLRP66EW6
JEM9HJGq50EFuGPlolpJT+nUTD29uA3zpCV+FGeALthwAiuAhEp7Z1CLGOZlbkvubWljwdBnMAzJ
6vGWdkA+WrF0jKQYaHtFt16wscafXzzbn3wWDOfQOBSWL4xS2Qm1O0tweD2GhWPI4H1loms/lIt4
PoH31YhUjW8w4QgzBnvMRWZhmxGwsskAiU/ot2y4Kn5sqlWzo1lLcmN27MNFqMUFJssYLGuprf6q
Mk4yezneyqn4m3yZH0V2bKpOw9atU1fybO3aZSZhXYcjnjxXUY78HxxsjPyz329paUtC9+dDwHxn
cTF8fLciMXw9nsA5Um5939SoVXuuhJJq9lF5pYgPn4HbghXMdhBXLW6oBa8HyfCvr+17dsFwbULF
hj+En3OjgL3kqCIPZRz8UncxsCuTV4mH/g0u/KPG9FFd5SiuJBT7tBTg+jX5hufhsRXjteA/2tAN
U8DBfUHh7y5+ZTjwEMx7MleKxQPjcdj14GvSCzBQtHtLyvoONoJfmyvlovxoXku1MgNa1l1ghot4
361iwsRu4vXOGCMYNdIuvym3ccUQ5mm6Rbr5hIGaWv1RWnUnxNy3SSMuI1ChFJ5G9DaCmIHaNNYY
iBwhxd7xZwzuhrSzu7TL3FRffflxq2BNt4zPkHfzkIWzfxGlovYxnxiXNGXMg8U54mIBWRrSq///
SG/MB07PKqaS5+ovLtnLXucDwFZ61V4PTZxLJoQpkLYI8QPg1HE4NAjT8gt9/E4vUc4Tv7+NZUI+
cUtGNwStBVeq2jlvpZ/HjUHjq1RnQzpZQXusx33Rv0W7NpC1WAIqADAtI7HNmlKj8JAow0l0T2fq
i9mHFaYi2G1R1/IiUiVcIWxs5djL/FDA80XrAXkrtciza9U8SmIe33PNWaL3fKyYsxz4eHncRxcd
tgG6DmTYMc1P5aZiiKN8GI+LlDPjVRMr4Xbf2owaYLfSNPb9rNYEfcR87hX0uXqHUaqz+q+eHPzH
Eniv0dhVaRWSQOgQuXkcSqaloy5+3IU/Z/jPazBMdb943qvuqgTbG112RDavbcRTYkP5dqRKmUl3
VvU064ThsIog1MYLc7dJ9as+R+ideu0yhDKx7kejP6+sQ+equ/xviFzYsNYtVBYQHhG4Jk8yxReo
/finfZH9xHLfqCwqJYsXgL/W45XitoaDLQvvTyCCZFZbLmLgQrLJKx63lZP49WpLRANhhtoYT3Rj
GPYqHEwbyyHth2oB14rvMkwI6f+2Doozs4k1PSbX3a7iE7XrvBOR+DK38MUVA3EYtZp4yxuGamJS
uh4wc8ZoQO/N/8s4jZIkwi8h8KNilJOD9T5uX9S3gOuKPdgFd1+ZtJezRg3Q9dRhBebbrXME7+eV
LmsspnQ7otgXosDUU1bSDpr8mmW1CAotO/X76uUb89HyuXZYDZtWNv7gTnD6rbzEZvYRmExeOzmY
aIIgjHNYyZO9GCyeBtCeWYsgBBv/tamGibSDE0xv2Hv2nKepF6MYVVP/E4C8su8CwYY6uZWtp4Fw
Gd4tBvW5YtHIA+ekDuDcrnfB16/oTIypcULK3SLeWktQWP82Sx/pLIkM6DPT7srzVSgO0/UAZg+b
yfBWMQQS2uUdYM634Nbrn8SvS2m5bsbqch43+hmYGT6uAKnnAlaMkHuSQ/UTvPxuP3+zBE2yPP6Y
p/t9oEk+8GF0vt28k1/CDrMMIghKvov5pOO+yCUqBxaXc6/RCM1uy8wyTIZSGVA7rLMdO24RJ2fr
xoYwQM1hwNbSetouLfzZrrEFPg6ww958xjAqtkJ2qA87PTEWXRYAiWayO19oLSur8qBC4mLPQmw6
scS41zJWk0DsXtvzWn6AS2+/c0XAr7Y/14ObBNL+46URBaPrXYcwGiefISuTuxBt4Kte4O8lwjx2
fKejcDg5b9R0+XRZaPgwtb0a8yrG4GbNBJxOheXdzvwRqCi7tuIT5kksT3b7HFd/yC7l9F9DEhjf
A089TsULp6Ycm1du1B/SPhQN/NneDPEYdggcCse4K/TdQ6suBv40tNP2E0glGnSIntObUYT8KpRo
IOVs/vvFsQV8kUPeGeHCzIZWvSGmIFb8E6LzUjpsGZdVaWLwaP3dku29SpsnFd9nrG1hRlr612BH
SivssiSJnQJsaNMYGq7chYamJMSRsVuR745585Kcv7nAQI8VKZWeZSaBlk5rZJPHuC4h1y/N2EEJ
QnDhFX2dexItnPMX7Vbv14NpVGkJL6yxsG/r7Qml1J4GuaDFlkd9NOJ2YKRsdVAcQtiGlKrjcD+T
6TimE3XU1LuRXDrit8Tae8GPIhm13eH2jw2n9OKNTp0Q46DoEJl/y+dqczNdjfiCx16M7oD3uxDT
xiudgEL+vyTF7HUOSL1ZACqvHChHo25fokviRyqdF+VVclVigYr5KtveaKyImHi4k2EHyiVhvLFj
XJtlmO6VBEFhLPDDsiGp+zugK50IRzyfAysnwhpbfxG3fXIbxtPbVF++0dAXXFVwU8kDLaFhLx2Y
Nt9pip4s8NwrB/0hv+TDfsgALGXWDobeY9N31stdyVEpRrlh+UJVZF7Ls6IH7q+I2lJYu91CPXY9
XLw6FJlIOiIPNSu4jLoC+DIM6j54fF5yv9etNYjXs2+4bmQ5L4NSzH5jHx9BKfApMGcN8xMGbSAQ
+tsunWj8QD1lU8cKKtUTMACghboxEQJRiIZ6DWzDusX3CySNtvW1eQjBV1ZH+AAWGQOIiO+nAPmj
SSfuuW/uP7EOUdwUPinUGBiJ9Ux+nGBZkNzfDpG75urzIZSmrkahG8IW2MFpDosf1J7jKznAmkNQ
lnJR2Varr4qt9pWQ6WFVLtrNoV1Yk+A61nHI+eMcmCpv4xhydTUL5kXNu0ZfjyWJ5pJrGOC5OXtC
j1nYizkmAkEhnET+4X+LWvPk5UoE434IokSNQpC6W16gvKOjHpkxfmOSXrm92yvsYhjSdfm4YNzE
gRwgVCObgWz41vHFbok+hVJD1vzKUrNh0K3U9h6q//laymkblqvZoXEqO7ozkeLDTA89B+Chx/C9
JdujXdgh6UmzHu2dIMrp/DeMVZX+MKORbIJr//cV9cv74OPNscsgJGcMWLh8hW02UXYcw+f7nqR9
4AB4tSc38DRR1UkGAOfcwEJWUapdGkuZd6l1Q0NguCgiOjqHTMTtyDCeDrS9qAmqGE5hEIk7ZUC7
ljANIthNIs30uxbK5GGtPSJA/osZPjyvuqIQtP7k2LVtOGzOI4RrA4CAzEhmcxDupiK354bVj35T
JRLm8u2rrjZqj8qpGof35cMZJpEHt4HXiQmo9Ki6afY5o7SKJrKHuM8PmBN8mjm4ZW3ihOyTbP7y
omgIEGVQXHqpcsCQ+i/47HPlK2U2x7tMJXgUwjIdygGFagSKzYxDV1b7jfD0hR3NR3/8Dw2eABn0
gampqpgTgiJPwdvH6Pfbg+CcHYKh27nIWirZomRPeC3Z71ukz45rG290K6jGh+MC5zJtUGANS+6b
UAmaF0DG4fAAJcgpZ58Sx02xc8PP/ZxuxrTjRrWLK9w9dSK8Rx1d8fKldwfRTkLsZIfJBEBBWFOI
4elEUsRGgfPcVbpMa9C3GFwOzsgXw7VtIF9Rn9RZEMrtRK/wkcgX2P85DR09uFIIA6zpgd8p4ym8
p4AtDCU0ixxpBckPyQRkaIF3ut2Ic02P6BWrk3v2/YRmFwpLvJO+VWge3QlplAB98h0vrcHw1X64
y6vH5RxaNd7dAu3tEmMgooFr+shZkgvB6Msq8xPnxhHkESBBGR6yW9FXOTrAAcXvqVwuK6Hytw4P
+SWNeq/o22xM9l/Z9bEsHlbFbP2TzwGYvPYHO67WR1+taIfYATzY67nKvJHP32QOeJyoTC7v7iS1
lCUcTmv3TweZdLSVfR/OvhmEWZdZf8OKtX8yX/7Zy3FdDb1EiTEalDeh0399XuluXZpmzGCxrmN1
FchAJmWCujtxwin0jNmbSIOQVL1HB3rWmwFPN+dHEig3biHIEoZ+HOdhwVKhfvECoZOU2uRjB1F1
K/XSRU4hT4x63k0g+zndktIy3yN+CQmGN8MYBDLKBOrTkRWRPM1YndvF6HVhuLyyvFeMSDNCUmZF
Q8S3ArTarmYMun3yoUulP5lwVjFqT2rmmCTS4zm2ZohvTFA7D0/hApag+h8v2EFKT0fmEqnTr2cR
O70XDvQpDPEgN9EHAW9U/Ti0ZqSp1b31Jpfm/p2J4+DndKcqbfdNaxdLH8s1nnCuuPYnKlEIwF+8
+i9+s+dL9PSxob0G1katcTwltNnkg5RyasTtlvyYouW2xa0QE6Ri/qDYWHt/z1hyTT2367FyO7Uc
Js1rC2bZBrrVE6lgQyqes2C3t/nE+ILEz18XiNbqRpXBePytZQjvN+xAjsM9yDM9k7LFkDw7lAwh
LGu2/5dpewCmToRSYruMJBFV7Opc/phDk9KLZC68ppaFfxfAvhjx74P0mTRtPEwuti4/PdUjvzjD
Gyr/52MIb8FC3gE7VSzSzOwrPy/enzFIqSSc7R5DDa+zamdtAkMdMSXMaM564D5CHQvgzHkw7kG+
cXNP1NT7MmvWmCq9Jo+MaD3AHYbOgmig6huokry2s2Ha5FHaIm36USiuIVxd8Sw3TIeZKAAQ1XLg
k0aSpP6GiS3plmk1f9sd8FYxLl/1D2CR55SYD2d1sdZSAP25OxoYiBkT4/nudl2OaeQykQ1JSdaj
h08BDHzx1LDlxoFp2ZhkEhkxnDvjySh4Kty2XJpznGxLfP3K+vgegFAZ/F3+lcW4nZ4MobDLRmo8
ksRvXCgbi347PxoDA3Loylh3KQyNuFCPszQYtlTT/Rad4OnUUp8rzoWzI3mM1UbY4HWT1ubE/8Qs
cbyvncl+/tdjB+S0wbOkaswEKuI2zXTrWzLAsqr+tjnamKrtTG52GpjQHhVcn71wHHGvJIu7THdF
ugRRGmEKynXMOzMEl4sYfyuW4VBHdTd/E9ibBIJzApf0nH8gugm/76GsMFqJP6smRmmmm8VWB+vd
7SPglo/pSes6Zzvfj2mpTh/4yNW2NJfDXpi+2Rvl8nhGa+yxyA4TcRptONAbkvYIvSFXqC8bA3MV
tKUCZktIM0Y+7LfG4aI8vfhQWqrkRVhdr+W5ZVdxx1vLwEOCSCBJSNwnYKOcYUfD80Gu/lo5VDiI
NWKzboWg6tFmgByvPt+uhI/l2KlecaguNHoPPay+BZxq5FTmL9e5X7GaM5vPOXYlJsaDsmMQUtUA
VkKXoaBTy4TheYHlW+AXYKyRgBNoSbulfJothoM1bJFqahjlUIboJx3d9czz5tqtD4bMRKGGEYCt
Q9u25GbEfUVbSud/H+ub5urWrN94Wr5rsQkYV7bo75IH70OzuNn4LSjzihL88mE2erP1SW/6MF7Z
ygsBGkhSfU9pK0xBk5b/OFi8naqOAAb+uIs8IkH2C2+3ifVM8/tg94AZ4GwK5QzYdOileI+9pxCf
hoa0nq2b/Jxrt+1s4pNpz0tTAKFS/Mz2L7OmPHaQ6MtBpkoxJtpPKMorIO0KR+Ul8pvWNNNiaAbI
8shBjgTEwtUc/p0ZWA/AcaAzvJz/j8/XsI6GRY2RQ4nnV6RSvTc50p8U9reLA0YVJS8BF/UBY/hw
E56IEv303UWhtuAbsm27rJ53sSyF+qKtDW5APc7KCYc6hQ98Cm90L0m1bSWaMEbdljE4UtEjog62
duTJZxeVit7DKfo5ceLQK3JoXcHoy2i4+H8lbkbLR5Zgu/OsV7jmWVRa6y/zftCgarOBufVxXBC5
H/Xq5ObFysibEqcUwrhOscRXHmYXDsVjRNSRAOhNIlLiZhNvpwC9v3gCb0ivgBqagUYk2yIWnYd4
xYpb0tT2uHF/EuU5U+uvFJR2FM7aupsRiEAOMxCqVB73Td2QflrieeeSRs5a2Xy8ZPiVVAdsbDyz
idfwEd1wmzOmwi3K6eqUexMt4TQA88/5uHVSk5yvxDPxdtXspxRWh9NhyV5Mm4q9/zT2EXPrvpKb
KPNwk4tZmVAqEPdZz3xl+RsDzZTStqPamNzMOCzY3cfPQekxt4l1cyfiahcfKSeIjG47u/1wGapR
OpNj30MG6ifzGo+ObUsnhecbxPTjzp3+AGEoXFWSFOPj///xZ0cXah425MXGX4CES+zWZszdQOl/
TqQaP/0yH2n6zJxo0CiswZ8g13NMC1HMKnM7IbEbeL4kkObjx/pNNPE+wDsc82kHprK39ARisi7s
ZqpbC7scsUx0wDf59mpJsimHx9buyyXGVipoQL+gk/AKQB6TLKNnq/XDDf5CtaD4j59Qp1GGm8dx
PgsEk6rBHt5RLV29q4410hxvoUD8HkJql7B4BvXIcnnDhmUli+jtEZ8MjXRJClk7kgci+5FQfPQ/
RGzGnLYDtOA0HzyJSQ86FprKEOkgpy8b+o+FHSs+pdHOuZyvd5p88Ev+BzOizna+OxnsHYA+SIZD
dm7YFYklOIE+Oj/KCo3BvbY8qr+LU4sQrYF8ov0YA44tJCdWzQV44/wtS/q2nRpn+M73LfCM4k8D
hQEPM8oX7pxX7kK+lZjXLqC98r/e8KS+l1hTEwwm3DZF/QbOTYDGZ66k6Gnd+HefCmn2ooI6hQ6P
y26jxHP6+XkOfVwRhripKWcE2Lsz4LT8suOcEDxTaV15811Xr8V13n+Cv2aosBMfitAKbbqyhgvR
zr980PDok+6bsYFhhNubcK+bUGUiyBVurT/5f3FhrWKMd2uKIoRmpA+UQ+tHMlsSIvAG74fExXof
CPguNoV0ipqyeqyavPLg0I4TwIzDcZ9Rba2RkUg+IPIxLxx1w0h0D6cui4PLc5cceFqc8WdqblSo
g2FQekNHxtBnYXc6C1AzP/6pM1aY4y1Oa1e9RBZHa1+jmuA6t9Q2SzFz6t2BMKWi0F9V/VPdCX4/
Y9pEXo9u58QR9eWddEgrYkUW3ZH1zipnyohFdvP/AVoFuIIQMuW7Bqe+KUDTqGOv0ImMMG/qLLXn
kv9Zm4hsiewDFnrNcIZrlR2nqTtT0nmbhG6A+bw3h62GCo1Ga7RELWCKpieNMMPo0n2HOXE9NpKA
GehKosvz2tvuijbMK32AqSea7lWZ7gNLpfmWab9z/RA9onOOdbJeGvtGY6Z3ZFKEnwZbplGc4PZp
6iza00qMg94gWfydxYwKgski8qQo6DzjBliyRh/cOmQ5pcojMnq7p6upx9/uqSODK/ymiQSVZkjV
n0+O0/GA6rjdwVTLSPlVxaWP4JF5LWpG1cI0mhAZCYsPsUGMUVRIqlubR0jnyGYFQFB1c/GPbbv/
gyATHTL31e5aTaiSsMqpZQimvYnnRzaKCH88DdkxJC7U5v2vUjXo+ozTi2bxLZiTd0mF21oQsd0g
NIixBXig/FGgcRg3dhjnKlo2rGNmmaCfnUG/Y64uJxTKjIHCyWjDgawVKKkyVqZwegaUdAWrDUm3
+FyD+LiFTmffvaFrW4EkQjJhD2QQGRPXmtg+lkbwGA4ts+zowzsJl8gMWtkA3/oL2mb6x/RD9CDE
36Ph0EplCZiMKyqHHvousM0t/qRFvJ8NNjST6FWTNNyFarN8q5bBwCPBzBPfX19lKBqXY4HOSDuG
raqJaGF6MS1l69rYSBzSLSyT0TF3j8929Nw4bEn56ycTPCwhr8DQtxVHUbMxzAd7ENZBKKjWOsVT
AWCgo8KFeecAP3gfvwTHfJnZWmbGxoZwJiJwlKMWhJUb5vLmCHWijVTmH9pjEW5p6uuQNqsMtynE
2ZHezFhIJRdADK+Bb72Zhzy4xWlKRNrzrEgvdjrtWNZ9ON0X1vi2KYFFTpZdRVWaMPl6Vlc3TOXq
P/KpCalGGVsTHe0QqVHBNtLPDgjq72o/i408fWDB+ml5LamO6hlmnpgV3UuoNtsg9dbwPzEV7/16
ScvAeDZANJIzmzwkDGlwyrjl07xrNj6+YVuWm1NiA8O9wRgnVIz/MZRdFVwYmaiQaeg2l5y8Mliv
cIWvu5Adwi0qC/wLa1FhqpRggctuN/9/E1j/AeMccqINorY5lmbs+1M4N4wT29jSplCCUnle/J6c
du6/DnJ3iJpAJj7Pwim/3lj3XFTAaMTXBL+s0GM/KonTeJtb/57rvAtWUQZQHQ8nc0y98XX8c+Vv
jl15py3neahZ68rXUA0WzXt80VEaRR64q5r4OeSoI9GEETMLkyUzw4IFs1u1p/Mq+GPBxW8a+PnB
S3vsK7WtcgwKDGt1DITVT7QXzhAQ07tBaW49Ym5DSlnARM1az7ScNMt4cFpRY+mPVbDy4ADWYdsI
H1xD0I3LB+vgSfRKXCcgSJ6EOl9UUxqchwv8DbAxQ0aMNnLLq03S4PL7FsQXkifnQ74ZCl9gsEL5
N9ADoGqzchwsp0KOMhXx8/eSL3RuqFYgP26Tno8TH7NxLMYm0UF9rLaH57aBEshIgB7GYWpAyHVY
Yp6i39hhczSimy+W3KuXceGDFRnDRjJGWYu/5FUwwAGMDTiJZIXVmnVV0ISnzBEA8Pl9iBsF1VPe
BxiuI167UeLg02HkVAfDt5i9WTAZMj8o7xgeci0n4A3WcgTm615pZVe2c+uTvjGTGouCkFH9PKf6
qLFvj11m/iquuASCA6CRZRta2TF2Wuw94s4UtXa7VZ7YDjO+OdbmVHAIXRrrYyYCermAmjZW6mxU
TP+NdCqoTrmnEYBW0mgPo56tHBPbdegopN5cN+0UhC2A07gMfJaQHO8FW6ydpwBuGVi9WO0PcXtd
p2Eus+JIOJkDsfEBzi5H7v6yEMDWxsU8YByP6gnDR7U5u0oC/4gi0lHF1q1BO1gYR/mrptj9MWlX
w9MsquxXt21RKzcgtCwuqp8d3znfYXHpy+So0ECVDppsF0vSjXp9MjvAN3E6mQaYJ/2QZIdMrflL
QIPl/MNW2Boa/cWQLa2pUoGM0GQmHeINqWopPWehpkBOSZOv0mF/U7o48UdqK76nbCSHYRnbV6Uv
Q+p5o6GRcbz67MFzKjpQ8YLRghilhlUBhXyaOQ4i3Mo30HWGqBRLrwG0mrNRFP9pLAAEboQV56c4
N7cb7KdB85xYOv5RFD7vjdKbfe5Nq5G8SYTiD2FkIWQAVTHyCUY9SNpYbNZhWgPdoY+9Ina52Der
9d6Yf8NPUUBIfStsKOspcncO1GFqf+IUg2eLO7B3A+vPmlGRQnHRlmM3GKXrjDx0FSNajR/YNnSs
zpIYiQNmWHD408ng4unbsHZA6Ff1oej+JsZ+ZvlESgNm7RSNid0DD7co/vR7N5WFLjoAQdKYmxDw
4LHXJ5Ulo5RNscUQP46HBD9Y7J+fksfd2mbjpC5ye+tIvHDFZCEW79dr0m4fHvgORuSZwos84lCl
xAHVmFV1rdeoQrWroj37D16hlDCRT2ONBAqxUK8ffR53jdy4GvZw+5J/90NjaHCmbRVxd8eU3va7
L0JN+lOHu3P0FjmpuV8fe7Yd4qzjHIrqUetgt1gqWpsgxaZ+111GoZaCmtekl+df3BvtFyxhpJWs
nvfPz7HnrR6cYanU7pxLX5kGEN8KCi/8G8ZSNnfl+B0bmwtq117Rq1S6Da0mLSEFKbvVP+GwttWr
NDQcKwl+DLzgoApWmKNZ2XVR/ea6mMHCyuBYDtajQ6XtvZkZeLk2lPLM029BcnsKIJUk0yPggJk2
mU+Eot/+8RNTHp6LxED9h0jSdjfRk3SILLcjxtUPN2HQb1kLjlRVJWlxteo674B490bNad4SHQ+i
gnbrXM2MeX5vuo/+0+Bv8UPX3FcjBQpUpXu4ILTgpgbC7VlxkuazwkOoZHv3SsJMx2gYZ5BrTF/Z
XCQyhgr/PR5OQB2+B7+GhfQ26vJ//+mocKpgZ1lHY+bKXJ+315PDdSVvR7QdNBZN6Vfzb0sr6/Oq
kYJxt0R3hVUOMpPy9OjKDeUanDbwrcQ9rZHWXph8JXidsNp5nviX9N8XXCCUCvgNXuhDB+HKj/Bx
Jtj7fFr6xFuSc+IBnKxl7rGpZBVFYxf4SeMvbfv2kUuO1AUl/DwPeyp6GUVch9AHrv4IbHVD4DKC
pg8lkwlgoVDPBPVzUZV6CXUODdLU92lAyHlN4LWf5kSE80kPm07saLh0oblMGJONC8M+28QKDyiT
AECNC5NzsyhFHqGbgz3LB4NBgadRLqxiFSlk4bE/isA0UGUHtQYTdFpwkuKXhBOgbbxTK9WhOn1n
sbREg7JUPbCsYkTkamrwith1ej1bGu12ddinJ7OHMBPS68RGExZrNU3Rdvr4A8eWm6UM0cB9dP2T
NkZGGKW9eIaFB7IzZTnzHQWu3FQXzk4dHc09AGIuNRRZJV0xPeFqnX09rk9jUQjP8pG7sqmrZbLO
5U80GxCztkD2VDRDS5YjNpg3CHvhQkb6T0mifx3eBvVns+1ZS3IruT8Z/DrpV9KZs/IoxDQ8Gh2N
c8afJgK5317zlaetMNVfTQ+lyFhv9RDrwW4yw/lHGZyfcVRRawLHE0e59MMHHPYLnXZTfaJuL3dg
Yl3T7TRG3jZgY0Gbal7d72fikn4Fc0s/Les0obVcGnAratNjmHMMMAqmemKgjqpTy7H5NhSsvcc6
WBJ4HUzThpH4FhWMX+Kwp2lVB8lhhzWrCe8ul3a+kbsId3AV7lfEzoN3wYbYJq0z3PpQ9zF8hEl1
hRu5rC4Q2G5iKFDHzo9fDRCQFsp4dO9ho+JHpHp2r9BRLe4/Ik4cwJInEpjD1wIURoUUDydH1H5b
AMS0DNgGSw9al16PXoWiLtehs9++w+prCxnCZDLG5hnNZfhYDjnZLjss2TaQnndwoWqfKsjX6EOr
hvLL0hTKlEiI9GEyWckVprau/yH1pA0pQSqfWUVjBwsbyhJ9KTBF0tqQCYCkYc+sT+xJ+zttBDVF
toEO6/B3qNey5d72vzc0kP2x/xtlnf9Y8k3njPEUF4/3cp1K/B4CMSkKpQ5kpbohUm7I9SgCOBXt
eSKy64RvCBPGZEjMjiWXnXTkKZfSnv6RtmPNec5FcKip14UvDEvZU2sqXpR/bKhQElDx6mevEoz6
vdMA05Pl5878PvvGOeIrd8ej9r0LtjOzbb+HzbneqWfh8vdBO/Kl71PZRP9kzcZifMNlgkVL+H8U
hICECk/lJ8aBhEbzUfcTWr+xS1LiphA1rABgADhoSStutSQsFt3Yi7yHkQR2Ker1ffd6ETu6XIZ5
IaPtifh560q2rfcMmQdC5FOa/q5xhfZFerZJPxqsVTfbG8pWU9ao+tzy3lBfPnd3jR6WaxsDePjD
0g6ZsL6KaXUpgwn8ycnSlKfeFOJ6q50pOmh1F1/6xu8vajJpaohRjdykFcuNb7YU1GN+Jmp2Mcl+
IfG/qJi9TUQFhbFnF1W03o+eTOhALEXo1Fhh5bxA6qmYnrDbyLWFb0/rKpajgqyKjn993wN7l9JF
cGk3cpJwx2Y6fNOokIQ8+b4O7X4VC6XqhL9q57HhbGNpO6pPWg6/rob0B+o8DJcSJIL8Cmqt8+BT
1NGbOqnXYGDjQc9ZYjGFEg+escILj5TmPiPOi62b8VGyM+RQLuRvFJuCIHRU6T0ZL1qZ4HaAvrOa
CNxwFl4l8l689Yqo64+UNyD7qxjU0yKiLEQiRHkFA6pCBkSF78id1RVehbMOjj/lgDe41fjuX7g1
1egqBycOjKr67Ag1QLS6CV+WZ/zGSPPstkbhJvv5WLMywJ9299IVbEJCFuUpnHqOAeNlX6vLuSMW
QnEjzohLwrOsm3444MQrXxMTAdgj58eQG3iy66HGbUIi+12ZkGy23Lk/B+uO2hNvlzSh4dSDu8fs
38GYhzhmmA0b/Lkd/vUYGexGNYBelQe54/ForfDSAT2g5ashS4GStYF8PWSqgBtTEOcLekYbKS72
3QdrmLxD8s5CSjJMNDV4P3H1Uu5T8uzyth8rtVLI/uk4KD0NenMxmiG5RaN8/8/YLLhFU/uDy8xR
kt5D52oY0b+oFvTSYuG1x3epGArmPEvGZxtPoPJzPF51xx8ulDb24CxGauthvwW474Z700ZvtyPv
TyVs6SP/hP/h5qWCNOeEBFZBERBRHOhPxVYQeW+tK07HkqEGeahzqTmGsUns5YdlCDd1ElGwttGs
1AJmnLgoHTM1L/V3rmGDb9zf7WU1ftRVTvgCKFXHNjivdq20VSsd0IBuvy8DL5jrWnkkurQpuc/P
cI2T7XaTen5X5HCWaz+fVByZEdFG7E8mV4Bz8GZ7FHpb0fa/8ioVs1AGUPzGP8+5aaXvRasYsUys
2L4mWnnRhitTZ+R05dScmf5TAQf1fcFYzmX13EI5O4TRvT7l/l3ZacFj+idkZKXtzr3Qeo+tBXI8
Gqxhk8jmiY8mjH80/OiyxmB6fADirlPk9LFdwR0gNNZjT2/ry/VeAcIp6zdVteo2xnZ4iILRYUPw
HQfS7gYd9M59SMMN3V2A8zc1MBC0SSgH9PePQ9cp7v0FKSfx/ExhO02FhJvXtWAyooV5ARP0G2wW
YD6PV92HZ7gLYWE3lphoWFOvqQybyqmiLoYrloIFRvXv3ULN215WBdaNPPQPEtbev0kWUM7UT06d
++7e6TzPadJHjuWJGRIU/OUdzrUMul3oUTSehJfhrJHivMHgwEcLKgX7RnWox+CQIDOQbzPy2a8s
30V9l5FfPSbh7XmLw79T6aDI2CRRcVZUNYiYlqBmS92mavfi3/x6h0KP49oP4yQQWghAtrlrciby
Itu0V6NUWP4hhi7MR4qQdSqFkF76sJwPIP5kfoCwafDxnmRi84YB6uBEr5U7eiJ2HLV5ZAyD8XSK
N2vDROCmmnNSGmQUBQ90DsIryL04HkwD+0S9BlT4bBP78wI8TNRZg4lByS2B3hTDBU+YdH5DQz3Q
qicYv1JiMgImuOukuRYUckCM8SV8RaeE5HZ4Nl7INrOolNC+mV3VYdhWvYZHbyaLFPU07YHQu0Fa
z3mC0kG5W9ZdcnIQTXCKf1QtSQbjrTYFIzLS0UD7Y3RJ7BEFxrPD+o42VDRTyXOmkni0xMfQ1bPu
ZaMbLU4BdI59Bu5l4FLAPD5StzHxXc3XwDhUEhrF/ETS5OYCnyL87/S9TM2wLDdkdUcoxPdTVzOT
154oALGaHU/7iqTP7j245BtqGRFoZF9c4hUo0T9HH0kGCooly4eZ2JF7lumJgLLhjAYV0+M2Hr9f
zfDhdItwtvGUW2XDpW7tiBn3Rm3Jhl0faMPIT5xrJv1vF6RNgDz+h8HEc5lqOoq8jzpu54dVdd1Q
08JZycd7B5v/ZkTqVOrS3BSQK5f7eQPtzs9m6H1Hv1meZ/M8/lWUYMNA5lL4/QXzgF/LFSKtk/I+
DjxyuE9aQiWghnj9XsMPla+Y74vczESWE8rflv0KvXH1JC5BcR3eWOm02KT+zHC/Snq3D9D1cEj4
fyfBpY/M3cy+DiTVqyErcdljmgqXAILyOKvqrKlBUOEBOFmC/LxSfIegrzu/ssfN3N7lIeY1Srwd
BEhGGoD9hAgSBcAfDalelH6vAFOa7yjO1pKuo1goLDVqBcWA2GQ9LKH5UHo39osiJF3J6okNeMp0
EMqnI7uDiTfspypqN1yTKZuw4k3fasSHjlm1PCOUw7Nw06ZMZn8NHbk+hPBnIXXj9AAk35woBMaH
QjzhnDgTyNE58Idn8oYuDGMJRgTM9R39ssKadvPCW8fNu0ptYqZ67R/nLfE6ybgXr8D+KarBhr4C
0RHFM5lkxzY0z6U9ZNcB3PpR2MAmSZwzw3ilTw44RVAcSIYR62m7qv1FSEHmqSbaK27tkFW1H8yA
8HLfGlzfpk+nkgmcj0c20TnxhPYfuAwT7ZJSHtiYiqLu5cZdXfSACy/4/UDxD4zT54VGi2rszXiB
6ejRBDn2kxhgiuPUAq4LCGyAY+nZxkspy8sbm2he+s507Uq7JoIK0Q61WcVE6NH5zo5xv4iNTo/E
dFnTxIJQrksqITh9AaiqSr5i3QPCXAWTHbRHkw4v6aqjJHYJ0+CgtqKevrnWndBH1BoIheGoxgj2
4HQvEDu+6FfBEAl4l1ZAVFK6atODKYHKEdokhBIhpk9Qvh9IKOJuRyqTGW7fO+UghjK+jN0CGq+n
LNlSA5we7tJcepH7nQZdh1La+mMyChaQFXaWyuBgfRkrLPVYDDcdxeFSwKbYU0jr3jULVAoQXNSt
7Fvq17+KzOZf0fokC1hgSD6qM2Tngyo7vLoW3023inCLM2IpTR5v9XntQai0l+CpYk+0EJ7iD7vP
8a76dtaKA3XiVJHtD+/hIdoxROI/axXjjL1YrpfK3U6hv9mQxkWOitQYgZy3M/Okhos4eznIYeDM
AB1cO1b7QNZ3CbeIhHcGYOiSAx2upHVxdJzPOPuXD+5xT4MoR0QZ5p93diHAHa7jDCzJ5+fQAwoY
fqMIYUmLFwYu3zy9hI/BXNl/mPWlclKDJ/vJITdR/Sl7KZm17Jzqnag9/o1wZLS4wRKKxzczXFUd
a5NUAmXuSCV4icZMjMiW7EJ9eMnvxhc9ZyxQj0V0JJsrmLCbDoP7xjRtiMC88ixAKm+r2Y1xGihg
cHjXbWq7uSwA54zMirfSSXJ/T/JwzzXhTghZV67a2dyfqMdBub/d/+PF5ctWwsNQH3bob6vWX5Lv
fw+YXOC+yXYxRuafQI4k4tHzBS5YkHYrT8CcW3zLwDbluSNpn3QoQSXBTDHLby9s7Qbo58hrpFra
lA/S2QqYhO5Gk5lRvRp3PMEzmkWG6IrzHxPJL4iP4FDD2JS2Z2A6rzxUoOOjki9nvaiRdwUfImdh
UTpDIaygT88HxN0O1qKxlekgZiGToAP1qVgVBYBO0gEbTwqmcenHYpnWr9XrkumYIxmd5FBRtXWK
N3dVBck5kWY3UNIYLegATCYnb+P5L6w7ogvcysBqcBFqC8kYpy9F+yrXZe3fU3DM1M9XdO9ZPzx0
A5gtOdnfQP0l5e+CbgVHD/gRxygYFssXidoe0XNOZPRqOkhEWZVq3bdNGpVbdUBUSW/QjmWMovfJ
Iswh0EV02Da2JQNJW/9h72Opm8E/JlKsKeH8/UMCtDyNTSAfL4H1Jy6qlKqD6BzvcLa235Hwdpoi
BgDEwdHrFbOcxXAkwTQZHGpcjriYYZoNHDXn/FW+stfuVKH0yPf9R6lTAgygq3w1ngG3QV6w5wdL
mMc1xWW7ac9cyEFqgdZj06hIpXO5Wt3fS0p+/k/5K6dG4IM3dZ9DJFstScPPuv80wDpaENEuVEIC
QrXVGcCxxIOWWWofAxgnHpP/NwHxw0MwQzigN/ly7CJOmw5+XZ81fEODrgwtO4byE8vjD5iGGHkf
B1VE5VNL0+du9We+btKPhnpDtm9DGSoSQK8zOTCqoIDBSsDZa94lhUUUnqE7qZ9OmGau4Yjk3koC
bcvshG3lTi/hxLdj0M75Svp9YiC60zw419U29A1t7o3DIY6LY49f9EQBK9KnNxqMSc/ir4z7EcAO
p90YYbBt5hdklL5VlsEwQBGwKVeQkzMasLZFDlOYFN8oWlHjAx2mZ13Nr+ZWWiQFgKLdh34jJ4mp
af22ljPhKFBIfUqGpcNXfx3G/nzJ0/mUqTxBwdvR3jN5bD+zBvlF1G39+TYg0KRlQHiHTZsNKJBk
kepBzzHBS+kmKPmPcYMv3wfuRg31qmWuAEbtoRlMz3uNanrzI62apPubaEBHvYHLPp9Jxgp1bXR5
WslsKMHBO0MF1TCyYAQmKoYw1cRNBRbqW+awRlaemPW30OWAjkmuE1lc/hyjcJkwjbcvWYLv/kyL
vmzF8dvS5i4L+1X0bQEtvQnsC0ecCv0y8ZZ/E+3C5Lnf0PHQB2gUOLWmX3FNNhmOhjalwIdIP67J
rh6umF00/xqAFGQMP4n2Jc4CqFOP/Fvvhd/m0G2SSEzyjFVzi+EKuVsAicrF2ItDD1gEBNBQA7Jt
myUqlxVO4cniEILtSd5gqgI3PUYOzw+kH3zb+IJILj1I1aS9R9HM1GQsrRX8nE7lnRsoja9ngX2I
DAW8MP7eu1MN0hkx8cJkz+c5aaQd1ak+BBXvaJIvrhmpznzXlzDjY+D0SV9ON6MZfwO70klhL7tK
t+/BnCEY7R7teHIeSZIPIqJ8hfIK+NUQD3cAfXjA7R3Wb0d7cHnplQDlX5nETkOs/spc3wNuSc7K
JWw5l7DrTBVQ6VjIFcK665XSBK1PXJqq5ewAJCePWOkh2irPiFBHIIiW4aFZ4Su4SDiuLNQnuS8Q
DYsWvneAlpRehm6UHUmlJIDqvSi+fGf4wgRfQ0xUTUdTpZ7q8rJAMa9sLlYSfCXAk/TFNrHndomU
6K1kWIos6heMcnVvCY/KD/W2oXG/zVypOWvmMj+/2ZkUxEeTwVyeUpQJwDbvCJi61Z3olcBsIqFA
VcvJPgYxeIJadtVDXNeFRdsOWalol7sihbwwCxwpK5Exy8tt3IDO374ctrNnIrvCRwOQKfPDpD5u
zaDmkO8EV3MVg8A3c2w8FQMWRTiXMUeGjjhBj0TEEHbaaayAMxS/O0z///TjLuHntQRpbP+sB9y0
VBdFqSAaQhXEMGttBY5gpqhNKA8zqFxzfb75kypCPfff+/xKsdsUaJCaP9xyNRw7tUud6oB8wJRk
gH6YL5MrmFXoydXRy1Rg/neTgoT13cRcEzYSSkLjuhzyk2hkMEAoO+fHvBHRzTiKYGrqRgHa2A79
VL7Pw9jc55bsB6KfJDloIWldRUuPVNsiBBD2aJWgOW3tPv+vd3Q7UwjD5meKnLXhchNgLjifk9zh
+F8WwMktdAdglMD0Qr92GyIpHrJmxmdePYD+zFTI2EZu1yBL4DcBdZQ/clNAMrJAcEHhvdES3rRM
ALUPYYNUZAaXXg7QQ88Rnc+hlF/206L4vT2alJkys+C4SspQCfc7ALFsT2pW4JV/iyZhMGCSnU5F
KKpZE6vpbxS0xn0ALWLoW4IK0QjKuez5In7zH4eSmtule5iCHcKmv8riL4pe5JPfmNkdHiYANh1U
cH5j7NW23biWclvGGNcaapZ6HgeoSEBbeCLggj4Q7kfxIZs3+DVskbiGD0gS8KYE9IEWqmLKyT70
d+rN0vgS0QR5xkHLoZocDaZCz60Y/RygzOnuqT/2wetoXos3uShX5rkzj5Vit2oPmQaI8AyOLK9M
NNTi7rCQaix7rXSOrmMsHhOypMm1eo4D55Lr3ZF9DZw0sra9jfXPkL5qOopzzVbUJJK1AkcNt8cb
2XB5aBQTNuL9aBVfwvR+M7hibzSS6v+TKMyjZN7VdkzrByhPBPYXr5OHkgDGsAe9cw/2gjAqzW+l
KMDuOeSCo++PThFufTni1gdSVAz4BFfxRTvtepE09FFvujti+5JZiELE1we0iG0w4naEhIctppwh
v1xWic+BJyhINs+cN6Mu8rNX7S7VfCDmsSa/PSP7Xwx9JG9A1xENyqYNkQ3yOXH4DSxhBXE+NbZ6
gbip9UkDqqhjUUDlM6tsQ5uQmCdSsd3B9SHyWE5fVrCfoFSsjLruXhk6DKBt++vPEkduW57nR2Tm
hmMXMmUFYalUjsizQolFm4Own5Ndeiwhge8QicgL0V9vDjbM/hFqQCR0FxKPeqJCIZ9ihe+dWIH1
lEsMudHFfnj+o7NLhLxXXGUticy7HVMF4i5wcOSYqN6OeGXUEgBsvdPeCgki18cJEugeFaxnq4fm
3Mv/IXndqsZcYbSvKx24//txYiPCs38mS6yik6dILq4qpUU2jo+fOAqnL/yDRlFzAIyMqvMvTGog
fu2dWkBW8r1RNcQKDSRMnk0jWkhYpwPjx4MMlyBpwD1OIAHm0RGlScAa4zDfjoRMZeeAMNXIHt7r
dI1Et7EM4KlkLgk//rRO4pFR+p6jc8oSlVUQEAw3cxin8FLyeWCfCPSx22hWaqtlQdgY4BrotzRc
joiW/7rsKp+hoGpbYTlMHcZ5YFeNZSlmb2JZWUOaz7YysfA+RRfE0+EhBpgvZK8SjAOujexyfE+K
jQxbyLiYgSk+xZRRdRrlAOWg7pD2Pm90DZNkgeUyOo38m6KerRQ8Nmybxb6MDYJe55ci/ScvUHAQ
3TsZc4gMDiFPy8bDrMbFY/kptio4ablwncgKhK3mEictqt6l5UQRgndv0OU2rvUISSk9KHKLpWV7
wlfPw4HBX4EpoGpQGwRqXCwUccxPJKACDvwcUqfypwKcK0LKzFsNUWQdomVLMeD6I+2pJgWgNZLs
VLNn/o7fQwUkwSyEgmN1oj8iTVFXwfvpKX77xriH8g83JWAKWMlQP24O3GyWlB9bZh474AWsrhw4
w1HAPcdgwE3oT3wCjMnx2tp9OFCEHDQKYPilHzSPXKUirR8wVLj+FB1kYK5Jdnd0ATVOIcv907ks
qcF8C3Hro8rOt4edaiPA5CLU79S4Y0ly+NJmrQjrUgueQHGRsF1PJ3I1RoojjMvX7r366a/z8Efr
s/RKAv9Iui7Psv8v2wt5LUe29PC8dd+bQCuAbq4rccqfseHnaN+sALM7U2/z5Enu4E3WZVojPsF9
7Rnaz731qR8x49fIE4vc5T2CNLO043OOTgTfsd90rImlUMeqZGwMCrwa8OUVW+3IoZlFAKm0oytU
gYRpGXZNgHknGy+NnMMhxUB4ZesXFhAgU5+F5C2iIK1ceaTJ5OjC5T3g7s8J2hYwcAyYTyqprLNs
MByEfejRm+FhHh5gxxU2XJsEE8Gr+Sky3OvlMieRgt+jR5FA2vHDXkXXVNBVj/E7pH5lLodVJsvP
prp4o87zM77tCZcLXKIaajnVrTionHjh+djwV91jMmTDEsBwRi0Pt9vizno0hVSBtvYwpzFNwBvY
mDZA0iILFVPBw01bXH/SVb8KM+tPxgH4WF9DLmvsPhQz/o8VTAg4VCtXpzNoTiqPCGomfEYVl608
CoN1UY0H4P4ZAq/zaPZFklXTkM4LPaCHG4TwA32TkSANwsarh1uLK3GhvvdQDqAJKp/tYUnzH8FT
hUr3Oc07P314ExtIBSsMBPcohdTLxc183YvfMXUKYn950FepAXXQt25Fpt1uZuHaLqJ2Tej6O1c/
UsegCkRhHn1HL89UMF+R9WmbHkEfX7XIDngTBvavXqyUq9VmZky7nq7kO6eo6Bw2mNx8qHXEnKVY
0NTkFMeEjVqXktk/MqDbjqGGZWD8HTWV1PRlCkY0dkdCLA15Uu4DMzsutIicpA2WCwu/GkHWf7+R
rRGtG3XVOqsvSCw9jgfluqK+WLj9SewmWg4aP8kSP6PWUUufKBp4Zcihcn/KnsKImNlQUCah4Ij3
8pP8T5ftp4P2dHlV7MVvtErfCPoo0ipXQOsneHIQxog0cxcWM9GC1fnL43G6O6xuf49kdgN18/VC
y8iOQ6/HDX4hklxES0yJftgpNjQhpEWCWQmI7nKDJqNvfxEbvHcZ7H5JD7KXs0EfOuPTb6o1Ifbg
XbcX11twzsihujC4ZzW5bzbS7C/wb7x76adTSZy7jDmmttbspk8Mu0v5gzEBHsdt1YfQAgEDubhT
CiPUi6qlHcMWEzmMNKeU7hsLD37eF8NsM3wBSNIs9Xi3/nRV/84OuhwAlSzaV4NTdud8Z1xq4KMq
GBbSDGqowijqAgq1xVDl20Yy5VDN8gTfuO2+2aJM76PCXuHZ8yUJ2uakrqwd3OA8ra12qecUDcu1
7Hh4Eq9VXrcKxGVw6cZWEvfYTWER3apayLmnS2D2j5B4CFALSw2LpCYBn8jHXZ+LDx0P6DYzroLS
0YOogcTVVsVvdNea9AWtVUaj2D2fKHQuYuDbX312i25iVyGP24Dcul91e6URDLXNfEJl6+k5wwSh
0ZZTIHJMro4eQN308AAF/C/aq64wDwZqwqb8mRjEpZX7qZcpNU4fpX9s+gqQ9yQYuJuWSscYm/Vs
LMmjDrzO+4GTN5kpNbrBS3KaPD4JbVVAvkSkyKfTLBtBArRjAwZ9OBbI+he272bz7wkJ3JW+4/1l
jTStlkmWMiK6y0LT5ZoP/wweGEkdD1ARAHBYvSVg/rbg/UT0GKIhxQ1L5sILCpQu8F3Xp7B15g4L
RoLYk1QrmXKYXoD6f85DU6DII486fpMAy+NlvMzx0ArESK0BcpOaYjgGuHpPQ0Fw8m/QohvOtptO
X1Mg/OS/kUy4WAr24EeQ7EfbNukriK+imXVdcJ1+T0+RWXu/HA1H4fm7nm48mCm13Kl5VzN5NqFi
iY+DxGB8QhkcnPanGm6jUoXt6MlaXembulEigqYYdYSZorHh0euXowagJrgUywpN41F70uQlXpOW
pTei3fsaUyxQ79nJaXqs4aZBrhU/ch3jCb7ftnak00SySEeS62QJTQaHAE7oX02VIM/ef/tD92tC
m4yQ02gZAg/NWgNGDEHba8wnMF/6MoW7k4xaAwk7aeeyU4id/Nd/nXH3KSuHJ38Xf29g5Nin720Q
HcPvQ0MpZ39Ge1OKy4+iZ/evWGL3D2MkyeSOceyrIquRr4PQ5FgxKYwCOUAbZrnNOf58x4UBIvEd
QmjP8DiCsZcn6TCxpKpiPwSsyhVBEQFn4xzpse0gTuHCcC9RsfXADm88Nrafitc6U34YfV2lvXSB
0VryX84YI09dIY88Qs9oPlkX1I3TCtbam9tQm2/BFEKF8JIo9Sih4rkddVaa190deQXKb78Bw9JH
TuGMk+AJWMFc/36OJ2z9DJ9+3Yg2jZPI37Ccge/yR+0E1HgfdKzUGL0FE4xrSNYnMpSutroi6XsB
WqI1sELVdE07wPsmkjURsBEnhXVP5vh93au2YmvccObiNB4SoE3ZwkfG25lVQN6owncrrlIVWqX7
/XpuEssnVLO7jRcX7R6Xz8ylWUNGNzVfzuH9tm52IBjLrrPMEfUf839Xovck+BWTo1vs7SwC2Iuu
vRHJmjMlMabcQhlguu3Nch1zLh5ioW56R+IdJ+6kbvmwXx0sGzHHX60hmPlTlIXCiMvrvCHjAlD2
pqr7x3EzK8PylMs88bJ/b3z+AA6P1MAewh4A9Vf8MVoMCh7OO+3uTyT/sTTw+dqV6PlDBuyhy6Js
xfzNshcmssxAPJHOPgy+7OrJvj7uGs4LGATiSAj1aF1igXCQHLGFrzNUqUd92CLRneGmfWg3q5Ji
FLMIPwMMzTft6/M8dsbwnfa2bKZv7qNauEpKHMUTUglHwjBKEkOTORboPaLy4v/mVjtsLhNgRcHf
a9BMpdm1bXlhKmGOreo99tCBZl9aVqEVnDfum7BBWFkSePBI4/K2JowljMP2UNjp3rCPwPamEbez
P07l6KfUlZP7HKVl70G+Ev9UdRC0tQIOIV9KFdiUmUvO6yWcEd7h5A1iyRrQYe0v5FF98dMefpaY
GEenH44QQu9le6cRoWzfXDnDuFmFpLOdT5+Pc8PcUu0xv85eBHkIAkKYki9hqQElAtW/61eV6dlO
I1kf2XrouK0hKx7h173NqpA7u0p0cm8v9IEo9yHQtRmseakkxGbhkZMqRB4P+lNwilVcC8sQ2v+J
P5RP2jtS/TMzRavNblWGio2TMyO/9urd95grpIFzASHTZKauD7PFKNY9Dj3GcpC8z0ZMH2DzJUHJ
q0cbZb2fLzDmNjxcNWP8qt6T2LYJHnC7w/Wb/5GZMGocmS++qEflZd0/VYPAmqfkWGjKYyxKQY2q
IbXDxdckB4ebe451y72JIAh6yHG5DWDB1KE5wgfdffEyqcLIXXOcklRiEo6JPAkqNmF5n9kfMzNJ
6C64LPP9o3qUD/ttfFwfvk0kosSn3EOHUiJPEkhQJOINpl8IWJLxyz6LvYR32ec8TzMAHyhzc00K
sq0q7hcSfJqvJC7EzgpDmWBJ+zPaje1Fl773XnYqQLSfvSMimt14NeFUYRVwbeYqT/foYbuZVt1t
VbVRvZ340BihZtNCx9LENNpQW0D4aQhHKvLTILOl2pMtqXtwkioIHh6I8HT3VENz2j9ONnVSltPT
ym9PtmqFnKIQVCWiOx8cQOGAosgPl81KrakK3KGOm6IbFy8KcF+2sJrmrZmyRfY3oHojPi/NqyQx
Oq7M6HZqfG1SK2BrkCbL605Ewt2MP1crpQoXkUWiVsEwThtXKb9eYkm1tQMk/JFVg7oDshkwBAu+
4CIodRCO5od4v87HRlVM/yzBDeNfl3V52dCdXglTyDrXV3vw8ayzN1Zo7fbzCBLKfHP/DNBgDf/n
FE0jmZDBrv5UmcgiH//7/va1bQl+dmxT+Urc1EBVeMtnKrZSPEKabQDBc2HTmyLrKm8vpsL4JQbe
iGBFmR4kVmW/CeBmq7opD56WEkdh5Vn7gTT9EigfGx3LlMOZfE/njTREVCOU9rrhv3N+jyT8lKYq
PngtCSwl1V2Yrhl9wlApCW9GtHSJLh7iVRFdAwVW7f4cx6PO4Doucs6y6/GNlL4pYpV3kmYgme78
ZOorvp1/xvZqjhDtAi4ZUYqI0mG1w/sFhi37z7P62ni9vvyDfsISDr03TJrLwGsxJE3VFUMt78jV
b6m5rXRw7Nd0EtELk8NpHxLh6OoDwI7FQqViuRjpoZL4yf5NgzS+MiuwTANRfwq+phN4NVzGUGLF
l10Siy51xpbfC7YJ+er4iVIZPoO0SJtOJOyHVGDEcI4QQiqbQ3uSl3hacvkcHkwF1WbSHEjGkr1h
lMbhD4EdpyG4P3xuFBIsEBJmKMqKkh58JkmgfcaSgFR5rJMl6oMdmBMvFnBye+MkY/Najn/3RULI
anW8IBaYqVCWjxHqZAA5eUaiNjtuwjZ38/kSUN49ZCcOdKmxRW/SXNsyIAZbwrmsRJzv0HnQKztY
vdsCwPw23hqAVWZsW/r89yxZQoM+B0NtUJp+7tvYzlQB7UixE8Oz3E9ar9vAf3gkjO9q4OHKKoHw
BTZgSHty6S8WVuWZnjFHU8vj/0vF45UO9deVMIiat/4iMO13okhtX/yyUWVRZbuI3OwJj4smlPaU
mCZrVpGPhYf44+1ncDLUldZSdvkbtkgHnNDgQ5giovtcWki7qGsxAxYER9vEf6r0jdbtEaESgdof
SsBjgE48hTdiRv2WK40P/cV2XvY23Zo4EtGzzIsYI6KmdP3eFK6XZi6HfhSSL67szUYGFkYtB0xj
DV7/bMfIzt6NlC+9A55HWJiFyoetkv6EZafo48tYigQ9zJbwF8HHssotB/PHTANLvKBQOF3/vixe
hTqleIvZjyUGOglj9UR+O7em5SzMD3BogVaeI0VnSyMIxt28+hENEtAMu0eJ5g6Nms4rIuaoNfh2
xYkikFuoQzJC5Ab1xgmhQkk5NQCdUoCX/86OQLUEv2Rd2KAdXlvAoAAkKBCsxqV4F/BILaTUtgc2
AuGJ04Z26kdmM6l+Jb82DMEXUq5hgTCFiAcs3N02q0l5iY5HX8kGQGJW7n+g+EosW6egYOKVTcdn
+6zxWhP3gzVL8BV5OAh0MoFgzkUCwmPRhClwmd8JKN1VI2WSEy3gcpT3XMxCtwsf0jkx/Zcn7UKB
qwxpo6hmdJyj+693bUKJsrBEWJdZaOKWTMz4GJ3Z0hGm0WsAPbNEoh1NgEk3cMZZbH5+owdvzCdw
W9K5gMt/zECK1hcoOt87Ya7NBHt+oOzMPIMH67x/TQlK7tS8rHBkk6lQIFoFt425eBojJErLs7ci
xDlUzmLA50KthWPw0UbHkpcxDDIn4Q55UDvW7OW78YL9llfIRPYz9xkQYj/UT7qgP4iJAD4dRRMD
oTXj8uGXn5n7v0kCvYquT57bsJ1mwD+bUYvOLoOx9M+rSBqSnrcQWgo0GvQGIQ5VgIJbMWYjKAt2
pCe+LzZWPRcZlJR3jzdLZwPwG1C3TTEqtDg+wW0qHmgVtZDVKvVjm0hyfFGzuOq95AD97+mWuHeW
kX/MtnELSLsBCbe6VG+UCAvt7BNr5E1pEvnnIEf3pvvL2/YB0dLf3aY4BHmysiQ29HYgPdx3ubuw
xI2oVvRp2QOw6QlGgELJHGQKQYG5Ml/IXHx8xH3tEPOYj0uw2J8cFBSIM3jd1yjgABD+z2dd6Hbv
bX8mtkmoRIMrQKL73LAayBIYlWl+bMMUg+wJckbIp0uaqkAFpN8J0/glLKhSEwf01XuGXtK17y6y
tOcg0qzl/n1V9F5Otc2dVvW7DtjvT/rjfnThxwu1jVuGE1J8obuP08Jkjy7YZCyizW0UVp1c0tIe
6/QiXzSAfO4UPdlpspu+Uxb4kcngm2P21zkZ4iaQok3Ml/fWVS0/QwWthAuV7t9JGb4cwDh1ljXw
9M72YkyE1c3m/0cprrPrMz9DStHobKsEYua2Goo3zL334FvFPV1Rk0dhapP9ksG3zxb4fPgxpIX8
jt3c7CXX+pGjsyYF7D8K7aXP6SQOBVCc6/XShEFrHU1mMVmEtgiiKhrzxmiR08U4D2tePab8wDVv
MXClFSNLsq1ZJ7rkzSnce0PnFeGbXwtNk486u4wrcSDbznEcYfp0GNlX6A7o1kFCP42lthJw8jot
0oWnLHtVIYaZuS8Y1W5C0g0Y4XstTptHxzHuit+7FcM37mIjUJSTFZwDBLQg+NtKOBCSftqACLzs
CqEbE5bylLMEt/kKwGVGu0aqDlrYLcKkoIafUlIJOIZdstU7hzeMfF2E044it1gbJLOIBpeI3PIe
4qv4mYbb4vwGxoYvrrk2k4khV3wp3QA95vpMUssH4NVS98CDFjWZraZUk8Jlon10RvGSNcU84isG
v0BhHSGtBH9SC3vgfTG0d52wo2jFJKS/+/Y/zFg0dTpvx2YqUri/AXFbSgxtqFVCbbg6g2z0vy0g
ORcpL7wylpHEbZzteRQm4rsSVbB8y1ty2qvLnOBuVLvYdftl23uVMhsAi4SLsnfQBNe3jGGGoIRs
SE8Fjjvq7vfxuR/aOAxUF/Ub2ZkNGDE/wVjC+VqP6bWjlaQpRmGEu3Cm3r5A4BxfOj1G4sjcprOk
otP4yF0N0WaePlMuZAtQUk1rfvp7N6l4QtjKkyoiB7QAvGA1WJ6pSCxYw5+5/0WFwVLjbfBd+eq4
URPsOFWqavVMIBbrGrJX96gh+wbPbV6QS2IqbNn7/E1VzsYDYsPFmEI+HqfcyJjEK87XAKgEMv3d
KeQ8joMrMGQ4SMee803gGe9rW/3Jl8ENTVBgAdakAazVlDOB2hCrrBvfqwuJ6GrHHGLMLE7nT7jn
IboaNsSSmbraomhmjIq9vxMHVFPDhE9SF9dCQzox3QqplnAJE461/3AYGzHn9eLfScqmTst/UFs2
Ow0T9GDBTdLBkWNT6dseBUslJhewj+zRLCGfWdNYBKnBWIsDmRubBHRMJ4H+qU0tCHA88eQpM35Y
EsSg+QqCL+ZHjeFdHDvTeE8DeJVAA801EUC74BQqocaRINXgX/G9Kcclo9SZl388408tFeL4uYN8
F1BemyUQqixGBRlDFofhB9Wk7bDUuJ4JhVH6hFyMDswUhvX+dKfCOfnBbalOzjUUt2zLYnDwitAb
KOWNfue2jzmj1Ukm6sn5PrZIoF6E+6N18FmN/Ln8KnnN7kcHkeo7DwmD5kte1USYvhVa1BSAUZu8
2XCEGjWJe/wp79atFNz4g6YRy3LCgIIuB2YGA69WqLjyEKMLqdFnOEC0tmI/VU1EoB6fhNBDnhuS
KNBQ/AxfsM4UiGc31IXa7Rh54lbdKfOUEj1zjPgbyg9BrP7vpOIBZSjXLf+E/6rMGbMbo785UvKb
UddZqy18QQ5BeEAgxe5+7D8CoF0M9UY5FgkFEisnDL1QbwTCvFMuB5sYOx5TSjyHQgc6cWGjeNck
klKZRPDxT3qS3IN/zg8m2I7LXDdmya18sFAPSHOyY5vLQ2ei7rOH/sPu0R4ot/90njP+Ug5n3y/R
NEhx0zg4TE76QhJ2VEydzGVZp5U0wJdm/YYW+ryPOxyUDCYsJzpcXyLx+l2sd9Y4zswk8SsGZEio
eF0D6AONjqFutWk/3u/XrqJZhrhWenJrp2ZM6DsCqkv3cps2EYltCmow/vH4ZH+mmt3Zvlfh+pRr
EXwAq3PqcSPeM2bDqNPv0kryVdsoSQ5gTtpVw2qbqbiEf64LfSF5c1rERDWtJF/u7U4hlXQRGRZW
cvM6FIv1fjwpMo1cSOGXVrTtlhH6pUUeKV8vw3kc5/ZT0+WJjPn2IVIjO44w/htcHP02FZZMnW72
XeY8jCJBLg8F2iLa+cGys8XqQKh5cEiYqnwfMeN0BoNVJmRkMO8iuWgTfsCZl4MFLk+DrwlNWJSZ
7hQPwKDKLfIzcFhcpfIPdCV9GucWUeG5iQkSymNa5DM/e7SAW8jMHFT98A8+4vhsZGucc9yByXV8
mdLa6J8L1m2JZ1Bmnh5krPQGYxgvOSNCuIbEmfVHvqEJE6fKeX5bt/4quePq7TZmlLVytr4nZFbE
5c/KCPeub2eWIfR0F0ZavB1NLhfvLVE375e9pY7Yd2Abg0JtquNKNx0Pe+M6aTmilC9xy03YZ40L
3mfZaZqKjRviCBOkKp1seyc3o2cAKs5oY6ptYFs8MkWgl1Dc+6SUkNgxzzRF10BrrfkQJlsMzBMs
/40dliaAoF99wMpTJDgfc61T0PdysECEWF5Zgd4USS5QDSlBb9et9uVeRgvqIMwpAam4WIoWu+y7
dOJB7TuBYCLWci/bwJ2DD7CAoY+80dru06JoPOrdWbJv4q7reA01pOF+N9RgseFZ89wAhdMx7wXf
2vgLMG3uPA6bME9yJZJkLxtxUqr9JqV4qYokRWbeyPf8vJc2KVNW+KMZpRIEQ06u36W0+DvEnjY/
Fcalz+1fRL7UJKlFj/+UYz9+HKxHwrvKuYVFDKDlVYukkIb+VJ+Bt3spLwTbuZaN74bwNOgnyaeW
IhaRySyN7F26+6YQtYDmGwH/cnvMZ7D3AsziTL825d1xTLYmoaFzXrEZCvbXdRSIdg0HBQH1hUiY
b6phaxs6kbtg6kIsePgRpLbOMemhFu6wUTiSInsC7307GyECckiFdliVkcA+GsKshi7+Dj+sk0Ow
kCELHNPh/KGgJ1K1828PTXXYaugbYtMV3LMxNA2DK3UO/jlfQC4qn2nKeI/L9/dDAQdJXVoJaXc8
PplzqGQ43jdh+XofbooDGdu9jswI/mNQlppAtXBGtKzjoNUMdJMvN3+0N9eqMHydRSdaGriOz3KZ
qIBdtPthoe0U6Ef5YR4eGpskp10vuy6/YR+ouCN3TVTdTEoH9yrabkcxLgxuuLjbCxobJ5CCbmjs
+O6eZxb2TkjDbw6ib+XJwsqy0VkW0QIVykk6LotXX+vrL6GsgJYUpFSXxPZ1m+0bbVm+I7pibnar
Dl0A4UiZFcmuzQ6K6LZQNR3nZ5iYqDPE2pIoDc7hhqDDedK6wB2xs3CGBnCKG2sU0f6gpOVueK6h
xgHjW6h1d9tn96PMXAZFAysXWtIVUXQKw2+M5V3Qt8/s0LCgh9XEmS3xsWJeXUMDpmVSXbE1SCXF
TDw3ulAGRKGgR5HGBc/mqsa1e5gj9Ohh3Q0cFbk7pHl9NOhDahJdYvh4BkbpR6YHm5zsYGgKBLbW
PpjLz8c0cCYrtoLF4GMyXXb9ORJ+FxUcnSPvLe0Epoemo/HuYh55517V1eVSXHs9ihhQd/H5eX8P
pb5XRvbFrN7jdKgT0YbC/CFRPOzx/5W/OXKCt0nZ6rg+4exUNtK+CfRKDOxT0e2g+U+lqSLTnP8r
qpGSq2K2nFaX1BjabVWuBdoEIXmdh5Pvi/QeNjPqZ2Jwg/OPE1gMDD+WF6wgD+y7ryV09+Er6wF7
Cq0v2fA0G+ZNC0AzDuxJfHg03hYHLqGPcQ3JJM15pi536CurLIqZIZsVP2ZPTVgBsdVtkBMgfMBq
ZtyffwMphp6rggYzXl30gDDFEpifnUjD6rXmxBuYLAfuOhzHbgQbxSAjkPnvcdpKid6X+GKG0Ulp
w8+8OTYJ3dyJLschqgUDXcapxErMfojrVjzB/tqK/7KSfdghcFw+iSU9UoXwEB/BC8g5OOvg7/7P
OZ4VEbr5dsdGHj7ep67iJR4xUMaUT/xI0W2OcBLowycrdZ5o8F2tdsxkAaQ7LwTseeBwgg7+ThUZ
PY9MqPnpb4hlwqKO1VR9Hdsuxc8GGLJPGI5gtSm4bh/TDx7FKBurIPJQH5yqGCR4Y1OsZNL9RP3E
DzVBM6AeTNcnApcvLsbBX+/RqM/UFBOY0XwPl+N/zQCsBqE8fAV+pJdL5cgdFjLLO4dwoAlHiZiB
BF6fYRnR7LWRbCVKHKah8Ab/zW3Re24r1R/B6dfIMuVPh8vI9ndR73kAnmUzQKJHdrK/OWUjqWEP
Dp/QsM/W6i+kESWbYebE2Po2FbAcKYhRENrJBG97g8mX53WFfR4F6R7oWRiypw0+uN3sZBfGo2ln
tq/j5O0JYIoBn0fwKRO1s/Jg1R/DPxR4/WC9QB80vQdiQ2RVVgWwNpsNuU7ifjtuJC88bJ44yODk
Mux9bBbsbpeKfZaIJgOFK4kboMxD/07HhehKL0VZMGJDBukLivkR15ZHPSw/iwOYSqghkDnTsbAN
RS03jEcMQJPv1wxUo9lA50E6VZG5Jpaq1TRJP8o5QdxtW3s/4YSCybEsYswA+p11+z1QJYXIA4Ie
eok/qBZGmrIeZb+wayIzrGbASHqWR8LMF4yzf32ptoeV1YVFS+kZpydEmAogHiIAS3bvrFzgu3VB
BGrnszzU9kpDjytj1UtfD79lJcr0AAlGi4aYXPXPldUyVv3ouqqXdOGVxX5FwyUgLXSCcyCnd794
QpVL5PPbUrpZjKN1ybW4gwUlfDYWpmgFY8Dh25uk5ruTPNIODkmKAAY8E2DqHNQavem94VIaatJv
yULfU4pP6Xr3GnakbpTI7J47QsfvPpyfKVSPRdrqKawgqmpu5ZxwI93oEDUsF8grxv0BHAqSGvlb
pHq/z13tTsl07TRoN1iArFGQ5tIXiNhoNHzq3jsop5PWuiKr0VGu/jV+FOnZ3bZb2alqunsdrI59
dL+eRsV68MRag68kAlNAB1QKd4TyoAAyGdY0LQlhwweFIPyJAh08TXvfCEbr93x2IkygFqJqg/Jt
lSNQzWeaXRktWFn0yY5ZmYPF8ZJFc0KY4AhYTp1I3JDatMEpytUGvAqW0/rsogR/LrblYPu3q+qJ
1fgAC5IaZupZUIHTwR4KN67iEPSpm/a5IM4YJIoygDQ7lwfdKvQo4NQoEY8XQd4q9FrmEj4BLtx2
l9HIe1tSqxmlbm7MatM5FabC0uxujF7HXG6QmWSavPKkgu8FJcnlnMZ/LBW9HH/R8NzJeMPchmkM
qNgV63W0M83BSSWUGlZfGgexWhQ+MM6CAsb8JgaXrYobbPJmMV0eNrd8BxlMBYWQ14LY4S5mqwcs
lodJQnFfHDPruzVsNantaCIahP4mv3Q9OGTUmry7mRMu8Iw3pJzJ18Deva8TD4VBvI0i1CyLmBE5
tzeHQL1yjEEbbLPX6jc+ZSh5XJfZRC1RH4s4MFJWNG864oqdasRJA9W8+Dt7blb1anI9mgLczxN+
pCpIWCDpJxmdx6Uz2X3D9TSJoGYFB4Ecil9J4OwMM3LznNFBDtsUxok4tJbXlQVLwLk//P8TTDUV
8ubJgJpKkabrSz10Qz8TMYCkauIfI8Y2m2IFYtvFvU+tUSeI2WrhDTA6f0V6YzL3OKPWyeDdKG9K
u5ncPlqNlBYAA1MlLlQF7NZWx0Q81M4SP6f7x7IHm6LVeG3iZ91JRV6132xDdmBM7usmbPPnzmEG
+qOK8TCaMAqpBYJzoVRM0tCaTgqXvQZZD8qwzSdx1pXFjCR42kKyMOVJWTQ6AcbXLz7S5+soXy5w
3bEP6Hoq+7A/0wLGDOrTDXvtkhlS9eUDPVTMiZHgdwH/soSR2btZLFyl0xUULTGxUp5xFMNsK0RF
Ef5wtN7P99mzKewpzi9NyAN28BmMv+MRnO4E7PMJgdZ7TBfKF9Vq2Ka88ndElBzomVUhXLB1mJ47
1/4juz2exW+gEDAXospOpy8ugEjO6L6EuE6pXc4dcvPibn4lNHtychvaCiK6A6GMeiQssxlJBunv
/EOtoNds8O0llOgTtd8qWaSWksN1MDeKEmGimRwnRj/sXRgQqPDKAfMMpmejRFJ4kV5OHmtOlCcZ
0kAnoeZ9BNuwOLznLdE8kWDHSz+G9oEz8YwDJfm/g0RGMPIqSb1Ftlon8yA9aqNaIWAH2me7Cepf
vaT127gNf7OhbUIFMnV2N/C8zA/PNaLXcpQ9DIlZ8bFRMU0J1fEUrDJgql5uTmxA7vrH4d10Etwr
Dde8cfwDiVtJrZgUt/myrykcb2LQRNEL2bKXRg6MiCKY5ffunE2DtPco9Hoze7c1sdmvDUvb9/Ze
FZBjRH5rREuTviV5ma9tcBx8kccDFo69XfrWExZ/M2ITAMm2yLL7GL6HrnEfhf1T/giR8Hc7YN0v
pih1WIRXsPdzknwHI6F42uwTHRHvLM4IHVftyW2DNe/a8YaJQVI5rah1EyA5BoDDL2wfrjQPCbux
c7DYlxX35D7oFFdbupE5jR62fG9XUFS7lUX3KUrQXWH+ujnKrNH51FxC5GTnwaZL/N2tURtCwrtm
fqu/YKe69izZeoYBrNXNEPubkdTj3eWljKce5QAe3rJVwPpkETgoxqz75n/Sg1pBnHclC/pGBBOA
ZSRxdudMJVvwmgY+aFa/Bk6sim0DcteBlCLBLtF9Y9f8V3nYVo4VZFntfpVXejbrV89WP8VXr2yg
yrSi0MFuWJ0CKrcZQo/D9T+HBqKkrL3Bx76TJtcgutvSrrph+nJ7a42aHdb3/VN+Q39S3mGD0JkS
RvlrYc1Tn0NxE36BXunOvbkycIe003kx7yYqq8hF72sv4yI0j2CvJgTOUWxD9DeW5I9JIMnoLoUq
Q7DbHkMn4uNeHQXPUDtHZgDTBi3mYaAAq3dmqYR3Bd8CSV3M1BEYxTx1ZHo1Yt6q7Z8e1Mne6ieP
nmydknlw4NIvfXOrDs8QdqO/GeBtWAewuI66EQN0LtfyVp2P0tztAufTU6EoTg2NNBlsL2Ye+VVd
fQSF9YLr7xNCdMOuK5rCPvuqIEdGBAZ7ulNyb1JRPv0022WA82ABa5rqgG0JI612u8SShsLVnzZ6
Ct85ioxsC+29S6HITooK/sooCAE9TBzmVIbCBPSizm/cvhcRNvLRSVDa5jr8fTikEMBzYXDsCGag
zqZSVhikcK2Xv5g8kCBdbjxfRWSWRbuMD3u1FpUrTRS2wTRN1zpxxgEI5IyQodeaDcW9ilR/Sp3q
afxEzUzLOFGskJhCUZrx2nMxT4ZK3AUGyy+gxQADghuA51z35cmjuCqUY6HVYQOakhygiaqBjtTo
TJtwn14pmUa2rr0xszQi4Ql8HfEZ7kc4x/HwKRX84abQ/xIlJz6L8KpL4IgZ/qQ+UocplpAtpQaW
z2FV6I1sOGtQt7jGjWolgRByU5iqU2VwekpWy3uib2pfxjC1Ptyp74A60vTbmtY9lQIB/r+XfBSR
9fATvddbDmWkKHVlVBe1/76n4RdsTQAUq+ehKmJiCYn+910L3DKjjOUIOyVuf5W5VfAldxowmoSQ
IcHu9at2Ii4fDHI0N687f6vghEaYORv61EsaOeRy/bL+jFxsoQFf5eG8NqZNVzdO5P8l9CZ6wCFl
iPSkuRo9s1QOxNo3/bjrNNSDkPhkD8QbPQPSghCtxyjNBgLkixW4j0GgnfKUgZV1mwvmU9gvnTPi
7LGh7ZfLpG4grkjamj+vXXtkbYNRk4/ZuusEav4h7lzGrWIpS5trvSw0LeZ0M34uLsDnMnNhPGvH
msGQhyKeniP3y9btjUddNRmfemztBPROan+YU1s+fRs+HSDdStrLHmW+TW4xSzPR8M5eBbfP/hWy
WaOY8rBzoNYGG9Fldo1J36XCAKKFq/M3PpM/0XCMoc+E9CE1+Fw+0wrMs8/9s+GNta3bL+U3vlED
QhSeLCMhPPh/YBfaG6S8+hig+MI11DVm6GoftgP7UIsLzm+ZV8WmR3JiJzfBBo8UEUexXuzXPfYk
ICTTYUH+YztzMiMh7WvcGkRFeFXBTOpKjiiHW+Nr8PF3RfWosLOGsncOtYlK0xn9q2iXj46OKLYG
MuQqG+4ygXlunbXJ63Jb3i7Vc2zTSQpisSXC0pQBK8qbo0u/2trYeJR2RiwOZr/dMA0uVds0TlLW
CqZLlJlsnJz0LrewCuPc3pE6M8FnWilyjqvJ8z3R/thta/IDf7yHXFavZZ2bOs8o2HroFxw/WccL
ioadAQRZ3z0v8OG6KWVIjpDs8Dj631MCRabmnB1trRt4yISiP6k8V0ME9xNb7rigOwZ9vV2oJMPe
aheQBS3rtg9e5oIMx4QZ6XEFX6PLKcECYMaI3mSrgjm2d2ZxK88Z3POUqkxkS0Mc7zw9socESTo+
anj/M0doFhNX0x7CdDbpXksPMOZlZZuZH7fnXE1GF6hWK7Uq4GaxW+IrPj1IQVc+cSLYdiDD5HNw
DKrwFFzx5ooNQO5IMFdRKX8R+schQoDnj04R6puPGPbJE99Mhje7ZC2HHgXo+tMMcnxJBBhh3geQ
+c7ZZPt7opouk/oJDqd6O3tUPgwQ7RbaEq+eP3OwV1+VNVHDlqTzWa1ia1nXbnq/IUM6Nt/d4r2p
9LrFp7PEPzdl+e5S2TJyy4t5TXdDWiMnMgqd8SH7YCfWYxSIlcZjifeCB6Qyd0tsApqS/D7uGJ79
X+9O7jjjCaoJJEFbrrjmhgq3YUWWZj40fug/RhI2pNOve+x0qnQ/uEJdjHxhit+eIlFOZgmZPE6e
qzCYSMzrne/a5f7xRrT1WueIQf2JkDJfdd/cNaH9bN+ZxaPq6lDJfNVl2x7egQYpOOmx9pTuva8+
Lj59sYtVZxClLDliQQg3pXT99bjrTvEd0/mpHAa/E1NnWiOrA71T/whvMWU7XtBKNvtTmo85lIzN
kD4mrb00g7mavYmI307PtnMuUuDKyQ4JzAjpQy/YmDY9V7vHFZoifAipQJJUGA727QYY7HwGi/ol
mraPuLA/l61nrRaO1II17CpolZIOzlwCYTxG4HxGQlTH63ABtfkA04wcdyHVgcBH3OrEtCgCkMdB
0Ei1mosoZzu7VRgU9p1CYicJ6UvGbiYmgi4jyeaSGkFYjCtzN+RnokdjWAjBClTazZiMjKQ07Muo
1ikCsSUTuZC6wbqzWtvTaufb2C8IDs+05yqNlPOJemXT3r2/zt9T3vG6eJZnnpKQSBVvkFBXsW8v
GTzcTtb3SFWg8NJB715NkcRut1glj0oMN9o0BC7OLKbIQW1aY5XqBP254i4qjU6ptJNOqkXTrJDI
QR7tg5Fkl0kxWJd3zE287Pjqaam9GW1S8hFyI9Dj1ZuGAcGbRMOj4WMVV0d2OiY/muAb6uFA+HDO
jrE4mA2Vp1CTHM3EHtrLL9XYCNuoXNRfv7hO/L8MzW6ig0gDoclhBbhzf22y7naGnsZqOpm3yF2Y
KrAgBxVHy3kzz/g3oMBkzYzGkiy2XcbHu84x0PgJ+V3HZ5pP0uxpr2X2f+moaMe2sxAk4Lh9rRxn
xe+lev+Zfw+NaL91htl4koKMHuKJjrJtGnNAeOzX51eifN3nFIkMaEfSfd9X3N3199dt2Jrw/l1P
Mk3GrQXWI6Vkwk18Apg1VFCOsFNEonmvAC5rkXXL+crgB2Jy8hYhd4vFAtI++5wmjKcAEG2Jd46m
QslbbgtrGW/hZbz4w4qmbfjTy1Q7AqxiGYF0w775UeG8znqRteVCxnF7C6HsfKObRPcv5lr88F0B
iFkRqUK+ertGZhc+HCaxp50UIrLW4vL3Xr1tIydXIQ+IHM8g1vT417Te9yXXhqZeUWzoOGYMsi7C
H8ksVtDJFkj+btFfK1XC9e6im5mR6UflwqevNUmfYx9Kd4QMBY1bCUtxfJGCdQAdkZSti6lLCWuB
sXGp25+1hde8nhO0Kclc/LwHPbqqlDThQu+OOOUOmYerrU4HwVDrDwxn1Nze9YdOutgi0YB2FjaV
txyO6SgCt2kLukoomoOL57SYIAljO+/zbu1B4XWtCQoOoqE6zTwM4MK1qa0kRfp2LXPITae8pjBi
gJdqNjYxHeOeNlJZ4oFk+J1zA7Uh94rRxKfxl1jTD2kGH1yNY/63l6kOU1oqwIQAbMfz/omMTi7L
Yc2D2xb2tCAyG4QlHhaZeiTOJOX+JszHeJMv6gIH3gLL8p3DLneRW1RxvqHQFr+xWnrAvJC2kIbY
iyWhh5U1fBHoQ2m8og8w6uXyP03bjr/yUeqg/2wookBod/52aOlqx6cLQZZ4SnDp3Rr4hs3+ViXW
gsunzsp0JAw0HRnhXeHVCN4uLopQW/3kbU9d+W0oyE1HYP855Zp/OZw6DLqaouUyIoO53fCtbg2r
dUpp0PJ7uoUN3k56jUCgUolHPWMLbR4KZx39D22IP78vuRBAHQCQBM6O5C3CPeij5KQ0z5NcrWPg
TPUd9CNk9Y/rJv1BD5S1E9Hsu6PdfoJYqXZw36Ph9W8O6ruKEF8NoPeRIUEYRQ7whcvPYlxgfnhs
DuWm93bCUU92lsdHCmflpeZ6ITvlx48V18cwyrH3lYOc4ljaFgfuM2PO4yRILu8J0UwD2lQXSqBe
6kRpC2TUwbsbTky3wkmqWIy1yNe05y7r4xZxycS0/6wRvD4TWqEfLbF8yM2KAfM/vf0LzcKTNLfm
RZKsAi1FWLniZ0Ln8S1TOxZInrYkp+3HhkgHOgUb3Hx2+X5GE5SoXc38k+q6EF5hqsYOysbfVI/H
ScCQ4zoILKzALKBM+TMZJM7GD0ta/rvT6XYFuY1eDBkW/j4673mcvD5e0rJ+lDDYZptGUv32sL+A
0O54pA8R5/6JhE5K3gNFa3t4GotzFU7kIfCs1VGI5VsEV7N46hJtGT3UDvEXIqJ6iBe8Z4/OhWmi
EOH3IyyFXnbuOi87Sv1SDfMuQ67ntLNhm4HdcPQdwP6YuioBJLj31xiC53CHzvdR/cEdMxnP0xnK
27aTdRYlp1H2rQCAnScJKodd2stMftVq0/Jy3i77TcRnnoYOSTw0o4vrfSC0SXZgJ6WJf35CvN7x
hLI0WBiSl8D04k3gvyI+8GAdY4FU0KUCqOY48tuS6WfWH2aljjukd01n6p0hjYNIAgu3j+Xxm/F/
LepG0QOEc6lqL0gVTss5V+ZwToLcKk/0u75MjmIQ1Labq7UllwQDNb7/VlXDpFlurXMwZg2Q7hpI
UvvmjK125esTXoXa3lQwHf3sAZSUxNywwtZ3vP0vU1om20sre/bVzcawVVMzUpJGe6uJRaOM8uKO
NSwa8KALx4CfwkzwclGFd5RjhFTkmynD0fO1CvpKZ9V4YxjHTsNj2l2CSAhVqEkbZhoTMcMX05yb
6SvHNrL0EsvbrWOFr0jPJU5orkQXgKE2RtzSDiFAu0kU9KZyE9R4qCw4w2ptuW0vY8bxgt7K0QXU
dgSpt+NQ+JtriY82ImDeMVjsIPwJrBlQPxdsvn5KXWw7mEelsOuDitph6e+iKFOTuyCDkOJ++eOs
rhLGHB2CD8PbudusBBeBdUkC7O8yHM5NsBzP3PI8uTOeSfKOaIfilDiTsjQxywCKLoQ7tdKJKa09
H2w+J38KKs+QWedovjraoQWbyomcAAotxaC/nYoUvwN8K5B4pbuZ5/yAN4NLT4x2KhbJ2F/wMMzc
Gu+gT4aq5QmD7ZBRCOPoFGbS7AGu9jcVZKdRUzkr5X6b3qtK2ZpJYGiozF5uKJe+xbeTd0LQFEeg
nb/ITRauNkoHCQ6RJkZ0aeIbEv16bNUcXw1KYMdbHhYcTgtlQwC/Pugqv7TdQvMXxjF1KHKSFRPr
z34G0xkn7O0QwEmt0GDGLAOTPWBb+1Cw8OshgnEmQem8iYbHkgwKOqhf8mtainTFEZ3yjPF8qQDp
Q9VnrjyRD8/409Vck5JwJNMK40NS0K/mgqYAtRwiHbhQ9wENWD3jbWvbkQMvGoVs0ft4eOJ+Z44P
ZY/V31dNt6tDN4HplCSk89uvcQp5yKGo2I2OHXyuhs3Y7c5SBeYG8V5j+xJZhhwL1quruIgKnKhL
6kB1DYZqam0xOXcLhIm+Ip/9AxS8v0Z6U4MmuzbL6+e/iSRODVbB9h9McHP2IIJAAI2s1M1PR56M
HNs5gH4axHvGEzbCaUYf9UN2tv3E1tbrJk9ggia8xde+8EBy5YJgKePR0pb1AJaksFupIokfxyqQ
axzQT37rhgRdzhrovPabclXNEktBjVxrJLas2aXG6FOhBZKuTySZhm2t9x5bDMckq0tJPboQDl5s
gzzFWmU4OCfgIwtiLGJdYhcxYjRDyOhW7MvxTfAcm5zTKjWGV7Vdw2jsZ9C2dx311fJd4zr0OxTC
DgCUQqbroFkKO8ajA7TPuQV2FtH5yBKgacOkISUsvFnFAmW2a9mWcqZyoM9pG2q8DCawvUNpHk1d
mEOjTgjy1cvYUic+u5PDUjhnAIFPxtw+V2R5bDSMhZalklvQCDPjlWNKeR9nLKZernTy9CzcetQ2
UPPNrJlsfzYN6qxr209sAThkwZx0hUp1lYwqobXcG87gFlzqeflPRCxCpQYjs0B2iNzCDjVi/tBe
V7mKT/oYlXZtcGS1+H9SP+Z6B1vXAxmFifORCRNCpZGD1wVwSC8Fgpe8eJ1XKrk42RM5IEkvKfrY
02VhkSsk++wNzxzso0P7fmR7KIpd37JAdBF5wYBM+FN9nCqQ7S2QvNFwZZXuFIMSDzXF840rdAvP
C7g3Y46qWXu0Lfe2XFBECvgRivxobU+dBcdN+dQxz1TpMcggR50awfPU8ZxJzVhOB4smjNTz2AWV
1XtE361hUHJUFn/h+OGmrR6MggTYNRhYRtuyOwexm2DbpBMM3MAwYX17rHXXQ76PI1gpDLo9W53o
7sJHNJDEpk9hDJOhKVl6ufpAiJRS+vZu6wctYSS1IMnAMiE8uCyV5uZad2swR9Y1qq9Rq4kRw6Qt
jQM2Tem5rzQ3qArZ6jySY96J1esErKGirqoI6DEgKegVHoe/9CIt51WEy4cWjb6MBmgxrtVL3TXX
AL/G3vkcJZcfbCWvnqVHA0Kif0m1dJ1/tV+nWJetpY/aHZMfBa7htCe0VacalE4n/OVTV35w2wPk
cLonC9wwnAQyOBOoAP9UoLnNPFgTS8xfaBiliOR6DtB2y0SLiud0vHncf2UFQmsoyIPrDULhuYWg
3zM7jOPSNIvUY0myjAgREJmVwkbEjGibPy4wnNr0jYcjc0i67zGjLuzIQP/aRSgEaOlfBpI8iyda
0VPYfQS9q6GRkZpqGOGS9/iN1JNakk9IB8AdGJ06kyrU529NjY24hn87PxgbHSkDAIlYjIGdKS56
UmvOEcQtDe3y4i5YTflfvg4X6PSCgwT/ouxB9mSCKTqtzMsNAU1DYqt/YgSeF+UAo8Sb6z/uSovF
DU0TmRAmqso6+wUbBXVvzk6zhSuwP9npvWWfcuhPwwKSRK82Re4vTRHlgGbp5lMPz4vmaisBpaYq
cC+wI9lPzubuedzG5wCFahITeMYgoYvTBc9Z6kGj/5L3wsbeSbBtPY0Mek2dvFJ7tKR0z3rXqieh
hYreN2gOg44mco59hM1dZFqAaaWD3TAFYkw+keUguywqAEzQbV4DGj5MLrjODdpoKtsoVMd+RXuc
DYibPsKYqhdEf4g0sP8DDMRkskgxkbLcCtyOXAezc0YVt98ACSorqZi783TTzqy1kkv1NHO7swTF
Sf0BRk17nPjeKfiwimVKRZfgQsI7910l85YzXv0GLDYynG8f7Agn2exVOxMOQBrUMebihSe9nPze
0RrHKwldMVtFi4onzn+fKP6rqOYfg7TyUgBCz1tLT0QcJdXdyHCpx0ZHRebtppvukshg1ulr0oqW
p5tX25k+vtzNpuYrqhNmoCJ/74cCN+ClqJ3VIB17ziXfw0nJzJgYiWaUJJWNL5ZsrnI2eJC5VeXm
/XGNuXJ4UTjDTZZULImPo5qsAZnOO/pL+AVBOzoEQeB37CaS/O5ziaexeRRyRj4UpSsdypkQLi+e
YGWJYNUiR3CCDqKk7MfFYFAUJiZcqQ7SY49qWRbUmjhXnwjAD4OI6sZz8dnK8bvlS7XzSky0ydqM
NYrhLgvD8XbHoxdOHTDnhaXzByT9SoHoys2b5d/Z4uWgGhHzLBs/+FgOqtLo8Vfhf9YbWSCuqYl0
4K6Nk9x0AN/NfEBPhD4b5y3IiG4Dz8fPDQmHNA5C+GAbNehW4D4CcJSy6QIINKFm9pY2rdw8Hh3s
5Pq/D4zydQ74hItSE47/tw73cjZrlUZt0NqZQmVnTWbQn+oQraezpkX4BmY95ogpt1+FjnqltbNi
nKRjOdnXzHzgIkWqtjjhbMO3y3m+asiSl6QbX85p+t8XPTBrvinOdGFca2X2+hRxbiygUnYD/8aw
Te2roVPWKho0fFTWvvwg9gntTdDfZ1d6SVlF/nzAVqv5G1Vipx8CA+R8w/txbaORt7kthObM+jjy
GhGfyrAHLR10aBtcmNpdgkibaMJ9Mzi/pLoVNviFvvSLeXWqPAF3m104b5jbiHCPLv7uPadnlhu4
rl6AoKjRVQLPoqLDhGteLHJoIc3pVHxszLx4xpdGgLACIvFv0rZrMEhlDsdMNOfeUQJPQxpT61Xy
rGzTbXkdLPwHVqFOuD/0XfvyH3J29+SoC76Ian9BXrgP5AXX3XRTKlH/kxBUKln6QHenJ2ziaF90
BSqP1G2UwML8NcjBbEbUYEVPvU7J2VPT4u3PW3IyBskXBSZpiYtQHB0muKgVU6NKKDisPy+LAYb4
TcTrRhHFPnq+nuUH948FKgWht1yjCKSZOCLyqUjkb8LVeKaZ0RS30cbqSZjBGN3L+c+4ZSEu0nP/
tO2mtM7/mHE73SbdPDyrp9RwW6W11DhpG0ORrLqTcd3DtT19BA0H01IzFs5LQhdG9BJFfMwgNFU2
x29h+IaUhIqHlhaPeCEVm2UBbY74vVeNfQ8ZZniuIvofaoT9kRfJdVEYvQvPd4zHz88WlXh5qA/e
AgqD0m137wHEyD3PXBbbSj5o4WT0xkQBI7d55NH+KW0xP+QEQIbWzeqd+17T4vvu4EuJ0OjUuQAz
jzgaa15eJt0mCH2w4ze+j0GNc2jrqalf2pAgCdCjIlRrFWVvCyOl2wWbkWybEpinJ4Wvr4fdb2U4
aILJX3NUecMJnTVMwY1M9O/B3dECPzXqn28l80Nh4orjihEVblweF+sY8s0KRvE1GGe5BlphiYAJ
bR3AyA3sbYcYymqMsE0q+/t/x741hdgHhylR83z4rjmq/qUfDtOGKAUvqT11PrCsgKsoXb5SYhJp
R/5rYXQUS/MJnGZakeDyIEOEg44C5A3Cck+7K83N0J8nla/CVzdrUk+CuI9BT3Jy2AGZfCn8yGP8
GZO5cVlENIOSjYLOOhhPFHJxk9xiMKX8RqQ8qEViZZNuYSBQWaVaGE6f9uYAakXdyd56gn89narC
LXk66nhMvdUcATLmyQS7Xi6EYQh4i5IvP1COtZLx10u/EEuSboFjA/alfhSIudR8KT6JV6H9wVjH
Awq9mxlOjcGTcURuJD7srW2v377bdz/dPNf3kEIqGQs6D++Iwjv/IJ1h/lB8axyU3VrDdpoOoG5W
XJYgPsb8phoMrTrCtAbZmb9hoeeBH7zELT/593Qv+GlaEoJzuYNlCuubeh86U2pTVIQ7dLFpT9BA
y+9faFOcNk70cHPnhlwEM9F89FiXk+al/H26p8P5LIyf/vb5j+N5B2vJYLN0P5v2hxt1uxdF2nDH
HtF/h7d55c7yXxUBa49x5lM+XPOY67Hl1g5N/KzDX5bfHh+ZTHaSETlctESbMsdeemh9+JfyrNVT
kfq4UkjbSNK7aBeGEEPSrkIUOy0/GrQxE3uB0dMTYzd3z9Mqb8ctGMk8xlU1f9t+GUF3gpA/LV7D
cjiytoKq/0Dq7WFldImpxGbrxUPuOdEVJMTihioosg8QNO72mKlv3ace14dF1JhOPmZNgf3kL+bd
xyxlAI3vnAKaYDmfzqblXAMdxQ+ite8tYwEsLhX5qj5CCX+VOPtfeh1dL/aTGWPuopiY4zNhHfJ0
MMQONCZEJ6Mj0V+k2sFWw80FNJPaNmyKnw9gCdf/NVhQAS9FRjt9pAYccC2QmcnqXg/zz+QRZVRx
MPSJjUimqV18U+B24E5MSUK5wgIsFjRZSccnCei7nywaS1koEC6YRYw/rGbs6VnXWNvNWCi/mRhZ
SHoeJI8k8fLzByKO0UjjBj2ewnbXi6CL1BIPNY1XNNQ1ENOetNjlMAcXp6OCj85dMYxBFBsrUbSR
/woHsxCIWCy85YCXp7EH7tSBIDd0/uz0SG+i78qWMYOeLYURZKtTD3qra1ADVF7KgEFjrB77+xBj
BdTGkMJHV4bo0JssBhjMaaAdcJWva4vM8PxxC73TzQyMqUb33Q0R+DXgO++nybA8LHRJVGxvBaZP
HW0LkviyaSC8BNG3A4QofrJ1ywuyL3fXU/18NXfrIpJEy16vbpvnjHWtkCaTRgSsfmivPttbUEro
OOKyg9i1PUb05lk1ekTN6KLhLjFr8kzbwUfx11LMGY/cfmGukF1h/kcNaAEcLsbYFC5CEkCJ0Aex
4NoPz6Y2+RC8evJR595nhMcmCjInbSREkvxCMgroaB1WzdhZNMghlb6CagnxyNu/lmXKIKlbt50d
baMle6vXZ4Mn0wE29qp5/6iOBh0MYmIo6KDGJjHOfMd3XehuiOxb4eA1SyhQyCwcUmbJ1Xsciz4+
x/7l3qKrNdiZQQonwvr6CxOLQscCSbdcuQuyve09syXxldRU4l93qgZrggTS3I9/bNYyXHxgGNKg
1PvNwG/eMujRQzgadkW/AoocvYo8oGDNPo2nfLpkTtwXCTJU5O8UgMG02TGzubhzVDszqvDhFBYh
OzxLlB5Lps6eRd8EQLmrvodsO5kveF2vUL3FULWnwXC3I0Pio7ZAxxHa+jD7rPXrIqGSVwB1ITSC
74NimrFUF1SrA/g4MnhhZ8Jx73UlHwMFmSXq8xwu5nS70iJxNhEijSd+a3oIzWoz29e+putc4BuU
0SiotamAmKsl+N+FW4wiiXLqdqeCSJg9EUsh6IZImprlXANbpBtPYgQSVqlRC0HlQIpkCSXa+WoV
jGuhzB2WXS1L54FlJ3/uRhHaePqKmyU/5ucgJ+wI5mqC1iTtLmhpOlsXezebOlvdWGHbSB6z3p8R
TXUrsFAWIY85osGHM/8Mnqf+2NwWK87aGKt1PDrfvVWatuHanu1eUMhN1ixPGmn/N6bQ5JBE7gYw
sTTqSVnqfsIazrQjPp+bA2cVR72x5YcXVDDN9Z2dzSzH4iL6VtNcB5jHiDT6AzeVWoL6GxCaqOc6
9B2Ucyi2nHVJO53oH9GJyZ5kfrRJamm2qNjIe6C3DQX5yX98qKrHo9OmPjU3zngXe/OI8v857dAj
WYxLJMvVDlvq/np5Vl90jusfJ7J+7Kb6WYZ7tzSYUOKzZWy5VrSVnuSV3Zdk+t34uCAMQ60icMCw
/PzlWgwx0ciUhwG9jimdRsilciM8DnbKeqFLv6iGbiQ2VRloobP6alVmrn8Df07FTLw3BlzUQT8c
HyxE+6orEvNQKjj1+XeHqzMaC8KZkHBlqP1Ks6cMtGx327SVdnAIGgl45LzvSJ0FFSG0NDKmGvsG
3i1XcqHKzoayYB9lcoy6hiTv7vDP6hKTgnr+3NfbJlhbTfh04lPljuLL9HaMevP6Hq6nL/xKpL//
8po5k2ELX7kDq6TlwICFdgh2QLBHxz/5qMPfS9LNFKgFfUOQ72A7YSs/sEjTQnDbqsX3jzx2Ub/N
UktII6AxnaRK2rD2YCtmcgQphZ7mUI9WkDm5nEb2aPLrNWziPojD78mMpvzFynX0PauQ8X76YwvW
oj1gvHbaYAteDZ4NG9tq1wFu9IeNLLX5cxl7ZdFklmQ82ybHxHfqaxiLZ1+QbB5OapfG2iFX7NvM
NN36mbtk5fbUNa4dO7NMTbf6p0G2/NaIUOXA8+nqBRVNVYNZtYlwxLJ6Q1XNfcaZhpGF4J4pgKXo
ZXrjPzd+Q8lL5Tme6XwTWpNGCLfCTrTPOXWmKoqZN151UJdx9V/AuCSG0pK54NgRPk5L23tAUwRW
jXSVcUnQt+gG0gLFmm8FG+CHbYFS5Y5IHu901ZbCQyG9O40WbS/49Y1HeK/TYmqPJ5/HVCOVh0qA
Trv5erj6fwAEAwQICFNakRKmB10XySZrFBf732ri2SmfPt1DgxM+jFXDWdzPuAPLNr/woKOM4ue7
dlpV3Zib2vWsNVZo+UiUo3L7CJ5liMQymYabWGBbE7NWHtBvY9l1zGL9fYWfy2UoJwBE4HW1hjI6
OaYJrlKqLbq+srfH5D1NPPgFNAzVLEo9it3dqZb57lbRO0sT83q/+woOFwpMC2z+Bg2d+kOqai0y
duSm1IGAFqx+6whInFYCxYIH/9L7uaKiBS/VX2j/wg3xC240kDbCyr7eelJYVfhXZ8dkKNQwai+z
OfMyXBXJKkDxKRJLwE4vj7n3OUPsi45ICpaKoyxa+I4NYnUxJlK43Og+5HqGmzVXKUnTdcJlNfv4
64GHrO/+xhZgB2zgAA6Ov3IOG1Y2VdlQmjFtyuPH1yRl46zG2mu1y8b/idl5loCZcw0aFjmKULhI
GHBesV2GYiav6VXCNRQHPH936dczyuds4yrRXHFLaUhUBDZNoehiHERhbO3gGJ97pGaIQFcA/43y
f3qyz0UKxE11/97w8oLH+FP5aQaNFdR3nPcIrV8WjS5aOE0gXB2GWhxnJwlzvUfg5d944Ohfy+uF
Cp7fL+OPq9fDDLhdKfEHXJe2ND8I9EJuM0XP8QclYndy5VUZtsnUZczmAnUTCujWGeXi+rjbDMX6
oX9JGDVnlVS8HzVett7nni7dQaO4ntfnvFGasrLoOjf/cqBBJ9Ae1d/gck8KB6gbFETVlUrTkEIy
b1h039SHWIwuFqXoVL4/PxDQ+E0c3MWUvsjIB7wN0Y5tseOa2pADaR40RsUiDmUY22SBujZbQBT+
pAREbskVVceXeVYbXPD0hg4tUn6m2qEvE2jxlew/KFvJEPHXvRnFV6vNXdEst9yuIOoig+Hv40pL
cfpzFN8bt4wtrEqBeeswpIW4GuE5n4LFZWTVo1oZCjrLOIX56Brh4gkn2uk3SG7TN5esPnHWB8lx
xHfdLB5LgnPJXjY7Z5pRu3WSbUCGc8w7DlB048njO/uaASnpKCdA0vFmE5dmJzagP0RBmV5hziHo
wkTo9UZC9vR0uT+/OhkT+9tvXKj60BlvK51e/UWk4IVDT8dahfEUv8X6JlukzNy/SZqFg/yHPmDk
eJd1soEGkClmNOJC2nHGL8HEm70TJntgGLhY9fP07TTuSCv2LBPZXl3jzkLKDzjqaZvx8On2lJRb
xdVoOKBCf2SBcbQ4kyUBbqs9J5BxXcguAc5xd8IO52lUfTXasJe6Tj9msPdKRj6ZJK2L58lIo7RS
WEZ3KfF8WatTYa9zxGTst1absjLf6G7ajUoaVBbjEbpY+DlJ7gpTnEHLvubw/kdWAY5kS67rLiKe
9Ij2K/0o9CLHWCnAbrjYECdtli1RShVPaBFRFzQPQkqrJf2H3Ce0RI0Hs9X93on94t1rjLxDnDuJ
GzyeAQfxzV1+1xo7JvhZMjFJ5cA8mDkHnhyKZCF7PHIiVukHMpvGvd1xl/rzw7DSxQm5VfQhN3/h
YxY0tb7N2GSPi+NETICl0AqhpH2T3Lv8grF3ZAy4heHU25NMHBVJ8UZyYaFjQSd8d6D6GCJv23b0
6c2Xtb2UTHQpZPL9KIfVINdGRHUyFIOc829REa9KzbLCBZe5AUoNgrURBWCBu8weK4JxT/VNOuxw
Fen24/5+LvMCzmk4JfCN9SXFzEeLkoshEmPRGLnr75t3HgyiOJva4H8E8jcNDaa16ywKKuCtgvUu
mIxWaQRKujiuL/iFtWsi2zxxz5CKDahsgXT06WR/auf69U73g44kF+uabTdgNQYALr6tRxxW+G8B
hICjkVF4eahHagIeOolZFFzaCOibK4hX0a7F9vcTakUCQYr7KsAvuDtxQPbOk/3UsOTHHQgxjTns
EmDji+MGvuODpAg9T7Solpzo9JyNSJQ556kYHsILeV4XkohV8qlPXFuEpf5zHL2g3GNzG6+T5VEc
yMkrJnYUK+qv9TzGXnwN34szxvtiok9ljWjUlV/9YuqXvAXv44iqfkOBJy9s/w9/k6CCihJIXKSW
B40NQdVYN31PBa1jOr2k5RxcYZLOMVCp4fsNcoqbVu1YCWGpTBawKLFYtTEfAhP21EJkcK/FnyMq
F+92FaAIEl/xANTpwQijlp6ohGXmA6mfrEKS7xecHHyLWjyk58cwZn0ojlSt3sXJimj4Y4g+Ogfj
shTf9UT+kJzPFAFG6YtAez5oG+L6/pYzu+NSjw7iVVaHjyeKK1B3WHp6rY7XNIu0D0QsuLZvjgVL
lx1ulso1e5BzdmVKQwUHDx+uUwrYaRfNC7d2yowWlj/80OPkFWyjErcO8KRBCqAZpOdrUuMFMy5R
s0LUUHVMSIhtMCdMmnjsDFZfjcPSC3AXtxxlhPWR8PbIv1G5a3X7BBa1c97sNxZ7hEVQ7fBE4Ybd
gnSpSKubRF62ByS6R4Xgupd8cgAsz5Evap/8mKjMRwY3EMY601rNo8WJF2AY3CFzTnB554ZXsWY1
QiYijipIDyrAmDqVXnQ5PQ7fIw+V131x7rCw+10cDnfKo8bZmOPENp1XtALjUMWHhuMYv+ALQFi6
OtwXgfnmIXuh2Tjusl4skmLEI5l1zNU1FnQnnI/+C8rKSRH5uVimIDSF964BpIzG1PojDEXnWrHS
fTGOTWft6dxNArcwYAUSzTZfT640l+jlABNsRSib3/nCOscb9c9yvoY5MWM1x4MG2YLflpqkIq/P
33f1C4IbeMCBiTbMKOxAC7EIyGdROY+D+enRWFu6R+89y4ICjKdGLSCQzGhHd20/VLGjYKLCG8/l
MRz3XpmK78DqBy5MBgA/Z/DpT/zA1CT1qZcytucVClqM59q4p1W1I+5JJGLNQw2YV7Il+YNxOhlX
HqmtyQFzP07lMMQPdWUvE9ZDTP4XToHtm2Gy4Z4ojlGg6YH4O1Y8a8lkaPTNBFjj7sNRbGX0sYLq
bjcKJNL2nZLn4Wxi6lPVWODOFbefK/l4Lv+mS8Ax/f31AElQmcfQfGW9YKSLjexLY0cxg5q5occe
+Mv/gXmr/kkH4+oDg/woMEh8OET8V48kyV/twLadNam3/pLNLbq9DuA/Zj4v2UvbJPtxgiiU/G6Y
NLLvCeMjMM1F0M9OBOH0rLFugMkMdH+cMQ4dAYhu9E40mlGUquo22mJL/dt3bLLytJmoUYgRXZFr
pxltwxCytlg9+FxjUi/FbNl0ZSubdtXRheWflOZrgeNZe/7td549zZLZurWzgbOmom9Yfbh55Mgl
sET5z5RNQbelwLVGTpW9vUyIxq9qRqBVpnhCdH4ge5PvOQWGZsHz/mu3WdN5MwV9JIjK1mkqtG9N
59Mc0mE0LlURj5Yv7v8LF8jVZBQJa4bZq9KTkm9MMkv7fx+4edwwY3MOWWy3GrbY15lgNyv1dgKJ
DY4XJTDxaOtweoy0wh4lPrK/YxsVdnXh2GYt+yh7J7Qh8V74b1a7vtEwy9IP3RNDMvOArVxYHkyz
nKsrk/G5r8O93yFeZpaAwauVh2la3FFiGqUQitnA1kE2VPWSBsZhqYlQQVjpBbv0IYHbO6TDpcbL
8WzJtMzD7u21hUZVGfNWPAgIeK8q0jlumsfh0aYpBhFlKKP2O2k5JHyrL5DD61A084QrjgArRSeM
1yFGsO3YEQ2xENPSCpZMCMwOlFHoHENEcs4kuyX7dPjlRQ4D8xnArb1N6G/4OgkwtRAZf1sXU7SR
gIM7KWkZBcBcmAD+4Og9i2lWp2C3SJXcea2AN4NKn6QDhcMVxcrNBdQGu08gnEAuLbM5gzgCY2vC
Hb9en7niZQDeL8fPqwcZOyPr8TfzLOpO2J0Wz3vJ6PoINb55XjDzuyWS6A6oOeXozQS1c46R9BOe
+TWIfyMX5vPmp1dst/2OmMJDqgKCn/aD9C/Km4PqpUs+wDHXXz0ho7tIny2xbNpM9wadE1/OcRgR
LIHtxSJwhfw/LG1uVtWWWP4L00xvUpBQtabp2e4IntQdyZBVaV5ai7iBRG6RUvb1R4r/PdRIfptV
dpdjgFkDXUq/IGdZFfzze0I8WvaAkuz1t3RFw2Czy4Z8tXAkT+t15yboJPS8PpBluTYtg2olT6iT
+99yxnf1GI2u3ftRo9d8GVKQAd+Xy30U/Eh0he+FJacrl0dP5jjtECKQrrBA+YI1kW3i//IDaqce
jAcDfBu4coyaEegifmTSO9j/rVJkrTaysQB5Nsz/xzmnYxE9/znIekI9b0DTGog4wj8yLK15JLIv
g0EhGTy67/+aPV94MVp1qP7WZOi7p97F2cr1kOx0oXKFOf9EItZVpNVlkyS+s3kL6C+cT/sprgmW
z3axwgzFjQ7R0OvThabn9EDwtXfpUmUzqpNiKXguQJJwmyA09I2gtjAljbu7wOv8SPH7kwiP0Y34
Qfq2K1dhJgO6K+ckI3uPnkduIZ8P2PfD7v5kXXbDoV9C+YjwRc9GsZG8IHyFC2F4pmiupXF8+xqe
2JhW6PbsIHpbtmE7iCIS4a0KTF85mEkMzrjfVPmGoBKNOxdo6JgZpETL90IRLG9oupy0wFy8yNzi
9nq8yfw21HzxKc8gfQ8MK1Xy0WCoEO/pNvLV7PPtRHJ1iDhuEFezIxLCmGpm6PmYt3deeZvl55Oy
xSf1yQgDvx9i5aIjw7oo7N0mXII8RCVo4JGISLi3VWQ1t+Bq8CnWUBDooFc0yag8dxA5FdGl+mgR
EZkD7+xzYfNpR05gOBD4d5Zl/R+7QLDGvj+fdpt28iQgDq4rPYLMpexxP6NLM0GUdYvE/m75y7Q8
YRL3m4EsAb8gVFFf4jS5NYih0QBsbGcz4l48ASwZynB7D/dmKps+2OHv5hS7Tqq+tB0uEuj1WSCF
oKrZBcsovdSU2ne+LkQeVSOjIfszJxpdV/NvDm5bkmEldRBIYvtxrpse7J78Pwym6xpxEWUcObkF
SzY9ZUFKIfDRxBLS0it0UPy1+0QrQH57Wl8fVBcopFprNoVUqSP7SW8CUhBU/Vk627LuDgUM6Ncb
HMIPRSHx44R9U4MJOuX3jFlu0WwSIk3Fq+eFauYsrwclXfXPoFJOO23YCyKssACYCv213kfasSMB
rwR5Xdzj6C9wyDUx11iV+BLmtXi2q93+cZ9mFxdy+Ajx9TZC9LeAS1wA4iY5dfOhzJDh167Yzfr/
jab6+P06H0QrNDCtM9WNZHh87ZU4iRZKIzV13DbR/W5ZkHCaprsYhXoizYCt7MWJw6fgAb9NFE4b
o/2KAj9hQcXRlL6ceYxN6tyMOlGThOeg7O4wqKEvb6rvFo02Q1w6+eI7yxUHcSi1ieY4FanIaZzF
JQjW1ayWI/dHVCnr1Ki+T8Og+KmsJQPeS9I23FTqmYc+Z887JuckYke8EtmzcvIIj5IYiB1oqP1l
MWvtpKB4C9TUAc6wZww3el+5dTnYEc0OPeN7yjwnDrtTmrNAQ9eCSsOUwhcVntEj3TzDX51HRqMU
OKd6JYtuWwfGgrm/LKIfcCXf3KGNrKqyMO0RIXcrVrqna6Kh8nZaCMsrkYvhEZzld2e49XdcNs/w
8GpiT+9nyIk56UUsiDlhThaCoUK3oc9HrMxaIXz3A3Im98kP4bsx+VFRKw29mEFW0MLe9CZIYBfH
LrjTCyANeSEWJKsuaj2Oi97cYL6N8znYFsOmvJQZVdxvkvf5JIyJP7F9OTRvwa2rXoRTViMBMR20
9IXIygcyeyiQn4spn/zu9nmjQ602WE/Dys5ZdKDQGfAf6NUr4FzkO8xDFDIRDJke1U5mUPmoGS7I
MfLiC002gF5CT67xCKO4CrOhp0/69D77tVNgu3lFnLNGCW9O0w0m1zmDBZAXk/ynCwtrJYUwZpxB
la5xR6D7SXuhKazwk98I3GPDZdaZOloW4f84UTiDZ27kt7ZaUcym73w/BCe4MzL1Rjev3MLYZjzy
yCHwgMsBIvyr1hpf7U5NCRbzfCPhiyFmkyjY89IovQabjHAuu4YOnrIlgXzuzIsDJNxpEbC7/EqJ
soq+TZGvcZ9vbnw1Wnx7ZZai1Q3LheLS5pnBx0sTLfZeLqRTMFvv3GMFRRy6xlu28p3BRfUQ32pO
MLrsT5tKbbKPUb/I2r3h79/mefh1Xh2hCCCPhwxQiIOKa98iwml+ecVsN6uSCiKDy4Kv+IgXOQyb
gGbLWRZIz5DAn5ZEzNPOFMsLaGfC7C3GsGjHRpxNwlw/L0aGOC4yjJuExH7HmDk13dcZkdKVe/VW
AyXOhiZmiR4pqoQxqQL6V/5iRI0XrC8I1qYgVeOmsh5XIqTV/ex0Ng8ZgGPpSFhjr/TCyQoWAExe
X1MnG5AGKR2wS7wxb1S7qtPfqvY6Sk+JiGRRg3hQyLEZbdlcynxdVrUIgFftwjeIsl2eSNmc9bGq
fJJ2jL3Op4rgrl8b+LdD2agT0CkzJFgyaqrf94FS5k9tRiu8R1nxDFX4hFpogUgDHvO/5qSeJq9p
UoOFk9eTVmup3KSReMTjyfkBgXn0DGJFJUxgDOa1wYzjvXrBthw+yLwIEsrRsJXo+9YHUpFT7OUv
jmwgDG9W8qOGkL7H2CJ6JTkdPbGLrCFDTY/iASYiHekZrQ5tdRr2zCuk6DjMubEauURbbZmS27tk
M0z3UyuI22vVQ0czCv38OqPktbfggCQYtE1+YKW+bg4V3LzB+HhCRsZtrneMRU6wa8you0CEH2QC
I14I8oL3NUWCCqMFaLTVdfS2FbcxncsgmzX+E6FvnVoZzzbxg4dw0fvpEy9G0co5YD3CDGA6u7mq
qdNPRBqfnjDAd0csLyEBlPzjEcGJ+zK+HfpBVITwNF/8QraM0K763pH5s/VlHiX7exPM+c0rrqCt
yJiJ4ie5H5qIUomWG4G0j9pkws7Fm9AbEgnwSydFVpoz+QfpuiDzVLZJl6wAC8Kciw/YRMTlAu3h
IDxw41GerzIwci+0xWxHed8oDWiUrq0pFwNG9qIyEkeHFM6oLtfRX7sx79UgFAbaUky5Uxk36QfG
Bln+vuu5zwuPcP07HfK8jCBQHZjKcB8hY0d0/1DUP7dd++Ma7Ndg9S1L2BrKr9SmfH5tbq6uHN00
lu6w1MzFDGCaPRS+HmpnfeMQ0l6Q0ATbyoNGHyKyrdAW4HA6VlB+HvnoBVHHNP77+62VZvULC8Ti
QX37sDwQ6BOh+r9ZoFsgJIcGuaAUAGvEaUd5k9P2mDYBkHXgX6dvhyHEFauansfOBw7RWExFtsiY
rNNy3baXBVxbiJP2CSVJcU8n62Sb3L7lNlbhgSZjbbX1ZK16j+/peItgeCAb1fM4HEzAC5qqo2/6
iJNqTgsvdJeiudEUs70xm1j3Gs7uV3WBcgEGtlqyFMIuqOS2ycWaGJcp8lJOMxEF3EyBWTGINRbB
LOboukEWqH7fhGKeOB7iewYAZ5l5SfInpg2I4WUYZQWm5oB5S+bXpa4xP/fIrIx+uiiuLmJj1Z1i
BZViW218C/6l4t9vYI0CmER48Oq9r4+qMHMmRijr1wICZ4zII6RnSvdli0poydjL8aBruqv8wYaG
AdqjG47YdAtYjJRXieH69UjwC2fmaLYXo5afFK9KV0X6M0sfthlvgv5PdaoziDE4PrudW9RwkPQj
jX+BRMQ9xjwWic5RlmfsKDmOm4A2GZs8QvY5bCfX+p+pgXtfrl2wnvJoV3RPwpuVbUDvo8iDYo4A
YJN0jD+AwGSwliovk6wQBnOqdlX5tkpfXyvyqe8r0E82pYFUqynpq/5YQaaoxnrvwESsZ3zzpLCp
ZbYOyiMNdcHLFLN0gD1uTZKRb/7vfe2PRO2WOoojm4NdI4TIQ5b0tZ+67DjKB64Uapt1LjIyodc0
HINmJ15RQ+EtCdeVniRGFGKBf7Aw6UDG/jViRbq5JyWPHahvC4dVZ6JhqWblbKib2KRN7PB6k4Ob
moguBKQZoTWJIE1qvzH6kbRX2we97dD5PtgbEgsp6lWa/uPdPulniTsEjxc7YYJlzkh90x1uQ6lf
AZncv0Gfz0Prvbg0WADSJnG1aJlMkCVo9/XMknk8isFE2OW2hl03qmLFHAFMpyo9Wc4hVa/jk3ej
MWwiD+qL4Lm/cb6zUmoYzyvF30MSWoET9q4otXS9jKFDFPRXrqIXjq7liKTLr+elMtQQFCWqrEoW
90KU1/LljwG2zsjG3btyArIxh1kGPrL5iptIjSbiNZy4ZOGv43A74tvL2yB1wK819o/QHlm9sZdt
Fci9aDMZ4QiNUE+bUqcfC5RkmN4ctZFfhnBFWvSgXtW+EnWwN4XnezNFnttiewMcPZTJQAoBtwER
nF8B8BiuqRmQANPVoM17AvLsyZzv/Ye0wVVs1i5NjEFVhKGohr42HOC5J0jm/a36IRQ4OGZyg/lA
Elc1/9fyGhJEaMGBB+GybVS4DNHov9H6up+rrEJq04DnNL8vc3jpKxKL5qM9IrdZv5NGRtPL8ss6
L8z5J2FjkZK084prcAZklCwM+dHaO8SsOUfK7m4cAyz48QPw5g1QvhkOQnYMT++rN8oYN1z++lTN
IyvPD/4UqDfCD4BfVzjckEPmd550FOlrBgf5chMTaUjSgBG4FqPKrvWMRHLr3rw6hlYTkWvs+Mc3
Z6yp3ey72Yi2fRj0+Ypcx+BxYvgNihXQ+xg/KIiQ1X4SorC0SDrNUYZo6GPU8iR030SWcT8sPdMa
PJRsUZX798+GnyxNyrcgYH5IaPyr5dUmTAxx9dPssBAjpk1A6MRWSXY6RXfMsDZsm7Oy7FpIIsiR
s7H7LFX9hXaqKHqjftI0fuHTZR1BSHhGJxz0sBWtLN2lfeb4X6r+RfgQQTc/VJ+YX3RtwR1rlK8T
ilxYAMuXDnBo+anTQ/LNU4pqLrPdtw1ztbAUoDSu0FVjmEd7B8tljaqTK0bKjSOgtZ+BguCX58tL
f+0Wjnpg0NwTH7yF7f4uyJv2DzRWiLno9DCtwl83UKXVR//8OBruLii13zCNOP3g24Cy+6+kXHnE
MbMkgQKUYjYNTZs9nvwDz5wk/EoiKsQ/Rz3VpJiCkil0/AC/O4qslrAxRiTwNq1FHiLMsUu9igvk
zfQO6jUZordAP9rvHezttNCffnn9av0JG6RUtimB24AVaS84BQaUdCBv/4zyNZTUd1LciRLDbtWF
QzE3RcAaBfscQf5cfSq1vBJJqbma12bM/0rwYlEPBbn0XuNyUPOEI+kTvYqgYtZDXjH9zkb4X0hK
14EDBIYv5dhX2a5mqaiL84u4PIbx3xXgJoNf1dQT5RlP9BKpRbD8Vbh/6Z5fsUEP1DB5+VobiyXN
+uaAOSvK7/yNLucHmOOrU6dppgAwwtoHPTOiRB9Ji81KH/i8cTr6EVZ8USp6RygjJXCp/OjeP0SW
SFLePB/J9LzICNHREorOgoiiWkjxq8cJzfQzp+0NdaM8uWF3+1S8vp5O6i7bVBefJ8oksm62hVPn
F3zzuhpzCzMqmM4VP/dCGEofYX5/hlGbD5IxH3zYtBM4YD0iq/ZbRSSeHqY0Az+zL/b8MtRxaAra
jDqO8f7t/+ywrXDENzigBAJIx4Ti2kNZOsK1YlXthKjXeZrf9MSG6ihTLYD1LvUlgon23uxo57Wu
2GsAxAjZd+YK+vRxZAKtVfgXu0NidQpy3kU7H6xGTqB5v/F66gvsQyfl4Xge36vf0uBan8tMl1wX
MAqQKGKU0tS9+0pQtK0/tPoZ2H4qEV49El0dpy8+d01S1Kzc9oCB7LkWOi6N65q2/O5xpTmTXbRc
5oMvu00FbZPSFEHKG6VGlkurfZVIJ/0PafinIXMFhapjKrOwsDtzibAfwMrGZReZrCsM0rIUhFzy
NLkBLO/vXvhJqyGjwQkj5+nx8jUmV7CUKkekBkZP7k0DDC27KnjeL2BBOyRp2a6eRay+eKlKXm9V
XRvgCv1OGITpYfCCd2saw/hAOyqvtFKD4wwBgq9WD369O35f8XsFBzRrFjE31P6z89TCW1L6Y5u9
Vzu4ulBS9a+lrrYxvAbtaKRUtLTBxsrYKHSdIdhX4Atguil63Sfm8m3vdtpznzc/o1aut2arXIWD
zPVGCILab85aJTwJkiQM1JXpIFnld02anjF/iCg6Ff5mL0ojd9rhNkICc6zqq+b8/GUhdddjew3L
9GSNwALlNPWjxPHZu/0WS+SyWZcxA3y9e/vePexVWI/yzcqdFa59TwZSuaZq2ofm+D2yKZuV+Lge
ABgD4uSIDthDxY6t6VDcMs1UNesR8tNYbXN44RNFawPCs6jgs9PE9RdOEVva+6j+kRlfNjdZe0+j
hiZa6q1nQE8TohmGKM26n5hno8fruugDPDfsc6V73QxB4F2HNlLMG55XaKQ0dHPoo4aNnHVsJ/ZA
8z4/0zCGOPEaRwT8f/cY4UtXfCcqia1kYJeHF80/FbNYfju/lQsdvghW1iImoRV1uYh6UCh5FFYv
3E6g6LxOiWPUgqgaMCMrXOjzeYgqCXcAtzEKZPDb7xyz1BxVkUxjrco5br+Kdr3nwAeKZJPLEuql
ByWglaTDFHetegNAuI1AakJ6mGSRbVlNK0t4oVy5DW/ptBPB5I5r5tTQdYFhZMHT0VfJ5uJdY/Hn
R/8UNLMHDjWSlWYVrOEKe9OK/YWo5j2ECFXxib7wI9ac+OiDnv1k9CELcXMRKOtKsyeZvTW2E7MM
wbHD3WvNcBO4Evc3ADQW7MSf4CVp2rBHOqJXHK+H4rcEkL690RvpiRrLbb3/rtZKsro7M1ifN/Ug
lN+BksYqevQ0Zo14cIebb9yiWkUFdeaLwzkEVH6cdZRIBqzIxEPKH7LnVI/i1QCcp8ABxAhyVvGG
rRuqOcLavwrP3HEQpA7pxg8W9PMKBKeLFBcML26i4s/j1/GMA+aMHxTaLFiJDeqK84l2jZgzsTM6
Min/qGu4oHutCVudawiGD+x1zAJhtnfFC0u6+kjwGTC6YAIZFpuIimyzMda/eWhMF9XsDtM4ASfZ
9KmQuewCZ0e/a3B5g92j7FnnG0ezWCQoTvjZTNMbghUguZ1vpwsMCku/JdqtycaLZH1w0O0v2Fnc
/SSSvfFB59Xavo5aOimsADE4inC/ii3+z1Eum+uea+SMTC9f1X/bVri6Ummz77ZgC+OCYpoeqqXU
5rC98Dicl5fwatZEqmqLj5ZMZBswkhNg0/pYOw7sn1qQngfR+QPgQm0DhPvPxhgHvi1AtVSX3Y1t
N5OLaLcBMOCXfA+03lZSlnTpNAzdtbNtoe1wYXQ89B69AnUOyGF8lf9waRBQFOLnD2FZzPKHjMRI
v9YknZGq2a3lxWBpWk2C2ckhArvh3V0lAyK4IE1C1gGB1zF/4Jnm5FynSbQDcqIS/cpPHCVALN0B
7P32rE4cgn2ImO42n30GTLxc8hnkNnVhtVVY66ZU3tOzaCov1oYa6kDrT/AbZSqXCdKBdS26rl9Y
i4Varu8S9In4BlA117n2apB6jW616HuwgHSWJEzMj4EA4OS1/SuAlWwR1gnsmSHnJCIZ12wPe83i
ITosB/4cLAkmhl2b+ew4S7/jnFAgbmUaBFTVnNPt0yWI/P3BN0ja+wnWhan/4s5lHYC8oopifLwt
LNeNgZKtByLAcSYdMSXAn9aEWk8szQ4e5HHV+Gatek3/eEIoxu3CG/5+XYeXi88tSUqqdZyhHKN4
DqvFEBXkwpMh2ppPFmDliP/7mU+DkXvdKdyMwyvBSarwlUiXBJfMTprk6ZbY11t28B9QvTI5aTvx
uJ9q7wYivd4EsAc4mVAb2OTlWFLlr/8xzA+kXs0CpQOI516XayQMxiqC79emNYmiOcZGDTCmRJhb
JvpDG1TbUCMgZz5HrFhw4zkKqIBT3QpgW0d7SVAjamcejRUUkT5eWnRZoTra0yHuxO3PaEcF/PM8
9LC2kNaAjzupd7iXIbfLsPDOOpXNdTaploGvHfRGEy+4IFIa4vI4HCnvT58EjkV99DazlxdnpiUo
BAihc++dZqsTTlWKWKPBNrwI/mW+HZewW5LtLGne2L6sxE6DgFvph53QjG2fsMy7V1OPWPuw87m5
BPhy+fAEopEOeS6NBrFwM0hHca2MI7NP21MZHBxfltj0N3N9cZcoOvV9i86vpXUQoK16oSSKJB84
axF6nG27f9n+IDVmvoESEtVySZydnIVYtIihHlknuLpNFmgOTR3RRupfSt36AKS3EgW/+KrB53yU
nkDcVt7Rb4FrRkV5jJkHSlozEEUX8NNP/TDy57rCoWxRenAixk5DSw7F+gyPFSxj8zfe0UjcU/5M
zi5HJwTv+6u1VDC9KSVL0U3Ed90yyCN3TThi5no2ez1zutLs1tiQlZ3QD7zWKZ6DXfZD9/pXceUj
T/1UKux1JK4JIn1W5Go+7khnc1zKIW2ua8pddoDhwTZkztOm4A8SSa69lSQE28RCneyFuBAhqCd9
2ViO7GbstnQMWwoEX4n0Xrd2jPuFr29f+edSHazenc+DyYlxdkiqVdpNhWDYDmvuGmI4A2j24KCO
tiUMoRcx9N5EMvsjW2NbSD7MXYLnR4YjXuGzRo0Yct4alTVUOyXVmNf4PFnJfQSvIn8ODr8R2W5j
xTI/P6T97PUeh0ka4W7EnaWf+4RfGEW+LsmtyJXa/I797h+6ApLi7GwD+lkjuS4WSVBGC59hFPch
Ae1B3H382p4queZeh9qWO80rwCpAi/5jPwDTe79spDI9WaeH2j7Lk4R9UzPRCogv4AKp0CT5Zxl9
ewwTXGOcZkHSYXR7MDH9VCfQFlZpe2keoyxx4JH4YTzkehbmBQbhHcKlEi9yYsxR9RQgziq2BC1x
waKL0TyjucPirBieFKyfw7oa9D6tnDaWb1cJ3/NO2JFF5ve7pzNedN4I6RR/U0OmhlWvpMtvDZ5u
kwRI9S9FHzkw66siXhz1wrTCh+aaucqkUAk+aULd9cSKV0Rlk469f3nwJENLlxnyI7eHDRU/dZeS
bYPRoGTep6E//lnVE7WkvWgyHLzntW6WyLlsTZx/bb6uZAP1LeGiMGtN3z45H8y1L+XEtTTKsMkK
uC/z58MtsJET5nURyPbKWn5oha+twL+R5KRwnRmg1cvFQOjjog8Hj3Ox445VnYtbnz6D2ZdhUqGr
t+6Z/6qHrnoeN03vHwGzh6Lzy/pvwZAsc1+2oYsimCFEI07gOBvzmq5g/zDVG1pEAEbSrjZWS7UM
ke2LMmvSqDEKt0VPs27rm2yYUDgBDAmYYLSd6m/AUCo2vPgQf5CNXLry8bb3OnCBgr0sJY61j2z7
smHpU0bHVlfy0JCB9kzUsTnGTXw/vOJJaYHqcDKTjc+ygy6QVCTri3X6d2896/jH5WcKAeomJdXX
7ZhOyVrxd5eBaNSgaYYTQAbQ1kdoi3Ciwgqo0LkAFiC++BcSurhnYNpAjJHZAaO4MZrjoylZbQZm
17RCGxXMEHvy743EJ6Q3rCHkhaW9PRiNCt2Vy9My5xJcQQwKNTDuNYR4I8w3DR+OHybK1yGzlGOM
9VyAwIA+vhggoOBNwOmrrdh1c0hXqvDgqLIK/Bxl9ijeheB4TJO4BxESjcfsvhxJgsB64OHDutzP
GwpdviyLCkgBgFs8FAuAUy5vnhD7gW/RISkmodPAeDiBUz9jdMBSEbHXKF9sumCM7CjCWDdl50KZ
15UOAyPjg/nV4fgQYknvCyOhjQWYvo+hMq/umTpGdXIQ6pK+c1vmBlXMIFLQ1QRZB9D1geMw6IPV
5XEYiSlkyycclEn+TLQwC6RWcpgg8BlElnsYXGEvXU9xbgDbIz70r2P7C6SG3N8qH/hoShWkPjoZ
+xtAabz0oG08UZSdSziBy4Qbjqr1UaZRsqtSSelPjzGK3HECiBS3oWtIxzvVd77yOzQkXTDlEr8c
egYwKsstv0avz8EhyW2QNOrFFSXOjU6MISLUha9DyoRXzqpXfbMUTKyNwXjt7Iu0SVxtatS9sAWY
AlFVyD/Zpu4mDME2qxmIEEj1OcQJUlKUwC9zTNLejjjDLqNoaTC8glDbQH0K0ZbaF2sc3N3PpOlR
9d/ozTT6vXw0wgDmhj6b99alaDrf+G0m0At6euSv3spdcUyy42A/wXEcF5toc7SUIcllseZTDSb/
Zu3R7zNJ0Z1xL3F24lO7CqIknIb46H2+T43OMcAQOoS/H5gITyw40cZg4dOgxEo2AvVFH2r8Fx7W
XqdK3KQF8V3IWHMKNtAjn9iZIb2MUNWs+CjUvsD9d6VIdFPeIixmXaFhJJ0KraXr2LGrdNsTyGGn
HvbpA6ZMcEN5jehuP7yZuYYMfThti7hVLy3YN5DX+Gy6IWupHk97cgBTlsYiHM50gAa/hwei0xam
kRaocVOL+thwwcD6iMl2P/h0h6B6XIIgSGMkBvOTqe1KuNKphYrmhE1+/rzz2sHEorysmihHfSjj
njZPI+YrN4WsoQllPkX1UzlpMB1tgLbnGQpnFjXTf/uxiLBOhEAqdZIUVC0M6qjQLcJJzRdjqbs2
1OnE/GxFo7mm3mRqGcnyU7z1o8T8oRGPyd0LiLNUGmuHjtp78SWWwQwRZORqyDbh8/KM7d1AISn3
Cerl84XukJoPTDPlp8cXQP9qO3suSSqO+/Nt/lT4008GFoRTHWNLCMbsVDoMhiWLxYRjixaRq+SS
6f+BzUAnWxs9KjSr/Pnw48chdZbJVr6xcQ5CZZJET8C5swv/QaAJAnhyz9YigKVmXufg+oTAerhC
BO72xmlfg/gVw86EAlIkeDGnct7vMbkgXHoM0NR8tDe/Gd5/3sEbYaoZN3xogmii3KB+XmVMTb9l
k1FSgTsfd4md7ZgSc4fXPaNDm4jfS7/1xi7dRubTynAfCQ/QHTLevAe646Th+XZC08Agm/JShoLy
KTqHYh8QQHwgWzY+/KUmZf5aF20zgiK56n4uWv5k+Rr4if8134JNvK1c46u7vsUCNsBdgOCf0ujp
pbKErrgBblmULUp5V3rwT7l+Xfbm0Qq+T8gb76Kxkebx1ecpCf/n7QtkEDBEAEY6Z1p5DlIjlLHc
kvDx3feu3IoszJ8DebkuY0EkVleD+bnctJNHQpsjja7+4ZbbwJ2/EIiSMds7i2B8kY71jGwgt8E0
abDyMRwP2PPDFXFj8XyEIX7RfMW75sb0ov5+jcJjThi4BY51IFt/u5tmvh0aQ7ZDOUuLKnxmtnM+
D123Z4p7q4XcKkHIdqY6lSDpanY09EXdx+wPWpNtNTx9VycsKVDZD7nfP/DOgEO2syKjHVdCgig8
p8MA+lFmR3meBm/4wzfHFObPDEmoNaRLULlpXOiSSaXLznMg1MII/xlw3pk2a2lCr4xPEZiL1Gop
cvm01H+5xKsw/nUFl+lSOsBSqYpjg9A+BAyk7t/AyUNTrr8cVcy9SCH0E9OUZ3vTc2dQGjzleTPb
1M4B6aWwH8X7qCWQ2JDEDX5eVtKiLBfGw3+A3cPoDYSOV7DSZN+6ZjwPlAm32+dtHSCa//jfU6Fv
AuCj7vEE37zKnFrhi9ZtU7UR2/AuZIQIo0RLT+zCDBbJuvW1yt7+iu26wc62+QWk+gVVpI/7du6R
l93+DSDMh3dQdFdUwbMk7kA80kidfFObHpMYW1WsnLFKdg3a9odtqyqRM1VOnXR1kNVu1PJuGn/H
7ftn7fAcaB0HN6SMEeUlkWHkIILLCkkuQD9IlEyYvNzbECfSPCdzPlFq5+aWSwZ8wnUmbOQ0pOx6
dEeOMOzN9XVCan4RTaLztMjDC4ZNMbh5FUE5Oq/40QYf3PqCdIcMAcwOoUcxpz8w95RA94kPptTx
99yMbNz7a7fHTO7DBc1pZI7EOaNWR9bBMp7Cu2NNrpWpmTwVa79RI+TpAN5XEaBQo6F4U4i5mjZ9
Pl83i3Utq05gXSiggidsccbmBjzFWFlfIxeo15Al8AzsTUY62r1+o4VSi9FlzpHOSIWSg0t4E20C
WuFKx5jBDzLGZzLT3lujc+DQWbMBy1mi2nkDsGlVdXRAKnNNbEXHCsjEzY9vugyVq543rCSNcnIn
SDpWdbusAQJXvTsNSMcjDAKk0VIgHFitfe9lWyjfguqdXsHcRzJfSmqrijA2orXtKr4r+NmyjUw1
pWD4MU6U0p5MfhJDzBw0XDtEybvMtypvCJZ0hUBviXUt236PGDwmFOtd1a1dvFV89jfplcMm0qao
IBLuQXY1U34uxHtzjv7vpWPXyXKv6OoCRePDVtGLPXry+kVbY3nGd27GZowE3jMbxIwdZfEuekdA
QxlVxvLywvPV3y8/eGV+tch15miPx15ChTz2jv1i2McO207+TcOEezhjnZwYHiI94XMlI2FW3zsU
b0/kJ5wKg4ob+c3rL++mrqB6ZB3xsc6KzekfqqVNEPdIqfO4Gp1w9+pXUDrw0qfFEMpoEK7OqS9Y
ugJQgwHvmlg9GtFp0SCBLfIDt2Jw/6JIiF6nykGfDaUk3BSqhRHps2DFrcpt2E6qt9oznGzxhAJv
3deYJwXFY+bi/f0A2b8OWVyjHKk2yD44BiGXiEMrg6JlxeJBTwcAelSfpcVnYOTgS4/PTBcnLJv4
Vps+rwIwxRygopBMMF70RsMTRS+iUfzB3f02Ab8jlrogEVQWI2rqyX6aKmtcbpkP88hFsV0zzZkP
eI7hEV4wvuL+wwLKn4z8knOOa/1VJ9IUe8ocmBxO7R7J+Ga/8mG5+Jl1R+M8Sig4JDBIfJ4YEKwK
AmwctHzRqGf4i0sXDtGLl9UON5gBu/T0V+lFPC7M4mON4TjNp4BYe5e83T9RZKsvkkTBB4MRj54E
hl++Fl/BZSMOSOP8wIswZxK2UODBaz5LoQ9NLm6GCcJ2xIQhOOlPdHnVCUC90sWOqR7ZIGd9X6O6
/ALOXGFINx0HTYA6clP8Dek8OPN036K+fKUBP4X8IxYztCFMp88UaU68Me7x4864Uw4vncBjUwBj
nVlSgZoweLtV49gChSCwYcQiCX352DT+XPAl31Lfi6GkOTCLGA33GowL7fLEB/hGG1VWO+99bbBB
GkZMlmhgxJPU3pAYlWFqIjWtWkfefY9qQ+BlhrxkT3rR2iaehXaQ8qV+JR/Q5HKwTPXLCp32546i
ZnUB+Ed8qkeSupxpKzwQk4nA9UzEvOaji1v1EkTAAUDAn3pQOhIrPpMqWBD/xPq1TigE5cxxqXKY
QNTvKOuX2wMM1kK4BBUug0GZVee0SJRq2sSMLvEjJgnk/QsAR3V/vu8MQMHCzRpw+Wrzss8SgUPq
2EmWA1HQFt8nf/cDGnTY7bvng5JqXNHmSzTX2eT9uMLvFXxe81K78Xa7H6FGezA1DEq4TmFXwscI
vaYRpwiHK/WBTT29rguhHhMCHreqBmQsuAjpDsvB9KTjEC5kqroRI9fiS/Sb4VzqhruPXKo3S2Xq
4YZJUeGr6UP81j6o8Wmsg2Yanw87PfDL238TPlAodO7PdDnWO860NJ3IEX5v+AcLs+u1qjvPWeSD
ciOIUbXlGv8H0Ex3l5pmcCE6qeFrqHXll/UxP0AwbynZt+IqM1Q8eikSGIShcbVF+HHhOhUGcCdB
VJ+hxtp4dO+QKgligr4BiLAzW0Fxnulkw34NCTb3lOdGpUuDL3Hw9sVXEiMiInW6+rQ1OYmXQ1sV
Laj4a6b9nPd1C6co5A+RHW2OGreaVm9OAVqFoWFB9PHakQJcKIsjgFRIQuIfZTneHasMwaCyOSeU
5s9+uXdzwdrjqO5JQE+KKxKBFfUEzIpXsJeuGR4FU+nVeoDYOlTgm70Qndb4IycdlTOr5mtUIZVv
wMMLCSW2l611Xla66FOMCs1YNV1TUhWcDa/P3fxvnHn/kmrRBjQZhJaLctwo2BawecQvKEypYZmj
B1n6bjTgfttHgSx0Q+MGggY8t6m+fi9gwHqgRYH0Aghe/Xm3bTQKo5rBtoESIPFaEVr6fIpeqGaA
a+tsCbsNVr3YyTuFNK5E5DqD5wfJ2x9mWrKbA1ZM9V6gzDFSG0B0BU055VcnSIDcpHI2QyK6G8wf
1mA9lGrU3bodpI0k2tw1UC1TmzDJNH+yyzoWPIDnjvtr7bMoA8vbV5dL1v9Ogexm49FmxwZ3UB3R
v68hvsemtLKFDDptOGhRZeglnOfANOfp2SUB40HoB20iIk+/bGUvQtpQiynsZ8rWo0mgV7Jp4+y+
jsf9aagtjaEgbG02ob75JJ8esXMdiHLlWWDWm55qAcbUm5lQR64q3Spf3E9g6+tY3oUZfNYGOqF9
pAXEsXjySvjctIBMUwsVaK6dLwrcIjg13lXuP5yCtY+gI+mIYDXBzvHTnCubsCB7XNSzMD2c7rjy
NpiW5iwPRJKzlg++OqtHgFLgtd9hUhncuTI4g6lrWrg1wzpSjut/CjNvA90jq6O0FqkRPmIF0zC1
W0cKk5IePm7VEvrZAsuaKo8qPt+Nz+HQwBDo73+TMpHIODAlQevLZ/7LIEZv4EYxyMgzlefvguxl
pjHy2uUb1td4hbw+EB7DkHyyFmeXxKAZO9qAWwjmglUonzwiacjTkps3Qny7eLTSmMtjXQ0as/8w
cmbvIFjdLFP0KYjyWf7LtPlYlsdy+yXwDsVV64GpblgjfIhC6SV7bIOicJZWDTCJ0sNj5QP5/fwI
JVZv9buEE3XqUDlJ4Lv7Y14IqacI8wa+T0+CbIwfjfwW2vYETwTVKAQ04dh1mME98o9j7TC9vTRz
08kiRVDDfjooDed4q7roonlDlb08v7wb5kRrCkhqwxaQXwqht4JowW3eB2UfwvciJ2DvwNVZ7+vM
RIJ++ABmm2pqCVUejt/48T/o3qPQBbPgOOd9cmyvC7cu+oky09aNDGYzmNxhlpFimMZ+jeXousND
hxH4l2ES8n9E6tUM7JjvvcNkVB1ZGHQrHLm4QEXCZRD1js0ylMaZrO6H2uUCdWTLHvznfQLws8o3
Pq0Mx140MGFzhZpGrfuPF8XJ70So+046YVFCFB0vl++kci+m/E2KFuI9eje+tgpyNdJntKYaMqwa
axjj0sPlpVKJ2tnpbzzG7ZkMEjfJ+PaUNqL1NhOnCGj+K3PllFBNHPQ0Pp1PhuUvGB7zL17P1V6s
cvSUuQ5BI8RX56oD28PZUIoXWUfrvu6ZNjZeqAOjj/IfR1D2GflFtKaJZKE+rRtXqIuy01rD6EAI
dPJfumRPjFbZ7kReSWOchUoChLHuy9RhwnKlLa8U72V8JcJMNbXuiTOe9jpqgGZK25M61nuAhe5W
Ehf1104Ih9EVQJSEUIM+7qzdHaDAeWVzcOKzpz9GBMtHcG642KiAYz+wPrxzaUdU/yTlCvylShhU
HxeVMUq2pVXkTRtrPela+qUca65l8Y6Eq9//YxJxmW22ghTUI1CCt3NL5kYmKRVZ/NnliCzUJ95e
c+mwhiHAHL79LO5m0ofpyhFrywb2anghUDK79akJlEM5UX8WCtbuvrpHcLxsnourYH1vokg5bsQw
KH4TSPvZrGPNrE9EHL7ZisXzXenn+IlKjvk13N5tNC//E4i/XqzsdM7QjWxuAUt3FEuJN1uaAUY0
wS1NznyopHaBYGgelfutleoqEc4iLO5Wa0/dGFk69ab40Vs5aUTfP/V4syrEwmubgAEpkhMi8hmY
XE6G4wX2tKSLEX8LZyEgQrsKG1xEqtSYFti64OgU+w6aNBUZrxQXqjRr5ML1kv0bgtAyUtctASRc
zQy+PAG7OmW3wqiFd7aHPa3o9HRyI8uokujYYJSZUNuc5tVCQb5cqVrqsZTKpsnTDba/fDNYd6Xl
JVafG+tMD/RINnBnfa69OVz38GLQWs+VtvVH4XWb7tHE0uFr9Ik1E3jOAIKT1nnvivCnChnDFxd0
8DQvEgCDGmCdtrBEdHYNcBBz7ySNJW6Itnw0cZ5294GRit0QTYbXe9kGd5/XnBXnUusxq2Fk6F3M
JhkcidJiFYOIJIGLNYCBrDoTcMsPzgIzOlKUD9EqlUVoZUQEAFV5CzEiyM+4/rlNhevwzz20wyKI
EkMVtTdOsPFphKQ6kBdBwpB9feVBSjmTypzewCA5LGw44ebNShGG0L/NQuhKwi7uX8RYH13HLGbn
us1XKYtnFgCFXTKi4admy7yVQtYYbvmCVzE0xAbE98RiqpRZnqbPfIB02WriH4nvogb3oXpXb1Zw
lJC2XcJjgjrsT3dv3ePcrTAIQQpVJ+Ab8bOlTPOeymuM+c4D4hiH1n0bPQT/1tNJUBHeeYk81bgg
+/DC6SE/LK6zhaRvLI6AkKJrxLq7dtFLjzbiXQRVMp0+SIQ2H/IZ1vCETpzrMCg5gB5eKCBzKpCA
MAgvRNdNw5h4diHVPyjedwt2C9QvmCrrdmzORuhe/V3CR7fdOK+NBTRkC7TVY+DhUXl1yW6lO6Ce
1xhQ1fiWOFJ1nyNqRl1jBUI+Sj6IfTS3JO/ebm7aHhVpV4d7s852KjWzt+a7GdoG8ECx5qjy2imF
8tplR7wSvzPU+6+l60+vK5YE+CA6FFfeQYJtkZHkb3RHTU7lyPzEkaSjM4i7rL60eo4O580Mw0ay
S8cG63R3bvtzQIuF+3udDAckMgjGkx/qZzKf4il8M3bcU0GA7xZNDj+ChviwEvXPYzl3njTFW/Qe
VBMIOjmTV9gOZhAcx1AmURXT60E5kAAm04wehEcGsJfxy4crHJ5t1rQENr758+P9ZHwJLMRucoIP
KJtsV3zplvzj0KBoHhl++3Tssrvie+UIU/1gXmqMFHFy91rOyZmykqpItRrrtXw5LWzcvoBG36Fr
G9kh73GGYVu93IONGeSe77L7LUugXj4eIyMzMvPgTokHPzHYBOn3Ns6ZkoWC3vgM0aAcnpPJ2meP
D7vfOTjZ+iZLdyikvLo/wBUHxG/UbhdQo1uuV9gTAZFS94RolW9WA8oVrWq+/NdHmRxxWfoenFW7
nf5KPHBNGti0iCp4tesXw0NX8c2f3QUWfdjDWhoGyzI4XUk5PBHBputPsD1VDUb6lIcsyy47FYwo
ZI9aIMBilI6Wc4eCOa1YGSCiNul4LzlDoysNZ531WW6M4hTtmMzjU0tElEr5wJ1sKc+D3EA3JqjV
MdclFgssjt+JYXzbsrQa2H9F4CfX2OlgFG0PCSsumYH2blt0cy2tEwmk7jbq6YCv6BrrrSt1xWfZ
jD0WqGEhqCJfDS+G6IjQojzuclZoFMFetEKK4psyHVqdWiXdJ7YcrUiQsGGg/nsaQH01vgulXqpF
F8mqWEOzk/x9/uBf9117N2KKqn5KUDbb4ZCtNwRBV14/Z3cu98c4+FACRTw8jzCVIR3/9LuiftCK
WY8VHXlhWOAH72PYI0aTdjMEsJbqc0KxK5iB0YNcFGsvYNtbSQRLqbHZpf/JsCCdPq3ol47RBYqD
KWE2EPzlC00xYLUrAb++PhHAdb6UYAva0Z8isrb4dHA8BmKbcNJneJAlXYWfueaKfh370cG8eCfK
66k7K5YQd3HEqNWpRxhT2odU0aGYm06N9rcE9V1VgYehyKB7tXK0rXcfOSXv5vZqbQt4oDeBmt29
+VC8FQoAEw4wD7ExQFVf2QGl0ZuYzYbJ/lgB6WbXvn2UfTcEIVau9DZIy8Af/NZL4oc6SK6BoDcp
pMgWnd60YbQYi/UBmyYMS0AIaHEH5lNrsL9vunrFWSsFci+yeScpz8xckPNN95QzL73HLimDhZ+c
R2Epimf5dEh/1opl6w08S5zJhlBZ+JM1M8wI2jkXf9mAZhkCrvy6wD8tUWPQZtUw+S5bbl9ZaDvD
I2FBLof3OwtOAba+GOWhNftzRH3KD1qn6MWOzalphai9maEIJz6UjBH/gXbwxGAw3xCLKclCB8qV
jLAxgpNnnNB/BQjp/J+njBQfcN7cDM8QzVpqALb3aM4epl7DdZFQwlXCAMCbj+Q8OoopdFAh/ubZ
UciYvNC3vBA1PIm/nL9G5eZkuZVbwM6U6FMjh7D69xE7/gNncIfKJcAzZvDbDZ18KYm30FQ76Ymr
gWSmA90jITHj0vuMAczGuxa9wcvgx50jXxYNgdnjYioJjptQ+pisxvSTCvtbLfWRw404ojjNBIPA
G3fvZXkrUsR/lLwNmarzKLByLwTWrQiEuuvu7LgTZPrYJYxJSBuat+Jy5MYCTZtkjs+xHgfpGL1o
X+552dHLM5Rcpjt4/SpYBLomqgkvwpCLUwS91rpZV2Sf49rsafOY0DzHvlV3yw5zuqah3qLT/gnB
+FmngwbOgvttKup+HDMPsG9fBrOGtv9EmnNyRd0O73/o9F1mMe+DKYM/K678Jzj9mmUJaHvpC27g
dlQhw7bAi0UPZonQ+V3TDE1+58R+uEUawaWKAYgvRvcmPvpHvr8UmMTvRr0ToeYSM01zcvZWUVtV
ZoobeqEvuKWQmiisRZdi+GYxwxsSpFR4QAgrddO/5kU/KXqJ0wNHADi2iqWoFwPaQB+lqQON6sDj
bNb/bH/YLexZuut0Yw81Xk+Yt7HmBGN2F79f1G84v7jrE1g0x7ns2BlSeQvN8CcK1MfGQqK6ELVp
ISXSvdeCb9zo8TGhdLrnzlSfKDOV74VDwL5HKmrbJ84ScQPfMuzeFJbawp3Do6+bQxcv/IKuLZMZ
Et/hHxdARvCp9ryKS2Nc0njwmCXQMwrg11HS4zBJ+XVgYpkCZ4rAmy0biXPj/EW5LzXUE/9wPPjf
y3z9xqUv2BJKX1bpnH4/4XdjP8kH61IUAZ/Ga7Wo0wVwIglgH36/qSC0DIvrbK355oSGOgRSF0Yb
bphkSnofmriUg66xJol0fGzxpY6/4mBCu/imwCVf7Sh7VX6AzCh/8b5V3nIvyaU33tMMyzVh4TnG
nS2COWmglb5uEYTLDZt31Wh6RSuog1SnhrSQXVFDMUEKQL55rx/+AJDcg7EfkQM33OPfwmKVENpn
asA7TqqJSgszuM41d+ZbHj6CA0dZ3aX9F9cEFuFe7hFw+GV7x2AsN7NXCHWIqHnb+ld6Jt7R2keX
KG5sRm0w+HQSpioSHoxxRIvdmNQGHLL8deM6ft1VuFcGC4BnIJMwT6g9GRougJ8BfE1zqS7wiMww
+3huqteLRMlGSSUsE2iwxuUxLc3FiDSe7aNyH8t5H6TFw/l+Tl07zoiGw2Qltu9d9kvf60EJYy0K
WSILQn0u0ddFAwTQLUmOKcIJ6s3QjpjFxHP8VicLPtC5WGkv0b/v/8bqhRxmZT2A6bfpkkuJOiKC
7RGJ7Iugjhjny2jQE8lS7jImJy3x/ZGBXYjMD85ZeAFnPE8QH9ccjpLAcD9iJLKcYfcShBbEWmWr
XYb/rcsa1JoqAkDWsT1cM/OcX2cJT4Ovbnau1oetHC9vPvgnBjFAOh5p7xr6lSXw64DP/ZtODEaQ
RtHWtG5Rz9sgRuaSXtCYoG6sEUebdxXDDYj9V1b3mOAJLJbYM5r9Qm5YLKQVTbO8zndc6ftK0v5Q
SrNNAvIe/P/ocpGgsQA8prFXw8LXHRwwbDmu3bMZ4KQW7qd7iWnEcwimjtgaB76qsjUVBQXwLEMM
/3vrDOdkdx07+58tT5r9SmtKOBuV0zJCO+zcQw7w1FbzkYkBspvBBiXWdZFrIIMvhEk5XVo+Cv8X
lfVQ8y+Y930sN3YVfMRWYolhAZAL5gL0+8P8/fEbOxln/+YHCEmZLPvtewRSvBY+M3tk1pTdIL2X
/tYF0r/7EiPE2ckxqGbi+Q5kjtv4x1CN5t1XOjgpL2sfGQe3EP3il+g75P7h+Ozg3L3kdCWJ8WIB
dTdVyT0CXPpjYfaz1U7DN4GpC0Hi+Wz+bUfQrCtFzXOcd3yMHy77x1CiwowCA47BX0fhtdfphj/S
q/e/9YFolA+VU0FqFYUc/N7QuDKn3zbfV+GJCdYmG2t2DaI/L9xAoYQB3hfqzi31Na19dN1lIl0v
6OJUkJWIb3opJqLNkNLG/6OHmTy+5fUMwYMg52tb+uPhZsXv2rFX5T3OJHYFZ0DXpn/6N6+hc8GN
wKh/QmOXgBspBGCERBZZttQLLe5gdqeHxVoKokcdQo9uShyafJkcR9Gei6lEeC2BzyMwPqp0zeRR
8w5c9lrhaLFczytKm0Krk0g1e9e3dLYllQtihslbBQp7plVpHKoc6edheGafBd4sHGGLaRYxUtXs
NdJ+nGcJINflJ6dlQG4DplafQA3fCcMiBzNcsNj4LHX4vee45ouXDAC1ptFgJU9t9QLXFZouGBhE
n042o4ZRiaAmzcqW8BCKgGC5IG5IJUITkgJSZUyn8fR9WMUf32GjYMF49YJRP892BfwRnQp/63hj
BpErm2Z+BOmBk6/pc/dYESDvhv+y0P7XVroM2twY/fVdD21hYSaco0e/376syAiVgQ+/5Gujspui
DdBnNVvUWp/RyVE0QwdrYqBXaCbJwac/lZ5NENjQuu3icFokOXuYWyhDcZgo6R0ntyd5u2wsb7CK
uYKHtrObTCo7tymLehPESl/49J+IPib3Tl5I/C2QVTVAMFEMWo5vlvb7qLQpO4F9FRiZTXU+mSWG
GIWXFcqqSd/PtvyBs6byaTjPnYNgVF6+ihPv7tpIbJ8pjshkMgOEfekPq1PLzX/5lUY8rCo2PeVr
F5ix2Q1F9l64EnaBl8Onq9NLE2Kgnbh2E08S2lv0kX1beaQB1Nzp5RhDdjsTE+3FajVa1SAYnlp+
nDOd9Ldao4obQH+JQXlTcpgU+DKbPXpJVnZRWCvOV/7CECrQg4ZZe99nhYcbsPKfevdBdQUOB1Kk
Ao879q/CO4Gh9wgSHftWWmOskkZN+/gBAaGmWmYTqIZirJLE+1erwujUKDkx3l2By5v8VPD+6gRH
rjI1rsXXC+kH070Qm5EyzqeAUJepBANf/s6dbndXWzM8OzRs7ubOHZmmmkBzy+bf2BtSwFF2EiDK
dklQ4rXV0HsqcrmiidipfRCX34FpNoVxfjtpOaumaDSU3/dh0MCdb68nH74oxZG2MFMcIi2rUyAX
tlVAZIBe1SEnlLNd07Yz6BybQXv/mVx8bfO7rtZQQgXA5M+O4a0YWyJ95zs0yktgA9jbI+Gh5LpX
25rV+0pHk6DGsx0hEUkD9a4LmAb+6XN4/gIKSunalGL+n4BpEzszSqji3bv2BxuYyajbunZ0CRSh
ODcD3hPjmtjnNnjpk6cu6chhVnRDSlmOqDjx3+Xt3/5WxWK9bVXzCS2QSyizS1mURWydd4FugVR5
tFLTsqxZBPuYdARIKwDJWyb1oA48ROx0DKYYJeOUY+GrVA4zfHtfAoq+xLhIOwtSSlcmslchGDuc
9VRvC3zcGtGx+3lFGP6koJoNuSNAWp2N+cTQlNGBoEWqUVsdHJzzb5yOPZau3m7Dp1dJYlGITAFN
sMEuRmZUG00uJstJbZrdJMVob7nkVsgQdT8k5sz3ot03hP4UbhJmbLMbXs6TnkY51yHevcXXYGRb
uZyJKTN89x7k6uMbE13KFWU8CXbpSZAWj1loxj8dR1nEekY+XbuJTDVJyDZeijJ9+Is6cM/C0o+9
CvvnMIsoEZsnzeumv6PvwzgzT8SRrFNWwXeMvqztqyzkwy7mwLzNwcy62+noT2qFS/lpgw94PLWo
K4jJ2Pi1rqE04wRR+eGsf03knvF7nXWoreaa1dM4DbSwKSDD970PDZuq/il6BAAxdG7tUSJuMmb8
9Pc3p/HzI1z+Ip6zGSYfI8MLGwM0XuY9ueB+Jg6br7RcfVZNyy338Vad9i1LqL61aimBHoCFiKEb
O7IjhJ0oAsid2+8XgczUXg3xta43N2TIlaqcfDQU+ySU0MLMIWPxDhV+DBoTQkgD4n8V6Qb045P8
PkgjcUqlYXi+EfLOOOAZsvbOlLiDptA+2/BGoepM/ZaHFNOvwz00tXhtTc5J/spFbnO8ApN63mwP
0+Jk4ICbUdoW2s7ezsghLVn53qTif4H6IgWa2eTEFxcJhd9zYD/dfBR8FnbDzM55lp4BVAU0DOqX
WJeAlRng4t2p61PAt5z9C5rw0ZSd8VpkktBz5hGJX+nY5md0YhENF1jQGHMyMSLgm9sw2jFqcLB0
/PzNSI9jDLURy0uMhb5ZnpmcK1fpZ5DzBvJQs7b/OPepTi/QyEq1UtLf26MD5smRD0qm3zegxgTy
ODJWMu/SFQRZbgdMgvRch2wF36nDwVvJFK4w+dLY7utQGmWRRkjFZFAPy+06P1ivNUPqdx7jMdby
mKmGzZk2omIPHIxABl7o7dzH1+mH8M18fBsIt3lQ7QCQuqw7GG4FGbXZyiX8s0Rq0GLItZBaZ34X
hNu+7bRGr6vaKYwR8NbPiKd6PuS/o8cpQPVyB/S6os3LGZcUdrwSLQb6j1HyWp4UPZDVcc84Ng7L
bxY+Yq+jrpW7/6gbGMU1jCLyZorQSNT5LLqIAKwF4J/Hh/Bn1G1ykKmqXcTP8WfbMqysz9JbAF0W
qwTQgj6Lf+cf2nTjrhv83sjzhfLSqBGHfUe6ngG4lau5u5IUZry/fWSjQIDxacIdTWQA9ah5ZwuD
z9YW52zk91weqmK3fUFbIU6RZO96/RDnemGHrxUpj9sjADqyluRTRFsANMRDmcIGODlFfWRf9kOl
Gw+inkmoCgu5viJcMNi1zicluUfeWJsdXFMgg9dVX8e2QoURVyNndA/npDQ+MKLvsnU1zeTemULi
MLg0aIlsmBumMbqCx/SEkP4DYY0e5Uz4hgJi33TEcWTmWlm8l9UEt7INeNOhGFbnAf4kT3eVMrHh
4in7W0P7vwdm2Qg/Yw8LYeBtOPzivplwzFRJ4TzzgmHnunigPq2gBAsToPc7HhT236tvHgBrfG/n
N0QSRJHdKnnGqSxg0g07Ywk0+7zJudmkIWx1GlupAjRUdVQO83cnCtd2GrA23AYRhjSI+daH0NHx
2j3AWACNlHEFGsQ8Wt287eDOXDH42+FNMVIgfm3EBBruGIxI/9nUEcPWi4+bHO6EsN9NCWPaxIlJ
nMZhThl0WplSbvCzmqEqV0iGGDnrhezJmvrJo4w8GsCaY1XYWdM8AmMq4OVa5VUPOGC0p7HxQQc9
KExvzhgYBjcIhoPVy4eaxmhEowNzbXIY9VrI4hZ4yRUTjHWrAgCWX6pfcn696VqOBIl9gpqKqjTa
6Q0VUmiyrCaGHEV9exRj0LZQp/REUyvhPt6OTsHAoiS3rrUUcvLkBOcNQkhHyOelcgJim67TGtDi
J+jVV+2ilGd5zZExTUuA8n+DtxkPwMHCwjj5ZxtgNmAOD+Eb8VHzH4yjUQ8cFayw2hNjHKI0nzqL
UxNb4o8BWfe1PTrhZbjynUxIFFMQaX7rb2aHxv6R83oiCu6dJk57/ZQode54sLl6ErT9VJ67iTEW
IkXE8S9Kwqmbra2ZBA9JAwSUUcsqsN4KdXiZI/r4BK2i3cxTd43jCUjR2ad5dY/Kg3p/o7KIxFGY
np0o8fSxFutcHdJq2d0AeImPjCcRdh5MNO6Tn0G3hzALPyIazIUUU3Jxf/ReWJ7lyP6w54n2G3Us
7nh2VjxaeDqSMAAMxX7a0dBeLJTfh3K36mcDyKnOaG4NKUZd1GNJT2u72uVl20SUmlenpLJ08biD
V9cg876E+xYT4vNOcnCOy1A3jh4XLI3m2UqpbjNno5rmcUXEu69CKKQ6Ifu7ZVdAb3N+sqLdUQkO
34tWUgKHJk9BOoyO2LQ4kT7l57djbe9KK9e0jDyMd0cnL//uNshUQZ6WZNtmpcAQ4dG2uITvVhyr
SirnV3yBV7I2DqXOliMF4whYSgJ8dkodWL2TTqfq+C/cRgfDGCXN3mNMdfxWa6RQCdYNkKnlVHDJ
N0BYdwu3UUxbY/WzDVoctmGrjV4lNjg18jU5lmDStaVsLvHKVM6BACy+hy5rgQ2qTZVWsU2SqL8a
GAri3EGHZe1cr0t80OLHwigNyhx8opgev7LsGzsdvXINbRoKNHOa+fRVKnp/pHtzGMTvMkR+iszf
NiwJmwxNcPhTvwhy9yx4BFUdW68nq1Y4kZRwapyW5Iwx9dE6AT2cdC2mm/a9Ge63g513B/E3S4bD
Wzhb2+mbIfVQvXVjktQ0tUxEahTnOQdqk7z7wNEOdtWfcjwq3LH9oENvdqqo2zvXZEe3C/hx6Ay5
fFRfS1JGRj/LSJG3eNkhl/IeROu5kUy1uqKgvkKXgz87a07tHSW611l8dPFC8CmKdII64quJptXZ
OVG2pdLeZ0t1EQGVMSR8OefIg7Jv4s6s4LDuCYFf+YOELSR5rOg2jKWFq0VE8hAc1zOM0gvaEIn4
vXJynhmMt9AIHzgLVU4/7+HbNsn74bQbS2tOE+fgl2C1poxPQArIbwTNbdP6xfyFrE/gQ6aIWXpm
lucAMy/BeKuI++6IDrCmeopFHu2pcx7sXu1qP+1AJoxiTLhOUAQjvI3+cGVGm0t8XdBFZ9+Ys6mv
fGnV7fRejlFJpZ1Peoypi0emwQD3lRsMty3dFJCupsbrc2a3QBum/AI8lepuEjVFrJOSNFheucnD
mSCRaSJ+/ikDsNiLkBym+4teiKs4JDV4RR+QEpimubtHQYxm2P/af1LZLlWW9SRD8YcOzpTWl6F6
kl6CRmNYlVlRS6CMvkRoTLIFXonnPnTtM8NKlIxEdhxTC6WotcumXjwAEKNH8wl8AGqp3ev9Mogk
U1M1VNr0m+fHzGbDW92RIHXMj0hG359cPz3bgPB9J87K3IfPmbLl4RaKkyepJIxH87rRqiciGn+V
C1Fb0UWsQ1h+QX8aY9HjM5m88thgq94TNrWDzj88uk72mJYhTDXds+L5NqOZ+NCx4w4h71tobBNy
tX4YTamhvXDHNPbeqQVQVLilVHzLsVaBqA0ig6YJaZY2D9XU5ubySQUOC5BPeQ8+ZLmJbIFTe4lg
ZgUJb2jOn2LFDZFO4W/J6tkz1aab2CEO+QgWv/P6KW9IOj97KuiAYY8+kTTHH0s0/Lr+Y1sOcjiL
LWZ5whxXp780PMKwm9Qq7xt35bPKTCK5k5zDtkOmY/0l3xy6e1K2hrqF/absg83bcAOPVaqcOEC1
WNuhbdWm2d1u1K6eCsqZI0K0RKaQ45WSeaWHYCB7NNbAMuq+wH/ksFXaWF1TEmiuyVXPBpjHNJyR
1LvchMHNvrTuXUv2UsaXsUcK6jl/PxyKTLcRa+2F3l70njIGuJPpeQXWhKMAF3YHS4KBVUa7TdF2
dyv2OH29iJ9oMKhGdiZRtfWOBUTF37Axa832nWjQF2KQa5FFm7f+Q4073DcmfeQMTnGgPHYUgGKK
f69jCXGS9vobCsFs0iuYyXNS4Dg4u/RcNa7Q2SO4sMzkd6cRUwpKYV0F5V7r7LvmihMg6Pnps1KQ
qxbs1++DWTIv4Ngrj3VAPH987kEQ7engBfME+GIbw8C0OPow6+j+oi8U1UvybCJkyj9AuW7CO2/F
uyNMf5SsOxbWP4yT6vQqQ5A5wRXgOWL8y1yaNDzp5sl7v1XyNF8luTVWcMqJ8lJPjoQ7x7voV+my
oxxoAZh7EdBqjUSEO0va6t6FqE4TNYM7VYWU+hIvS6XHfxR9yTtTMr7nee0VYzRvAY4scEcavp0t
xwPt8JNjn0xC/ZwMp0y7+nVZWCC9A/lfsz5ZbmMGW+rLywvh69QIXhsBZoElvy5zh2tupSf4me3I
Qglaz5AP5cIYlZNve2MGLF7hf9G34giDaZsw6HiJcG/xKvNIyZKQaijVC8QWbUlXTwKLbR9udk3Z
0VK/lqLolXaAQ3RUreWsfVSsWQY4v+QqFV51mR2dKt9oZ8W6isWcV47NWlelobTzBhthjHAzMrRT
RggtoLidQdbKQZANNtAHk+F6I5h6kN6NikdK8WrnjXt6No9SeZtKwWHOXa4mBXNBXxrUP4CIVoP7
UmdhsClXPLnoA4AX43cV5JAA0Y2p0AI14kzlQTrnjec4nPnvvnaTYh5JYQGY2sxsAwulcJjxbfVr
/blJN5AQQnVQiAQCQuw2jEeV+SJeEmk6+F1rdLWZY1ghT43+da9JA3bw64Czcxe0RIwxSwHXIR8p
UfMcAHHfAE6WuKocpuZ3Fe9GFtaT+CKpLmUNQ3QM4Ju3K10OxVy2uVYqInVPt0eRj74H8q63dlbc
d4nx/111yyrEcyVT5SW7R/bdlwxqBimuhCPJtKvnNI6/eMhZzTOoKL8V6CAI1PAI3lXnvAk4WEO1
QZE7jA25DXYLWHa7TGRmPZgVRbZSGI3GL6HOdelpOm8HOPds94es0SLmnoW+dvG7J2Cnz9Kp8w8K
rzbDVx3Nb+zHqBmgZWMsCa5+5/7vFnDbGZfiA/Mcx1Dg3N8G2wFm405gLBdFxJUBuI4J7Ql0IORN
PnEgnryFDvyH9rO+RGNyMCmTxKAzioo7mLxB/PDUeQda3t+O6JL1nHO7iIVn6VSp5L3Rv6/NUJYT
rqICXFgfpeLWF7EOEdyFF2CAsBbDT5q8vnjd0q70BQFj6VNUh8VZJFHACbiF41zRsgHefOSw7cFh
YaWOnChUGUZw1jWwDyeeCAyHsRdHxKIA/sqXlxBx3ipxoW/EY3yqy+2Ry7LUHSXkknAL2hzT+Rwc
ouADpuHBdfSoOFYRypZhILfSsNhmxmD+sWyWV1hxOPq/kdZzpB+jua2yvZS305ReACIu5YL+S2Yo
/GHmLfDBiXw+d81+c99Sg9ZoUfb5Cpr+j0CNoETjGC2twglJsFp+tMsVWTSAEz/qutyGxG8fPvE/
WjatWASgv4ZkCRkCLOcORGBwVIs7wwd90bVLDBc8FtN217pALuG2tw5TDLwSHiiZMCcVP30TFk4e
NewIYhBVEiWcEmMbgida0NXV3Fqq8NAtKyf2NBNvUc6c2fO2/PEquUHktN320gcbQrp9CA7Wr30g
+WijbYLQypk4lnlx8xQ/hIfK3477+FYpCPYy+cLKDIKYZPRwcBuRS44qauFK4qn8oFTNaXWk5Prr
tA7hmKUf0Q5aZb7jpUXEMnvvQb3ofyYOnEGmR6jHpfxn3GKQn5pLcG86kLthfIfvZ4UK5yoyyX1S
Ue0DRV7LWMDJk+GIvPBs53Y171tHfgAOv1YzzHmWrXaLGzzzNxkQeqdRcAYA7DmWY94rXnWHGNXo
y++S0lU0bdk0BDqLEhKwqG7xF+wPXlEm2KekHO4ePn0CkRtSje4kQRNdO9SeWUZBOl5sUh+hMu3R
pVuZjulExSJfNCLMidG3ce78I/8/7nlnFASb+Amorqsh0YW4I/Zpvuf7zOXPcu5q/EL9b21V+i1w
Rmeo/0gnOY+qilrbphhmKKNCoJo3NEpueqNBdOzI3qcq1pkMLBNoMFd4ePdL8K6accfxyIOejsGZ
rRUAdIwKEGKIgOpxFeaui8JYU9Sk77EMl1TaJ4ETkw02Ox66yVGZV/wjTWsu4YwtHMq8g2Z8JXao
ODOZTsCjgSovMA6TWfJJ1vSthP5h81BTizLhtPD5phcuM4hGZ3WNWKvzAPbLjSBucr2f055OL6zx
umBpLWNE6UTjgexIkPmP9QV5NRpUCejo9V3E3uaF3tL6rlfiPM/biqAqBE8dcvnp8o4NLHcwjXho
uIT6JPNc9w1M3k/xNhHYSkwPLHiLABp7jmbMI6ZAFC94Xrl40EZH9uJwBG23ITZAxD7ww227nkzO
DG+PFzv10Awdn/PgyHLp/hC/OnwkY0uqMyPknCJ0jy6vdysyP5tTPI9bFsniYTvVcLG1yteWJiwM
xLA/77sOnJ9o5va9NcnrU0WkYGy7Efy8P1Ee04G4AftXzLRY9iDhKVVvSBN2qjn8CIRwI0gG3x31
lYMpEzh4ImLzJC0Xyi3XdZvzAQJStQIb7uevTuUxtobuCHFRTc/MwypvNrj9PiwN/dzchUby8We4
gMkdS0+d11RWexvgRGEgRtrSdRox0zHS7Jble7Zsh5n6NNEMbBtzIbMokiiAPkiv3X5sMwTEvt+s
oQ/vk55Ih8X4XJS5L3F3tgLguLTeuqrS4U/uqnTDpFIC/sl5iyMVh9Ga1e3SjQM2uHvraJF/Va7J
7fqN7hkIkLHVF0nt5vlfMTFFUHsa7eUcKi4RKtfhSZvTkHVEg/cKmGkWyvFBd5JIDJ+f7jPGL+c7
oINJtSLyy9PXWo5pR11FbhTqUu2lsQugae+1iUDLLV2eTz6ko1m/qXZrF0a4VAc46XO898ft3CyQ
PwmUe4qWqWCN3qEoVrZKZRHOu+l40jt1t1H94zBPVcJIZL7DtPU1/PrdkvpvtDPRmpsrV7/TYa9S
RCFEiTzsRpWN0/ZN9qHSg56RzZ6B7XduefZdnjTFQ4NTVqxAn0EkXnZVxW1d1YvahT9XhvfXfzZC
zulKGlffuvHlFrBDQQo7FeWC1/zmFfEJfuWmIfJpAuS8uinIzT/7uzxYYy7khIkqOD608gC7H7jg
Cf/US68s5UUArJqq4QAnhGMarr71jMklS+NglRFxsjN/fQv5ZmdzbnsE50F9j77JhS0nGQJfhpKv
w5TdAnOhy+bSQVx9dcXIERKTqTGnMCH1PsVbTJrRB6jR4aGeP45hdwE6u7cdl8oMeBxXsmvdVXUm
6nyyqz2QZNDI0nCU8CfzRghtM5KQODp9eiV5so4JR+aInpdaulHc4zPBWnBOFp2TQsPN/mMH7nP4
7ZHYMSTFWKKoRhx75jrRA6jOTOFdZPd7zTN5nKequoR54cCRyUJMrrTw8jvPBSYIhQWrAvUe+51m
o6iVfEfcCvbPS0ZCq/y5m9SzcdUczZPjf61k0jxQ3qqV6lrzHV032FSvoVAjiDlKL/ATa02L5c8c
CK3Co8ubne8yGR2RxZ+rfJE02J+EiAxVvzkLCQsj/mE0jI7xoJeuJWIhY0vbEZp/vJ3rxRWxKcBj
nnhzXoE2hRsHR774UYMA9SaHkO8fJRVV77Y7tZ8mMvGcRC9m+wLGpO4MX6AQJGXcp7K+REAzNwEy
OGRTVsIJiCcD3Edck0IMVkgHBa2/upX19HdybYyvi5XLwSeZUv2SEhC9qmHrBZ/o0UD7KmYGyXcM
5jK1Yal6gjnTvo7kjcDKGuhIKy+X6jgjcUDTZBj+qD9sSvdLP/5IndWUVzoGU5SNO2UEhEdIU888
5FAGsUou2MdCTHRjihY2KU52vBKhZFocT0xnd2dsjnM6Wxs1Yc5Bjwc8JmrexaM3bYR5FTLg128t
xzlgj2/5abDyh6DDCtW2tAzVbObd5cOOFwLZ9VC2a/F7niLHqDBuQ3fP5imqthJaRSo6COdlNfMw
YwHwDZ6locKvWjAS0LnLPeeyoB9mynl6uePlIB+N6CY8fViuJk9RuKA2DR4Cuppwrd7f0Jamax8g
aMONI/5ealsXBYUzV6fO20CgQ9Qguh60c7xLHylI1AzKch60ITlvMvrJFafk1PDo/ILDGeBoZ0uP
qm19abjRvAkbKNgl0Z03vZ/+gLc9Q8qmO9FQjNDUMj/HjFKiWzuUA9P+gMH6lV0FWFFKXIUcIax/
DSswjetfls1DGiQcXB36XUgqVe5NQVHRvU/WPt8+vKUCECIYaJWR+V6Zam2WKJpTKyWr1MfHh8qv
ZQc5pAusVQQgb7JBwB1w8OZ+5ym4dIxHkTIjvxoTDURZ/LKTq8/tE/DyG2vkA4f491vHeaW23ZEx
GtkrUCSEzSp0XxE1Gxc1O2A29nHvEnWgmrwz1frS2P5arxlrcvcFM/1sWFgYBRHcGtlAYNfj+HWG
+aoGMVJ3ycdSvnZmm8idWr+qFAbD415KgUYpdjySgETrRdtBoFhQscvBp1++83nJruM5GOxjVubG
d2BvWzW0rIn4WamfIIZFhr4vtTO35nASOM1loS2xdhPLibtxDB0VWRAqgh5wqDJGpcDDZoiBEl0e
RkbyC2FXZj5reSCH/mfMVndm/g3oSPCLC9ZmRHsM10YHX/hgUUNyXM9Lr7jTU9+RUfU9kVvxx+l1
jwT58oT3YmZX7lhAO0mbDDMUk+57ZAFz1Khfmp5A4uzgkcv/feDMtkBg/w3Cz+1YqzYzfpr+fkxG
9PT4IfyPEmNHXR+a+Ta7fkclpKAhEW37J0Feyc6s0yIi47nd7++tmNJ35fdIgoTVp9wZ2kmOeL2s
GenZyWVcLQI2hwhnAiAVeryb0BdHQXSnw8eMHAVSr7DyL4ia0Fwkthzy3UoVT9IuWANYzKWdRYdF
7IyJt1uqPuU4M5Rr0gEu/HWCOg8rDyzLuMB1NertpHsI+FfFeiY/svcJ0JssETy3x1t5AAglYYpr
jpxfU9G1yBW45UWZxL2t0OozgWZkczi7IkZPxx3vQvxXiokQvzGi/pmaGy+fd+S8MJVRxqlFIRcE
AQDIRTIrxefcroCndaMzWbZ70fQlgDORmmGlBd1G0Vm8h+2mSbMfAgB+IKwKmxNOeV1orcL1gCVo
KdAmUT3j7Hu/gIYRPL5itRxCxFz4CXFRga184w8TH0T6PnbPMuboW4C32O85ApIxth9Kjg5toTMX
MwQEwWELeLN8IpXFQw/yage/1TDk8XDOKOZoxQyse3CW8X0GZG5fVNayro4H11oBGbxtPMack7W8
EbhXWt9AYFVRxs/HsDQJGPl/8HwGWUDmHJhcrZTXq/cdBGo7gtyUtviZ3aWefrtlYUJZIbKu+c3G
Tep3JomkNYYho5HIZOGtdqDXOZ4ICgECuwezTTY3dojba8Fn0fa5JCYTPhbtqQZBO2HGVukfG6gy
D+r6mEBSGU/73kbNa/iOObJMTM6g8nPs0tceHdwtNB4waSThs2THb0GrRQWDpUDoFyfV1HYfH4L2
p3V7DxrIYBGNQ0iwUju0tEo782mm/WfdtZpA+oyRQCLnEjnyPiC22mYmu/K8++y2DCLBNo5KwKOm
69s4YXGQKwT/M3nA8rzrzfeTiis5qUg9tD4HmQg3uMgMP/7YyLKeSeaDdxTIPLsn2bIsjNwxvxMC
Z2HNIwtTl4xhG8Hg5Yu+Afa1OPeQ198tHovet+oMNWn6MtFIvy4EC4tHuqFLNWhu37PrdK6YIqM8
/QgITfpivoCGEMtEt/xngggXhM2nyi2vSIB07EJejTE7NHf8MBfeb3yh5RvJj2iCgZmRoWSEkgF7
e4SsBh2OpD61AXIqkMQqeptRV820ErpxXf6Jt9LlzKJ268KuIUPmZoMHbqlHQ3XSlO9mzJdy/7eN
h5q8Hi0FkUEEP44LVjlOoBD6SW1y6DL0/W+9JF03FTpnk/paFlWmcVw+vMMWMMyGgC2HDP0WddqW
T+qb4+OMCtNXSxIqW1YdjlmvqZFNOnQdsWA0qK2hmr4NSOczyL15kr3DFGbfXvHedQ9f8+QDqgct
VlEIaDHm7a+3QjoDWwt5QDylN2lCVuZUFih6uNGDTsJGRlgJF+8OwQ0tZYBgGtu0gqtCkj3ZTX4+
r64NIU/2Xh/PEc6HPHMSs02aMVcCleeIH6Jwhk6bKGSFkkixfXvNlBcdpcPdGrJFR6NLh/NLaE53
YFXUqIO5JjTU4HM4bw//q+eO3YJ0gCllqWZiS0ml2NTUQbouK2JdycmbEIaM3kqVZ5Uqq5qoYV3w
oSE9sISottLa3xdWupwxuJ6UNT9goQbbYSMeLlz0irVf0BmVmIvMK7jG8M9btzIIKQu9E0mtwzdO
fACgIT5kx4trcq+AfLRSAvsN3d/VZ0LEC2/1KBWhiqR2s/BRE/YFQ90NhaACwxmxY67KMCDVabIP
JO0q9dtJnxLtelOdHyRNnuYplUivdsw1STMgPN1grdYqlUg6EEpiRaVwKg9cQ5rn6blfgregIj5K
65cfUxaT2flBB9tpXEqo174D1aV8IY2yFrayYgcGVtUxGiOVHrYxEn2wDLT6ydhvpCBhTGA3gDwo
+1QiWXRNQQ1YF2nnVoOCaJgHRYKsmlsLQ+5mVGpdfGyl50pcNUks/bPMYNrr+kgIfhxISH53BlD4
dXburO0I/DQTKPA+wkwN+/+n7kj1Nu7eGJRImF/TbpPc2z+KCH5PG3UYa7f6I7nN72CSgNJUlEyS
DQHFWFAFtFJEDvlX7pB+mJrSL0e3EDgJs3e7i0d47AwAqM81epkzj/Z0hrwf9hSOoMURte1ND3ps
ZwEyauEJphk6HOAQO+5kOyDOHXS2SPk1npf8GB1bvzcp+rbOMlV7d6n1E8MGt5k/CYEr8ao37Ivn
z5V+9+TRKBDklr0g7MNAUI7pelMMwkybPpM/6xmUtfVL4kXEhckEJlInfRSb1RPfZ4G9hUVWajDA
SkYGfInm9wFFxUJpLOxs5tYLnJ82OK9WocB5pAtCMoYaIWO7Ybd/EFB4IFr7ppj1EzvZIrQtKIng
ASAGyx8qVJIlcMR4OKeWaq1B2O46C9atQ+hujAEhUOWrvj4+yQ5LGhyKWDASUftwL/11VZpFSQZT
Q5zbXH1fqPYARrtzmUmY5IaqpvHbpvCyMPoRoxIWnXRMB+xqlUmI4GeQHc8hEwTDu4eOxRr3ulZX
2pH/zbvQXcqfIPTStx60qEB0Zb0Lj2uWrHEuXTjnqXxZ2/kMF44N3GaT2wkqnkaENmHSki0pIaBj
tHz/gTDcNIIELdqcjh2EKwOGxp+i50dwLKxI08O1y913R4kmk5WAUI8Sw+KN5gl0nSfX+Rnb+c63
XDE7Nd48W1NSM0TUGPHmXpsjuhu443o+wIQPbTKrAEQKIeMA0hI0y0qVu2SiCmInJzkIquzrdph2
fcnSkDsEVctmj1fKUyGaOC8689lcFAUxkYBpS/KS9558xjCjKPjQXuRwIkCkefpSY0CYL/vLGcww
Lxj32Pc1sknBlbLLW/DWrDyM5aRW94Ox0U4/PPpTEjedqfyB7x1+SPdWuMMLJH0T3wMXA3O2tLZr
LdQ1x6bJbvGMPRoGGeaKHd/NiDWy+qudaPKgv2iB+f2BGvaZmAzs+QTlTLbWFVgjC0FO/iBCfm8K
/5s2u3GcHLcm5pibA8ZxsE5dk5VwbYg4BwJsA6ib9LuoHboOgFEsalsfZo1M7W36nH55cv8v6wYW
5pFDAQTqRYKXXoaNXi8vZ1Fuv8HhYlGN11g3fxPVfq+YnR3r/UjHcCbdNlfA6klse8LaVxsNYJQG
qPu7ypg77g19rZV+ydA1RGju9MeHUwCEzKlNbQm1cORfkbKY5UySIEuD7ZmAtVmYzj8PAZnPIGot
+P439NpFTZRgvJ16WPnxrDEOomg2yfOsgTlAVjSI0MCeuYiqxI4iqVmPC/vligSRy0OTEEMsruFV
7mtGoaWa/pIqKeTyM+LeMGRk2OOKlOiPO0vVYZ5yAe5mu2a31lfCQZNROHJQ2YYvpOvVqE9BZb/a
MoPhAKUoUcDPjJE9NP8ySNIJrEKAa+nbGWUkyevtcwbOZI/MPIW1/TGrawEggRZ4nZaMc60BtHQN
cfVtc7bHaxCTvi+HZO1WeiATsO57VE8j3J6MhA8sUwTAig4fGRQTOtzr0KkMu2vn3/EnvxTuRSQA
B8bA2qVrwsPPGq1JhlInY6mPmO6uWofS/PrZQEmMsEAvUgDYWZb9wra2wihCp12Fa7Gpuwx82kvh
UqF3dZmD032BzF6dMRd0XiAs7GcKbCSHTRt7N3gUdfAswDpiik1+KXFN+F98qm5cYtoZ4M400uPk
vDN9u4UEwplhV+lB+n7D5+Wve4lm+8Pq6EbktX81rz6CXSSu+3wcY0kMfITVP79ckQuJl7smDcKb
Ff3p7f62OqSPSjieMb8nc0X62ueJFRsLohxYwWlBQXc7VSJR3G1htDatre7JZMUvvmpg1Fwzpesr
0JGAVp0VLK28HOUvJO719quivsBu6L4WAn597JROxfEGjt5WOculAFxH8v1bs9+c9G9DLFVK/Ob8
HOX0QHfrOCtyB/hfClfYC/QpmmrMXHhyIRItmJGMjfGFD8OvfgGKAqCEeCq96td9taYtM5OMa8ZQ
Y0ORn8OB1qr0rxiVPXry8v8RUVytKi2pKD5HbOPvQzFTlvaPovdEg3x2GcSvM1fvHiLm782T+roY
8fzrC7m4g2tVvvbE21K2SYz9LZk3iW7ZqEIXRmulGFRKVJ0Bq2OIMj4D/9XedsJwX+m88LenpUQP
IweiaX1icvS7LO/7RCeVtaHwN3fMSyoCM4afWyx4yH2F9SgyF0hXlm8NeL6tYULCqsrLmnXxy7gy
3btAam3BYiy8kJlXhARj/Rcajo22Jt5fgeA+qyI63DkW6w+f/sXAKu1hF58sa7GV2Z9mp3w6e9xL
H0RA25WaSEwZLnqHviG02Y69VGHH7selL0sLT5SvOJzTUjbbxjWqrXGXnA5HzSY9CPIna2RrRxv6
sXyOFyR516wGGWAS9qW2bgGPH85OuXyvGzn3YSfnphi+SD7u1J/6qwqriU08vZo9FssijsWG69gj
NTzYGBCHvQA6sckuMA8g2bMEmpF9htZ+rc5DwTZwwlRnZ4lAh23H+XHbZti9A9YQq4q7Il7HBo84
MtKECMcEqgsSLwunqTSj6Em/ab55G4TBke8x0qZWPFdXo3RjOtjLyLm1raAHVqw+/YfDoGb/4w1n
NhKb3LzFA/WHnPLVjHvV4FvKsa8rNCURREIKn8D049Jg/bFIo8pLjl8a3BAmRZ1xE9R7B6YIKOl0
qLaabref1YW/RnNRHDMVO+MqvVWtSkbvravm6X6bTpqipUO0/TE6fxXEtc+gpCsU3RmwhIeNeBJc
VFcg9TwyDoO8ipyVv2gCfU67zsusVLPS20Z7l6AEzAWKU8AuOtxvpIbomnA7YSyZEfid3WGSFOW6
5ItoR48XBSHBL2scF+oUVBCS6rYsOAyCBg/mCL7gpqsla/CNXFxCasIAGEvV6UJ/U2+mLJqJjYsK
6L/VWWGtG60hYD5Jr2qfbZCt4NRZpYJ8grdD1oO4g+DK5BNYm8d4qdYuTUeBQVnvTkrpd4rXbKyz
p1W6/sC/WwO1FxVtwQ7w70eLtGI2mWbN1OfpU87CcwCsBRryTCK1IYabq4MpyYcpP5OK5KgygJyl
k3jD5kWDkiGe5btqQjj91Uun2m/1EIMSMCAf1um6VCN6O+myHKEBRKz2TdeKuSzn5lJgIBFNT6AM
R/GMK35zG5p4ylK5/saPYK0yDqbR/9TZr9tzE56prOdB1BfxM1ekhFxPCFj/6aqpaM+KN9sh1oz5
HWFdKWChAWG7W5zCkBuPwl9VA+1ajwPfcG1WFtmIdkvESp1uf4fmHkyPDMk4mCOYT6w0gIjXZOV0
1kp/W6T/G/lkPW66y+UhUN40lHMP475RiAk5LWMTwPY1RjXKp6QaSpzsxMYen6rCa5d2A/+6x/me
WrbOsXRPyNbWESdAVHpKG8tWo32b1RsJsfKwj+ztgOad6tMZSRq42sLQubT7wYhiyjF2xNpGKARi
NtUWYp29lVFBHYmDB+ZEgSvDzFbu0LP/9vWmyAmyVfM587SrPlSDa6ti2WklqufsW2zcAb2S/VmE
RM8v+UtwYp/CizmGgGiEeEhCur/aiMT+vvwJOnU8BCCdigYh2M3SnopFxLzvZjx/fhsxL1HlYaTc
XfELh0pQzq+ydPvcwW5SivrHaLviSXzkDP2ILi6v9L4uxAx+eDsKBJu5VQH8O5mYVb2PPZpzNY6Z
U12rLcqE9ikljrKIm4EbaylXv9absxsDwEfRG0omnIoDEI245BxjKo/u2I+0kCKkNYkb0CrsK1hy
H+/EcOga+COuOZBiuLds20yM+jNJzKUdwp3q5QYAD/Kk0oO0NPqUFqZgCxbwX0D6cUmuPCbSSODa
MG1H655tmkLr1iAIH46ok5gXEYwWjU4l6eSzLJZD0+AYdLjIO4JLVQ+D2+/ZD2f1zQEW6xiVOOt/
kiVT+VzmPQbqdYbW4yVqFUEeM9BN3NIqyJZ2hsAC6Em4gPaf3WCWyAPXGyfMlg5mFTyDkqzsqpR6
WRVIVilmlCSidvmNvL6gRJcic8NvyN7xcQmftybqEkYxZ3t+6/HT9TTD6Oke0yCUG3+2Xq/+FCBb
4TpUicZX3Q5mF3brSt67WV0e5vRLfp+pB1aPO6onON4Z+qpTT+PR7U09nDyNV8T0//T3gZeUV/GA
C2s8i816QJE0FiMIwhE7C3QA75f0uMVFZ71F7DA870LPTiwICCzom48IskoojrNsdhtyTFnWMqVX
XIVnb9jNCvn0yZH5pHH97QSXeIXjZfsQTgLHkd6s6gf0RCkqU9CrAlO0f7zTra85zQ6Q7cCVqzyV
/o+WKjbHK9fK8xtDBzoqfDOKVEQ7LRUzs7uqbQiPRhjjAi9SXQgq4M2FZ+M+xOx1RuRXktazD0Ls
F3uKkfZA11yQuqcb+JXLyY8LBaNgTEXCAEh2gYkB5Qvt/EvrYG10iefEy3HEAqmSGAD50oZ0jIeB
aj8oebXVJ5mc4Vy6KS4s9+ERQkrVwHu7dDnOVowLyrA/7jc3AzczcROXTWhI/6owfg4FO2kuvnnA
npgnN0U3+KlLs75w2CDZnuwpFQEPdwKDtXasD1Www9FEa+4Qon1APuBptuZAiNJEXpkuwG5E6EnL
aDj1LYycygx/AeLb4s1S2khkwIcK1XjVzc1U7KPoZ/kdhuc7UEkn0JDKW3dt6VJk35ied2YyvmYE
o3BFT9LZvEPzMsQfCc+GbEIqtrUr/grrw/9vczoxobgwdjpQPfaTVtlUqXQCaeQ2+Tt3C+9XsWwV
GBww4pplZMLDxxj/+pmiSgd4/hBxphVijyVgWUiklCwXzyVxQLi5NNO0XN69hYbs5U4E1gzFbBBv
cJmKPjRrSL8gXAb2/otFW20REntY0PUy0+394YhvtsDIb8ma8Gu8DWecjyUGUixQt2U7p8bEHzh0
MvCB4ZZtkIOiH+630aqN2uEfYlAyNNYJA1et4hib6mJuz0nwqShHq2IwwzYGWPpb+LsxcaTvKEcm
xYWhEvalwwTWTbXgfpTJ4XLhUFG/iFRKwA234KIJTTUzWVspnYYcH5SCYetGrMGo/8vAcDx2XOad
NjCF3pauJuNbvdv6LKcjnMs6hmpEKm3C2iCqtnpt0LBDXev3mA+CIHISfxGtUHXBYanuZZyvTjii
aKe0PY0duCImfb1beT8/TYc+GnbWEilyGanPtJDDtnh8gD0IJowwrXZ+1YHftCqfvwjU9bCnz+xP
ML2qt8pkuHZK1DKlsp4DxAOHUEXVAE7pu9kde+7L9dn85iex+Ouuv3DpRvfqLnMKTe1eSkSzxSK6
ki7sFoFxbzpURbOd1JPkPxy5qPgZbWYtGVba5dEIFaMkkFGGQPFlEDIS6rCJLh9+10Z8J8S7G3oY
DkyDL7Dw0KuGdvx7b2FhbNyDyf5ExCdi6gY9BdmRiSVgBK/8aXxbGl4uljb2S8TsPiMyP5mRA/ch
6Ttdp2js3foCXYYw0r8eZ9AyAsOVAEeMTvJMb8gt0UonPGgtSx6DDPqb4j4CXhnzsl/vCkqwcFkP
LsXF2CR0x4t0Ncryzr5zmJidcm2H9jq3QGNEFAnpIVtDk+kAlqmKswzggBTV2/rI8VnlWDvADwuw
3GC7Tn8FrR9Batbz10HHh6MWPhVq83vEu1x6aC+uT7wMnUC00eNvKdm/w3aH+jYIy0+6wFKvTIOQ
LUbm1skessyzPRzX7B4Q7lhppNXElRHxpyxiEvgW85tftIgvEMygzFedwM1kfMosTUVz1NU5a/C9
l7rSA7A1iztq5ocntCvFHO3KkjRPFVGLsCL3uRS7Ze9iYpaqkh9lSuQY40H+LEFE4IdNefin1L7f
N/JCGllSTmSAqADeYbvjJTEuDvfMvaop9RJvftXl3+1Hr8Q8ps2/33O4UbxuOHfg9AZQV6jCREYD
PJ42d8iu2Vr1st1yMvsHEka1Oop4uue64U9J7JPO9Fsc6yRPU2uPtn16ZrsVwUwf62+Z3xMy9M9O
GAtTiAzbC+x3D9kCE0We6vEnclIjRGxxlkaxjYct5jrVXy5PLVB4sSArj+0RU1n27QGFlt4Gt0fM
qztRTEoGAUOxISCzeWGJe9wQj5VxkAO0MbIgjcAWQT6j9zdITTe3jYgonY4JslIc65Otff7NBczM
F/fhXuDLPpOoFGwXvpBWmZwPNh3vR1yK+/rttFq1N6iWhRPmRLakoykOGbVESJfEeW5C+MoSpErY
hIkMexP3cYOMwNnAdY7gVgOzqRaJye27xL0avkwlgN9dFP8un7WANxAkxsK4/5b+0Eu3NTPU9a9d
KFfyafd9/aARbKQcpgbgHcAF6F0vrhL9N4BRGiMIArEU9LAO+JefCxd+COafzzkV9wB6w9weQuC/
/brDnjrPtG8iZ6J85gRM82GKxATtkErDimPdPt2rwgI85dzB6I83XdgF0p3onjoeDqH+eFKAEPlw
8eFaQ8/GwARCghloiglGjvfVKtgJ9aoiZqFt5AYmZqaF+PIIa58BvFA4nTb3jCRo0YLVXzx9A2bu
gMUYIa6N3Qj6dHqD06sT/IqTR70JdNDlpQivte7f49DTkgsucuwrVZUWJOt6Qnvw26WrjPwry7ur
OU0m7CujiyxlMuysXRBQVr3Czr3XFGS/MCU/D6IAwo1+gUa5wD89+rp1SzCt31MAOnljzLe1oa1u
c7CKiBhcXQCzcGjMrKl1Huj5JZ2eP3aNB1rflZ45sKKK37vC3U6cmXyeM3geyqag1A7D2mWikFJy
egSbPjFmgpTdk1de5aljppP4I2mXwQj2zUIhpUhJHGwJBQKfFTAaWNAUO+BEqFyGsjQgyX9/YVOy
qo/2C6kLSfmOnzA4vnwK8djxYgRybVc/4o/dt789TIx6L89+SoBwPz7aB3xgcASAClm/Z+akBqhO
KJuTiTyjm5/cr0EZsRWaY4ibSic9Tk3Dw1dRWfix9JBAic3eULMFc2/zVw2auOk5ncjZ6rAFFmfx
jY0vlFaGxWCwDjpbhoWNNFKXs3nVe1c+dtgIlPNlP3FevFc2o5bmsNpXWYsSJZx4wryay+hUR3h9
b866A8fTct+LmEjHpb1/9tlhXyv9FV4y6IoT/6+OzPTX+45R8fT54r4p0qy4A92aMVf69eA8de5N
z/FDulaAPT8mGoMwyp+1+ZBeLqy6yEcrPefr+WqIJqPiOrLHGF9UWHl22QJf7Wh1EJKhG1W3LA0l
806kLX6B4adZ4EKOLG4iCzFihbdQVFaY8qoK+ilZ3AcuWyQ9CDGzRM31hbP95dhP3Fv7bENVn0bR
7/NFH5MT90SNosvv10zN6grodNe4hQaU/ifQcWrNOOZlP9DjAZtPBPbbruKat1hp7AwTAm4SHAFa
jULsIwhhjigG/knJxxv9+iG414jAf3ZsESf7KAMW4ALvz/k1jSG7kCYStAJ/heO5mXMkQnf8a8vz
RwZEjiXj9rWw3E5Ae8fRqlTpsfQINVa4z6STCD6KxQOsUMsmDY0/TCDcnlj1v5NjRMH3i30tk0ew
S4tYjeOOmYOrRGAv+TvMQhBpgmVeInT39RI2YA+8R+4TMPw3Lr5H+AJrUTgX1QKWHT+dSgAnJnGl
D/+gccix1xZ2Xrxz7t4nha1aXCsdNqSOnerwpWm1yT0wCLqLqI6QQHFaoskmGSLNWwSsfFZvU+uk
gEYMP9qI8No9AjYP9KGg+GYbI2/+Fcr5KNqkzHFQ29MtbJ7A1wBm1gzREXErTTYCtBZugRTvVZLE
2m4JhowDenRFo9lS/H6uugLeWfBe80BXpnbEWre7U2QU3ByvrPz2cs/9IzUqdew7myXj4QHbdK0+
Dd14Fayfeaj27e/JayP+4LUg0D/yun1A9eFVofUaVX/lw+9oeXg/Ad7HSqLICG3X5piXYCPVbrZB
qx0l0Te7PUN+R0AabuP8mNclEGF92ZRjoZpZi6KnkEPGjMjqM7q8WqQChE5M7Q4jTeNoTwzA4BZR
RNotjt6pkwEnQOqYk7cD7MYwSKn/S73DwynbzmtXfub3Ni8oBit0UnbPqc/ee5uQDRn7Yx1BRdRZ
wqXgNt7I1zDmo9QK3qEG+vO3vanGGSGYiL0SgL+cZ3pUQTotm7geJ+WYgZOr3hLpzkzDvGchPQAp
JlrN1f8/rbM7XIAPc91RZFdP8cQ19vhdTreSu6QXJKgYYZAm/XLkJLPZD4u1B0poev3pWO6a0N1e
IWwRqymJgNMOOqENMXxiUMhTeZjrIAPcx4H/5a5Y3a6FrvgzFgooBH2lSTWOXpQ5XhuORPPuD2C/
BvYVcR4zIkC2RruLfEoaKTLRZeVH0qOTKsp3rqRfXiFtaQilMSVGk0FD8zv2u7ap2N2D8+pGxwcg
hlN5d1cMwuAfXsIe9jUFHsxUyS25gE1cDqTMO7+uu975aZATEeTKjfLJUEoGgS9UoOYwJWT5uznZ
Fj47I01+jr+tgVHlPxJfHL5HrktdPCfV6xDNQ1fXYIUaEJOu+OQoaSjn66z6vePw4LaN1e03Y4Zt
GNrjQ+0rvtJhh6/gu/nX2MW4Xj09uSKYrdF/aEoOyN1QUvO7+U/M8BTtnJAEtuGPTKB+68hyq1Sp
hFDfX3LA4zuaRoebob1eQyymudPGOsMoruwmJa2juNDn7nWypNI3QY3CqRls/kXtFw6nPh/kdU3/
AHJTlt6AlU0MVYE9oEUDKeWpcHDHWRSyuwsngpilVCwp+21Zc0aFu95eoL/0kltrt66DvZeFP6pp
Bbwi+Ujv+qSUf1IHg4VUY9ZL+/1Sqg8olNy+p7jKKEwzl25Zwk5YdRfbo8QaRB84NcnTKFy0I4LE
YXT3v2+b+sCFif+arcVLhmIvwOun6cPl4E8zYmWAEnEtNUtmwKwn+HoxeiEkUIZcFHvznZi/0GLi
df1En9ixBITEU8pbAKrFxy03nqjp2v/n32yPMSvpQm6Vobt+f2u2TSsC0j0HLAkjj1DePavHtCZL
GDQvpxY0hwZ1Seulg9COWOgsMT5JWQl6w5kxZXYP2lGsZ17o5PZZwPdS0xNwLIQw/3PsIY3yrHbr
kpHppzcClopAvnoWbjyRJGRLtyeL1q0L188o3LXHhWxKUnP45LwW3VCvymcSvhs6muUk7hfo9YOn
Az2okOcaOWVTiznG9T6DI0p7Y4pOrXkNgYR+5NyPfbMsHl1WuRZ0dHxkjx5F0Oq4l/5/rX9HRfhE
HjcbXd0eE0FA8hFCC1sU+xdcaxoS4a1+zUdDw36YkTOR3zWhwbFqGw+aHC/cbsbWLJToVyUua/Id
ocYnZaJM9kp7XgKul7ZczenkRLgD/VpIhGNS8dAkJ7m/5qlN1a2Td/YAZnNNAxZ4PeEB2AIWSKbu
r/4J0ySLx/Yy8SCaTX5ml6LIIWVcn6wpGqiMe3NyXlDmbYi9qknYHeuLTqzWBXZydU56XNPBc6Ij
7g+ARb0m5geU8c0c1CAplgGQD5YTELdoq2DpzFOZLNbHXgQ/xogE3AO4SYtbRwRiD4P+ADGbt+Wh
uEplZplutSugUXetywV0D36uUrwjnDk3l6xvIz5Ie3B5g0poLYl8ySKOTz3/8CGsLYFE8ZM5RsO1
9qZaDiBwuEynXOlSaLo/RsjNIl/Z3BEzSXTclYRGl08uZdCgK1SiHzJ2fOoyo9p3YreXYOgPkPW8
BPezIgfjv3mRO6biplN8rR/DB8KdChLWIMpTTLSfRUtVxkRmCp7RbxZ7vLXdAtFCue60cU0lyk+X
M29VTE6mCCqT6eS/UhxLfMWCOpAqaCXaIgExK5LsVYVVDyvHUcSzl9e4+RTZXJmgs9NPzWIESmj3
t9AxOBIJSKKrgwcxPOV4UBI/gYSLZ9R9MAwN3JWtT4dbiSr6f//dHyijArddKJkuivMDCZ52irsA
L9zyhh6ThfaFaOVY+ETob9T7uW4c28KUF4TZ+k1jDGD/NLW1oQImx2TscsrWXti7D6AalQEPR+Bx
DpgDlBanYL2aN4S9eM7/QRtimY4tbxE1+ZmyPJT7qElv9dTW7K1IgP452F3w5ssL9nBRVvwFyX1F
lEAolu/wCdp5K3r4qhdf/xAYE5f3dBsCM0fvI7eyRWPNPOs3HYN1wYSB7s2j1d6kDn89MgLS6NbU
2BAxL5tDX512mvnEo8HaT2MVUS89stoz/7XElwOgZw9BMREn8sMO/urR5rOhlMcl9EBFq9HxA5d7
J6b2P+HvRBJSSl9yYo44qKcrG1i0dLJi4JfVzPxE+G6SvBb0vVhio9uO4Sia0G4V2md1huxtWM7Z
LRojRWjpr610xmcCOXi9M1jFtU4WUoYZz6N5HYrtEsvqgLnJqtwXyRVy6+HP5QqWG65w1xZgRHJa
pT67li+SqbkrPoSl64laEoR037quobdyAvlfrcshQZnnHbrF9ufdEI6mJyj3G/S/Ng0Ej3MXifdf
cBnSVTegmZP8S0XvKhssuzKEFsRE0GFlUVcSjqVlLPG0O7anbBICWuDN2/vnfKlMGfTwgAn5gJUr
uSgThDtbs5b2EwkX6SFG8A85zMXHZ1h2OIuuMJmC+HR8wa46TaQ641mTgEwNobZkvnMc2fOe7Y4h
y0xao3lTXdNdwnjAeXakhu6yw5MaIk6dG9hlJQmADMD96SbOZodgDSTTrxyTlhjKgjUje6v3TUoa
Xc+FIWVRq7gU7UsqvzfIdhSPXlX058abH5dDDBGFReXSQYwfGS0KfPS5XeLyA+wOT8y/LZwi2P8j
HCqqoQxPvi21XhjUqs+kRyuMpYgyaXt90TNxeqI0MRDFnJEBp/aVSIznU04Md6bB4gcy6nTWM/zV
GQPnqFHcsmynu8T6Pw9yrRC6MsY+JLp/hfH/Jd3hgH/igDd+VctemJGbb9AJpgfcjr/xfnGXzHsC
yfSQ/mylpItop82d8DxmrRs5GzA5jT4P0wDGxckXE/DVsRDtzh7BgKYFP2gXW+iA1wrGcgJe+Uqd
i7sBWl18l1DJ0q+SyhPbCRnwdZrHoNe6MCSfdQVoLml72kkFvjD9u1ENQ9jCYqzGY/xeDTkzhL5g
ZivBmniGirCbOuGRoEswlfodbIDwzRKvzFG/mKBqIfqe85bekKquJPSAMTJp7xCFScJcTZ04CFBf
bHRbwpEAU8EDlGXgGQQu7Uyl+XbyFnmXhmd4dLxwapDI8ZKNSdy23kF95huCx/666GvrSKYM1v7c
UIdK2/HIxIQqYy/IkSgW4eNV3xTPCVbNgV5qf6+nLxorNs+kB8FO2dw4ptTyK5MfgfqgII7KZSJa
Pyyb5LK8P2IsXIixpmK11u5dmspBfbx22ox+tnQlr2Sj5nbkkcnwURwqHgtSIP4z2XiDchLMC/qm
YuCzlAANfy2TBIScppccVXsLtDs6qxhOhl8GNKmMGDST5M4Zi3kUBxz0nmDOz8GpkdCyDXlGbA1S
wtB+9mLrce8WrLY+Wv6wMIS9eefFmxf337kiLV/YAQ70oGBeyxRiDg+nuLk6L54bkqufVgqwOW/1
4VUvlGsQHSZzR+J3vf8GaRFgpKMQaquaePqGkBKZbSxaBvHAyd4qbHlyORkWHI5ftBjXjDbJ4doH
IWJNG+hZP4KN/fJlnucgsAqgzqEyU6ZhMnw5UrbXNm6ohfoR1kLMSSrxv/OPyyZOtWiaieCUQDmL
9JCJYHtG3k+xgPw5lvOuN3krKpXj3H0mEjuVmgxDbKa+2LnpWAcNq/tjV9kJhm0PGdr2TcKBxgef
bC8wsGweejnGjmoFWawq9VMLesBCCwj26jBA75mP1Eb7E6U5K4/G6iGQ82gadMk8MZt/yi7faBHT
nHmiXuttX3c2NR/6nveOzqB8WSE6IbhmrDawAWucXv95RL0Tdrmeu4Z7RUkwjuxfZdzlos2Y823U
GvN3bkNrhDta2IfRqj5DckcSGhRBBzvB/NLCWjYQsXSgXt3CVFPb0r6slye3ihR1XT8O7QA5m9aS
WesTbHs1BlCfsZtGgvcRmcGH9isKVB44fleq1W/xU7xjF3vSaZ8lCsmnSNFl2aQmbFxGV5uhgdIu
Il05+LOMVk6rF0X494QQjEwZI+L5b9Zpohr1nOj3dPmFFZzbU9jzbE3hD++rAS7Qsj0dqAPT8cpV
5P/DdbhGGrmH4OdaF5fe2VGlCBKhjN1PaLP6ZpdcEkHV62NUuJp9Suwdy3w26R9l3sZf2DzPikwI
d1lmdKmSdYShIx4q4rhCceMkanXa1Z642lq2nqdrP+IpVmXuEpPbQnfO6+xxhumPQcAn61XyG+Pz
fHSdNE6DXxb7vEhDNqIiQxsjnz9xjK9udog7mbjwfGj8dHIKVLBq3Jqga0E5TeoUM5wbnrsMfqZH
lt5JZrFvUa2ThBv20u6M6q/DLjxGae+CQUYND28EwamPhlofF+s9FW7p6cZ7VvGOKLa2GaYeYqQr
9uQmxkkzvcHi66fMERqJs7SD4hw309g+z+bA//7xGprbl8B46yngW5/RUP4rKznDWUDed8rOQu1p
ITRn5whmS5zmE9Vu0UIWU/+8qnAoxxQmhWqJBSIaud4HZJjo1oRt3Ix8SxzznzMtsJ49Dk0ByVa6
KUVEPxDqETAQPat5BV9OQXmL+Px3F1xu1lkq17hP8hNzCwQtmNSdJvyYGv0N5CyOn42FGSqUAQQo
pygJUKe5NPMop3XPGnNREizB/F5+C3kgrrOyHjXzSRgnLdXbjC64ThjNuwRVD5YB0zVHGXAfOzW7
/YBC/eCajqiBPN0RaDU6APp5Wc6rsOnjnEkIXJsbtvQPNqw5NobkyXNUuADRhaqSvizDCW+2pmpa
1xI10AM2JyAWkpTfKbTdAVO/WdOCYHqnM579A4gmNXv2PS2qQMjX7yuRbmSC6FBrzNiBrz/Kt5XZ
NXLfL8NbKAWlIirMrL+Bkk0DmHjuPdUOffJaN7Z2w8S9ibHmM0NIOefasv1UTjX/QzUw7km2LT5X
42s1jKJEiyBv5Szdyewi0PA81vxX4uhos1axhi9X6XyVX4Jj269W0ZSDFEVXjCxMy8CRAAZbFcdF
jPBfoPFzZteQblrPl6JYAmgPrjOCaQJC/K2waN3hKLQr8eR8Fn9tYNVIuqHblonAtluaU0ob87Fv
uleQG3eIizlJBzM9nIzeAUUD9L231D/+j384MaMlOZEOmwalweFPp5913IiIB2gZ12tUyDwrAwcr
NiYwhHyypFxXG23yxSLZYMCEDxDbRjn6ryLGf46f71OwqvWI3nZuX6DSdPoduKoHEAVQ8fFNUzho
fJGZB95Nnc72qYJV5dTOfTwWusXRcE9uzCB1AE0cvBTbY7UJCNCrxHJnyN4nkn7hn+FLXBP3jEDS
bR/31CUMAbUPX0qibFzPAVFgNYRTRA3/ASYUz2Ug4cghu+njTA5w/SEftIbCJVMKt2jlBb7KLDOq
wytoBgkPccEo600hectGHP8zv/jF6UgGS6iA5XC1mcSway5czVaSZkDAdfQt6citCQR9Jtnu7DM0
PXVm+1kihiFZatlLkUY0lSxVG8rweWtel6Qrhow032QoPo0kKHfXgH4yT+8+OOykl9btP3uzYve3
i/tdunw8dLq3XHczd3g70yTNOzfpm2rTBvM4r1Wi9jNnQeELkano8Ka/+ciRgMZZot+u8tM4Tjme
SoY7HGC1/wAGhBhWCgtqIoNOr65kukHJF77LwG/3bc7+MlkG9hnKjG/22iWTUVG+Z9bxfwLUrh1E
IpVwVpxLHUVv21Ynfo3njM6DXKysnJP6hqJu4Dl5XiloybGRz01Evl8HVrTElLERdcnGHsOaLrvv
3TzfuMYDYHqA6hnFsUpafvqcWcjl97c7iWtc4zTxiasoY078imv38b+ktppw6mdir5wYLS0Azypu
PE3HC3hkiV0pf6jlb/vnR/2oBH3yvxIsjCHKb/1gRBemYhywBm/e7CQmwfZy8ResF5QEH+dsFu5u
G94wmjC3JvJ3+XKLl7a3WODTi97T5OkDB0fIkp1OLroaPIRUpp2vls8bChVURSf1anLpyX9yy7vr
fanhTB3jl9OZra026V0cpVVWlrJzc5MTzWwP6m2lexbnh6j1Lni26DTMW8ndyvq+TpQQXdsO5pTe
hXsXJvqmW2lze8cWxFBceqngkMI/ueS4+ndExr5uwg29PsN6czg/2VFPC0chr/m0FhJo73iE/Ujo
LLcnDXFo50hnvqvGZ41/uwAOByV9AGFwAZjlG4ncgHlDZS7hkfc0yEegDxb/xw8GXbnXFVEoRwi5
K1o7J3wWUShdpTRbwIIcYIzvWH/A+PxsbfPkMmsZk9fXZrRhDJRdxVAgs/Hw8DTZyZwu+L4iaX2u
OvuIwjgN0MzQebEGxZoZB8pH2hpl36h2la/FS02AgMuVXdbpRH3EFLKg5twuRl4SwcdTg8xknprM
OXSPhdcpYrkRGa+I0o32dIs9arbSAaBHAorqDUX6t7OgUZNDCYmoqD2sgKJ0YJp76ITGeMGWKnWp
aA5tRLB6746+8/e/TXloegRri9s3LwmbQwpEpWdr5oNxyETCfU6aEgYlQuUg9fpIj/VZZMuxOziJ
1Kp2GHzcVyTdKduRoyIISw3lvdAMaLExmMSbFaqDeOqWyoJFHT8D/Ro1Ua8MlA7lg3qwjjBmIrEZ
kVBx2f8wQHGOB2fh26BQ4FL706UnpbZ0KBhOaLDTCB8fmSGyyFhlEhIALOPU4rN31SMbd0TNNVwa
VQ/rv9/NmpzkeMlUDdPrqglSFoZVRDQpIGsvhBFXiwcQAv8a5YVuR2fd6gEJN6hULO4f72cYAl9k
DiyWHLXpwUyRzMtMpwC8Bb4fLCWMc05Dj5bcTY8WAYCq8jixwBnRwa4lmmnj8+3nkIvJ4NMDsPxm
Y/YtIffEsgvnb1CfVsfZngmQGFDisuRa97BaMqKscroY85KCTdJvIhd4Fsnr5zjdc+MNIagMuHUk
DDojdxUOVZJmq6wAN7aTT+z5AYPEPo1XbNszPYdOiBuWIyOhXsjH1B8NPIgTrMzmH0amNQIik3Vr
PgZIypqIty1U0Jq2bQ9EfxQGrSVGfT1tLL/9RAAXotTDK+Lfqn75Zdi9U7IAvgknDypUdxwQKOrL
MSM9yiOc0bpMgt1Ekp+rtgh5NSm0xKwlEKxhac56+D39qhmI4nNCue8Q63V4Acww4N+WKhpwGndR
8btvdyxigQVQx7MrNeliK581tTgGjta3BdOLNXzvdop/LB8cPX28Plxj3wW8PaYX9QRtuCfopV2P
IJFQ+++XVzgk19/G1fRYsVt6EOEQnhYk61kHACXKO+XrYDMO0QgOeEHUWyA01kCVBGZOZxucMWJa
0C5pZ/hg5Cn6EaBZVVB1Adym+r5Vx+OplCHp4KBGLItrNrudAslaLKwfV6kxen84gD5Pe8oC1st/
a5jodfdTd7G0pcgGU9YM5Q0TeFfTkkX6QTO3Mh2nffFyrAseQ/rzgOAKqzGsbJFPdvZH5/YGi1Kd
O1zKD1MfCyeDTDkKijmKg3/gcng+0jutPAV/bfGHI2RganjMSvbHiq0KZ4SK2/K5Ipr0KSbo3fLv
y09Xi3pjq1nQ6E4cL5z8Coq0yQyArh7UMNzbVrVBJrTGOwB8belVlg2tBJNgljF/1zqlnOnEMRig
VBxxveXWDP4oYsuZ2melM0QesaigwTYOgUxvtFVCrWU9ZBek4841u98wwc1vTqIM6slHB0qbOAHo
KICEYwYqQJ+ks3viPTKnmyQSZEVrSGYexOgK+kmCwSCv9k4LEYvR6KxDLg4yOXzzwANm/HgZcDr/
AYGtjpvvlCAwmAgi6dFgMCF14m09NMpsAEZOwSjhvsct3uwLfRHS+xp8rMwqVLIDD8gfmBwCWgVM
1m5EBzYb2lXm2PEUl+9A5Ivgsws1enVkf/dOhVvwfs5B6oFu8Fyu/v36l7AQ0gKef1PK5NLkdZn8
4xEhrpSeJPOFuXxTZdYt1hdxUm5HEb15vi079oYBKgmcqgnHyz+4MaAlXGSbeYdpkBZYrq1IVCHT
/8Nk+NYOreacWjkmtEC7b7HNevd8OA1zZH9iV0nfxhfbEtotk2mkiyVPIF58vXdKT56osgVpSixU
+tWC+DZhfVtHDcMK9sgmSrsOLF4GgA4u1UX4RWhu/EedyWblnbWfAOCsy2FjyRSCDfDofD3Xq/zr
H88g0A4+ttYxUuAp2I1sR8ay2qhuVcUgbvGe4ORl+688JC3fNDxw7tEQaifPkGdS3FeZGw31IDTL
ChLaBEOnAVqsi86zYCuViBfAOxKWZxKnkAdxdfTotjvKUqWrh6LR8gI4cUB+D6q4F67C+ni0G/po
kvhBQFJ3s7zg3yZmONw7cMg0jcIuIGMBjbKYUuihZ/kYATsxFx3wzIAbuCy7wl55LkP9sJhO4y9e
GmAyKPAxl72VnEVh+O5UJOKwVOuHI43jUuUwXAmMU+Kims4/Gap+6seRt1KtXaSad69EKPn3H1ID
pnbwOZACAoHaLeN2TMOpghtJIbCFZNcxxz/cqSkZMWg3q60Po3cDsmHHQXADT6TdUEn4FEWVNk9y
yNoUH2CHNuGP4DMUnodwPXAtB3NWPETn11T/T0N14tWEii5AO1CHJa8qI4jUwdsc45ANmo4o3vKu
7GH1bPoPswq72hbRKk87m7qXhujzfIHevoq9pI4WBD1Yv6poWfJ0xvZLMOqG5Pw3sFmzwG42c4vz
VQzP3JoKSTWtZAUK+2sxMiPA69Wp++KEgddq+g4CQ/tKTkhtAMxrwd9Tgh4zdT3edYR84skYGina
bLtk6vbcYLvZgDlRKn/hLNLUZwaB5XKb3RAkHWoE7HAJu+P0GH41dKeZ/UE47ggVJaCpO2/62j4U
/PIa/3WLG6ng/cqoPNr0v8MQXAmwwgLjc/Pvjv975FZrcYldJpXnax1+j4P2LuxKRuqqxV5W3Cvg
oqwpXO4xOFCrS0H+eJ9Q6K+hP8aaVnFStbU329w0hgvAyAlINRONWOhbw6yA6u7rUaIXu0THKRA6
GS7EjEGlJXlr09QBYwGtfaw7Hfz8PZWB2JBtOd1NfeEOddRrilLPea93IHYkkS83pgvXN5dvZHld
hYeQUVZUkMN1jqjp8zZY6Qx6XHw/eevM1RwgVNlfOTCv03b3u4tobzgV6l3wI8FfK/ztwn7urf7d
mVo3o0iHTSIdnexdk4lItC+tAgRXgaId15T9bpznsiAs+eg5ZTV7XWq7sn9tISTjJg61SRXKzqXu
G/nF2uzOuLTytUNIzxyciaEeVpNZdRmEqxQKDbK7kV6J4wr2nn1tCIk7G3PFazqLG/YLEiJjaP3l
LnhdJzqkl5K4zBKmT1hDUqk0i0R4spAuWNO76V2v2Y8WaFJJubrxe5uGUO2KSnmdeM9g23g2HM4c
E3ZS1VLnwLsiH5aaC/g6uPidIASU/2KYDcIoj6XwX6bCLH/SfHU/ZtFYza16owfsPQAa3iW1eWtD
4HiGJPjZ/lLdQPrj9RveEj0SmB+WDiXhS+kfhbD3ZaZLFfbaeBThXaSuX7Zf2CiglEMsuYM5MebO
gWmfY/M34/SqMIywwbMFNPBllG2mGxrO1cvizwqhdiwp2mbS+q8CcjZu4PpFYK6Rjns39RQGg9bh
hIt01hV97Rlh+iI5MyZeau/i9jPrbyInQ6kgsQDEwY4HxKOB2eN+z+caHPnEY4CbezU+IlAAkI3Q
fbvQB3mOzSHGoUZPSOF4f2bjxPpx602d4Hj53ur1WWZ/QcLCnuLTCER7TMYuICGUFwiI9hXNqedw
TTJXk8PL9Ip2Xp+9OggLOnxeVkN7jkdQfIa6Lt5suSORo8W0Ur0bBTJHYBNzvBvCYBJc5vugjzJW
e358wX3z1uf+WuGpMC1VDRfKvzViXEZd0xB+HY5PpA9tmdSVwGlc7jVr65UEfQZzCQ6wp3+2zUwM
AwEA2yNPh04ddd8gingI1ZePREDZNKO/H3gouVinkKMLW6y9NvDLsMiXWw1a9DKIZu3n4HAfU4Xd
LzkRXgNHA3RCuXCSe6jqNYVJfRMuM7zeSCy0I6oui3jmHG1bi4O2EjBvuoaa9Ga9JxVJKjfRvUWm
2LGDfV1srgWpX18i4Q1GQbDc0VCHxRG8oPl2TmPadpubzwcSoYhKDMlmlvBdfPY58gZ0RUlY02en
kUJ1qVG7sZ5pYRDlKnRSGV5EbBAGkJ17TutWRjrJr/6qApBGh72NXJI9pK/dgN0r0E3dDGXcqhC8
IcnsI6I7f0JXn+S/Bj2dGg84388E4Nw9NEEEA69ioYTSbrh9nhipEGsWlHx7uwDlPuaRrAnOx43Q
4VYqoNsLeNz8asU8oVf+vK9hQL8tniBOb4MDD7QS93wNYtlNZ9ZIDhQmWkwK/nTRo+7Nwdg03CKm
QOEi5JRGg28zURg2EdStZUqYybDSIDWKZlY2EWKQY5RPpFudJxQFFca0rW5VRmfrt//ve+scA/x4
A5LoHpRso5HCeEEyCpG6C5MLliuzAB1l6jXkTNIDZJaZQ0PLhm7AR7jZdOpHosFXnzVRHFwS/7l7
E0tjuoZYVXccdFIkK99VGNn7MnSv5/skbPKxKOK6IV+Z2bm3LFL7juKj3hHl0Ehv8BQ0XU1i12ZR
sGGnAgRlNqvL2Yq1aQsLbX9wzKIpqbX3jc2or2QaxCeeHUXxb9mP6EBSTfrgSTHiFT8HPanQOVWb
IjOZF8TEQyj4AqpxFF9cRy7I+AfA0mjlLu6bb2OViJxWWMy7opLmTdJEJ+4qoh9tAU4t/CvUDfUA
F+an9kbzzbVpTmWiK5GzbaZYF+HGVdhoyjWO1jyJ+sSHdlyVyWHnrCzvCJkSQbX9Xkv8B87wlL6T
u+F0Qr+aeCeGkF2SufqwN52AOcM+PlSVF05L+9+GjuBukG5OskX/1iykW8RIrPPIeXyRrYeus6sz
NwEFqjS/bhfc7Ra+avLepMXEfnaqJv9S6ZRa6XGc5lo8VA2eJYl5ZvlpCnlbsNh2LcFxsOtxy7/D
5rjGpuBXm1oKCeF6ydRrRlj0Tyus05NovusZSjymju2BIag1WkJ0L7+JhfpiTghwTmM3F9qnG74B
hZeCRBgS+rjjSWaxyQaxpu4wZr0bdlegKcJsvuR/eqvJLTaCW8nPHxDLmMBqnnBE92KxkGZwMVUm
t3iZUmWvBIw/1+ilS4mBNGXW3rEijcAqziz4Q2QnMFd0AaQ+hq9PriTYwPoHOJ1KJTePL0KkP2uU
ruKnHM0vU98a5u8plXqP3XZRAhCLWAokFZvWTMG7GYS/4Z6fWaTIpNcaoY3ZroVwJbtTzASCqaCU
NSvedwPrVqacoQePMpvpoAqOiKq5/+BmRFntUJUn0pQeKQntBW5Loeg2JxhMe8pdrtZRS4H0CZNO
qh8jqZNo9boiXBcpmHf8Ui73iIxRENdL8zQ4o3JK/SoGGBm4Rr0D/cc+8LBassX0bE6TNNEQzuRt
wYV+wEzVAG+qg7KGxaZKex9y/jY1EWp0Brc3M7wUNymf8lpY5YHAsHsCqfTuvZMZ2NirndkjjSA+
R3lNSU0MjqqnqnxszgMLdL+7FqOcVaHSI+Zw5wlxu92qBnhkPWwBB4ygOPqUzCT3Uh+OBHcz48zD
IwXZGE9rIs/oGeDoP1FQnMXvp3+iUSAqxXVQGWwVvue4U1aQhvYVdXgEI6QklWBhYsI++HcKXzlh
d9EtV9XNsncZdga86nE0sdUL4TnB2gA2DZ/+aEVP/Jm1nKbtCZbeckDUL2OZ022xeprC5hQ1X8dz
vvx+KuiEy1fIlrLN46iGSuYuu1/hc+PwO8KCtXXax8IZM9VNKjJl8yJCGyVxGCKq5f6PrLTvqtx8
8TznxlEPLw6KKI4b3zJDhsLcW1M2zvu4Fc7NttNGf0nhQZwlNhxMTU6UeYfn6WXgTmvY8DQgKt9q
e673g68eoNjgCYtro/RLN37Ig5cB9MUUPgn2Xc+B/RHEiOdXDi22OdPejCzqGZSuX/1GZCK3VVF0
r4/fEzym6tQNCwy5/wQqpEO1DHzbOpj0D9H5puOF4LPaAA5K4wwvTM4GQQX1E2YKa0AogI0MVqL1
/HHcGWancUS5hka+4agrlm5rVyb1a+NvyZnHlcZy4nm6JukTi1qWGlTuLsNWCLp9vP0+OpAbp8gA
40UOKgQeLNYfMXWQ7hjvbnHzIEBWw7erFrugzvDzYPn7S79szSnKa6lxgVI1/lmKZFloZyfPDmhK
8MoLjHc/VGwG40FxgT5qRpzMxPATJtCTlmBdgkRvnKBLbaE2ZnyGFxAYmzRUKdoSZMCux7KCt7v8
yOWRI37J2pyITgDUY5+gbzfjxxqXOvoMcwXM0huyHTx5iXPgHqg5neiuWdU+4zgOJ6X8GoI1l30/
kmYGGX80HuI6pAawsVESj48qhy2p3GV4/OiVmuEyk/V8D7DvG8WLwWidwkZjZw3yCgv6GBXigmpb
zpBCl/Cv/yinIpOt/HdVelQAU6/0VWf3ZQ/IfuxqeeLp/BAhawWC2f46hF0h/aoB/vDezfQzrqYH
JVkEh5Os30rQSXNuTGS8yzJDCx87TMh+HhDlRBrpN9E4k+8Z79UHvp/XVTs0gAYoqnX3RelGEIdn
brJzfcqbTUxOieqqZ+9SgS1EgVCATxv6dWRlBCQTMy3ke94FdJ5xOsU2gZlLpSZ/1Dbn0tGAr9zQ
KNUu+ia2xYqDBu2Mf90CkU4PZAf5NRGUhoUVpye98CjFFVcNxspLv7RNbgjRVbx2MK0J6WQIFkP4
+Mi50OWVDNNoMeeCf3OUvkGoBnQQHPUUk8zTE8ArMQSR4XDoQTDNy56Y7Gwz//ZbCQ9+9iQB8cOc
tUzo8AC5VzmtsWmiRK1wfW/Eq2c/Mbs3Qfw3WwwGKYRGNvjtPEacjV9FuK27Ou5ozHWrE+jVvMlP
YFN6KYb+mlFhayzIV8P2HMAaHTh9OpFeHM7d2vDjl+h4edDYZE/wm9m/1tk/I5nUnPXfacBcMuVP
hORDoCWk7/j3z4v6sLrXH4ZatBJqwYTxvdT0kkF6rctvQjnLI2jtLTkhhJiGysM/P13U8TTOoRgk
DIpl4OrNRRlcoIpmGffvUmTLjdirD9E8iNqbTt+mldyafTrMQ9q1vseoRttZ8ymizh0zgeWfoPSS
ozYxSHHdfnMP4WNAV8nWzqSM3rjgv0I1l0qvyfdV5Dw+fqC2kzZBgHKh7LdBeC9FywdRoT1+N5+O
olz4QSIwF4fai9d6XKcnGGdJYDunBVDlLFBQKNZgtj19x7rMW1kHTn4ambth1tuhp8XL9jtTUiyW
pRBMX+Pk7OsG5YvtA0faqPnWdDN8uB78/rPk3YVLlcEKJUUrjHt8rS/ghjSerAUGGzv7RwgJwYva
gnfvJ2z0Nf80Hlhs1BM6ri++O5jKeywxz/dTwk7rrOzDI07NNeUJm13GGUbMWxE579YlAjHYX6KO
8a6jX3JK9T5fY6f8SUTDfriw24YBWVpCMc7fHWf7oNDDqeQNJ7i2ZjZoNe2ZY1HvauCMtZl/QFQ8
isVMtnrnR2AUn3VQJ5pAkIUBbgR5fZd5YkiRm22PDKdVvsOLcReDGBqiogFXy7rXfHO9AdsA/t2A
Avbrp3Lz9025KHaHf+/naqWThu9z4/bMZ94gq9d+az3716p6Av8+LDGW1EHVvu4VH7aVmP4PahWL
l655o17coQNTvQVMMVlcRlb206f6jGS4FYUpA23MMpYvULShpr4YX7u3lgGz899mT38vd9LEKHq0
ArkdEh8egoLf+YMphZQ3/Xw/aOcE38hHKblV4IYFy1ro4v8ZHkFQCVF57JW93iBddGEHdJkHVMVx
sSOPRYWKB89BzTyIIuR4ahjW0VeMKQsZBVmtZEpbH1K0PZSybeDKMyanufKO76l3WLJbPzjZGQqq
2FEHWVVe1rmXX6lJ4ruAa6wwrJVPv4z1SeEEqsGb0vDgQfY+sCtErjFumonpnEtnCxrzJNitTSY2
xwzYdFtW428PpFkx2SZaUq9mXnCb5AVfEg9mf9u2FMkCRRn8tohzyJ/mn45vvlKE7WaHYdUaZTFN
AeFT565f9WhrBr4THfh4AzakI2frr6RjL02JVY4uc+aGY/e8azT760MNOEhwO6a6FS+bv1Nl2Ohu
3dBLtfvmngH7iEToaa71lqEFJ5n0MU4p5QWOFKd2OeCGJttDPyezpLJyBg0I1NVzeEurO4Dd0Yi9
YdjjaNimDDp0KUH9bbOX+lthKIoqEDvxnRs5dlBGWb5zmiWVjLMaPQeqSy9+1vqjQHyHpzKkXKZ1
ixcFX7lFww21lHe+foHYvXvqwq5/A/7ZFV9Y4NMtY89IbYrVQb0co2qzM8oqreca91JGWI6k6PMB
G96v26DLuDwWNl633BlnDOo3GDB6svVDmi7tYQpKdbXjVRe1cLcKHj2TVHzopZLGQqHc65qOEB8f
GYjPYeeWrYUmX5ZiNG4C9aMnWyvNXPUZHLpiySQ9sBDoyvr03HW3CIqw4sqQPBL+Z1CPVrKdO8op
Hasy1771Bhm8R3RoIOqAEuAQFERhe2DQ5XoHHKsuSJ/hFW8qdHl/LYym/uPlknExTFsCw1DexHox
yRnFHbNLHaAW7a+Dj/tI2/SZjj7tc3JHSLkaPcF45t6IPKx6lJVgZTHjPfViSNrwmlP3zxp8LS8m
VvP08wsNkgfXu7h/QcEVQ4LnTflqolbvsT1VhbrOqWXfvOxHw9/y3ucDSRD/uUkIBj/vZlhu98F+
fjcvO3bpxBXXs3C11J88mY/YiTc9VlTzmheMWY90P6xh1QzjO0NzeeIhTv6ivdGt7S8SNVbPAvjs
znNc8S8f8n6sItqhPZnJGT+8mO3os2DMQrdSta1OSaTNyDADHRt5yMAdubRs1vK8IFep5NwvTOFY
bIZPvdJtIU7xTgAG0TBOHaS03FjKv8bCPbtIymV3wM6ZAghDmgt5z9CDE9i6vxDTdfA8WL+gENcY
BR7if+0tydEEg4UM9jLSDVS9BMVJei9AHwdwYhsUDhehCa7mp1a5UoZ1K+rCu2CJE0WscPnbgpzm
3A34yPBZjGt1UJsZ8RR+OomBOOOvjFJg27ui/kjsGfs8RWK9ePlnRWS9M7Vs0/C33Mwoubp1WTl2
v070S5tMI0hAqJ4xGe9TukwKuPeYmBir7zqVQHaK2A8syUc3k+UzjZnl7O0OtYWJC/Crv0nfDgSD
4AxcYmPdsg/oj6Ap2bhxr2rYRdI11qDI9j87xVrGTqWqe/HiMiO5nBFxEf+7FRw1f6SNGrpEBzUh
1inVT3YaA7+ROybGg+9aYV/NeIQWIN6GVNh/pHHYpg4GKQVQkIQTeWAbTmT3t7irU7ppL6Mni2Ty
PP6Inb/xZA5RCenZ8hXz0KF4sby8j+Ku2Ig8lYEU/7U4nqrQ41GNYM7qZ31IJOtMze2xHNazAZCx
Y73euz85EBoggW2FRHBorFAsik+qIF2RH7LEzj75PgZykFg6dv0DwpO6CUEODdfUNtGhqHNgyF3L
0TdYxUHzejQ+KKDm4/livfAOWura7TN8M+gp2T1t5Mf3qvxzOjukCPraRc3v9ML7/WjXdJpwanE1
vlKyGG6OkbqG+V9Jo5KtcBHmwgRmziEw7P9GlHZjOuwAvDTgc67WTiV00msUuxpSgfpRlWFkKIyJ
3tU7ztBDo4i3ULrx2A7bEIfTqaZ/UJh8xINKm1vVrXJRSOmsHuD/Ahcw9w7bbE4yND6cMwcKpkBu
MMBfs79CsGzJrHN2Bc2w5FO4ugq8f4VH9dxt+NCv743y/bSirBLxZN/IFYEHlfZStMLWpycPeCLe
f5R4KUxv8q2uWLqgGUOMQ91WdvTXgYxzTdTr0HXjWWrgFiND3fm8isonrjqbnKpvygOCRWHDe6F5
oBCKpnbBHNG+0uUZ2NtQEUm0qHQAEJw2M1hwjxPFyuft3rdSwSEua5/5PCeOgvY6wLd7SjXduMVG
5B9hfNEqUxSQXp0rfKiHeIHVqZVBKpGa3P8iOgk8+qkktImGAvw6Um7Cmg18qbmvg+p+aCKQl7vE
0jzRHwGMwQjZ+XzsALHblPLrk1PvLz1BSxR+vl0k2/UUudHFmKeXAyYkTC+F0CzXlCzV8JpkyQFL
yqX0hBBss9vdQcGS2xdPZR8XMTTBCUJATOzmlU5jtzoeUS1TBvgqgvKVrtsHCqvI8OeHDCkVvChQ
EUP+sxgyzrxIpg62SBNiVrxzL9GrJ4W/ZTlQaESzun50oBXywd2Q7lEhGXJsObnIJ7s1mxtN4q3Z
qUvBMQHiPjssZVsDUS+X3g84aTyzj490owFCsfztKhfEjRdApjA8B1IMcSCU7V5gP2aH2uVFXkkA
74OxR5zlQp7bZkv0AH7qjweR2bERcLra9jrrnzTHU5zhni9Q6wtciw7HO8Wy4WlUhXPRvLKBHmiE
xL95XaqolOaVgfqOlCFxxXe033RhrdwJGdladG4bmKEEh2uzbBFwEcCGJW70LKav/BWXXrtDTOiK
hRaqYakHWCQ2z2Q7jRCVp2EUjj8a8Qv8nmICG1pWCK86qTPQpHEKg75AHxbjd4CXe+D5mLcc2zvC
BwSqPzjDP0xcDYrGQQi8vf+6t5pWa8JgMcGfv4rGq5/F3YpAb4hFLbjXXhVePVdiYu0X2agBxdOI
PoKlvGIMI/ErXtD6fKUc6DFopI8rXc/Opylv/oinmRvIOXUuFqGifc26h3GIpRkmM9NmmO2SRDjM
seB3YVoTsjHiEXNHx6sl7Z8EOsomeju/WpcLOeq+qZULsnW7yDzZQ6Ag6WlwpUaFKUkaQ8MRpWUr
YmtJf8LdFwMqPf71HklktDK6jDoyCOC15FD2Rgx2J9XQ5qSyfVvlsFutlkWrY9Fb1GQ2XEuHLQvH
dWz9uzlGqoeaFiy1BiZUTxgEnV50IsYYXzPiLzA4tDcv/FLc5IdZ1UraSKoKqMhV5gpfmvNSO1bQ
OCYBJZtQHNQSiFCaOChG+utZFK4iF0zKUrg7P/R59krMmS7d3odiff4ob0sWf7z5fntNUXh1NYqJ
aKbZsvnfA/NLSAj/wH8Ec3ac0v/F5iGMHNnr9cloanFX4WDwuLagKRMj26/NtrzH0TJdMAgqZAq1
RnVACqCtB0Ko4OW/DIxtkVvshGVFMvKLRsMmRV7Rp8wdgP2N1+nsLeFI9eCZDrNt7LmiZ1Vj5Svl
058l+pHt9pg23jWc2ys0THKjEGUIDlpA3bYf1O4vE1lKhUXBR+6fA8j45gytbvZH298PBCg+cDAU
loWiLVN4HxPBjoqZ9u1H4T5cowRkzd5gB0Ym+9qqBx4NmZrpGo6jYQAP//GZIL1Jdo5ExtIMuVjy
I/brNrJVeE3ShCb7ih5MeDYU130Qih5dAhYW76vFKy3dkrunnLtTGW5RzrITKV0HWcJBfn6aNe5i
+jgFWYkU0bS1C3nKxERq4PaImrBYDj5z5BrVYUbvBus7YGUTuI9Qa2YPngPo5Efec/HDHUm7+ttb
01SLZGRx8TFDwK1LDSlm6/HkmSgwB2Z/3ki8PAHwhWLcOVhlNi2RwAT3HrwoBtOq/wNVOIvUvkwn
J3hjb0zYYwO/Ho7AkeYePcnenR4KzBLqUQSc/lUSxx8ijMNuE5vlfDS2x2kWpe4qjjWH3vKhxMnT
RdFWgwa+kvYc3F6zj4AEEnV+iURr7aha9Lk6uYMy2XUFl4fUDcA1e19HrfX0gZkypoX/gKoBRunE
ZKECnvWkIFsU1UEAwV2tDr9j+3O6LsQAspK1A1+i5FnQcHECa7tQpCIXNd2zwmyW1n3KHqoOp6CD
r5NCjWkta33YXQMIteQQ9mmzazgp/pBrVIzyumsSnHhJNFB5S/DeNKNXiwigNZEDDbSlA+Dj4pP0
6JysS0wU7gqoDuiKW3t+CIS1EpGBKJyBWSfA9mYhukYY25cW7UxLJwK6kvN3nA2xl2KmA8wCQ6rI
aytjugvKjWyhoE7KKbGwPHsXerBJJA9gK3HkCokeyX4J30+DK/w22AhgAPZ2HZRms2RWGDfFbOdy
FVZ3EXP/rTld6I2ZVtwbNanctLKJw+Uv5TTqoLZR5o1r0C5FKp2jHEOBDSchI6k5BHfwj0sUWVJ6
Oy/Wks0JiWn/5+mjAFF3SosHGuIhbsfcKHNmXLHFT8TAbUKEHAdSc4WvQM1Yo/GnDyjpiJpEvwIR
iYXRwdL2v0aqImHg+JeIkdD62dfW3/DJjh0wXIFbKKcKCnIRVyiFSbByqgcs9VC7MXHfaOKrGghw
naOath3831L3NiSdSal2S9CykP3/p47oIDxSlxQaL1xH4HepmgjEkqnFfOeVplmIR7D8dLUiieoT
YP+YWegzEQkSY/002kmXe03U0/gm7p9uDEefv7dFotx5m09igTRzXI8V/MGNR4K9so7zzfDlq/UW
+nxSlYY1eCXnt2gOQroNMv14gmFmCYreOvrQyq11zyHrOtaUupqyZIKi0xdMex2b4qH14IONcnmB
Jjqr1XnSHkn8UUvP0vKk3CFFIMl2fHIRvQQvcwGfN5yYn8pu3xVuRb5XdIAmFBP3hrr6tTUV4XHM
fbJurfTHsJYiJceKa3xi1h40QjckD1gwUcUUcakr6bL79G3QlffgEVkgl0vLw61EtdpCkEN2W3XN
2qO51pS3tDmWysYX+ryKDktfQY6rCr25ZfaLBhR+0mCUbp+CmrtmzeDCVvL7A/+N9owEprHJ+E4L
y7AlIcHX9rIJL52BbKMLDFUFWcKzPMbn0fA7KpVBqz84VxbD7vuw3Aj+I6UrjKmulta0R2+XMw+9
ILsbPrVAbEc0d7kynXC75nL4CPnwUBkWNjV+kB4cjOoAOsii1y/Fodwx6gQ/Cm3xWM8qX9Zp6s/T
E8NI96Y8XdjXfMYJb8+6NsAJjNVWGdtNkdXaoGz+FVDpKmzMWTv2LZwTw4AV+rtd7ntWTa2Zg/m6
NdXLZygFdrDjjPd24us298dv6gb7dHNmqDpJCVxSz+Z+T/Lxr4Mhhd7xyz9zrmWQoi6j/QjeG4IN
ot1j68TXgeDTnI96tzEuet6Pph2tJK3j9rzlSBSiFdRa5I42+ikVg46XWxNerhK9tHn7NtIfjNvX
4VaoQUbSOD02kCMpnNxo67+9lnrzokd5BTibN0ii5yHsWrYdpRPKpiFSfopqFcDzkOvf0PZtdHYS
rAV8in4Qt07iLvFNt01swdjxtmBxRhyqievUNQ8l8e/cDF4tzLWVyfmHJZCLcritkt0/f17L+vjq
4ZAe+ZAA+ywzn4jd2uQALz84c/OLDitmYkh3HUEn1PwK1GcccgzbB+exFFqEQ1qw38dnbw08i01D
BmAZLo4J5pJtITnRfcbfzk7A9uyAFs6XzlKgj1cSh/nAOu3JA83+MU/FXpf6Swz2afbxjM05H4+H
g9eD0h9PRjQ3FKK8/Tpz+zJOR4fRWTt84bw3yBaEMwL5Itn0CrNuj3NRgyfL/rC6mPQOJ4FmIb51
tqYSk1ybioD1iziGzxSntcti1WZiIbYXLQ9sw5yT3FwORCjGAGiV1IGPUAZHIiX7u9AxOOAtA5Aw
7CbB7hzUq4LkJM1TDIKnaNcqs7P2Rw9PuyBQ+3SnQu4YAgvafc1UIgHC9R83VlZb1HBaMjlN0lK4
sJYoS9JwaoqbpDjhNcUlbusTuLROpSCcz7GfZPhBo6ueL93F6bXIfaeNAGGJJlkO13dZJ3uuAsbG
RVsk1omkDK6y8x+6kiIuV8Fm/vvk+GUN34AVSToNyKKtBEMtHojhOBKQHhgkN6vWcg80pJlEgQIH
6BUMqVP+ewPgTouSOOGfqh/kXyknqg6yJFWH7HrRnJitPuusHgMa0AmNYU2PxoFB8T4Pg5SDZJfY
IvlSpeakFW+ZPnDL7lmn+jiCZButPX0K/zVqkIZuhAgCXDGDykc9gqnjuvnfCGkQ73JZMDauintY
1/GI+EmoUwePFCuw5zOuG098zdSIYTn3cOuhk3rCj5ursXLpYPRpg5IqwBPzYSfCiDM3I3gT9YOL
dMXIWU7qAxVe7GCQO7SV9qe/siXGNALGEuJfXSt4UtDCd4fodvzf4FrCE6vcYcbM9AxtEcbD36YW
H1k0DtLoovqcCNIbiZDPeWa9qTxtlRgPvJAGIk39eMW9j/rKlh0WLsa0PnS1Wg8r0x0onbI4k586
hXa2bSzzqWmYHvSLlqW6SiH1+66DISZsRCbvNDqMJSFXIjYUU9qVWgC64kT8fI0Cgitoj0IoX20w
5z9ZxOHVvUVtbk2pttwYSanAIKqYKiiyZPIBbM4S7BcgVwyqMFeXfFc2UDlnWrYKDjpbpapOrNp4
NHOHg3YjJIMSTvp3kf+piPNlK//a5fk7sdzbFe1PJeN42Wm+cUCYbk6AIJt3ENkdRLyCojHaWTVK
WoI57HVdRr1IrSfg71ee/iVsDc8bi1XAgnCjjbAfA7q5N6wujYC7b4+2c5VTzGPV+F+fhDKmEE/O
9laitjF7AZB0y8y9nPCYp6scYwHerFrs65aICbtwUO58MzbeD6paTddMiEvxrbnJ8O/NNEmYmJBR
FCadqu+4Wmlx08hxIEdBITDftlTX8SLyiwdVpRMSQINR99TFgD6D5S78IvoKQowdd54ooxw7/Gq1
smWYB2tcevdsQvZkDCIwqZydhWrYH0Y7QFctgsf8vOwuQN5MPN4QIGyKlsKmcECZQmKf5tO3sUM1
7EpgZ8hn2PNalDrO/9EEpRJ2BBW1aJXZWPFYofCb2qKbEBuZUfSntU3ZmIwKHf/93WN3M07ardyu
ukfbXheEYboeUIHSLKjGg6aEFsM4W6fk1cG7oVIdOM2FqABtGxjhgtm78CCGm09yOehz5ASa0r/q
umDozdgPd8k1cKqF5T34jorPeSVrfXwWn3B4XHqbtDVR44kAPUXHamJXrFlQglL1zCI02DYKTgLH
wWzhBda4qAURIDEsQRXCMp1MToi++69Xh3GuypBOCpaato97+xzhWTQ4NVySnjpSLk9d05xGalLv
RX92XQvPRn6RLQa57QHh8qfLirpHW5mgjPzOAHpTBvfeRfnsFceS0O20fZzGIJm0eDpf4skRKbhk
MNfHV3T/3g25LD8yUT7dop4GdOM1yc50UA0ZyOfYHGGn2Gtkac4hCdAOZ85u2uo5SV1xoYCRLSwQ
ioT7Ty9zyjfQJ3TvCqQVfVWPMCFqXVwDGBTrdb64GebSFotCUX2yXkAjQJqim56w1d/x/ibzzKGR
TMKO/icCPeo25IGkPcVmPMUFNRs/e8LBKIMt20vQC/zx1SHBS5P07f5OjoAs+1VGkQYwRMqbgpoI
Q21Q7IL7twIBo2vIeKMW1CpDvdgRZIRMNP7WnxK2ka+0vBdKp1SrkuTV1R0iQEPRNsxwGGUpOdKS
8qenm5LzsE7Rt+q+QyhBsiN+v+iSZ9cHCh/7owQlbi2OzcDbrv57AS5ta/HtyjPZynHF2moBOCgX
Lok031qwhsiWf33FS+RRFFu1z7qBfeYuJltVeHZg0cC1mtJ4PKlEN9gep/4dbRW8L5i9SNHY4ox1
jfGHw1gtFc2Hra06DHI6/lULZx7PkJJv7LXWMpfyLTNk10uhBFqQYwWGwVjeyt9QfRKxCZIYvHCa
Nl3M5f8rviCEEl9imezigZzw5QiaqbZwkHEvuLHqAqN6klYAEGRl/ipx/jtXHwpariIG7++KsVwc
PdIqPPTWhPILeLim0qL2ekaw4k0zU5PpDMCaMxcpqWQqhFhdk4ci45DHz5dp7DL1PUU8CwRTfHLY
HVBVHoNjO0yfcpqvGTZOT+98BMJVGTNR5/6lZlXwFquneuv61Extl0bm9+O80W2HeqznIzREXWIq
x/pJGaBBOz/2gSI7gTlv+xr//X6IecNOH0LMQ7ettzSxkNCXoN4ZdNalDayYesl3AhF/7AJc6TLv
lPHAh9iFvcNPyX5UMqYYQ/2iC6smmsVBSET9nAeq9EQT0hY0u1RZgV1JSmNR9eXbGO/wh2NlLYDd
hGlRpfL7+bhj+3C4t7lhq/KduQJot4mQa4du70A+ij3PvpTpbHS0A/04v+5x/1pfV4MD8JxTR53N
p6xc96NYeOQG+ggfTSIWQRWoSemRtSQJLOFk4hekgQrwtqsP4ovE7RUGCcqopZxlu6ndhBJRf7dq
JYF+PgJAc9Q2nifUTq5GCtzX+cOAc8umWmbdr0YvQccPEoGrOOU58nAuNCj+6VVNKolpgQppW1Qp
0VjKDLNSod47wzQIfg4L3uvClAdgnE7ycZ3Q1tINyry9RX1Yjm5777mzLfsPGrt5naq0ri1IGPWw
sR6Eb83I+uNPoOROhrVyzAm2mU2ou970ab8HH8k/Sy8bgwwVqUos8c2IgGx6BWJyAM67WxUY68fz
mvWlPZ8YanoHYy8oiwsTXUwGp1alFit7ZmLQjVxPoSrXCV6i9TtX1MLlCbIwh72DWBsBh2Kh+6xt
COzCCyWWrX+JkZ8FJkKuIrloH/3TlAVy7LKAD4nk7pT8mpbFC2PVL6ibvndEQSVs/u84HCFosXAA
SekJXZtcyy1vSFHHFuSGj7/4vfQXINCEB7FXh/heqvHRrTwfR8hGS1oheKpC+zBnolsYCrcfEb7k
2D7aL1jmDEbcXUMbkARDPPJqcmwQs2c8wv3njgzUrNW5d+tD7IfDrK0nYk4AGuv5paKroDxibkuG
1r7iGqytLRHfcNx73YMlxxFropfo1TOoa9awyNSYJuzwYTy+9oUsSLhkTqTIRibdNxTyxZzzBWwO
Yp5qo+91AZEN/cN4ZiweF8IGVUgkm0rKGAeIpd2kzzvpNjch8na2TXNQdH1lDBLJ7mEpIXaqFKxb
fExGJ7h1LojCCEV2MEGK/lErKJbkJTTyJSpuAL+VpeYzkOWxgOmIwAYZe72XBceo5VXFodIWC+a6
2fPDOD3ab9QR15PuhhBlDfaBug/Nl4MPiUi3kV7T+1zhST0fZSc7onNTZfeYHGmkdawNZDZInoJE
ENDGGgtCGVfpkMIOIsNP8tGkTFIwAD8ERBFzdwGjioWpRu2lfyJWN8lBdJC+KuqFFxZFkqe7OblL
GVTetUTjApc9g0u88E65UGdavlyqem5hZy9AaokgCgTIFykbeHK2SPjZ60se3QYz5uEmEpiomb/B
vvu9YMWJQH3528AcxytiAMYBGuC+/erE/W4gu6sjDQX+a6HA/GLClce2uazg0CWnctysRrx33w0y
f/r97YSTdBGgQodayPwwRFzMlslFb0xMsCIl8f1rMlbU8yaIiw88wjpbIwqog+NfhNuwsA+QcE0z
piza+Fwq4YZHXRPrRk70b/iJUAIolEyRuVvcQyfoWP6u7pWzF4wJaLfw1xOOUY5nIfx4UkR6ubaq
TgoW6+enf/9VhZApFalw32kbwfYZ+k8eJm/Yu3zK8lSSTCuimLe5rELCRef7PlrA37fAT3WcBsSD
v/NHXctUNTQ48tTiZgul3CbuUS7GTP/gGqqbVAj7XbE0MPPH6XNsu/lqEvA17lQZ9uqPeecfqOEl
sOmbUwkI9bWWYUTiLlKN/j+9yl6B0whi+oOKQN8WzYyDAOfD2jiMjlXKJZQSTuflIqT1Y+2JerPI
NL019krw0+iqz2EjuL296u9N4AFv/q6gHl5/mZ3cLAeNE5vOx+1lcHs4Y5w5IApIbJfBw+VHQhBq
9NEb8+GCZ+EML9n3HNtGslNxdKadaniQsfQ0JwV+L6h2ec/DHAaNpMyK3vTXMunYZVdFxjHKUdfn
ArP7SqILhXqiyi/BuyMaLTjAYzHbvOw2pzPCAnsrH90M491xNL2qHG5w06yjPLukmLCGqIiA3Ylm
u2VCAc3IMlQjIqiEVzGiGM+MIO5oWJ0jgPpyiUYhqXsdOFxfQY26BaAnp2V2+8cPOMqSjPEN5LCJ
nZ+x9vB+G+2h9nLryxuZzKxVv8aOeerrniQKZqzK84SHMYsRBxDXUEdXbXsurSvPswh72evUqAqY
AgTIN9/5NUZ034upMXxTZYpsKuvzGV/wsJ0bmydGuLCw5qa/HX3lBMXxl4SG1ZJC93d2Y8w8bS4h
zZDnyRszvd9rVe1t8L0OBtHt5cv3TM2JHwaIQDot9BiS7WkM7x/38Oe2vPah5YdXl0hVlKwthwzA
b6d2w36eFTfZbEzke50/fuuTi8la653APoeFi0FdgPCbM9KFihfs4vkB+Al5dEWQLkp7adPZ9rzy
aUDo34d2LKPlP6OVPXuM4LDWTv/imklpgvVL/ctWKqOq8ADCdbm13OZnG06k/Z1Yx9PGyW8dbmuL
T6Bg2sysF7eImNSF0oow6D0d9l/AczqUNM5KNPUHkSjDlvJgWCikuLVBSpUTFjzqnr1SHOHRiyPa
oDiUa+7YUhOvd8jsvxsHpwfzv+4JccOVLIN81iYLcH3Tvl5tBNe1HulTj8/rqUUlhKBDJlhJjT7S
wfXwB6FisCJgvz29Klcm3h2g5tTP9YswA+MscIJLMlKhjcT1LFPDujl/zVk7nwo+QD5fbGkdPCiB
209fvNbuCNfwgN787j9NLL38D54NBueCChIom6bOpcukmqbxUmxB7g03cUCLTjrnS6iwZBSIpwqp
uqKOgtCldeEhPcFGx64hfHsyXZo2ghStkhxM08d5zjtGbVsucnXb3LOP9DTZyMGvaGK1Dg6skfSu
TnwRhLro6C8ycqGE63vXVqTdwsgd1xGMkPIBB2WsgZilkBMPTDdf3HIe8N2DHwD1JheBLQfaAlVP
LTxBTlW4Mw1iO1vpeQoXJDCcW4F19PMf04yoikmHbylQikU9CL3/1c8R2XMXLIbKzzvkUfY8xJEW
SfbNziKU/tiqIwPPbCQ+ScgzJJvLm7mWbUTkOVGlCsWpec5BfE+cPjvbwiwfs6lIpd/Z2pE6k9ao
8nn9gIwAQMBl4BlcMiI4CPIdTQjAO9hEzsllq31KhrBiueK2EMWKVFC6WTya7rRfukrUs39cpzet
Ze3P8cX1j/6l/mkk56kg435AkLfYxis3YhfEX8ceX8sUW/YOYAI8s/uxZ0qLa//zsxIhM69h4ptF
lTyYWlCdEC/FhB2/9Q1g6i4ziOfZvqndCk3FkxQ9RMmt44msWYbhcddjD3azvCKFoxYI9gHeYNnT
DFE9R5ku8pdvHV6QyDdqR52P6WfHmrA/KmU5ywhlZp9Mdaj/g/P5+ZhCnw4BacSDIdFc2MmhHZ9W
rbMbmmmKNd2zTzvcdvwkwHySw6gOQb4yra17ZhBFjC7z9FaDNnB4SrO/AkdJnngDYE+Di8mWOBD0
4q5U6prJbSUSYjudFaZjDC7XyMibv9WjJItJaA8nUheIZdWeLjlLJCNtDdjxXJ29iG9m4Ht3+cxr
lbyjJOXhYlyY25J+GCP6ocUHu/hgHJqPYWEJ7A1BSwCo/FTlxJhvV5SviTNjzG5cSlF0/nYtP/7X
bqhan24cmdL3toLhHBRPfkRfT7a+DyA61dh2/YSuiSIxtVlGVPUBsDSL2/pCPiSZDk0gZENhTics
XhwIWXd1S+kNJ/sz+OsEf1FaIZQl0eCoH1dwv0rxSHrAAtfI7Mrtu9mt0Pv7rivGY+e94OsjXgyu
nksKr267pilokUlWgRW0zZXe7Vv5q6Xg0Z+uxn3OpyEkeHv68iwiG7kI+gWhoAAhPxWDWgL+fRJ3
tAXP7aMjRGBlM0ccrRkypuSix+Phq1foDoJa1RRlRAVdKxN1X9jNNVEzAdaQWICluN66l4AYSTtZ
1urxVV84FloKes8heyusXzkFCCJXlxecRmmFwMn7CLMW1ytOAF2fnCZeDxvUk3KJpKdVBnBOEFbS
2s0KzVucSF+QqslODy9prLUatS69BrZA0Okbx4Ybcmups9vjBDkvHk0MPxsDexRhk35HQNiKYltJ
MCQNc4BQZStqPhcDWvpfaMxM/h6VmmWfbADd1hyJvRMCHmWgcfS5ATPAjX40mscD2wsKHNege++s
LNUfAYSGaeSwNpy0EYf5BFOSTFzvLsvfeb1SAH1ApKXzSpt7gW1qho/bYmsQZ8LVT9c+AnY7SIa4
958sj5lQKFI/NIPV7WSWdLE/BMibpv5ei1DA9XcYrFd2UOqNTKQdfTSTFvgnI8uZbQ5M6c8X0pDz
6GzLgniJmG510WPhfY3StfgfuPsy+McrLCQY62XmIwtOThAO5Qh8eea6VE4g30YAoHc0uv1iOx5G
rWkYiAC32fAg8D3v0S+a4fMR3iBaxrSu2SHSe3c71KXonS4PDROMleYMmhNbvZIwmTDclmFwK3qB
V8sRayZZkctKNHDuMl2xbl4ue9vItc3dqeC3GqB5HZOnqSM87sVOYe2BcpnhXqy6DSSzjb9DbtId
GJ1jNXGUNzf/Gyzb8usDvhkQbXxwf0WYpB6xLRm1kX+HwIpNXKwHCY/qN7TlBmH3n4fgBUnWkKpm
dA49rL3R2QDwxSHfOjWET8ru2I7WVKXgkK3DEWfwt/D7i6nvv4qtV0cgE2sVdTfY8SCnuU6ROn6K
PyGLsM+MZbWxzi2sztTZ3d1VJ30m94wqZcSLcSJmxTNlg8Y4AC4zZJihlOCa5j3unSZlZSUj6Yco
RiXZJjcAHt8AmC6TswevYUEDRpe9rfx6ZhIbSwsivOaFDvGrq5u1vCpPPjuj/+EpiPOM3VONLLxR
N3wKP9W27qQOIL3cgKxlsLfBnFjelEQOX3Tv9tq0O9fwJjlEDswbGzyIMrpXBMqKdexWyCZspc3r
NSq/4mTqaD6ITaWAHPeltZXVbVtkhvAq57ajidWEI5yQsftW8oCAptpVV6F9vG+T3CiaV34RrfBY
ZJjXup8++hYJ7N3hEk/UerOr+5xbbTqFKPeRRYfTB/s40Jtyg/1rb0iz6EoW5vUoNnrrrhUECyB7
FlHvLMXYNEjImV0mrMNHbkA6yZwQExLR8iyyZ5zOqSrCyHvPmMjabYE3d3qMb2Qne9cgvISbmSV8
bjkqEqbBSR9eSk/ihgvpRCRUcjYE12KvNtsIGtcbvAKnKysuxi0VgeOT5T81Y8WFcUAGkvnJk0TW
NfS4uk4VU1ZZe7wlSGhXvjYBtbA5j7cZXKgFRzAHcAUDj1yg33h2SNJTFKJKR4olpgipCuHlOX6k
OrrPZaQGLfK5atDGmcMuPyh79UlrUHfYhbiOLpnP4vPAtVphsKqiV4MSHN3DExWv2RlS6Tz9zrPy
e4MhLLXKVvy2VeuIwyG/cqFhTka4W2DMKXKRCJUHd0ZgSyKpWoELNYPQk8TSa5XO/pc6yCQvCrqz
YnLILV4FCTZZVsLvQI/1SjtSw642cQ46uAX7QcZ7jG+ug/Ip10gn3leIDzmzbOIY2BhEbk1Ue8Af
z43RfIsKyR4+P5KPq/oLwMFYwV6BovHyBgjsJHEdiJhCGsmRXf9MuT2+CH9j7qOnoMOGLhthPTRw
EYUYcVJ9OuQIWu+D0pYVRjKroIiLZiPLs/jZmjsixjgnaY7ibLBztD5RLF/fH+JVB02iSC6ytNyZ
JbyEqXW3gN5sgjIKsK/Kx4LKX1aYOY8sewSt31o1aDhL8nD/9sijVB6Hs3bVllqbPT7yaJLe7UnD
47nrjh1nqZ0vWu/fGeFC4E3uWRE74xBXedaYAfvCAO0FINnACgLqLidb3ItbRMkzu/kGKh7ZFdiE
/+R76KRAAUJzsx8TWclxhehrDGANApt6XIVuSkLLbYNlWHzWnf9HQnkP5M58lZVyCgSRy/vRIezd
Hi+ZXMX8i6+D7FzeFraImX9rA7ibLU/elHo9ZA3CiCBdut8OhRvdPi4iU9CPD/SOYGXmsc1O58Yx
NiylXmUAB5L8wpYeMRoAnyblPAsOAshsJU/VgxUQmKasFWvd+WHNY8FINrQ5Xr1DLOrLvc2PuWbt
aBTY2FzJA9gYUT3OB9pizOHRMayBztGpRsKb0vMlTNUWWMgmBV/I5T95V1cPFC5uYUtnvHGLLyrY
DlLXOWerzTC67iawstNfUMPdPDFB9RbKZUvjWm1LYLQTI4CVZuwg3pVco0B/CxpgjreOK5ToxEaL
h96uEDMnJjSOIRvLUw1amy2dT4N/CrsXqKpMgksG23pKs4W5MFYynpczz/+UDNklWBRASiLJLtQ3
2p2OfWi7lFyXJZPRTmkaB9mPepEOSNRd6v1Mx0dEa8LMd9awJuTQcoQ5J2PyyhZojsPQ1iMAf2T1
qR1YW6DY9HBswNPBnhePQ18o//qrQKiiRiqpKFP00kEI+ktCBkcEs0KGoG1UiDP4M0bHc7plBUXi
/vmytV/XbRsPv4WcSz6rpSBr/5jwzadoBneBHrMFQ+ZSwcoJlXcKacQSY3WpCwssVsmkg11ZyLz6
nhE9JMgxUWFmPG6kSyHJ8AbiilzhvxRM9HsDEsFzeDCkxtPb7f/WDEp2c622gB+gl60quPR95YKY
zAMEha0Z9mrKLSFhM7PqfABc66s5QI/+2GIg3FMGW0hMx9DyqxdVtfk7m+uW+whkFCqqfK7dLoHX
gCXR0BRFEiwptEQXxxZS6k5ttu0+atSuOFBnwCxveSrRRCgA0DMZ4P9BSr+6aHN3SrKBemw+qXeM
VXH202xE1GNcHJhag715VKv8iK2owyXuQed6SCBvV77MYeouqmk+5qsZ4vH/GCBy2qzK9zGgPfRm
3iURwZEQm4MiZvUcOVYM7SC2MjbeexZXLrFhUSJ6yZ4IleD1aTSxjKhCq3DW4OtgmfK7KRyVYqB2
gHEs5qZKCL76t3tEgnJ91H3lBeMwhwI7qjrBZ5rT7uvHLLOsfT8zl337Ug7/g4v3Q11UdV6C7AtT
mZq912BYDc0hoTu3e0ozi7gtHQ8TJBe5A6mxQTt1ArHcRvl800Bph8QxL4HYkKk07/Y1CEiZSuRf
pMg6DmX+tANbswCV67iHdZcRyXsg1SDTOIFvvbhNx8hrdFVHnUjgjQRbSv8Gj5OVzbb35tC0UjYW
ZuZ7Cly964Ex43fouS8TI7jM4PZAxFJUl3YwEUWe3m5Sn9+3nTuq7xBpzUtTa4KHoxHEZRHwOMyz
VXLbXPK7uyw0/F7dHEnTeRHENduddLi7tPtRpzqQb5u1/oocEdGamaumN8YbI0/L5Zv7SEdF+sde
p6wr5EOnBXiHHUj9qyPInI3kkHz443EF96zZV8mRRBCbBbDj7GD6UJ8yd9+tYgJ/V0HT0VyZ2ZJd
pWc6E6BuxJxvZiF8AQuF8vWM4bJL5asZmAZA4eO9n3YTp8erAnMUwHiGKQCS4R3EYpA0CwlGFJZk
RomIEj26huDxuRb3A5CvLKjgJrDpB1JwE3i0qxC0U575uYhAmlzqK7qlwHgkY/hEOkwmbtZuzso8
cjGHLWAjX3tHLh8oX7s4LG0QP8yTmem0ej1s7Ik8I600fXGIb20wM8ETI6n5UYBVucphfJOQXCXH
i4eSE6YMGCFO2/go0o8p+pJldAkscHUbSxHWRJL3bE2NAeMnOdQsCmF1Q2IY+OGcyaTVvBToNlTO
uAsttDWF5jyK91V+z98+/K8kF60D4HsTJUgmPO/dXGGz7kDFmvWUD5Pkby1mbt3Kos3n/j/SYgLY
BRp7qbzCDhh+X/elb+/3T9StR4vWGVNss/GQhkyfSiaKLE0nObT3rtG5jgjlg1tTXYWSM13NBxqg
ji5uCIoB3ib61ZjIrTP2soGl5TI/XrwlFUDB/ZAJYV/PMSWrLHh99l4P2tuiJ5w48c3HVCROIPsT
vN/1Pjl3byW9gL//dEPeDPcFdiOHuUHDcHKynACmH6omLaYNnitqaJldCrtNJtdqO7v11jWwM9bq
TfQxbrE3ZVnXf1vmF4aglC2uIt1f0JD9uazNuuQk57LL8oBmG5SH/8F5ZA+cPX+wGPiALvIONiq/
cXdY+VjswVRTKBUWFDaPdl5Mi4NA9mw5XN8T/KGZ+tiVO1FCKDmhs3Ola7eXAkRJ2QWM2Vt2HGr1
di6xV4t8me7QPhJ+pHGc7saddBm7BxrjsYt2nQBkJeJ6dZVVej4+vZeUw70ZKel85JhZnTu6BG5a
Vx5QxXlIg+6a3lLn/O8rXH/lKjJ4oCWv2j0t8Ui2Gd7Tf72Kn4NDDcFSU24RUaSqQ8Q4qcJPjsxM
zPM6ab8rNcGev0AUBvBYcUmsK6Sv1ZlPGYZu/4M2VFRHyUTQ667+HB8/T+/i2kll+m9Spaqm5K1U
LJHd8RyI2/OIy2qFy291GDPtYp+YDs3AnFXXyJaSqiCPvI6mfT+LYWLcBSNT7lrxKFKBqiEARMOH
en7l4tQd8eJMw8gTRR4NfRxNWFIjRm9Ccm81MDNCkPXyBKMZv+LnuiFikpeZrB1lErMrsrtiMTbY
KJ6c+5qmSKSSRz7N+XRQtz29Loelerhe3Pi1H9daikKK3/XUsjYc8iKLDqxcS4VzZi0SjdNXY7zV
HPue3erKIteaOKiGfIpT+EmmTvOuidJoj3Bb7PpAk2xkFxO8Xq3X9/PyxXsjvtp4MpSAi7wHMWhj
uo/83+JW+qSKb9QB6sWqm1+MjKTHjRp/s6XsyUDFGtg4FWONqRz1lqNcVe755eTbZqreMrWNL2gb
fEviCLxwCRPJqLNqWXC2N32wbzkD/gRkJ7NZOQngeHpuoto/CInc5PscWtkPsCCvbJXEIXFmGxh5
0exFgOzcJRYwmKKGmldeNfZBMbON97MkC1fIzAjkvXZFnC/zr/5gMMTPKF9z0UJ5gA+isTw6IS1H
vOKePFIIELEB2i7/uz/MLIVIGPSeHV1MZv5DojBmENJ0uSXvoKXmaC9T+r5HASlPYwbr8Ip+4AEm
ggP2LXKIXhcNX3s+1sUL52EQq7aMdfSXBqJsA2mbCYQMabnY+Nq0nStwOA6nzWllSH88OUCY/QH3
ycdyLG/awkQf47TRNU19sV60gWW7AO5XPkgRUy3kfkvT43Nzexuc0Jd3/WGBFi3vR4ODPbAZX5CA
N39yda1Iu9ma++/S/ISuWZvBLsFZYH6RJt4Cj9V9W78VDlt/9I4dfRVJcx33Tq2LB28X2o6W54+4
Ls5K+3PCOkftFljUrEkYx9d1sM0fCa6fB4etJSruARuxv1eyfbQ9g0Eerpz65brgRljorHl+4u+u
XpzvsQU5bT08oBj6qBSm66wV12c2m/su6LDxWQgylo19bPmBHHe4kQf2C1gXH/YnxfhvPHfOJzUY
NJ6aMKkjRzfneZCbFBxURX7KqzY0LeEq90I6pP4/EX9nYGqPvsOL43YgMjbqRS9Q4Cm1/XNCl+B2
CVLhryW6n+yACctD69TOO75QZp+KBxcn78SmM6b66R4VQEqulVUD+kuexUJeCuY9ACs1EXaeJBzc
BD4EXR5sRz2ueoRZoRXhc+QzjLEzCnr24T2LToJOUqREFNmu1WTAUKBet0bDxXZl2MmEY0s4tiIH
N8Q7WL7BaXLxY/SzEacFd8E1f65IWgj8QX8PyGWExg21+kUmk7rT0R7ewDPhkBon3DS+TBiMVQ5t
rn1N+A6bAcdDCVV+ZQu2r9JfUTTxKOMvV/fdE0/p3pJdyeDK7x/I4gQKZwHztrnRJAF1mUJx2TzM
lcWf/Ta8WP3xqmq16+rmKeu+3gRcqKpSbMNZbNBii58BLEx/f7FRUPXFc+zJXLpUmu5sT4L/DMLG
WcML5i7m4PBxlr6PKxgx2px1eeCqvUU0/02Ts0k0bkhT5aIlWeStVteIJdaZvUXz1JqwYBXLhPS/
iLCHlRoGW5pmh5aXacp77oQi/SW1Gx4uOS2Z2vefIHjn1n+RIacWnUjC4ORZWJmcPV5u8Y7YTq2t
ZzRodm5nILR4iRBwUZE23Tn8lVB0jGsPzrrmRm6o0Lg1vMYZhsRMzB8SnDcICMnZCAR86oxlNFwG
QAhHzlJ+/9hF7FJgi/xCOAAz7QWifZC+WQATuP2sh2PgzYq1TY8tGHy9TvK9MOiIkxDluSrz0XWZ
+8N/76aSoWL4bcxE6SsLViMjemej4x548x/GRQ8UBm2RT74LyCjFi+7d9M9k9hpGw7o0vCg7Zss5
MEXbSZQ3GnpwjTv7EeAQygGFobClbNZAW7bjgKf9ZTLd9jqdBklgOrwomXGdndKy+Hi0bBau/Ibt
qGHHHz4c76zejK7/KqKmB1s+jPr8cfp9x7gL/t2ytvd/PCKTDBSEfWHSGKo1aYJCbANeYm+7NWUQ
J0jahCdOJ3Pu0wkbi/vE5A5rrLKiFkMfeRmmjPNyQhQ7fRQG0vbK+33T9P8Y0/2INXe++JRt43vq
6P6gFanZv+iX7/lY9pRl1Wg9tIOAZjqJ22k0pNwuGdBOiNy8bxsj63hr2jGsx4JT+ouf3KCrmCCo
SS1ic5syKHVVNfHF+ohqAh+v1UYIPuGbiBU2HVX/QW5aXByUAwQ8W/uJEFX7BV1mDwME0RaUWxvD
t5EQscG7tK4k+Qx92faPDhY2qhdYYGBz3LjjL4veJ8VqBblqNas+9ou+Lx02VK16YFbclVWIu9+i
xizfhDTPtSbXDup3dndElPh6kf+YbdDilibekAF7gFNvYbespczfxfh8dXa5VYAzx3Y/8mIYcXCy
+jHsmzyk/Fc0znOQy5rmtfHuKGPp70kPXzn+f3lsZBQtgEIF+svmFz3ulu2C4TJf5X1RNHBfUkyb
y8eaJsihCn0Zmy7qDO2uuNhlObmNsqTF5qbmfL08vQDkHEVhTom7a6RVWQrcYzN1Raeh+jw1PA3I
nnAReaPcF69D3a3esLT5vKwRjlgmoIlhkIq5JA4BUHD8Tg661CJ+08P8aF0h+PY2aFKgM9UGkHi3
OX2hjMmZEaAg/+WZja4tttySROtj68BpOrlBIw+HHctKtgA2A0+B8jeZ1KDDlE4wHQaiHRUG3xJ+
hPn+lw6t9PYRoQ9Vj9ycoyMvno8ovMXeWFwZjULB5zipO8Lfe4zRx5yf8bqQopktMYgzBmSrXF4f
sX788w28qCjQUuISSBNPDUQE9v4ZE0HFPnQO/UX0t1lHOmk8XgNkoYEwuwQb22ZYHymW5td7z+3j
cs0SW8+qcgDO+sp27w67MdaP3Y4PjKGvVqRHVyW1m6lrEg27E3ubix3D1/SPaUkuN/S/oO9p6yjr
rUdTPwpFEtzKneTmO51xsO6t8wXx6GexlrHLaQlIzFUtBPJgaKlNJ0jzGUeDp2RlA4wQhXm7Cgxp
O5SAWv7gdJqlXn3HHQ11PnIxyzAPu6+VAPui8l2oKiT6ARDPyUXlExhQ1gM2Bz6B3d6K6QSR4SpB
3Pn/W8Wu9VcW7eh/Kt6ba70d+pqZD2E2T+kf42RdYX0Fz7FtKf4+oDTX7ppFoxEyugQmJ1HaPFLb
wC1lS64g9qMwRIexpGxQuLii3NnChfscH8E5+g5MiwXRrIjj0it+U073VTj1UNLuE+Pq9QJGQSvL
yXSdbxBkFhSnU46dCapgFXjneSc7oOGoKzMvEbCTrQOgIWIHxZfJe/2R1fahyWIj0SzwWjDdQwUd
37f6Qd9sH+Yqv8MTQGgSM7GlD3DtjS6q3MG9lj/DzO1+bFtSgzs91T6XOMavZ6kDrSBAC5xchrWF
yM7kBhL106R9kcr1tGa+5oiAp8GdThEum9bui9p7ydBacnCjcjUUP0L6U414JTeEqrJaIc6OI6xz
sNcpndq1eKvfowM6S+qk2UuwFwu/QmWMIBJ7qb31bYA4XkgBE3YV4jNeh0sMEYHGDgIcgDejF6Yp
6h5uQR2F4+riwsmitkvNASaF3NFeqfdxnrzUS728s0mR/GOBN5KrvPR4lvK8FKLg4ED+VUFhr7Zh
JYMqeyyTfxpcrPRq8ggcLz0GqjI/kW9LmE4U6l5TOD+3zF/+3cMj78U9LoZgP5nhD32FR92oc6sE
+uMWlG4bilHrS3hZYq6zJhvbDkSJsLCnJtePohoFnCIoeT9QQnqPNIxAhRsjuIpHEk0lc9Za2386
8o6GGNOP4RHOhjMJxtycaMfSRLj29x69isKmohfEJodNTYO80SKIEJwHbb76DzXwiuhmystDiEbC
APKZG5ALeIYPzAt/R1wx6snfMDCMyCdDHoTolpf+NQLiiPDmJHgPjNrzYIVveu8HRwVyC1plBJGw
Y5R8yQ0d5Sdrx2pl5ittqMqx5naWIpB2KjyzwizD7sqPg1IA0XUER+1fV2TgPf/+1Jt2sidid5u0
ucskND4W8IGF86zhDXbfNCwS4TNwKMODLG8VnrJskrEj4GgVGUtR0zpRr4NelebBmp5Skl3zVSvt
WXFmWdrVQ+DGa6SUvAEMd6z7iyfsvmdixjBl6khS4N4goM6+1y49rp+iibgAQrL37FB3BvwBUdFe
Le20feGCLt9QLzyOuPsrtp/SPwKWkPbgVDeptUPKLd9/V7XTJmjoH7x7KDhqO6bCvBqWOqqO/g/P
8qLocDH954Ed19TipJN1/Q7VsvRvTVX3AS7w5j0Dwwl26nc788RxLUH9ShJebGLINQ2f0pnF+PoQ
y+j0XjGBnD1N95+Rd/LgWzhDsszLmXvobiRfCeqCR43Fs2bSuKV8o39pY1G4M1rjgcELbgH6rWq1
1U3QkuRdqs3zkziIYD2x9WeSidAjEQLtRvPDpZoR2/RIS2nPIAgUQoT8HnP6iAFOa4qbKdAB49Cp
1es+Zg2Nojpx+424jXN+qwrJ91xlsCtb1YqOU5IJ0xf1fUXh03WE4CIere3E1mrv3nNqBEhshY1T
fPwVvDUR0vumPlyjok7HFDX3LqnEhG/IKbR5fuDEcV29JGwu+ESFuo/Txa1XpJctqzzSlaF3NpjN
nhnLKAI7U3nydG/Ap1pkPulo7TS/n76V0lBpZcwMSnSVGocTI1PcIMcqK5MB66y+9A3UZqUCCxG9
/dwnqIWOoaBOUnfVySIBSR/vhYzLJPqyGWtNyTMrRXa/G5u1IXoewXA8EsiSH56YodFaSppBhMol
FTrttV0zQ2u/IkiSR09o1FmWE9ZK8PyLvb1JcR/KP3tIYV8Rmtvn9ci3/UOWw7pcHsdEnOfGrQzQ
Hx6AWQy/C5G0eIbjsIba3nCHu3rGiLx0Zv7LaSN4evERaG9OOKfcbOLnEk4sb1tycwtkbw2V8MBb
31KScsAI+osuVcmVNCpfM2j1AAEryhUYHWzMwC4s1pb5rW5JIAn55yULAmhfyDHuQferwaPnHMgX
iEFgzlLyy3hEXgK1J9W65gMDzEqHaHtKlK7lHFv+qpwxS6fsGY+GyMeOrEYkSnclLWGl0x92y2Pk
RMpNGQhf09RaWg5kFzj7u/DyNsGqyq8C+EV16NB1qqqjvMPoLQD3Xu5XLU0fq7mpPgl+R0KJo0zz
Cb18R4EIqPWICNBPsyweslN27uX67oZ/X+R86xkxzdNZWzBc1Bw1hq+Y6QOrLpNMVeW8FiDAgUh5
Q6kGgG5oVLbBsrmWFq4PKADLKexvEIS90gEf6DhTg9RC4wHl7xxdsR8yEwxeigLvNJKpkA4U7O2t
npFQjAiYFD8e2jliPrkIZeMORw17klbgYJLEHtLjtWLRD/tdW+uXym6xeKzIvkc24W0ieAv9Vw6/
wCSZ5w6BkO2pjlKWotJacdFsl0VABEOiz+4oE2uS9bLzb+fZAkZW0NruGHTMwfHVf4b/r+sn9jKj
PIl2IPiLidw0/1zvK1rPaUA18g+p5tkAzwsMpBEx4svF6lTju8MNCTfH+eExVIZMj03x64kIiqkM
AFlLIe86Mzwkn6yRs/pN8R/rEGeqMlvSd5VfmSLt+ilVklpj6bZwrsFwOacBZJbMvoQqNbzJpSLz
FB28o+YOE6GA+tCOZitmlWnEbLrgKZs75TtSZK/+GqikgmAUbwKzqBwqVQM6Kp/OG1vmQ3Of2cHE
FvKELRZZgkXzlx2fJjEmEqvbSA1YIMFuS60TiWdX/INz/2m/Pij2a1fScIKkOqR/1IaevqImS5WJ
v8s+7JzyjA7MndRVZ+Q/Y566fdBUBrZOk1m5a4UC3lpOpyPVALufOtytL3gfcFn8AgsMik+m1Zb8
UGlJ/zrFLQkaEDv3/Sy796aqk7KRyU0pBHed7Ui4duj83SaFNvlNmST88UywD3vAa+CtnEmsJxnh
oPVilkFL1psYHGpOooecID17YaitObKKIo47cLSQh9VR2jXV0vLxDE3oBS+1A4ve7PM5G3qGsvDQ
GGnZeaKW8z21CKnAuZ6PlnqRo6pASibLCrTGMk0n764SXICGrX6O+7NxX1wZouaTV9IRKpdZP/7v
sXMVuFgt9Kp5CEFqWKWaWJeAOiu63C//eTjb49YL74UzpxtfI7Dem7RAtmAFMQDiHwXkUYaVEwz7
wDRcJ+sPVqIvxjDxZplB28t9xsq5avVCuYm+sahwjMl898CiJD83upn3xTguOt3VSaBXVfXziYi9
zg6DhNM1whhe8BRKJo4uus5UcDXX5nu8JTWnsyZnhzvMESBOLoyNumcKtdibS5fB53onNhuT/GFQ
YMhI0V7AQ5umSA5GFD0jZBLdgHX4t3lAE3celoSegAtkCtAWVPdIxx1gzEmhBPnfQ4GRam88sAua
zApowHBU/ByD4WlKgYovrR2GxRN7+msJBjxaIyHvoZ1H2YhcJy89I43FDh55YIqj62+u2UoEc4WR
fZHfJEObzpL9o2O0I6bWYHsj68oTifi6DAwiA7c7L04Uk89n9ilcKi7U1SM1ZcYBHwiE2l0P/DW7
qZ2mvvtnMgjN32ViwK/LKj6s5FB1FIL9N7zmRpTxfps/2XhDp/JRukWu5hPY8OG8Aqs/CmTfnbYS
kBBcj+aQ6PZqtPWpYdNcdrqWo/RmR+GqHDTowTzP6+2Kvikbpso9HqpucIOQX1ARqkx25FfNag1Q
QWg4dqmJoafN+/L3EK6bfD54P306dGBcsX2o2zD53uwzWxdKUjFVwoe8ssQutZ69d8bI5/Qj7Sod
7o5MMVqV0Uy5sJe0/a4U1YwT4TVh52UBujD6fDELa/9q60k5rsnXMaqiuyp1KwRaljJP1ZJkyz7F
VKy0ESDpW5EHYM7tqjqerZokm0n53VexqBhCfiWrbVX6qQFOY50/sylxyfIuE1Qez6bafzGJAm/Q
5dtv7mM1RfezXhQVUq7BuDzpoSEiK89Y+4EZYhlhLC7zWyedH4m30yyw2rhjP3hGlvOBu3kwQhoX
vnRqAJBvu9iIiTi+rj5Rh5z2MZwZrcvFmtaXzwVq2AlKxGyGC5MO4Qof2js3C/8jwI2KM44hg/kt
oz6FHk5Dv4Vd1inoAg5+JVeVSB14JcNb+1dC4EIRg7MjecxbCiZbJk9i5terMeV5P7yXaj3b1v+Z
OZOiXlcY7ml0ZhiwFExPLSB49KEuU4OxqE+bAZVGsvtOjnXQgOkiS9tzAGX3uFc74YJ/Whr6tjzj
cH/KQeLEHC+y86FVuufhkPGNhwcA5gNGZmmpLlBfuyNwz0jEecgIPukfMI/ylxbMo2t28rr2stAD
DetVoSKbgILtxuW4wk0kaQJnG3mEZDcWOi9IR5aDYXc7q4D8ZkHirDVB4eHes1xxWY+3FVISbfp4
nblMc5PHH6c4bBmV5P/WT3sHbBswqqpwwAlWDmxbyE9eObxDNIi46jdxXysoTZa4BCt1Uqs5Icvr
PIWLtTtfoEYPkYwBntVwV7+B7Gy4IvuI1H0N+zgf1zLcez+a4iZnQLREu7vxK0+l+8AdlA5Mu0u6
uuzCP7Vsx72/KYhDvxp9LktPHvYNwTDxSb07fdHvkp9udPFH68Xd/DjuGjgTXE/TklV4//p6kIqX
ysOGLXBUwBA02d8BhrI5FOGlzZthJu0DmHJaQwlSz2seThoYItFSPrhH+EgoV44G1veeCSx8GYCt
hAUxc8VTtdhIXMNjU532YB9UURufjVPOzQbN1b/PfqhEV6JawJfOWfHLcx0W5b16KpXzyAIICTyX
pAdpaIzzOJXcWxU7hAWkoEWrOnCtk/qugyQSYMjF7D50oTVrBJB4XXeTlE1pmHdvozsXh7bA7lv8
bxwqTY6ZWfzth7Ty53TiSyFml1KLXpRVxV93Qa7RPgoVYJKABZUSMlFv1OW2u5KRj9PMxOkHmDEF
YbC+e9rRtRClCbUSDN5YG4BxNSLY6TyCs/74frRtt6KHFdnlkicK/i51cKMVIaR96RSc4SuvDaQ6
x3HkuCVaHyDTr8wu6xqXNMnItvLihSOkPuL08HsZbJ9OiTMzrP+C54yAZsjdMEyYYer79BuGHGrZ
rmH0j9p7LKUgZWCXSHZqefeOyZ/p/97Em6is7LClyTjo51lnrEVuqiXQ47wE16y37L9iGYTM47Xk
/weyPXwtYG2crM1TFmmLjMDPPdFw7ylTMVQ0SdVhH5jkyVauW8EajbroyziGtLGDWjxL6tMG182Q
ZhLllxmo/oSzBIapdP01rfHJN+lahaZEli1w5bLL7JuTmKkgz2GZKN5b6n551RslIQu0O6+6OeJB
3tTdWFfw3zQ+0cOnovHFRIZOzExO3AuppGaprI9FxwROtV+2BytdVzUEHmvVnbF8m2UVRvpVVTXU
4rPIPRXa/RT0W6jEg4p6fIlz1DgsIqWRgb1U7WkTQmSgq78SDyzanS71ln//pTDroHnJGiqiY8HL
6pPRtl0kXU2Upjm6wdFHBcfU9p/9tvalCCTgn00ItvobPrBtizV6BzMid06w8WNnubDxNmPUtFhu
YzVrv7jz58jQz447eQqvZ7mxZfzZDeGNEQnaY7b72lDKrOTBGLEREPfUNiL27NOZzqEm6Gi1gkcL
UK3AoDfISR9iFfZId0NwaUIEjwdqavjhOSRyy7VYEwl4Amx8UxWjqIJZ5ahAMmYlQ9/JKd5mhV/t
Yxn9FVrZ9cz5QQu2jJJu34PbPbLNtsR4EGoqL/pb5V29QkAAzXDdkSQV6sfWRiVD6sbG8o2zAkm6
KdxObDsaeQQGBNBAXewiTLhVd+hQTsiGsDdTqelGLJdrDeTr7FV/BRZ8Yk1AzGGXLJGWMU4H5Ayf
CCXEyyLeyXnM72TYC+ITdbacbGf5FlAChAfBPt4b+aPG4hwB7WT37jpWm1Qr2/wblRNaudYIfl4z
1EvjlojA4HX1o7kZdJUk0ooe87NALSOxI1h8YJAXT3B5pjU+jOLcOncgJgxDfg5tDCO7V82UpN/l
hIqla1InmVXmhXXdwovSeQg8mTe+fMAytaaWeRneXnENCt9YTDgl8YQL6twv5y9W820Ah0E1xqdW
WzPlq6+xA/HWKfSONPCOhOMUHZCTuBHHEeyEWYbLDFOsCHujXXrpFsXWQVOWNv0wViwDogz50hgd
3nEpAi/43dxZUx5eGD/VrY2Ovx+AU5qsMUU4Jeig843kfUuv92WIR9xBssoXD/Z7HOoLyZcerZh0
nQyyBbshPrratNqs31G1vi54Lp35k2/BQbUvGqV3LGXXYargr6bcqU8V4FmHDtEEXul4pPh8PF09
1g3u0qpj1eX1fndX7BDnsyRa5HcNlUdg09tIPv9+WyqT0HXyHTQaKbZbS2NTq2hABihT1UkJU7so
EUVFxQYUYMS5UkycLnMJMCcP8JzlXio13C/2EDM6HG8OTxCKsV/4X5pa41K+0spdHAQJ2QGhmf97
3dIefL6QK9+BfgLgQpy/p2khN52DlMorJPAfqeViJsyTxqaH/ksgrMhgQ0fYzvhCwY05qrG/1pBa
SN2KfOse5JBwZvrta5PCshAnoDXVQYNFUqcTluOZizh0LdGktvmWDN0spziZBDJ+2TsgLO8QWG33
8qcdcyfVosSlkCgmZR/lTFp4Z/D0dbF8sujLuvax1jFD0rx8A7+BEqyTN9oIwUQCOxcFgJSmpOBa
9WKc46v4x1xdkrjrlr2mNVdkKZ6XsauCATDVr/X30oLOqRRu6a61jYv38wrxHwTRVzCjvU6G4Vae
QzMDWunDNO5HrXYzJBvo/6UDQPEZ6SuH4Lllh0JUSu3q55FTprR8rsCq8SucVF1Z6XvoagBS4k/L
cfvAwPNTqTTz2Q457jsWeWlyCGVRHHH5XKKNzFhjY13zLXAh0i3d5K/mA5VDiejlaRQwsFOaDG0x
auTDjVArpLN0oc/ooqbhB5R0wxCmkhLMnMfNXpEVRAcl4F7GFnkr6A0ghSWeIcfQBV4dCwRf+VKK
+4mgvSmGsVPFCu/PevMdz91wNLU0L3SSLyxc+3BeT9X4U1NPzJIvb1qIUQ72aHfj9AezjplWsQCZ
P/u3nd/f/lcA3UHGFttRi3S0clQ5mxaOAUuGd/c9fZjR2HWfWR1S6NmIYsbE0L9W6aYC7ZUtRUKg
k3gowRaZU8CfGtDcrVZjN7TldDX58O6HnBz/mi15wl6GLT/P0THVt2Zd81F/d9+NgizlFo9tYqN+
ObrXdPumvDaR0tGGGFy4MGOPZslcM5ykn0OpZEE8pPwIVfuVbK0hQy/CYqqTstwvSVCPAlMC7OeF
wRmcteVhvxzJyHC0UE3NBIorVPbpmvS4zMSaozKExqn26Urk9Lf0ogWp8D1mgBDVFx58OrFpkpQp
bXRk48DzirtCvg5v/fEmV/qMJmmKpD2N4whq+OHHVLD/NqAUvWolcTA0N0TUojYVvNLMCc0nqJ7q
oQ6Dkx/Hl1X7/ssaR7HaZf02pzeEy9erjS9ZaHePLaUfSeYXVwCvn694sjm4VAFdFSwxr00oQnpU
NHrnLzpqbv1WVgTmFvV4h3W0vucoN1GWnR9AeXdV7Y/Hxd/TuQtgzP1nHKy974TJzi6siQR/1lcL
liq0jV/NaK2YZydJNHAfTSN26W5TqvC6SjqWAx00KLJu9FTwaYE0flCB7tM3NAUCXnKS3mspwVTd
UL8GHWyjA6CF47/uTnchSvArvNg8iLD9H7K/ALSPGyQaFZ6J+kZT93xzfTdFtnztQChBOvhYzkgx
wPzk90rGkww36fq+Q23IZuCmUOjyMV1uzTDWakGnwZ4VqvV8JVkQS0VpOlFtFOfydpQRgV/A0BlG
odHl849tW93lt7+vq+x6b1cCgGqsUGOYoGEpGTHvgDv3n5yAPaSlYIkBR61WHrSLhjz3qadU0pDW
pTPT5LSIKkE8Y0QEPfh9KPIEf4FyjUi/Unkpa+OykdFQhtCzV0rScFhT/uiroT1sTCGDfoB7kiZ1
Uy+nglBwY1EcfvPTiW7hNYsBaDKtggVegTvU9+qOiIFtnujwbSeKFNsCCzykuF9m7Vt7rNkK6hGC
lqVp+2bBYwv9fwTwCWgcAsvr2gL9J8KR5036wyrgQbjUvebBXShjfRDIch/1qv7AjsDLnKBBR9BJ
uoXVNUJ8GuCd3jeqCM4ofMumCVk+4uYjTY3FJU6X5mIAsmUuN+vmFTFbeYWekxYUIkbUTt8RbJz3
1/nJrDDAQN3YScliuyMjXiYFD36HPfjyBcg7fqF4nrXwknux9c2ryhqLn1C4zmGMESRnOiTCqZjt
FV1YjKEcsLYkV9d3P0hnsjpvGYTr/Z21h2NZOnemiegt2I9LQx8axjUbblMHGYo8vaXTLi5BY9zW
uT1lVFFjO7Jdns8oYG+FgXdNEHEdsgS5cSAvV3ieQGsdRNqpJVe3QQeusVWSxGtdSomsowK2upFU
WTwwXU59hLoCrXvA7ytYYjgrXolOxjJRewBoIKyQuJZz9a1VpdAd7zTyZ5SUmwrbxPX9NXtGzoS7
3bjuKJ6b1T54UQ59MWybjTyyQuvKCwQFkKbcwcSwzBqiK33xce3EUJpYuPddax9D+ooZURlQINFT
H+LwDyXPOkGzbwJh3la1Wrggsq/MYCgjhMSpElanShiOaO+R7cX1pXDOdQDbbwqEePdtM/NmaIPq
ZrroUwEgJPuug+PQsRPRQWn2avw8FKYaI20EKf5gSpz422qEA8yIHP7ORxVKA7O5cO+g59IkGYzA
FqjZMoeR9Vn8IBpwzLcNwqT+do4jxXHCGrkXvx+XAkrHWf9hIaKKk/w5DfUTmFe6oGxqY9sszykl
SFjXUHyl9hnZv2C0n/n2ry1W/zsGA+KTTR5YO4hKZ0sOg6ahuo3s17sBes4L8WMAvvUIQccBnQnH
VJIh3zPOrGbVHDdWui2nFpM3dLCerWyS6Z7/7GOiJg/AsnVZN1nmtLbuP7jPzGeHW7p+PnlNujhM
dLuEqmqrDtprlTC6PH1V0CAci28fXrkgwP+im/EAlI8WllZIkIlsKj6Ge5k2duascXqCkyZKzpnT
vg043EYGWsouy2LgRKEZcAXpDzXTDCshOvmZUd76xbOvqvwth1Ff7VGoJnNUMOMRwWhftD1Y3Mrp
DIT3dlRsw8+9kn7/qwZoi0qh9RUX/wCH+TPcww2rWHPR2Trln5W+6e0GP+sjTIJZt66C+65quRt1
bgJqSji2qwjM6lckiuVXWzEkdUjbCQ7AlBXIrUlmpEq6xfnG3l49uZ649JH2Q3Yp9R8cjhF96A+P
QI1DBglaidpufHwJYM2zGkCBN8JxMRCeoLqRzKPdNhCRStdYk/44J7Qx3BDdKH8dvLICM1wZBRJk
LdF863HOtQ25Fu0KY3/uMNvI4FTs4jO5aPuwWKea5YskoMxxSjxa8RF6CHj7oFQvmR0qj6Ob8FSD
ayEvs02H+LW/jNxni8pdejY2vOM10ZwbsIKr+hMKVb5tKE7tkfSfstUOfS1DkbYkNjb++cm2ssYl
QnAMR/Iktq6/riOqFBgGCV7JBdDtzGiH0x9oGYROSbXJiSUvPXCdss8Mo1K/qPq9vmloEBIC8Ddi
BZDC+Xjm5cusJK7wYOT60VFK05lMqNDu/pI7ft2Jl1XYZ3S3hCGF2DtXDqv6f3q/pyjFy8EvtUIA
vccQNr+eCFl1ZBcG77j2Jq0vj+c90Y4W4Mu0cmbroo3bPutjLXqT/yrjmW89Rj632jx+FSQouJS8
O2p/PD+pOV+CgOggjn5Kks8RgbYkutnqdJQdIj5zUymqxupKcRqC03t/Jlnn9iJ3UJxsXUOIGQZw
uRy3c6zZqTpuvwxCj9F8y5kswZMK3p8cOcYUQCYmKAeIo1NOpsPCd53gSuzOEzZIa6IdXG2qNZxc
pv9uW7oDZEcaO9tZaENfnh/rNot8AxLdOKznE0Q+NhziQ/EtWFjTK7WQMrcMoNQn1588ALB1bih7
sqdZg1z4bZ1JCnm7hou+c+36dkqCQLDhDwYiUZiPLKJ5JMzSIMeZCQ8XuZvzx8TSxmWgZzBhyIZm
DTJwtBFBvj297uiL8uG32hzKtFGAEaXIdvV8CRN8saTx6tUYUJgFE/4OD3mA3LK9gElwzfMAiW8D
U5eCjAZtiK0z9ElqY5VM2lmmzG+xTYX+Bv/cLOyJwPRh0EtPv+H4KbpOwKQpQH2rvjT1cGjnoxE+
AX6SDDaXoJTx+KJj2i5mnxUwLanlwaM/za1q3WGV2u7eTO+hK0sKOKzZQA3QxfBNp/j+P/S4RrsG
ub/Kg7NQmgcFEFuZkmSHdSSoP0ABAcqjqcD4zHFQzD2C0e4i4sfbkKok96NxyDFx4uJFrtFqxEQB
cJBI569NOD82uC296jMJHLCat5lalPmzb2oH5X6+/iNLJAbDy4xj0SyIOEubzVgFfiKXe5xvOhj4
i3fYC494XhRzCoWV+Nnne1cGd8okn00X6UTxMfkWQaiferALEOqdwUWO/FzoKiRWOQ2rRruDcGUg
TuLeCNNVN/jOB6PYSkL5hN4A1jUotyB0fbUCF5FH8hmkfSlKK6m7xdJitxpQPZXMJScomdCbKxYU
kRVLZ5Iu9ediNC5CTFWFmeg22xnooErYd0cLKXEt289JTnPM4/f74ZSPxgtjVjI5xkk3HdB9UruM
6XlGPW96fbgmN4Rj7Tz3jLC+XRSAkDXEanN4E8G5B9rGa3YqziaoJEYM092Wc8XnW1NL0XBOIi4r
UGPT5aruVpYM/XIovEO6QA9ZbcEZYVE8Raq27coGR+snqFn7y4L3AB/ufSa+eyh+CJpbptGiMytF
HWdbsTJMiPduJtBqcyqhdjii0gpat2i8cTq0ms+MbE6SCI0rflII2KGagZkH5QkBd9BGRHoqWRGr
Ex3FkbDWcibw+OIcr74wjtBputmqzc8SzrdKbdJOWb/mVRb0CRdsDQqfMUHnLEtAYNsrQGCoAZUU
lV+7sR2tw3nGkLOvUhVQJ09tpSwOCnZgZrZ5/+i84QnabkkM0hZEfzFZiI+QETFsF94wJ0wh/7yt
kDOcP6BKjFf9YVKXK+1ASalHNiDWzn3BcvzQnN6AxFqFNyyH/wz4M1GeozGG6vjyOiPUJTSsTuAP
4nzTPdAOiA/N/xpc/W4LLoXHZvuJSX3BsEyUhZkIF9C9cHPC4DU1HmZ6jRBiBcYwLSWwTvCBDl42
bGZbbN2MqfT2mTme54NtEdC0RBRNm5YvQryEYEd34h/GubByZVwGVxQS+YPX1gJxQrkLzCq8ySTh
r2ooqknj9+wUGw+Kd4l9mmkHCgt35fuepTa4kr0+DuBWi7VvGdFVGM3d4UaGfxR6D0ZLAVz3ufdG
cX2YakGwZM4pnH/vwSjNxDMkA9kkJYTLIzReZcOxrG1eaBl+I6PGr1N1nrpG0CvQq/tcljALYdd5
FsZWEX/hxP1HXGg5e4dkHHn4TpTWNI2wYChuVQJUU3qIPNMV8mxzEJAf3yIwkHDGKWEmJmMqY7Cq
gXdlO9gQwrgmrM+mUWBtl5OKNRaPgNgfCl4TJKcFcTnWZHlJdSPfUimg7BMI91gVBcz1D46tO7Tk
hCaQrzocMNMOtGinOZBOYqPIcsLW99Mi8rXNpU7c6BxyX/ZNMsc21DDrrKUGTt7IKF671Ar9yMLP
viL1L1Uy7C97txebF+Rf0vR3DMLrgk1+dshnjQNpU858oIh4OXYIz/pTnXTTGwyr/+dBA2z+DObF
Onowprw3HOecc05OVlcwYThKJSgBo+x6ICp2CWyi1mB93cTagAf8PyDDWZmb8j/5THeYdbv6a2Uk
wr37CKnKJ0IPJsNAdEUXWRSXuK1B0acd5K61afvkwl/LaUTSWOazOjEhzkBDImuop8AY5ebLDtwz
3vbILKDrrYzJxmvBmvl4AEmDuQnCg+P+3AVcDkCkoXXNL6iX6fm3vLyaulfySBdvtRhspiJGGA8/
e8rzFwVzCRlVHIBvfx5GFEnfYFVuxZEzFjAe+Y4QoVohAIWrlpu17M2kyYiGQBcc5R1WzSAnB9QV
61vIxdQ9quWdkYDhu7X+f9gWy/gYM+uap3OUQD1EfyST5z5VgyaFfsD3klE98eTFJbtIndLiRokF
TTgsHnIMI0lNsCzw9rQ/tUf/DhgfZSGipifZ35WFVWz0sO8zvLp4u41o/Y/Ja0FiwfzhilvJ6s77
4xvJVltMTfLIPvgPpz3nNoSIBZ5gknWAzz1ANeka6v3Ogy1JH8j2ZmsyuSuBKrNIrmM2VtS979PD
OcQlYv+X21mZarz8T2YvdBIWgosQSB05/U2MUd+/9iAf6N49oCk+IZz0iL5YAdvR3jArm55HC5gs
RJUu2H6v/qKKFYwFejMEY5uAkO753zCKX3lNBylGlJglAdhYnRj9qY0avN19AbNsLbKhs9mm/+wx
1l7PWfnxYVRnjGKLU4S7H/Iwl/7hcLGWnK6PYw+WbxiWRQxsagsLmWD2AqrNBfLKUtysCQowpFxa
QJ/XlqAA94uTNIj1I8lJpis4M3kXTyqXOoLHdGcu1SQ9oYW4Tbqwzd/79kB26diezrxy/a5p0pbz
iA0b3iqKcx7LoVQdk0Hg4Vko5dta5+DK69I22GDXM2QlIDXFffktepgdOHgSHaG666RhoTU6qMyy
YbkEF1foii4yhs9eUFzvUyiAjpa0VHAE5WsfMwi7uzNQcjdRao6AvYK3wW16gL0tlLb7uh3bH8iW
r9L5myUHTtkEC//S2pq+swvVwz9oyOnTAc5lzLs9V0hD9YPKUI7+3gaYU4mZE4hNDI+H0eoFIOmR
Lbpg0phkZF8zXcfrz+NYzpjG9/WwdZvRsMh71jwoJ3vvwMaDCU3Kii7S6GN40VmfcLNhgPdH3oP9
sqJCPK05XG8tj3Jcy6xKJLzsP2px9hkeM16NWjMDJAVI0avwb14HBcO8KhKBxdOcJn8t/LWMZ2TM
+HfzpvFtrUn6XkYVqTCI+AiXvTOgxwXWtGVKpfuY5yqXPCY6P2OIU8ZPnAoU+dvy41udWXQ8oFMg
xKCjhVmqfFU1/fxSKI0GvZsuuQC4KTEZmD1YmvE2hrkR2DDS14SsF/qN5zOyGCJRq3uEz0WvgmQT
V2GrsdXwxP4Z++6mPC2MHvQMqTBhH/G0UFHZR7SgblyATfWFvToQ2G4Wh2VheAfePDLqK/kcxvmi
Zwkkl/4utst99U/FCgxn3DzWUmlCCFm3AwIv0b5dpnjbgf3lLi1A3coRtmkYw2lXkeLTaeKX3j5/
olcyQmC70G8hOBYZMPy9K+CnR0qoDO21jJxG+r1Vk44brQRtcpCc3pC98cxr+K6rloSEFFX0hIn9
k/tO9A/JHZaImTpKQoLNFHY8RDMzzeNqhuGDqORiV1XtDBtCTvgYk9cT3gpTjTu9X9soPGFTVc15
cjYyaqNbuplWpaue3EglwkKu+rzoIpTcoPA2/kwUYUIWb5xzScHqvKlZ1We5RTc08BgC8m2hh2EO
NgjGZlTuI2KIwkz6PxuAspAh9vLU2H7Be8gsgo8X8dd/jkkLjoZlEw+Q5wGg2Wf4C2RGFuiI4YZi
sxaBDZ+UKTHjBtFHhPdU+tqbKryts4gFtEOFQP9YchOUNITSCBPMO3Snb3buAOmcT7qE4Cf4Up8c
Auzs4BnQ6Cw9Kx8FSCyz1stxBguhiK07t03THa0xp2Rwdu/JUp1lPReJkkxLEUswrXjkhMJRVCAs
bCPrl/q2zaX34pXrrcjjFlwrgJQaFSKDi43dGQ00hCg0AkXJUrHLNiTA/xgU6Ng2nTVxlmnoULAM
mOX629RkTWQ5Hhiaj4PVl/ZcWRel1juJrU2YYy8DBFytod1mQoW261MmAz5QWxQw9r2e1614GNF6
pmaVlOSv8KdLbnzPC3rJmEomHu1lgDzN8o1Cs/FjJOJW6bqWV2uiogYxyFrnxpp2ctybyKHOgZV1
eQXQYT11iR52KyMfS4fYH6l9nnRAFuyyUSf8LurrxS8FxTNCQcAFYQENToXuKJH6tAse0RQqeoJD
Wxc4Idblj4F3r9liNFntW4/X8iinW2JFqNMs7s/PZRnlnR1MVsrYYLs1I4MKaf0oy5+yR5RBB9vq
I24tAYC4F/5/SSOkwkfLba7qYMXqPAxMuokaNLMWT5j7GPZhTlhb2JbqoBO7zMY4kiyfIuWC2ORY
G9gZEf/Hf0MZYgde+lCo1wQaViN/4wtTBWB06I50/anh/R3WGCoKN4Cg8MOgeh2JOG7dw29ALHwX
IZIiVtaov/Yt3IMOT5Zcw2RnMBOU+w96Qvq85ZKLA9za2Q66SHFIkcx8Hhx03VN1cvixBbykIwX/
ZlONa1rQ/cWR/hKszWivduC0WMgMjSE9OyzYgUF2i+kec91zLEm4EZ9/h5FOTVMIJ1vqrAyWfURv
Ytesg7z0qTQO/eBzxDb22fkW3VKyB9aFLAMh3EO6bkV5mlkwaCYJNGRjABchMn2+HlTZMz1krRL4
xEXyEOyIjvaJD2GcvNb/KAES1Y13xY45jINt7AHmRDbGV9zGW+Oi8rEky1xzt0XkSHHmmHgh5nSs
wqptu6oiUO+xJCJ8MdE4tSvBoYP6eaeg23/soAFtPMocfG/IDKaouoHnbqrODWcvtHCoCffIkMh3
mTDezQ5YTNGEMQ15scC9xgc00KzbTJbhBjUAy5cRNugneUR5gVHmfKJ4UKearZsyKyiBOU67RrYK
pApeo4W7U4xc74VpetW/A3L9vqlgGinWiAdhzaQTcbJlAmzLmpvrNIzG7miHy6LBHGKTLnAegr/Z
RWdWA1zbXhBZE37jJGgHt8yfLWNdfFw/aUBF6XJY1GXwyLJTVThJ4kSmxdgGvRj/eAhcAaUZCG+L
OSHL2574C/77H71c+Ysm4uLiiADvMUV5MFqNjdxY+xeR1Jno1573LiUKICxSJ+BgTZQrxS6kwXzD
6/YvxgFLS7mttet0LfP520YOVQargH6CJyuRD2WZEA9CrAwNga5pHnk+9yVLZhUM4uyNT7bIOQuv
Fv6krEuztlqXNhINYC2CMDKDMdrACfA/FaaBEMczJOB+9fL6dQukkFlhjyjkitalCqv9rDt30uIH
nzVKmd0ZDGBUJ2T1ivOTabcfafdcCKxTJyMs9GwdHwRe/hEFZIs6Lj11QyEWhkEolvdF22cBmzPR
7WwGQjjjA/rXF8KYmXJYho4nlFcBMfSTcWNMYmwWlMcGyIeah2E5S25z6lwvguKp5/zngNGU+gON
tjuZU1b+WJq5W9+nTzEhPMcKHQbmIT3fjOgDI62FqoAdbDz/etvmcTJfeZPq7Lpijrpqc0JBc2xT
CffPNFbILd4pCFHXi8oPPxdLhoGaNb7XBmiCuK1/FvA6TCUaGQgNBJazAM4TopqBBwf/0v83NgRV
E2PzZXbMYqVBZqcGax0hk82y4Fd8GAYsCZ29KUd0o8aCmVrXQSwDviiiy+81FRBTTiyzZv9pjLVo
XdPmoH5SZoU5QYx+ID34rSW1Kgx4I4chGW19PFGuwHiegr9pAKN9vC88lWy+9ekVs5go7jr8s7Hv
zwgOVjjyb4gNm3Be3xM/7Lbm7IVOURtU4f67Ms2AfO3TCFuc12sQLuhNnWYtOLEa65qd4p0V8464
7KjyuVENa2SjRcY/Ni+0mVmw9i90IZE70bqgLvOLGBFNcxKmoCQt1l01epdRzSmlMEnTBNT+bGcz
5X6eq6JjwdIv2W1PKLqKUk3LjDhZ4UiwkvSMMAWb72p9zwJ1gTLtREH8U8Y0+MeRqKY5BpIT9pH7
/B40tlY8RCY4fpeGhkubfBYpI2QxHkYQr79Stj9XCf256AWwKsqGuuClHXqkD6IPhMJMMFU1ug7u
0dzZ1G4OiIYD3aBG9TqanKnHHG2RFf8oJHgIN86DSMThPWNTFZT/CIdUFZIWul3u2cwyG8xGHutj
0izPcoCzOadJxBboSRhKtQGhz+wKwJEYJP8xD5KoaJFceTa2WasYrQeftLzpYFAheRnQnZawuk7q
m7YGA2vg/oT9LSJnas9gB591/86jaWTtL3DUvg4LoODgDdnWNfikpTohGlBbUAX7EmqO4yN7yhAq
DMOpAo3u97mn6bg0+ixNHXWPa1p7WQHPlfizYnC/fKvg06K93f+tY8Wd1kzDJcHXkEWOCsKuqhvE
6PPwDPltWjI+Ga9JjcWH1jF7JRREw9Z1Y3qXIbMXRfd6fRL4Wpk6QELkFZ2OolsqxEHJcFoDAQ1m
BKmd1Zp4CdlZn6qEvplMGcOu2SQCF+lAwiFqkCHRuDJOeEdztn2NxX2qabDqcnP2eDKxneB4wj/S
2cDpfOBhiBg3Tl3RPSXat0PBPJAf9xwZC4c0O7Q2Sh1H8ub2CG8yDQpW3VnKSNIlx4Ao8LWVD8RK
rdHYbILRw5lzTL379phQYKBCJ9vz+y+2whRlgVb3LPdaWFnjol3wvnn5UcpTZi50EvshXenm2Ly4
f3Q+nV/q6dESVR8uZ5KtB6/fyug3R3YZ3w5y3wzEzeFZ/pabhJ8sj/lQwiMNKuAY4J+OfprbvBqp
IVYRgg6r76MCkkJEBhhHqIP4kcWgvroE0gZ8rbxftfeABqo4qRq+pYZ1UJUDtz++1QQIehpVrsh6
VeiaomtKAFLAfagfiN0HLCeMIdgmQwmNvpllqlehrmPXN5keiQLiKINkPmrE60sDLJllltBPMGfp
Op8ebWqZwn9RpgyH6yKjR6eWPhAOFZxo+j6KV+Umzvf8FWH2q3TzVgoBgoMgREuGQYIn3+azAIBF
MT19110napl+jghnnZ7IABdLB43TdZetPX3KmOGAHPvkGAfw1E71ha7QTejxLSR7EyS7ALBP5R3N
BLfOekpc2dkhd0lWvUiQgNk+PFhTnKQl/KOn2jYyjsqcXEjSEirf4LlhQ3a9+LZFvkTTPzCeqcqi
UqbkNRDbZfqDp9C9gLS/VsEum4CbtqeTxZOntsMxApzn+Cac5jUEWfQIso/3yQPxK2wUKYZHtG3u
cYpCg0V756kcuEEmD3eAYi9sEJaauQ7xpSQiRpx6CZ3VjyQmcnWopbaLHWnGtcOoQ7Il7MgiNeQV
O8585Zf5Hwyjv0cvOSV3QGpXWOIalWJbcfFrhMcDWctJ4uHwEs4nB6E/ToWP9ghsDzhy0zizDZCs
8w/VQnLGQ4Djx4EkYFQOPUZ3mLtpPDjY9AZgCBhUj3g5MtiRoVdJbqGxuMEL4iYIfIzIDNhLSUxS
eI9RjwY58UN6HIFKeI2TkRIbpfprzvGePKBXfK+djMDw1e+c0qVLGFTSnY7z5NGa4dqLqG9M6P9t
sPwTHRr+7FptxBPmb2vMH5jBteK4K1RkM2YexlGGcWkKgh7LUzdg5D3OS365nLLqcmtxu6uZuij0
lNNd8eyP4vrN8WbRfRcEHWrCCfYTcD36aHDBhwyeSj9WgGtfz3tX1COTH7tmASE5S7eewXrSaeds
L2103r+31JUicS1MQw5EUsKqG7Xko8tcUI6guPLNKRd5DM3NJPrUSZjcKuWbtM2QLKksovJ6sNfX
84dvByGLcs79B6vq6KqKCaDcCA3b1HpOIvWwJgohhZingdq0TJPyJyPCBJkfhMooNIq3OPjPTHDM
XHdfNGuEdU2JiEiD48AstLW8k5FKWKRM0OneJ0T4Aw0CEmWW7hcYH0PEP0vUCgwv7r7U56szE3wV
1kzR9x36aG5GfxGZYlcFuDMcNn3EMVs/edZDpjMlrXeL/D2fThvgg/N+L/xwU7xNkmLLXGRpl1EF
e9VVg06bl8tZv4S7cjpvG/FJTctD0ejun8XvMuGw5CIIlkybf6hxG11ZJ8lYpCbXzziLj453cbIF
VhsExiRzejpODl2WR6WfI462Q55Qb8YjAnQMHM+vL/JqrOiKYxeilxqj9LUImMV+JZRi9+kuAWPG
pAbXA0iGhHdL6i9qbVsjUIBKnCswTHafjGL627d51lGe7oYjdjYahKP8hM/Z1K4WHRonTuM55VYn
hxLilZOklbCE7bAOCiC1oQ6OodFzr53o2B8RlZHgd5sMHkg0U6+rZG/lbzWuo8F3//avAnmNeOjA
JQJBHIsiI5tDHJiklGGE+ASajRrb89ypMgepSjp2fQMO/KyCFmg8mg2aAT4si5y7UYTJbWl/PXeZ
D37p67TMNTFvheo1FxVO5MbYiGQ1kd/V0rqHmu0PwGH9/pdd+K6hsNcHBtpQf6ePLMw2qbitb2Za
2nWp3Jv7wZAXlSKtgIuAhZIE2pOcO7YSkRXwhK6AdS8Jljo4Q/2EDDVFjVUn+2GzAakso+efzRHN
odBlG/X9HRW3s6QYagR3yngY/MqYCf196tULHN5GpAzIMR2Iz1cdf3uCH+o7qPf595Axzk203o/0
Vlu+gKAjpo/2o9Xu7GLa0VavC64gaxiKC5dO/4fuS/S87/UEosbaz7eGjRBeBsvb41mD0JAhx+fa
faBI+cD+cBsFp//r4Lqvcd5QDfGwx6TRJ3/MzxXII2tSTN2NdixzJnBZmB2W8W3Zsaw03Sxy/w8E
Z4VNbWrzSE/I+++YIjuYwoEyiN8Dqxei7tBo9XQ224wEWpRmYjbUKXipkEFdT0YHHU0nDah6/wBk
+L6dWvbyHR2tJhXY8Cpy+zS4f4mV0kv6eANAojoeGqYTrnOhys9Ilh267DGFblbfrt7ooCZVRC9t
PQOGQohkvxvIbuBETARMhFwYmhaHmSou9BJEztourSoV4qFE9KHQwCcNvKqUU6iUkw4JQx8wulUe
M5xPHrNmqK7C+ehViQQHJEikM7QdQOO3q+cI0ou/eiJqjB8AUCNaVjO9vGDhkPpGFq6/CphFa4IK
dJx1raWAilmuWkIL6fh2fgiJSykZNTdvU6Ew13m2G50hbO98u8UKAZTVHaLuwZrY20RQghHnz6Hy
h/MyXi2KbKnpoRFEqGmtm4AaytqJd9k5m7nMdIoh9h7QlPqFUUQIm6+DGlDxPo7VGYK01rl107Nf
E4npTeP/oVBP8D4ss8NteEqsHjeBrdDK2LsqvxpjHNTLqSr2hIcEYiMuNwVp2DIURIbcj7US4diy
FThfly/qXhnXkSHgRhob3oHrzSZJm3+fcgqAOuVX7LLZ4h5WcsdTfxcXjrf7M7uO6TLjKvmn+pPB
rF2VgN7aXp6pqUX4jHLH+rGv2kneC33TIAMI711bdu5/q5XcAeLYIxLI6uH/rNVW93gOnhdKN5Ov
VqGv7xmO/UaWAiRgiMDDRrsQWarcQvJQgQXZQJ90XGCQItUOTvEejql5xO5Ep05xkzDMyArDmFg2
iM0RQyJFIPwCeF4P6yuPXXX6gxQ9Q7coOfV7seaOH3m7C7gsgrizwlW0jv6sgTOIS4vEug2HmY6Z
ik/cylyzrhrFnZIwhGR9M+iMnSqNux6mDlzhOFuyJFzeSZWH67Cw8mftuyISoJaGsQ/RDxfDm8LG
Jo5vQiJosKDAOz7XxiEbWlFgIDQ+1yFBvx5jzkiitJtCzNOuRPEmVatGXJijlfkXyUqYS5af+vpX
hJ5rYr/2H5PXIRPW/Pi7FjbkCdKwLDhJ800usYVNeiNG4eSYYmIuNzv6WAN6jww3i2oqWPD5aFhW
KePsHc34AECIdYXdslt1t0dCvGo2fXhTTbMjuXcR+TxmRdiGc35CtJBDA+r/QdlI/HpA3zwnjtpe
4razqmVNsftY1BfiJnev5CuMTtAAFxO4Z7QCq2JuCzq/rWtgi/PFRkeEpWNSGaxO+iApMV7IFG88
8onQWhDANAnAl8+BvYiR8Wl0ilH75FkjNWqz06Qu9rWNIicMd9Bvz+QQiiTTr3z4WyIlvuLVh0OL
CrUkApn+4POdWT70Sek/g1Owub9vSAqdM+T619gJbDe4bqektQRrN1G6fNoUWh5UYtafFO152Ol3
KXjPQ9zTA4kxtSaCilbLbsybFvC3wRbC8Sad+g64BZN1EV5QQGqF2Fkcj2E4FKnGcLlO5lWzv8eg
tbexiPBAm4gLDqgfShpc6Qi12cJtR4K20o8L6mjjDitjrGYu5vIIE206J3qI7sbgmmUvQiUKnciV
J8nnnuYbxIbdbuDL03Y64fnrWivExvmGZCCpM/hJlHxWP5MAvFKKSW7EA2PPlI30vDTURPfDeuYt
YZQ8b7cSVk49E8V3KxhrqxmAW5rlAw3HuMoZwLbycI/yPgJlzoOoYR8Gk/WtO1g5aQ6j0ZwJmtuv
5N5wSiOLStvgPjIFSQzOhsbm+0GuTmv+8ZulstIXHm8SlgiWR/9CX4DCKud7y65K45DIj1nq//dY
0Kcx8FmEUrNXjN5/Z3OFqFArP1OejAOPwRXU41qxkYGyN+C7zrwAs7LiTIQfbSTJ3NXmfH/3sdl3
nVviUi/qjBfFnvr1KiprRhwIf01qN9N3TG3H5ubZPkI2se5SpZ1lLNrv/JH7wDXuR1TpvxLm63Nm
qjsBUsvXzl8r6lk8u4hds0lYaOHgTtniJVzJIZ3+p9rHDN6SMUGLTWZOkV85X6SGWRykMeHMTeO8
GgXnU5aqiYUCZ73MH02buifhocCTVDEdyN69FdaFY+dcyLsmYyYGJu2TNpTBvbQhwimMXPvcG+pD
jc9e5fiSoAzn9K6jbezSr8VBpxRowWs/MhtwMF5aQMCYbu3D1TKPHnu1+ejjOjSqVcKTK8fRinZ3
AdRzeKVLij2T5knL6P5gIKOJmfgqxSPFNWiWpVkAVoHuYAL/TSLOJaCSzvP7BQVq45qWM7EpkEnh
1bRXOA7j2mr93PfMyMBysantlnE3/8CKXj1PHKRm9cINKtoiKQTUGT1tJcHXmwYAW45p+lfs2MAU
RjkZD65O1KKTh6HEyQ27Y++VDSBWsvl4wg2dnrTAVaYENFxfVTI37Qent3N1hDX/u35tvNYCtBIK
4JMp4vxlA6T8WEf6Gjgh90yOFpQZVz10emTdgbY7uaPPGl8zCdkcANmuOsU0ahBNSrZn3ZrbCZbA
XA+BS3oh2bpuMkQkHOOmNiBLE4h7XhoB6tG7rl9iR0xQV5unOlehBUVgqHQyp2x/kgUfWRQcw/3+
5G9JTxJ2GNsmIFm1SbjWbhKuBcWhyhedo2vVIzI7TOeKXVd+g3x552771RARHuzs858DvySSnGwU
7LoYD0vYv0gR/0VmBPcQeIaKAdGmtB/ONWbG8x1fWaww8yvQG4JrXOW1EMEMhJxM6UhnFQFyfCxj
Fx46hsI0WzfOOgEYye7i3ELxUvnAD9w7s9aNz6+9HoA0QjP7aD76k7AHYNQS6u+xWoFZOQKdoGWY
8dS8O4YW1GNQ8tRPcXY2ebTdgO5Asu+w+HtKR53Zf68fMi3/+9Oa223U1pCZaNBsMx13QJolNANO
bEZu4zzXUDCCnAvM5BBIYc7dA/LS/nxSibRfUWyjAukULBUz+TOYukMLiTqcjuLSVXcLPHWp4cuu
KxPnEKvZzuav9av5yeE73kuqvVO/wuMJYqjkPuIz0aBdWa6jS6StHv5eb2VvpePGb5KU/LegRWb9
X56Evw0Ux5dxgP/QUoYRUcjPOXfxGEe0wC3n4WFkaotBNCfRhT4tppU/wuW745m2R3/ggLJy3bk6
X6GZpOUX7ZwB2pT5JKu/xTCsTrSva6GerxLB2Y6AZfroalJuw/Hrpy/WXVJTodrXFixi5AWu+zH8
7drUSq4CIXcV2Hjwerx+M0mWRmcGTP5qYEYhRKRZ+RJnHSCG8a/4C8GhHdfDhHV6EdtphisTcyMo
MgMhTKg9flIqtiHv8YYavNzjLmVVhD7eTMSIUp0m5VTEfKrdH3vfhETLsveZ6gfg/p3oh/CfMk8m
YcC38DWZBV2mNe5EeXa0cXUUJ3nj3DJ6zthYnWg1YgPeer30p0/zK6Iyfhv9nu1IOEr2nwD8dg44
vjDvx/GRRaUWw4g781lqatTXbbzpBq6iToox797Gw9H51Za2XvUO6KBzVXBbvF4ep4F8+MppEDCk
fDNXl4xqQr1/WZ+CrXx0nBH62stMuszvpXs6dVWkAPxnUVeAunG1c5jwqyi6QwW+uU1c6Np3yP9I
h+EcxkktD9Ej9hZg4e9k5dA4HSNG7I3Ht87pqkQp6m+5JBx/8rLy49NVQ0kWcpAUj5uKRblXsXCM
i437JNDpCJ4fkwa4ZdP5DFu0lyYzmydywWoVyne88a3FwhqPlmnLOV0VrPDF5xLhQpLVcI2DaHs5
tryM35pPpUIKt4d70TzHWoDnyGasd3uNcDB25Ux1Y3SoNbrSbEHFz4xfFKmJHh0ofB+90MqAKnEq
1gRQ639Ggi9KtpzAicoicpdKY4npz5sWivGKg3Y1CbuvpposCF3eLieS5N48DLxk5YQQ2Lp8nJbj
SSCfgOklNV5DDr1WpaJWkprDLDL/07l4q2hqcP7Lg3tlwnQwqtojHM3+Mh+jil0FxpvpzRSwB7ew
Mwi7Uldc1l3wS+0fCFYc/r7+96jCxPZaufSv1zgo2Po4eZVkneJQ2feL5R/9DAPxTqa7IrJcDZrL
kvTwN+dd2Gx2dFh+oCzCNSDcmIiuRIDmDsTQ9stcNTXNQvvxkazr+/4Xf9BJfYuz7jssMP1Vuwir
cahzksjPmiQX0FCSdQcZ6bXSy8Ue9/N5NJxLjLc/YL6tZqKqWQTedZQVDx/ECiB5UwnAvwDVXTpE
3xaqpN3Gqjh57QleTPpdRuvvHFDWE6AyUFBV9YiUqq6yq5AGjVuE560MsVVnmBmmLY4n7asP42r7
ZZG1nLGhrA60me4zLw+X2V9e+4WsP6CADE2tpc3/mFLvff9TK9AXJXOrm7JgJsxchuZ9ahPvOiZn
Kin4lfWT4NbW6E85eWdMb+uHsfgUDUw0+5VNj17hGVq6nJ0R5wClkY6bPt2nDUjJG1oEFVjfUzxz
shDuTc/xd6v73zVv/h9xh18Q2ZHXKArzhPUTZBgpTi5ZPNINUoMi3E1+K1PHo+zilIYDt8hK6PLj
dglZHMtm6iZF38z1YXn7oHASd6dhQDBOEtuB0Vzi7my4CuIsATiZ3tpc86i77wHg4haWbTIb+F71
f80USIpWqikWGdtnUBsg44avcJDk0yI3N7OZF8An8+qH8QjIRg6MUOFe4aDDxrRPzHMu+HmCSahF
4fWXEyaH2Tb8t6oAJJGDn5WL9y6AMDLirQJMB6BBxSxCuZoe4ewBtV6ynD4Hc9oW+q3tKZ/oeHGO
mgRUE8I0T2ekW/xHGXdBuC6reY2rhFwG0dcLn1OOjTmh4VqP/jfYerscaxFvEnzO9UXswLWVY4LB
BbsmvWX4uIXLwwMnbXlYa79ZC9j4825FBYRpFW4jfes0VesY7P3OdEuD3wcWRjiIxPcswFm3rpgV
oeQ3UxzrDeubx0wtWPXmP2eela6LjghJYrq8M4a/jLi6Ti0aD/JFFMj67Uf4KmtSQTcwBIkjZiAk
lUVuxy1J94RcLXFYbukb7ymcP6CWggb9F0B7bbgTm/NlcNAQbM5kOkoI52aqJFq9jjZl5a+hOL8n
sSDdYmfIdlIIXhuM0I+y0udXANCealol5S3Ditxeupfdc2eTrmTMaYXMAMbuNlACuxJv6ANY/Op0
FIPRFnS/zIuecolBQiHA70APdPaLpoEZMjFL3AmCiwy0mpe2oElie55FawPM0JZqk+o+qE9Ac+7u
JPgs0FTgA5iEwYZj2PzGIj0qxwx7cpJsawaEmeZodRuqr1rM2CfLE2GcHtz/HUs843d6x+8YjDvt
Qq68hwQ2zqKlEmJ6ifrBWDf5gCITtMcm+I0B16pmEGfUgg9de5hYeNLcNxOrVhjOCx2BxlPcxrZv
fa4P3as6wnFoXb6ZrcoP/eHXmbQEJ0fCoPhk+hUqOstgJR9uMdBH+itLYytvFH/6T87atc2+RHZe
dhHAC8pix0gBwNFki2RktjkBic848qjSZfedcoeYBWpn3LaG6bpWIIzpwJ6UK/GQkHLIqWC6DNmj
nriFRXdc4R+Dm00lFQ+FWCq6q4tTfJNUAVn2E5mR1eitbEJ9PyBBse2bBUFIBoN8nWJpIBGt8GRZ
GF9Tk4zZzIeo2laCr6Tubax2dLVMKfDImb44FCHTYWmO0xEJZIsgjo+JvuU5bspsFgJ6ddMpfH8y
Y1dt8SS/9zBwomlblpjGCHXB4cjecajC9z5+NQfSC4+TPzpQxSg1n34PbnjKqFLa8W7hFB8gizDZ
UFoxS33pmvFw/TGHh5imFV7WWr1nMgT0VSbKo1gBvlaTYbMyIgBbeVOfVT11h64WAzAz9n8jWLRZ
rdDhhu7X7n586E23oW0uSfqfB2uRmdr0As/zWP2fvxPPSExuD1uMtWZ5k131B383mA2st9qHWzey
ybs+inDbX1wb6y9hJAfZbhjA8NeCAFmkG4hmZ7nnI7R4HXJNMma4ck9uctstxBWYomY+C6WpKpvp
iAMmwVfcx2HSxMOqOcOGEmj0BRE/ZVnjZakJbz4UNladjz5BPOimBeH6dub7hB2QEYfy2PMsC5Ba
jBhkhmQspD8Uv3sZ6Eu+rqu/4fGQMm3qkfEoarjGQhTqUqsLEmu8uxeks/bTGLDxnmhcLPlQZulg
8cfSM2NM+WzXzEPOesovpCgxUchHfNCwUSXjtVEDzYBksGK8ULAGSz8/1fTufxtNRAz067s0o9F6
zfX4v6Qw2//RNCg109o0HE0IKoZ8q5EmPmlfVc1SsOlzJmF20T8IhtyUZBexuEkd/BjEjf+qk1oJ
chIHu0eFd4dVsz6AD4+CmWf4zGtcNIiP1QbEHrEKcX0eD57n7gC3cnhTyFETTFaiVtnYOhiD8u7C
CVtlAzbj3fJFSAQtqOWPDIMy3qSVp9KQq0nM0BO2OeR5NNepXI7B1vQeDJS+8LK4JAO3/tMgcpJs
bBbVQhc0RjgkGGIYMZuZ8akI/jKEwPzi+t6os2iC4QoHNaUr+iflfR7Pa/CJxwYOnAXFKwX8EaDo
qei8VCHs/DFgXy8MF6NFTfo3PXn47TJl0aEiLf+91NQ1xeq0jSMdp8fzft0Fxfbpycah9+XNwN04
SvfF2seurKTRnEPiRt9AruSuzH1TuyH07y+HbNzr64IGShXuwvtIy5t2NlY1qNMd4Lm+WLLMmckX
OsXBxfoYBpm3LaNHdTeRNyd6G70BgglUatBJaBjt+u0IqtClpQqo/1Fbp3ZvQ52WeZ7Xc2GLkHG0
Ca1XBKNoj3HYntqhX6A2lmclR/ou9ks8ZWynn3DjfZUbU1JwvWard6AYYJA+LXiu92evtY+32Cxv
sTuh3ngLkDpfZSEUYzbVCYnqQfB6PzUfOr+EORj74GJ2Pwgi5RMLP6AemC0/JUZdKOWwyS9X3lkc
EYB/EKHIeySC3a76ljec6sSEfPqhc8h8xXPhIw6wM76Z/sviPOKz90RxVfiOfTf9NKMkBYFxnbqG
t8oV9wk6doSMH9fpKKpKtVvgUi7OwoTj8mbL/Q0w2n5ByL5XEjxU71WflqxTX1Y4FxWXYw2BRPQG
ast9ANULNAngXe3NSs94nYcm1NaJcSyLXzTplVHMvGmPnpgKOMGTmaw/aLZPs1TUatZ1NoG7atPO
ro2hyfjOHSn2Eh7I+C6nvW4g4J0aq4vpMbozg8JAg5yQKTpU+s+W6bjazZH5J0ttPR+n73qKR8NQ
P3v2oM7y9FRAmS43TvwjYZHn0xC/FBj1qAr81yyVHVLza/tGT0FnDaHiC5MH5GBU344uur0RQLX4
MV2wb+jgenGwKnfxTGfoaHRjbkU9VYeHm534NRMcxU+qjeUba3xyxbN3n+Jn1IAxywdQejLkXiZZ
VkPO01sy6Ln/P6mBDhKfUZ5Lx3r3use3popST8WPKL15j6FOQAtCdrjVJ++Z8VQEhYnHT6ZW/8uh
pCUu9CIUxJvwN47yWl+uMAVkvO1/TVWz9GKT+cyL0i8twSYktVLAAX9QK8excuZ2HAaRgjg/Or0T
q3SqRBOs4VvetgmyGh3COPcGdcX1FgzIBRS22qjhCKtoPdWt02Heu23RkQUSJ8la0Q4TKyQQReTh
U8P+/O6cqnKrh0Wf/DQ9EiUfpEatJSUN/RQQCJOw1nX6ObHLou4LrIjNlEXvFwXCywv6UDYTTaa7
pjVmHQESIeBt1ioVjXDlASSJeIhxFbq2ZWdkntBlKE5yKqSrW97BibV0GgMsuqSn2ms12YbCi6Ys
fXXk8qSH+FiIv9rrHdqfIgUYeHb7lvg5NXh3sg9mnhStbRHXGFf1zROFM5/4Y/sMJkLAZRuhIY+7
m5qSTtvCZ1w2LU90gEjlmcLrjUlvQUe+SWW+2WkdJQxGJaN+eERAFXXljVDvT8qwkdeBezaMQdjq
JmfQCxvlw2HyJ48a7C6yN1Eol/zZSiOBLgqLK/tvp5NwrALRfJCcmqJq15y1T5AS4mpRg+JqrjHO
jtlu8GQDGZboUR/l440vutP//L+d8GLPlv3YoEGWs8cPF1ewhvKpUwHNARgWGGraCPnkn8w4n5Wd
0KaT1BR6N0PBNGI+RtKOxo8TxVziX3GobUiFAk0P582NChbSiXe8YhPkQtIizV5OXB8/Pw5mAIk1
Wihw8CGbVQas+tGBk+SvauPM5j2WUUTY8d4Lz9qBuZUSrUG8OZAGmUdxj7GyFNmkIgyVLdy+AW0L
By/B4ZCSNBjWP6NgFlYFUzL2strOYQDkoOBzwBLBn3o9ru4qe4I/UximS4HZ/Th6qFxmhlFp9OJl
e1OiCxtC/WufRwHiC8MDWOXJ4uRdzWnIinW4TpYE2OqpNTl38mHbcZteerctLCTIM6EA1d8ByDvT
nzaz02Anp3h6dY1DyTz/XvxoBPBOpyIpZzbA4W3FUzPwbBlDapt98Z+r90wpUFSipG/6ZT/tt0sQ
rZvNXzN7Uh3sjtIDa2LdjDVTu6gxZ+OWWo5R3l9OoTk1ZJ4gt//iaT0JDtdhiJQ8sVOTAQJZOnW0
v7sn1n62BqsfS04b9WtrBgHapsmAiTxhiy8Qdq8bmx1bdpbn/Gu6gWrCjwC3CPqbPC21NCfGvpdl
LFcOQXxWvPHXNPSdNLEb/UIj/JNDyN0jG8DCgs5awsVmY4EPUH3wvkBXAvXYFk2+0BLOtedJKSFQ
dvcTsqhqzpJIorxklKHQwBFNG7zlPuHbYPuQdlj8cBov7YFeuCgVdSoQtxI2knByKMQFE+Qrk6Nq
Q+H6R6IhPvFagAruWjWpHQPJWrbkTN+98Bk1sOQvXVCqOdXtFc5MXUb0nK5JDLTuc4OUBfgDpTR5
AucSJyI94nrDaAYw5tCB/7KjtCcJvLWeRmhI19H8yGy01ottnQc1ExSf/G1c++LZg8YEAKoAJlNu
OPPKdM18A1OgNqIxUr6JZSx4bfwihHiOIuvWDxR0GGq0JpJfLfE5r5TY6HDuhaV+PM+M05PYGSd7
CvXHbA7znoTn8zcbLT3GkH36Bo9eTkEjmYOBz2FQOAWdkBwlD8LvNW9ah774X2ajV3aRdWgBvFm9
GydI+8rPfoNy0QchAOVNhfLKOL6C+QQJpnd4A7v3pYzeXEKJusKowgezrnn2raspuUiwwDQWYw4a
JNyTX37FFd7TZi6IWRPSAztnpSAgixIJWt0tPmAkcWbtAXnAfHj8dPzrJclpTlUHbYrIcAAs/IQW
mK5Gmbke0wlsbKBTfBzPMwCzdjoU8n505F5VSX/DJZce5N+93pfYRUp5YBesYI3Zf2xKuOENGjPe
LkHtDZ/obgCxdufLAT+NQIfIA390/ShMTVWs9BoEJsx5TibY+T8/EOvd+hA+d6kJ/NxAKZhEYtKG
ubm5mJy4ILs/AvAZFQAVesGsw4rQqzPqMTRaAeooFqr8uFREMm5WcOA5eCu1RLqx5rJ/TIIspBdu
GoUxzY9IlJSPqscjs/T0PILksXuQMDPNvgJVJxkj/dQuDyOe/aiXZ6ydps4bcf9vxPjTt3AF8KUb
wfhnfS/w+leUCJJlNZiV/qkwY6yFmIdOCDFspQBMBPnbv+fHPNLB8pM0VzuKWGMtEV+7WMa3wmGy
tLNyYr7eViL9UIjt8mOcbGRaQeoOSZ8jRSX3gt99pw7TEBi0lswyvPDe+60f/TwitZSPcw9yGWrr
ziUJhF2O/hKOsDuPzldthIPicHHFTBxA/zjemM69GoyrmlBBBHf1YQk4p/fMk+oqxatvERyf22po
jecSFGfFxnzaxamnD1lcKkSXAkj1R3adH/8tOKLFpp9i7wJxvVy6YF8v3l0Pf5xFryqGe4ykKbBj
p2FbWOaetioiMnFy2a7Xwiij0Fvc5sMC+sF209ylYPl08fti5vt5OZPEff/eQxox7vpe9p/8IIQ0
h1PUyzuYht+dzbHWteKoKGYT1m7GXAmAmixD6Xs4eilIt/g9mYVcS/hClhetgkmaUmCU3bRuUrMZ
Bx17SWaRhyB0cWzzuQ/9YDs5CPhstK9P06vrMUfzvxIC6Br4AzbDrHIjGvRjUEjJqWLTAn0XhwyM
i9O6ClDpNpxWgbk18klfda9RElXIqvTndeLR2NGeCMz/FrnBT7Q5+Ii1HTinr9sJ9yMRB64P2xrq
FQwCOMYm8eYVwgs0hniaiEvuMvSMGy2fSrXTN8hPr62QJZbqYlUB6exXJkqprWEl+4JGSum4RI8Q
Nh4+YxXTMjr84C9Y221D/iWRdMxdVyvzcmwV8N3ZQFym1og0CDu6pmNlH0sPmnS3Nj1H/B7ThWSh
1NchGOCB4bpKl0MLSuTwfFKprLIT8c/fUk1NA7UJ9M7+ULfTLuMbUnE6HEw4Srg2EjxgXCjqLCFK
0z08gVDWy1vPLFmjBDqXrJ0VBR/kYx+6USvuCiyCeOBSx0LQDdZLUF0r0B8k8bGzS6H926QBgu5j
cmKhWEzUP+B/FBjrCiY6aDwKcCgiECHFuMWfAwDokmzgRVob+5s4hnWlzEIPDsacwKuOKovOG0YE
vz+pMWDHDKs9Ym0KOr6by2P9YWKbbOlJ6QOuZTMHAbQOSZMSWrDSCgFVpH7SN5mCxaudujK6bzBV
yDmZYdGhmppeFBY1pYsEYId4VQ155tfdb2jHBWEbXyNuPpe7DPBvEyZxmu3C57qqbrfGQkfV8YQ7
amGUKR1FHNFB6vaAFRF282qsk/A6dxpDdBl/WFHdKXtBLVRcKDvl/EuD5aa9Rfc9AT7RTU9azMjd
eTgzjB8SM8dYtU8/WCYOnfvyalL1j9L7fH4CxdHvucI0AGJP88jdlrtN0TxpfMFf1MnxrBXuYNHb
EUHL0XX72Ha7HkCgydIwlN3luGT7haRcc+DuHLH+77dqUKJIYMoDBY2RbogxViWkV45Fp3LFSSxQ
n6SzmVaX5ugh8RZIGPr176qFzjng5EzBaf1aEkWcpTrNz5lJXoMauV3fIh9zLqH78jrS2KKqUJKB
rf87GLBqpyZ923lufIoOYECem40F+Gc0ACE4SnTYCdZZj43N7TNWEaPLInVb/AzPw9nvHcQAfNi4
Ue1btRB7fWTZ/wr3f2ija8p11rDyRXBomyvkWw0vpAKj1VQ9fLV9B1iKjWnbie9HwzP+r23qjQ/z
DL/xryvvZxzDaH2kvO1SbvYdC5mEUuuXQtao3swyoxDpck7vgBWC3gjD3lrFUSCfMMF3ZkZY+r7Z
a2/blo5C9Vcl1/EhLJeVVD/+gW87DU3DdpG4AlAkDcal/NXodjQM4BMryUnqtcs2ZPOqyx4GCNyG
UyPIregs8AZ7Rqh/F0j+dntOToiJ/cj5XK+tzJ+Vpbh2CzMlZZtJNZv6SJ/DAbT4UIo4I4GSHd1L
2b+hCY8rp74g9BgU4zKugqCxfavAbweCD/KzdmR2mHEoFBvtkVjOEHkSjqfYQCV6kEWJ/D7eY1+p
UGmB4nz6v+JA5xluT1VkNR3hEOKrTtwxt+Mjf2wZTVXtqs8fc+avBmPwl/fVUzsK47j1ufihbSuz
m/FFSmPY+nh3FEYa9N0/wy1muv3eAkIGiEvAvdW9FKGBiI6FL8xzMTl5RI9AsrK4tsVLVjk1EXNI
LCZSkNlzfMzDObB3RvKrLp534ienM96gqxV7riVPEr0ZXjgTyAR+x7/LTiyc5ArwNXYVPXLQjtqj
bKOZq0UYXvtVFBh1rejK9d8zMNvDxCsWsDeBSQSJCgkMDSOpAvdfY57ZgqSBF2db+Rrr6QZd0iW4
waQR196IN6+iNgBBQOAi9ioXl1mNQYb6rqzW7ahZQJI6fGG9Oi1z9gHGpOxLnlqYJIOpt1ltIpbT
36kx8Nci1wgsJBXyS4jPBDEbLd2kzzRtJSL/sJ4rhtoHxDmi4pZ7rTL8xmMhpnWuRjWtDpQTjtRo
G/qO8+mNq4JUC4ow+tnPxheobem0YnDMyGgjsFf1rkZ/kGjMM4tXCh7GTMj3nUnx5WaEPwGOsTdI
S/cVmK7F1DNSvgJT9WgUUXpfQwyTmKtZJY1/gnSxe8E7ZcPufbr7KjluVUFijZk9t7Rf+sp5SJZn
HYtwUxIndt16a363pHBTC7WdARbo8TI2jdP7X6O7NtJ8O4pa0tepKsw1Mz3TgSqZvOqchvWAdPEk
wX9d89aQci2PFXd40ydsh6OUD8fFOtTEwaZzfj9jno7ODiMt0NIyKjhsYd58uRo5am7ApPVNlkg1
rsUK2bvIad47hhLULYfcszpaZAbjMLV5obxT/YmDeLHCoG64uTXOwgI1TmqlRWfUbVyP8cVfreH2
NX/ADOKPDID8AEE7V3nvLaJ3NIHi18REiGFcoxqE3b0mVntcRUSnL8wY9xyMlUUtzXRCPJdM/VMq
9WdVF5us7Cj47VXgPADGLW9/OWGv7f3ef2fGWuQMz1QJoks2rUmjU7x3OefjyhPNbXacipB6O13K
SGGHrPn+45RC2gQbgcBhphY0nXqoyL3yo1WmX85TMYCltgah4aJJJ74egeU1Jrt1ukmRjdgTEMvL
7NO3tvOLsP3qhZoH/YtxgiNTnXrBifK60r+bLOCOAo/l/0BB/Qh/0sCKfG0Obm/gue/eJM/JXqk0
cteTjviohADjpQ4KwbIQLFtxRv9OPMZnuylsAYk9CQdAbyP+RUstcK2QZNVaeXSYKR1xCkyHHsbl
fgu70g215UFG6nw4pHvE6lZPp7E0SQ388XRLQmYcEASh8aHpxXlIrRzMu0gpd/EnsjnPGBk2mTuJ
h4iSoYfww1n6FmHoYeVntcDdA10XjNL+BTu2XBLqhhSwCzpJF+87u8GA0pa2SYiWxXtJWu0mOOCL
PpNiUKOajTQhTEwRHmBIBSjn7UKNkHWU8tkmQD2iJKm5lW1Wj8HD+XK2fArwIDU37KFp+tX3hgL6
rgK3tQ/WeHLOHqnqlimHBmSzUpq/tIXhheGBxZwt27AvtoPOfplJMUEKetFR98IIYk9y6fzEGu4A
wd8SCmOimvwJQxL74AH2ZIBrbKXE3BfA7CuzFXLAxkXk0NiVhKGnKE3/1yfY7eJkDdbZauash01x
2QVYbgPlxmP/i+CL8ffiIMQdcbNNryEzCkxSH/9/0VUOyE2axajoTJozZfJO3HFanitJQUB+nPpH
INjC14a8oFzLl0Eoey5cd+x4MvQCLyZ5RVhBozLNn3HBxXZhxC1Gqmw6bzpikTWbC198kViUnF6I
hLsbtKzaWLdDB79DtrUFikW9qVog3Zyd8kDNuVAHCcUvOkvOAyc9+6x/NMqte1d1FHXblbZMSc4R
OvzbOdbAA3PF26Ly8/BZwpn/coOcSaRvDfWSZkAE86H0nLf58pPPdn3bmIY0ZZREWPmzmNw+o/Tq
UqLU6+g9yidBxzBXdsqVzCd2chmkEbamq54Y6+F9PKyU2LD7nx6DfiYYMEDQ05y3LeiJvjbRlZtA
9OYJ5rKoIPeAbtvqauP/ib092El1WH8CRbYJhUukO2Ho1Y9Diq8ASgDVbtcDhimKte+eIMey2knw
QCF+cGbJeb3k/8+hA/XA3yCS2c6kIwBkaRjqfaSVScwfBkQ5zLJGaVwFazjLIaTQQjA26shtgoIk
j8n8QOAqKkg2pjmDEhtgnHch6rwzcjq5SPQQ5B6qCs4xw2lTilwrC1rmBJb+0w7HdtyYxXANxLSk
N4j5AIzn8Q2BPpmr3SD0AdPMz4sBI43i1T5CbUp48W69qefwzLd98168q4ltbHHlehui1BqnoPyU
plFEa2EsiHF+7UU5gOVU1LpBkx7pM8GYp19886jGELO24URhJc4Ax0+1RqndIhDWiEC5CL8hayBJ
t3L13zKsgjO/keMxaiJL+l1T4Q3bQ/ba2V1+eTuMFYlMbdb2uZVGhR13xYR+UftXhrA3oEcuK2xO
+59KjpJgVsuNQp7NNuuN8mCQYUjZCrli49In+kb2egjne88hWKhN7/D2yXyretba9mH5d6hbsB3H
GnLSa1Ts/kIPcg3F2snF2/dDGdJYKLS0gfHFGnK36fE3mu7sF0lN53RP9FOyCvb74vRB5bGcNVr9
Rwj1yrq/EApu10Ny+XDKOTI+BaFfHut5qx0TYVYYsRb/AFcW4XtnCVF9MjEz09q2XjHBOjEylQiF
g0LLFRDzNTpvjjlx1rmCsNx6xUSOI96PgaU8Qft6QJzf14nyk/9OH/a4S1iQICj6euJJumSm50Fo
pajTBYvFqQLGcKyr+9pz8Pwr2Omy+nSz+T4tXLB4dVkXJCTR9h9d+p/JyVVonjGCHGf6G2BGOM23
RQsWf/5fO6IcLsAPDk7iKGbiTfbO9BIP0k7hg00jk9dQqSarJNpqGcOCbwKnrVDrbZB3cRy0GjgC
NUiVysL6AY6FzMpECKNgtS1V8PtGl2/7u9/I8GWqLg7a43CSV2D1LfSxzLYr6L5/om21iw5fjW/W
fGaAeSX/f6ESwG3eHiBf0iez1KTBTwQKaPGDu0+i/euCxwWnkjwCfxsvyI85/0CYglWqVTMfKwbB
KjSGcSmihgFhAzJ0aor3C4mPGdOK1TOJVxphCFV/u7M5Gby9RFk7QFVcLoua2RF52z8oRhWQHNEf
uUJ21qZMBKOzy7y5M3ThyrPyXpF18An+1+5zBgp8u7l3/AWmb6GosSWSlOdaUQ1t2JlLnvbFx7p8
OmG1KxS+sAF6mRAJrklo/r3VpLFT8drox1+8Scgab9F6bHzfPNBJWfxsG4PxxqUeXYDlcWoDcC+e
GTSJtS2664KdGP5GXsyAxKN7kMiRGsdF5hP/lMmVRGA/G6lVwqVs6nYDEFycEcKaTzp0xMm4YAaK
VvdXhAzwpzbiZ3KoRW/RKugjoUfnBXyGSPWCRl+wfTsWvQDpff3oeW0zeaU6Dncf5N7hehC70M4U
0P4Otjhzt5yV1DVq9tC8DR5BC7vBEbo+J6Cf7DmItc6VrpxKJ/xmqFAgLAfXS4WVayJmmUSo5aAN
fKmu4kVZ64G8kcBnj1ZyP0cIAoD/3NE0jw9cyPvkqU6QTFTMFTXbD5Cd0wTqxeryLWx7UfovEK1D
GlufS6VJ3j0vGZ5Ylj0ruVNI8nY8yCvvGJdvq2g6xvBpekggt6QoDLs2i68WQCUMbvd556NfvN3M
dopFCkOOF0FckfQk94xf6Zo0FGYb19bYBUYGfaF9KGlCg6dDlEQFNwb9Yl+w4NMU4ow0hXgav71N
Wszqf4Pnp/UD8j5DM4lU2YCwIOa4XPJH5Fu6Fw/Jn+dNXkY4hXpVc0v1i3KSmxe8TgmCbpWRmZRM
X8l2hxoxaoUGnhBl9yH8cexMP0T3lU+cjYnNOtL3oG7wkBOFU6agGAOuztZWj6tHaWfZN+08YUs4
y6JnidNgRaDFYBPJjhm8de/UUbFh1xZw16myoFO/2/sdz07DXTYeJu6Ph+dLhFd0Jw4HAqmb5/fc
YZTIdWpI+ec4QdS0MFJkK7+76r2AnkYSLSMckqiwHsFy1cE2ELrnrOLukgX1sKZtbtR8vw2nZSg/
jzDx4F7eCFnGMX4FwVzOghILihPMA/fY0GILbz0fL1VSEv+FBZBF6hs+MineA+riNyzlK/Moxl6v
VgcYVU/sZej1a2FPVHWIm3rhnRndjL68Um61s3FmpeU1OohHxRrVejAACZtHw2lVQaZuQvVugO49
ZG/x8400lY6fPeomACdGxqYMIHl+Pj4q0FUCaUhUArX7I92W1M+toI6huRST/pbgQbqtwNRKiZkR
Tx58o5Iz2bh9x36phstFIdVG6kjbYT3KGTaJ6GSDkFTQfM+755Qw+I++9jvrxj0SFUQ7gEoXeFGN
tItvCuxG34Gu8BX45/Sn2OqCReYjjSeg/ICaBIFTCnJJSn/RUGwSE+mfYWcmczsx7XZDvAaVSwzZ
Dka+wgo56Ego3CBmJ3lR1TObMmj652ujMpXtIa1+u5fHWJwWBHWczKZru88Soa8PIsiY8syAr0hl
almu714PYvjeesTHAjTVz3z/UUR4Ny5fF5mtHpCHWpEFWU0SqFvWq5gesmzy1yuXKYd6id+wTJSM
FiljVN9qcp8cYy5yJXP+sslF4qvAID0SYG9i+Y5V2XLxHaN5zrNmAbvifvMiCdtZvldT5UZScLiV
gCYU03bc+fQtWIWQ0dwE6V5cDF8Og1oDH2oSluiDE9KNpZlP5dd/832w0fILLuM/2aHrJFvv4Df0
hgEQNKqvCsuk4w3XVoNwlyIoKLpk0LefJW8gpDmQKHLyh5TBVTUesmaQ5Fp1O5E9wlSvIGA9u+TF
+doftSbGvUiTzKbzYVQD9FBtI70Qjy9ZepKLq5MTD1Q0stsPctK+PbU0dbAYiLBWg5x2JeAlb/bE
zhJe02e9quj467sdmKlzru8oV4emctOJQaPhuB2CClwKRETT9Nc/VmhOc0YNm7zEozTQbRHnGLoF
sXW/zWbSlX/Nd7OgxAw5GPsaUJ94T8MQe6N2qV0a1bRPfJdoXUKLAmbD3jbBlr1um8w/IxCJWL/h
ZVRHZuh/GbX+Intf0LGw7/AFtaF4GtNDapIKV59cN43NMAlEI0vKlYMz4U2EHfgvM6gZ9HRoOA9z
gwzOSC2JVwfAOPhXaybXLftpYG35SbBF7ozVepGMMyqR63yqgSHTmJ89Q9n0XUvxaAggJfT8Vfrj
WT2fz7iFyx+p/uHy4PE6RUH41ywOsW0u/ENsAuG9Clv5zkMUrLG5BmzNmZnPs0ECYgNwRIuFPHeN
9kgd9jdR0r0qKlguFhfBIQ7KeZ9rc6dBYdYQhUvPMKIVwK4j6Fvppwo5BfEyZ2v4h2P+kvqlkhMC
JF2n6VUhuO95GUkbs/V1c50Ecqt4b0ILyZgghFauvVb4m8Bn1gnZBKfP2IN8ahtCqufIFlgq0Rsg
a1h9+TopkD6rU8rtxs2wQ9hhUU4o9j/g7l+f66u0t4o7qBFRXII2+tXjo9zwgbz2VYNoRnrozHr2
qlADe33g6UNYQ2pVlRLfSqr9RVymkEu+TXFqMsO1Caxug8JdFQDj54y+IStH/Ilc9aIpLhYfTk/Z
M2el0x1EZX5epfDH6jKHReZ2jHwrA0WXL3p4FW9fnSLy97zCwdE4UiltydSUoMEUXXWecbgsi7sa
rOW6prdujHJzN9UfE1ngNwwXgwwrsFM876/d9/6Adj/vJZPJYl7EiXwDVUS8BZD/KS8svFSZDj58
iFxYPAKOJicHQXz+YQjh+S7OPgONqQYEnT1SOIKIve9+kFYbgz0w2qfyHfOVdwFX3jWkuXD37Maa
3RFpQS6syZuAIxHddSsNlzzNGy2eq11lR23pEe7e7Jufag6gDDFYIrI45z93YQfA1wDyTzVI4Xni
CQ/RjGqJFQODNg2g1sR5VuBewbOK6/Qz1L6kd3OZftaXX2EW8b/SXq3RLb+jKBgEycCQhcqO7E8Q
4XJyU6l9PyfHnDp5JC9ekrDpVFZ+C1O5KwwKCljt+uV7W4guyc1Uz8a0TjHQ6rnnMw/K3ghtWXf6
37yf1aamVDebG0djHqkB27UMug3PjqQsGC5T1McAjXGKcY+KuGwFfK9ZQPJBDJ35YNtEyL6vMbMt
tDfbJBTJFzRapmkUMKL930wk4wFVUx3GMPXYi9iBe8VN1CGsng3owWHMjq4zt4A5fOO+33W+KLgu
D91qpiq3CJmGfOhW+z5xxGXv1UYQ4Fh+xgEGllZg6ftrNhkjzO2OexQr6M5e8H5XyXP6dynWrq7T
ckMCGQDybrGa08mQcbXdSGsrXQeR7sJPfWFWlOySmhG6dTF5gL4WzGxKzw43tvKDq2MWXK5fO7f9
l8EBfDvkObGDTztY97iXx6osj1g+RVRWZaWBw/pYl7TfsTUyyHrVvSHYFE9ySEfR/8Su2dsQA+h1
BKe6OjoBRnJ8LDMcQxFKboWc8TMFdWSOxWi/za3ka073cRYBK0vCR/jQq8USclAwMilLFpB0GlGf
JIgBZrceQYNh7as5i0MbdxJHGImWFtODboEJ9q139ZIRSdOT1/sxcgRAJL25M/NxoX4wY/xUBayS
+cwcqrWMqgftySRRq9TuoMoLtTlMEZizEGCVxD/FxyFzYmDJ9nFshqKlz20BuZYtX/nMJ0OiUbCR
+gVOshSMT1Yy8d1FyK03UQ9mas24BAEdPEeX6b/cNsoSUh3Nt4lsE9VR4NkM9/hHRhDoyIGzuv6c
QYicap9vE4X0TxQmH+WcsWIj1iSZgkrX+Hl1WytfgSKpWg5OKUlG1W04Rb9xHIK0BhuOHvLMnRj7
Sa6VjwApg8TCD43WvPCBrN4hdephc0iZvE6ktOgbvtEwi9/N8jMbczwWxh2YF0xuUXU/uotGjS1l
/ynNdz8t7Bk6MIIR0+yRVmm343s6pH+Ij8CFVQfyrrLuErTA+/rGNb2NupKin80VSf9GAY44F+kR
axyU9Lt3IxF5ch9eEnrePbrT5NIvii2k8fVUZh1gH6ImO9S5egiWWSNFUnrVvAHiwbwd6zA7Pi7a
joS79Dlwe1FPjQgm3s+aETcElBU/iFkM0WQ/wnumIN7r7WHUIbyd1VV5AVtHf5wjdG7i5kjxXC/1
YXaxMAQ6lbWnbG1XHgdBIrV1VuQRugxm9ZntxyCK77ofdSfAvlhQYVVsiiOo8HalXg+a8lvDyJ3f
cnIiUwR8in88jkKqQSRYTM1IF/mXBsIJM17apZDLYxwVHEzhMic9wDG1FknUTbLqU7kqp7Ke0uDN
KoFJijl9am7qMT2UGiKsPF3EEZ/DPshi38PfM7bR0LMoSukS9OI5M1i1k/UBTNsfofFX55VLGrMN
NQIT0XoBwxQkN9ttPPFbDXp5FBZ+E1LVolXhwq9Ii5hxfCr4BoTWXU0ZEgkEOP1lc4/1LKV3ajcm
5G3p8jmYMxcWUbfkZPmfk7PfR6x3+hwTw6ZshgpwZhZ5udMd4x1V6NIXJetffix5LcGn3fQRcAnB
HGPpw4lF5ELVLaE+lYnTom+qz8WqLhVpW2mgPQ9E9xciEaMEV5BvZqDkPzsjgB1tjzH/Ef6Y2bAd
Xan7QWBce2lHIK6hCbp1zsxIStp0o19VBbBn0O3zlMLvkNsJpRCHmqMMDX2rTU4rUkg0w/mYKc6h
75G4HRQpN631k8mv34xYhw35Qsk9sNEs41mvIAVWYDNzashYmXmVmSFIhqL8HTWS/t0gtqSHLTyk
UsyxLzqUPuIEWodmRfqD9nSTJHg5XyDX2lnxiH+4c5dbQZiYqczYRNQ49DkEuZ3tnmaGk6tueaLR
cs5tcrpAYV1EEBgtNpVcikWLTI67bzuUbTTRZO8XKP3QZ1gqkUmC6zs2dLClWyYr2N8CoA3f9qwm
kZnp/wA6Usp91jAqR0AM7nW05HuUL9pytEOvtRkMIkEUHxTfx9W4wSLvl1RZCdeEolabJWmIIUos
uNpAfVl1OHs8VElFMfNS0hyLRZsK0+mtkywNXYEjbOSaymorSxmmj1QhcoHzakBNLBRmCiIFjixK
dKKs27FvbDWu/bww2UXhmrNPtV0eizLRY+u8bo0eFFhVOEAtTB98hE1KymrcKwx4b6appCCiGZtw
T8c3OQIqCEqfMD/e7Pm9hbcChQOL2aqodlpoXuoelfxyuZkwXU4uBeEr2xyPejFMXm9y+iEGNg+D
q8uqp90wjVDeJAQ8fy9kvos31L9jmhT6OYxKQIHusvy6dqEUnA8QWq4xQCB+lxInutc9pKw7WM2E
WPoWDktx7zMaBLxNZ4r/N2dimXDVmszrhM4i/aPxDWC3Og0LBrC4CAmcDt1uEsndNQmE443sWJ5r
FA6dagCmOfudfcCDcYgvoOYmyOr3ZOiDTzaqc2OacJ+RHclQHjc8siNm9renwtULtYHV/iTgo5cr
6JzM7FQ2kHX/KyCfDIsXiRbKZWW75ixA9NlwQhurS31wbN1iw+G6M6s36PAYtSucI9X7Ygv9qysk
TpxoXb5jvjGfdEAowUEevjFMiUE0+g5M8RXIg4CfZ5dNCJrIMydDS79KG4TvCiIWVB/86mG6ys+K
BoFkH2EwCkmDP7EuRUSRtSXiLKab/ducjv9sAG1CYEpHiw4knZj6qW0KTq4Y1q2kK2x1KK6M/3fO
ZDGVB1TxuL3YV44d0wJrz0pnVt5Xob3C2BzUHQw+F4wtqJf4H21af07mAZ4dEtxIAg8cvw3Mds8+
sPcXvUkSaCE8avD7Orr0pBb6vIt8I4wBOZzNBO+DW3LliOaG+3/dS739K5zwzqyzud7QnLCrO2fR
96+2Ol5CbJG3owhrHdI045+MM6lDTCDJh2YCEnMM0QCErV9SbyffnHhqwbT503jAlPdXHFMZMlR3
jgrlMsOEoicpO2UMOzFGvjVh/l57m0JKCHCIXTNHZArekt0MZnrNQY8RVoxtPfLLEKk9ndt5rdkm
JCH74JcgMjch9mQ9ZX5Pep0tJnTEk01Q+1DynnGpdZ52Y19jEktzPf2tlEmb4CS4fH6FJCEjKMo1
czQSEXDSy4V1YpcvcmhMcbrRhn0KVdNimklV308DrVVttfY/6p8U5Jnint3DFX2t7qEpgP9eKC7e
F1aotTuc54Xs0SmviOAX7iWdTsCEAZPIEwbVJT3IB/9bykA84x1Rdjl00KuFkm3jF47BiCUOiMBG
7/Yqo950wy0Jef+WwB3k+c50HYuSUQAUf9Z0aG3MonxhD4WhwIe5fozyp5zNeiYJOWQ56pKATGlt
8+TErA39JvppAkXJHvActZlYymT/qtqyXMF0af7ca0ZbNLLrePmEYvrPPp/8e8G7d75pH4g8HFqn
mD1IxQ1ruf9cPb87JwOdV3DbO0WPFiXQVfv8tzrPNqrvt/UFURdQVUUBdg+9PqkqFjPt9yIcb7lC
2KM258yXWM33PB0qwLQlZjqWaHdEByWqnlR7iiUTwBrcinWh23qxttEun+f5uu1/JyrogXOUcM2A
Q1PCcBBX9E10cFjXDGStx4KPPKEpc+5FD3+a6D3AW/zBu/Reu+V6tDZFBzwYEoZ8NNjJTl0hVF9C
lxtho2VIOY1cWTtRnRv/3ErN/3sqAQ7QRJuE5FSTpcMV7q4NXi0Gna1+FizoSWWhP/QiEWKv+WU0
2vf1CXuIONp4NvGzBncMo9Xg9WoI1qEGTmN/Np4mgAV1siBUlb16xWUpkzeUcrEUi1YHZ3+/nySN
B60fzxtQXNYKp5oX+SEwoEtvOOZYuzacvWlQDfGtCLbxE6uEbZAB0p0OhmcGsDWzrokEyfjVDQu4
VKl5Dv7nboiJqlXpksYhrfvCZKNe6pvy5DSoYqaSYNobL9ba+UjSWnN9PZlfcgPh7Bsnf59EM9qB
gNfJy8OUKrLiJs+bd3UUo0xAtFyOvSQAjUJTn6BJLMKsxd2+WRs9dUjs5htHywhG1rkNvecZY+Mf
WRwrXt3aQB0omVnOCfd5Kyk6lB6IeuSqt+iet64PmBYug7hk2iI8V4yvxom6B4RwTJ4MIJc6ayAt
IQrNo2NddNLW81XMrke5r5ZQF6cBNX18QjrkxtHDeuPy/Cnnq1Fol+si0OH6YTw0h6NyI55iWVk6
3b8REZRgE5Re26uaw01zTPQHL/pE836L3IPISw3gxGK0PYmHxRisa5DW1jTXSqXGEcbfSyGdXHgr
X/olLzjj9rhueArLOqIMafM+P4Ipr+dgnLWGsX7OSEKOlMnmAyAbGiGlbUb57c4H/DkKKSFK5AvQ
ObZi8IM2mrRq4G8UumKWbh/2JaCQgquqDD4JbVwd+l+zHWkq9MP+EmnJVk3hj36NNccsmXVqtu++
xeY8rbpE5PLKL1ZUtNaWhWZzxtULvQO4yx9kuq2/LcZjh1lodxGx0yjZGvqZY8VY20iU1l8U1Pxk
jC07oT1uDWn2X/UCDt8t4QWVvJa0dL+oPk4SDya6o0pToTn0QLF8FylXgkfvHHKzJTxGRkG1TDFv
Xettvrj0MwmIoi0aBbuG7GkeWUrHwEFY75t0P2MAWmgpOszxtJlaR8QFlukmh8jr+xv6Ot+y4B1/
82KhX8V17/uJuACjBMHkphqGzAMi+EtWDxR26munuksHBPm7h8UgW/KgWF/wFOAMyTrXbMopMSn1
2/fsIjz7IqedW+lIh2BuKLFKizW/6VrngQZyVJGbzvsXlSevSKJq0NGV1Du3+2pJTgWPoS+dT9Hh
s+8sVE0juZVKO/DzyIhRgNnQCvB0yhORU9IIlt2uY1QNXTiOUjiJ8Aq4yzXisF9Q+fPPIez68s0C
hC4ityND/BiBsb2H66cNFhnoDQiA4AZO0hYpDXGd9CqsEks3Dc2j4+ju55/TCIIq7Uq5/j4bu4e1
315gy+y+rCPuTXNmePrEb4PSdVvVfkSwwJtx+prCSp4zx1zyDhaEvNIpm8XWVbS6cPOFtH8HLBqJ
rp1UcgeL047QoLjhxegqnzeRa3irRCMIFYLSu0GWRKlQpfa7AJpFCN4Pdo7GCUdle4byfj0Pt+k/
RviP96IeNJZjaMMc31g0xWq5HLpEueidlNFH8UCrW2wUGPr9x2kuBbeMZUKCAuldGVSDQ6ZI/tDv
qsY2U8WIXHp0/D5Q+tVY9QryGhpHWtteZi6KzMevbOT9/GoyWODF9Rl8/dmLIznS+2snbl2p1CzL
HaN7ff0hkfdiJhSUhI3klbdhsv9LbzFPvJoN1y8VGN+u2b6nIx6iyNufRJo0+0xM+stmpzMsGgXw
dezCMzFPbl2ZK4OqwdWV7ivX5TC5LoezrL4UecvBlFWwmOmwP9hzKQsBEGkeVzVVN6x5u866eLbH
wL6PQe393YxwlVPeOW2BKxdWf/qzuui0iEz/hts/LxQ40bPQDyVF1UM/NJ/OWxcO9iMbQ1/Mc1gf
jABSvEAMScncRbKw1Tp96dD3Om7Ujt2UWnDxPutq9SRnd/26Zg4UD6mXvQZzkwV+oVd/zTeuZ4uu
sSNqfJbkFBUmJXgk5slaw3H3cJc72Q4u0YtwfzXJfK7VpOqhfJSMrG1KdsaWT5paEfH/csBWEpNh
S9QpX9oz0hKyc7MXMB0nTR5qu2QapQCx6pLxHQmEhQ3N1kVjdiLptgRcARqObe++0uCU2rZYmOS/
1zQe5NSFK7DHg20Sa0Li2yY7S8QKwBbv9iIM46aXsavJfVg6/KhkF7W52ObZtiPhOG9Cq4lzq7l6
AhMJrVF42LR3Evt8IjNmEyXNrrYWgV50nxgxmyAwLxReT4TgdysXbc7+5nHNRjAQkL8VBK6Sz6CA
8den5OVWuQsZKi0A9g4rF5WROtU+Z+UOKBWdOKZguZQiCqasUYarZH3CwUevWeDrjnk6aEGeyUN/
hehKbR3SkuU5j1La2dBT3+CiYwcDvz2JIrWCGI+fR6MD27S2SbWpV1WkjtImQ1hBoKh7xjiIyVnB
zPNbaS9k9Qjm4KAR3m++EWZ3nGiezdiY5NiupE1dOpVFUQoJAQ3IL0p/FpBRTQiEzaLc+Nx+O8S1
b+vSOQlEjVIFbYl7CKeuEa8ooBtDOEXOT4pPwnLqb1nhclSzwUMHvwE+4yEcelM0FKUm1c0YNdjq
YbfXawIJm+3se1oqVHtD3LjIDo+rjmtdBGzlU+W50IV1iJtm4rkrrC225T4JuZSpxxBg0r9mQ78M
swAfZvJ9g+5gvMKJF0skb1kZFunUOvuZGb6uJOI39vO5ozyAhEdFoEv8XksYvvOXU/37HoC+kp0h
SuIpgtmJZne01Hw3AQXkSirN1j5JAAwjb6BzD0fv4odEEB9PRsj122NxtaGVnaZ65xEnDAlj6eb5
1pApbTkyc91lMvDOGwQJicXQ7Qa/oAc5C290qaMzEov0ryHTgLDd9RKQ/rjG/8rRoqetDo0Sa0Gr
BV2Hr6HeXPe9NhFmw08Li1dpEkKDpI3x1jZIY5ovO4hRx9SFljKt3u9+3CGFnkgiZcceUDx+JwJ1
NTAGFD4xMcLIE48wVG+x71lvWd1jEqYkj6rGLuoRaP/G6uGjro+rg/Q8Ay3viOMJUw+MVJQRgpaj
ovDenwHHh1yzX/AxxrP3OB8wT5U0G79lhRqxMLLh59XhQeX25JmCxXFA9KAKab4TM3z5Ja4Fty78
Q1+t263VbX8zFw5gt+R1fKCz93+UTdA5inKhJUMdUYr+q5VHzpyJ9YQcuZyNDPXkXIGdI6+IAcRn
L2Bz56udVkJLpxjQfRPgJGCIKYsp5bRIW3iKDZE7pYSUjXSTKRBNRk4MFh3b4F1oUUWtIUPoEPQq
qWvB6EbvEl2DmE+iCJFsex9zxU4kGSqdFUqU49V7y37T8Zecr1tVHwb5/Ciodg+JbIQl8OMWJM9M
tymwON2ap5GJwY09c2G328EVUz4rW+nWcTb/c7x4lNtMjMexNnvRCMaXgukk82C4eQ6PQmqGHznK
aR65BnHYQbMMv4QPQd82cWOz0BWlfrPgK5TWtv/L2H++a6xe+eR7ISoMcxXjY9Rxej/E3IDB6yyr
euirgfSDWt9KTtbw+PgzB0UphnFcDOeiV008tqTMKQ8edcGKOXOavStij0p58+EeH7AnRJDXlP2D
pJs2lejRejobb+CUr479gi51S4i5XlJAiWTijJuurlUlYDpQB76v0kjkaSyoLa4j5fwYLaBZBD4H
jNj/vLEHugvS1pUmr2+lSWIB1RVB9AFcW1IFkk9LrN+UijAtSvYSFQLTs90TnG6lZMaK4OE/I3py
MYRhrAWy0nVMuqr3ZB0AHxiLNu5t1qxnX1EvnUso91CVB+ophmZ2y3bDsXqpzlZVUxgjxmlQEQze
v7ajrI/ZdpcP7QOvi/O5EebS5kbuxrdFd3bhzks40+MDKzqu5qn5BK6b8ysyNj/gAxXCqUoiIpSX
7CC4MR72mZy+XgjwPTICSKsNoko+5s/XLAyqgF3Vavu190EdER2mTwZBPzox7a6TgSzomAUGU20H
oczwIgxxHRL2vjZHPkCNMnPcvDS0pP+UEYl56wSo+Wu640avUCJYhKsPZ4SAzbz3/scXSfla0Zvg
eo71poOBr2IzSKad4ebHrVoz76fxd+lTjp58fmztICnKhFRVlXJ8Rzv3QG1bM3bHLhslOOuotxDl
VLs0Vmcf+HK3NI9bOkNwBIxAseS6lf3dju5NNFBTsEqV/zTw/SB5BLfwOnPrhplkZzg7A/3lSLy/
P9wIj3JIlVIXkIirbrNrYWBKF/aVK5iRkIkXVEqNbfHmXsGOSBAgCsCC4zYIGtVHxQgYiBy7vDGX
uuKAEHylKnzp7cNyiFwr0oeUnU7mtCHSvqkuyvE3rME05pNRwxD/keTKYKQRbSZe71Z5H9MGy/f2
+60cm2mq7QmtuELJSWp+Soq7wU8k2zLf01wl0rWMuMJzOGwvvg+wOW6Diez10O+6qyTvzCdWSqyv
mckSIfozPk6TN3+VO1+uvccor0EcjMGvqvhylmfapdlkiNg7xxylS2DvKvYeFMHegHIAE1K2l6Zi
CqiwgBVeLMzLsUrnZYt8ka20xCXzuekxfQRoDK7GF75y5ElBxEDrgIyj/cmDFbtUfOo1UB4VmUOk
zjFG0PyYxNJUlgwevWJ6DUigOdatIidML0qfn4odvM+19pWwOq+ptceT0Ib3NCbjxKavR4spq7P8
BWO9i4/92bMS38lxGiynROy3DrxhaDtlIWvRbPoK4sBxKTWpKQmY1K2oZo4+nL6MGE3ArrObl+69
M9H2/NVFC0G3UfY9DRcudO4XV91wn2l3Nyokg0L5kZgSWEKbyRjpxm0l2XZl6Tkh4/HH2g6wPSSA
q9Pv4zo/x8czlsMrae9yHfXKtYhfp9L6eCKmBiAICW8AadlqsowhSDjvzmTbJIZh+kJp5n9Ti6KF
IX/yp7hu0aIQaB4WK3ShzgjKsSQZ18aEXJUuKlBU6ebSU3Q2tKOeFidYb7+/EvLQDlRluxdIAUWT
W3dceUvhCizTDIYLORjQi7j/BkVt6YgaTiQ/+sERTMMvy8B0VDrLbjxjr928rtk61Dn7v1iFO+Bp
0GXInVPeyOgptgv3FqYCXSWEuSq/s6uoCfcfsDwcei6eI3M4X6IxMMw8dWAhAOPtx/0v9Gj0RgfS
2yjHu2OTIDOUc+b1cgsHQv0kH242ow6U1x42vWbzLVAKxA/dFWePD96Zt+Tjdxfux3dWKdcxYJyq
YdH1M/g3njOb4I4Hsor+qtNn9YQXA0yXL1NbBcYQwseq4q1MVZh8sR0SicKcda5p6B6adzVaZPTB
nCNQdJIfuBel2TAIh5bixjZQATZFTa887NebYBVAx5ekexMwQOwrWqBBva+GpHTaLJEjgyIDcacy
abZSKfhICMI9NwbT9rMvpwvgreGgP4mGXCa5sFPDx1gOFiKvDOv//7PRtE6fj/igmt1ImCSRAZLq
UhavAK34FBvNgDiqOY/zmgK9jmdX0gT7OLSLh2XxnFB7+ChlVj1KovuXeD6R1JZlRK/r3siH4Fat
kCL4YzLGEkzv8a+Nq/2QkNSS08vB/1PZVuWw/OX8DC+XYyWYdYMc1ZF76TO4+UjLLAQ21kjCDG8o
+tgO0bE0y/zndD0O31CPmJLYQnMeBUaMIcqVBYRjiyNDDA+qYFj9X+YV+K5kciT9d1TE+ut6XzKN
0zbsFDiuuYVqWNy8PyGfLirQLoMSb4Qr1aF6wtAictSw5HplSDv82vb/i2VsAfi5duyyoryguZqk
ekSascjqFzMK36CwwnRBZrZlur8M2Htk9Gpws3CRqjY3c7Y3pGCFB6KQFd048YdB9xy9IyXkXxF4
Nyy9KQfBuFmM1vTfN7NcnoiRYid26Wj21EX0A4B4CVyjeyfDSAWVcgSmWphromAubbVo2oKWa/Oo
+v11d20Tm6CphcGGL/gUZ4AvcwhCoW8W1xkEHLK4xAkK82LN/JMP0b579QLPFYNsxy1HKvEp2yhE
VFwgxoXZLvhAB9e4wv/5ARWD9LMMRrH7nkGfTC+gHg2wygsq9h94Xl1i/+C7mlV27Fynn6f3IAGR
4Hug6QMEBwYI75jezTquE3NFOz80Rs9zQGpVSIaE4feRWTcCR1KqSZOqeswa6I9U9KLeT8rNZdcU
glx7M0AA6FJnJsIb+FcF+SuZhTaqw/oe3jfdsQ3sxzXIxcs1HX1JQgPsA1YkTQOQx5ErZXrykY/l
HbNzuB4NRSQsXLjsy2EmRrhktQCNghexmEEh8Rvo607SNDI1bBuZ1/izMEAhnKxUjXLmCra/gPA4
gfQztMCDix++H6CnH4FYq0ud7t8p/mrFtJ62J2cV8X5Ly+O+6vAKTihKrj8yI9HetE6DmKKhrh17
T1H5nFDtdaOhmQ3m+OOGcRmr9R/PhLL6LT691EgLORf//xUgAqRgcT90UpohS5nbT1TlvqRyNBEA
KhbTztRzwNT+a3FlCXNqcRO7pyGF8/tY4SWpqY1jruhb+htPNGL7ECLkFrqUzTe0c5Fu8hHE442D
hWc7dkLpoGkmbeS9rZQoGHUPUXgzz203tf9iWy4DvUYG/NThwpkh4NilC8dezkOEGN16E61vDNOU
EU8CvFnfPHQb16rYfrUUmGOUq6SCwdHxwexH0GkTTgMwZbVoO4RzC/VGZPh6rGUc1P2VGo9xO7ja
3FCifE7nHu7Uk6dBZZHZhwpY1gPv49Az5g7I0H4pTDgL/FC4RygSwYfO6Fs+iKB4ziuHk51Kz2yd
xUXbYcOG9Vzfy1HZg0ddho5n+kggDJywP4GgX/ayQKMAp0M+k6/9s2AZCz+Al5jFPgZMDIzGSjf0
tfZioImnicHmjH+uvQFuTqEEsGpT4Rm8H0TizlTga62vqCnWQjzZF6xU5mZH3d+fHTQzF5q8B+wE
HMVu4XMYxEUgrS88ZU8QWHHec/WzqrZWZux/mioduSQtY6sJKPd+ZKvNZdJjQn/N+bCv5j6i9rm7
KyBDXZ9W7g3MbRTA4Qw3QwL/9S3HUaaJdAOfwz1YIxHBktUPW8Es+bhZF3C2gJcF/37KfOcQNetG
/izD5xjAZXGTN4emA6R7C421+7sUszw8XfsxxT0hAmrFIt/oKNpecK3er6/7lTvAAAxrw9GkhUc7
KRZENawTxzT0JI/6UawWACG8A1tpHGIwOMBWplWaqRLljoS1AUNbpqxeQyxoTh9UppX1tbicWbG5
2IyEV4QKcokEcL7R8w2ZC6SeZv8jra6NXPKMaJBZXG9Ys0dc7NbX46v8k/W4132M8NlmXHcYpwl4
fsDMr7j5uqbptWNfeKgO/IjBUwkj9byUgEJiazQsnZiXRDKpTzWmhloMylqMEv4J27HHyRxyyM+j
54fqadw/fVWyiMIfO8opNNrBi3J+h3EWHdHBe6hav5oz5BnOoiABRLgV1Xwx6Qv5WAmerp7b5DVE
obT3n288HhuwMzbYn1u/gGJJ1ywNo+cIOeRVsScJ1eNppGB3YqzFCBEcPVjPRxFX6kZcNKWph0zZ
y4DRY9BXiXSmhX23mpZ9CJEskAhrTAKe4eApw6ywWOFuXpxG99ujZIm0cUZBsnSe0FuByNgMuQoC
r4wXPiiGHOAQNPbkWfdJIzFoHat7UWueRJYFDihQ6doJ5ttYeYrtI/zKcnuxedt6TFw9zbbfihor
RO3kOBEh1EBEjX8zjKfJAVycS8aJGCs3k24kKLSSwWJ3Gz/m8T2RV/Z9ufIYNk0AnhvlLaRtQhwL
AeoVH5KRlxcysKnwDJIEt+ndD2x2ymR3gI75UhLsihJtCeuE7BTniR/n+y9lKc9qm7Nx3bco0UWe
8XNGUn3s38csJMpQq9XkevSSR1Bc2u55sZ0/GaweNltMxQIaAl2I8pGr4ErQgwiYMY3xIDWUCSw0
QsjfN3TwQ2UC1VyKUdxJEXSb4YLLOGaiUPtdo29b9TUnfLwFNaxytUL1OGXHdYHRbKBXrSMeUu8Z
rUc1J+TYp66fzX46MlhZYlUgRw4WU3WJMgh7SpykyZhAcIaqsVRyOLMPI6smFHfp6tGic/iKiSW9
xOpEmUabeWPjr4+LIwxv1qLR5nkPde8ndswjTZ/Td1gWFwkFco+Fs7UuXhykyKG3VlewC4KBPGYL
b9YFPRCrbAcb9kORgm5ErsM49HVckGq5rcBixuD+Sz3IMQVm8ltt++ZG2bk8Z8Ff41Jl9Lzoq9WW
DXAO0zWRMBDq+x+yhKPsHLymQ9q42WT1cDhztc5H8ztsjq/mtZjYA9YK6X4Mp4urQDIEPv/6j+QI
FJ+3GlF6N8cwqNf9lWMamkTnhi7c3vYyi6d0Q6AT7Fm0Pk9N1trQsEExJrzYCjZ140Y13aY51yQ1
jmcP4MSdX9T1hQcBFWIbAXOjmOVku6BS2/Si89KMQqdbQYTboDJzsNx1SH1J5Snd04l+YEwBdz3H
WIkGed5qkxaiMbocnpDK23CyAB052KUoVQPzLh4hrwkIszDie+LMdKjbpff3RDm8+fJOIMc6u1PG
OErEkaMqUxqjSj8/3omNyaGxpi816hHzdNd0lgRvx0ie57q/hHhwFeVTtpjfGv7FtS2Kve/mPn3s
6Tt88Gd9njpOoJsWGNO8gbb84TKKQjQTz1gmMr+x7RfpOcQvxrS5rcl+gQMWRnd13zYrossM3U0m
T9MOgLQq4yM/51ZFv55kuQRv3b+qH3pP9Zo/UjowjvwJCMpetPjIkZ/rFIUAV1rtQCgeb+bXjI5j
yuz+AZJvhsCKXnF/xbM44D61JmLy2sz0vxRebjgSeTIfhkmMPO7ORUJVEMkzJ3jqS4Y/p8yqzb22
nLkOyjvYjBh5HQjYkTCbDcP8qg3Wigd/1e6nrjCDH6LMUt3yU9hefGq4XrnaRXdFNcFJe2bGH+9L
w9cAZfzPdXhWUPy5AzD/ujxewsN9LD+Y7ILJK/BqHSm7XiJ2epgtS4VFZj3gBEhM0Gbrj/mkWR3z
aYRBFJ0pJdwveswyoYnUnsNvTNa8W3fnh/88Jr5sbqhqboDfIp5ACcw5EoHZKHpYeceZ6LOfPBjF
T6B+tG+6NiF6Un/fxwT4kWy1jcnRHJa3i0Cgc74PeBlLJEd4vwa1nzsIb3gNCLG7y8kGOLfq+CWm
tjmVWXWFgntMjtOvbOidWBXNqMjAhExeXfkvH8fouE7EArzN99jsBw6MMWtgqXU9lbSHcFH86++x
9mL4Fm2AiiCcnAevMHNcAOpviK3lRoWJ9uMy8bmLiImqiGW9i1eBh4ixg2C8WpO0+x4VtOllMbj6
RgfSsBnJIPyjIyOUpJ87QbkYtu9Y3rYM0UKJIypCeUAdZeBZAQwhEDavAWeqlObs419pIhoJceTq
3lBQtSlZODgoCZI1uqk/MwI0hoFZIFhCLVyXaJnHvwDRHT5EkleYjemd5xgg3QVB7DOml2L2Zot1
Tzj0YMqyXuv0e7sak2lxA1UGzrBuhwDuW7eX7Ib0NJgbxG97s0MmmIWCbSVzeXoguJsw/wUACqJj
Oz0SOX3BgVa43m57XdEAYtz9RqqpUGvWVzZHSgvke4nV1wKhPFd28VWNCR0layKs7neXrvg2fHZO
+WnSMosEq0aPpsXh4qsSWNIFDrG0eWK9lzhyZPvPttQ7UGoBddyMxTW3pXrDoK/vjaT6snjEjfek
8CJWIEVFvs10FuEvX3ny0IWbY9p9g+VLinTmtRGcBDxM1OYcBYjxRjAviaailseprl8RKBmtzq0a
nh2oSBtOZEbJWkU2AoimPpJF4GBNWuSQGcg9cApnJ7Bh//OVMXwNUDBCs0IJKPsawGEIjX2W3ZjJ
kouxpHziam4NFd1ju7EQ0jFl9js3OL4YZhLkXbTPfjm5L0d7drHS5sqUfUZEdYKHD4X8y0ZiEplG
1hd8pO4me5dGOwzjrgzDZMsZKHvv9JXxVzUMAgGYRf/p6TkPwDCG1MtWp2LCb2VpZDrUwyozVYap
IPlz20fgOzyfXBKXV92D45ytx55VgEOVw0fi+CgtWefsTb/I0Zt0No4UB8scx4m/LwpEzZUXRPG2
6QSDtFZWMGRT18ZUvok8B6AmczbK4+tGmoI7NTElA5IoSUrVQ8NRdSfxiMyZorN6yZWeTdGUS6XU
OPZ9IJ5IHth/Rg2Fytio+ZmO2HzpDlJqfmKYfxPDwO3WiZ2VIDuDOq/0kbkm8+5Bkt2qOOxNE70n
ufCWI+tmy6K344D2Y51h8OtXfQtoj0WlcMTgpX7/Tc7mmu6tdgEnBU39yiQG+kHY0N0Q32yiuKyc
DCLxDSwSHk0g1a3D3hQt6K6K6WL0M+d4si1gfh6Kg+iKDpIeAkgToEiBIVDKunN68JHvt4NYdqjT
Ct7ZUOBUgtu8OKABoYOJpItzzykG1xOPxBuWtzBxLSvzbSPDMgLI+B0TQnRzbJ1mstSVPsaqeffr
ELH1083kUXnF+ygaayfnapfJSJV+yPsOiqBLLExS/xtZ2OuA2e3HeMFDV7Vcrtc/9G5ByhkF3kBq
YyqtF/DgTXLM9QCWCtLTGsFPq5Zh5k289Y/UJzBEtbZWwTlkzHsrg/r733eJ1VVNyWtjokA/385W
z9CkLAtwo2HmMPjHn7am2xyr5OJq4oxMk6imCScMEsJoZdSdtVdsOAa7zMNu3PoP5sjlCVkZ84+o
QXS8zwVCIVuddcslIehUmpzv1tgmazBQDoafRMhAPm/l71AOWrI6WfBXhyu5qotoAuYfFpzTb1Vd
s8g5Bw/Fd2+xN9+kWI3USy+4pDyMfsd2ulvLRKGhkpJU+Rl+/9XlsDa1PeQN2F1ZFHpZ/5YlsTww
ZD4k4z1fymlDAOCb0beQBY+ygEgEJ4wTyr6XqbI0paWct+bo6rGKftMypo7Qxkz2kHej4ekTD2Ew
vJQ1qaSC5mcor13NcdKQjMZrlkwtHVVFGsWkYBKwUtZaG1LoCig+4KPc6gtgs3yTbR0aRJHsv2bU
ttElqHL0YBT/AVsCENLxyoVs13Ieovrqu+ufamSebAkPjBaELz/X4BhnLQJtYe4CCJ4A43C/DbqL
CXcC8SSWGTi+VUkV4dpInBBmZFOD6/jTIrRyFuCNLqXYBRpcwp/Thy2bu3CCVnmfAhAnEauSrXZs
qyDQTvgHUcyFGkIcxPbUbOnddXtv4WSVycRy8zoxDyOlV5uQBJUesyxrM8a8UnAswAupsYMP9YSG
OacWe7+3MrA429N/W6dHaMwyw9DsSx1XZHUVmA1dYagN+ccrgPfROStt0xx1QM1XqmsLl4/j6DQo
HrgTHM64YdXKn5l3Q6hIYyUEX6UMAs6tgD7OiVkVdZhjuERo2j80MVJLaNaf8ABKt2SpbTltXP31
Upy6z6oG5bw5ZIwqi5u2qFGbceUZxKh8hNKtp/D3rxdKTHljUh96I5ZaxqJKDt6qVzV7aSzB041h
B8O4pQ12hoIHb88huDauywAmr+AQ+IBxxeSsSbmidl0Q+x4HwNPKd1Uq3UWrsIjljEgaSVeiJWhG
eJmdyuVfO3g3XZVppLAI46RMRAc1rNBs0w7JwLSXZshMTXmhsZrzPOGesUpDqYlXXFwwFMz4txqJ
2scQBNNGkiuy2auyREwNU5D2p8EaTldUiCFja2mtihole74WxLnT2nCa2WsgMXFVpCBja5VVUMRB
mMqZrZ3Pww0lApQEWxn+I95pnek1MY9sALj5nVK5QiaQe7MtaEZtv0rabzSVDdN3O2gMwWVghvSe
yBIPsyrfjgnL7+6u6tK0VgDvbBYamNxOrqoA4EMmcUfOr0hVsT4gxNOQS3NJdptHSq+TtlbReEp6
PNx/B0jHf4I0YGejE44Uo9BYlxADjZIkCHG6jQ1AwVbI2E3CdAWKPawlj8a7jz5Umw/ODHz7BHYj
yilentPe7aC8zY8IKRHcQQpt2SIIqHEhCjEVywlk/E4M81TciOKBNDXtdcRDma0WMh4PxSR3Gczy
RSe1AP/OAPXFpw/Lfue036Kyh05kAAQ4uaXCD5IJfcmf+i9s9/m8GsPbI08xja1GTkTLW6UGfGcS
Rlbtdd91+FLDdWPbMbcGRT8pCU5agfe7LElp9OSkYQtoFmoTFkVhEDaLxSO+/jxwyNeQmoNDVfDQ
8jy2ltwnGsFdVmimpQs/t83TENCaowSARvkXG6SB4CAC8LC+ltqCzjL7nGLFj7KqRKoSsaP7nuKq
jajiMVU7FiiA6UOJ62e7oSm3nrutDkL/lOTGMbguLifi60N58kAbC1GcwSR4PpqcYTZFTp5AGxkJ
d+56POb748mF/x1Hgs9UfSCBD2GNY44cYBQXxWGqlEMPNyTMGR5kBFargvBHH5SEGVP5TlIB2lSJ
Phw6yzzacDwyiL6N20a0RR6iBZYhZHRISAGAz2w9TTXvig8Hv4ANKnIRtiZa5Nm/NtLExoJM8iPR
+oxFnm58LliIUv0WJZghhnAOFQj9OBUJWuluJOdZqKiaTsq2o0yMG2jqya6DTuppyeR4E9wcMbud
hPzseE1KmDKrzZ67IGLnyLTqXWq7Al3tGKUEcb3NWn8D0PfNeAEYyUTVK/dr8IkP9UAfaBTJh6bh
teB8Va/U8+JHf4z1wrUytxSz7xVQfLAI77bMLP5cHka0ivYJLET+wvZjt3mfMbKfasY2pwc8EJMB
CP21j2/Ssjvi/hkFgWsVzu0SNlK4VBKNpDG789GDuxlmf2L4gX/qlDl7x5X2Js+/X5dr4G7Tuj6q
st4C9L2WbR/5usQiaZJFc7raOGvgtQf+H/wxoYKJhgdKKy6W6ztGWcccJh+TjOWKkj0OltfBes5L
RyHw3WOi8KFI6yMstqb0ITVc76fF6lxRBqhQMiS6++4pT3Y/UnAH0K4YJF8D3eWOYakn8Rw/PT53
2c+fZoq9fKDvb3Ztyxfck1wmLx9+BhXQpF0a8OcWyVfeIuIzSYudfR7/mPdTvjaX2JxUKVp9j0Nw
32GliP68Oi5BB9qoO1M/yq9Hce81DZZxx+jJcxPgrCPmd4bsc2PG9DHSmRc0y4ISSJpTR9a/Bwea
i0ZNYYVcbRAh0li9yXJEHpmqpADeU5huaxTfs13wgiFim0dCEAwHGI5U9HM47KBy2SWBYa9/ROKM
JI71jC8xGtzPOHZBgaPhbYtmAm9pje2BP5lp2qi8p3PF2Mur5tbFGEqfmWGixRgVihC1VQD06iia
3wDDaQit4Kk0DQz+ea01pLuu57dYWa/kHhSC56QCRMTe3zLD7kbFKYq5KTDAUjxwA8fm8sV2Vflm
rNTdm53r9/Z1+fKsrebeY5nngQghYX7dKoGwfZ/AmUCEX57m/gmnMkxauYqWBhOo5E2bMw5Q1aN/
y324vDIR+1q9srGVSrJbu2iBZwXCihomrM9XzDjcfC7ZuO9D0BkzwQs0M2ehKTQgdK2hUkTBDXbe
uziSXQheWwKYjHebpq6Qct34yOeIVovWfi3jY2avlIVapPpx85QzfKB8+8WeK+1v3pKA42589oRA
GhWuQxo+73Ti01a+6G0UvvaTHzSr0xvH3oNlQmSJ8bDt1YOxWntTP3Drjh0KzICMACGGLzyikLsX
LQYiYoZhRil0jwrFZoLYeKKB5jBqFix+2udCqqv0CaIjf0vnoYP1xvARuWdxx/oJg4hB/e5LclcU
RSUIPILgsc8TQf8Aky09TbvGa1D6VJ8qWy2wrfIAJPd3TJl7kGQwnYb/s/3BI5qRgBnFGxwwOnB4
vzfn/y+ci+25FOJUqK+dW3arChZmxUrZe0faqAxW7BQqx3bOnR+x6MoBP3ZjsR/mLaNRtAVZZoV+
jRdFrwIxdCkmRurwtpiqOwd8g69uS0j0HCcqX0wIlmmQ1pfNXn3135T5u983bAqBfj88MNCaG4Sj
LctVMCqZP/l+ynCCvs/0DH3mTPKHxilp+lpP+WcrjJati1yi4sfP6GOuDTOeJ3YcMkFbzd8gYekK
vzrrmGqhqauEaUwqhGCFXiUopH9fwtv4zqx8/O5uL1OwTDXIQ0ZF09+nB2gtSf2IWy3dk/ng+PGS
CrmWXghuLa2k4mlzdJuHSaml6RwlmLdJg5qMAr4eHPNRbfimsKH9sEg45gKsSkQF1uHU1ZZGavw0
qiVHp9dLa/+7M6acmQVEhLreY8XOMNnJbyLk5biCx+eS/wgFQ9jW2zI/f8YiZhsa+qhnzcA3FiNb
qxTR13rltyLJMuLVq2wtNH23fwkrrzm409mMojAN0t8WK7CEAGOvPD4ZfPim0QUkVUcFTCVPbVzl
ii/N2jYlnHbdQcr44J5H/6eRjFYL532U4rMwD4exNVMe5cPh3CkQMQk0J5deEX6W1vwF8p3xpZAp
ifl9N8mFguyms3WyhoOKYEV9rBGIjvx8nbm+wG0c0PjnBdYxLDx7mWqgdGv4kzI4UQ+IBaJFzI3C
SMmOmN1mtIzVioHqgB4KUFBfYB3NOFnMJN6+2iTvX74aY/TdRej3saCVwCNvBPTjk6jK5rpIX21V
WWU0Up504FmHzAcCoFKqJxVXxwgZi3xxBa8muL3kzw266Zt/NihUikgKIPRi43EPLcnNV+IYPkNM
PeAdEBqQVR6FtHrGQLTV3Cw9UiVG3UhuqPBovFxC2ryFXedxWP5AwLj74z5+6NLiAiIlPJxRH2qF
NMp2THBu8vuz2+17ih336xJNDd82GPiVEX4Jo4RGno0K4uiMe6v5kHrwKMhEXNdcr0V0hWV1mZUw
vH4jYY/sI3oqDp7tSF1QJSMAJxmmG0crnwpeLo/E+kWAqLOKAghyRzDOWlJ9uDTtLg4xHPuBaK+Z
noJHqrrFmh8Q5yltlaIBGXQEndGF2o95R+N7AQEFHSjRIEwW92xjgBhTG+Tx8G37i4f9gU/P4MT7
6rvtVtRLJF/o6cq+3buM/0EdhXJT2+MlHUvrlwbdL4FMijNc2x0fteo4iJsCmlgNFSOh7kqkh0Ma
d7ln+YgeBTpPOojgynsL+mcutpNEq4+raDHELPrPAyz8PQa0U0HOnGEMr8tETU66g6Snx6Q7GRZI
hSyqdhxr9bhcJ20SrLBv8nDZ3duDAPLHs+Oon+HlW1g5E5n21Q9PKLfMMMztpL58cFpu7qvPHpek
eO3EphDVnRj3rIV/MTdMdOyjNhgQbpRImSituOKLVMhIwv+AE2E/3HAYYo1NUer1xmii/iKOux2j
k/C+Ggala5bAE6Uza1MQg/DLwSDqoDFg9GXNpsOVKe/zc+VF9p6VwuItBsBlCBqklWRFeR0rV2XW
pyZklsdlkixxeHO9k/E6f2p5UPMiDXSKl1pyo6JftqY4xAcsP83ry5dTrOlXjEjwQWOTcqMUMRyg
ZDtE0kgFSLkIltD7gFkbhIbFTsXMcLXmsq9XT97+E9JRDEBjpLBHQAoo2Bea1mrBPCJttNk67WPC
ZJZsCA5xqFpHMP3cSxPH783JW3YkcjXwvpFLdFRrqsw9fIfL6Ym5SKmMyTmyrPRn/n981Becs5Fm
VAsikVdUtCek/thDIIn64d15nCnma3RgnMJBO5V8QQxoH7/BcLOhGUMVilnwid2nRcjo+/IBqmbf
nYOYZtrG+3duHq+1Ivo7k81drrlWbooVBb/9XsNBvmEfwdYhT+JmHT+vtqgGVR75/q/aogILMCsw
itT68d88Ws+QRVi/Erj0vyb5pX7kQCNOYfaaHZFNW/hIXtCrQjetDlZyb4JVHMeKA0u+SL2WtYzG
cdElnC2qT6pk6qhoHHPzEOi7TkzA5fUwmfAsB2d57HDebEslAQjSOeTDqK7lW1rUcnzJfPjw5Bxt
zrW2x1xlZzbHsTMu9mh8QrDqs/oZ4xYFfNRduUEEVU0eL3NhHkYNjoTI8UePGeyfGDgddHDRxbEz
PV4snCtO4IM8QGW1Sb3mOzohIxwHguSF2eTTJrdsqUvui2lJMa+VzXf8MXbhSzFkl+Tpdq+RjBV8
L+suekDrEe1R4FkobCV5hiU/Fvc2fYV0qCqi3UKhLtVZlOaDv6wSg/7ttfchNKErrgGnqB2AVQYE
jTo8Nwed5qiH2Y11zjPWgg15l10o8nZ77Xh7P3ZyyIRU7L9x5/y9dJn4aZ8tXhXKHwh7WKol9asA
RYVv71KpEFvknWD32NdI7FDTmKS8XenWr6sOiU+CAxpHspg53kietcYhsdZln+972nfOgMOzywSN
LT/hsYUgGD0dvwJpLmIBRc4HJ8G6R77MZlpJhZAjNISW8UXrsplR8Lo+xR6UyDSptxSImGL9dF3W
T5bex7L9qvpfnIiLdSyplstqiFRz5WBv8cr1raLS4UqY8W7IDAlOnSoYCmlzfkg+u/MroRcxuklb
TiSLoPnpHl4eUTTGDQb+YvgxyOPucoOiOnP4y+b9LVJ9WjiuMh+21GPjAUyjXxKM+TjouHY9QVEA
DEOVLW/4m7DsJewWzbiD4dByXx9UX0RgORIUJ2alX2A+G+ZrH1812WITdh95g34/Xrn0numyjCR9
vi8ddmKxHD/1VPwxX9WdE/tTLje31eiWwuiiRckDRxLWRzhLG+14zUW+RAhWXrtAaCb91sr2AL7z
mH/o5+s22zve0Dzu+u31sc0GglQ3cpNC9tf5ZhCIXji89Na9MStn2zncQVXMX7zbfMRyIeFOQy05
SJV1UZ9Bob21BqIKTkPT/HdJG0hy15uV3lL9kfiuVQEsaqmQMMeFSTowjUhPJ7kDzLmnSeYbW+QZ
nfLFwLZFH4zUGC1yOMR7aXCGrO7P5cYsRAei9AdyGYbqiQrKi7QHsD08EBWHhXWfEfEDupT7vW2k
7igmrWFXDuxUsppRAqQbO2zOFFoFAAElmxoosrGWEmqgfkEMj9nacV/mCApkBG5QedpAvmjEp4Pi
TDi78ybawRdA8pH6DJOda71GvplAJ/uUFFpYFlosP/aJ1eb3QZq327dZD40zWm3bJ5qU4XtOFSB0
N+6vp3kbcZ0GmK6Hpzle9JixdlJQpiS41fpHqfrDCBi457mFdJxPpOTT7t4BrRLvTshimPv/P9Ft
bHkE89OtQMP17iUl4tv+uUazgS31SHNlgmoWnGOhpZkBoIQMwnkk+zFoMdBkbPPo32hyEcesXyEK
y+3NerZjTdoK1FKw6kwrpnRDNQHe8Wfa1Dh77UPQDQ0/aUUQN9JS75KtObFKBVhFzu73ai2J1xHi
gGuq1oA7Yjx7Z4Mzz04+GT72d9IPvsZ5gAVMT24qxUcyHbqWnnpz6UrOkEfZMiIJuUaCze+IYx0G
zUuOsPXESxjmqRpLkzcpi4hyXJL/ZD1qnEDo2LXsRYqH4+nwggOgu3lX+0bzC9UVNK7lBU5hiGYD
mTroXYP+5Durk/zDDkbwtYynv+5FuD2bhM+uKImG5lLxBJXAZsSf9pzcuIEryIj61eKy8FeV9X+J
wg5dvhru7Ki6a+5nQrWd67jSs6vJDANCanGe5zZQ8BuuBsldsOr4QJnNE+AAL7KpBaduG/tUePKt
7JVuscIeJy+z/7gfQhGt/4GfG0r9W6XGPzhI/R718hlH4v1O1dV7oldhbjbgQY5RiatJiFrOeJuf
Hh3JMPX0qeGZQZL+q1qqDtv0wzVaev/RI3vukU8pW3+DdZzv+OT1mUG7nVs7XxKNqv0X2x/BLTn0
ACMhoXXJXIrFieHNdDvcSdVHGImum8sLtNBIFQUvXka4cck26bPHpAOyfeapzvUhx+RVKp6Pw+AT
WjxuboZp0p5tOm+rGYHRMSo9ZKZmBm4451bD8/aReVokD9Ff4DC3BUPsWfCBnuZ2DV8+lgMUgljI
pYutgKpQM1LemoOcAUXrlLd4YpBc7vq/587OYucE16ihgxkNdeOCuDuGZ+VURhpA1JG19pOXikGq
zgTdaw/35tMUWL5L5OfR2Z45fhoHKWPVh835WMS2q1iOvaq0KLlIApN3RBJSlqWWUY/nQnxYM3aU
jciMP4tledVlWiWMV3n6ESZmwgwxXyjYR8leK6riD/PX2lw4OmH9eze5Ph9j6BDpCqZHjTN23wS0
G39mZrA/+bG0uQLTHRtDUV4aiK5E3GRJ4DIgFucrJEoQDxwYf6KduHPFir/aQQDIcEKZd62wUpVz
qZrnddJj9HfoGHjzQn/UjvWrprdtFqo7cMMM7W7PMbAiW7cZcVRaGpDlDo3bkVVuyY3g5Zir/2Q7
tgpgVOKL7K0k5pCuBq8ExjOXbNnN1jIddlsMUj+6B6WeGBxhJWuzArXVKv+E1psSgdPL7zaNaFa4
5MF0xJ5DAspTyhIUB4DYO1IUvy6fnKtbTmY073dEEaGUY0+2B5QGpJoL6ZlC6AFrSOOg9id7+EUK
Ed/seQfszeu/ZN8hjIvB6+crQSPKVbQK8Xi97vniatK+DFP4UOjV7955/7U/aeaAT/R9yOtGWTJy
z9hBcS/sUdhgsT3yeX1fcfFiXcLYKfAgdd9mps7mcnuLEoxoxA/4ixP0/FXeYhxus+bo9UTMS4P0
U5mu496rJbqCEDcTInud/2xWP8SSyw1n29JzPY3Cc5hcgLOq8Qu00mNscS5+xr/GfHnmQKJyHq9U
UWeXG8mOGlZ7FJfziXKcJwyaH5YIy7LP/8Mj2XMo7Dz7m5vZ6uqMj1Zmtq6UtLX7aCErhv8QgK1D
uiabqrLof5c6VWjQHHyuTNog6aKZRljMVbqPO5MP3zIiJoQHdLvsX47TOkizf3uykZYC0AjH/aiX
GUAqx+qzRwsN5bLrUVXxv5Ol2c5cfLtpmI8tv/resmZfQpCtdvLrlSgvi66hIHYTt2DT3cVrA+Ha
mcv4SD9I5tvIQTjYyh2JR+57MLXNaXkqQ6jbLxv5IzsE7TI48U4lUSI4eJCgFs0uVaQZrFd1l8Po
cbUtsfsqFzdcdYKvhdxJll/TaORVZ8jikuVeYh0R6IlLIPBiK0fNj6E/aSd00vVCQs57DPkgFGMe
7B3HIRMl1sYQP3Q9zhCo6r5tl2YH4xCb3PcUBDc6FnrePH91uEOXWJ8ZkG6PeWRxdgoBxSv/zToi
kUt7b71qbEBcSELuaN5X0Ji1rrE75F4M8RgLmt5bWQzJE84LCovMmUuQXt9pC98WVPEWlTqJehX6
Ax+FQxdOEhaWvscRiknvbiXe6nd09Rss0Gc1AzjWyKqy0vx9DEhG3n1vN1WKabB81Vb5LmQk63vc
5VA5VZ5FjLGsM9GgQZl40jMpOCINFMA1XlWb13kEgVcdf0wHoDMhDrOo2fcSNmZb3kyQAyIYz7e6
RtrCRWi+eOeaEtjSeX1BCUB4oofHQr2Ddfm41uc+vsi5uC/tPwJ/7YHwc0YavrPzxgl0VARGy6zj
lmx4MCXip+W1TvHO7Nck+tCNcHaTB/El3qMoVV6/Y5yPB155YhgorBN5kqxNP5qQIMkS0gom1vR9
S8csiLYO+wGhAat2+zf3D1KbHNbD5QpspWvP/+IPBOChMrgBr8fqMfTbu+MoOU2DA7Uz6FwBSHMB
tMd33zkAekJ3yyoM1P3KM959HkTRYPL4fXXAKqvJvFH5xHKNpCToW/j7n7J7mJ7Ca+yvkgJUT6LJ
WP7s/lb2xqvSbqjs3bcCbCWSqdq3QrpfKY9zTjD3BcJ62Xpc3uNOp3QVo5s3UzjywVQznAN5A204
K3bmQbclw+6Ef4dfUrseGRt5GIZia4z9heN4/5gbfVzSXi4yN8H0x/xn13f5HJfM82F4lu0s0tLW
WsJMtCsaN98s6AyGh7t7LmpkE5Oai/VWOWqlkuAAPu5zVMq/wWyViVN52PZQbsinVQKzWDw4eeXj
JwN3UAdU+AVzlDIDXrkCNSeqPfVQ1H1Fd6nHx9hkQ5QUQIj7ADKMwyfCe2hCxe+Apy0vK9BGikgq
5H1wdhPjEoY/rGquDLe7Sguk8yZqXEqtsSwRIKejCxtqHAajn1WsPVYRXsy9o7eErms9Y1sWqpcj
xxJ0Ar+uf58HyKSCYhmiP34RVIF0YMiEHmZ00+WHQMEdQOTEYyM27ogF0qbw8l+ZbIZXi3UDUB+E
CRFhTdUm5fo8P+tn6Kwe7iMSMj1NbHX+uZGX/xDT+1PHTVqrLR32Au7eAxLcwQYqTSF6xn7gQFZ9
sYfSv6IyiLrs8eiAdDsMswV/DkEgtlN88x2EufYO9Y3ze8/Jiuj/O2y73ycc5sjwHal3I8XDs2o6
mSnfE/3jZQhoZJu8YE58WZk3gD28mpAACS/EVpEI1BoQH9ipgumxDSWWd7goqoqvDY9o7adgQ1cb
NzyO746QzNCp4pDsLAeEpss+RVuWZMZ/DJn05MreVWtTGo1/eHjlIK4X024ujKw85cOsfqDKR2c7
VOodYUxIet+zVuO+5jtPP8CYQnAEAr66NgKNaLei0Y5tBruPaPDunQFpefDOJfsoeFL6GKT3GKpD
eI3dkegX+hqMSDwAl6l33H/cpPIdf+JVw3T00vsjAVIM/0kU54T4n3iBkI/zWx5TWJfqwwTJJ4Zx
oMjNBpyByA9EC6N7yp0bPUtInnb9rATrYzpKEv9EGQwPlrxTPkm+m0v3GNphBx0WUOR/RnxRPRK/
8OS4GhdwyZy1kbDo+1KpF8ZRBcCE7FYiyPYFsOMSeTXAS7qx7XpWkkfL2d8Z+bHfmxmHg+C3lhvT
AqZmI+PVmAj0hmP/A1TdeJERsdfxVEmCgtyV9QFDZhYoJ7dWP3bNdgf+6JHv9d9DsmTp44IxclhJ
toZ1YLZrWLm8PoLTaCsOHWGeA0kFikMgxSmKM49a0CV/DiY3xk9zR3vD1cEB1ZtngWt9dp+QfB+F
WfUKQ54hXAgzSXZp2v++eZmKlFxWiI0GbQ5WysfXt9yxaJtG71lm8cv8Z2tt8uyThDY9k2iTm7p3
6roZKHB5IlyQvNlfC+r9zgjmVybqpF2WRiHGVMuBWoOpEql+ZNmprIed1W8in0FmCG5NlDJPfKIg
PsZ7SJ3bi79cgr7A0fj4v/4HAFiaZxA23ISNVAxU17OrsxVDD6njwciQkGjIUqqM+LTNXI+DtSr/
ZBhZRhFli0QKRwd4SiSyhCdYMIoRvEji/7AH13IKvTzvkBImT/yAfuuS7Og29pUtpqdpJ/2BYo31
mkMsCtfIQxyWAw5ri40bLl6leGOUTchIwKykNyody2s8A0Q57/rCLhkIu6fmdpN3qYCCBgaYkNmD
lu5TYb06nCyfQwfts5ZcoEjbd1Wcu+mi+i3MEUsryTX9m3o7YV1I3YNmWKvPNjwcPSTFWKygG2bw
mjtYePRM+eU49XM1ACBUJGhs+8TW+/9Dt+iKsDiaoNruCo+vEVDfsZ5htOTfAv8HE4BKWD0wjkxt
7cSIHGlqaDfW3p6t6PRne6/ogBSqCrXDZNHH34edDP1gPpsvGcfb9DeQrpCFzP3Kr6RBUYW1DbNU
52BRT+Jk/CvoCddA/wW3WrdXLm7m7D7qs4nrswyqkCRSTbR4ZANkOIyLOIa0qbXFXEjfh071Ojl/
Wd6SDbO5amGPgKrCmWp3Il8GYy9u4sQmIIMnMqfT2F0VwWjFlaFbB87D9xgpwCsdVEFRXT0GxewL
+YnGO1+zRekrS60CWiOdx/dxdDxXG4OPWx7UvIBfalviysVS0cqB0IMiTSifbDWH7PoOioCy2lsF
n3/4Ol5ou4wPVKZu7MyCjyWDemIyChE6z1rfGW0qdgoBDoZBmMprj4+su1C24OisdWETDuMVskwQ
Vs9dHHcBGo4hoMdIe+FtyRfPtovAjUkxkAxFxgVGKega0FW7JVhFcxq16PHrcPAswwyknEB3E4UD
URGwh1aQi1R6LdJZAy6B+a/bukVrepquZVJqWPEvp770QCIujSbLh1M76jYoVJJoKBxGpcYTCCBQ
xyUdMAnzN8Dej8vLo35iTl9tbMEtUb5hIFgbY7M+E42R7rhvp1ZFD1wz4M1UZlDqTa9nii89wc9x
t+X+aAXOz3h3lIebejgfpQ/ERv9mGeGlpmXxksaMWkBgEqq1qri1WSJvTcHC/T0CrEMoooNT7Efe
qJ35yVkuu8afTTLGrfLeeG6mQVA2OOjHJbzMm9on8+g/5hCq46qHGwc8/G4X/2nHK7wIgbWBhGfS
WiqQ9CqsW9vob1eTDQyQI34qvfi+7pW1oU577wD0nRic6fQfJj7VtG2zO0JkNA330jUBVEIli3Ze
77ddKNf7uhZGJ8cimoIVDGLzpLs23bQpuepsVDC8e9eIESZyCcY3YHWoFj7hFPFqbyxa0qTrLLCk
sycVU8VFZUMZqLEzE0tESjAJVgLeMcx5BZjyZ3+SZqc/Bkf3yX47fHIsTm+8OJqN9pdCEXuEhqwv
GFI+Pu2UWw5EHgsh3GIqG2R+iTiGiXBBUFdxpz2L9aek2H33vA949hsh7BWj/gj9cT+7vHvEARi7
sIvxpSYGwovo2zHIv6VTisROozjcEVfgj3S8WvaaTuN+G2NexHnkZfXPX+2w8DeyWSM64LLprHCN
y+TzrHX+UBeRsbN9yhFGXoyr56t2nm+euIaHHZmyf0ulMSyV9WBu0czN2KV9CJEh5xUTxMfD8y6j
ANAr6ltJ9VYHcDlLVIot/P8KJK7h8bzOie8eUslFAMYvTG0ogUBYyVUn0jo0CG4SQGVD3wJwQt2H
KLhfKSMQNc09Hu1PxwiUttj2I3CYHefpjs/FRanjodMjYNEehotAL9ip6TLCqbI8D/A2iQFmzIkk
DPzaM4/K+M56lpw8p7/jt5RsFUHv+8LC3SGKiajHJlHnTp3lVr+rUJd3480sORY8fZLKkvOIz77s
CgHrhqAqlOstdQufoYuV77qvOJIaHcTjodtzico0FpNeW3ZtxsD4PoxX94AecfH7xT8sxNvKAy/f
VGpnE3pA+teAgLiirhco9OVzjQVanG6XycN1kEuBJqomDNM0M+Z8rjMB8DogV0H5QlYMVuaofhgD
BXcdPMCqU6XPPDXNh3sUiClrOx3gbIQM1AVDs0qo94A3Bcu3rnUy4xxvPnjmmQ8OgpcLy90C1yGf
RYniccfhj56jT5pDBn1/8QsodOPMyBIUoGJSK5wGkpm+GCIA4cbE1dQGesWFB7vxXC2K4hVLD3E6
mFdy1hc2doBSLlrt1AMm7T+vr/uCfyjj5qW0dTLs8wPH7NrtkOGf32RqFIfl60q2Hpjpzk9zubZs
GG5JzJN1JuAMWi7Z/sryJeDfGOZtUiW0TN20FmcfighK6PUPY5Ku5QgiCNrcBbmv0/6wKkfotZHg
iLP1wi2nFTw6OQIgzqmBlxDlt2siuWfjNWlJxg+cuVM04p2+tlqB6kcJYBaL9IA6+pbms7QyCOiI
6l8qKME7dhVhonGiB8ZEOS3eCr2W9Ir3qm4RP0hTQsHGQSiXxEF4SB8z8FxdatrSsnJ2reJ9pNHE
yXB0yalGeFRsHs7tXZ/y0LabgIuKgyhi5dmk8U3dhqDtMqzmOeU5FXukWtjFn1kU/FbDJxURiagG
3E8R/YzzVwIU6Q1BKh3vI/1bAoi9Qi+7BsAfCM0jkN+FozEBQaINsejMNPr1C/3iA6Q4WFOk/u5v
ekdq3cPcn39JXsot6JpP++nh61ak8f+1Qmfa7OHzlWI/H57CnF+TPOzhMBhVg6a2K/fcw7mQyihX
3TVqUrVYBWVHxxwmP/uYWPFAeRJTuCPnJFl3l7ymaWo+TOQGEHII4YhcjsZa/0KI0v4R13wkmrcC
s2psQNcDIU9rWLGJ2JdSUMgAN4LnIdwa4xenZvkZhzmYEV2Xt9G+3xztOeaRv7SE1Y8DEjuV3jNm
EXqqHCAyAIK/irVvV1ebFFoqbZJbZk/97M31RWWVx85ele/MFCR9xOVNFXtnEViPgHOFv10tAqVf
uY520wAZY515YpGSXR8KAeGfT+qK0h6fF3QE7w6cMLPKCf23/88hwMxpsViQv9vBPpoX4wAMuiq8
lSjWLVT8jDkJcqFx9ZLMwkH1ojCGlXS1O5IeyDhX7d5Jt8881Jud0fM2d3xAq5Yi5/vCl2kzBJzG
0PghOxW4Z4xXM7y02aapZ80eyDyIWbKpuINnxyqPYSCaOQRHnnODyctpjS9985ATD81CzZ1G/bIJ
kRxn29mpIUs8BZNwVp6l3uMGUR42TnNJ2P2uuzhu32knTJPElnuovvJ/faRFcrWWyq64dyeVbFgC
3uE31Po9SuE/IkMQ0jO2rD1XwdwzrC1H6SNmCfp+48gDT4XJ7zGQRVM1f1OyLgLgdwcUDmh43d9u
UK2lhuA/1aQEy+/iIpF5PbhHge00jv9Ndrde7JI9rmKsoO0DdAqo7/B+RoQo62FiGRi5kDzy7u4T
AgE/2xZQXZF16lUsIc0QDl4rzZKeX5bY0K5vmIxXQKjPZ0TNQlJ6mIyStN4yddoM9RRdbTN5GZAU
XOHILmiMxN00MayrQbJAwSluH1kk0BpsldY5j9N3Hmk7N1v6+Fo+W6xk/Q84JJ/E+KNWkhvH9ztZ
xczBbRGKRRNDjrdrNBhBDkPXEVdSDKVpCk5hoH4eGTOnHjGhSE1r9Eb5JEE7xDtlVtk3A01Dt+3E
hU0s9icMB8Rc1QmdRmpA7vJI/zawgZkNVWKcV4Zf6HVyvjSLiN1moVH1vp4kuvfEtd1WhjkCGHzW
wUU8zaZK2KYyC0iXiJDrqb+3IjgGwtgt407ne/WTBg3If4ABXfiX4H7wZ6Uo+EVE56J/h/ShVjAw
lXpUVHafj8dHhtugv7lVB9EZLbsgQzTW8Fw0VAAQ+WotlGEXly4byegp0cqg0Ht+neIXlXX3yp2D
tGNccXD8zwsnFegiEKKU58JLRNrAvpmRdeBuWrWLqlSRV4R1iC7wkzTmo2/wf964Luc9T2unenXC
FTJSjsB0+Zr+NK06gZOX01viLvoByKMNr+CErNqpj88DWeAVEhM7Onocys2oMBW2atajBBb7KJZ4
Vp3Iqs4n6bt6KNhFjJnqnoxQn37qJaDjfYE6aMcIQISmp3s9b6Y+pJOOVDdZ5fhbU2eyEJNfYYGG
yYAe6J8cBAVMfM2/wjoxWyeDT3a4v9eiFm5zxVtY2YWyiunnULUDsxAenQGUXARKcOFmLw30KwQK
c5TeZpCxXp98XpX4bHi1t5aygZFUDVkCT9DlE3jHDozcU7fJlie7Off+VGaZVhjy1IgQJN2J3i9t
iq/gCZdiyck5rA9/+I/4GOamivdrJkfCZjbXw5FH5taOisYdyI+o0F+e0PcIAr0IXS9vPhcHJ1sy
GJEpXmXzmdIlhSXwjzYvmkuL6OHfGFw8H/pWxxYvOfa6sKu37+bRL67Df8OQHNCtvdF8XHQrN1YK
lWZPqoY/Mp3ibazgjuEpKhDvOw1jLD5vZ9dETPa6Vv5cuIJ6Rd9TKLAeGohRq+KzBU1Raz+2rWVq
s+hMTgh1xvCuqeT9K8k/y0E996bFUk98w8K/AC8hFWOiOf4MgHE6Ayvd9BXr7z7s98aH2LRvFRLn
hROt+he+lFl/AeB1731GzuvraQHpAWjbJQnomTwbKkwVqpF8oNoYpnDXby8KaI/nf7tTCxaj35V0
WPb7VBTCXxTRtPtShEVm4qiuqrijurUib45y6dNdQdW/q79C0yafh/4ne4aLuzV5eDUIp0TemqTg
LadxC3++xc9eHvIYnwzGfwSDqLEBrxqfS0fqq0pt1LhCZDTx+AfTg9LyhbrqlI3zrieWrxiybcdq
t7gn0hs7MOfQNh61Zwdr5xSNlLbyH8yLx72vciry76Fk38ayV8itcopf/lrY1gUZz3+pPVr6AoLp
IhegEqNuYHOC5NDoc41lAD7uwqwh5gWWHm74gZCOpjkVdW5hcOTOGjfxzjF9dbbzpFiO1hYdbKjH
vHaBuOjLDEiiQKrAet4IevjynawR3qrvgJujxsgEm38DVrNhFg2rI8k301HlBvdeVnkJzOHke689
a/19dym36yqf6FMJ/pZrP2WKpNDFCvSPAe0IZFnLMIgS/kHxkb/0QyeoMmuH511LOW6ZqDfYMSvu
B8F04A+qCUXzZN9RoggD4FBRvQx8jUxF4CXQrsi9DiA+EMNlZizLuc0walwGTfFUkvuZpdYnpuJx
65kVYvdPkLrn961kLoDrZCcMLjcU5SShiPa0XGrfMTNJ2fW04Gr1eCcc9B+6N03K0uq7Xowql/ed
daJtJfmRKvDs5fcK3himSsf2ARtASsbOd35YE3JVMXZucRa7thITd5yy6H/CuGmJAmqd94GuHLug
fuVy0iF6eJKtaBtUXpF7bwHsT2zEqms//7hiWYfkG8g/jidAhxS8fLx7JtbC1C9XebevYf5ChYGS
OpeYUQ79yjeIB7dj3dQQ/yAXdUgkogmw8yvovAmGz2HWgaFAa3gyjyCfY3rTF7X+4SM+OpSwaRNC
xnIWsqYcSHIWKCBB7ZO+A8zXthFaWS/hs4dYaNutyIQrTP0hKA+qH4OVOqor7UcJp7FL6rF9Th1j
zpfD+pfFW4yx6xGk8lG1ECzdjQhtdldqrVS9y5AP4yrQjm017KkCuHwHuk9JVZ4DD2WPejU/HKSy
rG2ne7WkjS+R6QLk52WT678YkjNxqdHpVK4GL6RzZ1WR6L+TRzaixVmTdY74LxL3C4C5I4mAyax1
AjjdmuKq0zVDQ0gX28WZUP/Izmt8Ozt0JAYI/iZ3k67uDngFr0pVzYbsMwvcRcHR+AWv9EjT3E/w
y1qUjQ0fmldi2LwNcUqxdpdJbtUuDmp6SabT+w4glFM2PxRjzHx9ZAbKVmdNZa9hUNpNvdNs75QO
I1XzmalzHcttDIUB/58IphVkDX6fUo5efEU5G7/AUgK9t3QzXapVfoS16aXmRgx3TgHI3cEX/irL
M0fT8U8ZOkOKKsfsYrKc3s6o6DRj66JvmRpkLazVD9LKfUk76IoD1aammw6X04R29XZsSQzpxZi5
VHjKrsvkSlXmjlhdDlgTR7KiWeJjtGIFue/SUqQhxhR3970s1uLRWKbo9PmRf2SDp67Yx1CEL5aT
Uht+0HH9RsqId+r0c9k6+7HVjrCSTiLKdBnt/tLuymPxX05sv7f7WnNh3SvcyIhC3xJKywzr1Igv
4eByA+yer5wVybC0xyiWL6MleKN709nUTzMXiSzQA0LyefWKgr9qYyUYI/JpaS3BJOWUEJ+1sT3L
/p7B3KPfzFmnVVEYJ79ecHmYeIQGOv8r+NJEkOE4K1yfSJxKXRQmwTAJqoYCIui2dIKdOkVuTpAF
29fqHCzTGWrGesU383iKmecrTHN1FbTeUx3Ct0H5L7daQOPNIwH2tauG1f00hPQYpGbpqcZuE+qn
8zUX78Mt4CuBEGR8KoaWXU1zT+dx5fIZDzw7y7a9MF8/NbmAE3DHrtipM3IZKYC2v31JGr3BKVQ5
Qcj+zhxe3EkOx3bY1SNrCaDYRB9VgcKQneJaKjBKUr4Es+N8SPCYyjmfV/1ea3G9Tofih+eTkGjb
VQH8GOomJJ1xp/CT0tdPitEab7NywQyUqjVFhCNJD8Mv0LhJZT25tcpoCMbrjQoLWER7qKfqx9IJ
oFEZkwN2frQyoJ0LcsFZXxa9iQ7D2HCnN6W98WwsqWUYB0N1N3vdSJ87VqLNAzn5w/o8EisxZgk9
9rTIY6cBQ4zqeqgTXyB9ryVZOG+KA3spgpssZE52yHyFJRgd17lGEUeye5IN1cwMnvyn59cImYZ3
NRongRLgOPBVyrawZgt3tYArewIOjPOVZ7uWsiDBSFb2vdKQ2JslvPliJsuumUFVef35bRdKgtk4
W4g47w1kYdHC7dOOCtDru1flx1Zzd+2/+HUqxJvUp9zTpfu1yf6OySuFo2M121Y/9KSlqTUv53Yy
Qy0i3NvtZ6ybNeCAIBF2D0TNNxjd16+Hv2HXQJYxSUN0aEmns/zo0l07HhuNLsSpFH15Yrkcx/fC
SyAzw3gJ91lVuGxpSQtadJxnA6bf9sr21xmYtEPyDGL7TBv1HB8YrGsCk2ipAQRHjFeeY+I2kB9d
kDiovY5jkEqsg/uhwp7WAlrjqzilJkeTiRAvTJo1cwNvvupHV+zU4fzBM95d15f+E/hH+43JaeKA
GJ7KASB6epeIV8HFqpHWMJV5VOqVuhocOHMnhCglxs/GVhjh18UK/tY8wSYOUJClc5bMpXtZchoZ
7TAuTIR2nEmlPagU9xvTuVQEsrkAMmoZ4Evnedm1V3W7hbSlaJGJgQhxGhvnjL70oas/yzG8nJwv
xJ6tnhC3av3/nD6JnMLkimQ2OwhtquSlsbc3Xw/XxmRnloEuoAj6Upj8I8paC/KmuBHRqCRGWYwk
dVMCXiEqNtQnqW8f8qYmXq9oQ6qTlLOeti4JDHXkzvVwL0XJuk0RNFNl6E8CgPU/sOuE/9OcGlNu
njyKKdNifXH5Zk/HVFYZ5kdHOSW3MlPBYVrmBC/q3sdD/CQa7/ABiUxyiIFlyuKMmnQcKXTtkw0V
WciscfRRrOxOwG8h3GbxyA1AfPDvsuKrD+PNTYVamhqpIVtxiBNovtsrroy2ZB68foMO0Mb9CAjg
spSbW0U/YQciYUJpW3ejpUHqLXx9oEa4MGc+PSYFCSCwJkJUGrpAj6z2zdouy8/5RdsgMGWTZ0rp
oHyDeoajKcIPsRK8tGk0lomW3V2rGFkZ1GAZ5d83u1P9iQ30koxZTgq8/CMF7EEem697trzgzjL/
9pVe36vLMQ+ZKZDZd7EOGyM9r0R5l1G5NDsQxXYePjUIi3dmDZAbGb9Ex2d0JD0OH6MvJaWXV3ea
XO1/ikLm03T7/ia8BgMzIqzBftFRMchV6YXq6kN2Gwex29D8Pu1+RSQ0hVZ6WzbemP6DOcPkNWbJ
5acgYyCglWzPo0XOMSHiUt1hsXYAWRPtlCeTXswBLK/PG27tKCxRMR6j0Cd8iSpizoJzg1TcjmzS
dPnE2xoaWXMhLhaj/TgI7tuCC5QTPNJijGFYsCMIfcWtr8v1S9y82wpXqQoLRVGrC98iHDBBCk4C
KSi4Xj9b9CzTE4tmFzLOS3LXtGwiXIPoBoOl0qH0mW0JjzYviqb3zuVrGxnfXQKF18mqiK3ePWFh
pZqhzE9qUaqBWjjsF+NJZ5bCq50s7FIi+707uHTLY7g8pnAvwaHHfpIFpHRSJUYBhw0UC30clDjd
USi35oAm83iaEqzdrnYIwLfouVb9rdvcBHqnFraUEX1DbLlePH0bUkO4GQ3K/UQflV0q4TXRoLtL
KNK5jJYiPmzS8MjZawDVw7V9qNjlb5WYzc5s6fvmxlQeo5bnfnpRnGMB2YghVFl3pW5N4OP4Zly3
2OE3v8Az4ImBfQrk3gkC5HcFMHnpCgUljNavva57SDyAvsApu/J0u0hUQAsqK82mad9da6vU6pAL
FVazNxw2imz057//fONDsZjcZpdBy5D6GwRzGP0doRb7+3dGvCn8gSt5Z583LhbzGX6sWb0neXXh
gc0lMeoNA2JVI7+WI9KWX0Si4lUr6k4xGCIbsjkpGPFOzVDAdGbQxfPCXaSDjugfM28Cin9EUos0
FC1sCoHEJ9q2igBaKqWHEZx1h2kWc7feVUTtKqxUV0FWyr28dmlP/8m6DvXtfEVWzzYjYMGnm2Hw
wpPHgPh2TA5c1eFZ7Ii80OFpD7nMAQt0rFKRT9FEXgiQ/0j4Fjy8m//PgcHaHTlNgOvK4D5EQrkC
jvSESZ0fc1pKVIo6/KtT9QFpji7U2eVHOcF5mcg7xPkyV13lKhoy0KDWfZvwJP/9q1kaLWd6KBKi
eErwUzTQ1mtrO2prXS8ndG12SZJiR32ZOplgMPrPClvj0O4KazZe2qEeahZN4mRTG5I33/3JtbzJ
CGAxPzJWlMJFjlPlnWQ6x/Ag2UmI75rM4kz74S5YMVZj9suNq/J4bQG0elqzSmBBeNMTjsCYFEyK
DkICliDiPz4w4/35FZIDb4Hz8J8CJ8nPRLv1TeWaEton1AgHZorOLHl4zXhsVIdCzsMQEj4GWxwu
/DbkTyUwGRINPe7km9Uub5FyQgalw4JdErRoFoBhVUI4mrUuc1gGeuz7+uO7fZeXze3jYCAYBmSw
RTkhi1eznr/K2YTlNJ7lq0+R6I1G7YvpBfNCGjAHtN67zp+qb0Gcau1G6nnfEd3v466t3klUcYNL
wzjoh4VL6dAqEaCuH23QCFRDqstYQ+gitdtOpBnImHU/RmQdreAx67bmlmqlJcQu/e6+F0PlAFYG
fu2iW6CVDuIv8Y42EpS+zIVpBnQthSS0hc5cTqwgBPIsTgGA64u70CjB9u9r+uX1KKmhi4mhoOjH
V6H+BovUSB76tiu690xBJIHUXlUHRRwQy6CtB7NZV1klB/vfuh/2BKv19G2qLTvEMeDvW2Z9BhEt
f7IbKUM0XFPwvPkmy0CJglC82qGSorpW/BznlInPOQnWoK/sHVo2mZTcLd72mEmaHlSpeJY0wGuR
4ZphCF3H96L55vKiNQfIMRhLblTBDD0Vs06ORWKoH25lVpxGEVfBrY+sIK6Ds8unw/X2W86htKw+
C3wY0QALOZnun4vz1r2GLdpaQze5YGv/6dGCG/FbaMXeRV6/Et7mcPKX2iqov8+9Bj4JDOWAyDjz
YZkbqolMtzmJVJD5uvXb4nNPau8WnkfOKHrhzvDNpSQV7BXff8yFca0aGDZZkFvmqIBBB4SiBRJ8
r5A7aL5WoYMoIQzx/lzcckyhk4eGLbPcb6bK0h9r3HF3bQgBUnkLHgf5Sd5QEZMGLHhxEQqmp18c
cbLd/9pC25wfNFi2YaG4j1cOFQMK8FRSwAkPS0YJtMOmvXbfrUKgwbV0aqBSrIwf9pjrCptI8RVI
U9VcjodBxITTyyk6H7zPW3XwdxX5NDsBQJknGgRWB3RIvo/47RGZhP3pJpB3tyTpBN1ND4cHZ3nv
JGw/FExnN072ogQMSQPIp/EvQisInjlhEWyUp2hAN04LSKkCZIqhBadEbD6V+xv/Y5XO6m/vCaaM
djui3lfaD7gCnvUo2J8sDA6VfbAWPKzaXD+563G8az1+OoaMi9IiP30CTHbN7LEZ5p3ZZKsqW8B4
oLKtvN4zysgVZUUG0Tm+SWEemVSgsvOm+PRXShZyho/DpX5SZNNAHfbRXo3GlnqXxsRmYWMd2cfe
c+zCvShk+JzkdL/SrUqN9vOuijC2fQ70kqTilN7yCD+kEdYWnih4QQezfAOPc8nJ5Ff99rAP6pjF
m2sW6oDqCOpu+j57L2R7IsXXLBj7A/jf7+vSizUMwZcK5YMMJ0HHH9og2caYtmr0XxS14ZtR5YxE
3P4h0zfae+JieIEzsZlvLyIeXhdiCDzeL62/K/JKRB1DRNfXaI2jL/oO9LVHyWE+9lzPkkqFivLd
97yhnNmyAkO0TsDQuNwKww1NYHNyocVjupf4PI1rYL8W5oBkION9GNeX09kkztXReoN/Zo/IjIGe
UFTC+cC/AdX2zzmqWZn2HY9JaftpgGeLbOEoFLrUWCSFS4uxJO4r9NQO2DWnpkp7aaQTfZ8tim6e
lxyjvA2sLvV1G9jZXTaALDK+zHiqBFKJbxf+3PRHb4nUzIFBCDKmuFnuk05cafZuTVU29HMyJvBu
/+IdVZDQ2K2gXXCo3gIYW0lmcXFwxthaSXW7+19/v1snkDfh19u4uew6wBsNrFMCFfLlHaNDPxPp
nWf/9LbUej3x/NR6JzykIk7BGjtZWvSQzXlaJLzf2atph71cjAexEauVzi5y9xfwGjEJV5soUotV
FmJJ/fdMN/UXzXFB0Ujpoo3ycmmF/ukE9LqBmd8KnbG1kNjlO9ybZmgGbC7GWdrmvGD1ffKWel+D
YAUn18FEP5ZZnZ2/BXqnb0Oe0/Gn73UgKn/sXjGPJNP7qTrXsneVCi8TlY9fs6EJMJipAQ3odVaK
TK2EIOwZ1CQPrPSvinLTO4Zyjqw+PCq4RyP16cNX+vwrjRyFbcGhczxN2WH6i0y41m2y3HlNwUzq
EbErFBtoIUQRujwSH9aMHb7PCOadcIo3GbUxlcs8vcMtnsDQVZRhw+W+IQtY9lrQs22iysid9WdV
HbNBID+SOiwc3j4IKcaliuWlLiN+43p/FFUVXfn9J8by2D7E/wjVVo2tJVTEIHbD8H6ukIGxGV/1
W8j05UJnG6tDK9w2BfqFWvpPgnkg8p2CAtrHfipoqnBHEqedtOroyO+k71dgYNtgwb2DsCY4jxkp
QjxMImDftQ9cLGz3Y4AU1/6muq1jyuUR2kPfq3A+9/j07swFh0l1U6SO1K9Q8qnxSMvIcBOhZ1Bq
LIEBWXKiT35WyEZm/lPHz9pEMvemQAAs6NgkcvJnOBnPnP+yAv8jnI3tswv5Iw8EhO86pJiMmGdT
b4gyQprFvkk9lhOUhnswp1JXOCzL8zeeFYNBOyr5S2N378DaK1W4oRJgEhfPGlolAXTtwsMwHKOM
p/L5zSSnZeVu8xyGT5/F3ZDizeAO/J2+HQL0SkSo7TCnw/HYGU/OUlia6b7IC3nxVv/x6OL2oA2x
hpsCQKZZjQ6euxgLdcUMKUJhTWRQgbIqywyrPhc4J2p6iPDczCRL501IhPuL0KuoT7SMEJjdpKc1
YxBUD1EwAYr4zPGhaZrdtJVyH7IXtdY0gU7OGIp8c0WQjc9XhXz4/ORVFBBcfY0DK4OlpnkQGYAc
ThMBKMQTN6q3ovJUX735vswviKvJuSAQzrR9b6ubI16NiNIG6E4Q01qvV7s8EhbCn9g4kaCk0+x1
FM1nBvQa7iW+5PpR8Moz4+2X7M72LDeIjBnDgKR+qCf6hCqUfG1MF73sxNuf918ErANn2xudREtR
DxrC4t+4Y5itp0J4Vhmgn1EupYOG0wAxYcXPbN8D+WlGccvrX9L5f+BJ1YqNy/vWLkFmjL6trn1r
mNG+MBrhvWR1b07W0HDlInNM8gH2Fp61dH9s4H5mEvLia9FyIRrKMh4PeJ5G98aZllLoPAsDuqRd
zw/2b7X5EivHskeVJqkfwLXLaVj9LQhfrfOEnrzVAg5etCTNbI0vcO7pCm8aCzh+neXKCH28i7kC
ETpmZd2iD8RcGhdxgXxDluXT0kpwMn/x4cSi7c8hNRAP03PXUMC8i/OeHKpa57dnGQZDvKD9JTIt
LHAFxbXBhmTRx9oE+YDcjtO6R6gGSe1dXrazUeW8ZlmgMf0D0JBfnegITx1Lq8/TvgkH3rNdtuda
tOTbJ4Wot/o2iM3eXRwuBPaF0qrahraHAykA8v9pXpWZg6v1siEvuAMc1tpri4lUZQGCWgJoT2ey
l1aFNnWJGaE2eqn89l69ep0XFvG4vERYJHOUdtWFR4gs/0Hpp8FZDbL9ubrEOiOEfhPmUM7hNkN3
/8YqL7BjyCY9YuGUWKPoMxaW/RWD6JQEp62hGEuDGmoAfcZeM7CKoYO+Zq3fl0eadsmblAvirvfb
hfff6bD+xE4oQ+QdcFyV/DDc40F381Dwk7mj+nSKqDmJF2dmai11igJO3t/aZCbra06SmOOkN7Zd
BmsDn7yZhe4YzU1CJohYbfHnC8wqi1DMt11eH74cqAvIGwmW70lyS3evyF/PUnuiboiw796ghKv8
Wo7xc0I8rJSTlG+2M0dQoWuZAvobRufDvCWoonZ/BKemf77aWP2uDdAfAmFE3sZD6ceWMgJ0QT0+
zVR3qmSriQP6Nuh0mWem2di0e07LfJmTbIFL/Sa+kpgSMNmAYe/jU2r1rWMYbClXR44xjR2PFmS6
SRlcAxscEvuWMXd1EeJM6p3vFWOxjVu7XQGUALv4WMvzLo25UHqQazj4pUf+KQPACBdHHdewydAT
xlRGrZ77b6FOt4qT2YE+RD8IfuCQEs8iFrUjKiUTitf8NklSRw0VaTl0edoYEwuR4MdXkc2FwNeu
oz/Zv0RusA2Hom4FVp06ALclax9zUk+ueRZSs+LIebGteafMw31LVvRpKAwgzzFFKdyGodSSuTM7
8ZlCrgXkYmEIxgIT7RGT+lwLQUkt5jDoTeKUOpZRXOolYs754uCEGhFR6ShideaJXGGfVAUcmzw3
gc6LEm7Miq6BIyXwUjD+QEYFYPq2neoIuo39ETD4LiIT71biwvmhFxL/f3cnWRAmvR4vJ0L5ZK/Q
/zFRIgm5/17Rgst+v2nUw2lHakkxjPrgCWOvvWKVMVo68fyZgsorz9AyGObRBOoMyvivEsWFg2gr
ffdtH4ceIBzUviH8Z0GnMoHhg2Kjo64K7sYWapeRoBBq2iaPOjvL1wJiM69b9DlFYmWA0JOBsHkZ
pPrbWWnB19N3pQ/fZM2yimcPNZhEEwUOwi9nczN/vScUpZAkr3U88nU5EjdRjDMMk+oIcwViDutg
X0QQmAjPy+8ctuz7aWRZIkMwxv8W5+Lgov41/7qDVwYkelOJ7CA1lt5kpK69CpIsK/lunhbUdaHM
F9hWo/vkiTOY9j/Pyb7pNfKvEsAt2AYGhgBJD3s8SNiCD6qhbWATe7CcG+RQD8rN8LD3LsgUEcUB
HQNdTICVeELQxhtBYJaJwFmq+ASVez1u0UDYpB0BlrsSqz1yzLw5D4ktcKDlaofJbgkk1lV3/Qw8
cfcvZQFIcjMep9ioDrXoRAfH4uFfMnt7mVYF7S6v7anI1P/iLBA7w3IO+QBmin7V1Q0RYmas4Uz9
tfT/vGlJb9A2wpGTNOjkvKu4xW6ubmbv4sXFRZWzDHHMZEIN3M4De+ArSRsL16I+nm7XhGR2LFcY
X5mf2cbSHQY6PjroDyvk7orAaJAI1d2IJhnUHChxsK31x3100ipyWbfZ0njcADwuA1qiVz61ZjCi
QBoB7fY4WrpBTvAqNZnN7CcwC51/DUu/Z1sDSB1pC+Dot8SBV9OqBfj15PMFpTWGruGVj583gsxY
WN154uvGcM3BZ2ZCHR0SVoDY5A2G28G5oq+CiCmUY7QorIbqxHeA9Ss3LrAnhuyUYd12AzbzR2es
bST6gn6tuV7FjSMBEQBQtBxwvic1CW5Z83nforwrr3rk12O523G9ToZtfAWr7UsfGuAexY2WdeHl
E60NCHZCtcP4QFo5EwxOHeweKcGL48hK0LkatOhYgjbfkaQ1bifhuGTmSwugfLkp0R6HXaXl+RzY
BIVEds23LSiUdHsRuhniXvRicCCEQ3IflzHjnHY5OujhM0BbrKD+hgECarGOj8fkRVCIjCO7G1gF
NUfr+00BFZ88dBQ4Cg+zs/O8kFEE2VUDCKp5TWORXa3wC7XSKuLn86gV5hv8R2k5gvTeoF+2IsnW
ZWN+ggB2Uaqv48qpyIS3Xn1/SI1HyC0hG+J7xE4xmkWlKU352dKxJtViCKoFej8VUzh+Jjgbc++8
qDhCBu/Y/w3ILhJIixvhAEBdu68Wc81DUwWz67ZKKZxvWftIbC3OVUieUgbfdXOIRUqNHtV04TRx
2nm5TzSyvKPr03KJdV7U6uTZCjPd0HKYU8VQFJpjG/TZiDmoUe45M0CpRMNy7QrdK9qcbpQTWX74
v4ZBRuWSEWCBtYzbZgWuFCQitf1Ui023mbSzvcE+WnFJ/PEhCqbRnqvh3Afuc/YXrCJl7UBJZKy+
RaZhTfTRGNxIWh0gIBXDZX5TLxFUaUdSUx+oWHFZZ6FMWWtiPgDRjCPgRnoYOTdteZbYmg1FacpI
5nph6646LsXG3SUHyTbLmw/b9TjkZnTkoiCMiqasvYeAmxQQyqqLu69G9AKOw7jUI0Nom4+2bjIF
4RDZqYcHEJ32+/xVZOOoWZK+i58KlVS/v7K4Ykuvk5AeM6171esiSJkvJmsjRM9MQVomYdoUMTJG
837jW0EEg9iPjN6SV8KOTreehOG3W9tAdRkF+W+GazdpPQSEeNO35rLmzdHCqRD+HAynExyPWeVP
ssG+F4bQvI4BBTYL7l1eeXvnKuZ0peBD2rd4oTYIrHvUrc2jw6Md1ZKB0wXAZ/W1LcQIpzWv5H1h
NIynfRmOB7PCwTiZyh0CGDsqPnPebpBUTl6/IYwOPNCEazZPPPINbace99twzyq5oJR8yIdukgwh
8xS5U8+Je6JaSCxVZd6to3Wf2+cREQECb2z3b2bDhnioZE8Lnd5qFrs7pQCG5ZEM7H94NfB7MHMM
7RAuUbGqLIUq2t1xkQ4VK8ImHeibGDFe19tayooGyO14TL0oTVrRjVBBt1y3Mub3fo8jPsvM4EXC
L8xZvLpr9CHKXGoH9cViCkqu1Fg3vidZeJT9W05jwXuag5HR1qhH3pkxTax6gh+G/b4iEdbd9B/3
ZeQ2Wx9DfjB0hmyDAu4AByjNHvtKAcnxyqNUzD1Tl/UG/7ZoCTXatD7Fs7oTpnikM9eKRNcndLrv
odYB+mUqZSZEUAC5gljeHhAOVVWdhxGFY/TK8U9+hpZkr5ys/6HppvKxbApaoLs+ddhbaa4M93Cs
jpL2cBqDAWLP8SVXwmRMyXUfMt8uZYiUoQisQCeaqOn7MBip1ScSfxlVRs+Du37hh8Us9a/O27Qd
qcCBTp+ZrsDr3mkUHEEkmR37JorUKkTg6+91R4klryvnpv9vBvJlX20Gewu9xnynhd0yI+eWaiiN
GPvT+rJnx462AURrG1bzWXlzYOqc6NieWyWckQpmozTN1IoaqiVht0/omXMBqE87SzNigD5AWhn8
J5I1XsPrJfxElCB9taohHTz2UqKWzRZ3agmRwNuzBwiRgG1/z2mhP76QG7WNQvcJGiCcm4nk42eS
YHailh45jysJGLCDw4ibUhCEFYtaGJIV4LhKCKJ5M9L/hcyDR2jmft390dVKDIXDMVe0pUx9myW9
5dZhe0Xd+zWWCC6hg27Lq1eG7Kx6pWaMVF/rsEmtNxpT8ZAc0lgHkXwL0ea9j7UYBZl7Tj0WsMGQ
cdXwbDNpdRPbVG5Winnt6igO8svA9WlmRhInDgcHn98iJVZURrozZ+zeRg+GHz9kJb92KwjuV9Uk
0p14i9JYFlhaF1qc2jH4DYnBoiD7YhMmxHZDThi0+rbhEBGrXwxuH440LI/LtiSGM6EloTJZ5nDC
c0QzTqUdlLjLMy4oa+Zz4rTGeIpRSsERUPs4NbgTQytUma0B1yW+hypSvYYKEtRzDn1M/zf7ZpeI
fNGD+KDo/taods7q4geoxO2wBBHp7XIZzUdp3g9Lltq3uUBOz6Ctz/G/b43/RuffLBplebX9PDZg
plkEqmADaWvC5tMZxYvqKJ1M/3eEYCvO5RNOrpejZwdS6lehOSGqrz3Kh/uHhQk/kKvHyQngCwKv
J6QYAflc3gs+23PC25m05HpNr0SVoucuB+XBw3ru3tgiOlDXp569SWgCi40eCMsggBLMQVv0VIMz
jYYjdSmjC8P0nswbNYi4s6NTeuB6CKdD5V3VMtupcADlEL6u0/wnA0iScrH6NMuz61ruFpmvgQpz
zq3jVASt+2UjVquoCB7dFoXo9urNLdsVr0tcGVPvj7thtdPDYceEGVHPPh2FAj1yIzpNwctZNRmL
uZ4Pjbc3aqy9Rahpp1Gn99IpxYldabGoNkWbn+KcK4HzLukJpIzmRSmo1o8VwuRGGjzGjZpphH6n
xA6DYrcexiODOZGNXlkYamz/S9vGKAX+bYvpLQ2Yk4zOi1VucvFutx8RT5C/irBtOxT1IBZQtIkM
ZQrbbJHv0vx2tLOjpYOaFZzSAjjWdolmy0mcs2mbzsuK+C3enmi1TSbuOpKtNydYTe2/zmUJiJfg
muAkF+ZZc/n/Zx+XFXKcJAr0PB6fZTjDeVtfZWh6fim+YBC/ymID17F8b7iMAPn78MuyYhvUiJ19
uc8xtPaoAzhJyKqqsiblUUYmkm9pr14bT1/DOCj6IqF05nAv9T1zUmD4tva+F6WTA7F0z5kNXeJs
DGGutdl536LX+WomRidN9GLQlcZm/L6+ck87raoIz55VlpNMtakuhkWYMiW+3+s6rb3MdiAw/Br+
oIEMKs6SPjnAIa5fhBLFvUvAKCd1+QTviSgRyZYKj2RWUJTUygmiScdV9E1tWSaATjiYNUuiYW8C
srJh685zHDTx/a6KKAFaWSpyzniEtwGRVbRzCp7f2Zfu4kzSKRQdsz9MMZ0mO80Jxp75J4Z864OM
ArgBXN4wU4NZ1bf4uOlfU7M/gAxe+n/azTa8CvpZarPi/UT+T8ncIJ9xEGARB1knShXYv51F1Kkk
J/qMI0jMdEqUL29lk0VR5RtsM83iosmnVZgDcLeq8qMmYXgVwVtnqSTjgNfhl8Rb5hENLPLnzDDC
MrN0GHyXAdYRHQFea3hr048zwsuqy2tXylP4++nPQW+OrZ6O7ZfdAIAKZuXkH/xKy2SJ9Paomm0i
Tw45m0aIo6hcZ/hAK+Lek9T1VlS8L/Sa5Wahj5yhEiOsm7DC2AtLtH37b/BQqrBlDeR4D3V3BMxp
Fg3OyYcwByDvMVLKKBU5BxyRe5uxAlrCtSiR05U7rHYDV/p7hGNbHLwOitjcDOEQob9ZnZlPx75+
8JhRCQvQUOMYzQ73gYyGj4uoZccB0kxvLoeBpJp1q//HnOTVqWdQH0PLMc6/55789eR4r1nEoBvC
h29RBecW2IJUC737f3yYsQzn0+2Glm7oXtWbSTwuIBLZhGihUq16BrnbRqw+xHNIjlzqGvbngsxw
jkWFXBOzCXxk5vcm6/aK72DDgK4VCLe9dKcTaOUyIAO9pVdPBhxVUHI4mtPaIVi0vByIfNFbAPY9
MLX268NX71/5dslfQfr1XGG9lHp8ssM+0bNKy8J2QT50vRnsw1IcN+zFMk3wm9rz7lTSjD67ahUq
y0Wtf1Z6VH/7GgIq8S6mIzvBQ0rmqMsGrBuQwsxkkhzhzTgOE02g5apUZE/sQS3Jr6uALF/sSY1O
ea4atooUJOn0N/dkF6LprlJt+OZGnh5MgkWvNbyTUxvFvAQjwOOGm0MpdJRhwzcfuXnzO8RLrRdu
0H5k+nDvCgtdl0/W/sFc5rPQGIG8tSBib9Khs5q7PCrX53DSSjWNSb/18ilHIH/N0kBAD9NHTa8N
MgLgGgu5D4pI32Yn5W3NCVVGteb8Z9PhsbAjob6kP/dBk5epi9ftKvHPzA1KrZ+BQyyPtRWusp+3
tKE/1lkjNx4yF2ER/PRSta2XnOWGS5Vvpny9SGkDfVIK+UVGbQNS7keOxjd2DYYRwg3MPLrrcM9X
o9u7K80BwCAYKOmx4svX/Oy/AVMZPtj8ukG8uZF0Bt0eyNH15NFzr+hcGJ9iE4OBIEXbMv7vwXVj
2mzdM5QNKyvEB2zf2G7ujZxp3x6EnCxqBYBeEgNY3w8ZhlPbikCvmECSj/V5VU0VqDVUNbjV1Y1X
EqxvtopBBKRga+J0Y/ib6izOC/5C8/o8FCaHlSpbltqVmuZKOJM2bADC7kErDGRY8udFBlyDV0ie
J5AWRVZummIIuL334178vLKMOmdzQWIDHtDaDGDcjzd+lbEMfNm6BiDFsL3ytoj5W8+1mcWgyajt
GNzEocumhna3IdukkVo02p/G7idOLNfGDgr+oYE9VGMB0oqlJqxx6WzO4YKGGlXTYoo/84kwT2pX
g4jJPLfvue7UJ0nPfBUEcpV49ZrCdcCLYa+2yZPyqrKzLZ8aJqqlcgbE/3sOQhEH2VMHiANMcx1/
rL3nDw+7tNZf/tiehAVzWgNSs1oVxRnvlhUqrm/GFAGI7709Hr1YPUtrtqvDuP9P4ZjUSa2zbyeR
v8ThmG3OtVXY5MY0ljwLSJ4/KNCuIOkdFZ/ScnQLuRQ5MwZx6nIqmCvVARMsZPFf2aJX++iOMDJB
IBHaQ5CIQu7WeEuB2T46fObgPukHt6hKURg7bzfOsj4Yv+m9252rh3X0Zs1efdS/oXRAPohe2CIf
lwmpV8A3ojf9TQDZOQv6dlJkHGsTlhqv3Y7XP82gcWU3uQLtmJFRFUClMXUCdow5gr6vP0RdirZC
mdAy09I4s+HSFYiOPpwZUTWWfytVMYUyS5LB0l0KbiZ7HDB19vG2KrP3ltg57hZdUS1b+EE3rKRX
VsVBo2/LvsS4twySIpLbVSZT8wIou8OjboIUGV8BvpEDCcqDiOIrNVk0I5ut1PyDKAEduaaWSy/f
bzOCwswkip+6gTZubBmSBNOkXiVVTyMji4WlNN/lmV3IV6quGZsK2wwwu4HlzHa3M2sNbRD1xvJg
HCZr6DLtW/1e0UtX0a4m4ppWS5FrCLHXQteJ5n8N8isJIiCZpKQnaFPvpCuqQzcGeKV4MRyGj1sb
5n8Kdd4QK2pZFHkaH2ea+K5KlSesDFo8kjVyI6SaOKsdVXXrsGBSfg4xaBY8zH9vlaGZ7vzQYRG8
oMt6yg75GAI3vwq3VerNWJtM1SC2Vqw7PINbI+Kz3UcQv7J7jhAZhVDLVQ6Yi9eMqPL9e1SI1pEJ
TXbPj+MfWkKzjbMGTAYV9liOw1SP5lsJ1d2dEoJT1lTAW6EAXlgrP+syHM2Ia3Vt1nUhyRmnRkRH
ZYvZVzz93SyZ96JMHPJfDx05dFVEPWRmnuL13MHMZPXzxYYrhIyUeJ/1RpYCFlzM9N83DD1O0t7m
YECxjvnxgg/eLe4+RIHf4fA5LF1X3TNH6bXs1i979h1zCpTQ2K3eE+nD9+Q10uf6GW2ZS8LbRRzf
Nl29k7kuLRy2e4iYtPk1ClOiTY36fkDygm8RbQ2pYQvYiXIrKU+j9aBDdT4FgEsXaj/WsU+s6kCd
ERM4xvI526w6d+oO4wYYPJMURXiBkz2aUKdB+eGZ9c+87P18TSA0bKSlrqYs5eXyESZ8fNg3dVnA
ZaPu9rqN35FZG1hL2O7AAIJV2aXuYwkow0Gp1VRG8bzRkl72Iiwupd9B9bv4UNfAEK/O/WQJeUI4
8AJjBtNu4ESIJqEQXOLOv33Cv+eAJpz48DSJ1DnML3wJC9sX3ZGMcN8qDIV4GrGfe3jL7/V4Ph/s
/jQfPst7m7HSO4B831OijRAEh4Mn9XK3pvH/r8N8D/mR5LgIsI6UQU0TQEfN8Akqj9SNrOkfqL3s
GTxDyNUux8a2JFDU9JHDUWG0yT5wINp3+swNr9duimgTK3ng3WpOiBGzfWIFvOGFs+7O7QM0VL8k
jX8E682jIRNZjICt3lgT2INwi0fwV+8bouFwpOzuQKVcRKH1BsOfIhobLaPpvxiZU0tcAKnU/tLn
NE6nYYXwB7KsHIrBaSO2yzRox2FRt5gEdsSWA2TyVHm/lk55ACYPSDFxKzF03O+9uMDuGEc0CzvW
1IbSROG1jyydY242K4+UriZUUGaZhzY16p1nFqkvspgLBE3zaV+fikBwKXhYzDDfCOqPzRYSB2Si
XpV+V2FpxaPy9nKsJZszla9Klwejq0DlUNVaiZASDkKuwAuqtN28TvHzKccgD2mXhf3xtFLmMMlv
OpfeAqNjfWYtwCIreq/4ZyXJRHbp0JoLvzjvP1zFT8PewtaOt9e/YRjlpA7MkbGN7JKvaMVnI6gB
yyB3tcQDUve2SLyHf/9ezXmjmoEd7XQQSGX8IJ323DRyBbQDQCXlPIghc/m7y84MH2tFMYhZIGgZ
SozDez0YJ0lyCiAvUvhdR5p25QkeEFhlyOP3SwOTIK9KitzDOUEgg2aeNoc/FCG3OTlYsBeGhfWU
TxEpFl2APHRSxgTzRrtmn41G9A9tO3GEOm0f9zYA3lzL1FZBKCb+L7Z3gOOtEzpWAE2ihgHw7siQ
RMfZf1UMHH03RZ1y+ajIRbYwCTEMRlQCE5RRMnFOCXABu3Y8zACZo5L3oMGeBDCFVC/uN5s7YkA9
Mpmgot6h3jTuGAC0XU1jxnuI0z3UdJLkgUD6ZTgJkAgbHTWWqhYqN8bIt0tyOX0r8l5UdFFfQ2DJ
2oWMRfmpS2PyP0aX6SmywX0/nfhzEBpris0W9Fu/5/lzTxqOXmOO4g1tGcRaDZes0Ryaf1SL8z5V
ucz+7BfTpd6bsZcJj8ZqzWjffrkc4g//Bv2IjATCXm0HUtP6APRDY1cJI24cCBiuqmYJS0Z6uwp1
hK3LbtH8O9WfyYXurBFtXtzm7TQjdP0tjSlwc9poYDloY3CcAP95rSpCGc//7VY+LnAmsKV4zCMS
YpdoIQrMsoeRUJk8AHsmutHFNRshREBkmrdFRFHCLPP+inyNZ04jTrN+3HBv7Y/cxs3IGRKf3xm9
fHfhAqTCby57O527ne/ks3dHR1wZ/W/bukfHJ71Y1kOS1reD4y9qs7dLvz1R3E6XyjnCkpfh1Eyd
rIIttzWgBJ5ojwHqte0WgAOEXqYU8meukFWXuOUqzoQePRQLH8bCdDXJCK0BEAafImt64SwRa9jD
uywl1OrrsEjy98XNyCB8S3+Qia4soFZbUuYJM6Ui4cond+EBip+iHza/nTqCnxz6eacrOIzVVbp7
0cuj5mIJFvKa0bEODT5xCjQw8Ph6s9SyQ84Bi8oaVY3LSCTY4da9I6Tqdf/XQ8n1r1c+OkazgIiP
lCYJpLji3eMGlmCJd9r4393Se7TZeV4VOjQtZMcvmvbVYC0hQ9xOP4o5pngAUxN3JHqFxXzLhlyK
EOjyM/jcFXi9VpS4z388A47frvQrIRsIUL7BecA+WwTO+aeFB2vLBdv27yqmafUCDv5KSwDcnbbF
d6V5HcJ1u8oyiZYwNkc8NgFoJ/nPiUergvKQnp/SxZ17vvaE3QSftRP58iWzXN4TjOMOnmir9orq
Jg7xSilRpl6hcazHcDp5QEWqxC8cJCaOslf7ejsGhZa2rhiBIB67Ip531mqSvWaC9a/jlA3Y7nJB
MJCNtqQtPg5B5CrM9+7ZrBIhxjMpomW257Y/KDhrY0MIoi5XXYTQDveF1M4txEdYLQd3j350DpkI
KdPaykIyeGk2oinVv2RD1rfqYPx1jZDtOZ73sKWsXODedSqHlh6dvhnSkfUY9ibUFdKeAa+FXRIP
HFimVRJnjjYs7gFknNALfrwMcpvfu5TsS2k0XxD8umkbiNL2Kc+s/v+T2snmecqyVE1vj43TlkN5
8Kg2rdC/wGlIKctowdnEDwdL4Yt08ywtvaCbvkyNmNxxXwAjZQ8K1AV7KtptAD3i+TnsxRXiSUNM
/NEDJ6NAahjiDZ790diYAnQP5JszaP9oL5tYtCxSMYLuc9S4uPwaJO164por+9kGPEBkDe93CVKv
6H9Yy9SFDtgEiUwpqmqcnFSkGdnOh6rHbBXqfsq05I3PAwd7HuMa3Ce976B13dQ58ZydJt078WDn
M7jusMtjpABIlbu62Uyms3iyRwTHGFgM1Wj2iy28aa96Fbl6kiDkb4oqaYh3+am3gBrv/86eEbDC
2q65LqRWw+rUxitA+HtDo/okEoJuWHPc75VFmSom0im6+zeQeS3HxVfQT0biIiG/sO0qLRosR383
BScREXrT87LYeKBAXdY1vKtqrBXy7Cu8wK+awjlLw4yywMxSgmjP5ADrWeN7qflJZfptniBykAH1
stdK2mjUjj3l31EQ5QRfv1LGCzpp6IwbtS8gFyYOmBlRm2EFLGlBhgBCpD/PXz4859TeZmAJujsG
LwW/zeJXxTKUJccB9jrvuTWDAP81N6VioWnMMlKUC7Ffuc6/rR5g5MzH/u1lmxSYj0LHWRaft5Xm
usJcxeIr1VYIyLLth4VJQNfimnQ5W/U3RuGeKgQa13BVU0kTrwZgSsUNHyZ0NlSKoCMiwxbVf0p9
md2n/CUsrMknP+V/j/Impfp5YvzSnlpaXC4v01PLoqkFHWT1JnDL0zzr+5UOKyJq6RfGtRNESB0i
iliuHzxCfK08FhQrvEeLLpmLVfQGd7khEBxdjWgVAwgWy0NJdRijiNTJy/VXe9Mm51e/4+uXyfLC
qTlUkNcePl1cDIQtVmJcDwcIVcs+vH1dcXqRQvI/6L49JlP20wufE/dhwzcbXLh51Uygr8NNQmrs
JXobUpsGnZnApTcZdt98dUUn4RljNw54zvuRwU56D/jeIuSbwey0PpG6n8XHD5io7/5DS4NeGuoW
bdXnL5eWeZ4paMhH36t3C+NYJedyriKGyZZGgAogqTWKsV4+zuBS/HyA0ZrVvddB/HSyx8X46mcn
EtRFZ3rW/aRWdpVSA9fcz8Myeh2bNfKIg5HFxK+86aVxKTTLiBWYhSCrsYWXuCVUvDzdQ66K2Ajv
bONNkV9TA9fBr9A0OnoT385s8MKpNIiozVs6avLZ5QlTzQS6WkdrZ4Pc48aT23mQ/WnBnJSLntsB
5FoYzBxsKvw/RUOzUtOLkNw2Qlz2EqOIRaUV/pggAuOxCA8EkjPqOvXvjCcyZZaSx0meIqgXFc0g
KzoOJ1wRQyfGE+eUCU4ddg4toeh0+Ii8K2Gu8OLr+ME1uNzIElqo7qIkshMbSFpOETdZKgoRyEi6
ODsu3rc3SU/kUbtnYwanmWdZW9fLyuvddlaCFYYmrpt/F2xt34sPRzHu301jItJOYWnf0pArmejI
BgUmeIsUNHXvMEZTwi8IW+uCaGRSFuFWm6+GC4ZVZxHN5UPVfAxKn4XWNhFqRh4O3uAFs4fGBWdW
YZeSFiTMwO4iUkXCqERtL5em8sRNQO8esqwyFJ9gJUf9f6r53i1IJ6ptVS84c92xSAPfUL6Sb3rk
ZcOgn3o59Ru2KhmxoBSODVDD1d9w3JFVg09NeGudkvnEcTUVitVneHuO36I2vYF41qttdc9UxNf/
cpgnLGEj6Xt9MWMFXuBSAlMtDeu+uPy9ZZPSgB2YgMJU9Jp2RtjjZHoXJoEuxwC49eSwm6f7fRMx
U0mmn9NH3dhinQQuYbheW5tDw0SYwetiWj6LRF1qdwe06o11M1d5W8k1dpjwcmolUrGrQm8Jn7rg
qym24C1HUOdwoBU1zW84LEUNh/WAH7lJUJwh8FeSTZGFD8hVyHj67CgCaHy/4scCLTa3tkizL1n7
CYDe0lMaDiCRwqctn/u6f1zrk6/kv1inIdY3a+CH4yCSF4CYoQzOjalDZH1uTYo0yyNwj63K/w3R
EG+Fm8LkR+sWh86rE4vQkk74VNbWJr7K4ryka1lb787E14y8/C4MnmZFCfkJxHutpiELZsLTL2Sp
YUpaTwntbCYSOeg1nZhp7fVYL2K4MtzhncISxOTh8AERpyXzCI/kVZ8GgYIka9WfI9UFVTloL4cc
aE6rnBIhxOwWP0b8zzsiR0ok+umrsThMjdkrc0g0hf+MVh+WyGS8ufDzIkl801bEiNNuI0+TY16y
P7HOztHJRmO4y+PcHlEFF44Bv/nDIyXZe+X9g2GBsXh5CERoe3ngB8fE4Bn24gs/6zmorQnDRQpS
3Qdr9UiHMubcZm/hAU9Lg4ZOe2niKp+alJgdbXUAF6r9cyDXFzeKK1icuWPYRfIcfku7KRBfLsgx
+u8/6Olpv3yEFZGzcXGv9qcorkJd9+hbFVEYiVNw9Fxm64p1sLkrkcu8+ek/+fVdivEKNBuPDyom
+qrVA3M4Nw+Atg6SGMyLFp2kOeg+SX2FFfvIyq+vrqyYexOCh2EKeFly/Vs8ADPMxr5zy7aDmP/Q
fujViN0D6+1qSsjwk0rBRWJvhTUoQl9/hbXT8okBFwLt/nz+nMMmkO8ehDRLn9r3cyUQcCb/fGEm
3bdWUwFjZo6JoxC/PnRcZenB08tkSnJZ+XxaC8oIxKe03MejVvbJnLPzKdQSvvcF6JY/zUCHCpSA
k9nc5cC408rJvjXQ/+Ok7j5/wW0HCTG86+03lhpl0gOFYqrF5spc/vih42UQBUTz1zbDP9WDSz3U
fb8mfOHlpbRTNdNUYTlVS9JcqtUi2M19UtHHsDVC8z5AFgiPZjLd4ZSwK3KLQYSkVdGZO1jW8V1V
Gs+Qej5p7KhtBNgkEVQuTap28NFRuoG+QIT+wn6/ZwCconoimozbHhh+9gPkHSOZFq59o1kvE+bG
W8o5Yfx2SR6M8IcNRq3zJfHaVezskohkxoYACG89w9Ek6wr2isFb58b+1pkVwGnfTJ/SWTdB42NW
Pi71HSpsJepccovjsyuAwU6bQr7O6GwWfyoKXZFdOMyAixZKXrLrUaT9oS5FLcpevmo/Riv0VIVH
dUHGFqgQUkqVmJ5sZzYSfT0/ptTOuXXbDOc6ACnEtMDVA58/KAiBhKrDxtnsWIckrrrcWSrabDFC
5D2XwIc2HrrrcNmKb+zHuvxjHhZqIiMme23eYCnSq+mbByz6QLsIWW4coMu3hISgy7zgnteI9Crj
5BOC5wmQFqlrhOsJcoWdrmr8QlOjV4AE7U43I82hnBgH9n4T9Mu5Y8S8PUnLyWLHjMT/TzNYjxTo
/DSptJ2+F++au7RlveSc1wEIftwUUFUMXFmpHSFYjALC0qTrS5ZmN1QdfUfeNm2XdpYJ2krGbBaG
dBwLaxkzxnn2OjULKzvPH+dYz12E5QcHAUS5bt6atPgUlAWDAton5gzJ+7AxPg4C2hai6Vr1A+V9
eUW8pp0cEoa9O/ryWOudN7rWQSjetU20N1hYJNdNbvwlzCHd5yYwDbdNInI80VK9U74LtxhmMMrr
DKLQo3THQo3XfTNUIEDZR9psJSVfIxRo7h7q7ob3h1cguweWLTRbF42I1+6OwhV/sr/drcwAP4wO
m/Xhn2Clf5ExEZoYrmq8xvPdE2uZwhUPB+n/ecp0WTcnDisJLAjhIde5SjgATc06rr32O59kObms
WG8EqkEi2KHmtlRjgaKVN6L4zNi6kZEb1NibpcIozjICFdR8bdVJY0K9yQ8skVUX+ELOO3N9HIKw
BY1dBbmE9hvD8udnJrc5TOvh9VQSg64Fre7KwdQIAvZKjW7crXSOkcQ2CXh/llRq8NqM0hhXs2Jz
6Cfmf9/+OVWW2Df3Umk6yExB2/tdoOEFwKnVDk7ULjfrB2LqFkwoYW1Ys3Le9OmP6e7SU6tsR3Jy
esrBGpf0HgaGGfMnTTF7MlgW3e93OZ12g9mbsZX7Q/ye2SmOnNbfWhfiizQzbfrDeM63YJOpLeaG
AmGQN0Y3PF0Nkc3y27Ad4tq9Lpy9uvMnbhigk/53K6Ged/9lDz1tExjDdWaCPvcxH6vMg00pUyYq
GNez1wIo4OfSvJfoi+WcRPjFuI4AaO+80vNLosszgAf8sXdFMzIutIeN5kO6YO43Jtbgfm8Nqou0
L8rYeTxnxsrCjPvM5DDqC4jbEJhsR196NoI2WuH7CLudny1Pa2AT/d/ow7L8zZ8QU7IKGSRjNbks
0j0XOJIZI/Q6YzZCNLvR09Teqlh6wXTK7B5lQR1cAsSnDAFcZnsqKjdseGxUiZtQDJWknYP/oIqt
4QMJjyJgSK9V0DG8D71XygoK+R4ue3bV4yVbjN6eqBuG13injfD8fo/udvTRuIn21e+yneG9BeHt
U1kvf+2n9H7m4YNOmEOdX9yI7QaHiTv+ooSMnLih9v2t3t47zx/dzpB/XEp1BI8WgpzkQKBbPI77
RBXZr6WF7bKzqKjXDCFNkdKDPoIk4l3+epUx04HZ9EZmNXuvvpwGw4wlONmW9cO7rMnrIpugAc+t
yyHI+YQmIIYeK0LRZ3qeFvkC0xiIuLIAybh4z3Xbxy1erPjRNuDUeQNP1ngXPl17muzYdX8zFwGk
ovl7mipA224m4W6qusDTTr8d9kQyWjITWZRGxjDRCWd3ukoqWpVoqXOuJlPg7E62Rm27CVOZ+WtX
RjtOimXyp8rtBoScCIEVQAYI3I8812BjV7por8UGB2K4pN3bCKPU4Pog860+2Q4KEcHUfUX7bpa3
F34NCotmFVk6rXpAzyXeqpxAGci4zky6E8ztVvZWCEyqmklFhIN43krZ8e/15IX+inTtMiafnAgU
cExPHpLLKuu2+9sX0YlCOfHua2EBAx5bcDTZJSMV7leZWyEo/8zxoBYUDyyLYTBEEi5Kd87F0go1
Sh99FC+nhMrq1PrekvOYoROUJ1jNA5Z65ptlopz8Q5q5CfeseO+xQe380FMqAQeryL6I8nju18zo
MWXg/VaRHSNNVIqepf4tFIkONfUiYUXiWmB/8qzZUch3sHTUo6IuBBbYHKcSrLwAqqx7SUlpSsFU
nYrx+qsixek3Kv94bmQBdds4V+p4xwQ1lShleu0WwL2ZcpKDMe1W3uKxmZENssXTu4mZAEXdoAiN
8+BZ/WG7zoTXZTYSQFT5wjwIycCd57IuhdQgNTy8DEC9bg0Jj305DshcPJz9cKHHeaLL1nvxhEC5
6XpqwGFEYPlYctAcz4IvWEKmG6PtKw8Hi8BJhMe548/d7w2izF/s+LbgXqsv3W9TiOsjmDUAejRy
vaWOVpsJ2mJDcWwDILOL6QxAnjEUfgzflkB4IAuG3F3sPQ40s/kcAdxPkgZJDCKUnnpTR3ILrApB
8EvZMx4vdKvuOWSvndWJGEYEv5I6e/fTbs4Y1z2pAQoYzm5Gn0ZIy3OuYjWh6wjUwTMGiJn9t/zw
fwGVhbUfmHwXjeLMlFHJTgXsNPWqLGPke6Dn3jqBhrCFKmhMH+8RUIgaIUJomaSuTBxM2a09FHEe
ehDRhaelNL4SSTiKQ0bqxdAGZzTmrbgeMzBkuoYn5vLWn5KGEfHHN3mmX6y2SIEuOP41PZTDSNor
w60HOwCie2MehT/sY9kxe0qmr7ie+G333/75aWZBFcWemvqxrKmHTNukhXZki2/+Ks9+ypZQmKjA
BuuvKBNK1Ax9jJrYZx8wmvx/9FGBHJ99RzoZdHP3lNZs+Wnw0tsDDwJuI6YX0HcHHlvMUEYANsk4
8d94AclRu3Dcz4PHENgCqdDuAPULUouvccrpNvTwelKFcY7JNwCBu0KWsoveKKhgJIL0X3lvbByR
btDblvpA5QZqt1j4OVBTRDxDj2+iQf37amirAxeUFH8oMhff1AUjP9UBEBA5wOfaoxDTqx4DG5TW
f3DVNodXoEeY4q1430LRzgyQFQVvms7qjzN9UypR+40hTObeRul+3AbOEQL84ONVV2yH7rrtbHHp
PSFGN22bSln+km/RadKplzb2rFfc/LmWbMZIwYpsC72bGtYfXPLglTFBrt9NwTpijAsmm01Y8FRS
BdxI3ndvy53PnsKKNrovka0trS67uPVIzbPg1rD5lDhi9UOHNflN4ZfCMkLkZNFCQa2aTc20SAhF
yHajK8ZVw1mcf0s1FSUqKUJG2ax+vIMPDOuaw6QZT1x5vlNSMf+JjM6pWylFv1LzPRcVmuQbGl36
+pyQG60qX2ZcIGXrmZ6KiEhOrLULcLWXdF2b3JTixaue+zZrx8S8PRoSSb3zyOg1sim6qKdG/pCg
8cf3i6dMz9m9GucXOAd4YeTOL4+ZnWBSWrTIK42eNIf2gJZLJfoBy8epXtaSDsHJM4now7Hn7XtI
BxF8WPdTPQO7I1jCCBdfQ5joCEsLI+sk4AxV+uQRxTeiD6pQgnSxcORk1aH4JIBXxH4IPYEDCgNs
MG+LFRfAcBQwkcG61XdvKfinLJxTLAbUJp+RfmvhxTLkdi4qb4/vW3plrr2uYp0kF86PDQpz4DWP
NN0Iq52pYAa40bCgqTghH8xJahfUaRMYA/86gtfn6z5S/b5e0A6CPpW+f1TH+1EcccPRdO7XBRmB
TWP+fNp1hASdnCUjxNj99idgsPjMGfJjjbhlezCrnNEGcunriNCkOBOsp+diKeVK6AboIflQLbZ7
2C7JOFi5mCHtsDB3A4WEPyeoeWJjP2HLNo+I86hHfbpvFt02kBj719zsWnQTsHBnDIoYikCzPAS4
56PqfAvfxbtW3c95WQBFYb/j7fr3C0CtUW/6bCE+a/u3kqxVyDoCWG3uXxRvkJ3Ku5uqlNa5haKx
5Lq1lwl1hyHGQopzbKu0uIT5G9xWzZUrPh/2RJCDXXinbaPhAWhzdK0O71hOExf77P5/qoW1bus2
C3EMrKfwrGDhtkpLtuBr8abXajA0k2QFdg5OdsLAmjnINCUmV8XFJEJGKlvZxzN2LqtVchp0YMcD
SQPb9kWJFjhXc6HVpQ6gPprzNbb5qps/kXK7Qrxp/klz7v3V0I9LASDsovksYkg8AppAfZWjUEJv
vpYF4ZaXECI2ELFX5ZCskcxxvrwWUH3IKF9vqcNDM9Rxp+X/cHINUowthLn41Uoi/8v3fJ5/82kM
kvDnjApFl+vFDUzwauQtlrm6Bzbk4OxXULzPVrNGxzUEd+Tj5Adxj322fRQ5E3SL3WsnPICFtJCf
971PysQuWYmOP6r+r1gGjk4CX6pHp2J1bI6Jfj45JYeMZFA3lJv6dBmKTRjbdmZ4QhnSgXyzqpNR
RrdGpsAyV6VQjLb5g9/voOXtvccT4HYOnxFc7egKa5N+jPqc6h0bMl/meVzvuVGtY3LZoOEmGxBe
H2wpBG+nxC5gpPh4li3cmvDpe6l3EhDUhnMjuzgjvuCEyVdcMt3EdHix4MNlZzi5Y/K5VojKJlSj
BOaBjHqkXYImJO4SBfpqGQ5WfT3suXk2YR5MY/mtI6WtOvlmTLnypv/zwh5cYKdYgL3UcEt1x4OZ
ZVuCP0YI4q70+FUnVCLCIv04cFYXQJvGSJMJblFuNyNq6vQ36OIQmzHmRXhAqPWqPdHOsejKQ+gE
8nBkT53LCsmkS0Nh+lQe1J+k4r6Spru+hojkKME7BwggwyyjXfzH8HYrjU970wxmXWY6x3+tPcL4
wgjACZcNoxUu+iEqqzabpqTne9vBHFglPutF24TqwJYxiWS4zvQUFgDM3pzqvblYAeiXFn/HRBlo
r+lZV1BJ0VwrwzG7u1LqEmYgr7yt/Iwqiv7VBFNqgkehJFikEeVgl9WCcB3pld4NCcFCuyjYDUbq
WXHpN4sIUhcJHTFLTMCLpygulMMJJw+TM4SPvkVmSlTav89IBbZLVS8Jnv0K9Mh79jZPWZYiBY5x
Az3XxeYz2rZ1CnHEr2d7IL7cFIIYcj9RF0Qz7SheVSfuVHZcnKgZireAYR07hIaqt9jY3zq7H9qM
86QuecUTwzl4ZQ1beGdUPXbXKTi+1VKGWThQidomGGezpLgsCno/n6ps9zPZ0ob1SmQo548pBWnA
mMCYXKF5ObobbSDN65EqoMflQniavrthL8J99l90D+UcP8DpcnZi5ubeGZFiXgJb59i3lgg8TcB+
i3Yedp+G5uzF36m848pTi4IB70r+E8JykUHYkxEN9h/v+/KpLHZt54/P6eWWwl3ydT/InejOGzWI
hAUJwq12YFvJndHcxAuXMvMUgCNWx5XJrpNe+l9+O0+LPMYjbzH5EaBmJ/SgOIhfsnvTUfTXpd78
5b0lHazIQ+CVAWq/P9E2dut0WWKNPBX6MM21PaTlPqd60xxb2/+JlzdGSARrCNvFU4Vz9ITTNJvG
kFPv3oJxPLWp1/VaGu0JIwMbmrOa7L3E3fESbKFVJ6zSqvfYEfRtp3g7hIcMkneRafx922SAw8Gs
xlHDRhn4UMDN79dli9mOBlqVeKEm1TpkBB1rKiSOMPOMMIion3aKXa3X7X87nV8pEyUjaeMhsEhW
NWNm+8+J9j97O8+RB5lCIxMpjNR2GV5EONy8Zqoo9PnoUmnncoyjNbMVamYc5ebv3cG+LY7C644q
D3rFqgKeJQWJ/R3NEPkO7FsF/zDDWKuQzGltWy9GYkOMPxBalwn81Txj3OD+tfy+nlb+nNjCmMv2
txbDhyFGEgagxLSA7FnN5eYP/u6aJPQyfgZn4LVov6sgjFtSvFPyM6uDDvja83YMi9mxxVbfQsyN
grjvZK4kLn2prLczZ3CE4hUa5AmAfTyarmruzzW6Skz1cFPGEpx8MJzKCMzGYClhQofAykzHAM4J
NpxKGsEN8eC2FhzGQ6yS5vbLekP5sIx3wzGDq6zoLvOmTRlYkhjObf2qWEHNDV7EHoG4e+BmWSeH
Zd/qZydEaN1+WqHmaqXr7onFnEwjCe7omKj05etARtD6fi5OZbiy+z+6IA+1f9Uy2lW8N8+k0tzt
6yeunWE6iPyyFwZnI0cLdO4BlwgEoF2SKN/wKXMx4mpFhooHKXSjZEiSaULaieBvE7FThnG40R4e
tpPn9KRYOx4j3LRvjsMUINT0bQldjTu7RDL/CTLYdFtNMikhKEEFFKrnDUD4wnDT0uHsu5V0b5Z5
ha7KLy+Hlsl6opVIMmPWFnFb0ydBY5J7kPuPvwfsAVuIX+/iKG9GHWaqp6do3BxpRYMMwiwQXM6+
xsc+qIuW6exnJpxtet9ABf2xav5dnZnfGM23xe20gNdMrzU7DhEBaHo15jUzEvimkDN/EaEuCcZe
ehUycTU7NQHLyUGFO2kp9fFf0DBIHDxHciQ866Elohw7cEKdIR+f+dVVFJq4Nd8QYlzPuASJ1R9/
p6XlHod4/OUx8qXPRomcpnSHOy7eD+nAoBnRUy12PjMbJQa6j5wx7VM+sbydIfq3k4SouZ4DR4EX
EZCBvgN9HSod2RgMuOyVmx4f9pT3R6SoUEie+ihvFIGLZPQBFwD9E+CBU6Qlgc7sSbY099amjNpb
NfW2tT8cxsZZyOoiOFGi0AkQd3tiD+tiZxxNQftTDVUX4sW/qNSSxgjqr8VM0TBh7MciU6xqs4fn
jVCwN1l7RSyAH1CSFKP++k+OLBh/f+cnHgRALTGe3vWYN2V609A3Ju+G/cnPi6R3pQOR6b9mtKFY
yre14Gv/eDHeZv04KYn14X48elgHC/n/JS1vQU3ZUJKuTwsMaLPz1YNKZZi7FLmNCzwldwUQIX/m
5tZre4K2tWQ/x72XvV22Ja+CvK5hIWwYMHJzCns2hYbKKZNNk3EVUCorFcr4mVSmUnn+0e40tdtS
w2YMWQvyZMUTnpmrXgVzaXaLhakRp3q457SDcr5DzDqtbDMN87YiosnggOr8u+05UwS+SGfRTLuC
zXktFo/tfCM4Jj8gZkObN9rotibItx+mCpzN8P3nmlNuNwB8Sj0/49ef06E4YU41SeXbYi7aeb1/
EAajTe+TJ/PUufVlRMT96cMJEjtzsLwEYZFPMxmV6PIDP0LW4+0iqCvTqkon1TKwLAJvsloWjwRh
vyvXkAgr+SJlVDc+b8dUxdD/munoQ2iooEf4MvlIia5TwM7Ayf38voWBe8mU1/MCTgxwmGWoTjYL
VG+sY02Kuz8d2BNHDZCAj2H9Y+xwQrCed2UsEez9J9DoeHXd3QRDmt3wgZEf99BfqpTsc+O4qdLh
prh6vjxuNddzXwx+E8toQZDUblgwc4HNtRUfu8VUUCY8PhSS2fmv29SzvpV3BD3pAlNEL36xmGQN
Z2sJXXutFHDPAgSHvJc+LxBbMLw/YZjiRmYETDhaEAw2fxg3qlxxOdm1BXqRotPylk8/M64l9b1x
XWQLqZ9SpLN/zwXZH8GxzdIhjNJs2z5AQK2jYc13D1kB9J2xxStWo880r3r5j5Kd6J1Z5EcZ0rsA
8K1L+vXXv5k/2XEqXfShbNXYOtQxRSkV9v1CMaj+c4911x4BmB/2wvRKwm+6fBfGVRQ6uYU+gx+n
MJtpTuqVeJVuu97HFZBOk9MztmQq4r/fn40vVOyaiw1S+Hns/rN3ALGkihFaxncRVHDBWqRt2d12
vz4b8F0BbFAgzHgJbLd2MBEIEknCy8DN9mtRT8QL1s2XvIAPos0yv95Kml4Ivr1zI3hKYrko0WPM
0PJCmN2YFFhs/RRehjzjzvwpdWtqOtTldLNkk98UbSkooQy72Vnx7HXRRIOqY87O0r/WofeKs1e/
hNAQveeHwD5qH1eNH+e5zm7QHPIr6DmYIfaa5d+6dREhMI6Y9tZIQiQQOoVgnmCyab5VkqE6tvOV
TE2rGmYTIBXa49O4Kef2XcRppF7fXGtQ91kLpFEh8z7ROM6MRX0+mOs5U5Hfi7jBTxs+mc84fJDj
A7+S5zTiW/aya0IPjSsbA9sxGfQRF3xMLSpHug6kNoe5LdiTrFdkeoD8A9xGNLNxrRtPcU0fg4dg
qKVwe/8AbpUx75k8RQXNTC5XRG/9btcD97f+L6Hp/tXvubjJSP6fQ4A7FlulgHwepnjrW3Z6/uka
4xJNYothXNzF9tCY4vV5JQgMGW5aVZ4UP0LmapXg9rAqxlo7c5sNkZoT/fGsxgqyCMvKL5o1EdMx
ZdgkIH0E0Mz+nJTGuQZ5a3s4vQKY3bW1+If7tApcVu8K7hRVOX/4JEjR6vNN9UTrwrqBpEbs0F0G
QqIg2WNvZHh+dY+57neT1mC5xFYLT/F0eyiIzkPUe9CLiuHOZR6xP3lhFlkdI5YsburyGZquphKZ
pVLsQo0pZcpwYkkCFj9VV1Wh7lQa0kgpA+utWkoJ0hP6S1vmmMQQOe4oPABCQU/xzEIkTc32hzfz
eD6NEhHd2cdqu65cVr9qYDlqiECaqQKqpktl9JVqoEJ0ZdSBICEFrydJc340R6KKmIQW5010mKXy
daVJMhjjf/uT60yp4C1ubmW1y0zTg1isaLBXFoYNy3XK87q2XQjLjugDbD2c7NL4sOztnOoAnbyz
6Pu06G8LtqBhsYVRQop+UfZ6Xs+8SSIRZIPALExlvufdup8uBEMkWvXFlUIhUw1QzXdVQC7H3G1B
uyYkbmZLHmD0US3twTl5iOMmxQXxEJ8CrEYNIFw6LXcuig7/QYWUrfWxOmnWA0nTrnq9nZgKkUqu
lyfyg9wFt+PGggmIZ1NyklPa7Hk7LPTCbqkJza6kun7CAzBuitWYRotNbptmnTcSXYo3fmrB2yBg
dUgI5W6JOyc80tABqs9htsoU/rjPpNEZTYKjr49GFuOlvVdaoqaQZptvLNphALL10xsG4cEXGONn
PnozWaKdU/bwBhSsAf7+wWkJrWKXM7QL2HaN1Q30Izn+da+7AcFd9MV/LlFCo4FbuZRMjZEwz36I
iry0iJZZEMfmPw4S7KbeFCffaJdkJSiiwH6T3jZCDHgFQ44L40kx2jKgRV+PC8ZhArStJsff3PBc
2r13jPefz1gXRB/4vyFaDsJ1Iq4KigDii3vuOvEig/+/HGGNzodf6CzNzZktUqrK8LDFJGrqC8ub
x/Gkj/+lUyXh6LjoHCf0ySk7HwHo4RrFloU1rnqLuLU1YlNF3TTgFPq32yAsapm5T278cAVegUPb
dQ/HdER13V8lKESEYuobM/Nh9swdU67Ryq+BYAggSWXj8N2bUcCpWXIocOAr92n7XEUDVBpmQl9w
wsLdOjvYIseh3JL5dwjlIA0qRj99czR78Hlib678HSi1f7Oy/WfEBffjngwwbwqwRNiJ9RKLJjUA
IlA7FXIuktTAdxZAaEIaj/yhb9pnY4GayhsELzreTi98BCdzHa9DP8/C8aIcHeEFZDHeryLGp00I
gMAEWsndQN64U0WA+DctShlgS9YuWLHvDpBkvCtM6v+6iKVHPCD5g0w/uSJ6MF5N6XEnNKEN/YpY
EIGPOtYkYVTJsBmh5KfYmWzXnYGvMNnoPPlod/g+dECOQAhhB203uLd7gOJs88ehjeK3ycaHqZYu
rAzaI5vqj0uB2uV5g04YWgCHrOYJOV60Bi5H3taRFt+tOVpMyzDj2FQjrbNOwxlux7kbQWM98tJ/
OYFsDBbeR8CgQbJVP/H0RaXAtKRn2WIazcgJoPmg1LUwYYOzSWlYXqvtTHVc6d4BvroYbc29/JgN
ia/R41MphlmeDC5cGSbEcUa4I9Kxv6UH72IIrRCjq77RuA7klTWJglBCqTCGL3yfhiJAr3kbX4+9
gUKYQrbW9Mu2UlO8YZ8kDZoVbMv74ridMsvLhfV8af4xJErpNun84Vp95HQ7Ppn/MMWj217iDdNL
q/sUxrSIf5F4Gc3CtMtnodcddxFSdN1FMkoc/wBjO7r+Hf0vhQuuDriG7mAlmmfnOwbl3CXS84xt
rapp3KXgGCU/UBNtQkJKNOkaICIB2KId9N6mPSLqL7DVt7+YKG4TGkMVc233qQ7pF+IrMbao4CCd
S/d5wVPwLW+xZmLe7JxP5hF/IAJafhvTMc9o4NT69MW7KMHN4OvkVlwzHJb6KKz7iQsqTLKFjItD
2u40geqy5zxzgRpmT6mutYgvcLXyLPf9RvivOwOtTY4kk7jYDSyLojtIYNBSK/G2zolOo2QpIUf+
AkD9+lRozlFvyV0JvoABbwrX7+nfmer0EU/OjIIkkcNNrZPRSZE3/sHohgj3uPPiaAzNzbtph9PZ
sidl3YIoc3r/XtrA/QllLxP7yXQvaavp/5OjJNNrKX6JSOUP5HNJinmogCQlgVyFXQKsBAMuRZR8
yOEfaIVMPR8yaXmmU0iZTQY9H1ihy3detPUWSTtiL1q6sm11NwORKYyr+Np7FIQck3FqFLs/RZjC
kO5kgI76igibYphBMXBgOPMWeBO3CcXSZK90e1/UT6nMpktYnfMGSVUYm6ArQUe82VmZrUrWv8SQ
lnHvjtupIdqAUmiQzEKtlpucJ1+H8ZtT1nKivNQU8Eylj2zJ9VtsJvyi4KEGzSNM4MJj+llO8SNd
nSTQ1CI0WZw29gHc6OF/KkzCY1qAnaRhAoHdrd0Ovuo2AN4JkCAk6FLpxaF1rp84TgvSQ8ZqGY4F
rarP/ask5S1n+eNNruzT0Kp7zJWXzPAJk+v1G6mZRm33UIvo21xvJi3+BE33mxNF6BrITv7R1vXg
VwL7zEmctt9QwbiL+mWzK9sFTLtWYmprDtam1cTd6Z/gzXe6MR+ywYGAGDt3d+ARGB4lBPOMU5c1
e98zo8YZKODR91G8uufqstwL9Q3zHxKE9z8YQ8eB46qxMYsDSBucJocOG3xfcYUVwnnJFSP/GeoV
qni8J2s0nbFY5kz0+S+tTX27MjakK7O6ubdP2Hwp14Dzm3FZyjkqrRUaaYb43npfKecbl417736v
GVhTN5iZpwycO/9KKPH2mMWrtt1iH7Uw5LpRmLHJF3klmL2Y1A82xT0ZcVDcOszzmHxH9GoMMvm4
SBMPMi2M7EU/sSfoYHCpSsRVUfHXDoM/zgMBUJOtvvHGymQ0JkdPkn7E1Hva1tAMgGvse1QgSEyZ
4JZc4yo2ikyZvWkAxBvKgwRLOsl2RuNYWffq9frIatJgCZgx1O+Il8MpPjCc8zGIndsI3HcmzFhd
sRj8NML67x96JvlpEOUGDc7PK/ryRvLj1p4GowJiBOaiU9FVGGWyvY7GzFxgR9d2TV5rH9rrcrAK
DHjasQgyKk2qDUK9iiMUvZq1fU1Va9Z/vTfxYy5pv59a2nxZqYoPg/8gbxCZ2THeHw2C0evTE8Qu
Oy/hJg+p0FGTVc0t92HvQPX2tRbUyzkf5+30rAsheJEWEcIVeUOKAD2cfBft28zeGXbUsTJIePMe
ClbCw7w7HRZVs9ISXPijVNW2Fjgqpl63HcfpqZnU2X5HzRS5a343z9+GX3LQWJrvbSRFLsJt1sL7
s/D899jjKSIkCYn2fwdOI2ekZNzYJ1PxNhn7mlFEL+RPul+amFshnNb6qQJV0AOkBYm1nwLMhNzB
Gq5pH0+LzOYWSoV6wNdBvWAfq9GO2EASCUyDA1r1KFyhsy4qDQvXjfXCUHG+/m3+3v/KisPqJP/Y
jGgPpPr16ou0zUP7R2G+pCti5vN4W3rPpJQTSTavjoOcdVL+V4DhQn83DC1dP7bSn3JyjnkA0h2R
pj009PIf4lFKrZsorjATd4yli+sWsxa8GPvm5m43mbcKjXydYnHWKm3gB+F1OqFt17WAVe57vixT
4ElJDBM+wm0yXqxbSpRyMXR7paRJbHvUVVkEDGiVC2OSKuW1cCNt+4G1xBM2L6f6YypS9MjzJVN7
Nwda+PYWDZjGsdvEGpd1KgX/Qt8mhDtXnvwbSUguhCkaRn1qkpRF75mOKklnu4wAjjO+77a3I8G0
fQ7002nfMB/0yExz3j71RgmRb+EZ7CEzmMEQqIGCFtHjYMRrHnQ4rB2V+fysNAqcL8BYFSNAh0pH
+ZLwXneKufBdnExwGWC3aTgwcRFCS9uE5yXWwOKN7CFMKNdSvkq2nMAZX3vXjCIREwEg5d31HXYp
bTekhM4tVMa4FS9/z/B+0uCj8UJ7xVjNbuqTzsuCNaISFSj9G+fzZzXnipd6EvYSgeCjLY5311gn
4XOQBMQvct1DRz3ZFvkfemZnw+S3UTOD9TH3OM/BfthtCoytl09CMyf15GJc7zLetKJPEP5pqMki
64xMz1CwePGx8wdfsuWr9jgqw2M9nhcFKtnDuN3ndYoPOkEA9g8r85Mdsn+ZT1MgeQyK5f5Mc/7H
K5Lya6Vvuvt3E4B6w0mxIBZMEnUrFUEX3ooOjkyDrI7IwX//OptbesPJHYHDtapMG6WEAvaJwp0X
WygM10TmM5z10KitxZpqHt3auRSO4N0L7nSX5W+mxA21LUjB9lUC0Nw02VWvbX++6c56EBoHVukM
w7XjEwwid0LXbeVDjAvLO7YwnmUhBJZqDbCffaJZ7hPQlsOlLHk7+l0dvqPe0DwIUZ+LW5yLx6TA
Cj4zNiuDiMmYYojuA2zNWAAXNig4rWWZvcyEGBUf3xg9qta9CqoShepeH2zvvHUvEKbKz1dQ0RG2
HLZXsKXvRdqvG7p55w45STiTohAsorWOogtgkQUm0okCH3pmkQD1kOylS5YYuW3/agh6MGRB3/n4
RPd2Tm75S2M6GatfYTpviedj8SYT6pOGfre4/LTnHdw1FSoJShgqh5xz+Q/dzX9vSBtYqntTTCpJ
aRpuMjn9o/MdAc2Nh8NQ1BLmM9jzjWwlbUdiptFq/TaYG2d4uIgeXIvorM72FYgp7gHsJfUzy6UF
IKjjsBZ5OYVirVUIKBrNh5gBjaKK4aiV+xX5YrWH7qeyd5lakyDJSQN6kgPrTQbYq5NRaKBNFsWH
8u0jOozX/AbSAE/Xqc43J6IpzYAVbUvUB1LuiBKcmI6eB0CtgzvWove7jPaUomQiBsz3yFxMt9YT
a2auyP/ahdsZet6hasDb5XoJEN+ueF1fClhzyGiDlYd+2YHeLNHj/95BPTO9IEPDp+m66LuPzS4g
1G2GePzpCNP0VgudY9/lPANk19k0XAN8w90XICagvDuXUBNI9nGsPO7jVMlnCaxrs/l8ERZwarjb
T7JF+iAe5hhyaK4WaBXIfIm6ZafcEI0c3LqIouAqU5n1rPjuheGIk+l1rD6qFiVVtUBxIovyPsv9
1zcaBW5BAAUXrp/ArKDVzMO2A6oh6RulPu9P4NXTjxCIfBWj0jgv9KjMHScXJdLab7ek4Nw4sBLz
tjlLsJUJOMg/3hDJnb0ZdEZPNoBDw7Pa7lwnf9BzejI4wLJUqLPJ8aMDpIHlakfIfYI8Tzq6OD/i
uL2SD5M0Y9+6vAMwgth2AafnN5T3md2S8BeS29YOZ6IrJcOMMVDgQ77NS3OGzoAviexvm7ujsuRh
BKuuSN2LMRG5G0AQPU7VvIGnF3LKjQKJFWSPtp5uhoCnWZi6GdINq4GzdZIXpCCKz4Whdm6vqgvZ
Pp8HNOq7O5EomOh43thqGvVy8WkXp3u4Yry76Q5xnudX939pmepar1KtijWvcJRqv3tZMW63MFv/
ELjwZr/ph8rttX2v09Zf/vVLkkrZCNuQvjeYycbE3eVGKXdtmsiacysUMlFGOBCkSYkuTPRWnkT6
VVJ197OgntqxrM0TWpj016SajbtvFx6H8g5B3PemM6MbrCvpNVNw5SqPyh0EhYI0p7r+hsUpkAtP
GBwjXqOC5rSAYv3pciSkD0q1+WkhbA64SknSwG5VHQ2tzhJ/q8dk8QGxN10gPVXshq4HyT8bywyv
HNywwDwxyAjZf5ruXPGQx9BX1zNoRemx3OGnPrFMj+NJTt4++ibLp8uHz4XHQiszbslCGs7htSDX
J3BbvoiQQXhy2QcoenF16UpaIniI5a2b4e95Z5KF1nsBs1mCuNF75Tkxp9tITUNShzQ0JYOK7G7I
zsQ0WIBBmMEfoirzwAKEXvaGSkcdUVmv1eGgSDMQ81g/I321yYfbSxDaYEmnmaPY3fAYGl2fxXqD
qiZsMFO31wePAxCieFFAItYlMWwocdhZXS9vn2UQSk+KGR/cqBEu+GZDydOvIvhVslUg1DWVlaOg
bSMbnens8oMZt5iGc/NhYqEQ1ABBbfxTZSfHE/JjSr48CLg19YP9i4zkm6By8QV5PXQFA1zVdhzW
2BNKdCTgD8P1nXLLwkI0KTPPEFYEqeTULodvwnjMfLOiBgVl9TiZC5amKld/qovhlsdLPENF0kYG
B6xTuoiRlb1TsKLkwxGNzm85fOhKfiS8dECOVZlVcW9xPl0/kFs3RHPmSCnsP6oxSGf/s3SnOelZ
c0e+LwJZs4Il/UUnmw3rE6mb4BMgKNobDGH4j4cZjzY9cHPYKALvTgwYITSFYZMpTEUzNoZCsB2T
jedsMZLaP4UrnmWh3RcpXlLdNBxefbZbLVktV5r5WJafg5TKuhMrJ2d/JdpsJU+1WxzyLWQNXs0X
oqO85PpZssHe4FuemhKFHIs61kol9DVUBfgbrx/GzCTWbOUVHfsuWiPUfPiF3e8u76oi4Xv4naBA
V9xrW8pqNwT/kfQOJGJXlcxidO9WI2zTjaqYQUDhD5bi9MguN/q5dMBGtY8colPphCfEN4KyBUCR
4VmM+JdJglFewzylxxAl87sL231IQ4lubviNlKyLBhyOhYSfEyTCMA7hP5X8UKihfAg/ybKaVo3e
kMEXdZn0iWPc0Y61EJXZd7K8c/Or/CRGZu9l4E6TZOBMuvpjSG5Olid+Ee9KxReGp8c8vTtU92mG
VuyrNuZuJmLkFIz4GqWYeqogbfL78a7rK3zyMrwqs2CQ5B/NqhKN/66TQAaCdmODx8wQyAtnJAUP
026ehLDpQTl8DzHaT78Fg6gsbHeMJesZtwoF8aRQB1fNZz1kXovBvvt/4njz9Sp2Lw3se+HiSLAT
q4CJk/0DVS9B8fbm9POwKk7I5qI9GVZlt6tKOT/y5hUWkYSmR6p/mo9BD9o1FfIrbeR9U1DVBChk
W86pfC4e7dqBQjOqcdpwTeKszSqcrfR5Yh5j5MlVed2A+TkzT8b3UOZTWEMwoj19WTv7RIX3kDQe
GVHk4SUZ2j015trVFaOsikvEYPo7YjVsZEi1qnndLtDIF4Q+8mudJFO7SvKkOO8IrkymTOvC3Md/
PQIjWHV2qQpNgqdeirL9SS5Kscg20NYMIsuXgE+JozCAFP2gy8UqYACp7cR1pQHUjrRJcLU/vOoq
PlD2cyTM264+aFDq4lgPW22ADeYl/Th4giHN+oLFZNrsBKi0jRcF8OVAwF+tzPQL/tiW4QuDqI1+
D/bOHtbdSa/4q5RO6EZ4HT5YRecMjgUxyPcLumsphDF5ONbklmuWb54xKPnHkaTgrD7fcgGkdBNI
xb+dQEwQQZcrGYMTONwdfZ3Ni+JT6UrhSIo3Fu/h0sSdTU1EK0s4SltiAjVgEeMZjyx1dLnLsxIu
r7R/ZDlLGRWhWUHpQxQnWnBkcPtSt+AZo4suRjCvzzP248F0ZWneuMmqiUVLHRo2SPbkEY92l47x
FTUuDcyQLSR3To5jKs0B1M8SsHxyQf8Bb4WvVOdk5oq4AEcQpO7lTVt3Gdgp++amXtvd0YyVQ5tz
X3GcsPP7OaSl6OunFxd1XIfd36nRN/7TWWQuGlvW3/pp+Dv6PpxbZvsI29S5r2GsjcX3Uir6QnUJ
UYUI4t0hcIGK2l/WbKMYUgQ/8hA/+8Hy5AXKbabKuHBV/4pjqpo+VSXFRCuxGNhLBX/LUc3f/u36
RYjz3pHBqI4Hv36azGBNWL1lO8AWio+DqBFWzhadHqe1SZEOh6TKz6Vsa3QOL6L7Dxn5utjQmA1W
Qad31obM/m1oqDuuyC7ppWME5cYiR2W/GFqgcR5TR9B2Lz4UmNgOBsPZijaANC6DQNEvHvmo3pgR
h4aRdXV6GbmHPV944tV5rB8C7Ds5PBe7+kQrKT+MW7U/pTZNYJYjlUMJKPgOQdUg1+Icezgpk1Kw
3lqN6Pt8tP71o305jyd6LQi4iewy4qcu0I2TmRHolfjWHGB+JrilT2Z7k3/OyhVh4dfo5ppbM0q9
J/fa40DWoyCV3TtNfsEC8CtSMG5t4fcLCxKr5VXYMK1OiUAHXNe9SSb6YtX76F+suzxjlPuI7X1c
ljkre8UXGeMqVvLldwjbBYgyA7PQeySEAoBarglpEE/6UDifm94/bFed5b1xHnyLbimJBN+GXRip
vaA6idItwSi3JSdG4SmaLhEdhpabUM/8cRc1xs5L5oD523wvVXssvG2nlf85ARgDtsgVg4dt334w
r8//9J3Nqx63x3bBr/iU3AP4Jl4bfCD1iDdXoS9JLAybhwa+dO7s2/v0/+YYvczC1EHbZxnVeHEX
nWk7+t74q0YTmLJPqMLmM5inbfhOKEtnUBUMowtPxb5E2Ic75OR8E2yRc+mv3wXWTouHnyR1/XZR
3iGrM9snKG6IlvNt8YJVOvj3CzZ2rpfsqPMAfITQuhiv81jKqLsbbxR+atXNBLzgdAU8UkY7dwa7
kpsadCcAfIE/sgK+0SoGW3SOTZHLLvjoHguXAVL8+DlxhroaOzimEgboeWv/6mGZXhoQtxKHlUlt
F3zICcYI40C+bcyBTDyW7lrIhseqjBWgWDNzY0hqdWiuASpQp8+jAa1xnKquM0Hrf7oRweZP0Fnm
Jsfxt+IKolJToccHAIXrRJuqKXrqFzSgPGbHRb2r01afZ9cjMUux3W/Kw+qL+hZNlkCnXkktgXLR
w2J4zGDgwr2thPCaTZqj8osKXENR8QI15Mz2D1UV5goPMU2z6IyTGQg3IJqWE6aqWi5lIVyPWpUl
ekydTwT8MYfCVRcpRviLquVsSb3eYuY3mHkFXiZJd/W/+5IJfP4pVewTq/wcGYE0j5A7tTQ8Dk8g
2E77a6hTql/x8Phyf5F4lc+g1F1UIxmhOoFaIljFqK2paNg//cjqFUp4cmoDklHp6orf3ppwrVfd
vE6H61wRniyconQQ/u/1qm9v+pe1tgCH+SbsXu6xJgDyA9sM4IGgIHZhjR1EeRC1XkFNya4XM0Fg
AOXXxnWuKg/67NaOpnv2AvO2aK/YaEICAwWBJYgUMnANTFi3vN620j+0TbAD7rr5c/52hwKUA3Bg
dPtyouLJZRRA3cdHGfGShEs4ToXoJmpzKsR0RAJbPpDoW8gOeyAxzce4GVO7pcTpvWcVvIJ8CAZc
/3VWLU8qTYQM1E1C5VYBIaYrfAk0AM1B5cnACmkyZvYS00fKrIL95g5AFGBcw9ySIeS9n52rR/Qk
REh8nhtEMluLIljdoS3h40zjDIszpGLNa63tpuBrzce6FZugJi6eBQrehUaAb3obGcUxYuuJvy/b
i/L7pc0GEGwk9MtAEA1MZZ8i5cTp/pQney/gPCPyVPNxvIhll3BVpT1DL9AwGqBpJKfF2j5tfrU9
EpuZPIvme2aYtMFJRArpA/KALSSl6o8F2RmMAyqFcsmpO8X7R6C8YtOV98bk7j0u1eLqo1Aw9hYK
J2DWFSq/y5d0Q5EwojETkMIx7ZLgM7oQNg8pAiYXtaLv8UPbzTf1fLdos1h7UAYiUu22KA3fX8Za
/AijcJBE14sHEOxjEbfDHMUQjdKRb5GUIUQhikVK3cRLLhMc+LXTsHWZOvR7yBx6CBby3MerTNwg
dpvTH5CoLQjhO32zqpX3HDxsqN6oD3p+SXmlF6fnCQOrORLVn7NVgeoaAn7r/t/3l1M5A3NY+aqH
Acnpt1GcFYlmshFKChyHUClod/O9VaOVt7C+Y7OVPyiccp7DxrvSOapI0pwL5p4lJMz3uoztYC7L
xJ0jesvZu6AxiIBH0ZWZps8hPE4bgTmRBGfZcmoMnTmGcReHMjuc8/daGp/3JxHnLETvBbuZbWlJ
QHr35dgCkPdpAy29OoH22+4GFErHt2yUM/odPy5lHBZ1areHPxIx69AmQfRuO+llI2CeKWt0+FKS
aTAEMariV/dy02hSW58X2sGTx8Wbef6+LyrqHE4QgtwFVDNCH/6ZT6pW1BIS4Zht1cJa9aCw0UBZ
1OqB85aTwboOur6RKARQUNgr8RyOjyhfrJKWhvIaHiqFzRnU8XgYb0eQ1i+Ef4tJGvXMT5aUIqL3
5HCkGuq5LopHXG2udc73SIhowEN7S1QNAoUcMXVgG+yAQxgQpf/JqsYzH2yOcbwDIAvYWq6EUSI8
hR8oSukzZLEG38yg0NMInx+EhKMU42mQ7w9Fu7PEsjuCPpgLSxh/eMRpX76BWEJRNAQLprGXZDFM
aHcNXSfxIjwzmbDqRuTt93mNHkicEeROwodX1APD44kigaaNCa/TwnxJ7o2nHZ8XfMun3c3KuaSW
tncRX5xbR2KDXwhvfYgPjTCfJiZi7vBnhepbLGrmz/vowOctPA3yI7bFJ5pPDsZG+lBIwJg1agRm
TYZ9QMy31jCnPgUzQvPO3PHXWuaqlqE64O1+kfl/hPg7fZDKcFCH34VuqUglwGPR2Jvhv8tbe0Hl
/8FJPzIVAqXRPmFov9VyrorcZav7LBiAxdVufc1IfaxEBAprj/F9PhMsV9xvWeAO905TvzD0TfMU
kFtB264j8ZQoBA48MvhdWTPrYDVtTzVoDQ7RRw6g22kh1l8xaGosmrPXCuWbZJP7Sva9uOLmosfk
Hu3ZFoopQtxfoic1qVQzKk/UTOzULK/i3Nlb822W+O8m0sLiaY+qIYTqFX0Ib80xc0Z1pZjmwxiW
yf2u9P6M2eZNptJeWKyPEpAFMnTtwqx7nhXqlXQ0AMQD/wpM+mlJUgihBC9tmhh4v3t+Anz3fPJU
dI5Bae0szVlNpzi7MNuLKS3D/zNgNyIbDG7ldx2CXxPnN6uEHWgOO3zFFKezFeZZ4Lf5zIwFwjxT
lPRYuIbZYrYu7CTXzR/9gZk/gm+9XFD5yeUHu/U/iTYgU3pHklGAnU5NWXIL8yjbUerokuQc0ue0
BkrVrureGCtWaReLaHanZ4lrqRQznN2FLvQr/oKouuHcnOqbXVP1mwEMAGK2KB/dG/lh7HsHd/uP
NGf5H69LjoOXtOmkFNtOqebZpWL2z/fXTlJ/4i9+ppdupRXwRhC0+usHTerP4i8UDdHy5p7QXzup
ZeCvVlI5IOs2r9ICuUiRLL0rs+Y8vCGAELSmTULnpT635Pb8sATjc/xnPk+ht3WtwhdBVsV2Q2lS
R1vFCYjglMS8Fox5XcuOAjB6PZ4fbDu85BMUXcibCe6fIr29Z9H/vXQZVsrtcJ5brwiUykdRgwcK
uOmdwEsBMfsq7BvHeBLj5deiccT2LZ46ai8FYko4vCb94lu64zwjFKiOaTC4+8e6bi92S1ig6Xmd
NSrcWTkQPtUWvu/gMBo2UR8hWSZ9gtRP2dILwxQN3gioQVnuxkojIMXXHZPTN7ijOpPSWbdLDaXd
R3kbK/mFf2WyjqY5WeJ5zPfcgDtI30v8VtlSsuwdSCgUyI1Qy1R2jlsUdrPTC9o2OrOlZxGm9e1n
Z3k3+5J1kcEh0+npTSI/6ctdeI3AJ0Ad9yutmkC0wUUXCXlP/DVA/04O9R4Jr+ALhswYqhfQ4uLy
WVdXUzQRcvB1lR4Vhl+ddWDV8X+JvqN75mcPc9pSaFOUTCAhLqAQ/YoPmtA5D0ykDYgLsMltoUtE
hEiDRwJL0D+Scx7KSQEFK8+H67GsKxZcqhSYKYBBEPh1fV3oI3FNS9avS6CWQQbeb210Ivv3BK2C
kccXEcuDaFq4ESX+1s9FENTvkcWCOxT2BxyZQUBwW/pKgj3jjXrKU/NfVOyKCeG7bPZ5VsS/5idb
WVTu5ra84DiSzj97lYxsKxivW9tD84iW3pYioT+Jqj+Ju1DogI7YBOnIPaeIt8wBoihSQ1B4SENj
T+wzBTgNIlyRnGXGXWc9R1oRGCQHgUk0wR2c2a+A4EFbc0S0L3YToSN6bAdZgXtyQP8psaSWaEHb
qfUxTj4aHVHHjrAFsfuQDubuvRCdce2uQJfpG28voaEL9Sbnpbk4S+CKH22DsmiQoV+gSwDooZow
cumBclBWF/bDm380cQMnbnDVfwgTS/7EhdHND2Kue/g3a9PQPaJS+byMzdxob+OhQOuy20680eu4
4C10dtJRuyBkM4jXX7fLxZ6zfwcCgfUADLIHsKtC5CjYjXi6E8CaDAnyHROmRz3CxQ/9Il8Vo/Xn
lDXZjoURBqXSefXdlt0UQ2se3KEqRQ3WOtyOctF+d6WXBNX+mlVDymrpbcmHUze7CvGsj608vLuD
lh3SVHWDvwqugMEBO4DRJfc1tniqaklV711vGjz1zc50nFw2C0jDCE+BvASoNowcoPuXWs9LNvzW
jvPLBl35PFnd0NB2vm4rKwPOI1ciDf/aIW7NzaL7dcqG9vfhpa3LD5lhl6nn6SFAWf4n3n2BZtXB
bVWx0Sh7rxX6aF4y827Y4W388W2qHPpCggyivQ5jsQ7DivJkYh7JrcONln/5sAqeuRGORFIXTEMs
AxOZo3Ridp1n3ELejbpkKt0LDG6rFMFygmoZAeV9rMHs5iaa2fVEroiFFVVIUCqUDkfniiIRFllz
hHrBgdX8lMrqtrEpU1cPwUS0GDoUTc0mlpKBiwEa5h6mOyz2l9kwcwhp/SO1fnF/VZuvZqREacDJ
IwOdn+mlwbMqbeEosspqH4WVj7X7uvuLbHd3fM7M9GZVhvoa/PqasgCiqwndKHsp/C6NpAhF4SbW
Jd1UM7sIBkY/cDsGT9BQlSnlhLcdCCDbKxjd0/W/3MiOwQ6Epwv0h0m8whIK9lJv3l33GtOKH2Sk
T3R2plizQmjaNCFHKDCoywQ1c7LUgIbX1g9REaAuWol+rO7uP38/FEpqtkGPwGgHzrU4UGx8bC7T
D4gSY4AhuwiS9ym1ICy51c27VZ8t/C5BRcOWcoadBriQbpdXEH07QtGft0tfSwwKCT5Qw+lh9ria
aMRBjGoyiKwlUWcftSTt4uvbiZCt/tM8hldEn38U+DybQZeeN9vaJ1JEoynp1KorGCOpbMVX4Ck/
Szhk7aKYOSeEny4p6u4zQ/bkgg1ZMBQ5bySi5IpRC07EPKoua5JBsoISFgDquuteXXBrwpNVg6lf
uGKcx5fdCBoZvfEX9r7wKl49djq58w1UVpFXyc741O9FJ5xY9nFD4YF0UFqpcpqpejSsTGnm10sd
KeiMtt/ROYd6fu1h0UYWv0/s7sXYaf0zDc8QbF3WIadyHS8NdQrLcsu6pmQEC3YhLpw+tLl2veyX
BunNJ4Xs+gIYb6f99LdrL5CX7ofEgnIdkqfXO5g9DS+/CE7ceaf3P8f0VCKVX3JAHrrDAV9N+3Yg
BuP3VGMHApUzCqE9ovPY/PyF5bCkOkb92DMzQ+hUaBKkp0RbuSH1Mw+tnfjQLXwuHwLIso/9br2f
08TWQdqDWWyLodeGGdN2rjnHqPNj5iZpRi+16r/WYe6xLt1CX+qWS7aMHLAJiiFfzxBqEp/rrnAw
jXSxtlj5PAU9TcbyyAwaSbdGInxqhGnUnV7bEYVOYYxPwOXBDWmE0CTnYh46ANrDRmyG28H+u7by
dgGqIewWzLrqP5WyseDjTH2sL0KdEL8fRs+x+QCGJbutR/MHnQHaJ9Q54hWBZtYkWlx33QMHdimP
GdlMVR7TU0OSQN2rPAPJzII7iNFlCLolriNe5tuuansvB9amv2t/kaWEwqkJDjOJmSKIIs60aR6R
Xzxe+GMQ2c+kyDeB2DPPjGfYBjt5GcT6QsdMZJjuL9ZcDZD4Gvx9QkJvzgGqf93DnQbz26av6ThS
8eiZd+c3L7toWWZuJdVK+t0MN7cWCxfwPbcqURxPLrmRjrlh7QcHkZHm6aGZQECntJIdaj5arP7t
ZWV8UsaM+OQZOHhgTM6DXjbyYyUe8RL961db7slx22yOVoNIgH2U/fGqdOMDAUQqJvYB9yycwNAz
DNnZwhybkc3mWAxVXLx7KCZr1ERhDu3XuIy7IQfP6zEZabZ5/9IPR16hKMOvkexyxirfOR+ZnjJW
rOAGpyI/MXxb3t/bPWk7W+QNYVdWdzpFVBQx42LNPNQ0Uqd7+ti+FnTISbZ8KRNd+c5wcJXWC90H
eulrAWezt714mYOYsf32LT4tuH3SoolHWGpwFkvR45F6Q9S7UHr8uV7tv0CEOrEIALT7JkSsAOZ7
rD05wnFn/QCLGTrqAwcHPfApDDhK3rQN6PVEOPapa/yrCUCJ2aWw0dGFMLNA4bL2t07B4pJD/5/h
tzmaZGgYnT5qv5QSramP1KfpdFnSoXP8n/dCc4DVBVdLp/9OY/5TIlr//qaDV3+G6Ww+fh0tPoUE
5ba56JURhS0yjH/y7O6UBJz2uKY2KK+o/UMf3fHihiPzs+UO4ipGIdwKM01AlrfyD2hG0ey2wGrM
SUCU3aMaAuFjkS6ySiyiRRIy0094z9t2nc/gXUhrAZuVOmpT6HOapbhysk40NRJsQT1vuOcchoT/
bjecZk4ZBma8ftOgqOyzDODQF+KqfYidTvenU9ktR/jcU/gA8TwvRVedHROpFv3azJP/HE1a3tCk
beq/3MzUnPAtaTzr0iGf2hm9SkuHJ9Nc18c32elNzKct9YTJQNzwGAtP+k5bxT5hOmYPHcp72qr0
2yGosg8olK61gEF21HgfXLCO5arK4Kqif8zt4s0iHCcxsCUHglVV6fzY12973tT//+MbX+2TP9Kl
P+S1m6zBcCskhrXcEL6vmd3u3IojSehBJHsygRvkER1nWnvbBxUWxIJhVZw9uMjrZ8V6yMZKTDOS
f4lbpuJoWvyo21L+GXzxKNJUf6/JG8wQDGWqUCyK6WsZr70QuuOCRdkByAuQ7H80tM5LwdjCqZ5p
QbzJkHRboAS5INep/3/h45rxNSBP30Wd+bWNs89TtZF31t+XsicBFvYSj3jeDuagHq1w+5K10KH7
MpZ1ncVqMnnmWohDGdjayixeE4irbJT1OcnFeHGeyWbVmGVGAaCDGqX9k0TOUHmAteFXXmHAghx4
wCTiyWP81rGt37RktmaVhsM/V35fbNa2iD8jsX9xMRqunCQEX5s8o0YqJhbf3zhxSvQ1UrDOqdqB
YYv0zbocmVCCBkEs2rtVWD8TVqVwAv73209+Qfrp/ZD3gc/sZtS4wojdPHPgM9WPN1XRSzmUVTEV
+L5DXHx7bwbpn830u1IJ7HuSvP7+VO24M4pYBiEP8PNhL+hl/fng27PoPV7P4/DaNNPCvB2ug2T2
Z6apvn7RDOiZdqLEtjMGfHJLlaJm9sa/sWigY8yFwf+zdRE9fqHfwkfhmccfcoWVTqaMJp+uOwn+
A2IuL/AR3R+ljh6vKOH3kXipOgBYyfTjMNKJTS5R5bh2b4XMFahqmqlAGhKFdifWzi3W7f8b0uBZ
BHmApdK8O81FVlYKPfXWk5WFW8HpJIznppXDKuHeqBezUb9x9PS5z5vJhXVj9JNJ4TcduD5nLoup
s6Z0UPUPxn0t0QpDzYm231UW6NGnmfDphb6UTCfrufNq4aaRxWYbXPqMPN71zloHzgxLVylv9p3s
SiMUDXh9p4tPTGz1w3ct9feeiFUH9SwbFhQGMEQDMSRRKSR9ltCPBskcrTyUkRp2jw9BmW2JwSnA
OM7KUrHtjzQO787yyYEHk2YqgbiLHV18/4LQ8N23MM4jiZ6/vSde92UZGdHRTTPlSE+ft0Qcz5fZ
6DrlpFHPTLVwOWRo1xqOsfTJeMnVqWO4FIzqR6tZ/cWCRbKGVOLjC0T5s+PTR0BKacQBrg+YOPbx
o+NfsWsZKpUTrLN+BYGKH/zY5QR3fpS/lJHQyiFM0I5cdZYa5MJWnQwkEWc/R+tDXgD/J9/xvQSB
CNKalTbAV6V2uTJFnFXyHj8vKloVVfq7mj1S1Wx9536aY0CCocIxw+xq6bMk2yRDo8eWVp8NH175
sZyKGinSIxU/F8GPzMTr3v6OG/nRx18Ro9BnKenEa05iVrvoHFUjwIneWlobTs2MJBAzW1OnXm8R
Ay+Cv9M/nvYaund2ZiTvdXlXrfUXZRLgQpvmnIR/2n3sU/+xdXAPE/Og7LislAWb8gvAweKpneps
ufi6UEwhDTNAcbdrjnCtTBRonvJPwk9CJdwfdyCSk8R1vX3bLhBqWznrhTSbRQhQY+fauOoOjMGi
nsSq0JaojwDK4V2LQAP4iJAeWmokr4SJEW6+4XyV4yJDmAIQRsO0IoUAiJjwycZCn1IEROYIut5d
PkpsfiGKybmYJvHKCUPCw/lJ50HA5KX2UuJge8+K/28cNcvDnLqojFrvXAzrQ0WpOml99JBt7M+R
KcbWR0sGemXdN9fZpsUeK5ME3c77VzfgIdaLCzjaykHqg+v7mPS4JBeIfNn/gRXRmZ+jGg7lM5ru
HNg1wQlwUh9tIRJZXQHg7MSV6oMLPnCeagUw0GMcHkzyTSCE9zPpt4Fz/sUR+gDoeS1iUBHizhlD
0UBpv80Vprjyc7SfHWYuEZKBBBL7rBv6yVYFO3X0hoWL2TT2+XjaeoHjhW4bj33qM8GaviP0cunZ
lrjxyBLjPdGqxmqVZQF2xun7m6+j+vEi5hCGGFTj4cAmqcewzEPQ5IbRBEzvxfDIOEUpdfIFVeER
EEUbEGivyj43YILL/AT30d2Pa9QGA54V+59Yao+yWxSKUNuAeSgNm7A51sXLr8temRctz/a3dPDi
tBeNInyFavnZUqc+qzTm6aEMJkOK+8Ftnn2to2dJ0Jqzvhg6EnN8dBsXGIYgXPG+6TO6tqhg3WKw
VnwJKHTpg5tSuWlX19RcbCz0+CGcd1lghUvW3KYnFz6A3LIq/eF8y9VFXfUeCu+d8hmhiC+qBXMR
EVYsPnA9YkJA8q+OPvltyHFZxq2RxApkDyRx5ZLaXLU3AAiENtUo+ZOjR/LbglI5MaGJxm9f6ZfL
MWhCmTLsSV45BWVAmI7O0bSt2p7ItI1pT3r1UzLJuCsU1LM8BzEELFmXDmuhU5Mnm0JxpQcrRnoG
Wbvs8xhuUAAbKVOTn3MG3jjekBS8fZd0vfA3o8Oc4dXWA4GeqCmw7Xym+F4FajENynXP+6kkzLoB
r8moR8ssVcu92q3BthrpzuXqPycjZYIOYu1z0pXV8GpANET9Is0dEczXmJZ73gizAMLT0CwfGzhL
QzA/t2UzT2diS6/kBUj0Qbuyq0PRpZmlyT2MsULFSmR9p//7bga/DB2+9aJ4lB38TgvTQY7gJEav
PL0VLpmP+ZFcKP+J5fIrc0B4oPoB6BcjYBpaDKPzsN2kxSnH4/E4x3daw/0O1T8ioc1jkKgfVj5m
dFi776Q6ihMucjZxiGEihWLbMjYPz3ExNt1b/d25kbMq4rlndNl0ebzxjylYgZzPi1tkOnxFF9rf
vAtsVvcruac+crI+PSAeFZoFeVaarSlKgM5yL3F+FcCwSDtj/FGfSReTH+asXsvtVWziC3oXBHUc
be68jkh22v/TGYbY68izv8K1Jeh6PEewQhj9UWFBKRZVyKrIY3fwY2KHM3OfW6Gkzpv8c69aZvnp
VVwdwHk6Nh2D73rKsU3J5cfllwEamVsJSngGtP096wmy40z+LWI+6utZlbSkumBohq1KOEe/TPjL
PdGLqFq7y/HhD33lN5hSHrc9lUBjTSMrOZyc8iikfO2bHHC/dla3rNN/M9CnpyaRAYHUBoMAuaQx
DF13+YWX4Bugz0p6LeU/HBoyZv2E5pJnq2gxp7QAyIk9U3v33hwSOWxMLT1GeF7SUpNraeWAPidk
M1MY5n54aPa6JW/+ulXIuGuaTuz7jlndyaz8lxiOx3CVagw2eWJIn3nDolWT9ad4+NuZWAx+fSlQ
ATFAY0ygI+62Ti0WotnmfFYLSUlfreM2N4fCGFNZNeF5AbTeIXxwgvzSZh/urX4aKsK9c1789RtD
3zCUbejEx4q5Sh/vnlOM8B+21gHLWj15dqNpNBo9wsw16tfWCzgaEZbWVDzwk1b1V13SLVSO4/S1
oA5+tOO3oAWa8ZCCYcCtHeAuihB1Em80MindVH1vYpvhYC9qpas/TNJZoiEmM9+dsUJefDi2H//v
uLvd6AS9JU8+0Sp58aDGUD9ZDL2VBSSQUFR16ku8ut2LDIOPiXQh1HOSIRSWNO5sGrT72QdB2OmN
hgGo2uxq5MYKRLpkL+hmu9LckyzA9xHsCA9WzCyfx04pMRB6WK3XcJ6r7p2Cq2i0xHSYBTpkcNA7
qURkA0Nd/6yJU9Ii+/qVJYH8zPHPkJ5M112LIknK1kCuIfzJlnQgIVejgtH7yd0DA8iVlofKh3sE
N86RfqegOjpWRPZ7Zan53eT1AXmQZT/JyCJBIpBVImXq2hXDOX2/eeA10OfkoJUkjd4kmLKAVx4+
w7680AUdFbxJRIT14NyJOLRWrusFDBHdpn4f2pQvpM+R09ohZJdTbeYYtpa0HIFTday3XdgPPOoe
/BkPl06kT+2sgcXLkYX6TzxjZt21gzp49Jngbu77YRmNTkzn3e9QnHO7ViPIrvohZvBcnpihGWhk
tVANaSWdhKmXYMc4qEhE70+94SMCYs29iojXZwG6AvOJdOPvmLCQQnt1xC0jl1Su4mzT0/LzmcYx
3FFC2hUW5O5sXwkO/RdLlGg8xRalPfD1if+NGq+p68qkrckuoJI9B2d5CAf+kb/1L6VK4ySGvW7c
TvkrM7auvXEm/9mXTvH6YD7+rvyaqeyf3PI0gG6U1cQ3vHy/uUSOn6NR9N9nedTkhfkzOdapRhf5
aFfMGX1ARF+3QhhZKarvOm4C3xt6b/UWhHzVJy3zQOEktgYiaUm2MEN3gf4lHh6ummL5w/hltdjZ
YORs1zg/U2O8oe32wdLUtPJj5H9UF0r7uJGOvCXdVrsn300PvKF2ucPOL4OJLiQf/ToGi1/m0tpT
DYKsrtaf3jJ38xiRd1s1qQd4sYVqopGIQWazBgoHb9KSzH7zDH3xdqOz8v2eMrg5FZchqrZ1j/C1
HSi6PrN6mckF82PHILLm999H5yyFxJEyFl1vTi0jmilnPQD1KkXF7KxU5Op9zrhorkj19HwEMV0Z
XoNRuvf/GY6RKdOaDttEJnuU6VEFwlY7ayBqtx1xnwkhR/oTSA1w1wfSIqx54o0g/T4GopGvB0Lk
7qzgfxwk33NZJsKOIDTc4i2wegbuq8FLSx59g0HTeT72GKsldOQNl3XWJSzfz4boNgDHMOEoc1c9
AXx1Weq/sJ7ZYsUWKlphXXYSpuzUQs/DJXEx72FIWS4+r8tIa2tDLLukw2qVkK8JDO6GSG664W7i
nN2NlTP/ablvevclqcvsmYTP+3IP0aW3vvPXMWG6GbMSnowiPO3Kd1AQN5iGrmx6LJVocfCVR4U5
+ZLcWOMPnHLNnBJJ8t56nDSUpdY0qAtZJt3OVSr6lmf+FsDVLq9NQJS2XpyEqwF1CC4+cwyElZ9X
V62Lb7raYhP3phaUzHiGlcV1oytUTwJnp9ZQ8dGe/OfiZAfgi0Zrj45hOpOfVgVg4OIS9SNO0Qfi
Z+DXxzpD2XGYW89TaGvxdMDhWCpYCZ9n/DJ/i2y9Yg5xCjN4Kw84SWOePBkzJZ4OC0fhDlCdZo5D
N+6/+jZqd59meCS8mU+QdFkloVtuJ2FFuEphNpQdJ6entHA9+9ovoYCQj9y485sehYinUjsi8drY
+mEWF9bdS1zOaetV0Dj//dVvKm29I3087g0rBoPdtvtYzM3k6q/QvmSTxeC7vLfWaapQ5/BFSyMv
+orCbfBdr2ikKYvFdFcEwdacreyVm1a1Cyo85GZ+V6FB7TQln4W/I6cw9c2TSCrqgSUysh1FctVE
vTGE9vr2YtbvVsiNA+5aFOJ78qZ4nHnHgIcHpUoJejjtc7qb8j+a313cdfO0d+m7T2O8oNRCshBx
mRbnNAQ3NSLeHatxMmnR8nymluAZ0UmPO06c9ArbtWa4kJqyQNsRbH4/fFpY0mQdfgy/vZoIiGe3
EECgkwj7nwnJaV0AbImxZEs0qtpB28XlwkxbkKGY0U82HVFMNEGRDMoQVfrFPIsK2rCQ01xK1ZBR
TjgvuItEEHn3EoYP+WD+OdinyugBQ5P2Dp6OZ0Pf1FWO24twgQU5mTd5xf4qqTUXl8e6mDCe2K50
6cl/EZMWLMODwpG3vdcJUvGiPVIoVxDBPATpnQqk+NX+pc1/zBVIeu129je92t4qKm81XYLtapej
HeZrvz1CD00TuANP2arngwfejgjzbOpJBE3R6iVwrlGUD8t/VHYLbyskStoiqXg7i1RvW4PnZZ+M
rCu3CHJp97RucjOzW3X0QdVqCKRXNiLxR6EItxW/j+Wt3JbTaqYEkRfoIhAyxtSSBp9iwuDth3B5
W2VwAyJmch0cTENuIkOfw4pUJBjOpK0SIF6Yo2CkuBKoGuUJEociEdV8ZnnsYuIasRYxA77enAVB
34fVnAoLzKpMF0/zH4gzWisNcfRUNrhZKcU3TWK+0VtO95c7yfKsBTEb19q+MXFNnVB+L2MdrFRx
FzUksyu4d6xXXpfeEE7IrlsouknM4NU5EloVFMISn+s+VT36V8RnwWRsSgGGsQSz0wJWg0q/Dbnl
iq8480Hl/8ZnYJAizSKOKaofwKKc0Z7CMp+Sd1ToUmfIFGm+0VHJftXFfEMtFl40hwdvaFddVd6d
9OH7+j9CSDiCOFvr7dA51LbLSL4tkvLGgVa6Ojm68w9jyPw73N8Vc9m1LLTFEnTid4cFvjArEtSg
PEOGayx2mvty/SF4/VoVXhxubJPXJkw5CJ7OZKp42g4eJrM5k6CfcifNCn7G1XMIuBk4iBSJDc/g
FK8b5Bym2l5Z/LKIcdeYwAyI+n7+MVW8SXFjNk6UipRZEoZlym8nhqNWcv1wX1FIoYcN/pqMHoT6
55VlGCoKYMfg1WJomgKA3QvrZBbIAgWCopRMSvpeUW3KXY6e8Wzkg7XEQTT04yarueGHEgjfpvI2
XOx1h6mOPteJ6kXNGKDu3+/PWXBm72omxLSsYZrAMlO83IIh55OeuBIacH4x5ovpiXEfAjt5nbsO
AOQk6NBuoUEuzqFsuVztHifjbKXTzis73bLujonlbq3o/2QZN1AzpT+tOF9BRG8j09yjSVutP90V
TUeGoyixk1iCe9UnJx8cUW+HpTXpXhEwNiacY5LG/3ln3PTOZ6bRFSGoeTtYxSHFdAckVkJVqOdP
nExAuXzRMEOleRoXv82mQeydkDEwGaF1mloOPVnf+k5ZDL8JrTbD7UF964o97UgBYkJajTjn32Af
jPy74asfy9L4aIs3j2O6cLXnDBQFdUFhSV2i6vjCsYMJU+QWvl+sK7ah7YuKu+gjr7BwgseCD6wV
jPGsifykjAVG4myPjt7gropR52sbbS6uJ7Nt/zGIqz/G345jBeTKEe3uxVwM1VKkmfuyVane4S1n
0LlDP+Dgo77/INp4HQfvQKnXsLquQPp6tX/4KR6l80RtV2QZowdb1K/wWv8wyBt5eMIClC244I8/
+26FVfwiXi8JYrXO7e9dwPSw7+G1CXq6H04MEA3t10S46yS4EFGDtTBKAcHsfaFbR9S3R01hcuJW
+Gc/nUSMzmLT6jXExiN++tfkBpBt0S78xtZZ2JErDZCQzJeJxr4xKgCfx6knlgpPSeZeXbsHNj2i
02o+fS6zXdmmOpcCnIrPe1gwlzU+tJ81Er8HY+fyZAS9Lab3BYCkCrMtpnxDR7mGamrt8HKof09Y
35Td+bYphDeAg3m4BxnLxioKqjYQthCqozjGpUr+L4qQ8zCkySjAP5OwagGCTrpCTHt1qkqUIO0u
Hu10ekoFmBHbG3lghTbr1rHcYzBGyQ2ltICyZA1lUYWEnRaQyIr7cFC3JGwO2b5j91grsY8kJuSU
I6hZkfrWY20V0u687qXFSX/t29AGr0bUeY02Vm8lueiMoAWr50w5Ug3ma713rrohxNHvOPclNqko
ux1sKdK/qmDViIaA7OLUwcujj54qx1b5jqAzZgl3ml+2q0/IAg082Ei+GcMzOdLi+lwb8IoHgTJL
0aTzLv7xcTnHZX1g7n3HvvMObjK9ZEepIB+GqBEUNBROGIYdxYKsAYCxIsP+JYOJG2s0t9yDm7FY
Wpx+9083ZfuetUro5L7ont9H/9fmReyysh8Y+d0iAoSltSSlS7s3Dba2YJa/cG+3XzcsHrH0w2PW
0lniR1hIzoZO44qdRAV4XPbtpQ/55nHUzVYNjL3XOo5oQbz7KswobAY+EF1DdEve189lag9JVYEX
WyI7b1y5nOCky+jnNo725tQWU23P8tOKk1JzaHGgpBc6mwH2YaajdTBYWg51DD1BmZ89jOSyrO3I
2+ZqqOUKQxeBoYJUGTnJa7m5+1ola2mcy7Yd7u22asLPryytrutkg+cv2TZU7ch+vwtQI6GTTm72
Xft42DLRnSrHw1umk/l9Q+1lj9Pr71XT/HLXCuKf3Jzj/SqehcKDcqW0nhsSeTBTIrFMcypi3EoZ
dDbszHYt2NpCdTIgEEyZHGGBJDdgXLYxpoArXMzCSD4t9UtgJZiP9YhkdiGO9qSuJ3rpzT8wimjN
isHjGxdQ5I/8K8Bkjs8IBolhR68Phy2ZQsaXOmGp2zzwbtA54fAusSOHVURKJp49bMpW2e7ymYdp
l6ntdoBxUvnC5bITPN7TTAL5YXQoqTb+VuXAiiDw6BYbSwfWpWJaQlsWvs9LT3NCsWbDWiwYVp9g
ArFdoIhyXSaOC2dsK+Y+CTLm4J80nNAmwbhvvCg5QnuOb+aqhXOwWlbCB7yAXqUZXH7hl3sO5kx/
BETLf5UfWDMgnI9SqDVkoGd2F1ljqVLs2ECtxiFSVh12Lvl37KKNkydttMMBUe0GdPEa9iO69Beb
hIZGr7RChHq00hGJ5GGKdK+AjN3u3/7RU00NsIoD4hF9eHzi6R+3h72Ah+LX/ZhhiqbDu1/6oZRh
fjdjX+oFCGOUTJQDJ5dUa1Jgm3GJvppNM0R1xzwpDo1pK56amDmnZMY95FjELKlPXSCkKilmN3HI
LNStU+ciCppFehIAngJeHr3rZ93mZgbLiEPbsHjsZ4L8C1+YJ2VIP8A5RuvQ0BkztvsBGhGjJzFA
3SSZmg7/E23IJqtmvyJTcV0VCKAYMRhiMitAUlPiLlcH/A0WxrmhPRLw7KuOSskYuvwXk29BRh/r
mFGSzx5reMmh8mIQrt28I+ro2R7EPIJ3NC5zHdioqlTj95xpOfKqKdSaCSMZmnBrEqVQJNGhvjcr
XtZf8kTzosXX32a2yB7JGeOqj6G7O6RBZvwRvs4CHC4HOD5kLDOARofT5a7MjEab142I0iV83WSf
Xq/LYyE7+gZ+hVgcgPXz2+rfGz8bEbzgfAX1XVjyiQD7WZICCFvJ0mLauWbEHXeV3jy4GaRy6LGn
9An8GxZlBddiQAfEAkyMdHR7FkpmZkE/j+mAo1MLdsZm198nVp+9ySfHXx2PsM6quVcQswkdG+77
HinfV7UmiU3ZarCZp2AeZtvd75E2sPKi4jn8xIrqViAJHlteQuOx0h/uf957A0BBf2g3Ndtacv1B
76nhYKxlZCxHearEdVUzPJjSjZQrcq/rUyKCTAqu2SS/oaqocOnyZbuvO4UqOS60a+bdfdAlb3BJ
Lnj4GhjenuNFdhrzPBYT4wim/rAf1YOCm80gPEOZ8OaGg7lNIsr1UZs19y7g9DWUJ4If9IOtCrhI
yKc/xwpJ4yHiv3ahGDWUVw+3x7UJn/0yF3BOk1XbyD5y+pQXeSUk3vfFahvDDVWqts7GAh9Uczvl
bQeEILe/9K49SbVHbGSWDfN7kNKbgryPQ7E0j+nEGOp43K5WKP6fyTDIqk8/v+koY/J58g/YfjiO
SBygBji9Y00x79Zkue8ZXViSjCpltku1dSSUJJzr43NlYllg5jVdwA4gUaF9pq98iNhzOpz2g9Vx
56GjUtk2TiclE+NduDo0Sv4dfONAJTR4XrjR91s/6oAcq4PBWte2qvBBrERRcOcbrAk/mdPOiWoc
1soSUxApghksV+vdwhMKzcd0AZjHeupo8zjS+tX3356XVfcRkPyxAbzMTFxDY7l9bUI810VSQkM7
Cgd6GziEo25Nn9ODC60HWY/TUexK31DIMv8c85ClkJM7ZQ36BCTKKwIvWKMCnlhhCyPSYROkSwFl
BzptKu9pOTZx3RCh8r2MS8zUyL00wHwYjGNKNQadzKEtM2TgtI6GSn4OFLuXhWSOVvxYJ0n1UVLR
oz6Y21WNPuqYH2wlQQOCLSpZpGttNRs+emHFI4EjOXEcvroY0JfD+xbGlliOv+Qqx+RTWfVnszmc
xWb5PxqJkvQpz/XK8klni0d5i/la0edNpZaBIJa984RW47o4mB4NhRNsu7Jjd8VyOogVrqUMzhp1
+eDIaPHSqJWWs8/X46cQm700gplsomwCje7dA6SdVEmQpRlDreieJ7TVUI/1mpG6lvnKNAgRFjaS
w0qXnMcgsF2vE08bgrE9zzuDZIv9zlsZgwVOcP/3Bb5oRCf3eek/Y+ITdBX++WX6ofE4GLGsiypo
d1iAYUFlPa3jaan8JwGB3enU2Lhm7gEvO1H+pHUQuOxPJaIr25ZDFBHYzrDGn1BXESoUw2d7Kr7r
k3E5GC1rcNKaiM8F95tEwUxMJoapI+Ffo29hHzhFRlcLnTPvoDJA0lth5PPLbznhdwlY5pUR8GCU
1LF9FXDT/c7nju1XMnJC6pH2Ee0Y7rOfkWIGkjViFecFcfn0C6h2XFNSoQpAYGH3uZ0DqKk92QYc
o3O1QkC2SgBRoFD0KsqpAsUw5tb48ZlJszaK+hPq45Fip7g8xXeFTahJJxBdiV668GsJTcCgEncn
BbcNuj1diROxKU/pAitFBjJdNUxEUwU+aC4RLlY3fc7B3XISkmN8O+jxGAaDmZDL0h7nQdwqPOCd
5NL2ht8mVefK7/mLuAYJ1nfsX0dtdzoEY6kjMMQwyZIfwktuDEuT+DitQ/QKSLQ375m2b0PKf8SB
Gr/z0y9Xn4Gl8qbyFAFNDgw7pa2Oqbxld9UtpfRYvoa8E9L2kK+WnXThm9a3nGp//7b14jTxZPvW
UfV9Anbmsr++aXmQlIe68WprJtRXH5KXH78Si3aa1YwxXbxLdky+UuWBGFkTqL8rNhDzpKl2DW5z
oDgz5oT88m8wyd4/aHHexG2SSkyXzIh+wmXh1b6mlCfXfV7g2KpqfUTC5KvFTkTHq1+j09EYuZSM
jyIWaNPaGrMxWqx1TpSVHl9rgnHuYlQA/dzRJDFbjfpj7RnLAdRxcWgzP+TgIjQelVHe5iKN3BhD
+/ST8VKzPdNhu0aUVVNtjEOGukghiX7ZEUZzLfPWnfGtf9bhg93Jc8EO6exZ5NN7VI1vl3g8dnTW
krUQDTHW6yqX487jpoH/J5EJ4bYc51EXv5bKyfupjENB1kyquyNcwKt/ZCqYRm+HKK+Jtrn4QKR6
konubtzVG4aWBpMLze4et4OHPUk1BNgo8e5fdxBU3hGvVDAiDRlbl9UEKVzfOupYNz+APOFhoVNO
S9hPOTvq6uRbfu+VmuFz/fe+UeOZXBs3wfpb7P9IowLOCPE5U3uNMu7E7G+4YKWr76JmyxM0h67X
PXD/MGHRTwUU3AlNSrCLNGZe7nBCBQgPll733FYo2G8w/dqCcK3e8ZJw2k+Az8P0kWv1M6F/hCmQ
GN/J1MiGI4qwgpcC/p6t6ri7XOUQOTwN833MgfLCISDxSLFQ/HOJNFYYsqX+2+asn8vUQceFykHX
BX3N8VGT52adVq7h9s3jKkq4TvIKzrjtPFBH0UpRr9ItZ5EhHYEzmlW+Y4zMh7JumhU5rWwoYiok
FnNt+qG+4vlS8mf4BgWZlSjJZjbv0mjH6PEf4hgpb6mNaPJ+dQE1WaGDPeLk6X2YWvfXL1MuojZR
aSaWSishLXT3jihRo3XfFdpy6nW/DQg4El3/XqOhJxGP9TlpdwuhrojXIuoUt7em/4e6GpHALSmS
9OsZsUZtlfAyho55lS4gqESlz5+9EBbeq9C0nDywUV05k37Fi3twZaiX+DvxRvaMc/64D54wLGg/
qOWONy5oiWBauzHyk999LaiTH3q1E31BGYsfqqzWE7dgS6YtOKsHSoz56ZbivOjmAJDxGJfGecbV
jOZXYPonjI6CXw0MBcIjrgeb6RANEW0nnl6/zkpR+wdSn8nI6b6/HSbAJSEFKI30DxOW65FVqIlZ
k/HKSCTSsqsERrXdUICgTZXcuyXx59LdPdZsMVXKhHhVRnXj70JTVq/ezpHm6IhqSql7p32iXine
VinTN3TyRn4ciG+XzriXrExw09So2pIpNs6+czxQz3tZ1mpe2C9aFngj8qzNZOWQbi+rRUqAyvOM
Muz97Rl9A9lM+Rjib4y+8e/HUusDALngDOxx6TQd0MZ/rObABbKZICFzN8IDmjnMOaHQp70YcHHJ
tkSqseICyBVfYMYWyZxloLXxbutFcxDaS0mOjklgxva8P1HLBj5Ed7X5bhIi0ICGiDvx6GN4+nNe
AgNR3+ipIyvzazRP1HLUK/4//2KpFtdOUBI2L+GKZf0GaVZ2pKemfMUBVbvjL1UefpMVmmets/+m
QvLHl2QNGXptjNMBtSvYmaeHF+/0cTUPHT3fSUnbZb9kFZ4uozeIa9HUjXKVmZqnoqhVqP/R6PD8
prAMGStVh/ObTPjcHPKGmaBxPv8HZECby5Tbxx23z7UItqQoJaHXBqhp5RyCSZ9LSfP1j3QK8eOZ
YZuwfvAM225noi5z3uNQgfCZznHC10RP8tgT6fgwdwxcH8Z23YWyfYqHpoYFxVbYV1wtZ7aiu6AU
2QHU5gGogkzqDoRNmIPQV5NLhifRxiadkURN5LPP0HE/gyBwlZHvXQ4jrbbe4xVzPC2gopCitPfS
vWzwqwkU+/7wBqJagnWDPAqLjFcxiHYT/JRg1XQQxzfl/SuTW965wVslKiVk1fav0BYxPxoY+xda
pvI77PtXdWWrFy663xRrMsvUaza+vk6S7wVYInSbajrJSM0bhteDZ8lfVB+UdlbTdcZKewLuD5Tu
Uqta2z1JlunrmuCl0JFi5Cdx80tL5C9M/3EmxSSRxi1laRcQ3PLHcD0sK0DUMCTSDTJ7EBXCJnOy
67TmLVM5W2ypEHOS+CurahLaT8h0QXSJcsmxKhtElyccReJaCqnJU+ratU3YLhoSYjVc/YkJHtlv
pFwieMujo1moVSMiX0wYOaVWIUsooSUMCOP/Pu/oTCyCccl3E+lI5ejOeDR9ECRGdi+Id7kST+6P
lStpCFwlxoSogpShwOEoIGmEX0I4TS6Tw4Tk5Y0xWqBb3UKb+rZ+HUuTnyitGVJO825aclcuFw4U
+5nU8NGBk/uuK4JtTk8evohThtNwsWjlKlXShQZ8gpbLGR3Pc+pQaClfSNMy9vrxbn6cbFwVQDy+
D8EM3ScTCLAzT5pxVx/MmsRt/c1VECiCL1V1IdOqx87cp0keT3k5TGc25VuLKiyT1HMg++u9p0b6
7sGLFqInYkBL3E3Xms59IfN98udjvfavv3a/JMOnOI1gdkDHsBMNw1SykcRx09ft6dsor8aHXnBh
U9vTtboGoGF4WuEfQMrAHMNEcxDNt/FNtLG6B9UojKP0oSXI12/NnZzs2dnS1DzA24uw8W3htLkb
CMbq80wUvkb25EIP0itDtGIx2ZNFF2yFJ0o/iIji+P5s7IE7U4vdSb/Hv45ncx/WQu3T/hid0Ob8
ZcEemQARq0PP1zX/l++jkDloO4C9SQd4hqyXHjw4CIi6WLFwuCyzMGyUD9Ulx7p94ESdjBNkaYA1
NNx+O+g7K0rX6IkzU+emfC3/sVQWXtXVSzWoUKf2cb7ckHwfTTNB90oeCHAFud36LQcpz9L4T2Ke
u9M57szwt5WmL/xfV6v4Rao8c2iHtZhG8v73cb84zrFr8H1y1y4ay1qK6mqZBhFzUFy6Gru88wTW
x898kB560F9UIlz+Ujkn8abuyLzZVr+QDFtPYRlNrhuxqVEQme6CLZQvywoyvc/X+jicq+KBBjQu
IP1cEkbm+zbtxMazErigzi6hiWd1l2EoyaMJuAXgOK8dUWhrjKCnALRIODFC9FozMyowm6vcRUL0
MGBoHyGWmLAUiK+tfj59ZR427AuDVlUGuWhKm+FQG9vR0Fs93ejL5h425/eIVyrkAjl8tiIuDxax
36qJ9n+Zq/7a/bKoaAedI6LIQYUk+caPUByIhuilgu0eiloo57Vesn1wRBLuNZA/zeSS9KNzY+Iq
1JDRR0u3/6qhCrGQE3hwrzW69BhGRQTbZlbFKAbyD9NqmX4ptFq0FrKhZ9/5pYmUCbPeKk0wedGH
m1/z7OMFRzAf56whQyxFCwGGu51ylxdyVTWm4Mo2QTHOMkyR0wgwctRhRHMnfeX0WvEctWN0NdyY
3ktTpXP5aCBXEV8Pbg0TJ3bJmRp5TYsYEEfTq7KR4D1zteYXdJBEN22BCFAyXnBDvj7Vb7V7zizy
6HEl3RbYM6pjnd0bJNqIMBadlKU0jqGmA8aysN+vRonNbSy43GYw54SrTgn/rWthyhZGQUdgAXCP
v7QmovM9ShIQ4nNf/NtcCJzmmSCidAfOX9UZJbiTxolqg6WhOTe2CuFetrnoidgE9jJV1f1yNOXP
fuw8ackCZzrB0tPhMlhT3h6ftsrq4a/HaOs5JPexZ41t3y4Q9yj/g15Bp7AMA0FPQfjM66PHKyNt
Pn8VLT+ckjHTrAg8hIi7n7Sl0Ur5q5vdwVrXMke6SFuZTBwZ7J6VqVACx+pI/RJQkj7IDj/a3iPk
w2b1uhI0G17kM4ZRh3v8QLWQTTI7V5HXl5WfbxiA6C8fAw6/Vgd3jQWj4bNIHaIPuuPxKJ8Ncgo0
iO0HzzvvTJKDkiq9G8jzfQPSju3tnCSs5dua9x2tKB2WWGTu2WUXLXKDXePJeVtvFK/HVbm/9KOz
xeMgGASCX9t7staKMnA46XnCPcxJFJvEOO7ZUygF7EQo0/eRD/l/7TdAqN1yOzv+t3sHDGpEW28b
00wQ8AWD1rdWfNgZVL0Jz4Q9Z0Mrsma8VbiVOLSiZXvHtWkU/UtsuzLIPAl2Y+OzMXBNXxScj5Dx
6yqa30RQ19DUL4FSBbU77kWeCrlG/UFoYGGZpwN0oZ7pSAXWUodAlWYxTIktidmmrQ1juQudrqHN
g1/GSqMewhs019MlePtA92hOdRP/Hm3aWGygPHYmA/F1drQ2VkI8L3xUCe9BDGsWKjXy9/Hcq8NV
hfe61VcSLUvbUoYEPgrKCU3usPCNTlQ0/UvSj5U32ZMz8LL5fkZ0Inuv7so7HN9BWGz6ZAygihF4
Zy2WGlPEiQaCr4GJFSlW49wzUPVsbudmGFdWq9XwquEQ1qQbyDsE3q+/OYrdqyTFxCjk7DRSZjkP
NjD1mS1paQKgPPNj70gl4iCi6/K/CH6tdqK87pcTo4F7A5m+XASgN/En/PHTsgRwkeq3ALUE33oc
ZGgK3vxopTRQeWVCisQnOu3MR0URh2T+IC0e9AzVS2zGHaZ5G25816m8h5gv5stC+Zfnn8bwAASo
t1IHAt4tw9ugyKyo0Zv+uITtuQO0zq81mTe18axhB5CO4TLI1K35xJdFVGfC/+pL6qrf99WsOA/I
b9Xi2qhtrfAJ8K4RV/MS1rYO4XbV9Ll64ZqCKS1TwAeutS1uLXaxqrDlfZS16lw2fPe01rB65Dwm
FvlCHyy29tEHiYkl/0Cz1SrLq63ej6QeTSKxn4HEqddFvcYtxjg/taVV83ypaaoTuNE5cgIIvWUw
/ooyDjpHyMMGsTkaYnYmeQ/EAVG9Qv0tT8msyip5tpTAF6WQgewgvdUQqyQsoa8kKsCkEUWsKwdX
oJmr4nWGsIrM0zdP+r4CSR70rOrrL/mVpXq2d5nX9QnciXfCTId6E83+4LOcCRZ3AtklCVwho5t8
l490cnu2/GxC9f9M+tm5kx1XZ4/qt4q+vNyeYfAumVPB34qwMsAQCFzgBsalxWc4xC5o/iRwKU4Y
3Zmu1FdwOPYjcIwthk+yGOrPRhWqs1uNO2xBuhRrwqDSZ/+QV/q2k2rbdGB6tICCY3kgrMuVqbII
ooLVv0jyJwZ04gqS3eS9oQygvtv2PCUlxis9avd1RpiWOjBiL0HZLRI5vgsHQEpKmu0gi1Uj23yw
Opmi2aBtdfd1+UJdyI4CLm/uncTiZ7StWMygVtb0cZRTEyV589jb338xXv/jVdgetmscdhVDBJ8R
AVRknmVguVeone71eQ1ulmwYW54B2gZqN7tYum5IIruPIhKtaBzgGqwwu6ikQrc0Q7wAVsMuv4Xt
X+UZ2T3Hm2sAtrusem3b/JvR9jKHpDsp7PZ7/RqDvln7cnRfhS77YsB+SWnseoLg5YEHsl5WCLNW
EVLEANZMgMWUij20hHKh3D5/S6KnBDKQkmxWQ4NYUikqSQfZK1pUs1ko+a9aQ4QNQeK4cs7E7giW
r9E03yWvpI8r448ScXe3v9W0MgUBvpdjxJYaq/Byg9qa11Z54f6yW7467fSVoQbWPEKbLbtp7wGL
+5nZlVesYZbkQmpkGUFRgMILZgjXYVkvvAP+582LHCTs7SoHD8rxvarSmL/HevVZQHNaHXO6NaSA
4JOrjNmknSsQc/EuyT7oW2b2cVtB7kwV87XWUaeZZ4PVqtcSskycygXBqM74ONJq0ZOnFLMDzyNH
cDO0oPzVYjh5phNs/36rY5Q2ad6wQAhh1Gw2crifM5A2UxiaL9UbKm6SWJPowbLahGofl/DmNUr7
D+Pph1+YpUJmeqtwLyevOfwCk/HU4eGDC6T0BaqGKbFLca3GG0fD0KWkmSs+wc/wpzIb+bIyMaSQ
iv2cjqU+dKzpAKniS7MLQrh0Ws3qj1RrSEGGBuj3WCQXhDnlJhGv3/0tnNNydR4N9XiS5K8c/a03
ccq927m59NuTKTbBbugzZLJBqUYTaUJNuh07yw2zItJa47GwB0P6iJmgrgacvAUpaZmmSAm8Vqc5
Z4QjxaNRcMgX8ErVV5De89qXomaWYg+r5chuBQMiUDm96EBpJbrbaMrJsYbEOjgvysZkub8SQ4Lj
y308o4QKXddWZwwAH7BnkAARCgOXRz9Cj5JEPBCyPHCMgaHRi78a+ljkblr1+AMTKgd3kpuefhKf
Lx+1/9xEYUMEoEVNbq4BZfqnoGh8ELVmZTq//BMMQxGH5CR0QOVYggYJO4CNC1tr+ZU2QOe0jWAg
tkJMNNMDW4qcBiQmmU+D0OlYWRbnv3DzH6vmuOHk7viyxZKsXHK/TC4uGD1L1dvJzp/7Jw57w8jH
Lt2UfOqz8Lstt+TywlQ04cEPPfyOMG/f34Ht6EydIZnwiErG7DHdP1MkXwXTz8Xpv2BjWneL1rHb
uf/yC5DcMpFs+axfOW9RsDqCt3ejYn/EVYNKls/7uBrC7cR/3HZRiJrEqTqFw+BIX0ZYzVxqPtpj
qw9dr4EybsB6fT8GnzPFt5CBRM/TKwzcEXtzqbRcxabEGqv6oVnOGVqanT6honAQ+ALG7abs6Dy0
47Zkoi3dTAvQKuNmw7MTrtVPeshRNxBo5WWuY6hLYhS9pDWz7U9B4T5oSIYKWVt3pbUk12IWUg3O
2KpZGf+pcMoJgiskde9SY0eENXuXSWFkZv5fqo0lN6rIFEz/AcetJTXIf4boSoW/nMta6yXaZ9UL
I4d9hmEMGg3JkIesCuL12VUagi/a3wDhEr5ahlnz3HL+kiiH/8fltnzaYEL/fLdab6zYxxoyE0A8
7XejQv/XcABvUlCC6H3iXpTh0DbzKoYdWcM+pFY9dLLDaY7+oTfd/ZfZhGTSdVqHQAsO1FeEiMLF
GuCLHYU7q6OxUPcoiaF+5GCXjh+22C+/3rl75NHaU9l21FY+TUQF/lMasWsiImbZaKOo1JvqSc/y
KRJ+FFVFCvNVpAeUwu+PEIIbhWB0rG5CabC4Wv5IacUrk0GLX2ioehSq1gGAmzNI17ePD38l+JJE
F8znimyuCwQkrnofM2nm3A2bYHuoG9PUMtg8pQXRmMqxr7Hh6/V/VHB+TaE32FRq9uzKj/X2wwwl
YtHKhA2AoZCvB1OaaUKycvfmAMfNyiCTxPGPuhc8Ry+tBM3k0Hs8jKTjKUBS9398j/CEADK3IPIZ
OmPMmYza9CcsXTXd5Ah82NsWnUv2llIe6JKeo70yI3z9b3jD4lxa/Ukhc8iuch07rqaLJvAd37Fg
HQptLaiy6FPg5gyqEgU06xhO9vVdz9IjVzxHQHcyHG6+ChPu/Daj2zownhboYoOaXupV5BmRTOut
eATrno5jDZd1n7P+yE1VeCatIafx3iIfa0zpTEOWzQXiRrpuYE/+6WiUwjetd5rbqE0ya87eRp65
oUpISrTFAdVpTCN6kXvTrEWiBdY5oCltUXDdzzy8Fwm68zMOWG1VW6cOLQkzsuXZwDRexQjYzWQv
6dVZHQyNVp1N9nNeeiOWOCIG1SnB3SJsUoK8I5i+fKxjInlq3xzVUizSMcc4szMG5TYHqOGCM9mK
cbLf2S3rYJ5UzwBwhP56DQoWNUKHrHYNwKgruKJXHw6bUZkc/lP2Y8tHTndqTu+IzS8SAwxcNs9j
ujm1rfvUauX8omKYSfbfnXIa/PMCVexJk1Ag99FOj0613ybtpEzwya05TjWjKHnjDhd9tyPbM41a
VHLVZ7ioog0TDpZ4FyLsYCHC/xm98Lyp6RH8LjfDeFsabkuKp4JXKPHJPeqdltO3NYK4icD8bEfT
RCPB4L63el1L0l1V+tNNWY+TjMRG+vmcFS6MgIT4+/76sl8Eypv0hgnw8TqQJHY54t34FAsIADSf
2Arp5/H+sW8gKqTFLolpZxRA0WxT8MqRcJ+GMwPN1d6KWIfKYLGH5XzoNBhaeiLndLRe0xUyjo7B
i/GFX2rJRApJvj74Pe9SPtZJRX/L9/20cWd6ygC9bpgV6zE+U9ZvKPdq0i+60JVVfpjlZSUN/JLe
pnOdq76mxxZQ7poyco8jO9P4f9WKJUQuO7Etan5Jz/eR1pPTtVSBrKlkY7OWCKuJEtgU+PXsZogT
lsAtgl3Zf7i/Xpz9fs/+W+e3KWe7IhDRvWC93UKMMCWBAnQxdaOjStTghx3kIRJmSk1nGrOoknGv
jdn0kOBGw7mddPnIR/tk7THJzqqyJLnRk8BOsfjOTN+DfrUvdIQL+4L1zIMFdsrwBRqnSU7eQ5yT
jf9wJ1l7JwtFPGYQxf7fNWm3luo8wuoVbtSdbDp2LQ2bpL1FTuaAzhj4SF/cai3lu4vKXwGCsJQD
Q1O7HegMa3dfXyvunHbKrB1dzdvs11DCuhwdF016XhUN0MMTlcVAbfacdIXj6ExHUsPqTEFJN4BV
cEjO3QgiEUWe6nwCBuOXNv9TtztUK0M9ofyWQDkCY2V7XrmIwmj7OgTfLAtyjAWW7k2Xs0QclMx/
McYKDHRhlo5qlQ+JiBSDahMABdg8ywrQA+AHC0KcS5jb0B1G35tlbBvOvIF8C1ekXpP6AkJxpBEQ
a4MuiMIbawhOhshtJp8kQ7AsMCW8sLog+XFyHF3vhNa+E5OV1St4xICEpJ/TL7cw1IphoaOy+kRQ
C1qPzfc0GH+wfic35Ffos7t49O/7763MtvpYKwpPUHU64SxJnxlx1BgSjZDZfhvqgZF+K74tDd6m
7qGsc3p7MzZIAhtcbOLmRXHPeek6VLqlujzR0le6fk8k2+WNz2miVmP6OlAkpEyV1XBZMWtlLtod
prqG65umsgqTQnBORcqs971PKpYquB3j0oGt76bEPYrmuQ3LQ4oLGbgg4rzgDQTLlnb9Wl9krk46
ryJMTVWoY7G0uJZ0DpxpVFUSjfKzleJ4Qz1nNE0ggLxEnX4JdmkvEft2YuvjUihnOeWXOYq7jK1B
QcT69N/gg150H7WhGouKmV7zktxr29uIOpTNvna2Y6XVgjuUHOdkRyRkGh3yn7hmIdwAtOoPSgdl
PqRnNYKWseRRZoG65RLzA/ieSn2EAy6y38jAnLZnKHmmzspb4+cgfESVbBwedwM4LkMufXUprYow
zsuedswpZ21vG6lPyzaf8U90cG9UGIXVxRZvMc55sYbmp37i5SrutPXBz2SDua7tVeRwmZXcaL5W
xdtRs3BCGFmGEtRIzatSh+W60tZHCHhJiZElCdmhKaXRkW/PXC0FO/o5OJZncA402IpMawieT35o
S1dFTlMYqKe9uZ3q/wnEd8Yb6Hw1EXRT+KGM1Jv6i2XqHUcIqq++EGegHaIwG1AFLywx7opTvRc8
SpwvEMX4DFxKnqIJSWfmL2RKaAOq9HcNH9k7zXJ80ZygM/wNK55hQ1+dVarB73q9oRbSMgxBVISZ
SDH5ydzKXC9Z7RXeUU4cpCJHm/z7I9TuMaxI5intRE1FXhTdp6FKb4ojOG1tOKjCd6Dpdhgcs27X
O4H4gDML2BJ3X6/DDslX/ERjAgTYH2DHMt/ofOjFnmcYBwe2ifAvHbLbQl/we/XwyOJfNcvS7EH3
f70VyXisjUHgBxstikayzGmWOS2YKjWHfbvM6TRrVAZGshclRd9kF2IFvfia/FLdrCIhOo9Ba/uQ
v2/06DOLv5bo/IvXMZ0qt4bWxd6froj6/2SA0UnGFAPRb4Uk5G7cz+gP1hoA8cmIbxKqzrDNY8g6
lKtidEfvPKBHdznXJF35MAdF+dUWuiHUHcfTyXeC2DawBqdK16jB+ilZ9AzC2MXaGmlzudDobyES
sK1vfrqGrJkLDuMlhEzfo2843F6c9HGGFu3//iJP5cWqGAUodFULjIQr80R8Mj2PnxXlsZVcGiJn
WRmsjLm2CiyLhxIInzcaGAuNyJSmpHVWTh48y1NjPqUcWbA1jsKUvPFe4AOyidW1Q0WE5llqIrH5
BpwFl+lRDhJ919FMeWcyT+8wJcCXEqgynEgvIhcb1bhTK7cQ5Sa0s2YeJpaoDXHYEo6HaV1EdNjv
wzZ8oTWFoG4UoW4r8BQzxMklPr5aoBKt3G+9x2r0HY1P0H8TQ68jTSIb+0vEGYLItXMp24CqB1O5
0CGfRxhKuNuh+tLXXqwCCfAtcTDNAgzm0S1dVObKIEsA7sH0FDYwyi6aJN9gBWNNP61PPoy9pX26
WpeAnSNoPEZ+hfsKXnE/Ok2dd1CeqCXr20kLp/TvOuqVRp1Pj5IBJ2TA2l3LYxLD6ONsJyyb+m1A
GgMBCrWhToo0dD3PyYcLf469E1oeS9PquZzpXPQ2GJhh4RWXkRm0xyWMFI83MElewXn98zcR/PEl
WHtQoroK7VPt3CrSSaiBQfTQtmMixs8gPRz2PiojzoNF5LBbhfRX6AOSeK7ZAwyz/5wwrDJX9p7m
cOiAej1AjDjzio1sk5AVFWtp9uGWtqsr63CB+4r7JgT++g1ljoHCrP2oxvSvy81i0ZSyi4za7u0f
gSjxnElYET0Jd3DksiG6ZPLvScRT+x3FxMaWMer7Kyd6XWm6tZQrPebtWHnmb7EbBKRTcoyhLzCo
Nqh++XDfK1dxYSQ5t7aPHFj4xrZg5htcrKZevKA/FaieVB6pdRUxuzfpEzrzdynEupOPvkvTvaeY
Ce/+gqsQdoiEF8F7ovMCCAIVhr4SYNPyOFHc6b788Kx6kAE0j/cj79nbDK66lHYSha6RpgrU/xsl
wpUyWKxVHhHuXEG08+lX8pAoKrIuohMZTjK2EA3/H34jxWS9CsJBkh6pOgtCT1kB48a9N/JONrVT
S45MYxdIN/N6rIg9DV2iiKpDaSx9hJ/rQks357emZ9EgIFVRVFjn501Z9dOBc6UFdnvrjm0BQNu1
9JJFi/4+wUx4DLHNXm78C2jVd0CefTFD/JRtNe4HYJbbnvQ07nh/NRaMpsG0F3eY9IVCHav0XLL9
KyEC7blYe1oxl0SDF19uQmuLCfG1xmX/QtOI/uzPdn6N7BM/iInF2ED1CtZ3sKQ9cwZ0qyyC7iB5
U+KBy6cZjmU0BoNMlBANEJwhufHZ/rd4AfcFZVS7TX2ImURCe3EyO/N6vR5is3QIZAx8zfNy/FxV
IjcA7/cF0m40qbIk5+hxAWv5lEvLAXswWSQv8UKLaumgwcemhKOB6rzS8buLu/VvfkLWqkR28V3f
nh+ws74Tr6vO0TPWFyaizw3+dXQVL38Ki1SrhdTc6kQHATqpth3mQTrMaRCbgjUZSDNKgnh8+bTR
5RjeUcg/2QkGUCZoxYOWl/QLJGMhIgs9/owjWocyYxx5nghuK/p1mmb8aXCl4IEhsmP6QKyMWBt9
Sffklft/Fnp2BqBYt8YY1VI2lU6EgJoywB3uLeHMlvBZxN8QLPYa4wcdMzhlNt/ngV5SWERMu+ue
7WUHJXNUijf7VS+++PCp6TK76YNdK5AkYcT+bFb+Hiss/7Pc20L2vtm3+29uP9GR2sbLs3yuqpNG
c5Dz32455mou9Go+/goENu4XEl/uyCLY6zqdtbtLSrT6TqKVqrCct+6FxvJQZPMmEimMqbkPCAEd
7BF1fqwWojqo6OTd6Nl8TEz8jnK1X0EwX+4s0L194zaquh7gStczqCiyznq+QG6JMVTowmNF8aRQ
MxqulZRjCtzdIyQWyVDDnFsBbO7aMZaUf/0r8f1Vymh6FGxHEzyLHFil8Uryk7j/fKdg9NbdH2VX
5MWGe6IjmGbT+3DFViSGEJJlNgf2F6hWve9fKNlBVR6P9v9wwFkL7muXvzRtIrJS6o1bf7jY7YYp
YdyKfCo0Xi1/KJ9ej/eOltg226PYqUQDx/wH5ECES5Pzzu6BehcBQXs+xGLa2AzZ/Wv7P5HxBv0o
5avODDxy7gqaw6/MtxiHyCjKKM7qI1rG8L1wflWGIBv56LVWYv1uJp3KsXYRp7Xsk+b37Tjfgrq/
zhJladQrCVOQcpa9kVqMBtcfOdruJ4PMFETY0PKa3fiJ06/SwXoMZ8+eF+AdIM9qqKsfra8rnaZ7
UA7PAmcAqnjymIQRRLKWsgwMBR3lxXEUEqQCDLL0VeaAHE4PMXz7X7nwUwIyjqSDNe5kthl7njgh
8SrdYcgjnmOQTEDM98QqTvY/SUwMi1Dt7bX9b7dFdl+yB/NXFZP9Z/g18lIGHYd55qCNQ0qaDnTO
+Ikbqynf+TchvULU+JbHKUXrlB/P9J2kCZHMefghueXQEAUn5QCWGnf8oTMBie15dvG0S5afhKtX
YT5PF2EEdtztF4g7Yx4NlYnd6uNkAykTplc7Z/RfZfXu4j+gHn0sViZ6UPJ8o8uJGhldZ1cVJMTn
qRukVwGQGsBmAgvcy/sr1EM1KYm1eZwQuuCTc1/ti8UJCYD3lyUEYCQ/vJX6mRw/F1t/JWV9+Z6N
rBgjFexo6Kuhonqu64JNJ7DfMUIoGQGnO0Fd4a/E5NkbU5pChEjaaxxNuXDBq7MWZ/0MqWPA8LE8
NxGF/LNnP2hdCit9hwHdR/fYKoy4h2ag0cme9fBqc7YfDcxZ45hu6Ck13ErrCjb7v/4Pz3LrmvF1
sxA/NR8hQzo0EGQEtfORMmc11H14aL1gRdBapvX+Yn3udXZNBdW6OiiAt4uipOejYsd1jDdD5wKB
/wVYBU+45c7frp2c+HFcPlKHIhyHAzo+vbFHNtO0iLwZa9dXjOyaVb1/hJQ8m+pVhnNQ0k49634x
kcETGHQNmJVYx9fuTCMvgEDL5ySKwPO3ueyefWYYJSFNs2Yq8UK3oVM6zskv5LPl1UYEQyRLl6kS
QfgP8blO9Dg9xkdYBg2G8e8spRuSAdgu8ErYje9BpVsvHkI1FPoULgJGfCLBzBajSUgm4jVAxJZC
zdICmXb/6R6ke8nzXWM5iq0NRFwl4owr+jTPN8FB7z8+Pkue3JjBI5pGsID3v0bSSG3esoQ1TMVu
gqzhot0MiUl8F84dH7Hna3YLdSaMwL73o6BICzmHJnH/N1IfJm8bMPy+XZ0Z68ZoFrUUKUJcY5ZG
lLaa36lFbhCt+un9JWTm/7OE2EaiWC5Xm2QhnXxiZ80Jvu+IAs6PRkbHsIqE+QOzPYuMi0+DgPEV
x3pLPka1JAvcRHcYHzK9nyCvPFma2fmwX7wkY+kQJYBabzAanCyRG7zPj10esO841uF49N4aTGoc
8L4RH8/Xa+dFBSq+bLcoVORXAzivpo3e97KKViXHTBlXtz5a9w4V+8C/uFU8P098sx+QDnP6Kod7
6jQHZ6EDGC+WgrqolnP91zP7oRRJa22QJ4+DkU2v0XG5gxaKyaIR/V5bO1sN2wQ8cLRUuBQ9vQ5L
5RcBAHfkEE6MzMVY3n5SPPrUEKJJLJOA9vq3cbbATL1x3CA0VIFdvKa8d5Dv++RVnKz+/ThT5aJm
wFAXZb9c6K8Z+5nFLChsuf1zSW54OvVcvhGXIV3fEGmvBWYF1fto+POav+K/4QPkVrCLsZP4+ULZ
R6Fm3NFnFcDL97nPftiRTvJwFhNlBe6dFVsodywYGgf8sgsN6guXQCuJfgMajWhs7XniFyZHhdov
QC2WuZzb1KMf0u64JS6E6m8Ff3tjcfhmLwxAmz4m47LuMRI5DzsZIJvKA3M0lmGu+ZNLWLTttGNX
ei3YiMnHbIjvpA6+H8nnAsb/IEk2N2dREn9z6c5DDKd1c5mBuSJCuUQ8XDT6Iq/kpTlmeplBQo2Z
DCvqTI3NmstuJBQWwRVNUw03Eo/0yXhAseCGhx7ohTLJSS5SqKjt64ba0MGG7CsvN+ivZALvJYZP
77dvi/1gyl3Lil2B3xtkh1ydIt9vJbZHZRviJckhUNkqOCSDNqFxMd7tezLKXTpo0R/sabHK4Zqz
rxJiiY4x2Bxd90xYbeSuOlf+1H9XR1IY+3z7um2jjTgp4pxnvtwCRd5hlzv/znD4unPzWlhgtEuS
t+w8BFzhG2FJPdjnegqY/5WLVoDGi+BzvTAm0+QIROtEURv92rndIYpAXfNkalncq/SzBoqtUtfK
UdOTAgQ6ZXepPlBjcOsuf5wqkjDWvmM8MeL4ekC+pClfaTxQTs72f4AiMPFV54PK6nBXTyEOp1HF
i8RnP+MbjAWKUYhvjcZWAECVQMucmYNxbIduYbhfoWNOFRbCd7RItneukMKAhzv2+nkqD0itt4D+
VHio7qWiJT4qv+4lgEmbMZtnSCdhFyA1ak2KsWFI9EcJLM7DkBdH55VFGn6uRUhJulmFRKGxdeYf
Wl+8hyE/VMnB0Ryl5hzr/cqBWshbnDBO6fKoZhPCcpx0YAfGtyG0RiL+3cb0LwRdfyKXuCi1qSP9
poqReOoWWn0OpD7H1ua+eMpbiICzFkzdOJlgy54Jd4qGlRpc8ZFNNIiI+Jae7pnoLS8FbzWwB9S7
ftlS0NGtCNhza7acexEGbZt2y1M2q6fLHeKT/MfT3RAjlSb4Y0ZWLvAAlJI9M9jxPt6RAefvat2i
WuF6HYQB0eGINuPgLi5oZFHpgjcEmtI2R8LlfkDk7TRQ3r6Rt8B2NkwxOwHvTPxZ/tkWFnDzekuj
2hCEebC8iA3njEUGByEnEm5zaKaIOblRAJAMoO+AXU3AySqhlyjvdxVn4mPNjQfkK/Ymz4pOY1GR
9gnv3ABEcxV7unzrTKRxi0KdSepKqirf+ouEsUtnthnEVmo3g0bs8ku0FnvoiO7P8M6jDvugtZ+B
Re/0QXYbPBRTSO//I5PAw0iFUZ1+bOFL2h5kdA7gFiR/GeVeCpSvh8t5iF4BlSier5N8OTn3B0cI
x4kGyJvw2bmuehRyOI4DqbSVt4lNdRYuWXzBYAfM/BxfxbsrwLlyGPcogF/2hp/4r/EQYrBnxYtW
1bXc0KhhPqnZWC+pAuzGbgTbKAbpiBeDea9k8GJMei4GQXiqHfir03Y+KT8zK/YLLE4J/LEc24x+
Ikq48CK7aIBhDyLqPj3Ul/btmNb3+ivZZqCGczLpIVll4vHSXIrujESMPuDCX/aqI38IepSF9zq/
Sm6fovJSgMxf/Kb02ZiEW2vGMsw/5O8MBN0nLZfUEn/L4zswO/WrmGakAVoDi5lXlN58zztxs17H
Udmc0TXuC+sYaek2Tp+R9W0TQlQE9ajLb4Oi6NO4yOgs6tTTxdRyIFy0W8RT7UnnBUAGNH57Nw07
dnV8VyhRSaksocfRFxN8Zh47z9IUYCWFakR4dC+1OjdTOwKNuZyMMtbOEl88rn6kWW3IudYJ0tGL
fkjzwO9JSKArUz8yUtqiTH40Co/6yeinQHbYkgtCyN7z+PtO0I+BlMyjTJdFODHrNqJvKKmup+3j
eyJNqa8Jtkjysx/3kYrv4CdkEl/eT+JYAEj1MCVLAMBhtlonSc4PK/RVZx3w2SQkLXiH/j3wK8UZ
eXMYYtRLnRK0nrxkRvp49r3vPfZWndGdaRwVgdgIgKoUGutehvWN64em3wIxpFeWB6ExG5BBXRBt
L1ieiWlEu3H2i14+/wWESuZwSWozgTXEPVWq5pYTrXBINvXDzckxqbOAq2xFrihXZi372gpZ3OUl
+dT0IcCmqA0AZa6J4Vq9+8VP7pHCXDNJA6ssFWcD47SQQofr04o884zb8HDTBBteiHR6Do2m7Fjp
IrbSNx9X+FYw4MObykyfuuleHscL2+s7S236lJ6JWJbp9rdle8AywtWODDHbSLAFdLJO61XMoLG6
PHMPSKsik7WyfjCvAVIJK1eMdc+PZsIN89h6QsGiosS1LkCEEHSkyqNLuyLSyqkyUz2ujgK9K5Rh
WqfwYjt7/UatfMl335oGSvdgFm24ZmCwOIHHUS/ER+ispCgDDSpiR0MwRuqPpCtwrf9LqUuq8mJL
sdvIkfYSsHOKt7OCU3yOKgsg/mhaSHlt3Pb4b7LM1YBR4zCBtbeEQ9PMgnRLMwycqAG7wQWGq8to
uX6m0B4ai/Bxh1c742Il7dn1T+o6gojqZLUxbDzdFw3KQEn+C3t8pMD60qo+NpR0r7VYf8mLhMne
DqCwGHIC7ui87xg77Qufy2bB4eSxPo8zoQNoTmXrm+u/ckzPX7Wxxowrx4MJyRFHtSbz94jS/xjG
9wccdceSXan093cvw5aiEfuOx6J3hOTNRwK9wSFyAKVkC5ChqGI3J4c8CUZtqbb/VHxx5HBcSsBF
TCj/guRwtmMnix6JWiOoBCZ113GixKxujtjEDW+DrigFBM7clsHqQXIxnLQ2vTKRj5QsADDjKz4u
UlySlGIBHZ6ZJpg3LtbsaMNhzFGhcMc1aWKYwxhFlRuMfBF/+xuPQrRaJC5r7hVqn12ZOmRBnBns
aQ30lEM6IevXb0I9y9MUvKLTb4O521GQg4FHPYgb0cF+uO6sJCeiUPGuEt46fQbUfTlXq9GASpef
lXxIeVZD4E97j7RZg7DXjL0mbDO7KHJpc1j98QQhhT4UD/tfqu5cTz4gBuSw7dzH9RiJXHZtqLEy
5/hcdGcKRGa/7gKx2/AFT40qFm9Zw23BxohHZfMz/LyXBwVdgQvXliirb9UhJhRTIU7xyTHqZp7t
k63Up1KpVzjWjczHLOLk/JrB06Hr+kOYAdKxHb+EOSYB9jiTAbFbfyfge+E0zHJnx7UMt0wsBxhG
I/I8abzCbTrp7/8MyoxurbCJxg82HyUwK0ZQ7CbeXuie6SHIXkaALCG9m4yStg8Ie9jvDwwLE3uv
aqfDxKcuAxo2nA6C+SqQ1kBYEut7jq1yz3TWawLBXe0N9jIw2t44cf/UROcS/T9yHXbshV1uQf46
zFqgW0FHLgTCME59nL++LbXH4Ywcc/jDeUDLI8pen9R3V4Z7SDJNNMJRJoRzVrLOMoLbI6a8VO0A
qF+Mvam7qXzMZ5vnHpdlYWjX3JCthXaHNNiYkVHJJZcTBF76eN5yY5DY+T3q+53WbpnkqNHbPeKt
ryuBpLGhGROvwRpZXdks9NmVBHu3O+FZXZOC14RaY2i+qxcP6+pciwoiCH+W6u4JbqVj75Iy6h1E
K0VWoAEX2Vu9Z/8AVssdR/CfPgvBEbjX5n4gprxBmedGmNdTsS5LDUfa/XP+sFhBYdIu66UxfcPP
srucqCsJqY9HEcRxwIA8F40Qzn+rgdrDAzqX3YsM+uQ9NDEkL0jpRRREXc78IGSeyjJ6OZ9FhMXb
2MwL6zFWQ6EBgdmwRJnPYjaieNecP4Pmv3IBC5j960H+V6qXG+PtkfiAyY+2YhGzrkoIcABXLKST
BCeIikD56XeLyRH6bsZZebgu+UsFYce7pnwHyqlaGjVNhF9wlk2HZt+P88gVS1F0JtE0T3g7Zjo7
6F8SWPoUxv3jhBCcfsEQyeP8g3XmVfKGaKXcm7jS09BwV8SoAf8CmLwLO52UXiKGPelEikBcXP8b
AncvDzNQwRAkVxeBLijcHjneMPennEXizo5GjoHxAksVCfppMSRrjnikF6brWmZRwBty0ZUKB5SS
g01FMgXqh7BYYMMZ2O9yfzTmnCr6DG2y6TuzKxU4rZGj1Y5+JbHRBxxlEVpdSF3GpTg2ozxWjima
LqlFQZtcH6vck6pK4LyhakqbGpLvm1Vh8IEqdFTwmJhg/qkuqukM0VxhxiBlToivJHFdDi5NSumb
c7HZZ4cDpIBsaFcenhDzcvQPyCh5TtzYtUolIZFEL2AbdNZfTnxBqAemBv1XCoyFf9+lvF61CgUx
OQZPNplsdSQSCdGJYS5j9rArjwsMweSWP2/W05GBKjsec+1I0RBvMrQszdLASl9wp6ALOs6qzk7T
UOMzd2t1RYN06aP3HhOmkuErIMqw9esnR6gfXvQM/tzfKAX9ZB03TH/mYf6GlH0UPtMLMRhTjitY
QisvY1SNrZhnIdsVbpKmbQ16oaGJeSuTJi/h6GszWgS9U0LdAsZTA10TOmRQQcoPo6lMPzd5Iy0r
dMoOXZWImwAwax1YMGIQLd2b8UIIqPbaEvc5u/o6721H2qNTTRRU8Y6cExUq0WWx8nTtZ2EAYHwf
uuhzKr5H1L8apUwPYT5zvciVooIZZBVyM0tOscWjFiwR/dgyyE27+LHObHaapHSuEUt23bxzBPxl
r0TnAGDbAk2bB1YvzkmVfzxk7v/wi1R80XZjCqsEVVJ6BVYmOLKZt3HcYkA0o85Ez4aeI8uuM40W
SFKKinn6D8374uxFVnpGSR3L6J21/3OqWQqmVPt1qM/PsLA+4MA6o43sEhqfYpBmHv4/ynH/lGWC
dCFX0smCeXlgG9U0clJeXT0H+FgTQUMEg8j315djHkMazxo3WUKwjHvQCCD8zTD4HwQ086AvrLX6
BOP/YNhhXeBHtVlhZYCpSDyVKAcPcEyVz1TweuVcMQWvPziZOSrkSoeErk8s9zGgwD+ZQLrgDRxQ
SZD5nhpM5eURxq/o4x8Cqv2NE1FM4U4BPkoCo99dl/IOPhqkQbl/2EDie0HNCS9mVeoUEBE6lpbW
eaK8wg0EGq5yWF/bpZNWmT2UlmrQKBPHLNkDcUvbj8/V9BTTeKPVZSPEDshWINL8+EaHgf1XBkhr
xfhxJehg3a/suj/novIGZV2dLBLR8+JsLWG0zO8KSwVzeqa82N2n6zde2m23ZV/c/jlL1BlmpeO8
clFRtGZGps7cP0Xl76Y7SXvEcJr+gOwGubDp4iponacr7lgBTrZ9nBJODxSZf8K2/Ldk24GT9Rdv
hVbR1uUUVrqroUNGs87gMUsMfUazn1aYiz1ys2dFT/mDu/LktKT/anaLRMRMYoJD74UAWLzwWDTk
uEa2j/C0R4UurEE85arWbI7QWuXrOAd6hBTuf534UrusLjeXJWkdPd3R4qvL4N0Z81ndWLm8Gvxq
wf7T7lak5aHu9CSo1ZAqx9+l2vf8cbLpDv8kg5eT593sMGlHZg4OCIe2HltZkHlGyzUO4uPGa8ib
xmdFPOiaSItA3nb/QZAbiGFKzYZYc32rNGs7J4Bl7hEC3AH8cj8LR50l5+3QmWDvfkNLNKmFqBdq
07C7h9FBPv6uf/b/ZpHX/jry901KeSGTSRfi0f/wU+3yE09vUiOt2y0MQ1A77Aqfe1vR4OYvXOl7
g0mXccmQ0brwChlT8WmNlNA0DRpodOJt9wZmDi5n0dYvbWGzAi5q3QQayeHxxqkmueDxxSqqFYcA
L4rAI/W9O+lXNAyrgNt3Tott+v7pAZzNeQDevYyJ4iH/l3rOLA/cjy+1BLVWAWY3USiB288z8qrf
BEGQSlqjy2ofQqCGqs1m306NA+9+y4rKLUn8W0MiV+WRMt1hIS2Q+q8k/guy0QVgXxYnQ1wM9XHh
oRQbFZfkMf67JE999sTqFOvPQ51c4VIAhcRETQ6abCLg/I91l1BJL2wHWT+a+Nc/HaJuaZ6GHZOs
OtTb6LbB9Ff/JBQsoIzo5KvfQ9YF5nP5tOPAgvUkWPV7B0mMulYcE6J3hJzFepEVT6vV8R3B8+Ee
Ig0Ln76Id+z6DAn6biCQzELYbPNvtzaueB+K9a0Qp0awRmQw0t8IGoiT0xh2fWUwm4y9MW5IEnfx
kCVOilRAfL1EwPrGP7EC2j1wTTW8vXEtvleDHcYIVkocZHZgN0nPDq572iMFc7n2KjAYX/8vxfwL
tsFYrcqKkLZzezvz4oLKwXZB5/+QQviEwzWc62mGwem/FqNcmDZ15SjTrB/3+FoDUHoKKtDu7adY
6iL4ga7MYL6LrZWwcF2m0bxbJHdNfhvXlWwA2A4exqhQiJg9viisHAqwGy5ltrO6mA4nQrmZqjfp
ZFL5KiGacf/khCxB7yNns5ZeKDu2JXK0y8+oJtSDI7m3hc/lKa1MYgvyBYBwtlJ7KcRrRP45m3x1
x4wvfHeuk6fECE7JGO7nAUQ0k7N0IauVPmI/xDFMuIE8DtNU/dk3fAkA7PxlBcjrFeqeeeOAhfG+
nyvkaUZ+ELZnUjpRTceiXIBalhsO84j+kSFjwoUiM3ca3ra3QAf3kWcTXoZDpQ6Fm7THothv1AYq
UiqKeVAKzhBzLqZKvLJG6iW0kNI9he7y/qYfyMs44PPmdLIb1y4wWL0RdkS4DqdHjp9f4DI45/wp
5ineS89UzPS17fi/C/j5tu6KS6EAiRc3KK5yJLEa2dqMvsR7rXEUscxGH+sq7xPkXCso4x1gcupv
koGaizmeHpl2eLAY+3z+c0XVAP3CxA4EJBioJ0dFj6YzDc+KI8S7F3NARMxSZa8ovqSwY1C3Mccm
gbbjnTvGaUS5EAWuH9dFmvJyanlMKlx3Ln/yFlvS6K3Ho7WMOjq99sEoLh7YQKdyDdEdzHoFkw+F
1ixtCE+BfR8TNPSZ6AwgLKtyUK7h+7zNYcUNXViinr68u/QZkrXm9wms7ld2qfBo/TCRv3x1VzOf
D6W2t/tg5K1uwxhhw/+x4BbpQ4Pfw0ot0Mim+gmOmbELH8fQipuK38kwUDGw2dkfdVJ5ljYCGdgf
0TgJ1PC9A92CqqrAOY4YsHyb4mGhv746CGGgdhlrlQS9FhhZ/fi2KsYBfneh/Jg3B++esAVS2d/c
4THMxaLl+5qBrEGAZM5snOkYRxMVvmfVr94qJ8NxuuRvpwAycaIIdsu2O/M+U6nBog28zZ2m53Pa
AX2yI4RpHAIAONEPPwHLJNjYWtzcp533iTAQbtGfvLbK/B1a3PZYYPsH/8r5yk42xOJgpIWAx1jn
wyUOU/hnyOizPTCP4xtadEF6bqKbY6CKVU6RYQ10JO/t/geRqdn5NvLC3a/puGuf2NvFii3118X4
pAl31hutn7IoLKpUI0pNSV+SzMKvd55lWonOdkH+1M8CBRYkT2dtGdJlkBv51Q73gCL2dI5e8AMd
/P31FBod6uI4df1s4fB+ly2WAK9+ir+lD+E9HcP5yz7xAkHom6nDedhauehhaRYZdTKGzvokVFEh
uPY5PkQyfC+BhTFUWs5J4CJTodCBiypwNFL9hvkk5JTjhrbxWrwsGxymnOMZp6HqxRlm1GUNEAoL
27Bt0+hMnWELTv3G7a1ZqS5zs9hmY2aluCk6mBhDWyYXbTKBA+njJI5Zb7EsTF4Ov21douTTUHQf
lRzmM4VOk07tFnULXf1q6Yc/R/uqxvNXGR4dcsyNoa8T/fhUmW9tCAH/F02GNKlhS/mACZkEGfGB
wAvv820PpjDVK+oMXUZQpnnxrM9Y0X3/Cdf3ixvppHzYLs/mMyEYeuH7w6fCIHIQxswN761i+3oz
t+uW7Q8PK/mQsyW2Afk2bHln0Fvi1kB8qKcB3qQh0A4Yguu+bsYuwQswwbbDxSTsdkSYUqcDfE4V
vZLSbU3nZQn+LOG0Miw0b6SMyfyEtV/kmdYomdCc4SMTqktB+RCCjLAUtWjtLFrQry1Qt8KJLPL4
Jqzd0Vz/C+gwi4urvkh5bxk64yMiBF9i9FZw+Z77qMubDwiiuIY6/HKuNr3MAre+y5LZP7WZPCNN
hsHq4C6s7nynVO2qfIZ7zuqTffmMJ/WvBvuQBPZoojy1VSURW9hVviiR9nLA1XLr2rCj6+fP9G/F
0JMhHsTLebDztR/V3zE+/aqRADJnGD64VC1zJvp54ma39mEOljs/8bnaneK5OwkIs6qsGRjKzjvS
MvaY6pDIZJM/rg5f7alzDJETtVQqeLpdIimM710lhIuSIlc6M9rGcp4wa8jbZWQtJn75whLRZ/TL
lzxLm1A+mjEKtbwni9K0RqjeLMj+d5PKhDeCTGrZdoxjRwagjBl8VPl/P4A+ey0NbUSNQE/KL2hj
Pj1I3aFpcpNQZvCfgx1pe4x2rJDXGM8hd5umWqLUe62ePAqPmLY8zNAH1V5mxPj3x9QTdT+MJxBK
QI6B37aSkjEqRfduRw3RHmghjntNPQr+nKqO+ckCLRW1++jGwjyqYPVWfpNiFuOpIEEafUfabaZP
VCi2ii6dQXj2v7xvhsTvJEK+wsxA1vIrHz25PHD576C9frhdsw0VX+844rrZ/uF3GE7iO1uL89Ty
3evKDeGEp5jtJV8mDZyZ/eyLjm4wrSB0mzpXMdrufhGZol/cQA356WO5gGVrEmWrHMav2Nr7kPmN
bDYW5BO1cvyW5khj+pxM+a/fP7IhHAwUJuIj2KyGhfaRzOoexjCURhQlMKR1xcS76y+LvRV6mByL
TalzUoAAPjAUPRt/52EWPBYe9Yx1NBPEvfdUukj3aMx+LsDVfoO94NrpaVPnXFFZ1WgdH190Bc6T
nTA7hnszS17ZiTcWF9/WwJDSddMG1jsihPo1vvbGiWydT8evs9dJdIQ/RhgOLf8JUg/WxHwG04ja
VdYIPsS42xu1QUGryoZP3ZQs7gPk6Yx8vTm00Vqyq0j3ridtcqExUVx0cgKIP0VkIgw6IyYGsftN
7WlSpXaWMKbDg0471cc7Fc4J6PvbITkF9jxvDDhYfQ9d61gUWeHp6QmhPdRq/cRgc4fEne+1veKk
zYpQ6zdKwIO7d35X2buAZ0sxDLYeCl/E3sF3wnaIwhweDVN0LbbnbLpMaVbDao8vyRmZDpB6bpRh
xC6SMIOFqxoZ61/O68a97OJTByPeE9Ea5dZ1jhou2O0//ZKYpsZtslxJahw+RNgjmQ/1A3hSKbuE
UUElbib6EJTEzkpX3XV1umTWv7ZvSs7atWB7GmmFFqQFkpl4zOWYFRrwKN5SmL5ZJmpE8P2bRgdP
CoB5XWFZbxywwxDzyydsyG0snvinss4Jkcg4cO3r/EzPrXkpJpU9KZPWMY2aiJeTbwvLUgl54Evx
5aa3SpcoO7BDrUXcA7afiFsDj5c72trHuUf3T6mYMhzkyqGDgVEW2d0N2UlHhGm7NQHucoFW+GfK
TU6e75f9beAncqiCMS6mbovB/+4bDwNvsKMYBsBiMwj4STSj5xERIuTCNrEaDLjzmH+GVZ3vqqJ0
AA1pdkIQKdjHbVa8FFsc/gcevAVBwVT6fNPNsJnIMSO50jgo2LhgtyrmY3rvahdBDA6v0pADu/Bt
k7XfTkfuc1pL4kjMBTjAQLfme6JeWF1mEG4czPXBJvtcXZZe8nLggzC1lN+BXfEaOise/nnGafvF
A8cJBX684/GVY0Dsqvgk+DfYmyZa/qgX/7M9eWS0o8GWoPTVG/6tPqGHbRXcR4xYqMavnMUbNI3p
jeeGkh2YwRri2Ng7SHhG4qr11MlZ+CgHqAyL8+FgehOsj/n8YfLDoHPXxJ7ETH1bfvfDc0hprgtX
LyHfoCSx8ukqXJnBM4DugRgoto9VitgNhqhtAWmgxNJSfsWEb3VyeXk+gfFH+gq7PTGmidK8RRyT
HP+GsmVwwAfPRmqK/PhDwbrC3Uc/THoAo+4t0bE/Xzkp8uwkvbs4xqlUXA+JW+AL/DWLuUPNnRAP
++uKt+y+xGc910XPPqTZlL5/OA4WEojoeaPCgMlm1efPiigxkS/Br1ugY6MY4IKcq139/77qrFWP
fLDQ2K6MztR4tOtruaa3lwHYaoBsn+tPoFOMBjyeRPF1fMh0Jdkx299o8g3dHiq1/RX7Q1qImlPO
9fxx6IdemMRJkzcKYjU3eWxO9c3swpG/pkXdqD63DTcVO80Ei5OW14mCroCwqFiRM9iVSG3sUwrn
6IN5fnc0e+VYdOrn0r15Cqsdy2wNk5KivV1Zo6dw3XZaLb+9jSENzGQwV+PFw2XPyRmrkSx2QJaD
sz5iHf25YBHMGcR7nvMfKI4FGDxZLhB+13ZdcpZe6Eq4sE/I01l0yczxPSxO6epOAVt9nd1D/QNf
yLzplz+DJScs05i52farFTy2LsFpqqfXkcINsE/TGwQspS9eQbqqND6At1bk4Iuc3q4bUHE9iyxW
5aAqYTLPzQghRaDgmMmM6jqNGO8e5HEfWslmrq2aZu15uq9VaT+K8FiJWsj1kcaGc88uYN7fSXmZ
uTrn6mbBM+VzP/Le502yZuQ4r6MYjlP1a4fmflCqkarBVJ9tHLx99IU2sut7zG9pj+LxeFEdoL1z
e7Xg5x4Klg2vYrL30l5ghF9mpYWj95z9QQFDGPhh9DqWYY846mi94h1V4yYMeOvwu32qq+PgRkD0
DQZ1WTLHxN2tdt2Zsg66hrNjVfu/ekNxhgpkRcuI1gUkDxqkVjYRLG+6qcaIqe3nEw9g06jBWQsR
9nV5k6scSldNyhr15DpBxSb3UY2wVIXHPCSbCCJfOkwczZnxKClgSZQuvx6SusWkHIG2ueliXxFm
c73rGlyp1bjCCEj9izOeRj0gu/nh8IVayhJVfbTcS9IeEZSWSSY7vI/kFKaObfUAm1pOOX8rHAtt
yKMbayrwPkFbiEyXAZESJn82ICUJL0yNM9zwdb79uyPmPK5IG8TDbnXovmmvzv6FWybn+LPKtbdh
YT7+khkLYKASf9Fx0g8A8kmtQVptjp0K2bWDMHeKzR92eg/SUGw+g+qQbJq3yDIBqTVjWMc6raT5
qan4hBgwjzqTyYNi1vW6Y6EQLH5s4i9m04YYbpMHjOYruHIdDd9QbiHnqfNCaTAIn0w3BMokUFfi
vJ7W7c4ly1jtvOUj/VcafNw61yyxfTJ3YMz1q/P2ElwFYmbTHErxpbeGASHgfrFKG1baVoEgHma+
grVDRHXER03Co6ubqxIa3rausQkacs1M7RNGKzvcxw44uHAjKMuZmixGxProzk2oN3ZbQTGLDc6J
EIk1p1juwdReoQzxpoZnRHfDPniMQq9bkTa7ApdbgdSFHdA65cwD1U4GOOVLOnKg7pGt4tzSGeoF
agpZeDekfZDpUIiZ3bMkuiP6m+D+Uugqq0HEtp0pmrJ/YopAbf11pI8YElttXbIiXmVRhsaE66bP
G3xy4kBTwpO6OrEBba1zNk3p5ovHPuTC1qYCcnXWUtapI9iVOT8OOnKY1cznDIYf/d6l7pqYJRl5
8zI2HzxbDs4qFloW6Aw2bPdpIUKUYSLtJygf7lEZJ8t3lu6HVge4SvotWPCSkoSc7nhLucpZXg0g
nq4ZqSvdmgXd6km2sLj5mO+kTF1AbEOCPBIGX5bMvm1eEI3kMm+ampHaM0svCcnwUWcFcmCoA/Pp
2IY0tRkRfGdmaazCMtNlIofAIPy7EMy3IeQOUwx1BbGo8eX3wKEdMUxo2CdneHqjC/QfkbHKnWZ9
QROkOgz/m1jKiAMqsMrP9pSUWfH9bu/8GezFw7R8sJISrqFJNig4zDwE/QN69W6xC5T+i3DVxn82
YxjY2l4SjoItB0O3nIhNCD88oNQ0neGWKC9ckwJ35ZLqV28Wwdx8GXDq8IA7cTZHcbb1Vk5n4aGN
GZLlROAyYiFx5z+JMy1fhbF8eYeGyXDu7EthxHpo3atAPn0XqbksFb5elLcxdMcxNoVLAm1FmUya
PW8U0bHDH9yM215g4AlsTuudgeG3SlGz3r7X/zw7y72Pfs0I5zz/kgQQUY8TAGLAZmC0jtxMoqKd
eaPLgdsaISf9VzlroWJUXPqYbxSONYAsw3nRk9n8cWxbZgjlQboSMz4BF7xkbVFqmOJ8XvwS/ryB
EmfFhXDG/e1K3GvuFvdhvNMMl0mzZf8aFxnhXkhl3I9aDpERSD7ZwZsBUmEbjlWsEc/LGtwd/JpK
iN0FUafO1hyf/fINEGZs7wIyzXoZ4hSVhxreDQhwGvlzkvywPS02j//WCPCnn23ejkHrJad9i4cD
OAMIYhwysm6u6if9t3eewFSL5EhFbBGMglgkJekay+l9Lg1eLKViBmjYJDlWmYYgTinPJZbJ/QZx
6O3LOQji9s74es6A/5GuiT1weMUmirc2eubxVCQqR0H0ZTpKKKcqLdUw5P+JjAQJHhMLTvY2dfWj
cJx/nw1JKxq8nEWy5szq0KugCzuaVUtMjcrDybYY6wm0tDgaDGu9m4NPoaf/ab8SoG9iHJBoIMqJ
Ynhb8X4LZ0dLOJMcjRQC3Hdt1fNY2M/DCjM5FRttjldrt2zCofA8/snfYQ2r2q5iEpmIrTqssqTV
sitVQmchU3Mpm0faCgjK6Idko+YdkyWGKOMJ1Zwk8GMTN4mMitbXqPCydExeFC32Udjv0nUsHri7
G7vqjmmuSX0jggGgmpJFloni9eMsO2Jfr4pBoq1Dwd2bwzqy68nxc9crBquhXrdDdYR9BxxuriTE
dHJN8p6GltCzJTZtpqgEhp5WUDJ4nEtpvhp4kU4hOQe5jfP/gPT92R0/Kmbb3HaMF/qo1SEn8YUM
Jeh+o/LtnkTM+oIwAQGd2io64oNzoncpfi1LDv4F1M62chle++6ePWvoB+PgT4LW58olh+gOdO15
2qVwmvRlsX7jxt3tP5fAPqF1YuOJgfCnH4XDazkbesKgxf0qeY7TCV0reUE3dGCQoouwBN9kyZhS
pB1ps7JpKIN/0OcJosqClxdoPqScy0zzxQZK0TtMREhYfZ96n8E9pDA9ZK8OLDXKY/SeexWryOF3
/lHyrHkXJ0oMlRbb0roeLzewcpiXjTkaKnOykcQB040SVK8bNsoi8J3dD8CIkpUrCNuI5fR7XpOk
b7IqC4Sd5etmi/RDED1Hfe8LvX9ATv9ldfFTEYmat6DnL2mM4bT7LjetPmktFydpiXSuTwTKt2GJ
PJopLoy3uOTdYqjMLSB9D1uQw3XumFqjZEPfHKGQREsHiDglguvAQLFYDXfQasuSedSj3D7J5FZB
prFKk5vz4bNl1LgkBMHaThmipJHe/47HlGHdwBLZ3s4MTEmwz7+rx/d9FYvu/U/F5YhEAcCdnwK8
FNnla6gFnG5I8SSpEI8TE/K9Mdl00u12x1vFe8qBrdhhsoS4WYtkqYB8exnRprhUPBMJq/3bWQwH
BStetR84qBOBKoOaIrYaOuaDuOQXw0J/VwKxUUMc9gd84Hoxkos7mOyXCjsvRiJBGOiF8jbArYJ7
lF9hd/IArQep/aM9M4kIhcDbzT284HBsa9vIc0ji1H/eG8wt9oTZr9XApHEupwIl9kJqvl5zItpE
ja1arUu/WMKiflVnRZCrMpQwvW9Qcf41omfLk/XTnBZeIEM2Vst4AOKhUupj8qtPmqJCQZyioApH
gj3o6obIqmXPjO1HB6cu40DeL9ihHsniOW44bG8cyDZBHvz4AQ53ZDuFbC9buBBSFlV1l4sI6mow
gsVWr70lFH4KvFxAbTBAHp971Ku7XkMW+NmTbJhzEBoNIv9QJCv3L8Y+UD6SWovzJkGEYxVfaI2E
pwguFBQV3GeBEUqZbJjOUzDNUKtv/FxI9rZGmK/WoNWW7MIjQis8p+Z88EH18dNUgwLL8NSNCxRE
gXSViBuHIv1BB8DyClWkzAhdEVi6BEiTYwOST27b2tGAHmwcCRH8OZqYu2uveCPF5fdPUgAaviQM
2IEiQiYf8qv2yjdsgSk8J4Zu3BuuVg4eevjIiF8JjsBcJkk0Xh93qyOpTp2fHX79mLb/l+v224GG
GgOP2x4EZ0uNrD6r6Ok20/b12ket03CNILg5wy4x/i0PMKDQA+XERSpyjuGWv7Wr0hVZSunk3BXe
Qql1J/rQPtg+6MjqkkP4sCK2YjvGj+7hUrGjJDuzfAkuO1mQzdsgayvL5NTBxmWDdTtZSVs2z98i
yZK5kICqQGeVbgnIEDcF6xCxE9MAdosmkPsQ1rYij0x1amG4tCgslMcX4i6n5cvobRSOzUvvJjCA
sfDW4q5wGgHaHUBoshF+s9Z4G21g8+rFsav6goazEyBTDKfjvN7Vg0Jd4wfCyEiUuMVhqGLLn31r
+eFQwQVmLxmDJGwMcbwA2yN/fjkrLPtMIcZbJFvHare+bM4LQwYxJ3DgztyafwgMiD0MM4QKE9TG
fEtSOTNfm8Bep7ogOaZi04pHFWiavqoR5OuqFjFDEYqds+TQWrdigbvs3vmzgHyfOpu3lc/+NGrZ
z5DYpm350Z6fBagWjW1Df4AzTafYO1q/+nXd3rrw63jV3DaVkASAU5opCVAIgt7HtOzazHQSZnFm
JVK1lU7+GjMnggpNvhyLFjfFZMeRTfwGYoUyMLwVkrwyrGY0kC8YySuZE1qHCx5Y7zGG9rv4lszp
cVdBm4unuS15jDUieJ7UagnUj1/eDQI8kXwsGJ5syAQRT/HKBwSMNsLozV8oD2HOiYjzjNHt5+yH
smc26F88sK7tvSqAN+pB3GtaEO92PiviCDbst9VpEl4R2P5IybAbiDDIqxeBcsNY3RXuy/vgip5m
nQFAtkrc5fHJMNZpVlHgPXkslWs4EKxq1DRg/M0qUMOrbRllAFAyfG+2E01fCke9WN5Ye4j7FQW/
T+co6cIMFRCcUYLWPCzmA371nM6LwsmLTagB6AObfRgrFlEwmmJDqe5dKan++QMrlaxLDBU1TXkd
G7PEsmeqD2qOPbquwUNm1BMIv60UvKqK+U9xovBjiuyBLGs+cb5O6cm/Als9nNzjUCDhyIM5ACAf
TardgJY8IE0D24EEeacln0tgW4eMg6PI6REVOzJ8lHFOnqPVqdFsBvVBc8fdyOWsEQ9TdzYuMnbk
UtAQMRGGItfVbgcp4LkvZtgMWgV6iaWhvTiAEnaTS/JKqrsGTCyGR3oKQtYSg0YeahSRo42kc+dY
VnrqeNP5oOpswyebCv68/cXf7tOjljfncBANb5cMhQDMA51R8U3NxuZI1eziln2Ti47DThGh+MJL
fWeqWCXltsWRF9FLgUfXjrBQFImkL9oSTMgayn7fNpT3CzCNmTeHCDddJeaXBEoej5vD+BRSc4wU
q7OHXcY+Qt56ijIT10iHeE+6WxrTI6riO1fVKjQOrUkc9YRHN0Ge55bPfyn5fZBgd4r8+ELU1F+R
TSsBeo7XnZirVo69i8E9gFo0zTNrPIvRzs1SoX+MHlMdHSbHqv1wuzSe0G1xcvHfb5cNfgv/yodB
eP+5EsIE9rE9AExJvrJUyelH+fxc0T3p2aIsjbYwMEjZAxCKYUVrjQgRZUOtP3Y8k1i4uperlIQj
g0TUJYZW3rCeTM89bLMzOgeP85NRXyNypjxtUrr/fal3tLxy771aAm97leQ9OgoyUhxO2MJKGuwo
gFu10GQvXpjcV2M6VVmX5idrp2RLgOy4LwaGtfEJXLu4+ofbwQ1rv1eRIbCslQLMtg+QG6r9f+Ya
7ZAW6gFp3gJ4wq9hi2Nk35k7St/IIPpP34KT5dNVt9DuS4DZrOszTAQxTPvnvKeXopsXPcDVSXAv
Uic4X4dVrZwVrRq1mZtwYNeDew0Y3Ypx6lzf7NWlUtQYusyukrmDMZwV4ut63Gs+UHL6HbcpPjwm
f+GCbjBpT5g373+Q3Jj4iyNXatATMnvbB1pBMxXE/4m2LhV7dOzI4OUAkD6hlh7tbfo9l8NI6EU9
5KnxUsIBmhLeTk8dChdhqXXO204av+AAf6k13ZsI7Yvh4g7L0S6DWaEWngKXQAO4osjKsC3SVQgi
pS9I5nv9UL3xSwF9bN1Wy9dzh8OpNIVV3dICUN2fuDqNfk+GRB3ZeZwylt2tuABPcvabrTObkPD0
nl/I6vJNtTc6GNMLDjUp1GinAQ9gYPLB1CwfWOdA8BUANtpj1OIa4cPmvmycHHFCb57OnWaZA1UK
Vtun/11//btU5D+uxuLMYJFeV3CJ2M4eXFtfpiybykYlzOm0SqRGYpqf3JoNBqeEavB990LpnySH
+iKwUFAbcmD0NgnNLxiizkxsdR502+29zxeafXyJgThM39CrpisbdomFSmwfJXQavKBirr7QQbO5
lGGJWgHMvyR7Eietu2lvsCo3dgb41wWZtgGEo6Np6++dCjCuGL1dUliIIRsB0zKTU24EMVr3CGPh
HH+qDYnOEtrXuPnEAlrUxekdSUPVrLFCugaCvZGvCPb+zHXDVZ4VgbYfhf7GHlgLOl6wt15ax0Wr
L3MafcFx2iQ/wBZE76JCS1rmYKNJogZ3JcJcnAgcPuAj/pWZNciIzlORCmtq6QIXKMcmI/aFpJ6w
eu/ilaD8RWtBtW2diLvvhslKo/P/zwX6hii5WCiPnxl7a7Qatwup+N88cuaa6GSm53Sq63vyiwi4
lDoFP7+R7vzS5HLWk5oANHutg6hJ0C/AKceZeZJF+ZRJBzCu4Z6ZG+Wwo1w3/Lf0Ea0UYhfIW6Ke
vMUjYlLC96zJL7lO0uMM6IMo6XK8kDxr1x4kp1HNz1xKXYMR6sVYEjwBmR2MQtThuoy+/RMFXEFW
eBr509OuBLxmrDOhDFKbc+cxLyQlJblA6DGy8NKTuYQ0mzSqj18WDcvTaH1qFQzMnoG6O7qJTu/M
h7r4vJYjzVyteEuQiomsoGK0+LShmMcnUe+aNHvqUjIQLMOGt7zEOO5RJ3sbdQ00gbBrm1ycDOHj
iIdYRXhEHpDMwxob7bHSdpLLHdcQl2jseQmZE7ZvttxfvombSkp55JN+AklZVyzoejvM+CSg2904
L5lC6M708/tEpDNivUlknxNe7+04qx89w+951tE2QGWtXZmbAeAkgR2gMggTqFJnaVTOC/qhNADj
TPKZIxxxcCs8LP0I6eTpxsV9flEYTGRpyXWGZbzLesjWIiVEMdhZryQRjFCVD334Ch1CLYj9xKKx
KiyBCFQStxPuO1Zae/DiezH93iACq+nip/7DSE4dtxnH2XgmGzqp4kxLB1j2r1FwVHCwbbaOFwPF
HBxNd/wzjYD2oMguhpRxs/g7T5sUNxnNRrYTZducy05Eq3+AWAzyRm3UGKrSbUG40zIBl6L+HNlE
MlsbVDvoxrLBk89kiWLvEVPYi/TpgzMFiszsfn+n6OzqvkV3X6mng1PleBeJ6z4MqlMEEZ0EhNFP
LCKLdZVZKQGopKDQo3BYfaxIGR84lGI5riECc0P9C1/q/FqfPfNWeTX3CgyRUZKsj1vGDomcS2S/
qCRjirwYOtqDc7cseTxTKpgueWmf/MRu805TvveG8rjwyTJryVGkwPTfdl5XCHZGFnQ889DFM5w3
CHq1girkDvrCZAaCH8gEzzLTSH+4jqJYP528x0xmeIwTNncuAqCGsLPNJZQcE5UKV4aDgDfbFnWj
zMHNRLQOCnHXI3fV1aNYy4YE5zERtWalp+sV5SJnFiQEHLxiGa5oGYWe6tQ3vciLM/fby+xl+raG
yJO9i+UKyfUOoBqmViyPJW6Cjd23hB6WSV+gC7FFMlKPFjUvX9WndnbgImvABePtBg/3PHVzYrbl
Bp9FfzDchRFJNG+/duXAj+bD2EfRyiIR3LXSFfeuU+HFhCvEr/ahermhC+26Ywwy2epDnp8ksnYF
y1ynwva8YMrthCdRJOcvY79wiEBfauF+0+/BIORuMJ/4j/u76qEHZUYakOFqt1rykAYFHGX0igeB
zBFvTpFuhvoJbo1P0EoftOec0w3Xg/g7LdISL8mX5TokDOetDPGe66L5CJ69NhD2D5/coDkil0UF
qgYwa8eFTXoNdJAOaseNPsbAMTPhUiMU8eexk2XRe2Ws+orqMkvdr/K0atwwOt/UpFT9e5ZbPiZR
PyThZh8xh2T6NiulENNVAmhII4yMml9KOwefq5LniaNdvQGC0GI76JTCQCVcPFGye4003u7Gg4Lu
zIWug9cpOnlsmkqCyqYjM0vq1nVSL3E0CVVaTxO1fwL+FdRTZfcdzpvXzVuGAgUCKu+T2vJ49ZK7
laBMqt9ZHjaP8iFGhs08atCL1GKDPW3NST88rIeDqol5fPiz1GJYFAEPtJCapRmhHIdG3y1zgl4Q
0d7pg8qt/P0Jye4M9hdkYksO/XIc89fNWCxHJKYkXA3LXgQuEyMtUXlPzbhg8s5SOqJom62abwCz
QNE/yDzEM2ZoMFSmBM07IYEkTWOtIrWNsInH0s6GMXwt8sqPJ6d1V5nPWDCsImMRBjOv+nfzuejF
zMgCrQWPltTrDLCvqDhsRJT+uPN1Gri9HPK94tqFI6sv3g8lgBR2Lo0aPzp8oSGd62GIti+JeXZf
U/agRVmGp7uyeiCb6VyilkW4UHG6PAfF7gKIhg6XiHZedeaHJ+gEaLBYB/yFufXKdAwci2VZk0Wc
O/8ABufC56P0suu5NKl34BXu/Lno3GhFJIn5x9uqJVYFcsO8EPCE3DZ/mks81HauIgPgLnxV6jZ0
dRqPdeEXqcXrjOXYAtgAcQS7aYP1dtypw3rJXjLsorhrj7SUinLbbZD5jqU7FVDsWqfuuRxAZPkx
5KHg2m3M8BTleQFFRXsXpeVqu40zs8EjnoewJsrEpFKYrNQnjX5EdG+rGbK24gVQhNQ6Yo5fmon/
8pxb4LkMVAOBU54FftweVDcxLnn7LCceE05ICgP5W0wusTFCMbgPuh7bI2x/uANe5h56tpcnC61p
eYbMQN9ioZrztJ4oNpYhccIJ0qDF8dSLIYq7gwbUjpBL7jVy5gQPw0kMr/1mxngYP0iK+1nDzwHI
n6kKDBVD0cFTlIYpZoJ/AkeJWHpFG5YZpMPnfZa0/C+2SzYFrtzqsTlEpuz8d0//qVallNljAE5p
7fh67zAiDrWYp3FrnZkx06kEA38jTcPxoMY0RX6l+D3dLJb1MyKdxkD2Q0eFgWoApW9gLm+U4FQY
O2BbGluiqT4OZNXUGYLz0S0CyRhF6l1AZoU+AFYITp3aXkKHuIxwqBkGJNiL/V194TWpLpvkCZCr
+BJZeROl4+IH2ub7ECRSJLkzS5/g5gHHHPue2mGvt8xYWdX2m2UKBKBcuIZ4jUvyIMMr9TuXAJ4r
iT3M7xc82SBoPdQLwj5eGpR7mRinL+kSevTJVGvbW9eN5ZPllquLYRFeMwMHGPpheGOmMij9Ep6V
0iSa9zZwzlKIByhD2ap58sTLtb/BuJQ/gfKI03RfyXiMNVu7fsJWqK27MzsaVHzlXtAnFuHF6y3B
vY9Otr4cIvGD0J/kH/Kuim8l3ujfDpUWE6tAw3+IoHQCO0wurCN9TSxVu1Ch3xnb/oM5BbcSkjZ1
mXk8uZFjHXePq7lWDg1SQRznMFXFoG+O4/d3Ko8LUn2Y5Nb/wR6qPaV0RPOlR68jPlI916tPAH7l
/UcvCxXUOD786+r7xlABVv7mjGSMf+HizHIkLuU0HvrYBpcK+HLsFdmKrB3oVob8joQ71a+1tCIL
PStarW+altw9DJ36OWRi2wDJShlyPgnZ4yVRntKSpX+ujdPgKB2K9fXP1SsLFQSsZtvRdbcHYEPj
ld73k+DyIVKRO0bFIAPp66rxRvSU8Z1unV+JTF0aCvrZ7zssqx3eKQNq3Q6VkYzDRd42cYBBd/08
3aEGlQHji9XEbVC67mH34F3PsxhPZ5iNVfT3j1FneMjiJzovTKUxMKemUCuo6kp7XXbyqCEs9G2g
4HnB8nqqlrf7N9ujDwY0qotIbLKPt8aiPloPSPhlC1j9fob9LPvEAS0Ca9joCxim7KfC81Ub6nW7
dGzFHa2tWTPXIOM3F2TrZO6cIcw14hzv2nVJ9Mbtzfoo/hw3Jyvb1RzA2SRKXtzoBbWXhwI75evU
sBANSjw8VXDaVLxrUG8pYUcOkpcebt6T5qwOy+3p9w4cb1if7XuTJo+dvWyVwZUenO9MxsB14Thg
971VCmDBhN+CUbE4cuPej7ap5/6MMhsdSbeUvV3DZI9LUOHVQA25oXkaW8lieT2o5OzNmMNYAoY+
JZ/fliyByZmaq1Yr4diyYw8DvnsvFM7Xib08zuFbOCW2kayVcf/3iIOjftI5PfXgpUhtwuzHO8lO
b/5HrN4VJ5jaO7W9gYNCJ48OHOwZhwwR1Uap+WcOCOyBHE4lc7t4ZdyNbW5jkv55M4UXsp7bxI3Z
0QfJ9CCW57P99UR03JMVo2I6NmwVIf6Q14yZrR2AsjBju8rkmzwDUg71g/aBg7psLlU5OKhwAvyt
rXgJkQxkyVVAjv1emWCH/fM54NIpKNdMgFtDhrTs36FaBibNp7ph1tuoEcZBeaxgKlh+0PHh3u0z
e9sTdCeqBV8x5k4mKYKmnIeB2F89nxnqKWQs6JbBnaQ6pNq7Ui5ZRNcziYLdSTq95MoXct15C6yl
6j3EaFymEWLBM/PxTckjUoxdKbR2PpVoPN0EM1D7asBkk9XE/LAt5sKY3SHCDKUoq18f4XkzAz1P
ngtsQiNzggIw/+tZgwr83zBf9hCoev3TKpZN7w4NsLbfSeqpWWj0EpaHeag63fDdXBRsgPm/tDZW
7AgTr1uBXaVGCPMgQCP8VQBG19uyHMhXtoSule3WO9oJLIA1I1lSHn6tV672UJaZRAZjnXty6u+J
xqLvoAhiIHM+eD4Znh4l/TcfHFyst7IBDPqQqRS66X4ePRDzXpELnqbyIGE7+CCu74KUpUUvpBUC
ZlwhPypQI2my7sKWk7O2m/i6gZTXEXxwJoijo2SnGkX9fF2+JBbRGv9pvigMGf6n713LOvTQ81KL
hYD/H/Ex/ZTL95KD39Omqh+b4NYdSH1mTNZYQX4S2yJMe4wnb1qOqQ8+A12UaJncNmY0bsZFYYz9
AkDeyKLgYMdamMBzn3wy4PwScTft8/B0/1UUqBY7ibgO5mgXh0jRm6shdUrGwkilnNyKC3pt5SEX
hXwQ0Lna8wWogsdGkzAWefBJ5LBvHWV61cwXJS9gW88qUmLMbYwIrj1nRMVVtUOl6y9npUqIFLf+
TqdxLMCBtFhPKqynRLbadQaeN/UXlWfh/Yxl0s+xIjJyAnbifP/f2wbSqwaLMYyDXp/clOyraneI
qBapy5YZ1KDbGjHi29bdBmJqY1ttm+7oA22VbySLGVCqG7Z0GCOOskhIApRede5ezxnFe0Fjt/1r
GXD+AEbtWuxocHup5WuEO48w9y6CT/yGSP9Spd97DvNoWxafd8zBEUwRLkdo9wBipRlt1R68leI4
ogqfz0kMysIf3/3oD8qDFmxKiB6av06jMSI1C9eyUuoWs0r8/Z3m83SYnxIqXJCRDNcKIn246yDi
zlN4CKDE3XiKtydOwTH74dPjPBD73a+W93oKKg8GxMfpIhF3FGTFqKQvEx1B7CrxVkW3CfrSmNxi
XLaZO1/81zoaQv21C5qgGcU06WQNQmUD276JzAgbGxAI1X1Biz4iBV9HhrlK2boVn4j3VuEOb3BD
OFgJn2zUXVjYR1yhw6rZ6uXLeVYAzKGoADlqryrCulchl8Lr3TcO08qRrS0QFS9dLx//CVovI786
QKySBuwHfwh0lsQx/WWFIy8ht738ffIekxObVzFki8Qo4aprv414EsKuFsUBehjuWAfFD9ZYj9Vc
/eB4BhbQuBQSkaMvpLF159OXuV2+bbA+37P1JFi1Yk6/0Hj+0MNw/IFTokhPU6o4NDYWRNMjUNRr
uAi2WT60exX01YXLdvEfmvNw6cJcchNrUQCsRDMCO9G1wrSCFr+dQi1HflLHn7BqKL/aMnlPf7DS
Akj8F9o2ecGrbU4M4Z9fdVsxM/5rP28jUnpMq1hXdvVgsn+tkvFWRW7O7RrZELZyrecVCKjjh46a
7jv7l7E42BuPjkWzXnCnI4howSLTPkraqXTbB4MdH8D756CAKo38+bcXkdWBtJ7p+sA7EKstAU26
GdvUkE/iLY9yeSgZe8u5xERwqQ8uwZWIpj3Xkp4g/ExC674jr9oPLmXGzCDDMi14CcUFSEfuaslB
T8PQA/oTFAbdpMyBdy2+7j7sAhQGS/KWR1WbLqC7drNDmSQMWgeo2/jXj6YzKStJ/NURHWbjrGtR
1dFRRJDOyacVmZOZgO01FL0a2Vq3LlT4L4oaemVkATrDBG7RgPnZrbkQgtrcZt/A6ZLlzAHIer5f
BDDJSO/CzOczAYFxXgs4w42teTqOCnw+XqaiLBJvgYkYIgG4ZqB3gTAcaW4xWvWKEfTIEOkpEJvx
K85MIJ/PM6Ls5bIuGneiwQUG2NmIA7Fs6je6naqtYJtr/50+gPk4RX2+k2S46fsAsqOJ519TBSgQ
GBxJ62rAzFgo7qucfKsbQmlX+lOBnJtUMETjnk3+u+1hnPMTxjZGP2fpN70lQnwkf4k8S42zvUq/
XyV/X3paiVDx1UVXOkvYEteNYEf5rW9m5ydCn95wGaLXvKzQg6+vGz7WYJR5ZBCPmzCuZsECfj8/
cTVngjoMrWX8Zr6RM0hd2ws2wOFqtnrDPKMM0Wlu31F/+CYtf01jZderKVKteQ5JTkDE5IvVYZ7Y
+48EOfkwMvg/Yqs3hsD/DfAxApoG2F2k0HQdTvjj/x9pfx3ry4Scc5vGHvD70VMzwTqOJLV6kb2X
KdR1WwnNRboTLdGqbxfLzIc9HuqBCsDWchmHZGJreUtYtj8sl40v2sJUTTLGMY+H8fF9kpxTk5l8
3GtKUx2VNCekOZ4P6T+jDBhwAPG3VHp2rUwoulAhfw1BErL/smjySn/V7rKOWC/4ESnMdnZTHXnL
I6mBcY3dCvVqumzRLDt7Fd5fyOW04PO4ESaH+TLsf3fOx4J66BHwPV+fC+30QX7GC8Gdvt2wrjKg
7cOD5F4HHBvRclJrmy8zbUgVhvl8+6P+BDVkzVdudvpMLRqq0p5JmG3Zfm0/Br2t724Zj75zs3io
rctzdDkANDlbCh/Rk7JeVpDC1lgulOkzNrLfZwRMKp3Y50ZKsRm91hp3fX4HrfyI9UDUj4PvTlL4
fjtrbdXO4nej0bfX4ofYwK27nfMhbbL9I3S4IqePKahNc+xE9H36ARbSPjjA9ss8CnoET0LJ320O
DTqtZNIMrgfNNH1EIr2ft3z/jCYXBkmBuHCwVlZAqFilbiyOaQOEnTdCThOZ3KMmg3Pjc406SNaz
YIu0fSLnoS+jLbFtTHLyagICaJws8BChi+OMmapy0W7BlaNELgU0XcMzadZcQY57mZ8r2Z8JgCRm
+qt+/9veQU6B0VrTpw8qpUm1nKzhn4FHp3Rg2awMN1215DvbCg3QA1U3BTOhXwbpvu4doH2cXVnU
1jegWgviBD5N7qN/oiRZVPKohCq9x0bcQRkOKWFrsPhAuQ2BQ30eNX/3SAGnITbBJylPm9HlC/tJ
Mfkuj83Evtta5k3LZmkL66i478WAeZK0K3IxRW3wmrBPwmCTUc4b5qpZtI5ek4Dv+0B61JnOqFPS
a5jPKeOsaYNVZKsbuyX/uvk6w0SW6l8Rbe0+lJqwSgDf9Hav+sQ1/fcocXuHzeTEko1KPRMMkO8a
36lkQ8lkui9MJc67MeQybZlOoEsjgJH8oFoDunJoysRxbmTLWqtBfLXms8qkn4Ug4F68NmZC55QP
GKuQn4ucADCqb2IZ+IESFWwPRrELx9ryqAlCgYcaZj7ZhwlH0VekMRdhHzI2gvf1VeQ5Zm8KFQPh
AULSh1jUXpeAQQ0qn4gcV3Qai/DBWcBmzObqxU1+KH4hR0pYJNa4TIGdU7OT6Dl5ovwypqmaCZJp
1H96ICF4rGi4iexky4fvcwLACaiKtd1n/oekx8j216XuCNzNzrv7ZHiHBhJaHGGMbARJM88GwJfz
sSx1dhVSy5bzq3Nnz6W0dnNEZVCCUY907tFwnYH5AjMXFZ0hMofbQGa3HIJRrP/8RTSepDHhDDCl
m+xRN6+wPgwAO/BI0SK1BktyqL9wsHmGNz2TXwhp5j8zb4BP2oRoHR5cTUcI7BhXXMEKgTfnbXZb
zGV6dT6RL8Nnz9Hb2PEkesEeHEwH+hXQNX4YktBGFS8uzL+9N/cf8USETU78NLyWzuEbykFESOKl
KeRMWNnN7ONVElSCqc3V6R6cdRf63/MJpcsFsdGTaDOPW5sjC7gzoJqielO43Z7slr8kAradVHEo
KJhaO2M1i4rEe0/sUoFbWWOW4kxmfQG12pnuTs06maUJskFREEtx32ajqiqNLM54t7uvzZZrZRSN
ov62PQm+35Wn3RRLxBMCSRteY3BF9TPWKZs+WMQm6e5PmygiEHddggBBYfKrxKQwQz8oU14TtWTK
njUIgEWm+dniU1FHGfYQS7Ragl7lFjIrumZeseu4x3pq5gregjUgaWMtCzDSPLABVmOJmAYRENrY
NjSjQX9/cHXF0IQ6EcWqLomeZGnZ3A2FDtF/6roJzFjhA0sKGiHRVJBC1Sec4SIlwNi+p4PHBROp
S4dsm/2Nq9qRWMVC+0v6FRzS6XXRnoZdc+bDYFMNxr4acns1x3HRvUO10ourZcZRkYyaW4L2jlRE
vQJp2mmKQioS1nhmU/UeSAUxWjIyfbUR29Q17q1Kw6LlrK5e2jZyCe87UITvRY5LpbpaONuBOZOK
vtN5CTgtn3M52B2NV7xCjusMlnbFLcmkxlQlsM8ooYoNtCxA1S1gU2GkN8oCibZemHbkYDgg2lKE
FVAn+MwfzGVRCCSaA8IOfHxSQruMFrPG1ckMliSJv0XHmYgZg8dD1T0fj6Q0ISnoicJJwKVsOgna
gCoEvF/hioa6Cp3HZaDFNaqVFfKdeQdC8y3+WUBVROvJ1apaVrIGek8KoFiutFsxQy+HxHtLmtHm
xz66UtYZLBzzu6yrq7FgoDihTUeKhnf0MIoR8z6irYfJOEZExBOg8DnxNLOI6J/5R1R776ulrN7I
ww6kO2/FAuLpduZ4HQDWPznqG2miJm1w5fNJqtdlKFs/okUPArcb2olUw+gBtq89oY8CK7dsuoqa
/i3XH2HJHLmweAVTu4MFus65iRcWeZyNfQ0y0I6axC0Z8Uzb8ySoS65HZtQ08SUh25Sd7CWWGn2N
rpNhZt8pYgWBHFRx358VEQ0pywIuAYOsoPfH30zbClp/apm5pBh7HEcKa6S1NboHybs1A7eEsQvX
FdldbGp+P8Az5jwJR6+s5okbCLMCKiDH8v3Oyf2Tw/Ffg3Z6Needvs9CeEDdDE0PG/2e3G/7uQnG
cYemLSblEeomZDFI+ogwI4clFHoKQvNCJFWRFBfpzjFH3NAbHGB5dPgGQ+KY8DvizIednPxRoiKr
/j+ldrOgCrrZuSsh++qIw0RYFkzBqgMY7XQUwy0Wr7aFjyYwnKb6WjS0dEMVmJQDfKgL3G+4l52H
vYtUqbT2naefrk/K/sv3AqtLOiNJEmv/IZT2GCnc/NjsaWm72ab4s1onDqcT74mh61N4fVxHmCWp
JiI/1ybc/Tyt+GTyeyz+4LTpN1p7J5BfUX+pzdZoEeCyqo0yDUtMdUCzcqJeBb6VkhSQUk4txrsa
zQR3F8DL9mLGWmVrPoErYHWnTIHC7PQ75LFI/j553uwP5NlJS8JrIbVX6c4rlkbNWSloWeyNNuHC
kH2vF+xkE1p1SfnOeyX9PvPxi2e3Jl4y+KOv9bn5QoWxRMzRgPwnAZAJoqPUaalcxs/c0+uYuEfW
WCw7jdSj5vubxPMfDcyYLU4SZedJxRvXLNBw1td7r1dzWK4aJUHmZ6DS/cPiB7Yr8rugCDMH0eLK
Uy7hsn4IWGNMn7qr/x3PcgInjBiD3/9nRzWR+Lp0SQ3BL3LwgQeXKivs6/hRf8cUeNsX0KE+DP/5
xCfwMfFRAigvXwtQ5Z784k70riCyaBw7khyWmLYmTJl2OWHLrIbE7QgzEnYrqVoXwaLtkjwioAnj
78W3C2ytwtL7M8OKWbo3cuWGLIqLdsPDz0wFaUJTZzXjoKnJ5kL4vnXMmW77PfzuAWh5/ghV7wVc
tzRvqIJxx7uj7/thx0/7qdeToVZYt65FuzNm6ch5gFlntDmqPmUpIFdwCVg/gkiOZOMP1kuyif/9
knCvvn3Q5aqaj+6Lu2/g3Z7VsZNcMaSIcDY5Tytj6NDgJr8BR7qA/Rr5b5/APhXyhEg0gM1O5FZb
FGvAQ0/OhF7E7gTJgfgZwXGvs9tt2hEtmoaeCfOp8ycsNrn+HZFAvVOT0EGmKaR2duMJfI+T4Kwh
F/cZu8nU06fnzLuOX2fmpQZqt46fs6YJ+nRz3ydgJi73CX/mkXHE3Oi1fiNM5fS6enWQcXY+Pp77
fspgmVPtwP9XAwXbtB44biGFRARUjhJR6rtggwdHgOVzD45Zamxr55BOeZNocJB2xliy6lp+r8/5
WFQ593VugoybpEEizeEpNuNlPFEf9pVNut4pekMtcKux0Nfylok/j8UlOe4wz0t2XAY/ItXSYnoY
1mGmvV5E8WGftAWUWivxzfIMDfYBjc3iMOSgPRye8fW68uzyWx8ojaOzM6kG97XJbbmRFW2fVWaI
nPlByKdt7bkyoIPN74LoVdgK0PEmMeKjwEPBmFkE/Tt0jigXgJbyWFKVoGbpL0RYH2y7xyeShMEq
zkkMDWVncpjMMqms0RbzKB+yqBQ/H7zipEW++nSaNFNlwtuIdDzcwoWRxCeJXHDtz2IYss+koXqf
ORDspMnDpF6Y/gT0gGlx3l01Ql0rj3+CHyN8UF8SYxqE8/rkBUquRkzItWeujaQY6h2tY29pxm54
fOVZDKRBne1eTdkJNGaipLGdBipUK6HIP0FLpK9bMnGKnlULqHa617vYYSj7350myNzj83VXvJoB
5G+CBkyeIdbmJJd7zLxsBXuDJPrQjNXcD26v+K9oq6HBhE9M3BqsQvMbY1cvURE3LhrRkPFXgf3i
GQ12wPGSyejwXw3BEDQOa8nWzXI2oRtvEuxPsNWWS6AfNsP2jPp3iHvl7yAmb0TVP26ngb4h0RfR
xHSVF8Y6pctrCTDtcvlLQVpIiraq8RKmCF0p1sOMsw9VXtu5Chwr3RzI5g/zA4iRxlBcB6Tcx9U7
Rgs6b//k6SFHuW8QBLmnJG+FgcSabRbOYNdQUKB0w61/AnWsQ1mCgEhlsLehXTeB4OB+8Mp6ptUV
t5+r+NHXB+eBhq8fQxzFtsdXtgqP4JbCwxZjiCKODLXSVw15i6TLuPnAlN2+hKJmPrSYrmDGfJZr
zS0TBn14D3VE2NDS9bFVovoLE4J2mALTmHS2iYzE75j9ZKLqTxCH/HcO3v3TRLzJQberyAuSw2Rz
YN1RXz60M2i99IV+ifdz5cE5EqAEtbvN9gCWaN5xOkaX0RRyvG6apVp5//jVC2nrH8Z3dpECW23+
WxlaTeryMN8clUs+SJXfwQyCrDLhGHIweuIMGQZSowkZav6gZyRIOmNXRwVSBg4DhF+lDW9OcwrP
Qba29LpIqkmZAy8xoZYzsAKtO2I8LgvbAGEp6Vbtai+zXZNAbRCXc0IU3J+5yvggs3hzctwH5lRi
3C1ym+XWSXo/qclKrkqmpi29ibBuj8YZOEG75YMa94qkStXYMbwlBEIZPuOJrIv3z5DjXIqKARV6
qO9dbLVIPBDNJ7C9tLXyxy/TLjdeeh2HkhnDZPa4ZKNXeg7WrIyANJ4IA9kmo/5DohUGO2q4bnQW
Si1ESd5uT/K869A3PvpXYh9ODGq95bq+Y6n+j7j3f+6wzm0DbVyk2szDNxvCYPcA9K1aCZ/NthSs
CSW5PIhtcZ7KlS+Y/sLvukgf+v+hIpSrhYKXySFoi5gXJq6mCpsxNiZpg4eyB1lhU1AQhcjbuO6B
RvMP10YphAt9RwogsBMCUJRANnQpku+33KZJw018H0OHbeEBsgOyT8zOQXjMOanOQWSvW/B/PXUJ
a/6BY/pdajeB1vC8iz5Yq8cYrBoZ/HKtxZui/tKyU40yEIW/P+WhQQWHdtVsSz1HQXNqfZMUZHdf
EWiII56JOUaHHsPMVhSjgBH1Q+BU0cYBhUXbGyCvMf7a6edn06MDJ4d9PEVgKqX1Uju9Cin5xGzu
4i9nRKnbBPFx1LlNXdjaKhtLzUUwO+4vTbiXF3unLOAzraE5fmihnZl0Qn4FijqrIV7JeLO0NOcL
TpfdTC2gyGABB/mAIFO/KoeW1mb+bwwJUzhuHZ5mr2LULbqjec47JQ95e5BlpGpydN9gV31QJ7WI
T4Zfnqe2eHMmUd2+58otnHmA4mTOHVZC/2YSiRy8SlHz6oyifhqxbl3DZjW6Dkv6YIxZyXFi3wjT
J3VOlDNGHkPi1DEjhkyUuhtZf5joHJ0XrxMvtBVq802fxVMFvPxwKAHH6T9J+g+LcnxLbsSe9MZ3
6BxY+rWjNflCKRb12a94ky5LeZPVbvSZtoSbC64kPoctWHt8y0c6t89Qn5UpVHNCldUQxlP9eL0X
rCW22rdSnLPupy17waZ7DkOlhdyRkE1rHw19rmY6AK+ACl6lpxL9fH444/QdOgCcXQcvL93Ehvpx
ZbtcLDqo59qdphOD9tN6ihGVl0XUJ7zVwRMWgDQI95ZiLjFc+peOsvAfaDKVO9syUeaGG9ZXC2Iw
FLXssrFBo8IMGXCwmGCYFUPfMi+x36Zz0p6yRj1aMQbFXDFPQyZu3irUOuErWROljKJso7mpIPQU
ROmWAX4qCBABf2ZZNq6qxsSokfvAh968aGAq7V4y5tVXcSrBpPc0O0uaoPP35syjnqNKVydmH1uJ
PYp8mIO3S7WXW+DL2mq3SalgfzQtV/BxD4CSMb2HFruLC+zEPyqvy6ECEOiIX2ElXpLz/d5G3z97
TPgLEi0vwzdvFpsRYWyQ/IbDQl0q7fj7DB2BknKlVDJJ3md7P9n5nyXMf4ccklsnwBAEWASB87L6
I1dgUVT/vzBRx1nwEDyf+/6QBVXPh9rBWjZU/2OWkNqbCWzx+6TFhOxDWOhtJxngYDwix9G6SMYn
AGsZlSOAT6oGc/zpDZKhFYBq86AV5MDFnGIPkPfvXKC1CtVkQnfAdDtKGYn4K63FHzi1xBxxfiNZ
Ias3UoSOU6t/eqgLVzFTj3VAxci7cxclJZud19Yg9hPzjy9uLr3D2pO17WaMpwMqGxLdpFa5pN+A
DBKObzTATSKlc6OaUgD07bNYRe0iDrRWmaKCr1ietYh532nNo4yCARfokgbj7gO+9qRUnF58Oczf
dYrcfwOr2UP5EQsG4Qhb4qT7vMHp1gz7ojpukYaMKeyJ5800dC/bJZHGLmqz2Vz8XL/NcK7bG/O1
rt9JVioj7YkjLDCcVE/8GJ0IjdkGL3uCLgsRQ5KLtjlLDw86Yu2YI+ToW3yQY+hDkplbvift6wB2
XVXgjjai/SrmzipwJ4v11MONw6trL3aGdmBdzq+8n+tyDBpBKpHlfMLn6dZ65mlX6B/m1xW2eHhY
hgQdAJGNmOf3PfZjkLEw8D+RSorTP6cRgpO2B3PFZOGN/FQxej1iiwhtqcWS3qAadhoCxRvuEZvW
FgTK6If5RGGfu4CvrW77sAPkTRybzXtPcoUSujQmRGHVctW0smsXiLXK4doAzK3JvAf4I0Du7Z0d
cbfdOchb5EHsgLf8GDlhbMwTAbwMO/D2DNRkvuGnnHaoucZEG3ijnGB2csb2SDXo1bGEUylKCYc9
uxDXIO+70esFXzKECwxH8+jILcztdJ4/hwxunU5W+UkFWR55+TxJlTEfhC7SxhL3szH1x7C2adD2
4qZiXwIPUbw0aKXnhl3E/QWpwtHsvREWTaMC1eZIgG7/SYKM92FdTrDvKOqcRNRK4d4d4hwu9tyS
xEFKsjUAiXlfn0gewpeqKYk/MRdTzdz/7wa1PflMgwkat2LqMV3Fz+v+coQe1btST6RLWdp7DHwT
VykvjGiTPNSwvVvPK4B2/NK1VuFEIwDsGrUHk99Jjvy6oJNQncTv3/fMzCnFWUP9zjEbC4Om8N4p
w4TwQWMCX7ujkyJMuvdY/gOki8i8Rpzhpmq7jzkX/ogXdY1dePDIXA4xqzJsqhb7uAkpbVUwqUEI
zKRu9O208+cdUaGr1EN5TRf4RX1eaqh+WY388Z521YBDvVgyzMxEdUGzgFZz0P3ikXxzVN7tx0d9
q/oZs0ZqKHAWDz1fUPV4Qqj9lze1LSgdCfSASYNre6nlIco9PKQ/tApj0LM/+n0C1mNK8OewbBP8
BGshbKntwhb2TF4YxEVTRHIpY5YQBZKphSxRgyLI6EJMEAvL1C4Cc8ulQzmtIzGVd9ba89GRLrIf
+I1yvgL4jjjfJIlADc6BMA962J+TlTWiFPLeYsSEFhSJvpBC8YTAb2lQ04bmGdBsq1cqSeEVN2xf
M+15iaOqyNKGzt3Xibuf/wgNRfOF7VSJsvXc6s3ZMxfKhOsnCgJ3TH0UYG87ld7KtlQUQz+37gi5
ZgkchJ/O3O6ZXCkiD0CevUzqFziFi1jqlzgT/ZXUaKYXbnyuUzfLU+EOTzR9LHMkRAIdXowa5Ifo
/+TYGajn+cC25PVF/lQbbkDrX/V0vuVm3T9uhH/KK36grlKZAiDOcgLTBZDMJd5omotm+en6l+d8
3eLf91o0XLHsHsleWHbaHnIlSkdqeXLkZHAPZBLPG2ATRwOIHPFdEJi0QdtsHpqCFWXHfs4ZfezX
ASH528dKosyrplBcUpaPC4OmRFaYhLVfX9lgKeATXgvcyKDueUZpnLspzIl53YM3duWf0kDmweG5
CNQ4ZkhwLt/wAxmm3i0XY2cOWa3JisFBQ5NbWBBZH+DAbLgg9woMm6uO3tm7hp/T5fXVt6UkWakU
7FTUpuyZFVPLVCopctjgtX2RqgJxfVkHoh3ndX5/FNZiFHB9SigjCoUViCBDxYiCuXQJ/Q9Eio/e
uia52K5yQM/KKrqEnxUvqrmvBpWwK0jkB+yslLK6e0W5i+dPGAha6X6z56xgjAKXdi/TBqGabQCA
m7c/TzfqIUd1QfWyTcpXwcnMCMoU0l4mcJFsNC6PQlPKiedkky327+R7lFqZzM+EeAiYKymOxn0v
lgTjnSmWA8kPTWYPRIHdd4ryP37vH6Onr2jry4PTzSPSNHaWbEuvxULINSXUE+k72Tn32H/6JHmc
gcW4ZMArtx/6bMaH/ADYLX8F01CXjVE6ryCoaweIyoEFNiVv1TeDzdcTige3ynm+NPoroxssVXk3
9qQmn2udbj7fTE2MwSTFQFQfP2XcBfYeV72kWziz4PHEZKs38BW9wQ7wLKlQ5N+UageYGkQzcxCa
z4X9aCioluRhQjtJ8qahQ4qm2r8rwcchX9w3rkdKgr+N1ZAObG8Vn3QlmGwvn0ag9yGs9aqa77W+
9ncDGeJh/8KDDkunTF9wzxlrpGiDtqZqwm9DrBje83W26RuxqLhxioJLHt0FM7qn7b1k3tcTdOCr
L6/wRJG4bVfd76vXY5SlWn3dVgTCyc9jp3ydIPh3TzmbBJO9zJkckr3G4FFri5XBtgl7qsSg/Nxd
pFYtMp65cHABT7DMe8DN4toeG39tGCRWtpmSazfSX0jKkIcl8ZAMKDRQLyGB1TmWEyYZ43SkJzwU
FnpeeUxdckjGmOAd03aCTC0I6K1YkjYjcLI2OKlzaKkaviarsFGqsxchHw8lU3y7dpNp2VMxE3G9
sABZ8jVllfKkilOD8D1Ag3f8WmFJ3ctiThCOrYTLTEwi/e1IaM6QJUizFJ9bM6RI7/kDOGgpbAou
0HKqzqrrl57UWQ7cqXLR/nZAfcLdJKlL4XggJIEpWHErKZiTqRbM28gdh6Owjs5j7X7Ktz3FrtVR
P6pvAAcTr3wOVcD/zD+xc5uOvjprHZTBU9Ns0SzxxzQCmPtAWlLxlal4DbV8pZ/InwKl5/HfVtWO
QPyAftIMZ6C5eQzU9V7w7l7pDM5c41yOFq306VyeN+XfNP3Fm4tghr6q+0MI84YuooPnR6XKXRVG
vhpdPs9vlEjIsVCb7HCKOR56gwCUKWSyRgGrqKFhCgYwswWvMWJwMe/bdsQETR2rXCEPnNnyX+fa
XYJk9+ISw4zSJaq8znNBQIfnEXr4gorU2QgKyRXsOKzvK4fHYS9eKhRsuFoM5CAXzFxIZ/F97PnR
KOol1mA74yhjnZWR/cWzXi4pSeykPGLA44eYBZAoBQW5KnR9dOZzybHOui+0p2v41AaBYPlOG0MV
7futscNanJxVykqsMBkxB1bzvZOyDtlesd/Q6FuSBMIWLWTfHeD9Y+AIok72a56cPODHvfbpOBHA
QEqjDNCarEcpiYF4Y5LZmavWLE/vjMaEnaWvxB7QhnhsF6dWJSgbePmudxQ/2h2J7RD64g5vboG3
LOUCB/z7tIuvVaYmnGHSt5I+o3clR5f+sOkdkegAPho/9TgvDWGJTwbnHCi5oU/gf1524GvwIBWa
ekTpcOiFJ9vaSHWaiS68Q7tbdM9DzkxA4J9DwRU6lx1oy3LYI0SLJXDRHSCB8KL5IT9HteGezCDA
QJglZUjuF8gAaqAD5SYADRYa8iljVr+S0J5aN4a6gm6oyZxiMRvVBF0ncp3QMSDJ0VbKgzZWT50f
szmwiB5E7f3hRWqEof/dqC7JVJztF9txlb9yW2jay2NnkKUniMsh++tpko9YO8HN5+SAQGPdbZwv
/paYDFgGiVJqCELlerqxZMWPlIeYaRquxzjaB/v/5HaZmrf30GZsyx+eiVC1CFrVAa8kwzFR6L3n
r1of/vRi1ULlT/IdEe22dRFiPc3GEqQeA+bsga2jaOhIQdnPNwYGQPJgS7VOIU7rXW9ssgsS1K8N
LW62dV7lLe1hvdDXFAnKWf+j73CTfERf6GcB8N/EBSyWsuhyzCGTnsYDoZ02moxOYXhwX8WiInMy
8XTdmxjx3oCuQK+faKrIP2YoZPqOhEA6JoVdmG8wcKB56PS561XqM3GBBfeO5fjuVUxW3fSByC23
zl1cAXYP1/wFpIh+mRQEg0jNQIzorn6h7vep53EZMiWpcRPN+7ncV2zLBsZK6gEP5I8TU01W7j/X
3TlFupPk1dG1zYKQQAydVM2HwKG0Mp+BjSc9443Wf2quADnFEvjFfEHHwEgK2K7QJTMuov/4NhNs
fTKRcuMowHb7N4kbTcUNEGZ71bwpd6CoFdcmUHRbQXEb9Xcjqt+pnAuAm8I8AsCHqRAmckyYDU/1
pT5Kkt650Fz34BiZGbgA7aiLCtEHyFBoCRejvZ6Ae4SFvI8oBPDbBa1P+RmxbrK0BPcqmAMypOvX
HzifN/3GeJNI9j4NNO2CDqD1a+8eABgknoHB4d1/kCtnqrJzqVf8LpFNi9YbAzGzdldtwwcJaqxw
UhdtwGaSWtf6vEi5bQo0YXyyhAZDmKhTjOq37GMtWSILzsrmAnR1sYjA9W91/UD4Q83NSQZ2D5/U
fzN7g8idCFbLWN5hVC7INB2liLnPU4QWUlF3vL9mkLuEKTXmG632TBGvYhgLoJ7Ous+ioYvC+/qR
g8z+rDmJq3lf4aTkx+QxQEex6iGnTTg711/pHJYd+iHd8HCI0OUkcYUbyuzoe1j7dauzEthbwRzY
Iu2F2E1IpfFqLA/BkzzrWlmF8snB6L5+UaQ7lORXBE7RHd7h6QE577DoChweY6H8/M9kpyqGxf62
clv5PBJRyWlVal5E6h3/KJtyblcBgGV0dv7MjjgdNLaVpqqd9KjuuMPNUX4BFQjfbOdFSWKXK1Ee
aY2T5xTxM1CMSW/7q2Odk5HrHMEiaIVh6V3IOsdZYftzMtv6LeVvOb/EUwwg8Pl2dxWlerritZT5
km9QZhZk8DpnxjUXBZCuja6JYL6iUpftm/jerUHoeu2k3zW+eMKut2wkc9MU+LcKlwwYkA5BrmQH
aAp7TOXQICn2/mIn5jCl7XJZbe5JDC4IUo9Lz9mzCwP48TAtD3qk2NDS7XUdnz0L7mom6ylktUJg
JRkRiG1jE1hD+8vP/Evzn9OTGJ2mXVIMuUm3NIMBcOZCzW27RCqVrwB+Tqu7D/CTcIkrBwffg5+r
FkTEwLXddMpQn6bGLhxr6R2BYtP5RxIOZdaGtHUjRpFwSyH9rCoMLFBAqboIaNrdfxZqW5LwgWAK
SJEcbYkxueAfOMF5608RVotvQLM9aWbuREE+Q+H0Kil1zKdrQSRukp2x5UjqsHHEyqutQl351vX1
lUNsCa5BNnbNL4CVhd4UljrEaFzHUdlC3hji2pKi21P4Sgk9Mdf+BiG4QklrJM1JOkDW3cI0+JR0
c5VLl+GbdcNPmjnMa+Q9ui3z3bV4oq8yIaOIkDb/iT2dHP20QlMeB7BKPaz1PQDtVQTpjP0HkCjk
zuLaK61GX5p0xVe3rl4kcnWpBvXYnEBFb9xUvMZC2/2EsnVD+t1dlpZ4W5jilUyR/0zunHPL1V3g
kooGvorrp5ggNCdQ7cdNkV2wDjTzcpWMD+ji0IEw6nCcF0yw8sWxQA7lQp+OGnZxg2z97CD5JcgV
w0I/e4bO1NXlKIfE7SslztAmhXfVva/Vg7XOVJC/VWeoiOUtbG6MrgBI6vQeVH/jmk3ngJovMUlD
d3Nyq0BcKWDAvtUPVOp32svSoDub7TooekEU5Nd/CD+Y8LQVfEzWUdm1lkrtp+b5cn8QHBtd6NFS
oLFRjtYMwDw1+lDQVFj1skqnTFp4rvHmS6rkrtDWUtj0/sHZC5S0NzyvvlpAQpTPoUkTj1/VIUDl
Ow5vov8RsRyzQh+Jc5eX3WJvuss2q9NNJcLTbjwn3em6SCBQP0TttqOV52UUZFHWeILw0WI9M6OZ
/3iWQxUZY4GH3XM1Ye+OQdY0VRV5VxKtVq5/XSOAXt/yy6K9bGpQfrClq+5+Rie/izJU7LNw1YCX
nYOWUiRfLO8K8Wggl8MhhyOc+jnUNxtgTwYIv15dkhI9EObsTue1PIMOu7zMSxY1TEvK5Ph+3VuJ
kik88Xzgw8ZdEOjvhCjEiLSxuYspJap0zNtanZ5P7fY0g4O4PZBib9MREgFWLV/FcrqIbD5tjgkd
px0nbMfRr8kiJrJ0iMfC+Tp2siijhJfz/r/wo5CNBGc3QQfd//QT+CvoIg0pRdWgXOm3pY65Fpei
OpaTWJX8lbadeZo6NQJPeHJnLNhQ8Gc4J0HCwu8wQetpkMyJ7DvAv2/uue0V7JFnnC6c8/bhPHJs
2Xp8o2eG0YqHwOitROur16a5NJ4NKFcV6c5rRfeXMTJadmGSIazBFwqb/PqV7IRmfFmwxGm1JXMV
KgpIiEu2dwpic8E+2IuAa3SmxWUqQXjK6vrphbjniVhSJXFWgTx9XMOq77H5udGwFdoRE4c5FX3Q
O3+hsH/YYPF0FPghb9RHfKKxpAl7n61R1eFwfVY60lZYa1vH5XMo3jSAYTtTi2umaiwsy2XaWnws
POal10fANA6qFyqbLdVwNpUOfNoUiy7MqzHGAnnDsR7R0aY+hI46f2XB/PaNrhgXwlM31zAvTRtN
Fio1luwagqJfNg6wKZoKcopAXn5HGNCDLUk6IqDb36Dx9BWFJUlXg1ZwiXpiTACJkKdaqW5CRuy6
X+UhsNvmucCFrY+3UsI878YMWy5HrpBrpLg37ssRjxzSxxeVSmgbGfgzQ3Tc6X3CAmMhv8Ot7/1T
x6Mtvqtlr/IglVM/ejnmvpkRWSdbGiQODRd/kUdLALuP6C//n7WZUvADtZWbqSqAYmhTwXD/upma
4LGkgnaR2Cq2d2TVUnHiRF5wU5fUWOo1LIIiW1SvOI9B0xBhjgr0PsF4vdfsnfHHlvMt8aPyVUh3
C71f8sdyenU64pzd+N8m4yaJBjt938F2v1I0Vo9H/Vw2cIgQS2PgDWZmzUvo2bEeZ40B6v5b6OcD
1JfzjUZgx9JzhJEqo88tn6nF8cc2P7+VsCb3nkOD0Sb83dTz9Jeblg9GlAHH9L6YP+aXlq+zLwBw
+lWqAsIDUEtGg9qH+bZxx2bmRts/AcNHpvMAS+wQx4v5844BOMDZ5lkp2dkogqGd2ZWEebU1VHMa
Ux9817S63gvEi3cbJDGo3jiZrIThofDVmNkYbnxAufJzFKmVVJ1HiNeFsuiNka6Ld1/jsTJtLkjK
zdk2T0GQ+dxEnxA/QVoWTZYYnjgKNQD57tqLB9KeD9JFdoB85VFuOh2B9tyijhKs+TD7SNlIAvQW
Ug4URG9hL27/G2DxK5m9Se96FuySDgYiSqagidVvG0Xuc9/7pEIzWrhFSwvamWmvwB+M4s1AGGcw
q8Qvy76/+mLYQabdwQ5SwV6v81mImfrDgeqDRIleRJnU1CG2WOmXc3avFMlahE8Lxz/5vkap1Sj6
Vy+EKQr56WeukRjUWovlachs9oWXA56Cm80pl4/xyHEQWxD/yHnAUsBIocAwnJLlZ253NCuSXShd
S8CXVWnA1vs0iz2ZOjF4S7aaMoE40Fyfn9ClKuNAH42SRB1TBWI4esqvLw5jzbjmQXMIavKAn0C4
L9GmaGm3OfLqhALZgJTaZUR+gMUBayU29O6PBA8O2hvxO7/pkJIVk3Q+UkRh/LXN1iUgTYZG/Bwr
CY/Fx5fbBwToKBRopJuz3Qc08bZfFBMHm0GO+UHSckDr9+n8fziHrsJ1Vpk1s/Tnw1SWdT7jaIOV
0TsUKBssmwaABkiVGGO4xacu+bXjInktoCkVoeFjRD0jdRSW/oEdJs+69S8ifI6bpTqcAE8yWKxX
RcSMmAUCM1EOj2RFO+GUU7sCevXLvkt623MC27+k054BdgPtXCSYVCjYFbRSdjPN+YpM+Yww0Bio
j+o9ThJyG91kcnREtuJDECO3jgZ79vsK2Iu5oyq5vCnxMG9GTQF5iaU+oMLQ8nDZRmBhMnShDecq
2fOcuFAX9lQ2SLhdFdTSZh9/FCIIcM3MvO3/IZ6DUdtyb14wQczWA82yUzaOYYO0UOYD7QAmevIe
UxObEWodFW227TlttoIJxRm09XOYKK6VU3YRsywgg0Z4hYbv+kYjmbB/8/ZvuJkazRhtPnG+3riB
prjRY7da+Z2DIYB9Sy6I27ok2rLQuX3DMB4GNH2tf3In+QlOcYn1XOF/UQbYiSOR8rCsWJP1fmCt
+xznlF2N1nAdBgfyvP0PR1DvlR3KBHoQkQmtfqVLph/Zf6mX41006mfMJqQI4cExYMDe8RGO/mlT
faEAs7DWpU0CjGJZxBROOaRjt7cRfLSthwZSe8/jakoEnBg9jLr0/bPEwteEUOmfFalQ7mOdsmeQ
otUYbFWxcZMCJN/RjClGG5XxHvJOE6XkQwD74iPuqb49IbxBE479BsFLqRUY8NhRinszcd4Q1B8L
LiEiRA77D7zRyWDg28vZDakCoYXOsg9Wr9RXr3UU06k6WByEVsR8q91Ha5TND4rUmRNGgGlalzR+
yyUjbQlBwcXwT89e5Pivc3AQ1ry+1pP/WClwCP71Rz7A6w8+rXUjRSwF2fXwFqaoKVe4cZol4RXm
QE8/JnhD+N6ch1rtHWEqYq2R8B0kryhxFgvVyCol14uglutBibj3akbxVqemnKOs2oqrxt0baM23
SX/ePhAToy+7gvKFjUVtzW9GdUG80CnU/FnFiX0pdJkEe/F/wKUms6Feqgo65X+MQNKZdhCWZKEr
lxvRWYF5GNNEThrdWmRwwPVlJCl61DetIOXuugVyxNklFL2rq0sgImiyuq1qD9UGr1Yy1um/jneN
zB4H66Ej5ejiy5RFAJQ2WYU5NocnkzDdIt0elpyzR18XWL4t2H3f/TtImL97mU1H8/BzvS5ytuWV
/8i5CfneQ9BwxOgHLZKgnRpcjy70JaK66hkEGjmu31QS3jbo8TIEM6sA9WRV9xizo0rlCw6q9bdB
rRkpWCaZ+3MDGgUNB3cqsc9RZHAgD1tTf/jR7SZrcsbLRV+dcJBiJLBapmopGSXR9jc0zqITqjAk
uzX1wnLGmMH0+ITn/7iTAcRoJ6vhgfZqcKPEVFovNlLEJtIjd69KBBN/14WTB+ity0HDBsr9RxnN
/9h4HYSMMnvtYaZSN1PVKw5DOK8L8JsFNil5A7hqvGt0g+U5DPP/dB+8kLIIe2KstZr+jIbyJWl7
UfyP+Qhr21vWQpmSUFVKsDde3bFisvji2oaOXA6i+owg8njlwP0Agj0D/1CLN7a4H5OTuol9Z2Bd
K5j1HQcGQtjl/a1XoAy3028vSbxwMdWE2d7L8VO5HXHkNWa3gY9TqJRNb57OCJETnhHVU9Y/BPva
Qdp0xmiXwYpM3tCtuckPLj66Nn5XOWlyl1mq7/KD1JH582Pxq29UAzLTMPcO3IiNuQ/7q9sdLE1S
qUUwXf+RtvgukotNYXBtVwADW2NFP2NtvDPgPLbzimjBCx7DmxOyq8J6KWUNHczLgrPcVjQC4RSy
0Ibs7g+GUHZiOM67d3092Ezy62tlfkWO8K+aI9VZFuDydDEDWoPcF/HNhFuUgCV16HQtrZwjkmfX
b5JoCCexuPpbNGVEDqSyTJ5O3IebeExYDe5XRdojh6b4rkBNDWd0IeMfqWk542j+PZ6pHoLfPe46
iWv+HbJzOQ8+b4GdSH0zPpUO38/JlUgNbC5O4Egyc9Iktuuw2n29BnA/KJcN1QhbdkXFEzFZuy5D
ARm5mAboBFAKayT6DxmXl+8SxZP34Lj7FGK2cTJV62CN3anOb6dxpx2JUyHDDC3Nai97/f2A58k8
r//lYnDWkmOYadlmO8L/PdExMnhvI5zGp6GPxlA6RZNFAg9t+P2B0btld50sG9k7E8mLAr7fGO6F
duUee30Sh9UhaQRE/E7RC0LReZEnk4G64+guNh/NjDDkgnGCCxtxPY1JOVOQ0AE4MLW73ZOP+aVP
SIoMc5SgtsDVmpF6mhjf6Uqc5irSBbtZ9r36880VL0bvzavrAZPD+HVfE2T1HOjmc1wnOLfVn7Gf
cv029FNJ6zR+K9ehHmjUPhRNqhnESTNqKd8O9e/3oUDSMH8MJFXW4I6XOZuSlKbVc0/lBjGl3OIO
W56ItbgzG5ptbN7Nf4FQODafInBca0UCw2Jl1cKRXF4nxoyfN9/NJ1504O2I8MvAt8gq1g5Klpss
H8y62vLRvzT4coKbppI7RsRxQwknA7hYa+fTzvJgSyZo4j16tSO8Rfd+YysuQFF/l9lZ/q0SiYtg
FxtmG2i//B5g2JK4vR0CUh5az4a3Eb0HEpA0HVdktHL8945w5U650weuKHDzRsN8Knk6B4nNUdvG
5UjJgsCluTEr/F2dwFxGAkKwnoz9yF9097hj8YeXOrcrrrRDHu6ps/CZaIEh9ttypbjMXWGGKNlE
8Fo2VpjLFv+jeuasfsYKhfchsXkYOIrHiSvOUFEKRiaT0GiqRynuxgqy1hvbke0Sea9/LB9tosv0
Lj7AdC74XR1BLM8Csi0n/0z9CUknvqbv43KMtV8Td21aqWOpwwufKKo0XpAtGuJbhHaYA/EnHq8M
YboWexFcH2oa0VkXVJkyfXbKxyN7f/F9O1IDTzvQRPLhCPo4u3i3y4pPCI8fOTNoTgDD3GUIQm3r
tKqXd5oCdq6zs22zYiBMD8wXbJOUF8M0eKCCUlKPJdBzh4VOp9VmSjzCDJVYd40Pns/klDlDTKzo
FyeS8Llcd6qf4+aGyQnKE4z4sC3J/HQoHSiKfY3Qzc27HZPGdKGjE9273iGqp+8pjSzWKJdppZRJ
yFHk8CpVhPqDtoezL3LIfKZj5o1EyxPnNIc7AsnVR5M7CC4479xXBqV1dIyRWZgo5LMzm+n6MQQ3
oHDWEw0N7Vw4S1k2J/OeBtGwdh+EnRoJs9rx1LSJnPslxcSkx3CVX+NNM6apynO4YOiijvE09kP7
YL+syNlZMu+of0USrY4D7+zQZvjdbO4YO5WYPzYKAGUWQokwildL2uz0grvIronIwEw2c3vd29YT
+5XcNhuuGDKHYjjdy/gbKWXztrlrP5aoQzsexnkFD8oaOAAfiYmRHqGnF1XfgZiV2iNgDOdGXo9p
EEHEz8HRZ4F4bRum7Mo9DcEKVOp+IrO96ndYmOlFiyUFQCbzs/JWIZ1Dj8Fx7fbO7YlAe9OKQn1B
Hrhk7ld/qgK94cUDiw8tY6rRa8zQ6IDRbzjF8RB/j98StthQbEQ1HZL6Gc2sXGRXLYu8Af0EUarr
Db8BnXeZ6GGVGFwJvG5SuPlxrp4CZfSO0JzZrlmIBjy+/fh7+Kj0FXour1koDxVkADQd3r2gykGN
WA9h/qSO+hHot/IyN2WQQYbCz38IUnr2has5q+DOgy5OVvOls4JZqr7kCclnjjxZbhBpFvCngUHN
e9jLfThOakxLgqkQs79Df5ep8xa9xlflFTEGjIpaO74BJ/klbP5GJbFJZ9iz/BBucO9CSdYKv9dc
ro9Ad0M9n0Mpj3mKUYC9X6dUcy/0RznWfAIZE4slSGLk6kyHuGCg7iUukF/ORqcf6s6FpbhxdsGe
T9ejUIdy7Az79QJjBG6TIBQdIET0/AXFGS/nrtZCzPQkkGpHYJWAVexh/g0eLAYSN0/RVKCFxTvj
w+xxYa3dIC3o18RCSjU76dK65lbdxbtNfASq2UaOQ5R3sw9XtfqSJEcIyhosRFIGqcnmiNkqSfGT
WUlGjGjOMiBTo4MjsmH2Xg2Ohlhyc4UFNC3C45URgNk5yA5ydjrSwvOwAeC6/EorltKnjNc9Asvm
XoUsl20fo4MAlJ7qNtkUxaHmvC6lZi8Se/P/FooYxF5+krxjoWDbUyyV0vDZexOLwukPj4HhfQwI
tvN0birrJSkqttuz+wC+c6eL9vY5uGwOw/8iOtyjjfyfw0NTK6USnlz479Jxe1Cy1G0oS3e7o0wn
k9GrwMGNaHni0dn6oLQB+ORYxETRwRZj1/3lLVoRvbubDsLjGy033sIWNnVAqgC3DQo8a/xCRyqs
NKV+H0k1CNzJ61UX3GmDlbQabpunjezITypRubINpbLkC+yHfMV1xzYwxR1h5yBxTQQfuRSo3r45
yN8rkVLlF79VHkWq7vyuIENWAJv2d0x/Rx8Z34bAiCG91r7T0mFk5wS5yxIQ97eOycQL50Zd9Qbq
fIJFj0J1WdWyOFAdyMdnT0OA4sFHXr3XIwtnnbbmQYnA9OWayADYqLmtl+tqf9yVNv8ANvG8R1ee
MSWeMpXhlD48G5Ml3PHQNIQxMrtQgPQX+fX4bLC2e9/B6eJNg/UyMZHJ1EE+DTIC/vmj7pbKZ54m
/Zww/OH4PLvLc0AdlvodOiBquLKHFn145JYIjyVQIaXOT9UICN+IxQZAkxHcCHptGg4QFJkJ+TL2
GTPELHi/owntur/3xAxn26W63b8maO61M+skDERPhnZGbzBqY1rwj59CDTCNsnO/cUAGTpUG5Agj
6f6DbrRDhHpbPYb9TtHwkfHckS6oE+8WjVS3fhq9nuIgr4NEz8fccjbscNe/dkIxraZZnrgG+iZZ
UW6e1sLmjzq7VmMzY5VgbvtU3k5/+7yt2Hpt8VTO/lVjPd40clUM9UKVtQ8q6j+kLM1sUPQWwKjR
f7sPePNTUEWximtelGSX0VHJV5n5PW3uplY6AxpQUzHYyi7KRsYh0HigTrYym0aq1rsneTIH13VF
kKRax9uyilUKfzmVtyKxPy9T9PFvaompcUJ5087guTw1ZO6DrJBjdgFs9PrTxDVj7FN8Vm74wqhN
q8pJECBuDohyYRD8ofmPgtqFZ5Vc/gI5EACvkqqZQfjBdxuM3kKXbrcXu+5l16D1isZiJeMjnIJP
tbtdMKHyVGlbGJANOYVQTAQbiDhSLaZ10EqC8qZZhun+kbXgwPXGjEn0Ntt3y4J4NYWXR6E5wc91
YCpYunOGDiw4sEQYTLCZJx6+MDqX1H43GQIrYFTopaJ9Gq21xByVt65c3cSyw/NBPaJdGuwz1xmh
lUlAfpSdRimy3OT10iY+UJqCw2FxAbFijbD/3RMmEvsiZp4eHzk0j7QcbeXpVL7Y2wFZXYfjE1BT
M/EnOfLxttS4ODQ0lmR7JZo2AKxOjfBHToz5qJtxD5PAXQzRD6MaSnMLrGo6N4iR85jBpfwMe6AM
bm7E/Gfk4aIG3iJxTf8lekZe/fcBlkvl8Cgo1Wn7+RRx0gZruaPUnRnMBDPpZQjotDkhkTWmnpQe
m1cxRVmQO05jifTFtXX7jd2BZmCnMVV1MZW7Qy6MKkFnOgMTjXmMYC7dPcTVAhsJyeGmSBrLPhPC
QPoDn483TNJziLlQ8U+InZ3tC2kiBSGJYu2vlwvsHHiZfwszP+V/uRDPk+rgP9+5PPXWd1mLwYPC
iTGAnqd1rslbKkAFM7552YUHXIJXCEhsST+0ni51PKlFYvcQZPVAqjECE1q0nAG5dS+kW/FEe3Gp
ZeZjVhgkI/j5f2Ksqe+ST9zCZmev/1afTYKOFeIS1NkqE/uEHvmZMXyLxzrGPZj5BqQehjEUicm9
uQKs0Kjgf7AoOP0BbmnyT1Z0/M0AI9AOWlTMcdcfkUp2pWEYsbqpH3F8yF9ecgj5cExUjkk4u4bm
g83Dxb0Zp2h9uV1vJiEiaBvkw8bAM++bUzcvBky3N7C9qJRI8uEB6ueiKiz/VJHG7K6ZE4nsnRb2
gebs4xNXYSmuTjrMWXRz1v82ULY1yUCtIyzLHqWd12LszPK0zWvFcnZlkqOFRofc1ES5NWuvEwuv
XDmwRuPbEa9kNLlSW1JP4OxId8V5HAS4qmWtfUDOhFCk/4CsMpdVm9bvD4KDVm2yRHxAj/r2VCOH
8HcPXjuCEnhadGE/z0akokjZB+9ThHhhSUvsvR8W5/CmL8kgia4FNLK/aLPwgb/ymR8fJJhfqSHP
q2xUTSeobKtfppkVnCK+OYjs0taLe1+qyZazqSeeeQBE3sUWmZ2OHw9GvuqfCQCDWFhgi+jrX0Jx
L6Ephcs5nxbtirfBk/bcGchMaWUg4qu6Bes26uFq0s2218o3yHj1tc+RkUd0VNegHGA0ExUmPdos
jYp2p1ynhhBPMJH3HUOvVpDmSf1TQIYvd11EDM5OBd9+cakWo8qqDaltMDmYKsojmGwyjOD+PEhv
PAASza9kmZ1Cc6AsEyRLxudM0zYB+scATRar0x8mBA9NjaZfAHTX23LeALqu6soJUQuSqqP91y+f
pn5IjLJcCGCBtcNE/0Ywa7YlipKIuI6V0gUOCE/fVQbyRzwTxa4Dyldli7egwvYRT4uray7Q6AxI
3FBcptyxWeFb6RNsFNChJiKlfmTD2hw6pz01z6urG1fcM/pZe8dLDIbmw74S7fOrYFfWZln6JkH8
/+tqnjoixvpsvsLuyqIusrxbIamAxanugEwy6k8uWGuO7leC4VtYFRe/5o7up0gp4kBFnMhqBFnD
HCpQ2XciT+yluC/FnSdM0mBy0NwYRF0TftSYRRNy6gd4hhyhEgzRMu1vcTtI4mJaQzQlJVzvbaai
bPulDaRQ3xA3aoqqFnl5UWM0gk2UHV6VwmcdqlIf+vHJ/MSK7i58Id26/lGyCD5OVXpDV9nMA9+j
Dq5pFfn+PeF1t2Fa8FXWrQdVazRd544SwhHykrC4py7s02rldxCoK6VPkV9TYUqkYokqDQNrbNqu
Nu88Zt/q6x8Dm5NTsTlcMrqB7lvQhQ7LhvmKI9bNWHEzZTX50aJE67RK5m6J9HgB+eF89dUvnzz3
F3Sr7APIsoT0qYfM85euB2DTt9E6+N4qyEokYC9d9nAn67pvaAT4eQTuQEnunwMk9v75aKhrL2rl
YSVkv0FctdtxPWeFdm+3tbeYbywIP7IPf80XMQRVN6tV/gq4RI0QjxgRIB1/unLLQvNDcwldK7ud
9P3UAHnhYTQzY+r4ViV8fHcuRzJ6PXKTS6cMlbR6YVDuxqHSr1dTTt8fAwFrrv13AsIz56HmUgtu
HGhqwHrdTjK4KdXB+66pqjuVyaL3ilpmgCAMbpaouiXyZVDqmFyW6k1GORiAMJKr4GuXQJnaQEfx
LXE5Ga/TziSFcKGOINcv5j/6jCjIQ2vdTh0zQLvC89p6rGsxRXUw1uOZ+ytMAHaAHmJu/sOpVuDr
Hu3dZHRsTBj57hFFB9bOScL+qYaii7RAkOhUAyrSo40FTINUgfhTNQtebn99ZQmNhN9YlFtdxqze
et7yRhk2G3RWCTtmtSVvcCPLwL+81sq5IGC3d9YEpQxLoTm7elCZ1/uSM8TWD2x63B9ij8ezGprJ
5sYxnwTXr6+Syh5Q7HX9P5LXIvMZvppFMpsA6wWFwQZFEyt2yWXpPcwEV68Ju0nIfQ7sd9O55sb5
Z5U2vpna2VOe/TekoTl63OlXm7eOVqdx5nFXQe04viTNy8FBh+nmS6eLCu0RJ4M0RSjZ1F405TVG
LQVg/qwYEhzrS7Qa5/CaJl5uUjiUE4gqiCQKc97eYFoqvt0Lw9nbAaamXTUsaHSZaz2EIQ10RjT9
ZCi+XzUOnVmZWzEu0toYDQK4waXcUmU22hQIimcJdMJzYFzQaviK02yU0wI8K7ytnxoqmZrzgm22
zGAMjJP3h67a5SfK2BS6OrzD2HYzwGLfCgVnVEFOIUq6LI0iM3iyr22W8+9aExiNjcioAnB/xwz4
/LPnnBvV9hix/sVWj3xeSRm4kbwYOsuB30NyQNGCcuzPXNUIjSSyGRm0ZtJbFpTQZzYIEJerWrA9
d/+eYpffKkwkg3FDpVLpAS06chFNUuu49ZpOfVQuJa2Qiyv4rYvi/DNIHj3LvlnMn2IjSk0d7BFb
9WdsN/Ox8pcBQ0forIBBMWlsXXKrutSDYsC93414IKcJiW1JIlOOO5qb3Syzx6Vw7F+np3zH/fdG
X4txLIbBhcVd8j4gMxZ2S9SgzBpD1f/Wx/PWEy7D/7w7B4S2NDycTnzZ/FC8eZcKKHg7z7OK05Os
Z4CCkeqzwwv9tLnZNxZR6knEbAuo891b07yo/5cYkZLeTjIwv4U0sbS+evFuU1C5EnRv+Ao5qH0H
G93GgIOzUl0elZU6BhtqAHzpXlxbZuk33mMMKB4+iiPQkhQFCbhkCigwDPRfPy73ZIfdVO9eqcUe
E0c8iSy3C29x1fqiMDv3WF4DQkNsVKxyp1HqhbCCwpg78amnVKcyiVKr1yntpWbOOJzDi1UltbJL
Df41NirL6gy+8XC2xf3Dd9s18YOHuvXzqyclhCh7X0lL8EBEcwwZmXd6B0NglWUn9DeRbYhvw70A
R2BqNg6i4tc9D4TFEvn1cAqne2ECMrPqgSH8OWVHEtgVn59Mc2frJqbnSsZgnq/sdVqlmYvf7eNU
LhZMQ8J8XoP4ub+gHuHZ9tL8JdvUm5lR/kM6GobJwoCoxTo6lssbXHCW3ucZMS44/jGfOcXijOzb
4ZJOLEr9TephV7XSUFUvHean/ecBpXytvMtnS6oK9hQjRYgCVfqHhl8KumduUV31jl35/fzyQ+UG
AyPfHi1Hn0wUb/fSAm179vPNGyhYjuEgDjh8lRdaC24ea71JALz/SsNyGkc/sHlAWImKJ1WtU01h
8+k9wt/jNQwA6emKvDdKZtIK42awcfQ/ffeKfcMzgUEzDauyHhW8TAcv7SAEBGxJVZGGg5/H7sW+
963n/4KQ5abKDgtBTI61GJGLicLCo2jrIqvSYX82EvT+LmkrXuN+G3MO2nz8Od/jnFi6sHKbXlM1
bDtHqpFiSw99Tpti6a4/l/r2Il5Gt8Q6M5Z7sFNZOQ48c1CYhXuNiu5s3uysS6DbrVWof4Oc0POP
cDIPbvc0M31sGnDTf9uZz9VjBDpGjFwJn8ce2TvAhbIn0H6xZ6bOq47qq8+dJ+5WO85ngf2FNPGV
Yk1HvjX/7UJyMSliPSJ9QrDfngQUkls8Wm6bU3Yl1KnboTm2TyuZNRk9wFbxSareEF7GCVaDNa85
Ab3IGbgvjtWj+cyzuz7OOdYjtHqlRdKjPgZe9ZeQREXndjzMTu6hcFZ2uZYLDi1OuLJRrqU8+vdL
84FNgCD6ne9/Y8U7lGa2U0pGdFiPVusqNzkwKXZGksGwswF3WQa7gnSoB35U8CQJ6gyfIuJOBhgN
Deyz8wqvP7juixUDyHtvUAFbMXdB/td0noFC860MoKN3xy6yTCd88RRCoPvkMwvwWHCV8n7aUP5A
d48Q7gG7YeuhvKRSs7RvhhLp1gTV7EIRCGts4QDcHAY0uiW3PDDn12rdOMLFryhPFB7g3XBad3Il
iGJufXcc/8+twgsBHVsJ0ECrTkXLzFO7k5SJNL2kUQtLZEjx3lNFM23JFMvjnvEzhOlN9svMXbrQ
28kd4FbAbHAGuihGzVsRV6Gknwyf8Mq6HVrumwDOUdp6MN9H8LaPxPmeTBKSguy3cHQT07/EFEE7
xE0sobMzww3XQlMa1qeCmykUfUox0HSmH3pg9iw28ALR2Mt5jYOjhB3Y0DsCD4ZIc7hMUs8G/ECk
22FIDmrVgqyHaOm/xAGrRS+BwEiVn7hCZrrQ5k2zvjfULEdAOMB9RQk0bkMfKlDeQaMil3aEGZdO
CDUvysepWrUKJrdg0EJNa+86rEE3Cu2dJ2e2GJtG/gnnhMk4sivf6j0o27BrGa20mTkenax/IoQ6
yqll2NqKKVT60fmfZwe4L2oR+xLkcWzTp8rV8NLO0oR9zhJS0AdDxomhRj3cBhDN0bxsB85JmSC7
QTueNu/gKKhNU5B5i+8h1DzI6XpISyjeQL10Ys3aGrNWY6EeLM0C5RZdBG6IqxDzSlV1+SbsvtR7
DpVF64FJuHc4oQiBGuJTDj9fmy7PzUhm41X7zKc2vXiMXA64iAGCtsNHBQgUGytIMwwLDkfzMqoy
KrOCrYJKyB43x6qeOdAS9WhiGR4nMtvn2kdwQpzj4kiQ62GHNqxYuvqVHAvb5bZs4UNLRp/S1Uoj
ewOO1fdfo/jRYRTqJ6btvc01Cn3EnbXw+gWNFKZPa+sSLPSvsqXwRZVavMoo/HHQ4dfuVpu8a5QB
akUdP97Sk5f/b8BWs+ILiO4jZlkaSO43RaiopfY5BB4OZxK8X2WJWwKv/oMfPJ0QNuO3/RYOWCAr
Rg1iYKxe0wRv/eIzr2qwWBau/GJx4ipMBuNAPDXbgfVRKOy8ztZ+WNf4I8z2ga3RpC5nNJwd2zbU
YVVEJBywM8l+ZHplbvlYpmZJTnugjDuTfivmAd5CRkSehkFK8UakKx5Ps3gGm6xGxfM15EQ2FM4q
oJANuW4Y0BPnjm+aQoBEjG0e0YZCAWoPt/9AIPn+TIU2qapwBLxhZ0TR14bCtJAmR8pz4IVqxyAy
40ihVmMEoYFeZZXMzVGjZWt/Ycn/RahKhweBQQOedef24Ynze8VgJPgSHxgpiMEOk08g6pJFn3qB
jkhyzQ9bzCq0Sg1sD/u37OTUMwPaxP/Xpvjx51j6LewLYqr26Xna4W6FkUcevhzYwIhML3SyPAR3
ZtQFL0PmfnPYc+ASPDukb7yRmQ/xInHyM71KeZ/rW1QMBRUEh5x9LRRyrDd19Ll7UEPUO8MA0gmi
JPrObo7uMo3Chqm8c8Ntimo5qHxXtKO3HyXzmph7Y/pPiCT7mUwRv7lsaK4vW/1vdIs28GUoDw+4
TPHDfIkUIjaCP/IUQEZjGMDZfiF9KDsWDGsDz4qhSZp7+YK6MezXbAX8N4pvhdB+obiPb7xyG7/8
pnTKjR92K7VnXeDiQqF+gavPzfNVTs4RqAB9+7lfUBppl9YH+KjUSGdT+31Pz16dG+AMZ2Tlzgpc
LK0O6M0UtwHKg2owb9PdELncZVMyuk4tSwbuOk6GKLCFq5JSIpH22jHtX2C9+hFtQB5UKJiNpiw6
DjCFAF09E3tUUOcngYmRuaTIud2ClovNuErWLtietvpRQsnz69qoGD9hOtmXIjfpeeFcF/1q3UOU
pKhsQ9GJ4wIoRYvqvq/mqFa+c82sDyNOA3OFuWlutBG7BNLvzPGmL7kAfR326tUSBzF+C1hjhO6u
w3q8G4Xj8FEOPMCMqkxu9+jgFlKBSF7NaJe0DeFXfN1D29uj879fKrNmCWREzhXU0UynLmH98jxK
pj5RyTmzi/vkOHpOXadDKkLg6FpM/d0uh1cGiG5eIFVuKCPt1tpN1Al7h+YKVleb1yzzJZ4dSIct
ofX4XiaJpYtbaG89oKaqV/Xp15qoLnLpvjYl+NWZoKYMktagtXVUgFA5DkELgzM0k+ajRBO63JZ/
z6CzjE+0Mgr/LsMkMlg1N/zwwYQWgMbYHc/qAWplr6LWNjHEPkLa1EugheJ7UHEhpuTSUty/4yR3
Fc7ar01eagP2xFvP8TBtSLUNh4y0irp0hIH+mHFB/3He8t28kimfPW97jLr84++SAzOj55+728D4
Gp+LSOowK68YXRgMLjbhD6plkT26YzdPSroGWNH7qkVe6hnoRNUWZ3Nj/wzhLrCMSPk1JGllGFaX
uAAFZzjEOoHV9gjBk9XrAJL1l6S/kau3uJEtVUodjyQpywwmcL6cifeDeMyq9VsJFh2B388Ed1Ya
knxlNKhlUvItrbFdD6LPN9Ya39rlDVBKuiVlFXsjNZoZ0U7gt02N1JU2qqQLjGTQWBlTZCEN/zQT
yIfXnlBddoLd7Vn7WgdRQjho/12YB+Ng1sZIywc+nbjE7J3QbsR1PkRkNXfQmOp6vRn5s5dPLWjp
eEvTDG6Vn1dOlcees3rGVGlPpAWFR5bVqKJDubMJUyTzOVh+nyZrRDPhoBq3MUfDg/1UhaXuabHp
N+MEenPn2bxZIRdtQkwtgSY+gX+3wNjXFVnfkp3iQ9Ig/Mou18izdEctTlxa0N7xYuaOAzqxfAfK
INm8Xm3C02i2sLL/5WC6gIAJnd5LziyWY+42h7lRIM6OqaoDOqhKRQ30gL9EEPvKygj37egedTB6
Mu2L5ccG/msJHG1LLdXzgAeIKvhIIBy9hMdYxIR3OKcaVmGP8mQH9R1DmyUy/J1M73upBZcIa71a
GQG0Gw/z9SY78lfkyYqwAmyiTGjOaHZvRzyENFw82YaG12xls+8WUiPF9+OIHvHjDk4dYq7ebgSa
9MJinCg6KSpkjIGnpOmhrIXXdCljRG5UyR4ZY7tINwMsDnIfPkUUVhZA49daTjGEGLQdqi+5Lbf5
BG5FLrJS3iGbdAniIOEzGa3h12ts41F8IpAGmJp5Q/h+0yM3YCQNHosdFtDn2imQ5k93H0/D4RKs
imvczF34a6DzrJkLx//RJq4EPcZS4WmxBd1DswStijFHCN9KDvEW57zdiq2afnHMM6jBIVtyp6J3
FGhAcgtP15dckviWczACRVfBS9YAlfGV0+yJcT+D4Bs+PSlaIat8rhddvrSjvy67UXx3Yvg/oR0e
DCDkT2LotB2tKKqj1WlpLNJDddDroTBfdJVhYiNkoV02yNp1BE8j/4309k00cZHPOi4b6KnZk0od
pAtdiOEEimvaQFwgvcxC+r3w8+WMlQnJodq7iCsa1MdG6gaKGWnl2zhxqqApxoANpsU9DxUw9O2M
zUs87TyEkJp0931gPIevlTC6UiZi9ftck3GfmDnkflC4tHE/VdgdRFKA0a1U5xpyx7xjeRSVKpoF
fI4ZDbEcDRnlfSshIvxa6HzG9R1g239qqVxA9kPN57m+48wa2Z7kYXTZ0Wugu3Fbv3cWPBPaeCGh
FHM3aWHkdnDi6SbkbQcBa+x39nnffGnXDFRBwjT3nRwt8NpH8AJqUaeWFeCEw/42VZEo9OAC6+W9
Sj+40ufV5GvCCD4B7nXI1xjLv3p3jtusbVnTuJGBwCh+xn4aA5B6HhVy5jZnIFNcsJgCcQNiHr0p
oApB+hPqDoWVEbH0avurY7vgjYJWP7phvv7YqfFIkuT/vhuG+U5+qrHisupdvdv0OQNUv0aCEsGu
MnIs9ZlcPXQA6T//TzvTZ1U+zqYG+crL+I7b68oo5s++QHNY9+YKQNVxJqxSjJmvtIxh1cyjijDg
44Fdy4z8FxIYM4eYEpiWeOFCDinDT/KP68xx/Xw/pHKyTyTkPEJXLuu/tZLa2VIhLSmCKJeLFy3h
EbrWMQHJOh8vwTsVPW32xSVk+9IzvdpN5Bqt9Ta6muLd7E7ymUuIStfp3LBWI6PzxmCwZyCFxpHp
b8mmdUC3hu7xwdkn6oQ2AOOPqMf84Zo28h4B0pLbXv7A7a3BQpRzIsEg+6yqd45fHiJJTqzGc/8g
+L/B1G8s2xeYGg3inQbtG8O9PWAU0AR+vA3OGgkb0i4hKpt4Ymb/KjMe5A9X9FtiQbe8E9i/rqKX
eBZRgObYC9wr7JStaogss/VIUsAouhw79SsB8wGx3VrEVzgTWJ0Ydxx2BAOGeACP9U3JtyENlD4w
kh5xYrtcb7rWWnwqCsaPz31aeHngaaTcNFhgrcEBCYpwwROntLNpKqBDqKHvZqCqt0EYogiWTjHg
OYn4KZnujp+0tbd8AuIuCuh4xesUiLnib8MjvstBiShY1igiDWqsOr6gMy6+NlwYyNuEHcXtY4p9
3jCPVGEFIUdLq99BRcxdtVozYFnra2JyEmZ9MguVeJu+JxDC+wqzZr8RpFyfKut/LersatbqpP31
QggyWdTReJ51Ii9Ik/ee6fJme9hsYwGwCogWIA9ASjEvGoIGz6cSjKAb+GU2A7O/HC3loszPEQMg
Rhl2o7c9Pk/N0nXDRqagirKvavfD0Jd9AnI+v3An8b6uysGhzjRbXdlg2HtixbuXWjL6jLaKKPWr
7JfseS5QP+rgYYAwA81n0T9yX5/rvEZE5U5bwcsQY+WQIA/0MPW+dH4hjgFtME6S7bgBsqRfr5Vc
ZuYsb0X6dzw9rqGPhhwTYpo1qXZq5qx0O9Xj71nKIPBTf+5kQONdhfprinsiXQI+2LDo56O9zq4n
JVLgAXFRzipBMwfPYV5/qJS+tAtOWyy6bomEDBlkQGBUoyEBd6IWKaw7hnbn6BIg2txeuPwd2kSH
JmoeR+xnde1piT863ZQWsZXQP629wKtQA32UWIMUMyJTx1hGf9lhNqXGa22/H3ZN2IPqR3zjZA5E
utuj/NWYKZtGQVg1uRmOEu2PJYgKHbtmP7/ZKyctquuLXV1J/DkSfQE+pdiFvCJPvfMbbUwG5Y9w
2Lpuw4Jhv9FcjoxeBsrqJ12txsf97Hpkms1mFAx2E+bILHTpZfW+B5XwhOvaBIB8zQ7mUtrrHIwu
MjVoud6DBoSmS5eBgN/l+J+5QcCZ9LaIHZS8I9j6vLhCgf2SC64KdeJ7rRhg18aT99KLKaXWJXiA
XQ6oZQnQLeGo6Npd0An5RO+QJcg3cLmZYUcbteaySY/2cYN1y5cOX8NGr2dsD334LUa/Z47dRca5
g55IeqyHHf+MbA7c4SWoCpJ6Dscypd9MY1yRES0Uvi/se4ok7uUOB2YxdJd7dzkAnkdFocYkFnWN
FP7VQ79F6ZG4hbZQmJW4K3GSR7yLLc1e1rkg9gCpBB0fpHISuk6IpiBeEnQR4z/qCMJMeI9xKlo5
Kjwksak/Dk+iFJ1LmihZzZS1dCWXFA0fS/A/Lp4N0Hs9b4H/S2ao3ZcSWLhSG/EykMe1qOLFwLM1
kQlAJ6EaB9Jga1y/DJl8ok6fT0MG4LEX4zyJGE+uSnbhf0BGkrM8Ua+v5H9sU0ljGpy/5IhcquF+
Z4euIXekHtInlFnMfJnRUFX904mlbHq5m1ptRq8jtn2m+HjHh0OZdDLpaaTAqTbymRCSw0jQ7u8w
T3j+3PpXnROsZsvH8k3EcnNwi5MPqndGaBrKn/7f/zi6AnYFpTsmfTUUbw5Z2jMDYm+Lb6XrPjKm
neSDvaz26U6UJlHCrZNC0pQHMl8pmfU9rE1KNXWasLhbS036I4rBJRTg37Xx6NStkqa+Lgx0Cvm4
zDQO9Q7vGIMoiVe4q0Og/+kk3xr3z1hGOjO6D2rt92oce4bGVyjX7SbsmeILFkufaYPTjWuCGzGf
GUIytcTD81HAeauLzEptObh5PASScb3+rlKlzM5SDMtEFJwMoTgDlDNbTgpd5SXPnWVYbHVXgoSS
xI4Lqqc6erskaKpsII5EF80nRyt2VFlZTcJsXG36fil+KbkNN8gbphAkDXjB1BXnepjTd5e3FyVt
9yRAd5tyf5YAShfyLyisVuoRda14EWwymcLjW1GT20tdT6grkQ1ktIi+YvxnbiGGcPigMHbDHR/3
wFnvWY+zikrNAbiwr/zSurmDO9LjzcgTMB5nszQJg5wbPpLz3tcTLgaH8K3wXoLeipfw81DbNGWZ
WjEcI4uinkwd7n+kIUdd0WdgrjMfP/GeLAfySMX9VdfRDUtHLDiriCAH0MEV4hM9Se3BShlew5tS
jbaDcQ1XzScl+4I1pOOgg6sk40iywKZeJA3MGEYw2nFzsI1luqD0JNDlBE1eY1Xvqf1TKlkTuFwT
DynHNP7XUSorCyKpmBh54JVFAHrd81vXTzvOQPaYn9CjYC0AnVhRqbT1MFKplIXg9NMMMLpbLYjr
MUGQbZBZYOmPgVaSnTX9uYxwNIeGR8Y1vgl7V0A3zhGDOlFM4pBMJJYr79bAxaVcUwiaRALnkh0U
cF78/Tu8Q48QDpz4iDR6XBNRi23IkU1z8YFRslr2dIhCRBGwUhLxSIjz4kRrmhIEbIIH0TtmXmED
A1MXu39nteUg8AyT1E+hxYHN1TK6+w3chxbZT331bqbTTFhzKkxSDAyEfb094KHqAHoZwaGPAq4j
xal2ZtBteQeioDoeFS7k+iGFYhJnOpTG70NFjVxMRybpnCV1XGzUgoYeuwzSZDKqjaRNbAyCLtev
E1ENvF6VeaV9/p+4LNTgRIMlrK2ENHEM5u+UjqwNG8+aXXZ2CScGlx8U+/BZm0B1kvr/spfowenc
kEY9gncn8WTJDAQRbkDUksLwhRmg9NrgqPfPnK54/iVZGf7ljJ05PyOA8+K2wQ8xt0uloGbtpNSc
wNS1JutoONe2VIxt+Lwm9sefopv0ekyw2BI5SY8XZtzwaxlAhG9rUo2BYocpRlo4h1VystMCRoqf
AnLiMgDOIxKMaIYTMedQ6eyAwQqFokdyqlgbWzl+AutLeQMdl+AqGSYvoMWREybfw5mgWEPz11wP
KRmHHOsQjzUT7bdnBtiQtgfDT2yLCQNpr5xcy1gTVH9vmC8gROolVmjO/x5PLEW3FiJ53XwE0SQw
PO6TnD1ZeEjO21lY5k89EoogeEpQJVUecPd4ch0HfDHa/Hf93k0c3rcfaywZewM44QlmTj2kIfGc
Anzv/2RA9mQma9DKVO1Cdo2tLRYtWWrFfCSiBIqyLJehavDzwofoO+rtjbR/QHSobSFMnW1I+jmu
GOG3h8UuNJhMWs3EKaviAdgvOPqOnqrcnTcWUKY+zwiuag4phUVxQ8eBtkxwpkaeFFl6n0awf5CG
QS7xLzkqPf8c5OF6giliiGhtoeyAlrFzLVgx6LgSTlmZWmcNr5eOTLa/hrGsiGNUsjqtNBGoGuVz
xfDafhnWy2m7mSIwFF6lZnISE5K0KoR5GDORV8hoWTudlvh6A6O/XsteoRsXZ4Lz1wKz+POYE9wm
v1ae58UtXJvUjj4374nJrDFgG+xcc1mikS6hQGxqB3mmM7x2IMpiStrJPKckHtYmmFwbdw2y3lkL
5Ko26jD+DZIqzNdD6Y9jxyISg5cfnIvqVtYEWnQMjPUaCVqHcFZ8lGUEDNxRn9dvM6ihj6PmOh3w
fL43g9efTs+5Fz2n2S9wgjwjnPRRpo1mY0UMC4svwUKTBMIEZ56yUOVlSRLhuOjQucoJr4wkDMg+
X8wILFlgESMXGK2T9d6loN4D6ND+XqAtBXWwqKTNhWMg0a/zyT4rsMkLN4295WY/bgguFS/D+sCp
TO24hFKicBHGSP/KuPSdwH0Cz/2zRrTCCvN4Uh+y4B6FVk7EjBfwLjPmjP2FtkcNWxARU77LHtlW
wGMRoTknEqLfvsUJMiUvxOY1bJUmGRg/80eJYipTyadSYTy1XFZ0eHChzyV9E2FZT3w9YTAMqk2T
s+9i6Trqq1jbAeG8QrcQQrOG2KUtnTGJKqM0kzpTfuwriiRy0bEIojhjY46vipHV/9LakC38Tsn9
/3Sb3Od7Hh260qht5xBGjoM0s7PebOSlBe6SXbEDefkaFsRWPjo3awMnlhBCk7i/F7/BPjRkcO8o
2DrUYLPgk3yU3aHz6jpoAnmiEN1vXj85SLepViEnGBr9bafhJgGGrj9OhErf3Yey2/5g3Vt3kFo1
4zvZhl4hUw5cz9GuOZPcERyQVFJppWSYXqJuMVTZyuOwrLvAZEua+Og1zCt2K4E5EtFUvZw+3uVa
jc6Hlv3DQTArhENAgLiH57dESPJX4TdJQf8ghKk35TD6j0MyTRfLcPeHKBNXHZvUX9h9YMr0ne45
5ymOXkwxu1kDPN/Q4DHuauKzB1vw/09Uy8UAZuagbEuX5RTPzNlIFkURr3AiG+bSgwSzqYzbvEpA
+d6BkRLavRuRrKr63tG/sTdua4u/xvw5xRNG36snf3fTJv+KxizR6Bwm5mzDVin8qb5SKmn5wODE
Kxd8jV5RNKi/OESKVMQk6wDT5QLpvMlQEFDr9177QBBjEQQ14etaeBGvtyC3WPpGY+MOKCqwLnjH
66wvZ3egS2qaWhulpy/O3B2t/5qm4zveClMR3nyAW7T1wTmdBqC+oxv/Qxh58wskyODobhtMOQmf
dv5ffjVE8BbSzI5CkfebBeuI6xdKTf1brTipsROM4KQlNDdqRzBvMBipD2cyUHeTdX1CrsLkRx4+
yI341LqsO0Zx3t8urf88WHqppdAmCElcihAy0B3yKAO+nOoF7SNopXLaL1NcHCjIIOiV3hwX2w1M
gSvIZr10g1RI+7gBsjwmWK4z0rFPMrWhg+vRTnStfLzqe/miw05f4PHB6P4L3PqlwHoR7ANowA01
RFP9nm8W/TXPw91wxnGNGHqTwLppxLs0ObRTWbbQ1BuMeybFdWYwxuJhPLVZgvbxjlaojMPgimR7
RxlachIFeQkKWjWNJdGxrhzWuTekfFGxT3w5LpBfs23jja+mbKsf26dU2BlCPwJwVB0ItES3F3pQ
rjpcgh4HsoZBp9Qzk16JvAd2zt+VSmvzKo2MAitLp+OuKneaU8H5fjbDVXYD/eoEiWnTIZ27PI4K
IJ1UsulA9esjo4F5E9/u+XjeyJV1tankadyJcnnt4vMADDbXxG4vHGXDBHqSwvkKo5+BO6FQ87Ew
cafOBqLDTgE0K/ZsvtbqlJ0UYE7mH0zi4AzZn6mx7+tcKZcuw8XYKvYnMY6aviMXC/6OR58we3UK
Xhm3u5y9E7T8eL6yJ0YdDEKQKhm2eKc1TguAtIKVkSOhIih6lLg3DDNBW6ZmiNiTgrYwy+wt0Z2j
HT+15Cww7gNMmNDZEBHflDljhIGuIbarIANrj46GHU5OnEEbddWyvYxVhYiysjJTlAkaPBIe8bT3
ZS8fyCxcnX+6m/5hfBjPnrxx+nLhssUCyqnB0/20i/eKDqpCjt04Iurv0048x8jANnkHr2WKVJvz
6eT8Q2g2oqTfxxgTyFQQVtcV/pDhh1GQOwKWOdeYm0kTdVYCjj95LsRBJi9toUDA0UM5p+VnC88y
/r8HGEcuYlws6HFL04YmD8gMJ7dDRetv9awDmo1G34dhGGX8pGk1Hfx6PSayanGmN4K66GtV54sg
Ij5+Nv2fFrlgcUztYRRp4dSxjlwPl5N/eBNaBRdhXh8L9mrilPwQZ6BnTe1x5QZ3Iw2sh4jS/uhK
gO9Z1vZnQoC02T/Fm+P/LGA9OvLvjEluQdBkIGVvJQd+jGSubrchGctCKFAStXI01nB56OD7K1+G
cimtXHcRqM1tXGW5KoUsmnEhASrduXC56l5a2JbcISfuns2kYmKWcf2VO/kWcS4Df7po8io4s/n/
9IYDnB3OMVF+ropslVmAshtHARvB8UvxN3NQvHfnJvRZ/tmaTv7rkjpoLQe7xe1wI1x6eASEGicR
ivbNhlEFuPlPKbf0NqCETW+GbiGaonXLlyppBO38z937NB5jDvmxqzhFkQYCiVRRsWYiMQ5sQJjY
xnztYzVydKxq5AjccdnD3H8Gy0sGokveX5uNPN6GUwcXsUkk3RSl8M13JyNVZfNpwJgPtYMBrB0D
MmPKcm6X/YadZF6F+sOKHC3+HIQuQMjcJSeiAaItIE03p5/LdgktwV4+wvGsEIqY1myvkx+pNB4m
yMo4vuHVGl2ER860pnTtuxe5nayds+BvGkYGGeK1mPTpOgMevW+u80ewAadjM0HfAmGgXsmJJT0L
rlsiAeluGTbcU95qiJkLXjuRDqS6MyOSTjcJXrKvzebG/B0va4egs2y84fCXL7UEowPOvhUdXgfa
nNDgW2NAdmYOkCaMHeOj8CfonBDi78wO9DZgrniKbHNZK8T0dNKkAWPQ4gb2o6GKh6iTI4hTwD7e
Yomc7hh21OPo97UZC0WtTu0A9S7LE+HmKhy97VufQxRgfQiVdUOrYHEVUfM6057xKbmlMIn1cXoe
gaMEQKjdCJNlpOYYu/yU2Dt7vI99ZcRxZsUv85TlmVJ8kG70hzd0W1607sFxZNN6eK6QgGI7NyH6
jEGNPD4+fiWWR/oDk68BPcBlUE6zmtBWjH7yfYKY0kvjEypCC7Yjo8/i2MQeY0u1pX2lrVUnOal0
0ijrMCAWi2hqAbGJ+zosYmBQMXH+UQlLh/wG1CeT4j+ozC0gJ1qOcn5EJ7S9kIy3xDPJ4Z16A0AB
hwwCVurbgIHEdmhS6jg/8Kt279HNZpMS/CWj+Ftd69I3zOPhw+KIzgh+TjwG992LDqM0S9uZ+vVx
aBELmjOgtKIlyT9uD6O8i5V8ZNVvl/g8PbPrKYsVKEFBprg7TjuWo6bfU58M5SzYvy1V13kTUz+q
fID2pn76HH8sHKUDPJcoRZAgeeHsrx34jFrLpXt64X2HsQEAljZ5CA7L9Vm1xzVymCk6kCpSSSwv
8cG7WtFVr6/gU5cfgPeYacPGWW/uf6RfaHCEL1W91XT2CZUXkUQPFxsOws1xeamDVY4TAq9+zCmU
hJVRcYzVXzyr7tuwkMIEa3cL64JgzyyU9aDmtF3NbilDDri2cVgAHoHL+2TKWTeiIjsVjMa/FIo8
2zEBw+44jnsl2JMMP0nem/eCANA1C+dmaeVT548tt6gtaSLaqROiTNwK/GvDI0KxhC82L7FjDFwv
z+avwd27SG7LJ6+Jm28KTD03YdnUGBA4WeG6sofzPolvLRIk6KtfIW2oyyOBivBH2FJpU5KhZa5r
ILJd1Qm1Hj0NZ2LIELcdrET+/z8PqFc2EBbCdjA1/kweeDIjE8xqhHzwgQcET7fdPCjQ3A2FiLEd
MQBacYU2LxfDLMaNX3PCNUcfjFgvjyiRZvOf4RbBcEKw9cBTtf3gvPcj1puLvClJjAAVsvQFIlVN
TAhXiDfUQel2tXI7D33YR/jK8DlIqKe2eRbnK7FOuQm11QQOq93AgsJwBtQAOIoxh8kcLvcs1jJA
PSIV8OEWNZQ1qyFSAgzVrpVSm/OSvtDeFwySwCctO5t9zJsRqkoKiH5BGe7gKvfQIGwFEKwhaq9+
T+K5BmHdATpEqNbilPl5JayPQnzZYJQu0rE8UjRkOoSVjaVrWGHWLkLhXAbK7eTuCFthG+rdgGNn
pO2UqmRBSNkcUEh8A3xZcLb0JgZmcbdrKmdwUN84b8IbAG3xO4NQtpEpp2QssjQqiCyK9Vcf4UXX
aj7Ln6zXgeGkNig/zVeeDBJ7FSsKV0xG4cukvD/ipbEslUTWlyvb0F1a+HNmV96kIl+l+x9+WyhI
EZ6S7/kZezXSXqo1nUlMfz+9qmqWUy+gnU8bElmVMT8HdE0nXGnYmBJG0+mdcFH/KBJKG9hPfQ3p
u77TSTRYIrS92JEBiLeLdMTce7aZHv4i99CWU1Soa2WESoe0X6RnUc/KIMHvMNS+VznzZa2lgFtr
3MDzovuZv9gsM3k3Pb/sVwHYfVf7Sgz/URa8gfs+kwhJHFgUvD9G+baJqvEavTAQnU/IacGPnCKE
pM/Qw5B8Z33Aj6uu6PBGa+3asV3bDt27uFMOuc3WON7Ly7yDEIxupZJOkuEI4ok7kPSYYwb6WDwO
zT03j+hDpWnm/EMx4VQEQ+VA4AqBzsw+/vEgbGztdRp/iXoUWdtNw077PeUvDLKwKdWzjiN0Qe4W
/zeXZREjmNf/DotMoZGCao4G/ThbklUDBEdMS2tTRRDKpCaZUouivZ8IeyYbTW3d0RS5WKXiezDA
aQlYw8kpN+7Fpq3GBxi41bkF3NbsJUBFkXJFdHjGasDOQ8UCEzNU767VgLNLubjbho0F+1gWWVho
zA/S9CRJPK/Y9F+aYRGXgIhnmCiQSdoScs4XtYGJkhwU5k4b+K91dBN7n+POG2LTr0eRnKBoAsmu
EYMREmbE4MNIUWbH8ubwX451+1mlF3q2gr5F7IeebjkgLR03d1FGzysxsDuBDfHVfpI/6TZcm4P4
uJ75SI2Qg6CPqPUgPOxIBdNIG+ciHTWs4b81fr7A+ohbP1h6sJFaWerW0bMKbKCDikJN6mI5QJpY
Z4ixRb7e5VZSJd1TvkTApuFe68fLGSM/ZUCb3fBjXm8xobo2cTLxI8BBJbSLV9HeIhSAnZXpgDB+
Zf/k8uXJaQKEcyyZRzLsyYV90pUUIAmAD7LBWS5r4vcNh0mCuOYRfn/n8mba3haYap2amL0z6yED
Lf7BmQRnb2FzOeCa88TlELPklE5gaaVMa48699hATLu5IB2vsC3m1ma5ymQDioICYn6dQiwd5RM+
IuAquwagJ510/Z0QKpB8h5iiu/CpOxG+xAjc6kwV3TuPpofhCCHa9wXhT22JtHufL7Ey+Z4BgZ8A
pWEHCO2S+nUlHgGg7jYtoXnEyI9dlKZhagHmgIx48hDu6WUn7+IjOqEphfMwaS0hX9OfJ28wioBn
TkNypevFcz8E1iMMnir022TOq0IYUHLxytvleV7msjF60J1u9x0GDwV967CtNj5axZNT0G1CoSu8
IaSCCC9E8dXgaCMR0cHGYzQ4EyeOc6VR/XhXvjgR1hfh2QNFyglwn0f8x14wuLaVdEcSHS1YNzCz
30TzfgEBGIr8ZGwUOv2SniwQKyRJjRwcJ+f9bjBPMCbjKUDuC0Zwb8aF6Mtn66cWIEHdJ+RsylP8
rln7XSm1Lggg+m/nurKOtoVeEGLO0j39tvPJY0argNJx5ohDisAaotpHTJAMQtJ+3JERXEqsjO7M
MNcXs2fjpMcPCikLl616TBtUwjGmrATymTSTJExqudvvHox2lm63nRTXHjhLIKXaANGZ8eUmU4Lh
MuGSaVjIHFqcjz+BCDHkN2OJS+WDhx5tFmSxzJ6k72nlSBnndRl47c8xpFh/C4ykdUKUUgWTOdeb
9xOYQXG2wPrQLkV1GpQ2mhR223bw0PsBBsEjH6ZmOH7UXvdqIbZU4YVykMIWY5vR0b7TLjMUWXvM
wi/kmVaUdEHc7Qg8H6QQTJGAqEJAjyUrk/Jlhm6Q1MKgDiJ5uXMQuGA6TTI8inHOKDNfDeos1D1x
Mlq66ZPjjcwo7XF68GXk6Da6pTq3jMSiAd9YmJ28DOVhF+6FutkEVW9MqYtlQ+PxdcMbKmwT9Mcv
bLY4yUnoU8lezEtQyW8l3+vpEsaJ10D9vMulX3nDRW0asyXBRAe0X8I7ojY6gt3JthKvpUDIwfiH
2UMIebmuxBoFduRPPf/EjhqZ4gNuMVi8TlrmFQsGxLSGSvsmj2vImHHtsazY9Y8DHjVqf9+nn3iJ
oyIRN5nPVS9yYbxA7hA7+akdiHVjuhb7NOBekptGU68m/O34zzh15VqCmO8GjLFFSANbpCMHXiba
RS55PplIOqwOQj0Fyp1t1skYw4q6UsWgW4LVP2WYffE3TyXYceFBiiTJxZjHYRuDfuA1x5qCZaXy
m2rZTR7rzP91dty0CRTzaDR8a2T0yXCf2TcrSMb3a0uX/9UxD2SWX2aPvgf7DMHoc5S5xrvfvMjR
fX1I/R+7xe0sz6oqwo3aHZdI/lja+ZphKJuK1SUG+qoZkyySOzAxcyQl0n9GLHI3RBNJjC6D6mu6
tFtTZkPveSxxpxPW0OE11e4Nv+hSbut2topSME0+nGc80NdrZszdj7cI+I1pfm0GN26+vfN4zvS5
8MROoXQsmlIpne85jYrXnbmYfEdd136t5FXlFfFF/dCWEEivQlvb/OgdWMTE53XVV9LqS66LiNhp
eR2WVDGfKu+6mgZOP/88Eo5ebEjjGZTfMZuk3LmpChHRjAJHa1ah+1A1CMswO0vabzWjNfkJ8uGO
boNNj2+SXx/jrxVkhJcm40kNGfA6XNOGzEp+WzZ9Pe5VYBd3qZSa4U7zPLs9/FL4wAcmdbHJMJRC
hwV+DQle/15X5esKSwu7+7wnq7WJzk3ooDANVz5W7DltczOsc9n97jg3m4HTf+1RdUCYM4/GUo2R
U3Gy8FW9DB+qZBXzHYK15qVlI2xnWcrqp7kszObxVOfOUCqumaNnI0uawKWWPjH/2NWaJlHa78kE
XeZbJS9YgrWUwo2e10iOcwJoLGbol5l9mxnz3qu/r2LePC0vRPWGYWNCbchK6/L70DOI4aWSjzpE
3kDEs3fqIzaS96X+tiFT/VoCknxNjAJR0U4OaKfnk01sidJE6GQdEY1pj5Mp2VKxcaXuZTF6LU5H
5KYoFD3knyLV8h1UAMRBfumt/+5++mNffdpmFTPczy+N3lFNGotjOdR7xqN0MCmwqB6UNm2V3tvY
fMcQk3KzfzQ2VHSjPPByAjn3xsojS5M4K/aDhSbTFOIDLGcGB7aUPcCC+gNosVlbzI2O/hQmbGzO
4nl2g9OeqpnJ8gZJrFMq7ok4ozW0dvAzieVzzfwLkYR7LyN/UHQcB5DgrUA6RZviTjmRIQ+0iy6Z
knkplTWGUA8fDX/s5zHlfP3lkiLhcVYmHKiFfGvyKYrY70mG58itDE6Vp9Nl+hWmdKb7u1VtB9wT
ZCz43nFydCzRRLYbhYEa7AX6zB/lnc7+TVcPACSkBpAVZHNqGP1OFVNeAVaRwmf7epcL6+kjGO5r
2ggAMZaS2hFqv+YJo+ZKZjWOsgsT6DUn8ZpUAiIWtBvEAbpknExQ+ZzImOcD/75fK6GAOIph6/dC
LGdL7a2p/2chBgG7SOzEcDvvdYRuRfqijr0conntGySyVjqJu3dRdV25IQBZi02/f+djTyKrj++R
ZOo9lWjthzGQQ1gzKWP22avYLqJr7jAbD/jDy6ZaK0aKH4gqdvtWM0V0Jh35IslXQW8HvMNJ9HzZ
Gb47Db/XDyft2++hU6I/VvYwlyNoPdX1aOM4/C/Rza5C3nOb3IIE+ZN2Jx/7x4z0FrCMxBG0qrxH
zkdfB4S/CwFz8dt+OvmPETLU1ilrIbYihtVnmpiu3kle+f/gsFx9/hc9Q3yz4yM5lqyuTuvnmYVl
+TEqbupHWtbY2e4ra5BANOB/xzO0TQYgUo+1kKbFJWAj/2FMLn0AyHHozFK91m0C7pL37xnolc3k
QK3+uEeoC5dgiQNddxG2UVoNB2yk/rnq3qZDg88Zcp4pMLS5PM2+k+hHcgts9kImz45qkN+3x26G
4qvJ9ndVqnkF1hjNh2fwaIqKbg+dNWSokUfoZdE6f2GsgiAs5pNAsBU4wKDa7i6Y/R4+dXvx2HyL
2S+Ev288chJVMf43uQQV64757Q/9qAFTuwLrKpETDe3iog18unkhI20MFhmRgXXiYis4e2ieExN4
qhCVY5eLhiT1OjYmwKpD0KMiztLIuvUjtw3NuJjuL6GhzdoMbmYjpLV33xko1kFCPrH3nBRLYuH/
WgmZEhd1yfd5BoOJY6epE7CPVB1nrGF+05W+JuKkWG4L8mB8WTJCTG6ordXDIznRPlqrw6xxxmNg
5cuJ5nRwMruBZvWrhUd/ouOLUsuU5NH6tF/O3lmPqsdRjHY/JehJXF8dpf2nXu12viAZWUfk9W5z
YDcy4PqESF39102SkZfq8pv+jZ8Cf1s45D86T4xUBqLeCsFlZJUCqzhzSsIitWpHGqsTkdU2gVNA
ZuXNnxB2c7NuPDNq47eXvWTvhpr137T/WvSd04PBKUAK2RHDIsIxN7pjNgpJUQQvGQTJVjp7Q1NX
lyjvEUAkYQ3SFjyCZlnt40VY2o9igYu2phIVnWmqlQHZqHUKhrOzqFeU4xMHwH5D148eMKAylbZA
B4hMKFYUCAd+lmES8USGgfqGax+I64K4SlCl+mB+nlXw2DibqeP8E3zggkhZfitDpdt8jBnoYilp
wghFHeMnfdDxtYXskSRsj0sMcndwiiH1Zb+CCbNKzm+RreMiE24YuXAKBSNDywUa/rZPNN1Ba6Sd
aFj2ExyzZHQlRscMhQPHuPR5vVblxZWBTkIE+DyWOpN7Ajrrie4Xtvz9VhWIRVLGv+2x0BX+NLIM
R/mdfzLk1aav5+G3TlfQB18J8H+CvtoleofAXIeFDITwQAq/wNieO5ENeLWQVT+ZXnmxO4j3JpGS
Gyv8byj5O0v6/APRDoKIVQRTaD9E1Vk7bNWQAYl29aJr9MBFTKg28RR2Sf7ECzem7ja9gEoKJ0zt
tB9UWtoIbO8klbhYFXU0RJd8CSozVWk4ZoptxpZN21CKpRBmmOIw7A/B58/CyP902E+xUQJennN6
/GqMk82AFZWy8CqpxVStSNemaRc2W8EbCRMehOAinjiaADI0eYR6qbR4XJQLgr6M2TJ8/ELeP9E8
FuVQ+OdX1xQYG7Dg1Gq0Xz/q3RFCWwQOQc8B9IaxX/SzyHl7mhrXRdtxH4zjiBENWndZwcsDhrAj
/yQPMSvdYMSYO+bqwEMrOQVvT3i2+oTuWkLhwoGAlS6lLq+7B0X8SAb0yr+sr1lYbEJOwqjHhNIx
qFjC5ZjUluo8eqkaHofg7tyA4vzxYxkjmfxou8bqDBESiAd7iJnR1oGi+Z6qz3/Ht1kRNqe+ZHGM
PBZMj50koL6/d455qk3SVhX+DTtB1VbHgRl9BT5JHgnAmvPoLRuYvippNcnMqMDD3t+0SlB2v4lg
nCPXAuBksf9alRp/bPkr5bSWTQbm25jGruncUT6bRl96iXq0D5zh+4MG/HU84oRBfBF+Tlcw/VB6
kuqwh9QhUKdeH1KUhsO7UQwIxm++FQpk5Rkcdmwz+mysy0X/m/ZIBOgUoKOS7U5bKHifnV+9CBFb
YHRpV9Bef1cn+GYUn5SPSeZ7HwR6NgWtbzI2X7OZAFdozFekVWXaeoq8h3UvjwFD0HBDxGBmhVK2
jxEMv27PRpg9h++PcM+7pLjOx01KP1L/b9wNuOT/BvyCZ48LQBniLXN5gBu4yqYdxf0o47oHnuqY
qpTEvw8djE5aowZFEbOtXkpA0vHkYQ8FvDf+niEGtmRfHw37+8BZZMlNpIa7Xo8sAs4iOh1pe0uF
FRVM7kNY8Y53EfLoRxLBh2Px3odQQ9fukmeNn0cdj+Or8wS9k7qRaBZFS64+vza7oMBmJan4X5zJ
m+ZhM4ofZFy6gaDS4AYLfJnkVH/9Ivwi265ooEyk1b1eNk3kucIGfFHfnrZP4aN1LI73giygTjjp
qKK0pbkpfFmQsswUdFklsLNf01OP4P2EfRRtawOftO9q4IiwLg4fnTcu/7gyZA+Pw9YmmJyEw0be
RDlvMb2DdtkAFixLO8gr8j40yzCzOTv4apRuj5fnNwLNOOj9p87z1Gzxcfr2RhChFR+0pO3QXSt9
0FwRg3N9i46FSz2k/RkmeARYmxb0MvCzIpj30vvEZ1q5ygSybbLrJIQNFJdMHxh8nyE1KcOPplEH
83NnlYmWMFJokxwrTVbrusXlwOqMD2Xx0BWlqLRTPueJ9+bPySbyMySUNYUE60nSsvnJ6ETtCC5N
RQYxZiizgy7u2pNHiVA8sTi5GykPEUcwYM4JlFm1jc/rBbOFRWck3U6ekMx98uleUCsDh3VMYrch
BgQbMOU6nbO+2FfKRG2PCRZkVpJ8vfaQG6nZLdk2cDdTZAmE8D3PZeiWlNMrojveVY3WPvMIv8lk
XN+D5/C45fx4F0wTLg/YqZjJSe0y3JywO6ef1vnNflfGdIb1gBoGQOOTC4Eqg3MBCW54rjlAD7dC
jHZVWOUp4v/+8XDJZuDUmOkYKIsNHkYDWFY8UF6ns6P+bV/akZWBUmCF8TjWO+759OLSiVMYloTF
lKj0PjxSMMWEwmIP2lInhZQPXRfyN9+S3LWpwCj1zKD63tnau1XOTWyHAJlwwdx/m1aa7Kiez1zV
QHkiN8N6/9f/a7M/7gok4kD9asApHrT/OXY1FQszxmsLPuDPqvgggIvUfizcOmoMb/4/M4cLuxwP
KYuGOJ9cPwMPT+bJlM8bCl58ai4V116b6AI1uZwsq7abvzAQ0KPzqYGn82qxoGOEvWWZuQcxR86+
bfTLxfgXQKnWfnsBwL/7o840rl+LyErRT7ltDcE1/iUpP0t54D0fKeSbup9ILo74NPjHJWiRv2Ml
ZsmkDvAoic4fZFvhgq8TSeL5RObJIFtvnpeTf2QOPLWr904pWx0Qt0e4ddBrQRq9+Gl6JqsV9XcV
VPCiSyUn2MLlwyJuNJWMtVzSQvmGowHapVfchB7hFHZLgQP0Szn0gB+VKVNDZGlkwI2axoH5rPFu
RNDdLvrNWNCzqIjcBDg/gBEuvPJ4D6wnjCz6yg3kjYuzEVGBMv50SwOqn4PdJ0u5DkWnrbP7MHAA
07fvzwInbDfEm71aLx8Wq1araPGHglfyQG8FpxZtjgfPD4cwe/NNwkaKVnA4eSlKKyFrZ/Rqw2RJ
55vEkfEiZoTMYYS55UBPMOISLp0i993z7Osenl+oHZlLmYk/7l+8SKBseyVRaD9mu7vKQdNLO4O/
a4AHLhzmD8cMnZJ+JrCaCJBH0IMluuC8k8OyNHJOga6Xa6relOq8uBLx0XOrpO145T/gWuLzFLlJ
JklY8+ScIysi/tgD0/o6JemhbL6ngTrjtudU99l4KTMGE6KFqCmMF1KuzgFhtS5POyfk4UBZzBcY
bfZ0kmcOlmIN2WlmdeK8MbdBZEPGRhwoMw6lkrs5BcZeGFqUBQDRrRsbjyqb1U+KnujtR6BcpVBW
dilCmNDvuij7csS3psuUU0M6WAkau05hnhrMWCVKvlACjJNvzK86n1NnTYQN489ChmxVyk0Z/YRd
9jnJHluEUUlYoX24KyX0y2Old/mMlW6w+WGh6IbF7/PyhPKCnOX5JaU9bF+E0fjMLp80Fs5gVWpF
BD09MXsOHQ+RG2cUEUJIluMWa1mv+3w+1zg2bkeYWr7MGfqvRUhsJk5BrE4erWVlveX1w6MBZsvJ
7XF7QSutDNi6YFFmhxFDQ0QdNvD1ALSPD4pR1KSjVf8nyEixzZCI0w10yS7KwqsvDrJGWPLQvbhl
NKymohboHFVuOQi2vXE3nL11aJ5QW9fTcuJE7g8cCm6tR6xx7JRtZ9Evr1T2yd3idRMn+vGsL4ig
PWE+MneXxnvuo4EPTJ17XuBrtqlnsGspHGD+3cHjHcW2scUTCgUeMgabqJfYRggc9zOe15Y9QzvU
w5ptDT/lytnDYejpsnNrsHA9SLgWuXpnB1NdR5YTUBqMgH30yN2do2EUwDuMzMGupxoX+0vFSdkY
3on3cea7XNYms4KJdW+Vm+mXp4PcqXVq3Y3AGIUl8FUTIvdK5z5tNuUXZMupZIrwtsn7TTMrQI4p
ZMqNc60Crv/UH9vGKcMxlmst4htNtrIC5mDgJimqhFY90T9WVD4uZPs+aZwzzpMtQhuZIS3fz1Lc
B6RaZFbc1NyAvM7/4PAFagd3m3hVjvXp4l+UdnEywqCVkY3VZ619PGuu2fI6scCMP72XplEz+SAB
smUPkVIA1mwrAbWqpZoexhvPMkooTtkMMZjUHdtbY1FfthDFQG6PSp++4iqhXck2ckHgXqWtxH1d
VUCSvoN9fagh7g9KG84Fz1X10l735MDVa3C1EsXb3KB6Cnjp6muu/VanqiE7b+6TSbrA1Qg7ETuf
xenCe8b6i2KD++zV9xSYUvDhIYCg2cHKIV1O1HAxWi8e+M3P+R9DV2Qn2RtV9Rc5pRIumGxJ9+lF
RCMl4EX1ROuMc1p5o3TH0tAUlNLSza8xYF1XYx0pjbdcY/lsFQUp7Os3kM50zWAAqTVGvAe/feSv
SREo4BbEwpKQeAMsxfD8XgfxSOqYwxTMTMhD1xsDwvswh5A+rBAebpqZ0Z6CDH/lzVXwuv+Qr5pR
UUkLSCBe1Ulhi232XDOXEbqRYJCC2gE2rYoBNZNAC8fSxXDxRfvge0/rGUniJTrCOF3stZY/7Cr/
PLM7JEuc8+Dx+HzFfVuhgtdhrtM+cSKcBE1anTw1901GyUDlXkjcnW1TP99loVazp0YZN37/cDBl
9gr8c+s4P+ZGqUcnpk7WBJyKbyNly90EKzB1i9CCAvtxEdzM+sbr1qAdWs3tPc2ttaak/80GT+yY
Ap8ixPPkJNvV/0lg6WLnz/s+XmQa+0Xs6lJpVfWUevg3raBcHDgoXs4pYDZRbnbLXJyze5hXAAkc
zHathSs5JwucI41ThKWBlZOSiGgzvlGSidvyeJb632U40HvaWbsARLMCG8ZSs/dHWwLPj1CuC/eW
kJBVgfOokxG7Xogyaej2Dj03o6WD4q6r2HaCOUFCSXb/mLw2nJ6MTFKWmDhLgQyunrvUwC/JSDjZ
n/LPDAKWV5SiBMIBERPt7GlntewGqZB0JKFdpuEFyqTrxYc/e4QvVBVTi8uMDVt+Rs6NsRw8ORtb
iy8yJVBxnCIEkeU4XwPIApXxIannBa1Vm1C40OKJ5z4Uj4+FvpUPGvxvXmtUY5UWoh6QPKXTXpnj
0BDHLmQUtC1oPdChrDKURA+po88ztfiESbnGD7AWMcMgSKXvE4uNNp21BH+3hFIu+Hxe/H2nOqSG
uqwVpObfaTaqJSTe8KM7yYRdeoQTQWkBxw7g/jjFbKbdr+IkOWxYALfVY74xhYyP0iGM6uVNJycw
HVN5rO9pNoGhgFUAzwd1D/cJyo+XIbnswJ0sk/3Rr9zfwn3DNTg5Du7YclhICxwBOj8WabfrHiQR
YCO4y6t3eSE+m3ZgD7hGj2+Rn9HKNs8d34irWGHtYCAxTK72L+dCEOltPvcjFOIZLvOXUzoTMKwR
lV/sGv9gndLjMgJK0zPYFod59sU3QuI3a2EHSfW6+So2jQp2I5n4iS6bhScfjMj8dFzFj0iPVHjD
FMw0ElYhjpjU8rSakyMvAztwPHRxrg1qZfuK1gZFHLg8uFa4j8tMc9BB1Gnk4Lj73IBCvVRcnKlh
ezUHoLQogle3BxZPPuXQ2Ie7UId4vgbiKLvt/dV+r/bpiW5JeLEIa4ci3XipWDvsqvXbFb7qWc0j
26hNNtlVR/aKFqWW8xVQHtsuTzQJngVnWYKuszgyYmAt+Yxs2w1yLKpbALsAVhzW1Bdrst3jeWl0
lpl88TmJSNzIIYP0VhY9eQuJCvmFZvxh+UqTYnCMl8TeOWCc4x0+JkH2HACn/Fmdfm1SsCN4StzU
lAPU823HWpJKmobc+5WHh4DyUhFf9sbGs6kffostCfyXPOAxw5xwF5biqg26YUW8cbaUpF+Agjuz
j2XwqZWtsWAIaOUQR9LkU3BUP7WfkC7JFNHm3reC1O6moKzyITDFKjL+b4El8TCTq8jEm40pclNz
neVdH/Mn8yNDNBHbk0Tinr0N6tyJ2NyUTSA5VdoHQqBWUF3I6FJ2gjCgj3z2A7H0jxZTb1z4DGy9
5IeVp20ohc0WxD98yzIdx+tVp0F3Hf69o9oKWlZE44mdy+5skhdc6M4vRKMh0aIQU5T0Dh6J+DmV
+VJE4qOTymWRG4mYEURr1yVP+gldbngUjT6kuf2UjQ/f6Dbfyg4wnYPsynfThptb/v3TRu3eRJM7
7YqKglFwQiQ9V2FbeKffqwTCOJjihaAMrF6SyiVvIlSUQDQXWAQK+ER7PQhulqPxu9TZiTIKntBN
VhmvTMIPPhlBogvDU5Mh49gtuM919enTz/DcDbyeCo5DofYUmDJFBBHouUBNyabJTUJwJIoNRFhI
HDDDnW1+swiIQbOjdKgPbRKNB7Vmz9jCnMUGz7kK+WKFbAst4ih+kiLri8BkWLc+PZMtsxeJTFUQ
LkKQ+ugdNCkho2+14gFPC39W7di8ZFCQMzcZDfcAJeBdaZNffDfsb0ODVFRTdGWJTiqfxo/k+zkA
6V3BOoPkDKT6myGhjqImYThdqmWJYr1YixpqZKK+XUwNHc7nrWSsMrq4VA8v6Ps6V0RagN0u/Y3+
IFhOBPOc9VW5nGSmp8w9EXPIvHxrUem7f9PWb/qoCsCf31mqio7tt3w9rHTpxhKrMawxsCI5415M
GQ1Hh73l1EawFFJVnMeAuAYljlqP10VmYLne302jrO8D0Yy2fejv341x2PBPxrYNfyNLlepJGF9E
9b6fzjurBhBSuvtbC2i17va3gaNN57DzqeVPwWuhr0W6KG9E3BJ2rd826+M9riC4DuRZNwjGtCZy
qIs2io9A0yftdzVF3MiiR7WPvmFBKk5r7rC12Kj7BPxO3cVdZdx5LAGweY1sxO+7jAohrD6LJJqO
NBfxIazUDN6b6tNedTcUFmdpdjbMJaGWzkNTw6lhxaq/zdsABUY+LZn/ix23UnPlp9EVRxxPDqKq
lWnBsVE6r0CvtZ7iri20yaF7rXqP55vEjjY7eYAxazWrhe72cxTEeY7JUAJ/SsJaolCDvnb2ooG+
t7bU2s2SfpZNLaguEVYYKvDHBQS7flUopYUOPsf9V7lW6cwAIkwS/6Btr3F1qArnlo/62U1deSHg
v6WMc9rwHQEiTWwSassfDplno7ShwR2O18i87CmJfNHzf4K+eKe+MF2s3PHuNCUHcu7yVfbrdVG+
oSJuSWnUnTBnYKYlOrQ+wFvriqAJexQMRa7hQfQ28yvbVKmj51tDDx5jbIfWOh2qpO9zX0Px4Igu
ZnurF/yx3Fgs1RYU1YSwyjl/sGBYb/tpiq9hZldnEzAj+qzJbCSRBwBDZNXBXXQxkaNmuoz8lZQj
7eLB4ctYPakbbp97o7P4qo11PR0Hsa4STF6kn+pXcLred9DXH2ZrO9wtt40IAE3jM4zU6PJlRqQq
XnWpXhJCcWUePrWu+3QdMcXQZEQ2r/W/NoysEYJnq/qBhBGoc3MmJjJ0q8hztc/NEHomlbzHJwH4
Afq3xTc2oHxzZVhqbJnAgboG3ysfPMS4/8bOXxsqQ6+pXnxwkXrfBRY+1apWeNbSjL0mYWd5AiP5
5W9+MAb6ejiCFtdUTmd9Id/onJHQRJ0tAnKMs13wlINbkvLPC06pdnYr48x9D1XZDOjdPTaVXOXc
Lw8m1cOa15pkvTlb/tiy/V/2pBSbQsjGIceUCY0I3BR44R9E0M4JWjpEHixXVmCaV67o/LtP4eXe
RWkMDO03wIsM/HDqq7U9j7Zf1hiJyl2q7JTBuUbmBiwZ11wWcTSC0a7UqIxC4Nju5dRPNSxdk7t9
Rp9PaZld1looBhTZLSB1hO1YLehBGxFfXU9HmUPGYx+EgBAXUscLL6/C2MIc+bxfqsuh+Rsze5bT
LWKCiFfN6+LwKmIr+WXMncDMmhA6LL/7dXKPVe16xYES7i02WyMZ2ykSnz4LiISFyHWrh3+48pID
ZBHB3+PKzIMNR3yrqfJ8od8gSJ68W8DwChF0BL5N35hAyFto+xK3GgO2zqu+MDeMscDxfTsDmP5M
WJUfFs03b1aSvHxZadR6xpmll8q2WhdFLuAvF+vmpW5S2+6nUzYKi4Nbp2GeTzhsHd4ikKSIZt8j
QYG0b9iRFalAqefK9aTw3tcUFx3kmn86hD5uMD1DFoioTYx8qvpC62Kunx2R2NsRzClcXqKYVyos
CGAtVJafTBrrjp01vxIJLBg5G+3QIlyXurlV7PuY2r67bkFOc+pZXfttT+D+corFI+U1N+OfNO0s
J6/Aj8/FbZ3IPhwQAe9bt+q5A07gny/fmTkAH/u4z2HgoFJbo75FRol+J0UllMNaa4AYP8bI/rlG
LCM0AT7KSfqYMfCsy8t7fvTArzJUrw/FdiOGlLkaPskAvN2WFZOBpyDFoTvgniY1coaL/W1KzlPT
C/xXblTmPlkJ3b33WvhYrjx1D9F8+033U6XyRzfqGtwlUKzLEnctlk7/FwVH062ljPA5IBx3b8Ok
06R8CpgMcdoU16zMOf7yjfeXv68rzdzWmsb56hknP0pATqgRuVZKaCAaCeKWLQ++u1IPHUbywKd8
RDHaMENquvh/TtAk3hkuPoGplJV/0CIdL7l8dGeZkndsvfF2yr4fkNfjA8fewFFdzAS+nkb5Ip7Z
4jp6O6sfUXEVxH/yTTh7FjY1XBXUDl4/ENFKzwygpT1UJyHWnF17Z4q6qAY3emXXj2T8VDShCJs0
v6zXMnMW9wvYf5ZddRWnzNXgt3eXcW4yuxziDNTysBNOFqghGcyLxSm/DLbX1zWejVUaSeo/yKj0
jLNw/lnLajc94kTyw07EmUBKI0q8bGT26VArlJniJ7C4ryfLEROXgxVY1pwdKIsQkQVPIeZ7Mb2D
0aMY5Il+Ce6HPQPNlYSEzuyxQjuELbHcZlg/+OMkGgD38trtmgHAQ+OPgyqVTPgHZMdC5SEPvfZ9
6whgfN/SyWJdYW6OViFGzU158Uzrb+VPnt+iEMKF79eH8Ya3Lq+oO1yUfRwiK26EhHgGgck7LwbN
TvKhRACKwZSDrZU+RcdCOdvlXAEqZV0y86sEQzxF9d2/pdL2MKitefMxMjwMYUrQkj3RyT3gQvh7
MNHlMwyBmQfQbcKS1sAhtjWcHHhh8xi1NeE153uzWQTOJ1LteyPeiO95wJEUolvL3D3a3FC/vEPd
Y11qiW3CL2YEfufDpg4AEVJpCfmyCPip+zlPIDYvp3o9CuUsYVj5T9GUHmimdLpMrge5lvjIAJ2h
Yiz/h9PPsjK7oPRbEt0RmNMpXmCMDVRlwwFgkHWwsNkNCr8Ks41WJvM5VyDI03+8HwhbUBkndV3k
wwiYCT/3B+nWMvS8KcAG83GxOdRMmwjbyvqHHuJyqnJK/nMkEPGi/QIl4BEKdFY9
`protect end_protected
