`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
dlnK0IJK3QgRDFdrEBcTOPzxDfGVk4BB1Pk6oOzt0z2aZJmhgW8uvUf3E1hKWU4G9fKojBIvuj8I
Gl2KasV3fg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
bWdqgHDyHTwDxcaDjfg4EaPj2r4MU1PcPzBsf8E1I1w+Cv7WJ0j4hTfUoDIaFWurQ4t/2VZHWyZs
olS4rDrMujanL91QLTmsJRfCXED50Ljeq66Mmp0rz6r1Kkr5hgxef3BhQI3ZQZ2/DghM5hvpip/E
wRG/1buWbc3Z8VfE0D4=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
XV6lpMqdYehAsK41LL9E8lv83ma0J9oMf98zlfOjZIi8QvWgFHrpPe15L1Klq6RCDSlgLJlWOnRp
1+MNafPwlgkeKoeKlqcpn7h3kF6sduZXVK/PAPYN4C29YsYSI7EFhC7glJEA4Lk+4PYVCPpmOHHF
AZ587E+XiqoG0BCwfKqP5lsfBafpIdNci1mw7FZO2qGFykd0OUM4XH0+A80GA5PG0yHbZxwJzRCW
oGzQd9+6yfctb57cO/b5Se8icOPGrb7wiSEpRXLimxWzqhJYBwIO6ZEJbwdvMpRHgwl0PUIR4kcM
5Cezz7ckm4uoFydCgcFT+N9ggz3mzLsApwOZ/Q==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
TTgJpXEFykuTTrcOH0tYDSJBDR48mSIPN+ED2qe0Q6gnmaLL9AD+WdCcKnYiFI2anrCvh4GWwf25
vqaf67paDmZ7Hjomu5kUr9CWvzUttD8TKeHvUoqKJqf9uwrQZ7f1bP80l8Hl45l0K6UJmuyS+vbz
gInCm4rgaBYxVCVx5Vo=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
NewOtClYb18ngXhSXwCXpgvYitnFNVX0yF+ZO9gn6DGBKYWHgnbTHPJ5iGJ+0PFvPNYGucYx5br9
cO7i81Hu/zlUUxyxRpu4kL1nK+4IJAGf/RZEfhhsBy3yL9DMqrI8rkh6tOHIuswgHEn/crSyXjOy
9CVBjBTKydPYdjUnqzkHFi1pQ3h1fiUSV9LOT8hMAkes30gGWBbg/g3Yj73AulkVnvVg3vknkzlz
ahZgQblc44TPvGBAGIRgeB7sC4q/RCV/m53KGHTe+EkK3q3PdZlxq4Uaja5ZTaqN8C76/dj1dP12
aLWREY5z9MtJrADvbLoBgmJsh1qY4eN4T29IxA==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
GVRegYYsxLi7caNL0HcXs+//tU2Mnd/bOF84nxPikM38TYfKleJ7dsGIc3Cc4hQfeIsG+mCjTm+V
nQHeuGbH+8z2UuvGkhBgc9xZXdUAwZ8N2p6PuqWvokeFB1LbBfWlEVZnWyAFK+xeCwr4feRvSARI
ByaokX19jq5hIiqtdGLh2T0iYgmWr6J5j2H0r8F5rQf59sW09/DopDPKSZILm//I7o1EtnjSvOWq
5SL7qd569gMWwzMt2nyWfxmAB/OMPpxCYk4KI+8hc9wVitr4BR6lz1BpJyKeNeejzHUHlj93IfpV
dKU/KAdpGqx+SFtOl5evynWuWB6DlWkH1QYzbg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4784)
`protect data_block
2485/cuSVk1XFaPrmRWYxIafB9Ybd+zYtZ4OwPzoO/Ajw9kkcIUP1QAEe2HLvn6tz3JEvMUp3KVR
4vhD9WTlSt/egtis6xTCQk8cZmcVUzI/7hQwaxQBLf+9Zv7N6B6I1RpywX07js+BBnTSatDgydYZ
4t/oV9RDkIp0PFLbOpcvsIy5LVT5MUcaBMy3xmMjuBRD68VaPNUeoOrKEryrscez1NadB3GMMjjH
CzOEMu5EELDae9IaKOwNgX0KZtKY495jDsS2dvkobXJTpgW5lXwM8ANJRc6+q3opwUIYzdjv4B8u
8Ph1SfMrybFQLz8Yuq2LnHabIpDkfL3KA6EOfqbXsU/M3LvEFoQVeGS/gz1LrNg/+MO/7mGZcsmI
bF0ahttX1xAmBPWrZVD8iHXcwl5WjWv5+SsrLQiOnuclx5+SUGqWMHruw+cXXHsz7gBZfC23CnqC
9DMxwixMhDbBGk5FanJPvVxcKesnPpeu9vzLb7vUr4Ui4z/jLyikhRv9JmICaIexhNNCQV+PxFy1
WMiOpX3aU3Z4Jm1yhbNqqAXdsXwP3xfaFZc6Lt4Hi5BqJhMohDZrfSqTwfJl/I0rNGA6BG8ndPLM
IDiZ+T+HuxF67SVcp223p2QYl/fFtodcTfKUdGIbDwMtY3nenvn6YRMn1RqMTUVe6tRP5cPcAjOC
Vz8F6HhyjKI45xl1vuHPdSsdDCvLBQ5C/CRXOdqvcukLWYid6TDztmmw1OBOPzYWOQb/YpEabBTc
tctlAVHTZEbKBzwPUQEVpcA/vRMG4ddcNnAgz2VquAFi89HmksXBj+raC0cWAsks6677cJBl/E0G
xhsmweSkiQXFk/YdQersYGbIA8mmSiAriqzk/Afu9hEGXmJWPImsGC4B2F+n0NTG5RvRCrRdXGXW
ZtGWX3Hcq3bB/Za4Sh+x0oN/8h/zIJb2axtOfLKrEiaR0QLzdr85NjZ5MyQuNxPXyDkXXJQ/Gegk
hC83AmkI+s9aEDXyYE7kdmzBtG/WBohCYNAHiNH65Vk584IssKDJnJ5UOt6h5oZoKqe6eZpWabsS
XoWQT7wN6vLPzQpEjL64qzMo+o2ZoqvG0GjQFlnYCUXC2NL3G/FB0TKkrG87p8LPmjO+gYbe7FCg
TDBErq+4w2pu+yl9/jptYKRXLbg6q6K6CufPBPynmqSo88kdn5lHHDsFlFDKikEcge9Svg2lpomi
AhD/yhzUphBKhTqnTkJEPBTTkcUuhVGDjRt/SsV1bX55awPwggcDbUQp5EVDps6q+TKupwx7aB/g
OYpdGcqOXzMOMuhNm8r+g238dpvSRW/RKuJIkbk6DRsaz6s9lUrNsiSNfSYoVDJUigK2uouIyNZ6
5yTQwmxIGkvCEzXh5V3/r88vGS6F+MrABB7OPwP0QBfzaycSVfJBknm5C0SbM6tmEBB7BIAU4DSR
LW+xJFoZHDq2JvusXUALX2+gpNChgwjUo7lK8DmVeL+FLK8gymMzk8vU5n2ier6sN9H7c2hWcHxm
+VpwL35U3bzpzDDzHbizH+JgklqQtYWKh8uJK7DUnS0ae3o2MY2CYw/yrPQRiuNyd0/R8LZbfyRC
4UTAhBI1TkNFIrIHCV50Jdhi/RUfuMniNOxsDShgB3Oc+um+eLi3iDlonYT2OYB8Ge6dCQaImvz+
ie3/Wnw9yvmH0kbC2WHtupLhDpjZEf+tPLDYZlW1OlQUEd3SYdNmG2buYrbo/xUoAr/zD0MyHY9w
M7ouEg8hbRY7YDd0SSTFGW3hPjul/xW6gH/BUozJ15lCTcVwpICx9ouSR6X05cpg9cw//PyPwuSF
OdBHd4VXilwuCee9oZEaabnmLG2RorjGmy3HTvKZ1BEsMtbZdwK0rEQGcFMX/Sv3S1u5jCau3Lym
e8R/RmISJjf1qU38urv6qbHbEslUlpr0X1OIJpUoDirzkPghvFwiE6mLhGaV+0f97iybODOGdzU5
KKuG2K6+abiUm+PEj/vLdAiAQEEmNxUHfD6AtghiNg3vkzv1LbfHdDBTazN0bYQUkHadW9JTfWU1
HHtWFHXurt9aea0lBzB5xRsoqUzd1jfIzXCwxSoZUM9qdVwMQhWPjG6IN8kunOpNiRswKxKb9z1D
arbwbxl2ELkW8q/rk0w6pNhQ6xPbFhADYs409G7Ym+7Jii2V+iw7wx/xoVXY0EbRPrKDQVlBj/5j
JFPCO/yu3jW1a7EGYIKV6NNDsCAKMCqoYiyqkpbX30KgdJn2Q96b2dIvqKmvs+UuEBdW87AQPGpg
airhwExlF6Z9qZj0tQJ6bRNZ/7UyFDDiGRTm9PVu5No9WJhPNJRHsEwgQoYXrOlK0lTh/GqGq6Dn
Mc4uNtCJ8glTbAs/7R1Dv7sJEjVA3aN6NmmfTJMRz4G2LZyDWXWcqzpZ+IVo+n+Kre44mWmC3EV9
mXtnxkSDLc5myWDTMJIAntrQXZS5jqKDchlb4c5J3dpvHuXbV6+YiVmiVRWqqBNZGQ8e6XT6GJRo
PULj6fCV7OW48HbQJJz57lTub/afljpSNAgwYJ+5FtYOyZQj00cu3b05/+sEEYWXQ+UsYWvaHB3f
RSM4aF2RzgTc/s4x9VGZo0N5xA+LgdAWiakHL01GxZVegPe2iGFcxV/Hdl+kIng8UE+IC8tiqmhO
hw35oPWqKwYQtCqRBGbr/nbzLcGZAKhXOTf7VS4y1EJmW8NbBP0z7MJNkGXF/p+cL1jGeAcwwcJu
jKuP/spgpZwnr5A799EOznRLUnrIC6BkgGDYE+LpI02HQTXLDiH6/2sixNDNH9jxc8akpvu+0gcR
o/hjsuuLGHk2Z67oV7Aj5Xg4PN2ygvLiE7ZM/kjD+sexwDgfYuSnX5HXVJ1GAaluOJE+5WlSO1vY
P3SLfhruwO5SRB1MgvSFVqqP94FP1f1cgcQkZhEZQSgWbXAJgfwfmQNej5VrZ3yBYmFAlMvtzhAO
wAwgFAJBcAe7oOgY7YlCOKwXbLIedRPLiS7/Iefmr90OPgKfYibhVvg9UsULR0IMo6YBZHfOznHb
nRLfF5mowuyxmDOOaFWbQBDTKucqW7FL2Fl9lMrNB7lqPEYPd4WqJSd7uB44lZWREj6wJ0/zQgYT
AU1cfJwDXoznVISfEDDy89QaKwaiI/oqnGovu+bgCSiFiSWQE/V3CmyxhmQHrcPyKUOQYIuzLa6Z
fqwuw/Y+T0v2KCMvwDzw25A8nf7fuXNo/lOX7fTlzUFODzCfL67211KPQmxsZkWES1UDvhhzfTIi
7UJ2RmWcSwyzjrUp1EtIAqMK51yiuAoy+JP4+LkqkQczDGv/f4KXfXY1jKtX+TYLDwBPow5scSbg
HcnKrt7UAW0RcubjCuIIo8M9sTvGOGnFAzVY4HrihhNGMNKcH1cds2eZVWOIg9jdac93zklNocTy
fMXYJyfC0iVjWcKojt0mkQ8jotwKB9AgczvXcCmCIJwMfgLfMM7wF7iFvThhvq8OVZR/FBav6pFH
VmscQOHWe2+ShXMp6++ecm9esy8GfNEbXsABRizziHgljDrMxaX+9TmXDh1sTqs3N/55hSQnDlF4
97tIdpEWDnUZci2n2fk8mvMga1UPe0G5ZkrYiUF2DdVP94SaC4qnHmd/U4UtiZhkkjvJFm+D5x++
6duiwR/xwc7XhPQXZHcXuYzBU58ueyMtZdA30/DbRHhM6vu1Z6FkY5Ur8gX+Md6rd4MPICt6Yk88
ewsTbnmdcgYn6PPu3hBSh6I7hpQA0ia9Qx/9G1YdtTxUWsH7FfFMgVbeTLEZmxeJ0Hwsbu4yyuyP
AE3fr3DszdCF791fRopnY+1QjJgcsSSExR3Wfoj2HU18jvnb5lqWNQYD2pE+yXPpRwhhCMiqDZvZ
Y0tGNBwE+TyWjokj6bPH9HbCX4LL1yJc1swqGOlw4JsnSEddAcQnjXE5Gysdv2632HnkM7uj0bKO
YQDmDFb6L4S3hld6Av8wRk/AUS659C1k2wRmMXgxpm9NvEcCD9PgkC9gBmIF8mAcj27euh54KqKR
2TmjOHdgZ4H8xUdNSzIVTRRx+ACQYJNuGh+3sUIRS446XLMCJC5DEmMoPUKfGbNQKWw/12mzV+LC
jwhz3YamMDPT0EmV20pnszIR7zsLB3GEJcUuYyIh4HUHKCl1awh/lGpW0VPQoCl0p3HYFSjJSYVP
+HoJ3sP3QNODn0GqIm8C89JsVRytLGOhitB8FlPD9e816bs5P7BugJpBKemVumRP+HRoaJ7UqvFp
Fb3V/iVvH6DQp/t1LJEGn4Ar5dIuJNaBISfgYqBPJDCxpt18KW2Aue9SfvyOwlYEIJuKdyKnJ7Az
bRlxeFKWNgVIDnGGof0bgOcWQwUEOM8XKHT1kc+GvrWwkqeA4JtwZ/vFcRrTwKZ6bw1A5shp4w7p
Q9BcJaA5vXCMlxQmeqHdLRYtAkQ/ZViInKtcaxNsTDPWhza8gzGs1hU81ODS4V3gtUAACVJ7rJFK
a6vFcPOiHz0jVF7mO6FjCWaJkmwECs2Wmu46+VXg489xyu4MEu+YpKWv4TAoXGOI1FoksZpagzgm
Ny/9mFOJFpq8DzXoiIGIOwBmHWfzLbxNqBO8RJhkkauSr1/vmHbAm2D40C60FvMaVicPK++nzkWn
kIC4p1RJytXksUSNPo046J9ntDH+8WF5FL3cpGk18RsnEG1zqXxPr0FDRWVMbxZ00drk0KazhTWK
M8RUzm+5Y28nS0M6eVlXjJvF8ls9tpwi6uUdHqmFu/2oglqKAbgIPvWMgK6e6o984RhSc3itoLCi
IlHnrW0JBo2G3y5AiWcI64OT6gCufHsAmfzq6bvQHqX/nNT12uTkzruvZQt/VBlHipa62rTFBCmh
teoCH8+XbufVOfX4ryOqbR++0cejbHDCWvYxPrwyBCi4P+QytF2IHgYWFiAyLjLs8wx60KKutM6K
wwZ7SmYXymbzNCPnUMTjHMHGE7AUNn4vIeFPFLbg0e9T+3bLGqtFfypWsMgcTEcTcX94KyHxo7na
wgmBvGDQ+jme4CzD56tA/dyKHIxkYPh3ZME/E73zitt9K/qQrLx+QzmGrU1p3ddCdANo2w3QwHyh
HqRCdsAOWL+8Lt9Op39UGidi7F9qHDwEutoupK+BEJ7tVSdwX8fGagxVxp7e7vbVBlRPNVCj5W71
aJ5+7eNs7MeSpZXaEMZ5B4tdbj0lujawhJ1a6sJi9wm/s0juYkvQx158xQ6jCG13b46XpebJQJyW
Ig1s16UJVzpwiI9KV9eoTk3yQrO36MoVQdOLlpsvFe9p48o2/AOeA3MYw/4k8qnlF1gDik9pcVS5
+BWxYhQKsm9y7Sp2kFTnPWHwEHAw5NWqRuI44OGHfRDxbhEqD2gW8V3by7nbbApPrJtl5BLAo4CA
vXxgjF3ok6jEf/eDZPKMmAVn1tT3BbDj+mdqKR++LjvAhWSAVw5trSYafo939LHOeeMXbh+DAeSF
+NDaC88kgW3QcQ8fXhvPz1dO3CsjhK9Hejlzd5WOWKwscLsohrrpBPxz1FwtSTZZA6k8AG3ltFiu
QIyviOpnue/gVvs4hPVFk8pIOnYA917is65vVh2rYWwj8LrMRV/8RktuFwOc3HBdSHuGsydN/L+h
rAiWcIndZGgoWG9sQ/atEACovWmyuUWCPhTNj6KBjCwwVEMzKe+KQrd5VWh7jy/lCzpOmot8EmWO
b9g0GCp9uAVs1k0JmTvZ5LeiP//g7DnZyrLariexDKSxaGBFTKArZYrAI4XjdFDQVQhoR9ORTD+6
o8ZnrVcMa2++DreN7fCdpY4493L2fatI0VbnUO3D7uVfjBBw8dKRCNYEcn3BFWdoIN/J38RfHr2d
QPp2zvcqeqT3WiG6UOMJl0wNAY2FdhyrRty1IDC2kysxGHclRkxrCKBneiH6bFjmMQ9n4nIKZ5ZZ
8TdKbiYFySbWP6Gnq9i53b2+my5fKHdVwfT/GW2m6QlL81y2keN7E98bryC53ZFiZLsJPPip+LFd
LBKnKgGBXPh4ScN/jC3d/BO2hSnO1sIx5DSad1sll2T8yrt6w1llkwwPrRKZj0qNEjtFYS6bHih1
3FV1il3QLn8CslVLYdZlP4ZlUyINVTJA/6JsZgv3fASJpzm6E1/Oa+nBQ1dNS5C2Ct/NWh+Yr2Gq
jHbbIH6MrpuZA8l8XpUwSmKCmB0eCzCazMOKzTkLWmYTo7rRzj0G35x93YKD7wDpoxMmzIFGuRl+
bXMokgVqulPFi3dpIKd50grAgWHhFj58n3nr+PvjCaHm+Wc5OyZVnvB8EwP+RtZ1DT4wpx/FFZtA
YzMh9B+8C1q1WoDYOUnNwDcH032cNG8/8dARsra7lkpNtWWpJb+yjmTshrN+12DWdWXaQ5E=
`protect end_protected
