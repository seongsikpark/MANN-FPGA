`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
dlnK0IJK3QgRDFdrEBcTOPzxDfGVk4BB1Pk6oOzt0z2aZJmhgW8uvUf3E1hKWU4G9fKojBIvuj8I
Gl2KasV3fg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
bWdqgHDyHTwDxcaDjfg4EaPj2r4MU1PcPzBsf8E1I1w+Cv7WJ0j4hTfUoDIaFWurQ4t/2VZHWyZs
olS4rDrMujanL91QLTmsJRfCXED50Ljeq66Mmp0rz6r1Kkr5hgxef3BhQI3ZQZ2/DghM5hvpip/E
wRG/1buWbc3Z8VfE0D4=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
XV6lpMqdYehAsK41LL9E8lv83ma0J9oMf98zlfOjZIi8QvWgFHrpPe15L1Klq6RCDSlgLJlWOnRp
1+MNafPwlgkeKoeKlqcpn7h3kF6sduZXVK/PAPYN4C29YsYSI7EFhC7glJEA4Lk+4PYVCPpmOHHF
AZ587E+XiqoG0BCwfKqP5lsfBafpIdNci1mw7FZO2qGFykd0OUM4XH0+A80GA5PG0yHbZxwJzRCW
oGzQd9+6yfctb57cO/b5Se8icOPGrb7wiSEpRXLimxWzqhJYBwIO6ZEJbwdvMpRHgwl0PUIR4kcM
5Cezz7ckm4uoFydCgcFT+N9ggz3mzLsApwOZ/Q==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
TTgJpXEFykuTTrcOH0tYDSJBDR48mSIPN+ED2qe0Q6gnmaLL9AD+WdCcKnYiFI2anrCvh4GWwf25
vqaf67paDmZ7Hjomu5kUr9CWvzUttD8TKeHvUoqKJqf9uwrQZ7f1bP80l8Hl45l0K6UJmuyS+vbz
gInCm4rgaBYxVCVx5Vo=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
NewOtClYb18ngXhSXwCXpgvYitnFNVX0yF+ZO9gn6DGBKYWHgnbTHPJ5iGJ+0PFvPNYGucYx5br9
cO7i81Hu/zlUUxyxRpu4kL1nK+4IJAGf/RZEfhhsBy3yL9DMqrI8rkh6tOHIuswgHEn/crSyXjOy
9CVBjBTKydPYdjUnqzkHFi1pQ3h1fiUSV9LOT8hMAkes30gGWBbg/g3Yj73AulkVnvVg3vknkzlz
ahZgQblc44TPvGBAGIRgeB7sC4q/RCV/m53KGHTe+EkK3q3PdZlxq4Uaja5ZTaqN8C76/dj1dP12
aLWREY5z9MtJrADvbLoBgmJsh1qY4eN4T29IxA==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
GVRegYYsxLi7caNL0HcXs+//tU2Mnd/bOF84nxPikM38TYfKleJ7dsGIc3Cc4hQfeIsG+mCjTm+V
nQHeuGbH+8z2UuvGkhBgc9xZXdUAwZ8N2p6PuqWvokeFB1LbBfWlEVZnWyAFK+xeCwr4feRvSARI
ByaokX19jq5hIiqtdGLh2T0iYgmWr6J5j2H0r8F5rQf59sW09/DopDPKSZILm//I7o1EtnjSvOWq
5SL7qd569gMWwzMt2nyWfxmAB/OMPpxCYk4KI+8hc9wVitr4BR6lz1BpJyKeNeejzHUHlj93IfpV
dKU/KAdpGqx+SFtOl5evynWuWB6DlWkH1QYzbg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 69472)
`protect data_block
2485/cuSVk1XFaPrmRWYxDzK3tBuPiTiSM6MlCDHoe5Z07I4MSOnH6Hkbvo8AmVtaCzyNX1mZf+8
SYU0j+FYDCXgwSot8T9VDNjuNydTV8+RGyIGdeCUraYQDat3LoXjAhiRv99oWvrMbLCHCDxYcfo5
quDmNefSuUKXYMIcQpd1XH3dde+o2CiSYSmFeiacI+qycm2ZPtWOS3J0mFpbAEc7dGGrQNyR9kZy
14CqP9gonjJijbcNGJkFXXNoICNraXOmW7kJPrLF1w1L+vCsbVLujzFwHyqUjs30eQOMbW7wNBsO
S2vDwXvtTqhazB8btADZHCbOkEXyRN+Z9yPeyH/AkLrcNmOfw76RmuRFiWU+1n1KZJobCFWdlvOR
X0CPO5vzKyD0Dtuax7SYqMJI6BO2YQN0EadGRjr1Pe4M4fPhfzEAtEGoDwOITzXKd2Xmq0UXphnw
aSc+96tj9edwggHKJ54zQApdA/5VDcJwSMBtEUx4wrY0u9ryd5knSIH1QLU3uGyXIpyC8MRxrzE+
Uu7Rv7iLZ88fKCvtbeBh9scxaMn9FJn4miGoofKWE3IwsJ67L+eY2g7OwJ4ZdjR7tTI1nMZegI7b
fFBnBH4wkeKFQkDyTp/Mwpws2zBRCgOid+Z6JjRCheajsm/k2A4qxidnwDWe8KaYSKUgvBT0miaX
Kollhj5tnBObU29cJpa8qq4YnsVDxM8HcVe1Zo9Mt6JSxOZ9z7tNKI/tuJKiWT6Ghr1BZXt02rgA
AjtVFNAbHc35Mat0SMBjX06iF8tZh0+NMAuAkEt6/z+d7EkX87xg5cYAJVVi/6pWgwrslaY2zNKF
Bu5dUoy6zgXb0QttUq4yDa9WXRdZUZ1Ha3bh7/MZVZE5OSO1lYydtiU2fz+O8sqjZKOjv+H2sqlx
8sFgq6nq2pYDBs399ocFHDxwrp4oZNds0XD646KK5j/jCHNxByY/eT5yDZRgVi+1J4ZXYH/peb6i
geoW2gjy4kTxe4rOZZ71BHW82DRBuglnGCLdGPbRVN0FJmAcqP2SaJW/N7Hs86LlbGj9NaRZIRO5
jZa49wqfzdJ5m9sCx/ET3ZKRt4nV3Fe9iCrsBg3iSl+DsM6JtgiTX9tFsskj7hJ2xEolVh93L2/E
6U1gf/rGbapu/42fZIkY/Eaa/zd5Nh4RWF6C7sOtDNHeJW6WqYt0dPLIcuG1arPCunxLZzsTFls0
xMldMux51ccX7robhlsV5u7UNDDi9ulq8tLsfOd6ZkjwRqlaLGLWNVMNPsQcPy5RssQB6/1A2Egj
5cg8jniAHT9qiakmtL7m7pp4ZzUPBAHtw8POInDz1TRsoXhWn47WNqvBg+grc/gx4zpzZlW+QVTt
93Cpl90bevbjiWR+nK5d35SW9ECH255Jsq1sajBJ8FAQQI5MmyEoViXSCOhjb4P1klPn2Dsa/PqG
76jbiRpHL2Lc7/N68Sf+XPy41jhOhhD/g2T83XihDDjMvnAJ0/EyC5dBNOPZJsKQdDImQ5WTPnG3
8Q8R8iib7fnRSHWrMDi98aQLJEypYr9euHQ/M6z1k2bdIiHfy2bKjx3bYdt+zVzORZ+oW0rR/X5N
VpLPrYyJyARQ838ZmVwOEUgZJJBY9aQRsmv1UuX2DDwdBXM9JUE3RqPuicuVm750dDd6ftaYXuTf
lRxX2r3iu0Il7nfndQrFhNjaWF/IkPsIowr89ilZVjSh8X429KAGYnXG5VmuFpNTxAT6rUax0Mny
ngoQhx6yWKwa9XKOV88oQsAfiHPc8IuXxu/x1SUCjggA7IygcUETXMBnYF30PnRqi58obZY6aEPv
XPGHBqO1exCAMVOEF8vYVc427tKLytqM/9TbC5UNOHyyAvlUmoTXfk/tQjd2TAkgK8rgj2iVRSh0
o6TPBqY25Ln8vfDmG2+kPVWSPN3rTO79dIM2/OjBvO2akhMNxlTUhLG+ovQ2y9nK9mr8Td8yKz7c
dxoumNWgKsD4r4BYc9YM3BYV0vSzSg0c8+mEutm+O7aVk7gAF4zyesZO6S+GkEvqz1KNhAvKx6Vx
+tI1TU95tq1tQWVFV56sGmtDOfJ+vyplpZiO/C1UAmvU0wHG4C5xZ57qA5gk8Ctj/rZnRkKpSdiq
xK35a2ob6nXa89+WGIWxQHQ01KolWraiXfTc5LZ77rS1k5RuinlGu7fYk0Ryq9dVeTTY9++MdY0b
jAmJI/jdIntzgeCJEFsDTlCO+lJAUcSaNKUWonDLtw7LvGP1ipve6larbFYC5hsJlg1SAffExzf6
tBnVM2kh7IxqKFU8QcHigRDeXoVTdPnr5Awmw3Bc0Y05QfVeRO/lnnDegrKj4NewH18knEmbL4RQ
B6s1u2MWTCTywfPG+r1RPqu6D0hhj1hxC9LQbcOTn2CzhAjbpYQVNx8gVfporoLD3Nu2TXsSZsm6
G4tb90mY0WRab+LasvUcuM8PyoO6Q+WB+KWlqoRAXzE85FZMV4k3BMSMZi2IT4HVArRPUHy+sSrs
qPGU7qL/FgQKbw5F5deF921kc4ND1+hx+M4kIDB23+Kix/VksC1ANOL+Miz93fZ5Szf7Q2i0gb+I
gp8T07XACv0VEQXfrlVnrtKuX+nnEO7Wf+Cytxarhh0079XT1A4fe0X31Jlv6kPHvx0zKgPYrVlB
g/uLOFqYaGheua7XYYL77ql1rXdKgtI4p6wKhwceb8h085A7jXrt+ysd6muokGDcfEYOmhZuN4lf
qWXytqsg9/NG/9cMALyeReYlO07uHAL58D/9V8SXLDuEXG+RH91NG2ZWp6gLD2twJebQVyr695Y/
MYwTYbrSi1ytaiAJZ8HU7fzF4Vl3tybuWn13WXaOYDaUMZogkvVah/M1VBW46zdqFf7WVw7kuDQv
daw+9B0yFUX8nSoxzJPxcIGKaJCQQLPDXPgWz+3NHrVxTjaMDd3LuyGTDH8TMmcufNPkXV57W5TV
eU0F0HZQzD30ENlTwSohzXLYpav99NbEN9ZBtjxNdaxExvUd3H9HaphE7skJ+dDqJJJdHKzxURi0
rSiyDG8PzK9NcW6aPE6j3XcLw4VzgY2BfkrPFOaGIPpWFqnAoSUz+D7uiM6LrO2NFsS2d1hkfX25
2nvcSr1bqonEOZWRdYoYWXxqhVoJtqIELJTsLvxU4MXfcxdNPj7FE6ihuaLsVe6BcmLDr8zE5w97
pXbC/P4vNdOQMNaXxPXUOQAY4G7cnJLVa0JGo9kRrAE7FwupHn/4DNR1zfPj+WRT5gtQo/T0qKia
LPhphznK6fd+phefnf6Kect6shqJJ73dEQwVZP01CZQg+mxQ6Hs6jX4tAF5NcH5VyHs9LUX+Skuo
s39WY1DjZurK7YQmH4gL6tifDj+KS65hVYPMtw1kmZ10dW2OGnGG/l38n0mghzt2Win4YEg6YMOm
LfjDzvB3ElG5n+22nnl0AOKVZzzXGo1+W69zWKd6jMSMlD3sYvKH38WDYhaf+h9zFQu8Peu5AXHR
fD7/y8C3KZjQ8HHIgY7mKiCBv+FWo1m3aAIRFBSidHEH4VyKfXyOJ5YOvjpRM7N44GidZ+uHEMGI
9cLdqCFzZKMhDlLU/Ro3Ap+y73g3gWvD+aC5Spqw9Mw24vygWq9IQPsZ/eTUs1E2ddWYVCjLnPjy
C3NTpllZMI6SEjjXwQ5/onZhIHijdDm0jhHckt95+3RMoTGb1fPqKylDgtESPp06lBRweAagrhEW
ZkXAd1dYXMV6xlYQAVHVJ2GAuJpTPbZ8hlqBpB7/UU4E0aqNsfkzzYUykjQBEBBAUwE4hpQ4j1OT
PklWWr2YOpvKgmRljHhBIKi0vmH6y622O9kFC3FyD2xx/xe0kDWcNmbb4zcAJ0JfQ6PuRLPyHT5g
ut4UyoaMFN5UN6gurrOrNoTy58TJNKxuPRhktEGWHXF1bk8S8gjME0wXl6+hi01aGYURfL841xuQ
XJUFHjrsQFyGomeRGIQKzZqxAq+Tea04tPEzGXri/JF3ciafAY9ceDJPZTy3yU7Tdsg4xvXEKdwK
ALhXi2iXurWkzjX0O8tsmhsjYWhfDNcMDOZa2/OGltu//Rlfw/JWMPhIlaDF3ZczMaKG3/NKL+T5
er5fGknK2BINOOGuna0MJqPCqiENljANY1uJgavXxc2/bUfWCzCAr429O50XbWbwU084bZc6SniY
Ml7cMyqXqOgcNA5n7/0rcUii5r4hJKUXXz2kStfFIKXvXJJBel6WbP328QQhO+VJZ2JQQ6wHLbAa
twPY/U+wLr239dJaWUzx+6SHipbxx2bSjjV165V9hi5Nlf37ij2WUHGEhTRSQ+TejNXhABXOYrco
wr8AHcrvg42s7DnsstoS11qmBJUFT/Dxs+EEb7mBbOFDTnks028IZQMPULYWscOjf+YuWjxK0mOe
15QGsf3y3J1onMsV3SQx//H3qVpgFXkysy0Bys9YOfEKEj7Miwrag7A7mT5u7ZCGv5XsBpD1HIW+
IWKJob+JGjUAMkztV/S/h8Zz/N36TBAu8RSZ5rfW5EvqFICxVDYrltzYLYE368BazdjmQUOyKEUN
CIxy0DgnN7vWy3Shor9GXy6JK0UKwsc/KelUIJe1F+08TZhaxvkBn/2av2NjFPGGBCsxPpyPyYbJ
g9u8cc++s7W5ofg2/vJsxbPnXCUgkMThIrImPA1wspBIdG+V4qDLD3V9yj5XaMW/PbzmjeHFachU
5BZ7gM0F8X7SplpSFPwJsWMaRRbCtvRBWy/OEHhCQIjWf9/Uo1retOdzINpYdaEuVKIzDWZ2MCsU
Pf04IOpudA1bXtJRnos0HD5WxKyl+A+w9FnJuAytXTvFdoiL/tAkLAvdfy9MJgjvmThOTZG97y8y
dzNc9tKeACnozrvOpZTLqk/zkQfl087BzaQENCYmzmZmeVZ4zP5kZPzImipT0V4wXCh4j9YkG1zI
Fyn3UO09pSxy9vVq3z0zPa3GOpn/V7dQLIxJksxV7WLkJf3F92xSVtF0blyEYtLq/2fKTJP5+w04
yi1pjm2MnhbuuVWpsAwmAI2Wviv3Tt3MnQJJvmVbQtfz7PDKG0k207hIuHtHrtpD3w9BYdZ+J42V
bAcovA/M7wP0qAQozc6MuzoHHfJJb47/VZabIPT49aJ2tVdgrZ9JfrZG2Nd7ahuiu1Fr4EHDlgVi
FBQcmy8lfsu7mujecKfQ776A/JmYrf3bZ1Lke9eOaAYgtBU3jXO3qhlyGWNoc2U/rnouSt9fw0nD
OU+xZBCVVJlD0epqAJS5JE0VvlaSSHkKWQQ1FRL4nIXPS0Gh1CKJNLnWMkXCk3Wpz5JXMHtnyzC+
XS62vBZ7xnAVe2hdGJVh3U+Zj+96EsB2h3hu68ZNaeMIrWnKCzBfzatwN/ZyIVnS0A4pqbA/xo7R
tQS1U9AtUm7xSqPj5+a1OYL92ji3q4mZqTraY+yC1b9if86xE7+zOivkC8PzjmPeSzf2o9nJibbR
amJmZUOn/y0xlMjxKvkHIDNjrOGgvUr1GEYSjH1erHuyZE1YRgJyvoCDhwu3QHIHmjlWQKseNEXL
RDDL99DWMBx4CVlXuq9ZOzRJ11fnT1g8H+e/hYQvTvKSeVbIB4Ad09sjquXQpKqSN2g79yo5DbhH
Lz+5NJfMpbfRxsrXJpUAEM6khEk9/kHSAf2GPSP73j/h3+P8JStY6GZ4Q2sGBdLHYF+7OncYvgbo
7Ij2xmyA9G+4hzSDhzZtgUs771PPqUiMY94Y0JvCSsCSHrwn8TKEPOR5zTPeBM9bZYYSQehDCmMc
BcUFgw88zPyqBGv3NDnzryYmvc8Mp8nyk9RR/DrnA3FdoUk2+RiYH+TEcokHiWgBLShtrZJOnW8G
c2FMuz/mtuXTj6RLvhuwU+N5+oFtjfkjAob7iCyRb0pLhk0dDB3WtUYBbMG/R4y3nEo1U+O68iCW
O8D2w3Pwn+/mUN/WFKAK9teNEN2CEr5HLgIeEwyXcKiFwxTGs4U/Ed1BM/qQg53i2o5ZUrUqeRWf
dg686M5XFCwuAsrsKqBqrNjKkfLeEqp/cfWLWnDZGksZQqJ7mJjFH00ZDEYNZbvceNDd2sfizXYa
arlpvEEDDr5SgN4iuxbOVDkul/h6xMUsDz27NXzR6ZmMfqT4yxzqulXFAMvd0l1VbaXouFas0Duj
BnMoJ9BQTj95Ir8cf0Femz/+wWzbl8fI7uTH1n1JKyzgcH1101TgJyyOmPyVLPhNbJw90BRu14Zf
FORaPKTTTjru0bhbn57dapxi1CocRARAZeaPIHtOAoQcrsktgHANiMgmz1O4UM/zo+L4ju4RlduE
Q5V1bK9zLAlaAN/Xt+qQELcLFONJQm8JXpeyuiDAEWhbX50zcOdRZC9wekQKfX3wjlpC/NMqC8Bg
cjGb9jr5Kxm3HL8VG8MgvbzrraPMg/7wfl+a8VT9B2n5AfzgrloC2qlnTSDgg74SMEdqsSt7yYvg
rTYop8H4/5Mke+kUikaGcAO+g6PY/cK38+CMDUl2lZQbL+poyHAlThtLaVsc+EL/yM7m+Bo+h95E
9iN9G/ycHYQWFkECEeck5r60ZZWqGmVS7wQdefNGOcGGwyUfPNUFx/zAJ/GG4maAS09kb7SOjTm6
suxOH19jiWqf1kPWmBSEAYSvqoa2DgCxVhVdvOPLefKADS7ZYsU2j90TZVMt19Vtv/1tNG6a0l7g
N6FZZ1bII4d2iehgMeOtaLaz9nxfVeAM2Tq652Bw01OvAmnyJed8lcFbwFd0HxN3fpVORPENYhaV
qVUUHZMjaxaI6ZwkeO4RWeqCEipPa/feVwkSONv9Kpg+w6WwCAk2bDVJngD4ZJjJh0iO29X/s165
gLk+pPJZRjku/Hvx0mLtYPLMBKWrI8E8VTpTlCs7en7ttRvsiFKianXHXPM0bhhUlLl5+MnSVB9C
A/DZqp+cGMmrQfdN8xMx+L0b3YLDmMJIACWYLXZGIeyO8DBhmvBFFVxXfoZoPqM8JfVC3pfEcmrs
bZIUXpMv1aTrENnrxZRCzq4s2XfHSxX6UK16+FHPvyugrhngu6qItNsmwkFVb1/mt7+fk1xBoLGd
183hTDeG0rNqH5z8XwQsfP3u2ds2ZxXK475Bvf9T/nd6lTCRSzeTG0Td6KPzZAfMGAPppFSgbrHV
y3MDUnC3xh33xcGCTZP7cX0DWJQ2AUcuuO6roQrxNvjn67nozlikwxujdmG73MoOgNnOlXWIaQne
vEUwLb1i2x+QEQwclkuCfr63X3xWihEGY69xJimxLmaTAHCyHgOfHPAM2AzW7Fo/eS3IRjZMMsQK
IznQAtc3jkqa2ArNAicwFxvm5y1NKr99hjVkWvEQf4z9KnJB+QmkZVBeGxmjd/4I/tUSrwQNNtsa
UBLh33AQisgAjTICyIYzMrpu52Y1wletE5MctItACmfrdJOvE/0voH9xAkIXJBuiQHqjJZbHtHRx
5LI7ddPmO3FRNF+GAZhZwwidlVWnTO6zfMm3/h16pt62/WXnKTTFm8RoDTPsDdut6PUxzf+vaJxA
Jty8aa6KirfW+Si7471KcYYg1LqK26Ua2XkZ5G5Du2u94AKgJFcuoqe3M2yJ/pncH/lNTnMHjk6w
+g71uM2iFs3QJ0cSbIej1Shv74Nh9LZJemFFfAU9lycL0WpB8xim9GBFBQdNn4IM9HGZs6tb6EYz
aL8N1p692Swhy9KZN/XYjDFw/2/mjNlUlZJ/h0YdmDmGFOQIt9h0fBCMKfmpkMsZlLIIQ8mdvIFr
PjYct9Eiy7ECM/CqPzPju9RjL8fjQor20mRr/RVGooF1YHobHV18Dmt4skpMrhsF7eW0iHO6Dw+t
tx1AiFLKDxy/230yQnKb+LgkupUVSdh2FWQwkt9KBfFWLPF6pty/ZTdzrSQCqt0gOeC2QK0SFNZs
M07n2SQn8+RUbYdb3OEMTbmQoHVNyPHTbm9B++ADsf2XEqNa8GP7UHOtE8njW/ybMfd53CmEiA69
mFCneeE1biGGCzahME8yChnY6FIlAwCEG5mMxZz/LNZB1CR986758JbATQ6LbuyoC4Bl9ca8ytWP
x44xBtLJlMRtComGQ0DmHmMxTh2xYfNqEItn6wbUdoK2Oy12/y3X48jNA+hRywqrMohlKgzw5psH
ryAQ2UMOnEKNP488C47qXgCFuKcxGGl6OtnIHQCfCesPVF3x03J1bM7R/fjNm/IT+UDVBwQXh8aj
L7Bu1nuzsyNqMBQ98yGM4h/DgQ9AbS3KZmKk0/I5hhZi6TvhtrfGMaHfzgjd25qW1v1FsMHBV9po
KLQ5KSyicrTlD2WW9aJYmGB+6dXmXpiNKaqhyVbcmZwdSgrENbqKX0J8WIqx6eeeZIwXEyMxfawr
+NoB6rWEtRJZ5Wh36/cVLzQuezDxZDQ5JL/RO4bvWlRCk9z1DirPk5RRpA8tUHAp2cvKcSQ9qjSZ
HSx0XikrrJN23VFk71xu0j0XLfGLwNYWEgAigJDKFXTNQ56ZZaDpwWOK/9PxXBfvC+ozuOd21j0w
z2msjVs4uv3+BEYYxLTV2BiojYl+mBzdQFBbtqHAegUCjEN+qLssvuw0k8mQEXr5l7xp820vE07/
CzpheLooOPj8F/jqv/QIuKYKacoNDCvx+t2rqUKcf4cPpZdswmBrF42vSJWPRTTXGjpdoer5BhQ+
SK5tIjB9b48ib3nrFzCjzukuB/FO2LwARLP3sbN0kkvB0zQghuIKxlVeHzGCmUQIavVLuEFWSK5G
5blYQsu16yxPCI+upfxP3Nn7nxiIt7LKI+xwxDy9UC0pKiuwzZs+4q5z/MTAusicxzZ3x975Trer
ewLmMZvfv1c/YIvf+a7rHlMsmuM3O96O6dxhF57vPu6wYFV+S/RSWlAZSiWuwE/qt8l3Qe39TPK2
tmTPZIfgTSKN9rkXPVXYm5kU2hOpXJjmmFdvTBz40rzXPBYYoz52l+jLho+AeyLDUznbHd2CJqN8
vf8/gTLpfNoUPDLo7dDjwuyGbBpZzMCHvQZupSThrEu1Q45o3umgXhlg8zXGQZT0OapG5Lzs3ONR
GoNz4WTB3pYxlZGsJTdyuFH2JScitTjgpXNjeA3WcK/mcTaOvEA81azG9e2NibqjBjJ7Lv5NoKPV
uicCGpwtWbaboKHCDro0qzKTabISrsh2gT03LjEF690ExLWHkiJvG5i3RNSZuulj/Kz5AsL5WvLM
slO558opdqF8KtXMTaQnAX4kWwHA4WQTyCqjpzc74w0JHWzh6fA2RLQphJOBf7uvH3X5zDfcdqC0
0NOsAl/TtsEnpmjGLObgHkN03TnpOBFZ8KZu7dtORZZbBLjXKxUk1qMjzsAdnrpz68PF7phX1BuA
rQ3LBfbqtqVB79n5Sk0Ng+CggWn9rsvbiPVBLAtA8vSE2lCBVQHHVoScGjN2Z5Jbsb+ELB7V9O1W
rr0hC/laj20lYVcfX5y0zbSG6EZ2aZO2r81+ekp9PmZmmE5xOc7szWAP6LiCCIHb1KNeMqZq4cH6
oEFVoihWcaPtJXdTjIZ6wdqfOzY7uoOdozZaOzUZincM8iG4akpPfZRUevlx5C1MDuOEzeXmjVSS
cwodaPInIsGFEZZHhdYGCTj3iWtZjBNrQvdv1VJ7uwuuEH86xBNKNnx9gB3/EWu1+0hxAi+El1jA
DifdXtPYYj2QgiZxl+SIRSLbZrG6o+DwmOaK6yD/xBIi54qtQmESR6bYVfokpyoJiTreYa5jpujN
HDgxVjqmTS8pMpuUKgNdKMx3lCipaV8Sl3D8MdIH2omz16ftt52eMFbVTHArFCvf13zXb6dcNgYo
2YXRRlgYRz0hL5WuC5czBqPFb5S9UuNFiALF9UVEh+a0fi4HlLJz6E5F3+9zjhnrw01vowugFrB8
R01e16ZpkpDBeco7N17SNJXZrsblHJxU1Xh/ZMxxhHN8CBd+I/K2D1cWDi8E9eA9a+1IOdeNIt/C
KOffuCQbcdhYUO7zZLNoUegoyDoMDmW5PldvOzC+tzg7DflX5z/XhEw9KT4sos3x2fmcFF83jeFE
7Zgx/PDy2lSpM8X2Lm3RzRP0U2OFVjUXx7SPGQXRDxw4bJ1H9Kia8E6f9QuEWm521r6Ulib6vdbC
oPEBhve8JjhriT/CLm+I7E/XN0vxTe3Udzc3RxwIIg3n9pKP0dUDMSqroD5sLwh4xOBaj0xaMhUs
Tj3mNL27/ZXIAVvBKvV2JzcHKs8W/PXBG/f4x54AO5/5ogAn79MHfSCn9ED2ScwPTxNswkMsQf/4
iNGcfxDL0GIcrfk/JlWZS9wU/c7SfYWsitSpNFh0/TWMOvsbNT+kAg2wNlKlatJoEXukKWcZm7us
S/s/ntnOcnCo8qsDg5HhNQUVwPDEIRiRrBzxZnDjFB/bNjyM4WQu5AY5jeQ+/GGbTe7Ab2W8ztFV
+UxgIgoQ3Emt08MO9IO9bnelixSB6UNkXwFfui3hSTUK5AoyrKVK92NKeVooE5AAzX4PRBypd/R1
vs12bsBULuDO77f8QQCWgRQ0Xkn7iR2PDsVZoFqZfxH6d8BaPX68ZnJLiqEPBZqk38U+OGWyU6AN
qn54RwaTi4xw/RMo0LL232Xrnu6wZy1Xe0TfB0/oE5BHJogNr7vBuH7+j2dXInpoJAWK9djTXqh5
hzL6zTsnLkm1hu9xQqmYWrBC76tZb11vW5JugPiIZCwOgBz35uFrqteV/XeEUown1jEaJc3QYOzo
c4gyj1tuLZz3TpFwdE1Txs2KwCARChhF0Xdmpcdu3bR2n6MMcsKWlIOSS5qcX65gFe642JAtbvOa
9w/F+YHLSlu+S4XGQtC86VilrL6I+bJsGWhBD9eqeg6zB2mgwAYZhfLoauNncsMsQvAndeq/pNyk
IjloIB9XZDsbwloICbQtz/hUaGeZGQZ7JjiaGv7gGvkqJgtwrGvJtlMnlGFf8FvlPIKc+w6xa53+
NrKuFj7JDlvkIet2fFzMU5MoNprMGfTsmJxn72OWFPIwpSOqLsKnUdTvO54cwHKE/RfaTGpxPe+N
k7o6B6sHCpniZuff7BJGjsJrwqRpUE594lUckVxzZCKkL01T9OVKNlyFbmF4tEFRLo53FgiNnCq6
HWA5tGmDJWBgmpKxrEL8+3vEucpMgqlosmv5uv94jI2wi+IQR5SKpcuNszdj5Hjd7bu1wRUPHCfX
SqkmEZgu2NUTAhcjB7AdgmG68/X4/ArHc7Ku4XReZWRrR7KAA/p9ODS2QCZzqvQcU1r0CvVN28/f
NjP8b29DiUTe7Rpv/NhWrBvALW+FjOBxNNCZzowMyNfeMG2cNoc47X4p4bBcrEoqYGi+M5Klw3Mh
yUBikyOpX6ZWpB91VSECc/XImr3DK14S2pcrK1HbpLNLuvXEPOpmpFOiyMlrOzdYe69s2zjt82Gz
wiihBpHMd7xlmK12aSIhqKbCCFl8Kz6CuRsCzsCQnd8/EriSDb7xbUR0E8+GUnIO93i5Ifpw8xZd
L+hhzamR4kkmtMjLUwT1x/utlpxCpQcWI/TF7ZnFe2xF7oGyaTHoJLcbK8FfqLjhi28xhz1kU95D
xwnJ7sX8QDhA2tBC9m8U9avx3OhF4PBvb4LtTgsaQbFkYBvFJgyJxgmqMUwdpPnqzR2/eglcitWB
zgbJWhkdsp7q0h3aI27PsMiA07ht4DKoQgYLIdr6KJnFqRq/YnSJmYT8HTnfNI2EbNwgPZkgpChT
p3+cMx3l4uepauc57xqmNKGYo8LMeajFM0J/r6qqUxSg6DWaMPKtyCdjZNhupAtfzBhq3a0Ldqrh
upp2Dyi1F6x+IPnJGU18OXvttESfclFhQSoeEGPHUC8+uRQ/9YOM0xP+1gakwBbuNBboPBN4bCT0
gMs5YkzM0F2mGoxDR1CMJrGcxi1FzsNXlO/bzChHeCZdioOrNFgF6VVzjJkq6VZuwBIEcJrrwKcT
p41cCUJZfLIQUbAwMsBtmikBJ7OCsGtgfSgiqJxStHqfRwn5cHzGr7641QIB8yFeuqKTUSQ0gbcA
aN8zSjhp+CVupIPFVYonXfwYl0OlkuokkOd52XYOJlrvuWAMzYqcfHNbO/z/J7h7KxULpqI1dUkg
8PDpssImB6GWT8MHxGAnfy+tqb2fy4uVt6fl4VN0YiISwDb6kxWx5lehFF6eT4wlK979WZKcLX86
Y8c8IhKLLf/4Gm7j8V6bawIKSNcaWGvTzH4g3/ldlMh+HJxZg91PzgLp/qvJJQFwS/CrILtGkg7G
tbFzJrJZwgMXBAQSU+DPTV/yoeHkEI1CHnfGWbFZZH4Wh2sAsU2rKKIMZTQt3Bhqy7rD0Wxuimy8
EX7DLcVyfGaqGPE4AUbQg9lp4Bl7DmR8yar/G9uUDaAAfETDzz8FYFQKam3v+/OFCerwQFtXoZRu
iWEtWfE1uSnPoK0pbvwYprti++IFzIF9JeQCNd3aDHdZH9JbYUDDZwiO4glO06212QCnGEC8rakN
vAJk+bdnKtYoJZVhWK95bX7ibo2zVvR/KWTVkW55UGtWBh8YGv2HDJpksb+pwJ0G0tQFcyBRXJpe
YXWCyL6+GONjd+lMtTB9s9UIdCh3OvkgpoSp6IAO6jS0yE7sWBrp3Nj2lwfTOVegBT2AhHw0Uy0b
rdB6+hB4WCbctw97v7N2WiPX75eFvYA52N2DIFX26kf7QgfNqH9IftAUMpuXFL4dxmxTUq6RrXln
6ej58IRP1AHOZRvWkhgGCUWI1ZvDn1oyD9USObIsRJtsoc6kqoETWoa5xzT+4RnDobOZ+k3GQkZk
xQBGPv+vOVrMZ164kXkSm1UdDgAQv8ALntp9atlWcnDK8MY3T/4sTe0csHxHg3+gDVSeyBOTCaDO
+uwJ53iP9zOFXzplIJOoGaBRyOVmwMwgFkG3VKjVYpDiX/VdHXFyhKTnBoeZwoVSQ25vFSqD4xkq
jkJZP/TEqaVS7NWSZo8z6zMMEnv/8Q4hdyZ1RIdEsNgQPeeE6jWAvROIg0NPgcnpAmuBbBFvEhIA
uI6xGqFmjWrgYuzslGO0RNWySwjPqqTbuLbIdeq0m1OqfZSjzDDfR9FzHeKhUK1TVAcF8ICUb8V0
bWUiMg4r4NzHLZSc9jBMoBmr9CEYnVIG+RB46IJ1Na8tPXwkPRgZxX+6mUMHcMfQ6loayvJ7Vty8
JOvqfWZJGGRiGAYYKzzkPVMH7ibKSp6lRcZiHu4A05sJIN6KmwP1hgGLWfoFAXwCArukJrIoYNyB
JIsAkyN+3BpJWa1+3/Z5JwxtuerVauYGlywckY6csxtmzMx3mY13e0kHcSoBYE/CW87PzH2VCObv
j7l0E4y3qxyriNMY02zZvaBGOXxln88+vv61TzO4QzxkbLwi2JILA5MlgRN25Rn4FLsnrZJYCuV2
3OWAwNDiI5MlrCUu3+do4qeo5ooTVC7w22LiADaRRWQISW7/ghQTSy/hOrrJtBEoHnpkoPiDpj32
0r/t0ePJyVENVH0YXPwr8rrwmgmdtV9vNTsraOjllkD4zxPqhFczin/MiqmSDBP2p0oiWp8dHCCT
jAXmaaGRFmoq26gLhQ8KbmqY4m/k1QIXWT4jXpQF4Lax7LrFpcHDiNbxnf92Tub5hMSiVK61sEZi
Q/QkduoAaczNVqwy5mTcBn6sXrJhz9SpYNd8aR3FIFXYpgBKGpapoPkcCWhRk1J20xl/bAb/OxuG
z7GV1yPA1bjPt1xe87vdMDjjBcnf2GEnfwPyssL74f+h8BCMZTd38XhvlfrgbhLFp/jJKKMUPCKy
mj8/2uY6XFURSms6tp1CKjPDaLuLWOzl4cKsxiM8RtEZesO3aq1CuZEHbSMJCvNURevCEY1mhtQr
NMmfIsiKmXbbvSwg+iweYDuWlJWHjlA1JvjmjVEE8f5b9E0GU8HDu53cXxKgB7gKUNImbFI44sm9
ast4nKswbNAjCRZR0Rf5PjIeMt6nO79L4e3xvHWMCIPq8KPx/Dm4IZIhhvfdKHUm300MJRAeUSc0
aYJjF8daSmmffI/edwhp7fUAjmn4D6M4qW7ZSRJ0j0EicTgCQMN2SX6iWT91pcJX4hDOobaMZm5C
slhOHoFdRKnXcb0CvgwKDSNG1IQF+DUdfBr/c+y13netO7Bp06YPSirv3HOczL23RFa22wmqXwMl
KYjbL0duDlVccslCqixV36x/UFrFz6EDLBs6XzgcpZcWuCrk2azoVnwteAy71jioE7jivSMppRDp
5NfkMZNwwm1BUmIxNzBt0M4O39dTmfkJ+DHhg4lpTAXBgYXkeIKzYavSeYK2JQ1jsobqELBpjYCF
mNNldMztPRgWPFxi996dEoFQ4Lu1o3Z3kxk647EkKMeuEk4XhmPiV0UqDD9r6DVTy18nWIsU28N+
bPkIgB1y5lZZwRCrhJyvd0tNhJ3I8EcuViYKW9kFIKYRIPj3OC//+B5PO8YakaTGmWCeyuCYZike
OkqIT2nFxkaWIV5DT9105yJGrgPeQ9uBC7Q4lJ3eKu3Ggk9nwiZdj7D8x0ULRc8W9rIXuuKVVJSV
sIIqCirp93VKPzCqanl81/TuJxbRiX7X3uunVaIR9xnaCOF2OWm1QAW6MqFjacmLHYMk9CcpyHGG
ccR2d4n3dPc8cXVxS3KAWslBk6hpUqe3YylRmIzZD/GQyQjh6SYWrgLZddnz/k2JbpC9T26v+A8z
Q7a4g+IYOEv1IlvOkJGJ6wrEheAQHDssg8iz8DwqyfeD6n8h2+AmOZ5Pyf0khr+YmNZvc69xANNz
/vuWGry3a1ea57Z+t6TC+K9y2KNmAjfzTw/kYKSAOgRshyQSQ2MpsthLnZPmjsaAash9PBb+aa3v
idu7FhbcLipqXuZAzIDrEGqdKxYRcqy+iWJfLKOpNLMSo3LCYks5xIMEwVkmQs+ScDJz6L1OBU4f
p/ZQzAVGUzUyKj+BgQu07CKiVbzh3PYpJW0uyOaRFW9KYHvJS17LVCrXBv8kbDOSq892I1aiqjo4
z+pCke9i8d0mtdOEsQcfwuoY/FiJrMOcBPve6lPwOkBj7oghdKKIdQzus0bNfomEPydSTrM3Gn0w
IvbPOXrZ9RpfD4QiUYLz23maQ7+YFel8Y7x3IpaN35qG4dq5gtaKjPxkk95nAgOW3M3guaMaR/qj
CeCiRTfgfhTbk1alxS4HOBpTWYoa1q4365KxGEukQyW3I5Sq9mNqGEy4riExCiPH0D+bh/IAjo/H
fuZ1r4QdPG4lcfA9jEwIyFoQ6QjMFXScDavmq5gYDb2b29QiwBRlLUw3afiIfmXbC6rN0a7AxkGx
YYsQ4uFHYpzHPzbwzKxPawtuHgeD4n4OFBT+VCrohIq47SX6WtvzKIPx+5shUsR9itTQxRwQxP1V
ERCfNP6/nGIfBMJsePsE0R1gzuqB023fbxWIP/WTLX8frppyaFBOEwu7LpBWr0NiiAao2s8xApH0
eigHeMo0yTUf2NMBgMNRigXDTQSoxtXvygHCYs9qc0ABSrNondfuAhuElOobXvfeSk6P3AklREZ7
1jLdGuGAo3I7j3ADEL8ruDki7J2pg/tqOJe5DLOLL/XUOR06qNSUR2i8JfgY+bXk/OtqNNg5fJKM
U7SeXGN5Gjj7l46LwtdSJKilyWO44p5fUjcpglh0/YjccGE+kxqkukdelF0JxiAQrx4phCv1sO2B
saXYYIgOqPeUOJjFpX6x3xgsF711be/DUD+CqyyO/Ox1shcqGtT4mOMSq8/mu2i2IuMkVcpUY0TO
FM9Shfxl+MyV2QKxcNYgSL+UHy5B6Zo/kv3iKFfsc4kbaWG8Qx/9W5IDh294Thwu79FzlVrQyTZi
P0q8pRojuud9rhLAfI8jRZlZmBGbOzGPyPnri8VgnagwYJiLOuUcNa2phMxLX7YoYPTmVLUpKico
IBZizLT7rrTCCtihSqRegcApcs+LKcOb7zP41BPRDyUb70eqg/jGkkAHmuhQlKa94TmhYZfGeT+u
jX16WYaOGMCWv0fpkpGGx0bmLzSKVxH44kUxoTwljXVszlRMhEZ3IxnND79Vf6mYla69YmMoYrJK
ZnHmx2Rqp4uOgItXRqSSpl7IcUT7VfdZl6dKlMua0XGpRU9SD4+1qi4ockbBOwsyftGsvkSZ9CU5
FrJ0+Z4Fxb+P13/wFsJFuJWjlVpQyuqklpXG455VA034arydsrWdwYtHcdJFDK1tHkH7tkr9Y9VW
yoKRGmc7qPXvttqqQR39Xrh+cJcV8NhnPd+qfss91USAu2i2mV10lilrCkRyPaKZqzH7ehnP7lvN
YZmpZ8eyAN/iZPzL9J2wvAuWWrDq2POzlTcCdE5x6BvZc/Jc8awA159HBC1bI88RgW7FitSDs/lF
z1sa0uJuJzRvFwwG1g2VWfZmOwsGUKFNMY9XeYlJFaFnqucTmzOElC7wORRlniL+CuBwzQ+HSkwF
JdcT6tn1u6L5mATNynf8fdrM9MkWlGL28QGRFohQKIwjdKQWGYFxCuq+9cgGUequ7kDVgXsSwZ6a
o58cZluiakZxeq5xLvFtvbQznXU3e/To4Rp/UqruOpgengCmp+iwvz9hyB0lNEs1oemZOgbxB6Na
vl5F2YvPsQ8xEQmT1/8AZPTjnKbCemfcVrjgad+8NtceKZWF7108NRW3KuXYo2NCPOFqddURe8WB
sadZi3jNoRPwn3w+B801kft1GjVQMoyrXmEWfUUndEMGm/jDeONfkZK3YF8ZD5muW+zYlEtHTaqE
0pJXgEEpOpYPmGvJz+y0FzbzzsyRhKg2blHq/JnTgxA2wzCoDjOFUZC0C+Jb/nUyWHO1kH7easI2
yBWj0ccmXAbLXweyQnqQaS9sjUWTtnkZHKNAHrXT0MafTEsmmzl489wDAZ66bgxR78Nh4k1/oU1p
/SDfJnBDo0KZZjAoyTaiYZp2NhAfPgrKxAQBvUa7d/k0TTAo+R8fnOv9V+YmTlAWMteT+bUH+QmE
OFddX0kZS7bP9WC5eNcEoLRPC2PCL0Y2NmLGbmU0IPC26+Y+6qBmWniURV3hXCOfDtvD+Ru+LmOA
ipbWSL6R4JYOC7GFFfvAf+gObD2+DmEzvtGrj9xPCZmlnuFQ/HK032uhu3PA/H+Yj87IZx7Pi6Vp
WxY+PnYgirYCqpPPq33ErMv+VR4Gcv45+JSXV5NbgPsY/pfUJfyApm8THWC8sFfDjR8EzRPgKt6S
oiSVlatYTXwK4JAJ01P9a+0l+5hR7tW9Nv9hxPMEruyyY/Wf1Yv/Voq4vWeoUk4XDuSyyp5owAYi
JFYWRo/FK1uBqaj39N92/V/0TrNWHYG4g4J95WeSNZ8WH2cZmGKQ8wF8XC7UtLt1hp8d2aSDk4f5
jvDS4dTEK4epgXKpw5rwq3Dh4Zc8KMpnlibGghr57Vu6jqjoTVKYyYHiayE2sjhx6LwWWsi/s9UG
/8IxKF27RmEZdAPcMAlhC2NjQUkb1Hygr+AhzdPXrbNEX2xlteZhbIfLZGj1p/NNUxTEiucgmhkD
Aq0UANkcSITVqR7bOAcl4puUMTBf40NurtQSD/ljiAiXK0PVdjZSEbfugR/hl+clWkKxZ+7OOK8x
k5r3PsWRn5XM1HP7FxZGxuTIdLUV/p3TB6mz/+wwX39h+EVhDIf787p6CBHALM4QtbyUzlDD1NCl
ttjFH1ejtvLeLXAs+BBymCsVqAhyH6NxPGHq4Tsa6Ef5Q/5ELer5aAkobQxVcK3DHQAOVtRuu3r9
yAC3AlZcpmbXQUWdpVmsrvbXUbZ9TKPURQTVcgVxSxh2P45CY4EdvkRvlZ+vGlTwW8W1CpVStkdN
9O8r9brmE/NyaZPZqvfTMGhQwTh89aymopIyofj88XTdToxegKCntyphQr4nnrrjF/svtXOricOu
/jxTWsri2P29/ZQ2cTK2xAUexVfFBcoqiciQ4tBbmSCULmMstNO3rE7x8I+SrJ5BDsCDzkM90zYx
wpBKnCUy8HXmU5I3UzjeZHGesB7aXhE1uapp3q6yb/Nw9A5gWWryos9cN+qWc006ACr3Bsi0MsUV
K75WcvUTXIZOvHg+G6xV+RvuG2qYySZBQyrErfE8z8tiAFQxCtrmG0YnLDbqYJFaKozxQ839xZRX
zUPq5/kTooqa2oVe/hJF7zJxPAaJHOhzPorKmpzfbPjODW5pyILu5a3+Z4ybuqpIpr3cKeIZJRXz
SagxechsOjtl6AAd3fuYm3hPJtiIiM6yZ0X2fcKV/0OXrvd3eR+vT3n0+IVpgfvcMjRptojzPcsL
e5/5jBw7bDUJy5LvK6Yp53V26/nwjrcNFVBFrzfZ8Pq37o5MnzqpqFMgsjpdgypLct96j2YAmpiR
UHtJksXwUjAfWxVYhpCEXf7LD0CKeTjGBuC9zeavQgMYYFuuWw91sEg19G6xs6DmjeEVbKgW3M76
0+ZT5jQEXIWf64aCXToJTOJHl8hky2iehAvSeSIJKCZ7zza1YHltcPVE41MHzg1xVbslXnDLW+/C
CVlCLEI6g7FHbRu0RgPDJ2t0fFZ7QP+vz/xeHDecEmr3Wz5VHOKULWh307SLjFyltHZmJ6UAzxkr
HctYVr+6WpuQp18gAVN29icHbh6BExzuKZhw4uXNN60AG6QeM55G5LrJkJEnkXBoyy05l1Wwzjk0
3+rTbn5dJe8ZtXxWwn5dxCPBTNNjnMW9N4en6DYUIZ8DWC1wooXXlhUTfsjKftH4UDpzkeYjzDNn
DrdUS7r2khuadeAGyM/jK2nhN7djWfmj1/6qQexQQ3FP9JJtoAcZ2BTUKCpuw97esbGsZcbf5x+4
/1nZHZX5T2toHK87lAGcB29BxHLUtvq7+BQpyM5EzwKDq+QYnJNpFO8VVY64af8rpiF+biy2o2UD
fmRMxYotK60oJLZT8qLtP1yzIk5x2h+dbWUfkBvF0yEae8maVmUmdELBIcZePesVJSFOTfg2i13O
UpVieMQTUPy1xW0p146Y26Ta4DpKbhixrd/uGafE+iMjutSK+F+SKwBr7yhm+5NQyN/RxKmiiZHK
ZBHVHCQkxGEgD85/LdIIJ8wdDSr5rMiVMin6gDmFGW6bmaDOTpzeKs9bmw6I0OjzUXaqcBRPyeHh
GmZ5qNTyCC2Dy5ovOljrhrhEOoXSFtNAXpMDrx5ZEnbtoKjRfD8Q4TayK/2/vEUub4zF1c5Iyj5s
ij5b4M8wv6A3P5eXqON39aqq6+xyExviDK3lBBfh/WA8hVSt4kY8irC+auTpEKsNGZKMm3C63Zi5
6P0OI2vvsHG3AW6MI5gUbzj1qvB+KtDx9mdLYRSoB6XXw1ChlH8+yK6XutfB1ZGbyYpUQplZWgLT
ORsiMYMkXANLuR7N6ejZ31UxWnVlb3fHFIAiLVfCXRJN3wQi1O0Dct/KDAugc9dXP9bYSHkbizAW
dpoZlFLO77K5hKCcHjQOo53GL2LXpC/1SzuvJ5+lU8kPhCqXJUDr0pQ06gXELlgCzvg73q6WQFQT
4uCqlWguEqBcYfFyS0KQ6VpkaHTLz6+lrbRRDYn5SanJcEK1271DCrp5gBVJvGhvMC4YjUeJWmOU
sNl6Y9wozeXhNNk6eqXtiF4GHksNOruTutq5twfotOPda3iEWNiGy5zbd6fR3Zr/UMG8nOVZtBPg
qeb4Z+VjTZbJlJv9wV56BG9yPMQPANT/JbiZ2ZkZduMI3jG28Rh0cAizU7d9WRf/OEKdx8mUT3Og
aLs1YkStclc2P7MZneS35Hudc5kzidemuFobk5XoRIOWpkNcPzuhajv4VA2Ui4QnSr6myss/KQm6
ZU3aQqz+C/yQJdxWfOz77+ZJNqLnybxctd7muDs3dGn9gKmTHvBCkII5impyyOyzX51Mee0rVWE+
Ft0KpQg31sqZZ9KClH77+wkeyU3lQ/x1YHB++MKyRwy58v3KQ9HW5g4IgrzSZYO3vMd7+aFtxOBF
Nd2aLl5xxTY2aOhd0bOBO+LLCsM+M5++RD6zqjSS57dsUq+v5axE3nboKhjdWWHmmYor+7MEsLKA
D8DetHZo9Fril3cTp9gWzlrti/FVseBsJmm3L/lZ3yPDztVTlQSUdz7Wo4Cgv4AfdxtG37qlfYC5
Q0Ycw6pdrogh0J3TtwUWhi1Cz7/FKWZz0b2Uu3DpycnrA1tCaKCaZl1x05BtbarDWBIcV/GH8FAc
LfDIHLxwsUXhCeijVz/kFao41sHO3kXnqnynwukglTBR5LD/DPGySO/l/HWN7n/++bF2hw2GI6SR
2iFLs2qpK87SQNQM123m1wLbsh04b6ut5fjukoEpgw8uf7Erg6awGbkjKxm8grA8pVKnNVUbmiN9
/F+qlNAI4eX88SmzABBCr3gTVY/gOeHTP5e7KED2ajd/oC+9MWa840H2ifYB81BPMtgkA5U2K11L
2qdYU4MRt4Bf4xPjQMybIyYOoR0EmohsIlLKLvdgxkbRLRo+oBtr+YaX8LFp0w+qRETUcVZrm+vU
ibDdKIWs433TsiYlQg3D3owAkc+9LLckzMkpD/hpFF8tarZtq2dLHV5Rru5tqUZP3ky75zNnbr7m
OQmYLH2Rzz6YNrS5QIrJugqGEahb4Vj1+8Gw9kUiVJQdboXENamFZDDSFA8v5HHHRMJDkW9cr5lf
yAs+SbilEBu+W9vTf1xxqb084SyXYDyZouggJi+7ptkgV/Sp1nLEt0BuJ4FEB9CT5TEjwP4tHQ0X
mg2B3PcM6VTt0V3puhxZzQcW6Ho2o7i0c/0nR8I8rBjZJ5cFe2ujYbqSluAt5677w2jtck4MVlcr
oyq0AWRY6xZG38/WZB9CoHffVsOmFt6txuPEGc/Ha8CXP1ySJVa1SzKNpeZwlQbJdyJDdtwCjjhx
gqmOFqvLbAbVcBWs1qaFzhtvIBmLFSMB9wE4hKmrOFcnv/0SKBYYw8ygijqmzyvd3P3AU7vz2msX
Rkuc0uthuZgeeoWw28HKDvzS/FvQ6in4FSXfuqNfyIIGrxsqulYsziZqaEgrR75uAXQ1emoqgkMS
ggi4B6ybH3GhKrG8IrR09Ian7p259KJWsmGvvVWoDSz8IjvJ6hy5GfRXSbHJbECIwN7IqsClZQBE
Ke1IIdq+YR72d2rcld5AxMCAhAAuZPf5A4+0jhweaInt8bRupsGlY8UnjYR+l5djSWWYg1tBjl5f
zOTLjJelS8/b+xv+OcH6oZSmDUsdtW7crmHDettaMDnkb5P/8Uu9YY/llTSE5X9UhwPwFDal3AOs
iqf/0Tx3jmeJ2PMlqZaTEIc39mVLRGTMszZ6xuFX9Us2tXgtmJCfHSG7+qQI9OxeW+gYZb20lHdV
D/H0cJIM4CLMP1mbu1YweZgLL6lcD5hTX/GydbmXKdb5gEgBTpkVC5vV3FIxzx/cmwCglVrfAqzs
mqfVUecLz7GRNy3XbZgGYerHkqWDPTNtmxPWsBaSBd0M7APkcNW19mhTep3UrBDtx/mxnvhFPwmx
04laY3OzTkvSndNjpQ6zFDXbhsDBsV/DXrR9zTwdrZZoAfMoQ/QH3Xfo0wnaLxHA5NFnOaE/AUkc
4g98guNjnFyfobG25WJl8woOHSzZ6mfhrKfkq1r1U51+oUuz0LRh8j5fbD3ilb+ZFTvqPrzrXTUH
uL456rjNrzqGRHaSuRpCn9RVzd4ZnwuyIHKLhX8iiEqMLAPeybgnT0xvFhztF6U8V1s4CaZyiIrp
RMll0khmnSSwk1nrdF+0AeoVElVKUq1j+s9aHRnZLdH4fTHK0yrBkDADer+wZmo8esZmDiP2vZgW
a8U7A96gUa/ldXKaWj4BLjxFBVB3Wa9T2aXgS8NOXTNI7S2hKIK19R5cgm7SjXCv35jC6z1aCNcI
/IZfbmpLXJs78Ntsi4yTsXxM9HPx4nnDhcdk2RliXr8G7TYjTQhMBaIWr9vyrpaMX9W8XGYaXNcD
6sOq6lBX3D/wGgG7zyTrcsyZge3bnbwLTe//Y+CPH7ovq1O4A5XG3k7P89kk6472kjJ8vVGs01U8
Wgb5lQWFBLZKJjJ/Dr3NdtWBoPWSlhILSiyocYiTEAoJyKzzly5Rhr+dNPNCZhnf13z3Dhy++QZx
B0CDj3c48pqfvtTV28XLvVQ2rtFU0OOtn8wQchTFp/29qHFagS2ESla9xx78KLBGmol23finG05x
IlnHWzza/2BQnrpOLzWj9nKAm6nCdf1S4v1e/b2GYZNspS7RjjBWuThuXS55/BDFXl681cavZ5Oy
bNKNTpqW91NBjeSpQlndbbgO17KAZ3srGyrj8a9u9ivVw09IKL9jdaCNgkQT54yoSBLAoQS0ZAOM
Q1wk71BVih0/j0to0t7/m8Mc2OaiK76GGeU9ix//ravWCFJ4Hra/6qwYgBUKJbwHtGxFtNOJ24xi
Lvd7pc9qiq8Crj7zBcUYmfq7Y2mG+srO89iVkXAQqYgNW+GKMBJazPNdUbiyE8fWDgY/RoJHKfZe
qLPAn9trVeVckaMWGHd4TBvhOAAPp/OBMAUAkPnH7L4IAP7zSv6xZH9JgCCelkzE4oV1c6VyFiIH
Owgp5ku9jTF1gDtn0iv1ry6Kbvp+LFu8OZa3Cr/xzh2QfNCwP3HXYp4QnHTX+lim1qdJqW8Ridhe
7v1wRqJsdfWUkvJkn3UH3yLXmqSm0LOs5DyVUwQ8xEJV1XFPz4b+JcZ6H9unDkyP09HSyTwT5FRE
cLBd8iMlO2cFyzISeg9I8wmMdLL/s4oCucLyiIseH0KSFus7bQlLXwa2lKV7TSfGJt+FsfWJJaq+
Z1PwvQgTPU5hjlyjw5BC3lT5MEgvhUC/ztNBvxlNAc2N0TIrGZnfV4LNoA+WYOcIRNz5ti3oKyhZ
uoBuaETx7AQcAgUUb3p51ruf8EADBK3+RJ0qTwelfDpaAMH0Wp7Dz6OYJ5ptdryyLD13V3rYMcQ8
cifx6E9C1B/S2w5P6sf3GiBasFLvLJOIJOMHMZXzJLlLKv3BS3AvvDGV/7S/caXgm0JJ5pZ619zu
spU3OvgooNmSZNMzcNofppBy+t4VBMGaF0a+lyyJeZzNk4CHPyBdeqj8I1cx5YUzMfrjOvvsfJ0w
j74fxojVf9/S37TJJpCRWCq1PtG0Vwsz7R448Rz5pqgZ9230Vy4nBwA1wOGhAr/PLlMDcUp3iwWt
D9VTQc/nlVg5vTRfdtkWx8jZCZKxKGBa3HuT0toGGGvyc1/7KEIcOb17fpGNCoX8ZQ8bdjXoSoJi
Rw43QTLrc/zgNHAAojtBr9U9MZfmfakGNybaMiAjCQdJxv4Wf4i2hKLVe/F00wqaP3rymca0VDiP
Or86G5XPqHVHfGqcShzR0UCMxpqWJNOu4Y2wEp1snAifNfEQxENs0jwtv4/A8hAa/NsJ6zDOL1Al
A5JmDgXCxN3vkW+eoJHL8tX7sQ76WGGHUezwFZ4EyPEaT/hUH15E7yMhVSjwLJQzzxcESei/ukkN
jc+A6bBOv+kMBvD964k+ESD9zkn8NSOf3ddFpznyLat8GDSTyWZgq7d4cDkGZgwfvMDi4Xd62JZ1
Gz1xA9dQ2gesXSHs/nVHLQUbaqZYKfs1x+8Ct+c7IN71X6XGDRnOWBCpbXCqEmxbJLEJXvWUe/pr
nQy4EyTBV6wJn7uRevdJnWnOJrTUN4a/dQo7+5mBbgy20lLSU+w07IG1npUq3HDXgdnIGvYNGXEx
+tGC5wtNR2MaT5tPgo9cMBnbU2r2eahOI+KlIS1HYg/E/FmwknqIRu01VtiqJypTxbVukPR7CPI5
8mKi1JiHL/wEVjB0EXpXhwKegc1n8olr/1A0wnPOVCgzGRUdJ9nLRL54RFdm4z6Y38okfq1EYy0h
A8MC8gi5p+8kOmfL05E8ULb/vL1pIajuKsxKKyZHRcBDzLKj2in/vteKCIGZcKIgmkjVcLkv1y9J
Al1p543DPPiXQ8hxYvYAw6CFTpqyk1kg7RHU9/XvY3R2UDy+S80MnUw/B94qwIO77wzDxZBcx4OD
WOeae5HTNzcdQrs/b8amMlS1OIZzbz5HHoonEVK6kEBR3cg4RD9WGrM9wiWmTWj+hSGFnotwADVX
1f6mVWPakgMnJgN5IrcZChqUQLx4kxTRdRGQ8aP5AtMB2Lj5nCPBV1xYbe5MVt/XuCT4RXjLBx9M
Avd+GtcjCDoZdJKJqbAJy6Zbmborx08hvmZP3hgJaBXsF07563++xMm20vykIitQDcOhJSjui1p3
WrQHcLb0etsmpulVeW7CewsFm7/91e7YR2ol3ZWozaICJeYPFZtWemMmAZCCKnDkTYCpjywcxFjg
XBAFal5BEuwz6cLKyvCNjM1X7YMK6h3BdaNtkQmHcmbk3aC+hnKZjwXkk3TDun92Q7hzPGKUX4ot
8uKXk/5A7ClCvx3IohpYBx8LbJcxlqzbwCxUBZs4y6JyH4weKUIb5WFYBQ9VLbXfzVy1l2Mb641o
cQaaJf+8x8+bXBnLIAokXj4RgcFQVacgAR/ubuQcU2xB4CtDn++4lrsJo1BG6fUytXvns0CCGiXa
ZFWxw2K0RBFnyhQeaz8w+ecWUB/rBvU54vJE42moS2NiVnDcRuxdt0icGFZAL7/4imlXkxqX/J31
ZYlBRW7rauBk/OfcKu7TxUqvV5tpKPDDmkD+Cb1hVhCJsfdcBXa7U7KGghn/kZl+tP88Jcd6/VLc
A1kOyNtd+Qc666PgtKAzmSOS3jvzXIlZSwmaWWpzh2Tzp7ltM3kiJ2Ezgg2qL5B5vQCASPo55G6P
8ukOV5HiiVjMtt7ntXK9tgIthc7P5dRFuTf/61T75z8TMyPAlI/wI/r/5icBOc6roVrs6h7ZkW6h
Wp+fsscXNB8EXLOtEJ0H48T3O5NhPWZ2/2yN3jhhkXEM2s4osLAg0zDAa1X8+/+puvdwhQPBuGLI
J2lVPGaMP61hzsZcVG7uapfGAEwtiyZcuHIDWxhdzC/fBMDFKQAP6GxK/01m2VGL4CO6QVBxui7H
q2m7LzQFn4rCr6lXXIBHLUO0K8pMxFlvHjJBlvRfBwcWqXbIWqx9SomVG+NYpeBWpiNP6oxcQ4fo
bfv3wOHDqOV8UbKMISx+Y3kIDNG0nwMjcjO6OFizcT94vnBiQjAZ/lsu2moG8OuRJ2Xu2lbvdcuc
3CiMiILSkZ5sYkn6XOFH9cc3U2fRifKdfs2LTMw+Ab3Wq6iiod65QJtAZ+nCCg3yjcGc9o/s4Vbm
nrmxxRrahZpUyI95OVRpDZWQAG7hfchAMU8OFufKPQaI+Sb3IygzPhq2iwhz+0z0xGFU1bqiVcqt
YpudKXZOBmP5d3sgen5j0efWai98VG2Siy50+9xu1GilYWOMDnrkubeTMCJAOmKVnAKxFlDo//aY
zLy3PE0bjV7JRXeNnlkNzZmAJhTtyoCFnD7/9huUJbhmsFH6qKvUIzMPJWZfCITEk9BvKl4u+nOs
aj3gCAzxEHF6dU4G8VwAwwZbNv2Ae9jUGBJ80izqydLsU33xpWrdECoqdQ25pFC4UfxBUPZ/G07A
7O4Y691yUkwgYXPbU+cAaO51sR94ybti8D2/gDhkIyqUkOp21SrtFJe0R2OGwd2Smvbd4XdWSEn4
DDEItLQZB1uuXnFpi7qBcJB3b8LH20vh7TXxYZiMGCky4/GiGTlgiK4RyJ9dm0j48bfdTu9esvaj
jwi5hcCd4MEv3NtAayPl72sLMBptJLd7GMic4weE5ieDxZRkf+EJNJ2eLegsX8/jXLNdvz3XuSIW
d+lDnjl3r8MbxYpTUbqQSKsKJP5kUva8QsnIZS5W3UTUm71ouUnb6quxegBQCAGpHyltxIqapY9m
p7w4Ecnvc7M+7/zI265htaEp6+VIzFcrTbg43OaGbTsDoRSFdGoBw0kiN359oHlSkwxUz1M2lJrd
NlwK6bAaO4AlDKAD6AyeLyyoyZaGtxNwHZq04gB1uU0ovW7dV+9HjGOS1k1H6OwZVtv/c5XrWD0M
t/gkgPgPgWuGYNr97ss75jZE3GVmmQ1P048e24r1tWUo//Wmkbkzf3lp2Ygwzk8m3PSsK2GIOnCp
p4NwZUJ5l0SdD44h3d7oOKu+Y+hhUWshSaFWo9hWa+TMjP0/AKR0UDZWnY2gKnYKfmbSwvX0Nbc+
gN0yGfosYTSWGInoBB6oOaqyeDvjfXNUBko+Ytqzxkfm0QWpWMpV1f81CXsdyhtyrNudGwpZMoZd
HZzxRd/psSoG/zContIDNCPM9Iyk13ccCBY7ee2MB6NgLqDlF+9JhnFj2V6onrY62vhO9bAaVN9A
9Hvi86ldNvcJDWM6NcrylOWRSCzN06T/yX46llJjytmifFXqnXpL/DEIIFXPwnzAvC9+MKHU3fnJ
OoBNNtvAfVYMsA24+LWA+eEEmv5FMmeFm9MpRLmnx7HsNYakHybSLtc9NqljD28oLcOIfhh687EX
sNJadVSnkMiG6v1edlf2ZUIb/Ll90Nh9B7YlmuPIfkSH1kGuClBk8ZLYIDYbuivPVDgrqddxD0Kt
FiuzNkbM/5nN0kpZPoPE306Uqz678MThxhPu0RikKYgemU1JEsvmkjw7GJhqbNLHH/RK8B3JFAe5
dOJ6tLhfh8fPp97D98NmU1XiATpMvfi4uBKyrC8eyfh4j0S3a1MzW9KGpyfL5OwHMZTxoa+FXEJ1
UsFadmYD6RrwftVnJCy4GwY0i0teKA5GzDjcHteZuZmri+efji+rq6HyJQ4zblp+7bOTHUNYng78
h5A9Su4TR8EbI43sQuXdNaJG8EQ58kIYdnqy1aBWAdTJ55P1kHzDpmTUb50MwaFZb+mPaGIS2iu6
uw4K9+GQjjSztlMhjbIUutc20onwId2Nq+MZ4dyXW23G3PKPihvZFfs1kKcHy2ZyRr1Hh1MaHCJR
D0JsU1vdO5qKmtenSAl4Lp2ZldsFfcd9jZsPLFFnf1sQp8gMJiAwy1DY0QVz1Y2KS3siAqk3puqw
ag0ORkm2i+ODgOXXJQs1ch06S+Eo0I2neXL47UYMPkoi8Z9pPWXp2SeYI5xTTNU8leua/T8ye3cG
NGeRWT4NIDi7Dh28WV50d9rE+XJYFt31yiS01duJACR8Xrln07LNi+x4TXhR/OyslTac+T6bu6AU
GLAjKi7fJ1kJUuR/p3hPdGskm/7ivBMfQnxODeAp20m3nChe7/HnWu7p0N875N58Eiro2btTaDoI
kiQOgxTXNQZhIsIJSKjTVI6mYRDwfSEQZkdFa1aAsEVlLSfInEmogjMRnhJab8iAXSSZtsEqlGMy
eOrAzGyOoBu3lfZwZdAT9F/hgUCAuxfFRxdGyne3ImVGahxMDU5vz7JJJCDEYRiYqcSXLr6+XQE3
bPGuHrsMpokuu+km6rooQSHroEUH1mC9fxiPyDk/4lY60EWpp947TO9Fd4D51x52kn7NDYq9I7aT
LezMiWKmV6N+eM+om+vCFS600K520xGt7r5wX4VRJrMdwSWiojxre5c0zPEtOTDn2uH26Inu+x51
sW2J4Gc72A0v/NmYw2ffNFHOoBVjz9geWzmYFE7Ie0qYRWrYOKKkPbhZeC3B6FFeLSqN5Gj9+hJv
4KJS1oPSiM7jbeGZENof63G2a2VLwunI0VnutBE16irdqhJecRSh3DY+sJVYy0faKLwGIoio7FZK
LRC/tYTGewrjxNLVoHFlJRVhVK4A42nzKyI7YDMoXQDnM68WyM8ye90uPLgOA0N/D7T3C3UNhX0A
rL28apA+QAhSmDRfiaP8qjBCAncSAZzIbQi+z2ve6x0EN1xwIaAo64G5WZvEtRhJ+4vBqbcT+WPw
bMU516Wb7kVBUxjau+d1OjN01fp8AWHHfBL99L9pcO6+ubG3cUILSfwfTMAj8WfSGa/PZMAc9JvO
Z3EC3EPVvC75uM56+esErYCGk8E6UjaMBwWs3MxxrwUU+2ys4m8Tj7ufw2kI20xMekIXnqeEDz6o
Lbu40HzzuiQJTdO0RrP7pwqhH6Ne82CxwrLSUE3PZM89DQggf1i7D4Dz2TYARbK0BUOLhYAn4aDP
Mo2vbvKc3A0dkcUie95TrEYwBldD5DimXtA3Wm4gzrdFvAA3MGjFFX7F/u1VAcwW/2E5z0xKtg5O
1fA7NuE1iDVO4oPRdRHnDXvjHwWfwVA5EcOXfei5T13rT7bonDovzzFcMLoSmbZOLeWOZdC4oMfm
GpUYfTQ0Mt8girnnxN5BjOLbjppt7LZWLqCgasDeTgGQXGx/va4om8KXiGD8Mcfj97mr1R927fVz
OzO3Kj0Nhj9WK3Z6YxAsWAnXK6pH3qM6XZcdLjvjB8PGMF3rP+bOkAFP8KwVMfdSNOBzwtjs5MON
T+N2LftfXgVrkzf+IrTv9SH8GVkDLK8XSluTSE9ybLv8t771KNaocSXtPCtV9mdh9n3zLhxTqB23
y/wzYtKqpSlhRYu+bKEmcGpA/XVBppKD0Yx8SYR1ZDYlBJxKObntFKynSqNxmgEyTsAnBUUGzZ5q
1jqd/rJ4K87UdPF1Oj9a8hwNa852jkPYRgF7aLzMygaK87vJ+/POSJq5wTLLvUDoJByz++9u1CvE
XivrhPjua/UHvUWxTuV0l48Js+noNpZ2Kub6xStMnDC+HSDgcuEUk8SLwD25V/T6jT7AXaN14N2g
PrVm3HvStr0hrq0YT/xrQx1BSdwFIrte9/TM6Ig9seb+xyq3bGdem2w4w4lggqoHb9/luvVEYoEW
RYMUEif7nsiT4RR7fnbfX0m75ug+h17SvtebBdO4B6m0Svgaj1lnLh+vdP1sIOUX/SvdkHMPE+dU
ceLRjQ2yatgT55o9zx0KXjVXv8EvT9P5MFvnUWDa8W+VsMXKXZzJTUCstByCNOUacMDPXfO9dj5j
EiwtpaBdREcBW9M3CcLxm2N5sq50NI3S1/mjSFO/CLE75OKAOn+6gKTH99IJWn5lf7StBTzTfAKj
jfrOxQd2BPtFTthdlyKWSJh8s7xPsZkVFJD8jiF3Pf3vZSRRFMXHfrUOq/nu+bOHlXmdU5i6kmX2
OONq1aVUpcV8M3QkSxxCx4fX2/8KzTp6IamqnXWrlNKxWpnrrtCC7xH5tp2DoUi1ejzucD9etcXe
JHObq41pIoBkdjWt5a9Ni9v6S5lZVIKefxRYCIQ4UExCTFk7ubuGeMvwFYTgu515Lrax3UfdYaBc
BLGxnHcGrsIdZ/eoD3VgQjQ0Xoct1L3qW1NJIAUIWQh3AS4v3V35EASGNRgvfMLpVVyzoVMdLkud
hYsYwXpcFaAvW1+5ucRjveoLI1YqAVQsA2uG+ZOwSaBMHd1F8k1lwpcju0wfArEPbalt3n9+529r
d7eDtaqUzXT91ScS3B2FhAij/K3bMVUyYgA88MqgDZ5ySE1I1buglZxBEfob/1JzYamWKuQxdCuB
PrNZYrSLS2RH7BWjr20PjL9rhUxYYvimnh3p3/3udHyCIh15d3rw/+k5fbwpvHjKbP3Qi+U1IGxs
uvB8dUxKAi0e+D6gBhsOPd+/Udp7IeUnmx4XImnfianhD+/eNXKeDase+HpqXz0ppS8ej/r1afEC
6qOGNWH4CgYNu32WXDuayeTzj3KEqkLnLHYptsYZCiJQynyNxP2A3PwvJCl+DeCgjdgWpLd229iZ
dtBrMJg0twSS2CeRFG3948+N1zC/tm+cbUhQJSVmP8TCrJLbiriR8mhTQVwFkErjf9htOsCYmG99
gO+IZ4rgYNtiBmVh83c10W0HoWjRdvtHVZS+2bdssL/DNbotWYyJIeFN+GEbbCl1niJXXj52QoIu
h00RDf31tJfho1TGuqxZNGRu6q4cnxHrH3dUA6uq9w7N6Rm1ot3GY8i/hN7wD+0demBbq8axGOrt
EC6ibuNaeDSBuUuURpxiIyW5oq+VWx1xwU/d/Af9fyI7XBYZJDU45/ZIt24pZYrCLsyukLBx2yDv
1lyhDXuC1gtPQqvGuCgfIJtBLX1IUaDueXw44kEQa5Qk8AYIgHg7tJdBWwufWpQChg3Q08+dK1gB
9pTT1NqsOFlr82iX0crMwgsdb/ug7w0lfG1mTAhuz23U7qHnBLw6/dQ7uvQTUHHmc6XgWfvpvXFV
Cn8YAt1ocMOMGls33c9kv8ThkmxGYv6h7OEPq6gmzzQahdFoq6CesUQqrDtI1OKVlQ7w9Q7jhi8x
eNqEZxJr7dBof8l6sqWq5H6ucZvwvvjj9OGXcB6TWreYQYrL4Psap665bfse91oe+52Bi2+jYsOG
ZkPliiKiP6LBINvasa/Yqh5ZDXiLPHxvHNPZGamM/oSjiidrClcA2dNZ+AQVmVVtL2VRRBjRyyzY
CEUFHHBPVSFxn08V5k/nHL8uCPwX00ZaDwvx6CWFMITHFIPhXGPXvoX6eT2TP7+nDvlqdShicHNi
P4+tIDsAT2xNaTL6EEygn8UZgvVSYMN7Ck7fyfijhzF02/cc7xupJcXsIcTalt6GYSyx1jxe0aeZ
eqnslqlRsuvA9+/jxA676M1EXljJ+bbXCewCPN7ERxbwL3sJsAhNQkQFXCCUw/P14jWvuvMuhpqk
BQn6S4VhW1Uj8avF/AgFLE1zFCOcsQNn7Typl5DaC0ul0gHJO/NJAR+bH5zX0sIkjkDHb89dinNZ
QRjuprvDkmhnRazSAuRjTgSzmF+X1cQM/UMvy7Skm1tH7CEkZ1tONGYOqeoD1AWqvOd5/NfOpq5x
+e3fgp7nz4Wd0uJeiwSxaBX1CNbL+cP/FuwkEF0actV+ykzpSZrcQHAFBDZFpiaRI29MwiE/gz3G
gnCNQtWAyBwtoF0s6xdc9oo5pxtLbCqdSrABgYnUz6eiTIwZUH2OndFQEMkANKHW55K2FRjO/2/e
AOeWdrTJ0nlxjlJS7WQCy8wKFEgWjoMxfTv0iajQAtCw8lOlrO8yaGoivJV6h4l0MX0b49JNvYIP
eO88Y3uuliZxhsdWeQthNDtsdcn6U6jtCmoAqy0R9ZKeSGBt+7aH/3zNy2DdzF9Dnfm1XuTQcI+8
zJXUXwrASyATs72NFeDPkxYMLW07iBQ4wv+Gx8rxYG6/INXbzOETtLbIvGr2MnLNgecvDo7obiVX
8JiWtz37IaHKXC0BQzwuIbnOYKRI4FXDe9dD2ewUffnjrU0CtS1bbmChLT3+J4zxfCvOWhNEpfi0
2O5z7NqWDx+ypDNOnT9xrTF5DVdCI1Mr+GczQWPfVqa+UwM4wzSOo9qxGDsCDFar3Y6jxFQB/PQt
paF/Ltzxf0/gf1x8+BF26x1AHoHaCvcgo6EycVRWhqwJOgRbuu/9uuyrT/G2Hld0dVC1M5VR0ZAK
w2dqpqlyxLC5x4vsn1j8nn6clKh0wDj2Sirkb3SszhnoM141GuQd/BIbSmIPbGUAWK4SnbeFY7na
nbgjkSa609o9gMbPTStHB7OEFdkwrJoi/65Jw/hrVJV+rQbbmy0RUGo/eTow9qoAJ9hhN5g6go3t
jVy+5OUivpzSml+bOEOkLWAxnETWXa32pvIp0zqUCVFLaCcDdGGCiztPZ0oFnATZNsyUp/DLLYyu
GKPviDsDkJAhyCaq2OLpxdKfEHnFIqCYuPC0YQht77G+Uhid1NMLAHGWhv6zFsveBh1d+yPd4cEK
bFwgUAubv9OhuYNrBk37lnO69pu0Zjfnvhd03UoU3YaCX2WNWB/lqWn/nIfyZ6EkE5jOFAzktFGA
32CHyMY69ru5RCCrdIDwObJkgk9ifl3AERpoWUmN0gk9/laZIWUCCzgcKce7nnyDbVeJFAMjWW32
4ZUFRD6Mlj5O0oicCRWujDcq1K7lG7ePzsKkytuiHmCS8xDsOs0dprqCXmV0jNWbGX/eQxLJ8I8O
N3yxFnjkDiH61lyjX0KKNxUXMUOnPAXLvpTFTXQAro6HUz32xy5xCWOWAc3zK31e41OKk+geULr0
kBJ9YktPJvmzUf+rG51Tp77YA+gs7Qa2t8AcGL9EFMoh1DOsEJ+MGYb5hxXmp78eFDsQiaWKI0W1
OzcdODVB55aC/L84OXRVBqg1Khkk2fMZqFyW9aCe+uLavTVJ71IMg7r57c25Fy1Mwij+3kGAD9uW
byHXzK3/AssGeayLvitiGr/qAKbcOSdJ/3tPrtvMiQkwC0z1SP8wvFsl0iJOrShVGAOrw0jlgddE
KqvyNmhzn2ljpF4dnjo5dNk7IE/qdq7BrIs7Sg49HzYyDhE+Ne9UzBiXTtOQRBdrzxRo+iCuicPT
UFz81ZYXdNbWwQoOH/ZXEWiMj3TKvwF4xZVYGQPM5aqVFLn4iOPKceVeQhuaT5Z+dmp1k7JeoUdy
z+4sL4t+WQCVbv5UEsnnKgY3XzLTVDZg5iHRCVwLrL7wHvR0GzyKJVtL17g7c//rnrMIrnT3vvMA
2IaDEWrS8uFJPlUueTBr/nZjc86Qot+mXix7ytyJnpu+rb2sto57f0+iVveZBdJ46t+TehkrL3Q8
hwvGIXpcUWRFU7aei6kQ+OkEY0sJhDRaIddtXTJVO5FxYVhhY1hjCk7S526qwqgH29ire6I9VnB8
ee2fEml9Lom8CQui+kD3mbYhHqqjRCoecgAQspX7nTvVjCvezt3SQk87cjgXSnGlIRPfIYh7PAG3
QPhJfqFQG6Zq7pdvIP1V0axYrvvOFzYhikdoEewNaW4IcnWBcXCE96ZygIpXCgfKTioqqq8RqHZo
h83iZ7POxzhKQDYGdABW99R3TPk9BGdp85arKa/q140JT4yZIaZqmL7VWRiik3264PG2Uu786DZZ
zGkWM8c+On9zPrEIR0JfmX6Wh8WBTlVOLq9BLU7B8MHOpfo+nVxwU9PwnAJ0/FSE0ZHnycX6vcdu
Z10Ej/fm8drOE3xiRU/Jrm+VurVekOtfJOEaeq/qwryNFkuFWeC/oed2pViZprpeYt44lPSTJr5l
fG1GpOiJesEr1avXSOv8Uwam1INv/xJD4+CsNDCySGXATmK2qBjh88QQmo03TBC4dkNLULpXVo8G
ipP/PpErF6wseUw4eaTpOhf0UtlZ7vWQEg4jpZBqFPXS2+/jXOEZiJDPvwjwl7ttjog/wFv2UCzs
Xds+E6HtjsS2zDzRa7pDmsXhFfTM0MN4bO+Kc/s/2krVy5imuPhkyLDOMAQwuqooojjE8H9UgBlQ
jjGrLQPIRgjgNmdG5zHHdj0mlES1dps3eGQLpg/Va1fxYELty/E4/dqxO4J4IAu3rRVEnzZzXIAW
m+fWJ6sU86G1AT3oXklMCjKwu9z0tnKol4CalG5wJY47y1jW9n//FlWcrjP9y+d6UI4A6t+L4yUT
1IdQ3QIWa/7MfLHQPt2jX3hMg0lb1p2nREUHpa3XJHMvbanIE0NYaE/PiJy0fA1uexvDDdNDSbzl
JlkyhtFMApfMP5xd7kmzj+h2t6NfhcKCRs4WQWY2STPjCJ3Bt/mYsAivX+HoPadu2v5eX/P0Cskb
vNuzOizzu2hnrLyPTGEtvFTs/U4Zt5TlSGq4nhzBb6dYnjFlQo3F0J0+UjZWU7I2bzx1vbjcO6an
yoeLNTdoFBKPatfOSuKqLYvHbpWq8yefelfi2SObk4ek7BiQW9BLbezzzDaBvndKn7cfE+h9ffXK
3vbWKYk4WOnVPzpuOlxehegUhvI/AR5FMhF9Ms22SQvRq2zLtQTb4nJZAxSjVXTPbY7ImVwO3ZTC
3NlqyXONcxFeBb93Dk9C769SLXJgu7Ajp6YmHOoG8W/B66aehYHF13buR+AyMl07CCGAaIrj6YwI
+P22ycl3W8MZMgzvB38Ryfwri5lHmHPemRj4vBnHQEOoNVQFhrrILFws2OUU5tiCbzTMfJh1dp/D
2lkxbBpBdxqMx4vDNkRWsw2tSjOCJm5cmeKhFwljw/OeHpFaWpIC+CbqaAC6onaLZ9ZEXHDLJHdc
cbRk2KMXw0pmyTJn0eqreaZj4h4ZMYjY8M7FXYAnGI4qSiKANRo3klD+TwQJAk+QgLDmfBPyGEX3
UI0fHfvc5XBzuDrnSvI3ZJRvb+F1/ciDYCqSYE4myZW+9etQLude+30KGZ9NtBmMRw+6xXMjQFah
G2cxFduKJ1acZIjEbDVQMTPlS9BtdFX8lrcgsV58PwcTPU4WgSL1BoEPTwl/61OlgSqh3IEjA3E0
CFsLfEDKEwfYppqnlQA3s1AEIMYqmqt8GUvozV1zd5/XuEOB/2UyDipVJGV0E03pJEDQsfT3N8xD
ULIgKrwAoVuWjkDHYiymVH3nu2q1yym8QOV4GlrhY9XJVshusrXybB9SYHY3EPFlPbGFSUXSheyz
TkItO/9ZLnnakaSf8Cqv/BsQFkiZcplCRNJoJHGWjUYRnOTbjhEuSPxz8ZaVuDPDU9yfP6iKGUBm
cE9aisdHyzLOsOySGIzosO7YHe35QYM8FjXcQO/fy4Gamiwrd4PZz1w+bif4nlXkLk/A4SgWeT4a
DVgu9lZx/Tco8ujJjnCBkp6FFXrOoYljQkcDX9bR1VQo+jZsNQyWFzeX0EHo6R/f9kkNGsP2Fkp0
EnKr8pzLFc94wCGBDyKwvi72Zq168RhIbI4HjnpTRLwwYH3750T1AKccU5WIX/6iRDUmIq/ouI3C
W4fLBAJ+GtEvO+ssuBvD3fpoo14swi1gYn7TcCEYdIjS43vhr6IRDOrOSkLAHbS8lijpf18srCsx
Cc01saGF7iapuG3Y0ARUUL6JNPjhalxbWLexSWivOQtkRxFCN4S9mmqIaafvNry4tQTj89wOrUuH
L/p28AGszlB645Ib7pHUh0puxUHO9llihRR1QIbtat3cncI+PLOHZFCkBdzhOHHNWlhY1F5SXdYM
dkwjoeqNEsW6ZtX7yj5dELxWRBuMBx23Dw7YSx7UL2cKvZzwUxbaW9MmErEDkGs3CVyamd0y4BA/
0pWH7/xbss8Hpmu2qP2/vc2y7+ab2cwto0cKtfwnONX12LRGEKXT21a66dt3bzEIYx6z35T0t5F7
qsCw4mMYS4ZFIRjzXJDm7si1diddGq/vYimG0aog18BjY1KsL5F0fTyeg//JgYAtsXCex0IjP2pM
WOq+c67m3+zc8Kx5S2/HICwZNMhF+3oA9vIoeFFFc+aFx1ClWBpGnrNUNRIPuQ1hOTduAtFI4bFc
zvM1h6/Rf3rVjsibn4Z2YCbUHymPHJhhmsfOjXoPT7GfSaj2cB8aVrSOAqdBC72L4yoGyLEnMzRP
coGcwpBHOwDmi07cWwCsbolKMLZP9mCQUOirVZwwrRSP8Ocv/ZHygcFX0qbqnK9AKaofwAIBn+Ym
j9IuL3X2O6Xo4WD81ZkqxzEOW0wYj20rwQHO45IcXcikHTD3RPrcHPEtNF15MgeXVNsKEKxttwLP
LYYKyHgJxbYghU32jHWnB7SOiVh9lyRtdynCNRacHlIwkPPqLatP/pRLONUZ6NJwhqU+gyeofycr
torO3STgdwjswQFF0RT5URy/uFs011hTdkhR5WVQxRz3FxbSyjzG/F0JPqG77N4q86W14wtRQWfH
K1j1o63e083cn2rhBvw/lTc1hKtAEmO3RQEsmNzPQfELkznwBJmXCi/gXiwbZ3iu0W6sUiaGVGzu
SS08fOxof2EWFZa3oMnMAfrLQlgDv5KjpG+e7BqPvUTeQpcCYB0V3lLdbzoasXYjiudVw85l5lBs
TDcwK87QN1EtcxLHa30TbpS2DW0KJM/huChU0QtyGtMvRgjVkoF4LLyzO1YP4i61rYZqFKKx1j6n
zI07a+gljhM+Ies3yvXtjJfe9cdgfPD5rPiGTC0EkK286rjTGZ/thNdAVIeN87wkbmW+GBiVbgEh
w6RsN8Md6pM0mzgZqhBowQ3eo9/sIPoPbsuw+OYuZPd+AoGiKw4IK2E627gVata8IrY8vCCeqiNK
VNa155TGdUBoOdzAxxeRPKnQy5Vo2AY1WoIkwEPk3GVIVRa7bZrtLA0FkBNvzmOLi8Jq7sr6n3Bh
Y0MPYiSjh72roCUTSdTfkHMCZj6nLK5xKjV5J7yPFZ5cSxX1aDoXGX9ZdAq409DEfX68wrb34lL7
4/03tj+9jKdoWLiesQkF7DAyBMKu7q+++QWZRhgfkrcLYw4kn0qckVBGOqwgiE95dNaEEfWuLKjw
5lkc68FNGbTQv9ptCzMylwAyQ59W30s9RpoMHaudrBx/kX4Lsifvm3WBLqLlV1pVFYOhbIL1nZ4q
gb+uFeqNgyBdAM6GNYlUzPaXXENvHYor4Sv16qH00w/Ij0ztL5n/HEpGQwkwsXLgyxf6pZxuhm+J
EwZUB7zWv7BazXs21vgKXegGUDSav+sJeMvZ2dlMBkNzDRSsb4Z6jSTVjrXB7h2jXZPx5kzAFxGe
FmEo7Oq6f8VhTqqy3bzQQ+CflNyOh65GPJzTT/c7yqJCpRmpnMdwN01G52lu2ixFXyeKnDq+vXXU
KiPryWCjZTgJHD76IErAIC/t0aGYpjmyp7i3NfZJLo3153TGQ3mk+vXXb5/bgcugCltlj/NsTFuA
Dzz8UCxgrTWfRwqcM2+9fyOk+JmHci4xkalT8r90fCAplFEJPy5zAge//Ht0Opv9DD4JpSiPSlWG
7RW0tBP9wVBeO79OCS9jKFlAOKSkxv9R1yPpYBFhqDe7sG+UOL27+y/hPQ5j4foqQq3jJkaQgn3X
3TXv58o3EpPcfbwfoDmjYelRI/fPEL/9Rp49rQLHFROYxYN/Gxhz9Kdkh46XqagOmFDemrxTDsQg
9XuB0pEuLfcJFhjlv+u2d+ChXBGAuuE8eSiA12+pBU3JYPyq/pciH9HoVlltnEBxQCV+4pAvbf5Z
vO01MYFV4kD6zOe5DrlPiv2XdSq3UTlqHbylH6a941L7jRxlJml+lTk9VNvrw722j/9kO4Qs3IVJ
fKzdgofag0wDJArT7LCAp9y/Ky8Il3lkIs4D8pquiCcxaPPrA0aDiyw1cU8PEOGOuzMg/ARihmOe
4iNJPlhFBog4OkRpHswO8QNZSjn8r4T5XKF7VpQFECc2aqLGxKhxUV6z+j5k1/m58YTcC1o+NMVq
znqr08cAYaEcGHCcPeD5fO5F6smDLZX3KR5M4QP1W+9JBnIiq+2wCGDyqkX7HCMIppklS56cabAT
H5nyGxOMRAUOCGKVs5v6CzyUIzWMLK6imKMZ+mGonhEIYRY38cbP0XvN0pPiwpwxsDCDu8IHa8dX
NxL912/3KzYK8ZL3joZWjS7JnzHw2bkJo49ca7wWs2sOe6+Txb7CooU82XwBqTm7zFsT+74n6WM7
slFj40CFcKIVF9D1eZSxof9cFPFaLbXWD7GywJbvQJDW1LI/7vV9dRT1e+os3yATHsKCq5SzuTz8
EvG9bELeRVGT2y5eVJ1gsChPVBzuQd4QHuOiCKVkBEkcM3swMLIkq2QkFkvIDNwbVuaarsVfOO84
Y2euwSQ5sqfLLsDd5CTDYiavj/MtBMam6F7fcfLplJFjMxP0HjxiG2u4lwzv7/teCYB1qcRth0aJ
DeEtBnY2o+80tR7o58wuVRPs6031tbwpY/+v7Jj70gpQE0CHh7ejclWP5UwKtIOcs7i955Q6DIRH
L1Tpu8ViDaePXgnChp9nT2WQRJjXoHLoSnBHVVnxp/albgw+8Pi1SZH8H/Cz0rOOylS6hs1YLZ1X
+otjjc/v7W85qGboDv1xL/4U2N+16Ok+UCIIjVvml+6DZKiMByt83JS8SJVVECVPgk493i0bZCEz
zG4QYtfQqE2FqXKCQvq0QXquHxJcJ9r+FEx/5WSFVVunE/NlODjZ31nhwuz1OVG0gS7KnhNjnauP
Pc5Bj7rxHyqffWAUYi8cgzyONAthaQZx6Zectn+mE7lRU3AStEcHlu8wUeji9DEO+eerUgG9O9cL
Xvm8EYEm7NlomLbJMwwz/N0uewt29v8zLGpLqyE00HkZIlhKP5t8yqZ4PoQSs8nwlS/RrI808C9s
Wg+X/3rScjBWmZifCM7PHMMed1AyJoBmyjB9GP7uZFB2RI/W1rvwYLUzK9z2kzVC+8bE6qcHepzP
OvL2fAy+ArAfZnKuawipVoC4xuTZF34gvV/BeZYPbpl/DlUVU6HKTC0tk0r9azykuxKRVWH71Ggd
X+q064iwT0Hsj4nX1ev0oWRU8hiisnFOpC/yphujFjH2PZbWMceNCB0NJH+8Pu3ee1nMh0BxwCB1
3xvySsBK4YyG1L6wBsViMFF9FT+L0Kh0hSKSjVDNo63/idU5u2gMp7SuFBK41w44WxrlFTk7MrJW
C2yHCoyFwndy+ffFKxWPJ5cRTG3cXbmjLWc6FrkcmnaJDb4z29HtZIPx1iSvD7tkOfvFLgWEq3OY
enLkvexFIfYcA0YBv6ASjQvJyvVoove0qKMBl06ClRGtGN6L0zONbYRAnpzaemuRgibtw9cDAndE
bh79z4zrUlLw94P6nEvycCKsD+Wvk1ly5PFbRTU/bO6hFDkoh2d7bewYVrtzdfxLiDIntHWMkOYJ
d7vxkQwbb/ik7MBELwJhoS+E0Kxt2Eg5rdkp/85zm48k0/p7q8tBh0TgJR4Lm/noiWR+52TTqHtS
9KHsYOxdUwGYmF8NZYXIc3y/rac2sfzPObvU9D1txsINaN6MlrJI04WfdiMzilSYSSBvWmzPL+fb
2TPJOwB46VMw6PzBxFQ65TW+/ROBRQhTXWZ9U/sJvhLewUwj4GCfHv/XFuH3Cgs26FqXPOxIlqfs
1c051o1/XWaM5QqIv0BNWzEWgWYXaINlrxTA5p3qkxHwmvOO0hHaI1dNHdX6gteE69LaOI1GsQVi
B2wOhji25zy7F/I+plr7xfZNasNpZ7qlkfOKWPEzEOgTKXR78Gzf2Hwqdlzsdjm1adFFxO779PGx
oHsqlQY7h4Gy1lkBoUVyd25OD14tArbdhMQJtovWba16Ifj78UJs3sXqFXh1QOMGhyfQFzaO6ws3
Zf4DcsU2guTh8qnt/7z2yvyoVlY6Mprmvl64mg1vOYe/vjKIW1N319WlS+xu7N3VgwkpPP+9gFd/
S/i+ssIR37OYZ/NUCZKkFMJel5cwZM3Ya8QYWRt+U4+pliIk/RqI/IvHrXkjib2sX/3x8n7WUdTp
612L+Rmt7Eu5MjkKZjPgLiERfdNMw4YSsiZLX4N7JH+wKJ2xNMB3DHAsDHqONmap8gvHKJCBloGH
H6ezMknx4Vr4mVjemZRBndB8RYKNz76tHwzHOBB89N1BQmgVrb4jM/1lLeloHvhj70K4OEQbMsDy
16EtsUeXjsXhK5+JYvy6lA7F76VMBx6b6N8z4VfcHwrmenJaO11P43l7raPXlM6Dm380y4mcW87p
Kbj8BVstRShHW/tUXxtOwPQ1GWApEngGSNKuakuoyMIBhd7ZbM1a1uADaJdMXyH8sFnZpJkITmy3
jeMgqGsHhRHEC5i9c/pj6idtz6P8iseE+e3Iw+T6kNWahCto8hHGu0jBaaP30E1LhXERrrxDsTAe
8C6LXYpiejJEW/7ulE3twYigIHhFLteTcpiH325x8IvfIhocRKWNLpjqIn1VfOZWXVvurT+h++4F
zi6ma0xr7HQlLyo4vAT/KigNpzZsYh86GR+27rCOakqf1M55krM0AbttXkOEB10DM8re1DX0sn4u
P5/TlQR+nklkM1JhlJqT0TqtjsyoNbxnd63Jhz7tj/aQjNbXSFgjwYFghpm6aVpluXjVKowo0xFV
WuBMIPqvbbQON/ScZt0NsisVCP64AX3SsmFUbq0rji7BZ8Hd1Pspf8mVT88X190yaH8XVwaabj1q
b6aBilehHoUHRqMTUmvX0b0RixGi1Kh47Prg25T9D91c34nQN8bBGjjtwkTGIa6AV2ejDI/Hn6Ht
RG6Y5SMVdXvjPRHegs6gXyx2KSwvyx0r963JqRfIfsIRQXsDUs98a85SoTZ70QYg5J07VmDScbdc
KWjT+PMv+ZEhlU3/VWW7L4e++VVe/gkAhYSpvIhLWrPtf+B6CPHwSBmVlP2w+sQ6akAO/CHhf8vU
uY1DRhUnvw3FvdEbKJX9IuM/7VFmwKg5q7U7SOn/D4CBpGnliMPW5WF2xmbbM2lE27uokeq7QhSR
Ap6EX7Niu/mN+4iq9dj5uCtxmqrt6EcBa824Nu4gvw2qoyU/D60EBSVn16cXnrM65dcs0FUWPomC
hzwFZyNcbAuEu0xwNxEp/xOhkWzMqKVCBID/7MpPErCV4LLKA7ncZIjFbBJCuszmZLrgO7TSa4S0
Ih7ZiDAftumJO92K25PK8BqD34lAtUD5atHyrQHOAOa22czTxeCsoK/qzeB+99TGGTrKqUAZcjst
RuG5yk9lrFo1xlCnpszud5Wykf7TwtHhFhzi3dj7RMWGaVxoTb2Gn5jTosty7/1EQJiI21th+8sW
geCNodJ3ruIH6pYrsRXgKj3rI/FTqu+87p66f25FaC76ztMrUgFE9jtki8OpyAQ8MYQY/hTYgl8t
G++l8RipLkcsMRBX6u064+SvnrOhF1l63VNrNOc1CsyIb67Tj2ct2E5rr4QPSlA8wDQ33gACoIzQ
GJO3tK4Gq9JQZI7SBjsmVP8o25CKx58t8z6n4eznFpe48dTquCNzDhXAD5dySyFDlHsuqtRLIFtS
cRiD177HeECN7Eqs0Xa63mpThscaMnY61vw5j7MqT34PISdGTkmoPyl9PR/5VkNaF+R8EA/oB5Zo
Ixx4a4djt44XxuN0WXYGkP6ZLGI5YhbWk8Mg0mXOKHb+irqH2GQaEciPR7iPtgeL/kaPFVa/WTF1
1ksekmCiX11WG/O7aJyR5Orxb2HvfUqW8a8Uwi4aS/mTyK25eN84UIhAthmP+k/hU2TzfZ39YyTG
oW+LDr5zDPHPR2BnsvIbZ7HeBO+zvCVsLa4+qFiL4uztJAGPblohDsWYmhNFkjzI19Y23ZtTJq0l
9cOgqyTqrMlw6mrVRl9TFY4y7tGLTooqEN+Y5qbAwszJFimt9CDpJRzkNZ0OWbzL5oItctGjzqxD
p+riu+R3+BZPNxRsuPFJidJ9tzB6eGsK8rrjDDpio7FvKVrENLTq5dSsQmjidiv9CDHV1mGFf0PE
qpm0YK0iYMtXQ4ueU6aWh+G0bCvqbyetmKdaSKu9ASn5+doD+UPr2PMbwr0UE4yjHUnqv8Wu+wXX
6BaVXfF6uq7pYUZp+ajV+wEK/Qol27YbzJNlvEfJvjiyZogyD7m1/pCMDWwL8hSiYjQt69Zwn5V3
2oTmA3KFbgoP2lgxuFrBatHKsNCY7FXrzyw60iqzWyOPsC8t7UZ8E8arv5qJd1gzIOeUcfvfYv4X
oswy047MtM4VdjArFTthH4o51DcyRBA/ZnD3rxqAy0zmzDnpbhYXqbViUpVOJJoS2bbywAZbruva
+TNW35JkrKx2EJjWrwhqkajpd/BNrV4AHeqw6CkFme811EYRkHxt9FFWllfxbbvjTL/z9VKufNTg
76UcJVuBZR2Eksz+SyVvXxHKmukUMGl1dsjRDPzDG30VzrjBsOemj8A9a+qHRIs+RqMtV//v+IGG
WyFdXcxwrEpB8uVE3lVSgGPCu/9JFhdNI56gaRsAixrTtnv2TyH+CJvVdQQkFWG7qNlX5W5wJGji
6WjRxvoR+apV8lCUpDoYU8xn8b6zvda3m3GramK6A8p23u0VoYq+IukwLWm6gBTB7bUFsXeBdE+f
V3+XmHTLVdS3FapazKmBSVYJ26m6+zIYvGffdw8/PJ92qN54XZJogMVDjvNsJ7tdl4xIIrMp3pls
NkR/t4aGOHOdDLU75M1RFGq85Krd4pWSRLiaHV/wtzsbLSuEPa8VnjoeLhoQgC6QCvk5R0PLlfVl
oUqMnXpJTCU/TRtu3MTuSO2qk+bIYhA26zDxi5wa3nt8pktjMquINoMu05dCT/2FdeJqzSR3YBJI
wDF7ha6YE4MhQLuii9eRgEU3jZljKuSwBUnXmcpEKZjkax0uhXa7IDJ8WLeaD1kZz8BbELRE/utk
kIEnQlTzGZvjv8nQ9sFV3d8ome7CC5g2dClRMHs+FwcvIpmD1AoXf22Ke+/0MtUfHcPGoKDb6n6C
iJ5xpQR8jt2opjzAmp4VhJuXf0C4CfkJ4j+X9waXn3cOaf+yyuxlUNIFTHn8LjqcMs9I2iOF1kyz
u0T0z1+396Rb/n+VZA/eB+/qmNk7nGwvJVXotXanoZ9ZCz1QxS9sTlM8uYryqT+A8QX3EbqVlORG
X6aGPcFD9i1RtbQzJEAaHkQDOUk8B0PqnqhxqoHjRPFoDPW7SQNQaRaEHko6ezgMS0p9iA5C/+RK
OqVxnlaNBK4uzd0Ebx3QPAlGHEM4Ej1MbiQiqm172IqmrawTFvGCW4ksa9kAbVPIGpoiGULiFpvN
meYXtJScp7ny/p7FVsrRohzBoXaFBEH0gw+saE4RhtOyCE2iRZykfAALdAX847S0fEr9jaCHdzwi
BqZTb4HtYPWQvdunwS/OYyQ6YqEXCW6wV2VG/PWrlVOa8gBCuomTE1dbrCl4tFC/lLttDdrRaqwb
R9fcgX5UK2Sbqufktpl10WGPJxGryVya8VGkwjYLXKmPihsLQeJ4LoDFUXsNUy+ap4kDOK3f3WGr
ZfVI0ld7X5WfLC2wLKI/w2Zhiy5QV2VxVDADGxRDcngUHJxQL0lyxNcPmzQYC+zw3N4Or9gqhHd1
ElyKtqN+PH8IY4KT1QPMglCFKjJm9LhN8E+GdqLvHSzTkizPvsjAVCQG4n56eAdeioG2McXDNqwZ
QoyLy+k5g+NsFau7Oc/ZbLDryy4sZr3Fbt8HZU3ZQLc7xDBQ4BNI/x3EB+/kTMRVV94pLwgenH67
UQEX36B2L+q1IGgD1D0Lz02sYmHNlfebdD3YkHHKr73EtfE2q3bTsc/ly8on04Qj9xhV+kQJ4bs3
mXrwbPuboV3dlGB5o0vus15MKbp69FKUVzOKLpmCM9ViBJk6x6n4pT4z5Ykw7qonjMaKUQcpv8VE
U+fFBJuOL5qdoEHuKvj4R5nQcG8M5WxEfIudHTrY5LkeojS+ix6C9BrZPfeK1ep1m0TknAM64KvO
T2Dviuz5xwTtg2djmXkNgUxE3PNmuK3jYKAn8lQAyxHZtoKDruFpcGeI/6NQ7aKmZsz+cShT89TQ
jad8GcTaie5hHQTLKAj1uycTMNzpxoWyJQQeyHyfVaa/0QLS170W0b3/ZA0myPeRsB7ZHMH6+XqJ
iGJ/MSm/prvrCQEPIyXXH/S4K+Ci5jPBM0ZiIijPGbIHVTQXhvCnAjYegoZ5aqKtRccsqbuRTcxk
F6K3z6l5kT00k2wGStlet2+4y3RbAN0aOz6FclKvtQCmh5HdH3fFO2jAqPGaxx3iFVEuCp6FRBDr
exg8yeQWQeAHJ7Y0Y38+mKUar7GbOFH8oekb5ch927odRUJDSyEe5wUjOhj2X6sUR9QvoD8gDAyC
6PAcqLWNXFUEeSkhb8Zg6W+Kxrk0P6Wwpz0VQC2MUjD35yM1zaPaeQzGq4mECjGyD48mp5VcU2CY
UT4pWjKwrli+St/ggBX5AVm9Y17QxYh4maRvmhUn8sbRk09tsoy0fDpji4QZY1iFBleJA+bphLe/
fnnNFVwvRhHQs8yhXg06br9LIHUj1cXL89H1GFZ9eM6jjZPXrHlZqxN15GYUJClMW6mspezBXhe2
J5haB4vvXUahqyZtTCL6CspzQ/iwYYSOZvi5kDlPbg23K1nqSQt+l8QvBnBqqXNcNHMkU3Vpl8MU
bkUwsJyX0YBeJm81AjOaLc+0opV1Lw+LjrrUGNjSAthzgh1ARiJiWsMJAJktVcNR2OoBDqE6QrpO
TNYFFiaoKpbgXyYX4sIrqQb/bH7mp6oXvfrXN2mG1oWUrXaNZGeh3YnBkzV78h7uoeyHraZLPdUe
ZoxEMXEkimAZjg4nkGSVTiNhiTgI9itrh2LsI6gzti6bT4YniNwsAetm4EG9uqSafMYpcDALDN1G
iC/dnPmkCdu4TMPDR41sc/ukO7vFcvq9JVZCPxPIqX0aENVO36UkfxW7rytK92mNGIvzlokPmaO7
GIT/9t/zxCVX/JkqTxk6pO7r+IkPAsMYNqvOkGOgzojqxmToxxDs2vvIDoEily+yDh2pulukp8o6
6H5R2MItGk5prJVvbbOrkL7wN6Jbi9PAqC6V12tzKLFlqVyxwPE40bE1h6U6kOmhLi+ZS2rEO1lq
qztNZYpMoESIvooOgcTFW7/V0YQIEnoGz5n/gmKDqhCYaWFWU1UbJPFvO+h5vwW6zrpSN7jT6K9S
h8FBv4oOsxQE0zZRzyI84gH9XuRrm97cDYqzm6B4+p0nhIx+qxN6g+OkdTQpltspybCEczxqjg2f
4OqwK/w+2M3cyQip/wr7SJEQCynxppgnxv96dLnCx5MwYff6enMztG/5Mv34NnpJeGCFvWDzC6R8
kGVT8zw9AdB0WrFWtgUkG4cH0ZEg0nPFDPNGDX5zkTlFMJUTaEfB6u3WMKdaRfKe/9pfYnNZP/sq
btosroGt5NTM2GIX9uywkUQpjBoDw5s9zdx6y+iVkLvHwwn5bUlPcAbownbFhSAfhpBQVUGmrr8m
xUjOtRVW1287mNDAWGKeq387YB8iHhLX/LpNqV/qIb8bsZYdcabE3HflIASPYy0JcsXtWDmd1QIE
MoavwzUFZmzPlHLFBgsVOsZx8kP/gYSk6hxJ06oprowkMdpxV3gb3aw/Q8A4nZuZRXPpXYJIN9QY
Sb03df5FCPtHcWkFBB+EfNc8QW9fQy99plIydj6M/dQOh3ydYNtx0RXxV22qVfpaIX3ZTe74NUSC
8WzqSGzGD8gT6zErxKBb8wuuqvJi1iNHVg7kQu6KPIssS+CP/C5nTNvV2O4O5sUeSxgeNpahqcnJ
4WFG4wga+Y6qySNdLqGBvAVRfNwT3BWWQDgOpS5WNOhZcusZQGpbc8kadssTL26FS7QV49SKp27F
zNR1xIZf8S7Y9GDZj0sVsq/PkS5zQOwvXSZT2lb3hWIYN5LmaWqhYiiT+q4bnldyovdF+0riqpOu
cARBkNbspxaOUU4Ke2lqaFRZXe0cYyL5eh1TUQP64E3aCM0ENQPt1HHDwh5kPQkZ2iyZReZBwM+b
kAaawwOAxA0l2tZPMSQ8/bvFSHedtudeaAoF/mB28zFSx6F222oobJVu9ZAR4gQdvOboIRDRK8Gt
wyiFFRuxP8f5rMus4Ytfc6j/v8jMNp1QJM/JZoMXvU2ZDMz47EMEtQ8VbupEJWNXwzbVrYr3M7sb
XQ/VIzyWNrNy4kP49QjhfZW0aw91tYHiPSOroavNKQEhiFOdkG7dNayunxjHw8tqQ1+fdHUe/XKb
I3mpdG7RH+60rp2j4oo4R+SZa6196rRS8mFVueWRG4EhXyPjPhIoorf21IGTQnoIJOtuLYPkDkKn
U5yu4jBGsCbf8OT9K0oIM1gd4/Iv0mlly8TfXIiTCd9NjklYA22fvQMeP2JwdhLtFT+D80pPbbRp
xBYQna51gw6tTYbrf7kVYKqHpO0otc7bP6y1oOyYabDcm+521swUV6plpsoTnU16HNFVFmSJyhSp
gAokasVeCMRpwAtR9Rf7koNFFAbpgXnSuuZC6BlLarZJ/ymz6iVIPsK0sYgwAic/gVSno2u7gDW3
H5ikCxGXpdYwflNWUe8pxWNv284wxpKybJ0ZlSTKVtIpJmenz/+WUb5f5mHoPUCDTkUBGK6acvFJ
OrFBnef3cIL90meQis9CXb+l6NBVTSQw8P+KaKnBygshCDJpeRKaJUJffKsUGmmb3p2ojvMW9hcH
C4jVPxaGHYuMhoIR73dzBsrusn/MJfI9FcDqmXMPhexXzKKqTWEvCNeATU58CrMKTb/evh7Ftsc+
2tzDrNIVac3JIzty1LvTgOFyWO7R0ZCN4Xk4aFLayRaPO5f15NHHTO7Qup3luH+omVZRJ71jyTe2
fVqmeEIRcELzewRsd0AVzPR0NyvXkd9Q52C1TIO2E4MpNqn3VydwQ65UrPkzwSPMokFTPsxEVIlE
Y3j/7uvylvsiKF+zTIWzBSSuF3l4aNU6uMi3F61rdkwXvQkzAvJA+ixH/nVS3aVQ7iJvmRACA1ZT
fFSviWj8mJmUZYQpkgc5UJc4qnhpYzJzitt5d9ZeEsRoJN8B0at/OZohwvBMYyQV32ZN1M27knNF
+nQL/skzIBUjbkNCjOENr2wl430z+6179FzO9TyTXuUVRl3Dqr7pTwIGdrJR4uafMuWsznRksZrM
71uthMZXv8hxM64xo4KjzPsUx3KWAmlm18aQGcEpAwei8yqMgSiXvE4Ap86BqYJHDXlgoGPl2sFF
y0wIUNLlirYupt+oxZeeY2sRtj6n2nxrl7BtB1yJsRVxhpy6f7FF6/wOsjANZC0Kp3AUhU62fKgc
4rmfgatWv3F/D7//ItJe4twBMQ0gnUxmNcVW1D+M43euq6EowMsxl2uYL+Os8nq52CTDf4SrEDpE
ChHxnn/LuvVahBv6q9ei4c8duO1eI0cw03LqXRP0/aqF0YyJSNUD7mCtgFLXxv9h/Z9kiS/W5hr7
Wtgz1uaRJHDscUgcvnqmlLEHYphFqEBowDI6HubC/rt3cstSvAh4eu6E6n1t+ZGG9lkiTE+T7TGf
Gzud7RXxwZaaffk9NGr2S2fzvPD3rsZH1PHVNgP8qAuLSO8qkwbKbnJ2sRhluOZwA1csIobEcrdV
OhUpa8S6JuapBd1tdiEjLq7UHwuH2rpt4qDyR/jYyunFqDe30GaNNSY20qwsibo0XSdZq3cu4psk
DtTL85A6nM8dQT6YHO5mxwAc95VWzagM+5Bi5EaJUuVVLJKmYZ3ZexG/8arCouUZQYvA1NWQziGs
HtTRWqzp7ex2W6a9qrKGPj9cJWia1GkPkBIG0hbKLmOHF0vNEifImxcL4brdpPjGdXn4ouccqPDU
mzpiTI4khl1oWvrSzBG7rjEgRWFNzUEGxbdMSTZIcZad0KA6TbpY7or76FpjZDCT4ctMLqLsTGnR
kPju/1v5HVsbLoiOkv8gA1bMF5m6yEUssmeRn2gIx0z//aKKocbmJSovwnX6sghLVd6HV7LLAJFa
UHNk7/IbBrHhtiUcwcDi+/RLKr/OxzyCzKeSJ02Ch4sS2IgCfymBqwUTaSGMhQZmjfVyBFEqOjaV
nH7JBSmZ2zqcxavWsaTvhQTcQB+sH9mdrylfh/0iWZvaZ+6LKYvFc5No1ABvvjnTJkiowLQwuyLw
aEkWgamw83xoKrW+dp4SSE2ZwkTUSVrBsM11OOzpCdUgh7mIdkWR6Hamoi1Tyu6ttEvVdQ3o11pn
i/NJI42ugLoIQZOwsOibbFpUSU7mB3Nk3jkF+jFJ3kAGH5G22k9q2jwd6jm9hLIIx+dANWJr+an7
Fs+HzwrXZ7yFpJPIdkICPnoGNkHSHz2LdJJUhFJvjRLVij2YvJO+bWYZ71oNNBzMIgGtdaGOu5TN
s8H0vEmDlgBW6jsFzjcPrhKptLQVF/gexwUrPDuQS+3nh44Az7f19/5IyqHKXMHpA223etMp+w70
Kc5v26mubjDZ9AObJ791y4KP+EVZ6STrUcW+mnSYoxbfHl4YVcBJji0E7FOsXYto0i+y7vxGunBW
ONMaecIeQfzRsTUiB07zXLUnpdW9sk34Owq8We0fdQMSGy5gy8HTDhjpg+xRiBEb4lVY8fTmFBek
BLY4nYYjFkdOMI9KcMVum2ieCA4NlMMLF3BuJC0sQqIABGp5rlybTYfwFw5RRMcrMMIXVqp9kfbx
JiVlzA5CH6GVnVJzgzW4YuFn/RrOOplqFfAXXOAvLT1ae4cXJAfZFCVY8aZwKWdWzwplaXg7pGd/
Dw1RayySaOan9nFvf9nMJx7OrYTpvVDiMZ5ZYGiE9UOPag11jFWehyAJK+cEYUs0qLdLz5aSTEdG
USb3hUCmmS904XPoGyFGxhO0jheluXQyJr2Fc1VMtr352IY13CdJXERlWdnUPut3OzUXRwdPtezV
fR9dPcSz7Am5WF0lH+lpJOesIki2plkFiqPxs6GTq/+6sE2SeilfBdnPHmQOBV3QcUShkU02JJ4D
O34Vv14xqE4j5iLlETywIHO/8OMZ9DmmP8N1xaw/IyfrN2bDZYJqXDkMvkA2JRrEyygKJW94mkui
XnM8GRbOrR9bQ9hCP+MWiMPsEddKBc7s1WHuw6UhtQFZCfe+YZsKRNmHJsASSok/exiVkHXg9vtl
JnSkO3zWWLPQOO7RkAuwiChkhnTevRJdUsL/n4bOS7NarKWU3O3y84OwxedR66yOCV4iEItgHDon
XJ8mSV0Zl54Z3ARG3qoG3pY0FZwwiqGMKYg1U3+SbO5N9ezeU8u2jesxM8Xs/JQxqNLFm/1Uy0Km
4tFy2GUdIuCiL53sUyc9QVq0KgZTr0h0WcjF2IUyDokhw+d6G0LpdcGe2PoR/vFk7RwM9Zlu7BZv
8pu7Co1O+JiedvTF+buoMJ2UADOCLOb/3Zsix5uBYnV9oZ8yurMOo3VO4TgcDeHEn2Dvvo/AYwau
hFyyNiusMVf1dnBrEn1sWkuq8jJiCNlM8lGalnMxhGePlWI7ltHINf/euuGkeB7vCoVDauYDcnhR
ICv4TTsoANhPLenSfxi4cT29slBdz4Y8XJ9qqvlli3axdP8AJH0BfYKK7riEpT5YIh1HnW2S97Tl
5lgHykHhuonSvCaSSIs9++dC6CPUrXP2HyhTE2bfzuBryshrNGa3jqdZ8G0D/1WjY1wCEvJ50YkM
UFwcb3cPBjzy7s1CLr3+Uyl6kOo7+J+2bgA2LMDTFAdz3i+xh1IMIvlQZPWraNW2cBUMk1oE2fTJ
VjgTYjOSGRLV1KlLDq6uxSy73gvOLyg6FSOXtPv4zd2pfSSHrFOt9Nf7m4ggAqId2YQu79r62rOO
GNm5k2nU3jGZLscBK+duHxZXvJOL5eEW9buBNlixIQ1ytt+mtAc/NS/1JHBjqlTXOOJgl7jjmfoo
YiYEULUUWQv+V53STAqe0rg4ofgDfvLph6zlQkdu+EfdhzF6nWR5UbecUVTWAqHsk3/mSfxtQnAH
+sg3YPQ4JCXE1mxL7rDLsMs4AscByutm2oQwngig5NrDkysdxcShupsqSyUkFUvUHvKPURR5aQwj
s6axcPeFFUPM8plw1Tx3ytCW9HXl3CVpIYP70YC+OBawPTuK2TTGKNpU2fAs/Sk2zbsPBh7aVxr4
oZ3csiTJo+mMEQFXox2R6H3Z9ibrTJAS+vhocXqvgwxLBfDPIsQBN/RzS0YOz45q3NQZA8exyp0e
ABkl20Gyf3DNN6U/9LYc4ItBqHelocImQh/X+HRrzA9DY2PvximC6rg3qkVzxA9pdsVkVO7av7oh
8Wy3ImLGyZ7zcqnx5Zroo71j8idOXMQCc6SdHLYPe3/oO8EtqSlVozgYiQxFLS30ERqMdAI8aZtN
wzQIkUVhLRTtZCpfohpoyxGo7jDpIsFIQvFkq7JZ/bT3ia/GL0tV18OOGsNpeWJXefDa9Vt/GmEe
8UTn2sg+4Iu7ciFnWAXgr2JTzvrsxx/2Lc1nAHvoKe/NkZp1809ixye7ZQ2SUvfH9wkkwPvu7UnN
vjPaG1kpW4J1ObTBbqHLeijZJY4rwB1W5Mzw4bYMY1fCp0GkGgcO5BN4gKy/0/chiL9NFTeSEMRW
OTWnt/0rjRjrX7qZs15MwMkq0r+loJeAkwdpMbeCvbkLhp0chxf5rw3OwDg1dKSjxxAye4OWJSTK
iB7gLlFm69aUO4iHs4e0GoX7X3GWETnOeD0XRzW3pRZSRxUcbql8q6hWaoT/A+L5IyZhZDB7e6sw
aZfJMGgwz2mlgDLPZjZ2qzfNNg6FSbZ5l861hL8OUlG5yLbjLtGh3Ll6X6DbQ9PD9Fq9US6CsraN
X01ZFlK69WDrxb4tytfb9VLkp6eIKahBfX4vPalooaoGIhQQJVUEWf6dU9lnuFh5C/V/0EMFFHWs
8JTD9kKOBYAZVOvo7WkWogfMq9GjgwsmvIggDcUkYLVveb4f3ZiulgPYJKXAy07izipAd8PlkfKT
7yTL8py3B5lJvKTl3YskALdsLCFqSZ724XzpplEhjEHYqCSlVb5EG3FaLW/g9lrsoIG3dSDNxBi3
eypxVvAyAGHyV5tRCO6S3inWngdZRrSxnERruOBSm37i62jQSh+DNiRUrJLN/myR7GuJmg6dcFZ7
kT6DFmWAagkq2ssg6ro6TZf0Tb6Qq7mKzDN4oafWAZLEYQapJM++YoLpWRgZGIjP8ayeqbNeokVi
jZyg/Re0/c8KrGqSGxxHxC72LLPqun8EX/FiTK049TiYJdnJuVix/ZmFlmg1ihUAxLkJVhxZW2WC
u4zG2oQIbS3gnnvUlkkl8/+t7MJi+C5UNeCL9DaKkeI0UmxC4oezVA7noA5g6N5HjSnECCR8J8HM
JWETOYVoUttAUMGXcTqUH3H5vIs1vZgrl4ihDSsJT5Jy4+ku9PB1y6/KDVZOYN4kXB2/QUElzDV0
r75AeYU8kSlWNIlwxRZi1Xbh9SnOA6HYodn2db1PTBpJhpqXrrL3lrFNEyPpyL/UMhDmut1bVHYY
uQJzfB8x/ehVFJpf/EwXbs8rkuE08jkD/flq3Jnv7+ROYTAUE0fR/S7Py+UWXoS2f/+st6qwrFwH
/V9pQqmFRTuiVQ2g+7LKpE6++YQ9JUREs2bagcIF/SvX+0EdvgEkXYm55ujllSwTkD/gWvidqXEg
Ee79aefcp54UE0Cq9pF/a0o02pOPOmHatzti6Pr/PKUXhZI6bKPNtOWYzklGHy1sMMsv/QNQe14N
H4Tm4GGtVC5dvyS8LIrWOWx1eq6GwTAiQZEEJtctpkEQyEtBLK93LptIzZ2DWAeAiHemS0fs469e
gIP6FwxGVSGylOR3VtNZ1+WWHfZ/r+RSkfLPxAbZQktwUPR6HXMritZC74OgPH8uVjPUjGggQcdZ
w22FZ/fBy1/iiz6uPnwBNm0ztXzYrHBW04ujcJygbbby1EdQbukKwnrLJW+u+4PUcDOgZtEINZr1
ofJ55QBrMrDDHBM5h3i9KNJ5YYuB7G4jYxdKGqgvcfUwcY/VcXcPkzIOWbCt2m31+JjRCCQ9eN7i
0a9UFEoT1vUhMurN63PSGcXXua4NVjVh1x1QvZN3XUmGoFLmpyFLkJBxvsjRtrUpoZNn8roKb2wo
SArpwJLr0cxAKg+kqNCG6Ql3nqcKHw/UBQd70OrElYV3JLQYe7MU1fJnts9thE82UdLfG4ssNMbo
mdf3iZfzTtwBHkGMygyrdqLz3oqoXlI2q1nY/ODFCjUDLvqn6lLnZA6tzgxchPCLcPanUTquQ2U1
cmOonmA9l0Vwt2odK14OQPJ6eF57SK66YiJIUp6rISsu58fetCx1Df3fFVLkTYOC0T+LrcKtWDHB
Vj5kuGZB/jxI9kjTixGmmkkVKb/F1Q9ACIpTef061orwo2IejmT9YhENc2NUtWvzEwFIDqd3B/r8
V4nyaxA/n+erHPjyvjFHZWBlt66yhWtJUWYXA0UrbSy+e2nvbGw0CYglGRmtO+kXK9qwaD+7Wfbq
zP5oww+ek8icWDDHLwiifGXU2rxRHQNOuDnEfgAIAzKxHedFBaGEHq6ClyJBb/7B4p5m1s0WYvYQ
m933MICPa+8ZdmxF820aUmeheEvBE7y/scKsZX/wU5BtyXRwi2S4HFLpQVF5NMydpDLEu/ruV1jf
zq6t+Xy81ZTm51GHomyCWG0JmtgyyfHw2DcGlZ1ekqRF4LM+4z7KVYhl43sxnrXBkOekaxM6CJLK
5x8lcRYDsbD2Tty/JcRxP4fWkOk7J3jZ2iRjLLh/XbLHx1Jv6pVX1zbk9BpxxMpocERqZyjkHdSq
adws1449mYsifB/E37Q8EkYulDWgjLxS8seN+Yq7fgwRrlG8xJCRYwtp3NhwSOb+Bbpy4xyZp8dZ
QCRwrs4YeF8yT9XotgfAHveuQONO6dnO3IiXhqq7j5GtkK8A/fCBZjpjXdlcB9VV4FbylCXgBWqM
ync08y2av4/0/nFrl/YHCOXapshB5yElbwd60N4N8GjrbCNeBruAfOxlQf49fh0Ed0SIXl9GEb4n
yPZwn00dgyLgAR3lvbcWUfrMFqL4sYlYaf8HlWWh1RkBAfscbfOdLbhYz4OH0pOWPV+QOWh67MkS
cepuI14Z8gAOivtfzBpOjsFMnukLTb6R6Pt+fIFgVAN7S3xJnDPEnlV0KIxxvT5BJ0zM7CmtQOuG
pcSY/6qxQFdt4oX0YkSiefPlxWO/fEXpzErpGMoiIlVyTH8wzbmckVCwki9zMwKvo33nZPn2q8BJ
+XN/1mVnPIt8OrIFEBt+8P2Fsz6h9DHh9h74O7+14VNZgQx+Rop16QDFk/K7dn+cgrvIchQV4Kp5
kACDLKvsyRhkdTVdVkSNW9zXOUq+tpSyI+kNScqHglUv9eYk8a7mlK6nEumryTcDzClozs+8I3m2
4JFwi7zX97jazjebpL3PWonbuMLVg9rxhtw6+yut/NMOif7guMkdawQR8lQUy0xtNt26yD8RoOAK
m3Fhfd1rIZFg8Rnmqw9X+I0o6dbm2WQIUVmUqsB8PgtKGk86ZqQWceBvQ1MsMc6PM5Z+QkV93A1U
WRICvSKCNF27BrhdqsrqDBvVP6ZUNzu9LcUCyI2u18ie6TvS1oudMgCp7Vqgtt2jgfrUmr3GOT51
yn8/efAaWb9Q8t7njxJ2rqlIQ9jOMGghzGfFZm0W5s13JBu0HfCyg4CepkveQV38Q7TlMgidYVax
vqj25SaD2lt/BS8yXK7UQxu1ryYi/RHXHoSMsPEV817RkbdNLhvqPH+A0hQmK8I2kPEZWlXiDXVK
R8kx7sihH4mzEfLEP3Wdqfw5uRhKJRRmk5fNTIiBTh50IMLbLLMfus7m9AAixGVZ1qyhc+rb9oeB
w2v8hZrVcpQXe2+pMiYE1UQayZCx9KzAt6LiZKIXejQeZbewNtwIp/Pbp4binROvFNqOrUF6KgaY
aSyXz3UdNbc+LewjVr6UHF+TIETyWFcV570yMHu7uMHB3wWj7b1725UlBiosuzdaoEGPkZKbzxkk
/B8sH76eGhyikASCnac7t/AdlnSdx0CCPrBwpu4pjAjFsKzciMtRf+Xr99Njg/0MXzpF63q8hTX8
izaOMPitHxILkw1o/J+aQSEgw3+2sZmtLF88/8aNc7PXkmgAMyMDpYgpPB2cFjO7BbrdW5mTIpeG
PfJ/pPdqZK+jemCPBF1uZrkLy+lFLuHwQ26QPHXQSMzJpTofwFinfB5ePbK/rcY5XFJnY0FEWPL1
ci2Zcc+WgNopjyBIo4AK5U1VJ0AqQT/Olg+iIG4IbAVCxOi9OIHpZwyc4EudlzE4nlujeGvWsh2u
2XisP4Xc9Q7B2Tn8DblXiRazgQO8Yu7IXkKXi2fq/RMNW4yn3FyOdp2bCffzRh/rkoX+IeXzEED2
7C55jJAlFQO6L9FBNIFKoy3msj57QXQ6fMv/+nsZhXq1Zuiyk4qP98JfoFvadH1VBnxALTNwZHWr
OTkQCEgTBHunUiKCeCaLT5CedwXHY78Diuori2gwwPgX6ULzJ51ST0reme6m8mKzLS1TEseX8qj7
3ZTtWCOzpyLS7zLeQj/upWEVCU4jZDSAAQfRYVDGHulg5pY7v7VfjJ/kqAXHm3n+z2G2I6usd9dP
5mawRYA6DHxnNCKhWiYKlFQNgb9sh50FrBeGE+Ud+492WDB3R1/H5RcD9WkVDMXDeS8re9xeKArl
pXf+iINFM04WukLX89SDPD9gqtz4sfq4nqGPYEua0LhNp/OuRix/Z+1hhGU/HBS4p+lR2RmzFjfM
cwLe/sALDRQceVNlUzK/8wAcNdqFAMjDBnfNiKSm9fHf9csjt8epX9O4xDTj4nvIGW1hNFhL1FZ+
qESnVysQa3XKVEppzxx8L61K9Ktr3EPm4xMWfFZCtZKKCfZ+2F1UMEZinGJMSFPOL0P64UWNwW3f
jpGmShq06yTyl6kE3cZ4rkPMwuXGWM/iA9G9oLZiRXwkJAWq1YqfvMgo85RuUFyHylzItw5VU0qq
Cokun3lO9C32ys8zKccOJgS/J0XD4sd6sGiGNORRTh+cR3oX099mwDXpcsBxgBoLMFa3YSWxSytb
evGMT4Q9eKk04HvvlNj7wlPZ7EArnNzM+r51I/xqte+2CHMOkLTZ/lGrOZfy3CNd8YQ2inVDbFvZ
iOwFLQLcuGoN7QhPQtiPmDpKEe3KA4ApqAdTwenNzECo8DZA05muXVyTy/Sv2/eASjoVkUZXyCGo
e/hlwMlIw0QQNroRT9VU4H6yVeS3Kw38G+Qsv6TM5L75Tew3sWsyB5LcVoaqwuD5o2fzRgMvGuXF
Ql9eJS/cF1SK/1bM0be8lPXcycYruDN9qCe9Q2s/EwQSBqTIMdUCeJ4nnQ2drJI24QmvQQPCdUtG
PbGnN6kCIX0gjyr6u73bTq+30If2+o4zxTfUPGMyZcZMJsdxDAjxIThtbKBGLQTtjZd8QPEUsy/3
jf3eNfsIUpx3hs5dBdXYzLR3teMD6qiMnXaTCjCHSGg8K8avUaoDEtprvSPMighDkmZgI4gLLTyg
oX0bqo2nPoSzin/UTyD6sGf4AU/9x6700ba5LP+WSQFJR5EVNdI+k2VXD1YCn50p89XBXp27Oz8W
xb1u4YpAiSItlML19M2fKOvk9Vujtwb6w9e7+eCl+JPkZlp7IY3KycZMQlL2wvhVMCZXrX1rWWDk
XRjchIAL2m0kDC1HyAMbrJaA1p9VSA1WIJah+IemceUJtoTXl6og6QNnKaxP2cfvXvlB1Gcc474F
UY0PH+afzrJTDLzZRYH4/IpnCdk34uSt380xpks3veDqcxC4Lk40RUo1UiseLQvI0dwuNTmdDS4C
QzpiAYBEQGYLzanbmDePCu7qHtY3myPa6/oE8kTVqVClmVVvqfHvo/Vm1MqseI55ixV0i6ihrkr0
hh8kGxZWGX3tP7nWK18azRCutbsht2KPTvVm84orRCupfBPuzvvK/W3BJ3e422R8UbldLJo0Wmgj
z7UmmJrSSPgBnMI5s6k+f3g0oQH/w2oRz4LIBezBAXg/iLCtdvFBPgm/Oce3sTK0zrOQQhGWxni5
/8PIb0v00/Ej5bJSqsGzQkueaIm5NCRvwiA0unkDao5rRCHPKf2oWkXcMmjzkx9O7Ijax9+nYav/
BpgK25cz4BAC4GKQaDCzFUnQFmDid1smP+EZqxoARB738U5oD0rhJvD8R+1YUHM2vXaA01zDM7hd
sRcZNcA7ovYzKGPWeioi1IwnZ6KkEpQc9gcjST4/DGuxg1rHHTmDFsZDD5pZJcLKqeBj9TYqg8LC
adkpyFXSeUjHX/JLzMtcZUuURFLniCs0Pv5WZquAuYHUr89gHpDsgcXSSwMF0oqjO8XKvdNeDcCR
Fgq4bgv8kpiB1WKXCl+8rI9DCESMmyeaUBF1WWG6AkUo3LoGQaWmU/hbZhxauLItQr1OyqE3hZTU
uZpcSnf4SmRFnLkCH2qqqu1phq92xQv5swp2ppKdV9R/0iGPXQf0ti3Z/AaGfPLW6dZQ4k64mWdR
E7H5W+zAywNKKtGN3tHjNQ/22DgGH+BD3vejLUTQr4m5gy4PhI4U61XZfBP0fC8sQ+5yCehddS5h
Lr6Q45iSarzpAPOQJSgWuETOwQww6swLU0nd2407FxQBBsEONluP0SWYGHupTeZyTHbfQA98UkBX
a9GjdPjbqfquK0asmW6Yyi8eLWtKXVSA/aP1mrkLeRItFt2s876ebAM8FepapKQnM1xYyZWRFJnP
iZaDfVsgj+gl5UxOzwpbTDTfPfkoSpwA8Pk7Non0ntyFJWTXlXEeZ03tOug9uz1r7CQka43iG+l4
ZhuUgJ12l8Jzo8AvWCDIz9V5uuEsilVcH9N/CI7ZmJ1Ob/AA3EYTz7WcQVANFkl70a6w1i9GIwOa
pe344xV4DKWfAq+aR/ZTFCRkhdbj0qIje+RiE4cygmlI1txp4rfoPf2C0uts/qwjAdpWaGf7msh2
edcYdf7Y4t95Zo11uKG6K4vDiYK41cjPo085BIC8O7uslSOExQi7ZA3hv2JrtZFg9kRZvk+aiVDw
5VyuXTsuZoZkQA8nS3vUE7iyXdavmS0X1rM/lflFPhEDZ+TxSCaFwMkXNSHM9+hUJeBpPycsxPA5
zQYPE2nFkyNzAIydu87LYwvClwi7+Y3RdQ2mQ3SXbXSGi2Lf4x9r38H/Zq9OVXz6RIWl8tKgU97z
Uqo643Fh7qrFJ3hUP7aXkYMlhDLfj8gs8qkqT34RPCtXhz/PmuIm4eO875M9dU5TNWafkzRqYuqc
BpK40m5I0M3teFX2cw50mJKn+DdAuDk/hUXefIxMANnCD1Da6Qo7AWGZaTskIGGu3+raHZg2JO8E
gk24OgSY0ARQ5cPCrXdSQkHlRaZrLFFz4EXvNs/gHncqBRhN12LrM66WRxpXLPtszzaWTBWJ0Dkp
Qwdfu2kBQZcboe1zMSO6iiAgBBi9oB2A7qEjatsWFZOAx9fbP9njJhPa1e88FC1TSQ4Fm6ovFdCG
7yYaZA1qXRKUa38EAjjAd0K6NIR/mD6KCHlc8RbSdxvTf6eiQAciFBv52TxLBvZYrZGH22nXO1tN
52PCogRZMTnTjEHuEU+slipPYmM4NRzm1vHgR+wio7Bc685gtjMvIxEtuH0TRp1jej76+vFbTr0P
AKwkouKq9wS2ii5pYm/hY97c3woz4b2lUsB1uIUnlYwsTqNO1CKD+74PZz3TPw9In5q2VE125NfN
QcElccjYQ8YVahDKKa9i09iHMV8oTDerc8s70tHahkLGaCPB2Av4pJSNEr5FAvnaWljxAl7WBSww
CdlqxLxghohlpPat2Nhks/ak7ocMHAQSNCu9E+pHPR+as65QUAFQ7LVdmUhnLvGJxVa3M02Ufgv8
Os4XRqkiWGFgII809f9YwP0s2rJGUZZHoyWvUZL/TjZv00i0el/B7nNDLu9KYoGwVuZ/oR/6UAww
nFTcXgHzFkdSwqBkiEw7+dJFlP7BMnS3NsZoMDZrAnylnE134KH4bCPQrL7aMqPNmaL9WSwTV0Qu
nrZk0kakzMI/PHO5VnDsyUnPXXrXHVe2090/73BNrqTrB6JP858FM8uP2+P0qWqJgMojvojTcMyL
ao/KDVjuKgjFZQB0yhaBvLTCBaMbwX3jj/W/s9eOW1x/HPFhjGnR5BnTvAcDSsSlGZbXyVZjXwPz
nRnRZq6bOenPZ8Q7bZijCoRCq38MVCC6PKeZCAABApwlUaaYIxHj5jUX1fykeabwLJv31qP/fPo8
4YU6Vr6SSTvLEeRvolZ1gc9ghJXi9TC1cZSoYeC2M40F/jZ//nQO/DB428MmlVoZ1d+SzLeYaVyh
H8lHnlAIm9KhkU/rjRBuFSfd0WN4Bo/gBXFS0MCPzGGvhsdiAD1wzaFA95HY2L96FFTN3fURr2nF
VRQKBjW8xpZzxMB2uLIUnE0NZKW0rIpewo2wW6JokT+gZiSXCG3e1Qul4WPmpxQec1zA1uEoOeNq
eaWN21j0UbsOSKHrKdkW0vqv8lY7UAyBbnSuvCGS+fBqZL+bl53QDM+rPw4NXrVwSMdfE5awEcjp
0WFlGCCQZBv0/slkqK9IoTMvosofgAlq8lZcRFJXFij3Zn+L5O1eFg95qO3wMMnkt/r12WvYOBFy
K+RJmL2n01HncFOnVPtnYmXlqFHi9KiXdhtSvFVYnfkcHd17VtdMcbfWnyHGAo/WlaIqv75cfX+t
wFu8Zd5/Ck5986Ge/bd1Nop99Hkm+Y29dzMlw3dfiBDLDdvfWaPB99ogE1EWgByh9NeGhKhzkGYZ
fE8D079oKHLACMFASrubaLTHmXmLWhK0OR5bkJXyZIi/YCQRsyEwxx8HY3G9vaGla0kT1fCjlj/b
HSXpHgPoW3WhjL5Nr4/IsMgyT3YFuFB9uX4dYcICwNT8bwog6eCXBP+dGRXqYvMtWWnkUyuAdkOf
snoLIWY7pTiOgKj8HBbT/fAg+U3nd/DEN86ML8Eirqm9CLrZKIHy8p9gIiOUHIRJpEAxEV/13S9U
L+9thz10NYogYSK5tJnb8msk5wPBcyrqtiqsdm8P2Hop+NyirN7gRsDcgoKaUB/KGlVsvwG4Mu7b
NK0GWkH5YhEOLkkjRybNfWQpryEedpYQCGL+y5zkXJuveGsRIKAqG1WD+6brpwbcEgSP6vVnrOqp
ZSTELxDA/MH698J+s3lW6dXAELaSE5XfDZ0OI8x1QgKUuIU2Y9+Xve8qlYQmSyWcr+U0HVNH9TKa
jPOF8ct3uy+HkMHaQ38MoNLpDSu3v6n9PvSSIRmtBszMmxObI1PBNGbe/zsRjJK4gOOTcfZZGSSc
Y5o0Se1M2IochHnnYTGGvHgqqTmo8EL0UvkOHYsE3GC0+FHSNZzhHW69jXC9ARHi77e1p67m2FLP
rTqiqXhucAQIc6M4yp9RyrIRtGJCUvyYPNxK1eXvTIX3/wU4oAv4ht/24IWMV3TCm7l4bQqluth1
7O6JA5bfABXNNYDYbwN+od7MNdIYz69eEd1HiNS0RMNyeg63QqhNaETcs1UDQ+TNzz5Sw0Gw1mCU
HDZWFpIMKHu8WrhewW8H3C+1JxvoOyQ6lXm0y1SnOsbV8cQ8HLg7SKjGGx7lYuWWU+CzpXPnN4Dl
jAEdzhluS56Ceo67eHc7ElgEtE+ctSRRaDRHos8ygHheFDXBmmQ8LLTCahrBYSFI82zP62sfsJ9k
OGis4ZfLS5JckE/+4iODWrt3/1RZY/ZAm8wiTxuFf8PS4y6mUDudFVioseZUJllfpiXFAHcYY/nF
87Meu2qlEsWGK8tFa34maIH3SAntBHPAbxR5gi8wi6XHbIViMdRKQe680YLj00ZPnVjDJpNV6+Wp
c13VFda9UjXVWIG5TyQS9IQ+lyUUA4sG3Z60VMqIBlaVwcgZ6UcXn0cyJkfTqKBp150iPZ9MKjeG
dKIfY1dcB29MBj1dyhwxQeyN4H9DxI58Zpc16Y/VWDdDKwpajej3rVLJdnM+7r2IX3x9ZEdPIoSV
ueGwRg2er+6tVgp75J7nfrnh7TZrEwe+g8nfUPfBU4imgCeK3+twPiqzyvZSVz0D22A+CQPEIxso
gyC7EmF9d2gwhSAyXxEZW/8oSBWbwZHrrcj+JtLrPgbl4jcSgijZrsxiakIPenfi/4lXWE+sPAwr
xYs4COzMvmFoaGrwWQmPUBB+JxEmNqF1YmvCOHMPcps9O+jtX6ASqOFJbC/XjgnLPkzrKW8tnvL/
7B3TEEdXlyFAgAw1ZD/9dF03eFktgUfU/RbwRttzfOVfsjrJWfDTkm97YZcW+EP0Wz9WSkz+lVFP
1IpK2emFXd0dL/BMVioIQQHnnwbvZSdSTjPcQndgHDtbZ5ztYS1h/7VcTS4/aHQHN7OD2z0B3z84
iO2iGlGXofULS5QHzRN82njaxNSEwv8XbOkp/WVlXX8wwHJW3pNfoFRRj3QwKpUhlf3sazfeq3ny
eX3CFX3NlLtBYsz9l9KNpMdaooy5Yeudj8Sf08NoMhXDfLLg/hm79COLIVG+mseepgDO9RngNo08
mU3iqUribZJMFj46GG/ZrHc+VXcqZWemFOUK1Ji11Avdd7HgIx4nzrNHFI1VDfhnPCU8eSHbyeDI
VuKJZyvvcPkr5J/mzcf61kGFg5PcXT91KxOcDMlBe410+lYIg/RvsbnMLHUDjvJ6DMvai4g1rNQM
JDAcDh+0PQO7JpwN2BhUsmM1Oyx13Nk0+rpLB9qxh1CztS8d/wGM2pkes/UxIHr45nfsntkV1AkQ
R07I6znjBQmWJeIRtuc31j5bs/pSDtE4A2e5MVGH9kt1jQivqHeYfgxi1ali4/XWxcJHSS1KdzhX
VViDtyQtrCWvDxuQTnM8puhlz5Wor1vqgr7Wd4E+Onswa5+BZ9I4blFWJWgxCn+k4WsBEzZ4q2P+
RmiatsDlyHlT6MEMw15TQI/3kI6HFO2IrFiMOPqOzOSQk0tF5o5XwQtI0lMWHxvIpdNUuxejI5DB
Kxdx9BDm+Q/sC5hfXseIgeZVDQ2pHadnEtMtDzg6+uEy5k8N372T8HllcIoPtGvabxWVLKrFLSZq
BMx2Qd6fSyX/394ApfzjKLqKturPWtVT0HBjTKZw+J0YrpH81RJO+kwsrbL6U+lRmEKb6OMTe9uw
0Cpfz800TTObFjwzG5jon7jU6QfzMQeT3OZyi8FE75a0mg0KurNA1VYRYbZx3y5OIIrm5fOy9Act
t/6HIX1svmxSt1sLxA3HjP1LtpGuZNrxXzj1dlHaZxWscYJ/D+MSnd6tWt59K1vW7mDJzUcNa4Ow
yASTOtPWT4+3/sW6AdXyM9dQDBN9Rl/ldmoIgCAck6OlUN1b07mBglVCqp8Y07pRNxqy/wZwSxFt
JHzql7p1q9y5W0YYEpfXEXoy+vKgOj9OYfl1hzq2zv5e0vh/Xmvy8PwyyWcQ2Ot8QaC7bHZmtvuk
JKeOXJRTzgp0SfYZ/sUaPNchXGDRENBllAGXWaFYEm6LAV55QE5HdVWfPWQl/OYPM8u9UuG0C5AY
/qS8jhPBNIeBhz76Uo0vKeb5BsBvkwKsqd9BBVO3mOVbGMJZuAg8eZ71ExghyFcVpZqffIaFNSj1
uqzW4winhqwxkYbIZ8rYNZhHpdilFmkgFRkB5SSfWoB9pUxrdCMj105UZXiioIFL5R6l5LVi4bon
1R4XvQD5awTSuCquGhJGHFsPDB+Iq/SafMj8Cp45QePYsTWGNBuFiC18VPhpY6YEi8UHZ2b3H/8f
uZa9++bIYYf9mL2WHn40o15RmdQoTNCkKBVvuGigiExKp51X2YbtaDz7t1sBX+B6/AsmcRwZQkER
HRbqqtrTwtkizXZdVKhQtm3k75eWVAoKeV8Yi+ouKr0H5U63c7WqiZ9APdfKWA6RKIaLgXrdrTL6
GzA2e80sVjot4nMVe4t/KLYo3bSN/QVB+U+td+1+ccqnDwKbjHcLgl3O8P1x1fTs5r3ucmAArRuz
zaZRf+r2yzEtPCabqI0dzQLlhmvD1rsAkfVro7QsQMo1kIR0QGNTqDi90ObMgm8bSTyhyymJttvV
JTNOZ9n7JOYV1dZ3PnlnRLmZWcfYmDuGHQw+aW+1QmeIgjuaI+tnWtw0pzW0ACtZnc8ag/Ad+q8Y
8eHBeLEHrOq4W5ZxYsTSgHiMGnaP0fskRoMjvsL7qiGqqCEcgrSeQAXa847CKu71V+1Q0xVTgTnw
eZLsO9YBBc8hM77A2rPmLKOnRRRDhdwe0n4t97aJaHefJgSskTvFSMwRkMsEsG8FdRkvA+ItHdlC
O3eki2M2YS03o1fid/QKzMjE9edFZ502VghR1/mUKvvQ71fTme//fGx8fSz3yg2h2iEm0F3r5OdQ
Z8ILfTZt5VD7ZecXXAGJ89rfUKbLPKF/QS/b7p1tfWcV+Y2uLhAGtT9Y0mAfJsrHVUzpFUp0GGaR
b9bI0TlKp5tdoS6JTg/zMm5HUxNwrPrtwBFJFcoRbH4AwGoXDuHU/5vQy6JgBsIqbxMMKUHC86Qm
yKbGTVEvdJSxlZcdmLyq2xPcSGrwk+jvrFjKjyyRxH+JbUZmrGVEIhx8cQJzD7luOEeKHj5kMaIq
WbAVZsaY4NRU5WSPNDTdvkJA+JRRVmF5g/aRI34a3QOuzMr4vOHhLNqz+C3bVWvP7RJcyTWJ8vyr
ir4HnT3duGvBc7UvxZX55zFblIfD9TvBUUj0Ff5V+S9//ZJi8Uy0cmhqRPN/rGH3zBzFz8Uq+kWI
X93yiqR90DXO4SOBcmyV0sheEmlfo4zL1hcfnjl8X+sQmskfjClAZLfF0XAIna5jqYRpcf2o3ksD
Oo16MR4GEWSxUPNrHWlOrysVSoHjA+bdNz8gEA7DxU/ZFupGURNEonsooRMF9BMfKQcElKhXyvcA
B5kLv3dupF4o6PGmWUKQ28QZx8k7DtR4KAOnbje4DmCDh3P3SMRtY3xdE4jCwJNOevr2NYpDoEjG
gleg8ti8zXPvC048K4WqwNYodrvqrF8LMijbEbDNtt+RhRCFrbOrE8tnTGu4Vy1MjjFJhaxdZlZo
dktmsNV2dwLdtLLfwuTc0Lo4NYL3jzIent6BN37UBQTwHb0n1RtuQZlLXvJD6wAuKHzUTXbJYqhD
hBo1DWV5BqEmATXHbRLlWD5zvfwPXW4GQANU9A8Ip3t91OrkKAJRCX36L2McAIv199N2h6JtAW1/
KN9BTC8fLL9VH0Ly1X0t7BM68rQ5pLossvnOaSD9mMEKCi6e+LOcwIUH9tQuyWB2Vzj6VlQLafXM
A55BnjilMFSaYq0V25Z3aRNMVI9HEu0IoGW9OAFbK4BZUJmrlYi53XUJjELD+vLIQpWZMTg/eq7k
IZy3GKz8FnudAzuSIrp1Y4WepITPUemwHLJZiaMd1fE5NZss155SgwA8VdItxdWGW8dKr2bxkOLz
hBDO55LTBlf4pYovXXZ0REa6Fr570ImFzIjlcwNRRrXwCSrQej99zNdITJv7AnQmoQffiiXjofy9
1QmAs8SFJbQjUDups1wRr1yoNRqTPfeInDosB0ykmR2TWfrEGqbT9LLiMyuOAVtq0ZVyQfks2E4T
rh6BDdL6h94vgdYCWE1K/nRXcmfJI4zVKTz24erX3RV9kjKNy+GHabetV0gUlU0ApjvKvjO4DIn8
hgR2Ew/QKXNStV0ksde/yKpjk4JDHiw8f8DNFuocz3oq6B3BDZbAfwPWhbShX964YsK7wDpgqk3j
o4mDgCY/iYkP/YZ3QL5oX/bgQ09OUEjp7Ln/GzOsba9B2ewRpvNL0NnR+34nhjOZRkVxEH/ABW+U
9xBYQBqpzsARoc0gFmln3qkv3Kh3UdR2OpnLAEtFUMsLA/ZmtX40iyA0RzDAkadGYQQc7K4pnZyh
AtOLX9fyXpogxArzSIalTPgKC64h2H3luGB3jcxhKDK6fEF6wcgvS+aV83VgzPk24CKl3K5hUTlH
mkthzAxFXMmuNhyNybydVw3wbt29thDKfPm2WzC771qag5N4s+F37Z6cv5q1JuUcrdfxITnleum9
X3Y+0vnNTDbY91vR2L4N6gL3O16ilF3tVAcoBEqsCO1AY0DtbY/WmOIyHBE11+T3hi9TBELjI4zx
NC5bpMDF5jpUX74ivhgg6js57UOY4ChLqEfpy3BJt/hCCC7Fzm0Ajj0/Y+yyQNhxuw9E/iNMki2E
930aErziWywtGNnhNvj6ceI27v5MrVmhIZujZK8pg7S6xxJS1jhbX8q64M/0e8cTfzvuSYId3YJ+
F/5Ax9Yvi104ru9hftKrNKpa0bY5jYphjxQYz7qjMi0uHjAALeYsvmwD7bVjSDOcpyP5dgJsKlLU
NhVllIpScgtZiiKdMJQCByCwutFCTdqPKU0lUAwwJbHh8eKFNOiU1qJKH1Hl78QzpqxD+xUobtaT
BMnpdLAGMnFHclfNrpYsxGBeagbwzME3kk/hxQDmGd+GMC1TXsF02fFDtgjjnQDGnFzOLkngokBS
mRbirqjusyn7DcZaqQU/57c+LFIMncAiNa1IEPd+yMQMBDhao/Ghxfg0HD/jLu3d3hP06zz0Q9qC
oFG/DM1cSiBbdIXZmBcOr3jbkRCxspmUerQNzSxUl5a6O/88yqYmALQ0jN6y5ESFprOIU7enYwuB
qDnQwRSOdSRlwwEIMwR22z+xtgp1et/BIoTbxFu3gD25cc+CqrAgY1Df+UNi9UEc56fGpjokQMnc
GWdlVH8NLNqfVxgR/QBTiRDVnk4G376obaWwQlszehxEwarXYcrtC4jkWTf53/wjjo6kdohudZIz
fxG/Ho5jRQnsh6IljDXb124wHm1+uvFnYx7/uRG5GskgC6jLZ27sVjecXG85LeD0dwQwSc/q9aOm
6LUrLJg+RXzUypHX8Yb96bUrkabqFRhk7cuXNr2aDsACiJDeDWWVv2WnDdLkJ2Dsd9xhcT1tozO9
QmNLG00Md/ecR8K7Ivl7MGRHUaW/JFcQ+gaW/jBlD+P/Dqu3J0G1P2VreAMeeXZDrScUwnS7skus
GkLg+BN+kNSlqb33O5qukjQr6s7T0Yi7INqrVoScEhZYMj8RQwBG0edRKn/6TZJPXFnkpdML60vh
kqbCmEpmK6dDRozuRdmXLrCW11iplV/BI8FP3a8nXtbOzHt23RCB7YtnykUNxEUf/w/Gyu9vn7YG
tYnX19I0c4ujz4m1Ycqn4MmourZm+0bs+J/C6AFu4CivNwRJmnuFp3qmMExM90Mbl5ntzsZqXeB8
rMrRBmA6zeWzP+BdNQ43/g6ojPlHNsOJCwOZyQuQjhGSbbSCjnWR7g55angGJe6fzYTAHzHvrVjU
pQjTIsx9h2mI5COp0D0uUgZY+l9Xirq/LURwralB3qxtt2ML7rLnWPDhdsNQSgFVWZ+ZSQrjuAd1
4NKBbsMxMcXWqKRgBeWqW6dI6G1psHU2KsLXKB5MEPT3rD0Nahth3Rc2RuNplvyy1as1PwESM0ca
OVK50vJ+4t7nU1YFyYf0SH91UiOrJrexDCmOwbdhWsCwRguy1bbMGn7AU5PNw5YFazFU4V+3lqwF
VEy7PrSYzyuCB+tghKOr9t2RByOPfhps9745djpqkkS6uNI7V9/JDm5oRCdSMwkjmWdARxMcX4UU
iSBcmoyb4TgAwO84rQgeADKWlYktlQt9o/T1aZ0yFdj4REy8H75ecwxC67erjRA3uxIkaeoIQvA1
xQVSo3MBWZ8inLjf6iy5LfujS7p5Kw53UX0d81hxvecilYAlYw+eow2hahCFkHtnlTocOJj9pkDM
U1IbItXTanaFESuvgYzhcpO5bDDBfbuLxiRqxlCSEDldbN/ym+hW7wVj92dFAT9xYPULmdUFtd9D
f0w1kSU7M0NcDWBmdTHZ0TCxf4mSTuFV09K2YZRlNK2qkvcDItulk9SkDzGrltsH5pGhMIH5YUhU
YoUDYllwbgtiRLBElwrWWrEaWPgqiPJ8S5osYIEhSnaKrV+6tpqM2TPCeFi8o+Fde9a1dVKJ1Efu
89LWbi6Ve0C0AvcfbyZB/9BRYFmmMRZvLp/D5q5eULJU2a0wkFw5wATXuz7D1VMS7lDo5Bzaqwkh
ntnX/PdKEK7HJN87dEX4Frq3W43j7UfOySq4A7SnoFglk0sipP7TnXqtPRZKNgVoRyjce8AF2MUf
p0y361zwbI21kPipsX4kbA4LBHeuSKSJxsFVhiEhniT1pxlXcGd8R3ztGhTPyLn+VPHPwRJg8l3U
VFKo9TS/2PU0Q5+HBTXGiSCzrqgQOyfXYqtnivULyZ+Q2QQC8iMTkPqCuD4gX0EKU34diHyG0CC7
uRIFKjOo8b0NHZsWNryOMkCxNx6kVoLAinfhj3/zEqDiiXnSg++JMT8neS9EFyS7cuqQmfdAozxR
YXFCDjkOtTtPiCbPW/9mKdQrNwDOCBSwlE/gpanbYJ1T6DNOfXazE6oR5ndcJ3EQG3s22CxCGd/0
YSeCrRKkjhM80GLJJGmVI1fKyp7jF4Uo4kracOwMHCSTPZpiHRWcE8g71hJsMyC97UGFCKMLxGRl
8NhYua4zfoaW4mJUNGArd+0gD0398mETxv5IPLSKCsL1VgMmMWtbSCCTdA9FCgaaXiWXd6JJ7GyS
7cdJ6pwSTFTrLIVE/uqiN6S2eGhc5HwVHLgl+QiwcPU/4ktvV9tFiOm1qIj+Xatm8If+VIsQHSd6
pEOFg2+E5WVqSotOajpWibyKBtCEoupx6Lo9FszpLjUhCdzsrVLHOrLHEHQxmgfp6ua9ympf6SjO
vXkZ8pfdUtCMgkuG5evnlNeKIxjypArgHoUlVDy+eb0tj4+ZVNpeXF6NhoaSicZwBgo8foxNTxDb
WR2p7YJ47JNwgMBDOtft2j0A64upZNILkwrjG3CgkAD1P5Y1UlWKZd9XaUfWp7JoPLYzRnQ8uXWZ
vNVhx1qlenf80Gt7U9eOKffKLaa4wqXRCRzV6kgwPR5lbIojNemtDDS7q4U+PQl3dQkq8ebZ6Nrl
0xu+CBWWP1Oupcwf1Kjm7ezbjHxKYvwVkTFBtDHNWlbFSNvsImDxkx3ulCkgWio5NLwlKSTDNH82
xeVv9pwRg+tKl65m7P7gcvA4qmBzdcqIermziXNG/ajwPLpNIlBANG5ZdxkrUG6jdY1tcg6CUGdL
DZH9n7u7vJXU1Y7qRRy77tgGzk3jdsHifVfmVEWyR520j5ZJu+eltMkwN3K0lUweq9ff/xA3Ll0d
i+KkzWmmY28FCLJff2/wFVUtIiN2nvTmQPU8Q+4GBWliut8T/n4yUb5tK0P/YZAS1/JW3YFNy6ew
BgUZtW8KGqyw4BZuMlMrJi4IVxcbFB6GOhAewVgaeWWcRJ7IvcI9s4rIOqmR4GBRCYO6basuecu4
NAyP+a8in4rOfyMUqBLo2tMbjks535RKc8mU+6Y8hSGEcVE8OdAacwxYeOvHzotb5PAsGHcm2wbN
hN63XqhO0WkHpz+0odaeYnW0KdvfVo+bkvlD36LMkh4WkwMyK9X1Dx8Zh1aezfNpoeX5mfLAaNdu
SSVkR+ycAcfJMyK+AnyT1/AXP7oLzJQatSuc4nCL1N6hghQr5F3/LfmYNDRn77PEBkMaFxkXCArm
7FI1owsD0NMVhJNEWD951VcGinAXzxszQyevkHcwRza6dZhq11ssfKny4S0/jTNeGqVojD9erC9q
TQbkcfF62STRSjRizefa+A0WbsV329oJedEmbchafJYw/+2J2jx8X/Y0Z+ed44tjn/5ndMnpWSvt
T/JURlfs2bR0EHFLsKC0YtYncM3R7TwamvdTiTywYRZN3+Y7/VZtu9ZrXhsIIykpjzeuH2aAPhEX
DKtwiu798rg3aYc5owHqj9E5EXA7hb/I8PgbMSknqZsVW00ngNSvfyouaxErmwZD/GiJHwwP/nFT
4ejN/FffILJBE1CI7DPjsHAqJYZSPnp5R83vhPXwnP8Ry4zwvJsWc5lJmwgBsvThYeVv1tYNY5Bd
AgA2XLl6PLW3fJsXVbucbFXudDCh56HiIxpQ70DiulkHoqXTzov4Cp+d1OHUE98Dve9OaWVqR6Id
zKnzB9F7CjfoSn696kNLaH7/9RoSlnbMIvjNy9S7QJfXTLzRXd6/ZW7nHzSA/N8wkc0j2rnJnIIL
W6AR52URuKg0733OD1sm4TmG72hZBs2gzGxl8EJPs/htZFyXoWT5mb1iH0MlNZ3z5Ivj4/asG6s4
Gtb7DeGK+JrnPYYhuC8I6GSlRuZcffGef99jw1YyvAuk3KmBahfmPpJPBpOEBaefnzOz0lYS8/s8
24IkPh4AuUjK1gCcfqIWdozwfSx3fFVMGk6CDnthTEtS751yK8oIrOn8nhzshDA9uPtKvbH5xOHf
3S+midKCReGibMeBsmILpxFab5Krx2n4mZ8UPa3CzTm47l2G/8UKVutOF8DUYq5wlFmK+NSMS/kP
VIXM0OA+HoHbZt3TjEV2eU2c1hnIZ+E7VcjNZ8lXlHd2Z38YcRAUdYPaJwEDWHux74kY8qJShWIG
Dv9sCg6UedAB4Vw5D4B9pcjnqO8OnyLqK/D6PpafOrH/4KLMvufWnEPVPV3HAnYeAVz5IwoFVyhq
J1w05AA2X61bB9VLzK8AIzo1dtkdNBZ0AVNPHDtWHThatNjb+VTBgO1JMFugmMSg6uCUGypyI2wL
Oc/VYDmPiINdLErkxJtJiZQaiJEJJ3uAsBJVWDfMsL1ItIAv5eZpgrLsxxto9ozqIwl1KfMQJnDX
L+hRStzPors57Qn2ZCYpU4s8aHlxPff9mOYdBR4rJXGBuXTiWZtUo7Zn7IXI7/WxTVyJrdHdeZb9
jMoPxXABmDeSD4hJHxhVyK+Qpgey9JffiydzmXX25J+2w2gEhmHrosLaYcnP7qryaoUYEYbInpID
y0h2FF5ziIsZoArPtwO3505srkC6ahE+5q6WjwbuvvMbk/LWAPwX6bweXyBS55jUrA1vLCV6gMdZ
aMRv6zzXIogjkMt3o5hTmJ+lLuxWxhb/1j82aBOvQ7DplOFDjBuTBWu0/Iyf1kyLoVnzYJ6unmlL
CCeIip7BbD+U0wsA3LyU7LQaqlB+dBsRJTs3Ol4dwsaXLtu9Lku39m6sKgHVBGClRtcwyG5YkgS0
qbYe8khyqmNYKQ6XpcXePCYuUSInlvgNJuu3gl9jOf+RFQqSKqx97bIOE6gYwy2/4f15gc6AIACn
MlW11euc2YZdWvA0fDDXfVv0WiUSPAQPXNMtvDAthH/9turLUAxzEEEHnDiBClf2+ZAg+YIPseWt
thjCvyDhba8+6v+DQLHCAy+UPOfONlkwokaDK7j2Ti+jw/l1SWMXqut7plP8mrmoG63NgJXcOahg
DbgFw0u43mlKznIM8S6RFsuqOCWuQLvtmfJZB1Sh+qEeE0epOshfehbf0bES3UD0c88WQfDVsCXq
3Qw4QpUmmk/5+O2XEJVa8CuMz2mmptb8iRre6Wpu13VSFeiPJ3EefBx86g16TrLeKUaoamKT0JwT
1RQRv3qJKCa9IsFmIE9pKrEH5UlghFP2NzK5o4ayDC6ENyVZsUUszbT9w2WMdoJcLuVeHZwIhkyh
uIHYwCFt/2yqRNYx1I8ZT+ETSZD1OKn9K+Glf77K3scN+YySHHHgX2SHSBUwNY9JYnYcRiDK8PPe
vnJg6FKPM71t2SrBD/zND6RgldKaJ/Xp3CvWf4oMiemjEuVCWVu+CqaDCPj5mkFihYSRzpa02PFA
GssMH8ij30JErr0xs80usAUPI+cz0+lClvikx2BHV9m+CO1425rRcYoqH/5bRy4kPNCxOUjnZznw
lowxA7tjPRzL5VQeh4ZHH46rKe42/ln76k+G17oKumrV4RYMARANbW/6bCRY1eGxpxAiPEsEgIoC
Ep4suIbjTAsd9zAklRNWZx3Ac6zwknGuxZcsyYXSveiQAN7EBRtgouaWiN7n/V3ZW+4GL/jm5Uym
6LNvvlT5aggUce7kDSKsTB3bADcx6y0fEvWbn92KthK2x4Z81xUJ2yzUO7vjKuwuTLvGUGIJ/ziP
jQiNhk1MTp9hgWridl3E2ixYJThbKCMAsXQsxjcOpYhITP0DWLtz/gj/C3lwQKDdx5kFd3/YZg29
/f8UlXBQtu/gh/FmXXZ0C3cWEmQM5M9bDwxgP/hH+p4qVSS/f5wRIpk9eUZPgS7HOfPTfqRdMwiZ
p+apEfYKzMzX7W5ZMqkU7GiLOQ0gRedDz67DzmWQBjtGQQE4+n0a03eTLr2oF6GRF1mekyD1qL6i
2u840sc/V+NrwbffjSxfwcd/xLqCB7kNuX71LkF2lXKmWiXPNeWFnqDsQn+7FBHryHThlFTtLH5k
p+jCmGWZh/Zwd5b0qYoi1rwk6geaJISftDG1Nyja4ynA8ClnXZr8HH8JKA6hEF3k3YtlccCkgMuM
e+1XG8Cig5d3DVkU+1cSntKOama8hN/8SjA8tuETPvyZaJlH/SVrP/1mQu88M0EPhfyYhV49XZb9
Xizhg24aT6nFdqwrHgp/1QR7SMQsBgC7P+NRilHUO5uzmI1askHjAjQLKJX25UXp4xr1Tk/7NQar
IBvHSDnYJO1m9T8ZQIc/nNuaaQ1Y2urXpR8kUlL/w62uSpwqmwOZWz6ZaJI2g7/CNnbF4KAxNjGD
8EQaNZzVt/5gTvQFHnYJEUiH6a0HRTEXjS+1U8iC+s/UkrzyY0OOf69RSnfTd2+WTq0Hrqc5PzB/
u/+Y0raPlRB8TTQ2nRtbNnX7V6nRWZyexZMLv9O/x+AzqH02oIPe8GD3T1xCuOLl1nEl0x+hJ7Yv
ROZWkynmWXrdj5aJYwqN9FxvrEET7fKYuL/4Gz2CVxipBiwUVgTTGPXRxVoOBNtHnYUZQfWgjDK8
J+M4itUTg6MpEEwz59608OJmC2B1dHT5DyhhsxPRL+HM4EyrtS25XsBOudNxYtoFlxfL+CE4cjym
3TVmV0BzeuLgOV/R7lwCrDhMr7Weoe6Oyer/QEJpXAK6r68e8bk31zLhqchxygfDaB9H9o+unEwo
IuTwpLPmdgrAXgSjfipjjP7S1OLqVRQ8yJGIEioxNediLPvzvjBt1Lg9yfyvRJUKnqBvb+nL+49c
MzTzzXs1OPrgo8SIAlArFQrgTHb/KXaqZvBfTYwnbo7hI2Ng7zjRWYZDXEZtiUZwH2cbLj5tM5V+
WYEMOOjvzdjvo5O2SlB5veOXO9AopgxPJxgmLylvtioMW6Gw85aCIbDeiH1B7Crm1zHRwqQS7SvR
C1NYAICWZz5CdFaZyCOxs0pfZMvN+elz0U8V6XWBAdzKI7g/nfdTs4l/zkA7Ddf24JOhnTMzHveA
0T5NoZaUViCfw5mMQFGhnrOQ2vislAdfgTEo4XFkwKOlsisqrWiZpRA6uK4DRSwBI5t4JwC4AG9m
+gA4LLYQn7dnzuBgPeoh6ix/DhevCrwg1yA5FrbT6t5F+RRZz19TUqH+fcHXaYDbREHqGEsa5InM
eOwHtJOxzSsojGsipDDQNpUnvq/wcBTCmlJgxH30dU0Q1Rno5q0p5ABo5JzF/AiXI4AkWjJe/2su
i5V6WT3KK+AoWj5sTvoVgXR5OjetaBSM67p4Tygmbv7bYff4QaoeoqvXOgFBEMbjZ1vXzqu5br12
jprbPYsYYtXKx82WnOe0TCP/y/jl7J/83sUv44uKezwJE4g/1neX+E5IrnuLEaWQg5XwCW08i4HX
/kGYIXUA82ZCxwRrCLzYxy2P3LDJRKl8YproGXrnNeEcIxDPEIdpIlcSCnXoQ0Uh9HLbKbEDw0ED
nLZ9yeUtPr1PEmfe5zJeNVUD8tNxF44+cOd8Vb8anJ4aFd1In/xxlv6ECZ3ME3THT6pbqFLaes+9
KJC/XXH8QfqvWjauDv3bfWGJAT4XTFophAvQT9fTnejQLp9XmpFL/r4G3BDOik+HfkXe9+/pX/q5
nCx6eM0owWk0/ovA/CMs6EcV7Q0oAPKBvgpiajkspBI/V/3PdSid38nHSJ1AeIHRyUKYhoWVHFXP
zOG1qrx/qsvstS3L1YeyQn2vaaa3RdY/64ShOvhurba933QOgV5X/FoAX5WxvNTUQ0sI8gGQf70P
NyrEwrJNGO2uRdYjemTs20WeezXOm2eusGpSRHiVrfkxEYYXLYWKta0dyLXs099A3oslvVqBfrT/
7zTQFt6ED7WdGERYMkWPnoLJlBVKJhbMwhfc7rA5N96WsosBmbNKMA1x0Wgm5JJ0RjHqx3MTvzdR
DzTzg0sfwNOZ7CPSV1chV9LI4xqt8NjlKfW00uw08e3cRaGdwB6qyekxPKMZNkZgSamXbUX42gu4
uC6VIHbWJvAaG6go8p4SFlVgseyOR2KolIoDjdO9an3854G+h88/IHCkj45jRzs7V7RashBUloz1
sMgT7PENF+XTymxIR5EGM0oAR4huByZYKzCdWDjzIyF3R3LrIDm/mXnTjOo7iPozezkZRANPvJAs
qTKNM6BulFClFGoWIQGBUBvVFk6oIgyTTEvO34M97qymzCTjDMrJcwG70jC/4mUgO7etWd42CBt3
yz2S55ytXvzj1pwZ4eWJm5TEyjz7JPCucVYtMRhUFtRidXgiWnvMYo9oRbmtDTdX8sON2Zr0vVT5
iAefIHABihyUdNTdQTnF36UE26I1W41usH2FwkpNVGVz9Q1hyeAygmylh0JPI9pol6bdbK/18V/Q
YIyElk8M27H2VKzAWDQyJ4c4iP66eNUme23CjxDDlkGKBnl7/3LVf1Qksg0OPHx2bpML6Me/2JZZ
/4Eupy1Qih2HUW0dIYracyt4QbQ/XDsDchxID/OuyDL/PzAeizal2K9t/6+WiEFRRw5Tq1g1WZpK
TZdHauaM8s9ClwKdVakd6TtJ8MtA7oLoUFmuPvIxi71IPYhWUV9pBiL73htUK0FSdWY5rEqxD5Q1
PR/SDL5ctMnZ9XhpGcykDlT3uLpm4lMlSbuKji6j7+BkpRPrva/YiZebqOgaVyhF1Uui8LsbUo9I
RifqVqq9Z+qMH4tf2i43BWXxZ+7gBZOM4NH9+eR2Y02WHDg0oXpQPR5HR/Md6U7S8E2Ii4fn4pdb
UlkHC5pz/g8Chc/Zju7Ox5tzNpREo+ELOZrMs9uMSMhvnPvcSKtkfvOufKTQ+o04MsCmZngxu7lY
+OeqCewDQKja47uB64ssBrGpVHxoc7XaIJN3m5W7Kc7B+GUqCNRkSX1z6parb8oLagD1DpfE6xlT
JQjDYvceveW/caFH8B0hSeR+Dptx5bQ71We31TReqhmmpIIMH0V27PMTfpQh8PxmO6KqpNh9TZs4
0qlVFxxRrILrY8NHz1qPE+a6w39X4jSLY+zM2i7Ee/JYclRtZIcIOxgc7YR2nq0lowiAPjfSRiuW
ygUDb6zkE6LQVt2YN+Ngo+IxvYIS2iv2I9lSGhSZGzvhQeO7c48TtZr4ZEzJzG8YKOHXu/Riy+GA
Kp9+aotnFFwEiKVUEpNXvjv5HSXMI7xuSONLVIU3zi+sw6YhgxmgC7Fn5WWa4pvD81JmSwjm5ZbL
rwTbRW2h3XO1Vk3KeTHSXXltR/imdXBTDWfoA+d7/gabfQoag7Z6jct2zYvtr0YxOf6C9ymVVTw8
uvnXNRvLeM1hujXKsUiB7esOM8m1aOOeTCl+Sq3CodE0yyaM581Il0Hokda8GT2teGSj92ae3Z9d
EsT2Y/mFo8ZOjZO9O3lnsYF2Py6jlyPrNQ3Fds0m9V5bN8iq78mRqZ66uqMyYlNcaXhvF2H2DeUC
hiNtl7ADzL0wDGxbHh5bOj6OzyfaRZ+BTJkoWSxEoI1OO35rymBzljbk/dhs6xjE6YO0KSy381o3
kcskgwNz36GG4B2kBoeU+i0r59YL05ibpTXyHCFUFMih7gVHSQjgO3aDJmCGzIiVpZ+KpLyexKLQ
2AizZnizT0FzAmb3TVS3Ms4HpssI5v3Iy57mQCbsN6KnBJooZF0WXsHI2LAWpo9Ja6B+bEpV1fkv
br6s23m/O8LRzHOPfravCL/axMM2sno9Sr06QKo6TfL9MXStMo24CnbinyZUGZUwBrvlcuERnH1P
TxbUNXiHi5yxp9YCh8EipvFQFv3qx9wtKLoD4gFOxnlxNAyde71mU4Bgd21LupMakiFepuNyF8nO
FD/dRUOGnrnaIHT0bwROM6TApfq0mbXJzkeQaS2F45wCM10WrAojZTwsXWs+3eciZL3eKTLTtBbd
ThqR3tFKelTVhsmb/LzEnBvGVhFafE/x3wOjASKj8Xv94RpLioKVcQbB9cZjtRLLr2PuFcbfojUO
yexHoZu5T3Bp76k/GC2v+eMycrfTfoGnZIOZ8ovNzV6jQlLrlstLUvav6yVjC2NAY8ti+RHT6A9O
B8tPcOBvGPbMtWvy3COG4rVjPgiuCKf4cqMMMxzDMIpIaRHZ/jzUJH0RxPUZjfteVKhOcx4D9psM
lMFRu2ZyN8OfBgFEaiZc4IhLFpxhYIL2L/uYwJYAtiwI2zbOz8gQZCnDMu5R3WBhaRqZq+EU4LbK
g3a0gOZPqi17Yzw9IA6SDW8QBK6PdeeyocQwfpgpmwMZ9I7Qu2F/ipgEfQV+m417pgEhagdVZQ07
XkQlECh+XQ3Vo/VR8fiIDyhzClPlgzPJyVLgDJxvL0lcXLt9cH33cvzgPxpDikf6i5VZoxj9+78E
O360G3/DEJ7q7mTZzoaoai3AOanoekKK7/ObGH0mzItX+tFH2bpfwmDL6GkA53GZ5EA1uK0cWy4V
a9nnhc7dGqSdXZUDbtbDXmARvPfEStA5WLbKdZyz1N9PQ64SOyG6QxrDYwZfwpeOGrfHVNG8vnhl
6UwLNFzqGevAMIvTZYq/CEi+EVHPH2Shcuebr4lgmpl4tD4BSnMpfgtUcklKTHMgKFkUjtI5hQ9/
SNVaCF7X5vg1l7Dmy5Mtzu+bbVos7dNefh6n4FiCU5BqoHNr7U/DmgJVQsW0UEm7ruS5gkw3Azik
vMI0QUj0qGmztFgjUr4RGwC+fo05U+ZNwhHy12lXCoMKkgcglxfLhUAGUlwdwMRoTZVJsdNVKaIR
8s01Bcvz6/XK5/+92IMOl+ZcJjcEvrnL28xhuIqr/1EfaSUvW1uu0KjH3eM7fCkSprlCMhUfpVwG
Ptyb4xSu/S/BG0luGCKPcAyiKQarFHVsXiRmIJymhcCP51bdX8g+C+S/nlxko/CWJmY1AoAoNRr7
d4HHXlEk14/TPvu0fadL8zK2bsARH5QsTe+MwMZKMKC8fG+MLWzURnZ4KUKzqz+gyrETlWgUJqcN
RBFOHHzxZ3uivVsyDT1Hr+9B10FspzzEQmPg5sKdOhn5TvnL8o/s2dhGCZPqK/NZUZ4Ms9ZXMg8/
CKFFkvCeKWrwWfgf5+onoy7fIGBzTP+pIJBbeo1WVOb/8ZsveQC09uDBK2bxPsQkmp/4QhTSKl0V
AK8CCb8LZuC4Xh529Rix3rUbQO39FeB9gih9ABPCacZF1evKf7N+e/7FkvKH1UlfV2GT1c2xs3ds
9XQq0k2yu/L31BUwqTDm9TASxi2cRID3ZrB2tL271tqbAjS4TblwmGKr1cFG4QGB/WVtq95FhdBo
vtKEiHwSpxsJuf7kU5a92mqxQNyF4FoTAaG5rqUhxxf5JdfjH1Z8IV8+tQlW6L1c+i5U0dyDLkdG
jPVnU1JTDDN27/qcGxAdryHlOBQoVGCMkQroj6TYhrq6zJJ1ydhAnj3Zd+LnPSKTIk/xk3FfBxaI
R6S9YoiEU5alBMMAlna8amloUzgymixqUT+KIafc/jI04ksDRgQLwLyI41Gb298elFqA4r9EWEpr
8Z4939U0XA/rhkQh8zXmulnHAEotCkEQY/AqMnLs3vFIQI6K8D8fw+n8wBrf4HWTuOQMT5Ysbtn+
KFimS8m/VnStTquCDI4P4ifn4tPlc44LHsAFc6l/p2eEbmNxnxsMMdPlo3qXXqQ5uTLwllqBV1jw
17ov/DkRenFd3B8Avq34zGHcOzYReaJZU11e2ZcrY1E4d3BkouHjor30d2/mPkRW1BlzI3s4In8E
bHUq6eb51p6weHCkBvKISJPPZW8EIokPIYWAuxIOrtpJkWy0ZaXxmN6mvHVvbasmBW8k7BalYvuw
2vQmY80wgTDBDhVACz7rOchywmG82ZRsQKMRJPgzgmEfd1pAfWgESTcTpKzAKzrapqhtBrPljENR
RNwKilCKj+VShobtcLpGpMBibWCsiUBJ7ZwXhJlAYIVqmXG9PDaalFA6DjDu2W7b5vIXfRa8m80U
2SDgfVIeRCOd41JEh6hVacP2wfgR3IehCMty8R94EmgocevrKShB00Jf37bC0cgtSk/rVbw716lO
ZGB+/HzLlJtDZben4z+o8qXPClhHhBanhnTu5giz46tMxT6Qen0qpRY89TJ0a5Z491miaAHMV7TA
t7kdZtKnCYMtLP3ceIEaaEwcGCqWch3jYbMO75/Dx5uJJ1NmKhHdqMnkjfR0A3t6SzHe7BJbeFy0
UpApS+3bKGcgY4q/MKJfsXi8RidpR10wB3qxUbsGYgvbtvki7aRvmnX+7KY6f4D725DsYLduoeO0
uQKc0mQFmj3B9uOJhWqZuTeY7JTrOlzrlUnPGBrPVqLbitOh/te5UYFDrrKfkLvli9Bzo5eCpX4k
MXqSIN8q4IBOiBG0dPrpqkQl77sEY9JDr83KMTcIpQJi4BmHm1KVO+CiObyooo9wFmt+XvmD1cE8
k4QeZ7N3fQRbEvTZ5lVJPpW24gWn5HggNv2IvomVe6kkugj7FToZPjIp48u0D+jFoWUsA9f3ZTvr
PFjox4h6+hxFL90K+PPP3Iu2ETx4RfhT2mIGg8msYOtx3yQpA5V0qSbmqcT6fko9NNK1ch8+nG59
sy0y6avWXK90aeDjAOFHApIzloWjmi+pkIv1/1pSbuIEFqQONeS/Jikq9S47Ubk+dDk7p/gkUXRm
uBWvJPUQyxIiU+sxWH4GpAy2TgExcgrpwibiv4DcPntPRCoRDlVwTDnLWiaQLzPKNVyqxopv/QiB
vQorumXo5QnD8TZ6UXXSyl6v1u8ZA/5f8LKyiR9UcSfwqvEkYHT41/sGSursTDye62BXXaiYpPCm
E36pr0wasRTTnfcyJZMhdEakV988F6kVYy8ywhjGquwjN9kefjFtizz5zMBW9I4/8tEl4R5qIsTK
x2d+PIiAqXw++ZLlc96pVyZyEIW277y5LYRse2jYbK7K0+47wlOkfgE5MH35xtTcHRLbLE+t4jCG
iUBxbEkwhJYuOyIB0Hfb30MdE0zyJwr1aolz5Upva3rhftajzwh5K7Q/H8cnNmvcegsFPxxwZ7QZ
0/mmA3NtU2uYldK1Yt5oW70GI5Ms4mLBT7UGsPDB0A2LtP1yHiWkjja8HWUWtJAfaJP9fFC/jhX1
4p7fJUUN1QFLA9k4aYSNmi4ZclRrmIYsDx/WCXNPe7EhVE9Z4ZaMzZqt1R12tvbZigdkTwXRX7MZ
ZcCinTmsU0xwjGp9oMi1fnqoXGCSaMDVUDlosD+36y1mThX07Wp6qkrm8scO0cGgDnMVPk3lZn1Z
dhFlOjjHyUje6rMmhnWCXf1pRbZkvdyobgSD6ek9aklgA3G0mG89iHGt96AH5Hi0n4ZlPXSDn3kk
uXEPULLzLS1cSErfjk/pqXCzeAeYzvFrhPqhtKq3pLBNjlYpnseGpUMrNtAf5VaghPBapI5fFXtk
3dMmnEKgiC3zpXVP4mkEuMfmhZjMVaBsS1poUg0s3qCkuIsTibtQTFkI6NlaJr80+gvY4NbrxnDd
xMZbNVd7eOL5i9/VvSkMnoHK8SH37+aKuBTj9GVkH03IwzJPz0s7i9L3USJTnm8yhCuiDAFEqRSK
JIOPY1p8QoZ65uealVUyRDWPJ0nosExxUX8ut/kmNvQQImVTg+pS0sZPTCQWfOOZ+gd9Hi9Ulj0F
FPY0g+fZLIzeLmw76ANC7fWpeIqGMEZcTZCEZvhIh1uoUXoRPOCJHDyqZtmGHFj9lpr7UmSwIkdA
6AXaZdLq4bCWvvqBAZqSLZ9vaBvnZsB8hf/TXaJB7ZC+sXGZpBgzbMCFUWy5fcniIyyGnhpqdtU8
uuKWVWAtldwhfNHkwWeMF5ceELz8ZplcsOuK1lxfTklGFnjp0KmUdPq8NVmK+OjMtTGM57J0IFc6
eXwEmguk/qUJHtLzrjaiU+UbHp3OztM7th/Zb1BY/NBamcJyn/7eiap/w/6mtJDkeWlet04M7y6o
AvXaisChrUb8CZ1xn+EGA2pgGAxkwdHnFz/1HiAvnijVigJVY26XWZyhfbeZMuhp424G+pNbRYz/
RQZKMPnftjl4hXtutTYBG34nWvmtnFCBemkeQR87GL6SufRKl5S41xTTFZhOa0C2yfcF1WjQ3H2u
JVsTf92gNXHF+1g1YF1+1t7PFdNmj3nMvN9eOt76WDzjYcTAm0LsDG//GXukBpol7YDcISr1pzS9
ytoPWtIuOZZl9yqPO0KP7R/spfNCcCDL4HFiFEfOad+ZsOcvahg96QOCArK4PvZfiQzVfE5R/Mu7
KKbw6Jai8mA9FFTkUI+FsYaHJyrL0ZJMJYCvHbehxK0gV2pWxeHIfldB4TQZN+xdwYllnt7dRveQ
vMhsZpczQDkAfi6iSviwewy39Ubf5wRLMJAPkpeZWHbqpuDQMi5eaip1bRAqaNKDsDZDtBSzwlUs
dHZll6XC6Y6UX/1zSCbqF2q/HmJhLBqjGJ0dmitaxbjMcaOeaL4Mq/UFy3s89a2EczXEVzwUaDXu
nrhjtBl366KIsCod2PChdoZkoutXijIGXNIu5bAFATugh3xfFM6sThnzAchO3kWu4HEtTfxHSVe5
zmgLI3KE/M6jkfH38sU/Eoww684Bt1QuLAFP5NB7l9R2xJwqgzjRhBH0udd6NgGn+2sAWZTV5l7a
nOiBTayyythNHIQ41/rigA9GlomugVa21lo2CmRIMePm7FqAuDi8OrsDaJBYhw4pJFJJn5mGSs8v
osshVHjGyWuPkbl+jNcOPa/Z5ZhfgOrgZNWV6A8I0v6TZX18vbqsA9rbA+0XXZaDIewG6EIIg+mP
MUQT2ac2i8KjvQr+VEuNoa7wXHRzrRUCGDD4J2hnkwGbBRftoAKj4G8fh80NswYD/6qlZ9+FWrtq
1/P/eUpeuzAm+jj9F27gZwuYBDn0qI4DyKxtXUgR6RUid+gRlzCf86refksxtVyFn+j8/FiZC7ma
/v3v4mzRzo/qeDM+2r+UpMFXKHJNWK+DEFmw6KslEBfeZPtECeMdTEry1YXf2lPfqPZwv3jSAwfs
gD7dpLKw79hZ6pgK98VCuf9opJxjMY2joPXs2YwiKdDauQT34ZZXKpG9LyHxqQlEH9WBtSDmGpcw
uvkwZlqSw400INjkWxFJfCG0oiAEqeF4iDsINuajmRydORn7Lg3CbOrbqQsSZM5ZCrTOwCR0dtGX
yca6zisJOBKuwD4nzliBNkGK/tF33hDHsoCzTvflrRHBufybEqCWxNQBkt4wn3wgjs1DvO1irHq5
/ZeInSQm6lB/QTm2QXsE/sOXbSwlgTsfEpPR8n86kR5RAisNnnBT9TIG1IEZgOlakzX4xnD1jjh8
GjWcRm7RSVyrYc/je84bnm48WFp4cozaeaFmFBd4Q7z634cAAzbL4DSutsaJjpt2Bg6iIh9U6jLe
IUel7dgDjjIXXjKODJLsut6ueGA/ZyqfOo3WzgEaekeDLTBcJKXiKrvyBoGrhPZNWmbJhpn6hU4X
zrfSA11PefS/Xfm0Tt5Vt07E/l2dNDb6wPrix+1sOuUkLXnougQxNPdrbZio62X1nXGNKsd1pkuG
L0b+uKtLuI48J1Gg9t1VFN73+4Ov2z2utZVtttJToLs1r6RVztC2kB9k5ziUWm2Q5CPmejPFJ8wd
y3iZnZpZHqkUw9g9QIuFL3ZcNHjeN10U92/AeVKi1NJ+1DqJwSm29DyeFy26RZhScGGX3gyulG+q
qyRYOEvLBMIPOuxj/VexZJczjRAG46OD9X5mzF/fGg6yh9N6Z50Gfc64XS3U5AF5Ft24nuoDZeap
G7vxmqOi3gOa513UEV6/iLG8yPF/+h9LKm+JrDLIJTFysnW36Jn7bMxfLH5S6rP4BLeGxxD49P+E
jKsgMtkIj5iwMxCSr52/t8xOjUF9+9l/o1gTu9z3f9J4uX2vnMlBfh6GpgzU6MCxArExXraWihmg
uGdXq0rxSgx+aVD2YQ4Vm28pj7CP+IIdnwPeEFlX811zXgrJ+fNqzIoAAeYG4NPWF8iDX+8o6oUS
y2N4GYnah4mrquNwiVcB5wPS2TlZIhCInw2+rwYlhPna44DqfwBLPHH5UpcAHe0M7g2j1r9Fntg3
Z5IR+pGbP30uhm4I1QamhsHa2iwXKPk9IPez9bDfbVm+9DpPUEqko2bm7nGwdiu7jCwjUi3pQB5s
0c5cWWkzJ5gFWc2gU/gFOWMzVrqNS1KoSTgdoaxDFljYnd91j8nXmBHyMzG6687Mpat+nZyO7yAu
3+8SgDRu6JbtbdVRkRV9QysgV/0SnWX3nO16AQCF+V0n5K4VT3Nd3Vhby1Onv2ubTnvtBNwl61mY
4XCgDT/XyO/EMbM5xoBE15fdYRFrFka9BMKoZIrWl30YW27BTp2HgD7I6Soo3WK29mBN2X9nQDrT
7PdrqIe7/FnaXgxvX2j+r88rH8zIadQME4rNejByM6WlUsRT4mclIGeBqXFF4MLE9W6hXiYu/Mzn
u4G1ETCCEsZ5NwDbthlHRioBmBEVj4jP+gXg0NVpSZKLM1yrwYaVC+L3cUveJOlwfX85xcNBmSgX
TWX8d8Lmf3vW9XN08eO4LaogbehoByJ/UHkP4AJqxlzPBHvxK3n5DTSgptrJ/koQOwNjEegw4tRT
v7FuDBLT+kiQhymy7O8YK0jqlKAW3f1/5HZDDmxf/P0Ac3XefsV0RfTqa8BwIzpc990LDlBppQHy
NqYKEo30N6ZQxGRWtvl9eWtTXGs0PhxnzoeNMPyhuyEPba678dkzvlcI9Mgmc2gmk5uBWwyowNsy
FD0VhXoMlcD2nkAUnCcGLMHuFrRbyf7M6Gd6zrUQfmW6S1CapwJfjKHFNxDPSj9A32sgVyoX++K6
B2/gUYRqdCEoT2kEdq4wBINcYPokxdOF0dIv6YMTLP8hA+Z824LAsZYXhlC72M69WIKfRNi9ZG7W
gTnw01RymLdXeosrUrM8JbPLg72C/VhdB/itXemx82FCofQByWBq20b4suS0peEBCe6E3mlOPmYf
/JGMH2cNmULEtNEHzOqXrHVPzqif2TJchgz3JknIRr09VO1qwKw/4dAFviAqsdXb6ZnEFGMRzKSP
B8egQ0f6xJb7PHXVYpiCZQD2KEv8Zl/5OE/XzPaOPGlRrLbuoJ8FvjeewMJpLdDe5OgYfxMKwYYK
FNsAsjdN7BsZqOqwwDQZ/XDg71+7/p2D8mGwVIhVY945NWok/5GESuqF7TF9R3RmFS6j4KlEgq4y
Jb56FOq1qB/vXlmqrDX889zsOEEGea3jJ4zVOYZXu8b1FAHg7ker8V32W7s7+nz1PWklXYfB85P4
tlTFV5FcW9WnaYEcTB/V6Xdd2d/lN/WU/moRBIyA6rGLHOuhZ/UBu9pqKJUizaG194PJk5Wp6PWT
3Gi7ZVmPHDSxiHWTv1bdunw/wxgc615bQO0P8n1IOfPhykOUdHha5DyyV+BqEhP8JUeDP1clTSxw
2mKJkgPWIfcmMsR4wDQ/5tKyrsFCvmbzYxi+NI5OF+9YUbTVVYCI4kZOh8STAIBGnn3aWyI9kPsr
vNccGl3iPwr4StBJ/9oZPh7fjRyFRvRNM3BzJY30XyMP0CAvSheYHwkF8aNQQrYvL5DeOgK5DQjR
4zWf21yqIJE0Fn89xYACVBq7zicnSmB6la4VKgN1dTUPRroJlFfRqY/dnmhXgRgeNemhNmW8+VWs
13YdoLDFUwI40hibEJFbUjsT4vSmNdaaWcNyBayCS0NVL2lFzwhFjdbH9RHVRaI2PlW2DqoqDBNP
u4nS0iujOip0dk60vQp6noI8mAFI/uyPT1Tr4BFcjcV1rD4hhkCHTIgOMe7xcbz2OkGlaRLo8H38
cU5FwiAKUs31HeYEsSerHKI1HTH9ZwasaWL4VlX4Jj8EWE9oAtC/fNkDnnh17AYqdwseQ+bwzZQr
8L3RggPv0g06xp6nwT7XSltd1Av1dOm6o2KCZgwtks96wINCCZDEZqmX2yJgkffVIQ2KBeeHVGJ3
Xma5iMrsJYMMrQupk8W6SPOMq29Ipn4VzMDeWrXKgJW/cyDWqtwxHQ8/R6qusZk6fh0kIBn+gy41
AO0uR17oys7Fpv0kxREP5noIVgbQAkzvMTDf4P6Y+sVl4psK2KAfCJjLYz8w/kj/kUuWRkSFFG0o
RWXtxG/CaeotK5PlqSDabh415oW0wPFc5OHHvGDE90dmWoToH6IfTvXrR4MhgqzxZtsfT0S9syDp
9i32iYv5me8ysZoEGsMMNgr9RyhWeE2kZQT4EJ6ow/vGd9ySx/wG6/5rwVc7xTuq3ogsbH+Rz+WZ
cvB6EnhuiDJHfjq64SPCxHFsR6Xm3c8NRyrlWTC06RxZdIqTVjHojbQV0ypXAWwQ6gt2Hm/JNOFq
LwliGeGdb6ESkiwdA/kyM3h49dCRusvGKwxKMYkun5T2vKcsMBvFl1eAznaEWW4d+uLR8yWAuHSN
pmJdXm361wkTyZaycZHLP86P4nUb7VM7PFCcviVgJx5hyqW6Vm6nPnRu/8/A6XIOHLIWgZCYUMC4
G6ROtlozdbNahpe4FADpuofVouwvf/tgzwDXD85F1FpmCoOTo4VS8YvwN8woGXGIMxlGcUnHgMQ0
fyBgkx27OAzCygWVojg4oyU/6hRwnG5/39wjl0GvZkwF91ThDT1nJfynLnO7FSiNhhH28RI6Ys13
+5O0ckrjFGxs1vEn3jYkc5LGiGyCg1+2VmjpyoA+qOjl9qIIQ/PpwCfnrW/7criNAXpDkzd/S5ue
OxvySJp0jj30IX3GxE7Dsh9ilh25P8zQZWH/J8MuIaQNhigxtdmPDSsUTeacX1oakMVgsrbPGuF/
3vgQELqwF0DG4tKxmjAsTsb6wilSu8Oskgt9K46/Vt7+uFVFdbfgnLdLUmDzZ4ClUE+FWi24qv40
3lz8x5Sn9eUXceP2i7gKjXPLaZmfM3HjBVLrs+OMyVMFkWnjUuRbfFuYtvWpHGNsQ5ZZ7ERZaNM3
cEhzuUZ6OwmsIe7YygwbEKzJrE+PnGpsBrwsWrYay2mVPItiWJWczucCFlpHync/aMtKOQjreBcD
UJu5EJZh0NHU5OmRy7MojfFbEDrE2CxVGkrronQglt+YiMLCcpe4Ohqxha6DpbjapNtswroagcwi
c8HVaJuITlBvo009LH1TYnZupp13XvtHqMjWH+m+YxFieQkB8hJKD+oal1glH6ipPp8TPGLIEaOz
uc+5GXcN1lrDT5+WO58EimVqtllsAw0kjqZBb2PQOXclUGwD6FUjkSB1Kkfouc2nEAJ/z+vtWvSt
CifsBy9DAPGfqwgnWtlk3CSHQ7wQTNXZ88zNoeOpG1qmChRfhLu9JRCuFpLUauvGklSPml5CBOcT
aYd2WLep0/BrsSOLQetXKZmEz4qs0oy5unN7zqj309QcA0JC4yOsMdOa4xJAqCZrlrOiciGvqiEY
LFoQd7AYxk1eR4ccqawx36xWP8fR8pIds/TQgdcjYMcGP4Z40PcTaGcGRH0kpEOg7SIQEe1s0ka2
DMbzMgDqWRdkBgGgo4kf7DiHqAUwwDQ94lInMPiKkcsK2oxO2LA/RDu47zWSSV+4fQPVLYTYFu7k
TLfb/TQfrX0BvZPgvXv3fbKT2iJtXxNjF04Xwnev02ovef4xApjL4PrMCRaWmE1knjM/srGWU3gg
egdgyGVN8JY527KIeDkViOKqfYEL/ly3dxkzgl/B+UGTwaU8vNCzroEP1uds6za/JSp3Dw7TDDfN
K5tWkFcUroaCSqWO2NF5Aj8lZ6iYOV00LbfPh1EEEf+/RxcZHGXPCh+u/PVFQWt4om46jvh3LgmP
rbIUecOnp7tPo+bKGWV54ivH3Q8G6LXQ8h0k8MVGQI/avSErv3n4Pp0RmqDc3ffy1A69a8w4B3Ti
UW7/CGk6juLm1HPxkT5noLyPZ0G4FbplU6RoU6F7b4KL+boYUY+Obn69ANFFDLhlqyY2r96X2X36
V5juLb5aywwcPivAsZ11QOnl+DBC7vhCeg+W+zDivnNUaJIhoxTzt+ViFd7eayXB4ekkCQT9c6Qv
0R6d1VlbdXyg1GzSBDp26tUB1aRnEFDmQhaVzARsbYyQq+Jf5W6b9QMSx9aQyRGKmdBuIfjwaqwn
Hg14o1ObP/mvdgfQibTWHCedQAL50Um/WhLR+Jz6YEBDlszEgXGIaTXAsTEVdPqDcHLYdlKkuosT
wuXBbeP6zCcGSLUlmNguczVgjeV3MXoXiJhzWiPKBiLtaxYtwKB29FXyjVe9jj+Ur5dx1R0B4MY5
K4eieDMkyPLO+IUkVCnGvnQQxovq7hXGCGoWAQoFC32mwM8F7cXXgsDxLSta+Bc3mHDf2DENR5uQ
JBxfqm27/Dj4W1CRimmqcj86iJ5dskyIQSvxlzHyn2FNLN6VIqvoGhHokgneDylZ+HaI8C46wBX+
51MdOl1InG7M1qQAI3J92Zw6ThoP7u7F07BVvvD30FLWF/UrxlK+RxNl9Dx8gIqxfG4ATzJsF0Xj
Cw/qmGCpazu1Ue0454VW2SD/Fo7r0dIHJbMCm9ay6hMyECZ8aiD8xffSgWJCSDlEshOU9CEUH4/g
0Uh+YCBvIUb0y0ErGD7tdf03PsQBWFL52UpB2m0tdFu9h+daAcg1CF4dX2nUqYSCXLwmxhsewJPr
OBW3EMNAD8oHI4UUdxTVrjjecbtrxJgu0e+AwiZUISg4/S22MgxulExX+A/XAlpkgSF4OBHPZ5Gl
JV2vJeg0OaPfMQ8sNV/uLKBeufDoH7PsuNuPEj1T1DLASw8OkhQKs6rNOFdcqhbRidrdK7XQ5kbf
Vc7OLASkjH+duQrB66eiQ/D7bqoYIu4rLXVaD1KpKDRbiN2SpYOnlfnDu3ua1rkV2cCI9JpTT+o/
1WYZvQQBPgOUk/wD6sQrGt4CKerhV9s52gWKxSGJhyXN842GjtdsoeRU7PKJEYfTIaTZuQz2XuTh
nWPQjyE8pkddIJzwOTf/otRHwjhBVZ0gX0mB8dHsReVkWWDv1yzUQRuaaPSPWyU8wgXAqFC+w0yt
+a6PdBYSb4I2g6wlPApfBqGPPJFH4qxwwbteik5GZGfFtn44DmpY6aZAOxCXRy2a62algISPDnSK
bqeVzZ2s1Oa1nuOgXggvnN8FnLb/OIz2pZhUw3DeAHq7i/mZhSE7PWec2wwnPXLdjW7jorMIdpL6
V/Hhms7bvczZLM9AlotvgcnK4h+Ag+2/d2OKZVVhpopAo2o5xMWi2MOgsn/Kogxyzlu+6C/+8z36
wnUggOmHARxodcehF/nmMIM0Cr8XVnfI9Ug+thnSBX361Iap2BH3PAhDck3bmTOCHPgh4NpDcnZx
x8hpa/XK82cMCoUCbju0pkQw7d+1u2cAFkQzfxaC9QlgIStcRYRO3oU1ArWJb24JtmoOHVEBcyXe
LEo6wB8eEsLAg/adFqoyHkgAcV5i57UsVrvBk+f+rikDj3jEtIL+9dtZEvSQ/h7kKRfqUCTw7VZz
4yHfRvQKklnUuBQeyT2Kc4qNEEZnOB2hhArUblPMovtSXuX8vB+dEFB9wdROXAB8vPM42fzltuRg
Q3DlAEXKfaa4zJ7/632DaCQVSw6KJoDa1eHi9x3MY026Dpy4nLFldFaM/ECuMX9o93Eyl1AbUlf7
T8OoU4g676EcQPDRj919xaKWALf3RogD1fcKucWG6ywHIpPb910Xok6brphxs0NluCs2lTKoMOWC
OxEHzUErXJLoTudzWqXS9+FVZa32RVM1DkXE5jbXzaVbzD4aUIAL0ngCL4iYpGj/AFcJ7/5+bbzu
kP+FAFuke9fwhpcRqU6hFnzIHpYs6fwQG2OY6DcR1Oyob9HYpuontpt5v4ns4NhZ4Yg1y53V/OOQ
YFfNvSz6O+niZ6PIbUGDm3BrIjcBsBIWvyPU/ZZrK7+5v5cXwagsOL6BusIB92ZeH+nOXu0faLKK
Lbg0p+ewyIFNdmeNOE9vFFUA4o0FP4h9gL8+BivkM4X2cLkl3YNDj/4MjcMcF62dVrEMPCh7mJBk
w7pxthQyKUEfHqciO2ScwvDvNLpBftjGa4ekPtcTTxAxrkOdy/GHjOr3/qJkMfuT6M1yVi3nvrqo
AvQ1xzlVTW6YdIznpQ0J9X0JAFvVHOKtSMTF7GXCKqzYwjdg2Ki2549+l8lkvwoVDMMTwzxXhVOd
sBEzCgHcbx8HPLQmQ9U5av0eNZwnA83VuTif3VIsjzbhWSZS2LkEcZqL6bi9kuwbBsxnhM4sa9mb
YYv+3rs8joC3HzhAO+ojjETHyUQmSZtMFCsyiNudbPTzY5KZTwSnv4zSwBSTL9p6q8n6qq0UH4sw
+ykCoLV8nKeUerMCZecHTMTFSgWFNTYZACEkoLOESpzWAt9na+sxRraYgB2K2VX0ag7lxPXcFiXy
rvyxHACrnmbkNzig+QmsxLSqJezl3YXtzLb7FpxAoWhXvvn57/SftbnBZiuYvfI+uOidC0dxQTMc
mvzt2Y9MxP9SdY/Uuth9rrqCZdvRd56XeduTAMSBlOHcFGw9XZaU3Twp0De7Oo+bMKcvEslDdecQ
BFbX9PO6Ir1RH+P7Z2buraHnF3Aw/GNixUBw6qtFDbz7hDJ8Kwy2b6v+ox7ydT5AXIxmBBaSE0Ub
9rzYdp8YXDqKIRc/1EG7US+5T3G3NkEWryliRrEHYtZymTW9oI4LVu9x0LFMvFMQtJnJD7XgIHYs
zrRnfzPFK9pbg6M/2EfC/O85urZxLQAxecek4ogWFtoBzzG5azLOiufzBLHZSSS5KMqAQOpj4xir
s/qYOlrHgsAoa7GykNeB7FkRHA7F2m8Zh8po7kKYpHecZXpN683R6gGP6FMTPbFjs+3UQBTdYQFr
TBlB+vg9sGCJ4V8Y9//M5cxxoEPd6khddR4Z8mldHljf+Op3J5IyZT1FjnvEE8s9GuOvos4TfTmM
XANhCUNAdT/UIy7R2wIvNoG5cRp7ti+DzLJEV+yqzxMxsWneHUS7Awpp6jXvTjqIcyJXRQonAAe2
pLkNIV/DIAZ3VQEk8gAwOJgppBYlrcFYLePkEMG59XfB5LuNYd8IEnfdaSbjiqMfv327Mg4Ehwy3
C/OV6mC87LEljH2+K4rh8Iqfi/95F6JtkkbPyB5QE4zE2wBkaExYzuwm7ite13i/M8ou8t/aoIPh
NKPzSY+i2+/2Dm56BYwqLuyVgkZQohDZfoy3QrRxCxqQgHwk+0Q1BdfuI2KkyAOBKLbWGCflukO4
lANJnR+3lcKolV4ChB23m9dR2FgVF1FUne7F/bZHR4EkO5Q4q4BCmZUeNU9JUDkz82O79AxPd30K
2jFIJ9cg/L1lGDXfBmMlzltJ3574xZYrqKCye2jLP5pk/aTGN66C+DS/m15l1mw2c7G9+AfdGFUA
HZAuMjSKmhWxhcq56un1TXOFaujnt5rG0bPQ16VNes+SmLhiko9cLhOQJTJaew9gxSYsjYx+2Klt
HQiWVod5OjCRCGcGGO7irIF6NmvxpSSxozHDRBIPT2eIHnSb3UtBShmFr8qa+TookhWfzH8SeK/n
nNRAldJ6T+tnek84wd/6izw07yG9RGCzafnMfcxFa8GhJmZPr8YiVMuP9aazTTDOZhPRpAfZhba8
Mn8zsXBgfeDWsRL9jBg3PiXLtkvgFvWgNTJkJZDsurXfRyIWcL2qPDNdGhWDA/MAaLEHJ4hAflIg
26SZJMGXvr3EMuus6W9SHB5j0Do8XUTA125lrtJOah5ie7/LScHuwqoylgfPjiKOrgQd++1/chWr
sVLnZ54oQhkZXS+uzpiNa1GmmQksW7+M9PAqzm5zqm3sVN7D4ppEzZcA5DwuQfV8ul9EjOy9ivc1
hNJ4rmf5C2XL2wor7QN/44XDxwnMDbz63XhdCcBLKEfhnV/9YI2/q8IMaEHLnNmfJigFEmGroHrL
yDrR1EMHeDysI0SGS6HeH660XXeIGoaTZzu6+RsOgMA65BNvsQaFgUWRJLQMtZivSICqcZ3/RBrC
rXUH2SL7za3ympTKZfc8puC9MU3pp5F7fqWgo3hQxheLMWa66ajer+N2FwJ6qsqBAJwwYpVJi1PF
D+yfBzjG+8CoYm58tS3TBdYe3XGp8CnncXbhVtGGa3vDljnzQOxTPuSBYpD1w9GXVpTjGrzlwp4E
/9+iM740wQCfNkxPMunVtH0ZQoBQZHlEuIa9WS9h0xPPGwSvvikhaSKO5a0TzFsksxF6gSB3nnls
+cQo7gEWu1VYsreAfQh1jPQI6U460HREeN0t/B+Id+Xfp0gSrzkmwhrTMlAB+j1DfLHMO4obrJcA
FhWf80CwT2psykozWo8Cfz0SkBUUquO1x53olx2JHaosgxacqkBdjFg5FOxIilBIhDkqEcXIcvJw
Sepbo38AfddtS2kDDfWEEhgZReLbZjyXofPAbpk/RdsV0DpQ5NoNsfZrjnt+HCrqe0EKUqvgWGKo
M0DSbntmj0GAGI0JeDQIa04PzcqIhZ04KYUngR3ilgO1Rhanl5K2sLxkpEJJa+besC7M/n23HOLl
GtSkpSptAKKYjF68qu9QOOmJdatx8xmkMvtB2HyHhvmQ1brTqGNckskQAHiCibC/jbPst7IpU3HZ
tucOuevECFtFtZGWorh1i6AFXHpg0O7uT7ToeJoI1QCRGRGD+pIm2O1c2MJ62e1QiLq2c8gJ7IKZ
4EXER+VHJBzppXbXjab/RWqn/kVHwsuhBMDR+OJ8TjWxfEbYTg7lUNDVoTLW6wku/MmcubEVyCVG
NkWzNzf5RL+UmNerrKF328McUDXZgwNC8IPDuUTGXqf3plbnSCZbM20s99JcD1XA3UU4cA4+P3RV
kcwInYDKAWu4FJ0/DuFUodpAcYmYhlssGAwWbNOFNwiTm7hmTg2V9KXRCX3/fE+TObZhcsft1oqs
5hZpdMzW5t5+3vFESQMm1kHsR0j/0kSU1iRqeBcYGj9QQ4G4nDXGq5/yLKVx/SMryoHGAFjs9Tyg
JyWXBFgi5JD/UJj5vVbNyJn+hgchyqM7lG20wEN4oVqfvbdWDr5Ev2wKAernv0jN9CRUKxdNZrk9
8NNZc9RDgiazXCZD6EmgMSF/TWDCqU/EGW8HJ1xCBLkrz+90dassPlY4fp8nUsA8wEj3xEJ/l3mJ
xFK37Pk8Hl+BsCcYuO7lkDWkfwmjEu7fS3ZGpKnNCAQm2sUDjQoesntWtlGFaYDdgED9zxQ/3kyR
eRTgKoQHNL3W9tB22Tu5EaXRo8n5yvh7svSBt0iLeIqfnLWLzqSL56X/gG1K1R9oExe+nBubq1p8
MHF/tqiL68dDcCqrU8HM4Z9fAUwuGm+iGn+NfevKK56DzE55uv+c8DsyNg5j9YeQ21h5uJkylek6
MGfzzCHeaBKiM9YGT2vW0Nyb4K9rYHwoILFwTLFzT5URAdf8OuFXkksItKW0ds8nDObdDTO7K/Qm
P6qnGvUq25zabREXYxfWKqml9YYksTuzMVlNEzE+ECy4EMmDT+sF+r5XAO+WuwjlCy5bZ2oeBOGj
42OrFcUbpT93P3x+6urafTavcnMtcJ2uYWJhnHEPpu5NwlusHuRR1xhsBsK8+v1JMy3Ox1Ar2X8k
dAh5S+CevEYa4p/69fgdznD0Q5azHAtMhRGlRxWazxaT9XoMcuLsv+/t2e8e/Prp/KpALKSBTEy+
T+MHoNTIfwBvlHxUtqS1xtcd+vuPrs+O9ZQcYHq8zI2q9g17+ZLUmDLCOojBnTTw4Y4B0Q4S4oCF
XxWs4ZGopjgESNLLXeMPFx4L/ZqMOL1svgIZjtSl9VIM50HRU2lUof+nBrM2FME7y8XNisY3HUdS
2ZJattQDPQ/NdhsZyVHQAoumadWInpAR5awfH82bCDtDaa17akllXDoUE4mshLD3bbPLc3jUdT+Y
SOHf/RU5DbBwUjDEw4SboQZqj7EIpoViJgbKvFGyGLhvhkGqlpa+KiyYeoQVfM7zBE/CBJr9HdAK
pmqLnvduI1zQSyqqJXsQ9ie4jIZu1TrnoIXDL+g20YgVUQ5V1A0AeA5NmPvWjcYCAF8dRJzZEKFf
tBPPGON7Nl5EKB/jkLCp6FUmRecui9psLXshXcqdmWJdD9tUHkVdCsOdZe9swZSYiGLy9F2JbKvf
kwr+CXPatV5paVLAQZrCupOAzHDre1oUy04w+R+PUHDl/X8K21cixvNmNu3Fxu4MkrmbRI9+a8wF
oma7dGW5BQ/JDDq1eGrs92VU4y9MbnSwb5fTVYn3k4c0ziidNUXMAjeAYs+0VT/g8Da5HymgYlum
YgirpzZj5EHgqQneXLS/qyV21vDzSFnvk6RJB/BREvgGcFyG6l6bwzX5i9UAB4NDdBFvyc/5NoNJ
2nnOzgt5vo65iXB1UUE4kPLBIHvRiBqyASrcH2e5akp7kFz6Fbl/ZtNC7RazF5QaENindPFurZVN
SISVUPczDjzXSUOmJMjiMLDFMd8dDWSFuz690gG7vKxaeb5qsvlIWF2oWLE4ELyxsPHPsFKlM7Cf
bpbIlyZ5RJ9YSkC9ofLxYUyPuzf55EIonSModYnOF/cYVZnZMfm/G8CJQV79wZiDVllJE/80eMiO
CQ3lRIjHVBYEY/08uoTWO+MzwcHyzLdWrger6QKYpSL8eFF3xOU30mLRHJ1H7YEGT2ISulkNyrBN
j0eGzcqp/9u5B07qwLbZd9h5b2Ic8EY8LFgIhcaE99r854DL1/1pZq5ipXcaB34crGtWcINqHp97
jZ0jmxcLS5lNPO9dinCywAUfsb3bydhUzwjuCsPU9VEzsaPQKLE/QiJ7j+3QyMc9W9grQDGMvPDK
p361ThmswUdK2W1uoNcA9tlcjecpPl6XyyC1AwnhOPAw7PJVWQN3ml0laLHWE2GhFzkgCDIlxP6h
dwM3XIArsvzT02CoanJueUfNYwiFq7ABEjVyNndhyD8j+HWa5DlgBPfPFjByoq/2AdtZgVVa48PQ
wVaHLxvyxQ6ERgeifKOILoIRgli3/stayenCUH+pGNdadJaNTzXJFesQYk+zR/UI2HpwA7bvOUPc
T301q+oIC1WeBih2XD+/xSsHhtyYcbO2nDR4m3uDOUlt+tCkVTmRNLN7TzVhC3BbML3tL6dMywx6
+gL/Wzh/5msI2xg3aElCs/IupaLdtt0RsVrTMJ7IVF4QMZf4ZGK7PJOTft9nyyUCz7tPPLFbl1dZ
umV5twyj/488OWNJxPQovrHVGJYI2xeVwwukEG6oS+scBiPcREaQ+aCtE0HRJuXd4o5/bMcJz02T
3yqtSgH+vtjNOlv9Qoyi+yTzGgG6WJiXZ05IgqRR0z4BMq5yfACpRPnukprKcnBk/TMM6BLTlRrb
M2LK/u5cQ5uPgMn5ntdcBhX272KN04PmBbO+M4fXs8YPK+XutJTc0mxETUzxixEawx01g+abb3W5
44yU1sbgUWkQG64mRuoz4yi+9Z0W8TF2GQr1RByvojZC1E8elpYrLTcAkBEdtPgHwCM3yYg9HRpz
D3fRi40PVPUExfkN3oYJes/h8gErb+V/QLyY6jejdBu97q8vCZTe6YzD5jllxyeq2HRw2HYWPFLa
IDNNpdMI8cvb0IBHUS5yAo6LJfM2U1Z5yjogznkXTDrgkXLD8VAl6X7e0ucf6ACIue9DeqJLX3AH
kOf2iiyPxxcxq568MTyecqj2DXS7R3HPDMjjahg2wra58SFPs6GvEtNp4FfXaakUOUylPajc9NjS
OE6mG5Pe9WIukbSRItXXS0hL0Hj9C+X4XkTB45ZhdVR9DLG8IQfKoP0652CDM1zu4wkqSrjZk4TF
rbZzvZ37DKLaoH5WxAyr8e+hDJv2htzaw41ovIo93zldpo5riCok4N1JRAvvBNP36bqdYvcNUP7d
cXUT50/Jkf8/0RZ7H2/Je+5d6Ton7ma1XWeebtD/pPCHi7XGrHnMJh4bsacGFInhY+nFLGuoWd/Q
fBGLubYBuv/a98mgW7S3ydgzyuuyGTgu97TeSA3AoZ25h66og1HNi8DpAUIA1w5brkpR3JcNCi1U
JqPEFVIqOU48+y8dkpJSPZCyDJgVVD1bQaMr7GMG7TdFIgjXo3+0aa81c/GRz5PXtA9S5axFtOZf
68XGreZMFppI4PRyqwBWdM5VLaS9xCVcceOnjuLuWF+0ef2arRNM3XlcefTHB9Ict7vv07iRbp8m
GNutOL1S8B7J09l3ffoLtQBPab74mh6cggFGQachvbYHoXjyyl1h3dy8jN7s1cL44HmecHMNIeYo
NMM0Oiws7QATT02Q/1eHqz+WHHobYjM5i6S4tePYidDMwDpgGDpizU9YZcgFcX4iWsOdc/XriKel
j+RGfCkP4lt7oJj2vpeK9d0lt2RzcJKouIVubfFuRiK8W4GDl2ae4S7vKIrsgmqRGmgEC7hSrRwl
DxgjfD4+ohkQ3nbpEIxikhEYnBYs55WaoGQFixMxBDPFzeRqwq/C5W1sdwCgzsxm7CI/NX9FQBrr
3Ov5qc9V0gFe5d7kEm0iZhLlgRkH7GVUmi82BPzjf/NBMI4MVklnL1zG6q+zJinbovj3PsBdoGur
PpZ359ELT+LF6EzmatncjXpacWaUe+8iy8eM534VeIARINeLhtU17zCiLWDXqzBzIdT8fWD5YqAc
NqL4aazVJqSg6Hlfmm1yYXdk9nYGynPowvX2XzERmjcIUC/fBLBcs93WRlzM+EjBWtcij2xLjsr8
S1zt6VVXo2nsevRcGeKCeKnFCdAxlxtKShuDOZN0y64K6A4fLa51qUSEzkA/ubuj+Yzbsmss0dlk
7lYWi9pvAw/ONOtJZg70u7kKw6PLIYVcdFJ34I7WuW0GleB4HKkyIKZwbpFDQjtvk7HO+1kfoejw
O8jE0kqxBHOOwpaZ4VI5mVG00nOzfCr+NwZ8hSH+2uzlWBNsG0nAnAdrD7CvDwBJUSnTbYk/Ye69
1R8YZAgEqQ45IjJQ49VXDFXwEBspx5NZYIVi7KOmgPcZ/cVu70eH90WLUJkQsWnO9T5loKjoU7yM
B9BBQBRklzAZ35iAOE0ADpvARoH2Z/8m8v8Y0NgU7LfEDgA/NRqBm4R9EfnA4aD4Ee/7DXa71N/x
JjC9CVts7GHjsI5D+/9mRDuBojSwLj3rO5usnNSEHinVflDHwTm1fFZdbjXTYJBWNi7Cyxqeen/Q
t10z3Xb6Oezn5etfCnXoX1XEw3dPqqtwVuJU8D5mtS7A+WW3X8l1B5HH82uFaM7BDLnJQjNvKIgT
19WJZR4UmzCuuIREfBrKECQHHnB6Sn/51ISjx1JafcF/CVaeN8O87FbKHi/FH6XUoe783tLIOUzP
m1QVtXAVTm+YIH2e9ZI3LsqGLJ97+4h6FU7Wb1/yYSw2ptNCf/BF+w5Tmy7Tew==
`protect end_protected
