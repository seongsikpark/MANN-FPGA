`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
B9ZpeWvBQQjY4dr8OyQgCWD6kSA8+HY9SzJj88aCfo3JohYFlKYJblw60SIQaUnjOxXx8h6ELYIM
UjD1sVmQ8A==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
iwVbhZc2P9arGEbPkPDN2Ciczyqo1Bl+qfZPC8pPG4eteDJDMYhL4//JIPliW3+60AO7KZbyirpX
isgEMka3z8ObvLYO298sjCHDgs/FZfmZsyGmSoPOb9HHtHVciE4p3TjlqyIpvkIcyPdJ4/fD49Sc
nvJ9MvdAGyLQu3dwTZE=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
oMpLZGheLmkvkHecy891anqU/IxrSwqdYJi/BCqFCgNsgmImYYfizgd6jy5pHiJ60XGOPHkcnOTy
jxaGYxBI7Juc/kfJgViQFVV1aRuuXnLsEn9jAYeCNbXGjMOcxwPk3F6E5P+SRFJdfx0KMPcD/wM6
bmyeQUTBbAdhZX227QTipqzrOxkS0QaVhzCDUr2q4VKPQsqZcTtsxxafdT3X1+kJkg+J8PgudGXM
7bL6m5q4mAXKVyd0GJhD7Qi8vPhpRKok6azS8kpVpinGEW2jOl+g30xnHo34r1Y57zE7Hac3U3mE
kGglks8mYGbOgllRBqR8MUiayaf9z70qRFoHFA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
e+nYdllhcdKHJg0r1my/ydh7lhRKOoftD3bwWM6aLfXtcw02WfQ5kb3g9y9QOMp7sTQr6BHcJLPt
ngjNHJ9dYgrGajeUJ2ATpRvbTfhC0dOu8XDWytje16mCpWOwZ/hGr04rwbOHpcTXOPGdOE/VrnEe
X5hIFArmQ6cPSEF5nr0=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
zSjmKksidjShQsfA76nBwQ0teiFzoZZWQ+NicoSnGqsbWtnh1xC5oIQygAEkiJ7KViOh9n3kKUHn
T/7xc9+VdDMh4m77ilRe5mmwu0QDyeCK3aCjSZoU/zujjnRNCwncEiNjU+Gv2xu2Skb7GZ2pLHN/
r3bxm8sfL9KDPLKc9jA+Vo4EyJ2KkfE+MdKkuK/XVdTgh9PRlhFmAMvYUBNhWNbe+GfbAcQqFErh
Wo/ACLuJCjJUcZa4Z+vmEqQtU8uNZWUzI9IHtywU7ECvMX0j/BlC1BtXYBIYzozfRRe1iYXGiZkh
rHs7xrnQ611g57bj/SBA7p8lNIET4VbFnbxVig==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Oksyn1Lpp8o9+Nend2BRJah5VMeR8XjajkNcetZzZabaL63UOeUOV3m8kWRFtG+ALxcCfCl1m3XZ
RL/RbQaq5UobujWx5eieDvAIYrWHCxmWjy1EjcD7YuPi3VynYio+STtqql+Igru+3NjtjAZATsml
313AMJlgO8hvLTBcs3+r1Qx7i+2ulipkTg7bCX1sFywvBbYGmc+T/j6RXFVM0SaznzSl0PQYxxAz
yjjhfqBNDlAfLgRFjyyKSpGR9PWx3mC7aXsYJrTwQUQmd1jlXVRh8zCaqpZhaRQNbIlT6/ISEfAx
hJHHib4bco0Yfo3fQ+I+EtzPmOJztekW5j0x/w==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4032)
`protect data_block
ceU+yUO4VzpxiJsMsHIFnfWhnNW3rWYyYkn5K/eh4W27F7lbF1JTv9S6E0lw4LVSZIy0DuqusEN1
dXPTwgqmJaC035Wag4ALl8ElkVekRk+piUIR1V8oE81fY+LeB61ryATdg1ECdFSHlB1RuP0qpsfK
RYd6XyWJbPi3dwzreY9XpcEVNz4h1Ui+RMsWOHll7TY4TKAQ6njYpNq06t06OjDS0ZJhfpVF4A+t
nnS+NIZJITvjqoXYBMZqk+k002zLC7GNitvH4ehigRhBCzRIwNkaweUHnWAWK2e/t6BDyXHBlTn4
5DldkTqV0wF8kDaUOPOhw3mU1oJ1ICNM8kqmFUMTbJuVMLoMGycBxILQ3qc58pTfPEk7djcmmO77
J0U5qm08JddahZ+oeXddzcSPetd1Ogbx8G/UckX9HraLUxwbpjY9s/UgfrL30yOSITpSXy0rq9Jx
9mHSYothvt4s0OEvKCBUtbhaFaSZbFOy7/OsDwELjiJ8o6/515uuaZ5CcOpGZSRfoOdzs+KC0QRM
HKTLI8mNJbTcco90qgwIc8i+rpvXrkb6/MwyWdp8LLEGH6voR11b6t4KQvDX4ZaCXTrqkXiwN/pX
oE7GEaEr2uhpLjs9xOcuG74HR/pgAEUa/quiYcbIw4crXDMKNgzhCdvP9sQxbHIqp/SVYpPFZ16+
TqQMOxjIXrgSkZZwZxGY+2lTUI3rH4nGBmcwWj5jr6yILveoOY5UXGuH8PQkkyxmpRn1xe6lHWyR
fW8S1PK/10yFOU2yq/DsmZQ/iwMqhvbFa0/F/vrjjs0hiocj7XJRsqKtHUsblFt5fDwj1tBObT8w
hCoqyzbzFqMT6Tc0w2L9DgqQKPbXCNxomn6caOAbsEUCcyTtuMRV5z7EkrggI+zyLT1PRYJsGo06
ZdGMIWyMYl61qGajuum+rHuP18ymP2Wammj80BOU8G/wMJ5iy2nAVsfa5NN7PWCuxK7qtLFgSDZE
3SDqFvc3YtN1rJ2rg6fDNuXGvszi3PexrXfhfdmkcGcD66TR5VNbMQBsV7UzfLSfVU1TNA1wQVEt
yNM7YAhaYG8PB/yu09sTrV8chCvca1rBd797PRMCqYesJq4HMQamOgBbysGNjsMCbm4u5FKbEO2B
UZMZHEvW8oxIVbkBRPzH47jfXfW2xYHYyIdRjpHawT++kjFjhZA1bz3e+oGvA3bc/6EhDd2tUrcF
xAkIQYhShm6qsI0d5Zbx+hlVtertoifJpETP6YRPzPzAaH9OD3neWJzCAFpMHmufR7cChwJr7Zq3
QPz+uQhdNNTKCLNc1s8Clkfm05Q2KAaGCf5eJ1RGEesmcWqBt+XxDsHcgrxQ4QtbFq1T2gFB3t0D
QR1LbhJP72+JO0LyuVuD4thsJ8DHbHzbn/jiHHw6mtPNeEWM8y+Y6muOyr3UnRHgO++3YGStTzV0
8nEY4F5iVcNUja3SczLglVIyn4L8smQNJcY/EP7CFkcoSu1VL6LcHzTpyL/9ZM8M1bIH0NDR+OOT
DFpOm62h/RvOuvpfwhM3AS9aKxDn+quWOkOAnI3Ht/EOiGyV23Ed9hXyU+B8fxPUFAMCf+zKOviO
OSAo90Kj5bVbq1jnPGyCOjp7vgYT7y0WDg94xGOc0HOXpztdf8a4Ztk1V8MVANu1R7VUugRH2vfA
JACYOdhjj/hQrfMNfdqYeYisCDmT4wZD39vXtOv0IhBGdT1cfv9yfjB32rKNuJHvq2E/3GGiWjZI
/489qnZE6hxeLYd2W1fOuc8D6dvLy65y4LX6N3zZKRLiD0UNDTKKDxKXRQh+LIg65RYMK7XOSKkB
xzLIiBQi8phUHpUlZiJD5cidqc2f6+8hCrvYBQ5RuA1asiciOxBdkpnCLzsxphAEcU8tPoxHPQ6M
QKdz+fD9e5hPQAWXGvtmUE+nS0sRkMYdEdUWfl0U3NZQp+2K2CEPZO+FrIhcNSnWGeVidE5bYmAc
pTibS099aQYEphZgxlXz2weNvRZB/waPlC1w/OsV8En5urN+ZvlyGvjYZBNspGH350Fw36SVRR68
Q+Kpo2aQEjXn3qerH9owsRTFbDvjVK7/lmdqOPABQYRmzK/9IffqMZM9vTX/NQw1q/6iSQZPvT2E
X9H3vbqV+u5/sjmS+AHR+JaBEFAtYizy3xN4BIVg4eoKoGr+jV5ikPV55ROE1BSGAs5EbhJSITk4
g7xH5007SsSynagZN5c6yEt6PF1zkxyj6j1l07bDi9RVv/79B/kGPnci1yU0CyNUfQx1ZXhUgtBO
dK8w+xX8recNy7laQUuQ0/xp5iagnwBBpBC3C1kakzqqau/xOVZ189sE0i0RH3s7Xw+kOg4lLCfi
c8uyNwxMTRIwSLzfErXi3Ijy00teCaOpCaG7PIILhns6hG9AG8LKXfZVCDiuYCaJW7aWeZs8Kv5x
d81tQVvqVNh98N/2UqzfdHHqtyabqEUTEg/U5QedRBhQ20ofeDkcI4jr0yKN9myzMw0WtDuSx7Yl
/Jxw7n8/CZBzDDFTonTerfeTcmbC6YXvWlc9VyTEq3TYhJm2p67Y5nf+TDwTJA6Y/QVaEgNh3LKU
ULXUrepGvpN2iGrf0HtJxI7A2bgcxBf8JnPeKv5AejKomeBIwV0f+Bhx2VVfZGF//2FaLQQpyw4w
Gs2Xg8Nwh2MKwbHE7cDyB1LpVOE4H+M5fNW9rkfIwtKDltJmFEPzIjOkRKcNLiNKnbKf//SCBmZk
hLcaPx64L70rSOTlcDsuYg1dIduZYHxFRZ85a7qr1Ch3SAck/EKfINmgjUY6ZpCo55N00cCytqHv
nr6WEfURoTR2KgqfhzRnFiFtVDWz1HRd8LY+JXRT632I1T6tmpOKmw1GlYtTJjiojPqXguV19i/u
n50f10WLOFfdrl5vatS/tGcgHdSV5PuaixEUdqZ3JKYTSh/8I/tNijlO2Ta/fnqkQlDe+uTIwp2t
6dtyci4xB/JfZo04MIUlGfuTTX7jq0S7AheQjoMG3BrzmJ7VrohYl7H1KVLhhQjiArTvgedpO+fR
S26cVl3ytCU6CBbx1v1ngCJZyfy5rsP9XSAlH3ln6xSodVs6/Q2HvGPqYCCdV/SQ/m9+02NPKRXB
+qrTFZoD7ZFlptnFnEyr5fLAL/C23FcSHH2UCx2tMwupX5MU5oiJn1c6OUzAxEuXO6BdB1KOT5Xf
3tNIHa+VczcbxUxLvrGG1vtLpca5oA8TYgNdiDUPv/rzqZYGyex1I5b6f03orPoHLx9+OwFJ+fc5
OFwZgM3eGj2znmuIYrxTze8tiQ1T+mTCu9EEDxiCNO6p6hKBRrjHHClI3rQYFkclsYtJ2XerCwDY
M+Bh0GG7BLd2L1tC2EJVwvEh8eNKNJ7F69BAIxfh2hyGUvifk65TE3MvWF2xLy6S1nidcAhmgcfv
F2HvmRfZ5d73CJUQJR30MpSIbToHXwg6OimvxH+o9NIBwayYVqDMltkWvtIHVwUCts+bHKM/Sspf
XSR7KUmuiayTm1+jIEvBXsm+1sHDqqQs2qDqeznlk7b3JCqIPGURwz9oVqFxlH0rGjw7LajzdhN/
DX3IrVfsaiVfoXq/O8oVHlCnMBTu7OxijohTNRpfqlEjKIjAqfNVCtcGNnEPi0WnVPyhAdq8GsNT
NvwqCkCGNj2XzQ1jIrJf2cIT+7qvUwqYw10eu6D5TwY8IEjFUIQ8ramxtxFKiEGMxy6jEfknx0xi
VFy9z243wcwUkD2ML6bMk9dmsITs31JznfnykVTsO8tOBIPfcfML7TbBs4nXDq6xn8r+dIU22lEk
2rK/mDhWUD2ljKTSPCdAS9fn1YYdytuc8PpveRldLpwu6pW+bKC/3tVaHSIbkMSf5ouvm8t+U3pR
kBGwL9kR5rVQurTyI8sSzHDZS7mPffKss46Lbqf97sztWOQ1idFeLqq2Atw9mcYRJK06m9N/FNs5
FS7RCCg5iGK4ABvLE6XCx2qBdmUnxBRxLOvFgs9E9Z7x89EKwspMhr5Vwk2yLUxN+vXub3u0fXkO
7xm+v2w3kMEDNCuZsqCTu28SEDKiYpzVv9EZamIQEVLnwqNOWfeaER/bVpSzdgxi0OwC0pe7WVz+
wuR1LMt8UzBmM+2AswT558M30XrobPSW+BnhpekKJukcCEjg+jf7HYei6Ty7ZO0FsdxkEm1Ojzmg
2+ZoNc5Oy8PQ6AigDB43DuWjDJz5xQ9UZFXNkaOa9DH1llYgrIiWmPd4kfLq3WWnDQbJ93fAPoKb
qwtX8CcWUSg/ZKHgXsuegv14wj/1lT9Aa9EfZDzS17rAOd8yOklRgFzWwLwqP8/8F2g9vvunjtKe
KeBaEY/Ew5RpNbCnvPGdN26UbZes3SEhJ4emZP0jY/BXK6cvZ0LRpFAbpg8QVsOFai6xVPE61gJb
U3+jyrH68ZQ7sHqTiGus+Tlo5cBDBOrA+UhtXu0i4xQ/vFtXtap1s4InCHbEtXGWLRFqYMQOB3Fg
TVkfVUfXn37is/ACCxnXBf7S6jqpAG8drO2w/k1sJ9J9+0N75pi3dOFmXItupOH3zlxYCMmdTPXN
j4bwyg93BdNCW5gbqRS9mC0hxP591j9qevedCqN97X7hvCXUGVM3EpDSvFvZvoDztwqEWG5h+Sw0
kgcKRjBw71lpoXvvIKF2IFrEfahnaMiUjXM+3JbOxqLBepnfyU869kgNfmaeUqgmd/nYdd4bbs3O
N2B3mnutXRSnFa+GRiaw5jwJuAfGkB9spP1btpF3R7GBRm4OfUYiFmSJuN6pmjq7FnVySkQClTRS
NjyQK7f3r1gZ9H2qzAu9RQKjAuBJodUlJe7U5Ih1O860t1vfNfd2Gh2/fjyi9nNDG8C7tAGepAby
2HIlZCK+x8JQtjrHUsnlOEMmnQlvlYSoqdMNqTMhZD+iGGu5jPBKFwfJiMIo6Vqr1wiPDmr9LhMh
1GCCcM+4hP+vY25lg4FfmIJt9/Cu6UfRi6+oZz3tKuJcVuGVT6NY7VvE744plOWl/p5MuBuM8A4v
LFMvc6xmiEZKW2SwS/Yf0wgTxhm4SASunAPtLJqz+aIYGORdTVstDNxB+fdi1eeKg0NwEr/jiksH
5+ksRKwMs7EOog0pFwHy/yRxFU7VkljF4z3A3DtLJRTtlpVV6Kln2/i4sbijsQ/Wq+bURpJm8chb
eOif2nBvdCvGbCFC12dU9wxB18mMKpoiazbzCgFapGTEvwflMT2AQHD5qu7LOvBghsYEpkYtVtlv
dWgG8JUNlUGiSAQl/jITEPCChngfHTFUDB1W+s4b+UjkVkPZUmckqFnFlqDL+5HIUgrSIpAziz2A
ibViYLnJrBLY4EjwVq0OjyyD/xL/8/zPkFMFJERlMuU4FF7Yk0gpjvfR
`protect end_protected
