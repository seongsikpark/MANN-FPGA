`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
kA+ipdqYRQy3NPVtmKU6jfwN4NIHjjLzgZ2O0bBMa4aMY/FAqM8oS69YBmkohQPtuczhEAEqSxEy
5x7MB/PfBA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
AmgJ7JpCiiivwF43M3eDIuboCi/zvH9/C8VvRuHE30yW75cJJylOlFHPbHAOMRD0dv0SI7/fnQr9
MaE1uNXySOVyESLF03UH8V0QNNO+Kr5zj02fzhMrWVaGYbFPD+cEw88WXFAmXCx3JddQEMgB6MqG
4u3bce2OyeED2YgQGP4=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
h5y2BoDynYEBdK/Y8MiwopN4nNXYz3CekEbTJmm6pppvfFImdL4EVOnGP34dJ79i4gOHoFBeLhVb
5RL9b65DiQIW/nKNTSu0inNoOp+IvyFmqfjERJbJzrbPrRff6hEN22abX2dTfFzom2ObMjV0kEE7
gAnpMdeQz29Lnew2xe409+LIGuyG5q1Bk7/miDhvSyCVpeSrejtjSZpWyD3Bj8GASBVYrzCRWT8w
SCi8Vts8rJr2uiMt+ZSwfimaoddMgE9N5ytslN6hIxxymoeoH7fDmWLPvorWpaXxzE3O4rddpN82
2JVs6fWtbGiCXt0K31Vxeg1y+7awXFjdHggAqg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
JoESiuc05geZoBgHD6/E4dt4FKjaU3E3jDbfEV77HxVsIKX9bQ/xTpEKUytUMu3Spy0cREwG9qLu
wY9jm0i4XavNWQnLrJ+SAJyyAvfqgmwnADcD3xLHN/BfW9g1K5ENK2yo/J3hK7OAZEIVxFGAYU6J
f4NhDBNOM6EiNIlqc+g=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
1M4FfCyGwD8F+5mMM8Rexr3c/KMPn/MyTiR4sfjwlJq6BSXkeGmGpwWWmEerpCFtIhYL8rD/p7Hd
5AxKORNGcAv6aPSTV+3sX+6WpHI/XHmdhFrVdpcyJyLOp6eC9PSTy4XvmiW7AISDzeLO3/Ww0FmJ
uSBkqsrYiavxEvC/MXJ2pElAS0zd0n6QHxsfphgL3T2x/s0T39pWzsbZp8Oz2yZusKDtzuvQTTVH
Sy3M35sIlqqlqh3uU2MTg+LHjEy7uZHmHSACmJR5150UtQ02ZTT0gJaRnljxdZW5/1NfuPS2rIvP
y0XaLcssR7xHms5iu2Xwz+/nze5c08hhkprOeg==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qEUqfOScMNowQMFQ7cnHO0lSH6hy+wmkM5OVdcwFiW/oaXLND528bwpqkEuSlHnn6IZR4bvTB6L5
uCqhY0vXBfD1rYt5R/CHX8k4QFv48ILkmF3q5tHibdwwTSWxWHYvR9h0ho6gSC+9BR2WxnUU4yKK
ti4pytetgPHcBF+KKnc6DoMztDOmMD5bpwKPiSgEtHU6k8dU94xXedmyg1XIZv2xneyaMtkQuxX5
O2B3o2duDCpiZf3vW/Sklch3xgj4aMTf0F9U+/HJ1ytw9tgZBPZ7CADqQdr0M922p1jO1uSEdlDX
7Rv8e0e0+0ebQ32zeE0v/aSRTNio8FDIgGWC1A==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 8912)
`protect data_block
48Ug2gTs3BczygN62ETfI0IMnfR3zsRoaUV3S9ASUK4P1e2AXbh6NnRiAg7TFg6KZE5mUuWxlTZ5
xN++XR89d6ySHFQEYVwVf4Rae0ZNw0iQqqLIYdQAF6xn74WB3Z+waFGFwlTVGaTMz+q4O22fIbWB
fqgKsjtPs/LFfScRq0/3fGwautsldwATk18eFXAwo1QqV4yjHxwQHkUbLw07Om2br8gm6VedQ+nj
4n+hk3gcXjEz3LsNwxx0L56NX9/ufiwIWg8hbvnWo8xiRwJcuQDtluQFdMkqMpd3uTRHwoCsR2/f
Cm5PevHhzw6TTiTabLs/8MtZ3CzKiALsnTXucXETxtIOKMw5gaUKci4ufYdWH4oNjl7HaqzYNQaj
vao4mPhbsyxBhvom6zFhyJCpg7aqqzlgY1yXn022NDO297buT54e7dbI+0CU03JLSrIjpd0PQaRE
RlKmT+ml3oa649sntxNyKfitmCWuCl1yZfUx/Kcvo6msvZfiEhzwgSZ3aiDTBnX1Uem7RVCjYlYR
VcfSMFeOn2lkCOAXncMfe9OHr2RjtYzq6yVDFQp7+foQr48+iQaf0fOJ0ovDP+XDmAzmsct4/1Ig
O818lI46pDsUJjZqJlNnRPCQ8R4gyDD+QpK2OOLudkjicjQtST9n3yxx5QgkQd29muqY4yUZf2xE
818g3BHaGCvqZTkquevHqGeC4Wrwt42Rq7JkxufFG983qIbZ83OHdULEiaJsxAxXZVvYONvXsm9Q
u7+znWsPRFD/95ko1fVUVaBJHKtxQ+mXrlQSAUm1e8UflyLuRB8FnFOVnbeDrBUfxurY6/FMRk/2
xevYhe5GJUEf6atlX0bD/AOcIHSJQkIfKexhdgv/8lqeHbWfoWd/PpbQvPhj5WMiiRLKGBBYIevG
Cw0XrYdFUgXV+VCmiRGetfu4BeHx4dP6R1fFfAW/CjNAbMmgxlMRz8ce2FsjdXfKk1FQ+IHZ0PBG
eW+bhhDe1oEfo/+qcUvcU+BuUlDyebcK2GgkAT4yHCckACIDFLU7UFR6XNDMd1WQDuCC8GZSpYXN
8xug7XRRUelZS0YTYZqJCVtUza6g1dcgKBWmbpLmOiLZgQ5w4+4kfwIeUlf9oTsta4W3LZpVAILx
AHi8ha6kuHMOTMuC3Mn9Gi86e0gkZ2aG+Gkt1t9yhugUxLOyTHHScI1d2KwHFcxxWz3+rRO4yfpU
IeIQiLsvnspNDr9KIrxBizfzcw+Oh7bPXzWN1B9eMjO5S6TD1EMnnRq+HVBJ4YH3Mwuq7kNn6iSl
ObUpdxS2CdvowbV3EGKlSlaK4DsrHOQ0s4Gk+HgSHn8t6G9ou9QvEIeJMPi6KV6iSSmYAO+GoNGu
N/+WoSg4F/3TRkdowiXh4hf3iIPW491rQF4oulr/OW+goo2QS9VucDsiNb2VlYimlOLL3oOpbqb1
phJuaA4S5/FcxeOKdjHkewWk5l6dye4EglnwemVrsz2/qy4gFxDyFa0Hc3II6pbxRXGQN0YJ7osG
HoXiujtNRgtrNv2Nu5dcx9G/3pCsfOQdLlEO/Zg/jCqHFdX3H7yvqrD+pp25fmDxf4R45XC+s71R
WV+uP98Vj4KH9dPClS3MaATgSFfPYmukr5GEWfIMJ5jBkHLQdZdYSc+XxZFi40mrpDoRZZRdpreV
1pwKysVEOdzzxyu9P8n0WGuIAOkRjwRW8f0dKB8bXN82MWUF9xzXKFdALpc4xURI7vMmsPhOebGZ
vlCAfcvrZy+N8iCt6Q9QcOgpBwui2+8zQENfHY4h8HWsyv9qo6yvIbxzwXnmBYbK93XLjaHpBg0a
MpmP5POIHrHPzeHpwFAJveu0i9kpAPk/SmLqAAVURRxeMD6rnRTnQ3zn6lkX4BHAQfM6i2AP4Ic1
VeUWdG77eNll/YtRSAup6U+mwfJDw91eFCD5DpKAOGUcr8hsO5IODD4tzlMBAoouTxoi+WZxrkC1
Bu4moWcUHJhRChNtDcsFNnvAmc9y+5xZA2dyid4ISUUZC5EqW0udwkq9or/1u3ZUnpAHLTuaFg+G
8/9gsP6JLJLSYYzpyzwbRBMRopq/j+BW8XBt3Y3gN5ybRP0x46U4m4Nbeu1lQ+ucJp6O9yT226Xy
mo5BqEg3ctESCcDVyPf2BYMAvPwORrX8x6qeHruQXtAJP/YC72sOM5Z8xdBTt0pxI/A7s2H/Sfrq
P5u8/KivrVrNJ638DAfnjjWyv6g3P3AhRH+mZ/lOYecn5Xk/UtHMFjD8gBN4tN782POCyMqeE3qA
vuOwdfDoRBuNeGupQmjT4Tt/0NO0rvxXwk1OEldqzoehPxrzjPlNtYWi7pG6Xt7U+c7qbiUkHyKx
/PXxhA9EBYuvphrc1PCDOy+JU65VghD8yG3Q/b3TkwFpYHgPck/WerB+Vp0biOyXxD5OCo7Eqs2+
BYtQMS4x0bhOqa4yyftNTN9C2mxcCEENm6QX7Xzdm3VF0sJm7joXygGm32eMshbDwhd3LSotIFKT
VzmkzdrMIsfV/IGE/Pfh8YgW9XAgkAI9cdZRd1kpJ7DkbqF6qBKe5Hr/sj84gn8KBfQwYcjJlLoC
T4M6ExJFnYJ0yRy0tiqOT1YclC8gKY3mhsvkTA4jWEwdbyb0EBgWlo12MmQUJ52kTiDKqxPz9LcQ
JCzlwHkB++WmEprMTJmHqnlPJI+mir9AEKsM7FVF/FlsLl0UeBC7H7QqDMpJCQRa8fJ7nOviZ/4J
cd81Fe36Rw2mvRf0fc0eS3zWWAzPRQuYDHRL0KGAUOY05YZGTAwUMTic1nQ70QebWn55hMjtECNl
2QaU9xKX/I9gLGm0CyFoCUJ2lN3gf/je+tAAfSB6YuXMtde4LvMdAXZAW/KE8czQkP7nbtKlwetS
inpmJbD1RaCm6d6nn692btQqB7yWYAtN8VHI+ao179XxwUjUzNFoDt0BBsf8+iDJuZBxB2V9rQFr
lzuBaTOVjQjq1R9a8RcGVlt1zNzi7+9GO+fVTRYlHuzTqiLh1hH0yP4fJPcOTuabjV5JqV/wdKrC
amZAL9sd3Wce097hofItPfmanZcPNWTOA4Fj/siJtdLqJt0JJJKXsldvX2C1jKRVHH9+h2irrGEw
PI725f6u8LYasnEuTmmxJjeU71vCZE6wAP7i+/6Ee8vCnwi1Ka/YgThCR3NlZJWmoD/lsY84n1xI
Xq5l6C5ynEGVcqCSAZTbAvtqtPhn9UVTqq268TxrWsTPrrmjiE/asQ0A97o1/h4xfpNFow04hffa
3TFuX4HHZxBPcAsGAUGRcLt02qYtm7JjTLjNWbMZIB8HAKupZZp2j7O13kJAJgJ2FmikvDaC8Kcj
ghVzM1yaNTN/INKAQbjPHpy+z18NYCnyj6YTfrACyhe0+3t3cBcWGkOWsLbEuGGA7v+yj3pAk8/r
Dub8HRDZT5Wy71udoy0SVJMHZpQQbq/LuN7pqx8AvGGVNMCuCs9wMFgjoWbJHizQQ32bTxL165L8
iA2JzSod2QBRrJBEUZ+ohxgpBOn85J5WUIT5OA3s0z8L5gpmeUfHAJYBgHfB410C7nwovYGpFtm5
EXrXoZxDvhHpmOzzZ5hgfuZt1cq6t0Bh70BGth/gyhBdqE71w+0JkVO2QY7ruSNGERcAYpM8QKik
Vs21tW/KuznxOuCS8XDx7dFthZivJMt2c7+jIdcQ3Zf7mTXPemRYOwtJ/fwu1TlWQvaAtPkInkne
NlzTrLyd9UTFEwULDP2sNn8VwXY9bUmMw0SvtUY9cnZmxYek14rxvgzP0bk6sCcehTReUKExX8DY
pCzWtJyY3FCikNEFtc8Aa9oDtolEGuiNhGL4vprjbe9hzKs3Vu+vhtPDUBohnmEqxNFjliqiSKVg
5R5o3N2NWefu6ErlsgC80AVOcHMKzKXEO9ma/NqCl5ubXCsUst6xGhuZr5kIReIcHj1Dg8RBCBjo
ecLhH59OmYfCvHD+3dU7YBEr6ZQTSO37KvTfnvf8DQA7DLb6I+bO33FD5Wd7lbf+aTaik4/d8Ksp
7CwaEndbwiaZe3LnaAmBR3Jnb2lM2ZJG8DvHxmaIPCQyIQFCfwAVT2NwTbp/Ist9QL2VUB+KFGb+
uXFybs4i/xB66wkczU/ywiHRsayQ3WPmgPXRYGqPgo+XH1Is8GtFGjG+xZ/maVdtLBdd60U6Y09o
MMJ+0xURRk8Rwd0iCedy3hrHTUI+ECv+fK+9seinerAqcmedu8g7463k76JhlwGxwc97yFIr0bUf
UAxPyRn/y/ze6zENMEAOWJ66DpQWdXNqhnCQaHqFpQlgBAaEK7rWsZ2YDwxzW8PjbII3a50hdK4c
x+9YHG832FDnjtIWXodraUTJBJlV+LUVyjAkWtKuB1KpMp4EfsDxm6g20q3zYt0qQmzNavHNnEJf
dblJyAsRFYCFupj7NlTRlQ+2IfpT1/abpTqtB0GnpQIUH+kIrreup5h5t1r+3g03I0q8DjawypFD
XfL+G8vcdE5cXjr3QZr5mHcphmf9Mo6tzgU2eNHbw4cZhl9+nWkjs54tRa4fubv6JR7d4KWyeCae
xnMbWvuzhkgTf7669B6grB2RxNn6A7ThqO/QEcabRDvucYPHhAaUufRYo1oqU7drxuxU3B/JVjXb
7jSGap9tyrI3WlCmS0rdqXt1sLpkRYziKbFAuPOlNd5cTTEse6peFnlMNna7asdLpePR4jOksJu+
jvof47kPDTU6dJJnHjZq5lyxl2blu/1F7L+0QTKIX/aSBu4PzeGJuCnqzjmUKEFvXxzGqu56F04E
2Ku8r4ZoMDfkScBy5/LEMD4ePPYMF0aPOPaRYtwn4ZPbcbBManxF/r2TiQEePxb744QV7i3n6OQ7
KGJ+UfaoMK1VQT6WrRyMNahNmZZwMqhv0g8Z04aeQ5O1Pbu5YP6NA2gr5m6+sU70FPXvgoQnQAPb
wrfVTTxmUtb9PIDi7zBQdjffW+ZNUVAhTfMEtb4SyQLiV0m7fF2jYbOQr4a0e0YjqforKfbAG+3d
OFuDON56iDrQ7FnihVah1x90eJg7gB/10lQAvicMqO7tI2M7ThC7rZ2jqIHMptwDOF25IEp9g6mk
Tds74PPYQJggGRDfgcHmJahWhO3CJLUxHsQf0PYYIUijEC+I/IM5Gargc0Cl0ea3pzSOerZm9xtD
XZnw7rwnUsIHN5eipyhGcr6e7i43G3WBSlzge2fEDk7Pl0UDgRfKoTUUzcPhp7u+FqyUAffjYbKl
8fYCYwLjgMRGhIDBqw9YresjW9qQfS+7rO9BQjZs7C4aehO7ZZCKl9K66HXa09GTYDGIPSCpXZL3
Bz8eaWU+XB5FbUH768xZF6bPMkHg7u7/iVKvyAq38fGWiNQkKa3tCfR0hcT+uCl3oGASvruoGFmZ
YCRybHQMFev5C1oMixzqcM3vQVuMsd1oK27BNwjpBgnKGAQTBk3ggDv2pLVgzJWAfDGTmEv+Tk/+
OLwg+3ySeMPRLC8IWllQ9CwKB4RvyYjjjcyvch5+yWVIo4YcwHIvCuCTfwkKuET2BczcGQj62VPQ
pfcPYqhSb8hS75sqEtfhic7YIAqQfwAfnXOiZ+QXkV8KTOtKG9X2h6IDS6yZ4BC6TnlaJV/p8WDG
QkowA2vua1taYdZl0m7hxaHzzDjaYC7Rqp6YUIUe8P+wigt770BfaNQ9TdIc17w6WuFBixpGJYN0
oNvZ2b7PCf2VtzNO39OV/Y40Gs8PEZ+MrYWO3855BG/eDqTkX7JLvqFxQ3XdHc4/8rtCkoSb3YrB
JSlJa5GikE+eoI2yxQkERXWNal7pYmpXa4bh80212J/im7RARTHAKFm4ibgafoI7yT+wkIV6Bqd3
8C3tZrWGUcqx8kK0z4Kp9MWAWaOiOn7nW/jgwkvwDrbSUs9BXWfwl2L1EMU5wO7CgJvVKgfevktP
Wdat/2r1OI8iqzlkg6lOadZmzkquNZU/m5vYwXhPOPJcFaPZVxPH7IGLh0UrYKF47wlZvqF7mqhM
QyeTRKQieyD6iAJxsyPu94hqWDy3tUk1SahJxgiz7+b7K1fnq7/pNpW6Dh7tFpl2AEMqLaVhUNeK
hKOV0CuSWgPIz5MR0V5CFWlCkzK5ZcGZWNTJhqKfECO8S4AKAnCGnyTVBrkpK1jhk+7epXgmOCPV
/gVnhdwaFCqMy+vzQKXGpZb8+ZPfR6TGgqqXp8T+GP4lT/ULTo49Fw0hi+gVw/8aD5udLBR3bedR
I1bHFOByL/v6T52fJGpxRcBLRkX+GW46q9oXcblYE3hMy9ZmPL19/1fW0O33qnbGBz5QXuOua1aG
Mf+iNX28nAX/R5fjlmbh9ecBkxoUhFF1Ds9Ij/2pmPGeVDuYwPT6pyDZZgGUh/bcEI8JJcfiHTO6
Q1e5Wgvbiy6rOXQdF8fy+MuS1kecugh2RfratbOgUXeSJMYRieJcQyZpZatfB2KhL6H3ERFCqMCs
EuUmhExSqLeMJWDWi9pgsyLJzyuyWuH0K3y8chO48Gt4HU04pqjoDs5cD1BP4Jnbzkgv5ARTsHGp
5f8SzIWQaNZSXzycJVXmxWPa8c2UgA5+ftvlgzmebT+GbY3bJtvUyjkviVowgeeJaLUJLWtqESgB
aRCyHKvn8Gwnz/BxJWhpeEKYdPBKF9NxNhdQyKPdzwNBeJd942+628znoQavQeu2xWGCQcrt2pCd
L0jGrOyPyzrMA0IdZx5uK8GGH5N9jA9xqTWVn/gfqjUNWpf1V1/qukf4cf1jJ+rvIUKS+oTJhULg
9invHc28cPL6P05bQlyHG3DLuFAgED201LlVW8PAIld9dy9tvOQJhPmikXcBola21QvLNnNbcLl7
UpCturkAriQ+7oI4gu2FTgarklTWtJWKf97WkRgV5LtZx5GmD4/pBS7UY4FDj13pvvb0sE9aVkDC
+4f+CkDwZSe33QfRj+/XNWhvs6GIUnBJK8TApJ5wyNK1+5Jmog18bjBzcY9jNsPyMzIP0z5b3wiB
07o4DMDySRfus8ePI1ygD+nyAGE1yPzhLdwIGYEpigVSI+LUMfxd48cV6eNI2lsiXnbwKIQJcsR/
+4b1MX7ae26PBge12yvMHXwLUbiPOqh6dNbjpm8E5nL04KzMtHrP5gEhKafl4AsPqmsvzzGyUiaw
pFdtmDhQU1y7MLouuFMhMk6C4uiAcrpYkExGGdmqAEG2jx7TlLzuz+KB2/qE6jlc7rvYGG+hFxTH
gY1UuJ4qyCZqQB4IZasLpsqaZj5voMxtuFuuVZnTzwGh8DCERslcFrno32p+a6X3RqrOW+1cyQIl
0aGxXotkKyq6AM+3iQo04lu3NKWkP7WgREr0owDCY2Nls+WFyDFhpEnZTevhtET3Oj9ljE7AU513
oQnB/0ypSrwE9qw9U85VpqFmPlGz6Sg8hTx0T3OEjJoJW5JXwTJCTQ0FviEVS+uwntLniYd8zvvE
sC0SQUv9bG9a7FwfDJBTKlCdQ0bUc00pQmgyb+9MF5usmctPqcQthHzJ+B9BN2HM6i0cxGf0HGOe
/yVCeQOrE8sOoaYbuIc9W1apgmvRFzqfWOLgFDsU68u0UyC6G5wfuJTxmbiSVsHI4nWD7WF6pEGU
4DimBicWn0C5f9MG04St9g306V8uPCC9E5vm2pkWnhM9bUcygra2eSArSJLXKXP6b4atxHBhuz8S
1rPYqsdtLs0ZIDAyVqsGxDqRn+zmFMn8rRrK64V2jiMF7/NUIpKPHZ1Oxg607TTT8yg7PRIRQgdL
XBryWk7l/Cze++vUreAXewi1ESXTUyEjaysMhPqLY3av6PxBiC6zWTkc8WukQNLTorvpaEJkDdUV
bzXSI0ATKvs5tBvOWKA9YOZDQqGgyWZdh0ZnMnNPD8m0LYFPoHSrYRlrYhnwn8rN8w1C6RaJ9qGw
GDuLr0Z9/xHKPZyc/e2FK/JOCMM5zryIAsycSad4WAD5ccHZ2eNH+PxaIP30PxTNvA62hL8R4UVy
tZwnmHDq0QTQ7I8OtqDRkHoW2rgE762YncV5LKj+VAKqnyGRa3E4xge2FMXon1CVnz+2wnhQ3Ybm
p77zmmmBcIrkLLaON8u8S0A2jLmYfp4xhj5JaE2IZt/WASDLbzUAkIuvjFhAahT7vu4oc+QCPCgm
Rnpk/tDc79v11P3qYEVb6BvPRrxPTX403xSlWWqDpiey0dCkkfmPiT2hr/Jqj9S0li3my2yIv2pV
Aqrhu/2JIcgSA1EgBklDkZKe14Oucu/gYFM7qj5gPss0Xk1v3o9Rl/mXjt4aIAKio3hU2NglxFme
OqApJBOWYl4TArz5Ggca+AWz3S/OpQnOM90igz+DvLfRQw6hGEC73BUa6np6NQhhn7q6l8EGsDXT
bjLgVMh0y7pzDkASE3EpryB7wOeMoMcrVIkqWs6MLzgULhWRqZ6QfUO4Ig4ZX1Pp+P+FKp5cEWB+
kaXhxh3t+qFGI2T6E880aK2luM9M+0rCu0s00o5/JbzVyA5EXyHaDXHqGf9ubl21GSmKNwAMz17U
ACzROvuvNc0FHi863ZxJde61ESaOZ+sWdtyRzc8U3mhPhAdhqycJQsrUC5ixwD34JqeI3dAyn9uB
FIi2OvYM6zHYrvIo/9NbKt+lo6IBh3kkT/TTyoJZMulxG3KIJ092PfrLbNKXghqY7VUNlgiRKWbM
y3aWmQ/sYg8zeKawMV2Ir7cJS1LhEfeAaX9+SuUeE/34zsn1k/VzZxZNS3wsEabvqhQzaYLQo+fE
j2a4IgHpy9dNEsRfnLeAndCKF9/tklEB0JxjDJcGVMNxznUo+z9T2SC174WoRI58tIYfK4GmIb9l
SYAwSxGuE+2NhHIOacMyJOCbJxHrmHD70rcOUAgj/60fRFk4T3frAz9PDZEHiDjQpkSn8OmTm+SL
5heGqRM1w0w0Kt28B2oKaGjXXBkhwQGE0ReoL0srmzXOvp1SBfbFdAIMUAHYb/Rju/Kobp/nyAke
W5l74MR1mfsvKxOmuOPVpyvmu6ohPzVQCr1FtvUzKAXcp//cYUkGZRYf0JdtIgRgnCzAtBpA2o4T
JH0fQTM8nKC+WlYT2J/CVV/5wC+1nYKrBrdNrNCCCLmLwqnMvEsrXA7lk5sLEGkdtT5nzVsbdFxN
jhjjrAWpL8nQ6aUoy3hsnmJjBjFeovbyI6LjgPH/PGoz1GHJmA4ngZsez6+2ASArED4khPfgWweY
RXIqsM3k/sEfKGB9ZhEAPClMefjath5Ngs7sW2DmpIkAvAFquxu4cxiDC39dltjtnUpO697XJPuL
BV1yLTehSc6fD1tzyntv6cN2pDP6k22Yy4ViHfSMcC6eO6vHGVvxqy7LTmWj+5GITnvBdvORnlQy
vHZv1BsNmvmIxImTZ+ebJLyMPbEjIg/iT14Ejds51oA6zxMSAQJWujH7P3kETMaFRqPbn5+PVdtn
903fJasLdNiagBlRiM9YeJzZnuxY5f1iJCI22vOcgFVHMv4S/5WT3a95ynJviW/kpP2XCsJE1qTF
ZoipMOxUasszuc8BDUUO0iiJUAwTNlYRPPCsiWfJIHMonKqNez4ATL7xmcSZeQs2KT0DeCakoyb+
4NCtF1c6S8CtMDcRFeYW77CZVkanvDz2E0wqymaQFgZLiQ7FHDqCf6p9Oyxw4H1n0J1ldBy6lGFX
rdcLA6VaaECPjje1fx04PDMxXAzbTBh8i3ELAsAXw4ZaoiS7Tkm/TqM+uUHyi3+f4ezh3dMxTZee
LoP41oF51lpFJq0bSwFG5XdkjxkElhKBdrLzYrYaQawHu7+ArHMIsNCfV6PmJyJKostD4Z7Aiu+F
VkO4HBiewsmWb6mbXoet0updXV7FeS5UQrmv5d7zHRRahLVwOni6KL/IFQK6pc3pUjozIiKNGipJ
u0DvPTBsiPrY7o3vHWpjyv5bthxIRJirsCH/wktAJiElEn5PQDsobfz1qOJVUbVmQHItqM1y0yXx
L0jLAFetCM7IsZMbbOklxn2WOyVeNFQzbWxh97dEMHNQaVVD1pE2x1UXo+vQj83NiKLWgXCL5wAB
IZOynVEyPVAah0bJveVeB14MfpckKF5LtAmoXquq2f16qYSGFK/joNU+Ihh2mkgKjt3Z6qO7gTvA
qB9WFW9WtDqIHdg0QzwGQqCLtxh0/CVhOP9qn2xJeF7Wci+OILsel8uyZjrTEO7MsiGVKyAYJUUn
aFS9bBiszKDRMueVmiPg9uiKIoDWiTagkNdT3hBPBRQEUmsbCjG6FdxlGykKMQVBrgxcFpFgOe0+
z4b+pAgjqTzKbrzxY26paUhq8I2yHGJX6DDCPjywwd/Cczj3HMcJgucxa1RpGfePUZj/mkw3byxB
mp9STUGjaePV7jsHjKTu43DQKc5D5lvFF1Sd8A3teDvQgg2UrfjAN2SECDgZScfSNtvNw7Ji4l0B
oc+ppUi1FM1rbnjTMBLwyMhG++GVz6BQwc20ydX/U/HYz0nUekp5lnnheCRcnYF6B1vHbZKuTjbD
48zgmMQ8+D3xjhWJE22v6vWP5y+HyQY/+jjinzLGYwuEvvAie8tzyowGKvPBrv6kqHOh50dXiHRq
mCLPbE80Q2AT3n9NetrdLBr0huamp4HY2imEafiOVT+2bC80MAuBXJqYaoBusRXzwgJbt/GxUe8D
lXbM3Y2gWH3wAl0a/bFk0/LZ4PAUYIyAtVzCVl/UOyfZATvJdOR/38WeYPpsKOId8m1eC9+lMbuf
v41H6cQdqNVo77h9SwIZTgRej1uN/mdmwF6xHMUdR8uoSPx0VbzLABSGTdMWvIEFmyivII6i2/Y7
BLtspGoVGzBkQ2AmbALYgY+77lia7YgivMwXvk7RNlFxgtnOAgkFbBTjv6lVOZIBCe5hwh3z0945
yJgZcQ4ZE/tJBrU1Y7ZbI7pCKvZt+cxWm8tt0a3/tzKxxRtLGmvrJ8hIpY+s4qaKoeLtuOtIPUYE
5o+GclKhTJ7ZU7Uc4zIRGSK5zeEI8SXub9kO8eKZCJ1vQNgyVKf6kJYDqyIv/6z3SxXg/Rfolt4v
9Kh8tx/hBXx3B+NDG5oZ7rwoCU5UjlSwPIh6zRTKeCT2za8tqN82jrgknlBnmsPyS9sSHZJHU8oc
vPS1J/CYzOPANnLE4OvtAQpR/rNXLAq0zHUNBacZ32xivYVJEiRgMpSQcYjLrc4E2SjXzo8OMYY1
fpaxpxcw9zBJQ93kVwGXBMy03y9RvUB8leqLK+tgHM9hwcag2Rs5BTbKBiO/Fxz/jwbpXkvBMYb8
onlk85Dc8T5qaZkZOhstauxBoewLkkzpUQYE0GQJUEdpSCoo5H3HeTh6sqkJXMOnJxOJSRxYU16s
AaUCoCg5CXRcUCFzkM8KRPTw17s98ocgZVWBUUDnCBdbq+zrIjIqhk5Ckc0fbe1l6WLkcSDmHSzy
imYBgMczfHP4KWjzkLwFochNSB54Je+Elx0r7K0vad9Mi0hYbXwgKx8OeBTI8NtWxZnGFtfSnep6
fKVYOn1508Wt5ZDMWHis41Wo6DDWn1RJFM3Vcvy5V7kw9nFKEHMMwNnmhJNx3C/+MxXlw4OxClYe
W2CSGEJutEIKW8HJsTut9LEQacJekthUV103Kf60RSgkLfLzkm+BI8hpD5M+33cVjebxdsiKgbeq
Qtz3jv9zrFPdkT4yHV61Ta7T/Qt8QFmQcVLhJHtVRo5+BgJ8EZL0VSbZcF0Nbw4QOXRKNIi8lNKs
ED2m1dtHPh7KtF1Ty9qUJfcNSEhqFlG/emNXNiGbwuizCK89XPHKFBsUFRO6vWh5SIRMmrzs58SQ
LeXXTDmFOvCKG8jCXIouk79AJiqdJDttATyMmE/K3QbbMMIkjvLjwG+/0Xk0bbhxV2r5mryAL8qt
+I2/Q1VSlPbSrq2UD6o83c5qDrY=
`protect end_protected
