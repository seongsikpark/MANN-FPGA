`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
K6MLXsHy1mE/e+BDKQWWCf+4ivx+zNnJ8O6cBeb3pUw6btsYq6X7MtHOz2Oz8HDGPA6q9x8lkpvp
HcdJOMY+HA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
P6xTgR8Sldnm8Q2SDl0KldP8Mxalhk+FQ8DKI5wS3in+vTjwT+0Qnq+F+NLFFYSjCVLQsvICID2y
uDTWUrzC2hBYfXhSogTyPkvWjKOEUhadOtQFmXVRiaRRmDsmYIP0VfzBDciE/+KgDZ8IlUPPc2cU
WqlOcJ/eLogYE6zQYMI=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
QdKj0eSWfm5SMookhXL5Mfkv6ZPZaxlVqSnBQx6Zt0SW9kTejDuRAfDQp4EiCm9dC8Y0Q5g8DAto
xJWkPZTunorz0KoMjqzfZLgIPVA5PGWbf1yF86jDL7ftFfK1/8E+/7kecMymdPwvYYkrdFLOrl83
j0kjqGJFjwWrjZ8CVV09XjFElDr4v/W+DOpUjCphuOH5LKetNJs0j1z+JTO6XyruGaCJzAbl5xfA
R3li4pGfWu8XeN8gITkQImYGrrJF42U+3XtYru5NbH2wQlg+/uqFprJWP947IwURkztN7oj5DsqW
VGP0FCt12yKYCT2AceNJcCSCSfsK4Pc0HB0raw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
mPUaOpmvmhBtVYCiUSfFBnEWc/b/39RU8W3MPTyFNUhf8hLULjpBea+PhKmrbx+gPsC6jLfNd/Xy
itAaLl+gJoHCpcTd0fHd0QVx5zBysFQ96p8lvwTAzlgiIf3KJfmwt8iSojdq84xPq65iSh5WwHu/
tEAPVBe9eTqEsegw5OQ=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
jrmiVyp7fll8pzeg0coNDePx3gVSGIxJxJB6Bfv2T7tlCbnb88FAvJzHLMoMUWGpWm5r2zw8eCKa
Re0+GzIsqFVL4pR1zaSSapK4xk4ypME+FriinPALL2yVdhs/1J+jPO4gjFoISVOsvns5g2dSuY3P
GJVpKqvQHiraQr52fdpU9xAyUKpykZT8l/DaSAGnjzaVdxVj+HEfd2wVvaJm2IxmKgnNA1zzVFzv
P08LRfOwoyCo4MCVekMYpFXSZriE/BwYHLhQ0uJrHSez7UD9w9riANFGHIoCRiRg998RhA8HIHyB
SviozKjzIIihOUGyb/M6tsh5Yc/fya86iklPYQ==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
KLs19GN1d72xAG6XSs7/+R2FVv4B0ae56gDUM2+UPaYIMAruFbPejUIaZmGcPW74627oECmrLsqv
yMhGuqy2Y0ZAH3mvlDb2l/KsIFLZJZNfnjHfIqdh2ln71HiLa9iLYqMfDqFpjbsNmlibkeIK6Ye1
6tjFbBzcYUfGzxxN86GVKIyqUC32+XUgV9CY07BtadF/xu9ANU8romdQ3zqjalL6iPbVHMGpO+ri
zswv6sMOd1tX74Na1ibUuhZG1Pyqcpbo+mRkfRQN/QptsqOS9K+PrfdE7Vhte7nW2/xYzDgGdjP0
IIGZJzDtIH+iqkAC+Hw6/elB7pBRqkRDetaGzA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 65248)
`protect data_block
m32k8HPm27Xy1sF3XgmUllWh2GeMCSuFyEjY1hzs32tMeNEpfAZ4Oovnq+tV1PWWha9hRdAuo0fq
9oRGLvoZ+NRQ9MnEEFttErkOkQrF6qf8ljaXF078oHU8eCB/Hn8t21zeq2zY2CviqSv6xr8Hk/eM
0ou6s6anpMd1/aTvbftJsKp3Z26TKoGoCtj3zhAFp9esUUZx7LayVUjBTZ8V4iJrbOUqz5bRcPxF
qM2UvwjRjJ/WVhpOHmxKOCqo65DkJ0qRIzuXj9siRWZk0DgP2Noc8VO+v4TStF5SrUZ7emglm+SO
3zgfBnesxNSuozU65Z9gQPWEEuuRawsd/fLRELMDQPWuZSNXWuLqGMBdp+0xRDLPr7xqNELSP9kI
y0TX3bed/B1D74qMMAuSng4E4XzOy0f5PADKkB0TB+xGMtxMYgEsrVTfE1VD8jA8Q1+y0Y2nx+40
4DL3qLOKO7kAjRK3455sfB4vINpBaIYr6p3qWwErocNOsM8skA1gWaHePwuswTzzd9DE0uGF/Aen
0nhpq4suR9qPHZNpbQ6Es0pBhONOMfLYvCrYci7bXmefdBalfkb6+RwBULx6QsbnIQMvT0rbymEh
eSi8gaNWgIPK7EBj0N+REc7xLCa5V1GghJ5vK4GaCmYQ6gPw65emi0qJOzhZ5Ar4Gs/Mw751BGdA
9u/1KfSGLeJ3A0/KfvawzSL3+HYbIC/bTTCoPnU0HAj8ZA7yhYRpqW+GCxZBox/l9JdqSygIDnXG
KtdXRnLAuTzXq8ETTfXbEdw6pxTA+JI1UU5dkmmL2uT+so6PamxjpmoFQBLHDi1aA1UbBQf9LVsZ
k7PSTR4rDerZk8Ix6OAUEwVin/UrgsGL9HgKxLkDvnyi5W9BxBJk2mOcgEDMFDzf+CMDKm2qbg7m
HdHut4oluVDOfNZUnbNgW1JtNaRojF3/Aa9nbIvF809jpyTEt2zgJn3KNoWFHWVztq667uHr0z/g
CQz8knaeztMyrAXYGaSx8QStXumM/srA0X7MKHxYvgwK85NV7ePZ0NAEZsWv4rCMkIJSH4T1U2VS
5QF73qvQUyzvs+V52SWEwoOTIf6sqSYLOZQHrl61EDDdamxCa/IqllHAWhYVogVmMb3pTOq2gxFd
VuoR+epm32sf2AgJlYZO0C5tPKJWav0oxsInOFCHXeZCdBFDSTpzkJe39WFFruwCrbrw1z7nfDBX
MG/k0GFg/RMAT2Plx9066vpq+tn+Pv+LXMxqcBqCqx7U5DQ2xOk8AI8/0IXQTrLvWz1Kt5gIB8A/
OQsZccZ1NdP/nTXFCp92tGqHN8TKNl2ZpP9jiNdsAzyxpzj45sURfeQQ+QW8aXazUbCnH8LRHeEl
JeekC3WgBUnKaEUSu572fcCOqyJgiOb+iof5t3VoooaAFRu8kDncsqm9Gs9zqH+c4ZmERaJjtHhD
w8cAWkYR7Mx+fOtW230ucb32a2HFvzeoB9n0DOu+AgXeOUdHW21RJJOKRl8JjvFJsYcAJjrGfBBx
GjMSdv6JTgJvk72PwxdE8Sev6HQcof6ueKQ5qEpEUUhkPZte6oL8ZB74Y4T39DFDsh3pCWva7VKJ
GMMETrbaobZHusWSMbB4KA0cGV9pnVZ6xFBueJmJdX/HgSzUuw+HfgvJ11miDd5QBHcaL+veQ0dk
f7GPLKoC6HUfi+sblcj9zvD56Zh8LES6+mY1lOgE+mK+MYUP9/Ige/2MUxpFsobVlKaV/lWVmfmm
9BPRp4lb7bv5JHoZAnVPXp5V8z2cCJ6ZCSO1JXQd0wGxmDmkK3p/oN7RJLZfJZlKitvxREfHu3vX
VE8VIg/lXuaDFpcfgQwk5Tn6raPnvvIoexNoJKVp9jmPx1KGegPpUfFMCfva9730DKZpIIvSbl+f
AhEhirn/MtGxd851hdFdcHzswAtAcEsxaSbMtpolpQAw819VsO7I1+cD/Yivq9wt8Q6Ujo0Q9L8x
j6yAmxUDF+rZbN9Y9RDZGoofHgWlbx9mURjImjC9MQ5ljwl6QvA8F+deHoLGPi9gvLfiq5zwc7Og
ojy0cIcfUVL+/yqNsv3HXUZSP9vONhGgUs+SV+DcWw4DJf44zOEKIh1zWhRcRBlMOFAZxEIuIS5l
W/mvtnn9PYLmKREHzf4eVKYjTQXrEMSpy1a1ai7o+Rz0RsRb5jWyTVoa2BPn+vhMtsmy4fzxDpLG
+2oTQs3kKcmpXQL/L9LQf3mPPTtk+Wqr5FFwYaglhUiM3VjbYbK5GTUeDlBoR5Qkr8tkOcWNSkVP
p4qrnOnI3DQ2use4lXGAFvN2Yn1mc5ylEz8lNi06TYrDlgQszjG2KZB2WG5jHrcJ3IlQxV03NfFv
PYUKz7lrrxPdIY7ZxbPk3Hu7ppZCqzvFdz3f+66GoJmJWJr7QRvLz4EoZN7H7/Rk5TyuM5MOfrKA
VNR59y2Z0nKxw186ntGKwuDoIEd6U2FyVLtilZ3+7v/QUR/DMpMTxdZ9j/zux905OWRIV/mloIKS
JD7Q4ka1qmMomL7yAc/1lPS3J00RqsnGhjUiOhFiHjsij+BytDRHk5AILvVcItTwv1VqJGAalOSv
0fkH9k5d8UqP/wI8frKKkijOkC3cp0AJVMyyZ/9PQ7xDU7dedoSoty/tXqaW56vS6wxhAqzSmA49
STVoYR2230ngR4Gd3MIEUeUr1q6rTrLBSOaTtouunQ52LsOmGLqeIKvWl5ACwFgkWHd9PvUedKpR
8I237yi8KjgQXNX//AbsYEIH0lRkSma/up9U5pdPKeZwoSkrQRvfoa44a96iUR4b4nwM8j6biG38
Qli3SQaXfLxTpBUx5xNN66TjytC5noXbBOLmwVDUWDmQeNod7XtQr2fGBmGiTZbDnMICNve6Q0vo
JL0SiWLo4511xV0Jj8Mm2P6i03+deWYSBcsjrCNoSZ8Lt9fHvOpK3NMrw3Pl8qs7QHyzgeM3jK4L
nfowfoBS4DR4vgKZjPTPUhmF+OP2nHCFpqLCoUcliryHu4HOMBJEt1LFbUgui1zNUeYvJ8k+jvaU
Lw76zgdfHYKI5amx624LGxMVDIN3wOr4dKc0yMm3BWSDMT7RGpwKGbmZA5mxDiSe6E70WsXjW9zN
VuVRO6cl2yrbQrganumcAJ4CkTUDWkhoadEW66qGw9D9BeVTqJ0Av/+gO3FRR79nt72tQxRXwGnB
eGadn9XQUpMFgLOpzt6lgE3BEKW4VY2HJbBqiiZfMvhaAKA6wcAMkPr/u4Gi1uRyFXhB/FNsF6nC
7zekAu0bllWBf6mDpYsO3vBIC2q0N3ywYU6lJ6QlVXRspklIoEiwntFVlbyBtbmToP38d2rKf9r/
PPESfnv3zy8naRuese0nUi9EfiQtkrjjuIU2/TcGq4AetMBxoKCiAllQyOutK07n20uRlPHpZowj
d8jGbQv8DHAQVrB4pHkSWsSSDt3c0A2g+u2gMwS8QELpIj+6bZaGycxQ8WBHDEYzcTUmkTUmxyHF
GZyiUmCy+YP1YvTp297OnqcA4TwyPfLHYcm2XIBS1ZTEqP3LiEMFl9v1AYMvTWaOxqwPxAQdVWqX
32PWQ0Z6yzO7GRsvxjzFRme6cDmsNtW+6g7K8t5D0qP1AjEoOGgg+e+AxiFQSQ7PcThpzj89qawc
AZ4iDhSUJ/Qw2YVrwGoXni4JnG8zVYyNPIuCH3mg73nzSWjcUpgNDf0n752yjEFcDpLlWOqIc+23
Hwpxd9ZS3QxfZ8Zuy+H7+SBCQHswvRNJYqbd4NH7+TxeajIKi3voKqRKcxbec7nD767/h6gwv8t1
ttSMekS9fbqCjpxnttHvmEoWiTfPNijIpBOhnzscTuSyY0yDIxCh4+BRvsLn4n7kC5ZT/696Zaay
klu3E6Kd7l1bAimDlVYKv0I8R/kp5ujQdjBZyi1lrv4gdIf0VVLHHnsvuHF9qtaMu5w2VV0WgeHt
V3ZRUWEEOz3qmTEPTbUjJTcrXA/hg5HvjFPT4Zy45/HfvkjWOiRS1caARxPc/kxH5RW4opRbV3ju
p2jXg0sh0oYndxUCWLWiXg+hOntouUR2MV1MZ+hFEMkKeE9ekT6hZGoWp//vxEWoXl61j1iL88Yo
aqqTbzaZFY3bzZGY9ExShe2iEC/Vz3NcNd6U5lwBgmrhD6hj7Gy9crdkkkxc36T+gLijRhXbqvVd
kSW+Sim5ZsEzE+D2S2TAM68AfYfTHUuWoDxm+uYejH5HBl+iZjjCEebMAJrZKQy5UmD68ctwwMSY
QgiQCw6vXnhdYW/ikC5ZhN5OSw+8q6SbLPaYKOcUearFrYsRR0wfutAy8t3yumeLlmOHgezs7KFH
Xpf7gptkBZLxWaeTUwiu3NjuoY7QVsftRtzVm2F5JyLtVRc8Acw/1Smm96MBOjxtBOMEk0CZaWQd
ZLk2CQ6peAZyba2BFx5E1Zxb1Ta+A6HYy46uttOYP3tPxL1LotG09WSVOoXH8tY2kI5i8xWYMXmW
Ih55e5y2gE/ws+HdVPGsVnXzcVjMiV01Ff3Gv1cbjgC+FPY2WNmfNqrkJVayLrOqUp2bsJnZ6Bmw
UW8XYRw5NaFaT5CuBF4ukdUJw7JXQ0NbRzR/EwTiP4jI7gM629uOT8CHmov4gnr/e+H9zDeomMFv
QtftRUtiGHzBxGqexMZTFGMNh+14+W3Cr2c6zYen6AVfcnEB1aRNUUIBynfcJo0oU01zn1lsNqhW
9eunYNZkSCBMcsh89d4UP1FPofSan5m8ws16ygt3F2bg6K3SvovUYlgnTJhCjkZK/+nNtHl2Mk9b
ygI8SbS+r51OlSj/x3RNjfmxqtYg/k1PPcrOJd34bKYkNEG70fchVAPvofT5CS6QK9b+fRvg32bB
9+H//8WPoeLXN6ta+kR8s7IOl44C6FER/tnN645haE436OepzEdYLXCuFoROXK426nTsQvlIcEL1
W17mMSbI9aw6WlD1UjFx6k4qMF5FDAhje/8fvdkWPczxa566pfG6W8JBOs/GLJlqP8KiwnvBE3DV
KDCVWXeNNghNCXJzO/pfmir1K9ZDexDEBT5qmfXuByxEdur0RzIOwsz/89pkiFnnL7tLZSDVTrR5
Cojt5RYTzHU8kGAX2JcZovbuavLSBkSjfm8+pteAKKZKqP7unBhwZZFHAl1HC58cTC1OVUbKL2PA
BIMtfe/bYrBpOjUNR5T3Hmn4LWexJlZLVLralNRDtVsHHqgaC9PATmq+qWx7ISduQyzWJglNrx4m
nul9CbGm9SQyBRZhfGn21XQQTaf6KTdf5MiHNaHD6wuA25juG9FVt9hg3bI3hcsaEkvqGRoYQKn9
IP1lwOv/JqJBQejpaUo+LXc9Qjc0g3b5XXdf2SL+LrFO5Gi6afKKigbwZKC8kxYzrPxJYyizPAI3
K+pyH0ft+UDpxPkpjexXttwe1yVQvj1SWudXdkasMVJMvcRukkcP9FqtQe2UZ5dZMvnSGsZSpjnj
8P6PFgHSIusRqzYh6jdDHvigxFqqPaEf2aG9qVU70ul7nZU2F+5n1Kkx00Kvx1eVynH5i6FKa8ox
s8+xRWLkRR3ftMcv1cmb/xO3YdY11BwyDLzU5NsoBfzIOWxVS6oryy/G8BbnlRplZjgc3qDjSqqz
C3jlmmZ7Lm7op/aT/tEDfhXXHJ2kMK3ROuCujy44ih0/mB8orAjR/Hn/xu9KgrKg3ALqWFrSMAaL
kCs6W5CZ744dy3fKc/R0CiEiQViMGr0LxurdO3e0p2xvX0ZdoUQKiWHbiBzogo0mtb7s1Xnvf0op
EzFVIdzCi1Sa82Xcs40QjcVVv6akmo7nqLd3zawOwZbc/ZYAIpqIbQv3wWpkeuE6n/SJFjMkZpE1
61mZqtMQtMJsXvy43iEOfTs8Uo6+P4QlWc6KJrFb6UuZSBD3P7hdlZIZZ2gpFk1hFTiUTcJ7bs26
lQwt5s8Mjnt5aB0WSnaQHPncN18cg59U1O1/fnFbXRNAt2n0EiOYvwM8MBx2VBc2/wnw1l7ZNMXf
Az9LWsRJlo9V2vD5nmsj9ystN52X9pNKkMZerdyUKNjprmSWfSVEJxxTeG7irW1AUmoKPZVBoVlN
jL4/HLem0Y9GokBEtwXKBfb+2BHMqgQ/xJCA1alYAPdpHAw89DL7Q5VjEgb9cIW+uJJD2tCdpVZO
EDpsfHF3Qb/IwdYcRxWNS8VYAPu0Pov3Z7zQrq4g/4jPYvMd5xlaR61T9YJ/uzrjG9stR8t30f4h
q4r+b7voHjBRPRmoVa7/P0da7iaKqn7ApTqlYhepfr6jAlKgXu4hOwyEktwU+8+qEqRhnTNWbx+Z
wIWvxCZDnC/1ijXKOi0QVhUT3dyUC55jNIdH79D8ArA4thmRa+vSOhgCV22Kk9NkYXDOeBGc1FUK
txe5XOYUtJQvPjzksooTlokjcuK7BZXEAh5j9L5oC6BBSC6AWQI5kvw0P89dsVu4bRaHR92O9oEj
ShDcCLfrmlVcfqdodV8ve+ZHAJnxZ9COCYQTOBgVQW9KFNU4Udy4ZDcSDV1WDIIe2VuoZHG98Q6A
aJdOGsRFYt0qlk905UxgBmKYArl9w2WW2PTk6iihQW6U73cM8X3AZvph9oqwEWL46SlwcYVU+OeO
hmGV6+0ef1tyb6GeV0MGCNkJg8f30a5So5777ePX2aLNDyBLCSzAMmDbqbo/ZZaP6pfEWs2VkM+m
PnfMr4iUBEVQ/rKvdskdnQkO5uIQQ0qQSF5qY2amWBcPOUZK6tJ6KN8AOdpMilwqNjQjACdxC9zI
BjANWQfPkY4wfCjZCyyeNSPoCL99VDDpOLMCCZnb52a+FItNSEuQn4ZvrBfr1f2zrYGT4jLwyNjo
mMPvgVtLqIQxMcLoDncdLxq0hbOUpR2R7+3DKjyxrSwrulcLu+mDymgYxdSnY9WGIaXVYIJqeWGj
R63i/leOo4yXbc7BtUUtAjNDiNpdKgmFBLL/v+SfmSpwmbJ9U3e1ZH+zqZsttrbYVdyCr9T2u3YZ
rSmKfWCJDhtmvOqdUa3gxEfcMJUkSax8UVRaPnwa2O+5VcNpHIh9LD1+QxXBGq893fbHoVi4uxN8
q7Bz3KY2+w4Y+lFD+PWjOiWFpa/fUuZs9JZ+njn3B2FFZZ06yjb4LbpQFkNzz5JRBmLaaD6Cqqy/
Pe8QHBWJbOKXqrjJLV27fHNxELp571ioEIVv4lhjyQtiGtSEIbdZdBKVXqZXfwHhn/8iAH5my70N
Vjjl88E7uW/HFpWMh7EM7fMr2GrdRodV/XfAo2mpL/mMoJQVjWzRRM+XACdBLvP7xDh14d7pPEB3
4LxYwtS8ttXZz/EtBOPhf3yKFx2ngR5Cp1uX6H1wYwLE3FM/Le3uSJXzj/KgSJ8TYYKy+WdqCK/P
Lagqcw3i/ECDnSumBUy+91cz+ywnELocBG0+16fkvxvaboef7Kp0W9MVC0st9AVWXjtzVKNHvp8r
l1RlVL6cvPp5gC6jrKBQWkGOmnqU16uw3KoGPHGOeE/Gu2TPSd3OnUYnf2s6SC2pMiRjINC7g1Gd
NoeuB88hPDe0P9GLD/R8FAf6YwL4SefAQDEoJb1uxM7d6xaChQ5Qk9QKQxWn5Sr47Jpa4AaqGvBU
yziFjeergb7xE4+v6Uy0uOYb8t4ZGuxOn4vx+UFQcj525IVYKJ2x1Vlkm7YR6P+MOgPxqSla3LSu
AKhK/kU0QSR2wLul6EesX2g70c25ZL4P93zYj/1fqaok+dK0F6hHRp54ZumtTdnBjuyvFSXtZ0mb
WREQsgvVzv5Mo9Evf44EahG6p0KlaWsfy00Jwcpi3RgTlZC6MgKSlevQ/Lk9LB/IA2w7NFXdO1Cm
xQ/6C2B4DJzeoUId4V0Jg78EjXkKVf48BxdMrtI5Aa6kccPY2OCl92iANT1m0OD7OER9xKZK8xI+
CKTdPYGPF16PHqgDmLPh8/8yva07DgD8e4DRM48bpRGdLXjQ31+I8iZZ8GIPyVJtn+GklQfqNl6a
DGZKSS8HdJAF7hfq/1rIr9nmJhMYKA7QfhxIHMLvgtDrJYtE5jwN3f4WSAKRKz8we/Bsflpvc2L8
ubtJhPTWwsXA/0xN6GpdqN4zwYrN+M2nfTMxe0uSTzMQWkObaWjUsZcRJ2iVYJJFZeKOSsSS9HXd
Wp/WZ4ynMxV/rHQspk9I3f/904l2Js0WOQDrpLP6v7yfMDEzwbnvldWXZHcHz+vSfOVoZq4ksCn2
Hlx6A2UfpzYEslfdM23UCzKeFYItQcSYkg1tyymMD0FQaXNJazkGELiNzndh/Vqt/aO7eA6sNVFy
govz/tBu2YI+lgRaP/iR2i4LcVUFt0XXEldyTppDf+eQDV+8h4DNE/HNhM7PKwtxGZowPgVtzU5Y
/3C4Lj28hodOAKIdH1sMkqH2IWle5f+U8w19B+m1aGq1RNd1q56DIIcPsKwffop9oUuAKgckescr
tJoa7eKSxfhQkCqPbcZx3pgD5uO6vqP7tEX2oJSfuHGc2V6YQxGEJ0jSUQsvqiOsAwjgyfEIiGaj
hRjtxgbXGCxHBxx1I5uNSxNkcJNoUVs03xyzha53DGURFN8Z2Utv4gKNnGu6hkonV4j8+ftYDKQx
7Nlg9rv3WKB7+0ra193qRkXFgkAsVeIvGGKM0ia45PIzIU3QFffomHWpLNeyII+Hg2awnAiZNk/j
Ohj0ScIv4Wx57cTxomMah3s1hcAUn/OfJRXZcjcR8hGmXPyaRn5T8PY2/4TaGdU9tL20T72fBs7S
dd1czmAjAJsCaIciU+I2+K7M5VB0Me6MU7o75wKHdvLcIQbr/DVW7pxrWnpKptYil+Dgz1NqGWh6
2vKdI2M9guUmSQcGFUuUtiIwzZv/NFEQM2rwm4B/ip/EWGhEqy2dfTId3QDYZPsJ4Qs1eBRV6OXv
LOLb8HP4UrUCP0zMNVqaT61hDWozFC8u8LgQdZztqLN+WvdnibHfrlMeZELmwn209RjpSy/SZ8uf
9CwQ/lviNjRYnpk3vDR8M2PoORCZSHJW4LCdzPBlwFIY36UQO4Nja8dO6wQSAU+LQNTj+tzdA5KX
xvTB+pjICR5pLpAxd/AXfOar7n21P1lJ4LQK23mH18QLsc0zTyYJ5pjlNz6fNM/0s52U5Ff41cnh
v0Ayx56L9mDHq1vEeaPv2JYXr4BXKEvMxsdrJvY/FfG6rd1fcqWki//Ts8I5+H8fq3dkpWLpB1Cl
Z2ERVjvYVmfM4RSR9vIz5EtZyafa7pY7SmUUMA5hn+LZ7oHhkqo864DliAONt40nI7l+CD+qk5ZV
wv44NlhUougd5Q0yPbtp3EKlonKAGqE5F1cMrOS8IwFeuZ88chQBnOxApVp2bFiAQEQqZTL5qVm+
WCTHBDoVlwTLQFc35T67QYLOlxr7GWTZtanTWPC7OFBnpsZssmwRxUr7iHD5oSWkb2173Q/16aDc
NJ4ogSRwgH0MXUhzfqLegEK9NitHvhMNjv0+BH1EDYk1x7cwBTn6dH+CxqELfbZVA8z8acDXaDZ9
ficlQc40IbTgT5hKIQslkQP5im1Gtp5lMnRHbzhyhgkU4A9806QGAYL+F1S/q7pzsfsQVmeEG9LS
5iaeOb+ouBEWMrgRB71T1Pc37W9P7gcXx3rsRPAAFddeUEnzOaI48uzUOXUcPpU7fy7wUe7Kf+oU
RerYexDch/un2lPNI+1TLcN3PPiljhCY6GQtRDIqf81D82DIHwFmU3udiUU8um8dUZ7AxXRTuw1A
NfHwurRVpwK/I7HXC2ia+YUNy1D1a9jVPTNkf6uhbAaJl8uyCgm8jUs8yOO7oUyA2Ui5IZ8Zc9/X
l3iYqFfJA48mQThAE+Ue2CrGhezYrccpZ9mUUnwGKs6gWYsuqBnOkxxLbEXwwScJsx4FzHR7fGC3
j9lZt2UH9NpSmwgk0SPu7WToBsNfc4WGI6aGQXpcdTep/Kx5v17RDlBByauGvFdrfsnQ2kF/sXE/
lBGRTxaEIvluslmpJbDICF5wChZ3ATTlHdFB7LiADwmUb2eAp9wPvaMFn8jJglv7lV+H3zNpUBrU
RHCNcoNOKrS8ZKe6GydOeFyLTsw9kndBhBLy+dbfe7NsoUr6vgZwKBizbUSJYR48smN4z7i0IOw4
x9hj2B24pr2y2IKfidix6CLyC84/+Sxra+zBf2I9V90ySxG3+82aAcM0ebTQKbPhAGGMX5lKcgQH
GbFhHtp6bSeyRmSO0HEcjSu00tj+hMk3O+R6CKWcH2T/rj9jKW+fExX9mee2WaVUpAn7pcZFrYoY
yQo1ylecdmwU9GmXJIXUr8Qve+QLlARPJW1Y6nuz0jrG5RVQ+wBYX1nplqZzTsi3ePXR42p5NJ7q
PpVcmoc/Q/fJowAJ8cyAbG/LkrDidTpuzcZ5KDDmAZmFrYU3Xj8Qh75TpO4ReQeNp450Rcr8+930
OLtX3xcLSB4V12RYrq8i1jMVp9pFifx/JocEJO93r2kKKxZEy2VcTIZHdyIDkOFTTLssDjGfBcF/
32RfBmdVk2IKs0bMTgdIkI5oEU0pvlmDO5IXIja8UG9rR5sxrh038CalaMs8ZI5lgc1EEBPtih7s
dkBJVgQiFIrxEfR/UEoAvkIiAb2E1Bdvge1eIZOA1VbDKvuR/l/W/vXxwjxpa4e9a3hFyF0a0VgK
XK+Q0JOnAoBpAW7dqRBp/XSlUwJdkLJV8BXSTUp+RK8fY3u0t7EInFDowIRsdqU77w19KLn85wa2
M7OETA9j4eZnk/+qiy0pruDSbyDgSboeLmQyVNE8CGq3FrCuAgNW69zXPGvYA9PquRhPYHAqw0j5
g0Eh1F9Upzop8CYSCkwZ7HDYN9KfJP9TcRNXzn8NqX3w32GRopFegmCwhHFnQRQS5Rvw3fSCm2ed
7lG6GhvkN0jTaQQgHaZZJhL5ffYhWTVkPyKLg2Q4tue425LfF/PWiOzmU1n4UaY9OglxgA7Ud5KY
AiIeCIVCQgKEy5qmIliNp9e4izPnMbsSawuFD1igbZhYPArw+C7I2Wu8ptIdPg0gqTAhtc9nT9jQ
PTzZGJgLVBKh6MkzuW/nq/FDXfsbkghjY5b3NFAnDmMJekZUvixfdiCOB64aN2drGzKua7ZEPiOz
I1sAVawdmpaDGUO1QsnP/Go6KBlzjMJNEoMa7EdHg/H/Bx7L3iUkbaT/eJYihVcOo0Wprd5/Pz2A
4rqVKkId0BYGYhuamO0Y8TGNHdx05pesKXeNzTi+aRFh0cn56TRsqzLuVMAV6gXzGldtse6Ac4tI
C+xGn14yZaHgR9h/EMfbkn/A0iuhKdNhnOvO/VVmY5vObj9h3xAu0Oe3aV1iGLHAnRB8jNS65yd2
IHnEko1Eulp69wzoel0b+5Gddxj4zuOcvbN8520Nli2c8deIEiNaoNC5epbcMiEJtzI0MF+A4RGy
4Qk2ozIuol4LEuzDLgRVcc6/FvucuZzlexO3pxcmeJbkVs9AudnEkfZPMY1gGG0o+T3ytJRCTyhI
udlJrkko+Eyu4dRiM4nPJMMOaNODmhbx4/8InXhA8IjwQGfFuyWVYNtecfg4qQBFD+vzKn8oD+zL
4DyymdyzphcPVW7bcM+SJUhJXjcB6cWjFDjQECHt239rhnIwi/nSeiqdmmYd0wqjEBxPSMrpWPhv
d9smmbOKSKqcikue2b3vWLfM/CG69jMibfONa/5s4aWr0PwVkQ8VfGzQvcG0XKX1f0opPXNW2lL7
DkQAvekCFExgIESQVFI/nztw4BbqHJ8z6TI8jIVrFHMSN/UZ4cuBNZ0qU0LYro/LBSMj6f7ytxJ+
DfL+XRV7hM9Vnmh4pnuQT0P+cCXqHzriM4KwXVcvS0oAaalkkIAKbQUfuu7gV9vna4Y/nl5HtwpN
ZrxuVqZvosR9ImBqziymPMYgkM04Ty+DaSE/QOo5/R4TOOoPHLDa6V29hfzVofZSMI0P4ngfisb3
lRbkcUhxcCpxLb65Lqx9xazR7JmRyd1GG5QZhCsfQV19bVXnUfqTYyJ9R0LGCyJy2ogjg6xDH5pv
T/qLw7An/76nd4hspC15AlwM+MHVAQTl+XAjGgfHY1nEuNOnsaqVcBGilW+/M3worM8d5n3uF3Dk
um++2YG/rjJwarLoGRD0cI4NYf+Asev77Td76QSG/A4EbTKKD70ffcH5qmESgbJk/s3mYIQFhpVY
WneKQ4wyLfpuJ7eVWKn75se3MF6iPXHgPWzpiOA97YUnNNYAsTMA5Imlz9pwtUvaoA8fVKcL1Mk0
HObo8uj53A2OLHioSk2shy4n5myB9sXxp/kQP8g3e3fbPbz/iUwqOK/fdOZKIGTuCGdeGYNZUZMT
uR28cMO1tg4x1OuK74UcH5dvzD+MlZzJdDpqQBfeK6id3ahzj8avw48Xdl4ZuBGAXLBWfL/nJOGY
6+CqaXm5wO/TXJJJyNCm9CieSH7zOBMwuiLGPF1KTCCh4NLk+ZIFB4XxfuMwRBDXPYuMFwYT8rJ4
pDF9jN9mlm90JFDyWagI7fVH2pFdU3tmqoZpWyvkC9IwwZMkFnwUldJKpb2bqlrUnH33qlcG5sfG
XSn45yIxuQc+cUD80GJWNkbt5S9CSqm6E464JBFt1l1QA4EdkmBKz3V9e0sGEiEwFMukOATqxh9F
Z6SYmeM+1w3DJH8ws93tm3qY4xN4ROKAz+Kvvp+58I+cbmsSaxFo2Ne1aGo9OEG0Z3soCnfsd26d
2QoiVptJWlLgPwi370+5wrXzyoGMF9QiMkAUjsKbcpcSFsNAbyuCi4q0HX4XDYo5FLes+PDQ/G9e
OmnVGFUJEidVtvyQstDg6Xm6Q5ABLogVPvenzHLZVsqSKodsydUm2vJx62K37qJk+1Zo3c4LfCwo
MhyFsm1Kss62j/dLbKeusJq6TPA9ZnCgdqPs9i5oYOJljvmxucVDSiR962FaQNPo9LJkuOiJ7Z49
EakBMYYmLeKxU/IbKDwUuEezJQylm0yQEmCKqr+3Wiy15QyFNsuagwypp0BZAc3yPj4Ppi08Hd10
FRjfL8gdulZAbRE4ho/EYbn+AIYUkl2AEK9Q03dVqAGLqGsvPi5Vc68bYGOvxbmPzL8PvrOEXZoh
zSuIFCYw+lR6+9t2tUXJek5AOKhdQv9ciYmc+pRzJp38OijaoM08r7BB4g2usPvPwePvcBl6Ef20
YHachh9j/o0WPvcFMom/YitJoL12U8cd+CMNdPqomuHhFoGR4g5YBLCdaaVJj7eOseAOfLBaTsrl
799mEKP5ztJoZhnZlV3zk15/2N965KlHg8LZYlzX+ut19BMCV4GrMmPYzitN+uXP2DFy5MQ4dTJo
fbzTERHmqGzpsAnWCOnUfNg/i2NVnhoriEgIcfDSB3I/Qqfg/C6aY58rMnAVAnkuV629C+ovfyxQ
T7jAqbKmx/cvCf+PI6rhkOUG+HkMe4Md/T34fF2vLRPqA//DhoAe6HO3ZGmb4pYav7TbKbKK0BCF
gTXB1jdS/IORmpmry36WNcznlBOi9BJqKdbtMc19Z2cRuOTYIswe2QS/1uoWXYxGlWftAS9JPYuM
s832sWIIpNvSONJhHUOlP2z/4fg4TroQzJAY8zm/S7I3tNS2b/IZdnzas3Qr8SFLLzmUN1rESf/D
BgQjDrhJ1t4iT9i6O/UfOgTbK9jkVD7YdUAbgp5LqXoIX8gZJkmU5jvZw8fD5eW0vUnSyj+F4mj5
1jDo2SluKXZRordAem/UUj8Xypdbid3frE8gY3RNWEIeQtUHZWHpRzUGhvibBmoJJQb/E2H6rM+2
KsG8igoXCysp74T9MrUvuPgvWyfhnk5tXCzB40RerawqEQh+56XNtCM1awizhzledMU+CZDbXDkT
MI2sZ2Y8aBO+WhQlETHlf1SHIg6YgBqML2BTjrqnNrtDWqPrb1SRZmaITGQvyk+ieZSp7EL/yvNk
LSMKGzaJBdlP2cqyq/NFuuHhttqZu9upm803A5sSfb1kKMatBle9upYNibzFpl8qE4Y1spgDh0iX
YjdI3BD0L0gwEDad5p8FP2ckgzlK5fB8UQ5MGuvibm/ypTwzAPgfDNCHBX11xI30ZBI+7es8J/SD
F7aQ4ldrdXyHSALhsubJrz+jQsr57m/ITzkh3EaEaBhFWN3TVsoYm5gWzVlM4s8qMnIV8A91l5eW
Oty/sW2NENiBqGlaeekoUaZ7uyBAIYm7kCAIq5N9hIG+0uHrxLOhhbFwt1TakAummNHQttmR1XV5
odRk5ZuQSyEOldh7sNJZn/KHKvAJX4GLEkxijWMh2DSZYCawaFuxzXOqIcmGRS1WqKRjcrsfpOI9
m1K/aUrWqI7h/ynWGb5zmAr02B4Rs0vAmWtT7A+b7lzmgipLDfxt63XptgoUGaQgTxRvIDzfSgiz
EL88+eFv6g2G0QoOnSDZy3EWD8K0y+is8364eamgN6bdTKVPJDMEqGFvDIlyxtHnYBoLBpadDm8D
WoJUEvh4MHSFDDwfIiBzmtQfG9K8mdxKBvXI5hDc/eFrnRY7UJwM7I3884dwbI873Ax0V29eJBst
wdOrzo5LXhmvvb46mKXVKum/snNQkyxrpRjCfDNX2mx2PPNBTFFW/XQi1ny92zDiSuuSI1LaKHwl
GS9olmY+goNhEnqte3tTLQgA9AMjmleHYP5hkHyLx11YwVFSy8nGHFiQ54ITyrgSlnQQKw+/ibx+
fVRlrjIFNThRM5q5eFb5jPXXfILYmgs7UmQIJ/DIvyY7bVQTqsf09k87ja9lGdiGhcoNW7KX6zE9
ExgBoKpUXdbRNQ5DTRjk1FuIBAAuEnrsWx2DTqTdj1koTVWpByZwy7wP92GRDS+F48SkKfX1VHnS
AWq0nC0zi3UO0L/TvuAH3IK6BJXSFeR/0DskJybb8mIFVqFLSjounMrMLESR9voj3yKMUkUmRoP4
4Utb0P7YBExzpQ9glDIHtKmIja+2j0k3ZimBEEBjzSRGeIUylP2rM/lG9mq/Bxc11K3gXgBpxnMK
VxZMn0rvGi7tOCMh5GTZEJFk6MjHXKYXeusseCGdyjpt5sfOzytrAtTj0Wy8kfZibkXQ22qdpCh0
iNoy13ZEhrzVIokmfCYAexHB4pJUOii7hGj/NLnod9Ghy/U0WARWan/KLuxTFc9ol9Kwo8Umipo1
l8FE+usrwQS+/aB6bq9hCk0C7iJS2kXocbASn9o+/tkWcjmmTLEjeUcHMbjWvCbm70iMatX2yFlC
+k4wY1wodHwr8aTcdtZjG2FmeFAw3T2g/XccJClKDFIYZbI9T/0MgcFw0/N4kOfgfTOmYnzlP/HN
DSmGyFmrtZytLXHw8xQjWMi6aNy7ly6sAnPSQ8oSqv0FsXLJdY+gzLwsQ8z3PgR6RFaO4zQKLwgA
yY2O7rKstheBVpnm9RiUSoAYdcvuY91QQXij8zpGKECapRq4fysm/UEAYZKlN6JsmVTQqXy7lczf
4+SFIo5LQyFfcdm+ycQhCbh5AmfatBUyef4QSFfdwZLH5uugE3ujuSTYSpA4M7Qc7rlcjI9pMrgL
KFiNa3z4jjyHfMaoREzxkCB0yxStNsbQV0TCAFxLY3tHpGP8aZr2Q5xFWhGOBgW00F8zb3kg4Ti7
X26sPzTZ7eKusQQ88yb4Vo2S+3dfUy1cne2GTwH78ing0B3qxqbf1GroObSjY6wAMpdg8zjt/6GB
Qktdv/ZvWzP0b3B97odmLiP5JrI2r8dlQBD7SCErDeIWBwQrs4tLWyIILexdxbsr++pNVS2gg/1E
Z4ZQfVIxPSp7h+FQECgKCgCwVLwLd5iw7BRG0SSnLlom99CQ12xpkXNHRt3pa39zefJIrUuiTSBf
DRkNRQd3gFbpPw+xwQ4wi6osko8qP61l6/AYIK+06QcOSNCYrFNDUjZGgvxePCWq6FjdhHeVO/7m
VjJ8gGDswy32RMIBZzlP6MHlqx9x7pzrIfw5WwI0Hg1GNp1Ilhd3MT7Nw/J4xVbvHmbKW2b/zKSv
UjO52E+vUhWGTkHi0iWhfr8YvEkEjrg8Do5AR5rPfuS89+SEaDLt7cX9f7GHYWgFeLvXAc7olkgl
R6a8/2YsgrzSMDkEYx/oprRrV1/Q9PRIdqCD/TSZhEYALXc1/m5Vx4QOytZSbMRIGcyjBcdr++5L
mdD58fv0l9AN+CZF2sPZlf6PIn9y5ZBKcj/Fb3ZXezJvsq8F3jtG9Ohbl1k1DuckVsTInbnDAtp2
wJlUOb/mQlAk5zSUKDjDznLO/UlHc7EwxmBVikt4wTVyjqARkDcqWOwoEP3fDUiAeAgwd8lrSP0R
rU14OEH+UMHFnp/85c+ElQ8tCKJ8P3oA1yg/6xy/EHivaeO1wEV/GLEgxRNwP3Qyo7CiGKVQn8VC
nWk2WfEuNvMNhAqIfnIzTseeMq0H5BTJ8z8XVqmCg8WG3WqrSsauhyfWc9PZP+nMIh5kR8oZAkDR
//5NAQl7xPAw3Q7GoDtIDEh5JeqsYzPFkuJfrcEOVE687+sQ7/Fxxv6PDGgKnAhKGQJenwlncT8z
132zcYcmVXiR0s6KUWt6Pz1Nfx73xMogp3nKg8smgvwF2tTEs04bvnYZBASUGGG76y2nT1c4n+V3
tN3CNnt4JgN/8XrF8kbl8wT9TZWz8gyCIRYio3wBiiVJpAXI3Y9arFvSZCEK5nrlvV7lE0eIJLti
/efa/hPNl/Bc4Z96IPkVop1+PVquberSDZZX5fvIwGl59b823PzFncwrJp3r/mW4qYzEplJ18X0H
XWzV+AEL8pgvlarw5YU9p6r9iocO7w97OAgUcAqJd7ya9iC9FyS8UdyeZrvi7sfnBkjs0/V37Euc
NciIFU0l4GluOeP4rUYuCnad7h/bWJWM0qMHAeSOvpRv2WAhoErkXWx7Qo/6VIXfMw+XbwMFJW8Z
biGiPvaA+V3IABx8SpByXqLOSuM7BO3XPFJFCZSyoIDfZuxZ2zfMn+p+K//jVTMkgXx7VI0uyyXr
jWsR5fNkDBqSsAendGbEXiUjpFYJRdPKn3LhnxSDQVBkhlHlAwtxwo16IQc0csD4anLZK6KWBHOs
xbgpgUzVC85PCQR2+gav4dJdr2a2q9+BlrsJVmhu31q+zC2E1bZq0Ao7lsbvjC+uaDyqPyCK05EN
ZuaWJu6mf7QeancikxCOQqSugygYOV6bHGfECCaoqWOMjMEPaMi+z/cWwSaZIAJ/ssCEeAOEUGJ5
SZRSjla8FRcxB1NoVBvD7jH9LoBs/c6krdsU0ad8SAuaWhI1sTMLngLEQGPcUEDNSCuiIqFU8xkJ
+vJw45V5hmy4M95xuxXYkJ87aBRuU2jgLLZIRwwFP5H+PBitHlW0MCI8e1vdSHSH0AR3RUX25ST9
335F0EjZJHvbbTAyJSvpXIbNWEI64wYvBY+vAF3JOmJId3XR8o0ERLO9Dh5ZA47cVm6jCcmv7BFQ
SnWXnuotfsk6SDytAsK48VUMuTQ379lVJQ3R3rbj26J/O+MzrcdQ5kEGLP8DZ9HqzY/2tDTOjJYC
EsJ5p2Agjht9oMj1Nb2tAp+RmrMDmfUliXSvh4UQAf6FgLbvAe0t7ISxLTbjft+rIPDp2U8ZzOr9
bs0gG02+KyIBeRxQlLj1t7QqDqGC3M6EYz7v/Y92NC3J1ZI7ejTmXThbufa3maoD8GyMqMEyOVxh
cOYeZf2bxRycqnxXASVjAqbzM+OOLW+EgUSRRBW1na/2t8wDn5VfMZJ3e95wspu5bf3RwC9l/mt6
HnXMIlNuvoZYV8lwkVZap2/kfFAsh4tOBlw29tycsylYFweu8PPPfWwZMM64DMNrAGCbwP3AmSx6
hlExB5+pjHTTlnQHtSOP/Z5/zKKR+8uHyEc01Gn/4Mfov8e+gqVOjoGeDtD3/zMhi8GdQmfVx+xI
sdS7SlV5dx3jIRf6AGP/lMnk6Fa5Zk0hxuEk/iWyhxzqjxk8+MgNUt6VtO5BLP6VJjJ6gEXG0NC1
D+JojBxKZyJRC0FEmEH5LijO7wsAKeTfkSd2TZqmPgtJpeRZlGa+lxXnbM3RF4f1y5qjsnhEe2+I
u5R9+bPMqV/djBQ9PXgkHXM/+47hlOUlRoyzxfkVHLEVKOSICJk+AByUqQ32kAAIriCf+zWRb98D
gy/+LE3OnO2jsX4XC1Q4jfP7i4ELGHzAtHoo7sGScqwABA+EAVZxvxa0HW5z5xDJur8lfuXyR8Zs
7XdrUcS/AsbCmHlQ8VVl1pf3o6wI0D8WM8akMwQDGa51xBoHPsDKIe0RSNPjzutHuYvGWPALUwtc
28pYGPPWvzH+7vkWEymhnbgerZfY/lBdZ+/wDhA0PcA8vTMuXXeJBd96VzRa981up4zWNRkW3poO
r/kfKzp8bZfILhVKAhUojH9YHtCo3zjqjeHMl97ulp7Dn/d32MybjHHphhWiOmFI0zXF3zQziU/7
5inaA3oqy0TlB9cFIz9/PzrBlRaT3oXm2Db4UrPxIIAIDc+D94QF6ilpQphQVUqyX/I8fjf98Wcp
DCmuMJl58D3ZxH/W3W9HIwDUBWVp8LXa05cLHU02td7rp32bZh18IKk3ebuKyUEzyA9hzRfudCcG
0rkiCn22gUFCJnxGT6V2u5IcG+c/Zb9SQevpJ0FV0Q8PuJ3MR2cgp/XyHBuV2YXN3zFGIchpGpem
VXEwFmf4rhgqvsMwSr2RLgoEBVf852tBZhG7ENO2ukdqAKiXN2d6WhZxhCtXD/dff+xi7zmPjTVv
mbcf6Ej+ChNsy0KcantLJEk1DUnShHYV/ubzXJJaMZD1yD2vniZbS4H1b62MOezjSmQoDUnSguVn
F4HBdae3/2hnZllICFKzu0IpeimKHaKpw8SCd7TOlV0zfEl2wXWavsskeh/cJLvi8HYcyHiUzPro
OVs5XnXJeeOFvzM2R2ahaZo0hQpiV4VYz9YZb515cmAYwl9UMnUQRR2RmaOkTNvu1BIrozGa4tEA
JqqfTvmiiXvrWGz2pMO94fYkg0LVZJa1b9jX30oGqOFGkWI9c0stYg2Dgdrka1yF9XFW83X/yGOh
d4E+ZyRDqEX5TKm7TiZL/GnDiB5o2ih2kVPabwFjj0H3P7UYMzSks6SLYJZ8zKFDfzrwLYOnov0C
dLVHKwYfYsEschCISSYA9kZRAw46rHZB7SNHHeuPXZcpXw3SqHPKkFmV2wzSeCFPYWTYJ3Icerto
e08PmXMCD/HMq5rNcg9VUpTvfDNUTrldbis68V9Uiz8VBAFkSWD/ZcFIixw2sZlHP+6Yvb7ql3WU
PZwQxS9Gr+KDFFuKz0mFvAhGyarzZA4fyOkyjd+cvKUvvhfQ7jnhdnlSVy8zGxtZaDXTK8Ivvmi3
PO9pvl/k9jlogP6HwPAFzKsZJjGwKDfAnt5a0WknUZCflh1ofArK1/3czBnAv0zyXKyAGOuj3Tf0
IR1VrpdNA0mCEmwMuqbxdrtCvGHNh7EYYMT6ZZXbuoN3GaQhiuhhITYCtR9MkilXauQnakwX9Lrm
fdlDjVzaeliCL+30oEhftjL5JZpTYR7X7d0YRWmmSw+4Xrx/hVeU7r1zXEWVcEnGVW+imcktrmij
d20+oVxylihcdR8Ldo06ZGtqDbPe9hwOdM9tvyW0ZuWyaP/qKZu4+7Qgd+NiQU0J39aayTm7bF6s
iS02MB3cYl+QqIz723yhMVhnf5VLTC95UQlljuX62VStcDEbE4vMeZoQSl2DXgBaWk9/XFFHKhwI
AgDGawsZfl4KJkKUoY0IGY35XXgkrHbrKzKqiUun4zCfK2fO2fLTZPlbuL+0z3ZcR6/hUTCbMu97
UNhMFY0h+IA99ee5m82/Ng2ok7cjqd3YomBy89tXbg8QXHYm20cFNtlph4qAC9lDFcTANDHw9s4L
7QsMNsJQPNTjqJdoTJ2MLrFoZb8YZyaCF1Vio2YVME6nsIjv3UDKstnSn21Bf569Xu0OK7pjZExw
iGdPzprQX/DSORzZ6IqTCIaGfCwDgm+swkz64Ya9R1SY7916Yu9RmTWBJRPfWfvcymGkqMCdr3bO
jNaA5HZEv/IkSm1VO85fHFcociVExVlsNSrmuuJu4Oh14gdPWdrBoiulCcQ/lCjPRQ9IpjUORfst
qD+xyTJAg7NWzvL7dZppy0ez+HNg+QZXMrOljnbXdxIRTt6Z4HVdg4hY7Gr0HmOWFQGY/ZBcAYpa
X4wCVto5PXzK3xdONpFBtnmIv/tkiE+aTvldlVndCktgGIE1PvkY+Ilfh8mBccwwAzEAGKKEF9RS
pq1XAZx160mfa4AwUGo7aJEUz/zRcM/Dk+vhDr3W0zlSrTPpzQajDN504qso0XjQ6X71DiiW6BF8
F9DU19Z+/H3YNPQtV/gCyM/AlGaJsgJHccrZhfbnv+ssm2Q7gbRYkFE81iZoVeUHE12oure8O6Wh
AStFGLDMGacWSth/nQ29usasx+a4Zok0cIgVFTnfeVvWw8Pr2Si0cNis7ucfuQBwQdEx9vsaERxs
sWLuj9N/LrVzI70cF6LC59KOSeV3TE1O+zN9beDcpk1Rwou06u8mp62glu4UxRbbSHJyLVelzbt3
jD7U1Zczs4gbIffHfKgHNrrJ1wcXlcl2sqXNGAnBGQ1kVZSl1LPkmnE4OBJu4Dzn3i2FyMwMM4vn
kmbma45ulahruS46/LYrLhBG5OO03T8sUtynksy9SfbPxQ8UdmSG9byz/cq1olYE6m9TiIWC8ySx
oa/4ZoTfBP2i4UAACBlP/GK6bl6Kunt40DSt8XeO7T8lCkpms1Tm/KHVy/kMok6KSHIBSoE+WDXf
HZEv8/l+cgN6MOddtKFfEV1Czdt4qPv0bNIk40F4IYh4LTTg7mTND8beOUYbW1CqdpRMPd52zSkg
sbGRaz2+7ad1UvmvFWHKoitpdNrT4XGyG5MHa+t6TXHJoB8BNwDIAkWHSWkD9MXAHjBC3mUWPgKT
VhzjeDS4Vbyd19HzsyTY/ygHfNDMULMdlEK+QFAkq9W9HWTH59YilDDEcyRJVhibOI+mvPSbP12B
L/W27CF8W7k5X/noV8mcH6JUtLj2X+ZJF74seecJkCH0MU2N1AIRhnYMmyPKGmfFbFFzj+8ywjzh
rK0QxGFxhSoAQP/Lo5gRIUylYfA5hyBCbxtQpWOnElfw6s/QEOOwDDlRheIxv2QLyktsOU/z9hGu
ePdniIk28qlF92o1lDMRecugsaYvZt1Z44aStIG7w7D83rM0A9dZx5dacmtELQnMaqi/Iv6vLayx
7AkzBsKt/it5TLiTxGe6QyEkqhQZTKp5ybTAeNnLGsNF0CImHr9EziTuRlFsT8cr7c63E5Tv6xN6
XSvo3ngTxN431Gl1bJ4rfWUY7sK8fJqHY2PWStoCC6WBpd+mmu/eA5r3I0W23GqAgaR058qNwcIC
zB9Rz1MsDD1NZHPTnX6VJdEJJnl2Quyn4LC4U+rM526VbzrDAss0jGmBdB6wBnaMN38zjnvdVYsS
T1ejwjeeAcBL2asOWDNL9nZsJHuR5ZWeg/H3whpbzI2nEz+Ddf3dsBOX4u2F8BJuwyR3xGj2tie4
7MH2DApPfccEdQQdb6fCEC4XVuMW8W3a+EeBQmpNwN9ygNT6TVJmKSXcwekV8WQCkqaz4qAiZG2p
IHGgMiYCV2vC88VY0eDyUFoAR4AzfvtTD6E7jUHAZBX6gUkxnl1srfB+mDU86eAgEX1Q1S3GRbHq
2Ycpc0vnTabw2uNW7vmnaoEqk38VhTxOjv15KD0VFdT6nIRA067mwl5+MXhX1JfdOkPT00uaWd57
oufxXKxSAycCRA8g4Bbz8th2ZJ9oP2NI+8NHoo+7/ideVQugVzNxfOBlp3x5xXC2BJF7uktIadcO
M+USfzHGrUk6bPTdo5D8CPxJRUxk7d3NfsIAy5Uzi5myhOc5Tz+j5ab0N85Sr4VJbzEv4X27vcaJ
KRadNre3LHIm1N3HyqkwsxvfDd1QW+a7gR2KwBqAoMbV23AYwPHSHwZVX+DvKPEuTmphjgMgIDn1
AsJtMQCskvcco/0Mxa6NikbQ77qlW9l7knRKU4OPAjntb0zRqBLXnt6cLW0fXIWELBYezOQs86W0
kPxMlLdCk1SwARz2fcu5jR7ULIE5gNWjq8RNjeq2+O6ZesuhO8evYWD+R9zWirJHCsN3MOY+LD26
h7T/6RHSmzifA/xvpsQvSLm5T1rKTFz0zDTjdxSD67sFXFe4lwYLRwFENtDME7jy7W1KAoqfUzdS
YsN0cglckoG7zpXeht/wPCG9uVjTL5JmV1cr4tCiX1CO3cRWuego2jxuafXIPliPL923PDO0Rcch
LE/scMzohVY1u72dTX1QP/kRdDhFXtNU6s12r2nB49837W9ovUGwSEHodn/Qg+YSR2JHdHF9aQ+G
tQXfHQ6cMSEQIl8hskJsyt10etPw7d5V1IRnG0Z/PLp5DbBqGIJRN5QNKDa4qFxOYBgsYwvf3GK2
BP7iscuwLXJV4kQ/SZMWVYhm2Q0WlPjvOQKLd0ZGh3XjlbhXsQzyVFFRnTYfL4OVn0uhw+rieYRg
4kM4l2jUVusSpNrJid3pmHnUbb1xFFSMIBLx5aXz3/UV2Vy6Qyrg9jkBUzydOB9NzoJe70P+irAh
HAVJuU2cTWqFH+W5BsavadxTYtQrKMzuvQBol2mjVxWs48Dd4XC71JG/k1jhkDKHREmBIWLQYSP1
p2pMNjF1ki3+7nS+eD8P3MHgJvOU9aoMZz6bGQ3KOGMm55/TCgXjrR7V+8NE2MQFPGXOVwkqillT
+t/KhOsyAJeNAGw5F12em+ZWh0k0TD6v6AK2zok9aiMx+0KeR9mIk0JHR0OLgCrI7DWQS6QdJEGJ
2Pd8RBUO/OOEHwWWhvzlh0G+LV4I+fXwvOi0Exs2nlZ6y32XXvssliDNxThabjGHv/d7FAaPchix
dfJbEsphvFp4Smc9TEUK0dQGgAdXp4gkjVGfNEOKegABv9BjJKn5Z3wjuTz1WjPXrHoY+D6hHPro
nHwvFj78t8FJHE2Tiqmx5u4Cwqy70cy/h5JHprJrnYfX8X3MSO7v5j5vlofEKWREDcUz9kTME0Q3
PNDu7JjxMKOhmmIFO0OaySSccjfN9mqLuKMy2TONInQsCrXUEavDYo+tSEHVKTLF9Mi7C2NU/rBV
xnLBDBMvXQ9d7UeoXlvbvJYK+E1II7hhec7juZ/8SxR3GEB6Mntt+c8FH82nqq02LkLJ/bPL1NEQ
C2U1pMAOnoUYw671QgsjzzIyKLZIOuhV95wWIwet/pDuznW9BB44dVKz7yfi0Sa1jcRHkUF2KE8b
ffy8BjwCSgpRxwUzKTB36l80+A1zhqIrUvcmstUxcNeFcqnGjYogOTiBKHzlX/ylKR4v2drrOZBJ
uMNh7Af9N9l1MgG9XS46ZUrvNmAO1Ykq4n76UVO2ZG6ZvF3NAaqBMFnmtEG21vIuY69fojEQw+kc
uuRwlNJzIBobWl43UdIeDfm7GedR5c6Y6viINtDn+fFdfqYAE7j/9y0cbFr3VBdWJ4eaGGqx/NJW
nOv+ZTbibu8SZDogcjN369uiEAgapxieKkrXX7eON2q9hrBub9TucT/3L2TWmlZRcptR4uzNxTv3
d43ku6jp+k3rfPuuq0p5FY0lLlrOr+qVSxtNrj/PK0U2yhaYrl2HZGx47RwcHaiid2np6/+3TwXn
2etfeCHN4EsMsXKWxb+DzeXytwp0Bb4pyOW8nPoznX+db3I1u/WSG5+RR2HPFtUvazaRVt0ncfn0
MY17+wx5zbauqqcpmIbLpmztm2LQxRFwOX8PGfw1IPl6OUsi44jsYrU2n5Qdk3fHWXSZ7F/GPBBO
lr0cn3TrOccGmTq5unssara+PmHpe+LzxmuEtkx05dHSo3bQQH2tUo6Q/EDKlXOFmqpqqH3BQaf5
hVOUqSTK2tAH7894EV91ZP2Wu85BIcH6vt9uo1HSM7PetTGbM7TdswcAQd6NHQbKpvq2hbvzLo35
Qhas2NWhV2i0Sk5hbUTeiTxVST4eGXrNny7rqrHb92um5bDWC+EiwWtPj60JYAJakCzWJ6i3aJrI
c2j9NQJIfY07ujMqO0KoHpoA+VmlDT7FkUMpletXxSNpbHMT4Tg9YcvEUhBmpZpWgshWweB7BWr3
90aTMrFW0q7OQ1xvdFyaVEOraFI627gYkMdrZLmK/1BWM/lujYRaI8xip2gtny2m58GySbMBIFzN
YZdkngd2bcGWObliCFLn9Ch0owpI9Cv1RASzrlLzy7jQJ8BO13OW2jGQQiEjVMOPIIOpp+NS90+b
x/8gB0BzFAFRJy/wgMHJ44Q6yREBrr66nhum5WL0YTdNVjTmlDwY+e3+KbW0aJ0tUBgKdIWRFSlx
V/NjIshjJ2XwuB9YS/mdksgI0wOlW5yDSv3+rSBT+9l5XZ/ywUdyTnyQikaFrYP2t91nEruKaIYX
7OOcIzeNLmMYKXVXkduvLVwEuONLactda//yI8jnWiyd75zJvGJieAiO1vigFOUUwAN3fLH///aJ
NkXBQ6cWc9RK5ToxOe4JOxOoNsgz5b+EVgN0R2tdzRQbUD+wI1nW7dqVfmrOE42XMBmUSsAi2HcU
r3VFEudEp3hy4CdjPA6paRK2SiYSeUTLUxZW3a5Vz/PPyHcvrnfONyUyipu4eh+y/baPxcZ7oka/
pg7fcGGsy0Ufxq9LCUI/4rW7/tKatdzb7/B0v+jIK6+1wE493wyb86cnNv9EE0bndLYgGb32k5L0
L8v6fgKOZkHhRxe6lVezKOBpxecBR80rtV7p6OwpxXom0thS5ZiLbUtUSLThG2MOHDEi1RRiz2kf
ymt7M33JSzD7uypB4Hdo76h7kU9DTYJ+bb7hUenbLcaHJj8J/CmhWTY6qdPs3uc3yD3Q1XJub1iE
czyKSxpjdr3ThRksyjQuxv+zGVQ/lQi/9ODMi5AHIfRm7hnrLqXxid2lDdL8yfFoBqokXyjSAjfg
njb39Vq7UGnYFQuS7T0Gq5eDFIKd5/gx3rausbZnTX70IPAlmTo+ociZ22gwEMO3kEI1TUAOivwl
/51QoEG7QfmMBKriBMn6cqae2ZYJWdLgSKzMW9OBM9DdUB6VCNKrnQHtLKY0uJxN05BjRP98RDSJ
uyBnnSzOF5oaUHDsf/fa+XJ9+WPS1U2mAgYzDeKijS5pLI6aMmy3gjWGqkYEFamsQ+0KIZeRh2Tb
9cLH/SDkb8CgzAkkzPAFFK8kQv5do8XpB+TJRuVIj11+tUyXyCZuQy4uBIK9v101HcRqDj+D2AUw
c7xCQj49omQ0Q8QiszoUldvLZqG4srFgWWyjxIBvU3I1bU3PytJgfxaQ91eE0tVErabDuZI9yqNY
1s403h8WEhYkR+J6ljbWrBITOWN7A8VReN0OVbfy97p8GImdH8KAxTDENa16Ncgkg/tjzExn+sSk
VsWB+iaUui1wfdxB1QPC4WJ8AjIkjQBgx+RlLuGX3YfUa+3Gqr5IT4fKFe6bsT/pMsC+bP8b3bIw
eK3nvZPSuqx4LuaQoaeu7lTNZwWuqb8zyMIesCUxkcjcMExB/2BVrijVnGz/frMALJ6jLQj6GZCs
XUbzgNBYBXdcmAENA9j6BvdXdnURZkrfwql4KxUg0o0+nmem8rfSTTAq6XPdM2/JZHuLC1Ivb1qp
V2ePYoV5zNGfv4MM3vb6R2aYI/JgBl7BXXtqGqj+pvGqE+feS0qKOwmiLF6vGgDjWCenOy9U+LWc
6EF7hugIQKJSkRcF3ItriePdgMDFUqDi1cbAWfZVFyTs4GrKRLI0wm6AYPgY1Pw3PTTC/FFt7LgY
75Uko8cJVz52VcaquaOvOF9mlXONeWXKEF/twWCM/rFGmILYzwAKQLYDC7iJZ6xIdeelfl7/tIOP
fXjJ5k8yu+BKn0GJ+DFE60/CGKS/Dxa7afSEcUvJhzqAs1Zv/pq3kt1jgg7z++qkmlG4thUO9ZtM
GfRLyxqBUMdAddDh0xxxKOocFhGlW4z0NT7FvxoE74jWxYw78i8kJqehy+gS8QIAy8YdwMtPLBiD
IP/Fs4K5Dfz2+qjOD0hBXLgJTniGitXlXP8ZXFuHr2BCNsYGtcTm2qTtqXmOUa0+W1pTRSnqEjge
5Gk8Fs/anVtJcv552TvBjeztseMDzNGLORLyDmqG/PfrLkivU4R1I+C0eQpl8zDuKZb9lCtQJk8j
DD3NmW8iw+f2h9/njSlT6fuV1XgLbUGYkooYuho70IQUgBHXfORznSlS93QX2CAkR0uTjjD56Mas
MPc+ZlEQ2X/D45rJ/5vX1Xm8T6fMI/2NtIZ0RXJeIOhWYs+ECbStkvobwBiAkPJcaywVHvuTkhpA
71nfNrJnPUNJfRPjIsWFDaI5B90ukXJ5Hr515yn4+QKLCtDW0mmaStdTgxMKEwTWdWpeq4UFbeVv
izQLclMRX3vuFcObqflHq0QfW21tMmm8MbR9acNgdRf/LM3XIBnC+YanSBXRvFrCGanmpjgENchW
mbAK7ydiAk8/5l1ezBqk04s30U8zhkFnbt68lgEXXRVXV8GNOYlZUOkOAOmpBwYPbfH+29v7nrzZ
Lwtidz1gWU4tM219dpLyV8fUCO0Sul2kjhMMFkCeBCcUkF5Zki9r2gnGWUDHACNMLgJA+bYTbcB/
ULMm+TkynA7ediKM7qa0e05+O6oXgY2KnZfMeNBHusVlTlxuZXYPfgIUWh0o65VSwuzr8pEJOhX8
Id3XDfpL9BB7ThjjEk+7OAj6lHJjhH+m96wQcdcaqYd9LFpbHRy4RVc/LzWaVMwG4SiATOflikGJ
h5EYXgqOr+pRPe2u784Hy0pWp94YkR6e0JXASl+2rES9OWafy1yfPHyAbYKrCf893msk5eqGPFen
7ZyV2LFOEAQsCmGS4JJRH2duJgam8N1Z7S+Wm1mu4SVughuL4cv1fqeuWkJ+wKjIKPHo+SeBOpMX
fJpXNGkU7SVcZTCrKNKF9k6jxH471uOnxufaif1kKS3q1kJ8OcqXBIaRm320B3Iy/H+KesrHk+Wi
ivJb0GkhRIyPi1cHAr+4XRQXEEeeOlnYShHUjMezRatqB7z/E8eRKfE8Vb+6F62CUqjdQp9F5Odg
1tJDeloQf1BhNVxjGIpxt3OUA8qQUQqDvHsSstA7QoRr5JL0XC2SIJi9leUvo0ZGBG/XceqOhG4z
VrO109szXo/XIRTecFV2k2StwqHTOaCdy4+WAIQd9VUF/gshX1hsMGUOQ9Ip9oH/VGD0Suic0QL1
UzPxW0dgPa/LgivjHsd1dibfPockMhOBQsosjWC8SvmPdhe1zpdfhI33tCk96/jboPMu/Sp83o15
bvwop0wrX/6+IZ3Wgd89NWsXFNb82zeDajLDpCQwSiDztVNlOX2USKU1N3cIUK4gEig7os6ao/56
r6ny11Uw9G6FX1dnIMe4atQevJ9N7R8iIBOWNUtK25UGA4bp5fBDG+w155ePEtaYef+U9btlF01+
pqk/EgNdH4yT7avs+FCyD2PmK8qmfZx6LyjyXxv+jDe9WdY8Y5lqQZOUXjgFG4K+tGMwwls3Z5JX
X2O/K6+Qgf3i5HcEesfJEsFJpgV+tdei8q2D9VpiVjRYlI6XVmngYRAM8og+flCCErn7Pn+/93sU
Q/DxHoRGAwsTqIyfzkrwJHhkGnzIXkpPg7NCDziuRuFkHbybM/RjCN1wHScK3j03nBFvOAyzcIf8
jK+CN4d753ciC1jtXcCG/c5Gxk+U5JCBFU5mvbpG+UnRRfASi99ELHjA0QQz5gOoimm0mdZOr61F
HJd3bGbEbYUGuU26S7wIVQ0xvtU5FCRzQB+CNqQs89pTDkTK4t8NTnJ7KOIzC4OUA7Tjw7iiNxU4
V4GPTw4A8EMOURUchk6lLxXRI2Q9Aytv4VoUTuQ09PPpsQGuHuRdL1iP9g6FCrrt9LCse0CpCKAj
NMFAZoa3u/rDwzjc1smH3PR3P+T1yYjUjstrAGHUYx+yRmiW90++YvjLK5WCa5r4ptNdSIFTGSw9
u2ase4fFlkbEbhCJGh1SRSvTtletp9m3ShgAmR4GLvsn1Ya/A/cEcxpz5SuAxeb6yNb6ZTNeGKWg
4/fkNMPKZAUUiiQAfdJilGQ2Xp5hFHgc2TLSR7jIi6YgM+noV7h8x5AFAmj20l1ebyAc/N+pWGHf
o60fmMTg4CqczpPu9qgWVZ8xcfM77Au14RFpkU9mHD//DoFC43HYoqESPNVGxHzbO6AUhXljAL/B
6LEKk5PzxuffmoIgwiQBUqxwBLhoEqTeHNyG6mmrK0p9TveIb6NTF/W5bzReAeTQ1rB7KpxVzHPN
r1zY0akSVVp0Wrrza8FtNPGVT8OJd/W+q8rdLASxMCmhkm9iDk2nbdclR4oU0ilr1FRXu9U+SqQ2
s+Zt7GngJUXA1hC0beHxAVZHH3D6N0LyaCKlrg5zwWtuvjOzGc4DNjFCtLsTK7biQsS3yKmf3FWO
tNAjwx5bdADiA6OXlmRAFWOIHceoPaSamHb3/sjCPms98p1aqpRqZqiLBo6ZQDOS9FWS0luH1VqX
1HeDBPDkhGzGyrdEThHmL6Foxdz6G/GdMoMKgzkZipxuF6oiAFKCq5NZ+YCGCC1iieG+jnG46G9W
VAQAsIhf08Apo4pEUDOPsiiLfAkTk5IvUlBZdRvztEp5Qgn1FwQFwxwK7jkzoy+CfVjqHJztc2Gg
NxlJJxI6+QWc3MGbSTCvHfn7iBp8qcpufx86oYMfLzlTaxELx7lOZg8ekZABaC4wClLUukHj8izT
6PCQ4Lb+bm5fyHEVdbQiR5pD1uoLAU4//slD169OMq/7RcYUbvtG2mzwAPxPXW6HSHFs7Y3Xbbjr
cDEKynrtUyeS0HfhrE2dI7X3XxZ4O5QdH8JUQhIo+M7fU7wgz9s3f5vS3nb/3SfNker/+x0iFiID
/pWeJ2yp755c+1lDg+5J+97OPtQ51rkIMc1a3YP7SMwUo1LywaF0wBUgB3qGEt0n6RH86M7vUWC/
t0a+Zlr0GryqRwsrUIQDCFLJF6e06wQClgl9p/M27HQijkWDuH6fVHKTS9jUY/RiQA7f66nLPXlk
87qWBPgFU7CGoavBaFRlq6b6l52Cvar7mJyOggS9jpN9+PZCaZSDqA88V6My2eUKhA0l2HHHB9dj
6UYOGvYzKsYMLqWMsAobhmV/HWqtnFklmaKF3pzXUNUCu4YVJYgp/NqO7iySlryfw8zCPVtdZ7fd
V9Gpm85zDKrAoy+1vhcTGI21tjTQqrPOpfqhO8cjw8WiMm5BGE+dzkTmhwo84t255Bui6E2lpKzK
5ya6hRAOrPbFdgaLUnvoqL2wMbl+RTJ7MFyWXer4E1ubpdfhlsBL26SCyqcKNaaefvW1zRk/WAAh
k6IG5GCqw3KCb6BmeEDgZFdMeqKy1q/fKtlgA23MP7QDCxRjJZi9cOePsKxI9/1Bx3g1PsfPTBVp
S2cRT5BzBrFAsCTpoFnf9DzOFmcPdtnFUCdQMm9jIt4a0xz9Wn8PRr/Qt37EoEeHpCXkDCtHUpb6
RfVgCFIvQbo4B46T70b0/VQmpd1rrXYrtlNha6I6CzPbuR+F2/Stnk72mGo4Z1WX4ff7xDoyOQKM
V67ossDBQb3Q1WL5Ug7dATMf5ymCtNMxjB4G0fKpdWxsi7A2i5V63BQ0OhU+hfaTg9+z9ZsJQYwM
wvMU4nvXVLO/hayyvP4U0qb/P3JsMA0YWscFGmHdvs1Gmiix7S1a6ggE4ELXLW9z6kuZ7wd0aTVj
W9I5yfDcGBKRtCYAtdDO/bQs3mqZXL+dNUxpDXDCvb3D6St/4no+8xkkuEMSRS9rByP2v1mfDaF+
RPJH/5xHLxx1uNeDJQzQHFSEjOzntLktp6mBjB/+PBKS9HqssslZtrbnCiaQZ2xYw+1WdTAjuIEE
5niiCKyS4igivQyWPO5mvLNLq+5mcJVT25R/ibGrYNXBskA58g9O82WQqbe1M+qxBnHfu8b55yUJ
dJpmeyuD90MLQ1s//mFnp1wUOzQe0EyJJ8ZsLzInGur0Oj6n4lB2PDtnxfwSHy1jjDf9csX55SfF
wb19MWvTSqJxp9c5seCEaxEY8JQHaGoXKphh2eGWLJQ35M8PYUf6g3h4cUA3qgiQfKlkNKrHxgxU
Ms++cehmKRRCyLJiXgcwgckH9DFvUSrHa5TWBqmVxDhUZfFSOyQTE5tAtWpeFAggO0waBZh1omTR
L4NjISvbQ8W40z7mtR7kktD7Fv1WTfSQTEGeTd1iluaoHQQ9cr9H6eMWDa+iQV4K8kADzIrRfFjt
+XVZB/qtUwulAy3Kq4YCZ0W4TdHQkXAYvBsDLJDH1QFDGpi8zHmnvDmNh5+AqbAvw1igZwRxlspj
Dt9AIgCsmvcCCa+lHNV/HNeuK7KX9o2xTb9/zdlBRcIqbrd3dI7653kkboz/32RAlRtitIIQfR8g
47zH1mzXd3q+aADIv4kdEw4R3yFZhD+42IsQHBHnDUF9AREYJhT0JerEVmi+XedqmzGqhOyc4Z/P
3YbXsV+M/ewOV2rgkKvFDIgviwJp32RZeCGjw8b4gNw6CapK8iBtTNrDAVjv27KlDgZk87Klu1Zj
jleOYx0jIeMAFE8t0lK+52tLrrrBxXreTa72iZPvsIcqxyNRKCjHqh1XYiGn32Xx5w492sbSLaEj
At0q6TV5/qavxeKwT/SzsFZ3X3jgJGLNr/bDXR2xOcmmD4gVXMuWgKjsufKmVISZp5wtExIt6BuL
VryvMS7ZUUnbh4ByQURM6cBce4Z7onzeNYxz5ohKQzPTjdDZhYBg22BLdbf5NK7J5dLNpcFxyqv2
oX//XZJJGKUG04GWwejD0QZj8XIfOUyCV04f99wJ3v7Vw5gENCQtg/p/k0BR5urnndc8yUWsyUHL
Y8VVlJGxtcsooMx+aq8sUsBquivWQhvXHgoWHOX+VPd+hEaDniZZSldG3TK0WnO7Es/oTnf3lDCP
5gaSfFEzOOJhhSSR1dmsU8DaFys4+LXZV+VjTTlucQnYv6YqrWxlqse6lmw6PjLRp/5ahrj5RG6e
vb6+ixBDsLNRHiQZl2j8DMirhOaoy/wrQgPQpgUCrGLpePipx7XvAl6dZfF6HQkK23J7VDHW68IK
i/GsUVfoNdthb/+0uw25+09kWXHVbxpl819oOp97JmAu9N0fjmv9oaI476pMk/T1XEyaS5qMDBGv
foRwUONjg8tYbeDCYIT1DYh/IelUeEIcXN+hza6owtLGltmhvBWL4czgrWcabdw559FY2K93xdQu
I3TrNNvbA4UofVp9l740f8tqnDededMXD2VN4jIahefmvjO7GwdE1hAH4gzWug6CGVx4PpU7e9AD
jSrufsg3G0phL3KHRu5KKvpALukP4vhcb+Pz+cNeD9NxJtDdKyw9985g09Umlb3tMeC0274s4a9e
2O5nSD9yDvOVscdnJs5p3IjgmGFJhsOlTU9wXEpd75jZlrnBkRG0MsP4nyTOfWryLbBQaYKNkFb/
7Mr8zjXLbmY7ucIOXfyaq9YntidT0OiLGKQWqH4PW3Q4oQZ1JHT+oUhU7LXXpIcLhPvCO6y3F60O
CjALcof2mqIBWOeO3tDF54y5KgwpfPsRioD/upYOPmXhOdDSg/wbDTvG6TezvB6rTU79u2mlkBMB
m0C+NBU5Aqtm2/9j7KatSbHdTlpyKsBnlbJFW5NxcTiqHjzp02FfYu/HqkJkaEJyH9jTbPe/CEU8
THZ6AZoiOlsScHQivP8S1LIB+Lx5QMYWyKBJF1a7BT2z4ue20awkv5X3By1lEm2neuX3Wgz1t8RB
QIFSmPeaHmfKYPA6be+snVOr2gkpZOsOS/Ykic6BquC/Gb4NWbkixQSwJUsI/lDhz7q8VhjX55Dh
wAO/NpPbnBY9CldxigX6mNEJMjW56SokC5LE3ZD6i9EvdQJNhUlAdD84v4fbj71vonPro0na2yX4
SomQ0tUJFDaqSht+xvRXYueqVGKl7CjYwTFIQBquFbBp4vnt8qoRmk1dD8NJBAvQ8+RMIdK2Hl5j
xnB5C/GBqCvJBLSXFBqHwsrZUWkETOvPosiXcgd4n9SvYoTXYUbhqwxFdPT0yaJl2vhVwswbXsrG
l7GloIq1TNsS6gkTGQSuYnRBqADzuXGRep6miWIh9DzOIKiNujolh7o1bTeVqTu8T0HVgwNWxYlE
78LvSYleEseO+w5jjyONF0yNthoW4XdI4QMOkv1IwNWH5FlIx/X40oy9UGMS8Zf+14eIR+pkGmbL
sFp0pKRt0VyXyTUF6FGp1c7czFbYa7LT+51+y87LsvmA6QQtMPSpek9AnMqAHCBx3O5e6gDCNP8I
PncjbkmM6Bd6FcIfCoPKUoyU3mDzP0XwVOc4GnJ3nVOTpnGVDDnMABIol4Rllv1fdgQKNKX6zs1R
gXUBGXVJ4L8jqfI+DfvjfOhpMwIKdZiCSckvrg3zgXkig+Sb1SvCQlLVKccS1XbEOc7oFF+jzP69
7I5m5qzevNVA6qVSwJEZ9eFs/I+f4x+jlGZ7cuI8ACOjXgFNMNflYRoMbOFWBJ9udtRuttQn+I+m
S4lR8ORP2miqXcTXUHHpedW9VIVP/a9gz4QYiRmYgS+pzoTuwZXc9WLmjDD71Dgfc9kocWPT8PV1
hF8ayriH5LYPDfojp+ynNjEX9+BgE8vQ2LtViWREA9pOEonjqJ7bpwCw+xQu611+wNilRBcG2Of1
dGsBI9iLT1/nlApFc2X3nlEjZS01aBrnCXjLwvTYsgZJVzB06jcrPGHkfpxTxSRAbKuRQcPVKSpq
lKXLxUc/KOwuZvizudDU4FGBPwFtee7V4Itar525fzHVmfkMlXdQWHLq94ZkPzo9qG3AtXPhe5Mo
JSwbqcR55nl0+4a8wyUJzIsLLlZ5491MCbqFM7FBRxwpRb6oIkwOOIxfn1nnMLmrHbYesxx4TOSg
2Lp2nSClYJONFptm23ahlosBxS2IAhrEvKfnx4p3Lg7uFIh2EwVbzeZTT2j3IBqYt9yDJXHAljV6
1K2EPGpb/nOv2DsKRx/4xV+t62aHZS+8AkdqVa1MZzbF3suZRLhvlxv+/vVwRrr4GDTaYcbU4ld8
fi9O4sKyzxfHLezgeSUuX6ITlK677tiLrsdLG5GNPivAwqI65Q+rKQpEv9hZrq8XJsoKcBpjpn4w
mg0qcWRtCIdreAxjPAYtLOHbCTVx2CIfOcOQ2eq7IRv+uUp/B0+XlcfXpZt2Ktrjp7gGC/N3U+dP
pF1P9lqyKHcj6xEXafC5vyY5wlU5KLjsZLnvGDy2SZLtVoOieAgHGDoi032VtsfuLn7C7E6F/ssu
oOSFcY8PIIDPu2ZNoPBJvDpNEjNZzmJv5sY2HnovNnrtU/Th0Pmcwlz/TOGGQr4b/HgZ8+VRky2D
/KWr+zevN+ck71tBGzdGmVSeoE9RHElpD5Yh7TSO9iYqO6TaZzCVP+N22r90GJXcbyTmfuIgs+uF
GfN4IYpS0OhL8wzQdVsloPfkn9kPFAx+5zRfpP3FlrBgG0na7TReJM/PHMgocp1Jf7jTCsjUoJMY
BVqc0c7J4vQIXLn75jzgYJcfvKRJhmUfb3Rb5tzbM3ewsFckSrc6wY7omjwhc2GKJEiyBl0OMOPy
0ONQ4N/qjRSn6tUi6r+Nvab4qkp3o7FLis6zD6OWQD38svYYgSg10d5oSBUC199YQtC/kVJlPuXo
GmnkGDpFz9bGX7Cdt7syLYtUpeTPXcjmH4rj1k8ST+NRtYRSxSwb6OufW48zhLNV4+Pufrd1cbuA
IdTaeODvGwKlaTOJ17Zb0mFi42ugcWW6dhbEeo3txgYsVwzVVLd7IbBQWuTfcRqQjVWnUnVvKC4t
OBRyocTzkG//4eosFRT6Ki7Y+emCh8MUytP52e2LjPkkj5Qq9C69XKgNL4RSHU/loi0eT6wMTVjI
oKUXFYTWvpYIilmV2sky4M8C1HURPO54SfT7A33W3Fv5cQFyfgOkogAFl6kvQCS8/0Y5OZnhMvKO
OWMcf20NwMLWgazEZ/ODQYbBCcOyfMCwMPe/sifZBpbCW0lH1hXhg37i+wEKGyMj86KopzpVs24r
zre7m7DvCbL3cUTfHIzwjqD0hx3t9/hPwTbHN/Ki0TnlFb7qy4xjxfvY8zMAsdO1W9QL5/qdrylp
jOhkS/8dgrKFY1SVSM6y3fS5LxoZxJgvkunMhiAv0RnO8WZk3ZSSQ4QaobChoWY0j/NxQLf7uiLa
m1QD1W6pp50vR0OT3TkHNNL3AuK+EKjBZH/NIhRctzFDlEFn0+0/0K5FWAClBkUMtaIzja7YwaSZ
ZVPJnxm6pvoYFdwjjfoMQwUYdO1IpOGG5+VjonDZVMMd6fTAnVzfiSPH3eusttrSLJELK2lPP+gv
Ex8zA9npCUbMnW0fxtie5+GTlYMGkjDZygC0BLaLtAsC1ntUKHlgum606xpcaQ/zAo5QByav2F3W
XK2e4FZNptAG3VpyxkzRay7vymFKcCE7l0VgUEM2TkWMlGvozNApBx4k64f9Bes40PBdXKnXVsRF
4DwA+iIX2r4wdzV6tZqry4abayrBxjHw+MOxsOV+jfIJtt/g3XFgdhVEeHgFZ/UEV6ynIvuYsDez
7MArzbuHVxFZ6UgF27eGUBGUBvcc0OHCvDqZzEbkBVG+90/hFh4XorRha2rZR85Gh7QwbGImy4kK
obsxHovxSOLUi7+EWiZtZFD5EVCiLQcw9+rwDyDZvD4a3/A7ipEH5zOdjgr7+nV14yR50fwyIZXX
8xfQk2fL/FAn7p1WBLD2FwCxu8iY1aZMUiMv5PmPwQ2Ds9JykyPtyO1PNK8tuO2KC9K5doeNFpjS
9M1r5Z5dIhNkwZ/r4lFtbfRHVffliFCoUmmmGBdk+HowoUPiCrx7epud7Cf5fD2mVhXGSBOSCPE5
Gsjrt8eKwb0q2+A2QFWJPZ5OMZUEPiNdI4E/mBoQg9FMc/PRvj/da+JRM9sFrsE/MOzdoKtM5yrf
/Xjv4T2OO8ib4JAfwQgSroRWwQqxJ7z/n6BS43ZlX9vW80QT+6eyq59WnAOSGtXotSNHMZr4VsA6
2PkIn0hEfAveW4XM6h5IQ6TL7VOzCUAwD+pTJzRDwVcK7IX9LPGRiPodUmHU8R3uOudcm71DkBgk
NLfREcEIfzl6p0MdgT4l2NeLf8DURi1+Pc45ffKeT/6Kr0wVzdgyBfEbU6UcPkY1QGLnGe/+tcG4
6FJdO6DVzUS5JsWqufZwj+kbdWNvpNQ9MKYp3iqQ5x22PQhw0g/+3vhEZZ5KTNzerysQbKSqjdxi
B4v8ZrhI3Xd7X2v5gTz1EPQR3wm9o9GOAqo9uNFyJGIRsW6zsC6NmrqDgtQFiS9yOuB6nd+2fLYq
0JAhWFlUqonXanVWvCw55a/YfC5ZT9h/GFc0emycZFZCC24CHJmyjtQ8InMK1BOYOHWy4ylwFa6W
+SzJtnijcHj5Gf4eJzCK9vx9zI8kE2kRXeQTBX5GjT+MC5ATw7dGhHSZTMrsvZWHNJKUtK3eMHAP
0LJdx0z3SN9O9M49/n7K8K/51LLjxQPnqz4I5wMfmmQIVEUB2SmT35sY6GeSw99PCVNUOKg2gutb
HZ70OnuggjA8m7d+gye8AIEvcdIgA7Wt0ppdrQwqCSCmbpII5LNy9Ectfzzy8Oyszny1VS/PN5V2
6WL6QzC8yxzoaVb5ul0mSdyZMupEFQn80Td371cXFMWkjQGRi9h+14iMU4Mx4Jth9Gdi7/axztHM
aPnCl99nTeJZwY8x3ZuKzY8/JVfZhmnjVeqgqD9+S7L4XetE7LsksY2NazHJNuUwXAT8dAxBOJf2
xpGBdS2NI+AHgXv9x0AgBE4iDghvH3CKV3RsGZdRooWWOkdG3mvYH0H4K5V0EpWKQMNasXZh7c9X
hSBajNR1QHHSZfFPUiK77PO5/x9JqcpxXZ3My2x4CoBNPfctt91xJAL019g16k3ss68Q9dXvyiye
WX2i3yGjaB8JGE5pmrznNhsrXvl8VY4OSjeNz9KQ1rjez/ektlgEWba0376KJNWKJoFEkgZGzLC0
OLlXZU9GSpgwUbIxTrlrZYJr6WenAyTwioXNZBcR7SKOD/O3nJIGEFznK8R07hjjaA3Ozbh0UQ7Q
qQZIbAkmrS1T0YTUYGBryMycDwc0WjIxrfTwkYytDqmV4BZvzvZWk5ecAXWrhpiNr/qBvQhmcSo6
zNrRukDMI3ns04sBfK8rCK4/+mLSR/4jlEjFd0gN9x+lNieIxwKtGYs/+h3hxjjrUYXnSba7phr8
Ou6xI4+z3XJC6ZFVz2xBndjjp/fqo6a1HzFKmYgcO325NtHojldJO0Vtf62SbtxEj001zncb+aw7
UDQxM1fGXN94RNY+JH5Jm7RNDEpkOknVGTzQW3sDJh9g5ou1W5ZY7fsJQop2Jbo2xbBKzaYiUz5M
RgDiQdepU5SWn53JcmjxAm6swqFMoFckwQzaAykNtUQKENkukf2r2vsfSovr/dMJ53fjPCt5saGS
81kNOJszjQ4IZ5jJd8T/1tjSYq23ERGoIL/nIbQjOaRYc61jZGFDK4wGuuKL/mr/wdHYnoIHWsIY
/EPNuJldbah1soAqCiiezg4KDpN8CtERhkT+uHMiWftApgbuKKrahowP8gjr2OvvQ5AzhIPN707S
uJGfYQdPNPwcT6VAd5UjEM/zbJFUE+ZmqS/HBM+UX43FzFWZB1bJzWQhcXibXDUonJe2EiN3BuaX
rKz6xLEXUsVE+U0USC5YJpfZMEbhX00vx11NsdJiNcfwuF/JNCbAz/trWUu+w0/YFlAk33XBmKLD
jKpyCp+UxfFZQfPh2cwcY3cngOl2RLlvzQxQZC/TQpWuTczY1SMCb3Bz4sb+tuNrA4PUUQoU3FWB
PDXSxQySs1bJCUtG4hOvMPe5vfanPeaoV4x+tB0Yi21KbdEmvanOUtJRN8FTy/Oze++vdakUdSGb
2HH6/5aWqSSzAJT9kCGEV9RnqJSLjQbKQAyb/Fkw08L/5cxUS8znc5aMrpLbhLZguwYXLhMsCB9P
VhrJMUBVDIjSXR5GES55+zzDWMcTWvE7DI6khqvXRZvURwwZki4JD/RhwPUA6EA6l63wAxmB7Y4m
hkPZ8VSlP+pF76UJyUXLq5fM1x2Fk00ELlXJ4JovnW0YCRCtab8vxkg6gWmw6S9Zn31qDz8swMov
hSvHpNZfJkjUnBDIwbTxm6R1JajONNcI7sRg8GubdkiltOW/aAjvckhHLMxvLE/HAaxfjLJub0qS
tj0sNuZYUG2cEpMvI3tnBgY1NnR/uhV2KpnPSgfxGAf3et00qcIWeawwjTIdEfqSf3vpCs9Dzkv2
+F0hWEsVj4M22c81Jgg1LX6R1kvIp5PqPId+h5YS36Z2iwR82x4Z/I2CEfh/KFIwhrKqN/JwmwVn
vjI6M1Gi4kNWKNc00xkS2e4Zh3HUti9uN5s4aCMZ/8t1FCB9djNeST1r/zKzsEn5WF3Y02ccXB+g
t4yOzubUpEl1rsgn28JADF74ste1Zy+QJs94AYJw8tR72u9/9vFJGbag7agIu1fZp0mY2J6yOuGE
Sd5P4BfsOnRU1s3/6RH3EDwxrAP7C04T7rlki5hjWE8Qga0bfTkt2uG4ioJapJ0o4hiv/2c+bMjP
+WoQBstaW4WF9poeL0o+nvFKHIeQkj/s53U0LFfTEoOwIvgu699LA7yyUJrWPuya6jgRNFAKfzV2
/ypXanyO8LW/lQKM8tQNm/RnUXSIzGCdWDk5p9Zg+k2ow7365PROdRX4ro2lEOwHElBSawP7rrTE
BXiljtLtWT2dne93QysNbjlh/ieUOf4mwAIJdHizt6m5Un4Q/7vChGarHJRhGRjBW0XEJRDoI7fH
hz0TgxkUFDmh6UOiq48b0PbZHRuXfVdD96X9mnOr8doMnazo/NwBqAJGqZIiujIsBqOp8ZMQG8yX
26fj6rjRdK1e1emw/vCUM0gFW7AJ+rpgU2jc23ShiCE33TKZsd/oL/BXEfPYvBktWGNCZeXF9247
x+l9KdIv9pUQUNPIWks1PI1XdZklkh+GVsTlOWAAAhgA0jHtPX+Zv7XaNLH2WqrmVJqhWM+81Vvh
fHOh0Rs0j2tOEPNgkzysg+2fIqcjuMM0bvrUxQmbVEUbIIX/hmF0c+N8AATBiliGWf5wKg5rnG2I
u/0Z2dq+Wj+1/U5zbsmHlyN22po3+JbLFekA5+PoZZ2h57W2x+BDdLwa1zdYRWVfL7ShiBTdGYzV
H09wkyBhws5vZ9+cfnRrPZWqR7RPFjcasXyxtF2bTvW/jR1YeaXnuEWKqiTZ8zxy2ht52K0v7gga
KO8mE5BNO0KAtk1Wae5ey23Jd7ljpUuv6DCnPeG12zbIrtWDG+s+zuy/q0iEBiJm2eZWQ0hpKbNl
A1zeCGko9VL3Zy1xkT6IIQcYyYsjHPSpbfvQkOnLy0/zcC88Ss0UNAxs4PcFVbEFUNlBIYGV/w/0
jaR+RS2lYoYoqjLptROi9GSEx8OzqvX6b4VnGvJl99BxsiNnWhEEUew4t5gKatWdqCiQBPbwecKg
oUpMHkd3tqlExQDTBl8FeXSQ+CIJYgqFpmnR6TY3TwU3K1Ijzn+bNfqjfpPDWa9Ugk4axQnF6//j
fVy9XrZtgl1JMjuOnlKyjRYpTgaVQWinaExlZNI2R/FjxcPLBnj4Dcfr2UDtf9k2HOkKAOOJt7aE
wXr8rK+MJJXDSQVbcnEwIyXe2iWb7QkiSJ0a0wQ+8lKeafd3RM1VlXCBUdDl5tspDe3M+hAlr442
oe8EmuzVGtdUhqguR5hzIDt0a47fj1fMFSPKejOiaIxbRBBgVImhX+wXdh19+CvmaczIZpx7Hzlv
Nu56X75XfFGAbDR7lOUI0UY4/52rjrN9YCeQoUl9mRQtlrRpDviPbCurNrLChvCF+3w1XjFfm1po
GUnos3TTahI0LeuI3zSGqLq/Xc5vMaztUUVLUpmk/sQtzarCTZzJp1Nu+un9HIkQhF/17JdqERx7
/r+BeInMq777T15BKs40DEL6DiHLli4xuMXIvtK/9B2//dXFqJlsXEmn8a7fdlDj8GO+OH02Pf8I
TS7pSBla4dDcBYmNrt03gCoAqRIs2dUZchMUGnU1BTGbmPkL2t4n84ExD62lg4c1s0eueLnrD366
lM18j6L0+9kFLnN4jRHvAxzv/KDHkiRqfv7lTh8ydO18UnoS9BagPLqMGI7O9ru7B00Rr99PlSjq
RgfOAmvNOzBpOWa+4SGU8l2Vi1qO1yQWE0h6dE1LskuZu3gtLJGRZJa1hqdzH117Q9JKhp0I5SX7
hhLM0cK1k5RmcekCPTtM5yRS/bvbRkjKsihWrpTZ4Ti++ABOLKE3JQ9H/v78JJMkaaAEb4ovwV4U
fOZjDp8xNuv+RsKqGv3oIH6DQ6+L5CobI5LKHYlJe9LQD7ihNuvQYDwDwq8uEFP3CJHWVOYY/KU3
PVolc2d9LukMzY/i0wc9jDnhKf+djvXMuriz8qAjKjHn585/lWrHdHccACGkvRCuxe9ZgwU/TPLm
N6xqUvl8RlaoqOdSEje6D7kkRqHfSFns9Kq1o61rvf227dsX//QxFH1SGsC5wVvSfE8nstebCHZ/
blO7Jp4EcAnF5vbcSn0HfK4Nzp3WlEuyFfgB0+ojQo/BLL/p/VAddSVJS1g2pn4hXUTx9hvKVzoH
S0QLeh8ejxiI2JunUn7T4FpET/8qLelCChyOBaklhYj3S7IlLq2rs4G6SuJH8x6dy8crtuaPbUL5
MBDKxf/9OVrff19qGDGFNIfcfAlpgDSQDmveu5qYlA8eIWu3Mr74ZzMeoFE+LcNwwLnqvFjdrBRV
olRdgWauOku/DxvoPi8+uQvUV/0wAvXnaKwDlsfDbKnWAM8I2ajK7RKpgs1gmJ34BLBMAY/RQihO
KJMaTUhIpeLWJnRgluBKNOTrz3qX4rI/TPrmBjIY6g0HSkV23GKjOYjK4pnsO9Dg55N5M0iL+QYT
3hNusq5QGhqaMsgnfgKXwUy8CzQq/6kmScwnHyfLvlyskDuuNi24IghxOnnIdytpksycvB/oekRJ
rY60x/BZUW6TDbHEwDJFy8rIh7GuAk+856ApwYAf/RSgCiuWoG3+8/T+DkULfIJLslIvXfDJH2Oi
u0hBM4klLa1nifeuV6r+CXWJishhAFr9UD4aZhweAEUHNxyUrXX1cNtKg5wtyMCBtVDK5Ohxmjf6
gZZsan6xW2qDOldAL2F3J9UqdPr7gXlRSox6jssJHEDygbT9yNNXCIqmL6o9a+E4X0MO14GUFfWA
LeLO5blU8+qNFPtkGf8EsRnOmvPCP2O44PMRaQPCPHqaFF0ru4ITldbqIIAvyWJrLCcifcOu1maS
Gpc1pS2Gz94UuxlgxZa86Tz/U9bL04HXfGE7emnaPZFG8ykkf0bJqS48b0MSCuWuDeVlVWPVEYBo
bARm20GJVv+V4nRZtDBn/Wu54+QBm91+tndhzS1ddgIxgVznzCGNnH+j/gwxgIx+jtJ7Cu7Hf5ba
q0wKsY1mK7hQkUrmRfn6+qs8+U6+7uvaItiNyRbfwtTw+Gb+Xqh2KUETCcF7qZD5Otv+ECuQjYaY
3Zo9Ny0RkUT4QrHaoqpuWLKPK4STIVlPt69LU84RKFfUzjnD6c4SKM6tGbf7sVEdUnWzOX28tQpj
LX/GobuhSH0w3u8N5gCgp/ckEIBOlSico2W+pRbZ28Uxw7/II7QR0FqqR7yhZ3v3Uyzcl6w1aUtx
vvmrtJvd21hwuEfc3QaMlRzz3lP+f8/O/AKXEC8in8fSSz6icJGX+Gdg4wOAR0A34FvIn6RdQZa+
T30lLa/tIaf4g6EhAZLX8jFRzHKx1Qzi/qIH15eV+AB6VVZ8kVzgpZHMS63R+USwCqiOE/yfS8v5
CGdxNVHCq/Z7Frkx6jvfaNA52s+UNm5h/Em1OCXxfpUXECQYkCHpfrS4rKDpR7fz0WpI3Cuy6dEl
JjarP2/nx9+p83BZqjHMTEiHp8MFpWFONiyi1mNW38n7TBSiFi2MkBT0sYTKfvhIXeStUUrz8bUr
YRoIXZ2JC+os2z3CwFYOSrogZdt+SDoaw5WQ7Nlepl6sT7DaaQA/7mae4EciVOOjq8XXiXkRKTtI
j+XIwNlxnhzqkWcW2XDqxQ+OhMCkZ7CGMvPCWk9ooZzS2k3PSiyKaumPiOECZxkIwkwaY5/VG9uP
K7nCDA/cpcQZ81NynRbDabq3NcPLm/s+6zTPTYk2xLqIpLTifn9bIWE5hEcJVsTHf4JsYwI+p6um
fghWnqRj411fbArNuBK2t1Az47nXESsZ5FW6KILqX5YME2fDyTU53Fd8+TwJ+E2VCcyo5q3CWNTL
LN1V9igNn1R6fRC7n0vUuixeXuZOQYvbc7SkUTlxa0BBTZJr22v0gbAJoqdv0r37lhT790PoZJhR
av84Lmjq4050YeCwwi0oIYy6b7rG50PvfkTdqKvOxCUgY+Mx6I6OlSsDc4n/B0HXPRvnr6mjaXXv
jNCB1zLHb0ZfpvcTfHiX3n4SfmehtoQlSTCCmoAJ0ESfKe4n68TjEzTL6MOhk+J+pQ9Ve6EbsFuq
dD24Ut7ueM2IPqlXsYQUWTlB8lqO2GjXA/vEmr3T52zjfOjNKBX01T0a94ZLZPqYG2ptQx6NYFeM
YUSGQmVKvMmxatMzJf69mxruUYV85eeufmXKgGSn6Q/DOKD9/kPg1MdgT99LbW+1yGzH2IXzBeDO
+jSxyVBVrG4MyQ7icseagZbKSw5vVzRadGAkcz9MnlTp36ANxwmrlhZI/rFIDsCRd03LovfMAc2i
libi9/2JuFheT7xkqdN8Q3iGcH8ViT7w8V83RyLYyRHG5Tg72whUKSDcRTZLzArbcGfNsvbMsOkz
OTlBbOnULd57AXdLmbE8r0RSrtY1OFQBuFnnxvysujE23LmE7GknhUSRYOlMGBSMMnPnW2UtlE9q
Jlc5GXhD33ZeGq8Mb9OKgHjJnz7Mw8dcRpDT9JW9+0swkOATocWtBuaVrH3+CFLDe6B7nFoYUi/5
Mi6diVUobS9sQaM1qYtZlF8pfIqcWlLSDkZcnDy+Ke/AZ+hEApKR5Jd/5rXbBeChqWk95Ja8yQxY
DmhDUd4d1GyMROsxrwm6H4G9+96WxcN0W3sXHgLMqqE3WQy9ysumiKG26TFIPKk5xqs7FU4ikHPQ
pv0fBdf/MWVX+0dxCMIR6paxw3a1n3HMtJnP4dzD5JqfDdm1wtk8X51X7QN4gpDUwy5G5wH0H36e
Sq/eJFINcKFW8GHKHgjfHzfORFPoSnXw6JCpm+gznWnnn5v4fgXV+e+yJwgrHnwfo3+J3Ubz04+b
X/V6xg93Ss+x0MTawFULdKhzhz3w9qQQyoi8ukizSpYo+I/72oTr0trXkBiXQamfGXEdqFqsf1bD
FrRVDSXGBaPdYwmGQfeE0EoVNqoHb8thSFfg9A00J2XoxmWwgZWKBkR8+2nsfsIuhorUz/wqPGiH
yUcnbpTKsGJHztDqxqMOsfhFTi9ap/9ATynvXmDvHB8KqW67S2ZKC1pFz2IrGzFK+Ba6UPlRWzs8
/vAWd/mMeUsp8dLJ4aWZKzgvX+R1GGrGj5HLfvXefBgy5GQOX/5+4xsxmS965+YzGW1tdA8NyNsi
OmswchlKQtY7XYE72lIadLwcERbBiVXTwq7xeDcWW7bq0wbeJGxI943FYkRKLhkwltriDC8kbs84
hk3WOdvLT1luTUDfBPxgG+mcKJZnUG9nJZwihl0xrcRV59J+cbL3FcPMka7mSf3o1OvZvQz0mE4z
H3durANCxGxz1LYB9+0H+4CalHefLKDVhffLoLOXrPConYB0KVz0EeT/4dXOon7aAwyloKWSZHXg
QpGRRqpZR0YUa72FAA8Fwxu+Pv7NOqaBB/tqH9gILIAMMYJwWWSkQcTrOgOcEASjwensLFqfnx03
SGdDD5BCf9jmfyRtwdYKX2+fj6CpMG8XUAO6wKF1XRwkI3GFiKkHhIosPDioUw7HrPjFr4OWWWv5
q5VJwJXI1JLY8/bHJulveqd6D16TrOdiznrGPTmvM6sgQqSQa8VBCGxh5p7KwE6QjPbeEBauYSez
yrw8b0tAsoq15qC4u5Hk/jKdEx6HYEX42a0c4zsLJmNbqpNHfZfeL6hQUy0UJ/uZjSgB6MIQPW71
r/6I2Tf3SHkzKacG9O2MMwnajsjfDrWKT23Pnf0KQbxF/3toOAOn1e4ladZTlOA1oqp7V/dY+xwS
SzAckZ7w1tIUrdQOZNOGiBrKpaNco6p/RnxFaEKVR0v2z1OAhLJ/WRF9X5INADX0yDtN0eL+SC1h
BBmFlgwGSZ4F7G299BetJN9lhZASSgH9V0fOd8noTX+MLxS02bbFFOCZKvTccq4a/EbsFk/o39H3
9o50O9EDnfXQpzxCmOx+PPUoabIqQOidY0My+xq4Fu3Vui7lP5fgKrsFtknTDGV9Pf1pwFmUYSQN
p8uLhuBaqxQSrTqSBrEjg1Q523YVsKwbjJbAjzMN+r66tBacK+SCdJUH9Sh3X2pyzSwV7o2moPoM
/AKDarW1Dfo3FzUk6jQlOu4joltad6cUPrTh1oxj5flE1zYLIQwMgQv4u3MhF2qELYoC0ytEdM8I
OYZ0eI/skpL6D9/22NhKe79ixJ+0H8Jpgy9wHpJ+N+uxOHhmZpqix2L5qsYQBy4ITVPckwZfE0st
twrolyUKsCvWbjsFiUb37AjXBhKt3hGQaOpbzFnTkPhDf/kao/j+YJeLGzWcU9rYiAxLpFXmzS21
D11QDPPqfkSYcVPjcfJnH0peoekC2wcUSAfSvE/UfzCwkdAHkRHXmVCIoVDsM7CBVKsE4PIEgiRD
VUV78Y94LkQar2TY3w6tV9S9dIbSkuxqun9q5W9LwKh8xKtfjutX5GyKxdW1UREY+GCUD5Ve4N4Q
4mz/MWsille7JlIqGVZ1NL3qDavf8flv7PgAQLQoVpxJGNRb7jn1wJxJVuhTqr2lF8NjJ7s2sXcl
ALGvbFQ7P8h/4ImXbOrzXapcdz1Y38g3IMwH5O5zXVwNtbOq81bD93Ztx6Q5IiCacEJprQhseFO7
1yN022eBg0pRtvfXcFbNwrcs2KAxFv6eqv0LfK37Q2+NpX0nm8ti/HwFoimHhy8nL5c6J5/yKOTz
toqD4QBaZD2sihmIg5H8fyRiu7C7r8J8ZyyDfjbgU62uaeUpApLGH/1BEXuVUatZE7ago8j/IK9C
ZWFv3N634AG+X3X0KGFrL0URgwyeLbCz3eCWI1Ot7DjbB7tkRUTwhnhhUxC8BwMl5qYiTYyXJ7cW
5bsjT0QYKIXb39mhUEkBwD25R71bZqm7R7ylvI2OhogMGeRyvPDircwMWHS0X1TpB83aIxb5UkuA
JL9Pst3x8n86C+Nwz7qLfjJbyNRnZ83TaAc87fI4r+2FIE9p9ryYjNg0si8APMkVmFTBBNq3rkNC
1Tyjk2pvDWwn0ZfgfyAouI0+aVNpDLK9rL5xJ9KAgtljcxTTx+b13bwV3qFzB1YaCt8pFvJSXd7/
hDppqYVOj0n3LE168jL1tY6k8Dahq7mQu9hL2518zFjYe1Vl+jXUdMdP9XDBSJK3UwL87ursEkEF
jMSFNd0IOuxw2j1AJ+BZDbmef+mVskwDosKopBuyJr1Ph6487Vq94/giOJJJcfjL6YrUszQb6dlF
KV9DHQGsUNP3F58ok6MQ5Yew39Fcs6Y2E2CVqZIj3FylJcBs4Gg1tE055ekTYo4ewLwZSstH2jop
Pc/IEV47tb605vm+brdvC5HJw1iIdQ6kG/dT5qkbDRe6UNhoLfO6/ASrXAgMR1QMwW8vpc91Hh/j
m7lY6Q8XZP4wXqXdGzNA8z7h9PRvGhLYxQFSiiu8yfA3Ki9H6aQEfvwpyRB1UcXJxrAwd/qcFDFK
GNArm5hpYSFftZU9EC7ahMcWp9CL4nx/PYm07y1kK9pYvaAr97FHUq/dxDpnJRfk+LoI93rLOKSK
uEiXKTTLZQIw7BeXFK73+r/5N/zOufZDHxKPhrLsvvMXfdWdi8Xxdm/PwrjKMKYtkxaYW9kTbKhQ
1c90VtNiQGbhAL2/i51rJEXBs4yW4R93gwAfXlrxkRdw7xk8lMpLFtUGzQJo0E21qCm3BaL1GcP8
V155AVPvKFRcBR/1c8lbEhxIwOGioiH0jaaoy87p5JvDm75oq9frchR4FQAslAeeI8U3Zkxdm3T/
ofTZrjMIZE+5P/R6UqiJ3jL/+0YSw9X0XCEKbQ4tJEfiM4CUVF+8x7F4zhs9qfuy1BXOcqxqzcwj
HzhmkDYFG8eKq8hTUwkq1U/CNdnvAsSf4/AxhYIvhTaHYXGoNjvdXbdAtdlw2IQgo7yjMyNoADRQ
eXTVjSKwO9etYRzGNmVcq4AV/Or4mVNh5GnPjexmcOtf8gnWnUjCpBWs/b01P8SXQz/y5aE2u7Lj
jp88EOdQBfi9pX2JtkZrYGVsxUUSQ4nqqBJFyZUNCYdrXPP+7aJc7eIiEmnRE5sZ797sn0Zt04TX
hs6iscsYUCcP7taOpiKRen9GG+ATJOfoG9ufVVhGeP9RSqtaUwERKTHELgTnKJngEetYDuGIxEy2
V3rmT+U7o7KO3QcPB/e54SOhiyK/XnFeJ7x+NXHOqFT6V/KzhkGIAbIEZKjmu0YzV824fMkV2pn8
94e8aTjvqe9z83RVUWCBEUD0lgL/5FNCN1uYieloCUDQIbs1Q7+hu0qnAcPsz/VK9slpNvoDMMxV
nguYPU74n44tLJiJJUPBlHTpGMiX2i418Ensd/8rdOj9gBHx1HWJXWZZFKCjlthyQ716xHGf06b6
Cuhhvl/VBoI0SnOsUVsXi5/u4HXToofNSthH5qp/842FFAQ2vB7iTAwpMRhRltN8uYqE06FCL2w7
i86mpRP4l/JBOcTgr45uNsnCO4mSWU+dNBCXcpK0+SlB1lNWzIdvu2dnwpDdSzccfR5CWP8hbtgx
8AnwzkzVK0jiTmVUSLURxAgetI/06Gbr+A+zRunZpmu/BCa3i0rG2ihW+Ml0uv6JXrl0+Raudlv2
v3iQJGaDoPXsCg5mF8QNoGazWu6iZYozIg+NBjfhSbW0m1sV0jxyUWN2cho3LkwbqIdzQm2m37by
j2n7JKOJk9kxm5Quwp63r8ArOtXYWwDcunun5w6DD/UqX0LhGBK9GnnECwwLoz+Kxp/CBvcy1LD1
/G/nrPTe67usJyZfvfBZduABs22JAlhaTQY3uByHcoe7JPQh6GitUvZ9xBSkWp/MfKO7DiYynFV1
+gQ7xaMwOcyGdcM26d4h70pZF7UhVXp1R/GAMjj6K/X0gpQuKpKzpn5pl3LL41A+Mt5yC9PGR6we
5gUXScZQ8Az+3LmcJIZemd99fQ7MIiwjgIxcp9ADcMGsxIvTs/i6rB2vyImoQ+bLNPEtrUSY/R1y
F0ktXQ6Uo4THu1ZSyBA7JuX/xu/BclFAa7w/+JXPgXROu2qh4lSizclkTUmmovlRz7oncS1t5R27
JScXhSBmIQ4+KuG+RezUfdUPOxZcFI7aaqghpBAPIbhvY5gKerQ1BirLw8M7qX7qmmvMyfYp12Lp
n1Hc2cC5jkLz3dPDWLD3HHGKxtHNtGaW+t9Fc8i5RGxWyN8HaGGIY/Sbtg2VoSaklMYUKZ6+3e6o
JZH14kUhjzKn8b+WBmYJ/L8ydj7uvNK2ccOky7FMkHhdstFlvQyCvi4RxoQ5wK8of8Rv6mZRxW0G
gyXopZ2MgPT//jqB2HFswDyZdZTQAFnStAUMhgjaxYODZd0w/fQOHrbAObbLuE7mOHlCRcoLT0oz
0ZpBO4ADx9EB8OSRkOAavSNmSuov4KJIZZLqiw7wX94CgTp2nOz7RUUnK91yLXACkBOiAflydGHi
XiayJfTjf4QSEHlKRXxgT3YnYHxToPOPIfqRc6aGLuKyjtQW6/7aoSEjFhPuA4KR8GeJpfwpoTRO
QzUG0TIWhICdhUTzXrC+7JOgdBCL2UcQBy/hgUKSPQAT8uXZgXF1kLe9IH6ukTupGS0JSVE3L0fm
2VWw8d9Mt1jaeA9GYZuEjrgTOBt+PLw0pbbyPfEzPiHb9UT2lARkcGlVlofFbbjvt0OSnI/xhVjO
bBwQVf3SmLgYjkdHyZnzazuKT415jrCEIl9pfJ9AnEDIYoTCp6lAm0PMQq14TAUVVuToaT2DpufX
UWvn6VsVnvh2YCkF46k2qYp0H+LXOOMYr3QTXNIdy76oIF4uzm8p4Vy0DK6hZnNMxbLGfZRaojKU
pyFVjTzJH2ohKfiZUFdhFek57YGQhN2myB16YZyGfcBfsI82iVEOQtbmWGM71aYgcF2z4GC9yQ4S
QKFN/c+Q9xXBUHjEKywr8OU3cUt/mhugCfbMwz1SMl4sKh5ReLomfk+qVjIVyQqWRaZCPofrrP0s
rcogMs4JI2PYz8XrCp0cio+cViTRBR4g0HmwRdHTIo8ajSr+jaTjZyJq1py3NwQ3LQGEV3dqyQ5P
KXtqy1iXQgtUqU4p6HApas6zNSLhpDE9czFToQaUVEA/66nPCUAOKG7GyTxadNNeb/yp/JDieIka
yx4ELSPItZubikjoJMDBC2mHgJ9tCXtKcuxTFQjxqj1aUPMRv4n0xSGgb6rnTpRgez48uiz4qIDd
9yzjlpU+v1uQylQr2cZqo8ob5I+S+2gNXDGli4Co9rSeO+1tOJ2TEL1nb+U76mKtsfNa0+mSVcV+
XMWMKePP6YewS87YDkUuyrzXqBJPD12Q/wvhkAHiZUHyBOtEx/edt2ju0SYK3PFiosttIrJDW1KL
8s0MyN60c4ogrcnySgTBtGfJF/3I35K9IvFLik+Hzv2l+ZhodGFMQotYjf0ITcUxxtDuVXAMCds4
WF9PcxBC3eMztnQazQZb5DLG3v1F2LXm9/RVpLK9h6n/Uyx5tGjGHMmv8RAgrAuIDcxEjICndHva
a5WRP4KeYuLcKF7HLLYippWcJ+Z84S/pZhY9JSv1nP9ibtGOSSim23hgNU1K8jonT2Cj6rfl0aPw
TtdOQDtEZkgxj94JSewlGJVvSIFfOWpqwAKgFBWmQVw9QSlQqAUc5N7iqQSxC7hXcdhlGv777WKn
wn9kTeM/B2CmsroMKzkXAfwLUmahJ6CyjIxaVmx/N6d97OXptCDpdWVT+q7pvVeF7sS4VCo/mn3h
BKcMbkHuguhsW2+A+BWQBLV3Q/MynQpbakkOe7AKH7OBdBUKn1cekOQAZAXolHiSc76IA01GDOLJ
OMlb032nnX6sHUZxoH7feB+43qzxBAabWjB2IdUqIS5o1EABAoikw8Eni6byBfdhrTqKm6Zw2xNK
Jq7bMj7z2ywt26aSfdPec/kOAM1q7RvKgpHIp7gMCuxl71o8U+R09z+YHUUQcKBqPiuu8xpQEVXk
vp2E4rVEToVdXq+9huM4vFsxyFA8YOeJs/1cZmT+UkACyaDNJI9so70/3jgtSyZmaF6S5+MdfUh6
XGEumOWlqxBiBexiz93tNO2FO9A9jXtiE2uJTnC0ZQwrIAjqEy4WaZ8vCFYdmBWjQfLJAw9/kkjR
2TodK3+BkGBltaZnlpnsqxon8eodifDSypI1BNyGpiYk4E/aVL0o/i4x8f+KFQSl4mjQvA2iO2Qu
zDzdTQcbbDZLWCAOqEKFjN8CDBw6bF6TMe3XpIdxbPbHri6dJZ9gejC1zmjMY2FajpDxPlPVxMZI
5c9uqkXQ74CX3QEo6MQkSTlrJVKIP/H9juGY1UbfkHwONoyvYcF7sAizYCthmCIYJg/WFjOK+HyW
EqOGFjfIAxSrCWKbIwnc3N2KGzNVxk3DsIwxKZcueXZPge/px5FxqakHayq8qbmC7JRaKOlBYvI6
gsegHib8p+RgBxVxbgZtJ+5a4uT1nT7ez6+QNTGfzqYkD7SJofE7p3cJW44uXvAlyc0737HFujrh
hNnwhKdtbUQLLSyAuu5dWz+rYo5hGgDTlj1Ce0pWISdSq4BKP86AjOCi90Bw3G/SncGzmUgSB19c
XmGi0rLLTgXyRzZrWim/4Uw3ol+I4h5EZSGu0aSImybstgJsDbJT6MxuygBymXbCuQpllah/mj7F
mY85nsKRf3Hz0AHw5YhZUtsbPL93ORYiB6JWBbXFMVzyt+DlFcIpXvM+qav+3BM8KtxO1LbbY5wN
1Ln1LW74WnW8XYQQBLcuXtvUT/p2Tige4kFsoPIx0rwecagqAlOIevdUvniaEkl3LtqN++5u1dfy
MO2ZtGTgugfGIUUUjHmIUnm93aBYGlgVaS7f+vrHCu8BAsOX0ZPn7rdIyteVMgxOS8bSHrEnsZat
0K7ISxe59n4ZAxiJg7GNmXS0JXe27oBLgdvSYVCqOMUJ1QxrmVe1C29qpiCctF4Drk9INfg4Dg7/
wi+qgjwrx7DQG5qRookzI+Fn/lqvi/WO7u45bMmRr8nt4lj7+7QvepscUXRp3JfOpWwGY7Af1K6I
PcTDoXIPy68gJ2zzjbdq323KNlXxEROtY0r53OfMhBlI2BrYFraCroX4boNz8DceAmzd79CWwXP7
XCToQAtZViDnjGxxjBPcEz8iGWDmChbnnItXuqRKZnp89PUGedVDLGST5dABPgg5hvCg8It4+gu7
2SMo/EZAXwEv32hN5ipaB8frKpJPwW9MSBLIHxMeAyqgxT6KnId98TyEoeAo13IG28Pq4F6v9E7W
S1KEHgNTH4VahtzlnJWrIvDQrXS6ptHcWBKkfr3UtY71BSRW1nSDr4QWaNMrGAiBsqISQFUiaN0l
1uFf0/Iop4qhBKSpZOKOBUV7ptkkRbmv6oSNwE+FXxNg6ATwVQ7eDd1gTszeIQ00OmN3rnHlsPgF
OmG16ZdeF1p/aLT32YbctPRLdRw5GQedBmqDYateXKIQ9T0o3aIRIsGau+v1grX6KoUz9YACZLJG
tl6UNAIkIN6o5y/buby2Apu8FdW28o34KRRPCXERu52kupoCxcbB7b8F28+IDwkv8KLbQTJa1i5l
gSqAUbDanl5hoLVu7t7nRgRivC3VhI1nPSz/5WHx8c70paWHWOy/GtSBgjS8X1ZdyHkuZrgxIAGy
SonceKfjtuC3twdVfV7KwWUPBCD+/p5c5YkS3WWtyoJG1QHUxsZCLHTZzGhuaCGfkkiJN6Kx3GPM
RUIA+AbaZPiklxyv3k3PO/f8xjlZaodCQ6zsC+S2iAPvfih1x9Y6NayNa3H2BYujiHxACmOM987F
4oqQ10w8q7sCyyCrjLSd+GyLBb47T7nLgE8gN6jaX2hRfeJE1d81KWoohgPJCsbBIto/zh8wWDSm
McQT3NCMt6jYCapFiXqL1LhlYc5+Itfj48tbGbcmvaz/BpXZfRu8QSb6X1stvNI6Lnp5oq4aA95s
9leEvooLVR6HFzJyxy61BquV+aTA+rpKdsuVRPyR9PeVj4szTkUwUEPY8IO3GegNWFOx3UdE3RSf
KtYmPxgACaH41swhFNQlm4aknEmZwHbq1Yeuwpv3ZH/vfz0r6bwGdj1H6KJnvVrb7EW2/C/YO37B
pOuT3YZ+Z4N+yMk4j0/AmSD9SOZihZBG3TLGtkS6wdmRtCYQK5pE9SeM6Aa9zJ7j7ob/Ou2m5iFm
aEVPNqP0NXvoKKVzLbniiPCRgA744ljERNcamHrcdon18KVf2tdLfwfx9wrEj3TzNmr/52KoaXPB
F7MhtI/ZbovdlS5Auub2TgVeBuiGIaGh4MclKEjuHQWa+d4c3qd4wYPcWWiKZ2oNRA5h1DbcD210
4Deu9FyDynLzfqhKbLUPAXlHO45/rb54+stzRG3DKbV6dpHXqRdnMqWEjnbEOFQY8xH2efDmpBOz
mgztX2SPW8835FcTtFs/R55zI8rePMmIdhAm0dJe+zblVfVryHoqJAyAEW2JeGUb2OGvmFCrPUq8
sF+zboDRqZvRyKbhAEF2xlt8JJRVz5FlBfWNfqFgHNeBoXNBX4101JhZ7wPEkGq46+CHf0KJKvvk
1olgUux+ug3BKoHSF7D0RrhXGJ/XmkarqJ4Gc7SkareA+DrG2rs5reqVeeSse2snMwS594hR6Nzw
7hf9ej4+mCyoOccU7CAYFhsCHHz/F0x7LUgRndDhRJ0oUq4KIreZFV+y5O/NN5rpTTpysdsC98Qk
DR2IUz8Pod8wkR3xzanIMhnzM2QElhk/bx5aIgCAs23wFHy7xWasHqCK4KkvxyU9KI0I2I/F92yP
Aopgebuepsoo+geoxRdlmHSfr1MJE4LHw0k0eMtHsSsN5mC6+JGfsp/6c6wWMCmEALA37dPxQGPg
OaqoDsv0u7PoaxDm4mfM8LNhEhSlz/BnrkRNA8J9M1UMt06ctbBDPc73aUHgz7bl/7mWivSPw+dx
ERDR/7K2GM8bZUNHYoZV82YxJZNM6VaHkm2RlK/mrEFUMFmV5j11ujGiOTxKVp5C1mb4UrxSxxVQ
0eV3QrdsVnmL+UITV63Rj4WstJT7HmMd/cmJJK2qeot2pAZuFYs8nUwT7OlGJsTa5HBfiYIci9tY
ThnK/o4pV9BNTQWrsjjIVLGARnOiaCtfsm+oMPMKQkiJPKtNvMy7cecJAkxpO0Fn0F5Gqb9V5frA
V7E9kL1BYvpvDqICa1wsUBbm+L+3Ejrc/gkYEpTVOhjQMKUyfruGxAim9iesTfYO4eeK0bncSDfY
jkOHoK2kHVJudw2vYYc+f0XJn03t88p5/j4rT6LqLicz68CDDNY7Z4YUg7ECpdgtaTZekd6a5Hp9
hLR6ZDeB5z9mU92+DmqQuflMxBjbXuJu5plhF0uneWOxs0wrVEOBNPi16ESZCk+hzoAaA1IY0oah
OfGiSqN3HVr4RFf3nlj604jN0CYP18stOgrC9fTCW9swfLc+kBxv4eudYXEtOlxXkkjahCg9Z8yS
8FMKoXOhhxqkrhNtclFabbrpSmo1Tkjgmd81GN6zeiVZx/0vBEbWZ4y/VJRKCO3vQbsA0XMcIGvq
0NERxkM2Ri3BZQV7QNsfWHxiWkiHKsSzswQs8aQgLibfOlXBzW7HqTlRqjlMdFxXvVAay38kgzKF
pZLEJ2fSWPlDsP6Da/PHjhR6OUs3puT9WB5YR5jw8ksebSbfVoS2y6V3YKH9w+9qMR8pc6AV1zq+
59pZkw4LkSnAYTANwjXp5lTr9SBuSTFKduzfZIViulz4OxbgbeFQ6ffMQZedIr0DuF6CrLjkt5Xx
se0k+37WeUBmbRgEqmL25n7W7G4QXuSbfQBfajrTmlpXm75AAa2PuGw9c1zUfZr35l555SWTCgx/
a8sTHbIwI+kOHkRcaLX6jxL5F+1O4tCCe7Xe8DIx99od3B49gUQeYFP4YVUYs91exIi1MFHTXKv1
CiaZXsvkyAqtq/PSzOUKA8fyZ+Bqu/rMMkutmHk+N+I9yeUjL2ZTHzMTcDNw2OvpdDybp7whucka
1ncvD4AkHOBZgGGopWiGlGfWa3RZR46W2BJSXpFkPSlToCkzps6K+GA2jNdrQZ1O/bZ+DTRYyLkf
kVZ4Wulg619eu31pcA51OcnasVBUS8nzj9yCIsGuXEnCuXsF73K2BiBy+WteuaWPb/eypzmV2etn
TC5kUUv29kgKQYF0zNuSvOhd24UjIwK5hMmdwIt9NvieTGBLXHVyVstXZL+5RSWjkc2cTwJ4uNGA
mipsEqsxmCbemo5q34SCFjVThFHQ5U9KEBfZU2qflcRyxvleNokslqyjCmNtaM8TbcL8qUHlhR6f
3NXCI/N1YqyllIK9zvqqgr8tBrn2+ucCBAqlCASMXhqA4N5oYG3WKyhYzg1DoFX1go9kxPW6zYci
V7jZZSxa9H4utGy0iTtKdw6eq+aHn1n1hWjYI0MQ/LPrOUFyzYEo6HiW3SReGh/xJKcxp9PnqVEP
yqyfHVsqtmFFN2KnMI3/qvt8Kq7qUUYs7/t2sXenFDynzg79YOXmj0Swq92U9InZiJrLiZXRZBVT
+lOhWqEp/w91uCbBVmKYFDlVAuM2MrgrKTv7Oo+0lZUtukj5/J/zBuObSxFeqvzLlvnfiVXipj99
UFj1jJpSec+5c6LPmzc5zA7sa4CWypOrEbSE5eng7Y7+oxhYV2RVwo10d9gPOQHeepWyO6jufvGi
V0JChSBtd8fNuwaEYCOzgfYwW46pfczKuPMXFzA4qGuewnQqYk7cHI6fA5KSfm7f1I6cP/4NTaiY
4jS/FTL7zQU0Ye+5rHopjDt7uKr3eOJ/Zk036SHdlIRJ00h2t6yhjdQajznSZuBWIAypp9q2CBMr
HJ3Xe47OXkALew3QUO5T508tGYxKCAI8V10qqcsUxSthNh3Pon8+nL7/d3dit2tiuQvhoieDGwLM
50UzoriRleHNGiWNxNaefQL6Z4dsJ2+9fZK19k4iVktlGFoVoqznoHJqB9fMmkVnKF1S5V/Jt4tj
7hoQvDqrPij3kOVNNxzCU0irvzFgLd3ZYwLAbXrPjYWvS6djds8QJoWkJsVOMnc+i6z1FbXb216w
dq/OxJF2LfmW4AJkaB4Ylv1yrsNUT1aILDTnv4fstrSkFrGws+w54GPsH2gAZXUCGRmLckj9hlKa
vF+Yp/T7z9xGe5+mbxY1/8mQJUE8rKPR8l34eEqTuFdItOywcVYx37XyeTzVQy8AqS5djxWw1BFY
DLbCACJnzPZ8ZbEXnyucbtmpnT64mgzz1AaUiPprwdi/tDRe6G4Mh0nibNgiN4GVsRygzBGs3KS6
ZK7QOf0/52cv2RS0Iwqf3GJRCo8YhpouOqrpXtbb5w4u1ug92Zxr38XTRx64eeVJ4pF1OjjGcq7a
ucM2+9iUsWxgWqRvmanI8aLQGn0zNQkKXqCUT+v7JVDHJk5bMNwzxLNyaSs/GRKSDnhqkhBzyyxO
WWTffVhVjYqk7dwKkuIgGYiEX4pAhPurOLxNFto6zQI6kwXKWirI0fe3yRNcaXAUvl0Um6eqAgqG
A2D6ZPypgPT95hlVv1cUhvgcSFS+InwBrV/xdEn5uEc3sIyQ8t5yM/kPLTdQxoP1qYadFGLfnmDE
2NK3Pr+Pjs0QHxCdR8MpvEu3IQnUsfmvRID0sVwRs0pgWIG7Y9N6m0AsRgL1v0bLWrZ8MXREXOO2
y/yvgJ2ntUEHsHHVobG3ceQRnrS2P0gZvaI76IQS8/Rp5B2OHsqpsOsuMJae3lWQnvTUOw++xQeR
vYe9qqSNtwD4C9a1sPUs2rjo3xZPp1/QblPpaFb6WBHnLX6P9K57fhK9jruUvoqnuP7iqRTyii1E
R7RtfOwVaHONXWbrhEwXH2jzabJMkrMGTSkw53E1uCfmZZrof7ujxWsN1ri7h8s/pgx8TXWEeUgF
de3SoJy4/yGYqLs5dJcmVQJwoXdQqxVE0oxI1+1A7AfW5p4IpKnYuckGgzqNpLqyVZzJ56r5UzLW
ebydPukKo8qrCdCnlaDZNRLm2BpQq1mmUTBXbUDeQYSyKAvqK20dGKLPKZFXBF0bztflFCCtNi+d
pDB8HnuY63SQUAdFFZYp3buAJ27lziWJtUQdxUAnEptYylHC0ejNd8DOsBBeam43jjjvAsPxZr8D
5TtegSamThP1b69JMBqGAVhAPjU+acLmQvS++R7kl0YziYlkWidyS13NF8ppmaL1258DaDKP7yh7
Vy9mbMHyvMPa735WSrCxk22ApYsX+Mc2fzLJaiN2cXYj057wXk4dht17bhXOxAT7jD9RG7WGBmyB
ADoapHWr0AnoaPJcSuOsqupP636sewyZTmqoB3bpNt0Sfpbw5UJsrNwa1QxooAcvtEEkbU/aaXMN
dsXd968VDBd472kAys+UPfW2CbwezkeqVaNal7ygZCjl3jYkld4LWp/KZxqIkBVuY1G45e3COqqo
7kwxOCucdLjYr1gKDRUhvcM7UgUfNZSeCr1ZtnajFwKVOWUx8AIX3O1gTB+SYzLVepqQulllKsC7
7Ve3BzfcBMs/zXq0D26vW2YZ6w2QGMrFg0WkYKiSDDjBiGAB+MtGS0Xuy9MdH5ood3dYeDUABuVg
97YWv4J8uj3CPEwBxlUCxQ5MN/dpaU4RABLPLHvBEuRZZDfxgyfdLjzG4FId2Mme3pqlQacwqp8Q
KRjCCvW5b/cZtddxAi12c93OXgEASnMbAPSGuoKIYumptGiVs6pVDbA7+D34Oov4BaNF36uOm3HB
H9eqO6XKq5PT1PdZWZEW0GnD0z6V6Mmbr2fZ339AhdBaPhFoa9uzJaD7KQ2B9GQei3mYu06u7XeI
lXScFFsyzVvaivcBMJQ1lv1h2mv32iNoVO3ZinO+/AHaNozI3GQTaGRvJAXE44gUUYaEVahObiCf
HEoJTSuOZoU4Jrnp7Tc3AeauqaLXVvGmRcRhT9mEOkIup2nNg2mmGhAiOEMqLJjp7uq0naJgsZWg
oM8MuHHKynp+sAFH3/x59NFS0KrWVNpHK6Z93mwRx9lllCP+COAG9KVh+gg1RNNaNFiwxFcfNNIv
IoPJuKnqsLgvhVmzNr8rZThNhiofyk1PjIX2c6P6O7G+WkG3HMldn8TXphgp6zUqY8AHgmJWfR+s
FCMPXLtkRqQhKBbCMNLxICSgeJAD5dWHeAdj8gJymmoIpEFPsV7oSL0sxvmmI3IK0+cqA6EfyFOO
Zuoc7BlswPx0a0XxsWKW0CMNtIKX3yMTqWW74yOEInfWpoDfDQr/wA6hFV0z1jyRAdMm0jUotONH
XYuFh7gKUtWmqb1pfZu4Do+IuyGDAWbmOZodOzte7HcsP1b25W+VfrWtZk5g5EiwA0o0XD38nY9E
rObyIEd+c/uiC4nk3GNyafvv7GJKNT39bJXU0opd9gKP8WdK3oqCDuKI79AmumSRFZtds8Iaxz3K
jjszqF1alWsZtSfwFHq/I87IGcHztHPts3a92lToEMA/6tCqI5z3FK6ne1hQ0jbynk1kJODuI29U
oXXa1qSmoHiecUsflBhtql5AKgIaGM8RbpBO8oSivchNuH2GsmB5zjR7+fnUv9eHA+XUmlpCzjNQ
fKmk5cE++lEjOXU9mgolRzEumkscTqjO+9xtqHMDfHHGZjkkEJoKWeXHBj/saDd8GyGH4BAuMPVx
ij/u1syRLqLC7T39LRZIkmtm2Dp82UvATmgMQmgO53Q5TVSKUz3+uhqcxg8xbAP44xebJIzfsU7P
PY+zOft76UQKtBv6/OnijzStyMjR+qs26VZqx8qxnIC338soT2vmF4ew3YtrqMbGLw92exskaTg7
nJU2N5MaymUn+Ykt+8+UWkutSrIJjSkJu5aRs3jpXg9m7G+XhB+1mCHZ039FfAl1xpXlNI6bEEg7
VqXb+nTb8Cjm0hsrlkDSy1JYUMDvW5/HpPjDk9+tHAjmUE/6zFITX5d101Be4WlWhYceTMvHqZQC
+6V1GHYTwnuzPoPUMOti+uyffCCX/VDmuuto+zAtRqcsTXUGLek87eJkg2sGQ9fYL+j/Bs4fNac2
3WRBYR0iZI9AAq0C6sBDsdgdPSchZ4DKQ1p3D/2UrrIyfZjhDvnu4Zl4bhUIIqm2nY2swEZQ+Bom
ycbDKFaezpEhEs7Sd4exnBuH1aE84NRY0W4fY5uI4t14wOoBhQrBrWp1ug87ABCz5g20X4XTR6a0
T+W0KzgpWen2rA5FMnLDqc0x9ewyLy7KUw34xka7d9S18K89Qc7cHJ371FRQZORa9kQtXRxZ7C0+
HNPpR+g/1F7aFU7knO17ROPnqLJ+vsnixDr8I55jzsBnO2b+zrNEs6VVTHxagFicTGe82wlZcqV5
gGdkdU0+DcY8K00nGwnqnXVl2hHCvzu94ADP377QRF1nuhRK8fHWwtF88yrci5FcJGAL+JpDT+qP
RGn/jEUNw/HT/EMxKMSiGgrP9kQb1+FQ3t5Bc1qGAdA+beGAAtwIWdLVYxPfo5VcAApdnP5sgYMR
jIli0zEXkjNecP/YGVK/zvaCKKcBKCNVaFlOKEww6W15KWdIKpUE2QTT9qh30456xNodYqfoBDOy
XPk5voCSelW1UY+C+1i9l0f6RHTRcyZjJfkwYWgQTu9sEyJbxo9E0VD2brIVDjCgybTnpWOmogLV
qiH1jpZxuMU6ohUd2KXLfsqfbDDh0/z8P4onbz3Z5wcRg3O/x0T8U44ulGf/OCFBdNf+mNM8MZ4X
wLi2FVTfAL2Ag+m8yRWCGhMJYXJvUk847chrUU/kf+AiGx3NqqS1Os+dxYWD12fT1vMMvNNYDZew
aetf13AWkbjIaDgrIICUbTc1fnjIvcn5JdpELiTevEbQW3uhnFiLKawiwCqYKGPkX55OpdeMoGF6
4Nse6uLKGI8HR1nbF0mEeBzWiOPEvlFXibM3isTILBYpvMa+JUS1Dm/tcifYgTF6EEe8zhaFtvjR
AGEyNDbaExPfIJjwNTxUnvafVq7WNxnOpR0612/ZJSQbt5F2j/syeprzz8OVtwx27mGtqSSqzE83
YFUh8+ndIkZfHxpBOOYYwOTKfUzWETdNl3bwDbXy2His8jB/fiKHnGtW++EnYO8xwvHDmaxD24+X
Ms8UopPLJaN7pvyJRy8lmrTIEJNsTOLD+KhkBPToxt5sF8gvY2EicVYpgmlA/rKiv4rc7cnw5voz
xjrtp/ElR9Ybf1f/R/BdYqXq75QlNxDeehodBxqpbKkuj2IlokxMe6kjJMTc6fbgdl7eAh1U2b77
NMjsrE3DeYheImqjAZAe/omJAicbM61CCHU2hsSzIx9uqm8AJ2sCOSqkxNk7HR/B6fG78GVJLmIW
4zxh6Lvzg0DcxH9jacaYRs3MW5LFlbIuw5rUhqHAggFEd1Z4Td6DAC5wnXVX7HOy54n+wd2R2+6A
qi6T9F2Jg1zKpIuLhDGNoDWNfCJp51l/pFYtVRt3DdiuOYw0wlQLaJymWw7+4AXNwy93bI6CKiwN
RQeR9o6r+KLmWfupn4Zbz8BesnTIOLKkKoM++RkvE3TZq+DTQc91rZ2+nheKb2J8tbbnmzua8KBe
c1o1buKQU/kJv4TbHNDNSfW3b0ZHvKmk2KjUeH43xVSqvvfDQvKNeRJKhupsWA2ZdUFjg/nKC7t3
vVVqaSCFjbJEtD1Tv2Fy91qESSSjlSNHmWaBZmtq/mOz270fnUmRkqqNhg13uk92yg/PmC8lmQA4
PLuHZvMMriXNWqmIgDNOUevwHZ1fS+RpoCPmi+7cPU6NCnkl5oyBtD/6HUscKSB2aROpHl5AqhKF
ZVOd93pEex+9vfqYO1EeAimBFpMIgur7vY3OT9DpfIHsw32rG06knT84KsxCGO1JK6VvtSIElOYj
bK/IO39s0YtkFruQs1aVE8rZcIG9p4XJ3o9k8bHXnEokQYQoVLdrl20d+wj3M2U3QUs7DWgEsYB+
Pqqw2SSC3MBMAuPq9krMusO2KUtHkxNOjiHzBARRIVNWChWZfeAEIjc65XFcSxVYlEo9NxyHNGRC
tZO4tAGe5hh6xheaBxz/fgZ8vEbfPsZ/lT3hcl09DX7OXtolZHhKg3Spj143rkzLiu0qTDBE1e0p
TcF5wTqE31Zwszuc0krcRrLHPRnhZXy95ASF5hD5WTqJdINlA1xmUebRJxfMQLsVekVbNUQdw3N1
Wpm1fWo5Rv7/QVBTUESsJLxZUmTVTI/MC7ch5q0tH65IwifAZcrdtWPj5y3dYu6Uts4IGNpJb0q+
kNwsYyum/cV12m74pB71+Jeb9rF933yOjpNxUHxOmbNKGJt1LH7vDGQcEoCs4ibMPiEcHaqwaDEr
UP6pBury7JQJpdeiCzhA+qyVAoB+p7yPlGACGoE2PWTt9SLdf8oLeS4wnJydYf2rgUjvXtLospzg
3mS0qKx5SgnaY1dokRgp+WjLUb0p7dq2VFeCcxsLxsPl4i3NUF+lUrJORdcL3Sn9jP+N1fMmbDvE
focZb2XwTGjUyLrg7rHBypmL0tlYSeVc2KzMRPmNnSuHKEjQCOQWXNhD0MZawBiMm+QldVfKobaI
P60//U5uDNgGNm7BYP+ne+hWI+O5ejtEhzkFSJ5GCtf4Xb2Il06pzlnljjXIWOtD4D22tB8cgo+I
5RkxVFrukBJ49mUFW0wxVlhlWVi1MkBjOuyKZvnYGu17PVDDFagVF9wbnzS8ciOjOEesjR0Lv7ym
4Nly+7U9WoU8MRw1CfSsn9cca3s8cTW3jm3QBzuEWUCm80ftgXdRSijqUY19u2v3Fz7/lHIoi9v1
lUUcsZwTywzZX38i60IKhel/iYOxRseER61c1eAWA7msLKXXCXLa0xft7W7U6uSqA9Kd16SbJC10
Ihu+W3Z0Y8LeTwe0MYzLFeInmhna+bIK/Z34dGvFQc0C/tHOx/WZJbHobITYcFc7BI8V+5C6PcUp
wuDj6SZ6MYA71Toc/xyKOwK++WgsO8W4tPOFH0qgjMveb2TayHVVKCnSaudZJM3vnc1SVKPvAoMl
1BK3F+G+aAfddpxZTA7hA9VSDcIYaTmIwoedNlzB5WDO3w9tnYFu8CKbQxJ9Qw5va+5xzhgaK+2S
crv6bREKDtgP7Zl/1C3zHQnYwQycTHMiLum2HjuNJQ7IrL94ZIa4VEgM+QlI32yeogopav80KSyr
iFPxkFvbqa7wwLglLkK3h1EBQY75cDesvGtKtnUJKTxMkAvJc9PrMX+7Ab5aDAmT4/+vqFX/LR2R
VW8b9wf1B0FCM/GD0ivtKoDivOds7L2QDTJrA7bD7Vg4YQyhfIwuh5QuiQW0sm+Q4blPEGGrcmg+
R/xEnoakIejKE6NK7jcahGX1hVt5MVSFjzkVbe5PGW+ouVUHHE40hjLACWNB7iizk+T43wsBKwbp
dNN60WlIQLt2rNnbXkD5Keg0JT3MR9vP7+xtr31OQsz+PRCzvKfaBXAdFssQ6E1vuXfoGCnXOueT
spVgkhq/FJnhew05tDzJqubb/FTTSUviBPtq9v430GZy+ZU1vP5z96vIHAFuoEP8DqMpKh4L5HAx
fD0n1fYXcmTrB3ThcLx+92+gg5lIk+FdcsUPOtxZY/KTxqvKzzYd6cNMXBQNop58Q6owe8j93VJg
hkgj2oa/Xxrz6TidpKkbLJEXeTjo3W1ZCPTuPyMvrNGKCEaAWkkGkOvL23KJqTWfRmCyLCLd3v0M
J3c93NF26+Iw0c2mQk/Pycn56jeaYjWXO5T4aPQgF/MbwySfNdyUIi3/Tfn15yM3tu+/uj17vW3D
cUEy9ZRVcro0bq82hcQPBYDw0Aj4QNXZ6bx8od2x8zZkxTq/tIJ0oCKt5AKVsljhV5Qcko5PwlJy
ZoCggqpW06YVCYMFaDxzldrSWBtw2nfQEaQJb7DRpAP/POZ917NcsCMUZSsCH3kArY8Gr8DZiIGf
Sy7pKAXnhzRy4d8cj5hr9le2Ni/ZL5dU6PQ/4m32O07eP26KFi4BQPpA2lkf7u5UXBI0jzaRS4b8
w4Q0aVDzxbii8Sfbf7h4z0/ffiWtdULvxgr06Bv1edCaLPQoNA2aQJz0LokheY+jfEtZiXeoQA2F
nizM6MFIkRcA/pIg7KKr0aa5ZqiIHyizf437dFNndJXMc/2KmS6LzPJggY2SJJQm201DuWca91MC
cA1So7YW67juZcj9wlkgYfbMnRoW9fY78NFccUYc1039avXuEAf98IfSmcAEICUwXraEcqbHJmkv
7jYmhVUCaYreHoTDhG5b0gIwSEeH5BqC4dhA0Gx6u1XgqCCy4WDpJGQfEAk1nMPuls7Yn68lGL1K
Xfls9NQBwQ9fOsWOh3ZscW13DSskh1gok2lUwwv0MZs/cROGfoBl/GRlmQaWhBBFaTRxosCoXCCO
MqRxplxthCWYVeDs9EwnyRf4PXO4I3S6+jb3ywm+cz1rHrBOIxLK/7FKdMcefqok54xiDpsYBTKA
LcbQygHRwJPsFoq2ZL/XENM9ghMyOqXBcPQro6TX1Z6EeIOi69XLapUnWczM48Ju5M73GQkhWS+R
L8ikExKY1p9Cy4arbKfKTsb0c2SHXAk75oj5uAjLR9uis9wiauqdZBFL8iEwRQO6+v75OnrolLcZ
tMZAMPJnRI1KDYUYOE5jFUClc8oxdrpgPExqcY76iTyEabrBcapJFEmN1ng9dz0+8WBLJiOYFG/F
AdNZZ6VrVQcJYynK3Pcaa56k8kB59NT3+Z6jVzB7rhLCUmP7fEGjqMTLRsu++zPPP2Y3fyrGwXz7
Ez4syEqyexjJO0qHjE/3MGqSZrY35KBiX2NwWVxcwTx8KGizcyklqk3kB6cC7IXmdo2f7sshu74w
QXzREaGEyHg2lsIE94ro+btK23tSCY5JLF+cQnjdDp+r6GnDymJvScxTOxvHY1p+IBg36IkgGQ9M
R+41pAta82UAlqvgLuvMowm8Wf+b1/uWKKPNXmWJZ6qnCAk6/iubTc734tLWV3KgAniMX85/y1bk
ySJYH3TPNf0+3M8TfR7jQCuF1Ce5cpXo7LwDxu3ZDiDyJZYO8jtxg5N3zn1c7i8W0QehERyaxHNH
O02O8zQklVfgPXMX6VZfyQ9l+l1yYrbufRkOfUgXNwCF+Co4ZoM8514+yIbJMKJz1fHsy4Kazdds
CxzZhOJA9KFTSK3+zV7g4Ablv84RgR+56O2qdFKgnGpv4GGfNULh8KtS7Ex3hbTacJVABLIgfo52
PLGQk+8W9grSk7/vnkXLjI0ip9vH+gZKZA3l9xL0MfO/rKhpCXNf757NdphvMvEsBv2JaUJYFpSY
6XiFFLA/Ql6jGc6Hpq6GLDjDNsxigKSKXQDhHDVOI5zoSOe+0ZbTay40AocjmABvfwuqv3TAt4qu
oVvtMU4/qgCCNx6WQgRV/xsGDoJnws4K7jFkI5Dro9sENmdI32h3t5LvGsfWWVBJcP3fiIkrAdbK
AD3hyKPpSmWzESMcpYvCPwErTxPPt+VeHEQVuVpvIauGqZGoKLA7BrTeCM5eDxuSc+qBL9+QdMFl
HfTrTvbl+ml4l7mVNtZJFU1u2gpg4jSnOqE+3wFOB5iVhQQxOKI1rPKdPUulGsRExHT+6ufhH9Ky
ke/Rc2PA/HBZQhG8L/ac7Zul7WfmLFyLioPtDGbMYvwWyIHKvJfTqPDHaPqraWfeZEOUggjPwkTt
VUotRgymMVGrmcCNeTiEvJJxuvQZjvsxQiH9iVT4fBACG3iesVDfgiBgR9xX0IXH2q2MTx8YcWbt
KPKDjjxaTw1pcvaVar+JZwHW85jDert0qauaZ9FgVWV82oFj/5s/lXpZeDBlMLfQjUxlpsENlcdp
1E/figIu/MhSLGFBGJopHUi/Dpu18JusNNIMJ1FYPX+qcWRGXxWvUDRzFAdabMN1BPSV8vLaiEHb
KjOUensXxRoEm5P+3+KQQMpyWnn2B+y+qjDmS2NFUsBUqNNplRfF6RL9BCJCMNvKgLzBVkF24uEi
lqWVkfB+37DFk4QOU1/zD8Uaz1aCmnRQsnA7T1wd04JQIBXpRi434rw5JXZJXxFRy0zz1FwPrdml
RG5HQ66v/i+IEY/pp+7oHq7LtMxeN4ThfEZUgNoj4IXXZ+lbB0y1uRcHY5G/N726sDXEFVOB6N5H
MrAubh0zXfhNi61NtPxAAR/44wPueQ+KGFWQzqemc8+YnOwTxIYoSBaPQr6KMNHx+JDyUmV5uSKZ
+KUGZCLIk5gQHb86spKNRvrBpd5n23QWUx+l4694jAEJwG+WuMrkR1IqTe58ulAZ4fOQwrDw6phD
eEeI8Yke5Zc0vFXE5XfaU3QLhwWqRNH5unOs88Um5BJjg376VE4Z8EO3r/JwL6w7512g/sEy1+Ym
bqWBQaXHPjLyzvkPnJUwlXsAZQbL7I0j/3qVX7YIoXZdBeNQrzku0mr4jbTZQaMw11tqQ90pXkUn
SRBQ4F6lCyIyk7YjxW0wxxeolStaOh0RMHOFgvIc3J3q05oOMdoiesCLw3mAhzRmihjkG3AgCrt4
tWsBeZ17+A0CEFua5GK+Z9DWILbxGcIOKnWrbe5KDthUzfyrzUxq0IRkfXs2M/3ZdWwEUDBcO0uE
MPQec/rG4O2FLp3Zt2a0kensUrmP6S6Raq+iDgkHRJ2KJ9tpoUQK27TeuQHS9r7axo5ml/0T9WlM
D+ItBRSPXlSBmI0LmcAykUBHfinUDj2bl9wiKuJkgCvpEqqJf848w5u2jjyBxvLBVDrnDaK1kn01
QHQq0PFjmtoA3afLbbr/GIvVrjGyX9moWMy5+znFFcbbvYWWeZG5dFA56742A+5pJhc9TF2ZIDKc
qKRyzwcxAA23Z98qdyzd5OrF2oZA80jr7tD1t7BV0H1Mvkb+ogabHR6Ihhl8Tf4QsPtGtD/HEum3
Cm7/Sf6BWZX1EIMwQFX71YbuEL4GoNKTAzpYeXrSNbli5A9wzzhKzDMPJZiS5vdDbAkuhfiaLnb0
HxV8AiDUiLqp5YbvuKY02I5OCMuLBc/REqW8xqPJQALGIl/OCbza3CRwBTToLSfBAioOdghGTKcU
dGHEZQeCxaYTSwhSpnYXpZWF/sEfvEH+Cmm6jskNSXTunNDlODqo5UT3DFX/rJ0kDoggzszKbM6l
0oP0oMPiy4zslwBZqV2jbDqc+S9txGDh8636goetyqssNI3uSEbjlYJvJp0rSDotcJP1RHVg/S9K
EBYsd8dndy1LNfJaEG37ld9Efd1iLF6pdC9zA8HEtYCZCdMgRQIjYsPPQkk/p89AH7ryEmon9bX0
gd7wZO1ykD/M4gibfs3D+8x0bXN20+0wtZhsZ5qYNJ0vTvxDE+GC70xz6N/DKyy9h/RRXYznJAE9
JcitUZYa5Y63ehAV7ckgpw85ULvg5p4aqBt8k54q6OwKGQrdyHuSQ7uKV3dLHW/FegE3klExi+ST
2NSk730VJhGiaJZ3xLbyh9VXjUr425nuUwEjubhtAadnVv/zhrxegbYwQIzJtYQPJ+mkBSppIZDx
lNzjdFfpYrHt6zrOxm7nwcqFtZSL7pa5DQQY2QeZfbC9bHgSeLVBF4hA9GKFNrUJCfF3QEmDvFSk
RKTijfuSQwRDJ62mKZpuYMV2x9MwYfPOLZNCjpwjcQ/CjzLRXYhSsnV+ZGjWGbb5WAH0EfXwOvtJ
473OsoBu90NAyrK3mhZfNgdnkeLTJVqKI65p0q3Vo1IbIMI6c3oMPji6bJjYVvmN9tDt692RW6x2
M5qaFDwf/55oAlsFFyRAcpvS4W6oDp19HseiD1D2yMcyIgLdGr7nqrHEz5Mkf75FdYb8+JNyaWgR
FjRnu1cwP5JJPvxxBK1To3oBEyVr4dk5zWDo2WIO6Pq7RvDM5AY3imXtI8g1Wg2+h9H9uhgkKMRx
0IhTwNmEh7fFydlX2JhghVoKopBdwYy7TL1HUpaUo9glKsAS51OXirtMEDoEq3OHDOKixdNUyTtS
nO7SOJZaoU8BSBBcHohMKKUSdtRWaM/DpM+RCabERjGYsHPGJVzkbYOby+BiYLclojE9RdjiOxh8
XfcvwxTl138Fq4eX0KNVyRMD3UOtp1lM15z4WectAsD33cqUARIg+C1sdtQXhGsocb/NvT76fwHt
G1hvTVq2UovPOXKCCcDbjDLwTpGsWb/pj72mKZHFFToBTLK8FnIEMlkWIi1J0Ab6kXMbD9wnzd6F
jsUhPEaJA1ylDAJHSDgwRNtPeCvQuu2JC/7YUhxOjB5RWF7YOHuojfdYPYsPbDCrrqcU18cJL2nL
tva5E8ORQgvoUU4Tid0yNP0A9kbAQgVFEmMDjciz1kgf9DQDXPCDT0Ar4DTtAL2XbKVLoxvrWYqf
N8qOGjsUf71ZAL1nt5wCP8h924PB+cdUoFB4Wxc1sa241lA3BrLwyh6TqabaGSYAvbU/Vy7Mfpbe
873J67gLdW5MjQAfbf5tpfjXUUcxhOYz3vTe4Qqh7cvat/0cCUTfsCWiuyyxecd8qBdQRNEuaJBC
GcR7Po93VJrTxh42fSd2uzZZcKqmmkDE3Yqi/8Wy1FJOdZjZIZatBSBzAjnla3TgvPqESeDfbcqA
UzyzamjZRMT7hIPZnigTgiYlqqck/NXIYMI7GlwkERYbvlOGlR6Xnnu9LJfOPhLAwqOjzKbQi042
lzP8Mzf1c29I6sB1QmjkV13M16tP1xv7AE+Wca2ua99oXDQD1kvfNtc1EQpG2I06PT9bjhWuYRXy
p3dzXsRD03P7spiwgD3ZdctXSVbRP37TgAZCtMMfg40DUlbjb2txnIO1xCoYwrNdX7o3j43TACFi
LEPNcfSde/h7qaV/v1L5wlH6tF3PjlUWJWh2HKEsz7EYWxh3zvAbzmUw9B/CA2UDoOe5TiLxBYET
bIp+i8mF3uoeABVQg1ipi6i8XoqOp6kTgT3N3Aji8kFOzioqxzYABjo2Oz1l3xXE3FfEDycD1gVn
SGo05KVylvW/AyytwgUb0l11/ja9h1udgNwAqDef0mFfsrrlON8oev0Zj68apdGjn+wLkFHBRWsN
9C1kmjuvBJcIEtrQ6kbGTsL8696864O/OjS/A1t1AoZs82Jv+YTrzdTip7qj5LlF7K1TxbWF9cDX
9wWw0YgsTBnjR3X2iouPolieFYUngH4GX6nR/eTeGAztC9GcCbE0xT8pIRsgs3Qu+1+iIagRs6n9
+o1nkGwQtCw4cNgMY2ODtKCnwiUR/I4bJFCYhDj7s8uwlZgHr+fK1ZCDa5PdfKjNAu6m8YnGqcmv
XYmOXALzphbyMPcNxsToySadWT1MWSdEK8ySGNuE3KBq6EQeI266VW/NP5SjxhChztAzP7sMrYC4
KAnIrt4vwGFGFDxyq6QvVY9tZbnxufvT+gty4vpatUFPsSSX+Y3qVurKvXxtLWizSvc9UdbpROjo
IgnaLbFKLlYpDJ7nbd/dJmOrb5TxBgACjh5PdBnEl7ra1CrOsxmWGRuz/GTh1SDgXOcN1+Kd/erD
SL5XWzmXQN9qKMYt19lrxfjRXgx3/33UImntelEqt6KlewfBiDarLjsrjcGkT59Mx6Yk1ALHlJdX
j10YW42r/Q81u3dofEa9oDpf0Q2hOgmgkJzs+fmQLI1UIvfq6kgVKIaVM3DaSqVBLj7K7z9dN9mh
uDMlhpZhIMukght9oRTJCHdWFw7kaJbKzjTZhqeY6MFTJvNqiG90GGB7XbqVLo16h3sywZzv9yY7
GEF+sIseDGYqqcGyQGfqrSGnznih2cvKTRrxcih8Ex9pw0M8QZEzbdNg2Qlf2I+pHFmej0vA5kri
rksEndJgQF7XLz8p8PlKW3SZwSYDws8293tytvrGXj8X36PilXHss1uG8B696M/MqSVtA+O5uPp2
rTJrufBtF1wCy+JrGSAdC9dAHqnRLrHYtIDuNyCrlkpyTvGcu/gc6jN47Hg2aX929/YHuE6YXFVr
FN7b+VXSCX2emLZ6HctkqMdItPm9BUMcihfxwHPgTPpbSSV11TFi4MZBEJy0jf0PHbYAlZigfmyl
NSbZpWr0ZUjLFqAd8lMH1j1H7KXNi7HKd6NkuYtvHsPiKjW7nwtMIqmXuKXvj5PyXJBjPOXPZVnX
fgC4yCKLX7p401OtXm/YksO96V6l3n+hfqhAWt6axELUsSTQ5Z/OPDGD6An0COs0LKA5eULEgK+l
rujk7WO2nWcMGQ9d7Ce3Tu14xgLme9iDmdKLd6WUlv2VmnotXL/QqyR2vB7pmw/luzh8jGm3ppIc
pWckeCLn7Wxii6frdlVzoFRnv2eHjYFQtbtfpHTrrFVN96qJLVZ8VCM8o+J4jMgis6+NWQP8nHTS
tp2aToWp21Cc0kK9aydrb+9b0CCxL184/hzBrsHoo/gRr1m0v+rA4/IL4VRhzk/JcHmXeLApk4jO
HYcX0Gnu4BvMZa5nY4mb+pJhfqggssLhsTJ/zGaMCPzrKkV2shcNWQ0iHRvTthqOl5X1csYkMsT/
UA91bnNRSuMyI6zEpJmsy/1jUUXCwalHt/8IfcLxgbWSc5QkyD0arssBxaELVuM2AABPlg4l6TPV
ZbGkWYqhDcFTwMiXw3uQFhcQOnTOA2Tc5HSS6XhAKKx1LGscYhykzSYk3wyz5wywZlHWN4AiIFOf
63LRGQMLyB45OA2331G1y87F69YfVfuSUkGkyPQiZERy2ntsZMDs1Z09WJenUireV4LvU7DDui4v
go6rQG52kBakK6+PRXdFJ62A8pEEfx7ZzgtXDqWNVzaNMdoQQxtvB5muR2+v5cYKozWqzh97Gilb
69C7kOc8iuYCWtHHA0YionAux9ukVmhLhdMIt+zZoc0RvQpo2Uw/HWBoxU7RJFOebqOYYqKCtzH2
16UQphJWGS8dEMo5HJFuOdpNOI7Rs1s1F1wacjOQxzq85zhI/zC/+/5c6DP3CxeJjbPkrsSvaKv1
YmJBL6OcpLZI2AeAqQyCQP+R0o4ImRXi2aIRdbXhbM0AOEly4Cr8KioyKYfupHc1oqvYttvTugcp
l3fAvnOS5/IOenmqKng8azi3yiUzkvMckaclVgv6UBbAkGjtli0C+6+6Z+tQpwAwRl+2mGp8+pUS
dBf1WPsh/b/3tPZYi+VJo0GTHwGNsNWj3u1hrZpUcAJNN9/NLJ4yF0kKqJxZ4BOE2bFC0oPNC+vG
H1LtLsiTs/kmV2rgRQTNxTTVcmMqKCLrnRTjUNkaXeefl6kNbScQkKmc7nKDfTc1qj8//p8wp/kb
hl6mdGg8eJ3c1RG8pe+tVEMUFpgkL/PXUsIjHsrsAKGO1CxbVkTtIL+OTD31J6272DbOxTnS6mar
xYVWBwxFMURLKx4+O6TInKg0f4i1md8BADkb3w+zDlUJUSkync1dzXQItEnNTTMIVSB6hmvhcvh8
AdE6hQ580/mk3eRYmZs7mEiZNrjF5bk/uJE7MQNhonN/DAiRI62grI9s6MNvUarqg8OEuDp0LQEx
Rw62VwB+WdhYvaJPAnxwGCT4Acfj3lkgfBVwde3BL/p5D9hsQU1TjQiLHIW9KQY1aIubv5jnuiHs
IXnh5FuHMO6uyw1vMQheK7WBdjJ6TYPESwqqFfqcDMtukKBZvUgnwZwr9Ay1KBqq20dcTHTmqXoE
X+XAThGSIEe5O7ZIcpGf6HVYT3bCuHNYh0FsyLkT0df6l9vqDka3YLoEPT6iEJFgI+hsPjmHnYdn
dSFsmutydzwrA3u52ElUOQ2PjiD5gBcSy5g4mRLlfCW5b8K7uwnyDkZVho92Qj0PDz166CvhU/Ar
9qaJVJqM7jTOGaUVLSZl/CMf6/YV44PcwDnPYa2aszbDD1PKkMAmA+obdblYgAZ0QgHi1Dr3LhaY
BkyI3smBxzjjZNCkf0lAMeimBbFUFcPFDuYZggTw9cOf+395toX3TaDV/JTmAEmtnv94vpFlnpTR
lX1MC8aUZdfI5gnkkbVhB1ShqEkX2OWaU4S0CbZGsYp2PzeB3BY1CteS06B16eWnM3+tiBRlAl5r
zE7te/Ui4ZF46IraxVhxEvkg0yA2dtrj10O6nyKRuN/0TI0eAdU0VV+0xteTYxTUtIVKNLevICEi
B6Jbbi1EIxSkFs74fLm+XoTWhDchSp1JW+VerjtXkc0iH8WScP8ra9PKdzIg2iTH/qW5UVoUc5ks
U+6QY0sLGJUn/JXl7e1i27xz4jEFwA/Eep34qIgAgF5vgSCQnPijbGeVgp+WLVFVgvKO257ZAUf3
ceX/AN9R5R5yeVHd14iiN6KWP3NjXqyBFhop8kHXc1T5TrEYnf0MRTxL2ocSrOxAKKphPR0EpdmF
FHT6SBUkAcy/ZfNnq8svSFGaB0Koc01iHQpDTYmP+7ecLljwp0qLO4r3bRYIf7ZtxZVLRYVcWs8K
Fb7S0KO1wcJSAOpEeBv6QxtEIda5ikgio+BZh+96hEH2JVhlpVlOGbSE2luaAnreXTBiVAhNsKeH
dJ6psz0bNeb1C0rabJIf0pyi89WyzA20F/CMM6ffzBc+SFjc4IjQt7dcTEP8tVLwpyROTNDD4BJb
GAk4Uxhcw83Zfe/FVXhD96NI1Q+m4koUdQ6P14a2yAO2xsSGXINIukLyBH51NFs2PJ/01P9v3DRz
tXsFxP7bZE4HHMS45xX1O47StvpUUvKb5xQn6QK+gpl8aneOA0ZsFJvrx8oyW9A7Ha9QzPn5dWCS
3EMVErv2aShvwPCrPtstZAs5pMmakY8nAmcdmy4KPzrsn+pzj31tYce0NFUbXyu+AuySLAVbh5Pd
9G2R1oVroZrrIwmp9NAx+aJHUFCCv//2IS7GY6IoWSNVJtaAW4tveqg98AH1leLzaT5QmlluWFNr
Ak8qBgnts9+dnCSQIF1PktVoNgBL3AGjxVlr3AtjkUb76HYrGufxahQhsAAD3AykuLbRsZCBSdfT
hRhrKKz4FFdzx4BlNacPUlF1rxhTWBLVciBwWZl8efJ6X5CGe3a7eqZuP/8i6sx9K1tU+jbUnbFL
OQSnOmulpsZRfVkG3GZsdIX02REoy3rxlouyiMiuZKxZDu+yoxf80yuz3S/aHJ6+iyYGIJtTGdeh
tbf3N6DOSilA8q1TNkbcnt9amaK+Ry//c9duuVHKX9Y1uCKJ/2acME/QoNHWqOCrJKbx3Yk/nJeY
xGtaYQh3z7Hkwpl6IUGvftj95ulHzogQk2S08wIX606ITqGEUltMlUrBgRzJCmbOHuWgLfo0bXuE
sX4pk8EiAZojWqw+UN7EWdgWcYBv3Jxfd0pI9ABPbXD0TPUW9WVYFFF2w3cgtLXgUr9v5Htuwctd
N5BUK2pE0yHtYpgqO5xckwt3wOKZzu8LuO277uzYsnBIZQbKxSvRbm693HPq9SNqVUDa7kwy1hdy
AvupQRSCURrKtgP05y8DFMhuWlCCER3BXrsBuPqhN8eRz6ud9OHMu7qiCh4Ycjc5U/R9x1V2Y4gU
ay6cwUJfWow7si3FAp4zfHLnvorqHqzaGOWLUrE57tRXPzyRVwxr3ATO0A6pwjRFUqJ6Ez2x58XI
iLcQKHGuTYd7Z8wF4DPyUQG81ZutQbr0djy8OW/S/HFJHXSNsDle+qu4v+37KZkLl+SeLzV1Yn8r
3d9xsrF8aU6EOSP5D4fcp5SQikmQVKVZt6uzCILcuqfmpXEgyRcKHi1qMAkR6LYvcCbMCOe/ALME
vXgafBuzpAhnUzYdyGXpjzpLGfpZm0L/wm81hHmhnGc2Dt9M+NUpQpzDtrVflh/ketMlxKiKH99e
XiC74DluGcwmEowbJfXP0qW685YKGqaDJfGIUJX9It9ox9Fw1w6kfqUc3HPirj9+vCt1ygNaAtEd
pb2yv6QDBolorLZkU4aTKaqA8gI1IHuC+B2yDs1q6Z+hEtsdfKcLZ6nuOZPwEE0hdYbeTeUdyboA
gWhgpWBHpWD1Srm8xmWzk49IJkapBmyDOVNBRd8nxk+ZVXulpDIZ87rHwCrxDLHFKovYTAIMykL8
gFmHU/EPHLA8biOllf4vHkips+IYS1aIfa3+/8jkGFBlksenVZ7D1gxeUQ0c3Vj+hSe+1gBvRFAV
YxIEkh7sRSJNrAbW6GPO8FXobHL4PdNLQmGhAfXAyLSNXjyBXcvPa16kBNcP5sYqcd59Op5T/SFY
Y+CB5Q2IA43Mb5wZwnj3p4L53NEgZF15FJZE+cs/c0OIz4ARhgzJTKQSjkhzP+n3iRmnetRME2Im
9uJOSRcuw7hVREGp0DxZaLmxo2QQJlDEw1XEHeL/kgWN52OPwT06YDCVPmLIRwqt1PC5WHNIavrA
ERp5fplwLG+iuvSznfiTZuUh+pXDsX/9+G91yIUHdiQ21my0YAqMKLaesue8DKJ772zeUvLoHCmc
EL8VhzLJOlhfjDp/SLRDmJ/zlOd2FmtP55TyPbpDgKGSTbehsmlB8XY+1OtzoxAMh7dmk4YrhukD
/ifYSBFjGIl4kRERbAOUaL0BX6xhuxo/WSnoR588u3aQXYuFw9MrNs7qLiSCxtQntgUh69NIs8Rk
X/Qr3Vcsu5xtuz+zqeRhpIfUDYziDWgLz0J2cRBbnFZNSKbjKgxn5bQ1JRyZvOXpnxhDI0CsQXRm
74tgKh1hz87AZKOeyDXXl7tE+vWqRA6SSX4pD0EqmGvr5jmoT93qR8S8Z4X7yHK8UXx70Gz0FLDn
nALZPn90CpqQ/jM8/dibwBRkoD5w8ZDoX/fUVtAv+ArrAZgl2IF+yKvAtrKaPVQcYAlK1/NpGD6f
s3YtkUdUvkwseYc5inyRHX8cUiUbSEc2AGc8WadtkhYIM/GTDI5xykjF6ambBA07wYpwUSzsfsUA
NGjn2xuR3VNGVyw6LNlf2Js1w65KluK1BZBznsRWUP7Wi38BR56ACVbyJwH4clUKmCLLWV+unT1n
59n05i1z7yM3yDvBq6uSc2U348Hr81GcISCp6y5lzkOxc/IfUqUiPxT5tBhCFLSjqmVXdtADfh9K
D76zDR2X3ML5lOaWz1w2VnupX03a9Tn7F4k7mLDR9x/wcBq187gHCLjFXKmOEzzwdIDO+kJHBYNq
56qG5rChiS9c7ypCX92bHd5Ob+VWTK3QgJeP1YQEZhmCf8AATzEgXhezquzlh6zZ0U9E1QBoZY/y
dmSNn/V3JBKmLX42pB5TJgbHpBgGiwaUuKVI/4VJm4MbKAX3NGrncFtEhTsslJYMGuPLet3rKEis
fkgKtSxHH1OvAOi2FNTtgI3qdnT6E0SJc+Wt7EtTenU2KpHtyeY3yQiJdUPZYF3iCO9WeTKNF3lg
zDJX8IjIRlR9f4N86pgIW5Vb389XIr5Pd4QYPZxC8+RzAnGjrOmjKA0lHF+kwCa8l7SO1RIN8zh7
fe7zgVVkh/7hOyPh2SuuRph+hlcQIITFzGLEH+Ix38As69eG55g4RjQu+AjJnNajDyRKSzvJVFi4
lnwgoJfxR97oWsrKCqOg5XZSM8Wz78TcPNAs7kRRYir6M6r+3qsUOT5aq5xEqnWF8F4S5wFa8w44
BegpW84uvo2IXJfaLMikb5RAggNXsk6gk1ZVUYisS6bdXXpTwEdDcD6tuFAUzExuT42wTnTXEe0y
NS2kOxSCipz81iQ3H+G0zWiVgQDubqS760kFCUU6sLa3Tp9w9rZT8m7O+iMDzw0p+FWjpCLuZYLB
opIX2nKSAHGjBBgmdnQqf96R/fb47ldfWic/nJ33tRkbvLlIHhLCJ+JH11GXDMVayRZ3SC3x+ypu
k51W7Hb16vWHO7TkOSBE2s4+bgRbN73ftqSOFVyo1kX83BIxAlgDDTB66FmV25cPd4N67lLjUTAP
Bs00CZqblx9VN2jjZE5NMYgJf7LsT3T0IgvnXmv+7fQRuxwlObRp076p6LclcGXpYJuIInWsYBkJ
sNv1A+V/emoptnVLc1SbseNL7JkGMep9BuZ+I1Qk3C0JW5hiz/enOPUqacqiueWGR3TOFD4NLgS7
Gt3lJDU1QU2rY9wUBgRrX60jFsilGXO7/UoycdtATp+wb8+TFSK9TQaLr/nkSpJ/DEY/MCsV9O1n
atNBwdnLGYq89YIKLfm+v5b+I4H3+uMfmCbYsILtvia5J1AaaG7jefY41EgvQVNDanQYnsg2c2X7
8T0/zBGTdqgbogpasz0uhRPDLkbIN9qLPCMQohy1moM5ENGdNpZwuHuYVl1Gl8LLSYjIO4Fz8svY
ilIbMggednivD6ivB6cMWQASnLL9C7gsu0qPJNA0zInaIrNcSV7GDRRPpqjRrHCB3RJVHJIUJtRi
PiGWn5Lj84ZM/bcKoLfsrOaFohrqFqOt0pkUrJpaPg8Oo4kN3qhs6aB1AnPAwqqRKS3XGs2E3XuV
t2unkjAsYdYLPvZa2l9CQy4Fj34V6pkgv8DBg2+XiXZBKRcBp9koJVA+x18MgIbgzs75Be3q0r68
ssSrCYb2Mq35raYjl/Zccv+vP5Yz5i5alDtua50AcEA3HWl915T9ywYwrFIysaZncr28qzY0JeCy
qbAPuclRIz1bTT4S+xDUS6614FnxF0mhjbUK7xY66Sz7NZDmn2l85AJjLbAprLjYOf+TfFY7pXlv
TQ8G3LQbQLNzDHoLA1bncAF8R4DcunTJ2fRrbjNNMKKB+DdB8IyYhYT6TlUc3O8QlqPoOFkFsgRr
GxxNBWj87LjABm8JUD6ZUltfOhNhORyqcxFqE6GsnxL4BI8UxLCeWISc6B4wPxj/7cm8fm7VPZ3Y
q5cKdt0oYocJ6cZ5ygzQfraOp7j4Y6BKZNxZJxpE2wU23mYw/dU0+a4cSAVHzAJ7hAdFA5GZBEVM
/rM8N3+BNahfCLvu+juHdGIFzoO5+5My5V9oYx3cZQbEXCyMlt+ztUa9zuIPW18OZFqTLa+RRa6z
RhQ1kkrsuZC0igCbjqysu9avHx8l5j5vX1GI9VC4WfhFJAvmzbKXmH9ba/32uQYuMZrmgA6nOLaV
GXteHNR+ZxHG+5FvbyIXUXme25ohpDeu4g5gx/rmtJqpydnA88lN4X1j+MNAKm+BQ/Zsw8Iv45YD
bQH0pQngQH3pCugxcyI5Wh51x9h65yuk3Of/FMYglSq/IJpIioqd3S7Meey5K0KHOA11RFbqs/93
S6wFycwXLv7uerUy6dqbVJrta10Pu0BfuQS4zwGj0yElTn/1uF8kBzzmxblTkc9c3dxStiXTdAZC
ChzCjCjwQJp9SRmdG4bUUBp/qR4LU3juIl2sPJjp0lg/jRja3799suAJFc4QRNZ+DUpbCN0lRhcD
T77RIgUp7XaI4cZSzobeyLdmroinRcdtIJiTHTOKlwWgcI8xAeJqJea0fABTJti+PUExj7WdXeCH
KJ0D+bQ+IPClab21AEmkm0wpSmAnyQ7NVy6FtjbZ+le4tsylf7HRyenOB5PGfRR6DQc72fJFC4a7
NS6blNsdyDcIGbK4p4zwMFSjTM1I2Di2OSeENPYdd+A82gKvfb3ztPUGDPt2u+ta2CtgEKHqrExC
dOMSHXv25b1TQSZUThDdjLdC5lAHEvUB6AbAFY7xjrbnLlEAW/AWk94KLWv5d87BfpIYrcqFJGTI
odx2ZzI7oMyiquy0C28oDk9kFpy+khEayXX1w843KD9i8Y7OWvvKc5zuRwEPjULkFCB8q/zw44DN
6A716U12zZ/5JSbX8NJ0P2zdvHWMt1v0BdXT5Tn//ukAHsPas8aMoOaMsewxXKAZJW9zgsTtuEhr
vek9dzcwQPutHEGJIIg4THZr6mj9PZ9ESqpS8I7o5Lb+2IWruiUQ4nsBjZsVQCC+x/MVZfHgUn27
Kvvswxf82pME1sWi8hAYXpwS9uZNvQmxaDVT3AeNPjBoMuq6OcDkfljdwxAPOSQ6B5WN6SDkG8Jv
sIDR1sUHhIKP8oCqfOMlE6mq1gVCf2q+mcQ9tfou2RRr2mG8eAic3VFnuHBD/gvwNPd962YowLar
NcsCYs1byVQo+rsjP87BSeOrIbhnaihjPRIqTi3mQFVJ3z+U1B7lftrkwQzsf81++QmHMPjiuKUm
yjdhnDLTJnDq3mhga3+T+nlUvnCr1TtaxQF4dBAICVDDe9W/Mx1BxWhjsptU2NfqszexLioJmifw
VLJ/EFFO4Pcj6U7T5Tl9WSxhmKvPx5SIdt07a09wnTk0LlbyJaqHLuR2RltN8opoS4a4Ny15cGts
xaoONT8YdVNw1UjdaLNCKFZEUTYimUr0rWZWGjMr5I7gcgRGc4vMm2P88iAyPA8JnsY+qH5o+bM7
F/lJNZJD086LaET/WTJ/oDVOcIUzZBuIFDip9BWDmdor3a4peaVTvrlHwlmzxEOZLRt6M5Qk2A0Q
jyuG7rnhyRm0+KOeO3fQUG3yUl1FBBWw6q1rTVPsv/a4jJC0HCc0Fwy7x9v5eIRnAl1Ut5E6iNw3
6nYedo8mQHtbCdbK8TP3kUDOnwIe1OK09JcyPpWjWjUCV8WZVFqhkEY7/E6fYpbI2LpGtDyDhYFJ
INwiu5wmQph4HJn3yBpr+CVUCXnnx33Lp1Lwbm64IJJG+3dqlIRs7YrUuOw/WI8d6NfZtdmC8ZaC
T5KFgU6/9gRfEP+t7Pwqv559CTxhjRkuUzgRdxdPQKJKQ7ZW9eDfrmTyk8MuhJ5pC71mEqAT9SkV
6BGlB/LakVjz3LxG8hEv2oHkgqsE38q5AQBX+6l9EDSjlksQcgPRdyr8hMX76lXvAFeROVrTLhwY
MRZS7bvmqSYlstWbYX1T7FOBi7HBNqttRg97xg1hgsFfawM7K3ZYnKnA1MJPhMo6e3vR/1lW50Wo
XXCaoo5It3mKzii1HFvm0MrPvrF0ln4rwuHZ/fTZ36DlnZ8mo5Nn3bYMrVQ3wxddF4+IvWRvpYNQ
H4fIzfCevmbBag96HLMh5FiVlr5oDlgRxu+pRgUiQXAxTi10rVdYGKIiFhh1jLZpQyhvYTwcb0pP
go0dx3LQeRn5bIH62XGRGHmuG6b9g1vl8O1+9bi4WQeJUMoq4CFJkwXpgCuNrYXn2hy97hocIHwD
ZapBlOOmWx6juezJJfdL2kpbKw+3fp5ptM4Jj3yrBYwpLx1GEowDdk/BscspEjMR6khkMRSR93rx
xM6UrPrtCOO4zqjSPN2/40RwOQ0u1pB7XkmSgtp5mqsKGu+wEbqnt6mAeWAQqtFkWW0naLIebaqo
4dpU2ERu0wg++WiPFzmNeoJqpdAMBHbmXOf56hy8PsknSABBfsAjEdoQYI3UuZVJzYI7H87Bccnq
7CdUsSGf1N0RPJrcfkimrfRihYAyFDvpJpQQIiF/Tm0+vENnvQ3C0aqT4BLHG/A6YGHa1mMQxeNW
QbOgbteW+IDAQkISysAGljDbn20wCR1nQt4zpshLXyXWVaEKPwduK0a5g4DCoruQXYMAtV0w9/OH
flcXQi6kQ14tvrG8/gCLCLtToUElq0hg8IfeUGRTs/ft3o2PEnLgHhs0S8hwa3Y3PiGSiBuU+tSX
m30LjjPXv6RHvTfAleCrFT04x0NDJT/5ZJdrDBzhMP6tUmoVYpOVX8J7tfmqagZuXqSsyQ6BaV6r
qLNhu1WCtaZXjxj6dTr9wviOcFuWwIWvn/5KQYsy8K8wd8KOgaitgQhx9nGWbdIR+9Azgvz9hsH9
/KIzYrjaaJAHzDICkD5/ZLeRk9YBsOeN62G46TUbIxWAnhihVGCyQSzUR6ZgsVqLSaKjwOLlxVcC
cmkwhOeX/l9VkKQQhWY3Lkqp8SPVv5hKia8cXK/Qw4w2C20vCwZnpvvrKxgeITancXkpvQpOuQp3
5A/UpIcSbFRcHB9LO2AdqCKsfHmL7aIhN9mHJpptoHtvWgUiZTstzssjNDgYzEZ+1E/Z7nc58wZK
3cWJdFBIURfKKJ6A/tCNpOQAPOBdRysWRURkFFtYSZqPUvJ4XWlotdLxf7v9urf0gxBp9NUktdqn
+M1rNLeJv+I03u/9Q/Tf0/oxjKlH5z8fVa6K8k7CGjdLxoet671n/0IK84WDdSD9ImXtcrEetpAR
GUvFfJUQOfUX+2fM4ttpZdflbPIqSu/jeK1C9Q2t2VHN0A/rO0/LhTM9DbIGAD/E41DrYBjmSr0f
2u7Mf2lFkCSUhkRjy+wiQC0nJQNLyT6HVv/SXgZrMGApJm3Q2gQ/p6ByLTgPF17zsLM9JCW4oYUL
ZS5kOU+Kekhfs4MGCYDmeX+L5seTLg1hpPSGT9HES7m3+nzsb4lbHXI0oiUdcub4ZUu7gc4uWQam
eXXNQAK0oyeryQEYSvX56kaRaTsjtdT7EDN+9GQYPXZW/GeUQm9dMcFaDFhSiZ/g4zmKpv1NB6gj
S8/X8nH/GqpyeF0bhZ19NEtap72H7RqIHRBh8+Ft6n4wqnzycTrxc4gRakhgBuNHCO+4yLRwaTe4
Jy65/PzSoWkWMGmXRK1g6B1rihX0CbR2CIKJyN24uNkXFP+IsQOYm6wBW/f1DTGCWFWLQ2YuM1Yg
H33HxzkV0PptvDSMLipj3FYE3GfCgEXALm0Np0vBDEdM01K+A6NxsWg3uxODCZumvb5zAZsH0cE/
9f1TAiM000A5xrt7TRcl3txDZMVpZ3OffVZBXPESbf2KpdYFYuwH7O6HR/UX3zIv6HkvzDpQJvv2
fngs4arA4eUsRmHzgjlakMfJ/WrNos0gchflbwGrfY1C78jD38kVkYM9R0NVUkoecOLPVUwJ0GdW
W0ls8qmenFC4DWFMMq3AQW20vzJ55GER+HOnXmBRkcf5MZBI2oNgxkFOJT6mIy5y+hKOiWr/4bg0
Qkhz3ac6WSsylEIvSibx2TgF5HSKsXZpTs1KnVkq8jY0ntMJDedt73OZYLtbCO17aTtlKCVnwL8p
skfLxREWif2XPSUAcWzW/kcHNi7by5izCcFDNjRKKqWiUDhLA6txL4s38dVGgvHoe3IAY/uqN168
+K3b0Fa6yWeg6RAvM5oL1GDk19nN8yMjke01oBnJ4NcqRp14/tLHhcT1ZPHRkDNNFOp4GDTQrkRI
gSFaaBiF/J2kt5au3wIIjxDuBdtnWGt0aB2Oeoscb21QB1bC0APhY009cZYsxpP+mZoSDyBgYcS5
TxGORS2qeQcpBIVWkBF7oPvaytLWKR+/WV+5YxOyqxC3FM2Nt/EMMICRo0CsfMRzbhIvZWxMQjYm
Se/00T1X6ahnjhQ3zLtbTQE7KWH3weyrUeYKfV0RM7/tbGvbxOJ1xi7BiNWpzkNRY1zjpahuYIz1
CPLE3Jb9UpXq/udUZfjaDappDX0DjKpV1IsA0wcScy4hNNPOu4ZtY9mBv/ItDHquJsF8cS87CNDm
o3Vldr7bIvOouQS1U7aVfOiB3TJXEsXP1TRbhigcl3SiWtdA5I2mY51+yE+zmybiuSF4hHD0M38O
P0o78fNmjA0q5RpVLDmiIzZssYVQY3xKBvK5272MXoB9JC1xRZhlGsejQv6tvx0nXg/J1pQbstYl
JhhLNn55L8GttQBQwybksebnbA77XA9jLAFihmcj2eLn8zpBycB45xsjsJ0ANa+j3Ln967mm0ASb
Vz8L5Lh78Yz3REHA/P4+g1yWensbCszl4Ok5yCpTZ06y2hl/Wmwzn9j0dUosK0XJYATv5mg9tsy1
gKNai0D9RP51ze6g9Ainx5PY1S11KLWpPB+PHwOcyl3qtJhmBxuvpJM7+1THn3TR7qhnhkYcQv15
bPbFw7idVknWFmgMzlZWbkWVcc8VkjixV1wECPnBEmH8FG9Cxw9nOUpKmTVo1SWGS7ymCsNwxGyC
LhsV93q08W0vs0CFP/uqnMTo3RHcrJH87h2Tn/1j3WH1eKq7Icl4NVuAxuovKddMb31jOXKbkbXV
GOLCW5igswS9n9dVEULcoJV6z/TWASo1aKNXhFiYoEwvqi5bCz+YIe+rZWzv8KOPHZZHJB0gi+wV
fdcURoxW00szTJ3/4r6Ij5QcTXM55xrc/AyQl70yQyAuCqmGRPKGqusUswDgQnY+hsfGaCzgOBcW
L1IDT0XNeFN2OvkYlC3QANjUjDCG4SXY1QO/0j2mABbwL4QKgitbFuxo4TB+Gdb7iSGmjcXFLaTN
8Bkwhql1zYdzOBB0pehcLxbOHHbznKS9/NvKWZOCw5nSpLtYzCTpFi9Yv09rA0DANOebVSxCdIpM
txcxixzReWFhka8BzOUucKKdyDfDqWDNjfIJduev9PhLAOIAPJpZE1VSesjXI72D653SVnYPpQzV
6F/0Z/jX4xWXurxLdYScVLCarqFq8x63ErJ6CEhw2HtmL/j1Ixl2DWYUKVlE5Vk/222gKDzQCED3
UmS+qDQ4s3fpEZtUZjtqraOh9n3yYDbFIDjB7nWPXeHZE0hDo3sCAdb7df5RvGlpwZwjWK01MWlT
Zqyd4Ue+wV9zAIsw4YRh9BEDoieXdGtb4SNuknJqJl6k4jXAa9y6G2CJsn63S0KKlKQ6gF2h/e1S
Z3HIYhJVVLd0LQ70LkI+dewKpZ2gImaia4mfBY0uqiB5eBeVmORfE70KfVMd3njwemCmsMDspQRn
DHkypOBOcZbjTFwg/B98ZRmHQqRN1wXF8oY2hkO8YvEtR3Adn7HNzV2ULFJkHqGosL7ZEPLsIhoh
ooLi6H9QOtIjKRa/la7OF+6mlimUMYusOXpDWnnBQjb0hDyBimn8AUcMWCVDOeTJiO+Rt1xVPA9p
dDMxDNCnGuqc738FyT6x+DfvMW60ZbbxOhygxT2ToRUF3gNHtxoAnOdoBRrtf+lUORsz8dTyW9mF
izBN0oLdbW2xvgndTeUUZx+Awq5WYJLggs3XwJUiU13xib91vejcWFu7lQ/rejf+v65R9qzE98H6
Z/h6cm6MN0CL8ElFyZ1scPhF65nGmClRjz7YNBpMmLAV3Y6kvhUDxof/Fd915ogLKKC/zvxrC3a0
dT2lf5EJAuSV89lzUnStlehGu7MHFdFmjEFw529tI7QLUBIebWgVhmckGKJ7SzeTckr6WazPijGN
rEV+Zr9ArPVkm8dZKDx+1e70Ri/Ap1NeEfkeXxDLvb/e7IkvRnIhRmNZVHZFfmXzW4ndjtrg34bj
Li96syZH5XcIByH8DApjIa0yyM1byEbHZ3K6zl6d81kNXKU2Kmljp40bYSsjE3A5ixYFYeu+bXoI
b8QyxzqJBJu7fwDou0VUCtcsZr4EjV0+G9QEFqVLkqrptj3/vrwVsTfZO+a76M2UGP9sdO4AHoSW
5oXufudyMXePwVUT7SLEteFcE+sGKU3TXjhoiPUquwp1tP0IYRn5wzT9LaNp8qhYQH9oNcEcnA5M
nkXhSTQhbRs82s/zQ+MLoovIUi2vXBiRNWO24vXMdxg7pj+Xl4VWmQoKZl1Va3Zb7TS9PF13IhfE
Hwi9MQCsWF/VemkfPfPZSNytVXQxebJKaLJFwoeVTtSF6WQ4BSpIivuNUF9M142h9c4XMg+Sq2WR
iJVkK1mijy2Lc6ffrhpyGPnICMxBCoVVpIYEeB8Yo9CpDKK39F6+sW6f0M+9FTFGs2tywKV97t8h
JY5piWwoBmSDtZ4RzAf/XbBZ3G2fp0aNCYfXkCXRnNAQSDjmOgNf7+FjvPyvPP8rKWIZU9RlR8oi
9TnSLlJUTrbbwPfcAY/++W3nTP2TXsxqiTkbwsuYAFKBKjcZnkkmdbwcOngvC3nsdIGUZEc9QH3/
DBcnFlUjy44zMNBANwSPY+RzK9wLF5ADoQ4OXUONz+igG62E8BpXw22JRNTYwum8aqWAfgzn3wKK
X3sA04v0wt+aCAKAL8fqdDH8OBqDXJt6NqIqz8gRc0IrJRd7XZ2rzJI/N4DpTV/XNo2Y9KsK8yko
/KYJw4ZA/WT/mUjmJTRbljntNDhxYW3Av5p6oIEyCda2Gun/Rr4aR+sHCZ2vkVXf9czaDAlnqMjn
4NrMyMBSvL+J3hNnPyiwMEtiHojNdWpqD0K1R7f/g69i59rQuI+N+NGXPMpzp9dvKBq2dm4U2dmi
Hfu+84lL3DgR3ebLrH8MhyZxaHYBrluE5KHjbNKF8qjwmmlDf3PfHe76c8kHfSYjsiRg8BH+xD4P
bkodNg1i6IYCyZaNqbGhwv4KFXVaEMHWqv/jXkBBXgogV/wwqvlqxdPeQuNKQ0KTOn0Ot+3v1/+h
OzCg/pFzlMfCXxjuLpmz/MOTo6J+vIxCFFBe4E3LpktcxtY7Uo0XjTe4vChzWyFKGkYdDkN25yp8
PeVzA6XFdl/rC4J8Ab0Sw9gVVQb/IFwCgw8m9y9lOI0LUurPCLAeTQ8b7f7e+pxUMLQdBTVCg0nb
ZVtWqWOoobsEUtNcpDY00nYB3Zh6JL/O0RKhyNqi45ULvI0lT97Dtu5EVcjmBTMLmn1jk46Dv9Hc
QXuIFFdvh7GDys7yBUpQYVKsv8bIh9ieiQ6iJifsyypBHAxGC0dJfKi6fsFp2cejXuGV95smGVSA
ufoW8HnyV/fizO1YwoxFsJSF99csuOY7r6EiDNbfz+EyYrzJo2lg9NHUMrrzx4yszNbSZaw2a5tX
OMJ4s7LuQDyvXxOOlPxOIcdmdY8qJpUHapawKLArlbNAP4JqB/4YLQdF0jtURHCdH0nbhOsxDY+m
qVdzfwMb4XKKRp5O/lr/EoCDBsyBMHH1L7i+eeD6VJKT4eHujyufF8/g0x8ezrfMirVEN3rdMQpW
leOp8jR7tI7s4bd45pd+/29NzXxpZnl+F3rU5vyDTkf6Lmrx2EEKAysORCRbqixGJTzlwcbB3A34
OYJQGZ2/vZt0y1cKgLIHkPPc/+4/4DaVYuIRxNVHTKGxyRpkaxje54kCpcBKxwlDX8yP9AwMqAq2
CeD3fipDbOnFmJBCYHJA6/N781YC0J2MZNlslFMHOUya4R3wS6R1j+RWseWvcDszUUCWEA3DoD9U
QQEBXSevjpfOGejCG/toWMtcT3Yh01LKDmE8iqo8Gd++Jr6n9Xu+HjMGKaECcJiogKzTlmzAUhGh
mgfI+rKAhMkEaMzGHpAeLHou4xRorrDPEpFt5KFO9BQ+lZrcqUtYJtwsfrNGrO1NspMaJybLpc26
l6pBof6fc6jsBq09ktogxWoEW4lpFnibxvcct2IKsF73vIBcg80BKWqUwScRBqZC8vgUCMnrjmYC
iC/dJs+cuW0sByGDMfXlBAfWsN2rkghkpUZOCbLQrmE1kblpAsyOHP58WEPy5/xpRlENsxo5wJYh
GBwlxppw/O1IRvx+QuAbSKGLVrIrnc+I85VDw9tdTsDHshZa8qVXR/JfnPMZDJuvr441ddDlzZID
TZSkZCjGQe4Kt9N7pETqVnG1svl8NBBeOT9RhfRJII6F78X8YbuL0yi032Ix5jM53PesjthLog4s
m/natYC/xNO3DtbkuojXBD2C+CxoS3WYMWkyVUnrOYMmemunspejPmCp2fFvsB/6UHzVzPtjvhrv
TN98Y2yIizhdqNQylcotwWLOCc1VYxVJoDT/RlRFhKU7FQAPMhlINzZLn4QSW7n1UYlygj10XzYD
JgwCoXp2GZFJgV/feb3h5XgoZW1zQ5Zqsgt+Zk/N0zswupYaZDc8lT3/Iei1a5FL9EO2zRHnUcgD
MBrcwUhdmWkumsVUaPinK3nZ3XfNwGSXOe7c0y8weTdS+R2dyFrDIL3Q45nsTEr2cGz4qvkLAljw
mJ0RsbpDv6jMfG2rntU2g0sJDUfYy2VKJqlzNhwQsRjOtWUcImhDMMaGvAxZ8WlXKdPPuYcZJ12p
sYI62RgVDdmNri7ovziXrI+CCgzXC8+OrVLthE1sC0t+nQ97/Rl9oANILx2eKtvPF5Bgf5iqrfCx
8ad6FrWpUfKExnCKrukQmC66340QgV0aBm8v2JL63mwx27eBZOXPEpkj88J4q+T8omnE5osZsXzx
DWHGwYdqY/egVUKCK1yaWSL1bo5YGHofWevls/LsO8pByouvxA/Khhy6DbiLYUVMvmcxEl8aIB5Y
GhBy3kUARnFz8qOTmiD4gW+f701FMBpqPHT36eqTa6Htj5iRBUF6F1UE0EOKOa1Q7Kn13ugBOWEr
VfmiwSeYYcvlGUfmEB4s7FXUNi7vZQiVIQCUOuRt0fcE/AmJyri5fGR1iDRLK3T8K31exQ06YRzu
Zwbc3tfGq1dA/almTKLEJ/zt4Y3dNFLmQ/e7UVYb2cQ1XtQLxcCIJCk7M8B3Iwstrsjwpdt1mStM
xQpo1lpUwrnBkpPewVoIIrR0RQAPIZ8iOQES5qKn41xbDDGlxlAh/nMA5u1aknKhHGQzmzhNdyQt
nhcVrSKmldtcL4elWXDpG5nriUegJyYJA6UuBll1hVAyc8KzCWTvBennVPwdf0tbXmwe+Psoggzl
W+wAzbFTZwiA7GC5EQe3Kq/eUlmUq+9p8SfE4wwLqnhsI/6RPkVqOKRLt5VgPe+baanbPvACgFQR
DTuQxACxL3p1NmTivM5iDpdBalt7zOnoXxwMW2F/xmJy/m2P8nn9lHO96KkEND4QVJbUrY/+ubKO
ZoEIHiAz1TEm0IeKBdHhTIY1EZGXN65LkA1nqsJ9DNzRS7UeoofyOvWNVQDTdQTUuQg2a6eNfZIO
VsnpUFoVL0m3f5q7OWHgwc9Kv8K7GRCQlYhrX4f1IIBgCd0ofkEQwCu9LGkqv69BGJjd/SBzr4/u
bouGfWzNkdMKL/b6PIVtm67mBpwlX0xN3rcxhBYkV/tcbFl3TfX/p1caATD4UQyDocn/c/wlEpsY
1tgDaYJvwKkk59As15rO5gw3WzETpWFyEJSPtKxQMXqn4Czo1AzEOC3Dny8DJTtDcpj8y296ic+K
sqnBEm3gBu2crHyO9gaGpbnhgMe1Vn2auZGjj+V029F8A84fP0ymMq4ciMUk9c1eMyR+lfqFgqGM
b7xmtGxE8wbRad8HZd0mqfNgmBqJRUoWkGc2/3lJujhIi9Jh6mNtjv/Ual0fwyNrCBkmpvPn+Tkm
a3gV2Cs1Sb18huIp92nvnyhLdAAx94/o0Mr/iTgkPbAJqixkyc6A+j/B7CqStz+5b12BMJJ90lp/
gTAfExUrdr5wdM5bQmDqDGmuCvzIAgCnWF27Hg8xrSg2DcSPIuRC6CKxXicT2OeLQ3Yyp2lODnPR
4HZJnQ1FhuFrlqGD/hXJN+mtKGOmjt1riIxLuAQJjPDrM9bRJj+JkFHJ2dSCpS2BgegMrSoEKuO+
gi3rLy+PmNByAKc1yIf8kIq3AFtrcQ9jXGusv8VirIcdhfOXV9Z5sM0hirrzi3KYO2WQToxFBHiU
DmiYOMJADK7WaXUZS4Z/SHUwMcJuQWw+KM3hET942tmVgV9RZfliB9Z6EYbZG+TtyEoPNrrY/fwf
AV5kmc5X/lfFmIFFjmeVfWXIn8994WWxa1DKEmnGokRBK8a20lCeLcWIai2Dp1aFEYBCNmpFGLx7
RJhq7+YoxgBp79Q0/nJ9hPuAw+bBSRkkmNJBVHPF8FGGYGoZfiX8YCqX3tzCkwYa78x+zlit+BWh
a05eDNey5egDpVD2JI66zh53gK9tC5vD+J41w8mpagms0qAm3C1o67zeeh3U4fvG0eo52Ir96TJm
Kg6FJ9vsW1Ka+o9ytXXa2qUVxv7ytgEpTQ/8VLIFx0NOkLtAE+3SNt367VihJcm37sNL9XH9Owuz
xS71N3BshbS8h3NADBBiBkqxgVuJu38sepNPHydsiHK+A1spwQ+JF1q7nM+5kCIcHwwesYcBnvsz
iia2WdRM7P+uBQWCQaTS9D0K66fCHRzLEsmeo3dWu4lJpsOV1ng35Nl6pnVL8km9zk5+VvTjDiJU
zzf7JefC3Ne9cFfdIfFpIjBzcUojOl9foJjf67XZH3vQaScsiihmHLwBf1Bn+ZUWs9Ya9chXrUTh
B8sxWAZFDOmaj7aOtftpKtae3rh/VB8hvYWYJn9uS3JRv1YT7Rp/pwwyJvMDSK4YtkyDRBHGDENE
75Jr7pHgKJJ1BBUK0pR9lxBGkNKfTK7lpKxeHasJlDVZwg/cQeE8ekAbw9EIOOr5S2oZyU4YQzVg
swmpPm3wgT46f27yJMpgl1iWpUfxuyYFK5/TDtyh46ObmFgNQ9YbVsgOeXSOVUZIDNy9FGOGGIIW
I/9EhC7mDtBaNPMoXdKlS0MiohVUHJoobpnc5kzSFaH/ihX2zlj+lquRaRIsUVSLw78/tHHIizWv
JvobuyvMNcIHcv6CM6TLS2c607G5Ic4vNlYAO+krY/TGuyB5u+t0Upemvn9fsjoaqeouywR7O8C2
wXai5PvhzMb3U7ypj6HTR2TBi4qN2g2JIeCd5oJKPMH4ENDxeT7LpYODflIJIcgA2rcfFq45wE3k
ZKzVdz1JDKp+1L8DtpPbHOVyGpfe3Y+gWUORW8nGL2AuRgNltMB12V2zoozSHwcmYNrijAwsAORK
LP/1VT7BLUtiEdaP+QmR7FBgHe0lXtTYARoF2Hj2VfFz1VS/Jl12/5VBE4k77TgsEzElzP25+cYA
ctnpoo4XzMqqyxnytGbcaPVBLj00IHpBVPzsNTQqqe13zfp4bir4c+RBA+3MqapW5yNshsP0GRsd
dcgxlS8Aj0MJWGUfSqmvsTqveYS6cm01FnpnNVvzuFVDnt9Q87F+n4RpxBw4s0rJmw/C9DBVhSMs
/FxznAt0k6ChHGgqoMbvMYprp+cdlXeCuPVYioyI0s7FQObIheAUfV/kHp6MFESiaCHHoIEieZKU
8eaRAjkPOuP51d1r7yA8baSwc0fXDKGHYc6Rm0Wg30/6ldzycDgS2YU/+HmbIpgPLIfVozDUmuzD
AyG0mnHIr6u6JeqmZxaei+4/rquEwM0hSZ0z+lCVVMNve8VeaT2CUtPCRuJbpnG/J6z97pMegH8M
Uukf5LBHyjLp4g+DLzRET2Rz86S6ZjyN3wF0QGlYH7cb+5rSyB5Hm3ATTAiNl+9Aww8fb2OIZh8Q
wX2pN8cBqCt6J8ljQ/vorkE67xKDFC0DSAqwthw1H+aW1to92eQEE03qJsgjzu0SkCwY6+eXYFn2
vVxXKq+//I06AtaOfvEYe1XZcdC60XCVyQdahbVs829L71wbjHlYM7oNYtzfGKBSb+5NmN7hVj07
ADbBJjxTXsLHHGEU3qfs/Fo5Hntv/PyK4trFbnO5fgbqivdy7QSXZf+fyyGHvEAEVFicIEUq+eKX
FH4xJFEFLdttvVzqmPOcIgu+IYNDRmIPqGrCoMcfAaBJnEwt740n8Otw8FewLN49psWond7PlPHo
dv4AvAZSMJdQHZ1wMQyIs1Xro9qlHh7lmAbbbAeuT9DLwgUVV2/4KMABUjzZKOeb6yYzcg/fxbnj
413lFgNs+wJmDjy9aaR7clcZeKntdzN2lBP0LhK1da8ooY63FnefFcM+28JANKCOys7l5/b2sijA
pKjn2oG02+3HU9DBcWH8eFXXPCnJcmY35KIabH783MvVcccZOTZMyBWGC12iJxmDVi2MWe/gAnu9
VZaFpH7hCYdKd3VpJg5vqF6Ao/ba4p2POgSJ8oQH6YlPR45iwxMoCrjtatBxE625ZOzI6WE+GhOn
QB4Vy1DAwXZsspVHdcn6v2yEKHOTbRmZBFBC6GbG3W44Cd1cIRx/BJvIfm3olR1E+0yyabDS9cFh
t3jLJTgey11ZlKnUQYC2JpVSiPgR4nzHr58/HanoQxHH2FnmqykveVIwxk4KAXEJQ+LkY1vHqJDE
ye516LspHm0oTYnuy6nFI/kFaFVJdJ8TA647YEtvF2b1BuClGbZ72a2Py3yamYmSuY7kdPPMDqTj
x0Uqa06K8tOmqr7Tq00npTYnWakWbNIUZlU0/8wgMp03a6WXQBzdeWth1tf3cxOlBERBigqoamhg
dcR6TjCsZ9S80LkL+RS8DlzWapffCSaEUAx50kxqyhmfJru1wZhaE7Bl4h3WEceQiKyldJrpWYX0
XeEi7SBTGCi8pEZcEuv6WilqAWiew56A79rYpqMzT1SoKsofn+kuoQW77T97n6mtXsop1miR4j/a
ry9wgxlIhrKVj40+jBpgNSsKjuFiwY2KzO+sNDrB/dKogJv/gKXtrx+d+r0jr7oBNiEO3JkWYSxF
JyvvypXy0YA5esjpXpIaKfrtUpfhgDNy/4SSbW0UkTUZtlI7JZNuBrObobPGqPzsFTXHMuPAJA3d
QeZyWu4zryqJuN6fyEfRibsOwVJBD0+Y9ymhExOduDqjub93bi4+95of2pM3uxpgAUGzUuGHZ1Jk
F4yd9J9kT6edUw5oV2XNzfvc6rXRdQ0IWlNJoMmwoGzWRb8ERv6V5wPWmVY+OFUIkQO+t8DE4QNN
r9ZBR4tlBYS3IYHTpbpG/XB7D0IxgFo9EBt8fwTDPgymh4CPZXRQ3SvbJT6VXqgji/uC0zdxo5ya
PO8HmARTh3ZX198oiD9P+izt+OsKUhpzaZi6VhRw8ofqFWPm4YvgCYi/No/FTGPS2Zd1sZ8aHx/K
2rmFy7qYGs3+r11NqJQEDKXXkHN9qEwVPOQ+CU8IHvFWineRnvHvFv0Kt0otNCUhvqGG+KTHp6fa
mhlNw5aCgkB6qsmH3E04s5krd8BnSfc5wH5cqeoqJmhYCJhaWBZD1GLbHfecD9aLQQj7eEjWrl6x
Xx2Nvcn3cNhrh6Pj6HnDT194MmLX7CqoMP1dKqXJQV1720q7qQW3pw==
`protect end_protected
