`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
CqVA2OrUEw3rS2L7wrnupzM2b8ryA3Bu+lnJvxgVgrjNcEfookBm3yP7nJiadlfzz4GXwIp9iz2p
s3/zJCpagw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
PGdlKzNiAp+RfljaUz/4qWu4UrsaDdcb5I8m2pHEh9Dw5NlzkSTUrehmIwXHdNZusEIuykWSAGWZ
/B64COg99vwXbChOMVOzpixzv2mQr+HqmujYKEqSPvVqZcYkaJU+XC13dHTzB+nF8v5xP9lv8O4r
vnd1MJemao4IqJNNJS0=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
O9C7HpJnOAPQ7vXXyALA4SPMh/k2S46Hh5XdLMUYWYp17VipkHtaPGZ/6KFccH6RFn58ICZGO3KG
sGL5WYBNemFQqBq0y8svyUk+CP71thqm1XgysiiwK+cLbzasmWv6gd72IZaDJ0Dm/koqglZz9rGr
Yy1oI9Hp83u8w0ZrJCUozxT9sRuP6Hk4NriTgdm1bEZtEe/2gsoRGZ4uypGCTZ83caU77u5XkSG+
sY0WMUN4I9JDArAXRZlcZzwLEYJek3pwzASxa3Ss4SHc2/ugyBQEnz0u03Ct8/oB8h+AKz/WBsKk
FtYCRL0FkFN7NG6Rp1n4otCijlZmPDy0sb+V4Q==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
UYTymsFhvRnh93jsBmiwdgozSwCEH1PzuBioTnilEvHeHSSg1Ob7Oi1NUv6bQneX5bC/xEpsrKCF
ZzOktRibPyX+3Jk6BpXtTU3T5z4D8X9+eQTazzRLlGFkOR25EDBRMKSnXfl6zR1c91u9+kYZpCtD
tT41G9m2iVNn0qwHADM=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
EKb6oPxzLBvAKIrzC7UNBK8eY5ryi5iGJ7/BdocCXYMaivf2xcPKTIiYIkE0Hv8PshEsJ9YIK1VC
T6c/GEUGhuDsDpN8XNAiNGvxpcj+TImzhi0UBgHdiDVLhkJAtmhW7fOxixaqronVrRDaXAhWqA6z
eRM9XDYWonBS/l0El/PUUSoDAWcnU5LoHeBeSG8Z1TM+qyUa7w6WDqALs5O4HEYB8EIMehKvTcBS
pzbXxQ5k2wT+39vCq7Vncv5YubiSbq19B/yvttj/idZ0/y9fFAXYHF6USm2KGjPUs3+CmdnaA+hm
Q9TgqJDQ8e3agIUv19cQIAqFNQpoClnjhD3haQ==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
VT15/X4T4V3jrHxVnZkn6UrAuaA2quR8EdrkmUFjWmWdJf2TkcB/YHt56tVEUMbBtX0cu4OhICAV
5m4ThUbdpGUSaVYCFzK9V/BGPk159BTr9sJRQ450Co5g/TE3faaAIaUcLrZ3NPDqDbB8RYHXBpv4
SzpcX46ohjmLqHyCiSUO9tAg3SQcUm6kjbRntvPdE/PWVqx8jie33+EUwa1OD+KsIwM3co577bv/
C4E0EyQrjR6YYD7VCJNxl2h7GqVjE2qMqA0zrYZxk7F6DpgH8zWoSyd32pPOkBTg3YVuftBqGZWi
Vb6Jg33JUZNlOQqE0SjOJRpR8BExFJ8BGHwy0w==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 57296)
`protect data_block
yJR42fHc5CAsXyeEoKbA5A8ApJ9SCVRK3c1RrDrhzDoMSwonsfHavwO8SsGKzDnFDonM1I7DsSoN
GYVarhE0hDF7U4Hd5vhFCzqq4MJSr/l2ci6xSK0/6u2C7oEJT6qjKmooHgMlo57fM0eJDBFkuX+A
UqJ7B97NIFvW9zcSRTFNqKe7G+y+Rq38PzjUjUMQ0TPeAftsAJLTagrJNq6DHQUjWuYVvVxRV33H
/Rp3dj4PA447v9bkXeNH2+dv8vu07k+zNxpAuv8DgzJQvR9b+zFFgsW8dzafbp+dc+b/GSptbnv6
Af/E9ltvjV85gePD+LkRztPf7fHMYkcDShrRI5vT0ZBJz8cQ9z4cgFKiZQL7XHRrZAMpA4L2Egx7
DInL4YsoI7IHAJ7xtiSQuE/nQu+Z8n9rzesRw8YNvxPvUPDa9pJRvR3Ji/mU9rbhq6LwCQcek9Nt
+Ku5PKrZx7HoQX8Xtq8HoZGk/y46WRTnssjwrEMSMoHTvUFx4pqT00j6L/XmDx0luN8xlMg1IsBw
SKhIDYSN0XJEVVQbSB9Whg05YAJRRMOrXlAUHGuONeWoqMGVh338VStRJSNKTYzitoI4x4zC6vuq
s5UHHDpv9XXW2sanIdVlOjwSFWZwG86J7vH9Bh7yR1d2Ph14o7Wh1n+S36d/KohB0m0y4jnS//+3
oWVKkc9+M18Obi26iu9ilSQ0qDfG+bPKO5BUL/zHXgP6apvYXsjqUZAinWYjBIAHmURirQUfBUsd
hwzfU97RBP6oUp+jfkCEdJKWo54bjiPtwzyF1IlzkWhy+wxhpQPMeHIQV4Uo8tSe3Mvt77skutVZ
LhPW8J9oc+aMwiBLdAVJ8S0VYAjFwMjTrong7Gha34b7Bub7wSZ1GYEX40nOjdtepJ3RvRzHzZ6W
tRdx7MJn2dOvNCgxVMdsJRaqoRWqSGsxM8yMJXrzV7aMKfScPWitmdrhRYY4X+SyU+Lv+DiAs0a/
+ACNOSVLYRelK4+YBQEvzjiJqstuKc1i2cq1JQs8kGpFCca3oi6oQOJW0l/7zbziEvlMbNJgCXdn
BF5ke67Ia/5ccuwP9Uo9YPCQaPA7AYzM7MkY4uoxR2tIgXrHO885vRT9POOte0O/q5Nkgac4owZb
mTPiLXWayfFVih+AZ5ncQaP929WzX1+KKS5LYCKKNfJiO2E1HVqZ8XbY8LxF4/KovMzruwpqcog4
bspa7683BZsZLaIQKcX8qEw/n0FssgN7DJl9CNDe4SuZROUdrWRehfs5jBe5J2OaKeY34XEUXuMZ
a7wvvXvm8EG9sRlqABYUF6+kQcP79WfqohRfFhG+iXBVS90v5u3mirhhL/qJilis2d9hBCZAJ7W2
XoqC4gQWU7FJ9TEI77KrxGBw2dprqoubr+yd6tEXMCXQfZdBlfDL5/ofoOHYyx9kS8AuLWBhtZJF
Z6b8D4QVPd6eFpZwmLeadBMlLrl8Kkhmp3ufL5yR2K04H1mJB0u6YRSD3GfpNTwkCwPB+vRCvrtQ
kee3kjIrLuo0d3CYWqHlr5h5a7PlL8l/IKWWgg3ZsW1tcx7xVt5MpF7VSQA9ygmWBVLZZEMTJM5v
VT2NtZJa/hVngOPycUlgfGG52OnQJ6r59s+gU7zEVmLYnAH0INbZmDRv20QnpGB5UhFF1qocBWZE
aX00FAUXqlgnVjvYaNLm+2uaar/bI3VI2iSOP9XAa699J4tVUMf/gg7sHL6uOZrUWSJVNxqgIWQV
y11EvqKda/wBBLYNse+xuioirMZi1acdJpzB0ZHUV7aUpDsSxiQXcFPnnWm2QhkmDYK3Q4KACRl+
gSDz5l4VnIVmyyfQWJFKDYzH999gbSnv9JlkpmViJmuMKhfB4JQnyhKlWiZTSysnTYgHAWXYhHlz
GoMfPsMPPN0CdstDcva9pUF2EW2wFzs/RrtdsZSjIqRpnWAqlpriaA80DQaJX0Ffikr4Nyiw4XGk
VZSax0pjVQbcRee9UaNZGpq08tEZlusFXWhSd86Axmrp1H9SqaehURpSwYSLn9plZjiI7R8arYTf
trexSGmsWfU2ynZQJsdGr+UHnC3cHNygjp1K9RdGjVACHVZHtgOTGxTZQNE2xe+mx6E2aFWnvqeG
bnjV6iaLZAr2WHyrCQ3PsNbOFLiPzy6OcpdjBHFgLIZsWykFCscS2antXxKNsUJsFkfavG9K3LKH
8UN/d8bbclUyThToekFs6TVuOxtFIVCoRLZwakcmXuR0uPlHojQVnV9BgMyxtY0mCMG1jGQc/sOq
xig34cypgtsBvmRWhknSOHBj8Grr6lYCb8M1rcSf7ZGvHwqup1YeoqjGUOyH85LWbd9d22kAq8zp
cK8y/ssg7Y30uAicZj8FRPui+el+PIGFQTq34TCadTwuNvfH/vv8NIliCD0aWD4TtJdhv2KulM/S
wGpR9iHg8USB48rPj8awXPcPJx6fFmAHI+WCFI8XURUF9wSq3mFU0uZJqES29ITNeGT3ReGSLPfS
NPyh9LE2I0xwVYyDv2nNHAHjoY9N49RJleBTm26b9GL+rvCY1keqkv3ChgOgcI3cfyGPUTG1B230
mGHg07vCeA1jEUUiCDKBCIaMry8FmV78Ei/1qQiDrZcatWM6PpOvflVe+ZtCtqkGqrObdWtZ/EjM
Y2ooOW+PpQX0Ek8EiabCK5wDBwBJmboy/6tkQUFsjDFQtRVMnx8G2+zwEp4r+q3MJGn94kRHoAjo
Ptki0wx5qCI9KGpa/q+d0cwqzSspg+H60HAOqYaHzNENTJ9Yq/Sj7L/31Mc8o/ngPF+aKLHcRANq
PNu1i01JO9TO0fjiCph8f4SOhEpiBNXlgLJXUOfyJ9foyx7o14J9R8Kp9k4wR0XLwRn6/+OCzFHY
6pP+SlgxUpcp8ChYREq1qEUPEtRmmGxphHfl70LjljOa9aqn9KK669cQc5ZdrMit2RvqiK7U07et
V+nGk86PkK3d7Ovo2jYlQUfACcagnErhBPV1IVS1FzEo0k/qCtNuIhny/U6xXz0cWYUbwT1BMhMP
L3zFRj95BruRQN6KvPwOU91KJ/yUEtDc/SM6mR0qigoAXVpGILa0K5/KPMKGeTbOBJ70KIKhjBO9
0Cu8kVHtidnQZEZMUIFJimUMj7Ha+my981c4BnUn4WmgkV99qhvgT7Nc7C3a7EyYp3tbPkOJRyM1
BDN9nHDHnl96SZ84/1S7nnsdV669a8vfAl8MmlQKr6MDyIE+1HyMqsg3v63+etuKTvHsEifcLj1l
5JgwftqcpDUPLr8hTfljUWE2vgtcQaim4yutyujmZt/k0qkuZBUARMLBCgpoxaFYBc60WOsHjNDI
PsPIE1OititNf9aOLYI2ImknKlEXKB1G2jBsu0qNSE79ooiZnjWcppKw91qW6NtwRcNhj6GY8gM7
W8ALGpE4mh3QczTZHBFMLvBSof25heH7gKT8j436uAun9edj3oymIWSiktkPwINfophROGRwR1XA
urDXjT4j1pf3RhmsEn5prZpOXmcbaMT5XPi9ZYceD1blK+KyqFpGlgMFORbigem+kj/LvlsEz/xF
AEpRTDxIyT7HTlb6sELlle6Hug6soLSRL21u6u5tYB+lvvVxsTqO0q8oM+q6h9P4s4z3ipixyM8X
ItsDPFriTmjFYnuoEyb35uo7DtaQlLtUGfUV220lHCx04oxH9wMR+tOgT8RclBaIl9g7Qycv1FvU
mfhTks7Qtj8C8zwSPKTJ31Q8tpc4rS5eX9BdlUCdXt8VqXpueSxJqCgyCPlU6uuNteTSxzkMV/R4
FKUj4ZvlpeK8Dwsmu0hIw+xTvKrIT9wXaFYmmWK6o+IkcKJBgUw+ZT8gj+BzvcM7GIM3zYN+jOqk
8IfMBod2Qz+fC0wP9G42GcWC7e3lhLRljzUMD7FYAPmAydjXFS2wxillkVGeqYk8JqGFK0Psmopx
B7tzdGeY86hrK//aslSnGy8v8n3USckVMzO4GW0H3go5oWjeK4r9iI0zqtu4jUyQvuTNKzCfV+eO
cNZWRpLI/Vp6801g7tItuBimgKWcPpiz81nQr15CUZdM1ZJZmsrM4/ykzbNU673zi3jsprQsNa/p
eekzqAn+3GDBmu6P6d8Ucqjmx+Pb1syjDsc2GB+7G1O9mo6tQTLl9H2WWxrxO1OGA9DoOk502R+O
UYg/40H8jiV86S8bZE9D0riUZjSiAHAcY7/DOszWTtIgFC+DRVt2TF64WyYM5M2vntjBw5xKtoI1
4vJCvtKLrVcxHwkFcMbURKlgHiPqHnWYf5z1uSA2lHu3m0l/fob+3Z3Shb8qPV58o9+pkZ0k2Knw
1tZPLhz920S25LSxNBzSRMeOC9EXT1d+M+bUJC4kopaAUEOTocU8hmjjYyQMKHRa58gGJD4PO53g
XGYZBgiRJZ/e/FgDMj78IYxKZkovvzalg/vUMfA7VHzX/mR/lAexjxKrqGQb6C7IfM7mcqTCptD1
tihNxU271P0zHxx83iXNO0Wh1cSeBTjL08BDXBg09uFutJXe3wkmGlPHSsspZ6/hAJhqZEevVkEX
x0zVBm0mIjqiezisUxfF8mONfm4I780zTs5vjwLQ+BzvL4aBJqpveGb55yEd5wNpwBEMsn2Md5Ug
bKPiYR4kVhkFqjoBXaSeXCGZ22yIW2pz2QOA1N2VodcgSEumBiiulPHTJWXA+2Oh/SXE4qRk9ujn
bAvtDrToEOUb2c6A/cv3inJ8n6RE+iJUeUbXTCpgvZj92r96Oo5V5/3rS6DbJzDKK1atagqp/czo
WtqxHFEoen73/qZsRtD4/On4ogC1u/VD2cZkZTCQmRN7TKrla3dtNsmo7lcFrgVdlkluOnZfpQsI
GAx7YY8Spe+XquTTLTtKFw31AjCu5bjpSa+zcQB1AM5QHl5JbZkuxkOpKdqNv+cO8K0ItkSc0nK2
v19la258/TfHOdhlZ2mRcasIPCwixOtfeuYa+H+DzcJNLOksmPUdLEUx+KtGIPVSvu1dF3OkUH51
tb6oRsf3XjKDLanYdDErzTZv3Jh0e/X50HQ6hZ9zzcsWzNOuFn5O6XqISqtPBCxVTHFPtu5ukbSe
kOe0rSxjTcrmQ7kVf4Ms91vWeq6ufbz8hMv/VmQ3Jt74iRmzukoOKgbB23M/VTsB2aW7F2KZ1Ey3
8haUixvsdM3ofGQw+ZDuj7kX2wT3qVVx8iewsset0Myd3kA6VDy8iNEmRSjQlFXXDTyfnvckqZB9
reoHrAXkYjcV24oSUJqj1VhnW7pZmiL2SlRPsVf2nw1wHyRgNY1X5vPlXR5enqhzVD9BkU3mwiu9
L6EyICLjpCts+8faTC2Qztq6bX2Snwg+L4Exgx8pJ9NnYYU9xWw/1yleJOEvrgG1cfUFS/N+L+ub
DAIl0peYaw79j7qypmFW0j353xPeBxdgMnP3xh5ZrYNGEF2RBJTS66MTWspaNi36HXsTZYnxUPQa
Tp3TAdLwQcyycIhkBW5H4RTWI1Sw4+8KEvSLHL2ao6OG4ZPbzAIICWukME3SPwBiksQVhfHhcr7T
u3uHhdUbkdSDkcWu3+qFNCPbtM6Xp6i1MmSbZ0vXeRxjC7fltjaRmBCpRTNTXmY9yuLHM4MBfp5l
IWcMqXXniM5HoEHLu0CDC7BxTMcPna6Cu9mouOsypOwB3MscZ/JsYv/24uhD0hBn8mieQaviS/A9
/d6Msa2UqjlBuV2465wzwZli71SVFdCH0mcOhu8YNgf2YtIc/uVSL51fIFdpobyNldPr6a4NXyoZ
QBkr/B/kurIqV3poxd39NKeqVA9NlsCAMfixVJStImC3YACdayw30kTZwvNPAq8og9/hXiqrp7/k
5KCjWLBFASYMVfX3BoyA27OsCHtD4PsrnURTx2HZSpW+JhJhH6XYhFh8r/nHM8joLRARytDTjYy4
rK0VVKgLMuZP1nVhBReJk+6f7IzolxDofWhpQKMJfeCuVs++faPWaNuxBsczKbT6t7WV2qYPHpHp
XZbgJrLD/12Tt4O0GstoSgU0JCCn+98Ig+S38XI20bxOha7kbjL+mX9a7ixjS66oA9O/we8ahZBZ
udkK2swUgC4JmSvy3HqQr4RG1QcM2xb1THDgoLlCbD+0nmrUuikv+FY4oM8L8V6KJ0LhDZxSjMCx
C6hLDrlSugl8KaIejdW+p1EYNuZCnnuMgxKJm04ibg2eScCnrffuMiDOqaVTv4DLgiRGzseV6kYe
EpDr3nKOXW4e9oCWd3HAl3rfGN5e7pmKuQDcfi2xzfkfNGtl3NpKQ1CRYse3nC3CaHOdpOHrOwIE
2weob9v67Qu5wAe3T9vrVZVWTV3XdOaN+/jifaTMSty57L6pm4Hu9Lw29W3euSe+HG0oI+16dVAs
X6O7K9eCimcIZzx1w1IW9YlaiUatzGSiyTTXAJbMvnW72yFgcK2RR1FUwonVDlY0X3R71bQ0SF/Q
K4oFyHZaSy5JNZbc5ZGRERCFb8ascRM4lyt60WPYUaC8+LsGc9I+XtYarQ0gWJ3gQv4JLNAu+XmQ
cwEKrfnF8Ib1xzdA93YzvLkJ5cnN12Dt5uHv1GQAHBRIcHkg9Chb1PSQnVU6SCb8DGpCDlunF/By
tcb0Ig6P/+rGrvZvbI14YDw35iq+rGwJ4+iCBvvCAc+M0ol9D5bYEBcP3LeWfrHhNEd44ot0HpLu
Q+GExeaF5kwcPUL1cfYEc47SNxCSMXRjZv5EFHNT6gk/zzIK9ZIQB2ByxgvCBjUgfYBe6QE9aAep
YpM5dD4lq1AE1UoKw4/9EDjfSw2AHw3FnDC+WturcWTElg5s9Ih1aMzi7CY/w1k3peBFj7/Seds1
ZTsWzbNDdoezyFOsv1fpE9ocDqlyLRSGt/mcTI0sRoB+63ebYDPC8x27PeQ5ux6uPBJFCQll1F+d
z1+1IoNe4xvLtuQxtU6fPI+nezuIgj2JtfQhEHUO8MEn4ylzDaN37XYl06aOj3p88cBIOGef3p0P
YJuwM59dlNXxLGUnz8zZNTqZjL0+0BtT593IJl0uPyypTPjLlVDH+DHRk1WuBqg/qYx5IQXBP5jw
rtuj22yJg1iDRqcRLpEI8cCwQ9qdGWD9CzM8FQC2nVwLNlhdA3xyD0b6zeoWUFYsO6NtTU2RF07F
xMv3jXtw7Ai/ZDFgXvQ2Pf7xdQMqBeWmxFtrvzCZrwLElzDIkhfUJkUVXaZgsKYg9x8/9KJvmXuH
YmuWcMKJdG4NYw1S0bS0seH3Bc5hXPTgIN8uV6SDir7OByvk/Ag9aCN+drT0PA7WgHLfQRKt37ng
k0ZPGRt4AtP9TlnlzIeePlBA5sZWefLJiAeGv6b/MJR+i5d81AwSC7KTEFBPEU4T27OeMh1NJ5+S
4Rhlw6y62/y/9vcltVcgAXzE81rbKkZyyAJR6Q6EDk+EixmEOTUBunJ5kFKpRS826kM63Qx5nkc8
rHNbhTeW+9i4QzPLa6F3cOSSjVSwqj0jTYZ16J/I5HDL7mavuBDBDV4/7GSl84AwAau+pAYjCNmX
yCXfr6GiH/AxFbuxo1UNCEe7F2lW2O8BYriWXFgD814ZAS3p+M+oiqpUM4r/8Mg3UFq64yXcnuCX
DZEZE3OMhDm1oYngEfdx/ZwgqRqX83tHbrHWsfizjxBsI3j6yw2Wmoy+yv/R+eOenpnUTwnn0Bd6
01sD5w/lOTqr5jULdpfOT+2XKhvw3gHKNce4te0MIELUbK9XcpVZd1+h7PKumfRjvZFxX30W35j3
Dhxrg5hYQ3lLRBu4XLyusXL/EmgMCzkq4pW5TWhbNQ6poXOAP7yQngWxuu41rRmg7sZdmu3Wl+yl
lhr5zDBRD160omk6pOc2LdoXMl8yQLH1vRYTiMscd82ZPlTQYN6S6NzO3oZ+GBiwL/r0OFAjel1T
qU8PyBceuGG+Qm5E1n2qVdXrFCu8D+EEg8uiIontRYPmu9QKeP+ok4iqsBqo5/bUHL6UcCive7bz
N1RIW4uyt0+392JgvOn4mOpCJ9n4EovVCClVacj0t2B+2myPKm4YDqgP5dOq9bIj56XBMXlDwc4x
efjYkPuodIYdlHr0OKcPDxQtqtUgNTNrTdMUlxyU2gzoRNa5MfW/b9tJU6REi7ahYSGk13fxzIHN
hybg3E5hk0ogahKiJnoJZN6JF+rBdcBZClINgHgX47WvgcxxE7MQ0tzuv6S8XFwU0+PpzCtDFB1r
b44PjPw2kLcS9hiMqVxiZO6Md1uxdE+jhlWgwkpe7tHGiKFj0uEmUMAljvQjddTKgm8yT4tMcmrm
qrSK8aC/lQ1ugwQP+4yKFLT1rSfyTG6SGQa4zzX7uUKJ0HDqc2VPtm5RME0lLomQH8aSsPxi7O/E
2dRasa9FlGhDyuU3sbRnC6NqQWFn2RCr5iQqCu103b8+KvMvxJm9aVhDLFYWXAP4mqVP30YH77SH
AOLLZH70MNhDmychGjITyRCv5ECYOvQtG3x9j19Bo8vgEQ8c7ktiT8aWtAU06zm0h77E2HYcIHzG
yoR8DFvAXJhc3LXlU9iPAw4n3WbyrDZv0D8wP0LEqM88kxNCAdD6eNmzeSbC20dG/CC45epVehnM
Xx7lQ+0NlDqvDqiGt2iUd5uM58g77C7S6zD45nRH/zPDkJYFXTtosLW1TXQr+SbwZdiU0//XG4++
f4ii68KoZ6fPGfePTsEv9biWT4WLzk2aJfXZ1vK8GMAKqbRw5978UpbTrEtWF/GObYJVKZlBtkQC
dDfyL5TR/kQT177nxfz9JWAWHr5cIo5aV6beIUHEyEBXYcfgTHsmZoyjaJn5fbqi2DfLUBeomI/I
V3/57yRawbpYSijREMqihwHPf40i9YJnxEEC2ih5SxbGND4J9WUNej/B0gBhyXSNxN6A4uXg1b15
HOFz2omP3hsaoTHrHwAGViHa9/iwaMEYjKo4kwj0fPFnHtWKaLEyW3Rh52xObGLV6JFA9J8aZx1I
hlcCpfOCtHza3kIuh5ddocuROnfOkCsCsGaFkCZHgsARBUJU7Ga+SLXGdwDdudJe1j8Y4pjgef/t
U8nMWzA98v54ChPzf+MFSZ8rRSFu5RwsvKMNJCA8qa7TTY3I7WHOe3FB/EEUL/WPMVPdkHVG0zzU
olDOBsSlY1KHCyeezjv3z8FeofUxCXSuaEHbaHH0oCnpg+8dOwwjb3/dDMLI7Le2H5a71LBAc2us
04AyHBSPzp9X4YageNZsayojkM+sbxjGeG8/pM+tdmC115c6kYiMcL27P6/J/TbC6cKgfMd5+nAn
clkgJe37Wm0/p1526Bp2ZLs7tIFcuVk2GAeRYM3TQPpupi1mb7xy1S742n1HvIm/Sfo7buTZgXDC
1jkiv145wfbtln5UUAN1CczLBL7DzSrG/hnp+H9wruDWz32c1s7rJx/SP0kw+upuKvW5oixuDNQX
h22asVyVViVmTsCOcfWLfGxAZerTi20G9L9FODiBtuEfGGovHIM95gcgEt3sqEL4GZksZPrzg+mw
meSQn0qGqnQpu0ihzgCAZoWk+X0fR4QawgGNb/AkOAtqCiDS1az1hiAImn0VlQo95Vb7Pnjmox7v
+Q2oEW7jwDuxrbwnHcRXt3steYMM3BPERwYPCHiTVU4VUA29K6HCCCMwpQLq+EB64srKuXWePqn4
WlmemErGCvus2LQ4KP26nKz+vAibKE9wVA5U41Xja+CKHYIqL4S50m4rCI+OAOGVT/sOLCHXMAgW
is5TAHU9tNyvX7Pzxf4BbIF7MgTfnkSbCEt4r+0RC7MZ6a3liUgB+u4EN/W6pxKIwdWThyOkn6aL
hwoXqnE0SphjeZs2r/dmS/SJ9vTbHaWcdc1CtEdah6B75Gkmyzw6eYoW54qjRKkUUoG1MBu5K3mh
K1gQrKZM/xB77SdvDjdMWnKEc4x4qq1KEzc9B/+rmEdc+ougo27NiseHhQU2gmGJ65rYkEraPgCc
YVrNhthwJRyZOuA+Fgx8i8Li6i2YYHLUzXYrQRFf44MCjoE1yuJPY2EEzqSxKAEP1wZVaopGghXj
J8qSoMx3amSVdqZGASVJYFNFzVmK3EYQDNlHknbB6KkEN2URvCAEHzvZRV6PZBN/I1xc8lFDwxWr
Z+dcp24S5/IYwF8BffKLbKTGcNjjEckGmCSft7uLdJTpxWhZ7wArV/ptAHatN0AazBp5YYa081r5
9pk7cyKSpiOstTbDTz+PlgytnMV2Vy3R0cVmq6jqQUXJQ1Iwx6WtW4ICBK0Bo0z8HTiz/5i1N3zf
vgxxKv8d63TbOVmK0nOXGNVQ8+s2r9seRb9N5w/N+ezHgC0xcuMQDw5eWOOLmd/gft1CIF6trD9s
B0K+K90BHDBpUgHMghUGrGICRfBvGontkC1hHZnpjs+jwUNxEXJ+cZmVuniGgUzoATDSobBsTIds
HXEGlQ3dJea2bC2gsPkus/R8wixmjHwmSYW48LBF0UrVZV6+y2xR2yyaF5Mp29ElePB870vplnw6
nOnnZrFvK4dzs4x4nsVRZ5tQbOT6nrs1yOODR+RNtc/yPhB7P+/o5WBneEAZeejGPX6sPxpu/F6T
bkjQPYunDs3N12Q6BEDluAW7NHV60hImBy8RTAMhCDUlFFpzX9azjjFVc755j+rwVLB0wr3S0A/B
A5H1AitwYbRuMpu4CW1r/3olnvWdDYsWjST0s/HLN67gX03+UyIWKiai/MmIzbeg8/srWTkfuxwK
ceObHsq2RhTd9xtc9uci98dNIkDHWS/JqCOARzchdrJI2N4qdl/iLYN0atKR9EGUPFJDO2G6GPu3
8gN/5uc1DvdzzwBnrzRf9y05gxWTlSXu7lkP2w7CFYaWST+MN7/LQ5yFANQfbFWmQQBqFVGAux+J
ITEYgOygyPapNxpzIceZaMFAmWm6fohtb8ZWMvgK5B4tbVasxHx/dEwZUy8GHBeR7gvMKrRG8r4r
pseXcxvFlXjx35SScKo1TwhhPmQtvS0q854/N4rPp+l1HeKs35z1NvzyBASYPiRXyd6irVURFrSE
Wm2OPdb6xI8U21bmZJ5JBJjTJtHlnNV5TtdqhA4Sc80DXw1INl30vTCLr011n7W9RoVVr7RZlfP9
6XEzWxC84pInZhk0el9g8K/XauiTAR4rYYba8YPFFDakcU73xJ5yk7JjFfS5PTRvsXA1mpmkb3L/
jtKVBmRe7F0e8+09SXXaZWoG5YfR7fOpMn6MSUckrObItyDiwxnn/SxrSEbhpfw+jsE5lnzDMYxe
2Liu46XADprq3JnWZKqW2h6i/eMaz4MoDJaP8x5/G04vYtbN3/lbYX1rhJFNmwcOGBf0bNzH/c4M
apHeCKCPpFS+7bCmnz9gdDXYGtoAm2zuOcv/upFpWUkikk/Xuftg+lA7yOCLNZq5WcQSS9kqDDZr
7uoBpPdVtXCnc+khgEg7JlJSSQVQ/XX1UjUF+F18c437DX7SnNO9BnOOrPLYVhXF7BxD+ela/Slj
jcodbLMhHtuf5BF3o0YpfgGwmk8maVSdySB2hjbkxY0bIZlLo0V0Mt99Q7nZ472LLICZzkd9AXpX
mbfMSrYJfhw4xdy37dgcnT3ByE8284acNmE+3xOasFbT95U0ve50CONCTeWdTjnE8xZgVBmIgPvq
IAVao9m+6z0Wnx9ShdA2lnx1iUIQlhr3bMOhM4DEdyhko/zgmdCcApx/+ueehXhf90QrjIpN7gGu
vtOjcrctySwrrV1wrW3Tp/FAYNzvdHHDKz1cs8eb0zK9YGbI5MVytx9iP5tavBTpdmb5kCpA/V/q
pSHKbGB8fa3qkA5/WCXQUZJ6XELp0K82r4wr5tyPKjKSZDUJpGJ5z4W5PBK9/ImcIB+EnVLd+x0Z
PRy9rUMmiSojJH38zKdHv5hDbygbAW58hlY/+qMtJTZtohX6/V4E341nUDf7bEJkIyzTexph9Brn
I1zUgQuM2xYIbjpLhujir0t96cCLCKpPQ9BfuK5kqYV743IOcM4mDB58vvG1XtlXy01e1bidARlA
FATAE7S2TZpbqpIafzr/5UAxsgLxsxoy0UCCyeUQYbcs1h8iHApDpl0WeP+a7leMhZ7CK5pX3qSt
rhX55FSXwXMsDRNWGhVwbPq1L082K2VKM1KQl56xWUjJo3f97SxLEgbatq9DO7nhN3XOGHdRJxfw
lwr38DymlazEuB7T2/zy/MnaMnQ4Ar9UMP80GvTnfEVO/HJ8HrkZ4wJ9r3Hj5tqgNijA+ujP+L5z
DzSaBC2lh0J1Ta00sZbwSnLXiDlXyYUTfNNCyhTtS3x99gVofnbPKWATQPJz72ZQbLfc+5snwMB4
7zrmJfqcKj3IrfAjwk6KcNulv1EzfDWns0ZmEaW7+QOeCTw+iJ6Ho6Z+6vQZ2gbWHP2X0X3PWnoi
pJTzN0XuBG6jIRJpauldqNIiXSisEEzybFY6Gl01gcLY7LSl3RnOqeY5m2nOTDJG5gmodiDMAV0R
LjNIyIHDqkMz7fQycOX9Ax/XcXnRKyGtERoLJejb72CbfxMs6ncgVy2ejOUIRTi6FsMpPqnWkHxo
ZhFKNFY1s5dGYZfREfaI9vBxGMayRvvvktcfxhJm5FONJ33+dvcfESD36qBlY0M2VOBsnRYsM8CD
YRLH2vpQtKvv6mzky9FkybQej+YLFzYWGSDAOK6q58b6Vw0XnM3giu6zrk8t958fxQ5RM0OY1Nrs
R/F02kqkA7OjchWrqfGEDlVswaWsLO+XiubXDr79LLk/a0AL4fd4MBpmdfW1m5x4uwS0VDMU7y2R
YoVk9VPNGV8CfVKpz/c1qIOD/Yj+NqjF1OL3H8jRpkJZpdrzYAlr77p9J9rb6jCOfUlHbsmpqglh
6mXZb+GoqSEfTw0Ef+DD+lNM0tkQ8cM9aOPTIs6UKMjINw1LE98NggE2MqHlv7BM463i5+th5+rG
1z11FEN8Wsm4iS9QSmf4I5kn1DeajXvWUaNE7KwH/wF7R5QterdOVBX9v2/Mp3mFP803Aj+07GW9
ujI33+LyWauABNkGIWd/o7OGBMda+xVvp7YXjhzFfl2fjy17iHFhaGJ3y2HoxOSybLRygcDlWt1a
MR1Ineboqc6B9qadWFEAqcnf7+rw1zThN0+ctEqqlI7paTuscKZcxqi1JtiXkS+HYPdhVIxqOPMH
eRo6nS85BvZXcSoH4j4T5FU41kcIeDNKTBeMMpXw5eNenZ9s/A9K1q40rIxpIZa/LKrfR0q2AGsy
tDxOuSBcwNywEQXS2gbhA2CuaJXBAQYmX3Izi5+IgMEHqVOMcSPOrfi+Y3a2AWr1R9q0s5tZwcrZ
VAySRb0Sj9Om02V2K7kX8wwP/tQxcAeD6Ycpxd4smGd9FpHOcFJVwhtEwoOFCyhCWneaq5pHyZ87
MTQTaUxXQuCqA2lihu8HDKLAXRDyt9fRXTeRW9bXvyUHFz1UwYJMUAxyb4TdlqCjMIZbfkdN/Ml3
ca627v9JZvFbB6iLiOEGV2kIdM8zQFYmo/RwY0Kb1zAAVVFibbrs3ULH6PUbW7Edl6ebXyxe4j6l
aRGDDb1X25fow+VRw39FpGD7e83eza62tDBa4lm/OLPU095V6PnAZMOL2Z/bR8reTXDZ8VKseMyM
sBV1ZkBVbjn6bW3v679IJCCV6q0mhF7//4jT6gFS6OQxnzTPaD/WoOmmGs6fG7JQcgwy3llRqdyl
6zhQJTAd8R8JZmW6wNUnk8C8zrJt1Lzi7XOmVsLRAnoALTGGUiVFZC39GMuqgDvpw3qtjFh72YPs
QLZ9gAC+yPVYtnSyjaCZUGv/7hXVf7GXy65Dzt3PIi0gwJHFpaCduV4o0C4EavXFmD8h/uZGzz7K
i6CLV4SmrQowIySrYe6FjsyRqHfYrYwIo7D6Kgui7jblK1rHIi4bpOUexQxmq4GL16+VQEUUk1+e
clK0lF7F+pFJ0LSXHioUhj2d3gM33RQCDzkWmX7mN5khXjKgH92qZaz1JZ/wfju5SVKSVc6/Uhsd
sqnwMblC2oL5yXb2bgAjVphaEkdxpimA7/k31099zkU080aUHW+QX+4vD47ZNpmzOaiQvCq4K2dZ
fuH4mcEBN8Za2lGt8zninRNJIq+XxvRSVygb+/xdJptjPu714rdl6SX4aSl6miHQ9dzY8qDEVGTK
WaEbxnuc739V2xcpFd5N2lZI8OWz/0HsylplTlSIbsNJ2IwcKn9ls2hLutXz41Vtlcpli91Z539H
je1YENAXI5nHgBuwxgVfAJOcq12CylIzIV+6pwC3X6G7+TI6vOPRFwaStrqGIl4MnalJ0FryZYbI
XsFf77xPVBJORAikVV3B31Q7WnlA16Tsgza7LL0cXH0o4WO8k9kYxWxjbnt1QxPF1p8QcrdhF+Q4
RE3F2RJCQi9dHGim5wwA2aAionQvEdASamUxeIDkXUpYMpCDyueKHIif/YGYSHYgyb2w3mp+sEkS
uICucsxrVX7R7T+1gxbwTYUS4lLW/N/xux9OjJrxs3gaoi1nUqQB7W6U1iSbff+H3fVNs0EbzNlS
BDFzrxXc+Ix1K6FxZLtCp3KCgVOCVlLrmAHY3/c7lA2dGEhAbwB7WbKeQddZe4EU9uE3bm/Llm44
TU05AAXHDd2+RNZeDOGbOH7vu93W/slOp4B0dJhV5gkm27WzXlvUSz7B0Mc42o674nxpfYXr0g99
dx2YG9+FOxvecOaJjoxaPaz73YD0cLnH/UK2caEtXtcQuGmf9Rj53ZOAwOF7w/LpfAOv0GArgtKe
BW5QmuvE8LBQK0hOJXKtVmF1QPpj83G20ouUypBrxNOyFtwGA8nj6JgBwH9quDzDPX0IdMMXDvBk
RVwBMhI87GDcb3l8KlvCbLeZk/BRDdOqcPuUedten84hTOXa7VknRNMQ3+pNFO9svKl/WE+9heIk
2/F53fBW7kL1uI5sm8JWoMJWKDBu7hmCXrJgTLX9VNnxdKwk8PYw7bMMSZw6SeINmdy38PII7+Jb
YJhvbuUz7zZjLN3WlDZiARSoTB8JJlKPnGcbV6MO9u4BMqTKKAmaQLOsXozB7WBoRFqZRJT9Ghhu
4Ki1UTRD/brw7oiKWYabuMJEuZXloLql6K5LHr8pWztQbGliA82DMAqhLOJeH8C9yPOSH2jiw8Pf
+yovkGY9WbWRszRFxTTEkHtKZchOHmHK2LfL3yTVVs1Ru9IGwjVPJog566S55IFdqQaS4aDwjKIj
z2JiuszTBIpgkiFYOcXK3OpVW1fdJ1bUJMlz29z2d2rLH6ogGCQvVycpLFmygCbUq8haxW7vmtpb
CsFiJsKSWMus0X+WGBy2nTPmWlmhtO/tkb5yAkOw4flECHDC7M/0YMiRAbofEJXjx+c6SI3zAEJv
yJUHabr6JPC4X44MWwOFD8GFOyMBirygSAwG7SqwV7JWBnp/GICjFssBlyGaob+7CuJiT0TP/ZRn
mrluCpn8WarykG48xstnJOqnkYe9794qEy1+0bD4Hn8aHO/SLssCqxyKWr9YGCqDDVgxTXsk5aiZ
06m6F4RZG9rU6s6GEec/HwIMFyYSpBFAUib/Rgc2nwGDAvoWywFBi0LgCJlggDEr5nCgmA6jtgIE
GsLALtAFWhFnz1uzINr8A+BkoN8WgEeQaOKtdpM8r8t1UrAFC74w4smm3OS3mdbFDGIoiyzP56Vw
NSvhjF7epdWAB8iLCQXvVebGGRSvOgUG+uMs6BW8E0vnfnXWyKedcjtxBLkpDhLxn6NkKRxyrkBK
NLN9nB2LM4Y3OBrE4dmGm+Ce4EVm4gO2vxVusOF8JNw5GGtnu9lRWb/oSiUK1iVRAu3YPzbVZsei
km0VtraEV/ecMejy4M6lXxt0VOYmLeRbNdUpj9Y/9fAzCeyznaDoVtlMjmrQ2XWsQBOMfXgS62Zg
zTAioJhDsaMnrFOfdqedugJjnQeULmEHiQzxhGZddEKKfMmPoiImOKLI+tLSfbLkI3rDYs5oHDtH
9FOMR1nxXP36YdWIFZD2FDBoH4BIfOEQGBJPc+02wPHnxW2pXo2RaYHWUw5ozR28vw/a55L8gbi1
WIdRenfUxkVe93x6WFu1jil1M54TiKTioN8wTs3g/EJJZa2YybXWu4GTiFyJkvbd2QXOXzllDWiJ
4EPmBRgRa6MpCxCNwb9jWssxk2cK75ixI6kjnSfQ4dRmcs74G8GKT+vFRdXWcL1ifCH5ybL2fo/3
ZKptoJ3vheQXfpblWgTTAzIok3Cg1OE4xGDsXkWL+vkrHTc6IPRTpczad5F3FubxkpexL5OW1NSh
LuvVt9wtHf9Yhm38/31P7xI3+hPCXik8lr04kW9nr26bm5yBn9sq25bIjePvxzc8bF5x2g0TElJR
P3wbiG6B0r8DPH9i1KHxW68JLT3HnlJ53LK+hLuOCjg62TILiGm4aHWXdINRQVmz9rDRJkPRPqs7
sxe+0502MUBsts+uDZ5YXqBbODkcdmtBZ/1vbwuwembhCr3+5nu4ka+76CvNVffWd3eumvs/7uCl
wEBwrBYCj6hukcxwNOwn/LdDJcGVjQtUFRLyoSPcK4dwiLV5Ysf6bxjeuUi5J24lGLll66COy99g
r2aBpcOxELYepE0W6dXi7/TSoDz6psFniJBgjhUhDu4V/5ZAYvTXRYpTRaORV4PjrSBNnyubB1vt
mNWtWlAf3RQAWpYuP9YMmJaXAr6wI4jbe8jlOTHmslY5WYHu9OYt+sCEGrERUJ93Ir4LIfW3TfZ/
Dg62xO0iY/7BjdN4lBmWGOJNyzIOHZ26n2icXP3ro8YNkgxIfOOrZ1MgT8EiJlu+QmNQ0nYEiWeR
1VdVSU/1C/qvWIgFt+LjhErcAx4KjNwblcnXtxks/1LcNh56PTwPAEl+UCI87eLXQkmJGY7xQ2eK
sY85gmS4YtAx6WVRwYZeF0NtXg3SgHWwRjL5ABmXJRQUxs40Gbjdxx4j602LZ4DjmkOmxr6bvXOl
rfVdnY6fobwuxbDpUwcDXgTuReKUuDKjGSTIfDhZJ0ZwCiqiEyNseZgOzBOBLm5C928l8lqvWYvF
FkdGKB+AG7iHzELn1iHdMmE2Qd5TTFkTwHeBUDQTYgNcrKMLwzfyb5VDCGriiHeE9kvnN4TaxQxN
Rbti55yNnpnfcp3uorItceSTwnOUNKSkI1msfk0/5B7H3oqA1l9x2wOiWGfhimc+i7GpV4ufTeaa
qCnbR+JUw5iM3vD9Q61SB7VIX1DZnSo6jWfEqEnCZhZmXrPSd6YN0si3vcsTdBDKoHj9DZpQi5Tb
b1bp4wF0T/J1eb0f3rPNNIinv4sIS+zs1eg/YTbByfM9FA+x4DA5/laksoQrVYuBXB1CORNr9X61
Gs3cp4IcPzduj+gdHwN9Hw5ym7eFT8pokYaR1OcXKSQ+ZheH/YXKd6xDVlzeQN+sOSCkeea9IJq0
dihbHEMpr93itUeRliEHofb3E0oxGR/Vf1bTdUwJEJUNmVUdeyAq93Su7IXhefC5F6yRO0SFhdmE
e6uspBS60H0t63Zx86IC+SLrzMTKd5yKMtL3Rou7hlVoWITKuZ0/uymu5SWCO9B/5Qt18V+Ky9RZ
uknZaPFixhmZSxoAeo3/zYILqbvmkm0VZpPlgsPx+0jPDc2RmUTx8+ECVDpikuBsrBLw/XroHIYk
UTzD34C/7JLfUpmijJgIcyieFDk+TXcPAI5FilJs0/0PiTy+1lcZpuA+Gtk8hpEVt2SshbEwQyYd
hFo4cYsgSSf+iMmd8C1xvQX13S0cYQ14ry7ewenpUiJ6TBl79kGGd+Zg3h5fLYfdZlT8l0SOvVEo
ay+8svlsj9C6EnD1hYH14H27dXllxt0UhuB8UQJhzYxudSceA0r6i1YJhe77azlMs2XzXnOXEQab
S3y/YoBnu8bjfe7VVyIiUj2zqDmAjfqYAMjv65HPHhsVL3AE/Efw51010whIh03H2PW6iPLG1n6z
JoChS/BjArrH0CWHudKT2LzKh2atg/+hnQntKMZqDBdDGSrVk+JKY0cIJWgDzF+im9xZLJV4DXjP
wg06P5+GObXSUANZ1/DlQEtn51q4ulTlDieIF6wVMUV/wl0VvX1hQofNZ99LQ9j8xwlO7kzjccEq
7G5HCNO5fF9x2Utmg0v9BZ2af325taZUgrdBO55wrVLysXfAO76/idFIPJrZhunYi5gzJ2Euv3SB
iUtMUUdhRbo2E4L+O0Z0eutzJ8XKKk+il2b4ZzE8H+BrrVHc9+DP3JNT5xVGQ2+ltgb56Ingadi9
hYz7dGFlOej7EZ7+SCnKvvINAOgd8or2t6nHXOiIAb66DQJyp1D2UJDIroNWkA68JdtPmSHAZEsi
xgBT5ANny2FnWGurWb73vB8OgrGHx7vTUc664Ek3hlwiIfe7OUSN1DABRpa2MqpIoMVZTl/NjOWI
PrQ9yQAeEXsMPgo6n0YPjvSrMtG5PbPg3BQvGDrbsJkzU6n6C/p3FOTO6sIUqGAt0yKLmLin4zgu
fvCL8PC66o9u+rLgaK7qxt99/fPBl9TVSLvd7xNKEY6PyDBdioUv5ANw5YovwB8BvSp0CAugOCaH
lWDFBeNJ6qQm+tHoc4xQKwVdAnIhEWQi15aAkOBH55ewLScUUnImkAXbJQ9yLTEsuZwL0ZBy2QYA
hfviiwXf/KUPkA99YDe9IiM1AXwVCCYF274r3JixRTV6z3kanTU2eA2N4bI4MSoDpLo+f0Et+0zl
j3QERWuXnsY0HlE3VwbAzrE8s6S8pnaS5DGkvTbup0XRXiMlYwzih7SNWEMH7Az68cckIdIhMoW5
XuZ/Lbthgehccb0bMj2lAHDMR+wGFxIof6CkU/N8DhhmvX5qQ+oW+9QzPO842FLnRWnMQ1GI7MM7
V5LDdhDr9TGf7DIWGRiN/fy01EYmcQFr61YM/xLTwV+eenL1XJn9OhGLxf2PTTWYqHZtFBEnzvl9
Uvlw5EkQiOgaOiTc9wMOOVIHqMLVL4683fgtJC2RuzoF6AW81jA5xMqXli/8p3/UWpSf+iTW5Q3v
uZ7MPTF3j03oqQdeepY9MiUbLNM7EadZJpQus37olRnp4H01t332b9Sh5zRGbUGxrXmtTej7PZcM
VvNNmAgcsgD49Nz3l9K9sw+VBxhsL+w+/3qg1jHd4jE3fDRlAbSmlrnsZdumu33jWbicxun3i3Ij
P9Ns+0s7leBLAQIuj2bEXLOF4pLnwJlHwIA+SmUT2kRcTtTCWknEuyxx1CzER1djJFdF/hz/5d2C
cLL7cbOXZrminJIm41Dm1A253K6mpc9YzMnxloch7ZPy/2A8VRMxntdGLgPEH1oqwniMZAQ5SDJl
H7e04GJcLKRzgMZoJvw7/CgyeQyDUKspILSH/f5OUo93QUe6rH0Qr7aRN5SzehtusSHjFLzR4+T7
+KHFqKeHayqN07GxMWnzd4CebqH1hh+mjV0a6SHxK6cAj4ZtaLdtRA/3tr7EJ/5NURD4Rou1URXn
E+OZgex996TRPa/iAwE3l0BzrwEUU2vzrDtfB/9Lr4JLXy8pttPN2Iy/rvFOZSAUwZuxUDsgDjTx
B8OEe/0Zkvf+CsnaA5bRDrMeEh3QbzxonL4668xaW0ULKt5YiEzVPVtwkrdN5FUSS1dtQmdAf28z
yaCPNlvUvaEVFPvmt8C2SlWVEqPTvqA0V2n54WnkRGodoEiySGsHjAl6+zEhykuOYz67Pm4fAGsu
MFFBrdw3nnULAd5lfZYJZpEQoegv/sCJEQnhwpGXOrS4RpeQcZMe4Za9+4ytx+r+F9STAqwu3e/H
SJWcJNY8R1yHQ5Ka1OCrv0e7bojsJoctMQ1kyyfJcHz47fI99r9qxptRMLg/rZ9xMsJGBMndUW2W
TJXRmKynQPbVguw1V85f0coTK2Ip4yYdcu2droaHM/Dh8CsBMX0CIK7Y2LJyB/5j/Mm/7ugMgpRO
5fkOPYaNqyrJNTYoBkmIu7+U9W1zlGno/0nMMgGTpIlZjr+bB2tKE/TXG7Zwf7yH4I2gkt6D6f5F
Yb5vx4SZcWj12AI+mstWFZCpy20srco2BErbKQJGPqOfYl236iDFGNQuedFQrpUNeJuQ/sSWtaao
WgXx3Zhaqie330QJqXWlO3nzOiDrB5n0NcVNBF/1VnH7P/Ox2HPZNnTdtEhTRApLkvyohSFz2hcn
0vj7Yq0zArkHvqu0hp5gTfmVDWVNd1CfE/60sHMCsL3sFFMe5KLQ5jX2qaolKCvgoWCBOXET7KxF
vonDjYT8yIon+VfOWDWM2frACpgv71elH0RxE6ysooLQxM4s2RqHtpPqKZpiafFcBas3GwbdjERj
bECO16z8cV95IDQTzy0CVU6Lj897sBc0wyERvzSz3tSkm6PbCuWyEd+GsFy6PVMVRO1iVRIDLPAV
7yy1pCnDToaV06/Yj5FiIxnUqWYUW8HmnfjJmsyqow4BT0P5/bsWjjyXIXA8eNzEfCjeMhprvpem
vxFU2MeKV09eAgDIh1LTKtkS8LgFWj3gbcrkDoIa1ZFWv3ZPPMyRdH35YbAJy2u61PkZog65E0xZ
6NM+Tjk1xpK2APKdy7nilL0LbzViWnsqw/0Ju9rVFeJqLZLNUSLYuyTfXRiWLUNlNTa7ZZ1XCZBH
+IEH/NX996UceIKvtpTm30AZtukYbix6syMVRBVAWi1Uclrl4XSYTvnE+QH4GDHjusfw67uzues4
SMGB75rmjQBFE2s6LyV9KZ3roEv/yaHolj9bbY4ufjHes4MblaJyzUmsovdWZAn2esggo+jkAkBk
GJEVbQriSvMg65jbSMCfaMNrPMpdzKVhcdpUrptx2G2/htmv2jlEN+c3qi0KMwiHsIovVi/slPkD
6x8oaCfn+mc59MiT3mLayGzuknAUAfBcz34e9uFqWfWFlYXGgwvV5OD2rX06rPUHj2AM2BEz8keB
yYLRAfzbR6TK+4LjjxIQUrKHXeH9GNeklvTJN0KL9O/HjwhzImYALObi28EonTTql9ZeR5TEnkTC
mPlR1hiVhWMwTUNBQziMTs4GBhzUmnSM6SYWVQgd0lfZx+14p3v2xxQaenoU7BtvVgCaWt5lPpul
7bo+pcvYGSB5H7sps5MrEWfl334N38wlrvqLWsDrvbsPMMeBHVCI0Fgv+yBd+wCASa/ExTUPAk65
BTjbbQ86diGGV4OZjNeLm6e184L9oAux0H+F60Qw+NXckiyWtl5UhFefIr/xsGPg6N+M9XUIqZZp
8a7k26DsgIbBmfghaCU6sTRmDXiP6HvfobwU0webPQScehKjeyAEq7RJiA3JZiHR7pox/NKwLtoU
zwPc5Un5WWLNgzTFWuPMHms9PcOS7Aa+/cjHVVZfeVSONAM4hVUmbJBrqqtKtyLbrpd/0/NFJg4V
GDjEK2GpkEEnCBgVnHY97zCn9K08QZVHavNqL9IqJEdjHiYMOl0pxbBeZEEJFhrsnGclUPZvuV37
NhUlJw3Brr9bhZ50PXvopfRTYzkzsGuwofyi/CfbuPxY6oNpDx3UJH/ArMK6mZBzqJCUxSAFMOWA
ukPAjGXmuRyWeK9r2stekg8l8aeMmHpeJxRb8TGvnx0dQ4+/uDmgkeGGIjsOb+hpGnoqwmdBxw2Q
iqjxxQAXU5GZLh39NGmEq8WNOWo9XR2cj0dZoIf/bJZbr5OUOpFGfaYnWlkuGEOAYWLdygKh/AjS
sF/X5Lurt6JsAo3nhuB9/eA46X/jNjZqZCpkltjv9XlE4I4EqwkFrCT0mIlc5ajF2Jc1HR840Fdj
hOEZ1rJamp/7TehJQa1nWn/Lv+7RgZNMgwx7BEDDy3l64rJXK1MaWa2IwGwuyzeIR0TVNR40xQB2
r43C0mSr3i2sSk93UGZ+f+kD8ZZTy/3p2lepHp85PQ7Y5DohHDw4UPrQHQyZhrNjKMt5FRJSgs+N
iWiHprEDNzsD3PmAC1Xt0mp1MPIkf8M4RJEdD2TmSThfeetHPOxJWJ4k1Io6QiWjyK5p45zkCxnw
oe3q/uRulUB5uqnjxD+g4tNofjR2aiEkpNwbIrEykoB93fpPzQnxAUItfdCcpPLEKpIUruIOhYIB
7xCwEchjDAZg39Ei1T8TfghdRhAvNcJ+fZ0GA7YYDPJcutwWOUy1rrm3pYfZ0p/PC2pV/D22WRZQ
Q0CdHB/tTgY6rQtorcBZ2D1UeTTCKve9tGVC/DVTaY8kEjQVEXdNPYz4ExHZaf6apojAEsFFMZPI
ySzq/akO/mBDFM4u+UxS+2UofouOo9t7edWQQ/l7KLT+pTEq7YvoGOxHyoRnQZuXou4uB+NuLQH9
EZneZId5rIAkhsglCV+m39ejfD3SWhiCvyo56KAq7hlIf5dlEDkDbTtW0YNEL/kd9GGDiWUVGWtS
PcGtuSheyBwmNHZNAul3HPC2ceS4wrjh9jjsHLje+6CTQpeyQCoioXGt6k7Xk/O0Y74qV4JvLXni
XqZWHI9WJQulI8Gs37MzitIxwIcYdafYF4WHjG1EfSDEo89/iAM4rjRXYd9rrjtRt8z7n/EopUNN
qOTwhrajPcmChSytMoknFgo8lJb1RB1lBrxajDYLG5O82anreIzZv2ETBtMue9yvN/TrLjoYWRos
lL9/gp4vM1OAvrjzVz8lYl4jvhTiODdhbnSDmaGGvC8AW4r6RIKn4sas/rDL4mR0yuchi6YpmYS/
DocWBrrM9p/MhK9NuDiYoZdQFD3xYLUyW0Yq4YtemCEUrIGtg0MzKGX+pc5fdGlByeOKq1m2hnNm
ZDcwj5euhSOF6SntWhIYu9nvao5LcjAC0I1ThZS6AyMUph8pOzVZuPGaswT6lSY7qLL9rVjRcaip
ZKCQLOPeZTmxe5a9holMB/5QjNg4a6VrE3JZQ8xT6j66C5lQoEMfVctg61QEFp2Lq+3XhpbPzjjZ
0DtRvkPxaoIV/9TuDwEQzvCR0d3Kcza3JNMeWzV483aJvId9N4+ZL6aFPQlbYFt+Ow7YS4zjmHSu
vK6V2oryYi/cZa54eHTBQhLZpmbVl3X9Vr18DbJtVJ0Huz9kFqfnSWK93LEtLh1qi2YRVeh5l8S9
tJWF7ljrkjKasaejWkX7xOGQ8MdJAX8ju8JYr+o4M04K8hhU/1qpBc835HB3H0afJMwTRAxybITC
ad+o4mvmva9Y49bkpZ4zW1ATrWZNF9q4VAsXlZo9/qQ+aykgCfjajibA8ZJ5m0YGKFZfK8Xnyv/r
iWInI89jmPtKIZyIL0jce3j5LTI/l6Rkute9Z5DkX0r1B53DZTenDbt48JOZQsoqOrO1yRae0lIf
fVzR+bEaEzvx0cquXxEnWt1YWHnlJFmhu7Hp9hM36WO9Szz1hf7qSXHKENLq6wVbFMbU4ikDW/5o
nIj3gIFCS86+nUg/4nxb7v++7J9xZNOnYMGJFNYfR6IiwrGGCcRyJP8pX2g8H89pkztGuQTSOEpe
S/HVO4uE88xdy4rdnqBRf2md2c0VXX7TNNrLkiuOpw4ZhzN2RAoemnHArQ6mGjUIXZM6k69xHL9x
uMwAR7EUsCn+6aAxVeCmnFSY4bZZP876KhP9tjwBoMAqKnXWy9uMDjg9R1zlllSKs4CVMMdNYG3m
knygrz7VIjHvYzzzWs2AFS7GtFtt8l+2FeC9lEuz86kgKGVmiUjx6Wo2r7+DHlvJ9iGzi+WJUVZw
c7XUSkeLd57SRLf6pA2Yu4hnt3SSJb67es8o5/N2E/Uo2vlgD7o1YICeTpK8OhrclTEPM0HGaLwh
eZTtcXW9LKwJULEQ3F3qrN1DMvdfF+CLWDtAimzlcAcB/NemYNb0k5RvfetQXfXDE9EsBbutwgDw
8xWeibyz2DHWVc36YsFVckhTTzMFSqkkJ0CmJ9Sk84vwC2NzjJeBOPypW6PotCmcXh686Cx5lg+i
tZFs7qA/oRbDt4doaoYw2P3uor86/uAysQqSrUv+FAvQ5DqD/6lNHDV9FOp3332J4ciby9hoY0I7
t9kJD0DOZC4f+sexKi1PkQKPdHslVdQMUyWydMIUgos7akrz6jnjRaN/g0JXbrKaQS3Dn2RGKiTd
CSIqJA6pcHbg2JPskTB+1ClOC5EBQfRIrjca1vNRkOUwAv30uZc6EQIjlrtaxQbf3ez2WCcIOQyp
RBsLIBBICXRlJ2ZxP9EYJc1t8dgsAc7WcyESzM5XLXMlxHed4Z8KETnnrqFgcHnSJ0mB/0ai1rt5
iU14wcdX91uLB6/DjvdbXGPUis9W9+Eqg0YfvfgeDBV3rHK3PwF1JdjwtwU/60rdFGS0+ERFSqc9
Vk6pq63IFsEDphIKOvtzgXzU7ItI4rhcm2CXbo0UKheO3i8d28AqBmAXNj7WqObMOAbLGmEaCPRK
+ojmBuLL7M5goK09AYWqQt7W+gKiS8C1TzTsfnOWKEUVPNH8BCtq6zOjV8u+lkjITdtrbQZp9ade
XcW51SvQzkYFWHeXwZjQ8lQrP6n7Nint9x1XgmXpYS9MDHoE/Nm0+kFwbiGPHy4HKxRLgJXqTmKL
tb2ef94ID4BvZkJIBzBV9v0xsFmIJsdmBIj3I1Zxf7gg9sL+viet8RTiTXhEjaxEfJYYWi1RPA6x
UY+MKShvJUmsGo/yOttXTFQN2F1iyhqM1AiQ/aZqgcciIZ9wV+DWZaIAKh7go0IOv8Gq+Bp895uw
ZM0ksuXSywOQPfKLIk4XnKq5MoyWgu1bVcf+mmXXuz9z22uVdSGrxuzdcvZDjRYcdEtIGznc86TJ
JTcka/BEjR7zFAL8rsbwXVvmQw2ncH2bKmAot7SY64pPH5p+cqFXqSR1KNooWlMw6hgWO0TRTW3F
VmYyaYOr4tIHmrDAnMRUwWJgXrjee5WGhEhjhAVagIe5Mzp5Qbizciw0It7mat0PCDAW/8+GMWb6
rfqYDnG3T92PdPQL4LW10sSHwAXoG86Wma/CF+HOHTzLH3r0HQ/ShiARbJfEftRI9pGin359GarA
YMpxWs5xXIhXVHUT7dvQ3LVc7TBlLqeInow4yzfU5/ZoEOGItJ2D6+EejCZUPWC3IG7R6IOlPlzS
ueDix5iKzKjv+GvxQp09WyyWoU5E6KR6750WJTqdOGlr/GAmDH38LT94HMT75Q85HlBzCEvsBGWa
aIF1+B0e4Y6iwlTtEzOyX8uqkdKUgMTFFI2u9jQEJeyXBfVCompS+LWUc8wh9Fq3X+W1RaECGfDF
/lRoeG895cQw9u6cnU4/mIoipy9G02ov/uWiufj35DrNAAdEN7o4/lydaUpIJsphuhY26S2Am4qM
iCSCT3/gBsStvOxduAQhP2ayIesj6WcYyU1K0qIcbn9paJ1nwBsNpn8AjrJNBZ5ypPhIgFIIvO/l
mFCz8dHkZKHhsbbWdsfXA/5nxmPAK6UXr83P5sMO7/SqInx2+izM6+0/NMxeFKJhRzARV/0oPtmW
HA8gQYB70gduNgJskNJgcPcOASVNqaE7vFRysLYHvL2b1BI65A0oqC5JbZXGfAFro9AfI5Eq+jFl
gwWG2n+2MYix2RwvUgcD8AjWrpygl3wKgGz9cZLkpYy8Pf29ELWbv2qx66YA30scm5YUOnGT9amc
tcWQDgfsBx6V6R2b/39semoWbcqN9KW51quR6CGD33eTb2gTEKGdWEdOncDvcieycrdxcUVcpyEm
rPxBSCWTtoqIU1eTaA/wfZtKhO8CLZw5Jod0D6s7jhTYdLVp009HhQpDOukVKTRWpu1AOz9R8A/f
NHuw5UQZ3mW8Y6ekhe52gOQFIWtubhFulgeVKcmak/Z262uzR11xMjF65wqKbwj7SGb4OmyubTBE
G6T4SjXxdxONQJtyFiFZTnWAp1KTTrhiDgGweFih1g92C+5aKcJRTh2BBQzjkMjdVSAYdHUsOXRH
v/sudEVKTcdQ9BKM8VUG0tLR/P9AEap25hMyFIwcGv2fR0bDU5mVP6Af5SfsoWVU4JVxlFF1lfh2
tYhI52vff6DzCJvCLt2oIrro8RnEVG+R7Rs+BqvFt0W7SmD2ki3cWALgEGnSqRuCD5Rc59lBP7bV
3ZFW9wAQacaPw0OZJQxkIV6BGQ3AX3+4L9xnEUDxJaDSIRogcXU1BLbsq8XeY1im8s+TndPCVs2M
rx4NULHcRb1cKO3J69ccJ7jV+OV4Ecn0jbkT9NIMuRiIJAwl+qV8BZyO5U89mkY8CqHYNPgNHWDM
Y7kSRTKyPTj+XAPqmouyiNVD+GphYkIwqR1SWfQVS5EYZA74zman2OAmKiWci3IQQVAVCQFEN4Dd
iAnf7ZrLHIJj7GWnKW3FJnMqwCttVGfuWCNtj47AKnryVOjgXUTeqX0hPB1izMHXGIOQLyd5yMrR
hfrMMfEc6ht3Ts/uUKOzb2V+eDWLz88YOfcnJbst0kZ2yBBA22tvrDPUvaL7LL37NxyvudhNZehg
Lyn73miL6kaA2TxDOTFi4vfibDd3Rg9EkrjoBUpyJo0fIW8vjvd4yFoIt29LKKS+06HODwQv7pt0
zes8mplKk58iDq7sM/DrTQXT7OAsE4JVI3hzpxRJc5Mi5BLCy3we6i3qDEN8xTO7XCakSstQnkmd
UW0AuqRut9+rknnYv7VmBfkyvDAhIJpFmQuMgWvukZL/b0+2jH0vh3BKuzsz2g4vv+hwPmx821tg
/nmPX5Hw5hr0uVusyH8Oh8mr2RSlbE+0mJPbVDyzxM+enQrg48zdGFePiWGQ03J89uh1MykkekrT
IUmPNLqQ/sI6D/HzMp+gt7rgnc1YilFCwLesWwEte963WQwV/47P72PSJuKknPIHVYgKiyHZE6Zb
ErJ2s0BSv8JQz4f02xLuavoBixShj994it0Q+5TpoCkb4ju07/MJIxk1bRPqvyAN88/5hi/vDLS4
q2aa4VDCu5tKkVK41EPTivafqe74h2q9JoJFs89xF3hsOIprjYCRocDjQWjMVdMloIxM2HhO+zRm
GtcwYP1Jc/2BroJsmZrIuB3JYq9+QrCRc1AA7tcB9quxpI+gOZ6y2KdwX8nskFhQEwtvEx0vVAsq
LM/poDCL1S6yyVcqP3gzrNpAk9x7o2xspju22MglCft11UJ+PaooJIeTZGrz2ZXkdcMDkO2YR53b
n4BVBZTLGZGLD0Tw9c5hQ/FVMfDgpLLQaw2t4MWltgR8m6sFcUMaXQSKgzHlQKrgMoy6ungTKalK
LHeRvzVnzspfd8wCcThzWpMzQZ3E33OF5liSZflMHasZnljuK1rexYSak9MQ7tgCVwcT3T/pxJsK
lxt+FztYeca1nCK4ucxQb41MohlaadLHhQcc4rWx0ittLiFfEgF6z+kGikklwDgfcLq1Xwr+q2ee
9UX2R3ZXXbI7jKhu+nBF661kSQyHk7ul0BrHwVvCwm3106WzdiLJlp7eMXbhZ302S2G7zMFNlQAU
ijVrKs8wz5Juv29JLLa+UfpL0HRzKCuIzxlFl7UCcUjM0NFFoNFkP4gNT5dSVPJp3K+63DkK++2j
Qhi7IeJbC1ePKtwBLrD5zAZtGth6m3cLdGl2FrlSYbYbrAZhGL77FSclu3Qc9fteSPJS3EUJzw87
laTTvs6yWxXwUBbVp6vc3kw8fEawrJddojiPPsA6CxlCQmcfrPI5gPPDmhv1jAszRyTOw6TvlfDj
HT0YKY6NE/5xCkfINpY81cXZ/mOEWy/dWf1vdYACrTMudJGW1X0y128V7mT7ojdQ1A4/PBdG8tdJ
NzoY2bLpmcExuaSX9RKkpxxLFaWxTg/1PvIQSLj4puDWAcTa5oJiVr/an1ZfxwwnBI5nQgKfK+4J
iE24xZWYdO6q1wZbZvnP5vQnrVWD185/X5fPhzoKoJI+sdCieZNHRaqLf3T3PxaMlNC4APJdcIg9
Uqiherx8wA/ZXKLZ0+gpCyf3kHEICrH4lZMBdLWry4yLgTQngo82kE8jilrTSAJIlnwuPYfkdGbS
/6oinoXs2ASQo+4TtTmFVMSIOn+ROY5nOjSGnXVUvjQhvkR1gk7gUHDgbEuRrbIghPLRE6u+JHZu
BF/DhDWPF6nmemq8lDEnbcHfFOszYnewkZZCZhUQ7MQVTToiir7i+5rXxFt9KwzZFlsusL8UTXQl
EF29+Fio1xJJvM4qLlMbYo9esVKSdXNPcKHW3J6emO3KMOVydljKhpvOYzpo0nNQY/NRbU+Gy3AO
wd4fApyaWNcPk2IH2LM0pizSoKxx1sy0W+5IIfzIFdFGHuslpT1OHSwkRtryTFAT6ie0duUGuJRp
Xxk0waQn/dS1fcqpk+95DNp46uqtJRoErnJXjfcvPs+uNaMvTUT+QdZ/4XaJWw4BUsnW5pexh0dz
xGglVpKkGP+S62q3KbscQkJoCB/Pp8/djHNNp8kmWvxf8D6REAXZBSmP0Nx2sePwfnkSSMKFhY45
RKSQrYSY7cutT0tzyAw7qHAK4q8LCHc7bh2giNFAhn//zzlnp0U30HRcyLEzHcdWAW+sIfQ744hW
JnCP8qN0wI+Sf/YsvvkFFwaRQg5RLuByJVr7/gGNmsR4+wHLn4f3k6Cue/gt99Jb7V7FTyZaKKu0
aA4TCwNIpyvBWbwSGoY7OZEXuehu6oBRjUDM4PFmzmhNNV3PnYiK+JvDU1IwdI1/xhum54ukajdP
sH1jFAP3bH5Noyda2f2CesAcufpbrzTzKHeTcinHj1X4EUNaPQB0lK7MNnrFvkoOYnYCQ0BTlaIM
yiaQkX6jDDWhtMoi3OqFxduPXcA2ZhHWnVl/Oe+8ZJeWd4Cm9cuKGV67e0T4Jh1rNLgtXRCCyr+Z
dC1RQ/fXlmkGMYWmm+0zkKXgrfdXW8AagWd3ISzKCI1OnfXz/CnIZZozSJ3mcexGtK2RTYq+58ZA
pO2rBIK0r1BIFQOZLHDX13zWSq+z0v2CBkBlUx0eymGyfHia2w66smA9dtCFeXGSzTl3Bg9p+Ann
6JhDK7nI8LB+JGVTSzcFUzcBEq9pJSXMHhOdIHb2QydwIw9X0aX6OMO5/Vfk7FNtdmcR6v7lgukp
htS33W5g7l2RbAg33uvQvcJzxZfB0adTU31rWeM3IrL/pQveEMO+6w/Hm3Nk3ti0/SlCJuHG+fpI
Cp/2g1H9YnPj9X3hF88nnBo3TOO1cJ0ZTy0mYevfDcgOu/ZT2rX81QyIgI5LLwYpxKOEjc6/H4vN
26J0H3WO75JixXLqHnayJ/vRRxbPC8DHfNt5pIk8MRDxxPq9JywL6Iahin3XVgelalpmtWteMhyQ
SoVF1dQ7HG/W+o4t9hCMGn8b/9wJbTigv6fI8mYsaMn9y5UJjYIjbtZOJi9l+wQoKzICPAy+FhVw
9ysfqCfN0w5aiXrX2XfMiMuo+By1NwHGoRs97+5GwsDVBVUL4iR1lZY/7RJf3Xge1UQoVfdYmN86
TKLoB2dx2GX0WYLFDxbn5bPIZQFZseFJ9vMrmKsoALax+lznD2ZmS1GrwIPOX2SgAI6/u9qINPd8
cB/4IfQPET6A0LFAoWjWpcM6eQaS+bLFQNQKy2SilJP73dZxWtD3NLaQZPQK5wGCc7KzYGVv3bHT
gN+HTLT7d/pwwbLz2JyWOCIUCu3WHnlm2zFvPVVdtUJgqpVSsmNdZoK4VD8OC783T5T1K+E8s9lD
M+nxBDu7w5lKDDaNP7NLjaY+zMOxHn8OtWJI9aKONQMlZyR7iemQojXsiPhTG9thQ3NXK1UN9Nmz
nI7LIpAftQ0ogvAs3RBHL8zA2pmGFmIVwCiwluMW/l21exv+8vmT5KfNgkmGWW3bSEcOVdW9LGFj
mMF/zdqEVLq5KSxbsJITY0wmnzxKeKhHJBdLplA3C22oZl1lauChQEr3Lpuq6YACHxDu7EPaK+PP
Jj4wkTwNkX+Zu4bxKNSSMNHMhm+kUZyGT1q73H6yYrq8slLElvKl26ZRG9QOdz2IFDxt1FjwZd1O
6g76NjvSrQUV0dFno4VZt2MNgjBD+1n+t1jBuZWtFlaffO6WsLRcNKxX+YwRQeWTS86V4nNObQwf
ijVzSAN9eS6bBJYAQGp4orNZl8Fr3NIWFF9HaJEE1eMNfgjtQL7LFCO+PqHxexX7YyZX94dvc3II
YWFj/7TDK/gmePFohqQuGAcWtA2yOrSVXewUkucnJN+bCvpAS9xNeQIDhf3nlGx6y91gMN0uxsdq
+cUoLqwX00yxsbh16FqjlQ5sfRMKT1vGR7luCMZ6jjvy46ZtXw7kwG0iSzBXwFsX1xAIQUOqctIr
wfDuQAT3UiIrUS77Z+TQnfUIL2LFjW35r+IOmPUc+h7noGWurTYSCHXlkKw4zlKGi/x9X05OgtAs
qEcj8u7g5KAnWyJE2dZiyn1Y2ZTde5y8g2gbhwlNaXxYADN2d9DKcs7l8KHykMuvQdRiwzgT5iiq
vQ3n8O0uOIfrMnzDOQKfzk3Lrqa7GvkW4FAmPIzU5SD4Scoz/wY996NCvs+JHnLSfRmdIrQnRNtf
t5vvRCQ4JizQOtadYQmt0AUfQIJQ/zU0oKcv6TNI6TFbEb9UTmg6kq7iA05exSFqusLzKma1M76V
gJ+LtW8Mc/opEdcN4xQX0WCeS4DvMVBNsXp5Nj7BHqxwsikDbTB3TZ+dq0L738CGahfQKWhKBKtK
SgpbR4fLDW5Dn1MOQqW4KyarJXDXZ3rT9U3+pJ/UQlHHEywcPAtsfJ9wVTYZZYltjctndLWf62Bz
igwGhaFce7slG+0H3BMynsXobSAQvJj+A6oTBejSRRg+v9rspQN9VY5lcty52c4QUQ8nsWG4J6RM
YejoTpM5qhXJx5vnUi95W4YrS+wfi7asjIbKTtc7e5MCN3wyKuBvbZ0qNoF/wJz4oTewCnQZOrZ6
JssJzv010gdrg3M+YAJ6uUqSwTh2DbY86v/jbyoN4CoSUp2Sm4WmuSY4FGMLwubOx2bV3N4c3R9c
GcVPoy+uU4bDX+FR23syQfXLbZXA5EjozhpDFmIBMJK9znquZn4JZ6hOC6Gles4Xl1RvxZD5Hk3Z
SPKi9SbxtIyJGVad1IVQ3CqP2pzx+AuGpRg84+EyS0V6J6eaivfMhne0mbOMYI1sxru8qCCeaxyR
KLYHR+P/CtxFjwjmBRgJtAvX3elk6aI8Rt2/TcFWPegPLxrbR/sorWlfQqb7q5g3r+0TFJgDjcE5
tHCk+kgVtxduVAPdEQwHC64i23Ifwsyz1n3qRUgmAJP2KROV624b04hfQOmkhLC8BMcx/Zcc2pYO
Z7yDFEW8xzF7S6KWcJhukyL3AyEmAq5dx2qJV3Z6UfMidshsb2neA5hY12Y3DDf+TOkCxmAQ/9et
bsvMVteTbRyXcdc8izC1r0j+4wcc7rz6s0/LU//IhrO/iS/HEJ/U70scMaQ2sKXGRYvAZTKvzSJv
Nw+lHjZCYUps6UGYK2YJvg8nVWr9r4t6yBDxtR2ladtplixR+N21rg+69Ys8cMvvSWbsBSvnQ725
mz2p7k3+fXQcfMXaIxjD2Ze/vxMsj+WE52gFXYgYb5sQkiut2u3+Ja9MXpwc2YXPvvQoXHNPMvTb
uzLRO7hWTbi+DaTA6ieQlhoed2EOZ46J95Qmy4FGG1af3gFpOrBubdhrM66c0cOzSyo1Ahs2KpJW
zAJ3URAf7V1kwgkmp0UQMPH2dOnxPy5MIj2gNNMOHt2hUnwg2UQDiIv1+3eA8gfxlR9cceC6RpcJ
7KEMU4vuINcYHW17G24uJUslbEfLGRAzjAbeEV0glw7rsKG2NljSVyvnXNClHoC7NTTlf/BiibxG
o8fKtAG7bE2rEYxdbelvr55/NLkHHpH9WFKnrPWG57bmR6f0fJbc1zB30vR+k71g3Pg6FKBgKUTL
DE12DWiCVpPGA+cq01oLkuzctaxCicg8LpvE+PjcDICvaqfaPyWC7YayPYyteF6Lmjw44CL2Cxyc
aXY8WG1blyV0xKY8Eae9uT//lHO6QSIcfQdRvFxTFvAJb7zjviuj3ZySN9bsTjPdjKZ9X8IhoMvM
l+pZRCybc5/MlS7ZZAfniXoM9zmtscrmO9deRoLlWPSl17EAKxWigD8bLBN9En7HsY9j0KV9vxiG
nVA2kjsfAKOCsiDi1w72733RRyoFBYykJxehRwspLLBKIrXuUtDrFv/P3TRaooEWbIJmyCtc2oda
P6i6rXkl4sfcTClyggibtIZmF50D5pHhWaEuRRbUgeKIgM8LG4g1Vgm8IQpXJVuHXzqj9TMpiEzD
0VH5Jvuo6bLUPVh0o3DTv/ZoRaMJ8O/a9Xj2aboBDWOsqlX+NLQHCUsNzAh+4WWKtZEKpJphr1oq
UTQsgL72SjKmY4AucqRGTKXFBrvfM+Cu6j+UxNff/huEQtUaCvyjncuFXu+GzJP2AH5Du5p9GYTw
nBx6leME4HLaPVYgd6mj2hnqL2jFlY49pvSkRVpf9+YqCoYPYkg+l/jtHbz3EMkqn3Q2G8yab+oA
4pbsfDzrkEwr+u8m6BlZD9yJXQZrptn0ttyi+SE8crlssOQk85823ejJyDctbp0q71VHqS0/+Aj9
cAHv0uaOJbbxwsA5z7vGKiZDDTFuXXEDTyrje9JtQVEN7dGWZrrKo7DJ8nS2ldzq9F/rgMMO5FVR
YR9ETMx+FKzAcg9aOFCgRQYXMUo3SNHRxKOULRQASUyu9MnwZ2tRrq75dHrXHRqzLsCJBJURk0MK
/D6TFIt8yOn5k5H1/bgid484C4e7hDebkXnXbDzxjMSq8AF1TpKiRqigDaXTgcIfS5KjcsBi5/B3
soyNiOQM+4yeCpxRk9OWye5D/+LX7Yt5B7aJ3PrkLXFVTKXNRrkvPfavl3r/Gtk34jeTaiqBkZg1
8TrBYHjl7kUrGMkLgLm+8OEAHvBFwnxL0TRVbUBA+ctlUSfuhH7wmETvnPTyGEw8ZF07BSXYWbDU
dWN1He2hkRwp9ssfCP19S2WrFVfm+cHy9jMI02SGlABwyvns+Us4XXsZrXx8ldOm4c/Y9y5TCkAW
CMBZFVDT/xGJqk5yZ8yYslhZhCvJXMSYmxs2H3j2JmqKX9MOHvGZ6NNw2BQeqnP8ektvDswvlbxa
MlTje8JSHIeLwqU7gtHhr+WYYj8HHMC7YvOqVBcRs94z68L7lKPZs8brLnu3MOGE05G/79KfqMnP
Da0k11iVkeTfLsAqoyuPsO75arPRkQoV1YtoHDj54j7EVx9UcHJfazqb7zSAanLaJoswfqq1kRw7
04S8fePX3MA4bozZukB1RuamoUrd0BSWRhqrqMPAU57aXTp/lrvZJLVPcu1CQgu0WaN9iIqhM/Gq
CKpXp5cA0P6Pjn/21b+CjpBRknHWUI8ovqQ4IGpX6Yg2rLxuNTmetDIf0gDej/6NLilIoQbGNQJm
bCcZtMJyUrg/JVgy13HLyX18BeXWfVYKZX0BAIfZu6Tqb2OTuLAuhDLqVqCOdt2gvapGQkrKmV4m
3moRI8QqxMXtBJ4w4MVArXf4NKsTryOijOtUDbhqlc4K/1aOdeVJtsdXJQ3AtYpVY15oj/TtL2lE
y77amufI8JbUkBY//yfeIjTYs7pMK09kafZc35dSNDfaPC2aCmBkqPRHXo/WJkqQnU7ESRZRtPYS
5hwBe7dv82odMWTPjQFmKKWrprUasDo5oEwQPbYqEZxerTcfB8TlF0zxvJHeqGdZ17Az4lLkflJY
5jWLqyWQl3Es0r9brUwUVZuWwt8XzPdtM2mpWCyVSa8TRIWUyJ/1cyaXBl/J3dMTGlDci9wulgB7
ESNp9t37hiLKOGS+iDM794Mu0sg5pmKUHROgQyrt9Qq34/gghp6RmXFBuX7RQVQ/oHzRQ92hzeuZ
E7qVhTFrusDFrHvoZgdOiJHcIYF/C9NwZ4i21w+CJjG3eMGAT+Tl7UFoRIowySkpZ0lv7W4DBPDC
JGKPhXF3HG58UI675Bw1FK4tpfaql0t4Qb8vBCHft81/qQN4VxJxRmSPMMdgiDIeAKE7TiNbZrGE
OdkQq8kS7Fo7Qq34oYvOx65XgKD3vFWU745cxG/KEA4zsZ/NmVFv+jvLKvRe+lxMPw3XqDZLJbIi
tXHDm1Vdy4vgxKUOB/dDgtpD2ZEv8uDXuI94kQ8B0blOFDMKY6k+L4rrYduOCITdNNkkdpZ7hf+O
oFNDhszz8DxvfDxSUAZp4fszPaA+IrnKvJyWIOrc2QAPFUG1U7SnLJ41U/5R0dcJw74VLWJeJxy6
maqMPICNHHdWBNNgy8YUAXOWuozEZWjyER6yLz6tcnqepOhZ9PoiA0TN7jMOPIYbXNHwjV9pQYl6
m/o92Li8VYi50173Lnx9IgB7d1q0Dwv7ohLN7f2wcds6FJSM6z0ET8syRk4Glk5ShEWH6XjO/7Zz
cBsEZX/SxJa1ehrnu3p90MxLHsvvWeDMsWl2EmS06AllTB+JYKY5z7mnmJn5TCd8b/UyfCvZAXtd
H7h/GCEv6gI05Jx2sFEhRiqO/9huVriscUJfhP7Teokk/xqQ7bZL80hbMQAP0ICYcxYUvLCjTvGN
c3bFFDvy+WYdGs4V3erqHk6OyK+8XV+ARtYeEz4RnTVCcQi9cQlEcaFwJgi4sFugUGQJ5ZKcLLq3
NUDHS7XvJHiGf2gBXjw+wPxs5kqY8JytocYA7nW14vLfvaw9wNF0aDD/RiCF6RWD70nfdDMxdOIv
u54kKWzHc+hPUZ21a3Rfc1Z/QkqEp20v6ldnZTu1a14fezOcc816B1/qHGehyEOd+YPMW1YggGSS
p9xFyl627mb2VnfBSIYfw5Z7B5lGZhMhiY7+CsGNhgsSUK9rnVrZC57NjxcY1nN3oywBa8pMvYzY
8ghNjHEcLONx659WqVlKmKWApOqVehWloH8zqhlbrzUgev4uiy7Km71hs8k3+LAZ5FqGJZ2wLti/
gX0mE/JM6hZNTyqFpUwvQIVkNIhQD5RxZzxU9hz49PpdDGGlBozuiUXOnvKRCrfgwjeB89GjLGRg
9BBL8QXDzdq3r+rVuJl6TjuBQnOijNQy4+b3S+cSNnjY3PxWuel1Jneg+Dk8+BqvpL34GHlJgVmx
s1XxXM2yT2t/rgy1Lub5Cik9p9+E+fQdwKI5jiZtg2FZ2uoy1FoXyxiX+n6RzKQRasREZLxKXYb4
CPTdpHsDCU7Pc0SngIyRdWhmwhJMpZj63aLTGt8vDq1jXSonQLtOqcBqacRoFYdl6GMLL6jE47UD
eYsaujPUb/NaexkSrk+oELC8PHJUQboAC1WuI93ELcspfbCwGpdPFncXxkZiwo8FcfLIUuQtSibR
adqei4z+THOL2DBcIPJaYzE0AhLm81DCzE3T8l51DYrDe/ncecwga/edOnhuxObf5t+ZDROJR3wu
kNwXvT7/QcY22imvh+qlIAywnC6jvXZo5Zy9+GwnTnGHKxORFwqoDeaHWRwDx/x3pmXSUtMi7z2I
jbkmBmpK5L3ZBQW+jE3uxU5TuUDrsRTH84XzaHv+olnBedIUU44rtdx/DNFrSXeYSMLfWGpaGkIb
mkej8O+q1GqWtyjSCV9Qie08oQC6pYGGyAGwyRJjeLHf+LgWjUrb5pgTXj47Yeg8yM/cnTFH5hpd
P+og9YDkkHF89uyJzW6gCCUSWhDnm9Ur1mAcB+w06FsZ1TD3/cmVTf6kKZViD4upxeS5mbbSZyWa
Lw+bAwPeTC6wdP4vC/GXNXbneqZPy4malzJdbBmOOKJqO3THjLDJ+vdbY6KDp74CwnUs6qnV+2CZ
lfiI3Kf7ejVSefEgJk9Lh2yZ8AU+Jt8/dHfrXhQSbT36FJ5DbFTPJwCAJV/yP+RWgBXdsDe/fkBz
AEk62eo0aiCfxl6jUUpX2kQsbcteCupfMhmGlrkiUcgm6sIytgbj0yx+Glp7Lk5zuiC3MO4v7Dde
BcjTUw59Z8V6qe9gQ7nHtIk1B4JzTfo1FeNJsNa59GrpZAlmxPoLc+pD8rgH0sE0Sh0mAbmpYyJL
RL2GPhNAKaAMNncHkTt58yfxoLgyeKuJSt9zGo7q025IgDgoxD9Xbbpp9u2jaYUS4rZTyakfZqjb
r+x/mfGNela2UlHe1cqBa3bk+EN7vs9OvBImU1zbu7m3vzMCV5Oy+OuzR5e+GT68026QUpBGEXLT
YX8blNOUINJ4Xut0+JxQUOKnqJyH7KcTSAA78S7Wpw2aQwyEyGhbXbGpQC+eq1md1ciR5pAIFzWP
nU1sIHZGjnNGkm8e5mlyUvnH5KVwbkvK4nxqDlZ1f2Kdxs2w1nDobwexiBehftCF6a8o2Th0knoC
nW1LpsgmfU91qZ9r1Ur6hoSR9Ie98IbUSL1om4u+oG8L1dF8ppwKISJbFJ+r1VhnJ9gPYB8lSrbb
TtgqbcM4yABoLQqLuWUTM7Uh4LWzZrq5pl2CIWfW8JnU397ACG9jPzZuTsWYsjK/BQsYqXZ2kACV
6/ZLNlp3yjjUbW66aRcVqiqwZYycNRNZmm6TS+/uSoQC0CFfy5bIVmjfAp1WxSQhXx/yEy/d7Noh
pF/o2E54tXgTdoFMBqda4PeotJfYSZSwiD/Mk7tc6MG1uUFHAW31bxV2tIgkAIMnQiFlV0v46onf
IEG2sJzwaTWrj8QvlIjkufrqv65jiq8Kk655xYPQ6RhkW1qPL0lrRYaHW5WSUeF5ZDp5/dumJYQr
JJEn1NIft7uOZ2ZamJli3Zd8c58mLOV1k03z3K0AFqdE5OPXIH2V3EI3FGrWCpr4/jKNAXSBma+W
F8yvK7rbaY6zDRt4kGmQsLjeVqedjbaANntJQH2iV2bDRlnq8/G5rucwqBydFdt+cHqC36W///cR
0G0To3a27xp74EkBxOYwCPcNjPneaS4cwwJGXbHgQEHHYyqem84mRnq2xJSUGpprpIinVV0CPO30
/33B669FJ96vDdtkoV6NzmdzAW8U7qMEkpHMW8Ot0Tt1PGUfTTvWyRVYFOUbEkPYU51ue/PHwkkx
DXop7YJgQqpdPjvVqkuhHyF0GpOzDOgyijRR/qzdXEDx5cO0RZA3h3NZeuVRsZaVFDCEmNTYcVAf
qDPusHhpir323ieuYlr3WMZq/YMSm81FW93z5SZ5xzgj75FDFfL8fQvK6zqb3Lna9mnrbey3LYDt
yVt9K5rlBrEtpZt/kmRmo9kpHXd3fH0rKQqgbdSYRM4kVKBwapptLCuQoou1/sGsAlGlXwlWgt+u
6nBYn1NIsJ9M2ZiPL/qqYXnssI9XI2DF8QBx4mP8PwEIWgWXZDTRXqnbDdgCH7/F3nUH1xGHNdBL
uCJfMI7UFbDC57NoB9zwLVVc2V2/cC8KaS5cUSDuubHQs+bnt78zpv2iJdLhyuewOSxx0fcvXLtZ
rjwU9rKGHso548EL+G57fW9512IYeEp293hbz5B602FnXbTjCbpcBJdlNAHRCJ2gdAHebGXAfQ0f
3TCXf38JjCFpV++1ZGBGUETwBZFl49hiExXutOQm+aKmqO/dtEvSmU9lCSYCxGgMEEeCWEe9FYlR
CkNft7pBlgaNdINw+VkMBHR4GNXgIckVD16D9WB1lSrLBvynpoichAtu5jbHwOe4/W37hmYsmejT
vZ4e/mdHUqYEzGxJtDJ3L+CngzT3GGVHr2TyI2vJaGC/hTVUP1oD95tsWKcTozRiuz9UBFkwaIN1
xk+LnsQ/MYNiQSvyF9mdz6g8trxx4lZJBJoS5JuBGsK28VyqPRJCaHghoY9VnFzWFFrn8DmkNNpR
D43GjVLc/H5xQjigQYrbU6S2tDurADJIOPch2k1qaOsiyvZmOn68ASWUrRH6XmNbSztLZw4TDFkJ
qGsmAfRBzC5bqvPCwG4GIGXf3MtfdHK2IPmgw0R+FXpmpPjHt6Snjn8ZiETrEGUrOm7sdshAumd0
V7xTv3e7MGepFC8k/u+toDGQS6aB2gJvvLEjOUXyPaLDIQhtCRNLnf0qIn22YS3zz08pGjETbu2V
bbtVHvU6AMFD10Xnoc1pmu1j/t3ZWbn+5v8kssatFkyQlGZ40PFmmWfsQu/vJaffTZNS7WYRnhd1
DRLvWUEvPsNcChHGLxoEpvMupoDx7l6cx3RLs6UK6bJvF6W/s1iodFaYaLtG4A083nLACGCEX7Rs
T0bWOoQ0im3XlEEcvmDQKsOGNOMZm7/UV+SJW9kqEodetEs2A2UtNnVzgWy8yHLauYlWSim+Gg9o
VItBZLAdmCXGQYjlWs9R+lTvHQpuqytriKEHl8XsLNyvfhT+ZePNSX0Z0ivKwdaF7HJqQ/kxF3MR
2uuAODpw4PosuLi0Fq9lmHzdVzwd1L5Xqd41NY2HqMhpWXLyYgGcE16dDTREFc8QoUS8M5v0XLIi
N015PaJkE6aYnKruFOS0BwUvYyzOXG1gF8DKn0HVqJDRPw28Kqen4zLa9NPdepl8IMJseI8TJC0R
42/qCPkBF1N4yF5W/iIdMGFoG2ItEX5AJzwc/LTNLGP4qS5I1D0Zy0FyQZupWUpS3mGcV/MDpACQ
s41bQiVljT+yZq8pjCVmi9OkdJia3IVFhnk9gHSlamdSj71iTQt8YVN69cYW8DOccD4MshDb7LpO
+Q0btx0dKX20A1NnnW594X5/g7fuIBY/yi9ClmFaPd5dwHDNcjJJEsWNIkcdSCYGSn6bhfsiqvq4
9WbNHwlq7wnsRHFOz145Tx+LHyZW0cSwYo3SZOKsFvNp0HTV+rk2LCeisQbR+PPQivngHjyshugY
7e1S8j2yAzfXfm+1Rs721UfxiybkE4zH5/lIxz9ScgnzJ2Rwt0P9B8Q0ltidHlavpNdvERpALaCA
MnSMqwRue5xGs/eQEiW/0vOhRkFSyz/iT59EDCCzjDQE+/QA5eIwCONuCc5tLsSuvfiIe7m4S7OV
iKCcZSBEHRLw7zbDbKCpildocBSYyTpdznw5YU0H465VZbo1X0PDQTwAPFG8pxi40LksyWFwHMnJ
JNPUzcZJyZxZVxGQqTM88Rd50X8+4u7smN2QEoitgrjhuiZnLncd9kcVdcD0rdSDKs96q1RAoc16
ZhUtJG2FOFbKaZLZmatt0SGRE/vrLyzquqwWLmjDqzuOjb1gBrOTu3tQ6ezdsBd3trej09/IwXbY
03iHLUKrA91Z5teZO/dsOyZLMOX0vFgQhQKTwMEtz6hj2t5EVZoVI6H2zFpxLxjtGsE4Eg7uGPYP
tgbIuUJj7HBvo0ZUCWcIuD+w0p4D3N5f7Q+fI8Zuy5h8X71f/pem8IWdUWcuRa9PPzC3dmwxXVPd
/g2sFOfPDMJlWv57LwMQ+aO3WlRTJgRbboZiqVvmNeYj+yo8tVSHipUVCadtwuWOpnjUgvJ3lTv2
quMfsyotX3+jIkTSmN9sJ2l/QwoJbA263gWQF6cxqYYI7Emrm/S94VnmBKKyLGyXy4UYqckZNVb3
JwFpkFZ0wiajcqWrkpniwWN+rE9bcSYDcBi+AQ0DdpnT5Vsaf1Ykv1MbzxsKcO9vFq2Tu5Cxn+Nj
V4dvLA+QvgnEGSRUD5gh0bH+6h93nVZauaKyl985grIVsNwflEDT/OA743WAZiN7umzvlCkbf9HT
VLiOO65VzdDjQpCtHiDEpz9yFvMAXtlRmPMWnrKFxZSHXbUBfSyHSUSqa8xd5asmPVj+fIYXa8Xp
4sEAf14qY7WBZKyqKEBw1WAV+Fvb/v7Yy/ZCVB6XuqCCBRyGSxyKD18uw7Yau13uhi+qao8p4ttF
+JLMXsdibu/uW642T5hTqu7eJPSIOp442c/lwlhYECHxtVfXGfeS2Iv78KF1ATi3Qh0QVg9uwXju
wskJNOn92qha5bGu+sx5JUk1AYW5gjz2jLciFnp0k1tWK1Fi/CjOEPEz/Y9MN4j5rotupk69xBI6
zbLhxcL8ktBOfwsv6Zq+xrZwlNZxIk2PY0fpVVunJh279iEbYOAgn0J+HONjz2aIss54mHAcoYBZ
qSV0W8y4+tQSZIhIOMF8T8+wEmWRuWEwz1EHARloJOMvqCiG1WJMi0LbByyulgf2iqipvOsKAohv
nKB6S6Hop/GUvj/NY42geGh+chUXyZ0eIeXbGCBmRWtwvikBM/xnH/aL95V5Z96lNW3fFXAC+BBI
iOYO6xnPCp1lCDCSdnctXAFYoZpwimuLo6db5oyHBVtDNP8nCP3JjSovL5cUdc8NhK5q3Lg5B+pq
IOJCYKSyCkh8VbBEPpcuPIal0t4OV5tWu0iVqMS2lA+M899ZipZF3YQ7PEBoVAorPLMqakWFu1q1
FD1LadEC11HLtW7zX9idBu3YJkKFJbD7k0tHMXV/iSXho+MXVFDQ9Jl70XjcqY0hrYUV4R5xz1i6
Vivbmdft2UW5OeQn02QgcXED7TB/6RM2BrHJmtWtSMqCxiBMsFn2zDGAs6C0bzG8HP2I2pMb+z8X
Gx+isz1NH8fgf4hTmojeYHQOK1wPnUigCCp2i5PVVLlvTZpYZuo50kpkFS2ipimLftWaGlJ+0Db5
nV34FcPB4ASVm7PgqUoxcM9BSJav3x7DYZKEtZ++WGmnRJwBKWPHcVTmJS/KChXQzJFaOzBOWDnK
XZnO3J1RIGkkadVOWeRUq+7qHA78RA5yl7hsbzZODgiyNQAP17YJnu1DJYWO4TTJ0Ulze35Ju9Mh
EC0uGnFnz8mzW3ff6MCP+C9Q821mhpRO7PPXEqNDYo1hW94APjpjzOFhumvhIR3/l8rcHvmPGPsR
Yd/hgOoaiYhLaiKToh8ZBScyjfbsksVlghDjPv8ugFJaritTZ7TD05YuTOopSDamyJefB0kGmG8e
6xk8YH977wFWRN7OiDADztTykyVg8jfHcw7LMgiZtgKrHmxcf94QNp4+lXHIuCa5UThnE+GYzjHE
Zt8nsvwZwUoi78v3UjHkwqyuBPwhmYdL1EizY55uFiP8EJUba5TBIFejQqDaIWgTW0fVUcKg2Mnl
ufNwmha1vIWrqMBDWdqw+wa8EThB4vJlLf+kvD+ptTYaYXGILAdEcY0WzJ6Lj++AGdMpLcMLxMU5
mQZWM95ogL1ujaOqAV9Qaak2RGEFR8o2JdFr1NzX4LuMVyCK2+eQ+gONx/SKLPhzHbBtGeN5gQcX
LSKRugJSgxTAGfc75fEVTg0Cj2LkUffN8q0f4XbS2HulWgym6NOyuHccLTYrCLA9oz0a3CAzALEF
kcdxra0x14Uw4gu0HGZPX6fZ6BejkLAbvmmD4Fd9aQcmjg9DQVzwMuWNSsE5D+VGanvhtOJ8hBYM
CZ5QWUttrHhGlARnrL99mBjNM4I3vFlNbTPWro9lcdVbOns7iaHyMuX20xqfRsT1B6YXJLEXD3bM
ookCQfqSvzaU10wnZUpFOrNLIEThiZ2NZxqrtaagSqxmgDOW9kP9Ky7kXahbqmO/WMGmXPIKXuIt
sdXiAERFBH+yH1K6LRjR44ToGddqCWmQRMhMUnzy2EWzPnUcGVhPcJIGncgclPmQtoxHMTMS1j62
KrHQD35OUoiwVdEhhsQf3hoiMG8mNxzodz+WF5703EecAilhDl/jD0A5x9V6ZpJhKeqBddZzlZHU
+KjRLkXLO0cTQJy1Ih1Pz7QAvFK/fsgKDZb7qAdQLNzhnHP89mh/xDYNoySZ06Xf7aryTkJIdOdT
OnGXBL1crslgvbw+yqtSyrJUS3S69tUtRwyVDO2CZIfQ6vb1NMOmsxYTsjvygytUTAVigY+RT4Iw
m1Br6TbRrLoTI7n58dKpe368quRx1bqh7rno55mfqDCYUBrhsOxJMjJjDpGyZG0VCrTYvVOa6na5
gf3SZtEOrqFWifloGDm0XO6D57i1xmCjusWm/ohEdZNrOimtq7e75gwY4nHkxy7pys5iod8CpXS/
lXth5M49W3UPMACf8cbX3Ydpk6F/C9DVQI9GpCpviwPPovV2VquLyLmbLy2J/LoMljx3ORW3yciQ
a693LXixDArWUSDfhxLXWI2A72odHqSPX6b5WnOZDUeqmJO3jNsNMLkId5s6uMeC783742tfdhzL
9CUVAa72I607goB3MWPkj6SzplMwYxlptwcT268dtzBySCUWlawZgP2V6miCWqt2GYU57Mos6Oj0
LXTxb8O5vGTXKIFH/aAYmq772CdxlBsApx7ddboVHekab8CXocs7b8RDjqjMO3iSnUZGwladXbmG
EL4EIZG0un+zA3BXKzR+pjjpLDv2nePbyBAqOxbMSzdkeE1M+F+6pMIseSChoDsrSVrb67u9FcMw
gxYzK4dLFlolXGWTfspFTjAYJQAluK4owE74Jl308zcYWIsZIE7R6gaJUuSQBkWTIs88t3sRUrBe
yiqWqHy4TP3HX6Dkr5NBSRlRwzwLQMOY3V0IT/cIsKou5VGiTEmMQt3E6mc15vpk3fgWGqoeWH4H
Oucm0kSb9sCQ5cBkmefngzMffWGZ5XwuPjh3cZ0lsecQqXXeh9HR+RMtaMA5fmauNwz8CgWbKaNH
TiDSC89hsjuxjXUgVvxZ/o4qTR2X7a3q6hyy8XwVfpsq7pzOfaDqmxL4H5Zfn1P8DcrSFAnbZyZt
vV4ri5O+qPScLqTuo+lsYQ0oHewjnJXXBcREcFYrBPAlKDx29bTf/BXW7tqmzfFkQ5rFmsnSVXZs
PKYrrvwxalrKeg+drsvXJ9y+yTWzxjobomaAWWE+9V1umO9Ngw2MvEB4Wo0oSShG+nroxmz1t2A8
HuDLpoDYK/tg+coZHSOiC25EbN8dzF/T2lvgbnpOs4UyWtbUbOX8Ev1sntesMZy+1Eh18hvumK6D
wk/iJup0Kz7usqDLq9EH/+bnvC9hkSLt6vkETmw5FT1WZFa9X1cw2ZRyw8gt9JlZVH1rhoWOV1B/
5hzuaIrsLdQr8njCEaBC5aUPXhC+ztFyV8CUf62BioZNHHCpmhovrrVgphTsF4xkwRQsPH9ifb0Q
yONFiWi2jYN8+etiPTBQD/ULecmuSo6z1KW2cTbc7/8XiO7xDa4k7UbZVXYXpRL+Qb5R8lHXGSF7
ZmlZ5a0pjP0inGZ8zSkg8yXptoxKHoOD9UsPTDWAB9K0NtPJP7UBjlrUEfY0BZqMu0Jyu29SpO9a
kX9LL8yefc9s5Upb4q3BIUGWyT4AXjCKdJKGjMqtrLtfzuDrh2d1cdUSdDsgloXQTz5JPX8cDLrv
io+SCE0olbBs2BcliVLrPZo6s/TZb/+E/dkpB2bggu4P8jwm4aMCa2obxYk9KvbAdV/Dr/I07fVh
RH4bOwFAw8icCD9zFtuzWZTefw98SWGUeE2mWoLopFmmpE0qb0dxD/yCsUrQ3HLpZUQATrqrL/h9
l1Z3G4bjiiVjwaTuAySL2UQ92UszR5doyeBPMfxZWjMu8wNCqK/ae1c+p6wixh0/9XKLrpUXJv+j
Lzb+5cbf1DwB5lx+S3AzZZyp2ISQUQS3xqMZp+VZtdWvGWpY9nMqDBJKm0I5QFdzMQM+ZgytNNbm
Nu1jVnuF1epcOpdatqfCPgVTivUM0q2GtVGZscNA6bRCQQaG6unbtZbKP5GLkI31WGlcfA1wvP6k
ps0IQMDV1x5xeqgU0zZ47Q5lRs2zS0e210skdRWnAABOO1S+w7Il/YIe6lLTfZUG0aaCNxQ8hT1u
7eQl8xqC9VGT9nosb2pdUzanAem/Osqb2OMTmiEUGrptvDdEhR3GotDgPmgdBkyu6s/1bC/vq0uG
4MY76CEvj1ifRE5NhIdtsGtO2RbuZ/WoYBPpXgEyssibU+WREyuBMgb2CYX1KBg2rRFJL9CFkdJD
msXbF9k3ssx3UG7W61hzPte3gszXIMj7ZUJ2VQATOEF6CH+6JMJVC0jsthTX21rSx6cKUi9QWubG
OTLgWWMMG5JPsPEXKERKpZAzZm9dPEj2YvGK2tq7OcSzpwbxyVWeDqcwwIl956CMZTzui77We6hy
9nN9Vy/mUTdX1eOeH9EHB0WtNbz+Z5hldqw3Y4k2i1K7CWFdeS45qoaBkDwyj4VlKRnKP9HKz6JF
ELFWnn7mToTAJRgkRQJqpFxpfy62yjhMAUM5uhHBGfLxbvgqhoAwNi+A1KF2+7UZRtIUNX9nHKx3
HdntO7yRBCXNPmEbZ7K5ETtCeZQKlHLNosy+94tdeHRsgnkhzTFr7ti0SGguzEgCmSN2IcxdwX+b
lS6u/wIKGtBoEZqq6/MO86wPF3yI96zJW7pvOrw9QYJGLZ8BexrJm0orVPfFP2EFdNEQg8dr5Uqs
fAGLjYVDFsbNyLOEATs9TV92SBraqylNbnKpqQ5AwxfajyRTxb1dnMtRqX78Su72q2zV5/aVkFhK
L+gLargD65RhYi2n3WD1zCuAu55Gno6jzirXvXBt/Y5jCycD8AN6gA6wHeSXMnOiIy397SOWDOQR
QUQwn0q9xvcrVDe69mppj5rdY31ycJ6D3PAN8Yc9fzu5TVLTT3xvZ9YfDC9YYPRzRigvNvCda6Ti
J0jcsm7We0gp8Ic0l1Fgs+VAZo8U4A9556Fmo/GVlEXOhaDRYOdr3neLQGDS++aozXIb0tA0CiPh
HTzDBz+KnPQgeaX+gju2MduZvAHgYiU8kpPF45+l+6caddyMCoPdWn2KcoV04vKYOd/rpLo8Io3S
l8dPoCaSAPhcg6TIqbOJK6nseFJYGJSzTyhpjJggkBFtFo9piwe4ejnQPHXseLzr1t8mPYwZ0Jth
OqG4o+lBqVyy7byqxT+lS7ezQSG6Hv3vY8fu8WkOaaf9I6CrImGirvu6sWtVC2TdFF63HcNigvLd
K+08lNpLhlb9DTcRQp472NDTtNWT2adTHFvib0Ymr2dHchHcsf8jZ+Hki871SeXyqTjcwAzgxOuO
Ft3II9fkUnHGXll+K1GTJgi19CkJEGzrU7a0jd8+BJnlpK7NotoUz6AXeXBPLAz0LM8ZrCp6q/Vg
HzBGrQkaY7RoeKb2srZYnJZ4hXp5/qdDW6/s3yKzHtV9M0lq7xjVdbihWElasdFhm/qcOGpdCUQt
lrbqnhx4HqhYR/HL3iq4dh5fQe3Tas3ZhdgFjSaaK/08FeZjGzOXEXoY9rjxVL6PffPoZl9GPsLX
ScSOX2mBHSCnhSgKMYCK8Txjt86dSnN7KbAV+iAYwX/fuDCNHUdWs+Y3bNivO4PG9vtLNNW0bbIO
kLBUl85fbFHaS7AsobkSFN7h4lPn86fCWOx1UPr/emm9IgH1sVg5RVKvzLhgib9KXP1Q31i2vLpL
RbOoUPrLlpOajzCeTGJHhBkil6+32MXROb/MThjCKHwuGOk627XxnlV5A+3e0XyBKeCuM9DJJoWO
oJ1H4xQlZ1SuKJkAMMG+tN1g2sU6wbkFlaqdKMOWSO0uDo4111JgI9qNpTmoBTAhZIdb4vH2EofZ
hm4+8W6iF/UDGpqmHuBHCFhBmVMdeUljPetax6VmBvZbVOsskrDm0h0hiK7xy5vppYb6rXcpQzin
00oCUB6NBjBo6cqqMzpyfYymLSeDJsLgcE/EClX4Mh1x62OHwsv4W8jLDTDehdt2KCdss/QjsyOJ
pwfjuSZ0JWHnZDuTAzTZrpnIjUaKYJCmk3c2q6o6q7yyAhykvaheM7G4r9anWCzdnYr5SgkPtNKS
fMmllEkMUYQMq6TlPYLDgoTFJb1PsdZEjfz5lkPdvl5lwa+h4RgB8+EQPese7VUkO2Zn0VH1e+Nc
sZ1acsqMQ2V/l1TDK7uPjtuNg+EUj5AgplDjE/qzFZZ8jdOCxM+k0yWmsql9tKivtgD7Z9iwoP2S
aEKeRIkxsr1Xluas3AsBe5QwzDRkLHYpjnXSw91mctTnRR2V7Ox5annyd2I5FGqNaknsSA3h+0uV
Pal4xwPLVOVHPjy3MXshVR0M8IH8R3dITEHAP1WJ8N4g9uTjGSJf+MCNbfRUlQPb0MizyiZsoJa1
K+RigwOjJnbv2Nxs0wmzcWGJapAUdEHtPDVB73MJnN9aZe955WVBNu0UYy3qxA/spbFngli68qSo
1VY3pHAFZ1o8n6ZlQ+Kn5QRODL2r0tLPwOHBc/K6TI0TtDf51u15Ncj9Njy/bjEJu6Ip0dMsyS5B
aECMO2BUzJoW5iuL1UJ3riDwSqHJ3QdEDgafvBAH0V2shfRRWWjlcIYsT06vbbXdYhvw1MbobOfZ
JQoCsz0VO/ssLS3Y28TZwq8duA1xNMbE49KPZnLNefkLP+/nysgphc9v2cQJ9JpcGp+jUdmHh1gr
VCzONsqU8n0cnSjpsWNEQRamTfBcuHkH0JG1J3zyBtU79MhvdVumonCDdNrftj1XiVOySYjiaFKX
XYSMVVUn4u9t6iSXmXwnRdVOaUdmLyVs0EwTsQrmHUtXnlyDa3THNeKWd+zql9TeyzTw6kp02nfq
YQgP+8X2BIECUsRLc5PQmtgbfbvaIiZBL1SrZGYPiDAW8oozKWUPK3m/L0OdZ/hjIdFdX9IlN4Ck
QDu8Q9tC/y64qQAeOCXrxeOq7Xo5JbY5mTPmlHyiQFhhPJbgnipZ0nwWJss6HDts7zjzhnTl3ueu
UGz9pz6Q8hthPT2oR5GQkdA7WyQC4TYm8b54nNxZlgltOsSG8l6O0J2We5Dd27Hw0EN5+K1ZxcrQ
0bJs3wuIK5c7pOpGifDMW1tObeD8/PsjqSvs9915FiyiFBEgFrsU75y8KOXGe3l7Hl0lx8GNWjPw
y5BYdH6AHuB/nOkjyAi0Yrs+rFJJqBYpV/Pd93IJoLWxf9021N442z12+/w92m010UoxWsGD8GTW
rbR6jqz4YjSH0KTe24FZvNyuZRqlYVDM1VevzfAmCa8p4A3ZhQDRtmK/YgQFMyccN4ETrSzVu2mo
Y8EvUxKHxZZvL6ABQjZc3eongIjHTCCH9HbqUkDtOqwaD3HOtSNrmLqb4BLlLpN5wskWV3hwvGGS
pxslKEgiPLkdg2spIqgKxaUQ3cKKHwXewLOJQ/LoABDlY/eF0tMHhurSkZ7vNn1Y2gg1zJp6E6rT
lhuO5pTBN2oSauHwcAns1fk5hGVoEL/+xi0nt+IuyxMaGmPcN3EpBsecESC5HcTwlODn8z8sZ2LM
DOBhH8dZBQG8tjvvPbkbE7jP64g5OfZqJyFG6eyVlE/oHur+yEOOvY64WbNUJE27IWqy/aK5CpQW
LrVOhiizPwno2/KSBpwmCFlOnSfXWyyB/j5hzJE3UqkRUWsiSd+wncJiyS0KIHPrg1aNGZJ+eGji
1Rp9uRKxkOJQ/NQROfvcazWxc9hgxq3vUedBakoJQxkSolJkPfgbxtGZUMuGKSYnNdfqgfF6Xez5
+SjNXIi/M07lqvbqM0nUyAokMvR2ry0nK2DZUvv729CnrORr28CIVoMtWfQlH4IpLFkPCdS0/7fM
ztPxOyKijyV4vmPizzIOSI93loRDlQG1q0Mq+4nOQwiDfPe4py+2Uagxqcy7ptDmoSR3kdCDuNKL
x9Ou9NLXs6XCi3cstsCYxUKdbaa5eKHdP/tJcWDS1zNRNkMEWBTnx/5SP9OBr5ZQgNwHtW6ZHNxh
GnZfjqasn2eB1GYSrP1I3ownHVMZJS9m5C+LksAsS1IBKqE/AJTYWADmKQeeQXKIKZ8nbBTUwgnL
yOY8QAhhMOj6aI2mXNBcg5/ZsZxwjKASg6SBhISEBQIMLyVIqpIFM0IfXodqzyRm0wtEAEPmK1J8
kmy3etXyngDOFXWYRHNlHrqr8wR+/yp6f4F92NKkRqNGAlbvZzBpfSwiq9dIXNfsnFzk2gwMdTdQ
3Ono4gbDfRk5tRzCID+FOome5aZ3FWFLtIAeH21bTdWjIWwNRCBPzPzUTBoNpyejNe0ieRsJLLOr
lKSvpyKAMxejV46E+5AX/Lc1os9Ou1LzE+/ucsjkq06BC0AQWX5H6IDCaaOfPGZaGuprtjHfgkgW
QYmzvokjnCX8c7Milzf7L4gIuDmyNa+M5wNtH5+defzlcE+vb5iah9X79lLXdcLT3nXLkOHjKGrT
yod+4ydze7JWU5mnOLaySRXzTyd7NTLQsIMj4GRO2zefDzB8ETN/iNxFlRD2pArD2ZonPHDJ0ZIy
VXjEXdJSU8FeYFudHjX1nE/l6umMMoQ/X126wAqMfuXM9/B3+s3b7NRvvNgscUr2hTW933QKL/S9
3q4yzvsVHnG3cz6A1izif6BHCa6iW6ENn/M6RsN3vQzxYCfEamrmornBmMCqHMGWud9tBf9NjpzQ
YxgLgR/ZP971Vo3epVLmF1hfH/jFeL5GdyAdo4mivexcR+t9SWxosOTWk30p6ZxjbOyF6NlPUkJj
wZl9uTVErH4CJEnF8DAsUv+ovJluWm7/aBWVwxXWnJpDm7677ogvFIP/gMnh0pDfxv38BKhu3Xr8
6nQJ3w2n8tr9XL5dqiLu4fR4uRvy7gVHo0FwKPzr3wo8CVmPHr+I8ALxTsTmnL58gNNGsrmXMH3e
YUnxi/HbKC2moyVG61hH2c01yAMfHbGI1FKBolXTDblAnEQzR8wZ8LyZPTCZah5DtfaRsW0Cca+L
+Dzm+GSvg0a6o86+xXDJqju63/0O6FgmqdhIaEQILWLRXmqHQVf1HoZYOEIA/9zfT5lXYsuTNtX5
0vOqEOx+M4tsmvfG4tcUO2S6RNO7tME9RK/p86s3fWUQSCPZX3hCT+6cqEwO4muu1hrC9wLmA7Hu
Z0AdvCPHiDElzOpt5olwagm6+5fDOutx6vKVS8/gX8fwmcnYS/EVUpZrR+lggayiUH6cMCFG9ViA
vNtJ8rd70lrKOMWQJ9GbdHe5/dqz2UE/T6BfVsydiEM5ztsP6FmOe7O/1MDH3/Sh0BBJ7vX5/Zr5
5Vh8aOgcjdg/Cgn0ycvUgHtPaJLAMHVgN3fYAB78zNfJNG6Hjgj3eCpVGG1VypdqRuqZTpA8Yqce
MnwI91BWmqHtaVT/WKKh0Ebg+Hz40EL6smtBhax+cv6JTGR/sTy5U/ryvYGtm678dEvkzeU3GRH1
qx6+WdxWoCnOJ2Kc1G/C7QhX6jFaYqhs+GFtl4exXZbYoYQjCVlfHGJLR3OAs07nFyYhRyNTFoCp
jncQE4rfK5bBInCBIjlN7vfuSxM9gHa57vhusudQtmkdco1HpNjOII2VyNBQR4e5ZjCkPQoAfxl7
xmNy18pVrVoF3aSUh8YLI/qfHf4AEaZWZGW/JP+0CoXbpBgL2Y+QCR8s3PdsbokF9YN806y4G4wH
ArHGcBlgy+pn5xsW5eTUJ7pquEyeX1u740+KFgEAAYIKCOQNx70cmA9l4fyPF2v3b2VXoTK2PWJ/
EQBJnLn7DnAlHoS31e8gqPRxItPejph1UJkQFILfOlAz1rkdRC0lbLXz1olRzdVGWNsilSilym57
2nkZMJ9dVu67tpFEDCbW9ULqABY9YICOTxTjqA4UwlUHlnQ4jTOIiPOUVbUZOT6Q2C1jTg+rjW5g
LW8m10qaDKUpup1GKCcMvzezArVhx/fjmKNzT2SrDypODT6RVsOCek8fS/1QQQ2ZGguPjAEfGgVI
yQ7/TZqnvJIAZt6uOZnoKZAmTPrx+0yvt1yEnAwNU2BqxtkcIHGQFIOjqNM0POchilsxFWftYTue
WwhV7lcrE7MSUBcAcO67h6YKpEY0pfttH2xgEE2gIWa3M1cBEDy/FZ/znrvvzahn5SdEGc8Spv7l
sTqgAUU8hI1PfCerWgofR8m++e6TXNAgU7Gwr4LGa4z36bKaeX2TG4nxJn8kIELiZPfa1lRt8zex
5lX9K5kjBCPj2QQCmeCRfvPnNG/plfXL1goaH582trZXixG3ZkOUux7elSjdn7u8QsFDkE0FDLwM
ujRHxnVqwQ5yi7hPD6BfdLzHPLV4Mp1wtdzuGd29eg38So5jrJoZhe3n/Fi1YLBEwT8+agETlMO/
xltBGm+AynHczjuhVx7iQA5Zt9efCT2oi39suhPAJRsOw6GF9J1prxiML34bPMdCBl/mBP9igAAw
rRUDka5emkM8eSnNyFqLBYRN32ZNkeZK/3QJpgUTkuWe1pKKtOpHlnbMm83dhfP2HtnRjrYoRbo+
LU9Ca0jp4oFoNpKO6BNxXmzge4c0UYHy5iAPszgX3aljTwH/sbTyB3mSFfCmdJzK8gl18znR5a8u
VZBkC2Rzm4UII2MSlZTiDr3juYOF2fMlQhtH3ofuwT+2F/W6GDMHarLGnSVjT8Nn237kdvuhx7hI
5gxB0WM+EKYAdCvx54/bPxxXkS7S0OvKCa8LiPvZ6kMnHmh2ZyRNz46ARWcHWkH3mUOQxGwXZzna
XGh6i14xW1TPwPnexyR8OpSjj2QMmtXR7I7JZMWDoXt/BiVUlUM4n/RZyCGkFxj6kuorx/d8UwnI
A1RZ+QlAOutHXWvczDHX1c/e1Mhyjkt5Rb+0NqdEEWyv0ZN36t03UR81zya/uBz5QpURxXW+9+Lk
gm00zxosFQj8ToWtqbtdE4wjat0Xf7h9aY3vkpYHCYC5UCaVUiV32vV1rONAchE7mHUkx7xEWrmY
GvH3RAwdrzVbtp9dFJ4+Mf7ZfExN4tKawJtPrVFTGZKe3yEveH6yW190+GvIENAIgTl0sNOzAj7N
pRgEMfNKAjzhUcmjVdjuihpIfNcaRZOB2qhxv+3QbmFigk89fWY+C4SaY+NlcOQvs6o4eGK5RZse
ThPEHPvR/5dBT9mQ6lDlOMmdrqsXF5pi5LXdkokrMJnuIyeJPnQy+jHEuA2KC+a62PqD2ohunMLy
EGFIj9wbxLRjMK+dYZflbpYJdBiIsthxjM3SJMk1rNurS/+Ufs0I4MMwagNVcdEA4ODMoX6y0m8D
qqJ/wXSRyOU0/8hIJb3ON/4w8HyjZYgUgLDXuuWeqTCgc7R/CO84lyA9xPTSNJURsDb+wkgoR7fC
r3JkHrpRxyGxPyXSa8XL8Nk6DvVMbU5nTRx7CE8KcogcilMGJwi5Dx4TIYBH9422Nlq2uVd8t6jo
15TPVb4bu6nkZZFVWkJWf2BvZYdHzCFuYeXgFJOuUy+iVZO8gVK+XYI46YlTYeG3IzOn6HLtMz/h
LYciA2PotZyoSWXoefY01cyFE/ifQNquWds/b1HGpXYFrQiCj2dblpHXeitQQGl1XCvNj/Ns8qg4
qacjZ/5MQQ3r0zpmftEjQtXf89jLfI/U/Vk+W1qBPrHcZYPedicyHqxJ8PkCFhtIU8LUZwMvlrKF
jOb0KgKVCmwvBKKpS6h62xxJPc37Yp8iHqiOCtZOUyNb+9iiO4XgLS9WZrA/6qo2DpBwqLZ3JiTj
9wMEWrmaZk94q1tSOLcJeF4/2f+V4txXT8Terl8cZeZCxbqhreqvbu63RkS9PPS4uEfgOHKiEC81
SKxozSoug2Cwj6K5AxHr8qhvIuQFT0462SAlgojJE4zZ/XVH4hAY0rQaN02pDrHXusPe/iediHYD
9qfxsNDZp182IbcVQBBaP5XEXk6H6VuqJhUMs4K5jMYCWTev7c4fj9a5q/D7r1iB6ocJ+0yBml6M
prf5FMu57C/s+pDeby47dWXH22+J9t1h+eFnOrU8T99F30xFECH68/2TMQdePB12ARK2zyYEZeun
s4g16CN4RccaNA1D6cy5odcqjk+lYmJu2jYNFB+rxCjBRmIs43j6fhZfTJOUlZGv2H7Fyamy/izL
Sk0N2JkF20UPYX0vguaVOA9g/l4YSsVwzsSPnv9tAqi3FqMneB/Nqxu8CqSFUMwAfMnK6lXrgeZ3
M0rg3ld7tbJVdLab0CV62FBI8RczNMR/XqkzJbiMq7rCRUuZpmyK/2gUlX7dFphYK3ZlMcFlZ6Tg
NJeFTefgi4MJmueDVaBrK7D7Aatmbg0j71XobmrTtBzH8zbp7C8Lk7aTkCio+u8p+tIg/3j4CDji
UMgGicsCNHutG1h/m6NVEsKSOCZH85s/8d4uoIymhqRXFh6l2xF2u1Zp5pPlLz8HvsMFEm1/6/It
VybhBPtSii+ejb9M9fugkA+BG3FHCalEjApyiJ6gW5AqZ2PpYl6i2RjbQfOv3lhNfp4f9cv0pBJp
7wQSa6N6cft4kV/NA94kQLK3iPTOBIiGwyu+3pqOXYYRlw1JlrlUavMVnLenAgJ1WmTn9e+NF9jZ
xKFVHx5/cAYArVSb8F/2LeOnYwBb1CCToNP5EouK5T6/0xFoigO+AUpIKory+oIT+T4TtIuA8I2G
moe4vJIRSo07ao1KqjrxAeNK5YkFw9akZNlnInSNNHH9m30ezr1r77OIq0EvZcjG1dx59T03b3xN
cRONRV1nUzWy1su9yxosMQq3Irzzdv7eNUqIIehOlZSsFM5sIt9MBFR9ngkMXBD6yoGN+8f20/rn
HKwsrIERbCBxsJAUU2mKNZHXm/pzfCyDrRVIoFcS/Gffc1t0mJ3mQKmUBAENjMrFOQUIV+CXcCCM
t0aDr1WyFWkUXNax3kWqhKQZHV+rIYzUCrZzoyd5sEwe8w7m9O3gJBWk2L0sa6nR8GygONPCJ+hU
VzPNcxiYSeBVH26LwRlgB1+XwqZzHTKBnO0qT8oDFZwWyu4vVYXHKY/YepWwelw9DXR+B4GLeHv+
+Y3jcxldvt3zNUKzWSVw6koWht0wuTVvvm6M+qYGFQ/kmpOAA1sJMvXdWsqX9xUIzHrAos6GKUNN
58YTSlPM5TftZKclJ2ASPrhCOA2zzVGuI87reyyoKYma9EO1sLOXEmfNFJxUiYVRmcr+czmuo1G0
7Qom+F0JC0rt6iMqLVBIuk4TMafRcP4yW0npqBhPeXjIx3YAvMM9g4D04B5QI/hA4FepmpHo7eMf
+NYY3rxf3XDQwGD6NhEQlCBKj7EtTTpkoJwQeVt2Om5dqtIGlIwhJyvVXOJj/wyLgXdp4GYwqyUW
x56IOwac8bEResc0Vw+IvApMzX53oZLig79+NZx25AnzEhzD1I+iNbcEfOLs1xe7f3S9AeMYHi6q
fGoJGtkJGWf5LVgs3Xc5bpHSnUssvIHZoX3TbnoogKCBXF4CHYkTzliC/Ax5GjZFyt3z7wPTwXZn
B11/YTlLVO5X9OOLxdbqEVnQuowT+jFrKELFFwOIGoYVNMF915oBF2X8WaGmBrvawWC1zr0L9SDj
qfd0O2QGEJN2XK0jjgQUnnQu71xGQrr3Aml5yADl4Wg6kJmZD+NH3tTzAt945LL/DyM2wDU6YP55
i5jdjuZyomhFufiWuWfhwu+mFnTp70UofU/mfvm+HQCfHwo3e1w4sEH8k03uOyDKKmYcwZ5nLjy6
0r3C+Fivybv0LFM53Yrn6JxiQoQaiGGtSAh20ABdIQ2BrXaxm/qQTLJT1+18dFfOoUTIdeCJLUjT
h0nKuV+Y9r5ifOqkKpqglQJuvGOLxjsOiJF/mP+7TgrwYMK/fbFqJSRh6BK0I/1+5glfdp+TqV79
eLzyPmToLMUEjlD46dAF60J5CP7xJNGJ41j1ZvWxzcWZ3u2/FLjsLS9G0qlP98CGkac5gLt9Kp79
HSYxPOd00hm+LhjE+lvkKrYId/0vIgyWkBLbprCzDPhRNRBoDneaHXT347EJJAz5AzHVkqtiTuYr
AP9Bu+/EwyE1z79DqsZVaDgL3A/zp0gI55yvobOZ7sqAIa4yTyTk+zEde7kinC5TEq1DbBgXupP8
Toa38tRfNuSuUiH7Yjmx0iJG+ne6d+zl+F7HnWDCOEuefzfdrQenKYqVvWfelDrYA4hXwXLdHUdf
lyzI5ExyfYEzlsSX7rkg9vNaXqagbe0v3GV+RLP9ROkb/paBSrB8zBWa2xYivUWGnCzd3uwPzk7o
SdwtSulZn7asgTXMg7+A2QYAlMSasK6pHyuFsLtyQZcNcS1a+Dl7VLdUxzayYAr7VBbrKQIcbO0g
koYc/4syOk6ToJok4YjVIqWY8Vg71HfeBVmSlG8uS+MPLle6rrf2QhX7VjnVxGx7DZcxklK4Kg6V
ZpKe5DG8ms/174WdYRJpkLLCLUYSMsLHl3iSNOTN7RH/gg70d1u/YqpoJi7TLo8PtQkW3vDi0kY8
S4CP+RrJhx3bmeq2aoDhzz3HKF7U5I/OfiFFFLx6oRdZV2/wB0Eu5sX/a1AhsU+urLJ3W00Zha4O
W3mT0jvl2LBoQvoVrwsaZcZGacbEwM1aaosmF/vSwlaGdHVcvwXhNX9dfg1sXxdwAiG68HaAoKTa
P0F6T++ZYO0SdeHs6gz3F90Cc5MO+302S+OXorcNNY4y8fMcOH8YoKJi3y4gtp1gJatlUbxX336x
l9S+HOWTc3+LCxDmdBUoH0cLQ8kP5TjiKHBuyEekgRoFSPpGDDIJt0iH/kMea/7KclugSdyBUp0a
A4bBs3Fnb+T/XOS2rXqYd64uv3Ylgg72Vgox6oNXGshixew28wsmyiUWTZqPf6R2VB+jP2cVKH7i
Vh18a0SNmuC5JRPIsTqipd7KRnmfT4w/VgSX8cLI0760172vP1lFabuF553etdPoRdqfZfR+E+sa
SkcSAbGbSIRKsBJF6LlrOIeOo30Hv2WKsF2OF/5elKgk8g8gbckVotIyO9DfF5dwPoFB1LuzvU0v
ev7qVrVkTS4IteGHJzXkZv2Z8Eb5c8punQ5gNgLNFSmkh+kneWiNKMZ9c/oi3V88s4LT8Br0KLaL
bZvOT4OEtU63N17WFghougAcJPOJb9mh+LlzL1XK3DxaGAwiNeBXtasv9bcFJ9Lv0AF02RZ/ccRD
6fea6vBRGWlLvbLCvTWizNg7+JNbKTvzUzyT+O3THd3Ct4whoNsz0gEbvTsaUr04xCRKIXAY7HDM
v1VF28xEk4g70yuoMzsiTautDNtKbJAdURWkvjXSG7HzuQHUrrGCte608PC7lGBBBHgJQL9SpqAj
oNvqPGy9KR00tZ9PQSacL0ASND374WnJ4nuB9eGeufpzoWEX+XkHdycJU9VQO5bK+Hif80if6zGJ
Gh3LsYZy/k7MaKh0/QYIELKYjenLSng7QWWYJUKkYAWU44g+XSRDTmPzssRxHD/nDs17floEptKz
k9Id1I7tD6Cro9NdvZLXsijLOeCbOnnT/dYrMd3Zf2g3ufJSqEhVoN8kwsE+uQMGsBr/D7/YPQCB
DoOBVqNeWP+A5+W1sTLI40pes1mfKELOWhH8pfJGT+tHmo6Y5ik9d6syulLJoxfZ62AJqTi/BgKp
WgyLYpmyu8/l3ZleIXRRArpqkCrjv5lJuZCuZ7R4+hPWw4BBdVVlH6YMQ/Wnh/yjNduqDVl2ioRy
3gjY476gk5FDJErk4bBwz57ACx/Mi4WPGkezx9u8keKh+zRP+7mU76250pncvW/5kJ4Vw0NNYPI/
jJnl7JQaOo17v1faZoDfB/zG+BfL6qlmJzeejesheA1AP9BV+YReAbfJWsEi7CikfEP4V3rE1G6u
CFhnMpq/tls1r6pND8k0n+1iIaNTlng8Vr4ItvTI9ADmG2BC/vxKUcIUIKEPol3Et66FlVYd7aKy
WgP4mA2amw78FGFrUUlIxzgeFd24C4W9LUkKjJYnQ6pkr6l0ud2/xXUx6fCinGCJGCZIJYM8e6qy
zOfQw6Dqw8NJWrKwbltYkrkK3qEpM0q/X87VwoadiDcYYCLuFoFrD2Za6OklqRtziHM736DUiPji
s4FE9xOslOEqHRdK2Jme1vXTR3eh71o0tseKQJtCBH9mu6I6pA7OBGJhznh1mG+3VjH3haYmgml/
sKLJKLLdzwcVceUFj1GbdDGmt4GK/iN8Oq/FdCkQgvIzXLgUGoONNTygVaE3wLO1Q224GEBbghBa
/0hsYRJAUdFSKa7umKD3d5jYh5eh1HLMMQdvzsqnBfLmqTtXOw+ewwvu5E+IU3biIbJcsHbolUNv
uXnJG0LKN4yBV1Khua12fiGmEfkYDAvxhig9qw29ABBTbHZSwBC2IlJGDBPjj2xMvthoF9LYxyuM
KQvayv7UWT381p14Cn1GZVK+jVFCwzEUPfO2nKAbH02dvunYmVD8tWO6xcTsIwy6uHBzG3hu1Deb
xT26wPE7TM60yKsxLE6rIucxdp7tr+5B8fjYjagb2yAoGbPCF9zccJlqi3rEbPrStrUM8Z/jXO+w
SwQrSNbl/5OchH8P0LTpKz/WAOYx7Xvli3m6JNOZ8MSbXg2/662rdfy7kP1Jcbw7LzbRNsAOGsUn
tnTdqmmAxIXRp1DKM7ruYg+AX/u1afHAF8YujAlVwpJrNUWmUL2AdvmkEMTQd1WnpxUXVBvjTsHM
f9ITiBv3OPUODTKeBO4tjKdV7cXcvXnmnINbBHcPo8AEKrQ2eQWruv4kUZ7S9o9mBZ6mHlWOb3F8
NF6VwF0TQ+/lng9ges1XzHApfGWXke6IjpulQ0uN0JB8AkdCwSQoqPGs0qb1gm0oUjXwTr09l0hS
C/OjNhhUU0MX1Pnl6oEtuETNxgRtLOd2Fr3GgRerO+BsEDtF+L3Ai660QOOv8OrDqmSUbHxmwV7F
xBvKTD86lFTH4VzKUC/HogKA9OhoaE8B5biLA8EeDyqNi6QxVS+WiJ6Ertn0cET1DCiosQ7kyIBx
9sihxb53wyCXBQwQZusxiWel2j1/zyWYz6RFfN0r3oojE+X1kzD1mq7g3vJKnWq53Kq8bTdCSh4T
UoD6U10+1oEhrUGix9Bgs34a+AzdMhWUMkeLmFL5mdjE24sI6gsVC9l2/fOTSzebeWWRgJdVq1/A
jXjqBfHW/oJgaPj7JsukO7JqgiGWNIq6figd8FMPxOjKEIiOKZWV8S5CbLudcZTbNWh1pXaP6ZTP
oo7NJpIZtrDqfSNjk8DeUdwQVMZGWZzynBkatY0TVgf0w4PgECrMgCfY+1dsgiqYRlJWaxQgs0vD
0sPqgzSYP93eQ+Zds5kdItEjkz9MRAV8gyU+bQYbOWVRVV+HBuGyosMa9atF093z3KR0L4vNXNKa
FzfKk3eLFWiHvUaetJukUuYGxFEwQtub+OznslWyRYv6FC9mAt9nitRoibNf48LzUgBSlZfSalqB
x5NwjwHiuzSwBegyy/kjculpOsG9DBqX3Ws/w8pjCdXUmJw4IpKWEJN6NEF2S74txkT/2gt3Xk76
goZ7/ut9SOMDGXY98pOcHRkVPGAXYdEZyctoCu8jmdnZIJiAnVIrNqYkirFyuruOgmjH2OLepJUB
YN5ASWRZ5RnPJlknp/lSDBU9VJcqXOsnmNp8lSZFZo2QI2Xvka95L7pOOXYCFj9QTiDyY9FzcI0f
4z7l28cpLhOTQHqmugIY9/6mOyr7RprGi7kDpvcBc5YNbgNI/BTE7gst1X5nYNCC4NlZSLxXrqau
u09V+1iAzUZwcthAASjybEvNMOb5wyUodGYeVVw7JDHuuI+o1JAXOb2SC5rMe3CiAET3y+fBC4dO
59NaOlaGJYBjX+N/PHi+YYrsbuOChbDCzCNjaMeQkP9y4b261gGuCv8D8sbxVg8RgCAi5ZAVDEfC
wurN3Yc9ipq8yXDk/T7LhyJJhpKKHN7rHItg4OtIMSx0oqqckWwsSI1LWRfWTUo3LZ8LBqSn/yFt
80tWaKPDzsZBFBO5D98s5kJZelBbeP3KwojaG7LtRZJJ5mdNmrZZB7ipRfzfoNCNlwfYQXIxoufi
CwDIwM5JLcd98yrSXvh/phJTHD0r5qqT/dNV/4dr9/XqjhHJlomQoL9zF+Uv6lPeRAPjZ9WjVIx/
5doGTDGOnBeEi65aManess1gkeFm+bNz7xLsQ7h29JQ3dx4nJdumS1mb6nUOMQkSscOQcD7lw0yX
kuByh2WnogEAdHIkDXrftXEAOU1D6mGX8W3GppHDsOa5qCeJi/PJB9HqolGgXhwZMTDDE5qRHkef
ipNjJ6nu3Ugg5CnNL8Ii2rC/aTT21GCquxJiaM08iif2aHsQSWTkvaG4w6OtexXrLEmPgs9EvqOm
LBc4GlVyAQkGPhzcqDu5dlFF6RkkWH/by1T8nfHLb+Z1XuHGg3D5VJMp1H4kYOQgriWPhIUHTsov
4f94gI4cRxV2PBTIWAcIwzVEf1UyIT5llJ/51eQwcRhdr2bJ9PhSOhl5pdAJ9Db4Y59mLpMlIiVf
qk+N5x+sHAMEK4sse1LHZicRFUvlp/VNyI/SVc6Bde24qjsyPp5Vv5dFKC/WrPmHte2CODHB0yKc
BBj9OA3JZPutg9qUyVDepM+KjsuZU0guVcptdHzHL2ARZSZe/abRNM7o74s8ntDjIjlGlKQZiyH4
Zy09oEpXoUu22plKGwMmv+AC7wPpYPJd33UrsUdc8iGPlS9G4fLNPWGBzLmyvYXIoG5HLgp2hoST
PV2Dqn3boP/nFlmHuXFdR6tiY7/KIkQzFNf8qZwjSKivIQQRnZX2XUAzEuvJvXjEOcEiAq1Lne8M
B17oUoC86kGWYtgNl+il9p++voEgOMAQZsEVF5q2x7bTXt6g+4h16DG0bR5WX/BmoIXF00m74Ewy
nfoXq04VXv7yzVnwBl1ewph+F2LB8GHbHINR4D4TmUiuOdB1cUe+qkaPFFYT4y6w/WLw+PPcTqvj
VeJIMvDj0ZP3/Hqph7CZ7OUjt3J5RorINaZ0KslL3nqWjx/Lb9VkXSP61dKURZO0TSgH3V+qa4lh
ALa9Gm4y90EnOz9ttYrKZegCOVsns16V32BdvL2m8fzzVdzjTXtpUECG9bokLVC1v3aCZcd6pGJS
2czJ87VFpl/I9sk31cX/4h/+KDjrTXY3NmABH6Ndoct8D1/KWox/x3JkZPT8pMTtUcLARM3Um9zF
Clty6LmxHCIGsB0HTFUWxg8qarULCL8gYncRbjh76yzWnPeetBlJCP2J91fUSeXqjQyb+gOmajeE
Zm3QtfWBFi5ZFTPBCI2im9yDkoUn/KQKIyMU5rzrOVx21jM8OlNHt+7pJky/o9Ck2nlzyawfalF4
CmaLv+gGNYaVXVwghN81YnY87FpIK4WLF/1H5wRR18zsLGj2fKixScQrtsBTRx/9y76nlABfM8bG
1L62s1wNHV0/oQUjDEhK0lpUAbrAUr03m82aXiSJE4JW7if4Ijv7pAMa3RPmFu0iGPgvQ2WPUYIA
tCqEnomoat+c1trBjcvPA+Xta7RF0fpoq449WsY95m8ntslJTZeIqcGNec+uGZExh6SibRAM9mqa
8bxWUMa8hF+aypnzC1PfFsBdidE0fb7wOVwZTgxjJkewuuPMDJWey/hFeuWMfOjEyFPjIGsqpR0J
U/rAvnfX+L8iArsbTrjJp2zmyEjjQowNNLYsNpmg0R6YegNOGKHS4wt81nxE4nQuJiXKq4hBGGWH
Vf3UOzBGZYp00vXI5Z/eDEJ/FxpONQzssEiw7m0/wqBwiZJVmGdQJ64TgiEr/mKgL5JnJVK+MBX0
l4bw3RL9HNspBhGw7AncOl8b+dQ4KOFmjPAbeg/g7WKPxWOa24k/EI98ZC+oxHn63mH54LPFKk94
ivoTRhoVio8G67+sBQKFCihGTceZMVET4cw4f9VxZkc3N5f/uutST8ukuLjPqSBfjs/KeIqCyYXE
PtLjF0kMaIK/0nqUtMlawzWe5DQCPZCBAopxsmeTIiiyJdSnoqqGt7UdjcKSacsK53ERL0GFcgA7
VrV3SyVdzmGzV+MOXAN6CBQMBAdSNHNE+MJI3Twgu6RH+vBt/uJnUTa9A2eq8UoiVeajSJsJA2TJ
l1kN0W7fvsuyULJMZuL26cJHQdkhCWZmdWhIPi5x8ECyg95Ge2sJiJAGf1T+lwJkbLJROyOIwxKA
I00sV95I15aIoO2PULDCZ+6z3BaLMACEq8tAx6moOSAZ9QSANgG12Ct4kQctXy1u03J3dJNVS1mS
zaWC4e+CtOceQEaGhV/1PcJfR8MSjmz2nh3wnNJdnt2hshg2kRqGCS7xOr8HUI7MzIOsv99jlJ5d
Lvb4zcEzQiAMaFkfsSPRUpa0f/AE9jN3hVAU/SBq/vbh2QKPnTzF7nY+pdz6f5ZP6v4asYbaZYvh
jx92j16Ka7l3M9AylhbVBhufZ41vb5ILdbsmR0nWYeWkARO1Z4VY1+UdHC2jxYOnuUwhwQkD/4HO
H6cKDov2qJrSfoa2BJJK+iSBnSiqw3fKfWTYh30SZnfxYFS6G7eYL0Pk2NvLD/qss8EL2NFmj5CC
QWj9GFJGqFP5Nru/P59EIwhAmaIrFG2Hz+BXVS35IMO+bHHWs8ALBWWFus9ko4RcEKE7hnz3xY3/
Qtoex+3UklzwciRIfq8aAStl6de0IHsaCKNRxT0FQB8UWQT9nNyaIA3YOiWPbtsT5cElNJq0UMFE
pjplLu5JdHua5F7G955ZeHZWXZ2vJgA0pqHmRjXjNaaR4CmTP6XCPyNlQ2ll7i1QaBrDS56frZ75
A2BfmwzONxiMwy4e9+q67LmPE5Y1+AjS4zpqUE0SZykrrD4f/Tct8uYtRjUtwIQs5NGxTmMnsDMr
xOiUB/ae56x5ti/uw1uOKH2XAU6ODUb5xDMx/tb0MmC8oeuSS3Fjz7RMOK3OQ6HGWPGmJ3sm8J3T
Xa4xdxYpEih2TXUSwV2QfQ4YDVSFaQ0CzcnG4kMcsGxQfiHWYwU+iWSJx2+u3zP8kAF+i8mKbdkF
XYIEVGNwez+G9Saq+5SYHTpveIPBZtLp3ST3o+mJgi0B0foq8cr1W9Ij8WfIbcUcJWdJ/TRd7L/E
0LXtgAA+4CRdBkQIlZO1gt8IqaNCZgxKpNPP3u8ki+xTSiMPbwZbqaWlv82bY0yKpqjXUpa7gH2n
H+HKehtvtsYL4mNE6t9V9ty9sE30chp5rj8jy8/6Wrd1MS9RaAxZRPNry1wnXOIExgjD62nTKvxW
LfsnjUCnD/UZPJYQTAohlyBq7XMNvNjsaTN6nQWZgn3q11JV/TV4tJBww6V0tnkFUSf6cgtRRsJ8
sjiIOwQY0qJK87Zki9zpXVp1GArFv6MYsq7k/2RUOTE2qxdzhANWZ7oLBwy5oHnQdcBWH2NZiEem
+Cet9NxDCqOOGNEun6uNTUxFtfM0Jm8OieXY53x6RdcfnSv4EfphPSqV7SYTU5cgJxNE4bjuOUBd
074rb6O/1y1caAjwSZMpsUejUDkZ0KHHO2TR+3Yy9OOayOMwVeIsJ3D5TG4qW3pFryui6Fn0bqSc
Gghujb9eEO2+2XSgwTEQUGnlBrk+7TFVCeSY4a3KQldNvx7yWZZFUxI+yGs3fm+coxvQP/6UCzZl
FoWEIRDz5i4aFv629soufXaB+rAOUL0OZkzmDRZaLWVpBB1MuOmapFsUBaoAmWfntTyETbzSrJYQ
HBmztJmRUCIrBJxSqAmPgmf4UQekvj/Hhx6c0jhOpcOWw6QvGtpcdkCJ9/f1VT2d0cbwu5wAGhjZ
ybP4bLU8N4QfKJCyOn+pz2+f3QLWl90hbI9kMBYCQsK84+LncE1SgjeBTSKJrv7BcBbT97JJ8QyA
d4V5XuVcdDkNiYefTk8t6RKlWjULEFA61F6j03JpzOKFBAG7GT5zIYEWMQaZXCihDXYr+1eXESvA
Lykz5blS2Hyy/IZTfwJaab9zvmRknfbmm9XtZH+FGSl4bOctAU5DaC0p7S52acUCfCs/hsRyB4Jg
rjCwr+Izf5ILTWdlIKK60BPgrCqT5d0Df1JNCv3op3oPehJe2zLgXlzK9eNfgXWVvXFX28TlO8Dg
ecHL8Xuxakg9kRTov7SuxkrUvhUnow5/cJSiKdzupOjfTs1rjTPt5/PXKRtEnBjt0Ju9aDQ//lgk
rd5kPP2SULNu/FQ18JZ4oAzCcExyjcyQGkNKNv5p07Zh1UuRx6t7YYG9GsA5ExvXRxcua9QcMJaW
WTNscJguQG8ZDRw5trDlOw855AlsfEMIya7wFgaxzxcDfMFgpdpU4M0r87Uifuildjx1Xi6OD7oL
kOM8Vn6NkQqEkQQ8Ete07Ff/q89QaBJSP5Dn42sseCtmztFqh25q6A+yipVoo1g6yeIjfpr8pMtR
FTaDKhOYkIf5Ta7dROEtqIEwo1ducjowpg7qksuKR15RK3gjVN7y6QAzgzB3lDYtEeV1fVZ4aDmc
V9+pyJUYl1YvyPzIGNOQXkvkXD7xT5VlXhaYcouMV1QyPSJmIH6W7tDuexEFCb+nShwc1+VaCBLg
qxkFHQaVBgGsJgDQSIj5t/sVBqTB5rCE7YWDUP00D2g9wRr06b5DCj70k+oZM8IEJw+kv180QvUy
aHvjwIdbKJ+Uw1ZFq7W9eyGGleyfQHLpco9GOP7tJBuwWDt/OHvaEzeMjGrIiPtvr122B5MPOB2A
qpo+XTIgKdADN53Dg8S5EW/ZAkjQEDr+IotweMIOeSRt/XGk4+1K1YNu8FMcS88AsbEZdZojBgQR
sV3dJnSxZ6G11jCMvvYk7d+83JXaSEjFNSXZ2mDm4E6K8KaSkr7k41MGvpmXZxm+L2DDa5IUx9wP
zoJm6IM395Vwg9us3U/JTCbbX3OSyQYkMow+NRPCituEuhX775AkCHTfLcoUBIgEFIxZYryRjK4x
E5VssJyQicq9TPZSMoYjcwdxnt748cGr+8T+uvkwfM9vWGhzoCc/pm7qyVrHN8Bfv14foohUdzho
oNIXhaWdze+8J4oHjKuhAg+Jckd3PMNVbt9aBhfNCOy1NeQCwIakDdtjTUoOm06FJ8AYGsohrCaM
Ub+LzediYmFxlinnkFt8kpdJB/Y/hnOiBMy5wX9UbPf1oogrB6wrOKcZAti+IwA6lpfvHNk1qLux
jRnX4UXGUXRVtBNa2APheR0mxVH9X3Q8WDaKUpphQPvuNmt1RoCLsc5tQH+iltya56vSCrYlOPXb
HK81ZilPRgkO44Hwld4vAvOw9LR15UjywW1BWIDxSLrlPdrEC1Y2oZ3DUP8dVp9JTDTspm5F4DgN
TBUMTeT4NdmPNbyvhA2Usk60j4ONBslUeCst263vdfpLpeZM+wPRZDTYi7Qp9ecUaaCdw5cnmUxm
tzy9K0P0KtncGMyaYWmWfJgu5GV2XRdwIfggUE9FzKSPRCsH4BmjVwDMH8Aws6j4oK1A8Kz0COWd
J2dB9Xw/W4WN9tOnOlUreycbim/Uv/y1WqGLnfebARRjb+ETnYBSndfz4PvVONlK6ASX8AgeKXCE
pdrL9bcHS6nKM0fmlWFdzVpcvJWMp2rEs2PKABEjrOpJP27QC/A1acFzE2BX7JTEiAJEEvLOWa7f
mBsMLYH5FADRqWk7qtJOuq1odxMnC9IPrFjeADEYlPnc5sS/eM8a1vqtVFloth1WPIRKwlgMnLSM
n+woPV6neB+2CHJji6CReRyX4p0XT6XkR9vDcs+7/Bd3weF3VFZtFKvI9N9YXssIc/yjz9jOm1fv
aCcbwHHfjmxzgrp269tpLBEiZFWt039ug93J2DvofgMVS4S0HKmAxUPcz4e2PqZl2XRenA6Cv1WA
Y2PsPM96GD+L/AA4f5FpLdGu0xXaGQ8RlIL4xxBGhu8zVe5h6EXVhODvQcRxZHDmcNYJqoSDrnBi
PXC4PX8l+oPRwTUQAeJnASngWg+dVKh8DEe8KEllV2ml3VI2C80wQGk9gOLxWine9rkFGVO39PhT
kUg/AQbACYBPg96OLS0EWk1kB3W1KbzKnxDamp/rktljt78q40JiGf9hmeMqIQ2rwYV6lv9U7fyu
AvIENi6+7C9t6QhdJFIWPJIFeCOwhaOHuG9luUot4Z1ikQNjyCQQ0Cgvc1k/AHn+CesRk8JlEOSY
zmYZhPktsyfrw8fc9YTjhxcfXTHZsd0G+0wqmI1ozE64SWwlrnUVioLJZSkBQ78AFgiZGU4VSBJT
kmiWzkJZjKedRz7vjtaxEdRcNXuVrZW/vSItShuNrVQm3Tu0vNeHtG+AENKpGe/N4eRhsmDt/JvU
h0UOU4W2Ya90xfpRlk3dJ/E9jdPwv11Lz0oB7VrvJQ6HRjL297cLeQx/ejA4K/PQBRrtrJf5mi5/
TPc501YBJ5s2iYDJ6gxiW/A/ZZ7otExxrE3vWhSu45ZQJZJWjNsvPrA0Evtc5bb1zfC3q+CCYCY5
L/Yf6K1m6ZYSt2KIEI9+THgkXUz/c8XskpUfSdhHqaiHprC9KLU/5ad11+JNTU2XHu1R6p7GFiPP
JJ5y9mTHH2sp1QW69mH0dorWwNQjc4X68dpX0RJLPMV//XWv0JJWd/sPrx0BdeX5Vtp3PFunmKSU
iFwf7Toe2QkeP7vAQCUc3bXInY/zzV3YoJ16ZTd/916zj9l9Sq4a/DnAb3R3ZE5+nk9BQvGcMtgN
0lKjN9cP4UyOk8XMXUv8ZpqkMBPrMwbarPvKyuZTAAe9xaeUoBwMZhGKvtlZllnTbD32AlCASDBf
+i0IZTurVxETuoPC4jVFR1U6DqNNZqFj9SGvrfa5EwOrVTgxbQdHBDo3xEzzfgL1lMUcAQ/UzxWt
7JcvSp4J6ZzgbkWS2GoTGfFPicfG/iwYeKI7J7jAnAi6tDNerigr153xCreFIVkpagL2jQfnrb9R
BKKsC4PhMNCg2BzauoqQm3o7KSSvr+NiEb130KeODePIm966MRw/kp7AiKuUMpYPLfr4+/BwIJ8I
GOQBI8fdQDd3+ba8iqAa+AP4Pxy+4PDpEZM7te5wGj5nLqV1fnzAW7XQLWbDfZpBj5lUerSlWFDJ
iA/CTMPEwa1Hb8haC2ta6wiiJYnB/XsRXpWyyZlYzi6V/i+WmaPMTU9K1H7szUuUNSKWRkRW4llR
PiyrZwDVlLeSU80+oRAXp2bSvoex/6gr0ScO6TNt0J8iKg+RlOOC46f0Hmz9N1UpqKMXtR0kVMeu
5yVuHXF9qUVjH1hE96lJTxU5d3mF9A+L/29563vMckxC4CcEN+Sz5wZUyvkPx0hj1yvniRfTpaZH
ZTj6J4u52+FcpVixOIz6K8e7LINMhj5UoANHAWmWq6cTJDBc94Lv4UOF4nd/5auJ6U6gSd3TuneU
aJbsQYsHUyF5DBxYOI0eZWEvsMwKt0AIby04A6VCetmxDnOYKhMYRrVvwgrVELZZb0d9Oo4j1UUR
YMktQ0zN3oI5Q5FZGYG2NZXUmpKVCOpcCbTNjuK/DrhSSo3JEmwbzYNWgbBhKqy4oYUZIUto2/IJ
hd6/yrJj9O4z+xL0DJMMkJBfWSiBr5oD51FOfT1VXT8TDqLHAIXizZbCq4WQSlpKJ9kT+wmtDlai
RSE+Q21zsAFG7RR/+l7fTtXSz37SgbuT5NM0o2X10sXRdJXFs2y89Vj/nGwOzDdQB/hXqwI3Vp0i
OBnamOrV80W6ni5tWPLZwZcsC1AkXON4Jf8hHZQ+rBTHggFwZ6YD8wftyWmoyZTxVdvi42k38PTV
6juFxleW/OQGdbJdvcon2+fwiCdMcmFVNzjXE5uFd/LeZZWjk3/ZKsRE3WPgqyHzPJ76/0Vivn98
rLBQxM+mrpMmDYbtS7s4jGKlHrhp9tpyeefWCxT666Fa4jQ0M9nbPjuz6Rnwzl5h7mdnVjzPSDd3
O7Iz95f2gSp5uPUxYStf/wjI1wc2hEmVaAjSdSB4ZSvdKznSb/0R+9m8kxDxH/5gfyW29F/pNxJj
eBILiuOgKhNGkS+Tvb9mQQmK2M4Wqpn7EJqLFzI7HdnNKHY1ZKOEXS+TOLQNjMOfP71qA6GJjp3N
HMJ45euwfoHxRKXIgq7nNeNYstPLDsq+ze9jqN4AM7KiOUGRYY+yT4X0UE1h/VlvdiZyPyQEFjgv
DesZLuHXrgmSS8Uq2fTXmiG7m6uN4kI0JGtf8Zc9YF4Pr+KUQaD5FGTLhj1o0d01X0+HP2M8F1qn
orga9JGI45fSpsdIu2Y355gxU/0XynZbTuSovIiEIdVynboZ+Pay2b3IiKzQixAnjiUlcrW7ZwzH
rqZo63QKzdjO3XSb79s0IPgknL1g0PTXSXfMMmlPT38RCjB22cAb0K3Uvj3Oyg9JftHdkvD5JHSS
aRRlv5RTClAtI0Ws67a65GEX9UbJ/J6CEO8O9/HTmMj7b7Khas0vuLzUv0mqGpylW7Zb8HxnRcNg
rMt0Fo4Df4ILKoOuN7wTDbXhSCZs83PlhVDsvTOgn/DlLaAwnyljYMF6el+QTTejvqAvtFja54Yk
xjjLNbIKPKBoaGV0+YuZqXfh3bmEN7O5EcqHeB28M9siARSzZ/eZRyO8ON174+ldy8hcy5iad3xV
Sp5OR+wq/Hh83NtxiCc9YmuVoWcy/ZuQp27uACtH/EL47g3/k07EqlB4pxt2yJtNdMRWeDgjuvdI
Tw256JaFkToEpfL90W1+J4UjwiEPYXFoQqSAqms33gldpRgGdD49lWwgDISRsLt5KYxDhEOOB890
qCJ5vKpVjebeskZkKH4IGmo9L6nuHugPhs4xL60yLUkou2oIrg/D9wk6PkDZBz2CBx0KaKVH3ogr
2gGUJa1548f7CwGeMW9FTXtB8Sm2gybXYbWfT3dV+D3nwdTPiJDdVjSICr+oV2JsVX13t5ZU9Szh
U+WYYqP/QVW0zT58XjA2m2KVK9rDObw/6pZCMpB9QNNoMAX7fG7/Wu7C0WA1E3ZVEdI7A+xrBcMV
pTWKS7vgvBXQa9mHL84PUFz9t+1TYEEZOU2nb1wDKxBRyOEUqYIjBCcTLMArCLlNbj1yVh6p3ztv
ifLhVCB+IelNJ5t7FLO7mPb1LNJ98cr3loDot+Cm0S0FFEJfHUcGWSCLzRzGMi9oGHKz/2Ns1t4t
2Ju4q0xftn9cGPYEZ/QnSDZ2pUfhxCnCPTdueI8bMhXmKM+5IdUUJzp4Yupojx7WWcZmIR637rw0
22gOwdekW6AWKshbqw0wVB6ICFiohvzTj9zgR2d4fGSVEiUV4Ptm9Y1fjx6/0pL9MmqNAXyPd5rx
gca2SJqP3hJoo9ptAcAvTGrhmNT/4FWGi2vmCwG7bfZtdDAhMm2wXjM484IDP7sLoQPue2sYuTBk
HPq9ScF7ikxXtzQ4eTpW1A+mZ1yEdSHwITGl6Gu9dgTyQDhY/8dCZQbxN59xsKKg93S0ogFNYq+q
Qu0AwJUn22hnF6Kr7YPEH7D7T4DAZDDa2q9Krka0R3yRLtE0PdRmAjc9O12fiuk8TJh06/wHGCNU
4wy3NGd/S5xwIOI25WyzdYdpmAY2bn9qrDUor7lYyanB74Wba/RCUw2lr5HCUyugD/52WNuGiBEd
XRUCTmln5UFIoTPQHcwu43g8SGa50SkTZMCHctq2gSYBBad/LRbycAXHKQ7l7OuDHpCi+N0QMBze
vLTZO3lL0VF1t4fM6inqx8Q71EXa3ap+N6PmVnQRQ+MEw1odwpaid857lZlNP/WJ/9LJzfzAhvOU
xUDkFe9Ql22IQhvtslrWzyIZ7zuve3HAkOk8GGbThlmG+OXA7tBRdHjJW1egnSe+3DnCW/MLWe6h
h3nL+bA+Q/ZXb0H3qR9M+qidHSu2umxLVF/9E+W0+GqRP+vsL00i+cu2DLDXPZuL9l7reIJu40mg
NNf0NZayzggBCaWD2KOoQMo/Z8Fwd2V/kz26gIWAQplsrCAvdAXKlhEwO3e+67cm/59CC9ERr8H7
hNTknmwQiTUo1eCUGr2IPz3wjSzbOFK4ofnxw9s4DWl6fRNvRJd8he7DE6jugTWk+P36BP0aB5u5
IDg4HUROrqlfslbeLKv/nd/R2o/JZSuC7B5k3jq7xgWiZ8o035W6VtuTFHjZVvthzNvvHaKUb+dS
tG3CoCSGwFGOhZvcuJA1FT+A9mQDBkBAuYqGh3GqnrcdI0cvxH49p3qtGUitpu8bHd/0QXHTJXdD
OsxF1LwFHhdgJUfgro7NLsSB7sooR0ZciYG/NcbKoX+79GEKDk8S6APt7hz101ovKCOxLKxBKHPY
oqG/5jKde+/vwtmx9TePwzHuHg/+/yRvtHn2WO4ANxbNOuNU3HtyMfcxm43RxnPze+4GHy072JcR
uhyMQTENPjWPNUurXotODP2jLjF2QtwN6L1fq3ERW2FGbpApXm8iTD6rNFtGxkFIWnIQ5QylI5kZ
iD4E7BynOZvJygL80pfr+OBuEtZl7gb1/YpDqTm5QmQ24aK0j15C9+PALprCPRGi1b+QrgpXtc9y
fXVdp0cuzcUZvKknSwXXbt2V0amQJkK2eps2cA2Qwy2fNKfgM2ObINSay0nY/raqnlIbsd0A47rz
FBU4wamwWO7Dxg33CKf6btvTqShvAuEV6+6zJJFkyye163oh8UE1CM6FA/YaAVt7HQceMaPe0Zu4
28jI6XV/iXDQTds9PFme7qaYu3bKGkrQ2mOyBf2c2YtnwN3T9tb6EiPf50P/x+AfJUe1HPInbGw6
MgShaHpG75HDcBs1owdRpWyh0EbgD+lFEdfkzv9gY4ke92oeALySNz9+J1WaN93lfbyi2CwZN5oj
7FMHPnZfGpjOZWlFgjmdOoPhOSQqebEiwv/81/VY9lj5Kokw8Kjy7El2AZakzRgaFwLhgJbUrhbV
W1Y+C5WtXvWhuB8D5NFsZLdOp7vBezc5J+oVYVqNrr7dW5HKc2MfsylfkQtBty6NHRlBCxq/eDps
Pjx9GOGsd74POR0FGL54ayxwtk5hlmPjkZhSxHhcaF7ZzD+iLgOnKsQ059kBfX73cEIi3QVzJ9Cq
I2c9dDS0pHuYY9NcSgZabVLs4ZJY41MI0vfby/Wuamy7Bhcpx7762hFS0tzYJdKkiTQ8fgt301lC
qynGJks6bfFB6RVD9ZidexmW9fKZLxfEWyfdwk5um4atA6BZFjLT91thva2YaIU9Rdr3ZgRhlLzz
+wTO0p6OjiVfUcL+QC2vdONL8Rz4kkullNyjaNkamb+n3L9A6qr5lm8Q+bbcl+PAn6NX50XGamL9
iRd3Bgtoer5nPBPduDPZI76qQR7pOz4HlBOtb5pHAI6qGuFIBISHicUq//VDFKAsH1jcZ5gzoF+F
yT0BqGUAvQN2UGq7nfw9JtkuunLiD63BzkkP5xC1hXR/0WbAYzSXn6VsBYZBes7UnG4g5Zy70BR8
ksQOxiJ1FNXMZ2JVKaj1lFM3BinCJy46lFNG28tA1sJrXdHuJzFeCFniOiJ6UqzN8mLqxOBerh30
dWwtzTtLwkLH/GgGstKe+g9CVgegzeGYV7hvFMNfHd2B12ZgvBqaOZkPuBgSVuWRwuvVjPYcEILm
DLJdGAg5A6HyhdquyObSLlsp9XXgiIWqptI7Yya1eNsYditKBkQl2v0SXRy86crYsi3ZIlEPkJXu
IGZKAoMs8cgebGCrkJK7H6ZD6kD8uR8MUIG4c18gICTG2fybogJL7s+rTACeEscH/Nt24GyYUrZW
Kp6jlOYMTON7mARqWrs0JQzT/zF8OYbaw+2N3GjnguJJlenIewql6/6h9TdI75VMp59es9YnoViM
ZbGpZt9YCn6qeAwWW1GbXQaVAxtg2aj1eESRErD5ZZlCWOYBz4pbz1+sQ39ND7aIHPXVLKYJM/HJ
EoJlFIqen1AvdVUpc4HFq+ziAEKw4v6MtQ7ixWq5BGa4WLDkRbITIbSycEBWo0HiflUzPdyq315i
6ZCtPSXjp2yYgFWDPD+8ZrbuOYz8pYakVYFbimEKdb032ybQoM8MtyRIu5dTlxkXz2ishQDbD7sS
9T0+floyJ+bF8OFVHn3uVs7lJ//tac79xAEWgXzVgIZdrny5pSs8ElnW0yHufA4CggZR5jIp8sTJ
iPXEpNUA6/rusm4BmRXu2+Rb3zv73ZBDIuHoExgTTPtyHNfmW6UGn2KN4lN3xYKqBHOCjpC/3P+v
/AC9s1xqJZgLEeKBvE1Z7TaPwz9f0Fgszy8bExvKiWUnY8It+tg1m+xFYM1cGsIKEtmQIAImyIyy
aASQAwZCipFQ2793EH7KT3QtpwIHFO34Yxt3mFGEDHTwUudKiqmbKM7c64udim7YtnJxZbJdlZ86
wDOyaGPzz+opwxqlFbeW67DBXWKolzmGPzBVmhsvTwTZjU0R7Iu5xxRsT3CeywYvZqL1JZScdCoP
2sKTKba3aWb2M64ie7zXZ4/8lE0ROZIuTx6/PvezNTx5pk3DQT9i6Lg2A7RPSxq7bvTDQiehmbxw
5LOm1zwV0UVOQBg59+XPSUia4AkG5kmINN3ybWzDFMwdO1QPj4dfcPILSpBNWR/gSxiBaHx1gv1G
gCzS1gq5QT/i6rl0oPD6NeLBP2G/tzLOnSS4Ivx2vgE10q4H34rI/s7Jn32BBjyAXNY4u4dvZFtQ
KF/fR0m7jjAt2aGkBc4CdILbD3Ht39/k9aRD8mJ8AVv2Al2sgd4EOsalkvn0gac84RRwa9B1rjTy
f7Mb9jnoFVsZ0sWmxLWEi9lhKhTy0PrGlfWjtZ9d0zIXHdwv6LWVvGgpTeN6fn/zIDwcBmlal3FR
9xytrdHpFMwXSwFDDOI3SBK5jVPUdwreJbPyVE0dgBO8X4ROMd5aGsOyQXRI0WP5RYoGVx7kzcN9
kqXRis/tpmuKPMWtadnsnCJX4mWyG6U/T4oYJz0MvLK3KGg0Z4XLKQXl2FGb16QlnQ0FPE0ToIIu
UlY3M/sbC1YoAo56pJrC6TS50sOt1A4CW1xAlT1Wj0Sd0hew/On5rURnyTX1G6FTyqXZadMTi6FK
TZcOS5rf9w1U+SLIROo4peNDY4G6KUpLVWRp7cExOCf6oUmVueHTE83cIklyM5rs2yZjC9UHknr7
ecHB9Hsjwg7cKquJMmdtMojx+RbuDzHpBozjoDZYSfQBl3eZMUXA4SMWNrxToUjkoi1D+ZLxRmKn
Ldj7WvIxH0ruuoyTw0P7Ag3tZggMkFWXaY0T9uDjj0xTm1lJvpDSy8MMb0do4mkB0BywudjxcdSs
LynBnOx0Vu2D560QL/iVKstZ8dWA20sFNMYprSriEl7WvwhZ+T0jNsZpBljD7mp7sSI2nVhrKRVT
Hxpjv/qnx88zSaOaOW6y0nF6z0JeA5utvXP+DCUo1jvX9KEyVUhlJDpkT9UYaAki8KPDE9cGrGSv
R3a7/NAOHxJgl2RDArn0MqpQ/Bd3EuVh0mcUhPC+Cw/kJCeFslUQ/ujIgq4ke+ktCdJWlin0jpp8
llDt/rOIs+45CVmFQplvU+ALpVORKOTTJN/EPT4xBGSzRy3YJXBDZZuBohuXx4PExmq7mZv3grrO
xs0Gn2ZjDXF3/ct9CihdFRmqXzc5cOwEmk0+3A53rIZCJjhqHo46MGL6QqHwMJS2K9VoEDEdmGum
8kOrScTLSJz5GnoS1Yrb8FWTB1No77zBFgZEOKX7Z8F1uDhdAFBUGAnDxiETkEDY2vocLYdDGQ8R
3Eoh3NLhrL7m5Bxmu9FdPRStngL8SN5wSMDTCe+YxQTfDQLg/6URGzIbVo2tTMkbazEQG2Y1XrIS
bSOHHBoFQdMfaxPky8/Uk9LtwUqZXD0+XGSq2DKSrF9oeGfeV/4g4klS5ttYqAF0nu+6vbcpuTQo
lnhoQjOXbCXxKOxmxPdDXjO3LwREeBGFWH4/a6C3GkxV9BR0zFDB7vU9uCFYV2fVgwHwn9T0/23T
ERV5AspDyq93Po8dVg5NKkHfpABNH17w+J5YP1HVIVM9nF7UKZNiztig1HJya9QN2NalmbaDyRQf
SLfWwKjkZFISt7fgmPoC4/+HBN2ZdehF+rq8DHFnOi6THsMYhILdQP3eavvMXIPyeobmEDDfdj23
6LtINi2f6jXiR0Ix5k43eEk/KxZzntJZfA8r1ugAYn3uuKzM0pi6YVBz78Bf1fyc2qozOEYXunus
lHLmXbbphT4Umh7ILlEiQetgYMrveKkFpiVZbLClzdl0Tgc9WjCId2Lw6qQkhZzs9kdlguoxrW6q
zgYmFVuU5AxpBgGK2VIo/mJXmMGdFMTYocOHsEGYeW5p2m35atT+KjWmsk6+RtXPO3ImBTJFR5YK
kk82PQFVnCENs1MPxOTwIqlwe/9C40B35+pA/txFrShs6kCPotyxjyaaWpKuWJU/fvU0IG1Epe4y
uH7Y8SfAxKKZ3fJlPX4O1tQbPXccJ1HEHo/VqDx6k0fZnDv7Y/M0ysOUY6FOcyk4UjUMLb5Qc7w1
RmrANVX6xf0jKy31osA7m2xL0DxL26iYhHB556PaISFSOo1jaZO00udJAXzelfm6ycgubuwJsmHh
GJZYScqKkl1oWs7ovuwn5n/2b9jm3Bw+QQxkXHBI8e4bGp2+3w3LuRY4xt0oOs6/oIq4+IvUYYDk
D5o93/rR/BJcoO3rYXlPFKQbRNpcDRblrnoLDaiZ2IUmgDWxagW4hDFwI7dgjHkZ/EgrJyg14JMc
eTfa3KrUyzWIwfPKAGW9oLGZ7orw3GfHFLf26SBBboum2SmfJ+paGyKJyrsAiOpM1IzY3gpKR88q
XEQuwrHn7Jc2OPYMhTroxOdVsoTJNwoAop/a55lIHq91wiOx+U1kXwVdLsZyHFE21rqHT87q3sZ5
qVyyYRvRyx2Kgf1ou00UvZm+ltklQQfuMeMTM9W+sSc5fELUcyYtddNk7NZD2SlXAd58D+CV+5Hh
OsooJUgSwnvm9HEKhj2BUJjdBBfB59gZc9L58Av2LO6a8onQlz4zLeWidHiubwlneP5aqE9Skauo
tGC4ticV7Kdj7x9RrKp8YC9SMAQbVpePBRW6PoP+ntVCCGsYgMNnDivUhQhTsJgzVX2SpDahtEa7
bhLtW2tUVpye1YAk5Op4hmZsJEurMZDRbH4IlXEQbNXhvF4zbyOkk0mWvYMcz3WHIL6OM1gYnzkd
GuoJyoquvEBx3sjf2Z5g/Jax5Tk/iIQ5tYYyBWkfpN4fHoDdekymORMiUzjgbAie0i44bVdSwvmQ
pKkRlGfLSwSXbgipBiZPRWtPFWxgrhV7+88Gq6nB8f/4cwf/S0lGTYTeWW5reDqKEvjTxZPVciS9
+BnjbXCyrPg6/W0IoMVkXKK4+NwWtHMuLF2jZA11q/EvyXXXWwr6BUdmJwSBkOsDFDxmxkmx8SWi
WqEvO7+wecS0tV4thMuRn/tWzhR4NncLQCtmbaQwrIFf2imEJ1JQeh8aFoTV0E0shMjpIcyAwaXZ
YwJDoCb5EpF2QFxiGZfnoZF4+B7Mcy+WY9sxJHKa1/n/KxeA/I0eBEdmPz2wOFTFlxwansnEr61y
j9L/FPSjFCzkYYfeDguhCq9CYi4+y3i1f2vWtl543Jtn5hho4ZW+Y0P9KUR9l4oIyQKFfn9ErOGw
QLJst6WqB+o2DEC7yKcaLFl/x6ARdXdI0InwYskzok04QwDwnrekANfyABdCyS/39o6N//cZdRpt
RbjJaB+79yn6jAGaTjfL8Qboo9Ezs5qD7KB7asrJYJ7eISICTpVVtOKwznw7q9c26hucthQKVdg4
AJeGAw64kDrrsb+OjWYVO/KrEQGqckjkF9kRRQXZPE95gXN2CmPw3UmJFF83dxPCEGQ3ArTb+Pei
ChhjM/YlaL50j2y3SvOmsWgxDuUuHiOaww8lNQhLIjEAwZH+DLFXjTuN8Q+TqBNEkmW7Ee6UaDjY
jWEUx/pPDjaMeHF47IjYp445Zjvk70HYCxqLH8BjlqCjA9NWymsyO2Rya07lN+0o1Qj1SAAN9HcY
SeCq7rzgtsmuVF0qfBojiCFuoGOMCrPmZ53YH6ezaoYWZ/b7MJEcyh7AygY35iaiklSmhn4WVNb5
034ktsVdKA0prmRTWgv/GJuRn1xUAPY3qK2trBWRygSrXFL2MRbAg3FtEFDQaM0kOUryvYpjA38Z
cZHWD0FV7NqapmxyeXT3dKLc9xLAv9SDfAcz2EfGAC83xPz8WALD2I6KFaJYoSUsez8zBaYPSvfV
RWWz16zR06ny8Zn6jhpDX+4lhHqMprsZX5wyMMKTS177mw0UFk0RPpr0UKv0y0TdIViWrz4cwssV
t2TwAtjhzITw8mq6QPhtSQhTKkgGPaooPhVvVfs93RLBHpAiC30z5lQHFNykE6Wjrhy8w41ROya1
taTNTcy5mYBMa0dvv9qSNTB3w04QSQnwvgxSNB3AT8jS/kyV05MWKQHhBzFomHlvG4+HYRi936w5
ifUmk1572TJjSmIq3hTlH3fva8vk2ZvRsc+CI7p/F4yS819cJfOydPBLfssE+B13TPLvKidkm6tu
tJz/w5viPpj0l8kaeR3J9TKdN7hBeSBxg4OdJKlZn3NEFTjBJfKyZjhpt8GjJRXb7A9xU7HP0j08
z2Iu3zqDpr5BmLHWZ5xPWpacDcn7LRIKixXWe2b8ALi38vyJ3KFYNBF9ubnzRslspXRNbN0IBBz4
tRrufIHH8o/CfM/BIPcyKovWDL6ZYVB3O+bXkzNlAk+ARyMp+el8KwvRfK0Ty4t8QB3ExkrxDrF3
otKOlTNAknztYJ9+wyDP15q5imSdNUuhf3dQh0ijDAoDijj//jvz1Hcx98lyToItSXwqtZYI35y/
m5TXLVUNzWCm/MpF9Oa5747pvPDFSh8MB7I5QzlBnaP7KABzeow0esAoo6TlZasPXavzfW4wpne5
wG2MZXkT5syAkmxyIfbowZNQI3J+voCoBF1TQWnT+Ux4zzp9kdw+7ykThooJ4ckljulnA70iboSC
HYhNyJSZG3lpQx33AWtTmYWWrUZ70967utk/4qDKLNdtw2bKNKbi+eJEyuuGYwDfLhxAV0A7n06A
qYK6pL/Wmp2IFg6afrZeO+2U0n7zNVcGZ2gHLw9mesVV3oRQaFnvbub1YoDFqJHaXpeHtOuMxAqn
G9EoXnGPK57w803uEjJe1gczEhTCLkAuFmBm7hlDT2AcBJKoHMsQO9Fo8Ga/g4FfY9J5s9kHFNkf
fLw6OU2uuLdeTqWq4+fzZ48k0r7lc5n2/2Yi5vYNiDRNntvNKKn353pwLS50Y48tlc0dFbUu8T+T
jT3eP755pfq/v/GuhC/7P29afevasI/dRSVeOjhdvF0NASTeGcnO8D9uSXaFGVxIgVVh+HbpgZ4e
2+2qFRbU3HQToBdqwCWD1JqQxKjiafOG8q8d5gnwm2ba3UMqGWop+4aF5BqJpal9zX+JQwQa3ZZ2
u3rLMsJpQ0JihEruQnPoPcac0ArsF9H8HaKdkupbnrVp2u7hPioG6KYq5bHHD+6AVwY4bs72rw2b
0YYqJjJg/5CUQ+LXji+uVh7QmwagziWBnXKS8zx0UPU+ENEVjvDfqC74ssP0307OH4+tBPRl0HHn
KpyrbmyPSsU04hQ0robVWDocjXsqNXfGDVTmQK0ZMZRtP5++Zp8v5OhT6UI71TDUCvi3GqHM+WxH
yRkWCQYunHditRdKWlM7ZHaeGtrpRziH//1PDPhbp6B2KBaLgOo1CvA8vj5czZhPJ1BUgXknplaB
6akEhBlalqwYAqeX1pH/XKeylbYtKcUY2ZrDz/lH9Z3bfW5pcC7YERgFBffxPj3E79SM0g8NIB24
E0XbHFE74oIL4pKnXyqt6B/Mw4ZCM8WA/Yvwqw9NRyGW5hFhwTP4p/wGvSBmPQrpyZldm7l914ol
UEDUp4dpWu7Xg/dpBrMLK40bwvvgAbIbPvZEDdtGt9P657I1Ol+y4uHwdALUxleYYOeaMX1jSb6S
7+aScMz2JR8LD03zqrV/XJf5Ntt1M3CcGE5cjxFAQK+/JoIkJCuBiGcEGQ/Si+/8SGr01bIPn8sP
825YRxeaxhZ4VLFLIrCXsnAEBOT/Pi5Px9Som5r1QBUAaPtAQltXT9I1rCAceDpuhImxHOh0gEO/
GZ49x4Ly6/HcF6xFNXx4JQJ7mm7Jg9zWygVTlEOzFlVC1MPCw5hxZ++iPeYBjOEMl1HEgvrKGhCM
Z1ne1RO6yiEPKk/Q0yu9PIUZY21b8QVeUvBREJX2yj7ZsVsZBwiwHhTP2qqmm7J0Z59QU8ylCPl9
c9SODOAA/fZRcDSQMxIXH+zsMKRjBrInO1h3k2x4envTtyHBMQU9gxDtfUf0uoN+ZA55NvS1tpmW
643pLRKgPfV13N8TZCw2BN8b+6r3yIz3uZ9fO3/w6TwOMcld+Z+UlE57nsDH0ObAr8dohUOZ8MkU
gvDGJIqdCoaxLwid8Y8QICsvPqKHKEB6Jp0LDfrGuGfj/6lAdz65auFg6OyqaXNUxybFjnqzeBBj
4FuAkuMswh015J2k45roprpGaHGJewBlv5GlsWjA87IKK99won5u5pvo6Q42Uj/TKG4s8O7kopr2
fy//r0GZVdLnSXX8LpdI4Mfct6DEt3E8SXKPCjDldQslaPVxHGyKUVO4125RhU1zlDMGVyWxKFue
bR8pQqfldYHJTROoySCYx0Pto2QqURyPhZ2uYpD7cspKXMTxIlNSEFBu57Vvd127IpgSw0QAeSdB
A7fZg8XCf4WnOxZ6M6VUjKOqVbA7ziT5fuXZPHARx7HxNtBkpX9twPDQyUXAuHizHV59cP0h56Q3
CoguueSnAs+Kmw5PTz+fqqjkuxmBg6hCAodqWgVetPX7kXOP47aBkBuEMKSkJ2NxeV4WFu4nVxaE
qAhNQhOcjoGqDU52TwX3jlEn+qbla/jL7c+blb6b+MVBGU68SKtS21NM8RGfhp+vlTHyumAdxGZE
g5J/sMUcOPHvNyZGSMdh02aC2gpSbmC80t8iquXdpBBMBnIYKh6p28ODOmLNfJez2UHNYM09/CMZ
AW0ITvpHAO7iauCcoJ0+kpt1w4yLCxzHQss2nF3tti9xQdgbH89f6yg18wvjVcOf2qr7v4mDresl
QOOk4sr1vuCBVKg=
`protect end_protected
