`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
aw3gwA0pkA1KM0EzU0fWDqpDBmki2pv9wCQV47fFme4JKsq63WG+ADCE+vbn7Hi+Z3/OAuKb4EEX
dGenh3gQNg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
GigQBufnZO7EfSHP0Y6uevwpckWE0sKJaS4js+xivY48qGBeSuRBIXwcnXUOYHc1ZK9okdNAvJwQ
JPNh76bftVump10ReYTgvWpCGfLwjQCmMQgfqzTuUx7v6mXzXkHNM3AF9yPZCD3vpvtPZgQmT472
s+pvZ7tu9fma2LULf98=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
psR10jh5pgqZ3xweJkjl9fsr4y2yU1lL9FJOcMraSNIpnfe7ZuXdAFUVc4ih4K8UlWax/IkXIlFZ
n1Go7PXhFKnwhLIovoHM5Jvl/aHMnonGGRE0o153utTtS+2xjpe5KLXNZCOOZkHt1iYsRJNgpalq
Ec60R/l2o2rx22M8MV2QI9VH5n6uir/9OOojjQSi0z76+QbzIix15clS2EM/KdTtUZ3N3oc+KXNb
M0WVoI19ToV40VprGKM01OBici2WucYGjiFP1kyi/Z0HoPHzjqKzAbwWnv2tw/U5nGwl8XzHIrqB
6RuMYMosIIDOeLH8KbgRiQ9dk+eXqTjkT6DaFA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
I33xl8KW5axmztpTK+QsmLAzENZuPcE7t41lhXfih+wjvg4ilv+yHoFmQGqQiA5OM8uI3vYwC4AM
uhXm/XO4za3bWTMKArTaogU8bQC3ob07Muh6+PRgnAPkCENTQno3WFMqNAT9VF4hta6Ms0fm8yCH
mYbJdYkWwfOzPCaNq6M=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
P5FwkKjf4Iwwox37r/di1HGRbWXhg6hz9YA6uwui7LGq8dcYaQkeLr/GG5TGCrlD0NrV37s2LSbX
7AfoQ0uPsN5S1snAl1OJw3RYmlGpl9ibMHbUN+3sJlFPQDBKtau5bG83kELMq4kfchkNasGTpkOE
dRYrbcvCIB/P8mfl5GpFxl8+QUwKwaWo0q5QQMl5zM1EUknMP/KD/TxvLLiVnpCvfUu8LhZGlPzT
mNjw5c3aMaPj/h7wJZc3woV3ipM+9dh+PE9NoHqZbgPHU6murBnDmTgvuL4kJuWVzDB54okyCb65
ivdndVdsfQ5rKcJcHoUkja+vdOnP5oizOryTpQ==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
CxoPsRKVWfSyg/9xz4OvBgE0/+1nmJV44iU931cbXYa8QCvRGQyc65x4pNqQX3xCsYGV6DapTCDt
vD4a6ao9+XAXblO1MzjeCgQ3dR9GgRVA1T40xYVGduF0uzm7xeFtct3ZQLoV2n5EURYqM7Lthpkq
m14yKvLy83eQwqPDs13ImaOVXdczOU6xX3ynkh65ShlRdsloyxNGOfXYpbb7r0IEad322Y3RP6hW
wacfZyIi2bmjbID/rU1qpxootV+r0jgb1/wWkBjvG45gLFr2NH2YbBFOr0w1OHD4SOYw9RZ+lPa2
/3iRUorjuHYcx/D50YSrKtQNMZZgT3U9/nU7hg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5872)
`protect data_block
VxqvZJEyVHWi54uYo0wJOQRTq7DwKUbpldXTlaQcVwDM+pfhyHh5WRy5zAFkJTel0iBIO+2lAjTt
Ug6eI6Md2Y1kYqM2/TQIVYGEmXXdq1LNVmAsIrWGTGoO4XLP+Z2Y7HCLlCcY0qW5mrSujMB03eLD
hX6gu+fy0Ozly1zL2wWfo8BgniAloEQrUDTRE3+8qZBrQEdWOjI5AMTfRJzO/XHISu6o9xSDGXUg
l8vk3lRm0Ylt983mRX3XoR3rfw/PC2E0S5Lq+hZMcL8osrWjXELP82sl1wm7n9o4t2C6uXUxgHdQ
Ow9nKIQ4XISBEhLh+FIC/AG7S7NTeF7DJn4yI3xEXXosenBYGTcBl3bLK6Et/C40exQNnUgezMva
WJxhPQV+ziQbVDyBV6RRM8mtaVyTusKn1hSEcFEV+k2n+zaBHLkt9iQGLnO9MX6UN/RVbIo5vHlQ
crRpNzASJrBdsaFm9+W4h4a/k26N5OjJvQf7Gl7dJJVBjU7kbd/toMFuREGAkNank9Db3IZN/sMV
ha0eFlNn1P6nIyXQlVRWHL7sqNUBFTsTzn43+2GjW3E05qRSeEoMRHvX82kWGakTmw1Ae6ABVM9L
mghSZAUxWHC3v8wWJuL0YAaoYMJetKrHHanKFvq7kAQL22vaRjkDyn7G+xW6pDUlxc5S0O+qqfyx
7SXdm/m/s+IlrRK09pRCNEkyZtk+jwA/GxCIQOUAOHEuJJUQ+AP56zOlq88pbPTq6IRleVchgsHW
zmp6O7XEBtiUcHDG83xJ/hnnOnZFYvHQtGMShHlLXD3Uon+2DigcgyFx0KrtwRK0Rk4CTmIvNm9W
HuLDd2ulvHICvHgRuPoqmYkTe/21c8n2hb8k9PvQhpR90kYcuy021Y9psF99WOTbG3uZUmJJwpQm
9PsaCLIfs6vO/4xMvzhIi9dq3f5uHdrDim49rRoUNkgBwv6uP1hk7Qh1wMBynJO7ihkaz4I4t8dy
ZTYIwAfIaF1QfWPM52z8iV26JNlVc5MUOnh1paAnbjFcSjYh5DIORWZW8VDC5AFSptEHkkVwB9if
+sbkZ7wYw1lCJUDii6pVxnWMgowA9aePtdrRaMJtrt5993W33aIKoGXmJHU7V6II6OR4zx7sGUPu
F17VUdaVqPpHf/xE10OqyiYOozgosEv/6rM6lc4who7g4c9d8MClrI0f1I1JCMHJ3RJXDMzHA1+b
EOOh6eTlXKrFegvUf/cVRWIc+xbR88/jvdxIyYzcOivoUWpyPKeNjxThtoYdJiYmbfW5yz9Y1tSn
FahNfTtiBzdIcdkjC94cPOq3YUi2bhxBBAUVPJhZwcQNhO1ZuSho5ySEouLETw5F2Jyyc6OjGAI+
8rMH3sX5ZjHKrYiJr9HdyCS2WZAk0vUwm7d+ZBWH06t+NdE3sWNLuE2m4VthRlP7U8pW6zEtxsGj
kTMVCjU9+7cQxUeRDPEG56Uq7uAT2xwyvpt4I9q+ob1radL1xaMOlRuFJxksa1h1xTo5cc/Oy2q0
0vrD8VgPftBYssAmbI+9/qDtRxjx0JseL7y1PS1TtrR5gOYE0HDcY1i/bj7XTZVuFM0aNmpD0zE5
SQAeiQziIOk7qP3Zki1WpbU/cVZe2yk17xWA0YiRmICIub+8+BpqMNgCIbIAO4a8uNRE7IcyvCjM
zI8hQDSAP+w8jy8wGbLagLt2KejqTtkwSdrsxbNnDcZt/rfAAIsQgQEJLPR1J2Rj0fOtkuy5FTsl
Dz/sDXyshJHJ+uMa80K3smYTxooo9J2AB7G3sLmm2cp9zNlulAl9clIbywMJs22fAPyj1MjjEg0L
qruYygiJ+NYaeGfjAMLXPWJlkhtE2kcTE4Wq7ETbm4p7Xt4Dn5OakdZvM9FF+so0tWjXJwlh+0CJ
mrUxi8GwYR15+QW4Twu6wAXn3q6DpRDOdMMVgJm8KYBIozmu8MiyT5666GgEMGKo2AeK2EFIc5GP
52bkqYp9BNPFGvMG1iVZojgmrvN1ywIVP5fQKJsNMUfycX5XptiiTAOMMZfah4jz2FUPVXdyl0XO
SERvGfLBAKJ5S3yis1o3tvSGTb28EmuqNpm3qfiSNWbMiciYoptfcRcF9hArvKue0S8lILYYq1kO
ZxQCr9SxcTEh4zTYvaDfcagYSr8Ltzbxrq8/PRwim+wErERSETDKAhuM8wVTURxSWBpYWLP3jEqi
SjffgfSfhKiaXu/oLtXUv+b+aU61Z9ddlpxxs0qQ58GZ7Lwo8skyEjVqjQLkSxfJ/q8RnmrJi4xJ
rtMsWHK4B0aOE0YzsVejWJqbDWVPlCT/7+8gvgeSx44IRNIwgCSjrn04fmnUMNIGH+zLwOzMUPxH
b56u0RpHDKugO2Rr6wTDoJPGi4WGS6EpXOGwpfCnKutW5qA0U4D9l/Pk5vKP/T302EXSXqToKuX2
NVaOWe9v+Pj6D+DHeYKDMl5+TndMmpTALPSJdnRj2ln35YpriMT32boKlAZqy1zsyQbTFVbFfUar
rgvLqGpnzEut9gnWXx3hBb0psdiDHkxwPCcHNv7NPpQPp4PlQblkzl2f1JUddqjh25DEDUsdbAT6
ppA5Eo5cPlO9NuOxfzXTubXw++qQoF9fQfkoiutTew+Q68BYylxF4eOUtsj1y+sjHBTuleOsvodZ
tDs8bEiGL+8QYJxMSw8e/aPAh1LR2wwj2AzGQQLwImYlgtuh/CBMkB10Wta3yybSzUqIEJofUxrb
w05idTV6VL+Y8qzv+Angf0hxSaSlVNKH95Rcy3qi42SHqE63QEqxbVE7APm6JRrOZgUwkdnnwaaJ
E7bCXYdolSCgq4CvfjUNlksSybJpd7bGem3xYQVmgpRwL4RZTmSxeWK4DeX2VmDX1xPzK6EcR8W1
G3gOwJLN7scBHqlSQ3hWqrwgV5UVIUizMXs1aEYO1ydUTpdHQhg7ooxNtkc6uTN21yiqZ6MyT0u+
zuLWILmBv2nRf2Sx0eu2a7OEvSWYykOewtWXLdPSw7zzbeCLxQTQkaqD+syKxLYvsR43ODf6WW4r
hYTYk89C7gO8GCVxuqFRAdpZ8T/ZZfmD9O+//GtK92fxXRe4OrvMxljVpjYLK+gqDbH6D8XNDN2Q
9HLZm50kSA9WY9xFNUAwAwNveFvdqIuVafZzGVE1CK2/fTp8WkHE2h1man7m4mTHXxacq4IoCpDJ
Kzte7eJQnqBnodnyLD3tAL3s+5A4SrOCvafJdgq9SxatWsx5Icpnp7ZuDxVa38FqxOqnSSRH2hjo
nO3YVe5lmCzKmf7IW52/IZibaMYDDjoLa4qpg/s/hqBUCrAScwfskbnCeby+DB37GIDiphV9RpHx
Zb2T3CmJfgVldJn5KkZJZbMxORyKIBzc09TjE6o+cLppOQJPAi3EoCRNiThhUaXbkMkjVHPU7GPC
lIUvnf2WphysRlcZlEpXsMV25gle1gr0cfbcRAJLKy7y1mjTEJZpTBkQjekmJab8CWMcdLg5+Eeh
ukG6iUDXmNbbByIIU0jFNUqNy5iS7ki2yGMWSrJsL16/C/0Ow0bWV2Cy2DLnZ01rua2j6P2eyUPG
B/y2PkuVB/PDk58cjGH65+6Ia6gne7F/zB7PbJNor6FNjM9Ix5CslPcpUpaacFz32k3wPjSSvMSb
FUZuu39NxoakCyRGzndeCkj7tiMr/hRIgkdeeryyFjZhzl1cgnFkk6OUUEkoPLkXmgb6T/gJp7uo
wL0yO2rSAgbQUyZuDBORXAr8Pm5HtHBVBwXBSqQssbvfak4wDsftmSF5TRb/Df90+1pocDM6AASP
KaOlSh867E+E7+x5Z9Zis7X8/UXBUOxlXS/V4xp2QRQk2BlNIrdnttGnkYAJA8+/k2K/gDHEgSMi
BHTlpoTtTF63v7A9dYUM7G8I52FKb5yeAtM8kAZATJQCfEIJ5s/hLdgSftDIJfbnKoriu9rO1Wlh
rvyzvsA7BNWG7UM1rhMx5kZZOqxY7Zjc8Q+653E2IdAk6x6u4RlyF7wBTU6t/e7zLQ7i5nFb+mcR
biomwSlL/MMoTZ/U6iUhImBoYPxL/XSXvG0UUU51HZYlyX2gjwF7TUe3YNrabMmdl8KCfVhoI+nL
HM7lMOrNyUgTK1CLyLRvTUSPCHaP9CMi43GjfZq7Q4T9gxbdADWVh70Wb0jO6Evzvjnuredhewjb
xPBYUFTMslbyCBAynlx8Di4v6X5yqSMcuWpcOEamtj12/4KlcPbsOhFgC3r0bx/uOrtBz9svjiRE
V9zCYtlxMUPziYCCA97JvuBMA7OqQt5VWO/ua4yvc1GN2X5l66didArKaXEsvDz8spOJsqMsTPtk
1+P1NWDjWZn88Rt5sauET6+0APY3Sh+OHBmf+/WNodVXRZod1VkmwDlrcJeq04VltSW3XZeW0BnS
VL6/hrJRbK52oaDNxyRwvFK8IPT7O7WvjHUMH9nedmhtKP/ekYa2dbazOAF+lN7Gci4WnynBSLkY
amVG3K5wVa/EN87MbcJ8Cyq+NgpG8nIcpUSRMI67bpPHtALm45WRTbDzaWO+Fr6xtkITUWD7zy2U
9OmY58VpK3k4sx556BpVUqQxZBTdppc9n0XGakimUF0G2cNjvr7ctmCybs+Do1+Q5CUs0Vu+jLCq
XP1NMFHFG3Ir4StMbVT3lPpIa9Ef/52yYx9yDjqxsvl70LPyv8qj5mAU6clIeD0qFdVfNJDtNjUs
xsNlyrexpyy0PQatlPJGWSSEiieP3FOiasdpxuOHrUXhmM0vomBqMjVMAGBLOZs9aAAcV29vY0oS
Bgw4JM4JNHrznKoPXZ+Fi/PAYr6Rgql0DcFgeAt1Wci8O6UZVxLlqWegWIUUn5T0QXoukUcu0t8r
2kNh1Dh1mwKmsGAguCIbu9khWzz+4LdFubchwHetJarPJ3PKKTaXAo9go+v7BwcEBIuRx/OSIsbr
ZaajtfUbB/2FaPeM/3FLcStwrU4LQ/VxeHGJt2iLvue8c5aExFw1PON4h83Wu5eQi1noijHVaOMd
qZGfRSeTNADlbIYf/CG5dZvtmRcI6lXiDbtu3ov6EKTK20mC4OaqtM32+Yiy/vYn1cUC/TPIKiPU
J0CMzhJ+pxZCdvn7D9+TtM04rSVT8eYw2HUlUwGqvbxc7rlIuhum+eWSuDD6DsU2JYdxz9qMX/W7
zqkYjY/FU8spIQxEC0V+Mp0xYcsfRgWAX0J6j+LCZzoyWvlNlOe3YQZd/K13QQvVJKvb2ZDQj90n
AwmyGoPBFzsOmvTSzxNNA8AuIlzjiAOUTyn18c1U5Aqvhpdz5cVIHATnI3tzeQD3y9PLG0ixogpQ
nruo9gSIWQOfAhHIAEKOoa/TIkD4c+UlFcemMIxDuRsetiCBPNLz9k1vrQSJEzhhL+dSb3ec2j4G
BYGkedRq3njplwbMlLX4xmVeT4gSscXuEjzmy73jRttbN9WLIe/VB9WEJmcNiVamD5wp/Jj2fx47
BYH5+bzYC/p3sKEp4XO9ppqDisAUw0h5sz7gX+w0sYeSG1XSem6X1mGq54fwWpzruTSR7RP5UI/b
0wOybcJM4R0PNihLYBV1ZZW6yrb9iQj/ZTydDiHX0DMVtUCiyTA7plWYCWJTQqS/0YFvPa8vAC9k
bTAktsIOrTqwBKWqqFdEyXurUGnxGNzIYOy5p9TQQevcedufG5EleY4q6JKkq0TCTrEanrrQaYQY
rqatEBYZbPrdgcv5nJQfPxTCSkcC2w4zqC5ekBxyXVtzLyK0xETj0Qa9oGrMG64LhYb+3j5QfaDH
7EmK6/ySs3Ght6ciVNXLVY6aPDO+SPt4gOdDQtz8fTHzhoOu9GCqT4Afav7LFIZfjN2+L5lIIomf
LH989TAoTsYfKUqILHwBY7J2n1bCB8obBW+FVe4IgcgO3TU+t8H07hFe0zgkSz8rM4hl92b0xFZ5
E/q3L0eMq7rAHIjHI/MCrPZzo+TI2NUDu3sfz+cxu4mh5kWKwPCEpyjG2yBlNODcfpM4UIEWbrnU
thxZl/oa597WO3z/YaQasrIae3IRxg16bcDXw2eDXMGaoYkMdg/R6T25MSWeZUqYxzsRMH8S77Po
8LpBJLC9durvwEnebT0G4cZ6J80pXVitT0oY6l0Gow5iRXsghKcJipHAL3SvI4ZKG4rWED9mD+ly
lP90GzHy6UV6LOFxdvJT3BVmaByBcZI7AQvqDWMNp7WQA5OQqYJDhsXgqIJ3e4hHFHVuiKdJ8c42
i8c5b2xECitRmP3HkX+9uLTIxJuXy5kqwukX8I6Jk+mO/syipL5GyAlHUmaBaZuMr0SYXIg9tVTc
q39vZTMY7IsNEUXRoVJpKESvLNRnFwxD5soTs3IV537UeJXcYEzaopiUaLlV6vBTqRAq3q5rJ8um
wO6JPPDSWjLivirCZFDrxcSwbTIPkWL2BQcS/FUsOZQMJ2AlY7GA56f3xdGiS4Ft2Zjmv3zhP+Tz
dR5VppRxyjrO+wE84q+9cAoerrgm2o6+437GNN4hTwBsNd8rkmsc0IOVcSYiYUSbvM+p+RnZz10i
tgt69jv7T7q+3BloMIaFImi52uE5dg6n/W1tutBxhsXQYYcLW+7DBeNaBib+MxxCeekERg7MGjE8
n/0RnceLIx3dKlB40e1pDRCtDA0d3BVIhNDpBgjW5s2KRwnMhHPQZJjAnc5y0tJK1xH69Zc4blcD
FuLcgSSjZ8bTu6s1nA8ur+fjYLMeHZP39OKvdCjPiW7Ddyb521YzwHHELJPjdGCxjZ7ERrhPeF3X
4f16seqXMWliqUCjaKxskxROlT+nlUYms2Qau5ovCO3fo47+BZMkdCHCzZLJhijxynv4/6o9qSoO
Gajz114sx2Mk4I33jzw1ELcdVV7lbTq6urs78C6TtRs0HE97ppxClVyMba8cYAZ/cfqOLZHVb1sB
HFY+CN7RE+cKB+K0ZzDOaNjiZze4nXUE1QwtOVGCo1rNUA2SPGmJ4i1Zp3mQZyiOWNIhd8g8APTr
zaanbJaSCjAGEELrSrUzObRCBVbzWao0bn3SZnTSv8hXeRPeJqIXXS7KZ1s3CGG85AqzZ9mMA2sh
5l6NrTtQl9yWXOIrSZg82TYIKAZIe6/3VSh0rBrkYXsBW8lJmveFHv5APhcArrWG5beSCc8PrM+/
SrBQ8ms5By1UJymQg+YVayRBtSrBFJiuDBosruHFJDl78eSAVbw6Pcx/FNLTTagPggvbfY2byjiG
jnEPV7Sw7wGp9e3gY+0w5UUIa1oan+QEoauBe9S3jPHa+El9cDCX6AV9Y3usdDBEZrcYYR/6l4E5
fgMC+aKOmwuhjpvoIBPOpdwhuWsGmMIlb1RkspNnfTuN2Nqgs6KIXBkyjgfZ9gD7Ka8vROWBm1/7
baZcPcE79JvMt6RTulzVwleYUz+TZ0gLpGMQgi1gZ/5ZkJftBNQj6Ou+qA7ikVBX6clpQCvd8/iV
PnZTFwfnWVApY72rTm80Njixhu6aNYXpcojobPSw50ahDAARpAYUrg+MSc1oRAQ4p6jb/GoqbU34
Rok97JottIPZzyg4Se8EWtdcYWCufJ6QAg/ltu5V4dbOy/2rGAXGuW0D0GeXqsEBATUTpzcrUavs
OSMQZ8vkJZ3wykcy6J7Xkj/Di1aJsZIJ6pSAu2u2eTH3AFB/pNcpG7LE0J/JzPGaa+3iK7ckbWDB
bc05VRwVWaEj0rUVhH3KbzoTb48kmM9mA43sQ03xUVkSN2Cdfv1JtiTLf8ufaM5v+yH/Q5b6meCI
vDRPsRcQhzwK6Dm26oQc0NfP3KN0xHRZQWZ4ihm3/oO7eE4y9PGBzqOT04W6RYDLC+FgUXjvE9j1
qQ==
`protect end_protected
