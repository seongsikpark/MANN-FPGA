`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
BOb04KJRoJudBEfc67qBMx8FwmTzerWgH+0+uj4+2TC+LGlzLcQRUB0OXt7HbNZ2n4IUxox2e6jq
ucRLREBvNg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
lH0gRqNvaFU1Qe0mme5jG2jtlvHn6qO4YSynPKrvVlR9oq4NdF1HapDzWTPaC+4q5CIpkGDp9CM1
HHNxNi2QTxqO4QuK6GOtgbVHEiYkuqfnd+cTvrfZOQigvUD/qqL4+rzteP+3gjv6AlmUjPQCBpjt
F+ZXXtA44cq7Wff9sgE=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
B5e8yQ/VR5u3iQcjQZqSUpATM18U2VkWBwbq7LdjY4b3/OzvG3xZcbckB2JS1rW1vweOxNbEaCPY
/Jizoi4EmRy1UyiGAZm2AdRSIwYTGrqS+BdnHvhdDLVMW6P5zah/3vCtv6BvIvNMk10rOTAPe8zB
BsXnzSnqvM3+ibDibNW6wyeDDYu53k9/jWCT2J1P7zk5B7517VkxLySq2BK31ccfA6Ac1yZglQFx
RXWpcxHS3We+LkV3c1i9zOrWwXQj7xZr2KGIBYwu03dXG5iUPr8PioYW1f8hHL7wHIZgqtI/IHZn
qv9my9/bGlR80tl/wbqa/3huS/nR9s4EqisgZA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ao/M3SPLH1bCKHknOdawe9XRFnMpNLWuIi5eGNbohGBxefMLSC1YnCgv3r/UqBqbOUTHi6qlZ0oN
zm10tq5HBMwJQYY99BEL9DBde0ZDFQ9i8rSmvWKBioJnj274Cl6O5LMcnBxfdZrJ5sCA6TvE8jC1
KH5ch5ogHkyyXH0i1Fg=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Z4xJBBQDsflv3TritnbaHiNUw8gbGWc44bYVBY2l4Q602T/JkeZY6h9rBijq+CRkyKxBOfnF7TOx
Kz3fUVVh8vmFixf0mO/lsLDjY6yAndkdro7d1XdlsYR0nYk40gBpto/KRxYYoiP0Ns1oqPDG1Xfy
L7PMmN77S2D6PtixwKs5nbWJR1IY9/kj/P+NqJ29uAgMOofsgEwRmJne1g0dTTi6fYSlxfwXpWpF
SruF0Fy1f8mmNWyi6m32HosjVmW/gUbljtMQOIBzIjoEMR0Mm4MYgrbjhotdc8d+zbOoQAjuE+b7
EsgEcTuSJlOh+vBbfOvctIZwhq1IIRqlnXLp7A==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JfOmnB7OrPsYkjrR2D4DpqJsTszKORckIVUffs8tEkV5t+uIBh2gbrFyPGCo3dq9R3U65vQ71EDE
AxBRVk8H0eUOiu1iwM9AALMz8Eyvg3LPW8YUG0cHC8hcp0jq0N2bGiLSK5OIhNx3KCOoDCXNFRss
v+bbip4xlA1u1CqcbnX4DjX7nkRu4IbdW1wko74lHhvA96qox7nNT05xFD7Izk9VAbLixY655gBQ
dX3Cj5lrzn/YmrtITOxzS+aP/bgCi3wgdsm9YMHzewos5vWCyqGX9tkGocRxBaXMiNGsIxa+Ruy7
N3zc6Lutjhag81i1aI+q7z0qca0LucLZxHIrJA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5392)
`protect data_block
SKPZOyLOb7zPzwQIaDX5TtkOpoo76AyhQEhuhq61dCeIPnCI9prTHt8/cyZQBf1F6QWr00PVfvkl
xz5te3qZbvfgcY6b32zeN+n+WEAezcyQ22B5FL1x1T3cm28aBuhCVlX/Es1/8lLe6sKQa+5Ii2r3
ju8nzylmEroFBeYR98WcezACZpewVeOixd+GytYZpsAXUcVRyMZJE/MrIcWgNUyb6HA4jIXfA5rA
kzJwFTXgYWjhcFS+rAPlK1tb6ZTKE7lASaK3FpvFGQpW9LjQWkNZfbCsvob9uQ9tTummZ/uP5pLf
t3jUf5LeyoooEMvFqxoZWnaG577MQatFEd/A827Q7V9okSkiMquWcSKkrifhQKHEdFOpJhhR70v3
iA/1b+nO/yBABdtaT15/k3ybZ7TxkvnUlrs3W8f8AkS8jmKD4QQGLalu7FsJq26vj5XFh5lUhzZg
a1KH0GTeHrTKAHBVGR519FQYl7AYKZYNJOoU61sUp1OIfWEwGmqRxxQkzUfdMSE20VhD6RgRsRJc
Lv0sUjigW6yhkf0M7s5NI/e/uvaOhz3pE5jIV2EgjMXBhvFksbTjjzacHyhg+oTUOniGxFQFQLcq
ShsQDsmYVtcsMWQSTkHyZFRaQ/Ah+mo0CxhYEA1yXeJ+FO4EG3/F6Qr8o3js9yOB8D0yWoQAZ9XY
vrdZU57RFcBznaEnn23VIU4Ft1+RbVlQ6Ff5Zt1C6wmZ1cooHk/SlhuJ7fxei0vhcYI46KcsQ6A1
ea+kIphO35mKUhd2Cis3WUQ/IVkq2yh6tXDWhmgyu/tJJJsK0kUhwpAoCq1tK9EChWqRHLaMMbro
1E9t5Vc3UcQpuoPFOppBw4WJtG0biyTshDEn7DAKvTGUV3PZHgROjSmokqfln0a/rg9xAZLHrWwf
DmD3vG9Z/StbWLGUKg5PKA/fkRmEwWjfWjWfR2YCtca4Xe2BzO7EMMSn4EAfAkdNLzW8mHlOUCnx
Dyik+RPvaQPeQkPvA+9W2GhxkJTOwQ68FDRtdTJPt4t/FASMkoSoXQUOAcYf7fLw3qwrIMHXKbT6
zcA7tafjWKaOV9KQ1MgKb/DzSg7eGaTKphHeSg95TOoYgeQ3yItop8S9fyO2ALorvbkZ+NHW3M1b
/gFQLp1YUwte5uFtNrrGMgxCFJ3SZ94xMzzaQAmsbAjG1LQPzA69mr0YqgzOZfPbGo7pEn8EY7h7
vzN+heFgr9HfxoTtFCd6iSgwBPDs1UHDhNp8l3XmZFx+we6rL/kghjHvwxjvbpLS19ZPqhYf+hf8
HjFg3TRVhf3rEMHJgUia1TJYuBM9NE/oIsJ4zJTEF99Od2gyv4A5hooEVRA6L5djSlRIE+m4uUPf
JigehTJiQN0HKOI22stb/poot0VA3mJQAfT/FOUDj/2y3gqUgPrVFL37aujP7uxKPeVEnZFiPE1E
X5Lk7hJbI94FPhHvameRTmq1TpshAR0VYNdiaaUJF6OmiTlIbakPZm6pN5Cs1U7Q6whxbqarbqsZ
JMpRi6gGg18TNWNp3JnGjB0Kst+JqD5ma0wKpBOH3LUEIYSDEK5zc4RhvjFdxeuGWP6XmcMuWQAj
K8H0SeKXS5uPPGcfIaVwBJXwI1bW8F0V0C1SpY/2heu8ZhYl4P9m5M0rBr4zlm/FJWfJSfwX7BP3
D4co1gwoCBUsmqEU8GqeHNRndzlEfA//eC6qYC76VBnkDWnqB1wAXz+biA3Y3uZ3KFX8Zl28ET33
bcYLydAMOyPGTJ5yHQ0AmVp7t5sslMADsagtZQkCmW07az1vsToNoIixiV/+ZP+2WPkV9kQ5rMf0
kS1EH+0ehX8hqsFVu5gorVZCT3GwljcKnyR2d+8y+LxzOVK49wDzwiDOyLjSyh/He1tMiLnxqzQx
kh1M/FMk8Pig6MPFRPTZKTj1rtbDmHknbWAxIrv7RQhSHzIL5yD7PEZUSRSPYmXRzm3DCQiFNcD/
/PqlQdZ48Jmjb8Mj9JacT+AYSD4Zw3kWnCZwvSZECI06mtiRgLqIvjYMxe9+gkhjmcqkJBracZBi
SzMhBnY5P4rU3XV5LcIPQiHkfkI0i/tuteU4K+3Z6CXz8Dv/0ylHso4XQvCILEY5coi8XAU0YpkP
xLZQudSsMQbtkBLiFti9g9w8C1bcQtm+dTmXeTYDBjkFXyA20ZwQTqzmXQz6eEXpStmNERqoHc8l
/zXp+c3a+6xovU0KV5B16DnXDSy6AzV1fgAXaWGaskzaaCjO4mVfMupqOFMRjYuHMadN7e34DU/4
4CP5eLQ1ZQbksSEXUaEDmIQUaMAnVOcDPouACGexN2tlr4a6H0EjgBauFvN+Ex0zjZKy0IgSYr8x
DXyLCHymIN7GPwxJSgY9QlkMPejniG6hrT21EzAUcZKQNSpyrIhinqYSy5mciTBL2v1qUh5d0Kiz
CFYkIP9GfwF0t2XN21x8tbHQLzOvatoezHwVAvUsf4MYn1HafV28yeML7oAnyD3k5MlOfZiK2y1b
4g45aHWt5+8CZ3CKj9HcTiHldxjQeqNgd2d1fLi6WqNANeYXEcRLSNvzAGS+ZwGLWN0TAXvZ571M
k74pDyVpo5erbYZkoUq9R9o2g3NK10VMrPuYJTUH0mZPrIpc66aHV+zTcgbcWiKc7BQTKcjHoKjc
4syq2DxShSxjyiu0Moi+wJPejx8SvA80howch2sb1seMAuPeOtv27qQDQPJsFTRuc4tTx/5/o6eX
qDbvpIKNMehAR6psPGltMylu1Ja/MY1IVbPmihWMtBqrYO6aOy3/+pkM7eLM6Rk/jeA9yHxa518a
M+LO2ySAiuvubSK/GU2JHz7u3PDxqZknU1qEzrEEjAKcT0V/FdQ+rpSV3e9nQ7trZqG6YzAqzADK
chY34/44JBZBw6QLOWzjoYqjHF0wqgsyjJyGEH1iwzqKp0yot01lOL6EbyrDvyTsPscH4oKITM4r
wMXirF7gYWpvhowqtdmgvyvFAVXZ8eu40MNeRbQCz6kePJXDrqm/ftndmdQeifyxCpxI/eDWgpV7
U1bAG+fAhMuMvl8Uia0UQ6aKo9qVTlLaQ9uglN6abjwrdJjgeakYxQ/foKXoUvfbHQSBU7oF4AjG
dlJz4V8ifyv1jhwGWfAFYYRVYFnkY+Q3Vv181lLCBE4oARjOmaBGGfVvDluk7mXKEPX1RYRQwY7U
2KMOOxV9PZv7U/xWRbr1SqNNpnnQOxInjmxGbh7QuYlw5MvkPssdHad+MZZ8z6bwaNEmUQgLtGge
6znyVTtF1gjATSUWs5N/acYCRL8et7mEoohHqmPsWm0bFLWrH3BlRj46nLZxB5qfEYLUWgrwlOlH
eZ45Sm8+gpynW7EZGTUmZ06VdpXh0/TRTv5tkUx/M4fkGL8mm2LyLJJU0uFpXDU+FQ/iOWuDKK7o
y/HS5+vzHE+hA5LfJEVm9duL0caf8zXjxsa3s6c6PfYJsWmPz9k4Z4HyzIiKyi5Bx/Jqr1whDXve
ax4QxpUJfKR4DXfUPkMLvUGkQcwuByMm+7UIrrybhgDPwWkWd8kinRSmrEOVIu6KD3ll1x0U7en9
1c83wlDKxgCqmvaHy4znZs0nVUqk8say6glw7fkTWM+skXZxh4zrHvHECM0ye8C3rxmZjCmPNQHX
iDVFKzIGBvcRp39+hQ2Pa3avaeHyHAjgB8/fI1dS1TSMEfSq/Vhv2+FMIFnUMKoZlqF+Nb+/e5Ab
3nPPyRV83QeDr0TAHhmvvTI1k/eG1iV8t/iNhqE/X4vjdSaSxqlsTEpFOCu6eZLYQUjewnq3JHBY
qMQHc38PUbfpV68G2+vzVIa6qHqFMvGdmAi2J9H1UaY6+bKqmSC43DY1mh+6ukQ2t6BCBU9ZwrOZ
hg3tHidntRXwMHqXzXHRCETfoAAZaeZibNyaLFEx1bfQZIj5fVUyybP7TnADho9zlkyPBM2OSHgZ
hCFJvd60j+6OpziNeG9VfZm7QIYfmEwzGF0DIc6NSCenIJ16hQgwYABjyygjZQStOIOG+DVOTcVj
JFRpO5FS9JjbZnP+Js+7ZGDACYPnnwpOJOEcBHGYhcBiTNpVBDZZG3yoGZJ+CJtGczS7MNeXloTL
swWBRFuyDbgAPtJSargYTvJ8e9FIt6tM8x8Wu2+605d4cb+F+5pOA/w8YVFT6aqNIWCmX0Q2xH8f
CLECrHi6yok3OY0Rgven5PYOKQtViuat/hmdkrOtZGMlCC0rg94ndAEqp9G9MOqPxILSdAIA/DVP
Slt2S9GHS0dlxdpqbXynqz/mfzrUqFN6C1smaRz0Rvkra6BA+/uQhNXb2qeH3vk5Hlm3GQFT8LjP
mjtZf9t8kdHUX4hmzq2xdGGEplyvTU2TMbzTiUMuqJP+v65huyFI9SYTrbcrLaTxXFX1EA92dq5H
unazuY6stpqrtyE4fXRVX3XejYUwHwtMLdPce1TYHKdt99fIChcOt72px9G524sZFJ5o8dF2sSMg
FLzYbqTR/9UEQBlGHjzYIQb25SAq3PQyYUfuS2RiAkJzXQZo2dANDCXraNmtwekXRSj7Bh05dEK+
vkdrN32mEd81R6Yw6DFWjH6/4kbTAsz6xSNMkNqFwmd5s94622CrZotk7CFR6MMbIQBgwMPQ1lOF
kF0FDG/LxotNu0iQMq1qqXY5XlgPat8McDJvmow0PGnj2oroPCqtE2ZEYKlFYcspdnyvfAUReLld
sdMZmbn+8Bg/RdfZlgDUuwA2cBshdMMgzIuqiHXVjNdObPx3+4dxxoFCju4FR1ERm5TH0tdPqtDt
bTF9zw00e1HJO4EdNJYdZ5Wg+bjaRw9u3NbnBA+2zB398WIFG2rFFYz1G+8TlCSVgVBmSCRzrtIw
Pfn48aBTLD8OosNfdb8Fc26ZTfTwZ74PL63c0dRjLFJQgulAPi8XrGu1zfwlOffSRhbd9ZmjlHHY
ypCoVCD96yvEXmhHdkuQ1+GBA72u40TMsvKg8U27RxPhvr3STlJOHiVltesXofFn+O0IrE/+MMbR
yQx9YBlXzYOjk0F4FzR2n0eG16gzD6TslcZatcV+wr/Svr9+Gwq1AEer2zSbfpQhGyK0tKA7e6TW
gzSYRJ46dR+aXmCsp2IPrVlpWY5SjOOZXF/Qdm+0om6x3mZdUW38JNfZjUcDjwrKidqU+bIkYatz
sEPPJ5/yegCpCYpYgHltjsTJRPRcD62pK4hEVFIYNHtrVlI7ge8Z4g4WQ5kjBbt3xzBaZWvP977+
L7OEUs6N2t5o0xVK6WScqKGq8FRF3nY8TJEgXGQkeP2ZIKKihrUItv3Xx9FdK8BNOOFlK2WqONpE
szjMarQeZEwvfYKBYiFi3c648hGJZOnmjxzXLMjkDuwayAps1q7HWycBP2VAcu5TXIrUyP2RXSOv
d+RUr/R/rq6f2dZ6eW5BFLAayALyqjX1dYWeOgc+83u8d8ehY2FVkHm4FbrkazC/K57SP1cBCf9J
StuBJe8hYLZkeCIWveD/oBiLbC1csMuEUGbSu97KoJjHnJI8+LZeDzNiXttG7MQWobSon8YXPNqN
5+Wzph1/h3TMPIKIe70E5p64fWOE+/mu9pesrfXdTUC2Xqll5s+TUe1lAKo4A4rZLqADxj6E2kvE
fgkPUF/blgZUU5kv+aWMMybOnQ7UHcSGu5gtClyEz5cxduKRGI2BW1OuSfhAcPv/QkB7gBkd3tWl
SJbB0B0AW923AfMGfvm9c8anuS5ZvWA9dGz3A7ZvewVx8bF031VarqKDTPEjTGWabbdw+EPSdfMP
QV8BUSbTQTNvjHGtfY5m60Vz8hWu8S8IdgeJTxqaTG+FoEvI9ZM26cGnb2yal6b5KYRp+APkUDYP
yXrY16KMyqGj1YksN5IjaHPumrChDJrEOUNUqe5qb4AB+bnov3xd0pLoocqB/D/Jq46HqQ38XgKN
5/iay8p69aETBQiJg8g0LEAmUW5qyVo42euz8y/7AqpETjX4HTu1i3So+nVra1LMF07dUEsGax+k
o7zONQ41yZdLDS+WCD+SbbN9HR4BavMo1+h+krEWPzrz26LSu6uPcyzrrg1o0yCOC+f+O8XYTqHQ
vT5D9NbBkETR+BI8kLF9d/QuSs+JB9mzisx83B00tR7gNqO90tdNPk/Uo3K+86kQ/UZRXnTXwDV7
axIHYXxeqc+4Qe32mn9yomlZj4cK3FTkiljuFO2xrwLWtqhuR7seL0l/Tvv6YPFUUQxjJldw/HMD
HEg4lvOuQEXe/BjKtY0B6EGt8oyPG0nrvSKDIiX0rMX+9pkMLZe2mSDOhb6fK1De/VWNogL6GqOn
fSLiTRpr8PC6+G6ZCaYisAP2Mk8XRZYO40SBFLYfEcWcOT7zZrLTB4JDz+fWG4ZYKvuKFh8n+OFR
tctNmiu0FMKkdWCO/nrcdtZG6lzbPbo8/CI/XasSSECMrRbZBFF1NiR4aVaGFxDTBf3AB1kU0brx
1HSSuvqwpQsI0OgBgzhx5yrO/xQ5ezRG2D+PGDibCvWNqbqgntImA5AfBGON1Mt6KHtVCY28nEAf
X+91s6K53k6KEiE+jvms+0D2W/LVWjcxB0gjeTDewDaTOCrnVKLqNO9+ZEbSwjwBnfrUepg+9jN7
YTZ7J93LcX7W9UbztRTorF3RiW3Vi08i6TNcoNJtIoMiJrlwZAPWkG+l+9MFWIonp/3VW06rpsbq
l6jox9UmT0zYNkJo/jnXTKyDlLQ6r6MCYYq373NEfOPwZ7GQWQ91/0CUoEl+KA1xIvqO1cJ17fvY
fevCWoQmt68+mWl7outJPPef/YYaBXBvDNldhqX4L7xGTLjAhfu54Xg/94ZjXJIQi+3/NqJhxzP5
ulcJQV/0t7cSW54mSjRpRqNHNMjAqusG1KMNGZPTuOc07krYOP30iuCsTMOerG6LXcyTbB6mqgKI
fDZPTiglhyo6/klm8rYMYyASZwBcYDq8xjU4Ij5inK6YbgxCnGF1uqfyht5e46wRFNxlAC6Q3k/M
EIE3+ql1m3XZh6X+mWNy922GIiGCwz4ju0JSeUNF9DJ0rhn9ky3ZlqYGbokKdptsjWlgola4HD/B
JQBfkkQJu/2sNbXnJa/udYihVJgJ22OiCQX2A6cwhJ/RGc+Rbl3irKR7hpfU1cYQzno8vwofDNq+
mTsBR1W/OING2jBw3+B4y18cmAeffiF7uTV/CnV6Gi9bcQ==
`protect end_protected
