`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
B9ZpeWvBQQjY4dr8OyQgCWD6kSA8+HY9SzJj88aCfo3JohYFlKYJblw60SIQaUnjOxXx8h6ELYIM
UjD1sVmQ8A==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
iwVbhZc2P9arGEbPkPDN2Ciczyqo1Bl+qfZPC8pPG4eteDJDMYhL4//JIPliW3+60AO7KZbyirpX
isgEMka3z8ObvLYO298sjCHDgs/FZfmZsyGmSoPOb9HHtHVciE4p3TjlqyIpvkIcyPdJ4/fD49Sc
nvJ9MvdAGyLQu3dwTZE=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
oMpLZGheLmkvkHecy891anqU/IxrSwqdYJi/BCqFCgNsgmImYYfizgd6jy5pHiJ60XGOPHkcnOTy
jxaGYxBI7Juc/kfJgViQFVV1aRuuXnLsEn9jAYeCNbXGjMOcxwPk3F6E5P+SRFJdfx0KMPcD/wM6
bmyeQUTBbAdhZX227QTipqzrOxkS0QaVhzCDUr2q4VKPQsqZcTtsxxafdT3X1+kJkg+J8PgudGXM
7bL6m5q4mAXKVyd0GJhD7Qi8vPhpRKok6azS8kpVpinGEW2jOl+g30xnHo34r1Y57zE7Hac3U3mE
kGglks8mYGbOgllRBqR8MUiayaf9z70qRFoHFA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
e+nYdllhcdKHJg0r1my/ydh7lhRKOoftD3bwWM6aLfXtcw02WfQ5kb3g9y9QOMp7sTQr6BHcJLPt
ngjNHJ9dYgrGajeUJ2ATpRvbTfhC0dOu8XDWytje16mCpWOwZ/hGr04rwbOHpcTXOPGdOE/VrnEe
X5hIFArmQ6cPSEF5nr0=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
zSjmKksidjShQsfA76nBwQ0teiFzoZZWQ+NicoSnGqsbWtnh1xC5oIQygAEkiJ7KViOh9n3kKUHn
T/7xc9+VdDMh4m77ilRe5mmwu0QDyeCK3aCjSZoU/zujjnRNCwncEiNjU+Gv2xu2Skb7GZ2pLHN/
r3bxm8sfL9KDPLKc9jA+Vo4EyJ2KkfE+MdKkuK/XVdTgh9PRlhFmAMvYUBNhWNbe+GfbAcQqFErh
Wo/ACLuJCjJUcZa4Z+vmEqQtU8uNZWUzI9IHtywU7ECvMX0j/BlC1BtXYBIYzozfRRe1iYXGiZkh
rHs7xrnQ611g57bj/SBA7p8lNIET4VbFnbxVig==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Oksyn1Lpp8o9+Nend2BRJah5VMeR8XjajkNcetZzZabaL63UOeUOV3m8kWRFtG+ALxcCfCl1m3XZ
RL/RbQaq5UobujWx5eieDvAIYrWHCxmWjy1EjcD7YuPi3VynYio+STtqql+Igru+3NjtjAZATsml
313AMJlgO8hvLTBcs3+r1Qx7i+2ulipkTg7bCX1sFywvBbYGmc+T/j6RXFVM0SaznzSl0PQYxxAz
yjjhfqBNDlAfLgRFjyyKSpGR9PWx3mC7aXsYJrTwQUQmd1jlXVRh8zCaqpZhaRQNbIlT6/ISEfAx
hJHHib4bco0Yfo3fQ+I+EtzPmOJztekW5j0x/w==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 16112)
`protect data_block
ceU+yUO4VzpxiJsMsHIFnSQic43DyzM95ScLRSFtqgaVOwkaPKz0m/sbvEZQYy6xJexkoMLnOC9o
/c7srIMGWMynBAosW81wKS+cRKlmDnwYox3LU1hWfFDRsWvOvdDruBDMIVbhen9Rq6qSTmfM0VwT
5Fko19gTNooC7o1YhqrsdqNMZvueZcOUb26Wq8UFJCpxU1EZEu+fvXrKcaXdF0wqcOj9WVXVtkDg
gnTvWKL0DhEVBGD6BZ6EsA4dJ0YLZV9MhNtEwevTXLHVLTxXtp3gR+872ulabEThKWmBKwjV+fb3
S14IGG8G/LBLCDvUYbuB6Na8fQlx6huG4MwLxegs8etRZofNOIlw+VEoYjdZ3Ov3BIfne0Szo36H
yozt1FZ+v0Oa/3vUEgA/qRd6LayW38gDRleIKN/zps7GSXoXs8u1aRGO71YlDtPsgVrMY9Szryss
+SJNwYr64+XQ6gE3S0oessIBc/05E4bGilrFwAOk1e4xZ1fd82kgFZO8eysBYO0cDVLAhbdj4XmE
Piq2t3r12GSevytWRxrSbPACGBd7IEYzp8L9mxNMSTSXgMdn7/0vON6OTxn3r3xbPP0OB91bRB2d
g2a9WkvFHEvxZIX3KCyN30O4DO3Axx6iE+OaqJF4R5Gvgw7QtYnTZrlTaNxkfNY4cKpQ9T+0aCnL
0hD0IVs6BJJlp8XlvUmQqBfteBRexK9cGRLXxjGBZNd7mR0lSXEdxHuefbQMNys6X6vmE2xo7eyI
mpxut3q44ZxeeF30kT8hSLSgKjObwc76zlZVo8wMGhQQWObr6iylsm6jYqRRMZta02vtAQ7f1KG7
OqifJFJlbwyygrDKTsVN4zdq7OFD0vDpFhwZZcma+OZeFkA2IVA+ZQiLydnLbAOxR6kZA1EGdhhb
Vpkqu+1AqwDbtWKjsYAbjDaYTgs4qmElZk3morNmHIhC+yGdTdh9MzTAUB6Tloax2R02Y0/i/IS9
ys1FN0FZuvv/WvElQMDgoWK4BkBkt8WN8ORsZs29trfv64gAi/dp8rQsJ2E5c8OJssz94jq1rvg5
DT6Yww7RBpmg28Gj2f6GxWCPwKpETrQ7+244Djk5NuBLXOVa3KdmD5yYeE0fW8BtXZAWSNHhOlGK
FYMnwTRJCi17PlcMJkohFqLJIxKLkTe/dHjdvT5+1r5BPQgsIv74WISew6eZV/6U5LCl8xT4fUNN
ybsvdr6WlXYxUz/0SWzieGSFdWA7HhUx3sIRLndgggyK+gx2IAHzNA1Hr/GBGzn7TnPK3PY84J37
A+pBaqv/IlQLQisg/eND3jxJ/VgRBNiP/Kn0HUETuxKlavFp15PUlfKYjfrvlvJSwZzqc7lql8hp
wMfuhU1okBo08D6yC/l9sVKD0+FbrgIs0it1h3JMjSBMoH4/wr235mKxVnVlTxSUl6jIwpuw/E0X
KJYIc1toNI39gTZ0LSuFkqftYNnXUxGsAd68kRxqeM7tDeBflvRJLz8rjUurYThR3To7gOr6XJUp
KzMWOhOyRNJFD0TvONnxIuE/hiBoFViMT+VMi32pOSrTO/eZoPQeSu56YGKGUkRaBxJFaLQzU/Yf
E0xlesWrvZuhDuSpYT4uMyA80iJUTMAI7D1qlBs3W9LNYFYv76L//5rX7pkX+SMqfcB4fuoLtZUs
uJRojv4+MTRJ7rB/4uwXDGVeJdN0PZzSItpTpAsQaUfstwZf2ykfzH5IE+ldvcKaA66tn5jqFWqT
AJR//RY69jIxa5gCMuobLeKjWq4ro7ZTXN8kcXLi0KoDU2XVmMF7KB7nxUkbGlxJSduo4uGwP9k0
i8urXD5tGiJ7Uk72MmNa+qXyGKxZU1AJ6hikYOukAn5lLitEzoZYIyi6Fpphm2MKHx65TyiHCdrc
Qk9GLKyX1vXGwpoY8eNqg8zGclyJkG1YWUaWDpHxp0SzmyUdCoXlIQRmnMFgbejnD0yvv1z4rGIt
f0r2q7NjsoALJMEjyOWSFqgNPS0L9m95yXSIrC/BMYqDC/Dc2KUhQncC91qw1nbqfqarvld71894
ByPV9UDiRLNoeWVV4/Jytrl1gkWOJ/r2bl7V0T8arws6udGX/BAKbCXaTKp1u9jAZFgcwInEON0G
/1SK+5KhwExrkBDgRYLVDNPEihnRGZIOf+mQi1IXNQUhCcOKm4dQoD/IxP9OnFe7n5cDuqbxBsbM
K8QV27ESIQ9N+gU9BJjrB3buLbZn0Cb9uZvH9vCYH3goGy8/MicOYeK+PFFwOMSxr5WuPWtIpYdn
zhBS/rMIuEIQspEf3YV7tBmafTt+pm0T1bVeNlpioGy7MoHfy0zPBt6JWn96NsIoXpGOWdwSdJpG
zbZ3/PRX1eWoy2WW8mRSDmzGgciJyml9nnjgJ+Tj9x/VjmCGElTVsBX9d/7sAktCHODxfMHhHS58
3Dk/IMaTePcmYwwjbYSZ0pfi84VtDDOyFIGemtPKSi1AP0/TkMu7W3WiFFG7mqll+Fzg2+A/jNWF
p2k5XazRdwJ/dDD5q4r4ZrV1DVaJyU05N3Dxr67QruVJIbUPQlrSADQeyQaozlcQ/CHDfc086v/W
FanIH9DRZrOJOPWoWAv4uZYehLGBMMP+G8YIGwhcEhPXUdWGgQ+4QtrEuBQ3T9wwsO7dExD3vUIl
LxIKfkXVg+j3TXqkD6xh1yHzPmrrfy7eJTMGZiQGWcNW8+76QUorV48DVADOeOay+UWcIefy/DZL
7su9010rCEBhnfuqk4zSHvyUdQzGRZMrtxT/tGRNaD2Em9yyf1d7dHOikxpnbv6RRRiCBPggm8nf
oFb8SKTcR3e44z7PtAVLGjna+utL5oZ96+5rW4t0GA/q7P3+4xUGJqQGjxf1l8Oi3reaP4LG65G5
6nDRdkun+w/K4HIH+SXkSSfleaRT61X8uhbJzstsuvmiuemZmcJ9Q2aNMdp7pasptHCS/Og4zyJw
fcPOp/c3AsmVmrwN3ikHSjPpbv4FrXMhblUfSrrw/QNwcDtDSp0V0z2xg6f8DZa92XyEhA8iiI+d
XILQaEkKJwziVTEi2ZaMyOPK92SjEwIwmQ+baN2rb0hS1lHkISZGZ5yoDn4Qs0gpdm4CRL487lkz
oxvdwNbyJ6pSCbM1cFPQipZNmHq5HG1zTscfsDbZ1g2JmMQjHOOq4h3m2Pj7Ls2yVIM0KVjXiSSb
ZvBU8jQ+UH5OrlObgyXHd/rynBGlfohsGYKYtBeLOJpn/Z/lSxFyjMX+D2QRwr1kulrUaLojpcsi
bpJyPCigweprtnID4SLVj7kneYEHGSXD3qwvrmsz5PC3Q7jWR1DiO0fHRtIrGBlInPrnSqXUKXqh
PGtjg+0gBiAOUJmDIFBayeW0OkJSOf9SDkZwHv6f88LFhEDQhmnR1b2lm6HFvAda+UBCx2Dw/C0F
c+a4q5/9jUolyudONWTyMCbm7Qh++SLTZrZoZ+bnjrDld/e59HTUf5VAZ1jKgPjPThEpVxdQYjzt
Xs2sv3auDTLUmXmKRN1ESnoicu6o83kkJPwicKwk+Oid7+vDlTNsIhG12syzHj9FzPmlKhayh7TO
wQ2jcF2YykAmuSrl9pjW8VUNJIA+h72D5IgeReh706jm/FbOP0dexfBWyzZCVb1A8fd0JktMmAiX
gYR4nVaP1AzF5qvi1D4q4HuEzUOyhj3Y93bM7IT4I13N1vCGFdk2bS/hR1RT9gLSEnq/8Az6OxUh
IthpvpwQWkVcpAS5r2YK9frtoWnwvoSSYzvxE5gPg6T0yU3EWMPtIRas4CovjYlf6H0KifAX9IUZ
eIgxq7Xwx7k0pR3dnqfoOMMXK8Y5k2q6nSo1ub4fGbXAMe0ZYh+tHsjEdgIkZgW+5cVEbdiSOKe5
9TCt79WXzo7aj8d9iJqsGomehQdBuMMZc6KCdHKYqrjMxoD74rrVNHBOzaBhfT/Gk92/2sCFOOYk
mEQ7vG0x6zXW2Malohqzrh7tIGoqTYhcocp/kFT9rDrrJDvRtjxd0gvVDKBhr76i9hSakHL2sDzY
1yjyPN4SVpq5fNCvdxgK9BWF0psy8XvQpuPjKC8gXWVFy5I8jjz1NWbuTr51UaBN5DD91cFiqKLz
UWMmYBk7KoodxaB+1D61Z5IuJm42Zvk3nT/4OruyfjCMefjEXblzVqwXDHHyUjpmnNtO/cPdch6Q
LZB98v7bK+nh109uCwKbTEjFiE/Ej+QXF0TGu1UdyQmaTzWUHXVKrHLna2M+EjofYx7At2iOZ+k3
rzaLCcoKeJP02gT1hNESo1auvfXPG/xLEMMJ5VwY3zhyB2v4QGlyVqUOVkeKx40UjrD5gO7z6Slu
fL5rrd0AbU2GxQIxkWBG9pNP5v0/NFwboMrR7xDGFx8JfJNaeEEIxgC1gLjOcNcrpS4Sxd/hqiW3
xHWne+Si4NmCDVlA0nWtg7lPjE5gI8cSpny3buVNgwLMSV2bpELb0ok6q61YI4ejSYlUUqYfLIfd
NY9xucGgozdo7l2zQ+eKdxGeVFCPLSpwk4DGWfkRQXGCuqmR/W39Pm2vW4vw64PT9KBTF6tCqask
nG6QAsqCnhGSkOhiDdmMUReSkjGORdO51gA0Lm+EidKSCd1LPGwdkMuq4DwU3e+6SQmcB0cKOzv8
UvM9fDbgUV04O/8v6DSkEIh4a1JO/hLU6AGMcIrOsL2+5iCcz1BpR2ShFm/mcxzlTMZ7iNYCi+i/
nfuDjiHb8AivVCCEGmtloVPbCpqfG+lVBhrruIjsQjIbji3ExVrXZAukPiNuso8ckIjW40fHhb3f
ws9S30Qkk7gTQSw8SAXosSIOKinVJYOPUWyLhDZRr+XdZ4vkgJZ2cGgrduiNmPdlKgv85cHBavbc
MGH6kwY+TuRqu0KD99iKVx3Rovl2txLOevzn4gwYVVnPeg4ChK0HGuJVi9Tk15wXOp1ly31ECPW0
ezjAc8qK8J8+SlKXdnkRwTNyyXLMRxTeeH0pucKT0HGKSXl0IdV/6YU3q8VjQP0Aa9qgsE4L5dqG
xl4p06ur0Z19eJ1gyqk3JEiR29LW4nR1x0WBkekfCfdW4VvxBRfVEtlmMMt9NYOFrE9LnwYAThNR
QNK2PsWZHIUbjeV27JkLKzyaYJha/RlHe5Z9OXhcJzogIg1b/dS69zeClRFD9BFt47ZlZtLjNIpJ
RA6WZO/Lm7c66U+9sVH1pENYUpXng9W/tzXX6Yg5HZXICuKVczH08gOYLcf+Uaymz1E1pft082br
LtBwarc+d2FPyr2oT8TW4pm2SdvwF2PXRi0IFikltWTiOPP9V8+PUdsEOMy34+B0zRg2ndlg+iyf
hXUstKwzDiishyKPG+K/WIjBydaQW3P05TV7iL0lk2tgwo7ACBgazuBWMaObAWM5JkJ+6CI5QQTC
hcSaVhKggZxERnghCfOZIgPJdt6t2ierxnMtclLutkld134g/hjf9xEEtzuUlGOR3TocbSWd+NmO
XKf+aKIeMU3LuWSYygeQmK7sFL4lzpZJt6u6DTP5pL1T7ZB47wkAhAE7gPo+FuNPbwxgnvvQ961B
9Xyp9aSaiPO+4eWd7RCE8nbDaeAwypit6IRiEcidYSp6K3JSh0FW5oZNc0OnpddaafHYPKbndbFN
0P0pE0lc5AHqHf5x4qxp8FUp4surYUIl1wVWihgErn67mX3KWSCuazkLcu/+7Du6MJCb5hfwnKhQ
WlnK8bQ0qPfEKg9E6TYpTMPUILXETWW7lJvQ7BpfZVywX6IiofxWluZFUKqL3QMiAw1dWLXciD+P
Ur8+sPKbDikZrN60tqFha4JX2VP51aQZx3h7FI5ENkX0bUx5NhDMlQxYT3q6PwNI3AeRuafz0UoG
NOL52Zb6yGKiTKJQuk6LE6ybTSxSeEpWy2hqRIlSrFJoPRJpyiXYyVlp0GxXvmXMW3/uk7TZLi17
OUIx8hLrlje+AIEGuit9HXQmSUk9XWXXZHJ2gBgLPeQnx9dtxVbiIP7gTpSJSK47CtkTkyHBTE6+
BW4o8+M6UgWK0nBaUszC9UD5gnJ2eIkjdfJLx6Cb7p+XyWFvTU1eRBVCBxTSw+UIGiGqAoOVlhmQ
OnMl/qNQ4ijN7HuHi31HICMDSsjUvz5e1NZEJBPfHTAPfbgu+vkDNGMVOnSfKssON8/ors6CYbEV
lpPIiw/0F/bJiNixqGFbXZdmYQ2Rt5w+/591dYeOMFs9eYbPkB7+S8HmPpQyflgcVdxztTHmPP2M
78BSIplI3m1Day05AZOxIpW3fUdAh/r1U4tEf6+El9YSo0CZ0QE8Y2f/G0u9/kO+KyuSKkGD3RWS
50a27C6+Iyqz4OyeOnDr39WJ4CpzcGKOlO8U+y8YvbbfWTmsFXVDSt+J8IYbZve0gDY+RpWsiwJ6
6LTHnHA8DPqx60F75DnNtIeFChqKVr6IX7sxXzFNeM1wCzgXTf3YkFLPU2jnV+BTPf/V7tEPBn5G
m6TyNUuBAfLRTwKEvJTrHq59SF/NgyFY5x39b7hsJJL/AR0QoH7uhBfgV/8J/xuALYqt0RqVtHTd
o2VInIgUdJnLm1zhn1gpM9NzUQY73SiICYn2u1yLlx2tQ+8GpbpEEnauBr4ZY3L40H4AvYao0qMe
XAfTNZ8NUNOGwpOOMBm+PWW8SpT+lCLQMCSgnAwhN249MyB/Sm8LqjbjKm+bjiwAt1eoFad1v93V
uhAv4E7f30p97FfcoEv3IKillyM4jepUspDv26PaDCe/Vn+QWCPeHOtyvrfwHRhOp6A94g8lgiKE
7l/X2cFwFfDrXP00l4+OWRygx4zAWko5zE+HUAnnqpQ4nDGVUBVhJo9//xDIrBIR2gCLRHw6hdDg
td368PE9Upjz2cutrbuQHCCESv25JGilp7suOJh1xLTVgD6IVDW4I0hbVzBhxEnoKNEOgm6pN8Vz
vnaCPEHDATdov/JiyZ7FlIRIyeC7NPbiBNO5zN+Cy1UtI8SW6PikX9FHPQTqnYrMfKn1Fli7kkaX
x8AlNdqR1YtNtE/pBoRcfDvlGrfnJfUTlCX6LlEpTnBU/nCCToa8LoiEkgMPoTGXXMVL1wHTRwNJ
eO9sPPK/IV3SWopoBvGOynzIkwd6nz8gPJvAk/D9Wega6khBbdl9KrPG3hVOMudeGx8FxWzOkzNe
ASyq1BfuE/hczmI0CZEAePZsQGWIvQ3Rmee4N0/aOcRt+bakIi/l9ANZZ97tMMIi+Kk0hLmmq30S
y28Pxao5DieHpH4kxgXkV7u2uqq/N3CC6sr+i472xDS83rhGFFodekfQMPA5wJVwdP57RQMCfT9p
cggGGOKxNlk46TgyI+Re0m+1xM6ic35f/KyLu238WecbDt1DePmLh50x2lwJyC8OzHR1oNiYR42B
Cw6QI5AXIyrQej3SEZDUHySBnMhMkWs1X8xS7E52uR5G5iaANwr2qfEciuYjyc6SbfZVyRy1LMLZ
FyEDWakfAvAM0PnRsvT5gWOgWALJ5vpyajDCpkN72ccXQoTfNq364lSaOzRwpN/wJ8FUTMocMglj
OUD2jkWaK+nk3hU6cyeONezO0HbHVZVai+q2WinSAWgxNsu6LqM8lIQimokQpmn34hJgU8DwmZaC
VZ/bqvMVOSQ/9OMmVUWBMdut1/MJpha/GMnadkWgLHhWtMxfTodE2S4drUJJvyVSwLiaO6CQGh6B
JTAUQjOM2cDVXBYL8dWZMRVBumgAwIr/TyetyY0uCx0JLOP1weOzKw/wq4kfwr/muJDDUCL5mG5C
euYT19Cl+EolQEqMpxfDWhLwIKuYCbtL8o/km2iBIQUoMFlcY6yur17mSbvzUEMMcMfcL18uWhXU
KGO0L/Og6gGqKNG4i/YSx7bC7mvFmESnSGKYPciwjscSt8XHUvKEGJ4E+bZ6inczIKtsUmbWodnT
ADoZIZ2QsLy0ZeBRhN0f3XwpoF0iKsgoOsUStNJqwq6QGQEyXyzYsJrwVekQqpQXGarq7e38dVk4
11YhaC0xG3B6TXHBjDZnSp6t41r6omKym55bpAfAcA8vrMECnRB05R2GDHclCQBYzooMQc2DEgMV
KYgBvds9O8iucIc4B47M+YrgdXhn7p/Ga6vWTPOqvzE7eEDk/WXhHSYVdfsLikLZTnD5RulKw7J/
f14MdOI3ckiNV8EMgTqsofqlPqUopfIg+f3KG0Ltz11ZS7jC5DbGDfrn2CPM7oBxAuMsklyTMH14
BD/gug5GR3twWxov7slPyiISUEe6MWDtpNva8xlu6yxhobNH/DJZkpsD1yTiPzz06NPwdhiicPFg
li4BXNaL0hqP76kJDYNn2eEOzGpgGv5MnAAKsqMywXmtAZn6KzpZ/R5MLIiBuxH9yVWP/DFjaNha
NKV3bYs5U5+U94hIpV6RPrxkWRaBp+XYEQ0+XEcShezLBamx8no32+yB6l0+dxO94rSLLYRrqVBi
qAF1/zQBhtDpPHzJTXLa1Al6G8MqDqAx6p4VHhjNSTfPMAAgezgU5qge9k4YHdF7IoNexyaYxbu9
elKb2ZIzHTgvdFI9pvATfUSG4ljRPvSzv3Ck5Z2MId0Sj9D6GyXBRpAMUIMvUErHTR3hLpRvRXQv
jYyfhmKmlBLDwLyhFkOyS7wMLl5XJo07Uoqnd7+JGwrib18tu9xYVW8evza+aHUv5St5PZBwaa5Z
6NWLH5FY/nNXbqJ+G97zqDnwXDywqeRCz44Gvj4GaeZbe0opAiB8cPQk4caRUujajmGLL7LeL6p7
OhQIPsEU8zHaMWIR/39PgLtmfa1EHnY/2hoCEuxbYsiLbjM/inj1A6LyJ7ZFJjyGDALJffuguGQc
W5Ezw0zSLdwBfziJnQGm7upbl6+sPS6hWjuDCD4hIXNUTYqtoKgs4/dkD93eyQuE1HlwjJbf1aLO
MToEmNK7JEfk557A+KvKqNVSKMdUbOt1OyhY+0UjWxQ20ymMl88eG+KmathP5QpKc5D3UIuPV7VZ
EaVuFuOSMg1tlVOuPZkzlRUFJl1HWEMjWXXxFRf7K/rNpGjYCmMgQW4nJwJsKboBN8ZWwARYfh8d
+AzUgv2OIpWz8RWnSNXVDR5FOieRci/T9k30GIU+9wBxt1moKEk8XdWWbCgcd/ifLBVtP/ktZt+I
CkPw0UvvCkENObDn0XSZpDF+RTdPC4XWYZhOlmGMC/zjb2DTPDArLr4BvLB15UiVIFr74xwgBeBf
XtV68KyTASt5EWBhjlJobi66zV5XHWyr1vTL/tajoy0sLTmgynkE9YBQ69SojYV6I91GV+gG7Qqo
Bi76k4G0p7zqO9CYXVXglt9fUWwExTiTWz5U9DjfhdDDy1ooNLF6lRoODfZTj488EutYGwdFLStu
bH4VxfUsYlTIiBgRzwlXzI+d8+OX1WIoYz76fEk1SK3aGC4u4VV83WteNwx6Onq9wYmrQSlOHly9
+prIakZSrUYh8scpQ3Sob0+XBxTaOa1Q6br5nII1vXHhk7FOhZz/FLUOmTLY6ag1ZjsVsB2eFODD
3ZeF+0S9V+Okb/wfpxLj8T00mizKUg5tw79UDIvmdgsuTi9Ly41p2aWu+VZnKr2KDrZCojsFa3Te
SlqLMNvDec0i9ZOZsU/bOWfcYigOA50uBLprowjqL4cPQOS1OdwRnzIsfC0HQu5xqMCtZpMaM4Lo
Bh19fHbKvC/t6Yk1kxgXMW810tJF9QMSJtR/BJsO3Ybd2bmKGKXzWMSQvus8vpjbxY5SsRKYqN9N
pAGnk42ZkRrKC7XLvazZdGHAEaqTXLGLOO65846PLgmNAIOptIjBDb9/QjLjPedEXU670wIWjgWx
nfP+WnpKhcgs1dWG4wy49QT/M3PZGW5MTjMPwWu+cO0VhuunF9Sy7vRXL3ZSZqUGitb/1KsfhrEQ
cgfIqcsL9nDEqneSFKO4BDtBvML9jzbjpsJYrlY844sFuVatGqggUUnFVcndWZFMeaXddCdhsxKE
OqfLBNttiwaBDgicC10vltHbvpScqsdRfGjIf88v049BV5hH+M41vclFeTniayBKYwB7TYI3Z9Kc
nqF9MXzzc8+VvTdP5aCN8cTl9W5aV5l2KrSuMa45qIi+LKUR2Q+HVepqdCDHRzBGYhrrHvzqLTit
1gEZ0i9PLhOUDbSqXv+XPTyVunn70bLq0wtw5i8Lqe9+ZljaG8WBP3xUVrdMqDKUtzpbhBCF9Wqz
WJtZ7paGcEg6c8fUB1uchEdNslrirH/HnJTDYbN/zjbXjgjWdbiuSI+Fcr5OFJx4CC2G+0+FgEyX
oLkDBW2RHzb83gSTTYKgV/K+dgfRW8Nr87p4t60v57zgVGuyrO4Lb7zYqJ2Z9pazlHC62cWXWhrX
0SnEQ42cLSO7JwFW36LlFqJnTpwBTAlrqsA3HUlUuEgK53o5SBGvZ/g0IAnrh3IskTAOrq1M6OeA
/t2fQp42ftdzWjTh7WTIxSI0StNEpEQ51ziLCu+ZDyQb1xOAVybDag2Hp8ZB8KFpzUSk/I32CW5C
jwTHsVF7RGyjL9BiN8xVcmzhIQjxuZwOs9k0pLUNxbgL4dIpw9zflNfIhc8mrSrZp0BHa5WNVj22
fnPx687OrDBlfmNaHx6lqldbgcnuUnaCuPlZAdjWW3doj+D68v7GYOhYvjekV1GkaUM4JMtKkAja
POva40Gx6/pfthhOQblHdaPsI1JaE4x5MZITfCqP/l+GFrbSRTY6OjqgKlqIBz1qt0huwiSw4zCk
jYVR9MJCwqvlA/rdvBmy8BKsPnnbw5WLUI4gZ7sy536vv0KIssnNeV413bJXYNkDQAchbMgS95Nw
PSjjKPcW1PqvXyx578qUZX/CodpsZI5mUEyzvXmC8lVeziKkoLwMn0/hzer1ZCi7AKkzEUsPlrHf
zDFNS9CaMyq30gEFfKIKQ4mJWpUcHFbCUNLKjGpHpS0QGUohWNtfSokygDnp1Rccg7PxRlCjVWRb
irVj/Cm1wfLlPnz8gmbE9AivTTTkX6utBbeeEPLV9wGgW/dq22JH/m9u6U+EbmqJjxWPUZZpL2zh
DHbTc0Qb5i4d+QJKlORp/2CHwkwbqRyv/rDEAh0r+keShVC84D6pRUCqy7/HL7yAm/AjzkxumlnJ
s/uinOBrQBONEZ2kBDXun7MXP8PMnPDDQazEdw73qrb/awbU+t/L2wSSQAvidcp4N2wFKYipIi3g
1EESU0FgHHxtn3SP/iswIGZVOrsjuaGSXNIZcO7an/RaQ8gg32D66l6OA0kSBlmMo4CrMJOTR2to
PK3wPWOTlTQ/r/o8tlOKWQNB6gEtzB6G+51UXP+GeSivCKMvFRwt9re3s7x1Y7+Ra6r5G26tX5n4
zb/AArgiPyplOdT7ZY1S2yWY5SygJO2RTKza5baLh8/Ue4B6UU3/DI7ib5CXa9o+I/lTBHBesvKr
5u5diiaNRFHQdFlLj7kgRg2bryeKQ/DFhwcysP94gQRCbDTiikylJuQWtpGg5wgXXhg65/rnFut/
p1owe0fZ6Y1p5lLXK0LQKFdJk0aMhgH7fgrZ003s9Dvu4ETSuEnhSSrn2cF3qmWVi8QeiqrfMN/T
RWawyr3Kz2SWi55D+Q/mkYU0MIeVjC+C4En6ajX2Pn0BHFuy5GavcPtVmHM1QopWGScMJKoeXFGz
iSwBE7BL9tI7896tqWEO+vXU5vFZNfBLRDq4iGEz3S61JuKCulbTBWzyEDYi4LHg1k2m/FeD2Sau
Ff+bj/zgAj1fKM2KsMNp8YrXTMxqnxhhthwk/Dv76kXdEi9PL976BirMvLxqZvGrK1WhNiVghofA
GENWBoWJ8SlUt9jbgQnsCFkryk01FYeVkjYpC5BtMvgmGLXycjhk9MkwylUf0uIekHITRK7ixvJD
dF9Zbei16l28T0SkLZLETW6rS6cIx2wM2pIatkvpUZpzdHXPh9JnTTQvfyIJt9O2no+GLCxEVD8F
TeWPSpjZW9f8ewhgQSRTNT76UeZcxvudIeWstZs5DrtpRPj1bTi4JmHOCiCh5hQvFZf8o89MwHDW
yGN6GmHp1kU8ww5ZKGAyqV93FEpIj9rzI78UUCqS5SWkqEoXAkwIbP5/UAUJb/robaqSeAcaNvrX
Pjse+avrtYrYwxrru/0C6A0u8O3bvCAr2JglsYI+h+6kaSvz8BaogbxB8USBbyVa2YY1ChrQie5T
4ZXvxSZQYZu87R+bIuDD4vqMPktLxefPrKuRjAGCnQJbXwBmteFAi5ryHLlx7ITGgQlWwv3CDMqN
LVz1kiw0QcqRNkIKDsjdMSbTUCLicsBqbER1vebqgO8ZN390fIoEWr0r1JpNEd1lNxzJnQaFzy5O
4B12G2EgvatkFgzfj9ZDvSKvGKdn/9hpnq/iZIF/Y3DwzyyJATMh0BuuKb+brFRr5peWFRdmQgVS
ev36cz/L/45WlxLph/iEmjG8UaQ3kBDETnGjCGHzkO60+mxS/jv4K0i4BPD/liiWfkdIbjAiOBP2
zHK9rpnJrh8u18RDwWhKgVG4GJLihJiXDpLIeVQTaVKNzlPhCcM1xI/nvDALeM1faRjY/Vnl5nHn
ZCqWdGmPWR/NyRCJ0Hoh82NVzjrEQlUvvwW5NpK9wQdWjCfP6Z4IgnqVX/0lbei3b5AhXcPu7pgZ
bPZDMdMj3usVk7xb3SbKPaxjSseSLEe6KKRR+uCD9qYeXVD+6q/qVL4J3Xm+wl0EfwlHeccfSbRS
IBCJlkIPlJfEQTywZ+32H9xtrGI9NapRBxp07TVIUs9nr3VsHABosJmg3ZgS/jDTHa21JTz80Nxg
d3we2QJ76XV2EgfGO+ESjs8mDeFMijmyC4t61gbl5BFlv2PFkg50tN4rwuwNJ0PS7UCmo1YYuDkE
SMr5aSyT0blAfpMUjvkvlGIJZE+s4xLMkJBXttI7Reh75FA79MYFaDJuoAlWzl9C2bRhjvLKp3/k
ZSpbN2IINGxnqtYkPavaxmhTUyOyNeGfPlGWQPYXxdediT8kdzbNCJY2YAArX02nLmRcp9vVsFiE
v2humGhIvnfvjNFlC9SQy/JfeWqXObVkPrDt+mTF/y1/LXGedZYCreC7BSEodKLVzLNILtFCCVc6
NXatYUlNwDyieVJMLBU57GB6BBxznXCz7CPktnkUUkoZKqcuXYPDlD3m6d/UE82svCHFLvOQVuD1
ypF9VFU1H23tycrYcBbZkDuMPp/+U2Wz6mW6yfNgRGYD5j5hlVAbTfojeIM4VPfaGqiL/i3/tz7X
QESxc8y4QP9F4pAJ6HlCIy6AOx2I31qLvxIoKR20RF87ndopQxZ1psOahieUEpvRHuc7zlVTF+mQ
QKnS5AoOF3yeaOl3GIhOqdsVkMduzfBH14zGI6PUao8LYZHigP4aTz8oRcm0VfiVKoXVnONVfyIw
ICW7diIQuNZQhaJnWHYZUAUOkPtizOH+qj89G3PxGkG4VF9aaIJ9Ly5S9pr5sJhIinylGLoiwNFB
nj0cuVsK70MzmFFC7ljYo1qcJI3ItFkNNVJCCXihSFy0yntY9JxfYmiI5jlmzMjsVqFZoTktk297
dhm8jD5zt8MO31q8k3KiuuSYRMNBh4WtBs09rla/5BZiTWGUVYWbiOUOmTXQSLQoCmlIAZRYesDv
kiKmZyLvQt7RP2kLQFKGp6k5YIayGiA2UfqovASGvOgYwOPgwC8MOK3vwXLiqojOhK/hNyFXp9oC
lTjF5i0JWeRgNBrdpx1L6N5WlD8LLPFipurpVFyAUbERe/ZN0+rv95M8/VvPIMe9WBmKqKYd/0A2
b1l8TbNDo5eEeLfFr57DJsUTQjhDtytK/dOeb1n9wZXMcro9xNOVBAMJd/rIGcKr/KreVzwBzbUq
OoV+Z7MgPr8EaVQE5do0G4kormJkMojn7EUGi8XWMdXiOWrOxqyn7mGJz9lQEj8dvUoJliB7ptbY
TlCS8vdErFAwmmHJvY9Pb1SFlp32hCe4Koofs0ph4bN2d3k4SG4D4l2jbdzMhEynPOEwbsEC9WB+
Xaf0+aJqtUJ3ukqq8+qy92j8YYYLcgB4HW32lyskjyQ9IQB1Je9NgWuNcJ2EQeGrzXXlPSrK/2E6
LnuLAKmG3w20ySOq1Dopzas+mUD2IB/dkrMRBKjexNRlo5//7JvJzziiTgIXcRtLucCCRPV4AgzD
qYTY8gIgIJQeDQyhcAgn3qDjmNa12NR+QTjshGXlHcfW5jipf1FYJFB9MBsivCFgqZReIyaNUjZo
zkW+D43A1XO8H2mw+jvKfKHgall+o9QtCaWwf4NV2y/ZsNfi41w7ih3D2gMrIkDYgS/Rm+h78RQH
KfDYUd1MKDl4rHxTj3LkKUv16A6s8TcFWHLLz9EtSxPiJOWtIzWZXSLamyawhoVoJ3n7D/umoE/n
schKgL4VBgOeCGBNhONQxPk5wblWki26likt/CozwliF9pL8xOoFiKpYatrTZfBIKuXYQqi7Oek0
HbDgTsOVWd0XbPY0WhIoRzr+PfOq/JU7SBkD50UkcfdiYtOCmA48+BRSjc8lNZRw87jMLu2M3Lpo
J5h/d7v6gIopLM2nUlfywa9YRbNNmVnZETmQ2BMIVd0sjrlIJ6F7zJZOWERHkrEl/ZPnM/ljYJkb
CGsHwO9CtXVZ1bMG0EjLGkuGQQzq/Tjqk4Ftaw1x8L1lCGCdKPdw946yr3yaRYmoTEhBZAA2iFwT
v4Rm2CwfSUTugepZyX9XfvRSniJbkTspPtnCluvb0v3CnOyqGNeAgTb5H6do1WNKscolPsJbTaZl
S5qhoVNJzKL+vHb3nTg8EBDuvIaMs9MP+RkKViKB61FDIiwKFl9mfS/kv55D3W/OJ731/PgNe012
v4zasJbzkwQ7UoP39exWN0ZRE9NXHMZqFfbLQzMLPUkg6gw1AQuQ/OYwPnt3REv24JDNI2dykIfY
OGJ0SLQ+cy8Km3AQtjHq5vDSBXmmp46Gqs7lRqeTdt8xl2MwKEYpt5cqVzrOgUCexSI2S88P3pAS
xVKaw1XxXODCLof3achkKApPEHbtWTn+XSUI9RWIAcYVLspX+Ehno89GuNOws700utAVSh08nbi/
KYXWDJ+gpOD4ooGK8tNmmzqJ/76lq0W0tU0F3xAxvHjtwAu45KzWwP3yff9AaV1jQSC7fBB5IqNK
HBL6CBH6qHpT8FNIHzw8x0f3zHISMKJK0vjLQquTkPMHhnUsoIBjJpAobaUl56hI68kSFB5OZksd
u5picYbP7bikTvWe2/d4JGw3v/bEiVuC3IVl3+LNW6rYNdhkzidMtVlA0+HIi+dzHMCSp9MW8PXz
nE5eCtDtr/yDgygN0pOqO/i0v1DbUbOQiqIB5urVS5DCo4RwEkUDLmTyMi7iGYEAV9AuqDqRb/sG
H1g6Wjt3hMGfyW5zw8XOpM+7M1kaIxORZj8uvEJPCjb9ueXoYIYR88Lc+LVNobS/61YDfZ9AcV/r
F+tGe1VcPzxQR0zFSw6CbeGLPoL167j6n/iLY6cJ/eNwjI0mXB81ovkLM5WZmdtlFx07o45HWfjR
Wg5K0f2HquyrSi1koIHhOlWHSt58tQ+iHoHjuyotzMIVY7+dcWoGaXTPD6x+aHMu8A2Slo+5xwYS
D77AAvl+PaA0c+zFADDSRrfGyTr5He61yxKdaSE0boaj2OmtKT4ZR1yDMfXm0RdOWE8O/y1DRLW8
bpu8vwgtAQyMOktuWWIc6yDAwPlTsfbvekEFGZXB44KOFCLPzoKqiYIcUGFLeEYovBa0kVEed8S+
Rdm2x5Da94hFN8Ag3QlnlLIdTiKPzTmz6jbETqD9x2fV+n7A41gzh9D9f9qWce7fstq/UfKv+qnY
BE2oVrK5U+BioKoKdrmYtQaH3co2PaHT4RkGwjvurnK+qKQVNtIDVWI0ZpSM+mOfPPirSsMeHEmK
SZMjcLlwymAurOduY9ozsS1s/iRh+yS4o2ehjaV0sdms6kkT/PVl7Fjzq7apJxuVo3qEHLtdg+Kg
geEePZqsZtnDFB9VHlzx475HlfWLG+eLuZRvCS4znCGEB8syEDMh5K+5Q1/hrhR1L+ttSGyV/DHi
EOYa22hUeoS8K/UHdXWi2791oQyWM3cY8KIVLap6gxMeoJVXD2f6ZVVIYnCAQwUcNuLM8+EZsoCu
d2ekXlx55v+eTYDF5XDd3uAvnjWSDLX18z+jSJvHKVjlOhgt3a2RBBXSmBxagJ9svF78lY1zvtYe
mcdEmCdAAFmD96+YcqGh/HEoC6MRcNZPK+f6DFSClFv3wT5rKARRRxq2ZtfPNPZxX23/rOr3umOH
ojOJu2Yp3zDH/MBmESbCtRNxlfPgfc/ohlyzfYCFLad+V1y79Fnc5dhfzwJbTOG2awcRJqoeeNxq
goT69CaXRF/XYqh8FzmAJxpoYvcBvgw85ldmuKt5GjU75dc6jjapaiBjej9jchXOoGnwaSgnbjZm
RPeRr0sYCkR7qVJxdk1zij2FBB8DiCem3nOOCc1+HsbK0DNoWjKYQenvfRNf2Mb/ckdafZSibeBj
lT4tyP6btYXMpauzjEZounoEQeGcn4QKj4l8X2k8g5Vtgb81huMJMBOmkmDwnzbb96/Dzn2vtJ5Z
M3WQXWe3gXC3tS19o26Ksia1DGzK3uNBVdaS5x9Q+V1Ko4ELYB1f26IvlC0wQ+PRMyyjP7XFefKz
OiseiS69Ym2tpcMIeUGwkxCcVOsMoSsIu6nsEYCvSAHUgV2sj14hAKFAnqJy2bZ1qWyIE2XjB8xf
NETufbzv/SzYA6h4M0ykvAuwCn3egE25Aewws3IcbgpVf9p0TQs3Bn/SMxHYH4BsRJ1bObvOSxNh
i18JKrV2g2I/NBKVkf8cIh5rdxXndyqSvcEB/ZZCoalYY0RD46vr0AkGjBy1kQk+fPW1F9gM6ixC
NJ9B1jtEoJw/Xz1MWep6+j7nj6hxylZIzNO/sAri37px7n3TPUgTZk07UBOFh+/AwmojCFLwqHur
pWynrvohlvFiSMaqJk+alaKCDsSN+HbdSJYRhxljQqY6QGMdBO5jARP2XsX1IQCdFKmSo2xqpkGi
YsF6bo8h8CqZSfsPefwYixRVSB3J3+L666ICR/x6naHFyWYOKWFc4jDA0goF14kPoom3OTcpLaT/
9Y4VPHIajh2QhQwcWB1tnimIU/D86lwLESgVwsygrrRdxVvvAmwEtaDCj/e5Rhzl4mG/OSl6Z6hm
WGuhDqJjpmmnZIEHdd4rRRXBWzoDIsAkjVzTXk/K2MCetxsu5s1ZlOqB+Dl12OoAXd7RIhWmK+DW
xeMOSpSY3TGmIDzfV5YQRoZvTPr4IDZyRlnboZrJj5e05/CrMzbfm4XUWA8o3EyGijC88Gz/j4pp
tsEGKCJG+uQVVUvgb/3ZupFAX0tOITuppL40oEqOk1fdwJJgjA91S/qNGLGXBEj6fI6vr8GNPxVW
9BYxAed1+qha1n3rkxLGJ7agMKe6OmRq5pj5CMZRRmjHN+g4zzSrlsvGk+Z9k4xgA6048ZC/zvx7
xNIU8Dg3f4Fn+neJjEChhqGaTS0kt9hA/zf/OsOSU6RNlaJCXPX5I9jH2z9hAOh7w+K/o8B/Qu2g
EJ3oS/UEngy+ZHOr32q2JzPRU2dcAjifMa8wheYq2mu/v7rmvzWQ+PyoAaJfHItCt0QuJy1POHB7
xabPrqDmSStBZ/6h/fGlbYLb5UQTbaFXRg/jTbnyF3o+rJoz4Qa1ail7EumJiCjfClOewLEgDtBN
rsyMPg08fGaNbmRq3CwKINadP35lf0/e112iX8bt9xZ02DrZCNJLXZBEaYyRu4+d58CV7VkZz1Cj
V9ljJfD2nJKUpAxDoM5ROxsnEtjeMcGmC3es1uzW0Lgok24hEKk2kEf6l8mKS23hR/Yc1mT2hhJi
/YguouVKM2iMvBxper0ilJGbBNq1h3pgCU/q2HFRxTllIX8sk7Sm4owjRmvBgT0i1PMpUCHK1as4
TjaVvqLsmbEljhacHvlWIdwF387dRJNrmWXoY26Yo+OvwXPFJ7liWzzwT/uyzUfCBc6fr2qgNw8I
v6StaT85Z+c2c31d4mEnAzqtWoeE9CQIhSAIgA13XJrrbmXoZNfCHnlNGTLR4lZpeG3Vqd92jyhO
n95DvWQC4yH1x4067APCEtaEwh+fYlFC/aUMzIsgzd+maz9FZ39XkQH2WOCIv8ui5e2X2O1tR7no
AoJu3b51SZp61YkCP1hDfikePWpqyQbFqmx7rWBGSvueK++F7oKmhzISp183LknHLtHvW0JGLGhd
vzRw0oi0YgsY7sgPkh4ZW3FEV549FMGSZ16brtXKhe1JpGXPLD7L/zjXNco+P6PzhBaKxvhdHT34
5lJdGuRYZtIOaZ9SI8NPA+SYzmAjfV2f2Bxs/qnCgxlRnZFHDOwXM2tEE11zJ3Hz8P3MdELftr9D
LUQ0Qu9vJ3328cPs4/UV4+p4/KU+sho4dyeJ2xIAoAcg3Ti0u6djO1OSn0jpjkocv+ZS/nN0Y0bg
+4ilj3BjLFDZUZvNoiEZORVZfYk/3Qohr5B6vW2Aks/k6pqGWTwaO3OdjYnoQHcX64Wp/LL68HQM
gX7OyxnU8WsT5lXtasKm/IhV/t4veadmqNGvZjH2L7pBsyzkf5U5Pqhn6+lO88cTKm2M4RhzPK1F
RoHK1kwN/kGDzRjMkIWm0bRScmD+tXAeUQnchYqVzm2tkr14NFCZG8MEJq3oSRbFmTzFf8Frmdem
CuvFGa6P+G8kTCF7uJG32N2Q5/9Cu0IWTJLiWySrDpj1qS0c5fNvaKMEAWTbfY9nnesTOGnUgCkz
+QM3Fthtd4qmZ5Ise23G6/saEim/8K1FYPe34z5t9HEap+uaSvghnJvtU7I6HmxXc897rwyDfVvX
h7iF1QZxp0cj2aBOlD1LOYGM6RhDADPb5An7Do5s3qnADlJTHl8CCQMlX3G1ElRP6TaG9BVlpcra
goUKg5ZUAqvheWEsaLZilcao0dWm5r//ggIHq68rCGXpzJ+a7/YNlclzoHs+Qiv1RsdNSoNNMU9u
irim64RGLRYMjp0v5PXFHPC7ptL9Qgjib/9ZYJ3gGlQL9lljVLHS0WhYGeF7qAbVqgMLunfAHWb0
6JzFXi3iFjQIdm4gNyI0/9GUrrRrf4Am36BUA9Xez1NZlsKtQ3I0pUo5XWOgLRfvZwdr/Wd78/Nv
hb+Xzmf3IW8qzaPCAK/qj+g5QFLd7KEJb1lbXQg2ClAedzW3X5FRxEnzQS4t4c2YTc3oVYLPtU6q
V9Axuuh76agglSPNSakgzIRlYmDHLlPw3VzyPVk/p/Q1BDcpPwT/kLNKZx327EcmizDAy5SooAAF
XOQdN22N1ERmK9sn8celtFyAdQJL11Tgzz0dUIsmGH+TwGkUEUSsGHpmHphtWW6YOdGD1mmHzCI/
jAoEE48oYthfBXuKubs5Xl4rRoU8nYjRp14d4uaxteXWD6QnuPpoLqI95u7ovpKw7iNn3fpjNm29
IGd7UsRsgcXqWhB1Q2X/ATwnzByADVczCVuSyQVSlCcPM4rnONlTgQOfn2k5wPCrv/sgtbWKqRyM
SW7vknuJuGCnlC00GbHkCiIdLiQxh6wOD0EG6uXwVhu+Gn2Za+2yscPbXDxm2gXXKvlTB+k0PfM3
5j+QuIbLSrLFQ2PRYpven1ElBOZdkHczIaRYiGaQcTFPvlBPU07WL6klhtZ2Z1DHEA3U3SQsugpL
pHBWuNCPVu+iaOjFVYFwie4J2AyBC8ielVBvmJq6iJrJCzAj5e3b+IVIC5qfnpj+U3hBQHvXDC6z
L/74j8PJtZMBe1wM+YmrTnINU3L2XG4h321oQf0TCHS89BWPpItGjkefqj+Wm4KYlaYWUhQaCL4w
cdCWJMPODs6zY4d6vh7j7MPqduHf43iaHdMowfFRUit8XErbj94gPRWDFRQH+Vj05bct+4aHCMh9
6oTdh7M9eG3hU3H0IGDzCstJ2rmbeDz/Pjk0mYbaTbSM/eDEeYQO62dlFtrxEOyvXss3DL2pOHii
tAFTsdRgjGFK4VEQ7JccmepoTbM9DPWfNqh5p63lf+TgxeEzihivzYCermk2FAiKLxPx/rh+jSh9
kFwlQllyOZ0Hu2M9LpnrL7lWiPyl4AWw7QRiTBYQzaOZTIZlkt6O8FiFqeHJLdff8DEXhgLf7ntd
TbBiLwMJbYJxiXU99wReBxKN1xOw4X4SsxEuEJO0ULnuTVa9D+IuDYGHd9vd+PlZ7a2cQhP0+8LZ
GvvuH9Fm/beSHzcbjLUKIhQBygjy9q76+y1I8hXe/WImIzPfy51HpPZNjjIFduxu9hYMGZYNwiWU
Tl+JERxLPKtENDrhgp2SesrvCMXumFPknZEV424IQaxZeYFaNiccP5BgK+lF2ZVhYmS+LyRhAwAI
Sk7u4TsT6qGjgWiSsKxOJE+3NpeFm9LO6X+G2N3vlb93Xe20xTmtcsD3UqeUk5vqBGOBAhGtZpIX
kqa//psojhC+xNbhdKf4XW50C16guKRRy3+b6Fqg/iqz+sGjGeyM4HXkxXCoaYw4kWSU5l4FNMIo
rxXSLTj2adI/rQFWyZUpO28DNaDWMJJIxZTOm1kcedbA5OiJakP0o9hs5qZs04Bxj4dO4nPhoGFQ
IThHpdsVdrVM1TdJglfJnK6FThWp4mxL967EUXMK1qCr6ZCyhKFyk2OqIWNg9wfYDC8oFN1dswRr
Z5RXEGOwmNdurv6UlfC76s0V44b59wjwX+Yszp4SjC1JVkzbj4Wd6iOu5ZJkrOnUYmhxq7af+JQC
1xRz1NJ9qLEgdwqvj3IQNIlmSuxK47A+6Xfog94votJ8nq6kc0ZnbY5LMdFNVE6Si1gY8e1Jc06X
KdMTqSUfdHdSuRHli1THq3KH14dd/YEktgcjnkq1BwoHYex+cqoD0mgme/I220cU7mtIrBq1CExO
jZv059YUbcuahOQ4rc6pXgKjsJbAWe64OMXwuTV4SRhoTx9sSDRh3iZfJkDpeFIlb1Pt98jCMyvU
rwdRG4vDdMiG0akZY7sQV76IHiysLRK/2ym00AtdUKK+SxIWRQe7obYxa0yl3QQ8H/TgTZ2kuSUa
VFC9UGaAgIoSoqyt51gMl4CXBb2biOMU0Xjryibo3s+31kLJYwvpH56e57LAwC2hC3ccRiKGFbL9
syarNXI8dQmpnGX+Q1ULDow7+ZzmHjpuH7gjX3IDZH//4A/bkLJvqdsXgfhshfUNsevJxhs3XT56
c63OyMypsAqmv8E+9/Suc0MVnG6mxZwT1IXQPb7TENu+6Flkm+oh2plfqTTMYWKG0quP+i2vI0Cx
i7uIJtMkxmpAiWsSIFxlFIql3Ws/zdo3AREYsWuYIainKYnODqe2lff0+27tieoehArOT7zM3sbF
jPSw8Z8xK+T2jRwpGNdhUcLx7Rfo/ZkSN6ktbd3lvgT9Xu+LLPT9YQvUgowKgIS17zBMTkZq7Yuq
Y0pmB2LwTADWnsk4byjVN99J5DaJeujxqOEn6RMevelX5LlPxUA=
`protect end_protected
