`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
kA+ipdqYRQy3NPVtmKU6jfwN4NIHjjLzgZ2O0bBMa4aMY/FAqM8oS69YBmkohQPtuczhEAEqSxEy
5x7MB/PfBA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
AmgJ7JpCiiivwF43M3eDIuboCi/zvH9/C8VvRuHE30yW75cJJylOlFHPbHAOMRD0dv0SI7/fnQr9
MaE1uNXySOVyESLF03UH8V0QNNO+Kr5zj02fzhMrWVaGYbFPD+cEw88WXFAmXCx3JddQEMgB6MqG
4u3bce2OyeED2YgQGP4=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
h5y2BoDynYEBdK/Y8MiwopN4nNXYz3CekEbTJmm6pppvfFImdL4EVOnGP34dJ79i4gOHoFBeLhVb
5RL9b65DiQIW/nKNTSu0inNoOp+IvyFmqfjERJbJzrbPrRff6hEN22abX2dTfFzom2ObMjV0kEE7
gAnpMdeQz29Lnew2xe409+LIGuyG5q1Bk7/miDhvSyCVpeSrejtjSZpWyD3Bj8GASBVYrzCRWT8w
SCi8Vts8rJr2uiMt+ZSwfimaoddMgE9N5ytslN6hIxxymoeoH7fDmWLPvorWpaXxzE3O4rddpN82
2JVs6fWtbGiCXt0K31Vxeg1y+7awXFjdHggAqg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
JoESiuc05geZoBgHD6/E4dt4FKjaU3E3jDbfEV77HxVsIKX9bQ/xTpEKUytUMu3Spy0cREwG9qLu
wY9jm0i4XavNWQnLrJ+SAJyyAvfqgmwnADcD3xLHN/BfW9g1K5ENK2yo/J3hK7OAZEIVxFGAYU6J
f4NhDBNOM6EiNIlqc+g=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
1M4FfCyGwD8F+5mMM8Rexr3c/KMPn/MyTiR4sfjwlJq6BSXkeGmGpwWWmEerpCFtIhYL8rD/p7Hd
5AxKORNGcAv6aPSTV+3sX+6WpHI/XHmdhFrVdpcyJyLOp6eC9PSTy4XvmiW7AISDzeLO3/Ww0FmJ
uSBkqsrYiavxEvC/MXJ2pElAS0zd0n6QHxsfphgL3T2x/s0T39pWzsbZp8Oz2yZusKDtzuvQTTVH
Sy3M35sIlqqlqh3uU2MTg+LHjEy7uZHmHSACmJR5150UtQ02ZTT0gJaRnljxdZW5/1NfuPS2rIvP
y0XaLcssR7xHms5iu2Xwz+/nze5c08hhkprOeg==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qEUqfOScMNowQMFQ7cnHO0lSH6hy+wmkM5OVdcwFiW/oaXLND528bwpqkEuSlHnn6IZR4bvTB6L5
uCqhY0vXBfD1rYt5R/CHX8k4QFv48ILkmF3q5tHibdwwTSWxWHYvR9h0ho6gSC+9BR2WxnUU4yKK
ti4pytetgPHcBF+KKnc6DoMztDOmMD5bpwKPiSgEtHU6k8dU94xXedmyg1XIZv2xneyaMtkQuxX5
O2B3o2duDCpiZf3vW/Sklch3xgj4aMTf0F9U+/HJ1ytw9tgZBPZ7CADqQdr0M922p1jO1uSEdlDX
7Rv8e0e0+0ebQ32zeE0v/aSRTNio8FDIgGWC1A==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 556736)
`protect data_block
48Ug2gTs3BczygN62ETfI7P20o5e3mFF10Lc3ZhLPrqgJWZYnkTQNHzZ8k9ufwxiE0VGlyoKkYEZ
7jJ+21pnLcUfYdPZFDr1MLpkY0wkpmi91KFoTdYx7JyzFNGv0qkIljFFl8DHmfhmj4WGmgAJ4fJy
wj1bdqd5OgdPGoilj+jVtjvOSSWiD4MIW0w6ox2s3/YdZuFxKNRW3b37z3xsQMJGRRb7njQ7yoR4
QYnftypArdivtxfmcESLoy/Qrijep/j0qiDmrqEBvzWgEkppJEj9ZRQ2MfIEauCwv8j7nc7aM5qf
R+x1ZOwGn/Z5boMyAP+6CGLD44AsGRdQMXpEyFRoyhkDHkgSu5KZXEI+FvS8wtdaQz3MksneECkj
aA4IqHUddZg4kY8Jcat/E+jWWDHkztsluu+UMJmJJ2xDvgZppgnBLTSOJKEPZ7YRk2gABq1z05nW
YTJ8bmnpS4/feD52cUL5rUo9mMl4w5DKH4l/xJxtFzch7k4BLgIEdodtJgIkDKrlGuFWoXjMmEhS
GYQFSV6tmjEM0fONj5PK5ejE0W+SHChW5d41KXRWcgGZz3qCk8i+lhF2PPq3FMlGvYo18TxPOTJ7
6ZW+jz9ToNyt8jNk/wr36oBR/alnIdLXuxmPkaKwtKGhOUM52//VuEdO/6RWoHvT1/JlZ/0BxI+G
8EQNjPeSjc8Y/tvanJlvPW73Um7Hoamez19aFhYP84OkeEfPsPO4Tkrfjz6+F1IiZuiTFqXJTf9N
oFqn7KwKb9nI7ntQA9P15b8++b6s2OTSNozTdObz1GuER2UkkUH0kH/vhdDzoHBL9XbYzp6NU7QY
oo2f1cYp1QLnUzP1ILS3B8Jnw8jjrA30iJmFQXE4l8McB0Zm7PfOd+5nLJtm+hHeidZognHDZ/u7
xRSt4Feje8HSFA6O+Co4y0ChLgjjKsvHOfUGWTqgwaf9GUg5+kMTz5Bqb//ccgI/jDkAQOliBgOz
d3yxzsH3K92jO5Y9THkbJmJp1sKIXAaWp/UUYJo7bbLNTwKTtRh2djMXOwDv3luS4PpXwIOTEmh9
RBg7vRgajU+MV+Czgp0KWoVZgQJe3KSZbQH3yHjgpB/iYTUU6AVp8/jk9gSnR+GydeJxITaZq8yT
Dc7q6kxMDzMb9eIwB6/gkDQBsga7Q7C1bZ950FoJafgQ5DyI1jntafO0mBC34vUDHKnrqZMavOhH
ddkHOm2FFDsC22+adbbmJi0U4dFUUJI8/0v8p2WwvH3is0Vm8Y0TS4veCjn6Z8xHIbpO61EAsL3K
xXNKmm7/vJ8srpNsKBZtz+ctuygGdoV7bUl8XD78EJH0clEPa4UqhUeKTeEOJ3Urr5GfmCblQFTE
V9Jxoa4C+PPDsvT78ve87lfBPitPqG7LpeFU8qiK1E6/6XOL6oz513U3QH1w9znSlL5PCBk03BJd
4JdD/+pFWmwH1BBUJcJcdN2SKbHT5Iy9FFcswkYNLOBfrsasdVN0wH1BHB92kiaVIdALxiY1d7Al
WLEVXKVQ8AK60zo5UBpmzcRcjwJ9ZM9ze5SfCjPtXANhSF9V83sSDjOkDQjG5CdB4johAlCAok6W
EmWr2xxPCdhydZCcewAw2wauSmDXYVHWQRbfi537fkWWGFSK6FmXcUACDAfB9+hDocfgZa4Vno8K
vYnNcDTIHOmVm5U0HMCsb3Acr1KT9GwGttg7H2lQt9PBsInoBb7gRuJKniK4ZRA/alL3wdPh8h2c
o7iYRKbdXCMoOEROTug8hXvqNEMnsgOzLCWkWI2E3A6I8wwdXdVJh7Nk0IpnyQPWqi0S8u0/Vvdm
2iyGVwmcLJI2NSE3bjrhppFWEQ6/hl0X+aB3EjXI2q7fdnHp1A/fu42mrSX0grm7JlfW3BFzW3Yp
WL4o3K4F93Z/D4LOvPMRa43gcmrD4g8ck//Ve3jPIcblhSUIOlokt2nFzFzePEvRFMi4OzU+3M8+
UfuD+s6yLghBfDW6kC0gxlGGVE/+W9P1WMzT34xD/dGDxwMe9K2FFP7KN8tvq2/LTHl+Vue66LmR
q+vLLC+HjYeN6QwnPy+GUkNP6NAG0GL91srTp05jiuhcOUM9i3Btje3fv1B/yvyZ/RCqC8e0OAoJ
B2dZoTJ/z32+qBFaNe027X9ozWMqzUSP7p86RhYbo1tWjfY9Sh9qe0n3/Il6fUnbse1PEG4NPGwd
WIcNqNrGrpDYsBRw+CiPR2S5PsC31ZURsso0zZ3P/tHn1p9eg45qiOOra4QGyyhphqNmExmevmmJ
FKIkVhtTvraEhpSjPlLzGvA4jb93tGNg9yiMiqqLUAMf8s5n+86zKdJy0vNKZ8BIpuMwKMgBw0i2
eZEMTxkCF/J1bl2qdQoXHZY3Yq4dW1Zhx7O+fnODYTiK3aPQ/9EFrtQtp+EAbi8a3DpY+SaigqhJ
3SV2NjDZJa9nDdtR5+8ADU66fdSw+zgClqUzmNMzUqfcJWcOI6TiWF0jQ5vQ+PL6ivcum4Pp3lB+
D3sROZN1lWuZEaJtHFUOLyHtXyMEEfdredlbVHNK/s+/6ew4r4FmlM0zdG/bePzVMzkBg/nQsQOO
JVFwbFjmR2Op46MtrLSL0YCsWrSk4bsh/IcKXtWOE5Z/k9tBdpIcD43f0A+FFXCKysgh2n4J7xLx
wIechTGch7QGzXuDc6FM2PyE6HwXFgMK5fsyW1sMdgRMLSxnNFLZIGMvAgZHJUOgMmr/a4lwjBaz
2xSyDMv5eDI50gbLaI2mwfpJFVeWZFZhN3CvcEwSCvDNX3Mj9ijX1k6dj8XdnFSJIp2V12qkZaAn
DeUp0n+UYkelch/rP5a6DoML0+YVUT/EKeTz1SLyEBM7VNmcvXbLgB1+/jjCMtxVLd/zshXImVwL
FNN7EXFFSRzu9UWmX9f9ZTh4qDT2hQWf1OsmchZzwtUjgM4QapXuW3k1YJooj7UFJ1MIPUi+Q0DK
Pyz3ya/oChSqRbl+/ZG7prAPJKTb91hqNOoKUs6mwLt8fOE0z9NUaYHVNIQ2s6MnJXW7yZ/N2j1x
g+/m40x0S2Aq+S10CBFOi3GAf8WKPrDXrfqodS7Sb7XIgDq6HVLSKLBOG0+cg1WtSwJ1ufmibFf0
Eb04vyiQSZvggbg9ia6cHg569PzMENx+E2gYoxaUImz2LT50zQfRf9rcqik15pCdC3a1BRaxYqMw
qH7ZLofk/q4gHyeN1wQx8AcJFzGoZFKXzwhalv8odcug9HuygQmRlfF6fISPkw2dN/TMgRR3fYO/
7teysoKXHhvhIPpTyYwCJq9hOKvNgXQfwQbgKHbL1p2K/L6JJiJKqQ6Nc7tR5Rz5yUF35eNCzpuM
2x4ju+itgfVTE1Z0dTUYVSxOQ/UhZ9SSajQgQIvwqh2xC53FMAt3KaCt/YephyigSsUZRx8bYfXL
zAYJDWzby2IGuWjAfgCfuEKy8Fxx5yK+7znQ03plNwa9K7VYByAB0DdjR3gIKV79Yqvu9H3SX2ZJ
26PAS3Sd9y1xco17yG0HOXyS+GcEWWRWJv3nxaFQfo1wdL166vs77zrHqbY5dn7x4LAdAx1qzOwY
CuErgM7+Q9PvbIoO28YedAFkPDoLpl+4+DGL3P4ZEXORTpiwu6IH83GZLzDrr/gXJZ7jdp92loqn
FGrsyZi4JRdmNyb1ntxQF3zFH/ETaXJYuYx8Tm3RQH6Ro9k3dgpdtjlBY0O1/N2+fXNDn5tjR9Jb
UKAvGuqyp+Ez9w5KuHOaQRngxR+/CN9prIAqxi+SGOJ/r2K6TJ/KDh4bqNviwG8bauEKM1IyWiEI
9jXlb78jFTZgdrQNka4P+CUVrmbw1kjIeV04xMyQIn7AdgwFIQzwRVYC4xnBdgHTtCY0VrMV/AH7
+XPNd0/LhcR68Sin5bklFpFS5QpjCvLvFF9VTfqVvDE/wsf/smIHzHkLZ2pavBO04NfkboXOMGTO
yBZg1Q+p2Jc8JyoDftLr25JIwir4XbGC37RrtULOIna9R0T3gTf1BNV+MKpY6uERx3RZzYbR8483
Z8mL+DXJnpG4N1HSFvlU0tDD9pFINyvrPpUqEViVGLAYYXuYAuD8Ozm66/1kqdbuvtZ0lPN1hgpq
IS5bJGH27ULXxw1YRJZ3Aw7/RW9qIUsQDRnjJwYy9ed9K19ei8ZaLotzMqA+2wFBJAIO/JPULyKy
zyKJRROPRueLpZ/nBE6dqOqiK6t9HoDcppYKg7zKD9X2a8/7EVo7yS5Iv9BbQpqIXwRByZjNo9KC
N+BHS8kaQFVow4MFGu/qpWO/99bRzpW1BNOrxw9UFXDDpdXXBpMxtSLmMrsHlmJdXpPbfCdPwKTG
K5lEbMQRFVbFu+N9bxBR1lLPVvoBEmABqRncEiy8KBhgRJYv3mgQbkS03vRuLwaJNU9uUKfvdkH6
lLwZ/WKXncEertuKZknft7UYhfuecANKOv/8UBMuo4450Hovj1R+2xO6y5saPxsi0BwbqjXGoIGf
vqcWVEkTp8hvCkIQSfmIyKNdMb9f5jADKGDe9oCJHtAp33QMc2ZDRb4os3/y9DCMGgpcyLQrLrVD
iQsX1pMI3gy+XzVk43H/GizQPusND3a1iRItp4HHuXu+Hg8k2Mj4VbhF93BeeoKllpqmjx4drxHP
kJr7JmgS6nFNCJKletLszYG8+J2RgR1Ruyd87gQcA30mGUxql5FV0l1Zfi46VNZj+l6n8Ou8mIgX
xuqbZM8RrBjuEp61C8DlwxCGEVNGdwru9Z1N9tn6xya73b5MPQFh8o1+p8WxfTBjOp7N8sLjQunM
MJUCGgJdw7as6fhRU0XQmS46owx8G7ML/oaNoBEDtBcDjlTt4ZlQSttpK+LXmeoc0QK3gNRpLZIJ
9I8FSXeftf3Wz/lEmjGcEzws1UOAxUVCeLGUsMXJzmHvBD2K2+fRlA2fZ3pQ9i1XoiB4Xhy0VarF
pBYTDkLW553XzEsWo/mtciWU+qDPHUqGKbnWwFU4sbjB/vBPIiOlgbXwUnnUNcv7om0G0oX6TYEh
TgqFPqAEmyLFKOrTd6PCQ+iK7MyUMl/JcbpI6ReF9wGUQ0Znw+eLG6gJrmZLRkCeJkmphfbz3tB2
6+oWKaj2vagFfyAysw6cXjsnCkd3V261ob0NfZ5aFd55wrVi4e5vk6GLSYr8evKvaoi8VfA19ju0
gGAHSUTBXnDOsta9i5hCVxbSxvvfd5eSqClX8Wv4xb1FmJI1DqvAM8qCYRllAn1RrEuGYyKC9X6e
5ZOdA+lX/xgwBB0eFKx9PKmzDk8/mFt61Tr6EWGqOjKIs9/OUf69RNKtnUR0CzPHM+pPWJxy+MM2
qBktm3UWMMOuMZAy9deytvRtxXfHPVWvJTlK/w5L/KB1yJY9vyL5OiSNC/WBmBUSyOlQ4SsD55+G
aEYvZuKM55foGreNtkE+nlje0ZjnqsP7oRbNPFIz35WUxlvuS8lDVG5di5DBdfCDhXS5e1ObFH1l
sG7ZZF8LOwPDEJUVR+CFxTJXe88YtDx5UY7shPFWM/24vQxRzuaLMu5jbp1IHsLkpPqNzEQahEga
tmlkpcl6kdBL0JdqT7z/Jw0yDjNTHlsFBGsY15ZRQ5Mqbb8XlwUUHqzzuFEnzejg/hFtJQqigac3
0kNqoDJvq/qXUdAFZqIfIswtMQWhPy10uFcKkgpzVHM0Hx7v7zkAbfYo5w66gCvNq7B4oo5T1CJ0
HTKwdmkIF4Wj7P1MrcQPNipyt80BxRuSNCVjpbCsKvaOwoPSe7jedbZtlTxYDd1hcNDgAHT/Wwet
t/Eb57M7ooXBik+PEB/ej4TZkDNJBLW62liWluy5wRASvgJDrmctnI1NkbO2bUtx+oaQWLbplA1y
eTaYsjc84tPlF9L2DuxFRXIEeSvqzurT4YYE1b0tcyrN/kM8qNlSB5EKVTwCe1E8Nd7nRja1NzrG
QLspBhjgT6ZWMteT4hzVMTlrGBviyxAYY/+r6NnZlb7c7NDTDpCeqyCjGzfys5+dPEgWsH3V6W0P
zdOXD0POyet7AY1XznWfUTdF5mIcOLvq5KnhwvuJosbtqAGWXOjpMlTUjF+316nrFJdgpqSAi4Co
bLgS5BAXgm3CTzt8DQYioynYIyv27BBm4yxYvrisrGL6/BzTrzZPrIrQDviU580Aghjve9TpQ8Yn
q0WUEY/iwbCec6VEsc3w/4WaqlidgL1wIv6kIxLsjJxHHGDGQZSmGpt7FhBEz0pzSNfXIG6Z9tSc
OdgWVC9o7PMyQr2YF4vMfLP4WqutWpyBn9ljNRRIngSRbQ48O4786NU4OCON8MdRlem16Tw/H1b4
ivWbVVFR6C/hUH84sRrWu9WY5qzhg8dU6dLp0TD58b/wV74AwkQqAmOuxWmHUnVNHurrfs0UR+kG
MS2u70sPZfUuav3gfMF7h8i15cwHFNl8MhwdJT4IHdmUBDP+AHc3aiAsZR1UiEao+cyntENVrTiA
qMRTKd1UFe6ayRg2cHrDjJVrzgMJH1M77wDvTBjenEE+tJu71P9HeARqhsz5ObTdunmBUrS0doNI
gZ6idycGHJDmJwV99RVh3rapiltDqadYNYAyUHBNLAczdg6JmPL+2UI7gLX8ben283t9oX0AS/Lu
n6wbeV+0/yWbb76VmMZjBeBNMjX8aYn+nOEuuchtLpHWC+hJ2XucQY8hoFLyU2zbWDR2KX1PEdoM
5Se46n2V6Imbil6x3UsYLjtYWm3bXmOjbRn0LnYtvzG2gu2bQU0TQxAMU+QUzk0YM897VQN6tpKU
dnY399OTV3e6BNF4fGLu/cKtDl+Xx1tErPAYjmMIoSWaod7FTRFP9+4DjsYc1Grw47fgP69HS7hV
+8b5Xb2PZkuxaSWaHxc5s38bjc6px5rrq8lCVuRZpM7RmJ0nWDORtHh6U/mlqVjwbUA8QqcERMIX
a4b+TgYVYt4ZCEaZGfwnFLzviGS60p4Hy475tk+T2ca/x4XYbKS5/cpR5jKQrBfAUV/F+vv0UwMe
6yRMXtAwOTHDILiBHFCXBlUUTTXDgqxYj56iJkx0/fghICVNWyqtYOQxKaymXUb+Ic+vsQhXkcvN
bW6CS3Qz7tzKr6bw/1ku6tGmi7ViwgRAK5G1OiFmPMUqotEc8//63GDhQXQccUQECZo5OfHpItr2
pe97ROJhYo2qpg6MfsBJETtMxCXdn59I4LigEyVGJFTejIEIKhjF/TAmuAar0tOuoiOahLMlohRW
yh0ZGhl7l8f3ppHotHteQ44I2EHELopJvJBMNRS4mgwQqQJPkw/k9hV2L2DL8y/YhFRxu+Pf7FzQ
k2xjwyzadsI4Dy31fs+mfPHPnSrX8h0XLm41umJFvJU+jsOJiiTbwV2jgMP7jB/URMDN/O72kB3c
BIOvrE40PXtj83NVxJAYJ+VOxFyuD+OD3FC3FXIzcszyOlRBHv0nqCsGV+0BHlX17oT9lPxPi5aD
dZdotm7Zij2OzLcpBGD+/3HhFUHOgbjIzT2T/mr3jhc1OJkNLk5txwaj51PJly1HNTEl2uT5zwwK
wpJbXe6yvHKX3g2yYIS4YCN7/B95O2diQGoalc75HFmRGbO6jGvlZnrjezdJ2UkrLDcAg0DEaydq
0V0aoLNlWgyjY1xfS1b67q2AdFPKfEI83Q0wW+Bv+6rXlo4mTkCPk/3jf6THVse5vRIjXzl0WRZ2
v/lY2ZrZj7+42AAlZLtJhoNQHNU9XtZ19EyKWAW6ZkTiib7WfD85a6pBoj6kRpvt/fBPnGIHRVKv
f2mgprxv9TIDLPm6h+hzTzSto1JbopNcTXJw9n1QAIVgpvJwq9ro6EmlD7eLai8MSYqodq8J7iWO
RqurrCXUMim1GNrC8HHUSZJ1JILzbseX92s3UFS1oXqPM3RxKEVDjmCbhNUDshaXjhvRezPNejTO
ZXa2ZY0P0ShBooWj48K0vY04/Glb1lMQj9Vi6ya78yJyR6zHx/apF5DEAQskGuYvpFncKpR4M+95
PIl3pvBNnyC0Q5/F9bOig2HV7xDToTQ407PRacWJ6w38KuONIKXMMwQtzhTw3qZQ76Q8s5robhDM
kbCBwZHcDMwnHC5asYSgKVswfTMrzyVL/8D6VmvuCwellrbRLP6E1sd5e5QmpwZKV3ruYtwrLeCc
pDKp/qpXaihADt7FCQe1kfgw5yT4I0pR8z8lEECzslPFN02ETc8wLqSgKPqhBtywFWXCgBBP6Wys
UygwffxHQMtPK55BnJ1MFXh/Dn0iOdsJWZOtp57BJL2rb2Efaojeyc2hzxeSUOXbGr9yRJWQAxmq
rorP6/5ps31rWEAOfVVmMPyHYB7YLw7vqRCD9MEaVGL/acp2NcnNlPFqD1Cg02VQmgM31MS70anf
3kshL61N9Dm8dE93ur0XGCTBPrsUO0tpbyLfomnrZEnQXL3ruyfgHZWlF9p5lwsJiT2S+D2rXKlP
YuSLhhQRzRcGBp7V+MWMc1BI0eRCmcdxBfOBDJFbYNFGdmqJpj75dDP0pGaiQY/pegfJ4/0AiEOh
jLCemTOG/NUcA2D32YMAfcEWmqPrKbQ301fV6xZCI+O6W+LZrSrdUldUBmnNknw+OtfBCEVVuHC1
V+vX9EYBk3haHIBBY78HbFz5IR8ehT9wYOCBs9LuibWXEaMflTY5pNiyo7HrYNOq0ewoqgFpzoj1
1IzCa0wNsOIriVNn4Y5oJ+l0JC4aoyEXwKj8PpgO3jlYAt8zam7ne0hDCRv0fkyqC2qeGLwH9CUO
HQwhvpLAUYePNLGZeX0W++xUHch9tnQ/L7LT8b+wqPXnFabN2vo4D4yrIfriV0XvwObWPbVa8Hlj
Qn7mYhMziZw6XK8iakzZNXVDNynd4g/wD9iNW8s9plf0qO/Q9hFjVbNOyuvrad7a22vBml/9FrW9
mE3TToSzpQNZXSvLO/8QP0XDJqxQlgx82S0yQ/rNik1glwKmp0JPqmOHZA/Cuqug5M9GOG/Ta7BI
QK16TzV0JmpAUYxXZJuOdebuSJJCX4lUkavHnmqTGDKJM8eXF2neaXBwV8j1JaNtV5GxSj+RQDmD
tHde3xnC4yNFj+t7bnIh219kiN07qqgLNhf0Eo4h86Nthe3FFkgCHANAG0Z4UOx6NRlnBv6qt2iN
7N/GbplpQ3guWaqWiKNXchoTvjXY6by8+91VNUu1K4fGY77/MRioyzw9hsHQLEppTSMZ5H285j70
vgzFkWGiZfypCazChQOiOCYap/KynETP1fRIHPy+ApG/uraVjwMXdy6SYyhM8d53pKPa33DrQGp0
rY2pnkPyKXnGa2yxbWRhtdM4bLt7tXOzYrfZEiw/4+5qCGLZDhaQ9r4XNfz6HmJzhFxlk60FCzVX
LbalUiOyu3hN5Hg4SuwX8jUdilIwnkkZygacQl8OqkgHXFLqKk/SORs48n6Vy7hka6zNfCTj57Ru
51/oqkN7wJ1hxocS664AgqQnTv28XrGnH2X1vuRzKUN2WKZOAyfTLMs1KhFjyn6Bpxx05FAP4cTw
z344sLxLh3bG8b1cIKyXdCcGsdtd6B4U1pt4v0i94DUZotDlSzaNjRVQhG6idybQ4ccSuqOUsd8j
dhMxsFFM8E/j+gGbMKLtAaQ4I6vV+gOax1g1+KnBVOFeTVWwrjd2rhDwoUjNlrIDdGJAymOlOOo9
k1zioM08go2RC1nXab+XDYI4PTeYtbm6fInvuSGosoGWiXRoiGa89twT0ksObIzoH4q+yZzr/QJi
wn2IA+msDkin05NAxcobkZToyuvXBkfXScTtVfUnVKhOFTNXmw8RGIawG/BciB6MlkN2fQkFwj3P
IjlKalMHgqi6j0wrwdHTcHv/X8uBD3y5EUSX8lKtWuC28pxS8cLOwCdhsf1jNpcYc39eysYSOLMc
xqkPPxzqR0QtsDvlCN6gI4VsTwYUgH9tVqjJT4DGJNUBPW/cFAmzsEq0rVTM4nhFFD2vnRxsILdV
l9EZS5xdYHELDrSz3Is3aB1NQw5fdNqWFAsvTdZpq46gSvk+W7W21zoGQLefFigei8A0rA/cQfoy
Hx/dPvR8zWUIQKseV5nxCijY8qwJuTnN2KcWgjGhgkNMw/guPh0xy9tayd9aRpa19X00AIK5aYLo
PNu18szMaoypwfE1pWisTNuuUMJwIPm/CGnsUKRh7IAwbkRRu+uCkf+VJ8DigbvlKiVFgw44BVsk
jve7hAC83olJ9E5rLxBSZZLcRFBzuUAemCCbiOL9Hd4UnB97d/9rQ+ojJFPucT7ZWVls3VspxR7j
uvzKxxO6obmqes6t3VByfZf0IEX8+O+tDL5Bh+lPoPcftz+2ABMpX5XYPXeyj85uDZy7xZi/RyhC
p9Iyekt0biM97plFrfZKYICBLl+AoNjyyYB8CykznNCflPjRL9woHpkIyIHQKoxbnFOwb9JGmeGF
rnt4Q76UE6JbB+XHQnF++selXBhO43As9IE+CodX2yBFkYx5kngqKtL4pFfV39FaDRAslQ7guByn
okk33XnZnuV5xp4Bn0iXzeYlwXKHSi920C3ru0wpDxOPyuHnZQUAGttNYs7mSGh5lW/60EhI4xHf
ciNAxZT1UVRd7yya+Pk2Pczr01GiBFJntv0jftMRw/hwXJlPL2+eHiX4YlYcw6ygr0J9552c6TDt
LR1mZ723+gyo9+L/PJG+YUnXxfoE1aJeep6w/nRYoE+TMnuSh1oNTA68DdAjfQmW5+ztmNXZdA+5
JxA7XO09EkcBr9ZE1ay+dLsYn4Kw4K3UfdwpHW9GFHLiRBZgL4o3lYEapL+Kx0iBAPFXSIAgT2CP
EB4h4/QNpXJe4hp81VA+MIpyPxHWVV+BW4zVJiQ/I8EiHTvru1rO0c51VWSu4nba4rnIpLlJTRJb
qGIynnK6IoO84/KibnTtB/DoKthk6tfhgBe0Dbatzp8QyzIiHF8PEH2YLmK2EsYBc5RpwcwF56iy
i/bV5orD0BCR1u/po1LkdIY/wSXegaf1sdyLkXSVcuUc04CKmbQSVpx+8yYf5epf9yBfIQtRJAYa
jT5OHemsx4hpmOgdWvogU5ccMPW1fbLSLs8uU/rFGchlwB9GOCe1SeV+aylEyfOdLdb/SuLjPHkg
ySXK5nru4tGBCeWOlm7G3TXOoOqO/ytaWV4Q2+4JT5vxT8inuTFd0EtWvy8B/DKfkAAO3ehHVVCE
8yug/HKnaKTql6q6zhOxvV2LGskgGNAwwhCmhJz/vp1ErktVJoDDcTMUZc+7ifdclQB/O9og1ksi
4KTicngBKasTCab6+Uz1IWkI824cYezgREYfobTuEB0H4wVKFFWxApbb06hNwwiuV8F7dxihhGbE
bVgqmpmTh1xRyqvMjcqOR++lqhWYEkm21PrL3ea1by0LWthMQrbxprJAihBy+xvtuiOai/A5vdR/
3KFj+dm3AYCu0e8K9KXV+dElbjBAGCBTWsMV43EP5CqSAm03U8bImBBUFoGCYOcT0JEzwc2SFG44
KQh/WDR8awWo3AK5p45lYU/InsD9K6O7Seai1F2MQJGWBNewTquV+YS4fi+GBKQ1hpbGc7o8MZdA
H5tX5Yg4ojoDWGrQ2vxtoGxc/iN18MpiebHnvzAnI0VtOnKcMYnBi22A3bDqEZufs/1zUVm0bt+d
HJyw7uzOE3zlJo5ma8CFCEN53ZYAN6O9POqa447CHi6k0cywRGXdAorwM7Pgp0ZMCcjJ10MwIYIX
6//xm+e0ocT1kcBJfUvjB37q92VDgwPYlakK/FNle+A30r1nS/Ub9fU3JsOD24StD7De9EPxcm5m
Y6KUZjAB5ockfEpA1y8C1/2z5o/STvWoi2EJTPWIS6rrdxdnfi3RsqTJxRgjM3tu4ht+sN1I0na4
louLgb3ioqB/ZauR+39SCwdXP1nvo2v6PAf9t9PgFTuZ7HT8m/KfjfL1GH0rm1Y/q0Zo71nd0OW3
bx9sOjzifLlOVbqhabsTQdEAUg8ldFqjuKkGrj4xQyp4ImKa4bZLanmW5MrDPxzEwVRvUer1kZRW
iaR/3ZumUKAvFU0GJNTuZvdvpfqzwxvFk48z6iVj5P4S7Xh55ql4pOE1IIe5TV7SAW9ga16fH7BC
IMfU9KGwMOqNEpHcsWWsVMt2EpQUX+SKFZH6UXMxY/gG+8tSL7FDzGwJmBNa+Fl1ABejOFURmlNr
P0efilajespiWTGf9FEadYTldsXwkQtJbsbc5UCvMvNOCFdYq/h/t2YYCEtphXsp2f9ufnRGON2Q
eOwz126SG4eSjAjCafcyLNO+lP5sgBWtts6n7JwC5pUU1hrWgHQXd0cI4qnnCJwYk1pHHXIqjk1a
dmEFFK6R+g9VqmVFUR8l6d/AMFqz6l0w2sYVR5BwCWvjUjiPN1VOHK3h2wDPrgCfhxy5XEAd3KKK
/BhY3E1m+cHX6DuRxTg6MBWWglxruXJBpJeugktIa9530nuoO1Nki8g+meEr4UGDxMI6tj581bRb
mndTgIZIttazHl4qJllT80AaARmtllFCNui86N7GW9gtCFh7s1hTW7cDAB0RLSk2wGZqefZWslf3
TLYV2TQHqP2Bvg/e0NLMzL1FourJWY0/i3y4rxuN5Sn0UxxfufM+30wnbapWWM8YSlFbrxunBmbe
Rw6aD64b/IFEEfv1YXgDWfOW0pJm6DkDpra/QOcm07bOaKePyRd1PceVGMpymdqXPzKFmbZau/y7
vagJrjCsCzfE9EDQ5MKtsv3r9mcwfdKk+7OCQpMWJ4l72XZBnGfkvoYsGzDS6dl37vQoAY+j7XZL
DDSvEsXV/wbbdFY6NKCVRYjJj3vBo+kr72To74NDXfbYL6gLR6tLJ66bPs43N9sRqPQ5SeDlhugx
vc58DsOtQfHgOWVxOSIvsjpxRQDxGshN6AZhdE/ZrHoqoQG37BOCK4OVX0/RwFXbQ2QVVipAeuIP
O2+kQmon18okyi52y+JYsh63GxJFbIuHazESOPwUR2gBr3892rSKKpDhylQb717kdRwtKJLZcKzg
D3Vdtdm1JT5hZlc/aMuVY5vFlhBEsSQpywJQy+YrVZEYnuQyX4N4R8qyMXSHjJtfXumFKuo7L5da
l/+6a39XxtqUT+2O++/vueF3D36E4VHBbIxKYj+KLmpXepfEzcF5t5GXi75SKJXvDt/XxwCzlpM+
5psCHcwsuRMfKkyHNJvUkQOGr7Ihxp2q9iNe/DUC3PIJ3g03URpDlbgigEYT+9MQ1eIo+iMgMjcc
ZABP7Nkm06wsJ6mQ03pSC3GiOtLiikAmjPaBmtCdgnSAsSf7OkLa/i4WN4PS2LaBPq+mQ/dUaxKH
pqtp3qpXvwya3GU5LJ2UhwGfBiyamcfoIZdbOMAMR8XpOYpDojT/pQ947bMMe6HtmNHw2xepcRH9
WhI+jnJLCr1hAWFjLnP1V5wLKKMDdYSgs85shlgQkWlsZXQTuDJ1BS3ifa1BB05+9lpVR6IgEQIj
wSEBJfZNr2s9lL8bTW49CegirDZhIRuD8tflowsLskoHveeHjYCKekfPBu/MCQcsP/+9aJk3h69y
wXeDtUNhtDJhu84A9tPSof4qR/ghyCV3Lwly5wkAjSbUoUAmhYdb9yJl90PJZVL/2d8bFC60ld+3
FGR+rJ1jIUYDjQQusOa7SA4dS2EfBIA1aweB80Cye8N41v6r0v1pRROTJliRA/4l/GK1NtEVFujl
7rwZhJOK9UtXInyj+hBFuhRsWEtt8HZKfQ5py7rEwI7rZGk4MRHKCv++gRsugT05cY55rLorhkCJ
A1UWtjtBK656ytJq0wjqae+9y2QHn9AqCqKTfGwTwVUUNktDh2/M8XKAvBitLWOO9BG0HueqmzbM
Vff1vp+UzLp7V691VvfS/mBpf6q+08Laz/4TsbDGNfouU7r7cNveDTXy09oQLY6q4mYG/wkyhKm+
rVQMAOmCqV2BloSN08IJPi1Dpduyg/mifNBiKWuZDuDIH+mc/KrWpoiTFbHxHuCZCIUFodbzGnIz
R501P3LeRT33ThmyF2goHHoahC92HMVVHTijqyykNmCRGsO7wwWmGQdYzUyVdsXZPiX/TWB9lTnb
cMPRDyaf/tP1/Js0dharPH5yU4g81A/QTTe5vrScG3pFDHILdHsSnykddCctl8ZgNxSiUajLnwcA
Co56kR+V91RFa6I3F1FPQl2fFM3A1OJBJ+SAr5i5v56QnKTgefDQtxI9u5MjFWSUsyFSF6tBJWZc
ZXf7BozrGk0RzYBob5XuqF5E9qpgLln98P9HzGQhNYtcsBKp+aWQXxxe2uff64d8zPQREZlxI7vM
JjHiT4VSE3loSMAOMUELcJvCHfhpdclqAQ3rZDH3kRPmNpVGOAwyHiDjHHDkH+cS7znsbCENMJyF
oupxMM4/VbVh1JqVFvBA0XcyKXcegoAAbGzfp4+4RiGv85XBssqCyqtGaQV1X1+gOoNVkfe+FTFw
B328efNX0Saspi5hcEQnFXpqccsCcVM7EBukeHBEGFk2/YHDXdBZn7U8ma1w7OKpPTnBD0SmG41H
fCrfkmRoXtau78cOColrJUrf3FimzL2/fu5NSZ8oJwGmAtmqcSv8Yu/Xl+L8oN3/RxJn3jp9sIy2
J4wsiA+SwKqhQtT6+2dAeBFERGRy97l9UPS/dqJoafFTRAyTK4oOQDi4Wf1fn7r1cF9aCpo//aSo
Qr66VLLvR4mAZhDuNiGs8vxrSgwmu35uym5zV2oqYGvjmFlLLygqSkTxUWydxnzofgBWW5fg3vbu
LE9cLzE2EbYE8q8iPqWNHO6/IiVfr1lC61yYjhDLL1tJ83CWKeBrn1hSunlnj0Sfwscp+WYPTraT
lliMOYA0JPlPQAngv01I+357n1PXxlmSR8hJ7f6IdBXLpvbFz8Xa57+fs3cIrK7flTdypUbSI1vS
pxyElK9SomeyT4KIkIoUcLacoiT5tJPR+Cmp8WBDqgvU6LRlZW/erTmyr5X/FIdO9ZGt2lY6ufGJ
kQAw0Pzus+FZqK3as8XXzm0DvA833j3z66MWJZmfFKs4W9UiE9OK0z4gmEruvnkiuttV7pStb1+0
v09t5DaxtPQNb5PGImSPzEiVEKOIfUkrWISYYoiBV2Irw3+KEV7vPOasgXzc+9J6sC040iTCLERL
+d5V59bWZIPWKaj32GDOdXWQtJnQLLid50/9lYIObJ5BzHX8z3Z7O0j1J9Rkr8ibVItDKKbWLgdZ
NN+9+aPS6c+sYncihFmIyplujeEMSILL+QwlNAkt0FWBgMWZF+ZgvW9Xgl+zld90qYHfBMhWUXb4
0renaR0xL+tCSHFh7qqQ4MQjqAQ7q7OgtSvL2n95VxTcUG7k1r/TS9NQHwyLAWeynD1SaY58JAgt
LIoAzF6uLe9uMyITS6mn7r5S6AvcttToiuHK2aPtSirCaelkBJXfqkCwFmcxzhC+DynEs0HNgErr
KmUmk+pSR/Xm5rMxd9nzELhsiAtEeGpxL24R27YU4yl3ktfBV6p/AIlk7K+J7hMqmv2KUycgefLl
14qxV0DG+SptZJ6jN+zZ9Kg8kjDKsrewz+gMVRSWALR/6a9pp6pq4ebLEpPL1g+HZbGSB2pwWmN4
/7d9JepiDq0wWY16wKnpq0cn8T7IeSLm9c+daS6FpPy9Lb0wkFiEuPj07kkBsxj+7GwhKt2BtSHp
S7NfX0ICDD5KxFxloXxxmE+5desjb/F1l5XLPNgBZr+m81ZkxiLa8ck2mgtqC1sofch2P+pF8Lv6
9c3GiuJnevfbqQLXJfNQ9YlhVbfIavno3GxpgUMJvXf646ks/t19UJR7AgD6Cp8BF5OP+99qTOwC
A3W47LmKpTNE+bfg4gLGOr5H4jwjr0XCY3r7SZbUDF9w3m9sbIuq6wcxJLo5EYHLZRwZomhZuU8f
W69CFwQCp/dql/cd5DBcPUi5e9p778bsFK00/b6lGT0KtCGeIg0z+43CmcHXkJhqtpSO1dqSGKZN
Z+dBSJogUeVr7tUw/BRy/jT/v9MH4W7hB13SRcWx2z1ci39KEjhAE+kNxs2UWRWZeWs7DLrazr3W
MB6uyeEiJPr8lKvgA5MpvF20LDUTFLirQPEH+P3rnCBHWPxLlPGf2kDWu0aqphZHGfCC58prhsre
rpQE5YCPn7LrlCKpzmbPcmW22daOy32tre3OYBoq5qKfxmAggCoOGUx7vqYY1gUqns5d0VfE6RqA
bkdg3nps43BPAAU4g6m4OmK8Mz+6Lf4d+mwQjVz6IXkVQ5wAiGMC4WeSRjAB1geDHp5PeooG2DyT
oA38SansLYfbktJhcMTktizDjyNFWsWb5+HNoE0V5kbfbbgShbrdNJdoImzyaQGpZGWCqhEAz82m
jA/Pnp6oVnOqmLRj8fI+IEIzvwc8YYKoXXUfdINdlyBAr0E4zCn7f2lto5MKWmFuxFhtRqAStXwh
DPTKPHrf18VlvStdCZ0/xJ3Oi8g2GN4NqJNmyqLKYkPpmW2ZnK+V3exFMEnedldjRvSiKJHc+TNb
LElxmrt0+98q0wHsHbWu/Fej83Zqd3xMCxYo0yj282n5QI7qfT0bYYvory3zmuEzs3it86CyR9Fq
DjKXz9eHDjfehPvj9LlSR64BDih+2bp5+oTjA2Y986XCu80FMYQsuc51B5hLSS8MhK3+nLAo4dH9
FndlQISEgfH3f92+cX1HG+FRq6gtIzIcrgdKrqJlJ1rKUX2ncpcoeSaPPDHUresPKOyNX86sZebn
wSpU6i8VPp9GUYYKzlkW7AEv2fBpq2xlDfkcns5EtArKhdAb/XT/dsBl706aYW2fa0GzhFEo01HB
RbM9fLGPhq6IIc0pYMkjGz/M7d7/bkoXGJA14RTe7/gTvq28hcoXqecJgz0+8aPPZhNPRXEBhyfI
aWZIILjJDnlhY3hmaoG331vV0cMgZT/yODI4+IO4DNVWLoeTh37z9udsN/heBq+ZO2DCwy4136K8
xCYyPcLHdIGpJqw6DdH/mNws49ZgD9U4Recd5riIDXnyJfEWSGBhzkcRUNdXyANlvVVj5uKTDnTt
yQr9LG18TNUqT6o/I2Ru1L/TMnM6feeTiTPUD8BXqeeijbz4LKd5rQeYLOVwjNhzQhHBHNEkwjz+
qMGhnDe63/O0/Zdhcr3ovKgsENDz6JPbxrCHRY/Z8IVnDmZolpi0+3fhW0bWiMMQN0hZD1/qgjb0
Sd3xu6P8+2BV7B69DEq+mMw2BylNW+1I6Oh8l+DC2gBMksQcJMmSl+zQkA776izwXF8bm8SkMpjo
jBnJNHR4qNPF+4a6iZ/fK0YIdmqEKyfDDeJndw7j0tvLPHmUgyUg92YQmUeh1Iv//UAcWd66+YEy
Qo6qkcSvrK5WdVE2KmSp9kZd2VHbpvQbRtNiIl4iETSZZgrVF7k8pM5nBh/RVvHAZl/5BLxrDwjU
+y2V5/CXhxCL91Y9YJ2WO0AfNOrJiTThtF2TEIyuLvu/XgQK0+X8vCbCOlWP76boRYJfBW5Wcga8
goZ+DjywAbXIo70lEAnCU4XV9pFRS8/OvWfyPQFaJCjWULr0RFlCewHcLPhvdDh1h5PFW5T6jc+8
6Hz+a/WNc0SXON/R6vlMJfPuOfYAx4CahcoiRSp/+6cQ11eXzHqgwl3xBY70NFUVp2FfJLRjSEK2
kM50X51E8R6mj5IPrhgiyVBlHpGXSZK0CbHGRFZUwdRskFBaQ855LPucIh9kQ2pWnE/tuPZduPEQ
u64h7v85jl9haMtzDPXaoPkyON+ftYoR0+0jKNUNIDBVUkmAmn4daD2GUYKhlEGpI0oipjacb8ne
xiy/hpSxYVVJEvMYhg1F/9we1D/Ffxwk7NurMKtMTFzddCUo5ztKBI7aTjAsB969HQqOpq8pHpmk
vZyQX9WY9vC1o7ANTDahT1a0Ghdvy99VYWgPqT00fNWIE5heooMIvxUMKR6LjtCpjmTCtwQoZ4cl
G7yc99KIlmfwrYKzuImnZ5dvgvwCr086mip8+5GGou1VgoDoZnFfS4jdmVxZYpXkRLA+xObvWIdR
gbU0ptZpTS5Cx4/l9/qka5n01j59xSWXzWdF3d8eNWbakQw+f84Qw9I14oYQx1QfhycL+xcYv0rh
995++8vfeBdj/RN6fxw2fCTzaeKc8Xizn9Vg9rrO2yhOxUvA7P/PR+RJkOe6t2ppqyKbNvA6fvUD
XA7yUt9M7KrGJeDK3ddr39wzRFym1Oa6qyMe5jqseQlIQBk1YoC7dPv2KkQtmOWT+87sMAR7CW0W
mtbC6c0HRfaVNH6RuSDSu4TZhh8Ft3fyeFyGuTtn8Y4mthY7MY9kN+S7EQ8Ik0V6LhXgqrP8mtdF
BKV9NMcVSZsKTAlmvN1zvXP/wrDlN1bDEeMX3sFxK2ZPn+V3+LWIHX0BWX7WHqgKjei8E7RtaARF
xO3NRJLzih78LavSuUs/r6vEnKvy3/xK0ImYiNI01v2dC/trbM1v8RIIUpPADPGTXYnGzbae2SKj
oWkijqRWTAIKc4J17FHfGcm6X/FFYzJWXUbj7pz2f5sc+5u/zaa34w/CQ5zR7lMGr6NI3+W06ASC
SnqlQVnbX3vx8KaVGUw5xgORp3NIO3aM/mbFNDbz5IzKhgAWW0QvusGVmmjrgNEUZ5dAAGajJNCm
lYb/7uoYSEJW7xLessAUitwaaT0GL6OGaG6ZpVm+43tDxzsoI6PMc4KkkcvE3neUkfgTan6MEd6o
pBj6JzCTl6j7Im9StTabQBuetMU/vpL3fGomQo4RgMU9AUc8Yndh5zMK8jM6cXB2WQCbVL865+RM
JnwEBFEJULeQ71KrFrKUZh06LP2THgwyPYj1FG6gYyi9WUdi42gvYTvHmLa9sQd41dBYcTmCJfiA
dE464f5kt/Xs6bK7vO+QyjuoBdtxFytU7cDQ3FuJphpPg5jsJZU8BEInSwkK8Ajn+ABfXIYUxF6C
Vbel1fkeaiFVat7U7QGnnMYpSGw3D1q3Tf45dnlqwySSF4QGraE3Fbvqpfft8VdsPbQM86TQtqdn
lfYEXxWDWiSEAfCwU9f6IauEf+PzP/6VmNsP10ysAiSe/d1u9bKKNHic/VzKSX0QobLtqFwCEXRI
EbYI5EvA6WRcSTIVbm3vfkQ2mZ1m6GSZtQ0GPsL6tYByVr3XUOHjRGdNO98V3qDWbHg1zd4+zW6P
PZfakPDMAQbqengl2qhrQP6hl1Mu5ZmTeh0adLflA3vdcOQgxySf3zrtO2pMlSuffOlnU21WSZR4
x0Bp3uLqR05xn+dJrv2k1YHmt5SlVGDXRfVnISrBXErYPMkP/GYxN8FKodA6V3rUyt7OMabwkhDU
3IRSqJiwxhsy7zHRiHIVS5nGNUteDsC3MfWhWvqTHti3L6wWiDtrImewcv7daCi39SHv6TMkAGeq
xixdo+NHs8Pa6ZI6F1JAUi6SR0VeBvD2KLYhdc/4qytSdbTiLozTB5lz/Nv8XnSOsGhDMeUKZuV1
WwZCWzBWMChMeRh2pBUUF4V9VRY2eqBMT/kP2nwiIx4giA3+AVrbmT3mcMUawtVE8emb+NzQzv/I
jGpkFH67I81vAmvnArpQZbQU2o+fCG1/58qEYEwXfGNT5xgB0PROOqn9af+gUoo6lTj5X8GFlNy9
5whou2SZ8O4/E4yhfB35E6xGHpATsGcT+c0lTh+MQeAGLuZbdVW/l+0iwl5oDBPPuJl+sZ5rN++K
SIyH6fVMJTrJuNmZIwNnXEZVKqZnMQsOpOcDnGnWUu1mUDLVvkZBbp6srGTdWSE+f9iHRpI4RulQ
woOBpwWSqkzlHv5l0RZpChDsFQsUZcKwjPNmLshOJf7od7AuMRY0dfJ/HHE+xqMY2HJzvgsiWAQp
/UB6h0btQrhKXOxgfKCfysrMBOMInvpO0L3xmfQ9UN5MRgBmgrhRyGThRcblFAQfCb8P9mWEd7Q7
qBZB7MsWCG1u1Q9V0bQOnC6M+Xw33MunsJdGxj+t08NhxM7YC+ReyoygvFAjU4fat0gaxmjS+8D6
avqFntsr48sLX99rUbX5KrMCk+5lcJm8ddQQnHIN6e/A0DPl6Hvn0bjL3F7CJWrWhEu8XByUN/5f
39Fbs7CjlcQscw38d7a6zCsLeA+sCSYz2tPD6v682Pni56WIrdS79K2lBMTTEVwxixYWSjlqLqmh
qmMn7x8vvmifTr/CLZ0BhckylMmLIh+BPsbH2pURMUyMGMYHCiCU7g8iRJ4VhlPZmlNOitL97qKD
QCFW+crx9HKefi9XYYEzrcu+issA2PABBmzH2In1VIPMeYlHW4GHVCwlFeD/K4jLvHgUZSwjfLXI
6Yo83wmanbWED01G7zOZpsAjdnI7rlWD7btj/96re8eth5kuiOWn87VAlSBI+TyFTGnxHQy5Yond
Uuu5iB4Q/8CJt+qiDhgX/BOY40kaR6dmYYI4clNRYK2ibptnRsKmYG0a2NJcmPuIVwGT6Fg08ooB
SuKcTZZcCO8PtMIKKVBnsbFzsWNWqCwFGGhm57z+vhf25pYuwbkTUgUDitID3bDPSgepRjBBG4nw
p2DNoYL24wBfyAtvT4DhWkuR0hSMkeyep4naJfgjkBTgXyExDWCpp2BB7lh5dFICg0qevoLJpMhC
cq/aZA9+Iz0AwIDYoIwwuQIWO0dBSeuVWEAs/xE70z4CKc/SYRjTZOU05y1J+PyrWVrIK90zOGTW
En4TffIiSisj1rXRYp/pUYZWyUy2TQxoCbUiqvWGERNvlsxg0oq3E9UTeXgfRVilTxw0MAtX42Ib
mCUoU+rrky1Ivm3sz2ZNVAMCl2myDNYfmUlmPQIK+lvH8psqTMeOlr2TjUzOE6vtnveKN0XPY3aJ
P5yz6b9R3AJiQDkbB+sdtDKkE1+loycBPlVaadC5Fhpt7Llf9WAOxIpmqCiaHcqyYxIB1c/ELh70
YTqFLeoRggY6S4u7diy02A/1LRfG9id57uj6OZKBR0vbL74PgDKLrBU1wsTbV9z7IwABeT1ph31L
QwZxWAZ8VpRfhBMdzkdbzqn2RGmhYrguBzQ4K55LGGkM/EFKBdgD1ZtJM/XZUtCi9AnRlbCEL4qG
1oBpOS7XFBatjZkc37XmS9Zsg/Y6GZ3i++C4dFLF6m3JFozb/sDFmaC+1U6z75ZUqD1DPj6gQtOH
u6rudEueG9yucTQaqAZB5WoOdJfqWD0Fx7gFAjsAwck3ETSqxyRNXcOqXZnHQpWZIr00itOlHGet
Ug7hv2FKsGWBXSMAYQ+JhCtGurhlGE+LFFGGDp3ViYS8nb7dlkyMAfab9XVhPMwEdL0MoaGpvnpS
2ctNFXFV9dwjHHCO/DIAbVSsKdw/Z1Ab6lYgKiARwt3SvNwJAVi2xmi4ne7mgcm3drCHQn1fcpF+
YHjHNziyNhgnUDpuWGztkVk8xWMtHXM9TbAFlKeEpHdnPijPIfswGSkhuq5TI+OJdPTahQMnRaUK
x/NouooBL9gBnKLKsC0af3xmWu2ucQ3qpC4Jwyxfs2m0lho3YlOnfyv3tlWNtQnI+nYL7UaZ5hIr
GppXiFOMpiuwGHoBBQ2rzLEAUnlTrz4jAiBZwdDNPxfFXYqpZTPp2fYdZHRaIR5ap7giZR/JwZQC
cFbCJuVgaqlsf8pHSqMeVpgzzIXGmCIx0NVj2KjovlPlu1NDWG2D8W2Y9bAu4urwSlSfOZjCH6Q0
WGnxf+EDEtFL5vFGykmS0wy1cJNu/DL+gUesDr4J2Za0tqwlc2DteHRn7xBAMBC8moSfqz/tws/D
1Y/2x2NlNQeeu3nBA81Ne3xG3hDQXQL5huWspDt4sCuwYCep9cHLcSoXJd19X4yFPg7oF3m5GiJj
Efv7vyQXPH3jSmZsRFmIObQZb4q2K2PTzqptpdVpCPxKF17i/Q2v+XLWhHRXOcIEQxb5gWE1rHG7
+aY9kpSF/oSFaiszzdtJvk9dI+ebP3DYqJ/uALd/gdeunyOxNGF4+NHrWzcfzkwXTS/dcsNGsV/C
y8qkiI7j1IZ8NVZCfAzunj0WBvGl2XeLb+QnLT4csZ7blnReDQV1CQq0Yr1x+cHBkz1khJDN9DXd
es88kF6pDR/uQ2TZS7sxjcAcbB8iA8JXsCLWMevOOvQdbXGvg8sdsqksg176ckPgN8STKHeWyBoN
oQE+OUWmeh/IjFJAygmIyj4eBFAv1uX5r9dMPzQZyKmK1varEdAY4xVhHHgORWATM6dlMXYBcXGy
SJOnXwDfFyGioANl9ShHJ6m53Yxw4eX6BQzg0jo4Pi63UQ50o9vZgPUPLnBk86QjQ9P4AIJ2DOet
Vh0KBIjJOpiGBvgqA/4i1726STVDypswB+JbmoTPlTOYEg8vrwhjK0+XNzXoMs7z+rKMteThfy2j
HM2vZ69toWzidCiOHGIRvkvPLcSs2UDjTebw9PSHCKZUOsRnorcLqPn5nkaoAbPxVdFQDVnMgpxb
A9gPCjHhH7jd6yv5lsSL7wvETjIVE9D2jMMn6bEln9v+doG5A+rGDMx5wu/TZIJpgf8JUPxxIzWB
FFCbmgPZu9+DohrA5RIY5pJKgkDv26IG+wdz3pLqXnd6HwZ8OO0LHSqwnsyxOYVnqF8yehwmATDD
nGFRAMfG+KrKlYLTMacbovxgVK2s5VGhI93tu3ww0/A5fcz9otfX5+ovB5oOpOsjvtA50IvaHlAY
/QUOUW3Ahyzr16sMNSlbpfBFyC4sWhaCXGBkgeZKjXNYyybjiOGRkiOdx1WDV/qOD+0/cIMFoFKE
RyOpxfTnNRIhbYE1ApOdUs3jfOF7S6FTo6bWPGMKrZ7Xzika2XLWMLOypFr8fergj5TY8Q11Or8l
GSHOlJdNOLbbzTv4zw1PAP3yQmsD0llwi9S9d/AKns+vJk2p+3l0BZVk2te8qzrnv7V/DVbNKHiL
MvOXCVGRCk9LlGunHUeQd80qxHhWOxkjMfiRXUzAtdGD6LkgOwaBp2vT+6KL+YyGzOT+Stfx/aaD
0a3TcqFymd8uLjHhH6ztq0XAK1UVJBLRcx3MNgnHa8stXmc8PD0KeKFvOF1i0qouKFMSJQn4hTfs
rHCKoGu1xmxjVtgzGNH4CsaobWTvT4YY2JQw7PXsWTpB95VjYO53pTF9XZW+bgPV5cPasmdsKmIa
e4b/eek2G4KJkEGAiiMA0KM3BO4t1TTkSVrV0to3H4PxvdpnlzRaz0pRniXo4HWHL0lwviIasA4R
y9yPimKjrSAKj+vWeIOA8VawmwPKbnj78AKSMsXFcQuoSEvCln3vTIeC7Fv/90ZegpQQbqO/CapY
GA77kg5VfppWNfA3ldERX2gkE4M7lQT8yJpIUTdAOfr7aSpi+YcA1Yb9tu5iDNR2rIvCu/rC/AOu
JMwzNtNM1zC2hqXTqhYiUiEvB9kIrfAdtTmO1t8QpyAdM/jdsoDbxLtC6JwD4N2OOpZfel+FAVYg
CByW1yEC3Hf3wvAt8LcndKwJdXmMoxEU3ER+pfGPwdHX0wE5gTqCeKDjCOKKJ7LN1IDSPn/hijHw
ojve1Zw02+7nyPkY77/a0LupYBM/5/gR3TNNyPfOUtV7uJ3Ll9hLgocEWTaJ3LrrrxJT3o8mII+H
n+tEVq6+34LPyqbQRhfaeyRL8f4TJyCGNrW9jaU5fIcB0iv3Gu38MGcBTqXLScOQh4EFGnQtTYVl
yNf48iZSHdYBj4G7KP6mGDJ+RysR6i0ZQ1GsJ3HiYe4SktYkLD/XSxsJIOyjDihlnmnNFAo0ZLU4
AXHDuJonmeWeEae3J2gpN1iiC8hQ3fSP4E0VbuxdvMoi2lc/Yo/DaJovtUg5RqDtg3sGXYOusskW
w4zzfBJyAHVh/JBRn6T5+iYrG9FvVG8zS6d7PQAVAipskJSwKoKnWi75N6b0z2QdhhcxLUB1UmKg
db7OD2i576lxm6e0qBiZl9m0M2vF5K9mziVqJ+OljRtoLzN65hCgUs1ios+D0pduz4XT2wY4oLXw
8HKKKmcwedLuJexlMLIMHrRvTkNnunwXehPil4kQ+yMaHTQBpP3ysX4c7CeYUCgnp7DtKG2TDmoY
waXXZP/ri/C1j7dcDUvic6Q/yJbm6QTWNFkj7+PgK3z2pAYAc6tayfMA0o+JnHGag/rCioveKsMr
i3Ijk0iCkabRWTegamKp/cxV/QUc6rsl/+eG9cGDTJd+WlR2SWw/cn4n3CvvLA2md/AWN2oLGUmB
NSUjNO+zdyOH/NifQ2L45p6AFU9Bcp1roqByX1riH6wBHa6diykfTfOp1qQimqdtQHT0kRhGdt6e
bQyBdBvQqOIvynorIQU5mH2Zi44RntiiVwSBIzWx1uGpN3inMQ+0/Ln64OgThMioRQAN/7gesHI/
0SXf45Yhhd4yH4BJbfUIli9g0E/2C48sWvynwx75UnSRzOr64FkbK5rZRwJ/ANVHXa7zavcxV0XI
5rl+3s8pSYSYBugC7sOQ68ztmVWhmiLPlNTjpjv+bGuV7+vYG5M2i1EJV2rVHpUxHSkHLf8vTbqv
GkFaLCOMvhdLzvG/vJKBfYU0UTTnNJF+b7b481VVOLqmnuMzFJLlVGNMoP4Kl2ikvg8ywp9cHP+y
4pUWzCNRMyJLHHzTaRMObfDXSuWWxv/ywo7c0sszM80MyJ6KatQ1HksK8LULmBt2CRnvmpVQdSO0
EZ1ppA9e2N1EU1cWbvwpDjU4C/2PyxUyPx5F7djkOSWeAIfNVpd0rbI1/MdYhoT/7ifx8H22vP1y
0C1m4dmJsEkBvxf7SRIYqavT3z5YxY8qWDWl8tQA4O30zIOCtUbxXMxjvxrcVtOHdZYFo4jVhVNP
G5qm+tojKjNod6mwZqPXENyIXAeqzXGT2KNpe0oFMeU/tya63TEgIw6DbEM9LbO6DjOHbiYpVCHN
OuXeDf51GfzCyFnr1jMVsHcs838bmwOQ9R0nRWyvUpW1YVM9u1sRqDzRAR8Wjkv1m6UdkAZvUPVM
zNHsMaOWr0+DTvrhwTyHmRHqgDC7Jc7H+WZvbZPwopGtOfNB4sg+q3nDG2Xr9YvXUuogw0ZadNY/
4jfSeWeXn0M8Z6DQ8za6Md71ToS3LkBxH/xbHC+ujxnL5Wo6ZMHFcUmQiCpS5+wXMb3S/FjsPQua
Mnne4pgBUPGGAhe+QLDpyCodlkf9SbD0eQej4bfcIwC5abRrKD44YptCxF4vGiOa7jj6aQkBdSKG
O2Ka9JsGiFZVYg2Xgv8fJl+25iwGAfqGFPYjT7aWESRLHGliR6XeEQHNAzonqJJV08jNXf/kurdG
Na2zl5g69tgeH4H4zzMhUP9macg9aTxg+hXKH3Hu9KngmzlF3asIuRbVoI2lT10u/hvZQ7vlSNrT
v9AyYarnVXPUkkMqfusaK8i5IkMQZ6hDUNO36sQ2cs7z+VXjrXpEHtpgPFY/MIyIN3hJsMQD2cgz
iDlVd/j9iHsvHSGCzKWOxBwK8+Cs5HgFIZxuehoUXRLVGZmycr5N4sQpWvcxp+RDhsAdEpXUTncB
fRFShNa47GalRxH5NoKY/kkv4qa1P5ntyCZyUva3Sf+zWG1olIWvOUGOW06zB56u762NLlRQDW6V
KdkxeQX+sehyZgYGSaVImGY4ZJr7t0IcnIaIdhMvSyLTtvqbRtmRB2kgBWnBijVRH2GgeV1/tVF7
OsNZsGnLkTQSF9rq3+oQF5UyktVlRr+Q427rjzrHUASVe2ewI481I9Z1u2yIzIEmtd3JqUl/wBUp
q7TWlDQLyw+JkmyshuKSh9DdLBTcSB0ahtlf4pIOm4w/qqgqbS3GN4E5tkG/IJQBxZZS6+IwADyt
/4gm0wAwo76vQ9qOcpsCOySOEKNdNhzJ/uIFP/fyKT+TdnGC+I2ljYAykHv/IZMmq22Txf+UtiBH
IA0xaDR07dFa492Abh5BaIHuVozUGCajF9DVWJO8DJfG3Wri39WeyJq+p4mXW44ixsPhnIWQsg0M
RsMo71ylFzS9gQVQdGYMhaRnYyUVbT6cB5vdCG9FNsqQC0jTyEvWmTjJX32JJY83XXjR/EqYqqZp
AgG1Ftwvd/GRQk1vSF3kpvUDKt2SJhMHbn/Mlr6ES0APKVIv30qX4lUi4bqlM83LykFQXb2DfQ/n
dAWGLwCbMdguX/LdBQNrXeSQHmPlMRyEDFHX79/g7//y+cKq/ORYikYkilJtxhSV48/qJqvDOPGV
xeFpgNuWs863WW7XSORoTMxhfbMrw4n2N89OWOxOy2E4L71R8uuIjpq+tQ3km5bo5Ul0dDiS71RG
bfAdmqf2CUJdTzmiIqHCf20+QCqN2gB1mZol9TlK8OKXUZoTGyKkm5Qru8pmXYjz7tkyC0yYWNOc
y+Wz75QVmOIZhz8EYge1aJIxqHsRq8zpdRjDzjEZoqQFvwE3benI5pe0YNq5gVjAuea8qgp7djwX
Bfkw7I1weLV23wOK7+iH0WkDB/lvykcBOyd4X2qrksZTDRU9BVZ7kvV2DXu3D84xsNZkLVu6s0yg
uyoXiKs4glJ8BCY243xk6sIvZXCIjIasub/SMEindiQyRJl2JaAkjQr6WuyOzWVcARjbPNEGCCC6
3GKfIeDMqNZSZfHHyg/fk5X2VtvSHtCfN/3bbe7JFTOUAq4qGg39K2zclfY8X51VRmoeao/7ide6
L09El6dB3crHatNct7opyoeOXUNByNb9PYgQq7qdvuj9vUnu3CniQz361O7QVl5FGa4kOM+zZ77F
Kf67fbgRD1lqX7mRGFeP52x4Qp0bo588xVqgtjEjB18GZ6YFk2bZne7gVLGwZ+1bJlWE42Sw8lk7
RJzmPeW244QXbnL3kzyA9yCMJsD3nsbyPHOgNL7JO6qqC6EtPbdL4FOnA/sbfC2Y92L9LzgUc1+V
9Q3HCVNKvGCJQ3vmq72XfanNdkwiBFe4FbjiCDczPWLRzU2nHBtiNjcbukut03jhUflhY0bWJo9D
yG/gkllQ0Hhaq/4bStI07ZLflxDWFv2lJjgmcK6Zo9pT9bcN8pxpmII0GkheTrSs/h1KqlDi0bXB
ornwY61YLB2TlVPsLR1mEAv7g9OlN4DhxcW/EY/ZQfbx6YVTadU1zQ/QllIezCj2k1XV9xxVCAIc
9G+qdvVBtR5ez3/igvGOka8iSxdjWTBQxwt6x+0cjOgVFlXASdCFrsq5E8ApQQywF0oerX96XWeR
t3y8FcsEbVOK8S3fSpItduf7FUW4OKTYFf+lFtX6yBZw18KgvPyMBk+xdIJFR0AyDGkKCRfCnF9d
cqoFIRtrqOHyQ3O/ar55QKm7SbnxmmA3HqLayolb+/ppGt5gGjxRl5lZvqWXQMIeMqPvQr0QSOt/
d3kldXnwjg8uAQWroeKmw/ztHZ21qu+BG8oQ31QFrXA0ywjeoFDjm7CXs23hmKalcpQcu6Q8p8s3
cqKvVRolJKgKP6C6rXXjCpvBZRWRhkoKh6hNJxSEbkGnpMcbF/t7Uk8EwEfm5NcoFNrhAh9g3kHq
8lkFt29PHjqm55LPs1sFabfrj++mqvCYFJn6m4K2XRVXhKK+G97TPkLPu/5jwPYaTstn1sloLDvN
iBYa3FjhhPAM+wcImVdaMBx749k6RXtJnPI3lV7QYvBy0RfUAyiZ7lDiptSkwUkFz4VmWHWt50gG
GQd4pe8i4WGHhnsVP3RYoFcSC4aa/gqS8cdAY3CGaWBKE3w3SEdTadlFOeaEUPl/Udyfu8yzdUFD
mJ3Nsw0FPFzn4SxxGiusW7XqKJXK6y05tSmtBAl+/zmAeRHxxNi/ktimL1Ul1ks3a/9Q7Z9tzNSO
dM8phmi+EUYF85difcSlhew0QwcKooudmDoxeEvSQ9ee/W4Ftg0DG+3igHQ9cyTypBywPyarOwko
SJYjaiLCsvqWD5z6igE+rH7JaEkU0E926pISeyFp+8vL2+tKwDeS1kAvRpQxqqXAfxm5rdcUdWcU
iILeANBl4NSL3ggnwRE+oJ5948OcZmDtMhqndfIITCIUT6ifoJ4oaDRVpuqpFjVib2/jp7+dznp7
fsyKlemiOMgWSeP82CP33u2sTcaSJ5NyeWTcs29lRZuJ5M2xC/zZb1y9ozcwKhAl7bPcBCZrgWhX
RIznXZkALX42STaawRUcrYtCSCYAgBbISC0u1KHALPJcIqp1HOacK7RsA11zO7BPz1yK7nIsezhg
EnU0d5Pu01d07MvWzbqZDXEMocg99cURk2Ju2WTT1yGwNnECh3ZE/BsuG+ypokrYsvRZ01kQ+prB
Ww3jv2MVFE25In8V7N2xA7xWNW3J+3crZD1EQKiT4sW4f1r6d1DH++RALpDdHjZCXZseFsbODd1x
xyEKcGtVhEyR0x8Ad5OuxnhEb6VfCZEbatqMkSDuV/10QA5k6OOz98nZjhLnRtk8Cs30eyw2T288
Zk2CmEMdxReedE/AgQ2pCH0bNZFl5hWl5RVFTDr6XIwEOg1R5e7SdBzKnwfVXUcktHOZ2nZ+Imn/
sbo9kGmLeBExT5KzMoQ+damS24vkIHDl37e2Z+6UHfDh5YA7vUlBEyxd98zC8UCO030z4TnvM9t9
GJG6xyeDcyvn/IZ2NSUSkFz8e/eiWRRjxfAHamkTjacOy/KZlCeJsYLMN2dy2u69AbRTVbwhVyY8
6ega7/m7FIBmlAsVrHf/l0R1yBOMhBOLuqnyDR9yB25znMcmIiUgIOf3WO7kukiPw5lQETVveqLZ
6R2Lx5Mwj3G0U9bWttE31oLkodujnIHz2pkoTgjTCGe6y8zOUcebUDfn2xnz1Nyj+B2ljix0ROx3
d4TK2LpZpCg+FiMygIeYS9pMo4cKimC4Jp/50f7PYtdyJxYQ2TIjcqz3mbGptEag26cxXPTmwwLM
b16KSnWWmbb7Y9yzY73zxBlODGSa2FMcZ3xaC1C2yCD8D56hPZDe1w4LZFLzgQH7I3q9S3vfgw3E
uat6cYKs2/I7/axloJITM90gOvOSYjvkjqAm+zYwGEN6STAHglTY2Rxw2zmUOG2sKQgnGJHbM4Uc
81/uaa8W3cJG8PO74U6oFy1/xzb7pVDeUyKiCk2FfFgkO5CxbohZ/Efj95ImgwpcSATMwZ+R6CFo
IayhVLnyCEttLFdWIuqI8TsvYbhntvLaEgpRAwmRuOfyaZmsHJROi9V7By+pQ+tHz8QosCpLNqYe
Fvp7ESH2pBRmGc19dOiXL0qXT2zYmYCoy/Uubg0hJffjG8QuE+bk8JT3JOil5vMZjAlksOi/+VAW
h1PN+zcfaI7yNAGWNs2zhd0PmFQ18gnEGzL7i9w6oVvfo7QR264ecfDgr+wAPnhq93GTHmSOItzV
dJzVyLj73Ckzk66WOzZXAq5qz3loTCaIR+sECpCrrevhObmtahxgALj3tJqVn2WuO1zcD83yg0lz
oOSsb36aEqszlbVU6XaBnDb+kuLHjZ9JHSabcUO6KXGF4MRRZFkrMSRvrCfcnvoYC0quwCo8RUAU
9KaErjTc/mPwt2n2XHXP7klHsvWyvjtRJIu8w1VJ85klYuKELa8H2b+qQR+zjYBVXj0zcGqjjeF3
MJ5UvOXrvEU5nZwJ3VYPjklZg/0qWGIDaKG6wRFkbJkpm5Fb2rdjycwyVExEe7CCsh1w+6/OW/zP
HlesVmJo3ttj8Z9XZQknMb3+I9cZ13U6in2lSIfp0xY1/zEBYe+ajQwr8wybVMOEyql37cnC/GWE
657YwY/m9gnADYy2vcD8xSgx4xkKM+er/bdiicruvjTrL0sB/oGw5deycPfttKaFJWXThGBvApyB
LD/k/0hHliJPLdyoSMFUojdafUcUZBEfbBdggOfS8up3u/hkbyQhrj7l4gCHFXWDmJJTHleNpV/f
PVPnkKs7ZqKBuWL8qA5q50fxAjHT9zd4qlJac5NrKEEWlfzloJYxo6/Kt28/fuuN1bcAYH/bhRBW
XeWTGhRDsUuxjQo1L9QmA3DL56tNWAAa//YLIo7wGq1WJactbw/eQAErCI/NpJztFnIqbj2BiP2Z
8HWB1THU9oIsO59VO+ybLGW2aXUQjYZf9vW+8wStKPIR69fWrAjh7+wATEx5PXOO4mxTiBbSAvNx
CVWaPJOCav97X01raeunKoM/MUwQ5QYiaaswxkZu6RqvOuY0PM+7v6F41QRUqFFMNZRlKDkC3dU0
xM57FJyvzJACJCfl51QQ8LehqAJw8AkjG0Zf855GIkQrxsPJ24e70jEpTn/U+DYX79fnRxUALDsg
Pt25FJ0joTzmic3a93SZ6uEzzR+0PgibME6Q1sK8S4mWo1buHsQE3SZJguRi1RUrXufYSBX5a8LT
KfrmS1eeQH/a+pX2UXEuGQoJby2wUVTjCP27aV2OGLk1JgG77R40zjd/SwV/HyW3NpiKs+B9xyxt
oZ9/+jkG3gnH5Zf0TWgtyC2ruUCNptKv+wd6cXEwdW2MdtoDVjY/itfSYZGXoARDysS9XyNG3Kg/
XSC2IVxOb7Iy0p0JPtVAVt/8kyG2f1aK6Wz9neK1aicROQM10yOhIZ7eMXHaJjqxvMjx65lyDl0h
7frufaJwSew+mdf9iV7uVu/2uhtyDihFLyfTn5XmazqX3b87wM1VP2ryBrkDroO+vfUXFknhr5dj
JfkUqT9tDrl1l96+ePjLWVkA6ZB7ytCcOqF8cT40Eap3eSrmyiZLZMicJgcATqy5FeTMnak40My7
RGyR0c9cOUyZLFW2smYCLP/vUBMiX6DES1M5hWRfeRIEabwwnvlDWGB3jLylLwofRr7p4nGCpN+Y
Ds8E3QeX2oAImjQBTj9hwV19JbwAp3j73hR7mVYC8W4+05cHwqKVjL5STrl3HoK8zJ3R5VdX0W1K
Vzd1Q1HZzOMq7HYR53DLCnYE7WiqS+AXNtST3ebOdt0uCkAokq2c6ZwgvXMfiDwzPNu9+C0JB0W+
GLxIHLr/Po+goigOY93iWHQnf675+yPOQ/kpRYYESepR63Wwh/+HRTx9sysHBdS4a1h0iGZz8wVo
leYAaTN7eEmifoeOJK9QhKdQvTENz+dX49pUHb4jzjmvyXxFBIZS/B2iFa5f2kOz8xDdxvk1Qp0r
nDs4eXG8SuajQcfR4BUxp7bnKZXj1fQC3qcvM3iWqhcjkc6kUx6eCmhJ4cmpZRp4tIkOmvktoREH
q04poinjXC78/u4bd4hCzX06P2H3rwnqpLLcmEnITUFuRrNiGY4zFOAvK3Lzh/SOavvikBnFHCAS
G1Sta36P7ST5YR/DFp/+9DOO+ofcuIvFeqJ+VdOsXSQJNE6mdPS5MfgxBcnHpcmAwwu2xn2l2Qoj
1nJcYs+VKyhyOhIocPYwSxZmP7NibTSwP5kpEkMkqZlu4LTyVhlYPXGQ5uj8yylylmqIHcMpqaDd
ttnMaDe2tVahcdczAM21iy8K0k2jCZBKknJLjTslS4iNM1dofhwrHtZxL0wm/1jGwr7y171IbLHX
VoUGE8YcpzTcGXdLamx9m/II6shSJeBGiT5VLHnzjDcrLAeHVSAMGw0tRYNEK6fe10TCGSlWzOTL
c9Rv/GNbCHUWHncwZ+yWGmy3vyXm9MFEf4/ckiMJ1gxFGNJvIkpL7x3MwP4spdgM4jkB3Czgikhq
bDjUuZiWB026VcftnOoxfZjrtZI3c0K/lbbHZVsIfLF0JtdPVu6cfuF4zLFxE/sK5YWPf+M+p6zp
i6NCYr6CPY7TQ/lTHUNEAwV887Hv97QY38RMV+3pA64mzI/QMVLJM2rQDD3dPq0v22c4h8poIUtb
bVwCLLXZTJcLTSViHEZ2OPyfv7B92GKPEVWBxdf8VCWpPtbgzdv7GMV8VhGO5pnHUVcWctNmkX7c
DYzWIwM9FNsf3np8Xc+vxH5Y/qSHyNsiFZRQ5HReQg6OO1TlKYyd9OKcanTRscqfHiuJMoh/WpDN
qt2XBSAux6ZK5q1tmUyvJJJ5k81THV1rWa0X+Zd6G4tTkQUA31RJY+LqJRlEnnl7Re7mZ4hLAnyx
RBv9Vu2boL1PNncPQ5PekW/FQoRPaRyrmVSeS1qWSE2O8mcwrcVy/nvDmANf4ZlaeMDpVX+EM5dl
xBZavPPz2sIYZL419iar5da/jO0q+ygOViJk7XVLGXz9gljcrf4LKiSBMNxbAX4fFxnFrXwD3H/P
KpMD5QwKyctb0KMRdu9a4wdOD2Ty6D4Ljt33xHc1iv+ocvuR6oXkhaPTpZrzdX/D+4x8fXniGWXZ
qzZj2WDjZtOccg6eOUQun/IG1M5Q4sjKsDGRd8nT+ANfGHdiwqj5UtifDOiR0cP0/oOSV7PjIcS+
Cl0UJrEHajzNXOWlY5JuqIOFLD4H0Y+ebQg3uu6uLQVTPz3yqz63MHCq/jKPqKDBZ7HV/yrCelwD
pZaaMcnIqSlNzADnjlP9q0djEQFNRZCkwPAHa1zrZTf2yp6tgitDt3+sJHsSvH7P8x6xXlgyOtCY
5ZJQu7K04aDJ+mGNpYbr0YkoOCbGraJFlPREzttL8HfRKic0wnb5PvbXT+wCgqWVgAhbypnZ7QKx
SZZHk3dAJCYscML3cutkWXNUnqejhPptTWb38mHRoIuqi1FNyPI8I8QtLGcRpo7Db+CPyRDaMMoT
uCTY6ykNzYtdsVgiHdZSQRUePKTb3Ngk72Mjvl6Ze01OXGjuuO2sxn4fOiC6LoCjxbmI9hSbYcB7
9JbtfvJbsqHcIkD+XysYuhnAPNXcI+97D1azWU6m+bRbQG2RJMNC/x253qeZMvKk+VUoTxwyrnv9
Ev0ZhZK1cCpIxozBgE0ptM4ekkQSkUF59/J1a1gyXWVrMmx6nVFosVNfNmHKCkhjcF7UzbZH3EFE
U/Jq7cbhmQYWpwkegbBqB+QMONYoUUDNxikuDRF36mlZC8HwHBrIbWVh1OK+vdMypB75T3Cy8BQ+
x4AYD9/lW0F5E6AfENCPfXfQeCBVE/GySkOH+h2nJtRdceYNM7tuZ9DcfzJuN8F0nXITSJAdPpL7
JkKcKYvtFV18pSRtK4TUeQa9DSKNYRFAkGbQbZFRzKqUpBprVMtxcD6NfGqMbVE1P0O43hFiU49n
PM+DFDqtIojY/pYtXipgs7VBuNFJkUK6+tI4lxx3pMOo+uWzrGOUet35DcTYOhfPJnL5225BNa86
e3mS1bXUK4nWgVXM9cS/WzrFy5t63eyjEGwDwybAROJoaOQAzIV4QSLXdUjTx8jHSWR6WnhYUOoN
hSMXDp1c1x6MllUiL2WFt7AQyLr4+P4j54hLrtNrJhX8/YSNkGdXYzb/iACISXuBE1OzO/F9Rhgr
R6gExgonQNCx4A2o5WvyPFBIj6qMVEU/7ajJr2AHKTf5BIU+JP9JJqqVfpZYVnH6g2vMoNk2nQnb
YbuF7yEhIdf8rxYFLbqPLB5L2Mhm8myrjq6eFO+QYga6wxGV7jv5WpNKImd/Yki8ZPaaIxAMXmh4
gG7y3BSr6yew47fHUS6GmRtzeubNIG+SXlHVeSCHWhf8Aca1021g4pIE55N5NrIShRaW4FaRX6lk
K3jIoJ7WWZEaYxHu4VhFovkahshUU4tVT1kRLatYn0MJj49UK3P5dyy6vZgDklt6DTXqe2S7ZsfG
ggT++4XqOMTpbhSMfBShKS79m2bYGCiwXkmZ74hs6heUEDgDkum6y0f/6SbY24NUpQuhHnWufqin
OwDiKuO5pqnFkPwbmYzl6wrbCLkhvR/YM3gqGUJURxIA/P8ZP2xeTVrkIkaQqm782L2gL0A8BBnS
CRU6QCnwOPrV2bwYjyMK2Sx48DpcfINhiTX6VInXLQVrC5WOWNz6Z4rtGvjxHDVj+Fi7+aXMneC8
WU49v3d1/pYSX4kOzcVlJRq1ybuomN4J23rDrV4yOqwbLIGt6P+UGLO8Yo3jb3VZsZbXlHGLzSy2
Gkot9uIpfQ1nOXqM8FDR5fmsjEk/sOtKkwZ6hc01tg0iY3jUeG6uU/MJj3NetWPInsCgoeapEjKV
eW1JDDZLqjNJRr1O+T5I65K78C/OtKDaMjo2Kw7NGOvxplmtvJ/92x+RtB+n66div/bqmhF+qQKb
VgAHSk+e/+q1YOer+Ug7YJl0kqM9bB78OMQY+F6Q7QazNac39t/FS8r+o62hbQp2ZZ4y6Opn5QK0
B2KJUWtL+x+tfvUMOIE95k+zV3jxA/48U5RS5GOpSk7cmg4EUthleXDsS8JmTC1no7jCB1PmN/1h
mriStIi7H903WbmBpCvlfNbTTYCBnA/VwttODxcHW2gFVv1ReldV3ao9QAba21zmh0dmknqeBn+L
wHxOQFrXqNDBUg4Q0wxqyBA34feiIxY2pJ1xkxj0DJxK3YdBpTjxOhZ+uC0CdnxoZtjkjtNYKEB5
3QNrZhv32hc0llWI3mGkxPpcsEuAHOv5Pvk7h6zz51gHJ9RNsuEZJN3J52c9iujemtRlw+KcBqfp
C0kVVj0uPAuBixQvw5r/mjCh0HGrk0Pdpll4q3eORhaw2VgLXADylz4T9zazvJpa7hF8wucai4io
xotIVLjk73OSrOmgI/lr7jomrSMZNXp3+02GUNVzfqL4z5mgyuvCu7KXsUjrDCkXlKFfebT/gUpv
k936eJrl4ne05J/wCePCaMGnm6z/k0s9WXSfLTwQEwCDcTqMgs9yz8t3qxQtyPnZ5o5dOmD7JBxc
rk+JmB/vNRIl4yjFWrQh8qtNAf2yy6Wnm4RwcVaSmnJA4l/iLg2C0qSCU0KVmUDNiHbhVOrLMy5p
j3j/TulvhvPSHxpQg98q+KTEcNBpDmHsREAqSgwU5KZZxBnKdq9qdu37BLFXdAqsJwejg85NV1i4
AxuAuAsmWm2r8X6Pb5mgBEQTZif5hNtLBihSY9iIshrrBa2nZNFCQyL3pNQ15ANVZZ7+fcTWEhO0
u0uvH05YqS1mgFi+7DbI4uNAmBW7+WFk6kNTw6AVEAD0vOZVxxA/CIQTdpID+eTG5uyX1svAiGmJ
lgeWF6ofMZAMLwxGqmV+x+nKWyUgzFA6a+z+QxblY8oqnJrJbCzy2nnpCTff+GJKe7PAw4Y7jcEl
LqxzPOag01je37+R2pgz78UQqJnr7Gqm5qJ7+gDkEssKNkUva/yL+2hZIIcGcE7xe263+gId6geB
8e9THeGvQx1EtPjVuklmEOYcKwF+OndAcVucEsUhnqXd2sNtj5xQCjGxVyGZrxM8QKuDaQnkz9q1
1Y78XpCuZZzkET34ZOfwEX+SnX/rzG1pQ+pjIIaKQTJ6X7z3jedWazPSjHox4q2Y7xsi0GfUGPqf
KV6AfSQIf89fiBME28qxE2OBjzF4u74LO7T4HdugCTEOOrLc4yiMLzR1HnryI4X2xV73zqXqq3uW
o0urNMkReUYCAIeY9lOlY2rrXt38pR0pHG40T63ALwQ1tUkgb5hihIdaMFdl620xz+VuVGG5BAEh
m7MKRH6zjvz8xo0g9V8tJyuj5G0dL61MfLJdhvaHfnB8xGxLPwtSdZyeLeKls0mMnhh+kxI3Sbdd
RkQ/1VWO0hg1ouHBQnTiQaMiwnD6fesAVLEXGUl/n1grls3FUBpAKh8GWpWRMzEJ1rPreRtyjFx2
ibJKPtmZxeOQeSQuCrwSr1Oq1+2IeIAP0hgVkZmDCJSs+uTeIlDCsKVN7miBQ4v4R2qMEtoJ/3we
oxj48lqDFALeZRnCnvn59Xh8ewVFIj/Y3OT+p7PbOiuAjBe3EG1BwS1KvYlusWcmYA5iLq0RrXj2
RhDaCZv/mOVNAHhTDiU+Vu/6nsNB400ytbQZpm9h2eXkyGMAj4LmgGyNV7s2d3pIwXg4Oj3M4mqq
4nPBI4NH1b7uEd3/YHNeW6xPtNFDhPNCAdgrn1yfMNW1VR6KSFk2FxWE7T3iAhW1Vq1y/dH5Mohy
0/DKirg27wRv49yWn7Ym6qCZFVPw2/ISs+I/qhcqLsBsQ1cCmzTBXJyJXiSx663k/9CjdtvEfPvo
pnlFcPQwG8jedtYVH7CEnRpQEHKAngS5J1bBK+v4JhQTAXeXqacn/L4FTFDwXZbslYf26Zqg9Qcd
Xp6pa41wlEODiQSttoLwFISoKuPaVQQG/jS2O7HwzlXYtQ0uCEMKGM7tycNPCZ3vnXNJ0FY8Usnm
xWede7ZpQ2YYgJyxn4U8CJezmKLV5xNN3uj0kGFGv0gl2QN3fW0peqhRybinNGjxrMnVD4JjFQ+A
719alZqR8wBgu1ZPBmdaj3hHSO8O6U3cQKgt25eOA5gpsXvQQCqso5l5tR0j/DTLbRR4sW8Xja1D
ZWaqKeyxz2MGiCADlfPC0dpyZhG8T3h10S7H5y6QwMv071S0oyUaOBa145Kq9etoNv+oZFMNdGt/
vVAhOsezTv0YQovTa95L4ACO73Y7P09viEFEOYyu6B1oRlk0qhAUcBf02/XK/XFU3NvPR4kD1OfG
r/FQI3YbJGIpfGLSbFv84vHjTQBxfajtS1h8Y4XEgqn7xSq4o0KdMV5RIqFa17lVJHRCVopJqq/8
Erb1pG47bn1tm7StqgiYk/emVPxwKdYe3jFz+5Up7lK7m0QleGnAcAJjWXuRBjvjELtznJ2rf6Bs
IA/GNsEThhrAUGiYdBcTBuVPtn4C71hZ9Y/14VrE6KZ32PzmeJHbo3akSp209kpZDcwe0cXPY8Qe
Anrb5/0tRYj2krtuubZ6d8FMG95e7k+Qn6QnCLNbCFjFRlwgHzUltsnkUWp43H6LWqOtEYiQTBh1
leUWc0LjVS4IfWS9rLWeEwc1TGilVWJxcaC//HVEDtnA6KKbWLOjMzuJBGCuT1uOlQ3Krij187Uo
tiwXNb+FnzY8SMQZbhTLtBHInEZFQ5ZQ6udrGuUro3fQs1FPUpq0KQq1g8BTuyNUhMMNPI8S8ena
I3NFtFx61ovgYz3Uqptijl5vUgx3nA9w6GwublYJ4g1CaY+mXdqvgQyc3xcN1i3unFrFsYt784sV
TFgYwkHQGuWiTE81BoajVx+aCzQZLlzZ2VQPRoRESbMkJtzxw0FM9b8xrUkR48YUT+pFNPdThqHL
vKAkb3Avtk7lXlNO7kWSuM1+jpRpwIkZCKFW8GqKPpo98HFacXzUmdRt8rGhY1RbfTQiKsA4G5nC
4Yq9RVOubdUT/5lylMJxLo0LOtkUEjZQxW4aYLn5e3jOMPVjAouHvVo/e2JmDW0ciJfLsP5mZJT9
XrVzjzeht9vjG6Rs1AT0y1X8SlezcTJo/TMZT5Mf1kg6t4TmFWz+Uj4Kq8boVtFu2pBd1z9H7l6X
WeoIVuQDlyu7CvPw7MAsaxhz6UJhaRdw2el6m/FcxT+XznVIjWh75S/eYwjki2K79z1BEE1yYPeg
7TeIjOO7HohswyudonUgF35Rll/ibEp0uc5xdUt9EtF4zwAB8fg+LWf9pQMh7qKzH7JkgURH1AZC
2ucNjM9ItvVy9R0rH3HS6t3K2CU5YxCGDFmjNv63E616XaXZ/T2KMNDRtxCHchu9Q2hKLwSxDUNZ
WX81kuFOHVzEjJTDIPjbB/P1+o3UAEIhRcxrRzd6XJIqDlqRXrQc24Bk8rajre99BkBDYmghSWfx
I20Z7cxSK7sLALJ9Cum60CYhALg4OHx3Vo7/Z75c3cX/aOUvKDtqJqLOH5yTWbKCdfcxn4igGbU4
jbFfqZhwhL8abNoAR3t/6jEi3D4R061W5VzYKOIh00smWkpcBBQwVjvcxcFd6BREIIndJEEOVLYD
e4ooat1h5pjFbeHIQSQ8W48v1zO4Yok5xXmudmY+ko+6lTCCpuKuHaR28i57hxWln/JktHue4CMn
P8hACrMZGN8wwkUGwuv07DfMTxevsO+2o3rJ9dTJbIlVPj76mR/x+KH7lPsciTQMyHS2i6pVRTaN
2WdENvtVLiP0bB3C15rujEGO4agfZRedes0dEqBI5wKFmT4/9dz7013fSTeigcZI/1HupjkjbEjy
MqWVuDhjDYsACtL8aQqpesKlKCM/MniVe5Qt48AZNt4txV/QtkakSJ1rmLp7+kLRf3swffvuu+ib
LuWCI6v84Sqmhq+QFc97K66jTTS9hsxbu3ncqwciTyltFa1+NWreBQBpvXwieBP66PW4RdgYMr+a
a6ehMPTOGcWGlzH/U4rxIAv+TR+K6NAY62moQnTMaZK+ffnBpG5CmTRsq6iei0mboriMl6Mice/e
zlMN1NHB9Pa6hitvYg36I0G83QbLiTH/NC2LA/u81qYQW30O4iUhSGJHxUr0bVKjJfUAHsJSS+xR
1cW5v5ywxpPbAYkNRJ3XOfVMRee4vdjjwm9AwE1JshwRQ4ZI1aAfQ6sFmGRW/UTZwdHRBLimxvZA
XFOuerqTszdhbYjRYXuxz+Z8AORpOUox5JQ3BaF7JWDxdIi72M0OEmJ4SoqOL/hMqw4pQ4gkks6Z
bjm/GAm0aOq62ZPeLDg7NFdQDVSPZUwF8XO79UMF6LGu4hyGT6gUyf5tSvqaDsZ1lhB6DitKMpoO
g2xhI1tgZNEV7ZeyowmJkCghmM4Fzsp71PygYPIuVHPPtqKnQzKbbhGVtN+iBM4g5n3xrdRaU0se
C93iLaL8UMbqEG2ViCareN7UkoJdlVxh+dNzrkoaJquZz8yGu7badYVoQPvKk4++fMKCqgQ6Q/Ef
COazLTiylW0n8ezlqhHMWB5XHLr9xzXMDTNQIxuWX7Q2wbKMNaCKrvlvNdI6ZgfAl4Duuq/E84yi
s7tQMcJE19CUJH6H2nSCqV0vz4+gjTX0om8P3OA+dYHNDDUSjW5v6rawjSxOOsicYkahQ5tpsDEW
7A2Yw3xDLXPS8yB8MoSTX4Gby0Uv983IA77lNW39rILUVQ7U/FMdpprNnfsWG6UuudIg2Wz4dYfd
/9ra5gmiAnFTw6Uev8UJYRyPhC0ZCsKPs4cGHcACyDYLdDECCVSHNHTDXxiU4OXu8rhc6Bsf0KQi
YE5O3RYw393seN/4bsObSnjrFo9AWKVC7hQ3wEXVtYSJ7nA9Qe2FM7vRlmkpHalrc33S0GNrp06G
jSlJVObLS6pjoIsrWj5Ji2v4wc/GU+hRcel+t22WHyFUD75U7/2bY7T/MUo8GANw4rbprdlv0Lk3
p/9k7VnyAz4j9WUIHH5Nsyes9FtZzGpWUodM4vSClET2VRePTY6uyYCDY2ofIkJlthugxFxqmsSk
wBZFMyDxuqHdzPQUWbdcLMUkF8ozI05n/F+HFVAAg4xN0tRYxP7avI4n5F2clI0cGrzb8aXeUjvF
ohHDhTUaoMB4WgQPwusmZDyu0FIfeff0x1+pZyY5uIvxkpMtRHsljZnA+JoZdmLSEhpV43C/hm77
PJTcf/Xppmp79Lxg86zIoZ973gW+qVPAU2GjaoPHDVVRclBkpZTUX3rbhDxTT2dD0tW+Ex2RTjXb
OyZo+idTTBbiyVfGyzq+hBppCNimBRNcTTdIWnBg3Vd0Vwrp2i9avrBnYPVX8ueLz2lA3TUd0Ee5
cZlSbCtg6W3kvNDfx7GeUF9PHf9MVjg3sjaaYlrrd5Aik/Fhge9R709ZqtyjiKAGMi9ZaXDTV7RX
Or/54FJ8QizSkQXCO7C0yQ0SkA/2x3utzBx5C+OTXBwjPIr1C88MZ4QJ/yRD4vN0YmSvMh8S3QHS
OeQHo7ByW7sDSS7wr5yjU0h3nu7OWG0dj67V0RlLpmolwVN8tQcnJkC8MSa6ArkxEiUzeVPobmSA
f30E/754jqpkjqg7E/kNLlBGjVxao+li9Z8MOFuCyK442hCW+O5Mb5MMuLnSYUZcFXH/x7h2elS+
2N3085IDW1CEE8+4X8SKtCmOeaA6C/Jlsqoi+VxFZ07zlagDZ5kjZFuGGKubH5N2iJDieTRr8X2h
RvjwszksauoqzpQTQtDhH3rVbI0gmLSENiS3sxhso9oYZdCuqXPHtQpSxa88SO39n1FqdgCa569i
c4rSNRIu4dUaxBiZLaPSJk10wxoclUGpemLD8NMWny1UFe9b7OhVHQ5Q7iv7S0/5YTrjiHVLIQPW
adjdWqXflfdHm3tDtY5qcS3V2RfZs/TWL/NtBgYUMIRMjJVOMpfYtpPoeELlCZ2FdxNfShsYNV7K
WHZ+sxYg8stGJ9iD/LnBIT+DohzzVP7vCU9bhrlcUBpNtVW99KuSxHAWf+eUSwilYS/bF6vQFinU
x4XvwWHQ8muFOMC0rSWaX/7T8tq6n0AMpq44wvd73ca2IY7xMxlfP1bvIfzGt2yYLfHHT6s00N14
xpFK1gdZJW/nM9odsaH5DTnrQXvj9RtlGvZdUUuCNAYPplpE7bFRI8DpVkMgL8nUzGdKy813SKPR
fabJecMC0SGNKMSn1ZHSISuUQwU0q2KQOn+p02DHHrNccRiRkDdZZgh/ReWlk3hWUHoRB2CZxgo2
wxViC8pPC4eYj47sz0oKwKiUHx9B4juwNr5Stnjs4sSvbr0z+rgyGFMV9B18eUJSNIXDCy7r1DS8
WCIJP8pnDCJL1dDhCACJl54kkHvUlog/O0q5fvQwblTmR1Dn4gymUn59JYlR8vtfB7B2okVzT12E
3cC2KomckvmBJgezTN6o367FovbUY02kNkH8N3RHtX0bENpcGy5kXBy2uZKX3W1eqCEO+tG0xDTE
CeO7O9P0At0PVnoqhUSVMxaPpt3l9UIaDE/wnxepWmNDYjHnl1zkZFF2eruoCyXbNOc8JwLORtB6
jCjwFRbdHuOI0v9LH0HY34ATKDcTUOTGagff71GQIBZOmHtfWqymiwbizrUCnamYrqnk69wfmFiC
ltxF0OZaKIPVY8yIG1Nt50C5AkKorIF+SR4Ldate8Qhlwh55/3zD7Z1AbM+cAxrg6br4FYn/UoA+
+M2wxGN5NqD9mpHm7kMTQwCtGcTxjxjHYUMVtR35zEuOsJo34z7Wdqc73Sf0DEWCYjGnmgLwYu58
RgOdlZxS95+KlbOBCzvuIzDKSDoKQqRYioetLhLR4wfPUk3Yn4aYdN2kq1A1ITaTD4HcmHtDssyV
0ToFKHjeNtFn5XaFZhK3TTrAu9GZnFjPe+xShgqKwe+GSjKkO1ZiUsPcJfZaGaA6fVZfWlHdoRt7
JDBc0iZ3I5O7iISojP6G6Sy3ChaKKcD8kRzsYqGI96OmKBMesDXqgZjTl9q3XITkBNmeNXnVeO7E
/esRTTujEkLbQuz/cWvbWkIAFf9FgxYGXeD/eoUluCGOKW/vC3cr1xpvqGFCT/8rzm7iiQkgz0KT
4RlZKyhQhBW65Z93VX3A+X3Ovx8pCUuwAXS34BFXZ5gIv/lXL3SX/9EYW9cRU4Qv9EmbTMWnFc6H
dN0XVY4f+KsRfySQQ7bBZeVi8xkOh5z8pxnYY18yZYZCmgVgMipwp7R+FyDheOmynCasqkzZFwdz
OC0NTD8N+B80izBRo2IUhOZKsCInVwzhcpbiaX5LhKGh32odVZUqzgeseZ5krmH5WKZuac6XITQK
d6VejCcHGPbwmY5n98CS3KaDvNSfldxtuS79hsGtGP83yEQgC0LOHzT+3vAcNlmbYDH4ogLjt1La
1YMgunUdvEycoM0UcUVfWjF4T8xwvDkEGvP/qJ17faEgpGAFoVi7oUCn1R7plh0KS075jU8JWpJq
9zFwnPfYEvCSOK/7ZnIsznbVwW1uVpF9xa+gAZLVHwleGrvGuUXothp+ECa6OAeee46McrVUG0ow
oV+fsS0P0XT00/ne/GhOkxwJ++uDjmVwElxLt44r59mSx38BG7fdwlCSqigHy11P5FASWwn9ROYd
A9zVLFJax0zg4UfRZAIMr2ETSF3me7btXP8bWrWMAtTxe4z998I2FgKkQm8YJH4T+fqKgSuRyfg0
lVMydrFnr4RPm0JXoLrYGvazWJPe+zLuqw6mTAVWMYobJflsgRSplD9MmJ9glPXo1D4N72FcZyxh
3wCInAi1Auq39ZVmDD1M3A50mtYrQe5QiKBp6eDr3/TWxZ0hr/1p8hGZzgjr2GhuY+jAH5SPvPwd
WCx6Gh6Lg66ihDzGAd+dhCwSLcsT6lf1qi8BxB+0+xUhMV74BxCQgFz55EHduIMtnoB7VTqLnuRn
8zE5OP607pG8jraMwnVyzqZxcp41e1Btv1VcvnuN2xgeP6AT02ChAGhzJgCdLmqlDxw21NPmDaNW
r0MORMftLnRh9x0N+Xrf7Rg/T2lBRrvXwqjrcnQZt9+7TJt4j7NJrMaxY3s7EiU+186SzT/dSbM/
y0OtqdOGVmxnzMQlkCx/V0tn9kY6aMuViiAtlQVoPQwr2up8kvZl/cdfDvNb5q/2zE+C7hWpvqi6
OVw2wfMeaHT1bU9kyK45mJafkootnkb9+fKDk/FPI13Mmg7jzvFeyxJkGqlB/p1f9JVUE6dIOJTM
7ShdovrUbAUmaQYnlnuH86XPlb1Ko2MqQfWK0JVbtzXulmonNK7KdMCg8YCac1gsE73Gz64xZ6op
ZWjPOJDmFiIVLid9nrcVFDtzyfzZJbFcyGQUCX4pLg8x+Ndk3yBcl5GQjIjptnbwEnhwGBN2wAw0
UpD/yjgaf3Felm2wMOfW7Ww+bIsw2KvneVUiH1i7QmZFEKh+pTYZDPmmnQQkfX2sTi6uoBZ/gYND
BHg/N7fdNjhTSnJzAjiWAr54PTQ9PUOAG+N3LcUsCjUCn8eEees/ljzmCXeHapTlvnFmsDHIX0L9
PS4f3CuNhVZeKhZ+TEcAikKVz3d3PIKKDNHh4zFNeVwEeQqhlSiMn/DGHG01kAdel2rk9R1Pa7XY
+oimP2gkKahBGYRRWaGooovXC28V32mTu8NL6Mih7usYYZVqqM7komlvfliZG/1FshrPOSXywLem
KmmrA1QweMHpq9o8OgX59LSDkDlanN+VbGM5BNmWraeEhpx5SxUSS82qUKju4SlkiUkIQIy0cCA3
eRVT50aHv9oZTHgzWIHjXJ0YDVa54FzqLtpuwrbr1+cT3EBz7jFCGuNHCk3MiYuEL4t1dVENc7gu
ZIFH2nwsmBFb2ZeLthKMLoFrKio9XrnTuBVIZwMxGwGT3o5zfMvA1Kr11ZHLewOLWKa5/98N5i0J
EBTaGRTCa53EaRUZnyXepQB0efyjBBvm9LGLZLk4ZhueUeBvDvV4ivTasv3CtjFiF3JgkJSvsVKV
yG94dnuOWZ2lwp7aWo+X+2E9k3dWuXEnSxeLK/eupQ7vJ4QN2H+QJiBpxXASVpFb/pcXuOv5Hagz
alzdofOKVU03nd5qd9sUdoY+OQUaRayntxO4PIgBNbLvseMVv2rKIzWlUMYuZdZbSfORZQfu+xJI
W52zazviYSXEB3vls4UnFIdHo3ZFt+yMMWdoUgnEQYBkM2BbzyEPh2thNpmHDpOOyD6u772uZwgX
mboPwAiBPZi5ZnIsrU9LZs8qSnGo+chr2sgOrW8+4UOa/w7OzmDh7zty0UlOP3gswdvXUZcmuiuI
nYypFyzb/5u2lBA3H3+RosRGnYX3o9RjYVAIMq/FRyJvIkJxh6ysA0Pb0A//9GcqVQlQHmfvr6f6
lx3tFabBa3sU3WoPvNCWCdz+mNqPiiIdQm5O92PNw0bOBHx9QHuprYgheGtUSflnn1u2rvN1hbHm
elsnPsVJ9nikDqMrjlDxhFUjlJqdnQBBdWMhlDBJztNDAtWNurGZCpl1q4dN9t0UBjMvnQh4zXWC
Tf64v4ZxVuhfXgcLTO/f9i8GLgYnSct/fXla7MQYS7afQKgAKTVsXYE8s8SbBrocCbocxHRY4+jw
wkIlKluX0fEem7lOOFzaIw9okQKd9iVDI08fS2uTetyvLErOl1j+CdOiimuXsKcTdF9LOcF0dI1I
AhNNwOLFH+hKJMMc10OlVV/rEbN0MT5kKyPmpwMN3Uiv2DDA2xjzvJLm0yA0vWWJ5XWL1ZmyqSBM
ZcTxUtsCIrsawNt6K3W90TToLM+9g7z+0umNAM5AhjkSJdbUyHJ9JDEVzD508fOViuJe4mz3i2za
JGy3VQaEx49H5poU8UQXidsWuTcLA7kCxH+3j/PZj+W0EbE6p4CZxscNV3sie0yu1voroSADhOd5
JJ5tcEnhAhL8OqrJftydB/DsX1eDnCzS8gkaeiF9yLq3ed604x4SdXNrWB2swKwCwuDkA5ACAuMY
w3Dzkqwe0P1gPpH0FogydZzjmHJ5fTE34ZicHfe2/Jm8bo3EfT6mdSg2CfvoxD5yP2a0I2co+rRQ
Fx0tqjFwzVIGLA3NlrwEuU+FOzv4bX9Q7Vx5OtZ0gCyUqEuthi7kOKU4fSasiZ/Yr+Oh5tvLhB63
06YjF7TN/VElYAnN0bsFG4PbXU4IVnfm8AdDxGSfq3mtnhbyMLYrS9wVxx45iVK3NdAxbFQFgLKE
zlIF4nof+v+7SuP0y2SPR/CKPA74Ue2mmrAaJGTe2efSEbORoQyqMUbx9VhJ2yhiiqV1cjqVjrQ5
SoNMYsH2Wa1opaYcko0HEblspOR2HQ7I6v0bhykOLX1ix3OA2k+53NWyQzdXwQOOWEGuG9lKWLhO
VqLHxggBUPvZGkacoj9Ycy8XvCHXB6c+pt8cAqSTobXDnn+CEWbf4rp3hrB0k2t9GW14MYR3Jcah
QGJtrSTQrvmDnepqJX/JZuXtrydKkxwJUWt9KqcSvFRM8op5KKKMnIYDyuRfWa28kvnqJg9Pu2Rn
8DccKSsxsLog74J2o3HecNVySWpkr2ES30iGHmmpreZ3dxk9n9wMCaXVfxPCiG8x2AQ7enAbOjgQ
1W1J4HHHYyLtOQpNkyIdoF2puQc81atp470LPj47v4+gck2pjgZQMeSkLREmt7wt6LC61M1te05I
95UPJNTt05lg8rx1ZJwCdkIOf++V3uV+TocJ+0Bz7TIKUIVCp42sYqKE7Uz6FQaN1bLTVWo5RfNH
JLFsnqOZMm4knrPifH7zL4+60v/xHUrgux9D4JjWTmYH7R34SOHTcrhhiTFIX+KW+595kdT703HT
e7Gmo1Oe6U7ZeGjaSHAAewN/S7gesY/q4VWrQxc76uOUGtGq8PnXdnwwn5gkUA/J7wVod1zKBZ+F
5w+ChRulYT+lMyMigXx1EniQqpXJgTfS+v7yA9LNGF3UQjy4apD7YgH3v/nT735mqpZ8As+KkfZr
wEcEGZT1toXFMjtGLs/lYvdXIDXhEsfGJKCKX9l2YLgKNcXmzca3WIO0ckPr+l4BiV2dEMf9B84K
hXNKPLOFvc1LvAiu1xhDtILfshGVjmPS7SILIpD4IPosfPlLpWgn2MdUw1WuilOaJe/zjKyOg3xt
b2kngOlQkA7GqRTP6996VHLTuJlp+lw1gng5I7ZNUw3aD8NOWxek7st6Y0peL3MHF87fA0p7gILE
vmt/Y5x0y5p1BGMVC787yId6XtG2nct2FxtDhNxZ4lpDPqpop+sYsJTG9Y1fgjKXj3U4sKVkKdnr
Ds7aYdWa1yvyqcK3nRSl9Mw3zRJ27KEzzOlf88Xvalgk+gzRfcTusYW7xg27m3Nlbqk+ibce13Si
AqIRGybTYxSdNg+NqyBbVgnRO5wXQNelgkBjl5GpIH67GTd/1272ly9+h/CsV+WVevzLIBu9HKpn
Ub0r1n+iFg1P4oMek8HvyO4Ai5efZVpHmdvwmYZhnxS7xKWr/hi73TFijwEPuD9hBxjxUBQGOIj/
+7Z7EwEoKRwi/5EOPVpA/5xxpDsdJ/XhTlQ5Xq2d2lQISugNgsCLx1OZJ9XvjxPe/oGdqy7M4v/U
hCK/uiASLX+4ob2uBdlQ9ZN8qRC3isyzMujHx44+pQM6EuCH/TWnKG1Xq8AAIRFWR/6j9vHggzep
S+Zk+xbGTmGC+AKk77XDMcY2w5/2ETPhGMC703njF8vasIS1KxOXZGWsQGlFm+dPEPTU3rlGAkOg
UH1Q0vFV9CP6hEMRZk19DSvXOHAYItUoEkCHu9YHZjiIbnrlL9/ZM/CwDVhIFRpBw4gJUoleaGio
UQ80hN8RBSKTJP6Z+cmcPp8KKlwjHxd2RKTmrIWSqAw72wSgaBLrmND8P97rMXh7bym/uPXm2YZV
4py0p8oBbxq6V4INAdN7V821D4ffEDqFzhbYCApT1eOzqZPOd3txBeK7Wa+yxOQDljjYSyYhZQ0N
GhkEbUeUqCDZ7CCUZPZFjrFNs2PHrIMB+GuhcRDHuwDdWNl8bBCMpqOOUlqps7Rkabl2tpZY7apz
94Y50cfyQvpXnBvRbYEFFesxvu43TEtHMu8FOLJ+t8eGTQJ1yaEUpv8PVwVS6pYrTcCGL4TMIQWo
+KGAf/eglViW+MQO+CgE0YT3/d8JszfpjoAqG//T7zpk+FUuYedJaSsVSbFEs0isQ7pOt2wvZCYV
u+6lW6QgvUusuQEIrIieHUWbnois/xmHZzYfuonrU+KZ5rg2uRQ1fuvldyIEKFzGpgVNSenOjTiK
Fy/KLGhS1j4J8NXlKBExnTHIKNrN9B1LuVD2yQiobETtADN/TPcFcVLniwHn7LKurx4ml9Wumgjj
v6g7LBmsxhmiUxw0C3AJHum0mLXKpJE3mKF+g7OfP8fLz7TL877VLcdKKBAmWosTXwKf0NjvChgG
ecKscr7ySndU/waV1RYZ9STlNhsABIVg6ug9n44nScr+jNkmY6pWG+4dytePgNzVQAeeK9VH4l/s
9bsyt6z1g8NzlqyjvMtJr6DBeTOE8TJaLE3H0G+68Cd4vrSSVJHYim0tbrIY85HKIW69I5mdeSXF
sK9PuDprzAMhotsvHlwel4vn+GPf4ct5oJwO4/1ayHpV/NDWRUjZA20XMm3IUV+l5Fq48JhAXGK9
sHr/jxKUHk2a/8xtoyxWJpSz2WDwUaWsPyZuWvI+l1U2m664UjN8Nk1q5/jYekNoU6FwXPeR2sL/
vAraFfQh3CXfOxjf++j6g6cFFqGP5xf7/gFRkvSffJvsKv1P2ugB8J5FOflYHkWHHuV9M4D/Whox
SYfnC5giUuxuvI8SrLckFwldoe584MSowOheUjTxSiLq/UWPgFOI+kn5LN2hA+W7PPbdHmVRult7
hzkgCrUHe1rLvPpGWXJAWXTaCsCp/nYaEuDCzDc0ZU2R6scLaj/5znJpyNRLf7l4DHFAr5gZh8he
cQ6G92j/KFskpJ97mG+ORj0ksmDuq6vjIROhNKgz6maSpCbyrvDrq4OE1w13GwhRGZnat0FThVFm
W1+TjAfIqCOMsD9rjxWx2XtLUJGuukRO3Xy9ayAYpPWkd4095OJE51fCmUFlDh3zUOn9BE02z40a
VAcKDEpJJrX/esHB/0rcr4DaqlblzprgOoGZdsZ6MT0z+/7KFIAD7lI7e0/DFd3fmrJKC/qslO5C
BHS3dINH7tFwhs2VncJOL5ZkU31tsmmdHWzRMVjdmM7hTVI8mbf8dlgeqwbHUY/xCGzcs1wJXFSt
5hjGAHZcIlSqNNBIxGxpvbwBfuKdn+LZGWKiyEc25BRPy7l8AUB7qOsGNnXh/L4GOeQ3wlepP4Yh
E1UZiFsUDCMqE6Dyk3P9VF3UoLya95CahCMv5VINl3odsIYqsCiXpathtRR0CwyHc8R99JfP2hg8
nqjSvC2HoybiGglcZda1qfCY9T7YkJhWAC2v7qKBan85mbpEq7IVO/9DjV4V0pKwTWnPrW90hCyK
FhTmsn64V7WoUXRjmCBtZE1xDilJY820wMBbz5SZ0G3HnD8XwMUo1mdJpnCHu3E8QtnQVIt4KMgw
Z7+mxYyXJ9dqXGJWDqSoy3RUDxMCOvZS2AmqWRR0xgkDkzQWeCRMzt0h/seahj/+9zsQixBTlEmD
MO9cHCvWAG/C7tM93ZGAt/WRyug93XWACXJwViLT1ew09tdhUC60z321NPvnnLix6HTLjNoQkwkD
+K9oXSgezCCCuFWZuUGeOH7/s9DtHLlBDksTWAH9d8FMfwiLAK4AoETOF+rF6fAW0kNDvw6XjRY6
FA9gLcKTbjzYAhmmMEX24W7QAf3BupFxiOU/ZIjGiVv0d7l86bvasRg8w1zf4z7toTMC0pIf6kC/
73yscGLFL+XULnRiM+OziLWk1BArcP/0orUvrQSZiC4cMEwToRLJRPW7HDMybJhN8KEMxv9RfuMr
ufOiAGkXi1gtgUe0RlnkcsRd+1uto1UqH7hltl47fdnf90BVinlni2FIhtaXH3XFm6Mx4ETW1snB
LlBBc5CUZY/OkcROhSCicH3QH3Z1qZutA6+dI/PBNtJoOgIylRnL5IQGd7Zn8gEJwRzQTXNb1p2/
6IpQhIeTjxq8C5n5gv52E5wMZgx0bguNZVSP66QabKPnmtv/ydiPYGSVY/0yWNirkT2P9DayMFTJ
o2z2uSVZkcu1Pu2/QXytKK3vrOiqd9YEPrzy79+ZBabe/doiNjZImxMxvbaa07MDAG3HrtEHZ4mg
LSvtHqJOchGqQGI/UyYIW8zlPmC4eeHoGRxj0SABZDrVP4x+Xeytr61PEloS0PHS4F9buij1hVxU
m3bJsud7Z59s5XNIT/ngkD4kgZy9pCqgvy/aemd9mC0DRTuCzH881FHdQTRboqEmji2fti84LXwn
XsVDtQV4NiW5k8WvlCNThZS842YPOnzwEXjblyZEFSe16XaHB/Y+OS1ypzdr4FNWXMzohAAN4bRu
CX/o5wmm3m9rFqdhY8VR9LK+fya0STHzPMzPWfDdFi/y7sI+mEaTnXm/NP1t3VGd30Dc28u68Mkz
+/mgFB+0L3jrML+wo0IfSrxjbj+Kx0xhRQYOXx0IaLdbrvD4kpNgXBFxKYG6eWVJ8uX7BNocBpUd
pbukAIwpR0BCdalwR6S2flPzDk/gwWHyXQcgOZguB1AZ/MCHPqMsxOymoEER8yXDa9gguWdpKJiF
pqG7okbMIrAIg/qrIdazElFc4NB9MRZg6p7G/zJkKhsqXNp79Heh2Lk/neVWTEVEh2xvuSChiJUM
m42vslUTLttOTf7L3c9plPqpR0VCkM1aswvZcZKwPgr4GBcZR5AHMNtWWJt2PjawqyhwuZeoKIHC
qNis7yvW7JIcAXzRWzFCiocbAKZXvRHMSvNtt/E8hmjdwTEPLfL3n4r/ry1zJ3cb0QuWIyaNaW/V
XUyJVUxEnyRyLqBNXN4NCnPCx/cjyhPXxX48TpfKYXNlmeththjDw+vxyYCFFo6ieUh1tM/aGD4S
UtrDUlE+jUsyFzlZCFCri/sQ8WF09+JweJcbl1r71d5Xg5ih00jmh1cPQzRZAC47tLXY4WqLjTPz
+yUqe0jZ0xOutOvMdgA7LDXtVlgS8zn85kjWouDLqkW+sk5tX9UfzxJyXo6NHUN0EkabNNT6BYJf
eM10MjNguaW66mJmz3KSDH+cOeme9/Gt0k3XeW8GIPpuj2gi/Q8x2Cdg2WIosTpwm8eMCDTq5hHp
PYB0suTqIBgmR+JEP38aWvBlgVRLb8d1iRRkf5oYFYRyubr1aTV/LpGQMJu2jTCM2d1aPYMyNzHi
cOvwruS9vwFfiMRHnqPLySTnYkjSzuRTase4By+Xj3ZJAgRD/HKv6xnXDzsfFC5qdKOthZyBuS1q
jFP1b5BNHv2Muvg77IcrxnDMacfr1kTbATAPZBipqkZkuM4Ctt78jXFyZVzuc4iQQM/uPStO+9EX
fwvPdfQHpP8etigpNnx+U0Mc4dnvf4QjnpsuX9pYj/BcXzCg0/SZ/aaHO055ItnwuAVn64FoxI27
Ei7dXDQdcJXMjudCv0tULe3g1bSio/yovRz3G1QQalH1vZeHI77z1ecYm69ToisIvwADv2qhNpJU
mJU2ZDSd/gP+sbE3BLhT0FQLo3ietx9xuXCiU8PMAGdryte2aAKmH/iD0BxFBJRv5QpDIYHAYUpO
kdGpVMpYa1H+JsGtR/ONg1WV72Oj7M60/GC9P6uAJjoUGjLknydvMQIWDqVrHgbWyLuHv5AK+mW/
ZviV1gGkJQjMx+lNspaJGFQ3/pCWDcuPt+Csqw8wpk7WNcQQuVKcv+PZJDwsW+WbW06CowDqVvfP
LF9cgt2JjIFGsMPIPcCBQS7yJs+VO1+0gSITImY8GqHHVal9WMNpIErhIwq/3gnyQaJ3EepIyQka
b0K+bMbt0AhQm3HM74U8a6N75ejei49mvZdYy7OvTp5q7H3UkCi+o6muFr95c/LQtgZcFSwEaUTB
yox1iJffuXuZJaZCZqLR59ToYHaCJw0Q2GFI8hMIuljCjIssswLnGUyIuhB5lII46pVCBfIdHVRB
tUoVdAyu3b/BgFGW6vI7femXPynBjsKsjk+JZdtGbLfKOlUq+2If80XTFJrlc3/igq3JXBsYTFwA
iseyvPgV3ZQrHbeZUQPuLbFPkxBi7uztlnUXE+dTpRGizJKxWaM6YAUremhlhiFV0+G8VtCMrOG4
jnQaqmYGxBEJRvDRhQUMvRVORUPYlNuXU/ioHbNcet+NFhsmBpejRxU75LCGMCNkjBKo1r5BHgqh
8am6uJMXmK8DjICWZFavxWoI79ADW0sSOGWLsHIHsHVzvHFz8bJjW0wMvxkz2apgaDWkTeUDUNLu
3ZDJjYvtRwQnD26T9PQveeExNScpvf9oPA83rZ9dK86rORcTF4mj6OUEBf2GXUUhj7eBaDY6+os0
6kdjtMIuh7a9vhIPtYqx8eD/NaVAe8CNcK10aMc2NAloaosSdCd+GD8ng48B0CXSIQrJTVLx/6Rr
81o5WvwcYQD/9rAraEVn0wjAmaJKBwTSyc2pJhKOGZo002bVanUS0JJPoaXRjksCI5+pOcfZV6P6
a3qkTWS68nczbIdvSVdVCedDkMxw7n0EhXExaOcyC5SAbaUxVo+W8ICAovAksjKpL+aR8jlDYFG4
NlW4LA27FN9tqrNI2TIJNZey3uv0TTVXSQjA9ONlRqWaVqYhHjw+MOBO3O+GmSe0NXVOMTmR35Ig
S0Td4j1MB3oEZi+FQnxRvmJFaWjHLPEW0k7IHUdhJnUZNAF7ikdO40TyNRdhZIDS/wJtACbZmnW8
nWGQhMw3uaLpWIkDtY6ZWbtvWqtcPO51vZRqf9mkpF4f8sYEFBZvScJAw6D+o/MnUh3LnE6SOFP0
n7RRsrcT7zJMTlBCuoBnZzZgDHufxcpIzQBKw0ISnjhs42qDZE/fXfA4wsx8D9vOrUQFWUKYlDkz
wUAJVREfTPYRuvLoRt0PYm+fSGiKa+FhHLwOBngTEIdxoC4QKfd1tJtKRSy4Ls4F6iJGNEz65fhF
Ms0nHX5aCZVCAFxlXADIGNS1zFINvxLDXRGLKnhEzqCvH2s4ilDK/3Te1UW2cmEntz+zJlmIoYZg
OoJrgiAlgMhAmvBO+KOSwkFA1hq8mh7vcaJuCjW2d7H5qlpY/xgTe2xRRTrrZAQev2x+FD90gV7r
+K2jeStCGbPioCclVZQZdpdPejSwtc9KGCR1+Th+djkFl3UO128iNNK2OgMfBZfoC7jKCB+/Uc2a
X5dqPuUDsx38tzmP6eF64lFYXzQOF7A263FfIEPbKlo+X7VQ3tUplUx2rCroDI7YsiFlVPxO0O49
zPBPuni+r/DxwZQrB2ZfWeCSUyjqiqh1P0gzZo0sY9XSKEuWqCkBAsJU/HsH/b6/ZXYAq7yEb6dF
rfzwHnL7o7VW9khmVAoPNjpNTQeZZJSzhLIiH6YXtfFfvaMedUTNx1xYuWGBRq66DjYzHR77h2W9
CPIvg4e522HZJ4jxo62rEW/hGCjqjDDC9ygHoJgeb6Ohxb+DThpuD5osY2JbLdeHiH9MunymWq7L
klZfrRTdW48odrBuYx0iV/IgiW1JAbNkWCoASPVlR9GA/7HHvaOjEQrTtGY48+tA4iDBw3ltXg0M
jNSR/ybC1fi9tYjnDqcsqBDuH/i+1FR6KzRQT68RmNykDRD9rMGlVtDgB9RqQ9KySHMFaqzU05et
tYIo6fqy+1Z7s6hBqI2J/IcLqDlzZGi28NBqoJu5dAWC0CjvATS97282Va/W/G0uNDMJ2GMejzSb
Gex64YHTT9EzFtlYuD7eVw0XFJzcasGk22xEEgCr1oC5aZUWEEsUYMLx6NK+vl2mhH32I9pqq4P2
X8Py0k9zfjEcgwvK2LfWjXacvRKK0rchpWHjTxRctjUGZVGrX//aZ3WahbwghUfca5TF1NukQiOj
zxHMA63GjV8ZLEjXr3eqlNWUkMCPijUDzTnc5jXWLJe1tb2C49SF4bCfGF1f0kwoEC75uovc0n/s
nvFV3z8/WBzOnB1lLqAltmlcTAf59zcXfOcRWEVHtgxZiQe58lqHt2KWb8tRlBHmfqhLDg0bikVw
OSgUpDmbICbG3GKB4+vWNoQsACIV2BkjX65buipj6OQ73+hym+UYq2IFWKK1FckFYnuG5L5rWl/B
Cv9hRK/6Rrmc3lsj4qrja1dw1e3BJnJGwB1YdKufgjJdMaGvvQHpHajoiW9DFbXNaYzcBXdeLrOl
7ZyuDlgMw9aTFJLMMTCEF9k4yxAuMwfuu7N5MkDhiwmj3oTxmoUTMLwH6xFcZ4uxivf6LID8SPGH
t84rJFyD6h3SsdY/raBWGjLl8l6ZZhhmYLN82IK/kwvgMvHpOhSqDg89B3mEQ/jkc8C1LI9/NbGz
eh+t68gU4pIyWi78W6jjNfm0EyMa8aYWpenDy6DhMYyCmfHC98/jXvgUskx0L/m+w0PhkvSxCiX0
+Nz/JFNKbQTAGWae8udBgCDR2F38i8tlebd5ZvxFM3jFVwPFDXIjvy7P6c1lirAPQi+R8C5wXePb
JiaflC4s5tcBPxFZPfUeH9mZUC+2Lw7ZI60+J9TOW32ziN606KvxCCCoQctxoTIf2+YetaeANN6n
kznF8l5P9aHj8cUSTyO1/5QuCfyG8Jnsx7iG7xZzulhtVHQX35EsQBF54csAW+rk7HSZaIUIdde9
RMXKG/uJefBN97Mbmi6OxvEqoGiXjpDPTsG7I52l24BvdfRA6VhqBDmY4f2HEUcN3HVu4UkAxWGO
pLTkHTJEEl1aJlBO+zzb+Dk2Ata1kfr/y4nOcZjea5A+4o48U9DEHZ2usA4uD63HDLkwEbTYR1Zb
7EufokYdsVWaboKYCX92DlbnJ1I/p6XifV8GRevLn6naP/b2S7VkFtILMJ5KaL7wBOkJSukyGVqj
5EvA+uEBENbWEEasz/r2X257Pwz/j9plg/NzvSuBykLBdsoZXU13azKJ56v7xRquOok3whhsUZwm
jwrLYlilmoDXn6hSNsLO0JTc5Z82yXjWoIXJnabjn3dyhLDfOI0MjupenmI8orZ7j9e7TxptUYbf
nUAdP7+lTXyRjFc8TZ/8Nx7Y7PwCiTmbEQ098Yp2ka+3xCrUtTSxU/q3xKpwb+JhvZJRCVHpyj0P
YMdM6gRAmAN4fO1xvlqr/X43y/eFjSaxq+OGwayzNO9IahqXDQknveZWDZoRNmnTzzsKD8Zkx2MB
MA9x480pwwFL/SejxAER3WFNbgVAbi2T2rT+Q8wCOYHWX/N7Bx8NK8rOeCc/OoryeMHmJJ9JUPut
L83USe/SqLlo1acrM+KS4UANxw1fU/smQuITVaXdh3Hnan+dxtKBudFqFtq29qp0/TYql6IROGtU
Tidct3+XRa+tM5898FtnFzNodMfqEpa9d4KxZYLbTESafE6hGVjk0xEIGBqSyKTwlFZX5xcCVmLG
FdQH8JLyH3s8du6aCgv/v1TYZxGJyI3m1lKuPdLjPtlNf2UzlgeIQTQpNvCoVgtxwtzz7ONWkanp
PYysncC1OQrGJ6tsZBjFhj5PxG1zWeO7/E6oWZPs3EtOBBgJlf5KADWXbmGyDUvgqJSBVcOAcWIX
R45mVKKLV5LzVYvvflxCN4i9Wcj8JDvR8UwMRa15rEDM0YB+fRJaUpW7lgx43CPp8o+xWQkmR329
AwNaGLR+3pjTnUhTJF/RuTs7fov6pv+cH+uZIOZOOIAOmIoZXTpCXSxPF0QXAEnz3kOK7n0oskI1
3/nwUxwbqQAtW6orr1GXq7sJ6BML6iDUW3LvxnAUBxlxjCUClwHLpR97nhgN2KzxU/fEpXxq8WAb
UlVb9Bn51jP+kEREXxdg7JORMVBiaqj3FmpzlcUvCt+kMK2It54IZ/LYO0+NQII5qt4ji0DDah7X
UQvJCZ7vRlGzMgTNz3pHWIXoLEU8ya5D7BWZqlkJtzGaKEZ7jGu3dpSIDey8dgSV2GdbPX+cXQKZ
zf+qJTdpWu51BuUQZRvz100Gt5vx6hJHNnh6pUGTdyPaGzeCuiZbyEOfbZUjd1rtxvf4lHp8cPmX
xROKWgSKhwRbiLVp8874B3kMURqoM2N3SxO7a9i+Kohsld/2261Um8t9hHn7PUrkRXUfLXYtl/e2
FetmWpkzaTMi0+usnqHobxWyZzKmjTwqRTRUuvgFmV3PQvkP7zxe3A+fhG+RSBJpsABIJnRFCmaY
IfYTdCabhpfZ94A6FoNX8Cq6eOkRmqEGHTYA5H296WSx3BYhcIFZL7JU+MhW2XPgWzO1M0JCHQua
7PndL1KUyx7qEA2sfV8g1CvIHuwAjCng7PyjZMTFfxzUbAvlRmA6N1+cxgdfHY9na1WE0QFPa148
OjEcJITp88yCedGbgofzK7DF7kSM0Z8T0nyCJc04rt4eAtTgDu3RXggQKvYz7weQg1kixilX1vzU
bXSSPWRu6W7u18x0a4ncKZC+mhT5cAzGDmd9cXNsZDrws2tajk17NOs8TyqSaXREpTUGZh/nZvMZ
0RQ0i8i0Pn0wFNCLN/rT9WpuOPVXeSCvHk7ftjPPoNZdFI53jPXDNzIzwqSA6Y11OKK9YlfV24d9
DmiHR80i7WCC/YdS2SABUAU+DjEn6xaIkNGapMh7dLthtZFFY1sN1bq7yUVT1/I0dcIf6fzSv3Zn
adcFEDptSWcEQEqavLdYqdfbwkU1cJ47IK/V2vZGuQtpEl61lo7biWxz7zq+8YXkM9V2hhhtfDV8
xKP3DI8IvJAgCJZ6NuxJ1PA3pZ+wuBkbXvwE8FMh7qQo9g19kW+VjAphUd8dDJpzTc4CIxxvUgjB
xCjgCnYaDsAM0HwHSg1YAcZKNoCEfVWCeYIAEEw+hJkQdODA/Pg1bfkGcDi/p+uVuvcfOPXgpLtm
AxRrtxZ9swh5kv9ycVOsTdrd4JB6oix4pw5dHIXruKbgaEAKjTVXJCqRq/BIH/cSnFh21aIrSJL+
OfuoF0rclE2XKo4SgG09KfXlRbUN3JqzkacCatVziIEe3l75/rm16bR+utVWB31BeSIPx4Bv/h4a
8bWeowLZa/E01afMqUFAiV+LmlSzvmC2EdC+3+SCCieiQohqEhWXBCOfjVSSWTH2tdC8ICqSElN6
z2LRom/N4vhlkWUaVtxTDqGVEX39QWsrFsMuWrK0qfV6EZra2hrqRVjJ9q+AC4zZYJ0yQnecrnfl
VKzMAZEvEKkIHF03fQiyJ+DlxbyVy/5RJZq7mN/CHpTDNk2dnBy5mYASM7YKZpii6Yz7Ltj62Lcz
cVEHLJwi2iAKVPb0hEhEOPpC5qBB2wnvrQnIur0JboxwMUPtlXMNKjYE9rdOkg2li2hKbH/e7juN
8N67Kv29gS5towkCN38humKRjyhC424Sg0dbWvOc0F2Qu5Vm/gdUpKFAU6+1DLHBNKi1IGv9BQrq
AtkTWgREQKIoPNvsEv7dNIOb+c1VLSkoCB3+oy890JDbb+KWliDV6uz3AyxPoSLrfcF077aT+/il
/uhViKD7S1fuVyeXxodbpy2aCnXWGRFTBh/eGtbB7IQouzsZAr2rZUxRID9pBXvujV0ho4MXwope
+5GObA6nvljMaHn90v34nAwkOttLU7FPf9ve52z5h17tWKq3Fx7JG6CZ+6yz2kcaUWpuNY48rIjh
ss7EAhf3ROfslkEgv7uYK3IFNJUK3LW6wKB7gmdcDb/OWouZFTVKVU+JC0xO0oT/rXvepWgGWInD
wS5Z3p3UVUlZBV+96DNQ9+FyR4G+2ldAsW3Vd785MG+kSkE0asfTTG6ujBVIJt7LU39dgYpADbgP
p8sf+/UouUK0WbkUi1la+5oJAF8dqBlTK5PNuVDUdZgUVrEARfena/RAi9701t+6yJrGXEhWYkiH
XrnrFQCerlPNP3eV459f46Pf6+RG7lofE/q4HDjMAaZamL/0VVCwniwn1jDMF7AJjGsO9qjI68Ma
1ccV2z4bQju5sixF0jbEiGB8Zlb6hz211OexK6isR7utigsQ0y7SYWvh+baqaHQ9Cwauz4mvv887
hdWoLeFX6OhVWUtVEipI4+H7KQ9IbpyGjaZMBnkVXdDR2rkUF+P5U38xl/aedEJH1B2lNF0Z2+sE
5rBUxyz7FzOGczfUAFpXU2eriAw33q5z2vpdSY9PBgat+kRNLdCUBdslMgsczJkvS5zqUfrheK34
b52XAwvIoEKwCNsUneNeJVhb8WtHXFQxd4k456Hrpq8L6fwgJDOaji9eZFWMfCBAG2IQxVlksuxw
QiMxjhCnhDG9MDeS4pjv0FY+O592uJmXCb10qZyd1/QDhl/e2VR2JSZypRzHTtx7YTNyKxpy7lKS
1mpo+WtUaRL6EgubsBlxInWRBLFp6hPJUeQVi4qEGVmZlXFK1VyUCkPZqZJUByVO/nDYQBDN2jgM
g4U38GZCuUOlm8IsY7WtuiRSEq04xMeKTFMAl18+I6LwkZp8lwrqGM+12ei3LzKHRv/OJ2QnbIDz
zd1JjP0WSHfmHrDPs14AdKGR1BCaw86Ane4glVSisaBNzR0kBoOhddbcMZHLfXgZyDjEQKIa5OiG
RAvGfxT9aK8AEbNIcqq2+nq6ef/qeavccaIQFwEbbh/OOjKf88+wNgnWZDgn0q7KJYMX4R0Ogpfw
XghKnxHLeRDTJYMzgCnFs0TVYZO488o2hiv+g//8KDe91wfE3saR5JsCJp6o4VLa9afIyp3gHO3l
09BI5qW2+8IpdYaWdhlBw/V4l0gmBZn9eDMg/QnvV/Y/UIDYQa8ELIGc17HwrBYqdS0euRxv4aR9
YVUVV8ggPAz9nVfIihxNZ8nSiW6mNk+eV5pva61U9/V86gIzeci4014qE3L5BFm9LouKinbOcwJ0
iVX/GaL92eN4k6CE8acHISS9GQPznbeKAo35q3/inB3IPIYeNo8ncL/LXYcwUr0vjPNUjxY+R2VH
BJW86v/iyV162PuCrTyKcjjFK+MJzIsOES8gfEw2wW5gYwo/n/+kV69UqPhLbzrjmRj86FwK1RU6
nlAwI9Y1lqWuYUDrZYnm6yQmHEKEh2qawir4gveWGDIje9l7KhJpLxCM6WV3TqwPcaD3n9Vk/S79
VhWqpUEjIaQ8YU22HsMKxvcfNy4fDFzMHmON/utsC444/A7eTf7NHxGmR7RS3ORLhua9jfjhc8ee
5HqyDr4pTemFWf7gXm5tSF1KPxJ61LuvfqrqWaoLZ1QdFKRrkpxgWpbrgBvl9zSoTvkZ8PlBQIx2
fZ5KvrMul00gEoyxQ6PEB7YXo3z2vlOMLS7WpZWNucI4jBwM9Tc+Jy0/6OCw30yZB19Mylkhr9qx
V4Y0/oS0vDUO6CbgBw5kmpFU9wnOIvhFKAsNko3qdcOjUnS94mf1/SEFT6M3rnwg2KI0e/hi4Uqp
6GVA/lgNZXDW81/8XdFx7QsLte4lzLnepBsJ6wW36AA9uAYy0ioN7mc7HDUq5gWII7cZq7KdvpKE
OUEVKukEqQEyRe/zihHIHZpE4ce28DgaxvILBB5LPTkz1cW/99ptBxI0aDuJ4tae6BbnO5QjrKV0
OWa7HzNfflyXc1vGWWQZsBJdei+XjL45ZSx4IGXiUo15HGqr33lGLtkanwxnHzE9YOfHfcyPp2bM
zX/Cm88JR6OzIcV2zPPD5jjzUYJqmKKgIpsY/OyLureaAq5lkW+jSohCSNhb+LFTM+l0K/yv4zpU
fQrjl1zXzMeNiS377oB/HyE6ANtQo1rU4Ca/tzTXHNRrxFIXeAY43fFO+f0QIumaYKn73a/D5sQf
3CcxJbJ6XmsIzNDa9A4VmkEnWvdaW/QbQWwgRWsG3zNX1TXSwbyO5cjf47r1Km63OesFUM7ZuuEh
ETvswY/Ej0MPkyRs82ZJvQ7MEvSGRLfgelYJKvWKJLLmFeP82XiHfUxmL3Oix5sV3D+dGBEhqzlQ
o4jDT/QbeNApO8lQ4y1rbCPz8R34OuO3IyHr/KLTV0Lq8q1OGeTj1VWBpfRiaWEd2TtlFvzau4Zz
JxpWKiwJ3hjVz2Ih6JINH3EVbwcIJ/vwHucsQtPFsjQz7Rrwy+XftL/aY83xINXekmGL5juals7f
47HtAm8umOgksVZcZb0Jh/ZrtrY7gZzfAqKCK3IiYKEC1hu4dRENX3qTEX6uyjU/+yOzCoxsSHVm
8uyroCZYb3tafcRK5dTaxdfCXskYoMSFsEK3787c9bn2ENNt+FEe6jDGpDKY79uUoVCbKOD4OY/a
RboBSNz+E9Z4VIW3GxMap6DBYal2b+rzpKYvGLiJFW7f9xWV69KWoB441VHHgLPKR7qm68AnuMz5
xkMFwyFTrLIB855RuGUDMsbqy3iqZM9Cpj3f3nImu5o+evKQq0GPX/aRTR+cilLZ/Qe7c/IDFua/
22WqehSQFjXR5WFYbFI9Kgl1U4vSxYgGuCEi4/ssd8qKkN5Tk/lu3h9iVJrGD+K8IWDi9HAI83s9
xXmfZ4JYC9y6MnYkIg2qB9QURNNT3BOG7+RY72gbuNTAtj73LnuC5t5wBoLEPkSVVJy7Ym3Sq37X
8CVvjY0THSdEwJoW2Bvclaa4PGW/eQ3T1NSEVI5guyJAZYRLFSEItU7mWaxgGT5pfnGzmR1R1eGR
SwVAbPsfLNgLSS7R4qkjpyHFoDU1NmeeQXgR6huQWl8jqJTLN7pxeiytwO+bRA2YWdJ+W51Mdi4/
YzV0iatvXJo2RHxdUdnOUfXWjoYkJZHtwSRQ0AXfz/Y0RW4Ue+Xuy96/8t4NGhue6Oo3rmZqjknB
QHzTrcuFUOTCw3HKACAcvCp3VRf17qg1VNBqiwGL8cy/axMMrtqDywcKKlzBi5/c57OwuAhwUvol
MXCc3ltQW5Hc5JZGJrNBxX9M/yssya7iqJQo/6K5AbDlcCMWry/pzcsAsu0F+x2MQgvxoSi983VH
yhMaF7PtRYgCkx9m8wTnf4rw5NputJR8uXU26CX0gkYF4HYhn/mmHlGiZDcunWEpyxOEAsqgMk73
wUvVWx4OxXjl+mv4eJulNkC3nFgl0uLE+XPHerGNuH80QMJLCpaBGQV9q1yyzLWoESdL1PrcMLQK
QD1kaqisvTAPL2WNlBkWhw43EMGHx4Xw/wcLq4XTtXkssgkZUyMbstQANcbrfyr/qq2pbLNRFND4
DjACmCqegjED+fwrE00Daz2eK4oKFD9yoXFaBmYtDLQdb6hazWg+WV7gLXFj4h4ifZ9g5YB1kd1T
Af1GjSPMabKcqK1lyRVmmyuAXRn9GqVmM7PkuXTmJVsH//BEivOwX26EiHvXihOiJrFKrA81Pn72
ZLmcrz/RTDyCjET2Y24+2b8OnK/YgxVpj+SQcpgZIWVrDDudEVi04kpCplTzLAuoUY9UIiCH/41T
FzeWGRPTJ0qfYncN6LYRnKCEFgpVV+u8hrTHED97vNTarOpoavQkJsFiEhpXYKxsPrGAre8K6HyH
sYhE3gegTcpDyj055HCM0taK+wpp0csKA6g6/a7rYj4w7uluo5J0DlklVGp1HQb7VfsAM64x7rbg
qE9IdCFj86qb5xGRcHbcZ+VBf0UBxWJMN3Q7Lo4lqnICvX9LFhEDh8wVd1O9o1CZoDgYdpimfA4H
2LxR3nH6tO5wHTQrrZ7x5T/2Wm33RJ4zZ2gnMo45hhENZ+iiR5ViwZ+ALkani7mPDcDqBwpkavcZ
szofk9pPVI7VytvNA9zcxokYRe+zcvR0ew267m9U/SRJDYYSxUsCJQVK9foQcLI17Y70ogOcw3n3
I4sGJl8ZIOM77lxH20JNYKBopCBPn/TK2mXlYMGvsdEJtG/Ih6prGg+whyL9N58luujQhtvIZ6Xz
Rx9SSwuJCsW4P4/kZAkT1/UiIIaIK8wdc6Jiz7VuAbjwV8LUtyvGmiGLb+qHpE/W/d8gyZqeSF2s
86KCv5k/7Rbs1JTDe0pJospXzn59SSIvev5qmqZCX+aSL1Nj5Vgye0W0U1IgaIIc2PlCmSny+He9
R1X1vtcbwtKkAQFnmvreLsEHg+xCf2q030/fA5uQ2OrLpi4CH5M3Sem1zyPqiY+6AqmZC6e9rg6J
DVthJ+/JfQvfCS0X4/2sLgb4fTx+Cs08JEoacHFTrdvtILoSDndf7YvifDjJJnyytfjYS88SpjAd
AsQmiVohfaHKlZy2bDKeAUnnjNtw+e+ovGqFhtWpnnijTfMWgPddjNcog4wSPdVZ9oBHXuSDcu3U
qAyFUnYh3p0yOrKJ09yoJ2ilFzLTbRHTW2ZSYgS5oRt+UxHxKPabHgKAX3nW+O49glk87r+WUucI
30fwlnZ/P9YUa+EC8cAsA5gur+I7x8OkfRpz9P/IMqXuHMHHA2Ph1xIMdf0ZLPs+dQioJgkvv3TB
bGdJsZkyFvjwEpBVQp14KQNYD93kx5UYeZE0MkwiomuRdCueSC6K+Yuoca2TJ9ZFOnMpvay9L6NC
ef1riHa8dfcAxCNRU5AYVWvkyXTYJuRJ924LwdifzljM7oW2WZtMVwkZjumM5U+9BOeRmb17725K
kzE9U9meeRnGf95H25/fL2plbb2MVXHOT14EMnSCeW2S1i9W/Kp0oMXUMxU0CYKNJLqZFlcBaDIm
7QjKT6xydhRJCDsMnZu1x6EiyJVP3nrPLH9K10gX/+hHAQMe5tnVNbBhvd6Ye39k6Cq3R+eHajcp
CSyoGuB8aeGanbNX7cCm2xuhMWJuASArRPDgvhy0qSG7aGBcw16dzKruy2KBMsdHUlEimdPlaS9b
iMbbL28uALeq5txkaEhgqmQcXhb3n3E3kaG/2f/sPKeQclETn88F+ZVgrtuEQEoTRenqaCumMgHi
aIJmyXTX+FvsB2d/XdMXLWJRFQxI7V1rJvX3GKxKBlQllo1ckxgB4RMhLmE0jGNaiSDMLQgtLRZa
wC9erLeG6hv3BGZpPCI98BM9sPi1F6uM1eOBhDi2gLTYfqlWYrI0d8mUJ3DfZivvj1CYujY/8pD+
3GFVoDfTXEGA3hl/tg33u6qimtl8LZ/BadaJLTVmhggOeFQuGyTaRbfx9M6fB8Q967BMS+cyx/PN
CF2skD7dx0QSSj29KHIfhb2bTVEL/J/PWCpo7Op2fg4qXoxV7kFS4luDi7QUfvBm0z7nT9HSzUgc
20woRHPrwI1j4xc6efg2V1JwmXMoIqz6g9yoWa9AhX/VoaRTvoY5Nw1Geh4jcJoPPTmtRjCMNNKB
hySudsXNxabXdaNB5rECZ5ywrwvFCTNCuymXIUnSFeP8WhyGqUK6mTy2ki2cRjtWM8aeg0F1foAE
/vJX5n319OG+mN9e79JY4yvGpO+FC05DxiLSrXqaSvQn4xn7taoVM0C70WOlVBsyKqOyfBU4Dy+R
NULxisaPTmzPdp0IAV1f4sIVm1x9T69ak6bQb5QjnLyYAmu6U1xTMpaDPbjb33vomb4U/EjVQGtV
YmxzWyW4iB4LiDUK/+eOvJ9x7xhwQH12JGXO15QhEqKKe1FB2P+pyMIi577pmYbp3421Ic/VxJAk
AYgWIoEv9BgGkABMZsLUBNnLe7a4d1ku0Z753m4IHb68zdBtlWqn88pjQn4gtrj57qlNPHqhNnO5
KhuFJmVx056KqWwiRtGqbX8RnBaLjOZQfYHj1b3X72wcfh0K+SspDUGvz71RRhSCo04g6HkNZ7W8
KTC1HGa1fTlww6PsVxoYKiMDHFwcM2jN2cx0pXBfvIc+ObPCIO03Hm+DwzKLyWWg3MWmK+mGI2EH
Xwr5yDS1nusY6dH0Ibj0MaxeOo5xMihPrfnUa8OZ3/O5+IgdiOhEhEiekVJn3A8fqq2IvfNGvjmp
a184l5BKQaHHwkQToZ9K8c5EVjzAAAqIP8dx6uL76pkYZSKdgrnJTi7YOSFRpmoS8w7NyFf3GMtz
g4+AO6aH1yIslSDVB/TxI68bpzwbooPVgk2KLRHyN2Cen+5jVpAz2SBpc7iCVJm9y77wOsnIVFH+
QzCtk/+b26uxVaTUVIz78dYBXgi0GvyEvuivB9CBygLEefuTwzdfWyViQuKI9Rk0U/+xEkg3D7BN
WVXpZZS2NjDCkmcqPmzBBhgjoU/Y4D6QQUKqEW3SItlJIjz8lYfjaIynrHUGVjlxum5fTiwkgWIu
mGVgIlLfI7kFaHDN2UOnPFWtM0DkKNrTLycKErmcg1xBHIbpPssYnv6krz/frRCyzS3v0GMuaufp
xnP6yE9GPaNg8Q7WwDzJm5T7tBq8e6kFFkDLkTvxPaMF3oWfIRmqGLDTcPe4SoG1tNoI+1boOvy8
neEaXBmEfyRisA4CxsLqukjg4APzD4pApx3kd725D2Vml4hcuRu6ss9cKvch5e7MiEzbFLmMXUj8
95Bbt8bATkYQITYpD9UNa3jNqorNM8DhUmOYUkFOt27+4LXrthITkjT9/lbAFO7/XERyEj/8iLZU
Ur74ImFDl3IQe3jyKbIXSceyJEefhtBMSmv7KBTmrFv0JqYkZA0ybfbSEOrHKqsujyaQGdZgUb4T
Edg7etD/j6M8bMUhKJR8G8/XmRc6l/cznglS6xFxLfOxAoNkAC9QmXZ3x3Suxx9HiAexIYr6dg7x
X3LHsRaMoX99TcAU1wmhTVqYTm60L6iJUkolQv0KZkcmF56NEsIfXJbEJOZmXVe3AxELiba7NFTd
f+CpUOMlgq8Ri5fu0gIc1Qi8zqFuIrkn3nIBHng+e2iBanut5nIaXbaupfhybWmnz6GsHAoqAMfG
g+UjG//4O3zJr4CCBFkK1pldooXLQdVO93PbWLQBpcQeflpunbVyf1RoET7UegAsaX+Q4CsS0LQx
16yQTUTpZOKzjkI5A83hN2vzQLRw1jGZUliZYNOqrAM4Vlcv0W/SdsdB7NlJ1wjnoVcrfUX92Gko
Dubmje0qE9mgYF/1ZtMCSL+AYX7gp3b+NYc3/tStziP0IrK9ck//MMkY51F/D8Z5RUkmoJgLJLfB
wVgzsw0PtSQ6CLxiieU34zvr9T9TvpipGjSUhXm2NJUznEmag0Q7zYgyx7BzK6zQYNm1jGm94k4F
lb7VM9isR15wXVipzL80YIhVMF1tZG6mTjKHbbLWo9AfrbrB78H/YA6Ph/mitRZHK36yk1y8PdYM
UY/RWHCIK07/foNrELzKT7ikMcF11NC74Y22CIB3ZoFWJ8J70Ed5ppjMnSt6x8wP+FUXwCBmohhe
23vRc1Y9C9SWKiWhjlQCC5ihIkb2IALmDtdk8xwpC6tlx/jr5QZQiwLR8TQruqK7J4208iuTzmtk
IUF4M7HYHjZCgGUmR1umdtX2bV9jDYtqGl3OHU9GEDx5dCwAB32Thntv15kZSMNSlKEaOuesnFEx
Yz3CxJS3MHNc1MTLQhGajtN0OCaVmYkSOWZXIXR+UqvwhgatPCD8BDnOuV+tXjvKn2GyQP89w23d
Uxj/3sAGxgTQjBNafq4CN5LawvW5DuO+ogGfhpR6qqHKm5mdlCb6MHoylNmDWF1jCkSw1iJvKwtB
O6ZvpDmmLGglpcwqYKTjtwK37mvBLCw7qz0pWaffX31mgHgx3ELL44ftRKNut7KlkxJAkujaY4TA
NuQV/ymEP0LTFTnfMNv7wCguY/Xhd9FBn+fmGg+Mnc90jLYfTnmz1n+N6OmvmFFlJ/BizwDtdzzb
bpGh6baO1cnzbev1iIUZO7PyoCg1jtNXfY8/NlwdEFciEBeuxy2l5JZqx0lcSF+iZ++6K2lJxbgJ
IZiFFVgxMLR2naNYn8bQG5Lx5z2JKEJQGKVIZc/RNz7Owkk25O74iZtHtMLE7kamkFdqFzKbMxBC
h5u7O3cbPbUp5ZVR/iU8XfbAgiomEkdUuHsnAqVkYFhnDQd4p+auMJCxBgpAhS32/rYyZHp6GgNK
hC5Vd/QWaC7+05PVw8EWw4Rds2JceX5r+Lw15va3FC66+TCT+4wgFwTyHlYumkkvCISWOY4Il47o
ILZtXt0+lnf/VxtP4FcSt7V1oHTd6sOVvUVlamwb/MwalaXwOZSDSBNQ+CEjr77mS8WXEiVhx2HL
qRfTH9cGKTf6Mpept/+AuTEu/UZ8C10sUVFB0WdvMOtYkcjG4thbv6o7vsN+e+owLaIaqZ96ZDx8
y7+IG4CPt13E115iHLi/SezDYwrvLV3FcOdLTLjRzon88Vb3+hdtYFBBE0BpVr9rxULdCd4neNQq
ZgCkYs6VoyEBbE2VvWjLZ+Bt1WCSNqvwSKADWTJS7DGNlwpdS6+DHweCWbIS7QsiozIcdbn2KcpY
Le/heHtH7EpSOsH0ed6+brOj8IGhfKbrBjz73cS70zV/plZKYaDzNyvk+Y9J6o21RLen7uy4+nze
tvcYj8cI9mmn97tqrNXLu/TPr+9d3UExAJVnnYb8b5oCef2P/469N3+CSlAlP/EIEjkiTv3Po0rp
xShbYgo7KJwetjOauF8nuypw83BflNepPOpM9xKNFe3imMe7Q3qAof3LtoPN9CqQFoDGkKOBa8K0
sqiOnnBEHMh/hHSqOBqK82P4j5zejPVgiT8KHkk+T7+xmBo8oQ9VAWZlS+ZJDANFCgm69Ru54AD3
UWVwoTaxGMMA4WTmZ+4hVYvJO7cOEudazkPMO4HeML4elzu95WTumpU42xoHR8Ac58EvVqvrYPcC
cD4ct5JO4efNhmofSN0uxP2h05k5Y4z83Ue+1uSWgskz4yNHyOHJC+zq8t1vgG4vo3xx+0krACfw
uPH4bzLTDeqpYSpvIpeBK4L2Ay8N1Dkfno0vi72iKlp1xYPHu5Z5U+Rqx9VbrJ95x7Hl/9frxywk
9qVC4EX+fpsBTu5K1fj4tDmUeeJjCi4ke+xET+J2qDP/L9HJzMhSIRpNPnmSgUIDOL5inB+cs4ap
9JB2KX7zPuuV4vOCbu45p/tKlDK0nkV16Em0CNpKl2AQlXEYmp3pzlr/dbtcaGMhiPzxRGj5r94F
w7qGLjAcxHYSr/4OIWRtx2TWPSiicfsZZF7ppcPOfO+9tczLVWUw9wv8JeYMJSxdN4MCFiKTLwET
nz05/NbvcjqyU+2jllQpJ8Ym6HOn1sFjqwA5NVBnAhxnnwCuL7oegjmvRSS6mZyFcZbmGEzYMxbt
cvqqnWB/ha5T7sEdA0MImjbMmIiT3qn6muU8LA4Oloy7ut4SD3fhqg6SKJqCa62UiQIssW3PJP+Z
C52HNxsYxiJCn3zzQYsM5eZRsM3KYCWyadP1qwKdB04TSaaPoa0i17EFQbnQoF3e7v7tD2oAJ1fR
bH8oaWjsiSMlcMZbOLILKZpmMEOAHB/hux2VuLzlszieTOEGTM5lc38Oju1T48mrl4QdsCYmDZlR
Rjay+rkDs5NE+XsatC8HBxmHJErar2Dtm5v5FhKw69jOC34BcfHZ1S4z4fGzROt8y9hbULyH2y5P
uhphaSixsr1lmF/iHR/Tu0HNoyY5XjxlcUQgE1KeC8JmxzN6MRjsbYMQFfPYUOEbNjskRDhWWWvu
lfsRv2el6RYlc9jj+KUnMuWmXCTlZGrsB9cztSVj46DRbJFO+cEbvOoIdKEzlh/p5LNmyJ2TUkKx
oZmHwQQTPqe203+6cqf0fc5tn4nxQbzVq6KhHCyX5Qm7njdXXzrwGfqoP6Xj4+eLu/NNh1XvGGMR
OIOxnh2LYeBcVj2aKjThNlRagJQPO/FXjuZ3djDb5J5cT+4k68y8df74omNUQCaKQ5f7vW1bv57J
An/t2th777ofm/kYJABO44Yw0AB9LGa9ngvwZvRlHUQjiJfrPgRfZRPXiuOd/egZbq5T8RzHoKlX
OBvETYH0lOjvaZ4bfgYTDX8vzQx8Boeo8Ho0jjUKOMF4fXkXaNhmgtHVr2oGsA5wHHHmy/PHrtkP
WflWEpwTu8aESwh/kq7PoC4FTG0lFwZVFTHRvd3EaZG/bUIUR7Er3NZLtXyzQQf7hjIHYjHiiQVK
JjoZw8nKZNsojzlEsyVM42Vh6S+vRo1GhH6CgeoWBUz3JXQb1Px/OQnFHmQF4Mwj/yUuPhdCOOX2
QSUutgeTMGVB4htvKixm7OBjmniuKpNsYVQ6qsb3wllXjHXoR4ulRbbyI3YPS2GCRymFmSAen6PL
D12ykfvv+/dMHl5hSg9LEOZMzC8wYG8/zL9GM0dlLFw+rD+89RWHwO2ja9WBW/4Htx2fa0ZixLA0
9NDbx0RR092IZ7E50YE4UAVaAfUk96covRLwq/9FaSTGdF46/ZU9Mkl9tqRarOaqmYTLApvwrNcH
9ncJDh2wE2PBq7WKmULEv1dJPLzUiwYzo2vXzpSddeKyJ0IK2KzMYezwjthm755EC0oT11SOeBYD
w4YusD5zg2mJCPl4vtPWTo7Qq2TBEryQjJU+nKlY95jTHFS451EMqi1X66J2pdMgsZ/HlGFFsFsx
TRFLqA7SqwW9uh1yyyzBph2rC0mA+gGnwhT6os8tO5Cm7SjhQC1WcXDCSade6tIFMNTwjqM1FHaj
oJ6XB3+Yf5BLWcUmSbEaSZJc4FcJD5pTHPnhzdf8tlGrnxhXolKESynZ2vsXla5YSyYZZSuHwF39
vmDZSM/M1Q7cVwyfClWSucoZlTpWsFmprA1s3DyElWufOZYHaW3kxFBQyRN0ljWeD4cUw05hOtjX
Rg9b3TsyGygsCl3i/pDzNzif6YWKG2mslEqqC7QlhUA/D5NdhNhy/+++FPOCJDdOAIX3jRlCFWQB
P2t8DrR1K0VKNGdZf3kAWJSUuqEECzbg2WR3CtO8R+7DVYP3t98HBYJARyH8yJMXG+pIjiB4MBky
6eK0lKXVLMq7h0ULiKCDm6OFQVDHoJ+L3/spccCdWmdCw7KTc8XIswmOkPrq0FmKzQHYpUXVeGI/
A4FlYRKCfEiYpTGQj8BY7VP3MrqP4+w9+/hgXBb6pfGj71aE0Vh1pmJVxCxo2/uqLGvECiAT+Q1A
Rtdkvymx6cSigdxAJToKBNxav/bmPddypX1Ucj6A2HMRfFHWx1Vjdyg9VdrBCQRSd06eq1p4PWNS
rmni7ZJbG0WdBQIrk5nEHfeIRY2oSP8pgR8VFFlXfYktBwtDlYYks1FB6eARW+eI0pZq606iXkGy
oxSfw3M03zPJCuzPWCFCwKtUUOXx18HXg8nTCXim5fnvTsqmZELzJ05BeKVZnuRfr3IsWTfIXkA1
tKWYSw1HdC/ODKMD/OptAjQz+EOS1aaIOWWhrigjAF+07JzjunN+CCoO+lELagldPplDG23IUaHQ
SGWnYgk74pNlFMP/4IHto3qdwxR+mwk8JYz6iswXr3RocxEsMna8nckc49WmKZ1IwJBjMXr7O6QR
WheZMENaxoZuLYEsw9gmk7sjK55la/IslKOeJ1ZdX7U3O6OYdmb2VuMDqC7vfgViDlGmKD2ZwRGv
rVqDGJfWBvUTD/5GJMievabFtQo+4SMZmfnMgzA1hOuC49yt4KgdYEbUUm25bsYVxjddQxGKqm2L
VwUkL25EbivljWWfZJR9o+86y/RTR7GbiXIgXOeJ9lwqqTo87vUOddtMCPdtutCiN/ExnMwNdfsN
vLVjMG43yyYQXwNrsfDr9PVgr2YSuOGHXmSl8uFBTTNhOgSgCMZS40JPTGXS0TbguceBchqpZseE
x1CMitcEWWSXisVm1okJ/zANhx3Yd5ruVhEaUqLoEACUzJUCctzUcu60Qn3EmKjNNd35ItaKrM2v
J1F3Oc1KuTHLKgpYyhd833NagIAkMdJ+GeLb2wNHQEvd/ErfYxZuxCxXfAcoM0xsnlbr4kLM70XU
dLIFmUl2rixas8cWeYaEgnQ7aho0jt5aydTB8Iv7q0yVoR+0ISWpf7yMScIA2wOb/mrUUNG6QV0Q
JRhX+tfTcFjJd+GoXB72cCxErKQOwsf+tUDW1w8hPZFS28L1yEInwe++3R2IfC4qIRvvki0qsKTa
cRI2kkPFL7+svY9M3ImceX2EeLzTfAFQh68t8M8ISDAweVvZBe1c/7UpNUlToTOqsNAc6CAO2z/m
XrjmUQYPeieVaPSYk56GgVBVolS+pwtIZJ+zoIW6nnV4EpY9PTY3a3KU58iktMpSWvigHXrAE1AY
jhgb0kf58y+iRyiYJ1zFiRAWg765ewJt20ESgNoysrhr7HrFIK7PtDNfYssEWLN7QOo58sQ9G/cR
svIaW1RfwrgjMCfcO2GncNUhSrHArCDBhFzt+Q+CfBFJTBEFADljzRJjSvwS9LBg7+7KroLjWCA+
5+8oun1mqs79QyHI6LmkTY3+pGkTRrf+WDC7Hsg/Tndcu3oEYV/ZAJ0GaLWMURNVXWL149rAg8sS
XtEaEKcXJHGEWrFGsY9llggGLRYRj3ZbybiAQBWLTnS0q2JS8jjyYtWYLJJmuhwh0FQ8FEtRqwqI
oNJcHSQqAx3bCU1DEQnk0Al6J20fQS7zIv/fS2/EvioSV0wwoz+jdAeSAjKCBWMPuRbFasheG6On
hbOtJI8V9bpZpI+vVVCTJnW2mXsPg0FCaxQ/q584Y3V+kfdpPGf4n60qaQWIcs/WsD+crREJBH/m
E3P1knad6LvexGYh2tSiqyLLxZCfDXqaUwx+FLCFQclC+xR6wV9YydnrDAF5asz3vK4BBAR/pyWH
0Rthd+T9K7pDXCozgh8nI1Kkjnm65AQhASDzWRuFl+Xkz706hnhPeD/aQmu20VtfF0Al2iIMPzid
l3764EFRqTjh4VsdcNaYXqNkhEKaNvl9PQA3nBxrECkv89+RPGwLLEgZCuL/T+dtm4zYePfAkX9F
4h46u0eLKLdYC+TxNS6vKqnnojYUntSKxQJCyTa9UWjW63BgmnCVorOhRxAptWMfLCPWAnXOCtyJ
rbCM8J6FwuP7oKSlmhcZIyVbAoH4hRwHI0n68nlfQanx6cMTjE3g8PHN5kWsaYRSio6pV+mORLe1
wL4xLBaJ0M22X9zJ8sjmL0ehhgq884g3kGJaE6IXSLdJsfZ6BY91Sh803vDVtCPb4eIME01/X5cb
rhV4UTj/p1i2lZ9spKomGzhNMIFcrOsuinXI38/sGg+tOMrZh7d+cT+NVmgxFVZAXE3vLYNmLiK/
Cdj8gsnMdeF/oq8rC5ZDtm+3GnDgMP+aQNanjaIRUYbUpEbQpWU45Ur1DQj0l5wquTMIJh+SJ6vY
0U1rgSzltgppxP6yVJUwyEdJxqMQgQQqEXzqg3src7n4A1xP2ExML/RO2YKaQlszREDhnn6RoJ0B
9NQIhwXwG0fLwUlnF0jWjkC0UwPcyV5ok1rD5+U1KVdBgpecg7NrwdmYet2toMzsDNzDPFHYHVbz
0KA6doJks22AzKWSfuAOmLixq5lYot9VzZP/5WEcFKMmM0c7BaulYuzBue8Nefn/1QE5QrJMYM4D
x6loPY1TCQNkXJ2GwpOH4AK826oHpRnIilb2Q47pJ10VVeZqZSvxWznBJ9aivnmDTzjitQ37JqDv
pQ5K8Lid5WCUjgWsWjyrqJ/JlGS3twq757+pXbHCA39avVn6KhrDBsSMBNUSqMKkf4S0D5IFFdLR
uKmoJqYcBZbYU/tl/+Yg78GelEe1p36xB5mMit3GHSBqEXDWJmuDosouxLYdh2uNAEH7ESCciwZe
OLbaYi6djdzGuFD0znJQ6KW4RyCHp6ZQugXWS+HWi42L9w+Gg50i+1ROavOfi4bd7tloSR5ygept
fmCTWA2DBfFqr0EEbeemF71Swa4aTD0vOwzeyD1uo/XOpqumXg0ZRniUREbeiPfzpqfpptXiq9h4
KApMlPSJZMpAPs2/DAzScNX3PgwiQnpJNNl75rlXWwtfnvSK35+6X/sxMfjZ17Kiv0oXMGkYr9Bt
yJLAD9AEoHMFGgj/FqcdloSHbTNWA1kYYpSDajXInG4IJ97CkYRGgg9VUvfsq21Y3etZkQCNyNB1
cE55shYdmW08itlB2JWOGm8Z8BOZFHBg1uR7WMP0DAUje9PEOoXe3wLUlWpuYsaaFpQMjHfxRNxi
2sj3Tk/aeit72NhBmV9RuI1Z5i6zl524wCi35cxNkSkmjeeaEXNxDFbrumKTLje6kLNFyKmwM/RA
0xqREdF9f4/BV0hVmDu0GE1DQ6MZqNgkQdJekTLrtnoc+kUtGzNw/Y0X8yseQKJ3zLJY2sFGFkt8
NVhA0d+tFUm9M6Un4k0fSCVMBUJNyVEsSCz0oDffrCvh0G7SwZJbJ63OOPeOnFYfN4PwMrwDBtga
ZCHcjo5FCjyyQsWcVXMxBlBwbSC9nJR8VN/1Ah4LhtnhOpcwJsEmEzJetLLdvtK4m337EWCDnklx
2F5emelNwF4ltY2ZUlkvUv9RRU8EEzKGjq/yUopb08FXC0tZDgTPGIl79gG/jrKTTEDvkJDXoFBe
bvijOTYfZSd/A/w9xaQGVV5Ln0KOG7pjMtZU6PRs5J36gApTaYnyunTYp53ffHfkkv98Z7Nu64mi
31n/R4Z2VnFgwPmZNTanAsrEVg9a7RidTHsDMGy+MAOnvj1Xw3vRcV7Nejm+ZJr+rP6200EPvIFM
p4CtKQixTBXVZFlsOmszY1zr4SngMmPjeA7yMMm5XykL77omHwMa3mA6Ry/P2HyWd3hzcjsJrgQY
Rmcm8fNa3YvBV/KLVjaqMrP/xuYXu2KTZASSgP+0WNRge51bEArloaCkl1LuQoDHwFFJtU4tfgwR
gF60+6BqY1hxLlaim63TyDhosSP+LlzrhIoMamozeFey2IKOOE0X5KU4SAh19aW6xzj4L3GzJltz
n/ao3Hdi1ElM8UxJ5xLF1hv0HVg5iETHkNxLuJnfDPQpLP+1NmUddnjHzfqhaj3q2hS1+Z58YnmE
WcgLrcnZCyUrB2ruX6n1bLeMyYDBidZiFLfDhoG3uxAZkzHS1hseauR9bafL+WD6tdbl6cQALw45
Vfw+9nKAVgCGYjOgkfQzsWsfwA95Sh1EaqYxM5jynZbq/JoIGJ+fCfQf2Fk1l8u1kaS6XszmXowe
amSv8hyiReSegeNYOpg5BbIg8JfcOLBRNYnDXsVLw0rJaydVKuD56PLg5R8lgkErbFTDKhyV743A
4GTRZqoCy03swx6YAH96Y12oCX18yjMgu8b4C8xeh5EhRAQdqKoy3aPONiWB1shDYANteRrKOZVR
FBXOK7qkW1Gew1kjHkEl1dd4uv2o7aurbds7/Qa7gjPzSKlg41rYNcAeQKjZYvZaXfEBvlq2ZXAS
cm//iclqseJcidxGFHwDZ1PI9jp+/3KVs/qVUisj0h1DF3hQQaS9FUPa0qzOlQGM0fhDfPkPAb0j
lFj1aU/sBd+1R28KsKFXiuPRqGUNpaKYruk6B0bBk9XAiHaUlw4KGPF5g8tw5Qnp8qMkBwt2yMYG
ept1t782z0DyME6dEYlUauoNSR4984kKir/6LQHLgMWIN/BxESP2d0TuPFq/8VV/JDRDMxn/abQS
Idff8vpPJ8WDKQqWJPwEbvpKfm0J9DXe5GTG6sItWz+wRDawVVDshyBnItjYUXxTxqxP9goCTf2r
vIDY2AY9mE7EGo01ypOUfBLx8I2S+qXLV0gIi7HIIAbno0+JWl4wPTpDXyDFLzDDzQGpGRVfyOLq
6qwsY/vZDEBzpvoPZwwLFFFQ51z0DWozta1nkBq3RWZDj7GlK3ttU1o/TFB9XcUmPYiRHxNAV8yy
8ZMh3Rq/BIBmClMVv+bghwAW9ELvj9S/o+/SRAkaqE+S1uIxxterAystkTKhWJP+l7okRUmEkNJk
g+iQY18SmJlEKupsDZh3DE2CAfQsMtJrlEq4xxHzY1qhLSqV9cnGcH1BTpPYE+3MmCY4UXyAiS8s
uQQxbaBWFPV9d8wMXdgwkivr7etts5bpJIMaf5mgSUlAiiu2yzOUhc3fvX2Eu8Sp92aP/GeKTc+y
ZsLebiel4zaPvtWBkK30kIauzWjfmt22H8Z7kntv6nW/Ll7hMgclmbF70t7XgCeGMk1YIwQHG/fh
TITypJ90MOuBS5hRoh3ZEQQWWo6gN30Rw4fVJFhz9QkddUcdDVgDBSg+XQx9f8JuvmFX4WHKs90U
mrBXyrvl/xaTsLPWm6IYZsGP7J9OX8qvtDdweJ5vu2A2J41ZsMQ6S+jDaLYaVcoP/RSYFk3ct6FS
tvUQb90CN6Q0PDOC3KA1wk23811Q8cY6SXiOtvFN8dX/49qlQRrAAI/4cgjlTTvdMUcZ2KKeZI6N
0BvhHxpw78YoShrlC0diCUoDSfPfMOEhV0zJjZHt3a6Ugkbx4DK/7a71Tty0CgrL3VPwHtQYFy3R
GVX8jLJo39kJVaikb/6waKaB7AyhgQTSG/lUpC2U/JqX4Lc8fls5LAHfHinodgQAFy+9aR82s557
3+mTtVdlLcVyIFwZoJViwuQXYKNQNTveCVt+nIADxRxh2RBlchMzef2oTuBpacQBK5yBxU8zJM5U
iz7f1MttfcvGW1GPjKS3aMpMRMDsdAowHuhNNVGYqYJcnJ2QRSABJqmcbZjDp/nBppOJi1d97kwI
/N8dJf4L4H69UDD8srqSs80KqdrFCQyGtu0damGvXQTVYrPrLPv0mhj0+jgSGiV2YFYbQ8givEQ0
JzasFWSEG8e9gayNlNDMtTUu/kLKSzdD8KBbVfI6HNz+79ESrnodwqaThAyvM7YeoNJ1q6VhMg4p
UXh0opZbUHCAJDdDva7WW4c3FanN1ES7TYwdFJcypiOSQax9QRqx+4TA3dxjGL1S5Rzgrb+BHSQB
r2fhCOMYQ0m2b16JVxtdtvorAPu9xRCmE52SE8EMNYoUgz+hg79IeHW9oC2CZDughkn6rIw5hu2F
eY5bl1Ada8TbeiDs6M9n02p5J6G15ea4/SJtIIDAQxoDGtfKY9FsREOgI96NzFwVF5k26aVKkOig
L4a8ZkK50RONqjr+221330ewDQdnwiDagyKwFI7KeH42VNlIhXojP9StKBdAzKyE1IhQHJVMNT2V
h2DIqhOR3O3q1chXAsfzO/t0vs7RTD23R/Xm7yqNugiyAm8h9cEk/L1qP0BX2eaSKBrTD+FgBpYa
iCR3Q5rHPVFDcQ+j6q41OU0I7oiln9uCEE8j8/OAJFr7PB8is+fpuhJ65npEfcc/6lXaFDT5JDXN
OmqQNwUrARFpKYg/atLbStmbwKQW0iqfKTbPPYwOyncD3oarCgZN8N35IrH36rSBUnJPL1PFqJQn
kbmDPBJ7T4YPtenirpp+RLcRTbiOK4bwZUylBjREE7zOeJ0IKsyn2jpQ2W6mVHnd3DieP2QUG6rL
NcP3sGYAwUA7deshtahQrdkyt1qYw3KKysLt8vJTkcgwf+fOMq4Hc8XcAbYwFg4Yaxs1ZgezdXey
1c87OxPWfJY6VpjZfruaMYLyhpqPMEpOaoOtjQOKJFPXOeqWD8+OJV9Bld31aGMYr6NUPEB+Di3Y
DaGKPSJzV2u7GWyuy7fyKuloO2tl/Z2ym1kkrSQmrvMj/OzM1Dl1wf/dqIjKzPaLA/UiBiNWURMe
uFzvBoCPpI3YnOGND0WUUKBG+1fF4ud2HohR13W3/Cnpd4WlFmz7HkH99D+K39gsCSgBHPxDyLSC
Cv7ym459EdvMWpsZ0Yxg8mkgtWJwDHn/pyPLKhkLCpb4eovgTmGIDaWImnZDiLMmjo0OJArp5ClW
XnjP4CNjMB/ugeLo3w9fbuA2oDrbCXFk3EX7Jb9uZs+5Ru4hu900bjni5Gse8N9jKAjMNmy8hhl5
eXf1NgnymtXe9VlSBO0OXyMzvyTFqMMP2l3xM2ewEAev+v2I3VNiJx0C6UuvsdN0wLN4sLOcvrS6
PITTVunaeF4fW72McHdSUsCLn6AxIPtwGhD24fXZ8ojjY5UgLb3rPrkgUvx74VeWEdnBlBGvsvxz
eaUCebAY7FzYZ3P5pSV6iAMOhgn7XlRasnIfP/dZnsCvWcBL045rdS53YAG5D1mPFYiT9xaPq+65
VI+GTCe+9SDYqooQ7OW++VuBkkRX2bpg26GxVXUZkyoH306pl/b7Pr86QCs5fVa38gsmpgFr2ZuG
A/3KmDrJyxAxacw5q9kd7addI9OltTYJc5GQDUaRdmED8qaHGELyc+qLfNY5sUqXpRN8+qEvJEvb
QGiZ/U2Eq4MmrvN2+aB+RKTaTr+hNibn+b1SUQI7i2vueoLRIyz4kLV54AXyb4hlB+nBw136FqQx
4keyXr6jU07RjRkzv7nzVTzc6LXRNmaBG9F5L4l/5hRDtR2fwDdIJx9jihJM9LOY9qN6kvd5y577
Z/qmjno/h1fWr2s+FLJhg0L8TBBxzfcJ4UxoseO13Zhk+IobHimjhbpRANKJqnyB99IcDraKrq3o
F2aSP2viOmznbUWCITBw/IAs+QNb5JumkS4r5rKGfxaISnUpZ9sVRRIoi2CvmwRf5oHn3rcyc4sI
95Tafe5rzKkI28csYOtMOMDl1ZkbVT1hgg1Q0SjobcuWNoaEZ7B/yMBWz5kyHb2BKAjoVpty00EV
MRcFrTzi0UWOpsPCKJe0HKlKhHhGhZT3l1rfCHBmbfDKefCox1T04g32g7ok/fOjB4usRoOxvG3d
3q2EbTCZ3QerPNsyH7zFG7pTZL+7HzCXM4v8qt55LZ8aStm2xSMGlGwaxNNA0EEsxcEg9aYlUk03
hoS8+4Jg0CAaVHiFfcOYuJ/x+pTNqQ7aCe2z2OH2vabGbIJUsqtPcuaYGKzstgvbTZ99ARLl02pj
85jRVGYBFbuZ666PhhBXHIwslFxbmDwMQdoIHGqEL1w5DSsylg2+UrL9OsQiQuX82GPwAu3uFCkt
a/2OcCY6MGpezLLW4ZmycpYOamnoeccc2OnEb++4RDHB48gwqgmVeIeDfVQuMWayH8kJ7d8S1l3g
ZsETAlwnxn2/O2kAO1llJ9xad7xHX+D9ppW/AwK6U58sJcJIjN0Sx0+Cx5rHUVu4BZqmp9/2SOdK
hNkSXDXLu4/jOznE4pvy0KtqIRlOsnlUglTJHpHcFDC7IFmjdzNHC89BT9A22Xt5IWKfzPeXZ1R0
craaG3XUkbXNfTcxoxzKWUomFgMc1ZiaxsG27MSat4tCU6561Sw+s+T/khWvwLCk6QnEakZGKU2W
d3gk6r29OUBfbyf8IqL0qJLRk2l5d+ZcpND3w7GSkk/EPDY8D84hkaYDyhIrppdzAl5IXeapwv5D
EX/2ama+DY2oXqefXc5tLBYQIcOddeP6/872qXJWpGqO2/6a98ObO6BdWMHTBGxsTUMmPARwtORV
C69HdQY+W5X4E0W8YA7WYkx9nOcEx6/dMullEV0+TDRw6SZPfDqyj22zgb/orvyPRvmIfmpegbvC
1aDYbnnMENo2SG8gF76moOMcyGHCeiHiPEprZ4KnB5eh6WIzhncG0uXETHBInRhnDEHSPUb38tAF
aqrKq7buNXX/B7Uyt1hN/wHkZ6FVyWZK8v1ZsMyFZtrfCdPBMJrIhMNXLm8ieCkB9Ko5neZCXorq
QEjXW7zJK6cwGlP/2LH+8cHlyYiwXR4YZpsqlQ58XbyUEtT/AXA9/gclG2OWbz9X8HmqCUq1+PDm
+b+JncGLS35GjUy/vbUT3vTjCx6G8fjyB3KC6/H5k79tzn5pxRzGVXKglq5Bjoit1QBneRsdcdww
/SFmJwR+dNxPYviW7+S9oLzI4aS+QSZViNHJ6oV7I4vxJ3qF5d5PhawjhW1yBc7SLLU007LNBWBe
PhRX5AHJ6DmcudSTdS97mitV2J4AQLye5qvZUPh7zS9EoRQIxwxjm5YZFU6/HhljnUIRmi3ZEqeH
+rt2KhYfsbdKD8qVZW3z/tigU0mBszxT3iN/UJ3Gxa1eiGRqnAcyPZBLfdlVcmlsInfyNUOCFfX9
gwaBJfn2bANodf51NrjGC1Jb8MNUib70rFom8EuS6X6Zlm9yoQaEDWgAtztMWIB9UZ83qba1fLf4
zWLG8OfgQ5kxJXZLpg/WF1SJMXMG6Q9+QX3hHSGiOK0RLmehgBc2kBxaB3vtO1LAuQojW+4wGehr
bREJSASo5fAZrPvAj3muO9giA+0ULis7GsBwM8hghpnVPtuddF9ij1IK6EBdfFaqZlcUae47ogCW
RTDKodUwQ+tFm5XyT9vSVqsHyebo/GN20l3B2fhdVh36unIBia7fmnLq0O7mymHMcrwNJQx49RF2
SZzykbBp3lZr8taBi6ngGfrwMQ9v58QoU/89p1vH4OvcyxDdkL42hD3n8v1d/TPsX0DJ8P7RMyzF
zTLlgwYCDUnNn9OzIfomKFh3VcrPXmcgC7XcZuzvsA2rV6mbHKaHbj+BzqalpXOjbfhndWAXX6vQ
FMmp5Wps+RUuLKR/XZ95dzc9jk7CxFKEf5S2aP/ZL9Auo9032jxEiYrMXfsIoDhduf0phc3BeCtb
rkV21OFhTjUVg6+JCWcph6cAO9wt+2sXz4mxL6/vV36MSyvbxVeJonqS1aczA3UYev0tNHGYxUw2
zSYcXMK7Ww0YaUyfRP8Ftqk3MftXB1lDJGB5sYqj+0Ha7XISZD7frwesbiBMD/nF9fEg2UjE69lO
czHWubSaUw45pUmpazAY6/qI8zpGScZBASxhTRsQgi5EgcIrzyop2SOyg7DQg2plUePLajfYiB/J
TpJKLPxIuuZ+DxbSAecfgJcJ+u0+9v9k1/+OJaug+l+JYmYlgntlSasefYA5ZM23LmkzP2YDDKqV
TsSV/7pSy9PzBrrIe1AFUxuBexWwyjmEGhEwlgxIpp+QedgCF5JfSxXOWArT3MwP58+5F/NYBPmN
NM7ttVImRr5VIFHMO9Dw6azQjAoauPuXy08bjy4Y3PIRNKHBPriM/csMfVATs61mxFslc4Eu/fxK
5kWvIpSEEcqQNruJ7q+gdgHH57AuHDIvny5GV+Df6Ff0RkV73U6wyFTM0H6EFo05LUxHbde3dZbR
Xqw4vS1IagNYcbP1SoMN4SfZvuBsBquGAA0Q6A3ss+Arg7HRjYOUts8h6v0lQKYS3J2EvyML5J1O
sMQK7UEK6F+xGeoUrtkZsl7DX6xWrP91QC0Y2rwMnYq97nP0QDdG9QmzjHmufx/1cjE3m2158boJ
Hi1WxbeGwaKqAqlRIn5IRfeHWS7ZXf7ng1+KN6hkky44LYjwKPng03OoDEffJXjXiRSRcdvUo79r
WibGIPpT9hWYsiCmNXthfMWaUBwLeizW/1nYI4pkDYD2kEXj+pwN6XP/G1Uq/rPmh49ftHu/4mLw
FuT3UTwQZ+SNctMbjBH/gUjuM54MnqD2P8Zjt1pvA3vMTyP6jaBz+QVmuEVOIFIAKeefgHcG+l17
OjpVB4r3+C4gFyq48n4jfbVfLHbBcOyGnnSKeeO20/4ZFWwK/ErYDuZjgwL2tNA04gsyzgfoJdyO
B5FFM3q6IbcOcKNcONPyWf3L18upxSUQGs8Hefss9mP2eIWtIFzXzBgKIjG1YOgTe5oz1CwpzcZU
K60wQKYvNlXhSe5snx6bckyDZZ/HqHgUfbDKS2RE5TeoFA/lsIgAauvZ96wSnoXn4beQaTJ75HO7
yDsw8immvLnM36RhyO253f0HUi22KXOF/Iaa25avEC3P6PpDS98B9GIFTaw3y5JD9W+kvgYdkf01
UCcGuiS/nCGe/nDsNM7OspqGiDmajIDxMGEEeWd6Ep5EmJuxQlYFAH/XM8Z7QJSJosLpyEXHPgMi
wnUkfciup9ESJamjTItHRMh7nGVkb2GaaaAdTFv9B1Grxa0zFc8r3HsYgqHijUVFskUOPTTQm+D0
PjoeBAuJvmeqNicWB/04FdVUTXrQmWgbsF6OSFV6s/rIdbJbcKZ875a4S6DOiu4pNvyAfIym/qud
MkrvMS/1jjGaDGy3RtfrC0/fTXkWg50rpXDUzXsraJPV1FiLz05ZMhfFGO+qFz/dfbwBlrPHGgxi
4jJoAOuPsE48El6iODYxrCR884L2OXW+9QUPk8XtmC41aUnt5QK5Al1L3EFhjlkzh4MSmAThXa0D
9OWQJMZRpbrUs71ue/Epq/EggzB5rrPGzltxbh423OvVVDko6QSRbjFMGZS2vPw3e27PbUYJGX33
AkNn+TKP84lp0xT009ROuO9imiZxD4LJ4IsOFftEacoTcMeHpWF0kGLkqzjXKElP523hOZt9eKos
IChOehItwS2/FjVa8m1/EQznlomvdCsPo5cXzimWJ8xAP0Ft4Itg+WZwbIG5g8w9S0CRqRW1DQ7I
L36Egp1uE8eEswbzQDnefLHcLWpHL8LtaHZ0t5D2FaDFZjtS0WuOUGMkEx3euvN5HXiH8lQeX5A8
O4YX6sR2qOT2ZftzpaxxxspZJbdIihGKvg4NdjlorVRuPtypMELzN3+TRzEqKmHMrXfFZzbT8K2p
IdAusBi/OxcZSlkYdraYVlPS8969Oii+4ABrWV7wsInv/zV+WT6hACr2rJ2VsVRxh4aodDOJqjWE
qN5NHLHlrNuEPtcM/jCkD8jKBEm+v50zlAKZjSnyj6SZf0+9bIMj9EU/GRpWXBsDfxeM5LwcYpfH
Hw9ZFA9XUuSMGsdfsF+9dKFkbv1lodG6ljsuIweqEoSCnQOdxmMJJIDHm0rKFYtZ2DGf9mskeYKn
EDCarJbjnbgd5sGOITfSa3TFsErcer04RMtdPCdqeeaw2ylNuNYUZvDkz6V5MElHjBaB2Lw3gSLS
NPA6BNaRHq8YmG5v5CCC43DahVdKIsePdHNZOf59p/k6SV6U5+ikAx1A5i6hscLgAjdAwf9gIqBP
9mPbheSdZWOHq1nU/KT7/nmQLQe37zrJgOQutH89KP3kOOd75reEBPM2TY4hAssU/XMYToszPyl0
Ym8zTLLo90JR/rUzXfkRQlaz72GgNWO7LLMIsvGaGWNqV8cQ6CYy/qgfwbygGjAx+h+vHfJLcodm
sN6dN084ZLd5e8vXX/GcEuxDh2tLm3QhG9mZOElXHKk7xerX/RmQo2dULlwZApK7d6r92ZEPTJzp
CF7PM/nuEeLs+I85CKW+doubgW6+m7jcY6qwXoJgEy0vB6bSzfpwtgsgx4CCjtu/PwwgR8G6JnB5
Z8lt2tJ9rxfzsI/Pz4WzlJvfjgrRgkuz2y9uks7MQidooYsaxze+72wulsQOoPjXBkXq1vPsv4KL
GFPtkFfVe4cb6HCjICWkQLa69WuvYJs0egrRV2X1GozgBI2U5kVu7+gHe2wequgvLzxQalEdB112
DF8Rvdq8jUgMr/li9iV5LYLUZyonVJJDBuFE0HSs+tQBrZbGJmiOknciAD6yX1nTwg6SfsiGhgyo
ImWsWkjExsaNVEWfEUcA5dk9Yly6O5zTzZVzZMuKprgd+sQPwx4DzEr58mXcw+DERv9NHoQhy+D1
PsHDSbviXpcRTf9ExwFDp30vtw5C68r5QwuKaNmAyRrljLtD/xqdA8iJtl4qSKfe0ZGL1eTNATvk
Nn54OK/je5qnG2KTsXqh+sq9lzwOJExdbhg7KXmxZCfUOhjXHsGn9+M2cYGrfnrEGK9Y8v8I3G1I
GNWT++BfnFS48dQtFsVmmdesS+v15GUi+QFNaE5eK2KhHB1N98Ph85QWP993NhIZHgzPFuNBAquN
TOtifmNalfBgU+PvuT2eaRG9xP9jL994LrSbt/ZOVtBm2/wLmgssfsM1m5XdslkV5jUmpsA+UrnM
rgFy8jKAhFQ8dKz2pebIMhbTm7VxJ078PsJGYPEHkbiwKlcnDD8miq6hB7yYJ/0k7DtYAAiwR6Ws
odPe9xPwA6W7IFFZimIgMtoNpiF8N9s7CtvbhUTBqIQO57+TpP6MpjjmnANMEuhNEK/z/6wa/wrV
DjmxMgS87VQdJ19eJamvu01Ez2ea0J1sPBpNADoztl3NhuFs3SHIZTqM1AeGV6srhyK7CpD5jlbN
Fy0ruBIh8MLzWICUZafVZEaaG226l8D5XFyBtAkVzuOh5f040pxGasQwrFUjWc5c6u3WiQj1vZw7
ldf5ng6sAReRUsVhN1GlHYB2QycS5Dxjp9Ixo/9ChPDPSnwA0/0Z1sJRRVekK1goyuReNyfAmVk5
870oOMf565gZKz8LgUX+PBqMp1EyjDOuid6ItV834+iCNyadLzXbiMWZPO0SxdaPlywHdzkMcp8Y
Yj9JgpVEE7q0XD1qEFgFGVZ80AuXxnNb2174h0P+Jay9jxXWRMTMBAImsrqqCWk4yQZQTsjgQ7mV
JtmsljBN4vsSIvpKemFT4VGzOyVASrzfU7RmsJ3axWtePeQhzwgRs0eDMuYLVUZ6YJor9cdLufMZ
/D546O12gz3RBX6Y3CTIHeWQXmkqav5nDUzwBzqLg98uIC+EWcEwnP+YVJyez0Cge1pPmauBBTcE
q2kIGn3cbO97X9wzeQJqPyvBgCZElP+SshxnUoOv3G+dRrDfNaiLWqjnbMGgEouIII8L8GEifjG0
agh/EeSUVVzzcsMtoMLGMj5qiFsQJuyqGGiFzL13i2exLSbnN8bMRbStvvFhfB9I2ZTtFiRQeoxR
U9BKEXLpHqYOhlcTkihSEE9hoK34ucPjPJLQNfqxmezAEa6/rpw47nV+XykJCPskAQPYFUV62E1w
zK4FZyZ/x3xknTqqjC0SVikTUj9wiTPutePANnakv7eJpUaCgNdRUgz2VhuId7Fk/wAiZO97/fxt
wPa9+gWIoVmACbHYytS7YZ/yjpHvqQoawGKhZIvGfQ0rc7Sz1LFYhbFSLjo5HwVwYqNkHmukbFfK
rKJEYkhxQne36TJF8NqP9KomUYpRsln/T+9tQ/uwy+i3m56DsC3l3ui8vsjc/H5R0f1uYghFjLgY
DnLIfWr1jwWK8yQEpfQWDDGLfusA8nOeeWfjbRQaWEcz6lt+rvTSP63FGZ7KgW914yrTE6pe+4k6
JRvffAdkVh855TbZK1ozK7WeplC8K1nKZZIVbwG38U9PTtvaH5V0VDkZwxLvhd6ZPXfKAsDYLITS
iB1F0zL1B1irdgwlFPjoi4iugvyGHaEbjcjhldIn9BSwJWTA1y/ooer00Ne6P9OaOuvYBxD3mRBp
p0Pw8cVnG50XdxG82wjEdQnQohjbVc2FdF8vO/NIgNUcu/jRidZbgcw2en0mO938CYZJcSHK4kDX
Sz7wV0v+eHnkcmkTN+1Fu30obwFWnG3afLnIjoWHlPY4KGR8uw1IZD87bhvwpldvIUCEB1hH9tNg
wZxziOF6tu/U6OYtX6FSn4tGnlT5Dqh4GH756kVmXEXMSn+UjEdAXzc9lHNJ/GbdKwlWaWoTjiG2
WU8ZVivAb/FRFbfQ4KofBkaPCu4UQJg9eAISjhnAqNaN5CuWBtHpBEHXMt95Tk3oFZmSnbJpyCoE
/2f54lxKvc421/MT2XfnNZnElKx1Ms5/cyMcxN8oVu4kUE/WHmVVsAQvVsRPs84n8sqSaAk+2naI
pF3uK1FlEkUdsic0ZcsZ9DZeOpefrEMxY3bGhUaSQ7YP+fuiq4HlRbPz7udqYWJaiI4xLVRGEFKY
tZOzVUhXWngLl/tl76TxlF7hYtEdMTEyHXFV5TXCqKzrMjY+2LbR8M74n6tmCdJKlT3Md8sCNJXU
C0jS2rIL76hcNoGlU5049mF+13KakL+4mDGqkR0ETjeNX9ZzykaBeMcgOSAOu7nJLsUP9QG3Yfeu
gkQb7ynFPmx2EQfDHBdFzftd212Rp9NRKNkFGHEJnQA2fqdj+fnNnEUzr/9MuzQxxNbL+wxxd4hD
Ua9qhbXbuMSRoHAM5O8GmoBLc8psWws2ffEE2QNRhFufA7oWrU8vYLw9MrE7xwZdQi8TNwFjse2/
/dlJen1rNG13AOqS504Qj75DsFgpNVJ9bdsRORGQo07aPbrAODKxzQyheF2QiLQqFCohlMJxbTPf
4jdRhjjTwPV3VN7NfHgNzBqeSfjpsEQok6ERZXeaTTtVe8XtOeTujd9cRtNzCMUgYE4P/j1vzpW3
GeCSaIkur8+lDApHrQhsotesmkOZMbcc8Nbu1kT8PKB65sAifQw2OBVRaSYhxF2rWyq9OYRv6mER
p9Ssx5uKYtmNVJrQSeC/qIFrV4Utmh/+G+25oKwSnuyihe57LUvefHDNrD6Q3TjhzyCNTzmCBk3Z
cAw4sQEQ2eZ7QgEX7lydtzaPdK/Go5dX6RdQDXEGBmTnHdf5q7iPNvblXQ5WyCDocp5Xncmv1Ua8
X2YMo589BYPEdg41UvoMd9nV9A4DU8QI1g2U5Ks/GSP7SkP6FvRIfaILXhyXZs8+Yeq/sX8DAjEv
KFNTWTVE0/sgEtPhtOaP1WHsP4DwBbN5kAXR2HN/r2KkD/If7t7CPDQccaQmbNwkkhQeM1tJdNm5
hn4HmaGx2Pfe+Uc2xVgY8ADYmZw5rSneHU9rEKcZtM7kEbY2fe32CI1Xdn3VTPz+7KgPqOJd9cp5
ExHmrYZExxnlzt9Uk8Jqij8/ZYny94I+7CMf0jyWIdY9pE6Q+XMZhiwx3d8nezVN5/fq+HWVvOUB
h/zm7WjcfZVdSVwCDtRrQJoElrgFCEf4iFx1XDN8VR1aNtEjspTz5xWYyOvbMCCQrMPgziddKftM
lg4fgMqG/1j3tz9sBVciQhniigOElY1RK2S8BFBwMJs0nWzqf0YnF1U04jXsqCtUZHMBX8ujjIa4
D+8RKvmR5tLWVvJhpkGwGEqfkY2onhcHjuKo1GEwmhZfg5OhOePmuZSzAuYbfdObslamdLc4hsuD
EZOdtEajYLX44jMfaHXDddqssPaxwSFnZaym0+Wbyhp8/rtduZIA0EgPDEQsuy59DGFtZmbmrwzv
hrI2HgHwVGp/gVl2XaXtFsWttWbtKHjhlDDpTcrIKv7L5Omb4CgwgJmK7p+bujMmUicWgJBbH1SB
0/BRJjYIyfFYZwfue98acWf1BcF7Mus0MO64JRLR5SGuuiRhpKr77a1uv3FigBz7lU682YrOv3jC
ckI49NA2Et5RDoyxBO24t8X94YPtlCLZdMyaauzYbTM2zKO16o+PGDVLZ36O9URSc6A49vSd9nyy
HPGGQiOkzG3dZ/0f6YvUc0mBR4aB+QvwUlvalNHE1rfOjC86rkf3jhSxrnyr41Jt+cqp6yfiY1/1
GZaym5V5v+Xuo+qdyrSfvgM6bziTi4Y/o1DKUr3XsGt2UmOlF9DLmIuIrsJGaysuOSEw0c2wC/W0
bw1y7Ht+DB4I3Hv4npC6Wl2Wrz/w3k+AsYOKpyPY540g1I5XWWATjruPMgC33SNuFB/9BISj4ffT
oFdkO71YoYcYWNidaoNlF30Fp0W8D6VUkueWwdauQHdk0KI+TBZXjwrhk0WvuiQeWwezW/Hd6KSl
QCP5rpfXuZWPs/Rztw9SRXGbToYBdnTVlkeHTn4HxrYGOFANbtJbbBGF7J7riFXvaWbasv6W9ABM
1T0z7op/ysxW0GQB08Zw7GJpsE4nIhhPdCmDaYJvnTfl3AkGSguidH0SZbUD2wiBBKlUtg4sE42B
euNdr79olv5knLS4gorEHHL8Ha9FTXD25hBU+RE23B09nm5RKavJmjC1eraMEos3fvFlF1fWMbAg
rdZyzx5Ue40r9pEvb7AnrPfAl/pGYg+Xye9o3UApkS39NnbNGy1MDYb8XTRqMVBOAvXFDznwuMW5
M0n5gkJpsOAcPGeGFXw3P73Ld4IM5iHPAp164lsw1JDFSNdrVYs8Yb97IXZj7rOMIYBK/PHDhfNA
0oz//PIzcwSOXc0Agv+wiz/ckpUjCZo7D6y2H5ow+z8Ubao94gbKbbD2ewZdUV+sT1tHbTlCsmSD
u9Qq3vgqxx7OREQwg+K5WZTGzB7/TI1NwmdlbVgl/nGGVsEytq9xZV1cbPBznsaOEEG2bszzCBuI
LKG6zoNX9JATNWNGmk2aKXWNVXUx40nBCicZPOE3FSSN1ybLpPKbZwkkFY9k7bz0HQH8zkpV77OB
8TTDklRTrfux/yQQS6ZG/75/R9zWItNtizXXiM1uOcVlCVppYKoHIo2kG9aDHvUfl2KHcSjbw6ci
rLnIIFWuagcpcEaJMy8HdoclQDdz2h/2IibcW02xEFdMV96VbEJqi9OHrrHoigNBfXmsG+Wl3nbW
gzQn3qq9h7ZDBZhbJSc3OytsRXZwZ98OOXjasdLLd3IlAwMOLiRNwRrk/GgYCu4DbFx0bJlXZZ6W
siB7AJ1qMXEU1CQUW6DOBge3zejgKjeiGVaPPAKD7NQjIYsGkFMOENEAysVswBXr//pCgEEZrPxj
rLZ/pfWToyfHL5w044X4FTEvEERerAPoa6Md5GkH/01TzJf+h579D4L4bf7MXBbz4+DSzyWSW+7W
PCfcgBe+ygGQZ8nCBvFfeqqPhxGAgA4PjUbVMgLYuZQCb2tmD1qo0jfC8t4x2azj5ow26biB44By
ptK7eC+Z+llaNpIs9q6Y84NGjlTYtzJ1zqNa1pm9mC9iPWMvDn+SNwPfnyo/zCrPBpEfBajVCqnE
CTMEGmi1+aBx13HxEe8hlZNbY1vdnfg3aAD/vTy5NUj+KJosdqTUjPejCHuiG9fDVIGm1/2W4wjB
PMxbtLrxFbLCx68K63R00W9xMnurCrAdkHgq/i18rUjlrVCInP20RM8jISP87hquu3yRT4sUjHad
gwdG0xKsCGbcoaSRdvrXfYJRty+JC19LzcM3IB3XuByvM2ZJ1OWmPI6uL3oze1h5ULl7IgjaH8K9
dzDKlAOBTbCRmmxkT5gJ5NiaEtJ0GG7vPnGutL6r7DXLXm1PIHfa2JgmjgDbdilcV+NHVhT6bTbY
Za5Wxh36MmEJXs5zoBarrS/uUBcEdlfSbLtw2TDi1/QVSGgjGt6HlIDwuct1wEI2fq1l74iAnOHq
o46cnilW7C9k7MB/Sn6oOfhkIEJSYrcdVl69rAo+/hYoX5Ihhc4zQ0gp99qBHm24cDZHN+sQjoUB
4sejYLL8iz2jB/V2lqiaRCHD2CiuCOZVpMPMu9UIyEMJ9sWrLGpqbmT4tg5J1u4CLxx3/vvJhrFp
3qrKXQhis20a9ARzp7BF9s987jF91iZx8PP8qn5VzmmL3MFkhVXfA51Ock5niz+sD174mMl7NhND
ofvPkrvA066gYaotxhJU+ozfT00qFwNzR8DfH9WphM8pAyZDpOl0HHVY8xKZkpPBl1+y8+jUThY4
pS/KUNT5+ja32Prfrmhihf7unNi7l4Aeq7dOhTyse8IhLdCT47wzd7VGcDXqBFSQY+te/RMVQE51
BtwReYs7WhFP0ozsgSlItXBU1ywC4CpwD/PZUhDvngM8hmLuVqcay6XqHGREogV/hxIk9AG067jK
Nx0sNLnlo9c2eDUny/XNymZZOclFQT6SlLyv8X2MhLGYb0jnLsi54MR417FRbZmnZ5/cCHTEyxlH
DaT5gNI3lDY1CeXj2pULByMCfBfoAg1BDZLy9qkI7O6ecaKOLxApvjGGe3dIqX5TJUljNnPo+0H2
jBqfckG4GGFdBagUismIv/01CONQiOFeFossDfYhxE+MISVynLXX8ifTt8spxDj+lcj3s6/i7LXo
OEnIYge9Xf963ycam0e2uYcoEGfz9w9swqIogZnKYb3TA/NNEB7ynOHs2HK0G6IMa4QSaD48Ss/E
Qjr424Gc1N2FdASDfw1iHOTvNvMvsSZyEdYip2iN4XaqlefaJdNjbhxzW8p+RaheV20Kw2u0xooG
EFuE14LuQ+NM4kq2O8fh4RCAsWHb8L2/ah3gn5mwoZqFDS47GRLp/06lTllaubCUfhmi8seX6Cuo
CsstCjyw8MlE5kfolzrxwnh7txB4f8I4gY6HDlWpAXkN5L03zBgaiB73Y5SomfliV+tEJv432d6H
p/rnx8KuxrD5MT+KRZlorFRssqij3Z51lLdEyxtkSTaNarPzAX4G18Ma6MMF8rI4ek/YpFK47muy
Qq6R9Q5p8jUNdmH6T/DyctLVElt/xORH2GYWoxGBdsrVYk2g+NtSEFeJmgpord+mmOXOgxY5hWYR
6DxhtAXa1TH3Wdriy6PzZlEgTJAdJoSPwC4sEOt0bw8Si20W9g41zJF54q/GhAqGbAd/yrgmt7zg
jzyHajngafHGtp7+IzqCS3EpscObX7WshPfEWH3kD0ceOaancSiVB0vpdNqPljyAJybUOXBs3yPc
sb6OBFHqhSTNIVoEemddqsL56vaLoW8oD3KM+cuc4dqv1IPvReZTRYdM2qbN+qNfsoj88rjqua/2
fBja45xVdfNAFGiTuVav9QtDEXnWAKVJUTE1L57U1R16DlSVYd2OkhIYw8cM9jEHCVhpsFlpBlxs
ojo2urltPwHIVPb/68sbLFB7sHMfbCX45iakUOuk1seXgkXbDkTRzgYlJiUaaF04XDEx0jBs0hnp
sdGwsaStc+hujNToK1h/5w4dYubmA6jz9X9KVgCuw0bD9MBGchpLeUSW8HyunowM68WUOJtimc+u
nAeaK/Ki4aBHcf5vHinPcao6mBtRI2tyNFUlSYeH8BzxyE4+ECCFpOkvPG+1CJty04idKE8W0r82
ExjrxjsRTOEIens6b6RYM+hDs5ov7MjpoSRdXKjVqwF5Br0eTZRmAFvHM3bfQEBrL53o0YZUUEjf
olno9yzjc4dL+UakNTQPV+74EcCOTHkQp0nTgBBpR+okLSFTqziqcdJwS5gr7S+TTFW9AosGGK8+
SmPG/Zs03aqFv3tTMRepTIw2lU1CTPjF1EtXqP5kKMsbE9waxYxyKMRu46GWEfkLn4Zq/mYmUyl5
IcbuDUz7LpgkM6Av7LJ3EJHJ8IsD1BIDzioVZyMQKzIwU6I00J/HG+ikJu81Y205p9t33EIqHXpG
sY3jcrVu6kqUkTL0DYMbo/vNsnlWiItSm3CcW0h7IJjhsA8XSTstCMF6jlDqjXFJneIEob7NRHKQ
Nsxgt3fI36cw3nfw/C/jTpBbjXUdYi451mb7PHOdiYkjuw09zxcINQmlxbGVpNLIn1qp/wgUKa6k
4v9qxiaYQl9R63krVbFGi/+cq9mY9gTTKG4OTsHFDT+GkbUivnK/8gvs28osiZ8ZczeDznQQQps/
Hp+OMMxXIGblM4YNBKRFnD3n/c9WuJ1QgrY9hvmrMXbSvUR3hPx6P28VuI/apZsBGiqHKjfaQdW8
TvOz3t50vxOp1ZM7PkMnYBoNz1u3kEfL1AB+QiI04PpxilmmQFKgO+ykchQPre83Q0zUY/7K2px4
usOK2gGJYSXoSUalcjvCB7St+bHYMcM3VCE8FscISBlQZpSAQ3N9Yl1lhiG1J/hHppa0Zf0d/F6j
QtmGGX5WFaLRXT+e+tTcrrr26deB6/bL4OUSapuDE5S9XJQctdeVRSjPMu8taoUUo8qYx31sGDGh
2nP1QxqaGW6V+m+MHlEHjoK7uFkM5642K5IFXJcgbaIfHhyrfUQSpJjEMWvQjBie2P976NmLa4mV
dksWqbiQco2IIysQCv2joPcMRUZKBTbZnEAukFdWvBNOOHjCxAP0Vb5+It4ast1AuUvmUPj2IK+3
wzSwOy+paxFWBX8LQ4gmKcN6+J4XZXiftmcDqOHAehm/p6C+zhRHS9PGOHCUdW+e+Po8B6h0XOM6
KUyXIHdC+B/UAgr7eVqxxjIEsdWldDoovZyHHRfNW+OBUibffbNeTzlXnOfy6SkYpBhBHqHZgVLB
x2kR4lc0Q3BWxu44pQzUes5sR4TLnV/e54uE3PEbajY/WxmgKjBkioqiZvyRfp7AL7fNFkHQ/KCV
aT4N67yLkUqIft/S3HXS5rq4D3nIodw2E/zQRduhojBeyxA++OCEATfSEjsjvsxyH2rEC0yt+BGZ
HQNPTmjE5GmLzYKbCYsiGP9emORdGWlB41rxRlKYRw4EIM5Z+VWeQIA3iKYVX6F9yQS0ps+maMjY
0jdEMY+oaShvaeGWKADNM48P6kTaDTqVUq/0TZqgEcbcvowEGmkzyu5jwVZXRPiWB5/lEMozah1g
RaQFIs4nMahu36Tc1jn2qM11Bcxwsnq8M6z2S1JklkqDSxIH5V/o+xbS5/snlyDWO4/E8nHuS+RZ
V98GZntjtFWcvTi6LZrzWxV/bBYJJe3/BtnT+QgLT8AfUXJDP8qY5Vv8bYn1+0Cy6qZiOlj90nSZ
yqyIcwdPM5nFr3ucofplJd2WDW+hz4GjAOZoiImiSgIEQ80lqZYuDvpI5oHjlrl56O7z+6rD3ZZH
7pJxKULlyLwzYnAYOfStvo/yg4eKv4Jg00r/IuyRz+p2EbsoXPtqrEyUrS7k+Q4yef4uhX44jsQI
8B6rQKPClRRNTWRl5nCKyFPeECXiXNxIwNu7ZWZE+gVR9g2a/lQTgIPgom6K0rDasqnk2Bqba3He
Gr3O1pRvvCFqZPl6waQ00IGQG++NuB2y11reylrkV4RJ8RbnKbM3urcvMHVqu19fv+SRpXOIB6it
KJCtnQQR9ZHMhOLxFkoEngITD6tan7Y87lG2hF6Htwi9+x/RwvHMEy+vDhZdNFKmpPWdR8t1hMXv
H+WK4Z4irvua7ratCUAi2g1nNcvWmu0pwIyWaiorWpiTEIvNm0xXuPUPUOsFU2PgGUwFzsaVYKpF
rcT/KLMrqSk3SLVCm5IHWp43w2pip9qkht3aJYGld5Wx0LkxrdXnTbuibFXvXr9oDeckbAfq65QQ
Poq06DMHrLat/w3Wq4KUjwqDewnjYRMRm1m6EFiZLKEYoAoyv8I94QobG2M3Fgniy59xJIiLSGE9
bT1aPNgbRr5tB1weLaRjXS00V6gECSlGZ1vTU8W43o/76/eox8j+9AWonPIWLJ/rKO5mFHBYmk7y
zcwVNH0FK3k9oqPK5CHJI6NH5/fbdZAFs7WVuWHfGjPwtidLb7nv0opie/tX27xtSwIj4592DyIA
6KzvsalJHTpKMvWxDkG8BzvefaTqbq18gWqrACHO++v1zBblsGG4Ir3YLM3yYM9NmaVFz46XMyXB
HfI9O1XqR6sN8TFbO2VSqzP+Njwc3asPPaQ6SQk2A6ZluiXAG16OyPAd22XUrIqxzzqL1ysreM3y
j67zSYOnTWYvLihELIGgbEyn9zuJmHQrykNmiUFKFn/JpxqvEi+7h1rCHs+99kVh698qV7kNNYJJ
JX43Kn7hV7xxOwS3Fo1keUQy9BoM0LXS3IKRWB3AA4Zt54vcatecaXTt++orTBIvcPactjjgahnr
1IZzSu26WUqd5HpCuZdms7d2Fzcu5fwgEL6TEo5k+SI76nY12rHuh8VdB+X3KPqmnxC1bE+gHI4t
Yz92w8wI2eIdS3Qk3rYCVG99JUJYVzg0+dM7EkDc9nmPmizkrZE/yGqDXxXTJyAhAn+i1H4BR4pv
L9UqGZJVVJyFrXWezRogPGnye7Wad/SyUhOtYOd7w0e8mrcSu9ueiuFWoIXnU7XKc/dtP0f1+3vA
JTgkCt09UkvMHZTxoewKqylBGaaNPc80pX/3vuAyR3yvnAUD9ugpVR51Jxh6pvi9ku9jl9sGlmLz
RJ6RVOclNrm4P1bGN157Si0IG9oJqmCdYBTyILy55okgsrNfDjeKQDOkCkJCTQhkPJzBusyLHyn6
kedFgegMdL2iGHaKTyV3hgx7ZYGWpd7gz+yYxbP7W7hOulMOm2wEkR0UB92lRQLsBrH6hC8u0TUX
wYhdZuT0bm9PY6Cai/2kaofwyFHIiouPyUQJoL+0cEgpoW+DePpk+1Yo1biGJc+rdHWJCL6XzS5c
89OvWDH4bTaxqMnGWKu6xFmevmX0FlIjgeCvkYL/3NjIlS1kawbQoUVrD4/L9UTJJTY6+LZKGIl+
/tfMyfVzL3wtP8Xk8Uc4xn1SwDoRVgsvroQYmzOeNSZVH2ihRvSGIjTmLa7n0TZf+NjggxTN0ApW
kSLnHv4LkZaTwa1oi2jMFew8g8vvg1/yIoXwXe3bQ0W/fTXqvxcZLN7NuMbU0suM3wYLhrubCsBP
15h/vPlkSPBxXaKsUP2leuTdqthEa/HpwtHV0TXW3en0eFouNG8wy6+Q8+UvZ0XElo5260l47DX9
01hZijIIEYqxigq56FE2kjGy6RTUGTNVV+/kgDkEVVcN1q0/8Vj7uR6tVsE+cyROdhdl4tp/wE+B
hDnCuXDmIJpmsqaeZj+Cb7HsrXtS/xxlBsOxjTY1hZwkAOCPRtP2Jt7mV8nU6KvhRsKm0swf/NAC
bBEZp3KwbPPHCpmCaZUXYvjwqB/OZiK3pJBq4Zhs1hva3ml0ueBGEI4ovRd51V/RosaOk9GiM+UW
yI7tyfZTvEOoR6N2WACVEiWivoCi+oN26BUd2pQEGKBVfqqV4raQrdSD9dxZlBlyPIFaVAOstVkl
J/WDIafSN/hl+TtRtwDCifoPK6Rb9hXaJjhPmbBNT7dFYJCByRdEPz55Qj+6JPTAoNKoSkex+nDN
BKrujmWZpxClGfhSCQgpIz+SRgTlkLRgmy/H8Igr61jNyMlxlurAtEJE94+GnZekwai3RUFB+V1g
qQmEUg8Txj17DMoaQF1PKzF04t4pYIBl9D+nn3MgW3RyOXZvT0ueF2/hIPgtNKfvxMK6mXrCefvg
vQuiFNuu8ZaC4xgeXH4BEVJUcfsWHH4YReOu65y/DxWBVg8+j1/6q2QHouT8raFBBDugz8ww59mx
JNeZuQBsPU39qaeeSNMb+Lfjr1SirpwSrQJoo+a1K4nY8S9GRZqeCQfrUWW+i9G6p5IG1mK1L9X8
jd59QhwL+FatjCg4jk0XlqIydS2bUY43nVNXKlq5jJi7yzzg3lLnnl/DlnwqzJL06wBw5yxL27+t
LMUTcTKqpTRk6gjzvu3H3YUad9nGd6BeTM2lV+SaBPrbQPGFKjF+80iNTHhmHTiYS2Exi54Z2miJ
QhaS9NjwaYhvHmsJFXQ59Iu9MZOKNfvMppCWtPRZwmSdhXV6im2ihC0ihdyTJNwBgHU0lt7mCKqf
S966BLFhc1PCagltbEpbAB29dZce6fiXh8NQOsep39RveXc8XH66aYvph3tKVTGL2h6gmFv/unRK
kffV3tvp/ndugTC1nZ97GvbrNl+SP8OSHiDa4n/LluLr+1NRucEAx32hoeVkIu+ZcxsU6rvy6uMr
QT0FbmrPe3JqSWSSuZEKReFoS59rW0oSszGVkT+YYA8+FRsaSEBQBwzaZYCib7IVe9+iruFCcK4A
RGtEjdcQjRoqxSvhWOrtOpM816fCj45Ywin/+zhJRt/zcCAy8qq3TcdBk+HYcxPyWIJVbet8gwoV
5lzw5rOrryqZ0RFwyOFvjrIyr/XuDMZfaJ4PJrfiv5E3/vSDVEbqM21+dKvrGYZcM2KTOtGigHmy
pyP36yygNpi1yHqIHVjhH/5HNn7kHRwqSZC2PY32ewBGgeN3epVGEPMQFsUQ5hyV6oEs7EWmnEpC
nO0bbazvwkHioCY2DI9gEa6BdkfNitS9LvuR0h0bzPzizHcKsVr5VIuvljvUJ6wlf/cnvHGldEh6
BUdl6Vn8P9Csr/rwa0oK+9Xu8cNp7dunj2ks+KG72rJlw4kfsifsWtrn0EmUSvQKRRG3pahP30ym
S1RYV+AzoDOXHWh7CEUltGHeKMZCpm5eE9C57oVxG7z2qqNG1HXpKkCaVOHIKIS5LXgI9RBRi9mv
vq2wB/W02bB0pO6uiIqpnBUyGOlPHGeH9otYNPryzJT9Nr1hyQtDCsAyPSJyfF2CWo2Rb/J28tQ3
SlusVGIt4qsuVkzYgIYUW/Br0Vejnbo8x0Ja+QBLEfr7L8kNtNrDdC7u61/i95Gv1AQ2CySf6RI4
zUj45SCh7CmxvYFl9rrczeMI2k8fJWjXrG//QQYnrErjGMIIUF+fvRnBk1E3qfTSYty2O2VwQ9eg
tkFkDi6GhmwLt0jm90yasK+WoQb6lMEEbyjj+e6lEW8Pw9I+diGFUa+5SD5GA6ZQKXcltBAy+cPZ
oJdma/H2EzoBQjyjrkWcA5LVuhKU3JW4IgltnNpn8wtio+I7kZwcEmQd+6wkrh1/7I6hpYaGdP0z
ONYWqBaRVMShFR1p3LuOy03h2GVA/cMoZ3K/6RWrs+Uim7bZsCi6oeiTqAFV8zEMFq5p7qR6ETZm
5vZw/f+tKmQsxHVZXwZMy3YgeMQkC9rxN4qQFJ/0fTwAaBfiGHk8uCut0/blHBwW0H5fJNvevy/W
sSHqA5BuasG6jgsZ1xR4x5ftUrSHUEtfQMc4Zo7AW14madL7D569bHTGKUgaIaLkQ29AlJW8g3pN
pLOQ7w6W8eePubEsTd3FOpSY9kMEqtD/00BgDuKmIjJWxG6HV1w4t4alMwOjlSz9RWtffbG2gYbL
F9PgdfuUFyGUOPS2hfzN4nstg+vnTapu8Sex1MVdyIZeGKB775wz0duWXi7fkId9WpK0n0Lli5fD
+fImCJl7Cqwpxcq4zBvlbFX1qLuaq6K7CjgpzGHX79NZb57grOMyBAkNW8Z2bqqazTfQkbebXp6v
oqhvVxQlv3ZCiFKfSyCBT10LswAtT3XLme/d0v4VffBoNdIVHookXMcRPyRD13S2KBe8qWdB5/Ze
xIY08etZeZ+yoNCCgWYbLZ6pvYzKO7SD+xPLmjDKNMlsK2nURlyJdX2VziIiaVT0KefNI2wlXtb4
HKbRDi2QJdTWVVeC02h7LLGbIIRrZ+YBROZmmjf6VD+IUFrGybgTJO/vtlRoDnRUotzYmcLYYDG6
cYeAC3t37I9H1PYlWKTShj6BECqnmbg9CyTrww7hpc4T89ktTWtB0heYDHa1jMXo/neKZDXZz4YK
qa0vda+s9bXuATf83ll/K7oqIPWuasTiG3IuiTQbVBc60R4GagyNysrQ3uSFTlQIzbC+o396Iq1g
O15kcZozFjx1CKz+nnRvTbYtqLcLenBhMRcTRlKG7y2nHutrnz7hwr/wE2SkNKSTPsLcl2TiYp8d
tlKufVirTg5X3AFL98kVqeBxjFc0fEW/3kUGjOd+z4loS7nNdk9mhUFiXZAf5C27HwvNvCBJVdWs
KcmgFiaPqHJRSc9JSS+OnUv3BgVfFamj5ocxbLiC7nf9XbWwhFsB2HUgrcXrf++Dd3xjNGGhUZYU
A85cht9pOlMquOjj6ZgpO8orXKZjC6hxe8lv0HPPvJyPt/gR4P4aSbSNz709zZnMqNrdosKnzhN2
yJLEZJbn0U4AWn8Wm5fMFeTlYS+nTr8oTZsgVG011w9vKeBGZIVKz8D72XLJDTO+H0fOAoEI2JRM
iGbuiXrUKV/S/pDHNPUYIeGa8PVsruHGATb8N+6vqS64VDJqBrO/QYhSIcymgHYuQ5yr3m1xgKag
BzfGzYWeUn3N9wz814+a2DRawc/lQ6Om7OqybmqfxAh6x+kjUgpyAx36H7MYkXWfA2+QIdQtzGNn
2cEzvzHh75HLEbAa+GG4A5l298+FQNUcfdUgxcCr8mfbEIc+/pQPZfdn+JKlB3nPKPdQT3tPn8rP
xTJZ0HGpo4YLI+tSehkJ4Xl4QJK37RNlsWDpsoZUaSmT9abyx4D8OqA6roiEbqJJjpci0shBJQ9K
2uA258jwPLcAzzVuF4gsY5CPc/QG9Z1M1iG2IUApS012yJ1/US3Fo+J5GP47+h+hq9tHPXzCmSw+
jvjeiXcfzRLBXNQ4Qci9qY/vGAYRJhglpxYULVLcZcoBi8h1AzbdPGuTfr7O4GzymHB1yVaUeJgl
do3NxnYTZdxbWvHQSrgJq8oIUXmDjncXTyrVwH7RvW5edHSpJvdIiN3woqbjNR/N//yNO8tfGNVs
ZPNwylWjlrVU9PPSWADPIi6ZiKGhIJ8ZuS2EHytx0GQqvDNGjah2Mwda8QwLjWPnYbBXiyCHu2Js
B0VxDNgTRtdXNTct8vv60tx7u0lU8g6j+1DWYNUDJefAQ6iTAUPLosERknfax76DLFxjvKVCtTWI
p5Ki8pUQjhFMgVHUWEG71K2S68qBHoylBSZ2Kg1tLXdBdrrT+DP4+SjstvD/5snogPcXhaJjn1zM
WL2NQMKpR+MfHJd5SF5PN8aHesca9dyjo+HUjREgM/n/dSCccn5fxF+mNSbksXgCrLusA/n/V3ox
qVMzLkDw9IYltcnI9vTD+FGb7dlm+iaEUObKWNGJz3jKy/PfP9LyYe2CaO1EH3p+L+BVkIP+Sq2u
n21eLpLnPAVN6jPBpAVC90xH3BruawWRDxeEsLYBowefsCYvAZNXlk/KKkbdHo9Jyeoe1KmNiSg9
V/MQQ/hPQkGOG/ZpSw5ayuXDJeMefnZll5Galquu8GW6M8NgmnArXyVCwAbn0h3+nVSIrVSm3RWz
Eqfrd/xuaMxphVyzWo5FnjRNhPJVlKmRSYWbSo9EmoGXFJz8DsEjAh4GVsafDLo/L6UgG945DOzZ
56LUqFCazVjZ5hb+oMHM68CBHNjlAV3+6hUeHUFIXFehimWt2HvqeC3ZZOgAMKUBpiHUegVOmabq
extexBYVgU57taUc/hkGHivGE0/6nN+FOpeeFVoOaQNRghtpadNxA7/ViEEac5uBdiNzfSKJdcTn
WNyJ+dDPswKEbeo1EpTYvlEp2oLPfiuWJBdGS6p2c6YzbmdzCVHhKQ5lwAwTmMxHzL/at+FE2sv9
efsIs2Lqlau4bj42ApgBvP0dXxjEpfjKCTAZWCB3gUmI/S3scJJyUfq5OJr/xrO/d2j6LUCwJxQW
xVQKKafoBY3QYlist8lF/NRv+zjfwbK1U6iMjr7SMiUruvjcftiKrzIRJm8cY2wseSEr+DEMt23B
E513bZuYMinQjwm4lepWt65IlGKvU5ZiuQcFfZsFNJvW9MBr2w7cdI1ATPhNVYDeAy/7Xa6YkLQ5
eZrxFnKohU+/bDCpHuCeXBmCHXnUwVsQh3yp0PVJPaxCT7O4u5wzOPfW/tz4phYoSbNPPMZwUKS/
Gkyt8Olq7K36PbHnHJ9+UI6PAFwY1peENKwZJNuOOEYwvaNDZxOmG/0hEJdkxcks/p+/KzoIDcR6
EvB2GbuinAQseb51ZQKG6P71HTiCtSLBQRvgeB3ukqGEvEIbhCFO5q9iaxHcbL92QHfPht5WmRc1
nouhaE8kXQ5T/2vqnwjy5Pbc2+UriJSd/jJdOLqCTEETT+L70UesYc2DPW2DUn/gBscrtmTlUkkc
sZPtnLpW8kNw504FYzIHnu27eX5YEwrlfUmUsjOX3egijICHl/Am53fhAH50mOYdInel1k2CKG9B
74D6+7RyEd3M1bFSSSTSuodDTJ9Yf2pT/pLnzxsZpRw4jhqa/hDItnXHLIvYPI7E9M3J/EhOzvRF
19tNQlevQGDyRiBMDkFXDDHOoJX7P0RBb4/+jUtO04MgfZgQknnmyD4uyCi6l1K8YZXsJbTllA2D
mN7jNKZwk7tgEBTJy1A5GSH/gOiyCB0KJ818kpXIcY52caoiLozfunn9vDG2RGSdy1H+foveOPTM
vaijljvdaoRmKtvrIo64qzZnSDb11xIFnNFLoWaG2AgTUXx2eO7CwCWBa6Q3WVQl6jkyfQA+2/+6
/p5CXDtXwwmjV2Rwi3Q0hB27y6Hknj0m/fgziSXMgtYq8nADuNU3rJSU1dyXHhmkjFo8UTZOnnL3
wddPoQclnElqq15+gcDOZdtdu4jE2EiHZ4bsDfXf5IC40qAQksXeKSOvEtcZ+eUD3Ae80DD+9iDV
5hptIDCEh1G+X528WOuQdvLHuoa+GnGzJ4CUtIHIRB/w2Fko5HYirIEagWzRzQRml5UNZamrZ/B9
hy9WJONR/7QBOetFa6Xn2pU4Mc1rE1hN6GwdaGBMZhHIPx7BN171VVL1Y+nEXO2Nuq8qe1hrnC9J
sy//X79YwQpA5pmCLzY9eCdCqUJCZxCx4pqsZKR5qNOWQ0xSs8HWZ6k/QIBA7qrTzBB+eB2G+moZ
HPoMbhZuuNFQXXE0igoOUwoRDnbuYMvdEBYeVw8syhhufJP8QewjA7ixnnzEX0IAj3pJFwKgtBk8
9RpA3KnEZMeUPKG0NhwcrCLNx21Tn82fZayozBG1g8n1wJnmkdWlMx4TJ5YBHutuBis3D7Cuuf14
apLtgP2VHHTJLZfFeDUAnnpfZXeogwKFhK1zzhtrlpvVLbHVRM2DvmwOydsWvcUDK0jgYWd3PRA3
o2ZHR79NH7NQUWZkmBzwdgUzbL3WH/rIMPvmHYXBowThZOeiLuzh+kAzB4wzLJZ5utev0/CehALD
m+1XvtKrD7t+BT1peUuLtCpvUKO8UAqTM8puhLTzTh4mzUpIMusk8U+Bb/bgU4AD/EkMTB+qPmxU
kva9YDgkDWYsoCnk2nuXxCaR7nVO08asdOpN6zSvGdswxO73BXN57nneMTG+bFEPUz4LnyUkR6z4
qI4yS3CM+CBekHB77guyl95Q5ClRNt8M3VuQsGthYg/K0NZt/DoumvQdnlW2UWk6G2b+yGcYqxBh
2u+/BAeVmftJBXz10zooUrNYVw99AVFs1tj1nXH8bjojjBIfF15AGl53htfIU93h7yEa2tGzzceF
r/LOjGlkMptAReZm4s7ax74T4eqPf5QWBPjkYai3gp944zmOErvGp1qSE5yXnOIjKs1vvCQEfOiO
Jn0+HIifKx4VekprkS8ArNrWJsDPOdJZGsKShd7NYKJkh/c4X6sNpPiT5O/emld97JEtInCLG/ja
abDYKTjwuCJHH3jCVvNYcfRwi1x8TRKrGJ3vzVpkEAysMNZaTIL7TPoyhIzckgeChjdiL3CHJiJ4
sRRBk+lNPE+bFoXSnPRFeJv5dtGZ/S6d7fkrobekoEsyAXMf54LzugF19z5TfbaPBxRIHHY28GOH
W3Tfdy+IdSkKKgmFTXBAX5ZQubHvz7EFEvVxMn8NrjfS2ju77Rh5p1nW8+DeRsZKhGR3y/Yegmiu
4fB/uLuECoxbS4/G6UQ5lJG0GL2wQ+MFPegqF4wraibKsxyE7gjBqlpQX+phnyV6UfPVqul0U6kP
y3xw5Fpk3be+n2Fvn2ufEQf02hMvbA6XFxKqFtKnG/eEAThjXaVhgQmTWdsMn/ZvVyPlFWsD/R2i
G9c8EWfHxubNaZWT/BCgYHZtkUITTIPQNXQvareW5SykosCYj74Zzc2SSMbfqH2xuMVMltsDH6I2
wODms8qFLjPtwTE1kzNvgn+38rKIJKHtsP8K1NB81rK4UfCuAo9QGGCjIhfoWa+uXzmEaeFLwp69
+hkZ95jyEvSfRPQL2l86URIUXNnLeOIZ2J+T0ryx5I0kGMQCHL8Del7Zm0NL2tnMOVpwB/d+UHd/
PBtGZ6TNJpZo/2l/NpV63Suol5o+iw88weRtNlbu/CL3zuKDEq/1EnAD8gbM85Sr2kGYx2DrJo3Q
7/zrgZfvigT0bZT0TJelXUwXOmOPGRsWQdWGcfC4V4YkOg1yLpsxFPm/Zv3UlnfnahX9uFpvArpk
qRN2xHzf1NiLBvFWMkTJqfl0V7UyiXvWEgV9JPCgYC3f2JbPhu2Ah44YdMW1DIRRQWhd6WqdGwFD
rkzMnVxwKqnhyA/0zCLlyeOvDf3BiTX9MfNRys50vaBSf41PUXTH/9T0f9dr94OahK4MkwiLBL+T
CL24GYdQXn+s2MtxxLba0ntKDJMkik5sV1xUdiAfG23b0vTzliS1NVzKidyEyhwXbQDApSo5FkJj
r+P7bk3LbgqV4r6rOrTJWBTC4tbGeY48nhEa6MOQnLFjBYpEe9laF0KJ9qD/1hd8H/92zzzQ+BOr
zf1y3ptJ3j9FIteV8RG+wKQh7tTo3i2J3sLAX5D4gyCAs34/CerDBtpKeqmrllI9mGM3L/GHdiKo
84Bmv90raIDEuCkDvRlXyXLDRuwI3XmgZqkKQvvKjO2OcjUTpBJpXqPD2YMhGLOgbxCxwI4vhmzL
U+k/drX7NBjUG44lBursfBPIfOp2oCnZmLUrPqWqp3Cm149UEJTT0OMrVH9gBmv2eCXpXkCTrsJ8
xeU2/8rtPdkvzEitJmyA2x5dRpae6sigPVQQmbrAVRKonhu2781NK6znvq0NsAJW5JQf9YaDdGpA
2r1ERHVE8FgKbVW9HExPRihxHBAIEQallrvIy3uxcjVsrBIqTF49gUV9UgiVHtZnFRVmUjQtI0pd
hZBDCxBXeqHBPFle0IPigzZ4NEA8FcTiiRvvcqp8PCvKsJBliZqvBZPYD4kAiJPzRFXV7CzMnplB
ARwmt4/XFhyE1OwNlTM1UGxgnMNrUGaubP5LAIVbmrXw5mMv+zZAubPYtG1pOoW09w7ULfgnFr9O
S7gk/9cmwZ1nsoW+gdhbOwg7JIgd4RLO3eq+pDG7pCMQCnis9JN+IGmiX6UtCLwtn2zTgKXLAqVF
kL5yPV55dqZ3zBTrzxwOxywr+Gpq/kgR/KUka8/1yUcum7TQKeqGEjrwSHupeTGQUHJRxuBvpGY5
jOpWNDXebrsa68uWEfLVoQOgpzFITIuGjDX2869neALvaXvjJf1DW6xU0lM3aKidhTP55i1WWXng
5Tvw8+tqkEunr+3UV8k2PHbJIClfu9aI3jwmK12CBrwYNdDY6iMSl1DQNTbvzGEBZZKS1daAaCFu
OaFAeL8gYbkkaW/x+eWUMFXDVlLmB5nhkohTgZiHGVxTfBy0OlqOwrQfQk6xZ5Rsvx78aLilGsY8
id8OJjD/Xlh7juQUvJAatioEUBmJJx2qt79Eikk5TVoJs3PKNKWBUGp7FllkALzTWiLN4AFIMPB2
wEl79vRtGxnNNBa/04zjMOr4ZaWIUV5mA0EYH++viZ7LhnusOy/uDim/qocFiLagfQLm0MJGnNpn
s5Gm8menlkWvB5tTKXctqTofnMg2SvFeM/QFddHkignR8JjjlQ7EgCpcogHqeuY1ZhRd87+etLnY
w9VqvOGoy0uMNlqyrg4ckFPpxlASRCD0LkPS+VYZ5nN/2ektGc8ZdkhPoTUUWzDmLrcfY8f4upR2
P99Sq0aUBLvnERI3iHjgACnsEhwZoCLQa2e1n9sy2/ts3nRo5SanStcqCYISSyUBaJhpxJa6gzg7
c5QKCycYwN3L7QJiWAzVIj7l2mVubjuFvMT36ChZMhDjOVCcudtogEywjT+KyALFNIkHIo55Lh3C
yirpSJnfOXzPjSixWDgRxQCdY1xxjlc0MPBfeX8EZQB8YIMQXEIcLLUZcU0mgl4+O5qfcmHvYNyC
p6nCJNvrX/8GVH/PFuNaI212PTHYFEb9hdM7Biu4jxVF68TT5nGy+dvlSv4ZwZz1AOBWgU1FxgJW
M6gMDCzZPyIZ+rthtwqz9vDd+OIKsdOi11j2smUNdYlm5hVWAwtPgViMeJ5EzCInhBm2xRjltMiH
rDwWcMKDYI/lp/dHzAMiZvV3LDv+Jh+Mk2Au6e4FE+H78Lm8tLGFsNH8KRf86JZy9QhHDCbQEhfA
A0Thsp5w8a8zqpVIUJrKbeb8T8w9yO0gBGjNfOza54PwinLxd0FOWt8JztwCP2qTzCpxSp/2ZuPc
iovY9hmd+UNIOd2Lb0K6I23wozm/Zlbf+zxPFnZTttZl+9+jJ8XULAqtTotFgpFzp/NYiU2zcm5C
3MOmG+RNqDKfpW+aT8ZJgB8QhOxnnV8PK50prNzizhuQ5kWNXnYcGtcQg4TjaAooTBSBFEiTzJaG
h4EvxzenvSmaMAEfP04Ws6iCrxHrrnihsDXUhIAYlmzYdsOuYboN31HsDlHsHNbksm6NhHDt9yZb
Fg1hM39ea50mmmNm0rw8kLgcS7wqWBBhKWFt7x261rZVGbtTawgRtaXfz+w+D4BRP/Ny/XBctUAm
0/9ICTRZqU+lsLIWYPRVjTNPucjaRf2NlLj/0fTWKRMtV0i3uNb9a9GUomOTQcwiN2U6Rcz9Ojg+
ZEu+IQpOuY5RbmBJPodkm1U+ahLnnSpdU8cOrYUe18tcQNuUS81dHJ4EwBnrof0kYWa94jBS7vJz
q15JbtriDGJjbS3/Bf0kqxerSo+0k71GV03bAFwAwHjG6AsAK7Z6sCnjbankGaroOABL5zTtgvSb
4ZA7nxXcxwHfImiFtqCzHzXPEyPLrTKwI0NrP/g48FRjqSu9/7XwHoBbPpRfj6s4UzR47PTVxVd1
uo/tEhqX2Mqje+1A3HCDfZBzAnU1yLRnb7MVXL/N7HrNIXV67IIkUPsZBG0mK1dX5ND8dAVTl317
BVTmYnZwQD5CMe0uUvZnwO+dvQhOb79SlROSZEcP3wb9LmS5bXuOrmpB+3ty233Fe+I2c91eDtKd
9o85djD/T12z2MWljFoR9zB3mrN+aAi6vnkMcs9mixJ0Qkwk0YcE4JhBqfJk0/cNMqHWpc0RRKdo
pmxKMlcVwkJsnWCAQS5HGnGWEks2RmWMhw3VtFz1d1+8YxThH4nO3e87QGyE41P52nwJED8BRA5i
636jpme9vFlklSmQjl5q8tMzzmd8QgHOj/k7Q/cT6ypeUdXBj4crj5+px5KP5Snq8/UfEMK+CHXC
MxfGQcjLXlSg1lNaErxF6F4elSQJbShDHHdHTNXDZyrJyFypS3Je035nlaPmLmFx6UAI4u/Kf3vD
6/4bgMkWtLlU0Pxlv75bLdM7zhBTl9fMM05wOEBbjWjPQr84FuPhAC7D791a2+zw+h0a2BEgvJ64
2DSIe1gejNr4LmTCZRxhShDrD0ju5TQl7sFTGfoqpc5ma/tdnZoBdHTa1AJT9dT6/fixH7OSOsOP
kD23a9WBeKshfHPgOK456m4GQdM/u2frK61gVY3Y09nfcJcREBUihL0B3ZylymVP6jYNQ3Nfzo1v
Poxi1oMw+x9U3HY9V3x/OThnFWrBCwILDt8Q2ZeY0pUalJNUEuEeXqY4cjnsoB3RLY7CtjC5vZ8g
RhxjB348JfUvvrGEB3SQd/sbDLbxqY5syYySKOj2fhsbQQlBQQdczkaKY4w9ggczUzH+wB+fvw8G
fOOdbwOZ0D2VPIqNrX1B/EyKqfDk9ODRRiYd3Ko8Y303gcZQeOqgLgCu2JkcHpcLdcshgbBUS4wS
4mFI/39RN7chdPrGx+qqpqJ068Oxj0GlTlf1WP4WUQp4mOklIiaMl7/3i5AESKDxPfVsCNMcH4jS
CTqXf2KEwdjsZ1cSBt7xwmHRC4jV6b1BgMejXTDH8zcrszpdlFSV/lHrF5Apehmn4csMPWYYj7eY
h6rLjyejIzL9w35n3gGbHzz80RY5nc9ftHH2ffR1DCSNsQ69dL/9vu7UjUpV1Im5M/AeGiJq/j0l
HVskXm9I82emQo+RVbRrQmMNihRHVwVpys6+gRqqLV6evn8zwAaMwpXr3V9fzKndlgs33aLHviSZ
vPQuurQSLivPDwSwayUlUt5wIxA8hnYEQDfULTJoNF/lQoN3/9CXSdW9qAzgKbo/c8IwNzX7rxqv
ne5QVDKaaOVcAdwiB3uKpKEv4S9F/QW5G3wkb3aBnfxQf+ARvV5Vbs4YOzwW/c2eS61/FT0uua5Q
Vc5hWiLeaB4UpKlLQ3w0mWS1S4RrtM3XJkUWzvWdzN2IlcFqs8GqoMsOg+Mk27+We7ykFLp28T4b
wlK0QECOWlygjv+dDIZswlRjZcbcHj68+d1On2TWkkfXcqLryCCWJuzwpNXXAwYzMsHhLun4wcY/
EwXFuy+HoGgyScB+w0r4SNKMHdim5t+5JfgsV6uP4VDVjU/KPi+OABlD7RpkGwU/GVPEcfEYIijA
7UoMHN2TZpSSRakVsDkdiDQrWMFP529G5gek4gg33NBBNmASX4Ao4wKLBmCiRRGNc86Wnti2NxQx
oqZXfxvGiS6TCeIPMaqCRN4GvY4uA6qw3HOisO7cfhjM6g3CnhMTIjVML3tz5H8cK20Xvom+F12b
alYqCLLLzzHIJwDS4yyjpxkwh+fPsuj1iEFBcxlDjyIrHpd9Q8afoKPAKzU1tXM0toOYTCrwxwiP
AsgAatzfUQ/+dRZ83vO+HhG0NU+tU85/rmrVoem08eoanQWvjG3XPAjf+fpFS4ZWg0wT38fA1Tr3
TDzMdU3OlQQYodJEYcddoTaSvS/FybnlFp20+eWlrjcr4GAIghDUp9kq+KWVq6fTm9FhW89BKGzq
l2aEIQtm1T0+qDu+7/8E6jSY/aBDRz3HKo06meW/o0B0gaaiMignyHWzr0J78jEYhRhg6EX/wdRJ
l9LasNHaC3MbIf+4ThZLModDjVavnuQ5pgo79iQ9kVTBR1ew9bMpIkZrEcHEsuBlSquDkKFyjaK8
gT+ZTmxPLW7MeyKcW2g0P0dmVFyuqIXMZGcVFLY4UpDB1o6vdRCt46XwpcJMPoz9+TPXlCxcD+qq
IYUMkJlt+1TwRnQ6BHsuyy7bTvXWmneBMqjniqN/ryr69cWMEOnLd0xmIoDODFvEGia7+A9FmpFR
sk+rRSTn5QpzBe1+46qTbtZMeQ2qAFaYSdI1b8SNp5tzIuf7Wpv2N+08ogiWS/4FBft/gPywbvoB
K0xSE4ZNPDF6dmiIId/A6ZwJphVIgI33ej96QrsUKBqTPpsGBk+4QMruJG/D7mV6/QMfH0/KKyZH
jCgVb5LxrHQ5rcYu5j2443EN+wKkqOgapvAUS6vN5pXmgouKbzhlYDT6x2F4pFqtCs6iIBxN/4VH
Uld0QMHot7STa1zp80Klfh0yw0oMUeNpqwIymwNMmmcKoloYKTX26Y3Nuqdcd+kkTz533FwX9a25
6/E/C2i5kaIXhNd1p+1a8cmFfjXtUoOJ6ozHEL0mKNJueRUNo41n6JNdtVD/izBBLz+4uos+q1CQ
ugE3WqC5bZIGojJHbZzKMkzfwvd4jU9ksii1OBJ9i+8VgnVQ9vvgKVQtelGj692vNdf4xvacSz4B
u335zuSXMHrhNoU//YcIrcbMEgzagn9C5gbqOYVFibR7hpcAfT/45a8jejl9M0/uXAPnJ5T79XUJ
V2WldSlg0CCMDl0JrLgn32jaBPFb+GqKPqn/CVuFPNTaDcnJKQS7aBaHprFi6CVfMFcZOrGzj2yf
utYnjWjVOtGZ73kU76LR53YbryBmOm64GfgGg83tAoqIex2euEOG5B60QuKHIWBJuH3ot5Zxz35S
m4Ohtlx97K0AOLIPZwnyp3h+0QytMRjAidEB1LECvOlyxkHYIVMbOrG1B+r4k/vgXZ10Wmbi7l3E
LUPapPQj1vhLyjw6oWPO8sxgO8buQmPQUFF+GBFwREnmQYXvp+lHo5QbvSEBf8DX36kZbbTDVMap
Zspt2lp07hCd3YTqEm2hhX3Vk1gN6mmqG8QPCnwQ0iK917VpUFkUd/zk5GeXoMx6IjZgm5uXq71M
2qvCDvwbdAuOJ93KmsIP2+196Nrr82IaGdSVyhWZXbKT3x+Mjay7sa2H9max5bhdd9fK4sl7Vuqh
VrYU62+5wv6mjYbrYi75AvwienXRjPF7ngtfJO7ZqWunPdajvDKFkGdfMTRyN5T8QKC8PDhJx+0N
WwO0z5WK9V1GetpTi2Emvn7hpg9zon4nsRbgK3i7F0KFw3+2VmAKxMERv8loD3Bf6T6NiQ15fAZk
ZQ+BtJ8sB3lQm30+77+xwwCumqeE1gEksMUEdUOj/PlEeyOnlrIvWC4hya4C9mFDRy0Qx9lXyjBY
cinAkfaiMGoNQRn5aaSYihvzapy6Kv9/HLPPcwMe3tbJsM6DbU89oI9iHDYt+UDpAdGUlok/6/Aq
g4byx4arXEDkviFZ/kBQ69Uct2M4dGcA69bwFEqhXDngVCzliYfqSw3qbrUMOHbdMJ95xXuc6Yua
EaAgFVMN0ri5okjt83W/UbcScRRKLzmOLZza15iLrQQw3tsKiu/s/JrchiJMDzKRmCY6Kv+kvbCU
+Zd9xQ5tOSsj4bb0VG6ghjIo2MMy51UN+Bk9QVGwptaXsaN0JYRO+VC8VulANEJukEWUyqT9Oqz1
hiPmfCcKzKfh9FrNDjzQLkqTufsG71rYj9HozxIqJJdcGNicB/AXynpGsZxSWjLdnoqv03QqsJob
V6DU/G0wGsxXxFxtPi4SjBGOZHtMrgc5hIkYJL1ZGYjpZk4bCLzT7VgNmbUbl6bqSfmEJ8NLO2Im
jiO1J31YB3WBgd4dcMWR7NJexpPnsz6zLMgI1PNYVxOKCz5uOKeaduzY0hu8gPpDh6FTGG3p9qsq
5WJeaMQq58qFY8hjkFhXUC/7FwhDnkD1kzw+gNYcgeNSODq6zUuheKVLWNPawUGL7qfbfshH0vY4
/sqMunWiT/xbvzwecsE5vJl9BMsMqmcYX+HWEbPR62gncE2wW9iNNa2loXXXzUn4/ZvdQvcg30DX
pn6qS5GPi/Feuhfd5C/5Dd96SrrlGPMiATuYPfFFyq6D8vQeDdkzWWtbQNnRzwKiU6Z4m3E7bG5l
hdr8UN38DJuvUtZl0VthaDyQsSa9AcZiWIGPZcl6lx8zfUjlfxlFUoU+TNX32Kj0xrWspf7WZjYF
hpHJ2p4YC/vRa0Z5fu25oTnrYAzdLSKVsCudP9iRRKc2VxJbCCaBmtwaftSbVfN8eSdgSW/ny8SR
9pOBz/64vv0YVVSpIONkEOotjIyXiyKpBq5uD3ZQ5F6NBLzMNkpkAZDDgkyV6T7KGgw3q/OkaWei
PDOxiQ9XZdC72D59nVgAXOiunBFX0zAIVFUCVVxwa7MMXSGOc4yVhzohPzLraaVNV2cxYuuxrNvY
TwSKpAmOGec/jUYDKiL+/w8YU5x1oo1+f8iNww2fUykLxG0bNKqYpcoiwRBdS7Sdhht6ICEU6fOX
OlXcijEFJE8JX7NeeBiG+bI+LcMYVR33A7Avga5zSk/3QCHbbSpu7bhLan4WGlcIqJ6CWrEb00yc
hMvUOFmA2TiLaDH/vHPkw4+f3BRPJZtHFkDNjQ+8JLmUkMGuCN3P8agzdhseTdcHKHXzA7QDP94C
vF2P9ZBjwhc49UG3fFjEgZiW80Vq5sBET4uoeJscOk9VT2tLcO8bYHNDLHMt8ShKtbOBUV9QtWTz
8DT8ljdzNudvm1D/boFAgPHihI1PxjyFJUK/8KQIXCqcEPshmBh+lEFM7yYQYqDcKvBoIvPl7+jE
9USStrbOWcPEetGtt+Y0DF9mXe275p29FGbNXcby6YoeKrseiAHRV13Nh2fLNCermjGyVqD++IhX
D6N8mp1AulWUlac+/6gpnQDmjmZGu4dKHImvxssOd38GyLKtj4yqBc1rLQts8o9/3hK99LggdLts
OYBdK0Xl+Gd4QKH3ymBnsKr/q7hnj9laApo+mwXrjVDzJkDAwlcBapdzZWDb7lpqZi9T5IbfXFPp
Jo6slaPZ5MIR1EotLUvfipqAkLQxYvsEmUjH94WxyRLl0ZTsO1hWolHTEVrwiiDDJUBYbLIY5WUr
pwid+9b97z/3OAxgS5D185tkHgfgvqKohax1Yy+PiR0PF9Sm7q/rdVufjBLXZlEpsF/Xeb0e5CrX
iAeZWRcR5XsPGmJExkhGrQw8R0PwpgP3Qq6C9yeDY/gB+1xNC/XZuTf2CYMWsvg0Vd88rLeIhxMr
cEXNSYgV/+QFt06EczcFjCI8xog/twVtQYT3Fc8Ek3ebpq+FXVVQt6GgYQ9jgi0Ve6iFq3gRmRcA
LU/Bt8CK1JxC0oOiPvDkDlqdXnMyV/Tnf9IcKOb8nYnWx4CIj+ke1SeLWzGGVnAv1sQAv/EZu0Sw
/OHimtC0d6paJkk7SaGun6kPgBLEZgF/iCGl5K7lkuYr51L3NAoho9D/vB13h4+QwPxpX9dppdYR
y0GnfMbTEFAI5lWCyBHCKcc/Rt57dlBx/NUNhExFA35YbACl3EiOGEgdrz4bvg2UtxE6D6tJef/3
Lr5N9W1jMhK2sh01CGOTV9WUUEYUvmFCV8vrEC+i9V6ogDVdTZvDjIOny6sa8rnyFSdCjgMCG59d
IaEC/MQ19ZuL0mh68VhO3lelggwA2bIku4gIdBw47Tsl53S9K9+zINy+d/CaLS2T4tBqU2ORC+0+
OTtQk4IZTNBhHmisoyhlWss76AwZhyRClg7hNZxnwn19qM0Kg42wEibDS0WX0dbtu8PTTfm0pfbU
Y8XEbFAy2hEmb8WTQx0F1M1IPYNrKAZGPg0eD1SByYAY9JEoJNpfcDagzPcknf4NaV3E9XcNze5R
hxuHfrZTGzXW0zW3V+ZnvL9LjwGl7cmcYF2stKTfEiNskcFL7/W4Iw7qD0eVcnv5ORjysk6MvNPv
3tx0zXu8Z4xvybB0Pdt3LCgehy6YqT6qiNkby+ynbA/Vlb4fMA7K+fnQk1Cfpx4zBOh/ESU2DVzU
OLmLyrnHADvjycOKitWKP6kvX0t5aKgrM8jmmz0UoQ9uMDrgxoORAS2kHqWZdduCQq2dpVQKGVSR
+MHwx8k67ftrX1TaWLUrxgt5iscFGd9+TU2zkgL0LpaJ38CiA5L8zkQ8Kht0wDiG6NiViTGoTMAj
NjWEpg5VLYi6RflDXi4Q/zoihplyNGsIiw1uKsPRG0T3jWr4LdtsE6OHwgetUzrKm1SXjiKA8x6A
XaR7pWPXsQs8itejMnOeoiZRD9Q9el8CB758q9m0N9qGrOOIxcwpGsKQbmKxmtpW1G0fONWZPiQ8
V9oWx707XM8SfPeiWNtV4TksaAbZ3gV55OGtIf62mziSxsK+Mn6d/JdvAgaMb2+jYj7+ynLp5J14
83lIKp0oabqRbPkgzTZnWq0mNsrsYknPQMzqlEGjlbO4JPfsjxqLGn+CN6pCU3Pz1jYzeKtWbyzi
HURW2KjGmOQTQGgrSXcXsKmb8NY8gs1cscrnxmNSMdXwHOZt2VEfgFj/rLHemV74c/+/VAjtngwt
ZV2JpCgtSt3UZBHWapUhILP6zJE5vBUIgifzpgwvXOR9Eg/UN0IZdYa8uoD83d5/zOUcSXVDeDV3
ny36meBh7UAhuKzo5binehOFwgilUXJXK5qYuQpZnGpOUJTS4zaRGqPkjjpk95zONkp1wkij5M4P
kRORwrPfY5wabGz2C+yugM81lLYgA8V7voNiXzh4q0dUQhKcoGkNaEYpZgAu3BYQqaliBU89r3qv
2TZ0+7HiYH8nI0EQcfPPzQJpR89aLu6MMgF4h01+eXeYoHImheDpRV4XWmn8mrg9PGssRxjHguPt
UatlcKvCfxhv9V/9Wwl7pEPwaV7BwzRGMl2+ow1snIQnAwDQ55LfdqpfrlrSswiLI6AC0XVFwZTC
83FQm/yEjua4DLXG8DBJMfwiTR6izJ6JRDMbxvDU2nYdsu/E8DbZ6u+Ow+1H8qAsXcTGwux6dr/P
s+wRSApegbuCoMkN3uaD/tqOj3AcjJs7ULAbUSIHWyiBWdpaZYox2+ce26kDbyVBJFcC9sloEIP8
l3HwItqeu1eGYz/oU3+Y6kb07dufmGb/lfhI30hXs8BbDc+rpd02BS5u1hVqTdHI9D1cxqJk0cGU
d26ZIy1VIcrwgkGpy2i9pDxqesNx65qu4VBpVQiMUcww5eT8pzypQjnqEnqKyij253LYwLz65jyj
lN0/sRyUQcvalvV7NIahlXWWjZYH+enQO5RVbwYjTZbZoZBDkt/h5cn+wG0K8AGZiJc12GhPDKKv
vi52W0L6rzawyN08NQwB6kywnX5dG08GYxEvkSccjEFw98q0xgwnJ9kSWla3Oc/J/hnIftpfk7zj
IwgPGYctcXZ1bFAZ++DiOrEoTGUZgknF+yp9pW7KyJyMvny8bgOmcJuy2N4rHkEPpuuuh5mo6zvu
BLm4+EWzSrcxC8bQt2ueVbYnwYe0NxixXLkSBnwXMXuM8Ld5NAFGlB4d3PpBv5AusklXD4F3VD2o
3x3CKiMhYcFxJswa0UCSgBZ+gYWU58Dg5lsMG9HeYBUhkhc6+VuYWBBBjmFKXV6h6TaLOnWYxm7/
Ne5RfdoSsPwMRE8PXwVbiDClqCRj0jsnDBcCs8Zz+vVVAeBr6mwJN5/1/F7YNbVwSgeo8pw9QT/Y
6hTU7zHtuqKKaYpREmMs/Uf5GyCCPtjwwvFC7j1zDR/5DIa6Gul3d+M5NeLr3mmN8P/B3vo86SIX
977ehOAUHNvZJGaPMkinHCRoFEhy65sLL9trZxpbukEyl0qYwAdgQVIwvA90ANNY5pC3ozg8zEv8
tB87Jo1/N0yXxnMeAZHPciLPPpu9kDztVCUzXSoliWciujts3zyoCmNegKYRHM2WwFIQ8APt1Rw8
bOynAPtRuACgt0EP7Z8fw2t3YS9410Oh1W0xxuFKge3RwcEUOq2rNdNJL/QxeR9ZfSlE7wyHD57T
CaSgoq/Cjoy8Q+BUJ43JhTQLbRICbdFGnzFaTFTVVPSpXioQaIQ+SDt1Mkx3B4hWlwkbhRrDENDk
quOBSULwgBs6GpahyqXwHkMkwrnKY2t1o9f49l6xUr2hlp9bx4s6cDhpF5QMiUXmIhveS/bTtuzj
cVm+DMwaIw+GwmBzAXkjjIs8hctHdnWWJxTBFd2tBErmHeCrsZ8bsunWg7/baqE1QVxEl9LNubBc
WDTXR/35TRyxXMxtKSHLEQOxt0/YZQHOrAZUPQT5Gs7kTN6fWw0sLpxPcZxi9KSLkDRgwTJcbV9d
dthS6vvebIqYiq/xY1MMc1FpEgU+qfIOj4FF2cgb9j+VYUKWcqB1Jfi8OQLLLh43zxI762yVgYCE
fAeQ4LFVzxCFzLzbYG/8D6PWxjXu/CmPlewjtV5lcoYQPpsABAgRTrJuYXZEe+5GvhfNs+OoG2yA
On4s9ytB0iMszDflrNwqNc1Qv+dHaRmC9MFpEOVHM5EWD20TytG6yj6OZm8ynWkwePUOEqzAkaXF
MD/juogemWxYm7L/nlznq59PKmWnhl2bmJR1iGOERGuJ3oi8FWPwASTocIpndiYDb3RhfLW5BLsR
dFrIXTmVoKqtPfrHroQ7wpiiuxc2yL4o7lQ5WpXT9SXew+AZwGpbP4CJaTi686jrSiNFZbV0/BnF
A4+7RlIi5DfNwQqOrVrdBBouM7dMaah9O2neBhLS2mE5GZNglI+l8AsN/Xv/qS0dsJ+X7F8Cd/ze
frCvw7DTYZQqr6dJzv2ln7PNSK1UlBRoWQ4l2NXXny9qQi10NXwQELX1ij7T2gG1v7jEHvluL0ot
X3/JhUbKC//1U+xuK/R0FKQz6UWQ93JHZMfpNf3Yqev5Lf1KtKStW0+faMH9bdTdOFtXo/lgVewu
yivTQV1Jc0K3mzJZn9giwelguykwM8oa1IJp/Nne7e8C2eKwpaJPdIBuCs28+ckHDT8nwpe3MZTI
0WFooJyJhZV0wElB7rQvMNsMIbzzhBnW8INh5NpoQRZIkTkm0PtjE3AQG1+ZRpz0sbYehFu9TliR
SexufJbWJyWNKpg4GgiFXpIx/tD2hGnTwOSKpLcoKUE1Cc8RzF18CyYsgmXN2Wa+lcEBErsE09rl
zmSR264S+Nx/Hxp8iDX1xIPELuMCjwQjHRnpy4nhvEntQdyuAdEwbk6Fb1XjEnylqlcrr5Bh+XrY
9mbRT+iJpeNAZ0WTIQDmzVA1x2Jw9kmtCozhvNn3/rHxd9mzm4BCE9g/CD0IFJFOLjarg2ePAVtr
9IyDUt1/x6uW31lt0kAm7dp3k8GQOMYRZxfg03v/Ok+/LoKmB0MGkbiA27HzpDNXFxuQJvAdAaRV
6ecz7ocF+dWf4WQ6jgKTpM4AJaCOjMCkZ4kaBLt3B+hbSYzz0KBH0/HgPZU/Fs8e8uafhKQNhG5s
hAznXM37wi2DTaQjubnV8zxqPQ5vcnn4KO2VtOxizYW1BzcXhH17XOFsAmYhEXqF6UEpGxJ7bYo3
wcF2huCcmiNrCV81Gx1P6RQaQVU9Znkv+LGJCtjykVcfK6SHzGJsooEvNk4EnXbjOA4u1IksTb5x
01n6WYPOeaudbmulq1dIjW53LvzOLM1nVb9Wct+4aGipQs20uK56ptcF7bTlJGPxmwFEiXg5ywg8
DrtxEwFF/cSKZg5t2IGmwKq2BE1WCXe5KI3w2lKHD8eGe46wkWlfEC0l0fGVNCFRwyriS0tPslTd
nNP8RtrYF53Uj01efvpstvA52Y+Hf6/hhDEsJCeBAcOnowVC80QdPhDJ/AWKM3EFeHtkzOOJ4mfU
YeGsaSAC3tzVtueEWEp4OtuK2WoTnnSL0zKM0bT76Ta6MpweA6zynKtuGqKet4nP3m/BWKyWLOnQ
hirRUF0VSAB3bhF84lA1RYxgyYWLgTG6/Tb8wASjjbFTipxoa8p44BaPhl8xDNFvl4tY2cxYpLFJ
XjUvv+BsoLYgFsQd+QUooLEVuqhKsPkFIX9GqQpfBG0CjaMp0c0eXm+HqtuExvRGUa61JMEbbinX
+h2NYG/p+KSzQWdDcWa/gdKR+68AZMkObGVyRSLcJuxLAR1BHfB40UdLtMtLOLRbOYq8fK6FO6SP
5aE40yjNa/RRpWJp7KYDaUlPiyjSkqwjR17Jr0C3xNObmMI9ptyoI7rQy34C1Rj1fno6058k7EoN
ttXjm1eezoTSs0Fdxdcpa8EiW/iMfo41ylK2a/LOcxfa6fOagjYrthTdOq2JB0WGOfwxGzYUYGRZ
2mTcCrywWGzmqhK/1CLXUkNRnCCaD6ydQ0Xh2Ep88gcT6W5llquS/CCy8XEAmAsqZLP1OZZjf4+8
FqaCgtmodY7CA1GuCWMC+szuOsDGjjX5C9snnr9ZVlaSDYRUUusvJQXY1EuHYIFom4g+hAJYmuOG
NVy/oSSXF6OgDmXCx9nCjE8yN2jwXEkzLUw/jnGw9S7y/m3zw0baVIHM7BBByJDJqIgocbV1ThQs
ApoKO0wWMeG37G7kUPo9G6jFdX53Qko+toVgMyM1XxwxxZWPOxswcHU1xTMFqZKf4iDBsckoGRrZ
UjuPw5KpNAOAj4L02a1eNIIjc7rmxj/KMotQ5fcY7faC1IIh0dTjr8RzvQCOcFOt4U4xWhhGEsgc
fNfjFncOS4ShiTPuh9O60KhrCjSulJBSCmdPk4bSpoH9clhx76qjZwdzTFkHi7cQfMJswDomilel
404LLgsHQt29qQ6lT2MF/Xgk+lUnT1mJDLyNJrcGW523FNzM7wjX415gfIEvr4mmzT210fVRzfp2
nVCiCj6IS+nsau3KAGEf5vd6N+yn5i1ToSSKLouC7QJybqKHvQOjLTvOO6hizOwwZ2NUzDfWI0p6
dy83q/q8KcT0+5gblrpq6eP/aUVH2+4hHPq3gBJjfD428a34sUKU/hz7LPAR6RGpZRPCsjn6P2Md
bel3B63tofpBJVT1syMrkjiA6N2eyrtB4eeBaVJYBELDm8Npx6yKPaHyMSoH78c0Uu3rr1yeUS35
aO5H9gp3mzY6jZt/tHBCUyBPKRADlnxWUoAARfs7iLuh+ZvjIk0dFFMPAEmnfg+TnRJpRLYdyhR3
geCU8p1YFwVvOwYgiiJlEOo883Da4q1J4mh8aFdOfnGkYOtQSyMP+Pv/eC1kSaoFiWHFfNyzGyO0
myG7r+ker18rzoK9QMWcIf/0z+xCw1WjgfNx7U4RvYIy4IvE0vCua8MRyN0P6CxW6XqyqVWNPY+o
mAesuAaq/hEpGIWEo47+JWfuuiRvTf43aHuEUGf2znKrSV6FEcCkib0IG3BAgiVDvXocrlmBOO16
GMRoJ2ZuhAN2rxRVuVJ2zcBxj39kyQsaF3/yr8OE402Y2EhNtnL2+pxpPYB2qh0tqzSgw61o8D6+
TXPyIPjihfWpbEsTkTfH5uSCD7j4tIqMQXjttqbsHTOz8KRSgIgmuM/Zr7U8TkaY3xCjbsptqjIS
j8dudTfS/x9qRWoJ6sLDblAaqcvLKoiHlCCoIjo3ih1niAjyN4/dd0X5tjTA4inntHyufI/yzavj
m8owx3sJ9l/ell/cyvpLgjY8Uz2N37ZANttGQBnhGRN9gYxXYqKFgeh8autENhpM4Uvi5rBNxNvr
9PdIRxjl/t8d2bzu05HmoRUH7EhzpRRcYjVihas4RkRp7VThjfE+6jY6uSR7IAVawR16Y/NWgTvN
/vrJKcqEgG92QjEmGiArtMfcKxTAWkex6zHniWJV/olsDz6RfpSrqurqZgwf47gFj8/zWLoKLNFu
S3kVeh4CQ+uQPMYztWVO/DSGeHPEkBiv8L0RIDGI4aAnkAck9SLtKwUx+wWMkSIj9PlmnqgDcnQI
lAb5A8JeNnsQU5E6SvPFkiYLyii8qXyZG5ElZavJLYmAY5jbgAKDjLj77nY95J6sqFmkWPL4C0Uv
mZJVeIAQy2kOvltcyutmp+y4WwO/r9zOPnpNp5TStfxDqRPBQCsycTnsSGE67MY8zpK1vlHv35rr
xkZ4oMx0fbAUr4saFrrWGpwRK56pusq/YiDckRXCRgkxxJXkwQ/h2t+cPdp58PfYLK7sYY6sLjUX
oRCKFiZEpzhC8clAAbGsr3zMMvPZWFI96c8HZLRRr/+GnyWgvePIJwHUWiYdJfyZ9KgRxqSimhwh
NiO9mocw7h5obvQ0WRfQ7gtgMtf+FEmBbs3xWT5iQRnumkmLFhNd3Lza/Ys3IMllZN+u5WaUsKfd
/E5tJpL4cvDC3t94h0cFk5yTrGD1PcPyXIR5VfG8FtHA0NLLZCQuC8o3mB91FS79ayVCSmiRQtq0
pK+8owQFvBqC2IPE/g202kWnAu5yShysqlid3BJUDz1E3lDUShzH3vh42vO68+lLLyhNF6OZ+k3x
svI7st0VQh7EzSmsnFMkcLkBJXPvy9h6SLCdQu/LHTtyShpe42XPnuDCgh8HtnTEzsePsJd5iUPA
sm2zSgbJK5Zb7SNZvg4U7I/S4BR/nfHF2RGPgnNGCMDwH3w3Vhh9Ul0403WMZseBpmhgSX55uvLR
vQm9iewkAOS87fcqap/6l7BcncqsfQH7u4VOWqE1ZIQJumByH00CVcUsyJkB6OBzdX4lMdgbwMyk
X1dnxEu6/9o85zlgkparzva4LdqdoD+vd5syPFLIYAfCFEHayDnuNBtqsZbJEHSuJwOXN6ZPR6us
Vq/EyVdANt2aY+2eTxWEeNilimgaxq9V1rQPa+AwyqLQmDYyTigMTqydF7y7onPbwkaqtKy/X9U7
oZOIEYVnP3mTt/Wg7xCq45OoicAVKd/kr7XlGj+toqnuPUHpQ7kURrOb8AAg9/IMtPtk5PHdMAp6
6n0cbwi9KyVsbb9a5p9FummobpE5O6u1xf8hPfU3WU+7p4qUhWaCCdCLXN2Ly0TCmR32Kn38+A2k
6uMCq/wC+ZIweBzvZQnMF6fm/5YHijc9x/6qlSQMy6oLfXv+d6gQPqEhpgLE1CPjCAgQkc7M5MX4
r/lN48qmLuOCVihlTYBk0sWFGYGG6lfyJ9f4mKjopiRsipCPlOTHoJvvjM+TP1p7q1EOekIPrl6t
flRRVm0zWW+hkL58U8noax7X7mCzsaReXuwEihFSAexFc7Qco010+B42LP+yp1z6X16IZWqs4klp
njJX93+6W0vm2HOAPptO4J8ILa+XK0tfv7tI84IlO0y+2kFnBgKCo0SFHp6kSAD5wcUuoZGYWnsE
UsGWWJ+/5c8IzYKJjKGdT+m43eFaxDbNPQlkabElVL1JU2k4RFTel46lgktuQ55ju2+GdmheGJyn
MUWTpOxAF5CMkERd0UnepW5GJzeJerIXcxTTIjcRbC5BzjlMBdqzzKTCMWKJRxpYA9AxurFrPdFj
ITmM97cERXUQ55igupKWwPAf6qqNQcMmOPW8LDSizQSXaAOF6urmdkuKQnIEEKTjtsPOW1kWkKtO
HdOzd3341wIT6EE73Y5fpg/bNJ5fnBXenwk/pAVNuGhPslGP63nyJiDhOpkx0RsST09z+82uXR1R
XWnvXV8U00qxF9nSai9PacwT0D/FbyahFquVitYLa9LM0fRzVmt3hC21RNo6+ylqE6E+ixWQGep3
aIeZ6+tkxoxIXvh+2NeqEslNJ7Br1GHAySkd9NqwZPTL+9MzX1zXm4TaWUBq4MB0m47vfeogavmM
g6M6Ym5JKMMYLJWa2vj2vTT623pnR1GAogsnis/pI+1qPVmCeuzM4msrwSc/ek0RVYTPNGBrRYQm
2dOP3Ot71Xskz54xsRWBFpWxbLnFinlg0gxFUXD2u3uwozi1UsdSTvHqoltRugOw/1PV0V0fSerb
+PiQOXcEpL7vyb41/plZMtrUi3nQSq4qM7LiFkLDnaqRdG2jNbhaQYajtbM9F4ysaHELLaXQJyDA
TasH1SHaZEtu7iQ18WJOVrzF3HDDk9aeEu6antmvguznb7Fc5IQvTjEkv4Qui9lGBc5mSC74g3Z1
HoD2SMdRBQrEDp5pYcM8X/C2ktRCdqsZzpbgybzM7OjrcHaht95H7CeyCAtnetCRjLdJ6BU/Y8X8
oCiZjST27iuL1LWiEihW1Id8Kerp6r+QDHK9z7zA1xMkwH383p+6JupsBzl6uW53wDMCj01cuCt/
BfY06V6YXjvmtBPMWAjxc1oqPPVJtM9sBB9mFKs7KviIfWFzEsAfUt3i6g0snoWKYN7iykiQmFES
kfojTfXkK/ouwTrAi9xufGcdaQvXkqMqkv7D8uMSD1rEs6vJGryBhVZ3Q/3xsypT6MH01WT8pviG
Gl06Vr3ISftjwtWUKBPubgdJuy41PrrMOInmB2CTKQ6tHDiEm+lGV+VcMWi8mwJbjvC5Ai8rhFo3
/QJ0sHrykh6FgaM4KmyhANqXrQdQHc7n51tnk+yChiYtrBsm4UOsuYa+XaGdJ365zA7/CpuXzBWg
UnIqhRfRmdm9JVUGjd7MIFJDToeb37+pIl3Yeb6Eip6ooOgEKTwZBHJK5d7iohOAsKAQzOQjX2oC
JWtQhc8Bq/6spdNp5FRrVBLKcxWDC64Hpw3UVRoa52BOd6UE6MYyGPpPY5i/SxTdvhrLzKzSixgl
KpszaCGb6hxBJTIxLtovPRlo2fqi4YPO1Pd+pQCHHXOlmfa/KxwmYdiHBcxCaBxQs5QJQ9uk/+Yo
5O6nZyZ4GjISrBUULD+HLkVusnBKezt3+sPS7fRE728QuQqtqCR9b6yh0uySYYuN83u/mwuzwu0o
HJP+xEpWZsnkwtMIcEQ3bmSc9GIUczPAu5fx3tUxmG6iF8QZcH++zDs1NQrfW+RCUjqZbQiya6l6
oGolDHISVthE+fEhn8kx3HVC8vU2PH+4IuVa+nYGpjsx7TnJ+i/eJxWcc0kBnG/3wjjHii2rnIkE
OxAuGSrNX3tPD1G68JWqIj3pRPycDcbOZStaYbvH7BxxGN4pBBcp5ddpK4LNDit2ipexoVXKChw8
Aq/FmaDCeE1MFgnXuYjJhUae/dnUW3Wc0jMEkuYhd1XHfp34IgmG7hSPTHxPMzult5n7kr29Cb4n
dgWkPaImknUL68A+am07yqHwQOlJIb/jW1ox3czo3yiH2Kv0OVc9N7PY0Tf8FcZSVCjD5LlDWIy/
QTWK4b70FxGL+eOu2+H63HK5B2FjJhyrQQt7Oob5VZLCA+sDtS1vmQW1MS3oj6LcDjnOKaprRZWh
Hl+DThsAZl4CuNj+TKKOQRP9D7WbGZYdDF8zO3AVUewDj7ZXWsf+sjDqLRC1IpC0n7gD+lPZPQyW
U5mhcXeTi/DE66w5d8h0Z2eopDCDTJ4vv9UrhcL/i/HGA2SQ5eKiGC8+AVjGmE0feeoymHUuq0f3
xc48ux8ji3qXPJonfsgaxN5EeGmLHiJqm6jGAusoA+aw/imTgggxEZkLZyEXBFWweOEhvbbdLSBN
gwTxU3eoZ6Vt7/Mvo3RrKnvYFNpn/Ezl7TxNYOf525W6L5oXBN/PaiHbMeXM7IslOKS8bESmsSky
QtZpb+uE4r3Yg6EUAjHuIr20UVV0A31bHSrfQL5IcR6A3PDceihVQX02D3SgHeQupG60ieZD5Oqe
ZIKJuWiNSvvZYvodmTJulwlGpPyKX981SI6pjRXpvu9mNL3VmVGn69GzLrhZTS0E3o/xBRPMUcOm
/V1IrgQppaan+HryLzFHcom2bFOMBjJvSPWgLgo3EXEzgxgiFXv428+2xLHPdDUbMGxJETg68MjK
tH6YaDgIRjKM6qNgBtYzRytcx+54gZxbkoAJnCCEPrZ2udIUUCZQg1WtraA1JMnFph6AWwrUkSXY
Db0fLLQ1gtSrf4DwTbsxqtZRk3iYBU2jGyEZyorPlqypviCNeiV7gzsaV7Sl7LUTYuMee5Ln+Tgx
HZxISW3IrvaOZg7Y6+wUITLof/EWEIMWA8MCJc8BN4oZZ+jtz9cGLahq1S0FdeS7CXExm4Im9Ahd
0qV9L0Sl+4kZyEb+2U2Gd3xcTnFspX2KpJX/WT1PKCxeHY52PzvKq6fzbuWRiIpF/gjjpx+KCbyY
6sN5BTbjkRaDjwPYA+KzsPDhC1tdiHJYwaNNRMetXH3D2OCf5YGDVFktJ1Me++++YaqBgjUJApQp
QiWuVSSBO80ht9F2VOvqSAYdOYfKEW+P4obWxztkdhu1SF/bcV6a+uubgel7sEWK2eTMfyaegfFE
zw8Lrh+uGMltoZQ8gfxjihhdozDnnXsFTycwNlBvqHULV31uUtDJL6UWIyDW5XiJ17Tvv0XBZ2Zn
8nsXdY+EItI0YsT5aCg31gAWcoAk+X4N6cBC1OHk8RH6Qo9tsOZgOTavDrFXxNan9T+cssnyzdWD
gX75uNlO74IgVZkHHDn75BCaOB7trLtngNouepFqx9n1W4TtBWp22CzWcrzvJYz8bpqK6AVyAucu
cj/5LC2T0AjGgpROeAO7e5xKzmlYsO1QRbE8X3SOZh8STecImsLJk4gILlkkJ+Hiu13xqx8amsJO
bwrWNzspc2KxedfuT5PJdYMThVyr0PyGX8I1w68CJGmukZ74eojhqhhRUL0YauTo7/WPheSZjFj0
8Ds4UnTthfNqpYIgd9egoeNZEOIOUFQ/FAnADZ9YrLxULYUaYXCrz+gmJeTCtSnmtAES1mnGcF9f
F88Qt4rQjUBrgOB+lF9yxtuPZNos4qtAuWO3Rs+qKpKSTV2M1Wr0KNYdJPJv7naXIFkpnmfTniU3
/GmMWyGLLjSjv2f5Vap53rmZOiT+EsouAVVdTHk2IobL09l3c9qZfAXuAxGByQ/9/FeyeLMzWIfa
54AUHaY8eZgMXrD5JuFafNDFNj5MWl2bTT98BB7Arv9gD5sy9dBxsgElLf6EiGBSmncZ6cHAngPl
2WLdBib3hHu61z02BdKMT3NBlpiBkm6xvl8OrN/MrGsN6RifoUb8QB11aQ68ColnT/d5Wocy+Xzl
BfI39AXsVXbYGn/tc3J86cpuCumwJTXNhYqBsSeYj1AkTw37iAAVusvGeDpbeFQpUSKSjosjuVH7
XSKEjVvXQS7xfY+tdu3vPxA3mAfIItyguzd8Wgu4/jeSXl6qAjvJM0vNpzRIXO7QVtcw9iwmESvp
o8CjNxgNJGunqxv3HzLiP5MMX2XzBP3HwipjyKSkJqUMSB27KdkZ9hnU9koD4KiteDf7NutcAnjB
wcTB+hGkC89v1QVP3HQMdtYeh6vtUxrS4LsOzkscHX1y0FCU7E+vrcWIX8m0Er7QAHfa+LrJje1E
xHk7FP7Pts2yCoj+B5TINgsO9WyBjOweumemPa1bNegGpjvOkXCsC4JF4U1u5AVWN/mnwYX2Valx
OP7yvHUOFOPeoKviYWZ2a1d5pJ05TrCd3JQPIg/JkChL2y3WlIz71plV1n8pXaXXfeBPbnrD8zl/
/TKj7F1Z+FqQ57E2B5hvtkzAw0GdnwNY0WmRB02GNCcB0vFAzPgiN3NahjaEgfszh1KLu6uj1P/V
9alHcNZui6La0QIisytGs3xtYEPat6EtwOsgdsdufWzQ2keGNFHKaDs5xM7ilTfyndewWeG73ShF
oTLOitWSa3BZ/7HL9SjEWdA1BqG7vwhUJqHf6LAHyLrH7wNk7DGrzEGMEqH7hpPKzr7qSVKq5Fxt
MUQU1q0EkbSaCtOnqq+fkKah91VGwfrnGMdH1zVQYBECh/kbbtymKKfbasC9CkZMX35F++IXz1vC
5Vef8oqupAGn3Li7UIBRRXd7bRBswKtkZbCanKIEtxg7g/3sCqzD0UKPUQjCS6JRXBnHoxhZAVcG
SzZVhv529IJS3WPx+1Go16T59KEiuOTvygqpqUsSJf4Vd8OcGTE4D4RxIF3DAXS0xyBCOGvRmezS
WGqWBwARWyAR71VRpVMnHfVRTlIH0z1sXhmYTAOYu5+v71HuCwN9xn6SDq9tLKkY9FP8RJFiP3h6
KmPlODf9WbWaJhVhC5kDCU4cPfZMBhQAYXKJLzy9l3Lk0HJe6x29m4ossmzmU3lWxFCUFqmKhdiw
TObUrNJQ9YJgKOolxlXyWPDdAQz7K3lFXNJQ3Wzi+mr/UceDGnAJj/DvtwnmZ9H7U+E53MrtUSCU
CWs55CyPuMmJpVCCE75nm2IRU7p1CiX91wbJsn9tWF5XHi3IN//PC9GDm4yF8Rm1YXA1AcLqk6zj
G+X0O4kjQA6ZJXpqlp6phCbf22Rmo6Cb6jrhQcKrqu4VkjRvdhbTU1olXG7Fdv3EFxQJv3XeG1Uh
tRuxg4DtAHc9ZA32NDf2hUzYPfFXHzxfB+ExgJhHDI6FnMSWB3cZdZaBzTJMofvVjyyPPsh0+OBC
YcC+RF4xqcjmyhI6qjwSfXxsLI8TK0LRQR4lSYP0VyzRbGbUWONnDVWZqLppY7YaEeI+bJKVcWeb
UZp4ch556TJrQjdBZhutdJyWrIDOEeq6mAx9NyXT3Xqge/qt3as2zugJUa9ehkJA3BeYGFQrApWo
rDvm/eMbrOmrr7n1u5dICv2xngxiTsuppJsVxrbPUSDI2ilZU5tF0OeahbHajeaqXlfxicV0NJpU
PhRsoBFnJ67BdAKmX4RcqRDTu2NEu97kz7w8tgonArRdJrDO9QoBpt9vPK2zJK421xX6A/yifiTm
8C63xm3gKnjLduWR97iFHzAzN6iVkYXwbfMzJMrVYqbsFwamIDunTP0qBGTrgBn3ifW4mL09Zlmh
fzPNawYwx6YnuMT0ziQjHUdzr3P2ruZGwSOfYCOODJgW/DwKVvGcL6p4hJ61eX+O0uUzc8tqtfuk
7BXDIYvelZEAGlO+Fo4zywOAYc9SdAY6gFUbdv+XxdgI8u0pvzE5exlZnu4tJKWHj6+9QDabaiNw
0extDs78xHQMmHroe9AbuxRWjnY3OXYD85HqxOtK2gkuJnEC5uZD5yrn2wga4av7i4W80/13rGwI
a003ed/6FGmqJ2IIa0cRvbwP7dKuiQSxqlImCi/Z90UphVcd3vuJNIyKbcyhRbYkwa22QNaZcQ53
F2DLtrXBVc8PlhT/ZDicIq+VFdzM+HVAL7dmM4fxLbJMg3sM6LkSmhCa4iMeK+2vQ+YmZ0CySuXx
dC+Q5ZYJrJTTMLauc0RGHiqA88V+1jyvaNXEDBCUiyTXmkR30rcXqlgq3nlfuaWb0nbWadUi0XKU
y3L0KTDvVzUtoyaNalqZ8bW3uVD0Q2MOhDuC5o3/F6gaAQXdRdziflijtyla82adfX+ei+w6nEpK
8AFrws/pREfapMgDLsssWybP6re6YsXrVCyZlGKQT+kQOBWZjltVBSCnJmH6brcSuikgZaj/boAE
wmDjEyIxa5H11+8+PucyxGJZUJvMnlHc/O7NELsDDtQgrsp3to81s3FqPxrUGLhM3xd/hBW++Mjn
9QNvbSNUWXB/vwxPU4hJy0H6GbdoOOtCP5i43EtKcxjWAbFLa5YPKgXcU2UI+OsqUMtiuwLeFN6C
CutW/+lrbGLp94zTJTWZLz2WJLsRpqwdVH7vneXYxhlIsqvG/1xz7PKfxLRX4te7hiWKDQq5hOE9
5vlTxCYgFRcQqM5BSfWsU2rCSWIq6INzFQuVUfST/FtXjphdjgib90WhUjvNdJDYYGxVWdL3Pr9x
K/PT6hDSm0wo604rMFwM2uwwIftvbo51t16BHdNNdSd2/KehXoDkNnaxFMU+Gr4RMRPIblnz5SZG
LvJql/UCyzgj8L6YSQ2RuGYdxRTquYDDb7tHZmR6ylKc7XmxOzwO6OEyTGTCrKvAJ95KJZXTfLbz
1GBypSKG3PIPpylQBwramX1FqcSH2RWIp7CiucfzQJQEUDp2rrBpSNB0AYtq6JlWc2YjJTeOXg3m
lwwvKkRVJv4PMWguEKcCCfyPMmJkc6cZlkir3Ie2fDjVn6Ls8BjyGZwwJHpuPK2obFAMbvDdyOJX
krNrSlfPwkzg+rTVznvike76wMoXVCchw4TZZJvSlgKY9bLUVytyzA5bvUaeA3IcGkCvc4o2l2//
FbjzD9g/nNT2hUVxLM5Ih0bUxvK96LAadkm2RNiZOtAYhY7yI+rylnzPWYhxxvUoQ3qJqI4XZpMD
Vhumd0t3TrAarfFS1yXKnvWmXSNIwWFfwTx7qKusw7uBqeUMeqobMhGZE5IQFTfwPDREDaeIYaHc
zOdVsNCcnlgarV4/aQG3/TA3CqBaljiW65fjg1PLlLxBwKH//Cg5IznVR1CRyxGdbGF/iUHKY5mD
dK0w/MAOWGAWYtZc4nX1u7o/1ieDKhDyQ53fPhwe7M8aaf+ofBeR+vheo+sBM8gRkzXTDhrR9ZcC
7lbVCcb7+6b3bwe6n57mVZBk/2yHom0FIThsBfBau1A+fSplj83p2uID5IXE82iR8cRoW9y1FTTC
9az73RxOJmDXCI4o1UAN4QonHaXgySXkAm5+R5RuEqs7HOPMPwcWcAN1+A2CCo5rDzJQvg8ugjqm
XAMJUfbUoQBRtXriRx7VotA8zIJioLSJ5ZIgLRLDrU1pORMTs7UWmJBrSNmFI6P/T2kXXSj9gvIW
JmIHFVv71yDruVs71aLJesVJAc4Wa7SE/fZbDPak1RvMAxziCijlFdVDAZ0NdmkabVwWXWsdriJc
ai9oXPu/bRZsfW0cZrlViL0ce87mrmR5i23tf383+XqdcJZpvzY0A7zwZVBsFrQ++y9jk6ToaE6k
26/ryLJDCK8GrB8Q2YDkLzbh1uCbb/X47E58aRKW2l5SZRGT+kt4vs+zj6CQnLAilLTT0gOO8/9q
UPVL2AEzk4+RqYWmwKi3psVVb5hG3mDKFfpMkWcnp5OCYk2gOoUs/NF8Y2XkxyU+xeqrhpx9px0l
liea9OiO6m2a2gXfY5XZKkhWm/IG8HC2taapIU1NEDXWtqYOL+EP1RPVmnqprbbn+h/0L5p1JjYc
ZoBsaWvfOWtCTUQr9sOGu7ioFjTzVgsBi4IkCG7Y+8cdKdXxaOD8DmVtsprwqGfr3056MajaB+up
3E17/O4JSlLQqpfnfynAVU0kTHJlqwLw1zeTccFw8FQTJvGxobus11nrYChQB9Ai/piOa4MlDpg0
gMhQYfF41rdBWAnUM+v5XdYhX41cTkJ6y0vOD9ioA+YJnRvmNBVuyOr9a5y6xZ7oryKoL8NtAAFv
pjFoVt5n7vuaELXyrEX7XgNDhfp7uKAlz21tNq7vuAulPQngMR1jVrl/umrYqmOGJ4QPDXWvHqqc
GtZ+NWsfQbHbB7AfyO+OYpMUq5BENAPkxRT/+erhVF8ikb5IwoAfCay+AdMEh99u5k0G05hHrrDp
7F5zCcZ2XNJHZsp97J2PiSwlQ3RqXLSrNuAKlkV9N0KXiLYd3ldtGjgNAGlcXfa1PdRA2Sy5QOQP
9NUMfp6wmwdSEQ4bl+xSlnA9MekONEY9J2RTR1L7gqoJyhHdd0n5PPaT9HDCtmm1g/4+I0oKnx9N
lkcxklOPP5M1KLgbb8KA+9Tp8u8duYNgv4ddjiGosc3ScIGT1oEoD2WqYeumCUzfBjhEZIE/F5Yr
GpT2IIFnl2HLy9oZwC+AE5kFF6ucHFYt0GlnIHdEPaPVPp80drFB/Y1I6tvWdJd4uZRBtBo6TefA
ytlLfCZVXzWmOt6bg023aSFBKUkPl2BrX0/LDCQuMBSZFKTXA3UkXNERwTq9MiJV7wSOLgbWF8xC
PO2ssomEDc3Anb+iS2hEHO7Dh20TS3qZMjoOrSm5fHNcyQ3Cn7usGIYpbU+Knq1lPROLTyrhg1yC
hoGrA4TYh531Mcz+uGJsDYeVAOhU5pk7h/jzvKzzKzGw0GjnRsKWEUxO0639D40UxtW05mj8nOFk
wvGdzAhKnKIFW5UEK85r6T7LwPq8KfZK7L3ll5p950uk1FOactNZtSM0NRofSyhBwBJ7aZXAlG04
+GQu6PtgA8fq0nl2AugDSjx9x2WF4zWQosQZBRSQDEWlgaCZfnsgd3K4mWm9ElKDs7Ryxuivrfgp
mfX87boXCCVvsr8o1t2M6i4RiimDvXlnHyEsfaLGtPqBzCzx/MO3VsBK1Z03zVMfroPNpKRct+bS
cC8iOKFJ/WsnChurU6IPKKvKO0xI70IUGG+8Cc2B0BXjgYJpq/KVFZrDmtbhTA+8SexZSVvr3OG2
K1xUr2G/+xzkS4FgOnib4zLxJO2lj/gsZl4FC1r/c1E9xSVPdnlThZEyuTLpwogdkjLIsTkkjg/w
+zF1JBKHmEtsvdwcUbtSg2CeNhsAUu1bz193JfL4r4prqY6sRtvLCT+Nu7OBUoqyyecCNjF6teRg
86pvA7LgkR4yOJatYBKu8+rNg5uIlTcjBFcRhSvIPdokaS+RfPMvJNJ67WV6flUcSKHKHuc60MMA
Of63WDR5fL597VpZUjksCb0+vS/n5wq58h9y3Vn/QP5hT8J/+ifCplTPj3NvAI8N8rV0cjiFomFt
caKH4GT0FdtZP1eQvFxY3Y/spAzskOIVHaECcY/mV2mFjQvdZhPvGkbFhU2t2WpUreJ52ocAcqse
SR0fB/5uGjIJxkA5NVNsovqoOuDcsa6/GTg/LVFxGtzoexL7ymLEHC4vlRxoBMGv/sb+sX7VdBmA
n+ZrxaTYw8Q4WHIPThSL8cZIZ69jye3hujmcnM/jV9Bh3vhq4/AQzGrhxujc/2wVF5i802kGbqMu
S0t0vKAeRxbLpmDqnBb8ehndN4l1hBJcbzh3N46o8cZvMMY7gqevPI/JLCVUWgfsgGEnHVOSFLNL
5hL9XGqWH7Jt8oBPVrKsI1gVPBL0XYIelcCunu/XPWX5CaLjgNQGADOU1hgWOYxgI0axh8jaXPpJ
mRyBDKrBpMUMc5oeCVjf+xBUJxLv/kvTBkcxBP9RGj9Yt503Cb7aiviI+5JrC4Q+H8szTJZtTkc4
WX4pvNN6mvTNf0ebwUKfYjQikwDMRbI0c0NELAweIfvmy6wv4kDPuJbFsKNoaDoNugVmietYh3k2
AYyRcXNSrWQ8MGPB5wHOfS/Ke2BN+Bd5uSQDG9bScvZQ0WROk56Dwj90s+hPN2fxQeqhoc2OhUio
iJehPB0bXQHqWoD8Nl5tt1D5QRngBPvYRqcpdhuRoyaB14VuIVh/C6fGUAp0G2D9hBiVHaPC3o/Z
mNPmleqwP/d3aju1SJb7NSJyLaxLlm1doZ7e/JsxNvVL6MBk2Nvio/15RFuKYwLnZX3UhjQo9DM6
Mg3zKQws6wjrRNUiAONJLzqzf3zLh/9g8IodHVOmuiUo7Tx3EkM9QhCaVrlEfhn5u1Ni4HufUIKb
M+06+2oq38NpnmWdr8KxADQJq4+JKXK57NntJHOviN+30qTIJ0KjRe7e/Y7VSSsv+FJpkEN29e6W
eVg52B8cuuTG5UEk+7m/CPoGGZtcZ380wpTZBXz1eRjGTssB0qSJWRsqoF3Un6WWBDZ6ZhD6+kr8
cSOBT/JjX7p6CH92z35dsrOqEvf5jgYyYho2rMPiOS/LmOuAx25yY1ww8dktfAPYsBsGQHXK0b9r
KQu1ofMlM1fyZXDamxB8YYEPOkK11/D2CfKy2wHMsgk7z3ZnXJC+wFO9E7j0Zm28TJyhRyzTIgJ2
rOMCZSMzQf2zrEnOpJma2grxGZHZAMbY7FGqqwurJBwFHuk0o6iRWElbE7bJdi53IHdegsWgNZ/5
UtG5yBfzDQJLYfJNNwlMKbO2h8onxTckhT69yqc9DGPb9cDcl80uK2R1ypZXXo0CbiphCC4FBHBP
Dvmsc/NsvXV9eJxvklGosKU1B7yiF6AZSGXRYIrAxb0bTp6rhrJ8qQN7C5HEoVVSO/Y6FTMJuVuA
zPikJq9b67i0GxBKkzwqur4Oq9QP3Fdd077GTP36HEpybFo8wofxV+OnZiLKCEd9QP22yT248HO8
gCGY+mr61nr9QnpAUsapSJYmrkZqVBhYWgM5x0ncgmlnERQTXxH7eYQpQXmMVAdArFHIsFigMRWk
hDo4CMJxsmTVlLITuR+WcL8uHaXr7uyB/sqpK9RC6T1oxlZYcRDWx9RLac6SdUnaSAmTuJLaV0JY
pBWxg6Mj3uT8sziKmAbAtV+ghNRHGekgTH+tqj3QYBSZqSHrzErcoEw6JUWVC8iv3bD1ROfu/qzc
nf/zGSg4Z2TbENKIpoEADZ27gIo6R6neV02PpOYnE27OW94KJ7VumwsI+4C29YRU8LHKkzKZ11+1
l5z3TnzoQ7R3q8FTk8xQsTnNKuA4//b9xMCLD2xDE6Ihd4fGxcmg1uBRCeEJbCVlHhLyduXn/n3t
GP0ZmNfyGkoAkuDI3iod8/Qc8gJ7Lp8EFVfi5TPowu6QrrZAOxqPVB6Hbg3yfRva0VDxbyk7OZQq
PjLYi3/aLuoydfWiLp2OHNs70mCEkdCR4qBQfyfGRq4eL5+ameVz2IbZ98pbxDYEOg21bwPjAJ18
9N2UsADp+ybjeDBfuLyrPI+tSuIuibU433l8z82nBVONE7qT4yNItShcwAQHGb49MLpCGggxJoCD
WOaxIk1NUZS5rxtXbJv+falh4kg3YOBWagEC+vwxC2Z3s/7k8a2w2uujV4wJVqaJKOOgFmifEQhm
ZAJyzKzbUCLgpHr7Cy3LcWsdGVPEamZ4wCopt6oCNhae7nK2k4+mMPFA2p/HHeQqiAtPWEnMy/Fp
9JTmKfbnMHbjZW55niCrCrJUyBx3dj5VlILr5FrZu1XUHITkxZH9dfXXbXXa4yaeIJlnZDj1zew8
nATo6syW/t/ehv48Plsi90FTtZq4Zx3RatJGzvVGiBc+BA83XW1M8P8gCTaRCE2s8PYg7ji+UAi8
UrdGeZMku+qt9+GJmh8N/MAEUGgm7sLny8muVPIW70ojhCXWKIEe/rvPZ3UQQKWJPdi28GzVhYdI
Pa0Jp8e4Y47Ua4ar8q7LUOQussWU8qaP3RVFXY769+DZBi91S2jWQdDriPMS+akLqq/QG7coz0uB
3ZBDsDzpVjzuZkSvD9XQmkrfIzXODAxdeoVF0/y1dQkAy8q/h7IEg85/BEIvjOHQfDVz6dI5i0lJ
gxZweQc0B6ZQ8NDVL9/zVvA4mmZcHc8XBmStLJfXyC42pvM+gVcWy0ZV3M+6Gr41HejTjvpExSDo
EPQh1YIfo9aa2eYGbXlx3kt0irR+ijiDZ28WmyeBJna+M/WjHH9OyWCNQgXpwFewjGkX0N7ApSIK
ZuRm9ZHQQS59euqy/xmjqINvDnduJLourRvVIB/REYh1bJtLPoUTgYCQ0SQ0i3Xzr8ICGQ0Uw7p0
f1ETTQWNtwgz1NhTtBPC+UFhD3BClGdICv3JC5ZzMh98qV8Lf+1I/bOpZWgC9N/FRTA6UxsflN2K
zwRyu6MZb8e/rCYpxXoYIXLdJ2hGxL97heE3DfilCRd71Csq6q82sYusROZPq7eH3DAdlhVPWzYI
YvJpzj+WXJTyQcDY/fkPfNAZN1Tlwv9dPZC5XdeKmHQvh6nDvjMxEkPNWo9uDG+K55k9kOgeyoWG
4tv7odbYfUzT8U3NBhgWnZISbqenwsk/wqaWbTep4q/L8+ay025J4apStqB68yaT/+FAxHA0jIVS
0p3/bl3CAR5EdVBPORrX4qNn/YCx4Jtbsd6mnIVyuQspHvS7NyW+hYQYpBmWqYobWDYj/x7KR1DK
U5jF+8boUxxfoFlkJ7puWSjF6DMx0KTR/aHX2fre5ECxNEe7C8cRZLfg63fpsqPaykQBLAy/qTyN
iA7bomoR2+HI10vsU0TZrHp0jBytyzh/+SUYARH7eFmXTHFjfwbym9Le+9xpRCqcBRvSriPnXbYH
bkUj4u/G4RyWdhOf3d+YLKG9OasPXBzIKatOA22lB9pxKbQVhSmm8bVIXiSG76ojjsF9+9tdKpfV
5bGOwhdlF3GndBNR7PlCuKJBY2in48gy7Q7Rwq6jQnObizkgyLzglbybRTKzK1fQIxHYB+Y0G5np
gFLf7T8a03nQWsrgs+Ps24ncUcNxY5CeLfX9NNwhLysIHZIi5ImxqMNIq1R9GkEKj0EWSwDlzBph
+snTcQWYJk/4B8Tqwj/agno62lNlRr7AvDyYwDT8MX/ZcMAu2j9NOX0InGNfAxVfG/XMc7uZeNJb
3MfBoJ+86noOCf/G36U5LJNQ32LAfnlWWyhj4Co7NYufnSBe1IwfJTQkQK54JiRbfvSp4LSVzm9J
qz8xyte1fTR4Zm3XAZSUO3gOiGSVnjun57l45jcv+i53iKbXiiS+HyirC5WMuagESDyG7t7bV+P3
fYbsY50/wsqhYez6YDWjDFlo5N3heKWpi4A0SnzlKWhTJ8hBwxr1dC6knF6Nq/in6HqaVfEM2zOE
66tbXnBtr1dPYBdGh/iuW2Fnb/2qEPnhrMyCV/aN5BNJ8yzROLH9H6/eHSUu5eP7MMtASRJ0f4gd
HGuou46+aUrx7CfiisY6ksppWvWfbAe+q4kSCCUFYLlzAhG69NOl+DlwoG/xO99VkH/F6npLdviT
nkJvNWw4Wrxi7QQaftrYpPXyYukErYn9vwmXmG0sIaXdplgOCW0/25BwjwtZlR/0Mlq0Tn3su7OU
jrIRzswt04RQWD1/OQgt6wJ/hEHqfMhsoRRjGqxlMEt9LKvXUwzMovf72W9rLeVCdUDE4W8iZqgK
Ey0/dUfeRuK1wvAuKvwE6zezfeR22TRxd12V5I83M5C7xmYPa6eJbxbOsNJe1LK/f3EUiu0mpJSX
J1USDOS1f2L+05AR4Kw9nMp/a2oHM6wiETaRTUOYgB5fqUWCW4mJEiVZpzV5lHMRlixJoNu8S0cS
CxARvBXgeFo8x+vfP5xV2NxVLyFdbHllIB+fS3MzChkfLz67TN8cqe3vsjw0o7k9c7Qj/F0OM4uU
y1vLcQC9IS3JPGj9X3Jx3j/xJCFtm8ZFpL/+hnty+cIL5Qm6wF5pXn7LUQmWpwRGX28Sz4zFl0DB
X+Vr6pl0uI36riUPZHt83qHDlp+ieZx0Tz5HAZB/espbjsyL4lzwYyaCul1yqE5rAxb5C05Wh0S2
zW0CRTcKMbMVRCCP537jY7laeHKWf7W2vkD2SrfHfTmu4clOWpADFGICS2AaLRvgbnhKdGbFmbcc
MrBobX8Pot/wdspY+VruN5WO5rhO6SgLfAlFl4AHHzPx5x2ehCqzYdeE71dtKfhJGvo5m2sUJtaD
2xm0d8hjLFFkP75tsxHADJW7+xk4Eux+PVir2gV7d05XDT7GsmNiHx6RM5CRScB83qCuZIifr2N5
wEe19erFZ+iMW3yNbTDv+7m7snw3V6XYx8pnnZ9r83/93yUX8vU0JXdF+nHzVXdydksvYkwF8avX
/xDsmyA2SoDET7LgtRdNKGv6jwVU4oBwztI4/kUm5yfqzZ4+qclXg62F3++Rzbx58l/lQXfzwpz3
nh8cczZ60jGXeKGJ9R5CVHg6O2cz0TS5pEliuvJyaR0bq98UNem15Tnh5h1kPPDa6alhzBu5ccg/
5EeuKODqdYYyDnzEDdzpht85FUWg2IWXVwvNkSzxFDxgc+pwjobleFqFHrAEn70M6ZNZn3z+iNKy
wCvXMfJ2zzWOxK/N+9VDGHDkTzNAe1NQMNuk1p23nhmoL4rSMuTMufWSX9NZAOao3V1AaZyRfXbX
GCO3hHePqewCN2lPMj8RyJrsf+p6r9MQ0msATfvt6tR0T4jUcbhWoSU63kAUyXwgdnW3da98Ebag
jz48mU2A8tTER75Vbz+QFWgVHi3gTLrf3B4G5goc0pKx13m97Rdgrog59XFGJ6/Dk4MoXXtAfDRM
Z79xjmi198CqcTW4raOck2Kyf1919CVZWsnz2grZjymDm/EgWNtQ4H/ckA31utrZdKLkUnijxZBv
RoKsBfXCAKyIGn0dcDS8OGPQZxALT8pGtlUqhaOTFI0vRAPT/VKDQxs8GBsklow2VKy7YhgdJ8RD
GvdXTv0y+w/ZRYiuaCly9rNo+AN0ZRAtVW3gHDI5YHHN8rugjCOlhr+zHMiHSwnDzqGzUwLTQXQJ
JIVyHECsW8TH21z5WXMRYXyvjeqkPz0CLAJx8oHq5Wqqll4EqaXD/9PHf+7ar3QJIXctxWbWmID1
w2KBfRtBNXXVOcWR8WQ3H8fxgrgW/TwIVNT06x/IRx+7ncAq01Zgktqm+borB9/GfSZcb243o7Ld
0nr/0trClIsEmrVUrNlljtEaG+B2iDmEokzX++/Q9Z/tb8Uu8SIOeTd3AzZLLtyi6Ogb74Ca2buU
rxM72rNpyKLdvsZpcmKIw1EzDWI6zDowqv28+AMbGd7jRkXdQf6I7Q+rhUBMmgl8b1pKtpsqhIIV
znIsskmaIhqytsvLP48gLAli4nmXf4C3WqhZJrXFnp+R7DvlLUxvSij5Cjr8z8bi7QTOcjQu+SEf
4CKAht3BB1HNUbJ2MG3B4IAML6rCAbW70pwYqJWN3cprTtTuiM5gq0FkCGxp7KIbsefpoQANXkYw
FxhUGuCWgV4NJkiN/BGiLXv+ORnE0Q075T5jvHqPxJ7k7x2x0mHxY20jerIEFUIEF5iAXnUtby8V
8N/NhIX83Y/1rw0SNmQ3tQZhQj4xy4p2Dxs3TTup/8iphRpy8AmEevJ8U/acQ3GgKrUE5ZG0w0Uz
vUrgHEkIvXO7+TX7fwJDx/WeKwBYQ4xAZWJziwQkiUC4B54xZ2ryJZcfTp3AxpsL8bsbg5FpWrC5
HexIiB+amTjhx5TGYjTphXXgksHYdBNUk/ZLCgzCiPtk4Z6BSRwHXEs2689vTNBPer5tmVcj66hm
kHmZp0EfaeHrq31pRIEnrAxNrvgIaTkE5H7ukXwnpoyd1AeUtDqK0pJmXikA6B6oMCm6GgmOXu2H
4QPXbJkrjOUAg+yEptnI+O0u8nuUfDi10x1Z7rfNd0+SFswH/yANJTvduehEoTw/I/yB5Ljdg86E
ORqSgYEF4jU9dLn7cLwV8tNk01LbvPi+uwnw6txFZaDxsB8Xz6GA3/08oQoybrpmIueA3C3lIYKv
iC5sHGAvxGsrQ2Z8lLpCYGajtiA32T2iHh01fWlU7NtBbB/KnzEL4Np8KxxFHfPJri5pUV9uphfy
b4B8IiSX25ipaGENVGOVcFn/PY2iC+hsEkTq7qZWLU5S9adY6nZbS3nfhoXXeLZbCMOywEL7RgK4
MSRjnkTXaEmaNmHTH3LelnmCWbFsUmXgY7Kn9sVFpy+3/kJ1qAFXf8e/Iot5uAvozJhKcckEr/1p
13vUV/wsTkMyw1Hb3Zc1jOcOBGayq0b5SApfiB3IywwciM1+nd46+8iGEchONJLPCnbpDD+c+6Qj
T082SeeLM8FmlZVhZfhnijNDwcktiueS+IDp9jaY7OEElqpucGdPl1xpMcvftNPv7r98b0i9zzfq
WXLwsLvh8d1aJAACp4ELK+QkmKRU+z8hWjb91B3S6Zjvmbdi6wzyEm9fZXMSpwojk8SZ5CPkjULR
thQniRTffcd4G+jss2XO2d+34xMragepkHrBg3rq43SqQWIplqZRtzrjDd1IksxIPJi7ZOdEypF4
E8nEODOlADjMkYr4afQf7LptdMYvtuOlFNlmzQqwZVysEpT2oansrsL1VNftSAsek7LKJqpbYZ43
kLkLz8Gu3U4j+hrncdXLV7F+ORHWwPUs1IuNFLqkESNfjxfSpy4lx4RJxmBc6ObdliuG9lo1T834
AOX67UU0NDBoqRCLTKrVj56mhHpG+FqkhH9EJA5x2ih9vmj/MljMd9LjljNKDKIYXtMt3RrH35+4
is0whb0y+1acG9DWRub6eUDbT1Ihfjq+95PEAIyfXlEs8su27WRE6ge13nY3lOwcNPH4EH0X2v0Z
1sM26S9Ftqskrqbk2EVcGrpTu6jyJIOoY2QaG5JI6Nv2QUysZ8/pN591xlRkEScyuV4mexeaJcAR
IF/9ilbF0pvbdB+md8qh7GmznkVZJBGkoz56kTGECI0xkVDcAaYSzGFHlGMg7vLN4WqihanUQcsW
0ZNorqTXoRdly+PrrgOPrNO8UI7hXSoyedoHfAuk4JueTWwhSzMh7VRk6SqKddip7QcKyJrOyJzY
a0sw0ELj++8hCimD/o6jhdXyq0jNqdYe00RjooJRzfWTYrw+RksUkqUrgiOoruniFQ7kNREDotst
rpfag8x3FL0CfzWF9BZH41QCCE3BIRIUzVNeyo9izVZiMWD4rliCAkJhfXzOLN1kUdQAVMUT4DUK
b51p+eFFLP/OlP/3muNaDTFub65NoLutPGXYy18Rk9UTSx+ahZCny1C4GZESdaV9VITilcV44RPG
CgFHSO5NCaZzvszyZURZqye89OIK643P6TLZd3xAVKQsdaK0cv73Bbsr3zI7RjqtCsgbQB2ryC1A
vpKfpcQnXRlALPPtLiAPIm3q8AgcKb0pafFDgD6wEuptHWoUmNJw+0g8W+boxFf/0uG5G3Ccg6En
B5jnHQvpdAUNaY99vFJiHPMrpez0L0nDOPpi8CJOzlGF8pO9QoMSHCMD0rgKTdWeG6dWioWVBb9T
HGrXNQSY7zORpCyk1uTFukZBsX1eHmRCBA4dR4hmjDgfBTe2FrJNFz+60AH64s8tw7pk17kAWEre
G7NZ2saHfnjXUjrTHuVKpVXw0eV5awWM/zfRSYkAs5raicgz+nC0UhYYWbI72KoKdFZRDR+ljkwi
5Owq1rjfbtQWRYOKbUvBpGpVcHd8Wtvd8IdFnDQHh+OU4wNf0feRhgHLc3UxYpkp5pNqxtc4pKBC
kUz3SQvQcNDgbc5X4oHo9Hf4Wdd8bh7idQIRydRSm5YHTuZaiPWRmi+C0Dj3Qb9OgI1oDA3bljWU
wok5oRicqfMZFrOM1/AEWgJPO2tsu9X7f41w+LV/24ZncZe8GqMKwjU7xIfotKr2P8gjxOL7m2OW
Dgk/Ri0ennkR8yZQJuVxVJeb2jB4qXT2TkH24H8grUCZdb+IzyLCjh/ljBika+A9l6Q4j/nErZwW
WAsLMsZ4coSVrXiT2hX0V0iMM1DKQGV53LHfbryCzmAU3tcw50KHJ6M6Y61xV5COO4r4mf8sfCuv
aNckZUzCOBgPcZLRWLxxCTHme70/CRMsVsYwwFVCydjpj0/LWlt3FqpK2aFe3Q/SSIk7Noy+Wzwk
925Y2lY3DBlwItNA8aHI2oTsb/skLC3TZ/JgySLX/QbZ4kZlD0BnA5zQ2dIzN9+ixCyzxRgtERWV
BnQByVH+uF7pFnwlzai3izJZVP38JAYm4z066TAwvXRzQuaj3tSzn3FakhuRWzdq0IChomkQRyY4
eJOrRuMshQFj7viaiIvuT7hC4v/8/kMIxDTTGFR1k59pgDFLwa2KiZd87kIZ5YmM2EU2xLYpljrm
3uFF9od5T0gBamMtRl9ofDzbNUSbOWnCd/G+T+2gT5QtIZsYLZQ60OX66Jea+83+u8baFB683SjO
+ayVeoLmn+DJK7agnXXtw1UArg2KOtiNZ3M922KtVu6vG+gWmG+dedWBaILjDcE9KrSaB1gaWJkO
uirk9moiLlV2lE02R13YUy8vE1jUcSnX6D0QAKNGzLS2en6CSQNkF6inCB8bat5r2RWBJvajtC3B
WItI9EQnzDDJGYNoRCycR+cRE3DkYtbEBR/U6BfzmWynV73J8Qh2PGLk0DtWhrE2iWCiEycr6WL4
2Q9BT7uglbqZMb1eX6bG9rujR2NxVpukrbrfq2qXj9/wcYMn204LR3pO6NWIGTUJsD8hNjjfB9Vo
iknNgF9nUM5D1jXJf1AmU1ELD38hWmNbjfkNusrtz7/Lnl/Nt9lg8+6Elb1ORhIIAOpn0mApVUMd
URERrP4wSQ/cQP4mdagPv8VELtb5MKCohVpvFU9UcgcSZvzxuxn210UcO6+2uBp7u8wEr9PCjoLd
bPs8+3RRpE+wI9Pt6f6d6r3qGWk3WUbEn8WMHzB3PokHCghTZcBTz2luTSP9whV8IEfsliHBVLY+
zNYFRCFdh24QfFVE3hPJjJACq2u21AyglQIc9c6s61USIYfyVOME8uFJOMOrSd4ElD2apMP7AzgK
2MgCboSPQU6dlg+1SXC11qfc+K1HceXrooG2OoWe6AJbL8hOVo4TnFRjDNafJoJIkk7qnM9LArGr
jSAZTZDcpxTbr5F9uLeB/naH1Cg1pk0vCCSk+hkkiDwHyZq2//lhi8Oi8XlUXsAIXO2dE2mKwkyh
PyF807Ol1hB5E8s8aOJvjUuKgeU7M5p+Xkf3sj5agF0dwQVGjh22QGMV8InJSDnBOYKJlz80CENC
gT9wwpPUVn61Tk/XH88OrUgcPSlO1t3AEZucB9P6ZdqDyuZeVW2wDYCIgNnrA0YwWVC7GsGK6+wZ
2Cy7JQCa3USob914R51RXq+OsHVOWWLmoV2EmJ4pmGkn+Irrr8l2/9GGBsxz5/40Ef5QqoWqy/Zj
hdOnaJiuH1D8gkRbi11H5kXebx2owykmS7UQrv/9/8PNsQnX8368R5MBNy26qlZBkQD+es52Slyg
zSYgrdFnEwv8zRPQCVurcJLVbj5Ua6H8/5pwuvuFkT6NP8IeR028hikBEjCsUbzQ66vod0vQX5x/
KjFFzK9WMTTLge4p/RxFooE7FbwlxtZzF/iyKK5TYjRfb3sLs0fMbntwdR5WJ6gqK59gAYN1J3ym
kBX+rtHCwoO1mwuSjGHIeiJRyy/fCfkZwXlIXDGOFrKfK7y+/PnEkYpJDiRVJB4euEI8z0Zbz0hy
fG8dmRyHsEzd37shwpPz5Tx4vo193JZrl05C+EVVwCel88vYjiZqFJUumFUJNzIrQ3Llj4h2o8bE
yIYEZ1m2UV/C96rwdknM7wu/LW2I/Wf0CYXa4a0Fm2rzFGIa6Wb88yr22Qxj4d8C9HK9v6IJJdn+
Q+l0m8do33HRMJ+zpI/vYA2viAOnJyTmuivJRM+XXmsB3iAInwQeqIaPwsQUpb0p445bqyOIDqGr
lc46cZ/rX+KUIGEQ3fyzB0sSa3wZnC8tYWcrDXiSNIQN+d9ActphZNkZjdy0if79VZGC59dRZEZ6
j9x8cvmlwUyvhDZnWAtSUCT82/wcWf5gEhTs/TbLdDTNz8323On4WyuNrDnXkDDihwjl5JK3sr2X
ZxDMM+M4GRct65NUC8V7K3F6lK3wRs2wQsjmtSDN4nDol9XRCvBK342STIUgepVaQl4iXUmHfov+
jlkC6h8wdC9qrU+Iyg7kl1BHiPnzAf6Y3pDWkMJ3W48JM7yANStbhfiCx984DhQR/ZB9mJGlcIkx
LGxd47foaSmy+P3BuZOdjBBnwilp9GZJedDs0HN+dEpyRVINL7XbxdUV6hww0EPkA6Se4NMwTe4r
xzYlesF5au40jghBnHuPlchcH4SzcVPM7nrqQfRaHY7OjH+pMrQNnkUz/rPvIlZKht7KhbCfL/EZ
FgMxkW/Pz2iA0VArGclutQcSN5HxDUap++yxS0EI6mxXYnvbTDQdDsKeMEKDjAh2kpQHebCX+fpP
uxe4OgC18+bThN2zMwHe27rUZIhgY/KS6fT22c+UJ5QNpAJoj73w9c+Vjf+gihv2mZ7aCK778Xxy
3pIp0HLOFkFR/VXbddv+zFqPtMgxz1z6bffCie6fJ/cfypsYzH0PRmDRsOakig1MyPeWNJBgRXSO
F6o5yrWQsOEh3pAzYpx7Jp9QF30TzOnWpTkD+hs45bG0incTrCQBZg022UbcEPj064VwqyE5h3KF
qYY2ranhLNgCBVHaOHyJjBbvsoksh93XP3M4s/wlIhKIznQ9oqg7OdPvBJ1PkVvP4AKOJZ1kmndT
mbvRMp3+tnBn8VPWY36VjTgvLeMAd9yzfcOTVZl/SkKVM7tEoP5bV5VvDXbOKF+4p88M6ohdBxKK
Uro1lgP9gl3DJQye52l+Ab8xigzUFh7lkeHlkBz1IZ6N90JnkP6Zv3XdG5tNf7jpMp6igaKjilLa
PWEVof7CpBnPwx559fXQhE0EG4xJe/uVPK1GrLN5IGhSnS/H0Ix8aEgqFXnTDmeCdBeOCH6eeE9W
SA9zw//g4XjUnjTszPUCFH3NSQe0VwZ2rouNb007oz1+UDdpYSvokG9O8wzOnS24VqGMV4gZBPjp
p907+T8QDXzSoIML5vjaEz9/rIli7Ili7m/PAhqOZOiYx/u07F8J/HK6LbALB2MsqJDf8nnAhxEM
zoma2DtLZ0Y2xNuh3jVHysogPNxAmZiDZPOl0tlRJEmAC4s3B54MYbsLHCCJ9QOrVAO5a8aa7aLB
aRSdjiBpiCjvhu+eZdiWb+NsNu26c3gKEkUnoI47PtFlwThhj1+HV5jfTaSL1MCY1V0BzcyY23mB
uOdeka3Ok5Mg9XbZrptuQ/FZlxTS4maQGw676RqW9IhALpVnrTQMavrP0U2axcXAiVFV4591f3BU
Zs9mLOQZWZ0OMHTqd8xo8ScKRTsNjwPaklAkUyg8aFZyWOt0chSLq6oztn1ExijmJ6rp4G224Ijk
DN59iV0y6HiKCfVYpyf8r7UGKkJJkICiZrfRVzQs0IC0CEK1+t7IE47Hod/TO+Dhtd8M8IsLPubp
zQjY98cnGrzF6LxvXXsl7GFo3V2INA3zFq9RGdla69NcvkTlklwato6ykG+xklDrWd/4jY9r7d6d
eu4Wb3143re9TcldCGg5pGIgz2T8rpZBD2bqSMJhYovwM9FjBCa5XncIOVjOjiU4AQzN/SqeKfQA
5u10Re/xPiiZGjF8CYlGnrSsNcvcnPmAS4Lx3WSf/S5j8XlD+Lso7PWKxISm3bHKq7YACs9NhOh6
tTgLnLll/fThaPBqrcej8+NEHFWXrJOLnA3IW7c7uZjaSxxINVk4I4k45/iJDG21gMtb3DV4q09H
FbWnIcZfVARyTlAj/sH2exY3y2KBi0LbFjRZVPQu4aYi4t+XAq8t2CqCq32nwvKVFzyQgppoYnIM
r+PZW9GHfqRi135S15S1HhVauBSrJ40prgBPCElP1dYrIJF6e3jyncQnuyZeyWF6rsKH2A3ChEIr
7D9DpOw3kun8EEpQd1zuCSxTwxAEP0R3c0Zg6ppHL50sXyg1x8X2rQetlnEsMdt1LnjZRksALB0i
RkFORWSYJQxIEFrhxfwQ6iHG9WN1T7Raru7xMCotlm/V0KKzCfhFJFOue60lBMCp8PaSLMVvBqQ5
wVYZzzwLQ47MYsa560e7d/MvLZZEetWaCwnJc4q1l0Po3SvKqhx4i9AeX19BZxdf3hQZjliaiva8
b1KhHoP6GFAYYPaZgEVFBUMkuDMI1ggaRKpdZEQBjrtRdZ6cHQSvz6eXMA7qRzXb5TPRcu74JVyx
YHI1L2ZDPotwrZPBOhNWCJ+MQewPc697/VU5yy20PUFAztoPhFu9E5cxCqTvHcnxoppEyDjnx0Sx
lDuZkEtbri3ZghSBXjwHR1SH31fvHnLtAVy39lKbX/aCcehPluv/dvsZ9L/H+C5q3ssamWEX/0ch
PZQqA/fymgnjUlx7CiIIPef/4s8ZCvchbCzZWJycLTVkLo1ZC9+zuwwdiIArpQAc++bxM3rRoUzZ
fojEsxuMMvdatzG30l+usxnPDKCMjyHaGmWT+c84Lw3dwnLkc6pA9HDr7VsdxdqgJ90n6sVqAurp
2pSJxITYwMlQ3K+NSr79sMr/4NJB8G72hDkb+O9T9mrvlQcUhAgiDUlFLIQY+yWVFIWnVSr9frTz
otse50ldOEoOvpYN7TWyM04fAlWvVZl3/eAXqLRFDunqPoomIzj8P0b3Teimx4zmGOX1LMJfxGnW
ddSOx+eXYLmO7H3q1yGvKXaEQ12PjHGMv16yh5oc3rI64MuXuXlI9EaKiKjgAkN6koGWlBzyU3NF
OHPLYLmUWmyW6HHNPRbxyc3RirskmIg0zbcqvGGOUqO2xaLqI2KkCCuI83DPIsNM3QaliekvFyWw
J1ogpPywwpGUqge1pI90TCeKlezeht6KvZKY2QivLoUW7YEh1XMdxtXRehVVLAUwfyj1WlWHKDqK
9u3n8FjIsUGyixKAggvhnDSNp36t+gM/hU8uX20CfRJBjQKyRcaiPu4Aat5ROA0n9q/N8/wYbJIe
jDgMUtJUkE/l5/w/TL7ioYWT/DR2JOXYu/fIlX0J1fZ04oNjGIzoKNH17B6NeOoVX4wh5QnKN71p
n0TxNqVqtl2l4zTTcpF/vZFV3cB10GKhuKCR+QODc+Yd6FRvdLtpeXFJJ+vhzRrJXjrkEv7rFJjD
RypUt73ugigiAHKtT3hBhwxytk5V2Bhc0qPxiQ/Vt8liJ4P7FLjZr1xtTrW5+Bm01Hv97qUQT/qL
691MwQMObtz8j8kDyqHCjLLSO88l00P8+fK8pekPjOaBTjP29EilZTQ8fpvgHIzMzqHjmRqtKFhD
rcZwF4dRYo8sd2EQUIgy9qD5rkhr1Q0+sV6DDNJDYT53K73EYlTQlYZsKi7b45ki0d4N9BWq8gIk
smYRkPQcsdFBuuLkiSr1nKClqwdo5SW05UXVWdPTv0eqAt0W9JZIlBn2KlJ0hgDYfrUd2f09LrBk
6CLTi/J5NaYwpjZYK/QiTFqFWFLjAyC8sj/YK8lXH2IX4etyOir6mscfY+f6oU/1WxcMxtGlinLp
uzVYfFDR8Mgo5kTPidUmnQqM1Zq8FaSXSof9EToKofCVq9vmN/+zHsAHwBEoXcZS6HeynMgxPfco
DI6yX5f3dKKWs7HftEdBBNjiV3o0aZP5/7v3gb32T4/rN65HWs0XK2YL0OvswJA6/LSOWM8f+7uZ
3Trft7cUmRpPV5EdrIS8AGSW98wDW7NyHkdrefOmlLzpSGJmOWxwvwSEcutkKfryqL/USYPc5Ex7
IxX1cMH7aTJdB6Vz7ISK7b5AN5A0jevu2ZD25WDtIeJod8t6WQtVE2yTiot+1qmb720b58Nt0CSI
PwaZ+mXbuay97/cIc04A4Xf4EZ3EZYxTe6yRRhnjGyo/E0lJ75kBHLYUG/txI2kSEZIOW2CKWlAG
YyzrnwX+Wok9b1YmM8pRWSs3RfeCgh9qfWhl/umZ7WvFrWNPRkiHm31E65QAXpInIHHcKLTvtE2n
3XX3X0PDCxlVQJuHggSM5eHkgIf7QPwv7Y7ma5ze3GeUEFxlc/jdDGc5+HqU6t5mD+msIb1BvV8M
10I+u9H+AsJROJQPdKL8/LohIl6IQXe3FfdNCetFdFAf6qcRbTAGJba561lLkqjsF8HbWjbUCyrF
kjsv9sp9VX3sZAB//oPPIEc4eXUqiW2NW2ugRPiZGbIH4HNHeCih65RANZDWW+8AItulYBtjym14
l9jL03xbPwtw6yUl2qjCy6san6kaa2LI9ae8+xR3ZfKT+vdAE2Jwlgn9uP66EdLvPF2Zs6s4Yoqt
x38B9G5UCezGq3C9W+1xec91nuEuJP+yAgFjWwDOm9d4Aa1hB5j96kS42Wz3durcItiyyng8Asqa
DKAN4r+z/6AgollQvt3zAOpRD95fbgUEUTKWnWRAoftqlHzJPTigAQb/RBWaogKLBsBUFdu3h101
NtF+w6eI4EQSWul4dHmjuDR8GRcX67CZ8zHIW6azlvVECv/Racboq3y7KgGBer3y3no0HlAhJoGH
T5j5DANEHHzHYWiAaIQ/nfnCd6lrUPdcPRWU1j6SbscNymfv12UuMCBBIwtAT432zQQ7NRiC5af7
xW7NXTxnWasixYh8jSIEnbI8S+X720qvfDzdsAcQlSiIw+85W0F6BUz4MCUxIzIJp2ef7P1X91mX
6T6WmjJp5KJCeC6+bXxmuxKH2RWACwg/mbTOXQs62TbzsbeB1qtdqEo1wwJfg/Rqxj3PlXRFoGl/
zp7rXeJ1u8M8OqmHhRZob/JcaZ3x6BY0PmDt+6YjoA+H/nfAMzPLHEzLSM8SXhkpccgpzIaaY8r9
zyiwayj1ROybY2zugYOWlNS44ePzBoq9XABN2rfM7Zxwhg7YYjjZf3bFA0GlfHx1ypn7FbmPV2tx
Hkad4VOavysvbIZpmma6SQMA+jygjGItRxOSP75CPsHFW/HjczgGRFITF1VeWxuRGrg2dN1QxWWZ
kFD7fFOqwxRFZh0oJMHEDXLhQAXkJAgqjsR1aiI3ALIQ3ThJjt5DUGdw9sIrfT8yao3PY/fBbGC6
Wg6XWOrdgAe2Vf6eqiZNrFHyRMME2myhuNBJrb9F9Oxbvf/5GEl2SCaOxOyhoNR2yVir028FQYJk
7DP+xQGBnpaoQyOcN0clEb4gOvVS/N9E6Sl669FpVfj6j62DuEO0XKsejqcNAVxBxSlIgAYO5DfD
yBP6nKE4C8z04sEtDXM4q28b9AqQmi2z2ohNchwSrDD+euE+dUfRti0dfSYQmO6yDz97I2mMsP3H
8kqll8euVzQ4s96DuFf14q7kZKy4pO/D8HRIWIojQaU1cvzAOe42xf7GWwskccDrKs0jLC44xi1c
jlaHq0JYYy50s0ZTyPyLsAappLjrxT7FXy93jnhskfB1NF9/bCV4d3/skb5+yWkb89dBJo6meodd
hMIm2BTnbtDQIpEvf+rBxjW+gfHyIbbOgtHH03MDb4IGEolNoLuOTuxCd8vc/z7X9a/WwzCAVk9u
2Sv1hZprOdykOrfUZNPMoFoPGd9zSSuXeDKgmgFB+cLZ39zlxJ5oDm/tL8D2HT6QjFUiLL8lxbOR
yt/eFu4dNu/wNwIlqUNUwYNTeWdjzIi0I9j0+8JmU7QQy/D7Lyz7JViwlx0yQf4pUujZ8H1ahQYd
9t9Rsvy3rnB43xsDI5Gev+YyfApsFha7HGLnAPwsrV+UrIb6/swl1B+MS/jCIEx9MQIFSzY8v9se
stAo8gcWHUMVAo7aWAqOjqsFAog2xDVfshdWD2Iz5SIPukXY/z0j327UCaX+rgvfAOHT1g1kPcwX
hgaJoqCncmwb3KkGOOmqg92BD+cTkiHrSGKMpp6p6XjX0XJRRBPIAbLRbrEl7Jwlb9Np6gz9csIL
HRu9CTWSvH0srIzRkp9TGAgCKjD0iofXS5wmhLDlZCNayJ/oJZtzH0is7y/+8R8J91547TYsVSQr
9fdTrnCDu6aQxMg35jfkfsq4ZM8zV7hhuI+0zKzvp1jWSpPEyUOjKCZuCjB9fZZpJ11KjMRLrLPS
U0SGj1Y6d3mhY9i2pVyaTUBHzQ6D6Anoybja2ZWYxD1khvT1aP7oWdj4Ifx96M1Y4PyqOyxHtnWi
x3y4pYx11yh530yR/qw6u5olbvm0Z2B3Q8te/2eaFMkZdaXPu6Dk37tBSd6k/T28NcuuJlQ4Aow3
xTXkdPkL438L2ZBMiOaEQskfZ4BoZonHjV2/pOY2qrqSm1Sg5QfN5Jy+wqUbqIaZ0lHbKQsQUOtc
veAE7oh2oR1BF+oz+7XXJbNAr5/vb0CiFVhB9f3ZozqyFYZ3DZVSTVmwA8DzjtBh9cxtHol8NzC1
zvYVuDKVZ/yKNLH6rkrAH7HS2KhdJnaqXg0qnsD1TBUDdGgA7wbfnMi4W75BuhwKl3eRabcfuAbo
nat1dZrQuQWImYPUtATARlyzPe6Bn4RSHJcm/0tQ+qn9LKrQX6gGTpQV7KVoCMVGwGzuH9qGIpv2
1DMCGND0bfNz3UnAUJ/FBOkld0I4F5uMgU3EhcxbF5Zqf6M80UolOWZw+mQoBc6fP7taJc/XgEPE
fdGRqUc8gAzhwlFoXnHE+Z2AcG1LJQv/KZDePTKiBUiPq3ztTAC4obDmVeoU+mFl1TkjnUBX1jEQ
aDw7tzywLF0JAJOCKlZlAB2ACRTWc/Me2M+FozVgzEX+m1RmmI0CnkWqAZZ8oEX5/f1Z8J+9k01a
wSoCDv6VKWOKhZgTTK8UGo0PZ2WVoA7VUeSWfjqHWrUZogrP4EminD0IeF59Ki9BF1WuWtEo5e41
PJ7aA5re7ZLMQOmCQVDKNq/2F6xBoNr9zXGd+efgp0+xe5DqawB0Nf4G+ZHCQnla3ITUsbf8CINl
/Za6bP1pzh4vseLgLpqSbbK/4vsO+DIrCDtMUxuGt7fLZn3thy4/Ss2u8mcgxARao/S3RpvBTI70
EPpmSCNC+O0hF7t7MUjE+/5Dp3t5mEneoPl8JFWrwY9SYURPj5BI34kgh82b/TXjdzISpTHX8GSF
5dDdBdV3RCiNdxwjP5KJepoD14FhE6OdlPQQC24BpW0gOFaADIwMDjQGIyqWtSdiUHKOiuibze7t
IFAumhI8pTvRrsQkhmgu1aS6hGU2AtKEwsxhl1cS/bY2Jm5qL31P7b33YFPysafu0rGetuEj7iMF
VzA9W8jiXBWsNvm8ozYwlCoyyUGIGY6d8db3WHS9xrgfOY01zg8U3f1tIdzFARwLChBR3drHbdxK
Nrr7xvxv9RUB6UblL5zfTHiPZMrNudRZb8Tgg2hVlmQ8sas1buwhbH/vVOMkUwCa6FlUbaTG1XT5
Ed+iKSfrw1V8wCxFy/qaEgTts2BvR60ORXHXGBIRhKSoPk9hhHIl0VSbjb3535x0xuF58Z67RJ2+
/rGesqjvqQCmta0DVVmCRGa4kjguUzV2bO9n3WNu8ubzSGaBvFAIGBT4+CwzRYtNFE36HRLmdUmw
/OZhL8wLmlDHrUvLDavMnkTbQ4TMTqOpXdQMO4kaXssxy0/tzV7DQ2WOLXI7Bc6Vs7Pie6hxXqgM
CquWfkRXys87wRDiYsRlHVB7kw5VQ9PtDfywxae86ZhE4RE2tCpcF73GSX16abN8vHvNrjqOUDmh
QjV8FDv3bNNOo54lRXLlEpbDq++pyZ1tGVqkjFOMrflT8LEbxv4AJUhndSWXQ5JmCgmsAgU+OHlA
AfjXFFMopFhMwek8SFm3uq8mU3HejAtCGxXDjWASTnJ3v6SGRmeHYVyEZ4p3JUdNNBczye+anT9H
+H0gAnFdexfnV8vg9dAtElYpGaZI4e6TmSCpD6ZVNoGjtCekThnSLrQG5UYOugBN9aT4vSDJp2Xm
pNheqtPo2g20ykZ8JcwEAz/HBr07ljox7wixRwKanHiy54mIG01kuAgDmN2RuQ2tBnQPS4acaGNS
VLIWwyUploJGyy50VuDgtxdvAq1huxsgciv9xsI1xWLBdcqDYYpA6avRbGCWs+jSFBXQdoO9mnZU
LrAazip4DG9Juq6npMDQwzUsqD41t97IEwBbYE8E+y7wOi/IDxXSt2TvpArOfQXGLVn+vcsHwzft
9YNxtb5xy36WlDrB+d63ZLlmHhJujplrUOMJN5Ukmnh+R6TpWo4yOkP8G7R4tGk1SnsfXgki0Fwa
NrlsQlP/EoJ49C0+HwPcyec3Y65Ts90sthofUJFuP+QPcytyWuA/ly+OZtBNvFXXuKY6lJYKyTZ4
bltauKY+LZz/9Ftui/KU0wwZgG88QMWe5mcudKMee6W5WPNZURCN1E/GvsmMfDPhCn17JfsdWSeE
XX7pvIdGR760GaXaXBOvu8ngregvrAWFNWP3PicV4s7+eK0RMZ217ACO/0uJ7Uo7Jcmwy8UupCZf
tFcDGUu0Cpxvob58UaNN1UO9xAq5chdoI46jul/0/pCr9J80HQjChOPnTJPURAzXRW/xlKm4dU/P
ya5whMXhr4zcDYIcKw2/rfsAwT3p427V1H8ZfMYFQIVg1DYFFHu/DMxMGomTTEVZJV7NS1GnV07o
jrAj5pahvrWY0q4PqxGLBs27L1xlgVdA+UZaOcwIEjDhy3TG+exQEXfhxzN+OzenCdtC/kpLKQMk
XdSLDjYwSg2yk6RxJPdmHvMWkfrV59Tf6I/s/4pLXP4Ykno/gXk8OqXH1afughAvGcNAWnmtK4gJ
iRVm5sWhOq7vT2LPbkW8af42RtIl+tstKXGu0JFY+ovgSC/asqUMDDXAwUumPcqRkmq/9oUZg7Ua
9sbEPUiZHQuiR6xfpW/pZLHzQixkzT3pWi0QGPBBUOqXlqYc/bqgvrudvEpaZn7AMnR/EbAbZQEH
89MW7Jbc0LgeyC1ZT70xeGrFu6gLHz8jDPZEMqM8fycfxGgLIxkimoDAXknJ/pchnSaOCGVqF1Dl
yxF2J5LHjhLu0cY7rHHQPrpyiOFANweXx8xywfsAH54dnDJaEPeVvdtSp83UovvTMNBVb5V13BxE
MjgHSx0Jp9bUqrtcmh4X0K/rlcAuVO7/r13RtLm1HOIbnl6mlx/+ufSVEU8U/9xhbIcBTnMVk9hu
Nm0ddntaI/zPXC/oFFfsIRlQZqL8lODBQFxIcCHQAuDAup5B31dyPDnRXrBUxIoMWnaOmGALtaAD
Sd+U1YTBeg2gE1dVBaon96ZBPBRX+AQ6jIRLbOS0uqLEB9/Y+BmDSDLXHICQ0ShQ3nCpd7p+6BYx
HCExLw0kKG2bXZTsRTCNeXwM5RB6pT7AosVyjsm2EEzI9bgTQiyaCCcMSINeiYG4JUtONlEBv3eJ
quOUTc1dKN1UWWR61uGlImz5cRpzd5mYyQOIplpOFaRDwTl8W/il4t0MWhzuho3IbWpHYtqCvokB
xjA3JWMa2gaHCwTyxXRfnJiHQBQjv0WLWjjyXU2j8s2bzISUITU/GHkVYkYID1dE1P7fCAp2SieY
UJIL+TJ1NzKLcYfejPMyYJz4G/ecL5zg+1/nvooahKQ1lvELSYUC6TjL3Q5nDQUIdkon1boqzDte
s0Xec68XfGbvlq2pY7LsQgSn1MxNXwmbGXerzG7ivvCRVawwqez+aBUuz9p9XHl8fbDxmzHFe4Al
O7Gaj6OXTi7kNnafbTVqpua3mRnSpArnXNsmdaRV1az4Yow4XWgleuqebvf7p9YU1BgPAgKgqMsG
ATPN1qs1Vbwde3i3bpykwWQhVW129ykYm6INKYG0X9Wn79F51keVcnvhqF1bhx5XB4K8MhmzIUp0
BMGB7+1QUMrQomO3TlbFVdMuiA5JsD9gZnt1pzsWspF0/fNdh1jSVleiOE6AsrmIhzRI3bwgxRr8
uT6eJFAmppl2ZgCzOifsYQz6rUvvm6IJEuA5ycZ/bQNEd1aOwlIyBfS36UPLhvbvnHQt4msz1AeP
PKGw8ARDHnAfweK3fzA1icUE2JMSAviLjNZA3puDEXsVv9r036U+AEmhTp2OLtEimmEqtIjkukPe
lTdyQ9NJJGY3I874a/lVv6jYd4UVAitOrfbjp7l5OQ9pFnfKXvinePqljWXdlKMy/hfIET8OFzVf
mZrevzPZ/Wi607d0jSqHShv61fmSr62oYne066VIKVr41JcHJsbb6OroWjrULkgvRuZww5DhnNHX
k6C66LgdPI+pX6zIxrTPu13SFhMJFmXORPGxNZYeg7yoVsr0FUHN9iyweZNW04K7lVh3H9IOQAd+
330zstd9gicVpWMjl9GxNoALqJySjLCfi82ABPgW74jkpYAwXN6TJMTGBDJva7c/DVK+mdiFFv7q
74nYtsd54reRBUGm1orcVUcREM/EnGs/GlajvWXi/OnuzaKEicQntAnEsEQOwWiyCvzQOlYXFGiI
7RE8M1k6PMVVqM5SN2oEoGlxAQ4LYVvuSWlalvYmMaNWrgcgd7SXY/AlhdoAcP/JXAFkyXLlnGXs
iO/7v+S0eUMty99FxrJ2qCwkCtpYJ2BTEV4ij4B9s1xJSbnAGz0N87OH+l3jCxZaR0/+a2xnos5X
DLO3HlNF58UfxyNlCxPxQcfcNqi4JJGhx52Xm32AhZCkbK0JfSmt2CVUqc//j9qe6QBf2h2annFl
Id3Lh+K5NM5NFUXe3AMfFfkqH4x3ctBJ65mB4FsQl+0b1BzTeA5e5ObEKKwEsh4XaxKc/1R3G/PY
BujMAwJldu/RMj/WTdTmbCM+nMMbYhJ9ZLYoL7akaDpiyLjWlYzMwt4osgnd7dVrrAh9xFcQnvRh
z1N/ukkcJAwmg3HEyfNbPkjw1U7uEu0R9vnnS38W54c+9gBf3aCBjyutKOsLyNiukaRVeAWXxYjb
ie2geVnHUZdMNGjhSB+Tw4AM1qWvGRpRr93TmzUwmJ+PA90gnBcDPqCPPjsCZ2rccAIMW3wWfuIQ
57HwhamOK+QsVteNh8o2dyTW3PifZ1iTyG070Ej2BYzhmk4Dn3iqxm/3FuBrhu1G4z7yGwyWqfYh
ktphrZQqCwIvR+hHdJChVPFSj3rvWGsJB05WXiWShz043CDJd6Yy7M1f5x+DxqV+xZZp72yRaAaj
NSVroJMBWxBoLGs11p+N1AqlMwQHHn1GJzDF9+2QRGbwEq+RvduwdhWGnQz8z4/WGddQbzybM0jP
6x2uApvQs1r5AqsrVR+IsDdNr56e7LZbOzVEMm4JI22nOBxY9gZQ3m70Hlwjk1wTASObc/KkMnO3
pSzFmxA82Ku6r0nwG9w4SnqIOACfjPxiy3rTv2MJxMVnlYaiO9714JLvY0edefrAxyqD299zT9BQ
SfHKhTjN6N+fMO/L4qrSKkk9P0q7NtfAfaVN9YN5XxPI4iDS+nR3aSsVYtu3ieiYwGWx4MU+Ajsf
n3KOevAvJsPjFeuSmuKQxN7WO+kJ5Gq2+uahdTHosnsuR7YbpAXsmlAZIrhkrEDe8yE79IhsdHOy
PstN5e8JhgZ2Yi+GaTEOYKdttGxziKLHzSzEgMxECP2foiR1imOn/mK7BvZU8lUSed0TQ0Et0vca
izInc81ZxJbhX7/d1fA7fT/6kWoOKF05NIEUr18bqDoJt20jb8cMxwpK+Dx39Iyg5cW1hsbEoQtL
6XrMvzD7qwPF7C2SNR0+zzJ0doSnaPagAOYeub8TkzYocB6hO2tw/Z18nEOuYnTAJ8QbM8I6f9Xj
Dbr15nU/z9UE7y2Rdrog5Kxpna7LSapbjFsuuWWSpxa0DE4qPoyRw6y6SEGkQxA8Z8+LCb3923bw
q8QC2ycTjEyOGpeZbv+RMsDK94+GMUrxpTDAVI8Vhe691BIMZtCJZaNU8the+/DlLnLhDkQPdabI
sUCvhv4ZD0xL5HgIIBX9rpisoj896Gd4VFVOPaKGNzMwg8MEX8vbPz/PZ2YgxgOnJD23T0A3Cu6t
g64qi/mo0jaq9yUMPyqUz0yIHjV2LxTPR4K3N2+npRlvtZl9zbXDKRGAXZTp/XPfQMNvMLSQsBl5
xFn7ARWbmpiwydEtez+e0v2ABWahePyU3T/iPtKWtwhRenpKCE1olNaCg6HYPD8v6B84tIagoija
nr0b986Ly2pDT8hwBZ9s9nuKmR445pkrmYvOp2ZeZS2vl/eGry6vExXQmcDdHkLdxrGibMtZEENK
yr4CK8vReE3WubJHzTtXVTdKBLUkIRfYStgFdFPmfkLkpT7otl1Ki12GDqniCTjXY+KVtSl+j6wp
difLN+2gyNq1Bi3xZMigGTAK6hC0EfcHy2TqXBq1HXkGycXmBZ66CPXSG+YFQgyGXu5RfQzYI+xZ
5c2RSaITpGRJf+g90jm/g7uWkyr3N0ZrAdFJ/OTlW46oryrOB3SSY5HQ8dOmtc5Jik/D9t7ueBcO
pJbOUr00m+F8jHgJo0XOMXc/nCgMZynygoFTDmteHn5JbcjbgJVCQmgMUpC4dinrkwdhIhB7C6RM
8kCdKfxC/+YgggT+bnlE/SK7/GYyjXHVMc048MC+XMIiJHhxDbtL8YWNoO/OBxWydov070lyy/Dw
iHcrv5QDGQpLRrjdXlru6gsGVPClXV+EsHk1vjzGuva/YfjU5iy5L6JfP8LH6xiI/zFc6o8CgqV1
Oypm06849z/WhIeFDuLI8Ysd4w4N8+FZdKr+b+xsAmWKdIW90cYs48+wmuot5GPXROEvudzHer1x
Aaz90JfyXU2AMbWfyCco5nz2FUODSgHTgOG4J/zoSQDxwOqNnQqc9rXHhB412+Jl5eqPy1XipMZu
TmMOLFOr0klVX6/8ygkUB6uxwKrxX5hJ8kYXVAvu3NhzXzC9i0Qf4mzJQj+8Ggp2HAt1TaRYQDcI
h8/uAY3KO36ibes/mSldZjAXvokWFFHBCI/FO5uCw6nKDiCLijiihTr1eBgp16c8Oo7IlM6wobvC
sU5Hcg5wQ50MbgWeQbwZDiz9Nsm+BD3FRK6Q/7eDENLqNK7HX9syghf+wgDEexXkM74MAh4sxIDF
WjQyACLXPO0Zv92Cub4o2EKA7we8EH7tKP26rPpIr1VNABG+xg7IpY6mIx6J41HwU6YuUUtYrMlm
sq0z8XvKCKpY+EXQ68xTPq+Yggc08T+USGwe7SWZ4w3bAAizREQBeHs22i3kPPoQoP14ryibe5zC
6xmRJDiaGsHmUzBJ7SZsSl7EumYJfYCEwXi+FsQKrzJhYKBheps0MiQ0C+Z3Fao0IygRNziCotXw
oGM0PD7HFzNI6WpNNOfU1UOoakO51FOVI5NTZN7EkPLbi++NARvqyFmBiJ2ElgASrbYSYMTkGdHQ
1rATGXF3dQHiipmhJxDcxLyvU97zWfmaEnNwacdslr2obt6OK44pGq1bIRyF0/2TBMxPo2lEfmCy
6XzMXb9jqpFpyOMUlfhyFvskOHFFndfEilqFj4MCHI2p5LeHkafsVvffuoXvVFGvIj8tmx7tQpZm
hvia7CqElPsTjj5k+28YzrafvIi2c7rLaD1FdqFpr4w21bSU6Uy6bLfPgWeZkpOW4D/3EL4OK8Bi
/jMTKvYy9XZcn7gp4xcmky1TH/4Y80hSUU9Q+u70NjWMaLc1wzMaY3dA9Thv3AIou1Xr75L8L/gx
8XfLaMHKQvaFWfZHMxn7kM6PaHsQ0AGomd/p+lxG++TGQ+xfOvGxXvh1Jptsi3eIfmb7sfVaHqhq
P7785BD7qZ3ty31AcHqEB7W/FFOj8HuiuZLjSz26eXs1PkxhOsErcBxjAJlQBlwZFgnng7EYLB5u
N7S1pKhDpl6Xm24KNNU2l5b0ViVEMPUoZo6aRgB0lxWH+shWL+V2icb/7uUVWXve5DmU3SrBdwfT
Pt4dl0dbD4ji8kwzD8CslC0JEN8y/GlCQEJ6Fv0OKpi7nrszKO4h0tMP9AjAm5OjrTSuE7TOTm3n
g3LAbaWjtWdNOQIlMDmdMDyT694nSNuJvNDWZxsa6cq3zU28C4vrYZwTmeAqlo2KM4OlIAq5aaJ5
OILatoxHB6GNb4smRGg4pzGL8j59WpeLIQJ0sv7mopJcbPyPa1RyqH/BqvYZ9N2GGnONS/02acuk
XKPb2VB9m/bky1xVnwVKw18urXk4P+Liqfq9y9Np2HX4fHMo0gv9CKOvAzRGI2f1U9q0xJyECTXT
6YmlA0O9+p9ybbrKBiSkbR8UpUpH+oxo4S4fataaUC4YMkk39n63ZFvMiH1O/r2wXiGv1kU/+gsq
kpEVKtLhY4JC+BwO4AHhJi3CodEZ1bG04GNIO3QncEdOqBAmLr7xieTxq2mBkwVBGCDACKRmwqjH
hv9pLRePfsD2hYDop7LLeY8v6Sc+/7/ZKNfthvmWHhmWJfJhIeJweljQdoFJ9AykTMQKD/mDA6uF
ksFKpsyxiCuscIr0zvKA67PfyaT7w9wn2M0ohgoGNA5e7K93lcxA1V5wNVvpN2SZ2TpXySW0kxpa
V1TlqmxeU2SOttA+/rfC19Fpb50Ger7TocPkL0a0sK94tUYYmN7f5ZLzMMlvg86eB/FVl3CyfIHi
jq4cvwwChJctVXB610/ubEG7aJ42B4I56COMsoFRneBRyPNVygJfIV75tweQApUrfJVsuYbO3ZC6
BtdBN48UTqI722STKqimzRJeg2oHtO+aJSiK6/ngmnOA8XkT978YAnRq39juTu3FTSBBesuM9Ieq
VkPnaTki63oX4VtNyFQ3UMwDw7ECNd7z8K1SNMa8O6+fZHgJQNV1i7sjnPQ8N/pzFOoIPJB4TrbH
6rk3cz8LX3LR2+HgLvu+70aYfOTDJD5Jbl3DbDfrq8yymce3cZoye2xfR9+WucTwKqA99nEKPrM0
nlMygrDBEgs5k36kxHvUpvhkKk0WseoTf5FymEEPWqBLpHKPejED/CXD/oMZcDf4tPcHWb7WoRjp
yCb7Z9+ThytrhB4sfOaZvOnDZO2wQGOrHKpT0dF8H0dePFnj3h/LMOmVBx26L4Ckx6AS++WSp9Xz
kRJCMbXcoc85E+qNWBKcXDPf0cI7bzApc5cPXQ2YceXHvjd56bFbZ+4J4E1G4fAl86pz6w/+e2z7
R6R6xHM6Ot14BgKGWmrLkPsHvouD83D7cXJhmur74gcRIRlehyx75AgigfJAuzcr4QOj2omUB1Et
Sr8hOKTRnG+cRuK8/zsc5eNkvFNuwDjJcYPuifBm0axJRNZsbFzgh84EdzUbRB/X8gPlkhmdhBLd
Mg1RsWK0PE7f2rrhd6giORuMclxfPp9ZDabbI75GZiRRUc+BLln3ymFX5Rhqfa6ELorLVYMZ1Uid
cMzfRuqVYHZMVmkUyi3PJVnxxzFSlutl+Fo+fmPdPE046GA71hvDewZik96AtIUzE/NL5C/79ywn
LJRnQ3M7nVcZv3Z9EcEyuE5l1LZNpZme8aXZq38P1wPf8+RVo6NmF/xlNqvHcQt0jGZHBCIDWh4Y
eXx+Ci9Q8H3kKRHwJfteOqyXIuNAEFB7tLPpqfk3P2hWSXMgDlKWIAS3QJ07ESRCyQoue8mTDGmq
/nvdNTqeMqBf0LweqFgK3ZlS7nEbGQuTCAa37Hl3ahI28Dm2nC1tiYRHweCY6jPHLjSGR9h4ijmI
99Qv4P4CR2oJsBYFEnlPS5kDus4rOuWCtEfqfxgJs8u9JqjxrVUe0un2A/ODucRWQEt5vmppWzgW
z1agZBmK3dqa3jKyOB1Tbuuo3fm9fdLfsyfCTxWG4H1gDXL2tF0pDMd/v+Zxsm+DYec9EQrpt5tw
cDtznFDZt3WY6EkyOMNsH9t4+buho0dGgYbIuH3l77YsxhpAsi+Ph7NRWCd7eyKaqMllSU05cUcz
k5YcYVXR93OF0l4ug+FWAp/UTQ8UUmaM9F0SK9qgAFeyYezSPxNilNxhBnsgkJnhlYieR8ZrBXuD
4GkL/shSpGeIxeuMC4fXyTGcIpc0lwgcUgObYlZ5FxgRG7c/k+3KfYAvCVQVsjUoArQa7qfKD0g5
kdLuONlzMKkwCKztvhZNevYcQ+ffFPZhzKLfSwvO8cTB66IlvKBZaPt+NaIERUxEhNNsB37LPjFP
DXxRm8ZtQ3lbKgmlkjjkSsMsb1I07yY6h10+RXfkBw8hrC3feKhrYz250RSRJa7yVN8u0mD0X9Ou
adc5qvHzpF8UPSm4Viw7ARIAt3eGEcx/ARPe4hvUsRfdgA58sEQ3GfnaIN/dexIaq6HuyuZAGXfg
pTrxJJXdre9vk2VtdylgGpeVBD/h1DFfQ44ir+C3ezpDPZJRqGp6HzISgm4EmlDx45m8zcvtUNzt
ngDnlzgA/ZlTNjJ1o9TcHE72+fxpcDrzL96qd5XHpjnKsKTHHj9UmRExojHhrfRbIkGfeS9TwCZW
xIDWDQTmL5bNleQs1RfKJXBoxAWpohGdqNceKdV+tnoJ2afsMps8zBmZJ4MSu+fWITxPUeOkfoDN
hNy/1Dulw94acKdzahCnGBYV7GwbIuUqvrRrDvW4QygtvK8aUZuVICB5qBN6IdNTJqXoBcySIMqt
uK3rzLoV+7MRq12gSDOawaiujnlLvHDTOdRaMfoTA+D/0IhYIl8+wRJ9opbqcGqPBPmHfM84qRa1
EV4OvEDU2BPPvN6QfxUQFv3Sshs4mKeug99Z3dJT/PUvUshf5Ge7ur+uAPFROATup+SV1y7EYvp1
u8Zx24XVhP57jY6ILluiKdsTcCYggLqhO+ekd/z3YJiZDV3Q5peoSHYCBVPd2I29kMBjXl/+1/66
NhuPRehKRaRP61ob+vTPAJCCLBEi+rwLZ/UNMlMmIyszjoqM4A1uBZC391vkOrD0aUqfunesfpPZ
pKLuhMT0EVzMWlNZoLvgLqusf+uRKJyDaJ9PXjq9p8jNfV233DDZHraM6VjHroFQ0AucbuZF/FPp
ip+pP3PWrIjnowuwnbiqf0GlzUkKKMs+Eq3IEB1R5MeEDu9nnKLPNuhRcIaVOC961ZJK6q7ukahl
tP5Y/ASqO5xBndAE7ik6krp8g+n7IqbehItArelDXOW8JmGHN4/r7iz+Z7uSyLgWfiKgUr4HMylH
lKBN4G4w0Gu9LhFeb8yQn41dTgomYJvs/zYjyXm4vynTXo7RD6BS+AbQjMeksf7P/ywUmZstOjb0
7CaEToHBPSejd0ifbUKeUBtDxgvwv9ZJ3ATql9tg0wD+y0teDKMXx2G+XT82fVrVavJ8939IRpif
RVB/jc4yab4QzMts6T8f9raQPfO0J4+L02bWcwOr6FszmRA/ltDuHGv+ykY8jwFL/fwxvsmUrAR5
yQUcqAJNGoM18iYoN8bBxHomHDdy4fJE0APyQQ300JL76xflx+BmwJJTMy0RpxKFPagb40XIhNQe
k9pIDF5fLuG+/NL8LE2WWQfUgijXs83WMn5CeP34ul/hZYNrMCcL4Kp7SF8sWhJgj/DR7usTErOh
PSDXqXBD4RwTma2IWwRABZKm2T+rfl7Ff4x7dS6gijC7556tYgyBztgu8GYmcZDdxPy/cia0Cadu
P5vCvyfmc4idaL9BceRnktzO9x2/07omjbZXZIE3uTzo0C8GqtP2vacayL6z032utiySG/1+Sk/N
F0whWPmdKQ1UVZEtDswkOhdsTvl8HjeuAXFJXkXxs5jtuKj3ogmNcl1dD+GEZREy9bHNcSQBXEWQ
6ydnA4OLj/VB2v+vRrJSFdcoqEpDSJNrERYeUnlMZLiyYQMnMURA2GWMW6LFoN3pYCIvT80wM0Cx
uIcBv8a924EEC76jFmfEKD0hyabnFY+NwXammcIYs0Sq+vetAaGqKKQgnTOyyG8P6yQ4gWc22iFr
Cg/KqEdv87W/GzAXh31ePO4No/oi1/ddkCl0tGiEFkVByugDJWbd+9BpomJIhRZLqgDqLUVX0kaM
ebOzFUPgwa5KiuPpbJzMUAcAYNfkx1BFf0GG+C0Nu/S4QBikA+7Y0eFz2ilsMKSbHKZp8KtXLUI5
dD6e8rf/Z40gkYVjHNw4utZlVTEdljiqynA36KQfu9x70Rfq8e4x9FdtDOF2KLP54gCunDtk6ca0
HPm/k2khCEXLbVQEqM8qG8j6UDeEVA3/MHgkw6fkJX9rTkAzLyWQo1bvwdCl22YDro6IxjYz+8j0
aBun+aAzDXeHaN9a5RoUFyZ7beZjyqOs7Jo/y/E7a8HHssPljyq3kJn2buEi8FawYHo3eT7r7+5T
TICRXPDIyxuoWneXN9lAd8oe+mO0n6mJOsb5IQ5youmD7pF1DJpHtrQj3a6lLOffn2AFrMVZzcLq
+4Q813yr8qalx3mg5LzJj3hvJJpn9ufyeWyySkZ5IeVE37EhGXYDkkRdHThZAwqhHDKI1eEncMyE
p9JENpyiUwEEVnlMCZan7Xq4ac0eK6CQRD8Juz5tHyDc1UkQ7nR4QcE7bTYiR9MR1ZBGGPYAGiib
5nkoD+RD67vRMa3PUaYa5NCQmh61ioEIpzlXPhUIIFoT+HOx8mGtDVNInzI93u+HAjTUZ2u5kSbk
xyY1dLEUKrMK8E5abdo03U/alWbKLtRqvohsEXR0hxiWhxFMkufSQNhJ+6XydkhQx1cC30nVV228
wcxuONdbOhs7A2blcScEs5fe9pWW2buJ7QmEwxd/8s+odPKXZMhHlojkiEmDlpqnIVc6ss7VeKun
gEnmZLulr3hXsUMjXZ6X7mnuVY85QAZ+Wq4yK9XhsnE5tpgNTb1Zw2hknl5OAlk8K51kmCT7B5WK
m02DeRdGy6ztOB5eWhoMUW3BoqCQ5KMoaGFG6FYywy0JrItyDJC32dnpiAxPIGbWnxDa2teOZG8s
G0oPlZJerjD6gqp3d51oi3hSsNAff9N/xYYooPKrPp9QRyCG6lsepb+dhmssCK/V/kgFup32gcMn
s7C8TvbPe5SJW799SdJ0VqFevqSeK5muPbcMj7HZuAL71m3FHSBhnafNlWdz5pBqqziG5MjVXaGs
SuC6JaNytxuwxCwqx1F2PnY1Ewvq0ZH/dIEGn1TCMpPLCXY9ZzTkbKy5Se4Poi7XCos3AWdi2raX
I9hHftwnW9nvAiurrJU2/1xrhcYQx4DgJo+q4izRTei2oyULCuSjBWYrNkc+dyyfWEmlz2sdgTLV
c5MJlOrg8lVe7xK8eLBkblGWNMhMKCST1BHR3sYZeVI+vmyDzHkFyrL3OK7yywQd8Ga4mSZtiwRd
5RmMNH/4l8xVdmYny4La8K92fzlm+Bwb3G1s/09RxWHVijpDPhqwrTvMry5d8CqWOUkZUQrMCNAm
FQXFLqVxechcYxOpcjuFpXTaZjTgf6r7/W/pyM31cquES2JL5TGtSvAeOP0DN9gBIfVcDEbJhlBo
vlA46wUEk5qyK6xtY9JduuxQNY8OjZLEcWKiDq7cRURE3euLc+iNfa42UfOqPUKjGjEFGg7LtmrX
XIiZQDpzFPQVuWggxwV6c26n5yU1van5Do+kzcpC2Fqzr9eEINRrUIUIwzZcaADEZr7HgbKJd9cm
1c1Pp6tSU7yJ/mvVy2TW+sN3jylQiA6Gn/zSROlA9ysjMe/0LrORLV7Y819wmm/VgYsu8nbmxMUf
9bs1GxplrkNth92yRZP71VCFG10OGkSV2t9QnQU0qADv9qMEPGt+i2aF9ipTyAaPnezD4RmbgMcb
EEs9oepOr2ijk0yLNjAUBO62/PcnZj/GLVCvsmIWv9javZ2Jo2MCOHnPlAVjqRHRuFvK2Ncl2klC
8XKbR2H96nitIv5eBOdvAgAb2Ooga6F0XeUAs9bee7n8YTzCmhjS0tUXMheyxaOIu0d09ztTYe51
NxGMLLBUJkS3wLl+CLXoN7Jq4RMJLzzG8AsMR1VqRVo+JusdnYeUB+x9HacQW0DPqxIw++pMbQXq
uxERe7VtGXOxz90EwfsKUhH/ZuEoDBHhfsNhs0I9l5DRj5nkEdF2HR9oGQFfmZc87ic/WQJVMsOU
Gyktwj+AYbjszFCOGJ5D0vqeskaBeK6zHYN+7ZYHji+taoAotAUU535wNmzKhevxNVl0PE08BsmO
eWWLNlehNC7ceKOvP9W/v5db3uYBJC0BLqiw7AIKiM3hMc5vP14PdYgtIx+Y/aBie/LVeeUj9Ihv
0NRmX5e+GPiKHhHWsXXoaXTcTV7Kr7fyNbS0+3DVMSM2i6PweUGggJ6GZcqyLhMzNFR9YvaLqKxa
w1GxWjrnl+0F5US1x2KMUOxb9VrvqvKoLLBxfGbOwcPfWHQAO6Y3MxIBT7lWmUz3bOzc9zZTFtB8
WkOBPFORycHqRPfUHOqHyKBZ2UO8dMXz9SNCbAcapPEXMbov2ESO6kJdrbPYQ7Gl9JVYcXmm3G9f
ygkg9BK2pDsdASCGWt0mRXgc8SoCzQdT/wn3x+BC49JzkjStZttg/5SnpRlPj0v1FqZg+2KATsJB
yJKJaBWDUzDOm0h0dLs2KEN2YQZeer3zJzcq4CpdAWpHw/7hB7owSn90jc2dasdAgRoXlimjpav2
/kEvdfxJBo/lrOf8gtp1fYRfClRptVlP1YygniJk3LN0awGXo74XsOtrYsGVuWARscZezbf3L5U0
Wxkjxn5om7OXpoMU+8D5MCrFDfrULkqofgk/thyPxA+vPnOP7Xfhk8xk/3loXC5XSPfqsnCxBLyB
GC3ISpnVZfXvXDP53zLg5l8tUX0i0pLXxGQ7m/UOhmrwFuDhk4YMB66e1BgnqxFeROPJpx6/D01c
ObVuuDiWG8Zwm2wcR28YyzM00lCFeZkdaJu+IdN7HVKSZhrdtDgrwzoIYQUWh0+l98lz4xXpNw5L
ePE/UdpiRzLBZDBR4ps36V0t0OLr2qTprylrmhASsVbd7atJZwXoXHmLxmMKNjiuumZgxpsQvJ+M
SqkOIT7JFjauvP8lPOfaRQ6ZcAIfh36jdq+/Ni6E+s20uvmQSdyGcBMNkglBmm4F7eFMe6eHMBXf
s1ZYkouXAi+kfFlGU+aaaltIm4r7hWnHyt/nSKzKtdO8cF92qWL3o9jhjDHDHdo0mlpuvxI/5bvC
ASgnmGscQ5Ie2wrgaEt26lZp7QVJnZ18BJ1dRKtenNphPoLedNNiNm6R4yEsN6jZia7A58icbrGH
ubtJsG1UCeB65bVteMx6HEWkrZ32r1+i4BSp4pD6wjzZiit21+yOfOnQgxAEovyxR+juE6XMD814
wJ0SVwsZvepfDaesv3QPEmaCozeWf4CAlpt419UhHP/TQNkrrJy88TyAFy0f6HLnFG5ll0l+UDWF
s2IF6b/8MRaygrmR6vdp6G6twzJGndgEuLSXmsi2y+CWeYxrvFInhyhQ4Ih78IttcIFEr5izk1qj
wRrt/oC9j3w7vo9fTarcpcinsmTtfpeERGfQdoC4YLBX6H3OnujrGGIqMqTuPtdKlA773I4xdrDv
0GMXAgT+2qZ6osyLxMlw0wdfkRcwGA5R7e/OmrtXg0rqdpS7AHdIKF7hkpAXn0dAiVbDP+VDggNI
3Kx2ZUZr7bGSQJGgkAon7k8KFJOL9R7jwWKhLjStL7pg4wH7yJAondnS3qfVl5Gmq7rNvatD3i6B
UQzlj2NqpIP2T16njnu0B1AKrPoRwndMN7nx2H/fsR4W/rNO0Cp1IXLyswd7oed0CstM2zX5YpnU
6gKVsTdqpKsXkc3QIz9S3t+EKczIMRBYSRxK8JiREWP5d/qWiNJaZdsLttuEErDS2W0tCUD3ywhc
+0TdipBuhXvIZe66e3ZscMBFiyF8NhKv9J8FtAQ7yuuer//hEhhz3P1J8tKe9JyIdGnOutRqtBIM
9YslIN0Di/fXWfj9CNtgGYtA8egfkd67HCO8xIA0K+J5RsMw1J5XULI48vPZuJkqb6giS1Q/l7WN
vUH5FTK2yvL26hgl9D1a2cZHE+lybjXSkAD2lXA4SQabs7B68HzX/RSe6zK7LIluFW1BcD1gu1z2
xgc8xtm3LB8RgSaUNx/F4b3o+8UKQo2xR/uK1BNr0CnwogUbC+adtRM/NswhDRNRmboHekWIAff5
KurCOG3wJOIdnPfVZ5/2SCeyT/iMbIykFno9L66xWyI2OO/yYkRXP9wGsmYsODRXmAue/gyHS4wh
iqDfPcgPBX3t0fuJyTPA5Tl47NJ9RInzzSsG35ay+fCP064ELDNYvtjd2yNQVh1ArUNLKsOYjbai
CtPC9Hk8cl+WrEt3zeoeP+pM43wQTVvPh4Qk51zsg2tcZuMKM3BE3sLYHH/FFZt7zRaIadvehBbE
4n7SDJFgSWsMplslYgghr1KN72MfRfQEH0QLXMXUDOQnlunVGcLssFI1sZw1kESmET55UQzpj6qO
oiA8VPsHnYc1A5umpvi7ATILPfuMB7+MVmp7fu4XG+MRB0Z5lV4nSCl6dsOvCT/nr+Mgy9WJH3Jt
H0F7idPNMR1NyS+r7Zjm5Px/kI7VEZTKVxiqMDws6WDzWDFRlQxKC+hLsPYOdySyteUCXIh1vFP/
GbmXFDneu75uG11vKsmaui3IQKpi+HnmpQqrj5RddiP8MGQijw6v8Vk37CoE2ogrFke08ssSUAwM
p/BiUWtvMcDXtpOY81jUqSdrbZr/Uk9bLQlU7M9Vm7+5c2mtLHhURoIRW3Qlfe835prKY/xVPSyb
v9qKWqs/Z0eKM+C2rxFQy+pQlNqezUIGXR4kQCVjDCni2VAAPjFO7HmAXFUSmN0N3nq7yJE5eG2t
eD7fzFNXgwspGt6AkTb3fXm3u8oLVdH4PIuZ3R05P30KLr8wWB66hWb+gyu/iYua7DRRXFxljWev
NIOTfujnrphduBHcuPAFpja9p2xbwy8uW7+2/xRnSBjpiPT97CFCnCzwQYFvyGjgJSuqkr2YJ3zx
r6cn1pgWCEV+MycwrmTGO0eAozl2R3l6jnUjS4fZtQvcw9ADQlFHjtN32vGDlrv/irU9o+8QGb65
C4m9j0uryS2bu4QlWgAg7seDp0r70Zn6jOaEIfiXSOMjQ+6fM9qKqk9qadsfshWKCtQTqRCGsuOi
x2SnbQVFoDch4ANmj1qa5wC8M7yyJDgl7lobjODSorRCvXpygdNJe0r6BDvuB0wf4s8CIifX+pG1
0t4gLsIdOB/NtmijuQYBKoT1hXZy1kAsAPqYO6FdeAhDTz2CfxhjiCnK53GHYrTn3NlD0rgA5pzo
pBR/4KitaBGimF7tOk+CskLhP0iNmYfxsTns0NGFT1ixaIYbcYzt5skDo6xyF9DkdxVBxsVGCLPz
Dnl+RoQAIgTk8mz1a0LokydKuYCgPYnl4evr70ITcda2+pHpFDwTfsTIoAPooi+5SUHvgDRNwODE
uws/QZimZTIUTQt1XyGZo5so9Vam/u0IO1K7l0KT5r0ONROt61i78A3lFPHvH0L/devB4ZC4UOq3
t8Wi83wAIfpMMuJIz3gkl0ApOjygQFJaGXc174Yj2pbYLz+XIBUxorkEY7GRG+lZwXk5sk7X2JI7
DMLUypxqU4wXylGlyMhy3eQOMXCCSiBrxA9aUacunH+5r33ttV8c7EqFskACbBBOGkqldI71aXwW
PSwpLL5M93i/TjcNSM/mOV2rNuj2wldI7OpOaeHxxxdOpYlGPneJviGS2r0RVFr8gJZcBSjcwSwQ
bi+8S/vMQz6IJpg8Jelf6s5vNWeMNazptVw6utFP+ao7hkUCUONNb/Ei8Qo8crBsn1JkX108AqwJ
5AKs4ILqYs+9yGmmDjtNPkNK2I5aqPJbtG28RqMgqhbpcMbWDidGxJpvdxSFHubxVdVsOt6Wsrq5
zp4yigGYu6VlBO2Wu9+XlE99+ykKCmOBBoKo6AD6qJ3kjamhIEaPDBEfU3O11BS6l8o3ghvP4gnn
5btoDds+YSThwrqkdYNcbnTdmGuQgUVf76aDIX7hMuU6LlY3yY0V1wpo/I7dBbTbubVqaY+R8m10
Wp0gOii+ZEu5xsJizFk+4VmZrFHe26xCZzGUTm25qcQF/TAus89d/i4TVokrmp/kfK5Iao3zyvKO
FSfh/L4fB24Ct6pDvYx1jZYCuOccxasgHciNpkJFvWuE68Yfq30WrJxbFWtcwSk7XdkchZeEVYpY
OrcZbATibJyOP5qQ8PBy/W5kEMVZ5vm9WxdU5wAFaEb7PuUwqX0cBiGSiwHHGiUCKGkt6YikOyuC
GSHD/IHer4aou6VzkSNK+F18QgykyKqMauj0UWulPnap9RtoavbG11bkyox7fYymfrOmS55jKZhH
WiMsookAfC8CcpHtQcMQ11cAsmQafT/p6RIIw5uiNTsJLrR6oOpbgJrWjAUd5IskzTsBsz2M74bJ
nh4ELiFwSMEwO2ffbfsxb+DNoeaIjuu/NwKfMgIrokEEEOvc1vAUiiHZMvvRjqOmWHiI+0JcM+jk
AKa9BdIYvduWAVHrwPLtrGPVY8xAker5/tt3RrNUrVQs+hbxD4xUeQRHHKrirQYa4L9YTATYsbhZ
7zxgGDmzbyR48U5G9YqN0HPCqcBJUCrfcQldOrO6wRxUaqAyCw+gsEF7D+dZHiH4j0plfrCrzmH0
nbwQ70MHytGCDYBKwLiIRQrUm3j92nkdeSIe31Ibu5jutHcQvRubpvk71iaHPgbi0WEcIPfXui58
VSePdQlKmMwh9JDRYl6CIQT1SeJg5h2tLRjtBrAS+mlVdjpntFEgmZxfqjHPS2M0Bx82PqM0Rv0p
q1WxCLfv0/JD8IcTR9aJTLMQseQc3LANdND1M/qrtmZWgy2IngSg26dzKeD8lbxmrQhnQ6SnyI5w
RxznQVj71ry+TpMukCHVzaBYPVbk2jgs/QFX+CuR7nIkQkYr3rHHYf0KJ4B1GsYQLopVbC7/hB8A
zJfBrd9HkeyGmZ0YsvacdVD/8RtN0oD/KuPTvnQXapLEPQUf1OLvbFbxFb+TzwfEy8JBuSdb3S+5
yg1CqK6Z4vGUQVJWNU9H6CxAQ6tsGs6Gnt9A1CxRN1JudLBn/kXaaEwiKTVRsi4Nel4wrebUo1iR
IL4CBgMCqT3JKwkmBBAlmQVUiLFsM0nu14zQS7UlsmeWjr2YuW32AEg/9b49/iFcL3KKXfobR84w
TLj7pZUi1jJjrXyVidnSpz9mBqb5H8f0nkIQPLjFb2ZJWXW80xqz6in+u67OieM+J+5XCqJif9Hd
kht6hb5askBF0KKfx6uvar1caeTwhqLQQRYAAV2U3Eftmbyr4pUOHCiYZnkPzIw0+yZeOJUkQFuO
TUrGn6xjuB6DU5jnROfULr9htwTgNCihgrnsjdGzbzFcSiOouSyEJ/SqcWRgjjTWwSGTHx/3Yf4h
SUirdTwzntyuIKuIAsVvp+BpZ9HA1ads3Q+mzOmv3BJLDoR4fp0GTB3247Bll1KY414Hm+3UJk5u
FXUQP6gvqUFKbjlthSmPmAy+qfI8aYHV25E0VfByxwUVj5CmKjpuB3BGkQzMxse/E9ddhw3Y6nwm
g3FKtq5++Fx9lfMc2ZXbBDpmz0QsvyDfHlkHnr7wxl62D8dZAfqLFBoAnRDveXb7vXPd8mN9bMi2
pvAhuPv5fDeUHS+EcVh9cqJ/ue47wsDMmGzeRgScgr3cLgyCH3+ztEg328ZlcKN0FSfkOveT0NSa
pftUPU8Vgte7+OAY0ESUE2R6Gcn1Q/ulJFzfEmCJOkKU9jCI6P7wuiAxQ6nR6JtrjMce4LZamB46
Kg0tT2eUn/B70WtFBh0EF1ctlZytepagil+6BKnrarA0DIO9FVLIrj1XrcakbeCGMEF69Ji0Wfws
kHT5tE2e2WusLNADhW8+f++GdG2INjuFvZW8yWPGlbbab0EwrN4vvjnz2Z8jSQ0WhKSqbb6WB9Fj
G4PhD0sqkcHSghDHegIIvd6WoEnltqtzTYrsc48UPELWIjRh4yDy9eXrtNufKVReV2qj9FTK2DcC
Mud4ZKV7nDRB5ZCjaUQSAfO6a7YxTj1zBEiFNCd1HbiqpBGLmwDP97Fe8vOWyBU9KU7FfZYaABTS
2KIfOzNlj6JDDrupPXrDBOalKAwOp/3uR2BYESCa9IlHOE3uLu8EzI0iT90och5u5U5EOXX+79bS
24hPKnkQMBWbA3VLEJGkt3ODBETPl9CAf5m55As2V6LXIvT96jJnD9CQk9y3odjVkkSn4itW5v/t
ikDmuVEDmJAF/zmr1j6TrDTvbQCDNlEu9x6vgsOnh/XGer0+m/GmY60PZf1XlUSL8Po69M4ol4OX
Gr8k0zvVPEiEnNuW5HgsVbYTZuHhMz1iEZSqolDo7EUwlGXvYS3vpyHo3bQxb3/w8YPkM0Rq3HhL
kd67XhNoaO6I5WMPfaI5t3acMYHsLj+lIjQ5B2aXY11P0z4AOiAyiX1O01uNZGjBvM3KfJDwBRDU
XRMx25evc9fFKEmMTHRbPD8j11ntNFbxsaPIMI/d9HzMXWuaW4FN8tmqbCrdO3mkdQrCOZhNMcnV
KQSSmdv3R9hY5XTGcnZjHVyh8FeettOQx4rgdHyyK+yEoomx8/7Ah951nCz6yc6kml5c55aPFxUq
EBjlYyBsAwWgK3SFtt1VlK8b8mrgbacR4tcMMK3YMccEdMLQaf7k7ezWTzjPncFxR2xKtWLhTLL4
/UvoMxXCVMD99yUuAEElBNEWMaRl9wbPzts67zHI6ClH5l6NCSx1aolWtS4CA0K3EiKRMf4Ex+0I
kVShS0L+NOD2gsQnuZm2X1mDo9mHHbdccObaLeaiJ5zC6cPhCqNymx7BTCZzZw0ycCaDZdYrooIJ
DJmPv1T9muPeXvu+sbVna5VCF+sz/cN7/bDgFUWrJO1g5FkCDMtJoDbLob32LcIktTrpGNP4k1V0
cYBFkja3YqvveiZ+GNLO/gHZtEhIfKSqo+yxRC6vsoDpJwgRQSMvzDd7QwV5bCFrD+fvcu2jZ4DD
LY2AehFe6jP5noHzPPhOO+/fSoyYDOgTCgoNC3hIllMFKsuwXvaFs3YnwMryDW3RP9/O/fM90mw4
bVd49zh7kaAtZxfa5aUJ+dOzrS5Z9EfBj3k2zP9kbztGgU+BGscirrexQQvFH1hBIJ2FbTDmvk2r
3IEYtyoofxW50XyNWOlH7O7AgU+sAFHSsb55yYAJJx+i3feA0BG5fae54MVJfm5LxdUOCKYSPOUs
7tfgwpe/YRonXwZ1KLHP+51T8Yo+REktRzvXMQTUVo+HkWQeqzSaqaOYkOiMw51dKAwCVAXSaUBP
LtosGainyodzQN6FJh3cG113mk1eIsAtT1UeEEl3GICYHs7bMqKCRKgT7Cda4DhthF4SMMbsw/v4
b8uu6zbKm6C7Q27YsgrQZDdQlDwu1sHpPpREjEp8sRnc5bJhujrbemOysDTSvTdDGA1X/ouRFxih
wtgrZH1qbl2VOOi+VH+rMSEuPIPaqNRzCHkd2veGxUpJPRiHF/dCw+qlEj6Sgfq9JCyxTy55G1SX
KWRxiEpKVBW8ZAeEVgYoRMjY42MGa5+HJCWs+SKtOn0Q3adA7nThGog+TcQHZNtYTDDBCVNaSV6W
vt7kvw0Sowuw6Wb8JxOz2vDVkzxECZ0ihyPeNOGQ4k+wcd52gyA9FHgUr0uRGQ9h/+uP0whX+RBd
U7hqAD3fSk5yYx7Z57pHB9FcNTBygN9No7ut0l3Dq7LpDhxjnODyYRHSQKIg5uzew3qktIGREvJm
HEeKtUDDNBBbtHnnggMsFaSOvLp7+tVprXZW3VmKWFjtBS1lUDQ/GjyN7+86fmo5snkC3QvgiT0i
o9Qalrf4yROP4ujWql6ejPDxFTBfLfsLrwATfx11CKqyPyfm29tVkotaQbHi0539s3GdB772siZa
C+h+kYSRBRfVB7iVqt8pgYfjH3MdWHN3xlH1/sxCnadMkOUqt+jglUuvFcFAJItEXJF8Ds+2T+b8
ryJlJ2cIZPKXHXBFt8I3LgERlE1G9Bs8g8e5zOBXYvhd5Rf3bsA6fe7XC91G0nwICFqFwi8JwtMa
gc/jV3A2nMaIcNXODBiLv8HRHeVeTrMjkldxbS0oiCaadlOa+kdL1uWAVPwXaR66wc7a9w2gZgtA
qykHcpCzoj5wiL7+za2nYIvaZE8xCkq28SvyCh0IeQkuNewarrwkjL+vWJNEFemAOXeNvl1P2Eri
/FQ7TyIcr9S+OJJaVbB0sjNKzirODRAhNpZqkgkT49DPyp0AFiU/28sf/fMYhc+xHnt21egikxwn
eiGjCRNCb4bVlw+iPnLC1tIPRuYknFfhUCCc600t+mlFK75/SsYcK1q543isYguw+3kvEcKq/qrT
EmGVrdKnX3M5rDf8+TsiZnJ06CTAmE/8Y8zQSj/1+4nOtMgZRoftQWBQGmfNqZCPviDUc0AxfwqJ
81VnEnu/wdIfhy0qQnTUNUJMVz7MhjUGTPrEQxjruXv7wMCd/AE6Z0jMeE/c7kkRreLD4NPsWdmX
M9PESssI0zQ4V7ANnOBGFXQD8SE0dhA+ObFJ//pbgWo5ESQCKWU0oj+n4VrTegVfiu/ENW78C4zt
3vxrbsDPbAE3tB3laKy6WuFWEUr3WqH02XVVGadSnVfDO9v+ewYHFjEfQM/ypF8N9RtMtC0f7z4y
7ddH3gvpmhK+GQerDYv0JbcCy3my4G+m2pacHyazqRmKtIZgIV8MAkOwgI/CIVF/4iqWMywLDQXJ
XTZ8tHk4GwKrO1dZXAu/gHw/i0dNg597D5Xyitrloph1fp0U7pg0RXCiObNZlt+uyQGU6tcifkNB
Zi0JtXdyKXJ4mR2P37XG9Bbos/EchOuiAB83rxedDdwKli2re0fWi26TH9lVgLIYtjI7BBCxxEX3
yDv3CuVN7B0AXvRiVtOqx93Dc4D2nj9RGmToN4u9JPyDtXfQrV8llJrZPuwq511p4/dobc5q13yS
pDwQqSNcyI5GhU/z/NZvuQutt0f6v/gxrtKjg7jo85DsRzbC2wlPejLrG9n/UXaAbPxJuwT6l5+d
old926r6cddCjQ3msGimRCSB+2FJlcXp1MszAKbZplvmQDsm67czBC5S5MY1xRoGOGdptzpUaDz0
2Wa5CxkxCWS/oki4GPuMkz26jiaOSuM8kaTwHnhBgq8qt5UX1wL4AItzi73HbVe3X12IO/zVK+JP
JiVncWW+HvGqmdrbi37jjkUujsv1lHf4Rv5urFSj1DkTfbmNx9JXAKVIMl9vhFLbQ34fCkccg20G
hYbTCAcozVBPSwOwhD79Cee5aH3oBWds839p9ZlBluyQq89cmlW1I538liJQgAINL7QJzuMjoN91
PIzt8URctjfNVB8Js8boT1AHFxNqipp44Vr2F9nh8/gD1QW27wSZKz2P1KqnI00cD0lD6lDVd2rI
1APBFtb3KMwwMP6edH6dcGzVk6qNr4ckhmBmPMURd4AkPAVzZVjjOvvTJd16VTbQwJqH7nOVOw5K
dRzFvAzAOb+PlQ3tLRZ4oYr3Lb4q4CtVUfGm1v5nm5HxIMXFV5i7N0LzLt/Sghg4rraf/Mmc6UWl
+TugitBqJmP4kou36kDlZMWy53REMZmvipWjEsUy6RBdiudaSs4FIPvnB4ws5+Hxevg8ZDfXOd9U
3ov/tocs71Iyt0NawTrgddoPLgJFNuwcYDB4niDTQjvBIAU9T7Wey51vIZSZNqJ1/lFJb+YV+aBI
LilygHhqrQ5V5bzC1xATzygg7E1IbJxWskDiKsdyJ274M4t+1Io49cjbgQS/xd/G/iRBLSO2c6I5
sSdXzsTvrKa0rkXPbuEgLoAc8MjQa794jayDAVR26oDFRCGkNceqLMfR1jBTC8UuDaDbn8UQjRwC
neMZa5vW7NPxde1GkEFBIjmPajss3gIkpItxY93XF2W2Qy8uQUHA+lO5yhmENbrg29SuPyFSY67s
xd5fA94A9MUwVdJ1TyKhi1+C/eygg8+27M8ff/27ipifiVg3sf31xZdsZKzX6XwPrqDIBQnS/9pv
6Xgfa/CB7uG7aItYGOlhI4mgUGxwFpZiZUjmE3BBJl61al8/QGjt4bE/gEBp8/jckn9q9+0CkDxC
KWSh8ZInLC+q4/tP7qvTr3XBLyI/5PJFlQ9GsDXqIuDQKU6hYzNPv41+fApUBikoZys9Q26q0x2A
aaKktGNHZrfeAu1QOxSs6AKd4l1tmpxL2E0cIiXt3E3I2MfMT7X5zwYMmfH4bZ1Qrr85TnqNhD83
TyHBXqQpqclmxo9Kab5sz7DyHNzLgtUAc3xEBwZZzlPJosSDW2k8RObSP0d08nFFQ1gOz2d+Em5h
VikSXSeWd+GIvVfMUktkcYvbwK3FHJ4tSGdSkcBtCDmo9sYoFQ0uruCUqk8oHlazRA5zNu+H3Ykz
xKWuyw/EexgZbF9l5uAAGHr0V15JZKwUMPIgUWmqIBN8wtR9feJC8gMscGbFtnXDEyT4TgGhB1zz
9HHh5yd6GQ1uCQSTcZ2/28lIxj3JN3mZ3DtnsswG/FwyFxyE1erRVQxniQaP40d0IIVErdBkYs6j
qQ3BCdKuRoBfSjCDjx52kSJ0MKL+on23MbDcaveYEomXe50AXmZrexw1FON9PoVxzCR4BliOxTVN
6zwDIOpd4afaJ3ATPxmIWQFgCLqtHyiKnfxm3q0vTsNTw/HhQW6tfS4EH9EQGLrF3l6oJOSnLSQu
zHf1Z5JLmLKf8vkH6/r4wHgtUdVKmm+stw4vyKwN6OFfknHgcYj+wDNjcZpBFV2Pi6HUmq25qLtZ
FXyLsNHZ+9BgUaF3b/LK6hDR6ODXVlrmCbVcIBPiSnaH79Q8moCcsBLxIiITYgfX1MwzVvE4EDHy
E/1tCaOlPzsMXYAbpkVDcN8I0vv8VeITK79giIlbUaW2YU7ScuC/EuRmO7RV/NEPhQYFnhMyPZF/
q/CkVVcrFld/76v18QXkM5Q8Wb0fLfE0iO4V3KEiU7db2Gq6UGidc53KJjRo2tkfUqFzIKa2Vx0Z
kv+ASvK+RKzVsRWKGLo2i6ggGHoD5zkoKhQncwbV4zNqabHTlMGU1kDIvFtFAzIKTzrbZrabqrHF
qqn0y/YKkcuWdzlZTqPnvv3O3JPGih1g80oJdUD7b3pkECk3NKA5IQ5ftLhWnMXO+JhUTS0do0vn
Q6f6fZsaxd9w4whvLrtabVRbdAL3Wc+QANNTeFGO8F/CUzQJufuuj/tLnNuphhfSpepjWaxoMwum
8Q3SxbLCoNRn2hTtM8FlTV+vajJa5SAef8HHShfR2/HdDnoCX0ZcxaTPQ8zhJDK3xnJaxU82CDJX
udngAwQRh8LxjnEGu1iaNw/VFUf6M+Ph4ZcVG5PumJgd/Dve9yoP91N2QMXFRDGd9ARGGXgK5Rnd
Rb+PRJ6Vavk/0BXa5c2KvZxRbajcSYHdNAy2e5f1c7RslOslHZHFmORz8co6wPnWhsB5jlz80cAq
yxIOqa4/sRwLnwxDvNxWx87IG0aE4PblRELYSgcN7j3K0TywcCStu7yxVU1SZeX81JCnMa/+aCA0
afAirlaX9F2tVMeJTE74TvW8ej3Ipr2FQ2beKH+ibbB8hgsl4N8Zt9UN0s5YitG88/yaMhDbcbTJ
ZJWBaD4IlBRXcgRkh73qNPpQ9ADJsO3tuIrTpY4b3TfyjCqxzOb/33N/x34iRzvSBiCJO0+iGKyw
gyytK6xbGY+V428RMz8+XEHWruFosuP2MWlDeNuJr8qgZahWVXuoaMKWxF5F8FVMCQXfCnpqkic9
wexeBNrW+KwWlAwM5OU6u43zEYt3IAjidZmuYOFevzAt649VxqxuiCu1R2YDGKse5kBIIVgIZ++2
AZ5XBabK6N+sINDJFmSFQOl6HPgmRJwILv4CWdC1TVadTTQCrJvqh0gES+wHHZ9pmp0eO5mKAua3
11PeWxS76K5ebB4ceG746PYQdb/7EB23BMsLNjqc6cgyo8lELFDm0bJRsfI+amlvG3ZmJtT6cTrQ
qamcoBhGAJR2fOVWqCKLdpaCvS5bXDzPfiAAe4eXQ7QHVQIaJKir72Lq7djP2hs6CPNigrLvNNQa
s+Ou0pdKDSi/QJZsOrtBK1rHaLnAlep9oWTzQeOFuYzqkeKqBcHUjyAuY7gfJHP7QBayY0W5gZDQ
WDb/W87s8/s9v2IDJYL12HmXULqdJGK5ebMLTDAESbf2Pd5VAw2IsVOgx5k0EtYP8v46D+pdPooA
O4oypEu5UqMUlnD49CWjGGoCueGg0wVlZaxN7VszghgWjy5McTvyg2lJ/OIjCd+s3mO8QyqA/iPq
eG9oTopnUHoBR9BpztMb3EHsEcV5udU3fIzh+wKzKFU7TrHcjc0iPvHmjmlzucoxEu9IyftHEQr6
JkbNNg2okkXchFFVgymor8rVL/FtOo9GtH0kjGX+Iy8c4O3GrBKU6g5usjRIp1e+vp+YYdK0lAHj
TyfZCcsehzb/sVUDdEpFaqbJdE+wr7p8tgH/HLEfOu+bk3ozUxWjxtodkrni2IjeD9At9kGIkeUn
zN9kSQ1Igajuf922duSgLyawHtTzUnAszK2t8iunjHbFRIA5Jmx/2UEh3kSCRRhMFBWaR7pmu+0R
O4SWH3RfizDaXtC0249fRyhybTqZZ8qhvKsUI+1GrhHZsZbJzCUP8MXoJO2lIhkglKiggLKyBfYt
pwlGx93OnQRsQ5+cG4JxAvfySwr28r8v5bPo9q5OI0TmcOPZaIszQ4e+juLufuqzD7fp5ncspEoS
j5gUKcNnKGVbZWgOiVoxqOkBXZsR0/CFQFXkqUW5s0iFlWoYltxX4LL5/XhUW5/a1s/2v3mK0L5e
boNJ6rYvpbCRtR5Hq5y2sNejbhth5UQzwHTq/+EUW16SrkBMbtih4Og3Zu0CmLcWdo3+L+VKMRs0
66lBZ28rh9Wx4Po8sfrHloqzjb3fOGM9HnXSPu2V6DDL2+aaIFWpka697tPdqQQ06hBAyHtfYMV9
RSv/Ibj8pf77GGdt/jTF0rnkHCvZQvXefbA/YZbU9RaI78B/c3t9+OiYkPd0Yzup5EtHEpiQEEH6
E2v2gbCajELjNj02zeLXAmQ+ZW28ESHfogUQ9RpzYuB47Batpmuiwj/wica9QEbrAAZu57GjLwP7
R5sT7oSjDiVdmftsG3IwNtkQ+8EaUbOwKXLvgPFUxGj5XhxPq5f7VvmIXlriKBiDGn5bneQlOmRv
OiVPsKI7VRl3Y/u9x44J7lh551sVIvVWN9PRNLXQDClEx1sv4mAGAqCian/H1xwsMl9LuGFp95qD
Tk2vjcjbl1IdugiFlhby4p5FicxsXpdZ7HsKfxcnx5sL53pfj0rTMlf0RGB2Ik0VT1I43JkeYJv2
/9l25ZXdC0ENKMqiQLFEOB57EtjdNU8CyggbKhmiFcuxzIZ/hL4Gdva2iNDHlaZFkVBWXv3/fCmX
2msW7XCvgXHL1bXWA0OVBDBQ1cRKC8KLM+A5/t9hgBpu6uryCkwMknt4+dSFS2UKtkYSdO8JYUyr
9BdkyWfEXQ+EPe5UUH9JkmmNvc5n1qn/jwYloDKJOmEr1ASQsmtODPUyDmId5z+Zd7PuTH8wnLHC
giPB+hxQPTDEW3YZF0+pSROjhB+5v+zU50LQZ0HS78wk0cqZ/9FeIU7vukvn8D9zts15eVNGd/Ry
dqrj4GJscdec220EX0HHzteF2Qfv/rXuy5uzKK13VcrE2rnIFZPU7IzgrLI4SHeJtl3KtwdAPNXt
X4HVHAWqb6IpjNFlGBIkxF+udsz4ywKdqvgj5k/1j4gWnF8Fpu+QSTyimdqhmHQnvKpb/8cCbYt/
FY1nSAbDARUvdFxne3nGAUC719sF5dOCvOKKBZ2l53EfBETcTyK3lrE8UP8u87sMELDubSm59kaS
Q5Y3hMNwXBBHi4doHWHbieS8kmen7T2pAVquXpaAjB3QPDtRWF2S32UVimvVHTyj2cnuf5aCH14y
YvvpesZojmqyR40crKM/pH8QFXsZK5jOSIxjn6SthzyDubEUY5iQ+hy0JyU6OXgtLLQFYZPCwYt/
OOtIYP0oEhkAh3u2IQTAtd8ZQmufzZJfgsfEaraquyE7bRDXhdAy8lE3VUKSTFjXGKyfBy0lt8MX
0lQUx32iraPuJeJkES/9Ge70BEVqmw0llT9DVxEKLPM0jroOneS9n7v1cTEiEQ/ObAcjZ4Ar8BZg
1ogg6VMKVZp356MNDReb3IB5dnKk2p9LAOjiQ3R6YpGkZd2+GNAkNZkiGz6mCAvL/G2/QnRzyDrm
vEXonM6pqClREmOZIN6pb7XRFP1YkfJ9/hs/bcGYYG4mz0gA3qsK6lxBZSbSJj40J8vTdQAJK/PV
Zc2CRhwXvKtStSIwX+0phj+y9h2gsLa9WTz8TmYZbqYZLcoIf1KqjvhsKcUEy+vdlvOefKtOegP7
epObDDfR/d+5QOVYi2v5ZZHBYakg1AgsUxYA/s4kCsMabuyrF73VOp+xB4QH4v8vWxSbRgUnPQsW
YeuqUMQiNMSDVrakRNWAzGc4CANzl8HhdkFeKAM08CmhicQTA8d/uP47QJnS9L59b6XY8SxZWbFK
EG+dDLQM71bB/gwRbUSnFGxvicaTrFsqf2kIIb9l70zq6GietoRG+XGA218WIBa8X30gNEqp1+fK
X3Ig7Jd4XbZT/Dsk5AsErxO48IPZr97pUmoQl23F/wdnJF57CnBazsRXm4hiOwizeAd1AjQvjniJ
rQKykqsid64aaGUXUlJgXhumMgdvSL3MJFTxcfMxbPJuzUxBpyKkcWTntgmjRhmdS5myB+y5z0Sx
iWziZs1EZL1tg1xLeXWeKPhEBen9TroW9o+irXNJfi2GvdNqdGMjXlxOGTBfAqhdNyVqPUFm9GP5
hJRUvlWg26UQ6FuDyZPwS3WJCN1SHeymFibs6kDEfQVKuv9O16Otzz5u4+OVg/yX84nTvwrgWKRP
aP3o7gjAH4eV6K8qJJSjJN9xAXzam//J6i+ipGmpr0c+UUz8td+ZkEVxt/pdsPi7+Gr/KLYJ308k
aLzuFr69A/15Su6Yv0Jl/hA99AgTAmyvuTqp3FukZpqunEG5Pwp6lTWOaRrV9ziLED6Zrn0V87b5
Z2DzXJhIAdSOoFMnHgrDu23F1tNS6go6sb9BjU2JW18Em3ZM7JpsV6k3zus94yr9hqfi5dgiP5pc
d6SnVOW40jeIsPKmA/hB1m9FbYSqK/6oVXvCGQCQ1hQTzXdWTZcDzCPlsgL6X80G4vQzYH92Z7H7
ensHvlkbXjR1FQvwBQnd32NgrqPjSsC7mgpZfmqvelk+0KDbu0i4p/kgvdLisRnRAGalKU1BaATj
c4wg+Mi/+fACB0SZjkGLtMWYM60r4o9VTRpI9+WLjeT91FAEinbJbNY//rD4lSoN2/rqng7MziYK
zDDgvgycwTIA71qvDr/l1WcwuwKWnsBZ81vqjGKuHMBPVKvlnyW0jxvpB8iCVoWyMYgcojp7Ag5H
GOIrX58sueqcJo8QQADXevyuBfabbHseAF63btJDo5a6BM8M1gDkKzEgQJTYZUuudfu5ZNYIG1A+
N7wacjqVAzVhFY+lDF6nC+OVDqEIYShUuIyXiQuJuCowcaPwe0D7NgQ+4e9TmyHfPOzk9fKEhVU/
R/EfLVGCJSWRH4wswziq1tCak3Y6e1fxfI5HFiBTiigGLzJFihEB7vLNjCpJg1Cg+H2NmYAssxZW
EgfiUWTrmxMZ4D2lA3jxbksfTc/WJcn3dJPM42oKBYnqGv8TnbJN1OVIQcu2fvyWaoLbrg2ov6+w
40IQZFwEAeros9ky3kPwDMkxpW2EUlt3lha9EIsWSuXpf9RtglhznDzmYZbqtYQ5seozvhuPVqZR
y1gkES9qReYPTMR212VixdWzlT15uP7mtMKTztNqTo26aSSHPQG6diju2FWqv8UPtYz4nFnML7CP
B9Mqv93Nc/yelmN7GTWw3x0+hT2nWQoOG0+cloD/HMZnbUcYMnPw9XT4TqZKnTqiKzU/dn5fJoFZ
RL5IRmr662L0D00IX5i4eir44uYSdjV6A8gXLfEEKBGTzK0IsE1QT7qFr1Et3TRK+W6pvLoEYVwp
Bti7l/s9MN6iAGMz+WnSgngfi8f2k4NWfUDDpdlZU5Sm3MEq0wLGODQU6fQY2HBvd5L/BsN9CQ/E
482BYHEpCQG4ara2xRhZL1IXZgaS13ZWJ2F6VLZd+VVIz8os9ytSIn9CYLk7s2jC7a24t8hFZmrc
PAzMkh1g4kJ5F0jpL+5Q/+Ntezc0sRfTLvuvVCExTFr90p+fKrn0glbd5A9pkiD0EHGV44VojGq1
eOAzm0Ae2d8Blfr4FWwupoQRjt1xJsb14cFux+MI2yCTAzv0q/CctO+bZHdCCY0wN9jO0wSvDxD+
4VOATtqNllMbxOd/hPuC283rIe3avSwHLK0e6IP+TrQO9HePOVqvp8lwA/+vi1sX2uh5drM7XxJq
p7/Eej0UXgUHV3xDUyFOSr33/Ita0I+aBiYcp9L05pVud9HKghUCFN2jSC8efMtlm2ucN0q7EKf0
u9qEmK4zK8mGEgNQe/0am1VxbqVKaiVc4PIzv6DrM5NoCiBpQGrSh/KznP0zHOfi7yYrWAKmbf74
mIEe42a9l/p3BMOVNHG8lWwDPICfHEI+iGsogAhOpzxxu1KuBhw6+tbIzSNkh99/cpvv4mclLw8I
cShZfUxEm2oNKWSqRSC1840n6hVf2ArpD2D7NjhjBqWHnpwIokVEPevRkNJ45F+VwxmpR8+eMcOz
oWfc7wb3Pxo+xqxQj5HoWA3aa6w667JooSZJE5MkjpLQ+BHHs4BUxqRJ4hLnDLuZzO8TpIozKnxE
f0XVQBKJCTAAiyvASmdFKV43rgCWBk6kFdKpoi+N+8dakVVTTVXdZwUw+RDSxKj+z/ekZTrLijhM
h5ckFrhb2WAWVnJLXfLOwBWM9+4M9Vy9SD2E5hdwaKOPiqsm6ySlvQt5tWhYV/M4FvuCSaloir7n
g9ci9BC7RfGJeNPX4AQ9v93ukx8HD5MeJZtIiX9XJMj0xkY+Pp4haPke8F0RLyGUdg+bk5Cy9rWH
nHsYXcvyYEOywc9SFY0AOaqu9TJ+xqQrXGRfZ6ittm0ZIvJDGl09RyHbgMmwFZCsn2dm/hdMKDVw
pZ70+wbck8s4DChlwbMd5CQtHoc/7yuSPgl2JcF4dCK8eQHRbt1lvA86i7GBhWU3Nt5QNWpoccNU
yLm/x9oSMpaojOur//MTKf70UEbYRa7hHqKPj8Tq3uLz6pu9NOXZExexLd06pjlrhkCxoAqhoAZv
sUV2EzoYvYa5xQlvryMPImIQ5HhYNCUjLppByF8/LPlMHbGkrg8ZVWdWgeVlcanM9/uX4nj17mfo
dH3tJO26Ye1PDv1M6RW68WCgPbqLKY07x2Im6TudQmsPw8xzlRYXb2Omchscu8PQmJQFlQtsjP+d
oWD2okBFmjv3uL2VpdnMC3OBFTylICp0hk4tlSwMaceJRRWZYnmjQ45A56SzyuerxnaP08oKF1ot
U6DmxKyJ/hlNkrNac2iSrgxDGSW2l1Sc6TGYvSq0tR8wCnlZfIQWQbpL+qFIWoFJ0fLP6D7j80pr
RaOmISmcFJRe7PT9ip/40Xc3nzuBp+m5BR3L3GNa3+uXDRFbdwG8OUj9ZzNHZwxzoT2wWvO49vO2
q0oJpxfAmuQS3vh9NLEpV13vEcqDyb86kP8lJee/4FAjZeaQio89bWOf5L+Gou0CS9LpairWK+4P
R6//ophjtEckdoCai6axSltsI5LTAhlePmCMGYZhniZ4goCYqf2vxoqLVYcbKNvAnLSTQLAN6yOu
bll1h2BaKwRcscrYWjok88gTZOkrAfa+7Fb2QC5ya4FKEzpA5mnsGUzSSWynkadqRaFEyjbEwWmF
X99OCKLgrxX0mM55JRbvlORWQKycWLC4u1YxusoS29vqmGoSYySo1azXLeqvjYO7TUr1KCtmyvJW
/9r9V4WlQcGis2Vtgi6HI1Nmzy8HDL3Tdm6EdxPsocZhGtEYQuAAlmhFs8BVtK0Xdmca9DeT8d1i
GGE2QRyQCVFOeVl1Rq4TxQe+Za6tSmEPFMpXs9AW23G+IHZLauzxfOyJDO/z1IPvdXMpwMMwXFsM
0Jn4XnGRFM92+80zHtxGhdF6B4Q/E3jZk99Bm3BhMVZrWuDjDgSWfgLqwm0etUedaAbsPEe513pf
PtltahQ7JcDAcpRGsDT4laxtt4j2UaLIbZxEv873M4o+b0ZKi29mo8b0bSASH4RqI2oCakRZ12CL
6+AQOy5PUJCRlar/nkgXBJp/yev4RqMBFoZiOUqxnREVpIo7HMNypcfNJSsP7edu2lRt5ciUokan
UC8LVBThpVAFamzNFmgqsQ6WZuWF1yCtJz7pG5x4ez0A1sKyntYcd1adYTBQjBqjJrwLG9d94ygR
iQ0+wGpfE6abZcSnE62EIWa5fw1y9qBqQYd1HHAk3Tr4WGrLZ8r0nJUJ4G4zv2GZ0YLGVUzIihoc
It1aeusLsGLACUBlfI+kB8prC1aUIN2SFS4XYhRGOiflOKA/3C6FnAVzxSe3olGxsl4wYxliyFUR
VFhClZEPXgn3kLl+ZAqM0X+EHw+f/NMZwdEhChEIf7SnAxiJn+kVBQo45yj1we8fC2e0d9Yy8V+x
+ektef1vZ8G4XGWNAPMoQ1Q6ZIzBOYX9suO0atHROB42WbJ0Haz64wsTj8061/8cQgvyf8hdjHkg
4WUruWAPkb+IqioiHiK4lzO8FLG2dgk296hpHOrWkbSPs/S2YW19FE5EWcLrYXPB4W+mHU8zV+6P
w7NCdWcmwSz3IdFIvCDeOKXqpUyLKGGb2fd49LRJnXFQ6F0m6dxhFikdPfl9Mk301NOdSB5SeZPq
VtObNOhbPp7FckBoVAPN74bZp3MFOM2CI9mExsQ2W3yumjYN7k47luhxNju8mH3Pg1b1nwttVK5Y
cu6z3w3E6dZaV5Gd7zFHtSNNScuCmAHnQCPakg+2oUMFadMRLxVE3fwfWoxAtW5Fjo3jiRqPSXP2
xrM3b95r6S1GX0kCKzYjX77PRMcDjZIf83n03j3jeSem+xClMMRy+m6BHxIrwcC4wS1R9X16CeeW
Vq6MaT2yYMQI77zjkIwkik4QiKBpQQ1hqWg8ydEbo1QdSQNoboZQ7Yl+e3TVtBXLkZ2qthaDY6VA
aaFfAFEB9N9uzENj+j+gCAqwajrN3tf8c0PMrdkQnU2HQAhamQKisLDYCkjpIv18qnankjs4sOlE
DVckY81/0LxEGjbgQJuDJsgt6yAhWcvZB8KYIgO9EkSNQo+DmoRGT4qqFplB9S15Iom+uEsxLW2y
NYcKcpgRK8A5pdcvhmsbBXMsD1PrDlz9JkITjjoSXTHhpkwBH80+FCJnclAZWeeh4IRzJvPftzjS
030h1+xKeS3vcIO5p0P+3YQSekAmILqVtxctDK0jcLh5Bqb76tsFNbCuV/5zB1IVb6jnoEHK1JHv
NK8D7gDUDCP8j4qVQrDxqNDYDRpujGFw7xOPIs1+sokrD8dG57gGA6tgUBlLlRPUAIsXTA8NsnTo
NzUIPE4QvYWccTak/+JG5THkSXrS998NjPVZHzAQkG+63O3Zkr1OUuFL3Tbj8PV4FDChxNhgfB/e
cjliN9+H46jpum6dK37BqWOSQi1oD1D1oLd2d/kAZ7rRwxcT9Lk948CPl0MehX2e7Fr+ZzNPGlLa
vtJY7RCX9AonCqk6yiPKwJ6nybl5PgZAUjuL6ztxIHGB4AQmicHWowcdPXD0UUMqCA7dKSdCJaF7
Ooagd4D79P5ZsqGPMA+D5Yc8KFtlGPWGrhtLuowMnNDTLRMu6DkT0vzY3Vy8m/9J7AViy8OUluX/
X1XHR7qdfPGA0asd7rFfdmq1+DHDajHtubyUtV5nGXnMao0LutSd93YTFtQ9TyTUkyvE7DhJGAud
KrAxJB9b7TLldbVqjlBphS/2Wkqnus20irPhCjXAZxNpyQyMVSsAmt0Y0MWg1GIQOyt3GXeVbxp4
400hSqZ2WuMjYjernOcgp54WmiiTuOEv/+dEd+FNFBsb9v1jVefTvXRhi0PiYRpRXV0KNo7rfY+g
asqI2sDzGhgBoQVdP3YwLA3DcgSZAE65n6fJHxgimSItmomtS8nYeP8czQRFoE5FrnxOQaezCDe6
6rzJHWtEHB0vPxBl/c94UjJz9tGSgmsZN82ExaFEWZZY+xVj9rmbwVdwj0ht+RLLRx8I3El8rwSY
crbQh1YHz3La5noteUVSHcdg1Fooq54F72UCd6Gegr9TO0MCKdgMsO7MkevWSDItmLF73W2eNTpe
DVkbABBxE/0oPeAm4o1tS738ZduSBOt6nt9lJDNaLgzZRe8GYMGAEnCZkXL44mwPqpkbnSCiEWF5
TK1ymFzxSuNvIjqgnYNaLd8wh62x3nmd/9/5a7ixY0V3DGeZYLkEuuba3J+juY2RItlBMapuFk0H
9eZ1YLAVhQr/IzNI08FwTnZWX8fm2BJIU94+0sQe8jVbxgQjYNARRR/ICgihzXivUQI0mIi4kRml
/JT2Mg7RcsIh6uKdyPCTbEHWVfrGHCGE2mxG+oM64AYYuYDR7HorKsRvzmzW+4cXvepV1yl+K/Di
/VfEHkgP2ArGw81aNLzYWE6O1ip6i1895n7zs+dOR66biR43gibIOuNHqflxX4OHGojqw+ibumiy
jFlOI6m7dO8gNJrl8pl0bt086OCoi//PVEDrcgkkpFHPaWJ3yzEcAV3hR5Al5XW7x6Hj+vCAe3VW
9ntwt4NSLMGdc2mJGg4d0nfozKeTR7qPmI2id9JRiH1jwYqkDZRezbJgW+JYaCScz48lpM5v2MnX
9gp+4n/+0AyGU6pS1AV4jhdOUjpDFfKy2vfTQqGkHpgBB71Zv/isf8Ys7UedPYSdGXlxZwr92cMe
oMVXEjfegrtoU3ydfIMSc67IrlmU5ydUk7E9WKUi67MSfAEJPX60Hf81HS7PqfhiJ70uCOuJarrt
lrTYA2cLD5N/DGXSyZU3kodP6mAVVNxDgOAQg6Ffb21a1H3vH3Mbbl7E6qSON+G3K/MmtCCf/zAZ
b1uFcLugJgurFDFDMDtVCI6C6tpsvHdcWikT5nyoKtr3xgYqPUbHbJbDd/Ll3i1maKqkqM+o4YKN
pqboZ0H/Z+JhPle8kMbAqBbZTmpORV4IOqxkXU1fvRAJSoOkeq4jjryOmWsyDTgPJ399r/A2tuop
l1KwO67n7qKl+5XdwMcPZf4oiMfY4tvhNWAxF4l1/Qlyf0Y/ZXJw4fS3aIBExU4mgVvymrioe4mw
Muwn684ytu1pyCDWCtjqH+Zsfvbn7I38/JUQ6VdTNdu73wNpsIYETEK/76JlAYlfwdc/rR4+i/Nv
zP5Onp05HJ3/nQZqTve105KQ1hdnnfybfyCQJFlOMbBXj8/6ypXyazoaY9ImcmNr8wvbbFwFX+6o
FwomUZ6YUhTE2Z481Mqm/aHjKG/DSJdmwic8FLAExIuFE280GoM4/4euqna0jUP39mmf1vTpt+GT
Wunb2SEE6vv4R5zJ683RL9HMROYKe/r9qsy6h/13ROES/VWlc7BwXruqaWc6ijINcwGicjnHOwMh
KLBR1lH/ve3S6id9fKbb9IhhRXACVTRklrm9EcLv9E/0XwQZlbNSzlSlvrl6dP7w9yCLaSTr1UVb
M/T/4zJ5XRIKs2lP7mU5pcoGr5AP3WK/ezIy3BjrS+SP+2b03efV72dcv1kkzXDziFaHfwhE6tlM
OR4ZAZe2lP36of6R9JnAYsuRoWvwU2sorYIipWE26lqyBe4/ycShtxke3AKbXgbWJElEieCCJezl
QlbtacZnjg54OlmCxhOVfYdKrtaGOsvqYIz43QaYVlDxk2Os0eFOMqJdsw14mL31E/cJuVCkqkMZ
gD2Zy8ENCPY6ViI+BF4PThXzzV6dzKiXwTbxg5neHkvW4u+DgDxQgHinsIPnYskTTcovAxWol2qh
BHmv1wUuX20ldOho9Ng5aM5BwhK/oO65jBv7o83LWAL65R6agSDm77g36mv79lKQcqloPXUdUlfU
CRySYm8dc8Y9hbsqBDgOCaLjbYdb2fnoAsgkTgz6C5/ZjNX6QM70It3Dn8bo9IRIpPxGNJk8m8Ov
pguH8VOjtvtZcFlNEvr+linesyE0E8xp8Dp8skI3jWsktwWIZ/RyCeVJsVLOHidrFAXHrK9RpD59
lp7XVFFvA9Sh2FCcg8SrIFAdU9++HvibYA85yGykwG0wvakryuonsKCioeAEpuBb+mRH3gEfgDoc
a9Es+fv/rbLeutpBhVhJoxKlgboiyzGnWhf9bN3Ti5dSHznC24HRZ8AzL0S6XQ/p2Ie9ButVAE9T
38YwQ78ll1zmmQvU/q5IcWmatdCvbLkqFzPozPlUfaubGZFRGD2goTOdbcqIeoT58F7FRXbPJ6gE
Gvs6VjRw5au74eLytvIAS5jF5B6AmTWW2VqT4wjbnujayJDcnGJ/Kt4UN1EezWCsBbANC+0noW+d
JyrDmx2mOZpZFre5qxIutAoQq61mMdMrmWhOl550MY8XkIEe+P8lQTTq2kpuOWFCdeaEAlnOUpVX
ClVfsiT7DSX6NwiFIn3ZspzIp3nQVFaNDcE/RWFEbGwxbUJQylDTASAgurL694wT+6cPjO8DRH66
JbKyPrakyf9qzWeTqL5Tm4wRqCtBqlfnj+KMIVw75e9qrRnM6gmtMxc2hAzdpJiwfcfq9fGUEM/A
A/ZmLiq4A++Hpg7KTdecTGRb+L37djNsCvHcLwVEvZnqAvGjK1wGlUgb/LyW8Ykpsj7iIEJQZXQM
1XC3bgaltoGM7dVO1jlMGyD5o6DFECrIXKVmE04CU4911vz7o7VhOeRmpxpusXOQfNluzkdkLW/Z
YNyyFBehzw/o9wZx4IS/7AfpOzXFbgT0fYo3PnIa4KdQLGhErP18S02PDhm8WphNwDtDWPIn9XDQ
SjIgiABlO/meBTrko98qFr0X7cdH4yE1cHXyKCDHTD1F//1xmlgTRhWaNJ/Pu196RwTRxEoTiGQt
V4v1Ba0v32hTl6lNI0WmiRNk/7cN9i7F2HGgP0F4carQU7ZGdgvSoSsZI8CyLfumMW66fUtdJuAM
hu0p09amDeav6siqt72NvxHA/0rD2/6zXSR8prWqD+kyYsUmng7kDBWSLjbp0WeOULo0K1kMlYiW
Tc/orbe7cL0abQyq0FBlWUWX5pCx6tTJs1Acu66seBhn1Q1FUV4wOJsTlOK0bFtKGrSajR9aAnVJ
YIvaJ7iSGG0+MZhQuLcpa8S3a6ZK2wrSKMqI6vUu95XERXxeVGCTiMuj5YEQaCCNkZuURxRBG3xU
EcGRq3/lsyTx/i6/M9YJkVUfstwnSODlSlPpzXcarXx8hBlKuOwHFtXy0SUTPNMP1dExB9AVKW+y
3bVE0gui0wVyvmQf8vW66cq9g26+50s6l4YQFt7UzEfdM79AUuiDrYyWkTiGbffquHG8DWN3omPC
Gqrr6yXLUkYhs44TxCrweWLpYxDxhRcJavTqlhLyAhngL2+R2jmZPcHWlbDjP0nMAR574h0hMfDp
0sjZ67ZsYz9PurkqkCSD86I9/r8MmQKLdxnj7nLfZVmEXJH8nitPa/zx4nMXdukO/IZdLp9gmiqY
btXxGvoKw+nMBOrG7+gt3VxewFyCQ/D+odI4NTlv8zJAtref7IaegkyqY7zuBOygVInvdeEnbsxZ
GvRrWkdPXSTM0dHqwpttscRD6QygVOdWFnGqmnlnOqO9k3YqV0okBamXNzkJgDol4jX7K3amSKhK
BeZlJC6hmEwVn0KOEMK18n9NIUpbbRC8VOuikMBFki0Ny5ZtWAUSzBERm4JojwqgrXcJq9hEaYzy
VVqjA4zOijmsmUFJqPVJm9EqlsmzBNGsqS5vJTlcaYwdt3TSiEIYTlCw8p690nDGngsgfwCOgIzn
H8nUvLACVCpAPVykV/WsbxbXFckvvD9cn3xBkb104FXwBdXn2iAhehwJoI0Dg4RfRgW4Mo0e11F9
4Qrs7C4L4pdkRpUcPgW5/+vRtTlwL/hfUnjTUzk2pXNrJMMj5n+n+mZpYyBCeFHD+/0OfTFiC1wX
8tV5dPSEoaPmG/d0Z1pSKHYL5oLawvK3wntVaQNdrwQujfhkh7DD5B5wyOrO8vcpHtvbMtz8a72G
Y2CMqNkx5YnNyvESzfoRTHA9Db7QfscAfwW8X+EbFZnpWWKc8HGB/jsfvNIz8E6regO3zaiLwozI
CVn54WChFsDM/+BS6t94PIAkPEFxWAUu8ybtUUMO8DZ1Xb6qjk1bMAF4ZGISbK47XeluGguJxahO
KetbHv8bo1hdGkJDTaUFmLLw8/UuCciwUH4gwed9sEOpeHR2UEGrzYhgSjIcS/iT9H1Q99cHIR85
b162/M41YWMnY3Qf4+9hlOTBHCgBuAue4MhV9SEiPeCdZ4zQa5ImpqDjulqW9ouDP39dU5j64uYn
UeQByY9AsD9tBtMbo4bpPRv7MG03EChWJlEmoHV7Y9QJs2CeMNqbdmgTI2E8QWvb9pOIbiEbWt8K
6bFs1+Dd4S297+tNukLitM+Kn1NwoXxjKD85clp8eVQFn/NKAshMH1vxsaqws5VjjzCq4X00Ltfd
MW1zntJQt5uG2xVC5vNMNftDCIG65V1W+vRi3uaBFYMget3MrA5rGhEr/zDpj5Q0m0KItV1tPk4j
VLX8nNw3HHUnQADJ4K/SzdkXG8mCapjoCmMBVzZQ9fft5uWQ6ER38x9cQZOR1qi4Z8HCNSXdqCWP
VYEEcSmCCdcV+Fn0n1QygIdn3ps00+QI5at2Ijdz9xJ+GKt8OtkqaIyOfDphE67uCzMY0GXSSVDa
MFByfTT7D1o6MGmjtNezCy8cIPLvr3fSRBzlKLb/NDKiSrDL4VKK5J/wr4Gddke5Xd+IqFjU0WKv
PYff/8uDCTYh47BgTa9gZvdkRoOH59pE5+yhkMUmA0p80dJGhz/1YdPGbpYtJKBW3R0BDYRXRJgb
Zu8sF+S/EXcozgGdR8X4x/rbI8gRmRzoVu6yWEZyeAC4s46nF6MjoDebABxcVnZT/zvs4OPG0u8P
OJNrqo5FB7xqWsNJeRk2Xh947Ltc6710/S/2qagYG8mcIDyZ9jAQYhKeyzmM3XJSInXxZOT2bY2y
55FHIm3lHuW+m62zkdJ+jbBFMDGmgq6eFQXMEnwojL/ZypViasu+Nh6vfAB7KU+898PthbdR7FFN
SUnLlWxlYE0bCno1lqkLGX1tc+QGUMF6W8RO5Quu6biQtprwI9aX4uc9BXxw4TraGDaGKbW06nWc
mm8xZZVoPbnwknv8mP+wqfCDtjvjOv9VctvWPQkPyJ5wvSUy3SPGG6k/Wh7JvXn7JKuNtAQAb0kx
2oCOIdAPQJq2EBPRlPELo7x2zIQ5MkXZI6v8Ra8CGq981dCrZ1VV2pt54uDF6ZhKN8rKmDQ//BWq
ro7bLfZKya7tGJ1vD1RVp7J2V5/XfG6NIEDA4BGIk0wxHVpXMLgybJKXv+LNh4CoT6NhreNB/9hn
pxmhYJ8xVhe2ceIIAMzGoyEhWSHhUCZTFif1LAPy7YvuU/YeKxz80e5vpTQTXKCvglok95DPqC/u
RZG9BOqRvSxvD4eBb9HW4vCLpzd4ueaf3atP/UTWCAeauhph9Xr0/5w+DaZRBmwkoYgjpfHqdaAS
WG2f2hbtVT1OUkhaOo75oaZ9S8++W+NEL+Xuz1G9gtxzKhbsKP6DNci8JhakG4yCfrbyRzg4ZlGI
XADEQ/HW7NrmI9BaAzZ8kyqaBAbtmYrF4V9iE5nMqBTQqh17HM7UuMjbcV5xjQ91GAKHFCLQApX7
ZXJyF1UmJeJ1g2pqJBe1dOzN97P06HC29Pi9Sb1ubrqACNWR6s5o3JImaWL/sHDCdi8SSb+83Nid
sQyHty8S7e7FsiPZDUNW28hrgzpgNsny/DymUlRmiyz4RUmh0pDcjvn3b83pu3fz97AUZmiDQHUV
j/D+mjvMK02YJiR26/hRoawtSfzvMc56eYNkby9k1V1mfLIfOwOJOBzYpq4IwxamEOno4XEr3PrS
uoWD1iYLPULZ360C22f6QKvSsHHIX1jprbZAA+fKibUu7SB9qsWrpXhLPYjZuXJ7QcTFZfDwk5+w
NhM959fIv9epIBYxUEqlzRtx7CEBtLet/5FQ18OkoAzQDh/JGAojxI6rp/TZeASsVSThwcT5OBhK
sHJRFjLlO3AjWWvIi64jtm1/BReDWus9MXa4wIGMYH0mDV+UZ68MZHDgXbBt3w2HpdBi2/gJsVmE
k6JDrvGCMBtxEjCn261UcojbbUGXYwA4TTOe18trxXOCMn8y68GPwuzRywociNCbtZoLKc5OmBLa
HdwGRZYkNQ9jGneivAK8P3rxvy8tQLEmMNU3igFgSaCALxdWofy0AwJZbfK103jEqHgaC3GONkMO
87FMiLRfwRlbmoUFx6s/0xy7nqEUdxHJicpqnptRBxS3FVWokYtptSpmMyzj4AvK8RayT22LYxau
vj0tUKFiZ79A85KFGeu+k7fxIOhXy2vP09TUS5bMqXhEWoogxJt+anfnGNp1cwaAFlgBYHXH4YPM
CDgNmNEM0Z1oEm92nNy+mrB4ldrdcPMw5hINlhDDBFz/HJw4i3wW9Alxg7MRf5hIEcZgYmyxOkKb
cntMsJ2QURcsBF85NMRPi6+1shfqO7EcPgNiUj7YFMvjS4YfnEne0L9mlrjOC0JSePOJMZZbYd0G
m6fuurc7bEJ/y5T7z7gRzH14Guyg5AsaggWQCupLtg27C/FyuSHc5HEvuRf6MMM85mtUGPg1bYQf
MRypfdfZwbsLomjujvJcr3IjJF3Po9tZF++aq+qnbFkMffTQwOayl/j2zYH/H/NelMV15a5XvGI9
Oy96dRLBS9p+2Sxz3uiznMY8VTukT2OzcQ0JG2vpwL6BdcMB4VJopGOo1NVN9h8S7ckMw/mDd+xS
wpPFRIgoMJua/lLvxg14z5XwXLlNln4ymTvxMEs3M47WPLEH0GxsRBSgzj7Xx06+L08rflcvUcBy
4UZ+nXyTdUKHgWuVTgcRUBtE2q+Bwq3dAfFrn5ejB5JXX3FRlhubaUu03kbpRtuzdP/NKHmbwwlr
PIZHVTEPncu2iqClvVUhfjIArRW1ErbiE/6Qd3HBxuFxQyK1CPHJy93cLbiXiVZJ6RhzAKiyZioI
cyu6qQ24l9gf/98Sm9vGYNHvwNDRuQQ5pqE0RoMZeeZ00rE33PQG3p358g5n89eLgwiolzNiGNo7
InXGlX8AnP0lVPIX/GB41A1jSIJ6U//5RGfYLydxqKoAnx6UlKIeohvL2Is9osJ9FHQLAlhAZ8IE
0DWrswsZ6Q1KBjVAOdy+24awozLxR3UBUtHFeUkSREBPfVVVBbnmnv4xLGEXZ6BHK12enyXV8Tvi
Bq2z+szvgWd7pkJ5dz1Dlx0JnZnVdv6NG0WzMYkleadEodQZppTbYTB8KdklZu7nVzZrCJjc7Yk3
/PyDUbUP4NPu28RIXxAxbw2B5ifgAkMnToN8Gt8aqZvejFC5fJP/Ym7mVOsi2J2/S0l0VHyWhI/n
Wn0/9tsuRqWg4vdXs4LTmixRbEIFI6nB2QOEQnPrCZ9a86rVUZk02lCeaoUsyAvqm/jOAF6y4mU0
a3MXMgfGvAUvaUnKsoA+KKzUxSj6bqtLWVs0T2QSyrxHt4AW9FUX5Dqq7H4bHL5kOWbLkRrae8kY
stIj9ys9LB1c0l7HRi2728CgLK1+aImaUPWzGDWBzUn0HCCRLV9C9KIseQPT2Qg4QTD8qRiykIx/
R757YXUBW/k/LrfV21LkpAY0vYemiJJkjGUtr9YHB3g2Y7J6i/jbZdC/3EuwEEEP3xBI7Vsd0La/
CyIolYXW4gHKksqJIB2RVjw47wHs+LocGzoCJYEq34I2Hz6ukTgLpBeqSEcydEUS6M7s4uNJroVL
1U9WicdLWGXpSr+UnKwPtKx+yFm6w/AGtCSLh28dTZpiFyQNAPH7ccgsF2LQtYtfzlKzipo/RqCc
ihoP4Vg8lgJ9VavoODjktD7WFvs+7YwvHGnH7SpPZMseKRuAvXaXRanpFVJ7H86wB0emT561zF5T
d0LdGB0oGat1530YXZk9Ps2KRtqa+vItHTE3+nxrI6k9+XiudFSyXJIsj/OLPMPzZdu+RqMjUU+X
EilUQgd8ZAsvl9bXpfer60giljiYRGoipNIDTIi24fFkdXwXEhT29OLfTF31AXp9b7RgMZtfTcz0
l+wEluL9nD7qWWT2/JyeOHF/FQ431ReUt0KUdH3vVHYZ5SBnxpREAgu8j599n0PprqY8dY2GW80q
2rK9Pgbpi7CNNE5yBJZU9CSOX5qV7deGgFd15fb0hOWE51giz6mxkILMonR4Uv++/IPAA1YT14ey
uBacI5zScuZd4hlE5oTbIEbdSLEydauiozk2IrmZeOkuWJX311uNVJsOtSUlj1pCQx51kInu9jZ4
04Zw7cGE3xU9MH1kBTYJ0ogPPCuJS+nJfQpVTHGoyG3VKt/WMfe4NM5n8OG063O3JqOvbJoYS8lg
zgn1ZU4T3LKKWIeRbRifBp6mzZW/3RQXhVQUu+pVeoFGhT9zRwk7dAVYdndPJ4r/pW1berBGcJJc
EZ8x9jrJDtz/gr0kM26ms3Lxe2jRX3KYaS0biEnjloaarwYYHPpy/lquBt2MLteVQ8GpCFhtEnoK
Ca0txryB2zoSNqGSgyzEYHQ8Lw3yUxAPNjfy5/MxEZgQTZ7N0jq/XYtJDvkp6cl867ct9i3CogiV
5jsvAobo75QJnZDfuHpgv7i04VqBXf1nn/l2wKxtWW9aeocGdgFQNF+1M/ynW27EqZENRZpaDpm6
rzwRDz16QT6OEeU+cfg+SQORLvsxwTUkVaDDpjaOICybe/UqGEIabla/N36hC+aU414dMZ1vWM36
OGdK4TeIA3x7T+Qd666jY6FyhP2xkXvJ4wiw1UwIfqVf8IrZQVHXEXpTbzHQQzhIBC0Ox6ljgSRm
9ltxI4bNfT2WgiT3Mhwfp+f8Zo0Zd9sl0eyCkiMMNZuJGOqqT93da7SKpiv56W5m+biPek3DNegv
Kd5givn5AmN+akl1ib7ZC9jrcKFuH/WEgL2dP7r9G+fZXBKGWVSNqfFzZ8qzwDB37SKXuveahSP2
gdeBy/livUWgG+F6R3viIhu2mIzQJiTkiw1n4qHApymxUQNInOAX9Zi78QUXZ3OkL5MfaTOfIqMa
BQMA2IE95QU3xuenZShTS6UxbmOJnHzMJTfaMz7KWaBqteVYAhgEXG3oJ3J92Pxew0/MB1mAS7Y2
TRbwShbvMeUdssjpDeKqIadbF2Qsv2zp11uiFzNzeHAyvHJYHR3Y8PeSFD4qru0FRACneqGmz4NQ
dXfOvfe96Fy0if2aOHwuPZdPzGQGBXP/weB2CC4dSO8JvmuvG+DmjVsGRL2Bntj8/mkTbZITcSaF
lCViBeO7JKtwSqhPOyBDFVPYXpqNP6LctwHMXZwYfvehI1lLt8Xb6XuCTUBS0I3QjUBPgzdp6sWW
8UfoAX1EIZalcpzlbPnTMeuA0NNFx3UVGJJdYC5vRk65ZnE5ATQ+B5VsRaSQ4/+X0KVx6HjpVghL
aaEqpAfYDt3d5w84oog5F3vhgBv0SH8SFkdQuhqNmiEtUaSPMw6J4mC0Wan5HfRfBSG5Jgx0KgG8
gpHduLd15JkXKZEuwrupxgDXOXYcvfx0FHK0eH3u/Phf/MhMg6ccPlJblYsHrbG+QADH55Tzjqh8
B/cff3svPoSaA92dGcmjIbePro/4/gzePvnWUmXZZlkJFTwgkYjcMm2xJKjdRNBPrBskj2wK9RDc
f6KQsd2Xak7Hl1Bx4r1pG+dXLkZMCZ+6qIDoYjAHIejbkrRWU2RXVi5gogB2++jXsPAPBnGAPThR
Bv7AwyuNJwM7Dw2heBsta6PszJ4fllCkRs/JM/Th9YLvPxtMYIoBxdTur6UfT4mJfAIwxMswyinW
QQYUAQmh00VC11uGqtcd3YtjWuEo9jdRuiOmLPMlsGnUUetQfWSEewLVJMCVarFeHiVAKSaMpsRC
J5IV2SF2n9EDRmhVXyYrJaQDHNEiUpwfJw2dJD7gDcre1o2I+Mf/BIx1Z3VO79LDs0Zpy+vx4r1P
J/50J8S6RdoHK343xyBgi0HhBkyjpqasKPnK2KYybAvKhKMvqko0sZy2LWVLeA/Xdr9gmfp+fwxr
3eUN0T5r/aKRrVOCEBBbGVma2yO6GDPqi/KoCN7KgTuaJYH9Fatw5VZDQx8rQfxOkvAfeGHbJQt6
g7jT941takm1zGpzTD0Sil24TpuojpLGh2UGfglDYV9ZHoQJHvBVayhzEeSl1V94+I39nFk7GtRX
9EJqrK2ioOi4cb1StKJFfwRryLUp1sDa+ehh3m5CI4ohMuwlcgjGVKsxPmz5Z9iCiGtjkPtE96vA
G86RtGIlvjPjiuTlarGGJJNG60QNuyDhHm2n/DGtlXIx2NhTBOWzVzWZFHhqqeZ7kcz4e/2tc6id
g/2bkHG9IP4ILqUPOZfiog6qWhxb62vh9tfokITY3cP7QKcbUawylzs3cvOmqeBAh5bFYPLu6Pjt
QaSEoxtLp+EbKK6SnFn7sPDuG8R7IBa3A6MVgBQOP4yTWGwGAKMjzvvnwLuvwWHFht1WrxF4WEEL
BEhPOQeQlgoIE/0mBlpYqC6Dssez3e5H38ZLL5LNDBZH3V/hiIv+Y0uWlZ+qW4nMDsCu5V7tVKUm
Bf7EamZL3kHI+H4+D7ZfhIGreoneLg17TDGtLmTPAMhBFl/JW1tG7/nA8j3qandqpBa/ZYQGLWLm
eR45qYHSwLoP/QTaknCCHSRx+5NoXAA7HeGZouVpDSU9Cci/XzHNBc2F2faBJOyIDNRDOcFXOqyi
s+HFOG6LseBb7YSCIBkr3qlW3Jk2YuvHsrY1vZ4p5+xwx+Bh3QaIuSfiq2HjzC+M6TqYG8G2+ATr
yPVOrnM4dZum1sL1hSzN340ibGSKz6/soQyQreNiYEm5GCb1nuFkb9XIbNWiX6vhthvPBclbnYD6
tcWFgduvLJ8DAHD0otVd+xIG1P0CxUteB0OV7xfo5+a5LTOsIgNl4Zlc8LiaXZhivFo8PJCjjKrE
TxBBFTB0lLIhDj3pWdAix6R0XWh2gitfM9Z312+Vfag9XwHBiyuT7CmrKeiSatyBSc+2t6NCP3vw
ZWdvvHRhxHx6R+sPEtOwutTKAaQhIdeON1VAQ3nGW55Y5aGj9lBMT2bS6f+tbvvNwSo9xK/lkLJK
1YMceKMFKJd8I0+7EanAj5mgOfuNpAwLSEhWIyRA52GOv5mE7mu3OF9kEEoY+AcJXUT6+OwwBeHN
k0FH2oovdu8Q72T1q6rPYvt6WLxDW46xOaa4meayl1urqRwlYBgb+d36lWEmRKJL1gmOd3fC+Vng
fWKxJgKUjtAyS7eCHF5Mt8/jXjBshFYmgfo+IK64MQUUfXnLkolShutBMD9YTbQ0/Fpurfw52Ath
2bfPtIlmU4JDOz3nybWoNbFocMUmRmNaG/weYwbPE1Ci63+xLStaHB21mk8VDWS03AXtvJnYOm71
aC4Op4rQZ/2zXH9weXEQ2Iu8VTGWLcAgu3wzcQQkRHujW8ChKbBDKGNS6yMIcbcl5b4lBJIKyvrc
m/jtFe84LpoccnX4zrAtcnHii3FzMFXAzhHJxQGkkblsK8s1AVKi3j5Ove73Y6Bj8+J/RpPlULvE
yeNvWhNiJxSLxYwAzeVwsIjdEZV9ohRESqo61l9dc4bJOBwGeCiG1eULVsSg2Ho55Dhn4PO3iZAA
L04nRLOk5aFkuR8QnHJoprd3TTPopSmT8VrsQNrtFQujSvqcMfYsSuR1mYbF5D5sP4ZgREst8F4g
KyTsOIZLURAjWVbPn6gfVQ7epE8XDbKfYEeKtf61LsnW1HypdJ49OywOE0PNSn10yrBH7le81KCY
nBRY42esrHGP9hDUg1JP0f3gY1kG109PLJpShAOIqI9o7gy3AppLD7QlW/fOKcx0ERih9oc8KS8t
SMPkBGeqX1y0zlBLi4ngYaown6TjlHB+TR7cnIoFsLrbI1+6796QhVm5R9maCth+3Yv3ztxKsSRn
lavOrlDRLwNrvIzPnvTH3XnA0lPcKPP5OnJIK4VpW2QYtooA2+algH73iriC8PgLiOmfOQUevnrg
HT9NTR+czgG0KZ53sf0/ZA9vTKgK3EBvzjKI5xC0E1CpNw4Sr20Qx5cPKMzlqetatvB03fhFtOim
WaR0mXQYUb/ksEVoYg8SSgXKTNwGmHRVsCEtmgGI4NhLTc8V3KsFTb08pj9UMTEXRq7HdCbtx4ev
ijK8ApVj8v+eIc2f+W1gy2iMYfLJYDhAAjkyNKmFnsoDuqcD71P0sVJrJJWvVZ+oM9E0n0I85Pc7
eb18r/9r02jItErqhWV9nR6FHLJCglP2DerdQKkMbvWCp+zJSPDKXtM8GQOwiPe6+o1AyC1ySIz1
TM8QbKDLPMDaJiBr3clU5jzO+vSF15Lx3apbaJQYpkjXQiE0V1FT1GanA05PVH+JmfM5GX1+QIyV
UbMhebjaso3rrLlvvEy8Jr+CsiiFxq0L7SOqH8cuh/2jvOp3bBD8Znh9u4tWaiG0ximlcbrGyKQq
oLXIyCsCSWZ40L5cTQHNfiyiCQPZt7DhjuTwqdMI27q8inYBOiWlIKL3CJLogEXhEmsxHyay1taf
bIKMnxu8lyfw2BfaBjYFZ+eVKpn2yr477+L4hbCWJzT3HieD2WBr/Jx4HeDBG4GJf3YnGrsQTh05
mC7lejj+LVrmB50qqcO2K/F/eYwp7ARxqfS/H/aRCGzTekgDCf5OyEWXSB79b0/nlVEg86W/uU7H
GswIOY63jl4o9ZbyHZu3L/YMRDW+6cbstoRmMxKQiuuXxd7FmnR9SC556xV2WUmhcgXC4VQChZQH
9ce+g/3DPRfxPS5oeQTXJtXnTt8wW8/J88QAypW5FV4BU8rX3YxWSEh/OU1G8bDWH0ihBPp0x/cp
UBfotzbrxsL/DX+IjdZtQXkholEZXRYKQJggWPl7tCH+h0FM+0Qi4s/PhtyhdDiJUzGCiz8tzi8+
AlCXO+wG4gKsJiqUW4jY1RmiZURUG2Yr2pEsI+O5icXaax1UJozPX+n2e5W+mgAKEpKSQHVA5P+1
S/jBtsZ7GwVp7XW+cWObjKM1rAWTnialhD4v64XyKNaiGQ4Mzm+mAPmI0XRUeZhD8JrPaT6yJJJu
E/w9H/NFyKEC1zAilAN48boYJZn57osiiiE74e7/tQ8vYKFFm/GXk/k1+9jSHbGJ9Vd4cJoC+7xN
7RaW+47gMyoIqKdo7pLzU/KGO9EMjgJC7uNJC8qPmKW5KbmYMTs2MEt+j2F2ggrNO9JfEbSYVDtc
Qk11NEH3DGFcyBI4HCbc9ZGk+htQi9D6utCtVpiSlD8q25gxH/xWjno00mXH5hdvW+5ffEUlf9Q5
/WG4x+I5KMhPJ9wtdWilVNaxmP+mHeCwYHDQK28SIZlIYkkkxOgMxS1Z6Dxn0l/P9LQ+zMEJOdxT
51vh9mvIfCD9AWs/dFjeU6MInNtXiiGVV25TB/yGeRJI1SFgdh6SMj5BPWDjHPH4ft9Bv1snMpTQ
rTNJ7G5mnUWy6r4JYZ5MJVBu0JCGN6NfvSFMgStSQG69eGnUV/BqxPqkdjLw7hweyUuQ+k3nOuxL
fk2ZyZONQ96zS+8V5YscquQ3Iueo+KNLtpe/twuWMoox2rLfMy/QFTPS4CDze939Y6UfIuhjDPiK
ELpbD9iqaESgW9hGPXtD2w6czYXTBoLOYKgPi83iObv9gyLFvRC0laN2Z6OSdkZx/1OjOgpbUQ3C
XNTnfW/lwrAF5tF+Pizg0Lfe+IFyNin1vGJjX4Xt5bKwZnSY3SvaLP1B5UTam41DD5+5fouXTEva
LhXfYYl3eOYpHmyj4CeeuLZ6p3tK8WpLa6/yW9wta/SHioGPhCOyT5Q9W+aa/c9EjwsO159gpxXb
Dy/g3Ye5k2vdK1UtQeMbHrj9IToWwNTvZ0tPKQP41ArnMgsRs6LwSbYAjjB6EZr6NjG69Z70DqM7
hdZUer9tl7z0iDwJksiaJ759F6CQ7dO5raXJjsmaj0ieRS+x/dok/re0qkBvW1GAIsWBMeeE3jk5
ydmBjHANV0hrnB3PgVsq/cB+/F0cX2A80G/18esWCoYbhDNJpePevo87OT/VhztMuMI2+VBZM9Io
UCou1+ttf846Mxtdz3GqWK27DPnhxkvLTYUYKF7cQLkGRDhLrMYby1kAdom9RWyv/w5lCRvsg5ZU
IfLvTpFdEY3Ogii8S4yCSDA+VbnmzWnSfOyxk4XMXrxQsSU+IDDy95dnU3Fegwd68+SIw6vCcnvM
XYLTy0NngvMevGfYrv5TiEUXTp/wdJxo9CLMdujup0fU12p2jQhk3saPWVM8eP2NTw3VzyoVF45k
udTOZBftjqcKoRJERlO98Kgr6sJQ37LkzbZWimyOLADhuLH1UmWKlMEdTOU+G4+muAwUcy74GBGG
wXFcAEOxi197spru3SmBvLE6XXyRxZ8W1jnii5mCxt5UVKwFtLeIBOsG3gtSUmmR6fcxHgqR+zXC
6StYp6nSGqQsVdO/7YC3egZ3Zz+85N5Njnw5KLCxXEFVTzY1zdfAL4KefARKbLWdY/+u39ySCJxb
hF7B9oZtuy4jk4XSMYOTbL2ukbGtwQ4QoWLuR59aHoM9bbW+qqWTdct/Nw1WcVw78g9bKHS5UI2+
veX+jas0ngPG6EcY4E+KJmkk82yHD8jLnagjGEXL1+8kzFyetMITjzNN9RD1owzmMd6DbKIGjLCk
FpHr5v28fmPMHuK/Z8CC2uVyAeYAiGbfVmXNOfFuMwxZ/lwL8SpvpQ1Ypsanfoxx6l0zqmTtwTeI
F53+xJ4EC+vFTWi5z3sGHcQZtcMNm184VowACGTHeE+Z5UBgW0yNuqLPnX7OYbc7Vh0CnFl8qB4A
vackLoBXO7ng75bEbaZgsvPMs1QREhnkp68hdC+WFh3IoUSJwdpPGujwE1MAzyQ8aI8m60DV5YIV
VOZe1aWZVQpQvwnh+zEeEbrHsNyoe/iHb+piyGu2zBaVcbi+IZ0BTLxqng7ldvNKZomt+nruk+nc
vSuprKJRbi//Z1XDGFGlTp6EPl58Ej7NSAVoNO5tO6Nrmg5b6sxE4xZBcsmjPxfr2Flw6co70n1B
Gmoaclp0rzTKHTLNUUWpSdu8uZMeUscGpQjoML6o9fzgdKo4v1VP8BGobxtquMbMPQeFYVeOoiTo
XIWac62MlG7FJWgcv4emL32TWIrjWIQqwp4Dct+ihe+yt/EiVRl9L+W7OyJcCVtQQZpWVHyxIFL5
AevhXvlhOcBrAV9VTU1W/YtTtFXM6dVtZ11k9qFJq2juTo/4LBiFUCLUDCuTB0YCW95AJbM9Xx55
s6v96cJHYDLd5APCaB/hks4VX85LC/ORjWvquRn33tKRXzGjzpZ52sfXrfmFgbgw54lYSIMlch/H
CBWcv4Wb1qSdCffw+5OUZuHBKOb8cJpox+Z6xbvVAwNIkqHAEH+nFf0KBX66Pd78kX/XnbgRe8uk
1XTrBA6cgMYzY2L7UN+u8c32HWTSdzzc1CVwovJxjs7cet701rpn5UnqDrPdLCjpUBr3W4sQ+sX0
DYUaPc+zy+8H9poE/BF3p6I4BSEAzPtvtPVrpWk/pxt+rs3ob2pAvpbxABWuMzvKMY1eFTe2ff+d
VjR6w9kGxrQGi+FZRDqdS4aZzSIZqeMXK+vJ228IldDxvH/hMbOIM/hqnVwTgRpaqtHdDlbp+1c6
WsJ0LAxf9vPKz24lAHHa79qoyUqx7GfgO8WAvXRIlftbmLqBgx8eivNNGVa3IC2VE3jv5sbxC3YI
g5a9e+OQE4GV8C8Mhhgg/WgXy2quTcmRO6DtoP4cuEhZlFBJRuRWOrhQ5Ckq8j7ngbSIvxhKIcsu
riGa91FPbCXKo9MqulkQ+/Pix9pwrWlzh71C9ObjrHL0Of0/+lFvk8DS5luZPjOAO/mW2f7t0eH9
N1sZBuFEH60F5ie3IWOxBDdUsyZrKCbgka3o44PfrgDP11pCP2LIOKSqiGlFE4toL2gJYBGrtA1o
H+kYZ2hMofe9McHpBrpnlm347/1sDFGlQavYMs0zgDYC90mSfX4ZkoU8lnAFX6SqufSf22e9ErSx
k5RepAALLoZS/w22MoNz5jBFnKZIk+2vWJOd1C7qoT4NYxtSgeG+G4PQQTnv0pIPezhpVFFtPKk9
J9488JWwzNv1r0bq2wVwJc3h30vPsbfOkirfmz1npQDDX0g4qe8trBHSjShuHMnCMDnwIFy9L+F4
fjsk85hbZ/rTGS8GO8l7/pP0nxlM1tEhrg0wOdMmFMLZQs/vR4uSbP3vtIi5lIFvq3Fo3GA2c0rx
MIvX8e5P2fqONVhNvqW1T4Ak2K7cEHnSHQO3FYHYG3Ct+MjKOS34szJXxaOQURUhkfkMr+9hrAo9
ZDHZ+i5cYn9VBFBBHmrZb0vbdyp2RpzBjCBlfH2o/dsw3sk/CpH5Kc3XMwDmC9hB+Ca4erj8I33b
XP4jdMp1QDgmY/QSGx/Igy5W4ZbFnKlWKyD3JxPBsw1+SCHhUh7K3Dk4MxbCkSnaycsnM4hcUqXZ
sM/4cllh85gz4ne7ageDBbJwd9laA4VrxU1Wy3ZXk7lZG3NAk5HrQEAc2KzbMO3Rz2Qr9uI4rdNy
Sj0R8ZovT8FXj9hDvRQq4Tad8fU4IV3lG4zlRE7YxzlAXgjWi3NuZ/rQVjR/g8TZtD6AmefCeTVB
bHpfaZMoVyhfW0Go5ob7FDbCZacXGitZNo2ofU//fksfhRoC3uXhp9gkRXhTMpTJUZDbjUVfvvyu
9R12+CfNH5Ack6tHY4kSfcuyVGZl+f26RAcUXHBPIAabpb6XkMvRDsDNybmS4uLjrokavJp8jokZ
ppCN+h3owS+I6F2+RXTnMzq7ey8e8mvYgsJyX3j4sXxIRvs6ac4gnjMd5O95pF4Kei9js+RuJlzf
PkzqaCqAHgFK+RTfX3cvah4fwOY04BSr4H4DA754EqpsrRseGq0qgepU6USQhhTyBoYV7/VXyLAU
XkVdbhirQo7c5MxXn5JrDw4EikF+i5Nfk5Mivve4cBhThQk3veCbPkZir2S4LtPLQAf8MCr3m83v
1ZeMlUCONquIrLTOYATBtENTxpZEEjWIJHjMwyrR7m9gg1i47LO8Oo6gyJ1kI+tPnzgRXyPJhnYR
K8F6Vr+yiOfyubWf8QHU8hCpch623ManeaFqKx/ELf6wKyWA+C7sAFs+fx5ljFnvs76DjGJx7Wxl
q7aoX4iN3r9d0bD2jl9qnF36hhOByC97dR++S8sQ/at+kJgxxMJytUTEmGe7bp+2CWgAv07IHCi8
YTVSw1CeBXgNZFeYwZF8T8AxVSGIglWDbPILOAUp8jRDEUdRSlXn1AzqQP3bCBPZhFwT/WeLPEmA
rD4jDvmMwCaSvlqCjmmZVYTMJIk1mb8MyInryoUq45nuXCDn5s6Ecj8EUi3kMlfdUo7S8FJsuXTm
V/fSwiuq2MYsGN09JmVdG7fgAsy3JNulk/JvoEmWF6hLxAZXJ3Raue8VVRymjZ21PyEFfvvVe6on
eTVrILn1F54yYEDwlhdPKGV1rz5L7kK4SCzIBSJEaarAKomceSAGbVWZvlnM0qnPwBkCSsIha9fq
iQbagqTpIVC01YzgTlYFHiIkN+8iUbZCINFRKmKAaKXAPqpNBk1HVopR6pN+lD7C0EIp2jLL85ot
k8ZA1pRKbhoymquJLrmIClYKu3jRJEf9udmLi6+and+nZT3GpI1CdBIS3PkFTE1bS5ezcoMbiXQU
hOxTmKedQC6tEYBJSpoOt4uAFe+pKfC6vq2hOPf9gFntEi1jCTLaPayk27AfIa3CawLaleyPs302
P7sB94eZZRDUaUCSmIEio4ocFCqlO7BEE3Bf4tfzGWUwon3lB+sveZhKk/0ilCQG96hY0+tPLC5q
bUHxWdX0GVIAwuh1sIhsTdNL/uA33mHNw5nXxxmullXP7uUC/gZrIb3yoAZHV6Gp43xg0vbsTqqk
Og7gjo/oz52gGOK95Wgdva8ikGUWul4PpS+lkmVUckoQ8TkdUXy8DfmeYWWZVOrHAFfRhtxQC58A
ovct0FU70MC6Be1QSYqsJP9lejbJsiMHWuT4Lm5uXv7SM64Uz+Dfr6H+fFPFnFwhUbhQgh+IHbc8
KVoPOhRE+pRL2gH0SUjGJd3FnXquZwZzzVil3MI6et9LLdyoeh69pRpZIP7x+y3PZwcj6NNngnvC
76oaJYAzMyz1qHZmcwVpaCEDnuipRxZzJJ1leykWD0lx46Bbde0Lopi5+kaV1DbYtmiKzWWoVlrm
TE2Z3vIQKM8+Do4bX0l+lb2hkchoG2MqqNEVatIxJd2SOuORR8uOx7I/89cjv2+K0QNfTvaDRgPN
w0VHbbKDkO0deGhXljw8gUjrN9JVMecG+SurL24IL7f++v2mIVvLWgwNrtiJ6a0P0pa54kJpv0Cd
lXO9yfk+6gTRTElTKeIAfxN9PURkAn4trJ58woOrwjUR+JydEaS2/xFKZl7GCKOOpGCH+2VvZmML
zNWBA5Iwhja/ZFp1Bpgl9Lr8NR2EGqFW60L9hkofQ7aklvJSEJ4R07+SD8GQn9j2mP2jbXE6xDAd
DhKfTIz6WgPINXO1SEdp1TvN7s+ZE2KgPJTZ6Jnygiw3BJM5U7++qxAJ+P15qu8Opv8N4TSXEydP
f2KdrWcqrx50fWsBwted+31/9t3wuxryQxbCX400sedDlEyYWlS6uQxw9zOaaX30VCBVsoPnQhoU
2y2fXHTqwQ30cF4a2akApPFYJ68NimBJWmg2QtlnVT/+LOuFHRSF+PQ27hBlhpkG+KgULNAIWYSr
iDDIrZuDZJ5LdKydhg2Q0M+0gGKXSL2Y0NhKYDmGmcjsXGU/GnfOtIVTBN/XAEhPi2CAd/rh4zRR
SDQMkoJ6ZCYMSChXqaCEJ1DR9ezj1Wo5v/KLbWZMH7ZKbRhWvtbviC1OVUa+JjqERuw44o5MdrYo
4NruC0mA8L1FlThonP36u94JIgYn07prILcapl/2CWPYkF6PxVJRS3bIqf0O79j3C4fUTl//R2ri
XJFsKyjYtN9KCuY+Gr/jJrUeBVgpygha7lJz7+6ZUWvP1zgyPs2J++TeZC4TNGVNYKfZ/k9uOfOo
+XrQp8jzwIOIDc5zar+6b+CY1ABYEyDDzO7KHB7wrKu1eVMNpnrXZmDKBXt3N8d5HMbQ6jDSv9ri
MHuj0u4TDTZzBOp42D5Cw3PKYKz7YUcBwJ8kk5TUkDAuWTMEh6GDJxzKEY/P6oIW45lMbwBl1HSp
RGokAiH8FY/ctmblCHnj0Yfx0xhKXB+UMELCeAUWagnk+f/De3cr0Owkhv/VCwRGbX/Qq4ICMEJg
MtHfOy+WPe1sElJL4TSOp5uPVkMoYKst8FAobWiQnlL6Hava9QdL15OYt/ln4ZqGY3y9H7kTWX4N
3HxrlAeyENGj46CxxYHLn5agK0slOaxt7R+r6WUQEyN4cN481D+9wayNO9VYIOI3IKs+/GkwaTDg
OUFI6ZRAnyigvFRXqwZuZf8RmQgEGn8MG/viGczAAbBkYvHNBE6c/uKrhiUbLUiJhgY0/sjRVHiw
FLqWTaa/O1vOX/XPwxq9NlD2AY71G6yeiedY/S2WuPH4unsXPjgjNzHcZBZFE2J0vDA90oUSDvW+
lA5HGT9Omk5ooLilUXds2nnmOA02gHWPN+xmxoNtmz+heKZAkLMsuqPm85z5IrAOElTjPc7KJduz
cWoKcbt8qgJRXHS0n6uI3LEXyR80t5jdnufruK+OxzK7nNmLyuozqQKxGU0regQiWoaLNAwaPoQ0
m9u/cOA8FQYewVjxR35Ibd7saSHeFtnn5to+wZc1sOkt+m3EXUi/2xSfsb66wgQg4cnDYPUQGMsW
2iyPdIsFKKNqE2fXrOma+YZAe9Y7nRbNeWVZUmljWzGyZShQTXvqg6xCs80hOi7HUjESixxGAtkx
Mse2vdSFBDyiQLIh9E0cg4QLX9lAs8aLnoAvQ6fja00zmZbpxwyt4ggEgJpOliXnJZAhGPOBmorB
e3d2h8O/cXO1nHrL9TBPgUMVYzxlydU3f+E1d1TGASsO0cPw7wGAxOHKSw35pvyKuaPu24LdrpV3
z3867QRBw7sRvkMtHoj28osGH6QqOy1RCB9TxgoOe9TwYEsviQrwHkc3HoTTMaQ9HUcqw7ivuqQ8
4qF85MFf0FA6z2i4/CAd8vkm86KuX4/WLF4lANLsmw14xYwpyCn2wNCTtZ/DtPio02vPyO3Rwntu
hXJxdhV9bHpR1NYV9g2FYFJp4ZEdnD1uWmmqHFgO6aIzPFregBRZMqj8jSKxhRxCuplYMLDcrbHD
dmBJcPbqvi08hxJ8FqY2ro/nuL0H+A+vet8TKVBd+HSgJYTPe0R94gLOHWvNSJNan48ITf3TE9fc
CFRzPvNxJdhJ4Sn3YclWMVdyEBbf4JaMKIhhBbCMkGLjuinMJJqad04a/MVpp3xBdJ3bbBg2Qqm6
ak3rURcX3SIQ7aPUaRNYQEdpJAANTZE0+q5c/7+U+SzfjyzcJKW2xK1dftnbUoDIFVj3p04DPGLV
PHEedbtn8Um5+hmaK7+5u66pChid4mwiS76mVL3DYbV8f+FFCtarn2midYg42qYS0IFwuwADt8JT
/YaPcFGxx7NaaFKnryjuiRMqRWbfI61BprIVnJ+a8tQM5fssz/nE0l82+RHRzPAnT074opEvte3d
w2M3ftk6c4tWjS99fXTP/q7+FCjKGbvxj/BeUoQ2xP6xc4yTxrG4i0ejUP9XcY175/lnj61K3yVP
ao5QPwJWdwSNFUenZmKPQ9jneiWYXisC1VvlXgy2/XLenc+qCTcv3iCsVmATBEuorppZ/a4qRbXB
KFa4eNrcGTUfgcA2RdCjQo+GaoQFTYPMmE96mCk4YBaJPvNXMfhOoRZlFDJl4FjPBZbT2mk2TbUV
ug00uU+QxZDOFXBJdFNrKd56fKSLt3bG77O6HZFjrIHUFXzffr5fZmKnQPTXwbvQMmqAhd47nGk6
jJKa9B6Np+r+8Jus7Q0PcjeINJ8NrUAJbg+KIv5iVFT9JlxYr9IUTmB9IK3Lr38TilES8GNYRajT
5wlDWM3iUA+5xp6T6NtAb4SerYwEVo9kUamPaN1tP3vflvtW37Q8Zxy2yUQG7wKOLqprzprv8I4x
LKH/6eZQIY9t+gMbP7Hw7XQdfH+ha3fq64rijK5FKSm7Xxq/Bt5Y0jtC4jhYbxb7eTMzLbQyytjm
mhEpdE89Q+JPAh4Et4/DRa1oB8xICFEMG5NDH6I4etIdHAOpMWa6zTgy1+jxkKRGe2Vvks4OFg3b
B8WtUOoQqixNTRUY4tYYeXWqBrvihTB0dAO/4nUi5lPKPYonFxKXwy2hcEB428sNzRwLXB1LpWoj
USLg2ZTKT7gZQMyoOq0xL01OlSdhaObUC4NSuqqrVMwr1GMtPDBxkRYRXRBDqq83uGwzdQIv7FE6
5VbzulJx++SNBXFVgyb0tczodGxJmLq+ovkKZqbclwNhkuCA0+eQDneOTF3I/I60oOrYuCmxkPtR
OFIcS9iK0rXmm8Mj0Cb5FhyMzWukZHQIYnrrRRMWxlbu1XYuXmnb+G9e6Ez1ft/M7FvS+4BRFLN5
5ItNqR8LtSJdQKOpikdJSibmBqzWOTSmDsqJUiC7SFibPi6ep72P1t4US0cCfZKCQ0F/ScBoQkTz
78KMv1DpFKfAy1ZNgH/pSyG6C2zGhC9QxmMc42R+NIzZPGAgEf09FiOrFfxkzgrGdeLKUDDjcgka
CcIr6mMK4VA6RgkyGjWjIUoLcf27yKrcc/2kUwH6cxCltZhOSTJITcq7dBe3rbBFi+Zz7Xv6l48F
hhiUgBugB4bXvAhkK4u6JTrTX944KmNXSM+B0QNdPRl+DiD6KNaL9Ky72kuCt/03NODvJPCRwwPS
tRxhOGYJElQlMZj28wppBcVbfSjlsh/M/BDpvf7ScGYHBjfALQB5EPXoXlxwMNA5TPaMvGc5AxtG
ft+TZDjrwCxsFDBAIwdRfuX66SxOCJbU20kOekWvbPkSIeu3k63mD0y9zezsfJuHfwkgHLswf6wk
ZVZ2YFdxEQo1yXDqUYYsB6HEGbisxqzVma8x3vyhBDEtPkYObel4xlpwi4pmbvceRJgUbCIVU14O
Eht/h724UqJOB0icFlqshF606G8japZJ10x3UCD/8M4KFU0OcmSbKwjn2gh4cNh58PP+e1AvgbcC
aZdr9Z5T2mwCoFECUwUe/tsZ0STT7Xhfc0ytzTlvJlQR8fJQOTJzN+kl0hdtBARxZucnzpMA+rFw
TSS829Oj7PkBURzOUNMg4jONtpkNhLwTJxTEZlUdgv8fZgpYZkLrO5/7JQm9ILFyJvOjQwym2Lhk
u2hAzuoFkl7M9Bq8gpH/D5r/7EUmeXLuuYe/uYl05A5vbO3XJSDGwqCI/PzF08vwE+utOg4D2nbD
ATbG94AhA6wOjuLsLyemSCXRo+SNWvwqhumj3o607O3L3VuRGOBJUjN7LrcCI1X5ElqyVLnbDW3w
/MKEFgFBhRuRSlwQikrHGve1CooMiSNKGv126dZs9NFQoG38KzZ0UyaMyPetfVkku5eEFNafCmOX
HqQlXrUFDWhAlPzxpkknxwoFZlbnlA8PuG/5azyYkiwYt1iB512sowGfi7pSiJPuwiVwZGl72G57
Z9BEgn7byV6r3AOQmjROe5whbpJEnz1xn5Xhq1UBYFTbjH+n/HzF/Oc9atYd+3ol4g5YhZt2zDoL
P50jolFsQSC4/pWl+NiMjiMPMFfk94aJferliF9Q6N719AToFSCGI2vBE9F3tyNpFJfODDFrQtT+
U040jVyxT7R7gOo2WN2bBqGMxhPLMtFSYaxDVM5JflXcj6Pqz9NxlqaE1jdd+woj/kT1uqVV0p5D
vteR8XL75HjTmUkPdgzc55WCXpdutdhCJt6JMDPD1UsVdONEe5L7t99AE+gEHjqVnM14iDpX/qE6
373Q/TiHqlqzHG3ml5MLwx1TvqCTMomcZT7lKRHrXCiHP3yQLOfFaMRXHtH6/rUYWykNI7PghAmH
UrLI2PqdQfZn2gja5tFVhh2SpQHOPIISfnjtIP6QHZKjtXup5o0U8tWW3fzbbPc2G4wjQ4jV49TJ
NmknwkRRjrEsbkGtSgafEijBgIZETx7W1w46yY2/D1eNEKNXku4t1BL1MFzGilF3BLb//PF6Y3mD
mmV9DX7OBDHVm+mQbSaZ+cL9HKz2TyC4jzxi+t4wABlmDmq+hXiUEddSMzsE4YQvz7ebwyL2HZG+
BvaGoKMDAo32zbCouEX88FdQJMpCGW3orp2XcB4kl7oFBD2KOZV8mqoHIF29TLrnsDXSr4+o1Vab
qSMVEyOmBGkA5ra/7Kwikie7fiP1BK+RmK5a61RWzfFSJUpaYlcGIDHG64BE8Dz/XAjZSqKn/IjZ
nU8+HjIfevYKTRBFzwvdArYPppeUrcMtt+02z+sgcRld2Yca2zG4cKYE5maWHSS2XToMODOoDvAD
qZ1YhsN4/mWow+bPHLT6QSwuC2DADp//dVbxJkx5Wo3fyhLsnmfww6e5Fn+To1mLFQ+LmY/RMbRr
VWyn4+B9zfGvxanIg6R/5tsaNdd7GGYHH8Wk0RGRujfOXpKBClUPuHmcMZ/DddljAlnZOy6E4Xdg
P9HowGkYOK9QXeYshk/0hyeAJxN2sknCMzpgJc+QoQKqm2TFP2dZeXPzsBofdO/2CsfudQB3L22F
mBjCqtCSXkbDw/vOxbWhWLrq+d7Rz7winE8rXf0JLTHiThgS/mLCmux++mBJhQtwKZTZaCxupdob
3srGm8e4Gi2rMyNP3hyHoT0RaARRxaAK6kl99MEzgUEH4VRt6fxSALmoPRWIf2ghOBU8aLz9ImnP
BwPkM8NzT5vMJc/FDI0wjhsQyPkkMsilkAk5qdN13gBFKhJ2v9bv0PGQVhZtuKg9VPgjzmKDPYgi
LsP+Zc4Zw2hxYpUUuXku5Fzz1wA7qvzsLKWnCHBSsymNM0pa2/YuL0k7avsD6Ej3I7iusaRZ6moJ
fsS00DQXnSZHsiIKPtONXRk+DnA/D5bWisuqSd5AP4B3hM+WOe5Cgbo6XLU2y2uI3LQaDDs10Vda
415foEU2z2deMumtD0vfcy6tNYe1WNhTaB/wO/2IBPXEtHIn4pTPdIuew2vuo3GdzjlCiw42NLr9
1V3gh/BVQzDozVTHuRUuAsgcSnEdefiI+YyT1gJZ82wISJRXtUUESg+O0RFCUG+3IbPi/YOFP5Jh
KeOp8pmzvVDo2jMyiFpxSckdRid0RSX8uhxLCnVjlziPwEMKCnek/7jGlBLl1sN20481oHOs4lWb
fC6mRj+8YnheHAQTdj7j8o8BEvs/8ufGrhOflwSE2c+oPaDCEFmtBQpzOljb/gvmQGHan8HhrruT
cjfO0XRf4F8AcU3OFc2mzhQIYoU6tctn/TGptr7sQAlYJ/ztJrDlVx/9Se4c9mUyIg7wd7BZqZfV
KPv5O9mjijvNp5stz+vQYy2/hV6R+LoXWH4MPgfd/tzgnnoPGaeURxReVhENcB0FdXEOE0R9T/Wn
t9bfV4Pikr3Po1jLiSgRR3xDuCaHqIb1osNme6v8zHrxLVq/VyzaXA3+SNADwekK2CaXdygQxSxK
xfCWprl/50TEFPcFQxwwu4HZZ/roWMN8/qr8pZ61eJK8m5ZBy+zjLmu6WYIklTD4sS5xkwKDG1Lb
L0keBsC1PFX9hbaET+hER2iAq58CU3QMgZLUR5wy/xr764u6Zv+rpD5fAaIDqW5XgDkcuQf4xUlr
uPm1Ud15WnaELpDIgnAijRrK6xGL6bu/tPO7Zw30QqKJEtLxUUUPYn9ZBTvEkeMLIOCCQOuQ73rp
p9N9VVryaphUHyo4QAlcQcj0StrxAhcQ4Vvo8Ju0APZ89nJZ/pFT0tDCOJBpxK85J+mCA0IMFygC
GwjNcIbatwoJUTSVwBRHppLWVdgJJVmtkxrjXHzQONIdYWGp7HPEnPvdDEJ7rPkHFl+TDMH9Eq1D
ldzMpdEXp+vWrnUdF0/9wH+mwXr64kqxWVGoR8wQXtRBLnVVzC2Kh3nNzRdu01qDx6iMcfqTJIyw
ObM8wusloHSvO5EN44SF6QkS3ELKSdstTpqZe6o/fE/J7Xue4LuZX2Aa36+w8V7+B16/PfwqNb70
lYsrRHEuG5WtGRGFm+43dXNwimJXX4TvNwiMUjOs59XCuekOkkndXiNKmteViEaT9lG9k3xMODf6
NTz3NGUws6y4KRvs8MZdNgB8o+V+5v2iss+g+V2VucQWbkZo6LU+HYtnypYSKPWrWR3KuO3koTcf
QjsauTTjCwB4InVA2LnTMRXUESZ6H1p31u1NS/dzJHVx++KJxuLunnzDH2BCSgRNtR1GoPlmyJE9
/taqY6G8ja6L2h/iBl9aOG552pFla3MpvsWbcQx87LD9MmZzMA/+GrpW7ndRbi0tHDMisekIQlhU
T/e3ALOaGoHOJL5XX7t8IqT6QAVSHwUIFoSlz8o3Xfg0iynfIejkzQ2+tdWV4eNTa2mFmApG1+f5
QvDNeochxq40+nbAfBrI8Mu9Mgc/MDaSNWCtSqPfd/YjX8xoJlK350Xd6gpiTKi6sNb2TRv6APCZ
kHxw0WwvjArHjRsXwAiwcX/AbM4Wnac+Ssi8y0PkLHQa+r+idnx2zzLie4Jv56RWEJxhkx5Kmtli
w94dABN9tqCv4KpfvFLNr/otJnzcS4ELfy5muX7P9KGtEJNI7EAO7mOJ8Ow564bWy6JgWkuSrVH2
sMhfOteSA/C8DrEf25LQUvzvyIyw2L8r1PdNvY9zAzvtObP+0zHIhi5EiLywN3axDxlew/eg2COy
+CCFs83MwT1gzfKAmy4o5kGL8iRk/oT/w8JjFBasYYXvHq8Qw+qi9MP8uWpxXT5XEgJmucxOuKuk
iVGtHlVnTsdD2UOOtMRw+3OrRWB7FgorGXlZFAvkVG2dLZQa2UGu7Bj1Vvo/tbfmLL2GI1kLBX/K
/IOiIGpz718F8xhXRNCxCzUwvV5DxW1y4RIFjxEaKPMrVyAL8ysYyLK8UJ9WE2TwS3e20zh5HVWy
5mviC83vJusNhJrYEvRQ2O3Ff+GtRlRGDVohO4gls9OV4FwtLMyjUX6KYFBDyDJFrqnE/23ovEFl
0rJVIFlaBwHl6BJBvcbU2rQKcRZ15CYb7Hh6czZZnxM1X7VlTQs9T7e8+r+HK9bOH8j2CUTMQfqA
qQs8E4azN56I5tZ3DnE/9ZS9lsHEs8YkZWWa4ZKK7BH4YGDQKTiiUVgpR1mDWELOwl4MV9S3BfgV
XLY76M24VvZnTIrJRGfs8C5NcwbUAHnK8HqZemiRFzduT5yutV0O00AOAdXcmaiNJCuC0febMm/t
SOoUdi2Jm14w73ijIBEZWzjJiXCsjLYJg2lzAVazd0f31hwCGxG7IctDJQ4Dadnb0llxzDKOJpAB
WPmNRseCjM8gwRXeckdyxAkKAX41kaCVPQR2JhXG6cwZI25RB4bImH/rykZN/HQwboFzXv1UoG5m
x9eAJU0WV5DZmmRTDf9kAJVVRR5ZasneS5vC20tOvwYvNlq1UcTuYI5UJbGBMywsFyyIpd3LkhZX
LjRBefhwWqmyyBoU2eunn31PKN7LmF8xL8UdGorkukQLeqREip2yaz4sPzbV7YHSPgzvc9A0TLhz
knis0nBICGHBrESwsRba5Vj304m4E60ipkSfhxFtL+k92+qGJwqPRmyxGI8Fb5qXW4pejbs1xMCd
8viACWuVt+/GTCWFtseT7eWXTerCfivK2NnLVmwnRavtQq9MrkfQSDUzqi5cckOJ7gVm+mryZ2U0
BXPZIooazovUp7OTUNZuzstsfZ7uu3GE/eZ9VVrEL0lZGMwuG0m05MNoIvZf4LqASvsPg7NFMlaF
U6TfnYrhd2BD8yE96ToQP3v7146HwkLChXQsAsfmnZDrGSWXJlMnTyVQrQPZXsM4TczvADLmazjL
iDXojge+za5eNvPCYjFxfaWodv12LtnaOUPP8+ruY3s7VgwuVv82vdMSvxlRpJyU6TczCpDtHlwl
w4HeTkHP/PYfzAOxvv/qrNo7DQme5TNqB73BCmjW8Qu/bDgp+A+d2Lp6g+M63afIRr5SkVRWRzCk
9Spb4liEhPRBxa3u1lU40pTPS3BC1C8gutgWPPlYkEQMZ6XSJLEZaR71sZ/MYp6OvsPQc3cdCjd6
Y5ZrwdqCRJAi0FBFYGdT4BEdfWSlBPrdzThkZejq5PApGxCft2x0SyT+mzUTbmDLRzsfIXbGvYVf
X6o1WY1wR5rTjs3mMj47eaF5lrsDnOgQI/XXma0LZKdd4rnY0Y1q4jfjP9pwi4zSGCWOoxbU+Jdw
dKxJ0A4CytvXDRORNcLv8ed8NMhRD7vdSz7IRytvvxedX5d3Z/kKSxrq7amqjLK5k7KMK5lx8zLt
8dI1NcaGILe8WbhqEc3hZUZ8sYlS2kXqJaoSz7V8enTwpPvXRSI07dX2iS19UQA8f+FmLkDLB/5R
wz+7bjUVGqy8zYjDKiTBQCP2tXS8t1Qn2wYk0T5BxmhaisSRFBg7TOAOegpMJfgRoYP+l3/rELWU
5b1Lpk1gnNxOB6jVk7iQG2ruOaCfuveBwWDkbjp1dkdu5BgZWpV+otHQAJQAPsGBWqkT+ivDtHmU
MyqX991dYTz2UTYaiwRrwQNepNgKnLklDXhcS9r+IeSOBU5p8YI0ZW52/Xs9iAMeG8IXfJrTbE5e
IuJ1Jh7dMz3U3O6DWtYcG3EUE7YbNTMuEvYlkWnyIxamzWuMamv0FZTAy+FU72bemGxNYg/6KobG
qtQ4Njm/yWr8mpk5mwBBr6p+/CYp9NJJ80+ItMUv9sprlSYN6itg7zYI7PsCE7e43yxNf8Og1fLE
JTL93uFWg9Oyf9gNhAIp/NrpRC3wRLSUc2xpVMPEo/pQ7R8QABjSLfvCECPtQbUVGdLosZhRYmF1
S2tqUXTdBK1NVJr0GEuI2fYM54tWH9fT8U4RcyjlgA+W/2GRVd/fAgVm0FqlTkgBoXfN9V9SbF5f
3C85M56rGTT0735K+ePGFqyjWrmJlbz7YO9XFXdaG17JvyUOZDI688eileBbQybwAy/+DDxfwGp1
cMKKtyhK3rdMGvaMRLT9QvPMQGNpqGiXnWcUD5Eewz0Z9iw3qYlVqbu7ZildlPOmn/xGlHAdAUfu
1pw4Oijp8Pk+SKDxeT2XZLUv8PnM+IoJgPws82Vzp0sF0WNVNFXyFLWQnla++VA/InqxYjCoqAdS
cxkYggoXYId/ef4o/TWoF+zpNAkKrpBlaApV63Pt47s9siVVxc32Sht13OHQUPDsFg3wYGIG4DNU
V8fo+oykwC5ZgffjRZZMyS202SE56p2fFN3Knin0OlUOa3BvZ7/ANWe1CeXmgjYvnwLl6Dmbt5lK
IzKs1c+PtzV1sKI5YnBzDRYG3dirsaDs3tJSINPAsWj6Hlnp9f+7GDbmxotRS9IyNKF69IFMvhy4
KgVaCahPELmEUAKYJAWWcLY19uUt9lqD8Qqb6srQ4zjLMhGqyXDge6e+dQIBiiKIu5Npweq+0k72
aIrTjg0aHhHK0awQFes/JnevQCl7zCAYSPi7Fz5wvYTI71xdTk8h6kpVXh3TQFIM8IL1Jt0d5uxL
t6d1y5KRbe608D0WcEwlMgAcc1CpGCevPdgpKp8k97VYQ8UOdW+GG3Fh7QhPHXexdUNO2GBwX0oJ
Wf4U9ol6Rear+aXNzMKKFzbJStIB3NRw96MXQ5n0Qn2TNu1toBfsCTEf2Tu3NPemW3H6EM5+mC+o
7afY+lICe37IRJH7we9rkaFbP2oLA/hTbkioUCaOJ3FarnYRdo0N8xV4Jh1wWb95DWXm+GW2A0Hl
tQg/4T7WrhPN9oWit/9f1G1D8QC/Xx1zeQOYKERtPDZEkENUNjw0uzKq7RX5eNDDLP5fsLPdC0Bt
6bLGHDA0ZRMDiuRiUSEBsVHjT9LW8BoQK2lgy7RkDOq/Xtqrh3qcylgAtM8CUBnMwS2F9rIwjTxM
c7H6VoH8E9IfFf34vTRsjQWYXV2xuRystNciQR8lQontWJFHGMUu0PT0+jmHBzCaPwp/vI3MBk0F
7es8bL7DUmp1RZXrjCHHH2H058MjDg68sjO+hvYeijnqEe6xxO7LM75pyubHTuDn6OLFNe+s7sdE
vi8EonImAZ6/Orlx2EKCxXqhu13QkGoL2Ap7uVXPG+NKWWuyHv6CRO0WnwepS176Nv9NSDmERh5Q
/o+xy+v0i+1+lvRB/1aY8bEPie6iFSWbaE2s3/fTs4R5zTSPlBcOE9bH1ZB+AUNwiI9r/Wp9mIUv
iDZKwxPYpLQGhbZmkjaJSnHEdb6k6g2jZYZwIj6SRGvoj5DqwclNgnFz2SaAuo56sycaLrx3VJtl
uiMCzYrenQBsMbukWCGWCkJkZAtisuEUOrcofRb3Fj/JcY6lnv6xJvipzydRGc1lvjUjrq7XtJGc
qH1u/uU8upZEXgtWemoqjbZc9+vW/HkjukaTNzYjEb7Arv6fpvube9citPyEspMOt1wWvcMOBToG
LT/l3DcyMu3vtDrXB8ujZG9qcQtcBrIQeiuQrvx0A/HVhjZM0/x9ItrIWRaUxBIZm4YplyOGE/TW
9TYxYBdTYEJBQ6YUMCAOqMSYeUdYUORLP1gQBQ/Km0DgnQJQ19KCjpXNUYY02CGRgEQfwuXHXKQi
Cap/wYexWZjBix7B4TgFzuJWls/0GO4Ej7365qlWCKsV46CO9tQ887wLMqneoDpKJfjApT2Dh2i1
gwpnjxa8CsyYOgIBCFrpn/+Q7kUPTw6urlDXI3NCGX58O2Vt0HQrCECq4ICB6Vkdgxdx1t6RpI4y
1iH0fXqdcpubrU57MeurXcp4EvpE/MunaEnjUdEDUWp/PMVnkCmdGR64xaGCjBaQ66t5hedQZSGH
54b8Qg8JC3lS26IDm5MGdV4sQP3NGtrCzfDi+/d3CJfFDHGd7PRi5onFPdjzxWPEX+A8lj1C+pfx
ZQPM3cWY6iJkXorUtUx2drqGO7b4FLz3FI8BBleXDmKAAau/UL6hVMzWKQayg+TpxtxnnJlbr2Cy
vsXHEtUIkzEvuWrKpCnDtNHBijcX4CFun49dgXWFULeI6DViOjAXvC7tKaNTZL7WPLVWnpla814F
Uwd5r9Fi/2KnheGu8jDjwH2fIILWjpC40JrUCgUvSsVCeTDbjTKHOCTwcFcA3una6Uo7TAGWGtGI
KO6iFuXqXLrDh3k3APBweokkLL3EexDm/txvBPFkJgeDN6j1OqakUOM8GQahOpbXt55j+jraTdP+
nXyUWFS8Sq9Q5xfoTwilZJDv9gjv9vOZUPU+zICAbkIzkKB87AXWHFCUvXA9c5hwMpSlAe25V5Nh
f7uoVZqsebOYg5fBDI9f1q7PigazAWpPiNler15rB60rp3Ruq4+v0pIfTEhXqnkgvAjoS2igZWF6
INYERjcZ2WmBEV4OCDAdiC80mNBQnsZyv289qREjAnMszGWCD4N6oAzbJAukuYYPS6P0J3NQlgXZ
ZWbjQTjcG6VbD+X4mHLuDcUQbj5WYvRgo2meSiTpN9JvGuhu5nmCHZmMyipDGCeT76O8DYtuqRwG
s5DDWnlj/6w7bdMOkYkgy1t2+AsiZUtpuKkBWInbj3K1ttp6tsDxFF+JoUba7jN1IjRCj44Z414M
qcIOIMtJtyTCyFSouTQe9u76vZAT4v2b+d0VO1uEXOlC5TNzpP85NIudultPgh+kzWp8efvuX0wl
dWuhwI/H8crD8hYnHGL/x19RKfzvi82tRnBT7q3dPf9SdBB6o/CTQx4ZXM5btkrFE2tS5w3M8mVu
rdT7MWaR77d1PsWsc0BHP3RILWy6W9Yge/pulaBtIYQQ5wZmGaQPyyPMa1WJ5cXq9wd1qcTON+J5
cwbltEoNJYirHteHB5PYyqLC6mxuwxzPK81E6d7ouhWFjrW0LhdAcQQXejA+5k+XVdPqGdbNlviL
zOH1AoeWg41Ri7fPQLmUoHyM8GWpLfHAntNdAwatTq49TJocEd039YBEvkHZLdBzM89FUsxAQ9IS
jZbFe5qH+wS7/Lrw8Hh8tn9+79E8NcEQK61MppqcGvBH+l9XPFP26k4xld8V0g+9f+P3xxxIvqOv
Y8l56hn7I/UQhYXFTV3Or3OYdLWE5u2ofVdwJlkm5zWNmvtTeI4n1GcPC5Pdoccj15Xqy9YoaIYa
47q2n0J3O8bVQIPNBO2d2EPKvLQXRluWK+8muJtixnNdJAVz9Iy9XKDz+MRdAo6o8sonlBsPzHe7
ySgPhrD1eZ12TRFZKU+P9G+rR9H1a7ZFsLheFEaKUg3JId50aYm2f/TptCMpb+P+ptv8Gz7uFlMl
OQqrFPvYhk+RzosTykU6s54rNfom8qBQgCjJRGUo6mz+gV9dXQHxW5PIY/kfa86WR6uCkcbzmqQS
NjvGV7ezoXXIlqKG4ODT9ALyuWaKGwzk5J7iMrCgOi69aFElwuTFfRtnRFfMd4N39MBaerAvuAq4
qQIhUEIxS6k6CTJkom+LrnyqUSVJK9JK1ovVeN5sJFHIPKj0xyeUbsmowWfgdCXyuqJqrWyDzAuB
cg8IPbi02RZIrDAoaXvCP/xKd//ghAZGvaxY7wKvl92HLXy31x6gNI9mXyVl7WjEg38JC8C3qeL/
9gBnosRweKMtPGR/Y5XoiZ31yIcACQV6FmXuuXMlYQx0YXkMBKoa707YxmbOrZoqnyP/ukGXO2sY
TJSLjxCjGtOrUhTp8yaCWfg1RcJE0xgCkVnpBVHH3UV+vz9eqdDkuj6cnXHDdxkaNapfiX/wwylg
xOpOj71gLnC/e8vj0rR8VrWwgAOHxdwGPZ4hpI40nFnT6Wx8p6cHd2p72f0kyNfexFE315Kqq7Mi
Rd9SP62wv9m44dpISlnTVR40bVoWYPGgrFO635Zc0MC/+Iamrf2In5H5IgUts4o7BBoehZAV997C
3FGwhvASQ7npfjkvi4FdPqH8HqOgJdkmDNNujuX4BEnTkWmYyZ1FNJm1SPi5R/bg2bS0CbnGMkjW
UJ/eyOJ9f8gwtwRdsn2EyMwt5ZbzUqowXiuuYKzd3kl5BZEELbs8zoz+b6gaVMzjp7pbPn82klDb
YZWxnYRZRyLlNSFAJAQU9EBFiy8ngruHQ82NjxBjMMy0avzdEMtLAgokEiCaVRpqTz/AeK+sJLF4
p8gcdZZG6YVpLZIzUW7vqAU5wiC3/E8+bxkjlk5DUvl8Id3jU+LjRyDe6Dt+DrLy6YWxPZ7FGrtI
hWxsjKwIXb46Xpswx58JaCM0GdLtDVVz5r9ecrPgtKtVHhQTJBodYD7N0DJgUFtrbehv8/ZSNAu5
aUvMWvdeao3z9hJtFQI13+xfWxAQRbvtjAq7olA/D4nn8rxdLjTA6xKUdY3mky/2fNzW8oNnl91q
BuSJfzQxNaaxP3I36mn4SbdntAGnccGJWWOCMagAeSE973Vagry4FnfbHZHW3DY+0xBZf8CD1/K+
O/lpaX641VwfPxsBwwbvnyJlluLElgTRdpTdYfdXwQyuOf3OpR0X4Y6mCBU9IZv+90huDuyxumoA
GnCVr4e2HdnqnGExJea+r4vHx+FI+ikK+Rg53+CPdHFIPtYHtuHPcMH3eFGdsHLC5wNwUmue3IT4
kNhkElBXRFIxyFJJLoklIPvbVZ3KzcUNFQW3HUaq2Zih+rnvYeaknydJVE8W1G3CRP8GogyVsbHv
0JlPZ+IXtXtcICHq/Rm5h99LSz4PHGC2KTR4xOQvcyCspvtsRUrQrPNuoBdzQf85Z6aot5hGGm4x
oS+W9oO61oTYBbQY9mtH/SbLJPfJz2pEwrfF8iF+UTfle6vJCcPZe2b1n46xotTC501mhv98xaVX
nwlKjlAiWX9sKJPdEFZyfcxOt454hFOrEUr3a0GGrCkxNiZF98zFnuPh1qnJTsw3ewAN8CUPEGQJ
A2gYmbmOSFLDrmRlbz65caiu+gtO6CYINmWzNYxT4sNKC4sxrOdksgcTC6ADg4r04dery1ozp6BY
5iOacI+nPPUYmV5HGpbUPPPeNC7c/sIw3GUu9jqBKuo5WfHW8wr3KD904+TJRpCcdvR+Q8pDvb3H
KZ1avVam4nsNF5Lr8neB75sWf7xPwMS835mOMP9wG69qJ5zRLAb8Q2ftCUH4Q3kZX3aUOKMo7Jjd
pwek+aZqNZL9zq+DDq0K9BTxjn4Na2bqLYrAldXAMKmQ30MAh2xjS4fxZLjaD0dF7tJ6mkP71E1P
EivLugqMYFlQxONt+25cRKSzGnf14ZSMoRZDZ0GBGritxSnxtGIBFUzj4A9r9LXGPft2j2I3BUI7
2ABdx/AUlhi9fEq8NV8wwfWzQ45/1ONacq1eSvSgCFhH+gvtXR73ZficsB+LPjqlqQx2rGp5ZZO/
yhrvvKKUJYSDWRL6lGY9CyOT4kdj2noVFWyOEVWGi/H92pWvac7a9AY+AQIavqk4FjLG+8IDT49k
GdbZ05KXeaWzmlrgLroAHN51nbVQ1al3vSFpdAZ32vRM+QfA7Fm7PUikxKIMnFkAXZ4W2EleaRtq
w9xncTQMd6bnIjOXOsSS2uHsHc/jNntwX5jYUJrQtYgSgr+WpqyAGEPwU1VnwZtqoQ9wxtNXYuMH
dZwyksLfIRCIW1889HPbTakyXrbQzcX+2kO9uEV7ntqc2z7McdbcAnZC6Tn4SJeLO6IJZapoEINi
uIJdFWFy0suOGtk7FXP/J+c/SJUSwaB3D1qxwJlw/3k+Zg+BEtaI0KMO0vra1TSa7d82/FOeIDwk
ji4fKE1bZY7UyITsCRUYvCaSgPSTCdmiUxkx5FOqY1A0nrgjF2roeOXh9KyDXmCivsrGtpVsR2nn
VN7Npdcpu3NwD7jElrLpjC1ndoWz9QFV10TcID+TOEeK6xCuT9MydQqszgJbkMfe3iLyGiFA9gWv
719DQSZXVOaG/ylJ45Ej35MjsgCbh0gl6Nldo7Nqkd3A0KLc6KTcNVdEOEPauj5aVk/iUAygByU5
0neyoWDUA/Kq4Tj13e1r22CfbqFekI21dhsrI4orq38p90DNfzKo76XAfs5ZcZhQA7DgUMoUhoa1
d8sjOJkPxE+3bmuOF7U+f4TGHdOipiPY5SWNbFU6G7fkaFrUAnzURpurFeFQAZx6h5M/hdsAsLCr
REASHsG+YiOXUR1eFzqaErXDRJltvuysplvoEFNYfb9g3PrGUTl4EujZIzCcpAZC+EfjOhlI2bKJ
VTW9QxSZI3Hi3cd+moTFsOStGptF/CZt0GJrVT8geZlMLTHhEbnFMLARVcup75WnpK5dxlNePm2j
RZzEUugwfLjtBGQ/UOJpqRAFjOgXfEbRC2sLy515+C3NuKTa1DIDzTFFkfTxthlKCttMHbCmgpbQ
PZKwbYssBlDZ00usLjshjXDmUZu5vnpJNEFhDDwLcTBQjHL3uzyijfSyYJZJpK3RHZOw1QOhPqyG
S3IBA31qzdHvT+epmwC7GJaGhza0EkvZ/oa83Y1xAt/3mIoCIGpFm7FXOphgB+djoGd2wcwjiRy9
28RZRDlzhkNl+8Zpalx27Iq3cUKS1nkEUmrYJ3eiwBoo2ioUG+K+U/dmgVQgPaGC4DnAZZuNI1x3
a34Kx3dS/Rb8Wdy/KhohMRPox20c2/DcGbGYxHWe2oM4L0mEbLEMnSOWRgKGBpEY/cQo+UjbN/hS
xJL8zSBrlQR9FZIacacBceROBPkbPBQovA2wDJujjffn0wRYquzFm+Yqx0g2pF85krV3SCXr6CPl
PipUn7sHZmbRXF6vMMdIANm/WtyCyqUWFE5z/ha3vUYKrv3T0buNNlaRS2QAgl0paEyWnmnrHm2Y
iyUJoup21/ghXSb5DZQTEgCofqDP5TKCL8w0hB3BF9isWz5miwdTtRIHAFvS0t73ZNREKWR699+K
ALGtEUWOzX8cbW+MEptY938uCVLtoHZhNUIqJcgA0/V3j1pIycsY+0ID9dDWhMoytX9GatRycmjs
P+WfCJ8Z/OhDsqBaSM209piYerU2H2RrUfi6uZBwQ26SGtXahlCtTyPCgzJluD9khUl9vtb+F6bV
3OmVFP7hYsuFI9yDBEfCAfw25O0EYJmFNvmxYW2ODLeIonwcfaRK4+rF6h03f+EOpBNYLdDMMOlo
tqDRfFQWhc13cOshpt6FoBhkwocKSDZxwt2psbXRqfG5Eikk/LbzUji6E/xpCkn1WNKJPSikpLsG
dIF8QPAq92hPy7Cfj3Y3iM0H4lyGw1ywHx0400S2FBSE1yy43UUVWvkVcEutERCadPsOo1X19nU7
PhD5Oowj+6gznpqVab8PHNrRwx2EFpkPZ6cCVr32Xpx4E5CpHMjOef5qCxJKjor4rgmE4gCzYF38
MHaojd7vskm/r8fRIHEzLMMHhDkQmdvPEkRkr8Heqp4hvtkzq3QsreHhFchd0gmZRcqx5vnNPdHU
eXFnG1Nm2gfunHiMDBOswAkB3mZ+QV533x3SjdMhlTFcejbqaYZkmcPRdsxFRT4SVRQzBG/AWDXZ
5H+hNVw3mwvD7bL07LSOHiMDlMEb21jmeXkvcRGlfxyfmPVHg4ZikIHIcWuiurRa9p9w1SudATRU
hGc/zz6/YGLd6F4zaFUhI5og/9RE6LLcfa8Vm8ww1x5jrk9x8HGP9Et2ypXpwQoEhovl4VgmpfCZ
J+itIsBpPtJGvDpWZwV/kc3yoY14uORs/YpV+SPeb5QJtlWRLGQfWse0zUZwTJyQ+U9lwDydqiBF
j5pfVgXyNyhsi+Xb6dRUGnZn3xZpDe1sjfDXW1xkX4akRtnbF+EClqf1lLMp3JkrKeZuXvKxPIYG
ntpS6GcwuKJoDE9ewCKLqm+8drwGfEVKOo11asvQo085uCqrlSFvRMBhC4k0wjT26yd5Vp+Th2mi
5PBQP6HBaVDTTGONNBCTC6wj90gZYqz9YnE1BQ5fA4pfCxAAvM+qRImWDJMh8/BFIOqGh+Gv/pUn
+9RjeABq2WQosgwOVX90cZsK3d1xcLQvf5UcVH+qlHYEX6/gK4R+rsFn5EwhUqToln1HizT4KKya
Uk3Gx99bR16IK/Offr1dD5xKgZ8VdcYvpgjP+MLcXcO0dMyFicvJQZTkBh9y9X/x9/4h2ubQl/67
52DG4S4lQVb7AxQQkq9MGwJ4m0Ljcaqn0Fq5M+38TZJ7mqGHYJqFbVHBf4ML1SAE1GyZUHMtOh4U
hvxv2gsMOVtrQypv6ZPgVFKdgPK7cMiB4/y1Xs0ycaySfXLywYz/rKm15yCRiDf+yFuApDmzWGzK
ZrZEGkLLMOBGARBn0FaEcI7nF0drm+TRFA0PZyb4DG6GM7QZ7twICdnJOXswe0qxqYuN5qNqWEoe
ELw1xUJhJ9f10F/KgiZWq32OqARyVgGQOW/8ZNnOV2rRfnYVZ04w0T9wyTVJk6UmGazVW06nU2D3
mg4wEuLWQlKc/6Lkf8G2XtEMKTINYdZ0NtAD85+7cydnsUhqLCHsokgx8C/nLsLpMmsQ7NIdUovT
m4mESI9H5YC52pESNETlWfOSrtT+8FonOlqlwvaua7Wy1XyzYX02deIYOfFaRu2/ZmOgn6l3hNfS
puv/A4la/lhc0o4I+u+9VBtgWK48W0EOohHuzRiMXgUpxH8rkEOV+okjRrUagMm2od+2r+tDlz3m
PvPjrAOevav682ROMA9eFvcZE6PTx8fimlWjCAZbVEe++OKFi3kSFjzbQBicQINgg0AnP/s034Sd
XHlvcCpZWFVKJ6sZm4/mPgO/el1qYZ3DRIWNUh5u5J40UyI5EfX2k5hDVnBDoB8LefRcmkX4K/Up
9Jy57J1f0JcaREk3xRBPa014uOaGJ71XAa8kbD7tp+l4z3BcZweXzIOSAXSQN7iVVmGKViGeWJ2E
2OCqFVb6MoM0mw8oezWd7+5PTm9WaQzYtcwlIPFtb3Ab3Pnm8/ztgwUA7amWi5+r+bSxv/iyvNmq
HNnYTeTPbja73mKh4o3HfJxYNgm+YP91DXIBkpcJnBjYfoOv82xSsBWC5iNJ3rwR6I6Kj2IhB98t
bE0hpgtnGLt24eqxedhqJ4y+yubVWlwXrcZE8xS04XuGRm656rGoHrIynQVWxVlKZqRNRIuDD5gs
fd3zGh5FFfZ5KDX5C+WBVj02ayA9le52RIyodetJHZ+hvGM8G+AUVdJTjato3pDb/6BljCo/A3vv
0/t6Nz4gt4RKRA8wAP0B2MDRVUmo87i+SRyNoCy8n9N7pt8sbBlNe0Ws1UDwM28wPWCZNeAApuNd
bXFYUXOKljqX6kJDGIsgo+UqA34D0g3lC9tr6GDE2xGGpLR0xi2WPf0qXU0fUxQ4LMbOA4gv/qsz
kjXyNMn0xJA7CT2/E9W5f35IN/zNATU1aRyx7rqFnYRsnFWqE66w5rhYzAAaL2ak66DOMs/Is5CW
gagSqvCRnEjT90xFLC0z+HtQgEctyi9Q8E8sKVph++VFLXiho73p8LUAiIZS6rHJDugwAoWbIWcK
IsMtza0w0QzJqpHGEXsfxoAXmr3C+T1Mjsw8QFTuCkOhbKDJxK+hZ8e4eQa/R2gh0pZb2IbGj7wl
6BxrMgemUwD6M830Nao/CW+uPWY57CcEbFNWH26FdsOpONnX7jEbWuXVt7a8s6zBD6iN1v5ezoYf
OCH93zXy0/HLqxbO74GJmFewvps1pDVQ6p0Swrnb0LAmNbGj9iChET9Yrp/jRuf4dRTgNLCUCK+K
p3npo4tcjJTBv/voCwHDQtJFhkBFXPK4kMBpjfrSGcKT0oh9KpF/vrh1UNZo2kvvbsL+5h62QSYF
s2BLEYow6RYJNVb9xnHqAdeL1PX6sJzEEIibeLH8ogw1rEuVYCn4WpBh+5+kcIIWEJ+hmqkBzkYf
RJHWc72J02T2Mx1forB/hYdDHbSEhwWgaWmFPzcmqIqjXSuxws9SPCZglRvspksn/i4Eqp9ehOEI
Ux0omyiyN0UoHKVkW9zRezGCChpHoEwYmTOm+rsJHeY030ck/FQVoMExMZLxOVEHhXMc1NqYbYHL
WmRt5o0IyRVnuMIoWM7SEsQVmFweiam0qNd5ObURSv0iYo8q0a4JlUhGyR1AqNe6Dw5GZL0j/KXt
ALiGgG+b956pk6dVwg261xeLVLu2Ooqa27PJyhDUfncOGR9vCU4R0p39XWMLT7RttnZDHjm0NA8E
C61wKvOOZXN733ZwZ54hJ0XHYxT3mNmcGtMNMKSFpsW4Pl3KzgRF7iKBd5A79GbLs6RKcZ840uTi
+wZQed9Vzf3d9Ud115ud83Fs/S9L6jODEqzKmDTa6mrgjnki/HvBlgyPdad40CAJEsXOwWdfVZbt
6KHMcW76SnCcx+lkCU1rOpvO4colNyD3Z/NY8584c+Edx+T8g63YRxO3avwSL4xas5CG9stVuZ95
GpwnRmatEDI7rM1E3NXOEidRWz4MA46FfHu/lfDC6+EeKmAFD5gA4+byHAdIrAmbcZ5dGqfpbEko
xtsyZVsH2E12xsA7EZvu8gdq1CxiP39n8MHixE/RabhA5d+V0vZYTibwWFVUpAuLPOVDAShppL6k
KMh/SmopVcxYzQEqD3MinC6otNTh6ktYQfx03oI7WTRqHDkGuGvqNuynkQsCg4j6dR0T7bZKZPVE
9iAgCG+ehoBwRx/zGyMJWRMI1bvCe1GuqdBUHLp/vP4zUgbLVAaxBs5Qs5gHwrhibsujwprHaVDp
+8aJ2eiX9yHuy6McY6g96Ew6axYfoPYICbSbNp86k0ZXGh+nqm3ntq/QVqBdBBuRWjXrTPao9IuV
F4REr1mJoN3WegnGRhneqIq8MHsey+vr6wobXz87LjGjamNkYECkFYubGn9SX0CleBPRT6hl7QXG
gpVor8t2gjbuIiqDV6vMga1dS65uUyt2TomGdHGDzzsnlp0NTuILBo+cjSHPrjjFXrIzGzp/WyVm
4T2koA7vH8lbmc7PenfbiwNcimiOBNvudm1VuZIYvmMqmn61gKlb7mjwqtTTtwGomBNfNdBRxigU
nE+dNU5mAobCaPEQ4g7AS+amJdweCyuI86/WeHUmz2HRZvcewQMarhUIy5Sn4EpdSrarzEZXGh9V
fBslsKXZOoMJdyV3poTkqsOYVrzJ2o7v0tlaXzWn0pYHqRyIvR46uvVORiItwf+kTJZI5JVzr40j
q+V0VIPvzEKB6cC7cMfE1ruWdGFtZ2CxxMumfb62G7n1owEWnllrU86raZG1rl7/5kC0w7J5pzhC
+uv/4epZFC3f7vlV/d/XJ50pREVBZWpWoIQO/T/PfdU2eIrFsNfyc/laWDkxgbfnQDXbDxOwUYff
8QcorTPLz5xCDNSjSysyPdasbh0Mva00rLWxa5qmVirjp0KJZmKwHVo9gMDc3e0z5h2lhQ6sT69B
XHyEDpj+T0JAIieM2lX2XBFa0hR+fw4TCgmzfFGP6WcJAsmQRiW0ReG08z/1IAffk3NTROHb38qa
6Ugclge4SlVFO0ECX8JHMbmPQKKWmgoguFOYdfuHIqcWt3gqZ/oHS/ABEtcfNmrcKZnkMC/9rSq3
6gIHCeXxMidqWUxJ+0ZTe/WXHJlv+/g9qC9HEgW4G6MfDFQ0nGFg7Q2TpxVuSgIej1ULlk1U7tSC
YEYX/H7bZTBEMDx8y7Szfjl5fB4bQdKzN044NiNho2T8hahjr8ryn8scfLEXwi3Wqv6TBrVv3mCy
aRuKf2ZPagVRrBVuVzuBeD1BziyXkc0jjmWNFydbNLtxU49blxEK+g3S24Ag2hlFp9783BX6hO/Y
eoYosRDHZAsAmBqq/lCXZUAJ59lqLZ5czi6PGMggYQQ66Cy+bh2GrlKdBapl5x+FFXUlmzGY5DZB
b8dCkOm8uOofb1r/i5gnp1neQrHwklCUR5aVN4goWm7kXwxiNq8/XoxZYLm8JKJqVEtJ1OjHNjRO
1YGuZa4kSww4DMoOfPIj39A19kRPFnDsYw3GgtlQ7FoQn3v0T0b2I98d00UWXFr+CkQi59Pbgdvn
32BQleFKv8ua8Wz2VmQaS3XNARzazpPN00NZHdkdzwEiRKejAnAKlGZ69jjwh/dHTO2N0hzFNJ/5
pyGhnRhLXWDv7jZC+WqDSrrz9nVMBnP5avViL+4IqXYHfF/GyqW4ummR6WqtQlA8o48MnHQAOS59
Q11NrjD8gQgrlzVEtTxZc7QsI7nN8XdODtQFQKBYMe1PJSyoxk79q+vULdnZn4qqyZdbLxEPegDN
1WoaBuaQ8HFuiPVGlExchkV84M9YSJQGiwqvoXlVXVN+hofQYkgD0d/WvdItfTMG+EeMHZyaTOui
Hxv0CA5sYEvX9Y4kOPu8W6ivRpBm31yGgMCCF3zTdUa9jCAfR4cRbJA6/shBI2ryguqQDCQYE4hS
rUXNj4rDmUCFIW+XC3HLX7N9qdMWVY1FuG5o/JwrMjna7E4fLayIwwJhuwPlNP8rP++jd0COc8cR
0Q/sjwSmf10taTLvelB42+B0kq31dX2pg8cJ00IwklKJ/GkO/Il8/DXmzKbYDtn89jzw1sZJ9gkQ
dj4jytEp51OUnvzV8ekEbNs1jx3ARfVcwk7QKTs9UGF5PVu29NKWwq3di+lX4AF96CKxa5m622Ky
c1+Har4F+tIZL1L6tqDkdaoXwym/B/qzSdAU2uCVWcRqT+KTo2k0MFPJOlAJoVSGuSDaez+psqoQ
/iGp/tmWFAdkGQl4D8J6AIxLJ5vzsdz5xFoGTcq6dOn0LzxR9tKFV37FTt749vJgxN5QehK+Vr9j
yf044dZ17k194qJ878N/A1r8H5aNxIots84WMPt1OTjQHW6eeFP3+ey79T3kcmrbV7swzH5Ls+24
zvhYXM5ySP0W5Itv3/Of+PpvRstuT93r1xJfc4Xm8m7h+Wcg/uSyBQDo6sqg6yidaWlxmn+meCaz
0S4YvyeXjYFtLRk/KNk3nBx94F3BKCaL2kqJaOnBt2Y1XDXcI6SxydWBM7kX1F0jKFP9fiIISm+Y
/hQFd0Xxvt7ne7plZ19Z6gTJj9M+mTdd0rQ7cBUAE3pkyqk8YYbdLlkQkiRIENb6nDFF2/JNqMd8
Sswfy4CmCrr8hJS2kpUvHjAnCeac5ImU6yiQ6oXyc09qtWRYX3CQ1fZ4P7wfoNfszVzCQdw7VVuI
Dl6oQzSgVPgKjNr5KGElMqBp2/Yxfu8x3G5bT5Lm5LAm/Kk8YEXm41NynKgqd5Xpduo4hME2A9+z
lCL48sqd2O1gaOdrNP88geoH/ppFe1dmVei8bfR/7evYYPcMKp68uC9mUjFivBedyGl1SfurIE7+
/PfeqbDM0pWIHRHp/usyHDfingKvOClLkUr6unMoHLmZJGKVHHsEMF3o+ExTcWX20he1HeUCAsIM
F6r8B5iqstVkh42gBKDqo2XIcIhzUhHRy7xGQL80nJJWmxdSD5wkb3ixMQnFnL0ezZDK+2MMZzUa
6QhcTlHdp1Qq576i3rAuhAdE0dh/HnbplpxOB+bkrgtqE9Gr3Vci9jJyUNgco269HGB2ecn2vSXR
LeElJpj6yQ/4aAC1tdyKXTmp/SZBgPdr8g7AkhdNB7NEN49nqZeoD3D6vKng47SPsEDkjkHMZyHi
kgcu3OwVOyYv93LdC5SC7oA6dRh58CZj6YtMqFgGpNjvgxtBpFYnzZ3NCDGap7zuHU6/t6YqVzNS
ONoAhg9qO5keU5xkDTpabUb7oKWvX+gXvBT5RHMxxkJirw7RfJoEodkPHbxWDFaKNQmxV6WDMHtE
qoV0k6HRxNH9LOfisXHqcC0Mc9ZWQyJJAIeLLOx9HQ2C+adeSw1iihW5OaaIb1uZiSpiUrP7Z7Ze
dxP2e6vidyNhS6VNAt6yYd5qovhUErwwUur8FZXjoxqApB0MSt+qj72ztARkllbWrVN6flV9FK96
WsDBeLoWZ+hlwmAEZ2gbGieQZWGXi6RJY0O5h16pP0ZEwdJkJoIrgaU5P8zEefL2Ku58iAZRHwJ+
QcXOvHRfrSE7FTJWqhSsHfKw6yGbvM4wxIdQcJsxTOLDa7pWRdbs37o4doAORFNZjYFT89GP8c1M
3Je+mKBctiBVkepS3uqVA8jMtpuW8YY1B0fyVO+jNcXtgkuCzX9gknK18mRBRpXkJlNzMDW09UiL
X4vR6hzmDqlT9putJxQred9PJgKThkZwbfgYxUb2INxx4hpgQghln4w9UTvsjHiQv9gVwuYM3Idn
RARWZE6GOuSVd/rveylNw8NjfOk85oOlTgIXlqNesS8rH0aa3qnEIV6HvqemezyOlYYo0AUMEe/G
JrzoZO33yUGq37damiP1cjC0ZcO+Hv+zd49MTlCJu3j4RbHie8oUHfVfFolNq+siYAInLQmVSOj4
EfIdB5f+nZt8nj2B/vwe9be7SKRgEBsO0+ITwAKwgdA88hcA+RWVX3ZiZBCn8rcbsAb624efjrzx
awu0+OizBFJyLVY+oSPUe+gaYpf2uVMoB7ZeGgixtlTx0PLJHU9fIEz3URy9wTONmtDEFsgFqhfX
kS1FxTmaufRBMzuySUO/SvuNfTQDnkHVgVbbwJ8heDnUNmjhtSK8PVTq0DWW1gZ2tKNb3vxv0cvG
KGBJXAAQNathxgXxXe1rIIeJhaXWTM18Y7uKiSLXTMlyk0e56Wbkhl5FBHSGtAOA5CJGCZX392IB
jHlDvG5VMePlivmcVJFzBP9RtBJLbxonLWfSIGXx2xPUNZsfGmgB/kpw3YrymrvuwW8E7AsIUDsE
Sq94zaFWh0+4iyS1LcthacHs1A8fZg0hbIpUxRkYRghMKPj0Da1j/vsLef4mqvOsy2qRuZMKBs8V
CXRUKb4wU9gxoJSKpgoOCGJ+08ngRwCdR4COIj1LN6UQA/KGhYQI5Py/5bfsVi1mYjgA60jzg/e3
FvfoDCcgMRJbh6tKiPCoJ4e6DiQxeizc0dhzbx1EKKC0EvGh0+AXwQVGuklVxXnfbc5qWRNfhH9K
A8H14Pk/nhUgobupN7GaJuJLLV7i7QgLPM1PtJ+h+bR07O6xFYyCN9hsDyJI2TXD4M5rE9IAHkQ0
Vuxgnsv65F0VnaOyKoVPy0gNbAC8pXq9X6DJJg+s4lFk1O+up3cJNc9DGLKQax7oWYL+EiuVakK2
kJn8BJPcJ8ebxPQMiuajFBTQe52Xm5bwSPmI/sREcgQ1uvfFlB0CW57/ep+neD1j2O8jdgu6TgKo
W3JKrSssW5fnoysO5AZdM3GPTcsScFAOT9RhMuI2cNlHvM2fReIdjX1Gu7buJHKjY0EFhq7Tkw6W
lbmXWq7/aqA+jiJnKrODnS42mO829ATbVqWKVhw1ka1smVbraDWZ6urL5CZMDCYDceFUAVJPmEpW
F15/YuLA2424OmJZRgUKPL2xoPZbDcRp2Ey9De261fMkrhDfml/FD5xdE+wGzPeFSc65npYHuDAl
KRnBzHJyoId+ISE+uWeuuDOB0T+XUbeEh61/WMHPNgN13cQc+cojTl/UJAhMqxolas2xMIpM6zSQ
LZu0lAQAg9w5qaqHIdGFMFfDjztQY2D8pTy23Qgn6+aiGJg8yOHPymiko8H2FHOEXDliLSwRR60j
pDeqA2W7g7jSO2FLkxggtC8esZuKSsCSXK1NztZS3mRt0XHFdJhRnWXN8BM6zs7a/n1MyXpx5yM7
OXtS5llS3Q9Si7uqOqjaUcxNHeU3fIo7IKWGR/8iQwhO/5Rn9Zi1tb+/jt1VFO+RgKCbED3VTh6T
gtGwHhEXnTfg+2RxMe2zp0R8VfxUVK+janz2Ca9ge8sJQ5fFrwD8WGyLdISdOthpl80ZzWcq77qw
o3zJ+uOgR+w27O07vCHaohNEGcT3xGexrLocj5omB0RefUdJX0PK0TBpdm1x+ym5PJqHdEVEPkIJ
fXGpo2B8opLq90EcjpKUpFAsKUIe1ovjOjdqn4IY0ZpbyxtWkpjxxpTy3jXO+eN7ktKV5okN+N4O
PlEUGUHtE0Ne2/j3mGWKa8WdbOi1iwp0BESfQKHg3hSRJFHCyvuwdBJcfE3uFFTDlM9qAj0S0JDh
UawP7X3fMFHiZnv+yi7Q/C0lvqm2emhy58b+1HSIJjmNCVtHO2o/hyZrUXGyKBY+429VyjhIN6L+
0jOby7t59HyvYxo9drJWcdI+iIIu4aF19yyWV6jMkdilHHzixMcRMy1neMN95R4GPlVmhEHYmtJy
lwg2OMYInN6BzJj7JUQKiMZeB7XSeeWDzTC7NmY29uGyCZQKwHeKJ5SBsA1qVu327/6YqCZmrkjv
t2Q/pe1VI5JVMJIXjuvT5RZsxZEw0Yve1AA59rJefLKDk+hJaWUPyhNDsPgXEuoincJyVHbZXu5O
ZGvAJOgdYyxeXO+fSmxCxnCsOmzO1wRGYwBv3cSXfQsO1czgOmiGuuJc/59GNJRBmKOXX1VMlpyg
KaLAJ+30HzRh6vSJv2FrGyQ1KQIFb3q5qjbgn3QcI90EpJHmtRk2hlxDfFIuarF7VXX6in12cMBZ
z/iOQ9OFWlgr4fvD8JS+WBYWCkjL2Rs4s7oqOqU51sXoI0gEWTzEOE262rNBJ8h98IL8TpzKM+N6
tFE4VTPfmDpPRMjBzlIGp1t2oLV+atF3HvmD42pA2+t+plUpLfFNi2GsrnUzcO4clMiUDnF3mBP0
ap7NSb8GJxVKphPG88BR+Ah1OVosxgR7wc7iQV1/VZUyVenkg/o9qys1Edo6zJNQ0OvquJ1Jhg/Y
JLHoz/9VU3XoPjdxT/uTDHvuPAMaLrt5qpPdkZpPpjeTD3x+AVDQtB65+ddhTfVpcs+fs7saanNq
I3Mtw9G6k02uDKZc3AUolx7ja2K4RtXaJnSROwTRgHFXdwc8JBRBSYMpPAPV0NQ990YmDu2BOCCl
OlfZ/opeNshfLwQBLc/rnC+44XLUGoiNW63vqQpsyxrRaqozqpIYf83EUepNGh9EEYm/b5/5rBGk
LVHiMWtAQm8UEGLDwo8UnriMasL72QjQzhazmcjMqBgvlKixbVNZq5NDr6P/PG2SD6M8V5L/X84C
q+e2g1vW/p/Dtd+3whTJJ45xa6ONPR0gRN6gtSta8sX+S1hzzPx1EOgGpEDK4kAWzBmwdpgcUPgj
J3HB6if1hA+XU6fPb0pp95p06m5WRMbxxHv1iaHHBwwI65MIJvTbeUK3D4vEePwzD0nynoIqwdhn
z73d9v4xAJDxM6LT/QroUEHZbmcjmfyQdRdrcCcTLZo5EQtFsEcDOh2x2fFgSuFJWLdRWrrL+Mka
RTYqMnM90VFUkyRR2I+FmpC2RGiJcBSLGcYOzAcSgR7NkmWodD2nZyZL481DPt6ByN3GZ9t2Yyqj
IZ/w0/CUjyD9Uzrq1JHybd4kWd+X6YzoS6UP7PseSjduR3T9neLPIO5AGmsohtVHr5XvY/HwFe66
D95++Ppl0lwuOSjkgHJONxmcWU3UgC/5ncdX6kVoRdDtCxaC/ILfqYzXGj8u3VYoA+gxWMvndg4A
U6dIL/VnPDRgG2r0SyOD4lne5bh4ccGJk1MhJleB7XV8Hj1IptfcvQiQ0+cgYFKW8ezr0jdPDjSR
mODELoKoo4Se/8Y/ntqkns5Xq7LX53gXMSiu+hKNWVc6bpHAtJ//rvDmjUvEx+GRdEcUkWkNJUoX
z4QK6BvOkfro8GXr/bgXa5VuyRzGvAyANrbeGFw8JL+iukGtHKA/WzJWiIhYepEwOjD2ClBs0IV5
4SzEe6rDWHK6aSCZZuOYcJpPc+pg5CTKqR3KqlLbWzw+z+NxiMzVH61hZSDsV84cRysb1D9b9p09
vIB/JdAac87Kfu7vNeR1RfOPejOKXOqfLfDw0OWBn4q33PiyiFMZfRK2IPMEx1xXYduBngsPCPAq
+CppOmPx6jD+7khgs72Rq2+WxgvCegB1niD/wEQjwoKRS8qYe8mBgJ0AEejltIQeOxOibCKm4O3I
oTiBjMkCsEqEU3vKqNC6N5gyRjqdjzoRHDMRuGBj139yr+JSHOPyeAR5z5LR1+Sd6MbwtvG3t/qD
DO/AfRClwAm4yurXonyV2Lvoqp5kIub2TqsGZWRh78kuni72rtQQFABPrsphfbOUvTsoYqaDhs+o
N124kEsG+wWAu6ryNjogYDV1NwnpRV/gcU9LFFI7tsIOV3R8SwO3Es4Xj6Wexer1vUtE/U+SDRxV
WEXh4v3w729cgL65WCFkwc7QI3S57JqlNKMWfyVKipQ7LJI+KmVmbD30TxpBozImZuGeQBOIKAfb
4eL4fSTYHAaD69TqdwwiVn/teuGIplGNZSZHp1WAtr4wSTmR1OCqQzq5r81MLOC/MOQWp/J3NWPf
ICMrGFVUD415rZUe7hQVTxkUO3ZLZ0BhuoHfeYIumXMNQVw2zIcN83HJIcJB2+Tkt46ahKniWBaA
EIVgWBuqFTg0hGEYU1cMnI2mxcjZZwdduirfQc5qBMY3ZUMZ8mt+HcyvdUVHyV2trj7jjXfG1X20
dxQi0hyfEElzdzYCyW3pg/EMnrVYEHZRg87DthddJ0ID1ywN5ScoQZTsBijVovEHPif943pO7vXc
hHe3yxGJ4m/0EHtR1BmdqtNZa+wK2Ab0Hm5Lv7VFlZXXM+E+2dSBDspxxwti901QVJ/yijbl1+hM
G/ZZhibl4iAzs2jc+XQxZTUqwJEbNckM3WKWNJNBNXQ+PujV5la0dJUxzd0MktWgQbe1LKqyxU/N
2+SJSJOueauRkSkrDt+QWg+O7IpcbxDxMFs4pR8eXgr/8Oa7bgQTP0aEPaSD49COdIsaLvn/rHW+
M3hByXRdoCcHcKlbEmcs0LfxtkGBpk4qd/w1BeX6PhdVJJyqqmZnPoMLn9Ze6Tf7MhBUWXCvRbuM
7ucjm39VH0WqTByXTotTX8d321kohtng5hsC+u4WA7gSsa8vHTTquFnV1rjgNEzK805IBgcAdca8
DkIvjhAIJG0Qsz6qodovSkWeXvFdynv4cYk/Lj0ULjiUMIrDXpMDg7YhhdnCqqrEKPbg6Th3ymQH
Ets/RsoMu9Iu+0qTjUUroCjuAX9rmQwEyxadCE7xjKig5/jpJnqfnMJ+jSgA0DlFyrgladh59hpR
Xa/1WAjCLG7igoy/cI2WZIt2TOPlR8BzMY9VStMocO03Xt/79TjZnsuC6zAQ5hoqSvTwUj3PLEwG
WjpRfTH1inYiN4GhA4IYFVHPclwI5zP47HjMyQ+OWkRxfX17B9lM0zsPht5AFcQU2pfySPQ82H9W
baVBTRDrD8OWw5ZRaCs+f1CzWrntp/j7GG9eUkIYS6P+v8w4/Y57wEpH1dYEHlufS5QtLLOAsJEK
dccGmK3xvROKEgkAEb3mMaIS2HdEv5DWZbw5ub4z2XzO2DMxQJ2XCecs37vpE80hCrWsP+FlJlPd
8lbzReLpNRP85eqUGOWx13YJNNufKOc6ztWkD9aWEnu8MAVrgO85SgatbQR6t/VkWFM0vWzPhSGr
JPgOaQLNHEvl3I+jXmPIlmy0N3A6rBlDPgY/RUcPy5drlBaI9uMLID4HkRL4f/1Df4yyKpfVpwSf
W+zEb0thxU81ccqFDGLWgEI1xsnXqwnzOb310+eZwifAnc7i50Lhmy439M8Va8aYxaNnVFZlBhJ8
wPI3jFOkC8o7oS9SGxz7TZ4Ac+b+hG/ymVx1JIIQBZ4lw3iDJ8YZa5kkRy7Xv7plY1if2EVlpBwI
WQjP2KB4IDgz9lf0E/b7uVyvs6j+XDHVugNyxhdOC2xbbvpGteQL/GVPQFUGUKskzCFefLg+kyXh
9W56dsc6tl/owhLjxbMUjE+nqAuPKMCnIyouRlliY3ElyRioqTRakRwS17ljyIpSf9CEL3tQSPFe
v59ZX+V+CjATTCeW4v2X50MJhVLXihdY1amJuJjFSzrM6mtQe3P1I9ECLk7tLaqt8gYvyL5vP4Ph
vHv74zOC3Y20Nsr5jVSQfWXfLbNco74EIVMa6azbVXFuCIfZeXh17Kk4gdHhQfFkwEl4FmyriLMc
AAsSQg0N/bw/7cUCDQzVhVgwL3nYAJAldWjAN7Mtr/Nvxirtkkt1VEzP8NEeP24o+wEuVZKnVG8k
Mn1hi4blcsDi4fjxKQwmDd6l1elr3gC94nsbc71GSpAk9CsCY849orMfi8JH2G/HY8jTAvYLYdbY
8eML8kDdftU1PTvBnjwVcG4hrP+opEp175ve/QiOK7bfe8T+c+EoHXxx+NW1NIPOPDZSkJ+azxwt
NNB6fc45qVS30bAWlit38Xp2h71UQ7qemBeWPMkbJHP1RZXGepAlvqbXJ0XT5/Bwo+dmQfBtt0Lp
3tbo61cNolimfqU1ukFdftdxjePfc6TBtF0eTqzGQiASOkf8kpWY8B4A7dtjPiNb91XTFmvmWUqg
4QBCUauLSa6qeiDeJ1uyXkCIUZIgsoIxJCbhzOeZbNSULn+1NKmGn9KmvX+EcKvOZTMhIX+XIGnh
+5j6qsl/AWICsb+/0+5cr108SDkN4soFio6NJ8Id8PAuKf+iEpDpVay4XRd4I4NJxovZH2Fi3jTO
jr39h22qB2DFdcT/0tuDP/Xk0j73qaAI+Ev5xdZ6jDQTNLrKft4eCJwb/ODeX1BXXMkoxK/PFYi5
8UP5x9+kJ+017n01LmawVITJaQN2g/EC0vo/7kb7OrHLvms98w6lcHSy7zUeaALeXmpqX1rJ+ivq
Gixgy2dnaLasCaqLS9Ws9qRDqn6gdKwFFgbz3IWLtBcRx4eQAalN/1lPdkyM3XGSdiZlX8TPpjbh
ohY+O8Se3GbWJzEgjWyCq72JOed2Qoa7eGYfhN6ICW/N5CgIV3IpEQAM61/CIdGfCBzl5VmnmSnl
gjsgRvj00K7GWv7GhtbY+u8q+FbE7nPtJ60D0i6eSoeo7wvPkcvUFqBMvu13i/koNNa0Ij3xZHbX
ITxcJLLmhv0ei0u/gWFEgeFFrVCW1xRvc3oTFo6GAUnNX27UWJ4zkuxjK1Ou8/7RnLRXcXxWFWBV
ZLuRJpSEqmRmCENBTrPH/YhJGm0xUoN8e6q1GBSwV44jj1P1b69gGEYvM+KN3pZfY+2FlWCZqIVA
nMJ3IEpEHaO/canY9Thz4V/R6wWMalX6Mq8sX6Ge38vQC2mobOzhcsjP+5XLNE0kkeXvCxc0UQk9
rpy2NpD9xzoYDN3qnajyP5Zxq+gL9htANLJBTGLqKy7PJsVcukIJzzYKwnatAOb27X+YAiyQJ3fG
FCAMI1VsuCCyAXhU4L7lQbISJ7Iqw0FJhqMbMcQYCTmVjw800fRCof1mEi2YponeOvQxqOLEQCAl
c+aMb2cb9+cV+IHZnbcfvOO3sF/8gCTYk22O2nNYBh81TKlgGEyd0dbdfFb+a2J06ruVIKlEGdul
805riIbQ8USLpr2w+BqV4BOGe3oBUNKVdYr9JyYH/vvmPxuUyqs8GyVHQYKwxtb7CiWECZ/zeY/8
q7rDQ2RnHQUlpr6bQDp4UAOlxIqehD/N14E6l9+gm6wOPoZERRE7NJnMwEyaD7T99L03SEDW9N/v
Ll0D58fAPxY6pVKN9FLKix3elEwPNtTrebFoW5vW4I9+YjPHFT4+neNXZWUj9VqiKf0Up2GhUlkD
t8NiAlC3Xo9KGrG+vmv9foCCcnoYtUVZE/lTMxSs5dhYW80saGH5UYr3LELWjg3srg9BqZkwcuN1
8VEgj9V+x7vfTTP4HqMJ1I1zzVZWVyXdNshLh4qsYMsX5JNBuYIDA6IpFCqFO1PF5Z5xN3ltj74s
a8iJ+N+N5UV3nQMsK+lbobfl1nZInCgZIBpg5mGW9c7iQjzyJPNTXMUOaICWBtwVKSwzhG5t+11i
SwafwdaxzBwkAWSAHfhqnuDvLD1IxlQiVmKDrLnupNv2nKgzCbDUKscTD8PrJ0yvRjmNnT21oCJr
JbXHtTnXGeacj+dCQrTMHQdDrICSsDPM5Pv5KyvzQNQvsEQGdr662GXgaEQTuwkB/KM+DcsXo7ZO
+P55Ub38ELd6PNzxQK5ZnfwI14qG8hI0fGnhkPxOi6Xf4rk8cQ/lpxhQfJJGfdxw29AdTaWo+Cua
S3gWgEeIdMw2JNJ+Elg7Xip3wVNvbe92J/y5o3iB9MiE+cO5ufxfDrpKa3jSB/bS8f7M4YfeXMlE
m6wOPxgw28BK7lWudQBeuH+0QIw45xgLHTKHiUSgEOa3Bb5OZtuQvr/T/vSseXW+cjZMSCmhEa+V
pUMKN4HW/Nh49JXx+wy+5sLv2GAEYen9vlv/MOGmjg0OcVk5UI6PoGHKWp58pDGHSj5Gas0GI4La
U8KKuS9r/Rf8YLA2X2+RhnNtrZYRbuYmxMo5WLQzzF6p37efAZc6GwGwPh8Cl7kQFOn+zxL2+Jog
tNkBGIv1wIleoty/vOMaTTiYiSCCpGXGuZK+ROfKRegvZTUGZ6BVRgIc2CQ/q716648sjBzltFlH
28h+zg1BxRYgwq990y7kGcMkq16erhUOtvSxy2TDasnHIi1UfST6wLxSJobYxm8syV6iPkOyRGRH
U1/TLoY6erwDIlKx+j85GpEaSecpLEgbvFt2vw/8RQNwuJxGxXTWnmEcF/Bdq2eUu6dH4ElngXBK
yI9UbKJ1mQ1HoIe5sM7QwkSdO0hUJC/TWl9CJsDUYGD53C8DwgE3Iid0jqUHWtnWgSRB72gyroBP
lr9GgeKhgy1drmhIdP2wyVGjNtu/g7hqXC+F2O1KhsXy40s/08rw4SiQ1M4IVRF92Zghh/vAV3hn
DLtaJbie68kr+gapDQ9x/N7U80F7evB/MpVbK2emGQ4pDtMPPN6tyzrOmU74O0S/KeJJg4IslTdl
fDuFz3WDGy1SehbXVXK2KxkI21qJXMYl5viTyohRGnx61VU5mEmgs/4ipDxvH4ajenTvciXZRYwG
xjM84uRT2XKeeTLB2FzZ8TgKVbligqcpxNRbnSqjal6V8yc0a0yo1BwVxEh2Lf34g6OQzk8B5DsS
UIuyL7isPP8YdAqZ+ua1TcBs8GWZrWdiw6h7ZDq5XTQX7svp2mgHXYgxmR/zCUXXjz5Wt+aZ5aqm
6UTovEVojvdGGC4cm/dPEKM4UN70sP8IU8h4CUf+Y9/YfkWxRmDk0TE8zRhQnO8PeEVPJXBEmvfs
3l3LpEoLw64nYw0czQEN0mAe77sDaDx0brINnI63mus/0iE5V0GqIqLdFaXUUEMlRGu4SO+TqR0K
PyHyVEeNnbzBwse+QyzlTQZ8nVqdJKO2tqOCQRCVZaaKKgnw6Cxq6RP+6bMvdmpI3l8nY3IJuQ3b
VZh9z1Q53ltVXw3udmefEi0mBAwvqpMaEYIpof8uBQa/9v+2+ES4Dq9of12e7Sw7RgABd09ZgzIr
2OVCWYez8JKovvsUibTPHsFuZYFOqVX3Zihou8DTpbcLGg22TNaqiGaEjhoL+Eh5FIDF1yCcwoyK
rrcP9oeEs9I4Z1TGwwn2Hg8e3Oe/a7Q0HuY3Yh//xCsxIkhfHT0KuBC0DD5OdYB7bToTFDpYzIGg
5tzDziqbu8mYRludnKt93voHq+Qc4jNiwF/ex78/qtGklBcugS3q902KRogPl3j7+0E42b6ryEOJ
8/hDdKt0xn84oVmtbqerhgM0roa5GxhBLZciK3fMehmu4l6PPtBxi7vTG6Z4OcRHqTMm6RWRQB9b
pOuGAbxZVkjOSMJrxbUEn6vBe1/n+pJ3v5SunClmoJKylCJM83Jp/zJaNKFKpG2LyA7e4vj+3Lrc
q1qWRv0oVBYyMmXK8Rgi+SGdZdMrecfWxFhxAtyt7r1vnLUDTyg+9s3BgxdA0LnhVzAeBAx0KX2E
x02IQQYaSodgVrsy/qwe2+7pwuuAyu6OUou78OzR8Sniq3jx1axjOWlcAXikybJV84DCtz4b0ygl
glJ6+T59iwIwv8L5q9onMdJVvVyk4AGgtw4HqXFCdZyigw2nTRhk3zLsCQEoWq+hBQmYWBh4qg5A
Mq4o6ouAwThcV98nrH82ZULjry6/yxl3ep24qXQ4fio18QlKSiaI8OSoHVa97dbW/SPIgnU6Zdkp
wjTCyHAjlfxwJ1mITfgG0ab1h6gYVSXjVVDRDthHio3DlbnubPgN5Pgtk8gzf2ngA0tGreQI980Y
MmJ72aJk+meGaVs7bcNn2kqBTUijgHZLUo53EbWR9g2jjo4Y//K0VGlRBFND5fEIfP5xOe90aMOW
GtG0cw+r+leTP8asGotBOWsAu/+j1nBh1Hq0G8BTqC2crzzwHryDjIY5mvbjlQp7tOIRYUJEznFX
geqJ441ZIkPz+dZ3WXG6izt56SStUSnMuNg3nfUs4EMgTdB1kojvJDGKiKKe5YKaG/+5G+5y3q1d
BRo81kJ4LPQl3nAMo42CiCtaC/4Hc57mU5/p3V2Igcqutl5JuP5+kB1fqmHa4itisYomyVeNCiaT
ic8RWcl4DymI0hoYoOKzs3qIWXYPrMnXdQxuptgWj/iR0ma5ofE3b5KVjbfM8oa2X8/ct0wZiFvI
nnXYlpkr3ynh80wtInPPZPg6dCJRyDTga/yOpJTaJ+yL0kzchVxXFrUX6itgaq1ohaC3ZwQSWRRq
zqHLfIFWozcCp8gEE90oinySI9ti6roAkRdED9mZSnKcH9lmx4s12qE8leB8trBYJjDWxc3AxMMx
hcUDyTa8bGxA6b6jeknNdSv3eq6B1aP1n9a17KG4XLN9zfa1RTKrS92izghK0S11EDkEK1EO40G3
+Xard7/4zFjTzFVbT7b7IBbezsqmY5X8KlXQjH7hUUrTsDBY/LbqqzWHTOP2mKm8CJtTonQJGWl8
GTd5XeE1288AWcwTv+gjdPVh6dxvV/idzi5+eXNh8yB3x0ecZcXKvTk5ZJgIFugaKWrY3SHE7i/L
1MIarFZPSS8bGHg70gqHyY0OfBUaJiKKbReZY4RSTcvxrCbhD0sH0ggFn/Mc4AYWMwEI62smShJ6
8fzeO+LeuJ1siZ7BA+ZMZCZeB57g3yRpiNbsgpUOwXWGpfVtnZ4lSiFsesBf7sjDjte3KRB723+S
SLzKpTfUced7KBw3pKL+/VNkLwr3z1hfgGr/zB5AUREvI4tXA37AbBEExSndxmspM1kKrGER9oIZ
OZyhE2rkvRdDbk9/VrQl57be7FZ9YcKMvq0kbpKLIRXe34rSzOTNFkWGOaqaBiljBq2/ShgArHzF
GjWVyp54GAoTCNGaHt31Cp320YnBZPBXb2jPXbuarmIOw6yr770yeaYUbUwDsI59IzBxhcKXq62d
FXbqyqTxzefRGfCZUHSDVf1KDM97WBWy5yWeFtvNwrdGv0jQi68ypVcZknJSmemmZhc3DlEE+wI+
GvyQvkO3tHmTm+KCryqc3odtEHzDxkwdHfBGMb/Bv+T8n5BBnmKVV/DBGNpe+vfAuZolNA1e1XcH
L/aCL5iB0vmAILrqhj+YOyIQv+3gZ90ZJLwgd1tc6MDafxWHRfwr49XW8GkrYo5diD6ZrWPXNT6d
0Alzs0v0YUJM+mLEYJijOYhCC5xTI3cqQh3bgLyTjveSD4jsDdoNyEhCxdRfAaWgPl3nIzCVaeac
bNNnAG1piObHfRe55Zatd4zMjLFntbQyvAJF5Ln/2P9Rg7GlXpg9eyebatq5qWq4e8JlThISJn5m
a9BnFYWU8bLbU/UR+gjDVb/9gIhqY1JB6439P6T5zMUTdKX5DSAQPNuIjhSxHNA4w0fryGe+sQFL
lmNYW7TX26MqmFB2K1k0KUNFnv0bXHb7nF9kf3kxA/BchAdeVBLxuocAIpXTnCX//qTNXZjEgfSi
wKlIETUxGs6q2Z6bVOIRmPWwXLGHWv5kjfdFhUKrB/MoEWAN8KpaQzCaR7pcJ+DOFF8tzACmHlPO
LjLM5yZzvftvwhDL8Kkev1n04/zdyjwDH9D9vnVsukwChwHJ391jrtCUs0TWP4dRF9ZcvtwCkboO
aP2lpWACPk5UkJ+9NJ1SakBZdM3iyZdTrCb64ujOqpKdi7tWOYRzI4umGP5iNuwi1OTdAysukx3M
fZUX7ZY19WfMsIbY3I7U/P3Iv39cOFHAQoVkQ8d70C9P0hhzYyJBT0YNyRbrGQQ3OsLzIaFfHHvb
duDkA5h1chkVoDNeVM14VEAfNPI6xkbc7+Mt1wuKP6M5WS02RIDJSpucwWRhvEqeraXhHPAaHgkT
wdoy0ZqdNsjS2Lcoi7I0nW0kc2HcAb8dmGx+Q0lSUTCg+aeESxV4Q1UD2XDiXeW+M0BhFlTvkDNi
JGwalcS6I7wbCuvRB2RYFCs18oWXEaOS4GS+67lLFDmNcqcBDl3MOtr3VATt7/QZlaYzRyupWhpz
InkQ5Oza/GMSyJRDGOeXF8CA0VeqvJlgsjZkMWbTahkoK536pgOiDhWTBoBXRPO8PwTHsf2KMPhe
/p5208a4AakFYUs4IxDJ1ZKTHFemE1ubbJO7Nz3aims8HUINiM/tab//cQ78hNevSAQUl9G88qjb
RHK3fd7gSoQTJao6/RM7WL6ie/kNcYPMcDwF/oF89zkfI80ucdFNvoU7v9IJK2mvFoU1OC8odOUN
GE01NtQAmacL6PqOPiSBebrAMbOpSMCUMQNTlImtqdqsm9olK5baqXyglcY1BUmkkBevSU4kTTqn
0dLreNwsZzD4kzAcKk4dongBHQGzHCawXjbWu1a8g3OCiSn6HR8CrzWMF8MHNzUjCUZ97nfeSGDg
4nCKNpNINTORmnggopCsc5CUGHK6AT/CC1V0TNkBWFff7sBKf6s/ut7NLNwL3Np4SzTEQjlirtba
GGsDZgYyIU3ogrWcuK/uYb0zqeQ4FYTcxg4B6CWhgBfqLwntxwnZgD7DKsZIHGcvQSeZRcEMP6jx
UW3bcXptz/ChH4fXpHnXNlSVfwGdVvyoRA8h3l9q/PNUpVIF0KuB8/BsFcGx4bAQDuBcuSHVnL6H
10u9lxUBfZCe6b4BHwYqAPMkBGktb01Apcmovf9m6AoEfGX5EC6HY7PcCEJUpokgxGUB/o6UMjmJ
Q5CIAmFJgBeC27FxIWDcRS1CdyDhRWWaKfeDdLV+FLS3eXLJ2ZMPKj0hCs+RUty3xGWw6aYmq4Cb
HbPenxg43FEEYwSngamUlxlAtlCj+8F1ZSa/03BsVvUZYhfykGxR6aM/5JkuUC8BYfPLGCMtOZ2I
5SUpqo+ktrJueIcajMU4XduJI+bVd6SbSxqduPNIYEqJlzVkWhmklCeF4WT0H8Ym6/kKl61bUXKh
yWPr7XRwHOgATRHsAhztrddFuUUypcAhuJdyqpH/MAbwpojVuoXo5u6Sw14zySX+GM9ML3okIBqX
jfpTFsQyhdDXoWHs96WNUv7NltRWSJMHcIBUSUkmIMdNQdHHq/e1QLWRuxjt7fd3sRtLQ/j6Ew1X
Yw+VtkULro6RAIk9tqDEBmtDwOoqlRxiGqcoWqRyFzd70IvwqpT3KJ7GDWIKWz4nNjz3W0LT++bK
GdNFLlPIL7+H06kJ6yweJiFHVnNRCDR2F5FgDRQLemXuS00ZUBkqXhpePfXtxjdXDvp4cKjZq5Oo
zRi8/ZYvK4rFJ92FzDPtkfxH00ZapjO5gGjwNYRdfa8BPD0M1BdI39e2Qif8HK6Y75XQI6SyhpQ0
iIVYP0+770dJT9DtE5KizAEwFyN+D+dcNjtCZvQ38dujl+iXX0iXalKAc+mDqIzhLQO7x6eE/5B5
s3gZ+Sf0xm35BpcYsCfZEVzrp2oU1m8UoCiGRjSCeEt1rRhg/6KdtX8wq7PGxzDxvAonGy7GNAsG
maT0qKk8pcuC8IJjdsYKxAd+y4YfMl50T5QqGpHUb3MQl+PyVMJcUYbnAcUXS/99IvaUa3Gy35HC
hQOa6mmthoiBbAHQqEWK+tRT1i7UjvcBvoDFzSRLatkCZ0Vd6JlI+AMwQO+RJZuqhBZuvMBEZmYb
Zx9KBOBmnJeYsaqvmsJ7xXfg90E2mBXjhWGz6SXvRr7Nw1e3iGvdUTcLpgkqqNScofSmW6hlFers
KKUx+aNyNQe2iSvfxPCLViEKKGymk6inGP0VJbLRpUzJJveD2MqeV2jkjoJv9JvlZZrRRczDPv/T
LgLcGohf76LK8HS/CSnq2RbtA1lCggy3e5ShfEpErQZYpCJb1dE3dz45u8nZBMoWf3Qb9/VTPj02
q+XYdavxtXXE+pAmORhxq/sETtHaw56IiONcAodwchbkbQSpt0tkF3UXxLrTWIqiFl0Hy+lcuyLn
al2tkbVkgc7+pkA5l1MZ8NA0Hb3DTKvr/cRPtL82blnRfdqM4Xyy3warjUzQtvKOm1kDIjJ/jMnh
S3nz+NoV8Cp8QqSaiK0RqvcEZCBxBndXPqos55OfBtTdspyl5tWTpYGtpIOh7n+41CyD/41M796i
P6LZz7g+Y07GOGsj2UhkrSP9ALFn1+naew9WTyrHWbROTf+cnUAzS05L/wEMVgiH5EwjyUsDxH5s
nN2CI7aTl1mTMeDH1NPJedWNjE7Kq4p3biQ3PDGnf4iXDsiMOCLnECN69Vcp19Sjyhu8+ap/qkNc
Ef0YFwy5WZYW4UiNU5N8ad91nJDJXI0nT6oFxDnSRJgcjR+MEG2kGKYeJ2oBk3KFwtcFVexCnzMC
O1c3G2uOgsp+gEb5Etz3cHxV/5n0Uh3zvieOlylmenMOauqNJmcfjegnBTU+A1fXIupn/OKHydGQ
/d5WWALNS+NTaTCGchfXtUOJfsUbdS9Mm+rnqv2IpJAxuB6RPE2e0n6FO+oTjiA1TiGhcJ6C8fn5
FYlRxjASFacgOx5VcmKhDh2Igj/Bei57KIzfNfj6kO109w18G03m2u5vZ+z1WdzmSh5PvgOaakXQ
etxwoFMg0q0J/CXVFcQarjhRLfSre7qDWTw8vGLl+Zv0oGEJtbthgQa0bJDnuvBgV3OsYqDlSq7a
5F3hMQ4zYinhc8x/bf3jHg+q9YvTRp+qhpeDlXMSPUYedkOFujOywgD7M6XjCTUygxAheY3rJNrO
cAFxpMBpTJTJq+zVta4VWC9afcfEb6hq1ImBtoPBWKNRg2c57o/kMyvZ2bkItj+2Rxo+/AyJjCAh
jnpbDZ2dL5yrgIjc+qplLmeemGulPcyip0L6GdLv5ISeUTSNLa6GrG+M04Rb2Oli8TAUuyR2hIkb
WA4e9zXk0semEypS5EPD7vNSnz4gauja4nm8z2SUovH+dmYvCDdgMvzowhgNdKgv74TvygD1ukZV
c7dKM8SKUbRxiihVO91U0dbarn2h/9wJOty60cQhC2INA/sDJtn8xdtyB8axgRHjHHRc9pcD0RTD
tAVq20a7ox15LGyjcqua3+PsRBPUpyEZhon8p1ZheMgsYFskxS4B7FvhEB4QBrL2Vv4CI9TVtXkZ
YGSCk+g5uwDEBFIBz7ri8TMYmUAH4MU+d0emzQtEAJe+IF1OtkJI1a6ioWhVtFpDFSu6wsGiuIbA
B+TALqKK94fTItNQOlaUAOXz2o2RIpgc6Oaul5FtthYHfSggU9KAHOw+VyFS4wwHOwhXUyUpgkwf
Q7GhLccw0Q2PxwU3IQlcJJH5/HoVnEmnb28gf61/g8qfKo838IpfuBnWopk4ppOI1JnM4toEON6d
i2ldC7dOCi5eUNtU2Q0FQII1y3rwhig1v/u8WW+7gYP/TrL2igJJ+P8Xg6UeopaTmj9cJyDq1Ty7
f3gSorSz1isx3OHteuJ844uLwiFSHyiu1Xh86/90HHVWC4/bdBQvtCy6lwDSaAal9FUAsT4T1V0z
AOkRI1/JH0fKoOPW3sXkxquC2Qnl9AwxE1leuiipD2dCBrnVnVG8zaLtwxRB6iqv9wIXuK17PBsz
1K9G+Abl7lvcyUF8Zy5mhebw9DJA3Pmp4cQME0S7dg5IHv8NWhPh8rKxBqyY5fGKaHw/m8O37Y3G
y85oz5V3fjAZKPZohwyPTsJF9QYdRXU43tKdp+W/e8fLiAFjPNo0hg+8Yo0SXmuTNK/zVR7NmHXN
kM5spm1qp+h9XUNxBQsowwvf7IjVoRzXz3+8zNsW3QUDRCWsVXZeeTTma3o07kFfUfuIPdNgwPnQ
Bg4yf565P3xTRgWbv32DQI/mgk+t7vVv1+pP/VTkElrcOpUnzhNTpBqrRiOBA3D3ztKRfZ2Exa2T
UVaRKfZmscW8aPoDWYfQhgGHQCMfAJOR4FiOwMzNOgSrSJCRQYeUX/EHaz5I8LpjVCKtPlHDgfdN
BL7jJPdIy6AkLgcgMBL0i+xJFdsSoGIPaNq1WGY0UPeAi/fgOEhLDqM+HjRbXjSrB0EyIXSJfid5
UJnwY59ZrB89yeOEtgxNsm0lnEx5nxnB2hUjJYIacESmJzVvEnRNn77b+3wz+ydBEsmmsTk+Smip
T/C1dOvu0IMXeBFruY+LhfZwMoOjGXpBRor7zpE/j4g6e3gDMzUnOOmSlMp0F4hE4jhm5UB8Hn1M
1IUY8zJszSpkdwMhwBFJwpMB4OwGzGuFXtN+oEIdR1LWgmE9gOhqaLc+bYSnXFbO8jjzqO4/zhV/
LFJf+zHiR3sWIHZXlnokdZaXFnZr/dTbKAoei5PC1+Wnd3BR+QCcdpxfVKdg3s4L/JqG4pZXrZj+
L/LVWnsICkNGmAOuh9ginQDnQFkJKtGlgbsHekRJ2ySbbHRLSXrNP6CDPO4OS32OYNRqe8o4e0R2
fpjdVK3WVvLumNjKK1c0kOI6fB89HunDfbc3xvbnXX5QUSmUVny3k4uD+uwZVdNik+qzf1THk+S+
4GWB2tzM5kLXUpSt/eBmkcMGVyCBw2W/bmYto9CzP2Mnn++l+LJMJnI9972G1udvRCLzWPRVUkPx
1f0pm+v+GBm2tkr/qy8+rKQ4U+KWnELZfeThYoqyuAUsS/ZSa1+zoz/fim4r7Xoe9XHQQKX7aybn
SdNE/bYYM/YP+0cKiX/miqLhrvgvuwVgQvcxis64rrJKdMEb68O7tL5xY6lXIAb5ez2v/Y7asdpy
JHWU40nHfdPy16D+UGLeZVhjxVxq2n/9Bm6bLYLb6KWVbSjzb58gAPe8BjuiyoQOn4vTf57DNMu9
nOZubGHhVFOda0AAKAfVEaeJd0iaboj1ORMw+bTVwb4ltl6wPhaAraLUxUw7OCTlkm2OZef8F6zb
Mh1upV3/Gfz0fJ1SPRf3/hvFo1iiz1YThIydM5eZxyTfx/GhqJ2KyDUA0sUup7HTcIYb4LxeQ7fo
9e4FQVypUI257shJ0IkUiSO04cGI/BcfAwM8TKg2BsgUVOFH5yM5mBEg5qkCkQVEd/vx8/L2BCV8
CEzKToicWWwY2mxzvOZvcfmqyip/cxnIR2jH4Ep0/tRJ1dyBmYjyQJEuGtr07MS0oXWEiNAh/kF1
7d6TJr/A4bNXtjM6PkQ0jnrZPwG+npv40SmbQFgtGDqvqWZzUc5h/z3SGIrC1ov9pVwhR482/wXv
3SNCDBgpoeVftRUlwi0Z4OsfcgkI7rW6LReJZisIItWOgFWOP5xFyNVlInBwKijHEZlwd/MHYFHm
ZP4imJMNDKtcP2MjQT6MJsWM/cIHfoJGUZ7TD81Bm9Mhgop9ji9nZKjvAs+IbDWrsf6TxWTPVxbM
/p+viiXgmMEnqQOnlr31HTTAMnCSOX+EpRjMhAlqfWkqqMe7MjZc2PQ9pmfOQOGMTSZD/BflMqZ4
Yag0GQG9l/36z7viE38x2Z2Q9I809DzzE7rAv52Sux3dnSXBRPmqwoMe2cYsYn25TzOY0zJauoq0
ouOzr6YjlwCJhzEi0udV62Au5VM/issWuN460NYNn28TE1zBjkaHDCNciONn1M0ydpJes9qhTTXV
OvS81oacRXTprvkz8IwqN1KjkF80MBnGUMlP+SuVEiwsHeCBM8pEGgHMmjze4ehLuzkZf50RibG0
q/Z3CeltDtwBZUpRITV99O+bzpOwmgXhzOs1iXYFg0B/yNg3T33tGRPo19b9+nJRldh6FZvNz32n
c8apnrKNi3Dlsdd2k2gqbcjnxUrptmmhEteVFHzdByyR5ww8XoZkUuCypcy37VIStiyk14+6+2M0
1SLbrgEZ06uW9XN2I2//qzSEWvkotESH/l2H+V52gYLhuXshv4UrnAJEnbzdfbzuBjfTnurVBv7T
L0IWOjQA3PVeZzJXz2FMNNmJ1r2WT1nZkpDyWtqCMWfWgSBsgeVj+fZyQ4CGJ43BL8JWGXxQyMkp
Pxh417vSqFWoEUCeZVAUhzYqoGkB7OdUej0TOxv3g84bGv4PoBD+RowYmD5xlKgR+D2T0Z5pcCl4
wuFIUo4gn2cOOTJxPkGFNCtzXdgkRkJJSN2B2M3j/IVCvFAinTg3ML0GNyYlpvGmEuwFvfd1vqGX
CxIqjFFrAIcqqqxUdigCgYx+2tscy3mcdnP1YRxj2X7aTLFf6BDS0JqeLNylEXBhWV9zZa4MstLW
P0JBch7MvEN1zZHcuV3yfER8ZBsZycPQHUZb6krP6TYQZGLH1pJ8SDO9NlMrCOXy49Y9uLFf7yRp
I10XHCPBj2ZGXN6bKLDo6Lk82A8pQD3D1V4SATFlUVH38LQGpHJI8CvxAh0VsAiEvwWF7J8lw4wr
vR6IlfOm6k2rOmJyjShoGKRQgLcP3uzVdyeOgZs4H2KwXSjpe6vTRpO+q+QC58S9VRU6t7Xaq4gr
RGuPeY8Uw/6ijgrIOlUG2v/ZlmqtyVkNERlRqWPeyvHdfjYbZiYbFM9VPSGpU16VqX9yuVBYCySa
Mu2Nh+CSfK7jyzNAo4Cqcds9aGyXiHvFnkjVm02Mu+1ocKYjKDUDav/fGEZPj/+nleNxV5fP5Q27
+ypi01oBAHSQz5CvnCoTEKWnga8/FdBEUut4k1F/2BVawsgRlDmHw2ttd3yV1CIdJ4pbccLfaXZ1
rbAOqYYsINVTdtI41IN7INQ11XCe5k8P/AFLDYDLPnzKw8qBqzOGCjdsNTBn6fLPANa+4EEDu6xX
bJLHUfsnjIFNY5A7pnRdmmIPRfZCB0k3t6LRArxJOsJ6Z4qORY0Rko03rYr9WmlyDtRmEED8NXTC
Uq9zLK7pt7SqqYEKZVX/7hbf7riuexVAlBVQ0PhGkx45wQJ7pQbW/yyeoSp+G3qSwt2VgLmkY2Tc
hspeQU7hJWDM1+TvlozUgF1TwX+uzQpOr1AWoCrq9oRQx7+Ol59IqZjSYMKYLxc7wiDmiyIqHIwX
oX/mJyHI3s34JGd2xumLwhEraufCbGzAtTX0IOEvaXoodIIlmX5ZvqJrIes8iIa1ePmUtxjWjhVV
FQrg7MAMQMV21H5SdPUofrFcMNd9A/CItnu7ayL63aOp6Zfs3GQushBJPgZa8VFIjEJS9TO3zhnf
bglrte8syAsK9vBZMZAKaALzcSYaYnOgReGLX8BNT7leLHucqTIUbTXnKak8on9po074gEnmNHlP
F0goHWlD5J//DkPW1S49Xja/JkFPAb5P7rQiDu54q1kEAYsNOb4Fun/zlHy49CsaXcT74Fljz7la
k9zZSelEH7pGtwbg9Upa0456ofDasRkG9Mpca72NnHq2+FOh8SR1ieiDzM/P+ONIf+vRviRePJre
XiHaO1e7+/ciQQL9ugoDWpZik9fVVlmN2fNYlGLTFbKM5upbZ+1GUkroOXOJ/+ARN49g/yLUnrpj
GjZFOiHMeF5KYvXxDl4gvaohjOmXP3A5wiDio3hTnPdLoetNDNd7phbWcaaxGpLkGIrQN31TS3u+
is4ggpKBMLdZTDiT/mHDIy/HrTwFVqK9qlHshkw/H0oMHhEElS4/B9ZeEDTAtzogvpD5Pgrj0NGS
HE4J7mMUggcJ5PE0aLcn6W6pw/oE17Ga4ybivuSKv+VXYIoToYOYkzeVbkhibSqiw/ln715uyP2R
xd9zSqRHnJW+BXfVihAVImcjBTMYg/DjSyKlcRzdq/YUg27doGfKSGcgIot7+QibY9sStm5HrCAx
YLymcKgU9pc4q6YSBOAGmUYhN3wDyfxxzjlr5oppNqXmiw8QmGALzrA5dPIeZeghRXcnGrszigrw
+hII9iFOz6kbMxvZWzzNG12LrTASMRKsdDyqkWga7Jt4nSKWNwjHuHbxFULwKtCnH/nCnl+pN7LU
CeC6vU3C7fqcUCn28cqKb0flBLGrRqUi2adhTW1CHbBWxSpRuxEO7wRc4nq1vkfkt7hgKshSTCHR
TDrNN77VZ/UbctWcyV/a8TDZIIIj9SFQ5cT1FcuKG3WETp+nKDEZy2mlin6fcjmu38q5ca8AKBER
Kj8ug/eY1Ds5RlsczxdpOFheyyuaa9LLoG3qHD8TpKVY8sMiHkArhmD3LVvcDMPSGMMK6YcUfDE/
cRUpLmqk7y++i/PTY991h5eYEhKo4bGTHdAvXAY0xY7my0CSVsDv3YLVmfon4kxex3UVHxTD8keY
k0K7wPjehJXad05Fp4JRWdxzjLdcVggB0KDJe3BlFbvQZkYUd75h8sGGJk5d7BoLKhcz+tp95M/G
JM9OfBTIxv4l2WOFo0ASc4u9uC1Ojcp5SJorjY9WpYE3Q8WgxP3+RKT4wFYLJHjnJsQT6d99Tiht
8n/KWSbEqw1mS3G+rkcOqbYXaeWqi7hNa9PTBK7byjaWIr5BHdYlRwBxt8BtCa6bZo58x9f6I93p
tMoyR7St0ZyrDD4WsbmmkytESeaoLpbDj6fOEagOtQqZpjNYihKULiAeFU3j5YsiUteUyMyyO3BK
uR/JhrS+m/m+4solSvFmKV4/UCK0Sl66IbKqO0RouAdJQ1z4xs7pmJhaWA/3Qv+EQCACK6hDGduh
omVb4VaM375VLTlBYeDPAyJsBeXc6VFtMKl1gVzLpNbBMom4fOsFUKZ5t4A00VcA4vMDd07llbXO
gKWHClYLjIxvdMfqilxUH260AFoMAwo3zccL5Xh/4CuyH9Sxy9TXwVapUkond8J8ZjCj718VqqF3
2jqFSgk3anMCtNA3KC9NIDlQc13Yg2jNHqdKH+Z+JUg9cT0VKuUvClSz+AADh3YdSFO5PaEVRhHA
L8x5bOIx7BxrOKH8ZWy+CR0v/9wWnUXnFGQKJAHTPSLXWXD6m1unRygNabMO+r6yJyPb/iuLtC1Y
sHQePAgeoFHwisLshGwzq4mh3xHxYUTm1epHXkXzbwCVtVGxPmQJk/XqvOtXwJzHZRAJzsIMF43B
szMJa5A91OrBBhptxRvYqeYyyWdkHXU/iYlmucPc9F2L41qlRYMOt4it4ukcHkQZYBc88AtReEGq
S3Pd88HWZVB/oPliwi9Jb9xRCOdurBfCOaOmEIKyRPZdKkc9UWRCvd8VSNmppWRF/i548tR0rg68
HlVQ3Dxa9wNkSmMp106DK4k06qSzvAd5XPWfSHcOH+N3/DVPvYjNWPWsCYrKKr5Z7Rj63Tjseyp2
RH10a+o2imvLzR7GT0pW24HM4kYgyiHdLgHk8xVzNLxFQIPLte2FrrAWp6ufmxTV34B6GCmOIgjA
5TQrfZq7uwdSDJw1PiP0s61SG3y4OtEQPyb7LCXyneNsENTqy2cCQ6mWBFH6mEWaVdd9gl17x6or
PQybWeMyOMQV6aHn5jLupM2JCWufvIHt5G/+trngX0mTSFl6PRvDUzSmwFgD3PHsnM4kmb5cHjnw
MFlUTOU3wXV5dQH9qVlPuquGlc3X9HC7iRZqJqDpKkFzL3sS6BKkNWm1BqVs05+3Kg6PBepNA/u4
UPNnp1PBetp4wfA9nEWxd8f7xYUvAlDbuci6u/lSqj7gEiSXSZsyFP+pVLmCfdki85wT6vbLvjko
v7OL6lkzkdIQ/lUIU0XZ07HX7CrsawlywZMbx5j57uXYS91ovFcu5MibW/eOuRURlwH3zXmdA4DE
+3WKpUKnEK8HOOZDKvpNF0wagfCOOxCkmIdPJqOOaIC2XTOKbUzwqLAxOHRdILUamqQ9pzXrqJPD
etJWg2UnYlutltULJD41gHss14Cf2QnoYg+gmI17yWfU8O6cLGxWI7bxZ4H6rtk91GfT4UR89E3k
WvlclfqrDszvgY5ZLQrvTjxvRZrs2N5ur0zAD+j+G4btonk4lhnfXZzZKslTLxa/Mql45X9TqjmZ
8uwRZ6/8ljWHuEdtjBYgyIg0PXRZImQzCkhvp2e/NVcIg+3J1IcjxMKuGHPNSeiSZkEVsZaziKFZ
3lKaVHt82EYrfZk4mY0nqwywY3bthBtHCOJp9y2ealS4z7ddlwOZo/sJ6KSorQLYNDO8gT3F561v
gYo03kQAMkJP4vt4tZ1nVnZPiYbJn/GEw/bPAgGV2dNW+4NmW8E9TTAdXsuFQgnm6pnN9ORSMLlw
Fwr8GTgtPxo4bk623Uwv/7emWgCJ2jUC78pdsT8Ar5qd2Gfz/CCteYVRYA7AppQgGNzgdg43gMW8
92TlP9yibus/ncs0JaeH6/FVaKF6/T1u0inP4O7KUXZ4UZUfYXc2Gv2bcI833hv1X2/dnU9z8ade
Rt817K0Z/XciyYWcAStuQhf+lQIZQeoMzX2hw1QAVpecJdBB3KlaOyt+P0j3qmixWmzY5pMyBZvG
Q04qwUUE//RZWSq9DcBt5bw6EFNaK45VATUUkjxU5thWNyLlr5G/ce9lWgfDw8dYGBEYHZ8NIwWG
8yNwKZ/Ptq9/EW9hLtmGPqQKwLKTnxhBE4u2zmYw1F3erLjRL1vW22a0eeAEvcn2VT5OuDWepJFy
9JCiPbqKVJpN2xECC2Yxzt6NGuixj9ljoYfXYvJ4GD/OpiHYNRGpxsZP+FPJmScuGw024LQyiLQT
ueV1GaJi4/ldJE2dYF+L2TQrrGWB1E7tpgFljIzz6Jw3pJ/tGQ1Hv9E019e16lgF/Rl3n6yb1Fmo
ppVTooFuHTjFzBYJGNYAFjhUL+r9K4f53inFKpxXpy7IrpG7rmJyrSuQV/wpUqxxtVL5tnl8n4Tc
j6DJXyyMnMrM6Zeq+41kz/a5qtLZ1ybDzeG0uMy3emNaHxQ+d7zZ4qLvX6FU+f8Scp2Z4Cr7lmVO
0v8a77C0AckHvlCP88NFTitspEO+lKz3I9TiWogtDZbAYhQt1tBKMJDy6WJl1YaZ+2eomCnSqJnV
iZB+Um/TqTna2OJmHRlcdmUkIOR/wsJMWcKLV1+u4r0dfry3UA1y2C+SCGrXZirAmfQOrKjc9V+o
xvYX6SDsvJNUd9IRZ3c9bw0zsERIvHmfTp6w1GcifV+d7VACafGZ3iuKp3uSDr9DGjd+Cteh72tS
Zq445ZSE17Jbf+xQ/NrQuKi/Vl+Rh2RQgIL6qDN4HShLC1iT6sM9gHgqyY7tbHpXJRLvUxERcs4p
1RVxHY6yE27noKxHgHLo1nMrPn3iebV4x3w1YBk8PhngzYxSP9qXRqxWWJsTTIuVVIEbKU1Wun4w
trYSh2PgW7ZZowOBBvJJgoeR5+mU5sm3GABpe+WJIfhDbyGryrBeGwIxX88JT4e3/E1CHi+9lB3b
+ExWoxJvfyz6Ho82dVTFZssuw4CdbYU1Q2Qw6VcN3B48R/QT5XByh/+IPjtZ1bsvj6wLhF4dBTnn
mTMtIifq/Xwo2TAoAznDQM/DZaqjuKzT0cUmQvZosSN7yQVxR/rwITTfm5XRi58i/bvD5CD8UULh
GhErMt0lYwBSpmKtEI6Nl4eybSFXXJUkzODAsscMVrifXKld7N7MvAZh533gygTvK1XvBzX7F8RM
Bf8hAQS1LRgI04ZQBgFlAVKN5RKUXZramOG/CBQOpgQN+fgUy+jZjhQWEYnbWUCoaC+S9Gt7BbsK
H5kFYtLCdSJLqKRgtihENGuwezhOL2Z2Z6qHH4tnIare6cyNxDavE2OR7gfKBKK17BM4TASKtg33
+7LEb6poQPz23ucrZwDeXb/3T0fMFtkpnCaasT8XfTmni2s14TlCbpV93H+8tOj3p931wuf7O2c8
LyU6wye+FYfkmm6NC/LgSWX8ybk8Jl6HD1HPfMr2aFtmwgh6zqUAuAYtWg39c1raJjoQV/jhe67B
1V3NgvcI+TKgMWdb8GZkogrkAb2DdjQDd2UEGWsgiZWvCg+r6jzvcy8KowYHCAsQ5Zj4MHyycI7y
RggX3i0SmLrh1R0aOEOim6wZrlb5Awj1g6K2uZuYuYDurFyirmn7mDxiybuqoCGrjIFgkeyXxhNc
35ZfsD71otYcs4hDNjA1rpyBMZbwnxVc1nArYyYKDiG7zJmONtQW/ftonRjOSdJYeIKiAJc50z0X
g7n8DDrjR8q+HurO1VFTgmqXy5rr79SMY2ZKU7YN0oIvFn7X0TXrF2xUZ5dpsw19YT3MyBmApxp8
XPgrNoDfcd63GAQuVsd4oprgeijDvwWNe29nhqXuw3xAsbHfFkXTTmCfuwM5kNOCR+P02J46nVgo
DjcYy6QroWzlueh3cwPdqlr8knagwPizjtBsINIvuwG/KTuHLbvWwwYqVZwKc0x0WlJqEjQFttIw
vHa9vLL/NYpF11CgDmwY10uJgaLrsZJTS6r6jKRWto3jKg8OoQenCClmsfvTkcJEithYVdACFXOW
ukWdHNdbBvha8wFX0WB1RNBbC652DD8m+NpU/OcIWExrcNMrz+u2gLCs+8sWGxrexbc/wvK0gPw+
RsTlm57jBJRo9vYF2L7Z8YJvx+ILD71KjZoO3Yli38a7pTeqtD/f6DYcrVn/dzRNbTa5jMYLRdLf
fuqZ7l04Zebbv/xo4e/BMm637rZC8/CMpQ+22j3fYMhy6lIke22C1g5AW2hWRiABi3Ndkbiji9FD
30oZc4DxAL4OzMCapzXuU5KHNmD2fs7khz/3roze+mKsXYuARcHXdZqPMN1JoHFOjVmLroHR/zyL
c1q8r+qEkSd9FQP+dQibD6EvEiIAEW5fQx+tV+57xSXGNVtsvU3KtL08rgVu6AVMA+Q/RLvEale/
KIKybm/chNpSaaHU1Uq/Lauox2w3y5zU0vZ42LHo0LPx8YD+3WaNtpLyFDedluqBBHA5fWdyJiZr
yK6dLzbz6wooU0uEaHyTSjsQu0j06GeJWu9e7zBnZyDKomYnFMTRfEYhCp5/1rw/BjQQdCQhc+/M
PgPyR8bApizyYFZgJP45r7UpTPx0nAORVGs+KEMoHRFhX9XoTx6GrgIpntfARmhnMBwFc1cbHmCX
9I2ujBYb+XkbdYwjRJr4KuDVRyELVZgCSZRh/uoGTatcJKV/Xe8OLvHwI8SVjay4vUweMVqPhVfQ
G0UQFjc73S6KjUibTSKhtYK21vkil+OxlhD56n5cfpx+DiiSHLvMT0cpdKV9hBbfb0jpkBXBBVJz
3J8qousPTx4tOTalPuDjEwe2sa7efajesw379pEO5NMEJLI8NSTBB3pmVKvSIXQ5VGEq4O/NtMDs
jmdLKYC2gFTqfyoGsLMuREhgo2neISgC96Yp3MWmKMHa0NxgEcGaA7wjuAFcIRs7OO/b158R2Hyx
Ue/vjODPS7Xzdjdo0HkUc12OhoeBE1PBLPyslg1TrxD2Ghb0wi7twGQ1ipteIS7DP3bgZ39hb3X4
B7r/1bLq8aluNxBmdY3PqPDeBNDyA0kZ3u6O3oEcgBZ1GuXqkd3kTLQzgEgtpSei1zA4OFuMTDhT
+5hOFrW6+p2uIWJUmw+suXL35xNhJcRITnR7S9sxjch1+l3XrPrBZuy3BrB/mBozmsl9kMuV22y8
7jGQNzrq0c91Y5s5Br5R1Bw+tyx1SV94wwEMAyRrFh/ffnFOG6NLDtdp3F32srTSQCjRd92JGHdn
6pGc/9Jn3mLpiN/MxpFb0A+nnMif/atbkLIfBCS3UCcNEDkqipbvNTbAuhx9I00eexYV1IeOEUQ7
RcajdqJbGYcA5WaqAiKQinHSqXiBa967BFHC1peFw2K0mWN9uImDi5NO+t3XT48uXxubb2In5txZ
Lzd/gtZ1fDjJ51hDYEguktrN1iDtUbv5d7ZmymEVXlyYqtvW6x5is9MEtaL6LPZkCQKn+QAJm59A
7crpznyPkYPHTDvCmjOEK0PaqdanUJGi/NCrq2eavQRmlw0sqhbT60yMNRpWtEJCCqN1VWVWqecf
twPJ2lIiZrw3G5/haoD5b5t4rq29aruRh12twOsesbISZATdOKUFcYlqH3gRw6Xxjvm8C1XGbGRc
PFk35kugo1RsxkhhcczuUb9UtUv61qsuXcaZLtQpZs58iMuKt+pHC0ks1yCXABsbmrxdahKD4HFs
BcF39OgqSYG7hiGrzQ9KUSuCfpJgfyaiwgVmud7zePubwmwCH4Sbo4mf6+I+Lu96gQFpnRopfAur
uVUkfUXCPC6XVVWvYBmQILoeNOg2T0DZRc44Vfthg2G8F4YNo6foU8i3UiLU1cKz9nz8piDsJIfs
6WDylc3yUa2NkUaZtUx+XEcuIh3EMW09APNWSjb1RqMNp9/f3QtCiQ5SNwOYBxiIRkakMa9p5iwz
ivkBD60He34HK9rZTMAYvzh/Hz7229mVidqJhRIA2BamBJY6luSds9PuNNzVk3uJNsSGhtuMH+uz
hzid5K14ywh/zHAnRX64u5BmWA1UNmPxR0buqyqzL4qLUIjoBgK8yARjsYS4tP70PV7n7nxFG69S
SuJCooGkGJkiWOikFTPw6sGMSKsllvBSsCF5HkF3yJ9IJAanojUnE2hIulTkhv1QCmXbHQWncPb0
r0EObGPEPt6V9uc81xY087Q7IoMbAWKsgfwkOFX+sFKJuwaO97gbEN5MYGJ8Pj1dMYaw3HhwR5l3
O8SqpL6d0tM2kPxQ6eyJ26Ohst2dybb1Iv3MFmH84tG++iU1zd3pxN0UUWVOfJZewlk2HAq+kleS
qKhDVWBARq9DxheSkA6n5tOe8qCM8zdaa6JZEyDYIaiYRr9t4vzUIl7iI0Ot575+GsVHUoLz8nCH
vUkiEqr7w1Uiy21gsQDnea1lqXmxtAy2he/6YDxYO48X8EeOQnHM0o70sDZ0Vx9Mbc7AXRsL1yV9
fSEcCpCnxEQ7NT5l6P6VREhaN8q8uZwSeg8fKG2RRSFH0qxJ0RotiR4OLPz8M8FBo9ypTJgP/3YJ
NLJ0PzvxEA0/krzwHyAA5gXSjP6CRf7tHujS52+yj9OC2APzTlXxo44hCMSA8GHPjZVhLhv7UDgQ
4tmvP+b61lhbGUS/5Bykm5VkPISKEYnVwZPi2BAu0TX/bu7u5NXT1q7YP8HK0oMxCrNcC8lKcmrj
z4s5XFh0i0b9m6DEO5IHDnlvcB7xTokwFJJcgnAWUTkPCMtXv7vOZi9hzDSOwfruyaGy+vHuUnRr
ulwB/Tn1ZPnODJTQg4eWTe4JQb3CtORtISHpGkvERLMAAw6ArQD5GMmvIEp6R2l3u9iFMH410N1b
Ys+hSfyO60JmZPADNXsRu+7sHb9TehqvajIieZernB9p1UtZbRN3RrIOv+NmVJwMe8YoHFwN1iMz
LlnkCLcRYNG3LqnpqLrwCjHuWNECrhzRtLtuG0PynwHuACHs/gmeBPYTWDTOPldkFXBUJJpqYlq9
ZKeqa0yg8DLU5wLHDHHLYnWqaajdpu17QVZNC4ek/XpoXG1caxHqJZmNRpLJvFWyzZHbDsICMG6L
O7CMmaqOLYAGMwJlLAIKb/N5Va+C2RYF0Y5Gzkw/aTQYN9oMe848rv6cThVuWTrhM2ONxo4VmYEH
f3wHVIAZ1xHGqV/ojQiVEwvr6RwgetgrAl9hzBH/aX4vfI8wu4PcEzMPVF8JjcgNzuOa/T8tDVKe
5DLXZRRkb0wsgwFY4HRtfos8PrZfCd6nlX1R1yqgQTeYUJ+XKwFYRmnLdvBMkPjmNoSiJ2p1DnoT
4wP3PDcAcQhB8mnT/nhtonLQD8sO+1a2BVMDntKvw74FyLDllyHQYAyAEMQ+ycgXLRSlifb4BM+/
9N1RT9iMQZU7nzMudZ641rUrMO17qvdmQgNxNllg8vRiqnRyn2WBHYmsz3i0lVzmEYwZH+x6ndUJ
I4P8d3A1gykw1GkBrVPRJhq+G2VOMeJ7lPq5nh/sXKb9xLaywUWDuj6ojN1xd0iJ+ki9nZWFHcoq
+6etrOm+wPVVzcqImX+hVWPe2sIDXmbccca5KGJaeWj0nk+7HZsMzpOcDlwOxVcBaRWtp+fc/w76
c4UcKvJkBNFp4s/mvZ16mh3IaEqkui1ipm3jouET4LuQz/u/9SS318eiAyPNXvpWbfqqDfzQYg6h
UdbKaNBS3Gs91OeEtEXnujWFGcW37j1CRA9P/KIZ46JlCCTocBSvfpPWh/fQuPdj7GAtnVli9r2V
fVAWfx7Xo9dGvA7fJcECiEYFLh8DekSHihoNqh6NKdWW/bYWRvZQuoDJatNvs7pFRFbEIxmalfq/
O8xXzOxtn0/MhSJoaAyXbcDXYeEC1Vf9E2VM3qaoES1+/tBVYcoa6tse1kkvmmWkD5corP38gl2x
sX2S/f7mzpLDIrgEpn1pxvef1ZPS/w/+qlx3WIw7ZJSoR7yARJ5QmG+4cqPuvEsCMYh4ZQgGQLDI
yJ66q2B0A/M0x4ArpVG5/GdySuVhGNBEh2JHi80UI2tIpRvXe4Ywapg9bq35jCVEbT6iur+AzjEN
omjR9SllkKJSLsNMGU5fGZUJQciDtT5Fc0MvK2P2dbJQqCc5fVh/xxCcExNl9YByDNmjXIwXtddL
hVZwD4uyELColqOMXe93sSjXkx6kmpajmCfbygJYnuFOn17is0ou6XURiCsCZ8FlO1bELappplPM
E2Nj3coi7UpxkDY4Z8be7LFHSUN1DYnaFKTTq8U/0v9d3o+E6CvReBxLhltcI9wLkQm4uS9pU/K+
PVIlir46M9clipLNG44LZ7v13MC7LLvQPRB7ZlX/2h6e8LU2rsGhxSUbC3SmgZUPlWqYVAFQBOiP
XWuo1FcapXMmPr+UJUWj5V6CnaEpxbxI/Lp7piE6PoDEGd8nDU/wYxs+GPXK28Xal4tahBw3/ue5
1vzOAT0SyXJJmpphkgjv1oZT9kDWBT6A5KLVNsUZ+cnsLG8y658rSnrZgWhyXrR2Dh5b54vykoPJ
7z4WuPOYARsAnyFc80+2kBXOHO/7/iuyofUpDPCb7v/5JK1UZgFhLjZZS/Gvm4cs5v/yC4jvmM1F
2y4iOeu4ggNa+27OpaoDpjENqDY64XhxXP/qkexhD2RRgHqdOPTXdVl4eOPJabk/VKHecQDtW2fe
ViWLGYs5j6ef6h93BIC+mq2bFDBpxMfJkyHV9M6fw8eK8GRFJxEB3e5h+5GWPv/VtcyTHwhgF3Wz
2UE2XEffdGgUhY9zoV716TsxDXvhpbvrsmESu3f6ckpirliJpLbX3M2N+A85zjoZesGVoc4WOZtc
9vZjoQ3J/DHxIdZEd4DyyZMiU4M8E4/56ftUtmkX875TkeAKr7CAwoPJ761LvFgHTmZYnN7iYL6s
0byynZhH0MBYxZclCbWO71P/daHm64E1XVW3Dg3lOWe+Q3SYEPYX8bk+RzSCdqHeGzKAQNbxqjW/
ff+aXstk2p7VvC7xKlWLK0Bd/hEuMlnxHHaIxK7zqLoKwI324BP9wnunCT3hR2hKqVSzsmJ0r438
ahGRh1DQ+1gairA3Ni38zevukcSVB3OTDyUnXsYDVgsYGbQunKw2eWhq5si8Aqf5t8o94qd5WYYZ
iwS8mxuRXL/4Wrc6uKbqbpNXZJqfr1RGA1nehO3A01K2nekNY9Hx3+fsQtjOZIOxDSzrIlP1jeZU
Rcm9nl15R1QPTnxSJIKxgc86E/FkwbTPh0gWNjIWLHJRm7VWQVePScs98XmsXRMWbQ7Lzsli/faC
e6ZpZlwtymM/D+W7edT4IW7zYau5Ubv+T75NZBB1QWNKa3qqP0ecOW8Kji/+KSoD8mDwVJZwEqYi
Cvw2s3HUZJjATewq3f4ov3KAMdevGgBotxTkNztdYTZk+DTskgU2LtkO1+eqabyRHZmBJT44h95y
q0BEfyUNF/eihNWyxhTD/0Nee459wa6/DY4dGAqa15U4Z60gVO74AvuUmawlm4R3WtJtlF8Wn4mG
ZxSPyaHZ/GfEOVhcPY1hpmJCkzpEanAJ/dLvqwjjFcJFs6vm33DJz/Lx3Nvgu32uncV2Dt7oP0y9
iAtHblD+6pdVxekOydpa556+05KT7dgb3htSr/0gFnr1ytMgAaoQKMUGGFyuKgkyCEGrjesEOqeK
6GIF0/nZzAdkjygi03MHDSMZuzIz+9uzqk1X2hcojSugvVXjLfL64UFdWtutwnSptaGFL+JErZcP
yNrilzsTn4oRQpKE5Lhd4rdL0QCTc5mTTgMOU/9BHjautEX0xJMPpP/8WLhPgpMvYr9Xy5FrWy1Y
OW/gn5WKodPZ6dUvizeZYfvpCeQozYTX8iRIo8v/4H0jA00cE3xcnFoGknhI5bR80WYJaR/n6Ded
UU4P59nYYAi52mlwcUEKekPvP2gLF/6pqzxQhbYj8pBIaJDftdBpG76S9kcfaOrxi94SCSEoj4Pk
f/46iC6LzvgwqPJyPEFrUid7CuFnQBqZf++GDK+luqLrGfX17Smyo4yHX3j8J62hUt+yOgcDvn9G
CiRMABBKUNlDJzxPMxb9+SIe6xtVxZ0AVtOigqDk/4TbUC4OFwWzkYr1HFGJlK6TDYDab4C0ZuKb
6tJmjy9tNCei5vMlk3+2VRh0HexQZqMBrHYxr0HwfWfwzQwwf+W8X39a0Ju+D1G+NzK70ty7ApIS
2Ge6wNt+iIb1ItfPz5IBVs49WfQBc+atH+qshjp6tI3v7fJ+gFgrn+Wy3du7EC+HWgAgkiMQIMpU
/3HgJeMyO1gred9EsyW8Q5XACIZrBQ/KJHjCK05+98uxh6gUT2mBg8m6HRE0whz7AfV1pz+gOV8M
VWk3by5qmdeSSxqmJMTFgyxIge2EWnoFmgPL37yeIX7jcYePj9DirayqEBS22zDXBgc1UwYENf3m
aTRSBevuQY37GwYxZ+g06jCPvi9z5iS7YGw1PeGojj9MeNnJBEuIf2f6zlgc1FpDH2W/8yWT0vba
2GSyEd1fcFcDzs06MWUJWT/KTv/CP4/cuxl9U/ehpYq6l+k6MTPQS4AODuY2zquIENPLzv8tygix
wBUztEpC/hRXB+PqvffYeYC1Yw7mogH/a+eiH+Y2bmzhdK4F4AwygGUhnghztH2pP+0JiqO9ScVa
PneUeJIBKq7DO11jLTSJERnYnv1rk3pwf7LTI8irXo96g9i18jQrahOsyomxzyNHI5Rr/xACDwsS
31o9darZ6cJ3lAlegHimP6jtirV7s4IM2zl1o/dZHeaPTw6I8FP4uPpIf894OfdRyyXUiqQHdYlR
npqGAiH8ZFvCjWsq0IwczDiILcda2EFjPEhMMenZa5p6z2RGGoVcT4XcBTbPNBVcoICEROyd45vJ
zjDrwXXZnUCMfMtkfgCg66MpEfo96kOqU+4PIycvyfPHPu/xg2jPIkc76dn0OvESItkMV8hWiNmE
1YIzv0NsrhNMwsCvsB1ukxu3jgTa6pxyFdMI0smpjalYqSe+GQrpLASzvAIFDk1FE4a14HbqPHqv
jDyHB0vb8Y6zi+Y6R/6xEXEOR7yleiJ610dalcxhR7jXEzPOEULQYTufaRSJ6GddOfim1S6zB6qr
RB+s+LdugSXyz9GXx7WzxjvQhdmuo8XtF3cryc2mFWdwphA1C7WaxSjlgd/9PofM4AV4kQhVHUyk
NEin+Bzzb+AtltvPNAJW5ITPRGVa0IAkdGahKNtrplKcmEfC3VfAUTAlRv2EafDKVKry6Tp3+bAB
cAt81psLab0Rm0lmCFfBVP6yp4xI9Hd9SCA87LahZqUtcpHbf+pZIeLaqUn/s8BT6htErKMNwBmg
sR1g7daWzo0RlgNvliUSVbQd1+fuhK6i7q+ccUsi9y+qz81k+KPqM4MY0O23mnk639ts7o08pqM3
AkBfB+w76RgQ/vIhTVu8IZpJabiuroBUUsp0F6WfBmU+hXRxtjEB0hmltxeRs4ShVtzUScBFq6mn
cd7H2vzt7emLdNix9c8US8Kvn122ZiaxxnpDT0Ko8CJT96YF2pgG9wKCtQn9ZnJeeIAlfc1BaZuB
L5tLyQoU1tHiouEjyjBDO48dqL501izqK0bYAcJHfXlcRYaC/9qJ5vmBtpjWpf1ifG3Sl5dlpEjd
3mGdvCc8TkJf5tZzWq8EhcZoL6IkxFQLuMnOGy3tCy/iehSxDfFqCuGhEillmuWVSbMtA8bVTD16
32Lsp7QRo9/2RCOnLiugwWNziGdeoBzQECWxXbkp7H8wtpUR9RmMXg/y34wHsorj1O7hk1nZNNZ1
bRM7cz7ukvyeT3Goc/h3f3uetydUr8dUjBurehAauBe6R7Vu4Kqe1nCNRj0jUrnsglhMO4BMQ+22
bnug0neizUDgRQpAQy/CBq17e/zLK1MRZdaiH3OR84nNEKGcV1MubC/ElvNB79og2mKQPsauUfJB
UyLGKCyfiSIAZNysKlefRxdrvFAqDImslwKMtytSfM9KD4frbEm6HvcD2/ONJRQE1k4/2uP83FUr
HKgcYe7MiFB7SbpeGekUWh3f3mkQCdb/C98+lpfuWwWVPSPWvXegyNL+qbyxy5YhBlsqNO80BrdY
mA4u1SLt4EgmbFMMNdOdBEH1Nb1hRkt8RRpXHyyAIVruNa8RDtAXEMybk1SV3Y85ny0+oYwIvao1
N5mI7+2Bg+iGqXimd8f12LXHDcGz6VTxuT3ZBlMoazteLwC/ZG+vVUbXd0lJMO50Xb0oZKbwGmsr
9fGiYltzBIpBjy+rjcsnBStFy6Kshb30E+zefYlyMvuxrg8rWK9Mi/V1SdWe3hZslD7xZeZyWCBR
2DYAZkBgEKfTqRC17HX3+JFTY5EfBCL+h5v75tA55ZgV34z47NHDoUe7bP6VXnoMgbMSX+ohhJET
H1+jRietLrmNySBQWvfXpwhp/4tszrx/1bZW61x/IisqJJMW1l2tgFX89a2ovGCqMMcv0ik8b8Fm
FLbsAIU3uE5xOZdV7dp7qV5wGjp84blci4HBP9oUeEhPehxn/0/glyRjelrdWOh/i4GWg2hAgzD7
V/0sC4js31ZlTBFLHLx8j0dqwePjLL1J//wYHDEUr4Sj/2RWIGF9mGf7yk/Hd86/4FbnZb5zxOeq
jtqTKt5CLR5bOqms8XAbt3+cCJY2rybWxBetV65pWPHvSmmi3s2+8oXrI/wqRJpkhZoZz5QAmYDS
FINuEs/CgsrXmCfxMothbmDl7klBvUxAbZhr7wCCWe0s8M3Sxi7fknMo/BjU56G3We5Bet3w1bmZ
mi8nK+h7Lava4jEgXA8S08pIBPuMHloeQXc7XfF34zyhb+C0Sz4XmjPlUXZlFIgQhWmTHnj2YNs6
Bf2B3BayQbc8RT8DRVIggQm1y/cF34+qo17xtL1+PNrIr0l+EbNRsXsiQ8DSEZbZsTNL0vf2mzJA
qoKScmbt70GWylM7ggL5xJxs6OuU2Nv2Vqkuv14Adk7UXSbwH/vczRK7YYlcK5btPORKznCMaxWD
PwfSL+1qGuzF6gj5uth1InMNP37OWmqHUmPb11qlryG3DGBWI2vO/UlereockMqTMvP1kE9JrAJG
ErPJ6EaRt9n2EIvTwL0NRHa89Y3cDoN4snktuUuSZI6oiBZFA+iLC1pSl27UAwVkMhxKgMglKD0O
dGE0yelw29AnAr/HmddXU5B0CEyXixLI3Y87zV3NF9diiRkoxEJO7TWw0q690GPpdaNLoYTEKcpq
Pjej1poHQLa9a1mb4/wdXLURWkJ+hXTEISVvh6yJPfrUG/1+tj/gc+gEyE1UMpsZhLHqGKm+Cfil
iq55jn1CNwS9LE++hdIMKJySJycpvvtFkFBOg2va7U/F2KyvYZUKn8yHEjFWuqOWqNN4uI1BGS17
juP5WNIXVpTiv+IuP6aGrJ9CglULa1ks0ZNC6Ydu9gz9VK8f+qo2DFnYvZuXSoxgUN+qafQhBDof
NI4e1RVL8nuk+lrwfa1BGu3zn053w6cWuU1HQwV/tcf5JjMpF147jRUGrTqRr2LNUa/oHWB8p6lM
VLyIHAOLa7y3sDE73I03+AwSMD5MNQ548GlWGC29kSGDJh91oiFF7Akb/T816qoVQ0mWzPQEoggF
QOBipLqeZVOnF0QiHMH9C4IYi8sR3qNlncttvmNZX36BM2tWUO+oc8u2ydMss3NgCfZfEii4jteE
a0tDruzIEvAO1zMz44927HGc5OUXtCjzug6ihHtxRwDCY0Z/scR8tvzBBNpy34Qq347KlZownAvb
DXxix8C1CNJadravUm2riMajUHen9JNJ59hL0jzIuZ1ud92ylH/VJoYAmnbPJ9TrFzLTF9PAaZwU
1bJUssZ8cnkAA0AFF+QOFkV7SB6EQU6B3jLKsC9hVz5VJ95FAHk7kVgmDdLY+jp6Q6kp9iBsqy0B
UEHHLoWi5ZyqLI21e4kIlSHvOGJB7GdMFim92jIkDUKFYD0F+mKMAUkFXlE4b6srpLH3mJ1h7CgK
rvvTypSOD0T3aR86SxhsXrAARPIERfJisYMe6KTxF5EnXhYu/ijGoXTQqCnaSgU5TmeYyoynJK05
mOpqr3QzsBAFDbi5GfgyeJD44Q5ys7XAiW0Q6vYrFrH0RYNLhxtQ9xPa1dXDi25MgxVVOU0c5ZIx
UY5WtpewNRLErN4o7rYdevUU060+0AlHWLdH1k61Ur4JNVJ/3NISD06LC5IUXR3QfM2Duk5qgj00
tNuzWy5RpmuaVY1Q2hJ1U0LjpwvvH0aNeFk7pLOmRhRtv9bWGR7JcYlP8T9RiRJ/vi16Gqjm8PhO
pFq/PvObRaNLRuDR/8MM+Y1mk3SyfkLYK84E+8BZzfSad5KwpqDpD+A/k2f/q9VQsOzqMyn+kUxt
fmEz+Tl0m4M02sqQYgsGb1Pd9vpIkoDcJ1bl4dedLh453eYLliEZDc3I9lWctg3pcswgfsveBikT
Z8NGbW/zMFyQyulkaK3BrBx7Z9bS8oGsD3dX+c1k0qdk41+8t0IrhekrU2htDYpdvP+Qo4uP1oLR
WHq4Kma7ObTeABsmI+sNZ3E6mWmK2Zn8RTg/cmVgeetP4Sc/sobtOIeq4zINNgNZY/A9ojowrFJG
mFDnbdFRAxfJO66GJEKT+Zu90RKA+PyODY97aDqoWVt+tr6mim61ij5Eb0Xvtu9VFbH8UzS+y1G+
1yGeJ1UczIZkLibxF8qmlO9QUnpohu/CHnm1scVPFB0E0IFwbZPkPdCipwa+bxxTHj0kGOxh3A1m
803EZyWy9Y5M37r5KfyESxCjckpCs2xzC7ObAetjVXVFBcf7iCfRPHaI02sABmAhqXUpERFlMVLJ
VyhECmg841zGE/xipC4Pws49j/22HVUh0dg/tOpqj7v8PwuByu00DKI7k8sKieO99yiIQo0NHVMQ
iHYsdD1Fqfr0D2o+IjPINnSJgiUHIJtVM4WwWc/OesQa524jQ54pVpB4NRMASk8o7Lzc1cm0kytP
Ofh8cWc7dJ8GX/8zT+GriLaxKmloHJXfC1mzkLtv3C3VG2jPOPVs6rML39dE/DIgbblOgMRyFqKi
vGrcMe67J9nrHZUqPAsOiunjrBA/jLOH+v5sD1jqhxiUgyE1uFDak7bEmEb7EovRhidUE4FTw4u3
aDXAP1P8kHy4tmLdcHLJXifoW3cIG05vkoUTyv0Qu5zyjCK3bfguOJneskkEhITmrvoeUQV0G8o7
W/rVcHG3l1BphPcl17cXgBT0u69FwKPTQdWv4ncnQLPh9t0TgIaCzMsrKG36qNAzGaTS9ZC/mJoA
UxVp973Z+WbtYJAIZ80D6KjfGu9q06jU5NE1G53vMCGXut8y+Q9CIvT4EliQe6vJeXbJ2+VImP5X
t+OG5EHCf59wbTSSyR47vuQx6hIuQFlLu6FEABsVXmascAKiwF3/c2l6GiF+sNL7JYoyHfipEq+w
kzXSLG/vm9RbgOToUEcz3SVVQwfIhS7c/tm4Bk4daRLE320dsYJDq4S7SH8J5jaB8lC+9TIXCImb
PlpPCqgYvYAftkCtE8cos25nRvFpFrSbS/Rw9D+DCQaugejiYZe4qiTUMQ9fqzxcZXbFMmfUHFzy
vD2pQYxCxz7VAs7v4m9pcPJgYjO6YLl6G9PWUtvIx+NSPfhDSWzaQOHMZZPM2IOZrNSm5Nr7Nziv
LgaXjaHO59HvYvSbgu5zEbrPmxgCmxVgSqtdWz8e202LnnfYGfRDJFoDM0o+3C9CjK4vfZfaNWQp
zcbPfj7cv7PxGBaQgSikoYT6VtVSzN4lSDjXehzo7SFrR23tdLNLTDQMSWkHEAn1B7K8/REjFOwp
RSiUs59HveaCpLVmD9tQUufzP2f+7OEFdgJBWA8q6RZPyD4VCdvD/URsuLLtpfJuIGSoXP8Ke70G
2etBkZ3StvS04wEoPQlkL1dejQO5sqb4tvAnixS4Q510yf6NYiYyjGM+Fxa4NnIHXDZ5SsoeL/zW
Nrb9ERGk0GGiGPHSQV67j0el/dTLaIbPc/AEKyYQ2h+Ht81Y3K7eIFyEdUmKV+FvsjjtcsPW2xGE
aoE4inkhsCPhTx9c0MZlnZI7eJm/IwAKnPyGex8sOT2ENpfgq+J0PvMWC/yOlNDsblz+h2OtpTfa
hwhMfyyVO82TPvsqJ54N/d531yUAAkg1WwyylfN0FNILI9YA+L6Qw41uk597RTit+2YbqXg25l6l
sbJSM32TLNOZTs7epu/H04wglE1qBneQMwTVLMm83hta2LfhBS0u+SF7fRciPOnp+QbXdq4nb7oF
2aJ57ryXjH6EHcMmXz9xzyZSqBSjijEjNA9QyZTBo71rqE+r7dDmf8QKbj7mSw+bDIDb2vdEMBK5
tBUOdNx79Drrnpu3NSA6RDsbmPQKS0/Cwm1HFmukD3qPYOzt6Pe+RodXp58PPVlJugvDG85IteYG
NTvBhpM1zT40KhyK0YJ3DpgehZCVe4yt4uh6BoUD5BYEuh0HqpUni79NXdYJO9pRmT20iU9E6qci
C5Y8IVTYV1LCGvdDjB4FGZkKdKcUEHcGHI3WUJAOBlkAx/ZLTvsEx86ntBFL5PDNqZ3q/fKeAOFn
KMM/HEE5LTAVg5GNWjUTHeXPuEIbvs+LnAgbkoo/ghMdvBWZPP2ZuUecpGJwkMubyXiHOknEdQ3B
Iu3uZIx8u08kD6ExR9wFg6WuhhH3M8f19sgQ2gqqADFgA3NQQ+JUB66vTOOjUaWjrpw6r95FRy5L
Fvjuen7dQA6ws7rOrbYwAtirHgMTmJtN/8gk/3FGBhKo75UnxfZql14Evk0m4U+Fw00AI6UyFCBO
uzKWE+IPS+0UfFW4jk0VvWuG1KyRx13+QCd903kzXNPxX/BMOpNNQmnXI3hd8sqBTr3fTeAevtCA
2PfcrpZ0TnhM14oMK9SuQjvEWl/Qe8+IsFdR4P+Yb+FxYxSMSAuAmKhlA9IGHC7HyCXIbUxFEoai
Ms7Qjwom1giCpzVqVbbALuteyxGjqI1Vkzu4QuIh5vDSMeEwIQcGKpmir+tdVYPcYB924fkgTejz
sTSVeyp5JjvxPgAASZ7eZEoNDDpH0UsMj+UyMVsmItNehNLbaHDSJmwxMTOkckSVBlkEiyO9K3Dl
wfrBNAzq34oSH6s3B5lOKQlQ2I5VYwNyS0Q37a6aitEUzhfY3FL5Ya6RtIWdYVBgh9TSpHu2Wlr9
ghQw3tPz7mATFqN952gloZjEmJgeNz4Rec1eFvWlgLxIJPTb2rLm4Ll9h4sfBIp1EH41d7SmJHt4
/Rczlf3XI6D2LtZMle6nsxZy6yvhz68fcEgiHMmDh5KFTq0Rarzfec9LYbM8kEWGpUAzSY/hqTLy
AJpIEPMYJJDiSneGqt37s0AkeiF61cu+WF/qi+yoZ8cGP9y4ytyi5qjTUobF803InXysGduKFPGY
kGOMtCKEfaigrTMuc0a+EKUhhybLvjI/JXXTk0vnIWOFoMFUkhpS/7/TDMj6MXmlSjuyoSMG42MI
fpgMcfDrj0ZDyqtjVm4b2cnRBjHVr5PPo0OO2C8Rnf8HzB/iDEvGN/RrZD9VAFuxxG26bJUDdY+N
WTbAicM4VL3VpY/ggLOnSHN4p7jJqaRKU5kWxQdgWJ5J4Ah4sB/yhDlGZygb6Qoj4hB4c01KT2WO
Swh40oS4OMmV7f8EjTAtL6mDbhBY5eJ5VFx3uq0nGjGbrJlRvchpOIsVDI86kbg0pYRtVeOq514m
QjKPQCJoEuCXxxkz8OaJg9bRhD9msmdMTPiOX1NT7cVOoxM/P9Z0yfsU3fecZCeN7MxgO7lWo6gn
9BVl27Z0TR6p5NTHY+hZgdVqdCIdWcElza0TsRqDPwsyEPnOEyeOjPiQOWkHqW1uQsnLsxYNInHF
B1pGe9kjwVmVX4O19OrcPxTNzJVcy26OwvfLuPyUX9Joh5gMAYG1EA6bXCG4Cknw5GTU1rpo79LY
herLHvBoeJrKX9HOg6e+zeAVHM8SbYIL/sR/MyJ0G24nP9Mxz046aTafm4kSsFwEjW28C6ur2RFz
ZDEtUtFQsoYI4BKmX6WVZQA5lUZd4msZDk9uXNlR0KWlqflS9h1w3Be5cnuYrba417rHxdhUaeas
w90SU/YZaz9D/IGpSTkjLMFjrPyal5cj4BrpgOc5GAQGqQAtd+teORXFlYMOH3IrZ+766NXJgFD5
f6Piq3kKjXc0dyMp/hyMiDU3kLCPjKe2yQjXhvUNW4t4Jw52ReTKdBa3+zshGizjWg9JKyExi74j
B0PSx8pzHgdYrogGrrVNw9eGpVU421FWFpjhKc+HWsjk0McCN00tp9beM0/IyhpmT4kRrQQUzGZd
SHhzhYnptEnvloOZj/DRjn3K4pIdKAkOmspb+XLZyuBuqCY0HtXSGRifwaH0mSXGKrpR+bVEdnhN
E/CSarVuwYXeOgVTqc23jcnAr9l6CGw75aQpViMVM0OS1hB9DxTwOV8zU6goduwLErDevW7ilFlk
5AcZd5cIvCmDdAmMydwmkzWjC+9uWlW2NNYRdMlOR6VBZpqoN1KKHprwU/La6bZMLYRaPJVp9KIN
ATUy5Oj3iBplzOWF87v0MF69x/a4kl3/kj+m/lYzY3WJO8tYCLdeRBwnapbBLseObeengl9JiV8q
nOfj0TeOQu78tKkHnzR3dLwR1kc5YAjVINktz4CFdGDNtC+lKhi3u81pgLWrQDT70oftXmPDlwym
gt9mvkqlAbNQq932ZvP0oS2QlNPd5IS3yfvyDwszfS8wac+3lvyWTfth/nkRvQU6EUJ8yf2PfAFh
QyMmzrT4BZTObJ7gSFlFlOcW9xEZzSG9ioVdDMT52uZqzOBqN+r90HGJ2vMMWm3jOZhzi2F4GVV6
HiisnaVbOk9k5kNxqHS/ba22X1IcYkotINwcRsLFG019add5uzPzgGJPY4AeCeU2659hMjtqKlBC
Rg00vfSYQoBDxHRsvPsAhg2E2V1by2tG6T5nAN3IfKGo0u1XMFe7xRbUk/WuxAeRKB69cluFVFgX
8CCKpk2bo/YWwbNr631qeAcXVVzh54ma2bHhX/k3SLGVih3oMj1/jFZtQbS1hI6nCGTOx6IgQoIF
qpZk3jN6stSPSpPVNc0EFWCoRLVB1oF9emjwIP4QVIpiEBNsrMxY+a0rt2308ZTECDO8wqIMLTGq
zmMeaYb5bmFOiVvvML12TgO0yYobjZVEDrGzd3W4XiHC2O0BDei2vZ+YaaUCpXyKu0I0iHRjbyPl
ZKKAppHty5XG21a7NUkPQqnZ5P30/pm7tHF2UyI25MGTThTp3XbCmNAhZrs7R4Ysvahluj1HfKGK
BH2ygxYxqb5EuLK9RuK8SiCJlhtXWFiZSaKs16VaGYZLWCiyKQhzq88Rt2BeO/w7H5Rc4CuCqTUV
Tz2j5AJQOCcjWEPKgChsBOLLPMsuEUkvTwBh+CNhdg5L9Y0oVQYeaahN55P+f6aZCdQnFrsNXJ7I
e/51N0w3oZPivOMyqoUhtviFncWlEq7bdc5aTFX6qs8Ow2Mlufg2P34bglEahAygxb4wQgqW0JhT
CbFu7ox3mFxpy9Y5oUKN+CEn+7SWK9vTaswB+6MtGOKf1oLdQq5qspmK1xiZeboYMC39k7kTqE0U
7q0tyJQQoFz8rZtihNEJm8YvVxZHvChh3UpdMMyoYENwChYAssOcjQWIn0QuQM92jULW111IB1Wu
6dN/ooOVZJEyDVg8I8Wh3CG5V+djIhgDI5h7B+NIL1SVf0Y8xCMr1X7NVvsEOvYw8dJHGM1ioagW
YqVr5ynrGNccTCeVAs9WLD5qdjOvVPf5ccEc7PFLfgAYNuI0DvUzUGuo+HBx31C5MXU5X0N9nPFu
f8W1EFwt1F6wxzmk99J9MhVqXOV4euFO2AT6q2E0W8lCPXmj28w5Xa/ot+lAsm3Q1txtg2Qtp/Ud
6FZdWpYaYx4rsKDQaSdw2FcIsi8wy2qLwMjLsaZOLd2a4iaMrMH3LnaK1zx8Mr6O+TVFv0CqFoGJ
YRXrIg37zKicZToJxHje2vmIcuIpnNajT9LXGLdunU6FUl8CpLIULRe3obts2H6wL7uGL/PoKGgr
CT1sgsnii9LfX9XVwlj6awluzTRaFgNWfBDt45JE9dY3ZevQo16CvM1JCZ6IIzn9DUXVCONRoNnd
LHZ8zzTbiGEBTxVSSxp28HaMJNYe6x4Z41EU6V+UILT6z+rhDXxI7DegU6o34vjDW2Tp5/aMRyO1
J7AdUVdua6y4nDKKc0VXwXyuqKvDOBDuZDpiTIEkWyKjufZhWD8LV8OmXq9E0QREBOo2y5e4firT
WHUdLLcvej2vmStLjV73SGqV0NxpoyGPW35oG5wtWPDlGDUyhwcvvDs33/AaO5I/5KV0DYJHa0tO
fTBhAUTGl3bRDub+A47m0Qj4Om5+tTpQFqgUglMSH/92IdZpAu9TTFzKTasMRnHzNLKwCzGGaZd6
SM3piL5Ccd9X/O8ov0k7ryFwEhSExH+deJ4QNY9RjFlMXxHJOfdc1KxCG+oNG+i7ZA76AT2zsqYJ
xijOEjfMvT6opPXaXrvp7fILAZtG2W08aLpD63TDOGpMQljXAgn73090Fg3NoqIgfNpwJBzUYfBF
7BkX5IRxZ5qAqdKGPCk5/tkrOItyXWUvirjSvwCg4h+uug7spChGtDRUDNnVii91kLdtmFuDUqac
4tIuHqRVT9ESoOnDgd9wWOen9mUvvLvSieJcugF0b14SBE/mdFyG6xLY/1ngPR/ARq3sRgxFl6EQ
Aou12mVQW/rg2q0VCL0ncrxO6BLgeUck3Pc7zAUz7WifRkdTVKWsU1TLtAf+vJOAxHrzq01yuo/O
ewXligu00N/cvCezy5blmh1lV57hRoeK+Uui3DLVbF1/pCg7HZkbPxjrTeluK3X8N36buc0gREWp
YTavFCxIRRKnx9Wxz03M5JJYTpfalK3xfWqIYTMg4YJJ/qSLSPC0n9Hhk5OuX8tF2sI0NJgK1WdG
iF2zxE0CHrle1HSjWeqv6/OfXwSb5XZAsMle4aLiXMkBU/Jh/HxmExFRuYBoY+UZICWWHUO3vJXd
wvWxKVYfF1bszH+XGAJfwF++k/YC06HsjrWF9YvtiLwIVpABo2yM30v2EbPJPGj+lIvnh/6Q7vd6
pTPrZ7AhNxPrpH0GfN38h9IdEZQiDq8+5y1kF+IIcjIhbptDa6WMANrO36l2I2TzltzBVsgd7kaI
AU/i+R6aPTDoH1BtvmsgV0rCFSU46E3nIbftibr/T45M4XUY/TzFa9IhlQnfzS+dqNNgq2cAFLXk
X1eNXc+aRBHCQaGHJp11nLuq5ptLPkhy6a7GlKIBNf4SyNi0UFwe4g//11EJlggntZ9HPdIeb52d
V3egEFt653p4bkC/+kFu5zhzxcxj71qH/YH/i4ZthrELLY5ZkZ49z4dUieArvyd325VENhldoBZG
kcB43LaWKYNabiKC6MkCX4/KWB7l/yUjgbnPUwz8sIYw1zSnKBKwfku8rQZLkUx2m73hTr2ouuEu
RFEhi3qMdhikXyceXqNulTFSUl/p/+grruEqyCxRW6qrmniUNSHxXLKeqG5NcfYltGrzpY0VQFHW
eb8ELpx2qo+WYmIRevmS1Jdm3/lFwbGN+mf5EycQ7v5ouBZtrP9CyrdLHX+5V0Y2UPefcFC35I0C
K28p+LQsUQxz/MIj3Mn4mHDmtLEFAQjBjlGJM40QRM6din6UpE+OWrE9J1DqnYb0EZuf3Ar2xLvM
ZMLl1dDkVNVXArDk8l/vT9Z2M8uey+9wS8KSAtrgS2nXTMBM5wSqjxVDkxJLLAFhrFk0LjWIpVSJ
NZXlXTdsV+6vaQX5XVvHVsOVuagrXCblq4DhjoQM2exUiioY2DH4F2PJoqnRQ+DAXrim+yn8Sc3E
3JGxDGEkLcOnXm25eP28GUtL+IeEYZKbeUqIY8tnpVjtzL+z0hV6QYuZJUysBi9vD70GGLEvxV5i
0i3sdQbrb3aTeSSujzHOn7urP476Jm5j69+04+GSqJlVif7wJwi1BAzK+czFS8Phvl6HXX086QI0
uznc3nvFB/0fhJHZYqjDOnmMpTM/F+bW+0F+ueL2JqlDinFcwMk2ANVrwxED4U3KNXx5YjLdXaJ9
fTFGA6ic2djVG4o7CmSBzJZqKt1Yw+/5ycgLYYvGo5bCVkuEvp0olim5AICTzNQAkXDsFujqnRB+
wbZru6PwAj3xuE3P5Ytiukh/151CsPPeY9YBIqj/em1r+91yvQxnmmde0vIPFeKnESW3QWnuZdy4
yPKvNTNZoeRjoLukqgf6KJENge1AQN7bAARVSXdil0XVbQuDg0GQs9eYZgq9kXXLrnpy+wT2lP2u
VDx/g1pU69dktzHYVFzDDI8CNxWWHjFKICjgNrKDM1pVL3C7I6jZth/MLASQ1ZI1MceQAPiwRXkc
W/xBUcZZxH5b9uEcC2Pv3PMX5uAZ4tOmWTyFCwXQkhUcCreUx5s/+j6R0AJ1XBemVmexnyZzFLIR
YYXVQFvQ5OS4+AfR1GYwjBFhNq2hZduY8joL++gltDgHGhv2dG/27/Ip+jDuY0ivsXrvzDfFPtQx
RdxK3drvjqWdR8nEMXijO2KIBeRtj74GcRKfUD+R4b7yWswE+n8Key7QjXemj9gE1QZIqj0Bq151
kWnu+CQr4LkaomhZ9Pxsf7/WkrSK7l02yoJr6/YWHuYT9Q8fcQKOaw9mQI3dcP5pFZRRBESr2djO
9ihLp2QguvQprGaZjybUdQnZmaQLNE+7AAyGJMoGmjhZZeDAXJYgUnvwulWWvyeroazhWwrlNcy2
4+v/2kMYlatuPZkvHnmWffLGVHU0NTgICb6ITNlBfGcIUk2nt2m9bF9TZVepL9EFJMz8VT2HFWLD
RUPGJ8lxLNfOx4m8pK/GS5OvUmI1VE2htWI8g022bRaEEnVm1Lnp8ykz/Uo25+K9rki/95btbJtE
X4dayV2SB+4Rr3C9/pIT8O4c29BDM0Q6bOm4uck8NgYCSGUsxkNuBMskDGUmQsa7mGAo/3ZsrH0m
g1/WnQk4DOfwNiJ93SUan68LPJO3+f+BvvigasMfGHVMUC0J2UUqYDbQiHEu9FQ4f8rpQAuJcZ/R
5nKRbHqxmKoegI54h08q4hVUMyj8oWjBV4NHJD63tWQvu5QTMVIx0uISFsT1yRAki6m6sMAsUGg1
4v1kaOHQ1tVgbpRARqOWvzl3dbz7M5BLHomhHVnlitFojjS5i/8Zanw6BT3VlB0qOCkmQkwCWNLt
17WkqS6ti20etsQcT/lD1A7jB7BbmIzRSjy728IfEq9f1UdZOHbUUnlAbX4eYZIi7D6P8doAUbA6
+wYY+CmLPD4GHe+mzRB2uYXxSIJT0M4nZeKBwz49bLHuVABIdUj2y4w23PvimbWuQiZkCadYs6aV
R0fzlVLWkxykV+ESYviby8EmHAdopXxImnESDNoMaLtSax8NktvK2h9HrbC0BH+hqetWNyhOs1DJ
YMX764wMOtr6JujvVCj5MTLuU8pAmhU2Zm5JecAQSRgvis86/xLHViFsK1rBXG487XVPB0AtFpSe
TH5QJ+Bd+zg2qk5m8nE2v3qZPp4pxGnaVneT5Z/8TbdHiP5iDgRF8qUSC/5Brn5xklg7xFeMOI1v
cxpZCsEIoq4XgDg+3JhjQdF9umZUu5Ph6IvNhU0mEFYJilsasxTzUuJZoBE80Jw7x2SsTDTuUR24
KKPqowhrKfHurn72kuPjN3PUl9a7lCqZl+Ya2H/62efbLslFfN/98l4hs0c4wkXNK0IxbUkJkeDc
gxCIQRTHFVOCfGRgS+fxwyRa49/TXAE+VKLSoWI1uBfGCXHZQtGjEpexh4Wb+XFF6G6pEoO+wJpV
l1xsjRVbmSItsutkGYYHLLHlT+3uVe7I9o6vQhe2JHpk4P/6+/TLePR84uInp4UwqT0xlhWlStt2
3l2Uqqrzryd8dpdiINhxuaa3D2wK77dRhlvjXx2AQTqWqgzXxOnQ5LYA9sKYgfbsG5G9ikMElmnz
1+vHECoq9J6eiAoPbRje6RHOk5UENNLVNZiaHYtcpJ0M2NQgIasogmeFeWyrliuBWS+O4GVsZuUW
Hc8z3iqVTn2rV1QHi9NhtrJr+JsgcC9DLxzpbWAL3dUwgFEb+QtwgGFebVDVtLtbP4D0uQ15zHBQ
180C+qoKfgfKNIaitBRFokO2wu5qb2d28PEzjWKAbvoJV0pbzMESCzPoVa6hBRNHuMPmYFpaTVK+
207nODe7KUyvBs3bybdmiYucJCQSPX7OEc/yAUx6fBbPTxaoSmdyGjUbL6NBs6MBrjOjWHNrBGeT
xv/a4Agyz7ThqDs7t5hVrH2U8L40s9YxkUeupOVOmglYFFsI7202QVm1/VbbEXGDQ7dA+QToljb6
0DSHCEnGQ7gyBpsB3HJRr/6Y/Wer0/xlCEVozhl1v9Ifr2S4SdfreDjv62wNxdZDSyC60UpAfdGq
MeJiEaNKQyd1BtgOA3UEOvu+hLfN7q7r2nfy2tnDW1yKLp9P/9/LtU2tp6khWeN8i97dFb1GB9dy
vhfTIEPXqeXDx78So9ucOHpipdU3SdYvUU+KlzU/5AVQLmZ4vTBBjCdvkfnOynHpZzns5Zns2G9x
TnaGd+PSTEv8lAUadxGoFopadtwI4yT9jCWLaryHXszog4SK0e80MvGGnh9S1mc1gv1ArX9tI0b7
J7nydH6V3V3QjvGAOVL5mO4RKwGrelhbnFfCfhFUPWASyXDN8lpwLA253Oxe5oqo5yQhp1+wxPCb
OCu2Lsn73dnlzG5PFUuqtjsux+ntB7MoYn1ponhKEJNi5U2Y6YMvDE7xckegfEvUAw1wQ5OFbj83
/2bsnsRLjVhfvX1GTRBT9A7dzNbJsNN6eRqX/snN1ArAJIL8PWFaSRn+zZp6bny5Fp/zI0PQPLrN
ZAXy9u7tjdMKDZyff8+bjYkycMpe6NT2skpwO8A/iM5e5IB+k1yo/D28hX+zGQYC5x/dP8S8+6Ut
kBSZv2iKtWbFJOUQ1rTHAQKyLoylys6mUt2iGJnncdf+tab2RSp7YhGpFKnsWGELO+MycVc/qW5M
tFh9wLaCjP7mMSxPaTMP+HYmo3iIkCC0uhdLwAq012/nIdie0L/Gux1xpUdhzPGZ8L55uNPNS3Rq
zwKvCo+ZepMt0D5keLCeE1iQS1/kpMERsYHJVBUO0TTsi/dHTAISUFV9X/y1bioXdR32pfL210I4
5rTAPLMCRMZFd4TdZqUls19K6uxvq9AL3BVPKSoeLgkP+VWUsow/2GBm9q7iHXHXHQ5e1Pu8cmGH
nwYXcMZ3biaVN6H9mbo3rl0y+d/mrjUsrsKa/qNCFNcjrdRJg9wCqzXvXJ46razGt3tiCeth3GS6
tZAHHdo5JPACf/Zeam3XHvq6ip76yuOm0vY5CU/SQuh5SpJ8tPWff/ncaph6DvKpyYd7ot9IR0dN
RbnPYL426hjQbC/4WA/8MXEMqoiqHpoxN4zFx54G2HvyZmLnIBSBmHtIs798Pq8XGg+GSbFaesIo
Gj5wKWFv4RVTuxx9CLw4yW7qe/QMXXVepNs/FnWcAFMW3H9nfxoOCklaQMMKLDOJsLMbSPPAkfji
7v6xs7zMtSRzBNFPtiuriTC2yWpLhwX/DmI/SvB1bMfoNSNBYgcPrw9L/aONpHWm7Sg/aJKtyk3l
NSeX12nkHWW4JJCkrSA/7EH5/IY/w4P6xk8xfQMEka5ZPttTfvJ5ZROHSIUvuobKyTI4h/oyO9Nh
/j8Y2wYFTX0xw8RjvqjkYU+gK1rx5p4e9XSZD34F0797z5a3AVW/pJ459XGxxP78kuYubRZD8S/3
/GQd3JG3lWjUzwJEaB7eT0nsqsk3RCw4jWfUoH5OS75DCFudl09Yly/UqpT+eVpSHva8zBenpmoD
dpUxjw9JuYby9CjAaunUngNFfH/yTIm//y7xSqyiBJS0zB2bjmVG3jZuJ7DzZLdgbMCfzzV/GIzB
i+HlObLfpqUsfEeHPqBR5wvVPFrcHdtWiU6wPYIUgn9v9QMP65xVhNEyw73pftEF5sa812p755/W
yVN2OHeVhI1YaoChWRyCcLWAY5OI+7mwDk6pYWRZqRbLi+oaURTZ9a07t0AANKmnFk9hqttXM/jq
Vl5A0+cA/tfJ5qgbRNsnGpc3N1f66/NWi2M9wg0NBdkT9+jn9gGvUuqoK57y0t+pvEoQFNLraLYQ
K7JX+nxYl6axlCE9h/AGwyqsglefJSjGTYTjUpZX4YofUMMUGSXSpVmX2sFPKYHHTmhw5YCXlegi
8nYT5BX0IIoTsgmzAVmhO7dzLddA32u99kXs8k8U5BGp15C1BE6LQw0B4Zz6WIFuMsx422jebp8m
8qeE9RX6e885fz0fHTSJNyXn+hoqSlTxKtypnduGWNDjdSGiY7LKn35/PjAOtEUdd9tQSjyI2HVI
bdGShSozaWyj6Q69c7Ap95loyvnM8n0CulmXLTOpsQT52BbxkDI+4sT1HsFRPrMJDfTUEoL7gNCs
dWvEMRLleZIX4iBOeVqqhOOL3ObQClebJyX3UlnfTp4oRaSCLouoVXfossYFVXL8OChp+NvxFDs2
80z9C11RLrZ3FolJ9FkQ9lPq8FTDLqBUSsRFpe5roeu7e7rStgW2Yt1xBT/0mw+yKa8DDXtkxrKy
ZUrvG/Rqi2++opACu/UJXJ/JsYxGiIm2JIJb5Nw5XXSko8+XHQH/aM8oCw0sdyehMl6C6O/PNzTk
kS4/afG3Rnd+0mLt7d2l3jCAQMs5570e/3S181pPUNbaD9w27mCmXMIJ69cGZRsGDLjeH/mJSp9d
UdFM8dgAFFV0Hu84zuod4Tgz7lhkF0sXy0TISUcNfokMQPPFojbIctvcILeb5P6RCv+HoTy9q+8n
DvugPPw1T2JDmFhzozaAGSHQ6na/ab2CIUxotPoQzYMOJqGKMiGAUhhKdRBEqgNkLZmSjjhHtx/r
k936SmEVoOAVV6N4mMJcNSYGsk4Qe7IcUMN3hdUnfbw6QUB06rmZETUOnEmZ/gvnl7xodrKttcr1
kdXnPRPELxnSvi0e4mVB8mr8MpVmjjAy+H4JLbG6pvLcrVVKLQO9H15bhUMyAh0BrjA+JRwkvVL+
OnPanSrKu4ZmCbdaZ3bpZ/pFV6JPv50BHUuCK56l3ScEtMZxpkwoX1sOXAFvKS0FCEIYWY0nd14s
SBAgATC6dznB7FHivKCTHbm19+8GWWW2Il+iKkR65QLmdxIwf1OD3nIEwnmWCQh3KiZ+t5gxjjb9
HpcGn9/w+AFVCiSPKFzPTBnCMEuIxz7uhZsGkrADQfeuAhTI/87Z75P487dj+YL2YOOuCdY5t8Ry
2FSaM/IA53Awctr39QVxNzdKb2dSExZV6U14cldSafG4tUoFqyfD0ShNWqkzl/xwFNUITxJRdm2w
AEMC6VpdEq/I37EawuS8KWHs3KUBJsla9mRQNPQ4oCObgIthE70rpUgh9SelFcoFV51iYVReYFY7
GETkXKMnPFdqF4s/yPDrRJvvkW8qPZE5ZviyvPXJGedzOVRQSk/whw93/XlMw7f3o+JaTO6JaeOR
X+WfiFThfISfOboeOJ1JPcGYdvAnhY9x1G8Hc7EDY/6RbSl2NpiMHS1FAPEeEZmVPbhFc6rcV4ch
Jm+vm4Knw40BCG1ORsCgOpGQetPUJhuAdU07OeZT7cLxDPAxBl8IFgfF+Dcjo1BBQ4PVibS6bb0C
798nZsCRUA/J7lfPSBzd0VavnGkHFC4coWZQ3mGFzwT/ss1wtDdJxoctVknmt2H1WjOF0oqMeYan
6FCbnlS3v2VGYBy7fs3ZeG3fl78rrhqszIch7zRxQxvHQX9vaOSpIpPKrYVTlduxEeRFhbnyNv/m
7WdrIn7n93xD8CgkYr3wQquUGF8p3n0/XmI/3oIivD5oI/gQYkbazdCEwDBA6a0sVsawjdbbCUGT
auqvKflGqYhYZ1NhAo5P7Cwqv47ATi6/cB42A/M6itzg6rjrYM/IVER5yoa9SVFGS2L1w/DHPbnw
5VoQ4n3QTHiFgK8QUJgy9rm09WhYvBYkwzeLJrNnB/dlcMsNOSJZMmASyVY3r3MyusNFGD0PY6zx
pYxES33JK25TlY0uJqyVVuH40SgoqVAfFg7S+JKGCwgHelBhrZ4DX4k0XeqheV2yoZ1ZdB6iNqu0
EztLJ5+cGnvjoIGcmpImj9QxwW52k5v+ltkHZIy9/0ju6LoAqCu/0Y8YUnWWZJIEDhaOVOLrv+RU
WJvhSgZWOFx9y3zpJjb6fUwKmd5KLNYhmdJvcg3woxPlO1zFUUPeI2l04aoDeYi5/Lf4Id8077d4
0M8AnHQ5g1EozxWmE14u8EJO3Nna/84+SLr5ReHZ4S2MBmXnK/og7n/PdAgwyjECM9sXH8nQUwgX
QnKQ8jO1HAIVEfsJ4cHSICrFqMNH0aqi6GFwjqDf27SaJ8y+hXoyYe27C0RrorH/0+CoJsRum14W
8/Ll4GFt/K1Sn6x3Ex1sabH0j/+/X4CEx7en5q7zwZQtzwPCR3UbAqIxPsetlU7jrg3mpN1eYULN
ynZc6JokNyOueAxvQEtfUXGieaLtPJI4O4fGxDo2qsySHTp9L1SLmiJG+OvpbFXJoEWL2jfyka7J
C3hwfVBzJidKENlOvXare8h9ozt5DWMoG2M8+YtzN2/dL+EoAYTJqJB45wLrmjL9a8TnfjXnTsns
9mY2EO1O+hmf3uQ4nBMQVGvQglfOrgHj9CtWmPDY1ovyh+xjWRR4z5p/9s6dPg8TFSxDnx6Xnalo
Ae/T2Mw5qkU+2yoTYbr2qYzGsuhBcEBhIP6xCKxCUNG6Z80WnMPH1PDGOTgqpF+beZ8kIGPNzl0F
ekhJZd/i0fGGg+lZFGlw0O4Zv2MsXDxNF+TPRCIGgtvv0DzSbRSzkTuu82kfa+j/URT4+DfdEfuv
rnHc/UkEVvteyyL3Ijw1pWtwZPMaa+2FxX4z3gbe0U1qRoxSeZZILI0YaAMJh6NsaHKLEWRmtFeG
Jnp8tb8HS3dMrQCkNbl8XvQFiXPSzgNR8odHli/lFIRm0xaYtvZ0ZIpub/36L2/GBlUsIKgcIofH
RKY7N1pI6BUm/b60hzZ/wlB/MoXVOa7oQqI5iI+WNdpM0dCbX7d9tieGprEYjFkByuCPlQ7VjXVA
oqVJFo5pPY9N4gs7dLd6UpvGQofkXE/Qylm1DevyKVy9PrZGGmHffNi6KOCwukPGYhHupI/f4Zbn
gvnZjwNXy36oJDmArvDjyHz3lOoxlafW8ATJy0ZG6UV4l5/d6WIM2+2MUqX8Osh8Bg7YAFM/VEa6
N/qT8hhCMWLQS2AMnP0mqcqV7uOXTH2FC27NDbyG7/bp7kU0v0RmGspg4HPS2Ewf69pWMgs2fTTP
DeQ3NtcRM2ycyXn5byUNgF4Lnp5gpYhCu0DGRpaMD5fuS/EcTTHnpsg4fvsY3qk6YaD3V0/2ouGq
gg0VnpkJs7gKhwe5v+HQpCJX5CmVQrNxEbrKvJIIWEbcyya4607Q18e4H69sHVrZvGxonVtsTXKP
u0mE1JJaB+d4aSHyZyfxWTq33jvFSeQW1QBt7JedysGQcRGqD6ALsEJbwo21s2kw7B3DP7Y6SYwT
tMTYglxk8AF62rNrPhdsMr3kxq1ZmGca+pPAa1ga87qeKdaEXP5VC4vrEs3EiUmsTGY0ho1zb5/x
/qxf9gBud0Fdsrp45gLAyOybRaEGM3QZce02YNxTcTw0kx6ZYTSSEFLst+59MP3DO7wBkjjlD9uS
r9nJWQBpZpsnl5SQHPm9veusKZ8lppuwZUaLmSfeOxRrB6LS25zNa6u3VmGdYUkvt7+uMjOMG0kx
JRphfLI5fCCBz0WBObaKuvCWeTyVItiMHyI4tHO+upb+npErsa9dp4KiT9LGSTa7fXwcleNM0QGx
WBytIrwQnOnjjBLrtBsdPUnT0fxIzDzzoUIzA0QkQJu3Dr3/jjTarPJIOpYRuDyZqADalhD7bCEj
oI9EqHwux/NVaEdiKkgRRIF0H4CmdUp/y/fqYcLYCRv6n3Fmp+mjj+AXFFLGBglnXOEe/sAV0MmM
hQjkRHRVNhGrPxLGaNGW3TF8SoPMFx91zMqlXoigGeVkyaOOWkaRuEBWIVQkE4herWQpYcH9YK+t
+XhJ7Jt/+YD1OFj/pPivmbDokSklds7gFgB/NPmQye1OKVUkVFkPFJQsmAxFJRp2e72aZuXjlKdx
OthynEtUn3/oBsObVH0TIuBNyLXfiVzdHqT+AIZSl816hsBlYg9oTmf4JvPHzv6dP3BzxQLVkv8g
gG8vm4ALB6irl42U24OfpBpp/6HIIhmGQ+v5S5IIPlEId+rp2InL5QVflrtrniHkkXV58P917DDH
jI553BgKGoQ04UflUKvSmyZjW4zeWOkddhGsKBbzSQmLiwWhm9BnB21zPqitfwPNDOWH01fQcFAm
4FtncZMh+cj6+4fXcCvWnAYcfMhhp1flT1heY49XSswBEZKdSz2BcPWS8uAsohvSlwUzn2yOrWvZ
OC8yXu4zfgulQBAu7ljTpdhPaN8ktKCLYefvUEVCYFNE2S72ygYlwmWSvLJRviO+MXtlcoNla/L4
FzsR/5evG0sdTuWhH5auf1ZsITJbbNQj0LOp/GplimkMTKPPL9emh1Srvp+W6sLTSpINnbnTR6bE
FHcKgd8YyABnnEF94IGilzjQyQhD8d8zwEpIonS4N08Gct4/r5eAZUWbjKoKhRP4oQnuS6PEF6ef
cnbBuaqRcK/kmGisvIDX5GU2PkQBcVNuXZLqdCiMUjevZsRLt8dUqVEuhXvj2z1LiwlKPtCGpfOT
BziZ+qF9ak3JPMXzAhNu9M1oWfHoyBkgq3rznk0BFUmB247yVFu2O6/g4WTbgOhaxHfJIQElVbNJ
WpwMnDNAbP1+DcXHiAqONsy9HWELY27+0+fmaNsaPe+D1bqtNe4WhsNdvIC1IcrULjFQXY+Cz2lV
rrZokByEwC1Xux1rv5+2xn7G3Yq/WC34ey/HM/i15EFch3FXk4niAD7QfmY4cNYKOReppy473xHW
Td9ysFfBbRFvmztacBox5qtfEKjiV108t7vJmRb0kiAyQ03MW/XIFeH6aBI4vojWYoptTQ1sXHyR
QX9Z9e5SdDLaHRDyogtvmTvXCx/sOQP0fLRjVw/IZNi7jfHL3RT3MNF94RCnYaaswO7gWpSWKmRB
q+Oc0yU6e0gpv0sRI5WYexY1J72gUbe4PR0d4uGTK4nrRB505abgBjmpTU3fV0b926wg7RrYH3gQ
B8htHkza/9oI754DGp5vi9t1DRIbxdxbrgaZo/3If/tX7glUcp9OC0S7R9d6hKP1C07cTbUd+ica
VLfDbBVcCflna6Mp594dt5RTL0EOEb6k+0gpuXHUvwV1WhitQ/MSvHhz+w9fRQ7CwfwHf6TOFF6/
w9YU++734wj2E6rTRDHRXQgdYxavDQTRwUclq44lGzM5M/rg7/OYYILh6LL8C5cN+xEPGRdqNj8Y
ZhaMMi4edAP/y4cnzNvAdPNDlTlt1mrQbGfhRbKS1Q+rcCadp/CnkijSzsJPiZ6tf2qXeNAbcH+q
a41PABpLHNTIewimSRbx8JV9AbiYwBm0g0JiPus3Qhmcj+PLocvUVAYjagdPqVmiVkbHBVUWOJqR
2/9daoLuraonv2Ajt+NTMDZnvk0DB3g2xrE3bqz52Il+9P8qY3eWIJLifO6KRqFbBFl0nUjXf/+E
lO8cw/zaN1T3sN548848SnqFnee4Z7wscdH9GN+EKMzCHFTHdXLWFoXzwq9CDxXFRUfNSMm9+Q2K
Q0U32v0LNUqWji+xVzIkWXIjp67qYx7DKSQ6I3F7B2YtsoWQq8Il2YacFb0sqh/NwAqJPd+JN9LO
ADrP508iiRRn3kjOFUn206Fh6kJCx15AC9GZ6MFFkq+3qQocE5DR1PS9lMb2NnOZ5u2Pjb6+tGLL
E1HPtldxchTdEMO3qlfAeKzJFrNTzCaL+0rqjFOrQ8RV++bQX3HKcodG0hPVMyaqd7c+H14fBpyW
Wn2pyTR68SACBVk5aH4UsXnZFGy+93DOeISxLwOXFIYQLy5rZ7hQUvNBuVKhQxhj1PAMzmefmHOi
J9Y8F04WwA08xpjA6b+npKCQuiLG14uyJowMLXVay4XFw9g0To9xc1/eLNDABzxZPsPj69VwqDZm
a0+xC+tl6oOqAwA1ZFAfJeGgsLyUebdu/L05NxQQJs/cJbnB6sf7dTwXf0HVlWkyQBBTaHWwms1V
fkWx3IDg02JsUpEPjylR9oIlyvBkU/BFBaf9zhXlmw4CLertykBo6w5Jkz2niO2dyxTDKVRFRpAZ
L515N0ZTG69aGkz4zLcapIKUZMj+TJzgocKdnrYAEkyN65y1LyrzwPHNIbFc8bkFgkjMELYa0Ncc
v75pEaWK3Z14SswuwACyAgAF/OIGeD6dk04XzCfQyiBYhkaP44lJ6FpfCYAfp1OoSHR5I3NqFV/4
x2C20Y02M0EK/SDMy3Oa1ugdu6+K1aGqDWcr9PFNdNnjg8kmzkOIKmILDfs3jHUDeV9aosXgK6Ot
ibROl7c7jcKkm8GYEp/2LCGYNZ4UKoJSS6ec0VaOqc3GRhQouakzxt3v8g3O1AB6T03h0H1hPUbb
rSklykz61bC6//LVBRG0vjoLJ2kWNb8rQKQ7XWCoOxkzVTnqwXRcuDNIeh6Wc0uSJ++W9T6u11XU
z4TX9RyKLM3HWxr7hBb2PDx035HoSkvLOuT3N7sm4vlO1tAXmNarg0IESxha5FWU9JM8Y6bt8BU2
rLcqdY5N+WpZLCk80DqoL+GI90StBYNP1ORBxwbUaenQlwJgCJn77nzV+nzRXm4hGQgcKh/SJm0S
b9K03lFyG90mcVcH5kN8jP6OFZFVCAoChOByGYX07u4LTW2jH4L3+WE8YXARnyX6RdoGqlqMw3ni
vA22KhUtf9e9mlBUQIkIKOHO6iARVcvhJkzVIU9m9tpKSB6oH0yY6bO3iGiBvlCBGsg8PTKOnOfc
Oeq3a+yghyqoW1XxwxoYbg/UfUlhplHGGU5E0w/KRJPaOR8Ektg7zlkpfi/dQ7ipN04Klqb4NjGp
C/c8Go73xl9HdGlylIrLCOsQnmxx8SSsj3nwf460IDy78NDHBbHomyKlWU+igUaHQDZIG20bvqcV
2bbiyzKPUGWbeSDaNhpAkLv4xlFKoAG+8mBBRvh/gkGOsSKq3wcoBZTQ3vf3SY8Bv9Uou8yEATYt
MJt8L8ZT23NDyTbK3hfg73JUN0W+d9omo5RW8/WxFriZ1Fncjzq7hGB7+GBCMzqWprIQHa8SE92P
5tb4zjOTvN49PP/Z2xx9oFUPYNQDcp3FzGWkwRJAs8h5oVhLxR0VJAXkVU5mba3gp54Y2LhtTmNM
CYytFjho90xltBHiHV0x881QuoPFjaILgPKUO9oQYgMr37BFcMfX0qK6Tdg+l+B8Tfu4y3trOd78
v70NMDdHgDkZVESbYNeSZMBD9YTQhXRk1nD7gD4rIQbv4rnOLe446pw8P6giDxAvxYC5uml06Fz9
9bFBc0MMN4mshjvYQTtVmtEBwm1WMyNqyULknMw2T2J/YOYrejNuUdaXt629ZYtJ31tk6k74Iww4
ny5+xuxzhOvw7Vj8GjKGTLawMz5Eui7AdPRjHgdPw3I+Xtd+muqBXKQ1eB/sYkYlbkdmt1A7xAAO
SyWSdiNMMiUpdjtrwY8tm+tKYh0d8cPuXKDGO2HaF5NAmcd400AyzlFQMChnPGmOZ0Ia06PKdYwY
0l5c3/txkOpTmC8yYkn0w1nDWCF5vEVcN/HKLks1ruXYYHdVCULTkc+G9sWtVFSPHe8JhtcVUfG1
/5dTwnYmEXGoWlq+T8EABCXVyXFjo3ogFL4ZEf4lZZP/w5Xsqpgw2WCrRYryB9yCUubPVXnqflnM
r+izm+GXnQwFhjYrx13N6a0M4Bv5P84THrE1lgzmrDw6I2uikYkFjlqt4WqzGr/DtMIdtqraDDp5
U0LS9JESnmQ7yinYCGsXrBw6GgkusVQpGYtaNWmbTjVrwr6kQAvG2TQJXtshKZpmcjtftLFOo8u2
OSAm2CWOyQFq7TB1iZFY5bF1W9JXMeHEb/9pwwNaqbomYZc4+yauS8Ap8MRjLFXSkwvLGLQOlF/e
7n+TfroVT6P+44h999fjTfx9uXAdpwwGCN1AnFm4b2FJCuwMKIJsCk6qGQEecaQuJOwZ1dbtS++d
788gs/qMUDXVuCV+qS17rLSSKBckpEjiS+9mRza4q8Gv7H5nC2HBHocgBZasaKQzFOF/jhM1nS0l
pozoiuPFVeAePzvPq4XXwwR2xfElzmFSn9LXVQbb1s/PP6ZLQMqd9ybXs/25Y/t2yUmB55kwDNiH
uKr3hTtg3gF6qgU0COnjmMcZVo0d2pzsIX/HkUpjsyFKf5u/J2MxxfjAxMvTMqBgHBwe137S7LbM
WiBT+ySngNOg/XmJ5qcag9qGOVtE04kI+upOUjxL8E2jAjTaDnDYQJ9Gg31yFWSPG5/WZsCsbTPW
syGxpZwm+m50qclmeAF7UkCsvkcbg766etxtU1ivh4VdbIACJhID8eUtjf/faLX29eisutdqOj6E
8F/o/m9fWx9JoGHP4TCzz+m5MgjNMsrkEyhUVO+kUKQV/ivDpd2jepGTtTI/dcFUU4DtyFEL51FD
Yzqd0Cwa8MsDsZZLijc9VTVVB67BXVh+jbX2IJRU6CuquHxXHLW0zarcOqOBf7KUu5dSWYBEiSgm
S9ukwzLqlAP6oRHUSqDjeITBe5MKskY6bVTtoZ1+WmO7rSoe6BDI/LfatbdRIzM76B+MmHR/D93a
8h2HuzuwRP0JDFmYt5yNmVGnO2G30vOZ23hbg6Lewac8OPKBJssNwR2owpnt88oUtH9NAC+9/NGN
sjHxJmbIYdm9Ys0n32qWcO5nr2cK4oTifY594hDGBe4sfp6wG0bBHH/McWoCndfdgimI1FWQwho8
ZhHrMNzKjv6E++nnsKFS6+mdFYGYngy022be6y4mgRVr9WWn9gApEqchqpjEF6H+KRWBxG7iVxlA
cs8UFwmeLr7JOVmu66XOyBXpbe3hsPTig94ql1WHJoqnVHZvK+oQ2NtTmWw6JO4nApCxp7J/anm7
RSkhCexLe2jnt+tM6/ETHUd24JRvpnpyU33eHwXQLgVDqXxLkMqoQKaakj+MVYkWw0TwiPor2JcT
a9E1h/3T/Bio4IpTHFxEtVWak3xcM658O+9+xlH5k03hH2yGQ3QBHoGVzZpKBl6V52Tf/McCn5K0
n63cZKdBsHPjFqMX+W3ZWcT7Mm4o68+wBDvPtuH7XjpIFYi42UOQbltcxrcO44jpNoel2A+wqZRx
v+SagQpe/764q+0Rn6KYKW1Jth75do6a1J6D2A3KZMdHilmDWkGW/xNIM2PHPyk/D4Eq+CON22UE
KLZa2FzJ6qRJbRxq6sz3akJ/af63MxMQBeJ7AwfSWpPP5crS2WXlGNinqGtt6wAkc61NJDn5dJQy
NsUH47SIVxLkosNRgiszcChGKyMU0X2t9oUrIHQmfE02xDIdcNt4PBYXsvgbCgeMxGO2V/63zKsw
sFyDYtcUXt195rLJxXBu7jviTXo+Htk5xH72cOs3cNohHUaQfftnMsRR6Z7B+Q3jL0IEJy4HrnC5
xKVEtsDtI0OtxsLgJod3CWJCS2qGOia079OulB4zT/ktsDuMcYhStvcEozZpn/2hgDYE2XFfk/H9
xPX0NL+wiFdpGN9ZlZp2mLW9iaYf6FubEwfRS26+/AgzKOCIM0l1yJ8iawbSsrmBOJ5fR6uICIxW
rSSBIBnL3J7ekVmVfZfl9mB9sZiV4ucBNZEd+y0k6x8LxE5HnBDW25qMvupUHQ0ZbmS/9qSiBKCp
W48ZQ+W0EpmNbNZqe5Jetz3T5Px+IrWKGjIxyj5t5PbsHE5r6AMJUfaS7uWbgDrVoQqoaWc2gvT/
6HLBoOO/bEunyRW74o0cnso89FUrnDQSrCCgVne8xn9kdTLqZBPMgHOs96dwR8vssSzCFVRJTCxV
DIpAM/ImzyYjHeStC3gtQhOyHIpsZvl2+IqOt6ZjN5jFzRlL4GxgBtw/ElGgE0uNsbyICpytnzMq
3HZWT0UMqc/9QYOeZVOOXtaZCU9Je3zjVSjP/kTAgEKiAquOQFjhY7cUROc4fmIRrqGA20N/Xx5h
peIyXuss9GxO4EX6XKhsUAM1RxDBHrihirhp8JrIKpaD63pZAqQm7OourDbPHAXIVqOGwDhvhcg0
2h9ooPmw/Gr0OzI06KXr5dfDWhuf/6wwG+tCNaVAalYZ9JyCZjWtRnc60s5pBdxBZsK8jSMauOLF
p5hexGoXGu0BuuJA/UqKdF5TtevAdKfDFrEAtepbYwhYU3MtkYZkicduKAququ9wg1L74IKwteSg
ITS6RsokHFmqt/xH75ADZdbgJfl7QThttuj0AvadzV5lGq24sNrMEkMlZriFyiCKk1agU0hdYtOy
k/ceErc5Du+d/VUACbEX+pDXGSpUMyB25/iuPCSOwj83QeQ1DttzoIURsZaia1DYM2zVQCTbdCHm
G/3HdufUFN1yWhXLCRD05OWCfUecJ4gw7E9r4zta0wo/gKhHloddNMsdhHyC/DyCvLvYAoF9gBTi
PksC3SPhkcyl/6/XsuuKYeAbBGrFzMV4juuJFHJ/MvAQYZ7vfuXOjiIA1Rp6HrjrLnyX8kSKoAqe
EkgJcCwX/k5IW3Rij7Rv337PBJcBkJFypVHcPtSbpenLk4lbZZ25aDJIpNdF9UI+0e+4xdGPtc41
JZdWwTG8Czg2MQU9JmKToT1YoZF2LDiLEZRgX3g+Ndlv96K5XmKfG3n0WIM9WFRqSM11SoCCrgzS
AQ61vBpqpnJxyHMiqJGLloH+RXG6lC8yXZwcDycl3tELNru97LLNDSCEWIIwfbxwE8K3/VlS2+Wy
CvjXUwRN8HPCu76B1bjSTYFDuOvyR8F0SyxF7cXGeLIuwHXNY3ZiV9P2d3TcJeMPnq0MOAjygc/J
hv4kKT2jmI0cZl+5ZYZYSauE/0sCrVfMwQ4CO61OAydTB3+CLOebQAdQyiHEN5pqVO5FJqMY//4N
PRYj06LqLGuFavyVzR1FO5EZTmMIku07mDNhp3uORf3EoVgHnn4vb7fXK0OhDFrnhxhmaJrtc7gI
LYWBiAX2ixXyey/ZCj/7+GP3QTpjk6tSHNYvMv5n+vSV/aMbnDbIK+4vNU5YRcD4JXJxJhFt47LC
BZIMVG64I0za7sk9oBIU9Ujo5R7HuSiy7bQZUFVnXbACVP71zQtzE+3YKXWj3GmLUpB0sTNPtQv7
pr7iFR7GMINIwJA7fkup0Y9bGwzSJt6yetX6zdqwKK8mjrujd+Zoa37Ss3eZKzuoL8oZaNHfLmfY
lCX3qFshIaUG5o0yCg7BStF2EV8fiQN+6j9m0hErOhMTXGatFsxMV9XKBh1JmYAlhwH1ZXl+0I+G
WlgK45Byi0rt3ipcWb07hhkxP80XYg0fGPwM97FRKEgtVgXIHS20Kwk/xtmWx0rQ1uyqDvd0qX9M
mkWzFgrq/Ei+cDFKIdVuM9AaK821/gKiWWsdLbBwPVjfRqS/D7WWyeEbGx+Q0LmU4cgC5FU+C/x1
Nuc6wlc7KBVGziJjjNKlvyihLlGOj5L7a5xzVDZW0EmXviBXwYmPdGnwgDPzsZ2+kq+pgBkSiQox
iMs75t/KI+SMzW3jVk1J+S1W2SNGpTEBH/V5gyKe5KmV+oJkqWyp3CRDopXY9vkhA+XzuB2FJwfV
VTUpC770S5Tdl7BDGLiBUPbDDLIQerSA3ALf+VNSPQhbsiQOfK6ObzZg9GcxDI8E3AxLiEOkO+Vn
SF+D6lJpF9qDCHQRAisR/2YfqOfxcNu0OL04jiTmPBidTdwxd5UFeJmy/cDztyClu6QJENsloEw0
qR2ifTmraFOfTE3iTbwzTlwZ0+C2GNGWKvQZD8UsIMk9ZqXn4muil8510FdqsFQO30iRnNEFRqko
DdFEOdkl5XLok2knNvzVhWC0/CS/IO7KS/LvfjlqqFUmQQOHSFO3FAnl75gnq03Fa2bcQxdSPPXc
FyrRk6sp6p/oqtYxX6N0zRiBXjohWLOrbvnUzyDeu9+L30xdoIciBVNTWTRskn41C90NuAcnu7xx
/3lcOKdpINKgLgNkqkXUOuco+Ei8sayLdsZT6Q4AEzbxKa4RWsYktnBx5cmYiXevO6M+qJS3cjga
rndBySLfHUbKf2EQdbKlde1RMsMa8HI4j/9UG5//88b9Yds24nHP4nTG8K57SfeLxp1iDdzqtI51
OrioEoFhzA7eiVn93UdWZbAa33UBJ9i+mr2hB8foHn1vf6gold28ZxoxFUo7uPOCo6oVERnWMIPD
4CNFD99Oy+AY/2dVXUXNr6verXHL3aEYDkT4c3KszGU9VT8BBZ81hmaA7AnL01idomLnVOIA63Hp
Smf3F3CgCbF3pDTHUJYaL5D+bI3x2hUlYtwgnUkvi3hxG42cO6c8HCe6YeOoWm3A5WQxIXLhiz87
LeNpN1mJw/IA0vBb6iMaJMkOx+TbQ9beBAMvLauf1vh0JXQxyEMWZKnwGTrZVjVLGJiaVoqbQf1l
ziXsh0FEmCD1fudUJvKMHmvZSQRoBprgfO70tj6J57HnWyY4KYcdk5IkO9GtLo9dCxujaKFcjOEg
beXyjlAabzUg4bKcuEkIEYNbJIOjKfEy1ouZRE4/Lh0NWzqhWgupAUhBQrbfCuRPNcxZCDmWb7Jc
Y1Zngn3x5FtMYZYapcs+c9SUGXF9juJBymnWYfBvAK1l7xpHDJY/esJknRLq5HgG6ABUF0/7zWgO
bgS2eh55JavBsAVmewEZCGEtvQndEBQ664t8h9TbJIb+RqGidBgifU0fHc/oRibPE9YV02ht1sT1
I711pBw8TSxtteodcIlaoOGr+rrR5os3KmWafo1SLKKMvTBDCZlMM6+iSUnH3NvcVOGZVpcog0Ct
p4hG2/9QqT1HIbTWGZm/0BGzz3XZ9gyyl7D8UJi7ds/TrNElhy4xQXF1+XxXKtGb6XO2RbDKsaGg
7EUmOnK2nyb3Z+Ug7ToAb/6LunjqwGe2CvLk+ASeV2M+ZBbQjZmZ5TYcoXA85ow9+J1epScWLd9Q
7xR9ughCMpx66lxKzznCG6rAipIo/pNWxXOoDH0N//V3QCqP5IjwXIdoxW3ZL65/wM1gzNGdw0Ps
KbIOZZvjhUBPOjo6Iluf2ejPCXU8w9aFreoj9mT83Yj6qbqaHjVPRyQP/10/knj5DnNMk42IaHvW
6fJeTNyYKx1IwfLwGpguv4lXitMvmDgURVj7WbeJidOAeJZ60QTyUdyfRv4/XW26ss6NmcDOCyfa
UvxljHArtb4GeRQwEOLkQbsGEc0SQBu71P9Q40PtQ25v9pJ7uppytEI4Cd+HPFcQpoiZWsi1p4Ll
PltyF7UtAIv4DJ6LHKbfbw5g6V8CfI2PC1BeE9VC7ZvaRhr3nsLHqYKmKZxiEG9rsth2u/wjt8t5
/4SyHzgd3JhNQ3r8EhvP9k7TgxBi+ldXqZMy4VL4GObfQ5kYQsaV1YThrTPnF3HQNDksLAajnyaK
MPplPD2FAV3CgyOm+/xm0Qd0rw71gmJHpY4t5kvIkseC+OSvxJBpUXSZXeEktHuHKtIeQE/Q3XxZ
bgNc6gu2KwH0fQbwTvUIGG6ofKc1lNgXjZSNKPKYfSREDIC2aqEPDyZ0DOyjIbysaG1mlyfeSGAh
RtccEaG7RBBHOVFroNR+Y17LovWgQZzk4g7Uib9A8FfNzktWfTsyTaV/1CMyPuCxT5vNpL46HCiz
F0BVH3frv+NuKjja5IRP+t49UMKkSBYJjLBCEkmpO7KOLDeYaWZGuq4fE8H1BXM9N/jewE/qD+/O
vad+Q0ibaKEpYoZahLyFrN7VDWeKB/zfeBVdfJuR871Nrkp7A2HxLQVDtNOFcwxtZQ/DNFcHtc9K
fIHI0kYNyLDpj9Qww+o7bzmjYpL6I7Xo4rbELFAGwSXEgvwQLAkZD9CFP2gI9k+pgz4Xn+Xn6bAg
HQLzmQHx0YNRDzfrpxY0pskFoh5ju2RyNm7G1yiTVRclccXkX0ZUBr3tkVaZ8aAVJwOQXV71xuDY
SL6A2mVR6WZLP+pcy2xP7Iy4ujffC0QbaFiGLsoq1nyM3Sz4WC11ChRmvGa8w7zaTXj1MA7GIq7e
/IVgtdRb20flwQq6IY5MdY6CChZ/JcMORhnZjUYgo975qvQpa9U3qX2dpgYRC/yWh75IHqBG+CYU
XUG9uz+sxyU54QXjUZ5L1LajbryMeP4rE/mjCLMZGEgWndbepMPaFcK8b/WYe23FvB/Jsv7AmTzs
Irs7yigO1Z6JS5KkErOtOK0mkdLii7D0ebIRd8w7tSdh6U6zOw+m9owa0yZvoPkqUWkXArXQMW6A
0+pg7xGbU6f1JkogDU+DjUyhtIpdtjoZDUNBR7adaP32ZkO1R8TVQO/AEyqXv4GBcFBNghpEHSpl
gP4eaLo0EhcadkDqmAYwXkB9he7HOviCyBRblWbMAAsDC2b1MhY5ePBAMwLDGcGzq0cphOAwjpWA
gI5/n336xOI2LqRnSZ17cg4uKd7cZVvcAEBnze4bjKQqA8LpBlVrAq57i/LFjwFdL2F+SHm42vLH
p1+StcyxrA5x6a+71Z9BhsUltltMiWuaFYUahmjwmq8JGFSNBnEg8SIRMOXexDO62ec3WqQnP59d
y9rgBu2D0rpqE3cF+CogmvOgJsOYaDw6Bw6oiELqmzWAnSzca/WP3oOpIzUY/pPis+kmUe7kQvq9
9MPpcRp0M1oq/bCheyAuWRYmNAfVkp9zWEHuPEtVGAXvfkDdEzXocVr+ueluormuzDydS/SaevPi
NyGUJQis00rvMpDjpXluZMWmdHvZXQMmAbhMbjVEdWSHliv78Q+2KYcMAMyUICphXDhcCbcUzw16
1adI1KwaHKYlpjPidJPYbhAyslnnnVdPK5I84MJs1YoPytf5Cos4/prH24V0bkxT643xIW4UgJgy
8rpza3EdsTNFxOcFuE8VdNImrdISdmdcPF44C6oWmT6AGbLPbjth2qEuCZP2GK/wYdf3AkvVvIc+
22H44tqXsLgBLWNP0SIVjlOK9Ruhmz3hs/Sg8VhR6wsyC5paGSAYdvs7qTqAHN76siS40tPkfPAD
Nmox+5V14wshvOlxJkjFnp6nFBa+cmfE0bE1Zn2w1g56DdhsYZPfsPsa+LZvF7c7BXfgDvOMeE/t
wA2MtAPAd+C0igan4uTqAIId0gKOgL+NYLwblQq5mEd1fZteOLMcuXEauu+8WcrHJsp7x9dFaKHX
xIMcgoIxCLVvmlOHeotUcwivB7tTcQWHjJtCctC+HFdUyO/ROtBa9roxMPYAHq2MchgJWtCGq4LX
vPOirVkbTJUrFnmxPEuTht3pZpDZ9rSdAkoosj4RzFWjauZhdAx/LjhTvl/kdqpEwkGG+Il8voUl
xDhrFu4ZKQp8vsg2PzhIIDWIk6mKDQDSeJxRtcl9QJlJpx7oVYjBW4bYJgNng9frnFSqCEH/Zlfv
nJnTAL2ayfmHl8Dn/jqeBZ8PirNwccBre01w3VCylafVKREMJOOSbXk4M3RaLWoeu+F85xptuysu
xEQ6iqfElpfnIehDdKs35siM95JoX3ZcyKjC8b40rgJT9Xs0Nhs7S3LPe0St/9Zj1WhBi4clnevs
sRY3tLZAyapw/ugaL0J9olh97MwjXuXELyaqdw81vIrr86CLJgX1NJsJo+hTzWSoy+9zxhg2Pg8L
KtdenJCJA1FlCLjMhS6A0dw4t3IbBT1pn/YHDRGPEUH6rXh1vW5CyubM4LWVtOn8BAHFt24PjOuW
B+IybtBOo2FWyC8SlfayeYxtN7gQasyMYWXF+2nX2Nl08vAyelgENSnM5nMSS4RXKeAlVsToindi
ryR+vPRlgFvUZP9l3V3M2Gph57s0oL0ONbC0s3CRs+kpXXZjcHm8D320HWSKDQ02CMOxLKMI6/IB
IAfDslR6qXbDCkguHbQbCX1BnNZiWnBjvFVl4ft5fdVkyY1vwoT2s9ughAFcK/i54UKKje5sxsbg
8g7mHxwiF+qBEun5ZEgU0EOwp0Kp0KiaCD3xJMtCkGaEH0ognm4zpBLrlm+MjXGKbGV0nqDUPJ7l
98/9ehzsJi7rT70QSiZnPt4laKJJrOVT9KJlUvYkEto+3eo5XNKS2POXRaMubHK3WuBtM5SCgGPM
tyrR/t+tPmJqoJaAGk7G8KIA/HF7XiNp6f75NAgT8W/rLkL1Eqn3P70JhkzafoMujLwOH3T1cdMt
0gA9wteXBNCljMNhzWofcBbwcBEnY0FKVwWwvafyMHQicfauP+nGhU8mvWXfERP4Hpr7upEiWsHa
J1EFXZx7rhn9huMHKm/iyuG5mSTa1arF+kroQsy8HGNH+imtnbyBDaBF89nzyk8fqgqWwlnhtk8g
ikURr3N0JrnJ8ae3jFnOiNEOj1ntEc6cYEnSbl2+1aX1qX3Uf3UqrEFcA7wcUvborBjTkYn2cunx
meTZbnQE17BJ3xgQu2amSKH3NW3MSH9GayB0fQOI7gTsuB3vYliuSMNLKxnAxBR4UAekBNZmI1zO
IY3uP8IJRtQHIuncf25rBuY57yx1deZ8UVyiy4Xaj4p5xotrX4j2bPjwzSylS6Mt74GKwOn1yYDQ
qEdqWJqNUMln9iU6yStiHhOXpoK0vr4nMitgLRgApLXgY+qCJPhfhVT5kIwNVvp8t68w63x2VD2a
8Sq5xXQttVIbJGR9NigEjtULtr/kYccoFgfiiJ28crQl2LWny1iiZTrAJSA4lVHyjx7na1jqb40m
ibmt0CPFFTZ5Vsynm3/noVRIDPvQG0Ehx3moMjW9m8Wg3v/BXu1+HFPFYwMIY98kncnmNyDV5eg2
N70iOpvjV9Ifgx9rx6jnEMJDP6O2AwolNxQxuLpJ7H9/oPmDbEG8yzRqG7xofZ3TvANcbHM2GCEq
DoVtIwEDNdz9UR0YidyhDUUWSrPnnWtD/R4xOKLd/CQVmkoMfJ/IBAKGeAXytF1QjvNkrnvqy+HQ
4VkLnXmspgAkK99fsXyPselzfw7tdw2tvb2SjXiDm/v5tf80xxLIS1xnR1JfkhoRyX0Qdms+Z4bv
kz4iq6pEm+vnpyQAlSWAastKRzZHJSmyaTMYVGrS57Bl9SQt+q+o0YLvd2edbWHOhLV0zH4Ycydo
kZVesMm+wppsLwG2E5nZF7duOCNUBsAS9Y9yjWaynohtGT4//KgrLKZMndanc217b02W//K2oBMo
AJLQpt0dXLvqf9+I/w2jWeM2tXO2Njc8JzXQv3jt5PW+ESnFWwTBSaOBwWaLc1mSQQe4sWK2wGw0
/8cpuLubfMJK28OzsZHSTOtDPOsT5PKkrhgysl81YnkCdVoOKXAtbGG5vzgVvs62Vmb/qZoyxeR3
zZmhuSnUD61QZpSaPdg/InpemSykNRbKBWsqvihp6+yeAfZ23m1Y961jOhc5q2FPW3DkEa2EXI38
34tRvvRHl6iHjtCg2ezG5s6suq7d4dgTs8tFS+RNuU82lLpdb+2MRlabgRlKNDtbKQ1kGlXZ70gz
tYxoJYcbyCKH9uY75Z3zGGSYgwTV5vNcfHsk8zmij3vPK9021/Ft+/um7vfazfGQEJqzXOEICTer
8J41OIkjz+HNb2nL4ux10zWnGT3Aw/mYrC3HuhR88GKwd6ql4Q0o6OHGZE42snzwl/8XtL8So2DX
LCvnxlfp+gMigeMWRM2+r4ZGGjFTeLrSQcpbGudGZEGqQnaHSVxh6vn037jqDy3jDmbK7dxNRvw0
+Eqj0j+bvJ9KxEwwFfYqTBAswohHhDsEDVZC1561dkZ+V13f+sVq/+qgL9dx5/GuTN7RTujpVnMa
HlPHwyg6NM0kpttYFHJxCsrTc8t11R+MiX0CZuNDqH3URJfC5TZwzuNDJnw8P8Yx3elOJxi6zYM4
W+lUS9wS+DmnhjaEtSYhB1BWW/V1KcWQi3TXtzGuEl5GgF6CYiW4q2Fh8PVzHCnrK0+a43mm2B9X
dIpRuCMNLBx8t2MfLt/b32Ufl/XlE3JRsw4X6gvkvkqZs3mnAT0WN7uuZFmYg1WncOgcFuggDHyk
TOIvSAq7lpjOc5GrYTE6GyR3hiSxLJ2X97xb5qn+Fw7RkO6uSad9K3U3Q2miKpin9o1V9CdQyjCE
i+5aoVOcIL9I36aG033QMa8zGG3nGLwE5WGEBnN2SuXJ7OjHTH1lETYICtW+J6OGEn+skZ8zqt/P
wOr9hn43HoOIiTcZ5m+VjJc7gqSZjPZ5zQ0cKbqcdRGsGkagL7U4oTLvWGmZLOq1LeRXsrURUbV8
gW9c655gU+Ak794OsOkoWDKxsg60Mfpqe/FFke59Cs1QV9iG1GvtiAN8sBDw0cZJNf1wU7x7cJed
LhRqVq0D6gg3gaywZu6mEIotJ18/N6yBtzUU+JDKMkIIe712Y1EEu7MAt/UY6MAE58Wzl5nId/1r
zcAIPztYnurHPkT5UFiOT2o9f/rbTG48Df0x5lIPiWF9w3QA6rVr2szy25K68pDPIw7JgsDNz1jN
F98MtG9FjansbmmAfiVsMDaUHkKYUO90UprlHoSzaSu9wudr70lb0Fcvu6I3F275UfO+hUUzsw/s
TNenwem8CJQ2Si6DxBlYMF6sQA8AOghHgisoS+ozuyqTx0464CzNGjSoUzPTjHq/QTmCwrJP/wVC
tP+F8bObl03dia4BYPEY9jaxvQ9CGA+mnxxlVcJYQRT3uwxoeKbYc52igluJQmGtxGriFuI/CITd
4L27o0zz4zOdKTqL9s9OuDWWH+cBpVOs/VDsvCD6Wtg/KKY/7AQLfucDgtvN0Scp5wRgLnFDHove
HCGP76yEGy/JNY9MHelUTMkga1Efgj4QzAeCnpQ8e0U4ADbMKYYBKcUVa24iCYRXMxeRh49kdw26
D5mD5BSvh5qbsns86n+2n5CD5QVzgh7/XKGPFIpXeqR7fIgYeLaUmbp9NueAvzQtgBvii03rfc1Q
2y0xMix8A3z4P2a5fd1HL9GnQu9vXt0m9ar7iGgtptFv2BeYgkVFMJ/YZ0RoagZem/YQMV8ktWka
K6TmbDZaj9Lyrq3UnTPNlG94jMHFpcn3//lG/7JvvF6XLuekZO8YH50yc4PDHcT37l5nHP2vEr0z
ZlyQ6H14sWFWl26XTDB+0dx+4ZRAIJ/G+vIG4gW9UMRhwjL05c1mrIza69vPYD9flymtEWlTLWPs
m0q5pKFvaq5E+bmAYbISZJSRvTozR8U8JDAOv5U/J+9xSZlSfOuJcwWZUbnIWKl1Do45fA/u0Iv+
nZjWe8SVVUtTU8+Bmectvo+qBrSHbDBX31VQL/6PiBBUQ0su1uGoVi14kpsKW97yn/F7y3OD0Icm
7dYfuSziWChnPIcXdSyovYqolUf4fdrw56qV3P8FNKelthKaA6tTt+YOyyO/VzfsbXyOot5WBYXX
Y8NzwkKNNz2c6GS5v4m2ySPjFgssB8fy4LXMZkCQJpTUFyRbVTJxLNm0QFr1+rrBF3Ds8BPYm6+1
15OKcJwgmHnRNjVONScvt9VgBdkHwaAnFIRyaWK5DS8Fimx5CsuAPqmg8i9MJB2wvHkhlqgKwC54
VwKqNG71i3obowmNVZMTXLc+7Muwy8uxak0FQiXZKquse62Tm8EaKeyhAHOzJtCCMRY6kEKIJTVD
fSdKHLDxvDWIAqRiLMOEqSiStQHpc+oks+kVjqyjStinXezEQx3bsalREUDBUWFB9pIajLloh/Lp
/Yn8bLfVXrfCtg8hQP35uhbfyhqTCKrq97FALSNwss3iZ1sf+heluMxIYTPFiZxVJQKL6eBr+Lgy
/aN43FRibBR5aLieZ7NFc5icAef85R6dmEyBhgS4HrNasd+RQBegNz2qhkxEeX3gJ7hfRNzTe1QQ
udY9IArsjSYTifhWgQNrw/Qs1aEaua9p9naEPR0zqaBjElu6KdlXDhooUMURpFiLSXv3tLSN2MqR
/4X0fNDapjJtpBypKamjgBzqYgTjKXGRB1G9Ckf8HbeKXHvSMe8Zu7mpP3hWyA+URIFiw4uEYHB8
1b6wOVmUx8kv9hqu05PSE2nx5/CDoQMJsPLCk4TEwC2DztsvRAIamga/hxEuRU7uGbNzFZBYKucR
0S41Qcpjjcv2mm0OsHJhfG7jdbs6szJ+GJubiwt63iVRVXAVZTv3r17Brz5ao+6KvVZeODY1eljB
MbwLSY+AXL7IJ5HiOynU3FjsQRpvoLb0zh6xixdYMvoSQ7dkwJjVKQju7qZDbOHa0VY1kWoVv+o0
LtoLPviQb6Q77RnUCRMKUnmBY8MkiPex+tbr5SGv7DsN8AP0xONbxf0vR/r9ArzLnMGjjN80QavA
Su72sqOjsZ4Dh70xtJ/xO+C/Gnaau8AoRSkRViCjnclQofTtcm7//oWu4XYyRm1FJDvcHPg8NGYP
9wWY4yo/QNa86mtBAnQVmuP6ep2By3o+10p8c+QqiP6Kcf9Ptc8l8ZcGpAulqLSIL5PL70yRKjD5
HQGn33DvVeCO0IMGGDE0IirWcEExAsEJeHV+QHpKXkE/rJODskZXm2M+ZTeYSfG/rxE6hQ/ZLL7k
24gBes1B6x3s86Tn7bz6QVcTQ9zDKwURu+FrJy0IObh7ge3md1NaWe3xWXyjCtu95OXQUsFTljE7
vAKFWZHUGF5aCsd2ZTnQWSaqkGTTGQGuqSUm/p33I73hboX+I3pj4b0M8RgiQ1YVvdVIv3ym1M9r
jOuK7AA6tN1N3PlaKBx549QgLMW/G2uSMlsfLb1JqPb7FPkh8/OBB/IPIOpAibjHiy9I4APKinvd
g1ac6ziE830oNX2tJjGurTow4AFbmVqQbaPtKR0KjtlBj+2Pi+2Gw4rQZhWJBXqCnpzQ4fxgQzp0
69uqAlXNn+OJ3PzotrGl6hOa8L0NrKuwz241ufre4Rs7JXMF9v1WsXOOYZ7E2DyjQTvTWjnzYCFw
qxLRExvnLZnyeMbhB3//GHksfQd/ydF10IJj0ZiX6EkZVBFX39HtannzNWDNk15SS0U7CHJRPYWq
VN+zNV89dKlwgHoNctvOv7cNBS1R10GcxSLgZ4p+umBElotovlan5/20TWOA3wIeb0Tpea4zomR2
5tAHb9JOIwLsXuQzdN3Tj8OV8X+4vbFOdHISQCwXc1qraq0a4USuErGM9aBkec+f4RpMsTg+CY1d
dHAZfcYKe3UMCDF0C2lvcT3GxQUuBbUnpx7bUcauINqTjJL0U1Y5IRbKnUyXWg0UJz4KCxsKYRZk
sJw2lA3a44DfCMskECmACGgt3jT6SfbU0chtp7UnNpUi/I7KdfM/NLBJirJo0cQfmL4buZTf3Luh
4cO1fNPMreH0nLmtML/UUJGNCUlCeXz0epQ8hQrore8wJvJaeLrw7urt7ATMA8R1MXg/48NjVCYu
RUljp1afcoe3RfHQgje4MaGQLegnEsF+3uSQV1hDrMaeTi/gYni3v9lQyLi6BhVqXpUshPn8owKz
JXPM9QqRfjLh33rrrbgR6/06LO3EPwwF0IcPfeXzuASfTmvdQ655VCzqRpjoRe1CRceHhRhy5SP0
xgCBPDHy6ALkKw25jJL+Pz7TQlyifw5TSoSsMd7OnW6KUZssIogHRfef9UdhmQE4gzjRwZHD7x8l
nYurBrgkP0nzjar4rs5wNfFRx2svkzJ5ztJIiKIuthYrrZ6oPV3VQChQIz+w/U+Fq7Fo1gVdN+q2
xmFNeglUxdLIqcDtwnBY1pg+PIJIDdJwMryoUHa6SJJJNemPBLpB4q6cyHluBcMzB52yL4U9neWq
QduJ6mdnqUHu+xeQ/4HJTDsWqrpXCSWpycR/EG9LoqL7Z4tzC5KWNu4xkaWZ1aWm0F54Y3kHCa5o
yugvuP47gqOI+Pbg1cBZkIbOUpwGKfpuPMIaF+EWRQH/+crFna7j7FPDE4EgXl4B+JuLZQY/qqi/
MAmcX52r+b8yGhwOQhlFut0PIy/6Qx494y1GphuyejdL8UoKLMLAvsJARVwnmGFXpAjKXzTf6SYk
//p/ltMJNKnaBAutfL4Ks/A7RrvHCZftXubZ8GeJz6RMUifYwFGUSmH9GcyZvi8ae/tXQT+HR1kl
YBN3bFKwWIEZApv/7gj9afZm4I4LESjJDfznlMXiHsEhl+0r0hEjQArIWGFrLKP1jArChM4hqCx0
jZCZbqES3Ck4X63ZWBEMDw+Z22j/HMDBE9sHAzejwzLxm/tvQtFyfRqIxG0tRm0JyGCQOKw37DOA
8znnxfmjOzwWHV+ybPXa1kpYBBiO4gN91c3o3JIw2ULp/vMttj+GslJZoKILHH6G3Eydp9bDHMOX
yqsWf+7NUt7Rj+Q+cDDEDfUignpx+88aukZZunG9Q2i5ZP/4IQHgSHHSLfXU7jYmuot/TDJ50m4y
qx4DVhNIUC6atK/3b38rFCirydLHDJC8brIMAGr1SJpIpb9FpSDogc2RwJZLJgVwJxCIh6nJhAU3
QXwqRQajq2othb/u2mhgpAoZLhG44a3JoOhQSXB2yrCF4ynGTzt5rBvX3bmkRMZSgNZgnxMe8HfJ
HitnL0vUEb5my7VA2clftJdQ5S4WNahxNObXvA9IdZQsQVSBhwYTZ5416CR30ePIxr279u3rwp1d
M6Kk2ttllppQc1SKBmC/DQjjfKRGUWxINsJw20rHcVH+LJPbvP0eEgFKK+69X4GCa9pk2TYXf+PC
BofeSR2AKFGdycnMjRvYuwCMpsNm6osfQ8C6IobqMRR0GNOXmP4Oj30IXXacdqObtuR8iO2iwo6V
RU6Yo3ghRzyt/M3fVpq8sLYOadIXmYIZgCN70r063N2eyzNi4e/n9qLO3SB/hm7mGWBcMtd8YVMc
vvKaOHu8WyDedpaaK/OAScPGq9R479AugySNCa7GDU6j0bfWWTvfe6Xc/hds3GOU1Q39Fr0DaWZQ
O9FAmjKO02QZ1nmQnaE+ZHv3um6RhU5IzPLRkj4ThaY7Pnoz3QuHpWqyUPC1lwnLeuwSPvk3qsZV
Q5ijWl9x3Qyotr1Bf1UgibCA3M3+TnjHjNhR7lAt1HrG4eelhSb/XjcIXyVfvvmiLu/7+FLnPl5K
C1JpAFPxUHHyJWnYVz6HCtAMXXaceQTCXPM01Khpwj7Qxg4K/jQrJ5pBRD3pm28LxEx0zZNQjrQg
Ob+6mlW3oGg95RjXHvL+vz+fTBb1Qex4OjsPIuNK0XcNdfifn0z99k2RqGqac9qhAmfzCPXbjg1y
ivWAdObZh3ADD+ulh6m/pyBWeT13M+Sy7n3DC88TlQShUW1lnacblgDvUgTJWzGXZQSDUp71hAaK
dlnYSeFtsFjmX5zZFibZGrLXc4PDxa1xHByAYC0z7PetgDbqLKe/fhyao/AUpUSUuLKoHzt3328p
3ssfMF7e8qYCW01qXxT+idDOALv1RYNosa9Tu9BsO1sA0q1U7X3PglfYwPJu0fmmSIMm+6ioZBCQ
WgkPVzojd+gKymiiuiH0GOPXo5OCKSsby7NY6X+mg+dGxcomzsiKOIRx1GxMqS+lOZQx1CVyi+a9
gsXuESAO7oVnfbNPYO38kvxHD0zySPSUzQ37dDWDWm6irGWVkheizESTAsm3i2Y7BtAGwyepGRlv
4ZNoFhfpJ86BOenDmacoMfFv27EoqMT0coSNEysOMy+e4Wqjzj8QZCOn6wh5cIjxwtruGEr5t3yy
yrlM0WX5SxiIu/fybglpryVAMOzuAoESmFuM4UEw8B74zjUEW+9mEX5cD7tdtcO1ih/zOI/EqLdW
8WLz0NePczGbhRuB6u1AH4FOIRV4RqB5iOYBUyEM6uzVlUyYla6Yrkj9TKCdKe/7kvrw9AUc/BKO
8/aPSXY/dFEUIq9LxAP3qrdTyCUz+AAlVHOneb8cGMnYeMdQqHPPUdoxLmOV8JU9NcVYblbnPZXl
z6loxJ9f3FPlMGdb61+G0LAE9/ybHRSFgbHpa6vmerQ6ZZizuNySe4PJcruQmU25cEhQyPRYSiif
c3ZUAiylwLU14d4gT0jgyTotk6r+jk6QPCvbv1UGA7nxE/2kAfjObuKUVSfxAUvr+3vWB1tih0Gq
DRW109+3p5h6q2/tBNbXFBeB3ja7lwwr+i1cr0lTAaqqxJtFRh9GcDh/APjN3Wdey7YR2b5eY8IO
NzWRRxOH9M5aVd5bfWhhp1YZ3khyeVk/tGtdhPo338gnWkfGu6hHENC6ryRAfLb5rf4uP+JMPZtq
/yWVOjy0KZSa3fQJ7q7jX7WGYQ/O4khj6xISg4AESxRt7ARwPO8fAwcaWD/lbN86rMEFp4PLXh4q
z5w3NIpAwqsagOd/CMr8mRqDx/Kjr5WB9xRAqQB0EuTSurkiQGGHdOgHiw1sXuYNimati0JwHwbO
9Nt9IWR99acI3XJQv/IfiAm5/GfLEhM5k9ni9yZ2EX9zaH8afxYsjoVcglnDzoc8LOmerztrfXvi
u57JqCFPsIpv8hlf3Ohb0OEftAapH6K4eK02adF8SnXzFOrfUap5zW/OB0F6K1GcQucUjFH6TufV
S+OvU3JOpZa5hu5YRGOFLE9sPkdCEzKo4bZNvQdOEqlm1acw2hKcw3+eLzP2XD7ueRR70uKqd/41
CzehjyrZrwyplZ22+akKw/1ahfkTyFZnN7PkTqM7+fumbN9xGiAK7sBJBw/0E1znWhJ4uDVSGiAv
KFrd7TGbFYGU7csuhTLC7gPPq6H7IBUWXYs50vJb7UwsGHJ9FODhhPBupdTJJseMjLxzDL04Guwl
TdzMixFfjBrDrT0O5b2Gs2B/M92KAFGIViqv3eyM4WKTYp8tkquknOydJl4KpZ1tyNAq69q2153B
HoMIj/MiULDT3v9RqaS/0BSBjp38nWoq2MUh9qdcL8ClB9pQ+hhV0KsFI/rMSWFT/ccp1ocbaCkK
oI7oeDADWuqb3EO+/zuHaXPBbMor4oosJjo0Iw2w5KCvoSzgO2k1tyvQ07TuE9fpv4TyZT7EfKqU
7W9y95a8hXu+9cdM+MgcMrYOSPMN9tWhXJaIN57u94VZNVkaiysEmGicka5BShQ/LvZLm7ko382G
n1OH0TuIQzLFwIOOF42I5lXwjXjRm2kufKMHOcSGtBMh33WTnqowuZnvPC4Nb0DNfD3pnE3SoMzk
ghPYv91Ot1aVgjMwLa3rdu+SEh0t0IbBXS5h9BUDnK4c9cdoHgLDeo2Umzq0MKAMz2ZIHp5zQIob
zU0LXxWc9dsRtWb7W0LCb/PfKf5gDLkv+wFb09yBYBDOPFBD8bmw5+Iyouna1i7dT3sW8WXswyf4
gvhy0iavOLbw8OFr/t/LSgsuXD7LW6RKPFQO5qlqoWDeesWBig7Jsa1FKCwUlX2N25PXJDJbYyAr
zAyJW1d+eUjefsBn3NRHhbWVHhT3cUfaXg2pUpAwvhYVs77A12uI19BUi+KLSCdQt17EzD0EWANs
To4pq70rELfMIa5Bv/aJWVG2OIpBK3TvgikPsQfPYjaXdox5tKxQE4T8vPRu5lcqH/7Eh6f70Bxb
SfE+82E2smIUEmMll2MObAhNBtOO7rPJQryzJ0IMSkn6XZXgLt7tQ7OX9aZcz+xHWPZED0FAWjxZ
/QRyXvecO0mcqJcqGNGejlJ/0CAPYCRLDvRWSft+9qlKw0oYo48knb5W+jyzdQCuyoqTuxpkgLbM
caB6rxyrjPiq0DiiWb7v6Mgip31eBlI4k8dMR1GsfRkdGVyjvuBpqiXMsqhUlo0qtC880R6RKeMz
TdxSN4m7bNVy8laDXYSzp1waAsoVTTQJMnCrNimrfx8OMVQPOUSTa7B1vcCJS5lp+/erjjkxVDIf
Anv9bkEZA8ao41io5XZUA5L0QVUBKbCq7nI0gKLrDjUdxQkQgZluX1zLx618OF/oz/QPK5gFtGU0
nLeJH5f1bKxxx/AqeECsAWV+0MMi7x0vRJOxlo49MW2x2drB51h/jOgWspxZ1geXzKJev660PF3m
Vkg0e62FS3lJWKv/pEVpOs29X+LInes1Cl8wZbiUcNfaJKE5+7FleaPb/rwNAA7vqUn8RXdtFjUT
MmuS358PdQjJs2T/qzl60lLtJnR6itS53+1J3867pwqqjVAC809TgUD3jq7y1XLGs2EhKsmIkhxS
Z7c0DZ4wqugTIkybQ5N0gyaOdSfVEmIenHccJq56v1XAaS4lH68Zaw8jWiuwPByC3zeITBo0vcGu
P+vvmEdJnxJXuAiTRa6DtzlJe9HfNy9fVWv4ogFnT8Qr/CXywoeDEBwOi48GnnGJEoj5Hbcc/B1j
p/pyo2XQ1W0XrgrLsmuxKqmaeeTBm3aS+00uN1BZxCknYrSpi5DYyd05YAcTvtm0Wt4Ppkier4X1
QDxfT1MOj7dCLP3IKMuMjGrdqbGvQh8Jf0hpUxAfTpPyFyzrc9DK1IRC3QeXjh5smZYeXm/QMPFY
7URYHFJB8Vn8/UuEqxxCyuz//KZN9rh/801xNhbEGWfbs5hcZsgLUtxFCRjLnm6vJV87gVnEfK6d
Nn4cfjqEGsEPOE7VlFVNI8Zu543BomnnKW7vQwpuESUo+sP7vGciyxH4j5/Is25hIO1WL9Fw71Cw
zcfsayzNIJeRz0t6TFhO9y/y/oZzTtAbf5WG1NC0TP23HrFie3iV4I+0WY0pCm68b/XfHiGXRyhB
72TygcbPjPbKU8XC4JvVd7twnOV93JEQNMU+7vXJIO0GMHg1I1lI4ymcebZWyT4tQod6tTDHOai+
z6RHbnuaR0DUIgjCktagQ9HYcaeP44uruOhc2RXEowpfzsRQK41p4dEarcjbpQVWMwJT7pAaSeO+
a8//BdjFLTOADrfdkktQSVAZzs5olsblxeyayRERQTQpsImf3/lb7evQmh4BLFgYxwFGWOw+c2XK
60tcRwKasuoThDZW++MJlDsHIxsuFdP94sw+zhSdaSmoe32IrevIhhsLCa/S0beaJEPVegtrQd0y
20tZcrNP8Vi0JdgDWTCpnnyQBHu4vvyeZMYNb1wASRa75mx9qtWMVDq/XZN0khvm/sBrqG2Oj0pr
GoTrCwP/lDzVinGKWxitHtpU7pJQeDWHlGoyVtpQrL8+j//wkj4OPNRDVh0pU/gyAHEUwE8gAGi9
K0x2uXAMStPMc2IYg36SVJ4GToaAgXdy+wIjjUbgeQPuoTCpt3dRfRfZ95G3Dy+WUxb+H7O3c+H/
Im23vf2HzZLvqFGvn077e/yTQnSdWwXTFDUCj9bRhvq3+6lrh9YbBMDoLnBLaM1VnWFIa0AUKxJt
KHUqnzXYHmc98+NY2a7UPdqaVJW0/fqX5bWIYWFLqEjBUuvj44LVtktBkVL3/N1mCV5kCHISuvVN
2fMwuXUSC3OdrQsCrGRUf+QzVCUE3dbtCwYDG1eze7+37qoa2Wc3E9vxIXxQLlF9KLR2qrzDKQZf
arKiGOUpvVH/HMlXBJ5t99sCxEeiPzXPXFEoiUoz3RIJM2o+SkT4U/NDa/OGmo3jNOfY97ncBKhG
bTXdTbdre36LCrjQemf/jfkwAmB//GBlQqlbUmGfUPoZQPTGhRLea4O/kvymZyS7EWANRfxE0/kk
S/tOPAslw3dPT4emXPxsBm2epOQ3EUt+lE+6571lWX8eN6DGYiaK042LBl98CSox4hWI9RkF98iA
oIXBi6NoC6CT3lu1H7iJYlvZ5cPEH9xvYDMKtALSwB/ojjW9XV/hNpMDpSa7Zvmdx8I2mkytRIUG
GmpchJ/ONSCKgaytooj5i6fY5xoZLRAhM11jPC0XmiUXMZe3e5iF9m7EpRMN2WE1WBrVNtpgLvn5
EDpzoBuXttIbXA2/oHIpogegUCnJsF7sCY7CGxtSpZ5h86TZmOT++UJ1+PmGjKZ9LJzh1SWNTLwk
qH4e5LeEE0SWO335d/77AnftilC1JH0sfAiDwaoUkQzcLGek2gvJuyoktC48FVTP76I5ojNMboj+
APln03XCqnwlzymkI1b0OD9wvxDTk/726StQBx1M9kJW1lfX57vMPSsBOgN11tGL2yKJs1k8/5ik
v51weN/Xj5XuUhT0hdebVtrRPEfMO2lC49wWyS5CToXfY02I5JIBjSLRJfxCdtaV9GhRQ2ckcz5o
Oz7KWQ93fQr7aWy28Ax4Hsj9imggrTCHv4N+ZGFvc3PsWj4kEspgXjo/pgekFiiuv6LIkg5ptmdt
4BKsfyFBHAqtleLXNlh6+nxagOxHu5RAm6AjYoFZjxJty0/fYaxKhipA77UKUmcDAtwXVW+09orb
AG5MmlF7JGBy8NrKtMnPPhCiamStEjAjgwf0Ksy+90xUS7Mm4ys4IFAipifCYZC+oLGgoOGPxUvr
W2zC+luWBITxT83HML60sL7X+9oAXUKFMMWTcJL4L9QnbhxBkl2FDFhcRrgk6oEkBlFY/gwrl/Cb
S5tZoSiZ45C+loIGLzJd5oYjmVfYGy37msASEqrjFK/zA9t1dzK6Z8pQCbqzWeqSOYCok0UwWQUQ
vQUu1s+3OK/wF9OIBXgIhEYgZdRFRRW51p4VGJhk3qu+1+Ie9RfmOGEwwmfBP/1UFkMQNdon0L0T
vedwbvoan8GJqGyekFDWXfQBZ1fYFEeFyfHn20NtxqxUAmsdW0Rs0vH8ri0KCRUcgM7x9+RPZhhI
ufpL12OSNiDLL8s/+mljjBCVIuk8xvR91jT23WJNXG7lCRiIoJtGR/oUzrv0RpY3zTN9+rgoy+0N
5ZeKIthvZHbo7twJCXiHUxgEFhHhryajaxy8ZqN8Q9EaePBTCZtu68xhTpIqYemEXt9ImS27u9cy
2hyhZudw2th9N+eYiBZwAskNCQZgGYluRd7DVHyo/633kMG+bVlw9PbqeFZcOeETuexKeQbNN+pf
kVL9jNazAbMvegs4IznBMpTiDwZ5OPXJgSAHrjfzfbnBpCqaRLCQiitHSZK4EhZSd9MQq8lbYIdG
lQwGpBNEZdz0a6M0POFjTSQWDl9c4iU4E0FKEYPMZbuannSyv2MzYe1g5YTwpygALjQONkkbv7oN
lzG8gxGWQEzzZ8BKHPSTQx9uKepmZD5OfeQSRw9+1PYIM4BCuGlZ+mQXg5o4NXJlhqSt43N7x/d/
3nI7wwsnqtgrRh//2FN5z7QVgmPj7UcbPbiCd2jpVWLe/WPXgNxdYkEWTM7vzhOhRvQ3gbHurv2j
gEJRmZ6l0JmnijxeK7CBIMEzZhPJ2tfHDSZfYAkOZ5+Td1UT6stj2shH/7vTm3YwY1UwxZqKe+HB
JFrNJ4PQHvatWoxuNOJHcb8sT53MN2YgHU2r6BeCLSpKo4VBsd+yZdABo0K52nVR0ar76DmpgP2Q
iX5cvFPhKJJ6kzNvY+icUdfLA+nxsiYK4q9BgLPkEQA/ErhJJNfoGKyFNERww+/pY3Ghg2ml2vG3
+bLTGhgD3clLX4XaLq3e8glq5AWkgqemYvRYSgsN0LSz7cvcHoHJawVgzqcddLzVHdksIpahQKqm
L+/lEgnCdaymmxBPRQaWTLCllIqNSzUGeIQssQQmVjFD5/fzgdVUss3bD44UvfmpD1w2u95uVqx1
cxgWzWhbSJE8CJ5imn89BFQSNO7HH6rlpHjls26LUq8EkgSDiCaIpPhG+x6m0WMyswgKV+5RANtE
ySdFHHurg5fToNFpn/OHgONJW7l3Q6bD7h/RePpJE2SWLy9hzzcI+HAdp69cMf8U3HvOLfUhg0YC
z4oG6ftRm8NRJax7Hp1avl367aQUwpemGPEtbyGtbC/4LzVmwcKWPZGfu1z7BAVBjwCz3vl3s6Uj
uL2g5JC9jAa8vhxhuiyZcyfJtUodsZMIA668R1pS5EjbNCo6XvQpAkniXpHDsc6g7wJge6nrvURh
WPdPsi3D3OdyhkL0VzS+Ti6GqDgd4reA2VmkYtxipYgtNudeCPum2sW0HEBLEbv2lkzl3PRGSkqZ
JGDbuSTwXqEXyL0/ESX1Swg6wx/T9OM3DEA8Xie8HBT30dlM4N5BNF3hpJloLT5JGk/bWW1OSCJB
DqFPIKmLnKDZiol8pkve7pYnCAYQtfX72Z6kQp85jbigL/SxFEyx8G0uxqDPa5+Q947AIBRr0qUT
Jmn22E3gmf0OXlOmvZGlsOJG321Ktp1kSRvPLdaJRWXDJf+VQ4HEFYp6ytS0X/n4rHWhUyTW/JxH
Kiqxu7xJOrXqOh/nR1Rvy/jrWXwCr+wGwrnhGhq9G2eGq8PtX/EWQ3/S+tQvb+Sr32NJP69m5Jkq
EQYM3Rfmuax46nN9FHEGQGC8zDfbT3ewsiJIy27OY8COvisoqubVn8PRm9SCsqpEYGF2FEE7AiSU
TplnelxdEjr4XqS3XIhumdy0vng6cyuNHC/4iI48fY5ummRSD96gKMucm3oHUwlaKlb6c4XnNgEx
q9wCKwVqW7oad8rsSYP3rSPfQ0BYwEmGfqocgryLDmM91Ahk2zXXcZE+kK82FKHOt6hg5a4eWEfC
8ihjbKfGxJJnAKfu6ps+l8QtJ07YX7KyXUSAVXQXv/ATRDG11TMcIJK24jkiqwYNmXQAMjTmF4YT
g/6eLrgw8RrTgfLRh4dtV7CEqh3qhjm9H0vkS1BLSi3JybHOFezi8zSfh973Jjqoue2F/xOloATF
UsUEkqDViFs0MzQQWHGr7IhoRyF+fHCuEnTW1zTOg6DmsU5LGAdkQ9gsd4R2Rf2EYZ49KElD6HBg
2UGz2kKP4z7gTjA3luL0flUnKVR0bJzuEaEGPASV2Bb8NyndCo5st7zgtdopIgjC0jSPbkUw0ST6
G4lWqvIu9MaxdGq/DTdTZu7u3GRoC0xlOiyQQjUQwmuX5Qr187qxf+KZiLDYsu5st7gTSK6eQQMa
yQZwuaYLoFCfKVS9AxgN2LkwqoiIwQJgCpyO/8w3YJM2dyY/PJai7eKGiOisK8Mwh0uUktlbGpFe
+nqxZXI5dlU/9L9hofW1lcbXRNUIvpJYhLJmib+U/WfmPsLGRtsribzTddO5G4o8kCy3KhAG6flw
mdgRweGN6Ax6SncnmReYCpgBVeVf0jy4jS8woDmPxGv5FjxjGg40Vv5J94n2PNltxE3c4doiL6SR
CH+ia+bq7XM6wvzRHYpJ3OOq4WN/xh/05AhY/roH0I2F7hhzH1zGb7ERfj0hJ8VcBKOGwyWej0XM
ZE7FFapnSpLPIXAhDLdQ26B/QAi3JFxAmN4gSi/7mAKF2XZbRTXEqFmReBBeDGsqtpjh+aa+vgz5
j9x5m4nD8+2BLhs/KJveSdoVPf7XaxSzlyIbORdVifP4yWtZgkTyp+aT1blBo3RUBRE8hzXYedmH
TOj9hBkkadTgOFCY5KIhTY0T+5bgKyn3n8u4o4exh2A60dHFax3Jq0DsyxDvm9dtp1owEWnsGZa7
47BF2tU1gXaA3cSwuskyOLfYYI/CgQHQkIpSlAu/YHkQTn7utd5rW7o5uFNR/wPm9ZZ/gRQOir5j
ozC4L/8OIhHwklUd7eWNLUGguKLOKcBSpwbK87OuWDR/YsS+BKoiSEW8p9xecPhQ1vouMhWdxDkm
eNBVPeMjFxDa/LUo4+en/NCkhL8+7JRKsAj+NlGQq2g+r/0l792njiW/fBE6Dolo19JPZe88VTFK
47fmYqMSVCBjj4pwnfTyRlPkF6xXgShDm/tk+jCLYbN5k0AgAamy2wtfKISH5SzV50lHs+2Z7lJg
AcypwPVJA/0v8PAZJUgIhyU01/Gc4e8laycBH7GcDqazEn0gI9GihjoVnvKVo1cBYBFoEs1CI9ok
MXp6ZAsbFET9BoV3uCGDOAI/F6CMgJ0fIEFrYnYcUrl4tY8cx7cKdMpWUmoI4xTiL5ntHvQpYJNv
Kaw+dnfi9Hve4l4BrFKojMFvZYImEmIFK8AO36kCF9ifuv/zDM4u8XXh3DQawc6XTtEFPgjGDEi7
czoL+6F869iT2zZJla/qchfW7YLZn5c3lzZ/227L2DuYTSDaqMZg4TsWE0OwaZNitFVUFkLzCNOF
HjATiYxQZrgcWzuEDNSgL72MkX/FEhFS7A6wmSrEVrcsw+t69SeCgTK31Gn+QGiylbuGf4xZfn8Y
uYxE3l7FFzIFOsa7/p0/f1O6tKSO0CRQLQn84bLiijsXoXRB/xz3YTytisURGI7QtkzaygnuAhAK
0oFgICPBBd3QdAn9rQpfn8P5gcxy3XfkbZ6E2osHx7T5lC58KFaWSiD7GyBVCMbDBUWvIqY3qB5N
gIjqUKqIi90WA6RCUPn8QFiacBj3av/Y7LLygud9WHarXcM9xyJml/Y/hiAJUdtZy1YAa9OTEhh/
AjuRCWXhfiMeK4WpswdeHB+tXm6wVxV2sbXqmtT/W6k5mWMTtnuuwhIuaQFhKeJTx5LgpBaMLBOj
3IFo+qLhuZ65umyqVdKOVZ2G+nm7PJaeAaKUuVXYyP7DcKirg1V0MDeAbfMgKkhZMtFUNMzQPWau
X4fz6AfJQxwTgw8D5quqTtM26uoFg1QVvsQ8ECn40wbFb1U8gJZbRawhyJAkWZ17nzOSlXyqbAYB
co2/Ekp+jJycHwlTP/2Gmg8o85jAz8/d+Y62XJk0VdU1jfS4EuIZe9OvkCpo6z0Pt+PAW18cNJPF
lA58DAcQuvxGa/bk01cEEQz/+A0FhwEg55LXOIMvajE5TPP7WngDSM9GHZOddciOM3aaanXDQPgL
Pav95UrEogqIW3wYaWaHDJ3GULm4ew3D3sj/eqx/pmPYf5dABPqlwlZRvkxRrTNvRJkwabwM7M0b
ohBLgNiaKbE79533omTYtDxb77rT++FXF0Zl/9LgkPafXTCa50apzL4/8JFTIL4d3KgHYvo4NhMc
9mA1Sh+nm5guzzvkr8DzlY88JSt8bkd8tbnrhKMxCaF2gYtMWoQQzjLe6JCbP8hGPOY3/be9adMi
TSkzpz8r42TMOK/eb/CyzJ2IxXQVPC4olmLJkny7yvTdEwlRl+YsnS8t17b+PfYWzYZaHVGgfD/A
asRufD8qJJmV4GtNvMhjzgDohuoc0wZwUdZwgWrlthGCVbmmyAGTJk4zPNy5fhfdlk96SoLpcRF9
1fPtzubylwR7uhazY06hz90Rwq8LmTDqo7P64PM4CFMN/9R2L4sK6BKO523sh6DzCj7HACVE3jrq
/ktEal6I5jFXkM4Ef8a/SzqfMQ/IcpFvmyjcnbnDAZeK+IuTl2BEc9aAXuYcrI9u/a+/Hvqw9S+n
qK74f5udo/I8gYzwZeslbIh67GaV2bU3bWGy+kXyvk0s5eZzPgwkw3fKBN4Kqc3+/aGEvdNZJDfg
WpSGDXFrGAGB6X3jmZEYcx6ubj4klauqndSsYb2G+Jv3LIxzKQ4gTDQLKrTsEKeLpJsAtu6ECPpF
uVFYMgOb2vdgiHyLc34LkXyrvtbQhOT1FZ3DJnI0H9EBl5HhuHhnEkQuOyf02pYS1myk39dKMFSW
DD/pUa8CHasXTzFxqL0pGgG2MOvR64Jv5b0d/mwbSt+KpASZPThGXwD3S6wAUXYX8c8M/sC3x6kA
XRRDOtK1VLwcIl2JIlFA91DARQufeZ4VifAA2w9jmgZNj6Di/E+IyU8KqAWGaDfRJwp5izGE11wY
MtyDkDvfoaY3bP1uz9QedIrUj3n/6zz+BqiKDCED3E/IuvS2YGAae0951KJDLh1eDbYsB4PiQFNh
wIGuVc1A3jZWqKAwK2uUK3Ho7HqganKCh8cBcoc+f91epRsU0mGVMyNDA2A6JWyyWzD0WCnWN17N
P3FG3i5bzx8dILEnDcvjxMUQTLK/D8FDmElXgDUr7eZH+tpF7jECH5QkZx5KbBlK7XjFyoQXLylO
Gn5uhwNbmBgGqHgshfQjeFYJtjIpn3/GpUjdigoi9X0uTeFVRw9r2BJCQSWqNHRtxXn7Myf9Ulxs
EnRTHVDaKnsPyQGepIwMHHk4a7KKU4wzCYIPaj2U3fhUovRC8gpTl0At1G6+BwIhD9vz/rIlU0Rv
S/lUFsMrHKNW7XS5vWmpLQzRd/ifa7BDuuRqgwWX9qGOam4axKT4n16lzfgyNL5AggYqkJn4S3Cu
T5xO4tGDWHVOAEU+DyG7Eh72e4xDgIWmC60uqoYaiaaOKUWnmgJSaKkeTqWHJA0F4RrOVR/5xG6+
+uJbcPzwNEFhLpq2domIxYzuIMi90uh5/rgsgJHlAcjWCGovpqde0qIxEWolgW0c5LWHoROpTzdt
XykZAcwjYyeQkzL9+OKuedKyToL6zhFyQAJIsiRuFR/QPxEeBF+ZB83Ti3ohSufTN56Z4VHefKs9
m3RVCHef+YVA2HmymBvvFjVnA3prT4otA2sJi754GZ6D+I2v4CGDPmXRRNZkX/TwxtcqjluU/JPh
MlhR4ODovkTSJ042UGJhveoCL7KZ9XkFrgSiohMzK3+4Xy/HIXJ/siQC2rTF1/XQuN8teA6IPNZt
LWnpa53GN/Z6qjzRndj+QO2mqJITer5+Ywq2e7f4oScQb3gFAvslU/2IApK3b9CejYiixtCZX7/R
TeHhLfHlP61srITdG7CF54Sxz6OUSIElw0sG24bBvk5isSiO8tXUKQOUKATQfvzXshAr6wDUz5J3
yuPaCINd+I2a2WmLo7IjbX0s09n96b4ipbLuz58wZ5zuS3t5b5Z6xQF4mT9+mEO8UwB05UC4qq7n
sfJI9ZK2H+uxLFgnOEBq0uGiZLHkQUQjUYvAlXZMjrrv5x1RBAACIQWp3KQq4wlxwrDpjOZqf/zy
8R8ReG9IH91m8jh/g/5aBGid/f9h04BIcorn3uPZ13aJh+cvVaeQ/Oix5PFJHA4QebZcNkwW+pG8
UsMCNAMgfrePrJcL9hLQPEIi0Jc84tm9PY42P6Y5hfUteTdx/PLz+HjGfy2ijrAnAH658cvX6AFn
togFK8aZ2yD1E06EzpB8KpyrgeV881CVv/5hybKGUSklXqTPRvMpfXGypUefRMh7tOf/epGWHT/a
sIwe1EaW0gC22Y2aX81j/0jSHtBE46vK1p3nEpo6i5MLByXEyPOehcJEWQYHuNxQ0PYilaW7ItOf
0Tsaz9z3V2xl4D3skVLcsI+0RXs0pYcMy1YqLf9TavpuIhAd0iIfWTqREy8B7OYY56F1n1tb+/Y8
aBJgWgENcGT1QtZx03hr9OJNo2MtioI3d/fDhA0x2HsZe96rMRmlHp0mfLbYHplydf/BxYvDdeTh
gVMiSRR2900nAmlpcLKQOQ52Bh6cwI1wYW2oVH60sGCP0zpneuk8a/90y+VFgV32aa23qDUfaJNT
xszkjS1eR3fdef//AKUDffUuHOsYLUMN4lh0wuVZ3GHBtxsOQHvrarTjJV2hMvPO/0DhCkFBhbz4
0kia5Ya+zIhMlqyLkiU338lT4KCyLA60y8f24msDylNHyW5jPnrtcsxX1OcbE92yj9XFExJTu92A
KuKcg7uv3ycMXLF4wJdlHqe00RdMbdFT4Q4jMzG8MzRpS4uTY9wxal9XSt0mfcLo5n0oeB8EAmR+
PJRFcn6JREx3GP+nCTURpO+6jfeGr/wWC6FM6o+yUOoj4B7R234QTGanp5H0UNalnZcYWM0sWblN
qdNZ9hfU1gjaSLLX00wmu3Gr6PgC6Ly/YAirytxzWWGgdtJHQ86jHJ1bnWEHbg+Ly8dvPj+e5D/j
ri0yaOlQdJ4fdbZT+a0sEVzCrFGqtgpIIY/38tMfiqN2KfNQXObfJOn/92UthjJrcZ8ESdJ2RFxE
3FGYJPN/I1Zmrn1nobHKmuqU/Vrz2g2+qrQHMCrwvPK+g1yKjad47FP6Qx6tfM0RSvl8CNYE5pNp
aGuEDwYtK98r0u293w1ud9H3bON5LxVim48RcJGY9jX7IWp4xWfTH9EZ74qqKYCFB2sF4TZw6udR
IiZz5tRAv98aR4tju0qf2zs9zmkwpwRcDPC1k9JDns0VTz93WLtM5X0NIwm178b3S2O1ZNtpTHa4
7Z9vpJhvIhQ7dM9J3MUMmB5HWbMgifxCqp+OIp14pFqXSDo9cLykOr9Ap3NvByxRf6kxdtH0Esc0
gTt8Ti3zGnNHDUR2HkjQzTevBio+bvNZCQ7NyXBjccNU69pMali8FMyINdUJB+OfDhrkXfPyceKK
+8qXwU6kvGKDM/jyNkSDKX6hyMRfMcoqkYKFWZsU7OgEjM8ZCUnApkeQRoAU/MCmo48M0qdaRNzW
BMyU9PVge8wDD+0HP/ayJUWpXBcCwsBRyBPupC3cQiVpbfOPhL+RVpYJhOKF9nVXBh5Kci8G2XCm
gGMHiXCisSddEjSWMPBPLcgYpfukKjj0XwCrzIL414ayZUyzkdI6KxZUacOCNmaOdfSz/GykEQBz
0L+osjDtNqsy2iu4bI6AWk6EhYwZvppy++oR0c8XL3P8z+PT8i0yOVqRWj0FTm4hm0bvRfwd9fZ+
Aikry5NeC0qKbZ81jVmNLD2q1bKIbX/2tgQaoGipYMMFGd0YY5ozwEsc3KICRq5qCyG7DzO8vqdP
F5lTziS9Wl9TvWVZgGfNT8MCZ7ETUYQOCliZoUmhVHs87RbB4gtwjzP7eOblWwn/zJxfc0RzR9dy
XJz14aXEwwYhVVqJ7IhPI2zeCdq7m/bXXTd/7tFyUKihH+WowHPbD7zQ/s3cgH480Is+8n2BL9EE
gz6iNHSOztlyhYdqdFYthIjah5cSiuuGBVk2BwYIEhPJgw8ncv568tE/JoyvPD4B1yZVuoQ9OfRL
rJQ+U1y78V19KHI325uKaSf2PyM4FNsSpXmm4Tasu8LZ97+JObzdD/kO26CqpJ2PKTeLOgB5b1ea
DqQXnnnEX5FVaKdYqatqLvSyEfTRrraFAIuExMGMC1g4y53JyoI0J3SS+78+AWqQFWfkYMVuSb2N
ISUmHJuVaf+OtCE9ptnkRCyC3KU1mu8RV0lTjSfFGrn2WyyGEzZumaDBlu/s85coQaV3rJhMG36n
xPHY2Z9noPBXc7eSPS5hBma1e8IlHSRytz7QlbOApuhZeAUGiWoiQXRviKV6cGljGewapLi7ettN
sjCHu5nTKy+JdtDVPBJ2j8SgDZ0YP+zbVD+Ig5YG6y9QmQ1pJXZrWYGiRLNRBVaKPmX48xY/Wn/K
Pfh9zGjo5lmVSU1tP+26ClGZYRxOzbF2qPLlxjMjxATJxnpKgBYPGL8SImz8Hsn1995C9rNCfk5v
JSBA1WnOA9QKMssVy2+XJDipZLFKEjZuVsfxuWWP3gPDCWN7vhMcyrKJ6SihjymbQtoKhYXVAryK
VkvE3u4BJPCJlu+rn2vSXCF20XjCVPrr1JG0lg/Qh6RncQlfd7XZTwBT/pOW+lEUQ+HmNBY3cIiU
Fkah8qxmfxd5HgscqSy+1rRHTBqKR8/opJIS7Qevsh1OPMBOl4YOz4c7Zdr25Gyhr5vG0Dt8wUZa
kRi8tkBaIwFP1+TazY9+d4+HKG0R7Z8+NK0kx1LJ/mjWLhDn02srqeEY3jnhh39Bp3eGahAhr8gT
eCdT1jKlY3pOdSshM+VbxuffQp8o2WvqqZFZSmwyoNARdmMkTB4waExu0C1f7bafM4j4W0BGsRd0
15kNtdJqi2AfUfRpdxNMAxDSfj3Z7ARMx1xLrxyJbYAyZWdR6HGJ7Pqp42SDLDbe3BxhPDIjkDih
PdHEj5xEkN4kmT14YVyjBNq4BGO0jBEozs5vOOLce3iTHIf8KwyZFtIiVMpGDP+e2JC4XtrreUDR
47utuW9cM+9IASpEe2JjZqBbGEeEzCv43mBkm15cvf3BXQDlkvyMkJKmQ6FqQBf6R/xutB71L0nP
7b00Z3PAc/9o3qbrd+mSK9igJodCPxo4R+AMXH+OioHbkzKBz0Tp2nEb/7dxZJbl+EYnniTsxDRW
FLH9Q80dS1BygoFgAEbJZIKRu5ol3du8+l3LzKAtFMBDnrUJYbbFriLxe20vzRikxMnIzLQ1GrEC
ne3j3dX2vK5ko/oGSX6bBZgu7F26DXr3ec+qD+BsBFZZ8ZNGuAZ54/x8nmXiOTlP1no271tOYsQJ
fGoAsSbkiySCYl+aDZP1jSVxMXY80l4LSdhhax/qwyySy5tEUlO9bBvTQiAmYwRLd6+D2b0/kDIK
qJ41zauAANwQJIEg9f0U2pZkt0b2AGAZqWzTI3mf2nRTDyQYOcQlt69oicrFYfgAOO1CsEzOXjix
zvLF0vYueNxuyPnAR8BK2qJF81NrhKHurrUsd6vt91HDpjopFsJEjXcT4JUdcYmZWZeKW/mGnESD
c5RIArlnfSHnuPmRliQc2qBTvFiJSE4/lbij43J6UdbBz5O/kVE0r4Y2c90TpkCOvVduidCSmX4c
FrKv/9v+59bNtmcADoyYn+/2LuTyqNCWSmeST1hRfvboMYqs0s2ZUyW9z9jtPv5nCgI8G0+nv5mV
BCeo33bIyk3EE8VAV8A3MzI4l8+8S5SFEDFJgKkyYLeMoUPOqQLnfIOPMPop5TAWZRFT7J5w4ZlU
WFkZqESVlGNtnPrpZIjg1FUnlmUWENaaV0v8QcPMFXTSi3xfoNaceUbKBBjf4b02tEfigJBR7TTs
gMXbDFz8/k1xQBswvOZMoyyylaMJMdo2TnDyBqToVnK5UecWfMP4Q5XjRKT/ym7SeLTQueWAxGUN
2PVbG6wF73/VIQF4jh9XkBoLmKSeOz4BEuWd1nYf5FAvGZv5MZsF4cZFc66FxkuMHNHrkr915fob
KZq+zlKbTwQgF43VfeNkFAmt+IgzYuSsK8Ju385UiAgTw27lj4p7+WVZaB+o9JwLjCk/5uA5bb7t
VTdzR76jlrcluM1xlfLqCIwubXf6HAk2QCiYOMMcnJ6RCYThsWDzIUQk3UjS7ONi0kzEKSh24nlH
E+Q9xlvDpRnYefmPbrPRmm3kpuq0H8mbMNQ4GhY41nU5BPL4k/bB0u37nokx+HQZestNnJfEw19L
TpwuAY8rXPS6yWVkEIj4oV2jVGLSFvCnnlgOEy0qcXYZKSJRrMKmVI0JNruZbpQ1Pxhk0F9awHCL
TsQtj/vTC3UBT0umMkt+0lR959+miUm1B2SLWK7Fwnu9WMxkOiem31UCJREdp/mEeIfo2VYfduWY
VKijitwtYoG+ywIKOgqIHaIFrZdpPrnB+k03qbBH3lROm6CRQhg6YQ6IZ9Angu3BG6a7Wmjwdb/a
Tt8zemH1yy4ceh0Wy7c+3IrHawdZLK3Xt8AmOlXqi7yhPcOJm0HWrIXeTbXx6BGqKI9nUAqxBZpN
+dtvauEIEziSijyVKmGuu/wGcelwPItzq/7PTtb+mlW5HeYOUgK8iuV5GUsXP85wQlKO16+X21dD
Jv4+Fo8Exm2Scu2/rh+uoltEqnN6S7clQE3mVwEejcTOLLXmi812U6FFNL48tLiSCWeOhOaPpKC8
FvzuGVzG/jakQ2xakhGRxWZ2R8PfdtVydbhCnsr+69fOurCu+zpISgmsexceGp2fiACODuHJWhtF
JG+dHKGx8ED6l4Ge4oa8PWEYJhJTTt2qL83k+jCuJM8QgC51mO3j7W7drBGZwdx9+U90Hv0Iui3z
3dl2mYR981Hxy6uiNgaOr3PEKNSuBxgVbNXMBGOrQX1paXfsPeDSNT0x0b2NhngQ45Drqr3sET7Q
n2ypQkLMzrwSIA51ZnOUjlfksq99XIFOLMiJXdw0aQto2oXO1R3VPIs18jKelzPTMRQW9eyguot9
D+j0FJwV643QnvneFbYbFxSCT9nDpnd9eaXg31vkMrxArM0LZT+qGYup/RI8Ulz71ca2GPZrVVy6
jUtPKUFI9gUp4TroHMNlMJBxMkIiLOmoWh0lCEAWjzdY8MV+mTa/lvV69MfPIP1s79kg8v3kED3x
vBSQkTA+vxa2iMehdPlRDOhWXcUowTUchG5IMIGVvwlu1DJWR17qpOV6K4IdJnqfgurQeRoPEVtl
qjN7HywDiUCb0nHxN0Fyeg125D4qiMyCV5kzjhxMIWXAx32nD1A8BBrrbCDezJE/7JHkmv3wwpUB
kYIBGR8LCA9Q2+MLhwV+jOLkjB27vbyKv1G1n/11vcCTlN4egtRrli/9M+tI7wDiuRpG2/tyORjU
zq5HNyzlnRyW59uNofzbUeDnUF22APPP3l9SdWAedZM9ToVoFGGZeeGEoYa+1UJZ5QOqHg9MQBgu
XT86DzaqjQjmGi8LgVP54uS0IIhm2f5lr4NBKSxKT4IUSNfXZ3pe2406I/7tThFWwBtSshidaYJB
yldkiUEhfKPK34xiUY8XGz7WamrkCY4yuLCxiDWzDPuvCyHZi50aTQejLtvaDWFIslrL/UgtHUBo
cZen9OamV99KIWWu88ogD19lFmrA2QwIkKSWbkxj9BTrkiDGgBvKwgRh49Lfpk94mGTXtF87ytpB
YzGBB2i522Vuyvki1SiXu1wn4lm5epGhyhv3irF5f/kbyqEoPrYlHzmv698Rbixi65f2avPVQUll
vgRtANt10mcu2gaNRo4/hj/sjbqyiv68YVveE10GthLp5TTOaJXOC6+i/g5VbcnV9bteqr2yuBhk
9Uc3gGR2wPgnaFwJHHpJFBWdDst2BwXWjlVG6J2ICOiOvvanmoI+nsZtAJPNtYAJ/AbnxpvxfNHz
j/UYhQ3YltaG0rnAQaLx95SnTOd/PKl3/CkXJ2LSe5gZY0UQ3chYVSq1Sd0tXlwv8EIbyjFATYrD
ASIirpL4IxGpMXqfhnOupdoaM4iTN72TtCtE+5Yi7xI3/HW4esA1m3bvpqBzT8fySGX05F8Lna88
61rlvBnVLo0/oE+ly+aeHwNN1c/SRpxfrWdAFBy19W7OzQMBaJelHdSMnrwC4/AOlwpWEdOSP8YM
/tN69Gn/wzTURZWkyuNCqDAzOrd+QG8SSKPaT17M5Nn7xmUt6ERKDsioGw5gsW/hGlROip2QCKh9
HYNQjlK41ADIrK1wIM0qZetYmFoky3Ak2O3iiLN9kTrjIrbmQuaQjbNtF5FY+aGjYgBPfhpDy5vG
QqD1A/9u70YvVjM6YH3GYLXKW+JV0giaABIr4ZdzVU/Lm21VveUQBpYV4UCIu0TZIvKYBQUb7w5o
+YztKv/9WS3DdaGOAYw/0K1+r6OLTK8FNZBwuerSJwL94WQUkVpuCLZ2v3beIklYFcXzFoN7qtt7
zigU9+A4X+0QCWnRucD72ZDW8HNMB7a30GOFGdUu9PUPyXKIGm9ili13MzddO5Qq8mf70HXpKmLa
73cRQU+Bmwzh3hguCh9b0TwBT8V5jk2iBRNZgR5kn42G+xoJrz/IVKTQcmrua6Fqw68E50LZS3yI
JF/qNOa/0KgPuvo1d/tU/C6g+D5hYsenflTlFy3zKTzakMInq/aGc/rinnwCQoWgVN7gI545o0yE
/JnVDnyXPgQisgAlxBi//ye2FZ9wwsgcDzI40Tlms+Upg51jDYdf/3R+xwkDHzBncSvsvfO9lryP
orKIG56KNSqhsTlO2tWdKTAcr8JldAGpgfA5AHDPnQ4JzS87/3/Mm+/S4gXXtIncO06VM0sKxN/A
MzUMPsN43azVgDX3fGUyw0WhQHuW3CZCaWZn3xxR4sQXVx4EH7YONxgcx6Ti5POUwhkrdkyWiZ5A
ODGRKxeRvOmgGYYpcBmx5NyfZFvI5Jx+SmmE/VkXQgFF7ZGTZ4U1CCHoIERpt1Z/oKm6SQg8+Jc/
+ztru/DyNBTbZtBT57DmnRlNzWajRsWs6Nz14qYSlqHwwSpDjnJgIJxOKhvMbuYw/Wtio6ih7C6S
ckRZ1gGrp0IP+782Ep9hZuyhBXbyOkruyPjF8e3xix6beLD5LfYebTSBJppnyICJ7qjwzwa8UIYI
SfWH/cZPyYF/QEvZ5Y5+BEmSE01osBfu2rH63NCNgWRwLyo44CtObxqyREnrJQHNljq7oDtnk0gF
LSAB9udCSif598Q3fh6D7AfpD4B2jcnmPx3Q9nD4IPOVroSKLTY5cbCuDmNUTtOl1hMsoqfn3rAp
IdcUubdT21/F/FHeYA0TUBWfiTwUvsOTXKzRUtK+EfXq/OskckhbbVT81GZQhNFEOJzCX/EWbVXV
jCgzBJMdLSSTh5Hb/q4nA5MhmPQsdY4/7uvTvtkCF9O+w5IFuEUsB2GD4AgyxqIa+FDb/sWL5RjF
zM3N8Wj4vurljqbvxuLgt4GouirXNc7TYK/1XQaXTadEvvL/HRIm5fsBvPxV+xQeByNHGt22PXf9
p2G/r6enTRQ3LZtGNtqCcBFK+KBASYY+31w6Hpzr9CC47I6tpgstaMOTcrGmykoglDDnN/XOYgG4
ZOyCR1MXcxeWPJ8r4kNeIdaLfUfpLy/3Y7nmDzIuZS/soHgl9odkf728YptCyDF6cL8DJOvCire8
3vCx5qhhpkYPxnx/GrKtLgTYcOmrNMeMp5s1xST+aV3zrckVZgyeODxIjvgVMyfKBYiA9cRhWqYl
uNqQTZZdAgoL3bAREoLaE4RjmSkn7er9hOnMk7OR0h7czWwFBdto14SiGw7O0faNaWmPq5htk/4c
ROCP6zhaTOlCPAGGZZL9go8Ga/2TDOiMWGTyLHR3Dwsb8afnEJUpUe8gpgYubohx4n6uJ92zYXDS
o/wVRVPtadS6EjCE1jwaHAn5NPWoh6dRIyPRrR8HOMQjj0kEYCq9sOYdetgM8y94b/pOTKZC3bCA
gKE8UUcd8QrwipxJbWKLy2dwtjUAKTa4Su1hBEmNeaHPIq8MiSjteZDej9c641uAerkY9dCRyeQi
zBaS+wmQCB5ssEGF0UFazteVkJHNF4f7CXHMEzDkKOiJ05h5jJafsks/dqggW6sCApg9NrctFqCp
392HmN2NUOYS4DWjRlZqDSNnC876ycXDOfmHr1ob/f/ZoOOulH+xJpCsJgIVzOGuEQnZeOzfW1wJ
5ekSBiI8BXsOzULEC1Q88JaXNDEzNz5rNe77HVOfvcn0K7lwatO7TT8WCB+P7c1N8cnmBE7w+zb6
nIfFRgpK10Kks8p0z/CsYJT7bPP0xEq58laF19y1fCUBKsDVosis/S9LyrqyNDdGDVtu5/3HPhM8
jvHoSakevFgpVNMWyBoJ+wX+WefALnOWdwLBJsKg61FY66AcYyrmm4RnxpXLqlqcroE9RpyY2sjy
13MpgtPpPwQlLruriE7HoMtoaJa0umVayiGa6vbEhpm4X6TDtY1X/oSml+Sy7ByZ5+BXkeARCf4t
zdpyXHmNn1vBuXBLwu+rYLTjtyOKg4J19yyfUgQpuQQhX+GYGkGT7sA5aEaW5rZpWXqgHMnfGgIS
J9cFK5/VRIUH81SA5uYF56P57d3H6MSTtj2gUgJdbn5DC+bFqaGWjEY93pfHSgZ9zgQWVTws2UQu
jeBqO0grKH45EhPhPemwLG6ul/wgOUeilWRfBCeHRrSHA6v8T1te/S3fxb5oGTbTealjJYPevpGE
LLnZ3KP119iBFpWfu+zPUWv15N7ArjBkZJKgYnXHr8MI+y8i6dPJMsaAVUCgGe05p3MPFZRjhHl/
sMgy/FnsAUsBXmOdpY8liko5UWx45SyZWnLsDP7AxELb+U1tCefVTGJuHIS9yet21qUirVKFA/4m
xruxILnKKOPAIUgJQzD2d3eCLk90ydkIPrzLzcR3zDzBPQc0fXl+oCpcmDszEeIMEriv6k6uxcLj
dLm3tAltNqWQ8JqWUpPxASmST8XuDmeWelYWdXViUbUNSZfbQXt1aPOf4iuJbKwt3SIQE5FW/vvD
dAHBCTC1XiMMjbtDgTmw16tMmF2ZYwihfonPf3esFUS/QI3Yu7I3jCzYMa+Sewe5HfbBtdzQZQG0
A079Fpc6+ACiwIm/Ze2I+ammDx625464z7mE2oDs2GvhqzgERFMy7/YsEablTVzl1ecxwelcYpF4
agEpTxlCWNoeRVS/Rljbax4iOy41kjhkSMwauybk3aLjpKCkrhzXz3yQRihBOro52v4ImH0CwCOp
XUNWLsf0t4f8rOFHIoDyOztty3gELM6z4PIBBu2K6dUFiyHNNjHALnlo1MUdyOlaXcXaIFENR/IU
p7x3nqPiT/g4t5Ko2FiqLJi94NQulsBbXQ3Na2+AWgUeEgvOa0cFYq/hCGv2C6vraesle3KAzt3L
e3ZWYoAReM7Tju3M0riv/cDeVQ4brQEgWtEPMBhl+z+oNLNzs50xohAdu3QB1UvvL3N+9za1OwTi
2/x8j36FhZu20M+6FT8bTo08vCUf+jwfkIZ7N9sKI4WJb9f9Xbk0KzVv6ux9crf0S9ftXcC/fQYK
JIphlKRPPXWaE7+9peOUgkd/bhuiZsvItjJLQy0GPWbgsJPbdxGf9A08y5t4R83yQWrogLBmGFiM
dc5gNmhDwDJbyQOeFurN++GgvWwn4xb89qZzfqIqa2dTUNAeCMNb/r2/VL7g2WOBw//PN+I/mLzf
ZrP/G2vOrCZkQBwLc8GAbCGC79hfLD7FE8AILt1U0bKH+NdPthGajD1lM+2iQQGJvsLKTEKrF5qH
tQX8qBwa694zeRzWO6b5tRAAN+cbXPUUZ3kH5qTbqkX6N39nYThLU+0NfOOPfvctEFybFyzyj7F1
kMwZXqJKVwn3sctrDg2i/NUBsBtVxjegzvmQCXrWU3X3Zh03UrR6b1ApR/v50hjVMHJlvKgLvupF
0dt7INi6vHoY2fGCFRarfyHijphkeeEsRr0CrmCj61ckmL48pp1FjlqonQzFn5SWzN8C7SDGxJ7J
5B/FCg2rM33izLMOpMCE2txcQEVThsr0FPetZmDG76ERVROnK69Q3lXrb5Zwo2vE82kOX0+Q+hz5
L7aBpkKxwj6IZZhCuzXxEdvWYpZk6S2QhTbUgq2UJd35yswjI1+IIsvbMTDQaTZ+UaNAaGAp3aU+
Gzk2wigE1h0vSesX0aXEzallfOYmRO3qWOmELSEzsGsPJ5ah96WtHefbDmWEBni4Ey6JngplRG8a
VWSw2bCbln0aYhx0bugpMxd+YPGhz5G76mGzvP7ah8V2G20pMpnNnzjUKoUWceLEGiEHfKcivzel
ScwKHjczfdo8uwou42oYjIwbM82Y3oCO1s+Mw5ULB8vSA3+1JHpsArR/adoj4adYK46fX4oRG6k9
Bd1GE0mSlsf31SmXQ9QQZyJftpAgn1Gu4+GE1K6QfHaVKL9ZsMc8B02QcTq/2mAIgH79J3h7tONq
CWHPtObC4jpFaGVo2BYF6uTjfyQgYvaHkLT0FUrwU47XZn/HtsqlcZ3a7MkoGSVlGdFprLIzZHw3
wmudPmSb3o7cHT5oYkrUd96xEWPXuCwVMs0xl1UHVbFkPZ6p/XrLhbfZlUDochA+Nv0SSkUS5b1v
jtQCy0xTTgHEZlAibaBmi30ENfheBFsQv/npCBgt9MUybtowP1BGKkzevt+SM70kalIbQRNfVTe1
UUPCKMnv0G5ksZU8XEvi4okQRubEcEPP64b3iqBkNZFGqMOdc5N8XEicd8EsFtFgnr0Bowy0uwLv
kHwnk2FNdeZs3LQN2dOGzzMCuLiRliO5Zqsn7aWNaBpLLiDE9RftaaF04juE3LnOremz4d69Ok6a
aAl+dDlCqzJLjRtpyQlDICRyIDu0QSCMd5+pz8wEDsoSUUo2us111dBLwXFnX96/dXvLStEKTbvV
YhyhAyvojGj0W6tSvrC7/Q/14OfkxoZfBAkakrApaPjQ8OP4QJJ0GhXeHvCQU2tgwDNF06LJ8jUl
H24Ret9YR3NySikKvgoGemKWTdzPOZDsp9Zg6vjVveYWbuKD2Cc2LWVFJ+5iddb5Y+Wko5W63pvE
vBufZpHd4f44HgMDpj/nQZIPB59GAtk54cqx4H5mV0OBOgjQlrMDLGA5tT5wqoOPKKcTBp/6Osxv
Dc7nU61Ulq6dlAe26sJkcENHg/r3hSvLo1Xz1p7vHrRHuE5i6sIQuQhU4fAZ7Qm5+B63PV+Zpnmy
Ydh8iBpYXLQoURYXS8kSQNuKcfLIwQmYYe6wyY+HZ3+qI2dcm469Yz9gX53aJ0Be3uFk/nGX2MK0
3OoVl0t5BmqBFDNHhVrA5kpst5gpyH5M+omJCDN7xCmSmkLkEEHdMzXmDThxUsJvfBr6tKt20ZJK
PoGt3DixqqmZiWbHGvsm0iGgFFSgj+0dCy2hg4R/L9vCLI3OfPnZizWW/0mMsKihOGtDpKZwe/NN
BVryyS4U4w+TsZ0qST+DbWDWjV0LXEs5ST07WESmTwoC+Q4Bw2rJCqxAi3ovsF1S1YWL1cOHqU6Z
fnpn58ZdM+BZ54zAB06pWg0wXsP83rmKkBcO2L/U2Vv0bKorFnCNwrbOIi0GWuf3h6Zteh1Qrz4j
sOnLtBPPdy0ZSgTY2tZOXk5GvylcFw9ko3gjtvqOBIsLA9MepiAof5wWMmPQBXLNZxi7mIwR31Uw
zJd8Ss2A6wgfpvsfIldSdbxGsiCl2lcVYnTLvEiMW7nc0NDmk14ytvWpygipUhVWNPOzsWjx1MiH
nUj9v+eXqens1pBlc9kLnj5ikCvlfP32DUNkx4c4dkCjKm/xBygDhFgLa36Eyf9+u7CasFhqpNyS
GTwLmuY9hetdrL+tgQa0SpuCqAqgQbBxchL5D+kqVeLihywG4duAHByxaAGVjeT4k5acQBWytgaA
YIMjB8oDaCrXnu7xraQIZPxkrUTsFE6JL81+laBXNqWlBYPFcZAWBUsFd6Eyi8WwwHKne4/CrPCk
1vlvIUmq/VBLDdPd4T/FyiQ36BbozchovuASr/xYqp8UtSAFQG4SLVAtq7I5tmvqxlHsscl8x+nI
FBKPKVnBmoAW2zcps+8QOFehurjbeZVW65a3Zshf4iVwhxz8aggmbuEf/eQc+ibBENBhHvi2Ve7F
w2DXfVSAO9AbwILGTTKd9dXvkJ4D3t6D/KsWSJP+zd4TpILrx1Ms4sg8sOviRJyfHM4fV0NhXSSb
un/nGthQYfbgN8nEaz4MA0HP/LI2ru7iNrz12ftVcoG6mEIBKT/GbA0clBGhZtcnSePlZrN+oFBH
+ZiPsQf4I8wmCACpnLKhRgaD7ewWsuzeO0WJZ3m9CUVJIs9bUtRif41bwj7a+2QaeQnLxBzXy+OW
nnRUCWn4PRp/t03PRPIUYci8m9yCHmwF4Q+IDuz/luSr3uHs7wkCvcAafSfg+c6FY1MxlRDN2EDf
7H7bTpiMMhGXifm3jgx8NSzrzdG9isjKW3FBo7JedX+v0R0J2OO7n1f299AT+xk38AaEOR0XHEvM
TYMEsSscS8ledYXZ4z90A58q+GTsLwUPthldLSnB33EKi2usjTexK0M1uEjlYr4rEeS4zgIIfMV+
iESTx+pFDorMIKzYT+o6h++J2NRqtAaU9NYzyehhiTmnlCcA8HFCRpUXNnewEb+5YFUJ00WkDAcS
NA8t1BfOHzQmGRiifF19wRaIgzciCCst3vQxZq1Gg+JP1WJDrMzHGQC985PcoXGR6oDf9wG18+27
c8FRvX78KGdSlYERQdM6XhRmppieNAXxsp7MrNLPPKQr+HM0T/NpGzRQF5+VcFEcEtY6IpBXIt2S
GqVAvm5hKSBnth++pfAMSww56TXhSAXZqddqGYV8PWfIpqDP4ft2KkxEPSOtBn8wlBuLh+C/bLzO
6aglqaOj1b5hNFP2fUAFVUwqyyVlXy2v6obUFN+AzqZUwrC8X27zaK3lhXDJYMRkMjMJBA/0hwd6
hL1342rDdNX8Gh7pQ1Csfi0muF7mnDUv2WMd+zYwpydESPhd5RSW23T3wDNHreobIgLiCnMtcWh9
qhu8+cs4hWt9gXhvlN7AOUAmDSgizsb8CGTwBB7/M95heWUWN/e2xDXkGaqguau1YB/lxlaqd1Lg
X9UiExyNLhRUGm7IK0UgWNL++vkeZmwtDt3MNVrI1J1JbHIBUK8KzUDdEZ6H6JBkc+4rLv8Sw10q
FjJvWTZ7MJfx/KJL9FMLv9wKFT/Eei0awBPeyrVb3C0OZyvoo4r+wW8Qav6dU0RMszP4u9fJDm4Y
GSxLbBAdelnSghKgabSFBqCORwjDYZq1gkQdO93w7NJf1cLqIrCN0rBb+1vbZPF2wNLxFXaAEXif
+4p8DPA4ivyAotRb9/6QiWyhwwgmf0CgpQplGhIvn4NVGvGJ5b+2A0jrFBGwe/JQv8RfnzcFcTTt
2joA+/5J01OxuxBSlJS7+2B3uY5V6esUcxEpJDNMkHdlnLNjWHTcm9FZjhZQic8txFypT3esvmMt
p4eiMolzWIQbLbujSUENpWEdYBXT+pDYml/cDmnoXwpw1Yn+lwL09oCrAn78Fm5syHcGikGXKwCr
q9WCao82QybqthyXuwfvdM3YHYvCtzTRMh8bZn6nF3+o6NR+BIjeawUnjsqht30Dc9SsMHTGooNV
rmcSaBxeR/4VRefKEmaGDjVgyvrCidKXS5qXTfuPuP6erDsjp8BWD261mYBoLiweyeyAOzpKUxBJ
xgv8ihcsDDsmljYpZc6gs9ZIwhQde7CRjax5eaaiPrLOyad+/TP3oQK64CjhDkTwVpdhztWgLN/A
hH180JUbz9V0UGRH3vvbK4r6m929fNktrqsdJCKeWzrkZXEPQiwXUx7+7OLco8cMT64JCJNz8aTf
PXxpjO2B5wxqIl+N2BxIiakTC6Fa3CjL1/fe2LISRbf/90M7e93xTUv7hpbebBVK7E02XXJbGlgt
UqyxhIGmn3CGsrTMyPGpjFNVDKHi5Q7SAfmRntCge2Sek62S/p974D7xTsVP6080Y9r+0kSuXm9x
qt+ncCUT/fdl91SqhO0gRyCuFmenef2MVqbj9yhz98pxqe+jPhbRvn7qCG5HuDclYj2BOW3J2jRR
NQeV13CN6BadJ08SjEYEKRhg/f/lx//pqiy2xHqoOTO3n3Qf/SZKi/NWRlnntVkGrHby58+WuksU
jpCd0KOQnGykrvxDkBrLsgVLIYvNMubOurkTULElJX3Y8kaLRRAJ8W/+3JnTUmagXRtnjbwa3iD9
Gt/MRc1ZrLWTwxVbsEitoC4JpseGl3WcCdb6ec5+IOh9v+HKFL7T/vU584SNO+aw1t9O5F5fRELl
idwM/oX9Rn65KUZM5d1Mybz4vfKYyQHaFz+Xg2Xz6/QSAaeXR1CXwxEPquc+KhRujL1ScI4lE+Vc
3FWdEiSdRz+xdG61KBJ4OwDXt2I3ivAnqnaom/HmXpdrqjRcsws9IWjhqDwblmXzShJxycoZ83HM
Q6t3Ym5HW+z7QrWTA9ZeRB8d8q+BdBL7+zupvruM5oFsEgJBys3TIq1Wv+YasR7p9hZhRy9GSDQU
yv/P1BAbZi60EeJHEh2LK5GzVEDMlJEb/XyGzStzkXDgI9GNuZEyNwnOtNY+rvLTFTH59BzL9izJ
TiRNHznlzrTXHBxUhKo6De0klsaqu1ZfJHe4sm1BMdAaLVJ0H/uF2p765L9Ms9C9s9bCZ41YfuXp
uuLULCmCGgcOC8m29aVx+2gbtxFeCcooXcAIKb4bSGy78YBIbw/yZkYEqlkxCqhtc4BADCmz4tjL
YfxCFEhSvlVLjDaI15v8eE1soar5vaWzBwwjF9LE2A11wpLMGB7y+M2GrjQeTwJbW8k/76g3yHc3
YUjPyroJmKI129g7LQhVcy7gUSor7IXi0q4HaF68YWA7CIcMh203YeZyX40qABI5K2tcpaQrhK5A
uW/ACc33Fw8HW9HC0Tx4G/U7JMid5niEHuhNTgUx51P+yF/RlDtZao6Cf+gUQJue2MzQcb+chCTj
3J4W1rcWkqY1xY793VuXmfKkfn1p2r/110YO/alVMRby6JLJ0DTfOCBd8N5RxeIiZWpGslM+vvZD
+w6tNow2gpzRYZzTCnnUejwjZs/YSUzVddaX4xPIRkEkXQMeHWr/5tlkacIps7vTqcyV1+hfYM/3
wdocgC9Ur8j09oLn0PvmRX/ajt98d+LfTU0Ew2DyKCEeVKEMYN555aZkCS9L9aW+FL+4U8jH893E
YjdFB4JFFZSSWHSGua09p2+sRc4UM9L8Kwe9GBrI6xSga8nBMC3+1Gk17c0VpcRWWarEpXmNcIxw
dP2q3p3vTfHCg6DlrhKUMJcctciE+Cl+c3pfD1nBUu6C4XcmOzRTK66FJBlKmemc0HagRn1K0iTT
KpctCJAwsiSPFmBaYyducZkH1I/2Zh3B3iDf/lmGqNCr2SnaN3P1zldVf3VbsJeZd9YnhQQHJHSY
RdlsgSeQDA3V9KqyCISEnxN04pIn7aNhc9I47D9ToHMWhhFxVohHtjEARoT70wEQzuUCMlpEVbr+
MU6LeWe32hAkNmKyxZjb5Zs/OMPtMsUgSvubVOxtXRzW2bk9q/jZGQ2/VTKdgP+fWU4Nt2Xq3BlI
NxRwnQwp4aKxLU8Wun2bQk3mDSTqocjt35CQ5BQ0js1gpYiMiShxhQH07vB1EHeqA1nTqfC+Vc+q
2e50dWo3GDupZGiQGQSMeDUkkSrvYf6tBFsqpeIAO7AtsoW5CZrNjraxrbOgZmplz7dqAW8Qs9ea
Ju2ewTZGEJGiNP4GYXNTDrFkrLeIJNlCqiFcHQGWzQFQFFTybIr/TLcVRPG+na4sab1ASeg3qeWn
Y6oDPiBRN8TNt0p+H9qc+m9sH3qUPVQStc0lvpVqiaGs55HZrFErLGM+PIfe0kWQJoHI893IeBKE
FdSHnTbCLa4hF/rbVOdR/iyeJ7NrlmqjmQHB+QnyFN92xc4zbkO7L4I6oMstbAjDOoITxvD3E+bs
fdrd89bNaqpRMJ4+Y/eN2vwXPD6mv6sgBHkj39odjglSzdu9ed6tprYI422uYeCzFnUJ4Tse9q0z
e7p0ZSQt42xcDF2dZfDVOjWkrLWISPcVzTAfYGQmXYMJgmTNq/GarXtOlmuNpKKvtSq9Yv8NWi7f
vFdRn5I0wcVOuLSAgfR7cvcc87THYpAA9TbzNbTd2w770ozMB0ZqxIGRkXXamkmOIgGaT61zYiae
S/eymayExVt8QHtABIhi/E8A/zzSQiTvLrjrZ+Z9lND2LkjvULpwLpGbw8niEEI+Hk082ipp8CIL
dmAo8MbC/nKJ9QGXAlVkJa63R54LRq07ZEhbVAFmA0XmJyRAsY6xpGKLtr2DfuUweaelDjxdsn+g
RHg0akOVSmHIzdvTYVNdaO8oRS/djcRXl9D2bXrxITXhntRqba5m4UoBv7JbvM61khdhXcFMOP/Z
GCldlx+TSGKY7ROGTM8qIkQvYdY9ymQPZakfdEKNU7OLutL1PlhjBE7fk7UBPqJLVYrdMSfOUBXu
Dzt437xihYCCK+UReP+XP413KkvNmqcWWXWYPhYR8B4r9H9xEmSj5PZfcZ6zAF1awOEAorWqcMPn
2uKW4c0CnYWZ4+xe5+pWco0T83sLQUbcBs/q/c7TwdUDSXQW2h0GgmqAuxatC801jMHTl58K6MAU
Lp4OLuBeGFKePJst5PFHMSOp48wdAl8DQ8xue5jxs9z7x2qk3hPdfquuJcweK3UPlFrMfB1gJ44f
WJcozviUNNJOR0ftW5Sfo5aKgRmfz5lPsNgJ9uhlQVcvr5HRlKzoDnFmgLnqhqHI0Ju/EJV+I9zx
1P8vuLfF/egKCQDdXeM6wFKhyDQMFQU1Y5Drv8LNCirjU4kMqFXl7d+Y4KSxRgivL8Be6bOQM52e
ySXbdC38WEsgPBnChAX5E+d36c5dEyUkGIbVKN/TUfJPAX2B6QkGDQ8ZKpISOYqFM5qFi6uEed2Z
zdLPPCBtyEx58mi9kbWWtbVTPgiUCF8yl44K38GJ61OYbqNjGh9aAPZJUYkBSqwGyd3PjT6nAN3U
5gDkp7jjavzT9bVGKlHlCWxjQP6+joPGNVwSZA1TRB3mOE4V8uClDO64dQxDzQlp5HGqXu50gZ/7
LCoRLGCk2DaE8HlljufvfyZvjzyphCFNvj67XToU675Wc2GLkZyY7rTOy3qhEYznAh0g2XYXn+D7
kBQizxn/E7WrUZsmdsY11HSYsfElGmxjPcLGUI1cZVCOTzRr4r4RN3BxgjIKds4ZNFTClUcil0y8
/Wz6N/fwovUGjfdU3qGROafIZ4wHCkn8zmPi0C3T9WedgnP1q/Bphp/H2CM/K3V9hyi+DqyQ9NMt
MnmqWt7FRbDZUSQUVzE/44qL65vgoUi/5yZ3ccaqD59FNK1cE+uPhztc8wfW6wIQl6HCnflIWe0i
EAz+w8yP+RgS1Ya/SD6ldyL7nyi1wHZ7g2n9/spxaXNa33gvVHeQ9MSvTFgSN0z4pWYQkB+jdoMJ
b13emyorcvPEu6eBgcGbsz+1qYx/v3/PWX0mfkMFYMXcEMC46hbxZpglFHDH76H0WS1e54D9zXY3
whq2heJH1+14H52Zk20HAZ5uheGUYNEUg1xnB3DbBYXC3pJKRFxFy+2Wx1vuk/bXJvut2zGAfxWs
w/YBew8T0YQMCViCx8EpAzEMmBpZXCxZHhnwmmNMgLIGf1b9ZNlZ5IK7UmZndojhRTlj7xGIF4ig
QR+L2oUUBY4rZfOspFUOOhLz42ck8UfnAYklez7AuVwXRSV/pjY/V7MNsnY4lKVEZgu30atjkupP
4nTS1bwvlDiMgHX0DMpEu/1PCBYuDlG5/GTd9lb3q+IxSTRtFQ0d6DjQ24XEh1do5ehXvFxe1zpn
K6nPfFUpsjUBNErSggmt/JPrvaPF56IqcUDpCgwBEGxcqRQhYWdChnpUuTqfJqM1B2vOLa4XGlIL
UqiEIAIZoAndm/rJYB+bz//rZ1riFX3R8TQsCJbB9dESuDH3pGNfDTGcSry7eTIbcQwrZYnJI/y9
CDSxQ8RnUiaJIDGyfNbMjhgGojlKV3RLKQLqQkzGFJBlRDSPLg6IMh5O7fbI8xjdpMtVhWFSj/ZB
kij3I0pIemH/j+RtdpYYj3TnYbBlK7jEfVf15UGvRxUncmHEKK+yaLkp1AhV8JnlUn8CjDNs287S
OJliqqBDAbEvGoARzRP6o9Wx+SU31widfP6d29FsARU9NeS/TMPn9OswYHhKQ0Yw+ow+cgzqiB7X
kMlX3aC/fisERqRGPMEajGirVD4lAJpy22ebnreQSzKAKh3+oGt540lnxmLrj0yYXJN+bUP4reWc
toF9mxLgH4ZHTB08vg0Wgorx2K0w5cMG/pzkLuaabPEopR+346SAzIIWMJfRIkSKtcgGkmA7/Oga
Ja+8t5l1bWVcGBnICydMFGJfdDoyh99Ihtf/bQFopdHIpGt/f2QPOlhb1tG3AcHNGK+Ks3Adl6Xy
xchF1kFJgyhYN+cLaMNFe4e+Xma91t3Nk0WjNwps94Z7IXoUwpNjyU+Abcihe8BLTvI+kDW54dTF
kEkHn/m9Cznpu4ipbRY/u6nE2xNUUcwbZgHg6C6gT88YwletALmPdbECp1rMU6ue7/yX3yKYt0Yq
13BxLQqR6p0ing4zLwT6fo1eftegXyjhnDEH4d1BZ0z5fpXnY/cStICqnGXMcAOcgIaPFqtYz8SG
RcPZZyBx8vUtV0TRbyTQOxENj+vEsyUk0qPscCR8TcT/qsRkc3qEz8MSojKtkUAy2n1NbIRDwj77
jzY0Mkm5y6CzVL9ZQ2+um9i9k9otpC1TeSKa7YDWy21d/wW9YHdlP1VShb5f736pCVB7LLlqmFc1
AEJw0Mypeenz2qMKeB7sR7VBG1oLIxKQ0GEiGRXZZEihEa0nTWnt3X7urAhuEZgFkJKGSpUPdmaG
1ybr54XyZRQ4XK380lrO78cPHvCWUnhJFOPje1nga8Xk8j1Q4kpr8fEsZxr1Iz2VhyDJjte6pjob
UEfkTWNmq3k4TJ8zIiQmLRIh6dqgJK2YEa0CDGn2avDIb8UzHye4yBsOQnqbyjZHMV/1f2H2U3Fq
bf+nJMp1fX4klbx5bLYagNzey+R1zhsuRqj7Pp26wXcIMyNEqrW13eybunoczzWpC48P4efJLIRJ
IGK6XchEeJ/jjAEdrI3ckXWhPDgYmdoq9yoI0xMUVkg/GaRLT/ZggmU8TTRNgiCsdo2fBKEhFQlM
Q7T8YCpvQfuDTx+3Js88mP008HH4bOTxPILZPyb6fnmzbx8VYkRJZuD2wxr3g8EezarqVYHMvd/6
BZmNq5Sy5udMKVQ/lGMXBYk/v2yzWcxb2LoGZn2ilx5m6Qs0GaTdBqnBRQv3+yNCk6caZNJBThak
abLkow9BzvpKWp04aGaQnbXV2OyjBKEqTR714uaiMpgy+1GYhwvHa7odhfsARtinoOToIo3bKiC5
21RPVZqVu+XWr/qF8osBk/Tf5RePYpvqiyvlJp8fGhoPdfweBu1D+6euzEC6Ynod1FhTpztlp+du
+YpGriT3xc3jnQaz5MDW4YzdiAsw4vZC4wjb5wry45b+1Yzpd7ZCv0OjG+JXpoFAU3PtFLFuA/k5
KdjlW8jrku3cYIGazn2RdOjXHPqG60fnQeliBv0cnmMrRzXZkbmjrjfsVW8v0BbhBvj/suwrw/Qo
6vg25x/2Mb+lQk+i6YaP8wzhwGAk/bn9f+4BEQj/j37RBTwcrNVC7E8V2onyIDx0rTdjCzdvxxbS
Te9F3f/l+K4BzOojuO/Mu9+1WOJvz+09qb1SZzct3IMGW/gmiGV+X/Xdy3YNwtffc1hPNdj38AN2
mcCk3Rc5KbinVBG0cZnrDu+mOEbIUwOga2hJBVDZK4icHxctuSFbXzGY4raJhRhVsXUTOu6WrQY4
yJ9r729fo2g/wqS2t38wewcf+n7O3dxr1avVVoWW0du5i+xDwwZkgr1FBE7iiJ/zLP1DkuGT7ghG
9QzCtTlXcHgIc67aIRYIifToKcHwYUtTfWwA6ffjtyoqZ/Gk6ZctTGl1uhCguJULYnC6vrxq/lMu
LmPe2/fxu4aqDbekkh+8Ykvc4fuaWpRLQK2uF8OzmlfO85aSrfhrRIHQC1eXaUNA1M7a3I39hxJl
y4BrBigAIGFg5EiT7133PBvOxnwNDtd0v4vy/yFKzmIjgi4A9TyS7zSc6VpK1Eut2egGsZTTBnok
wqpvkEI8MgCv1aGvJyqDRg5wx4fa7KMo9n6ws9sblecFQM5rgFzLbi1tagGVAI48cmuKvnbk/YFI
Y3PAZmVqPyNV0DRcIV1JfyZuYq7EshNRhqSuSisehOketXkQsghZLIM/e9oksw1l5TgJ1IuHvevf
k9JurM4XY/jz+7MYV7LTZLhcYSGPn9Cb4Fj/mi8YpiVbv2Sy5lSnHH8UTHNbt+i4wuVOd6snMmR9
i8V8+uA1pAcV8JdFDsCk7FnD0p+2p+1YKt63KlBhQ6wzNA1/L7LMxVRYQ8KJRUx9RodAPR7luUcZ
GLuCkwOmtdDcIV8X6I/S7KoaCkEnwj0JE5hd+9Uyn+ocow0gZGz6nJWWMLS3PUAVemaLT1fWdeAO
s3aWSpngPEfGH0OwqjXoQuJBh/fjDKb4qu4zhny6UF2qGbIRx2X3Ri5jV3h2o9byYGrCq6QVQJEQ
EsGC2U1+oMEgwPE2I6T+RIY1bYFTA4VMBJ76CyH1YZQggFvzLgJMnUAsYwpKorDiS5t/+Wby+CK/
R09yFMy3vGLSluM7C4gvGye7WBSnrn332UG5At93OlbM+0ZFBg9WrXE16rBhlBw4yVKAX7v7Rwcr
mBHBBwuNmTIAJ7/ypSN8obx1TLZauwS8Z7SX5kgFKgy7ALdrSakUE39/kcoevshtz5CxvI0kLr+H
cW2bqrFstavBvgyvstAjWxRHugG7gILV8+DFUQ1RmHnC4nWBwAR39pazzvAVNA6JTfw8niSJcd3J
on3Hom0VeIBPdNcc5gwvH9F13J7qhQWTQEZS/OND87HPpEvg4GcvMKliPW73wNa5EGsy2+2BfZ5i
nVffKzIyMp8JfefU5X4ok3JWrH443Kr4ub1f07o7a8dqxehpQd5GJ14KN372Kv7lrVaTCkYtK7p0
9f4YBgFwQCLvL7kfwREU4HoD5lDQL8GLHzeScFM7iQCiuLNBv8nEKyxuJdxrJgUthS7/aDhAdnLl
7myrwDLB9kyAC1qUh0778q0RyAZL6CfmnjEtiF4Q7E5v+jWICXauRpxOvY/VidQ7MWnTZoDmhz86
gyMX6+jt7H1m4g1pTWQ5FWaA4/kP1Ug0u5dB5ItAGizhNwGCovwkfug36srcTXqYGeghZOmb5cnL
t4Cmu13juIODdcpu98pET3+gJaiDELDYJsISmLnLCknh/afAQDSMaU/fw5/fK8TlYOplIybZQ7Mv
mi/6SJab8WIdCBNFsTfEWutLCbK7ebC54+nVY+490jz8V3BzsEotCU4JN0IYW8Lx8PMMAadekCcV
TW3PTsysyGVGTAk+NM6q3ke4teeuT9TS8aJS1HcIr3ljApyPsYeTzYY99Rp7dYkzSYCUfFQK8AJA
h0SvFjPsHHkGrMk4kXeYXsA4DYSGJcf+NgRuvzP9bMxR4OD9A32QYK9qcD9h4fkI31MEd7lkh9wa
CvYPd0IxXCnJ30AlGCYlwoBL/X3XOB/mdovz9TkmT9wxewTdYoVmXGq+BqeUf0/1Zqrhec6zakHd
ceTIz2GfxO30ttqWaTbDV+HtY1k+P1actcu+sLnR4ADliDachO7lTlCNBSl7xNLE0KqueZvTwtuv
6ecwBtaAmfJWgDbH95Ma/Q5sg/yp/JAMeEj8Rr9kIvUIlPt3nhNjnSybrYtE1UjE5w7B51ev18fY
Eu+Hzfc+cF8voMfDKLDTsqzjkDwnOiIPE0fSIwUOTO9ae5ik+TDGW9BR4wdSKq2g1QUu0IIxvhBu
aqBz5JhOKua5EL4E7On/+Xk3N09hFQz06X0o0mDA3HhKrBZ5xZM85Q0MGryFgDWhM2WvpOsJ949y
2W0F8wjn4ulUYduruCeEDL/FkCoQekN5/Cy9EJVrMSaF/DxX4/VGAI4c17liqNsbfX1UQ/BYxAi7
30Yacn2vNP6CfCA/QXIRnPe/95t1CS+7kaJ8Lr5FE+vnFyXRmQqEuKD6QGsiIfCmh1/KcihhOogN
OeGgwutQODedGwgUvNfKT/mz9QAjxk/R/3Us7xAKEvSJ3VVHfWhaNzPJ/0fzUqelASYrNlXEOJvK
OjMm5P0/X3XQ879IzfRorfkcIOV791pXNi2ecrLobhuC8z1iJ78+xJUa9ttLazXzeXpvuEcH65Id
4hyPfXJpf6egHrBacOHJUFcyrTxUcr/5C3pGwMdjnyOQjWMZu6IIpQ5gS02ieCBDRqkHex2ES3HJ
lr+jVjkw6+1/eITsk1m3XmT8hGc+kK5jKmRxP2kOAqzUZ9oTJTioalQR4dfUJiJgCN/cwP4czpnw
5Akyxtx4fwcJFO6YqnKwx7upOR7pJwclmyDu8gflJmBI6XeQOJE5z2D55WuOg/p/B37IsnRrGkHz
6Q/3Rt0Po+JKwZBAiTxN2blC7bY1SKzANNIiX82bmCm33+aXxbrJBerxm1Fmf8txQYS7ECp3ppW9
ZvyoJQOxvoX744/0YNiVboNnc3SbY8qC2hdd0asZwecMVeVYcDpY9pxH7JZrjixq5+I6PfQsdZq9
rFzk11zrrM0DHUCItIThfRQ/qWL2kGUi0A2yMQ4M9TtBMe2WPpmUquJYlLgMwfY9NBLYcJY5vOAt
+Tl01GjJG5uOKSL20LF/Ht0anCH8/TRCnmGgFagziPdRHk25XudI6yEKDOVbOADg0Ynsz+gtfbLz
V3mslb4YxN8ja+/8Yl7gG9LSRzdEEVJD6oVet4yxkomwx3ikyuOH1+m1I7cgt8ZxwwWjSpS0d4uX
8YUpGcDSAKdzuddjNd8dxf9AifvzCNdevrQBA9uPsGDu8BMCCO/hIc2wmt/MhexwcVRlMkbdFXOI
P8XldnvKhhHIzGqXv9UH3BM2jRRUCkuD0fWefk2bQZPQx2WM8MyhVOq+/87NbVG/sUSLDqhS1Djj
HlnDRXjG5MJQoilpXmQS6OXUdJc8+QTgwH7Q8Za7V+aJdbMUCkUj27G81Di3Y4UN+2FeUEaIz6mZ
OxIx05z/b6htpokwIEU4nVDRlU00K4zUoMbVqUB4EsCnScCJIRRRQZf8j55zkqN/gi9jB0FvGEGo
rterY/pY0HsvRFfvMVEOD9txrx1uDlHriLurgNTSrBxMacRQpRl2QRhlmhE53x+zMxzeCY5W0RFk
+cV6EgK0bSlSrfwQEum/FWWn5VqL1oHStNM17ORSHWRq7vDXkPSY3q0KzlbKA2EhVjETKUc+HetY
nzrSKkpjCLOJWBEvRGWYDEbsGT30DZsg8KSWihh3KpK3p7KcOMC1sWHdi/X4qigFHbgtkUI7k6kC
XKYtngoosmUobzYIIkPPcTlqsp0dkmS2Zq7BvnBu6Sek0BN7Hj4/LjrggZehO7slYKWdLdqHSPzO
MXobOiyNlfnydSasQytXrWJq+fh5WNs9FCmM4GGynkBzrBXuJT0LK1wyNYzIQKwH/Z8RX0NJb+Mv
/OAhNxWpcm2tc+G5PVyHHt1mv2wbFX1g8vX9dtil7y6FzqAYs2t47BPkdomHxfbkG/lBSDWpmyw+
Q52xiqsMyGkq6XS6itAOh1a3+PEsWxo9H8kycHJzinCynw37yV4XF5KbRtfhljYvHRjnPnCbcD5I
a0ajzG9hqDmC7cYqqJpwclDN3z1CCKE3hfKvlvBXzdoZTXla2lSJXkaYK0gC+ZTpClomTg6nt/S8
nIjiTaiHJtygs11xPWunY+Zb0oXYWfxx1925II0QRbECPzwPwXO2MpkNOxYQGvWd+jSNmz9iivmX
rTYslvI+UDvuMseWGlhBXNcdolKZEQq3kT823vNAJqNx8UEpgVysVZIDTmRL5JkVq+n9FSi7f+cB
AJ1N/DWYkcwfs2dAZIxtTYvevHeXUpnAfZAWd148ohqKS2Zj7/smO/3edrO+J0xTHOHWkBTGTUrT
KC5yHoVtQNdB8kGgllnxJUZgqzr7DhEMJgPH8AawyuS1QlFphsRm9pCtHulR9bwATpGOdz7X60mw
LNoXftgV7chNXhqYRCmr1rO6MHKjh9zsNAzQCIC2ycVNUt6P5R93NCROXRDS5MkRhVMPHDp4YF2z
VmUZS8zNOctK6qS2JcW6DF3pzwQaBpVTSP9ms846uHkoSTH+jUxrLF6zq1wiGA1tt9rduKsow0XC
zLG7lSOurVcLAxj7g7UAhCR1h4v6hKHQoSzvw1lErnwF2jPRm9D876PYLQj9QKQVHNY4bh55+4wX
TkC+STx0hByvzL8bA4j6IJlcGL8Z/TqMsD7vacVlD2E4ivtBSD8Gj22ms6mFyiKzzsjTGo9gTZvI
PMGmmPrLAKusdAZy1Pp4wWJ4YfZg1YyoawoViLaVbms7bGM7P4QWwdPd2Y4ewTNYHrzrzKXiHppS
hbfkeHUdFl4gcU7SoIa7RzvXLU6x1hc4hnzupvWfVGRaHzUwTOf7GTIdqLpfuM7ZKWnyvBpG4SlG
fO5x9A5G3US+vGXJdAsyYCe1n+LHtySLcAU3+yVJmL8FaY0QO5+axDPjdM0gMC5ymJPQWBTZ1Zfz
sirTBfXcPbmt4vTgrw66f3jZJXPM62/Z9jCet7bBdsjR36pqj/rfsJP5LHvCOjlllHQ73boWnYiO
zOEX/JQctbZRZ74ue2wEfmbzI0r00GUIHQfOxBijzghBq9eLL/6A/vQExRbHceoisLHBEQbgONsr
UC8TO4lWpy5Lw27Fk8gTAnJPNuLuXeS4hpu7ytMEEdj+ay9g2/8XWBJohPe5Bf/GE5bybIsKniaV
5Qr8W3JjG0ZDIPmOghc32sZIztfNm3xruMQroJ3BNlQNYamBnNwDbMihODUy2rOe9adZzUE5Vfh6
BpVpv8X2hZuhlPiPsJpok8muy0S52oeK3cKXAoQLg0F1UHPtJRYpU4v5YGsz8fLwL6ZfjH7UFMH9
krr6QYtTCKI0nQqFciX3EMADBjvy1gyNLTDPCBMqk4vhU8gQRVUnoATFlVeHgD4CfKY2i3c0KLh4
WUBXo1Mh7BnP8q72cRsbLJAbTKt2SA1AL3atHaPsOLHmD9UuS+MMLWY3KozUCGizCrsaOq+kIr21
3np94jfrppNGNOl0dCMfcWVfHOq95iMnvITswFt1qtyT2jdkmS7aiPdp1/3cPUOTIQq2/9os2yxe
K1Bb+oO8JP+Pc2CB1SN4a0AK/ZOcCgDcBJdssFxMx5SyohyuM0hE8yjRt6cKz0dNsjeSkjM45EM2
73a9R8+e9R4DUSP1hccqn5jzIu9cwBpYyhLyTyyMaKX6BikH3h5oUBvMCCyw59O3fDIVvO630wSG
2TaRyIRxfDCs0cZCN20LQ6CiiY1gIcFpcS03QYl8NkNe08vdwKfPF4y8/FBkHYpL6NnPeBsygv99
ezdRmUNQHQr4hojxiSuckaNh+uUd+RCa5+vtddC2tko2FoJGMByoguxZ1gnWn1YuzcmuDvdBxgvF
AnKDYOJBpB+syw8E2zIY/wTPsD60G2Jo+qsIxSJi2jZ4dvbrt5fo9sTm5RddBlBixmQY5VWtz2Iu
l2I4/kLZlTjZUGav8U90dFR9BohuM/nwGL0VY30iPB2j0HzsNss9+N4v2po1OXMBKeyZmkqB+682
h1mWjLTU5Tqlc6qnCVngrs2E9ar3PKvir8me2QX7wkIR1fE8LWgr26kVhtNfIIcYDyj/DSwN+U6A
yLeTFdobNvV6Om+vEnVas8BY77XkBspJ4Wqk53669IckbYBLL98BWbNXQu01ds6sS3KJWny7vYy2
PAvA1HmEHe13WsOmAOTNjcjXiX90+Kex9erc9gWlcJI/aUvjoi0QC8NNDQxR7L4cYQ/NHm84CD6m
do8CvwlG7I/PwE7AiQmazYmW7hD0RvkrB4WTYnzqUS/TRd9uNU9VN9QYGIY5jr8gAmWS/lF/kVOu
ock81C/no7oIDRQiv3PAALCmk8E+6uZpZLN/tJ3RVV33fK3PQDlNIo4iV4InSbSf3PHwc5cXOu0x
cnFD7L+Ek/0+tAtkLO40QccuVgqR7j3U8fxyQV5RyzwGxKhbQsbBd1ubh4kifIsDQqRN9ni317aK
XDQ9kFYRCxLXpws7uWtkfhIaIwM4yodiI2uuSpzNmkeUM53e0QC8hVNm0XB2B95Bdm/JItE9pBKT
ztbe7jE/KKQEEjJRrd85UM2T73mv7ZwccMMHW5SGxC4BgufBpO7oC9l/PN1a2LTX2v7se1FDD8fT
x++39nCHttFJuaxbJ2XNI/dXZGkADF0vKFIlURZOKTpM8h+k1/QQMWMycZluj6I/ON38bVJzq0YL
r4ym+cJWeBMa4/TdtfhFtxbKm5NAYPDBk4EtoOQiv8c55v7pu1GeXbF8jG8nN2q1lSbUMonEkivq
ZPcxMYl3YEFONyyuG9afxd6kjaxOv1kLJTt9mpK7g/1jHWNnDreakim4z6aTUje48J8qWG0k2wIP
EfkFBRjHFdEELq6yGXIvLZ8SQzrB+Vtf4pGCjyKEOCsi8Md9gWcFOP9/gFMGqMeg9TGMshLoIyuS
J8B8fnflmefgsFLhikR+Gk4iNl0AbLCHCNiTrR1gyxmofUAo+QkDKIbo2DKtyIDoLfeKek3sTucf
EkCzUG9gbQ5XSZTTraBvmInlDCorWThrDwoFm+v8jifHB0m/Nvg0TxKcibh7Jb4wWIiY6V4Ub6XH
QjBRAi+PxAWu57tVCnzNKxuj0C4isM/KPaJka6HvG0/4ZPaf4xyyzAegt5xruR8F3R7zbyeuMugA
gJY0qRNLnoVFLvFqFRRAZpTQ3ogRUJ0TF5fpNZzAZ6X0LWOrMFkVxK3JKWmmpJZtptW6oai5D3OR
/bVKCskrh5xXsqdV9PdviBpcE69HoBqrivMSTxisdjXX5U3F118s9DM32p+xZqzRBc3TGFNR2BGX
Jk388tu7kZI3INmV2oDBl5tLYdW/uM8B7Gys1pPvv06ZaMa+yYxBKBvHYvtAtMKw+J4B136xKj9v
8kBv8+h4KxZObY/ekh2WKeBBh/ZCSLCIspn8r146QxoTR7EYBxtgxdH2GuIMogk36u9vlQCCyHj3
NLqbxPipo7JpVJS2GRcequhAZwM4GRv4AiRGLt46mtHsLj8lbS05RM5GK5bCt4E/7WiGwu3+9xPV
r3jq+YAIhUyd/E4VbyxIZ1kChLo7M/LPb1BBY2G/Sh0P31ath6XDLvaZ363TzU6SRjgYPRHey5ua
oqtPbDDTVsG2FN7c0DyOQK8mtaaO8++YfxvrsEr0Rd5jRl4mQ94K9h3S8M4sMyGrlnKhmwN3EID4
D9SXXP0TdxhttM+yQo6PqXKwFjP/t9BjSSoMvZ7vOI+vzKaSCaTskavEAzRKqt5m+AR57P1u4x3j
DfhbR+0DdUMqgmSzNWqlm48Wn5W++AdSNTzUbZfOLhNJG5O4jFgVPO52aW/gARVko7aIbcBy7313
VbzNIRbjpglHUYMRKFUK9rtwTLS3KO1sh57AfZiIcoz3Ulzzb8Fpt1z5XWcrK5Y7wzdXVIeloEZG
C2KhR9w5ClRZVifw2I40XkUfc6222cnt3v/JQEkNYX5S5lARh2UrwX466dSp6VytQoXXY6PRh1j5
X+Sgb3I7ZjgeIAKzzczLWvy3QfTeMT5j9vphM2duRjtk59s3qp+qhP6siqWfufbwqTckjGWgTTKU
RIeFXZ1mxhSgMjVBKYQv8RzGvuQ1IbIKfTWa/CrVaciC1rmTYhpnwT7h5N/2S9xQW/90WGTSmFji
AjzGDxxmAQSpTbDgIK5g9pJRQnEhOP3btFxPoqG54xOomWbFy95G9De1FMec0wQqaltcb7jisg++
DTCV6A8lavp7waABzKXoA9K84mqv7fDUNrobdj5iYizxq+qytpBOmuDNngA1ryL3N/CL2jR6q3Po
MI/4yIK8cAUTLcN1wEJaKk0QPBRpPhI5rn489B96qN1X89aPzQzBQ5WJ+1f0fmPCJQzD36RrGKVD
9Fl3X/hDGd6DJ8mRH1KjVksNiXIlJCIRMqmntsEMbseItsP0gX42uOe3KDICbLwbuU7/NkxifU/r
SiCet9ZMLX9mZh+O25UMkHNUpqlg7GsyRBZaoArSQ6TXoPjnT6JjBWuaFTWRgLpM51latrTkVaV0
ySHv4FgOSiYfYCpRhqXzJxhTpi1De13FNu1c6by2S6kUc5HIbSIKHa4Rhh8wPhbqrw01GHZPPFQE
r0pu3RdpGhWSkK19DtxeVHnhrJzbV7w3oPEaH6mJWqi3PXjvCbWOB2aXDjPJrnbqrr0Y/HgGqf6p
U8qFhS2PBoDZbrKR5ICFeZ0j6sNBi1/Xxp3ocNDHj95RMjtAUFQH65V1I+JPZcz3OLFD9X67RH0R
l6bX8tPbN+QbcJNvtSHKsJ2F2zlwqhr1VknCAsFpveXv1soTn/sDV+Kd8RD/ksn3dISvl7mxaWaP
ALR3n7mMJ7PlD2tFPcW+nq1gR3PQCCCL+AP68ACeKuCOK4aAXcUt66PTsI+zl7TPWoaP4yXZEj5b
cBfkX4L9sKT7Lijr7qFPFOFADFMyuUlMd6wtxd2ZVodBgp5u/R1whbAqgsoNJCNgSLzo2wuqkH5Y
a3u9wUKmnCx/CRsiDwI8nEXhKNOxZ0unmzwPDzNLwG+xcIQnTIbIs2sIudrw/pIDSxdNiMluy/iQ
BzKJJ2mAiPHs0DzrU9AxMjfs8kB5g5MzsgutjDakG8dQS4Vp0Gq1G9O7Y72LZ33tEZZVEGbTGRZ+
FV0ByNGYU1K3oKV3p1MZGi9fmNA62vZ4TUB4VKU9ITDoUL4Tg+dPMXQq+9sjD5Ah+WSFubg/6UWi
7gTln9vNbua369wPgPSTAEOZdEoNchcXqgX/5uwsOQ+CRCUeGYA3HkO8XYHp5g/dPWeWjaWv5G3C
SI+h0lY4cLh8RLsdRWeRWGHp8n33bqbqpE8vivXwjkSwILIqp8CT79xFuVXuA0jL3SSWQnBuv1tc
ZGCnDei1tE377Njm6LtgYdx7vTUq9uDGkF+3rysNe+TCFslHx3VqB+gLLGML2bacS8pfOpLaFn3S
C83pXVo1/IuZSOKqM4hlnxB+/FTNO0sCI3UXKYRYvVn3+d1CZjGrzuHnIBf1fLxSodVhIrtP7246
5rEtZKtrua/47AKhZV+6Ky2n2ccPTjdDzRH0OGpE2rhdUHr71ncOw90m0VZQQd4FvzXa+CUiCh4B
mwAP9d/X/ZcG1x2xymHEkVgY8nm6IFYKLzR/XbFg2zLNG53boq9uIKkKMDoR/dNiRqRlmAidM7CB
sVx3Tiocva06/gA4qrTIOJ5I+SLOCFKD49uT018Vz5MfIC26Qg50Am773fGKKa8O1RJO/BlMCBLS
5wkyRyUxBYl94vs8Txs+QHmz+PZSZvOJACea6/B8+decnEqcYQBTUxMIKfYETvJ4/WvgQHrPTluE
WUE0SYkrUzVM+r6dVR5gQeHkMzEyZO2mNOTpbNl+d5cI2bwp8SDN4hzVCWe0auiUat/z4reRYNIH
R/YDA/YleUgVTwAfTR/DwPuvMP7RXe1dk2J69pDOSZtLH/MqZfNT2T5ebhyYadKAlufL1vO1r2Ka
TcJ9uqqTUQ1FlQ0eLjV6PGjboZueiqDSUwESwvzzH/l+Apnd1KU2/4OdO5swv5QGzGZU6XyzcfOG
AXKIwwlXxXiJXTyNLi5figEcz5BBrlmSON9/HAJjgPAroXg4ssqGlAdGiyC1kOGjnNH2gSvon9jG
Lvs9yunQygWBLJCUljRVbq6mETKedJnlzC1VDzNbqLYNECUYCVBo7IJp2TPG/PtqlJQ4YAwa/Cf3
qLunhRcO+P0Dg6oFWPStYu86nGK0AH+cRMfiQVTq/VyhavD3pxZfjl5ozdfnPa3as3Y9kSwowtsf
W7s5YmRxfDc6FG/ADTTBMgkXJDP+mURMn/SXqueP3ouQGg+XUyJMN/akDlvg36HP1ZgCYIphkubq
qTgCYSqrfvjwGxJRDltwPDN0J0wyKn93xl1V+8jo8rj4Usn8Pr5qH5jmDCl4m2yrs4pdEx0MtEhm
jrYIAHQQ6sjkAo/oQ8IYw8WItLNU408e/KkmAThO34L4TT0mRaLs2oygtcoIwfVYIA+ijKlb8B+B
n3MHp2TMD3zEUksTZcfZAuux4RJQw3hpA7iNF2ltJEKPa11VLjpx8OvG4Kz4H0x2LyDBKW5mqM1P
OkuzGThowijGv4AD5GCZoXVITUR+a0vDBEOWkFvXxqEZ1cFLb8Ce8K/CBFSOEIehBxe116QU4n1G
Q88gLiHbjvvN6grQuu7lzu+oPOITDsN1dM7tHM+tqciehyjLeUHU4VajljQWK9iQHEP+4PmYeozt
fNOXYIl6jmTKFkwhUPKEKXKkIId/Jdczv1f8ewv3NohNc2SysGvj78XCp+Bu2/CdTLPCf2frfCEx
PHoLKMn1asGvAtvlbO33VRufZAjFO+vPcw0qg1xCM+lzi2yGUY7UH8xLi3bAXeIP36+HbFCoG8sG
U22T0ZlDCgQNFvdAsBaQqgE37dZxGa7e9pgk0I31+fF9mHQ0Tp+4SetBtXZxJcgkgloaspxZFxNK
oNmpFvx+GmJhDkVaTTm6du0LyQLME3QZ6xQQYOuz1rWtMyIE6PnYlSF31ATM4Ro+p2jskLCw3OsN
chZKj3YJaSivuTEM20kTqMge6Dqw6iuWoNJ9ncMvR0ajIRWVX3f5wgwIVrwn/UgqgBClHJAmVPGp
CVLVH0YpFSrfUVYN40dfqR0f1dmvTBzXT1DMmr5p6/fxqctyRlfoXfRgFDDIyrjEk09x/Mz7GpiP
RvKKPG0agKAo/3jnLYswGBj6K56pEKwiArKonYNloz2aZCat81C/IUxrgghYuUaixQ+xLDXJbxfI
Sd7VaBYjdE1svnhKEFihh0llrzoamKhOM+Dqf0Sts3hP6QddcsBuxKrexmwwEbEAoAMldv8jZX9s
XrjAiW+4MPHvbXVzHNBw1LzoExQDw5mc9SLKE+ZXP6D+DuyLH9umXCw96mFnK3Xo4hwa1XYcwnOf
RuEruHxS77cigaUcHWNNrTXRV5jFOu6sqHnmA1q04HbZ+eAxuvrI0zYW1iDTJJTtJJF+nnCSKKMK
snH3KbRq72DtljN09tZUvevMvj+Qzpf3OPzlOSXP2r/CLD5R06JToxBiEFm5xUlL0srUqPq5eJHM
TT488RijoVBNGAi3neZEuG57pADNAV2X60QDhC820Df7IqYyYKg63Wlr50dgQcIMUHOQiS1xe26d
DlSBcufUiUA2pSEmkg5oxpBPbXDPd1S6xA3PkaYg/oG5ozZJGvwIeCr5ztDN2RyKHbIjwWTtwN7r
GquaMUdoKKlidG6D5ZnI4N8IeXNjsveznvTFQt8w9hLUiv2w5mq1vRmtUKodfUqN4RdsKlo6CoHO
cETtBbAYWBoLEkiR3eUqKvBlT9ogGYCrKuFz8vaX02ThJ4daR9Yol60j1y+gA9cLCUGUV2QR1ch0
4BVPM1EhSVNdmRYDiw6qkeUsmR0eNhbhE1M54u6wJeAD/72b79KFdKPJBnlZvhjIuaXwF6g+rT65
O/8bh/0GFCdX/6UFgwb+Usyb8Y47Gm+6jOPxylE2eLKmhxL3jizBga4kDnCVqPGrG2dnTGvqZxkM
myuBA3HbG+zclxT7kApY/Gli65LEYmdHB+ik0aaEqjyhrqqoJpdFNl47GlHFOmnR53/5gzCbDNOz
VAiUxGekfKae0QwVB9VFuDMxkZEYN6gnANUsupk0dT+Zl7qBtvYBeHFt2QZuVuJE4xLYvw9UxITI
scZ4pSD7juZvdHbyM6udBxRf+JauZtkMOipcu/gLjHXAHYGlvDsOKL9dUE9urTn53HYB0g73r5GR
EdYSJuzuji1Ixb+YgoV6+jZv2Lrs1TufD1dgFxVO/UEEh7PTxVXACs+/4FMPl5E/z222aNfyzMFQ
cAva6oDHR1OyPyHyJvpxJ6z7WK9JrKiQrZ/yO/SpTdxJCv3g3UM6qH72XLHapoJpdKLG1P6trqcE
p9Aak27GyLDaOujHZWsqRMURdEdBFYh2GH/KKasbnJ7KkNnKSQi50CE8ZwYyHt1SRH4fuH7Gfeq7
wfTUBP7uMBeymenhv8f0lS8MpMtjVKTR1zlwLRYRrCpxa4tZn1TJsibPvAZcP+rMCrV98TdGm1ZS
pr5LF165qY1XslsYs4+BCYf2c4QAu3UJRxMB4cUQOWyF+kllSiOBLUjwjNYu39DmtTQtNAi/f6QI
FXaXhgGVYw+uyQ6qGKaaagzL4WBTRgFe9MWdPlJXLbD8C/vk0jC0uzrmrNqu+whZoHuvMLSixk1q
JVHd+pbxVr+xIDat21e/0N3+4otm40tJi9hubfaLx8Eggrs70PlyM4XpChM3JlTjQWRvmP97BoiQ
ktxfxGGT7Gojhg4+VuPeBzI/YktDKoKJP2PRNcjug6dBEGnQERSf1N0WWrUU+Hz1bz6loCTgY6IT
SjJhO0LjIaGCAGOH2iCoZI/IwRTFnDBOSdKO8xvN2FN+RkcQ/okwuAYjc0O06fndtjBMwDvati7J
RS694YRu2kzDjsCO5xgsxFEiVOBLn/KnxcUw0qNoplJJ5uHsKCsiRxfuIlWbyH2ByBtoLV7OYfZ1
42Lx77SAlfZ2Oy1c8Yd2/Yz/zh5XyAUrf+PGTcT5OJqlofSxaeYCOxePtrkzjDRMNv0UL8AMGbMz
QALXjdk0+FtR0UWH6lonfUzXlg1xJ9MqFV/EIh5iI0pq6mrgoRXO2a4GMgGtima1FzVkMkj+XQSz
y/YMA5MRyimxL79G9cPdak3ENd+B52xoR7xhXwTpecuBYDyujkyvB7uOEAIicD+d6wAl7zy4KpT5
+zmMYoV5odUWjhAZ0bKqd+R2qszcAiXxnekJFa++ByFUP859WDhelnBPbxgc9zJ5PGwODuXseUzx
tK3bQysTmjAmR/kHASD14ceKVzyBhSZAIT/si8HVyJkMnjn4xDlAC8mNoDxCjm9ZW+fCEDpzGF/G
AWlJrEZJSAUBeAqEso+MpvbTAOo/OZDfD/US8ue0ErfXp772pv+awNSAynBZzyVBvAwcgNs6LAHK
MZHkR07h4P3tczyY8pucXURK82CX7kKnKYqnhnM/UTlv0L2GEY4EFidvm+BymWFb4+9VM50EPR9+
8Gdb7zqPF6RfaluM+QaIrg0v6cQzQxA/KVSiM+pcth432jvTKd7vXTq8Lg1aYm2Jg2MscNlIrsfR
9NtI3Xfp1Q9XJKixlEJV0JnL/OEapdLSWYmNi/fvjbq2wYH070ERiy0gpljRJMXv87QYC7MEBCgZ
uqfPHect+PEWsIU8f55lzTL7Ai/bh0sl1P1BM0zYv54AmLCIdAy0m/C1A4v20wWa8VijEfiBciRh
5cDfBnYj+O8+3WEEarnS1VCc9T+aVteaQVaWDbA/VhgcI61HmDjVXTujHkaIiqqO3JcLr/Fd8bmt
X0wdKhJV5WnPK7r3YrCOU2ehUSm4fPoy42eXZVCPWr7tclt/kMPuW4zZSc7uWYqptiTzwybTTIj/
2bJtJqY5a/84sJ3DIY6m9GzKO4h+CsUx9/rj7phVu1Bt0wGJXL2epL5Gg2IcBaCtLM61tJaZnwMh
A648IcpXNLKp+Ywj2XRn+Ir9nC3rKqNUAZP3b3GHZOf1cHcyf4cfMRuMxOlMWr4ONMGY32NdDZXq
+PqYABPEV2ru/4mchMFDpere9ZxUF2x2dgn+YVXCoo3X3r/n3buHCDuaA1N+b9bIL0Gbj+P89/kD
A5OIh2SY8rvIlYKEENT5n+tSr2SmoOoQDCrWO8t+A57NTNCVMgJp3oUFXbMcGUd1QI8is7dQEwyQ
FKMjuF9nP9Rxnws9gy/dDxvFO7oCPAVzthV7aX5YyYbGkB3Hp9dZrObYrv+VRMoPN6+rqpNZcj7H
ZagoDHz4SzOgH6ZbhWHbsN5orssi5nMkuvq4Gg5mBqF3NE1TSz+P+c7OrdRvnDWtvXERCLVar0m4
sMhbuSHor9RBtRsP5I/TJ3VaTGdjpQievTGzs2kLCd/Q+7SGchAKH7yhMfoPH+l1Kq3umLSovQnd
RGvEy1B9OsEZAwsT01P3NapflFnmP3gRh0Zym7lzuiWyxaxL+zbXnMZJoWC5k+GM4cd1RgoiwTec
0wjQEfX3WN/MxTj/ni5B6k2YtAv0C5BqIQB7F3/3kEnD6jJCy26NHfZG1yXl+KQCWsKxuEJpYmgH
LVX4ce1zevd0iirYSuJErUF2IINRAH6accrW/jlQ5lGyhiCougT30vfoGuk39FfBt4xT7JX2nQnH
8hOfmXCvW43G2aH+7lTZTe8MOkBOOmqq4covRoi7SlZz9KiIGoQuDtr77rbpJNS2SB/5Fn9k0amZ
seC2nyZZVXC1DxvNBPDZ+0jaJF2cBvVLLgHqKd8lru+NLI8blp/J/755cesqph8CSA4wKbVf8/vZ
4C0vhsF1C8ukQBnZNqKkbyxQwkqg0nfYarH66lMp0Bs2EjHrnGE3Q3lCEJrD+GLgq4nJ2YHsgXrF
av9hSSkofbLwL4aA0FiRfI5kqa/i1u2cFXs0KSTZlSzcMjRItUnRVhjAArjgVEeEThC+ARzoxSAU
df1HY26FbypiOtiuGsrTF8Vh9EZjGv2a5Jx7FHJXdCjZX0hWQVncW0O82Mo4VqBN00QgjMTh/A4E
sDf8Fzqwakh9W4ybm2kXbYGNdZUqNfUnZgCU6LcExgf/hJDWh9iNKZ/tnHraiwXyFONfBYnH/D0O
eM7p3SJYP9xAEldeXcDvsy1SbtmbPNOiJ0LuwN/B0FK//Wsr/ZQEaSrOsq+U0JRfsVtOHGlhi9Lx
lf5Zr43VgOjoo1W82DM1oO2lCBwnnxo1DHeTzhrQ8vqfI8jCoj/jL55TXR2oS3Ys8OjDGwWLHTnn
7DU1aA73smkBvYkqpseM/8HcGa0X61W6p5y//b4djJp0AzgLh7OLpvBJvC9Cy/lCiGTeCGkpHmOK
Z6HJF7cggV8rgNK2fVIIcMKfXR6KJrkcStIvgaUeD1dqYFDe1iGDmP/M0abTDmn+APeWroEVFxmR
COBBwqpaMOimju6q2hjIGbFtpM/aNI+sTWWIIbiAqHS79+T+a3UERtqLGDiI9Ezu9fBDZqrLf9EZ
xMp28A2qMKQ7jaTkNXC0WMN5LQD+35txwHIYqDuV5Q/sOTKIBXnNDWCdLyFCzLB0d8m9MfGAr+ta
yLTwLWSoC6HNWiQqyD3SRuIqn99YmPnb5Fd0omX17mLwL2HvfpcA0vtSUaL5CLiPCkXDX/vLQ60Q
umlvaf36p/wTBw1NtklSIDQjH/Qd6Ax17BKYKRnaXX+k4oW7uTavrx41qeGJN3VnoefNzzg8bqJ0
JBznFJ4N9nFy4jssxMklvi2UXFbOXox/bxoeS79WsyMVvd7y9yom+MHoCLnwBgwzCzEpklYQ2bB7
g+MeGplH92hy3OlEj4oDsAkNAUaaZSeuUMyS01LURPt2T3EMvdziDsPFZWC7HI1o7cPH5N9OCEzD
s8M6PmyodteXp7gUW3ySDUlo15GgoNyQbYiBoFm5nevHUY6ERLA1Gn0weBt2unUzOwgXJ9yYswi8
tID5Gx8oDsXuRdUTxMnN7RW/nFiP9KQYamNltfyaD2ju+zZNbJXjMCDromCmVXRw3kbJiTUWlW4O
eTPjyLBnmNCnu/cyUJL1ln+iAntzxb5HmMVP2bttoXTEm9EIg3oH6D/ruCCjtQrXgVk52ofspWhf
WH0uok/tFyv9xHP0PkoJA5lqGNhMaKHOz7eouyW2ePAP8LZiLfQpcWptLD8AGoE6HpK4ke8W3784
awdmjJHvV8xa8cIFWizJclT74gOXN75osVLgIOmAiI6hZGpVtO6NL9wNQgp2hlsjniDunucSFWYp
dYE7YieeflbKLuj6rBLyZC5O8K9C/TCMdQ4GswzbXo8bU7t5h9jjybDnkDwqak2PN31hDQepJBkE
j2S0YNc0GfJFmBf4QvMpBCcKEp8RXZhroMTSvNNqcciBLQaCE+yC8oSPkBxB1g5HxCAFpUt9nAiC
PZPSYDc59yMpso1qcJTqm6JeKC7Cyu0y3kNlTy+uTP1QqQx98/Rt7bBpLgdVQxfqei01ZdZS7boT
i5dTxQbVF1JJGdZEAfW87TFfMdqnlye4jWAbLR2u9Eht8UHY1v9nmZMo/LnDdsTvDcA3+TlVw8pm
kO2mhqd8IwEucK4UrXFADml2yVZkmQwcpT09SyJmwIerobQON5IUxRoxPat/wMOM99EDQTguiijN
nFj5GCQBn42ZpagC+ifdqPWiYXAVagVN7fvbHNx4bEySYK/DGyDXaziqiOdYF5vPHVYLHU/lPw/q
k48AcfalPbSvWqlLHGml4GzsLzUGNXqkee135IRoG7VhLEy0hGrWK84n7yk4sAPbKKMJoDR5P5YO
9FcWA0ejT0vc48dUwpJuraeDfshLdbaBrIr3RjjRbvHwkFATl0+2HqVu7wDqrOEB+ZW1c4sZTnrm
gidIHggdoHr8M9uoaUFYiV1ZEM5JsY5TJY6HtA4LvfwRdTAtY1rCqozfcbU1JDHMg9ZlMfpo+MW3
wlm0qiN6aPBGoDJ5Fi0gFxKSLMn6Ji8aX1zByELdqUe+rqGBsTs5ld9QuBdsCAcqgSwIms/ljr/t
gIHXHoCv8xOwd6NJLxcDpc8Fawd0z9043OA8YpzAbjgQotxpjILZs1G2ZlDxTyKRuSO47xjB8UrS
DGHuKZ50F+Nzn6pdge/jC6ErlW5A1YXS5xIESXojMQPIr2NRR8OJXvEJRmFJImeu9E3/3KcyhMxG
ZwvR45abaPqNFbUlZ9WBnTGpSMiJQFgsp1lVqg2rmW26Id9NG/XAxRgPH1uQR3dfnfBPP0OrO+1j
i+UoT7xwPKZpwp6KVRXeffcKrwKApRwrubhpSfyOipcnW3LWYWSH/NT2vxwF52R8hBH4dICo31HA
ubjvMbOXoTMm+vzAF+6i8qPyvNHYPIc/zBuwdzS7+YCBNd0fxaJlnlEL523D8TvNp240IXXgPKe1
mriP1hzjIh9qfQe5OJj12Wh0HaA9ohHbOs9/jgK2dPZPy/hvokDa6SD5ukSyiMQnyUCPv+rbkIuy
COjtXzIcd0AFpy7dLSGWPZK0McFKWhObciU2y/FAc537/4WR5ln7enVDT7f3mF+fbl8qCd3oir9c
S3oCUK5WRirxFbvZ6GJoMsPeoni2B9q2ILQrbCVEVjD/UnPR3xfnIMeI5/CeFe97UqYwAMlGc/Ca
BxdKXEEwWSR6xfWrQqDMzUsr0iLpuSYEAWF9H2iEFE10PF3hx20O6eUyNdCadHcttPQbhRR7lPr5
bWFb8yLlMRJRuyet5UO5MjaOyC64TuNJmS4O1sZYQlLg2db08ItkVPVwM+w8pUo+KAuyZzyvb0VL
xgWeG/OywbchM2fc2bWPOenHZkPKHG3xIlbE/N3jGskjHWZLhj4DAef7KICBfHfvd0ASyueLjSaw
ZzSom4wPn9TjWE6JmUR8R0Lky/5yvfLpYptt++OU8tmJDVccCZV6NwjKy0zJP1EAQVmt7nNgupx2
tEVvojPjiXu51X0ojmm02l6GrofsmDDac1DItyvBS9se0U9qsBVGbocngdHWCsEH4RPefJLs4BSa
ei1LQbjjgiW0TbvxD5F078Pde9QKT2AdsNc+sgEhuqilY4xRXO4qSpag690asNGrtGzQkR/1+vnM
yf4SSBvoGdyXIarkg8V3fl/iB6gP8nyq9fxqSDP7eUSHvuOqYueS20TU7rpHNNNoRxpHI8BleI4X
LPpq0jFj3/K8WP+ufjp4mO3IA7RE3x1tW9yYeHGv/+dfYn1UAIw1TnQL9R85CMGVT/o66ilTda/z
RrT8ORBYvWLCnF4Rluoh1Vfv9SoSeS/DzZY9h33jigImG11BvGdnsQ0Ch0FOQn31AFCcJTv2dwDU
qdD91OkN7HF6AilNMZkY/K940Rxo2ap+GgI1PYFqV09GAkwz0IBFji/kMv+szkRE8McGrDv7rlEk
lUF668k1pwmrcDzlKMYZIQhYtOf+g3exf5G0S9ssOrNbxjBe5L+fRFRmpltbwJ9ucaHzHd6jW+7a
cBs0iGp1/+9OCe9X8Mm4TbaFj+qsGwfCqJAgN2jzwViL+fg5RaNVRjJU15X0OD+Zb2DCYj6BYJgz
m5KpW+X6AP6Da9JQUYamfQgtjZYQOkBymq48gK/k8pVmVRADu6Lmopz/HF9IPhZPXTG1F76i38Bj
PWNAjk4TOXzwdyLeT1+2K+Dfj2n0X4pVdDA06h0qNwwzyA0+3kcKoli9Bc/u68pT1NIyM60Pe1o0
7+HoEaBVTmMLeFmtxOBUcbsF8+455dm3BKky0dl9UOBiVrbvqHb5+wmUbJq8b5UNdQ79YBVNC0Cu
yda6GqyeXgixdWIvNbFaj6EwqgIQyBZmyIQoDO4o9atP6xldUDgqT15TsCJZPGx4K14UorYqyiYB
6HFhtKwNxYSEudbu8MMmHNwwBc79n4NVVZz0mTN6j3oUVrM2uqpk9062XOlN1UO+OqNzN4XQu1RN
Z0x0gYF0+TWJhVNAiEqlU/2bai4DTAa48gR6EecYY34GXM8T/wM6yOVO+KNMX4EV6mIiw/nbWBV1
FcMD5cfPm8FGOwn6NprJ+TVv6G/BcMcVjKdTFTQKksIsDo1yCtegBsrAJ2KKIyHpPs+rZLYKM5r5
uo1dhXF6vJHD95g0hZIMwXey8l24lLHLc+XSJjdH9paot8/X38/QeTjd0uKwvaZ9WPjDijwYRhb1
0qa9nKtYiugCodLotnnO82Z56Pvyy0pS7Rw3h5t5O1FcfcEy4l9bU1KXIIEl0+31T3w69c1xlxhU
s6EqMZuAzBVcgQwONVoLOaWCduCj7eBhJHXN4gJXlVRhFhIXKBae4WtKVyCABXxTch+OlEkPYsAQ
l8N4n+ft5efnb1K2W8zV4P1iT0YyJqimYaNuR+vrLuDL7Vxj/+MmWUVjWvp0/70FJAPm/so1bZbG
r/zn+xVHU1yCI1C61aFVTY/LwgY4Kt9hqvzeJ/Agt9Z+SRyxI8w3G3b9XOt561Jl9yWrB3tq3jOD
YX2S0ims9eO+aaDaMzLX/vn49EVTjw0UE7Z33p1gLVApLXItachPyzfarVDWCPenNay07u8FWUEP
MbD9mnLoMZdAtaKDANoiMEaL1oSd2ScUZA9/cp6FDLJ2jdOQ9pOYLzIW3MlxqI300It+IZK5Z44i
0/gXNfKnVWXOBmFnOXLfvubm3nFHdLxsEWF4OMc79jbFGXQ9GiZj/BnZ8E8NG9qXEAP/p979rxFM
2Q6yKZ/+ONL7G6r8DHzhUY80VuRTiSI/7AYLR5LzhV4T0MHXz32Rao8DwWeW3ajYt0zdn3F5Eout
yU+fE+gL5519nH7+u1vx8JKbYNl/v2CpbdMRwV0V4Ju91ki1YIJHWJXuREAGBN1t8HYr2DfLQm4X
266hPAXcsF/DX1+WZSRVmoQWp1mskIhyhAX/dLRZpg7cR6bZutVkf9H6bUnqMJpVzLOHPu38nvD2
ez4Y4QxSnzKHXDYFr5/GUAVSBX/3Va3BJGAphVk85ucOKGfxkk1oiGtLM6FQ20H36NL33QD0wfPM
bgsvSg0sHXE0Qrfwp4UtMhIdEyvqBxhsxXTJrDmOzbqLawGzU20v6Timyb2Uj04Cy5H1mz7oXBDP
pud5b55H6hljI1h0gITk2ZaNCLkrrJ0cWI3kx2lGLg692DW7DMNbFxgFdhd4FnzAY3elwZb9FF+5
Xhip2sTz+wYKXKWGVxRHfzBwX+kR+SmG/gTGa9x/mwDpJ/dgZtav0nTMXospu4zYRmdFA/RDQuSE
spammMlorSesgi/R0s6Zwt7c1XdmVr2DaKi8YvrKNMCYt134+VK8R2DbcECWBBG/DGhmDCisaAU6
EHp/dGBS2SLJbPUIPnU/Pbl2rG62U74aog8Q41Q3/l0GtXkRew8sSYh9/gJ7+dWALBns+APY/Ssz
NzE5uqwrd/9gwbwmyEvbJzBbCv7IUu+7OBAbZslg6QZyIW9TJQr7FWbJPf2jbLNP7KSJ1Y7EFuYG
XiEcuaLg2hI+D0JJmjFizqSSGOFzh8zZ2wCgcQGN0s+gVYi+t/BkbQHX+xr543iOtwyAPyzsZCQ3
fMDc5mFLXyPWHPvxIhFNkfIBKOyGbH4aZHI/h1qw9GUl5UMQD9bnA5N9gtEqHzrSPy2K8Xq7SiMk
f4F14MUjqTJ4D7gsgFVlADgwNXkTiJdd5wi+6niaYLl1XuiYkYCH4JPz46pmtbceUxv7UU30X2e0
GIA5J3+eo8aoLeiG7JCsfJoDceR201Np0m7u6T8hk7sTJ5wOHgxjBnwOyp7ZQobqLtCtHkrYPft0
FriapgSHE5DlvTg3oAk6T8uUZtgqnH+rPKdticenwyCtHwygkkPuR3je/qSTaFU0rchB/dDGpKTG
wEZDAIWSLvjCJEjKCRZkFwNVwkN87GJHmxJbjmbpAgQsvl0znveX+4RF4SgiUpkk9QnZvjjS7OVP
t/uVXYF3Z9Pc+LY/KMTaRqVyinSZUbRLtSciLQ15d6PcLKGHuUolQqa2cFSbmyjdOvylViUPaOhy
5QSwVKLu3FcXkVJ0ogYkS+CPtQ07UKhuc22GzKpbpjfQa/WZvzngZvWv5tbr/zKEtCtKSMEC25OJ
7VMfRrGQ1l/HopYoOEdsvQGv2hXKqp8wKK4U7MKdMjrQbq6FHZbv50FG/ZgSiNbSXp+z+7btmGDZ
V518/AYvGOU42cfJDVnlL729AjNYySbZ4S3Uoxmxf8DLsz03v8xGl4oNuHE+35T/4QfV1M9zXpAq
fy98jaHQMWGjTo9z2Gko/rph697imjqjGnp6vMRrvE6+DGNog83SEHGgRMuV+lV2M4jZpkkmG+z1
DCJr++rZmBOz4SDBn/GOJPNIFYxQhHG5MGQRmd8IskzwoTj2w+l3rSTxvxjM9kwwYm8FOtf4UTLw
NoSoB5iPXy04bzYqjdMaHoqkYKvzESPeg95Uw8QZiscDX+s4zv9BZ9WlngsSy4qwvHAegyz+uF6E
DczuO2srDfdLEO1ULsChwRVYTXIDwDwLlWyxo/16pFlPwVXQAU0vlDd96mXjQQ1XJCJ72XX4W671
HI8Kd1DuVM7Gtoz1XVixMJwhTGLRF3eNihW+sS9GU9GI9qr9zxmuJrxrzqrDLDyOfeJoFt/1V3rH
RACs3He0Mtz38xdyaIAgmzcRWnYjXe5+7pModpWgEY7Au7wQF9A+F33CU5W52NGoAWoLqkj8uWZl
Wp/bub9ZK/OHar2UULgvD1D/Q4HgCIkFQMLLE20A0v3m+YxwCuFzBpIsV+4X+rPtZbmuM80tZVcy
x+NUehc5IgHohwaHHRiFrtH5QPDstOCUL+VeCUkW3J9cxv+HuqjUrGiVg1SyCRXcHZ/n+kB/TtqE
CLBF0NCyNsEi4aLgD55jB+iR5deNU1aJiAeml98ikZnUv0k9auAtf1CvDp9nhri2Yw0CE/513BwY
Zq8zbZGMbfVhtfa+vStbOhmEGbQydry0YRVffvPqZkZOPiEf9AcpSoPeduwvpECXW+CABrPHPgnO
HOgCQurj+yWpQgEitECwVnxhFpLEKJ3ngMq7HKPo7t1kGf5WlFNfwTkJSoVcRQTPigkWu2tsPMEX
8i/ucsrLMvBT7+AwhWtu4wfkGeqFqcwScm0cB6wcX+hK09R5I0F87a9qrtDwNf9kcM0D1mUqhUUm
eCFMPKvSp66o2mR2fccyHOY+LYi3MdDg3hmL4Ma737QBL2BvjxL0HnwDjdCkdHiPzoIdVyB0FlCx
j7Lq2KTClEEwGrAEQ3/yjaOGZpa7dI0jA6WFAjGa9yRjRsTySjpB9qJEaD0Yf0baAuArYYh82TYs
hlkiZ1AdLo3ZuIz+k5aEDXr++NBDcgqJ+p7UR1uncskNFiNINkDU7aAOeQBJ1OFSDCha9vK7hm8D
hnQnZ+LYLi8M2hpJJlZD3kXE93nE5ZZA0p+7JczYIOHqhpiq22CYEBJoiQJZnPrLVdf57XtInp4a
rvPYgPrhhb0cumkUTdFCuXUyUMLyaSSYiarHvKUX6RWbEJ9gol0jnkqjPxD/6Fsa6goTK9J+yiue
SZowlEDBYH+HGzMWxA65BVeB+1BDrFYG5WnmLDsgmwc1SN1wBEQuCOVqFwkJZRkZOx49AhWHT/+i
76/dyv2roZuj8Yy4pAlb57lc74tqFIul3kclaOEfQRA9c0xSappMHn/lhm2vDiUSbBm1bgPhtf9w
4Edll97K5Z9Jl3zBNPUKjbe0J8C09JsBkWNLnOoCMmkuWTFbtVsTtfgeQ/aI5OUIrHOs92JjcH4b
KX0/+m2+1NrxUFMzaejcLcz281nt/OEIUsg5nSi+adW5GQTTgreKONWvnQnvlHmOeqx6kQrdyPhX
uY2IsxAbRffln/rqh/gPkl4q/dPqNk3THUcdznRH8hDMREJyxMz8o5CU6GW1d4u9upTOGzY97gsO
QM3gfVPAPG1CMiQoCaelVfouEAaoHKTtwJI+G2H5wn0oTo14eBeYPglRmVvEtDpoxgO5fffQ8n9j
wxpptEOotYoLc5XwSk0SggyspACAXYEPkhK6RhPiWo8O4ARq8/q9sMNMC07+aGz7VIjDZ90celdK
FFHjSBeR7trYvrx6kT0dFgctJaKKdcCceGIkQ/BIr6CgwRErIsgNZgC0/W8h+KV8ojrF/IbnxBd1
xw3UqYPV2GEy7JKbM2Xx2UKE+M33U5ThxD0xW1AKvzqtH7c0hTTPc0BNiO/8csbkefx6moNTG/UO
/LQs3otNe1IU2cHB4bQjZ1mEEWRfOMIP8CJOSsCb5bvI9XX8O/RCmmWkTl6UPwDLMZS4Gqi/Iw+r
yW5Lws+tfCqsS4LZyiMHluzlHlImLWxCawEdy63kgmHXJZbE1XTYWgyCxvWXC+QjJuZE7n+pncmn
U10yS3qqTX9zGueRaT55xDY2cdlTAVGuYjWjRUTgsxKIbUF+e+7r7DxvRVusBadvrhwI3OkhcHjP
OJ1/Etvtp5u7TEk1bD9i80zviGpp2ji6sL3cuoP9Fh3C6nJO/W8V+f8xja6Rf4Mby9pgnmFMeyDY
MbNdVEhYvb+OvIw3XuZpEng3V4X9ePJUA+Sf08z4VAEN6x28TrmuPooF/zOs6GYeIzKIhCSpc99+
CatG4Y90R9ZnCg5VMee+ckAZ97ShvrBNZv0SRuju9szoMZCRGKi9E5JtydZ6ow1/qIbTAEexATMc
O3jVOzzWI4WujS5b495OKITe7t9OS2PjE4tFIyf8vlK0IdMWxTum9YtDuYTNP1Y6w7EZjm4/t2YF
Y/tLz1B2YZ9j0qQAMpvgoowSMIPuErK2BQN+nVx00n6SApIm2oglpZm4svRuu+FiwcKI5uEG7yZ7
UCeCqB3dvXIfFVgdA6pIcQB2JK3TlgCT/h7hMUZ0ihaONrEeYXuwUvXNpo3tfp0k2+kQWkp5DWFK
O9SNgLtaNNaYwnOfz6Bw8b2TF9qFZy1ISJ0+0v80t4ZzqJpABF7f99OlnLPzJMnBGd7OBNtVzj+t
cWUxWm6UvXVdZ3ZQeaLcIWFEdDsPEEVwJV17nynRFdedxJpr5cQIhfu6w/aLxy2VB1mCSByp82MX
7tRxTjSf2zJXN11/NJSkDuGKo4QIixsIQszeaJNugc2K+i3jmtOtYLYU16QhD0Bpsod5Ke7mkCny
XcEy5UBvZgjDdi5kqueroW8GLQ/Z7i4DEgNsCCbkPdTxhnv4lDmx/OaKGIXmGQibuQr2LzuOLiln
hD4B+gzJyWYLzDXkQTuePUpk0JR1eC7rrnbnPDR0r24plXAcQlZYiopN+tVi0FQqQfliwZ+j4IlL
dSGUM7l1xkUVyLpivWuA29XiCupSfs8/ZZI0C+ZwPCydxiIppAmxgHYNd/ugg9LKx8yTN6RLktPi
38TmB/jCp/lwoAsD74WD8qRvelcj55P59TpC+YyU17MR2gyqwUFDhgcVE7OrUkkBlC2EbwuCqnXO
Ezhb4d88NAK5QLQaJMM4w85IPFabwlHrfOVhhYITcoAQy5edfNcDZX+jjzveGSnA+nbV566Q1RN5
vYic/O8g0W/vXpG+IRnmepbPo42Rx2qcuktpm8/TMXX6cSN4fUlVpL7iF4TGJ6mKloJDiMq8pani
bzfQpgX4KZxgKyzMaIHnFrkMthDp25VfI00gOy1BDj2yWZfsb9vGbe1sr2qP48OXf8Z62JS82RzW
b2hKiox0ggqX4g3Bnfi0s8512QkwiiSDJ7wHl9Io1yZYq+yjTj/pf2EfMpdFNP5gZPbOk2J+D9QC
haTEmPhzfK+u52VBtomtp24o13I+EHINqtUUc/12+MX7yTHjh2bwFvONPyyebDpdkxF4AvVxWAyb
775cQaTEdNaISIzKTyOJhcW31I32K7IGEsmRFCC97iozefiLX04rJbyiQ4MRflZo80ZIlYVtweA1
fqhDKneert9kF+JYsOhI07HxoWdp3N8wbSenP1beMEK1ML8Bui3vQcMvn5SvYC9Z4N3pYP9DgydI
M12dPasWaWh97znDFxXPvc/E+vlx9PDXqQRRtn91mqBRjzFLz5vlYe4sReY00sTkZ0udVtfmRmB1
ihLkQ3/YEqIeEt6CMotgjDGyL5lU8rqOHqeo1kLy4FeQuzIDayx//CJ7FLAeOBiiiAih12zgluR/
HLvPak1+eULTgWBBsX2V3WXI3PS7oQd9V8xNRo/5bfXDxQk/AgoGKKHd3n5O7Frx9J8O5VhJO3uV
8NOIMW/Gs5ZJfMJcgWhj8Jb0yvYYDS6mRpHWihxiJIa8Ccgg7jpbbIo+owx6DLl0xFOOrq4IgcVT
0Nf+bz5RKWI0I72xKaOzlIdzoc2Vfga9JN+ZJaFdkn6zqI4cPBrIo6s9A2udvldKjXXbmWEQa5HC
27frLD0kITNuK5I04jYMOxjY/0VZ11BkYlmkKwzy3SNyj+YxCicO630Ll6EvuQmygfmfl6DjUQWV
BNKCZf4n+GM+3Hr+D1sg62si/wVdDr5DBOKlHuLFrjbb1Km7OqL4wUE56FsiFkzzHWgzMy6SfTsk
jN1LQU+OGrp9vnPFrxfBR5lyBe51EU4CsV8h3jM5nLXbPaQOw79NCmLKVCNS6nWu6CXiSG0R5qu7
f5vh4lQquuSkCc11C3F1soWte0lhaDOnOtO46dDL3YTqA677P7W0O0L1YAw/q3xy/qoEyP1YW2ti
Or1PNRWcm4GtKdFAnaeGu7zzLnsdg2NKxZT545+EbUeKhwYCJMSOLct4z88mQnG1A+u76WjdiByp
eJ1MH8Kc9VEtvCkumbu3rk/RpV6z8OZpiA7m5z5SQYWEfzKmjPc4nD0q+wbencwmc00Z0Dl+MC/7
LOYkxJ5gKSC5bp8E3dIX48yD/pcLY6GUDsHNpP3HIWVQoHlQjxX+dkIgmV+0aiLVK5Rsaj6YqQ1P
30/7kjk8n49YTkrIXxUHaXZjzmeNvemVuNw8DLRt8S1l3Wj3b/DRJxtRyOI8whFxsZiju6Y0jYRB
yvVnZ4m2hn4viBZLfXd+i8JSp7HaG7/7EQLp9we4sROnJVpB9zIOeMXLqzRr4nSKO7ugEeiBdNpp
RQxDx/8Fvi/VDJ79KjqjtgDDpZ+ezQ+LBw/xhvhN/ylPlMZIlWheXXOHfoqRva3mGwPxOmFvbFam
ZinNLVD6PbE0LBoynCDBM2meqvVLFdKf2DoPRHkCZEzyU9+Ecos6nygVFlLzOIlMkvr1iGL/Egrz
XwLbiEuJE6NperBd7ZNhpoD6SaKcQ/sXZ8jzeV5p+Hz7A0wF6lXT0AkoTu2v4+r1Rlh7qFHhyt6Q
tXQrC/2Luwo1DsT7e2ZlNdX9t4Bf1ZDbe++FowwtRJAtv0BXHrrKVdpYYYR0gy1zZrUHzFcYyD28
RgORQMujTzEj9Q/AGAl5r/BBQUGZMcgwU17fNjb8+Fx+fpX6ocBUnpLEmx61bBqKrzdgWggHZmft
QlW6kVh15jglCqravvknCLfGMUvGk+cO4JNqBCXxGnxXujxXZUMb6vod7IcAZ/LaS/e9d637yS1w
Ue74v+JvmaajNQGe0ZRFiCeGia5LDJKKP7r+iOQLaUKZBI+1FTqTVIdVBQQMhAHddAVN4/ocyOt6
D3Q7YKcfyY7VCZmJeQYniqP37cUvjoZLEyrt2pXn1WV2ivuvhk60Dh0pIn+WbKiT28dlxgh7VZft
n2Rg5OfSmz5gdB4rpLhhXFO52jbCNk7dcRHjEdzlnQEJZ2th5Ys7TiiLQIURsR3O3GET91iG/rqj
YbVAZIbuCo3fH8ynUHzFNc3P6IqWokTEkeOFH8DkrPc99kuFy8Rfr52YNd5VkM/5nqRkPEFbLFJh
o7+yZSlOiiLE3kUEKkYir/hMH6WwOdxV4T4NhJvVQqeaDRrjantMffVRZ3B4A/5xMShMtynjyZe6
bGYkKQfc4HQzKz2OqPT8gYFxfEuT5iIl5GOeGN5n6IrHuAZTGZUsXAgKtewCm3aAFcgvsCwHL99N
Wu03+oeHQXcy2ie9xbqCo0VsVN26OvrHg+4ave/pMr5e3BlrCjXcOqylFL2gN70zqQGSeadnxovG
5TNcVzCGxrDbHuiOqdub79kjGLp357/CAxJ84qJpz5nWScGshJroWyC8RtllQ80Bwqsic/p1ec5o
bC5DOeyJGQtpM2+ASUQLtMOTbydPM6BjNYSCEWwQOgAjcylg1iWErzJvMSsd/Fk2ZcztScnc6J/d
O2aDauLED5h7zf/QC/6vzhBIhiTBJjoZikjxU2Yj7cIn4eNypa/btLe3ly4F2DBz9d7p8Z185d/g
R8bWjp0kJuEUt1rQR0+OVgjwpyRNcyhiXZClq0ButHV3wf29p54f8jt/z6HUSXTnyN6toeCAXdaR
jLiplvHu9wIkAurfvC+MPRLzWAMApLeOjkyMcbuLB2+avUaZdhN/9T29Jwlp+aAmxwJByyrXJavs
sr++9pqw/JzWEqhlXAyD4OT09C/QUnF8ZH+fZdyfuGHKFtabqnMdAMK3MWYvvIRBnsnfFwRvOQqO
JPCT9Nfu/6rbVSTxc1lTGEb9crfhpHMI1cSNKpEMJFTiVtY38Higa22fQbG+HlYvcAushEomIWUy
W+COD5zH73FIJcU4MMv3BPez0+x7g8XkBt9ebXL03b7hXNXFFP1fl8PuUCeagnKpUF8DHZF6yYtj
5MjnCztxQ/10J1uoXT0R/YzhjLGzCaz6ewT8dEndKGZp5ulbQFmGQ3Qw0PZM9cnTFK6eu7XjpxcJ
L55HJwZPsfnjEFXTA5i2laAyDo46n3Qv+QEc7vRb+wubUThaFa6VPa+A6MslCM73H0qdS1k/9UVi
toINQ4sltRXiVjNRODdr1/7yjL72jriCsGU8rTqMgsfWNE6Dxo5GxuSMY11MEvomFRHD8fp5Lmd2
K6A0775sP4XpFwFNwl/lAh/XbpYR7smYtrUnfsXHVQ2qhIsyZpjhMM31GwY558xcxCEs6daLHAGZ
/xqYz5EDJi5DUPk/8rSu6FKyXHrHtcrHDa85rnzrvQtuJRthgdy3V0exZqbsua+vdf98QDHPiORn
kL2x+jqDRzxiovDYtJa4WQA4zmGZJ5PUAwYNq1X1HCp0+ndKNND0nmPOoRIXHVaw+SSMkdpWs6dN
JBclbyQmm92zqkdT139mieAsuIraJ9WzGftVnAVgER3UICIePKe0Cil3PCqd6+BNq+KTjsrKMZT+
nuvsE/itP7iDSmR5mptbyv//+owlNyJMknTQk8MP25SrZESHTGdb46IIOVmkFjL6TnV6tXdDs5Yi
LG+pmguvb6Wnw6KQ299WVftvNe35DJuBiK7azvLm7+sXE3Cr2x+fI4eCONiOfdfWoyIAaee6jALi
fWwiiLv+oVo9EICbqlZyyOmPYu17RAzwVISftgplsY/9DqdH+6vh4jYcJWasRKrGV/rgf3psh1uu
1ZwL+OwJ9Ri08zgmKk2QXrTsTVth2X7+HPRfvdTwXabjUf6yTaB4FoE/PByKPrLaWp7CEPwrG44x
wahHaK3UGCn1cK9UxBAaECWNnaKzS220np/5W4ZWTnpZZp857yYFgZWIEC2bcb6/KuIw0658DqLN
r5AH6Qf3HjMSytwsSUx73QG5XZM8HVla5dvVd+GxqW6RvM2Z8urbd7wLh3fdsoYOizHcYmycYmEG
LenTGt+EvuB0oAohCUR4xgke8Rm9XlRN9W2NCRlNbr/woypHAfnrgYAk2bgZNHRXc4bNExKSmuUR
YjcvCCFoUyIE+6YPEH09deHE5JUtJ/c7EULvl4ByHm1IUFugP2e031E0sPly7wO1okXUcC+9wbZa
tyYz5BFvzJVES4hHFN5HuinAeMHJnLideZ29NRum4TMC6Qw17jg6fAxBO1KhJFRZ5F46J4mXp6AZ
LfwjEtAGnczg2hU4XB5QryiWAtSkRlQldDegjJFIJyenQaK8K96Twlk09PM+s3+M1cS72m+KiGyb
S5ZlZ1wEMkHjQaa0OspMCP2XP8LKY7ha39JVk5fUksYmhqDggir5R2siULJ4JRl7vYdKJIRHntU8
uyaLGpoqj4LAw0DGqAVvQ2exsvKwxJ6woD2GjX60YMD9aqoTen99TRts90a0huWbFBClI2rhRhEk
G/L74JrDg2YehF/BKRP9Rgkww0bqAEfqW8/5AcJ23CTkMZtpOrngKhxU7sWe7IQ8u8UcSboDL4wN
6xVNe1SoRWkSwDY/TR4Q5m1rK5f5bwcDVbeAUlLBiKE0KLgQFmamQRwkFBE1FA+9DpDcQryBv+Ex
1H9+sQS2HeikHzyAxRa1A4QxSCWakRzY+cKhKS0yYCdVwjQtrAbHfJOvxafoJE89cTky0OgnEriy
swgGh5PoQtoVS1AIbkG2JJW3ta4FNwu7Ej+EPFmIm/bUnd8iBR6gFocHMB94zK4yCxECB481vj9z
xedycDlX4iFs8nGE+Tu1l0UGJRGLbXLeL/qq1kHVwrBcRg0e/FU5K7j1ziftZbNXb/9cVxW48ZFv
JndpC8pLIKp20i5aX7AIqouWKmOuDyqS604o5bnlEMlHYdHIsZXe3haq1Qk2al2bRBNSCz/saMx+
7VEh8JOF61GZfY+s2cVWjxtb4So8+gEaaY36R4AfhUlL2a7P1cjz3sGgfV61z3UVMC1DRHWKc5Xb
tbnaOUKLQoW5lMHmU4nYSAtUvy4s3h9NYaETg3/r03RFJQyvtZmaKorDK3gDKApyIy/l/AXcLhIx
WnoXFc9490VGPEdhTdDinMziYp2k5nzEfXbY/v/A+yrZyMtqCHzVJT+MU8Vei2PunEHK3+rLIezF
QtjzwjhzFWFHZX4JBUMRFLvzg2JfXpn3A1ZTjJ89aedeJzDYIC0JiO4tu8PxaNtvNAM8ivxL2cGP
SSiNJj32naeWpwCCkg2//yL6dGe4WatIvThP2uQu5PZJv/rlVnvsFoBhjYOM9FaesiG8TydRK/3b
hQTWS1qtF+vLEwC3FRpEx9FD/E5h5f0X9+8SYyJtT2zPtYwut0NvjIubFlW2EelDoV/f/U+x69CE
WCEjgoEXnSP9bfaFuRdXQKTyTlXbXHCY58gAsFAtuXK0KIhdaSj0zKKRc4Y6rMMULh8HYdvAyKuK
h0dNObgqRREt5YVZrgiy6hQP9fKqmxFWyP2J7OB/fGOG/650IfHTt51Ynb9sS24W9KnvMFDCn+Ca
NviwvZhqBtB1w1Cq4usIU19auc6aGyXtpsP4uL49/1Fz1HYoWAGd1gk9LOBFQP1GxxHls73jqccR
C50j29TIF4+dvTw9pipbwpM9vZrQY6zKKvfamboRTJbnDgie6S+h06cXovB+2zs1qLDfC6lNlRQ4
gsV3mFhu/r1RNEhaLQuNdjFAn6AWSf1UJffBKh7pp+ABjGBamyKav43RGaqgUyOESTUzsNnGPp9K
qYXYFgqTqQFKgu09JSPnkyb3bAU48nRY2MSp4/3OC11us7JFniJP75XZtmobybY64dX1qNjs1/Fj
7DnAumhylIlpAzwzCpEqKbak/QN96N3rXTSM1Syy5i2EwbiQtbcXgY6EsbWkYBKOIQEps5CBdOqX
7gB+bKNxf7ajVgi/oINsdfhoQZ8PQAWuzErnhYU9jcIxYH3h0GAf4q39CYCM3NDoae4Ox6+o6EXU
ou4ETkERFm3JBp9q5Chu3DfGW3svtqvNAwK4+hisj5SsZn9W8ASf2/yixQHsI8ya5HE1iYWXlkcC
GsccMWo4FjYErG38KGpMfvq/nk46/Q3HNTYRT9DA0fEDLIkwtUhhkEXIUyendBkAZ4dGDMTGFElL
OBtLTMI8WQd+9qJyCu3FvGRvwPjsYT2CwUTUwyCqlaE+hWAfJBP7eewYx5QG9c//qxXqjhPW3W2s
F3PGLuFnQPyxVH1P8ojuN2DO98TqPfwbBrbiDJ33Jl3MT6rj8XC1U3vG98RPg2q5jxqS0B4RA21q
PvGZjL+XVTnW2S5ecI3pH9N5x5E3IXzZ+UGQn5skhlVEyHCYGZUPCsDsnLqc8w1WbKruiae3jiqb
I4lBWAt5TiCnBR9tzctDn7e0AaQOovYlQ5AfGvtOuLh9ZmyTt6EZFMAHnBwXTsTvlom0oxJ/tuc4
O8c9I3fAqZWpu22bALyfWyH6yqCoBuctGJbSByq4KaacEYMkWod2y+IUkMjcVk2aTBuS+qAMkg8r
gzLqZrVy7ICfa5TcxaQOSCmAinizSAnmjGt/FxqENqm1cyfKe/i7QY8sAcH9rbYkBkEEWYBwbBVP
cIisHrTJzkOmfS9ikEVNtVVZs/mGd/oYkGRG8Get/IgjMewchq26gCP3KH5GHBmeJLuWYhkBvn66
Z866wFL8MvpXvqtgTzanz8p6puyvv1gL7l3+VQ7KNZ26Lw8NgMbiiGoLMH/FPfEQ3qPuEc6FWo3G
wOf3AcXKozMvDtAFFEc4Ku8dhaljQDp0LEUuROZz9o6ugH7fJT0fF9KQlMd3Kga34pzaR7V3nbB4
JhY/4QPUjLh0v9iqUHCqqPcy7bjKQQeqwvamIGPHq/qG/3OHLSJvfT5n844nfDHaocOJI0Sa8IWK
uS5Bhso5ah1w1VJddphN8UHdx6FFEfG7Rt1ZW0ViFo6psyH5/XxOEp4QtmK3mfgh6jrEJ2evhiLe
RloOQOPr2d3G5czgBBXeQXAjwdE/B69v0Ot4X9e8qVZH2t5DoJ1JUXzHobv4w8Usw8nSwRcFh0L4
Ix5Rp3ln2lvvaiMhB+XjFCz+MbSHGTvj3gOaF0miosAdgUMyzdl1C8aQv5zVea4NG/wNuVtaLHGf
TyDPSaBjeWfCUei8UurxhB4BjCFMGJj2s+enLEkXPcODrtpsfTniu7c7/KloQbklDrdtt3x5/V7W
3QQy7hiPKRVZI2v+fezJXgKBoUtwUNX831cG4bp9XvxPknHpxrp78odKqNndSp4CmO2NpRh4zSCl
+9gOpZTYrQg5O13fOFGDuGifBVZEMTWZfD/me+CyZf6hLkcy6rNDy3Hb03beKY5lC89ZfAG5Tlsr
9vtLXMEth2Sql1jpKUhm7/u7W8YMelrtvknUyc4bqj8CdLf+nkUeYxvvs4jgkTaP306LhCLimvsm
R2ut9IESrAzb9wjjlCnJl89gqKQeRe2Bac2Na1YoCQXjqAUTaYc8ldo4UxCQTXyWGw/8u51wdHQK
PVaHb7puYHYn8/caydqBL3qnu5hePp8H2mLmOdQoCog6Thqacr7PWpo9XJ+gupD5qFYXItNrk+iO
5RcWfrULC4Ou0uoZn3OW3qRlD644F27QI2m/ulnDJ/fgjXd2m8FpBE/bqVMbXGcgs0xIdtQsdcqX
Iqj6L9R+aQY55nIfOFd/VDu5JCLTaZTGeTYoYeBrawYlaUdMNLfkWDlthmsJZAiWrAPo06C0Zr0r
MHDMxpPm6k/NZYJ/noeFP3QYO9o4IL3t5JcOyQVMZsaHCmtwzPgvE8JzNtUoIxq2KY5wBPHS0wRY
OmMKMigLQqxu5vimvXhFAvrsDeEKeS/G5qSkWtvU+A1HPeHaRdBzpct60s7c14vL50jGnxNTie2H
GHKv7I810GmAALBcsI/LP8fyFKjnkjYyyxP7SK+E87WlNw4qvPnTyZlP4y+G3pvFq81eNSCjmq2T
l+4n6yvwrP5GyxuiEI9HHxZY6psB0SWInlyEK/onkPY7JOrhV40CJQqlXMg6KxE3eC0xPphmImOf
M7EQgH8w7oBdMElpOmyZpH/GTNMzXPcJa+9yE1NZH8t3S3UD228sOXkBDcjYW8eSn+CFW1SReLzb
TxZ5MC+pLNw3lNpgDle8DZtjSBjExMDX5S4Mt0I0EGCszvmnWhMOjN1Fbs65/SQtalEXqtEidbey
zNEsJhBwZqiS7lGBuVHVvrqHEZzJEduEY/ACJKJaB8KcLxtkTmqSSUH6saK1scCvdi6LquXO5fqR
uCmTR5nlMxKGuugobZBeFYoDTXimWQa5IQUpBp1MFQqFRx9v8hPNl/yKx2nUfssX39l7arf4qBvO
5964RYOlF2aMNELbVH9U0EwRBladyr0JLHsM8cQfvKyJAwyb1b/3KuxE7J33RoXZ27klQ4nWjX+s
Eo7EPTlwI8arFJB2tgVP8ZGhWR5hfeYVp4sqg0qKWfS8Pr7Z640v2rVlkGbKAoycxzYdDa3vXfHi
hDOni6akWlV3hr7a67jphXvIjvnL6LyhxHaaOt7xzToKvcJdInfMbIqThem6MRJw1pcWV2onNFlo
lQYCq5zuQ8Ifl5UBnnni6+b0MrAS17OXM5sVSBYVaoFaekP1zGTzMvtVohbqMjJlF5Lq44q5HI8e
B1kCQXKPW5zXfED22HmfYhiWe8Acc04oNBG+u0Sy9pE3Cc6+ANA9jAJ8GUO/67fGd5wgmcmu8LkX
8Rs852KOoNQjHhtiU8fDqAZ8xOzPd207YI9CIGvTHWBiW97Tq+GjZFpVOtnSBaP+YMX++2ZJGMn6
bpoEZnn0SHfTf1OGYCUaFT5aeBQP0xNb8tN1rtasIOyK5u634R+mQJkCkzGznC1RPyD8b86+mlQv
zn/jSamxOcIyixl8cDnAuSPuNs8VGS/qU2BMpf+SBNAgvn96H6VgQhYjxnbos9+39r/1llg3nHfN
h/gEQAeOKiyK4Zbmo2IbZPFhOCk6Wrr805xOg8xAwyS4GnCFuY4j0KzvLpzotbTibeS//6SZEbqO
ECQlCXA5xy8EBGv4FRbaYbdGaQQyln5CSgzN9llz7eM8NS8Z3pyXBf4G2nBG3rRHyDUhGfbaETMq
cHF200iUpQzgQlqNTAPQyUeN7Toc9H/l125XNc57zYIz05ifzTk955gnU4YR9v5wAgbfBPWEcWUE
rGn+FIVCh4JzIvTuzcvuMIG/jsPgGzjsChO17OdIQ0Ck/vgUoLiMD52nI0Ad0LsZ0XyNxs6qgUDc
zOmhy0yu2c716TPcUgQ3MqzCKrM7x0yHKpDl97AhHd0BccxkbsI4wGRoLeAu+p/AoDyg6hfyszNO
IV/2mCXU6ESkAwxYsgrS5Wysf/hrZhe6Fzq226wHVV7VOZEQ8uC6tggdhnQdAdVogHsqLnYX2MMk
W3ABP8l+qlHedDg0hgTYjtpWCfQyZ2IuJWUXLc7C6cCdLFh3NNjn9ahoOgzVHf+GDW/sLBthWHy0
9ZdiJNazagBrMdjcart14jRN/a4RXFhE0NdRfYHXMa+QvFplbGACvxFiwJWEUCFrwNnRJBxgkjLM
IxiYyTqu1WudAZyDC93gbA1PKd/yOsJ0jeiLXfsL5FDZaJ+wL0OC4LkqcddQYFb/PKymNk3kAQji
1L/G+gYujBIOU0p56QRr8qNso2yczcj8wtgY/ALlzlRUWwz37D7eH4F1Wt7BmcjIBuTSf0cWi9MZ
zXmV11DPa4Okh+KEQrBw6RAv8cvEZrO5uW2xTC+/c+KhoFsUDjovuaZZxwsggPQV30H7nmKepaUW
QkcnPSQkJEJMSGQv7/EYANR6OhHVvUvsvjeqrwSwW1pMb/kST/0DrFHyqRv+Wkp6yJELGSLtrLTS
xdJBsrxV92cr6GAwecwj70+aOekkNMBVLHjJgY9fJTpbWJDMSnQeBQsczI+qBDt8FJawVdq4APwM
lc/UrvGLDTVbKtig8isLjUjkqFHNdV9y7uU6qeb4LtTTJ3+RGjVD2WOeD4Gp7i85S6snUpLIJ8Au
eACfms2xGBbd+9BTKpRzjYpQkP+eQ1OPc6efwaNwt+lv0pNFlH9Mv/HQkLEk897P9AZOWMMLnzvt
jvb6V0NnonjAnh21FJdrmFlQ8JaF2QC8BGiYdmNJLKOhOAjrsNBpQBTrP/WcuXDUUgYU7Jg9KQsE
TKlchfTFVQsuVg1kvU0UI+nPTexjiD3htnQnTJ74Dxyri//KuakD21S9OJan/RXSPZ854ibjc6fP
Cm2v7D8MB5XieRdJlM1RRW2dddDH0aNDPn14rshJPboeN7HNsKTSxHhhmu9bo0vm6ngRIdS4XiLr
AmFnuqk9U1HLCr2CkVaevaZcp4tVNObdx+sUPi56jacoJCHEXkxy0R5/40oWPrZ509uZOfvDzukX
cHYicg2ZK8+SHfbxyaAsPY0yFjNzXs5UUGOvJSHd0MVOBaPIyYi8LOlfTT78daZTBTLLLDUyKLXt
OnzIV8I5oW9fTYNk/AMaDN/4m4lATDS4Ux00OapKOOhcT9uk0MEaiYaGYIrU2CoHpX7SXtNXWAtP
Zs4A//86XFCoF4+FSwesj9FzkDc/kbqwtQpv0PNUOveZ3pZbOQ2730zTfEYOqj9XOU51c6SFV2Ra
jHNFTXh4/BcF0nQ4yrnVNB+MWE8aZY1NJx2jxfba1muy9jvI0gtgtNgfwOdlK0F50Le2tvRQ9+2f
oOLb2Rlt4EMIG4oGn0MEkGY4YPWJgcstGmfnJ66/TiJvi5PpOj+DyVmoxRiHixKdI5U/CBg8AWOB
kqlB9eYjBExUpaUOy6WZBrzgAvtPIoOrUGLR05SjAncvELLEU5FcBDm80QcOVXPJsKO2qufVpeU/
zO92OC/cxFI9MA/g/hTmA3IU4XXRTtKb5QtSr3YC1V8ZCUzL8g+iJpKAxFy7PM5hZ52igrcMXXDP
k2wxUOEi1VmyZ/yCi5lUdZ4GAIdFo1yqinS64DltAcJ3fLNuFfGIKWNbEFJnnD+ww6ruNSaPgG+3
8rVa3p4F4bNCYavmAVNvlHhxRs5m796ycyCywOJSuVRQekL/egMT5ndeb3V0bIqQjHk1BsavY2fH
4khPX7WbAB0MuDSC5CinPwZNoJR68ivEZgftCW2cWFD8D7oC6N/7Y2Gztm3wvBhWahpziqEaonO6
qpbxUU6RjVmxnEwKunapO32lVX1cRyi8YLhOATbBhxdfEMXq7dW5GVC1LfeXoAaC/Qg1FiNqwQZh
xhVLxc4brfQXzKCMUDAB9lL9wuU1mN/+u7oyBWNaqmqrRaVXRKc9i6+kaU/QTMIUaZ1wdSeJwvwY
eejkrfdnH8iDd36jBu8/7AoTA+y2eKHRjYF5gQvDuzZ4GANkTxkRk2RuHU0OBeEJHBr+UVTnjwBa
JT1QyrXInvgyhwIfjukYZ8cO9EAPOBi7LXFZdxc08WXhbei3usEYyDGH3dTeiYBCIcwwcXVzx2Vv
+D7utiXAbXjR/5l9gpdKUyYLs2Z1kfJx9IJEfNweMpUwFUxmE/3YaAERLZGWrRae4MtMTptPwf2C
V85f/Z28y7ZZzvY3fmhlrdKxORU61iJ2ylTc+NVPeDHAphKI/7nAhlXqXVijLKTjLgN9jwOwpFNQ
rBezoEd8J1bN/gp12RWwK93dDn56MkCgMG3whO47aRPpbA9am/VNaRCn4jyK5E/VnSsQMNAKBwpq
Dqx5UrfhCuFHQSuJPDmtbGYJsYg2ry1YIgzJj4AW450A56duyMLA17z0HdgrA42PjshJiBt7/sPx
qqh6rvBdOqPUXRnIrgbCkB4Rb2B8C4Ivc3c7cOOADoIjq1edJy4jQqS4+xQV55pKIxKVim6LCm+Z
ddT7spV/3oBniD367wvwE+FLTqrGxsaNMek/TwOV1r/0mIF/vftT8G0JNQiy6rBnC0ZkpvZND9Qo
3X05L6SwI2tIGh/gpqGsSTdO3uA4Wp4fzT9PSjLu8lwpRuJH9d/aubdwB20Tfn7p3nODn1IOquHo
R4LOSJO4LV2a3lnWs55oe8WTvODQ6pNxy3ke2GYheSgw/v9XGJgoADf9TduD3cZ5JO2oBBdODFJ7
Jg6OEGzm8XPU6WNJVqKdTno/Ugh7/+K5NzLfRENWFvI3U1mVedjeqgvmxpQuXbArACdKZf7ENfZ3
wSIdASLSysH6xEyYsVaWpOvuXADdkUfF7RhuvavOjjjT48uW5i8/7uMbeQJyayF4OJmXuBOnu8+e
c7sRzuuAsDF6r/zvwaECF9GdCzqGfKpjusL1ZNGuo68NhX2e/k1hgR8WMddUtD1lqWA1IzF8TUZ/
9qX/lPWfoD8mFiCFrrvlrJWdI5/zeasScrNijt4eVNql/hg6CLY0rLADxT0XS8903K3sNQF6os5A
s6kyod6R+9XoUChGkiJG2pR3NyswYdO0iSCrY9SVZasu49Xonjmdi442JfkD+pVHV/oL/MId74wN
B1qH193U1xeXZz5XPZS+y7UkzwAZ62MMi8gkxtA1nP7ErqD/GaEnBcY5GnSueaik4g95WH2J3ysP
nT48UWUrkT7UyKYEBX8DlRsuKMm+ciN/EeBzRdD3CzBGz7gsG6utp1pMtfcLNOV28mduOVQDNUxF
yxGGUMjLQh9ufPhXv9IXr5Urv1WOcpU08SAPyJo72ymXTS57k5W6ZO4emUJRigiwg0krZ691oKYg
AdWJjspSjyqDbateNvLrG/AyUTZFYNRsEGAPGvRfBVfV5CEgAEJP0KqaGtUyNRZYhxHJAxFiAH9m
c5mL4G2/s46wRg2BHaHQLzdAIHB73zsReFXTaAssj/Nw2Nh5suG2dBEDBh2OJtGQ3fGNziJblAXG
/q6F3Bi5XjMeE0OP3DCfsBAcXtXyQIN/Hidd2vYWwn6cA2Q0FLjmq3TDzp6ktUAnv4dFQ+F8dgbV
QKfBgMMTsL6OBz6g94bAhzGtFTIoc4hFQc/zt2LWhlIC2mpEwib+I9YcFLq56DKkpx/cPOKuxzC/
4EDg2Xf7hBdZ3tDkSrPHLCPpuzFGC9jMcJRGO+zBtW7/c64kQZom87Z69eIrPzcebjwp01yaHsuq
HP4+4drrqHf9bwKaQyRZC1AO4SVo/IsvOGNknxlmlgOo9oHwuA6oXPDT5ljGixbDNrB+rMmxmaKS
Udj5lOfFAhHMAIZ1TAvfiyX3g/fg7hyTDvaDimNX6oVmkvLVpkV9q79O9/yHnua+YqeVJZ3b9SiM
0iHa6FC1YRuspR0GvgbWf12tkCNzfY/sIN1BPNHniJ8jw87dGojaPAVK8xbqpTI93RASwr/eXf34
ORRvousURnVrZr5XgnZA45SzTW4PPx73JqmPyouKeVMBpvM4oFvr37Vj8uDjCbsKWbNXtfEw43XQ
VGSG48Eagfdv7tACQteYRni10Kyaf23n72QTgwzvEsp3OfJXtUM4wzMquOmqGn3UlqoN4G59XiSJ
Nj9jUt2nrCrS1R09A1NrfMs0cP47D7l3XwhPe83pFAgU67YWbF8goES9qGU0yIJYGrCjj6hE2NXG
jRCpELi6TIggYWa8TxYcmBGEFTT1EqgaPaO9Ri4Au9BkIETmYcnCFvXUGlp+8n2qJHbuvMItzYl5
6lrQbATvWyH9RoyQ0nHKViBIHn0prUiX+URX0GHuucMl/KOcjhZrBqeVf7/whO5u1xuT4ePRoRan
eDqPZeSTihByt76yhoyOlmku3HEBJkOqT5MyJSsnImLXAcGJKXwTcliyzQfVW4ljtz6/XBaymHV3
789sBuR3awNUeII/786Cki0E/W2nM38bKmP//C8a7GGqWMfaxz8dKX+c3Ahbi8HnU6HfYv7n6/29
3DYYmtPA/UYFVP5ztMgsDNASZe7jmaTxWivTXj6VaZ+B+tYyF3jUEyA3bt/7xIvjP8e9KTwsIdtw
sw6MvPm+ml+LcJNyVONrQUiTkKsks/Qhx8orGT/ez3d8RZ/gqaxwk+PEBPORuHpZJ0TVWO/qql26
VHnJpaFWOX74qblAPJcd2Lkp/JNAkfpXT5zCrfdvncYAT/R5+dx0iO6wn3f8cOXsjrAEPRYGl24X
ZjFXyGjBo2dm7mBscUuEPwtdcrbHvz3qKDUVYOzXS8VEgRFKmLaRkJrNTmdF4c6E8zx8UlwbkJrQ
ByQgvd2vSkBeEwE3lIFXeyZY3horgDNO2upi+Oscp511kHnfHJRl5cPzldzYW89US12UlEE34IaB
w8yRnFIP9bGuHaLThcpzZHa3QM2b+7yqxWRCvXH6w1p71XclzwSrmXo4o3nUarjjSnMxkYx5Itvy
aTD0Hz/kivmF2bbg+upvBFc51ap6LuCuYq+JhOpvPRlg3KovjFXQnNcVcQvCuIYA3I/NiJIio1t4
ubOf9o8Qla9XKLo7SXJG26kQD4nmTBs8VnfCvRC73V0fTddvcruSflLiv8zRi0Sztudgyf2DZg/E
6cx/MgHLTYIajojxnb/SsR9Ob64TdrB5n+Jc0SiIEU61vyH1wvAM4qt9UAsxFaWg0kLG3UO8Qhn7
A5H7X7ju8Cuuz6S96kPJ43TL4XjdAsxXsOwIryIzsiWtgcJS0aitDHRxtwt+00Ddl8bxCeUGWcb6
clK28pnL0HtuZiGlgn7L/kLvSoiqxerDLFRvEwU4ciikpFKfLWFBNDVf+r1phPBjb3fagz7VJcS4
vbv7KEc/Nkv3VZfM4uUfFjr74Njk7yYCUuMqh9tYU2p3F1DFGF6i40YnI1AiA2rO42uF3DUgxv1x
u6EEgMPE2AiFGOAvB2RpGo3103AlahwCX4SX35N8scNNlPO7PcBFPEJEgsYOUCHCMFGb67abZNMm
RdX20dAEAVxo/J9KNoWqD7ewm6VCZquLsokJsJh+O8qhTSJ/PrP1wrLtqtalsQmtNw12DzYALxx7
aTQIN5/CRfzMlXCcqJbtjC8LihGRdczXHZ4X5z2sNokJe+IQRWWmTrrEQZTC+aq7MO/cUVTDYTjI
fEVlyGFUDZujyEc9rtujV8hPUZbWyGDy23ESpRF+25xnJZpOdc6va/obc0WS3j8NncQnGemNGAEG
/8xhtXx4cqqrlQW+qz1aHQB0rd7DaMm+v5HZIVW5gkGq/CVnazL/qMwmTsoenI9TyxD3x7/QCSbO
Dyhf1QPxZdMiyweVPafRs1xYwNl5WCmPK/p2n6+NamTtIfYtRi5HQobj7SIObE4AZlkcG9RHHAyk
57oWik2WqDzlqBfYxfTW+4j17ZlI31qxhAstvqjBzeCJJ9cTe9Rr3TC8prF7SWQ35Fdt2bYKyuGg
UK10RlR72isKioZdtKIe0FgYEuyEp+UcStmWY/HDpYCIY05j1BspQA4urjjDsXh3mZz2sa0cQgXO
yolQWMnRsQD4EkEzN1tK4tkUmf0Wg/A/e25RB92mG0bofaBDeTnbMQdDidHWfaCEPjA+heW+IL0u
6i0C0j8SRONnRtRfuFx9aOOggGQAJ54qEZFxpbvp1dMt8RSwhIH0bn1bO7Mn0DlzK/e+i0sUjAQg
EcubCg646S3yCXE9tCx5XCobLG6w+i0QKapx0hDEyP7CxiJl+WBy9+fPXY1KFx9wdED1zl47NXD+
lKD/KnETgm3PvWC6CYmMphCyOS1pP7ZYZeocoq28jfxSFMuNGRzSYaw7fULCXSQ1vhBrd1QX/GPt
s1wa7Rux3OEgGaa8aCPTA5pBrE+TTg/XWskKjabGwfoD/uQBHrPaw1DzDqZIatWFMVlFbDvpLEcJ
GXFeJjcuh5A9lJLapCY9AMy/SaDZ+RSvLAXs0FyDvUCP8Qc51xJyO88jMvmRTIiKQA5P+rPgUxA0
oO7QP4Jbzb91fBuS/4+9onqQaU4kbS2tMvlqAGeBAyR0+goEouQZncAxjhKDd/rjwbmRcT/2GRBe
7Ef49mzH2csiQKIu2q92aivMoNLrimAZekhdC2wHr2xmQYknytBsbLPAjn0PYMT1g207Aaup4IKq
WEflQvZ2pHPqlnXJr1WC39k/8as4kndWUcGi6vVAU/Ev1ra8zivfs+P9oiFD32ETqBhJ1MDIj4JA
UA3n0o7HXiLWQQiTwLwA1gsUrF8IbhCn1vM2hUPW4ClZAyO8lw2AatcqssGZ9Ob1uWQshIA7xG2E
mC9MBoC/9fTF/VlLlDJWZKNEaE9n3aGWR7EBNj89eq8FtIFBI/VswhECmW4ZXGuP/tM2XGsIgDOO
uJmsmcM8vc8CEfY6NZoS6YmjfltYuRk8xzAQxtOkt6Q20fuMnP9eHAw3aPrKahyQgiIixrcCoePL
3h9PoW1tehOPzQlZEMyOBmRd3rfUIYxzffI3AaKCogORAtjQJ3XZ9XJc62sYkezbflzmZHZ3mp5A
JH7I1+TAK9t6VRJsMwBPE1JxyTaamKng8Ix2KrCxs1UFg76hErsbIH5EaSmsJK8gJV7cxKf72Oxf
zHeIVR4In/FnK+cD40Y9V60c/zcv3bfwRjZxz5+eGcy5STbWhRRrBD1z22d6wKchsvRV34cDs2I+
vn+zQvk8qQbkpGFbs+RP3MI5/5OqAAqO3csybnHHsnPoIoBYd2rECjalwA8EUPW0lTW9syMIs2x/
B1U1nvNMn/ahGdlqHcFoAnIw22ngjKmQmZkS7pcJUcwOuIcu8Dt/edTnW2smuxez3AoNAannBfrr
fU5HE9c/ED6jRPL2yutiHcus12bHl7a5kyHCPHgCwHl5R69fWS6tJ+ew9fm+zposQTrwJFcRuhpn
i7u8zrAU8uMFvrqvZTszjSdjembJ4PCYpSQsqp4c20R+2XuSB1wcKBulFa43VkJqJSjVMHJX2EIM
h3JZSQn8Bt3J82Nls0fUwuctFgnwBmVQ3RXHfXLHXbWm0jrG7fHJlodyjBgfSdFl0qaBoo3THQe7
Uuibt5h4CubSSCG1KGIa5A5YkAoYh4mw4whiGJLGs7QYojEIHWNBiGpdLGAuPeuVncUheRVoBjE4
KAG60YSm8WgPj0CUgVEoLuTcrYxnz8TU3+zOfmUgWJKB5iJXsTaS744SDh/IlcoKFp22LL1So392
DJST1H5M0wZDuSMtGAi4cPzrOn1RfGKFHQETmHDk0Qs/piyN0cVY/rSyx+yE3TlGhtoDXqk0rkG1
Vakc5cBqupBy5ZDqFJwj7eZqEXC+1IqnlmspT/IIT8TaQ/rlV5Rf1TWdIlw3cVfeU0nPRWGfT3LN
oNdVJP2M+xH6M8TpAag3paGUbDTeWylq3ZjFuvdZU+clPTaA5iWczN3ZJ8H33FYQeCmTFr/82EQo
x29WepdHCABEJPQmDOmU/o9MeM2idAu6P+lTdS9mvAiP9qQizd4EitrHYYtIo/wV5tQVlUKdF32y
4Ak7s/JyrQJddVrMmanLeoVyRd/X983lEy3lxd5NFrBIRvQzbvSp3OjISinEPN8SNufpyCvb9eyo
6z8ma8ybht0RXcqpP2prcmK+g/in7Cp8jIVHjtvS0GiHl+KyitcT2jn7WY0PKT09WImbo74qViAv
dJxwB7sQisBvIryCVYmLeBu1UH8Q5F0i34bloP7lMsjaf5MpYp6h4dSb/zjFl7Chy6cL3ZFYZyZ0
gH1GqVtwPQZl50hvZ+2kzSBEOwARA9AXnhPcgiIoq4QoqMJs5dK4Mywc5hYDTI7QSmYMy7Ie93dq
JQ4spBkXlzOxAh3jSbje/SKvD6YgOEFUDLBFMKnTCP7ekDWpw0XsaiXO414KudplVbNQGnISWrh/
qNwFgSD6HH46pS+k+hhFNX/5qEc20eGFFpP2yuhLAEaiccBlPPnQGAnEfLz032rDEBDY5VCF+ED4
Fd/54kn6qi+zEIBefJlzZptalJwqFZGXSCPW8Ymct+ZaB4EtRuXC6bAZo0kJtcg4TWb2xrLvGWb9
WVCbGjl7hjZXL6BqJCNGyEunf93DwF+gg1iVSf3cqC5llsG9m9XwzgnAoUn+QLdv85EyiSterLW+
QeELGia15eH3/SIiPYHwHOIlWc0BWqI9GOJlk5wL4tA7mU5+8qODQMZU8v3inwYkvm5N6jYsht5R
LQoaukrXCTNE/aR6oVLYaiMpxCIBkm539/b/6aUkNcVz/E0cOLeRiof3/RfbBkB21/CRGrZ3poQM
9VJxyEViBmie/ULvMp62CHhNDxFHA0j2ftJNU0CxY64Tsj52Fnf9p2P+tjW56uqrX5F/tdwVPv0n
AqILAedhqNomtMxCH5eKm9+AEL2Yo8j2oHWVLYPmRwbwewdJSGIT0P9Ce2eExgI7G2fsGsEWQsEs
dvlfpOYJk7C20iBWJZECbWA7Cl29iW1y/0dYF7/5IPeJV+tXuDT0Dy2/EkH/Yo3t4Zkp+ngJcVi/
6KQLhcburAH1zXUga1pW/Nx8o5RL5P2YdCSluHQkT5gVT+YKm8fK7a05BtDy69C9emqgylfqhToj
Gv7L97aLQWDgRpsZbfmrw8zk4Z2J7vxPzh+UYyr/Kze3GV583fpoxtgBqb/yMWOZzhpO6o+hhnqq
J1S66pnYuQpa/6kaHwoD/IJ0xwLdmEFunEMo9UBPW496VeDECt50FiSpt1sIbI6fZbrufl/gC0+S
Q5WWaNF+RoFFJQCcFBxkkfK7LlMpXr0GDUc8dci43YI66xJgOnH82SubaBLYyQDnyJexOtEXLRVX
BqndxrXWg4WR83sikcIeSQeQfNipoGWBBEIxZPDm/xWHw0ufaKLkfyFW2WJ8vggRDSpBACJ9Gpm0
44EiHN3X+Iq/wtr+mr0eWepV+gzx94FCskviiPcC2KApxZQkp+Bax27uotsf++Ro6kBb8+G/jzQj
yCbZvhiE7WY6yFI1PUUATi0PeuXvpLgbAgr/EXCj7SGz52SvZmQ8cXpk8eRCqG9rfVKEhLDD7oUt
x5O717XZsEO9XVVHPwOO8QarCVSmMLO8h42YjpQbHug1jLzmkG5ywMjqSFtwOH77ixDSNJd5jJUC
ybmNmQPwRtDAFBHR5rnxdgIvWR14RIP+6q0NUcGm2iD7BJl4HuFjANHxD0Wsx/jJLFeCVh9twb6c
t5PWNHXVBg5HYU2xVEdVfysjk4MLelS8WYS8OfjNJAwZAXdKckYsf+a/DE9scy90cDdkIm/Ivusf
VtLtjsbRgHJV0n21VvsgkrYw3ijGrB5NloDyDnkIQCZ5LB0dMZe26P1Iom1G8S46cYE6bHTJoGCz
YiY23ZFLmWy2XCnVA40iJGsxu+u2nMTCDsHYpOBiIWIEK3fi9Z7KjsOzlfKDbKQatisKCX6JjIhd
Zf9s1i5spwRkA7+yf5Kea7QfxgkBCI8o6nenin7WhzZeu38Fc34h/jRSyWA06gy2EMwczmVqQZOp
YQnUSEO5D+57rCVlFeOdGA6gRWSkwiAi5WHqtqk/ckfHnSJCrcFtOQRTNMfPWeV0/g2XX6iupUSM
qWbaC4fheznPn7Suq6IUrtIiHLndYOWYBzim5C00NpFAISxsxczPyfVOxR+x4i5GOLebF4GRqcbd
a8QHKFOPTywwE8F/mUCx+96akflzh4LZtRjo/A9k7KiPymTlGIzh7nkDg3i39hBlBI5nXRjnJbdc
b68ePcQ34p77zemGjD4M0ak9IIJeu55nCDTo8wob+rp1baevfyuPbNkf3W2YXDfMKA5sb/Y0KuSh
Ya2rphLfQTEyTtUdftqHtaFf9xVMm5fM5mp1DNvpNXgR6LMewriyxJIYYgjLASeLbgZB7VrVYvUm
bIZh4w317SDIBXdp7+JQbDEFxKnGxDCu2z1cIDIBnh5tVVWKh2WY4VOZsggNA9fGiRbFr9V9gxOo
MDwhvzgc+I64eAAT92JT7ZTCoMJCGbfCNWhdFyjWyr6Z87rGnw0W/GR+NSQ8t6QG712hwlifb/eV
rvm+GQRF3Xq5u4zkkEuzv81zEszLq7qYMUYfkrUtjI/7G0h5Whqo7MPbNwJPi8W46QMfApDo2xRP
wdrSRlke6A8be81Sgeg6rsPlRorJpbuzHc3h7qGGr28Ndvrk0STmUzR+Ixozzu4jp2vRjQCdRO/I
LRmCtho2/0Dty/+2iG+ARU2pjWXMbEAXE0Vv90DncVd3EFbwb5pjITMrI86S8yz13lE0TyMOhcTq
jdMQ6ao0U0h0xr9G9N9Ks3ggayUSij/hA9jt/oUIrL4i5r/wFI9WIKq+NDY8nMLbVZieRyLRb67w
bpZrrW3cE0yEcutY9Ui9BaLM+MGpmDwGhSmShlv1ehDfwhHs1mRCwiQ0FeeSvzKsKMCQ3faTzNIP
5T6aQqMCByQvMfjX3AryFr+A4feO/hjsO+yEBzVIg8ME2OQOrUnaXPm4JU5CXfThuvh98D0keDyO
ErxeIwWCELsdiwnAEe0MPOzolleg+UppfyQ29WKOToL0HiPP/qDOnrb8sLni49UQsFza9Lyvieb/
u+fMA2Q9tY9d7ertGKwnIwadUj4XzEH8F/ce9ESgulqzviAxTUdsATAjJ6jp5mO+g2aCoFs6BNom
7qQ1i+W9Cho0N0lHS+0mGKEdu3kazBCgSMe3ry7sKs2xQz7yaw/4M1IbeTP02x1zV7Ur7mg1kPF/
quVuUdqHgQpTf8rKZetAaVqO/F68PZh/p2X433TWXuHt2whahF+xv/oxNOf5tBPBnFpYTZ0szOj8
mx8WAkYOGd3YfByBpYHZONJeppCwGjpQFiXcQYOozcXBb+sfRS17VUYcZtn4iGf63FzHtMi8NQ/g
RsxvcP0FLWhMYlYehUJAsgrMlLhzqNGAseV/t7fxCk3fobmqt32P83lYPSzzow/Kii/85wcuyuY1
fLrufF7Q6JWiccZICl7qhR+XN7J3HIPsz1SDAdjq8hdjxO8QbLEMmSPvOJiA7emWBZj8GkCoNV3o
OPNEWRwxPbYcUi3ZUiJxt4Spj0PxBeEtET2CRDHJdWbWDMcHayzkO8wv5CFrHRNIHIV5igGnlSIT
nGYGEvDkx4NtlFMRQLZx6fLLTHUIYPB45+3ZjseYKMrXqJfUoFbEwu1pTdkJOwcALBb/JiTEoC0K
9j6BAA4yzQiA4xVMo4wE6yvmqketnBqSm5q0XagKKS2tPRkmQkmPkLZdjaWZQKVF8pDP25TNckIy
p+WLHJom2fhdZcJf0r0kyX7mFxj09sxAMjC09YheCUnMSpuCnBarycP2hxM703gyBoDB7UWLs59R
xvo+TEX4xnlF5O6i8hVU07868+vDZoQNVCeFBfoI7kxINDG5+mnknaLrgCjhVTPVonEtEoVv11k3
fygl+PuE8PKv8mA7j+7RcJJ5i+WWuqO0x0Ua5iljkiO/BoDw1BQJYJIkqbn2GwfxZ1QCnmeRu2Cb
hGz1nQ1OUoeXAPdzOUeRaxbG26/v/n3fsNY+M+VGkoNxkF1MoahjDcy2Vn7fQZaLwVPU6Iq88s1G
1rTQdeCUnQirR6kmrgRxdUbdpv7hydb3Xzsr2GdLL/FQJwkcxFhzM7A48m6OkEsyQsRMyXHf60Wk
oPVS9NLEAf5SFFJVB3RTsw381ClB4ZJnowIbLESkkQI6HmO9N2LwBv79nd+9ZnhU2ChjDuImSCB8
uJS8S24jHOf7yCKYqewnOVwFUVju5E6ZTQbvQZDZduvYrXSVqGGhnv2SkOjdrpLqAjnW09fBZv/E
dc19i95+lzXY1k1JohkcBkWSzaiRbyBPlNKg30UZk07Xe8pQfCNKZbxgDxD2kwzsgX9UvaYBiQVX
vcqjXJbwKWsY8kUsIopPRYaQRieeLBO2JAsy3iDpSactHHnSgIn/BZ5Cs3THYSOosidCs3QCd+3m
wRpGnEUXdLA5HqOHuZpLS+iP3Ye/P9Tg1kePvazy9b4A+FOxvJH9RIuUs27Jkq4VSzkDZLzqtVvX
JXVeebCwjcYxTbV0jKIVkvMmWbe9hZPC5o9K8HNd1p4JzsOzPN2TWDnF+e1A1CoAtLFUIIZ8zcfE
FnO8JZoae3g7yfy5YKEcMZJGxtnfXEOcX8/0Bn5F+5R6dTSY0JQ89yXps3H2mBIB4rvLEHAxlKwz
A4l1UxQUGGgiVN+iq7TE99Apfpj7S1e53/PPKXxeq6NI0S1Krm4Dw1GC9m7ABHkOQ4OAvX7KRoy3
nbov3k0LeDU7N7TJKUzIuPK2dPFcjJhoWlYNMfeuvHycxbbY3jLS5dnm0Wh911UZAeDjLlLgrYJo
5dKUSieyivHfxHHsp96KNkcCM/EiV3O2u/KteN6txPpmzMxySkk4Cn8bJIV9maPJlrhbax9rE8oh
N502BcXgr1Oxb94uNQK4DBTgqTaJS57JBlyxsR2ywy8/TW1tRKiPOiDUihs60icaYIVZDGlZRdmU
XLOa3YWOy9rutGsfKlCVAt5QvEj8upMLfm6dP+apz6P/g3Ex/FG1GTJBlooW6P179DwFSH2P2T/w
F+Wbme5pBprp5O6q5RtWY2imUTBDSChwsVlhOoHC8AncCJu8opyZ/ezHcakDUFMgfOWvrr+NCzwt
AvsLT/28MUkwE0BfVJ8EvdLnaZo+vdTe4TG/YV/6KAy+RpLATfjscJZCiI6b8iLxZFM4be2eB2qA
nEEp+Ikm5kthERXeRa6pZl8fr01iN+eGWsL+JNlCyzvsbgomqDcrZ/kYTD6LhlRBpLWuYO1ROJ6N
9KTApdBTSPJ6hwuG5umCd5sJstwHVIFeshbTvGOfm2gogE7sZtsLB4O2iY08YF9UcDhDfYV5r9uG
d4+Dhvoc7Y8PhO73xln6SEWdLb8VojuMH1VsPWakk015OXZvfKD4IuHrANUOi9ZNu//Xy4exe1UM
aY+YUKfsr/sneqqf/YCt/Wvp2fFhiwGCPczpB98awj0o7/hHUEH4kcbs+GAlP91w8h+hrgkMlGzE
ne4wNfEMVU+EYsEmlpgA7NG4lTyFl1AT/OxaluYb44a2BHl0ZYG99NnQvna8RjlyHd9LhPw0xVLa
AAnRAGgRfVNAeUJawZAc4RODdh7s4rwq1Dpg79vGmic5Hh+/1L09c6C4agRa7O9B0k1CQ/lr9h/9
MD3WXw7C90i1Nwa1VrzHvDCToKX0E8g4R1+V9ugVbqq8qyxK/x9OitoFB1Iu/Ha3bMLlTeocHwwB
Ywcfkl1zawJ3l5xzCwynwZgvcffU3EAC/E14YG7WM5ntrFaJi2fLGl6h12HFpY9loNgVQ16K0bhK
6TFzf5mkH/9XScxRVrynEek93gnDF7EsfAaJnkCcOlI4IBp1Du698UH1Cvr5Xrx6qQi9HkGPZBnc
WHuTs5wKnqegS8lpVooEeOCx2awWnLpaXDWwhsVfvlGY+f1Ne02X/2O2UYXfAoKsS7kjRrfQjvvn
L8vjUp1c5whNSaGOxgiQRH15dePGfEighe9R7mJkxdYZVFYvcnTaBKD/ow4Q3DCeYgypIVx+4Ph8
z3teKTlX686ytb3TmfnJetYw6bp2JHVLPDvv8iaOU40sTJQ+2BacSF0ABAXAldGINAuCNNKhiDdI
2t2fSWxPjq/W/X8DCf73I2xt61jc8y/ll1Q3HmO3maFsKo+WXy1OQEGRYylKz0V0QlqyCypLOEHL
urtTop68metR3ccEyNMNszCyXz/CUz+nfsNtsRo3IhxFx6xe1C6udAWRCti2DjsBwhPrl8qyr+Q0
C/EdTqGx4Vp74BU4HKZqvljifapopf7Ur+MABQis84i/mYF5uv/RCO/zAK0KXeIgaliJlIv3eE6Z
oTQ2WhFZFJlG8LxwbdgvZNkXWtdy7C6arcWS/+k0sgL+Sh1rJQ1OAqQCo9/a0zyzutJnxJditz7c
HiFIn7Mkt3pR80wVTylyOcB79M+y83zftf8ESjdyWtf/N+FI0WivtdYFyR6GvABg4GbL1j6bCsNA
jO70Ky7K4wRNnHQiI97PL7goWQQ5Hqpz+YAoz9nbcfltAWYSXadMIaEC/REDgCRPFMUOTYIrIUFi
YikHbdrXLDDdpYpouh5rBu+YOUnl8MWHyIG54Lm48U34/qrumvVi8GZCS2tebciC2TE7d+hmzNRe
y0AysZjxS9MCyGFexS6Uk5H1v/a+cnscR92Rmx+mlhHCt5OS3HPFNQPM3sazfFXJRdJL7NQ7/WFC
8e9Y1CbbuEmsa3+BgBOfAAl+EXgXUTMZGJF4Q1p8ye6ZF7qI1MPd+LBIXiAZQilBT6yCRfKg9WRN
GCWUbqglqotnsSjPyQJ+nLw6ydamEPeOxKfhUNySUSLfgVIxpgefvmLUrVfoiQ5+/NDs/rfnRytf
CfNT2RSzzETNQSofsNuNPxbasZoPPC0HoUW9SKsYzsvGtrtqvoTJFk4ovu7xWRSdKvPt9/I/GePZ
1gHATQ1sKP64XW3x8XajkcHQb3I6oaM+3tWH35hKgMBvFHeJKHOR6nRU1swInZl07WHLjBFhl5Jf
iLPlXzdUZdXVMH72wzRdW6zvv8ncGNyOSIVaS7MCNbnvd5zlyY6ngTHyDvjCyke0jyth+jodYUdR
kArhIgbXwcPnj5lBxUF/82ppf1BaeCEreFm0RP2Zb3AVGZwvWx0BMajLVXmRGT0fGe5O4AECDE2+
dyTzMSnJE9uIhGwl8jidermxA0dHARFyRV+Lt/BEHLgzNulHqxlPkW46cgNbygnzX+W5JNjwROIe
79xDYdMgECezOHM5e76BYrXvatzl7yKf48LVP45WeNkDubJSbmnGp2bTMxo7hI6Y3o0+zESUGT8Q
WGbySERYJHOWYU871VHnd3Mew0e+Az56KJb7XWwombfWV8iFor8pH6dRc6u4NfruNp6ykfWK6qC0
1Wlgre//awELz7+vDxzCfrJl+UDVqivGrNaOTrlgSKl9F0fBXULP8zfgGkRRRScD09YWm6Jg40Ts
bMA+9xrakNn+IAviboo5UBIeIKScTkgdVSM1pzr3Bzp6NRE/+Lsgyy+Qhm8J7bL+YzFG2mXTtevp
F0v6DAU6EhvJFngB67jBMhZ2ZN+PfIeGjGuJtlaD23fQs8JnfE4z5Bq9r+QOZM8W59mR4Ez660Ru
5AyJjftbCBXLpE7djIteituf8WLGZr+YEUlpZn3u8c2dLAH+42wUOR0zz9Y+wQ+/SCjKdJu7cxZs
b+QEsgYJG6LI9itzFUSXyXIKChiLYM5CoUsJXNMM5CW3QaTIHWg9lkYaLQtA/V68SOZzlNURzCuR
fddsvml+ci4+17c7pPfgNK5gpSNZR/c8Wil01w7yobIc6kVIDZfc9+dN4QQTNWPWMk0NR23icbBs
TKI/LqMgHBRKZZpwVPKk7BWEDEECx9lkKDSqi5EGM3piQeIQcNzl8R9cTiCXb3MtYW3r0DUvCrdf
KFifOizGzuClbPrWNJg0cVcjEWoSPKixcTFk1We4IWYsaiY1ekKY+6sOF5vrXdwF6UNXeelcgLx0
qu3QL9ksg2KRs169MaME1ONcFOHRFj52QJbz5C5LFI4p1fduLpma7+wygD43Y5l++vJcNqVCZrq1
LJE1+wGKAOexoI/lLT2XmjaS+ts8e8C+M0dsjmbA6PtKUTMo2jQXRdUXWQMbh2UZDzz08vYakNPo
1gCU2XpMERNK85Mla13j/iok1YY2QTsd/5HC94IgbvEbm3Lgct0e1QSCGRfnqjJViIK4S7CZna0w
u4hBmM+ZgnZvk95/043WDBNJFbdNo478PNLWGFz/lUP/fqWbfe4cJ9R9n0hrEymdo4rq+yKbvE/M
4yhTgFaQ76BypsQo6uNSif7292QGRy3ZQ7WzuzuGt8loyg7OouiEhx1yA7iQpFh0QcGDvhEVR41S
koNiaMGD3YDdSIMOG0FPnIUHNQGe6uqk0LC10VtXNk1h3UwWFP7wFK+MX8QEKwnYAjMq9FKNJFcJ
VsDNqI3hMPOXlBjr+warJjb66ZsrQoPl3iRttvrdWf++XAk5cq3qJ6VTaZiZKtgr8WOqA9xsOHRN
YxlMSBq1AgWr7jHwguVyH1p8+JvnMQghofga2p2NLe5JCqUn+bHcoDYJEGQdfLZJ2UwfAGwh8rFL
nudUXb9CakDkJknNsi26VDzrytOkGpU0M2d45ibDjf5FbpKVWSIVFEcfxzU0DqMu5J4foslTXfAN
FFW+xRG8qluvdgkhA5jPL4zvjrcD4TGBnz3FkZv4CuDn+4rlgRU1+Q+n+IAJyryKanCYMMYDKaph
EOtVeq1I426pOP5nSVqqyf64MPEIH6wgXo2lRdIjETBE0VbbLxdRu3u39o0VdcRBfkvIOD1TF1dT
ap+hclr30C0bA1jVx35nCfN0ZOpEedFYsY/KQs6lspUdIvjJ35V68O5pd71/K0/kNpSG6GzNTi3R
SC2VK4FHnwMD/VLuUBrH92wMziVcj2do/WyvhF8D7TYlapYAYwnX+Vkv/2ZY12Qmosrs/xxWtNs8
bpiUyCt4abvd7/83g+CvO5vCHnoojFWwKn+3unjKbx/BJOv9ljcHUZjEWppD4eWPoL+rz73VD0RR
caAJYLF6mYM/ZVhe2xlKdXjXhbJ/ytwhSaxP2GwYVtD9CE2s+LnZWEPSfMi/jbSE2G7WetjI4BWU
dtRR6V8WVAsh2lus/hNj4u9wT6qJHAaVvclVkeUaqdB1eM4gfrRI5B38aVYhYfxhYWQACFdYKBuj
qb2OrP1MmglOMBjctcq+UIA23SbQhkgdCf8bCWK8/Kj31Oq7/Ckx0kOAndvGqznp0tQP1OxMnsxN
G1FGbaPPft/MCG9HovyiN0G/LjGSeoFELHao2aL+X3iLLIsI87blMP5kF3lcgp0BCCqZ31CZLBzT
ouhVR27ohnDbvjKJHSXMLffiTsPC+w1QijR0KjIhKoedBMLY40MN2D5EkpkQH/a7dRu7/jZCdg2W
EPN6u0qryV7/oqZYfDkGJ67zT8ysnTMIYlAcKLlN/CRHpqO2UOA3H6gqXYqrBjA+9MeIdcDNpYv5
Fy09iyrwMvnaRHlbiSoyhQNOtgBJCTLe8j7PW0vaVA5Qxqp7SuUQpxpCWN8I32z74NlM2xgZqKeg
U5IkquVQB+MAhen6ykp0T9G6CZt0YpXlFTAyGW3jtKHehpimahCfBHRHZyZ7jLHzTTsRTZ3daHl/
5QYPW5wUECoC3rJSfW0IzpCBpVhMI7HQS1odSd9a0GtitsAo967nCswAxPYLNNvVsPHsDEVsYUxX
9CsoGW5pE1ee0QUq8+ohnEpWZrxpOSN8uz0/tL9hRaULxozKZUEZpY3Dx1xIznEZDacH0IEJg6+D
SyoAgx0cWSBHYvoWSpymecBKSWyNWf9/jr55apqGXB27jwhetonKOss+6iMAS0NG989HiGhKvtAi
u/CtyPrfY9rTIvRcC86vcV85+1WhC+2QbKqh7JKFTznAzORSgkQwXFJgKVY8d9DLi8eO4tEIFj2Z
X1yrm0jjEd8frAWpTLRBhZ7KHrLoFB52bi+zVqEj6+VWS+OsnR1d91eEXsCEkcfYKxcgedXnidV3
lXsPmOhojDTyETsTgIzgDRyv+sf2Ys1iVSOik5n+IYcHMBTu7cyWJWk46Ml4KAgAIBTHgISbOAgM
E757yzveUR4h9XequNw2bGSfTPqQLLm3YWzfnEY75m7lKdHGPWaI4YE5Opo6gL1Es32zuSg1iCna
Vbm0F7CltJpnIhtLOy8JNzs5fEAptCVYukmVAWMGuq2EtdSCIZzFWk0sKXEmJCgttxmrrFnxjy6Z
KeenFZ1nUTijsugQEo6q8H7/4ITVYuJE/dvN25rOrctxVxUT42vdcS2b15Wua8qAZRuVIUa/dzqv
7Q4GSG0FSYNz7gvVxIRtwNq/jhBEJifHGiXeb/wXJfK0sbd3vMoE9W/MmDg32w27mlU3yovrhcPI
J9FBi5VLZOQFqvWPlPXtX+E70P3ygq/e+Nq1f4uzPij/kGb7ytrSQ8GgBPFtrPwbfaJrptocUvdW
+K/4fQTFuP6GQdR7OYXetozvePdd3cLPoiG7cddmNvMspq0qi4Hksh8L08xgakZ16oYjg7kVkA9m
bdwQZJz46QDYnKF5Z9aXyK7AmiVD0IMjf0/SuTKUBM0wbUn5cB43iFEE4w4rNbznw37sp0DGOp+b
2z8eNXoimtHiQRmpbXdFhTNMKz+D5SkfVZwdK7XAsOL7uDoIKV/czCaQHpgn/dvI7X9qaSaXRxG7
moJ8Z2PvxcUaNQ8Z3gkca+5dyX027cOXvcvRGQiqaYvGq8h+5mtjFDZHDOY2TZF25rzihA4WjnIi
2XUi2BB9ECJB2CDoJ7u0AKWv32ozvb3GEm8l9/IySmrWXw0NOAYkYC37ZBKu8F41NUk0f9hpfyTT
NRW07xccwaMgnkZAVCJUj1pI2kg5xqXotISFVADgpYPTlR+bHStRTjXiSYhfpNMQaE1C9E8GtDoI
cC0rbejUWTd6mgrU/MIklV2ZEBbq9NBPcI6Rh8sitjr/lGfgBHjrXhZmCxFTw2AF4hU7J0YbmSM1
91DlpILCZJolVqWDz9PPlB6EPke8+Ja0OHV8VCN/zqmCICllCvsEs1JfpVn0l7a8o7sqYkPp5bXy
AK/M8/LjfMFS1f3eI3752wPEdYMAHlG1TydquYXikj5SRWJd+HmjLqunKo+AueXhJllisltqMI9E
f/7a2ElqkT26pJcay9im1oYlGaf5rLSsRPPvvxqvBRUL1GGH+ff3Vaqix6wuAx4FguC1IhmamMwc
253eowGz5zSfXsqd3h/Whgsr2yhmEyZvclW9nlcMQZE6kwjuN0AQImGxaPNHDiXKaWhLkccOd+Bs
O54SpGT7HhdU6IBetqHaweaE16fmdrSX0Ejo3Ajlq2kgz7hZePInGwtEh6mUgmEK1xObEr8eKsB5
p647ZyTsY2d83xZB7V9xG6sLDkFv6XoVJF9oeV1VNApDc5Il6gi9LBOaH64+1y0xiuf1OCUX/S05
ywVId4UXHqHiO3XkLrvlrlaQ/UDEycq9g3cNGqhIp2b39F607vGhyXlOP2UpplhppwxroWz03c15
I/UyfkuyBJi9hhJbauGB5axQKEo53H5o42xUjpG8zScAD7InmFqkf306YQQBwtRInmQatZZo8tJO
YqbEtEtmCP6M6yrd1xmav2VxH7h2Ig5JVZuuxlnmW/zLWOtFacI64L3Ou9YOu+VcFTqq8z/UKlru
zBsE/hB3g7YIWSiazNYDSdTcrv2o14/JLJaPW+S05j/Bc/YrVf0T+gFx3XkN75c5ZyR6esAs62HC
qVftErADqGssExkSCpiazk/5PMcXblhsf7B9DI7H0nLBVFR7Vd1LIC3V9HPtlyAkxg3cO6FxyuCd
FNUYhfWNIE9wkEVMpsLVT3DZAVDYFHu0BgOS9FNrhk0+CR7z3wNqCr+aYko9dp3f4AcMXbGPt9DD
ZaGY2SkifD9vw9TmY6HMm/pcAL7LM1CXqTA0RX7DoWaorZ+L2DTynNn09AnA5wulEDLVgpfgovk9
vWtVuWAB1KDfDBGzTcxtiyfx7Ov2zjSYYji6MNpy2cw1S6+ufYt+Hky7h0CNOHtqbiAMRo5dfsbu
bjApHG1VZIpGh58DgaZoDw1de0+psXe157P54QX/3maNWDhECRvNgo8ANhvcue0GYjEWoYx25/xl
lq41El95dAHRqROLyqYOQI5c+nsnDmH3HPi7WzSDkp8VlaYkyT2j+S+stC4VvRTfuu9E3no9M/NW
QYuzWJflb1tPnwWitf8dOYVcAMB4q6dYGAzS1PfQbJm2UDk83BzJ4EUpXK89fdK5uRXYNSiszEwk
snFwGCJoDOAzVv+JcFU9Ghi/oySx3MFCAI0afaJklf6knWCp2DnAn0+zbCRfI2Tg0fQVnRn0GtRr
VG0V0FJOqXyOoGzMbhKotIzqAhXvWy+lExdMz7hszptq7AK58707Cibpwb1Qtrkclto2/OgJTHpE
XiMYL1BAkeCoel+3pbjiuARr1a2TZbLWsIZIyCPIeI+ery8KqJLzOfReeyiBc9CavtcAaYEkXxId
Pvbbq6wVG/7vyTMJL7HYYlY2/FWndO5ltpzv/mUNYK1FMwBWOh3Fxsvk4rlgCqRyhGf3NzOIdtvw
mZH2xDjKmBj5nazDO98c0xXdj+nYCO7h4Id+9XhDJ0Gn/PeLHwWwSeez3CZMYHBQON5O8d8Ms+9g
WrgiOCvKVe2WsmFQXvCaSXcJycggv7DDq8aGpcU22iIoULRPRc/PPrVhD8CXjTvRcH9ZiblyyHaK
Dl0AG9gyppIPn/7wJ0Q+qr92OiAhnVr3gD3JD1oXem4IfEEnIsxktFSheMVWrcZBzKbkBIIL+sou
JWgLoH9NFpjFtS82lpTMF7tI34c2EuMsJLkjXh8Avs8coR9TTLBMQCtNDWABlP3Szab8RoWX2Yqg
vxHHdmI5rW0I2GMi5QGM7kuTsOh6DPGZugtgBWbTf2CjmwNG6L6gvAA8NT4GjVoUaiYG5eytQ/Cg
3+Z9FEiADVNyOLoRoh4h0vB/He5bX7RzeiubSfeNazzAFjWq9kbu4SaqB/2ZV4UF1D4/wMGjyacp
PEXdiVY7zniJuOd7SkXswIqnIGItw7R3Ysg5B8bolBJzkqKAMhpWYqkWiIGg5xIcdPciM8PXFe4C
lrRbso06nrBmxWn4RPO1t2RhulZo5ZMCG9IYab4J+s9+IsR7smvbWSw8tVVVN8sfbXjc4PErHH9n
6bGjWqbuYEee7CmP5MJXt+4lhI/PvsfR/+RdlaAtI3WfWAhzzgsGdxn9Nb6GJ71mYaT+RrbNKLd/
KGosCho1GCW2SG7X7KD/C3ituBLN4HewZsrW2XrN4b6TILj1/Hul7rAX+gW3P9b2ikmnmtxrI4Az
H2rfVMZmzJ8wMmhrV5dODBSZdbIKYcmyXpJH+yozkEoWbjjw2V3+Dh9D2IuDLU4stggZZ1/h5W5W
IsBkc+QhNu8qRT2NN2yjFv4EC1MBNlGqITI9wejxWWKKd5ARKKGQQ3BG1j74Z+ZHJuVEUM7LlegY
vUpnxiYym9543BlLZ9eJOHcaOgaroPkSqSQMHxfz9bYJxpsySeicx5TTIdTXzkzujHlcspCW3xJe
MOM38qLmPaaoJti8PHjbYjjDX3wyef1b5JbbhB15wrkLxPGuN/0O1QfY3HqQCHgjLXjJM6uPZT9H
QqMoaa84gbJS3AMpiE9OjEO2qQ4zGpJItT41JtCnZFB0d0NoWT1uaW6V+6HI3tEVxZojc3Hm05TX
HdBZZAUt1xiLHLoF+DGA5KtkHEjGAW/f+0z7AEMQoOuSz+fnJe6O/qFLyJyw79aKNRROB8uhVjCt
kajbneiA0Q0oC6SHH5yzQ9HW0V2US2K2lEquDIc5woQ8fMVZy3qR/LFgZs4It6cyeI4rxOYaDhrV
PmqcZbl6fdoogb0Urhebxo4Y9hlCD5q6FhzZtdK60Ly/jAcxon0YYfduZwiYc53TOt1yY9LTCRQ8
ZlYvqyS5On/lvqdtxIsFyaVgSzPlIEB2DMzM0/WvHOOTvBmIIAxbjU6HTr/bnVylle72k+XjYQWM
bn0MwriASzSUKn2Ha19FB8CEzop8sVstfc0fwzDRLGZ6f/WEN7nnl0q+a06++0H77ABwe77BvLeI
jsa8h2I0/Gdp+r1OthSmnDbLOFalKevIxrANZXw7/rCUl/oNWKU+PJP/9HlUudja1ljr6GMhDF+U
ZBa0Ln+qBpy2LvocYv954Glber9OieKSej/BC45cgtxOlJIbuqPU/t+NZkffBgdUAGNjn18F1cgk
hlJcWTaS5Ct7Q8M2Dz7HQ38hqD+ESQUh64jKWeTn/uXbSyseT4XOFvwg7I3arpkKh+URACoC2WM7
dalT6xatDshqEAmWE+QtdYwoXSIomjXRAZx83ViCeq+MiH73yjgw385topI7sHW31qVT9w9ocY7v
w0hkJzejMOHJtVl2HinRpT+9L/Ij3SYdolEbW/M6Qr2hXxpM8YowAzck336Izs73om7QQI5C8Cbp
bRrel6jF10F95peS+4fpNgNR1itqijSPi3ANlJiH/AUZcTx5fRxn4xW5lcZtIfMZ4u3KAxaKvTY6
NNyOg3gDRjBLw18hUqvuUl16HPZLVo1s9m13mdYEW8vQpkvZgpHkVZ0bwV48Q0wtDb/gwgm13CYE
8sHGHEKs4BMOrcBXQg83iiJ5iGxXgjYhP3mVz59f7rHu+0fhsw/bpjoMVztX4cMoTxl0Q60mxP/R
cxTVr3PUV0/dzPHHLt4/rkqPIIpgW59BvE/mp2ZLd6xF80b7sWB25t+lzVMoP/4l0On0n3qRPwqZ
F++/Ij1aMljpU6f4sEea1sojjDebDLsZSUkAApee9/S/srOjUgc5qxjzZZGJYT7DSxvpvBvl6HIS
5A1snAxa4bKwPmV1GoPkG0THaqpyDtPCW+2n+buKcFYfD3JZ4vor95qcPtEfMtfjQ0GRBXMenLIh
+bUfmdYNl1y6DEzg7vMFT8ZNNQvA51yvBTDtHyZi2iAkTMoDhwFCVQFu1CEkn0gkYJ9umvdXfTmB
/Frmb22KTgSXIPydqh7kJKWznXesL+CqbHpEmnvKfY+JvpXJfU8Ec/b9aaOpLXl7tMv2bzi/rP1l
+Ifgyp0ExWL5CDW7VslKes5jnCD/aerE8Fx6L0j2MMsb0TtYA9kqypWdeTozROP7sQd8Kuh4gH7G
Aw80t7Mbrjs0VC/LaOWXg6ue23QKTI7PprwXVJ2ws6gXXInD4qaG4ATsO4l/dNwXSxrvkxi4Mdrb
ru8PW0cyQsxqOMLtWAnKabfJKCuke9AnOQpsWkIoT5v4sxu7VDRLWC+KocauqHkiSxlG96ATY22x
OWjWcQpS6oUjQ8h3pHuuHuZzU1QFkXhQbox7nT+cd7jKyVSjKH7FyHTOpg+T3bT5XgXzL/3YsYn6
ftkKqkPqwteNXELL/CiNNJaYEqDDiyvkNLQdbioMdyTKW1xOhMyzsoX+UpAxSyqmgyvnZXVXP878
Y5P3gecIqpRuA+cMq5bgUHlzNhkcncW8ZOyaNjWaGNoyCVPIewQdRCN2N/42OR8uSS6saSiKLpu3
2kJYs6k1n+5NweGp90HjJ2wycR+l/KXBO3U8qMzMxroL89Gq0MwhKSxqAtsw/ebw3mEvM6DEP+jE
pZToRs+OBMNkLUE1Gkw9LAcSyC6poz0eS/MaQSr/HaPkiGieiInfO7QSvRM7rc6sf+sPgBpS9ie3
hC3gjgFiCpKv0+jQAQuvLy6EljK20lfJPSg5OISKtUypc4Ge/qHTKy66rgvtrbcNn30VZqj+z3rO
dc9at7B6GVy1tTOgp828Hxa8JayfqmyxbBe7wyyCi4+pnaOLT9PHCjATKio6OsjSy6wZgu9LOVqL
3QxI+EAxcN4CRPEOgRqMjMUKjx0kGLPF13+O2+5RuUgbA00HzxGcYTsRi2cNQG9pzzbwZIgzyBZE
RM9++7H+dxGrUcriSrpXECIXm+n96Mcpyg/bynFObNjhPfAWFfq0I1Hp6+L0Xmh4K2DYkRG1e7I8
Lq4hDvHdwHO0DSoxwle0N6ha4mw8lOWvIbPTAlP+vMha3VqMzmpXMsQHYd0xilVZzfSqxz7ZFw2P
B62NwXqU3vOItBWS2as9bA6pohVCPXb8KcqkX0HVKpDNlpfz2RmQc29i5BtMmOW7DeBuwz6FisHQ
+Otok7Q5bwPwfWhRHcKMSVj/5SXP0Sp7mQ5ufCKKQOnnOiQLFbc/13RrZsuypJnpcIbctfettflp
eV8x5BSVJnJaMUVL8vmqwa66IrKWE5PznCAbwuixPXRZu0CCQspg2hfG6xbiA4V5JG8DJL3W3XZ1
raVZ3V8bmaH/jYPR5dwQ2kXeDEV/YUXVVl57u9LIXybGciWllj6iuVbnTLRjGWkadvXN/v9gF7Ts
mu3WoeuzAt2wvHcXhcQ42mHDnbaIc1AiwMhbUfKIGLrVWjIuLVZYAFrb2Lg/2M/OXG12oypEtgcp
TdJgJXvkjX+zAJBfuZq2DRlnzYtvYR3zEjwvJOpiFeMmmxhZkLK3INUX/jikq+6ESw2c36i0H92v
S/jLdgAZjeqMorN79td9ffpv2MLVt3FjBzLaE435x1gH6EbJBspwdkJ9pesv8s7otKfQKhbuFqK6
o1WMX+/RvOkWeaUB3TNe4y2gdNaUSyWQBDSXE25USryDPrerMMKegOF+oY6aMZ9tWYfXscHN7LHa
Mcj4ru9GGD6p927yMqhucL4dYC/Xmar+wywddlK0aesfEwtRN4mGQVdye5sOaU6tTZz3pnSyBOSe
rB4K77KkNMXn4SfH3/gCgUeXELz4vIYEAHT8P5Gz3u5xvrDS6hLi9uy9DbQNc0MT4jTRk95Peu5/
TTKfOia3sjyRoi0/qMBctVo5vPzNd16BL6WmTHcpXUnCA/KDCyuZL0IGACwclZom8PtGYKK2qWoc
nwdccQVwaL0xEdpD4wqfPWTEXpkdgaKUPMnY8xHkAEgpg1eYxLa/s0Eh0ibcTHdtlwod7lWChxq9
CNFAegM7RNVekejN4XmgUS4Vt7bodv/gkh2cq9UHdgsLrVAweSEM5zqH00LW8fH4VLLbvB0pvS5H
iZTfPJXKQkPBKNqMDs3vKL70PXP2LGeLlF5LZWIsJADBPsZbaWliAmbX/71CKBr101yMCc1+FFQ7
nxVAHLQpW3uUSC96z0MSe7z1vtzOPKI+cWcIpUTG/Y5QCuAXolq118n+weY9usvgfju5eSUkCLnu
c/OrUrAuq8+VT9fkdai2xacgc5BFfEoCJ/kqV2YXD2I06SZ47R9Hp8OXelohSv/IHAEx9eePxNPY
DijNo6Kt5+Sr4CQY+MnMW6GQhASLMEcw6RH4/rFBMMAdVqpZs3b54SQJvLAevdu9bWalmN7MrQ3+
szK8AZRK28xTTXphsD+T2xjC9wxNGzcq4dn5KA8t3dtglz7VVE6dWFNRTc4YmXGfguHtmFtTwiJI
r3PTaTMLiNX8HGoNHwFoYas9j0a80Z07tXNg9C0SU1FGqRanWXVrL+L5582/HsOPcNDxNHk5Yw+E
+eTRkQuu5bv8iOoXE6YC9yn6ccVLuteYbIzf87ZNQUYdn361Y2lVkkqmO6FL6xSd322+k9ou+cLF
/zxgjmw1DkyHYLVPKbGYdee2PvSNbnJ1zeT0qhWzY5uOByz6tgqyfpyl36n082eiy0lYnv6Xsz0Y
Zjse+cfBS7n2/TtB7GuzRnD2SiOQ8LQU58/1uiGBDWNf/1o6G2njlGlnVvBKf3kxNuxI5tcA2G0O
nILYlvKij6hc66Rl49QLpUQ2Xdtn2I6rAbeFlQvoXDCb+AhrvjjkhJKcMJB7sdzWu8MiOGh8VyFd
xaLzNDrVYF80p25uKE1an2HWStzikW9xMkBAxtI+LbP340hFupS7Gh9gzbSh4zMFIeN1Ql0vbkZT
6lGRSBsGyrvavJW1nxqNUcDV/tKa3McV/1/+NRreJTFG8i0rG3dK+5KejTyo5T2h7NNj4rt7ct07
xKDRdEQIv2os7jBZlgWJwJhjfh5edpb6diMrTQl/sHcwW0K7HfekA3b/fY72GX/bqbbTMQB+L2d4
VPOMjUqzU41OijFADNlZHpEm0zds6Gz9HPOZvuhf4Wh7QdEHhcjFLjrkgHshsGk5zhU/GQn8yndI
0IxHXXzsfsBReHIOcwAfkwwU43pre+of1XJzRm1AJgi7OeSZue5zLBDX5gV+WdpXWu6738hJYgDL
qRWNMxegGiAS54BlJHTzkz6ogp5EKTSm3SJiscBKyItVHq3F3xpcWoUME1pdeoW7AYPH+sQpzLW2
IBolCXurckOID5/yX3T994ZXEEVmsraQyIBcpahj1b1rvXjfb8cRdYzuRSHNTtMt1TVGld4Bmfv0
a7oXad3K6EuMk2BrdJx74NvAzr0qvNDoc/GCg+INCj/2g8bD7VlfxaDFxBmFr3qIU2C3srPLd9ak
Xe7yvo+I60yvRYnJ3ESyk2/6W8Xs/4/RGYowQrfeDpZujDDNZ89urXg7OM25wdTSdk9V1mSmSKTr
qCKu8vjBldwNtbZKYMqb9kcqpt/6xrRgtQDTZEc1ITS1z+I1SiECcZXSzYxLfgg4E8JLhj5MTiYt
muiUfQRUH4NWU9HR6sLoGrpRdixX/K/3/pwnAbaIgshU+l6IOKgH7WfTDEuG6tuTqFfeAH+1i5sr
0n/czVoi0JXAn+eT4KWoPQHGY68r4fkxn5lqtDRniNJhjjbNsTYGLgEvvpwkhy1niPuGA11nEjtZ
sEIoCzvASlfVP+uAsNEn14TFEpQn/BiAfQ+YBBcK+1bqyGyjVl7cCNN9gCqh5LrpYwMJMBdw8Ii/
2e5NCc717TW0ln5dc6UJNB314BvI7n2HKXKbuZh85/fVDdi/B1izdGU65kseNjb9JJ98A6cEpjKu
uW5/21UGQwwyCYfkbe1tyj5QXrNZERVX46BR9eZM2mWgAqCEgGiP3kFNYuKWsaXKWi5aHuTz5TXV
GS8Mt5qJmRvfCcuVqqZagNxITqeDFnYOylMGymZTls9vsroO+pq93FRAWYURLvmko0deWPLkwz90
z6qJyp1RYysG/I6fTBXcx9YKFc8+qfQ4zBu3x49MPbb98q8M2AxoNxIwS+i93iARGb7iFA/AAiO/
8gtBpXlvrDRNJadYidlGLnRaWIDJXtr4ASGuPdgreZl4Er3savkELnfB0pgJ3NwJU8Ln6NfZqMmh
C8NBFGiwl5GrfoUyR282UdgOn5kXh+SimqAudAr8/LFPPFBzVYzVJ5T6Y66X7Jg1ijV4XbUSmr4B
ckXNZAzRkxL4/vPQMQg7ofiM2Q9dCjbTAurIN4QD/Rzq90VZho25teUmzRc53mMhn6HutyzZEB1a
NRsX0bYAhraMxuXXxncKfJ24BgRSInMJ396UJt/X5EeE7UoJlDyJfu/o4BaIcNIcoMc9ufMGxGGh
RcjydUqtyjLBc4UF8KK+Q/93OLRyYw94Qy0yE/XpqeBk5/gTh2W+9Lh/qv7MPZSvs8qwvcrgxAWI
9ug/QKtDrD284yv9+5A7WX2wRIo5wFAqAO6MQU+FfI2FegHC5Id7pdSqYMmqiCkHmQtCzKSmUqpK
6KaTos+B5IaeleeDZGksIivWj6vv/SjEPqZ/fZvhpwGTl59R2n5ejIJEa/6unEY484EkRVlkvCk/
9QIqRWisQpzuWVNFToUjhYRrt4od2LlHJwHHiMmGNJ4I2iNhIiHhLWKfktFw6NCldS9z30lOHUzp
JVP6gKFTPieVer3ZGOGb1ZsMi11pT5DQTl4cQwwD209z52AsMTNH83d6I4tJACD4flktYKiZyw4L
Wv1Q1zhfaZO6Uc6k89q5T0w5w8fb+q9+1ELaW+7LfI3SU8aloTc96hBMsDt9IT6SP31Es4tkvazn
xjicF9ZxJqXIMYYbA1OqCFKyf+oghzyrTfe0u4FO27Tyd+GU5vYGwyylOFAfwf+emUK1oVJts6QG
3RRfQ8DJScO/XXnywDDt5oEEaSJRZ6DMAr1eBsvUYjw8vhLEBZumHVgh66RrZq4Dr2iyMlrznQG3
sSY/Pl+bUgnoj10HvM2D07UQ+MFzPaGXP9XafK7vyN+UAkt5qPnIvli/liM/tPcz+uNS5/+q0UC8
sK9ONXQ7g4MJ6Bzpb/Y7pAuiP7D/IU4avgfPwhpN3GZkGLA9R8QowTv5YnX7TW0PwWDLa2EspiDr
RhArEHCyYxYKwzOFbddOM4cHRq0neCctXvstWgYKmP5cEBH+PqyReDqrI9BOYfzG0RrV4AnsaBuy
+sNTakaUSkNbgg2Kh4YPZ8LTiHB7xx88aiull+Pw+BK3v9YNCn1nH/Mt3k9zEyiFJTTcG5hhyUkr
I6BsPMZ+YkpVRqKgzqg9gBNujaG4G3+4ByQ8+lpOgmQqQrxB4i0kLw07x+lpCiYcXn67NrrVYiUB
w+QKBrLtcvDSZX7ei+p5Va8PiiP7K4CAamld8yJczXbvIdv8qzqdtWBS1n+czTH8CfMbYaGw24DI
M02SC0kH5UszZsMU0C0RrEtS/3e4SO/qP7S0B16pZ7xsOMFCrdNs8C7altMxKrmvoDFXdEq7Dd3L
mCYpIzoECZQXZjBb+sK1QFY3DN+hwWwIw2pfUDoOO97K78DJYOIzSGiTpGkE46cgg/9wpfRJ9HLK
gFvFr7xvckCI6axTY5svn377Wo79QewuPfqXbZ9cdNwy8swpRHSMMI/FobS0NfiNxL1IHimkRVeU
YM5dmArfufl7YvUmoYOQ+tpsWVv+AZjp3KcGpaZ5BFe9/p8vb5aTrgM2bXyxR9AOwAYEYNkYNE1p
g9m7+EyB8FTfFbaJsgnEavPXQvjqNiTZc4opDYt+JqxgBjt+d3aBRPN8nTZlsnsnxDj2m9dfv7hw
gHIdpgOrYkL4u4cpJna/wi4jnwFt0rpoZVQdXpT4PKoqWR0EdciQ9/TTbCJFXIupN9MkegQwAzOg
CTjh44mANOIVm5SCx/AxPbHbS1QKomsvHWRPeZzxTW1yRtLmzur7UfXRrGzk43sJ7d/0bl4/L5Rz
dHvZrP2W6BNWy+8KOgHzjk97TZ86scXNNLklQYFuD6u0JPON9zl3m4McSQ1ObJd1h2he6+o3Vd2V
wA9Q/ABV3jYmKeWVQ0uWfXolqjtJCYYtDEvoiZXHKY/95Jrl86e/2ToCdA5V9FiGnGMYJkq4+Wwy
Ua6DRevVL/mAH4BAVK+pHPh8ANiYOgpLMBNrU5pwgDeZqW0BBx3dqujjz9aUk3INuQDVftDvzKb7
W6K9cr5GW3BNqzOh84P0jfPa2j5wK6/PEHmrQmeqr8pHEAu749RaV+wDHIxFepk/XpbhRpyV6o9u
y2CVXsdzTNmpDdOSoI2gHnX/Efa9zf47k7l58gAtmvA0ifH3SvhxeZ6qmdqb2zNanaS2i7rkyU5m
96Jf/y0d05W38XvL0jqzCgOeQChG64Qt3+yhgn7hNDzZtBvm2OU9KyB9TAa3mUWCswc4ZpGCjegE
a8qyatWuiSv3wYrhfvtoVCFMZ3oXQH2mqkPGli35DA3GDKj+nY7nmrJ3zITHSd/hqe7mTna9rNBR
6AzKsSGkj4/ciRmAI9tx6B1FcnpKg0yn36HqnUiSY5AA/gV3WNqzejSGG699nfSbJTtCqtSZV00H
cfJeXgUzfL7djT2EewX1bBgQOOztuDgInZjNxWCKVIS2awJVm0X5s+6CJyNskrxa3GwbFYDPT6MK
WCuPQil9A6Z1TrUJNwjiBA2OOyfXTdW5IhoGW+2fhp+bkw01rhGdstkg43Aj0CWapN5OILiDI/GO
FcW4cIpvIVhTJTISjKPRl47hrsxieUZnRJJHeSFqMMRoibcnyjsGHv7CxvJ8P+vV173OkRR6vbQq
7r+H5SGtRtcNB72yN+HiX7mEZ5/6oE9guHycF1bQyn8E3vm1Zs4j0CGyuOlotj1F4AbYlI3pMzzG
Q2vJmrUtN5EpNcjzdtcPIq3z4MiRCPlG81sXxhd0HCw8eJwRTcHVR6XzDAH/GYCMn1TJR2UB+jDq
s92mFuZxYwskknKo4CFFr+1EmwxkWRLkXdzalr9IA/sZS0yC3+ZbAJkX3Rhk5kaVGe3jBWBIC9b8
oV8TGEWlUC9nXACJPbhxj+/kVjA5Bbhsb+Zl79GrIXHEXEdR1srDRMLExCPnqwOtAYbQKZs8Bf6q
ayvkflP8Dvm848X0KRtgusIqBavjeja8O/XYYgYe6gL8sPTgdSLHPzrVtnzt740JahKww1BYkvp/
MTwFkdY5ZX3a2hWbigocTkNnp45RWzlxVuOFOt+Tg9xYEo9ezOfOJXYWGk8UPI91r/O06z8vw7yh
n3dgVVd1Gs3dsl+XVpm8U1ePLzl5KrSG/9Fyt2NXoQfE1owmyJU0/jRdQDYh6jFXlvZ2U8Qa1pKH
E3Vkip9cp6JKg5IEEUbk2N9HVu4P0/3wnp6uk6cHDRngBCEyrMsd4WfCy6q3ji/eL4cb1MpIwAsQ
3CXjqzPREr3d21WKQ67WzvvQHIcbOUFDBFofzmlFwuSY5U9VuNQcqHD6fEupvHFiBHHqA0Men1y4
IiRJviLxXdronZWfjjrsFdSv2oxuka7SKahshS7rpwod4wJk8yoK+RiqA8mRq0142vbeXnpWriBn
BkmLIwBEEkgcnBFfFaZT2p7lHjE3QiTnh218rwXnm/dUVlp2jvjb+CmnKKVd6wsBkjMsZxUJrcyJ
FiX/sYg1sbi4ycEY+y4qN4sGf8mPRiZYK+efCoIKpM7Bz2gEuOvVCPknTbUcq+GVAgkmcQF8UXj+
vEhYYHNj31ZXq19nHXMhfTr3xfjvhKYnAJyLcJ4HZTjrrMoL/OVDSO0waaWESMoQWcYHzPQ6iCtf
3ETsEwrAoyUU9zQ/DglDR68B/gSWeKGMP5ESeAi74L2/CwaCKH5Y7E0JEF0vDNFEOAnxoWwJyPnQ
ZqIF+zt9xDLHyQmho3un9bamt5qhb1vQL+J+IAKSpRIaKTEF6lsamB/K55hmU8K32og+Fv9wgWyR
0XazqaLV1X4YLrFS21lqDFvZnZfSGAOZK8Manl23h2bYVxVDdQewJvNrLNvZmHLZxXdyCIfPlDxT
+E2/rwvJyRzi1a2WUukXLjo3GK9HBCa8ExWFeeM5L638/hlmWeDaFlKX1ty6vzaUuRvBq4KHm8ho
CQ5vtFyIfAfDbrwg8Rc2/xeD6FIWh8+v6z40Tsd1lKd7BZ45AsscBDMJ+pUQYmRrCKSCEOb13Awh
QoWup06Y/1imwWM2cia+BK1/8gbyBMYoe0qxllozktnaHtjzVd8zNbrqz8QwmjKtQfUFFD9m2TtN
Y5hx2CNTEOC5vgM+KErhkiq/w9Tsd4JcOWZ1sEIBa+4dATDqjls3dp9V+Z4ysDuJqbvDt+rEce1N
5ySuRnUGF+rX95cFMztviWQNIsY3TwLeyKO41W0h/t4LVz3kZ7KvzKURwsT4iyfq2Itx5/1lp3lP
kFsIeH8w4UdYzkY7/QMo+7nZq6K5LlLnPbDnwIRiWWbUAH9dcFygH9XXkRfUSvy7IePAFcBbGRm5
PWwWzNP6Zzkca2mdBtw4VoM5ngtkPiG5o6K/YyHXL7rQ01tnXCWtTedvMpx+S0UrA2a1vtk/U17j
vZ/wD0cV5U+9cNDALZM11LRfxQcDRrD48i/mjghs0V+PBDeLnH0X38vgb8pl4Typ1M/eCioyvRnS
zMUiC7062Aw+L2fLk1v4iP0z6Ik06cR0L2u2J1W+x0uz7YQdyYwskXR1iLzqJWmGhyVYTyqHLDhg
lrqihvr7HpwisUYBDVkzfhh/Eu2ZOVxAQ+ZcyV/yDh18vk4FEohqdgs5xLyp9IHdA95BOpP84bEN
vJpUHTnA/RsnBq5ky7cqiZ0MCcZI6FhaQUT0CTidr3xkEdNbQMKWA2FcHI3B7JRdZXcEK+UCIVD8
izaZnNTsgnyOEBBKMVMUHP1URQMvcqS4QNexT6cLhesQPzJGY4XuawJbndhNDIP/k+Ul+V4iX8De
I2aERNaVou9xr5eYq6baSl3QQCIqk9VIaYbgeFSQsWf7nPuabm3FSnDIl75iPyk59cjHEPo03ki3
4eX3RhbkHsiTWTjqMxjAbgZvgPzjWhd5znkGWtdtrmFUo2wth8LLmTstVFsJVgzxwFD1+JUzfRYq
FUQY/3051uSfrPop4h6eVTuUg53i753b229LC7yxMUQKujMGSKwwEFBbBXe+Z0vsm+Ag7XVs7YSs
E7Hx/sZGwxjuJhGXZDjp46crkSXyNkt+e0hGIR04T8p7J6nT2ExMLgpPy0GY/9hQbTeNsPFvFfTE
fMTVNHmMuLUTqZ+VPOvFzGNKtXHoM/pCW3VZQPFBAFWTd2jYd1tAT25j/tz73BboPmV/tHO+jZhr
4cUp7sL5L3hwC2pjWMVCKhOC3wsp05K76m5jARM89bikW1kbHMmLVFrgPiCl3GkrhAPFfSFpx7Ac
UFVaqwc5Bd6JidngICjYhU7siEzieila5/2uE/kW/PFfc+uo3vWWnxcLFf3ex9+Qt4o95JTkbsxb
JwDSwc0x8YQ1fVGSd3vdQivzyG7GaxTvvrh9dVyomVa6ZpjRLxwCyGlMI0po/uh1fdfW3b90UBGL
xIcjh3l0XLI+D6T0NeVEPan77HA4fgkKdN+KMr0C2Uvstb4ygVZ/YqoWIDx8OFwUyqxhGwvSGx/v
whEofGhcxIWiNNifVdoJ3z0NU0PrnSWkbDQHmKPrChQcDGofK5EcIPeN7s/iNwVHppH29x8aBfHS
tc9/xnrhVa5Iqo1zzwWpjY9fLhOSLJTlvJYOABy5DXBL/xCGa7xCYr2DzZ93yX+LRXFjJY+OlGkT
f8ERrNLcPTiR79sZE2s6+RBoxZYzwC4r2vOl5jn6DSY3CGWJhCvDvwK8NQm9o5rVQKrI4HwXjVEy
Q3WyNGCyEvF579Rxz/5ZQ9t2I5XE8niDqFZ7DTnnxtxZaQsJcN8f4B/4bQ3bW4wB4dVVGJnJGwtW
mEt+rRUZV14eTfl+4nrPA+yOSUqLgtVlFNu766IqyYqizNpgRA1xMyuUlpZfuGN61RuhAFaF20k+
eVqhzgi135S5gLr8Rb/M7YahHCAVTyO3d2Slf2d+Vbj1NvVq5uo2M2PexIR27EfZ/MSyDdRrGOJl
MKasfHwgt1BgTO4sI0E71/qCP/IPofUhMswcYmo967QTlXFS31gdOIUuNGkiEarcldTp5LY/Wkdv
GxLqbTPGhsYDE6d+6SP04Nx699FbnnGhaATGan/TrA816F832Cv7zGGrubAOBlosUY/DGDHZ8H6K
kdC01qJWg3gsMfpuM9Qs3zgRTQD+Vw4h3ZL9V+e4oVZrkkrWa6TttiNjHsrwi6IdmBB/0gLsg3Lr
l/J4r90r/hzj1AA/5knj4Hmf4m6S+Q2afIyXS5YNi5mjYaN/nEom4ryDQwESiwhbe+YE8+oXGpPJ
3I+bR9/Tr1NME6/0/Ja4ryJHliRvSUozM4wde4tLn4yrziMBXpgkqx6e96OSD9pjnxVs9/KQ7Ao0
n/Jq7Jo33xL8wM6sbpgVxEdM0dlIC4U3DrKEVkLe4/Bxzs3w5LZI9T2OFMzprFGaT4NsG6dsXYQ4
wfWKnmxbiPhq4sxoZQMQ2Tl/dKKPVNH6QoValAvQ4wV/Eqc/IVuUVakGGZ2DjdbNuAO7dm+ibQGI
m8aCnZqouFrMQ/ltaI75uZPzP8bo9FAVKp6Uc0v4bQp4gWu4iS3xH9vr0a0DsyDYuGdDleh6fdFr
RAznxTgIfFY6aUBtjiZqNhNcxIFybEHqSfuzCuajADP/+T3t1388UIn/kJYt8BG0+Q7TLSlSQ0Et
hNKy0krHOcM453EeGcWBTKhBTCo0EmqkEx1EJXPewFAFLuwEl9nISfWEqvILEQKLEEL7lpwjSO/D
/YmdGy6CxsfEutmZeR026F/1KnoaRmzirHp1TW8xUiUS82ACA8tPL1BbsmF3urCEXLRVckjYBx/v
6MTxAsWLILMia9y30SYxlQ0H/EGAMvf/wbOMCMgxrSH/S6reH28wl1m1EPK8yA87B7EtQuSwxpkb
ELO23jnoCqGpCCXmy77CpxRU7NtiH7r9BzH4pDYmsuX2v9cIjuidTH1CR+X2acrw6AmgxBOqchuF
VN0qt7wwJ/WmRIwUVSBVFgQGiMF7/CfW4lj2k3b50sl5LnrwiwPG5p4XZcAO2tB4Ug/TFUPdwzly
0s6MpB2FUGvjRc6jVcwQ6lgC3vHvzXN5R9oxNsCsTAPKBudUoSv1gmlJJR6IAG5OS2jVVQ+qHHKp
W2QJPawDRnv4InWU4ptRU4gOMqYEVa0HuC7w4b/3YSvnQR9C6uqi12MWaLldtF/5pZSNLQySO0CO
TDNVS6sc1MSs+O5CIKPYoQ5MUpIBLFg0eY+8dFaSAg5iOaKhB1dQ6qdgBsleI6+wCBYlpxUzloFB
XiqBtiqBY+Q7TbKNsQEnMwVFUhSDTEIY0Kg1y6BmwsC2v7NRVBaF0G3GiyoReGa72bBaWV2z4nhq
ArBxoQqnWQUSw2ogCIcMrCzIa7E+Hb0a3mAZeCcf0nomNh+KnzBk1KTemdSdbmBRUbduByMqomgM
27tsgCCdRvLvpJbHZSJEo3Y760WlxZYLfz77Saf1RCmhiKiYAMUYz4DjTQn2GA8roV4kyIKk8Tco
/qTh6Do5JeIceO05fdvoVmPb8Z3VustY3oAqEyuUB69fXyZsb4Y9vDV0i4jITAZuHZ7b6m4vGvqt
I7Tmci8i6Yi+ByIWRpsS6AYgau5ZpNjG3+ne8RkdffImUPTiCfygpeJbFF39R94BnP6eLtqzeNxJ
BkS7zA+AX2JJ4yT7F4+cv8EiWuMn7WvhXGqHLQ8iJhalrxx/pAVof1l3LyRXtIMsFqVdW7KCT4az
m+XbD1JfcZ/DFjVPcEYRekqvz18Pv2gPBYORCOYI0tTouL6iB7+BtkwNdz7aUqstmUOh2M3W6WhA
qS5kI30UwVI0ciEN6TlouFm1mXm098GEEogKqT5fxftQMf95vlAUghcHaK673gQntJu/VunYmExR
uMOrEnH6nmyjRWVMEelM2t5naiUvvZFL5PmkH6xc0luhIOGK7jzIfDB/bg87gmwwCC0qq88YnTee
/nOQccpcBpSsZqgJ+6dzdc0Gjrje84eeQN5C72AEtE9TeitpEA8RlXOY4cmJCzcAfBUz2R/j1R4M
Ao1a3M7427xOK4Gf/p1MvU2TYWu6T1fp7MZLrnafpi5cbxEi8xfP/erdznDZhcL63jz8EdW3jQ7Y
t3u19CXYyQjkk8gYyOuuqAbXZoXaT/XsB1wJ6nwRzx414i2fKogtnl4iGkIwCPgB21tCeiQ6kndC
yoQp680SGafytpGf+vMd5FP3jrq0Lw/r6KlBWvO54ylAOcRyE2sTgixk3eZAVGwCzMuZioPX8CBN
+CcB6l8I54E1iQz4c2nJ9+LpXHDISh39lZ59Gef4M3Bj8DwjkK2x4IUynZknnnB9kQL2dNlDPKAo
UophJJud0ycwdokfejjeLG5e8m89H7/Cg6Ga3utVdG37XoGLQQHRzREX/YmJ4hYmiYDK2lbRKnnM
YFDpMjdB9p0tqGrxPQHFCo2IGRCNvVyfnt3pvMDTeZjBKOu6KS+4R0k0M9IaqkhtLo4MuKDsUg4K
RqsO+ZptomLXHqK6urpsQANoc1/VeSZHy9XoWFYU1INnV12jhIlMNC5AAiXr/XmyzVX10GtkV8Lp
qZCzd7PyO4KxQ2Loo02XxdAE0p6pzwkXiK2Vsk+bvPH41tlBD7R/4ysvk6nCc1I0VSm43ON3rhW+
I2JgRksny7Z8C5jQrkFOZRSobOUPwaGC/xvZN95DMkFsYuaWsSTc8GUTc7GimESZ886MpQZjbHiC
HMAzrACxPLx6WmeU4mgfzfvOwkx8PRRIkWaAQBe2mP/0GBTTUYoviyAp3+JbH2KUH6HIXywFLM+J
YZLjqYYW1S7XTj63xh9IzZqNXUhJX2CxIT0sPGtj9T4eAZ1YEzIaNnjdN/FlZIpMJby+P2AWcyyQ
JCW59K1DbPwoHBxO4qgw0XsyPRvoL4Lral9GkfEgUQ5HRYJ45fSoE6XKA/TfvIMoFyaa1YOtyVzH
Vr09CdF4vvFOSJyCrdsFVjFa8hfmSMbdsa3JL31UitwWZDEC5J6B+z0TReSwBcTC2Cl9qXmbdcJS
5PAbqaFxMx5hj+1OIz6ZnAkqQSZrA99M14a1T7dgvqXfwfXaxQz+nM5LmRJt3D/3LlvXL1b+tLdt
TSjUu0QEDeK2/5073IvGKEwZWqEs2n8QY0cQA5DA0JxGdcH5OC3qKf8FhnBXIUFKJwKWRFU3HOis
WQWcz8FtFkQgw6qC+H4wizk3r8LoHo6gyA75OW0emvWMT+WFOYF4pPCa7raUCKNqQWoTxq1Gu4ra
p4X9Ov1x9TnWo5MPAKw37ifq6q69iFzU0IhTCE/2xKl6cvlGScEHiuwkaX+1O67FT+6fNHBwbj/C
e1T6mKYLdFZGndAyOl1XTyRDLut96AZmUR347PSp/dKvPusCTj5bsFewBw/d2j6d8zqy9Fl5gIWI
LiB+ZVd5KBi6mdbVOKlBjt24uLfv+9jj1yVqkgcYZ3hfPdC0x9uXU0PrvFZ41tkA30QfX0pIS9QF
mzDebM+YY2l1LJ1aq2MStSDpGnq1v1dMNttU86W3orP1FounJy3/xStPtqhfKefLn9UacKe/H9mM
etxgwgw850g58NxK9oNBhoxKFcdAwqzlbeFEjhkr4/NqDyacjAzh8jdemjB0gkAF3JmX+oblPV9Z
wvMUtD9gVFv9zGcFt+09KTvqDUopalcr7tPV63yaOy4YRHdXuiLqt/eUyElYv1oZUQZpQMx7mBEJ
WXrCKMN63n2hG8sn2sbMnsIM6aldUQh5pIkx9JSoq5vEBHbOAM0NTKQ1ZoaVlZ/+dOuQjAoR20dG
6vBhlXwM5gdcwoQVcw5FuLyy/HIDetmZjraqhCOlQxeRIh96A9/zI+LdfC0G1VEJVr981ufIj5Hz
Qi29z5Oj0HrAPj2I6aogcATDfXCILU6whZzRSlrcXrPAX/g1GhNdsB7gyYILGLzzG4ZIxuIQhpqr
H8HukaYzGqEeeu9v8orGXdKFotsGjs4kwylBs8Gq2xGX4IkEBWHVGXle3mofTugOBCqm94p4pTkl
hPcFauVMV8aQYkbh47HtufKeyNYhCE8oxRYSh3tbVwwKdUnGH/mLHVEqBWxXtvh2wDoEUycvhzSl
7NDfykOu2xlEuJF89nHkf31yLA2MXwkO6yR8BP58zFhmqd7gCZBbdls5Ls+OZG9HOUUcmr+eqvNq
nbF0tXLY+tVck95+pdQr/NiRTpqQwob4tCcauF3BCY5iewd+4maMkw/c0pfoLpGvAfFGA7sf4rqZ
hAHqETe9VTy5wMe6gNHr1uAbZHe1/WtQJT/FyGGsyZ31U7qUSc5fSS41DkDRcqkwYKVOKssdJma+
b6VoLF+HOGbrJ8xNSTmlp4F2fnigHTmcmPewCIaMwEkKVwza1t0bD3vRTDLnzFh/CwwYm3FKgUyV
AkzzIxm3v1vKxcFyJfr7mKM9+boM33yVEL4i0pAO7Nw8ITTlJ2BhkAtFX7crF3IbsaZakJVasRTs
if7apHdV5mdNzSWMv82WkicPF24mc25crZb94F77mqxMAgV9L1t+o3OxNis4fPHab3bdINbpLEkZ
8POXqI6BDLtauBuGLEj9tHxgreYULnndhcAivQtL3shej/RJJq69O+mpnIlc076IZD7NkvZIJ5hD
XkkhogASscrbpZIlFYxHkiyDTZghae+GXBR5CH57X1X4a6ttFz08d8xuTBj956A3ABDAoChUdWsY
4v6dfQvqw0tQ2dvG412VoFpouFgCkY8zlii5MToz8R6WdgQ+GO2n9aqL0WahFDWDEKhFFHldZNmc
Mz+GvuwgIR7WBO+Lu605eQr4QiaGiYaw1mayiASKUfal9u7VO7I0jPq5V2azcvz96z9HVfWTGo9K
HKKGzO6PMGyX81jEccxbtVe/b/m/7gIVKvReK+zr/7nUGle+9bBp8/JqFG0KRSLUGmbhB2BatNRt
ojZIcV/++ry4SNw+NkmfW0fYW+kFzDW7vt94Q/14hnwDFU57uf8gk1gGTu+ZJoOSrjgVSJ4YCsOt
aLQ1S+igk1PXEsZ+Q8G4XXOQ9k6eKXHS5B1gBS0CJlHS7ttdVESJ3QE1qFScCsC8xRD/zB0547Kj
Y2wjCRzl/QFNS79/L2EfzpdwMap5fa1mRZ95Z0pK9kPsj2bCYG1nHxcblWXk+jdZVB6Ucs6sw++3
BeTZmK1ltCLXq+aTFOA3jryVgUWSLakWXVpwBwsGnfye/Czlv1pWts9nbTe6Iu2b6u4tYQ9wJ89S
I/7OsvJq2zUFA8vRX5C5T3Jrk5cjgLf5p1U7RDHpoevdtH+mkB7LARooaUawIqYTxXUfFtITQPYV
jxo5JU4yE8o7C3H8+/qpQ3ltGcyXrz+Yu/pp9+3xnbq4alyRAzFLKnAqNu6vca7t1wDhND4Xp/no
BlJ/Io8+0ocVvibIzK5xreNbFLpaQakeWyWNN9uxVOmV8urcMRS86ZE+SzD1kmE+mRh3TY+yB4Tu
MdLUqpYn7B/ksOPvkDVRi8sLQuT79l21Wc9GKqF8HUFJKlXBcENPtX3XV/kQLHSyx4bCcFPlKbkl
AG/Sul+j8c8bFR+zM2+eujT7cAxcN3/xBei7XsHeEdaQAwRxIkxJJ0uU2XXH5OhtTdGolNJr6uyC
v68Q5uv8abyGDJKpCBjqxsfMgW3CTHj4q5otfChjrS71sdD8shy1du+dGMZi8DGsmFbtGkqz4JSD
PXFzsx01rqcmzcMYeDdZtZ5kVQf2Z3P2wNfJekjkHrt8nr5mUGqnuo9xayOznf85SuDZLCEq67PE
EKgh1z29ATD+frQYDO7ggEmiDjH3684GgnnhJZIxXEezzrIVE+kFB8AArryywMCineYbi5v/yNsd
RwAXZGVTcXQd0fGX2kLS0tc+9TzUmDJ3t6XAJrQ9gFiTLt3v17WZKV51i1KmeYXJx4ykVIvLb4dG
TniBWAWZA7v90xF/+mS2hYIX1l7XZ8pT2PK8xYCkUFqkzrwgwieVTqVytNNH+IlJ7j4oq2DFabvi
CXTqZkiLYUKFW+WfeLWfnNqm11rg7FpcuznNCF1PPoSi/vA6EJPEV8Qr47Kiy5qWXFuDA03pG1ER
aBu8BCdwVpig29uK4waL49gRPVyrhRKMGX359Lg9KCNYtFLb5JTpK4cMKI8StHblLmr9OvyLzkCo
QwTxGqHPa/ufiY1AgsfkQqRDYfQdsZiffMDmhWQfaWrNDJzAtQMBIMErs/ynkv6mvJhQAPJdKXPT
t+XNgrDxH0C4z4Kdf+bjxU0UhNfM0x1JWgVRHIOhiOKm7lp/dGnZ54Fni1NzMQM3OzU5YX5ymp8N
1ZQRX4Ne3r5umXiYu30YxBPvhUnastXP22D1xQDGOkvI+dZL6N/1V04RV32qrax0pgdLABWbrBa+
hbIl/8dwclp8q4BObaWtMxk315E8x//FayzvziQo1nwn+OoKtZ6Oipx7wpz4EiLnrfyIMiFu7OxL
6N7ZMbye9xSSdJ4o0rNcmw1ZKIzwNrp93z+lFHXsVhlzmDOzlnvCEFHDmqrkWJLSOHkC555/S91B
X6QbLDf5PR5Efdi0oXY3oesf0ESEJ1npoTkXq+mkRZ2eFDWALKU4S5/EljxiUUU9511V3C8yNYWm
datNq2NOutTiaSesdyJZOnXEmv7gnHQ6wtf53OeWsISx9YKFqQJ9Tk4ItkY91Offqo4X1ozna448
pGGlJNIvWXMUAeHr/bGA40xrhzScHmnJ1dtBKtrNp//DZXR/MN2nGXA2awS9uHyyy3sbwmPVz9wi
K89p7dJSM+Ja6phisck8nm/qf74G8mVprMDdJAgVM1WEF487bvv3ik/UGwZOTiXMrVwYZ3c2Tqg6
34baJPBcvwisX4tOHX3ohJjPeSuRfDyLr1pyA+/GYIJOOu9+iB7tIt9BCgzukvhHJ4VdG5YpgrMX
TQwheGdqZXQdOKlBcMzj5bu1ypx7qpMvU7yoGfauonnA8l78e8OcRFJqNsCY9Q4HBAZvCzyEQSO2
ODezF1sdHwUur1xOZEJBwnVyVHFFJYlpUnLsxotKQMdiHxpgbHvl7EiA9Bgff5ic0c/6VWOp6LsV
tqpKyslkTxq4SjL6hRYtuCHhCqSqEuPLAvNZMOmLsxl2LQ7VzlRB41lKORJ5S49cZQglMZsJiVve
XIHN80Me+e/HKLSjfzvCTz0sTROFF2oRSx04n2Nq6FGdg/NJYRlEC3jd79y3PiBYdgURzEZtvbRA
LiXTWKLaev6HYheUCu9rsLrglcat4MupuLp/zVxwog5KzAhVghadaK50NjPVaPp49RIAkR9tv54Z
Rhf0CQxKKVfmxXiFqUcPJ+tEXVL7zuhd4AAunaNwVUmQ4bslTXo+nO/drJ9Cn0D81kNaTsLVvzvF
ePJcqKjxWaj0TNK1enkA3R2PMA2XQ+cMZkrqPoGdyMn5LxQmD8cBGASWPEIPqKv7Lcib6a8+pZwH
1R91/XQQvnfPjA5E6FSlmxhbTpIcNtANXsncEHvyyNmS903ogBX+DuS0FdEcVe5XLSi/WwvBZZg5
R8yq6pZizn+ARgz9owUqNgTgMno8IJBcUi5Bl5/jyTNGlGWzE9+A39yHMXBS46tOvq/ldxms6s7e
Qo2Fb5AvWQAxd4O6BjETh5wn4Laxxm0ooz9Hwjj054x+2sRLXxlEwzTq6AJNtttWWFlFgKafgjSA
TY3G0C0OjwITLtw3OsVmgE3N5Z30NDYzXFfwTGeJ1UwSG1jO0/KBxTfHeDGu/EcEMxyI7loyeLhB
lA4JAcWqOnQ4c59bfS2K8b80BsCQYp88hxTneyy0aIhHBjfbvLQsCUi0oSkEWVQaa3bvdYQop2Nv
I8asfJrtUmLpO6I6uZ3QLuK7FypS0dVDEgM++TZi3BDa4+qGXx0ZSxqkCZ6a5W4DgLGD6L8+R7qs
Kcrx7elnVhfLosmspKKFvGf9yhIEGmWMcoUwXzuGYhQN5zoNaN8t/PmqDm4SrNnIDQ6f0ZiVgnNH
sy1az4j6/+4XulhN8MNnR86S7Ql1ZX1CUPJnrTy4fKuUESbz2rTPXGPFMhaL4SZ3XToQmqkXs9jv
QtCN6TRTFh7P0jmhu9lgxeGlRRRllUP3OQ+vDsl5v3OUcZtKZ/jdftPMMIOmuejl2MY4y6GYn9+d
iBHCBphFWQtfIWLgnowYtPs/BBYHhrFBQnvipePITh/XaK9aYr6TyxQw1g6D74jsNQIkOdQCtPc0
Dbwt0b+JCS6pnwfrUuAXOyLEsWEPpMgiKagoA2cgEY2aZDuQpmm8OqeHXAlSer2rZxpYY9Q0F/Jv
11vA4q8dXpnxtm0RSeARrdTP54zwaAZJtcH/7zvrhVDHhChUhU7FrTfmbgB8KcfF4nLwE+1w4xeK
PJ1+9bYKJw0BytV9zeDCXYMA/0usoQyE9EEHYqLZ0RInFio35K2dEeNgnc4+6jMCldVW4HaO+fn+
41ucUn7TCaEsA0b4FI4zS5wH8LIT4eSRcrnEKvw/4Z8ZpqqmVWnnHLgxFMdaWdGiQIhySOExrWUD
uEnmCPWSOjpY4cj012HmRsauyQx4KDRH+jELVMy4rsFQtLD96jQUaTaF1WL4673uMcmHRXQiNiLg
E7owU91uFMTJMVGlD51SzLhiwVe8FV4Lut55JNqKt2chI6v3o5l15wA5pezbym0haDyCeqINbYv9
/AFE4gYeQOugGWnlaPAdgjCE9ioNQVWlaWWp2YlVKgPzkp1Pav16ujL6Bx7ardR4wObN7q5KQzm3
y09bjWfsz+hUXnuJbiBOEn/u9EGtvuIGep2vDyrMr/do3MHpMysX82160i4Xe+B55Yj+UHLUIIKu
x47ZWoZolBwS+zUC+2hpELi0JT+pHnwUC0cDwszOqLyzqd4PEVRbHlgyPUYoBD9NM7XIbyscZleH
tmboAzhCPWL6cmrvzmFwbRbJgziilKmdmPidfHk5wunCkemDuSJkRyjXY8LBNFAmpxG5txRQHl3i
HTKqhJg8jNkCPfo58GB3NU8pCugthNgWsWDBE3OqZ55xzvhu0Kt8DgLxEP7Nse0wcnKSrkEr6C+Q
2fDmrL1b/2Asb+YKKM3JXRwGeHV3NJMYi+Mgd+VH+PwiMUcaTeiiI1LzDUYQgVcCiXYJnoaW22jS
T3UWLrgHRWDa/cLHBXf/1f4N6CIzs5VFStS8n8bgGtWOd7cDs+My4qYydWgiNVjTNULRrdM7vYuQ
wMNEFUc2WINFtsV+gDcLnNdedLogxZ8lCj4SUEBO8mMVml6XyicdGWCp9QLwIj927drTBbuG+KAn
vd7sfzpQlTopRM0kB7E/i94IFipCZ+avUqjZXg/LVtFuJ26F+BKbKQhYV6HSY1qvC6Jh8/5h087f
ND5bPsBUpUzU2GVwd4CX+SS0QMpZ39tqoOd+M2pLuDI5SmpgW2Gd6kXjkCAVtlnmTSPZ5wW6HklB
fL3qxgmNDX8TzIH3IXMyr18yykk09jd8JAGjF7j1cnkEwGNTtFBR82dnicrUxT+ZDcJs2Aeg2lSz
RWA+qtxQ1ZXINQf2Qz8J1bnZgik2jczjYrhPOP0btuO9IKaea2ktzpq7o3pyo3eAA4Si9qjm5wzo
pyjoRnRv7se8VgqhfNMo2Y7DodA6w/WzSiO3sf38OCneaSskfb+sOmrZlLAolgqdFM3zf+43b7mQ
7yppJQNNG1OaD/+efk0KWwen1RzL4RGOYGvYO2yR/iWr0NOtNNHcooJKYwFj5st71CUP5voUqlSC
TwWBIIa8tKwmegs7w8wp/IOy5RyyirDFIXvD3kmkMpkXIN43CDcaO7KiNiJ5gxN7uMupg/sVndfF
kyZEW/O+v1zi0nGEetaPjjHxx/X8yRpDeDi47h+mkN2WgxPiGyQ1lG/sHdN2DESMsWuha7FrP1Ua
Cmtwy0YYPWVqLaFhdOauGr0ohrJLCdFHgao5BVdLzEMOwmtPTeJNIt0wiMpbsM0O6pmoO5Sq71bk
kM1/xJxaGkhVWMZHXk5WTee3x4xrI6mldKRLOypnt5lgp0ap3poTgzBK9D2eGDoi6emS4gUwu4N4
zUbtt/CZOvWSLCl8621i/4gYuEa6ZhcQ5jF1HhiticYnXuRCckVa9tpeVUEGRJSdhmHCirMQCpx3
zgjrlzCGRPysiz4lVGMjQ2CjT1X66S7ElCSDREyFCpJ/rdwoSNOMSnFlkxgamSXvEYbA0QJrtOgE
JWtQBLeloJV7YXz7vKq5LdGXUBzfd0kek9Q3kh/j9HTU3WLrQKkVmTUzK9WOLhw+ZzfAtKOIn1yB
YjYFFkY+KpnDOXtutdWuNi2s+hJZXoJ2AXGQm9+xguE4pxLJbIrFlxc8nTMHfNF92ThPtV0KC7Cw
AZUiskzaYLT2kxVcpZyHjaTQ8H4WeDaau+4GIvCvFk4GhPFJSHoSiA9NWi6pufeFTzSRHfGmd760
HsX9STGFn7+bT+VrXR85lMYtdLbyqQdziE1uQcrBXVmyK0TA3kgxRN16kpKcaIBhEgxmGjc86QRN
V9S7x+cd6598r1Af6FRpxOZ6fcHqwt6AIpeDEl0+j9mkZ9nQtZfWZbmBg5JulU7/ePPnEPtvoF+J
nwes3wSgHV019rk9WCDj2sgwjXP+JEp0YxZ8P6ymFrPHMv/YWO1UjyUoud5IyxpSG9qifE45BmHi
AHMRN2SSlZWV4NDl7rZy4mqAqHuxatCcsIagf0GjFgouaPilVpmTgUyS9HwbEbc+5XB+FjBGNuRQ
fNRZG731PaaI/h2otGj0RrydKOmg7H/t6XhdElNb0JOGsVnPhI07GNkUmln7spNUJljgJHs9KNdh
t1V4ktYliiWBDz8yLvkQ8f9fDzaQO7SsF3hNYQ4jem+XqI4DdayrIhIxZIoe417uwhRaDWvo0HrO
BVc0zERMrzN6vZGRI4r4JjPlsQEenDNSYFnNhnyUWhTYVKhcyTblsEw7DrVaN2ita3Hb/S2p68Yq
/pijJWpcIbhLaK5FpzkUjcpoWOq60KOtaKmItospoJzwLs1aFtTN62NPi43MmQvkiLB7gJ9dLBwR
ojd5ZbnmR2T7LAlp5ZyJwXesen8n68PVK59KLr5dgs16c0Ci9Na+wK4Nrm5LxNPHX7QfWnv204I3
3nTjq1eS9Uxi+R48wsYorvWWajP8KdO5GHG7IkdN3vGkiWa8RxD5TIFWz5hCD52JD+8prxkocM3e
uy6PxjLqYtP6enwPdAC6erY5WW1bDEv7RibJa67ZNKWWcJ688cecCbmA7UxcGM0UwJ8lRdZqIxTC
WgdDZHPoWbrHieMGSSYvUfVvjbXfOr3an/GOp7d8tOFnXnYGB5Oa1zhSOJZFFdYjFOmQ+hLkEtYF
zLfdYNpjMF5SiT3wKRikrzzZe5anzjar3CzBrEgsOnq1LI4Z6//b/F+hjeRUXx3wwfa+JFynGEZb
mjG8AgtlzqJXSvnR+hdE/66cErfNd14MrwptqXocqZij3jJn/LGK1q83EYYVZA5lp0gIJddUV1hK
YR3n/3xp3omwnoq5ZZAxi8rsju3+IVN1bEaw7QhOinfL8PmuS7dzR4mV0OFDL5AunVC+EQSHeD0O
BeBe0Bw/evRrfr+w0e/6hwNOu2Fj1PkF/r/NjQrqcZi2OMlrQUpiWBd6Rd+3I6mM/QbB1g0rOa3K
OsxpTnUKCw8+ho36tUtJjhRe6h+PPB/ns/fZhnANV8+pKAZUVoziQg4zi+ujv1cNkGd8zAibN3tV
GSNr4qZCCgumdEf7VoT9nJX2vWe9laVbACkE5gqxtOS20nnOW0jlD9ckE3be1ZOHj4qfF9X7iAd2
gMxp6EsYGe6/wp3giW7SZaxg40Z7cr6EIeIFESvRtxTym03tCKO7EUmMNiI67R9iuoLPkPXJFR8C
wuQw6MoogFBxXMhw+e2m7mg8KiWMpMZqf1VTqtslITWl/eR7GaEymuZAe8tCD/zncrGFivmKH3er
P9lv0ZEqmX02NDd5uHKC+SIv35r/pmiiEsSbZDGbxQR0RliNvcfm3DhRDSJ5ic6m1pR2I0Bxxwqr
xvt//wr6TgvPhYD9Jwrne8j/dzLsBB29G0ekLo6Ca2JSi3qwFQg8B163V8Bs21SWcE3PmcCVZGgi
oNT+T0UghOtwLx+bg3RPNfpUo5AM/TZluDJQtx8ShoVid71pwyp2ODTKOcp+nCGQjZlK0Jhhxg0M
iuxt3gR7N+d4RhN3yVWqvoqzHruyTXAGZQPsD43j0uChyxlQUr+/ZkSN+AQJ888inLVUjw4Sn1z0
KSJH6YWZB/QEIbjMSdxjFROYu7dR9bWB8mWmDA4ZuMrayD6sc/lqeBSOvaXu/nXRdmi3ShhyoxNO
+toZy2hI89Fscwx6H46VSLKQPwUakMk60cXNMqLiePzeQEVj11usSnnnYfC0EYGl0LV0MVEYxU4c
ITJSK+Le17kMgLwozBrh/AtbAjXz9zqPAaXGQb8b0VGzOEd5WZZTormdRGFh7cCZl568jnRMZWyn
bMYaovKFcXv3/oMl7Snz28ik12QjOf7V+BN+viehdf+5Hl3nw4h932IprZZ2qEGfO7lXIqkQ/Zse
UljU84VK19q7fVEpOSYSLRMYpaSwyWGTrGUEPUI/spceDroBaanJmNNZFgCtfTGd/nOQyuJQa4IJ
LAe5fx0V/bH8KHKHV7MD0uWNgOU0EQxsG8yIbV60wNOtcggZgwWPJlrjP9wBu37N7KNYNZ7KEgCi
W87ln9ml0T+JWMy+tPbe9lv+zpMQ8xPoUbKUtdJ1DPYiYmB+B3BzFUgfK+r8OxlLgq1lOSaWEg8I
2IbuWDeqraybYs6LTGWa/1b1p5tnbyR584WCcJIDFtGjVhRb4li7c0CH27ZviYLU77kEcSB/2PNC
cDbNKNt7O6r7NPYos8lN4Ae24v4gULv+jQxfnjlR4k52j+EZ/ezFf6pdX/sUXud6JQPPeY7lvZHV
mtUZwkq8IyUhxeOMLDoYLN5dcs05M2HLYRa4e/XM9ri6gUqgWmwpdIVnCEvXkEpDSK9TPKDbxbkn
JTa8VZ/gGYa/0fYdf8ebvWht+pE+m6/bJYbbCxQh4SllhOzV/jPBzXb9bkQRvhIrPKOAmdU37Blb
xgQPLBkCo2AqyvDM5Jwyx3rOQU6Ldd2cugW8dSN0s3UDhQXWHlhQHxQ3bqGS/pry/p4r0J5RajaS
Y3U09LontFLYxzv73i/h1j4NVD58LLx1jxlle609Tp+ppPGxMqpRXHUvlRe17k2WcxCV7ml4Vh3g
amfRsTrWDJi6hUPAfkujp3K/ef2nWtzl8aD47cZhaTMHltKoUMpG7XDCiZSn8AgHyPJ3xQxPkS0g
K3dpxOZOEUQ8tBwVdfYJ4x1D2FrGvvixDXs8qbjilo/RLjsVptdEnfzaXnb5/MUM5dLAbcHkzdRE
wleuIljyv4E+5fHw9GYr3ceQvC0IeQKGTkQeJ47RDoOn0dCUqm+6uTyAggXFkKT7S+C25tvczsua
U30hesuhhygb9HweA1OOoiRYmaYrNQlENOPukidriErEK/c/VL8uTdfhlIbENFnIYVx+ZXwW/MqV
K00VsA45th8e0XtSV22AUenkM+m3Frzw8f9qVvrMh0HeWfJeSvcLcjkKDEf4QCP7xHHcF5EyGrBU
/kuVP/RNhBtFKRIbDL+nNfOzZjzhK5xnMzjSAMOf0rZAyOUVI5/KtKlgKEz9DDsfkBFCqu9DyKKJ
cCnOeGzfA5DuG8K6+p/4BB+YQyh3FEZIUHWYfJ1v7jlzGA+e1D3P9OAJyB22ExPygDnNy/uHfzCE
AdbQYg9p01dAbA/CCod2S1/D3N/Vo1P7HvREwbOlXKA6JznOu6Hx4awQzsmZ7t4NHlmSEYOfQtVP
Mtl1coZLcDOVLCRnHkJlPBICGwpCor1MDpOuljHfsKT6aNNSM14H5zWcEIaIcsHgGK5S1kl0OlIw
4aotfi70U3JNUNrufJ5QTKdeeJnlTMOFDGICRtMC7WzlnOygrsbgOzTkCf/O47LVvxXEmJhwfnUM
H64DOtKboOQcBeuijVW4sZoiI4AgRaUcYkO6AdKi52DBUOuLf3jsyiOm+eSf8Ab6CmY8x3g/j3Ri
+FAT+zZNp/QgfCS7pZCQ+J6EgIEn9GqdYiXnUTf+VJe3zxUm+3kajDV8YHybc4luqsvvyVzg0ODU
mXhV08eiUietgt90qkkV4kMypD8pg41CIK/2yNAbjilsg6hIU4bhl6su8a48oMjT4rmRxR6j9xjE
jC6J0TqKpqzCp/nWSgmHAZ2GAVHR01AgrxFEQ5YOyNZ9KBIH+pn9ZfW9Mi/+JVkdcYbAzTdKtwv3
lHuPFSq/xbk4Y3ewINQBoAw/9j/3Q6pKvFuYN9z2KnXYBxI/5+w9MOLaf+ScpET72dTAdwhwpOYr
nfmMjLb2lNXyYl0krpsz+b+gQdjaUxB06SjLUPJUnPIw8GQ/4utdKTwh9TA88X6sJBpJ1N4z5M2Z
kAUNwiCiDrjYl7nJQ3lTLwvKUvgcxJyBBxjkBjcWfFsVVD4wnMD7DlPpkXNsyhTHDj3wx71h7vCS
KOH3Rre3Dc0D4DAtqJpchluWTRPe5ImEUwOh6ZgvLAEkH/A7aFdQ8c42SA+BXF7U1CA0EMKNPU9j
FGSQLjtEM1DuM5R5DdUi5zBxkuCE8zR0D4LrlZtaDNp3brWrrduiKZSpTbVGnri0pRL32XXHvsXx
WeaFJhoxxlFfVl3NEJgun0MMvB9jj7NPcAdvctr70952lhaRVcsM+uiknjoxpiv8R7neXX4jqAcA
IOS+ADcO9PzMdtEiBrRzFnAvvsUxjwqmfrAX1Ck8RLt/NnnwPeZ+R1SQ48f9uIN9TQ+YDxwa48QS
Cc/nC2VZouo3Cgp0I4i0ryr0V1OWeLbuhEq1rWYTvSBWJWOJ8JJn5eecekIbGj34lviYBX9yjJU3
/QhwlcjhUZtMHRBRbEW1Rcq9q35Fnh5GOLuvBzXZnZzNqBGfHJv3ScxUZrN6bz1jawSiOPMZqi6K
lJSbYDyRJuqoCapeX2T4guzQTfUCYkqP/H9+9CcihR1U+eEhR8PlRHs5yKiMJ+FLtitCaHrRYsoQ
4pIYacl5NQq/vF16XcwTLnOfiL/+mexXZZP4q5T+xRK7dCwupqK6kQPhTSD1F9K15vqiuSOuFz4C
+nZyeeht0zlG8kFgUsomJgD39eOSScDogGkrrj8JwpOr/rVMnSvMLqPDH7JI4i20uyz4WcyHHiHc
7e6WHG2Z/2ADPE6O4A0ZvLP9c7kfX3l9x1qCYNM8uVH5E/RVaNzPRBULXBPz+FB7VNdnWPknNhh1
28L/9IEueEjUog8s7rBpDcM7P+LH5FzL8YXgdoUOX1wOq4SkiqwhFqSUKRtvBavtB8L0v6ffzbVm
CuADTniinGOSUTzslw6VPX5C/Nw7+qrAa+0DJQx5TwJ+ZZj7n2uxRC6l8px1aW9hDeL2i5Cskhpr
mvx2yW3U+3jruJA6Ptr48q6yxAc8RgO7DBKxabddL75jZjVQ1yRv+HlCgE1wqg7O01W1IIyyk7xY
KHoCnzCUyvzy1QSK69rzFzaTAfxj+iC/hvvQtY8FO0qzPgoIqGHRUS3kFkQkfgvSx/SjpyoGC30z
6NfYKUZMqaOriM013ObCvCypISJX0pRom8GEMVI/rlLPU27nuLe3k6fREMUkEVAqc8jfT9MD/3wu
YCEFap+XB7WWp/SasyWEh4nH3kyBSFT3aE/UE6i8lMRozw9kdImm8dzrRm3+hDCsz2d/4TfkfWsS
oypPTSbMmbb9wZzwNigrN+iP6z17FxnIKUItGYp52D8lmvt2wFKk3wXc0fcw2sRv2R3uSsqEChjO
EQIIbQquST3RTfUNxYjRmhj9sF2cDSeCUKF/9Kf8RbuXhxvoiOr/5P0Pxx/rDGG+y2BjtGFlQxhQ
tCbYHCHuhz7AXN1fJKbHngOVko8jOkHsGZnWwrDgPqBwr7JjjIxPTacuKGCijAfultxShxZMsI+a
5QL8j2Lrha8zQP29Q/K8EXgM+G4VU2M1m8L+2l00Pp853M6Ci3fRzwLnsWWFLV23N9c12mclUQb8
bvwMpbUaZnDqK87xCB1Vo3s7BQK206LTLGWLloikXigs42jHqerjzmge9Xxqkn4tUrU3cxuyE8Si
Q6YDMW6OJOyBHmkYDIIAIVg+sGN5yWClTPDFwrVE/I96L1+nWV1ST+F3oijmxCEvS3f7CSdk75L0
O2UfvoA8IJk3MNHnuw0XujMq8rZhIDEAFM6mAVNXFOP1DWt7SAnrIPr++Q3SFixOe1ykmwR6n8BM
1FevSbRjzk2JXSaPWNNbOK3/6ogZsDgAbx/0CGqm7ObiSMSEyynD4b8N3SSBPIQ+mmCux8SY+FTA
e914tlod7JcDBoNZK/MvKfh6E3vh1OEH1uyuXGYzsOXMchKg/yRe+UCafXaoCX6b1pdQsX/AvH3k
TR+4YjttfypgfviNd18Wck6OimzsooRQhvayqBLYa3YqRQyA+z/WjWeNq1SaS9XiFFPkOJDtekw+
Xbl5zmee6OITMJG3HMO7gSjbJhO/jnnE7a9sbvdYJ3KnwEtOaZOWZbH0tUoznpjh0Sb2nVxpX0/P
jh73aN9pbFbnruZy2neLljqibmyIv0FRvau9a6NEXmGZ3wKhDl6OW+16KxDyMxrwDa6VXUaaTcDj
w/p9UfAL9UIV+Xti0AKeEd+MnI9WgN4rGSL7GU5R6YiaMxu+B2UIeHEDl08X7sB2qCrYboj3GspA
2I/Rp12tNLLNBOozeczz7EMY/nbmGX+0GByVYUb/hbyj3kei0XCwFLmciZD7AGPIB9k//gpSnmC4
5+9eNgDeVGBj9SXnWxHG526pBIYiFVx5VjN8p1KZ3rvsMF2SEYELNrvgi8bUIF9TDOrXfCYh8YZn
3pXD18CroaGb5hXq5F/scUKe1PHWh1K35P7DCDv1Y4fi4XmIA7JeNvoSEGM51PPH4sHkv1n7SD4M
CmoQR0pnz5Uv+VtKdkeIWqFlQntX+7E9Bl8k7Fgamek9Y5J9EFbaX7OGO/UI6ezTWwdAkrbVC7ai
/hePakow+hWTE0r72TlZn82DH7EgdwNvoFe5WZogqggfbVThtVwIa/lm/Qw9zFsVDmgxg4h9wQVx
lEjJzYjZHvJtPdWu5G8WlY+n2iAjWFu+gr/LqREfEWyBNy7i8YbCeBydbH5qFayCTSFJ7mcZ3RFo
4MUoSJc+1NvvgY/titarEnG4tWyBDDQicfBGyZMmOE8cdofUDi8mMyzjAVMO56dtsbJG3fGLLyG2
HAUT+2OtmDakEITkI3hv+m8JKmn19b2ixTkXYhC2a8Xu3Z24yw4So/fZ8aLzn1vVpvndEd6MF80k
wWiAjL1p9GeOuhe9/yKiPZyF+gkC8hoPc8fXIkHWNibyfCc7JkocaV8qHFuUsCTtL6VkHxwF5rmA
lTtf/CfD3rzxSltuBhyWZo3fRXpMATuqHV3BM10JRyB7W/fuQtugez1jrhFiVyw5BmJpaKJ+67ME
bnoUIouXTwg88ox0xU69GoKXgY4FD957usw1tUqep/+LyIwISbwJjXBQ838p0tfruVlAhX6FRWG8
6/Bjghpjcs0LG0u6kko2TaWlHQro0I6l1io6sRd66/mnz8kZvHiRW1EG2IVkcGCcM1W8bOVpSf5X
GFyh5iOLwEiB4lDjTB5w7UCCsc3LLI2mvP85QslxUSeESq3JJFpcV73fcTpC7G0NGoDJ8I+c51Qd
bCu2/zYC9twGau2O/kn3/JMWbO8Tx30+hWe0cxoYpSXB2f6IsOFWaAFwBMg8sZMQoh+iWdT5xug8
G2VYTa5TNxI924tQe0CWYJeNMQRBmcVdVcwjuprPwV+62qkHOHUpbNtzD13TL4ZVoMdJxX0/Tg56
KT5UW/Bj89fJv0/FwEuKlcFfLnIP5uuD00+AaA0fSsYInRUPxFmJc4kp+yteEnsSGYU1Jb5ha7oy
oTadPUnCrp7l90XwZx3zI8dQUKP5odsC7154yaB1YSpweZNKfwrEtqEs/sPP3vzp08Csh/9bH7uK
6r2YjvcuuPKqaT2dxEM0sGmOgndZEB+yqmRe1HOtkT2BGuDcyN2wmpuB+hi2g78YJ1Py8JQtgIDy
FVz4hJIJuIdhh7O5FjSXPPamCneqS+2gsBeJ0VoJeP9+Gk+jEMtWhMd6WdJcfkQ2eunSR+h6+TFY
O/mEDXgWiv+saRNByQhc5D50zcooNMNMFvttHwrCgwtMud23UdYajMmxWLk0FQJ777sioo2ap2v4
oau64N9FjZKosFOJmr6EAF87F8iGrF0ynvZdXQx/cgC1SVdI8BrZWf2+ZhODLefK0qVT6njpDKDa
rhwXnaDEMEgQ8+5fodWleNCoz/ZaJ/Z6Jb6vtf8iWNBwYtUGoI5IfBmQYoaroDH5L+zHf8+OtjTD
ZH1mGZNqxsxSeo711djHADYxUUaUws255ItzHnNrcvKO7v6TWV2Y5NU3gJ6/OVkaehaS7FBQDh15
zlRe0DNMLPCSAkq+8yX4KbCidq+yAT4+8J7kX8CUElWk9NBg7Yw1gwpF42Zmc3uZAvD7wakLB/r0
UMDm8EWakFvSq8J6ij0wEh+5Bf37+iA0RHkPf/ng+Rj5riBUFprZd/WDi8m90/rxiqtj2bOdkstc
pge0ivlTRiHQHh7eSHU/5ycBOsHEhqJsx51oCcdhrIjCf8WR4fsw8f9EFXELk0lvhprnSWJVEvfi
4DVco4hQMXU78ciDbOje6mXawK/9rPL2cH1O8aN4onUwyzoWsMtXplvZxDl+mh/hYqrnJ73VbCFz
8AQdu5FJP2TtcdJEkuB0G1NTBuA5w6QLJ4nxF8w6uzZxP9mRz6NUqiHkVH9UMOoF4Clj3+C1RoYK
t640LaQoSW6Y5M0hHrPfGgP+gabplecSTbULO8RflvlW5sJJLyglWW5M78HEjmSK5rHvq1GFRSJ/
7mbGBCjn4xv45mZvtWv7w1IYo4EB8TPjj7lIuocSgbXyYGAGBR1eX+/cws43Q/Lxsu1tZetySiVI
5ITpe9f7RHHg1kzjWFBxRkCtxn7nely/yMI7F//maPe0YsDj9tvuX2AdwBxDacebI3rw4tDV0VhR
RpYutXdevvvLRMLuS3xjOkMlzQXLx9YbEs2qbQnt9/pyWgQi20GRiAJdfyAH9FXTmsAybEIQ43m9
K3/jT5lp6hRQHTdyvK7rRHZFSJanYTbiFFEd6cjqYKuqscfqjpp7EivHSLitp4rhRxgbK+zaIwoj
s3lbKLk4nOrigukvxgQu+DYk04xazkS5fqGH2A7iY9JVyeGYmONErx03S5AuRl1wslROMypuKl1C
hbeZUIJuAb4RUyP71DV5/0geedM+6ZyzAEI5uEWFc6n8EZFgnyXU6Jga1gpyz3+emiJhxWx3DLC6
NzJhgHbTJb37nans3lBqrWBpBYDh9EoZGL61p4fgXgI1ESyfPF30Ug81is5OcOMGuKRLUXgkPCZi
VLMcPzGctAV+486OzfowEbc9B3ORpc5azkhVMHBTp/oqsCkiHGrsdulV6uEPIW6LGG5dnxh0yQsG
tgRCrK39nKo4JcoX7CVWW1kSasbiMrtPVOaoRVGcVdkJ1Nn1bTj8e3dUNoyyw2Ay6z7G1724ciHy
LSkOFqInhiWt0mDhCFhw7XVlqdHtPzZkG1NA+enkILs8++j/HOg5DIk/RB5VeYGZj/ewOvf+OQWC
dznED2QOasHPcTZsnl2uJ/qgKx0sUA98//hjHpZyB+JjviuR995JExCcC1RiYKGUCpro5ij0q39d
iJ0VS8VVo9l9GOEcJVxSmiZGwQ8HPB2/0QLc4Oat1PQQxs//5Dp5FMROsVmvwINbaNYjOn97i13F
Sp0LLhED84PzNizHfWh/PQO+D5Ek1TU5X2bf9PR06JH/dWFDKzYpN/IK76MFOUmGGJxNs6ZhMmeS
gzEUCdf4La5B4TN84v82ia3I4+X+SQ5aETyaVdD4gNU5OAAGfsiOGolAqywyOlM5yrCJrArC38X3
cFiyko14V00W0GgIKhBSbwFYdo/Doog0oUQ8eX8mbx02A3Hhlnk5+fnk9GC5Nef6BwLs4aiBXpjW
GNPEF7RgS+CaTocrJMOgGK2uwten8Ozmhk1FV9ZDustjtDpat6gqQ1w3zLtH37C+6pW6u0ne55/F
TsdSRDv2au6GJz/YdRnCfiKcYAB0l+e0//TNYSgUW9g/gmb5gPLMlJ7E52cTK3Y/FZTD8K8TPGDj
0bcdot9Ylh/9AQsDIpPx6VLHST9bKN2Jc2hl+E4+Rs9fScoiagLHY6ID1/w6rKNFjdKf4utMAIAl
sXNDIvCegEw8DVcWsdqH9jKoaPELIPPUIi53Fg+74Dp433DGyQVpzzoeZQe+qy3FKn5w2HwPGQVb
Dzsr64sjisATJKjZr7INAd9VjNQ0lpCuvZXAtSH42k6eOTRhnAj9bJ0ZJC3YeoZaulNjFoWAqmm0
NhCfhzaWP/IIU6ioGFJNoKd5YxGliT3p8zTIWXFd3mzlhgTrGCmvNh57cT8DHJ3C4GfQSlxtnxuf
exYJulhz0BzVPqti/lpkJr1bJllf4qIsj62J74XZ+q/kI+A8y1rQMySe1hIEE9x3DToKhk7BiT09
wWDKw16n33Pm1kE6x0eLoYy7iPx7veAqK3BA3L9l6uCXjP1gFIsPnEwRzHN16V2iBO3+f/HV2ZZs
P6LgqrW2AXrJr9+RNZO95Vk2rpNp7gF8qSBLTON35wYsjBBUHOHqXBx78XZJhRID7gBnEwX2gOfn
rVriYeKE6lmXbux8qK3XfGlpKet24PZWkA9zlwWRjofxyX+Ng4Z2epoEWRvCrbWbwq4INkqMUun1
6ZJaUnY6L3HNfWt+bdPSEfZwD6gGtRSDTpnSwrwbq57EIQlc8uWLyLG8uJjtLc1+lvf6wYHaBdR+
gCcHymkQYjFZIdSBeF3dGxLR2s81G5f3j/JtrSrqZTyRbhEbC9dLXbDXSFbLe5qHulZcOmwaKZu/
/wm12KIX4UTS7rVs3seuV2en8gPMgl0L3HLEmy10sgeuT8UeCXQ8lYsZAxtTFOuYnq76sb+vLKu2
BvRSnHUnw3pKT4gcLxrRM5MWFwjM6GOs3QL2ya4MEXhF/Debgk0gwNNZdNPY3rkN7Lxcr5FMILzg
zVrf28fBSEh5mlaQXgzzISSQujM5+UdQx3a6JWK/9ByejOWLDLYONaBFdnEc8+F3NDqyq2bGm9Xs
t4epXO+DT6sVU7xLejuWlvVYB9zPpBYRZopbmhDfSXdiRZLjYOJADStkHF2y1ZeUcckKpf7Edluz
BRjJNNMSkHEJ1DOrK+DJPt8nHIvgF/irp+tukgvNzkZUYLkbPIOn8Hb+Eh+Xcnv3zWpdMomENjrg
8U3WzSPry4lsK7I+HfpknzQkSTeiIDB3UoL81igOSHbacJumR/C9Tin1UQKPFRdlwZwLuHxSfwuz
iB5nVMXkSJSxpnt2kGJYHejvzupC4BCd+fddy2gMEOvMiqG1A6kudAH+1kg6iGFCYoaJJxhcRAjN
6yIJXy64BOZC/jrdOySnYNiH1nuQZu7O7X4tQeazRZe6BX8R/Zr0m/79OXPtx6irb3zYWy51MOQn
5H+LbdFychu527xvDI75wXWKKPePPGWlXsMVU6g9rB3Gns0gcVjvE2KWp6Lb77gjdNRm7AKMR4jI
Q8jN1H52H+kGqH1sAl0rpJ7lpkfnEhOgPMOovCqMvL37RLy1k80dnLQb15pLAuGh8u8CmoVmEJUc
NNsugn+7eYNZpQb+8vNEjknzx0bniYlBDe0niyP3Wwp2jiYgw5+qrE/qNCGG1hUU9Bs9eODmDZBk
Wzhwg1ez+gut1FkRdZK7o8c3Fh4INCJMxrZ42JLNETm6+/8A2/ieOZXjcuAZhvkYiUpUooFctiIQ
Uv8ErzQs4zDMEjFwFcBWYNed7Xg2GZVzcrYxryl1yNDa/hjE53TVTzb48binS566XMpO0g1i12Cp
/w0eDTitt/I2raZxdojR9CJR7V6fTurJRgOseFsAfo8Cq27Uxpf3WRgD4MQCC8VcLZMkm6H+LilZ
5vDoFDM3G5lH5/qzNY54n69YSFtRAQMJB7obuQGOBpSMWh8wyKSn1GPi8OIvlSUCxyWa7w/jQVMS
eUYZWT1OHXEd5FCmCjpY5gAxEMyM5U8ysaWhFPp6UpW9Sa3Q3yc7Z6TD3mi6BziXhgzs4Tz2jMRZ
xCSdnVTfWC6LV8JIyfyY2LwRfi7baBgZBBs211A8UBSR2mBaFyEgdVaGxAghfEQCzGkEJ/HbzDTs
Ir2HPRfEuXhs/QCHEVL76D+lLwUGvB94vCUOyny3pTeWVkykIL9Q/GvVJDRYo+6wXactTEjbQHHS
y6ycvNwXFrooyY77jTdxoc0WrmXsUZqqxU8nGJRFPECL8AUTnRErtH3RvD+cPT6wFVoDIOZ6hFqQ
n5SXdpscV88qLHFWf7NC+s2V5hrJpRbmVcvwSwMYwWgJdB0zM2wrs096c6OPf85NBZjcBHGuJLbz
veocvSsXrmU3fBLmTb6Oxj9ck/6h0VSDoAoKbF73ranrHNYA9Hkye1tK4fJp9UhAGz5XLKteJGQn
uxKsNnty90qxV1lIXVfUFi7DZvFN2Cs+mu4/LoBFFp4SNT8QN9xJ1oyWfqZyNefUYRGVe/gMSZO8
No8mzL321SoarXlJ0oH3KjanszSGSsoXR1boQylaWLVf7Lc3tv0crx+VFiJyUYbBHFZI+EpnUlWk
KrIO58tju0LTBJUY66SBMuntiMS/zGxOxqQtwBryBNhA1qE6duDuE+gyzuiTa2ikoX2O2JPPmSph
M4yG7rpYqBvQjGJXtTQWEJRY9b4xsy8uYUaxaudJ4NN4oJt9fNtQ1OTcCKCWZBtgWULMjwM3LWRE
J3BmULWcs+pwqU3aknTyyZN3I1T0Sv02rHRx5k/cy2fNsCPfVvK7F6AgLd7xm76S1Tl7XUdTlR+k
Nx4Pmu05CdQ1VbrBtnw8AmS4yh9ZZtgPp15L/X4w4HYEFedK2A23PG+IpdbIvMwbdeiqdNL/LsU4
rcolKBaDikVfQbsjbxrvImaP3nLodZ7uPWxcZQlxdqEwNHTpOuU1VhSfZmDZMSOfqFlBey6tGGTb
7e5YUYaBSvWydHVOz+bVdXvUIB8lfxrBtyEZUxQ6WdhKqtr2Rj+T+yAZL1+nfGU/4Y/U2oXL1nkE
hoZTsVM5V1MRlEeQidnErAMuY8vQUP3DswKsekdXf3H3aoGcxxfdq+SJW8+ISyoI8egZKMFoMEaS
ocMx1yUhzJw7+xZXLh9zbcmynvq5jaIblBWAvImcbyzjLbuZ7TsTw8pxa+jPwdE5zw5EIUzizBV9
R1oVKj46ha9X2ypp4IRz7FJB7ebB1ULu9Zy2gVtBxxXu4xDuInZE+XMJ66jfITNu6W1RjmK44mWe
U+jpxxLNDxIvOZ/OatxX1o8PEP4sHheiqJyRFwbyqOUnrJ8VlDH9FQLnH45uh45Y0VXmYM+mmM13
rqT7U7jMZIidzewVs2um8MqdUhsOTbGEP6HUvesUxZA2/FGrUN9a+iC+njWZTDQQbzhIsbFUAMHq
sqcEPsr/93qL/tw3F9VwNxs9zZEcRwW2GBaYTiuHnBJr/mQy5JPtycRhEJqFKHgAcpJus8dfxn9F
tGc9aSqBVyhKjnjgW3PDtB6IrHEKLlzQxaWWpiSSUDnv5olDfrHjZaCjPJKLi7SYHndsXIWEigkE
GFPVPWyAKctfwhgIMjgJD4T1QS2efUWVJ8WWmOwiuEBw+XPJQ12nkvDzwVj3GMSpj//zxpPrjPxx
8tBoAPNHktpAGCpdzaEL3D0RTq8XYE8nbQabAP6xu0H7B3SCQpLHvCUwrbUG9lWcoJG6FOfvZ7mk
mAZEIOXVnq/3w5Y+lKkXCsGBGiJEwq6X9o3NruhzGEe2TQBFOi30Ev00dSpEfhSepemGqEuoOL7H
fWVDqo2IbVF2904/0Z2P7Mii54EpvpWigre/g3ygXKefYZPEfUAqkEVmvExWjESzxsg7dxkex8w9
MA4KAZskuWMMD7YvAOgc3M6g3/K6tK9d+RO6sZk6BZ0EN64EUUm2ioWnEEfl8k/TbyafF2WZS1A9
nvFtu+OBrueishJkzY4FI72Nbi6P9snUzU/daARVbJjSvemJFdNCPd2MjQSywQYpHX+HuzfOVqyA
5YXp8tTXm6R4ra5bzCJsXgYl6h/BnmT4o/k0rzAWhdTpQGcS/bAgo9NBQujOddz8ENzjbSmAnTBz
Thm1Y7UWjYBTA2xy6AlHURhubPZb5fbWi5cBJ4Lz7qRgQSWk0r2T53wH7NR3nCJPiBIrwAg835yp
ZhH3YaNFbyn4/gn8i5EfB5zJZomD6i6oWj77gP+MAaVFccdC1/8uol/s03IgGdFP5DEUsUNnOPez
fGp4lFVcxRvQmee2qvj1TKJeTjMbQKx+cwJVzU7zROIGlzdHaZDwQFQC7p1sCf1N5bB19sYCiJkb
ZkGIVf6oyi2APR9G42bclTcoOrimul/U8hlHQCtjRL2uizZ00YMQLVwZCGRqQzkoa/DnQgWh1tvv
wRYbONYzv2hiUvnfWVPeS2t08ZpixAg+CAoQgbfpHS8D19k8eR//IRoIiIkZYW15V9YOa3YG96wX
qTzxP3TbafNS+w8Bw0Q5yud4XsvNxuWG2n/4Ek8vKBkzpEgs0gbne57hUwPn0iCtCFaFJicpbFzx
pd5Ob/zEPPzciJmK0pWq2EYcW8OwzuyNcoHOq4dkB8KNH/0SpvpdsLiJnM1STnLh8+ljdUicrVaw
oVUPsIYs0jnuacoAzL/QMV40cRXII9YvYvEuzLoh08JsqIdijpOpBitWgjYPXMw6PrrkNrh9Npie
CLB01tbUv1Ln4XTZde8+zs2e1M2n5P7W3k6A+yTw738HFSYBY5fYX7TDqtkmJ8J46v7kgzn/mWHr
C/YOHtCpdhpaKqIpoGWbDanbi9yMnq/meI3kynzFcqGItbeyjq/jt+wFIedl2yx5tH2n/hTes/so
vELMLfl5LSH7hmomAgivuIY7hD+3ROYBuyf9xjz3uuB2Cw5pROvjYnqfkndhTFArZxsPY86kP30m
/dWHOMLGfw4JBBPu67XFK9eL231pLpzxyPJIlcPq7yOwAFwJ9MvlP+XOAgrQIY+Uf33touM6eqk2
unqnhxuDMOm+VHPYIpQRYO8GQr3N+QC7tHaKqcLqsLXFOY18ewf3qTwb6VdqDn2/ArNTJ9FhitXt
th23GTAwAsEqtnfxUn1qU/8O0zsdr2GAParP1V9KRbhkSH3fB7SixiJRqTo33g8r8P9C6IaNwcgQ
Ieedrcr8FZxpGoIR9bZDyxWF4aJcP8sPW0PPgVB/FXn7Y2tM54hKFQAYF5w86ija6OhPNGgfbJMs
FTPqpPISMMQsyMSiOder+59g0U9N3sliSL7otAle+2xGk8UfmYTIDICdHAsVnvWXL5LW8AaGXRdN
Oq6AurVBMheg3iSmUgzFs3ge7yTVnEVfd39yp1M/6uYSsYb9TS/xXVjfs64gMZXYesLRLwF4aFsV
REXEQgVuMQJDt6VPbB6iQ4asNDDH5mYbDjaDWUtzTkQPDscC6GN+j1ITVmQf/jZhUdZnmioTwLCd
uklqB+K1elU91I45//o+Z8e1C34ay9TssgJIpxZCqCPuhcB0T4hhDPaV/g4JuFMi57C0j5e7P+Gc
LMp/c86oKGaZ9SgLxWcgs2LV6F5viTsUIPYNsM96zBmSMyXebaQRLQgW2fH9/AvJNeH1kPmg1nOI
MIQq/1EdrzLhO3/RpPfGiMwYcv9mEOnXxtIH9ZtQJM7pPJQXlc2GuRqEzHoCZOfyAHylTiqCrG1x
+Jovym3J3mC0DY3KzMlbi6znnBh8iqWwYzk13sXI0N4KOUKI7fTgtsgN1gZHbSSYzSWX0ir679Ni
15+9fUdZGTiTi6SLw7dRTwqb1QUpC/G+UyFuyPyDuUMDY18c2vfTHS9lBrSQ1kztt9WYD+MbdyXa
J0yImyc6gFGlHwnmMPLepx+6oky051wcx7G0oOtpb7av2ZCSsUv7i95A6ck6TA0x1hDLBeKyuL7S
k86Tf+QjJt060vkZbmmwQKwfiFncyYQlZX/qAyzA+pQ9Ijv9VgxDeT9U+g/HTX6mU20ZH0WarNKo
1Tg2S9Jjo4X/cspJ0bOklaVA30O0jbeaZxIYN9lEOl1qr3aN99hi5vOHASGKy1VgPKuaLC3xvWzU
+G34GmX5bruTAdfc3A+vZg8c/VQSVK9w0OH1aoeOSTo83Pd6JzwWcJfQ5Lx8DviNckm89jy36aJe
HPvWr3gNLgT0TGZk5uNE2dcJbd5P1VoinIif8gO0A3cZYmmkb9tkEVbZfPOa5FRnlW3fY80ZTCHf
tUfvAFGhIV7DpfKk1aHXhPqcWp0VnOPlF9V0T/Aqko/kGSP+2YV6/7KrTVwcJgxl5a1bBvuZfARK
3udoNkm12dGdKkt5iyxpEQBxBO4WK3tH0o5vkh1jVwi036DHnl8wkDcsustlqzcFs4I9GOH8i9UJ
Nnlt5XTi55cZ2ofpI8DB927X1p/AHMJ54HkTOwPhtXxpVJ1boNTCA/WV/KAkAP7/p5TvDL4M6L1k
tlIA3LuRkkmTwTroXUq7RmA7cUkj7AKbuOfdGv97idwOQvWhR1RgqXWiGCYe8p1b5e4uVKK0JAOc
E4gigvmz1a+1xAb5tuLaOGB+SRNnBo+Gj13GEtfFco+wNPlSf5khCANjkN1cL363vcBpBKs0k8of
yb6EcHydxBKJvPtN+JYXmR7qOoFTYtuDm5kz+d969EqkJkGycLvoWolcnqS6OI3SCI/65ChMtnOm
jX88xTER+RK2D3DvGY+nL9DCOao1MP+e+Gla8xqLvGkYD9N4Ojzk0j1AueGZnkXOcTWkfZpOaOmV
ya50lPKEVZ6wbYPoL4twE903R2SC35ECQxv1UYYe1cwX3XLI+PB139d50JFub6DkT+CZ4Sp/bW1D
oWn/Cz26bKomaSIadkJAQ6/KsXKFafhGBzWRe90gVapE8A7yhcC9H+uf7Pu8QYStn2e2+vid3jYg
X3Ddsivb0+xVhy71pYwO4bMWv7MYkZa+KvrTxzq4t4M8/uup4PJe6E9l25XHmfnf1zJ89Sr90VP5
294AVEFZxysLBYLYpTL49WGYCveUmyKHRzjMXK/tf675xOQT6eKNkpJpsj2z2Gp7qlD605Y1B87s
XVuoTYLPFo1vsLUb7B6lPUBJC2Pw7dNAc5NcH3ev6D+wVPh60RUO29ru13kReM2omTpzTzTjBwxc
Cf+pBlFhdhPY5YQ12rhIL2wCF/y+f0K5QZ/PyNM412tB6kH7mTVeos84Iv1/VEKX8gigFSlrfno9
S63Zci6QQllr7frgMtIOrcABJ+qtGGGmudlECLlpY+CeWnKQ850k3mBqQRVs7V2l7RzYiaZKy17R
ydSa4qmTDwb52LI/wT+uuJNXxpM7qm1oNVVXpfxxZBdBR90CMkP5Sv1vitGkk7r6rAx9od6reaJZ
imQPsiAs8CWQm8FQV5hhoydHTtGHpoId3YaGhjGg6l6/NViRt/UXZ9lwqK4bG6geEI/EzE67rD2Y
GQjkED4HYNxAWkpMvSceZbDMTI5PNp+z+aiWgrJDUUG5kL479W1oC0iczqNq+eUhubPofBGOqiiB
H7pPBV1e3ktX2ambwymD1U4Lc7KorhcS6fO4cXTg4BDJfOOj9KhRvQ3WdO9CShoRlaf9NkXa2QLw
mdIQITDW/8jFCQttEFrrtZY/x4v4pgbAqSPc98yL6hnLhvZVZsoDs/dp8JRpSOO2qBw9GXO6c+CW
GgiCXn/JLya/880AEGCgnWjJHbQ23uuNUfzUutCgsH2pjGemRLEEjVCSkgTWHRr/LFz3NLLCaTdk
q036gwgXggAtE6E2iO6CJYjGW6jorfTPgk2WtUSayOLMKevYY0OrINrcJSfKwMG8Uom4sf77GJUJ
hBqzUOJv1L0FqR//7bQy0viEuGInChtiICQaIf3tiJlukDyiV1ZgGA4HCSFUblz15s4oJHBXnqYf
m4r2rZ/nd1wJQlF4XtH5y0lqLdI2vpG9b8yRaom/KbwUxOcfrLolSvPifSy1nsgKtJEgzjOk1S8t
yxokANn9Xbnz2JcFNDausEO4l4os3oSupEKWI1x6zl88G2mh8KMFseFhBMuzojPE8qjMYfHskHXB
fblsbr/j8bqDS+AZLrTXVOhGyu3pJl++WNpUK75nWMS+uWE41NkvPt4+4ZLzY7sK+k74ENOtevUr
TyxJrGtYif7BXmsznYS7HeYEtv3fFLav4chZMFtRfKnY9pdWMECtrkDaDsjPtlss7Rk/NtwRWTL3
/V7iq26JQxqEpYV8dMjeC8yOrFbi6ihfWBPC+C+PotLrlKc1yw1H1CXhDK/INoJQ+Da0D7etwZg1
hGDIdK2PBX9wpF8vjLlb90npUnS5zU2G33YRyOBeUHVU1FXZRq29afDnjuvFE8Kv/Vhwn6ejAi++
TxiJS5upoucBmwcuh4E7GDvdfqLdQzqJ4Qe/MfdKOzBg3AcNYl5Brj1b9nSUNQQ2bC7t0JGegar1
5U9aRXKpZgEt5ia9oeKGlxKjEewfZP0yMfaFd2qyToNMvz56oZFFC75HkDVewaWKS3yCNM8/mSmn
uOI9y00PkSfM8FZVYYrmDWpSRlU1sIAR6Mahs8SF4xdqTbcOzVMvdm2uY4U9DPLyHsBaXEET65TW
8wuqUoy0rdGxNGKpyLtXl6sTC5riy+BEEaHV6RkSUhuuE9OxHcqToNxGtyLEFNFs9U/+Jrtg4uPx
5eRZUem1AedVhqU6YYbSpv8dc6syRvr2DOGTEw1VXZ8iNolQcmCLdfbG/S0F5ZdKMTan/wej3d77
dwwS96UADrvFbuqgPTBYGXLlriC/Dp/sXdTo7UzMddlZCn2jguzc0GvxwAzLF63nJyo565bb/t10
9kLspu6gh/fcqVxKyvEBJDaKtEHbH3xGMEn0AUTPcvpL9Ygd6C/4wMRYQLsjAolr37kt3AdqFfnj
f0zSF/VV7lpDbJQqmM0Wgz369z07BOFv3UMn7OHa+rdBwtT41DQmDD5InsuPG2S404fo4ilcTX8y
wyffMnC/QYiHxV6m+l/Hyw1HNzPfNHOVmMPTFdghpX27OGAm52G20N83cU8uYr5sZnibKZFoDKyz
Y88iB19sS6uuak0U5eKEUa9tmTlKz9zJa8XhAgjOrzS53TQJjAdpKgLqCRDjmGMHun2MsZL/R85a
cQxY65tu/+SSxHQISUZ9U7GS4IyQeNeXRPiWD5Yo4XddYByQ++1XsyLIYSRaxY4aHMRaZbLRGF56
Oy61/woy4KUmxbALY3aGgNgtNC/rqI1zfhKhxP9kVyuH9mugBhxO7PYcK1TgPlc0x/MwCW3ZYIh4
l9t4Bss9PgSvxBwHsVlLkCfhRJCBSI9v5xUzMff/nsrXFV74nIkqdlv6hE9wlg+YzHOObe0zTS34
GQVSv/ROIKHo059OVAmyK7uE7wSSzf08vVLsYm0s6L6/LleRQQLkPi9j+7MF8ZraQCpdPxOLwa/t
lyHjYq1t4FZ5vzdr4u1hgxWAn5HMh2c2rAoI20mha4A1QHijFL7W8Kuq0257Vk7W/KEC71l4wa0x
s/R3rKnYQD6iD3/i3srHoRGHRRykZ/5ybrrdXefJm1AhLtYOcp2oR0sNALZHksRQzlrd4m41H2sV
jSnZBJZ0kq0L35PkeFkqJYhMzoe0vuyY3Q/bJkzUE4YRb/F5dENm9wClrDt67C7Zc7SwM7Qm4TjW
DyUJu+DSEDpfHH+FZcIFgWHE+k4H6G7r6tRLIorG2xgi4hWsE33FZ6RL+t93XwP+oGv48XYIHN/k
fAIDIMcc0LnRM4xpOoY/5HFpVkfmT589Tyer5P4czIvImSXN7otJlkvEznylgIBJMKli9kJ44mPo
/n1NcSrpBIWeOFwuHOEzShUx36QkEfqtfq114ytzzfdmgjG6jTf1ld7WIKg8ay7CF90T+OpB+76B
wedIfadeVcTS8fKRoSJ9DVj8QA9HFcnESo1TC6SNQRwbwXdg/4Dux90eYwZ0GZRVJA0X8Sy5MPOt
U1yrVWX7mwbMbUJTUYX/+KwXX8AlibPcbpaZ+9gQCR8nkZYMCCOGS+biIkVQeUrFs9n6egqyusQR
N9YU8iAy/g4puS7UO1SdUbomPoSUq4L6ajYkqm7q/2eGhy/V5hOhpjj8w9+E461bgyEgwQtvACT+
9IXNgpwf9GI5kjk6CV1xm3hwG1p2E2L5/zcdex8IgiNMC2bd80aVogQt6P2lXjsE5XR8qjDnzvC3
6KcIITZHA3uZCFFRJO+snc7Hmgjsn7Po2QQ0Adsdn/7ChiHZoqALD8Bk8mu8mEiFLjUh38ZTk4lo
T6r3zrPBX/m8r2cuf7lNC7X+rqk+wdi/89BjghkaUZhrx0W2OubC3V5XC9u5id4XsCkWYk15DdFc
XmYsvytKtt6R1eR4N3eHhpSDnmvMYxEsHUK/mJA5izPxueE825KE/Y9YmvDX6zAqPRDewPtlIelJ
GlmbLYORrVsW1Z3wMudlXSB9fiSNwvwHfV4yhxwtHCXeRBVtEAOKpdsBHIHyh6MqNUFWPJC6UbL2
lWi3XA2P3yqEOByjk6mquHbni8G082XSqBNzlE1zW1YZYZQ7b/uQ1koCLAUjs7HFBiUsgmdobyK9
jUJutDAEgL/ET152gIoG/kztHU0Aav5nnrgATLksfIW99VVVgZgIY1vBV3YSYFXqRx9UC9XWGk+u
xLQTrrD0QG9PFpBY3+p9wjNDxW/a/b3nLbKI5pe7ewX7uiVvXd5I01ba2M5gmMmFS79CsSn2XWKc
C62ju3QxQKkIvR1LrDNFYNTjaZ0YLvdkiGv8RZbnYNQv0TXCpPI98Lb52uhHRbLzjKuV+0YKJkbL
j9R1PNNIXAZrn7g5iVAD6+bSA7+cjHFZfQNJYbfU6iDD4NS3ZlQ1pzIjip/cxrn80fTbCY0BOJhu
fy7N0E4kzOO7bgVAz1NGRAImsr48Uq859xJPEcPpTM3hBlZydyI2l3LGyxReFkaBYLyQ1Z7CEk5U
F5mNAhxz0IW/jxOr+X9QteZ1cVDp8XFLKIpSeRdo89gIW5H/b5CszZO/ajST/xnWOGxFbuk/gP13
P5Z0LeCoa1QnUiCIbXBUWs/MOZmPey3ucFcLqVDUUdlfgnzvtuTJhV3LwNvOn5hqkcEIUdNAY31S
g+3Lf5I3bQPosCMJv0I0769sCaXJDWbCe0srgwZKk6fuX7c7JfR6modbkbmzWh3iPVTtVfQtD+s4
COc/LMStuAW0jT/wp9euawHADWukqy3TcFcieKt3Bp8wnZD+wTMs8W4uRr5UNWuwvhBRruxhuERy
MtqrjRx7p7uCHAhBrQ2h/Muxn6OUTsbwytl8VSwtRqT0p25poJsVjDEJ/nEs8mL9LXtfJ4fxGhb4
9gNpHOqb9kBu+KYJY36vE978B4Ue+GXDZzJbPr+mapheEV1L5cOtuLLk+bNz4ddNGxwksNKDRdWC
QD39CztSGYzfvNP4XU4Js4NhuKJtSm2h1VO58qMF0YUTBLjYIYodPwrU5PQ7qFCmG32Awe+oTs8f
/U0E4bBoO5Zqyk0mp5YsMSxsQeKUwSHcEl4Dgf39GoZc0ZdJRvhOSvCyDbV9ICirNpkuGEuTzYOn
QeVZ0BPMbfP2/tv1ptu7YgDT4KHt3K5qV5sVTGPH4+nGqi+S2qrIXjWIsDHW+h+m4coFud+nDHs5
ff5Cb7vWpU/Lj+JiYPJau3VKzywy3StlPPopEJF+FJn5qB1p//iWsBKFlXTF5whgPPnrftf8582U
nct0rHEUzsOOlJtFw1jyVCR1X1BHKA7yG740Dr3P2U+uYttNJIaGen5Qzqiv6APzTi21qtKO8DwY
HKOGWafHu0qhp2W++5SeZ8XNIE9eH1zXTdH83GbHFrdPGTg8Y6Y3A3+K1Y5FvF8yG37i9qxJvBDq
8ZzOWb1AeHdVru2TZloa2UPyL85qa0ZeqNUGjBCFZLJcvIyWLhitdPsYzK0lwJqTSdq4oXKWwj5M
I86vWqa248BO6MdiXBcKYC7JocKpSZwDdItOWl0yFKxis+CDdcZYI1Xa8KraN3fqC/BomTBphWpA
KPImYx/fBs+ABRP5lTkSUVLvB/Xkyoyk1VH/63M+2KomXjzOan2JVCSHx+dgA2tKT20i6IsTycaO
wg5dzRqe4CXbTryI/J75ivFe5ACv1NFKPdJgxf3u5kOfkcK0FvAhGBTdXA724cxzkOWQ9FuGCYUZ
+a7iStmmqNqMIyCzTGfTr9Jwkcj69OYDOFUDA91lxdE5zLWf8aDwt2a8C9cy4oBq8s0patUwXiCD
7BS7AXhtgKOiFokiqvpC7UevBUqGdBaItVgDG5/CCWz0htHAgjJsxcEF1LmsqjGc+QW1s8F64Pnr
iqvdWA/Q8He9GHVruP6jzFfPk8iEChP+oQ7rSYiFENuxreNcBd6vbFtG34VpkGXJ96A/TERQiwFq
j5WSQSN1ZP4Y7+teGgKlZ0Vsw7d4INJol7Kk2euYQsJMkolkY7fP+hndewyUv784IzrbvwX+y9L/
tWKY6C2vIa0kJtfxYK2UFzL6GiPgglUJNqH0v3KRSkd5dKZtQVVLyEXenz0BSwA45wNkfRIY35cX
0kwYvhJ0u6PNEssbiPc3CxhUN3wfGfeiAuW7f6qWpY/Qo+LFXDOxrer3KqR8AeE9PVg6BwJIFngL
UG3A+ekbfnQRsl0e5IYKyY32ytMoPyijs2bg8ULb2mutMk3fItG0KY89rr9eqQOhZDX3Z14gorav
4EE/9fMVcsLtrJno/7SUgV+G0IW7DK/huvUnvVWgbwnvFVU4K6qgM4FKmSxlT3At3n8xv0Gbkrd/
TUtK9e0uQJ6WmMZuXeNy/o3WxsXYvvVEASjTVmNlyc7FbdBsCvfuDy4ilvKp/KzAyHtRrSdmU/ES
pKn/J1tCSr+wU1jm1S1rBWKWEO9fNotzDiqpkU5EX0EDrxAWlh8dqezIunZDZmxK+L6h6IiGGzbf
TsytLUsWNNEw7ztckq2Ggh+CeJfa0zhCfuOTaDw6jcQ9qBC4k1AI5pFE1imZk1U43FllxV4YhEaF
4DYjLNvUkEhgA3dMX08Flo8DqaxtmMvxAWRj2bYH5D75HoLfujcxjrjy0kDWFD9qh7MbF6Aw/9SY
0hzMhZVPRWzBSFCySGZH8K21n8enWzMf88/1vW2cHoe2lRdLzEA/BtL9Sn5IHYZUPLH39VqhSyUE
C2gUDgSYa9/6hRNuFvbIA4XRci6Vbah+m9SfHt9MQyOkw4tEtKp/wYhsqHOW8UnBTUJG1hWDX4DU
O04S8EDQ7ih6NXDY+G9aiSuNVO1E84b3ooB75mp7Wq33lBsQf+TBxGVeah0bZnW/JLIRuvhqMvP7
Y8dyVYVm5AuJ3PzLBeToxLPmEiAX9S9bmkJJf++1dmDl9E6LflnJFD3kU1BAYEKWIx6ff7i+NPOz
t5ITza1DW0Syhu4BwaU9gguwcZ1QiO8EvS58IE29Lws2jmhQDDRgD1PcAGsll6T/5W+Ey0VwzrDS
8CizZ/hCaJ6zBUltNTPGFE1Wgkt36sPGtZkLAmgnN438vs/P+5Pi3WyGaWSfyiGnmnMPq0+sLhAl
ro+uXelxpa8WQjnUVRtW8tKapVqsiPfw8WOkQgU2Jb4VszVQaAPo8GFkvXl9WxT75el7PJwlB684
V33BEYuFU7DcTvAvdKe+QBiOeYQo7vSGQzZtuCJuCSHdgcWSy7HZuDMbDo4lb4efEbX0n8ZAeEZi
yG7BqJ/e6OpmS6yUjeJYZiCrFcnavJpuKR9S7Myx7NHgRJC0cQwhhi7F2hRu95c6VzU4KU0mMaPM
g8zi/+WxoSOar+ibbQKDRU5D2eN2vgwkUYTywAp2zgwv1Y1LFnMm3ToWrE8TNFycr6XAQlYGr7GU
MOgPa8t9XHAeOux/deqhk7oonxzTDUxDOwSAIK7K/9Atdy8fM8R/UIR3ir9HyRlYkF4CrKJ+xQwQ
4+WLKDvEcxONLQwjyykDNsiLvon31tokNq+sBw5Mou1U490tyGsT7CCikmYDxxN9fO6cE50nzTEl
4A1wX40giZ6isqWXxAU0fB6w3iwK8md1qkzqjEulRwdoe70kFNoOALkHvyh87TsacdWVgX/5sbr/
EjgF82bYD010AtytfHJueXC/mWRH/NLCuKicwyzETJep1KNXjD4MeCWXb5HM8xsvA+6wfkK5y9ja
xPPW2ird1vbTuOjRaEveAXVkyDU+bvWQO04R6L7SnSM8dM7dLBRNenTtm7/+Kptz9nrZXMYqu29q
ZFBryI9cjq4YwZcSr8xJFgdCcT0JPRRquNY+P+ucKOCFZJjKAfSbYPFBERnHxdivvjIfMyLszFOD
VEFjYh9nxiHrGi6hCExkEGbR4A5+EgDW5jGbFUWidxJ3xNFQk0dOsNn2hUBJOc8u5GdkkjpP6g7w
XyWCu+szhUzwqwCGgnsalr+8Y+aYm7K9IqWM3fcyAmTQZeoWsHPPygqG0StOBBsRtGNJFgDZLMja
ulLX3JxofFHv6qaOI41nCMcKkvlL3L/BjCjWX4pqjkeUnTbXsba8f3hztV90B/a0D94DfsI/59/I
SbOYmjA1WPdZtclNjGToawzCF2ffSWXmWFkbgImt9sC/7tGyO878ycuu8g7Cv6mA5AcKHIDWiaTh
NmzlvQhPYbxsAzAxfxa/GSAe+qsZfpNwj9Asu7mX8L4EComGOc98kuqAUABazVJdUTwT/rLL1+Q8
4WcAcY5/kiYxgWxhlXtRDlJYGWfQNOLsOLzm5v5VKYZOK5da9+RCjmH1LfaRop/XGa5N5UJdSB2I
qlMHaW05kHpXVsVqcVvK+feGp1/W3tRSA2eB0XviId9p/kS075yBxs9Hi+sPPl90FXszV16fFio3
SNniqaPAQPsto7P0Njz0jEQLGn4uwE8nWEOeTtN7FEtvTbrcghKhiIlnlodrRtQc48WEUglTwldT
kFKVp6hZ/cl24pEsGruGdkYWsSYIRBrKPEyhgS8p9gixk7nBQS0lJc47YIn6VbNrjGAvdMHcd2hb
rvLEX9DHg+O8hxHgR95IkzJVwcIVhgd0XGpXL/vBAmZ4pRGJlO6cImiTLZPHuBSaYPnUvhJHkjTg
L4OgqEs4a8+1ik4LpF/CPFdlC64G4ZsHJJjGxFoH+xcWSFf3c9puhp3cDoy83pVpRUOflrn+p4W7
6jind3tyHttocx4xHV4NWLCYdod5VtwDY8TyS3m1wYWSZVlexhMk3uTUDY50w0IkDrn3mhkhKKdA
XdxlwlCRaOJ1Wk6o1JUGSGMxnF+DdsNyQHDhoLqEr6t0i+5dkheUoWulPZwgyvcw9biwP72kEmUq
zF8uZuQ2zjpofmeoEfwvMaSKIOhf7wCCUfD9uQPqJO8lpOejIVuWZGuFL7TinwjwEyI1OllEpsoi
W9Jr2QTfmJU9eJ2XXHEtTTUsPbsY3csc8VFsP8xepOuB1pSeO5aFpoxDglK1swNK0mBSjNjwRaGB
PZFj3iPa+NwFQT6OrF1Ejxf/ajB3ZUar78CChzDxEtLTb7bTjDIfkzuV2DDbDXvE7BJDkaLSu8jV
gLFbttEJAFuKBYbgj+vsx3fCtXeAqSOXOypXDG4KKl/M4r9hsWe+KeCaSZwDIKWjvJ4QRB12Y+5x
SAoYQYdcjUq8Ib/3zJ9/flIzKf2aLfhoSmHxVM1vS1wdPacrpsFLYEU2ODNL/yNaSxnrrZouemUb
lsoR3YdKca82ixsAVshJar6P6+WR9SFtz4rozZ0ilXh3wwBXwARMcbxxBXZ25OTtSVJegcttqvqv
AnA0yCVCPyYbrNGGpRMDjmod3eMWeUXOpmWWitPiE/8gIwS63SBUYP7jzgtQgC8UfA2BfcYEaIGn
2XhWFIXUambzZYbRZXHJtWgMTrA5JPuH6HgJLXIfowycJGXzDgNXHaTxSU3AnjjKxV3bqit6V816
mHXaNRHvck06HqASp1k+kU6m/UTT3TdwI2O3jjyYOQD34/j4crj0iRAEkw+Lk4xXO9X89wkQBnUY
1ZmwwKwcJ9hhWXSl4SPzQ81cLEzJmJmCW2eTtwV4Udzs1SmMN/jNZLdoP/eIVRgBGa/0HRTMuxN2
mvcX6bPvYMagqBythv9LuQb2u9VwlPOOp5r3x6OqylnxckkYpTVephQjEaTBGJk/e3Zo0p7EWblL
wTsQUbaIga66UAz63fP6DLzcSD89sam2sDkx6Ob/zn92/EGwfJaeeZkzcszVonmWEnBtN+RLaVSB
i9LuuIpwtzjkTVyWkwDjpukHgvvyTSbtvGdwlLEX4dtMmYQPR9OO4JppKKe1RkUOHuBbROM4aRUZ
2M4A4STwTywQpmmpFBKNNLmv6fikN+XvlwalSEde4WXtqU1SQ3F+X/91SyOrXMIDm04pSDz5UJXC
+7hkIrCtcUW3yqSLgF0EwmLDJa55glYeln+0zLnjs3+pj6nqqgeQJHyYwV2bmj3F0lTYQiF/IsjQ
NU6cXWYbiKFe/HAuntZI7MyMFKwtHLphymxzw9WWa4wCbHewV5nXBRfvihGtVMuJLA51wMA1XtDd
la9Q7mHmKbiFXrLi95WDCvcuRLIJNEhyrmSBkH6aGP2mkwD8tyK+CPVTB/Wm9/6X9ejlonKrY9ge
jDnkMg/5qksTl9+oZcoRxihUtZxJiYUVFrWOTTRsscMvEIFxSWBxJIaMB2mOyBJOnGtowKfj6SHy
yLd8njzB2+tj4i3hT72efkw1sfgsub8dEsl2/FHYD6rDOsogDrg/eJmyQ4D1hLQU7DNGZLmAWPiW
rHeQthcaRTwHhnGCT/ukKFhlHGizljAYx66TpiDmTftXc4TX11qvg9Ud0qEdzqki4rcT00HKNIcW
FdkAKvyXwS2avDrDvzj4VnBZI8C9Y467epgcjucPyWOLQT88CVsHWzogiNPI9x/U0c21RVvnRU4W
RwsGzMOFfm39AiKZLbuNHGou2zvKxIja5NPKmWbuNr/oOhId4e2djDyDl4Y/S885ih1PD1SzTj7k
+7+P3IsLG6CKPqMPRSB2FMABT3GV0qXP6xK1CNbAV4+9o/0d7z5XcVkmm3aPqLxvOmrOt2cf9N7e
RiAB8KkWlVJcdms9LdoLM6hdR339yH0t79rd6RiZTuPIeZYZKpOkTE4qitLKbuvBKkrv4E6FipoF
HgHX7rqHwpjr+upnxQCOZP2TPF59/THXGU8eBsAJnwjBt3vOQOpdQHMuRXNRnUIs2QJOPwntz6/f
7P01mDamycg4aPxvr9SeTb032f+FEs+EWuFf/9/LUf/h4r2SPafJ8biwOqxwSv+zbB6nUmRvOxtC
ZiZIvwIJ4ZYFGhdZ8ILr2DZEpWbw7RZ0pm/Y1ryup99DuXnSNhMf4oLx/v/G6bm78qShnmcLHBHn
jGT6jkZ8qbYglAX8wBRtbagNqT27hhqG+yQC+sua64Z/sCGoy5V3Rp94LzjjypBFIPZA1hmku8wO
di737ZQ0aivZaaHxLlP+COfH6YyD06E/HwQ0Zs4DQ+BaCycPXtjQRoAKaGcp9qhYpJANPFf7d0gl
BMr6OlIiOn3N2JG2hjSKm88aYTVylts+ofbv67nUDoHduUyER/lHRhUlZtlOhHjAD/CbEAYnsWBj
MVwjqt8rqovsBBeypdhuKjf2Y2GFpFFOXzmInJa7hTiuaEyjOFaoG25iML5v1CcApcE9hr5Notaj
Bol1eWAtVJ8t7oCM10Y/H8FkqA+11nNNf7634KBMLqqSpWOgxQTrFJ5MFw4tFH/89A9ielMcUAo1
pLiYq8yAsmjNo8wGIiJRcqGwU1QGMTIswTJpcVRBc1pOWawUiw814N+W/y9W+YhKsR+c8WflYoo8
8qKD0KAir7CGVktYHRF0LWEsD9DOvim6A0qu4HhUQdZpC8COp7sTbKZdz9PzUK0hBnmiYKfNsYVF
mpzImmsd8ruLK/QAq/B5+desGUW7eIDrrdxoXsEGChaEuheVVsuqMpIcHfweSKh3VwgiGyc5mAzt
qEUTy4Fp/sDrX4NVG3ttbqbA9jnRFvUXFcZYIm+Woo3mgmVbJ5Up12PT761jYcOLwCjRrBhqb9ME
hOQ/FiND2WIqpdtSv54YorGH/PU1WXhZoSd6ETaqioGYHYh/ew1jw7PjhAgIJTk6I31Rb215oUKA
3HYpu0dHgv9i0nwmP7C2nJWz3KSebawfdbkk/gj8fLS70lVXxXpJJAh6QBSp1fT/3UcoFrWQ0lgY
JD2YUPL5UxCjuWhbVz2mBU48DoBAjMYjQ0EC1J5WmR9bS/ZJdMlg+OKH1jgnfNNA+fxy/CtziZE6
7P7zChK8bSpyk28eGkFlrViVDRZ8ah+06sETf5YAjHbJZX16PvVT/QrtvZCDXxQGwNSpO5Fet8zQ
5GsGAN8TaQg3UfauQExOeJgcv7YGwaw1+qLgnJ7KUxf/7ypzhEvVUkDLyjL5cWRiuoLHlmLWsLxo
w8O3XCs54y5Pcc8S0aCUgeXSsHlLtNGd3Cho9jF0Vf2hlam8oeAyxR20+5pLDK5wkfHR5NbQ5IUe
jlIgk4xLxjhxUQnJEpsTWwxLBdgAkVld7FAEmZo7BaDXy+7QHH19vZE08F1oWXnixNdSE6ONSRIn
GMzWc9Thmpn6Ha4JWggpvGMlQ3jgtxZ4b5FSX4FwC3WTfNQkzchnKnFeKkmaq5TZFeVQh5mK99KC
kK8kquifpXjQeqeSAyCf60rnx3WGnGZw4z8M3QNWrBMkwJE2sw4Z9bKq40Ipuzi0s22SrMM5bNLZ
UfnnK9mQ2gcW8Qu1ZkWkV3U69ZTxjiMzq8TA2tAPRtvU9WAhzcqqzIdLqBfiU4TM2AMONS7LHJzP
8lTgiPmC/9Zg1J1sLjn5vv9+/+5P3JBFi6J9y7i8ygnupYl5diwHdnBs0OXOd0jwRglCyjIXHs0f
u6kV3KZINun4sXMUWJmcai4REot0P2AJcWCNRL0oYk79dQAHEKtTm1DhWi4tJ0kGQw4AreLWZ2rF
nTVsZU2aCt4jofmxO3nHuJwS0ZG54dh39PTOcKbFfd+DidWUmMbxfeXgc897ysm4xKMUFIDUtHqK
ydmSWs4ay9Wi7M7g4r9LiMN+p/KUeOHUzK9W17VEMYbJ7bIskCvf4qKnwB7jtrYFXeyBOOS1/zIS
bn4Vhod/9i7e8M3lmJD3AUykvcQUOgp1GgAYz+W+pPFdBc4xGWrgTS3eeEI8px5W5JYjijsdcofZ
VyjJ+FRtKYqQ9VFKQ/FNysWCtH7QM8d9vZykbs2mj/IvxEy/FzvpffWsaY81J2ulOH0mbKrs1HQO
Ilmjl8Dvx42xgV0ZwicNyLEm2WukSkHypJicSMaQFJqv2EAjXU+X2BdwFtYsKL01+uSoUoheWSEh
y2WXopicUBJ+LHqW267LTqKHwpnLK/zROIL/+KUGczLDzefWtA9UXTBJIMFFsXYLpcIq5XW0/mnW
g5AEsXPqvQe9MIdFh1kZut870ml2U0AO+MxjPUx8k9e/ZNbOI5AFgmdairB51TY4NXfgujUNVahg
CsQatckaAikcMHHXHLLgAP727JcDkPEk3rPYkw2fTYFMvOHYqGx1KVf0mUoqvBdzxHibgl0iq4yv
0sh8tyOy4AZ6nPVmYxidnMxY1ogRVZiqBObFZTFYeQJCJdIJnfRTvDORED/gxOJeji3D6vz/Qzuv
jYTLun4UNiqDd8KnSiQeQznH92ZDqfsh1tdJswzePr9+D7qaCi9Vl3VA6kka6+YfK0OEzsqJXCSN
Dxf4pJ/3KHNCEzYxtDWAEUdx7EjZNQWwR1Q4ai9eMM1iVNnZ+acUu9Pi4KHNltWV3ZmvhlrJLFYA
N1h+5m4o5oXK93qBeUkBfDbO3EINOvM0JmDlwSEIJ342D6lCKvh2Q6lJCv7d9ick30xD2xlqnOTy
SdJJe6xmMyqhbYiqAx5dJW+m+Q/+rVuwuKQKErRX8gRHQCmczYLYl8gkdiVHDrBqn0g0yrIYH4aZ
v6JjrJWOGlB9/8c+6atfyNcaddYgvBP3KcI0kKSdBwQHXRfMoR5kT6GpNcTP7qWP3aOevZ6IUubJ
K4185QqW1bE80dISNPM9qD//j5KVmlqQ3Zt5sf3fSJTFx7ZbVEAUtYurkQmWqxIaJP3wjOvordGv
QXTVsbu0bbY+zEWyncI45fGChZAzkMyY4wO4D6e5wxitfCfEBWqhafWIGKJH1twO+IN4ef46ufxe
krFa/m+eXWM8zojHVuw9dv8xT/9sShR2DyOrTxyFrH/1eTojk4e2AWFkBOf5C4xaZSLjlTl0k+xg
JinRPr4mwsbCUCjIERFqNCSE6FT3rJ6dJEzLO6z6kpj41ABG+eEyD435qW7ku2kt3SpSIaWQalbh
Si7gZs1iv6Nuih6pl6nkb0dFqwrDU7WmYJXQJKM1Y0kqFJhzVIjBmLXrjFlTiSTzNTsMrlK+ZTiU
kiPXFmavbHqLUKAf5klzxuWJaUEHVhrUMjqoErLVjoxRY9YyaqK+1aAd48cRxWQUfV8Apacfyzrx
MQMFzhY6kPN4JJyrVsEUXBNg6bMQrMeGRK83hePcSihieKvkYnettdicCz0U8S4DUsTWtSzRqQc4
O6MNVSUS5kNECtgmTCdTSbe5keGyXknEipmX7tk8STxiBdUf0FTpjyDylSQl3DVtGxKWGDahB1dS
MF82nYXXab9KGxZkhtJq0+EBVW3/xseVZVOcuX80KbKAB/7H1qPT1H+iCQkjDs+mihgok3DZeNQH
pXstjZAZlloKT8d1TDZ285TWt3VpqR8Jjnq2Z1hRYFQtyU6SQJRpKsi8DyUR9ZwQHfiyIf5orrJT
5nJMAac5/xJAAB8J0XIaKqQ8/V1Zlek1oHMzw9wz/FYqnrdq/wQ51QGTQtQBaGMtjVm/PeB1Q+5N
Z8rzAhWs+BDHm6DQx9v+I+ei/oHkB6z1rLCc/pTlVeAVNNrp1x5YdW+/t6yBQGHS9k/H3PuEXClK
TNQHsqq9ZLY5oqKcgVstzPi6QSk0ZQtFUL2B0q3GEduOhT8Odvx89leLQWlvfXe0gBfw42MGV7GQ
DmU6uoPJf/J/gcQwoXTOqwRHOW2tFg6CEzOr7G6D7dmxaELuL16OqEw5NWBNXEsfP/Uk+7SJjM0r
aJ4cmGHlLg05GOOfYrpN2LT/xRtkIe1/Ln+kGDkqfMqNL9iI5XRq+EPpRIAYbF+tiBxLfj/Rb2K/
Bc5v3Y5eXdR/PdVkY8Bcdw/4aeoamvBS7P8GjZuVMWcpmlq/ZLu0HAqQ+fTxVkmyipbRyWFtOhYo
6h2hd5DM7vfIhKAnKMpq+Q+XNG3bYgvi4AH0KTT+ZGxIobITQMZpI/agAraSM3b5Ozn412ij9Sti
qHEMcTsPfuxFZtQ8HHv1DuhtWOAMq+vklsJ8glluwuITFaBsv+IL4xrhKgevmzf2ZSwIr+9Gl5mo
0HxvJMPbWsNJmapsCSduz9y6lLfJ5EXRv38Qpk0c/hcd+s8xKwRuSmF/fBgVgtUjfmyLa3bv8TIO
XMwziyZl62c+rgkVRhpV8VZH3W4ymB6fqwEiwnqoS+UhCmBExZJO/pi9X1hFUbV3D6o4N0o9fpME
OcHlGOvTHtHDgb33Pg/vmx/+l5b7JJF23lMZwldlyuqWdLooa4rQb+XQ5dHPmNTRNTFpmioUI4lD
1P2PoY1YdH4In7GfI9fvl3zpD8NH16KIWWHBsON2kowKVpnawGZRzOjVIIjvJSL5rUXDicYxfvdx
U+bk+SyRQd0s3uklDferAi9NnVDslQuWqIsPyIMxTylX4/RLDNZFqNGAMKMHiA/zPUldmzB51C7v
0u+2LlyTHrLLOzWIgmYGVSskxApyR8IgyHP1ULGqkQX1/O4lb90BWaIdwWeOI2l9tUGVXxH7hUPi
9w5G2JJ7r9Yaug0TVHR5c30NUph8J8Iq4+RAzdUAsitQmUXacpNt3Y4PzVnwlis5HpkMhIB2yGBz
sf0VW3343VSjIJM+h8itMX4v0kGy3qr0ZZl+0ObnMSpGgzVGZNpujwtKIFeQxHWOr43xx8QshkUK
ECjVc8FhOwWadJfHfewnHKtHaL79+bMjEA+wVwJqP5OO1j1rMpZAbffkdVkDJGzbLW6qfuhcFZTy
OhewcByrhK/avGkDB+7x177VPkxzFviITuS8Rr8jigL+ULDDjGhkT/aCuAK/g0v55wDcFoaL4utH
mc5mDBTeW6v0PceLyw6hcW29jBP8rJ/44W9/j4HlFaUMwo4fvUW32F7wvtohTYaRK1yOyqmzec/J
44VNB7Q6KX/A9p6vfA4H9t6ujNrytIiXus2aLYRb5GJEiQMQ6FyDqCrBKW8Ql+KerrPtw6wmOJ4L
+SgGXrR1yj9j11UMsuUwk7ocZrzq3aV1fhA98Of6+rkhWzNrFbwq2LYExpNM+B5sDBXEQ1jGLvWS
PBEDwdrpzF+6oezRNWP43YQbCOMnea1amWDJZec93ISDsKIcPdCIXXnin8oiBuUznFNa/L2Tn43J
m+u6FRMhgRWCMIVVm41J6WJVzdoFVHZ+txGA/4dO6gkJO8Vpa+joUHojATD8KVC/MQLp09Dlo+jU
pLaQ5keRIYmKPyRsHnsznlC6V/WMvmDQII+NlKNgfrHoVHYKpGEeRvbksfDJBDRanL5FMqtmziby
4NcCjWLQ+Du/2uu67AIeCSRaVqwBRCujmbD7fTEuAco4w1dbf+fYSd0H4O/0WcVml+I2qKWUqKH5
44Us8oL5XfzybQ6IdouvfALfbZaSMDAcTezBez1RmhSXxdzQ2Lg/vnbh+dqEsKG5yTZo0KPCls9h
9vf9oTcvcfFFYnCf+uAgCYz6n5nOySK2LSh9iLU6dhvVhtpOrsLzyFrQU9vN18JOLgh0KqtAKLaQ
rP/Zg6QCiuwf/AY0dDqPPoSpArnpvB8sgfOdD1AZ17SSiaFDSZe4vTZVv8jMG5kKkvcXVQfSB+0g
ZTG4Chnu0Z63xlGT7GaFJv7ERG8bkEodGUFs/ue9nVhfcWe+WehgquVxxy9/9fXRylHfPFagIFNa
TVAWa37ObkbBumZyjLxpiOfSq7w5HEPREg9xzn1OInlcBYugJyfCiioWmPT/a+sADTO3EUvRd3bE
du2m52/icI/WttAu+6w/ah8ppLNHpW1Rh2g3XsbBWSlHLhmTy3Dy7QdK9aopxYkLq/1FnTdEv57G
usZiDdPq3zixf5C3rTMDC1qZDvbuR2XE7sO6ij9b90gZpGqsubL2IACixKIGs5sqvczbMe1Z3OQ6
ugFw7F+/t6gFssF6JR6TTBVoGIq1z657c8ynhvn9h2kJasmsAykT3HOqHd9QZwn6W3eHhLRdUB/s
sR7VYHVnjzdyfLHTbRwNpImDe37WfBWoK9J+xBuKcQCHkh96txekpDl+sPwmOSoQkR/0fQa8vKo1
OrO83tjyGBUimuaVpbzSpvOlEdmrxSUMPGm80sj+N8JFQjihGd1IZXWEMzZtAg+kd9fM81zw15VP
SVU/tVQ15TdrTEfnjjeUcdErKWGLQPLXLwXCsjzpILYS3mk06fCzZeFlJuQq+oLT7KNpF6a2UgQp
2hviAQ0pQBfEaPLQ5ofyh+g8RcA6bmuQ3MG4BQsfXdAf1o0b/4Eond2jqQbWVoBlk2IpFvsiMdlD
uXlBTR4x0LZRvSuHRo92igGo4SWYS0fw2FRuYVZlPLmgvOnUHFGsYjyFNKZywWRjdp9Rka+7ivq5
S8W26YnLfgjEV647XUfCI+qh9MjSGzTNcuaJ+zPlAd1SqRbhR+C6zmBaEdiAaUUQdwvvD3JPHZFV
ohZ6Na3b6QkQUBuewUx0IOI2gDwQXvQGdnRag0avM6rzx3xTrsAeohBmHzp0TjEK/QfMqYqrOqPD
9WXPo77fa7RMefBhrbS4LV44E0RGUFNj5XN97OR7fMvbSeCAaF0PXFiNmOoBAql2sFb4yC+yuqde
VgX7KnPvFtfUMqWLZQCGmR8/MyM0CD1GgK/yjuOeqmLwDSMA2RA3oq3UHuzFbt8/9PmFsCNF5dSM
4w0tMuT1j85PmczS+4KEZFuvcPNX/esQX6f1+bAVr8c07/3/Qiy+t3y7MRpKz3LzxijTjUxd6OqN
X1HbTpIViXmoS7BW/PjKXFgziZ6r3HMgPlPZK+ZRudxAWiMG1TydKkjav0v0sef0rrPSUv776miu
b0akF4Z67rK4EavcgbQSZ4KqLXu+uQErAKG9GWyFcJ7CGcfGDAMBzDhp7YR5+evngnptPRQ7uh/u
S4TDQ8ZGt2Xb7UrrSPGnXedSngMyKPI5BOFLt6wEjLuusVMeD29++QOtd7xTtMYUMghX8tEWcknx
La+PjnCDWzlVVjMvwU9YRJil2+8zn/qzffN9Qxu4SaLrwNbCLddHLHZ7yhLvBa0LIbFY4jgeueXK
1X/AqEGTeSus3Qw5yM/knCVnGX9Q6XYcw1HzbWa090LHi5d1r3FaCRYVnsbdlbqgnszBelezaItA
5NaxxKKC9ZIrCx5rPbotLQ9U3+kKGgsFFoRRjoi6za+2Nq2CHr3YpHAM9kWJwxEqHcgQYqXEpu8p
XzLzqyChs4tBdms95QBZAnV8keSNtQD+rxHOTnAhnpnHNmZHNd6oHo2Z1bkHs/djyfLf01FV8Hd/
pN+q5Rq6Xd0YEaGhxcAuJCxcdKbcx4isVsvGCpauURkILDSrcd7XTZWYfyGUtJUMNV+lbVjYLsqm
Dp8gZWKcAVFDiMfItQE+ElCVp0o+tePbbRoW4hTKVvumtEQ7kVGjuf46Qr9ntG4Sg3LPy2SdbERk
U6gKQ9Epu4iLeL1Zj71KKrF1LnP4y4vTuRtgvAG6GZDrEi8XRxohf9O3MgT/q28KbYCdYTBtkGJz
WXljX//Y12ggmtG2/Z0yp+8nh712HEDzDsTDBvO3ZRC8Ebq/6g1sxUhGNRlo2bs6qb26LmB9yeQX
O/bQ3GjnovBQJb5Lb8duBg/qdjZQlyeYX8jRLVDGhLpSklIzxkvuTeTS9D+UA1mIfb5Diq8oQeKp
dJDYS1sTXox5NrbSPb7rQ0GV5Xoxien5kG5bnvplmYg+bt+81ehurEx1kO5dA2YTVFEHOZW6Ec17
ORYta/tLlI2x3O0ANI/YwhLUreRaJRB6aPfUb1O7Wb+5gigmFSEy2IwMnR9b1cabEsfjmFVmR1fF
usY0jMQfGl96XoR+B5SMtbjmZalHYrlp3BUGniPLNfBIKmnSVXrcqf31vxW5rwyayWRAXqJqsBA/
VJCzSLIeIXfRulaGvoFKf9jCj/lT1W5rGxUw+do5PksR6Dm2dmAqJla3v41XEvf6if7clSOcyjNU
6rGrbEUC7c7e55QBqdNXJItGBR0NiqQZRwAjFbmrNiooBXlYRX+XF3TloXYUc8cp7p2di2CbIh35
4PcN0vgjRqJdzhKBgNQSZa7J4FPBIM2YZNDp5PNCKFjCvuVGKTLw0DD9kU4v4T8gxZcllwDGNfen
LC8uppEAg0DNj0PHEKr+wjhfPInTxpyTHQE7Ig0VLkq8sImNcxU8N+g23fDA0Q20LyQEOjMPZo7L
fPjhj9N37fMnJo2uPCMvB92mgGyiYEoF8uu/iCCv7JN373fknMBmE7irJOzUt41m0Fo9Sq67b6xs
+9EgReE1JFZ8SSJtYcEx59CXOeAxWxCo+euw/WjLm8c2OaEsa6H2+X2asyQL3LH4sM8xdzy+wv3I
62wEW9rlVzOEM26T0M7/8xwQXmXlN/O7nMEhPEPmg0LzjbyMSRTS6dNDuebPhpPYH5YhqPSLtMXV
AaPAkFm9GxSDie1QkkLSs3Ls7V3/otyK2YZCBrElAGLal1r6duzAH4SAbLKguWOJCjU6tyGgu7ge
qZYXUlfupfN4p6gbgZ5BhD/LlFjjvYx++y5iBTkxWGpdPP2lYECUOGa5zx6Mapx8GQfW7LgQgWtC
ms20FhukYn33hdnHLHUM58F9l/VGKZfHSvPEBOcURdL8IRijXWX8Kc3paNVBypx/Rdz7PBr4J3Om
hjVi0PaYZL7eSZh8G5l4vz4sk8KFGutmg2UHoDWxu+t0RZUSvTgCzTHxJ3UpiRjq22peVkytfeI1
P1w+iwiraoIOjEllBW9f5GMtjRQVnW/uk7OoKRRctzzBr3YbL3UBfH9uSuzKVdl2WkGugkERX4lX
vF00KB91PF4F+OpPC4GeY94zyOJqGvuMzanrfM9OyJCfrQMxp12WHiRpuEN+Hh9uR2Vp7SkKfYpS
f7F9HSiNlHEBlCmSLOl6+kyS5BPZwchUrfLGj+gN/JehGoTw2UOcs3oDz96W6E6QE5LIt5yDsPZH
OykFq//XS8C6XxnVwZn7bDXrFnBBvM5Fv5alQvi6OoriNSBDHFp/FPFzJ9kPVnFaKwSqxfMuqMga
myHPDw9HDMTnr/90ZsRZloXbZuZ8k5gPlgoZ7OyPsOPnUNJzxJIXnxfdFgP69kNTsdjOYDm/hrUw
wCk3aSU8AeVcIIAyK/AXhEycCAq04Vn0l3Hppk4MYrop+bVMSZVw8pItHkxmldclbL8Vw4PH9r76
CkMLs7tlFxuSgYHc/Vds91CZl6TtYL4Syih2v9asTaIU0WoEfZRDpw2c1sGJmXiTukdxU7IXW0Li
Jc5RFDsMjvxomie968bCYPF5ZoGO5cUFYNlp2XgEdyyMhLC1BnkC74i7P0w7B+QgXQAM+cMk0tKU
edxcfIADkGZS7B6ATUa5z4i9w9KzSPMgWSEGkNLb7y7dm612KW1bGphyUgGtm3SGYrfii5CByTlt
3HTXg4wuztRG/VPpX5NqxMv+HO21i5yhkSjCmgPn88k7kSXM3MPZuQCa09/Yxv6Iqeotyjgh8OjY
ozcRFP6R2oemrlaUlX7bjVxb81oUtA4qs42pTUP84TKhevy/EhUkuARCB7LmqagZ6bb3XTfDsxNX
5RT/qFAHrLqS+jk4vBDuJp0Jjlb4bS4KMMM6JSTzH2Bm9oW9TEhRPjf+KauNkj46SsB7+nJ7LM7z
1NFh3Bu4RGxsaV+VVXccg4kLeayfkVG90pUc0d8yweTS5hMYlZd1Y6Y/GD7U/1Xiy7AuJQhbBjv0
DceViu3850R4RKhurlaanT09hy7tp4fuucE6h+URcUFs2qo6rw+alI8vjYsVV6kSTno6CqEweOfS
cFfoO+YWUqJzFZljfNxuy2BKcgxaktFtsYBYCf0aib3Q/8JBa78jcqURWt0cPBDHpVVepwS4hCN5
Wp9UfA98uCm0kGzPzY556gTCRZFcpsy3JqA4Bq7Q8fmqeKvZakpe3TdIAALv4HPX/TcvnR1rioET
l03WMy5Y+yxXI1ev4FqJ91DQUIjnlxcsvBukTj+AyLi12azvw2VSigD6+YjKbRWLQZs5XREsetF4
xoA7TpqelAkTWq0zrrrmAAqmcTHWaBM89dfLDMBUYkwXhwozj8ucWzzooQeU0HX0zfVAk87aXU3M
4kQTA9pPT7Hnc86Q3+sH+whY4m4q9ny2xqa1RF/8vMkceCeENTqdbehD+sKc+WlfqOctQ7NnXCwN
DtUXcEw7si1aj16RvFYEMeN7GigslE9Ehc6lkHkGMKAHX2k1uOhn0abklA0bpsPAyv+4Nsxmd3O/
f/YHyBwA0fVmfnSNyS0bKxUQD6e1IaoahJsb3ZxZ7hjlHUP++X93v/NJMK6fVXiCTyptQI7feIOI
s+yD3dKu8BtXnICTV6n84Q6YI1Jdrnmq8m+oxQ0HZJYAVEcqIqys4k63ayH0XgV512FKKpKdmIBi
GNASmXk/bzSgJ7qTg+/3yuSVxSp/OWEzWIjZdHPyiZniaDOOpzJypeK1WshyedeJbbFX+/m9QTOx
zwPOo+b3M8O+LXxcP9FLcqkjnI68lHVkf9Z4BktkyAVd0WcoAyI8xePKvsCdqPDwLyen5zj2n+fD
8WZ6YByc2PwIgYVoCdv5soUOomr4NxTptdmd4fjgxdUWtul05NQZpRl4gYpEeh9ebqKBxnEXsYYP
B0BomI+0iZHiMa90bUW/S3B35/vjZlt/qFW7U9hNMuGWKPkeM8XNTmYVslYPPZY+ibJPqObaI1J/
YbmTMZOCZZyMy9jqRadaBakjcx3F0giYKsjsmOaIhfwhATWASxgv+Wrt6xyIKO/Jv47CJZtsyQ5m
ZwU55o6DUUOaLQcqfS10WMIFddQ6txVS/jJ565kbPMa65dtY8+1gW1wI3vajw0qRP0YBg3ZbzwWN
yX3OonMKHhkytrCEj2OsSQvHFXY3I4t9siAG3IM8AmuuMWlKcGxzKwFovmWTZYzWIP1GUnPfuomP
AclAbQGPlcSzZaWAh1fIK/VAXaez+bODi05sb7cjlIfityT63Lol9cpvVq2rbw6QB59RlxDHGe1F
TBQ2NOBKvACn7JfN0Ofw4ijixLqun8j7QEvHbyoc1k9skN7IBfRkMkM82sq0r14sRELxn3amxD3p
Ak0jhOWTMWxB8GjCAuYkg6sEiM4BjY4veyti/PPbMSD4+YtWWdGwsPJ57TUHh3eU++aUSqK30yvm
Ettv7hkK1HMgDxCA/UOtXG3wp1GUFgJ5TyGwDs44LBKEahb5LkjuWT97wVkqXym7G4UYXefF9/Ys
GunzvolGiloqIh8El43ZSQTuhwLJNdNxjt6VJBJZE/eWS5um67fhA11vrtPQ/kOirPBGX9cr78eA
OgcyDnDkDJRc/2didk40NsXSx2gKXkMX9arZ4DpYoA/s3WUFYMvoIbSPiV+394kL4F89xY0dSDRs
FTo++k0kWh+v6rMDhEESg8peDi311o8XfSsCstJglz4HuUWF0y5ISsgVNaomU1SCCS52MN/laI9a
1dmAgR0RBRaXNyn8RJz3eZVoshLlt8rfswXvALevUuuxpoR6TbnCIRcRHU8qYJC6KInNdJhZjNde
lc0GUhMzU1ia6I/iTZ4GARikKHnGnlTU0N9pKUm4x/c8ZFzoIuSPpSBk98VbygQfq8TeGKV/LrJU
yXRWK2oydggTVybxR8Z+gQst1gMqL09gOsV3c/eEo2lIJFYk1Hdci7OqRm4mnXLLIGpAvdnPKqNu
uIt6c1C+Cwl6K7q5eLTM8k+d+d/cCSAZ5k0BNb1+D+9kx2gtJ2seFXiB3BCHPH43blPnlv0XbtXN
hppdRV2W09ILHhOF/Qhf0E4R3GvDqdBh0O1qhHyQRHhB0Y9RY7Y3wa+iimhE/VwvvjQyFGYVv8Qv
JDF8mxi3K/cQUT/MkrATC9oHWw+5ytTpxXzl7fMrOksP+uAojCrMHkbFXU6+od25WnwoeugF/dMw
f54dVGPHL5/6zOYhHsbZic9uj+ZrKcy3JsYszKJAJg+doutq0p+wk3v0RkcKuWsujcsU5cb1DzYK
1c4Mm53pqUnuvD0LyD3M1DCu0+nQDtANP03SHF72qH0tblD5M+58jD49IWbmxlxO47LqM1zRFkm+
VxpHD9ZchWdcms0eSp/hbjSGnuxYEcNKIjp2/pUuiiMIVhi2kpbvsgToXk4LKpA9FL7tnRKrGI59
W8uxjiZ/usUYqdhWyysJ8lT7w7Yqo+pjPp4WAVWuxNS94f2qyKyV8xxLQMsKPU3PwMkyvo2VsBoa
xMnK0c5zBPBDazcRRuJteOY0w4N6nlgHR7UZd42VmyqLZEbv6hdKJNJK30iCaC6scU3XVe7tf2f8
B4reahyN0iKpZUxoMC3ab5+lrB6zick2UDuHHNZRcKySMPxz8bfoIMBqRPYZxYCwfzpVZX2Drx3a
j0VfNwmJVAkB67sXNohKHdAectYIucirVld+8UAtXP9T6MJwbflEz8QuZJVkX8BCkTNE0U1ojy2o
/poN0MxhVyUAeJf+Yck5SEnvGazXtmseQC7gMakNnS8znn23hVvfOJpP9ESxX5xNRfdWPRKnrue+
6bB7p5iDL5+RzHAIZeHedqFXWATPLpAz/X4wpzj+WZeByntwO7WWbDjxrrWc/UoW8yc7UkKFOHvg
jzNzewxSK7EOUfZ0c3z/ntgjlmGiw0zUe1G4XGAow2T7Xz90qkafEv4hxllhYm/WYJCryd5OAzH+
ZXjAJQWCTbgNIjaVUCcPu5hubOK/IuVgwCnVpCvgaCcHKt35pvT3Bk87VSDTghn9O/gm4SMgAcah
j1llx66ijjEvw/l/zx/JRpg7lzUeXbS3gm+YUFW397TMHSEEjEyQQx2a5f/oO7J4N63qWxJIKeOn
qOlFPwy6hOStfWqr1mkFwlKYQDhVBgfvb23n1XV48J7Knw9/yiMahHmAboyiMhUnXiTB9LVm138R
ZZokBq73ep2PBhqUzk7wGzPKzKS0j/LcWaBZMCL0tx8WzpybNyt+VVYLkL7VT33y+pW7beVqaRZb
fTzibUwzI7U0N5bfm8/+gzEg60Ww+iqrZpK3X998SBY++ZQiXGZ1j7W7clq20pFp9/lRM93F0bGM
D7DIApLJbgbSEgVwdZVlS33nqUpQ/K4VwRpaYmdlv/8yuK+2u+1MWpflLPtpJxdG1xH+ad3hLgSm
grRBdAJZDZOfLEjoOyFyzCqeMbpHwItinQlIKm+GeNNJgW4PhejPaoxnj2jJTqeaV7YNVQRtLejS
94uATmHDvjfM6O2011oZWVtQQfUA/B4oKeWkV1rkz3ignQI0o9/ffCO2fErEIVyt0yISOjZKyyKn
kg+vwnhVtLAqt0GzXiwaeOjecuR76JIc72DhZZWYSsg49N99BVE8uT6Pnmmee46aCmWCCxC/ams3
r40RTk73t+pAB0SI/Kp/RThsZhY+3D9YLp4ShT3TXUYxTJ8ti6aMhJw1pAiRfi5quWMrEOGx+6WX
arq8lPjO4nPs4pCNdQMUnv9mmhST6I1BLo+L/2+j7aMRO22/p9tC6y8x0ZYSWUw7MEsPdnukSF4q
KlrawT8P8sAzpPPiWjCoRMgQPAf/yt3zGyUW0Hn6KpWY+DYwWK+x7fbTdQ2ALz/ph+smIIE8erW3
WUis0jttao0h8g7P8FCXQIucH+mOZC4y0BicdpjwU6ppZydZWEm+NiPuGKf+QOI4tjuqPJCMsg7W
52CUyIDPr0nSy3kXGdS1hRkgsn1niCUJaJaGoP05DXsRE0HggSMBlsUuf2gcjhkvGSBDKrtyCXfB
aq1w3gBuj4Qe8I8lu97YihxVbJiSCJNlRMzIc2Lz+1+yG004ps504vTF9i5anqgO8M7lC9gfMiII
09R2t6VhBmxygiwNuXJtd4hnY7FwUgToAehpNeHmyl2SgeYkFDuCh6pbecP7nDSTiCP6trcrx7ZI
G104BLXv9nQYk7Hm2RQjRF2g6UpVjOVy2CHYfzURsAYZ8sEmBZVds2Vy5kSVkveG9NvlUq04n2N5
sr8nyfdVusOP3cz8lAOgfwp4nNY3NUR9gKgAIOUCfONcWvCvbB9qESSgnvEOQDOmy1mcR9hhrEtg
T7Ey48A1X6I59ePHzljXH6TfsYbNzPcEGTZmK1QZG0u0/wOjP4Mp5mfVrgHnfIKj7EOZ+4PlH5DA
R8PYLQ6L4LcF8zrC5cWrntD9ABSAwEbHZdhCf0VUdcpDnesNSGTxwp0rGO/mO3lLblMT6c923Acu
uGW1kqzYtjIMcnkY3p+ZbTEO0+vSl8FHEVUShzZoP0Tc9O7aYBcWw0uVVQl7wkY5i/S7rQiHm53Z
6vtq/DuPQpF6xfPNeT3hVEiA/xxiQru24cYd4iftCuCgvNCNTxM1zjLz1ggXb8zX7/j5JPCXTk85
zveNu+rsFnBoATiH57QvJZJwfIz8wTiEscdH3cSn7VgJI9samCgW5gxWPtmUe2UkPHcRDuTNzljG
pJHqGlcpy6uZoLNzf/pxL/QiuBKvSscq1tLvuduth0Qss9c5uwBFUQJtBqh2xhI+mNBTALNM0U2W
bUEKJqOCcR5AdW1pAfDolVcnDDKp/CaqRmm4z4g9qqd6jClNybTcuSX6BidyGf5ocMRM5axoFWnb
NIATG0DVpFTLQU/tCVy5/iGUO1nBMR0c7TvcHxG7GxJRLX5AzGLQz/MgFcR9vAdXSl9MscnszLya
8iKx6guRS/KmGV5yxYxkUXskx5xvDPWX9Z47Re18zpjB2quksC4gLwx9cL7Rjkli7PHx+8Ji2Bxg
sfI1/Oy+VAg+fmvlJa170yqkL9mwGx1p4PFqoP2DuwUpxV6VsxxMSwEI1s9KT+Zu7/ASO+yiCTWg
n76N2haSDI7evS+M6X+H2GFyQFYLs0v5RQmx0h3aZhmRf2FL6o16zC2QfCtRP+GFezOTCnpUx2ma
E1xx9usajLn/3sIS5Y7u39k6L6YyFiQ9T4xFejEq1GEUDtPCEflaxotovbzXRY2U2ZEJyXKL6gCA
n0gj4dWOy9gY8QJuq98/V1APq8AhvanjiZLAU7T5dpotFrJMQPXXCLtyPqmG11VLEzQdOWcSn5gs
tWvBfDe26f/Ub+AM+1Na6LpMbD/6cBdI5+Ji6AucBnaTk1vo1bQbtJVnNJIKPLBnnRlsJ5Jg8Izf
4iJNOIY2OFTEEplHAW/DYZG4rbIc+HHBMBNgdeq73I2rc5SMkxw+uUrftA5ijLiky5yExQrYbee8
inHfTujwn/FfDKKaocX0LaLFjZ8eF4uHRudHjPrUF2lAqFyctbi4he6wxYbeXeILjMvNdLAbF0Kg
5QWHB6L1ZVW4NY3VjImXiLj+GIcsTTGM1Q66srL9qTxxXflsfYIEoB6RvUJdDEpR9ETAk2wBOi2w
c1CzlBzC0S7Gi4bgsXNThsLYNMv22ypb4YWWniQ+Ab6kG4BI0snaGIZV+X5Dm6NKUdXOmIm1V7PV
IDweNNUy/7G8LJP+5YaZ8SUvYIyLvHA4CishDeZDXcEp5AXX8f9JOorqm0tuwlyK+mkU/SQLhQ2m
/cjevzmht1t8D60daVmK1XxIQjiR4/o9wPsT74l8HAAAFhli78mNtY92mtZogDWNDNCnB7IoHEsw
BngrieABjD95lygAg4AGBjO80f3AMB/iQLTeH1s/DdfvmeS891wDQ8WPXW/6ZrvLpppsF7WRyj2H
mNVZx9LWm54MSGaHHlNVBw1DQ+8BjH4xlu1qUUCBdfEgp0zv0pqXkrl0QzkkhV+Yd+B1t9uxVXtt
snNB7hjdc4kofY2l+VeB1/QoPWzwd6ZgHCCoXCjjKk6DZWiOs4lSYqJsIirYeD3gzAjFOnNesBUP
zQ+cAiH7HXkkjNtBFayVlBh4Id9kkeqg63Lj2WVouel+6M3FotACWY2PIsh4Gyt2kvw9aE5rNzAC
DRf83q47m5wa0zAKdhsD+TmlAQb236pteJOp5rE+tyWBRE7zDOBSAg8A2mEJlMvWMt/sNQBX8pIP
m5+6X6tJPj09tvUTOVjGtNNP2gKlTfcwnPfGga9fC+EdH57aCj9PF8twndlB1q5CYmTu6JCo8Svy
J7he5sa8ES1P7BkXmcLqEFDX06cVwfYMZG884UWfVxr3BgXCQS48wSGSYrTkOGpcotQmMS/G9CnK
yaqPOLY33KOj78gATJ296FBv6xBFM/0oVvsilOK5XUwlaCZEVq/6GjBFiD5pni3Bu/CVX9YQLKb7
HsrvoyXnzfiM+MamD0QyiKzfoZ+jR5SLWMS1wFed0ujEvLp5U9VDkSE6zfP/BopxASPbV6BVz6ES
IRChrAVQJ0TqHo5CqKCGK6L/dv8eC9F7ELJwPSvenGSYlsdwXCFW2gL0EnEhdS58GayGT0nIRqin
cis+raydieBgbwHwQ+fQr6jXTnCW7G46zHWpnTwO/wa/AH0Ne8O3rzIvw0vIDVCjEiFez7ty/KNL
reQUOgKudv3jCPZro3rJB8qK++o1kYN1pKTIED7Xy3tD9jeHofj8qh5UYVsJPEdEkTQwR2S0dFlH
A4dqbUGk3PKObpUZ+LxZTB+6JHhvTteufm7a0c+BCOc2jVWyDW91+BvTesk1tXXRJ1HzokLf+DcF
ZGoEJXNLunaN0zYlFSQn2TCUwTYkiKd+xn21GDZRsOTsdqHLWuZpQg1VzfcdbBL9Zhvn3fOkMSw3
vA+HwD88QaXcDmJ5O2Ju/Tg7b3JrMYWW/wtWQFn+d4xzLfL7EWeq9oqkRhWgM8A3BWjxmSBSHXfH
bMLafN0NpUQGa/8vGk1bGCe2PplVHoqnCONGwo7rRk23Sodx38/HRi/AVlNywiKIy5g9vE4AwVgS
ItyX/J2axeQSTzBXi8agPsEb0YivRSTm2SYkfEW3XON7e2LUK0q4S69WzR6fOS3ylSuL5xetUlYM
a/lsRMrzaBZoukRxZoyWbi7D3JtDgYWupoAiL+25oyxzmCn5jgDhGDvhlQh/GSJ0l9ds4ohL+C50
4OANEtlG5Rt2a7OaBzEvmaOCSjKUVnvhtEezM7Z/kasiAJRl0o3FwsLup5wzBM+/DnmtcwweyL2w
t6UBE1tK3NpdUoPXTQpXcVN13hge+99R2JgBQP/VWSz7D9MBNbqWR/Wsh3dv8TnJzDZdn7Bk6vXN
OazWpO9VV9CM0ZL7b57+yU3gPxFUmKpaO5pF2RytUJ1xz7DoWCIfNMgMuLz/CJJHgL1KXE6/LkNF
Cdv9hNGgJmD3OPWGc6R51OJF1Ypd4s7ohLNIayxrmYJiFneQhebKUsEd0uCCfKI6rfgvrvDsvQ1Q
fScUI6VKZUDfrL4Rm6pg7hz2a9/WnoxaV25fEJgAuNe1ETUpGfd8h9FDJ7XVbnYtFSEU9JuWvgqI
Ke0WloKdrXxXyNoPp+AOJ3yeqAehF3zTg01pgPjdYtBREymLScGwT+uVdTgtAwHU7atxj4PydBYs
7PyPA7ko/2NxOWCbEVPucb59JbqTGQFdFDA9LF0bgVOB07fOZvCVvvwI9Cmrgc5l4Pesv8mu8XrE
K/uJLGAR6V1MyVZQRH1zKbAjIQ1Z+uJ0lWqUyy6c1IKZX32B/J+UleCwVj5Trqukx4F5WtM2dlSW
xQzr7O5H24lv0Q4okAUL8wiNstmkbL4P2QPFncgVWSvk8IECKwQn3j52hCd3Y15nMUfrDQzSV3O4
bzyOH4fMZfR3s2EzyH5RQJQb2fy9OEyST2GAOqMf7xKw75qMcPBd97MyjzD5A1ZOG5/EGJTiiDY6
+EROIkHpni8kfvdzCTVRSXRdt711hxQ5ZeyhBEk2JZX/s8ICD7MPS29xE2/6L1Fib1wHPU0Tfxzr
Sx7SMUPIWWp5Qsjl5C0oOE18mFiSCwwQW4RGmuHfCfqxtGfXCejK+w42W5fOk8fnwoVOH2bbCL1B
//Jbb01G7xDFxzBg9ILbj2UHpLKea6G093LFwsy5UqeeFEEpadbm1NnKw0yktAfB0+PcUGqiyW1L
alvzDHyiq3EC+ZjqwprqnYYhax4Bv6VcIcDjN9aV4K379brZAQP29up0XFB+mqd+E1UUfckzz9ob
IqBxImN6AN7hd37yX9OA01o0rZkrmFdeC9FYyRIDAk8nH2cytlCwMCA5XIF+2hjM+ZfBQWrJPmy2
jdbDmvq2uwBrOsNg8RTeJrIJBm3xARoE03Dq6iAPbHGbdPQAdp2AWPAlMWkpZcnkfXZpOvoWYiTi
n7974x9mu9vPNwumC8ZCzkvH83O0As9/zTG5222L+M8p4Y3UH5+tb9qHRsb9gWGkKnV2zQ9QetVn
+aN/eEczK27wvvHs7dkql+1QwG8DhNTOfMypgN2gB6/+8QLhmDSScmIWro7OG00S5/TqGctOhv4Z
LQ7Ay/ok8eGjadtwq+KfkcvA5ESw8DPW2MarVLit5UyFXcAIMi/U5wz8esajdocusU+ITiM9VjZA
q/MYH9mMKyaf1cP+R7rBNPPe5FNnro77s8U9m/kCvkTYxxiIiH7sgxt9DKO193gXYUKgOM1iU0Qg
GVxOLCo/YulO8xqivFFQV1dvZH8b8FCvqzoaD56RZ+2SXncz3aleX7xvH5TstaCH7jRHz6A2OdSj
2k2t1rbHEkcP6fTG4V2AXDEhevBikREZ6PTPvfvwdmAh/BLOFQpuPiZDtYYvTz1FbZdeC1kCT66R
PkDrhXPw3tY9MGkRvnzFg+lmX8dvv6WVkXhpzxHl1QxEWa1tg+SXDnWzM8PTq1HpA9wvPojQ1qIi
41JHts/EYa+kEjdvQOsz81CWOCmg19vkUr79ZE16+7Lgj6f01LUkRtwWqN49tAQ6MxBGBpEY69a7
mZba57z2aL6sgsnNYoWQFGawV5JNqnrG9TWeRWV5DXnAzHFR/UmSfjIxfe8nQUvcw+F5AMj8Lzs/
iv7HVWbO9AyeFkMMhs1Maj3QlFdPXyHeKPfub4H/fcVCWanqM0tjWqmidTEn7rHYp2V6V6zDF7je
EhcLJFo0/SO+AIF04A/L19zxYe1SKLnbqcFz2N0cqD83P8Es4xkkrDkbzCvqu1oHD0xzWn+sdGEc
hqDQqIxEimNXz1p0YUwsd81CkGYPZSpTa6tBo7b3YW7LC0nI1jnnLrOSnt4xb3nzVIMZUEfOXfRA
DgQcnX2wx3IfFIddlUhrkfL5Hj2NEEDZiXDuWaNBjQLpHIYNkAobhJwRK0MPrVGJ0raL6fX7JlmD
JkjgyNVIpkhBRPPmnZmIJK6i4yEdHoveIn3SRY1wNO9n8P9zUQmTcVToWCfpV/e5CrNN2ubRpGoC
rFdKeQOPm8SxNfbqTcry4HTQWXPaNA7eOuaSEQgNrM80OQh+2YUKynEwanlFG+zeVzkrU2hIYtIt
Ytbvd5n989Xai+62W9GuPwS9wt+Dllea0/pOv96nv1wDsi2dUo89GsP4aMR3TEUVqcv+rr6wBC7T
7EGPEy0mTr1gwEnWWhlstLupnh4i+YbdKL7xATyh0+qKJSzTwcN25nUcLz/MJ0S0siGI9MKEwu46
6LYGXKl7Ha9tDmR1Ui9GaEbS6r7Lt32eBvPT3WJHfDSKx1w6kSRHUdY0J/5cwAjjR4qfOuoVT54x
WsRAvLTlFzZq7z4CHQjdv9Y62aWClKA6/QqCCvFxr4TZbch8eFSi2wt53unken+TjNU/JC5t6+kP
P5C/UgO+F68Ad2bjYJk2648uc4PaDkK2IDW/YCm0sOa8hfm7391AefoBjNR7dEwKAXQ9PJDqgIjv
rR2vX4enTgaT7YERYkZm4fVImCs4+F/mMbY3HvxAL1QOq1VtRLb6r1rkgIPqC9BOmDGuUeV+80yt
BNrAthrrddSbFbgOBb2bthiepMZBOBPCSjTBC7hoQjQrCUINv6rOTE0PluRKz5t7WFKsCtHJuyB4
u0HiWPcQdb2CAWpdzvNBKwfnJI++oSRgfCT+3Oc4mWtaPnE5JvtRzlQvIe2SOae1wcmV3lbcyoXP
VoR0VjIrTs+w0se9AH3ABItmALrjl7wn7NGduAi2898jlyeTmWV0QSvKWFvsrmZVIfdPRBFwXYgh
QSWm3VNhsvYjsjFFTeTBLAYCjatVEst2NlXQ5/sucCu5Rd13zVTw8+hmG8VDDjrX7+pXLZa8XCHY
x1C1B+z+drPV0X0a2Pp8hK0LdDO7oEFoHSbRj5nCP3/Fcy47WXnDkDoBi36GjV2dudz06hqx/JW3
/04xs2b1fgGvfIFHf1STiaVpX1/PzsaIohhiLV/ytUpX6LifJVmYj51voYyGwOuTkJAUNILck3d2
6fEeM4grUXN5kG1aKO/Xc/kUzyJgL+THmhXc6L/SNS5Q6TQnG+jW/1+2oZUYWFg93RsFeBrRhsCd
yxDp57X3Rbasx9d2uhDFGDOmTiPFMYbjH/V8TeS5OtqW7P+cwUIv4tNm2slaD6f8AMzGXiiMeleT
BxZ7/Hhb2Xoon7hCJ0Q4lU8wcB+hq6UZaSuc6BP4kKfkUNG7+wFjo6AtalqoTx+1M0v4w1QUXqsD
Y/AQ+8OqqpOWvstw1+IsDzNcu6Y4X3PeeNz2MrQzMAPfQvN22A6dJ0JtPpWaYrzgYNPr21/S+pSZ
jHeHBHcil/qlq2yx2LVpzxDUAe6kCNBqHWNsPP34aDEpFF1ZLyo6Ti0RDC/t9XqxSdH6aFYdarpb
tLuqKo2/HF841QY3EN9uKc8kO42Ofiv35ektjc4TC9xQynOFLhELFmXTDO9ULpFrTW2rFbdubyzh
lskJzAs9KEFt1t9pQyvb49cWj2og90gfCjn2mep27caS5kPjN4laYYhGJA3VMoF6Y6JWATvYIKwZ
lFpxOTtHVD3o1sECHv0THac535qoSJKVML8omMvq+RqTCvzXj9lv/lBk1nO98ehCplSA2uLsJtlQ
8e6lYNSvv545J+OEzIp6j/CeJ2qYaEdTSzf8QmGUtf+vaiWD6tqY00TLxWj4DZUGqLpkCwSCmf4u
FxHlav3HbMPcg8WaUlV3kvz+gBus0m5N9yN50J8/JZ7AzwK95YwsFzjf84GNsBBzMnGxc/VuVxqL
4FJlHGQsRb+Yn7WtQaWGAoOYeaFiJleDP3Ys6UkMJ8uF+8saFth6U1ulJiRK3xdijWTzmzqax2o6
a2tYrXkzKxkKuZwwNCbqBsHb0a17Qowp/2er1RWBRQsZveZDBEzNgLVM+ZDzMPlE7ykQoGPlznc9
jlGMECGPF3QeSUepl57OKDkitwllhZ/X/XXHsJX6Vem4WOfgk5uxxBRdg6W5/XPTIcmLbeoo9NE8
IHNr47rvBKsaR4UXR+Z8kA8G0Sj2cyZ92O+bg6twwIr7VhuvZTxMOrp+N9VLeefNkgnybPDRDwJO
Vn0ApINilZIj/RoGxbaqLzxlIiSBLqVujkTC2/QWvQUY8LP01wazImRJi0LJDFJ3yLZvusYBeVVT
HZL8VdDaq1DrrBoBrjmpT12xSElrlNiY5JPYZajm/hsMiu+NfJf8xmv5jqT43ZzS6rHhC5KkECQp
NXz/JO3CaNpAJLWhA2jHhVgJ2/3CGuqEHLI0bCtD/velaIoGRPnJAamSRueHpKnyNQBC9Z8b/mmX
kGUCHeRifuzWpFWwmHRYl1s6Nbx6Hx7I4+sLJoq7xQf6mWBJs4F4jwvTaOP/OafwnECkGhk3piE4
jTA1azI/xtQcYt4cZ+DYxdNYuMFMqbdIklbFVc1eV3udeHait/rBfimSH5BRSttbzoLmt2xWXgDY
D3ThGZBUKj/FbupHMgBe7kbVmc972kh0MYq0gZ3+UXwzkE/S1aoxpB+psUPRRJc0xamLDgWwkW42
XNtNIjAc8f8281kzNvcp+9D264PAJ9o8INqAwWEgqI7+lBcSYZ2wc1/uUmQNJolnWodabOr7YDBp
KJFVYyYWfxAFR0arWY5PxIvd+deQtMQ4s54AgWopHuu6FsJuv0kSASgUMJsuDt4UU/NAAoXZ8hdk
98GBIlc1CDuJKKRYKCYaov+3qqmSOEZAJ8NzDw+7DzhBSzJhhJueWhX+6qhc3waWljRrwVyOvxvT
Y9IvoXqWbl9jzsbdRPK85xGM3kGObcYKCT46KcR/mG7JBu7moJiEHVBz3RwlYX8w2KYY3yo75dSf
gS5TtLriEjmChJohz3PQ+mzgrgAij4bWxpXM+na9tyQygMV7ihgj5mFDDQkWAmFvbZKEuUF47Vqm
wHeKNstXKUJ41wks/Hq1zB6k4yNpeDJtk0P1Im6A4TZ/AIc4L0t47oFMgSCyBFPlNRLN15VN/ISv
JZk75FQGusjg4t3l7JxAeRbn9gJ6VO/2+WbncW6OC/5Dt2WaAR2DAZi8E/EzPwflCOE0LwR9RAaN
8rEXM2JvNDfQ3geRvq6a+91D6f9xKY4po0062xme0XXVE6wwX9zrUcqzOaHaQUijQLs5WSY6X03F
1+zdc/+xaOWtUcJKjjeU4LN/az5TkypgQdKNf6Ju/R6wvelGX0OK2YcSlvHk+nFUAFJqGhyaILmV
GMWYrdS+HRGknYsmi9QgH3SZTA9TL2iic5o+MzZllZB8RutNNPSxBh3ecwz9jGqBEwk3kSWzGw1F
9FeHtY/5PqU1GigxzZljHkQ9AohWvD53LYgC/C0lR053CUrgsYb/KVVKWkcEvMWDFhkW3PeH/h//
XNgx6Wteg9dX9C/sb0bM4LRb7m6Km8I0qhMdmHnDm0JRfUQPujp0pDov38VcJj1fbBw27s0WnMXy
1ar10Rrnc0SCYnOHjDaLCWgegPQ7+CAEkgRIieVAwcXdv3HxLvVXahbqw4MDCO6LDToZWq8MTpi3
YmoQyupGauzJ4DiZ/yoJwxNLfT3OGdcKuT2CC0zIbpkF7SnyD6+RvGWW/tPVdT3D8kRveUjqvzUy
fWGRIJco+/OL5/FhsVdcLLOH56PAzH7aCdJfst9sY/iiuM+m2mNos0ZYszQfufq2KLj2mm41gKAx
Gj0oelM/kW3WwkXOi6iU5humA8kP3wtqNqbRMaN6IDcv+78Bx3x+3jvsu1LK57c0lhuXXoSE58KD
dCPwtMd8xflswKIT15lYDSgdoXlVCNhYOnds4JVgqM1Pz9kKwyly4OcBDNO8l12bSDvPYB6zaIF1
9eqOE5UF/8GpRU78A+bAFIZfiSm853Ik54eyFAo88K47U+6Cb+bkOgwGi+kdRNnwLZlxyouQNMes
DcFYGgMm+AlYQQOhfZU5s9r00+ksNALy3Uhe09QXTPxb20w5k85TX9hY2Z1eyvR0NYMYsXK0HZWU
ogWHEM0y8M9XUiwBsdsG5bNECIuZtdIizPuBFMY1polfsLvVaSXvjGIhtLc9Qn6hd8Q2TEU38Ieh
8YfIczKHwXBQ07HcpqyXU/lxFpnW3LPdE+TGasyAHRuTZ02xRX9JrjQmrt/xcsB66FYOmwRhiYZk
o4RkkZqCQQwA18pXqPnyUgOQpaBZYKaKgWYY0gDj0p95nOUNbXtris5rztYSpUKnlqyiQtSAjr2D
pOrqN7esYQ1h98kIyIPS9GRBOKhlirFxDJxz5DQiREo1Ol+cLpn7K4VNvvzr+nh6Qjz3IL/9LR5W
X4COE/u1fW/nJp0xMoVkrCcxzoJh3v0OxeJkME7rxzGW3Fd32GZnEm75zxLxbKk7I9QtQALTjI8t
q54+ylKKQKjPt+WpL4RTrafrKhuMwD+akklod6MLzzTbt7qZUkao+oH+K+1x9AL2EJyVh5upnUDt
vXLmOJqngLFKVKlsXpRWJm9sdv9H0dcCvegYXvNGSutiigMK8msHfAclQKo5B8z1X9GHxEtoXDh+
J0Ru1mg0d5S33j9Dzui2w2xpdqN4WSTKRByM72NVNBrMrEBY0QF6d9O1m0U/xFNrj2e5LNp75rFX
5yN5jgkagTXXq1/3h/0DvjEgK4O2g6LDoaTklqX85XmkbZeHLTlsMS6G3J81ppapip9k7AQxCYYr
dIsyXwo23/ZJ4OWkbCwR4MlYMIIIvyacI3VTb7so38nUbkegdRbgbpyA3YNzlicuBJrFs8QBGtFK
l2X7DwPeARq/IcuATWPlmM10qKi7zfArkNRi+yx+NnngtikZ9Nd6BJq6i4DXTg0FAEsN6UvZzekw
k7JHTY6+EDutrqen0QhNmcnl1BW/SSYtPtYgTspQv8D+AzRWkDh7izW/lDQBkR6f0pHzZWrUkDE1
bkNBJg2T14UyZUtPdZP2A8hnaSOktE4uHwDlgtxsiOTGQ8NOJ9jz9QbPNqxDm/5giu0xhQ+H2sBu
OMMHB77IcpebpYYNLg0sohN234tElpT6K5QRYSd3i6Dbdq7B4Hix86DOF5jeognd2jtc/bfZi/OK
DuqZRWlTAluABzK7Je1zVaFHQ0et0FA7BF+MwZcBloUw0SyuqP5VIElOIQZfHxFhKQmFc1weLC4l
ZdPeegjNT6kJADWgjeleALtCvrxr/PlA9qf1iNoJ4JF+mH0AjPmaMCBcllOGGq6wZr3d5H6JHoWZ
oK30a+oZxzNIXg8FJuL44k5LzIsA/0Y23R5jIgy0Pg0j1UGJKrQESh/mZZT13FFTkGACiA1g8xM9
jC/lXabKTDk1MnD6iBeoqJUaFKxIPc0W2HD378AcjbNnm79hAy4V8eoXXlwvQBV6IIY1AcatSz7h
CwTf1LK2FhPRQCHYsq5++tUcchdoreoOW8eKzKEzVCu6ZGU7UCvSHLC4M0Q540FKfvsfDMqqQTCD
lUR6tppzHaMnTFPVYOcg/u6LscfUCm5n8Pe4AC3kHTDGICSuwPO6M25RKDQLunfn3Zv4T8h/pUXY
f9hE4E1L9mT0rXEZQUKCVmgObPQL+ac+xA88vf1tmUQVFDrehXETyzejhAw5T1OIFfhG39aSAX5h
h3y61Fy7Yxhe+mn3BQNBUWE6tAqaQK7394OwQ23IR2BKRpL5kMwoCyhYLfeyt5aDCDTdFfsu5+kR
FB2kcNFwALJIzxXTQedS6CoV35rQKJw09+RhhWYBZdQHKkpr09MXiDrNM7FVF/uFYoeuYKNKMeYV
t4phacUFILGXjvrd8lzzp7PTa5TX23edTByaJ2VHEYtHNc2sa00QtLwVgIAkZm/nr1JyZlj9+rzV
unL0hUVdTQcmtFrSwRN7QEAR+XSUVv61sDdNoTTacCSG+w2gWPJyu6KhxZY+v2NH4xPfarU4hV1U
7KlygWhTTg8WOVyl/cdoqNrGhyVbqJaV1H+PEPUavEgmUmiD2ehRKu/Xj6rul3w6Sh7DJwAJYVmT
vayx5fQn4YcSOxqBYixjLF0PACmFvkUfFUkH2KC/5HHKAtQo7NDgUookPv/2AOiiJuZfC+58My8e
syfvBZKhJ89qLHc/O3bzZmyz9uusjtn1o49wKqAlUH/IG3ZTb7aPWVaM8fnWlj+pvqABQkSWEyMs
JB+gJuCZ+9V9h021xULvH+bWpt/9ZzXw4aLgBnxjKvvY3FjAybUMlkaUNQlkpLuHLSk/DgFulWlc
CUrwbETjsHlK46JFzHFpp5yEooM2SKxlEuDRdeM0l29Y6xcgEdO/SwOklRF3hpQ4eD5PNrxKY8SV
hivnrwX/R6P5O0yr2F+OZiGJAbd74xehcxLxuAjnLmOlKEUI7kIKHgVqpFbE8LxnhgDzb66vvShf
TrLDgfQd9hqe+uLdJOGGnXBvemv6O70wz6DQ0W0xuGu7yVPuHRb4hcV4LsH1q+7Az4MCtEfL7VrG
MoLFTHLs+dva3bHsD2J9WumQ5WyjBOazJ8mQfc/j0Aa3SGIrTfFvBtaryxBsBKtxNhl9PKJNwUo1
HT0a6KS6D9H9KHCU1gVJwlZJDu26cLGQU2dUiSp7QNrlvcyZwVk/v5Qo2E29tDW+9t17iPJ7RU91
Kj+WKiD6CIP8zzdWSPnvTb4zOSlvK6frZUq5YOrolK57noY8bOGZefvL/+E3bdrqr2LGKXz9rfkv
rzyvq21++3qONSxDoZjT2jnKuGjTFqmKAEVN4tB72rwksTIyghilK5HO/25cyshS2wb0J5NrM3rz
+WEu0LuuUjGA9rnDhop1c6v044KgzviC/Myr1YovJ6n4KeL2S50LURNrt6ld1rVZEq7X8h4rEITN
xzS1uX0Q7FKcuc3qpwXm2QVbELXiSogQfzHE16LVND0I+51xezoI/QjsgScoiyOuWExnYkmLj+xd
GrDGkmR6ksF+y2yls+K9Yz1IkpXP72ESVMnRfNBZeMjzq11vAypJB1xDlo3BK/E45XhOVLtnEqou
oa9++zU3s/nOeB8NcAZxWcUlbv7TJN0F37lNQtZf3AImo8FxQM3DmjD2CvSisoM7IXscbmWSDRk8
c8ANiXvrHfvLZHVMm/QOOpfw1wO6HFtNXUhOV/BFUdeoS2MzL7b5gqza1ufGl0Rhj0AarpvqUj75
s5xQpMlkkLorgjg8hHatpy+uxB2GmxLqQ9KapyPyYy/5Xl71Gv6lAKJ6tj58aRMONSwBKfhPQzsi
CYeLPZ79/R6w/nlYdQTZePAAKDCkcT6JN8FwrapfHTZm1fTFVj4Xv5Rdh44RE7qOyDeK9kxzhvkr
Nl4WoSc4E9BwXlx7BI0/kCzh8W84HEfVbp6+1FBgZX+s9j/l9DE1u7YUd+l6t3niVicPyirUGWzM
r5QuDjT+KDTD5RcAxyYS96c/fwfLSA5eENmRJ1PS7OE7v7wCjCgtM3SPQqHeF4gWCPUyHy1qPr4r
yAxHMapzMGUTTdLUcbXx6C4VJkVYslVtKC8SIigyOwDLQHEXZQ4b6ZWc1kjXHojdpr9z2x93C8UH
k7DQ49f4UhQp2cA1FrT7UkkA27xHcKRHJfVTVWg6pbjTAXUgFQrAU38YtpOcnQHTnjd1wmQDKllI
J28KNgYRziwlYMKFz6kY1ildfPPHSL2PwyfgxLWZhETAlLZW4Yoqp5Fyjajxyub9X8f0FXxBKWP3
Tq15c4NS7WbDEwSdrkkKZNX/vNqjZ9/rP+ty88x/yRWnOSSxlTTQRTykGO8zytxQ2ovED5+VSE6s
esAAZcnO7Jjex84BUF+zwNETSj6JBGqqtf2UehNuoxijQZaJ6aY9EdC2KN0oSIq+jz3IxPOX31Rq
smEbB3SR/ajvf1s+LvR4oNyqumZt9FTq7wyrVU+yQH0F6a8jSO0Rz95skyIhFHy+K5rrng7oGKbn
wmKQxQScK5nyPqJAAR2f6Pb9GEWumZpcPNO3vD/k5wdE0ko033a4c1mRbekosH+0lbKij0d1Rzqv
5fWNAfaF9b0xIv7s6OUoPibWWQnPCDvnbxfudMkG52ZwLkMCecKia15oaz9Jk0Pm9rKfhQuKfilP
ORLfWElbWPnBaDVI1/iBIoucAa2811G6OHG+XsPfydgb7bGHaC/jxsDN+7lhZeY4ESxSbtFnQlP4
R5XMeerTtAILNN0rwrF3f6O+ZEtUM8j3/ezDvft/GnwNx/DVMmbmgZQpW6Rvv9ar7kE0ZmMr+gDN
7fcMQ1DxBiNsFbvhHNj9Wb9DR0ndNUwFi1+ICjLnYroacqdM5rAN3cCeFM/dHex1E3n9kkX6IakA
YuPRPu8vtR1FPmYR2b+b917nxy6y8pfJrHHOyHarlfN+ZSUYidRvGCZHf1bVCjrhSi3iJzwpLqmB
yeavJmSUi5NCWWQ5m67B1/lB6lCZIAK6mikff2ZtcHkQkC24C75ZCz4gfg6jQReT9wE/BWBiM5b0
5r+iGIpjeXSVu+UgWAkGzTBbxnnixp+nTYPE1WL9Z1jKt7HNFFczSpKG9Xfzt5SkqCv8vqA52Tgy
N+Uhmq5oq9KGI7KtFareY7fCOK3LU8DZ8opsydZ5XI2H4PJlokMkRj586Y1aMgOf8yZWBlT9VDme
81WV72CLL3IvA4OhYIM/hwG4dRvdsvgwZGDDNVYxv11Hg1Ay8fP3t47lVpqxiIIMrmbwlQJaQuRE
Y82QWQdxBXbTAD8VzkwNTujSbaTivt0mX+Xp0OHrXHtKp4k1Te2vOhveYDhM98DrESOvGhWu7kPx
1rmE7yEgIf2gfUHO1xmJ7NSsFh9arTRjtvZL38lvwRHQQkAnVBVEixB5eEDLvrKFJLNG+L5TZM55
gwvMwqTyL4xhisZHgTJuOeWJMibcEAAjU4g7y5LxeaTNc8SToebRE06LquwjljVrMtbmJuUKmHWe
V+GUxIKd/1IwLWBqe9Io6bQZ8bTqhglvNTXeiJH0zCrhrOxL7QNoal2H7kyF40B90VaL6cHxZD6S
KfHCpEWq0De3zLvpFXcKhvIUhssG08T96kRNm8sXtxEoXvsnRcgOXdSP5LD2gBSv/fFCA09Suq2n
IyWr+o5PjyPRRjoX+E2MbhiZ08AZDee2AarthxNdvjTDZLeev3u4r3YDpnNIfXW4Zc9tUdQAK1q1
kAX6+OhW0Y//aVn4Ro6XhHEg+uKjaZYFyKLQQconN1Pk51es6Uz8SEQYv/3ReuloW5svfch4FaFL
Jgx2PKT7HAIoOyKvNsFT7jq8LCayeJNPtnxjpH/qcLbUL56Qc1BZeD5toJExTk3JUhICBL/1f2BU
HXi0xH+kPm/q54VozN2CYIFGpeUMTbCn5cJBFOsfi2L0fJL5ObQEmtC9DgjtVx8VbG48oS5NKyVW
xJq68BFnopD3XAajdxK6+HQDvVbi90TCDb/Y3Mjv6tTH0VeVXWNCKJt4RegzTDzbp1BsF9fCodSY
XVLOJDHUdf74+L9kftWNRnnl6GfeYtAzrMLCdBwj6hT4XM5ZEJapOPudVLotfNCcWOd86IJWWaQI
UvQTx1RnrT/aPTiUGtCFyVcpvSFV3FZIlWyuQ+tSarHgYM5EJqdY14TD6/HQXIb+0hVvVZpGIkfK
/o2zZNXpZbwkBY3XvoEUdjLravJ70zXY9+yawVZ66pBJ7u6gsrPgUZvw+IW5XBZyrqJmQocebHqQ
V8a5tes5SmiiAGRPeTl9bUwiYSnejROKZyIu00+HCUIDOKmNZGhVbik+HAyFKNBowne/aa8VWWTY
SzRBCd+WcUPnJcrdAPwuedJ2Oh9+NaIeU13U7w4m24k2myx4P52Q+SSVPvLj7dRsmyd2BetSKMQA
ZJhbGIsoU/2XGD3OyFeg91jLNA5+B/2rThWTMXHDaD7qxOaxLrMSL6LBjik7B0neI7GxgD3IESp1
EHdlYmuANr8D7FBbVyZfTSmtDBCt4rTFOW0R6admAZJgE8bHVwmKZnyJUaX1lO5TE86Juwolz1xz
dK9aVs3jLvnI0C0wHnsM81nJB8g6K3S5nxxxIXI+SiMIH4bTsGJlZHKULLqeI8uEusSnNGXugruE
zisEDvc3GKmpcj+vrb6I6OPRLPTPobK1yTI33UfPabPsuf1v1mBb+BflHSiGOpPeJZPn5b5wquCS
QsX9L6u3yDE4ffpjNYuXdB6ci52vmVf0/YOOs8o9tKGx1bp3q/Hm822GStn7/Rw3TbnbTN4SNB5X
nI9JjNkDvjzx1M5BPPh0+eK4x3pc67RHwIg/wZGpKujr64Pbb+0y09upeoAiWdHzynLpYRZLadIR
j+P9RhP1q9UCHtPbtwR3QkeXFbHFM6UJMw1trXVkaemBHDAnMGIMJGIXoDUPOnpoZQI1BIzjmorc
UEs60kB5CeC+1Rx9W/yDN9fED3Ma50wLTh05kJBIwNNUefWOEj1XVpeMhj5F1+qyQQqnmrC2W7sz
GMb3Pkhr5bZh3N2acVOxYEjSC2VC27c7JWahOy+ezv1teFi8oAr6+gjCwAg3JfCc7Owa095PYywD
vXs4MEDyTHs0bxH4YHDsu/7YipblgPOwMz7XVbBPYo5a6N226BOM85sTA1qQhWhRx3grTXU+CHZT
JyP34HT7UeBkde1MWm++dSNTt/VMWqn+//JD265S5h/NgCzEHf4wqia5tnifOiN8EuKp0TRBQZ2X
EfF6blWkWwYms3SV2H7eWFYAGK7wytL7rdfEWj1WRNSPSvifLoeoACaYxF8HWrkRFRis1V/FCjDk
S947uPqUnB/5DBW/uFKfD8L70RJUvu6u1HvGEhD7xDJs2GT9vLa2My5OxBE5pYfEaa8+3XgWKk7a
OBYSI81TFV0LBWoPr+TWy+MKpeqCyyClgTX1asUc6ekoaL6xt6hHKEvz/IIgLBjgA7jbHMXrev2N
R/C/blWA2FQQu4lrKwJhXPvTKExTm3sCyH/eUW0k9tmCPABAUyljDK67GoXLkqPA1wvKnl4SZe15
BinXoWi+QS9eyeygFQVtYrZhMdkddOFl37Ok8pxT738jx1902pZOWhhaQM7XhZX7GG2ODZmBeV8I
pqfHvLgqz9em1zQKDI9ZM9EBqASftOOufJJc8A/S3s1C/mujRh19Ac15NSb7KQYR4W1YrOoasM43
cEFbU0GUJxH273EBkmZKA1GFdB/5UJufvbvEUhVQsJd+RZORe9ZSfk9ipWj05BaAIpv6K71q/yhy
NIY36knukhbKtu1dnPR8dJsRxhPYRSJMeoZ4Gr/259B0l0/QzcO7jes2T7hZfqTOF8wYNW+QEt8T
rloMtQZgFKbTXPgmj9vnBEoIEu8UV4sOhae3iM0SxJIBgbWq9b+0ftzAjzBhdQT7xXIOOVDTbcLe
is0bUscYVyo6GkD9kcV4g3YFGtM5dSnvKWwhavTRMO6CKz2MnmZQqYUp5D13ApYHxULK0Bmxa56K
mOO746nKvqWtizEjEQ0Erov6Ro/atkwCcWI/xlcv1Z/4PoUKaLPM9AxDv5Zi3u5y3lAKEHa1Q4sC
eeuHqlEM1gGDqZ2gWtT8L3l2Z1uUUlGCyOxt242OoT/PXbuKQLSqL0kAjBP/TzWXwlfOznOPLM5e
Q2oNBYUYiEUkgQnlN/ZnfB2poZYHVhb3DEjjS/WnWWwNGzbwS3NM9SAGhRfW/8H0MizmMuQfVbrD
GCWFlR9KNbGaks7G3O+CU8GrPc6LGtUo15cGVzYPEYQ7NVvdZap+S3f/Wez0AuVL7w9+tbL1oIQv
8yB65uk0X4oiU1SMSpROoulQObKDwMgqvvDSiOY4ezM1H35+GUN3r7WUdyTRC/m/eGUYpOsQ9ek5
lvtwH1rpg9P6SnPfcMyH3HQHTIyVDO1xQglg40nMS6uctIClrsyznrtrc1TMq2k4Lm6oebJHf89X
7/sEzLudeqX2tsSrhIegMrrxmk6y9hHMkC/npjH44JpkPTXZ9pYGIhLroAUm6S3fNic75KPNpxlF
MiTXCYRXpwQSie+RUzd0XFUUc3hYchAXCpOZUqZNYgb0VnQ8+sOfxQBCE21mUkyXxnuyQNRzHUms
1BYc80WOpvLbJcM4dzyx+qasSsEzjJm/HBUKIDlzrDfdKWMkAnT0Mw9mzcl7tdTImseURLCIHFVb
EUVAF49R2BfjLFzTo66U31rw8AtCelrBHDPCBgbLA+JfrL9tDSf7gvpVrY8M2PM3jd+a+H3/XhER
WR705zcVcg0elXeGmBjMqVK3Im+4stfYw0VCS0YRdOUIfMUS2th8q1eF73Za//LuhWJ9fZSfzWEr
GxPcIoP4MkZ1HSa0eA2S64GZD7dQna9Xv26KzgCOeadNr4a5G4Tnq1t0ebgc6Tp3UkdKh93Txyb5
sswap2nu/n6YcmFOZy28NI5vvaOjxFMH7yvCPV6MjgT82/OKGn95sEAvZFFFNamsTRZZ8MdjtdfI
a/NG5XeKBvNOawf2tpxQEpwubfAAhCY4CQLIQlDR7VqmlYtda7gHOs11T7oX2mzRS+2OPzyqwGkj
2NoeyS8xFR40pB1PYRBMJnxDywvDpuZTZ+PvkdCj0CS7HexY+O8bO8HCLvOxgWyA1RdPb7ySb58k
KMXv0xVIrEySb74QIMlkVFvzefPt3qhqI41vQ8WXs9E4ksLhVno8DXLarkK5EtP3H0FSrd2at8uK
gmROKguVJNOFY4Zjqjdix8scdEYiJjWwsUayjJylPmKwhGUOhNYGwt9vecXHVj4wdEZzUm2we12V
zXhZHIiCb/Ikd6CFk2WODDaT4NVL5vmVfJAMRdOQEqoOZB5G+VoT6piDpqskPk5CUmFwjRM0Uqif
IzIm847G4fwXLUESDz7XIoBdoevrj1KshXK7ArjeEgqKuInhfwMqTqVI5vo5Vr0t3T3FMdGeTUSM
H5wJX9AQE/wQs4PpWPVNhyllKFOpzo+SNtGVS5rMiq/KxA90S8zlE9JpHuH2HYCcaIehJp9DZnrC
zDfI7DP8yk2rgxMs9ArDo9dutdSp+FwV+8g2AAOcKAeNTInka+FPiehzkeR4JczXdJrTY8IJrePb
ZkK77XpoIonUV9HvgdZoslroX+ft5rUgkIL0aBoO7G4I7KWAsoqPJhKr9YUqnVksfYcNd229I+GK
R/jLNbsP9RIKRuRvIp4+qzReEMjCIqxUs12r8UPYf5C+1yWbgpj2GaEUbWfWhs0FrJWefxxYeyJ1
pwrJatvRAOEUuSfq8O1DWgotVDHUT1Q6pxbxRbeOW/VSjMGMB9CJPpR25y6hHxjGsvw355NMAzhU
WhDq1mfYj+pZJxrgABhVVRopR16DDPJTqdRYhAOqbBFy6+ScoIDUlxk3UYOKarK4WMkkMXzESM2z
QVrSqT40OujwOyo7oQ/o00hgJ3aBn9yekD9EHuThev4UmQABqchtBpXctVGuST3EamBrJClterng
472emfQKb/gGzW4VWvxyMfO476eZpPVj5/o/Ro9Bz3Rhu5aGUT0bxAuwRb1PR8IR2eB17dDe7FXT
4EA4Gk+0eN7ndpYFg+34VLBma7NoVUGTln15W6jzIHs2CDMf4fUfksO2ULsAun4pSDWbhjMAIbVa
AmZjOWrINVfsPl7qOMK4pFwRa1Tdn4YHEWDAI3Gax3hcMc0iocNLP74/d5DC8LnpNo4vo1T3NiHQ
VEKxn2m4oZxrRZJItYV2GYYv/lPkobotpEZlj0o+NaxZQBGgTG3el1Zqwiza4g/qAj2YFfQqb9RJ
dGsFlaw+EOP77kruO601qmvmHM/LcELBEU5Fsmqp0Gie4z7zyrPkoxxB1GcgTbnnN0s4UZ0sGMDH
xbZ6Z4Q6PGL/jlL6siJ6QwDnAzqOh1GKNzWM+Wz2N8ldVliNfOEuTEokq/kOnmj/cO/0nnTFF90y
hL00j63XAwP1psNalU6WVYGyuOl35hI1RPPToqGrtDYPMb4v2LFSLtDfXXa4Mb6O9kYLHeyq01qG
rm2Ai5IrOhDBuwqK/jUlc5VqxQLXLtmAOFfrOAIE8OQ+jWW45NYx/zaQg3t/6MKXlQl/pKndkI3K
x4lMUTNA1qklCBq3L+LS/KDfSZlZvOJ8pWmY0YEkdWlN2BUFdiWBsAYH3/Pr9Rihluzm0XOsQyve
rPV2JSdyHPi8i6OJXqkiED1IQp/fnvOzpukhzplDd/EBgCEbkcUrpRGIR7SFLfJnc5pEAUAecdIY
MulngZ6YSexXKyosu9/TG5XoOp8MmliBKIUcTxuJZ9FYnvbIIG7iuzJlIaxLQnjpEIBzMNxgoFjG
AERbvCLo6ETmsnLoSpbIKQUQCLmhM+iSFCqO5uvCC1MHzuIujBQ0W28tvlA3c+tMGUE2m3C7UBE8
Tl11ntRed8eFwoJHaEMkGMlQsQMPf+XHFMwjaXkwSAxew27BTPSGq/7qUa80w7bLO0ZTW7I05tWn
GLj7mukcZda4gdS6SJy0ILB2kzuMIVqQqPJhm4pSAHJAea6PQ4l2unxQvm4/QsHmJv9N4nG1vjWg
aqZUv6CPKsZ7TM2OWAT0pCBBqSHBWDlN0+oqrOpS2OqfmrUCrRupF+8th0APNiXxdNmysebMtWWc
IyyIe0TRsNVP6Khrpdni4TSWac1GyrPZigm++xH5yXxCXVpVw1z3LKfBou9uC16Kyo75XsOiU1Ki
xDrHg+Abtr/+1s7tneNTVnkg0dj3ttAL9OsIJAYk3vHs/KJnuxRGlZI1tDQcfxtVJrilMdw6Ntv+
msis8Vao22O3qiqxQOzmTPalEEH6GKxoyL8svhS1WxyXcEdLDqGjDsgPtsG1rZAIfLcGm7OLG3aA
dWC1Jb3wW8ROVRAtHSiB00v0Vh1YUJG2J3eG6bfvODpNpKJulh7JL9xtpJBMfprdKjDtlXemf2j0
InyvNrCF+YOERpqsFB7Sxl0x3jCgP5XRewasvo0rCjwvMwfvAX9VxPVKK2FjakSINNk8FfBIXI2o
R5EOguFPyeN3xtZjBfOwWgoH5+39H8T4NIa1b3RAlEMML0YMelMd7SfnQzeJPUYTHFOokh/Hx27A
Cw5++KTzX1o9YXsZhyaZbODke70SV7fnvRdPlKnKAL36KBPhsFULZQfkNJGQnwFruZ+BueqCGBP/
YAabzFtoOgDfiWurpViC4vNKVNpW1YtvnFfu397cY9N+G40UletCXdgXh9tDJCaLu9o4jIvLMKo1
L7k6zvscjjq/jb89cN992Mysqy/AycSuWk6VG9kPW4I1VyUX5hW4YM/KZ3NakhmjstBY6WDkW3e/
0dgjqnCoXurFaOEswyH2HxG5bkqiv/PmeBvYqd1njoCNH1uJ4ZBy94+KMkGGhUrzEJukkYzz9F2a
FUmaSMzpmiUMTijvVSoFY2WfI+lHv/+CBZIIhtVY1p5nDQbCGISXwKB/CBB+EoKFc+D6u2H6T9Yi
HNKZk905OfDzNjJkZw758yb8dFaN1tuVhuCZZvMIE3KHW8z9NL4jB5qLfOCA53lKwQ5MWSHgJ2s6
w1xy3bG8q+at1fd5Cmj1m5Om9se1qR5v0GXMe6snp27P2MDzMp1+MeUwJSTcAI1Bt4+sQ8Y8RGtn
yaEcZtJR0mpUJUf4416MGZnYs3/E2Rf71UYsbEMomll4BzmczlSbYElvXnLiKA2OxCMgnYZhtwak
2rb6nnsfkdrfkWU9Qgx6NkD21zMbtOcBsUWqqP3yJ321zm1wPFrwue8qJn060qtO3CYPDJgxOE9g
Hth35gGv5aVWUkkV9AHd+kwgNM7NYWKs2uXKQVmYWJDI2U5d31UMfvjRP1juEp4BucBh7LQ37pRJ
Cvpar8lKncWSoc7mtoymwETK7E4iySkh7NUNmNEDRyTVbzCqhYNT5t2FvstkZ0ockTG5PLHAR/DX
UWjHH3hwbaIWw+n1hwDtBxfq75MrH+4c+3PDQjWLSvUfOmT6bKyOcEXh0KUBNGPr1XxoUkDZpwFq
QzSP6FpPKpjUGkCcJJdGu82Xp+yxYoA6vImdg/sx+ywlQFrorCFXm4pbkcq1Ha8/2Jga3dboIN7k
6mtK8RPK6+ZjQrl1P2ALtNFQG9cjbes2oKR8wg7cGuq9bRGkf0dK0dewkj1JjoofrUADF5wlHfSI
mBsH56EcmLmylKTiiowHZTwBkGStLNiZoPii33HuusKm/0srWZIm6wPMq15Uxpji85evFDZdJYUL
xBPO6mPXIYAKhWCDtXvOhaJUxbZGhIDwrU40zeIgXYP8aga2TCUMXNeAebq5mOTIKew3YmsGvOC9
KJ+i3L3UioVgivItgR2tff32i+XXSKB+5zoWFH9/UJa/n2yBy3RCUtsm2EkvkS6SziVlIWSjccNE
PxKfhdlqulbhQp2l8opd3VfjaYts4m09Z7oTRyLPeIpCKdAW/V3ICiGcw9aP0dxR/DPMs8RrEIER
UBED1BnaaOrM/LrT4C1KpSbQUittPd62yBza0O09hoqbCkgBfLj6S/Y//N+FrzDyz57S3bxt6U6/
H2f0T4rXF8O4zRW9D6Fq5e1RzKB+6AE65R5gCjd6ulv6yl4RN+k+Zt7/A06taDHDnppPIsOk37be
RJnmodmUKp0OykK8yiSdsreV33kynPWdOdGtZp6SPT6DZgV55sfKazvIwGy+yLS0yhbzpKh7fvom
swvQ3ZWih7RWvAdBsZYZt3sCmXEq5lmssnItGVmGby4ULBYWdUuCujffWl08DJ1Wbp+Uoee8vVfD
oqOfiTui8UJGGINluR8+X0H0Qv+JTglNK8IyxDkUD1M1MDX7XW9xrwSXmI/ZCHKwC3Z382seFihn
kI50s1d9jiIzLfii+WEf3HSeqVpWrkf2U2SocFBoKv/+d7GGHp/dbRnW2hED/hEzQVjQsmq0cfR+
GVphX8neuwr2JN5nHp5L7fM3FcnAO3Gry1L+qkMkDUjGZJUSbh8g5cbktu5fpyuQzarpcypS4vDQ
fLUE8iO4loJo5HPoPwpZUt0ny0M+YF+TgUh/3Ns+UNCE6c0u0YPFc2wddzRJqtZPLNOOzS4BYMsp
yKAW7XZTFX/eKD6ph/Kq4pHyscyLwM1iJNCAw6Wc848XjVN0pc1IVZYaDyxLLhRojncxEWEWsQMc
bu1gRfA47VwqPQfAve6dJ+sgQwcVKzhOL8vFAXY+eJyegdRSxZrjBXAtQrCK/NtpSJ1enqZ/Mph9
LneAiJGtBFdIV7pDgUEWiqr1f90e5HhPBP4t4mMMhP5oLik2oamVhhhfR6eXdTMiezb60rnGbn19
/nD3p9m5QD+Uvc1ZKWqA4MfSPhHny+oUpgQaDEhU/yosOY3o2B1Be0viv5sIaoRQUK/JG53oA1Jg
tQ3r4YFZdY5zivV9xoA7ZCN+0GO/T1EUZ5+G3jfj8QZIquKm2YcA+uYc74iCUYdrv5cPdsIunN+m
qufjqBqg3Y+pIlUPhNrCAFyigE5R8VNH2/WpRGACaaDpQBZhx+jcxrki1Pe/MpAQRRYPQRkUdtvt
u+xPPRmwP15fmtK9kaPvpfO7W47nT6ak7wcPs46R4XukwSSoy+5Dj2VBHhtxC2SF6Zc0WtXmFhiO
4PXr5GwDgFEtfAH2hEDYmppuLev4S9GGCCTbSK4qd2z5VAlCuSntEzT1BNJzteJmw5d9KLKkp28M
FQF+oktA2qNu30uzRyP6eQpRFiYgyQL2m6V1Ml13tJXOR4syem+5db3t5ww7x0WlTS/FNz4V2Osq
1+M+Fl1cORomUtmGZnsFtjVCe/zOtyyamgnkIEHRp7pib9oSuawh/Fj3GVt4/i4sYNhgQU1E3tv5
zrDFO9DhRTjODxwWv5zrTQZUdHDiAW/YxbkdmHw+tOrPUsD7l1LcgKBooKS8Mt6ISUhtD9Bu7wV0
NFJylwlHr6VAjn8O++I6aWFS05VZ8Kf2YkMBL8NTntj05lpAXyQQwR72ZXQbBevyYYNUCs5brsn2
ChlDMshAzAwS3iBrp+VKetgHAo76+1Lh/h6Obyn/HSYikpp+C/dzx0CNDTDN71RL0fha9XuvgHB8
w8hsnZFLUmKni+R5Gowf0gTZFw4qh7QwpuHkFUw3qV3XbbbHo7/+08SnUX82RMGEzdTJyv03IM2s
tifNtVAE+KOnPDwEKFqi7xyArxno22uybKT5PNwdzA3mTO7LTANkaSEXUzyxs6G8YynNYQ78+Bpf
D/bEJjCn3ylSO2cGcCcclI6eD2mBhUtxsoxD1SFRMS2Ghobu2TDBVoJ8+V9tK+FbCzKzugQ6Y2Lj
IUhert3F6fuaf7P+rD4ptzRqXhbx71hUKEIphpYcHiSXkrCxmYoseYoulgz2dkk1AohNrqwL07V6
Jx6wnEcR5+OOWHuy5QAN4uzPdMp3+ayXOWF+e09lODtHMMDj4sISNA3IZWWL+FC310aa34T3ZRBL
eZdLhhobeCl3GFbTCwGn3E5W73tsFf97S+LMX5W9qYTmPqviGSmB+vFm+MOh8f1vSundjKcwwdoc
+kHhYXrRu8ktQKSdb8AhP8EW88RrwRMWIrmVnUCkd+mR34P/+GpippOa6qm6pTLRYAcDMlXYnbrC
fQd+nAdU+WOWrO9fDS9kPJ7wabDmetjuTg2GPTZwzs+2P+OwfOmeX3RWidn8T/CEIW+wLzvKCoxU
5NQrs/xJ5n+D2P+1T+AMd+ElqL5e8amrSq/YLcfJ67N/Z9BFyWiXspmZ0Mn14PcBycB+q+t1cAVF
Z424BLYS1GXqi6WqFezKfbPX3pJTDGtAqJ65QTplbozOXiQF39rCUz4x21WF200I1K5Hgd3lnrAP
TKr0BXYgPjJON4d5naWPiLeeuMzUGTKpfG7FfTsN/NK8zkGUPPuYF3iwU4FfZln8RlT/8WnjVnN8
O03RYvVfLd0vadG7vr033JQVjR+xsalEEbT8dYYTjuhRm3vRuar31pO/qqFPzyOQ5/Cc07ACXzMH
o0SWs8lQTHDoTAhFgVu0wzK3UYyv6kZOXkvFfMzhfI0jsWv47KPv3eZ6a9zrVCn8Fuve5zpF5IJX
aH3eJM6mM1aqmMm/c2jwpqe8OWhGGmgPNBjvpjawzlUVmF/uaraWL0odjHrljWk6kVm02613NQvm
mU7DDzYpiJSDT3hEracin7IZ0kZykq5foZg4vGZlku24dfzswRjJ0ivoMkjWkmVjaIJTujW07kxc
aQ3lB1ZED4XisaQXaX/HvxAtItyScN2rgcSpWB/iINnRHU2I9J28AFXqo075VpqqWh01v+tgL3Oa
/ZOPH3vK9+HmTl2+8zKolUCzdS6GteTso05VvqDDLXUkg1xdygylqI5Ndf+d6F/c8BXqvDXW7SaD
ysgTBPXre1TRj8D36lUofBQExtZ6xVRjpNQJrjgZ3Ai+FVc7pXsCw1fwENyMNCO+KwZFL1dYE3Z3
DZQ2vkHTBN3qZCLq2DwoBSgG6g5+GM8ov6Uf9SZnt+qZe7SZbY66ItaZCOOZ5WkVf7GId80chVtN
iJzw9ijf7xvFOBwzdYbV8b77YNKyc+EOVP1FQbag/nqFY8C1kvMcHFmGQO7rJhCACp6MEih0IS2B
BClWWsG1YbumntNjBaKsxuTUfF1N/iuZ8QiXlMQVrsrI7TGQyxPzpDhbXV8M43cSgKsAnkgsmxHZ
K5avukiqazGiGsKyjry2XvMJ2QMg/QSARBTd6okDD/CWJH3DkpmbE17kyMsu48z9jCLGjLS/m3o6
kubBYn+PMw5KW5RkX372pJqQ/SgY59It25pSJofgQ1ywO6AIRbxLrGJnkM2dhSYgNvUqhBsA3EOK
17Lq7ghm8yYb1Il72XrOzQO4JQlGiUbzQQxVrcFr29TEiXZP3WgXFDttymXccTdVXMaLo1/RV2nj
nVuAYLbRtnJcHzhhSfoTTB7GVkLBHWJT6j/ECp6Co1cNhgOVShAfqIFEOmOtxmz15GiwAkk0yhx0
CsP95g9Oro77CBC4A7/S3Ext3yGTsZUK0kvdnEZcDP5taa9XkFWuwnzk/AXt6jIctZSqn4VCAC7A
/GqXGPk2K7ZkS2OF/SeLRx0Y3ymQKIZlr+FMwt/Yd029kL2bJ6PXKohHWV1wuEE3oq5/P9TDpn1B
ww7m0RvUEJBFUOFX5yurq/rwJk7qdK1fitkOMU1is5eORH4wbvbMuQsAvC5glLrNfMQFImdMIhdU
7T6+YzdxPMV1v5XQmlf/qCMUZpVur/bZ0TXSxtwOwrEinw0V+asZ/YftlZnXp+edefpmsRIPpytr
6dP5K2DsAKP/2fKFmhlAnaRIyH91fTczWkq0V22pE5VYVg8xNNEyNBRI3rp7J0OLfSw+rM/zmGVd
jetOIs0aNFkZR4S6uV/qy66lt1rODT99eM6IcNHaZBzQLBRaSjsh8sCliDB1XoPKJCH8krxAtNpp
rmHUc4pctUK3hE5zloxTXtwRDUmvMTmclnFVQkCPHxyzWWT8iUUl49Lj1D2GuMb3eoiCX4YKiqwA
R6rwJT+NVRfrNOigGNVT4oZCdqCUatI4gr9vTlHNQb5NonvWes1PpmrbIipuo58RLlYj2ehu/2dz
Y7v5ggr3oQ/zTrJaglevawdLwtJ30mz7gwjU0hQu/bXa52/vQf7ix0cwaheD10GVk4hcw6ruYgYd
rRQo9BfxYT1eOhrckIKwqmRV/JvBDs9/1AsfVKX4AXu/lncaTQPbdKI/nynSd4Oy8Kv2DsV+RTPx
qDEjvnuWA9jwxF8x3a+0B+H5yHOIp0az5I4C5SudQgyDTvZheOqOpAFhd4W7dXpe8hH7mg3sC0oe
PgjYPNzIQ6xKL0+EQUEg2LsLViQBvihSsTm7n/kZRRMXd4hdizJAAev21Ctn27VH8rL2FYApO5yX
QErzN8QgB1DzPIdjbKmCirUAyMtmafAkNIG6Cao9LC6/ovpgWYY6WHnovBNQgd+as5pxIAEq8cii
EcdXqGtnD3ULDO+tRo8aL+WxFcUYSEQ6UqTu3khkMyv54hAxPWm0tByPRKtoegN45tNiSCkrzgwl
aaBvSnmIH1lrA3GS2ax84XrJrSXOxyWBgzBx+ikNrU3ph5DXHQK7+A32Bb8RUkK96K1sPsQCmAZQ
KbbJQrkCoMQpgNRBIaa/Hfk+uxq0ga0OF+Udq5NMA+nwbPOMCpn799jy7C9sofhelFywG0QvTVEn
alkDTa5hBeEVpNBiJ4ELgV0qK2M4oYLU7qRf0k1/JtI0lTKSuI4VCaepcOom1/gn9Wiw41+Ae+en
J5mvFru6s1VuI4Ch4da/dsCEboLP3rAkoUsobp2debPPjig3qbr8q7HmsjLK54j+EKUr5WO6yysk
30FS5Yqo9HakTjCPA0b7+2smSUZxUv3DkJGBGPhtQJaDjjyoO/1++HWvFwIAHnLDNmEa6D1AjCMN
LES2RrQDwEoazw3VzB5Lvfpv7UnKROJoOkZqkeruYj7N397ZBQpFzevoUyowxgRjE3zxx/ZKXJrp
ycB0BM0/7cFpx0NxfNqWaeUafouCPARgpeqyraKTzQ8dnbCUbCkprmWYUC9vGwM6unNrHgIYu+ap
VS1bw7f60F/sHywN1kQmHzQV896tpieJ6q8WT5Pt5fCj2XyO+DOYk+QkYZ1cTuBS4UOqZ7kBFDPC
2rmNMiabu4dPRtTQ6alrvzaMqxOGITfbt5ScE1XxenlosCtGjfLhwTAy0lgR6vEXug3huyP3pG17
8Mon8d80cgKMXhNFxg8iMyrw3y5n2P48+xbMntXRFB4MMrwWX2J9OpDMajFqhvNLzKVR0VivGjZa
TlcnQkx5InmmhQYreqL9x3D+hiesT83DQe08Qdr+1lonOrq6561640fUpRDU5bYhLWHNE6V25o61
SjocCLciAL+MOSdpwPTNU4giZzmnmIXCFsOf+h2ERA1P4NNQ0HJ3RoITn5+dDklEy/nAih5ZUAxa
OCG/JB+vrnjqZW72rErNjm85+yGxBIne4zXVYwPXia8KCs38EXK6r8n6TEzq1kG80d56dmUo6Klt
wkMMEFWsroaJ8hiVIueQq/tjkRTOy0aM4rx/vkn9Lhp3y/YsXYXeupJyGoqgXdcey6+/pXTTyWJJ
nDu3x7r8l4tdX0hzv10FiEf0FxkW7DWDxuknKJvCYbCn6D4N2ZS1FEDlvIVZZvfSBzWiv8mWcXJE
8Jg/iI9seGzXArN9jFtRdUtLPVfyKB4m3W3RC4UowVJKFa136sK5SA069/8gfN2t/RGON3hjVY4B
I6FhSX6Fw56rquldWR3DJnjiKWot6gIWZD8BqOxh4lQ7TRL9PwzMPoXReLLyppq/cF9RfrR/6WNB
RfupicupSbXor+gWQ/ToqTJ96Z5GwAoum4dVQOWcuxY8HgB4e8rXh8kb0SpYs35Uv+FbV3jFhaBh
YS7BG6swj9nipB5sj0D+bGtGU17mBZlapdn1dUgRwIxamre/eioGk3mU8z3pXTgdMQYFPCoLzC66
CxRiKrdaQs1yjM99bI/mwgeKvVb8BrigePupTRN6nyDfNG9c7zOhRDms8zk2WWQY2fqR5ICKRubF
4klPGLmdyjA5ORIJA2PRnetNMOU92jz5zMBRIjFpQ0cfkeREEw8KIN2eQbH+kXJ2gAE9REI7z4w/
44VIQW7rmNTgbJk+/M+DDVDC9E/X2nC71z2XMdB831cK2/zftZEmDSkLP5gO/PcQJfiecO1d1DO0
Be79PbzxKdbYR7kGNtUpmqSyXeESKeVwGbz+tu+3fMoAaavwkmqHG82Q91S8HQpUtYVQJyneVoYv
unybmliSQwaG/svpqkW8kEsM8q7Er02DJPBpggqzSUQOJWPEB8UqrT73+s1Y6J8mcxot1oHnTery
wQQUh879yX0GqtuwnoxAFjubbTGwwjzuEApXi/97Nm9OZVAix/ztSGRml5ZbZrNtNvt/3fEQKRh1
KLDoseX1zqH56nhVVhyetcyjEOAuVz/NNjuQzcvBePT/xRCO8zX9Hgb1BCGxEIpnEpuVn+U++8sa
YNxcrmWB7yTOwy/D2ptXw/DvczV8P3NQxtAjWs3zwEbB2Qd4L0KdoByO3pKvKJyJs89+yvEo55qu
2ftgknrx+zl37YN4ck4WDRhNIuotXAQNDFOvvEB0vT/9yGNky9/77W9+mkwZaIQYL2UsdyHdZJLQ
PQrZgQULDFMlLt33bqFVqHN7v8KRt3ULJrZzfE67FRkQer3MfMQ6Xxfu6Nw7AIIF+tfHCEvNFCrG
ITmeicPRFG/MGmTfQe7q2Hex8wf1h6juA7Q4hdHtxkMCteXDLvIn28Ak+RNzs/DiPHy2fSZXXRTC
pFTipSG0/hh8PjAhiQSTPnqoOdbEESoBBckc0uaIINoNMM/KBmhaxKhfOSvN1rAba6YOJUjRJG1K
48vB0bWjYmVtnwmBlVMhMWqmmnQUzKznK5UPIHxQWw+opIWhpkMNIJnSlHGjfen8LjAPT7fmfxQH
Nhn74QASsPAAo6qvjUVFVkgiZIG8ayuXj/2+Dlje7ZLrYEHqCW6yEjoIkjub0lFq1ic9HF77qYaK
kpJkYVIqxWuVoy4smN9R0yf1rHMJ12RJ2uwMjeR5BXDCzEhYx6BlZn2Jz80JsOQWjdqePdxP1Ttf
KSYNKj0wVXknU3FwtBbR5oDvhGaeHIcAt6TJxz3UVLNrNzb8lrCFL7g7KBTG8LI/AJF0i6XN/15i
gPQp1wWnzoYFnl1l3/gqZIOzrwZmMJMYfxgUi7e8Ev5vCkAKIrpnNJf4VADxVxEkhTG+sfXoNPY1
5BWX1mnlPzeM8T31Z3s8QNyZpKd9ALNJRZptfoGfCWSHWrSncTTk71BKIbw6Ye9+qhGRGb2zPIaY
jBtX+Uk+AK9xAxwZnq2D55RQxz5/0AZd9lS/a2bZyASdanTu47jiw1ocs8Ue6qJJOw2DKOLn01V0
5C65rIcJ3xsiBpZ8hXQ78A35KEAVCmTaTjs0XtIGR8abiPej8fe0lHgdW/BLklwNf4J5W8/8SzdK
Jho4iayWeAOZpMbXCwNn4yVrZYL6zSanBKgrx5oX/QDgOymafphBKW5nf+zqZcVlonc7xfOJi4C0
7lAvxhbxwMCQIwS7h9L/FSjmeDnXU+Ui+mjKOC4rHBOWzgXLu25TaCGvyVGGYlzDREQQJRPs07Bl
JnASkjSRyoFh0gYjWUVmBIm8qTnayOh36MwBv62omMVYl9RTo4A/FD1bFF8CkOETNarT0sGBdvdM
eCyL42IncyLZ214f7Q5uyuz9npKFSPom8hf/FXaJHZZDPqV1+1r7VNMBHr2iCu4DMWnI3SrzjwrQ
B1uCyZpVSRtmqKYWdHbFhnFErAKeLUDQ/MoEjdwoBuTJMbNt5PxqBJxhhgo//+Y1GApwt6294yu1
FVOsNnUiGsonT1FxDTFZsWVHFWIeibnx0puA6TfrZbXUTJM/pINys0DhUYyHW3/EF2TBlvJ40El9
IBXuYyQd7//TV0Am2iyilexekLHyMePUxMUX6/pYvBPCxZQCDsoFGo7L99rGa9ORjL5LwJICAbnn
WLilWx3lY9DnynhI0AV/5De6zk5LemSmxgY0eI7ow3taMTwwIbDKyigSIvJGfcTeEDv5hVDy2hBa
4xG1XL+WAaZ4aXZAEvX/iAmOPguMHoF1/5LJzuUT1JOx+X8joSG2idEL8YOfdXjEy+u3xnVOoGXh
mlTIltG6xKqPVoR7kTY6ClfE3xYiCj9Z+DZcakdogn774MML58x5dDcz5RvzbHSq3iiC8/XweoMp
VvtYWsM0Ts11pzI6oHynFZpjfvwWgWSMEdEjM9XgQ5Cr15kzAjzKC7MAR/4/KKlh6lZb3875J/pS
YgxWWxOg08JQTuoB2OwoCRMKH/6RxvXtv0qcHDZPzC7fcqpPgIXacXBPDZIvQVPMhFXQtPkLB2m3
SeO1pknNYETBPHI82LVLYlkxi9jENFCebujKdxxspjoVJP9diyavdTi6O2h2tOjqQ0WMDGKb3RUe
Rea9srgfI1sWg/aAxnrHxzRCbBOl6rdK/cSS4WTDL9bfag4fotXa3IqiIdpZCLW88WrW1TnqY9UF
0oE9c4NKlCFjbIGjHd4DRE1F/8WJeRL/v1bB3AGAAGz3JoXyrBeXnMTK5K1JxJH7tg2FlZyCI8/W
rhKWFN9ggdDrIyiJjH31m2cGHdun8jU21ctHAolbWuSm5B3WcUtAgHYcDDF/7jsQkNX9FvmEOpUn
OYBwDKpe6m2UG1QibfpxeDhhlBkeqvc816tb97BcqZ9rGYJYkZhZFHYjOtY72eZzgV4fOX4/mczf
DBcdMDdbUbT9UkBG0SOtPLzn6U9wa+C7IaBUyCIMhYn5OlEZGWuJkDBk+PaQIQ+hjbCPLHEYTYhf
fz0iZR3Re6VMPX+cJ+R0fOsfKleo0NbzVB1YpJ50Qu+GXyzrzZpwekD4uydSu/9DCxWzveJZukvL
rK+znR9GCEe1K1B7PZ1mNacyV9QRJA0l5pb767Oe9EFolV87tTh2xb7hOQL7q7ON8GmD/edvzHM4
X4Ql85e2ZU5mYyD5rcoKdR6VunML/KEktOWDr26a4keQ4pa80abQFXQpRlksWhKRuPIpRSHdb/d7
9ouIncMrYwRc9wQnytxHCjPWcoJ6tcZSZZIeOSH7mX5jTrARlmcZQ2JcoFWRqxLBAsDwXC0l6EAo
810AWuB0hnL0UR+D0M3kGRLdV2ID6m3QhneAczL1MSICiBRmkFvq9FYVNRoq92vpHVuJn/vaDB30
3dpD41I637sjfR3OcVZgYjfRthAwi8bH8dTi1FUNrOYKnTdnHZ8wu6Gb91rNNVaHlYrXHfeZCQwy
KD7xEpKX7Xxdb1+uGxe/iPaDfjaIjyJjV/LP/OCvrDKIcgT0ERFXiYmfDoRtsy1IXb6u67iGwQv3
IBXx3vjMpOJIWCLfJAbXYLLQp41AvtWMFqkLfRUDL5dTIK73M03cYGM5cAEt4TphfyBsD/fXhV88
sfGnDtMveLGA1gk43Ycj9N/iWAJtTSHKXaP8D4JHVa9SbiFnRGGl2JsmBJLXGo/jPqrGlS5YvJsF
e6wQkmzMs2Krc+q6eI62E5d9DOYC/v/IFEJBC5SeoBwso/Znr/lblDqEQtLTDm5BQO3+Lb3ZH8xH
ANuKkxJ3zg6ZYdSQHaSBtdUraxq6ggG5loMOwz7Z+qpqyCmRDzZkdTsu0LjA+loQkmYaTrhdX9L/
bIGU5uMaheVhcOkbhFsduI2GWHMzLJxZl2TfM5pc217iGfBneMx5OZRH1GbCCvGk3ERFBkhi8d2h
ikQUmDTseLKTbs++dQQ28s4h3t8iTgG2gyi/CSAjpzMeHtgblI65z0DiaF02XRC8HG/k3aA1Nkdi
irCNHdihhl9sVQ/QsCz17R9nBhQKYoucTFw0T5x16l5th5fj3c+2TSBzc9PjxU5Xc3cGiIgXdnJH
hFrC9zWp2/iS8qhecVQsjRGFW7jaZJVPgQmu/HzJMlhfo5VHulHSJGb/ucUcqcWgNvZVVgeRhxjs
6s5lpSmbNiYII/Uo1tWe2Lh9wGr3rOKJYfT/ToDs10rKz2bJW/9k4qPGQiRiT3wcMHszLSXGkwv2
2d5rq7jRFNqzYD733gh3WHplVIsJ77lbCW/osAKa2inxW+Xvl7nXywKd28kI57GlZ3wIdi07AFKc
lYOxZo3Rl4fMiGk9u0F31UXDcosU55z2MEwxZvzAfDuPyWyPLfGlBmQHhraosw2Vq7jDA3wwfemw
IU8k6kEXXAA+BpP8z++i0O7Hr1giDYqqKVzfo16Ojo9mPbjdjEOo0cyfxPyCmQKPdB5htE8QiFF/
KO2Fp3cVgH3ijAeQjp1qP9CYBTsjsPYijXIwR9aryyIQZIPThR4HKmzB4+fXE4z17H3OQ1+dRt5Y
2kS8HEryMF2/iCuPACs/uUTCmPCeA1OzLgu/ihq0A2+0dzRjbxRBRVn7ln0Qtwr9/67XixQUUGzo
sYCL9thGAPnAIAcjNF+z+SFRgF0nFsEYGQv2pLsUXCBC9UeOnr30BzyuDN3Cm8zVyDfv20uOzejp
UazBHXdpSgn4r25wC41qAj498jI8HqmE6mUGe74tzqwk+uCk7FVmRNfhPlEi5XDPE4/kRZ5OCISb
3w8FtsVZZBtErEnbI9rQ1L50EjqybuPCEyMKqZJFu/P5DGeOv5PB0yokfWb29I6HPtFi5X5KcLaP
HikCxuF9UnoSB18wWUzATASRrANss5031ht3yvCs6RzR12wpdp52Ua5hH7rXfeDdn/2+3E+hSXxC
s85m/+cXmqRsFYLgl6h1wCCUo2Mom+QlNS8nOAF8fa8SdNliWiGBbskP4n7qKG4wlYjI/6YCkL1a
tG4F4Or4QGpUcEBQEsdk7+7vsjGfKMW2C66stTcw10fjLW6jYL7To7sZ/XdfbLH/3fqWa5Uwv7iI
hTlsKgjXbCXbfpOlBal9JRra+LgaEmZ46eOlIB+KBLG9GOe6UwJLO7jNDh75Vyxdt3WC4sMuBcnO
IvuRkSeXfb4MQLu39PiIDuS8SzvzJS0Cl6viSxZeDO3dioaqKi6nHB93uiyhHUeJKKffYQQBMkpw
HK3OQXgfHH5xH9TbrYrzLP6mEbmITlKqYSXuWBLlQXHxGmLvAj0bS0q9m1krVeWxViNSrjf4zpGN
E+wHBytmXu9R210KwBf1iuBZDeSkZ4UWcrdBH4MnvgpBcQgK29CHpwUPKEXS9XMCHfvb3TJGbYPD
th9cdTcpIX4mGuG5pl2c6rELa+Wndy2X7XF5JEs1JoVC8jzoDWg9qoZwgiMcTzYBuPiGri+uiKEi
ki54JF+v/qdC5K4AtYyb6Y7PK59csyFrG2tbRpb7s5aG2SoDTrPvdV1dfLoBaSAS6Jv+qZedyjzy
6wfXh104STvqarcPmaW7Dz+0Up3VCXhsWb0vRbe2AhTcB92MHVOnpeIkm2AVjT+Y6KlLIQx88JcG
iHOxnpuqNEx2oXhgZvZZyHwajh+w2XLTpPdbT9zA7moF83Pd6e4IYm1rBVb57ci9DiC8kOITyJ5i
/Q1WEfPUvZto1T6qsMA5Hivq2mouvca9USUuipYEKFTgjnMr23c+frQPxVJcNnZXraPfaj5g7lT/
BhfZkyF2eXlImy1zj4iWtLOnrp3jB0KnpI3Ga7if+AC5UukbeQAPZhkQbJD534tb8IIPGjG5n/gt
S2y4/ecYuodoYlchRPPF32yImj0jVCKMx7DAK8TEFLSug3l6IwZp2K2m6EM9J4efist4fZhkpTZN
k+bm6dwC7+eXHuFqCdMHm4VcZEJIOuSCK21zffAQxAMf4DJj2x6yKiNDBizAsKXEM5AvbhZQwxCX
B30/mTUISw4QWw7YOYLKIWARtoq7vN0hUzrDwTcarAZXrdC9MlNrSLeSF97ufTNFVoUCFZQ3a6K6
bg0ufbiSrV0z01kQxyBxlGHjHiFmUI/mlk4a2gbIMKEKs/6DS0YT74O40sJT1qls8h5hWfKLEg4Q
W96IXnGNqwpYgYff4k3ALygMQWzSCvPQDEGRN0HYLkYEJrsCxbryOzE/mO8CKLUekHfXALfQ7waA
V7Tl1BnsmVuTA0Rs715k6q5tC/nI/WobwgtzByB5AF5ATLH3ded2dbZrwU4gvODP9RYWDdy+y+mM
yLQ9vWMIMUyEnYVXp+nH2imeAycBIhSUHfsgISd5/QgrDPgvoAd2dg4IAEXvd2XC2OTpOlrFWFI7
TDuLyXSj9PhPiQEKD2UX6h07KEO4PHe2PfBZYgfK/RVNYobsUaOHseWLNI0yCjAb/H91MzNtlwKX
T9QeZGDPA+Smlxtuw7gAFYw3PoKj1C65cLBbqc80S1GHZ5QARjsn1HzOTo5rpBhSVoUyRylialP5
nIqSQcoT8BP0mXMWXmKNPphA1suWjV2iSjgSzb5DqmJsEDzUvX7ADBeY5yulAyj2Gqi8U84QvAzL
YnnlXx0l/wQXCjARjJ+M/O0Bd09hVCYz40B9f6sMtBcZ4Tqo7yUiP5Q8oGymkl+vtuu6K8k7F/YA
2/1Pod23i4jM0mTho+FmhoQOKXKT+lyP9q8y0LDH/hHXljuuf2RgTcRWBbJNhMpqjIFQYaYCqPnq
3bq+lDKqSyxBBoftqAQBYE/VsxVtMB5KyL2Jh54JqP2z0X7uyoBeLzCy4UtxeaKD4ARf5d4RZe6c
81ceFrUqCpAtnI0nOJC44I9o5gfgQhKkaqBYqAwjwwF/HrhaVpleyqb7Z48a6MlfPbPOZaI249Oz
DEt0NotMw9acmwXXruWwykrGV46NCCn7zEFR5vGnXiAaYZfXPSmRzUkcbo8ukpXOG0sRHr60LFR5
4gNjRmeLVZ60qFoEAZM80S60MtIeM6pvOGPkez/n9ESeEvuZwh/Au2glAgB1Areyq3k2cnfR1CV9
cvupETBPPc9lUl7fIrgsM0RzB1P2g3+AdGcbcoAnbvRC1Y04OkP077ON+ZcrTi9U0e8TO4yGQPU8
dmHxQtkuc30yNFrqv9Fd6xc8pSsODsDOkmoJiEjk16nGQDt9IuZ7YXu0M39tkuS85rvAzvX+l2BC
0wid7vyL7L7wc3El89mup5ahzNe/gBbTBEmo3XQ6jE7t76MSCDgHZzzHOCDEqjgjR3I1zeivcWAu
+PohG1G4rR46d24SLoOYX8sOpECKBpJaKLReTk1mV/2rstIrhnr1Tmer3OeMl5Wmr9+CD3vUjtMG
sPxdxZS3NlkSMGGQICP53qPBjdc3x/LkwD7ppJUCso8WRDgPGZoLONO2goE3UL0/6zmsUmDFApoe
iW7KVpaKEYIQyW1Vj2xEmHupY6T4lmgiUB0+enD7Llro4yA/Kv5QK5yJYlycbewlv2DUhqLrR1jX
FhX3s0MASKYSJ4h1AgfIpZmP+p4+ltd8UZGTtTVl4FQahFUyApEdL22lCB/n36K0/f6kIm2z/S8t
KD3wLi5FAHXNxMknRLlCQ38zAAC9CD9cDY8rnnFNW/a62zu0Z5mNf3ot+nZxPEuxxuy3OCtUkFVU
XbrECEMOkIYzpQDQXO1pJOFGQIQPUrney6CeAjUVx3lvWIuRFQB/OpGKIBQ7b8zKvDWNQnu7hLoi
OeHJtCvdEO554tHsGC/MVPtEGV+KjWhpNP6UdDVj5zYP2r6IvPduXtw77ZSefPJ6uD6F7N00DRuj
N/Z5bAwKX/KwpDweuFlNTTU244VAxido4DkF9PKd4EcY2L+KBViRo8dOfv/E0ZnIc9pu8wfORHAr
1x12QQ52KrReLywWREFdBqwvThTFJJdfqg1w0GmUGY0vikmkVbsxENGTTt3phxN1U2MeK4jgjJyz
taePPTDBjudgvnG50IP6GHNp0TzdM4DtvXEnqX6uctCuObEQKEXSRJiSOxXT0zbC4CmhJVsRb9bm
XV2BGykkJm7qagExdWCoUU7oatCmsuKuhNKeMHwSVTeIz/m0qQNDVtUDJu1CysWJscLHrni5hD6S
6QOtYRuro16um0Ylz3otU6vgZ5Giv+LQYAHGvrrx7yDOwIGrcksvlF4iF9shHkpEt27wviEWLATO
ARPL3z/ij+VE2hdS0Y6uHzHPoqbNE3AEaibf967hwCfP/+6swXyebzYjwcW795V9NK/uSuPZmRI0
NdMt1EjVIUFS3gtlj5svaox8jHiEmIMUJJgWZS9yhrszV0VOnESTDtgHYgDfh7kMqQKx2KtfYgSq
KhczXQ8ZjF2rs2Uy3cKcG8+5pe6rvzE77K27S4t1v9XxXfy6zkUVjToVIes4zra0ruhNT90nJrDa
BGTaBIuWDSAPS4Olq79FUHKL+V5zfdsuFo1Vi6yV84QTivhfLDKQUa+cO2UZ4QvQ4OuromVC7YTs
QIa4c3DYkBLeM4OPCzLttHh4sOTkr/g8QE47SGw7B2YIHtfpLtaYSENK3zB379JfA4O0KaXpRR8z
KnRoocavQCVkT286cSu7fomvwbJdGlE0uS0BsRajlCRT27rrw3kRgU/ROs6OAiSqxefkMTtlE6SQ
QyuJDMaPH+lA1QLYjvUw6zDD4SHOiJESDXEgnhY2TziN09PBe7M83dPe4h5QoRXJiA1lAojxQVoc
I1rYNz+UEZ0NRqL91LXXP9j+H8stFnlZAQS/T1SkHOO4eFQ0AaSbItHTJ+PltlLST/istox1kCkd
BZBy3ms/VmZ47OVeCOX8Gfp1DsaDrbosw8eZs0e8DyQxfiPd0q0a+LjGywiaqKRVfam3rINNsVtQ
a4OLvxHPOJadRA/22+4h8HzyLgUObD2QDkAtdpOtZS8GN2Fau2dhsUEltdB195EqqfCjAcvNon3N
zr4WcXu3+eLPw50Pi9otam1O/JTrBEL6cLl7vDvQ+QEtu03VvuQjpHS+MfvKhHdkJPoZ8PZxx8rG
CHW3qdtrEHI2pOCxUpXs5dVOm00iRfym4e2OlUzuLbDruxVQY5TSjhwWi8YNOFcx4hPF7NMVg74o
Z/XAMALe5uefdSq+CtEAVxgNfx5Xv8/KJds8BOteOoEbNmvBTvDYIXcMvVgv3Q0DW6XJxFZK2I2T
/3XvkTCifxKJ8/zRDlbAeoqkuaWtbUs98NijyAL1/DbcYxJOmxC0HmVpClJasRc9OtbQzQFKEz/j
hXbzOtRJRX8kJ67iK9bUsjegxjYR6ufVXgH3YmTItSGysKib903Hy6FGK/FsKbsIKFvziCQatUMl
mtkq2jBhksy6cTYlEqBEEHu557z2cfPpbvVitIMKf9+YynXznFz01Il9T4Pg7sqG882n4gq0qXyb
1mE2aEB0R7IPz/HW+jWq9MGo8NvcAtZbX3hG4VvXHzRRaeQrjnhymbShAxjeuWzleJ3OGxqlUa4g
Cdw6iQ2dxoXtAwGnymk0P2XyKqSaKQTAwZbzDx3swUB9jjhuzQrtI3esocPLz7Cx9MVu3RrDUKQJ
GI3jYpo5Qa/Pw7ijCGkyy5nhuf/TINTy4K3WMpnHWzTT3DE2N57JwGiBTICs2NyDPb9HocLmrtk3
6G9wPcukzo7rg+cPeJ/n5baZTeqaSHP8s4K3J405wuqsnrnGLsVWDnHmvnZUzo2BuCVXkneYztmR
b1OdkgvuG2KmjBZU4PChJxBViiC4DQeBmcOYlBnjK1OZcM3tgYR7pbsJLvmnnUVp06shSOuYi2gv
SwfFYWUZk49bd9iTzySpSM695k6R9IByDdOOXpv+htWYDCYRC6JlAKCKG8zS5vUcs++ZMHuvZDKL
vzRot1+Vd1PnNKWacA8dKex7VrCPNB/1paN1A+Dz8Q9FcmyQ5wSUQJNTwyUgt2KJP9JHEh6gzk8d
QUZDUI4zH53jiJAv17YcIq/lIb7ztBRbFAauGwkeO5qVwYZ+GtTnSi6aMcczuTPxyhgeVjfjhg/y
DtgufO/RUzC/Xd2bPeh/wZMGAy8Xejpv9vbXwEGv3rELW789n5XogfKn4mq2YXvAu2Bwz+CGlqXZ
iLTF5hE8fLHDMFY19pdqcpA5UpmP71gtzVw4rmksHOP3X9oY6KGwTueo3Rq/rQJAO7N77nrkv7rz
0w2E7/RSo09KBR9qKJUO993PI1lPrgpcMAiOseRBekFeeFobRmg/GVCzg2kOPxoPw6d5uBB4xSA/
XcgAM5JGp0M13dtLC7a/aS8tMPXp9bXqDrqZ0f0cZBtOmifhK7Nb04223kUm3YlGlrYJ6C0i8B5w
y1V20dt5D8zBi23U0t8bZVSgnmPhu5zpLrzK5ANMNU+XowhjM9MX0jmyLXT2uDnyhLOdXELeJuVI
OyMvQXJf07FYcAzoGL18wygCP0GDn6A7Ec4CnRFA+LRoZ+CulGmOA6g1J72cQKJaIuH3ofVDkoRu
13DJKpjezink+9g0ItArtXAuwa2Dae+cWNaHeobYpVH5+9NwBPrKtbOwtvFhQWmMDdKtch73Sgs4
2mp4hyIaUuexpb0S/CCdIywzutunFZgWf2FaRcfefxEuyXKwRYrNrWieUHDQ28jacZW1Oi+OfN2s
7iO9EP5kMe/SweIRdHGd4owaKJlWQISn/ZtYhpGlHNxfw8oyHSxUgW5/0ItWB4Uty2T3Aa0VGXIF
aRAwnB4dQZcs8r7AZVlftjPchRfN3sffXSi1OHVa8kN/gMM3WFy18MKLKD28mcbd4PqNFHZ+lK83
BzWb5B7p32IBM7BALX/tO5vuHbwNVzq2CdOfFNcZrrkniDbqBiLtjzunAfDYk4Bin0WhmmG48Ozj
u+4eKL0KPAE2gj//WYly+TZOchmgqRGYJkxdYjKr8d4FVJxAieYbJ8pbTKnodw2xIDg7JBwdhlgk
aOyAXRHKFW1s16xohCxRKcSwN0S5xg8TwRVc+IpfYwKo59eazGvZeffbEXnrRu+gjb9IxzZrMw3y
Ow9/MlhZpJfrOrWQOve4p7OLgSPp7tyn01uDnV6P6hm5SsaiZFgubT4TVbDAeoEfrsfenvXBbbHK
QHEVFkRDZ4Ho57iUz+hTW327DmGvgb8OeDkJ/da34/s5ghzvtoWJGIpW9Y88i48j5bXWcu3Q1p4U
lvqfetD/VaIb7QQHvsNkpwRyhp1DPtdOTUp/Ssf+EhCQ++vPsg/XbM2DoGKeVgUr+jnI5GTze+fD
cXvBpygeSlmZYkNiXWoyfZKvstpZ6qchaqQPFJ30fiacMtsxX9ZvHhsXH6Q8DdNjV1dNZt+OeXId
Zfh0iw90O7D+OW/7p5+H8ygyP0SvM5wf3J4V1eJFk+7c1DpZkm0rJMxRlXs7U9LeVx88gI3Pen+v
EQBzwQgaJhHCDAT6TTg+b5x6rgL606emjWCBOfVtvNOXU0j3eeRLncD7xT3xbp24rwNylclF9LjS
1kYBbJoP7Wicfy+lRI3jhZQJOfOq0eU7Rcu/SZOkRpI0tl83NFirXX6kQgWi/amddQrf/VObfcyZ
HYOtQoRPrmT6NUoKxLjYeL0pe8kFCn/pTeDYT2uq+cXrepwTmN0IVwtums83TXx6Y2G7KtJZx608
qwmnKNhJFbYhZS1hQJ8V8qNtAn+tTceLiWvHsdMcN1sBl81aXbJ8HvCN9zrNRWoy2caDWjlzZOZf
ON0oHs99C5YgB1I1lD/rtC8/S+gvPO/S26rUrhUDw+WaMGNwZTaM+n1oRtdGmtQQ4dqoBUXb2Uhq
Fk0mtCwnJHTu57RYyNSsBrUKy9HFxmuEIefDiICA8sAeJnSBv1a6pkMEx2oQAfjJeEZwPi1V3pKE
NOAXJCqybuGJWJTS5daEeXIIOacvkNqoo9YCAEpNrMXIYXOqm3o5S0FX8RbMRG8kDFTBLIzife4V
76HjQtP9IXtX5upx07SBS+OOHqHr9sckv/hEyesJQ+UlrG+5YKIVPBFMYXwP+IzGVIjdWEeoakg/
58sAJdwPcom4VNP21xYgnlxHuS2UcWIQeVpdpqkPl8Ff3AdApVbnNtD+DrcUEgk6Ia0G6Xzm5w3/
DT/LONhJeoWnjAfrHaUSrQYpPC5gzXt3gwrHbP2GvWkLP1QJV6pErQ6TpVpeNuzGuv5KERpQmSDx
3CFjLYLA3WDQ9GlWde0ZgkKsE3BjoeutOBCETfOIXB5U9QjHXtukZqtp1euw1NYz1lNN8OL+KLND
47HdZiMkNUNNtpYdsLJ/1gRjJaPsKwR+jhZEBChNJ+4z28H9ioOZldBgBOMhSMLbYPdjR+SuqQa+
msywbRpVCfERdGnAluwcMmqbEwoSOUph1GHVpJGB4zDIqh0yZyAzatOeQr94I9rxYbJE0O1mBe7p
1IJLWQFrNVdO53uSUrHce/D5sV79tH1oQyMGNe4HfUQrUCDWE9zPIlNpWrRLGyrbU9ITIKLaIKnZ
u1+dy/rirehSfIgZwLWINksiqRNn2fj6glfjhYYcH74TemLYO79csR0CYa2dRDgY4sfNFqwQY7cx
Ca/YPZFYLHMJmPX4jr1Et7HyYvmVbtzkEjwf+/Gpantm8cJn9c/r5f753VrS+f5e29FulrWX/nNI
Ybk74eG6QSPp2NMQXCUgwUwvR3ygyUboIynK8mAmKhbdV5dR0IAoHv9rTrjA4Edl0DShn4bTSmJZ
xel1kJrMqyBOn/kuwE0ZIl7svgjr4HTfejxCe0k1CCyZFXbBbhjqGFpkdgJ5fbSGzxU3F8BqJRII
hZDcB8faswSPeWQOCgSBxtg2V0qHnEG7ZoOr2nO4oqxC3UA22GkF5tigdmh9yEGQ5Pab7O5X4vKE
st0kZ2ZI24w83Fs5FdVBlMX+hVGIF3mr2AymVW2qni1aOpVmiGxSmzzGftMpB3y+rfXzR9phvYZs
iviWSIfjFcCpAkW/z+pxbgd3mGqeLch8M7HUFCX4uVUTPgg0X4LxLJqWt+wyFUhnDckSAsKvAIrS
4QeKFp6ODTmpg0zuPwohJMc2d/XgAy97KaF9xcOCAM6TmeMgnEIg2Zb7TEHxIS0ufLkZI77YtNYY
+ECLtSW28E0/C2nAA/pQ4Tj0c8ZZo8TnYlX9G1HfhVzzVudJ89+U/b33/pZXEF4f6RK2T+YeIbOM
HFSsjR3XSx3R9CKCxTMluVFvTYMWYijFtSyKM81772NfQIg7XAmZDYGi5V465Ke8D3npXb4Cisvk
0PDxc3T2d5eWHdmYECCrMiPhq4fw5bOWtmMQWYCcpTrR0lfnYXq1WiysjX/S+Qm8eqYEuFEmqFTz
9N3902o3WoVyIDYnxwzW6uXnLRk23Z4S4dvWbRwg2Sn2GmlbEb2q2FcSZjcN4tfchyx56nD2Xdk3
6nR3af88bqCB9ZJ4QLWhSNQRx7+Kl1PIkb3GSU62iZmpI/vGYqqpuqEpjrr5DlWjcIuOaSfDq9CX
r+AI/xclflaKcuqDdFSxirOqBT6MgizaGqAvj4acqK5IRT4Qiai3GKRtVfa1cJJqHLJhnbuGFnYi
2tvolEEamWo1/km6ewdMd6WVOMwpU1vkQBgazQ+EWA8MVRSqMQQnBsSo3Vsq+6VxZbm9O5Rt5i7H
cYQr8wPXNrrN0E01yb113mP6mnQdDdIHOtXrG0fbBTXJjMR9mhjpH9Ysna8VVCdmcALxhnsbXykz
sOSRa4fjRU7xuXhIvvciDoohwBIrI2BZmokbezAUvKc0Hu/5w1vCvxag5/RJbw0SLlutRMHdzDUf
xb+wKpk9XPEiFNEr2G3tOFGQdsfFgbg5nmZL8Xivs4vMyZf83GDmKIpSeBHLt8nqUiLWRmxN0xid
+xr8jE3AMSeyDEzi2F11e72KlXn8gf9BxIYw+nqbhDRzrupzER5V/GZ9TjLwul/OtiTjx4J1H3G1
5NeuTiNuGM6xIz86MhlK4tzKs+n4asZTUqhJF+bUIWofncYb2PtJODGnIW2C3lQFc7DX3KFLTAGN
95JuSHx2aqnhi9QS9aC156hVAivAD4IUOeaEZFUtyImzrYupC6cpWUWnwbMw3DH5RcyLo2bv4QK5
bl30xS4nD32VMoRwZsxTZDWpfGGY36XdOvuTCFdXTN+M2WmGZwqVWfWyrNHTJtctxMQtWk/Jy4VX
vXebibjqi4XKZSIvpLGRwKYPejd+AWXQg5iWiFLqiJ94nXoHhf6MBQ/kS40UTsA4NAxdbspF6aBQ
z1gUnWGIC5PbzgKUPlXhwzHTPjmdYTB2vpG5gT0chx5o8mx6O1lBSm7BM3uN+sqvCA1qLLF7HCPN
wNYGoO/uMpdTkMjLX85gAxLoL5f2JZi8f9wM6qMvgim5hor1nGBdhQRrqQbswCCZCTlOmUBt6QC8
bZrpyKcmFaaVOwcShrsvaKCLii/Zv8zW28kRDrMtfxO5lhPmueqUI1fz92P0mudqMSSOKYEHODXK
LFuW6CyYyhPTDRrqMF5fdzEuFbjVCNcbjgfp+PzgBZF+phkdR3BmzwfdT0VrYCue2IQoLcA0NEcg
UCiCdw8aUDZuneFpU5vahCsA78Ed0q5q6x4RFiqqUdh4FNsYxiHo8FbpgA+mdXbxCE/c1ISuT+xH
jVE67+rNxP3Kb0xV6lFis9ocWExNt+RHH30a0Ok3IPsv7NVeuyQ16mHIW9gMn1y7G596m2c/Xznn
UONLleriRZSfEhAPmp2OxudM0SlLtkfwd/QlslNsy+jw2yXVWIDdwVF9MkLKtdvGeUjZcIXmCodZ
U/lCWDj6AfNX+CLcNbTQxAJU03/91iTG2YQP+PN/f669MfcJIapnODelj3cC+tsm6yMzf3U3seoO
Ksg4uStkIDIuAeHQUlRp0+yFwtI6BM+3+/GCNuxwwBb/rXK/wCIIKhq7cPxasE4fOrZzSoCPVNDs
jVe5qXVRjSSULi8PtvRDZZlQN7bTKJt14NAsOqurLpfdUeW7KolmyUyZ69EGRetU7BfmreyM7Nqo
6JZWdQCRj+hSQ1zVAlkvhuk7VDlE9okEQ3EYU67IPb0Kqefwy8IaZ6MD+4CqvccwIDDmAkhZa5Ui
/z5c/cJ58Zgb4+MY68FDt/M+r73rT5HjPQ/4I+JbpsncyET91DlY1YHFzoDNsYlCST/a0dFkVUOd
WmMig7wyIOrwF15oYdPZB0/h2y1OlMgHAoTTXjSSUGMsBztpNs2qL3KI5Y02KxJfszhb/sSPZFzZ
ml839BAhWwJP/9LgLWNPhHHyOJU5tgbhTEad5bMinDddxS9j6vJLscwZi85D1FZo86K+NTtctXnz
cc0ymCB5hOwxomZtD7Yg0bQv7YSPlr8jLebycPKEk0RmWpcKNY4y5quY5gSACy6OBERoTtHRyC3T
sDAHFKG+IyPKy3nsPCIvJBpmx/Hc8u1RGU6VzAzjP+N/QjfNtt39d6mdOeikhlOjOobDnn/8SnEU
lVD9Le1/dq3r1IDnszlGDeMKB2LiS2uDnXeTKgPsLmduFXVXZRV9KZDQQdkelTo8+C9YlOaZsNKJ
jjd4pXe2lABTILoMTlweSubnBIxIWTchinV/MKlc6wYP3YYf5rYTQBtK90z2LB5YNsJOu7JvTv27
LcDFyJRX9KvGdy5Nfju7MTTLTpIbAXidnTPBe2loO3+aII2YXBb8t2qVN6SUY9A2SxkNTFKbBubB
G80ZKYHStDKM+QY1dIIeeL2TPOqDZPEaxoa0RTJIpA7/0v6QqVzLrFg/Rr1og1C8E+99C0gxKSvN
XwlCNvFhfxDrYjAbvfpQRS+GsrIcRoIwRPvjAhoNa7cklyF4H1e1ug6Se5mvEVyTFTKFMkx74wKx
0zHB5v/dne5B3CgCgdM52/7K7I6yLAdsxxfbsNqJrlrsuLakK2vUD/OY5Ypgtz5TpZCOuZAiTAVL
eXmu+gmQ0V5/E5fEjl4JKej6Tf8aUHGbPFUPROw8Hxp9ETeJh3YNP0F/Qb1ryaUUAoOhk2qTWqz4
UC2sLqcoY1lQ0NRv5zWNf34G6xilQ5wjR7Wj6T2ADiGT/qKYxHs5uOFHHAn2i6brl2uSUc0gN4DE
4svxYL70HoR1ax8DE4RVt9+ewb7+Snmc8Nl8Ynyaq9JYF9Ay9HAx+SnfMsW6KJFy083oQjyxp8e2
5IGHLYe26DOg0KO9Hpnpah7UPL8cIXcV4HTnUKIhI4rvMfvG7W/3U66aTrjcSdfZEPfWRs4iBBwS
YJ/q8SrOd9vDc2HKiazkRtT58wcfhi1R434OuZ0Horw6SHXogOwjdedPYbyz9BxGk8VhcR8yl3Mi
O121nRK78HLwZtFlqK9Qe1xjD4LbvV1ypk+9h/rd4GFMZTCsy1Sr9sTRgJW64WQqPxFu25aCopsZ
6PzILMzWgBs5k0ayW2Lp9XCozhdidvdChTyvrGQAUERmC6r4PUsSCsxUP3KK3mbF+IE73IeOABcD
origdCBKeirKbvQo0kdEWxbclD7Et7e4ZtrSrFVsXLKVbj56yn9tHoO6u6UzhUceFMdLhEk5213d
BIDUFoY/oByCthtkUKpbikbwpkvd3o+/rH5PebUwALnn9m2EJ6TYoHZx96uS/atqbwuGkxwS7KJz
70ZnzLT6JjkdMv1bwyxR0N/P4eXj6qzVOWhs1O17EEe1wwhjGZybHydlHJoYOb7UeoIihAcRgxi5
xratLwKwwHojaWsMWKRHaL5XuNaNXR7pi1clA+l9j3dawVTakVWQj/1ssqY+HlinGKOIhzNS0PHo
t6HaG+y1xh3qtJDBBzf5hDaaH3HPu1CSPuIVYEPn6nrCEjL6U8FiDeocQNxmTh9cz0jSeW3fitlS
D7WgDzV2+TMNgkuLKriakwlUtCujLxhjDY0tlTX9DrRyiSj5T/syzymFqV+HpzjxqSHfAQMeuft8
rwcFiRcO1ZaP2AmWY6pYRCNoVr7UX4vRfWILTVZbqATVYJIhO+ZbnlJ8AaNmG6KnlzG4+s6uSsW0
Td4LHblaajvRHYOHxdPsVNmzaNZ7XJKFq1khmVSHIshYii086VCqLv7A0Iywp1CK6Vm1PouABzNF
Qpn8evw3C5XZLIoYgvYCUSPF3xRxOz5vOMiPAadL+kJcZxGj1yfCOrXtjbxuqV31VImequpsdpv2
Rc56hoUVd3oOee0ZaJ2XlFSavW0lMzTJd4H+o5VLnwP8IYBsddIfCfT+jryAu7go9Ac4XvKDtU4A
biekIc2vmVZ0XbxsR9Obdot5traEvU33zLWUJdjp4mgWfLHYLTgcY7JodNnNGZokYYnfTukemjS+
CKD47kAC6Kqt0kJh4zD1dIgnv3kZQfS/E6hjfaRqQytxbWsccLVlYubtSlZXgR5rhVt3yCPrOiUK
mLZr39Z2x7MpcZl73qcj0GuzxIrcnkVWk8lHKZ1sJ5WktiEcXE1HWpzriRtQc6RGK6OcxHMf2Poy
K7n4k5EEpBrSlHc80nViQ2bndORf86Ll41tbtcx1JYhjWGU4joXdCtCZCCvSdQiJ8+U+1p9SFGF5
sTIQXAmpnz594ypvXduVx7Ds7Ec0cBnGxd0siyMTfNK/9EiIwoPBSIklyua7BweYcav5TrL4/eoC
kC4XSTcMreK1Vt3XCotEqHKO6oV4sl4CfSTXDiJywJkn445u558w0KeVIWpcJwJ7STeoTmr8SQau
20gr+6z3MG3QZLG+8jz9wjkXPO7Dt17VW7Gf2BQbmFqh0bAVEKvkSi0u6VWAd2pMPs9MtnE40AH9
8XmGPk6SwAN5b5Pf1kUGrOrzU0GjPf1aCVZq1Dvi9608vlM/ymeLs+9jeMkzZ+q0B9FaQ9iVO79l
TcXByt0vFmlc1vJqppfPlpAi807oWTqLXARtn4FcMxdvCjQ637UaAqTvhoLjO/oQdE6AIss5IUq1
jQnHQT2MES3GGbL1/Dkjl6nVrCPIqC6G7LIpSymzUEkNIKZXz697pTVhC90eOtRnomWGQ+XrNmGh
BMFyPPTGUGz7l4OT39tcIjrmK3GW5Dhc/gjrfpmna+Ed45IqB/t8wdw5+PMJqNHvrlAR3qc4E/tv
BuEzZ5Oh8ATbYu7Pp2NkA8XMuo3jaDbCtqShiLcVxIdYAJOalu+YcwtUw3ALoZbTnV9/GpKN+rVB
VgyluHtwMqRx8zjyMdIuoSVKSw3siE4RncT67apSLt6QFJ4m3k7kZzwf7IrLKHJAFicjytlwOA/c
s+lisR1KwthyJgTnlN2TbNHWjMDOGqywZOPfMgO3mpw1wk9v//Z/evP/eZ8R7jCzZ6jwMUnJhTsU
kn3+FjHm90EUC9rV0JlAKaKiEjQA2C2wWcZMOrJj1vD/rfNODsNeAaZQ576YB9Tvsp32uRg7ZhmY
OlahjsF1CuZ8yxK2u1FvnxSpBpu9YVFjhZsAN7huBCnNy8MCXd7XR5mpSAv01r+afRLevgz6+tcy
nz6io2AhW6torQpnltT/Xk9yhK0Z2sW/8u+W73S2QoHzxT9Lm9nDVmXrAK3GDFPVfNbIfXIjN7a5
cROgizXEWN4/4YP/5TMgQNF1fNS3lWkdN0HSU5wJ3Z7m1FasMxnMfoH4J+94T1zMdcSXRsrILkRj
YHvhLG/DHQkn47W9ixCZCZcQmYMwJBaSszD11mbZAg+KvaivNi05hFmEGLSXWWVjwGDIxlCSCjgf
krwm8Q1+jmHl6cbsyTb6dR5arIOPPANoCu8pDMz7oBg2jNzclauJ5AztZBalqlcLZe/8p+gbbZaf
LxRt9mi5zi9NSEKrrPdZycHhpeLAtkcts0Pojupu7J5jrwSYZoWKysrBVrN2/ALqQt+HZO8ihIBE
efX28PBrMdxUmjeG/n5BBKQeY3oQDThchw5/NIWwpR4i2CIQnyRVlIAnBb/70iKWhmfw1vYVhlJh
UEHW0d1Tl1LP4qogguNdZiuqPcMOkT68TyIgNecCp/XYAoLliSSAhX3JbP1YqJL7fCdCVctrzHAh
4tWHSW9OinXMJWpRjH+Nn9aB35Z8hp62I6+8yxh0FI6ddaE5Lb0StAeowp6SyXkNAL1an7SQjh92
OTFqFwTZ6og3gjVOKhap3lC1r3EahtPoDZQVy/Zr0n5oQkTXlQzAIYWmN2xXvZzam4eSP2GXQiol
IUsq9P4AvBDzmFZwT02yLjP18k/Zxg5x92QDlftzFXsWNQaOxIi9thF3hXmmo/pG/Zra+70Zsvba
u8Ip+/ryR0EkFJ1m7zbAqt2MqVNnj/ILc1yWT1fdB8nYu8WtQ3ghg7pzLfaOUhXBHEw+h0kAQGFU
Rw699S/GA/05mqSY3gQuFI+R3q+MvrU2DzJRnUDRrnHQpDr5OiTgCY/IyWLgjZSadnDYLdMmVOii
CzOa2u3kNDp+RnWQIiTPAXn+V6Wpw8hvXlR9zINKGa917LUBRi1B7ob3eqCBVkyTRWbbACrj7ujh
ndvNODAxZu50o0AgjWduWYXSgugB+O5Tik9DlzDwiqRVD0VwE/y3Q7YLDZ5urdJM8bJUoWITu7Ca
jz+NVwHaVqSOqRqpF8/SivLfA4JwhGX0FPkHTGqUjWBmnsqObvqzIlafqmMw1pyO/2GUuznzavRh
tiEfL39WJcm8w8IVq+KfRLLzbmGlKyRTIUNN0d6eTzhzQvxtK/drbIwpe72w4p64O4tsgPva2y9V
Vn8xvlDPFiX9foEhQFCqN5kQyWFGiaJ1QGT8YaeGVjcZe6VS/j/tQm29sFiFrcUggi6laeVRjosE
s1elrtS++XI1RUa4ekiCb/xU6JslTbrgaxjtFtCowYMBOVzP1YWPqvK1Pldd0gS6Bu98z9Ny2xRX
udYzPteNDSi3X8eCvzVwG0YZBO3K2ZFsTNfCbkqH2ijOR/Bqv3AkDsZzZ08U4MH2Hu2mqIvPmJBg
zlgwV5VCwH5gAkRCz7eknnllWjcnbcpZ8hsuRHc/GE/wplO+nFdByc6kQmtEWxggymyHPbFUADnv
FX5wPCkifVyb7MGTb3EpgfhNAvxINZAkJ2x6wyUYhLoD853MiNsbLPxorO/MJ48u1BfclZ9OEBRZ
FEbTcCSHORbh6YLNzVlwP8/2OCzkKdf7BtK4Gy1otLO5TF7dGXHWzUn/7967u7LcDVqEpEt+OMWY
fXJrzPSK6AS9zpxXtCVLZsqJO3ifyCfGOgOzPsUZ/5+VZl3FqLNHRhP5drapSVz7UpvLm26iXHfq
+hIrPP2IKs15Emwem8/blmDxxnyI4fx/YQQ5rEBoiSLZTpVgmFqc1ZFyHvlD+MjiaJ5ecmrxfv5H
4ep5is+CfB6XT+TlKr0DUy8LJDXoqrSLmMZe1Lk7wJ//kGsWQxrK4E69EhWVI9lWg67QOV0OOA8N
/g2F4hN22EBysErijaZGvjr0CoUf4N9Cm8IDaXJ0KBBcq2EN01KzuySbp+jAzDYF6MRKBEk/e1XT
p22s7Azi0HkGHKd7sl3a8HfHiH1bdkpA/V9jiyFoUXUrjTZU/JEckjToWn1tdMQ/kCvcqjK/6FVk
st79csWXC8+X4LPjTsih1Hhjukq90gKhLWWzRR2yXu30pieR+9gf7VcezbGYy/I0Kk4ylayoeaj7
L38VnNkcUO09ai3+Ut9WUmmgq7/9ouqtFFRjJYNz+QPXXsOteCtW4CwJgrDsnHhKoabshNA3cR+8
rLHhewCz0w6Ygn1Ww6DTl2SxPLygThYit8PtvN+TQJJs718LvJXMYEezCJl80asNqU96wq3dlwan
uhxHf6QAhL+hMdB669SRDQoO/rDOQP7Z74rjkJcuxs/JeIoor6J6m/pPjFhFfewKKvNLDRpc66ce
hjxbcIMO8frG8PgOnHwVk5npWw3nK4cCsXHXIAbag8LCvHjFmLg5XXe7HRZ541Z9LMcnqftLCKU8
UavVN6hZutoabsYRSGUpjUq/YT0JyifYQcSufL9S004QN2uS3u85ujiPXp6HY2At9StMPMDfpP6G
6GqoFStmq/Xeuf1AGe1SOyoX6R8snACd4hxoWR09kUaCg8h8CsuIw0crMPPCN+TiSZbygLxewJSZ
IjkfpN5den8zPq++MovNCTsnp8E4amzkTFM0Kw8zAvxS5TzEHcISCLb3s1UWxz0FGejk+Ew1knbx
uzrdu85H+1jMp7Olu6aFdU6YW/inTOoXPHYpG13ypCON0X6A3WlPC4ljA7foNzBUiOLvDYg9BqAt
wk02EMv2MwMRTNkU4zfH63zjgQTO241XqjYDGfdnjYl3vpHtko3omBjgrpYfA+ETxaTbhz7dotKv
Yp76Z+Wq55QBGzRPuA1Mgr4/F6gIScByJIb0TBdTego/pWd8427+l8Y4/S6/vJayHcZaOMtXD/9y
srDb6XDkDXuXow1K+11EJE0HOOVCTv56r9AO5AWyDjN6Re6HuwW0jHtfgaYCcxaPN4JOU/JDVctC
dR+X/4rPKBcExQm5F8uH3+WBhPsIlb+9kYvObrJZecO+/+kZZ5f+D4os6SgN0Ti1REr/a4bepjlH
wNkX5MpPnc3vfAHCLaKWXTn4+OPg2/O1MniXHW7xLUJWpTGK3YjgqoXwO/+OaYQ0WjURF1ZDEaFu
rUaU+lidTD7J7julAGa79ZZ7wmwFNayJViCoIlpTrkiHWF8xZiDMJwE2u0v0iTI6DFcI4AfTWspc
eC+mWUmWfL5FxzihgkDGAZ8WKWn/7RCc50qhOGw/7MemA478QaMzJEA6bR0PhB9QmEFltnZ/UQB0
6aGqD3PTPGPUN12ERmKdXWNhEbMBWlY2DLdJU5LBFm2yT1eY/t09uyVu+GHB+InEp37yAD0Obwiz
rHJh/vzCg1JUUllxBc6IANydpvxAFqZDLqh/suFFqVGe+8ac1nCYVqtD484hRZqF+pL8FAgDT7HD
1juX6BKfAxC3+8LV/Zcy9ZmeDq6j3Xb/G5sUw9YrHWIEtXNqZqPJbmjMy4t6Kim6PVQK93SkRvSv
/+dY4qkTj4aikT2QrGBUcghuBIY3hxi/82g6PROMQXNxw8N3tz2Dw9k9DeP2Anwur26xcvbwAFaX
Shyb2Cr1IdLckgweCcalgezakGYv3PHWmCVRnbjoEbnNtBCgTvGrhQF5SrL8ent0GGSgNJ1UBskE
lRZ36O9IJPAMjNqCqbKwn4GexVRvyonCP33pNaa3OX2K3jD/Xo0TncE2J5SlhUdYXYn9mb4n2VHz
HStzqf+XvA5vTZsuow66I1P1sF1u5SYGaCMjPraH2YCAW+vQ/5z8yj1bbY7KX/SecPI+a4E9Phle
ABQi4m4i/Kz0eaz1ovNL6h97kFsYbNo3ihkXZDg1sRfxZQRptfoo7HJFgsAm21PAmLAGN3Own5XG
Metm0mMG6B9jcECferZvQEY5lYglwvzEtKQdFbE/DDaVZ5+ho+HzyeVGV/MwsiBqqV94+yyzQ+S4
YobjDmx96JqUCyrNAM/b6EknPDWygwsnI5xVWjy2Ov3nOPVQ+R+0y1qWSvT0u2hri935NMZk810/
t3QIZBVso/iF9rXJ/xhBp3Fuzbd9/+yiBEeQ9W74WJyjkWjlSA2QZjpnI2uFpfyzPPmoCd4nb6tU
KDqICSOrLOo2137cc3uzu7zm5lotOW558BFpbJUvvFQR/MazlS+81Y/gMcQwWbxP7lRA+Qf2XhWN
w8htOg6pcudp1QnKnKXyUUahTFbE0Yn/VsQqpybFHTf54CjygGfFC4e+SER/5NmeZjv0tMP/8XRb
QCBzFXFFLxpfe7sjTLEg+S5zFLIhxck3wYdiLEH+dBC3COMv9ZNDNl5t0eveWUlnPWRUJLml3HrS
okDQCileiUZluv9aeGXdYhZsWg+JzwzhnD7CkCS8pXFefFCKY8J5yAoaSIGSkzWJQzk/seYXf9AH
cSwpiF3gG6SEMrILzzO0LSGqr5kUbSMB5JrlGvb3Icq16oOdyTg5slFXtrfK+5q31cBH4IZHTn4C
g5YCyK80kNDlUYHkAgBQwn14lFsjtP6U+5CuiDCOMF2v9f4wbtE5eXousdR9YedXqcPBSGR/b3Zl
Xpy44uEySMM2rMpG5U+begyqI078B5qGYByP8ocS52cdco0/84a5ci+5AVquwHZdOI7lF9A7Hn0m
9zKK4ga+sG1a9QUlSsoD+dczrdmXgorDiSZUDutJz/0ORgV8CfMguuiBv2Y10aUiInzcdJqlcDlW
qKXiA8xotOg7dYz2CsdKnthfjhYZOrUHM8LBg/NMFgu/5v1HdqA06DE5Ihlxs0/jX/aXagei1Z5D
q/+sLC4hiygJHKPg4BKKeojLfPMmJznvIUuQwrVk87SL16U/oCT1rqFwfsMIS2Q89dt2Zl5uRnxk
8MZTyfqke/gcbJr19AaEG6CtQEQrVa0l7QNoRz9YtuugcH7om8BSoZ2WWpu8L1IkTQ0cxVnG476P
rmho0/WBQyCp+kSp3VuFS5pcx9MA3tQLw30v3qJYhqYnx4YHbRkODZq1wjiDdzocaABnjBc4vWpg
TBFW1KmZQFV9othAUvtdhNS1ZOfZG8UwqAMDtTJbosWqbWzd/wO/dUei8fsZEY0qyXSe2lfTf1tD
tQEiSb7jtwmWmMw2ksXyHV4A55KEYLJAfDelOXmNiOvAKGkGmmeRPsnI8U7S8LdU701haF6zloOZ
QhWiUUsnRfV0WAITm/qIrSFYdrTfNLMwRVGsI4jnvw0foHJpD0o4ZcenMickhycHzUZpFwvrTQKG
4lVJnGJJ3OSmlMQfztK5Ci5kXVz61s5Y6zpGwd7o9Nrc0Xt5HmZ/EiHdELj6aQGLs5+zTTDd74p8
kGSIfjeXGAb0C+byfYoWbAGDZy3h3OutZqxU2aPgb706VCFsNfArNt+HNknATBoSRZMqZFRcmuP2
I6M5IN4oAkGKROBFi3SosUjmzVr67JRtdyI3r4Oyjm8cfZz7xHnOHvg/uIoC15VhaXx+q696COZW
dDy7ipiPwCempyThvARM9esIEdyr9jK2GxqSC/kR6QNEnjIQlV78Bws8tJ36bUN7vUjlr8hzELme
YPzWWaRmD94A25MoObcY+dnjBkRY8h8SI8Ni5WMaHN/cBz4OBTgKWyPy3WSae6zklIougMJoSAai
go4a+9UaFUJO8qf1btiPNWw/M0uEwwGTCXXtniOY9cjWXwwtGYUiM1ME64Pfo8d2dyV0baGN1ZNw
pSiPIWb5neJ6Vsp+SCgiFU5tuJ/cqQeYT78jnBQT9OPPlgP9CcyHu0QKtVetWE4e0T0+B27rO12W
tyw6ryEzlyRRtfjhgBidw1Hka79hYrJ/Fuoicq00Dz0TaDq+v2ETw/+LVIPTZvHKVsi//S6AAFQo
v7sIuTdik7xy2QjcoAtKjH+F3bXpRHuIa9ULNHMbYS4ISjFo1QYCWzg0AP3Ji1Krty3jEFw/wV5L
7oiY76HsasXDPEv2Cpq+mxfvNcntrbFcTXXb5NlshlGAe2gNqgqGyVVL7EthpB6OsnQ3b/nslrrU
wsfSVa3NJrlm4+WBne3tlwtFN3H2zNgWOsUzVro873VRI6iecI9EH3zSqHZU7yrz2qDnwpQgXJQO
WeveAgqzrLjZW5CWZ1qo6jyoNMAvZAsZ47fnKhhaMhXGeBHdJI20/ADv+zOCdUvWroc6dUvmgAo4
klS+Cayz0GCyjWfuiy3o792qEAczpNfYt//vwYrrVm4hdErl0aNMWQluP9Q24b98uNiLUFY8XpSu
F176O3d4GFpK8BGrWVg0nILr8SP1odltekWIEi0MRxuJbMKkGIqJG6bxiwqPa18XmnUH1AurnZLt
rWUDX/OgiMc8rfJ+mjSiUgg/l6Cn2Z2G3ZgBCdKqgEF7jP3vszZdpoxbN4Q5ycHajBnCUVV9KL9q
v/cyHQSKXkdRV0dzkb//GSkVu6gfVx2XTMnqfIr1sOjLr0nPESpKj/vxtEtZnGUTh8OHxgmdsav3
27k9LgSKO8Ptp6LyuWyVzPHiXff0+ubgwCa4ve1j2UQj1jDjVOWx2UHd+9UfQKumh5zx/RmzrihN
RpB+mbBJZSTiRwh13DeOrKLrHL3NnHrZ5mvsRJVV9gPmmKyL/xyKhNvjY6dxf+7hnTvjbgayFn6P
tZjj926iOsXBWQSqGNefu3SmMbo32h8NtIuA7fRoRRiEHNy51/9gJd3JmJKfiXthVFJAB3sz2DU0
qvOhTpu58YTynHnxJHSbl0MLAi5xPxzRbvsaBTIcQypG2yxTqX5RJRdXOot4uobgNIIexJkyXXSJ
wVQK08q34548meZ5N4uw8c5P3cJ/MaNnOjb4FZ5qsohSwvEcfY1Al6oek0adkuSkSWMYP3s23hoW
wSPUDiwzbdzOUvGp+Dovsb7ujR3mOosb8Yvhy+gbKdB3YUVxK5S9+NbefJCKwE7jIfWusQhaBbSq
NUuzuEYy0gTGUZIqmLya9zk73hiCU64Tn6tzbK7rF2GPBO/Wt2/ydKqcxJ01fXHVZKLPm5uXAMYV
SjO1ucW34FptRT6HpyWK/WsfZHuCGnvGeKlxyFlZa8J0+tWxy2IJFreovdaV5+os7OeUIc5P9H0a
yX3DCpsLLjd+e/w6vCikv2jTnMJYkR32K3MfVhRvVJvkDzIMYKf+J1Dh0zKa1/lC22s3/2fMb9TW
8D4GWIy97S7yoHaqzFwZ3Vca8/iYQfmRCz4l2o9OSpvEPebM9gAVn5Q8WaInzonl3NodJUHcyy1s
8vjvdp0N2rDNnpe25opOhVk/jOgzzv1a1LDHJ7RvKpHHbc8/GRD8xv/qXwmJ0mKF2+rm3lvzTZQq
Eq534vWSs5RHGDN+D9WYtKmfNKkAlpM1kCl9MKKKnKgLcj/zhWp6F3D+gsLbY8Q0vyRe0KPNCM5j
2PISvh5Bshk1HjL+rYCqyfnrgPL7BhGh9G09z5HuQy7GivZbi5dgtkWwAWSvjyFAYfoQ3V9I9hLZ
g9l6vUSzXMDj4z++gk9L5bPyabthp7nKa5yCvt7j04zh+rrfLtZApSv7g/1UQ8+J5uFDL4vmDfeL
nPRxaYbpCCCbOYtyg6LLfjZXRfb1KGLahYCQEf2se6bG5jGjrBJcmxYJF7fdMVQ3uqisuh6yzUmc
SR7KP2AoGgPo5Hh11xF3OxziLyEKqblx67LLFCxNWmvIDJBCLKYMy2P8xvkTP0RHvntPvsx2lSIu
Iz1fW79yEUhBbg6ihwjbFepc5l0SjjqqkGFpWYj0QgbNKEknCMufScA7h0OIpocNJTuVxb6r3qvh
bJ+8HNFBAUFhekaNya3DKLt3ML1x8Uccbq1utOr76zyFG8RVyV9RocqZVczvB0BnvtIFYycGxGex
PThbm9BNKqTu/49gCn8Ni7J4KhMWwbwgBT+iv1N58Gt/33iJBaz/e3eCFkVn4vKHQpw9+lZPWkdd
nstvFbU4mzo12uEM903PzlbzSrVzWHLz18GBQCj2zendd/QtaDyOsQFmKXF5Qq9uUORBKGAwj5yn
tUATGDyHJ/2CPOHpbJeo0S9xR4THHFUPIKy3sFWvp0ftNlB1ak6Ay3s54ba2bq9z50+3GbD81/Y7
kAXOVL16dFVw7HjFw5z24xN/TiDo7iotfQ84kLYTQupq9XXXxZ3V5jbTgNGnFg1bPmGVlssASB5a
yf23YsM54mSAv3jw69wMb1QGscBBkKHp8D1XwNSjiv63HYvYUKRXRi5SNYAFdtt2cqsvqnWgApeK
Du0eFnPZhPf1iGOb/QUjomDoUSoSE+kUJLgJPO/8e1xL3MYd1Ss/FsGZdnuAs/6E7J5Njv3y4lbt
sjcKpjSkEp6PCoOiAZQJ2bQVAqI2vhrm9ZitqqsNe/Xi82JrylXIEQJPEGo9ZNyKkuk/yfQj7qv9
7pYkLg+kI4LdSgGKBRGgpn6mWHXTwuTYJYGEyyeIb7Gy+uhvUxzOpgD0ibMDCwuHDkc46cNzRX2e
vMy9C8qK8aguCwhPqay61CZ8IumRGpReKqcauK3BBs8XGl8xmfL8hz1kZruVHQHDzsoVC24w3S12
NLZE7iHr+EK3WwspW30cv2p08KRokuNPKzyGTt6aVZYoP3Zzf/I5FBHVJSZL+GvKEaqEPcgjIbnV
pgA4dK59qs+Q7FCu6F7JDQvg83dO21k7/nX8QL6Wv0D+z3EhwhuMGjYnkRy0k1IxGRKuALZx3rrv
9pgGpbElu/DrU13z0XX0IIU0/2XDizA6cPgOc0siA/nuwe6wU597xqv/Tm/sePiYvD8JYeirliyq
rls19eDuRD4fDoG3f/lmChK0pL1WVqfOwVDFGzpLQr0g2uzrZNlYLXNEWnuY1L3efZonyTvGk+tg
3hj1MLB0weig/25YdGx8D+MODmUhXtpN7Z0ONWUsu2bYnkjqWM4SW9Dl8FSj6xS/qw8jkjDHvMlm
iL1LajmSwM5rSDBRnqiGhuMq6syXUWyeOMhpfC3DcLX2cEvNKLbVxBC5MoCvHjYO7MIfeM/YKEcP
0QysapnpucyToPPHgMN2SZLsprLIgrH+FF3E0NDQsBBgfwIYdC8sDzh+9oTq3SfVw1fi32BxGe6x
95D0VKRyak7jW2+XzJE8XXNwVl8yhEQnPmvFLsx0pwb3i14zA/Xq2QmcGwNLD5FRSWhH/FcnlaSE
DUtrH6o+rmIBFB9khGw//qNp86HpXfYJCAnv0ECrCzRyzv4x2FiAGjQtFvvjXBUvKLEOa1DtLlMu
VHkC4Cyhoc78z7TEfc1WvRwo1NjTkyv3r2BOZ6VCc8aQ+Fcjsh3a2mJwqWKFRFZPAwcwDLBR9i6Y
Oq5U4i57zPtYo/EvdzBxqGU6/l09PN6TxlWr8kCRHHf7mPs3lU1SdlTXPzwM6a5qqmeAiuZbxDip
m5k5l2Yuf5P/ZpinGP0L/mLrBVnLROeQ90qRvYLSDGwBVJV/x7/z2tkgZ/HW3kM+Hvsfi5oz6jZX
twvbH2NC/qANo3RMAc/GGR44b2Brl3/HRrq/3bq5zxksCmFLUGqhESXqL71e3bv5kmEKigoiWTfG
0gP3ZxzmQssFD8fsimnkvPDBxSvxvRR+0Uz5WJC5pb6v+Wlyw46UcAHIpzXZcGbyAaIoNwImN44i
SHDlO7nmqa2uy2hzMrxPwfJkxDgGC1wVR52teMAKfqzArpS46JY44s4OAI2JYxlsM/zE5MjZvkPQ
HTzcEbcZxcVMwbI6swjt2Y53I9aEgQDDxU+25emhlOeeyX1lQbf/FiOUR1vo53xsr9YrctT2io0N
q9+EbbKst22ZkeJrFXFoaf2MTQNCJRgMMdeW/a2Jfx3H6TQAMGdjjSIvHDoQvilSssoyjpN9zwK7
+94k3jsuWZ6EAIGb6ndouS5aiG9bzWxXEea0kBCf/YS0nygxYjeqgybeeG7WjnYWEN1W9HpS0Yhf
NwbcuNY3eH16oYtgdl+Tdy+2er7WfWQqFdRODKsPap4SIkJXZOQ2NTBTBbLd0hnjVNy1yz1m9uRv
EButawPMmoCCOIoEnTwuaOQDcrXMg6g+4J24+fjYZS/BuCUZp8lzCJHubuxlE9dmz+7bHjSCbJyp
21B/LU1pWqP8ySiCPLQpKd0Qxg+IPByoDoiCQAGlYE3rc+AuFRtgTjjem9JYRWTYRZyJcMpVPHVc
MHJ+5TCZy6UZaY0jbew5bXzPwdTxfDq8CaJcP/cJwmV6MLTmnC346OezzCeQWEFYEswF6WC9qfxP
jdIVLUPI3xYtty84D6LhXXwMU0SXaBwboYidvX8oi5XrVhuX/lOlx3UrdnJFJQ+s9fXdLvPRTapn
0X3ZP6hZGk5XIspalMpnE3rcVTKy1xSTNVFK/5fMVweVcygaUv+U/kWQd3Zos/8W/pn3+RCWhU2R
0VPTUdNCt7ZThD3QJVjDfjvj5W3aScpR/R6OpqG7AmX3hNCrWrOXTYWU6W2fot9MoL3w2r/C18qC
+/TiwkMsWPG4RAa9SqXAqzK9d9sDsLWUVemDyGmATQj1eceTxW9QJpFej/G09KiffhnqwR+dvqm1
wiDRWPfIZbb+C52TjRipU/ES4xrKfko2bYTAsgN8XthOEw45i5dVan8UOAW57veKyVKDhYymkZha
RAXA2WzHjWCWfCL1cPDHWaoGbknMGWZKFeXsVQ6GMn/ZQVBLkcUVtk+lbqN097eli7I8ZL9jf8WA
2ak61oK3PZqOio/z8B0TfqDfbNcn9KYw22elqd2ED6hgroKaH0jEFP3eg8ZRll1M/3gY3DcXmMVx
EPrW17nRk4KjEwwOGjmbnJyg8EhXrkp1M0StD2s7ruDM4Qho6qtbdTv+IvkuLEmRXZt4YdrsF5UU
P/rjRqoHclIGaDcOYJzxJew50Ru3PdqvHjZ8mWJpzISmirVcFDOqvwjOeOMDw43/kf3QgDmqXqfe
L/tCaqhThXzWb6hRbxz+YZW7siRCOuWU+Tm3yeZvjyYKSwCObgPrF9j/xdzuSWai6uWs+TuqFnAl
NsyN2Xl91EV0aUxWuVDPy/a0Pkr9Rl0jn+L1VFCbnslyv6W/NrlE1BISSJ6+0GjgFOAYoEtOvvXU
lIOh97YKHPnluwjXopQdTbkKnzjsf+ilb/W2Qq1TH1dxnjIpxHCUl2yk0TmF+udbuxXj9AmwAy2Y
6howgZ7aaaOOwOzVFNrfQp6ULs2q5bwYsMMjoe8F+gJkmVK4MXhV+c+BsmVfho1o2pbZiUEXr4sI
pjM4kPdYcw+fPkCn3Z9RtKvbwCInM9I2eQi7ItbPD6m33S2rz/DQmSMmRehIRgtRUcAiA/n/8LLF
93PgfbU8EN/cADuZpPvXeFS+Z1SUDu28RZmfQL+hQby5WM2rfQJskId6RvFH0/XHT4AIkhIhQ116
aNTczjfQTzet7Y47pVJrSvupmzEzRINeOuBMvgxwDbEHVJ67s1vzxxki8u27PSNQM5m5FQXabE//
Vb9l7CguCXF1m+AWbaPTsALTQnRdlGKxERav+RHewOWRNgjhnFPmld2VuMIA2Yy5sWWgw4UJIS+G
aNvsiTuaJJDaa8DKQCED2Mt9F4OKXrOfUPmxwVIP9qlVK6QOTMjpHS4qhLlcYeDCnE8/ylolcSlI
Pxm2nINK9mIO0LqyGCtZCSkIWuhp5xFFqka3p+tTG3xo6m3MeCTqMQazb6P2AeKmSAgt66shGKzx
rxxAiTEp3DOZanoSufLY2NBlkWmyGNxw0Hw7E0XGxIn5YRVMrHApiqHud9A0UuDNXLKLywV5G1jm
iq5ctsYRYZKEEk7OARXBC8ED2UpgbJDHSOjKS3f75IBbvQSXPIb1oNA9JYaSOfv6mOccb3YehCUd
U2mxeqiYgMsSpSv0PcDelFlhE3XaksguYssNwMoB5EVg3krNJRXgJSJQX9+NdynvK225CSPWG5lm
xfjT1lR5TsCjBcyRodgzFpfhkvXNjlG+e2SDrlaLB+BRWgtE87d6TYuPPL2CrsVCGqWepZWWjHUp
R8lz/lqUkknXZVHwYHqYBYdJ9fLO9ph1fmQvUNZFCch77TDDmt5FHBhI/uKokVVxukjLlgthlYDA
GdDuSs1kxXn/v/r0X/tXoLxu8qZpN+8lK+RPy6cnqvMMBzH6rs1N4ozbkQ0lttYuDfZn9fUlYlQY
kTy0/6sOx2EvP9/tagZ2JBYU6ydoXlpYDla7AM0rI2S1g+lxxhn5u41rhna63DTJwsJ9II8W/w28
7xCBouJOi1a1AQToVjruZox33lCYpBL3LLZSRUmt2wtHlU4UchuQsvimSSr82hgSLMwqa0fQE+iM
pJZdYOuxk/a0owAeIdsN/wxWhxffXDQvEyXsGXO+8BytTuZEdcyJI0GS3RuMHDo7lBsM2Du5nrdh
T4+tfzN4/Oo4gY7pP4AWpSKatUvubaMITZDtWhy1T59Vvd+QGhZGD3eAfDw1AYfajXHKFVwlMK7q
WYczXcp5Z+4wWvAOtvGhf6KeAIkNvXOzxTo+LEjYy9WmZd3sgjwF9xYMzhLZYh7ZSWOHrb0nZiwl
rYdb0M22/KfcVHkIS/UsTxSQV4jVbEfoDHYPyqT1j5mG21GivwY12roBWvX6ERFVUvHuf9AUtp5+
P36RMKhe+d4ooUwo4/3cOydXUCVkSMxALJngNIddAmLJu04kYBm0kEsBxerd72uqNmEAxjkhXSwN
LYFPpu9PQ0ngkCGvc3/oCTPPu937iz3W057NxTCL6KbrXNqCLiyV5TXXKNig6sV1UOWsK7Npj94S
ozrHGBiH6YtZ6wZq7gsWDSkbYD3iBR0ZGshGDGtHU9lGJ41dGLva2dAoKmOItV9K1Fr3DsiBzYTl
oaLr92kB44OMcX9oq6Y3sLTbBbcIlB7BOqitMR4s8ZUP5rXCmERLgq6pVLmWLmQc6u6520Zvw21M
Z2arPVpMdIGWdp4ArdV5jYeIqx1l8yWtmSNjLEVPcusjU1eCkJxOjmujb9AiVueNUC/vo7UDTMwP
J4a/qgbPGxBkyHiEbNlK9sI4J/hvEGTaazkbb1u5qLPCVu7sAOP+WulLWIoGSaUDGqvvTcRfnyoK
+CZBukNwkHRoiz/zw4C4D3XXHcfFZWRPF+CCaGpwgTrFr0mLZbeJWwNwFJ0tEQZTd9NtwBSgcIIT
NFwQ3NyAJnIKFoosEZFOS9knX1+dH76hBUJKC5KYD00JLvzBf+TdDkc80DVmjXo969237zyQKlLt
BBRRGz9IyqhMPA4DWkx/1sW0/hHpk9WlMtSN4IjDqBoEdTbUkRZKmHse/TuC0DvW5bUFhQO3ZN0f
hOpUpXlaHtRPfVlfVxTEmDLlxyJ1r5muj9MZxsObjOJ2ctw7pqFLh7jZdZkK/P81hQ0avSDIZXs7
wldbVnA2AO19lWU9TRte6BNh4NAX+5u1kFr5VX0Qir54+xVntsLt4v5UxjQc9Ng57mI3dIijprnH
eMDqy5OFumJ1Hq71x2tkgZqF8tMJRoxNBeLJTTbesbM3VjPxkYL0mCBYGpe2DqSngVsK2jCIKhlE
UL/Dagsxv7Fj31g6oV6z/OInxJr7+NjSPHbHQPpFkAHOmfI0iutl0234N0LQBbzo/EXUwMlUO0Er
HXV2RXf5czsRmkgfYkio1fuqt2X6Cu3TQ0WsyVgelio2evHGNkeeBAReU4m2D/mDhvYjzSVTCBHY
tRKIgKSLScg+42rNVt2Qc4F/AqJ4Yc/Tep/iaB+CBwGAtVmYxjt3gW2v2CEfcwq/xOjKvOFv8aX2
w52NKZ34nqUjP7byYMB0ADaoFuHaTKX4HvmqJjT5j1LQtUKJlzNEU0+CBStd6B222Tl8XL8drnKS
T9MNn0HxEpPu4FevKpcjQ3lFv4bkfnIwlSdOp6wYQWOJl60Qqs6EoSosSv/qgBjp5RHsimNb/9uU
CEqnHv5B+HN8TOWnnmjn3sX8V70Q54Xf0jnoTckB4slpzu8h0Y7bWbC+n6NIRWAzBcR/52uFApnz
IA2UZTOOo/nNaIj82Q1iuGBVWAsyeEiWh2KZy4Mf9OK8GyEBYHvPnH69jFV/QhOCxZKyluu1s4wN
gGZHJU+pngFY5Lvnf67M7AR07Es+ybExcct2aOSmc6688MIL/nQOdjybDAn2JCyC7Xk2mo4KnGfy
5CfTjl94R+iHkCgh1iN2+zovCsZC9hHCFFvuzdSybBb99YSFalWKB8NhYf1Ep+C9uL474P3P1FD9
3mim6jkQsJvZL2qhfq63QIuLn8nCMK6mkpGhqPhYmrwtqzxJbSpmLBeh+QmDOmov744eljd0aVa1
ixKTgNK9HRWX+FiSus+b/eYDJ0vklWecZhl2b2O9hxO2utM8cSKbE9s/Cz3mxWrCtzgILE25BiAn
AV2KkLRvmXYh08iW1UqeCksFKxexQG9VpyqhhBi5JU7ZAhRqSYKziYx7X14xJXyLyHMSo6Y7zqde
NsTxGI78ezWlR2ph2aP969g5xBDLI/CKESKoTKD0dtD+DGuF7U381xiqw/+Qmm9vJN8EeJ04KNAT
b0OZZF4J5xNfHY03fMg1yS5/r1Z1J7zu7fL470AfpUjA//5ZiB+slfHKNFUVNAjQETAaMo2SRy6a
eR2IZykKZLi6GPWCU6nSvP3Ltei/3QP8QU+2lWBROGZYiYfSH8C43qzUReGY9unwPBEPVNuK99+a
+v2zexOPNbx0gcp6hzPIbwdWYMfWtb9Wry9GznjxCwH3m0VqfeIUZSD1XN3YiVBg/7udQNSKcM00
tbwCgPx6RekU0SZDF+Qv/khVbWVsC8Tr+6TVG9SZYaN3iQhSHiL8eJaGbs6GkhHoZIS5y+2AM7X4
8+tXRoNrnI7yrVX/oUDRhjpMBvIEOCtE3iDFTY303ev6skjCnedL6zN9A0n/RaZwRvlSmfq+Ez7N
m8nRPDoGBqLo9z3mNGNKYWuUir8iOESelVoHFF3rFqDosTFhSdgJi8obQaSRDzYGTs+WnasOxXlI
cBolPp9edGElH8KeBrcWVx9Ho41rlTqsz4I+tTteUx2cNXCfGms3QLtSs3cZRUJhBqDHuzuofMVj
VZzzRKSfcqaBBAgnvI0wG2FdUKtae3699AyyT4T5aJBhaSqzmefKWVKi18ShwPcf5gpMWK9o2xl/
iB84o2+xvVajjjQNX/6uPfQchgLWSTEEct7GLXDM7IXF7+W1S3T+DuZ4gnbwvt092t698kLC6NsC
LxsaSRmA95iGh98kqi0DPhagY6CStu9iEHgYOooDinsAm6K0H2wwsaTFCYKuUlRt7lCI1lZdREJs
H2tF0IpF625W6mCZeRw4PrlmlWBKnrfwLn2cF8oiJJ5A+mMAdDq2Z05ZpkNK9NO+MmIOFYKKdV6x
FNvsb6kbnKVk6d8nA5PFC/W0zBLGaEm0dWaBvPh8eKJmDcIcvW9qIa/Pw5aGvjNeU5SQmNp7cKvD
cclFbQxXOn3Oh0OB2IZBulnz7K6EwYSRvLX4kH/8lMOqbbOL4EYgAon8hFcsVDWdxYdAKK3kZjb5
stPJEeeBJFpFzNRr8C9/hIzOBVXO8gYWWPGHqTjM2FqYC6SS1b9Y/eAPwRIGu82Gwei6ycYJpPzY
b4EKBdgt40U9XRIB0jipJ9KwSs0Bmez+GU0Dn2EGcE1IKYHCvH/8c/Z6+QkFiuKJLIZezjTTSagM
JXUPSo7HSv+wjzw04T9alnoUjGNQ3lIdm4En0uSVuqsi2ITkJY/AOhHmjAFbY1MMY+CTSh8/MJ1C
VSNEtgT9VY1gOXHHnxk0gtKutjRu0VhtF9PGrs2W6YVhMDdHhPgow176O6xxRJy5n8xRCPbIzK/r
KvluriKT+vkJZkWLeN5DN3t1G68pGfiB0NfYoVz9ThwRhiYwmi4miFO9Kh1hl4iVTGnpnsHixRP9
uREhdbbry6jbPDUUf1oDbS1tCOwR734KglIdvcRzzgJhArl4d8p1t++iwbYZuWEsq1AoLAL3zeTR
j3Yo+Ax6BbnJp+1uiASTUlE8/GicDGN36FyOg/kObS7FCXkK7yFPFNVwWIMuyT4ismgz6gB6k2Ys
AULM3gGEst3RD8JK3AWmeFO7l7geLlGaL0v98+oa1f2oMHB7m3E3V1OshDI1DnX7qsEN00sjQhqK
7uF9+TGpYUOhV2KOng3mUGTVQzhuVYQsjVFFLC474t46uNDbEXEoLb2ziaH50k4XtEtD+1fJ58iA
q/UJqIrVc1rhqUz1aW+SSg0hEsviVPZ4NSgsn8kcWRFuzn63acqHdSfESvZFboN53B1DfjiBOv3j
UMUBoH71pDba7Ra4sP4zV2ZwhR2rZos4xBXZBLu7qkU1PL9liQUzsYSkEAKOKBDIVjo3OTOLOjZ0
Aq3JARg5e0vRye+KFWeBws05zI7hxwqYAgyQXbqW6UO+wgEaysx+j1s4sjiJ8mtXK7yVZchwbQWs
3VWi6NnNgLB43PxYduHTovvuJZWKIyECD5cW+vlgGvfkb5d+XFn3xvOBu5NkdwLeG+COJkXeqU0H
bWHlMM0LEXFDFUh16KKwZVPSq3WZ7maykHfjX7JT3+AWgd37jUWKdQCeSJxglOM//c7vHDGnvNrj
cW9y/XoicBwtLgiWcmB1V/VyWnVfXNizV4/wHPskeEfM/LQjxAdwasYeSPVmZoYapgBo4OMnpi/f
vT75RC6/K+6vPYDdsw9nJK2l4zWCKPI1mhKOIjJ6HMY3+XnpS4VJiwBNjiUY26Y53+RilxXjBY8l
BrMBYN7PJowsRvf8CPCQTUq1HpQD/UoHeRohr056iLx/1Cb0pujzT49T1M4prSg+BXkWJoT0DxVY
TLKAqgptsF1YnKCggwYbtrMlAZ2RV3KoiLxmEegehmrL3wXXdF55fsuwsksY2DAitYGI8XNCHDHV
amzZQ20iCqxtHLGtmvnRGsmUSMgAfL5UvRjgREaBya0lWowptSKo+3rvvx1l+CBagP9qVYWljgwc
WsGC9WDdHEKYGoxoHc5CWyHfcyu6n2cHOCWRIm8OzKGqdsqEOWCbYQbYplEndFPnhew7OqywZwg5
ykar1WG9XL6ivWla0FoU09BI9UWeDs5wFkH63e3d65Dg0zwS7v6yyH4wFy8kvKOELoa7tlL0cIAb
JerNtBXbLIAdaILaqcDJW/No2jSNddND84HJJHDcVG6TYg8HbPAr3khiRhAwkt2Yc9Y93YT4TtdZ
dYh5LMBufCvRCNvfLQWyKAnVpxyZv+cnFqV5HQU+xeARJr6IisUnRsVQBEfGtlTZZvpkvfMGhiVN
b+QY7bBlq6JJVHzvt6vVBQD0uuPIbpfkgJ0dZn036hQ75okCexm2ULM+QEEnUh4JY2G5GQ2ofIjA
dNFQDuAsYnKP6kYuOTc2vG0OhEOr8Ozy0reG2mTOm4JmaP3SryEGa+l1X7wjJFgPv2Nndc7F56Oq
RmyuxNBmEtep/In0pErN/vXn6lFNqhx4l2syVWdsYQocTN/+sB2REI9EX+BlKzYjadiffpFHaRES
1jeUn8LHm2RQGv9P8vQIBeuJDFsDmdeNpL/R0sDz7uCvvv45VHGc8/k7AI+Uh2gh1jF+HVgezXYw
0Us2m4AvJ3GvPsi0KfMkJ//EeVHZTMea1zWI14mjnyZpeN6HgjQWfssiMPPh/picBfVKQAr+shSc
cm2yS5a39teF6fUaq8dJOuhkMZiuz238++3AnkQCZ6PUThpwpl770WTDhrvHE873mlLgBYduYRb8
Pn36qVg0hlz8JaOJzbTACkxNGJpv5xcijWYsVR8plGXGd0x0k1wgk1JsAj6YN2b0XlDDoe2ob7Rp
MOCgcexQrrZrZ3jt+ke2edA9olj4zecKOYnKfSBOldEZl9kPAnv2sNMVsJF+dgqWCQeS2gtQclyg
f2Wk2QGezdPdEMcfzcM6c4l8RPAT7PEQXjbWUfkmfdmlGaL5iQqsBS9nbtj7VCKSAXaPGjd2sLqk
Ptfmu+WwTPzi5eaQkvU7JIU42772N9KqWVS70v9JX8r3KMrbTmj3h22hAB8LgGyT+sm70C/Hu2O/
PoB71q+M0W3dFGThLcgGx69g/NeAzHRSZOmbulysTrTAEoBC2vbpmVSbbbltVleMGNIzhSc+bG+/
yL2fCcOkCenDZKeKzLpHe7ZMTcIvuTs7JYjCebbxBHNmhfxBj0GsolCHhasat9Teo9en/NWpOBez
mxzZlg3Te0J+nVHgpmq2nHwTz8ADBLfRPp3IJal0H2lXEX47gW7fmsZGcflUtfx0k63pHdsp3EL6
6C/EKTJGdah50UIho2xZjFhuMLRHaTVH4YAWivhe+ezCX1dfoXd9HDbQqPjNgZjnx04NUA4nJcqI
/jfOGvHvauooMbTQ08/8xQeNYk2Jy/oe4AvH4GyESyOQdlYagref39qgbgQji/r4gXPzg9yZuPju
aIBS92n5AE+L6fdbvB1IkwW1h0YNacSKLwb7j1RSzjL6GIYADUhBX450GMKn38qTkPNZ46iI8VjK
tIM2l2sQU4mnIQ8eQbXVZuOMXYJgh+Tfv5Ny7cvDNzoSKcuDrDzHyNMFIuplkA5sF9FaygO4dVdA
AyVcK7m5NLPtqiXHmiXxfqEsIcz8sHD6fYiRtW7eqewPK95I0o3hyqP8y0YmUu1U5cPVxeIxzUKZ
g4cGyxtsSE5FBJjyxr2TeIiP+6cmvzifXODwqpBfjuJijLtsCMEQxwLH2RbSUnFwkMbJ6/mcSjeE
hWr5Wr4hB8d3weKQSnjFq9rcyoVGU+P3iOxHCwz7Ar6p6TI5411OJs4aAqNeVNCKemCypS0oyl+i
YtBmY308qvyO3pjeURcrL6ehXV6SQiV9U3QuPzUgzXiHHnfYntZ3o64hcPeXKf2Ui65iyLaxyw15
eiufBGB9BImQki3Cbbsk/HruuxglhSGmI5NP1cY1HJ3Qy6fkQWZuCC5f99+qaKrqrsIkgfkH6M42
c6TdmT8kzJyU3MxgC80OGbKsFn8mqfVCxGoZyjB41+9dRGuMcMNMYWjEZ9nH1NuMIRHIJSwctyha
Povp5SwiW2Z1K9mNgqAc1HA24b5P6gb5bZnsefBabJ1jypkHSTRqr27exsgOnXNPvNxzOG/mCwKj
ZG8xarpugdBmQDSxizIWG89/ejFv3a/HouDmgU9XZTFl2t95jfurTCBzEXCWZ6pewF5xThz5l1V9
3Yb5rLSLaS2RJX1q+QPeizgkZCVdynuh28NGf9V7/jYTYD08JTPiopHF1goi+jJafpTxqoKVbUzP
t5NfGQN4eoEsxeepHdCZ7meXJ/zlHcFWUs8l6fTb2sglpUcsE5FNh0V2+sIk2s8qa+SHuPU2h5Im
j5ir4X/H+ViwivrehUK36f11A5TAaho6GEx4g6OkZowcx0QDvMe4c2v+CZ3nH6yakmeTKwmv1+RW
Y9BInttUYuAKsstGbTkcsmBDC0f/GL4XGQwZ5ARBXBcPN97HjjcDQlvQ5x8TH8/I/OWm/SQT0pCz
gOGkQgGvkvt4wK4Sg4SDkl2LjTA8LN1jBCeCaE+MX+RT4gy9FPEJeXHWh/ZyGGHuWt9wrVVHaPEI
apOX9kDW3JVpovgVUMnBY3PopiU9dMYc9AFSRcFQ6FbZdWfG6yiiSa90c/AQKY0+DxAnSVtVJBRH
sxLwSBBB2LoVTrGgS3zrURwQMIlWOpHlWGKQugDAoLZMaCJ69oA/JuPXZUxdGm+DhVSyY0D4g/xz
Ei/1tFziemsInD45JdHVW58gupPUskmzJxSiSd2knhZMceKOR+D9g4kt0ih6ToqKvP0QeQVci9Wi
iMZf/hxCgcnzDd3JVwG9u/eCgQGQp5aISgeqptbq9sPTW9O8ao6W0bRcEkpUU7i1ljlPEGxmih6o
NH8/cjw3N8dvy3Rt6RHFuypWIcvPUhIu463Z5eAQROu5vkVS4DZ6inohz5bfl8dPQRMVA0dtn9yZ
VJaf5wZT8AaEzLbKIFnbhbMj7jtBsC47DAn8a5P4GToW6xr0Y/5I823HPhUpYN1Q9WTgjPnKof2z
amtjvpll9rnMOnTdlyjwoJta2rirO4xCF+IDXNoGmpWY23bnvOgqt7QMY32RExRrOIe5WvXGHUb5
S6o7s0JVpJd0lEP70iSZZqQK92KKLQnmjVh9LQqpfeYCyK3eYKXX6n4szP2x9wGEpRsv3Gj5xCRn
d2mf8Qv3HPizl3yj9ftNIn1n6lGWDvBZeD4sLUtVRmYwwI0BJ1VREcsaaiqiX57RVxpsEFYiJtED
YLw+3SRJOC94Wffj6iXcwUHz3zss5xc1BJgrR8UTaubRovdxPIGW0kHEblaw7clL5snOTBnase9v
hMXbGa1WQdWrBBkYtTVXicv73pwCs6HZHamq7az9eOsrKi4TFxJLpPZC/mnK35DnC1DQZ6yXBqzA
NGOTNXGEjrsfF5oYg1ZxlphvDvnmBy28NSxk3xPRfzxLsfVKZD0SV5EHsIFTSwqS7vwzy8T9vOou
fnhjCOGfsWifk9xrjJ9vW2nUbHN99XQIYnKURThPNDRnfnRGE+OwmoK54AtYQFKfmu2e7xF/0SuX
PZ6Y6NM+SSzE0PhYhWDynSt6odDiNTt5vfJ2kRV/SP+Oo/VfCzHTXYyR3EabbFWdawjxJRHz0MKB
mzUdx8xNazG1Tduh3d6W9Mc0eg+jEdHK1r++yosDN/C5/iaaInPqc742ZdeqkAXSVghMqJIw58MJ
oeyCcdGKLL3Jh7zJONBHt2MImrDhxl3HiqIQc4eUjTWdn2OYrmBaagJpO3zTLwm9qaj7YNHG1nRO
Dxo1nRt27h9PqjSFOnBVVcu8JCG6O0XN30/Z6ZMIaswGN2szqovC/RMN5aYWdTBFqRX8MLqq2YCS
XSd55mmuN5K/RNGcARPPIKUcen0aK7OqJebvk5ZikD5XxJe1KRuIR9BU+W2UU6FwDmZA7xx1Jf/J
JjCZvUVgr3LsOGy4+iODuvpmEpR/9uRPPV2YMWPBkSyrwPw1GlzsdnvQFiQRk3PrSAdal0I3hzht
2bID55Lm/OtPiEfWvwN7P4pCytKXpf6HSIxrX3d9iuXRwSdhS5rGlEJbH61FEc6NxUBhSYaDrP+N
w5liCVzgo9UEhUNpyuBXXBRlPdBvLskvhHL03XLp2OjgzZjnEIfH7TgZUY5Ui9Y3smuyZW0sakgt
SYPVnL/gfKKXyZjEiiRcLfneTWdW9JBqbQuA/VADfqlABOhtNzqxIMcZbuif9ReIQgIxebEVQQBG
ODV2g2KcQQ9u9s0TlcLaBwwRt0q16rZ6BFic41EurHzOePLLv3NfTlAnoOC6zkmhAwFhtmQWZrql
lqjXLo7FiAiPtkDDFh9HvXtgwQJtcOfjrjfkBxMrPL794MFlST34Qor0kadeipKMm5fykhvSgOGQ
AtuSFf6VWzv7D0ukJHwiS5bkj6pX9OKNW1ckacQXvAoIfMqqKwdGi/nIV0eZasRpzF7aqBbnWpIO
uxF0V7//gazm5vW99NJzQ4ztH0AD8UlMsv0ELrh/LYnXlauckAXPuyKO8F/BOxDVQL/cSpQUxP7k
SgK0dF2LLk8Q+366zWUNE9FqlCAEz4SYgpDq24YFXMluHfD7FIGDxNgNNRWrRYU6gcT/x8pfn86f
lxDlAJ0C1zwA3s7nM0LqZ7iM6mx0Out7QlAqdJlW8tLBowq5/zv3sIxBGy+bIQNju8bjOHahKUd1
chfb1hXl4ZdrlQLDushHfjKc+vhROXmWy5/tIcBTXNQzQF1mQODvIsAH+ZZoJpRp+mIJ3lamOlw/
b6mNbFxwmvNzmU6gCy4x8Fntws58paei7qqRmcu1HgwVDG1eEeUR0Elu46oVUb5OtccQkNo7KIqd
1BcfCeY06Q85HoQ3o5eY01haW1pW5FizosEf2HqjcX2Nz4R19ZpUyA+3firqYylxa9EvQ2SZqFWz
CLzPBMsFSINRsKTTXl0mQD0rFgazNKLUK4GQk05QwOOr8h+pRgsc/ilEv6Y5fILjhs1kl7PttQBl
cAK9urWHgBHU71GhRfL1VkK/OknnWGyPnXNRf9t7cbAO0KKd1TQvMaEClBo+TH/npNOGwxouR2ii
CIq/wVNU02Atkl5KBLGLhZzY9RgiZ9zdOpCPpNvnumci0qGzFZSY3+uhvJ5+KmuFJxPzS34luFk5
MU2RawLsdwDNKNZw4SGiHvP1sIH3LGD8I8zQParw/1PNK+Cmm1q9O1/EoAZBRl0mcO9miwTuHO4A
vWhvgko3s8Wj0GJDJHC83926gx8EFWoxdGczytSCoDqWNQf2xMct4WMLFR3tJxZemRQkfBQHDvKr
Q4B7b4ljQn4cZhyCWuJm0STMLR4Q0LrvZ1I969yixAdOBdQgw4N08PguRkluIJLH5/LHRAU1AT5y
gNlERSIsEx2DfGtxZETTrUl/4bAkh75zecB1yXUMCBQOW1wP9C8BvpqRZjIosG7PEpsATLrK1zuF
E6fpJP1O91+m3j3YSwpbVBErhx2iOqA6Gv74BNlCoemLsT8Do7XohmqzJWC4/nlm/IP5c+Clgzh0
Dmzi5yEnTsDNp97nLpvx1JxgzfJYGMOULyoU/oSKMHk5Vp8pGHcL7ws7m7nwbe3Uogi1/qZGgfwV
72gqqfuhluhazEEHL42ma1emy0bQDw9ZQmts0TKfzzbj9ZG/9FS4A55ERNCxAhPoN3uuWArUsieJ
B1EOX3BaoEAyAjON3g9Je5qAo0TVgsWUz2qXgWRxdbbq3KpAdamsYpAztzV9m037l2b3gTSOPolO
twFnrzxTIqCyMSfhdrSa2RCygzfpz5fZr8fxFkrXq4t1OrDIWVN2hyD20GDN8Ss6Mcw2gtXZ5MTS
CLgvPOYrQ7pwvzIh9IZjIpYOrrSv93tKsj0hS/NAcfLgU5zIcg66EHyyf69H52RfPUFw0hwvNGoi
9owd+pDaNRamxXxphF8t3AiFd22T0bGbtaxxJ/J+k+0Zv2dKtExIsVGwi7ZhN7QVYO+hTDHD+42w
V1uWuvaAjeDcH83kaNw6I/rgVQKzpoQgqABp3WwpNPRPOCxKanVwxRXYidoEf7Mh3p/5/m+Dt4LS
SEqX5n6I6Sp9vxqPS3qaWMTN4kpAjnrP4vvIO/P4m2wvh2r3a7C1zXukLgyLBHtfXQI4g7r2CHWz
6tV2IBEWWMmQHTMPlyUKsObsFnA0wGNCgsdA1yU61aJbBsKM5LvY7X6h4qqDjbmWVgYn5HnSpEIT
X665Bm2eifnjf3MqdXhFpxLBemzXIaQPJGkejELiGv2U8qdDRjpFTAF38JXWagcI7VEHEwk6sgSi
WA5cfbj3ytO3LE0Mag7trQei/iWKpyvfknSmSdR2fjGA+VjfTIu2y/ut4rF+/QZP35DkZYK8IM/A
48TQ4PG3jzedeJeN4JTLl24T+148MZKZCJ+SMA+WS2xUv+f+3mTrNGDtu/9XBy7g4JrASjxJ/DKy
UIOR7FNjqR+tPaL8PWEAc5WntaPctnhZaOnoBEg6Jz54XLmJxJbE5bw3h9ceKkyzfObWrPwMMJNA
8nxtH7s2OPBhPX7BBv178H60LhqIdnCtt1PRCpcCr6akOMcRIEnd2O8CjZsinjo357WgPZauGst1
sn6RENX1bucQYF5H1CIFwVZ1X/50ho37EksIpwhqZu461YQAQOvnVVwG2cBozPxuozkDH/o45fzz
b+hDhBEdfdFg8bh8CxKHk5xBzsm0/vWqSoh99HwSvppYzO8C0dgmGmyOhTRwC5OCfanR+YUnWKpN
6tOF5YV9rGL7j8mJ0MEgSh2LWVxpXVw48oI3IG2UuDNIfcBKgApLer5EdZgcSrPLjIT7LNz6YhxM
kFF8kXbqN9IAoNPl0ymBjbf0hymSIlTw1mdezyqGH4oJF0RiWr1/LIBrHYtGVs02LU9Js6DkPf5z
TS/UnlLWrokDYai0mgGIoHss5V9hKqUTb2b1VZ3jhREyHffTNfSKI8bXNMFCtFgdypH9EdOfzSey
sNJ2DNqsNtm4WS670RPhbrQecKffDcH2TtFatLEddic4rF7yrseyqEPRfkB+H6zc+LlDPvDVtu6C
hjRpZWHPM0IQJYMzGDeRSGZtEB5Q3BpM7UQMHrKZ/taI9G2uMMtRR+qO+AZZE67Fz/ThElSflnm6
avMHGQfn/JzyPz7kAjk0DrJ6jmESDuJzXUqHqjd/r3U071jf1HaQmgZ8DJxQV+OWDJYKmGSqvp05
x+dpJaxx8LOXR1h6uyhFjAopKDXr4EWLkiUWjaLX/OMoIKE9FXmLUdUFx7w5ggBsL8hcBuD6ufXf
h3OWLTOvwQc15PJ/96yW9SNctQKWgh2juViYYdM7hVjF1ylCVAXUWvCnDWAGNNip2e8e6Tg5Jzez
vd2jaV7viuLX3UUwc3VAyQJ37rTvdZOaVkfxLUmm73ZNUZAOaz54XfldkoW7cVEbp21GES64dBRn
Eyh2wdFBoKyxMabAI788EmS1k74S21h+zQ+aE8KPT5VaIMj2c3ylq8MLzLZqqiyvPmTyBdAx9ngR
XDMuGNC+Om9gscQ4DePnTmdbZ/gTdN4lxxKjVSsR8V+8gLQjoJTE3VYbdi+f78YCKWWBTissQOw7
pA0OHysXNjy6Wa/LQfyWcBwmB8qBk1TSMv05rmPyJPsZ/ub80AcOtnmhveFgB7DCK1PgDiSLV1MJ
2UymCGANyYZwGTlJsdbiFAw2ot7+HOl26rhsQHLBRUhV7uVVUayIesqujjjJq8NE60flPBHpLGo5
ih0oHR64iyd/TfoBslcFEWML7uy3jehheBvgRGq56GsMBRlBZhcHDfdQbmu1SQ58revEn+cZvgSc
BiL+0LLqNs3X7ZUXWXcfAN3wQbuSjDeXLFiOTUoLI+4aTyZwDAx09CRIf3N1bKpaPBufm2SbBb48
nCaqayFmH9l7gAza+gEizjkW6OnQwAyr2wMvvbSYCD7aJj6+cKrI6yjYW5tyUZiqP299s2en976s
vjmHR3Svb1ERTB3ImUtWFGzL021fWF1UccxASui8GT3wzRM/GOnzQAsmdifBbxaG+t9EV7t6JoKm
N/JmVxuY5El2C+qOipNdyrMd861OHqTqZM+bVcDtxu+OwpyS2qNeVDt4GalQ1w4POz4kaRh2nDaq
ZPf+/tszUzl1BdU08YRQ/QI/+/XOzQLFeGTssdxzisf22cX7fBZUbVsT8jslKR2t7sKFL6aFAYY3
DJq/lx2rKYMzGLXR0NCM9UM0ZJ6ZvrRgWzjOw1Cg4sR3vad6kCXfpDOUBV9/oZIsqcyszyVgPFGc
KgZHo2pQ0jBxjDrLoD9XR298ilAM/8nS+uhL0I711XrqJg1KZc1sOrUHGiSExTF44X4QIIX//quf
AILdGpCSZGtNap40/UU/+Qs3xzInArUAMd4MEwUp+N/e2EUvreWX4+Pad20UmiSvg4Pl46KZxLX1
84hHisPTp4i4JH9Dd0ua0WiT1d0BNRRQutduXnNmkVdxTdjc5ggy/K4h2r/bos0WAETTtGJmksyS
9FWivZSd0LXzFs2kpUpJXHQfBrqZwmrGtysJqop+gNUVxxBd+f7RbttnyYjCGt4v4/+/z2NVvM1F
Q1rrBf1jVpKUqGMjCjAtIDrxeCwneHPzd7etOpAmxC3iugMdXzxZAcVhcAlDCa+au8N4f2fmlL/y
qeHHKwNqdjov/2YWD3WcCKZWCJaFMyg8JvwW1NaSgep+/N8UvyodTKmlPQ6i98ZiYkPm3AjZdy/Q
OVtYkEVjG07u3ve1tbt3t054KAEaRzZeIRdkrUSaKMeMj+NNbjfI/M1CSqzL0DaNsDzvj65AI0c8
gh78wceGValWHtNeQugTenl/DGzAhSasfLI4nvFFRNl59uypvatguh6wC5a853c+DiVkv2asWi93
134/L+cTOjJX6FAH+S4bIU5Tk3DxSq9bnkck7VLyYEO9NSjRUprSSpAaIjM7GKLitz+xfiCz/Ky0
yj7xzgdG0F1NXHmZTk7fKGHaqv7cmJFJs1HOo+tAxa6vmDd4D5abA4+BP505xG2FuIBgvtRwoj4H
oRcKVSTQmTHhXkFFfIq5hxw54UD+URTZ+lEJZnGBouK3QKtUKc0wAQyRmsVYN3S5RZbl/zuynpCp
R36iXI3Sd+WfjSKBitcxuRU0ejsnqBE7a3hgN1H1ARcfZUb3nvFgAP/n+D2vO5g9GfrY517dUKuh
18ndHCo9zUcWHwZjx375fqgvh4jlOE7t9vBHCgkogfma3VuXwN6CICQWPTZFFGTnZcj2GqXvDQD7
8kP3eTyLWO4dpB0k427po9ATw4Log3FjmcpXoBGCgXdi1U0aCtnsYo4FWiSI0F8cKCZQCOW/x0Jj
akwahBJFA5NZ924oUkTtwiwOfA5iYBIVc/XJjQ7s0B8TImlCyAbL+PLQzgGwSabj1rHQzlZCvrev
EYp6qq19p9w7e/XlEKfISHDohTvs++06RDFpWAPUAWRRK6qFPdaUNZmC9VqOw3HvFHXjG7X5aQRs
tC9VEDJd26F2EjLOImBg13+OqkdVSz+kul89CT1AnuA5ZYWPgSD/a3vxb6udTmR2OvYS25MjQCjG
TV66VWSVvHwa/Y5D3ag6Qoxc9cJ3Kt4JnPMDZNfdUXfuHeGAOC2R1W4s3vfZLEy5HBrav6wWskcw
tEUljPyYpmGF+VLthg8+o6Y5alvdnQV0HXC8Y6XGG+qc2VrFG5DPGiyw5svzKOssw7AKJGyOptYL
uIGZMgYCw1RLE5lbwZ0MaEb1Xnb192JM+6NeG6/esAUrBoc+BTz4X60SZWJ+f2zg3MmVgY0hgBJe
qyYwlc7CwMskgcnLJB9ARkVwz269IGtJAzR9PdK9oi11J0lmZ6Ob42ysN6kyDQ0GCyAhSEdhfHFo
v4NKQMv4Q7RG0K4MmSTy4LYm5pUzncRHjNw/B752jUDQbdHyrf1yDY8So4I/lSKexdwcvD30u9v4
Z+dD23ehZMb26UJCziYdnbipmAVp2aYtrFWb2mdYy0Wa7Qkg0Fn2nF0AMKbntOKZ1K6uXzg/P7ao
91CIFQ2m99Y9L5+BSVx6+Sj8sykUHufYnr6Zu/68opjVOBPnrQt6Rsgspc+4GDRAdXqPGDwRhAd+
98/Ip0+QMZiT4KYNOFu0rIgCfg3U1GVgd44gpmF240kqg3A8QW9HwmbEqehAU33ZGl18G1+D3PX0
8IQ2gd30K555ChLOgT5krr9k7WbYoS1rJi4T/JHqZWWvGdt2xt5uBf6/Aa+R/zgFT21Mrv8YLY7+
Ibbm4cVYmSCmuCWB9Qb842pJKfYAS9R2nOZaPK/rPOPYsKzt66tICTm6MoxdhFYOHBhQIo9FU3ED
6LD5h62DFkgJXOWmY8bmg0fg5U/COVPnL3rzoKsbJLvvKhdZuSrmRt5iImx4PagnOOgnety3qZAK
y7UH5JbONZ6ozbaqTHXqEDpcdQCzzzBMwBS87GZRq+/4kNS0fT3ij5hXe9SF0rvhXjKsxXSmiUxA
gexdkNnkHmytZjEW9pdAy+pICQl0fGRHmJ1RvWOGpHCf51C6GJn0m6at2uzgCX/Ogdv2VHLF19fH
FalnnZNhWabfXn1LC+MtZ3nAYhaXGCcNeq4NWVrgyBLG2JKY26NIJU8R9zBUxOdH9k8ilmGhVEc+
bd1tlyGz26ivZxZMrb7n3xJYekBqtJ2Wn/oXuu67uC6OtCihSsLftx6LKt7U24Yvb1FZA+U93ZwE
bcOWu1G4JZp+fYgQCOe//5SwMdr2rFzcvlUQdFgy6W2uYtOaLPyhTfsOKxNSYOYxdSKDG/xRGC3C
lmqhgF9IdM03JKsyVsugHMyyvyhjpvhqZkzepCCTsO4pS/X/wUUc/fEj09yi3PxV2Xcz0F+/1f5T
1uHbjuqHqhSZOmEpOXxSKKCHSfVDeISh/mEC4zGnvWVq0/wlJQdgkZ+Ms7WwkaHnBM2qfgHiIsv8
v4TeI75VI7KmA3pVvapgfEtldBEvmomWO+7koLbBUs1GjXFsEh99Tl5MEihR+7lE9C7wWIjK+W4N
lOvbYfDpKj6JilRg+PyEiLRMUyESANvDqXRAauQcDXvhFZNYnGhAq5Vz0Vi5cAL2x+5SUIo6VRFw
KRfkemnAyentiOk6H+ELmRKZrgneg+yvhfA7g5Nf0dWJAJ2vmlclyXLs487rOz04xq5V+WFwCyXI
pmeBfxNqlqfV03dLrixkAap/23iu/p+0kFg+7vCtafX+TgFB2swPLCtNEldutjOQjUlJS0XmaCN0
1BTGYQPDAAU8tkUvlR/5W35MkZ1M/V9E6L0bxNlDXnKjSMuzgVxMBCMfLCQkKgFGywagpEpOAd+b
dC6V3RavsLh6NX9+MCgw6cE41ogn6MRqd1IFFsgzw/e7bkfalEebuVBL0jnuY+IAtV4TSUJ8nMll
PAiE+KT2vitUEMOIfnlp1SFIede48QINEG+ACYP5McXdNvNEodS2MY5M4viBUHcMm2M5nLE6wEw5
C6VzeBzrC6qwHfsgHU24F+3dijWk05pUygIBmZadIb4XdggD33Kosr6wNsj+Ba8aCbQFuXUgPsRE
vTabGaU17B/jucap5u1WBW5cbJfJg4ZdhUCKPiRk8VPFH0OrGwoaeVJ0+pWwNgxg2+mKD7qx+7OM
zCs5qiz8FvM8rLrqfUcOY97Y+OwQr11MpQbYZCj0urlfKdvMd4Qul9k55gjxanREZ/gGhV+z1fHZ
VYIJbasH2Tr1kbbuwSs6AwUGXNFk2hGrk6ABDU1+cfhG+DiH7o6tg3cHWdmEaP0K3GanmMcV0u3E
JBhiCn2Y4ypW+PePpNMKig5YhCJoRLHQdWKp8H6+kTyl+vqx+T1FkQd6XO+N1as6Tn7oE2kBFsJd
1jYVvEHcVMdvwJwtV3mO3X2gbihZUBMApFF+s5a0OSAX/SbhXLvk1LX28BigOU2sakD6kcgHeSne
rZGxe4C3Bkg8l8JZP/lOJkqDzCC5t/ry087wSx3Eh2+QuiidoD45JCxTgFaeyg8bVgrQgjwtXJJu
uoiVV8TPXDbvIK5VtwwIH+bemX+fhHW/jXKaUqmrUhr2ZqI/P3HqVLzuAdhaSMtskmgBIDOyoixN
5pn/zIuERtSt62vmDRRe0Q7IFr0N3RbbyWzptQUyLtQTNm+BcGcpKxXihAhcXm/xn/UsSg+tt/9o
lSIBDXxWZlUZ17I9cFhmbkeDF/MTOa4nOW4xyfAlkKE7ncmMXzVtz5N33aRXZniW82omssO4NGTm
7lhx/lq+oJOgOrsBiY1c7a/S5H8oOY2tgtd+hiCRHqOS2rRooBcb2fMaFAVn65nq8GHgUug0KXDw
FxN8dcJvZrgaTmlt5HiSTfEJ97o9YVh6Gm4qo3mPF9mgrsswt0ZMwanzmgUAIGJIZFBcbrOUie+F
uRZqFyWrEA8hy2KyTt2S6RT2XlF/TuNoBfGnL8Fb/Lx7x+jPVKZZRm0KIwknTIBDklftKTX8KNP9
oUVq65movt/RCbxmTfHmouC1qgCoxAP4mNv/x62I6h+VwQ7JI1BDZD2PXx1AbCPicWUlgo7/pwZR
NyAQdFcXD/7WCp/fs/PBdXbITGoHJfuvLuGwSyzAb0xTpZvydQSABB6MPQPQnIMuezJ1Y4A+/XG/
e9AZcRwYkt4EbeRC29jzIlSdlQN+D8mr8Jnx+AVkzjrAh9QwvcHhN6cuHIO7WzGOcdIMtWsromDc
svbg26894JDS9Sogjg/owTiWCZXIsVrxgvUZ16HS8IVgXr5LB9xusgTZcHY8ZZY/AcnidSdZNVAQ
FCvFfllNgxsbCcNAR/xxWC0DjkIxV6o43AZi9816dFBhSj4cdyx8Fa5hbKvryZLojnxQJbFlWXBd
iNVb2PO6t8Lthpg69y/1r8t6d8kCLGaPYDywuvPKPjsxbGr3YDeadOsJ3rEobedhT75fvfEWWbst
yPMGEomwvKLuOorTgoWu5oZ0O4qVuZOMzXp1aeVAZCwVK/fjoQkSdwyH4aviGNwAO7mrQvtsONKQ
K4bTfpPVFqMma+K0XNVr5JMGBruXzu2/nr61C8RHysygXOOkBeYjZXfOmqSiRBmkRY+SNQPYvEb9
1OuIQxhr5YRZ6Ejhya7At7qnFtCV9SGrR+kSQSjaTQqwV04DPhJ4hquZ2z691dTEQXNhXrCltp1W
flx4H9vVU84S6E+9wRVBIEy3TUcGcZqhVwWDx4Ge37obfxyfrH/9TWXdcC0zMzXu0O4FhUq2vD0T
xJ0mlVLvVwuxUmsO/UrTaYeaAIBNgFOVKUfgFlvMsD+zjDJHMXiM99rPe5qyLq1y70Us3ZFT7Ib8
+yt7t7SI8e9CWXEzDjKeZhW35eFNHp4Qd2KwWJIulT/6tykZAmVG+GHrwDD/5WfBJ6VXy96+axHn
IS7IypDCeK937O74/jrrVzn/JbOU1WnomfCLYaYZLv9CVjoEVv+abkfYbs3XZJTGlhmfb9iZGZ5F
hGMPesyGvMHPqD/zaW34p494RMelgeqo9Ovm2v9LEe7yD8Xi5bCNdiGZs9A+PP0/Z3JzYl6gW4db
gEHBkXgfSfgUxitipkNGrSE/CT5gwEPtTAMTsNTuzybf6bqV9kT8QnK+uBxP/zeKmfDJ1ukfRTuo
3CT9d5BAsweMRzfZRJM/TmNc5/+ZVlIQt5EYdgvuZ6ziCxKw6ne7wPpaZQAelz5TYtTzCnrxbp4J
7B7u1uFtN6YJjF3UaeIEaWx1kaYCQnVlAhpJYAlvMOiXzZHb9yhtlWpmLfHlGQxi+d9BCDumSCGn
6bNkjOcKmG4ykHWxu0eo8o5ITLG1Vj6ipoDgJe19VuY1o3C40owOisYcduC5SpkD1rsmSyc/CgoI
AxihOJnIKdIjZTk7NGLgo2fOmXiXJWUTBnexnrTdGPN9au1oLwCcf1FSPv3hy/4eGSkDyU5a7cs3
iQsIR/Ao25JSaoXFWtNX3hZfHEy944BHXXshIf7IyrIa8Y3fTgLaGklKOxC1j19LXhd69QPXxDRo
3sWUfSrBGTdkFOXarN6QF5Ujew8+6oOedKy2kBCAVZJyAwdL37jseELVSQgMrmB7mS3JOAEWPTfh
MT9TKkBljKwKMcfiYXAqvru3v0LdWOtY5Cy3s6bBAm0LjL+06d3n4P+pto8Ws4WcPgqw8c/zQ3n/
C85HbXFynAsA+pAyXL4WNJ0dZ6rDmZUdx5rT1S0clr6C1GYC+6uwvhgKWZuYJpd2XWbieUQ83jVG
t0cgy0ELFbbEE64HtXMnx1BFMnRLv+OjAJnK4J/nYOukPZdq8MRsS1U6eqXSL4bQQ9xFYXakp7vT
Gxqj0jzhrfaX+LPbARahI4yeWXiicjXXTE3lEAV9Bs7E/sPiFebjrk7AeeTChO+qNdptGsjEvfVX
3daMpCz9hjv4D6AO05AdUtxW6jM44sp0HcjvzKd+hcpxSXnLj5x+WbcMCUe7qKXcnV3Au6jo7SNW
+9Lyp1aIdkTezDZERYrr3aawWgDZYxsrRq3CbFaXp7o5AnNC/qSFBu1EQP2NMyVGhVkRLk8/9IHK
wr5sjigxMIVvi8meR4vNh/iYNbX6AqBZN+PHLvkYonaZ6HgudJ7VcykwtccBlm/ORvS0GG/nmL0X
6R0IDK5cQNVpc/C566VOiuz2UDgArzZqBfNwD1ZZeKcsVHo0YyRoABlcyHeaMYjnUPXLxOdIwpJ+
ucWPASH+7dmgN7FBc2hzLxtb1dN/KEzDuHFyNb6bnMnuFnmKhgu0j6S9nExX2SBAec4RxF2dGSHf
E0mRkxUhHFIdQHL05UugSzuLbHNA7LUduieYNnKyufLslcDoWzR4qjlk4gJpoMDfkVXyz6H/sKBl
+gTgIYrHmeB9aTy4x55WnqDB+WmFWbBzWiizIO566buiAmY25T91s/Nmf2JEwkH3cykQ/T6UthRl
z0txRFCGSuobx14q3GhFAGpBfrkIk8gW3AJC2aZ4p9TwJaiLfl1Bcf95BDSPeQMx2TowG4aERh1Z
X+8wglP6Z63pIqcQmFAn5eGmNfiGoky5gpYKxEyuTM5t6KzumZePH67nfSxV7KcdjZ9lQoNw5lPp
PDTI/35T5WlQntNrENiHIUZc+DwjAJeiMY0n/k42qpN9QUA84MXC9oSsKBxz2iVS0uThVEaAsu9F
FXVSFlRL9Ms2KEGnXUyWa6prosdGUX03P/oKjqcxXNZZk3d3x8SSFV0Xix6eA5r8MdtiXKtqznro
Wf9Zbklz8GPb3LiJ6EyoypTJ7sYe/mmFTPDXl0Gm2uJz/Wi304SO68Mpg1K+6ocNizlRP3d+Cq3m
BQadW8qvLTmb5p09O0ObtQ/zp109fw8ln5FRCmnP5YKsbL2dUhH3H199slctv4usuOd/0ZpXi9qv
LnmOQ723VbJsCLZ/gn3qs17cgmfZoglUVC+pVVkIrZuWvoeht4hTUt+PC4PjbSBnD9BWu/z63Qj4
+m4GxvD918+iixfOLDeH7gisv13Q8dZuBSYfgtXV66ros1x3/Y1N29/VeoEsCVSnt1opLW56KjdT
QPeb51g46crawrIwb+XLV4Kph+6Fz6/gNaW4p6bw0l5U0PMbF0TJKZE0r9Qj/ZBMLT4nT0juwW0H
F0TJSCT1WXPJ32sh8uajJICc0lOcxaJ/Ro3W5IrKtKmTZgiBTQXaYdxnJ8Ub2Qy2o4w3r7DHtONc
p56BRV8bBvEAToLwLUHHrb7xI56U2Gre00LDWFByIJsXK2hmhzlcqoL8MavpZEJLi3zbCH2mf3M9
zWzjxWwYzJzhGtsADGfoYoBGO8SU6mbu2sRSMP1dmisGC69O1KDVG6KO2np939F46MgBl8HZSj9d
cLXY3ivw3bO5HNbVoeD8GFYb88NqhxOi10w1U8xHzGAOdQcQSVJZHPfiMVgsC53drlKWfrzDN9Ek
2i9+T8fIljhsWwOQz9RmgpNXcQSNBQagT4smhDaPEZMoJtLS6IhGR8eO8n48UjR318vkvbSfKIXW
tfctsS5/Vu24VQkxppqSW50W00m+/hd/LMrvW2dnGNkeoznxmq+mYxEtE6PxXrVjtYMl3tUOCONE
ibvnUxtDmd3fwC7A7x0mZIZmFZwVi3HoO0Vrj6cckyv2KpnxoxRlc8b1BtDFe8yJ0le8iXBYDVrg
rVCxAQ/LL4ZlmRWG4LVzVOZkQJICJA0HCWE9Qd1AP4WTT+0titOejGEnc+RNn/e/pVp+eS6r5wZR
FCRASs1gRVatQTQBSxWvgQQPzGEuLyMDGfPzPcgMQN+fqQIKSf0hiOzXBfv9ypzF35TUx+kX6vzA
M/AEmKtZ5ls0F+TGYLMfy2EgcH3HtTqyrg7AmyRG49L+8BpH9ZmzLVsL3nLi9v1VK2SN5qlhKSyd
r5Xvq4ZxStaFbCKF5hD6CxZTU8g13q82+8B8zFDQwaphJ6+vs9mn06AQ2TQS8quEJjtZyEDX2wCI
MoXbdr64TobORflprQ3VKRxbMnDg9yVXh+RwUXjsUigFtM2b5VKvP/Pxs6BuFqX61w/bhEd1S5hw
SU0v6Nsfj0uIJpt3kU3nN+XKo5IvcgHWM8wGIMeqvRJsf96VKe+Ryzs89RqogMGIfvAqUD3Ne3LA
EQAIcXc5JPEifcUmfISmJojgDsi1C4f7Ww1ZxFk3ZWRhxGbRf+H92CvYCMaqwXXVeSYEk3uC8asS
xunbzd+VLtUW8D1EIIp74eoCmrUn993GbZ0Xtlt4VJRcl6iPEvORMA7ivlfHrzmLKu6mGVge2iva
LjgOiBaTGNj6wvGKVs/ld825E/x6IjabPwdIH/bWSjtvXrX6iF0RxYd86kSDZ9jBE4npM3M+38JZ
WsZ15QtQrOUE2eu6BvBvCIZhypEQsXWTlGaa1NQZrVH6/xHbhzN7a7FmQvZMDMKmixMty/uAlEAF
phpRQdymq9Nn2qWw65yHO2xDidQWSMaTZKrAFeBaTCHrXZMDKPrPA6bR2W70qoDsZR2vCxMCjY9J
Fdm0a1jThNvuiBhXuxVFAxjMAM/2vxhy/NfL/voxFCGfYnOywCpKOb/WS67YOCpPSyY9Sa6gKg5M
lij6AH5vs/LsQ/p7U8CKjv/m/DQn0fHeQh2B4ZGPM92loS5WGuFno3/dXFzhT+zUgAWhyFx27zdV
FBNTL3X7RzXukjL/gt5wvRR/2nOot8FT/JdU/GcSAva5jQECsIrgdRcBrVMHNe8NfVULfNpkuyTM
NrrwdlCjBhdNwZ86evLseuQvB1rev+hHlB2sxFTCUchVN8ZV4zzmfATYn1iZKdCFhPpVGnzlx3Iy
wKupgA8Dga96JHsVYCi18k8RVWAF1UCt2oRigjQKyTC6cGdV9K66aOMYikQC7gBGqT9GEvK8Yp2h
r2wc2sukSt42edUZ54sce/+5kjFknC9MHHV2lMNHhpA0A7xYa41tJbopjAkpmEb86L0/omxZOt1A
3yDGc4YkhsPpbN0u1fSh6m1qCOYz2IC5qYS4fDM/IwyiE860F5+mvpiCUazavqQtdy+QvNzDPEFd
r4lFr8dqg0KtFCh2mF+TV06ePKKoewduS5ky1gzsoY9FDsPH9z6/+GQANHH+oqSv4BJJQb5HwOJU
rpUW1Z1QIX1J6k1Itj4gAtJ89o28conq914+eJgEeSYOxRJB6ILrxOfSBJUNgrBnIc2UmvEs0G1/
ThrUiWUJhmbAma7lSKLd7xojH7pQ9MQdqeOlEFhUmsC1USEePRyq7bMbdQWAXbFhoMh/lp4hI5y9
Rn/BK8CWwaF261Mhvj4x7LHNbfGZZ/zMF0OpHwJYGdMl8s1Qt/0wbcxGYsC0W3iSN3beYxphbLRN
oRFKTsiQPh1IfRQOxglFZWe6Vv0eycgmlMoZNycj+s8+m27YFM+VsaKS1eRg7PMjPiTOX9yD1CMW
GRR6T/1lkFAsRVbwZNtfYP3uR1NA9wbSH7FNpZQmtCU9ptdYjW0r4Cwrkb2TeOYoOZwwvozRQ8oP
CtgV54jOOaFNvr2hEtFmaGHKXUqrVCgsxL+z10M6LXgPE3DxfBGu5f6yDtvwLpzGOOfEh4YzQXDu
k1MC0Pva2wolxzJDlz7RxVIjMIaE3iLM/rXp2tODaDIuCIoyQcbhBgFerxp36Ivyx4TlverOlKP1
Hzm+IqL6L0eWho75hfiFECL3zSvw+4OCCDLx4Aro4UfM7/wu0YsKdl6FMnkv8miboTuB7QEbMjPO
F0vhPtE54MTrtbIuQaH4sB8m9VQ1eId9w0P+YCAqDdvNlcrkcIjN7ekwQJX+0bYxV8wLl/a2H7Lx
R+vEhqg5ntt/b6hWl3rdgsmhiK5F9cixMSDUB3pjc4jpQf+DEe+1/JFdkd4avvqYws2G8NfXjk08
hHwS4HUAjLq1RbRAQQbjw4vWQ0kBl8ZEc91EpfEiDbTr5TB8JIe4BPAmePtFRBVVsKPUZFOSrO58
+rd9imIEoWBtykfXmugqjWqGIQgIhIPby4rujAP0bmJhAn5HDVlgBW3A6gA2ztwSUlEc//hQ+Gl7
SXqzTDG07WR0oJ4H8LrlaHMElz+ICIdrmr/zOy/FGOsCpMQsIPNNpPPLdKar68zWwVxOYu/x5iEx
D/XpB9UD7aR+JfHYAw+f5ZM/bpG73TPMrQJUhPN/Npv5PvcA7d6VGI1pWGnq7wCaAK3D+ZjmG7Sz
1+GuF3DILnjcAzkoNfLkVhoGdsOr8CaMcbFqeXVngRGMAQ/83mwGEY7TmIuM0eZXfssrHJnnJoy+
stAGUrJ8Qyqa6vmQ78Ik7iIo3oMeY1xnrdSFGsuubDM5JnkfT7wwUOqpQIEiA5J0qo5WpHY2nC5/
8suxXPsvlGju1lwr237y2p9bzh+PBM8hDAq6f1A+3a4oMRHYZpWwaDcX9BJQl8hOwS2SQnII1cC0
twIqifQdta2slhkVLdLOoqwO73C+psEMGc/Md3kQCxI+0JQpGA2Y3ISG0DJqbQwDAgoYp3Ob5BA5
/qX2yiaNRIQdEeKWxgHu+RoxLlYSkqj1aVM4z8NTicxtmiQzdBrYag9b3IUDJKJmu0Fujf8JPARZ
hmraZfauXllEwUL24iFnljUoYt9NA5aCaDmSK8ipncfNYJDK7idj34tD0/EZaA+55Jx0xd4gdf0f
wAtOyhx5mNBgvgGahB0OQy5X3UyTAV/MU0VnibQKJcDnWX+7EPZ7tTtLXvcpCRgPkzM9tKBxzpao
0i33yEDp+UvpEQHa0AXGgXP8iwX4B/30uJ0LzM5+iyivSd7AK9rVvPpTl8+hp36iMx4EoRA7UlxL
iUAHfLS/x+99sQjZcg3OT0mBiaApncCEpIJhLM4kCep8c7mB2s55biP1caJNz6SD/7wIhmrjkZsp
vbJwpaDYEsP+wRCa/MqDnG7wKwXfTb4CBBZqVP1GWm1983V+FK5oIyX5H4Cx/hwmLv8EwxYYasZu
Tep1apmXtIxXjzOVkJZnnwa9JHPobLPyV2oTdTlszr6jcorkwHSAvC2wjHwu/iTsYxik9Au3KvO9
skNp7m/hSb9ksaCXN5364VLDIn9SW3gQOMwVpiTctEaCXnXkmNnm7+h0dFqs7QY9cA7t7h2LS/YU
t21IAXhQN9qYF6P/1J5U/7LO8/yIlofKTmx1milQUA8KWCtxsyl1qApwMrJj4LXrbZRbJnlR3Ygy
qrmk1vxA14U861hLTE+qiuRiBkjBLt/V1pcj01jGOYVOXEj/RWbRyykPYNX75gPDxs6LY9MO+/Vq
NHPIxuQk7VSG19QEkHJo2ueoU7wuBgwcDE8Vbkvv+F6r1y4zyHH1hkpfYApz3ORwLi90a6Xvk3Uy
muH1fFNO0zChNi0L/wOmuM/MB17FpX17uHKgTJ8on4nmG4iNWWL55USvtUxKCZO4J8b/bX64Wnma
qqkvu8m7RfqYdZfJ3cvnUam2k63bWr6II6rjZZ/QsLWpjSiJvPL0pWWBtOZq7Knw2Un8ihbtylSz
r58DYz8yb9ghRvby2wZIm546lETsA/rVBQF1lUHSgiHEKNP+iA+dSN1OIMx8mb8L3IhJZ2muJvMv
6L/uewC1mTPXU0/bpM+Ni7mRd0NILujIlgpCwPF3EkR6HMPKQzvGBAkMQ/b9CYIu4jl4QoKQ4Q/6
OHyv1c1xLaDv3iE3r3mJWGTeQE6WG+p7Gzry2U2yrADMoXz2mIwjXKc36zgLkSIKtrbS8ju1g+uS
2CjSsaYc55Ae6UraGuIbZD7t6sUpM02s5ysl/1pOGyI0iIc9QK9Stdmc7WDHVfKSRhAVv+wzuzmJ
LfVt0PBrSzlLeC4Xzs0ll2FH1E0q7LbrpqQnNnZuVlP972hOx2WGCiYnvGFOPphtjleLNVU4FJmi
YEriI9CNhNDBc69QmlSU49u2FZXwexT2mFbMNmqtUqs8d0DgzxuO66+bCLS3EWTN4F1Qmz80sUbK
HSz4AeYgqRek2sUX7ZC1frYKnbwWkR02mZ3gU+aFG+SkDP1WORARy50EhVYVbRBz7elu3E+14o2b
hvLRDlo/SDOj0uAb4BboauRFxXjMinYZM6LqKvt9/cJ0kv2172XZm5dr7lRcSB3x1QT1p434JKgQ
tWccO6nl7cmuDycI+AexwrjYMzQ9jag+6Mc3U9fh2/NNQflLy7o8cmAQBQCEOzjMX/41TMjn6R+2
T7U97IlhX1Bn4wxjDUIgx+2vO+uMZeK9ECEQKg3NPR+5iaN7XPVQjDZ5V+CwXU9SY2UiAlnfSLLR
ADd2JQTfHcCmc3hEoUR2f3WyooIDHf6FgCzRncvSr6MyMqENyZTu//RXxSdR6jd8urRxlqWpILMr
l/HMpzgdDT6BfaeIofpreXOiTWKbWnP2+oanMK2CpQkZ4gdyi5vENB7iWntTMqAEjEN43kUuijIz
2wr66MdsIB2aybudUtJnh5JS90rWMAd238dJmfQ2UtInr+crXzU4yqdv9K9PFs6utw1fXmcuplki
eoRbZxCeb7IasvNX2ozGRhKseka3++iFyIqefjZYcB2luCleyJrryDSKxEwa6Ias87P2i6NZ4czv
3QGLXDRc3OuKBd2FI1/IBOHKm8aW3pZTSpn000XF6doNA9jU0HvMSWzDHLWCkD1z2ekEkt5FzhDl
2B0KIwrHwBpNEEqaSSkGwQ2yKzZGwWeKBiz81uIDdWtq8lpSEkNkXzgodSwoeGA2TxpaE8x0y4gs
tfNAlH4vYVEZ5/sulDM2Vw13nnM9fJIbbtM45uzBKg/yK3sDvlQSU9H9nnyShjLZdmWOSLqwl4qs
DkFTNoj8yyaTi8ciCf/DfGRUZKQOXIx/SI/n2dJzzCOj/U6OttHXDmbu7RtZSEowOgLSJY2ahV3y
seg9HYeVNsQKvx+6jzx0FlFyZVomk3//vtiXrO3JQll8KuU6ckRHu42PvYXhAQvJD+b+Vr/ors6S
/vj2mYJZP66vGcPZyDAoQxE4ckkBAE0504eeGQvKlaTIHWlpvpSyNaUZm3VnfQBujgMVCoshMIOO
EvNOOg0RMpc5qhmCzaN7FDASGiEqKTHg1n446+x/YbT1UJiqdLecM+F3SMJ97S86aUl/9y/ZfYFC
BzbmFcjYAEF6KX4zzaaWp+UYEaSYW+BNMMFpewFx2sNbLsSnEI87o9KfNCiaLv6Liwnwbu/KDAKX
kBeFfOn3pb7M+S2BdXs/IjTwBF1Ya3jrKgTExdYDRPQxIHWa7ZFqzV6Fg0/4Hp6iZv4ATrKwxcVc
jEkxwZm552moaDJi/62u5/d/gJnk61F1YlJ+XVO0Ft7MRoZYpwLcs8QrA/PHQyzCsuPho7+mM0Xj
I+IgROsXRhGlHZfqf8IP2TtR9XndyxbHXiUwRYf80Is8qXYOxWuT67QyzwwYQbKYiFCsOBQSN61Y
NQxmMLq5mILGNeqK74/lP4GmmZJony2CPPiStl9tD3PqBvfCR6cRRlKoaFslxu1KT/Mu9e1xvOYj
g/8Y48UWSze0EnkioQday2tdOl0MCzHhqZjOEK2d4NP9Y9nmY+2sBKNF59VBLpaWSCq1oT/ZpIrk
15MpeYi73ctWz1UJKciAiqHOm7aO2rz9Sczt83aDRF4y1YeGM5A1gTkkBZgIMRFbn6UYuXBFcXjh
hQN9NnlXMmL2RWZocy0lZw5eXDGawgeyzL5uyBXm/tlejhZ0DlHuRRPJ3kBHXSd9wo5mEG/mLSWZ
vv0omlClzrQQjC8zArMHUnHcRC8MrAOIpsQEJ/I0G0rPP1Em5RxOleva91Ogk8eVZSDHxct1l0ZY
fGwl/M22AGSVPTJr0yGsIZyIx0lRij8oREfMlzjwI/l5slKpL9L1cZVm+6rcG9OH94FJn0fe/Hhe
YV46XFqsGLCDCpkO4BchU/eeEykSYF1StClPyxLgBv4ZmgPmGYiyrL7eD/geKTY/PMAKe1tA9Ecf
TtJJmgBIhPaVxtQgpOA+h5mzK21IHVyVlzPgIeYvM7QHh9yPBVm00q0J/JBMPeeSkyrB+37wPF2Z
Yx8dpq6+hW7o4tVJ+EIQnsqPRBWXfo0ko4ZCfwBipxYbe6lHRuBHZ4vyS0031/r5i+CZwwqPSD/N
vGIVYxigWB8vDVYW+LoPBG7CMBxtHsxNzTAcl8VfWkI+opkcXbLHoGXKQzR16Hc/2JCLd6BqnNdA
6Af8LpSiAqerQvbbR0DTXGlz5Cr+HdIZNIGRB0kjoEuryTh2L3Z0uVGulbhF6+qqR+Abd2x+YF7Z
fXp4ckWgkjIq4OVwM9PmWxm8F1oYdci87TGOA99kQKqdNHRrbC+T6I6UExhPxjkAGhQLQ5FPkqbY
6E5cLifozT2wtAcTQPVHz6k3zk1wWO8/hTaty6gvRqTGLpCNIAVbwZ4bEt45nrDPMgze95vu/59Y
wAazIyVT6JV0RnHsiUZouyRcw9fxjSzkCSgP99XfgDMwmGXUuE5OUnfxSYPkPEbD7l0V7z6jGtxv
qpoMiNgyIo4hLTosANmdByC+dJeIHCLI2oxSHmjhwBp39g2JPfYplMGDv6YswKBudvGGU1W1lrcW
ppm9UM7mSe02JLTRh7a4ybBvL9L6al0xQwNFRuBY0nV7Vyd9l8gYaiBKR81NRcZl8725wyYV5mer
+CgGw4NdASqx5CAzy9K3TF0qdCdKIk2c+2UcHHuI13E6ZA5Y2xMGYZ/E09V2LfvCd3W1JXFFZaBY
MzmQzzlyU01gKEmCIeN6bFxESMYOeUP96BiWLs/Dufj9X/O7237HeFiM/DiQ1/wTHf9eh1Hw/JRs
7Q6fqy1kKx46DXjeoDV1JgPWwszhi04ySql6BBiqr1ZKpwNp9efaEmMK7OvIQvUuFV0Xl2RY58If
fKtVtumFpVyP86YsjOkmretUejvnWeoE4ixgbaq8wvkLAfnZk8rr56rcIEyfiwkQxQSIxS5u5ryk
bYj+/OchZUGSwq29nIgjDpUg4b5jazqsLAln37jJO6yOQRSWBEQQJSA6op1C0lMiMEGrFewdz0Oy
97/F5CqgnIz8I9w0+DEow6y3c8CRTQY0xuDplbwnar+6VgdsvWYPt04lLVQ4V0gQq+9IoKZgWO9X
e1eg72HZ4qF1aKG7QCj3UFkgPi5S76rI2mEZwoCNLqSJbNtLep9zjlhhwHYOW/0gWiruPi/8fiCk
Rg1YLyM/gufToWNtDIHkjdJo8YS9l26y4wvU+gtn76cE55m213NP7jYnjniPN2exNahD5Ft8nE+C
oAAGWq50wjlTlpfgwsvvxRcp5RAUWUV2XHQXeWTOuSw+0veDpleJYRp7+HHahHZ1o27TUg1MPt9G
zcaoaivleRT4lQk621UIUCrGE793FMhQ2W1sZTBEJsfLjIr02W0P0IGNaJZ8gEeLZa9D1n3QcDhw
3iEj/0B5JRplNGxLsaZeg5OPG73xm8HtD6Vh3LzjmWMO/DYnN1l89Qnc7FC7ewjU7rdjUXObNrUL
PBwQ1njYPt8bBU0+PXZVTAWMbxIzeLTsb2NzsIYEICInSj5NGf1xMkOwIZ7sAAMbhJGZsMeaG1h4
bH9y9uLN7AM0lGUuseacIeFOZ7VOHRQQ6HlTqnOFSe/UH81x+9l7jvCHEB/sVZeFPmPpiPOaPvTp
r88gv+3oJIbKJjHbRAaGlTXMnAFOLeKCZ2b8US3N84um2YItAQL9JW4hflmW9jk/OKXcjw5WjWLS
MMYOCPGbeWOkcWwssMUjiMU+P2Jgm/Z8eOKBtqSGL1B7TYZ0aOLQxHGeU4UUCE2WkDOw0bhmNQxd
SSHuDW4RBiesSDbQ/2e2QYQiGLi4Cqk2P/bzb7QC2iPQnrSB61MnICvaVtgA+Kb7BFrYdd5IYhbD
x0uMpoI1G+K/WeKq0i8/BxmEXMSnT9iIZkYkciDvUZ0rm++8S0wTu1aLsZ4vIsfK4lBuDIeXvdmA
CeyHocyzk7lX1JbPRM65ST9Tscn7n2VQJcjVANcuwtKwRdbO5uBFw9ArGzPpfPqBm8qXUlBZQ1RD
o1YdHvfLNJ1b9B3x+euEiwqqlgLGv6GogEjuO4GCk7GIPmPX4cypUIHVRJjpPoTRogmRC6BDevFF
fYamn4W85NaaPVdbn6yyBkfobYRi4MLN9DUInmBqu4GOVOIDXQD493k92dkA9WAq2d/Kz0fdvUkR
sqS/F7QnTW6Z1j6MOZKVUwK3xl7M58PAxKvzGaxppcEom6QU9gM4DLyxBMUTliqSN+2HT4wfjiDk
EGjzaVwADrS821iEIj1WNWZ0ucVmLUk2LuxWAcof7oX55FTGIlHLfhJa9hTc2qssSBV9u6rPdZHr
39MABUrIszDdbnHBdVYZWE/X5tSb9ujCZ2ItIAOWSKORx+EKcOy4VTqCHzGiSilDq3KMu6lcOwsl
tGDajZVv89eQPQXs57DPjSq4KbZmVajDYd5Jjs1rTo+U4GproifCUZ84D9u0pKXXfST4GVkpMQVx
5zjuyAcj0j7RtgJCP9krTGiKuBVXnHE+Qmjgccw4ioKZxNBbs8xU7lz1Fc4Ni5J9nTA7rSe/o5O0
QjFeAZWeE/gmxIC4OX/c8oOPA0FzvwOwIi7Y0+9sYWTMuEBKJHD2aM4kkKLY9UGN7tvF69X3iF23
28Ra1AcmQsKfnrKJo/fcxCOGfK/U8l4j0y+09ZCwXSafPlkV1dnTMe5wdKw9hJXnfYmUaj7KLVVB
voaDh3pw9DdKku4zGbOnPVer1CWfmjz+ZaqG0Xa7tMnLLf7vlhY85Te6Bw5LDJMHP88dIiN/gmw9
TCnrlBrOLOryCa6n7jSKyBbsw2dDc1iJwiJuF1zfc0VeUlAoglHaGddWzJBvioaEHlGaS5eZFnOU
r7OcAaHil9uMAC16hVvRCg+uUFTgL49NU/1ewagZ1pPK/bPGZCzgSm2kWVhAYBUtG0ec+S7Eag2G
blPvz8Z7f+9PPklSMhxtMxvs6fywfDgYgv3MJgh8aJiHo3gvmyZQfXTh2fj36yb//9rt6931XT79
rbmDYJhHIfEDCYTbJLWpjs/d45a8Oc9KrOLKekFoLTxLXKMEyOGZ0v2dcv9Vj+9nDBEPzXdQRqku
KV8oFJtsv1gR3k7MU49YkGc/5w/lbkc8kIN+zrtuXhTtOmwjrxmIV8Q0pkRxQHkSgx/djkPT+r0k
kDYIVjRZkKQzZDwQwyUPs9Fvyrr+/Rd65W/Ta7XRBH7EX31sPUgw9xXjmwCV+03OTnd7b7gM9c7l
HwB5JPvLZbjUTRqyf1WZ4Ztl4rRLJFPZKNvb+1Jk5mla3KvDsHPGQCCoGyHZQos8eDYt2DVRck2w
j2bw03geAMowsGjm+8cm1xRYypYmQV8FrZbNTlPE61+qbV271/NCQGqDfNazXcioNIMF0Nciift1
q72OCUUHOfPHJNcdlRS5b74SkklJ1EwbMD6PXMBfmf+Akpfw/5cDB+VKdFCQfrxEbX9/J6J9ZypS
LEMrJ5uc4BJkEVwrGhVMLOAvnx5hqRtYGkZFJnQsCZcsmkLqC+64WJdZYBJQybuDw/YmHWv2An0P
FkaIbCSShLjpWuaEtIzlHcnfWCcfHLZwk4X7IGXDozHL5MXMxEYiextEPdIPHip5iX2fxyKHDRFZ
X8rVqoj8x7bYwocjN5Uo2a1xQoG6aji1SU5St//zJhMYQIaGLpCKXxkHuOlptsnHQea7H2mVKPQk
VpEwAwlSuDgIhk9DzkEechseJwLle7OaLeqV/kRhKH4ee/a2tQNdw049xq3G5AzBpD/1KRHqYktQ
vK/E/2wUZC44qqn8d0f24SsVex6cpnq4TExq398uxAfVcsP12e/YzlSen3RqGVJXX5G6Mg5hFmiW
OvdZpJh1qDlbL8E8/jI9k0r9w+RcnoGSx75egBqgRVffd7QYndFXuZGjBOleyCELCmrB6ujbcqvC
w+jDwWZPxDC97L7YhaQPr4Hx87ZEBO5m0/qPogizw6PXbMh87etRV4x6KuVoGcVIuXCt7qosq5dK
Y2/DYEmXUuD2mXpO4e5Wukz4X/0ug3sfbEO/OruGE7dbDujJgYxWo1kykyxDvYvzCNHkOyXK8M8j
+gSgfxILSrSV8/sp14l3qK9QGgge1h7X1ZhejvgOxc5xJIvaSfvNQbBJAFZ1YgmNSro9ZhIYyskm
2sTilPosd+7DsqRShdqWegp/KfLDlneee2lX50TpYE3IKhhUHV8pNNfVEMHmTa9nnrfqiUJdZVTT
YqSmGolya8zxunieSOrzVmH5/s1GCjkNS5JMRkOjK2pryuuoHGRm1H25Ad4jYIUh8l+eiKDjFwOx
V/NUEPJH8CcezJ0VWGxHeXVuio/DlvGTwnw3lnegRSJNmV1Sr2GVB7gf7RSSVwDnWkG0r0gMlqDx
+CqbqhK5Zm92PkgM+yHC/jVtvjojv55Fmeqd5hsSV7W9Eyyb8hM63OR5CfwocOy+wMJdfN4WBgda
qHnqgu2+WSGwMqJAzB62HmKHU0soCQnWz7L0SgtB4+NaPWkrNbe706hQGLlhez9xB1ewrOW6nL1t
Btb1yNjYvt0o+Yz+jETHc7SFmjS0rfRwi2asIxugtwg4cMrz5ZExYzuowmtUULbEahjpBxsWuba6
s3Id0hh9xKYJ6wkdPS8uYFHloDJd2Nbs+lVUwfP/f61aMRHpqA+yNLBZf8CpZ4ge6I9fHj0BDcNV
uxxuvatnyeGT0ixFDDyTD6BW4mppjurWozlh+8WJSQH58qPxJ0IcK1wDQJB0Yq0bblYU0uhoRSTQ
//mjnOH4MYS0TXJDrvQAaJ8VdujbZOXsYuUrRG3UeORzyRAp8KmsN3S9HAQ6xUDbMrsUnQ0kfDnD
MhqrbdZvFLF4fH/Xs4/A6KGl1UUzB+a5OMMcu4JPoX5iOILrxUbabJUK0KXW1xaGSUVecgN78R5E
LbQxJlBdPMBDWGL9ed/oZJcjD+FKqbvQ2rSk1gVB/75TcuQAUraNGGeSjxbWxi2YPCfIb1/VZQF3
WXsbwJPOsSrAO6lxikV2Zi+rjw3IkQQtDy7Gmfou5XB4fSk7B2h4a9bjLa5282OTU2p3XEkP0wZK
Rzqth+DdEHe80XIj3EFy1cKb3KaXseKy790jN2IgwKlK9QXnXycHenwJvB9YUeBZ8I/2FpLiZSb6
5SQHcIarip5dEslQkCJl714kcBBTFkBY801R0GoqWfoG8hhSyZrKDmh+b8+Du1BgEy3147W+ZMB0
kcDLstIZD5bmZ/Rd/MOKRq148EcsXMihUNyONRQMCAqNk+OvV0fndj34+7phXE9V4Xj+sX2xMPJ3
bR9GkX7lOV4w+qrwmTPfY7notMsBGGfWQyNfkOakY1OPm+8C/2A580GvMb3ZRow5QggI+GI5VYj0
DIKTCSQoK83HU+fsdx4hYmPJyGo15p5DERthXascgB32X1Pgn6Riu9yAYZEYPWXNzcRvWXeArlL8
Nj3IT9pJOACKnd3nqc83ojhrWllNLGC9N5qzny2eQmmwj3heSOWeMVTR5v3KPJvceSYQn0dlKG++
CVEVjLmu2T0A4fY/HRNQ5xOkbdldcnuFlz2uER0caDmhD+UuJGWqBMH+07h38idO+SicBjYG3Y+K
K3k2ZXUfpquTPy6JBBxV3AsPSlDv4m4Y9sw6E0ejHM58szjzv89K8kPqdavm/xVLiL/2rjSX1+vq
WZZs1DSa3we+y+xw8ULQGrYknrGFmarFEjj80IQxYwl78/NttKgm96CSTMqwAD3+UnJm058RQlGT
oebX2sfJnzLuXtpJxS9nMPJm0GgDG3PJkP1NTUKi0x7AHut/g5KTqfOLTlkjMImHhOHBNZXA+eFQ
tH7m5Wyh+RHRsCvjSdnxnOTGzmObVLeMmX3Yp5KwBLfd5ujZQxukbgBLGkuLpYxMw5HUWZix7p0E
FFCyG9RTxTF2iR0x8c1JfynmiEyiUtWxH5qUsyKxMzBc27FGm6UmELgkQGQMmaWw6Z2uJWy1xvYO
/FIF7IqTt/JCGV/YObivuwtiRLpka6SeFDv/i39QkmdwXrP97ZbB4HJbkNDKUysELeXbw1NusGN1
OYHzgiuCJih7s/wxC4hgc9pGkhIO3wrsK7yzrmQbWz2apuPRQ5ai2gDA4lfyIubmJv4YreKCA4Bi
UesSPbHpUW2goIMML902+HK3naAfbObVUx+jNYg5Qt5uHlumFFOtTWdtSwxInZOzDUWCIDyDfzBa
+xcMSx7Ul9iJTQUK1kmHuiQDSF4s2eOV0xZZbSMjLsQ5Ct9zpVbFwmJmB++P1nGg2h5H49l92gij
8VIB6BLm5Ge9sp98RQ7/9N24AA7BVNBxQOYYiuxTKLr0DMRr+CvTZfl8SkO06CZH7/2ZjxG7GfWl
w7t5PKxPec/YMEkni5wcs0caApKghO1zHNcBBf2vffz+E9Tlhc5k76UqxElob5l6GbaUaq2up1dG
sLPWB8cAIv725r3qIIA0nG6nKy+V85/c/gpElU+Bzp/1dXhW+ymWyEX87UvTVwD4dulqLkBKQy3g
BDTiLWAxdb2wel9JguH/mcrsS2wK4Zcjiw63qWYxslTVuzFEGqrZL49j4lx9g5887iES/Kmu8o9F
iceuWXM4N56dIUCP78eGnDFl6PHaJxi3RaCXirnTBizkLljN0NXzCLzTRDJY5ud23mrlUYnJ369o
snYcEDylD+NQvQlexawxwvcWq4Pt57pct4CN0HwrXFOtok4bWW7Sbe0JU1za/SLz8unbpDNZe4WI
GxBXv0fjM//MJr6VKe9KsykqJjvc3hdiqewwIzqDYbR5yqcQJdSk8MvN/76kDkQ7PLy4HZY6Bzaa
WHkR/HEWSMDYNGNMOIFxOINehYm0bhldNEHk0IFrtR5shFHA16fe90mtpcJ4USGL6sQZesj/C3TU
Lff1wSWEnbojKMCsqD5gar7ZNQ6PHjkTpMScO4h4snRipDm4iolvfS6yPQdnt20zierOeVHDJsG9
1Uisdwn7d7d1h1R2gUDrDkHwIQp6030/s3p/yEHH9aHaYaYuQzC1qGDhHv+x6N/61jjD1yI2dLWw
ylOx8boKK2hIj8AauWoj1wyKg3j6A7da71H4IIgi0OyNboIBSFSCq+NliomSDtOuV8Od0+StVzby
xJw1IpPneLoK0uJJN96wcM7L+Sq8CoKOLAhd5KqWFv9CaqrmWtLZ6ICdBlGJ4JamG23pJ9IMAwMW
ne1euZF5+tOQqD8cnvvMwOvx2tcsAnJ1BImc/5XIimxHAOOMGEhIpyMB9W+VyIAUZ4WgJaIglwoi
aS16G4jBwhzuchrmXWK0b3iQgTImnEF4OkeIgjS7bLk9g6BI14vj/IRLr33grceRvkG0wXFOkNLW
GyG+3g/i5Q94PaVs8ZPL/67rz6m+vli2A/AUCUp2ZOxjo3o9Lr/sdAQQO51o29fxmD7Wkc8HW8Cn
kYlPFzMMokJgpQ7+ZC2iQpqLq5wWOzBk7LK8Hr7eg9hPClKKxxb2CgnBQR3nPFdNR6+h4vVZpDwa
vBQfTrm1u3797WG81BgSTVw9/nsLTk9qfQqqeEMxB6X+ioDW9arrG28FaELBFtH8VlCCOGZcCBbS
T5EbJxfzJ4l4rn14tuo9uLzMJvhKa5zOgyIRTj1HcpHbaoVoXBI5UMb2TmDxXqzySng7cIsp5cP3
b1U2Pi4lc0V3zO6qZpFKAzaMlEBwkCPJM1rAwtvQuxwq+d02KkRgdqT5upmwPo2qs+6Yf4dI9U6Q
F9bgdGDkKrcCl+QK+/KW2UdeHFMud4PpLiMImUUIyYEwPbJ8xerWOUQITWr1OrXyGdltdH0xrh/g
8GuylkSf0HEHRGk6ysXZeyazjG7BgdPCea1AdRxwRSuVKJfs6TXWNoK+OobT134uA/SM8L4q+64d
J/ZZFaPqufcLggQdAn58qLjvsuio5mHic1yrqj86Mo1ARfC7uHgzfpCNUtTZe3Hi5h7rUiFrZ/Lc
xyIUQ4JnYH2qIQ6VeDaR9pkbjn2wMfJgB86ESSE/fqSTHvcxfPQZufQo9qkW4jXmevpbD62qWlBa
qgaucytGgwbDWka66DBro7Z3CIFRfDTW3530vT4t54FzJAXZ7wUohxfyrDWWEzHzB7ppk8mJnML3
NGGG3KdYNpPetbliRodphWXJF4fsut1enSeOhb43ZH8iYqQFBmnGsaLbErLPcqpKSs2pOco4hV/l
ssQmfs4Ot6vco0+rSpUOoW2Sbfq7atXyICFPuXicyxYt5Gff2OUbkqf4s5YkpvZ8MX2LdvRI3NLG
1Ox2ONhE6CocDwa2heTIXatoNJBowiHYno0qwlc/PoOvWAFBP4GAQwZeyvS42aGGL08+ei1zx4wS
96JAgc5Dh8bmQf5YbFT+vO01eoMbeKAP7ODIlwTmL/eg9y/pVAC2/0yqFuS4PHtdftIrZ/M1GgxS
hJHwKgz5tHg/lCya8uhr6r7Q1xgf5f7DV6vilwbEapl3hUmv6wUkmhezbJ07z53+PF0640oncmoR
ZUTnpEidoWm4ccfmsxfJeN5zwr2LA514vQkiehVCjsialtoQBasu/50VcIlo5d8ppdL4Escu+c4k
bus79o5CTQWwPo9Gkg9Sts7BmhtXOb5nFAda8RjXV0ZW8tp0K54l+EPnTZbYTE9+N/+uQZYNo2f4
i3QR2S1iIsls2bRXGrJmQUxTffFRDIs7sLkh+1KyLVnRDYMaLAjZd73TyYrNuZMTWCVhtLVy+jzs
mu8IR1LrqjSYJAkDyDXmmc27rtpmj0UM0oLAJ69EKFX71xRA93qIuenAPqDtCtZZJoRjovb+/A4Y
k7qNsnjPoBMX0nzIbofbaB4XBxr4voPaYrN4LdzBeqW6hOJS1CGaTq1zWjZgcziwwUdLV3hFE10z
zL1RoyNZHxpjtPbi48s9atLx33ExbzfUSH/mNYKpq+P/NFuC8hS8Y0Z/OT41KhyrVbN2yU55jL0j
D2zYR7O7/rGeNjFtASd/5UL03UfqT6TOZYkt3NB3K6eiP5AJ2lhPFnSGFmjxQCS4jwYioFGnoDpN
LyZiORTncMQD1AXifg69r15H6rULS+uz2sxJ4CgAyT4wbYiOyeM7KDBNbWM20jqYj6F+VNzSWGkl
P7qpDiyEiTdheUIlDAOwt1rVDVgOdgqwYGr7EabIi/ZzQT6goXY89c6xF9d/w8OuYfxy3iJ02fh+
YWMQ8j2chdsOpXEOVX6REQMDmrXNdkADKo1XDoA3/C16CMntSvmGDYVzyivKh7IIZrItGtsUFmr8
dKbaFwXcd40KKnbXaeucxgIAQz650+UloXsIjy7tq/Vl+vc8+UhKvT0kyxLhjbOkPPxANmlpYR38
xb6keW7fF3gIuO7X0Gw2QhbfFe9UULjJ+jRho18S1GC+n6c+qG7yKeZhhBrsmgKv3FtIACgG/aV0
Tqc/IVYBiOC57gn0J2khxzMC7xx4ddLMIEkvU3sTiT3gob/STYGntMUWqAKlONiU6SIitWQPJBcy
/G+9of3Isy++v0A+4g3dgsUk4w3nL34SfQ3w7wnew6nSuuM4uMEr74WmlX9TTkYoZPcWmn1KF19R
CPDVa2Q4X872knuUcmSwkUJtrMJGFGAd8R8O/fYxZ9w1kkNUDAQ+M1OBvdp44hxkRZuihw79usIE
ff+J2rHiDdYCRMbOJxVmTHrEcaeuHhx6iAr2vZxFKudGeusrAx1VDfsLlK3TqV3BR7J1cAVP6fW3
DtRCeGODovJQddyOXkYVx3gB0XrRgUMZWeYxWgCv8W5dAqBuwaWRmTFOC0hqzXgz0Fy2cXxm3eHx
b2H1hGbnjnDTN3TaWjkcKD1d+eDilDGyKZQjyBTcNin/YkAOP2AdG/LJ5QtbgP0Lgrwr0rjbz80s
E+m+mG1qSS0r6rlOz3aEmbhHSSFM2ysJ7qeuxf3KyXE4ePu3TR00IE8ENDtEClpdUnU6iTxbOodi
vuKDJzQPCy863+fPuH9XWEjGk+VBNTcwC74zIt2O0PPXD7Ic6HhmZTHKcaq1I3ySFYdsGS6PDzIp
YWbX3keZ3oAnsZh92KnVU+BdIsR0BJxW6vbOdRYX0KRpQ/+966UA8EgeNmfr83ODCv4Zoy1GnvFF
MtDIQkNVSg9D7LZk62Leu+Ezh0RWv67Fth0VPBIc0VV38poU3GFfcHXBLkD5IguHdnn8GOxPimA1
XJlhpFxqrOiN5vpW50gBHADTSuYFS0nwhvCMXqITQYtgK4HfbcrwD1HIGmA4Dsx9gO09vBlR0TJ+
ygSFxe82ToO5n1hVJ+lQcHUQNVz9AxhhQfHSxi/nSzdZZEsicnO2cmo/H8ERnhjmExIGm815NR7P
iZFzzRMe2G5RpKIbci1HkpB6IjxUgf7IDWYD8gxAA7PJv9GOOmuugZQ/T9No/cvb1InrSLTdaD3A
czsXya5b+DzKfcpe6iAYdwqwkgMJaWjGlIrq00vhgxT9WIeuDdApStuPS6LNLCrvYmKEKKXV02sD
hCeXTIrjYYTLMuelf/t87el8ZgDEr49mQpBe3sMyjtj2M3rMRCnGpCnAXbkA7tS//dCs4KTJkSOQ
ZAHeGEvnwkemLpeqifY0hSF9+8JGXJgXDHQ0QwZqZLVdQgnKVGOc5k0kZk7a6hNHh4B1G8ef1hgo
JhkxCeGCpGv/SY3XLS51JVBkBBbSmRVFu2G3iejZJnHZoZoC2h0jTT36fXa+gUJK+ddlYhneecA3
sY0DTzaR/NtriIN9+mSmj7B59/z3H1/HQHY56TC04t5ExvU/eVedpXvFCuB7YEclFPb7WlwxHW7F
BQ6Vz9MsVwuglezwWkFL5my+y+Z/MrzNGHdQgosM/knbkMV3ZwXbiKDGOUcNElxArV5kZALzfK7E
ili+Sq8wwipqGYrNGbZ8TD0mC7OTdVE5JfQdmH+xpJ+EjhS6FvZjeE+L8R1vN+mt1qyQPiQNAZeS
h/k1EHF8BBDEUNoGzfRK0GcAF+Kj9mgzmnMvagKNej80st5mX8p+TSUoNaBCBOKK3tT3JT/yP4wa
nxnxnLQlS/5IwtKzvet8q9BXWn3mBxG+JaZJ3e6vYRxgPvcRiPt68ly4AmHqszZMnpIAaVapXx2l
JnxBSR8Esdp2ucjPNTsoorVKT9xfiMWEGRvpHJBga82GoUdZi9T/dFBNZmMAsfFl6B8Ds0YJGG6E
AxiIXb0jded2asK+2kTlMTTeblmm0/AZbKnlbfRTF/DV6Ff61NnmixkBV5KRNlBrw85tBryXvYJp
lU2ktJ2skLK1ygOPN7qkedd52XwcQJlPAZArbRKtBkmYsPZ7qIksMMGe5K0Dv3sbG6qrkF9NLcJF
2Q9XotuY/M9iM0Z/iznsz20VPRasHVuVLi0WJMbhVuW+No9DKRHbyvqZ6k3s8zPrnQ5ZRKwL6PfE
Fe+bqDfB5iFbhsyBA5JU+qgFonKIPCgy1ShGyPepEoTyIaakwJH7r2D9RV+Sy85Ys8iBdgQAKA4W
s8VXRUWuaxlJL89FSAr0AzhZpL8md9r0kuMoKwEunDbvD36ESl1EUvMIfA353IHPrdIinynlwrUS
ZQEQPVRrvuL2cfkliBUEouNzOyJLid8RyzhojLiKd7WSgPnMt4ZviR+AB21ohCvHc++yiDh404R0
SHSFlZOsgxZVktZRQGwEUPuBwWt0c0Aa0qYYljQJrL7rXn4jeBH3jVn2TCFGB06sMAOF3b0s2yTi
Rubqm5S2+odSrmV9hhxpxmC7zlRXqsMwOQkScDFWRghKeLlhKPRuyU/E/AKn3Rf9YtDQjHhCkb9z
AYlvOj3nuHc3waKOdwVWpv9iS+VnssQ/xebREfzc5uAiwRrWsxPNJDS7G9QI7WGQQuaHXfExduxn
fSmSXpkhPsgslgJrSgOROWJRIaAHNDE5yVPxn9EwbG8nCg65SvJ9QLpjzi2YAxnGcWqfrS182UXx
GUBYf0Wc3VCgY65nvcAlaIt0ZD/yJMyVNt9JwJhtcT50luu9ux3J0i1GxdvGELdTFwqXe/rYI+Ow
zjhYyflZ9ILGDRC4MnhzvWtwoKK5p+mEXq64CzBeknUGxDY6aBAqgmDtruOqHDigxbGdS/Uy1JHW
FcN1JGUc+WI8oUdmVXKxArJRFu0KwmRljeIsYvsMtAuz/OYkmkWuKybG5pLEfeAb8T/AoaMRZTc4
jISFwIETWHD4O6moahj9ugCZd/ax8w+AUlcuXGX95BPAGjmGOQhtd5IuhHlV+YzUauFJxaTYeWM8
9J5Sb6+tcfEEr48s1fwbUD1fcdcF2YS5cUGCToS7RouRF6TQyxsC2/6HIgWcnlSEqjGGKWe6bWEX
dkyvOWp4fOKOrEeYwbgy1pEYlv8T+NYW+Ywfm8VEm3NO2OWX410zUVB8YAkWFDc3EJMy408Qc9/2
PwUhb1RaYLzhDa6y2Wz2sWMN1fryeVwF8j/YCx0e3gOfUMoVv8DGDdzzUPC+5y/5wA0Dh3AyoU8y
1tX++EHpzkwfmp6UF0fsZnNNMLgggmh9ScJzbFwQ6sM1fM55BfEfBQtU0Pvo6vUKRHGyz36wKqfJ
l/07OQWfnRnUxDsEgcXQr6QIr/cM77P3l+BfLhQaVQh5c9xA0TiV46SOEhkRSOdt7XyYhkC18Dd+
AWGgejAcYqlIu2IRfrMaaNG/IVi/CH2Bt4D0g+5gcjkQQxlPJkzeoF+dsT8MbdvkXrjP3Bo7KCv9
0O8vUke3S77XyuiS1E1I8UZqstSoq/l0uydlvdzBm6qmDyINu0osn6lSBKxZwtFLhNv/R+zMKO23
yhQAHDG2aZrsMK2lrCCH8JUPDQFWChpgeXb4goq5aiOEkStJsacj/2hpfZ0mhNvczbNiRSf8jNwS
/ozFFMUNAS+o3m/1KPPEDtUD8W+iwPIs5hOHO8riDuML7EtjEGeCSTXvkHnh6xmJNNwL3CQ5Htvq
AFU3naasVZ0sEzYHmBBKtc5GarzcCkDcOvkdphjPzb7+cpfxwnSY8N3gvSao+04VuzTnbhhgJHVN
9doYZQO60ck8FG7nqIxA3Bt084Xv5oKF58U/a182bKt9+wm5hS99t/ozciGgmpjLqz8KFUftx0e1
bfK/gZs498zSBEkuC6aNkXMsFPLO0V9Em6grXw453+FuRal8/qhG4HeC5ega2aAirHpNRPdWkKMX
+s15i+23wBGLUecYLsu3Wz/u58jsTDECBAqWlX2UUTYsSCQhekiSXfcHZui6CTgSGm8SnWbxWryb
IebC4qXcZeFxr7Vna7mn7DkDQ5hs01UvF6MP3mq2qSYdfdJvy7i8GyeDEt6Fsoryz/EHgkpWSRzE
36VaiyJDRoc3ecRnFFM1YjnWFS+CD2yZQVuOLeMSyXGYEeFECsn8WWebC6jtXL0rSP4F/9ZYlCdM
YhHw36LKN0QRcYAPpMaLOikX2r1YntUxJhcuHhFzzzxdcMhX3uGG5LxFJElFMhlvBNKYpZPX/A/i
XFkdII4f07Uzal0akZorIsnHnL44lSp9TyPTDTaLwv0qwGn19SDvdpru7mN2lmdqsT8a0BZD+yat
GsHX6npfuu3zdCUMLMjKJSuHcwYTLVEjFj3nuuIQpTjQuorKgBB+YIz505e+SQpU8wyg9CHIAMSz
CGs3c6Y9Mrcp0pdpmcTKk7ye6RFygUmW5YNHT4hPlL3Ey2TM26p0444JZ/Vvv6YycM6sOqE5jrhK
9KcNxQbtyI7ZwcRohdRFZuQdarELo/zbiTY4VLwTMg0gW0dQ8Gos77Ov5x9azjaNOiuuri36DWmn
zTOaJz+V/D+o/0WuDLzcfO06g2liDI5WLHWuXu5bAVdwsDpDP7rmr9mdWT53yXNqSLv4f1kzYVqv
sCqWWkBVfZlUf2Sc8b6gjkLRUji/7kwLYNvSUTrkogaIgpp7iajkSmjmTIUK/7P2zdPR47HEB+Z0
9q8povLJrzAnnd5txaAavSSjNTS20J1bQByrhK8QYbaMvcMd25gIsmjm4RS8IqkFOhdXTpKQIR64
E4tuXhN+JAMTKZpZaJ3AwADM/X11dasZnBYvV0ka0eZ151AyuvFG6aCzAFvzOXVkSFvbW/tUnadj
qDXBnHh/DMHid+mdXqFi3bbPt03Usm39oGqZo1g8pVxlKeQD6NIkNubA6cyA+bOmI6p3CP9pi/1J
SOFSrrqCLwiyWiVEcGoejJwOIgVWd99p7biz2NVFvR+PIY+7R2v8/b8CXZDK/0SpYO/dkRUBHC1l
81FegeeYyXmodsSAcJ0qD9aAwiZJPtlR6A9N2LkSSCQu2PVnUX+46GNhS5q99tRZSNJel9mYeLFS
FToHHzn9SDq32Z6BXUPZQaGPqtXYfDluu1+1JuFmYbiI2IjrwJblWzQk5l6Nus3q0ITIZpACwUss
/5xoHdNl4mpgbRHguIytx4HWthrjOfxZ2BH8ItqsCHRIlkJrHlyCSOtQAM2/359oNIy0/A4hKcvT
2t7S9YBQga3pA8po7WFvrw4zwfS+12zsjZHxj9fZYOAdDeAZtS7QlXE5KUhXvi+u0k99k10uWMhF
HYAyhXolu+f6iKg20bXYP3cTv9AT+z/mOH5pig0o1HBv+MN0T4n1MggLIH+Gwv2NiUGLjBObIsmw
xtFEtq5xCpUYlcd+7zOBv7zvJHdy5wv1zUZ/DzCE8NcemE536WTf+Ck9utJF384S/tOXHQqry4+Y
5sF/E+ikCbuUGBv6kKRrbV4ElJ+XVouLgNpmHncRSMmujrje6X8FGCMe+bcv7W4L6rQfwbllLD2q
eSAqTIikARAc9pqD+5ac8AWu/UX4ToX1EWAelZQCe7OAfO5M5sKJ5NaJ4EkdySEBnwB7Mt6sUquT
eRD8ej92W+LuEp1IMXrQKl8U/M4LhQSkYK/XkCOqH1KWj6wC7WKiLbQTH9h12jnIG6LsvthXi7ho
j4/vpLYHhi5i/uUjHGHyC8O9vZ9UvKYFlFTzMYOY3oNrk+OZQSLHoGT6yAV6eB/lZV97nxF4452K
volxQVRm1wKh5Ebv57vl8VTgsECxjxF306LFVDiIMjLLgiAD7h/Tauyu2ru2MLPhiUFVzE8DkSDf
34032TMDZglNWtcRyW4mhaaCKtBI3/5NFn9MJbCq5DDwioXPNqGicjuhWk5uTVxO0o1b8393XGaw
bcUOJGqVc26vqs5kESAumGEqiQZB4l3QrJg6K0opm4EFrBmCMdHxLCQBTU5f1K8G8qy9cSU3ZCkg
48tu5ZrxZUGVC0ZBX6gCVp2irs35O4HvoA6yiS0JPOSB5+UgHlzV4hJYka3c42oNahavwJmtzHsA
XMXh1ADCn9gWSwiIPW2MUeuQyqb8Jm79+FVn34Jowopxtj4uQ9V4q9XWyT1ezhYNANahB1pVl4Bx
RiDd4PWNs69Rc4rRcEprkgub2JOAXMcquWbVJDErit7Qy35u6BNiLKnNozQcIE6/JMCbjC3klLZ/
qzndoNeI5zSHfVkh95I4Y8OjBCD3/JGjqO//ObM9lN7PnkZoTtAGSbSneDV/CFxoB2kiRpZUTDP5
sfVDQweK6v5UZ/BIO4B7x36Qa8Uj6JDSpMd7+YVO+1FpWbhpyU2/irZdzF4IamD5DRncMbsFhDnn
0BTspm3X0W7980NfvEmcXYZMQ7TF6V1dXgbyjrhasdN2JJomALnTGTO381086pvB4qOq/x/N+hVY
xj1tPlMITokh6epyB5DufCaJguQWb1yBxoBmwzwbq6+JHN2AlBuhMYJ5DtYRWV2ZOKLoDc0D0en4
XpomBl3V/Om3rZE+ThblQXjgrk/u6XqleeITYP8PIqbQC0sykRoItgSIrVTI2ITfCZ7rCHxZqWaN
oIS2nhoWoFTNj2CdnB3kyY8Z36jGVbjqTd/8EMv7MlWwu3LqJvUOeboNuG9JEQeDrflO7xeS6YaZ
XtUf2GMkICzc64Hfo5fab7oMwrirl4ipIqG2+VxnP1bRh0QYnMJ6lgCahkNUDc5NKwmsnSFdIfvm
hKRcFKbsWnk73+cR1Iy9D3SLpirdxFK+edIPWVeWD3Ujc1Vjljv46MCY0YdXBKKIZ8IEMp8EqDUI
CsphOX8rNbQ1KvgtZqu64xoPDb/oxi3bbhRwVnGPGURkUWyoFBL3iWAqRd4hZ9L7hIts7DytCA4a
nIIIVcgHCsD4w82nNeDz2cdpQF3tIHmiw91KL4zu63cGdoeeDPHOne0RGn5FfDXYM4gueMOyIp7Z
sB496+MMWDmm0XZPGAhwAjBkCKaB/FjIjr/5HMC+XugOGSUVIMTRDvTWNqpkKCM2NkX56m/EG1Nj
7njeUmf2NBAiotF+lKO2/lLTg4zM8r2+mv2PXuiFWezinD5sZQRH4JzcogsqmorjYnxsqyOJGZC8
rUwHfFEyMNjpXACurIZlja1Huj2J6Vq/qmzn/9AYlWtCaKQzfi4XFOQYpAtdvYMfxroJWUf1gMtI
Dww9eDmlxmuzaPt/mmpkfbIJjx3QpBRga2ZjpH2D0mKG1vLb1fb1LQrRo8oTpOY/xPFHx9syJd+X
7mqXd/MN1AkGHrvHzIP21azBOQtlDd/vVqrwSAxODTfLNidFPY8Evyq14WiR2BJXqhd4RwvoOBnE
uRFhJqiqnsmVWSsXBtfSdsyEltf30NcwsAgEr1DgDFKfNlT+tzi7IkXyWdLFgpopD0MhQlm2IrRR
yVUaezSJF7y4WLqcqfqaSM36Jepn9xEhzyouXD7DzN3RnCZCLvJEePlR9jze5S1kh3dSHWwyMv9R
XQqSDScozHq+6a6BxrP26XJddzIvppXwYyk9NP10v4LGc3a0derYX4rjSJLBL2Gsmu1xBc63KiPI
JQ+OWm5oWirgCxvujpDzfTryWS5czhlGBTODyaIg3vpLOe5UYhkQj40NalHMJqcGDM72xqOK044n
S8g8RYC4jMuYtrOMOGJVly1OTRtBdjGa2+3ayEiGeuVhjmYH84J4l/aJ/VrEA+fYwDyh+zmvLTQa
VixWkvgdLcygsdM9WmrssuUq4S47LopoMKcZ6KTC4s7L4WMuWnICyqOXusB2NiWbcSpeocBe+0pn
fmwq7cQE4374lLKNE1C+X6X2vHHjXNyVPYdCB6VVoeUh3c7S0qixAIQ+iypxCxIWF8KulR2W3dEh
YrS1cFzMuMaxE1QRTZjBdV9Mkj20HQ6SfSROK5qJNGcPaeSEE0Z7xXsxPQ+Wd+qZL1E4aRRO2tog
nWrjyZkJ/diM2AaAG2kU0TEpmg6rth6DmbifvL1Y01hCNYnejztZBhs2w1yTsgaJ7qrc4Slm7yoL
QtO6g93xdUupLtS/Zi/ZKFlBz4t84Fr1vBgiEuisYeld3gn4jVLuLqtWujJNQuwcZXsrDbSr4pFn
LSC9zCFAeHenMZKe/iwcVtPSMO35i+IuusXJarPm/lKSWtoKPElsIWAkTLK+fMsc9gxNtjovD+nI
uvLxYDSddhm2LVwqFHaxcZbvdZF+HNDpJI4mbj8FKBb/TkG82o0d1vB6pqEbLXWvSThFq/LEphoT
NxLWmkrB6QsTCUql5mlX0yhCMjsW9N6U1Wrm+KzFa+XDBegfjo7wn8dV/IhTX3wyK11E0uZPyQaq
ZPgm307QFN5OgBDvp+cQBbkBeYiXFlsMwlrWfyxwlU8wvmx1rkMk0TlM6LXCwAyaNvXF1L96ixro
dCBoPxvM1n0fM6YPY9MRLGiqpAMJfq37efGGUOh/4XcKLM0rh8cgKvCh20VIKdQO/BnzgQrQHgou
wVvpBkPO4qlZDaGmU2+pI/tW1TyEtJdfmrIe0m2oN1LyCIVOolEn2456BIw2mWzeK7sbFFMLeezT
j42ODQ/eGQFCZ4CitJyvaQy2TtpXRYwZy7IX0hbBQoN2466oyHJRh+8ERs+mcq1Xsp/8pXTYhHI1
yH+4QjgLemBS9UnfIGGV3s+Bni3G5VilW959nEnl97XfoFGfYSlH0tIURVJGLh6JpnY7Afk9CYy7
eUUZaiWxtuCduvgk/poLIYZgoswIsHM7uEAFByDrqRWtWvQeZXck3lly/1tyBF3M+OPoGii0DNr5
5vbd1zduD9gmVNgDYxQKxYZvkNAkUry7UYba9jMhkd/AqGUL0vCwgNtMKu4aWqpw6G1tBTzzP71g
GrgmentGO0eVDay/srDHL96+J1KRtiXGWHlc7rk/grJK/yX9V08qMekpLT61RGEadwDddNfE/2/m
zBBhKchhJBDIxw0gJ5W0E8FFvkpL9KKViKV+YvssYrAPFTLIGqUZiC/lmLBCFBt/Dly7Z0sKgw3D
4LMff4vAtA2sQ98AGeKc+OdBT9kylGIJHm+bwcDssuT54HJAhMux8bztTQ3dwqy0YumnhvbNrCeV
AaxyrlvXg+l/8xrw+f9H/paKhFQD+S4Nj/0Y5pHDyfENyM9aaU+fkgXY/DOG5jMQap3HNHEXXiBo
ivFUG0l8/mSMiE9mO6a0nahWGJ8+SMar32RRs0z7gRPphE0LfOBBURCI3tHNaS9JrgMcAN528Php
RJZWCqVRYjeHGh4hSeNmuU242YXQB59nlNYN8EWVghXSpfG8713f7j4muSZnm5XXaLrM3Yswd54a
//BnXK3+kZ8wN+LOW2lncCezbNJbNwUzCcqT37apF1logr+K9gKrdcdb3ZcAZaLJV8cE4+AsMqc0
FxpuIZMQXctUhxoFfeTb4gRjz9FW2N53n8NjlkstR8jtxD+nlhs3WEC1DRMxuWqOwGhlaE2Hs5O2
QOvNbXU8pr0P1/80/GIdLMMWoQhLRdNtXzpewrcqUfCZI+XbLRF12eElBXWgU4ug4Zq0O3Z0vLiT
ZQYiRBkASuVRAB1JfLaqyfEqr8DlmBunXx2OFqAzqGVlb3fk1ipUvmtZNyIEgrmypB6nYXmj9XRb
eU0HyuX5rhSYxAy5VUnOJ4VfqpOGAcoGdN0r+vTrxMMES9Ntz/udl8Tpc1Y/oceU9rdG8u8VuzoF
ZRMc+9yTy4U9JOC37lUVFmKaMiWhSTsOqWfpBtzc0WoqfwmPNXrEVFSxGI4EbiitqAHvQviUNBfe
8ngFgJgSSdp8FG600TxKQFxAT4fDZ4tUN7untVtMz7qge95HnQHGT1H4YUsd/fgn7vDLn+Z6Zo4F
swW0/pRpqZKz/akBlclJc/GfYni81+uGdo/pIIXUtRWR0ONPhKZENRS0MXuLtOT+TSwrxA/Y8Osh
imVtU8R/9q01kPnpiYp+bBIb/F5YimRBu+bKi3OCbn7zYjx2rEAHovYyF0HIdWtF7FtfbVa7b3tW
vQNqqi+yeIe0o0bj4HQbBJkuFRs1bWiztyaN4bk6BcAeyMHUr4FEgbUP+pL6771kRPIwyTvVO20K
b59U1GqCRqPm4htwOoV/mnkw3nARaUv0knJPXsveB2RxyvvuB18BOv/qjJj4n+RWD5tKOb3MDEgU
GioDPgVUGoxaTZ/6i6P1aO/nXrWIlf0ceaUBjXkbEMIy8Fh75zK830EusKYyhi5f1I42hv9Hd6qL
vvNm7J9jmMdEouk1ZDzvdBA6Ix7HABQMkjuectrdPdDcRZA+6oJdJNLmueX504D/hZ47XxjfLINk
0jf7Q11N+BmSzjp1kaNLO28/V1IZ4rS2QQPCGF+lfHNgdQgW2bhfe1eZE2PCqdH9Zfq6CBJu5XvS
V6qRUR6c3Uo4JTffIR1znzaZKDf7BsPoUoAWM3Fj4FjyLcIRnR97GDgnL55VeC0/udc8EEjbPF0m
Wrs6zKGdHRRoYR4cpa0L2IGxmm1Pa1NgOZcWzrtrZ0Z+cwAMSt+65UOAQ+Of+1lOM66BARwwD+62
PIkY05dIxLmbKbXl36aJ5TUwALy1VRrL0yDHz7+qgC4rt4l9/2wezQyKtDdRv0hDwWbSF2RxK6ee
OE/y4y+FNZ6lDEKCW3OLvtG72tn2SL+K36RvPqFx1sSI5AJMqOuBChDa03xjefKVaLGxExy7Mv9L
oXUVz6Bn0x5HbdSbGTaYhBKDG/1/0hGU4P2jZ7g5AxKt6BRddECfckp3BwwRn/boBZUe14mh+hm8
hf5p5noYU1w10DMM1gQwNhdRe06nFiYczQtQ1JMG7cu0RYDl5f7riz6IYO1ovuox1nXMGw/1Mlxq
yXYyxLHxjOQGXNwE1uNPMOc7Awd417Smci8Lo1RyE5+jQgYSVdPVsMMbf3txZIKAN0z7y9i+wm87
y/q0cQ+TZxzRaCiZxmCng44fvcJzdwzGvii7dZwjj1p3lR/3bwbIdsmGqMlLbOjCbAic7loXGGRy
YVWCDRJ1VZkihceQHqJTSPWDGuQ/F0Q15bnCiXUcGYsIAPJ+wkwF5SMtn8GAkQ4t1TxgUObn3qJL
kGcayzg3oQW0+91fBPU33EhpIxp4J9jb8p5vjX2hWizzDTbSpfLUGZMcPdKahvDb9QJ/nuzPtNOB
pdi1n+uWzOdCTKjTSdqHORPsADtBdsl3lEr+v5OU4cs5qPxyMmJlWJn6yYmSVmxSxfU0Ev4Uh5xh
95k5G4SfCKkP/qP4hXFSx1mzUysoS/IjZ4P3IBcx6z2ivkYThYaXxUJaXW+qtbC1ZQO+CG5uc7sp
J0tqJN/FXjiTqPPqEpXbaVu4b/XOFC7ZMgiEiPToLiyB4uBGWve1HmvodFUiE2tY1czFm1hT79LD
Zb3ha3YaIbpwtVy0SzlE7qR9gAMD+DUOfE7VXTh0O++mXGjlRCcO4u/vNIM7D7nd0qCpyx+056dR
hKVY0VSJvo7abTwrGvZrS2J1X3JJv3TKJDvfO3hNqYXAz6Qw7QAm0Ej1WErfvLtVrTr59+oTTWs5
xGHxfP4LIZy+lznvfNNZBIEGnwE0gmriblw2AoROEI9BVbdavkaPa+HxUNYPYT/VhkQvaOE5ZXjn
KpzcCbKG38UarwdeYlXS2frmG1qRCaNOYZdLE+oeYyPXv1vkbUJ5QUUPs6vj5nR06RfixgJ8mujB
sBRIftBLEaaO6ApcRdLHRS9UR88ZXcJse0lkrAND4GFCfla/xleeqdmMZZAVFH7pZAYXsrk2VZCR
rkE9UMUgCcwZuMonHduzSZkj8yb8zs3Psk3PX7E0Jr8fgBClkCAKjDAfjgWsT4srzGeQvbsyBo6G
6fQrotsESfHlOrlCTVnefa76nKjdZEPO6boZmSFQCNHrkmtmdtesQuz6s+PWDPY+H+a41DMfUwqQ
k95ECKw/oGwGFUPypiMtGlVJo8FqCeX2lHaJnwAJm2crghEwPN/RL/iTn0oIwipAR9/0A0MK8WbR
1Ib9RsAfF44tkn2eeIEx9C7zG0Ml2g52gF3tymV9bWVnbympV8wls9M/I1uSaMy7RrkCmfDn0n3e
oe3hUMzIlPbBjzdn8X8Z/uBvdoD/nzRyiq7iqgVBD1rgODsazZMC1rrtU4F4aCQoO1ZMJLwRaCgu
ZSDCEU1lawk7rkSq5n7N+vQh5lHoh0ZilkxgdJ94qnmLmlMGRLUUVZuyKTL8HMj8mL72ln63uw9j
YdaeTLB7xIjMN6SIbVBEUYPfYmeaFtYXUJ4/zJkXw2E5ST9DF2TB4iVvWv6aPzibSL12ue9vvkXT
yuT7d5zPDeU+qwucGdNknvvv2lPMr0byeykxGMiHetlCu2v9oB9cV9A90DwfEjIWB/2quFsFC3H6
uvWlqAKSjbRqLcsxhEXyCgqjqXynqdsWu2IO0OJOgHa2FcH/+vrJl0+ARS50gfxv8VxjH9y6Zq6k
ktBzm7aYpwIG2D9Ba6Vv4C1hWUMblWp+l5uhvoVAX6+shZwoleYbDrTg+6lBzjaFZn7kmzaZzNnt
Hn2Wsr7XnCGF1WZZEZHjMRcB9JwnND+YsQgPF9167Dh22OBGRl+PLeVMl3d+B0RaZDZdxHsqVzFt
SJtJuSUVdiIjKs2IL5p9hyoMDyoZESrO72IwJMTUg3lI0XsGqVeMpqlKvOm8sUaaOK4Q0OeUr9Yq
NZEmd1CC4p1COSmQOEsjYXkhFkC8SCRSDPpArpNoX8eUKmRKBUM/kCuyQNuPsAeS5W6gPvI0OtvB
VT612whoDT/jA0PBuCDuFwIO6W+n9poAeupSGcGoSnkclsY75iGroQ24ya+sqUvHsHGd7odKKp/d
rEJx8DRs1UbP3OFbK36DNOU2dPDnFQO3Xxs7KmwPAPWNuhtdPMWQArp3/LwNcJTwZFfSZS9e8EI8
C7amgW0E7FjbJbZcZH+0tXWt5MI97jC1KRKZ0HvY1LTRQaJz/ahdSR40RzzdIRtyKZmi5iwatd9k
OmpmGFpPzhpLSNPcVJSHi+dAMQkh/+Ps9kHvVgMdn+K+4kTbrqmUtCC9CpqqRoWOtIHKxAoi8Jue
4H09f/SndSrAM5jUJOkpu8JV/xN8JGW/gzpH1+JdVH9bJonlL+JDbVgyfdZ5likg8Mmiuj3015zY
M0o1tEKUbOZ5OWxYfWaQF/WUdUZkIzQVEBCIPGQi+n7Q+EasUUe06yvN/JngZwWDqKR5w2Q96+ag
oTktyIi5woWEzQ+vlFNDmr5YXUQfu/aB6xEcjIdgMLzPnp1n8OhKW2LwGBmXHV1+9nFZvi0pl0OR
49BJJVAJVJBgszFojP5x2TrOAT3Wb2RCtozGQsOipT9rHfnjSiaZ006KCyrEV5TTpJe9fNYXfOHq
kV9Ih5pyjaZY7slEs80Mp43egmFR14mR9Rfdh8W6YvSk5QEImyvXPhhETFhn/mrjIHqdXTJeEq36
4VT4AlSE5HbzeanGFNstaQIouVAspSYh3vUfoNiuCAxdYqnAYEMQvwcwdUENR2ZWygFLUA/4o8fO
EQ8Sqw+SyEa6YyH0wYH+0pJ2deVvBsDhJTXUaDBavj4vxIBsPQ0NDHdGgCamxqxnHEVDFp8oij8O
ZLFGCQ1YPq2mHfk2TENH9X8ohgWPLUaIeVBp52l579a3tzwZ9qoNGRgrCKZ8fJlIWuXhygTeNkYG
Ydci5pW+udOe9E2tK6Crriwjdk9v3KD5R9CEsobL+YKBr3IDzuMbhgb4cen74PIucHM1xpQoSGJb
v8cs1xcMwN+mc1Swfa/f+a0I7BsEbN04w3bYoXFtwDvTp82HcQqwcivahOly/FAr2vX1DEsLy6nK
r9/5w0/WcgKPVJgOEh2pB0XcpMcAI28raVSbbiowkEH3e6HIydW7/gyscmM6hzJWdoL/R3SHZ1CL
7bmD9EkoIaNyeBXoaCLiTXOh1QfuJaFGOFU1nCtlMDP0Msxu9x5ub5r0zHzUvCt3W6nWyZ/5WUe/
yLaTFag5K33DG5R7LWsjuKN5eNHn5P1ojPM4hzYrExEg+OYU9Yph+2TmdvaJnHEgg5IQVOq5eHeO
P69ccpUvrnNaRZyfZAQg4NsIvL9idNwYFoxqdAuChWohfY71MIr3nnX1ivqmBaRz/NkED8HgkUoX
JW4zMUwrGWiK4tpYCvQUFQ+zL4O+41kdup1dxSHiY7dTl5FoepiB0y0n1g5oD3Qf9uXLlTgde2fv
zxlQ3YUhIeBGA9HFINEBck5ylm+YjktvuROWwgErYUfXEhxE3+xaFx/mQk0ZjYWyolmm0X5I8SSN
6tAVlGJLIY3u5pgKOOaSiuGNHdD1hjya0e5+rXpevBM+7HdK6gfJ1W6NAkEluLSAhEaSekq7S4XV
ONDfcxNBDynCj5zEgPJ0jQaliVPSCfovXbggIk/ui4neb3Mjj4Yq1fl08nNbFTc6/rhTOJoPeVrz
uMu3uP+YTP3OwYBS7lKAo3t7EYCdvs3eNoZYFJ85AzFvXaESDgVnqDCcfNRw9BMH8ixbGV0rxFDc
kG02xgd9596yctO0XrJGvC2tqcvk28NlPfn0I1+6/mtVLXTrZ7DzHbb4zTw9W1gFBR0e1xCwZaAP
IcuCM4/u6J66o4bCcbSDkpduq0DTIrRva5J4NIWsvE8CNHN4eaByYKyjg+vcMa0sRSMAAaFkGiLm
SB9bh8EVR8pI3JvYlxCBDSjdaxobZzBTAM/YnuTVMPVUnWCT7iiWqz62O239jrTT/5NdbzYp+Amf
PeWWQBnNmwHugpivGO8eaFvJA68thyDR24QjSQKmjPL+HUFu6xEj3XBQ0kOwRmn6O5PrVFqB501N
qPtnwv962EnFeKXLRUnhaWDKrGlz8TtGB1GWX0+7LJ5ENyj6LRIUL4HfnyC6ndz1wijNomiz1LRW
LS8kHjMC2MNtKPhqzt9PivCmSTDI8RvA1e1cqm7Jj824pBq6gYwb5Y9QHKPwWv33GuTDFGO8w2Jw
xy3llUw3qq8G6ZHqXlhbbo4yqDl9cxlsUzy1DAbpRqGjHdBC6G/MD1LGhPAURXaLWcXLI5C/g89p
HghSyYYR1udmyW0KYIMnXS9O2xsNvJZAxr/RmISy6zwAbQAQ+4uPZnre9cX9Z5m640JyXRSpDou/
ZVUK5EGd+SviaXBEgKQVLX40WAcOP2nY7qznzzFJ9Erig71kes0an6DUd5YgHrg7LqsdbPylrSMC
fwitT0hfGh3aHq/pPgCvuX3TLf5wx5Y9AjX3FBXACUITL8fgpFSG5JekzTzghiT3gg3035R9aODz
DC4HagEx/SVp+OU6lx2VH74nuwguSue6wXc1w4mT5+MC03cA+zF/T9lZCBqUEfLb6vylifI0dZQA
stP4OfgJqXcKgs05mHtgr8H72fndc94OHXTkdieSPqZ92rcusoq+FuvsuJo+SuDa/tC5aVtBoP4q
rrSqg1tZycksC5PLISBzB2i8nFPIjuOabZpwkyhSVpDhmAGYz7PzcR5/UQbkO952vrfvg50+HNL0
noO5OQ3lTpoB1N1CTvH2sBXRKnJWpz97YV5AJAIPVpiZjk8VMRzq8JeyeinpZNlnFQC0I2/9rVfD
PPUJDCiSXKpWmaYta+2QnSNEvrNcfONT7HoSEbIQ/r4JfnX0MEY5FOewAoJQSBdwcqG0SarTFpGY
e7Q7Aq5g3z2ui2E6Cfp61202qOaOuI4RloQY2W+SKG1/VihMC5W3p2F4MjIt8eZvCfWZHF3wbW6L
9Lx9agGQ43a/+4bf4YU/1P7malmdyyirK+Px4UXLwRS5sZylhI8OsjawVmQULuv0GvhICopkW9wb
PFYFT65pf1TKq4l7fX5eOEy/hgmKq6pvGbEbdmXFkk4JHyfLTBsD5BqsDrqzdOZ0rCOiRrNi78zr
MlCY5yNJ8oNOGEoqM0LsKIqWHALB8KmTIQyTjCUthRj6FWd4B8tZlKeOk8CiJLTg6TQCBzUgv9P+
zWfAOqTSwho00wK2LkjsDeYxtSLaFXMaiiUl/VgW55x+rgNp/xzgI5sHMqi5WSktmHrAhMUkoJnq
pzcqHnqhqNz9L+CuA/rWtLUgSHweuDJxsBJtgrXbSC2C62OkaJ2AJHoLa89iVSemrlQomZC9gpMn
kiux2lsxRCvbGNY9O43fOilZhwRXDMXzoWi2MHc4SsMuHhDM/9Q2wh+oUsAayqn1cDLgX2tb/F25
rVb9qnk4JVnEGPa9+veCjwxHdht10+wzv4Y2AiM2n29tVPN3uG6sAzCUiKnk/sr/tZA35RnaILIt
aiZqGhz6irE6+PKY40g2/yQYPV04EQCXcQMIprZEbz67vsivDcvBCom6U9tqYlAoGOWp69lem/d/
0lb2dkl5ztNlcNVMEIKw9E4FBCHkZAUqCp3uglf2LLO8ZmsPAEwAFV5Dc8V0ceOzqePSb+w96QAs
6glGPTa1hxu2/OTHu8z2QuA6Hf5hExqVBPM+BDtZpCKifILNvMLW9AMouduqghvZD5M+TFF1w1P+
3EyUcPpHvBX3Yo1Yh3aXckKRx8r7JbX/dhCLA8fBPZNTEUCtPhd40NUbZbxGdY88oa5s2o6ueJ3q
JDHNzcbFtPk3h3V+7ubOEPM2krI4GoxqLSfNsoefjVHfVIYm32BqgrCT7AaCfLRkBGRFkLsVFOHf
gWz6K6Z/Vn455TsVF0Xte+K7rcbjnx5Lfr1D5w9js7rlc6NBC52Y+qURE8FJD1A+rZ/ivCO4oGqJ
UMUeSlc7RADLFxhB7GDvgLh+VgPMSQlPwwb2mz9KzyBXQ4vFTY/Izb7RfhP0FuJw5eIK9EZ0vSlF
FH6hJhvaVnWqm0KzmUwGKVRVGlhpxsjRQCVbs5d2S+s4fwQL0Q0fTKwLRGhsBwdOZkDMq5ieNxUt
OKlK68M8zliy3gIUHnPCRXdcw6HGkRkjBAxdc5rDJb7XU19v3J3fBeQAuCN0z6j20zsjQb+oDECC
iQlkLlheHKsyqIecwZuXa7T3VibeNP/fuVsXoAV+DFMBVgDiNv/q24ARhXX2Xb9abV16IRM1WprR
iJQ9Bmr1xdhbDPkMunQ2zHCCJYQUyMp4dfh/Ir5inETc4wmG5t0FbNReCA79HSv8gQ8PI6XIHMDz
WiFErkKyxJHcz6YVTNCSR+gh4dZe0ln5j8dVEhdvUnvNGZO+NhHCBABwbmpfePD8+uCfQXY15aEC
CenJI49GvR76cxUnbGKuIFBPOBO50VS1P+BxFoA6H8lPgYhFy5vxMrymCG/WT6/aAJ3s6FFYc/bY
Gi1TqyC8qex0yZpLnEIBoJlTKZMtLf7+a7QyeLoCD49jRD9K2j9Hhba1w9FlleTA64urmdPhyUJK
vIx2T2+4U0n2RGRcD8/IfB48B5YZbk934tBE02UavqUmxq3HdDZjM3+f6zvfdy9bFTyN7hrDHo0r
7dSFtRMJAirgWgz2pj6a7Etvg1fyBCm27ibOsEmkcKUts22gwNR4hFUZTpgevwn4FhrAz/iaCzxh
rmscTyiVnMipG8+CnQrPGTUz6h7mjpkQoriN0uTtm6ucnL7BeZAA7eajjX1JEGXkp0Y1PJlgMgZu
zNeVlx9YsF4OU4psm1rmPsNlP+1QIeZAfYAQBVaXOhAHI2XS7L3U4y/dduPbeuWUotqFlQTlK+tR
CTdpDGDrh/gGLUQ7kahBgrXk+glV7QIO7JYFQ7xV6BJeD6QY0sRYW+lVxpiIZ7CD+ZVmMXX5C2Jb
VPM+v9OfM1Jsk5OZD0E0IzIy33yZvAblwQClpCDTCEfjyBH+zalQNtRjPsOmNMI1aApUnMZKYq41
mnt7BTFQThhha32x49mJTs9zTnStIxu0K6jhHnjgPsLu6hZxr2MpPve/1l2F+dLkCYNlKnVakkJh
A7mE72xKHwPfPINk9+Hk865diTx810uLqomX+1ytYEW2sX+3TXKeYUHLJGP2oNRVxiSVFeMVnlgz
vMuXZjJW1NlpEwoQJPTiGNDo5AamghOk/PvyqRHZkyRvqtLkNmvnu74m+MqqPeT+cwEYKF48IqwD
wJkVEoyttVyJ8Fisb8phMPat8P0SZWMEt9sm04LEg8b7YqTpj5hPtEw5v+ESyFh3ymaTVcQiNj+u
y6CTIU0INOrTK+bhPQ3aHvnd+DXZnVSF97glA6sMvXNVML99a82ScrHr9AXJI2bLYXT8PgQ6Q0mh
X7FbeMH26CJGF/qyH6svVUyIRugnjiErdfGJEERrR89o5wQ3fX8gIXKWOKeEag0HATu23NO4DJMn
/hSaI3V/pb4pqd4c9/G9TR7P1FIm8z0GYiAKHq3Pj5tLEfV0Y6aepFudbDyGDlIsYCG+4i8QEDwf
YtMfHi0lebAidjNLZtaToifu+TVHx/sNIJ3mu2bEEazr+lvvH5eo6QUaZWMWfgik94yz6loAimJk
1XJ0A3lbG043+wZj3IVTSEzrzk3DFaFmH8zyB4Du9DlBlkeGS7sbmpoQLq3eLCf8cgmLjlQ0IWFU
hZtbkD9qaIKeVtbn7LYspUv1TH+lxTEucKf2Z1m7AdKTElk95eHE7UcUBv6mKGjUHvMJ4Xr+CUEB
tGpPyt9kqWVkRzrURVdyoeA1eoNbyjHbsGCMKuYW5oaM77ydo/FBm0WRR2UCtmRdDgQrOgOh6EhQ
pZ0F0Efdm9FC6vKapIPxBMTu3NXRt4R8BPzhULqS5sqX9ZQEJV3T+wJL509MBx76GN57BYgqxWiL
O1YHNQlnvMxe/DkAi0NXLLuJzVmpIiWwA9NsDPtxC7wEoS8yN2BShvyfGvC5INVsXxkKMq1pskaJ
LHRMpkSANbyZoG2o4WnLvqoC42Smm652sDTRDUl3Ny3thM1zd9DmPapVXfFC9/+g0fcOcZBLxhlh
yKEBPPGLmNhdnSlA8dxWNi4jrJv+sMcoMfryTYk2xxYt3eXv+kLenLHmVWTni7ZRx8Npxp8l2yj3
bGGmyJbLkBSfT+wA/xI9qm4Ma/pHY1F/KPT4gEzi4RTlaxcnpvGNexDQogbfaaHHY+sLV5vusIGi
gIOtIT6KaPg7toFSQnJDD/LSfQvKO4/aIKeXJGv86aCBROFSQeOVa41Cdt0UvZdHO4JMgJ860Uet
rI3eFvY6sSFdFvQtOtrkFB3XWGRdCjRnajrW3RRTVeou+/RXYXRgmQtfxuz0rOv/d9aBgqvo7BfL
KrOF+PmyVOIEBXlwn3QF/zoaS2OT5h6PtEArVJieaP5V9t151S8XcLMeLZA2SNAEW8CVTIzwiITX
8Ri6aNA1U9Y9F8QRAgwGgETZ/uF/32NajwZ88JXCiQOQ+D7cTC1OoL8CqB6wXYUwyUYT2qzP1qZE
+29seuAy6lzgAydFeuI/iLiSf99WAdg9IEj0RKZpAZZRvTKquVTaRCE4wLS1/VcJcH2ATXhByPJZ
Ex04uTWdlNmHlRyzsfJ9CNpkYsMJ0Zx/o+Roxu9P6YuUb/z4tmXcdjt+3PTD0zVcWc08OF0eBSVe
aWA2k7CtVzxbhmKKzfxwQjLWaqlTciiq4sGKd0SI9JSAa0DonpDav01XLyFRTBUA2UpynUcjQ49P
0KpY5kXHWxJxYEegcwvSOQwXPM83ZDhlOyQ1eQZK89wb8bRF1QF4wY44ALuBS4Hf7aCbfKY/gvGI
7iaWlQB8XQomkkDIcPK7LiuvDq0ZCgqMlCZSDN8DkeOFaC7ajGXYpkc/ZH2OIapM1ywND3Wwuxyg
JCywS6bQiw1zWkydkxRdtaNwdpEABcl6ojxBYKKHFMkup/c3+h8GRZngtc7Ou/Og17gJklcpkiBR
O7BIbsfen9Js0T1V9wZZhJQ7nDvpq90AG526UXMj1E5V6Sgk5jDSFCSmcbx56E0MOhHYFiN0qOTS
d5ftxGjQDcxhf3o+xCUAnRurPR4o9B0d/R5CfjSfBet2DuavN9XGnnUZeJUsejk2MZ21a+WGyMa8
a/X32Gxql9YcSi0r6iZzgl/taM79CVG8ZyElUgm0nxbhsvKhczJmbyWxnBvv2UBMqe1SpvLmBOZE
QQSABxN7sqfn5KGOh3Iwg/FtaJ31Xs2RW7+0uB5+gTXzAYhdNVzlHWMhjzeA1scEg8fLIv5CHIzE
tdLbnzoCQwzW8UQP0fl2sYOWaAmKaNgD0jayD0I76pRWmhe3KDlW63zTfS/LAekQ25V4TGY7TC12
NFq1ZfjYnSBdxCxwBLmLCgQAkcjrVHvipjrxNgdBE4poMPNyGgre9bPLBzYM6i6iWgg42Sm5QG3Z
E71WHv/L/Haus6cwbrl8IBfyxYh0E38HWus0CVpMXyToDt9HWP92w6+vHStO0NGqDtrI1Rv+8YJX
/QZ7kzLjmJvMAgNh2UIIZXEDy/8KC4i2fyMeyrE1vb5kTKOyl8TEIW52LlkREeD/x+KTwJqBxaCC
QP9WGxyLvNVU63l7EwhJ9DrUEZpLfPG1FPAm0XbpNQI9gXCDa1+DhZqN4iI4CVq2zzNPxigZhVsw
6MOwgV7n8nqUEgqARA8Qy9zhQq2XuQPy2Ri00L7rAZmRywkoziX7ghkVNajUOOxzYZ/vKXhUTIVJ
inlCWCQryDX7vQv0sksaifXzC+PHW3PRVO8UH+HP1UmCTkfvf/w2OIKktNiGNXiVKFtHczU6v8tR
nA96l+vxFDcui0B11hmamVOtqDiglJsferSHwGlVXNGs7/dgBcjbHXmBV1QfqfqsZfhE9WEIlLcS
nPkSRFlaj3sG+8it4JObMFcRE2A5HU/eO910vwVu1m+GMIdBbVLXsYq7jxtRhBwOYXq6+b4tcQDG
pEiZGcSEyhj7vYJviZGqJkrCdrEUFr7F3++CX3LMpSrqorHikIzKFBq2WZUS2v9/PU/ru4fHjqXO
5elCrAr1MJep1+QoRCGLj24e433YN8Ynvy0RqIJv++vYTZIqBEDCL04ntJ7eqkNTBQ7R2Hs93jEN
cd6N9eNfUAJShCTE4VevJ6ft0mK4Q8AluDwlLZxWV95rm5gCf6PLxA1rjobjAXBeXPEHETgmYN1c
Qn9cN6RD1XNswYghvwUK+c4XrofRyA2dW8weaX9Pt+oL/iO8gxBX1HQGo8mQZ9YY2OPWcPQNDOFZ
YYCdTb8eG92aEFZfe7SLzmyVwaWxbzHGaNgOD7/1TbVP0EjOCbJWhnlmRdghyz0qYr5+YnQWtFx4
iy09DFKB5jj0kpCGltXNVXKrnN7XAiUBRwd+DXO9rU9juQ3TMPe4QfWTEuv2ZghvScn7T3X+DUYx
FKWwinXP52vXf+8Y4D7CU0TYtkk9NHnLmxITP4zGeuFLW+KqGCl6Yy8q4GQF13Kshv7l6V1QS4LY
zh1lyz+Is++qAvt3aZ4/xBJZutGwRdbRAweaQdLjYFKzfmbzbDpp0tbapqGsOGqQMhmTcbF/XFN4
V9OPvR3HKt2v8v4TfLBMPXjaU8V4ghVVh6g8uSgOR7aXMKKdMDUdlzbfE/a1IWOWJXHjRI8xuPC+
1aWqqwXwCwTra3VYJ1vqjXBDyUUfhnLSN+qnC8yVrj0npWKX7FNre+hnigff5yyDuSlblH7DX2pn
yIe9hETcgUnMD7XAuFuy3iSnNRi32v2kiIprZ3m6gZs02wDoCMxS1MQvkSLt3fNoiqKK2kdKKfHw
Yu6PkVNu9cdoGW7H6HGvZB/wfZep2oYUshr8XCGe7TVx2ybagsrQlUERmbHyYjq153TzSxpyRbzj
/mIXPhBVpNNvgEJrPPj9CcGqQOrLFLLX1F4CNO06SfOSRO5kVNesJDdPkA0BEU9S6D/GYIg/0BJb
t69ZxYYkhA+K5Hh/SwFOFjbjxinKnjtRHFsaS0mFtxIbtaN/JEMLgLV66x4C6oaeg7excd/fAZ2e
E2lupfyYGlS+zSlPnHvVkRn5j4c2REjKmfswxF4SRusMh4hj/QzfRoHkG6gaD/UIv6CJpIFMwLEy
juCia3l2aMGyGBt7e2qdHZRLoAC9U2fr6XZq3TYyPJPhEo1Ib3U70ty2Xs7qglpfzdKQ56p1Fybq
CmJplWDZTkGyfMlXcQ3jtLwhZV32l7/PcQY/UCEJdGjyncbdHm4xFxv43/Prl75KesVu6ZqPoPsy
rMAs0NdeyJC0yzmUcYrFnHTiw2/GgdVZCJSXpQcc8ZLzp6s3YRN3w615Afgpd0XyP3ikLpQEkuLo
Gh3t9zRpp50daavibwaEU3pDlkce8F3MAtCOosOgHNL6hM4acDDgcDQmxjKIygKAhQcK3uFm6J4I
F7WiAPMZU5ml0FEyqXkydzVXQmaV5n1RxJMOxgVAtE5/28wjmUd0xIf6GV6QfOGJXn6q8poHsL+I
jB1zbRMrSXxsgUYHpVGxT7KuCV6epkcEbnCeeyFsOwzUbPP+DZAh1LVqGUQb1GH2Y4jutCz15rEW
JKSHsSG6tDJc852R/y0NAD+YSD/T1R/2V2SNrjRbMe0loJYkcjYkHJgCJzIpE0MlnxRoQhAr4gDt
P70CLVIlGC0vhhzUTssVUf8O2jSJtgBU04S7MOPEmQWlx5sa+8rvqrBEFcJbOnS7K2FUAM3y4adZ
SH7YbbMU6lMD7RPRgdZTkuzXm91fr1+MzvijlU+MkwdrEosMVmba8c0qSnernmJI/igQq15Rk7RT
Vve+SkNNLBmDoqJlhm8bqnKflDp62Nr/ixSwQaFmYWR9kQ+7xOsqu+HXNQActE+HA0rnfNmA1be/
/DzZaEu3kCa9iUpSljAPL8k4OORyaPFzXpAGSfvxJRW6I4UR0UtX9jW4seGuaVPgy8EYzAZC/lzX
Rrnm6ganmHMytt94g46nMu8WjI4OMkQ6Eh0iXt/xFOcitUyqtL8Bw15AQ+u9fUAeDIQ/gb6O6DQw
TSj4TpOiQFnp3og1uVdh2alyr5zrHVMg/G//Zfx2+P6OGM9kq73L1f2B7mzrVG4dFleUULdzYkSx
oWEvGT5+x4Jgj/2KGyH4Th+6PbGgSWvDRKJHgwgCEB8zE8rIp779G1AeZr9InLwtB9NvWdLuSmZo
nmS1zqZxWBbhTCGiCRGhCx30i2RIU+/WXuecTv+oEi8QA3y9okbYLD6VVqy35Bp7H+xSUAGUYaX6
LGSuXpqJodD+J0ApPvpmVCxThqyPNepEQhpP+JMeln4kR2ib4htE4HVb4zVO7T6u5DE5PJI2t/BU
8efyl5PMv3QjULKQUSjDEqN1uZmrUBAWpwHvvy8r9/5R6c9pWI5wJvU9YDHjYGih2jdgQ5KRF8Kv
IRyqZ2sy5afFX9pZzguvHtsThTJT0rP+Ez/att2SPjjgCl2sC+MgK/2mob8/aAuUKzZuF9RXGhFI
LN6ENP5bZIw0MU4OILtwc8I9UIJl8QNTbgsr9eoX/WCtYmEyDZENDUjmqcNxKg/q1DTuQxzIATNK
eRcp6Qa7vUuo5CGjDe5QtRsMmzzVv0nlCRfR7QjNvL/CWUWYafEHJqjGvhAfgKpvxg3QSNsz/IdX
5jb2YPhOxE6+LfzPlDVm6hxZwjP/2wY20UIpSeZftO7wXpmfqaiz0hKoD/3cDA3qMrGsuWuWtKgn
Vcd4sXR2bFX7e0MGH0XA7YAZxIZOEB5ccEEV7ru1+P1ctdf9cPSBIU5gWeyaoSH9cXzu3ax5lYcZ
sai0nEW1w6NgoRNU06Fzc5mhzf+caBTOwpWUL+4QF7JvxIMrAtuCj34ODo68x4SEgUymjFkYFVKT
AOZ1RnV8XkUsysjuBP2/sM/punWLNgXOi9azpOMhIKFkFfNWTp7qjg+nImtiPLO6ZleW9QwVXEyM
xp8Or6H+FkBmqWPvi6qJWhlXkc2pVuToFnDJ3glDaPnaJt3BgzJz7fKsnGkf4v5hmBQCxP8To5kG
KCzkgPamkhQ35lgFGxA+xnSOroCeiR8MXrJrx/uxyeqLuBewUxTMbxdxGVTvqwYf8r0/yWFYBohd
Yl01KG/g7J3CEsP0KFh6csTsjIPVwB6DMey9Ra5qXAZZycwA1xyOJcRJvdi/0/pRP1Px3YZ8nELJ
UZ7b/hwGridrU6TC6yNYU8CNQMogydRb9e5ksBy2+C+QAiRTJErAj1lBd4GebVlmuLQxWNTmOgje
cvEdpzjWqS5q4b7M/11FOekUC816fQqunCSZsd6+niQtIunuzhx+VVc25tqJ2VZ4HZ0Ayeb0UMdi
XKhYeirHnKa8aENBLdjzWaZHcH7l3doh5EKTT/IbXujCuVlNFFT0jSoi3mJR8T1qVF40+MYHhivs
Z/MmUvFQBnIuEHRzQFYn0mTqb6ZY4nHXOjvJtYqLV2VO+zuVaFF2haCXVRyn+f73kc0NuybKqQZJ
tgUFVi2P3TYA0jBTfYm7uMtQmqfpwgnn7gS2vTPsSS1nnt4CBXmSed6G1etqhtL2dEfK6XLXNpuS
KfuS6YWXZKVB+aFZJADKe6gTcRE+QtxMLMQJWlQV4BMhf6y8KhWZXYB/lswkk++oal/FCwe46r3z
Do3CPq0G5nLH6f2gmH0p9rwTRJ2nSYJWBIM6YX6whd/k1jnuQ77q+HHPLThOXOjo+qlyfGb1iwl/
XBsL1g0WVIrSiBXzPF0/ESXZ5ejEpXjRaICLoJhjJf6JY3NYT5NcQfpoWMBVm914geoRsSV762OO
AX7cOraWhM/YP890Pg4BLRN+fkJI6ogH9Qco/wUdd58x14JI4IZJbwMPW6v4VxuSQija8SQ4DhcX
s2QpNLli/Z5C1BEFihoU9q2z5kl8QttVXxRwCGq0CZnT4oppYJT54xgc+V14m2jOO0yGPMKsublX
HIEeA1sMX62f/LRxgAmdKVy6NIdcOrsoxpqTj9t46RWrnM5SKEozrl7FexPzlvfpo/yWscKbarq1
LdFLSwul7oaMMJQTbvu6Um7+mF9hGMrl6DcX19d9apDOxsVg4qeSoOZVOytELqBSqqwrIsb74rjP
FvAA1Vhl03ElowMc6svdrPHB2y7sIWgobw63+i6HksUBOKZC5dWXTgyodd22NmxVUd/MeUoG1eVD
Jhs0nLbUj4Ws0jL2IHLGMWCIB6gti2x/LsYZcpgFSMx4bhE8Krg6mFVQfWYoS/0yYt6pcNaVDOzf
fYewjR3Q0Ni49GVEqLVKKE/u7nGDMwohJzKByV6kt9kqikuoaHcQhNVfV0+yDxaBPRT8D2fHKb9N
pUW0HFas6b8olw+gHcxEwlhEIKwZs2JxqJWZBZZm3UdVf6j0IbyhyP0lCxrAtU/e87C2EmaLGWZg
405LPFY/22ZYUUENE0jBss7N8/DNxR7jnqzsOXdRbU9seSdS+oV+HVdBiEXTE504BZPzCwpQh70e
Cz21o5/twTojgjz2uiMrHtrldW9Rnp7GZuItNCKqb1uC3QPmQI1NxFsm2IOXs1PvDR9O2E3tnVs+
JSKiQfA6pOqyT136EuXIva4eokjg/YRr+tgOLK/5qAuzKMsnSd670HCVnGF+lD8YSAFU8+O9shNa
yhlLcYSWmWAWeZ8N4pCtB/Ptn/JdnEM9QUHBuJ8U7pGOOxtlqdRzgR93pDNu3EGQcqWSB8TdL+FG
cqZRd/5IcJ7tTT4MQvxYhMK58gjzt+yWix1hxf3bFyxVrZ3o5uQVFXoXflppyWdEUgmEekjASs8m
Sf1a3n4mY410rP6EJf84djRPO9Y6scmS7RMmfXPAWkZ5Y6SjQ73FOzS5fRR1wBdz6AuiIZiMAgT/
RgupZmoEIyZ9ijcnhgI5SQIuX/LSqh/spXZZSmgAsbpIX/ZgCi65fDZSFF3YpdXkWzHvUCl5xP+M
eEPba+v4HPmCrvgFOyYCs3+NVtF2cgxFYnl1yGZJ21pYB6KIIzoz7rGGN/Y91ToiypK0D6zTKnrv
RAZSihWH01ZAwNxhEgxRXNMIcQbBasqcbrYjo7B+to6SOKH60CrJA7jWk5VfqKFzsAX7eFO6dQY5
eQdDQBGpxSTCPUujsw+idt5+gBpqjB/UhgWWA1y16YFZKIq50uXlwWkPIMWxB6bgx1B9ogDifjOt
YFSRn57L08JRj2uvw8U/GulPGAx+k9QcgFmZHjAAK3MjBsTAivKIXFGXAASodx7CWxB7Scld/ZiB
ki0VykCxPJOhZod1zzdwzGtRura/7xWg0jQWqhNnuJJVcyyPrGbZCVq81ivwlf3uzip5PEOFfemZ
bGOtpA9mdvzwQGXr/NE1unS1vkl536+L8fApfsocsy4ATVmlSeulWI1c5ZVO7ovIO8ntrVZ+Kb/P
K9WKQdpgvLVuvB3a3P0AUlcvhh/+EM02k0GtsKl3uCA+a2QGDT3uThASzUxWi/09ZhE6fyL6521G
v4MIZyfg3iMSI8By2RHay93MwfKlJIiXWE7sC4dPBkmO9+XMwH53HJERAVtgH05OFz/u2cJnSH08
5JWJR/eTjrp2PBbK+SZtgfdVWGOqC3BERsqio5NzW7pWGXs0gyS6LsYPBwA+oKrYzi8LgNQxUfEx
akYbX4ZG9AnwagX6PUQelUwejfQzHXBtYlB/UEQqx0Z62nsPc2NqdO5C2xr8YlWyACB5xDIS/lhk
CbN6jsXJQp2CWB9E3mFhUndmGFAU6onuA2RlY8kIZVXx9acrwUv8krtuXzjeno7i+PFb+ounRvRD
NAGYc0l+kxFlxoxDPewlu/VJD69fPsmnvZqE2AqEKMIXqm85BHy2HF/q8dXRPwiizsMzChxI5EPk
AEG3Yhp/R+oMZiPsQ0faE3a53p4zktpjHI7x7GwRzmVHK8CpbSxUIGmGGH1XsxuIClk9+VCJvI0S
X/RaipPzarHQD3eBAYintoZzstThqsGGoIaUz57xzSGCI/QMTYWf/crZapIpdYqEXvBbE3COfjZD
weBE0DdnL9dosh8r/xlHPgIFnBR0rD+iidzT3DwYXum/jY+8GbB6nyE+svps/svWSjAlpnxq3MkV
G7UiENwzLeSR/ASq0phzQpJKuGi+VRwz4/h6YZFP+jagXzWvXUqwHr8cQPN+aHOjaE/us5bqLBGJ
2UHP5auJ5Hl1adpJWGg2RddbOy6UgQ6NwBbhhbcwdPGn8WV46XHTihdOQDOkKlikyJ3tN4RPmpAR
hsMm6ugd7P+WPOLWxdqc2Qa2yg8O4jPxznWeU7duF1PyyPQ9A1whg/1snDJVDT1eyW4ANxkLM30H
AHtULH45URtvo0LsFuBPvAzbDH8qI5T1a3Yt8eooxDzylrVa7o9c9Bxe95LwUdm6q2sq07FKQb8D
C2FbW97A/Psgo8TEXVN1sjBOP4II7tZ+K6qwWzMYYufYHVi0EXtYI2Aqvj61Wc6NC0b0XE2cZRWh
TbLZSGLrZm4vV7ekbsC2SFEq8/dVv1ulK0TNtbKODPLz62uJgnW4vir6Pz2Sfbra4dqUkY0uusB0
LISMtatnghDnP6mDGS8vBimzLpPEKGEw7G4x4yGly6vdx5kE9NxUdGRVfPdZ3u+zgJF1ZXxiQ3sK
xHoNFbv436ygdRmqvKXzDm8HkYhvwTPn2bSoh4SaaN1+3fZveEIJXJQ/2JORPcOZAfb2D+W5eQ5l
Y5Hl2by1RbYABrxlSyPEtbNiCGf1eEosYnXOsnCNB9tSmnmyhIyWIfNgsCE+Xk72GAzwDD3mbp4Q
pNLjRxPpXEzZ2r/AxUkxFSgmb5owMoJ86Tj+VIFA0eRWJ+LbTxZuYIW7Y1PggycKSuIUlgJ7uMk0
zn02Ua3pYbJGAzJLyiksKvzE/CeXzfEJxebhaTUa6MArtD272es0jqzE7Y2Yo1ScZYva51vmC/4c
WZYbVutVG2V+uGIePWjvTRfl0D/5ExmHr3LdNlJkAP4fdAXf7NSYzE69cG+QxJbd9UNRMuFeZ/rK
1cV6cBd3877gJ1f8fTfupnj/dU6kghA77J+h5JBOJg9sPj3miXz+JtSre55F7jf2Vi7Si1uaZANa
y0aEYSAFKqxpxSxA/cxvfJfglzRE6i8GaBubJSkY2LuyrIEWHtiEodSusmKCeBf9K3SnYNgA/1zt
KRcrpaF3A92t4hoJxfhCmkD/QSt4K/rbZQftO+s2pSzUcFUT0Oao+z6ypvuWWADWqdxe93Wbn8Gg
8gKhK8BYXsF1qcn8/EOtMT8atS0My7sPA7PJv1p9/eU4mmMS1XPIKmsVHoLB1S0fWTYDV8PI6BA5
/Y/0dNtkt1akierK9YpS7kmX3SmhzYhswOLN2aKWIf+zqHh8tG4Fxfl3Y5zsMFaFhMqVSDEhhwyy
rSmP4tO/x4UxW4HwRNZLBdeETFcPXlz58YKipfioe21pZP2COG3mrC3KsmxfVgYsEp/uyp2PPeFE
uqCns440Ge1xsmYW+2TA4/EXusg9GTLy26tGtPOUEEjwqfmJsECJ8msjOga/hUfKMJsDOcZv+LDD
PCEPwV/fEisrBZaxl73MAEActAKWguQLwHM61MMTlZUo1k9+glGCk5OMtpfBSA8xaydJPve/CFjz
saGUgOGUrVnfXAyyUXnHNoz9DxEmD3MSPv677vnEtnWaDT6fWxibCIL2kQs3/44olVD8A6x6wcou
PiI91rs4xi6/7MLhaNJJiUYGuHRIxaXJJ4Wf5pz55F8E+CgZNwd4WXOeIAY9XXYEfiMYNm1AvcGg
BHjYDdpTniwRi8mvnN4DzUuduQT6fei4MZzz2drzGZEdJcB3LH8t3mf1dZjT0Mrk+pB+eBeSbEeM
VDsqQo5KotE+oqrjPDIzzxuGTE8OmRQhDfNkBCaJO+kueSJ9UukrjTHpRIEDQ2HprVNT4CXQhNfE
TeEgwz6LbTfGWFyKAwNjsvKXUFjQE8wQipAnm0qDov8bpL7E9YT8bMMt/P5GYxhqnkCLz46d4oKU
Quh4zHoiVDTkzfdepLtwhqTID7N1TsMY12TnTXNqZufz0b0BSfd9x8Qq+6YOdpxmkDZK+im4qs7E
BuDjHuACTllGoKM1Y/QBbtY9PZ2jfkBjsu5+4nda/XRrWJVnKPOmIv8M80NWZ1lOHckN3ILcezcE
BWHx8Yf7sHrHHYp0BatCMY+qD4LMw5s5FI9pxL2e63oGHgk7X3F8IAZcukKM1RbsRsfLSqOBNLS/
CVkARV4vie/8UUO/VSeGNw5l4SCI1kWz0YjtYlJMChwVMe3AiVioe7SkYFOqKAaQBwe6u1AnY49a
PT9BEDdZPcULC+36qYcl0KSMYWW3VOx1no02nAln9qlOdFHZiS24GnTR2q7ASSIczyhpzJiXvG0V
4U56tjTBbWfknn0hmairnFQpBkgwlcAelef1b6x0vcF2l+LX+QXaCEZbeD2JjXCVhpcDO1eDZUpt
IGFXaD82weVcv9pRzB//EyIRBhxaSII0iiR9EJMLN9YndXQ3JhRGb7exACEer9QwpKl4YLvtRhhA
ENilCAgQEHQ/FQIPE55O8Mm532ZyCGjHCqtpG07nMy4ApLAJgY2OlSBWU94OE92cAmb2qJXEJaqh
Fs9MgCK4n9JUNOkM3Jz6TFBov/s1c+ZpOjNCC/iT8/MQ4d9UZXLF4/mhJL2YIdkXzW/zMd2dJltX
L4xdXqyKI+wEIBwelBlH07F5UdWkEiiVqyNlUsmZ+hl1rS4iFC+1mkSv4CN9+xhyFxl64haf+T7B
DEvu/Dy3nP75zDjBwAqDEWI2y2IZFcFUjkkRrjSsVsN7wHbx3ZI3C8CBF/GyO2L8NWF9qUUagnM3
nWdGzytN39gi28DXL+8ptoAsLbzKdAPEKV8l7Pjb0SuIj82acQT+kdf34KofuXYNadQbnvySrrva
N74PsP/v8y2z+X2kPZ62gnpVpno3mV07AzVeUE33XPiLbYWq2/c/FofAagZXfTJEiDBuEVxbufAh
PDrhHv7fmJicXlYWCTNtBucKNV1GVQOUbr8fjpaCZJ647iw+LtjZjWsaFysSPYk6aKNQ8sGl71P4
UxoLO2wa3q0RuPY1tQCjoxa7pTDBZBCcn8pvQ6U509tZItUAhivS28p6Zq+r+inqqbcaAYOJkfyZ
PtbyU1maEcg51KEFjoBCEv4IjEUkfzS2T7OMyICwDOkQSNYXV9DqHtlQ0RZuSku+z0u7oMoU5TB0
aJiSRf0kiwOqmYo4sCRAZgpJRBzRxdc2ydmKh3XFNuWtdWjXWWJofQ1KFzM3dIqbBfrBdjIulXH5
sy3oWac5Omo7u2b7+urvPxa9TqqQS/bH+RwE4/xxrInV80SJoddI81nUMzTtcz6guyS2fBFQ8eww
1Mduanb452qUtNba2PbGL/CWVojuFDA5sHGVa8rpTfxOZpPHt4WoMXSrqOUeCeBKSSOVV7VWU1k6
o1rhZ/YFRQyd0VSKhBS/1uORrm2X+x3NWXfcWrA3rGL/+IgySFvd9DybVYJmCe6yt/0JmUOp5amm
M6lY3oymL0FdA26v8+FgE5HnTcNiVFGvFV+Nbf2rmIoWwSuVHoszKjinr+I2Dv7nDl/5f2LIgWiC
VYXm2JMbOd+z/SdHwFd8rsJbKRX6Wx+H88efV+OVXXJurS+IT1LEc+gqzmmlqAhk5dPYC4PradtM
wZGBac4qqBoxqSI6g2AANTzW7a70pzx28KP+WIK47awg1a8YEFw2UYK1ElE16o6vcge8/sYnVkBw
1IJlUoM/+ZjKKxYE8SUWEHUqSQLnd9mnhjcTNWyUSBYukV1ZDBkdaZzxH6RURArzprT2wsz++xmw
qWR89GkeJlo4vermm6vhZVfI5eDryrC9wpJY6qLobrxaDWkr9tJ9+tpF/32YceKGrOyVkaVr+YL1
vUl/Mm9DH/AcdEh48LtdrmBS0TVVcgb8/Yeo69wjH4ndZNHMlHZaZPqXN7VqbOPo06S3Z+n6SVE7
rpeZPAW6BSxX7NSioYNF+xcnUBTbs/DeZE7dSPI9tmIKzBFGomuJAAx2ptTPwoViGEa/Q5ONdXQm
Zgte0kdMcTfiXN/ViuvWRGXvyQUQkzBFIdx8LARe/pGVShFixiNs0WmAMPM93eh5AstuguzL8QFW
qU0sl/7lNm7Oo0fHt7f1gvQFl4sPqKvXFqE0UVUoFA1fcKrY3rVeQaF5zHoqDCLuQupnlPPaeT14
6aEJ+KkJFj+Vwd0ioU+kGeMF+egLsi5+WnmqxwcPYcTUIuCyzybM5+nrZIWc2YIngebhOduuD9iR
+nmtyIjRcQqkBUVDaaSMHJiTQwtujmUrGex7YXlBkygKx/Ul75uvfImzO/QEl5Sz7Td5xDWroWgC
eou1szCk+5NYsH1YIHslAVPF0L/cOzXo1IqnvuYcEoeZa8wjKCVlh5Ocg5Xf3aKK7A4QmX8i4DcT
qJINczY+/QIqfHcafTW4AbbAdQIB+TXjCH0FeF3ddRZyb03tkegQWsK+Dgu4ufHxOlNYyPLkB/Ie
vcJX+3IgT2NeL0djQ50I6VmoDu4A8Iu/4B/MwYekmQ1Xw1okhciXqlJYceDqMHRTdrpzYABhQLs6
kQqrVoRw7/FNTf3iIPWNUaBzet6IhFEY0DbG81/OKrnVSr3fVuO/+kiNQdAspFO8M0gEgW013KpI
KKEdPu99J/vtS97pidMwE8giJUPRG7A1aofxZM+yO2RMObVQZL0aJCeiBpqiFDI0uRUXW1e0QCGn
PgoFe4pMvlOq4MuAwsGhFlANpQ7g3rUFZEn0NK/iUsuRmz7zXzzEbmCblkdARS86eYbSCXGdlnmn
/WY+BGntjaHytKd8GnPScNUR6Qou1X8a8JGuaco1oGzaEnASd03AWEElJ2XEmdXB52HF9qdGcAuh
+oojkSrVL42aXge/lkD2OWz+D+S0LhW/8LBavcQVSzJ98+hz/bWA/T24Y0Zs8phHiBfNqL03kfww
xGXeCo/tlqmxYqQTB3bwojQBIAPAtgjBlcEZ12U2Sq0ttvfPcd6eO3l9L8IuK6oAjRURW7z3wq+m
NAdhLpU7dAswjqJhdr59ik1wj8vpYHbO7QoAEpyt65EAZdDDwblbFGES7JHByKKQ2OCNVlLFyjtc
WYCkR3GIH0x+hYFKuetoMY1FcK9BAGGU6cnxS4OAAod0IwFPnpWb5Hsoblhbn7KFCjY/WqQhjMoi
EhvnJbHGti+0CGdp2PG/6joU/XDgB16nqZnc0iPz0CraEw19dvTNNDl7B9jV3q1tIBQLHb2mYsen
3Bdr+chXreMpvv787R6apbCA2VUNXfpA71ILO+RKAdFzXHvB1V3EdW1LsQEaQqqcknps2lK3pxvu
vBaRLgNgyZkZ87jc94eBJysbq8brx0uB7TngmJ9uNhSvVSnkSnm83jmI+Gp0TofqUqnh7JjwoVnO
6xnsHmZxZHJeOBd617ymvYBh9uKfSjCeUdHbb1liFW7IBVxoknYHzFCPnGlHAtBKG8DSQhSIl1DW
MK3MrpO0hktGvWHH2zTSD6Dsx3hl3d1oqEnOGOvBF3xBWGvIqKk4gPaNlVu3p+GxYsa2MVQ2WXxW
jL6/VDldaoVSCSgmFc1GogNXcQCsQRMz+4z93DDkK2AzOGJseU7U/TH8IPPpSlWlyMXE33g99tRp
4zlxACOWg48Ki4REe6GfAXDO97wAf7zfxuOBcRYpkN9wVKWKkBTaHYUPDTixFAE0J5VuV2zKrXSC
rO4l3mxEz1M/RqD0T4G1ejlBgz0WB/Xgl7wB+iSt3J46oT7/StHwZN7tTpTHEteKypSfNoYaqo4s
gP7yVB6KmITXGfE8o9MkPPFWdA91xgSU592PwYeP1PYTab59s4+UzqpCwVwqZzXEHHsjcKw15c9Q
uFOWU45outhsBTihYfn8SLNTrPm+RI7eEbiUQOXlEMNsgO+YlARt61tK+FWOdVhvD9tvV4FFCdGG
A8wA9OtV0OqysuRBdWydu+iCodOTdOapao0f2dCw3bodrC2ZmoFiBEHbZFo41VpI6/SYeyz6yJbr
SgWjgW9GWG2zTP6/rpCee91YZzghIicQlEQUrhues4J5E8zgTcB4ygaJWNiXfPJ2IBc44AUWhMVi
8d8IkO9akhdjmMSL2nEFwSkR+Eo0BgI7VsdkQ4yWWcMJs8fQWbS2MnBxt6ke1TcXfd++usz0N+G1
IGV8BrEvrQLfaZp/8yKqrHo1YljkfQt5ybKHlWAkOGcvSSjmoL88Od3435kcyIeoabN386UnVhpW
d0HBzWHByV4GSfm3MxB4RxKDKe+2PMxF4sbTMduHhtn0qJEFGmMO31bEUguqqesPNK8zpUsP82GS
Olpob/nO19WCmcv+ZBenPrTO4zl75FUp4FthzrUMz6tYqt29D4TxkMyFYU57K3QXanbhS48JCsVW
hrBGg5P/XNaX7pLmm9pNSm9jYmhNCgg1uq95gY2UU2jzyyY0tSyQqSOr4zxXb41ES+RWuEqF80qc
haw3X3PWrb6xfngTKBQKwu+EKSi+i++kzxamrFukVXG3Y5IAN5cXEJ4+txStxGNEI9dIWsXBUTqb
5E0sWsIRxb877yo2DGcZhGuoCDFrhqEdL2GXnEH+JfvYyidkIgFRmMJrBhq3DeCHP32h30CyD0W1
WF6bln0RYptuzobka3heherFpLhrV+QJfLtYA86V+ZhFA+WiwlIh7LNKE1IO3yyDBdn87lktr/vT
lmLaEBKjHvStTFFM4fsMJoCxh4iqJ2pasAIQXro/iuEi5dEF+Z2gXryvgjxiCj13UFS5a7mp90Am
7h/VhI0q2MWFXuSSkV3mMUQ8YPnHi5N12nXlcBcUcRyT234ITHHWF9aYgP4aKCJRyhtOH1CFp1SH
M/XnAzUVL9mxPyfyoI/6btDP9GxkyTxhY/l2LkfgEEc5twU+R3f3Ylvf+pjyC7Ly48RT1QU/7cl4
TggRs1HksYYgSb3nzO1geETq3RxBZ7F4IDrUZFgJy5BRBLquHfy68buNr4At03kP6F94Foa+roZb
RLd9t10kQ7PXlolkZXhK79a6IHvyGL6s5CELAiGRNDOsO+bRVDp04KqWI3ir8axgr0x+dAqN9Fq/
2RaKW/ryOo1qWP471cHqY2Ws4C5Bn3Md44ckT7Ojp+D9Pn0WME4izjtOJopDjkRi1GuyjuNelOId
cyHxEdJkhSQOhoFKqYaJUqhjo3n99wM8mNMCmGEUyGb8dEvjPitOrRxdxfJnQFHp7BOKii5hObz1
GsdnIXx+KBLrUNxPRGF6GvC7xGASWF0jPknu9cNt0r2XpWvX1nSziAEpyadarsactoYXEPAMRtTT
73uRWczvccjcNxcSjEzjhGlgf0/FtJg5mGGBcIQmf0UPxYNBIMFV+BF15QbJ20otymE5rowi7uyn
+uFG+3j7Mk9UrwcisMofk570F/rYh1AHbWip+NR2eUk7dhT9qko/CgKFknbunYjr9fChxqxApbDn
llIcpXUS+1JuUOceSsQfMQoPnPSU+8X0GSYe1grI2RbQxoP+qtG+XOpXqgQGZ0l1n9KWzIAO2HxL
FRB8bCauvakabV71tkNp12tXk3eKIeQZklvMkLexzQ2OZ058fr4LkIRnGQwf2K3qraxSN9eLFgOg
x2xIy2EkwR+9/GuBX/s2avm0zkGxyaYVSSFqo5ohlhUZnXCFANZ+CGgFBl+PrjvVa+xDzslfoZKq
UM4x8zCQhEH/SBKkpPQY4+RlpSdU2+z/6xtFqmAW+EMYVemUCFxIbdO2r2MIqzZNIJ/J7obA+4+I
FH27RqTxvLeYLKpmpE77cH2R0Dvop+zAAaEkIjD1dqi433FNPdV80LjneGp4vSO/2gcdPu4nNo1z
BXkinmbg6Cl8mOPS7dCS3N1yeIyUxylFeP9Jg8WT2G96E+2c6a3avum+wXLxx11qIxkQu2+DZd6H
cwHLxCXEagaQVZKz/t8ewsSBN5LBaTCQEx5GzAL1IpQOypfQ+79F+L44o7C+ji/uT0ap7ipIWDtC
4nhto4SrHTxWQ3LTP1oGI9WTVKlrhOOs4vuyPOAahYYEDGvsKQJ+ixVOb/VG9/PUD1koi/tBuCVX
nofOguc3tGX4WmQu6mITxMY3zDN0VhRWqWIvIbohIN4gPEsdb1C5Mi9Y2zE0L/CiG9U2xydIetoB
kc1BJnSmn6Gos6wMiKx6LYqyCoUnEiC0Phds6bX4SN3WbTXLqaRfMR94uDynYqqGiOs6Tub3Py8F
U/FS7PKVR5rOxkCc/j8plDbpSZ8OU0dyVC2B8C/p2LovqlY8qQZNRVms0tiWMkS56+nW3/K7z5lK
T4WncCcSYRayEtA9Py+q7ZLWHtZ3jiCKgKhpi0dIKPC43UvO0WT6xyT1DLrFqxwuk9iS9pDyrerF
8lNEivHoHau+hApEUVxIA1eSAEzI7bmLBjX5BJ19J5wIOy27WFahz5DzcGp7Os2laMwGBLreJKt8
tFs9Nw7NaJTNsEsQOYx/hodcDrYm1hunoEoWEDvoxzVqFYYnqFwj+wvRICTa1CNkB9vplfgsodXe
4mVP9D7uMlvCJk6M7eAjEf9DnG9hsfNDtTPx6UWCzcnFok+n9hsXv7/wcStGAE/fjhk59oU81Zgn
GXOwGu8Miy1giU9mA6F+XkE814UYupgMb+yjUIajl+TQ++waYH769oXzzwWM/3G3zYf7iSVXIPdB
aOsufO5lf3qmV9MYc/+Kh6jBGLOLOyYxCs36y3Io1WLElhQm1pAO+ImVDGcbd7hSME6TOilGT0C+
zdNEi0albdbZkDNQ0zXQfIMIPSt53iy7jyeRntCbzsgJVJoATtkiZDr9+oScPIz2lS3Mzv9lMe+m
GfCt+iOVUjGyqoUQTW1J9UyBEKWTIO2t8+uCpwGmCVc0dp6JIbKbDPogmw6nN50T7G7P9sDmewQj
SriKGWdoVCM7jdnp869cy1cPF6gbQxET7xoU8ZCNBjNgq2AzSc45ty1Jdy4PEVe9KDAbsMri+AHJ
O+W7vu2Gdozyr9fLNhizw4iXhyQOC5AYjVD1lJhLR1inTAZPVhfqXKsgD+w+Se2p6B6PUrIKzkUp
8+jB3Vcz3e3PogHScpZatxqnzbEXWCKtwajD4sZQOzu540kIlVQJ88jq9ALTRAwXj6jo3/LQehIO
aYOM2Zz4IofqEt/aRlen3gkBgfo06ZACen0AbT+npEpivuxSIr/dsQLnCLK378lceGqD28A08BR6
MKH9CjJpssoNcJ8Acvw40gAaBSmrv/im9Msjh1nPbOOUhPNjFhVIwTM3pr7+BSkAppuaiFeuv/e6
qD6wtz9RShg+hnwTiMpaQqo6EIr1ebQBY+HlMHNRv05zGJL9H5HOUdNOIFfTBnxhoWnoi/yQYl8V
V8J/siw/S7bOvzoc0t7T454kOIR5rM1uhdJAUC86LA0gk5IiFmuh2ghhJ9c05MqZTdY1NwntWhCX
Ohv9gq+NeXp5gQ4mr0wz4ilOVvgX1u32JyosPdcMj15ftaqSK+pR8zDt9BanQgmtTrcvheM+Gt8K
tSmCEeQvWsrhTqt+40LnLNOb3sGtoofYX8a1O2vnUgaVXN65v10x92jvyxp1fLFYL9PMBQEfU9SX
ySFB5ZiiuaK14otb++3Ye5im2SQ+iip/uvNNMBJyFA1/I7xOzDqyargxFRoVwLCkXO5QYObjHd0L
vLZqCgbGD6H8GX6FX2VRvhzJU4qXmVI7A6InbKrbXPqPxj5w0rP0NiKw02w2gOCQijjbUAjGjQ5w
4toq0skmvfKDO+9ISjKTwPO4pcMyIjk8vLYqmH2FPctCdq4BBeIVLJGTDgLRFPq+70IQ8pRjYMgP
6GmDoSFJlIHqTfLGYGYrQDDzriGmS/11NLMcjpI5zxrXSUJi3RsDp+03OG425BqeD7eKaj/BF1y3
0AB4/GazauwlOfiUnPjfqOPDTG132tFW48r3g1KPiqC605a3MqqikVm90bwHjBiOYYwg9WpLe+AO
kulv5OZyK2qzlmSqGA9sF4/ISNYySoPV8vqnwRzbVfUw5L/09S+4gVPvmGa2uG6IFWvfwkASBgHF
Coo6HB6yrA+Ww5SJJppFPXLRDjbcKxmvo4ICM/HS78N2+YS6W3gHTj9QxcFoMzhBZxiCMM7q7WGt
kHqIHFM6a0WrfsGd7/0mjN35hyLoGX/AQrCFZkEcOVyD/0YW56hlsGbBUsD/a3nm6yx3YDeW3LAx
mHitXtbi9JiRzsp0RZjSZAHJJlpueCJmTObIXtAplbbJ7eFb4DtC5ZmWykeLPmXjqW9EGdPvVSPK
tXfEEQ5EdIlOxQMz6mpOuEEMEaZTTzzQUmdvOoY6JrMJ14Gls76BN+P4qyeRjiZ1fIfC88m5td2F
cjhBmrXV2jEK1erMiMz4LotvfaOiMnE40wdfvWeKFGsLjRVjQmrx75mTJsRv6CPARQOzpXZZLiTl
DyXcEOj+9NSbL3suA9fcFeRsZVckMJ3YgtbnHTEnvz/Nn9aEyidq8My/FeXn38+hGhrfiWxRbr80
zoCrYfTHYet97Yzp64HwPmclEaA+xhl1KHJbmyxIJqS85tCLf0pvfM2sxFiaLnVvzp1u30KU2xwh
n8Y6OOq4RDkCRxGSy//AkroN+mFdyn3W4x/CoTt3t/xxLFI1WbkzN+8HB146jqXh1r0fo+p/BIKH
KV5/VKgu5F/JRuUnQ3whwk+kpgbgwzv4jedpSIoaLEX1WnTxSXXYazOWM134fmqK3Xwq59evyu0h
vJJQPoWM/SkmC4LSgNQdjzrwRHa09pYkM6Oq9TROtkN1TOSgc5fPX6ozwERPDwys3Df3aMnWYqgn
HCQr73ZsBjGQhXHYxKfiTlEXgi8hUr0xawiCnVqESTIlc3N7y9rcKjrJ/bk+nNqiOmjwMCWUlYzD
LxstBmxxOXx57FUBS8RQEiO2taaPvV84XesLGZ9UfehlTzmZJXoyvY6TzfE5gmZHzuWPqRm90DpB
qS6N9QGWplaQzvFThg9KyQMnySdQkI+n3MpWSGISFfkliPg/aOcW7tZ2tDoNqsT+ALXgbfr9GO2g
pfTVQlhYGn/G3samzf9V57cHgPVP70NWhgsonzABoX9a8Na8npcdxaiPvyN4ns6bK7lg+gI9FBqp
phkznYG5uurR67GSSdRht51ABR9BTAi7j/bOMcUIp3ajKuoF5KBJz9BYdZF8JRrtTkZT5M2GS0cb
O5N2vLD4GGErLaFtSnlE95YWIRS09Q8H+UUmRRkcqutKC3GaWePC3LV4Rj4+ZK1pNgJyAm4ieShM
Jovh1tnJ0pbkU6F5cNZg/6VSy4Lv52S6OJ+nthnSUt/vgoXvAW1UpmPdu3Zv7bbfbbstTjgQusvy
1gocYw/0ui1OIP1DhLEFIdgveZ15CROHHcpRlr1O0kPseXT6bYUpN0Ctt+t5C9xcoz3v2aiHwH3y
9XW5yXIe/70tRClo8OaIKlKMHYAuxUnhr50LeF7UE8K3fL7a8IAg5yisMIAcEdgnPywwAGOsKF91
o3/chW9y7ciU+TXhtsltmoM/tybwvzxRhmubPmhhNnE4avZBCm7MVZUuaLRl71Tgj6m+GPwbm1aV
TuPjVhxIZ08XGrdYfWntmuitPaWkaF/Cpenq/3J1mYgP8hPFwOn+eSY9oWKmq5pLs3v362TLdKLg
dj+Bc0XDzl3LAxUuyoTg3QKqbgRRq6apYgjARKchWcOF0L3g05nY3WzeKhk+8I+Huks6NIQV5LWn
CDkK/nC9ZZRaVJsCyFA5dkZvLUrgtaHUvSz9ZvcFhB+z5phHK+uI8fqlBPlf4JzjXsfpEf/wwpAs
LZcPqDdXMrrfnfQOqnEPDXqM8P8uLqJFYE9Be1Hog9RrY2N2An8Pd39iHUDhs7xa7ihoNMyRuTuZ
tjJrAJzot7YJ54OwIoKLrBwy7OfDtXk/vBRHRxsI4Ba6HAOfQY2zHemwD2WH35aYwaC0wSp6msJT
7XjBinaQh6E6aQhmmxaWp5fDa1O1+x0JzrwbYhYkLLOIfkAygcqIShXseJhkUJjOycxE7LCxWrD2
ivdoiPH+YP6PkCHFYFRLt7MNAqQWvFPZRUvhGUmD4dFo3xS4Ftrao5MjggSiJ9EB7rq90/YzDq6s
8YuJFe4znQ+n3vYCos4wXVRVXBmNO8W3unp2mTccqDWcrRyukzQaq6DcjxFXRcK+sFOYDta/hPar
N/thLB0kC1FXzGHsI9nZBg2fH/tt5XLdKKtQv208c3aeb+GgbziaDSxFLTZUcNjMuRy8PnANzccb
nU/E2ql0+JzlaUFvWcNqByCRDzkGWRWm38+fkTPnC1HAG6gOz/KzZz02gZPf6bUO9XZcXVpQdCWd
XqSvZ1KIgOGrk3gxKO451tj052/Ouf3Wli6snefJgrKKQtQyKallXSaMncCa5bEk9Uc4nSmsicGf
C3CpWx0bfGj7qGOmvJRFYDFSny29SSgBokcnpFVwnr8eL/z9p87RIoUJBR3Ny9/7f4Dj4AGKDFrj
erzL+tzRLCE/8dOSG+848ZQn+S55fPXvQcCZ4QAURmVuCLrK4CG/Daa241haKnuZIW7Fo/Xisxrr
2z8AbBSevsY2az1VRES9uHgPNctmCcSmPo2tWBS2l95hojyvA65qa+vObtVlxrr6Xa3/0LcjZyrQ
3lIX6x0xyroNUo1j8uFgWUmsFwGv6bJ8ox+vBdZk8x4U4LvNTWznKclhvx+bO4kTgVs3MUNpWHuP
byBCq/2LoRZ/zh8WahfA2EsgsEMWXR0yO/VNxIeSLnuADLX2ohCxUPiMmNjw0ylvLSosP/p1hPBU
+DC8Wem1zOyGbePOX0SQbabXDUOUz8Cbc+UgSxqcikihIIxHdTvAdx/JtEAFKPgUBu5PA0J9HMIm
nayfKhAcFBMN17JgL2SMinSWd2sBavpgk8iRHsNDEvcRd3V+tJ189aMZKJCjltfkkxlWcXLu8wcP
3uZsDHX4CIe6C5pAokWMC/cYuJGgruEmuLtv+nlplExMR9WlbHgLp9ddl2UcE8Rv7rzJXhYAFSfU
wsz39lgypWv58tvVF4m05vZKozFVWrH+A5q8Rr71vyGJkqAAOIKBS14ZwlX9jZfPzm3LY4oWZ5oP
y53TXcP+T+7f8l11N5mSwaCBDkdrZkcY9Jg6UUsqDbhGpJgkHdeBHjOCBE88TaBnQC1wHfvQdlXx
qwVfUK+AUhXjd5EdkV0eLRi67NEIOvJ3lYFfdp628ULapSlC0eWGtvXkGdM5HW/G6NuDhApMjJWA
gR5zq9eicFWL6EJX+skrsaKLBa/5JzdBZVEn+11KdnLJGCDTNeFI501bgqhJZfF6uHGUmK/bE59s
dV2hhmvtHV4RgS22u15qPgebdgFMj7p9x+oLaOnyCwT8toeD1faxzU2Rmo5/XtwecbUQvmZHcO7H
NPO/65zOwH7Sm9cMOxam3u33fAuHjO+5Deo7xR4PKEcCJMy0S7PJHKi2o66xT2ny2oeUFNDVtOk1
REy5sfPZFpeeO5Njev+IM4ATsrWOG9gkAK6xXPbmSPCWHobG+ZsiJPwcAxY4Rjl287GnnzYv+U59
HuOHjZndfb7fthKXYtXkcS4xhJxKZClRylNFaHRzQ2PGcyrcuH4eSjF+4jinoBYnvp3I8kjq1B3e
JgyHifFwb1R137nI9bmXgeypCGZ/VbG7UCb+WXRvMntHDKhlw8rT0stwsS+rDvSVhkHrwQAmC4Z4
V2O0TX34U+Ar6QOkAoco56u16Xwbeo+lSUV5BVCYK4JXw3jg+EjH1t1br/NzGIztHOAkRps4Xbdq
j95Lsydo2VbuZMJDuvGf9J/OR+oPMSPud4wlw10r7a8Sx55ARorYSKw0hl1cnWDPe0wuHxw027VZ
zabfL8R21+8EiPUpuDfvBWPFJE3jLAbrB8SFB3k2arqLFPrhKUI0BIEdbCOE6ZnmLBoDYgY0+GD3
04RLFDLHcIiiTRStPPNCrndePTh5BLJID9vcTNxWJ8khBKxaqPACK+2BgzEd/vw8E1bMaYX8ldi7
j0QrT/JAK1uG/jD1z7R2OVKIuXi7TG4oH0tP0o/e0wH2GlDhtqaqDh3X/wG86UPOcFdoUTUpBCCy
UpliXt3BBZb6lGemLmz2JNyJoDONfmqksYbKNRm5m3wu/e/msEc2IKw9664rpYi8Hxcm0Bcmw6f+
ALD6HTTsHs7svAtxL3wKRins80y8ZgOZ/yV1d450rN6rTOaicIHeMRCeZDRxjZGO+RNJ7BY1vUck
fcNyDUJHbaPtIpOvsHpm7V5kZ4MThemgUedDAWy53W/4EtZmvDiSfhGoG4b8zjqcjS0ukvzRxIRi
1zlhL5a/5cKJE9Tx1sWQj7Bn6nPpLvL67aEVU7L59H/uasXdCYNGjOi5opD8Iw2sw+FlP/rU1IJI
Kim1VQj94TbXe9r7dzYZYQNFS4w4oMdIZuTWxtw32xZ7Tk5rKdcmGJvhBkSLcZsmn4JLAeaZIkf6
VwSYVNC+AMBs14WB0+A6b5c1d+ABONp6O0IxOIWz/N3PdAgjMxV+Bs8JxG1aE/pTnWwvF8PPA6p+
izB2DTJCuHA159aSAlFH+DsReKQOGRzGCzZ/S3AyF4zL/PcYO1Phj/XuZJ9G0PM358wYjQmafBKn
lOplasNz02dBJd3mcAjXjkK9/BpsOK4WxNc7q4rJB9kz8SKkwNmbgaUfrGXMslZZbvRM/TsJrFye
3PK4UVwkxOO3AEYntkcJJlRxygC/I8BiJkM7Fj/Dj3FXgBoS46Z89gBVSU2H24NuOXugdQDHyRyr
DDtGureyMxyrYavh+auU40j9Ob6uxQHpbcOdUllBehbBPs+72Ta7nkeNx5STHriwJeB1ArZ8DQr0
Vts7eqtmsEMMe/fBQXLoDp1s7YizDdaTK+F/FiDQAFUkwlCwHShQ9XnD2xCVhW4LTRd1FUJ4ld/s
ejJJTHC+yyRzYGvomUfJx3Sdn83Q7WBtKqa9wD8bODFnuJbFjhI6VgNDUoHkCKBUM0h79J427Qp1
3iusWSMUT6OQmUDfndtX0tTOtTyhlSH/qrClmFQesO3DQ2TLAAN4pamXFq98VXtHKoHyndRCuedy
1vvF4wIv4kEDLHDNdSgwdwibRFP6Kg1RChYOxEjepLGEXHyWysFcYyK2xM99WBHSIIMZElKuKfIJ
PQCcAGrDQf2hXovlqolilDuLmotck40EF2GYe5BnyDDCmlYtf4UyhjuObVsHFppqgpxz9NuFHqnn
uQNTZYbFsfmDeAuMpNSMznao3Yq24EVg0vUk7wOdRm5zqpphwLY+1i2ZRN2KLWzovFu+PVffTjrX
/L5olXDbRuCSJDgxuBMpRb/C9GQmyUMBP9Wz/jEe8rhmWdpyRXILnJyvESp8pNAAFAv0j2d0EW5j
mWT/xdR80O/H4qOs6yZFbLjIfYoTBqs1g3EdyOH5jFvXUii+JMcp2KQfTKiSvrygJeZacbqCpChL
Hl6HkwOiy/CeE90s6/iqT/tlk3RivCEdKIDNf3zsgVMA/rVHKCj3Vfq4dkkvoTn6520X6ksssg2m
5LyO5rAAYu1dHoAJJzk8tMNNx+vc1mvOr7f78Lb2stkBxSJ8Xr8RWlnuRotGhlODxGD1oWnmCZpf
NGmCQZUDfsVphfDFzvdWaYJZZ+Az8f3EikfYegdiTUa2oD0eeIOp7A/ZZ9URNcqmEVagrt2TtWt4
pbgD3UUXc5m1BUl5ziMCoWjuCVXurR+0lPluBcJeuYU2hi8j9iAsok8A+i0U3v7m10d41GEM6GTz
abo4rycEAHlIMwmNqrLObX8gSWXKiV9f+zLwLpnQ4dl57iw+PiIWdnE8GXNacx4sqe56LU6SrKlm
uRsr/RKjfObBS9FxS8Zt0QNyOW+/TuW3bI2oP53p4cahrj7RBbR7CTpcgY/i6U7L8bQLA/Vb6uMs
938LX1jQzA+OHKkXBVwAyWDL5wcdKKL5t8Fc9oFSA9GgjH4D5X94XbmJPJxT7474PGti0w733FpN
sIs/9ZM579DUg5v0C90w9daKd35K141FByejZYbQwkDhlSgLwb3SakokV3cUiuuht6l9P6KUahzX
g4ixuqSYFrOCIUrMHffsBBZc1BwDfA/bSYyHW1KlTHRTjPSGkQ8Pm/18ksY2wqkWSlop1yHr/Aws
caeo5XIsylbgJb3ByvyEZexCx+odU9dR/XLgBHk3iMD7LaLsD1va6R+oLxLl3GMCUn4Z/b6e5whi
MKOYtH75OmOEHlKSWykK5gZjaiXM2zy7KcENvqsZ3Oj7QGuS/I5sdd2JiCis+hzYeUbEfGzXtGHA
to30bNrGHgomuWGs0Mh48biI1ZX2MRKbGsGTkQESG0iEINeyUFM1hmDH2pB4Po7jczVU8hnuKumJ
yg0ENW7v3o3FaHwioyuAAJ5iUTpA4LL6lR5hEdtWt9BUZBn4anjh3H1QFuDXxckExiQkGr/Pi0cY
jkBdmcrZKpHz9CC8GXREwWIKw5m3KKSmp4PjJS0zlEeCPu1ZDEHAxW6t9z5oyq0LOcd6YM0YsDZb
BFCmcqQQc6p23ET6tSgSD8aqWrt7RHXsCsWindbJdeYh21wVId7zYl3C7lDbCmh5eR4lqzd8Q5tY
SGTD46LsP11W7fe6ggWhUmzUkMHgRvt8C2j+jiFu/1bskK3i1Qxr7WrNDlzI/mZSuSRH1jttEsZN
kr5rhwpW9esF3wPswdpZnB5b1+65hDS2MdusAHLtobKo1YUVDzs9sVTDy0WwnPBEYwG2i967VKgf
1vauuhn0uSe5W1xn/a7y6hrygIZgD/zxtOIdCcSEP0dKh1vHdHnj6U+ls3SXa7cGosZd/CuPHP8I
J4Bc7ovS16NfQqiX0n/oQJcF2kawzHILktIr/gSWLh2hyrObaF0/GGsL/xnQCzxBlKtJUu7VC/zv
M5Ga+uYPmQmlCF5SLkgneV1cpHwVdE1MNvjWOMJ8WUV1hyp+XXzoAphF6J9i9vGcwPWlH9bQaHV4
TukzkuqWZrg4CA/+fUzMOkvGzFAVs+DYZElzRxItgRNPzFhBSwu5f5voNlB0vSBEwilj1rwMsruV
GW05ojja3P2Wq7FqW8xtKVopZ1b+BaxzvNrNxIrZzlSvKLXVZWXE+gQ21p5Q1iUkTSyHDhtYTSvj
oHm5/RCvFsCIm254ZVw7RTqBskxrqTWgkE82KGN2cPXgbopn/wPISf4RBkkVFRXJmnXDo7umgNZ0
ea5HskSRpXfwtHHYUm9Upji98rvllKxRw9vX1hwIHSuEyWkywvvoerBuXzYhc4nDCZZF3xxn6c3I
lRAL57jIenyocbzzHv0Y2LuKOcPKyFs4vR2YnwoyIXE4dOTR0GlwtVCC0bbraS2LgKPy+WcNWOp1
U3hiebtKrLoECgfWb9WnOUni3tilqZHl9Mipg7+WnuYu9FZoxo0cxke0WbsR9mXcdtg7v8D+4f5g
m1aAuZe6R3BEldUsjZmp5+5jdG+MWyE/dPeXvRHGEwJatiSkpd4fDIEUzozjPoqdFDu7XNc7fs4j
SM8LRK+dCaFnqM3iiGL7EpSSg8OGWEC92KbNse+02u7IaZauPJsdrX1gOYfSQ4T36PqV00liEqTt
snO8gye+wH6nk0SxFz3Fcp9AQKUCkyr3+2fl2d3zky8uoNlc0bGYKdaZ0J7MVzQOkB4XSQ1gvqJh
2fCfG50VXjmWIbgYVZER4Hv3SJdZPcYh1hbqF3Xu4IsYpxoYIQ2KXnTzmpVGdMouppeB81UHMgmI
bKWGY++xJnuXIMcYbsXInPfvMCwlXujBVyJ+VClMb8BImBR8R6hCEKz4mx986uLop4Fj8Zr4brV3
qkx5d7A5O/N2ixF6JzaJOn4VMebuCE5JSyQiGgHGue+D+5C2bhW7k8lbn7oZjBwaZoDNMEwzFFIu
JfuaD3ojCaOi/YuvWwQsQ8hiCi13qaih9bBRclgbGXWPcXrOY8GXILTzus+b+VmdJ5ElZqr+2EB7
/0wCKyeeI0DvKKNpkSFgdLHsj61DKpgXhakE+c15mCBLnRbhdglzb7rT0mueriuRtYPy1QqzsMy9
TTSJz9T7903WMhKzgpiqs3STrpqIeFPxaYmo/ct1sJ1+e7sHSchrXVvwuHUHL1VefwdD3o3uO+eL
sojMS5MYQsaJeIhHYQTXyB3CxwKzkx7xbZ6xaCo8m8c8DY1sk9Xs3BvMGVQsyXPK9S5YApjaQfae
mR+6Pc5sd46qZPszRgByrDxBaVQBaGPw3htlstVRwET7P7LEfbO+K/EpmdEZBjIxi9YV6tcVA4CZ
L9K6aK+VQ3ON4rXr6EHW/2pW5YvTcyOXpPJbTmw9W11daMLqsTmmHzrqxt/1e2kFC7RGEr6i7cnt
wh7XJqSjci8cpA2W0Fr9cqA9IcOCaJ4SmgblFiDhySh3xaM8Zoqfc9lqxNF6cFi/uR2OYSwIcn4q
KEABkFFpYMlRwzOzya+Ecf6vKPWLas/lIxAo5IaWPh5xYGoMFVb1sIqCM72SapH9uw38b4f2Gnl0
1aOhC0t4zEnQffAra6pADdX0/mz+k49J7QC4FVpb5qqRyLNjFILXLY6QCt4cS7KzqHIkLR00FVuO
sVUfoZnJOK4QqFlUAyzCOHYTj5H+103a64DlZ0NVnqupBZD5qwEaiD3iYmwbVqZ9FSyvTyJt1CND
mRkDoxbO/oMpLvTK5eA6+K3+P5rzy8QQKI/TLGiBW4pdvRog/6lyiU3JnuCnTLE5hPoAerZTh2JY
k090pafMN/8AEGeN4ea1bcCe1C6WjpkTuWJ0GVHk9EjRylu4n84qTTsR8+qiX27E22oXAg//8VZ1
xeF/CRbt9S8Y+mOLUGJ4u/EtyIDPSf3CzGScq2jjhUj2BGGaiBJIJD5XiQyAEQ8HNSlCYLaJ7gBE
E7otRJj9c2W3Wf78s0AsxBLTAGKLm7d961IL+z3MaR0+FI6X1Szv3DNObs2aAvzMkKXbaOW3yGRq
P43wUFQncoy/V7RWm+ZAKWeA1u1kXMYjqa+K2z8JL7ILSP92girfi8DwW+jRL8e7f3KSHr82ii3b
dnIzA36DSO6sg4g6g4BsfpoXMBA8fQP8qnNTncZ6ICl915zS7/SfFwvqMARcMOtIDtd/JEmjR9Uc
2XkSa493I7lMmFQKxDvwX9/X69+OcVKkFy0Pe5tH9wU58coI/0XsCbFs263R0cqiIU4rleR9q4iz
LI5R0YgrV4CkSbmmGr9oo0e9P64flNAOwASp/kglr/jUipq5NFLRK9WIR0kajYrCXDXvamcd7aEM
L1m2H/Q2JU5f6NAX0Lr0LN2sksj8L/fEnjQ1xUoJFNhMtVlulPA/YC46xpkNtVE6PW83D/LznSqb
V7/6hYfjhYDflqQ7teJszXhmEcV4d/L4fHB0V9qfTOfB3moRICtiHg10e3HkjQ1V8WwQ5jRj4MVc
/adv3t6ixmESPHon6/7C6ZA5rxiihVRKzXjwgV0pGxvMhZODg4VnS6C3qecHVPcn46XJLyPm7JGz
UWjRVS0DyaegFlWiaWHSyJ5SE4sXH6+DjaL1yEwfGURWo0+wHRnmR5WQkwvI7+KIcFJxrEfDVtZk
OcP6UKelnorIJ0udGnA+4/WmxUNJ/ZwylTyNBsew03IGEMOvkW336pVjSPwfUyHdNp4mMZ3QX6Q8
bzRX1oqkVGwyN0WKM8gh8Ue+HbFBznULTNBeqylgVjDj/8WDWFvXFNBEwVQf1KM+XHE74rFvs2LK
8WCeU6wBxAy6ULeGl9Qm+MISf5ZqyX5vpbNHpWlKBlG0d83XYxUpb8LovvAwyrhvzEFIhLGPElXn
Og8mt5P6BJj9kVbWbB77pxU60+vF3F/fQv9mQSntdXvhF8wyEFei+SaVty6G19NxeAs9NmcUraUH
naaT8a+6GkCnkN3BXqyRB8zwm2hw3j549X8rtN7k44f0+ooYuf51GnU8MEP/MqMHCXy8nzWmAiqw
WSBda9aWsj4uBORzOIjtvdUl8GTNTh3FJ/jgYfQNH5pAHB+2I1sV2x4QKOEqXSM99RTI+qXsDuzG
17CUs8vuIVFxeRDRXsfd2jAND2FJn/VlcBL0v3ySaaGqVjKemFPwOYP0pEcQilRW1GPWTBKtAmmC
pIS9RwsPf9S3qYnjewbtc8BfCiZtlFtDFihq5djXcyzs+4Ya7CYDXT31VBkUbaOkZNcrgVwtfHTo
FaPQrpySETFvCJsKxcXyWbXfodUoRD9Z7oXJxSf5DpaFKFPlnHk6f1ycjLoepMYvwmA5HvMSqXkM
y+NvCxd134g4mq5J/8Jw30Os3WtTg7w7XNjwhZYqqCajsQlQFIS7QhBLOABypGEjiM+o5sABbQVz
p+vF8JBX2RGzMiaFbkZfJN9YTPwO8kaXoazKnBTiQUCUYs9dUMVtqQaYlrsChQg5keseMRxs/dwo
pOVKYdN/RXitGECfvViFk+zqLwfDLbe55ZwBwEKLJnEFEwwsmVzcJGOzCPDp21mEWG2TgvdAA5k7
Op1OUkAS7yIGOnMHvRhfsqzwGTiSdZGjWCeZwPA+7m5jnCU9xvEWIaEnIZzeSOcZ4tyCauUbHsxG
Tm0tyTeMvsOUxQIuauMT5SB0bpU2U3pMpLjk6lKeoRXKIRVOb5Rc+ltVkH1O0d+F4GnC2F8SmBwV
sUMkZ/sAQ7hIv92h75mXcHSupbHDa44zKJtzVUBvrQTaFZgHeVpxzB6xxNf8m63mLRdtS0Qp9TUt
ZOm6Vdt/4jqiay+Rol7uJ884JmJ+/66hK3FwAv+6Kcx5kfaw5fZo/tupz/akPxE6s2Uy7k/WB7Sf
BjzHsL0uFxnKnIX8ZNCCY2zYcgm9mE6OqRgegMXW7oX/1viuBk+CCGI8MwHNdTo4wg5xVCFFDzFI
IaEPl0EjQIOZzN7FW1+AaYC2rqcG7r5eYFeVFy1nFSMopX220FluRWhCDEeuKlPPhVp1twbXSzx4
eTCJTnNs9kXc19rfaeaoKAe4MaUmwgDVF/S0OwzN2FnJ9vd6m7zTrEUacu1zm/yV/c5RltmMDiu+
tNES3A9CTPLJ2Siv47i6xW3dLMkiTFZbPuplYKrwb8NvEhFeqDy9SfUeJOFCYNhtGi4OtBlKQH2w
YoMPiEB3dyLCoeVGqJVocvgeQfPs31hDr9oYXDc5EYFZSiynhkGDLdfnNQ/lly4xzt79J/5upwFC
G/NRZPT0v/CM7llUsDvQuMKGFT7q3jg1EEyfMmH3qMjCbYGY1k0AyIvDWRkSPVmvUVecccb9y2lx
EGYRxM9iv/CCc2YclYvLOW+OIe1NvrkzUgOuJjPDE0+ayYWsg16/3YGlDRFFDKkt0W37WbM72hAK
eRLEuFRmC9g4WTGZXhkggvHxBKgqdPfFEWAT0qvblegMIgvE1NXiNgi0AISSwj248mQlnkFmCMFe
trvZK78IEAYyjLpYnG5CWSosy5t6iN7hCnwlF3GAQseUvTE3zLPRHJj2Z/x/YHsqenhV1jOtm/O6
lefAzNA/Oy6gOCy7Hqtkxt6Ky4TSV2UdvXNPihxLsDQkr4sJ0fnxIO+fC9SCEjfgNY25YZA5W4gu
L5XKOeQkKWwRxgxrxPukT2TqQ2h9IG4P4yqRQufXdjHXNeCYolDPgEYN43WPb/PDhzehTcbGSQlJ
ug0R7AtUYRhxIqpnAHERe8ixA0OeVlNLzHhfGGlwxGodYOd6YGrUan1yzoTLofE91uGi+w6oeZC0
Y0W6uH0Vm0U16z+HtFDAh+Qk3RR4wXO1IDc1sSbXTbXd7b8F8lFWY1Djp+mzuqWsP0fQEEd4xYIT
4Zt+yQ8kRK1cv8WAFbxqBlTA9PJOXsewB3UHUc0WyYKKRc8zDVaTNU6vdPyJxBISLAyzUwsKt7Gr
24ia2aoGOm3JCHNHNRuYIzERGvp6F9ar8reZc1IECTxN5J+10CwYix3Lk2sJBLS/0vIMPA4xFqUQ
6CxHsn/jr3CYlbtTWjkHXwHm2r+xipAO/z5ZWRKgZRgF8Zc3dwt8S7HzwLIxIZ4z6sZX+19Uwe2K
Tc4KgKjrYrnbAIKpRQpflXbnVekKQlzOb/4Ob65mT5AxUuKJF1WzZQx0dNyutawPXST6xdXBru0u
BNuiqIEHajKxpzsVP27DCA4ttJWl+HxYl6SafdEpqVhQi6QcxwA31zcib75oKAFByAfrQz64nmho
6SHJj1aX+LM6s2D4TX8KucxhVx3iGpLXSDtfecAJOVVXGTc4kX+5yKDNd19Icd/bFPDYe+M9fTT2
WlqaQSNK/Bqr2yg4szB/dsdg0HxAZ5GRYA3jj+nnie7C1m7XQxUn4sWYzMtQPFZiIcKDMmu2TINh
3uc9e8Vdtdx6X2w/XQTYLgybkC07BLyx31TUDQEhopH1/8jEq22tYjPO2QeRkBYoztaEcCW9uRsm
K8hhc7ILLWRLjt7iGqkn5eghbyKaJZ72O0m+mImdXfwpfklleO9yOY4Ptdv8ESq11ptzqIOabo2Q
opoPbVDJWU7pagCQJ6nx0Z4luGOjjp+2mYR9PqVp4kA18KwGmSIpG0tY4eyqnnhgLeY2sZ1SfuvB
r9mH7n+9u9cn/W1KEoaCOepRFVzwvJG65HbzYRzRFr/xOByYSepCgF41BlIPRLu69kay1Y8Ydhib
+I8D6vqdqAExt5pA8Rv2yHpTM28LO17W3EYqYwUagD61gmilO6W8dscVu+sMq2hHE7t787tBrkbg
+b5ySdWStYzLTd7msMz7E6UQl45UQ1Gv8+ctl9OWb8fc8EWLypWkwSwQ29pRPZ2cyS+zzrawxZrR
O5MAg3N4r3MysUqQlvKfMginHHLrLA8neLCQoqDnpf8wtKcuk9fRA/xIcjJRA95SY+7toh2c559G
VLNLSZW9AoJID0m2SsabluTHLRx/ieYW8SLS04pi3YSU0R0OKLK7nW7nV3mbg1isdH5qaekpQWUm
ZOF3tJAJ5yqOP98E8rC80Nqbe1SpO5EFKrM3DH4SwBgc42dHDxPGXQtLo9G/yWsVTUm8uHBynBTP
tsGLE3EFY1AaCS2tkEDHEWd2xW3kIFSB5zqguQSpjqKV4esIL0ur3KkRKhM5dnI2DdULQrKCua2r
KuEgGL4JN9B11LrMLShojuGbhufxXSkh9rMeUe20kLlzBNGwJ7b8WXDPKwY8VrnC+k3IHreu/+Sl
3QHGNDoHKg3S47LOQc1ysAZO4hMIcBwXf/YEpTdVgS5EoiusAilfQ51BJZtt/j7pU8BIKzUygcar
zmG+nwu8N5xNjcoJDBrWKgbI4ESxpTo60vEygpoASaaabnrfyEt2B+V7Zv9QuExweP6TZ+u0fo2d
juUk9qk4mBAtkKBWls7pgW9ghTAgumSqoKH5QYSlvi7krU6eQxlc/rGG4dCLbwnp76pje33wJ+nv
TD2o2TuLMD0QN5lLxyvnTZZyKX3MhH5ieAONzMNC4zhFXrYdGg/GdldS9n5pbnj9CvPwSko3QrZe
ycm8VF3U4DW1SulWW6vC4B54ISeKSmy41RUXdqBFswfexlpi4OW187XSENEkaEzpe/UK7VP45tp4
HgYClhSQ9JDyYsMMqJD8/U33WCZN5KydJ9YUQPZ3p91VpXNJOJv5SL7EZGdq81nk81+7Xxxjo2fS
YETgLxv3XQDY5G/TonvyJj6YKZaw3HM2yQtYaXz0yy19vmQbytbn1dJFvcvC+F5XOHD1OAumbDyZ
Bi6lchEghBlS3Q/cMbHcUutwt3BXPUKaad8Lx5wtKH61RjWUTsCkyoLtBtXHFVJs/kG5utzi97va
nV3ZmhwP4O3xJgY6WymLi29DTiuUB8HsGzAu0tb96zEft3BN/HxiD+PglOiKSm+y2Y46uwiTr2t8
UcUsxDXmNs1Yu1JBg5UqP6RVUFPt2ZUeLtMZL0zGZ06ihe14ra4ByRX4+tMbqpCEII5Gnm/Bmeh7
Y5LIIUOk2A0KFxubznkeDI3T+VQGnffzkyhmhkOAUa/49wJHUCoBekAHEV5AIq4WFUdMm5CpB2eg
oulUwJCR4j+okZi2NtdFIbCISyCT6Wz7KLh6XT+39NXHNEwtUNqSZXStw6gETCYUTfl3er/yXLBg
G5OfqJtad/vYSYcYZaA0ARWUO3YrkylbFkgVZBi3WB+niQgNX7bfQvk6+WBdRpAcyTxPw6+Ps8f0
oQ/2SZzNNigV8KAzZrlwYSXL7DeX10AWTEPSyHGQmMGHpu+0pMtmBr7k8BkwRwg20AgYWkHUWDLk
r0O7bmQPS91vSHk/KduQ0xItGUr3br5rEa3QPDmMZdgP8HHjJMS4Mzeg4mSgLPRZd7PY3WLILStP
WfWg7X8C+EaRrhckhQKvqEB27Kec/ooAqGWcnhv8Sd/LKrtu+DX8YxREboXR4W+nq8l1yobEV1sh
2Cs+rzoHAFA6zCRo7jwfnY+BcvvN4+8vuNr8XRU/C/HFX+KdViXz6DLBEkZ8YoCBMHO+0xQHpw4O
5jyTXjh2IZKDg/dInaVHGgdDYt/tDD6z1uDA3wsHBndYzy7zsAkLBqkKw6m0A7YbRZLt3NLFeKcA
iLxDUXGWoj2U24QdN30WEcWxX1yXJIqI62M6mUEkE9mzenx6ChADxgLoMC2iDeG9Xb1XagaVRykC
lnl1O1G/I0rStZ/ZzcfwsU+C5SkRqRS1hchRkLpGfjFrcu2opDHL5MmlFcqYyCE9XjvZ5TmjZKZS
DIuSfHFBnAHbHIGBeg8XPD5wDXpTR2ik7TZFS9NAPmOa0RLlvdTjPDc/IJOPpBO+vUDBFPauTRpE
nKqe7IVZR+KSHzal13/6hyLd0Q9tMH6XMzYsydvw1CC64a4n2P+GeksBvbM5X5OFTG6eGNSCiFnq
olTlAu3uFLYBmcSHg17OMa7kSfHSPIDKmz0Tl6rQiL4gUq1RoARfkltdi8Dh3/V7icAH6YISd0E8
qtpdRvBh2WrugT0+ctZ/D/4jrsy0cjCbf59v1hyL8Dn90ttOSUtWEwdlWCHDG037ZPWuEnVUrV+z
NRlhu89x379eZPeVFFABxAJLmUHJBFie2hB1pDGpZKOKKrOCqQbDlmTyd6eJPTUs0f/D8XFgWwtq
uDrO8AZl/B5rVbuPl6vh/tJsY0I3m0kbuNVXEE0rBl99kXJ2WsHXPnqRqz39dHaLn+QWShPhTTYc
tNG8kqEgtWXv54pPc0BQMFlRMTKwd4v6alDTUZzO7FW6HSufD+0+ww4JUZ1wHBe1oRHlj3hh88BL
ytPVT2+KRWV3ye0Bb/Y12oLTV4JhkjCXIv8qVTkz2AUBOrgDFNaUvFl6A+/lkfIxpE9uxEs8JxSy
G6xlmr9ufGFieXi5X63z2u5tNnx1iZj3B+60LjDnPo1vXnXfHt3ZA9IcoIWZi4OcChlENgR0/PYW
WEkZ4mkRzt2EV+Iddx2r0xCuT5RoFgjxJ7I399x90On+sJ6Sq79+7eAI2GPLZ1+8OHqD4vQzb5Pk
cA+MEDn845buq22fy0YVpP52cEBfTLkjmmZa7EHUagp3K1OXCyUlDrQNfSKNZHncxObIwdxnQ+VM
5JNocAuAalHdnXk/XoN5rmjFMyCkCcnIXRlpmxB1j9S6fPmKEJSRLCGWJ7LH54P9J0JTBY+ApzYS
V8DnVjoChBm4V6DGuCz4S/TGmfrBLOjG3TgbgWEPWi0ie3FWsrJlz2O0XOI/0897Sj6Hn1Ri/vDF
2vo/EB/qBpDQ74ujZcya0Y9T8MBE1rkMdkUQ77W0Vhnz9FaHpBeanmvBFtSYt5KlMf5F6W7HcN8Z
zp1o9lhBMdtrwDQcEWymKv3p/p9zYYQls040FWfbhn7rX2rwxW5593mxFBUunuFU14HA7PyHnLLI
/tXPxcfaYc46bESm/4qte2hMbj6mYV5Cz0NLdXoMNiBgkZz79Ep4U7W++3wKMlbzUoV6BTTBvIvE
lQiKsTtzfXzXGUj0L3XOIq5drqAblBibxP/kJJOescNf8VkIkHFVuRvCz/H0onAJYtAjkwZJ7fIg
b4+jZjZdWuKyr61MKlwzEUVClDZuPlig1d8SUfmbZMclbLzgxv/DqYHvayP+NE5IVoF6vZvqiiuc
0glYb0FwK+9K71eOI2I7MbJuXFnxbuuMBwc0yfbpDiR2rZljV6Eq1USjnagrfzd84VWzpEoqEyt3
eJJGDIIxka0l80YdsSTZIWA8o7OdXJUqPELzWlNspiaCQx40mk6ViYsW99FOgPpaUjnN3mVyUHsE
VqgBRTgaxC1HATdrSkIFyvTXKLnplm2Nbf5fsZygADa3tmPU+JGN/tHcN9ABZep5aKRJTKz/20xd
xguBGFxt+O6D1r/Wd5qzmjj83CSnkh+6ZK6bJBylgMS0iulfgub/7Ch41/PPm0rDNEoTfnqARoEj
JkLLE2mXEEcnQm6Gas3e0N0tpg7P+YN/tb8dt1VyJwFKyAkhyT7+F078F5FRAlPrXhUqn50IlP5D
eKVsARJwlZ+Prn5qe/NnF2PJYbWUdSTuTnLrd/X1ldEGgMX9xDeuWQJ+3JL8mULcSdsWFtgDxNXh
yNMm+uxBeT5wWj9zFznsugDJggyQclTLpCI1WmrWWWk+ksOmE6UKESOggdLcGd1uzQIPNU/O7JNH
W8uR4MGr1wvtC8WwnWqxajLQt+eZTTM1JjNzPXv7Aq3e4pJthGrhmR10cOuTODYJUE1kqnf9cWwv
pcgS7TnZotT61XCEjK2oyS13M8tPOXBgfm7G2I3KTsiQhcW4uJfXGinhbuQubdRgxOFWjgHmy/1n
ZTkqgW7xucDUzqLR9gvLLLxKfhEjUYawXB7A9KQPK3F8rZFv5bpd5bpNNDJ5MOyDvhGIAJaSKnI1
teo3wJ8+pKMlFpVFGznUrzfhSDQiGnPynrkMZtDDw4jysehRlud/EhVVhzIFkwQIgLetxGJhO8jP
bzXfZFOCgG4ubWpnkWSd8O4GkRGGMMb/1Ns+KT96+lyjfHoPQ0rFr9WLZYsj/2+H/YB6pCoryMka
b8uF+0Pxo06Qz2pfuwfz/o4HRSXOdrCdSEHL77DUJoM4o/I8F1S7iN/se/yMMXoq9EYxsfrfCgLk
D/NiY3UKT0+7IDgezckGY8JyXiaaE8TRxM1aKxeLmza/0a8/fnmJQTO0mMsEyQGsWhf7xfcIaV92
R+sNwm8yizGioTBQriY9flyBssC8XSato2+Y1CtHs2PKcs0MjnjfECZEncwRmn52xK2K2up3/DLX
EgNTmZSAEa7tYi2bu1OaaEdn3Q3Ql0BqCy0lLenFGtQbXwftcMbtJz8t/IkipE/wZxR6u457uNZV
3/X6utRIi9Qqt56HXHAeoIOdnoMg+xccZmOrZp8n0yEblbCSbQO6RzgHB6VhMLDmGOuVdTCKFsEy
8MOTSf2zZqJM9VwKBv8WArs3FEQeVKXPi/NjPy3LMJQ/IJ68Apd8s7mLSyxukP4dng8P+dEdK0eN
jM1ZuEaOI303DZcyxkVSsL222ZuFeSt2xjuHMs+jKWFRz4t0kiAI6CDQx7dajmD98VbXJKP2vJL+
FOlrsjlsU0/osjbPW5FP8b21MHH4SkZDmvs7xZ/jiD9BjPRJT2HY9hhfoKLph9gyo9XV2uN/jFM9
9c07B+A61iK2Yj9Um/q3M0j2bNDyJ1UsYgwjcZwfUS1gJcEoPHfO8Kc0ZDp6gjEh1FOcG/4B/6Kk
/1l6tZ8riTOEkjzrnWmyEYjm7Q7e+3qnfd4dGqWKsBF4CDKk5s9MZOWUZKASu9kn2rb1oQyYggc3
58+a6BD83AlwHdlkONyJWCjF91qv0bRQTxPbb777alxtb7dDVe12td6tL2dkWhiQBHcNFX/RoS39
rWXVjTMWXWcK5z/UJ9ZrXk+mTI2sB2BFA8LTQQmDuLqS1r3msg6qoraNhZAfBJ5ksF7v7SGHpGfC
uBMZMhPv8WTyKAEQGpLLSwANjo6zzoLfSEjga7OJlFwreqT+rqisQpgZ9InDGbjqVQmiFGldwwUA
eUeeahDuPcyZoAITkB5pYjpd/FNtWcDFjxEFBjDegT85Ds3gpxkR0KXeEjlD2Wz+Cz8DdvGFMgPB
uPtnuwg0jxWdAHJt2sVi9o+iTeBv+oYp5JtFaWWnXL5S8BE4IldrxCA6Fu3DHMKBFuDwDEY2Wlci
mOB2oGv/R15rf6eam0RzZRrdQrLwOyhWh7+AfsUiKp9KQLolDBBIfgMHPrC0HCxf9IWFCZt44u3V
KSRl+V8KTl+2IcaE7Pd4M7wTReh3IxKTZ5ud2MojO5j1Pqjn8w3QgX+JOpu/CiMH8M7V+9K+JBd9
+n4w4Riah+zmmW0q0qxYLvOVcfcm00CJ5mXL/sL4qiVypGnnmXk5/Z5Su5aeLhLCWje3nLSaImaG
GtmBz3ap/G52k9BsRzeUj/+0DVTcaX+jSBZHXgi1FwhSCB0Mg8139HlYvz6PVXtVNWZcryFTScJg
Dr/hFS7XsemjAqLkeICc7vCm7DjFvCwIocbZx+eLBjjTDg3VLvgiXeD35/f0WShyAJh6u+7HAJFV
AiN0trRVjiZ5AVJrjsWv5mJhVVjagvrxSXt8pT/p3sA/iAEne4wsPSdMLEB7AjFTjLPGboOQtaO1
RmnRNbRhV+Cn9P3AYAzblyrmkh4hXf+1IVbim5wq3V4aA0J4Ze7suzuL7K+7FEXtE8EgHXdyG+rJ
Q3rShrZhNODGPby6oZevrS2QXK3Lw5rvkhK062aRZd1wS5BbGpDEKh4t4EJhGnuncmXNY87JK51y
4O3cf8hrWsmWEnbJMr0PH6xJ95sI4V7Qor8ckW6bglhllB2X3le/qvQlIzeQ5BGUce4SUBlO9IvI
M7tEgBqFzedHc3JeKfCxtryocNiTRvQ4JBEbHBs09EdYwcJJgLH77vbJvRTIN6s3gsg8pkGZDAp7
qD9QjM+efW295N1npihRoKWz1qD8Av1QiywMz1V+HZfuJ9o6YT4QfHp5U0m2SxAW7QFnHQ0ZfEjx
sozGhE+tSJ1leaG+wGi2QBteN/DEM+3NPb2S7fDJh5h25l1nQrnzDhI8aAZR/RzVSe9NHGlFMp1L
8TgpiolzfL/FJI20uiQlqNc8qyMpSvJcjpXdQeNOR2FStjab9E0+MtfSKwUs32gkCtDiagA1PZgd
gjn4Bwu27AKOerswQ0JuDf93jPTsCw3E6feIF17oxd/HiFgM9sHFyZFYvOb9NdELQu3FUPAU1Taw
o9ccOnBpWlRO7hNmiaqFIH8ipji9WeDILrI65t3V3UjxKOqdekcwuXD6Y2xdApju/lPs4xtwGDFr
lKSP2uivZQvdoNz7cHRO81CJnAGqpzabwqJhBUCdsWtq4s/I+ntwR+/jBSbUQpuKIwPWsoFpXMFk
0btu+uPne2qitFKjeO4nYbkTOeuKapo8zGu2i9sedAhP2Y6HXHAfLyt+MWnA3EWBP8gn5AB1Pdi7
UDLga3sF0YqrkSNHR+ArhdjXfHbMv/FZNoH36T4FHSZScTpXrptfnqELuUesT/q8WF0mG3MqqmeT
cljhRJFKMUqpQAHITucymAnGpp1U9jmKhettFTSqHe0ad4egBcZLgNEicj8hEg8zfl9TLmUaqeSm
UMT9UVJJFpCazt9qzin2KvgdmRki7NrHRApaog0bWPZiIRoN6Ne8WbNe0+ryIdwJUWoqLKHXk9vV
NOgFuUry1OKmY3lUyBIMhLyDR61zZd162MBIQZsdVq7+LZdzdFqmx721gc5MwnsJrAl/qKggtzxU
Amy90OwVMwZhD8hglxl1vAgy7MbytUuc2JzrYqy0ljy2ONK28zbaBwJlBmDLZoZARuATHBL5yl99
1F4z3rGXAvzpd018dtFfTLyklmLqucej3ln2og8Syd+A4hlTvyLSAKUPd9FjKmrb/okE8yjNj3my
Ph/YNlQY6TCAUacI9I+gSyDbMr6evYtF+T/hGv1JOpWh2m/WeYCbLMRLbd5N86tKlrWldWnJgnHV
/8wBF33UOJ6D3/xgkbL9giokqcBtsHsbHLrzhQPb5wAcJXiqmn5rS1WglOmZXCJIBFN5tR0yH3VY
QrYrYMTH74QWHlzk+j9A+gqKYauAWY7rpr3Tx74sjTGVeiPAPd6kckr2R1LZCa3aOsTc0pyp2j4K
FeGWL0FZggN1f8xSXgViV4ODinZ4uk43xu+alzQqjYY7qbGx+GbJQHpgjQDSBheTZhXtan/buEeP
Q2AbqlVvq4eMsvEsjwur0MJ+9KVCk9xcPv1LqI5LyzHvG4xB0skis+GVnR77y3aHEsleZ/IOefhQ
AxfikjaJ07ecLw9h2W81cp2jVN4jx12TzYYq1zqEwc9Tx1qTnmdO+WtXnDDBXzFtdUmE7REihEnV
7bvietEl60RXvwmajGoytMw1WTDiddif4WT/io6xWKqiqgwr8CxknGqlP2NArpEDtcXGERB4xBZi
9e4hcMAe7KLxhLYecBuU57ifOFPdWZ6ocCQTcKKqYx2IepzlBEG31IHgwA13hEfWIADKt+fET5Fy
WJaBlcLzYmAyisvCgKLFug7ms5iCFnIfPSS4b4pXbWW6ikCj4TguuRJb8rE5WsqLaCSWbqypiynI
ASLjDUb0sNyfBVOFeSLQstsWbO/1+5sRekOiEf83tYVazigcj5ZNbl+vd5Q3V2v5LJyqufGkk/+y
NGicJMds6cbbz79Huk0IOSPoj9r5zLzDM6bXLDFtTKq/dfGVeOYHGfxChfNOaAZYR/bKGddmLUQa
q458PPqkbyI0qIhK7w9ZiaQiPPIR4/4TauNSeaJ4aOStyU8eGz8CdcuC1y5QJULXqCIXQucpEcS/
YF6JF6pHXdEGUr0Kt4HW4g05EFCfoq4a879KwK1G884IRSOCmboUci9sJ3ZTM3cEd17WwyZOgyCP
K52gXRXsn5TQFOvDsK/k2WJ6u7VnxrISq36Ru9dYzm93NbsYZR58hQdz/JLRSPy0SWEuRSqu57uk
R61pkKxS+wO/Q1KqkW9ugA8iKhqXgAhmVSvnljGZG24SPHO2MRA5tMMruqV2iFQsm89JsKmkxwVM
Uamg0GXaJJNEApjs+hJ3eWkgGC6BDkdRieEXpf+kun5Ar8jsPRTi6h26mo+nVbp3JV7MRIM0sgKf
9i3QAYREidS72XOvpK15wqk/D2Gs5PRVMJdycA0TOr1tLMR7jsYzPPhOpFCrFBXUHlnxjcZFcfad
DFVKu8praIygEb7ITt1vYl6+HNu7AO/2iP3P2z+DQBdb5XCOeLErT1ZcrILBhZpqHplPvl+3mR67
zEtFrbUcP7pvWnpv6lLtNRsQp8DpV4x14xJUT1ZEeaC79ya59OMbzw/XDKxsDSNvDKW74T9bcXZ2
PcMv4sRmDZ1l3j4MC92h0LFInKieTDHjvvlZOLsQZJmRZKChIwv5GYPstsUMT/ohyuUDkwASFcA7
9HD7V8oQD/Ois8LEDBzLg9z0zHwalka/Kg6pUOYKfRZPTIHWi43uA0NFyUuhHQVr+z4EJdeKw8YG
Z1O40Dbna5Qfh5qa4Knj2kx0XDwrAUIWy8CucRNP5WZlVSmqTL5npAuFi7+TMoMhALHDoUyULs68
UTPYp64VOkDQoUCMHmAzPS526P4JluWODV1F45OtW/TZoPsRvmkeA33Ii/mQkJBYMm2qA/9zdXQQ
i6zXd05GZVZKxWedUf0zV73C6RbFeesFd/b9atcVwJRsB37DGDjJf2o9ZvM/GNaCva1Lpb/maUKd
fuqktZnyc7aLFEg9/POzvppOsbwJJwXa0fpG8yeq92nSdqnORI4MsInr5Lno7oSI4F+RQco8uw90
rYhWSNCKnkY985WJJNW9YLCnEqh8nlo5gOYbikBJ9zKbYKlER80yku13iUdxuut38IUTm+lrBUCJ
4nSiUWHRoGRmXPmqqad+oW6jt7SOh0sksQMrwh6NdhqwBpkd0M+IXQRO6sj0JLnFfeaAYAbPL9/I
+f+OzoMyIGWs9FL5Yb/NQY0yC1T5c9H/b/UHaO6tplWLNC0Kl09tZUoOwHr89CVaQELGvQcPh2ZH
iKxxGNKrlxocGVNQlRdP/b0OyMtqqun1eh33s4YolxQVpJQ86TtbErJz/33PwpBojRpTVX9p80bb
pcm9syf3V2cmUNxONKLuzBotmXdTJBclIYcUGhFBPrtu8WQUvWp6vpgpGKp7W6nn0tNqDvbRsek1
mFCZFBJIsvu2uxvoLmlxRwLUkrYQeWOcnUBweFmIMgakf+r2nnpzQ4MUrLvdhV/z9it28i2Ftl87
DMI+tXT8ZrrigcnhOCjndakVhioi7DwOz3dQD362VgAhR2/Uw1ICKZfdPGLKOpUt3tZK7JJkBeMg
jx2JXX9DeDxJL9cC869/4NJHY+6xLDv+6YF/5ZFQ0GbcbudHJyqn0zQbJvLQj6OHE6ay7wfMWrpH
Iw8tHANL+q+s+FfhAQsxCR2fErC/bLDjECjWomS0odBDFnCUK6BUhtWzBsM5z0Q8HazD07YvjbzG
tJ/J2m+c6qA+Qwev2+4wID98Pqt7lTwDhN/YO04og3o5mAha/9Q7Gs6YZD01zUZ6Rw2hh7HzEjDB
Q2xFpUR4ZPRmpPlKPP64MPxB1/82LysviDVrIUJ5ZmFn45zr6uWS+rNhNMaoPqvdFusB1KJKk98l
qga7J/vC+DZHnErRn3MK3DJYpc+bmE+UZ/1ZrdNtBbocmHxDj0BF98u+owpj0Gr3tKnBEgko4Is2
tM3IZ6qCnj9iXzqmLsRqbsujVyfKFLixz99nu4uQesGgbxvSPOGxU8RadognSPBPYovIL2HOSCwx
6a1i0XGSkRSn7jNKwyb3dQ+vbGnyuo9Au1k33jo7qMakFGkPhkmH7TYCGOMGhE1Fq1iXEadrKjsv
4MShq5efMNsulq8bgtHZgMW77WXl7mHL6Y2sLHAB3BbJTFOl8QSfJASLYburFHK6Kp4rKZ9AcF5O
EQetA8XTAoBHr9JcIvjJtEBrmS5+D1+h/Vt23mbfb+3+FD5sJGZLa5+hz9r8kAqJXHAoNngcPbEb
xAZyNeVrJw3s7Z2oBsbA97OfX4XQq9YNe1+IR/3yyjkWJ7gQ+f4t+4G7j95Oau87BfFyYFjDWtek
w4LMRPAY4reusUJCGB8Qh0uaTJw4SiWf0etvJlusjRcCPjuYMq95RRE4115QWaHR3MIMT4CVGK96
8bGLR2T4uYrWUodhUTLFVl34L2zfYw6Lqaua2JavqjUQ3RFcixfjU6BYNLWbGHsD4oE15p8lccso
iJOQBz1W830aTP0+4NjSSYYVKCwAsbTPg3P1Xg9QbEEG1psYXTfZ+Oetx7ykyhgGXYrImOk67hT9
pJ5G6SfZ94jxvimo+rWdUvCiGTnylWmPnTJ8J9usi6Enos24dfqWC4X0Pb+lA/c8aOVLxqMRHBq1
svD5QeXG6Jp8BhPqMc1Oo8O3SD+YVcwo9Cf3mz2+kI+LTKvJDovcjZd0DVqzf51ziO8TxyvUpGxg
hh84uvwqPoAz57yXDRt0+qbGU/XfvKXMB4xF0ehBPO8FYEIBPvXUT9894kSSsE9EnYZk+yalbhv5
xXVq/unlpsUXSl1A0fVIkDxKK/GWmHrqoCTZIzp0c7agN1mF9r6cX7xs8hy6DOBnPvKFw2+dJZrJ
w0mKWA5puyQxQQYCla+dVA8R1vcjygL4zlKIqUYemgWpbZr3kpaDEKmhL5cilwP/P0ok21Ytre9D
9lDNMJguWWO8qKpqckZPZ1g9B2JINwLr75N4rq+cMUIxFHvH+fjXc1Jv0nhIsPfQLuuBnTM5h55d
38htm/86g8V9R/ICbB+8MsXKk9mJMeZtWAcHxZxkP3LrHguQkhhkwEzZdtz1YOHpFIT0ePMy5192
WGUcKv7X6sD46QsbW2BoE0VOitT7nCkdQUefbaHSDHgKbQ6bpb6+co49jJmAHfp8dOksfIYLk6df
DYGSbwpG1i7BO7DT3ao7alACzk4XSNbIhnM60FI79UcDCWLL5MzmVATbj6SKmNrm/eaq7R7bdwQa
4HhfmyMAv9r/dBmwtkiFQYxqmA2/8SLvOG9kbxTfO3Br4PSJ5O1cFGuWyVP7787rfze/c3CSoo6o
qD0nbfdyW7OhKmeBH1NA6geyG4eKlVBINAXgSvzUu/XtKWMLs78mqUJxpxKFTBzuEjpPF215U3o+
IBPzdwt22VInoJ6IWrgAawwKSeYSGRFk2Xi49bvT9hb7SG8F5UlauMIc8Et3uDRtaOkKezM1O0lt
VuwlsXAuRoaZwjKCQthR172nHmUTJl69hPKvkDizNiZsSBWZJsEJhEcbtk88U/+Dutimt5o+0Mzr
2uMbzx4kJmYi23SAmog2gdhEn0CdEm6g2cu2qPYV7NQPLv9GwcYeoN/IhUd4vb+pTUI9cwThrajl
6JbTJX3pn4qmIj8RM6zxJUZ2wudiKE39hYYaRNWfzPQSbSKmd5WlhUGD0JzWvVXNxowW2DXSuCPb
loqGWYFnFh9vF0PcLrB3gptjP5OVFUGrxyOC+IrXCFHaMEph1Hh+quLdSuBHYekiOMVu/JCOo4XF
5haF+cPOxYBU7CyiWpvKJQQsIyLd66cQ9kCWvpt5DxvLzLBFTCHPmzq3Fa+Xqb7ZteeKdwZCbGkY
uOB0nrpOKzIcCVAzALZAV7xS1x3KqwnFa3pWD3NKvfPJQap+QiD1zNZ39dEIECJfJmMOXoF/yP7E
1jdbfYgsIoCjgl/TZOovXQKQdQlaKv+CcRXYy4xHF1KFSJD86YhKOlDIRMHG5uOv7W7Ag3GsB4Dv
zJA/LblEDUNckioc5lwYQnlvUAjD89uBeX8gNKwkj3hmgt8Sz69hQUKmv4C99V85F1GnTlbAYeEp
4mheGKXOePICbLS4fb69qVKoCpL0qPv5TvyBes0OU9oOfRdVlrinMUvypvwYbB5Rrmh8alXebzb3
qurlpRDzrwJ0oTvyBjm+OholWJAPuprHpxJ7h583BeL6EQkJWrukIzBhWY5wWk2vdFnKETbIXllu
Cf4X1RVHeI6X8lxZzuTou9tm4tuU6uxRFto3iQl97FiL3o9mRreJgf++eTx/rf09jSa3BERoKHEc
mwR4xCtAEqqo637S1v6Q2msb8MESELonMRRvAWI8Dz7nOj3YA/tY1Z7LVsYxHu13RZKr03DNerxK
Z+Coi0ZCK3vomvdUhriSi2P9Jf69ueHQBLcOdBgJbEpRrWz1s90gR8w6QxFl9Xpk4vqjeh8BEHTK
dvb3efonK1BhSLD5ZibMeHxdUTlfEjuInfruajXtOQUS1Hiv3UP8Uw2tJFPT0MnL4P7JdhQxqZYu
cMNU2ipWKqdi9h6ss9r9QD32ZSkH21pX7Di3K5olF39QR6gHcViVhc8QNTwvz0g6CrvR73JGRRWx
u6ld0okwUkuh/rqPxWoFtdVTZ/ttjlbvFls6F+5sU7pPkujCAYfWDUw8sR6wZb6Lag4XfGW7+UXo
ksrMPh6v8RuunjykRaH2QOBgIgXT4ymEW5WGkxu5P9iVW93k01RLtWNFoE5QMySMsvCo4SeBFErX
oqVPnRpiOimJ48SqgzA7+BC2gCB/KRzxi2iJbN5ZOxugH1NjwhqhVanTL0z5p08zm5FKdO9zsxhc
EAOoZxESa0BW0i6vkaM3FerPKxejz03/pwJcyiXlHuRrRkxKSoYd8N0rc2JeP+6u6vheMmAsM5dU
9hBLsmjnF9m/VUfuL+xB6kHHT4qoJA2Vijnwh6FX11avYxtQ6n6xgIaTm7POYZt/c0mM44np13Mf
Vc73gHw1GGP5Iq7ALPrGevzVX8zrfP87RNFbHQFIQDJmacoYkXIL0wpiYNILhBoLVqmFmG1HWsQ8
SesMzW1AouL5CiN3Ly4MsFD/KqSK3lsfKNyTF2XjsUzIYN+SSnNsP7MlmqUsCqupxIgZRj0XJ37M
Z2I6nwKCuJJjmls9MqlVK10pMVB6Lpeqlb5ooVbjd/Wl1sTSR06W2/asjieZR68KwX4FIPdOi0Qf
yYKOa6KSLhzBeruc1tAiw6UvPjqZtFRRGO9dgT8GEPR4n3f69USOu3RBXAQyTjCM7RWk/zhvwG6u
hQhgAP1GvaUnRmc6Ulpl6H7I2k9eYySR2rtlqgE+MvqzyrMl31pOw5nub0vCRxE42fkuf3ZWtpJC
O8kLQX78xzMv/kCD6IWSOPrCut9i8o5j0uDYH+eONSXTEPbt09FIMt+kzv4SiCzgilYUmlRe6zIB
W1KZgQZB8VhTsdpDMiEuBzh4fWq47ANYBvtwX0dI5kVDu3IfuP7rd8sA23jdOHVKNV/3TNovJW/L
HJv/DAdv0XyMRjQJJhFk+zzkZ8fi9yGJEMkMw9I7s06CqXNXuFMwjH3WI7a+Stq6M1PuN+GsTfpa
u9SjaF0L7XUzE8ZWO6vRFlYajXzkoZRK+XuY7fan7gyJSvXsVaNrGamZOEoQYGV1wZvlu1lbr5MN
TMWDNkvjG0lNJjWdzVZ05SIvbcQ9Y6vo3V538Kw6R51feJCq39ywZNC/TSkKO52pnL/9Xm2nc3ew
zvwslStdx6IAZNRPObGtqtUWwdhMroU25L6C6Z3nUwLhqXFfX1NYjskFAe3sua9JZGI2wQvTlYg2
R1CgqxGqvNl0EQQe38AdM4FeD4uAbL1FO5CzN5j6kTOzB88FhxRcY0E9k6ZPgegjVTgPRykBJ5AR
XlN2GavKqb5W+wSvL3VrrOJwuJcGF/Wx6khDIBkDJXxJUyKn5nptbzteIQuGjPZ07at1elLqo9MU
OG1sKBgsKz1Cpy33XbbQISnYxg9llVR9qHUNIUGxiQnCjDyLdfBbcrIN7HTyAiNVRqqU88coiHfM
9zx74Z1gvJoPbYPkNUDuWf2As0RSV/oSeg9gG+Q+vwoxAqsjZl8MfxfaqpCyptN45B4ppQb6WjoD
8pUlmNGWBf4wGXDQTqB1aM4/r7zzeQ3MOPrbpR4FRUP4CeFGmOTJsRp8SXp3FZJ4SDDGrduV4cMX
7eZgYp0fbCheCCHrJSTQ8AOvYdZssOWypzA7DrIM3GmmWu6YgCKOu8rO4esROU41H7Pur9+DaWba
ySwrLXB85jDuM3nGsWlj71tzVFIItrPEHHTJwxoxvpPCtdXuJzyiX1POiu6m7aqEqr2qGgbLahgO
zG9wwuoxvVaIkpCTtauZsSCCaA6zl+L72ApU8gBK/tGluc2tJIheST9XTndQx4+iNY4j0ByBD93z
8SsYZuO0QTIOihYFW2ivtU5Xsj2LxIsbWIzQNm7pVRh3ZTe/AWebuit9hYstFNsHsvnEdaDx1qZF
pAw1D2nK/UJ1vidOrwTHMEDvBp/zqSJbB7vPepa7GUiTblQGOvcByX2wlHjlqHimRbZB9vDWatql
Oskd/l9y8O3MaVBot+r/U0nAl7kNaHtQ0/50/cXavxXoFhvJ902I++rWhUWx4U3oYGzuPGjHfAPf
iuXxxlxLr914P8PMgAw7Rgpq9FG8J5LX5pCeqZ36MvyBZ+nCBLwwcVvpVX1JQEV17+PxiVS9sQth
oX3eIxBJ94AMn7aoBqW5xvMl1Ev5Es/pqZ4zqWYVJZfWIonsFwfbEr1hxu1s4nx7pQ+MyxCXYoh+
VyTeQvqDJMoQ5Veif4tRgHw1YEAiDooaRIdlGexiO90pjAJII+WqqxYEJgAD2dyWTMhK8PG3X3bJ
DNJJcXqA6d1mJe/MpsZq1IojGBl4KCiW8yiYBwKi+Eiwx3iFkTHnKOQNcNGR+ZIHPDR85nc9h7zK
k+MW9oIagqzO+QvupO+H5K6Nw7oK6b5ItAGtbejP8qOXdnm0obJ/lKjNNGA0NgLlG1MCNI7PdTWo
qiHe3mo0yr/aUyb2IFI8FbQRTgLQZSDQ3b0lGBvWCDxTj+Y0QZ6i1zoLEImq9kYLS3F6rZdkD5WJ
XG7q/sGRNy/2rMujP2YRUuvpfL1mN6T//PmJbMYdkX2Gz8oiQ9KfF2XkiYZxeXAOW+DDkGLzrDbE
K5nf1lNgsHQO+dxCvDudZ9aJbQe1z0LGQpVUODBLagko/1gPdJoMXLCVEJyLOTze1GtD1adcwLgG
1WDqPtHLuw/O7wTid1wunmpBBAami4tmOZkj1OfH8+KWZjOc6XuQZ56ruoH9/q8RjGej4t68U7lF
OLGADhuOJO7cFMzwO+5CTu+NSa7HHztD0qruE+Bh8ZQ3oyBLfPqKIlwZy5M4q4oRer7yPJ11ybBS
3DK0XDi17NR1viz/A4Ph3p2+c+UadgISzlNmj3aODFxpA42WjxfO92+O4sVwk497pf7Pu1kB1A3v
Ia3hJ6NNcCI6AX9S1OoF46E3m5h0CWrN/n+bjNSSaVgwlXrSNYWJrmq3EF6WyHWiWhsiU38noTnx
WvOlYlUjiHyWfDpplyhNOpVL9aj1LHzMutmVQzyvXuEjixavr/gFoHTeQpABoQkW6YZACw+Qkisf
BId/fDhFWr7ocxRPmivd+0eMGOvW9duJUAEfnve7BzbuWtxwWzaEkBZ5QwW0QFZuZIZT7PfBf7gE
ttDcnEpq5oOzwuyhDUuqLYfekLFqcSuyr9EY4KpOhKOP8nb5YD+3Mgj5gU/t6Ruerygd44aTa7wj
SHgirs+4ON2oOfhyB2z1xDAoR2QC5Rj4InvIqJlBfffElOGEx3nsl8/0q9xOvSAfdXWHhlB5uBji
olEwPQ9wWsJoWzo5H+2XtuvxSd9ArYkI8FXdADf5Ltv/Iap3RQmYBoe9RrnxAYhJOorZLV/9B2CH
gKTVVLkFYf06ztCZ1tVM5hseOBIQBd1PDN1sKekxkvQN3NfgQ77SnXF0slFa9xWD2SkyX/5eRKpF
uBT3KK8kqRlwSrTH6eb3cRdAk0Uhma8K3lQYUSaRZw3V+LX2Zhv9revX7esY55EA1EMZUz4kJnU6
CjpmZ/571bxms2oCYvX5IVGU6OcxRXg4p0ASl+k/Deaw4irkDCIZXg6w4LsQPQSIOG5IDmp6U6DL
rY4G6cWcvkOKE4tmCwWk+nfU+JvFXfOlhecuJeVUUJZCP6sol4M9YwcnL9pKnkwlYUALk8KAHJO+
/x3cDtdC5o3WoJGCug/6P2CoPOMUBxJyXpkftxPPJ3KjYOf21aZWk1tGba/mAfk+R7iOuvWuzXrf
PjBIEbd/okNMz6Y3psIlg0bd9zGyQBibf8hvZFS7UdKjE7YPZ1NuzUpjhSRnQ/YsNHDneFPwTdPn
p48i1jsT5RKpjQIzwXbjqcV1XVnVH9SE514X5tyPrmahmYszHPQEC/nsajhXul/hym/VLYE678de
wS5oeJ12WRtLiuTxkJiYNp8ZWgpJp8eL0FOLJgZ1C6lmyKVUrGvXkZ3JORAj1UV8PwueBVhtCKqi
pR2gS+qZpXtb7yEjBTRYkmyGhh4qq5rLDcM51WCPXlRAim3vEHZCVOYLysHKwfGfK4xNCdToLgON
skpHCPiEZHZN/XjYAaPasElSATx9MyUNmO+AYmpu7KMy9vVgpYkc2Qrfj4jPRf992D9VHaavIijA
EAir2IypAWHmW+niIMQavpiuF2XLZeB8Xt7QyQ82ElEqWBak1hS1bLXpNTXvgNrxCJRl64ZcTkgG
JOuEEzjtoYSOHPgtIyK18d7449uZnqaIvrg6YMdi0LkdCwCXT3llOQzgcOBD1WB8prFcVKD48W22
E6fV8ByZ16YKLChdgPL2DP1qNfRBZI449u0pekTthPs3ABZ4KMZJxV4hZu0C05eB91xynPHKuiv1
Vx3jD0/HBLF7yH7tPTt1ffEndfOPB0wv1XNwO89s4tceLLu3k5S5C7bdvjBHHZ9RiJ9ya5SAM+Nn
hxmetr5jpPxrrWOqWYH/nfMg5BZ82765TpBF2XQiL6v+h8ksTnbENMKK2tK8tXHsxVf9HyiUl04K
QXg587B3EfY0cWJtKHEcu6qSVDKzlYX7n6HwWsVvamAHKZLKS+0JtkPWbDYKIK9MU8dMzJdm7yBm
2Hn1OE+llr7qVIS89/47/SZLbX9h1gy7H/E+ixRajlt93S1t3amwHpPlVZ9KzrVEe8gB93Z/EvnH
RALZmWNdE6Z2WYMdoJy/glYQuW0pEqcqP/K/t3OQpz95RBmRrk2AQZSGpgf+648jwyjhry07jCiA
CjEagC7zXSazj3m1IDgsyitR3buaNT6Cyyv6/wfBlnfc0KuAyCxV693jjOBvntwKnUGAa3f4BHNZ
YgmbT/iElX8kMDk3WHBlVsfJuXOHD5SgQ3TesQViuXNVQMfqpQaxEglbkdMBfyOMmWmMhZwdP0Nt
rcU1HfCv4kxwxbLqTax/kg8iFl9+D9Tc3pDWOS4ccvWU+zKmdEd0yy86QvoOwlSfMnqBKfFw+U29
z71dld3YnRSUGg0KrgoS90UZn0hDXAQZCaKiQAaSgEJxeJHe3LyTbfIl2/68ncQIuj1TOawAV5xz
O3apmAbJG0rOlYDLeGCjQEWoyDbl2I2cOarAJ6mBqCKWKd+G6xlzT89Gj8IfND226kmkuZV7iPGr
UOUp0wTwLHaVCIhUN1YKt8xrq0JC2IYxwHse8Ui9aqoY8job9ehCqx7VZdAZTS5lm6oQYs7CIGz9
KEB0WgS6BpA5ljtAA4Ldi/mKKf5C7dVpJqEmN3H/yz0NfOGaO3KtKPRdfSOxKIjwr2yLDXZZ7yjt
2ZB2m/lFsdGXEk6qH14aOlSONi/3kMenZf7lsU4pzPARtcjZRFJAeydGXxdI1s3yCVqJQUKzJ8IM
O8EUGhjyf0m3/pFTlRScCF+ZSYUWYC32yAY4lzadRpTRlfoUx1L5oEOqQdvOYEvdF1nyOXID9GS9
VebQa9gAlv7MbOwTMD635IPrVi5iOLxecRHIH/8ynjJF4K3KXTHV8DtbtVvcBjNOa9qfrpDA8Sll
rQ2Zl3y+yst7sf4/TvXFx6GHWddteBp86eKFMevjUrez18pRN940C/AZebExNLaXdFiT4/IgIBob
YlgmcrPO7QVcqw8dZPUwgkmD01Unp4fradxgXjaOH3gDsnmudoTvYtswjCgCxALwfkL8YnMnujQS
/8rF7hjAjYZqqCaImvX320O3D1XlC5TwU/o2I4TLk9y2t9TKyO2Ubk9EXEF7lbenvgc+E/LZqEqy
jQ7XVGCbEviBPHtzlTHXAEmqBsx82/E8G+5ABZjbQJ6ruhBE5Wwfowpl3pHYc1MurAlIWfqJ70HT
4qxi/ufeWZjVIkIpXTDH6MR6iyzargAOx0eWPDFhFjju1qS1AFwn9WsRT/ucohM/dKSi2X7oAlIC
LZZwsf4blmBa1Lh9nprerpxQ0GOgcUJ/7B5kMcG5XSk3J4/nBrynwWD1k3a7kd61QEoiB0htfKOQ
pVbq4oMt2azoIV+KHzAXfGPL7/e9I+pFF43qNAhKftZN1AX32AvCWxSQXn8hC9jNfGBV9lXy8GeU
9yGmhuJ0biyEdZm3VkV5EByGyI4C7jqIfCRVZcBN8qOGIn+vJ3CyaDAKAy7T15sJU8p/cXwvvFU5
bazF3R45tM5Kmf3phTC3CEsiJf97G3luXzcnOHhnOOOjUlhF76p0/NcFwnMVimyjCo+NmMLCNF/r
y5dz9mDEgV8iGVQnNJ0VqHCK94u1OhXPIB1mNr92MSqn//LPiv51lPh2jB+hI29R5rcia4+rFFUb
MPBlhWiqED4EgphKpZHHweuWhGP5LlsP1rnQGLGo5c/fJpNV6X2yEIHbUe2PP5UnLsCOFLKWKJcu
23+Q04HvzASZuJEeirSeNZ+V5Mvm4SdZGcJTSylzdZ+ZMg+qj1v3ox7TJqyLQz0cY42/c/V3Eqj1
dfUhUOObQX0+lgyogsWvOxavh4FoULPkTRJ1VY2yxFEuWqw5NiX7itIYIxx2SlR/dYFPZ/MIVHgD
+JtSxENBpKLES0ltFNKqM5Nvk5/cc3SeYlU8IjRQ6WY9+fCeUzpT3jOJPcONcAuP7uCREty7As45
/hFI7ztRrm4pLLfeR/YR92+ifWupE2s/SsDJPY36Gi+0OgeekLZ0OeV1blVby2+/p1Ma7ctu/llL
ylLP+rea/CEzMfsbp3kdaWL9fPLJDQH0E/l22DiX0tGiruvA1vZ4Yy/KzhgAVkALazZxskgnAHcl
VdRqHEwyUP6RxIXY/f83Vyjcj9guVqHo+5sRXWenQqFU0iWtUPK2ME/S/Z9Xmpb83J+e9bHG5RwB
8/UBZ3gU7xMMTjorMlqqhCayEsEfVBSSqQiJswDJ1PXdWjCCvHCBDL3IqaJDpMq4QgumtIfSRLVb
LztWCYUe5s8ix0gfvCgXMB49HLBW72xMpkt3l/qTTNEB+nVn2p9ZH3eWxYlF+g7c8eMIhxOHtX7l
dCroVFgXjs8iecz5qAfDjMhFxFM7W5A7BxfRqtj7Ik6wIyvkpXBytC/eXE1RCB4eD7YqfD527L49
gEz81GMWVPZFlsaBxgFzBiLlohJOmulkwPWS4kPUGCZsFpWff02C415gDrpXW4oKNIZ5+776P2/1
73CQjnTirpMETSlOB+gFue56Na7kE7boaHj+3eP9VJOPAV+jWAgVdXjJYJYnhkVC4FNixcmFGa6n
kIf1eIv0qbdMg9Ie2uoYGmnSX8VLq2dWqZDVZAPwRJnR322NOt6mNLyiuAVNPhiOac9l4E86jrSF
HfFd+6Dh3ufbz7Ujd+NQ4MIOmPND1ux/vLSuqf3Hy0dXCL/AILuzGapFBfAiK48DsN9NXj0ZPEjt
U8scWgCgX0gagOR0nazdmPEc9AXqAjiAOJLZwAzztqSiSHbRqK+kzFg+KO+ptjFm5aAB9PrYjFRP
Cjwc5gVP40qLBRL1xiyRsWD/n3mQnoGymC71UjZTDhiUIAE+K3PZe0NjtJWsFDd8CPS5/Ii4aTAZ
2VyMnIFSyNAJkyR0ka34tGV5Op46virkM0JGTPDk/oxNSkUdOoDE7E5mJ+UevuuckA51rGkcIhnm
TAsZaj6OxOa+8L+yzoHr3vLnMTrD91J12fLrg0+TQmsDT9+9SmuSMdm6SbxWWPcuJVuffo4e0dYs
V7LWPotUByt/zGJ95qCbLKWSWtTZBUFwXedlq212aIPfjXfnQBgGg1GwAJfqyCkqmYhdvOeGzTaX
3cSHsAKDEoWl6kYh61m6ik2SYte/oeDK4lfxHO76BoOm4lzFA1+6juMjmQaGv7WnPIVr9lQpIYTo
PkM5sgiQ2kUeoyC4CqWJnaezNJP6L6AA/IoTgIJy0ClG1bz7+dfeuyGZHXmQlq3V+68/3cUqAUJ1
6MjsLl6AYryxF8KncQKglhoAMdbHCQns5wWHqdG+D9YeavOFT0mojzoy7TvbyLnQOsggh9fDI1zA
cKFNTVh5TBRcHspcX+1a6VoiCNzyWPYr8KUbqKpZas7K7CRAgUPPWaf4i7vT/j4rJptLCMQ7zVul
oNv+nyx1J+A4MKuZfKKaqQHj0F6cM4gPq3QIn7rouSqApfQzz8W3EZzMqTVYIJLWhk3c8eKGd/1v
rjfVHMMYUkmrcBi/eHG8aUYUueKKEjpKHqTFVXVUZoqW//6ne60MEHiGFO8Zw/LqT9ZYEwQvhUCk
XBYhTAjaDGxUB6mHVPx6Qgrum/11lxo08UJdkY85ZKfRbOOY6k8vo4qH/sr5x+wPSosTTBeKWx5v
6iHCXHHO92WxaF971cLEtAH/IviyFBFOR6eXgojhlsWanvT0BbFsZz8CjmkbqBB0Qor3bNLk2OYJ
kjJcVDeb+pYNt0+tiwqj7yXLExaxi80YcUQhzr/WLuS2+tJE1QEZqSRWVGx1YCf9phWC6mcYHrPz
mIPxmrGV0UE1oXd2aVwcM0MnXhNhMET+rrqLrvh4XIUSPcuZbODiCGU6jjs19IAp7ofjIAsr76AK
F5tKb+C+B24S9wMWnTAjHfZuGz92i2AU3N0sKnR+5S+WceuAVsHcEkWJ2JH3jXk1IsQfseULk7sk
p/nG+5Wpgoui5ANDXIB1v7n2NfRC2J+8VZNy/nsHreje3YUr4zZLQDCHdZj7rxduCQLM41FH7vaM
WLzeIFmgm41lfJPA7+ZPBM1xUpsSdMmBnrwRxXmebvaXzqPbIxBESuyC5FxD6IMzLt/zyGAK2RGk
X2+EhV0EmHkBUHYh9MCBZdUCc0GmI0IHKLS/0rSeqchOt1J/LbJLaH66eutcCvs9UoZxBpoA66lM
dM5pvQ1ZhElVcHa2A1rPK19qeFLUDqM/u7am5GoqxsJ4tazY/Uprmun2fk685poWZBygp3IhjLkp
xkqmcwsxfNd0dkViTy7tnRGyCNet/SALz65MGWCmc85NliWLVsWzzNygsyosO0qZw3eZtWTHzwcx
R4mL2EINyqcLdoGcqA/IqysvbXTKvHmMOi3xbGaFVuU5UOJbxzbg1Vtj6/K2iXpwiEBGkixhCs+G
D/0EDnk/NNick5yemu6IA5Hyx0GvmKIGBu6ttX/rjGJLkjDJmaXRTSDxW1N1XE8VzsHkDc9i6tno
tjKIxsEFQnFs36w4GiY8Uk2DgEd+zYmU3SCgyi+wnx1QVwXEZZvFkBOn0wbsVFndRd3mh2qg/mNi
/IzpHW6Pw7dO+pF2Owvj7vTjpoSvyCSsDS+bQmpOxS0B93N3GvTX97BC7EAxsK2eMsTcfc40z8Dv
7jJoL8X8y7P2tRy1EX/u39CePswz6AxpFGl3oh4dUltVm+2cKqcjyuLE+CtkN26r08Aj7ZVXQ6M1
RoVtTxEPs5A37Gcog0SIAQWbmUcqRNK/U/GSUDr57Q17um7icpcep4Lcbmxl4psaZ2kBq3xeJZov
dbkaKEg+9vWwF842VPSquB3VGojNuniOsXHUquIoT068MlyngyxOSRaeZw+KOTf+6/BW+HsZMrG9
JwQaAvTsnTiMHTfXovDCL/MjKCzJFgZRtHAN/gcvsXphRU0BToOHnMxEU1iyDzYuK2vle8zeNQe1
MLgbIpTTPu0Mcvc9EP8SKJkZWu2i+hiCLOsHuuhVBcO0m/KtCnPzjjPTn7q7f1KNiBfSDzKy/aNX
T8dbhN5IzJQXPC/2PxFZfV4rn9WaFZx3F4z7ZeRStInCEkE7CgmZelSQbnYWGY0zpdrqW7Zv78jO
X4MzRLOMikS1y71jxgGWssyPfqqL8aeXDgo5/lRMxpRaVU3ETT/unW945/1YOJyN4Kj0luxoIH7p
/ozEAK3EAxTrkFOeTASBqw1kqorrN0ys5xIsSKDIDGPCO4KRs3qkSZGrSUNXVqgTIV8ODSjZ+236
ZgLqfYhTFiZC175k8Qe6tx50j0NjECIsfp6iYcpJ62U3+ZUmCtkM0tNbWmCkFszj6fLmBk31QJOX
+684DI0dgy07Z1OajWNH8vOOTVu+E4pP4Smtob0rn0KyzNqi8vTPrSgkuNvMf+KPHSCdyEWrLfBq
xkTy/Xvh+44zrhTxuHpmrlql01rD8oyj+YSRjU6WvO1BjynSCWZwlNtj0x2hfIz1yFPQnrLgkuKd
76iznYE/o8jhaFvpfmm43ots6dRnKNa1AIDS5jAzeHGWB5zmCJ2UsjeaCGL7tpKm/pgMonAukb6i
YXUarpkGsERqv/y+EugkDzfk2ukPw8+AA22c7czfQbBjRFCs6e8zvkN/XEKyzV6ELPZ/oYZDqEcn
DMNnalEFwPqbyjR0C9ZvlD0fj15FuvBUJ7vP2CLC3B9e5fqIqiHeCBz5qopxp8NLplYDqEcZAKbb
o5nEpYIHDSadNFSpmASIgReyo9IXrea305TNOGueShv6n6TskgNuJVNx3DH2p9T/ZESdTFiFU71C
+arYki2FM9trsb7hdyrUtpwaLpXKyrMXHD1PLDBslEOVbQ6AWIDiZYmW6phtwyuAthx7bc/Y2ybM
gOnZVqRr3psvO0ZMtF434oMdgY161jIgOX4llqcKDhXycYAI4FLY3NEueJtAF8PVn7PWTi3xW+nB
Xr/xnLYaavjN1cbIT8RjRmW/rAD7QntKMAP2gkvzItQooDb2HUygP+sSoWOgtLfGM14VDdVT5chj
wFFPcdvldalRGBZ+HZzptleBuCBwWodTlIVRLD7cVsdTjKIJOAG+sJWwDXYDCFHP5Lkyjo/6UlVt
mYvMMKsd2PoBBXzzPTUT2v0M9SChvabHSumeAxCOwDDJswIYudPOH8hxL+NMWOi4LNrS3U+6dCAJ
KrlU86/L4/F6quDLKRdAIQyfRsI3zhF3467X7LT+AL4dCdY3Eoe40h7+tbrbuFK7KsbbLJt2B3ri
PZS0aSz7cm4GMLn8P36+peEP6DdvC3iQITz83KxirbdEkPvbvpyYjKL0CVMtYFZDwVU6e35RgVoe
odMd6z+M83/onqGC2HthTEdBOakAUgE3vHxjRDs2+Lk0l8hokbK2RKrpuNBmxK/PXfqBMz8cKHr1
YtWcQ85YJTwrbPA/zhgJXYZ86AZyy5Da5PAg/yXp33WgwWyKViMOFBA7F9KCFDj9Biqxdy+uAtTG
Yk9sQcLrbRwiVZqoe5WgRk6YOQOreWdkq7uMUX2l+6gxa8BOEQLlaisDuEJWxAMBC2kB2brgnsn9
7gcoxaCVrwP3lb4afPVoZsaCyUgwUPYpSta7KJ97PXsu5n+56li/eUXiYMYCcrgQ8zXFl1fcDhX2
T6i3qNW2nRY4i0/VrXKdSIqFJCOlL0VXCop7OknIkZEdKh+JUDqh1K4nPmu996dKa2PhAaGKyEGf
fEfLj6/jEr/0Tj78wJZcbNbUIADq2l2IhjlQfJvboqwumJtFMzOCu/2kr1O1hx5u+906CM6CGQKK
mdyFnO2M8hiSz5DKGDSsXVmUa5tw0AQy1Y4Hjqok8yIJcIQqC6WKj34j7nsfTcBSVJcFgSiFGMm6
Y0zGxbcgK30rQfAleIql593BKsQ3YT9uOeBMLASD2dlKLo/c+HUV7zW7hKjhB10BzP3Hcdq3Tnal
LgRn1W3RHIMWfNSyXdGrCKUlVvqzbKKZc8uK5UPjxRlcEWp2TgYOV94MN0Kkaw8s94U9N/5amLJM
1O8SftU3OBKqG3BejNAZlpcB77rMJWMyppl03BJu8Wq6ku2vgQXJYBCchcIY1wGGRLnKcv2EtVIo
HecCkM3kyBDHALfWzY3Ms8ww2oII60QXDQHND1acj/KvzKBgimZgWPVrmLQmmJ51DUcJS2jVmKEi
TZ1bLuZyo8lPwYmYfB6hKj9/zT7Fj0Mjj34HfNkVG67cHQEGhAwiYUrOU/iTkLG0lFohvTpXCguT
uUOiUsQsCW/CxVFwabQe32vSYB8tY0lVEci6XJ184qBlHTUj7A0dIBNMuBeB9W17B73+jniCWGMb
fN+pzUTmVjuwujdXC2l+Dm28tbmBrhlXLYHhwHJ0cgZnpE6eTvDNgQM97a+HWjyW+1J+UdklX0/X
YrZn0NVULP4dwbcbl1SMSzDWi9FgKB81CDE/gb20Iyykh0+fVruYDtnmXH8Jlgyoz29Vog5tEkod
1shXOwhpyp47ku4XAcet69IYnaJL7nv3E81c1mFquUx/afmFbjO73fIvqdEcCiR/E2/ydBNtjHpG
hySaiLs1ZiZrodoDYlwGL1ZI9XiYIQ7DfaAWuy1ni162Nw+wzF37YUyvGdgtz7DkAERqXqZgwegE
rofQz2PcXXA1XYiIXRDuSC2I+1W+eeQFmUd/pd16cKTCzavdUbMfkdQVNPjVjJvC+xILHNmpLjB+
LYbvAX0QuVnDXXHJFOoxy7sTo8hX3nPje6oJ7tf20OCbycGgC2Ai+mf2dGVxcomjeL6dN1edNa13
0/qZEU9MGbpKogNQUouCWIz9S71ZFLG7ME6DNRb1qXBtazPok1cZXkcD3muDSZ1eQJHf2O4iOswN
mxLTTuwuszWcPElWYFCw4JLxbmuqmpfvgTDGAXInt02+u/hFBXrByZaaqSU2ok2/JDd/su0zrFf5
tsMbv91RLOsgerdkW5oIXgsDYSKAPID4JV3WKc1n+BmFYQCgP7xwM17d2poR7FPA2qmCpd5cqrDp
kYKqRF8V2Uvnp1rN5fHEurlyhXbTXH+mv2amrO9UOjx6VLOTxOjkZQ/pU/EAbOCX92FB5v2xKBD/
TiQ+mMMU43jtUCsUm1TvG7IBpnXBBsNVzZrigDwjdbaFUzueLpG7cyYraMKF+VnW8M6c7uA1Ih72
5uYcIG89w6zGvxgV0HQ9j/iAMn1UWMcANPeU3CzrHVxyt29bAZF9kZXe0CrEwIErecNfB5oGg9xg
tgpAVSA7KdeDXjnWDAC+Iq1VKiIAVff8+4cvj716SgcyXcIqdOEhxBHzyV8WLUjj2dT/KiY2P2un
1ws5w3IatC1jsbw2FPn7rp8cctrcaYqhYRzGFwuD3J8q1p7mocVL4vf9WfAVVwzbmn36wIt7vlgd
e4jxm8Eb+EcD1aZ2JrzvcByKt3j6RY6a9foP2/tUODUsWZrxAcqABJgBY5HAs6H0OpH8zysBBKDu
DUlzTrToBOtgiUya9otrceSWkrGlnkiSyvZpkavbrRfl31M3r1oKaW2k0VkQowdf5LUedUHtV2LK
PyUO4PKKYVRC2gMz+b3ZLT2BLBJWxxLkCTU63l9f5okiTqmCYwwZ8oZoxd9TC8bXnaBLXEsMMF7b
ath3xKMdTP/ukRJ6DfqZUzmE9EhdN/3E01nII8akfTZ8wZLb/FGXTvqc0qlkhdFNzpKHY/jtRUPg
sxBN8bdFrBcnj1xFrtWtJWLxcZmghD3yj/LC/P4JzuWiOWUt99hUim82o2yW8oSUraS+1dHqYEQJ
8e/ze2kBPsiMOBwgvst6GIZhpNQEkxy31SvXHUN3Ybhs95f5TkybgNU3+brGA1vIz9fujrY+yXCq
WxWsxhPK+Fc10TJWtn52b5wVmPGE+V0oETUl/WpT8OEP1kFmlnrDDwPToctDhvLDDwwrqOWsNQ3b
ZrK27tT6JMWMm2/dYZbDlDGromGP3rCyZwLlI4QCpF2WG5Hc+QyZ5Cx7G9fWeTGrFydifpi72XKy
+OljHwgdh5BqfXAKYOlbqQP9d0y3+V00CpzxGs7dmucBEhs/MMNCXMMHEnCM5RCcwoyjkFFtht9M
m91KfaI593WKYicpw+zpLrKYoL6bYZZtSOIKYDr+2ZT3zQs3VEc8SbzIIvfXZOEFk3BxTtsTGTC+
PE7NcKPAka8g4QJRGmBkSHO9hVdUF9443GiKoHLKbg5rA5yiBTHIf3xxLvFYFNzR+r4SeWKqNCkP
aVx1IZgROItJYeLPUO/pDPg+mgV9BRAsqxAvXMNQaYOtPvW0mBlQdyvZecIDL2u0oTUeMNj3Dvkm
FsIzO9PXb2agCDRe77talPRfG71pkN5eDL5k8ZOsBhO6qS53TIfaJ9Ea8jPBiH2QEy67CXRwFQIv
Q+yLBUoB8iYC7G8t4OI+c45YdQjSTidKNuoMhgKyp8tSEKQMaEGTjAaMiuJSXsSCqAh2v4PoReWA
1Hd8ccbeQIVK+Os0g3iwdK/FJPFZDSLmLOw56AlpIWEN+I0Q35sQyUJVPAIEgphu698t+cxjLvzc
r4Kz3n+6ez2ci1n2Z6LtKo0sEBumg8/kIbvt7zXL4v3jwJchjx8rYIorL9Uww1cGUzQlJ+jemRlZ
afQuH9BK1ptqIrpmXuE9irBIs6rFUUKyp/UlIpIK24N7/q+n6aPQ3k+9U9CGu4W2agx7/xKX1UJ5
I5mYlZ4IO7Y4OTr91nhg8sUxpqV2aMH6v/aULBv7UZ0zY6xfOc0FJ142W5WHn6v2N0zTE0fI3P96
eGmDicCUb7L9qZILCiUMVFWsYwARPgovNLMq/Ec3nSTZpkHciyR5A63tArlaqAOf8KzrxOb4jlFZ
1jm0C+1Ld6zfqRfgZsc3tCGhiA+dphC1yOOP1OA9383tn3V2KJpGkuXQS6jYSB42+IahArgEcxQF
y5dfTmoNquZkWH8EHVm8idZsmCCJKJ9lBSr4WPslVcfBWMC0k1Adg/cPIRn109+4jyA7B9HkACPP
wfA0vKgBIhhSz8NzQf/dd2To6DztnJLtNdUA1rJEXxRqN+aBO8G9gPCAe7fJ8yk6nyDdETHbWIW7
yDWYJeSwgx8f2NiEdXtV7+vmIHVV/MbmS/821dHy/vip2FmiVChSnbAQCz3T7E7UjP5ppYOxsoL3
oxELNjOphqPBKwwm31hCnC0ut4NVRyTjptwGrWlVCm14N0ETgddqa/DjGqdtd50+Pw1DcdHVejK0
4kTpLaOKH2jDKi6sxRmr3xFx/iMatIDfyCVXBbjPr+OcUg2ur1S+ChwwxUHAu8sIlhl9wuH637Ed
Dt3zLxLNZbRlLrHL3ZCkx7b719l09jXChBV08/uDktM2SejBiFL06z2PP5WOvdERbuk/5WQ5AJ4F
KaBPetFjG6CitxLccFCKiwzGKganl/CrCgnN4qqy5sWU/k4lqzpR6AySSp3Zyrj4bEtn6J04WCdC
XEwRfr8K2ZUIKxl5+GpygpobC6KyEcpwcfA94s+A928WR0vty3j9p5tPZyS/m6G8usmdFk/e6qpu
S93hVbVD2emcsU6ufPE1CzUd9d6JovWHzUApcCKEz2S1WiNTq7htWHmvuU8tV/4afK418OuHB9Uu
sCbV50npllRr8LBf3pFFODlj2GTgpBMlVfT3HeHQKMrIESPwqep+CixiKWXaJrjlZZKrzc8wbGE7
md/duAtzoaIf0Oik4VcsXiEl/+U9L2m4EtnVp1pwprOPEBSf7cQVMXml69d374gkTveCYngYdWUH
yGWiyFYtR3XkjVAdNLVYOZYQjnNV48g7rGd6k2ns66lhD4xzCSEs8S3QsOsqkgNgUlHQOKHLiq6q
pHfk+2PfHkTIgwwMl97dnOjL4e6e83Wxo/WGfWv0VnvY54E9D566sQrnf9jlRw1MfyY3qFFu92O1
BPaZlH9PIwZZcyO1weevy6Ig6oz0vhiL7aU9e6mJv+Jwo4soSQbpLGt0ZcWRlO8R0i5ADpQ6MNU1
eHCxPcfRPgTVuRuTmudGJbn606S9h6eyxMFADVDGsd+8BC59x1YYxiHuNy2erTlLh/BnvOp8r+CW
aSjxlDlO7zeuInwctiSL0zWakXRRVWwQcXVrVhR9nsqa6qXlV8WebNz7pQxnN4xjQ6dJgOSbaThm
X1Lkwo0orPCLYUQFgyy5bIQmjxGuFyjO/2rIl2vMsYCHCmLYwrh6/ycew76Y1JjRalhXuynOPop1
5ajd4QCS+KUDbEmLxXmARHQoroBENanE4nGrppT1hL2iTgB7quyIvgEBGynj/VI0UNQ9osGu5kPB
y5YeW4EHQBCBmRGTiUwfCc/TY+PG2iyc7bboGb3sL3xHhNxlYB9A/n15IK88cRNyuAwV7NDX7QRa
BInr5hr2p9TVzirS+aU52j+dcEmTh+cH8QG93G3oymzQQhkUeV0b866pwGV5lPn594FoRsZoPLLC
QTng8Cmz5nx9hMTz6gnPXdy8/fSSZ2rb7iOosROdEJVbraEcnR6riOqYSSJKZT6dP9WZnfXIil1N
YxOPSsehPOZ6BAVuooaeh0NgdAS5qVG/Vn9FGjaMfDr8R9NF2455l1DLfnyuD/EGZwV+xP5ltLfQ
Fni97OtM1WCkbdo4T3xPPr1yqWD6bYZxIsHnKZkw67B8xXidhU4xE2jceg6Aq3ro0LYvR/3Rxm7Q
DgID4UIWuy1eyViYix2pvnO4x8aLxBZfuMR2U5mgVFvecjcJyGjfEcBCDWJDH6ZCU115ZHNzg5ue
fEHQ+fG2jYSIOz7GzpmLV7hfRAhBDM/tzMwtzuzsX2JX7BVPSo4ougbTe/yeAaNFsFyj+sNAo18K
8i650ho8UyavMrucmvCJELKX2VHbgtjZ6OQ9JppTbqqwcQ/2RXxjh3dnckxfcxyKGjS+o6TD0MTy
r+vS+grnEccB+yQVEJzboPptHTf0MUWwfPhqwEhL2/ikBa0lO44DKMsJN7g8klc8OBgvpfXg+kKX
tsMRfywcBPmmcZxznCuV97gv6dgoEErcXex2eun9pIRsKno/yAgvTcLz5ksgae7BPwq9cKpQ2svc
1qH9T/1rE0VPaDdUySvdFZLNWrXtwSh2uYA6Oul/sy0gd9XmkwuNhoMYMMVEQgfTCvyiTZh89iXM
1HFXC5O7sXHU6JKpZ/faDTMvjAZGC/grFhfLKT7bwhGLQsLrHKVp7g/VWDJy+Bfl0vyTwY6S33bR
hn5FGZnyYKbFWECC4fstJwpFVGbbLqpOdKaujcJ6qLkvao+H+2X8g+UlURllzueHCTA6A0Qz61I1
oMvcgRpXvObUg0PIDuy3L2yibF37iZB0nY7lrPdgkwBRJrtUQ4QV6iatyU4E+ohG6x2LYUE6MpbL
oqxUcsSwTWCzDd7RVi8eEy3Rui09tKPG65eg7UwoM9rIESfyMHemD8n7Idqif6PIvNDR+MpXoAPl
lpwdyvDRceBv6I+2L+xV0txFhqjd6ALqpxT6yi7JgdLRaUUcToIE+SfCEoQaRH21DNJN/gTBd/QZ
gU1Txl1+vu3W8HcRf8iGUlxHP1e6XWRqI5S99zUH385MO4GjVocDEwiYkMZPSQM98nExJMP6b1LJ
MGkZcsNTKyyuTe9SNwo/yxLg6DGhUg9bXIxuV2FE7XCMNbEwTBrDMhXSuj3Q94q38S1zlM12Ul6p
cFxLToK+ySFYpxXlXLicaZ2lueOL3twch4PBWyBXB04Qg1QaB+4o7E7qfgdSPP69IcbaRfvfXhFG
MncUkSVBzIZyNs+dLzU17rNiukTCFG/VqgVXFSOwp4eyiaAP6KL0Jb8Mnviu/xxxqP8M5DAaNPTE
cMJg674GIWtuyshhAouCoH/4bG97SXNgMGHEaBkObGrLSZUA+0Ig1xjgvcwfmGbyMza9vw0MTseX
8h+fcNNKuLtryXMsud0Y4hIlOlLbJVn2UtkGYpg686YvqThFP0bh93/HyY9pG4tdG0ccRVaj0BJ3
dXwz6Yu67mx1P601JAXXQcndoiW6Jy87l5QpmnZVvZjADxpDLdblCWf7+YA82qrq4iJYfJubf/xC
WiVOxNOVrcPaMGSJBNJo960NZkZfqFqQd853i4Csue0Q6/VqfxVWtHFNWPpLzTMw4DcLrC5U33L3
eXhn7YqixNyeuRfLn9hMkGde9VkDuRgSoN/fROVqewgYGGVJ8r47/PZWyU5/UyfY5XIVzNbrRDBs
7kDb+bXUalg3UQWnX0f56dw59TWCB0K/PRc7nV68d4iwC//DIYy+2t4S6w7xz2zX8uW0Rf3A3Z9r
fRSO409RpUYyiC5GO63jS86uxXRnFdPgXgU+s8VCF4oMmlWlFprjpUJ4kstm9I1G4V0kr9EuARot
oK4kRYCA3bs4QiRsGrMavWkcZ4N3VM4gU+R+n+JwJVS4SUEp8+DIe1XZRD6rJ3Yq+uM/1A5tfESZ
QqVwlIolWIGrhRviX/ckuXYEtGGDbpi1BmhrU0lNVqkBEdpfimPAUBdsVF/3LX/XzLAUkXSD7Edp
QttWkesKv8J9/twhCvw0cIq3JirGhyteEpjzewouRBU2shHH3b/xf+MAoFr1ptTsrMq6H7C8NowJ
ph0Bq0083zCR0yHoguH353oVcMYZf8yJjlHlXDsInjzOpisHhdmycM+ykse2akfvggaoVr24ZoWU
9AM1ZEFHYke8Ps1evZjeu7lXDAejwvGGxGsqCeone7tWBp4U4sdBsLAKGNo4LKF3J3UKRdODuGTO
G6f3LOCpVSyvD8GlVQBEPjuApG3kx2SCh6OejpRx1jfvZ4VU7nUTPnatEFkjvRAOe0MS2mH9+P6I
n8QpiaxYinDTUCZ21+DqVLfeyEjUOOHLJvhP27rkyVAKgRmUjmWOKm+5aw2I/8mOIbhrywlJ7dZY
7/w29oWOQ8c2KDMbE1S+KuXHrFICkxm2Hk8PTQP2ZrwYvusYdTpg/Fj0U/JqjRPwFWYjeyni9v7s
27ATj8PIgibnwVh863IUQbo64JxeZvya+E04G0UfR5ivHX5Ek/yItju7MCeoS8nE5kKqlNqBZGHR
+4doZsDOXAu3kD3C1wSI4juCFxCkQNwNY0gO6Ka9zC+LS1udFOMVYSd94Vz85/V/pe99PGB66xix
IhE/CPlZSn620nmJse1kdltZaXAj5J70OLmQUFgh3CcuUpWkdjN0jJFhCDxWVmGBNXz1EbS2LfQd
Iomh9pZV808NNBd7WmRAAa+ywyhm7RK7dAF14D5c8decD39kk03Zl5L0d76XvFy+WlXzGD7E3Rm5
92katIjFXPB4jrnx+po2ri4a7Ic1JMYd2krNXzwSNXoNYn7jAWau1RLXtUsUozRFzIPSYI3cfjkI
QDjJA/hUHR9/9UpDSMOYc+7AxAf8UC1o8b7PReFyqsY+tPOJwf1yPrhzzcFJtNumeHplcZuahnhX
qK3fJCRxJXH4atVQJF7TKkt53h/y6gJFEr4SPao2bVJGxrPCjyP8+wDrVhVnZ+goTtP+ABTBHJCC
liqvuifcOuhZFIjie1+T0tWgUIuaTpAxH/ZVLfKsinsiDOwk3N9DWNFrR0cTp9HhqLi9aJqpAFpN
ApwFtSrrrgW6rZ4RhjJVdm3w9eOIihLEZq9QwEhDdUyfJQQ2Ih6MUuYy6hSbENxw605RC6yRduqb
4BUGlqpDI2r6Pe9vC+8hZox1DCq6OTPKwFWnCQ2OLwSrkmlXW+dL7truTFp/iHNZrKbwho4o2pVn
mp3edYIxZDVDJkxQlWoDCp21PVEnJWz2eCg+CSaYpw8LZcPaKUDRCW+OaOtODo5bzzxWT1hnJ9xt
8hs+AjzlZJdEhUGRgCqAwLljXdAX7hLqw59rL2fFbQqmw0Rjf0xgqy+3sHIKt0F70IYXv8d17lLG
RgfFOG/RLUhFDx0owniruFUMfZkGrnDC6lWG+up3QKpAzlGliR/5VJZmsPqYK1ga2CgmxV/4PxfN
GP6S9B9IptMA1flzk9QhhmQskvQIt10uNfedtuJrEmscb4nZ04UbJV93UcHPVnY22/lZZBXRhr0e
1dLX4VeNKe0I0tF6T0D9kuxcA0Inp6W6jLKBSPK/VjIZ0Y/MmXUCXoyWo64DU90hHK/yLhP1Yb+Q
aCxcbhCVGcADiRmuLjXw4OyeA1wiMJryyvMWbtbzZ4XZRsN6s7wys6ViFqPGS0BCeukUFlZDGN1C
/UfkHAlsgwqZ0hW74sj/exwwFxtpYP8lXl47yxSxVK4WCXGyfkXSJagouOKqJMV3otukLtqg9FlG
noN57q+pda+RsbpN5brzBMNH42PupWegW2raW1U325dCiNmCetij0/ASWwaVUjRP1+wHM60vNQjN
GwL5wraIg1J9E5vv/jQD71txLPFUpxQt532TcsJoey+WyykrfezhNlMqNTjyCD0zldwBzbIJQeKn
nubvSITSBKWv1cMY529xxmJs+RmsV3Dvl3nrqARJBQOrMO0gPQzW+UC2xYP07VerSnmCy2v7gvOT
KILgLhvkS0jVhCfqU0bn0cvOOCbFzIOMqaCZe6XKofjtIKg6LWaRU3W52T/y7weE+NOH2xLd2iwW
gvxTXt0yLKJCBL8pQWDblsc3X3Bz4mfs2oBbED3OQ9dvxhW8aZMljn5V2UB3Jz4OEcEGcCe/PAf1
vcPPO9H/TVx0YVD9rLGU4x5A8B+gewMK8YA19SrScAOMHGcACmqrRmeD0HAhP6xc9LEjr1VLfQPb
wV66jV5gYYWlddLBckxnkBHQRpvRLd7wKdQwde9XS/N+ZVQlR/ppfTyIocV+rQT06JdrSaQeSeDD
lW9mtpUxmBFT79EnQW6PwykU0k7TX57etWQLvQXgBCVAhi27lbMF20o3bqKqvSUJ/sY7yzojwZ6Q
0lqX2r3c+3UdchcOxssV3U/OBE+eMDLgNOl+RduU5haY/QkXLczx8zHUm2N/kuygvtVLUJvHlH8/
HVG0yWuGzMgpy9lq2bYtnMPTglLoTX7+nvEmOqqTKAUzpujUto0OtSqbk+6AL4iS8+ODJbUGyxPC
h2YORhVd90dhGk6HO5PW4UxZTJYAu0IAdM0gnC8PBqWslZT5i34zBaTy25MJuzB1xe3DfVj1sCCx
WFbShy1dlGWu3Uii10uNInopx+QVb+x/8TA0GJGMddx9/7xfxTsStE7KWYgXmpTOuMw2Kr3V/wAT
4ysGa0XYP01d9GdtvxxixSAsYTbAI5u4V92c2/KSgCUPl3E21GXUHy9H5MlRTbVJ608iyEe9508m
rOytK0pK5RQI+OFhtyDv9JhHUQvC5mIF01n/N1COA1vKrQLjFsn3wWWZy3nmKO4IwZ8ptjvh/+pY
CQ7f3uxvR14T1Kwu+MtFZp2sna87B+SYdMGk6BIWeeukAQUogZPaaDsEvtd9GVjKqKMkP4rrYCUl
v9jCkZR111xlQxkT2SZyKgWR3MklFYLSc2tG9BojmchU3WN9NZRkNJWayF8YGYmmKaWCf5Fkxhbb
uBrTntSd9VVyxgethPAY+VUIGzv25ULw7iueVsSAp2Soc3D/VREoKR+xwDm4CMs+8i0+8JDqSDL0
S9mhdSP11aGpYy6YLg0Cj0ftxL8j1ZuIUdFPifi9YMq1ZBrgGY9gkVAOUVBqvsoTlNIA75J8ug6R
KwAKR5F3iUX8AWarez0I3AHTBfM0VS4RGawUolF+mV/eJB6eyZjJ4zw4wf8oVgLloe4RTy2vEHRP
60a+05m22JwzBxohY8R7kogeBq91TT5uMLnRTfs+3C+K5TYbH9ht7N7k5X0qvfhi9MF5uarHdK98
CjNrXbzADj3IArsORTTUsvtjLi4oKjPCyT5+ZR2/ouPSISyu79vw2lgPsGxnD51HK/d9EAiKGLah
Pg1Yxbwtot38H9vk38U8DBxHwOHcYvZU7ClRoFDg4oHAwUDb1t2v3yfh8jvGnjz87qhbkzmom0/C
bZDXSyTMxvTAciHCTUbgtwZ36g2jErTsV2qMSzEHU7XkUsEEgSmmlIzx8+H45/1UXizkymKrLJSB
F0fWiZ0QBBDgz6HsCYzs0knh045WnWs6xgpTCc12DXpXFa21AGb0QWOY4flSygnUgZNfSL0Ah5O5
85rU7jO6HTOG9/JAQ4Xw2fmWOiwribSFDBr/a9Nu87RtpFj+3jjmRhNKdLhYTK5gTu6QnMqxaf59
C6rx2YlBT0x7J64D3+/W6/MDCR29Y6zyGaWuyUELOpfQC0Zbee2L8h3R+B7qNw/8b/WJxfWrwlAC
0F9bUxi0Xczy8SP8w+OeZ7iNjWAXsO4Nv2BiFncAUJKBGLvsh+oWRfJNwXrkftlAL3jJ500rlLcT
k9rSW7tBxmoUbplRNU/s/qmzK0/nXPuW/z2JXHplCq3pVplVCFeyRMTJ3BlJ71jnbEBDaF/DN6fn
8PIJHUnRW2K5hzixFHgix0FrM1WcLYK7lULPRHQBTzzFv6GOYtPUoePkR+k3W7tlRpSrGr+vCqmU
CTcpZk+nD7sG22vWOt1iP4nFGfkW/SEjGh+T1VtTOEv6O3Kk2baPjRjtyqhA+G+17+X3gXZSpQMg
yOx2c0w4gJPi8QTUmBG/EbVkhRUR8WDUYvkerAqdK/fkh+srf86CqRQZCkog2HR1JlJlc1d2B8ez
qvCACKq/TxPjx9TiUyNuilebE5y5QyM3w/MHVDpoLvJulZ6VkT6vDtGx0JPadLvEop1X2JzCpgXK
wBpmSIkL4cJ8Rcw57fxweUxktDof6A0IUfYhARLQOhohoUuvpp2hemj/SfIrU1CnjkPp1GuUDDKH
tr8jBza7a3bPQtCXjD2A1b8de2LC9HSx3w6kqkoPXEslDIQGmVEux1FR1E56OcmiBehHKSqz9WxR
ShuY+oiYOIN18JHx355+AcxBCqw+s9fui7DQWLCEZ3h6ql8fmJdw3so/1ZerQwsark1Z+202p0Hk
yul89skk+R6TV6/xR+Z2h2GSB8Hoko50qtwP8AHIOKiYZ0+OGxZNG3eqkQoxcbTvFPQBidif/SUO
FTL6Xgw3F/3qEupNnr6bO72wNsBWNZl9m/1gwBFn3zu6qt5TL0BRU36mblvt5cGtZ3UUFWjvwjC/
QclyUN5oMyR1gV0CchzQA9svbQ25+cI5wKcpW9BzWLnlabtPRBuvzu+xrWjb+MDUmMptiUVJPx5f
zxDMNMQPkiJ6kTnQz4hi/Rt4Lal8n9Pdjbto8iI6dmHlrBprzW6xlLGKE3PQwS335lXeILwzLVgY
N+fDk4Nx7+7NpsxrcjzbJqZad0CwSJ9q2rLjyVBhjdBpF56wD055Nc4DnoFLx1KeTfPCKShD7qqB
Tsk7N32lwkj44X7UbfuwjagZrTk7h97UbGIxgHTFJiBqIVjaknoPZG9aUNR11b2vS3hHaFJizW9f
sfZ9jPi3GD9EPsS/9yFESb9gZ812Fe5GAzMh2tSIWM6gdCnKRbC/Muitp4mO0ghmFyRWpDBKcFBQ
4ZLDc81MIr1bDZMWF1kYQS066iSeF24W5KOzHeBQ74nKOaeconnnCvhRrtxHWe3hkBBFMKE8qgvA
Iy1y94rSemNpDx+VCIfUseqVsCzmpP/D6nV9DiausraaB0n6wApu/hnOeDOdAswGXY2lGYnLRAap
C2m1FDyxZVw4tZ2brlNWW1mRg7nu/y4z2UJ/1vIMcXuSBHjfQnW2J/Tj0cmJFt6iSxRUc87GVIgu
G8hoctaFVeJhFw6PbKTNpLa2Rk2iihaG7ajc3eXSA56XEiE7qgfXQ7qlx+qBjefG6HQTuwfR3IB5
7LVIsUJ+XxpTC3tXCWpp9NgUsu8J9h/K9LcZb514CSq/TBBkYJhs17tGtBloz6TzGaAhx2g1iawJ
HUhHte0CK0mfBBvB8/wCXxBlUmGByu4ybZYSluz/0/d7qCY7zT796Q+gP2oSScMTuibzz2/Mg3SB
Vi7Wj+gVgYtsSCMnpb7mK3smnSrQ71mCxm3H20qaz5paCRw+qLFw88d6vEMYEbkry48CaJnOjNVO
WvtwoByvfkq7C6FzkgQincoxU0NFoWxOjKsMOw5lv0S4T2MYdgnXDIfPz4/IN31t86/aGy1Dsy9S
m4ROpwRLatUZzpcuS1txiQ7l4ClVcUr7LYQb2P10OP/+YbJsLWuo6sH+xfYn/ZUgGW3U3Cl71txo
kxAJS7GiP11PLTyl5RoGEWwWxWBpzkqTPtSptEMG8BcmSQboB5wKyGl2vMHND3HvPNgtSEK80/8x
aRw4eLCmzJdePFHoffenfb+XyjvOr9OQUb06LBO4ZSSS8sEZftYgGkXJ8NIOjlbbvUkm5IBvDzaA
RZZlon7c3Xw4p5D/ecJBx1sjFlmeDYU8CgI79pBAzrOnPSAyxT5DCXj+ZR6pHoenmvALhhuNmeAk
io/v4QqnXOYiF93WxIasEAuGfntJnAFp2s50EkgNtrqbMx6xSVWmwyLWqsKRDhadWtgp2wkqTccB
gV6T40d4QjxjrPuWxl0oIbzGcKheFkIOlTwjyYtcHATPYhrrWUY6rst8/uJsWfTCkZVUwQA/5TMI
tNWue/qvHKS2Hueb4MBNeYdEK1h4QG+0i4kMBPZwwPsoAVo3oBooZhwZFIUAthjANYnwULSTBgG8
K03fbKHYQS2ZIPq0Kh80e4AThVBSUI1cnLAGnpyYRAm9BgeCkGc/b3iw6byadznaeLS9Wv+Dn9vH
Jr5fgt5RfbElNq9dNBIGaEgTkGE8/tRmPgUfGyNWcYNKtdtIweEaceMqcGZK8gMysAJcFFv18z9O
jDA45AAp/ieYZ2ClkyY/tA7vIKHTKsip2Y1iJCd9EefS1cJTu33Zp8xQe7K9NS73s81iaVFJdNb4
rDFLniUROgv41qKGGLupgqd3dxTlBbGFx2PNjQYmad7LdMWyW4INZCIoZGwI25kcrWt7z/4j+QHq
CPMY6yIKpOoL1+xeEcDg5XSLfrW+L8YYLyjj2ugEvaDrxvix00g1avuRIv3n3fPnO/YaiBIcFqP4
xxCafZskwvMBiEYDB45mRw47AI3Grb6PZtuQAUfr28SDtbs2xjDUKuZVLmUzkxOLMF1FaKJ8yakY
xpXslr5diTxKWQA5jbViNLs1K/v89WqRsk651AMkep6UdeVTTIG9iMDLwy6gI/MdDt+7PlbOMRQM
BfpnkRfp3QCm+4/gdxEbMJ/DZ/RQhMHAmiSNfcp8ryRTm3fsSWh78CkyDGP/cDlMPmQ8a8dGLO4y
LeR3RhfJTjAyfwzaxw8aLul3wdgyF6lLF2lFA2D3mopl+ks+XuWT0RddrpuNtVRQQDR7Y9JhjBHX
qN0+Wt7Dd+jnvuv9Uafgzi4ZsdH4CfYbzb2PKYf/N86GuZywitlcRiKKJfMkH6FNbQC3cRhUUaJ2
aeyq0+mDndGBzivFgm2pUn4dltdjbtETqEvZi+XRy2lqTs/PAzsxcpEkYOwRRDoqfTsFpHC1hLg4
HsWKiJUWwxatqvyZzZqbGmn+SvgCm8lObTtFr9kBSCgE4YZ4fOdBg1n2FpoyUnpugZ233CnDP4Zy
0H+3Gwn+EdjGMwApYuTFhrw+yO2IG1eJVu4omydHneKwvXBn8lsJEuz3pLFlhyVV9s9X4t/FOXqU
qrAzAx456BUTGYxqgHq2lqSK2x6EMJ10p7+0jEVfT6AX5Ezlx6V9Z6RuDp3gDbpJCatMsEOXkYGd
078MWW/0CkuNzplhgx8S118DlmG86jxpc5Uf1ayrSttB5uroIk5qT72vgY+1sy9wUIYCWdUCH+4A
W5mC90VjG/YeUA1SMf5KCDph2nKz1gSurETY3nz3ej6o24Ybn58NMKMTQZHKHlTXvu/tuvdTQ7pq
2uEsPWXbyryuUBawMn4Um+pYUZD2C6nhjfChmRrJGRVerMkvie8z14nEFyJfsrgWkNK0RcWz7FiP
ev4FEmrVbjxJp1WlRsXEhQiIEiZqUkEqQ5495T/VBlexEBBXYD1gwlyjyRqUBRFzXr4gUAS+7mMo
2dzVwbIT5uVEnXbvDDhSw+kq+McUYNenYZfqZQA625bBZA65SapK92OTQqwItHB7tVeNp1BHLzdl
oWFXsVu8psPRvCdLKaYf/552KxfVaQIvSp81WU/CPAcIy5Z2thKc02u88QnXidR8sd83zAbkJl2y
EJrVZDNOzUfDEsSbTvGHBAnfeydyq2NERS/6GPFojeI7ogN03kb0P7GczMFxEPTdzQWgWdCcr1pD
QCSY6Wy+uZD0MYLaNXsfMJLeYBXVkWbPBP1mGZJ+yjGxGPWJWoVU7xF4oPBq7z5vz1xGd1moudhK
/DqTdGqIeFNwyWEyW4CvYBWD4dEGwsh/3rceDc+aaIopteK0+zQgf9ptoXYb4TOew0nXYcdARs/Z
D4mO/DNVO11prmlCeCeZT1NuIR4K7PZ9BHHPiWxieTbQJE+O73OQJI1IcuKbr9kH4bD9xfHB9m3i
Tal71iy41vAsaHlaHVTFcnIG8+7LMOhb2IUqsEoqyeci6QEWYgr1RTgWQkc2bcUMGE37779tsjco
LgZ395YkFV3kizbRmP1pW7An9FEBSs1OjEzkBhYBVzFCcNU2UiYhTmlAhPzzRTQPdY7Bmkw/lxeu
Obr8kMBbPZ/dLXT28v1uiikeCymk/z21WnMJ97LALjRb82HyBUJE8xadaOxlE+d9UCkN706BdgDU
RvfF9QvmATpwbt3e5x+kXbqUVyS68BiF2Ls0jF1xy3efeadBC893YhiskllQfKekPDsuYW7/ONYz
Lq8/hj3sMXWyIlim45ropgaAmMEEoy9tXTopK1+3npf5X0e5mM83xF/VwYmP5PbIiVOHo87rc2xi
6t8Gvu7rd1epVWFBrCzW3JppmVYsT/owZd8a9Ej7wmbBSIvP32F92RXOexkySvOS9Z7w+P/dWDcz
6Y1Xtl013VAlxEoiJRU6HTUgT/jNvnjSljiLET0daMIkS83YbqM+kU/6p4DZxjy0yIhtnffGAFKQ
SDMBQZZRqUNSD2d9pHYXD2fmiO/qJ9SEeq60dGyzVa6sBWAwN5Up/0bHhnZrmJArlbiovlCLOpDG
llIgsmKPtcfGjrpa8F9wUgKT/Sr34TfETsNeDbXue0YWlup8TArALMCk6q3dAIvFrJA/4lWl8yGE
afpEnYbK906XKhQr1zUkvBwNFvyTHKCkgC0dGKua8fxxLo+9LR7Vi+OarFjJ0OtVf4O9ZY466H+c
MusS7Lh4TaKOvCyxBGbZ3utXXZ9+hLlN7doPVzbmoz6gJqFeUbyKiXkyY+XITMlSgYvjq4a9XZQ6
ACulwIoe649qULTrX+dbQm7HKlIUSHlJ/yLMtNR2iuzkxP55Q50opONWHLgJ/IAlpuEh3gp3BG6Q
6FGqUzu05G8yrbO8JR8198ksDLtM+EOjiJ7LxNXKZIVLvuOq8bF98uUfN0veWqrMdv7z2mc4W9lF
dJPKp0YiuSNksEpPE87ZNrOA9WzgP35cqKf2K3DJSmF15Of0wti5O1TmwZ2S4w/9smc9NhVzf/cF
cUL2DY+yxmYVNXAfIAMsbN9G7OBxUInMCqWWEK8k3FQcw8TBvDcXpTmYRi5j6ALRhLewPWcqniGE
ld4wpRg5tUBNzY1IIfvhgQ71xRklQkn3mxzVyPnESqnC4KaxQ7Be1BSlenU7d9GUaqo7GSwaAqCp
r8wgg98aigUyXNntyXWcHjXECaTYIRc7X60/5HM/R4/ZbT7iRnsbE/AF7XP3KQ/8wvfSPsLgM2Rv
0ncyCOulVBOa1dUaTxG7CrI7CwUtHLBGyqvROeRBEUFET9L12tAoLm+mZl5t2bhdMtl4Gs5ITQ8k
qV9vyczEJtty9QuneOcnPv8mkLpQCjVlab0/XasGqB5P/d97KsK/rfnX1nlw7Qvat+nHWDxDSU3c
nU3uWkl2P4oUGkMO4iQWNeQOi4miz4vWZv7sMkqKWmZAeHyKTjXnl8WjXq0fZHpWT0nuaj0Wyeib
z59ybrYdxTI7bJFlbgTqf/4ZZTUJHAhTFG8RT76ToNuOB47a2lJQwOCOac0wbHwNrzADxxQfATB7
c0sST1+rJWEpkYrqNP5c9Ob+dSKdt5rpZpCkSQB8LnwViXOfjhd4p3E6TH0fA5Gkc+NY41RkC3Li
+kmzWJEhm4ROK1wNSG7AfsoAYPJ36x5CLh9Ykc7hxwzhqAs/7QNojGNH0eAYKFpFTFJGAXuf3jeo
8W62QoGT0ZFBgpkcsNen1ElNvkX9TNUwPFKDjjZqeD23lMmAlJe/vUA03rY0vf7Iaz4Phy/a70tR
rOTRrBv2rLSR04ZsQzO+N24L0H5+EMO9ODc/0n96uXy5M7ze9X7ODeaV2KLLl6LCA5zHJ/+X71nn
JHVikCNXFxc9BSdm+kRlt9Q2pwlSnVcHdULw0rKnQdEjfnNjQNhtdte6tmZxsQVdaf1PUup2/Hp3
O0JXlPdJQs+v3PrKDX3GfhhrGMdK/73aOMSy3kmGdTi/5MBkd+82TVmX1LVV7VfZ5drz0/uHn8MJ
OQzEu8EAf9vdJN0tMhUS53PAapTSGK+ClDV8BsBEJi4/9THuZ3Tl/eiao8rXibz/bkNZd9mzciXp
ud8jCTJt40UMsNv09CulNc6Qbyh4Td3qNC2VAGEaNme8xPLLVlZ1Vrlc50yksCFGbaLtxhGVBgGr
BGOZwUc6HsyjPAPZQn4UTu4w0gktgYSBz2KDI1sNNDk/2GiVN+OQ6IhejkmrevBOdnghQf42hAXY
LPjSudqDoAd9jyG9ElW/fLtlkSqquJdvI88gX1JTJGBxCe+UUfSbsi0fgdwTirUdtMS1Uj9GWo6U
0hXD2+Gf7WRCYgnVCE81Db5C9LLwZsvzPL6Vj4z0iQtHlaegYoqCvAyBrktDU2yYibOUEr7FXx+b
uS+8oIHLtngZzs+8deLHAVe4Aac/C6JZrcBIYZKO4zOf3FVpC1sNzQjKGc3sZDzfC+4two1DzluV
Za/yW3Qnjvaex/nhWJEppqB7fUs2avdr/DdTyDB7uaenYn3sX7tJWyoVbsr3KIiGX4anuZn1VTUF
6YCahxA84/j0cGwwMUABzcK81ZFmy92Zk7fPq/aXcMjKJrQGu+BQRebduF1IulOYWzphfIa5LeBd
yrs6irwrgCobMJRfmRzvXOYI/rfMogfPcOY/48jiWsOeUPSak1VLeEOszUu73qWpL8Ojb/zAIqtv
P0oAXYL/8/WLBeaj/fTI8XIkb8AJlv3kxzKK/oDF5qDvgx4vO/uRmx74guGtZkt6tYniSdKFLme3
IYHw/qKrYKCv5bFdMWf/B5CKcmoaIuS2RlTmM5U/wN2PZJARGNjTmlTbOiKnfPj2Yl2KUkPwHY6A
ee3hkWvbIIFSQggRjUrzqDSG1I4g/byMzcqD5+lJNnvGs2XqlvSyud5vVkbxmzoEPvvWvcUnfD4W
2imQFMhLmnDdYbPgPvZNRWAgLgdmpZ0AXkZw3eAg5yoTkPhT38eOV6xKqeHQxyCEIxEotG06QX18
++fZTLUIyCMsyv7Bf4n/yDqcqgEXhHYcUxE/eh0usXWvRNDN+mdi3GGDpNh7bYlMJ7BBqnHC1WKt
8PnTH/dIpiJAx+JGDQVWdKHrHoMr6D5Q95a9kdXM0yFzC1ic5sSlEqwehZf/FaWupjv+ri5W2jMN
TWpPZqeanGQFScbpFnkdbi6QHypYzRkya1dS4khBokI850sACKUTLg3mDFrQUuM9BKQCkI38JVtS
uVfpgluJvjrc8r64KpZd68zN2Q8wrG9JC7izz9iC3qovihhNEuwERW4+JaUUGphJSCUWgkcE+7uI
wLgm+R517LNvY2r4x8pkYtVX2ddgzDumCTP1ZbP3qCsu4ioE2Ooci55MhcvR0PL+4rjXGllZLSqa
6wpbSpKTog2lapMBS9+MoCXMo2hw9VyVhgV+O98myGRSCGsKyzIAZELBcRqFiKXxrS6uIQBoy13N
QcgYgDlE7bwYTG6RKytomhvW4xk1d3xCNdpoyxNjShj6rgG4diYnC3IgBgsvEpGqOfK5cMbpXjnt
Bwjp0899JBwXx5zUk/G0tgxQ8F1BE1pRq18QVNw8BQEMZBqz3NpC0IH7XTy1pcB8eHAffkJS5jVv
TY1cZEPeeF+OJO6gkZ2OfvaTNqS53kzc3mlJbL+lxC+lIIE82PsM35I8x5k2bxQwTASR0sacWvvh
thSSmcpUD7LdQBegGR/496nd0rsT/kdf/xPcrSF4IOn2IXgbfb9WizUTkkr3I0KrvpSL/v+DZQX+
XQyKArq+whaK6MD939nrgwmaRcm7F2ZokC/eOU+jkmMjCt2gRHkTeRfBZoCOe8Daie7/APLKIbKm
oq61wuqb3Ady7rlcY9gpEUPUb/+k37eISvmFLl4wspKH4RGDckL/jPXYv5uQYzDyDumK7qPxPz+l
pL5vkjxdxigQk3LQdY/2ZHrcPc9IKjm95i/prf9Sv+WbGj5BK3WNJzdLFm0PGlIadQ088Ed1cUpk
/8BJ1/M6YmrLzr9RWPMOVUml5VqYqTeJUXGm9sngYw2fZoebEY0RhYU6Ap62ukNA+zJ8SUyvLj8C
C7sTlxNa29UokVPCXJHtDoVBoAZGSHX/8bnovpMzrzjJ5UEYe0doA7JDK6FAW3UBCgSpFQd8qcln
CiFWmg0coTAuq/nqT2YwIhZZJbXd+VQ5xVjckI8oTu3bIDMh2skz2q86M8mutjs0NkhzJTiEqf0e
LDJzqPhRo1NcLKky7lLE3bjpDVUDS1aUptpSTWw40vwte9CWcKPkopcNh+uEwdoUc9Kp40LUPvJ1
f8L4sXq3pwYNhWlJdO/7dndxOgZRrLnZMECzOlm+oCiHJD9e0ga2D7T4/sRMpTTC4s5znbM6JTO/
yiNtwkAWL3gjyWBN53Z2nfJY33P6BNkGNHOwXXcOe8yQmry60sR1loZhSo26tHosP14z428UIIhI
dibv/IHamVJE76NNclUqe0AnJrD90YJWjnWYu1QvhbzLL50lNgb7t+FQCRNSDTT4l9LIeHPE5jj+
BlZgHukZkVSDE+R5EgyZZSfyJRw3frnOZZOevwZ89ImG8RwZNrP7VCubbKZOY/4/RBx0qfDZMnr+
f2BMh4HsA3ZZEtJDZOjK35yr2AyCY2iEZ3JaKkAYfUedUXbwt+S8x9AiMKY66eqhaJpK6Mawum5F
1yxfKBFaXbTX/4xSr69VTdct2H1VmP4zqEaSfdZ/WN5iqTTNP8GTNTnD1McsWs1rzyKuCtIugnxZ
WUEZ2PQWO19Xt1nAL1xROofWt7jEMyZJKqxm2WvFHVrY9DXbM/5t/36edPzZ5PS47qKDjk7Bk/DV
xyFVkXKmz3tN8meQF/Nj0Xcmag4Rj1aRqIt5K5pZv+EFCGAWp65XyJuqT2oebgt0+x62WfW1Grqr
S0B6ClioHb4SJKEhp09BxjSg+UVjIcpWrDMaQXzFJFpwRS2R1wV0oGdG2ruqw1w3o7yKsL0Iw7bn
jm3dJAb9NDRtFtt9L9p6bFvQgotaXda+9sjHx8HZsAmyFvcaY8Z6w5OUejFJVc/P2c51dczVXaxP
QwPafe0+ORIva7q1qryKZ7bgZiqu3OuejcbdObjelDJrHHGb83IEWYZZjyYOjGAg9plOXl1i0tjI
gp9QCYdwtVGlIoeUOujroeBfd+XaxbHt5q/yG1wEpMJ5ZId2Zo45pi51EwM6dSfNKbRiI9evSZGj
4w94LVZ0SWgn5vQiKepsAAQpPcmezbvgvYJ2AyNqO5IiyM7U1qRtXaKKeGiRx17BduiP5/N1AW0b
REWaSJefh4CvEKVHRW19LIDDq4w8TkbskemTkRrGJlggSDNCND/DaG28NTRYzdAkhRU9clXpYr4B
GGYAcAmt3Jty/scmeWeRg7NRzak3OWTP6mYfEJ5ioSpQZ9J6MKvqm/tk5Y/x3U23Swmqx2RVhxRw
NJvY1keXQeanRQUtoYX7J+42CSLKgP5RKRV2/fb+nJ1axMEVc4kJfYhcz8ey3M0zKcAIDQRDxbBl
pKGvxR2lUgnoXEmwk3H+iLJTRJT08EWf7ckdAN3GyebvSFhWYAfAnr07RIN4egCpusBawq2nElEh
3HmL7SnRCkhsGOYwkFoDh1K4ibFFBRSHweiFuSH2/aMUQFxEqMND/3ow044LfKOTSyQ4xwJAPKxX
CIw21CNGhs66N0yZ1rIFHxfKV7yGep1/3dRUiMSk5VaL7aO83GZD1dzz3rLfbRgWjRjN6nhWn8f2
PEOPQpH2/cdwLrLARf3OWQpkGwtkbOegc14VtrRwZlnsMgtRsyT5H1qT6NRopGSRXE9ljOVcwj9/
ern2lhR41qkHW1tgiCPCV+MnCtKK4uIXv46zz7/lzXUulP/0IVw8laQQqxJc9XFxo3UJCYqG36zv
RQASPt2zjR07+maw+e5xUEVGzHcLO/hLXvvGShZPsmrSbYQJbDyLN1vIl1gSgu9OsPoG6C50XiE8
nxboIpd1MtMgYtPCKwbvqNbOR76Ac2+4kwnVW73CXCFRndzbY5tsoM5rrAc4zBMluR+dghjMesek
RxyDyftWYuvKyPzbiX3eQ7G6OLWs4hN3VhbbXrdoS/FHcslCyYt7NRY47y53uINa+x6CgdvyOaVs
0vuV+QLbQogyuVJ7dn0OpJKPLmYF9dxwfOsWSCPT4DpZX33GKQaQKb6Xre7ctJzyO8fKrHmMZOM6
ZKYVlxANPhb8FLT9YGt+e/Gd42LmaFnv76BPe3KZQAjtsIbbf3zybTEfAxXgXBYX55GIKcmrfoHX
UCJ8HKBxUrsoh+93S5sT8dSeTiffx4E1FD2dQ4J8D3K1uWa/mdd2IZwhkoYLkp+wOjpsPUwQIqtg
NDvNQLCv3AJ+HRWEcuhFXyZJrVyCd5mZAbjNZjIzLIZ6ldRojU4OLVxzDC8V+vjwkJD0LXj7iSvF
wca/UTCq25GtXtyzvzSkn8eIwADWufUQREtrQ4lbsDWbXtlldxGCS8X3o9JxEoQERw3AcBhZTc6l
R2Aq4qTsk9LWFx9O196WmQ4Msn3/dus/cOoQVyh9qKtacWyT0X/55P4YnF8fBmcbHsciJkHtmooz
uk1iMjcaxESdvYE253EWsbXWBfnjA8fVMfj5F9nJ57tvMMZwRg3jeEw3woDfx+t2MYPIXj5OjODq
e5kCTAA7AQ3RnAjPsTmEDLan7bu/0UR89K6lZDFpw5oe/IWmW8F2MTfEqyUf2V/Xui/vDz35S28W
5sOQaSzgkc6j2glQxmz7FZDqcwPXRCUtwqL8iXuhHlckrPQGixFkofd7WYeBKmR7bvnZ35tsDiQF
iggU5V4vB1pc8vu+y3ZccQq94E1F43hs94OYw6jAcG2g/tTIkaWCHknzZN4lG7/K4/RZxFGiQ56H
SYBRVTnCSmaIGq5VaFb8eVIDB8fr3joVKCwqLStoi8lXOtYVdTuJFg+ypQgdnPZpLNdl1YK4fd8T
aMhve27t4zBfZgKEtfbwda1NVDm5si+6MlZ1EThAFhVWq4vDyFxnpxW1pEWfC570fhgHr2kVJTe5
YkPpQbQQzEPFD7wIs+DQ0HiubgJQrd6hT5uGVRE27MYXHZeVBTq07GdfPG0Y5v7radJFaLEQPDyi
uqKv2gpMazhVtRKWSLwXsNVqA/vK8efjI07pioXMk7NxN9W3fJKB1j+h2MHNku/6QKu/BHBJ5XrU
ToXGDht+6TMPaq/UZ4evtHJgzhB/a+bV6Yc9KBgmdV90ZfwrBbgOUzPA0wVoZNAaEC7JW2YNdS7x
FzPz7D607IO5tHfeOsTRJA7LtTKgh+rv3pYaViQLzH+wjpbQwH3nBQRcuBEtGFGNJVP28C0nYqf8
tu7xmw+1K++NPIYdMzgTgiGrUQ026eKuL1/lP1PpiBLmjcYlyTYrUpeF0cJSjbOxhod4TTCwvybC
g1h358r37s6lrdfN6q+m95PJu+wh6LQfQ1XQ4g5T8lX6quaG/LDChP5Cw+flGHh1qMgdlBPgJyVT
R8c3f+bFYSy/YWgdPfJdR30uTQvoucY0+K0dpIEDix6i0KOofvV/PESOfqddJxFKTBmb8V7kRPtc
Eeo9iszPb0qRjLpTpe4bUDP+igWaWR86dC3exdDKVgQWkzibKqXjO9OlYP9tqDLx6i/u0XsgEYwZ
6rrgY97RrOUmvIqWaLkzNpan8MTIc2tchJkgXGd3a7dcIWozxSthDeZdNC6VTu0lf9v4Vj0fnJUQ
5LWi2BdP+BUPmIHn0VbMqVJlUVpcrg6gIJB2S/pquegbaaFPbjF6XTBKFR+NO0ynU4bDwXTl4q49
DbeBjVntBmD8pp3GsjE8v/bH6zLjbU4aDhEqqMD7q6qCLKAV9iDXYMRKEPeIXl+oT6BJWg18slHB
sCnsfz92h1FBoqQyA08t5QThoS3yc/LDXRkt42spEqhA4QZOrHBJhQms/PGN6CD7KzTL3Dh8zsr5
RpLgMiDIRmjSn/0a73PvELkQYgT5Unqx+7/NgtcCmxxy/+9jMlpESncOa2yaawPlpC4Pcqz80IWq
J1MmqvP1+NruV1HhCIlytZCJa2DpKt2LHfL45L20ohtrX24LXqLTapiHppS5HiziZdVGyMCayLDj
CO4OhRvaKf3pEXeNNGLxjdoPOAtgYs2akVsQUe6i0pkCk0YgrIooFLmqKbDHnOzjEgPF0TxM45Zx
XyRulf3Ogy955msgYmvUp5Luhy1Zv0eZQttYeTGAQzso75sMK+DHkWNSrF3h04dEFpksXeluVDPO
o76WAiXvTwuUuOxk70tO5ETxw2hYIotpO0RkANjjQf92abViusehVGxgX/OaVZd/NxncMEF408T5
70St+9GM7k+vKI38/X13a55tq84ctgfe3YGQN8+Rz3g90suqSziGRF9Fq+sWrHN7PSEkKElztbVM
np3NMwwqF7DIzvP6dFIhj1pBdumSRvJHDfDsjaFpROe50KXfdG02GKW1ND3AhkY/U9u2Ly8o2431
XoXkQSoB6kR+Qz6mgs6rikWl8Fv8nXNl0fWo03FNy8ArEztltwQFKmsLAAfA0803j1YojFKtVLua
obhHfiVpBKp18TWiFubDQ1/fhX7csnOmVaD8neKf+dttubyN1xe50qgC3t93iO7qLAKYIViz8vHB
SZSPKceX3M/biXHc7gfUTwmCLyt1PScAoDKTG2D2nW8REB04Nf8x5rbzOm/M9+HkupDCI9XGgg9L
lLPL990f0w4SvnXzcL41+VSBdKBCt9gVlPvJtAL2nWQcixFefG+YykjkGWg186GajFBG1MHM6UBU
P0KEgEY2AONoBF4+x8eOfAWJm5O2Jk8M3AroviS/joBgWUGjLSEiFc3AMBCBGKptF//eZaX4yBCj
83xARMwrqTbAd5JWVAYaQ6dvJZ+oYmegTvfXD/Kn8seGh4jfh2noBs9nETOTA2IfhevIQMhfzS8m
pCXz2XcDphz+hIPjQl3TcZY4t9feJZXdzri8nn06jh5UhNOZdFuCfLOYYPC6xOhgHTVcaU5wxYD4
VN43VPLdkosdgI8fDIswbbRar6jYkbC0DzFYxGRD+CK911tUe+VCW26e78jjhpj2YAUMZAY8Bn6e
IThnECl4EHN7ngKEUcg6YejcRqyfs5inz53gBEUEiTWDbDej+QltDyOyyojyN5WIWbMttFjEyl9Y
XAzkpDAO9AW1koDx+qc1FArQvhDNEBTyByAazgOhZxytuEu94czkgU2oT74tBK6QS344p6ygi2BK
i/T+SLf/dsAqv44CsrGeAhiDyiIiyq7u6qearbEijTcVtdmjuNS/H33JZBR6aPxbUN9lx/yv14Wg
Aq6gZQhN/nab0TkqoRmuIrpdlWo5TmDbzF+3zKKL94SgnVYpuKQAD/QuoY0WwSq/VgMdI8HNh9sQ
c1r6xxrzD5vo184Knu+1dLyF9F853yq+iyMpDfgRYCFxjrqUEfXW+Rau2V6C7tjAHZnTzMjG2RU1
5JW7F/wyjdrgSBlwzoKI1g/zoZQRo4cOixlovjNADU+GbFJfNdWkehpPJg5szQx5G3KiUa865iX0
bS5XCgdpHfjtkGdOBNtbfuj2/NF6J8vNFcCQZTXObSh5Ia9TCtsYcy3JrfKfPj+awhxv686k2WZA
6WciwpTGJ3Sd0K7dv/PCwuKGsih3t4w5GeWeaw1VckXA8g2YY8tSOkdyf+0t0itnRyYT8XIQCvgT
a5LYxusCjQcaTsODzhmC5OFxeSEGHr3YYTjp86yZg+SKLO9Tpo+3MVk5Ua2TCnpXs1OEeBYfJXD4
jIrVvw/nxkojrFVUVg52IJXXtIlxlhzDNYNHzGXv3dmG6tw++kKk4CVsx6i+GA3scnJpaIEL9ePG
jdzF5mIGXx73GHvmFpRHM+rz1ODW440e4JznzXrn4SWpeklYENMORjo/mwTcZMCJTnqconr5D06a
N8mLOxXcN7pnhr6u9IsEVgqIqe1lWoelFq2/YYX58sAb6iocajoubtRVgGiUyl+ma/uZO660VOKd
M2u3LPLR3bTKPoa2RM2gyWsxm4gZb6+sjiEDza7dkyY/et0y5bb0gBR27BWBTzKXexeiQe6g72kD
qDbxbmu+MtFbh5WYTVGWM1Ho7hOGNUX8ZMhRuCbEPW/CF1Y576Gco3sBoO435vNbq13mCDg6T9NZ
uYVZww0/GfpAEE415ciUh13iwQw8RnHlRz6hMKePSJt1YzNL58HmDR56ABjj2K2tZ+w1ZDkcGuuh
Xoex23+iUpe063UAfWhOqChtL3LItWbCTrqtErIurDKp7HhXu1TLjQmfo9j4YXhYsq/RO8FUxLu8
D+LHnOpYBuNVIuoAq5SfPRu3fTb/Qe5ZjI92HSQ2gIVh3LWJB2YFizkiJqeC5ki8EgLQIkRjxR+c
bOVKBrdxdO+dwBlJeKlSRzafs/IqQ9DZ1FrgdrJSZTkZ8JB6k9HA+Uf1w8RO8ePLBTJ01VlOBuDW
7Xd2bi2+7tiJhNBuXQdgZqZhabCVzCtH8y/rvYNZR1Hwj5SCrJ1gQLQLS14hgdMwElsdbInMl4Cv
4jvq6TI5dxB5MKqHzKhWrlmOz+21qM1fmcg2ci31ao67Txbyrsa5zGSQsUiCkZPNHl9TlmLmKcGp
LsPFSzxvGUZ5FATOVere0ca4Vj9Ox86bx4lBx9mvuWNdH5oXhGXrDvW+MXl5P0nziYqZCSxzg26L
0Gh5WQl0kGMnn0KdZ2H8dPaGtKSOBuwwc3WVKUDcp0Ag6kq9PsjQj+rKPhJQMcjnetIPyJlTybTF
3z9Mz17GFr4vb4ZwLznDousHvD1Mt7SbdY3mrYV6pNPhVv+2cEenHWeynnKomQGM7DxkxqGtoToA
sJwA7iAtKkifjpIbAluKWDu8mHXLMNB6ggtV0BbpCGJKN7LGec2s6HwXA3qYjEcX09n8E+SH7swy
irfucv/Zmac56206qU3sELOlhK2UH+kGOxc90lfEcrt1ezy3Mfj/uas90Q4OUkmoYi1tgA2ZEt+t
cN8LPqfWkiFueJR4otqIecluKObafGfXHrG0uDWDMzIAxxD+/uIlb0XbSwepuwkgpLj/QxTvJLVf
Os5+dnJ9s7rR0mLjGHVP+159it17z+sn8eYBfZ7eP31PKnOJ71fnShKNUDFRYPlNMq264dGs1Obg
b3vFV+farQbGX6tAIZVC+yiTGqId7vg20BOcuYy6vym7nDfakSETFWfSo10W+RYDJc/y1XEQATof
RH5l+Kzpl+e0SK92QoL8KMKQoG3keRvPV5KDfsbqwct/1Mt2rgujhoSCPKUFKVfyDcqYGACGf+Nw
pEYPMNeQsFlohhjZHbtXi4HSgrOIOws1KHgAfI/J3yjCL7XLBbgJIY7hBT1jK3a344Tw9CNBSL9r
W9pB6hUFBhO6GcDswnCMsy/gQSkTfqZpqsCMndy9fPvDkJnwl/oo1Mm5VccKqxlnflLRf+MES97Z
f9BYK5qFl0EhevUVp9Oxus9OWbBmVIT2Qh9mfWTmWOMccnVT0t4GFVSLSyXHUoCtUBio+ZwEg7ol
cCpXOsG6b7rZ+pBtAhtOVAPC6TaG76F76uO3/o2e2IpJoOaAGog/wWwktzhU7hWM4rVi3d3fXUY3
T9x2GvZNDBXf6NTRGGP0qOCVeyZRNstqB9xF9NuBmROO2ZapjMtn+DL0+cnVymTZoX9MTAuiLfwD
QdyJy3vfftxpflLGkyJxv4tDCQNeKt6s7RZlfxHjOJN7WYJFAO/DtEIsUax3RNep63PdS18t26Hf
zm6IXNGrUluutFI+a8uy7GezPPxNi+ODxCrIbCDciiIVAxw7jExeI/3JLskR3HPqRXdvExEHw6mF
ZLoZOSzbQiOuVxOSEXvoP6V90rbpy/bkXFTfKgI93G2GfZbI3CsqGkfcGJnRnny1yCgN8hC19K85
w+yMZPK0VuRw20Le8X/Wi33MtHDQm4A0Y0r3Wt67qx1tzs31m1jUW2LkNaw9E/+UIxMb5evSXIw2
+g/pUjQ7uo8rTm6WyB1k3TTRku0szSRr1DpUOsKlDe+BY7wMoVXuCEoPqJCBV9zfDLlhVEpAyIa4
qHeggAwyf1wAjIGuv9aOw4Pr7N5dSzeH9PfFA+I67eNCP9uNWBP4QpUtEyUp4yn6DZCIa6AETqZF
EtZ4BveWvLWVJWKZKY9CpDSXqhIT79uww1NX3at4MYfDxqe+FfWhIn16OR8894HYj91XgC3ykv1E
lf1h6iNxE+QtFV3iMRzKGeOyebea273nFTlIImZEs+BBhjsDBEMAZRln64TabylQLIjIVXIM0tFZ
FLllBYrMJLhdq4FXf4W32zLAEIYygAR0MZL4TnY8QYQlsSzYs3IVzJ6qJEw6gaAyE3I3CgRRmsbB
SEvm+iJcwRoz0szpgaydvVsON/VFY5sc5RKmIcV6qYH86TW/8d3/gKJy87vrj6UiP0+JiLOhFlvO
xSooU7gtqGAgBgDLd+V0Xwwz1rh7ifTrDZufeDDTJ4blJ2dF2XI/NZQsnigtE96x2espAs6O8+sg
Tqreui0+5Klnq2vU0uVhwObe/HWiDkU77+cMY3uzUfOgB8hREiQ3x7o2T3ZcLTv0+COl+4mgKwtb
3T8n92jC94TfHteX0Up8C6w8MKCGlYR6G7RrM9sP12MPk7M9ACyXzonUttmf7UhfSH3KC1470DFb
mP1ZsGODIJ1OUv3TO5BEl3pzypz4OOBks24+GRsb5K1g9Jk06EANigbSO032ciO3Ao+HdgVedETm
MGSeLz+I/imcyxg01uRrVKoSUFlqXuwLLJHOtC078hWYGpxA57BKV03R0W8GI9pUYLfPQwXpwNY+
UhXFlna0/rTFYHRSRANy5xHgxzq0hPQZ2qLk2yTJU9GFlvUU5hy8nKgntE6Dgp7Yd/wGHs7nhvdN
5+QrdLPfCsi0jV55wzYLkpgnCj6pPqyxXzt80rtihr129zSYDcCnxa9i/BWwr5vfmdXlq+7hEn4Z
YuqN2d8maPSSmPzgNiwCMn8AFXt9tV8xs8QFl+8Y3oRVs5pzlhmPLg9iuZOzt1HacFyoPfEivM/N
fxgqbnNlepobwDI8rGef71ecfOWUJTGs3QazYdfZ2onbZfT3aJ+QndWwwGTJbeDIWgGJ3OHDYZ1L
a3TnQ+gApyEh2oB/iS3GxHvAepEw11ni9KGvl1OHdDZIeXPUjb3V3hFN3eqOW6sM+lsYbXXTo42F
yiLMJwk0yZtBVB2gYlKfyJiO//tQ2NmgTKnsS2ujCOTsuR5lMN/KtM5Udn574Y1xhiKfFjhEysS/
B4rrSTh/wEmB1gs981JxN4isy6L+W/j6q2ovT87K+dCMN723o80s7OpxlE8uIH4HF3YDB2xgCyro
bz7uHtIYZf2xHlSwIdtVpuWXv3uNw/HTEA7M3tLW2Th/xdxkB31mtWoNAK40B3qEZZMfK8thvEVg
4WMRmO2AB5fyxt99D0qp9Yc4lrTLBBmDN7HPBJCw6n35JWY+SMtqNrZaBgQUu/S5SStPF3HpTr1j
bf73d7RlAmiTwvPG0JrFXilR3lz+hkqxudB68pQzzxxtaEokafKu9NT/jx1q51MEJW67Y0WhzYsN
noTfS8AN4ScghsH7j1utVw0IRjBJoTeLE3HwBeFdl7OzMWP7weYPdXWLLWJSL6smIgEQRhzCyv+O
MzuniXVl/o6cXbtxwNT6g3LJ7EiroTRNcJrTfzld/5+U0vsmKdzra4yFhz3fPoNOHyq5DmfCileg
Q2HHGT7r30pmsfj+AQmwL1kFRXAy8UijQAiJwUDDR9XFSmWZWgV9nquIKUZJnLuOV/3S2heopqWR
0oNU4/sbucSxxT2WRP/r7RXsf5BWlNw95qU/rrIGCQYlGegx+/uSWVun2IEiViKeu+BU82+Mh3zf
V4JbTDpcrRN+F/nNiEYWo0lUTbkbxSdDSXSjVQSo2bGLiYlMl1KEyhg2UX4WitbargHqFUp5wpZN
Jp4iymmMdwcpdOaDKrq+HQZnla0+ANQxhr6t9LuF9ZZ2wBryFKVearjJTPxF1qYf2XdumR/6kSlI
BOkl2OBd0bxgU5cSAJAyzbSEeR2c4MQT/xB0Qyhu+6wpw8/vimhmKpZV4TC5Wd9j49amv5BFRwVh
Byd8JpvRSs3V9k6CUMbJgJOR2KyAdUcJyfuDU7ksd3eLNe2FjcY21kA4HoeIYotJShwoPJ1u8dtz
fP5Ik1q2a0X/myEtzLvgoIA6JeDynLPy1mFTY5a60cgxqdtk6oSqdoV+3tL/cu/MRKtFjqsE4GG4
aaIW2yvEQjwlwPm+qQBS3WeUHJDj0o5DqHz4EvfxEaD0WuN093TNczObw/z4qK27l5VPfVfTk/wq
bFgpaqbT0JT23RJ6w0GbkfI85VpCmfaGXt0vFUtHMaCH+lS7sIzhlvF8QyoQbhjU46C1GO81RulZ
Pj1HJOMlfBpi4chtypmSdoC5PqGL8G4mt84yD4fZwf17JFl2+03ql8zSLrlG2b5KWa+HTMxjh2dY
D0BW8n4aoke77aJb2zzzpiH6LqrhZglTSLcFxR8gp4rdimyTB5h/1JWf7os+ZicJaPLeOr9/q9Bq
XO5RJ8ZE18nvkJA+yuvHfDn5jOX0RZa0M0Q6LdDzOCJoMgA1GfKM39ODlJp+6imVOBUBp6eLgyrg
7F34GcTJPljeT3IIz+agaoElMfdQgzU+UI1IE1SrCYRzfT9Hjqfvgb6HUY/H7HIoD/rvyyBLUTmR
BJCLM8O5Tryj5Eb2LB1p2cczZrnuIWAGwBhwbeLT12YrdDrvH2359eG84BSReadJB3uHWFIiijf9
K7Q+ACTsfmAkX6ZRntpUukknX6CB61XVeGC7d4tpyRg/jGB8kzE+s7boEai72wgupS+ASscsxYvX
Q1VmCD4kJJFHCe/m7FGc/CIESyfDru/3TfSW1izfYAFiCBhBwsaEVloph1q28pEU1JgBuwXTlyJi
zCh9pgp1qBJf594urEcmumLq1rX2B+u9dcBOenYmu36uHEspK+jLtN3FqtVfx6cpqN3L1gsTCCFg
ze691cN33PxydBl/I38+j3hBphB5EFflodW+thij+O6qixOakPMUuRsjfnD6L3yZxcK3IoJ22JNn
TARj16H/QgD1+LpStMU7JAHYeXHp1s0ytGrFBrzFNYJAi20aP9zLOjkvE68DJ64GZuxLIfvZEUzf
r/sQO8Urn7W0Oxj/KCbEwznm/20XiiU/7v3dGFAAoyvHxPLDPvQO24XZWjxjL0zikfYYjHEt8WjN
2Q0HSBwKHEaHjT9kjgmHgd0Po+XCcv/JkFzTlG30w0oAHY+XS94y7Mzchwi4Yy151RasSCqC/pIC
/EFcFJLHn7sC05SCxnJl0aQZ2H7gJGDwRyQmf1ZBPr7IeL5lfVsXPORihw3t1tLMbzKZ3p7NZzpc
Ghd29kot7Pyi/mV479Hh7kR3idOjnjVDwpdF5GFdRRczrtBpN0TEUSxeBfFqVdvn5RczJH8rfKFf
ntvciKKktp9WKSUv49xlkX2Fu+vOWuL55ii4XBUYOl8OW/Ggpd7H5ioS0L+/Mj9keubpO+lL8n0t
+P2g9+xv6v1DX3G7bHr0BWaTLqCC0UN5dS7fuThYCJp5DoR2UotLEUAbQEZDqTpwy4DbuufwVPnQ
ahotJqZPOQbDb5ppM3kiwyrRMCF5UcrfAINPYhtOaIYFkElzI035TTIYxrk6CHLshaKDq5jMF5QW
4iqE3hYJzgZk4uyaPhxHL7ZFJeEudDevO5u77n0kl+V9Tc91gxREFB5BhQIHnJ0kYg1/YVcYQbnR
Y2x0Fn7F6nTPDdx637CG4N3Q89PbOA73UxfF2Pa6krttASnsINs+0ea0q3RPMqHeqwFq+CvFyknr
MhaepYjrHDBSyAvX7t77/BlVdwj6KaW80jJxNi2C3oxvObKrwsL1Y4RIgpFNA2DDjnKsoyRv63a9
sBL8A6CLpfkkjzK2T+fEsrwZ0QSEsKLowKPhFJKZa0O+Ta+vWsfY5O03qsHzcOUM9AvkEOilIJvm
gSet5zvGwIvRoDnWVT1kIqkvtsaserijJ76lC1JlhaDEmbmWDp9KIU+/YW+RveeNx162EFlDUab5
AkBLQv8/v8RXXoQEuYi95aYCJOvXwSQuN5b3+WjqWCZQ+8KXy6yBBHD4TuAXauIp5rHTaESBJoeQ
o785RWFKDFfjfvmVElCziyvcCOqyK45YnncJJoPC8/i3hBygE2xXProxpl7to4fl4KKVNCRiN0yQ
J6quWWvV3tEuPZytF85H24biIAxGLoWtvC0yI//vyLF1/WWmGQhckIVMxxveb5Agqj8z8F81oEjJ
mVjQdm7QTPXd7vt5sj5xhHKazv3T9nzj6+u97DBSidMBHEmF+hFdRuOEd6QrAQSb+EeFBcCIRRrQ
RjBLX5zZVJoNl2y9OA2SJOgJdMEZf4AoPu3+SgI3+mqY4k4huH+riLF4MZ58pIGYrsBDtFCAtGGW
DXEcuEvzi/p3d0TJDsKV+vXcj98+xntRo9dLXz1UHhhhBLk7JuewFCvnO1vrorJdtQf/TDQRjBr4
UfUnZ4vBIMu9BHIQQcMlvyiciIXMlsOsUmuZz+CtVXREoLQd7JM4gy56ajdPGO4DjAcabosEm6Ql
Ruhd+uu/wKYEiq5g3LMGxFUg3ZPaV9ymyWI0DYBEod8wW5vEcibhf30CKMT09WhBHWoOuirswXvl
Xsfdh/D7F4c3Js5FJYYaIzVeS9eXeIx54T3AcJK7f+g9TulqufTs5BKNYOSYUYxHS6IKhLcpqHWy
hndveWbS+ViiFSMfcdXqeZ0vlN3Pu1INSJKTfeS5rswUaRnO6e0y5/nSq+kcErnEfBTjI8PiV/9B
xRnYpxeT8+Bot4qQTDw8kusB8GAWXNhzYxc7ozRKz4FKwaD8QAcDRNb7R1AMViXh3uXjiRT2R+eY
vqbl5iqbWXYjCunCU3XxWa/do2Y1eGG+pZ6Sx9H294eVAIunuBUzvqMO/1WvQQ1NKMSx0sPWtfNA
BLlHh1WDuMom32SW61d5fmkwOoa4HWOInj/sIixQNeBvBdgLulhlnPHPiRBLMzqxxVV21Rb9The9
qhbJJfgvGOKw9zROgM1zbAW3qM6+75W9Ta2PLs9uKA0sFH0YIKo22+QwtvU6eHX5Y1cOJ3Moo+ZU
0gIx5n1/GUt9GJ4ottSKiiiJKx6PLzgDe8YYNwUxOf4X9nqaakyCQ7CJ83hbktLT4dPNqHxDGlOu
HaFmaWqE/yBaoQfMoSNNkRqgSAowgmgnKz4hc0AoKImI4Fz6uWF1gyuOyma1HJAIfl+e272iNF5I
XjhhD7ORDqQ1RJU2VEGONv9Y0GDD2pNH87hX4G5jileinVQNTDlaNmCRkqVHyzTBVAm+a5/Ph1+K
skoKnjBgs7bIR4+fT0iIz504ehsOPPyh7VwxemCV2pFjZGYpI93n4f+svZBuTwlcp8f9ShhgwPpk
GxyH2/3mwts7sOV3m5pvLbj2Ep/13F4Q/MFbnpHz0HKdhIHhZfWCGDWVNN7mPbGTc1ZBbR03NrDV
Kd8xz2mLC2fDI8Tlk9DQYVALpv5V8GZzvAShUWGAWYjaNyUT7qYIriPNDldMXcY9Saom3aVgbVy9
+59r+kEF2di/GDdTCTrI/7QxX2/o4YTEJNkClObdramZoJSW9vcjvt8SjeSLGO6xZ2YRkz3FEh3y
iq34zqxZYoljKk4+H2BbguJmqCKzIgE/vhTrBtxw4fEXwXSp6IJY6cQggGNBVt6g7Yz+wBga3p4E
oWoDNr3sGjaC9LxEbAleS0GgNIQFYX6kGTvU0iT9UWyLubjbu2Ez/DgVrL1KoEq5SquTNS4kTW6o
mlylatlJxgiC/hefLnC+5Q50zXIBVNXrvrTG2uU1URHP7OXNaCYIgKHvGh5zCevrJ3wqDbRc0Tra
2aOqQZu761Z5SXIB3YOWvz8ZmNEcsWKICCWw1731sUfCAlRu9LeGokr64mICGotzlt40QMWQB/rH
f/ytMe6BoFZSkMdgi/l1YJtiUYp4s4uGlKwJx9fjxV8lq+RazViKXQqT5HXx6534Yw0R0cogoHVo
1+bRHA2jswkwiK+pE3iXOHzUdFRCpmQqgaBcWRucUsSaLcxwqvUDxrydm4jzUJo1BxXZFL5OT5++
Q22FDpUxcgBHVK2OT9DOJ7wCgUeACfzgHwLXyLKweOWgOGk9k4VqYCa+eo8Wl9zKJDN1kB6hMOB8
JmnkOj37jorXi/3r+jK2GrDwGx69mymHXVhDKfXpmM6AxW2GyiH+ifRHw+1IXlG91AVxnLK2haYA
Ir/jgAGU+yIcPJqE1T9aErJau5WOGG4KdvYRJFySoa0p4aXRQmw62A9cDtHG99QxVL2EtaVZp1wA
Rs2slrvpP+o0er48O3yZW+ZC8tqx4D+/rmR3t3KPLifK4e176htTdyx6PUuB2TSTn5de/iZIm8Lz
WMGQQveFzlKaYPsZgJAWIFxCJixQ9PNC9jNQfr5roHoR6tFuLqaOF4FZZsdUrK5nN3/r+IyTByfE
tCTtpIHG2JRxLH6G5W6AeL6Q2x3T6FbADPlMYzEcdYkFqkOiwJBjX1rnskaS1hXfbGKwVw5zR1p/
i71zyeHyr2wOFyrJ6/cMaTZD/CvSYVg1Gkt0cnfA3TzbAUuvkvdjmtM89ga62DaiWzXWnw3ZOQX1
555fMWe6BGwc36VdG0PMgh+9OnC3+FP1tzn6Z+EPlvQNQd0yP3sfq831M6J0cTYTlu593djgq+8R
FA7UMHwejijRhG8wvb/uzNA6NeGW1prmkk8IO7KGTzbJyJ3n78dYxej2p5bhyoCNXJf2V+RNhRE6
3SzB95VooCxs/eX3ruhL3Hz5sary2oW31rN/geFDXwo3FW8DKrk8txs/iBSB912r6j36WqNjMpgQ
Cd3cpW39k9v6koSIE1MmJO1QOlb4kyMD0xQCfOZoIKQO5g03Iv3B9tCZ6N2aCroxg1GLnYLIO1Lg
PyVGdinPbH+YaNUtmyH02fNiekxQ9wpCeCLcJeqWJJZqK/KLQKZyvjAzGULPu5hgvOCmowjOs2SB
NtFljp1k990IMXHiyxh2HjJlpLXuIZPCySk5ph1Vlccoy0kKK4J/OjHEHNiwV8l80YWr/e0tOnwI
sfof4OGLR5Q4jfl+vmvkzBJ7P0YDDkTvL2uWtnxJFXrH0yQqgEHIHNxH5w5f0Xi4/2WIFNAVXnVy
8z2OnYvHQM5TIxbMF5Ntgk5s3zUYl4cTw/blvbg1p0o+FMdECJc6apKpwELYC41OzgyH8aJefMtJ
unHm1n3K8oBEsnv+Zs6xqhKJUvvDT9mYv0t4hdSWP3x2z272hXwCw+XinuzeuPkq8l82nTlmZIVj
0k5s4n8MKQZVyLF9F5oi7sHRRR/NaLZsAJriQ9L+0T2LgN+Ml6okmd5BW054cxxhP2fID14Jh12t
3fQkwUb+0G+tty3xAi68eEih64+cOM5UP0n2H5KJgYtICar3gLaxQ7fzaDnFa+56N/dlDbvn3EUy
u0kklURxNJKQAtWJq2O+oJOHVgDzKCVQXMST89NMzUaVdqst/FmXrbMlkrozlUW4iWAwebeWbmTa
kvcMusi+eUJVsB+z3tqDwyLTzoqUA6cD3jFmRBt/P1RZ52wsRgaKgG46Z6luexz0L7Bs3o7cGu7y
JkoxjwSzRWYjv8si1Tytw7GN3L/5F6ZZ2U8PEiHh7fwFvUGlvIa5FLwNGulT+VlRqerKT6weYV7c
LoUYoPR/Twnzj41P+n3DMdyJSw7VSSXZiAFngl5WhTwjVzqbd1H1WNbU518kMv9V0t8uvAo8HW44
icVM93pd1fJ7WaHEv6z7VYVkXAr8PYLgnjdES1xYEzyj9Az8jW87nw6vu1pUm0ckpmIiiBtGQ4ax
n+Pj3ieveHfxH5OEYo9qcjsUhE5YsElArE7allYnlkn3oE51Gbui+cNRUnYwBSWxQRRAYwAMmDwA
tRFXuunFpe1Wj2wghwmo6vqkFcMJ9xhPopYBColtcLBxOUY5lwhsodraoEjYfzi4D6hFKpzkDwX8
6Y6zK6ixc2x+931IhEAJ9ZE9yqJitue36WP6YQWAoCzr+5BZCIH4Z8ZHDIUMNbYhM45aQgC6wQ8k
vVVmNaZ8MdpJwcP2Xc+ADa7gsYipVzU0ndmQodnMOSLxWs9rvaZqd1jkuMZLWsdgrgqTj+Y4LXYD
IkWYNVG0B1OFWXKmmRXhzSskVf+p987/13srHS+wAveUvMc0ZHw8vvxoxnZGwXPG6hYM1d9PmBac
roaCr8y0d93NJFb75tx2Rcz7gxdHmxEYfi0HU+Go6VUnyWFV72P1cz1gwH/JNaLEfyblbyfovj0Z
iPluTxJ6kmUgyIMfoqyicertmxDMFGtmx+j3KijbsWTELIAAoIj9xUI6alTz9uEvMXfUBuXYvKe5
j0Hcp92/hBUrSWHXv1VvZWhUXX4VHEg/Ex9nu7bPH9vGr5vxJ/a3jp4AnxETLJrTfIE8YoCSmKxb
j7+VQfF+Mdi44oeOgJjR/h61kZ561K7IllQ8NysaV5DIwC7OqM3jjID1wBZ6Zm6wjDYOsbQx5b7v
147yk+ffvI92r6RMtRv/kDRM7R22BG2vjD/WZf+3Tc/GBfHrClkR/hgj6luXzfeZqCY3ayWWub0r
vxr9/9CCqTLEdaMjLnWMB4Z8YzgvAIGU+PqpC/vbvINJtPcxc7WvEqMkEA06MNcp6PFvBOHatRdr
5FWIx5DfUZM8c/HT9PJEfMpTmEvK+WangKDawN46iMrVOqp3yGc+I2DFZ/T+LgLPgd3xUMcJHu/Q
e034KCP8z/j0V4cH2VqnD0A8+wlTQjaWQAwMlO0lzvlUQS+YZ01uQOGn9i7oX7ygIFgt+KNTCh+e
9cinv4og2zyWo1hbawQV1zEJO+sxigxK1TaTOKwRuCEwOD4bBUmZ/OWUOZVNf69pVeAg4+M70630
aCRrND3D4JB4ZB8GE3ewKhQR18hJbhT+4Fj4UZq1WP3mUROBskYo2Hk4V/K9ccUA40E5RJC1VdII
3FAXKct3LcEiV1MFJ/eUH2F0mkef1ARnHp55RNoHy2Mpmkaf8oIvtewi74nxI5YwkAblRQhZsPpj
7XJGJd07EDu/zRiY63Q48kmHS/0qKLuzx5gvOywbFBw95acLN6PgwVHznDZqre+qCmJh775bGicf
uCryQ1eQqZffi1ZfiKqiP0foI9EgfwPi8Ho+mayPCt16wzm1wmOIzHJqmqS1zKz/Uvutvamsl6Gd
Lj9stQsJ1JDHUfEKvlo8Ja3uTtLDpmFcEMEfqScK+3b/pxC4l8wW84JA1cDER/HwcmGGh3BGTd9L
Wzv/Rjm7JO7h5uR26rn0wirpK7alfOYCRKwQpc790evr8qaKgGz4wCI8AVlD7YIhu306nOQuy//8
iLEl7u9fE34LwZPPEtORHSgflmMAIx6o2qfSdGCRoi1AZg9gZBbOD33udHm041pIEEskmIdEIhYx
Ev2EVloKWfUCCavNmBA9gtTExerVypsdl1vwaIHsrnBGQnODvaif/q5pRLXOWy40sIqE25LAjB2t
/MhuTFUCJnVZNoDv9Yd7c9Lt2AGEebqD/LF4OafdEpL6YuhqaEEgePB6VCk3ZwB+uCsPebAWLIjv
+kxVD6MY+U8O6f/LHMXf7FjrszJ7QXF6IdId1EGNPbZtzWUkz1oWv/cLgctly9d2vzdoWnP0K5SN
ngdk4vfJvJSbgMQXfhM/ZVMs5hDSi9L5x9cyrtLQEh8A1yomGwJTQ9FKV5ZCEuW0BkU66DncShnc
cTI5IHlIdF9ULV65sFy4Db+Mr2pEnaIpwhCJYDxbE0hn9siBgyDs4a54GEmfB6krrUODzl5Ksy6H
HzkP29fFI4MkneDok3OitwEpXFh3egBzUa4ZBnUoS6WCfApKcRKA+Z9O2mG1RDwE3usb+G9TDt7/
hpAZE053XXcqKOdmdy6Rjg42S4KdOLxCDtQpbjkBEOIAO32leoOFWzEalCdExV3esXQ9NLSKMXNb
CYjwaEVEhiZfsU6Q1suXNvYVAjq4hSGdViCQRdkDwCAE2MzymLjCMTRG+4Ocvw2CQg2zivNDvBcS
wSHDW20itoSnc112xdSmq2MSkZIAqyxQaR9Tmm3Rf8GXbflcTCqLvJQkrMCangDTNaiBCbcnyctN
X8Bn+kfWYi5lJmz/sgpLGlkiHujGeiCNB3kuUpzoNiiZo+phvo7HSrqi7twIMfht7KTsF3oWJfCw
ah7JZyT2MhvwFUMQxz8l1AFa4WviiwFVfV33uR070A9EEVl4KqRUV5zIRWBdGkY6tnMvtvtpkFoc
cPjZUPMpnVBMEQGbyHVjbLdZIQZ8M+tTXL8Z2eauxkVDzLhtGJu+aF6LW+e42rMO4gOhyFhR/QIY
rVy4+4ZBNz4/khMRDyIQQiTLqqJJrgWSHhRl+ApQNIwYxnK/qfV0qYIWOjP4ByudESGxRQAEizaQ
u7o8UFjb+14Swgvd/megq21WNvTOsk7AecsZyQrJ73WrCwZFYn8MfOLjFjwe20CaPJC529ZqUpkp
iZd711lOaAhp0/axHnwE+G2DR7sASYQ/8BqwxAxmcBPWwQrmaLZ6+mrSE3Qb3YaKUzCg1HJUX/uW
YfmdoozPg0UmYa3Voz8xVCP/GQsuw35ono4qmIoYMphd935jJPbykaJSzR2YD/3zYjiN4ws5ZAUE
2YKHraEwNfBU7ugOx8MLo3FLqMyC+Kfxrt8LL9tchc8tBqbiRdUw2mYEHpIRTxHq/Ec2p5fpDPZk
b5EbdGJwZWKlrgQHsUIAIUGNXMqRyFjJRwWe1ann37TC+x6vs8LshsciGyUEoNdDQJ/nDbYmHSRW
RKICLefeK3XNp6mCH0uMTUL+kusmVeT6C4M7cFZ4rKn63zpcr6g0BXtA6tt+cG/D+MkfhbShp3Wt
4zsOfakpX/e/Rnoci+NqMLK0EotLxrT1cF2mjP5UTbGcKw1/bdKmmI1XcXiAaJ+mNuWuLzi62Mq+
DVWRxm54NXmz3ygx8EaOf6sV4zTHS3dQeIeBYg/PcBs1/lO6IEUjtC0H7JWdsxDQD6hRdFFvdANP
V0ZlrO20xoBKFU8F7Gw2STYaYfa6FaVu6W8BPUw7Mzc6dChl4VBoBN63tnlucr4qXeA5I1+vOJVc
PZLTIuTvx2fl1Lox8/F1gNxKeZ1vUFGTgTOBCWgEP5885W3TvNYLrBkMzXpYK3HRknSJMO7fAoXP
ddN1uKjuLzt9UA1mZGytOdn8f97m6y9/hn+a0JKnzxf2jS4yBQG5qsBMBnK2qlYoaLI/qLLmJxNf
ADXslIpLCLR8ELdW9rHxa1N58FSZIyiMf/IYoR0ChxNb/LX0PkHxCh9YeLLgE1IutnAImPAwR2yE
blbDfaytquvKRdrt9nebp8j7rQ2W6XDsPNegs/gg1z3CX/4t4c8slzIDWLz+f74QWFnDVZrR67Eq
9H3mGOi+onDDDTodV3VEWCRaSbqyks53l5vB9xhACvXcEbwlkYAI3xCStTf2qJiJFxhClzeBGhOS
iX7KabNOu8zjt9R39ZawNc3iUZTgoN7r4CI0z4omwX5NylWA0BEN12p5yvlsXMupoO7tAsfaGI1L
0H9BntHD8p2+6CjoPxdYtlD9G5lmFEA/MaFLs4vOvB07x4yGfGKjwvKJ/1ew1VG9HnpHmbZHrlZD
77WnL4ao8BJMzKAL4bvauWzyzjM9/trdppXZwxkhbKZupUJTl1abASMqrU9YFF1rhf3CjY6wSsEp
NkO8HRGjQWACzhMMdpi5VRcfWCNU+GhQxR2VB96svFSAWsU8CszgBXxdoI8p66Un5krVirBVEkOe
2YJEf7AvvZsWCoLcK3A/LuDhy8QVQQhb/ojZfRoIQOFolzZEbk+4n0vg9OlSCj/5CU7ihg6UNwZx
O58KVjVH6OeI6JpN++4qrldVJPWcEQdvHTQF4y7mG34hbeQ2xrz8MkhYMSPCOX29n4a2VvjLouR+
vlWer5JoJaHLUfKiYNzBIr7bLiTwJKkkPgktIfJxxeaHj34HQwJiRClgfewPlP5HKgirhG31JDkZ
X79Bqkato1NNe446FH2GoONKiTEy98i1YpEhhlIUR2V6CK47jZRXGnjazv6uZ3iBiPMx4DS6fIdq
4rzcKtxrXRuSs3/NoRa4bW+J0tagvX3QDL76A6gy/odueFlNaGfrKOJZTGmp/nZKsSYzhQkuKw2R
YQlpL3MHHQYc2Qtwv24vBgA822RY9LNC0dVmA7EUSox3B7ecIrTu0p/jyzRzL0wzaK9UMIbC334K
RGvhWB1HfOlB0jvb0WCzX5pbnL3HwFC6UI/Qap4MZSGj6DOjI1elyRrEmYgpwl+Ocq6SEJ3ASXkw
UWSJJx5g0WO5y+y7UpnIL3oAe79qXWZlSxF1CTAueSuHHvB4GRSWaKDSXEh0LE2+UGNWG9oWHGVJ
Zj2NM93PwmPl1KsSoaTdSCjDNlDNfITDy+N9Jf7POj0XQFvROXuXymMMDnsNugqV/Qki8/6Aa9Az
4YXNSIzBfMyHlogARQTUFq1/RuCFcmJppvUM/pVFMhCga2kfenleFo+noTz9PBNrL9k1XPPn1+3D
uD6LaIZgEu28qPilKY79VB21xX72TS1A7AJuLKGfjHBsiugITuIDx+VHKefFIY+1R9blsDh50FD5
APv8IZTmIlQbbYQhMiwZZkEx9lBv0WiwEldxhF7gdy6Fwe33BerFSAtCQOaZ+WA3PbkHPM6y425r
xfS03oF+EC3w8F1c6YFSaPX6xwUhYvzvjH3w6A1qmVYAZBS/Fn/y3CfBIaLY31rgCU2g+3aZ/KYD
/9KMJb3De+CyNHeCJq8tvSGo7a4OZtPZuk5u7HRr5RU117+XV+/vVe1gP4DS0JG4esefREhRnWvY
oLsH3iX+fZ+saSSqJlz/gzi/V5G0mFw9icRrvCc8yEHHXnPGo5eodUPlJhJQ1Lblt4qrfbx9JgOA
GlODuXgWTzIGBW71oYrINQzWsY1kvIqxECVncKGYnMmE4Y6pPTBTuXZoJqH8coeleo6UazqjjLlr
EMiR/IId86C3GDLC/o3mTTFWtdZJsgnJxPEfTPMKTYvBx9sbMcK9KWk9VMQascJ/uy6wgjXjNJfN
VzLCMTWEmkl4hkHYYp8ZUooy6IliazIZ1kkWL+HcmkhU0eHeoXgUXtQfJ7GyeV8qtzOpayebhEAS
PhS+ja6v/D9vuHHjODwtKWL//YJQxRL0sCOKT1xQVAFybBEj+m3JV1Jz+cjOE6ZhAfyFvQgdAT/2
RqAL6ZQI91PG/WNPVNAipmnsq97/4GldVYGYMawHRhnFY92A1MJzJkUv8RPNJsVlXuO7JPXYePB4
xrslKMhAhNiQjmeBfnHRrP3SUT00ISlltlwM0IPlez+blQvn/cxwUTf/zKnibgBLWmnwRCaoTWPv
kEFI59OL7ENHcZ7X489foKo4ClPx73BnDlvPXvtgiK/POfxETCW6mUaqFiCslKVNBAcyZn3PU1bQ
DYgIMDLvKz1lrCRi9jUUvWyTHVLk63XvcSk83jUXjm0ves3H34eY50yU3f/Zejzx1XL3Netry5ZO
k85ECQieJXo2qpvppNyFy6UvsX2ejvGI8YioMsJ/19VxGV3XQp/66JsYigQ/qiRaIR2+IR0hhfw5
We9/4xCMEfJeR/SPegGAJloUlqXvfIvbGK/lCr3I7frCv5Ut0jGTHjCB6fD4JG+m3aZfeAHONprs
Ew1GVD8Mp8MUObhrAEHAVHo7+IAWWwgRUBOII1zAe/cNHjU9bU3K5NYVb/Hqtowoai1weH2FbXeD
fX85uclZDKEg7YSHoO85jHOfiJopcVXyeE0Y2U2nbWMJdI/O72ZKgWenMGjto9EtfZ1Ll3Z7SAxR
2qnywHaa/gc9Y0ukmfNH8ybe5Wwzpi994Q1nOQeoTtfTwsIBkDvPIgMIG4o12449bBOhhOqj3XKZ
0072jYXzm877P4XA5vpOmiaZDJ7wDXhyB7NulyuX2lZHddpvX9mJ7t0HC22L7gthaI2cWs90dRLz
9RdUHQ+2voYtSbZLHVEJhomdGjTa+ciyPhOvAT+twdPXjRSYzAtjsfSGXy2eF9GZ8cBKVAE9k4yS
hi3NWGgc7sR5kRvtX1MRHVmjRnlWeklM/QFXazncp/CiN9G7yfRcHC8M/pucM/Pp4HNsf5Jsl499
/Vqodi+L6PMGLm0VW0bHAlLtxKiGqTDykZ/4mWkGNt53BIZ7YxJc/dpwBsvGz8orwi4m+2kO8eXp
1vPUi8FPUsEIIcA+TKOuKEM63eQuZqEj6uQzEj7X5SxXMtLEE5eS/wgeObfVsoX8HBTaQZq0lvQM
mR5cdYj6Yfv61+v5xkHErZ9qWAvt6UWx2Abmq/p9nNDL0oFMGytM22Zr8WpYmhllewipr+tnQzYZ
qQM5HoNRAMKTDfOBmCWF04FqxBXeE0t5ar3V+PQmCa9nOQEJCws6V3MS6A84S33qDGpBqJ8HdMTe
+WAQk8CNWN5d2J8zvuIipzqKcK48k4jryr70vp/8KuRqlELacZ1o/mdbEegyZqk1czexB1/HdHxM
IZ/bnSrU4+9tpx2IwHPfLrUYv44RzR6MQQ/SCWlmEWhgtdmrjcdhAOw6NapSvPgepNank7Fa25c9
tJN1mKA4RT+xyTA2om0uKAaW+w8f9+lphlnphuVDG4JWtuRRUnkZOLdkwvpp1X8XiiXuUNXGya8U
Q2VAhmc9ZuRiVmyq0evLBdcpCCxH54HgV2317xhv2pjXhX6/YpjwKWN9T/7sCdkPbPLWKy+uuQQw
S8UtxSVatEI4h/lsnaYrU+ojkh4NVLWQSyHqgGefj3kqXoYTk6Ysh3DFwJXPgSkohlYJv7mdRHPs
W8N2LoC0EQDDkTd1/txMdFZ/EZo5W4tiQAiaWFvCvlg5jtcrHRPRKN5I/vB6XtkI8RSuhCxVzYXO
Cs+mvm92Fc1pLMQDDRCTpsgL62sZa4XypA2708i2kmvk+U4ffx2nOyyJPVdcSXoVjfKUZ1+DRDw3
31Tzwsql2vmpPc1wEQbBpy+5lDLF9FCZiO5MrA8Vdw2K6PzX9i05GYHDw4ZLZXLVHTYWZqZP8vM8
TZBZ+zHgPwnVVPK2tudTrtgLDmdzqmO2u6BjWNeAAkS7Jbt26UV5FW/bZ8FlPgxLZ+VQWOzHaIR/
8cGHwM+UWsTrPFKkgT2zfrjHCZuVmGd/1j0lAlSqaucHab3Kc1j51kC5byH3qKxy/e+4PwFOLcTR
lcLFK5CYqhhytHwlGpAIz0NVWdlPpjdiSfKHYNYHViyp/13dqFfZ7Z384QAQcOPS8HvwrHZHFtfU
DS+3RzLo4sU9ixiBoSwz/AvF6pAGH5F1w3aCCcibOFluTb4zMJhH0IRFJ9riPn4qQKFjTuwxs776
nciluIVuZW/wBv4XaDWSgNz7AHQJhrWKBehR4THDKfW89cYkw96/VmsA8PjmTiKlQZw6xPexDBgX
QNzliVnOiJ29kkamUa8TwYpbJEp3uzaVtuoDxmsf2DoBoO+X9VJ5q8lULCC4JsxhczNUo5ByHWIr
id8Ts5wbOzSNrZH1zNpBCEgEnUtlfCSh79RLup2LtTo3kRhBLQuK7zMLfWsKaszv/lk140yncixQ
tKI8CBWiCDVEG3NZBSxsSln+GxceTqpXmQDYLQiLg2jS29yTtrtxou1mrOedpxm5qniDQxOVjgyW
x61i3VNgYUNsRIQ8XAlvo1kDbPhv0jZTglh5GgQpAruzXhKjhTBEdc9idsPwuC0d9m68Az3QW2nV
dLNVouqmppAECP8FteiNAMGmabo301jpdkJOW6rV4Mux9kfuAouui3Q6PH29agpMk8YX7O0LlSDj
MolTO8DRNCdr1omiamQE1/DjAfRhAnmIIkFnWkXofO+mlt/OBHIiENOU7iHzeFkJnTXAieAW7VCz
Y3v84LnKenwX3q3nkvfCthbQ+DODnsput6ShSBwoJUfrPGmayVIQo1w0Gf/+tGlWri10+N8H5ixJ
Cqs2ynqure54T1jr4MswVPShKSNAEYiUfpbK/NRWkDsXaMyNuqgJDMYmyQ0Rj6FQnDWwMYp7UoDK
kYxKpS+Mch1tMKWVTJz3pB+Sct4fs9NsOKNjNROg2NG1Um4sZBSSSvpdsmzlHEPncWwpMGJpZVE4
N93JbWoy+FUvQY3rBpXNbhveHr4LpRz6GTuA7cZ4MzYSmuH5dqB+SRv4CkVcMugwURjteNrqDUWd
pxsisCLVCv3OkOzt+kVeThVUtcIHLcwmCya7RrQagGekpWvwK9FnmmRn+NbTG/b/rzjee4fDq9i0
ignKuGZpcOnjF9Y9k2vI21kxcRXViCz+lLjzbIAkbYMS+9f6tq78juegBisSVv96boIVc53cw+E8
ZobVweA3Ou+Xit6uCgomj/kBDh95AdzW9M/nqvID2iiqIzIlhJvtgqLfEk9aeoqis5yiHI2U4Gvx
Dzo0KPFEcpMlkzCw8p7YC/yCFwy5DSJxGkzvUaN3XJHV0lwgyKkezvxPTiKym8BxYimTuQZB5eOE
48vFHbC3PxbhYtrTnNi7JEmeBY7KfLAas9m4rY0ws+Gfm2x1lpyJxALEsGqeUdjXa0fKrigrGiz2
pdUqMZGtMAmYWzDR1fI8A6rNzymGj2E6iTAFO8MVjiyAoaeoLxprvuiLElux5v8r72yQr/+L3h8Y
rBXKmhqwTQFdGZd2X2yKrbHkUKmb0SXeHtbMWliOY9GTTbdOUjr4vm3lzL1ZuKMA7ZVHOJfPi5yj
KyEOqeCxuCBTk85ey6Hz/+nBUlDRSqyKLPZZQMbAr3Wj7wbLBYYSJQfGOYMuNO+AvFuGIlt6grK/
YUrV+FZxNhUP8ePkPqPpn8mXkDZnaQTIQsCh9BJs2W0rYVmdgdsrH2o4EuRb9gpkCjUa9kUdHiQa
ynwsTmt9i1daiYT4cY1eflaL8h6AUg7dOprJkj/NTZwtt3gE6oxgLqanBV2XlqZ1es2AQxv0ojiI
Ziw0P+it/QExtXhfjeI+dOQwKTcxqJ/S3o4oguP4kGKoH+gZAsfyjrWESYZ6zD9jVJs0qAVxSbUB
+i7aHsfyUmLc3iOP68eDoaaDPrS3QHrOg5C6nyNQTB+eLQLM3CPlWxvgw7ujO3mGRN0NLqdBwKRw
O4oPb5G9e/C4LszP2RuS1Zi1/sgqXw/KkcnjkdryXQ35g7BP620sQxMSnO1cwyH0A7MkFgGOMb2W
eNqKajzscoLQbU2wmQ0slbOcwZPW/DjT35rgX2yUQYCJ1/qIE2fEU+D3cKa13nYLHrrpWvc9ecB6
o0izgyJZsOCmqtds82ZR8nDV6C23hSF6vnC0kTpWq5srqKnHVHxXtN1D9euV6rsAQsNY01m+QWEb
F3VUTu2ZF48sGUKIfw4BCFzCZFsbnFmbNKnaK6fg7sWniX3WTHnhoGZIs7JxelzbgqQ0PLmQJCZF
LYZk/8fV6ypanWHIbhRzh7+UKp5I++N7DZ1wgkg0Ogt6PuMa3qU/gnvImkoY6akWv/I+IWf2Piqt
RKmwhsz81LZPsAcs7qCFWsxgafz2iwORwiCRtVf1gu4nOGogWfcmO6oUmenc9glg7bqzdGGgGwvN
ehO/B+asmurF+Bn4qEE3gZYn5OkdSJ1ydQuTzKlgSIOS3TG1hajPF7bSJNDOz9JyA4u8TO8ymHQ8
XWHHrxW6Pw07TFWIH1fY6SDFg2YuR9foBICtU+GOg7Ps8v8HxfYKDFmfcg2tFBc4mYomCouocR5T
4Ylelgp0BWh4pZzAgHQznU3P9oXczZWJ/4mgJ/AuoulnW+ejx18Jz4tfAm78PhmMuzyQCY2YiXqG
zkjazdg/EVz+dIH2fuOM5ToXt/bECUJvE370X0MH/5qHoysEslHkTMtNzmp79PdMsqxMHpwYbRs+
Fu15MECPFFA8v+Z746+jxrteptxri7AVrfT9S9GMI5D5hKeVnVD+wTl9ivjKY22u6C48+qNei4o1
Plm230Vt1zzFNdetyeAU/NX0PXTfdSR6X16bpy1fsb6vRx75XXNjjLHPGcJHsd4CXLckGR8Fu5Uy
yHM25PCw74KmJ6HLnNPHrnsDpmL04zKEHtl+utNyDT0Ma7qbvxY5n1b2g1E9u1/AGGUiFh3Fo7/8
PuJhOxxQUEp+LLATA7cYu0SeV72EyH231F7t/JZ0LGL4O9AhdDhow2GZHBsyGmMAL3cBsuG6vDxs
kjWnTloabcdypg5XkgOdEaZVli2eEyApFORZUBE0tAWizlvHvGMz3cDfGuVuwRemkFlqif5RUcCD
E+7fBid6QK3wHkHA1NDnDOaVTBW+8sOjNsyf7AI8WqiKq/1ZaUj9A8yq7BDhuxXa4oYZ/Woxy4dC
rC3bODwx2ena98mElvS9CauGcb/Bnj+An/sYpEgVq5tZndHfTkEdecTBm2XArlp+A+oF1ipG8DS5
WngQhC42NDhE46PyXjQcIACKnXJCANaQTg3w0SLO+3JJpvOEQ/hHbSVs1P4l1CYwR+Dr7UneGH3D
f9uUzJbOuQo98a7Aw+ICEfdheEe3rBvNc43rTpBpd/n1BIt3oM4svioCKBSur6RkiuHH0KaMwMJN
kD476M0ZdYQvAZH+lCzXHsVDrOiwIZ2RnMF4XJ5puZaB0ungl/nX5LijofnCQ7N/++gND4gj3JOH
MaRbEfS35OgF/FYTALha1VwZ53MazGqAPJRtEd9fWzLovPFLuxBnb5H3kB9Za5/9yee7PgxXiMup
k3BztD2oOcZYLAh/mGaKvjwLB+wR6NLyaqIXdXpbdOozrQhdgAh+wPKKugcpVQknoO70e6XckHZ4
0HeLwGMmZuHyqkOoDAHaRbg6CCxL8VMWZPhimmCu8sU5bUG63g0/eC7R5ZygBk1g1Hv3xKf9CKiE
nAy9ZNz83XixkDm/zGgUFRcjSbCjupeCJ+lckgVfalycxGcxGGxCl5ifjjEFmmau5eThT14933cd
InxnjgPbLazCBeBTksPqpSB5VhXPRgiOtoq88WZ6I3I+avSbVsUvosLNQk0dYh8C05kkJcxBh0vM
bUS9/E+YVIG8tKUqyPjNfy9wH+WKK1KcyTH252OHuysYwE0x5Xq2ncvhVXL1MG289tb3HbB1lG2F
5vfCcArVWQwXqf3t8h7/om+mMnl/LITeBvs8lfdc5EjUudeNY9TOFNLcMcPOtijrITeHvqjRfgcC
s37sXb8/dvS6zr4ZqqVgQSDwPUhc0MphvcRKX4AqFaNA0326OOmiA5RCF4eTBQz35x7RzK8BKI1p
d/KM+3G3u6T8dpJ+hXP9PkZEDiv2zSBGtIHR9FT2Orc04T773D8G5G6Iph7AzRlp7S1+LQkNU0g4
io6YKmEFNqic7ZsMPIaEloyZOnXHdg0XJdQ1S7UsBfkUjCHtXTvF0ps7d1Rq2BUddEdm7t4vCett
XLSQRwBn9FyMndbXx8SSsmM54ts0F69/n5k3758GM+zGEIy7ZGqONupA/OigdLpU1xYWTFhKD58g
quXO029KskeO8yF3IrXmxRmr1u6iLJ+Ouuh6HyScDZIYTpi24C1D6ZxfxL8laDIPgudALagyKuys
f/CoDg0uBzIMTdEH3djERmBkDa2R16STcy4HeplogvvmgwftzZeA56czdftzXP9fWKwxXfJ+AeK0
YgWNjlrz2oBBSjMgnDmGuuMjJjfUA+I0dez8nvfw3WTpBgMrUURU7kzFQnuPLYh+kWIktFS0d48V
fsZzgMLn0JNu+w7jcuKbvkecCtXtB7lHXTzJvR84ELsn5Pli4a7QvS0YJVGQHPZIgrKAMna8vQkg
uv7xtFhTcgEtD0GyLT1GNaj3CpnDtc/KQ87AKGRGpG5MbWgN3YqsUws8Mqk8q+wJIaJwyFHWc6r1
wHd52Z5rKXEtT9aeSfvaoX19zTO/SZ8hcJjqzc4svxDf67FKEZ70OGctBGYf1T6QoxbQeX3R8rxW
PVKgNK5F62kTsex1vA5vtfh/r4+gqckTQx4lHaEpY/fpqQnnmrxqzh8kVFPG3PY/Xu8RWdwN4YCJ
WmN1DoCTGQQn97iILe1UfASTY3JdYWQIyOOl989YI7sE6fP+KMBwKXxp2UaGovac6h1aRlX8esVA
O5OxOVmz/jk9eF4j5SnBZDM5tqBoQA1ZE7oEn7mg0l48Q1Xkg4lElHJmyZEVIsuhofLM31gt9IRM
i38tzNNtQG+daAOyQ4l+iMq+v6ZpuMglj7x6Qf5l2/r3AS9pABZtmhGTnbX2+bzrwmEP1rXF13/k
0kVdd0+Vq4JPHgYENOGDq1P1Gwj5dTBb5Y8nV3KtAwyLCrIVxoProBtBI+QxSzkgGZ+OHNlrjgp6
g5gXjgOTmApMdGdmlsxwyIGfVtOCCsSvOyNe9A2Dnl2ZWTjLJy2IUp/kQCYFYRpz0lk3oTTR7iwD
DF/s/FK0V9Ca4pBfcMqgtNdkCjlnZPlxueYCUCP861eYJ2JwKMFciJZBcGeb+gBC++dx5liWszFy
KPsVG0FUqztTVClJ7qKlDFrH5rlSrRmePxkDC+ZcTNFNGXzrGhzpSgKc4N9G3NzBselEuVW2Z8wi
PtAt9LY1N6B6U63MCWZxLsWj6LcCs2mwmtCao3UI0GLxsZr8lf0qAQU6gtB5/xx7mUQgd5xDv7wm
XCXMfY53VKpTzyT6DFLwSlaxGmvc9jWBXnEmYW2IFWMkrdshzcunoldGVvyywdGVvu4lS/mVhAsv
vB+VUKR487wQf/ETV7Rtc36hVybt1U0dKcjI8LiiV5xjahLYaEEFH/BOx4QZ9bb+bAHQz1ymkjKP
jy8/3Ez5LLFnFBZiqPpcSH52c0gSIfBPQXSxqCj0g6TZQUQgIw0p8tVklw5MTt81AhZ5jFmuE7M/
pufqC40d8oqi0LQmefKzbddbc0ja5yZyCtHD/Eu5mNajcAENtwJe8HaDX7ltW7f6Uzp8C4L+kbSB
QFT6tYgZEzO64UoAip5+B850t+DJdwDCOajVfogSeZoVeRtCXloStLF0u28aJRDbPKPOD6asrqTI
b5vPqmjyMyCVrLZAvhPBe9h9ZDk5nc5TvS+3zT+HCW46ECtbhf/mchvKhP//UzJITdoQfVnKa+Do
0Eb5FA8gVurELRrDjckovDrcoM/wasejZulz+yEUhE3ZOdZXouNijXq/Z6ElKnfod6eX7JCGcDxX
fRXPcNLbvnP3WE7zhKC1pGI8VC2dnA2LZkbQjddnEQ0JSXafsfmiR794vBgfbaW0/ei0egYdBHc+
BnubEl/TG3cFnJteVnITK422aKkMnDqGj48gUi0JIRx8SnW3IMU8e//PALfSKU2PCGYJ/k1OrnBE
AGJ3oSyyqiD4zJDMJodAdx533IlSgxHve90OG8r+A7ilJpm3E4VLLPAL6u1BvHrKMqWSm9C0Cnrr
9aLSoQRxjrEWh1z2G5VK1+MDrN4xZkGwQpnGjU0sZmDl2N3tq6PQMWvNkUyLzu57G5gGPu+nObNn
PAKceJWmItlL+hdVp/KVenVYdcyv2DmqrKeLinMwbUc/QyKDF8t7LpZJ8ceOiTq5NBV7tt7H8g2f
9HJykTWpRSwt+/A3JiUEcO+vd4ZEoUtqAYtft3p5T0NJ6NQKeW/Xe/aAl85eK+Gp7FHHjFQdV3va
Mipti7J9ambUFPugdRiFOXiA2Nx/R6T7oRcAbaK2QmIPmEcDWJOQwiF9BZpUwKttVRe/UpO9r4/0
UdkY0B51LoaCTMZtmv1jw3v02p0SYd+aQFQfOkbi5eKSOiww7QEUrO9DvTbPQ+lrWwT73QBUKVnv
CvlyrID+Qt+rRNltaiHGEHiZYpjjv4mdGtQIBS3RT+ziaDnB1PyNdzQQPqJtNiIFCnsJ1y1t2dcL
Gpg5WGxVX2H6Zg5QEYB7iI9QveZwFVVNtLtoUtjIawxO/z6K1doUXxEmqSZzebj7UElfmvXGsXwW
pw2IOWJdvDKWGFpOZTvlFzX0390EBZK//HtwfYx9yKYwJaeRWwVx+1u6EdFK2VN2lavtmAJYVgIa
668NK+EJTxrzYEd15VbX532YIRaNOiKeDfvsMrbdxmuqlUC7oT9w6Hts+PpwEyJlrVdTUhGsfnQC
kkYsyYCRCRsAfyh8NuLH+z7hrrnewcmzSvHtIZ3lz1P5xTPo+aAxZi/03bZo87QVsftdvtFnGahc
G7L+bi/9TPZXGEExrETA2NyT0NKbEXpmD3NzV8SJs7Mkxsdi7MXnMSkThQpSNCi8+QarX8Hsrcih
nc3EE5wf3a1Dfe1YKvZKK63lyjk67VQfglJRmK/7UtSM/LpGmpsXoCl8AFgh/nCNBUyijcs0e+fX
IvIUJgfmNdATXjshrNgIfAnJCYKQV4MA5rqmCL8/ItsAAD9ARSfOIk0rWi/hSTSDohKOSTaO+ogb
DrtaB46+y0mJGY0qSpGy6vBmUzP1W+oBCKhXDJuG0s3Kpqcny4iwDIauTTW0AGM/VwnOjPkYQ6s6
/Yg42+OFd9t+dndZfOMaNVvGzyK0pX+2ku0Nh12/OxUaw37oAKA5FqwD7ZAXfwYf8bPid+aIidTA
67RRHGqQnxDgpGgT+oPqMNT7+PeyWCsVuJCzi7bY3IGU40wtlPEVo6/L9gTxrE4BNx57ElzUjcbt
xMFAvIUHT3c4ztzrfB+nfIVBAL7fRYwMOUGs1JJCQ7jo93JZoZzme7i1nNO0dRtZi6vnJgNmhMUC
Hs/YAmh1kNZP2lCu8SxosbecjGyEkbrrz0MsWHyqYEsZuUZrO/4McXfbwKP6KLNLeQB+UY+XqIGn
2BhFDUBaxU1lj6dmg5GlH5RD/Y9VyjfWJnpeLx/RMrVkRvhNfyCDBoTFMe+7dkmIMYWNRB9dSl6p
QQ6mr7vjLAJldrxaWTQ07fanNnc5aZk+em00g+vDXF97DuxTBXRleEcZQkogkwvJEsYDmj7xaK/s
O94myziwtPYsCkuwf/81zVWs0E37oqnUhgrE7RZucYjL9bunoL5a8HCapNFctFEmAeswjLdJe2R1
jybnYX3htVhNXJsXMlgqybg+HIJkvZp7FV5/2FXX+fzOx05DATPin9rfks5aAFgLzDzT5dh60SHy
Lx3coP/1Tol7TbxSeGpJxnZ8PLzHbzCTHxd1e67bmNWYiaiKPsjyPhb3A6gRxC+djL2JgXnoo6hN
RXhpmUHtGLivDzEuMFT/7ubYQFoRgQXLpwDOncXrBnGvEbqwrUtcgqQJcyaM4juKidjZio00878n
PJpDOnrS/jb/UnsApSLHgyPv/1Ckhq0wPUnpqi4Sl5bZriiAZgH7hmdVzLxofZ9YvfHuDPqIfyZJ
73YZVzR0uONwupXxFRWtVEtSgBCLnCU/63CzYe/b3z7sG5agxCq9wVkdYkjUdNjh2CCywkBpCShy
CmQRdaDCiQWyq2tPfMMf//lRZth3inMmEuNICK1GXkP3HNXRfhUc8HJmJKXZ/ZbNrGSYHMd1EVOL
OJ+YpG160ykSUpvrFTCUieLYgVfUCAjds5TBh7gJZY3B9NAX8ffi/MxuOpTrrdClCPrivduLRsaY
eqlq9nCng8CLz+WmQTI3Gak9eDuvFDzulYwEn1V3YalfBxB/k5V6KSYTO0aPUVYnaK7NS8U6NhR0
XOUzTAkFq9X9vExKK/Jn8FkM9ojY6qdJCZhZxn2HJ6hUGPr1zzuvECw3aUYeGGiCcuP6yIS/3FdO
0Up46Y/2iL4gV2dzrNn/T7qVzcTgqtoJ9BgA/yPIKKBf/i6Y2LGfN1V642D5I7xsJR4PsTlIjvZh
5+wOICAZpqMHEoNnRRJ9uHE01fCeLh4K6Xt65fEYHgqOEDAMNIm5zMzDGW89toII5PXOmRariCZ/
h2+P/SOt8woY0aE7Kui+YEYqi+Bu50egB8FZrmuDomo5CfTSvyXdJZiwiXPjY0m5FEpTyLUqP56H
gHrwCCFnLaNrkUnGc0Pir45+PP4OFHhrRebg2Wcv969bikXhb2jqoshWkQFmfznFCL1zroEoS+ze
/AJ5c/luUwONHlWRkYsI1lK9B4eRqZUu5PZH2JoEV3cVgwsXNcrjDcVtJjvUhOxmm2Bweb7OEzCr
oIZeTPFL/PMfXak3Hf8YvFMim20xK68VqC4I8pRHjXG7uk+GixO3pSmR43yf5mMCGXsIQxuuXIk4
6AUit5m18KnSOsIKwxvDghbOPpOJEhtg2f5Oje2OBZIrtmEBYCJD/zU4RtwZPy0MMjjqDyKnGTve
qZHYD0N2AyC1PlhWLyczSXLQlsrCKeCH5liC4CImPoe1qJbDWUjh0/CuBYLFi9y9YObAdM3fkr3x
R5zYZBezbVhnmJ4RbvQg9O4nXeEYzKWOQGSyGUHpvc1fpi1p+x7jjcQPKBX+3Iw60Q4sOUPh/EOG
hBoMqfyb274r7unNyTbS4NJ0pO1ISqejA8Qq8UuGDoFIOXq1pj8Zgxkr/S66MmQj/Pmdo3973vEz
M0dbI2+3f7MF6/NmeMOA+pRGz2nZ/Md7jf9ufpDQP/K1MT0PkzgM5HmrWubiGjNDCuicbVHO79bn
po95bN7HyH9mllgjtuycizhiBUnHtGPWRXdRkcyBh8LpSpP7o4V7kRVsAtKQQJ/2z0Cq8HMelRLG
dzRwXNeWPG6/F34t9KSrBI3AOCLHvIuia89rddHl/TxST1z4DzfMKmdU8pijTRH/DR5NhedgE/Q/
ualZB2T1/5EBEx9x1EnyyhV0cgS43z3hjWKUGk/gxsr6Zgw3MozkoB+D8vbY3tIqL7OXcwE3NK2S
erjXkKlYfq/4WDQ4kgGdb4tBOb6VihdqurYlXKoMz19PLna7T3sgtUakRr4YnV+OOXPQEURgDq0W
xCGEqMTOzC2nh3257/wPPq4hW/DqPuRH4mNkVPQ2eyAwursYxTnH33LgCm3OQq1H9PBg4W6F4+tV
WoF4w3skNZWixiypCqI+LwUX1h1IP9USz+2TamD0e2rfuOTsG+6oSeUo6A4muPEDgRvQI/ZafStG
OE7tNYo2zOsAXyQ5oQP3+GfF9H5lNhd6mz5Vwq7iMIJf2Tqqe59XSoNlp/8Ypv4U4TpCuhLPgwz9
P6FNjUDjhryXxMpylaUzbR6UAnU1WO5tFLno4lg1VeO0neJeFKpnv7CwgRFi4yG6I6dmu3FPRVJq
4lPPCPI5KnfCtf/fTEpNNQc8Oid5kbfJ9DPi0WVYTgB2B+z9QmmusX37QSalepmur6DGpq6jDdUZ
YGvW4KA7JVMnyLLXOk/Jo5nxajHLO/HY59oJU4BfH7qyedLHpOs5i8LS++hQ3oqVJOLh8SMijfNy
eU7Ple7vpSx/ALxd4dIHX+aq1QuoFMJpUK2R/DgbDj5TPih4v8jd2odTb6pPuD4oIucmsyTKBYmr
w01xS/r0OeJChFr+WEY/uj8xKyr5HU9f/Dfb7uPKpqhz0rOccMMMm9d0ZgqkdJhDd46GKex2GWFF
3BWuYNzVdcFTuTyDxIiChibYzyuUbiSBnXtLIpbKN/59RTyqZLfviYSQaLJcq3Jx8X9F5k2/T/G7
s73k3JVH6t4SHjYIrA8d2gHHDsb8SLE8qEGhrzB/NqNfhigaK6PhxmIOxSZaLrxABksGZdiD2jrs
LNFveokaGsEZS3dEx5EJOefmMxl5aE24+EpSiuyfumAgGYmchL8CvvqxHYlxxQ3Al6qNeUagJtnR
yz7qV+F2JOaW5a8XUVTociLhurgV02Y52304QsrXgQQs+l9NXBXryhRfiuDaKOn/emQUel7TXZq/
wCoGirkY8lXrsTa9ss/OS3P7IbcpPxZpOWD5S58821n6B/PL73VSAFXB7ntYySGh4rPKtsF48bXA
yRemiCieork5H746oHj0X8xjJyeTLH9tZIuDs870DBgBi2/XmKVqfG6dr1wEd1T8pP6fqF+fsr7P
VWg1nr0fCWXEeDUYWTV3OIjDdRs+43Bvr3TbivIfeGu9NVlLLeChAbkyDsaZxlWHJAQbgsO8WOhY
GkLBeuZUvD1guaUx32M7++T6bT7+Tl+zztg28Cx4yomgm/AirnWbqLCPsPhQwqW6KI296NMz3+oB
74d5/aaeJ1IL4dGQozuzRE1/jXLxq0RLzTEsb9+dhadtBKdAxp3asAFz32ByVb5vVVxu5gFsk+TN
Fo0T/blV4/QUQeTsKPhU7SlX2aAd/Vu/CidNTa4nTB6GDwE4Hvi8LBrRCHlWPiRUsGEvowfcNp5F
rhzG5x+5FKjpJfnVSiNur/a8YbdNDU6PfnvFVByz19GgR/d6RgnEqlJLZSlfGTRXN7SGVf0AhETJ
kcZf55zTxnoSqercAHjmbSEZaKhdzVRYAChu2X61BCaVFdDgmi40tsgKA1lDL1VvOOJDHD2dZz9z
Rakr1zVl0NGDR9lyKz4pdxe2VJbfWayFT5rHYy7EeGsUUQ9xVHBmFqyO9Q2N82g1qSDcaGxdEYAy
JLX9APK/ja6yP9ggOJAsIn2KtuNCffuFEHgCRkVVV8wfaVks0hrTlbp3PWX5bshsoqYvDtU0epXm
9mirZLuYrLuoXp8ECs2qCcMJbdop2Mnwk2MlYnV2H6/Q8JuRQSvJStclJUpmABDf2YC6fWv13MVL
8PnV6F0fXD70xgFdgCgJ9zXuo4G2AzsHtQBroEEVpHzeS1WPKOnZi0BWF3kl1bizJQpM9C1TYGVn
kUuGxwACaXm4TGHXZQ0PK9vqoGT6zaZxWWEpz941nO2l/BCUlXRDO/7qHPjxnHvJ4QapzUEi5G1L
vR5WHziSiisCeVZbobL6uRjk+7iU7KpXZ454pZ4q0eHffjh+n8w3yK5KdS3hW5MssM2Uzwjl12Qn
Nhf1t0PauYOKmPbqY8GyFE5Oix5jnNBRu95xxRE97kDLBS64MtUHnkIoF1X/AbxjvleczjhF9RPW
aSQ33rfEkTcbaMn5ASqNe5gvZqa+380ccrTwrmDC1uydkp6MauCIii3bO0xHyxY1RX6ePAMRZwV2
3edrFQKIiVVPqAI+nZMWw+qUi/Sg8KNg6Iyf4ohVxBSi+77Cgm+bNhdHIMrVb8wHz8dQvIn6UhB3
b4H/zP7mbAyPBMwG363YbI7ii+/iwqtW5UUBTw6kdUNWfiSV+dqkZsXkuDA1O89X/ey5bDBizGJN
978odI9lKhxU5mPQ4cBNJjah2jRtRmTCpDBeIC0gmbUGpJH6g9bg1583gQ6dkF4QhoDBGmQ3n0ss
VCqKBnMM2P6f4G3bqdvi4egymUhh6WPQV0vfOAU4eO/0HUzcKiavQc7mApcIzrW0dUKrVm2b9hM+
0nZ/px/5jPeFnyBrLaraKSpWvSGSoSeEDt+dTfCqvJ2S1uHwpW99lqKbYXXVrf4nCyfdyC31mUM7
FWqY3G8mkOYv/gvDn2y0e2vTZPEsRXmvQv4CWwTwUIPsQxe/J9NeGRtH1fQYAZpzCiKgr32EOBpI
2TRAKh9n1TOFUQ3IwmDUathCdyt3OHar/BUD5nP+hKRFgertKJPI8fI3dFSMSg61NyOhMeaF02j/
MkN6fDuVfFDunjXPxC2izKFmFwuWP7vrEBAMehTVlolIO00RyjOWW4ZPScW6q3C45WkX7ZJogldN
9cx2q/cJd5pRL/9cmRfYta/+jBxoGEjZQR5Em4NaQb7ZCviageW1OebnAGVEYR5dMwYHbV6F6mhk
ULGPMSeCQNeuG1kPtXjLFtAbK+YjzHK/EjZPJ89KId69z1CLKYUM2BCS4oXvwZrwB+/0rshIEoLg
ndh0EWoVbvpEjN5S5hJrJcFxWk7nry3wzXaHp9sXXB3tisjYX5FpGEB1XMBWO82tiqf9VVB+PSHP
1WwftNGrtjdERqJzKLP2nWw+JE10IiP6pbPNM6t0VnQWSFuWo5A2PI8IqgqL2N6gZIamlpvId8g6
CW3gXm4WFAQS+QWHKeUiAegM9ChzYkenhMcYh1n9GtQNfiNOJicK09qADRn9tPWsX3PbX1ertO99
r3TQEo1PVARBPPRLU1EoOKDiz0qqedW4JGtE47jwVMSaNaVEIqq90r1mI0ugi5hVHHZxIZw79rND
bc00FlQG+qEFnynRhrpBFsm3CncGmxeqzjZ1hBONxbSx8M3WjH8bdXceNaQCKByW6c+hMe8ACeDX
nY5zIJuYRl7o6EHWx4ReKboP35ntGsfIPq8sQvN6y+wQoXJMkHEm/X15nx21YAYLpLAVNC+G6Wnd
XGUXKhnCP8YiJ4fAFpKHaxI9B0uyUB+7rloNiIybJRf1RTcbUQtlioezqRHRKsEK6U+M095x9HUy
/RgUPYP46Mphjp93xXpuRVFa8EtrndhZo3L3ILCbmFDeZgGqfud+nbjjYWzPQWm2f1dksDaT0+9Z
TSVz0OZPX43kyyfSCY359ZiAJmSjkG+3k5KDEm+3zjghu9tsgb3KyBFhbKaog7rjoJMZstPKVDJt
5UE5N3ALLlzal7InA5oR5Za/7uA9JWUSH6fnfvr5UT8omlNdyqJBRRueS1HDCGANRpxWxMoFzXhj
ATH1c8itir4ifMdYN/W28guf4awR3l+znj8LRk0eRmV9Xo6nev8j2YJaYOLgEwTG6HQfzvzwA/ZD
X8oZatE/ToQHOpQ2ra+KBAN+5Xs4XXbdai0bee9ldSxreljm/6pcctHXQt/Z70kvSDfk0H0nji9Y
IeAAKMJrEelbNFUtvK0zUX88b0/9sJJ9whkyMNf2PkFzFcR9xfDYszZVgZpDNvCH7cMi3grOdsYQ
y8wX/omzg9BPTcHm57i58l9cBtDEwZxhHuLdQ8UlUYONL/WyzExlSHN2r9qfgn8J5CaIzLKgRmN+
5kA0rAg3wR+PXNXzPHOxXDL5tYJsWXjeNHyYmAjqOaNIlcj8bcgS+pNFiE/YueezwQNqxASkDi05
njIH310M9LQtx3tMvqLX1ZKeiImbhtaQ874McGppDvgtslLpZBOvBNXaDfAKsuM588TpMYCkJe8r
yg+tahdDEum22yfCo1f/pdKuPqelDV/8i1MaMMHZsLWNzMkWSzNQgXAUyCFh88ibWsTmILpnC4vo
edeRP8SYQSpJENAZ+E8M+P0iXMuqw828rwpoJLAjys+P2SBcVoaX5FXTFf1gKa5LJJ8hB1wXrOP5
Bi5g7OkxN2aKQYgfIOUUO/F1I3s6u8qp8+4S/W4E0+2VnvWToiiiIpEkkfhAA9yk/YvwvEDqHm5F
xNTwxNQ31poXWmP6x3ROAoGg+vEX28FHtpIT1zFNMJNHGAd0YPX7ZwV1FOgME5/ewFa6EOnHtyFM
ER6+Y1h7ID27urXmcowkjlq0rIjREBnj9z9ROzlNWowCDhr6jCTZJgMet1EZJHKAS6GFD7AG3Fj6
VyNnxzdOIxyC+y5skevoxYl9yXLxc20UY8ITg8MtR7xkXOkCMMJLOYkbNmp/yfNt2t8TRF8Hb42S
1O7fbjfhx9rZpY5jHOTd3IsCeoiZBuBgoFHaAGndbALu+lP+TcYV+enkurBBTCH5k65zaxAVM+iy
2MJnn7MTbpEaOXG27TmmgkRpyAveewlLOzIS/SCVx0jAWl0G0WqEVk2fEamaHgORfIy/wy0rFK2r
CRDyfgiXGhR5Fat6K5lNhC0bfKcrVIrHdAcmtUeoO7ape6WoCKkmj/hAUF0Oec4234KlvvoY4VKr
lAoalYjxLbu6IkJ1zDEgB0EmcpvcAVhoKlhTdBNkN4fG5TKChphYwImExadUOJd28Yfam/4cL5cn
keppl3pCQtqw7ImqwsnmOyh9/HuSdNfNebc7nq5y+1hjLKRbh2Pct2J0hgkxOyKFQ5HLyXktHyjY
hSvmq9lMJ4r5e6Nwv/akxXREuniBRB0uqPZ77GCMa4IZnPbjfnP3sV+fThFVCOtT52bzZ9Z37/65
O/l64nJgsiRN5jnI8CT9WxkUXKbuNRPpg75gr0rU16MwJ+GieqgQj1rr9k/SLulynuxOGJwlRIXK
TPHFSW/ePPCYDZLZdeLNcgR7tOeYV/jPciJUz6QaK+CRJbjLbeQYaPe6Q3j3Aa39HPJcYQj/DQ7I
+AcBOQX2x194hQAwK/mXR4KcBSL5f/FNGqEARKFzYZTtJLVNZd3Bo9hGV+dxuI8Mc7+W1V/VgRg4
6O7X/mmiNOg4YwYqnVmtp8EGI87uOAaAqdbBdCObtWq9WCl297keijcmiuUVheKogs2m7WoUjjkx
vdmwuNbgeGrRPW+3Umq/+Zp3HjLLLxAMb10YvduG4XU6F3WLKzxDtAkKBQryQmHvcRmeWT/vsJVq
nujQAL7nmpxYndFez9PHVOH7V2zBV3LjgU/6kpZERd8a8OPtGPwayNMI8pgiNzNds2S96gHS7e/Q
iCC6KTM2RkQV1mvIH+coAvugs0jlq/SSWIBzX23z0DmeVuZSXoOvkF/bZdxmlpW5+4bTV+hrk6HI
id4rKrK5D7S+m9vNkL3XdrMdfVzYYxwBQHhJgiN5PlHiu7TS+2AZyHi30TO+AHR1fejGT+nTE6sG
N5FcPTGyyKXWPoLKY4fkWjvuf+KfwDmtwzRLadZ6zDxCzJXSRW6IIw5uM3BzGhDm6Uf35GIyQdzR
cJsc+YbQ+kTe1X0yDXmvs1NOqgwtAfBRAFDtoOFJr9CKqWxadA7G3vvrAcjHEosA6SVPMOyHOeYI
UwXs0uLQ56p6ZX+q05rmbTGMNNY9NSqnWzhu0Rq23QQZvPDa+cOb/vbcvDL/SdcbOiyn7NQl4zl0
eR1ZT7SPrvA8Ti/kzhrWcUvnqp5T045CeiNK1ne1it/6qnmRZB1e7qfPx/giqT2sOKfZj0OsOePM
T3QCYCpY4oxMHOlf80fqdPxW5p8NP76OJALI1II6jrz6AqzSCYFga76PjgjnvraZNFInC5JhwU2v
Un2Cz1It3Fn3jk1kSCWys43zF3upnfsDWyMjtoGTksN7YfadvpwuftFDETrs/XSoq/HBVEUHl3EY
oXtC4Ir8L3lTPn59Dcf+F5aIKEb7eNB1/rVMzR0tUB4q5D4+g0aExikZLzGzaX3TIgEFXmoZM8Ln
HHdSZXMm2JoF3Cy8VWgafPpcsf9PQuwzdVLCMbtUoZShQ5uVGV2P+tQm2zcnDKXwvdhX80yFSZLH
tRjE2Q8iFXAKczmGnrSVGkaW7f0f71h+BokcI2v3D3xKa6RMk0uiW19RiMiFWxeD6+VzIiGIv/Y+
+C0tib1PbR7ls838ekQkmEX6o9WK1EiU8r8yaS9oT/WV+nZpfcjjLllsmJq3ynFg59k37BTLW7Qz
pLFf5GHX9DcS7zOa5ISf3QiS2FwQOKevfirQVEgPUFvCubaAPlveH9/nsOUacNFuS/bmd8gliS2S
2jHoIZO6CSGJK+WVNtu3SDrSbPoNnXfCkfztc4ERZg3i3RnyvLbv0enPWbntQBKdT9u6haR5RnGj
yEqRD4GloCEMMQf/5M8i3cCAwXjT+QCDblcS0anP2+7qY5ondTEg4maIL+OetG0UdE+Mc8mtD2wE
dxZkrgPcz4ALd4Kmh64e7PJb/a00IkNaSw03KGSd/o+rGslr4FoY3wRa2PE7ytKSFjmU487UlXg1
UwFdpr2Q27NpJg01n5WYk5zSdU0hSYDezhbqsUxvYVCh0y3+4gkk9rYjNLoDyvtw3ASE1Ol6U1ul
Y7YxcPfvRw67Xy8jxasscSGrS+Qi2lOX7H9b9JT/+yaDyZ8grMJgTFOIVIR96vVickC4hnmLNqEc
lf0AJ4oCihcnOZDNU0ddtjM7022qmFz6i9jA8hNJsV40Jg0zuW7SuYf8iPLv5RU8dKk8fwnuFrT0
VVAtNtakGiIeUSKuV6+H0K7I8CsEEd0Kur9XUwe4Y8FPk7Mdy3FbuTtILZnREJhaC1yQpN+jvWQg
Bj8gkEjZlWAbLdgTtN/I7MAOgLZA/75mqVf68Dd2uI9P556AxVVS/B6TGrkQb+DU+AOVnhMFKAny
u9gRfsZdmn4/LubRsQ4IyWMiHXr8jFf9byDZ/moI9EBkm38MMe6JqMYe+mWl+YOtNkqdjg3ikaDL
M3ltOwT64t8WcjNoAnBoBt/QP7lB8zIEC5NlAHdtDdghnFiMYJ1vdDApi/JUbXcHVQGso5Tsw0XF
8K+IYDXfiaKbHAElcxISk9eeZ+8m874xM9QhpKJ33cSUrWNuLQfhI5AoN4btBhDuLnRJ6hi7FNTF
/JPu4/yMWQL2bxP4Qhcm/pBSMJwF4Zd7vJv69w+vIEzQQURT89v/52rfjHG6XdUXL7z27wm9HaqI
6KP1bpqFXyOgWOneatoBtWwUcCBskpIgXF/iBo4NybY4TVGcDqLBS1yPP7Ud0RMyMwC3smOKc4Y1
Bkp9a2VDJwoWAm1XxH6hAh4wNsJNZnp3VBBCcQ/7laSO6MyULY8wj6slRQF5PUboq1Xv5Yx4/seq
EJA+6uNZm98zKsALdIpI6UamFmki/Q5+J90+BLRjzderBf25UNDMWJBRDOWOPsYViRs9FcZsr5Co
xwUNeZgVDiGTAmU+kINAZduiP1F2pq5DNiAzD4RxBDZwnk1P/O2OPSMKHhhQoQkckZwsIVgnYkB6
NjBtdLrogVzIIjSfyBbHwbw56GRqObkvqtpe5+SbE1Ec+hSCAzzFB88Td8OivBm8MAV3IoeOsDKq
3D1HJcUq3f7lto29QeRjQRapt67g4zvcmA7feU/Tq0lADx4D6ebpf/LAkBRmxxB8UOK27WHJbgpX
JsXXm1d516XkWc6v349J+189Vh6AuPCVia1IQIIWOqI/aQW7vR3bD+qf9XBFfzl01SshPZo/i28S
8b+199gMdYd4M5Y65XVXwviQWF4q9id4a/cdNgvi7osPjG4YwFm1iwEVP+IqNs+y5PcRSNXwPRy/
KO7/qg2NfAdM0xPSR2SBmUkm+HLSRb9S8OebD9h60KvZIDAyae1g7o2lXYmafwCRZZUwH2fuhtgk
+KK2Ve4Dp9eo99yLjMwgC0hgqO7qgC1Hw/4sgRvmRypplu36UBRdU2TBRMxocwAPKEv7kqhLskDO
P8ifOtBGsR2OzbsFBjWGqw032+B46Q429fhYP9vwltPexbkSd7WksBaHxBmUIVYv2NOryywlfReL
9goSvJQl7m7x0tzosIvOkWJfsEG7OXR1b6kf/kWyPyDT5EIEpfeM7KDyyFlqgG6cn3Pf6NH16PoK
c0H7pFTwsJ//Lity+zW7oUlWgbvB3XpDzcJ9k+t3FsYAllffY8Pc/ZIVFJzGLHnlV/KnoIQ70I1B
hJc0aHFRsfpWahVhYz0ArlHp/DNOKuJeua7p8MIIjxQvBPhKdUK2AoECsOOBrtiszUap697Oapr/
0FqPtOg7N/4cPZ6eKKBe4xdwFH4TNY2SM2T+1YRWFqAeuCighpWnVi1IGI506iejBr2Z5XpoQxr0
Dgbaja6ZPOO/WNKZ23odRx/thth8BO4tTe78o2JK//pUTNgmHDecuNxopqBLHzWn014dWWG1M/Vd
Xq+AB9V9p++GeKnxqwbfqb9g8VP8+sPAFu+75qV/m0ngBeBjncriBE+I/5TEhkeNaOM3Wt+JwIjx
Vlu6MBMVWF1zG2iVQczinp9Pnckca+c4sN0KEASSQEzcVYkSHIwMjT3y0U8TdyRmONoMBBZRlaj3
GEqFXlQJCJZZS9zp3BnmX3/7za6BnndtS+Fp/YkxAY7PeElYVrpaLbHhfJPkV8aTqWox7Cj9Y7zn
r1A85R/Y4Kv6DJX1jSULOPg4xxqSMuw4dVCx+m2pEo4PmqOPdrQQb8iBltHQil4ClclpGeLiew+y
sClnqU4Kfp7W9TkSMIsQ7oTcTfPfju3WpmgA7RNPRfO7+Vna0B2KBGz1+DVrDN5+JYcRps94zhaw
C48TB/fwQIYjKIL6RzCNNEHPIlJ6ZlvLg+V8BF3Zog0JtJUu1bb8kiMy8OBT1Yk32sIHQwLRwS6C
t8Nn3mGKWWP1YTGHv0Nvf4sIFJICLaEtAxi0po3sPe4QTr45lWLWb5ufkGy9CiE+QpBeF9sg0SI4
Pj4PWzvOQK1Nz+iXQyGcRyRl1AapR0OIZpDmqDBYRnfiLBAQDUVxzSgB+QMuywxoF9SG+6D73H0D
bASOrC1iJLBTYAnOGWyXDDJcqGAmT4WoMqPNGCyElu8FazYQRIbOfg5MP8pt42jmvgwOJZUgQt9u
yNF7gA+1to7mZc0wMyAv4oqWPrQBhzRZtddqmscC5zsZXx7UULhTsIKH0iEt5NlEHrHlR1FHgxbn
Hg9vdVgjqazRWretZdRE0WwNVgItVBGPOvr04Fn29dQPeSdf7+V3I0ZxnJzPrlOFaA5VB3waE+6G
IOzFBPomeE9YXs6Ky0qNvf1weIlGqN8XeeuM2DFqa2FGQ6Dr9S3TH9G/Lg84DXCoCBhzhXAIF3MS
fdUtefAD/lPpP6RejPBhPySyuybkqbWq68XrqLdJJG+rf6yFkUu02XYPEpeZ2TuelzQtZltC/qJk
AsIvZ43Ajuv5OuCSY7TtK8ZOMymKgaEm5zDCmCPESgGE2TkuPDbpnDbKKuUweOHAPlznDD5LoRp1
EEjqeEtFplrNB5HRIdijuMHb4/nhvON1reAEExfOfDLm0vxsyHC6IfItUlkzXSIuWLmm77CO+SE0
HGqIomruOgpLe4uZTMBo18HBq52+FSn25E3GB4t43yk4u2n0IWlUwgkNRo9RKSPP4nA8P2yQiyng
rhyHYUTr3QeLfsEE3EgeRz3ALZo7DGHfqGEo3OnI53esPQOgAD7nJggNnkOBXOsLwF2WFcItA2te
QcurzlJImgwIScytoll436lYVtcynJ6sKG97Kj/QY8Oi/23vir+j/PhKR5x5bN9Xn0mjNFdDd9g4
zlouPqCc1CXP2xyGnLTrASA9O14Z+lL7chYf9LIDMXOepz0RMnblZl1+O4vlA1oNAoy/lie+Z7v8
ytHaHkS+XZth/RthWeT5VoXOKusz3QQqMsjopc8f4K9OIPJxbCg9Z+cw077rUOWiklL6YO5cO8Nl
PQ5aP+Omo+DXqMANaXNjajtiz45eTtaggmDW2Ibn3/uQHuGYNVgrL1//cmNotnmYMHoKbI1Ps44q
vehSTIKAvy4FeaGA61kgGE0Y7unZwGYic0GJoG5Z6reKgVYz+QkjxUgsnTl93aqBtHJXjcsop709
VR9gi6Ma/8GC1ThenMnMOhScvoQrYnZVc/SAnHZf1CtS1UL3gcsTNGM2CSvY6ndGX5EzFvg8IpEC
5FyzCCP0xv7ukCUt36d6fOxm9PANoOSOH4YTpTEPxolgdd2eMsbmL7DyfgUdnLglJKrSO3km5qwE
gsnP1sIq7t5KCTG3LjGgnwZ01ea8sFdy8fWaEUgFLGZSp7j1PAy6iy8uvh6fYISKdn4CpSA79FEn
NC003XMcsAvsdBpji3tT/WhLZQ8tV3LPB3a01/TW061bN+CDPSTc58pjKFTJuqjM4hJHuuM9QAqV
DH4CrHLujYHyG+Jh0WEV4XqynT0BCdtf+0KObkLxgZCM9OwRfIMhKz2qHFn4umPiBqGVymXNb9QR
jUq6z1V4onzIrePzBObCrcayrEnRAy8HG66YpJyW2r0zle8W9Ykbt5O9p1QHm2enu5iugqDAxECd
UUy/wuDiqWi2TFj3W93/+NQQdFM6o6hoHKRA/Iaq/ZiKJu1sETT5hfjzHQn5Hrj7N2qq/bhZOc4Q
8NjhCnCKmTTlWTyhm+4jvQv/AyuBm6i0/XzIFO2LH7q7QLs5o7Th6S2niQcvrRvb1bWHJCg+y5I+
0xskAl0FgJgtHokMBq4WgIyMwt6WDpftVmAKCGcyT6PFWswxTpKufQ6xSILUfY5Asx0+Z2L3Nih+
ugXr3lo8iRsxFjsvRX7KQPYjDEw9Hi9rJKiq8I3Yw84ax2kBsipQIwr13ipYC7isChaSVKC0Mrdv
/iPrMjDBwl7gcG8gR5kyL8Wr0yvJt0+D1lR/rbEHA9MSbICCtK5w4q9AgmRK3kCKe2UIjhJkI7MR
+ahDKisxUS/eXDC8I93WLuVQKrTZr1pblFMOMZev0Or1EzlzJOZdQHslyBTiFyRUpo4J4LGDuvG4
nQg+pQkNqkg1bABxKwIAVpZCm9ISaCyf0pJj06rTAOOhlv+YKgVDRfUz4WbkbrbtXg4sD18EhFe6
flPZ/PWvUjG5bVQLO1E46kLmxmNY5/NjAyMUZRaIdSnYSNAEsKAIodhj1KE9eZqoxU8opXKU/G8z
Oy6izThbAum7ftsad2pE9GrNJVxPZzjLnDp8YGvTVJAlBR0d+OuvG2WzJDV8kAj7uWMVhwcPW9sU
GZ0oB41wG6+spt50VMimsw0cbZvI6tvh1hhQ4/v74vyHjhp5wYxB+p/YpQFuMDx7MZPFemCldX/4
3+BwTZAG8TA1UrCzco6KymF3oELL2Oyi3eWO3vmz6vzMKJJYprBVMqTfbVHEZOFF2ae/zgXDErpJ
gIHd8HKJ8MZhbLe8FODaTMrOQhpWmsAM7NCswy63yt/l2gsSnMFmZQOsQwUXRi0gMM8Kz/pLGO0i
UMCYLmVtkj+IXMSfaPJCo38n3zvlXFlf7jTeUufYr3c/QkG06/gn4qLB+msHX0tCW6aavUL+B9xs
vbQp8s5by+TzV9Z6rn4IxU11pA4no83AqGPA8wIsrETlqG58VX7qqUBIkF2dftqApoQuRw/k21k2
7nBpPtlcxz/9g1uqFTSdb1DeXSNWOJ/fLD9g7/95b+vC6hEdyC0UC2aHjunwyXgUE7NNhqGyIUhV
4c1P4Gy+ZmzyCOrHUZA6R/dgxOvRkCyiQepYhYmp0qgR7gxUkjv2tihcCWUz4NvcT3vsj/q8Mg6L
L24MZ3UJMTezVctCNMdiPMBApnrdLxOysdeXGDxrZim4rp0aKnXEvkWskCgexsA/skuXFD3W71/U
860a3TTez/lmKPmUGhHh5hn3NFuulAqG3YJYZMAir85Py7wmY8zMH0Eg02mjs750j5QpQbUciiy+
7WzTlLWhkBhoHVTpdRD7swFov3x7vjXcyEFzjtBdSs9jcKT4mTC0KQrlnDj6atLrm8i+X9EU4eIJ
YelEB2DsGzPbxNIy6+t7Kwg8IqVWV/AQiM9LJgwbuxBFeqjxSGijzObl4IEtFCPJfIxX9hP2CxBR
jRgrJ/bJZYBB9VYFFsEnpQks7hwMeTcASExd1yLxrZMy0aFMqJ1NHQDdjrL4bss4fpigiVh3szlZ
oZDXySW0TXD17cZgjyBBWlX5Cq4gilznOSAYy0wgwFzytRGG0Kb58eTXYJ17JrO5le0Xff8GCMZb
uK5yYmfDi4+09ugCHb6j1nscdg0wp8VLcVBYaceU8XwaFwQC3crHLgUhmoGqzUrJNi+dhRQcSDjg
Kr/vnHiSg3I66My2xh5I3ZZJ4J68Y62ptRmjqSZ9iow9fbNxb8lSEr/2uWjsEDD3Hl+RLFQ7jNtU
CyY57NcsXVbWtbuEn7KKuFoTVw08Ld8R7g7IwWaL3wKp/YtsvhBKY+LqMJ0GUTXbM2k+hvfWd/Oe
O5eN5dgSYMo/vPL4Cm7nVcTQZsuiyDb+lUYPBGx+DFdSD19dn80GD0MllX0EWL6Gm8XLIzvyEfZd
8aP1FdLhwru5j9vmgjk5wGQGM7l5/yEGq6ZbzWreSNlxRTvgwupYAp82T5eJlv0FRGJIR1xS2v5U
1CoSsdFElw7mdZlJplMYL1+VSiCsf2MEAHEXZ4FGMFSUgq9wuYWD6tEJbhz3jIk6F1o9hdCrABkX
UiI4ejzdKQIQ+Y7M81GX4gfXsRb1mBS8UIAaazCea9MlcfW+amdQXzJ183uXddPP/ZiUSabKsnGc
wUle6bwiGRHg1o8TySyqWR2lUEsR9sy347r7nyvAVISwl2GLRIlGwUf/sDUpK0Ym5MpQ5MmQMiHL
1Pd4bQ0217a4Rep07bp02u7aUZlBBhOynqXpf6Y8TmCSCBd3TudDPyumKTq/6OcneWlKIA3QML1Z
04/LnO4Okp+Y6fO+07GqTvlPgS8ZE+vDtahCnkRjWjsemkWEAxgQ7R0aWnSUhnUcdDQ9yozNatjg
XD0zBq8xmLlXyAjZxL/FfKj5zrNQcQbgP8PmKFUvkmcpYrKGfYQHqRxeHtylp/re42oPBAgNm59h
lSaeWCrp4GFewC0PX0YbEFXbqtZHH5wOqYoj4c8bj6f4v/dWNj8jXF/Tc51E8BXq8TigBH43qkUB
nOmTQHUCu5KqF0G1A2dpVzCPnc2VPRhM4nCsimN1YDO1B1Pm0Q7ZZS0QiN0LQyAj725nrzZbJGtn
szpkxNxojfQ66bw4jKtzbKkq1F3lLMQp/MTUag5kJLhhLpXS8DACo/NaO6kROwxWJV0NkPvPpz3P
1lAypCGI0ZgqrRJjZj+qXWD53mZDY8dHJgjcYPOrmgyCoHX9d2s9vy79uLYhXJDKLtK3EQFZSocc
KUL+xOyH8pCXOZJ3wjEmHi6uAAgE4Xs5J1D41zL1vzBvcwQ6Fv6bzn2QvIeXW+Cn+1m2ynRwEPoe
ZRD2WiRWd196kiuMnqhm98DWzluJoNjUTL3UVQvZeQ7//yZ9i8fLVInaClXwsEadbDkGcYGtO0Bv
xdxKoEJjX2Uf/SQfK+PyYPi3hHmAE6x6ZNdknZdz2zJdjCiFrcwgJuZ4BI4ZHx9ZOg/YJG/w//Il
gCmILYLr0cMl+VXGeqjJlkHiNRim4KgumzYpruuzR17ZSSJj/WgRsEXKS3kyEvYfGPybPhRtxn+V
e5duQbqjcyp9+my5cQRzEkrmF+NYBerxGbH4wtgdhM0Y/wl1ltJJYFWFeG8k5DfMije1F2dicwSX
t27Umw7skmmWIxKLQSZgpTmlNLxJ3cNx7XMlSz/PZEGDT1Rk8iQyjCoUfSADTx7I4HnPBwcoZK4Z
RKOPH57H0GcvEZ8kUlmCLk12XM4ugaaugzIPlk5Sip2R6DsnqJ9AUCbQxxBfmm4DyyS9TmK3N3zP
2tyFfQbabO5YcjymQpSUaI4Mbb4RDb4pRBSfmRULUyVx3Z0x3n9Lbh5j2+4ntwanucSYwiRKqrq4
WthmO2c5ftm5HijKSWIy8hUEDaiYnq5GMUswMn1qllrB0FZFkqelihkLklULXInI30n7N7/gQZTl
ZkNHAGgkYGd/SkULvUaVctzhmAnnYpL+P6ai2A+4UMdiCTwedHxih7G50LF0Jvd4lFFrAO/X+ze7
6049ffz+lq4rfphUkNvlPoLOQjukRUuaLaF/RfX9hWDmAXMWWDju3OBvppkztaPNYOhTe3Br4cf1
lzJHwugQYcP8QxHysfbAZfX9DIgUmwBNyKLet2GjRBjB0D6EQaeeNm+hNPl0FI90AHtUpPM1VhRW
6Rqvl13rzJH48Lbtim8nfCFHqkRHYMJdMHeA209bJtlqBd2/iyMBt567u1F1W6fPjQXTrYgqgbl+
atgfONy7HOpwc6t+0kPulMsv/a/sdCy6m5MV3Nn8HuSoObcpDZ3qd6zWn14m6nGu3p8v7oeqZ0wA
UT3D0hp6v+vVL2AOC4lgYHAN7NW8Mj9eUyW+Sm8oxaBnYGLjhVqF8LYAUFwHXqssCJrxHcTXdV/B
mf57VtywRpgrmylFZsFYdJbyLytii/a1fjV+YfGuis/1wRCAjfkF5UTsrF+77zHULSvTFapasHfl
TxUOVGlmUZS+oe5iQYJ2skIPjr14TFS0sQF17TyjeAgj5NhsbEcOkA1zXq7EQTE4bNI1ojmcnz/W
RpUriKTnYRT3IJKBHcT+W7tzOXm5Ks95bORh3e1Jnmkr3W10qSWWb7VokB/WRY9ICYoR9TTmsCQl
M7DCAADT2HYrjsLLfN8d8xDUVVH2XjV5AfjcQmj4brQav3pc4MvVfcuQNPo9+DY/l2YKSy9kMME/
mycBE4fUiPMD6qXK+P/afdrG8iOpOmfbi59sCmnZxxyhknoK/T76Id0rI6IwQOik2FNNAsLtQ2ch
pwzBO01lSAMXL+PSt+5XYKsD0cDyLdOEWvD5DbimZaj3v95tP0FUXm7DAEZrNegEO/XkAV4MQS7W
qLeSHEuk+LX1G0L15ksYiaUmhbZhBsrIHss2vVQTGUSvsWUruks4rXruv5lq1WjcsqjoxJiGG+Q3
TKKAGY0yTAWaTb5/B3Jqiu9WwXgF+zsAmaoRnTmJCDQ5IibhSkgYvJPUIQlU5z7uhalO3A/rj5DT
wz6o4R0UeU5yfhO7UlOjUg2QH1ym3tWTL2ZfV1v6DuSNJavjVEBbSXOH3WRLOJc7QApCxmNYi8uV
Hblk3kqJIho2jwxQSyX+QwUGZNzUSre4r0VEc+EMiTJI/yahGHrXLlNemGoA1T0/tK9IKJdTsE6s
2Ic0Ozzh6hlS/QhbVL4BZ8YtTUKuL2Xe8brQDwl/I3UOg6S5KvagJ52SY75KHgT9cSXUAePQXHPu
gRLjTZvdCxqEVWg1f9ALzljjeLfB0gOWCvJcKrLJ0HzBzRX6XkEpjgE7/fiEQ86ROIpW+yatk3KD
pTNfVWkOghvMdsna9KgZprNlUoQ9bqg9O84FtBdIUDNvS5pExEew2COLHuwGDZGQHzEipKhuA/DK
zE91Ig5BrKPYG9MyHDhQ+9JacwBw2RzuKiqtLP55gmxvrb2kXgj3TvANOi9xU8rDP+Ixbo40g4kR
BRlA20D81zZ7HW58dHZ/hsJrHWOpf/INcsbNJEw+2aWFK8atfmvjhYmtmew6zJrURuXAX3cEiMEx
MCh+I5bOUMIYSwmEyFaanCpBbIettfy7EoH2MuQCQVVkoema7TiKHsmQxd1qsj6U6eZS5i4FN1FI
fvFef2nCUjW2fEeoYw73842tAf3bZV8+4BaLHlEN39tjD+dE5IGeYyZHzVx4hCtO1tDNH/pC8NGr
6b02ILamhSTVyP+hoNxQQwq7Ma8US2hufbTEVEbvzFXnjE0JoPVGDzI2VSudEfKAwgQQEX1bdvdH
qvf+RJQiLCLIuoDTuILUZv3NFg+XGP8X64lL9VbK9eFy994HlM/Z7DkUrMIqnnwg7zk30rM89xbr
nXjbF2n5R9c3hB0s6jPJbosZlEsgFtmhWSOwDEOMgLCYyqzMGRSg7/jG2f6cW870493dIPUlOpSo
GvfkQ9AFfoEHTgnDZibWd6gtmvKrbNdwyr2ADe9pU1bOXfhQmyjC3DsPUowdRPDsmqLccB7kphlq
/R9lNo2dttMWlvampeCYk/lYSkB4gEpdf7cEiA6rlnNf+gPSk3IKyojgaMhJCRTroTh4COMCSEgY
BsGmu0p2BK0rDpN00Dt0r+98ZLRcqBJJVBDukbJvg7/ai7ENiedRHoEmAe8u3tIZr3zRbdIOj/2l
9i83S86650bfuEYoKyxkaLnKLFRYYUwHa1bpieLy9iUD575ei+x81Whp3CVkkar3ni3bDsvBQvor
Nc1cDOJe0Ysc2m6Dm9RA7bF1VFoMk8d7Sm4tTctC737up99KuLqvT7U9m/WpZtyKfURX0JNOItfb
Lft7EpWiaeEXKPr6F9X5kWGQKz3l4NAeCcjixDJ2+Q2evHLdCEQ3oszpmZW9yQ5FldFpAmxQ4ExH
82r5ngAcL9Ev255wtT6LnzCeBygo3h7yUx0/calG3p1RzqVygOPamjrnEquE7tfdxUDNHkS2CbY+
yjBRRyfS6L0U1C+SeAMeDdqEOzP6uxiSr0NPUzXhyE6I+m/iKKvUd8mt1uQ4BKTe41z59urEjoVd
U51gsLOW+vmNqPb0Dd/LOyYLheBi31hUO9gLyRJNq10oy3sZ00OfWOtWoXHx6cdGJtra367/bl3T
rTIh3ResLh7AeshgYq8JPx5bhLt3CnfmFoGJ+vSP26qhpIFCqrIAzu07AZKfQWLEnRlIdAr3mUr+
34KmsncaY3WYu3ZZVpfFg7s6JHR0plKF+y/302zBHaJ3gzzfAF6IdRXxtr08z/U0MmRkgbHlKTGA
nMY3d8qNOBksUu5+3FWeKz0Nv6qpkgWsWFejYwhQz7kbNkhBjaKp6AVQMl2EjQcSG1/siosjhQRA
zzbKR7b4msPIOduTPFeQNYSK5zF7HWEyvI0W+xNL9mumXDL6QKGnGSLaGEmNcVpUMeDvHQXIVNd7
+qrmKDqIPFEzkOWURxz6qDcryqYd9Iu36j7jwa15ehd4t28eLhMIk5RSfCJDMxnwnfzbrmuh5dG2
nJOL3A+QtrR/uNI3u5Y30Ff/FcG4niqkZf+STMSZ5/rL7I3TxJ2ndhQLv6yg/Qmdbg9if6FZ7S9C
Bh/z3Cyf+SaUlQAQa66II2HmUq8P61iVyAiUGqyi1SRo1V+UnhTU75RI3yCmoZGad1g7jW/ZKinB
talTMpyiRJgb4EUIUfPMjb7A+0FjMXKQVUefiqLdXQcWxTGfNedhHYANwS3XotUO8V1Ckfq7rzHg
sJ7ReJlnurv8TXjpvuPUjafQfYrIGvjoSxXwccCw836unafceMmhtfmxani05nAu4vF2JP6XgPSw
klxz60hJI16YiUaiOeBDsZWrMRUEk/Z/fewPmNv1SnI0O+MWpqiRNOAdjbrf5xLWeWSlZmkMWogG
a2AglMVC65nKUQCBTDIIS2GOcvISx/bMIiCrIQ/JKrD4YzES3bEYYNwgkUAGZwblUVmAiJxXVf5x
jNbMtebuN/Iyk2t+F2IT71JhvzmIDtH/Je8h7uktIFkiWrJQUf6+3ZLKKod5dkxuQTumBKdwS+U/
jlVvF08I6flzPuyEL6hIqWv4kEODiHMneEc12bVK7lkkyD+0z+leVKgz+vwcgIbLlNG0VS8IOsGT
QpqzQc4PSbkmOZUybjC9OtSRS7eHTVBFNS7ftTZzUOMxe58f68Ia4nIVi0CFBc1eS3r3zDmPh6yc
4nRb12J/VD/fVrhtfQs8z/RKYgxyfgNqVhL5RJmflo/xkcmdePEeBzsbvBnfPJe9J67E8x0O59pl
8cbHwV2Ozx0sMg12K71S8xZ7LvKYkohMCJbaHCGl85bbhapn/DeUNLnna3rKPOQE5Iz/hbgt4075
SVvAk3iFKks6pRdfnoFV1FBcJgjLyBopvevpeaJ0pdzp4gHEJb/ZV9f5PxyEfm0Kmavxham2WdiD
n32jrztywJo7OyWm6lRZ8TSJRi3BTzE39a760G3aFv53o/a5Fid/TPDYoXkji32NF2Vt60sPRVNY
feMhIMzaPWOGdpMyQKt41N1j5cQ04CxV8YW6cveGHgC/eT7BS65Vk588jaUt7L+r8gVZZ4GGEqnI
Zx56j7DidgTwQCdm2DpuHZOun4WdHdqKDta9aBkr7RI4rxsJ9ybQBMPEaYGzn5a4aeOqGIl8vRZp
KGsU8e8cEWRkGy8cuXkeWT+TxHZ95cv7UyUl7S7lq7INcVr/vLVjkvrxVHvkHylLey9enBTxY5KX
CGunlhX31x6yEyRm6dASmrLm8K4X+1DxcIolZoSbYgk1+Vyw5vbIi56WxIVkkjQgKzAs3TAal/F7
SkEFGhmukJKyjcTNwDn81nh4ioHJXbTgUUFkA20TxUnuPlbZdPyE6wImCf9xqi+VU/rh6BG0ASFo
UFEF2IrMyub3k3Wkxc/JZcJmb/cGfJKEOcMPXd15rXxvMwxq3RNZ+hVvA+XAe4ADs2iVAmNgNY53
KX7i9YfhtcG1wW3RRgE6ZX0QF/knl1Bg573qQe3HQp3KEjRK3IDfyIWCI5TWQBdMH285GJuqaWoK
8RQfCZHhKwUlXvA1jqa3piT+6K6ENtX7z/XPqoWKwIOOLcWBsd9trB3u4TTGGQX0pNaiqkVBPpuL
YrdpkDkXh5U3wPmYK1y7ARm8epIR+APRSSsfVM3oyZ/9saQdTWGqp8zDgSnKkikTZx6/ZSPOI7hq
iWYY0SXjEd6EaM8eudoJx+KvPJUgdIWuxdjJMlaVtSeOIDPdggON12ZlxBhwaIpvmUJpLapdNqms
Lgv7AHD4YNWkzJjafU6J7MPwvL42Topi9BG89VPSs6T3iLXZLUK8S9eDMJ1t5kkoaF0uzDXawfsR
/7o2xdbB6diVqISxOAZn9g3z/s6hf2Yvi5HIH+4eRw77nc2tHdHnZzLKKupGamHaRBv6o0a1wLWp
7Sq0IwyvxZ9MUxQq2zp10Msf6uS2BC0fPMJX71eRj/3Cqil/ai5dTpuTId2Rh4sDxr8JWTkvAJj0
2X97GaVIX8r7qVUZium/aXX8vCCgfozIGDH/R4s2J2uhGC7BOOmVsqPx7gc7bKYnWPosHG3lkOZO
8B+2TUd3wHlrP8kX1XALQl9UBmA10iP+Pf/Isez7dW4u3doE3Kvnuw0CGvSKdHP3zRjXlVjy0yYz
+nxk3lVkaE1x4dOvrJu/vVQs8u8tNAfasQevLhFT+ynFqK13QHZJU5GVTSGNE3O/Umo/i7/nG1xC
y9b3dwcfKaqZ0+Kx4eUzn1XpNK3ntxUrly9rCGWeRM/OmdmravhBHqvyrnGo1CoHKDDjne9lK9VD
0ewuETdCW4DcASDsM1JuXhHJBYEDhO51Rn4NTpmpNCJgapx4gMV/yk2Qxbjeh6nES/c5s0HNNGlZ
1QRtmV+qvsJUJ2Oy1ajlZCEZIqckFJYJL0jztAGXezPn2SziArzxjkodLJR0GFWyOqMS8ssD0R0C
Uj3T9UPxjvpDpIWcPx1oNpM5EJSrlG7slcClSBpHMcoZpmyhaxzTIRbr8bilz+R0Vm2PyGUq+zsM
72D6nUGlYBvgQujMdivxzYH0nU8qKnMpV6FG8j0ZDAAs9T4+ZPDqxlY+sYQYrXDKbV+pbdVrcDue
SjISAk+pBMxhChCF4KYx6sZjE3Ii3BSApkbymV1PvcQ6k3n5pSjXHnjR1dZ3EqROMKA5O9/QE7v9
FVJNriYQAUjS3NsxRO7P8SPc/I9qiAqx04RGZAE2V2x40PofoRalag28iCEVmf+9GRkRGeewEYAa
FieZg/XmamRet5LU8m2gtjMr6+PtNYz4BmxkPO/vitQ/kLbxIiDTOy+5a+RJK5zuau4z3MwC5rPs
i6m5XkPIWXq4QQ2XoTA8Yrps7HBZuBB9Ifllgg09Ir3FcvweKNuIoRomEzVqc3JSLxucknG0/eFx
zPy5vzLbehFCRMetf1XfJkrtiYkvIe8akFBsSA+De5GCXrlDIifw7uXTgU8cvKI2VK4M0hau9pNx
1xuDf3tD0KREX5Cr+/GxX+nL8vEXMwlDLQSDnrtZvk+/BWMwdbfCCk1zu1Yp0RBG1STdif9xxOGg
z2bHtpOF8yjuGdOS7k5faOyW/7bCzESN78hjC7YI1ndGUEdQLIqUmJUVE5ODDWKkblQjZRiAiIfX
mQzNQyTqRhd/zv5br/Bh/i0lhfjKxj5rYTyJ9Z8g6deD2olWVWIWDjiFeZiHtwyuzOmYFfTPMdOb
Um7s1xA4kAISzdIEj54Vx6hT+YmL5XhDzTiZceUJpKqE5WCjveQBfehDuVAuhGpgyK4/+4Jydt7V
GZutKfSEasERPmURKDIWuFG1bermmdQsbqOPL9H7RGlJYpbKW81tvzbZARY7VaZCkR9JVOANWCcF
UFimWEkcomMEi2QmdB4Kuy88MVO7GWoCkiKUWmXBH8PRlgXckyIdv7AK6kOyoWQbhlLv7MrAZYY7
mUU3J5613dC8Ve73O6F19kyDlwzJlWr2ZiBbd1NvyTKZS4zJeG+wqG0jm7I/PgP7jCpTBbHtTJf1
jO+Jb75aXRCbRkNq7p8E0/9MtemlLlKzKI9DpBnRCyLcrBDWewEaDVRkPZ0Cb91/AM7TaTfcODwC
iISA90xsjWfA8YOCOdO6ZIfAxR1wCgqw9eUpShA9j9XO4ISpRMWfaxzlfzZeUSW8I+hLLSa4scJs
PDOQcySFpQVKxj4+UsJsBUFFhsiMRjF+/DPqrmtY9BjJX/uD2pXHoHFZyuQ1INrFvXGJMwgXXtLw
HFzJjS5NwevLbWWc8yxkJHgNWwuhn/GUMgGqhVuIC1KK/AQztN90cA83O9rzlOJlq7zLSf/egalc
ZVCQtdQChKhT7AFudEWYi3wHE/HpZFsRXviXragqKpopeaDlkuJjn8VnIXgWngEZzgypSRBliHUl
ihufxCfhX8M5Z01cwpY/sce/7GOoSyQGEPGIlKjy7sEsRM2AsVUIC4X9lby5vi7bB81TldWRyzo9
6Rgw/ost3BmE1nvd+ovEkpZFa+uD9pf7FoAEKXr9Ih1+nDX/tF/zBNfNzUAZ5OAn9G1LS8yMLywL
7euIagyKqCR5E681m6c1WzCFyf0awGK49mH7HNY280AJqPnRPFYRp3o16ZytPdfGCZbmSRA1Vp5/
ATtnc5yi2sqCSupKA74UcjUtMSW9ijXNv7QjfRQVo/ef+RJBfvSqiY1rW4kPOJeeeluLI4P+pYt9
JnR2BlnTLcz+8Sgt3hZl06OcEgNfLSP5Zla1WUKg16uSyx+URAprHTxRujrj9w8LwJlbxglbtRSC
OmWBQXIJy+SmsP32elhhy7K7KcFHxlYR7176AHd8hIuZR96gJNdsgSugJwQky65/ooWmTU02ADJp
kgrCeftCIrOdNMHpBjLytJCWTdTEb2c1TD6+APTf4r8VCgOo4lPQ3d7KdqyBvQumRzxhqtskBqHs
D3QyXNYFAdl6EtDdun/SXD8m+FweFhgYkqee3142lErcb/cyAKFhRGXYxzTDBf2bqUFhMLpkx4ei
dHczX3Reb4DhxfDu6/3SAJNWsKgJn/AvUqiRwTFtJLSG9i+N67+Z7sHPUbvf+zOY1G+7yFXf1cUT
12ofDo687tu6wKVaS4XGo8UEAtgbUPJW4CneAelHr2mmIahqelCIDf5IjpVoxRrq9B4g4zW3ITo+
yqgeKuPMJq/cTMCIGNwyuW6JIkcznAQ/aomBfXPV4CN7bvp1o6CFkJfAq1q2HPBqAgDoeMrg6Vmk
KDalPqC0LGrKIpWjD00qRfoviFtedTUVgCx4EOsVCdzrSc49QPA/6daEqt/SwucZHUfnscWpzXSk
uMtTXXUjhopOBn8IBieM5Enuy98pmKGBXQ4gTUD0CMZ7kfqy6eN2nL7q9PL20AzUePkp/N/FRnC8
HnQFz3RrsTgfXMsyhGtSoNHwciDL4W2AWTwAZwMMgwSd1jz4T4+C1lF9VdXANZBloh2hKX9A4Fjt
4DG3fe/sROeY1YTXpMa5XysZm4EES52CDFqWovZvtm3GmyZnMNE63EbOyhdJxsaNgEV8MTkng4fu
fH+x5iJZ+VxxQD5kZnPpA87aCWFA6LfGBqLQBIPGi3h2xdZbePCHyNWJ9SI7hkVz+NbivvZFyYJJ
iHZCJMqUVOde0tNxSqPEQhhL/+l1O1AgUUl1t4Qfq713gYCGak93mYWIEYDMXiEC6eZ0Y906oCVR
c1LKOV8FkDLol8DZcinYunDjtimnVZ8SukFxhqo40q9GzXJyIPDs/LHEg4pCyEqtmZPB6DNrM6l8
RjZmurJPVllmK8WVBd3DtoG80gDWl8xXWX7MxYyH2m42l++njAKAaRGNNT0JMT+Vi/0zTI9xT6ZZ
qg3Q1kURe0wRdc6n5RTHH12LPAIsb+6D6Kg+4P/+QzsrwfP7+ChFIkeAYdULexCa2zF36kymuEgQ
pfMi254jrZEerj8m/f9KUjz2o7wzY4ObWvW9KfUZrABvG3IGosdXMWHuEKRo9f8VYh6Za62Im1Kb
xH2G5lPoMmVuiurtsVWHTr6mpzpFDHTiQ4vwdSTMuq53yvHJSPNTxWfDVXsTeJJL9FS/wAauBkNa
DEIfbt+89HH4ZM395yIW4eT827rq8mtg/izVmgdMz02jNB6NbNSuDSFZs7Xxw74dVBwwzhxf7CKO
Mqs3rntj1E5iAeNVcuIHBjI6OoEfTxpjrhQT8omsJ9v/srQ/o2R9Zt0oHJGqmVrwWbBmtCG2WadF
07QpMtdTWRDeVLt3G5r0572deZANSYuyiALg2EArxciRUlspxiPWdrPSbYXXyERiK0V67jOJnble
SECq3pSWP71xxEn43chkz6crrFu9Mgc/B8dFibyJcnnUzyKkHavs3EehAGR81oeODDjQVb/pm2zY
6umDnrjxNaQ/ro7EHIh6QCOhfDLGVK4cpT92k6yAH2gMDgDmhggGjKBdFHkG0MiZzFW30vTz3vz0
1vGuoTvrmoIa469oPSCxhYdRGYLGI7sq2IQOPqJ1UvtHs5S1/QYzgG5z1FUgKzYNQx5k7jHbSC9D
7zZKti1jGV74LWzlFs9sInAMW7i4gPhnJ1AFW5NKwjOHPeOYh+feEM/ZHxYzxoh/oF5gMx0dlXtF
OnCHpYobzYsfbDu8HADGUtUy5iS/jCuUwX9lRen3ZQpdJV1wMM2l9WgQsHjlp1ASCoEYF8kBR1Sx
Bi3981Ohg9RW5koMvW+jt3/34MBSxwxL/Gb99ckw5MRBVAWAnPQv0ZdvevSf0YEhQL5VntPeGLzc
bvSp8qOv8UYexwqTczkFkH7G+HaaetYWDHMwP2ZT/fMvmZFg4Ntjj4kL7bOdnzi0byCYG0D9hfn8
hktt9DcsDd1iSq34gqLeDyaQyW1NG30U8Eia/A/304gewfNg4ZUSKdvz76M6nwsg/E3dqjayEhy8
h7bluHAFI1Y1quN8U30wAsfi8qPrpv7GHcdJQpEAgslIgX5uEnHPFZV7ipEpmAuC4bAVKdf0OEow
VcC7UaE3GMdxA8dX6AbRd8VWjOfpm0gdTJ4OKeVnE1PmzeCm2FELKb3mE089Xj3QR8CRaS9ROfsF
oseLnGr0aKDUUr2612BTahq2cO1hhyxUSKqFELqGSQ+sEUUNjokbmXJWCvcO5toQAUGQQMbm7byS
AgUcG6p6uP9AAf8LRVjsDQHlXv44ud/4Kw7cLF/4DwfckZip5N3mWB/G2y2+La8/x2t6lGHPjftW
w2X/CP2tL1/Nwbe1x+C9hMgjPCg8ofkVU5RCvnqchvbziOTdg6OVj0EaTlEo+myLMF3f3/hJ3pU8
3/4d1Hp9/emnJPsxCmJcTgx8mRcCQkCC2Rjgq49qDv1k+AMj0SKLoctWyh1CphWRsJ+CqJo4IZId
MvwVrLmLsowGnwtZcqNoX5uYlSRW1PSK8sUC5iMH/rgiNwoFct8s8gs3hBTBQtBbHx3k5nqMbTpy
jbuddoeklNXR1DL4AmD5YX46EGYq83NNmQMC1ppVVWCVa05E5lpTjhxQcqgr3U1JUrfPLkfbXjd1
zPjasLCdHfBZIVBYdlnYCm0BqjCDxe7IzDDy9iuh7P57LQwDb/FSQxPayf0dpD8lxjCQyffCc1k5
1L9CZB0e2PSxm5Jvwoqh425vic+ePXuZZ3YHEby4NhFqOt/pfU6fuyGgxwR2sHnmhK/32CiTZSIA
I48KoA1kKq0AmZWDh6mtPc85SKmTVUtAG5xkP9KeTEEEqsQ7XuaMXwDD1SFVRWKEIJyA5MmcFtlv
StuwjOubiZdDmG0G7DwQKWpnSKJqREWky4LAnoGMe1twAbs73bOF4pbTCGYJjE1VgnNNsXSBZ6m0
ZdlqfxYlOWMTnBU7Dm2MeRMQ5Y+q/QvjkHuvD3tMCqCvhNFqJA2M3iEo49uwO/tDt71EUxWE/M4K
qWkRYeI7z3YsGxS+rfwWIBvEAVjqm5UhT/ft8S77MTE3I5JDT6rKy8u8zhJOxnFjUYHPB/LGP6TO
MXkA9zkyHY9tLzQ6FZJWkn0GgGyVlSD5Ov9tjfDC+FpvpjzyEQ0JBiSRgvw/j2zd0bxDlFqymvq+
qHS7Nmc82bdiWDuw0/e0jT4mzlK+YZxrUOZQiASiVoViGJCY0/BHg8Z4NoqwffYzRucAIyApF1KD
rDDi3FMgyepec/PBbf8ffwjjAuUQ8VY13gAvf4XFV3gqcgDl8O316AE2Vgb3od0ZNptLbdJM9yX+
/OUfCbjWpC6JLsLyMcyigvGl0rk4qzGQ6mYxlD+GyqSR/uVrFNBPswZy3iWreTc7uIoxq09ufWbh
abQtW47WHfsVosHB2EPyZswraTBAh6olhwFkvCQU3QcbEOC4vT95ML5UN/3rLmTJwxkm3/0hsOLK
s+4hA5dKoJbiCvYVnX6tSrzDcUWMD2FRvh+Ibwz+TqZByMbKLiWZUskEvhW7OPDHCmalkC94V4jA
AolTbP5+owgeEy7Acol2dKxFtE+SIEGs4RIu502J8tcKch5VhxbOxMbWTJ9hT08MZn03ZgbftVY/
Nwcflc9WsE3C+QcKMj4yDZ4lIo4rgZQP3N4TZPZjc6wpRTQGtDcsQ4GHu6bd7e41XiQdjyIEmJEV
T8lSFMMnebewKEJR4zs6+1/S9Q+3y6G0dsD1O5ivC+al4lA7VuVAhcrkD/q1Q5N2FWpoQiUzsf4v
WZq5TH8ECjnDl7E4Yh5VwL6xNMKho/biiTKgujj3nFPhAsqOwP2LiAttnh2fFZ8mebCDMBeuQKdH
SnfgPKaw3mFiUMM5kEfe/w20dk36vV1daCP6aw8wQYA2VObVLwVIWCoUOgrEw4w+uGIacZsRzFSF
nz0E7mqNw6nndmJE9ravExTKd8hmMdmPjcvO2GUpHr1C1F4V3EogIwlri2jRSzbKdLSQNHPNQx+X
3pm8iHH+S2itXeVpsFiAu2nm7Fj2dj4J/FMcD6wMucILX07grFbr7AZGiECrmPbI1Mtzts2Wfarf
SQ8SYELOgjR3Eubxel0TMAtGIPM8VDb6jz+2Lxo4kcu4Wh//SI2Zc1vzs+PgP96FrBaRofK+BU7C
edVaOskcvkgHhg6elV1z6dtsGgEGc3zdtHrLI1phsvrP+M2NFuMJ0a3MLxSkhAJsh/KAq9Yc0sMA
lW2dBTNHFFV61P1Bg42ewEtUbpwSQrCAl4JvUfRojnD8sxXTQa3r+kzfN9V0OTftiiG8YEyVlqVT
X5N4qHBVMAs8Lbn+JZ1fXiAdgS81lF78hBInvzP2nEPtoI/L+jTD7jr5bvAYTC1Z4XJXSCBGa700
zKeLQ3lH+gFmBcRBGxqM0b/btZbbhBn18a2vSGgiI8d+xK2iQ1sVjX5q3JrwXMTvjfMbxOWbeQNv
YDkMDdT8EIyr3E/hWA6BFZuSou5cpXxo1LuqNF13kCXu6ySHk7JS08O/Rio2Z3XnVYZU1uYSva6Z
BRj6tM6WQpHUz0s43bvg9o3WVnomB9G8zB4xb0Z96FszMvcK5mAOdZep6sGXCoF1EYzPhk2AguHG
WJp23SlAcXfgdHV0tu+S3NgZPW5N1fFaGcxhR/P9tIkhhlN6GB46MKRVkucmFBGS1FU1jJckPLWH
4i0ep7mLF3YvvRnM/2m1t4HzxHjHYd4ycDudETFRTX1QDxPM2wZ+XOwo5uZa5iQrV12lv+4Fh3up
CkelFtKEgY+q2U50Sc9Yvek7XvS5IeJ6SaqchaUNfJCRhrZO9uoXGi/jgWs6v0EuHsoCi0qsF0E6
qdha34F4WT8h1bbzfaPeB0f8OToXOvE/X+wMZB2elN91hgNpehtqgU6sx4eQgXrpgRSdBE6orXkg
H19w0SSneZHe+IAZEC/DtVtZ7mcZwjDULvh+X98R//9AdVJjOprnPDZz+4AfRGrcipCv7cy3eteb
D9I+qxHVCXivkcKC7w3jSEfY77oT8ViGfU+CAG8vLrj2YEZPN1HO7bCvESfcAwY7WZSejcKi6msS
SRgQ+yfs9yzc1Pyi8gkxu5PIrrJlWR0fU0qBqngcJkbkbLHyB0pAu05fGJMWB+3yf4FlG/KxGwG3
e9SiAy33Ai+WB6SIf0w0ljvvOrcia8YyanJ9tJOByRrxtOUfGbfH9UPNzl2IU9pcjK1UydC4SJNV
0mQtHzY9oNR4B++3a3UfZDu9DR5Ej0LfR9NS5WgSntnhyBNj0ZGCt2/1O2dsLBa7KBdH4JjYpgjS
SyxDEO42Ma4corX/otJeSLgkoVC0ozCFy299jqkz7evH47BBvqrtuT8MM+K+8cACRjbQaWXtTNaM
xRdElDJV0cLoXmhjXAJTXpwQaBIkSNqE6SX7FSPZ0y47z6MrdA/8fwDnHUGr2w45E7qEdwu4dh8w
GksO//qGN3t45IZU82yGAToITSM5AcKaXJ7JXC443FfuAdc8SZx9ryrqVLxZFW4UTHVCRU0Lx/pe
oji3LLqZNG/LCV1PPEXDLUK83sYwYeTFASRf/NsPwnOwkmBHkvqO5ubEGBdUIuMrivPOV6RFmJ4j
wbKqyHuWJsY+atH8Hy4QnbLguijBkNenlkOI5T9DfCCQy2nunZ6YRL6BPSaaDKeXv//14kQR6V9+
1lzmzPocDGu86hv2UVmHYcxoJ0c5XKlmvm8XsZzDTOeGdIUCrwRNf0JFbd+0gJRn4SN2+3aSsH7V
b/F4UwyLbUV4uW4In133tKava2+Dqfb1zzgQ7EchU6HUslom2vhdWLkkMKUEdfmONa3UdyU/vcze
vjYy+wE1cvim/iv3MGZiFk9H/K9a4fZ0P382czSX9m6eNQ34IRZMrIfYUTtVKrfqu83+2V1BHZFA
46HXlEmgfIhj2ZsQ6um+/qYZz8uhIk0IVCcyLwKtq4+UypYvyLFFSA3QFTTwkdMp0FmS6uPRkbPX
TshBIpszQ/TaBEMHM+tRkt7HdvH+NHyG8+9Sd8KyLz1ylY2+2upzw3urib7O+PYIrNaL5av4Vy5z
Anq5wZ0+pj24TAPOOTmrKhLJVcdE/n+urUaKzzdrqvDIoobMAWZHa/0kfFxjAgYnA9HSV9HUEFeK
UHIObPeM90HOHvK9vzlEYYP1rQycGqkdvJLiuRUqPno70hZ1BlAGymVfRAl9+ghpr9D9xyldU7ol
WQn9rAIIPsR1eRafM17gkx3KcQPyMZEugshlGo7I1RwFzb9V/tVfSVpitM4dPO4gM5Zs/b7sA2Bf
zGz5KPK0LftSsF5K7amNh65+nKFQHnTkpIYPiC5C2EY9IXp6P5tn5oCBOqPNZI1sNZ3FwZ/iUp1M
8Il2z+szpnInX+pIPhggLg4Ele4X4dfpDvtESCULeE+i8ak1EMNDuQMNWtFBNWT1oivUTaQgOOXB
mGEVVTf7H0XHDdaAL7/SgGDKPUIom63t2hy+hr2bbKaRnFuR2cGAvbbBrUb5+nq+s9jBG9KGTTkn
kFF6ugMvaCC02TRJ6YaKd6Z33OopNmd4WRH9+87r6yOx0elhHt/V7+MHSDiqGWvOwxzZJIK6JuCw
3m8lj/VVie+GEERooi+HTlc5wglw1uOlUyPk6DqPVje5XT7mz736bGtyCMZmAWhimgE9F7RXcMq3
1HKakvLP6okPaBAJCakDOqFok4YMott8wiSo6XEED7x42OB1UH0kuqCAqdzYmNxUdBVJRW0/fRMb
I2ib4lsLC0rIBMdIu0/QKniMxQLf7loXRFg8O3NDTqAOThcEbIoBkGPCqMNEoUzwhtT9WEv5rXTh
YP8rllH+rKCE31Pe9GK1QuFbt4PTiuo1K8WxBbxKojEc1CGe1P47xTdikXT4PuCHOLuEjt/WmqS7
G+CcOYfYtpfvNAbZ6MKQRHwCmflKlsfiGEFxvXPk/TgWLFgSS/781bLx5IMyrgqc8OukC8yqYj8G
s2wyHHjHZQQV83tAZkqPgSlv2yrruBwzXpf9LXVTf6OQXK5iI6AlQ6X86KWliMPlmVXC+hBR+Cqw
U0++4cgU5GrGTzeF3gNu8oalR15UZXbaFnHsWhM+VDQnzsYgjwVUd8ImWrX0z7vs4/XHj4Lc7njc
PbO88bMnSfby9O+I+1O26lGnmJTJ95a1WKzpu3cX9YmaRa4IXZVptyas+JiReZlGg8/dAwWh2F2p
JLjWjawXACNiIk5KrVay+NdWpAeC8pvpEANjssxW6AetsMuJOUlJjcQOSnNSEOd3SGaeobtyXqNy
s8YiMA4303TeuBD15T6Otwa6y1jMRu0Umi1xBPEIP2ctpnZksEj0deLVpKDVQB4oDE96NapYboDU
e7Iyqcg2RN1bdjSvmb/bvVcxKHzbmapxdmbyDgKPU877PqxYlk6gVIgDXdP+XzR8V72VPv1mgQms
zfEBL7CCwRg2yNuMlIOKFnMNxuIax3wiFQgfzhHhJ9XlLYFLWoRi7Zp44cVq1p9m0ZDlS6pM7L7B
psT6dlywoChkgGzYoJPYK1XwOhL7eAyRZWHrahJ9XMCCX04mIYnJ83oRPLgiMvva1ubyr7Av0Nva
38RE95Z7QndPy7BdYInp6ARUSvUGJeDv4Y9Dd1q5u1es9/29ny7akOeLqHrh3OE2toSlKU4+c9pz
H1jwC3Ah/OEH+G7P+n7uR+k6ETxxbFe7B+I7+vHUYGj0l9rurHXHGNPo0mAwVNURAjp/QN21bUV5
j3VPT3U6bgvlWjNldxYqLnXNz7xjscztDqGEakRSjTqY0F+ga7rq1FaU5lI4AoKbMcF18kByY21M
7zuWJTCJ/1kr2b522QIxVfAGKLxxnwdxXiY0nR+oJJd1uO1D/W3lH3c+JzopZdDDeCjBNOcaxtse
Na5GPGSPvvp2B2Oj2TLDdqOcmVsnygTiGBpCmboEja86a5iLg4ownK4h7606c/cTvi0+PwyRrj0M
2w23NBt59+c7sCrHTaZM/K+EqaM36fHLd1an6LE4m8W98M+8AGWAEd6WUcm7iLrPG5P8kbsYVVpe
SZLajHsdQ9a+4ekZW6xOPux6O+OgrbxDyUbnfZ0qk7Ek4p4NbYJOhBeUvme2vWeS7WYDhYQDKR8X
DSsbPBi45FG4xcX+Vko9R/xVsypRIaT3cGRKtxuTi/1IUATTL/ig/eE5upKIEin7FYCldRCPqzuN
OerrpwPpRcSsPYHCEFOl7GlN+KeBpWpwEvvQHrrQzRX4C9Ir2LdAV6bvn0sSdgI78j1TRQ05RF+/
5NGIvNFOMw+VX6qugGF3+AIX2HS5j1AfJUgl57u0+vHR9EIxRftySX76qxGYVBQV0+Skx2B6RL/B
HncN70MdHuREJXs50ymrEHSdldkZwzN3N3uvJYAk3Kv0K4/TIDbLKk4IUcfJwKK+WRJImzmxDOl2
tTDuJbEnVniCHoBiKjKI9s1FNZrDEaeFtAQ8zoCvPtsDGmK/GNljaYDK08CrN0r3ufmyrgY2DxfJ
8dFq5WfwD3qHxH7MGymqgNqz7iIgWloHZ92T83lAHCzeTTMMRC8CSjdEF14sOgaOFUXsjQC1lPze
JzuUp+BTftbl0IMmSZYra5XGhkcAgqnsiHnskWBABVxalBsxE0MVwWsFyaNbReEhXygESQW2tfgM
f14zxmcWmzK3a/93kEHTt6qVF4PFvaMSDvTr7VPNyGNoo1ixotJPNwR5XWJwodtYjBJ7fusM/OiF
ihvaazT2MGNDh7HhYdpmnr8ZEEaxoe34Mk3rREtMrm5pIHuLiFveQVDQxl1E6CCNCQIHD5DDRxWO
0OSQSiu1t5KmTpm5cF9rQX/9l8V+0O96SIov/lh6VuoS5UY3u5xkPqXGVtt34tNXiqaD9AiEhEkZ
i2pWxk2sLfwNRTqVS2m/6+bE9O2akuwDyIWfvaquPWGlm1rU6etlc5xe3iMO0F2vJpM3ejGlk4s6
98mTs89o+fYiToSaD9P8OkqABw3QLfcDjtMXk7cc1QrUgOE0DPvuUwHdQfHLEQAhn6mCM/KHGErJ
Uj2wfHyfdPMky6+h2sRXcmf2ebF33hzHgQ5PrYQYUZRiUM4J8XcUV7RW8YOZRezs8dfnbVLTAyRV
/3amGeamfGW9gnmmSGLubuVclE1zYzHEx1lFfNuu9h5S78Er/t+veiPNO18GPxJln3NLZ02RcOS1
9LWW4gUa87LsmHfAzx4Mc80EwtypQLCH2iq55smBDGzBoNHzFBpPz+AVFnrGXHKbgQZqpTMX5Zcf
J/gGWjsKoh3e0/XIhLvt0TFIDfFl6SmbUi0dcsH8pjRXqE6LOgY9OdTPnIbJguasPz/IpUWVkBL9
zLPJ2epabFPIol8r7xJOXeYymqlidaK6LlJccfOGB4DjNneB50tLLscziUcr+PUWLZze0fQPib98
e/6GJUyA7nW6zvAd5gIatfZn9KzO77JaNQ1USp69UOt9IutL9Jz+mSOL+INFAfcjlHkfaL+I/Vq6
9QLBO3TbukvnBXR9h/HXIoz+S9Oqnr0eOZVqHtg79UqQ6frc6oy2l/R1LzU18sh330A+bzvya7IG
KWxoP7EfhEwudfDcWGlajh3gEjrUwAGxImjbtNs94/9jIvrTKcqZtawjvT+VW0VDwYXS6naTfyaP
dtzhC75arT92ze/+xdoHUQJDGuO+o3hJk8t4sLkZpIfG96BWwwhxwBesJ4q9ndL218mfhENZz7RW
wiBMqtqiCWd+l/FUaYLT8utXrPx8DJ5J60zR977jqk0tvQfmZqSiV0cvAME0tnZkznz1XqpBPdcp
K6wEre+lNQS6MWSslLHm6UgjaYg90qXR/Tif2nmImC+XFqiUdwvSw4iG0jZzFMGzcqK6T0YrzoKF
NaxIn3HdGyoGIUtrklg1e05aHiQ0DpxAzi6hmdQrAe80Uvbm7ocI+/TAieD3jq34crlQ45LgdNX0
+EHVc1BwyB8b6OrK4dbS+pPtuqzC1Cv2vplVgHhsfe6soFK7W0o18BxmVAGg6FUyOOkBzC/SEMIy
ovWAZOlUDBu3rPhJRvrSrhsqpg7sy5Gn7BB3+BnklTSMvfoHe8nyn7tGps4tdX+ACUzK6kMG5FNd
EQkS1VIDUwozsb/SSGDSwLtBMobHeXasAeJbZRHmZRcQeAShM46GUhJRNfct6Tt06ne/Lbo8NQ7A
cMnl5vLQ+ZHAVIzxbzd1MxjyFr9t0QQEXna4klbzJri+QLBAniOK8qbq4vLX8s/BIIaSUU5w4d7M
I05/dowf/DGU6oKRnSBlRP7akYOXq6/Ab8yl+5WGFtDPX9tjMzZJziIp6FJUrr0FfQSO+zALrVDk
xl6GNC6RIcrOKsOEHAfma2b0lRngRdoZVcuIZjbA/eKtykbgwg7AosSq4WfyxYH3WsE0BG4uBg3S
cahhFlFuFlEILVWvXUCk4GENZPl/zinxwSDw75B7M/7k2r3f5+hMkLGkk+wcFM2uN3wdsx6GXC99
X8/gq0GeNpepb712VDnquL54RanACGEQU0A6G/FY4QyRc63MWcWnvDIb5GciCdVrvzbZNVOv6hG0
13W+Ir8yTOO1bHELg0taI5AMUQVaglzvwT9+wBwuISOQYHJHNUbjPA1vEsPHu60Pkplu3RTdOpj1
G4dbrkxOYVwRtpdYDy8QQiW/Nlfb04x02WSYauLmGUhp2VtWt/3dXsJ6BfTspNAFulqRtwhImCNQ
iSCOqXfdszPbf8prPkWkOf07uc9ikbenycUCQyCHrKaRjwyTXHf2gT4D7kzBOPzOxyTRzHjj/Ff/
fComHka1hcf00a87TOM3Q3sE1Sd1VVgVCAC7nP2saocniSfeGqS9tkWMSE3arg0qaPwUTc04Bt5C
E9kWcrPNd6SQ9wv7J28zl1pQoPdx9btmNxWd3K8kIl81tAqa75EcKbKkBLrdKqm1jcDlTVrNS6Kn
pL58R+B1UX39YEpg0CBfRF7Gc0jARMv5jGKCmdQ9pl/DHlcs8Gfcky1h0N1M3jKTK3Vq37GlCsy2
zrIp+iUcixVvxCKCSFXHQwyZA8aYn74Ny50HVKhelMfZtzgwQpC4t21byCB619qfRhDZFEY6LUdc
Aw5UpKLaXmb7bNsxLwXKME/B1LSJR/1iE4qBeGfCr5BK25nMSIX5AKvLynodJkHzvK5aPUZLlavC
mOzUbrFvVJFcmdJ/YmW7NTxPRd7JLKAZv1tp/4x9LQZ0U3tj1D8f7acJhTZcykX+AgvSRpw9Hmp2
a8hgBak7fvepmFW4N/LPTV8Nf/t4S6kNzPGcwB3GU5sViDlUfr0/IikUS13efLTq6ZIKwLsx0pBW
ZezhJzh50jmLZLsA/y7S/NDBNchBdRuhGLTKYiZz61g4JRQ37S01bYUQkh+KdAC/efOFsPIcd3vk
KB7okgww2XrKDyQCbSnBzAROnn54ACesBpl8CxfUhiuZoUoJBA9//zbzpwC3fjKZrBlcaK8scnmO
niDB4/Tt3PISZuBQSLBw9s476Y0BDkmxCaD4nNJSQwB3+vKVkWHJfR+D3wRgU15o4YisFISNUF1u
GdgRgGwPKp6z6Uk4HAVLwsCvVV1RNUforpPTf1qlFZDpdj5590lBoljyXHYG84bhHdEoMqr1y02w
ZVqfxg9iKz46xXODdKDLt/nWwa/dlAyaB3y/Bouh/DT9HmLJC2iAuuRYByKFP0I3Dy0+OlKE/06L
96TVXsztqTQgWAT0xZiEHR1VAUQs5iMiceUEmLKpRvjOROEQdKGIrKm5jo92M3/E5jjq6WEAomgS
LG/P+lGEr+/PjnaEdfYfrCcSq+0EPG0yU7S8EvCsq8gpyHm6njkn+UFGO6OTUjGfM3Q6W4T51Vc0
2jgciJDN2QA0uIWGj9ezGQuYvoSaEBOqXsizzNrH4Dzi1PxZVkxCXRZBACDH23mNwUNPxtYaB9Iu
ZzSeE3XV2Ja1IfxkQPXwHCgo6TCWG05FxJyUfpr7kzhx3hpu8OiZPx/WDyh1YhtRnPSXRcM2BWDn
MzcakiQQSsxRxgjxKQyl62TYU8DyrjEP9kym8EmIbDcyeHbWyGorS4UfQipzUp21W5EUFeI4ZTdM
h+v4sAJBWzq+BZcMFUH7WVehqhXrXo9DNsCjuGEwKgomRp2bI6pcOEXg+ecIqO+QKkCnGKJ0U3qj
wMReppruMCtpphvxDbBe5SbsNfWKoVZRG6HCT9dS8uAkyNkPgvKOevn/y0QHDnjMeu+S1T2FmFx1
VuLxtLIkczhl/0A8Q4sYq4lbLTLLUSQlWdXEaCi+n1DY3ap7bV18Vdr6YVEJJtONM8dN0bL+/90S
SqDL0UqekodMPUEMOubrLKKI1c5SX0KDNKFGijKLuF3wWo7aWi3V1fk1+2UnJEMrsgANvU2O+r52
4eeZ7c1Vza1vry8/85HB9LlCeUgrJH0rawXIcEnclNQ/DYNpUo6EpxSaEWOZ21HiPYq4aetdpfZ+
1VW09sYc3WF9EUifAfAcvHje/eoeIccMaI1ZowRDPacbfg65KnzUXgI+YFqOHcFSLkvt6cqSL2+Z
o/dbPiBya0J2vU9nGvXKjFQ1y7S9NNirgCw/Fm90XegwnP/Xyb9nWoI70ujNiPpsfa7OCJX/+dvX
GmydQyA68HBQo39LZytpb5bRSMDYRxEzmD32xfUlSuq2RgivckYBEbR9TRq8IqYW3Cplf2MuI6O9
uThNzl/kUFmhoEh45/jPpmrinLbhPfhIeujATD6elbZoz+Uwyh/3mFfD0WuiC2tS3g6X3Hl7VJss
+hIUk7OxVTNl9bIluKQwuXGY1Ug1yc85cY4onMuEa/i0bKaGf2MFmUXBXMiCK6d7fcnyaryRcqFa
LonGdcERUVhKCPByl3h9b6nkNqTgLxEFNlyhHDOPb82thY6eUdCUjqsyVvXwh3kSHboFTFhp/+3k
ct2GiaN44+INSYhVIzACCMRtt2Cnq18XE2RagqokUdHOQugJorWMfokoq5gHL/XUmkrdEh7EWfFB
C7bIrB6aHUcMdQp0R76+yg/RBe91y8smGt6mF6lPsph+E+5x6G+kdb1JJoOVw2t/w8nCXofqjxVK
cpL5XO82beHARrULp/rm3VDASduyGHYrTYqBDcRI0jycq3mMw0JfUTHfFOuRcEeg3EdiePu58wta
IgvtKIEDwg95UBLTH/Kivx8/RhFxwfDahprNAelAWgmeD6tcF1ZgZyM+A1Ul7vGJ2vFm3lvdmEla
vu6AWGL/ONo0g4gpkmDE6xbgmHmUuJzyeGf97vf87MBqtF/Bwx/XoHcQRqwk97TLNwkB3lki7seT
3xI3DU2zN4QmSvc1hFdNj0YxwLMwya2XYzhgG8+jtcVuhRG2k2X/L2eWLL28EvQIZKrsb0ZDFRm6
QnUaB/HqC9uNSomHsoqUR8IdsbmEEsKClBB/NiLtSFbDdOj+XtxQHSPRUP0SehQqQ8FDVkeYsPEj
iZTsHvbcmUUGtJoL+ek9CK+2B1yiOnhJ8NxCo78pR5p6r4K8kkUj2pfVTGF97Biax5jcl5SkohNJ
f0IAZSFpurb07I9GZX6VfkKndeUo8e6aKwQ7Bc0nn5gRXE2XwYLPzoCYxyZdY/INxNoKgasavKKv
MeHpMaOaG0yLMJp4VINMAxfs5WIvkgXF+e77Bw7XKMKNEUtBBgpmO/6prqLcdCxEfJ0+r0N6Lp08
RSMon4xas+CtagsQr2yeSYVm1xNPODiF6Y1hCcnmt+ZZkrMaKWmQ7uhIZ75pHVJcFGzvZ1r69tDL
1WG0lPpk2IEYpe46fZKxjHVTtdFevGiibPnFJzGjAmV6dET9d29vM1qEIgOiEPAo521vfE8aio5K
1lrIWHMmTxw6JI6z890whh7F9lcFcViEzznbMkA3JXTN38X+DvQIIPX0w6aXovfbC8J1yUMeBFmH
XWzFxUyRXY7NoxEiXvahEJRw6zYHjkOQz+d6YqqC4MVPz7h4r+3CaHp3R9OcvGlIQBF5uvokRGPM
HAygOFxL+PImjCxK2fNWzqBqeGMFGK+hIu/MReW6jRwBceMdc91S7bkMopdArB6ckN4/i2xHYVwZ
VdZka1ctIPwvlworR6vhb6aaAuJNxCQhEes85Ji6njiLGWahLPdRot4SgxOp8y/tdJBzmtD3FoCa
sbbc+L8pvCHP6EBvcbJY5dvLwZLMBpGWceTXYdCCwb1QJnagbllEw++IyJTQrwPU3+Pur8J8mzZD
9TK356H1GtJpC1MmlF6n8PU7lG7Np8vgoqhzBNRd3HIUMpugC4WPqKYWSHd6E38C0hm4Pxj5n4xI
kj71lhL5u2CTvFH7CgBSvaO2/uYnYa092mF7XLLNYEhfPLF9jCW/h+IeiBQK6aeyaUmPmh7H0luA
g0oA6v5G12F6L35hzpIC7kUnzdTfAg79jXTM7vOUsUjD/Mdt5Hgn5QkXhoQO9ShnnqlEfe5QVDSx
kztvvWV8/il7qitb7jGUU7nfCqsM7U2UsCYKsCdcmONH2kZjpn2iuNSgItpDGg1dmwvpQoZTDbjK
yUZp3D+rT+P/qkOFOwzHnW1mlD6ptnbPRLaK97RpRQa7pkYInL2wQlt5NzRFvzC7cG+FQVItvvmk
yzxq67lLMduufHQn7dq0DcvRPSRzK0ypdrabr/42GTg4wInN04aSFeA2ZrhuOeWIUE6BpMI0lElu
foSBtQSh9YUTQoIf9XArxWeyBDlnfjJ4ey/R+qfP7Qu8No2v6xcPukSvjLXDwb+zrewTvY6yxjNx
g75JrOUuQO+9251pfHpiKwAkzQKYeFxFsm8wR9LYxVFfdT5Tx21Rul3TQDwpoHZJ8RPT9NSh3hlf
X6lzdDn65cfdbMYMIBCNlGUpPnV5t0wmW2T28zP4LiNfPjSpeeZwdUSlj6IBLnQmhFy0veu5xJVt
FM0SzsoulrdlqEWUmoJFwOXmlq3FksZ+2y5dWDL0QOQHGcy61yzT5D8zDKZ/PzKeJ+zooMgPAsn9
ioVvtxgNO+Y5rAspHaibdniqPgMMzumcyXljQGB6xfNyidD/wUAssE+8/U8Bx8zNFpkkG2RpQrNG
N5gjVB096MENmDlWEgv20oJoSUGPMPCpx9pcJYeZfesJJLWUzqmDJptiWhcskwYa+Q1SjGpPN7ca
PC8MzjmRf5W5vWfezNdb79Yw9lqBu+UVHh1AjgioKk/ALouIu6IHzoB7xbpajzPNjDhGLra2uimh
yUAImAmzhpFyxh8iXaEvfk9LD35igLASKekM7QypcMCu+nSCqouFS1TqGXXHu1vrh2omIDQVUpRg
D3B95JkjGebftEayIU11bs5VeclIEONk7FD8aOWBuCIROA+Kg0bG9SHN428qLaq6cep7efjvqRzh
kia+v6eR8GgxGANiJ+q4qfUkLfdn9yr69WUGjyP1XAxv/NE0PRrX+M/NFx20s0g62seUAGqit7yS
+bnyxq7JZugIlD/CzQw/K6I/UmWPc+MW8TmNwmVS69RcF18J6GA/mfnlpe3NM/7FGQy7uXN1V0iM
BYOe/Mi8jKw+Kmoy1Bb9799Qa0Xyuda5qIliNXf5mZdhoeA954S37z6QHIF71Fic/s/pkVguiDZt
Vyu884i/lG/g0G/9R0wuZkiizOPIcIdfIXSgKVssgBhldHf61X+z0xbHtbhp1Agh+1JDL1AOvlad
zMyJ6JivUBui5XuZ3a97a99S99HInAnzD1BEmJq+IycKpvjl5B/kQmHwn6YDNoTP9XcWA+Ard/S5
isLkd0orHdGr7/6rGM4L3cNKZPzna71KiXUgZB19PK3IsLD6asFa2Xi64f+itCVqcvlqVlqawK8b
PB0YRaYS+Vr37GqX28IIaByAgwI0nllmgpUXmFng9ADVsGqfoprxZzebHeqh1jAndDywfb/OtE79
YMbA4Im5dhC+mfYYPsvlEAkAobpE6xC36LiCU59S6dezw5OTcknDmzU2f5etsWbX1xSoyJY5I+Uz
OCNM1nv73e9fKaHHs5Th79qAV248l4c2cLHLzZ8PwoJ03NJTBx/zD57eN2AriwJ6nP8ib9yO2HyW
GmvQtifxLxU1SOYazDNgH6O+/btbBMrNKM7USFSNnTG3E0KMh7abHqQdXylonBSeLEudtfBtDDx5
swAyUMF3/ReN08n+l8U8y7KlSO/iC5/6rGgeSozScfzX23ExKuIEuBNkE3ZupqoDBog4y0MaMikk
WzNxYtNJ8/zCqVfoUlZrLEZ/ONyX/9lrlp3Rxd0BExIZHBHC8iiwYnnOAF9cMvgeLUg15yivuDyT
l4YUBySt9/g7s53ObF4r6IlQGuV4tgULS0iiJ5iwe71Ags2pGwogkCZmT7XXsxmATmfCq+3jpjCJ
EgmfcW6ajQk+ScLXCEC086iAFpofHeFzyOitQVB1ei+Ah4yKG91GTWSwehW2REZnqr9rw3z2UYfs
12rwTEOFnTo/SLkD8wRYKkLhbpn1cuhuY/KCWeLxzdA5gDleGBffK13gtr8ABHxBq539b3kbS+7c
MFcgmXDINZ0OlvBxYWrIb/kDs54GBEEIjrurMxlPXtLlr9snk22Sr+PdPPyE+SzOWW5dDgOBC238
LdPFGta0aE/N+vNRvF0FRMva0uGrlOEyenSSxeZ1e3P4/bF81464+UboIl+pdIHKss12iYwiIfvW
JT6lWdwDhBFbYxZWU9P1ZvBgnQpzlVE5wJC2wHdzwMfu75Cii8pF2SgC9kXchFjAFQPMBfjmJs6s
d+/A7f0qzvOaZACj0wcGCNPuWvTMAQ7iT/ClgHAMM6u2XESKFld7YSQbQ4xrlj1g8vUOEEe4RNd5
+Z/npncbfVo+9eieE4hfctj6H/3/dLsinca/lWM7YdbMEPqB6WmBEV/XmdxK3uR7NxXHSu72UZxH
Wj9pE9EOhOoGfbOG7Ee6NwuyGuatQ6G8ET+FfXE3twQWvTO+gcy08yMPl6BWdeT1lFnuOnbPMQnY
2xalw/TyvNGw7+nQz8RJevxQ3PM6yKvCabs+s84+4a+NvqD1T3TH2nmmrGeMS38I7Y5BRnnXxSJr
k8xVgc83ZcpocfHZ2pcfDTnFUO+1WhG1aIABVC4nOVdSsWqSAUmYuyqKiny81KT8tS1QaUXa5FdN
/LRXho6uqT8Gp3aCq1/hUkrWV8aklfY+r9SzqMIuJ7OGbvNShQYw6USJoPkPXW4b04z8mN4zXNDl
Edefc5I5ic4VIhlzJ/cS5iDBv9USp73kVDbhKAPvOgJ59mqOVmbHfeFRPqw0rtJ4hV4HDtFb6ZCo
wJss1B2OH0QDhoDenawz2yOWfY1Hnx0fxbwEJCKuH540h7Gs3V/nuOH6UoFQH82o1yuS3Ptt6oSo
VMiwslTvjGTqlJjECN+ms3wEcbzGMnP437lxtHncUVy/vlkWlB+yRwtyu6sC5hMZOYaGjysHeul9
0IahTXd6Qq8KyGh59j7ew/xmUl+qIAUKC0A3A0Rpj+CJulXzs8tw55f7LAbka570ueGYdtxZcY61
Vs6M0dbJcskIIaCh6EmeBBE/83ow4Fez+dLwmw2CaHAmxDK5qrMD2S+cifEgeJ0lGl4bWVeOXcnG
YsTX7T/PVFDFk3BkQHRNFx6IEl5IS6ECWyLsm7GQoTIjPOdt0MZgnbkht97WTLPOb82qrqVwEiVK
y97jn7i4sf5TvG1TLO54DhIKIpEqGu/imdHtqVtO4szwNjx/2c4861SuM+8BN7PjF0oJRqjMPQq4
gTARJ67M+CCQ3vYwTal91TkZUQHqy8ioRBvnfAZzE7ppYsVEQP3yCmXnLz73jOSMKfUCRAsNIANL
Lz99GWI4FezoWBCxKScvOtTBxiAp6Qf1Kf1v3haBXQ/qirw+FOdGYeFK0F0qfKCGSCquiQDPlYkX
3bZz147RWibHH8oqM1Fm7hzUhJPrwHjEzJIkDoQ6kd/3CQMsmmtDrCdPEYpCt+uTVQwFaqWgalGN
yybsNWMJBazYPcnikn/fL+pMmM/ZHfCQwxHzXhC1JFgonoQrzunBX6Fnzogg1sxIG4G9CcIwkH80
M2QNZhHPgN/ipJePOdHFjtgWPnKzYoHuf8M87Pz9ZYGFBXF/QUIfnjioESRVeRSl8N3exjYzEE8w
oPTkh7MXMVJ+m1VLxakTL5bY5sV9TwxlrhDnharnh/cJKg6btnAHH0VudjJmo8WuGKJJVpsiSnQY
NgtWSiYkALaSFKQvF44ub9WkDLnNGSEy7sHUx9sdHkFN+P8HnEjBCW315LePW8/VPaNuoPOgEVLU
6wyU51e+Mmxfrtf57lbWchnAudqTzXu46mPoDB/qxmfXZTAsX58vOVUPildaQpyCyIkN18EtPOEE
UT7exryQjgm3oqofx+Eg+vfhLqiU8POHT2BYSRNAXfJtWhhN8NDJkhr1JOZ4YMEA6SlmyAbRgXoP
l6MOdXs9tSoR4ICYhwdnhIs5e5GarxD2qs1aF57MLlbOTv8W9jeK8mb9syf94gtZuwhHZ7OsU2op
MklDYnuOGdOvYpdZWSFkLjQrEKzZZnOrN3Gj1dHDHFyVNsqgD78TYExM9PNKlcSu9PhsTeeyfaFR
QQd32tq20GSv0lcuC8eujEr7akTFRJD51JTjIN17jgk36f5Gt8+ICWLMCR9NWaobMjfXPyUGl5eh
XVM0bM80FtDOIx69C/i48PkchlZLhgmqDMjxe+fA6Y9eRJ/Met5X7mAHOCWEwARrBc4LqmNGNZ9Z
G9zQi52HGaQU1djvatdJRzJyuILkaN2T1C/71ZF/ZpgZc48wL9CDgB413MpR1M0l6ZFoWr4Lzdel
fx2shetlSz5Z+67yqLehM+YM2oX8cqX3uYIGY28PnS64Ub4B/YzGW8G7fecD8Sv5FXMkYjqgpRE8
JrsMsYgftiTOGRw1F2zoFtQlYW+iFlLMf/in9twpDn5YTPnFDep//k22SDBdpU7bQHndWoXWg7KQ
6GseGyuXn5mOy1RP1SdDdgr/Ga51uFCyquTYdDdOzFdeKmvDMZ3zcLjgrlZY3hmLF6XGLTGAUFle
EdAP7XmgGeEDM7gKvwx6VdAfLI0liLPV/nQpb2LFg2CAZAc5BoPyiAvX7Sucg761yBOnrrQ7z3xm
oOv8naBFJ/Uh4j1vrRNOBtBQ3YaqQYyIEnLHYpW2j6yJzSMXImMuhkrQNbqi/0cQnhpmYd8dlUmj
v+3vGUi97PlFx/cmB9nkhRmLnJq7zZ0cZuTCr+6Vb7jQCm4cJg5byUI5wjok57OS8gWmWHlcXNga
2ZAh/UPKW0syQKqujxtsQbwjikFyGP1q7zzpEQXe9VLQTThUrzRaBF488GcF61XL+Q1hC2yJDAmf
Jc3a+nQbDGftrJXVQMNJ9DbtSI4mB14XyClBkm8MmW7LpO9C3cS5XTy15oXwh1bY1DnNBTD2Z6OB
WsQNRReDZHCYH3SGG7rYe0z+FncgJICD6C+pObWS9xHk0qfEjlTY8eJDFD+lvtt4Qo2E7Fw28qYP
D9Ka5dovAzBx3Si//wEg5+DRXBFHdicXva2v4WQG+ewq8gVKZajCzZ1S6Q/6AHpxh2/JEJ5Ts5KP
QMVhK7gcbA00xhQPQ4GQ2FiDpfvf5x6ocB8I2psD+AKKaDT2r/dOmWpn2+V5rkOXVgVyC8eFyS30
5EPHlZV6nMGS95kDklH/AVZmQ7dxp+HRWszvM/EsQfMn8E3VeVnHZ4vkrHXn209+VG5MYbeuNJZs
UNhnv715cek2zb1pf+FK6O7soEEk7mExQGwfCmEegRRrD3LNZ9a8IVOdXtKUfjnyqXk94FLGVfdR
FiOtanHuB8fE1a/1eGnhGQS2u8Tj4Yq9htFv7NTmhFVvL/CoQFBh5i6ne+fePH5QwcJCHXS+vmnK
KreeRx/Or+bw4/P84V2f6ZZ0SjywBrljfLDu4K4n+QwSwWUAlxjyYKi79hLWtuRWYjMYwjxAAiDY
vaPAlsvsHBbHlBdrn2vLrXVM/pKXHcKhRn51k+rCPHBHZd65Mk9HYlgZDkjZwjjMdhy1ajzuKIE8
e6nVhhIDhbPppfvJBK4+Dx/58OTlxqAebQczqm/mZHjo43+uQGH7ZyatZJDCjddErhaWcfCVnqxg
7aMIQkhYLID7ZixkEmOECe2O3kCH2FGDCPsvZSSafezUwHduDHS+iREeQh8+Pz5+DndbmkiP8GEX
4GruxWaMnMCdxyw9sXWJ7lTtO83tCxOHyodcep2ZFLyvRwu2mfwOfcWpzLaskMjm9O4rGiCoQXSr
geAfSfDZDacp5CjVtdHYJyZNNVeTCQqGAEFODEImPSFJ+qGCa5NoLWMIADcIQwfJ1qFTW5+PkVBJ
fxV0II2DfLWHZn8tSZ5tGc6kcFSD9KdxHPH2bgi68/WKk+pY+4rUzCeYXf5yvJvupr9sF1LVM+hb
sBss+msWy034qjQUNhluhswKwDoDoxQe+Vs2uS6bh9EJvPlitoTe8ZjC8+weJWJoQ7dkHF/CZTTp
GUfLXsBUePc2X4Pt5uqiOaLoqH1GLh9BT43ytywQJSe921CwiWFSRGG16I6DJsvz+tr+mVm+5+e1
ryaCix9YK3ReS01KSRPrpYdDF73kW/teVJSNSC7/aoHeBgFgePYuCekNpYOI7j5bBpheYWc5hPU8
1VfvzAWauF+hHaHkCdNP42feY2lFWQQaF8gCmYYer/R1mGSBu2UuiRiBMNy7XxWvdWGUvWUMStnx
grEqabEhoUUMQyN25kDGcka/eMvpB0QPiS9AHduDQe9GsRKGigMpY0mQx8FPI4mh3f7nXRfNrec6
PDBZBHEX9EPP3R5wJoM8tWnRSyW290Y/YNTftAxtKE/S4G52m5jOcNJqC4/tKzK3W+x8jXJjLyoj
kYV84SEUVn45tn9Pbm1J3L1RG3Dhk2u3f8vLorbrzWUA41YwGXbmPXz3buZRJMmRafMld1uAPOkb
td1Vb52wG5eVCjxK7oE2cS4lAzrkjR+2a47eAMN6Vs7i8wrUAABrchFYS81oMTEC5/bP1jx1DQT3
PMaPSsdk0FfsD4l+xyec19T76dD09RIBL0zwRxilmCwWrUKTQpIwBEtgIdmdqYAYTP7B+Y7emAR2
4uINsPYNY1IK4MVYxdMHqqGopdNygDtgr6VxhrC8OYm7qSwtDc20b3b62lUpg7xDrKeanz/b/5Et
tZPC6UwHWaNAhJLyHgeAVI8JZj1kd0ZHZ3+t7KfM+41Y5eFOgWQ0ghbqJsfBdqbnL9vxwCeOuAnY
folHKnRPnhuFypseLkPwu7RyBAa58OfChG3AoKXEFKt1s3NG9s94un8JgngLrry8yeg/qr7PwrSR
qklXXIQdoxm7IzgPl452PKPXRUkG39ZWtDssrGnK+4g1etctTHMsSERSbEK7Pe51e3U+cxu8VHFf
1lLrJxbldcGnk+ViTBfBBaH3Hm7MbUQuRMjBbZx+4k2tw99A/+eJNWXbY4JEKilJ0Iz/a4j0YE/O
76dxbcNb+COlkLXYe1mmLj13ufIfyqKUay6ZwU1redqanxllE4/rE4SxndbqR3Q1AFsnoIHPiCBH
+1HULzBrTDOS/ChGo3+N0WMFpYD0qKprxnptGZvaqHzLYYxJDIErDlPvOEFYhFnEqsrtJvPWlpiJ
fKEtA/3oxNDLNvxZurA7SSdpNojkNzQ/Mx7Uz0vaODMxMGclMuLsqQmtvzcUWqO8N1Kc6N160nLd
KlmLZLOiH+RKsL8Ut6PzvVdY6LxHjioYbWZCFDi9/rEerKw8A0qryjfEi4Zl+GDcA72uc3gFpbM0
j6zvl+6HJ/QadNiiaweul3uB/uW9SGKALBXhoDgXgfHDFLDArIfol4uz1ct3Fav7x8AgnsZ3ytcT
xmEIB/wy4/Vmw/Pfu578oIPRZ4LvOcmH7ukU1VKn8X2d8x3i1+v+noRFyz81Dn2s/x6IqIU90ax3
flOE4BpbHjT1s5u4gMW4tm20nhwG2+JnebPAuXzRXX3Nr6v8zuiBva4L2oLKwNH0hTYU4O8fj39F
ohiD2N2io9h2hsnWlJEBPjEL0DKKTO/zcZJkZx5YI5ZuTTtO8RBq7Xw1V4j/iCw5ZY8XWtHPu3at
Viwch0DQuhJEIVUIZ+AffK4VWnfnaV5JVHQH+PT4iPsYIaVhp+DnuJXXDhkZFXQRbrbf0fkrznE3
SYciWBLwmv02iJeF50SzjfQTaJf93TObnz0DNw6yXMF5t16VQiGuwoijjODV/0mN5KddvzMu1wyJ
NLqJRSeM4KvJowKtd6xprgxhM4aDM+4MS0bQIXxszWNy5AsL5qIFpIcajh3i5/AuqTUY6hEvKLZb
o+sVrVUOvoI1T69c4UECHcIlJJY6/0wF9mPErgj/coxLwYDUoFK4QCT3dtPi890oZolGovHHC48a
g/STN/JpUH9HvsBxSM5lPxKEYZfJ8sAs03Dy26n3iEv7/f1qWD1DZ/tVpv5cYqu562OSSO7f0+H7
FBMH5KbSzG+xqnJ0E6lscC4VARSgp2plYDCE4Cxq8kG3gaCnW4gJAA80rdPN+ve0xxHdJoiBz4VX
GgmE4nBDr3Kitur04buxZHpnF/IA5RQBAOI7RI69+IKv0Tt9AtfX5JLSzXxAsxsdWVGGJBKnM3oA
wPuC/kuqBEFiM2b/7ICiiOOQCENUQur8gOCU9y/wOp7/Mv4SHzfXYJgFsIeVTgLuiMgBJXe9bzIW
qTzlEyD6nc9DOV/IwU/16YgTJLf5raUXquMOrLpvRVHf44wGfIinD54ywWdbbU9Ukd50lwkvCIQW
ZPvfnJIeokspTQncNDV+W2ikN95E4Wzp2cXqWViJDebhT4x377GLDe5OkjD/JSR2DqIYZHQG138c
/6ioe9IG9WkBD+U4y955PMTxglA1eGqDcmrH8Fdfnh3J4MvYjGbAS/L+vmflwbTk66jXvlm8GTnU
jISAOwB/Xzg2noDi1w1x2uRIkHdRzMySfSWWhhgf40PzJaEpsHfbUkwoO2EcipTer687rnVctYdk
qowQu++omObP19DAV8fxjohbYMB9SHr/wP1aRhpw0+0OkRrGTODbGkVEMQqRa/z3l7TvUhMxa/c8
GW0/jYnv2CJsK64ttpCahpyonT22/e/f03ttKrOglP22/LVSrKRfrJ6qe4+Hw+mEQGPiVCJRgujf
oXAStHs3UU218kIvzVh1xjsJxn4WK/3kXV7QL1oXfmZxfNk2SeLGxhtDVgQr2mgeAanqX/7xS/rZ
4j2ARtnDGa8I8VfhmTWlNInMQuDygHYWUyf4mDF2HlwoJAC1Whgwvt3pcVCZxbXK7wfGuCC/PxQs
tdrVZCGmHdxMlCg5iXPaMtYtl+nSsgpFOvQ5PxDyxe+2jKZHqad3nkfUhzahOWrWezPSSlE0C1LO
vf7ZK0Yu2HumkOJW+UluSP+GsBuaq53Q1OGBIDlyIdxjFJoHbGsRucGIyy0QPQW2rw9VlgyengdW
EzyVlyT/StpAqQ924GIQ3jf1+IOpRYTW8Kpg9MwglvpQvbrqZOXKIee3s0uuEnoFya87P5IVUopR
fJMXRVb3FPcQk4wG1Q7wkist8GU/uxZSn9wV2ZBo909vnxEGFWtZg54VVRQ0dGgBPNPYndV2BwkX
LY8HfuSgWjwaXzR5SI3No1JCQ6Zb3QUZI0b6fJ2PTO1zNmnsbdyw9O8lYhz9vTITObcg/IgW8HVv
U2It9S8BQwNcvDh7EuaGT3/PNN8OM6yZVs/VuUlyTv3SwpggexnvbuQnjVldI5aCb7IG6wOQOia2
hjTRCkgtwE1xDwlXvCiE6aMdxGI7I0ZI7PNZunnJupfe5zxXQwat2nvMcyjTZqc03tQ73KnWfIHa
h9waYJwo5uVAaEE6SEO9A3WLznczkl2+Nx4klfcNY+J6rl0jjTU4T0buiUOxOG9wWcuhkCLhINb3
99mwkKxFDN82D1HenPEFYkQBLfUNozKn7ekzGHK8P7oiilRUelCnNQ8op7DSwhwH4qeZ+Xk3sX/X
cO61eTAjK/0zR1mMDwZ2vJehfy5ReBg15Oi8YFOQLhXzuOXIY4uMu6oP1bzvhuXL9HBzURYwmXJ/
J8p1ARRH1CTgtj94zqMu+u0ap3a/O0a5CCx5QpMGRQTLG5K31jeMEcrQwPsEMgjkZB1CBox6QFBb
B3GgHY43h10q/g/MgdciKqxZseme7aJ/JNshE63iPp2quXZyk8V07JRooIMwVhkVypwW49ha1jDJ
SppZDzuqgPmgc3pvf7eIIy7DRPrt/kI51Rs0zMiCMHUo7E/MSdlnuNdKXJ7GwOJbR1XsrEkppKs9
y1GhYXEVn/ygbzKG3GnmvJl5LxsIi7xkayaT0LNtTXQTaV7tDrSFMk/dBShUwg3AHY6a1Wxt8des
vA87iKSuf7G8ShJHPA8KBYo4V+MT2xxsbB/cZ4SOqx9EC367CVAOx8PYWfhKhXNqQWv+FDH2RS+l
rEvS0s/VkneLk0QXTfPLWqcD/q3eooQf4hxQT9LaOydVti+RVulpsADQEHz7ad01sQESvRL0gXZw
Brdok4FhBAUo/UUk8dpaZrW2tOtiA37tGg7dvQv46wb/IuFeF1SPdlFoCBLVmHqemLVlnmgB7NUc
gETargDrxw7KRttllztFFbnsWPmctYpES71HpbaxSz3GAu4F+SAA207mRxVMbfFUrWVJpMzxv5EW
5ytGq/h/Zsz9QLZH3oL7nMrfjJpwmTUbxElfd4EpVN5aEGzv7g6UXAsdE9Wdt1jCniFwwTbWcfLQ
P++JLpfiiKEdXU1V4fxgknzzB03OGeFJbFmR7odndLQQo8V8J5gaE5/b3shY9Zc5tWPbnqA5aVqW
GRwXLzeXXdivVG+fsr1C9mmee+eC2d+PvYSo7HFagP3hKyDD+KC7cn51LL7CwYnVZCY4nUEIWHZl
WNfoqaaxYHU964NjaqQdQYR/dcan7oyVJ21igz5YKWiW7ohW5GUMbsd3D6e9Tuw6MkluV4KVdXus
1mTKcdby6NcoRoHLy77whRpC8B1SLyRyKdYc7Oi4qIEBBJyJqpDqo3hQFYrZc+/Wcfcx0awPll53
ohjgQCOMrwFXCPdHEJm1Wj7/Q91uEs7jCM3c6kA7ib8PmSMiPCAlUtUy6MRyPWS0ZRlOWqMzdCmc
A0X315UdHCb2byipKa6cz0kGExNNyqAVKswaH6XuYQ9Rlkymin2QkXS9Y4SMqqutA0z+VpvL8E3E
H/9KIfb5Zp7EiuoTZMgNQ4i937gIZoFLoF2uJFCSZ7vJpRWvPHivb4GV48fuAwOd7JxGHYachFEt
+qM+DKn/TEltvLd6k+OVgalPyQGar5Q24CU/pF045NyshpXV29XPoXwNnA0CHEIDhvo9P9CNmLTb
vDNck7t3lpYMeZSkJPnN0QXVuQxBI7Pkg8LWzFX3JdlFkHWE1mKJjKAo3Ng7guPXST6hDzDcox9H
Ehrq24GhRNlYhId6EnGe16pTnwULLZ/h0nIgP6RinraffBO3jDpZDO9a86WvvO044mNlsEt7nH/6
FNWap+vt0Rh4oqLxPNOO1aKHilX9doff3uy2yS1OkQ1nin5+oubo38+N3Pv/E1JzZjRErzugQw60
A2TC5iRc59uT7H5nC9X27rH2iH2tpn3uuHCF77xmSeQaz5C+dXrWvFfWcl2foqV6DBBJncn/vinc
itfqtEmS8Pr5Cz8Tl+b3DJjITaGiAfA/WcFpmPYUbOsLJc43qFzPPu3eXA4GCXGgnDKHN8dDny6G
cM4BukcrZ9/DeXYX/xwZOgYLhoXcMTWgqUL/7YWcbOUN9IFZwReV1B6cwgPQQpmej0+/Rm9/i+Lw
L+wpk5EOdTMJMpUujwSm3x9kkw6dpqgIW0uYNOZsTOpiiE2GFzQn835l5ceybah2Y/49iHnghWUS
LbzUuKtQg8SM4qAAfZgSmFZU5uDsxobvR4YxDJLvMZzzphTMzcu3CaymmQVtI8kzB86kmsT0JwcQ
LGla1PR/CPhwu1Cz9VOy8hySY96u9rqgB+/UNqQlnjjW/80kqggfpwN2fDMEf1/TQGqBLAc3nB1R
p8vvXfvXPsC5OJijVv9c1Si3gPRjsGzPZlII32xmLLl1nGZ1IwCXIZLC0GbxfOI5xFCU0BGnVPlB
IAqk1eGrtU43NWJs/zEHMRFX0MqwRH/evsJi7cQXFYh+oPvpmpqGC7yRwNf6+5lycyM9IoVV0yBG
zTorpi9hvAspkg0OBAsJO8AlR4JwdPFJqsa6e92KGIfg/DSuCHadt1I2AG0ktXtBGoYDcyWTTJM9
IVVfSo7T3/6yAfQmLaWJ+SMLwHK9l/U1QvSuRpeWbPgqhmKmDEeIduuH62vyTWr3ToRRI6PewSEp
avInXfiGOGa5tzqk3VjsaKrVmC9FVoAPBa85T+TR8uHmYOjrpGdVndtvBoOSt35JtMMWWsrG1G8k
fsvHPlodwnGGyXQQOfawnBRNQdU7NIMW4HSV2Rztl3imDqf3QZz+UUBxv6E/zCS2MQ4vpc7hr/Zj
7Y75z7y+TVJ7U48n0HHpTZoZwrzihargmeQue7kipTvZ+/9vJjQ6BHRC/ldeYsvk4nWWJ+ARV77j
UZf5vBxWIOKDqOVFdXc49pUKKitAMG1FaaC3QUhVVYyB6HP26l0QHfaBs70xC2sLqr/EE2yYyf7t
psvTDpUUQaQbu4g258kQvwBqK6RvUZBq6f1jCMf4T/KHBG+Uk3v7FvfKKYmzI+CiidZIGvhcN8kX
2EJSxdbhVxE/JjGl4zKboKWcbkBNoh0BqGpdOgBIhBa55rLkm1kCivnzV3h9sCPydROuUyhuI42F
lp6vNO+eXh5FEG8avBn6vShtMrhuJQmpDF/PrOKNCcU3CLGr8X2H5EMUA4nhKJSqtFC0LAGkh9WR
cUXM0+f/A4e2Lv0GcLuii9fu6fP/Cpz4h3JUbGvyiZ7J82IyaAVgA1cnV1rdxuL4sKEYBk84u5wh
Ie5aX2m5xXBlB6WguZX0GZ2KRUH5Fa3B0AjwdeO9s6ZXcn7pkjL56D4i/qsyIT831ffED6CbSHSH
e4lKtlQNXAHMbOUsR+1qVuCvpshRRnTva0TiET5pmVDLqPX4WsX8FqSsKnkwzb+ifcli7zgxYK4W
wh/fLeilOHccaa6cnsYT6SYMH6U8jeGPPYPM8Q4FGX47LGopo8JQfAOIAxbFRd8rhciV+MMjRkAy
ximKQkW9TsKvgHoRr72VrbhfAFX1NGT5skZytn5iuV6eD4BD4pIruvKTS6mj4LnKAm7CS3Hund2G
oO/OKczcrqsp21i4Y9QlTngBgZ7EP5e/Ld8Z796jBIqrAOpAZzYLGAINBJ6O7VwPUaIuaIq36tRP
kmEwgtI2mDi3oo/wHVasWMhRXplGUKi374R5QpMwgKpz9+38ZzMFM+1vOpy6zyXw7yOTRoPBOxOu
l2Z5yT3t3q0SCOc9UrCjDwasxYNvDdnk4gylx/eq3/vz2n8yvG6gnJfDA/TPhm+1rNhn/c3BqIf/
X4wBOa3B4BBGz3AcW95iMBMXvWpgTvo3xYXf/YjV3aslZVCBsumXvFqzlRWCVbCqR3TjmY3Vf9ap
4OtUL8WVS0MraTXr/XecaQs2iB7yHNZaLcX7vbcv2s051JTPsQDs5DlYD8oeUQBB0/UBT8xJ7OVl
uxfJj3e4wEs79Dm2cVIUBaoSyJI/c29Ck9cKv7+RhVUErAB+1GMDWsh4YFuKFWf4X7XtGHjL6FWq
Rm4AFwP2AiOqMGsjqwsfHQsAtQrY69bxniyUWRah0wcolCNRZYMPVXLaoRwONal+rLSyQDyNUKKL
+6nVgPOLsbgYg5wf9mJKE/wiImZlX8ITUyBBYnm8DwOBrK0J2jsZsLK+PUCMDr6RqWBgCO2iCK2T
zqocCblHE/WhHA6/gyzSoDxzBe/vFvcsznLjInn972EgI7oylYddLMSM9W+XxAsJTBd5k5H1UZx1
6IZMMgCcQ0zFuyG4NM/6eS2Y5iaApT33ffK+gaY3DXD5kxkZ2TPqclGnKhjKoq+cclnLfKTKsjUR
TO4OCJcO2ghzDmCDyFuXg/feANDr+76U6mdJG/nUMZo6oXrp/IxIsGUg0cTF8bdd/1Wv6aQYWd6v
AoBYboJMmj5JKdaYBRqZHYFmdPrsT6Hz7ggXmiIWXjm7DmXn8JS5VR61C6OGYOGsL4y+nmfeDeNW
6gLiUCdq/6y3cCPDMEW4D0su0cxwXfh4oKaEaGVFJkCSOAVDE5wjTZf3YTaNEwnhYw8YL6WUvchS
qGGvw0JsZMngJS0e1Pair5AsCfYXOE18qaSQ2IR3V8XjL3x0VpWspOPfa2SbhqewNGslAt51TRuQ
FZmzlZQaWZwR8HckB83cQJzkdnPlgEqdnRoVr/VtO3R3dMrH6h0zPodXVYA84gKJ53wKTNuko45/
4ZKC5sp1Le40YhlgiUyd0Hk05/epJbg7aVSOplwn+Pt6KB9EEhHxW0fhcyhb+VJe6KzgfitN0ZxZ
5HhFMBnVtcETiSg8ajyK4CZcMuIqrV3auKw051a8VblUakdciWxSHLul/EMqWR95RREEUSZIsxoq
nrIpKtbRSy8u0WLLmtQ5S2muOtwy0V93Q62sIgprlOHaHl/QcJ98TpASE4DWIZm2oL66HIk0hanZ
w0HdZNpXXX0drzCjnCZaQTn/d2+sRESa7m0+o6a3/ll0saRmD1TqAsS04FbKvIMK42uB1EGmKW/2
yH8Zckb7pkV5WLVA3eaGPi+4t8OYV+JOsq8C1OpFDqKT/A/S5XyYFUkL5EHi0JCHsk4O4tw0VEjW
nExxX68OZlBgMoIotZEj1ySaFyTYW8Fke0maeK9vp+5ltZhm6YQ7ryf67jDfKEZhQ/JEihzrRZwZ
heK1iSoFapjX8P5dw/HJyH8qywjMcRlx+jlKVk86JbgjLImzBrvmkc5SPHb+jkXWc24RhHVKYAA/
vTyiA17jSWrYjUhAWtby7WxBHXTN/fRQ9lInDpJYlg+h13MoRa0PqRml6K9+HyWVwOXhnbZ9AlH3
BswvoELTF1kAV7xFLwIBzIb92TiFv88YbTvCyA6f/9aQ1LRO6KF6Mr8biBPnwCuudXvqjY/XrnSp
/PCEFdxNkKXL5oSxOtZmvwBE5TIw+rIm0MNqA63e8cTw8tR0M1f7f734cOgGuiX5WinVSzkleQ7G
nPRQbOeJdhq48cvR0GL9FRSWptgu1xbyoKruxWYBrWcO20X9CvpJ5NCkUnJbPsDaR7lZ1P+jszyI
vKHRzTe5e/O7Es6rJXmWzcugETjF3dizdiXkC7ZA7gU9GmVsRQKj/nS/WcLIbDBjRZ7elnwpPRkn
a4WmlEz+jcGo4wnSM++NGC0fIACM6aC8W2KihBMGVrwxv7ES5okqn4z+03e6/g/WJfjH2jgTEuJV
hsMUOEsX186+2H8/nkzZX3oyUEH6JGsLPeubK7VwhVmbJ3nj8Mfi8ugKUANg20e7DhpcCGv3b5px
KNoIjQ7lb+gg9LHRi4j2fVEk75L0c3JuRj3vXBUdQG87iLIhW4QBX0jHrN5dPbnehy9dEG62fAoa
IDQ8v9uixNCLPh3I2AXI5M1QeTPpT98q0JAqgw6+5lU8+OQNiLz3Jn6WI6mWoq+yxf+e7XWr6naA
RUhIcxzm0uWxGNvU9giH0i/LyPX3w/8vHY9f1rwB5nFXV3mwADq5UDNflICYy+kird7DfOlvs622
vSopVi/gW/bKGpnHxIhwWdwOTdhqDqY4eg8SPo0qbX9MrpyKG/ZguKbPnsgAVxBrfJznYLAEBGUm
TEwAUMvC/lSrB9+Hk+bfM4vH3YI1cL93M7ww1+/83vGh+ufGyI6wAwbR2+gziDaCwSW4HkgK13EJ
NX2nkQVkJsR/IylxSs1dej+qv3IR14pP5LW9ADD7NBcV6AZc9p0EMIHW7m2cRuWx1vaHUKhGd5LA
h2HjJg0S8zX6X43PsOuQWksm4batHieN9glKk21IVywXlsZwMLaMUaRhVANh1K3+ew+tDb49vUyQ
yIZHTckLa9wVrgUY6AzDwTPfCpq/hPMnB0jCdFDBwFY0uNG+cmQ2lvhV/imdw+wzCSx/h4E1pTQV
O4IsBxXQeM4MGHOYjYqEL+l+miNp53V1wMW7fZme4Rc+kd6w+0fJMVqBz+Ey46IDD6MrGqQftHW9
L1NYJqCUg8URTyOOt7KrwWyy5OkXbvxQkJT8STR1NuBZjeQ51G6hJ6jL7/7x9+CSq1D7YvENH7Z7
KN69su4aTP5RBpQH07MaA3vCrI3OLPnlR4/GnlzegZJGmKKrTwrcMZXh5EW4WRh6HM6xS2LmuAGI
f12IdmM1275KREODDj09TrdFZDmUBYAo6piaLpVyQIcaB5fnd7WASgxJS5q5WlTMs7cBADY82gSS
J0BZgwf17JUMrIOlXyedtbipDOpER5/1pcM4KsOf2C2+rgq9vF1pjOliZscUOVZ+YMzbHsmjikSr
qB+8hHOaMZnVGmDeMH+y2C8kjGGZdwJNPIZ0TUEPu8NJY5E54Wj8FCCe/ltyU7OSCqAo6CztEuHw
en8IQGfB7DdpnGI4mT7O2tqkVE0s9d8HyL0cMM+axnUUzRAJFAbnzViKL6rWRBbyKPiH9aOK0ZSS
6yrV6QF9e1dmI72IpXTaiM9LRNTNfmQl90lvShDHk3ln67HLgUA3s8jV3YQvhipqkCQ3jDNLOXGE
6OWIdotSsP340VWx6t7CgxGnCV/5ucVRzxH0bsS2jQYCZBVeKMA/P7hZJkEs5gGPc4OBN7xvEWKN
0cPpgkYlbawPxyh+r4MIMifBwCH0mLENjVVic/z5cHYJskqM47junXPYF01flJLDSLTaqTpeWHQM
1RRGd5QL8wRTRRFUIAGHb01DT2+Y1xU2MZFyWtcbssS9tTQ/b6PUJXdH5aXNJtrZOQdvUSonG7fQ
ZWni6XhX8QL4nsH8okIsPW8IZZ6CPho/iNdXxWxU/o/xpCTvrU05qR9rBAV5pRL8+Y3p8ULbdNek
pGfS+HLkLPTHv7nbOAhD6QxnPSymWIY67Atqcs8mlIXgoVOSel1/Nx9yGfWP4Y21NGKYEQFluG/f
0Zn/ZtkPtlnPAQyGsqorgzCnuTIcyBoVSGUHo71CgA0H7oxk+ebdIUZWklViXbT28KqOMngc6aKr
JounjVD5NdUxwgAp66yz5RVV2XZMkRaplLsOLbGR5ztyA8jGHbYq56803lCWJ1/rbSpNnfOxpJck
DywYn9+Mev9IN5oTBK8lD8WEWDNAuDaiHuvnrtRZnGV2lbq+zwzSIvxRQ11zmXwKPoppvkLbZeFW
OfNr9gOU/aVTmHd9IDsqr4xYQ8ETuNqcj8LAblDt+aig4uiPMrzdYsyPQgAJzzbE1PViyDVY04cE
mBveNd8Dlq3N6SDACSHV4Rm382NCIg4IsNZrcYQRg5JXvuUCZbJkOn1mgvYWSuLkBp8XJcMSDLA9
VWDC2XAvDtrT6wdqIO+uvvL4fkv4uN0D1VQk3Tl0gJB0F8OJGJwC7IqZvAA/qb9VOx6cAsEvf3x1
T3kM5PvbOgrRnQnHtjezpSknq/UcLdVl0fq59Dcu04ISg5kWKJcKkw0vXfuu2fLtvT6W4SQ55n8i
/q2IXzGNjoXuvY1OD0auKoygTj0vBSIMlvK6WNyeIC6F02sQ+sTf+suGc8vK53jAygBgOn0BTWUa
GmujdqriOwibgLQuV9osRLuS0JlliVNMcevKFXFo7UnztlrrV9FOXy8JWLxemDN6jV2r1xFugzZj
Ye3R4FmLgFVSiKi7/HLqgktVL10MelogSBY7YT4B/DXsmpPosj4anUtMHLrzC2xdHmxuT9cGJdUW
TfyQPwen3+hvXrHimtUldtA94aXwE4+IYH8VbS2KvYv1SxJDHYWkybSgJusU1UIYS1TfHRx7Anub
0yiuBZxz7G57fNRraGekTt4L6OquWzk/0nLz0gPCgfmKzH9sRP0gQJNFuoaPHdEQvc5Wxf2XZuOu
MUXRLRkTvQfuyPnWVAlkt1Wk34dFdNP+Ekxh884qVBD1y2yFNzcgIeQca6yiS0Kzbz9LDjd0MKUU
0B0mq/Q+vvqRCb1nngsSkx6yJumIGgzySasp290H8h5ujYCw/tjxB8+H2xh0wVHakdw+OrxCPlVl
Krey2D1lsbpzgtsydd4aDjMYhwpKD1X8oxOzAdxIGYPj0jC02Zd4dU1cjFdhoNmxm5/OBm293feV
/ilesWzDeea8pO5bplgeveCBqAnwJfXGNyIGoCUuTyi23GJ/BtofS+z9KuNQNZ0tdn3Qr5nDo8AL
xD2rIw2Cpy8gNTh9Erhywc6EbFH6L9PGLkgwtlN3tr07seCymcroBRmXnLTnFyXE/aVCOaFjT8B+
30+TarfWhf7aUiqQbIfb34pwTsLqDW4/kKbDCFSGD8QhHSOSR3cd4obNYgtUlih0udSwjOjhX9tf
3vTryAsucU8eLLT5Wd/F/nwt9McwIzPXrRCC2q52MEFGv9czXu91Lecuj/JVdIor9Qa9yAskEOZA
Jii+3LYKd5IYPAwyaGGMB+jHEL10wFaeEn+XYnKiNwAQmsNY3YkiEfXD8H9K1FKqvvAAbIjajrEp
+cwmf7MjQX7IaXzPEMgf8yzKoIn9A3fT4zbtwWQWnJBeZdv57Nwi6DM5wm1p+l3fDB8xq16V69XH
sJZS3GQ77ibZ1k+3tJGVXIFekIdMfBPIL9kNXHLYVDToRUIgxnzWUD01TH8WCs7kmtOGwDrTulC0
gyybxvPELlM2yDw8In9sbNd26Fb/IxIZgX6CbV72670VfgChliCccoCqXv6UmK4SNLgQ22BvhjBs
r7QSB7W//zMMlHy8oJLT6Dk0HgxzoaHnjFleVqf1jR1RM8Z2JJapJA9WiaPwhl5YLNKIEmpzonKY
vkTGFAfz3LY7gzmYByduFFBziurDGxiw7D/TJrK/dh7LYezMz0mASbvLRpiN/JhJfNnN72QYqjkP
pdUYWPzUsmQdDoH9dESnkKHUhVRtM26fxhzNiyZi/Fam597Hs7Mpi2nEKDglE2OW9tk9VDR+bJCa
+fPbLaZxhCw6mJU4YdKxenvkHEn5sVqyghA0l714t+FnMmkgVYzap3L36kVxs6LyJy4fd8JnI1yG
m3vlfau5W7HN1T3jWsReBq+WIdbfu3xEDw5zqisyBa9axH3xlwdzZUwsRZORqfcStRDgDN2B4dWC
99ca3MLzSoBCkfKtEESAVFBu4z4CZTkxoo0I84t/4d2fj+9XJWtQ5muZy/PUXCYP4VAvnNw10M9l
tbkCgqxJcFcV+b48XMTTOTCFeDrPhQLHj0hObjG/7lWjVfYvLiH+MPS0BG/6V7H7ow+wOLKQjgqE
GxBNI2xOr7Yz+54yLdQ4fFXCFdooTdiFXyx6n48rk3P95T/WRO0hoyLzNBoXPxTNuqjdmtwoJPb4
j5rBYSOylrldvGLr7tiVYkLQOZjAZ6ope3iIHJCQyoE5+KIOKCH8XMLVcDUSaPIVs8KP/IK0/41e
BPEmqbCUm0VK6jtGnxDjkjD+7XLBggMYlAqO41UkfNxZLIyjPm3iLQ3px90/4bP+NqShXpaidWb2
j6tTakeTLkGbuEajXXZFNaX1Jwu+LznuJUS5DLSjEJGOqNE+Hb42eSg/6kGYUiHBO9l+qd1hw6qx
6lr4bfOPYvPNHe6qDlIulLHimYsf5anszO+XwCrsOr4hz1DYM3wOdiEWBuDU8wb9i2opKchztN/z
hh0jeBkbM955LHsIX3H7L4tFRE1+q+37VtNwIvasqooFu+fzKV484xgTt0ZejXnCRGTrNA6LCheI
cL4TdaVBmNdxWMz0xLgG4xCWtKs1bd1OX25H+rRF4Fzw6rXj9+AEqK6M5uey4nAABg2GkN1sasJS
Ub6/Q5VwyhNuS85wQzGSyGTSgOktZEZVCV/ooewFVGhL7FvG+PQkfeqGpcXN8e2OE2rT30dFblEI
E+OXUkZYKbANHKbs1Cycpxh37TLMBFYQ1cpQzpkM77WZ/v63TRnhnsu1gAMnMSpU4j+Dor6l3irG
MMIgcITrSvxeL6ghWrhcnL/lA2elyrRZA+Nzbqs8i1lgL8C5WA7IwmS5WPpeoNKaH2is/JSUE9cO
2fw8hCx1q1W3WVfgg6eIptP7FkoIDxY5OGTQCQrPS0CD6bOkifEUdJmib+BFAN3ZqG2J0mEPpg80
9Eb6BmOQCPAJuIrogm7CwRMxulYZKVl6kkIpl1w/59gOneTZCNYdgcuyk1elbkRyADvAkBVM0Un+
21+eyhRPJ68Zc5T0steTkdF10hzvCKM8mx3toMvwm6r3sX3xafuA/TxIOwQhUkVfZc5BGRHsZDfx
UWWQlFSwGi1POJ+nqk/wAOjJATNC7IpF99hW87UaBhrTN7Q8zczToYHzecSKGBZmUY/RsTsfNAJu
6pUq8vAypoQj5NDLOkT0yA2JIN1PZVfma2Lr6NQh5qY2SNUE/JdN2/odgCDzbr+4CjzjoJ/Al+9x
k0to8mH8wTY75WxpdbHmy4MSobMygaUlu+duvGH7wOInmzx/ACaj88Z80rkqrwYeYChBSgnEvfxW
iE1EzpfskIxn6s2xgspEQRPnh54Byr+uQdxaWILIbuOBrEGJgC8/SkD6PsbiU4iA5gfmmm6mjrsl
HsN2rRT809vxF9RzImi0RrWvX+RGEYEFyS96MGuczv9d5IereDudiV0LJoR8Qp5BLrNLs3Zj6okp
10hiPfHI+QjH46N+7pKrbm55ry7DOvcm8eDEMRF3NtLRRIoxuL/cAKHMEW4TzI07r8/YN321N+nC
SG8OakPfC+j7dsNU5ev876rKOS8EjS3IaztPCCf8i4bD7et1c/uvpVzvxGNdQQ8uk8BKWRGoqB9t
oU+oVPbzluKxmKNpTMYbtF0MWlvlbBnxkThl4TOIIHaJR1sLz9te1JwMCTlSbwd7MdetW0gAUYnd
Iifr2+ZlSGzwF5gv2wpkRl8wXGDZLwlx4qv2EyctgX2yhVg/UtUV3gPVNWCNancPZK+SoNnxlYdn
gDqi/HBRhO/zvGP3QBesTSUCi30Ho5dd79faqU/ezFjZXrIa6apDAPCs4tuTmKEazIhK4h9mFqvV
lOhFMhu+KNCTwUwShskfj+RB7keJab4+XfQQRBh708W4GNlxZhQ8NImw4VPnQmYKxw2Fkn9maAwM
69T4Sq2ARq85VBAmmtYCHxnrVDCNdysFNXnxPej8BWBIuq5BgYgk7d8tscFMVQ/krJysK6nSvuCI
t3lgP+pIdrGIN3Gzny6nlHlCvxHLfSMXRn68HHWQ+i+XWWmdT9mNmOB2Tr96EjRYPTRRXJ+02bKs
IzS3VZRqGqWk5jOF3pDj+6f8A5psTU9++8Dwv8v2D//wsjrcAp7zU1kEF07rYiMqfTT1grTg6JjO
Yq+wxKGOuE6EtxYy1YgClySc0Um+P12i/WExv5YqIAjt7QU0lcDYjlz4y1KUhE56cKmxJyNaKmqi
/N5VWEDbs3jK161mmlCNm8YoIJlLWH4UuAoYb1fBsBJw53g6a0Wr3TL4JV9qlcIpfG09SWpUM2Vz
4HFn82Mql7XoLRDypBJxmZYMvyA53OT5z6UtuzdM9HtilxD3MVMN0G3H1D+3iZX/VdL/uHVWqTTE
41QXJM5/ngixOqFHpjmeN4sKbnlwzABJ0Eyw84FzB9gwaXilzwuCkOAaMvmOJWfyb+9UhbyvpwVS
nyYbORUIjlTYCP9Nn6xgQmOWBLN3du7MZlM8m6g0zaHozuZlek/bffj5/qjLBCijWJeYKAwILq7s
srWwxdNQLLuLgS08K2sYIwmefnwtzNL+CUQ+Xek0dQcv/hSq5VMjyvLCTAQ1jElCmbkrmf0pqyAC
P6hbawvi8WgZdZ605+Q06T4X///wzmUK2O/5sSrF4Thtot6cHabSjAOEHL5TiV1qNiZ3luDKv9oR
f/vRKnvibZsEis9dYlN5UDZbIxZbgCsRhsAnshmfQbB4MzPo3esvwAOk9yO+XsDXGzqTwcNmw5lF
slHVK/u00PzRGGD27oNHU1DiakXni/Bkm7E5HdfRPhS16jSmoTaOr2Ewr5g0opCC8eOUVpWkqFQ3
pTnbQoZLmdFwF6TELWB7QgDTb0coPTvnjWBJrGH+CmqeEJT7VEIweZ4b1Vx//xgu2S4vjwD7E97h
H63nHi/+MFz0vxhl+QAOz1jqlug8gOmHoGiiZ8ldlcRXs6JZ7hZbT+vIutDfY31+Ry0C5ousU8kb
XvQT6/2k5+AfO74x787EaDibydjbZ5vWI/afQgBZTs3kUtfgNVSiXjUHRcT0ZJdtNYw8uy5s8KS4
luEdpEFLiBGs6+ApTkIme9kUFCYP3612myi4fnbVCV6AOvGhyWNbVqErk7VxjeCCXCSN9nl35GOR
z5eoJgYFAkJdub2vIhCPKe8ZpGzR805HJBIw+bu1VtTf05tWweY2vKjfZkbi0bnNvqT721uYI+I3
u0KdJloajAMEaAFTxejrLi0ymeLtrBIRkC7prj0kT7VlCa9cLGODxEksEzZELT9JXT8vtstuHAtR
2ryD9Htu2swVhA1ZckAfJdfQMl0rAt6+hXmkiMtmyaadCMCGYX/DPr0biB+whi7g3w5AkYY03Uwr
58A3g3Q8JxJ1Czs0cU7ywVJRUV8FTmU9Wp+jM0PPsnNkMgJOO2+GtgE1brUyVjmQiScUoZKFrLTn
xTxVjDL0+1pG0au07J1wGrZt7NdHCKGYxrQ5O9dF1K6OyWg+uZoglFH8diKyRdzMnSpWxKR/aJaK
wBCf4ZQ2fEDUdIGzHy/unawPtrHxNdOclfWP5tkS9OeegydVWREQceiNrae/tQKICrREjIhHFUc9
QzpRWOxK7+pQZIQ/eHfr0V5LmU/3sz2nN7mX0WYVv8R2INC9jzSM0KR6z8eSH8rmkeE1IZyRoAxo
E2OboTkChlPvA5CPoOFaPF+dl5wDb0P1X9IbDZLb4T5RZlgwCIlQxQjL/sgC0Cq71pgZbDSyqGWr
cHxFDujr5MgsFlipXce/3LlFVQ+GagLdpIl8GDney3J9TlrML7L8NStXNpkUTLcINuciGPBcft1L
FisE9fVxJjzG1Cv0UWs+p2OyyQNGfQgJjcMzDG+J7U51Bq3OjDnEplD/4NSrJn5LAAK8MurqHWot
Yr1CQyblpG+703l/sSanflXVSoN4UdEpWCCBX4cxLBdlMtgONjPQE1/mi0xRcZhs7PhuvzczQYh6
uFTLlK97KBNBGrC/zsE5tk6KGTUfkEuzrKVi7b7FuBEu61JbJRAszAL1P90fo2Jh9eR4kW3HIOW0
jMYg1dwKfSM/BbrMYPhIlSjVAhLqCgESlLc6GGuRR0aJl2MYPR5gbb/qP51JlyrV9VbilAjqoFAv
BFc/Okfalo+Bxev7wb+pU5ApHuuGEloaFy6U0V/TQQ+wyuqjGtV+oAKyIECLII5bQrCUJ2DX5Vke
ofdOiqJPHMgGsbexzTO84dHk+HBYgPWspjA6MRhZrsBcUHyu0ktYFOgFv9wY8mk6CGOzPfkXtvcp
h6GGrB052nvVNiMRv8ZBbYr6QQVo/af7RKsSOCg6Awcf3HSpoaFZSG3YS/dDFtVX4hCeAgG6EBiM
H4DA2F7Y1L0abzlOSeInnyd2CKvPbY0gE5ZElvu5Rdk7ie3VrzYyjQ++OAi99bXzdPq9wIUBdeuQ
/ORW+UImPi8Jyaq08ReZ0F+6L/rQ1PctKsT5dBGqKbBuGCHNIITTPypavDmf8ybhsIu28nyufROK
plV6wucMCxfg3aEDtb92Eouq5b8nYuPj/Q/w2iVbA2zQh8MStSfLtzNe/FV+/ouy5rnGw+zw7dHV
2Ledqbrs53SO/zBXWf/jypW1hYpEx/efmbLmrHXrWCPI3abSyV9njViYGCMmuI8BzpoVmODWh+a7
5qaVKDeBLeN/gNMjC7e+VIIlHYZNKGONna4taWZ1iAsbEwQWrhWlY4p019gpQEtemMpk/MSIpabk
LfBLaWKCtCtdZmyDCBELXunVNI2zi1YgqCnEQU0N5q0nHx2/QDrxxIG3DkLxudRaKsXm/kaBptIc
CJ/U1P4ZhuEAv5sAtWWcyxN4uJzcx6kXv1YhGKQqIg4o29PQ43ZkmVlt1LMKBHCj3xnwujnS5UIk
TBOeTrrEYrLbUszBgq8plnS5mR+10FWUNCTpKRNEcrvtNDcPW5s6PaIcjefJfL/rlql7u6cGmjDG
RMeY5zY2LQmOP0gv8yAm1y45prpDr7v6u5Ro7CMdB1EZadtmVKo6Pm+tTUa8zF+Lb+0eM5wbdBn4
WbWA/oodrW8IP9ioIDPBCy75tWv56D0ZQoSBubCH8uzn/EXz6ldzu+6TRMMZR9xqIg78SieV/kkn
B8jEyimw98UX+469tGxqgj/31idX6OgNQ3GucofgK+rsz0eOfSE3SJAUImHQNtZrU4eOFlrIJgGa
iOyJ3HoLRniB2vBDj7U2b0bbwIdaUXI38gfGuJcHiSB63JyKVtb0BGUxp3U++hf0ayjiDPCR4KoJ
DEkqXMrGUKXhdluDNj04cfVacdaEAO0xOkfI/R6cNyT8+Yvuup08lCpBRR0Jyg65dZ8VhDVWXT40
QoMWuF6MFwv32ssaI5ys1tcwUiTaEH/2hANknOxYIl1OOEht3AuEQ9ThpsN554Muuju0k07tCrNi
alYzn9wRysEdLWIDNZbmp4B4oCjr48ex1X86yqz2TpyRHjTwZ1D1H+AGmQjL6UPI07SgLbONlG8I
CKL9znsm4fYAioGYFmbksJSeMTFq53vZtvqcrAxVDzb/ZKLSTlHxDbI40RNHhNHPM/MwOjmB2X6L
JUhhQv7Qix8Ax1lmy5YGwlXT4YlGdP7VZnoGZBsBoKIqKE4kl1+QYJpCEBadmm7JPreCeRDoz7cb
i/SVhTKFv6C+kItyvTSLS4hXooizBmlGjOo1o4b6f/kkcQ9Hs1rd5vC2ksZ3bakB3F5sk3DOb+JM
L7xcUCqEEQN1e8bONitcd4v+NiR8n9+HY1iAiSasDQVrTIkP6cJ1UZh/JZGzAQK+5vo52Oya46Wq
uRPJ9nLzTixjWTe71DUn3mZ98q6+HInIM/UHbjZAN2+JLoJeijDCiyP7GL+aZpb5yKKPd8gwHpVq
45jaGkCmvV1dIRLlp7tSazgKjEjFmGaQTcTaVAju+iOF3HhNYAFqcK/5UKlEenAg5cnqZCJ3OFgb
3oznv24o282pVgS17250iv3/cx8IWzJulOSvkPdEFPzWcUn9ekbQch4EAInafzscVHP91GLA3h8t
vFDXDNXAbvglZf3j8GnN1+mn4OZwt/btm+m5H4IIzRPPvmL5NgF1wBdyuw2Nd2tx3JdY+gTr1a5o
lIkTWUo8jZzcQo1K4ovCWJh0jszcfMETrr74mUidWugwbaXpFvRzLMM0a71Uou4iivkudZBiYf5Q
VfIQ6t/yXjjDuCCkjCuJ6JUIQb0DBOmo21FIDzuQd9cmn+YbB2Rv8rEIi+L1kboTXqg0clECa0+r
nAsIbmOAKwG4Ixi8Gml/CZBx9YaJyXDmtjzFOlR67D2Hzs1TZ5MFXMC2dsoNlX0BkiG96c6VqNho
eBoM3+75PD+VWCGkxLmZZWBaFkZGJ89Ajdtj9D6KbzN1VwWImWQEJravjswz++3qq+0dkIWwqmn0
H5LLXBxdWiQocICpHvFPUsvw0xz+7BGZ8hbbby6SuAyfigCVbNAnAo73vM6CyXItSG3ee6u46Hk5
DtgzBNjzes1ddKDMhpbbaUAs6ofR7K4VRaNUjR2j+d4z6RaRNVPc27zu2OB7Ql/9gWlzOLfQQcfn
DmnQw7kqHDaC664FyG3kEvTm+QIfpTGW+N+cltpt/EyoJzduh0dkUE7tGxDwx2wNpSg1rLVShGIs
NBJhjNQy+PPXrfK0xeE7maHs2A6FVKYzFiIyDz+GiwMB9PYmQuTN4FB7ojMs2GaWOUdfEUV1qf6d
vmYuqp0yCrtJ8/ehqqEyHD2kZ4sj542kTjemQsn+rLkw6fFlt0bNvxnxELRFij42HJqK1Ec7Nd8e
O3XN7HMg+yIGJJuHkmkEqS/70JmrQBqrremYJuOOUJF8878zJ4nQZhFhglG6NlK76/DrveIm9dX8
Q16k85bNhSbivYnyWajZoeI7jrgfrv7T7vKuy2vVEecs88IRzxtZV5lfjGx8ca0EQMBVO0+veeRZ
905fZUZSoDqSz/miklr0MuzIwnCT6QhWZZ2r3wYDye7lgtsAbbR2n6HRsICP2NhnnMG4qARM7CBY
E1kVAgTuhbSI6cJ561TYXktKCW8+xWQHHodBj18ZYmovx+P/g2BOTjtuUI2whK1TROXG41/ytGp3
BkV8a7tGcrRV9ZSw7Bb6GL9MuYik+1q+CtmUN7ctBrawyGkV2BMLhjYrfr7ibmFiB1J4bJbHDESP
vgZoEi0N+1rYz5jvTTGRBs1G8tZE41CbF5KoeGZNLA+i1I2oDYOpJO2PL6V0SWYndj77ttJmZE9N
0yaUBHziWMSED7Xmla37TOjzw7NFeZRsvS5f/PwPb1IrQncTSKYsvjeZWkzuwbhWlflgfhkTAmtl
AF4RkDNgcLeIhJ9HTUpUQnB6FWaqziWIokXk6iC/n0BuyzTMs6dsykhYpiPDpv37xyiZkCSAq/ez
yp4hBnl20pOW+nfnJ1++28DkXD9tAAUcdFynKNSFoXp68pdV0oeGKe8wQr0f8x4zh3LoWojstgCV
jhw4vplhO4LzPtY87/eQGQ7umow4G9WM7bksNyKfZR1NHyvbO3ke7qeh3PVmLCWw2awG4pT59XVw
bx3VbMv50hdS1U1jqj5JR1B/uukgmSRf1M0Oz1SJsl7iD+9pK50amkHZzC5B6j8HTGh7XkTLcD7m
w3RmsqhurAAkVPiJMEU72Y2V1NOEcfB7H7TxBP7b4GhZU37eadGZwJ+YjkAapZyacG1CCGESH7B4
jb7mr+/17RdP/VfIY3W9ebzEVO7/gG7PfGkYVMp6EbUDZ8txWTsj8iSoNU5a72ER+u8PgoEVhcI3
/8y1lJt+VGF1ugc8EsaviqeD/6LZk8Ive87oDFAZ3lSlC8k9ud9lwWcjCq6FEz43nnH0IkXwm/Sr
7B8xzf3bw/b1j/DjOUmp8KcX5ErAjgs6zNjD2jKI9oRMU9eHMPC59SB42moibJB5nCc6/QSO3qa6
VCF/+FB4BM62FIr/BxGxWS8VjupSZz9yY1Li7BOSgQHbtooOA9gEmWGClpVUluLyOPpx5bT4D/uZ
dujbO7cRDgiGoWxZzx7eMyvg4LfHpd0gMmsRjUfKuJb1icIFve6daeap5Rbyhp1cr8G+XA+NgQC4
xa95nLTECiasolYlbbytMhrQs7Ewdb3DYfgg3jSrB2XdNXKf7sGo00GV0z3pSZcgsheyjJ6H7DPu
wktfYOJV/1o7jj5KNFwW8AAFDh7AjJ1PGeDjRbONnMNBzuvt83dg+xnPQ5mzhZfVQlDY+0+KhoMo
1BPMhm+KSCvoJy1dv5SE0ErWBiv4NuM6zh0UsGDcDuBP4Lz//Y8YcziZLfNn702XO/Deb+ZwApwQ
YAy35qvorAJ6WNBxnZZdcVm8qAgH2mSF0MqqxF/Lc8v07NAs/85ODsien3jMy0N3sOrD+O9UKX4p
MEelOfWZHtYD9cshAMq4RZhqAIA2L+ofKWQJKdXsIV56VtfbNW85sCxKSDIPTFx3tSnsL9I9tI2E
tN4R7MXOn7BPkceyQynWrzLYX4uMcbdoo0Oi0y2L3hY540wi6MXiGp5HtC7Mj/XAgNyuhr05n7D9
9CWQm6bXfdS08JbQ8W/H65h5QRjf/3nMqCkQGXGDv8Q3jFZk2obLL61Bjq4ImHPJKP0VoJ4jbUYW
VNGfrnY8nnD/sE7NJJnNnGgYjHftqQT5B2H1r/nrucPG6iF9uzRF+MT7kG2oY//86MKqRUxFUaIX
KINirmokRL0z3JiRuZXqdswHp4NYMHBfdvILAvAl4Gg7L+x9Hh5o5uzKcxVI+XSc5vBf2nLG9i62
oXyc3l3uG+N1AQdWQhQMWD9MLUsQjmitE/u6ukhx43ok/oCGbXu8AJxjk6M9iob/UBOJM7ClbTqq
ZXKVURsWs9tuld/7RfHIL2AT+1m556ABv+XC7VXJle/dfbqi4df5t6ZoBc2T7firjpsgjULb4pKJ
xgK4isebf4AOTZz56yaD35u5v7oPMvV6I715ov/eSct9ZjmkyiK1HLiEu9QlRuyg/vcIeY056T0W
apeLimaMa+h8KJbhWTxkFdlqCEOUaAoeRe+3pVivLDsPA00K/cjEGghY2CrC0hoj/YPugk5SCHLG
PaWx6A4oxwX8mAseJs4LWcHyGW0nDWpZQmkw4b7YHCq5xRQiA653f6HLOQLTvgQi0k3Z354H7S6Y
kdK9Vw5pTcNj9DIWklYcxyKNIniSjgHaaiQpkcXdF0kv04mLL1tMspG7+QkIl8W9AK7cer5/8dnW
iM4/I+fOGl0eROOpDdDpFQxBSeeVQDQRK6Za3IHQ/Jd9jrXQkoDnRzXBkMUeK+9giVPWzAJ+IcNi
Uafxn6YY0soU09BatR/bzJfgnL+wArFP5oexN1WMorbzFkocwb+NFXyh8/wjX6K31fDgvhDLfuf3
yLjAzT/Ps+A+q287KTpEMOVawR7cLNTSBDjLjl9otDgTzrQSya6d7VGRh9N/57QDIjw9gkAkSwFe
BGYm69GYrGkMITjrBHiXI1BktQhasA8DdjYHsM80pAbK3PJvMBjNgfnlA7Pd1CKE9KBuzttwhLua
ZZgrvOPjoES7WDLczjSkgeJ/e0aMzgtjRH/0vc4gA/KCjfWDqDnra2fVIEP2XGuQfW8Oyfc9DyCU
dXb1E1MhHOcGFOO2+Sm0au5weE8I5q5EZWiEeNKipbcY3ymvA4dhmF9q1eDf/b2HnUtrc9TxXXVA
OMCK1+y35mCNDycgXeEmYaIkN4M2SDiBh6BiF8SuKxYl87ZchVWLxH3RKKRqRR7H0MTYgdt6jAvw
lsyPqhQcBut8dDOqqLU0ZmMF2gYJJ07zzEl6paQz4ewE02qzMqMKXbYQxitISEvyHAhJC3Fxftp8
tH9Ip2IbHa6QVa9WasFSG0+8qkvo5lBK0uwxfYClpD7rtaVctkQacLdmB6cNAZNKNu6I9Dlt+cYv
Kij+08/hk+tbNeylZIWnG6KsdxOg5CwEcOeXgi0PUJ9cHER2eyhd+v+W+ehxvrh3fFTh3Ln9+ZeK
7+xJsFoGCQ9wBlpq+PNAPdDbZzHiS8EWrmLEUluAdwPiY27tfoVsfv47VkjKrQV2W8lZUoa0i+HJ
hALx4/NH8/mB81R87vm2Z57WooMiEIg1tHz14TVJNyWcPeoYYoMfTKmT7sf1n8kA6cwIO1oax6WY
c2vpSS7geq6sNLN/PfujeQbgnq4cmWwqlhyn8zJcnUt1VsWjtEeOmISQ7UiWF+qVjzqRb5GTyJbx
8nb7O4nRWrhI8O4qRHyBuwhuFAKwldFIp5aA7HUlEwPrXQuucB0aw8y8sCMo9CJ+ZKsyOCAyLGCD
6aKJKpblZuTEbR44A0/1l6OezYAXxRuq6hTK9fg7qWu1zbxjEcLJeuVJbaH+EPSmWgot748dSUIr
iLhyadus6Zlv96I5AhmQEfSfOkXwJUbtXhzYfQ7YZ1uAFHf+qzCZBu68Wk0VFQ26ZhjFfwD8hOPW
K557O31Z/cHB9UKgbkqQnWFrNudEiX5xRVrjy7wDuyuKHOCgqG7TWx28J1ZYCs4rh+n0XpTjxFB0
HJeR12GzKy/N8TXUlFdFunKzeJFdGmJbB3YWkt8NVHisw8qv9nOy9Xa2jdhwXgc2JFkxJU7JVOfv
3UqBCTZxQ5tvGZTA0Z/p35/yXZ/ia6g19sG79ArlVefLFpWwZKnnRJhygun7vREuiSHnZ6JQTK04
Qxgy1LkHMJjqjHJuCbxEhMsM7WwOj7q8mB2vCiqOUdCRBO7MBMYT1GnC/TYgp6fRcKe9HFIEPHd4
TDyqc0wZLdcRzk+oRDr3eOm1/A7GF+iWMWZXMdpEJLpqTn5pTfyyr2/p5TNCNXcMd9qAQW/Ojca2
jHue+qQn7UtnnWoVXTW8oQC1R3jFJVZ2rI0UWkoLBHWmjEsM7mfz9AelHjJL76h76+C4BXFD8i/J
lXgubdmGviP57KaTQp/ShcS4IietXWs80asq+lf4ipWo7M+mKhcndy2ERAMjf955ORbN1t4lEQHs
b7slqupWfH3m7WMfy2ApohwBPnX7IJ/nKxKTPA1W0vrnOlup53znFZ1xJrYWKMOeSG1JB1mBVTaP
5zTNdLwblx0CUtOmOKM2v61HSnZ7WUfD0BVRMCH+pXdyhf3xYJaMWmFk4OF2EU4UILqm7aLVvl0a
oB7xF6teytx4vFYK3E8DE+E9hq676YEiTVr5cJlWSEX1VHnvDDUHU16CfyVse+QCH3CzN4v+8yXn
DK+C+PtKTQxuxQf2L+4mv/jweBmM9KlNOrR94AuzaSrikrCkzBEp3gveOG1/n+4U60JMyUADbEbv
p2hhnDBM2mz2gaookvSqivMqxVd9il8PSesRTa27NN74D8QJXwLcP7hmxKPV6tpNrwAPs0ExBiab
Be63YQWMU7H7PGsOH/pslrMp52iXm4fzfSdZnwMXeEeTNiOJpZ8x+mr/yLOEWfuWitLDlO/iP8Xd
1AE1j13UBk2VejXawZBjaqjJaRp/nvQGfk6+H/FL6/XKJtI2098pGPfna8zaRhRSDl5vbokKxnpA
6sWuhaSI7jkZ8F+OO3T4ePPHh3gJDKCiTMyiaqVXOlmlxH47sne3PEpkt7Lp2pp3CgDfFPO1LVXs
7jSACyxvQiyLAlAuc1gF93ElCx6Pc9j5bwheP1icFeYIK1RBbUiYbctUO3BXTSBf3UpNSDA7fdK6
H840XkyVQ+76jyp4QJIs44sPE22/6SWxinl1VVk6DHhCBwm12zguZ7d+ADIopIselutjT+eRvKL8
9PNCJl9ifsZdF3KoheCJUHkgeW9GISXV85x0AR/cIFGTXoudlW0pwH5QAf1wfSXpcErAkUsS7Ekr
UCebJ3mtubiyjOCBGUokyu9/Zvy4gZWU7Pu2WVR9gJXiNJCoUXfl35bkPC36lRpGwrEbVEc2OBg6
5S21q1vXZbzsdVenJT83tl5nsqyrENMsO7lqVFUHBZf94u1BSkmE8ByREWnmR6YcuWhaL7JA2h9L
pnyDy1ocZrDtEPQXI+JEZnrq/S0rN7jUB/MV6G8uIH2KGAEOFyUooyx+2cZcMV173ShcztRR+y7j
lrdjI3tyK/q/NMulM5YtTmvJYy5pptMNFTzRfZG/1LXnkk6dztm3pcnYPGYWHE9w1VOBiwbTg1t7
nql1oQ+PtQin56mG+qGIMhmZMLZOXoC2odFu27vNXH7MoMWM8NKo+IZ1fS+KymXE0SqLGvrjVQmF
255BJ//ZP114X/5KP5SmmSPBbH5W9+3j2n+3MrnO355YXGZKnxFeafba2sJutMQx3wKEDaqP2rYE
1z6IVzMf3SqwI1w6RxkY2Mhe5ajcVc7DtYV8Lb3mJ3LGRgV67pBqQYIPW7vxHG/UY/eY7x6SLqix
3liAJ0wZLRNhWjx06/XOC4soGc+nPgBwZx106SCDTjHoww/weWWJKl11TsJG8ElCNwWu0fnns8PE
n7mtfSgX3y8KRHcEfLvfRJtX27R3L+JZsSL8XmXT5hjinCqA17InYbtRmJmvLe5+2WrS+qB3Tq4f
V1wHT/fnmlKFTqclMbbjMB6kz9rqeJUVWyW+4EFVV9Z3Gx8RvSsLyQ9FTiC17bPo16rGCaYZvXfr
qfDZjUcpsnHl0sNrnJBxrKxUq2RPSYSeV+q8yqNQBUl9rr44oS0V3cgKT+TMCKgkaxePROmb5sSo
vdbtJh0aEJwwwaRfaq4u0wNnnoeezYAOvl8Ha/Cd+KEyr1r7piKX79vMD6BgfCt/pCZ/V2Yy+z8/
LGKP9Wcvwmnpky2cgIH/XpUbDQR3CnLG1LeysX0JowYFlul5nztbrAnG1Zx/yoK5J6N2V1LGyZFZ
DIZ/9ZTmCVAkxDFH4HgGZYYfZZqgrErO/gmpaQpjweUFi6HV1qvl+1f5Cw5n+TBp4HgCpi4WlVQ8
qnExM+AQnKV2Lx6MsyU9gO73C32mgSF1YdTP5cC6HofxNx5JW5xcV0q4+r/WiHYN8GWUZUNpkp27
VFR6RI3eUKKecMrQCSTdFPnjwQA96vHOM30asnsZBZlJKdoEG5otG+h2FFAqgmFnnPXa8JX/GMW4
RwA0stqmOZYjR3+syM2V1qtJBUnVOue6ihszui0IpwArmYqK05ldEv08Dq6N83/Ya8M58v9dJ0Z+
+CE8TCEG4ajbquSt9T4zsLm4f1SIhRv+7O2pk8qdr2q+jvBRj9eYr5o9OH7uTiojotcLrky3VZ8i
z1dIrJSyPTFWfzVj+ZTDZjZPZ27VETCxuFt6rxFKQJAEO3V7a396I1GRC+DldqNbCbR6RBye0QrW
2ad+K9VIDfjqM0eQf6LN1VH/zcy8a5TS/q3ksZ9ijdxKHbc/rOnXJbOYoYkWYwV983ko75U3LG61
k0UsljrV0WuuJmLSFXGesRD2ueJkLRg3xgPPs/MikTuUrBtUhXf4ycWcjyWp6OcnSbVUFRLEOIlj
gjpGFHJhePghekWH3yQi7bfPQDBxMmib1CHW0OAfZNpYN4yUx0b9juR7OxedycXTJrohq3WyyFKb
Q6RRhd3OnSoo/2gGhzN24Q730cHKOq2Vezzps1a52XwV0VwrxZRw7hfNWAnEv1dnqsP+UEGmtA9x
0cBbL4uq7LIgQMSpO6HvTHAjmsYg8RhJ0XwAhQsv7sreK1hySKnU6mhpZdMU4+XUT4e+V7VyfqIx
cmvhDsEf5GUnVPDHcM9s6wEt5TPM8rBVg9TTs8r3Za/RXfSDOwYUAc5YTd8EPo7F5LAXHgQ0ava4
qOrG96VwF1HinNoEDqhdPftlXZtxuxjsFrXcuiY5lX9AAE86TKTxfY++OiZE8HTaDyRbpS2DcJs1
Ymmn2hzljapOpk2QnS6FCI7enqG5OzvE5Pdbtzg+EvTtKbcLjYW/gPuttY7JGYl7+kdUB8BKN/oT
SBnPuOET8kV87bdPxScOazfMoLK8H8so5RzlspLzE4hVNnpnS3VbGHwSjkwAj+5kazyr3LasCb/W
dNUKSj4o5RNProhZVuMpiIJGA15+FjaSUZZ7yTOHpV5TTlGwgNpK9HLDTfcfVJq3tXiVNowcbjsY
kkgSqfdJo7PxU8GqVvSuhptHgG54ADeGXjowdjaUMMlq0ael853Tki7rJxe5uwUtN3wTnUK46Hp9
35hgcgLzutAPr0XjmCi2GTfSYPd5zsCvDMRa6nvFrn8PMx6DJfyxeQ2K7XEM373LPo0nVzhUjukp
7FimDI40HUhyr0Uclf9+KbbEE7j+3MH3uQtKg+eQKqI7VG3KWtq0aH46masJHRmu/eZKQW5lVSbk
K6E+z4uHQdzVpFbE3FRQ4dM8A4ywhAiCSLAIby6c4iDSo5XpJGGK+lqfD1GrIFih0MSVyKIV3nm7
Kc/8h8fAkJMwPQ8/BK6rhiMTwnlLNdQ7zo0rtyay1S/Go2sPJ156NlRHGXMeJ2PjWGAB0D9lvYpL
OzFUFKZk/1QsLJUA/2TslVXAxbXAkaORP19Iwj2kB4dxoW5bXTZT0RQyI2i1fZH2LfxA8K9nNXHf
I+qk+e9ozu65q1o+vWrhz+daSxkXDOZakGlTk/GbuqZOQc2bn6otXRuHgbyaWUgopqNQLbZm+6RT
RLtos8r+SD6r0Y8sdpcZs2kpxomLJ93OXokdZoGFDJXNFuEu0PRMl7mPHGb4GC00YW5upleMie0x
AjmRCtAsD25paIuY17s/i06iPiL+M4iIE5nYX26JamWkJkTTWSL5wyAcRGRSwr2Mxw0Bgap4o9yp
4t0QvlaKM22tUqk8Q4zKyoUBrICH6M+fy/Zx7pZ0niOVz0XWL2Lk2jrLPOpKKptrAKtnBKxmfoZX
o05BcwSP7AsD323Dw0Gfb5JbtEP0Vl+qkr6ypUkVY0YlOGR9cpGLpqvQ7DKJEqrNmFiwT2aFirit
tGLEJoFq+SgcApwLkuxLc1QctK0UBa+7qLn2ysqBT+JY4qKQk5FXPL5QsInpG3owNCxB4DrqbjTT
bd17frhew/rj4cHRRwa96iwkklWNpBNOerR0Ylp+ZSxUBCkCNBMQq2kQYEytZdKh4BIFqx+lyJSV
Y5g3/hgRo4RPkKbqBT7ljAzD3RLz3c+tZnjWIcQjxxIiZmadzmSsJqBeLm8sAVId84SWIFdIlOrI
laV+STJCtRKGwoIaz1tfizgzOTjzvVTZXS9464pz20KrjBseVG5s+dcgKEveVvh0KyCKLva8Vcw6
DRclqgbZXbbV+XwsVP4ZtMK9DBBu3bXhFWSQn8ww7SXQzzzRP2PUQoFgeb0GQJJAGXTtQg8OKXQI
a9owp01PR0qA6KyzgdJSrirk0W6Rqkdc3jMhsibwJPo6OFGrHbMDz4bYITiaWQXm0H0wDrxNGL7S
8q+dFIGWqrHszm76IxLKxGyP8Af236EJ7nxEFLWm36X1GPAlYPod05Es2bIaRflnrmH5k0i/KwnZ
cfAAejYrL8vMeRBrpDWfpCxQ9OsBxbp+HaoW3bcGhOEk7gkbj6DVxhm51t+IiN0iGzdw4DcWFOYg
2WtwgSPPPlx58nLHcoqsXFJALn1//OU1jdyjZfeSd8GCiOCf2ChA3X9i+8EgPDiyOjAD86hE37TJ
umMZKsYtg1IVnNqKIt9hBCQnbIZKQrDZcexxFqjq37w09F/Hbuw2GCsn7q/A6a2GTM4x0gkWSIM6
y8Mi0HgytLoYm7hKCY0zlyCtyX+TDcJX5kShhen0CLvJPq76tyT67FsbSHnp8mslOMjBjbh4urow
ag+DkASkTBJvMiEYB78qLWY8b6+zKJwRDR0iIA7ssM16cZbd+ntJ4fsk3e1u7RrCqo4KjpghZoii
udcR4cOh+gXWrNLOMAlFFPcGJiQl7xeVoIgwWM9yteGhsDT7fQpQ5GD5K1XgYw0ilqv6OQxwiMi3
Q8m0CDyAI/7ASR2Ufd67bFZiO6CbPYET3yXxVWz3krJVzNDFjm/gAn3ErFnzROgZR7/E51y9W3+R
JmD0YHHLhpUbiWx5cyc+LIPOfP6aAH24d8H4oV1oNnhydahc3N92k5Yzs8rXvpJV3nsTxHoliPLy
aOThc2+wc7kLIkdpZ1j1pz/m0t/5LtM32F/NodFXDVOEcm1aG3yMNlIHMuXUFn2mwQNWS3Zv9TKX
CpjSSHF+4eeYSBf54scbzYm5Npe3eLuVHG3X3rufM6b+UWESzrr1aV/ZQm2MEGMEvpHMzi2n0uKQ
BVQ46AZldUNQh7C66CjJUjtKmLtNnOaSGvfFFLJ+jK28E7VAEP6vjJtCuP7PcXSdsinUb7xW62gi
9UadHtJJmILtF3b30htqx4cgYJzMuOBwhDBYTfDveQBYyJ6EvtWggg3Vu3ys7XdRkoGPaRm0UwDd
FGfoYx2D2CehtmmK3pIpN2aVqE39EjGUZ/c4YocOaYAiXPDBr+ilk8Hei5mOXj0Lt74Fo2Y88Cv9
dj8w7OZU/IW6LMBhVs/7cNDiG++9sa8hxhA9VKwL7BRB2PHpwF85UtS3HZxUTLBzL/lsx/IN9mWP
H/aUBdtfISgtBrxHU2pWc3n/+vdJtO4ciapwlxXlTYpmKcklMrwhl/fCZ3cFHhNd5g2d/6cZTWV/
NEfk1nX6uKeuBazfPTYE15jre/+onDdDa7TExE9pLnoqu/5gJUI5InES8Z4hHVtOF8a8/oPHcuuW
dsX/x7nud2lL6ULJyZp4/eLO5e7/ykHGturwcgoy8eBIWxYkNegw6VZGOA/X9T3+mkZNPtnNj5nF
KzKcLESTaxeduzBLs+b6ktUkTsDxrv6M8sL6NimlTyVbqssO51v0wJ1vmdbEULzzpTgp+g56th93
temHm0MHvdYpCwLh5oYZbcJRk/4zuXotVv9K2pso6EIed1Cc+14TOXBtlRRJTq1O9i48uc7fP0Xh
1mnpyGm77afSn/LcCtX15+stLMJk87PJ7ukA4oVXV2T5DCVMsHvEdKWsTGOHdg0q9mvsb3dvslDq
Zo9gy+Q4K7XDTiM+5QG2nKosOQQnF4WckUeywv/vQb7L1r52lruQ0DPH94qMYLYWkHVs5z7XxZD6
xcelSpJQTtSO/7BWGs9gUng0IFeoEFKFS3s/AU89ix/A9of73j/66EJq+DYGZib7OEloml2SNsqr
fmXdVVGG7bdSCZZ/uBj4YmlLcXG+FRUil24QJ3GIPl6CbrCu/iTnCyczpUFyA5oRkmHFb9UdIim+
swDeY7MZrNSz+7UF76f8kEmZwrR9Chdb9s09Ktds0G2OCf74vnkzjnD+JjQfv8x968XmlX3V9TEu
rfc0xK4Fz7mBh4hra2VAc55J60VkPvaTl0wm4lc4kcSn/17Hvnn9pIo3ZbWigAOUyA0RgjVQtbFv
1Eft19ro3eH0tp9iFSZ1DYlRzEJPsv1OofpVrWIs1vwVIQ7Tlil2HkTV6+X0skqlfARlAnWQ4/2M
r7iIXp96W80IcknKMlTPbJyyJfwUe8QNsmPxMvqtTH67CHr9lTTOzUInuCK4XSL0hCIiX8H/N9jy
LAA96mfjeCRKFlQZh0hZNfPklF4cQG4TF0ZL1P0d7ARDbGmpCfi8he/qTMQuSm14c6M8UZxWIfTk
ujHTpKZToi5gHMYFWKC32EN2j3My/lKVncJdxbD+cFfahPNDvr4t/KrNSe9KSVd1Xuyl9cYLM2G2
TILiZXHYXL7uWJtKNxFqRRERr7oquVWAuW0DWZYxe5B0k7NxtFdo0jF+Avf3ok/08grZ8eguwUN4
QNEQORVmz0+WxBhog/WDn9dHssxnzRbj6e+NJWSXPh/FAihIq9gZkkp0HgPrGLiYmges/+lZ8zxP
OZpjpjyIhSl1IGGbOxjaHjahRjiRQH4q5t+K/AqG8s6gqnBDk8os3d8KUZQEtGE1oUDyfwM0bnKw
FgifdZsGJPflpPpRCn9+13N/+tcLpvNAfPH5x6T2444wrIFZ+7reCfAxjmMVPZSjvLqD77iGAkNX
hJaGuz9vPmHhdKRZ6qMoItF+/G4QVTzxLCe2xn+CYczPrxcY+5grTtpf19IB4mZcLi28CTlNhRdz
WWmBg4F/oQO4IjoZ+UvxOB0b/QuvDQ7iLjSSvFFQFJgpYtOyIFT8HxLd78eyZDECoMYKxw6tJfj+
ouEyHngQfhPyYRKNsXOuoPz82VXrIdIV5Y4uSb9PJalWdOG5+poMYMhv/is1qt/46DfSojrUHAcs
BhlBHRxM5i2+7+Zai2xZ1+DFTNSQnQWuzE8r//iAhT3eeTaxKk3QwAtSRYEL1lPluXd+PTnkbNMU
/cBQgDjBI20i24Y2XA7xylAuybtYJso4wAsno3YQL1FHksqy/SIF7409RSmuqt9rllRsJO4OnJVv
5K9hf6TwALdEsiteTGebue7ttMVp6p7NvM3lu4d8un969vt9Fxr2sCclfJ8SJpt9ucn2inTf6wog
aFnqzQ97o2Llb5Y3vilI/GZ+ZiMYr5XgNFvwkRcVuoO+b6YI4V18g1G3j88ChbbZ3Pn0PX9MIV/8
iagdVHZBN39DhektbAkMkqENOeoQynadaXFQfeYMucDe7xp/UyNG8LEigP2ORk+7JToPP2RQClqT
E87zSCkkVyzWWbFCPdv/sikMITiUduiGVc0IuG34favyWaR5TEcehN2kvK0ouakrS/lwiyEgko//
u3tmSVzvsIhv30DDr6CONZoOdx1AS49uTxlQWmyfUPLVZxJIqLDetLXjxhLROXjSLrwG6Z3tM5bi
BLCmiz286+fd4nHS0idnIQXl8PZVqOYA5KyEh2hD9Kj76yXUozWVoBI4ymXaLivwhbXSvvxU4R7L
nWp3t9ifFH2cLhCUxIZxGS0Fd1aZyGgpz9su/ZNuWk9O2/+udlGRj8HEOEOSFSrZM31OCTwIl1Ue
EWqKHiMuONvxKzSyAsAvRcdNGkCPEGF/qrq9mdBaGvcg6jZByCxj/Wl0ZaiXkkIeMQgZsj55heau
1fvbllGQ9xnTnvi1non4muw/rppLw6ENQdQb6MkkotDIZyEM2Zq0MIL/VInFRrE3pOMFhK4YcRwh
X8UdxbYS+T31elkNRiRuQ/Mz9LgGt6yIesidcrXimfNcg2yJRXlSnDjJ+PVkK0dBJ71qQ24r7unr
XRipy6iXNlSwZ+pSvY9PqMgUHZQ3JDbMXQS1LgeqtoV3Wi8uN/rA57U7pN7GG7Ba3CcEJTVvSdzB
5IHeeE06wbYgxLocs92cY56N5JqiCsOP1GTP3xomuY5DKDO0bN//ZyiijGRE4LJGgIEYU8mNqIul
tpknF0Yvy1jTKQoA9P9rjK+ryhkjzvfXayCxVgc+9HqllIDjby27x8EaHBIr/0AwebglQYs9Voij
/pI6jXsopTxjovHDkQ/qKeH1rCPw66jNy3/TRw9wsesAfODM+E7glBDxVU0okvfs5JGgRbVaG+ad
UEVYgwuiMtGKN9QJaJ1SDfewG85vYxzFIXzWmVado+eIyXSu4O+MRsQYk5pND57rJJhgiAA3Kwbj
LGz9YfOuZF+0elEo2ChkfniwAXAq+nTHNTg66c4EjaY7ewnsKXikOaC9AH05j8+VLTbRzZPO3MhF
Vt0jX7ag/53zJ0kCaGnIIy8UW2wfVR1JehaTgx4B0Z+jft6rvVnMjB/qLzlZbIq7FnRUEYl4p9tg
3st5QDyGZ1F1zCZSKsqMnnTYNNCyI7q7Qgw2aIgG/0oIpQD98Dm5zGVTg9pisAul1Jx9385RU8oc
Nw4eYdxtixlkUfY2IHmemoTeRqm8/GqLiMkrlyd13IyiuFK/dg5ofsx6/ZtX9k44H/nd8i8LIwk3
4UxVPMk4m50mZWI2ibAJtnuHKrJmc9IHOpHkauvlXweJXPrPlCqu9u/pOySUEW34UhuJbypnJg/6
PvhG1Tt/z2KxAyOmXEb/kEXm4QcTuNXVRCJjDeDswxu0pweGu/swovsCCxYColnYswg8gPtg+6oT
GD1HMYBKBcOze4rCM3CRf1iftRyN09rqQERoUGqq3NYRSjgepmmSnCHEDobgws/bRXytE1+6J65I
vQO7btIX3BmXj2XP/cz7KgGBIG9jptjZBi7CcTSjyrv3LT11TeAXEvB9/ZoLjG0dsvtjA8+PAn6/
Uaut1/3w9I1ImntvPa1P/RwtPWWShRGXQX9qwjpEePtH41l43En3+znOSnIA/PV8UwCujOkzNMsY
SRobJSUS/s/vEiw5U49ILmF71Ss8i8vi+jCasWY/liIfzBL7udDJJjAsJ19leq/hUmaRLkZba7Z3
8VioifsD03pgBj0OCwV/Nh8C72DefYQFyMCWVBRwSaDaqLvENiRzevX+coqISl6RJWjBO1cg+lXc
W4TuR9bXexBrgg6k/u+kMXw8DJVEPr/+YIwcFnspSkrDWSPkc/Lvi3sCgINs4Tw/RuhngZ2ZE19E
nCgvtdOnrUEMF1sS2mdpMHQQoGXIoJWE3fRsEUkbamnsdeArvhzvmjIhLKiuc4K9zO5oZIsN0xpp
JoWpk2BBmKIh8pz41MXxERaRU6/1Gzmg1N6dg2Yh2BJP71+iDvagrq7sz05yDtHqvypnVPmiPmpB
fW9qUGnvcbCM5xdvrWQtw/S/95Pv2UhCOTTKbu4LkIz6ORBOrDdexPPTp/cMsGwPQ5mO1wdPNVyD
neO7EuNBLAKK8VCbMHjI1zkuWTPlnCPdgS57hF5Jd/klzBnEq67yx2Ud0GI9I8U//y0FAd10QZRy
pmYlW6wAyP8dw8Qs5gnXLA4FJN09z3O3iZSSxzmTyxH8BP+wOfAqnw+bzfi6S3FQ7uU+X5MYr4kV
Pue8gCKiMdHO+aDy70vJ6MA3010ZZn0nr6SRtvwubpK85l+b+eaulBFYL7dSxE4RpP/cq7zuKnyx
EltW/ADWOAdBg8aUcolJl8Q5FMrRrpMopM/GRoyNSmPYdyszf7U8YYk+eQ8GbEgPoE/IqdWoZCdD
St0/CYEqUH1CaiflThRHpnlibmsPyqQN50TZ2LGNJIxhidYtaKnB/qoMxdtGYBznakjsZ+kaDczI
nci9yQpELyJ7UfODQqaFbEcA8AK7ujGERul3r8PgZdKTvQAmM+2nfh7awqVjMs0PINKZA8OlUOY+
bKGnzHyVmbvXq6DV2XxNTvX8PSJR3fOxnUu1ALqGuwUyKhuRhxj8BWfVsPcb43ixHBvVEWvM+hXy
O/Qs2mvjBni97W7+Wp3It9pAbJkdBcFrP2EInlQ8tiofwRdo/QvcPiDQ1AdHmPv6l1BEVB0MzMHR
a3lfavBfKgvcUn39cGdIbcop7/WgwCqkIpgtcKincFh/+Asc6cmy89XeSRPZboqDUprk6zM5fQB4
U5OlCgzeO8fl0WE1/r7+QX9BDrXIBCxoObPl74pP4l/4Sk0drBcuVLFIc08OlY4gE+GJfUNminOi
BDq8QQ76w8XoMPKkGVQbDtn6epfbriTmri3mb/Hl1XC46VBQfTbj51ycT0wJYs1Ujj82/Nw4Bx+1
Nzd2DlplD6HbHvODPijXc0ZohisNP2Cw3SwAlsfFW6qiUzDo/8gyL3Ax+udogmpoyCBKQjgaOzhY
6YohQbtN67XClC2asgNjW3ox3zYd/5JA7kt1l2LjIUBl37BmFo+DKAdzRjS4p7pPPAtkRZhazDzg
td8z6FQMqYpbcgXDOSCL/l6tkrQiIkxqpf21FY7pjWM19dwZv+b+xZYVm+8SEAO49APlaz6PGkM8
bkmMCv//eh0zCBzFlFP6oh9OhaihVvyWtzQwXN6pNqyi3VUUfTCarfNN1GHxBM6d5DosEcpX1d2y
MKTUF7cX1toGN3k3Jz4qHQPPkck1Eb77NI/mJaESrL5AS4q44l567UniUpH/KwB5+hB7sVqv6bLE
KWqg75YS7YzQNGodouAPcOhceiNk0GRzmu3tsebJ3aJkQgD0kelcfu5qrcWY/66AHTwJDGg7J/FF
5Fluq1BiWtApeORSOMm2OAbxIPfVKSM57j9Unl9Yr224FSUVc/mczBKSTkikgNnJgIfZH294dOuh
7iOnwr0JRVEMlaVQDePPtJNl9Ij7VH7iRvqhbiqahKI830/xOV9RNugWUmssRq6/yWyDgJmgO36t
tytxc4eHx8lmts9YPvcOiT9YNncFWAu2FuXlyFNyL6TZTxPrfnmmfs95tG73cYywRc7Ez+HU2tLa
kxVb/HbrUtLrYM8grjr1hXnGy81GA5lAzNoFFrp42WedV3h9/zlY2+5o5hatLpDY91LG2NEjmVO3
cyfwNfogp+hOQhBqE9loOItHeZVndUWs4majXtjWssIOCMENGhpzQf+Gvu1hCXBnk8+ZO0D9lYwD
EuYPan+oxC02f20KXG0ngHPDBJ2PVG8XkfaHPB52ATVz1TYdppJMMTZJ+WI82xLkkyMIDV5wWRFo
MUH1kmm9K+JYq9kznVrtl8dHnJ+Z9youXlehhC2xt90dHdNeU6pUaWUBDGlBelWEWF7+xlF3HIVk
6kX6puJxOzyktk6a4wyPpTCXNFyR8Q9Xj2XEOkd2ZzdkFKKM98TTscOHiXMsuZKhiAPJ2tsX3MAH
D6lIB+Ml/ja0CkUGtGBXMwjFX/nYhj/F4bjUJv5Nn4LS6E1QtMmzdC2QnLICIdBLjnv2andXGt/h
r6MLQe42QoHG+GZPllm52H866bgtOqQoGpErWupUQ1KYg5FfnTAv4EWqaRRL+BlR7QfBhEeg8/y2
Meju7gLNgiBLEjR1QN1ZSz4dSyq9QBuM/VTxpaZ6/Yz8zuE/8WyArDeLQZ40IQ2O2RSmUOVk342T
thzVANUgftsUwtbeCNGITxKffzoYCRPOAJpyDP0MDVa2CGDNxLOvicTLWUaKChlIM1xar3V8HrTB
QnTruKk5aMUoORkaQMptDMQDUVA423NnP2Tk5KxLgSuDQZaV+fKTpiWfodOWAPcGPGaCnyZOumKN
hSytw+hGa4FFc7brRetuI2y5PORC7TAIa+8xffyPG9PjewQy1oz+f6nquvBjZ4yCjXETpf6DE0Qa
DyzVLC6GmkAbGknMESUkJt6ylZZgDbIwwI46bd3MWk5RhHcxARWL8w00R8dgKfJgrCzUPYlCRXDn
LOd7dN/NuvYfOlF1NIomXc3G65fVB7cFiN9lL3COVSnCzDhKM+LIGSetP+FjgzReYuTpQe4mscVL
AY2mKSjCrIu/XMSMMCLtWWSjUg7YB+JUnm5WXh3wbSPIb5gZEl+9bLnmbbMGSIk8tjZUAyYLz8Nj
4jlY/rsRccZ8XNre8E4yaUwQ48YMnkJWpClWFSfu1DzVdvvsM6Ez3PdBPnIBxmWlvj0ZfCPTA5TN
om684Bv+1A/+5Cpui4/te93NYnC6VlhQqvdVLuLLRMDjrmWVVhFVm9lqf7a/pTkipLTIk6E+TrP6
FG6t7Vyd2XP9rDDSLUJ39Q3DH7gzak66WoEobc0MO4iQXNPErvC/ZMdtehnQdTSWkxD8mpZ2HCS4
sTulStytLu5HtVcqJTB96336KLx5vdsJTVm6jNsnEiYcyhUaDOl8WsIt9xhFF78lvKr30dT+yT8D
pz77tGs70v+jNK/ns/PH1hMnM2fJfNyqNe5LCVT2y20yCoz3h/EU7mj8BUM3wpg/WI1LXNLQbzqu
H3n6oWGeS40dWQEYQFFQT4/npF5oLRauf3Z0sfdrkB4035W2KFMxkMFqZQv48tu/eIFT14iEk/hI
RyZv0Cj2Lbashpjs1Z1IWIUf+VamVg40J2dpRF5WMp4pP2C8gjGBR6QDF5DDDJl7vBLYHTMm8+L/
YbpSpJm1vvYMkHblwetlFQiOWrFlPNg05Xi1lGnEl8fo7mAf08kwWbGgqHFqt1zGzV8Ch/Yaa29a
iEA3/SFZsQIEdSIzJ3ewPOVADaEZzDcoAdU1Z/ssW7zEN79ClNCmI6R0QRDURgeD6Cw0FFGMkV9R
LtakWcndcnFfDkO+2CikHEoAmrnCYWbisDQJ9PqZWnDHIjsQZ9bYDAdJtImcaovATVhyTfFJEXFl
iwFgNAZqErhSzdTjwCiozO6Y4DkLsLmR6mja4k8KBsUNXFMkgBqzJ3HVpkU6Ydgfm2djSItVNA27
wCBLmWcjbj8i4u4Ga3koKQpTs0Cd53DVL7Xq0P8A/GiSzpR/xh/4RmT7ivQ1LFDXtDF4DyNl7yGq
YbeZtxvIdFXc0aVL3nsXWWUcaDdaBQ7zTaRurng63Dk1/ZbYMGtDmZq3qZaNFBjViZKEgiBQve19
lO95gBWQcXFEZclAfCU9xr4isDLekJ+5DNEAse3Hd8ylbjpMjtntd3+nwku9jYyFM/GaGSM4Qnyl
DZEpqHLg735TTXCuXkkFl998OOI80kiX3hqwGpDKMDHUTvEdS47ppFCUpGxvNfwjwgbrw4GV3ViD
tNxpjNgdRlVjelVbD8WbU4UViooTnbMtenStUfuGKp0In7KXthjNBh5SlwXwYv4opAYHWtbvPd5c
r1C86JO8jylAXcrmOlixiekKd4BjoNvnwI392/8WLDSPrx1oMVotoDgSQEZ6OSZoRfjwPqqHoYPm
YptUkGhi3Yk/VvSEPaYgGBfQNEJh1cMnp5BQzQcRn2E+/ZOM69t0m3OpWPzyNW/TxUP0tNesiCin
U8ZOuXd59isCnEmzI7fPK1ALHTEQJFoWhHeHTVEGl4/0m1Rlli2nSX+ey77ba9jeu68afwcLgs/z
m2VSdZTcLcHbRH65TmyvH03jTs2Zj3+QQz2Sq/CDtDgzodwVJmXjVAnOxyRNCNMFGebpa6WT3bmD
QzsoHOnDlmlZaUm6wtfUzqAj9Y8t8h8zRI1kF1R+niv1VI8Io3yxuAqrTiFSauKyBZgWovU72mXR
LOJpqIdV6wzGKVVQsoMkvhcBtWhbT17KGTUyusXuRfbOYr3iDWEMA2GiwCza+kBnmbMXelmmQtrh
axOiOWPo2c5lyUdObqokM0Y85QMswcAPFlgwGkt4K02wI+4DMvA6ytyioR1VB0fz/MwBP1gQ3ICW
A2Aytxa4Nv4UHzfPj5H01Vom9ooEVGdZyFXWQfEpjVgfrbzBsrkK59cAV2ZcY/rTh5zVnNxs0OIS
yoMjAh94AlqVZYR8h2V6kHmpLMu3W4wRoXf5zXfGw2ErXntuIQ4RSU6njbg5WLz4P1ZuK8RgrvHZ
PJHXvK9EMd5tmBJ/K/oe1+dxI86jgO3gWDT7sjrM3Kf9mCGO/wTdzZcKlOYgJGiN7baWVue66cql
EDsvIUTdS1Fn/fpeDIoUk8530mg+h5jPDEi5mEMzCy4TjcJEFtpd4aGTu4hbdaJ5w8tpoTGb2Zs+
L0ZYaeotJ61MRqjtk6U+uEKd1jHVw8/wCcLPMuU0u/DlRA3QttbVZ4liUh3AwPLV+6wP1XwTokQH
fOOOrYQQISiH07CFxKDSwLu0I+HhGLIrPU0OIa7oEHyGhESdCIAvtRqQ9x2KGCxfhcDedur3VWy8
kM5cW2qJNGv0smkXemZ9K8YrmKeQfxVKK9MHd62bvu4TWHRlOutsqj2kWulk7MLJhnVwyxFhoZac
4Xy5pfWJ5CYulM4ROcI0y2HAOjEBYC0ZSbI/HRUkbVQXKmr885vCV0Lcn3qNCKsDwOF4VpqsCkmj
C5EAC7Oufn9jgx4vuq9DoGqfqRiPCJeUFF7GN9ztc2q+xwurR0/4+VekFItjukcC7ZtDpvckvSLN
RcxBMU/vXBMcCY2Wb1KPqR61osipOTWbWj/ySRGnIuEdAoXb8sdNtOZ+ZClUpW6Bh1AcZnTJq6eZ
y3SrWjs/qD+FyVT9jlKdWDFae8icNr1M61q/nV3OuOBh0FcewynDXnpLis5bX+7TcV+JeVdamRQO
+rVc1S8c+6p/ZZFZSKEKrDkqcVTfa0xo95XBLpPdhzIuGWOqIBa5EYfc+7o3B+voA87kAjst8fk4
0y59MaFTeDcFFEsolumhL8IDsQFo/+BIix9GxRBp04tC/kZ7gnFmp6tIsapQguGY+TmxNWDa8qny
XZcrwSuIxHiUP2gWvMU05V6U+ypSv++A9fiEJ8BJ00bnbXpATFyWdp26mGaaQ8lcYMQaAPQ9CkCn
cJEP/fDcaCfCi2VeOUsC2C0DLaAt/DUgT1YmTQxMmh7/rsJvuFzc325ft/j0zqzPlbJYV36IvPDp
+JnWZktnia0hMikoEu4iUWhI3ml9AURu5zPjqooh4hfbBk7iEhzyKSV10ucaZOGWT9btU8jCnVfi
5ZCwasighOk7CH0TM2470JvYtLLlJB/TycACYiDIybN+snZ8cZ70j1q6QE0CwWdBzdd2S6iRVSqz
3dDa5SJ7lcWMjWj+noYjl+g1i5+wIQmB+JGlHXZaOCQg47UUMrUELm0ruqDycdRhcT9MBwALeuno
dxBbPHm4YVFjXVRFORKDYFVXqsSnsIxz0h+nHrnWH1Tbem3w/DZyYauT/o1Csu167KM/kkqL8zlo
yuLX/qLeAwu4GBiJoU7wVabyEHh8tYg2sKOSl2915CKaHyivMY+ozQhyvTLoz4Y/yDf6uqLPO/M5
q2OGKTnMXbBPJIaB6brZInvk4GM25olPjcjKIIL9SDJfwVmvhvTvo7NTmWPrLASbcDLr3VfsUjB/
u3RPOMKhbgdg1tdKGVxYJzt0Ww0HYiC1CiHRtHrnCToGUrzjIF7HZNVLrx26Ch2FrRXYe8lnJrMZ
Um42czBSxqGiWVF7Eosg0cAfQVSQVWS5kMj1U2tcx6JUXl+33OxuXHpiXZv615fLkuFepVLuH1T6
NB8syokeDIV7HRbQ4T8mMQ+nodDYGtIEiE4KX5kwbh8zvv6Og1aB3tmm7/SSNgl0omRTnDTPzq14
WhyPsbNZvjZHDv4fajJTfLeYiM44V6ux9JwSM0aOxYkJptCUsPtuRX6PXZGnuLQVGa7lH2DQuS7U
bK7aQW/mLl3ALauKLLrHS75BLf9KgoeEL5EDg6n7kafojJnwtgBaBPnRNw1bw6NpnbUri4IwhJWw
obvA8N8xpMMxnMbAA0UoqVsEl9frQ4yzWPKGjU2EVh53AjhTW5RvxEcjyeYbQHxZ3x/xGrE8favi
+aDj6xiTCznhVee9J75eAiwZV9rbDLVntzf31NN865uDEKhJfCT2g4XXZrlVKf78nNI0N5kd68BR
JNzzngSCiHStHgV8wtHgZ+zHBt/aGSmvHuMQX0d68l5NnerabbXSHJfH4ShyBiANC1mTwOPg3QQG
5Pmz+5RbYSLrZ2nfulEsA6vN/Nvtve0jSvCqEmX9I4L6xrZSjqjRiHYSYWpLpehmglNfHWSLA8zc
uqNcpF1gg99MVFOsxLXkzlF7D3YldGPeS5JMhv9I/yW0HeeXeFAEpnQQMzdo1OpYtJogklfJbrAI
DdFl36jHhQdy1oRmhjkp46y73MrFtCizC+ASRlgu2AowABJXMQ8MiFW3SUVsY/HcEZ2Evox4diDl
ebNi5Ub/Mp7BttDYxYZ3Jompgan3IdIETDiaZd8uTzrn68V5kIYXeIo/ms8qXwvp5QnsZLq1QhNA
9Pm4/fGPeWfSmHIC1SEzak26Eoh49SZ2cj4pZl++dwqJnEabvZNOtqy2tvUANVBVrDr3tf3ZRaiC
Tc0ISyHnX8+0O6hLxQgUg3nDsCXN4KOr0uPqBIzHbMQ3hKwf8nhS/rakpQOak8ehcUgU6zW5Cr+2
hUk+YkHdD6w8wlijcoiLLQWw7Y8h5vcC6ElbW+8a5zSVXGicXWh//t8O1u32T+LSG2sesim+WgMC
LuJ9ltsrwrgj1DRSb38BcJN71Q+R3coEqiHpi9V+Wedv7iWiVgDcHaZvDxFn7ND/NihlWKG2tjay
8iWoA0eVJ20zr2e4OD+BRl/RdK3IKvObdb+H7YcpZJl/kmmfi6OYNvsSbuw2gTbcg4Y9KIKZJ1Rs
mkvcVVJGUM3VoD+wGwr1yyB+XCow+hLiEDNEHHUMkFpfnxNTByiA0mmQ+pv8gAf8jk0K3avMkJ9S
KAYr08ihLlAkrt6C1jTYd34wOEfX/WB38Y3gC6OeMdkFSW4iEE7TZFd4JNU59za+4GmzTMbJDtxB
ikLfRrGBx2S2NnboSliRCI7zvgeKK/CTj9a6tUoQkfI9UUwxmQQTtbhl6tACTt91r+k4ZXtKwUl1
RUnMUspdw1PkkvFLd9MQKUfKmHhFL5f7In5f5LGhY5PTlQG9W+E3CeNX9MVXmCTPQ57o+YhH8oyw
aU8G/po4DBDq98DVKyXOYC/6xy5Y8tZwAAXNO8zNWQXu9HSB2ETv0cct0GMiwSNiYUkJhQEMixaT
SkPwYMB2Xz8GU43CRKqCxVXLOeKzeO5L0YkZx6yweX6KBKOsmXaIKaA9zL3ZqhEDICNcx+8tqdUw
u49iKB68JW0q+Yhmk2hQDm9r2UrfOAGgHEyo3WsVuL/M1tUwN9t+lVsclXifWTCJIsIj/sNv1R/x
VSurL1ohldgWPLnPWPlWseQDzNy7F7xVWWdOXxN+pQfur2xFtt3PQSV9W/ohbfK5rS6/yfmtdLL+
RWbbZL1FC3cXgGbvlWXZKx/UCX5F5VY7orUmWqSx7sIWeYYceLktjWel18iKPz70hMEFGBXXng1m
xVv695+SRFgIjlMbJtRt7EHBLq1Q2QJF2YtmxTwv1nJyIPtF8L4CQvpFofoYYPsqb/B2EySCLW/B
C5Fd8QZaVRVKJYT6+M8e5Oh5AhmxPvbeKLOm6duq8IU0oQTd+7v+JfbHg9ZAEA1SnMO0/d8XptzA
wxOlIeQ74oFJKysP8najvHEphr7lo9LpptKEmqnnq1lPxi9vpU8g2/WBqgm+5hVDKMMB+eHgHaiI
9rePx+n6S5STvTiZw7gXIcbN5OmFOogapS+AH0nFTYGtVteC2xUcO/GZycJkbv/Oq2YIdYiCGhem
RGy2XZg7rRMRnojIXViWj2SNYL2b/axX3pf6eYdTvNCcYEmo7b+N0ikXUJRWu+n44Kpo0v2chDe/
nT9aP9tuW6ZN+5dYUxaFPb0ri8EXNfTX3quXQqFQyDAWm4jMGwQC83Vct9G38/treM7ywvNmXbGU
cpS69TNVrvrN7sP6oxHU/Tyjw4PmH+qNwIiNwAe2NHmPtQh1EZmK88RC07chUaDrqMvF7IjvlbQJ
IH1eunkOjsnDFCgbvot1KV58GgL4SaA+V1WzY9rt+9+HMBXBEG1skVaPe+aNw3WvrpXXPXrTQCIf
CePiRWJGcdcIK9fZGriNW8u4WhPZOj+mGN+VJ+0/3DnXfl9stnssugPo6kTd4HtJtsxrW4O8gTvq
MUvIKFFX+GvZhJxn0KLPD+GkZpFnUaqFMEu28x8rP7ZG0+uxjj8bAtWiziHoLGUile7kBynYM5+L
0EK8Jfp4opLerJwylPr1vAebeBjV1omFpO9KdAH/3F23xEjoGU/gZqETFIiUc4r3+UHDOdrcS4F2
ocZyMk2IRhY9GB84oCmak3HSU7HkDdrqcacVYM1uuWpRWPxFsKQIuWTXeNRLsORzakNupr/cxYGV
fd4YIWdPnrU91XAadc6EUC3JtelBo3zp+FcvmFC6Q/665S69LF+g4pUal0B2cTNzu5dhKE1a1Kxr
xFkEveBFoW6TLR7JdUvitahPUhFPlEvk0/Y+j/LXrCnJ00ST+P/EnRgtRz1sv5AMAXjK5s0Z72ME
OuKSG2zWRZ5ZdGZzd1UAhG2Y9+xxf9kcKq40RLHZV8tVzOmQ3CF35ZWjqj8675QrDKPMNYD0t5Tn
gTkXNPBc6gkc8LF0Ow4iFU3WQnlnPKkneDNsHCyeCbgljIutRObAemzpmMJJrQGcTitwBm/ss+AE
p44m79ptkpDcUnsyJ3y1BCOfPd4jj6eycIueJ6WhLGeUa6QYnFsUNi6aP2MfAN5vY+Gx9EFb3W0c
Hu2qF3iAlfWE5+3nxVftzul2atr7SQ5lU5O9jY2lvznerq5yYRhaCVh/Vt5cpndnHSApEUHKDYPD
kHm1c+x79fhNrYYp1c9rKHCvoqrcZcLLIQ1760APgDIsmI7M4VrfPOdBkN5xKgr9kMO9dYEFA/70
3h8Titc4YDToJwbxiVPrCP3ebNjTF61d6MKfLnpw1PaZ8oP9o3CdTvP776HtxAbucfZm0kb8Kyia
R2JrS64FpGbpzgWaj2DBBiq1D4HehKC9jwnUbsLTqw/fB4xMf6I3i8FOBUvTtGhrJRAfg1MJRML8
kEIjv4ZJ1CspD7HobzSAvygnibzhkVm9R0T2ZfVs8Su3LcrGmOb6xQeqzu/joMpae7WpvVfqB/7z
xBoz0iF/e4sWFazVoQOaqVzahIPucnrqMHGcBqrWx7CpGohiFHfSjuDg+bjwQFzOydJb3mlF5S4Q
Af3TbKOSJmhQ954yBKjQCPiqj4S2VWeFR/qeNv9LSzI8JVRtoL2gKkjjMenN0aMhWC4n5Xg8M8vv
W3Hzah9S88SiZ/NQ+iiJtQWxzF0WjxgFcTCQmqf+zSIGeLf1YN0ZTcr92LGDLvvkdB0XC92VqZnz
xXU1e1PRmu6gQSxsLOGnewKR/HVrcXhNgZGFN1hdEw8oT5gk53Y7iRL4vMz2037NDBdO5bU2y40g
944vbg4PzbiNz+RrmVkkfFtdMvVIffUpFi3Ao+nqanJEuRmUbpT7hnJAtx9fnrkyIna/N6mt3ikc
6mUXhIO8RF0wBThWkAyey6Ytu9THZ4bUd/2jiAMnnO+lhiLX6tKlSrPpj9e5Uus/zWKvifm1jOJZ
V36zI3Wh9ugynR9Wm+Pm6+TZuq4LQrJUzSFi0eQY3EgJJ4V9W9zsMC+iKSnQ+irAO5c2/uPNubZp
MfMAPYe1siE1K0LF8hlJgCgoxsF4aJ5b4JG4YZJYSI+Pqm765nch65c592xYZffjia3PRN3lxNKi
01OZ/KVn5yQancVFpbWqA0WXXGg+jGCzoO9Ca4QaljHwuj9j7p0F72XNoEQ9Ebtaywvo6OXqT11y
CFhlBjRTimkpZbyMPrbc0YmlD1SXsKrmweRwSXfKyNXZxvIebZ060zh4KHzX9r9T9R29jKxJ9R05
t54753b4H/ZJQHLWsoGIYWucGbMNImw+uzG/7zVCP2OauFpWaac2Up9KcfXkcoeNtDcnCwX0rzDG
bhMIxYkEbxyp7mrAM3zsPNRCbZSWty65aih7VXFNPP7gsbLm94do2qOYc6DpmCWJgUuXe2B+Vb/Z
Ktkli4ADM2sdMyDymwaHDYU+W2f6uTRB0VP/UolJOtjY8ZD3uAs7MwRqcFg7I8WiYb6/wXhxi8/a
KkQeM+NHloSIrpnwiMtnLEUpJUAEW7gbt8uMIQvlxDwWPtKxxqqJugrSyrFphDQsBZqGjUpvYFkU
F4E5L3daIMICRTucn0CT29crazabE4xMAtDO33Y04mSxN5/uc+DG9K3wcf+RrdvY28+4yoEXc2ke
/jeZQ89SbTKraIsx95VSx/zM0Aes/QFuKc1PGrXVa1AaQ7z/gZUOWFmfHGixWCYuGv2PUJb2qnrP
pimGrbcU2Ab9lPHMDzTytIKvR2HMaqMVqLQuFV00XXa6UxDDE5/Cynu8EhR6Aluh/yBwWcd+vNkx
M0pFdwQDF//ThrXzA5KXvSZ4dQ5giEqJlQ7UekcLeP5iYeQqXH+5zo6Wo+S1P+WHdR4hMkRTqwV3
0/37VPhnirxgUSzesTx6DZieP2OKN7jH2ljKQ8tgRkNBqQKsgk6k00zXpKaD66eNSupYVEZLC1vU
UeBNckGRxJVxjHyAwidS1O8ImYI5Vo/wsWRf2BlU7OA3iocBgTyR8Wi+ZSU1inYk7/X28cMlhuSv
Wc324gYQHR3DkZnRT3T7C7tGdYcQimyveokaoo//bHbCHiN9XlNvDOFm6XywEX92NuilBqKO1gGP
6PKnSX3g6p2LNHW9/zekylDp3TVFRSLrHTlrLlxpkk7JJ0NHvX/F0+poDY7JtqD6/D2dEfnf7+iy
u+p33zPryTU7z3QYlktPbocpiSJij561kNvHWqm/YJ8cPSYHMraVc/70fjSjXo459H/giYTdkORI
isIlu2uWqGdHhRkPicPNF2t7wZkPFqXfnFJkZmk2+ZGKHVllzXMFm7ezCDpUDJ8So6mhzN4EOpuE
m9EH4d7y1LiJ5msLzfbdt4b0aDMV9MuUoDDjGCLP3+NuHofAofTCZC1oOhfeBVQ9HbQEfX3TBD+J
2wL5AJbLpWDeerRqSpRF3bg7FtCgCqN0mN6b/HdyqL5jesp3e9GE4iPe/hFy9/v2VfCPja6KsrAj
1+UOh04v44Zfk5cwA5ThmBSr5aQlyt92duC3XcyCFRs+qrKIUS/OzMYUXY+YPLRdjJfUgdkXCkmp
iRYa+hqlKhOxsfKVHzCHU2lhn6xv1x4uP5KyCVYTVaQfr7rtzsJayDWdTN2Scyw8CpINgP3SWQXm
iI/pshKXwAdJ+0pDWwVsjLDo0aN91z+kOgBBS389x7fw4c/kjikLUMf4HcXi8Lu8TK18400xacSg
qsbLkcQumAh2YB1hqa5A6pt7dZcFb9sb50sysnZw4ZCY0vkMgbXQp5o/mWLwmB+4blbZa+AV8w5d
itItFgNl++QMj02YCGqLwLC0Cpa2b1XwFKnfWFTGVosgU2iGQ9GNK5JzV6479EPieLz8Yy14kDKF
pUySZ/xbDR43fnMIRKKsHoEAPJ5WSlP1z2bTFb38/c3vmtOPIVrTidavpv7nLBgIf6S5T1Go52zu
n7NgnUPVNA1OyAApIDYrOA8y+zfeEsODHN732WkpG9Qy7Fbs4/K/0XYY7qrlG01FInZCNoUqKGJz
WOrRIJVGZH2aerZraTGNK4bquf2Pi3rbJqVZUdgE4d1P7NSIGwM6lC28DCI5aBk2GBj8ZEbK22Oi
X9BfnUYyruPjQls54Feh//k/uEChyosSCCH/YSzVpu1qX3EcnkISeetkRyTMxqFkb5fXQdGYp6wx
mLym62dBc2fUO2ajhqV1vMs6qiX+LI6u6sRkkBI132V235DP1NKmNdxlRxMQgJ4haXNaTL3sAqjr
WsVelJxgt42kNDn7nuX89500N08yEYwg5o1E7PFjeSzaJyL8jDVX7khJ4LKOCw44aNZaosJYa4OY
uwzpWDG5FtEO39n3BYxlY6ZHQwQuTsOAsPKs8ULNvRSTIGSDROQW8F8zAuZpDFEEkESOW8sbb6VZ
AVS7uHwOZMI2CYW8n3B6yrFld7w8Tan7MgGd8aZCX7NptwX0jFHin7mmc/Lvqjg6PeM/fv2X6IoK
u3zbetDnvSvQBVm4iJN00PAkAo6Pgn0KJ9kDdzUe9+WqosTAjcccTP0y7VDNjIqDvjn74D7ZHwBW
nCyulW7HpEq/q9RR+4fK2qsNzClkejILrgrX+hS1gPBmesC1FU/GTZ1Dt0r3frtz1wTHRjHyXbOV
fTjU/uRRSK/ElArSr3S1fM7MDpYzngjVuhjs13oNWRGbs+XjCcv4wMI4XbUz3mFW25dPaUWcbzP6
9Sk6bPQ1MoiqxnrBaAzmKEhj7NgzWJ2zlbdJUeeugb0KaplwVqd1IKpI4hzJ9AZDA/WW1B5TxPtJ
FLJ1mi8mMP1otKFP5cMKq3e5Fv3WGPO9keXxLNKOHdDTUnAs3Xte+vy7vyLhv21f02hxb5nEmUBd
Wrs4NRRWB1/wK4oON6TxQXBjPhM4WlORvP8Ka2hBY5KmiQte7bcp70SAlJY1LM/wCooDUpRp4Ati
R39AyoQf5BO8I7TBOZ+OdfTsNe0vwnmqk4N4c7KIWg9HyXVpPRWquQkqsjPd17aJnqPSb2kMAvUB
O95XYG4drvdd2+WjozzQ8TRWP/Fwf8OU4fFCManDDJGDGxUcV2GqfkpWLA6C+jIbnmXdAlsle4Y3
S8ePhhRuj7/6FS21AGw7hVj3BkPeVeIqJ0+yMD4bsoCopn0R6pHXmaRULJEXUEINuOtx8xiKU1YR
YdP2fmXm/cnBgyZl3j6FiR0=
`protect end_protected
