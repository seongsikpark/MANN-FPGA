`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
aw3gwA0pkA1KM0EzU0fWDqpDBmki2pv9wCQV47fFme4JKsq63WG+ADCE+vbn7Hi+Z3/OAuKb4EEX
dGenh3gQNg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
GigQBufnZO7EfSHP0Y6uevwpckWE0sKJaS4js+xivY48qGBeSuRBIXwcnXUOYHc1ZK9okdNAvJwQ
JPNh76bftVump10ReYTgvWpCGfLwjQCmMQgfqzTuUx7v6mXzXkHNM3AF9yPZCD3vpvtPZgQmT472
s+pvZ7tu9fma2LULf98=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
psR10jh5pgqZ3xweJkjl9fsr4y2yU1lL9FJOcMraSNIpnfe7ZuXdAFUVc4ih4K8UlWax/IkXIlFZ
n1Go7PXhFKnwhLIovoHM5Jvl/aHMnonGGRE0o153utTtS+2xjpe5KLXNZCOOZkHt1iYsRJNgpalq
Ec60R/l2o2rx22M8MV2QI9VH5n6uir/9OOojjQSi0z76+QbzIix15clS2EM/KdTtUZ3N3oc+KXNb
M0WVoI19ToV40VprGKM01OBici2WucYGjiFP1kyi/Z0HoPHzjqKzAbwWnv2tw/U5nGwl8XzHIrqB
6RuMYMosIIDOeLH8KbgRiQ9dk+eXqTjkT6DaFA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
I33xl8KW5axmztpTK+QsmLAzENZuPcE7t41lhXfih+wjvg4ilv+yHoFmQGqQiA5OM8uI3vYwC4AM
uhXm/XO4za3bWTMKArTaogU8bQC3ob07Muh6+PRgnAPkCENTQno3WFMqNAT9VF4hta6Ms0fm8yCH
mYbJdYkWwfOzPCaNq6M=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
P5FwkKjf4Iwwox37r/di1HGRbWXhg6hz9YA6uwui7LGq8dcYaQkeLr/GG5TGCrlD0NrV37s2LSbX
7AfoQ0uPsN5S1snAl1OJw3RYmlGpl9ibMHbUN+3sJlFPQDBKtau5bG83kELMq4kfchkNasGTpkOE
dRYrbcvCIB/P8mfl5GpFxl8+QUwKwaWo0q5QQMl5zM1EUknMP/KD/TxvLLiVnpCvfUu8LhZGlPzT
mNjw5c3aMaPj/h7wJZc3woV3ipM+9dh+PE9NoHqZbgPHU6murBnDmTgvuL4kJuWVzDB54okyCb65
ivdndVdsfQ5rKcJcHoUkja+vdOnP5oizOryTpQ==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
CxoPsRKVWfSyg/9xz4OvBgE0/+1nmJV44iU931cbXYa8QCvRGQyc65x4pNqQX3xCsYGV6DapTCDt
vD4a6ao9+XAXblO1MzjeCgQ3dR9GgRVA1T40xYVGduF0uzm7xeFtct3ZQLoV2n5EURYqM7Lthpkq
m14yKvLy83eQwqPDs13ImaOVXdczOU6xX3ynkh65ShlRdsloyxNGOfXYpbb7r0IEad322Y3RP6hW
wacfZyIi2bmjbID/rU1qpxootV+r0jgb1/wWkBjvG45gLFr2NH2YbBFOr0w1OHD4SOYw9RZ+lPa2
/3iRUorjuHYcx/D50YSrKtQNMZZgT3U9/nU7hg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 62080)
`protect data_block
VxqvZJEyVHWi54uYo0wJOdzuSmKOlejy+55whx+aNDuo5utyaVe+ccmqek1l7nrg/7Yr82gBpMTa
6N98BDGxm8qkP9vHFWtiNmO2f/T8Ftbfjmgf9cWbNbw0uCpc6dOz49mN7aYxYB04dzNwveB5XSfC
ehvBmg6whAEPtXXqDrICFwTcOXFMlYie5vuVs7vUP0jXc6LHDDlcwJ4XjlYtDkisw2wHMdaevkIW
f9/x0LSE6EjHvd2+FwnzXuHPiC5DmocPUXO2uEHq1y8R6lKzvZAkw6Bb02aBnPuAeUrwp852HMv1
xG+Nc/kQPmWYSAKgUAdlvJTtq1rGR8PjPkkgUTmTI+pluXit6QdLx8Kb7v8PZkOcuxzVliX2OwQC
Fn31YDJJ3/5HWl4ftH54yGaR2XLKfrmYGf3UFK2DZf9P0PlrceettcBZCVj3aLFEupZp/J+//kwF
Ms2fIgxlc16SK9wtnaV0rMFlN50RIv5FaT1K0DEmyOcwDfCDpyME1pqg++qAU2F4WzyxME7d46Ws
/ksryzWe7OBe+h/u/7W55gyNUYgF0sh211HMLUA2NlRUFBouzIdXWysId4TO9wFuqJ4LoU+JE0PY
kGgA0abxAcT0uKUDeWIcOxrL4/Kukfoziz8tuM64f+T433burhCfH2VDgCc8ok85L0b6RjcTysVE
KugfwlP3Onp8ClxIqoes2pPzFCVB+yxHULvzcZ8yW1a/hhSk4hv2M1/QK93OCN6wwsu2ZmoSOPxT
JibC0lq3ZuMq5nJQ42i7ZfoGXvVhAp3bVkIOzEASii5qMmm5wtfv/6dthyIr6F2LAf2c0lzsLVjg
WFrL9zAhi4ox1DfACkfZa6sH337HAXwbUiPdVH/ATyy+BrLHbYuSmSLZtDsQ1SIgYXMYgZusZ3q/
3QRfn0/hadbh7fkTPL8vbB3Va/ZTt0/jFbRIpEsejiexGGeIVSodX+/YDpTDS5CNqLz7GArfXsJr
eslV4OK65a0NUkclmtO9AVyFKCySwGBN6ChI2stjZuAOvKkpJ6zl3A9wLa+EVhUrfq8R9TA0lkqL
8ADxYj/x9TUPsKKeoILm3BflPnSWXeQZrWKi9aQawZCrDEu7Xr9J1b71OESsWMo+3AEq2LMxcQCu
Jhl3yiZLBa3OVsGwZAtegekTGfiD0+PFnhjn2kOfTtGkS33DgAT4PNIQE9UllQ/Og3GraQ3R+HgM
kSS52XvxTSbMg1MjlB5ML+H0RA9s7ah1k7rAETKUMWq0T3/511qjGmQHH4L0zUqMBBpJRKE4ZbuA
hu5GfJ2meq7221IOz7FcMzfhEGJnNFZ/WSyl1GsHMDlL67k5hGET8kjGOAg3BYeUJPDBGe+dawa5
GsVkHcP+i0BioJld6P8Yn6kAlvGanfLkp72SKadpPZjlhyoiIM/ilMWwy2nH9RuRhmuJfx7EgMXm
linuNkLkMEuQQp/A2UMiRmkcbQaIc5+GTXbquzrdzf6yzlEYStTST+qNoN/h7cZERU+fxn8z9zEI
TTwIvaW8oFG2OFLpAYa9UstbpOPYzmLclaHZh3ATNtmP7PLrsFuQb8mcEOFzbqiQu1kSogRJeaHl
yOAJZMurtWPHIPAyxSYlwd/SsiOo8mHgBmUOGV0I2/Jvi+cb4dPedcHfsHYe4Ucb4btHh52QR8k5
yigrh9qHWJKuCCZSLOeRsc69T5hcEdJC4mLnaPNE8Vcn3vtwpyO58icoRIcBFALdpbC5aFAjQsuK
7WBddHu+NCTW8CJ8hHKjQOThHRMS8YWbnY89q9HJroZQTPM4uBEFZfjU7+/uT233Am8/wPRdXI3t
nJ9ySVCPAs1im+svkA4ia9M7i9wRtIgGytUT4ZD52eLcynv/kMPz1dWMIdaDepOENf8y7Vhntatw
kME/bau88n2TcOY+ehw2yXutPH5Wdsy9kNrZkebDyy0icmpT6sBrccR0ljzGBIp0/KBj6Qz4vv8Z
e0ELthhwXEivHJd+rcu/YDRiwoc2tbDkS7Iu6Ygn0IHQXARDq0EOB3VRUZ0480A3dRwjhDsf7Wnh
f9ZLmn1q90D4Yb14/oVhm1uwr+Lhbhy5CuzkSXMZlrgo+wAHn7a3hnntny+DYxmy1PB0dlx+5ALe
ELvJYpAGa8SIlbxGGekao2DM4GpmIXrzsnW//vhEpTolbsrJG6QvFLAWacADJex52WhLETEsrcoc
STsIEOlRTft1NKLWZ7kAmZeROkXQ+RlI1+JQ395UqoUxc6W7mqwXLNAWSDp+BE6h+tGEquW7kD04
FM/at7mi/38C+3SmMpnKW/9MN9KxpvIq0crupL2CiC9io9iBQOVswHgU8cVtku0TZObC3un6pSby
p4UZoZObvHQaPR1hHLMqipBGdp7NFUNygGW52Zjh1WlgG9pcIcypeDLvZw2bU7mF8A8Gg8bDomwe
/508ELnPup21oWO7cPtGHoqsx5DGrL3XlbXa0F8kNiOaDFY8UqIxPUubOMUn9YJeKQfJqSuArlz4
hllMvmPfH9vnGhC0BxZmyd+UQ836qLVxz3KkwE6KLo8HvMyaWKdLS0dg84Ks6cqWx62TbuASYulC
oRcFeoTcHNZtJNrI3EmaE/3mi93Acamxyrbc3XV2gbX/OefLIOBit/r6PrRTzMHiNQcDMkqFkZRH
FLDLfIqTFQE+O45wnP+SuxxRUv/GCZswO9QcpQTSmJrvHHhQurEHHqCYMDURzoGaejSUjKaC6/91
UBMGH03qaPS+OmhkDpfLV24JbV+fBP9qWzRR40KMcVwub3KFZFKoojPZglbZpbCCOs9aYQsTCvjG
Hc9rwEgYYeUVh7EE4ztmDzxoLankUmpe2HB1n9F7eCnr60XN3CXpofXcyCX5vAdpG/6861ed9TZ6
BY6XbSgNmaXZ30ewkdABvO57xELSTMGFa9GQM8OZ/E1hRoL8O+BD+9bFFMKCLH2HKbwXn8Awel57
m/Qnf/QCpybEdRkwvYYasNncPZUjkmSE27L8vCuEKP42U2xRK3k7fV76I8iwdLxCkFF5xlDoO85c
HzK+80J/iX7dLWCNq7ITsMKWhabrWgSoh+9ekbmoOZyn18YSRkgbxiLaEnUowxl8UD3NBKK4940X
yOVNS6nM33HM3a44pQk5cDK+0NPk4HfoCJ+mF3l6jMEkOiY91KcSv3JN/Xc6wlRJYo9V2dLMi9qA
iUe50xTQfJi6/h3r81dFFRoisGCwlkfceDew5/ihPy3R9/+1QZd1DmIVyJUkcnA8COr3JfIvrcgT
tGUr/Z6Cxhx0g2ar1bYW4hFgz/Ctdw/awBQUqmHx2dKQnDlaTYR+euL8xLoZUMOuQXDRP1yXw5uZ
jWANxbzM871xD0JgiTkQFtabixHyUenntvspd3+J5s+cS2UVZ91Kvx6ztD/UT8RwQ73e5GxTl093
sogyCpOQW8kgLp1E0w6z3dRs4oaT3vo0gidVJsBG3vRwyUd49/VfY6u6L+WCD0Z2vBL7Kv+rg3lX
E/OxLoGl8G6P2xj8MW1e2n6nIWp7SWhF26fPvRoVaUPfJ5zgWMWmV1q16CvTnjS8/QRmE4Nzk8hC
sNJwQvTeV4HGEBbgOPCwopXDEdEp++W/8zD2rUtPgPy8yd9PeJ0cVU2Vt97Y0YpzF+A9OkyKyN+t
x4Rt+B44QzNeJYkL7OSm+1u9U2FfQjlF6GEPDJ+HM0HvL/dZ0Z7oVzK6Xk5OTRFYOQLxOFMYvsMN
QCCijPh13a6d66nc1bJ9trv51wGZtABYlw5mRq++LVvKNYTEAYzjQIP91T0AFJa9gW4T9us3XXg7
v/oaWKhtIqcOBjp9cdoOl6bVSazHHPK794pcSB3B72ga71q1JGgkDwiOPqBeR/YCFNUVPXvevG+J
kxIQrrM4lZfm9jlNjAKYJy2LHnmV0VmexVSpQDTFbmNqWevT5XXTq0wCzQgdk+32ElBiDEV4vd78
iUOIdiJ2LtDSy1/m5/FWWV5Bkc+IY2V+mobBiN1AdiENegw2s9VluU7RI53tkMgwuDc0eRRkXwq6
BzDLGhdTwPHvwQ1toGVSley3yT5W5KTci++rQ5awAd/kZ2rXdr8Uf8dlNSIC+R6V38jg0t8vvfNh
kR1aO/oZebVIwzu+N7EcOkOsJ5H4vgxTA84PgNPFGQi6JA/kstSusOB/9g5JDnu9lcbl8V/fcpjk
EhjKDgxHqgggIRj1EhqvD+YYYNJrKCvA6Tal6FlmDB58Ojcl+mLqAKCznLnaP7szwV0+9n3Mrgvs
T23hk1ngQLiek4M+RA9R3um/98U75uhajrckp7kBuZgx5iX88U+T9vjIMrSjrHOPK0teViDHnqjH
gmAQBoHJsqvI21/Rr4m9AWUvo+LzMkvwXWegEIeXoVEOb2vInzOv1oTfUrWnKPUIO8wC5w2VPHZe
9N4uxRVQowi9LGCBolqqlZhg6o3Fg/iJag8WAassn7zTkrpQkSaJvokBRppLS46X9NwSGlOdPmGC
EWgjp211JVxptA4GH+MWyEBWR2zFk4ksegG5CNMROijkU6QBIkbZ9unHlMYGEgYdAtjTG4qUGLeL
Hy4XIp/qxAwct2CTGahmlHy5NluJya8V5V0EZS6Fb3RtJSVhgrpwt2P/vNDytF6rpThC6BrxkGxb
gmWgXwf6fW4ui9ahmraYh58TqNoaZPd1qBbx7Apm50gMm4JI5qzEGeV+zlHZODLepBd/w8CnUunV
t7S8gpW9GDTgAzM5RN1CUAmOVAg2kCL32WnLSIF9rn1AwksIR129vGnNZJY7CS5zH0AUlG6OST+Y
tGcXy+ALtow5nq/yei9Hcs4KL538NIsYmhEfZfYJx8XbJupbh6DxnqutwiOQLDiyoiE15F3KLhV9
QeeVF0KZ+3Zeak/Ulwn0Z6x8XVsV2prSsHzMzjqt39cz+6Y78i/7DqUDXld807ayFf4K09F3AJM/
E5h4V0jLcDEOj7uJOf3AyZm9UV60UM0/A3Pp1hMsQDU2g0XZXmRHeIs448mB/OF09jDazJOP8rHI
4LMuhXNdxdla7UtD1zEgQemo1r8ymZLGKYiRpCalwWZcGsR/VDCLkHFE/RiM54hEljo3ZTq2VQe2
2r38eE/1BfYL8vJ22RFQWwOjMWPi30dvMM3004A2LSkrhyDej0q3WH7/m0iKt+E02y4Zf5aIIWs1
nQprv4WPwUX1jWzLGraZ8qSis321sbrJugHibW4b/I5YXFtaO4i1ul2EnVGM9AkWtzxDr39e/Oup
zURQsA2TYUfNKERNz/l6iBXLtPyh1NTkktwxbvtf9enQMZpoa3t7ERtzh2jahTQSYd0ZrDJek4gu
8x3Gbly0wOpV9D5JfjzlDfzAMVolmp9tEZmHzuuiV2O2ISgczdiY0KhlLZuP9DqBBT/chhbkykbP
GZlPpedZ77UQBQsxBD9mXKUbhAdLhU4yOFxtd4z8rBWlMk9TFh8m+NRMT/7LSLToxLiTcF5O6+j4
Ft3ODNwhF8AlEVAJFO0oqQw8a6/AwFmxDKLZ6k37enoW1qjQD2nTzrWN2DXLHtgfKVo2BGiUGVJf
U2A2g/62ksJjTTDnvxW3/i36YIQw1t3AHspg2YAg2BcBPADLXA+cLFWrIVyW5fiGk5BQrSeiuFUm
e+oin+6XUcShAFClvP4jVZ/GKZuK3PpoBbTuJk7p6xXDRwUZ1r+UC2uI1GecvFnse/XtB1VU/mtB
JOqkUDo7uNrpzYIOGiv7rTdIWvrP7j9QwjFUKIkz94FpUcDB/ktxFrJNQ60Q/9VeXxmq13FVFIeY
pKe7NeeH6DxaBfGP4epVrGkHd8gTYv6OHt0aSTFXbEXQRxMJQBd/DxYf5Qhn1foVH8fIPPD8Ij/z
tYpXJtNf45vf2zds7cPvXEcz3eHQFPXzA8T/Bt6rn2TLukHPEknLml/qtwCcmawVIWFKym1A5IFB
bQTOyLuCX4wggiuqxqZQ9GOqMlVQB9icFWgFnbE7Ds/OLhcrxE5NLbmOTu65vXhc+/V9ixDZyoZ1
M2xtqdZEb/7SbleUZrqbxl37ZX6VJWZxxAlMdP7+zsqK5Kt4PwDj8BX5q/++LGQ67qwP1B/msY/D
XYp6JfX5T/3/yg1VXx5ymEd1A33uEi4qW81Y0t2E7qBM68AV1wQ8lRmJahdVrLeddXWGv9Lwt3Jp
DIUIP9NwkakPmR2XNQ+ERjVv3SE+iHc4Og8ZttKQl0dmA94oTvCy1j0KIJkyPdZcj0LMbCyxA+NT
C8XPVRPW2Zqn0zABTd/EqxFrELeVxLBQxIzyVKNLJZ3WQpQEUioo5o+mtpWpj7YbWANgacXOnFmW
jEgm0AyzsmlJkiAVxiBxQDdiJ4oNiFOuGAq4S/n66q/fjvDxnRhl6lBFEFdTmqhJNeCCZdELk2Fg
j+aAsfiKKVZaSMPBmix5k0cKNwDEEOAAhvSYsvYb5GQ/72c3kOWpM700FWTzS1tZYxMf62mkVQrd
UFovnd8ao2olvxpb64HuIz3O1Td0KN3TASfNFcg2TNacN/LvkXj4YXcBBGtkXasC+eXnWbqKG9GE
k87cTrGznar3hA4TunXogP2PsRIoC8/orJbTy9rUcKI2UWBsIqoFWf7zqvfTozOyfmgWNTR2tk6V
twgPST2qD50aEPJZcz12Pm3l9Htg1307ni3zhpyhrmDzcSJlfPQYQA1fx8XXRbpNegvXjiU0juSg
qXk5bk7RqNIfiMdKNW1nc70+SKYkOUvloA/vXJGybenWYTKIrveXnQkJlbsKKXFs6XbzHnAim3GL
G13Xgb7GFQNmufA+5kvlwvzBATNEma/ucmXPwEgaXXAp3gdY47VTMDXCrzsW4y+imY2gNx6b6fzi
XQbr58WsdDMJVVhsfaWM40k0K/2Pcz5kyQr3oBaHDUrpOQhKzEFouzRWXvtPHenBJsd1TaY9QdRS
Pui5PZp99Pn5kkCAhC8PYcDp5mkISQSJW0sKunptls9elfRtxi0/tDcZG3vgSItzZY0UkYNLtpqX
KHwXR717l+SApXxgvOLEiXehhEe+JVmolfaophPrhYFtaXqUzZQxJ/JaT38alX4Iag8+/iD9Azr5
0s3OnkBoM4EH/BThgqkKSXkTfU6SjXjb9WWHK5j5vaexEYvubJYL0LrD7c4iIxhdelaOOOmPIjuE
QstwtDWIglU1NdQkwjZyyOx/TWkKp63POHOlRoB29NsFYDZ8SQj9ZEf4a9z1mpwdZk2kQ25qcQnn
WBvfYSvVMU4qTTxxkLUczhcb/UB0/atGbhXnrFpF50VOEkoRju/CDJun8kWqLNjkcix9aaiIgVhe
1y5UgBpaslOjpwFmph5Fib5fWXUS5QDSRMS0UBb2wrWACtllUNr0efFEAlASrACdW5hd2AnrM1tP
QZwmNJXaHADL0vzTr9PXcA+C+OsV/SnZeThUV7qFOoFlySfn264mEM27aD0ij7+EYzQpwOnqTRIK
dbJI/QpoI9Rvy63LPutrByWv2rzWuY7zhQpmO7uUwZqx2uqHO2HsGGZNMzyz2y6uvOezddW7kIs6
W3B9YjpvtH+Ymr3AiWmHVSxAWroOgzuyLGtKNkOfuESAG4bwodSnTA+i11VPKES1QSRBPVRUOM6v
r2MJAwf42SiL4gNs72ESNG+XSc2KAEMwlV2y5rLAhhH19gkuX1DRmL4YiMu+2Jt5H1rXLOHFFqC3
7zLPQNJilrWVUXLNfyh+QhxSwaKylY6ixF/6TQWlmPLGsiuylIPw0HbM/GTG4Th/hmuQgKjUuve9
Gc5GHiuZpL2RQs3rhlVALl+cYeea5biXBwmbYAsjHIr6or7SGDy3Obx2VOvY/96WCmm0XES/CVot
Vc0l7EgKP0tzPrCa1TOZWkifxOiaMIjgfDbv5H+H+vPzZX7mTOrq8Os+10z4dvSwzAa3dK+H61Eo
KqThdV1jhywsCphW5JK3HxrYa0QMUZomPaEbBMlHYchgbn303hi555G95BbghZi4E34Lizme76IH
MRjLfYrHEqPli6XARjEUC+iwF/ZV+fIjEwAu5tInKIyP1iorXwjEj6sUyf/+9p4qc3UkkEG0jrhE
NCHW3ate8vAqXRwIO57hzWbwvCUX4jibO9AHJ8FuXe5RXSS2HdTgpKTcW2kQrS41u7hacbj4T3e4
zuw1REfKdJHOlz/hm/Z9jMymgOQyOnREMtGWaHgKidJfupCkeEh4QZ+ZoFmUfR8QV5v+Cs0o6wjW
bOzOk7GbNQvNh3tSNKpCrGAGGpFMLg0Y4OTpSm07lK7eUP6SrxUit7zNjAr/VbhdAbfc7qO2BvvQ
xVweq9MYfm410Ku08puUlP3FlxJrPZ2y00crbws7kY+RRrvz/XUWIwniZIN7UE9ukrWwACakAKSH
v3d+cGYCU8DlSLXEuvQGfQ+FR98sbqtc5lzyyR5tv/TU1nnmf4MNgJyKLpAskvAcjS0jCbk9TdlP
sY4xmX74pV+IZyePex/0bB4qO6gRAw3yTAJB37ud8YlVJgkVbC+vxS2mviCXGKsSAgRCmMC5uD5t
MHx424/8DD7fzjOLym3l2+mju+/Dw9ujX2OltbvtE3hkHu3lGb+EE+FhmyXMY5IlRHKL5NJBGb6O
GO+LwRJmVpFREKYqY1cyBTrTWx5jqN5JJfPRzUL884gsox00UNIwfbvJg4ixbn/8uSICR1egRaI8
w+0IBlUt1rowjCtCZ6diOeH0tLP+V5j+aw0xd6scHM7I9n52sCHj2kGnnv8rhEP3Tc3VttwfH47d
XoONJ+K7+fMuhW4Xw1KkKVkyZTEVbRacLfHqHfgznEhJ/6sMwzJIbdO3d7KWlDBlKnfR2pEJSRif
zMaaMhvb6FAxqRR6d/HF9Ek1Su4aZg3RyVPoG8nDrNdbRu0kg30lxVkhZyN0HEW8bGxJjkmU1kqQ
lhvrnLHfJZOr4h8aYKeMdU1KjVArxin3MDM2qUc6ZJkb+0VBJWE0JcPlCOkxqdsIzRn9JYlVB/ph
Slf+0Vq+E4r3iLb3vcD+6KG7u6DeQstPRJX4V5UGNtKw4tlzr5Nc4cc622CgBZSyYhp7p1jrko4s
px6HvbI2SlwBibX62m875D6gSzF9lF5HSQBZiJvWR1CtDi07cJKWVqx1jSNWd0b8OyFI4R6XiAPc
a2Ed0WQyvOHAxDvIrrG6NhG2f6+zA0u1A0vzBj7wpJHDh84idDDpeqgq+sSSf1YQ80RBARuTivUh
V3CnxoJ+6dNK3aBIW/BZIwkVxBAHx8KGO5fGmqUEFP+Sf8JHJTOrHYvBZJotYG+eszg0g14vUoZo
DRfLhhjOvFzrc8XfX/DVhjyoPqn6RodTSUjqQfx2952KvYw4gvzOW2dQEQdYcQWo/D47LeB63dYY
1WTJvAhfeWt5IdJROK7T0dZBsJq/B/pgcDhUM6EbAlcOCQHo/em/slJoyAi8wX7MMtqDgRLh03QW
7cVENVoyh8719UseJcyZnyuoCzkGPCVUbRyJGoQ2n+PzrloWFCYTAwopthynm9wz1AgzQoll3o3V
6nJO/DpLpO3A6h0wL2RMG+FJB2H5dFcUQccE5xMyi/2qEGVKLiJ3ydDTBRaVYSi7uknXgWwyGwcQ
8Sy6HBp0PHDj15F99LXBklznNCkFUPYZb7vjEr8zwhl5WFjbLej7WR2UxXrJJTF32M93m+qebRU/
mFH8xPIZrmavtqsYVGtIKGkE12+PDIiFjCeKO+hYVDAFfF2ri3axtcpBYC7HhM8pQSTJ+lB3EogY
4z4peSv5/x23pU9bS26yQd/QC/azQvfEWcaGrI82DWue4ne/2XwGNDtApQ3uenTFMa07TyF1iU8e
thlDuxoRJ76QdEyLdlmBFxIQx5+Pq08a80MRsbtIjmX1KiA+z8sxyiDsm0CWhIPpGGeJ3MMr21kA
ScQfS0cYW5DB1ks1aWhUcGuDgG9WYLKbNwlaDdfOa4Fq7GNbr/S9ZPTGAluC1P9S5leDKEBZiMuY
9KfrMhztN1ZetQneU4s1sSYL6eSXt+MOIA/j9eScMOC7gBgoPId8mKFmWTGHUytobEG6DbdkHwLS
6Gr+C/2E3Kqz9G8wW3GfwRdNLPQ921qy5CfSXXngzqXsLuU6J+rp2qPgluJOJjehGdBemP4c0vbZ
ap6A0FoDBmWrQHsef0nn+I+41frGQtGauJyBPUjuhRaltZOV4oO0FJsy4iKsToKFLjDl4RnuMJO8
WrlMV44S/7t7AnRRS5iJHC9YulC8Q5PXwhr/TM+zDsdOuPrEhdDB+97WumVLeWUaTAWdYMRvvbO7
BlQxGi6RaHQTjZW32RhgS63oAFIupf3ybMZpC9zqQJlbqMuKrzfBbq4PWIQ1mJGsxp0xGkQvxyPY
SW+J/1H/PizhicYGuY6Twnjm7zuy17kJSy55xAscvg2wxfGpTWI08yOSwsbcRIb60gp6zA/iHIhw
nOOJQqSAs4Vl4UL8qdv2GKscq+KxoyilfaE5uPZUgCLDyX3tgZfNZqgTljvCcWw2zVhE+JqyT5Gy
Vvhk0DCywzuu+QQ9NVnh7Aa7zyrvgmk+3Cz8XkaBFxziEBk9pTWjqZxo/6CjQUlcwRepkC9lmzT3
cYobcJvSzB1q9Qs+8egmSxXlr9N0uLTTeKdYz6i8Zsw+okhQsMwTssWhDEcoMCnEnar98zKvF6Dr
m4NTeEdjSdD9sUEMqItUV9WnxC1TonjzqKFXnwK4qYt0SN2Rdon0iZYDAVQqhyLeU+O/EnYlC5r6
cY3ZNSGAn3Lr7Gx29hn0Y5Yi7aAXGAPmRJq1GJwwOXaWFuugUzPA59+XLKSIOWPYT5Su92AemI68
qJ1x/99dcE2paIxAontZiHpb+K3eUvZEgkwJxn3EGaFWZKcnnKfZhug2b0t+ManOB3YXew+T4cO8
ker0tAmSCYJ1lAXjZec1ElDZ6tGYmFVB8NLTeN+FblZoGbZ2Myc8pCCa72VXRi9bKNWCTUCHmDH7
MZDgpMc8K3ggo2//IoZ5X5a3f1wWm4lAWR0RSFKs8hkDXusnfI1BFAI/hgTVri4KYGsy4EAiSPKt
3LwP9O9RezDTYAgdbkW97ap9APuMDfHF7bOO3eLRRLWtAAJgBgBlfEElrmsPdYw7/QzY+Tuk6/6c
xLhRvdMJ2lTKsS8VhjKL0XNVZn+U0oRwMMVzh2Z01xGKubhq2jSWEPd5O8HM7GPhV1JJOoFMq5qk
+JLvAsLDVwNPGhWSaPugVYZXuazqvMoBw2o1ZUMLDN0cLoU28gTMBQfUlqrk4IBSoskteTCnI7nM
m89zaN7zMMSX6sY7IYwCjXen/sf8ymaLdiaTxMS8M7Tm84YCxcMNE2+owVJT+w8FIflbXyqvNefz
CPJdqcFAJZuK58blxxMUE7pXOd/hz6sLFiwSsfZf7w0Ty7wUdDnXnw1KOk0wj7a5VbGsfnREkBeE
iY5oYYPwf9LbDmASpSeOdNCTS1iiijh21Do2EWatDpcaJZcovxMfwnbr7xKH8cSRdEl7JakzV6qi
gofi0FvGoxbEj3U5Q1w78sLrvtp5mv5beu6dtngMz/ULqSZzVW8SeuCVnQnKvFjBbbUTYbhuOci1
pmtfNT9xxO/xMOV1twiEtlhVJmpDWjVmxKLQVOx3K9/i9ed1/E1t6QVVrwmq7/QlItrV8q9XPu6f
j11hU9d9K8P+k6tWkvLHMCNWpHqacZAtiP3DqQAwIHdoDbKDq/YfRRUzvGC6DpsHX0yAHjEG4rhl
JwKddqCtlnaJDRivsQkggqqxv3qSBb9Lee449whO9SkYhz1SH1rYjYwBlm9/rXTLj2GXNnlW+XeK
iOFASqrdDQNGQ3cBS6DJkzv0QPqc3HSqRplfgTam/JqR/fNPCuEp3MgWg3Zeayd1iDD95nOlN9hT
zXjKuwCJH5UdxXbYrLNkWWPeS9jROJqYnQ4hECNnlNw60oTENQ61fEVnGmRu8nf5S1AuygPuokVd
Pb+RmheAxpaLDBYuxxxRgR98hUGMKewlirx3JGhIQxvDDudyYfg5eCN2lkBDmnOw6h08JyWESvOl
7XmzGHS+z5jeGeHFGAqxqHztM0eJaHFydUs9zuPzFPQC3kvf51RVuJlkDStWQrEBP7FvfoeqArdS
tLRs/e1AuspxSzkqxuztd4FhaSJSmG3/7K/qgM9+ZkOMj9BxYqB39gFwxZ3iNyC9oXgMzP5/9gDl
PHUcujZson9zvVK43KguuIidwQzegyue3vTTgekclaRT1jIi2XeU5ACvwbK/TTNylMALeI4qy2wZ
kbEVxGjwT9rsZhzn3yl6XmaCAiEz3a2uXp0jz0wOZl/odR8YUbvcgUYcTkRZpagr4K/otxZtuypH
GcUU2bwU7KVFTllElbiNBU/iE6bqfhHsZysO7SDkKDEi+t4x1+j4maZakkAZGt+KZwiE23mm4B6w
39NqvlGuzT5IS2G1QrEEboWVXNXOF21wMunbhQcGqwBgnYHPgBvHsQPkKCHYAFrhzz3iKciCnJSt
wPI2P3zC7wTrWP7NrcQvQweXEhCYUtP6hMbeDQBIHUpReGxUG30D9doGW0hqPWzCGZc+9vLLAvgP
oRBYwqn4VAPUaawCLxUo0zg8zGBBHtQ3C2dyKmTI6jXCWdEHSw+qjJhf0+e/1auwi14kD8qSbAkf
FLBRFGDeqx7VHH5eLCarWU+r1H29kjyAW62b2M5bFy6ZZTavEKN3cz9i20x+fpnEC44W7172h2wa
F+RN2/PHNy2MsCjdfaAsLfqo5fzzRVR+R3Ro5dosmVmzlw9UGmn5DLm7jYC9W9LLluMO/2UAo27u
s/ZscVyTKTCphnFMPUhUrAJ9MgmWNCfurqT5vpYaQooqguHO29QGCOOelYMjv/7t958YRZcM9OBV
UGwZk356HBjcowyawccrMDL/1cARwtWDL1bMYdL/YN3QV9uosZVjlsZ7OvJgbcvUc6Kwp+BZ4/wh
7jjAJ/W+agzvHG5NzTqSk1Pwu4Mbb7pTxvBD9je/9fQesI0RCfCvDG+m9pBybg3c1qD18cGc9SmH
9QrfaItOqPY/Wm1xwie/qpAIdAm6t5Wjcmavh75COKfyomvI2VJFkCTyT10qGCyIDUR/JJ8RxMc0
sV6NB+guZIEHAy80C8Czg3cewuBPWNXKCRSd4+3N3alCiQwbwQejmYlLAmCM8yZ1lGKrljDl5u+x
t2wwlO+mXpz1cvYU7eeRwW2kq+/gENcP+rj4zpyuGsA1kmRbiRUXZ5tOajVccyiZ4Pkri+CKY1BR
CK9HydMfjExlC9gqK6VN8E1g7veKa57rPCy2eNbz7j7883y7VBSpiTuc8e2VKOoy2e53dEEta6bL
7S9up2Gh+4hjoYwLxSQrpT7cTK6xSKkW8ZzJQta0l4AMXMgtYdv9Cn6ECMIjAFLwAIDvXdzdEuz9
a1gQ/lBlBisPk5g1HJ79iwHqSSuUwHov/RVOoK1s5Zd9uuigGDjxIGRodbVR6wHVjTIghWG770+x
JibXgjr/HwbpPV+/GXtPdCuKavNwVM01l4FNFXg/eY9G1fpQ3MX2v25omRycbm7KAp+pcOdZq9UY
U7iIXrUYI2OphPqTRZdE3OhcPIsDWzca4KSoLO1ZBYp3aqaWFvYFoCjP0EDw6sFjiZDQ+44e3ZMQ
/61BHXcpx0pc2sm4M9R9xYcJykDdswCBl9RAK540il3j9+7kd18Wi73OFtt7nX3Zvu5Errbaf8Cl
Rb/qhyI1iiI28Q0bmevzhMKSX/jyVmzYJTY7iruaoUx0nv+j2Gg/ghOjaTf15IJurDC8pefwBP+u
FmLT3fXo6P8QHcoMJcJeSWdWbAPeLA6pSugR61/i9DeStPRDXcCjyNrvjvYA/hL3gheJTAYk6+mZ
WBvLYmQwyBipr/14NQhZsKkp3lNm3nMYTYV0DhtD9LGE1/eIDCen7IYl0kko5uk4ElVtn0DnXb5f
3vDpjXy1wkRr1ZDQljNqx5bADcU+qMtlaALf6WRVHrXYqj15NZtiVU5tfOUjCW7v4/uUtBwYiuM5
o6QGWyQflWG06D0kfZ4KFydZtKqKnFAaUKaxSTpVhCXuEBaLsYThGyAtuQaqNLamlNauX6lyrEjk
KapUYOIJgEYlm2FJH+o+O6YZf8m4fEySFHsx/oJ82cOkm4xPre26tNhYkM+Vup9AZlFiPt8OR8+v
BdkB0DJ/z4tmvnRekJEpjIMHutkq442HhKXVMTLRvBNHx05cf857GUZe5vqBgg+lmjlJ0Y1yujJO
nnVZ0XwWzhEeT0er73DHvFWS3o1aGRF8Fi843Tdi4TgGhL/Cbv8Uq1PQ1Te3wBlJDBwvp4HrKHZ2
YGajuEqKaQ0ZpmvXoEQXga5xbCxUrQxUO+th24XEipQuAH/UynqcpGWlMxa6GqBh3qEZ4lvnbG2+
K6hGX2u2dABN14evUsCYIkezUYtcuAtJzlRbkxAw23gWMZq2s7i/VoVYtgEWlQ3i41N7J3yxp97f
kTEOIYD4Op9bmRaPDujv8fFpCWUSZ2g9a6rrWDrsOZY8FxJllEyoQ8WUSl5QBaTlmFCgEfWRB5vt
U96AFPpmTXcWYc5w8sqcYRhKlQZngZrVv9tmNVmYKGgJ5zTWlT6vAS5E9PF5Llq2BH5uCi99S/Co
GIMjQ06pOYYIyeFNhkwSI6ibSEMoZ3wxRzIuRwLkGnlX0N2JL7F2aSvytsPGHk3DjbTyI6Lsbk7y
Ib81OfYu7Y3cakSagLZcTh55M55yhvZpkodKoIhwl9FUPAncQfxp83dYf78TLrpA0jtqZtyWRxDV
+GnukSeKp1eogSFoPNbmKsUkOlf/RUfJsMAs0YZR9sXWpswMZqExDhGcezAEx8cfwr5FSOLhn6V6
1xHMchDpvNzDqRWOqBsJqEjyOhLHe42g5rlPDJr4LZUDJ6bK+LPHAg+SuscW/uvPjLXVvEnx900+
b+dN6ZKvcVXjUHbQkR3SJe4iC9AVoRJveTv9FgRJkS7QfGzVVnGDWHpm1O90/qn5NqEyxDbCRfbl
iy/yugReY6kur+M/O3FKYGVem1ybm4nWlI9wVlKQt+vJRWGyO3nttWgXDCp2nP43+eakGfcXEssC
Sjcu24R0n0dc7YZfVrTybdsiu8qWVc8/8lboRqSwCZY1fpxAZXC6lIy2kRmd0sRiF+4Vng8EmPwD
zHYzxqObb3IwEWOD8CHtNa3V/yTC3BSRbrxjQ8Ew3JodJk6gW8qFYNRVm6sQ/82js4ZVlvs7UuK2
JjgjMCovIVkBfTdOYd4MpeiPcZGd3KEoLBWw934P6r/Hw3xYbNjYY2lqATUUagYJvq0dre7/DRvh
KtmCvYSBugy8hzgoLO70sKYmU3xJk68JDNLasU4FQR0uxcb0t52ARcflYMyO8ZRIv8C/xAQyGNML
B6kEX/GKunT52rXoHXDsUqgmclHKRSAVxmHQo5bwbefJvvPKqfoztfKRgevus8RDntu6C+qW6aap
8Tsr4eGzjqegeiBJjjPY3x3WMUNM72lzhYi0qHjTbs8I0qWnbDZtkkOIOv26o0pFHG09rBXZFnpB
if5N7Z+lBv/JOZkpGHc8qEBENqZPqATG+yqsixCpJy8wrGQgPrsxLLRmcKjHR1diwkFtnIOLOBrK
/b4fORQ5Dwp8BD3SIZ7wo1DFYigH/z+0S+1Z+eEy7dsYaJz2O2KSrxuduluvzJVVzlYWrv5fYSK6
p9veb+JUyWLYl5oI3drdCsHAvpJQjojr1he34ARkzDM4ASK46oMHS24HMC2yEAOp7PR0ghxr7tsE
NDRkdZdlWnVY/orXZgwTJ95WrC5gIWAkw3mo8EU9+1BygxiLcPUjYC3iIjAkbxZscRJ/Y1eyZnL1
eBtNEiLAKLCku/sQw7jOvaxrkGO+GY9wdysxvYsQkoE6R5bOTclEx/35Izn1eJrxxULD/p8KQvnX
8N74yd27e8GN4PMUAhyCyw451uXobArTbQv8SH/BQgvxtKSkdinCwhQPUPGVORAD5ZH4aNnn00R1
k1YxrWyPuXezcb1Ok3HCm8KJF/CmAK30IbaPDTVCJ7SVWIZVWRthcmBxjBO2XlP6ftN3Q6Zi+pTS
TCP/r0f5PovU7tELKtksTrq1tHAit4UyK8c/ZlxzHATfG5nBuoc1KAuIQYeSssHgRmSuAEf3mYQF
04VSLco/xN8TW/MfWEW7+0HVTqcDG8dnIybG3J+ORAV5gPJR6sSk0vHUUCLcqJ8UP2VmJWIzXEax
p2go+HqFsyj4mYXhM1LU2Me6M8oHYrfJXuQsJcI/wGDsO4qk4NVIcFMu4ylKFy6Ko60Ln7ltcI6K
TcUnmpj5jrTA3XXVdm8C0mvGTAhZdN9K393usx8pr8pc820wght3eWEtf3Wlk3/yVzotTp4oIeIv
vbMm2foZ0scmGUMXW/tuAEuUoE/ftf21kKkZTt11nbE3aW2s8Ugnc3ct8WHj5j55MtIdRoHajOlu
vyF9usAaxic9VfkXx/Xz8gjKCmzsfUFFhAmJVOIQI5xtUdiDnalcoTheD7yCIfC/HTserZcZjBZ5
Valf4f62LAQJr99smyJ/KxFDBcu+Y5JgR0sIOK1bYMLC4NP82UTmPgX6tg7V4TgA/J5BbuLzA16v
kFfjEsTHj2uBaZsMMzY7oZqvkF8IfWkRUfEQMCE/2hOQxB/xSOsJosjYg3KPpRGfg06qNzvDVGGk
8kVso2Pbcgcqi25lvHMCweSVaXX8sIiOPcrqvbZWIGIbjm/vHvp5hc6QTTkHeL/o73HQXYisr58y
7QaBgTnVseodyQjVMLE1wo8c+OlZIyaBiOpIypl9VYhS/wwENjx9lh/GuKbJTz0VDZzRyKzFrz0z
t+S69UJkJx0HdY1bErJjmGnysKAYTw6WTxueEpUPE0roo3IuMH4yiYum8jBdeQXnuW2oFKFqgZjt
Cq4m14iAsdEWsgpNo+SOMLo5QXwIgpnzCrQMzey4IAXKBn2Z9vXUb5vVfJSW6du+lbiXm3VEcd+G
u1ZS/swt970TGqB5WA5v3Fmdb3HFAbbxfeV1Ke+oIko3snbu/skg7SwewENCNt74Q4f2hdu7kCi7
SCViYivVzO20jg1Cj1OonHUOntYlOFfaNbHLdbSO04ZYcmxg+203FNclNeCZoJhaezC+v0u3dAgY
I6EaiNQkVm9BFNOboKnBL1zkiMXaZlp5DF+LgPcaxEjaeTlPM0wIAjRZL9l7jQ4qOGvKJArgaKVw
OJdAEX98KqeGNZJR/2RX5endQt76OR8sIXtRJ2aor8GtYA2TUvD2yDnl6GzA5F8QPySGJodbn2Tw
eqt2f+5Rxwwpo0QNMxanN9ppm86eptRZd7PkPJD2O2CHYT7V48utnzVCpKvMtQhH3xLkd1KMD46I
J0HCTa0yeZsv7VVi+Yc2QnYETSQiXA6PnwtMotbC4zr1ALlGTUVKvunBoAgoyTbka+vMlYlyODZZ
SxqIJlnGqsdhif3nNnWrKmviAYb64IshtB6PvXbFQB5hyegHKAEhBB+gQDhXnfVPwc85+nykfHEx
6Xv1PQsqMYwXl2Y5QrKZpPCK6FdmCsh69hAGU+OoTP5JsTco5Amwj/E2EnMpTmH8SI6cBNUdd4IX
oyY2GVeyOCtPd6/JsHPpLimuNB4BlSliRq6BifbIpb9JSfZQPvXdMWMTVtaM2ow/nIlaqyNuNy/c
1RvnregRyewYZ5+8xZhRd0BNlP/cJ82i8L2qUIFppXxtiiulUB6saFZCNjIX0/4IUPoYsVMo31MI
rkgQxIOoamgjFAyMGeOgkkWdOoiFFWWIZ0dAWlMMQnOW9SzZ4jMdc4PRNN3JGygF0eKa1rJEGqXH
wHm7lvN5CwUlYL1zjGEd/h75k8j46Bmv9Zn+xe34xnPPkJa0N5AemVm/RJvEeriPkh+NPnWopgmV
TqhJCumYMVCxD457Gm3ZBSrNrE5uH3RyWPRVPSiWLYlVQk+TWnjwVfpgnZuBYkUix8fuYyQ1H0Jb
qp8BlZ4g9UHrmpZafGqzOnxrhgv4RqhNrgsABIQaNg11XZo4o7O09nDfvkyRxZlah+/05fM6SkOc
qrQWTfw7bym7byXmUkZlowtgebkFw9Gj7LpOZOqQecr7VKn6meJoEq62duBkxUQbpK3uWyDQUPjc
OumVmVlZSx+6iYl7uJOEIWOS0JZs3jzlsoZTMMCZo2MgsqfxH+sPF4c+iyLLxBXQ+dlEAuXt7hPd
rJ+o6jksODXQAmQhiUAqoh40J2InOAWvXZKUlzRE02tsDFey0dtnEfUeO0OxvruRT1VuOHDNg52l
yZNc2YIsmPslUj8QyE71Vr+EVbILB8LRAhkzLm25qTQHgGJHSLTQf3mVgblpx0uFsfQtdnSkaH+h
xibgQD66B9Zq9Tg2XXKRpYPZmX3PtJy0YIcELKzFrfqOIPhek+Qo4i2PRvZHqUPnrrXfWZ79dtl9
vv+TMWO/uHs+pmgtLtGcQcWINJFAjUTegDrH/Y8xRBYYURWViGUUO/aADG4QQxtIwO7yF7Ewd4MG
CtV4fikzmw2X0f1jdhvks4TFwR5rhVSKQ7HJWqixxG5IptNgQ9ooXBGTTE/YxbIi5KTsDkcghy3w
1w4yG+f2gQvhEIRhwCpCLImDHirB1CwrGyyVVdfK+yiPDu5OJnVzjXe/hE/IPYxVRvJnyI1jcE3K
jE8ddEEFfod7F9kYs84bkRCKsMSAfYp51h0kG7Vc80MzBazSam9qY+nFkPw7/odPiKBAF+TxVevh
3LwoVvl88aN4JvOjY7EVS+xpoiO/TL4oXfOiLGpCBfvgonqU1DMtN7hS6iD2eOyuYUQX6a3HwzIi
Ci+iR3p3Zau65lE+kbesezFBVuuE6zgFP4TMXrcHNe62e0K8PaN4ssa3s5we1HcbiN6qKtfc+qqH
YwVSE5X2mwjSCjQcEEYKPRAb5S8XE52Hw1td+qCrtrpy2cf/F9Stosvyt3ooUvpMx9L3Zv/8sbbY
0IKQh3A3sahvli5crh+vM7ghXXOoA/iRDm4XPOinwdpzoymjlKk/ljgjNvixpevmzj09Sjpqz0bE
6RjwDECQTbVJbVB2v3gfNRFsKwxfgFRT8cYM9KYcE12S2EjLwLO1UA71/ma7Qb1pc7H3eDLBpm6F
cawh/WET7nfsr9UMQe4TxaQkz9xJl4uJkxOoS42u52997t8Qj3YAAYtBl7uPRIxdqWUpzDH6P5Jq
sRj5EsfJE0J4yQPzN+tjQ3Zg1OXXqvbRhHzAfD0opR4fDGmvMIsnRrYwj1tBkFGreYwUiaCqcxzK
iowNT/HzTtEaoxB6oXiPJ123u9TNERrtOKhvcoODOPimIb24xmTzOWc5+wyA/WngizSZLHqWd2zh
AjkNo3Sl9XTTKBg6UHaSVWBhsOho5SDDcQCm91yneGnMfwU7o2oSlPd1GmjPghYxxXecctKFw91R
/qW0XqnckkcfI2/2JvrgXx8UQefGbbLeGn/yzwAV1oS0zsnUPlfP974btCh4OIR56O4Xv/tDvspD
qaYSACeZS1kiaW/lsBbxkImB88ol8ayHPMqJFJAU1NY9+YW6QyIiwi+QSrgPC4XcxWfEfiLmjM5w
wStOxi7hC2D/FJNWLy2LvH2WBx5JkfC4Qi/tkZnSDDOm8JbGTJoBMfFpjTr57J1ME4uU/MFOspVl
qJIRVu+VL9HkCyWIGiqDXpmO0kzEF8GPRj0VvabxaOz1P1j/cT18mcaxGg1UTx+B1+Bt6exdO6vY
IdbovKHzwgHew9G2gt0EIyPKbRflhmQKrpJj18IiHyQnPP3PH8h8VJQICk70iOsPjKe1UeQaP7+8
l5XeWOiYjFhi5pMaOxnVR+ukPSaZ4AdBrFeGcTWWdRo6NdzoDNQuZfuGsVv+9aBTtiyNNobSFEPh
DJ2+GAacAdQXBayKmfNy9YfQ6qKqHGlb3M/KZukrJHlw/PKJ5aMmJt/z27BaMkRBD1vIHJHMf0Vz
nXjeeQlemqavXTEHzWxd2Zpa8oyN58dBy0mNPMgqq61klu4ycTbe8eGi2WnU/YjLUQHy9nAeJ90T
Y+Sq79W1vRvp2hYWYQ6aNIFjkNRscoyerpIKTTz0PRXG1ptCfPiJYOuNbdx0e+QqSxpdtldgdGqd
XR0OohgQj/Xlg/RhNPUTfQnTkKhuA5xUFa3iqk+DPlDSyJHj0tQkYOBBRcIK61JT1ur2YWYg1LI6
MWWuRON7ZF0GdtnIFEDfMfL2ZISTL3p2MZvaJQNew8JMXdZjS1lsvf4Now3S6Q/rMM1ZUhPq/q0a
1YT0O8h6G5WsuW8woOoB+wUJcrBzgtEM87qKEORf2F3Q8QnPyvygLNHcnLiFRUGHmXDnvrRIecxZ
hXGXqzuMyjDUShOm7hgN94QzXAB0oaWk12qvpUAH8/UfPCCjfbig3PJlyzsh5tP7szn/eSQZCv1h
86XEADK+Cyohug+CH5wU13vMPKqPtN2XNmJwp/rJbuxVuKFxTwtj+8aoIzwtlWF28QjHKIarmGag
2U/xnfS+8PMB89T5j+2Ztho/VeiQctTWtY0H91/VO6ZzXdrHoJNQOTIGTsl5w4ZpL1aCZccmGiqZ
db8X/BIAXCSEts/rSNDcV/zvuK4ABg/ly1z39kcR8oyrg68ye3zicd+NcPsx5MXKlqkAPvlDa2xm
KvOZs5CWBgpDcvGnE7ne86U3GMOZkfPJpRmIMdBcFz1kG6dqSsxCR9WA7MEPPQWhWINpDIunA6m+
8GTpS3qzGqa4vyh93VhymzM3/1IeP8avzSZgcQz60Hgehp3FEjbP4vVZfH6Er/C7b81aiLGoIK6b
sBtDnBjk7KKf26qOcn/31imSpTqTuWODtGStN0IBGhEBFCAOwCW4RS4AWwlLF0ChIMah6O1sBzQ9
AsGD2+hk8oSBHv9k3wQ8W13Qm2ikrMEiK+kWEB04tLlQNen2uMfDJtLHxjv7bBkZfiygMoIlbFtt
6p2O2vDaWfCElFReMPBznMuhXyvl198Wjt+q7pyvi5cZgvfVxWMiOziO2fl8X9mS7xkBfjd1LXnq
1Crh8oiYHsjhm98HNmXfQLY1ijgTBzpFC2v4N5QEmfzFleGOwGy5ReRo56eJT6zQvcisNrbacfGV
aSrdOAp+EIc3PBk15v9Us166ccIgnzfhx57DZPb0HS9nuG4WMKhHaYSQE5L2TMLQgYD2zBawT6ie
WMD/Gw05T6juxunPQtSVzHAkT82GddoZ/nlr0XkIa2SovLwBnJjQ0Zcw3ry3TS9SALpkpOz9TACy
/4976QY3RsyOINLWI/jYGfuL+ri0wMD2SZ02VhpIrPRZWPJ5R+lOOYb0dCpQ4xMkAY4nmoW6L9l8
RjekpAlMp+wVWCSQq+0piV91bPcFkhXh51di5zwutEmpFDBckPBAjkIFQRP+7IVr3bzin5lg9gJX
FOec3AZ/JGhflFmkZYtlEXCo9a3RbRSLH/QNWjBXcBwmjgyucizlnW+TbKVorv2xqx0JfGSTVNi4
SKHU1fhWWFrOI8pp3DJr8Nhix/1Zfy1TmnRePQd7zJVtUG98M4EC47xnxL462bldmGqXBkGjgc6U
TOcXm1Hhrb6pcS/K3vaQqE7nuq3tmSRN1nY4cUHNUbRvgfc06Hqf3UdaZWJnKpxKDcUUB2s1jz81
oyN4Igy0jL81sBBwyhX1OaTf0aJzNFk1QE4rX0W3ISPx0Gc7Kdle/Mg/dgNhZ/C/wJdWrO06hCly
vX+1QNygut7coKAcvxVgNUqnELWcSbzkbQeTz9b/pIYC60ubuygnS/3HdKOpaWiDBlQJKe2X1+76
eseacJk6gcDwk/N0yuEM8WxlU86uEve2UGtGDkAfw+OpwIIlqFODQx3GqAcjS3Q7edY32jDQweDh
rXZFfKShtgJNKQNtSS3vsegTZAfLZSuOp044usMnDpxObj8eCag7/8QpXJ4aI0w4F5/GWeD180Am
gBEyZsD8cyr2MKNhVLR1Q7w5mviePPO9aG9vUVjCfSWPgKT+ECB9XKDi3NEEjgrk2P71x7E/znHX
k14cBJN6lyuHDwf9UQE2ZLlKA270mwpg9MO2U6zykf3Ko1aCoAw9uJduKXbStfHC0Nb/pzsHnlQu
KAcVK+RzTje2GYbhy9VnFS1bv7s6LX4hmcBpeQm3rh12L+oBH7XGRIPh4qXCgGh8IVAo8ZlOYDDY
9cyOk5idNqJlkmyBgTR/dY7u0OjstI/S7yA55oic2EfOz+q35v+cg7avmF8152kmrBI/XdMHu/Ej
g3WOfnsLr0TQnAZ1lp5gFNb6eF9fYIjiXtwqhBs8Yfn0I3MHREA5alZvGAlwl4Ih6VNimaChWEzv
VUZJKN6YPKozKrKvCmvW0tvkUlZvl4HEX9fTvWbggSwzyljSPTOjFndWzG6x8CyUNBzQGXURv10m
PfdB91eWIwzSFB7IB1IuAb9MaLGbRGY77SWpk47lsMvZgxv4XyMUKKjqdGfkb911XmdnuiU6wmM2
+ihTuCcGxo/KuPHBkCEDM6V6j0PjW/oapnbZzHFBPsnaQ8bfjGwr95gy+HRjDcZUwBdOLtPWPCPI
MhNOy1HQ3G4SdydpB7aZ7PoBc/DR8WhT1mTt52bpLQKcJ0Rnn75iy3ZgpKYXIr8jxaSUbazbEFl+
DWhKwAE8uaqrd0bmE6e/J6YovqgPQYgVt5m1hRyXxy+BLl4HqjQeLEQ6nMW6Tcd0l9tsGomsYyM2
iQ4N2diiqTy6Dck+1Ef8TEBbFkIyh4PIJ91z+s5W5DEf2sZwDvWULDqxxV6u7Hxv4GCfp3KccMIF
VrJVGGLqc64wUaPwCjfBGB8159OB3BJkGl14GbWof81mzL7kNYDQ0qEFAEmIrvHVYgX/39c5Ht71
Lak5lb37WHe1pxVWybhu2LP2VY6kViJuK8HfsYnBN09+3vFIb9QTA/1GcBhmjfdurSpFJ1Db9Wpr
HCARYV8TDPnaXJVUhAex8n4uhUkF84mW/jUYgQWU6AXJ2mlmK2FWWY+cNfKcTekeMdtua8RJ26SC
kCNfMSS31fvmGsKVY4f73Ymaj7fmB5T3flv+ZVgb0RiaSwgfqUCA+zPL1/XXekAV/DEBJ8aN6FLk
ROcldEfp7iz6pThl26b0EA65hsF5BJ1R/QsduRVzDik2/lTPdMtzkKTh57B6dnrgK0i/+yFEnNIl
Kz4VRINyokGwDvYSC75Vx9uNJzkXuTrgXZLtPv6rUgfjFvGEX0qLzYezI8uSmt6c65RIug41mXhi
KVhaCIP5K9vFFYRFo+yFtTZ/WA4oGvXIGKKpEpFGb2KPze0seecU/AWC6oESCImqi/vpP6xzvja9
Fgkv61ZnANHutPRKgh5G8JNpOFxMQGarMvO8D3cGeqgnqLVZRFLhRM27F5Y6Ok76phijZyZNsCx0
nLVwF+u5v1nlwPaVxhCUBGXO0DKuUCfMrZm0+YSgZ5qgZSOkL1ZmFagxEc1Ogdqy7/ksgMkKddD8
K7WnJGwOwslSqJJktMq+QaQiukl91QQ32o1Y5tHv4OKoTHWMW4kT1EYeGcGd0YOCONYi6oYdh1pU
qP0Gx2TJ94gdiq5s8dCi1N+qOLdTvnERS7sEUoyOE5WfWA9tpqyQM3u848xX5GWqADnxOkTwoHck
FWsV0g2GEXG79Co+juPt80KsLDocAQr0FrnPi8CpVvtmWxYgW4wyBQovMT6v9NjiM05r1aYXxFAb
b8aq9yaHj3m5w6YzuGu9NtlLfiJW8uYocLm8EockBNFtX/ek0vdRFEFJM4K2G5T7M0KI6LyalM9i
TSgP4Nd1bV3Lqs3mM8IEQXaDxKpMGTcRIEx8P6leuSdYshDoJ4tlNEKJkqFGdKYyeqaM/dW1r3eK
G5sGgIp/WfIjNIPIHuXn667W8mfc0Gi/Ru5c1xi0Qw3mMlbhnSjtKFjACUIgokc+bRvqPbcMpU1j
JrhOsBoX9+Rz8M8zOKxzwjiofpyTKYIIFRVGe1OsLg+rYiXKOCloSS4YGkFbYj7ngS5dUPnrd9ol
jEW/nKjtdzEvaMwgIAjb+qj9ZUipH8r4tbWdYJQbNniScexKE3Rm8wXM6EYPYw0ilttO/aWfK0X2
wQRVrigc+MREqTFs2dcaI/5ezad6my00asuREFXVi8KROnS0++c1KDH7oNMAoQp3DlAfjdlazGIS
SQ5TjPnin81c1RGzFTNPvpFVe3iANso/2qz02ditSOWVkI7R9fg5DAI/aUwFjG4oeGe1phO8il4d
qOrL7yZC/FPhG+803rumd/k+tKEQifcyi8fFq/VYCjz1bXvBjj8YxhGHrhb7Do6RhQiCXw6zJ/RE
Q9eoTP0PpCgYoVe5f8Qkk8pjdRjk9S9opK/almHmXCQEVsjLJkmOf8ue3RA1Y4xU3+PClFFwcoXo
XLl5xWiBJqj/a4lfxfN+V09Ql3PPJLlSS4P084rMORL2Z/W26VWa5BYSThf4Cp0ocNuSMp286ue1
PosIrmVPyQPYXH6aH5dOyGDJuzJK1pELjqcQQ2YrlWKcdT5Za2FQacrC8JjeC5gkMO0j/99pkyWB
bCwdKQwN7yla5DMLitE8Ts/OiXD9mrEwZFU9U6HqZn935JNrMPmZgLq7zkD3G20ZEseuXP7gXM68
sZhg6hGLVafkGBCKJtXhzGvBOFOR3rJfV0vFvUVxGyyI8iyxwsqNYcL/cqG8Hy7UUbKJj14DD/bW
UJoEXdPKtXIBsc9dvwDr6KL13DR7VCsZYajPsSV420u+cB3NMgUDacwLSB8DhOVHa9A/ytm/TRfR
BAzac1xCmAR3/QJeVxetmwQEqPKmeSCNSsTJOCUcoGqUiCEeQSdu9g+o9O+dGTBoZI/o/ltK79cK
CqTmh6mfevaB59qlSM1IwEh4+coo8nB+uoH8kajWUxh1JAGntSkPIZ0GQC33+igIg0HnVHbX3FM4
somguDehe7SbXGc5MYjNpOfhuT/rFAzc8RiJ3xJS9g1HdOMdScEr8xHpVfZsw7CSWbQG610Yvk+Y
TYn8xqddx9hOMgG3fAdthqEz+LuqAH1su27qvFYPfIapCLS2xhuu0wz/eYcmybKT6yvkSJBPfYm5
8kq0wgNU7MvVZpYnZbmguTveTBPj7qyb5dai1j8yTTK6HMKFFkZeB/0Crqzsbf+utb1qmvR5iLBc
45XP5fvHo1sQqocU/G34OIOug9BpgJ0KKNRGDk7jjDM4vgugjkDTBSPZLqqR4zoF+CcPkn8R8m7+
bVrRvven12bbTqhZW0fqLrS5MkvclZbZ6GgSZHizPL3cQ2s0FsMbL2jk9YklKx0GvOGT2AgCALTv
hxHQBHsq1QXEwIhL/kVCAZSMULgj2DbsdBoM5+uKUYduiMHdWT4JpXyO5aL/uioPO1H4Yb6IcJBt
w604nyMwkHVxXDVBAlUwL0cQAKa5u8VZ3mZHWa1LAFod54DbO/tM5O7hSKE4HUNP1kQE/imKgTib
05RR3Al0PTBZ2uoWCsE3LuZRbajlraxH6fhSBAUuEqYSlpwmqB5pPB8N7bBqZ+fzcxFq0t30WcN8
HRuuchKEr1hPTuJejrbCnwCzdk6f2WYkwmRig2Y3h7T6tkGZBdrnu2CWcHGCaNsENXGIsM3LFVcx
5Mdj4SvCMALXUsFZWqL8RkD5nYy9pNu43RuSflJPsaOxhLExJbIKzmtPNmnK6uuBSqdSJCxf8XUW
O0uQT1zGeiMqeRk40rQyBHLZbfJ1Tlhv8vZ2wL9Z4T+M9D8DBbvJKsyowjTEc73x/4tAh26I8GKu
pixcApfLhyNjb3ooTAUOVPHeguKoCCW8KPTLKY/3NFHY9yEaPLtbdQ05O2QccRoLRmwdL85aSMs1
Xg/NsFLL+ejzKggwaLjtcPuKCKnoUZrwKqKwcioBnA2HrQlOYT4McrbLdjGn9oITEwfQDhgQu8d2
Egn+6q1sbflOktmBeNfZ9wLoJ0NB00666o1Ug//3eXNp5+lHYTonOtyQzQ4zC7bJXWlhWDWikC6x
DW3NkwljlX8G5Bj0P7LFQDKOUdF8xxUYoMvoTM9DWV9UPCShYJ/7jOz1ZO2BNFNSA4k60mYVg0qI
u+AxEuHJ4qLjb61MOM8mpsSFZdLaWGQAeY5PpFLibVuZQtUVUPiYkjy2ZyQIJ94mdq1K5kgNeIO3
3EA1zhAzWQJTz33UWkd8JINAJ5XfMkQZIdJfJ3SV+wHhcBOUNj0XWm0/L/pPQD+QHuLNjYcjN3do
x2q7a50JmgcE1d8BvetWP1CsuFhoidnNn/B/672oot4vl4oCLlg62S5eP/lecC7qyyLojVOrqvFE
E2FgV/Z0qVHV39jdBg1+m1IaAtniBQma31BAs11c2ZT3uXM69X6xOSfKCSGn7/6AvAIl4cbLRmwM
/IKJ8codwkllzgdZlAkDE2dmfc6dPsFCqdO7TZhnylsgvoliWCYKZ54eDvA1alnj74eJmbY+V/LP
CtZUSqQmVAqSlZPU9kpQxyXJSkSKvNTZlcwhXdANBOoWpXaqJnczHozxnggW63eiG9i1OgjA9Dh5
z+3hn5MIqqDCzTybcf9yVUcKJuonC4Jw5LQ+RcuPQ3Meq6bdf23PK/4MyRqTFNB3F0JyZT3AXiJR
tAjiv9i6QZsdOJMqND823ARCjDkkYv6USeNpi3C+BGgM5Ntk9fvqlv62lNU1KJXYelSORAi6UZmj
N2AE01WXPsuVm6+NJkcWjwLDwfAstDUXp9+QMtC9SYGkUIYzI2OutP1MoZfLJTZbBZNr2JUpdCLk
GMk4WRgFEizEyPQskjT1ba7IXQSRsWGNKKTNtI+PPvvIwzhlDocM42QN2rl/d+EiCg/LYAigitDl
hSjrVdoKGAzlOE3UCMe7npoKP5YgQ1AzaK2W6cqPUB/OXcsktXLQW29nHOAWl3r5DmOCzmBE66zr
o65Xbuh7llL+5PqKxmNJ9aLBfA+XaRiYtojnTwJi9jF3OoeOYfZlATYAgMBh+lwzlZa22cnUymkn
0cmOhoQ9pvKHf9GQLZI4oPaG1LrDT3ezp4O1FggNAzO/J2dYitc+KOxUevatO4Z1km3quugo9f7l
XPCI1lHQE9HPMYf1kquKRnVFT+XTSmndd7PnKrnU0vFbu8ZwXWzH6QF+M3nvsUhjKCLVHVPPk5pD
sK6vw5LMzDNJkeSztGyz+rQOjVot/siNDmU1xfyb4Vv4nGBcppYl38M1Y59LQ6v2rZz08HwRpT7K
k/EVrZXNPq0DQae5bInzNlsbECinoSFvWlG/hwPws/myDyeI5/GisLcE1nw88hlf6jwVIE4S3+VJ
d0idks6x63LShqekLYrouuIz55fHCezldZXaD6PZFXrn+U4nP0pb4/x6+9nojwWUeuXwUamNTtpL
+IZMA5VxApzXFasfpJGrAmwZKxJihKafSQy3Dy4qQ76m8CwFqdFXGMwWDd6OMdTaM69P+UFh4NTE
++DTvBINQ4ObcgbqQVr0dpBK0wnD8TQtl7w31PUAC0OW1sQyrgz3C4nX1ffwmIVburWW6hr6ssSa
lla1Il907YgI5v2T4PnoSNgLJ7ereVpqCTprFjOHAudmmq8iYBTChOI8vJv24ApxJMxT7fVy/WWo
zHb28cQotvGOT+WBr3y5VW0eUqKclMmjY3ctzm+xDJHxmaG4B9pRh5oqRPA3uThmLb9OODYicx94
Xw3d/mieMnaTGiEVNIPlVWHybCVDeGzEbH1JnASNloIamEMR/+uGPhbHj+JhS+qBkyRP4yI9tYEA
XPp5cq5NBc1SavJMqO2ihMuF0IgHh3fOaruDlqqlnD/j0xyG62S5vLuNKmSkR783QXHzSCUn3GUn
FtLh5On8IA3E34pdcvD9VPn/SN3TXM1+woSpN9M1HoRqkYIcQfwQcHj+8a3UPbHDOkNzrfHPktkJ
obrpwL0pKI46amGqFX2vqU08p4IXohk3TXEWOoKfLox7eDa4km8QU2k3177FflFLk4BIrfl5yJSc
bkYy3tOc9uhov2/OJgIH+kbt+dqpUDrwo2CpE5O2hGRaT3Ql25wMU8w5Ctr2+xkysQB+y8iRVuIJ
1UHhJ3BAO8SZLT31vE6/VIXIBo11rex85bnJOT4NpK2Vc+SyaUDm6W9oHHa5qcTlraOKT7g/8ajU
juLP29nIyjW2zLh//lgOB45jdK3ZTTXG7zmGIDyAF6dXp67YVbmOEoQ/LcKyS2UWcX8stLRkF2J0
h5UexwGXUpnjF25ssK03VOuIevSNaQOkITfD7mXfD9SLL2QM3i83LyfrPBZLQWVXzXIfZAIoYs29
zaNEwEk7EjODKYeAVVWPMNBra6vBEr08BHoxFwGKZVgxpLZPw+EItimuLzyi5BMz1EdINYXIqT5R
y6nI7bH5Wr3Bc6QfwPgXeCJ1eFPUW2KOIIXCY8+TXmWDuM0Zk3HpG82wjGiSlK1Fd8qmxptiLIV/
+0eo2Jgo3oIVrvQNJAh3GIqc1SxQxETkJTXB+H4MdwC2ECTQSadGdyuFeypwHRI2FoX/OhVwlXP3
Kn1WjhQE4jey/ykOboYc/R2ZMCGHN+pbCnJencxV4aqc+QbDYCscWLvU3SMYOFRqBmjbUtByh43I
XGjVI6NsW+n46+lDInZZNZAInBparAA8Iwf+d3UnoKt0Vu95yOddnj/yLO5gHmVRYU6nfAcWoE1g
nesD2hWv8xjGoAthvc2YwYOw4zHer2F4dr+THtZOOySYDJ5I/g43dDI3Cr2tMwBVsVjZBA8FonHF
f2gT/9cts+wwfnyQjTmittrIw0SX9fdgBHUqyIICHKTKxYuHJxoy0jHIoHa+jRXAAcHwgtEBd8tJ
dUdiaZ4Q2c913Ef2/n4Df+BCs/oTc7uDkUqWzaMo02LLHXmscZICimUmbft2ORJxI6WuO9QyRFSD
AI1Iy7vjvXRgXVEiYGswt5GKlhxl8zm565lG0AmfCFyk/DEH0ConitFrtXiM46OeG0qtaSVgxaZn
g+z3qD2g7YrC61RgzM4WRjJGzaZ658Tpz6xSyHRVeZnehAzo+/+YkiXnMIFgioL/WN96Hx804Ufl
r2OQYM23rWIZhH64wWKLXQZ2RLgcxNJZJkdT77vkmnI22e8j1ZKQL9ETuwOSM4jWO0ZVnnIGaWCc
gcGr+16WJB+zoDuDgNyD0Ik+6BcSzADmTSeYnji8VN2c9g1uWXUz3misZbVoDaGXHwIsHYknjacq
ThNFALbV4eTIoOCFMigOhpupKJ8wpvkg4VhicbVANoXoVR+0o6UzM28u3k4ngU0JOVfCa08BYbHY
mPQ1viHwv9tnBhzAFRR7Wr0F+L9bXIa80lACxljTfBmwBXEPmP/14mhe27pTR1XoAgnYgGS9f44H
dd71btWqdAIs9+RcTtNq2NR+babkCSkscStE4FnzkcY9gwrEb/468dnT0KPIoMmAo9rJfbta9O/S
nCPIgQ3w60wfd3tiOz5I7CODm8pg5F73nDnDGhfqhU33z/ld+L3AG7pP2tx3m3jfSeCxJx+wwLFF
nMXp9E114Q6i+Lh86CcAZCScXM0B30j8vApXcKtbg3uywuleg5XCzKu4sg+9XMTNHVV7UrvcLvFu
GdUw3TS7BMFdUzXxjYpkII6QdRO5MdE6dmPuZrD75SZaicyYirFImkkhTCaMFeFuBgRr5pQKp2s9
j4Iw2wqaX0uK4AMRmVBm1fW0UOywDefP5km98JMhYGpyqezgtDWWVT//VBQcjLfozpPnKJA1oov+
n1ay5EEpBaUOpnnUQkfIUwQ69iSH42O+YnNTeq1WDizzgPROzS6ijCaRf2eQgFWNcj/3Z9s/gfmA
QGCAi7D4daDQkAPmvWbSMW/nrl9IKPt9BtHxivYFzRzsgIbHH1Ovb1KA/ZyVomE/QlChRVxCbEHc
+TDdZfhghi9NvszY6ate+TjP7nzfAquDdWOVT4U82vSW2qWx/i7GmGjyhpzptxe4Kcn7JJwRONZ3
ZOEUb37DXtQIstJxkpHzPWmxgnGRRyEsGnhKz9AxLgfY1Kbs5ooi5WSGtvzA/swM1WLKWtAM5vp2
ptgNzq0NXYrTgBnkO96xFJeFhECi+qIKcficOubjNyrmHRoXbPhAjC90kBPZIscF3J1UuIlmbD94
ckLGLZVyqVU5tiYE9+DrqShUOfAkviBNLePJ1Oqj6tfHhzFBgZFFTRMLfdW4jsAjDuIeAaET3tgH
jwBKRj/Z4Uau+bhIUP+5mjieuLD2033DIqHl5v2GuujFqLNzOFb5rq+QiMwAUc8Mcc6p5ZAyTWxf
XRbAcghGp5ZxAMd0TAYHf5EJ2gVlMOjXNTz0zVtKmq5r0ittJ3W9s1YzWP2+/HNVdGKQdKqABtyP
sDUrbwtzMFsqNBnfXJSFCYFfViACcbioG+KIQmwUq3l8ssK0Y1lsEN7q29sIA0qcxFok1W3KypBV
G/ZkJnDk5SxGLBUacsbi73yWQv4VmC0VQpirfVrj0eQamw3+efUCwqA4HWS2E0YqQo70fA2rxjDX
QTKaZi/Ti7q7AcjLugrel9Dy24A7TCQ3wc1HVu4MZvR1X1+rlpR711Ctb4VsFlykdShG6mXehA1T
K4Zy7wW/RxvdZ5cBt7PfVa3bF++7YAMNSobjkwmz+b3kdZ5MXpKwsfyIwOeNXelhGfLvW28BPOp+
WzNwpm8Hwo5GvaDv0EolOjI3Sv0tWteepKyaS5A7DEJw2nTOiiwNiHCpTiSXQgOSZWGXHfR8C2DP
VvRChhkTgANFIPXpQpeKikmQo3HTDXGZdswFoSWh9V+eExW2hM3xDzfF4tXxh/3iH2QfXpVxmxNq
ZzsbW1d8YbFV3mp/A1os/z69EBUnaK2GOXGxMzsjcnUU5HcxZ1YjuP8aIsNO5GC3ETCnH5Ciq2de
/N63CCxPwTsxYuLfjIR8pLRm+53BXrB09gn+yZw0Kpap9oI/CG1PvXOME5LNoWvesJIgAiqBi5lk
JK9WHAgQQOJsN8jCHq20+PiubDKloJ+XZKY3ym6Zvy1rJiJavcNRm5Y9kqjZFwGtdMjXFEtGSJKt
MduazJ58X5u7yP4BfiR9Fviy9wwPWp9v21hp9B8oF8XdxyFebQLvv5t3i1fvTYUal3gOrFiZUL9o
4bXhxSotxhuK3LQoaUnfH6nimego7JIU41PKYcjCs158sGwG30c1ewMmaFOjRpThcLnuqsacyKw9
v9+FhU+BLQgDwgwCoHGev1PqDk6ea0Fha/mm9EsrVuYE89OkFDXU6Ev3M5u6RFu4gIeOMETVsSDy
oo6F5wuwAJYqCdg2R1/YU7h+alyNot+CXZZ2E+THKlVsQhGf8zM0iaadbvpuOLZW0SlUSMl0/oLY
e8AC9whzZCu7hdIhhqTKCuolojXyDy2M9XGnDIw1FAoN/zhrm0ulIzpBSBOLW5N6SwCxyyF7ec90
A5gibxYNMmDUEVIAtsnWBwmjFOtkIr29n+Sv2lkWpGIeQ0AA3oqrZb6Pt8SCILeR14FoXJxJohWo
6hVtI58iHQZX7Pd3Dym/5KHAYv+5rlkTOKjKC1l/MYeJT0ZIq7HhVLmGT95aZT4gl+vZFoMWJ4Fx
uRxp76ETDUeRspX68rjYlGrq7pl0sBw1JMA5sH+B3QKkQ8SDzVVXmoM1IAeCuzxSmUwKsP2evvey
4SyOzMReUqh/1iuYFRgWr4r9Uz0nmtoX5B2u/HHAB+7stai3CYlLZn72E0eYnzeXnN+pJL1vHkH3
RtlIWp3Gcmwn7JqqrROyAot5TwpFCgswtSx97iTPnh1tTmcGTHsWah/S7VrK2Ndyd9++faZGoIPE
w5hETAFf/NM4rgPfM9/6Gh8E4CMTRqkO5HaEZxRVodSVA4l99HXWFwj6iqvuLUQTmkCOddvuaexv
ogZzavXRNodmBGAAPz59wF0/jZm5FhmnC/RUVWfmx8E9gbhqfdxCjOB8cU/UpTsstwJgIaUZtLb3
2GHCzBv+Xi+0FAIajNdd85s2/TsZV86+vFGh4DubAL2MgWiOnU3VNMe1iLUEuycZ1oQcLjNB8zZz
Cdrn5mZ70zHVWoLaWKS8xT2Ru3F2xBpIGQ7AxTBhysynfeoFCRzSMU9O4ccWYatwa56o0EEwSSuU
QSr4wcBjL5Qp26dRC10UodaLRR1tBw34tPomMcFqrnYPK8XglXg21230uEO+v7eXlJmbYZ7tGpv7
WQ2Okx2gUaq6517YlTI3U3qluoll4YYRkghQRfJdbsFakQb5K2p+FGjzQ25YaZo5IoW6IGHR9uoI
0JUMWukyHhvuwNaCQSt9e7uZ3YlPWF0FKpzTBnMY4a2HsGRUsdGAzPPDeQJyYmm+5PNIFkITKNFB
obf8+1TUHQUuX9ybTYse4tB46jZGfQehIIBpkgC3YEedWfSwPfS0HM7lk4dTNkr6MJL4vV/ZcS4J
Eog+Zk+GEFNXd/mveAP3aq8t85XttK95oSE5pYsagvZl+cCd7bdpWY6J1JmGpiTbOymyKc5jnnee
YBAs0nfA4SFWw5CqyxiAGsYKc0a8faxm3jQ8/AF9gXu8OGkmfL9E2w6l73XuU/Cao8Z3JS9zGN2E
Vi9nRC2AE6agsrW0mPpmjxrXCszdN+XsGM1stw6Zxk8zoDYYCtk8VWrt6kxJSb33lQm3atDL8UEN
pvQYGjU6ycoF0hRmniXFDWpQGrn1u2XeJiHYMBkTgqqxGM8xOhYeosAwlMGHUuTvLOcD3SlCISz3
zG7Fq66Ey5QYfkC9/pAuHWInniSNWTBD9CjKbAqFqvembfCrkQeDe9yipX74wEWo64spFGQPn49w
pR30v+YRpDwKI+7lFpirAnm+AIC6DtARHqI/fJCi3NBAfq0URvfZ4seoPLFQ1DlS3GqJRskgGl4g
/KQjmiBbjwmech6J4QTFl1Kk+nDCJaVHExsChhGEAku4JZtTWkQ9K38A+q995X5lxyHwD/BVISQu
KptRZcoSAt5e/VGsKx8YaYYT6kVwAR7554t0WbB63Up2gPXhefd50fiOayaELL/hAeEqgk/PPt/q
zeVw4GlFg59JzYyekle/W0PjiVIDENo0AfdjW2yt1hTarmw4fQJ7wB5lKZru3YFlkoOS1vLhFcq9
JP7YA3G7Z/tyEkXI8QUmHLTSr69VPNKHgq9J/5Ij398W/NQweeYGRFmfiGUJYCE+kVBD8qKQ29U2
witHMBVv54a12xCh3r8UBvz1IUPcHyVhFmg6kRzCTvZEhzcyMWXlO1sbuJL1b9H3+gbt60E4+nT3
RgNqTWOVTgkebqGMxamJDWwA2G0mdUunoMS1omJi7r0yf0SF0xuqUyzfFIbzsHvVLPsGPT5EUxC6
2gwPnVO15ecYQsc4r/RheBSHPHIHgwhshwJu2wyoC+tTsQ1BmJBPK6PetWx5Ghc94Bhb4hZHWgri
OXx53OG+gtsfH9JG9x4Cabc07BmKw5eg0VWeSpFZaKNyWp77iGasl9N4+XCWTUNduS6hr8GCtRrS
bEIcOd7ZAa9z3kUYpwm14hV6dH0ZoII3RXd35ofUkTMq/yMyjeaVepF6dBttoaWCvbbwSrPx+ICT
JBCSE1WCTD2hwtr7bmXUVhxR/lOq6c8AOjfkq9x2NejXqR67jPhRhi4w1N0x9Pj5UzautiSfkKjM
VjXkhYsxrPGYhcZ1JjZpVuohTSpjCdXUlDF8T2QGdFU4TS4HZPY3+V38A95CLNWJs1504VZ3mBvC
eiVbsZViGCh8Wprd2uOvDL3hDu8d7NHtEXoeZjDt1ExP56kKiEpGIy2MxfUpqDHAlyWvyUv+vMSm
LmDat67Fl8oIzBHFPnh/Z34rCsFE6Rq6EKoWEtppS5vQ6q+OtVVzhADNVrnnjNuxsh1U+CQjQ0/+
lkgqroG348m5jOxGkRLfsm+CkIvWznwmTwbhrg2DpZGB+vfJOT3afDzsbWv3Lr5ylXPc7kNJ/0G0
th7gr1BP25xdVUR6e2CI8Vi48Nt8f+7S6argwFQHQJO89OJm42tummsukWfI7+UplZAm2Fy56mZp
6IBNgvjqey9axUB4U9Xxp6aMIgvXQb2lUCxOm+4Xu4y4F9rqv5u8an5stbUsSVJheE+mSLJwmJt0
LsVAPbqxHYfFx9f3xuO6U6V1OytE1oIsEPU8ooryBzZsTbIgT5sSL3PDn6N+gq4V+SpYffs5eIxp
wG9BWmlrWv+TB2C9SxCfcgxxrGXIV1Tk77ht7r/f0wAzy5ThxLsWvtCLLi5UZyqbcql5koH4mPVT
90w6RXmJ2qdpUDXFQvLvrty1YW30RmeOqq+RG4pb/NyoH4txt/+mZRb+Z7zvi+34svsCgv6XKUQm
yMWKAnmU2DpYqsFesSU/Q+egAWDhjLGl9Jggonga3auYnWby5V8K7Zgij1+9ET23ng+YAqjdnCt6
xgx35A/70k1M3aRkzzfTqJSXbA60VGsuO5VkiushPTKvDWdZQot7S4FTDLUl4coeElz26YoKZEvy
j1XG9UQr9/CtK7Prs45dPif25Z57pc7oCzP+8hrqqrvPfTU/yxoLWSHRX2ROBuZPhJQ3/OsvwRL9
jx5iYW+SVw4JhsgPdRgUM7j6sJDS12+sP5uH1VQlW+MpB2x/aVH4PxfJ1GJ83DJCi/Dmevm4HO1l
aBJfYe4nXjsXZVzMXVEoA7KeR7teIxTBcbbdFo84QJQ1rNAd/SsT/FyEUeWiXpF3Ucv0cuW2g75B
bzH0qvrDEqThiQeMHFCS9xmGWjNPM2MFET9tUSClRVciDteK7Zkl/ZMlsRkAgrsXlxXxEyouDvkm
jlNolebdFsMWcK57AXJGdmy/pG4ih0DC0Oew0GFXdECezF39hXNqbgX0/5Nt8u9V0cY4wCyrDz3e
MpWOvuuzEd4TY6r7E97B/SX4+ZeCwqpe3cTgej6TWrAdLjKCm8H6fb+9d2Lzy01oO6+lkFKG0TqA
hh+SKT19/d1BD4j13WFOMVaeU9y+m/gX+aNQCL2e62aXLW9RlathEbPu5FUYpkEtytuHdJqmTqLM
CdcLVM6Q8I1tRyFza4b66d7h1hifUruTrxXFezCQP5Wr84tC7yCsPCo3jxg1Mralqt0kt1ZTpJ99
ktIwU4KRwrg3ShMY6k521ks8BQytvEnX9JiYZz+Y3yzV++nXKvClRarRf3rneP/hvZ2KCYzs/JxN
kW6QM1IgLksBfDDtGR0bVY3H1ZoH9vsgHuOetjKYwIdgSlzoE6iKhizfrd6whWI8g87JBRVkyRTz
mhB9h17TTPOIr6su469dMrFmoM7f2r7OeGEnp/jCwzWnViGqkOzH1sIiV04v74HDdfi6GJceYlnM
LAD+DcNOgULS98q1rdKUjI8qri6JX0stWpNzMqomctKQLKmH8aXz4RaoVSgsdFPtOQvd42IBYfmj
RXUYDGV5qhhZaeq1px8IQJCAbhzYluXUyuqlR2ALOzcJVK42sz6kOo6nkk5eTNMCxW4e2g3m82Cv
c3taVqcN8OusDQtzU+rCqW7uB56eSQ9UYNKarlsSsk5fHrpwY8at5HpM+oFEjMVXECOSP56HZuXN
VEahmLFVZOtV6tpl1QoSRAR8tiwlTGrACWDT5bbVXRexZd23CGBZe1kvba3NPLcYVSycRPs30hZD
jFdKsSI0VWzK52yE7663XSZ8UXCaERSk4ROprqZxiqyGvwsoov2XQkkPSSDLA44b4RLrn5Y7Vr9c
q4NXm60b6E38f+9I/PoiUeuW2N7qKjh9R7unCjDXzkuiGm+Odlf4L+sfp1YxBqb5GcNzmL6R52hu
+rDwRqANkLahbdS8bvqYHH7nPxJj7k8ryC+Q7qUCSwyLvpBBfn1q1LOyhTaEPcTMnuqODnKciPcX
fjn2Mq7W1ivzGQM5nygmDZVM8st8tlUQoSHPTV+K1GdtvPUlTnRUVfBunswIcJqa6b0l5t/dFzii
bPh1chIPzvFC3lKkq4yoZ/U5yN6bpPPENtw2XpQ6+BYX/igcpnJvQPf4hdzPChWakBocDdOzoHzw
ZPG0tYF58zEqscbhzTJcr9Fr1zqK5k16bmN3fwW/U6C7zA5rlxTM6Q0VVpEyU0QPWhfkSu4Q1aB3
L73AOyV6JVn4aydkz2ZOt4OEub/UowtJ6lGlBqIQxvXtTzDf0+vlzZUJMomSSrVripjtU30e/m9S
NjjlsiKC/6N8AvoZ8pnlN0s9/Wl8qwmOLRsSiByX4hTTb80X+ZpEYEptV8snInAVDG+5N/0bxS93
z7NPfEO6g6AkhXZr3l97lrTfxamMG03OouA4fexfJjDoZRmGBvt/IVHbwl9rRduEA7tRohX3H7LK
ZOnDPDIzhzgKBaxXnHLA1R4qhNHoKMCPSRqUCjAWedKQl1p2wHOgbKHQSowmLa5UWZ0ckA86BNx9
o0FmW4p0TsroZ3MVd+bwyviGr1n2fad0F6UM+jZKLlLUi8ilDKnnuAhk2J75HVbRsh/8su51SP+d
29NP96KoKCOEBW5reffURqQmV66+gA6rZOubqJk4YejZSxaa834WVNs49DTPwrv8ZRkzv8xkIwqF
q6UTZRLE7wDtjyEH3EdbExloUkdggzIy3b/PX7GEfY7eSl8QjBTFM8Tdllv02VcJyuyxhQ0xxyg9
SbZMYc2SyPWYLHQBVTX5AoJjLjTMyr2zcC+RESwFWPc25WLYBSCYru0QmO/oBvRT8sdRRX7nzBN8
+J7BNQQhKYl/NkBdaG6f1aXbMWUoCEbd2j2K2+K/wCx1Uz9AGyNr2veZ955Hk45TQYaWUOZ9nAB+
Q4SoufIuAmMV7rjvLGw//4erfRPLZ2KwDHneoyEVPEdMDASkKfrlgVdXw7XeLdZlOdpmZQCR8Owb
aY+FKJrPYsWdKxLFjJDtVU+oMVy6MRG828gDelY/8i66qOHCapxFMQfmnkjNXOm7ot0XmqiKiKxY
0SJHXGkG87qX5nkpIyCeiptLt+shhwaGFk+nX4mmj/hg/+P5yioou/ITtp84scE2czkCEG1hXfLD
QMsOC+9dqVkF39lWx78tjHck5TOgnfKjlV/YTShU5f17B04utOG3GqRHzJ8jQ82l+RPnv1DBKNYa
IYT/X+6HTQ2fZO1CH69mFU81uBy14x6wulAmXy2TipQ5YcbF/IjuK9e8VrKmqBhLnQqLaLqRC4sG
cbmqN9XOGXdLZCmJNNv7wkP3tFv/fGW8RiJgUNZG76GwGYNwv6oxwnWd5txh/MPe/VhNd2mzvWo1
QqzGtePsYF3ki5yojHBxodo6ZJtwi2nSnKS5lGk3rJpd3xPWg3FghtsnHG6UCAuQsK0Q4Ik2cClf
/ud2HYNmAPzaxNiuxwXcbATBpt247eu//O4b0RsylVHdH+SH1S1c39QzDxUZSQZQjyZUky3VFeim
E3IEZpSO6uOX/NHMSwJpnpqOuRZninpcEY6X+ZmyiRjQCmeVS7WLH9T9MwvciNSVzJKhQHYEEiFM
3vI1/lF2lhYyehxCeQmBSq1q8LGckOaa1+1gwotegMcEir9/1hNsttjahbHx0UpAoPm7ps7mLb2s
G7Kv2H8t5JgaZvB4a7gSdPdUXQbOaBEl7zDNUSu5WwtIRNsP1fRcwIg8W7f8qxNpbmwybinqd9jd
0+vbDwmiWjBqjUusHxpIqBcEb+4IZZMLE0YHG6auLeCmJUSmE431iRWjaEaYNctUd5PpsruEJx/2
wCZpQOp++gb0ndAEkvF98wRSBbNqQDA/jUCju2JiOczku4ujLqgTEtfkx69XLk94096/hg5tlEs7
FAIV50YOeohri1IwiFsJSzYbEgGpaSabMv+vyDbcmHeGZ4a+nNetuWs9FFjZAyk8WWZHO/eoKzoL
7pYDzBW2CENHXHHmyBjxj2U36FSX/Z4jB3vDyYHQelFZHPiechboQnXjFb+u9H9YLbVYy1+ubtWS
qZwhMHzic6uUPM+5PyMxBseRRd05juIcpACKm2k+TG9uAYaipvv4twWExhBwhYxvOXEVVYW5Y17A
xxt4nxFWsyB6REfb9i6bqZzlSauY3bkJhCDoowQGloLPzbIINlOHNopSsu+3LXIUmUq+5fysa1BY
EWwtWqQWNUlk4Ab41yrniCfVDsRUS0XSw49fEQXiBAewhhhEy/acWrjS+JvQ2FNKXgotiDNT9CKh
VcCZZqJ6gt3HSJzldShXSdvj6GSJYRaybke4YJNNbpecMdsdbsZTwX9yy+bLaMy5KJZioOCoNG38
RQ7CsObY5SHpWfHfeJp7IRsQXkQVQMfTNXcexnhi26F4C36Zs292dq4dnQ0J4ETGgN7rSMkzzxyg
gizw8efo8avjKBdqRT2T0zZaSfqTz87HQs5AfMyr2Oc7YU9aWIy69DgiPzcAAUPPuMLWwpIvS7hD
r9Dl2KIH4iRR6n1QpDGGuycDHgjrNP3u24XnOAmCv3pq58KPZPf2ij7y+C8MpKtNFEUG4VLBdKZR
5L3UPq+O9OppFuDVgjxuwevwtDMv7A4HUUi9j4NIzG52rNLEHf7rZq0pWmJes+6RKXzcS5LMETu5
P7/DDWGB4DIvGNN9NLlxWN/h/NhL08mlSDhrv/NL5byluMsL1gSPxhUOs1J62ZXaMzOi1qBuUJqC
gdcAwejkMNXhzFTuEIOBV+58tOZhQS78wrEDe0EsKeB7uwwCRcrxWao5B/1YJQBlsuviqybGzzMi
HgPnEU7GiLodZ76Zumdriz5sOfSwQnhaYpwsi1TD1bjOJR8oIfPMM8a1SYjs1PMLB5OjPwZ+6z0U
CWIv7BnYn3d+PXfXBFGv7xmze5mzBt1KQNC9BfkzB6AsPI5SNg64du2eu92hXj/I286OQ5rJADz3
MSrb/DqHLGqslKHz3SNDjdEuKEFcEOU8k4CV9acRrTPS+txo45z/Q6Fumzf+BEHf0LnzHZ5FPwsj
rBAiMMiCCWK+dpQrH5MVcpl5dOI+I/ACihq34Im1FlBPgavzfBHq5JyiuMd7C8SkZGZeuiR6j2OK
zRXHqxCmPejm5VstkdGeK+5B+WPvYCOHCby/ao7eQ9knP5/3RYy3bAScYXYRZckjOeLKNV7QPrLX
FjTu16JjA5DgH52b098Mv5NI3jOAxhYFi1+Fw1CF7xeMwsceLpN29iAmgOA0FC7lxjSsFxUL2iap
3/GAZv/1eU9Z646cNyT5UhEWcoWZQvEAlgJrQk/8o0QSQc4JBc8Nbs6/MkmGqkBcY6RzwAiPhZIx
ffqCJldwIO31vWzQzZJ4pyjdYThQRaSB3yKmLTeLzVEawYK3beh096Gi/4HqHVa93NbLzy7ADobK
2DxbxZT9HbbF27wEs74CvRwXDaKB/FtLY3K9TyVTL2fjESFne5BQi5f8MWZuuQXrBwh2DSgagcIb
RRWEuNGQCAs/jxeE3tftTY09/n349RDKK/pXBz+5DGwdEGSm0WVxpxWdztPq9AT/FlWk9gcxTLqG
CsZpJFnx2truFYOa09FJqLURSYQzZhZiWvit9E9X/DScX+ZpjDwgUiC9qQWJ7RDWFWgORrccV/Id
lXUNA8yWVdZcBvcIujvTvtVjuAVVDZTEJAhtMbLwriyUxgt7cc2vbBuJS9DNp5f8inD7gWf3qImz
cLIa1/QQVsmlpOEAqDNRunbFhPTtX8pLhmD3bxzZtOWSHEuCpgAKvBLLAEtI+7zq6eq8CD1u4RS/
XllzCVfdet9BbEiRHxDtYF3Zbo4amx+eQ8UWmf1mJMnFBjapS4wxPkjFESIxtN2Ag0IGuJ6FNlVb
dSlg4tXA+lo+0LgnuEz7DNXB3oNJrFyutejEAHtm1PT6uPotHlDHkQomNyshQ40vmh/odun3TNUu
JpqIaoJpXtuuo5mOe38LKTgWfl/P53OYyjtChuQ6umBwaBWFO6cKCKoKmXpbR6FjlqehttrbadhP
TmG/bhbub9FJ6a6mFuZbETjZrY8lUylqmXi2xHWaDctj6yYrIbjYzgXynxaAfttfoU2231qkaJB4
JaqLOMvuFby5kb5LdjrGk3l17fDHWQo7TIsbRSkIQvpNtA02H+MB4jlQCwwz0H7jFPAnMobv6dVE
nWZDEh5FZwQcshwMXi4FJa6wegWUIFJ1M3o9ZPyAmnBex8U7Ab//KYnih+VOYa/UsuPYTWWwRDOY
uJT3a43Urpz3zzOcpN4QNc+9iHC1CG1z0l088AGC+Am2IIvK8xn/E+l4CO2cxgSSrpdKAcae5jv7
2QDyQ0pFXFnfd2fvwnFbm2mQ0BHxXcMB2PlD5Sc8TpE40VPxC2m6T8kYugiZMuylEWyFA49L9SQi
vMJzOS991OQEpWyq0mave7abmLBTh1XhfqeApvn0G+rLnxvogZvT/EflczGTubugpBABg6zRfT0X
xTkjfnBMsgjmO2xmoyF+0k9BIC4u9mWV6oHS7h2/w+CS5dtQxoQttc9gfdJcE7KvRTkZO/QmJNG4
OXocdfpX3kI5TEfkc1y8tNlH8HBX1HZ3OExXEV96oLux/Z73BTwgJmgzkMKyw6UV/jf2leMCGpXl
9xujKTbSeD/xklUxg7nLv3+iQJngtL345GaquJAgNSPeGrbmuw46dHDL6OptxHAiQyz+KxvdpZDr
We02unu26HJkDyrqu1RvsCtci3xueKi6/d0jx2zP1n4DQWQIT/q8+k5tkOE2HHqkERW3fDHnvIZO
Khgj9uvS7CNdgr0vgWrf/VTpg3aEgzFriSzYIlkV2etTOl06LAQoscRg/aq5Md98tlWldZx4lLAb
RNJVQTCzjcIVoi1AeFmwE1gU3CNBbToDH69EKaR1qJdzQfdfyyoAw/JPGQWJXGw/zopj9x0oHriy
MHrFGmV4tR9KlUCVvCYmlAyi3eM0SWRpzUuJVX/+ah9N5jdsP335XjGMYxr9S/vRmpYn9wef5GcT
PSr9sQnF7gKG7RwwTLizmI32z3C45P1gMqM8lm2yrJAh6Z/NeYlzxmGF7v5/lLzghsPqTN+tFWhO
gQ+p98fT9BV2hciLFvq2fl0Fw9x4EVdXAWP5YYY8N+V9QUuRXPCBAwok9rXC8w0E16d+5kle4wuz
rOon23JQ6tphGTcFwWbsAqnXL0ZyjBNC/A4DJpY1GRyfVo2E8A/uH9DKEXqli4FBfJz6AwoGL6/f
7/ISE7SUxxe2EDL7oDKJ/fOJy6aPFv7Vol/vKv35/yzZ1764Dp9iELriLqYA6upoeHTjNKs4KpwP
P3IRab1UVkfvniTzXJnSozi7OLN1d6OXXgBrAt6cqCLi8vxVpuOQEyGeOjmNC0GAfJHv3Eqy6JY2
AT2v4+qCaJGD0dpLYKNZDhHrrZf0e880HbJqhJZHeOBqCJeuHCGnjhuFRYbOONbQCzgHAPjTx/4t
v7wk9MEq9WK+waAhHDKLA43z4qeq/f4J6p9x35bjJ4x1fJrW0vE5gT6AjgDBI/z/IED1C6XufS+5
WILV8svgtgSrGmpIRanHeXVE33Ylol0mnXVbbHJeq2yr/Y2DtAuL1LyHNjKzKint+kmjnNl90+xh
tG0MMjv8A9/2092bQOa2tbPR4qgklun2qOcfd3jrnt02AncLv6GLz4zhuw59zFP6HVQv2ZfsYNAq
kJFuJqAtT2ZZb4hgJ1FGPjDyfrUprAs2DylWZnhABcI/eCYSly5q4s+r0s4pYm7J0mvKQpeba3U+
QtKVq0Tl8MyvsXmwKvS4EaDM5eQMZyRh0dtYdA3k1IneLHBRCdMjqdUlvK8ygRj9qvb8/kWjGSaa
ob8P5DSjrCvmKDXGGfW4oniUP9Y9+e061njdCdbvotj73v/wsYn4b42L0YrRvfuVmgZ/yZaURDLT
MjqjqKLNk/aXOItCyUUV7gxQqlu9RV6i0TTZyMSTaIScNHhVRNyhm/FFm8CoU6/GcEdxgpQmj3ua
rLr/kU2hxewytRgqRZ9VkR08ncu9HSeD1xQKKE5R3XP8CLsZnPXte61dMmgCFy30/C5RsB0Bw4yg
kx4ZBZIA75Te7ory+uHcdb6Ps+36RihspYQEaTpxeL1MTVX1bKEYWIqC1MlLbxaEBI3AvoZhynR9
EsQ0pwqChUuNGBvrJPtN1521bG3i4s1dWyDAh8k/nZu+EkBTdRVt0UpMnYHZQA2lzzNkhqd0KE6x
b0wdWo2BhLncItx+NIoJgVbaxg+Dfv/gEgWmPsN2iLMwMKxwDq7F9NwyF4oYwfAri4tdbYMJxpTP
1MQ7lThLhkl2ZW8KUwEmyEPnOmFJPd2TO1okd81Pd+LzeBzbChHw0Do5DM8oYUgtZnujWsKwY7vE
K6+TkUcootLPlnohhBx8Ei61Tp7KC51WHiirToe2UwhdjfWZFu2vksg/YTR0Lzm+lVeTGhlnur8a
S1NMeJgOcGNqtFLJSMCT3Z5eVhLDVDt/AYn0mKwR1WOPjsHjf2kxWx32QA7dEMO9Oczuxl9Vv7Qh
cYeBJ9RmvRYui+oXIFmNSBIUJlXuK2JchiLcQABp6MzNA3RPBzDL68n8fUYZhO+dRcPmfiJYRETM
wEv1Kk40Fg/RznBeu70lRHDhsUsX2qo7ddaR5x7LlxTVTE5WSdTtksRfs7lEMHecuzjErH7wz2fH
Jc/H5Je4c72B7mPdqyNUX6o9zJew7dsFnjGslv2/3fLaE6MuaaLFDrYXpL53rUaIwbeb5GRDWpIT
Va9X4hWDvA/TAerxIsMgrLSssFOot3OwcqFmcJEZ4JMZNw6wMAVsJwLkMtLgm3sLRQtyn/eLdzd5
lUsMT1WDta/vZAAJDAw7RI369UP4Y+5hBXvRwjDVkNQLyXfaUmKDKylnx9YWK17b7ergRVVY42eQ
/gjwEcog6eUN2Zcs5/EMTfKxmBqjyo5FEPiWnQgnD8CUBjcpMt7IUnZHa0Oz7DYCTjfurApVc3mv
/40DmlEJm0Ly37cFgPw0gGobk3n18qmxcT3Dv9C/pkikFPrHK2y7oHvmtBf4eUiv/Hte/J10nieR
grCXLUS4hAkJVNVFW3JChfA8uP5B4im9ReLUKGCsMDqriep3bzAwb7zg6qnNZ1kwL46b0QVkFrdG
dR97sZy1LxHLghOLyU3Xjrm9jUw6pJMrbRt6QxfBAiw3en2azvKK92nZWqkMX6X908qZDK/fcmhM
D9b8XPR2ygNz22imU7QLJiR1r2hLf2G3fjJqwO/1rc2ntwSsziEj1hCT0Z3QyUQfNvHZTbGCBVHr
9hyml7SWRJZ0poCikhPZ0e9Q7Eg6rch8dJP2nooic32mhnP6dbaCLjl0kRY4OZLajYcafdqztHlG
Yv7xyah667SR+Xh+plTFsqNjPuFdaZLypVQfs6itVle/pHIbOXK02NxziwMqHVuM2LyJBVHbUZ9F
qvJiVS7gJk6Po+A654pUq0EBZBHrbbwXyx5WmVp/5Xy2d2Hes/glKexkRBqjgVhBFDJwy5uJKcnf
fXLrDnmWn8X1brgB7bq7MQiEjmUFJBFamPO7CbP/uQt/zv/96acEQRPjNdsrMCml74VR0iaxIKRt
fpLVE9fJvAlM0YsUw++zSlJKToSme5yEN1R3lsZ+KA/K7RWp8PyTdan70lZodE/hsHJriQDDxIWq
0PZyTCf9dNyL9LHWaTKsvrMVIVL2AJHErGwjPQhTEGgSStElQVGXDK7M2YTkya0Z3jIjak7F+/7h
6KYK1TBCY4nGYx1wygw0SV7nxUi0cQmJjYWAMPnet4kLmPui6PtKsKtz1h6UIGMjfASOoXo6gK/3
sclM4CxefTh5Q38hbci6tNKvBTbQsQW8Gi7uWxzk5uUq1ixdscP/RwA6yZQdWvOBuT1JMe+/kS7V
SPVyZPY/5JboJ7bHbdRQfUceSs2csq51WgtrpwqJZJpJUuNZ5nR1DKEnnoVQYgQJV+CdUMXjucHU
/r7mykFF9Djhlw8QyFwjFUrvHsfNa+JlVyRNYEFgtbPlx8RTUwh8jZX8gHNBnSGtnGLN7R6zxb+6
b2iWCOqNr1CndYYWdwaf+k5CA734jF6FrXeBOUCddTSPzMOIacdMWEZtAidnSspdJ5OwLet2qlKD
HSmE4axe3hHQl5X8zmrkWWSRVqKzZ8nstnwdt+jkHf1xKXQ2/fsIphLWKOzc4g8/dChdV87MsfcY
4GgQaoQqJUd6/BfwJE5WOadlb89g3VirzsNJPrwXTvJ4Usm9DhkuNP0REzxZDNk9mo0eqyIh4AAA
q7t92DQp8VyxW9Mg+TslWWLJNuoV1sA7lshf/lnZ/iE5L982P7x4z//JLv2BQPpQ/W+qLr/G6ywm
+1tdTmjy8cabf7jkWPki1VhWWNgXWqx4XO3LChCRJZcLRejwk5n58eGp+se8t32u9F+YR5um9XBr
wa3w5TD+16l+dU6/NlG7hYEL63wHtLb1ztXXQci1btQFyaubNUIyG0g88NhjtjCmHYkIWScHWuTf
vRdqT4VFN3DLzoTuO7EcST7OWQhvdmVSSwLAtkK7QgIpP8V7LIFR6+FdUZ1Qqso1jEmFn+zmesaB
F48ojFXtg5nhzxMa6Tgfrml75/ksxvQl7ld0jRoA1izjcew1hlsbDtbkDvJDMVKltfM8cxcmqLpS
7+rGBVhNBSa1I8coA3NNwVupIZIvfkpDURrbq5SeW56w7MqacfxUsYOkJB54qKIuYz2RrxV3U/FP
XLkAIM19k2faC/Re4vqCvmXNA84E5tv43MPS5PG7qR194WK3SFFj69YPr0D463S8bopnpGP7J8d1
PiwzZ7679uUMi2iS0KjG1vIXT0M+Wy19gsf9M2p42FGN96mxpPOJ4jf9XIsPFvC/eut12mpbqxum
InT/Bv5+xTLTvSkUjcHVh8BuNYwThyinNJEqcOU0jikTpEVydRGqWae7T6cUJv2iI7nWLE3/dDeA
QmQvN3XkufxrasmCp9/OzDy0GMF9EXqYYZGl2/8L+9JYxCDPUqbUU/tsjkxIzpc83lnd/Z22c9HB
zhO/3PIEIxFzVbUlCmBof2PiJt9iSn98GcF2lgBsi2kmk8GD3GIsMchkY7/ZJiOh4wmCjnt84Dmf
xwCTOLcjMQ9AbVhPWVCQp9g1DLlNlAsjI+S7UeOkER9Yn3oRsNiy1ySNjTvautJ9wFFP6hlxE/bi
LNtVXVVh4jm6b6ZFTgACHnxz4lnwXTaUorcqfpQ7tq+/OSOTOtNXQ1iBIHttY2ngJnEaxD8ito/f
ujWnHL76bIAqpv0GTy1ZIgyjJfDbdDqA32LolQwWJGvtW1XZId4DSelSgLMoX5L3pkyNxE6KfgB0
8xyjLAnJGsa4xBjwq/9i/DI8bZ4fsO72knMbg9ZyH8oLfzyc9oOqbdfI/C2rTULaYgNlSWVXw4ZG
32Tbpgk3IQN77uX1bfG0iOruv71g5flCstGWYzjfYV4vfjUxdIDy/5sGrpq+BzasTCEIrIdkQmrB
GEt4DnBMXphAOIf6r3YGnVfe5DGd5Pq1Ocl+JGhaiKub+0q0dDj5APBktR0GKeDnF2gziVbT7hRA
CS41TcqYt7kH8NsU6R7BJYFV9/N4y3WXaH+N/USiz66w+n7ykNnhBlFxMBb78RJj9CaY/U5gtkbl
Xb50cmd61BA1UN0NekE3K+VMeyxC1nbIk0Kggel6l9w5RIUKScYpXoDoZthnPxxkcpX0kZlnL5Vn
YDRmqshmNcHquVD8lSu+ii9ek91NeYkMbx+afk76xmpMq6Ni2l6Izt8NlfU1NnQVD35O3LVuEG1d
Fz74qDTQeTg66cLrGyVajtqrCn98dlQGV3Bcc925UZmDbbbmiCDvdFZu74xipiGSuLxVsg60n2GU
rBDtuGhsrlQ28DT2DXomVrBLP0O/QdmSKDB0nNxgjWPPv6ojqWwygw8P7x2f3N6imqVv3377iVIw
1DJ3WOV74CSDqCGLvRezNu9b5YK2dPn3c0cQY/X6T5rK3tbwJAVPGTvniHuGQTCEza0rFLh35dko
teO7vHq+i0WJjjdX4mrtM9gh2/R61YTUQVWwArUBNiNtYGVwHK9/HHO/5ADsBCDAX/kRsfqBWqUP
U/lLoC/oCsvBLuq+Er/OjWdq6uzIT3SET3rQ8/Ko8QbMBqSUrkNace+YOmXyt10q56VIQyByzLTo
/j639gYWi9JRWfCbgorRpm87oQORB7ViwHSNPqPX4+JH552qLmu91542DBXv8RcAOCjbfKtOCOw8
PRdUC8AZVIRqDMqcV5XI0Kf8rJK/326dl1j1+9tVYF0kiK5yePv60HzW19wIpS2HNgKT891iJMX3
R1dmL2tOLiwf5+q+UDXOGdcSB/Lrk1PR0uHCzxBpV13XrUoQB1oWbQO2X8OyA9oCEgrIX97Cz68g
LR0Iq2hsszuZMIciWdfdfd5nXbr0EffxmrvmNh8wg816vGmUPMml0XRi8VgGrab7WXq/gNcczIm1
8hZE2ouV+O7rbOx/x0YMoBAaVWAuz1yT6IU0e5m7xLb2k4W+kjKG9Vf4ZJrsglHR9DQlJQBv1s9u
NYBkH4LcpjNktyon/DCmzyK7q9j15xPfwb5qGkwtKbqlSL1HzhkQ4fz8VEfQCVbaDsrzI9cPRes9
df6UxiTKSex2ZNM08DEyvlGOdtLH7tHQc8qunwAEMPxP+6PUOjodh0/mfvTQuRRWwRvGmGQ67Wep
M7Ht/Igd8oZuHLF8Qhk4tZ/LL1CiF/GBxTMOmVET+x3lCFyYDI6RgnTotDXP4umjRPOrgrCW6r8o
RqsY/C1Iitr7kvOm6lc99IndGQZa8snrj66c4CvANRXzIENK2SSD0bw0yCmBixsuCbnfMOWF53jI
cskKAg3OM1cF8fgKjM9H6Fe6GYYhNACJt4bh3gDtHlVuy+j0afec4RR2nyOmR2HbFZ6TI9bOnMba
Mb1mbSy5ICIVb4zYUdURtf8Wa/9rnFSjzrybw/4ET8VKsKopyQBpgbyo29tBN2snH02P4+CDUole
n1c+2L/4sPJDAQ38f/pRavUnEUFLa1ugN6ZeSPk80Kgv0ikdiW0oPZVOz6lQNwI++68RYpAW+jrM
EoPEe+5fLzozjxTX0qZam0OSeEzdpCEKvCaff36GUojXqam3Aa2XrRC+KMVNDZOJqsjvlQIgY3rN
MEUGdlwjk5FaoCauB7vn8Q+C9vIPkM/Oeh+aVpA6TES8qAxX4nEok70iid3ZDnusVbDKQhnKqsKl
wI75Bc+7yGSeFfjNy9iSKZCF+A6hx2Tze8sYgkUrUTgVihtaPFB9vqaVfKb102Pb6jYZBQuRs5RH
wX2ouJ3DGUmwFOICUuPaRHrqgcmLr9YjpYb9ZGjWjXBRBo8/NDXvqv7gGCQ0hq1Sv1eKJjk2Oz56
XfzS+AudCnern9ftkYE4ynr0YqKlY01lwGYzavConZ5eQmVbCxJp11ywxjuXDGN/CIqqUYZxGl8r
FlnAmNkhHfT9qSVXZUbBswb8nh5mIbvVa1QB2AKx+SrfpJorbFc25s0nrZVLKuw2pCCLkQtYSMsD
QfHjeLo0yKTQyRzHaN39H/6LhziNqjmfirwg+pSGI9SrxvjEftCmUtOLNij2/1c969RRNCnfvFi2
E1S0fQuU0GVUvs9QQN1DdH4BPbrrcNma7iAY8kX/qdc0kCGI01XZnSdNqzmY9CdjxdI5V/0hqmfv
an32R5Bl5fJR6ZP+nShX69fpMCzR1l898URF7a+heErqf9UCcxdvzZ7eK4/r7AGrASQV+csyTHuW
cfWzGQPRc0UnYhBnn0p5FPCGiaj7E3wIO3mjzr0UHvCBmRqSGpQ1CCi2IqwUIj/5NSsDKyLTPS1a
9Jx1pCnpMNxx8mB/SOFKTnciShUol9tWug2gKgzoWi5y1EKyaREXR2nIUyAk8rT+KH3Hv+ulWF+Q
tExj9eBshWub4QmTGY0uXIenZqGYbtMqLS/FJ/PWQIwR10Snut9lOPriot3VRKZrxnlCqXTCs4gk
acoyvVDGP+G4GoBLXwWtQpfk4lYJH5JnwkmIylYjB8YAADQwPsGugmP7eowtIrDWqKq/jEx+LyqS
w/yBfAvuSgrsVSJdkeS1ojHa8bd7NgblUobpjcuejAeQukRlI+/yxzHbNpPVVCcqlDon+QwTwC7l
lLzVtbedFcpDmfqvq1q+Mmon/l+7Z/dqLHXf5yMFa/4+NYDy/znzWGaZcu0UFUGjXuG1r0y1omPh
wwxu6ObIVXIDBNFWkEAA2V01ZvP2Pz9nIWyEExUFq/L3w/c6R/S9/uHnvrpPWsy2X6FO+bMEvDTW
3/m16RKm/LeFBvs+WeJRRwVQmjlmKzi+WFz8mF02OOQGKhU6dPgzs2dnjvQqvzSdFalFbuJDV3+H
BzAbALcbah5KFcJOEAgyHff2jHY5ukKVQDZ9Z0/iNafWQcBNuGWWifjstBYbkqsOayyPuJXzIHfL
pacy1U3B7zXC+4+9l2UYV7zRCcBfI9YcVn1aiKWGULXd3czgKcGO2TrqKtmlDcnNuUtTzdmchSkJ
OMLoZnZyBt6W3QsYUCrWFXXKjNRe5MCFb3lP0IDC/EgmPIAgCxVlVdu3TWa3/2/u+ljtUB57dn+a
THWpc7rL5dTa5jNoyMTw8e9s73CQrnoxOKfHg5QVPHFq63mzAxaVSXSQvM25T9css3He2VokFD88
g5HvRj0yA9E22MY/3AEcbKMnHf+hyqpLjCNbDdfYOCuBGYN+O5b5WrW0xKMdEcnbXJjRgM4+b1SL
K2J1ECueuig5cNw0rZxvJU/ZaHxHSUd45zFwiKZfdUJuuRluQqW8wrn0iMMHVH2AG7xMfRgj7Clx
Y0Jc8NtyPtvBexKrteFCMDEsbRZKcdJfBxThMRpEY1/gr1c5DXO01nta/p9gN1Qpkxn5RbFK0WKk
yEB46jCdWIHGRSSwVJA1A3esp/cnOfEQc1GT6Ary5iKOQmfS9P0C+BJFriZsiiapSGmJ4WS0w2fT
x8qsSPEIPk52tvraL7+UTY+nMH/T0l365wHLh4DlkdwNCcH08oSrMFojDNJBnUm0igxbhKiiPqZX
0D4LCZa7Q5nZmnfx80omHt4RheHi1jHalNrpcGhFR4icH5P6b0W5OGAYSfTIIsGEUFhiAlg8dUvj
rm87Hyb1eKB2LscIqeGTWvyi+54PkPJCBzs5krWclJrV0yVbADkjSrh49VYrP9vC3V7Lx1dKfKG0
qLI5TTakPiMcVaEVaOeluHl3iqcNDuIWRe1xLoAVTtsu/jrYE9vozvaLExp6qiDevYAqvSMsIpO6
MLZKls6C4WSTvpDu8w7QpcwlwdtBiZ1EdEScUTjTcz5VF6Ukzdij2KskmaJeIfrpLL0osYqwO2MY
qZx5jJsAh2KOTkglhbB7hQxMSwI0i38YcXWFdOokq4WUGeq0W75f38j6TQFR/EYY1EmGHT5enlhQ
TdF7fbZ1fGZhzW+XomYgxdF2JVaeMqMFDmuyL6nJVh8ba3W/OO0iTAMlVzSRvvEvs4LW9446UaxC
w2jLMQOAji1l6SFOdezeQxwDVThvUDc7f2yuTRPdsxqNFnTOz48kCBFC/cL16+r/EVI+Y8QHtPzR
iUAhSa1sWmo4aApu6wLudGKKba0N2g5l1zQaGZwxkVkwyRybhfWkM4kPSkgxwDlQtZpPNrQXezxx
M1ahcSS7gataqVud5VGRQ470gJxiyirr6L9s4ptK2FzfAJafXhyASpgoENYj9eNo6LjmiG5UsEkA
HaaV/DbgO1pLaR9hlLF6CTekZdMIBlk0D/3AFvQOtRBcs5zvkDqjm+NpSMYTnzerAY6Yg8sUWiAg
0dTEAVGk52wkm9nKtVPjADAjiTSAWc9NapzGL4SdjwAla4aed+fco0uXZAugEhSYH4ey+eZA+2oF
Mffphc7SpzaRbzTe18aO7FFB0xS2LPBor9AjIC3v2yv/BjWKFK07+kInQg9ezp3UXMmTa0IJgRP/
8uTf2xXi8fyZcuLQauy7rKUL2o0a7qCPyVgUKcr7x09EKTh8SXJALDktXffAr4zzO1/t16pvPcpC
SWKm8edyBiLMZ1BE4mzMXhuVYzfhqWK1WVjSsGrKO8eGO66psCe7W3sCz59b9NCZGh8PaHNUKMan
ks7npGPxruOhCjClBCUO/G5RW/Q/QX0hhtz5Dg1J2hBsAr5F93IOqZuku1YtNZBWPT0+HRKlPmST
oK714vUuKo5yproa+hex1b2JWcSkXvWof3Fq47App3Gs+GYcXtWrk8T10mpgIS/nKTfxnar/srDc
JftZ2kuSqJuYmRlPkrdD/p2EzGWmQAUkGyIToDklSZqGvTbfOxBSoWmy9g8WFhFaIt0pyh9PnaLZ
oD8Qugv4i+0Ubu3arnmekBKwI7FzYViudvadf3wwZQEYhJ6E/QambwGmbftapRdQq/IDqRG5TeWg
zfeF5v+QWIMyHj8EcaLBUOQIN45phOHsz7mpeWgbKfBzK+REs8lZHNJfMfOzSWRu4Fez9kle+oKM
tXxhSf1CxkmmRNS1au6qUnWqzqQFkojNBrarBcdmAziZqmrO9Mql8sA3FiMnqWe4TAs5VSSDosO1
Tg6Kiw+x7o1UdBw/bMBzXu8MqIrFK2KzueLeqmLxNqAolP23EDVWnkxNQsQ0DUEi4D+hHWLxU4uv
5CiHvzeGgVQe7b/DZsqweysU5GnkHFXhZ2QEltTQ1szMDMeveGaberjDeYYrOYLKj//EmbHDECi9
lR7s5A5d44s4MNNIxYQJGjATQb/Qt6BNMm6Z450KuPuhx1nPai4vMPptnDQAoLNFW4Vu36DfTIIa
g+HcTk729JGq0QbWqD1ZQdQBhunWcpj3NdS74E4/tH2SXbWCg9X26WDtxMX78SrKsXZ9A4wWZH0Y
/RwgILpV3p8H7jRT8leOesHWuR5xRGzoxZOsxPCYQ6aRtHcQ6VRYO50WHH+8fPCYQhIwgz0KpIuC
FEHXuQQF2ymiOpjHg1yB5sE78n6gHTpP03SdhOHx2VZuBi8eMzu/S6WZ/IR4QMuGfT5nTv853a04
AQsXfYfV+gyfaU5QwfrFFPMTwRSrwHtH+F1Ew6MLg1Z9vQ6F1MD7p0sR/hPQFbTriDNLXiNNm65C
UYC0EUzIhCUuHofnOe85P7wp3g3Lrsue3411qNJKWbx1eTyjYj+u+QlQ1O8qMbyo/0Jh4l5XKGwy
0V4kFlCvPK9sS1oCphE3xC4fn6xh1z5g7NTnWF5geNb1gluHkcIHL8nLioxSBe/Nqxt6ju4GwbmY
kT+avxdzKeUutArS4Hd9fw8mHRzVs+/qjYCbsDdhE8I3B7WXxMQy7+9ERDUMH+7lF5I+Zy+nf4lX
DOU0F3iCATHz3EiJW/mRXb2MmH9j20bUSAydU6BbhhGBZsjibhyNN31gvZE6uT+97H6HaE8ST1JQ
V32JWyZ+/6i4SzSs99XvCfcXk7vRjPjHdZk7VdcaWDN9Ft2HjqSCxGWmYuH1PLVfv5cLQGFFIadw
ZvH2/0GwSKc67tG/9y7AWt5ZT08TilJ70Ad88j0LRun/ElEIuN8NnDMdQ3aAVJ1wbiPMmLMbtPta
CyYZELZFy6neKY/OYe+ThYYGfNwuX8aHx00nB5XLHeZCCZCn4OKSCl6oCrcvDOadsarxfeSuVoVu
oG2lNNfm8rWcAMA3ZIdLLMvAyRZxgWjseTLBmzG9dlrlRLm1p8U1COAiBThIBE/lruaDdnSHVyiE
FBoxJhbKqdIEO0QoWb/S1RdUu6dtFuomQqYR/VEf1d6C0sgYm1iDbcFQTw+pMfumuXFZJmXMgKeX
N/EqwzFtuOQwcFZCjweCJ0ldWgk5ZgPUtpLrr0dn7LJ1F7nSRiuvk9WWW+WHIKlEReLwpPewpxO4
M4uoh//xaggJ/uUeEcWANoMsd+qI5d6IQKc/X9WETZ97NGuUFj3dUu3/4CiX/3x0dN2GJmuzS/jj
6KHGGVqNzscEadrXl+1NKslQyDFY812MAk4049cNRG+wHw0sPO42Mh0EOQyGkB4QaI1UXZZjSKGN
PHpbmZTwfXR7qdjIaVnlWS9tHGVTkv3jyv1TvBKoaSqYw3awjYLWVeD/ke2mzAjyefJ+B7TBijJE
X3gWeIsdVbU+yvUKzdE00DiDcfMX4lAYNzeZATDehjfgMWa21DilVR12jvow36tFNNnyvadV0uSv
crP5p552PsdRIMqDe9MUaMKLL5YRC3BM2l2MVT9ty1mOh5wlHmjIoWpND1fcrboyRWoaGg0QHyx2
Q0KThpJcvis/HdHcPWYkZNmwwbP25CYc/LrS2VXm5Y/IwKfNVQs6VHb2OnaHKGYHvapHIyjQTxZN
NMgIyhiHsohe3kRi9sydX8JsLhDLAvCK61zCcrjMpLrY9Fih6m4xrV7xD1MDONA8aknCT02GFvYN
SVeTlpP9XYNgDCJq5hRDo7Pf3d/iB/oZ3F10d0NURNnhryq5VBn0cSzWtI8PP5XCF3Hq/OlFM33W
PlHKsgWZsVgEBbDZFnwi/4NqXljJlzTSYCdWN5OsOCaIiBM1i7ttRXRoIXFCvMdolXBO2stMnBoU
GZL5XrX1zdMOwxwnDjkCDCzQxT5Y54gFbRFOeHlxCx7h0E4BIC/YRNGOKvZjJdM/Opf5szuCWe4z
EouLUDQ31Tc2BpAhLwe9EvJbPnIXzEp/sozK1XtcV5Zns8M1ASBP/tJlmNOmvSxt5GvU/6kFo0l6
2i/1W8mUWpqroY5gMLQD0ys/G1tjqPJZQubgtyqa1VBnXX0hQqtLvR2tNs7upT+5ZrLBPXzo4g4g
LeYwqSQjBLdZTTHj/LRV/lA3sJr3OmayKyuvlK8CNkCnJUqq2jo7Tdi4KJgM/JAckpkpDFwN3P51
NLzGD8VnCVNdfGIeYgSRuFLMmsXhqjZlUK1qpDCNeQZHhnf27ICWUZGe225H0E9sr2LBbwVhW0IJ
KM3npmVbuCnadY+uUeIw2EC9mCehrRDPgZ7ktSxbPzEDtyPy3CCtHkOtUV289GR/WCkd0bSXzTkd
90wtulItt8mFsbXMSl9ItiHc1x5oN+F9V45Ch8dkdYPfrxvatEsstWGB+diXh/0HzGXVkgVraiLO
Ynf8a6PMxU9vcjAw9QJqOg8YAaTEbNob5TRfhi4uOjX+6NDaYsaA9anuJN4Vtdo0DHMhU4n+r5ID
LuA3m+CP6EM2AuEVWGSKG/ZN8EF6T1LT21JNrUC6hXjzgx64oZP7tI+J4om6MTs4ilo2WA00lMC6
bFy20u0A07h0Imgf705gimby0yzzP6/Q7+/q7H9cUS5u6DZOSNE9AX0GqaeYzdEc3+ljg2SqXUoM
0vG8ne3c898UiXRzj7/VmQOAPRqhmjz70+jrp8okpjoKSJ2Zz29ztPDb5Tbo7VEv8QpjqFLsrMgl
PeP9XoxEI27xZYLz/vyYaI+JxxaZBc3gMEtxFral8ydLJhqR70RsP9ynwS1a5SxDC+JsucBYmqNw
9ciOE3NrOTkd8mzWoJKYweGtFKi2dbHvUCVXy+b4gIKibUwKk/H7o3pFsj5ifAeFqyz3F5uwYF5R
Zo6f89vkKL49wFHCgx43EZ++NAvI5iPZJ1r8TDgVKDGT5Mbwr2ini03baof9n4iunBT2lwcyolVI
pLHUkVB+TLFY5Rup4KDhHYsIBTfe8QWGRzBGkVHMzuoNHK/X6S1DQscR67o6FCm7Px8DRhYBrI/U
GqxmzGREIIthRBxxDSmHpFTJxBj7T4soqApnpT1DZG/5roiOFMVvis2Wpz3AehAqsKEg2AHkP7XB
npjOnhnrL6FRtMtL/OymRJAA/5BOUThDxjEPz1UdwIlR4ismZa6hz9x67UHswEMR8SmZfxzjxPzd
pLrcRplM7XyhDXGmjdPwSqq66WCdbMUsMPFERPSSHkd0uxco9ajGu+47o7jxK3CzHH+SWt3fnrQ8
hOo5qwAa+yrv3iEVUeZbAKa8EpdSkEjZ6rPxHIa5nIsmdSaIKDy3l1bKAQJ0O3huWk2Tt+ZEoe3o
ffIvZxG+OGMLEg8LwABpUYi8iucgoKqL7xtYGtfMve5zH5Mm+K3k+TLC+LCGgW7BEDd0eEkPxxKJ
zpUsMslmf2uJvj3HsxMVcJ2N5Gl2p3nS4Fh/j2BgeNeEDiuibzbsFlpbCz7mUojMhrZ4S39tC0O8
7ll9p3z1ItfyqkMAnw9Noa77e9tDZSjrbG/5OHWe5sPIgXlXFSKer3z/0HLG50evwEu4A/PkEFYb
s5hkuRXTzGMjfY9ypdWD5/tTA3FO3muRXfrjDUsFrDkIwwbJ0T2jDIBc+OCm7tjZvwQTFDtsEMr3
zQFpye2XCKIS5Cp9vB6jKMs5plxgerXwWz/712bALYRlFxgo8IjRYNGd10VmNmneaigI/haWa7yq
Aot3gVwxWWEzjWdJfz+wjJ2segZgmcbx7FR447Nh4Bgfc/WX24TqdWzGdQOE6cY5f3FxoBklQ7R5
UidgN2Ot6RbdP9h7DpOuCx/bHfZizP7BUj4505NOXzfRo2MFsmD1T3vBPSZ69j8xGYfD0gRjPULP
eYf/B9anTJeL3Hfi4rfGqhXdCejMShDDi8xIM270utZ0xzg7q+IPVpgHIgbaQ4+iapbGcONzWtsx
wF3SXtqKEz+/TjwH2S/ePokai3vlaA/qd0kX0yrMwqd8tjrfhBAqhdgo2HS6kGWIzPrwch6+StfA
TdV6FOW4uYbuefo7ds3iuTya3jaI7I+2fK2dYLO4qxacgiCQ1cUnsA6TpgHx2ZZi98J1jpwyCLSQ
SOSXAtW1FAJuJ+POIIYoF9FLFySuMtSOCfsgQ9WHAsqxEHJsOqb27QXffYi4/9D/CGx9ozEfmO5b
sgwD15g1PSZsOJ+9qQLXUrT0fMHrRqicxhsGEN18M/CljHmCdMr3wwXpbT13NUpcndlhf/Ri8uIK
bn75E9ubSpXa4bCUVnVryvnOfRNv4gj2IY6oiHObnHNsh3Gva9ck5rG8VY+NYTM2BvRF6DbkXHZh
yIpdIdEQgXiEevonay5ug9RIncW8N2O7rcfZqKlW2ebZN/F43gqMxzlce9W53BdAclxXvHJBXZSj
xC1zFDWPN38QtEhx0lN46FhfB7G/XgRZOVjx4z1hQ+aXoZZgjrRrQNmWtjo8uJBzzUCl7PU7PnKu
prgBGwDuDm4ZPnleit25ovFyJ776YU8zzqUzd0Lw9LnZFd+eIxdYwvTL8plkgByEIKJT0V3yKnih
fpB0S1Vp8kG9rzJn/ZwazEUEFl++o46H4mb+MJf9ZCjzSTBsBAtmLLJTAJdmCflXEg5cpOlF2uIG
DGf7G4Ahn9Zl7tCkyy1upKNRJpzlM3vU5wibYthCGz+hxAdt5cTmlKy+V2jqRjwLqyoeUVyPpnkG
Q+5Xrcjif9n1318z4EBVxZckg6uosIEv+wQnM+fgbx6l61HI7LCvzJMAj+tSqWxdulPtO7J6p0Yc
sHcs5OCOSs2v7KhvbN+m1/H2Iyhctwo9xfIX4FoZuRqJ3L7Bz+Vz3eYKSqWfoh3DgIKEfa1SkLr2
x4yWUvZZX9ic+EILEd7t74tBKn/TUQP4NcNsgHN3Ebo7+Pe5zgRc0+57DwWnSTVsiPRW47evmWzL
Y6OISv9QwIytoMSiOsxAhEOcxycAvyAUILicjnsXc4ht7eUlxE6BS8liUk7QPpR7T2btfvNkmsd1
AiLKIa9O0sy0N/UmonTMbHZQeymaVxUWXbXLukSOEofQW9OWnn0ldolQ54I2ALBs/3AUSakXREq2
oHl/nUEYU4c04W+292nkTAosikKxDGQKxPmxNsHy7NIe1MNaVMtqId+vUMzhLzDJ31JWsoRAqqzm
rfglolOJeYNHUathk6TDlxmtMEOlrncNwwB5msqvTHUs6+rSB1hmvdZlDyHD8ixqT3+F+V5dq3RA
kGQa0kYJMlt6bl92lRionPp4TKXAPL3O8FAe/VJFR7TgGUd3pNYeCgpjoSRDEyKaD9ItyAJvz0In
7udcOOmSrIRoLot1WBdpPqurk539KG30VSz/jlyb1Wde2qKdGl4zcBSqNUB67x5sjIsCUXIQY9E+
MI4Jq7e3GpBagr72AGlecWFqwb00/AFGoCUp6//DTBKtBmK0poY+fKuZmpgoVcndn9GiQbYdzYTk
Z0ZskfOPgCT65RE5S2R35yu805dbVwbLzDYguEM50WihTJ5HRJiagaV3DOIPxB/kxOktE1HUOl8h
BUX4r7xs02Wpm1oMVFVi9i3dbTmWsqgqQ/XzlP+I9ECwb8p4zUzo2C5+pI3bFR0eAnM5CgW9awB5
K32xOpRK5/aJxGzB8BYA5K0EQTsPy9RKq678bczQBlRvEs/37Da8PHqWFWtuoqSvA7FZGkf+UWcR
a7JgFPIczv4ecOZMTgC3tmb3wPbShIQvLUJtxPinxetGEO2g3bwDIOyNAIIHZt3QYHF98rXTv0Qw
L1+MZ2g4dUjpA3rs6H0NPF3bMfa7Vw9fCPGkWbAyl/RYizYs28Br+9EoM3ZXrXVzDGQE3b98rqQ4
nMc9qgDgEx3306IzmBXP7xu7hjpZsVPyGhMCf4320dh++4y9xiaRvm+5orVdEAZq5xp8YNxDbAzT
ehbhH8Xfu0BevcxKeB7R6izC9fIYkhCrVuA72ZvZtMrrDSkat9SaGOiVccbZMNt9kKLAGh8+NRmd
/g6hpfbLvaWzksPfz2gmJtygoFM4j4OkiVm5ySyDCKcU4jMWZVM9j28XxDBfQnJXP3euNmPOq8Xc
deDDN4aX58OgzaWuCZUzeYyeK34Aq+gTBWtVG9qS7k5uspBX69vr8zfg+vNA5STfs+86OyYilRAL
QzM3Vso8GFitXaPAYyyzlSegqnGHfVBIeoo1gZZUpJTY1GazZ1GGUtqTCD4lJwkkhEPnkPZHrRCP
q3sjWYKAiGTFcMf/1g3rDGsV3Rvvl7CaAAQ5dWEBaf4YTjSTGPi+JKO8aj1/27fiznMrYEPX1Rg4
Mac6nhQze4nu9ipzmKwqbkffyQGd1ebeC2v4uKBV/AyBAFCC6C4/OgVvecO59cl3txF74NLehW9h
Sg4cf5MU9G8uO52lkFmIMW9LmXqLR3C4sdhVAesg6ap+ZXUElQx9wEAp5oS8vHAA19eemhyhBjw5
3CLuOY1KtvVQObOzP16YjK0Ppik3lW5/t1ogrI2yg1N4CnGZYdElymG5DrDGWGonuxsl3weL6cE8
xSfk8HXQqOLDifAAoTU3EGJAIcYkUUW4ZWMB5FrWt3wEF+H6KfAGc7FNUACqffP5yfI3fI9CeAAX
J8SBtATvSncxgT4G4pX0G1UzQTJ1HWzSeFGwRJUlE/0uu8BVNbnWXdoh8rwCJWyyYI6/F2dFfaou
k8WU2F3wjJUWlKzM1QCQ5+6S0A6VfAbYU1PWMx0FqZ5NuGb96jgAC2hVd0U+9Vfo7kSc7fG+coay
xxTndb7S5Ou/ZG0213dCOg19VXLYLoILdsPXYjfd8hJ4CtRyCdXuOt9G4kzLeGPcvnWLZk0l+aqH
PQibvaBmfiyUOw4JewzST0Ld06kPCpWlnpyfdOKndNDE6WwlxeMNNg77Ly6c8L9gk+HTRA/LbxuV
Ic5affAlCrDkldbJNktMpoMKNikGVWhXXoam1e5xth10JoPxzb0XiTdRsRHmgdglD5KViGkha9Eu
4TShh8m/r4k2YU2NALsrp/fna9tCgswhwzUOr4bqwMKlCFrulnyC2glYWH/pNg7uX7slX6y79b1C
CD3YKk8ChsjcE1hVsvhGphx+jcv2NgwyrBhiqA7sokSxtseMAcjl1b5U9Qlq1sZKvxPIoyuc8abw
v5R9Pwg6ka7mNn0TvHaIhOevinttY1GXCjMrjd0UAsJ3Kvry9GhKenW/lumDq9VsYz2nGwSEm7g8
rfHC4q2rVh0MiMRkexLLcTYDJffrb/GfP5FEN5XqZDBB85Fvj3FFhaRkWAiPUIkn2mntHHQFiBo1
Y6z9HXEjLdgB1kGRAo5vFJVTbM6sgGBVNOLZkvo3Cy/6Q4jq86ImfO2TyvOpnWzIP45pXHmEDOMK
gS5s8hrvMZRv4L36wkFMzvm9CBhOhDwirw4QG1msKPplPCsfqCZvPyy9Jl5bof5fJ6qFV4Y9vWGo
uZMQbK0sy9K5oeWxfZu7zO5VEBTTL5jGncHvlWm2zzeS37DkqZAcF3VntvNQEu8zvJ1DWuqoivfP
f2arCfY7QaHElSUbg4QYtg1yDBH3+K6cfR0kMnizatl8+VUyJYdSX5Jt18A1i8ONy7zvDs4ra6rm
I2JjCGGTbaLrJghHL57RMG/EDXIgL+4gYm1jhwE69zJB/L8rEHT5YQKSZ6lPFuW94VOujdy4D4GL
PBPMr6AisjWV1IBiMcDlpJ3wcjM7PVrrYsdarimJHgGNkLsuPhixQLD4QM738U9BFgxSDn4pVvF2
aNTMqji+O58isZLXB60Crl5lyoA4PxmyWATC2yMvtNQrNfketaNfSXDFXVgNwsRaYqMmfQbT+wao
iZ2W6ACmZEJ1u9RC4dKdJmlljkSs2O6XgHTpG+7wu9pi95MjF36pQjxyh059oOVbSzwx1GGj5bnJ
YYVI/ITMIiI9YuKpTQerxj3QtC/eMgLgDVvzXoustRFKlGaWBm7JE8JaO0NHCh96TaMWpvSfzcdU
xEYLp7WYTka9N/rmr/wKsS3/01/q7wnXsZNZEUtZMe7MVVPwHS9TT7mbiOWG23LA2F7/1v7WKk9+
DQl8Lk0gEhn4dXxGL9jpWcoYWYwsECmlHpPpRUS67w84r3UD0z4yc63Js4eVuQOhRcAX96utT+zI
JCUEtN6K7eIIk+N/kyBDJlslwkpJrgBriURFN/f/5zIbiKg0+UUn+q+628uMEPehpWmJDbzCSMQU
5rgV8ub1ihf4lFW5dDqS+i4gfidlnlCBQtz/wf0JLoueqSnzmQlC9lvnIgcsYPBLfbDnNZdh66qm
JwTfBo/n9tUC2+UuwnMNC0UdVFf8uHwt3tBTuca/gIB+epv/KvlJuL9hMWYEztSmi/8SP4BWy0eO
IFWm4CcBJ54gcz3/IoF7OnhRJ14jk4xK9r22xoMOvppCcHsefaQnc59mEnvtfM7/CQOFOhiEHQYN
+v7rQTpNluUwpfNUOJMluxQg8KSZutXMNkCZ+iv+iUgPGuGgnF+v3n7TiaHN5OPhacswo88bA7Lr
ySe556Mj5XO3spG7TleLJDn7K/uLh0Ym4JkjvYLwsiXATTCfKVO+QmSsVXx6qhQaa/k+ol4uXeCZ
Uc1nIlUOMq5UnBLj3HptR4U+jcfboWJjACxq7F2qS2C9Wot8rBM2yLfsQlWvO1F0Qs3pFUjXBcNH
39EYXHRFhXnrbLzB1NjKntiIgIQXbI1ysnxtPoBuqSJgi/MN0kFHhXAkwXqWiRv4B508eYg5/ncn
Cv60/ZUQtiyCnMMOPjSGZBtLyKZ94tByTnH9GorGZV6XkaZ/eHE6QrHEHsg3y9CNXfyzVgcdbo+8
04R/0arMHMnG+z91ToI2LkEStloxkjUD/9pPP4wv7QC/Rx7g4XeKUmWwcqnuSe2ubzQIT7JfcB9d
zfXWFQgYaxpjbPLwCKsuRUYjAtkVtLjf/J4WA8gkSBsIZ9ZobHGRBBQBYd7dBs8dPJgFFn5gF935
mXqpW5ql44udGeID/hk5u8iGVnLrzYDvLMPz0NsYzzgcjfFU6OaP/bbtlzEI4fS4xOOENP8wdAJk
oxDIz7eQjaJ2HDMT3q2DR2Rg56fAJKb4CO6IM0im6hYe5UgLzY43QZDvwSY6EYQgXht6UIpTazzO
Zum09LsHMP1yblgUCEE9z/r8HhBB8Sx9pnD//cvaIT71y10QvT/WHm/CIos259ndu/5PRri9wKgF
vBJUhgzEYT1fM/aWVkX2E2sjnwsRghEm0+B32eHud1ARuDnQ9a/L8dy5qkJqHS5vvqDbjXc41orU
gdJOX7DN78ml+SRmwCDv0jW9UI6Qd/gn9ikGqI+oK5o3b4L1frz4lvG4lp0I4FBhf6m+aePox3pS
akoI9/6TdkONjk0agdpQYYzCESgV0UKUu0KFfIxH289gSozrgiEzm4cCDOm/pHx1CbpPjQXvRuyz
xh0ftc0hiFtNbLj/Rq+W59UhZqE2now7P2clFUHnKYg0Hgo/Jojwz1b/GGQThPNlCio+lhtbD4B5
z697HE1QdfavMKTxqNVVxJI/Rvvn5ZUxCLncXrryLDeOhETlqOAZz8obncASadmPJ4g436fWw86c
/m2gf4Kya4C5vBxSFiNDkjDyznEZOEz3Yg3Arq7uhXjsQ/fh2gU2Y9CJpJIz5wnBIrBzBShNHueK
mx//nDAf/ZALS3Xonj8w5JZgxdXzNSCz6WiC7qg++qXT8lF2S9qNQ8SUGkLw9vXu0A8Ob2ztTu+T
DyXkYV7WDv9I1YUUDq+UvjBLzifC3zss9e13Sp6UjPPwDeYotulauhb7e70c4oY4BhGo5OHgHbKl
J255kU9wlaHQSNBVrsd3OiPvxVH6hTseYNs0Xms+BpGBKzAiUA2qhCDvRtgkXvxpDmG0aXKq6F2a
GvVikQ6jdfako1wyQw23mmS6Pxq94y+pEFWxrJQUGH1Xoh5Gv8yQ6T722+xpw/n4AD6kaaR4oC6L
dyYOj6Q6cTwI/BnNkBLYBB1KD60TjlqGxOe0MIY+hprMz4Xvj68rmtGKawzg2fCkHxJQUjG1H56n
mz73Pp6krQK3cH0I5KFdgTqqfSJXsfIGrt/rhabI0IJsLCwYhQUdlAw4h9gfkhY0EuDP5Y+CQmSw
pHoX42GPwIDkXYUtQegmK3Adjz7OKjJla0weWp/V8vdsSfD4tOgbfRQxhg0oKsBj51UaOPB7lX9P
4M7CZG3HxSks01Sjkvm0kXKuAsD+FO59HvL3xiq5BqrDGvjebjEk116QF0HEbKJuI5fWqmN9RPZH
Q4kGwlH8SdEvBYedpwMS3vxS0nXUZUZQxJz5O4uDjoDRgIwFBb4JkK0na1b8Gfge/cme83Q8mQFO
4Pwni9Eo0UGrlc64TQmlG8ZpEE+AI8wASjzIRPutMh8bVMrJw/IjnicaJR9MMOgZRENSwV628A81
f5UlqUA3VNcePWMD7y+6R0ms22ZP2Yk0N7M1h98QUFR2rgWO0knsVobgOytBkE1U/7vlJB7GRF/O
0HhU18sttOR8Cq/1hM9a2zRLYRQoF6eTfEJcN28omVMvVAWpZx7kQ62HxLrWPx/+mLanoPU+PgNc
mWdP1POuzOG6DbBlyr7wJc+Lm9nJeotBr4RZKU5Shzi8eMGri3drPONg+jHB0V0a2XNwwtP7nBfn
L/78Ki+6lYO1QHN0XrFy/BJBmrFvdYEHQQHi5Ra3ShitfPScbvpKCsHnyajHd0HLo9vpukKmvCw2
MQV1aRAe9mnK6cmrAyujMIX8lNbRykOaeAijfwcc52qEw9uv0l5vhI9rHLd6EAMLEK69R/yxF+pw
sFPy6lOTTVmgJqEK0N837YX72qwXs1GvU3I5hPdiMLxl2CECDaC8yw5VfxPqp+jVWDWMBrF+ozPq
Uo3TvS+uwZBnSKvpgK7QbkaqkqRaA2EoDZtZp0A3okrTsy+3ypKs4DdlUtAs+vYzEyk0/ugSkxXp
NVLYhQhAMlIkoimoIf56DAo2C5QK1rynd4edelOWco7DO0h2emoozklNb1lWg4Vp+gQrV5bgOPti
2eMxeMhLLXxHnlKvMFVv2GDsWA2f/dHnf9/sXnP+MztCeaHsBWqL+Zm3v2kIEw0FM5giPMdy/c3i
SbPzujle4GVfyDa0Eis1OsJ7cq8TbvKgmlLOsyTUCM54kYLiDI1xP7T67kz8S4UtLKK/sfe98SzE
AzCdofz3I+5mncpwbV539oGL/S2kXxTWirA799fDKeZDuEU7QzEgPi2cWM3s+wErOfyKWNqbQvGF
QplyIlEvK1ztDJvfnJ1fkvCgLxicx/71JnoyyaXyb8umsn8xb65eeUtAtJh5+7ajjrjv+B2dCmc3
zV6M4NkA7lOexvqA97A/H0mXQCp6gwSZp5czQk/Pw9bewztygT6AVflDXhxWOEJa6xAIHq3MxMdd
QCuPcSoQMKA3fhFBqLw/Vpaa5H5BT04QT8bH+yOvtpZJCDNEyqC92kuGLrgzh5KOjR2OXxiW/+s6
b04tTtF8lXyEspdFUTGQcodl6SUGXlZOozWQjuXudf/jzh2ktF6Qv1KXgooX0avpbrc7KsG8Xq4B
bB5wLiENWD8kdfk0x0FY0tWqgbVQLf6/3kmoTeSnE4C4CazkqVCe0y/E1ai7bRykZBVFDK04XHBc
Wq0skUifusI3K6jXGOQ7GZ0sEslaEp6ICCOYl9m8eLkna70czZ/3bqDQ/mcS592D9DEartC5ifpE
iquyX0pmLZSBqbn9Ty07bdeiqRohUnJgJRWAJbnaZ6CnjQnyOJGTeHPBFLRDvMI52UUYJttHEtl3
zLWQBQkKIyZZJZ9KXQMOnAiWJ2BipAHsn9Z8v5/BocbGl0LzWLICq3eSXYjGhm8wjtzpULOM2p82
4gfJeYsvcv2XsTPk0xBxpyansydJg8oNUKudp6AhCnB0UTNEK07okPK0vISOMHi/jq7Ct1AtjkCZ
9R9mgMnwfoVrtieA45g+uDrJpcKSX75s5kNctrcSTwP6hKVNxQF4PPBPxKWqvtHOhGajmYbNc8Ep
Ti1Qn2oH3VjtWAIoH/1xOyTqG0o4wDP6INMCGZRF4anhGepEEIfrw8zp5zjR2yp312fik3XF7pM9
Q3WxKWn3YXa/p/m4E3tuVtU6KLke5NFRmhCey2hhajKVy4I3Kf7kBhNpqAn/RGOo18tMbO1priqY
/Cl+MoeBqQd4I3mHd4DeuZ3yaR9rebfe8lRTbRHnNEU/wWy6vMgcSH4fTyEB8GG4vw8TMqBJ7MMl
32KVV8H9qIF0apR4AEoB49yEPAVNvUjfj1128S5ACWb6ggEFBL2Oq6I7T3KOC3AWWdmUELue3E0T
PBWBmEMtcnQ56KbUGc7E4V4LohQSDqG7zjMgkvOSF/10J33fKUgAyDXmEZ1xhdGchtxlzxI0mZjT
/mfhe/iXdXiDD9hEaMTyLiJmvVfo6jlTjVVykmVkLA87B1C9dZQdhj/zEWtv8bClu8mC5YAfzyWi
E+niNNwEmYrg/4kNmugh31omeYXpeR7v203YMBoy+GP9kvajHnoVVMxv7rksejg1aFucf74IwB/3
aKYA3gjsZScvMD0n31y3gV9WphmbsTVPV5YG97If8L0IBfJBotdQZdIX27NGT7ZaEL+KSsERls6M
Tj6IQxgZ/S4H5P+LhGq7+qtWsRJqQTwPZouSOuHIOAva4HIlS+p5l3lPhtHc84Gu++jAHH7TC7ew
EBdMYnHjjQgSAbE56rMDRJfF8eP6hEurI1R2DL7Rxx26HmI3iaFqaYOSZI4u5xzoXkBnQg/ivwrx
vRdHFMbPuXVJPMHRJy0vXw7qURyTCdIcmtchNDfBl8a6MGEOdULyQttDa50WOOBrpU+ZpSr339w+
uW16NFNWcLv2nID2a03EDDoFh0FOd0BRcr4yY6T9M1sdxGxxA4qZo8B5SpR4yqyhYnFZyIEY118B
Dk8rYl9X6lIwilEHOyJs8EfriL8iIxe2f4WHaKdBotwnl9AzKFDzaAd589hbtCd0e71mqEqSQa2c
QcJivmAZ51vdDUMu6ShtQMWqiWldfLWZT/t4ghU5Fju/OiRikEC10My3r4Y/gyfUHU4q78VKQYgE
K5nAn+5y5kMUJUIEN9gVINx89FMT+QBXkfzY1Y85uLAVXA8FfI0NmBLppEn7anR74HxdXGvGy3N7
mVzDl6ClmDrsxZUj/1uWtxt+I5AYxqrU+oDKuogcBFYYyMJv0Bruf8HAZcl0f/GNKSSDNn29WqCW
NgT0DmmXzdm8ItKrO/1vnTSjQEOyN6msOcWRG1NbiJhKYIFR8GYCPAtTnBW3vUXYV0OmPJ3XqE6A
c+ZupmB6mCI2J4+XRSBpFH0a18jrbmKVahYs2pLJCfBaYl5ZZnEHDvxV3GTsfwE6R9CqHtCexfpU
SdXYQTOsztiPd8SgopWqKi1RnlKFsN2SeIAEiIPT1Q6SllnebSZED4pxB3cnTqQc8Z/beWisDkWo
b7KdWmrPCKLcC9itLtliEQlqI4fk1atDYP4wseOk3kF62bzjdk2isX3FAsSzN30KekdIYlRmvbdQ
FBHQ9UE77FazOkK8DnBkL7Kys8ZVb/03oOWhxx1kfyhpIm58BicrGHKJb5W+RisGJWwBo38jgaX9
nl9oaJsows8lxfTAh3ug84WZ+jg6fEelXSvMS34G3wQtvVdgdVCC/kdM0+CL0sAy3EiZH9c0t70E
gcm0OtX1cUqeAo2c7VjFZYJkBrYfNCsLD2ELk4nIF0M+/2dKkiEwejsvROmBsjykC5V0HivLmFFA
Uj0ncXoWWBkn4n5vHvoqsu4lJosdFU2fIOgqy2AednyfVSbGUwNKyRypAqYkOkRGk7dfpMBnUeu3
Jligvcxw0NMwEgV6GLZJzgkoRftfKOwKUBLgSMxN0MB3VjGpsRMDSSyPK58ylbDAMWvnIZ/qeKuA
rMWfyLzeTU8f6F8pIKFE3jHMEKD6jlVirpZhhBqAxbRRNJ1QxJK1lowDsMuHQdVp/Y76/Nuh2kVO
PE/f4dKC4WljRBVQPz6OQsz2+Fp2GNSZshSzHIQrBzE0kYbLUPqh71OSouTPISeucbhaq8mvYCa8
c2J0JNq0FNWf600j89jkAvvcW5VtQud5di1IMOL2yYm03sQfyaKqUnZDEv/P/dSmTDO4g6Fitvdi
zSUoBJS0H4HUj/nHTu36e2oQa/jSODfNz+fT4EhajS4/THtFQo06CRCE6MWIxngB+UvSF6mhjYwJ
YFUMmayP0Aj7wg2jnMe6fiThxA8Q0pu+MxJMlmKGWkkMVtcsIXTm7alrWQqtGyez40KsWUAhvBrq
saxLaWou8IWWLpcS60SP0BwbEVZc5JFceqs4+xT6a4svtIF8YBIaIjrORfK2+lGTnQLJnJsXfxAk
N1JLkcJRuGCdf63yGgzDoD0YDI++KVJh/x+fCUPgQkCZ7fpsR995wrHv+aTGKPqCDCXNjZR9gAI6
mXtuh95vMY0wmP6xnMTcX/cTaQgReNrEBhFrNON2RKshh7YoPFC/dKjHsijR7BkJ9rwd3UhXwHHS
k/8MJiZ81Z/0n0Vpmf8r+Dp2nw0GjdALvmAJmlYA/YU8/mNj92UOgxUEBfk0hth/2xu2cOuTl8Nk
/Vxksn0UvXHBJoLprrfteTqptXSLTFx0A6DclgZOVGiLWE0ObUZzA6XOr1GfCLNzBH/OHGemNLCJ
qHeH41OrTn2Ck4k0mYE1o964R1ABg7DfXLUXuQx5QOuKoKd10k0rb2sLmpD3JALoM8YR1ItTwokx
wmF0EiXPj2KQVwah795RmmEQfk76XAT58xUTKJSJV4aXLX5JzIdqKVec17C2+324mwrSW10GYfW5
sL8/eupQcdKSfNlXFh+q0/P3Q3sNAHLw2t0nkgEHcNkGoTJnsXlNUCEhVMYH67nSp7O29/47k62L
lkXzj/KEiBwABi2qxJFSK3p28kDNI5qur/3A5asAklBPsY8b1MQK50CefPHVP0GW3a5N1/IUMssp
PUJ+wxWBi9tyCzJuMGDmpn+3pRQ2RAbfCiPC+0unCOErgAQnFIv9FdzzR3otUIllV6ENU26iSkMF
RhqJ5Sqn1gONUXQlATc8fDUadAJ8Wjz76MmykvhV3grxNalXnLJfTWsb93lWjjjB9YL5SwcNy2Hi
c+pdUJZX/LzW38Ip3URZRO9vwZP+GLNOyZ7MuzEe7hZdZnISxAyeVa1YLT/pwGDSqqRqh0iP8K8T
j6fO1h7e9Wj0i4IArrJzyGU4MOISiZVLrhPpZRchMo04agnPmjGUL7YDOpFyeaXHn3/ZtfjS1Tgz
dIg8/CR2Fjkk/zqM3TsDR5wMrM7AyhrnAk2Kkvcoa+goRcVF0rqwv8GyWcS/dGj3ZUmlTcn/lxfx
CPXg1EWaEI35mIJhcKewYmt7IJuMQSfQgFb+QU5EB1AQOSP6NNwboksZQdDDCoz+cRk9rzZca+yo
CyX+3UtV7qcYfT99pDJjz6aP1prvy0Vq4wxwKxPIUqTXzdkTe1zUSjIDfVS3yTVTDMI+wg6Qxt3W
239d4Pyxb8zQml74LrevoneLpTSJo6pqdzxGRi7OeDh+v4GYrZPQSXXNUn3c6MJ+ys0H4hueIXEe
uBAHxMibNzoJdyB+xOddL3wv/gKy6qOmUSTI9AyWTe7gId0xAUGnuBqY9KawVkh8C5rWke4p6j1l
fLBuKXvIwZkXCwV4KHykq3sMH9YyVtf/jrzSnh+U92SpzpcX4YmY+gGijlSKH/Qxhkm6rI75NCF9
/cx9oGCLp4EnwsgRDXdG1HIpz8KJ5wVVen8AXrRqffqVatbWIYKgong9P3K/m/pqNxageHJ42TD9
tMHuZAcoS8APC+N+4AeYAAKamOSnyatsIAT0swwBebTPwsL9zzJqCrTkkmtYIeKtRgr9nbP2cuDi
Ku3syQKDBZdMZ7Y3eqOZU/MuCifeT0jxKmfPX3eGhUQxhkp7ounYDFLzBsY159DbRvCY13sKYxWq
DutFtaP+5WJI/k9l9RhvYdBVAa1CXGMRq+GZV40hPFbNgOG22tvVZtgSNdfhFq5bgOUaiUEn19BZ
5TfHH4s06sTc/XJToC0Z5uOsGoyQmCW5Uld4w/G9xeyRV0+c2x66iwsvaboEH44XQNbxOOZW8G1I
CiIeg+zU96o/R6DLwv6lrD4kQFcSFqF3zl4/aRf/YB9c4IBbd39VDXbcDy14xSXI/o4s25VZ9MzJ
KYCNSA+wfZYCbFab6Ovv8tD7F/zAJOQNt30kP5xPAth3SSiQmzig0DNgZFc111FizvIvtHR4QPZ6
rBJtdXeLappz0B3TdixhYaZhetUv82IU3fwe16X8o4SgccNh3AsQz6sEDoIKo51vzi/dPY43KeS3
a5ORTMCpoT1uCPOOBpHZRFzll+UpADM/6lLH/JdZLPNt1PPuNHGUWUFniquYf0KtXU7zC3KGo2re
Hds0VfLXN9gOkrWg3lzp4U0QCVzOqadb8aS7J1qR32qdX4TTUfIf6cKCgd9iTCPSn1sC6dkW5wQ3
64+bTDF6H6xpRqm5ehi7fZvJKeT6FfKpNmYlC5iEgfRgNsKCnSzthhNxDFCWpArse1rIVdGpzh6L
VpFrEDSIq55xLx2UrLvQwDakrY6Tj+uGMnI7O5Dl4+yjzoqt90E3xt/gY/RQXttHzCJ6lX4uHd2l
Ho9pk9R75KxLccEMgOvXhQftD2CiW8y8/Fbtey6iBwKgekP7bYyTm/2zodzgF2gYA+N/VqpWesbQ
cBmsX/QcVBrn7QCucnB3oIYzM2FXs0essWpiVUEcGE1jVo25vCEi9E4XRC6ZGm6ttbwXUM40uNp9
G2KmB0g+VNHvcxkCbx8CCi15i722IEEPXoiu7TNfZXP+mO5eQX8d+VlisuSbNdbNSDCyQNxM0qSq
YjvXaYNXSNvv/b37zyPmmkUXt7mks6+vfaE2ItpzXhf/Te5DkNYyZOTmfMi8Xyz5TuaRkosId7W9
ZTJAHQ4e7jbiEE8xKu+mEgnc3BHHXkNj//hEE7s+wcEQ1bcxTsHQM6Iv4INwrbAtBjdX/aW+HMVz
p1JMgzLaCgTGlLyUXLe3RZSPf3VIa3MOvZNdl66cFR9Z9tZFaIIO6mea7HRqZPL9I/81e8Q42NJw
2vwfQxHamrZAkjL9GySIEAluhOLhCU2V+6JLoEMRT4FiW1Ws4b/DhCCAA0oB/xtHMv9NFk1q70Ho
o7EPCUKZDXTsEMyhy9ZAIHQ60/pmKBo+FUYIs5AT8JbsvCbmrZA5iasvqLb/YcksFQD+U+PAq6ya
fdk6y1fkEt40clvOcez1g/3ClGgWgwZVOqlF0ZN1n05j1NqpZ+y59H1ML+SFyz7CpQk0bPSqzM32
vklkmEL5L0MGnJwxDbl4QqkqV1CrdN47C7J74W9ihSAPDv1mEXSOES7A5wkDKCBZlz8/x7nyBX9G
6ZLrGCEbGAL0LfccMPSUZPd3m5mhWFtYdpHJ/Qnu+Ukf7zTutBs3SrXtys7V2UdG779keJZhstqk
sQ86BNRkx+kOZicRWQBZYPpDFYbnrbiTcZp7XkjBu1DmwA+D8/0W8PMMg2HgV5ZfSmjctsblLSGl
Af5VJcQMAIBzbGpSrqJbNKaFkAxPnxjWSXXZ2tq/OGfMVOFom6Wi+oWXHrSyKFw3RZHfo1oNh7xl
ECiZpeeQc+g9c3QCJbeTxwgXFITkj8PFKMa+aw6jXwv4fAXNUUAu6oryL/nuF2ADvdj6AJZfGW0S
u2nj5AJEO25LQMgoQ0pXkTdae42CVVKDx8T4lSFSmtP3RLg6TmRgsBlLnbM2BW/WCzj1g0KJ7msj
EUr6wNITcIvo44Hz9bRZq08uTkFCt5iFo5Qp5ugRPX5UZjx+mjgXlKcvbq6pMq3bG5U+Ybd9cwC8
17Q0hAg1vsdiBKWMQMrfx9y/NfHmaYX5b5Rs3tkkB79aQ/m3HcVGrrl8guHinbzh1Remuf39ITbr
cAXPWIg01KqBoOPA8Jhjcd1rk2F5fQMbPbgJI5tI6vH3jo4UXNdEp13wgB3jsXwnsQborNhYevi/
7dDPlzlicYqyEYOFYOf03eZztLUzm6xZYhU3IdzUaNhdpe2H6wnQX8My1rM9HS2IuL61WkRKDW2u
w3jvSc0BsDB42v3AlvP+DI3T+HJPdsVaZHU4X9pvQEBU2Ooo4LLrA/c90BhT1iwz8qxWbqen2wm3
7/d6vbHKS+JCt6A1QE6NPCuIBXZn7CjZKU/dZay2LKsqKcNY4aRKDvS7JHQq6CqCmDTnfDVy0qWG
oIAvWtj7CzU4K2ZvUSV6o3RjbbHCKluuxsEGsoYpHEYXsZeSBnSudGlmMzqa9cjbQ4H8jh/ScvXc
FoXCuaPSUODQyfWx5PAb20ROcmzLHLe5wbQhT21/XavbEHHzkOYjZc00gPNzHMSinBfBWgnxE9p1
9no2g9kkh/GEIG/1+bjPl8THCgEpxtMpR0dlAfCOAGZheae+AMh/3XqiLJIhZOPFhG2YSWDykawm
iqTA48EvA6w2d8YnMUw8bVkyyY0EZzn2utfifVr87nvUQLVmXU4PO5dKgscuIkUDsJ7lQsf6+Gb5
28gaEdyJlgNUC6K9ucvJ6KWdAsR0NgPn+lAtSJED0Yc83NdngAjEyaS2mt8bcT2Cf7P6YLGfFS4x
tXUtB/FUWSycFMagRNuevmvPKkL9D2U0y/qnLa2ZZCZNf5asZ5PsUVnqBleEaV7z6w1RphML16P8
jjUHABcdu8DbuSHqUDsVFtJa8XdtHzkbuT+PukVrQk+ekH3Pd/0f7w9xS7ldUi9LmnjCxSeWZDoM
AgyoRg8iBH8urLy9Pcr7IYBYtZUKTRgELZZEXbfCuErsZKP2C3byZiCii445WGWFDqbJGVl3Z3df
icoI21qaBUpJWYd0YcujmDTAUKJtzj3FJLCx/k2jJTMLoPYuQA+THog5rstE8h0/eMpK/eZ+9Jpx
kdCDYx6Sc2/p7Sx0w8pSbL9pD1ymbOH0Hu1gAIno7QXcq7qQaZOZ9z/vFxSI1tU66i0/fsrZRwZr
8Ql7REk5R6zxmKIgUGzfBEpf9taLl1NiFLibyw6KBkl22iAmkVH1AQPgnsOs/MRRLGq4/sxcFE2S
hFteDQn5xCqRXv6XMkoWN5fFOKwc/TO9U4eg0AFzSnzS1GM2ND7U9HLDIB87dkG0wwYjaUMfiNvh
FVLJYYfkNqq63h5jDa3wteq9UAeJPklkciauRFD+luesy9t3LDAodMB1lQP5qT+9Vq+H8jvYUVON
MiRzwLQwzvdEIGj+lPuDr/4j6GQatbe1Kwf7/YqnebBFWE3wmDSswDBIV1NLEBgBwfHR8Yr1pBpL
pIWUHclEHTTgpXiZ/3ucY7ZvzSyRb9uZ0ymUt18OM3YzB4E3pm0zOMVEan+kVyNjli4N5iXAGQig
Zxx26yZ34MEhqeHXHAtaEEUCpQfDR80AGQSnlFPtHwo2JAALfpm8EmtMxLDn32qHzyKkv+ICpUWC
iJ3CjANclhOAFKaLi42mZwmL8YzTKvvjH5baLJwdy0cWxZnSrB/LYVln9BFVIRb443iR82aJYDmG
kk8NdUzr5p1eaDQ8gCruwCknHMABg8/nz6heNyMx3SjWuCNX7+UK3l8WcHNbL65VDm1eCAbVfA8n
DyvDTDGIXXwjgIPC/Ya8UcOCSKAobGb8JduJstIqf5d/kCvzy6lz/QEwOzH3xEFYa68w63sbtoFe
jM61TX8wVjxDiAeeupMwbtKr92lLDRmU5H2adWDnhyyQZ0HT4ObMZpBfBBNcAyV3MUtcMyOYTDmG
Vmb21ZkOOQ8Q5m3TihWnIPlYgy+36HwyV7/wB1Y6JaRdoWLoJnGnLzJs/N7dFGE14RZmicjwlBKC
LrsmheMoIvv+w1tHYQCLDI+hV9PhuK+9pfUMqFMkPfVnqf17kXK7OiW6ilChjSjGNcEh4ZbDq77+
nbgVoBPsdaO+jOk4ydOagv8jb5R4XgyFbFqQjhfRS9FiAXvoU8yDw+7l012sGkD+sdqapmonuIwm
RuKtrgggjNjJc+zIFQnU1iHbcmGQXjG0xi+jR7a+6b7JDftZA1NlORDmXfy5g99EMfrc+WbMTUTX
hZVA2wYdgomenkzdJeKn2ijOsZbw48CWUU59gJkAdQ5BACx2VXdE72NIz2IBnygN0PHXXoSALKMr
FEc64NGG8Zgq0zii0xU3C8WF6JB/Cah19F2Hr7dsJw98Oznw2XDMM7MO75WUiEHoZ1k6v7M9ym5P
GF9yALiwbN6Y/qHtoqaBxzLA88mQI5O4lPVLsCmdYes5kcy02EGK22nDu7CEOOr8U9LQYQa/PAsc
PFmvjFKcRl8aQr0jbA40A3ty7pXdYqwxPUXaHUERPRgfxXQb0d7uxjIY8GpApfB64t8tyRjYbZeq
cDHpIkaACW36WcywGt9a1k9B9S/eNYwbLW75ObvElZQO2wO3gGKmh97zEX3IK5ZifB+Rs30rWRAh
WgBlT7Vh+ffCliOrABJ5Y5BuGwgewZ8T+vPdKoyd+RHFAInU/zrk+S/e0+SbDJB58tawC7gcVkON
gTj91B1kuVumjHVomB08t4WoJfl1ppvLfTWTmzNVlYn2WFh9GgPcvIJ62nokBYn5wnxhS+W4Mfr2
KL0JeeXrHyny4RQwkhy8IE2dmhZPaUgBunwY7qNOvSHgDHya7jPHGfADMqKx4O8UBOvKme0edop9
IhAO1PduW/vwtWseGFC4scXUe2EXdy+y/18l/CCldo2X9ahqZj7renTF9NujNZP4s1nydrpIKbaY
0fNf6eFA+gRFNd+pj+Aro8GO6Idn75sSd77VPg3hueVu2CupbGaKW8orWNuHGwcbncKi56AdcWHN
TleYHq+pyfydPHG45Q71xGprOL6VdaNYq2GII0E0gEBEZrZQbw6ZcaTVOuOn3h+QrR1cHoFNcz3p
+xGADNojDFZCtRrndHoTHh85LrI5vsIXSdVmgh1ufa/6/ACncnPO4kHqh+St1wL7H43CND18UFzW
liGNbv0Gtgvl6i1IU8mpQywOBuGZj0HRILEwzQ9pygfG+DthnfYKR8rguczHSRFliIx+2DgDAUqC
39QeN8Mrme7e0l4xP+U9PwsrSivxANYF1ADTG5s1YAo4hezaqIODtFcSGGV3rVRFg1ucnemG0A3M
onw+shCxXflmKJfonrRptssvM0uRFqakfgc6Zdz2TwKEN5ane5qKuR73xaP1QGTBZU/Xo8s4KTvW
LZBvfZrxrA/GkkNAIipcGAFseni8qouomT0775+OZc0BGW1FTxL82iyH2CX4m39eYbWkbd33mScn
IVX5dcRJSGteXAI7dxaSNGxkpvXS5vef3Mu8az0b8P3zUZaIrZPGKB/haz5drV0JB6sn5QwwcfkU
lGh3JDpLzUC5OI8I4rbFvUZVd4F74CbKNjo2h/GXawFUt5jX3XhFSvO/GxKr5Je/PZWP258B8zKI
d+ujiyjV59Ca3Wfd8YTcdf7XagybI4Pn/C1Tvd7aORZnhbQ4eyl9SK9ru0+Ddn59mJfe9plEggRd
UDOONIDpvafYrAv8fDB2eM1qMdwPxJmEPWNCuWXx8vJWM3XhEEb4opAYcRy0Ksb4hxIfxm89+s8Q
KrCuvC9mMDV+IlN4XKKFePrwSMY2dIv52HN/kHpsar70mixx0AJjEO9T/Cwo3wF/GkszCW4tSrAM
nVVs57VfLeaMh5RTzgMQLa0JRlxe3b/ieUcXKn1VUOSqX6ejKbjnsoJDjhaJajjpLZGiq2smnoyw
vpbC0+S2PIyTZDYLaDgTEnOf4VJhGcXGj49dvERQ2eKlKH549D63tglg5RoyWSLEHN3rNVfdAygS
vedGEZLgTAjylpcprKEZov3LBhp9M4FciSe86qXCiPVWeOC9vXcgsOhPohcckqEHVrdp/I+fLY0F
Yx3shh8aag3SZCxiK7QBLeZO6paz9gov/TVDrSfH+iDSDi6myF0549kk8aeeWh1HBsJUapjrAzEb
cVLyeZ8dZ9Pj0If+ny+4J/Bs6ZnRx3xggZ9V6g0+wU9nb/dwTj78EGLr409dCWwCeCLY9tZzrW/w
HbK+pIsTdpTXUCt72L226pqoS0j0qITQITeaA6wL09LoXzCwaFNvA7octseHlXBWyTgqsOKRuMUj
QO/C/DiU5FVXvnzpgw7aTeN06DM/HdzX7oIKaKGqB47k48SHrezCTFmQlkxZMeihT4DPqZjcjHLU
OGWkyA7XqbIy9ToheIlqRWvnpfwdXl7ble0kAqdCMXXn9WJARLNWz9ySuo9Hx5HyafsheJU6Ugqf
vH1BnYlOKhpL6/smjiciMIZoJvkJCk3axhm1Y/b3Plzob+3FJUETRS8Os9kcWGsWn/Yw3A+j2+kZ
r3lDLg3AxzaaQh+oe52IuBf0KJ6S6QYFdrDUTi1nxjXIfHvycXFWnE84feK14ZqFsLl4tv8QQQyD
kAKnh5Xbd4zpjNq6gwM79sGWpC20AzWcg7d26NCg+uNPznIVvpfyyzHVJlL414eFINJ3xk0U/bvT
fAGefg3J1XFdwZwQYNP6AOWPaEXe4ufOm1jZgeCjZE2VS55qhLVmOw1944PI4isDwlbvZnyP0bVX
hi8dDBhfQrZPb77pAzfDEkCWdUwjzRO9CyJxAbTNY3WFrWwAXkpDl2KXhXwx56h/59wL4irlXBXt
a33FoO+HN60to5jNaVNPjsuvPxeZSAoQn/qZ+GHaSYwf7b6F626kK3gymraQxjTESAG7UmHGYFgn
XM8YO2d11yobpTmHxQlp3d0059dv9ooNCevtfCxc8+7UhTU8CjvhY8GjyZRYoz/f/H9ly0OF/qWq
lc7HqddfJSwSe2DnTR4lnNaX6FWguwTA4WRPzUWWuQcBnexPJfy7HEEbBxFh7O1TeRsjlLFnyZ/o
yN+mvw2sGPiyr99CmR+aXH/KrromoO3y8GBbOrk6vMhK6R+CDDkPW27LUrqJLBqKwSS++JkjEVkE
r5kA3COxEfjuOtTYw/OLiq1BVWiPQmsTtJLxiMgIS4UNJljvUvgTNFXZn5H79c80G+Gq0grcH/ib
BAXUWVud836cc1Zir58rrakq0/z4KICWz4fCqyhpa9i0PLPhMP33SsrTvEruQK+NRr/R+mOQ7P1y
3P7NaNnFlZPoeyjyYZAqWDw61vJVHeiaBQ3VWXEeVtYqz1eDxTdSR6XTNz/j1MjDBj6XdBVTemMm
4+oPa4eLDwUtonGR0mDnaDnmNyiOux73wQpk5X7xD90CvksDJ6DEphGwHHA0L3kIz+5bR8sCczez
6YGEB1mC6bsaIxFaUfZwVQn2Sjat3yl/kjP2qwY02OUBR6evm8s7haFdJjDfDMiXhe67MfFq4LiJ
KwEdM3kYIVE1VLEft8LpA4xDeN30lz0XOOWtNbg+M5uvGeKukz/9cuog9zEnlIE6kKOry0XEl5JP
+N5wI2ehFdF/XM8rtMbbZmqGftsnz9DmbrNl63fPcsLsycnUhb61NvsL5NiKG6nwqZ9Af4WMLpi6
0kv8h0hNjP/awpsWz7vBV7gfwRnrO/fFhyXBVWXXvxtzg2p6YUCxdWKHU5qpsSI6+1iiMxSHO+6K
OWvfdM2b5oKZZSWrOJ2F/Qa7PuuMwVD4rS2o9m9YUL/Da7wDAjIgNpdbSnygQP1hg2PKbwWObxZt
hAPHLwWmoSJv6V/QUMfbcp0ePsRLAK1pll7HKgnLjEXxyE2RZPTQxIKgGhEKIEyIS//uJ8feZuEc
a7/ltP+Wl7RfVpI/szVUbHswjk1xk6Dfl2N+CciOL4NKa+Z709u4J/ZKOQzhX/HevC8tdWCSlaQV
aoXIragSMy/gGXB8LBo/AZM6ByWMzrZldFqB2mN7pASPrA+pEBYGJpPLKmNCtOvKlPnX/AUXpiUU
65XoGHoUIg/L8AhKiNUhdGH5Dt63CKK0duTz/ZG+HcIQWiPyoeyanlQFIQ35AbVEX239s7XpqGee
zPXQkfGwIDqJAjJzbhzPbtf1XaJzsWlyOzbcH7on9S3R9zE0fzkWMKvHNi8IhfaRBgQPmEc4LPfS
Dfo8Z9UW5h0wQ622rlHYQh5R+o68DK8zRFsvPKKgfaA4Z0UGEI4fB18+mwEJ1mSiI4u0DSM6lVmo
RfF76xbzlsJ5Lih1sHfXs2Q3GmhNCB7NY9AKyNjFjUvW8TjLZKox9SZC4a7FIX8alW3aiXyIRN/U
0qH9uFo7gi8u61nWoeHZTFsZl0dCM38ndmstgpaY681SOiYhEmtZuhujcUE8oBJqILDL7Br3eqQy
6kc+X5VTvSFCkrObc2QlN7nhOK6T+kB18TXGzAnxyZtlYO7JrUOQImdCr5gkG7VSRDoUkeUuygQM
dIvQqzT53GJktK+qQ7JpfE8lrFptyz49vAB3MoDmOS620lckMPJXz59yvsW1Aq8wBg0xuVtwYSYG
LmZhIHn6cTesyeuHCcASpcTid2QPw6h2aSYo12Dph+8xCKkn4fF68J3L1IATX9R7jxSM7jEQ1vzG
yHDT0yU6sIGW8uD99a5QlwLRIQnCLZV3O3WFIf1i0H7FYlVZXuFuBPqpcobow0M7SmvJyQHziGLq
wsTTCJcvaVOIf6FRze1yvX4/72Va1cruLhWwg8ihK4Nb0fbrj4kQnP7R+M1j4iF48M4qklygLwCc
/xELx4borxf41EZKLqnzPOz5UFcsoPK8kvk5zdIwGbX6AWhLmgb3JUOmpL+BeHMhThswZI6eUm9n
btTiCM1N06Rj7vOARZQJG0+hdVvLE2RcyCcu8yfk9UHhH+q/d2gSCVaa+dXcv3mHKd9ZI6hYJWDa
uYwf+HwTD1HsVwA5JNIqT1SiOeLs2oMJOOGtUkjINSYQFwj3Ane5K7uwrN3l0QIEPAU2DFVbUq6U
SMJ4w6D/FcuG+NNIZBAPZteSdEUddCz6h/0VaTc1G//9nTNwVOQzPUEV60a8usruB4YJD6p70qn1
4IFxDDXnakhr3GrSzVW+8Dsbdv3hPfvs8t89jphu6Vxhu6fp83BbdFXVp5+RTMXuxSVldOyrYaEm
lPDSo7v58iks1mHGVUZjJp7yHq/GeId9Jy3128bmb0WZbXKaR0n3iDz5NIJ796sJXsIG8u0q1xPy
iV+ZeN61+HK5M84Mf+IY82DmgVWa88CqqPcboRNRJO8/IZVNXvLlSZdzlQmxDi3Bki8cyA7q50lD
J1ciAaSQ8SVBtM5fLQ+5fjYzP2ieIVbU4FXnTHIPirq3/1ggMWT9/FeStnbOVwrzhHyzvEh91hq0
9DWZlq1DX2EeqqBxW21IiLDt/a0XM/tlMGs8msVEG/jKzmvVyX5dRxDgvS8vRPs4ArbQ1pAU6zuz
f5qm0v+3O52vuD+rUGqXAR4koKaX3+WQXnrPdzCkB62tdzBV2ZaMREvnABUa5W94QWeLtJbMl8Tj
lmPi/Bp96PEWUztl8HZKmsiRXKmXa3kNVIH+dbm+5ttSfzUCtbHbDoFiBOEm0aSpKHbv+N16KR0y
KipClaLPMcdk0c1hqMidYpBrC0KEc5IXfOgpLR8yQVK34QpQEJOsHdSQJG9fW5pRbIk8ZKVXhLHE
yhj/NKhHzso2madkBqrMxikYquJfNp+GxQZbmQQ5weRwfxcsUiT9oNB+GiXUOaQ/drtQEH5vFiL8
WEcLurq57yiVopzVFWJeuqqiT/uxz3W9TNtV0LKlqTRmW3O41S3/BVbVGnBT+h1GYBkltSbxosxW
Idj5LrlUusqMqBIivfovATKT4FzarEpoQfuZnAI5/jAbo40Gr18Jv+NqMEof/jv05Z1+Qo1KygUv
fodsnCzyRp0QSY9HQ6e7BmbxSo8BNhO6zcpvakz9VxSm8UDVj5wegLkZwkTLaExc2WY30nSXh5sv
kpzXY2nrs9kskj4T8dohQnAlEpURnK3nld1OeUzZGbueQflQlPQ2aIt5/DoXRxg0CbF2DgAmCrqE
y2q3Fdb8lFCA6b6WdxJBO/ZQ2EKzn6oMWtZAIRy38qU1IXfM931LidDsxvcaGpcSr0eCUo5uSvhl
mEsUrh4beB/h35LKSKwCSRFRKYGSRTl1LP0Y9a4DicLGsrms+4GgDzZtOviVs9vNZa+sX2OeaJvp
Nx2jCR7C+QLJpDAXCcsSxtoeZ+pZ0g0BaDNBVAZMM+xosemSMievIduX3fWtPKPu6mxaPxJQWy0T
/0OJJP6VBgiNDgZB6drNd2G/Cyh5H8fBEa4f36fnG0tN9bLJbqFbq2B/+mGWkYnZtNIV9GRNtkNH
Lrmq/+PDxYvEK6N7BqusgT1mH5ulxTGDaissMCiuvR+R0OzDK/rW+vaJWIuw4dP8SOdqnaWd9o7Y
dDPxlGAfnqCZFNcKr7sN+BIg2dqvYPpEQKsGCaRlqEXTTQZokWfnFzv8Coc06p9lb4cMJvnKt1VV
FDViD1Pb68kYIUNFMjSFXNaSVHUup1Jp+eE+vSE88Jvqn2GXE+IZbDJTB+NtYenXR6IVfXpr5/hG
y9enrnV1rLmrOsu2YFmwH3Am6HBS+8ktWt+hWvMvIHfBLgYIo2KV3sP25NvKqlg4nnDIh+9BqeIw
JyVLeAY88UbZ4vqnIKlGNQmpybEoWTXEiHMbxaTg5+9TLAEQ7JUmoDQq0IFXC2UlkaxoIw6Busn4
rLrZma5MNdj/bOI7xSm/+PfCXqNZj0fhNfCRSiE/Dwb1RnU3Blu4sWDtfMbh6mSCuO+TpLRg1lq6
37uDxiUUooClsRhHb6hX9vYuE5AydnOadb9pKMcF82PpNBcB0wmS3S5o+gwv885LeHNR5IHgii55
IXooP9VVP7pC02DVz5dH4sI1/nigm906vuWFdnurWX/n8g5W47QBN/VlhHpA3eq1iEylrszRqp1D
PAJ88Vqr2GGwq4fIIxnTnC95D7Akm6pGlYR03pOVZNX72kBtBTFyiID96T9ygIzUBU+5EtYKfgSp
nxOWz3kroBPsz27PLXoQ0DQbWsh7vpIaICE1NerKUesauVSj88CxQ2/y0RdJ4t6Uwiv5FWynWX0K
sHzEgCsz2VidOPbR836YldXsgoXFX90SF98NT6SPj8Jvf4kokY3DP2Joc4D+PLCQDFGVW6a1tfKl
VzEhF/xGlwtLIUf/36bpfQ2EH2XpHPElkQGQ58hZ3lA25d8V/G7T1SD16QQv4fhe6XDHktKOh0TS
SrgT6cSAVWNH0EHS9lNkgI7XdOMCIA7XFDbtjwUgB+e95vMQFw993LcJnLBag6Umvihh1/u84pwZ
mnT9ON/R8H7CzrHrqGqS/3y6TkgfxxICUj99xueE9l5MzLFJBMQy9cUMWig7TLmmDdwTCyUHHDgx
3eR/MiNkfaDMnSempel3Ev77lXu3AxUhFTD57y/1xnPUS71lbGUc9L1JudkyJytoAK0q1J9KKbsC
wpghlKGmHoCVrVRLZKTn2dj4/eXls4ky4lDOIbmxKWH/h9lLe3aF7kxFfWKZt4eHnaDQTz+Hf/EE
/rHjotmnTB8o3NlB61mYhREbEfDN35a9ENcg/gtei7dJ4Q/UesGtht/5RAHwnzXigAvQWmA+k4Vn
JjpwwNPzBfLxTVJgBcqpjHm46YHD2gUJX/5T5nIznfpUU7QDhC3NVHikenho6Z0w4aAZLjsd+xjq
MxWVOx1q0Sscuw8Yxwki+7yGsk6/VtXyUy4IXXFV6hD3qhvrZ/R+dhGE8MTw3Rvr+YavcazREs/C
2qDr5cWT8v1+sWsTYcMYic0O03/qPBjgQmCA+IiVwgP77KYiHEfW5A//ZD9YVfTP/oz/VG0620Hv
oNyyAFtu2P8e+7ZUBc97Xa5st0b3/OtNQvo7SZzt0cF5vw8zPCRfkUSdBuCzKXgbCteYs+xlNa2q
ceNsiNEZkoSi/nYp2LNkBIalke+C7L0aNq6//NxPjRdXICINoipktsRHZhqMlomqus+h/D03y70n
ytF3cYMuOPsbu0ZAqef99zD1DOIrBupZK3dMbM0jS8SewEp5VBzdeKgbO1WMlv6y8X2aYNvDAqXM
ExQuG7ldl4cO+bhoV97Gh/ODcgLIHxqd+jVi8PBe7NsuJZL/yJSa0geHyIu0tpDd6es1qGDpR84q
gsALEbpjKD+176C2EofheP0VmqzSLM5mY5pK+gLRrMeqv3QyPnh2FeeU2ZAj1YNO5Wihv7Trzmcz
khufwGDTlBmZK74Pa3293VD7GYPcPM/KLQ5epjIBTpsTPq/+zpmBCnTTXdV+z0jORVmtIsmOcGEQ
3SnEjW4ZDumzNvuipTUyBd7j91p1OYpB23Rn2aP8g83gvWgAO2SgnsPwrfoZ2c7U8YqOKAsznp/I
Pxc5tWENMeAbTqgrLnbsdBLDiBQ/dBP48X+dSMpCdOHUrCti5ogHUwiFDzGJ9vmJCJcdnnC3hJXU
tI86uvsjxAfpciIKhb3i8NqxJRnuqQNe8G6QsRlkrBTOofouwzL5QE0zxXctusiMVvwAbpBLUgCh
npUk8VcBJiKrH0hEl+RncPxjqTbAvhPk9mG/BCuMRb6s7EYgojUksfgs+Zf7TML5e3hPMDTJXUlq
btU57aN81WuaqeVl1O1uECdFcFPgg/1LuOxi9f3fdwNy+OiBg8kd8+zNm0IDbvf7MT9C3RK1TxWO
A7VusQnfRP1DcaW0rKD4uHfSmyQ/LuqASiJrKgp1UqioLemxZP84aPmkbVlLaUYkOXTmyVoUmihw
bJvpK8KlvTT0Ut3SNDfL8q9FRuExqtt/Lws8lyZ7qb3dcYo8u3RU8vEYRy5PScUrT1mqqBFpuR+7
+cZOB9dbancbyMmMbHCeIpHEYFfk/INODL6RvvPzEQqk768fA8o29NKmYKx7GAzxQyPdqFNDkPaY
YYWULezaEvY/EWZylDVNCKTZTVcVhCTJWRAKE3V++qY3lze/pghSBg0vdU2OiVhiM4CJCvDEsSv9
Ur7Q7HvEtrGLdLDwPTBjw61MmdS5qwCA6hlZBrKoMo5QEbXkeIbcYkUWo5boiSwipUyHjTdlaZ/Q
hCPwwtBNZKvJ/DaxmR9Jn1GMsP/YEGm/Igaa6VWVUpzFQs/gh4V4kIeNPpBJxBk2zm5fLNJWjvNR
yuMuOrzfJk05kRR/kehOGQfAIibxEInnC13IoU5Cg91d1aekrZOR+t0PdxcQIFQioUG12KbhaCDv
Ixoaf3YqZPOBVZK2Qqkcd4SHVyukmeU2M6Rd2eKBBC3M7KAol2+b91mgQQFKe6sVg2n8PHYzSEwV
JeGUzaQOQuN1x7rLVzkr1INrSvxJNRvIJ34QKiM2KvJJG+NuJrIxRO24cshYbmdcbo4W1KYUZ5/R
ink34Ax+01grnMA5qX1TnFv++1h64sArYeBzpPDCcNQ4DXSezKUK0NQILnVPlOTYZOhCUb88hWTE
gKxEJpzYRRnp2Jpziks2bh4mOxyUGCDVUmPqJfDsUmiEpxJxa/zUsuseD2/RQbC3CtxIj53hBcyS
TFjamUn49w8Wxa+TJi0kGHRjqRGxtpB+GGc0ONIKOMeNTUsILfDj2qVTPBqIibV2+hWcQqf/d8fo
BWyOfu023clWpB3RYsRdr/29xZPp1txv7prVC8zXD2H0S0Md49CEg4+hyTr/mThIWnyx2HY66inr
RvbQ1tcgPe0apyPzNcy+S84FrL14hG9irfln9/pYJPLaOmsUoE29NxBG940ds5EbXVy+TA8zQM5B
21z9DAt6EAyIkZdSYDCJV0JazZjv15hak+ZpQ8IhhJ+2ME0XXBYSislDhYvfoIu8rNObiZ7pyV4n
Gif0ky+iCsentVHjwcItP8C6v+HNV67Sa/wlt7UJzw1t3EuQ9jhwqGjT0hlO4uQW/bzwINZJ9I/R
2Z6dIsUcbexmvHG/rsj5K+gNJx5DVcULgPG9j3P97X+ksRITocNEpaspeAigk3UZ0O34AjUMNY7I
jdl3wo+e1G+iMO181P2Eccpf0f0AZxcCJeDKEOt0YIKp0NLd9OeES9NNSf2F3cYSC2Adtu43flSU
LEmFnJLf1drJQD+smL7mf8TZzJy9FqMHHZz/z6U/HJC0YkR7cLdSiUZVzZvVa9RqrgBY/cF/3hpj
mXJtY03FCotqefdrGn5/xTZAbxo9dbP3m8l1zCjsr19F4PyYDJncbYv3YI4BlLIkLR/wQBVeFnKd
nzGReAai7dr/8TggqHDv7Wr0GHjvesatA3jS0eyFO6kUxqQMX9cMa/mNJ5fHb+njz8jcQ+uRVSRp
ptXwJy3yrf3k0Li5bbVq6+70ucd2+bMHhjDWtQIyNFqqhy7SNFgGR8oxO4FwTlA0Y+a5e24dxl7x
4j72+gpzNxwwHNy2duE+uvKENpe4yU8PUqYxxqZ8nlE8Wp/5y/yB5N+MLpT7oooi/nn+UobvOseI
Q8Ily7AwJVEOmU0OgCZwvM8I3k6H+Zy7Mh6OgP5HgNolZhvEhRn//FWQ36SY2sg+L5o34ve/8sJP
pe1QFYo6UQ4ijDOfpZS4F+2UxEwFxq2e4vdjvlZLOY8ZzPyLcPtGLJTXWS8Tm35J52ADzspTmpuP
n/UFB+U7olGA9sCxr9w8ea+pZejkLZYwBXJsAS4inMukUCMFdh96/mq+NrW4VdIBN887AEyQ1sVb
82AsxgNAedscoee+mu20lh3xISRcBys31l5chX8+OOCfhMD6k5IHJPjy9UYhrWNfDu/khN9eNqxi
oC5aKX8Pna6rK4RaRMg2YM5pFhN23ydJZdgf1cpiJukXyZm98nXEH4iSBnPXZIX3JHQZd3sCAbze
YsX5bVcOJEijtARNs0oRBQduASu1/ZJJVJQDGkueF4AXT9GC7XIdsALS99npKq4+SAsQLetpeCG9
5+l3uSW4fl3EqmD71nOLqouQcZfN4/jebt5h+eoDHO5iKE2+BiyxjzxRTQvObOsuCb7NZVByDkan
YmiuV42YDEm43NAg5V4Za+lzAP55isBioDa8JawEMCbDZBxirVJy35pFmpYbu07t64fLjdqSYpnz
3M5GhibOX3s7UzXE7cSLURjcWBGziTspQwBE1D9ZWDj1lsnN9qWtkXA403Ck8oXa7zgMNoM6T5xS
xhwFYjve89gnfwg3/1/FiCtDRxmrRoETXijJFwLsFzBeOSDjlcWt5srnD5sOPzih1pCl+W90GG1h
59E7Bm1jC1MOGrWqXVZ3vE9GQQUhv9rQjHdpUBd9ki/aXvbvsk16voR2oa01W0BEbApLh/mlx0PF
IdjeDINRVdtC7AkAwNCVZOax3xzXimItSmIwJ4ZGsuQ/65T9+AKkYqDIlaHSkPptdWcFm5E7HBYo
ShNo4t+1Yej9X53fu6tjl0lELpOhJXQl/+Q4DViHZIKEiHxL978HLbVQrWKt4QVwzb8cRtEVjif+
LA5z7opfXPJ5eOEoc/J9tynk0ki0jM00Ba3mBOxFSsX/ZONqommBakbwR6hpkxfVDAyj2LzCAvsU
hoMIRoeBg8xk8EAzl7Iqp32Wm1ydjciETjG8MDo5MSVQEmtmJlfqeAhv/+FhQJLYLH23eu52QaUI
MZcrkefgjZcRg2Hfu59PbziCO7okxJCb2IJPy5vJZ/jXjfsMCd6Lxh3rvR7ePOYKHaWaYRZHhLNO
67vGXahhPgWPL/Uklgm07KGZS14LMkyJsBsQ7UX0YCufo3KknGM5wqr494QThzMuba4aKzsfoq0B
WjT2kfOKJf/XjT1mVHELjALO24HUjHAFtwRDQagfXzL/B7zLRIjEEecOzUt5EC9HPp2FW6iWhLFw
NUWpulXBMVJx4sgwNTL6EgC1yJGEMTa/WRwD+0kwmJWXuSriG1K+9kxAk3ejXOHd9MIk05REC/kC
mcEZxQ3UoGCra+HAnMGA6sfrCz6+3vhMnM7y2M2HhGH3kFJYwMaPLZTHhjdp5BjW0saVeFGwNkEN
MYZ3zIioQ1+uL2iJ62lYWh657HGRdwLBdf5SMS1xWZkGb7Vf3jla8cI9BOoMYkd1RwCDKo7dmG14
ztM+PCc3Pkk9SWmCv4c45Kl8SQXZCCeQ/+q7Cr4yL3vp76j8hQjhPHAGQW8tthFdnn9HZRI0G+v1
vmVZuks/772TsL6Vnku2NqUhk8fViScG4BD/ZZ5B2noREr4kzUn882Jw4qFIq+iymgBZ555PRCFj
GQtayZWif1lICZy4doKOSoctW6ihN6XPJ6ViEfdouDWlLH98J/afVy3U3m2+ghYaJRQ78bPCyFLh
fKiXrteNVEZYLgkfRQhNx/UEqcZ8upMSgK3y7lEp8vv4AKX7NwFJAtu7sJwiRs8x+D6/V5vZLBE3
687Q4Pp289xbRNflmj2ksGgCFPBeHIhEh9YvnFYPFscLJBmbG/CZ//arhqH9adVLNJTufqqv/oeq
axZ2PeFI0FApGnjIEdZ9wS/zjX3etlEf08yiJEdfZyDHKFgw7CUm47EA2CBhWvjHObGUmG2yNFPP
E3kz8SrLBw==
`protect end_protected
