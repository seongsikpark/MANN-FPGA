`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
dqfk9kqpHBtf6cHIzsspVJL7d4TJjeakayccql73lUuXXvWkQzlBQSFcyDaCslhAd394kVPvDfyZ
ylEwEPfUXA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
MjGKCxpS1CYuCcusXYMk7wgB5rcnHUJutA3ek5KzAXVJH6cX/ghNIr4Climvb8r7cln92LwINJ+T
+mKqJhOZ1lElekIi4y+R7DkN5r4gdyRBed8iaiCInvOf94LcQqdFTDoXLNJfsIOKn2P5Lwiei+lR
mYc0A+SB3WNqou1ki1E=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
GBm6o6T2sHP6AV/xYZPFXi1/VGlumot/faM0JUk9MvhbxVXTQqAbWbjqR351pjF1iYM2p1OGZbGI
l3PTOul6MhbkYDvdhpHXTz9KmG6JQmUCSiU2cCUKeeSgrvYPool4AWf8S50NfIcBZV3KicX2y+Km
6ZSgYW7HlXW4ZybOAcNPBEED+rIhzkLscmAgAOHLId6SLMu0M8X25tBxmOsAJmBJ+gk5upnVjwkI
oz2fsUV5MYngidBeJTD5BjHsGsir0tIsR74F4IsckhQg91fPdc1cpXiZTg6GuedJnt7Phmew15Dk
gWYLibPon8Fjyp5j8Tb0ndWC547WnNrcNEnFPQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Fcg3u8noyY94nbzwk7prn3WN6wuKEaxOnrxhhTpbWBZmMiQOl5TVAEDyW7/alyPh6d7QRFBeEGEM
zGtZwpTn/rHNuwo24NgImek9Qe7IlOndgOS0YabaIKFPrlkuUgO8/C77F041Z9RjRkb2Y5L8RhjJ
kAedm4X20sUOob04508=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
lRweFwJ37l/9bvPx7ZS+K6clRN+gmuGe2+Fu/tct0tKpKer8b0wh/J4tnv2kuB5nhdg0F5+9i2tl
5pCym4K7KOqaedHU1oRBMuXi+aQxPT5Xa3Y8eXUlXSVAttLhJv/FK4WwOrxeNzMz1oGrY8P2kLJC
6VkK9crtlnrdUYn1xtbCIvIUQGXmfhEEdwzMImsgeyiROtBpk4IOG3WGjSq599NEZ1T5mkEi8RBc
8kUR2U/kAgol+JVyeDQlk0QgLTqwnlRn4THeA38iztmUHKn4xxj9C2y93MzjyL1XC5ItXahq9pLF
YziwZ1nh3iyKr7qFAWZ3E1RFjf+3weHh88TZeg==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ooA4MsaOdUItQVTW8YDp6hI7u//4vhTsbvp+9knA4TwIe8BtkIdGFqnuhiuxw73bKvSzSXVlaKq7
kVI10wAvqsIR3UoPduTLoS1d8ht4BtIyzaLodQwose/0c8Wh/TCR/n0HrFk0S57FM4I9n0NHc5Gn
qOxEXY94q7aQXEFsymeaDe0sajjsx0gtbRzmSr1nJWCo4sLo/5Wou8I/Y/FfiAVbeZWJpjj6kocE
OiB4MttBLP70NQu1kcXCuW01gtaEPI/1EaDJJ6w9ab5h0x1qNwrsWn8uTDfdGGswZf/jQ38Y6PjI
CA0nHPAYrumt9mQLhIRJlD4k+jQfAas9YR9Zfw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 214080)
`protect data_block
cNu5ZAIlMM/gaAbICZtsv3nn2D6F5zVExhg/BETWW6fTZU5CL84TNooyHsfoGSBJnZdqVrkGiVPn
rxzj77nDtgCyQIpo6yuJ2e4RK3HhLiImj6hnATK2VDI9IieIGnalXP0EqV4dtzbHy2Y6ylgOIc76
1ljAHss/eoifUz2f708PxN+LEsrFGsOwoqovk3wxDh526WzigaNRytXEsbBZavwXQZ9E9OGqWF1D
fgoZreXYBQfmsnBiKPRot52b6AA+a6RvFnkESVplEIEdkGddJELfzDW/j80fhf/w7fbEECMGCtc8
mbPYEdAJXaOMQFkDY3Ij8FDJ7/5knIZ/vqv5UMfqbdj1nr7r6fde1AVAg9nBuUyVwFIDK1Rj1iCS
nKKtO4E2PDhaHESNrdq1wMZev1+eTpuCQoFpNiqe8HoYgMl7CskKBmrRSI95SGhR26aLtQvpKRUz
iJhBNJeDPc30l7FY0Rs9P8Pqkrg3it+9M0w9MkV9JlxfrDJQw3NdFuWhJs++b4TH7T844lNzuMz2
4WE8OcbJ6i6v6tOpomp19c94P+LCKPUI3hwglnIf75gjNDrgtdo+Qit01c0qw1yNPXNZRg7UH8G7
kRiRxMqUn+m0dRIAzRHuhkM8graW95meNNn4OmFcwfJ3tsV35g9t+AOXisE9TNkV5O1bL0bhb8sS
IDBSXj5mfwmxOQRKQgtISe//vcg/PPZYF9yeUj1CONMesnmlSVPCBGclauQtwK1BOb6Emw361zuI
qkXcauw1M/c0mfTVz1FVryFhSvNqnvi5ssdAw5OpvCPugY9YuguJnqzUVA68j9CJS6FhsQbHoY49
YUOHYFewulQ3Z4U17hQ10lO9dRQhCatwSkmxsnoTxms7DY0qYosG2+iMESBZt08sNtlbJAacpids
pwHpjJ+5f8B4h74zt9u6lhc0Yn/PERJ57EvmTKBOwhVxgpgtXu23oPfOOBjC9g79ZgE5/e/E0eN2
CBxtrqooYgYDjFerLQIednuu3uCHgyOsc4FLggW8KeVTbc0df4Xkh2ga8NPM2r3T95Iy1bLU8BVe
VoXZtIpFYQcfatz+53+6pDB7zuPvldptqnU+Q0T6DYU2Gp9ETfggRSTzUTUumA7O0kLKhqMLa4S/
kdI7ImDzcynY3KTNP02/fuiitm/qi1cflJuZe2/V6Aw3m1O6cY5s+UJz2H8kU6R3Y/q4MTubp434
JLKivCIeLdNAkyr0VeZmiq4ifg2qhRNTT4YhDm10IovcDss3qRWWItn3F7tVQUqkXXsFlRSIMck4
JJTA637T1CAfZPZ2BCpG/XPaAMhIS7ObtJT0egJ23QyPgik2FH/6JYDkNQ/KKlIk+0QVbKZankoA
Zia2HRCCDzcDjiTuXyOJncQqUW3bfPUpdBXtSrt5bRYikxN7D7UQMSezXe6csAfhZa9oIIHAwa0E
31qgwkRIB4fKXd3uXSrO0XoGe74UHzlAi0h/BBHuihaPSU1IFvpF9+aXBeBZm4CZRiSn9CsL/66i
+RnwJFgau2nuWh6GMNZPPo3SRj+Bq5+SkY1ZRq9fZWmqi9ji+mc6RWfCVJN4WLhHUOoi47YWplZ6
z++ymK/poElhVccLVPVJGFQQ0GE+jbH3bQXdsfQAmi3piq93AwgjLHpKrBhfUVm5qIOdPgrCCgb8
TIvrAmCC1eLq34Svn4z8pujk6J09Vqx4E3hZLUo7TWCKCk2g4HnkXzsmL5EUGK6iq7yeMzy+v84y
K9rF2/tRlRcFlcP64jbq1w4v6rEIRBiJo6AQUkcdp8PGLmDzYqvvI7aIFGnYLrPXJrDi4x7i5OVw
iKRAuvIwZGWSx/JVZjVWtdIk2MY2y+aJ3L5c8W3vIWDeOV4LLjNZQEJFc62FnhRHL4YpwaKVFhl4
GvAy/sEa9mBP6UH7eIKZC9fNalrAccBTiRIa2lCWWI8Fx1MWICB0mJNTaSbSvGBXBJVKxzlK3sMo
Ra9sNZDC2tEwWT4uHNVWTCGvRa+fgSN6CEDdwQhAiEdKMu3CCL75sD5PkkJT6VsvCYsxTJbmYtiG
4YOSUMROT4BcbKqGCADBfZixGOm1L5ATzOkPOOQr+FX/7CcG/rc3TWWqPVCcC+aZ6XtthLqRJeA4
439ESaropwN9cVWIbpM/zx1q3V3uFctm40D0BRAShBpqwtjAV1eAOeE+JJ4U61zpgT93djMRwGwH
J6+ValLcQO0WhhAyYbuxygRjUzx9HLFa8MkT2tfw+FXvYCCzHNUIHwFvOSUZ5pOQbewvSMrvljS4
jqYANmNC56oKlZthZdDEWo81ZKhS88j3Vl2JmzM4R+jqUZoUZbaGq9e46N/tN08hN3kwZMOxrpIC
OHos7NxWXhvxeiJlspuav66a3n/mnRIa7LAf6XmLCveqz0+Id+QiZtOLfw96SlpbLZeLTp5PdGEt
dGTMAxrC0G0hSn4NlZOrYURqY847a6EAM5dDtQlCVE13u0YqWn9yphYoMEVpNR9022lRlpAsHzY/
NH7mP/ZTEc0Xukl4Sf2WEGh/LHBbYBvFFLJaofmubos/6NGXgUySlN6fsXdyGESodEqyl33HzTIO
MRvtxwg4icxN6BHrQ0Te9BByMngzZIHzXmrjAH2Qv8m9FlbroJ5yFcN32IY/CEGOD+JoXQbdjW0u
b/FKjhINOYyxw4j8HvKuIGa96kf4sksRO8sQ7U09KpksrmqfZ5Nw3vGUVIze8NRWrDMdmb2Eeo3x
UgDDvyrni30J2gOSggN+ddDAMmy1Mj5bx0AVaKs+YxErVUSlivN3/w9BP4Dar8KjkEOVE2jWg2iE
mXiOtO0ABw51wYB43LcUVKbhYaJGADKeqZOidCUxB4DuXRKvdIKpvi0xLvLVktFdUXXnJU2oAlYM
LLI/q+aSHkR+kA7Zc7GFco52aEy1lw25a5qomjBAbeJeyxcTOTiZsWSXrQrD2t2dMOyhIiG6YhNZ
Cm6a8CqLMUOtYITADgShOHNGFfRW8wfQGiOEmPfg2xMogx532UzEwZCWVI3rxU/VxiB8+sTdfeVc
bxQesmbPbUJejKHR4Pgqai+ulF+hIPXul1dkko6x87bz7HR4Fp3K/5FSXSvU3DkeRDt0ZjqfNlqR
yPVeFvC4JPjTS5A+7KSWeqoTesjjAWySoEcO4G3bVmOmNZj1cNPstsfGBXy5zRXIpsxefKp/33VD
CplJ06H+JNrYVBtO22pmsVVX+YGEP8GhJPSVjWB1qVoq5kyuHt8U5uKW+zn1aX7uxN6UNL9isG2V
ZxxvSffThMNvgg0qU3MdduqzP+fJV0y6Qxtk8i9+QjkI3c7rPmA0xTrJwmT3Rso+evsgBbqtjOSO
bx87jdcWVNONA5fdbOSyX2JoWpSu6UcIx6QnN5f1OCtBrH3jozxON42QMBnjsYSseBy/VEdyOzRh
E3rAR3ZLy3/FmjOybYnff796cS3xzZ2VQQpivyf1YsV5/aY3zvDfFgTqh6jhc+z8FMEkyieDmDwr
Gq2zHbWvX4qMOopEiYZVjHDd0G/T5utVGWq74j4xyJSuR1S80365b9Xxn0bDCcBZ0ATsju27n9xW
rYSihg038Q4ko0WWvmgL8ITILQWk6B1iQ/GrZmSzT3+L9QaKeKMCkV6kCadUIDYgG2ItUXjdlW91
iVW1Kq9ungb2pM6JwgXiXoZhA3KPjGecwQlt61nJTzw+CGoC4o7tQVkWet66SiBBY+3BzOEr9NHu
7SaIQfCh63z+M6TB3VK8BxGpuFngljmdNuQbS/UKDtWPhuMW+aNIplCjm6O5UQWl7DeGRSpiWr9p
VtHumZd6+8KyKEG84iwXjVsN2yVo10pYFfHiplciJ4HXZYoF2hAF21jzZE7HNmvISuTIgnpbosC4
2+42ZPMKQRkJ0ImoDPc6Yyx88iiiqgRW2hBiDBoZFzf9vu2qXrOWQ7CUGAlJ2He7vhQvuPLJhSnK
X4p5VvECqmmKmsWKPd2wP5pvqUjMNTKHcZlzSMZ4zFvQvHwUr5T9D3qsQyoLpEI3KKvwTsV/IDQ7
LUUCAiD1xlRDOycIyIyWk/bkGioaKpMwR+0HN+KwZ2iSvk1JRCxgY4tX07ZErwP9lNqXIX14RddP
MPp4GZCPTMWZGRsTuLS9DdXj98WHvV8dwxTGt18iCn/rYRM4kLu94Q+TsXComhv03RA6wWXpxkg1
LDRGxqJzMy4kacpKuyUdsmp9t4nrwgqVlTZtOaXoxFsJeCPEt/omhIaa3sWLAdHVcertHSJ0frtO
eeQClBp753MDP+ZiTzSNyHwp5u3cB/C/bxmEl5gGhSlEcp6HSyfeZ67SnHwDOBzNRp2hyxt8EuZC
PWqaBh4ZW9TBLD1c2LVVk9X83arosplNa2qRp7AX/yQoVsgZkrsYhtpnYIpZjexapz4tMVgz+fHT
3MRs1Xe9GXnhFM+logxtkMLHTBVnb9tKo0BtjLA+SIKOPjBDLgvoPYbLXT+lIGOatnhj5Ua/S4ZE
8a+DmmWUo/HWT0z1fwHOHhmLZkNhzT6P2mrOjc4+wUVZENIsfN6d5YZzPFHj0ihpTVcOhVVwHl5k
GrdtW6sYrbCw95eMNhMimywbFu4W2yfu4B3Px0hLWj7lW5zKD+YR7MbMUFuEdFIXphyZvdMWJkph
25lnnQ6PVvHlfiw2MuPrlhJkOSdgbcCU9EY6aP6/rVdwGveiD+yGSTxTXxJk335mnJdOPz06WuLA
XivYsjxTOhkSRbLrAjYsYTB7CRi8l3orpy7NTL84M14T9fUcwOoKwefwoEDrxYUEwPnIYeQ+e+Yp
wvVqD1o2Gw+9TzaFUaY2evVRdjKJp5zOk2vmz834c4DgNHRk1cF8M7dNRoqp7pfNv1DdKKGOMHKA
B6AYihyHTWsuzg2zNIMrqkuFvlJnbM7Gaqi/0GZHQpUhveumoepoyNB3R06ubwpFKoOfDIg3Z1Y8
97/TDUv9SnibuN2OZTK+Z+9QujFwu0UkRte5voR5+FKeC7WR3ja7pfT3TVTt1ju5EXNeOxy+hCVa
MaE7/7Lm52xH3QUFf6D0awFBpCul8vUjHlbzKPfwbc3N9+O5glZdEoTAlcOOrIUST0EVkptiLNI9
5MGBJPDhkf/nNihrzPDwbo6wZ6fmIKWW47vyakU03sMbXMWiFgvF0P+HsE/CIRtBO/3lWBHdg4+g
H+l0QSu1NhEQLuMrfbwjifmYK3r1IZHjU/JH/PL7URmEks4ZPnf/vLoKbsYsKoCznz0ZfZqmhlsi
dceKj5XsJZR1/feyhWfCFZjOrOh8gMdZHrlJOJozDK8lMvEXVuSXBWyUjMWT8iPYGg2Szg7LWwBy
Acc+I5iZ21mN6+COjr5jeXQJ1eYsfDXocCVkp9Ccoq/0E3ANHbStjzsi7BIXF5zfjkaCTZDxunU9
JFuTLexKIrJacdQerNYHNXP/ntpPZ69SDTW0IfprRwAyWOhEQvWeTfC4YEIyfg41msx+Nu5ydyFN
DxfDZA/AzgpKHtcABRefDakAySdD2mQPmJ4L6Qntw+Hz9IH/FVWS8rKs2HWGZwLbmOIMavCYo/fH
BeBsp+eiFTNXYsL1u0UfAkXQwDBlw66p3VpzcsUgHVAuB+y0XINkpFrPgyfcU2L/tk689qZOVk0I
CT0fai1F30b81U8iCAjoerdI3kjJJlpTYXzRKssjxQs+9G9OmXoEbGtxsL0tU0ZxVVFUqy8ldhSE
6syp0tJV0ce2OG0sGZ86hF2MxnY7ZTd9GgHWKX4ElpOztlHNFhJk3HnzFp0e70ex2B3VO89MgCZV
MhmaSbZFcT7HWefhgo51jeoHmck6lJK6JlT+z2r2JD7Zuf6rGU/CMH40WaDKGoqeEqxfoaU2ujzJ
Sjgf2lbb7JBP2MTgASC3BPyTrF24275/BcPnE2aLryQ8vVvQAv3/QFc9XQ4rM1Vd76J9hJlnoNdh
hPyXFk/XrRNxP4SbmD91kgXvPa5rEGSQ8SlXeawQdUM3eCdcCS4mQxeEhR/1EbzdedqGWAgofVXo
WANpnQ21xb9z/MLcUW4ta5zKBkK8taRqIVJ5mQw7Hy8w6qYzbvqASCvtolW+ck7O/95eAWZbVsYx
K3albB3xahCah7qGmpDzo7ypZlxZyYA0+SNeyPC+xsLIDBbh8nN9nno6pf5/LXr3NEFKTpqHJVf7
QI6TWR/guigIgRIrVSGJJk64kccADKISlRwSSgzQy4bnikpcHHbUNQnS4d5ae3crKZLCrpXfmYHl
Ug4ZaH7K7qnB+iGAIwANcQicS3ckcxGs/mnz1hftVstdHb2ClqqzBifRpO93+oXGADyS2xXhzEIu
sRL7MOsKn11F7XOGco/2JRItZoyiUdrGer7GjrXK6NTBWInplZQTVsTYTh5mN6giWQLrelWu/qi8
TCtZPTc9tWz5On2LoQj/08xfG72sl5AL0Ylik101jTVYZ3HZLV23OSPihjDJsA5DBwniuPWgd4Na
01yTqbk9Mr2oKAgyNRb4bZzAmp4aIPwT4iFwkuHTe/da/aMgzv23wJozCeGcoKc8CRDSe0VvOqi1
K9op+QZxvlqDeeirdFg8QcDgUbyZ/BiWrXOYfZPRL3fH6yF4LUjKJt+CTDQQppAi2TnRlGvJm+Ym
HmaWatCn8F10rGYd5tDBMmZ2C2M/MYRQffcrzKPp2wWT1FZLmCBNNXN9csOPvPt0/DyqkLYJTgD8
oq9Ek8ZSGQtNC3hA7SlImNADUQH/gNk0xf1I/KXmiqEfo6PhDmBl9wXivCxc9IwyhNMtMKBUKz8C
1l/B6wS70OOcjwV8nmMn+FavqZEPiI8AMKyCKUcH/0Vxk179Dc7iFxR4YNWLfQuJR6MKY40nHE8s
20lSGuoAMhDrhbtYRccaaVo5W+ifBGl7YK4nY0Jzy3TiBhA1+Es7Jbgfsox+8WZji2n+OGGOrrPd
6PABMXoCP7yChbpVHtDVyeemQpoA8I8JUlConl9UJ4WNYkwYuHaycAKgjqHLDtLggIHhN7ssx1tP
S5SFRXmh1BItlhs+lznwo8+7qI/xVp4amQOdkE+xZ4N4N78FcYfYBQh/9jA1vnwzSH6iVjV661s9
1HbESKr6qWu7hyMlV+v+rXuYzvCCpI/eHMDu7M2mDI+W6a10Cj1R2jYUdMgRdjcx0Aa7FWXboAE6
bfRNGO3joa8zard++5xyKyeFqzsbZefmcWkpY8OLJxgbFibfML3v5bYMm5iMjUWfjI6dJrlP3L+G
U8RiySk9oH4yCXsY56ZBdI2X4Sgj2K93v9WBneDMdNEbOSMOwALW9lE4m3vfKr7tRxBGMCDDhNOY
0AUzfLUdi3ssFG/EjCO9wK/aQLyhvpmOlUQkc47tnBgeEdk0uWkanmIfdJEozxfbJcfMcBwgn/d9
ot/hAsMgw4qGlLCs/BB7gSDZTV1qkFuXLz5BeWVK+8QPmMbakglOUqXBZb+O/Sx0X6e2fg7nosyM
ZEE74qFPfiSQE9BMxRWE/N/yodFB5kVwx2UDkmDJWzsSscTW1nx2NyOTon9j25wpD9AwCpEr8qDl
q5DeJTHNBu2nLABE/D0SPjg9IpKrqkE+byqm2Fk+epDXD0oAGYiKfIIxY+L/DDgyqGHoG/TxNtLi
vpRHJ28MQGPW6oDhXuoIU31pHKpwmTlGBGKc9zIt6ieWOR28/CxBBpDVCht7YKpWS4r32cXqjbqL
wGEy8adt+qy21nDlVZvMUsEh+YXYV8wCFUcOzkQl+47Mky6ZD1TzL6FnubPSQxblkTyo+OYXsoRG
+a7SvbWxf1Lyp8B4f/1zdLGJSaKg3qq71NCRa0C3iKHusFA2nRLRCw9LolT4pOr+hJ1F5kGS6egE
IYqvinLnvQL8xlqBYcJl6pHk1/th1uAfgKsisz1rGvsAXHfLi6DXbpPBn8aPpGXw0eAjc/3rw+DF
wZxCHxKyZtZaywTm0xZtMSuNBvRyy5pttunlbEbus/hp19ZSvsTGmm+kqcIA7LAv4vmeM66pint/
pl1ny7N1toADFdHPaGcq60MenTk9v07d8cZkYZ8HwcqFfVJdmEvIkYsevyyB7fjXtcosb7mwizSK
wrpkaqtXuAUzJI7SY99pT/X74efCsKmRybO8cS/QI/yB8r5T/QLNwHymvBBI8QNIZBjD/j7JY2HP
Cy15Gioo0rL/pAj7ddRIP6UmCDRZzFLenwpuvwZgrybNp8sjO2ERri6rlb3irm8ngD87cAF7NZg0
q6iDPhM75dSVtQkMwhYB2zrLtm2gXgUwGLng2HRzJ5oefx65RUlQ/vy9Z++KBVwIr+hzr1i7kofb
UbRRgLvF2EKT8AdEkFu1EbmIl51lCv5oYO2B65tlR2vDrVD5ovQvilLXXf71QnLBi9Hy87fKpRJ5
ho5Gow09ROTshw9D4jV2w87FWGOQeX9ffbMLW1/5yb1oOSSBIEo2bghCmJUb2GlsWqDusEqIJpRZ
X23j2yAPvSOMEq6iC4TgxS+CnNIwZLr1dke8xUr1f698o38Ti0shKERzmQDU7BUZgwOjsmIRdqjn
F4HHBJfQJdCNyG7f1DqXkKyHg/qjZSHJA8JPDWCnFGjRR70cf8Ftcb8IWC+2qA7GAa/48gaNYEuM
bk8nlWHx8E1UfjoOksND2k8ekbZ+nwBaxWUKl2N7SSoG4XoBm8UiIySjH/rE+iLEOzNxq4O47CgJ
UVSVW+HL5iV4SGgaGv3N67CzJumtpGKaNLycSlCgukGV73lWG7Kpw7e8siVTN9UlLGKibe/LPwTK
IBLPeKWjSLDcjkBtKzJ6ih07F/FossPWH9jzYMEa1++Oqhz/tK/aGCnCW0XiBHkbsFmXlt+YCt6W
y3Slddx6kqyXBVeixz+VpFnGGAPt/E4D5jjBdFwSn43T0F/hXh4cCyGJ6fcAaP2RejS7I9zO7zaH
Nirlqv9tWYwcaSb5enF6q2NMoQtqNgtA9db+7GZu4AEJh6r8hz2/zdgQPpl5V5D77anjcugbRoD5
kk0QAgHpSimRJZrK/4/ZnnY9tu1GH6fQNi+nkhQjSyyWVlo4jkPZdqM0akR3BVvIQiADFBMRi9XX
HX0sTq+6mRxegd5Wzw//LP7UcwWSdGy2z2zhPBzxV6IyFtemf55/pcEDiZevxzHokB14xve3uRr8
FJ9w2zTUX2gPmzfr/yJLg7cP/8gWlblYmeEH8Rc9gijf1tlSXvbGwSXFkeVkwSxScbbJdanuT9Mw
ucNRbxvYA/uzG09awJ+8OsHw4oL9DPtZbSGF+geO1SuVzKxLasVG3JQIZIOqrstLOkCGWb9vSGHS
YGanZWivO5Mb25GzZAEfqaW9k6eLvMhcMNO2wD5JtdYRaK9iHeak1pH0Arfl1gFjc2lEOza2qplH
6RiFo9EB7Z1ePfdp/4BMsQuJa5Natq3PfYZ6oJ4zQvp61HRmmB2sWRTpACHNzlFEa1eCnDyAYIyx
9WvPbcwXl0jzHodBo3xkXpTgJN7ka0mNXZl8zCcjhcK9+KerZCPl0MMN/905aZzwms4tpkyqqCrT
L8bzgROsZTLLA5dIV222WlifN9M1CTzcxcMvcLtXvhdQC9laDiyc2zvwo/XG+L+aqGYtRW4egSDD
mxp0+uEb98tDT7/YPWJaVs0vhaErnJWvd9a1fxcZwPxol8Oddwt7ySHsx9uz5u93PMjXqpRnV0zo
9/Nc989Xc9PD6kJqoNnguSW9+V28ZsSv3qS7BSvH/1SQNsREidkA2i7FRCEf877OjcyLjEdxnea3
CYrpVqIwZrfE8IyH9rC/vG1D5PNxmRL2JAjbpMu0a/0CJdQ5sureIeuXnOMDdLYcotpI7GkZeqyS
4ypq4XmQJNkQ61vA7gWxZNRw2X2J5cTM5lrfPAAtrLwf/4S2e3S9OOG6YNJhVIo7B5v5v5BMtxpY
2yRmpgObbtGtGmfBqsNkqxRpGBC21h+lNRYxiTkBVg8n6hITbOCf5KBBfBgasPmTr+vojQoUVh3t
MW1XywZwIQflYDNbGt326sORgK1L5zwUQNmlT0oXykVn125661Vp8QZgLcD/bH30bJ1mCcOGJ9+k
Ki14d/kRxeVsfPEG+7Algm6BPBmLpGKTwzvaP9l1NMcNUUlSRwOR5zQ6bZIJh5kUw+kZ/orfuk3l
9IEwrXrfZc9I0+CNH0E4c/vRN3978Tvet2XdaPq5cvJQphcgwtWa+/52gGgqyHl5QIeFfq5unX5k
whLoTNW9XgPqEfDHVun2n2Vwpf0gdSyiK7+6NkvJQWkzeK2cLRiaoSMe5S3fadLKLCl6U3xcdRlI
RCWJt6Lgai2MAjYPoLZM1x8Q/irPkS0PEEcKtEqhdXuxiSB/lOyYH9I3ymf8wAAisBPdWXyJ+Ry1
yjVqzgVu8rmxr0oX92Hvay1pNSJteOwega5Yf8F5RovpIUltn1fhJgKWUmvROQRrEB9+bfaXehX2
kx0eAUrSIqygPoUcE+Hg5vJi4+6x/10aT3Fgh3zgudsLPZY2y3/uVxP4A+DAuEfxifcuUY6ELIO5
59EFyYoFaqFAXBiqgwHSVwlgbSVuUEgWuEtkO1abu7q8yIBqU7a/FwJN2qtqydHhDNCC6VghFJFD
JDW9QV+C2A7bpCHRunbXqsViSj93TYBzcn7yWsWpZBsmixkrKEFDtJIteD887xsGOpF4F12Qdb51
RHQt6+/Hqkw8Z0MLgLgjQZtacPiJJYN2wUJ5O6rQDeMwotr8dlZfQP7Wj1CfRICuJl15OQIecBly
WN6ebhbCbWn0g7GMME/ILzi7cG85qQ6ZHS4mjJdsRNzjp0f8F+WF4JTK4HKFtrNpi2gdOk4RpxC6
jDuhr4o70p6Drh6qq7IWcPe7PQ9r4NHz7drb4jW97Qd2ViDUj6rHA6M/atQiWkqD0/f7/fWPyG4H
LWtI/PacvbQzTHm0j16PdnmWOM6IGT5vWhXS1ufp1igzzKp+OFHcwt33VsPcnA24VsULvzzHZxju
agaVGEcJyzXP+nHE3tVP5lwrdWou4xHsMHh42IM2MqO1y2JDFgJ7hJjFyNZDwPrDrWT5bLjdYdQs
zZjEUFy1EcA4Ek3orkHMTN/PIqbDDsNWwjSzxSMLJwJzWzUwgy9WiX1Vn6Vmg8XtFhQqH7lEB91I
F1Fo61WWp7bBRHEL/S4w9WfQ9sK5tp+VYvK3p1S0zvPPVfX37rKLzDdkkLLkIKSXr9bNhHHKBnsk
gTmMLX2QyVpBoaLqb5EeJEF4HUug3rlrbe9FRQl3A1HEfoLX47h4SZu7SmNOW45ZEdE0Z22uyCZs
B1Ee0Y5uA/xvZVNpyKcduRvo+HjTWzygXFFv+GxdISJKA5x8vcd9KXxkhjOlVzUpXkX59IYfrjTv
0SjTQNxWPhd3uUXc49s6FTCqh6Ob9XQc68tRAIipk9lqMpEl0RVEvsGZmIZtBWARsSwMx36vwc4E
wo2txSzXXw4iZ1TbDBe1cUMuIy/BA3OD8+/lwxwpEKyVTlxlFEDHx18FLfjxM8dJt4BXPo8R6pE2
VIeUsNcEVqkP/zKgz38LQ9Ubm4RSPClwUJRwj5OH5Rpv1QTWaNBsVa9mj1wD08Z0EFkDj27fqWfG
BAG0KWzev3Mqbr9+gFZYeRR5yLe61p/J/Q6AVWubBq4hwueEiu+FRVYS3EEvqPfltMZNncPuL1hu
1NL3fTods5ppGRA/fq1cWy95cTK0qNH7Q6DLB1jl342xMnEfQYCq/cO7P+gKTmcfTv5pSzZdZKXq
BhykhO1dh7/3mywaXgOHoAhlU0jC+KPH+VXdOiRPnz4eUFgMTYD/LTBf/9JqoGjIfk36C8RqAjS4
4VCmYNDnl14GDcAdTJcNy2mVDlJ7mPFi3kMyABt13h+u7aQZfG2InMx9xj6JcnRmal701w2O/oSI
e9Daul6LRfkG6p0OiikOk3pFSvRWXTZOBy2quPg6uwM2cnvGFnynRVPQB1/5cMlAoIxwL2q4ERn0
KSN1NvBdlOzh/ZI+psEPOi2KpDcYA9HdPDoyAJVO0bIIjKIabCkHd08Aw4WDQ0nbvg0v4myR/RNO
QZUaFanl4iRtf++naUWdEc00pLqXZLWC6+ot0GVaZV0f8JI5OO+39ipvfditaG/aKnerwmjO+ARD
Oz7/d9FJ2NGC8yFXJ+NqzSwHTdFVLRGNEAO0LVHIQWajqyzhcd4yh/2LAOuCvEHyf6nE1uPVU4h2
WzDSmdEnpCF7alrr8VpCPlKy5QzuQ9Du5PZ8bc3TvF11fvv0nCrlhxr7PW91PNDk/Yln4AIlv23F
2WBjn45JQqh0BQBbyujSp5xyD3T2XM8fHDxkWd0jFdRGbGct0lw7LtZUtjxA4QtFCnMXinprxZvy
rMqK9uyb+lFPzq/4c57zNklILPGsfKoiz39LgsMjLJarIVL+v/lf4tcgQYEiCXmHQC5vMrSU2biE
PFI/Z8Ab6Z7+RSmanU9DwWOa8Ub+M1ZTKLJNGOWY/E/YQSuv4NnnDu3EnDLXxrbwNDtUz8vjDmqh
vdxyHx4Ei6Izv/Jn7FVajmzd/KP8akoOSXmR65opKLNYAuZGj75u2v40MYolZ62elu/yfSBSUNc8
9dVfj9N2ADgx6cqHRJ5Je+JXnHAFKpsbRJaGnjR/2QYyuUmDIlboDn1RTqvUWDZd+UDmWjjHUdF0
7J1T/Ao/PtvROsCbP2mpfcbFGqMOPZuCQQCx8amhCg7qQqAgtPKKEVdHIVUf9OsSaa2KxlTbttGn
txzACY8AGM+ORNAUA+AWbX2jdwxk2HJoS/G/GTunBf9QkYtJ+kBBdel8wHR5lVXEcTKpaxSL5+S4
rxPZl4LMVSxT1MYKpj5G7jcL7XBnwz5gWj488hr+o42CrhwDq6R+SnEaUF0GHR3gI9dWVGqFjoVD
AWw2JvREDhDMbvzb7fLCFfSC+4YPJuLddq0ohK71vTAi2yjTmIo1Aoj1fpKiN9PkmfBubkSnjZQv
wHWiPO8rcah3QEkeucm5obpUzLChpW/I/QZzmcqBq498lVJ7Na7KUqRZrrnCdkXklgczikrYf89x
qursP9/g/3F+7m1Ng80y/Cttney087DsgxLNvgZgmCibFJRSzU3+/HAeOgELA9ZshW1EH65vxO4u
pjmXuzKQiY17kAGafJVc3qVwji8EqTqxBCuC3UFtRMlqf9QKy4GLwlrydqi9t4ebwjcpd+n/pVho
8Klze9Sx55CMDCqpNnaq/5s6a4EnZw/p3hT1a7an2d0xvbbNUuESf9z72n2mlGfN6b4saRA2pbtd
6MEI6WbrlEkSpqz7Hoy/eKu27OdnJmiVfIT0IDaKHxaPmtN2VXdzrlU7HUc6GEWUq+8jMfahMK7W
0vyQOqh8hR6YuO9Jw+ww4VL80uFfUWWKlq+PjjwzACHd9K8lqPmrzXvwOZ9JneS9j+P6rH8Ex5BN
vDaWkolOlukBxRp9NDRVnjo07tcxRTGgsIQ9fM6QNQ1+yheBiEaKTiP2646A9/ZpREe6hpEYzjs+
n1zxHGVRqRFG6Ti2e6lMhMgmXkxy+UurYs/mSgkFW4SKhrjDYiIrPtWpMoFlU+PKi3A0TdiKp5U4
44tXOwgNdrJ/wO3sM7hFykcOtWJX5/8kHowBdUcbSzBfSFGc5gz39scAstgXIJGRdnLSziugk0oA
BEgmdecBKtxG0bnJyNhftztWuI7Un226hPgbvpDO0pFwiSrekcq1e49gNIfPWOEBMGBi6ZCcW2iL
gTgP8PdeIZEsBWrE1i3GC0DfYgnQOph6yTDqdRHkSrHBRN3iFB9xGl7ct03q3nuj3i6Bt/DZpGfU
W5/e6r7v8KPZtJEmoRJoOWghDD5XR4hsgPOo3Gpg8UAH/4LkSd/FNg2mHTdvnJs2Kv2NPVPlkrsg
BeCEmC2+U13hHzXMgWfCvnPoqMagmWZjlVH57+/rwauVitDyPvApQJwj7u5NfdjKYTBo8euOHivs
fLyLASX3bcl70JYqu25QfE4DFZX0BpHzQyKj2r2f72OaIdEtnbRhd+vP98HVRT4qXvvprGNaIEc0
TMlf5fHDUIQjx8RSdY/sNYqmnqzx1LRpfuPsSBEMgwsDbKYHNLOjz4sBwWIcmpHykqn2QYHRhLLv
IL8sSwhBZuUT4YT5BYd5H4xY+fjE8iJNlHOoRtZzUTNPpKvFAxk/SrhOLPFd6kUwXZk9k3Y7jMIb
8IuXI4NFkWBEo7yXuiFDNGRoZ+66LtNI4xbLKuhNgfrhPfgXuKVtKPe056+STWo2l6gBi6N6Q6ZX
vCQlAEr5ZhlingeYLsk/fjV4DDAN2Qzii9naQq2lUVfQ40RNof5LsteG/C2Vf/xG+55ucV3fP2L7
b7mayVYbrsshaLpDxS5GIryl0e6xYU+MVrrLXUwmvNask4/elMH9TlTaqjxd+vbye/6hCCbRfPbg
LWfmqr5YrdcLf2JQJfVdnuLEtvXZNFVLn6AZlxTVxDcB1+S+aVcVGSX+b8diJs0ItCPNRnRw/3Df
4de7xmIjYPb+PbALlKDb2fte2Bcejr9fk+IQONnxd3xXwkHy3pJR4x/uckaUA6m0yrFgw1uBYjdy
UnzOZce2n/qQ+cIvQXkPKaMyTLcgRf9XmUDZVudZXc4ZxRDM3m82cRkNaQ3TDcgtLBBbHUdogZHw
TLkO2J78zJlldnkjtd2C0km0yIw+avRCj5/gFXBoC+ROuwv3fBl5WWpZLbPKGUPvOY0wFYwS1Fv3
wyIHhSlkhUVoSOB1Lva79eudjF5MQ6rvOE3W5kMrS29C4JdAcVn9AUZiVI3/QUcLOAgqFla3OvD8
NLsNu9Josrfdn0fKrCa82qUiESIkNSs+/3t1QGBoMCiiIBm1QB3UoJkSOfvbDKJDSvU1HFfyaiH3
MF4oLc7R2xFvQ1hXdErMlmr45RqdFbA0Itl5HcCexjsvgKuDXnMOlJEjwsXDjkPk3Xf8z12atMrd
75+hZ7DPaeS6NtgxS+CaZmZmHgrdaLaVRCA6UytFneQiaPrWaFzfaFZ5LXllm629Wbj4kn8dzmmb
hRvv6OFukMmLBtlnIgy4NTp1xdjspp6WjKjHufv6QWRuy1hFV2sxC6GP8iFjYrtHddjFfNu1c/YF
Spf1S/5fJzGka2+gm0SVGNxgYMyqt3sFgc6JwMS+g6nMqgS1Y8b4jSG9QpRJSq/bLCXWIDPy5kio
1MFN0f2CaCyheKcEg47gzUjl9xNk47HjiJsAhhOQ7srtrmee04pUgo+mJcfqWFUB+kdNnAH/Xf0f
zY6TiScJ+ryIkVsymYwQtErbdMRhE5icNxGrSN3xxIt3FawsbRGuHAl0/UJp5TGwu+Vm4vjzR7C/
8CxGk08u+TrjhVJcAk3bSHH0UdgnJ7QBtR1u6ViR4lH2EZ6DEO3JqOPcc+DvlCgm2GkBW8hNi1Tx
mL4E95rd0SIrRgkqi09h5M3MEGSgWdW+ttwfM3bo4mC3HZwWExJV4HvJXYtJmjZ+Ks5L4mpXzbGh
AsfmB9LKtVFV3FB9VRSNDlwrqc3eLQsQ9LjC/lizz3StX+ehFd+gcO0RwNyAf6OfAx/W2foxyWgG
+yjKWBTiyrxiJhU4euLKQ3NTP16xO1Bc72LsD8zkijXYtyt5Zsxi8rL55XxuLbqLYC0MUqb4YdCC
Bb5RHaJTQ1bg9Db+T5svD2lCkVAjUZhHXrs/EkjzL3YVkwj20oLggYOo2ukgNunRfWiDp84I69na
pJ2K1jFqr4Z3ZNVCvI6pHdlW1bcZHWa8ASIAjm6IjJCBWRj6KDnbGek4vDL+pKK/KwVrkwCYSiA1
l6XDaVFMZq5nDXF79V/8nPX9Y2Exr1F/u5xnvAX/EZOUQcvmBWG1ddANTDCJXIi4vVcOuSNuv36X
yk6IVtreQAF6nDGYSg+FeXMc+U7D8gCRgOxKZhhuE0zfGkE2V+Hl4ZGLO8rorAc2JhnCzorfotE8
HK/C8kK2qyEsoxWP/EzhG97UQWM/35KW5AudNsUDGgFnDtCcHSq7gksU0Cs+ElujSNCBX0PZaczX
e4/xk5Zjc2hq/zXhWpx0y5rPhh0uj7pkQQJYv+qBA1dHY0kVXJ+9oMvwwpiPqlwN4jB68MKXOtDk
zFa3i+eOm1GMGNSRhdZV1tT+1Kgzo+pAfVzwkb0Ir+SQOySsbbBdoq1Lzy7x3rXhZs03STkkXRH3
CM+KFMMpIFrWrxPUL5jYrL6dxoe/f4PDRtoLehR2swPLOmxgE0HTHPej38TBl6kVHF5DU47t3em4
Mh9/ts63EyFzjFL2Xij2Qd5wF4XCIpN4bKorUo1CFf7a3xB+JvOHny6Wu6CT2iwQet6ZVLSwYmbS
LYD2pDmjIaF1TESRiwprQ2wxQrwoJbvc2IxFp4zks675474ZRYhT5Ld3V9uz33+Ei5/uhTSTiz91
GxwFVch/W50NVioHyDDfQQY5rwoKtuMyj1Ople0ngR9zCy2Ax+dwi8X5g07dmoruOqckEffKwmSZ
IFuGkn/9sdRmg6fSPS0S++LEcki9eqC44g/ddXVhiY1uKvIbopMCj2Bv+6iQbPlYgUFyx5dtNKsb
1JXLYlZIaPruWAZ4GqY/6VUQC27QiSs5b7QI7JkOqNQMJJkUw0igPn2wDuqrZDeobkhav53Lilxc
B4tWnKIADo9T+/75ocUwPQr5Gr6lASsvbCW7Kf8fYfRTpuqfMCWGqUm58zbs3GjNuQepdP3u5GVq
6XW89xI5/ZQFZxr3cbVJ70JzFfWFmXJZ5b+HQvfwUookB15jKyxOWWwakKiDRivhja5fW8TYUS/W
kC7uwnR2htKvcgCl/tYqCVOKomUmVDKMwpf4t6Y+CBIjvVXTN2NuIUrY+N3+rYVvCGK52c87kNwS
pj32uk9AyPoOjfbl/eR1VQIWJHLOoSk+uInKIYuKSswN0+6wEwlxzW+zXIx0e4NBR+dtCLtOmYfX
Z4ZAmtdHEKnwLQFFuizKi/q1Bhjhzs2PfAxa1wPM1JuYVmborUewYw0rA8TvgiwXaZEdKrD93w+P
0MDnBCoKpt2DbU3QB24q9WfyUCQDJ/EywTyXikxdJKgG3V1F9Y/ChoN5urGIUEZFkJtJDiRpWADL
dUgAoMg6eFsYRnILfHpIh9txIkeRa5NlY/YA4H+zUhitBab++LhFdp8PQCI69q5mrbECEXZ8RZrE
8swWx1myt+N23el7Dvo1ka9wyubEGwOSno+5YUl8RAgS+z+pciKGAbaG4+XK/e9CFvHzGK5Yzzv2
3rgzP+v7KyYyQRVmXJgPDsjhf5idcAEEgF3frKsgWx33Ilqje+DyivUJB674cpj1+a8ik0aiF/YD
ULmi1JoIFHDOYE9iSdubPVbVBvNoY4hMuHnmpHx3xKTf0Y3SDOb5WM2waj5SPt0HYOdHck56A+U/
0VecZwUbiHeNveOsTmeLWyTd7cx7EvX2BhXin4LnRgpLvBZCfVbSgVzf/tN3ROEwuxocgKFfmpKe
JUd7g4HihEjdBAfWwWXWgwx3TLYbr6fjvQ9fMWOQGW0/iIFBbEjO60GxIccGSHurct1xZuJvQ3up
ikATjzFPmEkh5Gp+9ldoEqTnGkQS2S6sZfmVpBkXZ1g+/to4PAYgMn2lF0E61IiPgUDi7bChpI/W
OvamxANjSNioekN7OVPpJYSE70ki92d8wKlU2DJgjhwLpRytMy5Dn451u88Ti6o06uHrqkOHJR0T
qnvyIlWZSxtulV737HVhFq6zG32M36YM+rpO7Hz9+8mApOPuBdrZ0oWKOFoPsFe7YMb1K7uAAx1u
xhaVyNKQSFORprfdNN/JQRNQ8Y8xbS+I7kP49kZ53QX4HnpG+O5+adQZuVcU0yVKxPewj1PkY3kv
m7Xvoc6FDqZhTKhfqO1RaKZZUZb4p7vcCLSNWoQRkFpfazbW5Ukg3Iq8IYX2i//4Ef3Zeva0Yp27
QuD7sCX6GQfVeu3zUjgXB0iwUPvRQ21yqZjc4PXsHtyBYS9viLc60SK+RYoAnFhzp2iyQuEMve6+
N3DlaFw9/fGrSgjq5Eq+SQ2k2WZV/gyMrABrS3+pW4QOfO3wGiUjHDA38Gv+iiuvYDBv9/Pu4+78
yTBQQKI/nw09PDiPYwiO9lA3MpS9IvKLmiLizXRwAHYjZHW5PaHVKaHDQpuNtttPqEUgXIvKUCZy
XgFAU/ODgyogSybcqhz0/m5mWt/dkDGS7oURd7i2zSAaev+5yl269MH+Ph+gtqjSitn1Cn5UArJJ
E5//4bEbxgZRd7diXP0TiX8U3ndnr8saGi0tuSdZ8bXHbieyoaskZ0u8Bl+z/STiDzX6tMOfVAKo
lbXdnINHyd8UeT5MkqJecJGCmMvwg/q1rb+yAFeGQeWRv92MlbzLiQobM1bTZUfQJOttWue5yFMf
Oyg6ncv6VLosHNC9kxUwMk7Qp9Hpr9wVFFdpcRqgKN65hPiq0nrEN8uHPR8lO2K04I2xSqec6CRd
EsnKcp0x8X/h6mGneBgbhQe7ip3Oc8Q8mtYh+tafjZ/sB5W2ZgS2NLtzkuGSaaI52KJn3Ddn5UyG
YY0LF6Ghkr+NAj5/8CCbizisgWmj4Df09pyWbqkItnmxDyxlVBg1e0D0lGU1ppCg6yZLOtVmb4I4
vgrxIpvVAlThoYwDad0qJhfpLIuKSPQ62CNAeq0TU2kOCisLEwq8KZcFC6xSIp7OXxo1bCGlCFWQ
6wWj867mPj9Xvq5HcJBP80xalZ/tOEz3iinRMI2NGBmHYLTZVeZr/8ZLLHV7Z1LBELJXQKulHNRB
eVtCxpk0U9xOSy0cRgPOjsLYrAGG9+ugn/vJbHehuBRF7PrifXpxFzQrtUgWpp4ujXjPO80fYb/N
4NSQ4IS7+pGQKjCCbA2ghk83LyXvwihquJcRQHpyKOmbwGngXpRqcSheQV4tYPg7a4uTfsqwxhcE
qlzfhCQ4DMdRfVeTp1kpYo2Zho4XMr8pPadUTs5F8JrGuNPEJdAHw02WNwP/CdrtcsGstJDdyj9f
O+xfOZbqjg+5ug6nvHcHDnnj150ajFq8US/ephRZ0B6q9TSI5lilSgiQC1ba22H2WEwnNtjjCwxM
F0/FGXFqzzE+cHIAhssjTI9EvIJOH861CS3rv+KG0bHZwC/clGiT/dAfZQIDcD7olzrm35R+MbqP
7sjYYYjaSIsT87LP+x3OeyxlpFQeSJsS3wdGrq3+JmLEzpi6GEfcmSz+WCpRYjFL/37pN6Eqa9ap
aNdxO9nn+15gT+8Sj/vyrOxz++SzIEQiFudGUniYmUNpjrNchQRl/YqWSd/C7ceWYu4TgKmb8BUA
57B8YBmEEwQnqBKHXVe3Y45XtIZrFlC32JaimPeC4FMl1QkaTgIru3r8EgwEaCPX88td0UMbnfE/
t/woZYmScJYEgH+xXf4JF3LntjP0GQSPDOTPL1A1KnX2k6SXzokkeMIMgU0YWoWpRpSAij9VzlfL
hUC05DtwmTtpRFdJ5hI67cyUshZmz6CpvETbRra5q2efioA4LqdunGUPMmT2PJ0EDG5fSVkjD40C
33ml1mdmGlQ3skvkGGkzDgY1MrDzNL9lGuoEVSWu/7Rx+CI9mYt9Qu+qAdyHDnTmK83hrl+j9K5r
E0d9hBuyuGbwzwwGVGiBxmjmUV+ZnIHs00w2iPqhQV4j2mHbYnzfEArMKfmu1MKn24Klli7uhLCd
UxoNiocuupmQphCgFC6t8GJcSWjXukjkdgfC0YGZrkUa8OIw9ri1rYrmYsycYj99F9YoHYSNHiLD
sqIkoAeMXbCiM+Gs5DtW5L1iNyqpwVtURnZzFGnRuuyOSXhJIRo5yVcaE/Dg2whrvrYtZ3R8sREF
KmDQNwGFuU6AV7wFzj/Vz8ABzRP6zdSkXTE052h1LisGqbyw8fmuFMNkOBQz5Qo/ZOXqX4MQ2xA1
uYRWq4g0sUo6VYnuPOOt/Mu4fjRa9WQDRKbGVxtDO8Gf1aFsVsfAg/zugjtxN5MrLvHGhfI/dGkp
jpaogo0N60i1QkX8KVl/atyRkYvjxdfuS9Ztbuz7a3TQTgGolXL+KlVOJkF3hlEVZc8QF/MISION
T7ou6RO7a1otBaeXavNqSC77BDRThW2qjwWcG487QoPJRikA1hgCVxr+WDBCKbWipiNotfKgo6DB
aboSxQ5v4LSrpFnsATlyGupl82WbvGVR5CJTG9lfAi3eLUKCpEuyZKpdPmlQSyiHK99ZgREq/jLN
Fn4fpiSc8b454JFgA50nV4BhfCOJbahjaMZk0FWXvxbtHCmamLM1lKvflmw5HRvFX55QZAAR+nM4
aznhdMh+jsu4rzcXlXLlb0LdD26xFq5jP+inAIicOMZBOqJlQLjlBdcLVNYifeLF1CKVgDsD+GWs
jUnCztsZw9ZPEvtS9IptNgaUacJMBOtzuNuo87hGMyFjxLDhJ0etXqZx4XBh5U1O8m6Rl8whx/FQ
1WuJv9i87J6LC6k6HG1yE1oJgQ5AHx0YxnQKYcSnHUlUpf184v8SwN3DPaMjEh3+fe61DXuPEMVS
OjjRq0hyjJClbADG72yq7B3D94atUAeEuiFOnlaa6avE7ewsXfKrJTbosqBaA3yQljwkQuJEoQQS
0DqWUZKJOQy0Ji1/IOsWgJ70WwmFrV5gBAazN6qiKL8FOzD2VJmgr8UD1OknVuUo6jwpS9ONHeXW
lIPetpld33wbMjlFYzn2ca52g73tBBUlgKfRvOO6ttRS4uaypTGaKWF9dJba3BM4DudYFXV7L+rw
ReqkvStEul1CRFEjrMrJn5lww2T7GKAtaQdRPW5YhP6y7YP9slHszNOpCt4RBVov06pXeQNec9oR
nzNy+hE3jaUrKFzf8D8OfTHCONEOs1UEybFXte2NQluw/mrC0E4YfKM62qtUzucOPvjkj73PN+hs
GzBfZ+uhiWBZhFuTCBXbEApC/BnzhZ2h9eBLkbViCtbDgNkrVxx6qPcYz6xARYQshh+kF95SBolg
Az4qLbPpnd4xeFDxtIRXE618z+zSg9U5W67S97lv7niDhZwb4gKkXK114CvosYDELKmPEOoYCdAv
MOEwt2h8DPb65qnB8Qv0abIKmfixIOUEEEz3XQ0JjA4rrTKdZn90fJzp5m6yRz78FmIq97kr6mTD
v7bpfb4TDEyMcC3wH0ZXXd0JTcMDh6sLDK6UeSpCigGxfxZRbMy/PLAz1w51vTnmiU6CIMBm5nNz
LW+8ak+INDy54pxTG7jHJoRiuoFLG/q+GroXkTfYJ8vQg26p3/UQayhxjOKMZSREzfOeT+jYsvBc
+/8pgFNPCbAzW55ELHmhmYl07CaRELFZ/BK2dKdZ29b29ygGNNzBuW86qtOUkssFXg3WFo1WkzxS
jh32fYX4G5e3Mcs7iU3g6JE68RIrFZfp9dRkbikiZZv6cm3DL01diOhJqpnW6EfUkDt2k+hivPVT
hXTr9ApUuNvwyWinTh9YM+gfuYCToDnS4OcPRxuBaLo7IYOResXvR7CiHuE7ogwDuCs+cbR0h49w
R1nJZbyVjiQuucpVRnyNyJ0tcAxXJqV0zRdZOY2kUod9JVcBzCFo9AegKh8edllSuOeoFQPudUja
mhFPiXnoF9ZYlVpjEd+oW95ndKjGsqor2ggnnazdtAAk9wsrkBTU3s84ubFUb5+VDaFYKFkfeVis
eYsikuUKv6OJBXdOIAPZIkrq9UyC2CXFGz/vj2dfIRjam8fRgts0gYyWTutXP1nQstDZjAsJxZ0R
to6DxJAOAvsQnLlG1XHH44O3QgL/HVotFyPIL2PxFTiS3+uOeSGZufXH6Ps86tM3xvEGJejmD77W
vk3VF+cKbhdt2yIEln1S4cG1vSHyM/p+YsIlxgIEwznVUBzTk0K5UnzaOj/AHo7Z7iQPtTJkt7sE
ayoq5dFVdBgAr3lCP1B+0tQ68D4WdiA4bX136GiRy8vuXzc0Wvb3ycm9vKEBHPuShLxCbQ7lD2Fg
/FvuZyrXsaa1Bs1t6V8z5BKh98ZlqdAPXpRx64JQ90nK7DF/pnN282UG1HUy6dHFHvE2e1jqDtAo
igOxI/cmYrNhxcsXBhVtqeSRRSsEe3vXhU4Mx0A0BziW2Tg42dpxrZrMVtfb+9UKA1d6bvMkGdqo
gGxRyMuVvlnqA94t8lJYFsbywaNruXL7gl7OxEpfd9dHOWaE40FQMG/brFRvMjmK69KuCsjRw9+L
PjQLLG933KGZ93h/C+m91C8nQg5wfPWgTvDTNxaJbD2SddICNsbtLc3gceMqQcxE6NBYsqfaFLny
Yw7xtJwZnB142OORLaCwTVXrlXOXZSMXyULhUd+hXbyqBaLmskPcpIdT1HF92KncZQL1iEJ6/79f
LRTgoWpPkYrgjU4CJDIsF7OCtwEhP497M9gej6zbyLi+ExLkO3j6zIYzUgIiV6X52KxRjenyOByg
qGM1/VN5ppBoGyYOgAf5R8igtsm5oEUqw7rYD8srzLF9eG1dx4vXmv/KsxulkCngM47jad177IqN
QaiHtqY9OYQIBvnWbJEwbzsLJLkGZ4nj8Ev6lOV4WPmAMFlahiBSs5Fe7mXKdGlYQqoVveo2AaJe
eKN0VPd17vQ3vmofCOTrAqdpbsC0maDcld31xlbWYOcAM5snomxD1WeBSomUfQB4XWPubJ83hRg8
LUK2PS7HkNjPhxrHxPZVMXRjQ20h10iGtzlPoPdM/0W9dk2b5M+J7uzMKX5OH7lFdcErv8ncVfeo
40n1OzZnRqS7K2oP485m3Gd9Z/tMz1YyVQFrbqK3h/jasUH5BNXo6wXqLbJC6osAyAQ+70xoC20F
YemDbvV1m/xiYj5jByoiiSLBM+vXIzDJq0hc3VlO3z5Rf8LjalzjfFwwOtqFr6DN7EntDLvfBCZk
/xDraaKFYDQbn6K14OhJOURFesEqDBTgz8pp576Y/JqJdagLaolY6WZYfO5AQE1hkbiJf3bUguUb
GxwErVBUcyMWhnNXE10HMM+WPze5SB6XnFiEAdiEArb5mRREPGGlxeNI0sQOl9GBqNN1zmuJ7He8
c4QRCJdJHp5QQe/Tq8n4DWsUEaao4PmluRChvw865Q63jk+gz6oU10OqJY3e+7J4nOo0xYfwA5N+
UYqSaozRzyP4kVJ1VRTO1S8bsrZzeuS3dAYkJbWqJ8AmIfhwxuRTsj0Vz00npEP4VA8TR0gokn3N
Vvmep400/felSRjVeyuozaYZ1mOpPC/bGoRHU7iX2JhShFApIMsu026iGFs0AHpcHmpPrwvzpFMF
PcH91h8KDpJhAW5gs7KLFc2KSiCi6DbiBYWqLss2YXN5U7nw6pYTLxM+LQMNV4lE70q25Cun9bSV
Gqa10Mn2iYB4E94EeM8hMqYbdTt/D6cH4/pXTt+sfPz1eeF6GaNYrEsgv75HifWwgLw6tN2WJbLk
TZT/SyYJjEVTMWHIErDOV7qL4ZrwAxqwAFA3jwWmBgIg1+oCmAQ7Ny3JnWeuULpTPzrBRU+Y0qYo
/GftrZjvAhBWlrkZx9bu8AS1cuJ1h2libahTazYnH8MFqqPUC9vXdK0+gPAU9NJjfhZgRSsGOCRH
5vouxSjJmhT6V5ycNCy0DHM1/gOKPhjy3WwLIazEgV61TZSMmyiAGL48KSzvA5p/WSo4bwKWmGci
q+yB/obX4VLk2lSNwBmeLvYlJpkBrWHCroE2S/11fpx1MLt6gAU1kdHEte9JV5Ed4wefypFOi4kk
8zc+8CGKG1+aM8m+bYanQDly/Zu50llPXQUNmnEjtkyvFcWoHXQt+fHXTIpO8wIi2m0IDkVwVGyA
gIBtwsiPB6JALzHdj8ptktrn3VFyEVNoeA2FEBgg5QypnL0hlWyFgGUOgu7rbmq8uF527RzHk+c7
jk1N49Z2sOdsUf8ZKSEcGfcaXhKhEk0kRTKyL8RgAiwWylmxfr+nGJAKYanFbnYSEib0d5vVyUXv
a4ghcf5fk59tIlLnKgHvEJahxo29G7Cl/mg+tdey9jgEV5rVgQk6db53IEAnm1d+wjdj7+ofakAy
LELypj8zOXtb8Qcqzv9Pc8dPZiTe5USl+cBhcuJhfullr2wOab1+jWqH3gtvfl8yesVUF9jDDfBP
wjl/Q3x7iY0K6dLuOpnlMDLn6MS4R4t33+uKTbFrrLi6kW16RCpeKcHYVWeBD3mrsvvbQOdoykeJ
mMFpkaCMRnZnoNixYxIeLSI+Ifx/HE80FONRBD6NhuEupx2cZst5PGZ1jgYGgG9KX8JxW4gl+q3l
QI0VFXSdiFl4MuOcDSLqlxXtzeNDVA60Tl41QJNaCjDvGYhxNBfXrp9/xeDgbWE03F591ZMEGSOQ
+o8ymxc+1oiUUOCUmsBWfL1sLck8zJL23mbr8TImxIU5MXFh2P26LQFide+0TvLDK6NvtZmvL7xG
EH6GbiWuzd0+M1BhOm01xWP0Wek541FJ0Ce/7yujRKygdnSvAiaG9nrTU5jdCizclLXOAZXJT7Gv
EiROCrZ0Ob9HVnCfctXChNZ9TIUaxbvXdDb2f/qtJYypkmCyE1ztjto4LEGsLU7WTnOlR6Xfy2cZ
tyANr6PKEvliDfKdHmE3YFlYbQ1Ml82Oxgb9R+cQvuFsAYABUoJZVhuJh+MxZKk/+J/ycQkA55Ze
ZE0yKiqxJWgSq/kdpAmf0zkVR978WPkqd7wDYRhKJ9vmlRllzFfQjb+3ynfPkGwl799J2kQ9LEKR
Fax2m+qqOVqpzldgMgR5iA55r9DKmekBBcdU/k2TaOOOEtNym8fdk7tPmeS6DNttD8ozPbmkVpPy
hysFRVYKQNmn/GMw2Zh3BOp17Z25xuknbJRd0Uu+l+RBeVA1tJDjcU3XGaVQGRnYRYpEi265nkY0
9K0NbQpu5iC+WStvu4FkBjkWCRFF7Sa+5LWkV9cicaZ17Vz6NhFx+jK9R5Ayx01+uJIjAHW93j0n
gO5cHdWCREoY7B/UTUrZbNFVqvOgPCo3WUCmMX33moLz++df5HMnKhrLzVmnu3IWHZlxNEczZIwT
cemqg3t5p36Wk9EA+cSL2yEbTSbpPantPGSHkagr3LVA1flG+v/FMSApGyV5biO5w/Rf82gMQeIW
qkIeswX7xsEvflXn/tKTwNMxfeXFak+IevQQ3JXkkTS9vsA1kcGoVqGTltuFkfqAKadcmXR7wW+q
sF/Wy1Hf2zXmmg7Jylhszps7WxBMwTpajLVPt1MRaNYBtJ38xLRoWqmvkXs2uncPkAPihmMqlVOA
JxYOqosnv8JjQ4+hmC+s782Ze4hNrRWt64spPZJ9iBZ4gh6RdvlXpru1k6bFmcC+1p2nf8RKqoFG
e3DffM8k5qA14P1TIkNpGZdm4mVhfiiign5DwOGByXqWUHqNNWke3P900sVKPGmVaLWxOJRSZIC2
MHiT8tpugQXWzzztil9tmNiPZFy68kwhVfQP45a4zKKjh4WMjFjLsPkmJ+DVABjZjEbzUZY61tkw
NeXyH1W7kf/3o3siYVGo2v+Ml+I/cn0PH3dXhK/WdqVh60lKvPhWwhDBA8FbRxzKNXlPQdy5pfL8
FpA7cGlSsGJcyy74Vlgu83vtYEkytV9VRFLiBdLmuyMTp1TU3gS9EEACrqH9ao7lMM3gy9GmmpJ2
dwot8435sMUJGhbIU4GreYWyr3wk0iDo7k3XJw7+W0cCqJor3TAHxJNb369ZRBR0qrkB975VKz9B
BY2WQn2SJa4V8J29LyoDUpK8wjPY6s5rs2qS0Pa+g2XjPDEo78/DnK9ZZMbDNBwq+cxCL99ragBz
WZyujrQOAR5qfp0d5cmTNQEqTZlX7vnkuKqRYL/GTX/ShKLHfikeqBrdG+RShoBxsFMRew+r1XV7
qbISrjZvNh3iqXnJYuNg4L/6/iROxkTFFXUvrZIKvYKEmOtBJoRO8pA0tmdCdAyyqRBAL03PiCu7
WfbR20aLeNbPFJPPWyT33O2TdRwsVtl6JqOjzGx03BPdZQzntX9dbDhmnfsOcN3gPXwh/y7SoL49
j8slFmOQ7jMJ4UiPoN9UqZEKciItt/TqeGnc5k+3OvYC9lHA1nVP4Q6i2GJScUZ4sSNJEcJj6QHP
9/3i4BSLCjE2wQoAn78JX6bOB9zqrEtN4u7NGOQsGon650Gm8DZEZ1JHVpV0uraQVW9kgKtq21Ht
NMMUVMHCfaesrqJ+Hv9rG0n6cx1k/MGcNyZBrF+SxmusTe5Lczkiy/274xhRccaCv+2gijy2GTuV
u9mGlUgTtAZGGrLzAsXbRU53HtSkJUSDYK65ahoUGxFXSU9IImx/vbfSyQmp9VJb58QAH6Jct4Qu
HC09Nd8A1RQ/RmJXgEsyB41/vWIvqwMKn8Xv6iUaE5txTgXjOxT5zrmkojwM9XBI0Uw7vbQ2OP5v
a9/IUKmhBDz5Qq+c68u2m6Q6/qytFpMylBSm1EwZF0xqboAm1L0wZO2KczH4r9iIyMzKGk2Ff8t1
V7ONT8yu2/cRycOUywYeJDQcL+WaPuQ6pZQWwqEC+vFDZx0O5B37oqz7pMYViDtoVZpy7LdtLBEQ
+QZVnb7x08nCg+l+pZKa0HjQdqgw+PdaWtsu76bL33Oz0WMX3omrK7PYC3Jw/Tkp8oyJ4mbqGF5f
GpCDVLVU/TpneZZYOK+l1dbGPVFHVbpgs+4poi8VNSCh/cFmwJbazTfF21RNm03SlRliZGpI4oe9
/73Ub1dcYD3diKCdY8lks3avC3UyUT3OQqyxlEtCJtbaAj0HntalA6sSYZXhr8EUj3BsWC+K/qP4
WwqKGmfXQ2rsFtq1gCCA9uzj4AH6B5zpc4xRNbAsD0zid6WihfCn0V8Kydg8ScNi1Jv6yFN8INc/
MLZ2RI9+r3WpL9UeH7XsUdFJRVem1VN+Y7NVE0MzmsUWE7rLrTwxA1fN05ZBE0K5agKD/wH65B8E
3stj2SXt415eU6zvusHvuFJnGtxXvua2rpord0BjDcMgXdzUyJ5bcIWPqiV6J5ia7hQYbRRdIzYd
KvW3Q598ujXe6/CzfaOlGpF1e+xzzXdOp+bQNF/+aK9Xb011SyxcFeWPJ5C3c0fT7hzDAT81W+2h
d79ByQcGf7t7QF3UxxOjL9N8C9SwgaTm3Kb0PseqmYkduhqogQUM2hQzHWmRbeXut+04aHKS1KJV
AGHScmLDoUnFy9iWZuoKAC/HoAce7luyEnWqr7fOVC1MkPRopst2GBvNRUv/f8mXTBpZUe3CyEJG
SCvsBDFLRndtiGUW4byrqm+w0hwklhZ73aXFd0YT4RLEUsBlD+hp8AhIHpH5IHLDCmSoY6ednViV
Wsr1eciMhV3R5smU1tH8RSVTVTtDIPsXb49QC2tKCCUIXs5i0Jx8jddOb4slPX7kOTzaVAwH38O9
1itjXOaAamRxodvtdPN3yUgzWph/HX1oEbaW26KIRJXcVfHWj/eQisFv4NmdaeF/EHVdg/4eRzve
2FwvfvpmAVoahYbrRarjeIzSV58bToBFw+rZTFvypso8U+H/TSJ8D76RH2tjgl4R6A7BgYUpuIW/
qUVxE0dzIsp2nPgsQRkRGQXebfLU1m+PxcbWY8pL6dHs77kH1zx0CPhiuaQgunksTAsDdeStFI07
afU0QFnCPHMLoH9BMZtKi7ZZh78ZbiSccNmudU3Cp6BgZHhVyx0nYPbbxagGSoWFBpDwrJ3RSCgB
6oXqN1qSqhPEiYI0L1BSUSPb2H3BdLrzMqiKXODdlbnMkXY7ru4Z7qbF+wA2gsvlNnovPXzZHGYF
uD17ITiBtlFtbl3VMTVXWAYBQmjwAES25v1xAjf8Dmq8HnplqE2uS6BhkgJhSOtM/HdI4IdyEH27
+E6jkUFMFwqwSjP0EvhSiM+r6mITVp+H+nrONKkrk1CA1dGBQBCaTQ0R01gZ/gL05vlXsf7nEib6
kTfjeA7tADiwyQ8ReEvSa3VDec0WNN+5b4dZSFSH1n2M9MIk3YwwS219BrGipQyLWbnHBHyHtfOI
NA11dfBfSY15kuUnXqS6L3wRvpiPoTEBnyOBZl5tSbax1C+vjBfMLuZyTnHAFjUil3+J/B9PGLhX
EJCG5lxQKh3Z4hJGkkKxfBkoEA+DTB3YPOhJe+T1WsTtU+8nBE4FQsQMZHDFmoH8r/i2VIP61gcs
cTdKfvUoSM+iJsyy1ONnM3GOfzYocG5vicGN3CbaFgDQoPUJOs7qYqfWuk79dn1US4kyPdoyOvKe
BXl0EvL7EI1tOUxc0FSkNmuGSua5yVyecLWFJd5GbKSm3V6Gsa8piX/qKKxRPvlr+KxNgcbV5fLt
ppGibauozdCTwxM3JoYXEjTi7rdHjTATc98me9chY0jnPQmJMKL0nz604l6+Fw9Gw/rwHIS2U8ok
Ce4FhsT0L/6E1aEKVsr9lQa1wZsQ4+fMAUltjyTWMTv9g8aqCnq6TDjbwteOOEBOQmzExRahTBw1
v7K0XytfPdNl2Y69TQ6/52DemsgBiwL1QDuHLPl6vqOCo/kZQlGbfClUhUhaY9ywFqmrC48/Ky/g
9YlR+KM2rQGfwlSN3g0U1Ucrci5ZDVAIEXKSKNHixbXFPZz7D0aLqBYXyfzvKsBrAr6sE8jwhvVS
4wXYWHbOjcN7iYchAnNiJC07op1twV7l58ujiuGOGCjALAzoc7ntctzQBWBIiaJKCjDSgFiUh0oi
iUyYHSGnxmcxjIhP/7cbpHzivo5qkcuHjWIDZp+K37newG8Rgd4xXf1uIywHWHtbP6qtHOpvHaeg
c6AwH/FQ+t5UrEdc9SWCXqTMWd5aWEd0KNBKQMhPRwAUD1XPL6uX57+GOp5ewB+/GcZw+ThrRa15
cdy7W07Gc5FCFHw0BZi112MmfW82FC7P2kKM87V+IQFXhSUT5PDgoLswIj+eg8UVDjOrnI4Ce319
bkxWYNbAN69QJefNTwndbiI53dYUI6FnTf/WwX6/fP3M3HnYOMPYIEUSXsA3RLmRW1Sq83H/LfP8
y1XM4Cs3xXdOWxDsbR9FvM/PugmtQCc38kph8B/oCGFm6HvKU6Ft2r+iMRXg6MZN3x0f+MqRECLG
uQJWaT8Vk03NlWalrGqZl1Z2aYbevcBUIteMrZUzH/lSotvRgOJA3GEN30tMbg8qpN7luY6hsBxI
aPwzHUmUJ3qtQRPb672ujAsVUcjCV+hnnM5/3BbPfhGwIU7TYXnnSu/52YV21bIhqrTXlrH0MGUe
hXGDlXdQXCuDllsC65G/ry4IltmHfOMMiuP4a8QwJ19gblatiXjJk5GbtxNd3Zmh2e5wP0LMMFKx
JFxgrb1ycGM+/q1FNwE/T/1648NPycCs3fC80sJBCgSt8w2ubCFq6wwd904vw/EL11Z/T4TBgtE5
5KeVcno0Y4A9PIRZCqFqRQ2CWO1Sx0mrQIxtGu/uPzOgY3t7nL/6PQlCeCNdIiB7VMTbKEcM30fU
67QNawfOgH0JQMtSu3dtnThlUD147knkHLWmq9NAcv9bli38hflsxyraVrLaLNlSpGLyRldv6750
Lk4129/+PPmqk5cYhhfnmzYYxX49oXO9pFuT4VTsbPYrEq54QIsCLF6dYD1gxm17Px05IY5Gnj0K
BGLnYbmn+/B3CpWDDJszuw89NlXYZkrrLDzCv2tc+Qg/nZgBjyx8l3DbxAxFTSF+KiYwEfxBCwCS
9SWBfWcm4Eob5HMFixW5w1GIehqs1QKuMoVlWkSQ8bwHUu8Vnzl4JwADs8NJ3bK80uxc8Xw/Rxc8
tvnet2WBSzUwqWfEN+oaci65U9huWIJ/7ZzQO75vhzNnZyeYNEEx5qnqRoGYzVhmFSESD6fRug3A
3H1OyIahpoYS8Jb6TYxRcXJQhWsMO358JV7X2m+KYp098GEGzB7idRNk7WuVXkiwTEVpBFHYzNNf
SkEIoDkdvYS1CkUcoPxlV//IWYoVFPkk2Evt5xHjogv0mINUGIC6a1rqjFZWWybr2Ax7xEPyLUFH
Hel1h6zIchXwyC+yrLZqNnTUF2YuzVWzMyh3UELLLPQbeqJjBXTDFCNn775g08rHos3npyF496W7
znN/yxphMbnNA6YfeECRCudGGW9m1dsSDO/yv+W3l1HlHkifNpRFqcm3vRQjwnmQU5tU2kZgFXL+
9bhP5KuwIYYqAsqeI/y/DhwVFxeb8G6K1gVaAi/w2Dpzo7A8kQLVMHo9P0y+IU9lYEsk/lCafWW2
EO4rNE8Q1zdHgQ6cc5ACPGUvIooSda4TIG90ggM2xMpVi0yMoKna00zeL50UgSFbbXk1rD5LnEod
vZy/ekUlQcOT9Rkp043Xy8E2BVi8VIXAuCY8zJIgzge2ZCt1fan3nOZK2/sKVZKKFkGaDYQwzdvm
/wCxYh4/VLVikbnzlPrxuGqPIwtigU+m4a1Eup651Kiijc98b7REvGBM6PFf+u+T9/GQVodjjNvx
9W+XgZL7bFcL74Eh5UE5FK1l1nxnHiZ0CSAoprWI/jkWCJB4XBYLj/L6hXTBn0Nhg3Fi96EZ5DJg
ynPyyoW159lD9gaNZlzwEQglOVnPplPhYvUEo6HoGj0t8eV2Gjh5QVhtFs99jfOsVGuCp/KAsmNA
z0+YR4T1VcsnpfpiJA6JDaixSFetV27buhIZ46yv7eBbZTEilSlyZcTT284Cwu/BZSttfN02K9RK
PuBxpChgsK/m5lyE/p6dUM4GimSTAerrzE6tuI5mBBRKvo63C3QBi6KAWfIwY3MYOQarr5Cb3wCk
K/lYHMUbZlgdpATxtTANbfN1ZECxBMUAG4JDrthXVmVUk5ILKGrk29ie88aQOuNJ6sQEFBwnjxmA
Sjk/EyCy2p+NYKoK8YrVsTqkGohAAs1kIGAYN7KTPK1VQ/bdAQcME7y/idQQBMDTrPcLvRZxv6eR
be50NQl/Fb9fcWgaWO9mvHaUsPzpaWuUFHgtlm9iH5m3S2WLnXDRMYwl7Lwp/gsCUfHdDGZB8Wgg
UxkV3W4TaDm/wCyhA7AUAG0oTgP5TdWimmUE119qQ9/KKBUfqbErWn9YGHWlozGF5YpGzYEbrYVz
VejZirf4tui+gqv3T68W/8Iu9slg5HNL9mHaAXzLOfkATGiS4USiPuayk+i5R5YP2Xmmqdp6UDEg
ggTMMJkU2/pQExqSvSYFzvRI/14se8bWSLrG+oWNkDjFyJoYJu8QYR6D8MznnUgBTmrj3NfJg1IC
5rsA9XGSHmcHLGodeU3stwJjZa6lFDhxm4hNJEkNHQZK0Qk5LB4c1n3OUSNl/E9rdQjTk6bZv87p
volCbLF0MVgB2b6mZnFMH80FhesZTC5Vo+HNbrLdnTvtk5/13tR+rQkeFSdUsevjL2MfQXzd5P9D
Zxp/hEnCUCfcSs9GwSm2IVxRfFtd2NsSf4CdP1t8mWJqA9km+6T1OPtBThVOFqfVV5YAo0N0FDW7
a2NYcM4/Z8XL7zi+Ee+olqVJC9pn7ExLzz5VkVh/u63NFmA0yULRgxXRELzW9qC8GzuZ3XPdeadX
iNkxJUTHXPKyoywTaKMMHfv6INLck0hd7zc+7/ExmQFD2aPEC5/456NmsUukcx2QhxhgnA+8xJma
Z1Mw814ciaBZ8tvYVC8Pj9w1x41GnZfzmwfByBCuSbS8JDa/45r4gY9wGmB9Ta8Ra46Bq/b7jwBy
u4b5xt2kgRQ8k2JK3S6undDGlr2i8coHSNvmuSiv4LVMewrg50ps08e/AkAtYQIgla3/ucvGGgTr
BSrbSBGxCRhO0alqqgSUljbLU29wNRyKSdfRl5V8ms9joYvYuuaiNfiJECnUe7+GZBGUAMiVy5LS
TPZFhOI0mIKH4q/i0VYqIccWLVt/C7yoycejA6vFYU0w+QuLj6pNzIGdgRJb37GRSCrJopmLSmIR
6z7QGZEMC/3n17Hm5M7rs8C7pm656tmBvyXEn5N/R6R0DzpTyBgz0W6KuLbNl9YBZAy/9RDZSBGg
w/p/3ulvyE1FbxnJbuUWPNFYh7er282GyKXWxkato73EfF4x0VhafUGCo2kjPPUg1OOInAYXHKfO
DzvL9dOi/vq2rCE9Khw2uzJyDNJeoQNXyqJvA5o953p0QiDg5QhAcOZ8/bYoDjlY4NAwIzTscsEy
5DHwQ3a8DVGzHAASVVr4QRGpTHsesEJjB7CbjuB4+m9FWkJdn3svZYCoq96IDL48k0/ffQZQ571e
iB0tC91eD6oGcdFjK5dP8Isl/x5a6Uty0y30ZbqTp5L2FrD0KxL4S3LsmJDo7vV0ku+tfq1Ct4b+
bGHiQ+eAzz23QY9w4SGlqayC/nIndN20G/8n+axm9rv2/7FR4jyLtC9dNOGNQDEiJ44urBN6T522
ovrCk2jjzgiWX1AxaKtRhy2PE3v4nf7daJwNepvU654qO71WJaz0DZ6v9Rzs5iHVcvrKnzUO3iWZ
FvM5JmpuPZD4DypcHNDzVCH+xvUIo+AizMEnurKL/RHNcDBLnaD8eTbiW3SxWtt+hjg8WnMpI00Z
Z78/2/vUozHzYU82Vamox/dVDuAQMmTB2D4eUmUGkw2qw041NuP2v7PbomPtOHtsFJFwyCV/Stv/
vach6ulE9qPrNQyKy23yUNEsDaESfCcWTeI0xFFD/JQDM09lmdgZKtmXBm5y09WXSJaQnRrc7xC2
UBaAsQtiAJ75Ksw5SZG7KTDQbfR0LrBRnWgNuOTADhNXALFhXtW4XzHniaTXbshpdRwPtvcl683J
iOfWPrDDNspRuT4ETojWOjC/UeV8vhk3Q4KQbi0LwVwE7nAeCGlqdo3xM9z4gpBs2x6EfkQ1z8V3
8jGkbl1h3A6OCwF4iHXT3PNNMC3WC+Pn1gK4Ieo2z02/xJG3OL5Z9RBu3hEJ03ifmaPuOomd1H4M
z3TFksxkQ/9jUsXA0uYEmfoYCaHGhboBYY9/A/KvctRaLgHVlst8hydorz3IQh1o/LneHzEkmLnI
45z9173UD3OtNLPFllXHcxzB+7kWZez3y6sh4B7Ez57EFeWyDgd/TTt9QkXuHBaMMRqR6L7FmPqi
+zTY0e9DfKqcniHaDnLetvdh+JHBb/nkx/lITLfX/mm2dhsYNDCOLq8A8Jwr33d5MXbkP90B3NdV
50NyBk2hUyuICB+joUCa4D7pIojhlEx8AOCroHetruVxNkCLkFB0sUjxeyoNXdCTxQkW5GIYvICv
BWwCN+bjGzHN7oqq9cDW5PjQdFg3+wME+MdJ/s57hyliq/s4wm1eSCuy9JVvhx1Q+vF+WcbwDLV7
FbTXRfX14n5aOQH8WEhGcEnt+JFZnIUrlMnDo7baehkAu7KWu5TdFsZJT0eVyJ3nsxp8LvKlLCoC
eYxBPJuCEhMj1qbzwfrP3++eN3JETE/i+FEVGq880+OMhTRcPtYhUvHLdqxNJpv+uHSegz68jXZd
hYhXtlYHOccknSmV8b26BNQE91fsKQ7lOsVXOMVLmRP4UVOIaFYhUkO6LTP4KNNNntBMlzzlPkag
xScOsBSm97cUlMdGgkS7+uejgrT53dCMwWCSB0jlwBS20e6SURHVyjrR63TBmzA1H5NaJ+lTIiDa
vFfV5zmf2C6OjNdQv2PiQhYEQPvWXSXOtliqNVZe5r/ImqYP2T/4IZUasvWcGV9WbKkznZZbWHM9
J6z7lcAd+0JQh6EuPcFvuO31Q1uE/WnKl9mKi9n/de86YJQuq5yB/s2OJ8pe33GVi3g19MTTVKYn
HnmAFYYgIGqM1JmvYi2qdopMj81waYbMXoeBEwveVpY2jtbVcqUnezoTU56iaAw+jigefw8EqDlw
iO/l34Q1I0/TNS1UZrcXceRVJMacKy1DGx0lNJwKXTOtXooSii9AVTrzBaoTlXo+pYe+Ht56WUOO
bdMITbUGd/abknUH1YWauxa7FoZ7zW+eoCHbI/IyxTylVRJvbcnIhbN6RGYI/zwRgUzqj8Dw+J8P
+bzQLw1eG3HF9twj50rIVFBAE1k4Z4jSth7XssP7eN3YfQt16lDfmGIiCr587wFnnJd/JKlObafq
DTI29ovzflPBV+H3xjM/vTe34LH3msOn4KGOko8xt+UipJc/p0wZ+RtaZGyHHpV7ASt3xutdimkQ
az8uN9fZasLFHYf3CcJu8psGn4+QKV+YzcNzJ4J6ELERfgW+fkIxBfp7Upu1jrgK8JG00cs4Le9e
gNe7Q4K9z9M/pFERGeAq4iFntSBMunzcBHNf9569hDBbAVtsvdQlZlgsnw70vQhXdp8NWgx4E7Z4
MspPjjvqVADR8BIbtsJGHmEgXla45W/UKSRGccL3mt9NK0MK2KEjfKks96OVdvU1yFPQ6jM6hciV
vhkcR1+KOD+zHVNwZu/XVPF+9dXVZPdYVyHak1pu0peBADrk9Pbeap88yADsF3YzfI6AVR9L4EIP
aLFN697opwgKU/oguAHHYYqv6Mg9Brql/nyRX+o6e7K6Qjxu2nNPB5A0YPc8o4N8uc7nwP1uMR/v
lvJysoJVvvV6bF+LY1xf0ZieqEUXuugPz1IRC2xF14aORatJeGQmHSzb+2qHCauFxj/E0/Bffd6H
oybVXJGZ76ophmpnvMF+ahnRFvfOsmICc4wReKbLpipBei1d7IVfU3H2C+Vn2RMea3FQPSL++8iH
rHszhSXgEYzb76lNjXwe7WVi5KGY9QU6VH842mvtayt6CgW0tcxk+DGrz8QoYeUbldzyw1mQzvKa
Y3kYNSje004zDS0niWVL2MwuU7xBW7+R4eCoBc3auLCry7k1x/4FyqhG+QTZ0Cp59ojT26staziJ
uqKKpgzNxxAL7QlsJVMSDe+NBc7tgbTg4c9ULQdfoqQHxCir1+yxDFJ2LJjqxhrS85CBDslj0CFp
cLnMpb0DWJ/5Q55GWSltoSHmp1igHfFM8+kHH1vZavAa9zFLeET/xDFK6K+2wVElqjXPxb1mqtDa
bZSifrD0oJ7khkzTuYl48YYH60MLJJUL03IqGfVYLAvvGMor/mrymfVXB5WdV/NOOLM8Fn//CNhV
SphBsI+wnybmrvq60RsvVnkaSZ1Ccl52ELJ304eRGFvcUaJQ4cjk4rQ8egWQIRnLAQ0oNzOn6M+x
PDToTf3+7kCbnxmgB47xhyHbady8BNOYyTFk6kUmr22+zi+ttE+r24VT9/ebtean6+Dz1yeuHCxr
jzn3COacztJXU6jP9185KBKvJcrhtqG5/zIgzUuulbM3hIndHod+fdtLSnoyHI2ABr1Qym+4Am7j
r0ov5kR2qaTuDBGR1MPzQMt9TZkhC2x5C5I/CFRH/RxLTQ1s9SrNMXbsdnlDow5PoqJhF/lGzV3R
7bUWhY9nIDWqoOo0xgbVmI/cZNpHGGmCNHaZ0Ww/Ckfganbi7EZparFVaNKYtlfpi+xI4TWV7YaF
G1GEUBl6SAJhin6vD8YMDnd1rTt+6e6jYmDqQh9BXPPUW3hv0SdQCn0jxWRvDi8RrSU6Zce+v2dP
ZofBMdY4FO4i+XPrylP1XWrC8okAdSURL16pNhicHeNxngmtEfvACqEzYTxCge9CjW+epOnhO9us
y+tCXY6mCkoFf8YFt4ZI9l3EKnpHjpTgFQoFDvdJUwNa8AzUzgedyULqLwkWDWqv3bSVgN8xZoKU
rX8Cs+HaUfC4M4i0eiKA9vJzPWMt6A1v8xwxGo9VjmWBVLOY5Uf1aeIdwHsx1dDSMRvRCOzxMbpO
4vsAVumW08z6IB2N/r0nG1Y4fmjS/U6YKp1jNGL580x2IkwzfCFeUbIL979NcC9v/fltDuDx13c4
jlMC8MZnkTb0qQkEqVoKQeHRqh01sdjiJG7NVh4Cf4gsZxavvVmphM7eeBBT+WqRY31BigZ1MPHF
OXM0J6Mmn3gRsukwtj0/COt6UZt2pziOwtPCjMJ9GZ48lnWi/Yursrn2WlU2QJKH6XNVq7fCIELs
XHft5ZegrFYLzjVQPfajq3UvUTcNWWC9POykYbU6dEA/hUQ3lvxHLNlZ4sz1ERNRv46Zwxdkb8aM
kh863Ho3s9Epy3Czq0tM+w8GMPxYbg8wVNRziIy3stJIuoZCs9IxfdB+uMK8+IQfez4m2FtDHKOr
54Y4DgoL7J30Tau6MSBqe9u35iBoGFrv7nl9Sf7cssopILTi4aQykrjhhV4151ZEld18iLSxNWpm
7RDcwDF9RW1bt1m/zOT5tp2vjviGZ101p7sz7sZaLKPXufUlht82AUO0tIC0xXwcd9MZb+uKf3bO
zlcSSFLTraQxENfN/7M5WM4TD5Ix+dohQ0mn1cfwh94b6mpzn5rTA5Z2FE94+hKXhp6jM4xtHOIa
GtMkywNUVeRoD8zNbJPv6fUwzwCCGI3y/eloujN7Ll3GS8xVQA0EE3Jde/BqfvTeLjtCy+ONqa2j
E6TeHyo75TVFHdW4RPVNVropOPudYQcRQd2AFDWeY6b61GRSIZHkZ5i75NQDpSIeXq97iwuqUv6i
Of0JjVqdOF70JAKj0sRjPoncF2clmj+xNp/iLN03eiuBqzakrfr8Tb0YgfaVJgBGcOCpy2k4hJnb
KXwQD4r3u54K2yy5YZkqq8Vnuumtt30imFZmerrQcV8vbRHMYrotzqXXOrLldVugJJP1NsQ/5jZi
xzeSUbtrBkPVBBwz2UKsGSXHlQ93DoFJ0QIs8U6+AjG3loBQAiUoQpvMf7FNJtIyc1vBBBvGnRD1
FB1JQWLt/cOLHxia/YBhWa+C5BFk7qTnk+KlzkzC2sz/gG2d98EHh8OaMbgGhNTJWcSMqIitdbrs
tvARgmvzyKaBnf+cH7ru3vUMD8FB/IMrr0Zk9RupuHQsrt3jFoi/lUOreU9CWhHzR2j13GtA8fMp
yxVsBpi0hB4DuBOL+Da5WmONFMS2qAxU28a9pRWNe4Dw0/ZdC6m8NQ8Hy2idbDCELGOpx6DjHPZh
JMQFo+KPAOzMM/RB/D7amIZSQXemXGgb4PTdL0mKE9hpzG3KtnUDQbsqe4hbOyxUWl4wBeusvAFO
Dr0yk6ExIg/Q6x8jHMiUJ4BCWSyjyQJUJ5DLmf6h39b3w5Zb1yIO1IDmoI9eiouDRTz/sj0qny+1
QCMN1mnw7Ay0hrucyJaLPLTdpMxG6cGC8yBOKQHShTChHQdgxHaFenle3KfaQqXfIEk/uu3UvDMZ
b5NeLZsrqEKu2oXHIpRn0b3jTvSvn1RYoqGsxWDC2zoXIU3JRmcsfG2oVoFWVTXPBz/L4DvbzBQx
xQIvoYexi2rJPYuJkdx9jOPoIO3YzLe+uBo+otVwPxq3CTRkNvXZp4g5pslio1yb0iTQAMQti7GJ
homxmmDfp+QKXLWRJwyK/8cIoo956Qaoj3PKuX9m1sxxNASolmObNN3+m/udtMmGnslZPeAtMmgH
JweCEVQQZ3N7nEMhW0ofr7N0yJOMoXr7lZLLbleZtEmRlrEh1XwQ/IDe3ztA7536YQEGtuXH7Fny
1cOwtq6C0UHMRBkhTyhEjqSbrCXhx6KruxJKxqqACyk4t6piUb39nsZErYQWPDXqWOJ+5CSa5+hm
e+wqpEVYzn5NfnmFEPhu72hxIKu/LJ7SoZg8k+kdIP7dDngImebWCUtw+EcGxjRJMjPAflAV4fLp
0dtrHat0qoTm6bgTbBMZyjz4P2hZE0QrN2lY1l6JcjwCWjcle0itxziT417hYZH+wbyiNP6AdfJj
46U6ED/WaLp/8pqT1cm4LZaK7SEdmE/UmlUtWVWH3pvuWGMb1Te630A20szTb7sWEIaNIa1y6BjY
MDxApRofMJ5Mpr8uzQcl5spUdLEYeGX7nDQTsPf+Of+pJ1PPP2LtaUiTMC+YMUUR8vuN2YCFseOo
VcHSoj3BQvAQPaJBNVbH/Fxp8J4dHycmclImgb9Xoc222KGd9BgS9q9PCqwPvMfnji5RM1AvqTwC
T7FWHppLeHhKwOuTPZCyGbT6ajyOxe9E9vKxpiq3cDrpRcutXw2ezYMIcJakjF1MLNPf3DV3ohvP
Dc3gwWVRE8PJOeSnhXpD4eFNB0ycsfUTCYzab5Nem6NpGtM5LN4vShlmLUGPFa0Ge1gbTZH80A9r
KopBRqn4EH7Et9c/8zbRh57q9fEGBjKLm6uj43bCEQiWfqZcCPCG0hFmOkXiD/nniSAyLum7jb/7
rp8eBn1wqmvMUSUs2GtPapEh5Duj09OoOjcny18AHoAbO7rfHVn9Jw0hzg1l0D31QPw9nElQWzi3
7FOH7TAEJN7i1uipUJdFwq8uQjUY5mXtxdi24rnumRzDCmveIcwt/PNp6Ev/SW+1qmsEppIVzVEr
VPEQGA2bjleP7OFI96qfe1mwaMiEOuHW1ncB5jFRIGbpcpoHnuPpJC2pg/uavJZfhs0owUBtz47h
/J9EP8B/AD7AQ+GANwHHg1ocjIV5TM+KClxcb7D0CUO1IfqWmpOSNm77DhNhHpgAjjge13J/m+NA
PYQJQ9W1XUGfJMFQW0R708IQft+nlof2LH5eM2je6qp14s1p5AeF0ALau8adkyvPziicdYp9Zh7E
iO8Jnijb3O63qqGgiwTJVPO1RwTfc7WslahHxTFvW91uYIE2BH+3dN7CWGSz7+9/kfkUwnPro0Yn
3RPxc6MwCcqNcoX7vNXKSODppooszJqWsB3CJykZPRU06owjYGyo3YfqTa0pdJ0Vpgyufox9XB8+
YH9bUNNg3fxdk07EbETbuFcvl2DzaRG+dXiOFNlqbjgLwqeArN25sc1RQEUnMCK975PaNmiMaG4s
1JgJvo5YvtHEhwjJky1UBIJ9s3Ir10hu+0IkpKemzf4p6M7bdHTX9ecm8sGJC0rL3zaJ9JDO50Qi
FN5lxyQMFEl6s0X/Nkbv9dLqniamEl6CArd4spML62GvT97XpweNl/t38WDp47IPRt4r2sE9IohO
H5bLYI6kTkZ4JzyDAWuipaeP6skE2PUOG6knZOzzIAMapaDzMT1ZYb7SDjlBqBkbiiVXqNjMKD9o
tehViDMgKA1Xkq2qtggts+JQ7HVawjLeskRonBzYt2lrF549rZLMaVtbxMSGKf66obVXFwndzQK7
UPJYW5RPpSgeYC8BhS8+kxB9WlC1Zms3LrYbM7M5HvHqx2DwoM4dAOD8YC//SG7kq+SNQ2Uur7Pl
nvKBfsDZORbhVdFMDOQaqEMga/J9XHINFUrdZ8fXURgjn2jNLQW8kC2kU7TYju2OPL7hyxDG27HU
3EREHw5tdYoOo47WixGWdV6tta1lUzeCS72MLXYylEZ62Yqxr1Zzont82a11Rk457bSAT6oSqANU
a8oiBMxhZLFEvI/f+sfuy3lwNkf6cZZrw9E8lfToRhlpBzuM1m+I/eAerAXV+xmsMCoP+NwaOFu1
3ocqqjX3UnWxjXE5cY2iAnq1LFe+MvDlb4zeYKveHNbMhvJjJdWkJYlQAkZ/ApDLUMf5UyY1ru3I
y4M3DgNb8cKh264GPmhGOfYZXBTxkkUukiZac+qcHysCS1Fqzz9onr/MJweRmkgyXZ3jH4LsPm+Y
mbMlTqb+h1fYL6gzSKz0cGHkwNdgPR7pI7W/mtD6lsO98FBioGSu2PbSu8B0ykPxAI4bpTkf5pgB
/Qk/DSR+rNgM5iEx3/xCpb6WrnGzMAmU2428Fa7pcm7lKblHibcbMLEzEQav7Sivm/67hKr7KXex
ktn1nKEQdsbw07aUbmQW829ER6cwNxhrE/D8cAcljLouwjbS6YhDt3zk8FjIMICd/CFkWz0zM88J
EWdIio5U+vEG2wTG2GoJGSQlSlcpTpR1uP0dYjkB6+LpZJtZBUzP9HzFq/KYcnxvBzPJ9zCsCcQA
3oAhqr3GqAS9pzNzVVoEALOAG0IJxwctD2LvgGJejMiBuxSZec64JQgq2KsljazwLMME85Z4ierz
qwN41xrt+SorkjbytIWoFhvqX9BWvo5NeVFnvecrneS8Rr3f7P9Hd+xETznpRKpDam7L/fKeX7D9
JoV0MCBS+2uazgJiuf3k+ZBU6a5eeo7fPV1vzlMWm1D1hmgsLHvnIG1jh365+SLl0G05p0F12iYs
dcRzKXHm644PsAfhDdnFfSJI0ZUzxckyWyalU1Jh1oohxGDI/rkLLxWr3/y18MhEKrRlKzUfvEeu
yJSHh/VUhpbN6Rp4NnVKlhKVFxr1016FzWPgdB1RUVYtZQ2GBsb0ihFoSrEKvYnzArZlLjVVc8su
9TadQeWF8K/9xUzrafgx/iWmy44bZnqTBSyhZyeAUoVdPJaFqR+5gQpAHHweIaApunZIFKemppWn
aMHQQoU0JnLoPASepdUztliDL/elfdWkmY8QQj06DY1Rkz4YsUAEnMFwHj3IzXePv+ChFRnYk0NT
MTmGdDcFWcIYgb3eaJnvWbCYHWi+b9GXMwIoeCUlWD7gJNfXBydEagAKxTD8DIuVAbzWsekl1t0u
PC1ULgeWPdAOksOmSNJnm4p2u6oMPhUS01TrYDP45m1Olg8ynCsMORsEgO75uowjYI5aekCiNcZC
MSMre9wOZTkwhzMMnVkOhuyYWyjOA5Kf+IomK7gK7EgLukOzeGU+pp7qj5BgUtLGE6lwDmWUtSNw
CI+whp5RdpysZd/Gx7BR4d8qfYMjgOIGtnkms5Gd2KRW0Ly0V03NE0ddAwc9R8pmLQracbMe6w8l
B5R1puCD5pDP8v5l6GjRz3cTwzCZH3WNnBOdhdwv0NVWzLqWmg37ColFJXGhPe/LAlWIkpt82BcY
Hvv0XU8clzuKGAJweJnTU1gKj/tC6PEKzM8EvE3yzTa7ppIivGXVhmt7OgUl6PcX4jjY4ynd0o/t
O0zFb7sC6CKxbHBXJ/i5hw2pE3nrpsvcFX1tF5vDqXPm1tERLYnGptGMGvTowtduKpPww0SynZrP
gbixdpDDtgXUnioLYwsBL/0k/UsfEHYgbjIGQRXoQyxZ4O+LYj03TIWnn8khVL3CQ8LcBn8ckfXo
DSRmDu8fuczITsE47+KHZFbeNaC4DO0SxZyNmgV29j0UH67YVBpOYnUUq+tVJNZJctNkOVyFhoIC
+3lQID2cJFhr2YYXF5O2N3AaAums4lO9H8h6dgLIv1+SORaGsRP185jJSJxuA75y8V28Cv0Xo/db
WXfAiYBRd+rUupm5LzU/ui5ABTJ5sucqrq690e8IRrWq2BB1geAlGS1w08J4HPhkHiDENvz4AHb/
XfHtBiqEZn0Um8w8h/bXE7zSsbd9hx1k3zrRvu47cWloD+b+8MKDexNeDTrMeb18sjSDuZY0cxht
cH1oyUzrZgCZuEYu6yZRxytOotGUchuSzC/5VhN34LT5uNwhxXBZcjo8So+K+0KjEgsH4tvt/AFi
wre3OfIOairqBOEqW4QXfU+w1vHg/0CgcER2wseR4XBxP4yPd/BEQS3YNk79OhowFE3GQvOT6y7i
2HTQUmjVTfR5j9vcVTiLDAVFLN9V3PCbupLTqMx8J1p/47rC5Nia4mndaUEf69KSSm2lLcUch+kw
nm98TaTkCeuY8apzvQlsZf87y2kyyi4T4lR++Lwf4wmisIIttUfYmWg0qa3TnvL/qo7Qljpywc1O
xWgfV5M8ngW9rcQPlQQdpZxzgCLmonvt49tAYQexh84MIqeX3W38jsmXdEIhav0sAcYyFSs5tckp
dUePEhKgHimqZfvZ3PSSBRgrn2vMonjlJMWKGWQAOoLxeQ9wQqsqUpChsw2gmyDFXUZeAA5xu4L5
3YhDgtkTE09um5uwfpw77kOpz+Nv5eJkImD2ZoeK9ZfvMr43B0W/Gs+VThwwFQkNxPvPWR3OLjU4
rl3C5pVifPByz293Jw6oPfJThanckdDT0C05N4QB1bdb4bwOXWqYPSRqrMbBheMzGTBcSNpxOLTQ
eOSn6S0qmn4vWSUzpzWXvh2PZhXjLEW+OBsqxujXdselsQBxF2N33IWexUUNPU8vf6H4OIblDw00
mk2hA1OqNRDG8XADZmx7oOMRfKUAMM7xmnEUZpCX/qLONhUjmbGbMd9h0aIVqGgj40wcRzE3iWNS
BZegKZgfANwYb21eXLCRqzqyYcQH5/NFzH3+PJJd72DsvsbDZ0KhMoRDrKfhFFc0MnNVLZSpAqoF
ziMy8tL1sl6gZq/Y/wtJFA9OKpKXTmngNo0Ar0dBeSYvhoI2SnCZ3T4KLGNY6/AUh4EfOt68jshW
sutVw6kDsJPnhxAjNWWzCJ6w2WyxZgQ0zh3Pb8EGngT1WH0lJoFokeXCqgLrHO3abY13g1y6nets
/1Dgyn8+DeakwyhdxSZgmCnQpuHfF654aBeRQpKeSnUZvisg93rDg578p/q9jsyVxD6r76S9Wa2B
Ccnz6c7AGwJ4Rk7GCQpZ+qwL+0nKq3q0CdNXxGedphmRD7328cYZtKX6Lmg2mHtkKWZtvfxRuqYR
yVv24aSeX88F4+v3x6ADwSIOMYNSN9Yh3M2Ikw344GNZcWW+GSYKgoQxq+OOq/5biIS2ROjEGjH7
g6iQW9p+q86tljTqIFAyHvj1xRr67OMLedV09adRXujMJSehiHyBXRG5tA6YkS7kLc4lltLSWIlJ
vXReKrpmKFnWa0TEqmD+0X+XUmOyOvkyGnpBTVCx0II6/Z6DbEieOiViWgsE82gI5/4auD5EkrEk
DeeLHIg6kYDJLZq6b+bkkrMQCrsXQokdG1lmX6OOZxk63dHwZIAzKCDONlfwq6QDtPSsNZABygBP
dLjdlCvcBQyAiOb49bJ44iX1O+v65eOT9Ijs0ElK985C+UAOyltcCnvdw1ehNetfP5QsHeQJF3fV
8vCniyAg06na7o/gkNVRNiDoVCBObT7mnIvS6yrVJhmk0pNFvCZsCuJ2lPhHhTP4Z4sVeASUjt74
bRQfCYZxIhkvxwyDeze8Ni5io2HBUGFKhbhV9GZ//J8eyy5jR1hYNXGDtul044XMzcIRkYSbCMLw
d8E72kzvK0IqTOeh8wKGGG8OAE/Cvno8YO0qcGWJWIXXYhMYCtH4XzgeZ+diMQem8nkTIvdeNHTK
LbZSa7N2kjADCg6x7INKWeYCvP3dPJZ4YCiUwUG/aOfnZAHwOaMXuzmq8YIGz1TxI9XIiwfLNTEi
PtO2QP+4ht6R52ArHeA36C3LcvDL/e3YAfai7car6pYFsk10650bRjxq+mZUXdMprM2GsFm1n9Uz
kiidaXwYMEs6PWFS9wfj/m9Kauo59uTCRVhIrUT2v/U9K5c2+K6lDNbiTgICJmj4/iZJ6vX00iHy
smGb2nuIfFCqAjZWP10ScB8QHsBK1RNaYtC+wLc3Cl8ZYxP0l5V99ZOBa+T4qxy8nOAujmxi8IgM
usrrGWPtdEQYEcj6bWHIrp2x18s2ZBgbTVEUD7Vv8kh8/Ose7elihwtQ39yOTnSc3GAqhl2NyjUF
BmlZiMSH1Xw5Cop7SKW2/0Y2A2jY0zRhNRj72ssJ8mabcKRkz4rTaHMerg6OQES8eYjALRdBAQp+
PJ8gp0ramGogvKPrJ8377rlBSJOL0xpEGZOIDeiUMtrn3+Y39+jQti0dMoFsHZQMJohaCsK4/Nhx
f8X4cL6drCh+NiAb6l4S2rYtymEGsJwKggSU3xNke+ZqWw8fRWVqDwNUxKFHy7rqU2ytKyntmD5+
v+l6iTfj8wJIhu9RMfSh3uXVRJYA+O0Pn0zxXE2k3FuovFPpS59XH/w2Nxq38baBQ4iara6pmyYs
KKUZj7sO9MLiLPGZXCrv2MlZ8GGDF3wcnOREHVN2AKCWHBAQhijL+EtHJZFSJvysAdAFtjfo16oL
wU8GJ485jB0O8pUV/VgPOkxNwzKDTp2D0oPTfI4RYIeaMykImeS9iQ4AsRHPidaFK4x9Yr+w1Z6j
kpoqrobHERUHW+5TC2yKXvYc2tuyQgEfWwdVxerKHi/LvnAdL49q1b5KmnyF6ijlFsmiQX3gstPq
Fc9V8kek6LxtxwSMiqypXHJOYbe4iZ1bwUnCZ91DjGUc25TdglPZx/E8RKN4rDHiE31JWsdL+cqO
uSONrnG/UIj4t4vd9rxP/cJUJHPmndSL4Jdmra0KFI1JUupfzAQ2MFzhEuf7QV/IvaeyCnOTtpLK
JIB8UicxJCqldhGLaT8PjnNqByz/7LnULAkGqzceMNqcjEiHMHd2OszrkSTA7Uausr72Iorlp/DL
T4ivSOxIS/XaiyALH96zyy2L2ODXMCqT+jNgItGPQyScW6vpz9R+B//9IodJHuowrCVJvszlr3bB
aAwbtvNM6vfCx91gGXedScrkkbjR4ktywX6ZTjG2gA8XUqPQX/p5RGJnTDCZbylSArDQYWg1V8tb
dCD07dlTZ4DTLa5wFexlLlSW7RPtkXrNyMQHE9aA4pfIVjjEj0DZ+JOFCQtoJlo4rIBWCZunpt0H
JoWHlr6kubCKOuGwVKYgFf3hMJ8D2IiQcfj8cGXH/ZcdZfwAjQizEBWbT4jJQfqrYArEiej7F/r5
EFc7Cl/NrIwUiiIiXaBFdsLiUZ/1gDEQLPUUZ0TN8vUzQFeEbkcZz8TcOQQ4SUyW6Uy5Vuq4U/0p
7dElQnVPdn2jn8Zx5MFE7442VAHVQ2aVcw52+boATJ2ulitHQ9lNxH+MDm3DzX/MFpyGszUCbcLR
EUNJG3GZUeEdoDpwF9VjmNLMUWwjMTq5YuVhIrO+d124cuJZqRruEBZoHesuEfv+fKja8zZB5vE5
cZrldH1NTtMm1UVw7UqdaFwkfTUSHPv58G3rZVYYtnf2EkaHQ+Cg1K9KoASJwtaDxJm5t4vqftD5
vTbjBkZoRniBr84P0FQD7IItFHXfW0CKzfJHuj6VzC4zlyY9fr0jl3/t6FYD8O7rcKgf/5J0zglO
b7ZY//whCiBGCC4lIFTm9sPs792v5/FPsme5P5qkUJM9Mq55LGG3uQQKlgTs7vtI++kaYNQmZ21y
805XZ11t1YAADKxO0OtGx+F9vkX8o09Iq8FcCLmST8Ano1S8DcBRopoHQhjoqN7QnzTVayzcTDd2
wzIUYSMEyoL+lFidXbDHJ72NrcFbY/0iTCGWRTQGBChf1LB4D+yDStMRmoK3dvJGMYD9awN7L7gf
ndeuis609TPyKAhkHs9/2vQBOfWhJfDc347UZMsVVhHI1EaSX7eg7clCCHvLoazK/2mMDEKVX+ni
cl5KLzs1tsunhI4tXGvKYeL3y0mNvCvBmPHmjxN98yaTGKEoE8xPjHzEjK1tfkMuirUpVQx/jZa/
dCp4jBWiHGWGsV5WHAHP/8kFs0Ey/Z1lGcg6TOMPMqFw053h9AvoMdWZFl8UO1IhG6FAD2CHV2Bb
skhpbga3L0zhszMDhuORtdBcVs/E1ii8OBIvLMsObxOdJM7wKOw5H6muOhlx7LzR7hyBM8zYV4/T
W9mauith1JtLG644t2Sf+nHCNZM6UznwLgoKQFSPwOMztcljXd4otCIcQgQxKggV1cfAyDx9dpdf
YKIVdJl4Z1bFIknztu5U6XpMs0zIG7MpDMOAllTOuY7bu22lo8NNsGHtn6Cty/t6a7+boMgBH2p8
IaBOG1jxeqnoi9h0vBsqkpoV2TBwUzeYyFfGl6PBM0pkmRtTwaNdh9hIRjb7fOA/7PWcUUVuI5oI
7lbUnKz62fqiMzhaRqqTWsSrbwMIyO11dwc+B4pMwJJfIKVnEEShaQpObKwjnlMsYFTvx2ZZm8Cw
XUqNLboSXiSLHYHHTOLPDZqrD2w17Nhdn82CsxpcNA/N3lUwg+HNZUH0OL/fedD2a/k3TB2nJ4wA
A4i46upzOkQMMswFTVPPJIP4bFnsHLWI26tfmeBbXIvrjNLvEVymEejq39Wf6SD/bpstfTxg19i+
2s3YWMQw9TnlyAeLDOTVwHIeUEdsbixnlQlBoGsT7at1JpssNrSrek5rB8MfJUzF6a18p/IwaiXf
vcgZH4gKZSw8IBs1Ig3weQSrCSqbZSVyHoyxlk892aFMRGB9dBtpzNIf6l8tdrkzihMi0Xg0AvX0
GFRCdUu5GTSMs4bvlMQAqeWGFWKDUHsFRU3VSVRIvMcRcNmb0cfNzn6zuR4IPMZvHv7G4Cs9Mvee
GeGJJ+Aa1Zm1H+p0Cam/3mwrZa5ozX4wqToI17sPdw7Ci3GgSIvsyprSBN2ZCZTPanEfXUsE6fvB
OnxnfSgm0DY+rqLLHlJFQhA36965G+61Zlxo2eu09Dtf+QGI1UohikQIX/ewWgZ7zJ8mF/Dbcltz
N+ZnIdRZrOzcBxjoIF81llvg1LiWAnNRSgqeEJB0p3CAX2OL4hATI2LTfKklyEfys3syMZ02CPLZ
RQ9+m5CwaMc6rZo6kpKhMZ7izcIiwK8QKU9shMYjub2wOew3bDXkQ6H3aM8w+9XnG4XCJ7JnUPsy
lExBTTBG704679f7UKNYZ4EacCOZnXxaAIK4PHwrBeVj7IeasJpuSzmPCEvTdr/MqRN3Kik01FuZ
Cggf/ocmYiFrk38L/t54br9jqjJKXyrWmROzfMGov9LhTCyGy6OZKUpxpFpDQKLYDvC8rLropG3a
FPZE0L3kciHqxL6SefV2337ac1Wao/RQcgb802jO1REtszlK/SogN7vtaDJA8fpknxGfiYpHmt1P
e3PzuDdqFLKKC9jLQy549wpeEoUYRRte00ZoYq/mKKCoN+3JGRYCll5qjcyRtzqTI+uO7tMSkDZx
fOwBddkf+RCJqP+oNhn6U8JTKfjiGXQeB9bPA9HjB9NT3e3PAtGQ5/hhkw0uGdv4n+mCLWV9Hl7I
UNoBDK1JkHwJAA4U9BufZnwDqkuRw3Js0Uoj9t0VbMmfpKOVTVpusBTqD6jR5IHPwEIP9QVuHg9Q
8OJoM+Xdozx1YHG88vtIncu8F/t1s/ledgdFXuf3a2HPsYlSgViPuuXgOFr5eSslG28H1Msr6j2a
vIz+sazMCwW5rhOAXcPtVdv9VgpGXJlCLk0A0PyB/VnzudR7I/ZOHigPGsEaOCxaSX8612WpxhII
3AaLYg5rYmh4RLKZxi4CdsTa6oc7PqzVDg7bhUeQ9Xe+bFaYknEpAPd5CmmN/TzzwdIvwRdqbmHG
tRTUeyjgYRSECHcny47c3D5kb3QWk4LTMrvJBobMaOnjAY3ZFx+HusqnuBUqMSRAd1l9dOif+wL1
nERMgPszvan6MqcnhgA6IUm4WLx2urR5on+ycf4vGuePVbUje78m1myz54OD5rbLhra7XIE6+3BI
Tgh61uj/ExFaqhiWaFBBiZIH9nDPVjwco/NEV6Wo9cLy1kdDpRQcCp21Dn6mv8K1rkZgUTyl1NKF
WyhnL8tuigrj4lsuYIr3jv4poxJfI0BBFcpFz6ZCH6sOFusmzMgiKMmlqgxfLqpHsSVp146/xJ3Q
VnDff9xKZnoduj7z4TpiuRa28PG56IkswvA0AsQBBYU5BPAQkdSpcRvT7doNyitfPpbKUp/j0HKC
tHd26jPxbFbly/SZAuxtJpwvsU/rMmPxncw+3TrEgKhQ+O2JpTxf4NftrqZJeY0OP+TaoRSLJSra
YAdaiPUaTyjsal9y8HwXw1kEOJH9rVF1AqWzLMvK9ecYi7onRQM1QCakBNKRpTshisUg0e5f38uu
oJy8lk4b0LMwiMF2bSaPQNyz42nBFWb4+nuI84tLCDmoTk4oOUyw7fSYEti1EA3MTW8QwHTeUp2y
qchbVk8rEc54QxNBsmw/DGeLZoHytb33WC8x4tWhcl2e2fw1fIFTm45LCamowh4IBW0WMTSJTnyk
8BPWc0FxkqGQDNPnDruBvipFTMhEr/hbX8tk8AqT3sXdvjXscJPauLX0KBPMzux/t94Ob0xMqAow
yDfQd9oQzyOGmcy1iB2uE8Oj2iPxKhrlLXQ8UVAXptR2urgqfG7sxzWhV0vgZ4Veh+r5QC56BqC9
he1lr2v/LMhH/X/JeDAUjmgerBxNx5x+0uwpSLNpDVCFmYiziuym679v+4jjvTITgVdzJegx/doK
RscOXiPDX1eBUnYBVesh0cihrWSunjySMFvEPCFI39Mx/3pUPiYG17Q3R9k8oQQjBAzWAYIDsokN
QAIVXZbrRwSC3oDqVLdWJ3h4fxltT35DHCA+4vP+BXtlcTiaIM4rTuZbeWeSYuJ6BXSsw5L01/zp
oqVzsk8UlWq0G5bG7+c/WB/ynfbFumgsfMj4875z8JroYhZRpfyvqpcNfpWtk532gdVPmSepCte2
F0/d4PCGTXJD66z0q+056Ctd9s73nIoXhczJvjndSQUpgawZP0YVUwrYRKvlV0h1R8fa0EZUZ3G4
aScLm/ZXjAkkQuw8JxZGPPpbPThY0cIrswdtnvHPyOewftj260+9KhGujUcXW0F3twTYxyaCrRpZ
VnjVoF3bOX7upogKAqIKSLpnx4NraqgKXHkuQganeAYQoyysLNl3/RbULCTmZRrXOFzelS6daopv
8KIArBvQ9PWyjmlGUJs4oBq39tgIdgFuWNP6IoH/DSb2x7W0AJSzPXpUQafLGC1J4KO7Qm+0PI4C
X2NNFnrGp7KkHa+A887mxlqbIXMyCAItTFcuATqAGvI0R5CqRu5kT7yTDoRh2pHj1A34oAH0p4UL
AIbI6w9CSq4egpOKdeLQuLVAjmT5Of2BOYEnXoWqw4aJitrayJiLsbSeNSCsSe4k4gnQFIqWMv5h
+SnE6K0dsDqf7NQv9VDuJdzM9yubHrHbuLh1JqsIyOPjQjUQ6yw/BIY1xIG5wwqDXfND/J8JUUwj
fgproJ6n1EwXZM98ArBZBmf1XXvWFMeyuRXJJGBgMJRgEhkxIikuicp1KVo0nUFHR9n7rXFRsURw
ocxYheMGNV8qoK1sdW7XqLqjC74jXkJ6k6KIYOLtAkf3iRGHXuUU4kbDIcoAhl4QSb1P8rYhH5Ez
54DZJXkfRGJeb0nfrxQ7RawlZAaKyoLqXxKVmhMM/x/QYp3H2foEJ5uJix/ZbOwLtkSbp53scGXj
a1j+B5ttOYFG2O0DW2xMbzTORpWD8R6a2N6jGWPpiX97OamUJYMVj6aTHuIhDCdq1xCSgBJ38eVB
kc4+c0DFp1WoQ4H9YdwtaxnvZWT8gm5r+up+QysH8neWoVWOWCowzAvfQ+vBfDg3Vq7IQ+dTxLGK
TvPUNv47PYZVH85Y2k5YJsTe74gCUqjFH/usgZqDpIIdu0cOkTibSdDRYGO9no3nygPZ+3RcDcJf
DsZwz8ukbRiIDSlYmEeykpyABCT6s4gia96WbXlv2eEvH3eQhnGUW6wFlk4CM5R1QtzsfJC6wVl+
US1GjYn2WWd1H3gZa4f9q0ig9ROhILMMbskWTgEjFAj6dWxIPIBjarhiwfi4xO5rVeivYEEp+W9P
o2cacIPSHdIa1P1C4X+ejbfJQZHAOx2iLdfuzJD24QujZeHuWqrDZzR7zigJnp8e2KH00R8+7wOD
JZcBYjOeOl1AEKbrKgrRXgj41Dd/VQhgix6FgphIZKQmGphDujhJc7qKZ3KjD8Uz91bTBho+l9Ze
zeUA3DAO0j+hU6HAsFgqT6O31M518KZv4GXUlpNf2o0VywfmSLRSiLm/x4BT1bt5/cWqxtP1BKjT
UbVqSRPsGGBqQPaR8+cXmUebK3Xqpgd/7u4iDsX1Mxw/LIudX6yCNu+qAxpr/UdY0bikK0KIW2Wa
ebQ/FY/6MfcxZOyrgh7wZ3STKabDknZ4SKxnBssbznDvSuKWiKNMNUeKmpP9GgMg5Ob2LNzDUg+J
4Kwl/4pEa1CXN67ZB1nWpZCwmHLk69c7pIpPW4fGpI5Dbw6QOAHffd3yW26erAVTQKDpXMl+Cd2Q
rQem4Ghtwc7Wt5BEq81+/XssFyj5TrnWluJZddP/5cGKRojGbiA49QryA+nIjAYldVGoST9+yCJT
2D2SJwMWzCSCZXD4z8RME1kJGYAaCI60KHs/vJ0QcTFB4MIlWONUaQTgv7v3lZICIn6gY+qwET1j
hq5Rv00dMTO3KUdeGcuXr1hjPrpEP3elpdh80x/4zPgSVuZk5hM8JlDsLSR72cRiY0JRdEDjjv1W
yT4lJbu8BT1NiS1wlYH+p/un6NbO/XLBJ/QktYhx7HjR9NL/ON4uzexxY+xQdUuopIAWPg4v1n4P
vxrat8NERAD0wU9wUOlpXlfLL6D9AA6rUCnvWdsjR919mPRWRqo4iKhGhNEzbee6Zx3A1FZVQ5Eh
oW3AhjZ8YdZj5qXyuoIvJPXePOKTZvP+5uftMP+utOoldC9vyE2j69xV+aF5j5KC91Gbs27SX9Jj
yC04kK9tKyCNzmPaXr0yEVlJidjl9iAvYAgIJL+J7syCuA0v4XR1u/bcNIqSTlqhMIuCK9MIlKDd
rKLAOwDawRIUme628i1pHA4Q9Lu/LZ1pxiZqi4sanagqBj3687DIMhTizpmMfYuy+546WPVQ/m++
dXEw7SiDJncD86o7C2TnzmT9EiW5OUAEixuZRIYKYJSgIZ3pibNYqFpIMuIv2RP/BbCLLVdIhL+S
kzKR4MAzaSIbczuqv7x7tUztAy71iZ3PaOrOSzVui0kGzTR1LzWuMw8RTFwfGMNkxWZn/0W7h5nd
gO2OKTsogZtgu9nsgAa+WeZLsh4/QsMNwuiDeUQkwMuuOqf8NQ/dDlAx0oUBavRh8DvuWVIOUKOK
OQK2ePCfjCAIrEu+YfnpcvIBuQShF7Oysiimci9MflQTJ82Sss3W2YLG2NpQPQ+MnnSNgVjVLaHK
NfHOFP56U7eSseWJP/AJZdNefYEf/yWlC1IRG9lWDFchvyS4lJeYjD5w9yzXUOxX7+vydJCELIVA
WI44R+9Pm1KtVfKlyCil4SFZQcTqRqoZlVDP1ldMNXxRNPMyzfeKh+aR/PxMAxpSVIKk4APPpi36
Ze+NP4kuk7WGiplz7RQCQT1IUrBh4sGK76VCwKE/KAd7GG9v1ZDB+SiinH6ruOa3n9cRWHhWWLpQ
gI3OQ0UbOI7dzTL5az7VsjJwWdCKfhikSZoKqXWpJn+tCbMqHRsrxNQa0daSWw3R0sHUdkUvMgmy
M0TSkgZxy0uz964NTTm1hy5V/p83BOGHRJa5fWN0jdO8rKUpOsNKpCO05lOwMndhq6q6mSLQrpzM
KmBM45IvD8yVEPCXM5KkAjTF0TGI1tY5FtD5TPzFpIwbKaAgvhfFrCh7GgD0BhjXejtBynKo+YuE
vfPa28D23NghI3OxPR9m+D9W9mGYBpovyfgrQpWiJZPOkB7IMthG45iIx2Dvz36DQz/cCq8PG+Qq
wqP0gpf8pHySuHVzNNk6U1AmneDlYWi8V/TrQk7zlcwMPrYPZd4HsW029DPR8IJ7xUaq+fdF4Y1w
tCbr9pfzSW6Z3JsBdYp0sU8GA8O3f4MO0a8+ePai8ISYBZwlpdveOD4xKf7jJhAIopfmJrMYa1E5
FsysuZmYr/L+tQF0PRNFT4CyyHJti9iBUGGO1G5p4xoqG1qWfNf9eTWzibeSW9IAWGYh3QRSwCCD
uJbTBu+omAQqnIhG+vWKnIU+NgVjsvyhzzDsUk7YkU01i971/kxihzXy9DfVb+yvydcOcyEPFm/e
EfmgWw6SYAZGAhRuHuv82BlFmIx9iUS/GLioLTnQuxnB4eFbN37sPzMoRLH7GgkfVZQVyduk+4Xs
skbeVUe76aMEQZqljzlcvDhsiku6Hm1DmLjzan/bq8JUYeiy8TSM7XE/yBiUv/tt1utnIqFaJRHh
+w0Bkz9ua/lj2ZBoHbWlzHeTPmi/yecXPngsKbTleBE+4puRgvIm5u1hwDFmzGkczP+ZfS1T0TGJ
NP/wOQ3MjRYDdNtKlYvf6lBNVK/Mwo3Cyy+6kzM+so3hSbO5sy4d+VAR128iTzFFK/4ZughO46+D
2d9gIzYHa9E6aOfj6Ns23dWKmMLZWaa1pqPxoP3nhOFU3qSnCwpqVbi5leHR/VQiqTcS1b5exhcA
3Zp7dCWUxQyWOV7op/o34DHiCJOm3b/Rf20dT2H5XI2flxXkaPPlfVuVcTjR9gyVAVc6rxOkSprZ
hl9JHOMOks5ILzmGasUkqZWROohrqzchw7WKRRfTseKI27rWdyy+3y9L1fJzKe4/lgK4MZPIJXoV
jY6byfBUK8ZNaZbMYLoKrwVTOb6NW1gMCQlYiRnEtgI/6uxv1n8t+GfmBIe/skXCP+3ko1R5P9yl
IIRPe0Y84jikzCCC03i5Gdr8NSobge8zYFfwnLnhPQNoljcdPH9oFuTSfoF9pj7pSgIFkVA5GXh/
Jewcl+IS6fM345nV+pqvRfIyc596IxXkivisL59eJa7jZThCH3Nh5P38SjTYdQV72vpQoxltad2r
Qs5hOZCY+GgBcT/jFhFfVJeiWu7WxeYZubsAvYBlzRmfUH/jiLGmyMXF2g6gyURE2EC3gFhi6RUC
VVgHLDfIdiA5bgfiGnjjzBf8i8ioXFXBn9bzTMuxwiTY/CM8iJXxHfrg6vKGdPYN1iuYX6RPHwNo
kAVmoCh2EVy74ltrd/6P6LKJFfk9JM/cbiBVTb+sBuAzczC5AFA+jZ9Y4v/fFhsFz7gdwykDUS9N
AWWA0qBNb8aFghdfZFSp0iNHPiotbnPhMVQC/0ripL+JC1KLz8DXU9tC9m16CepCTrRKKdPBjb2h
1G7g8QZuhCY2mYLw/gEVoNzP59d0k1JK+KzkPhN970lvdo6Zwic7geTr2o7eWGNJ2KoXXERjA242
xA66k7+aItxEpuzaC4m94XbzzvzafZN8EAHA5xAGBtj7YQbz2lrq86bxLpCLHcThXhKM1biBM2SJ
RtqnlYD5qKooVKRjb8YRQ/cvSPHSA5aIT2cwmW5f8rNxTgyAB3DalK8nCgeZQdD52v/fxQMkD6/z
WZEcCu4BVA4Tv+ikM1bDzB31YTnOrWwIADl++7kfw+8O8ffPOVm7YBa2MIjqUacY4oB56rxi27pK
rQvEtcinAPUxnNnxsmGyN5oIkfjQ4uiRKNKabAmCLVE4an79LtaHesKY/dOkAwROZAU+epLjTDzy
OshGcleqvr7NI3O5d5VBWRWgg8GCYg0kuM4M/DJ86Fe75e2d8kT//KQM1lG/c/yztB86DLo6MQDb
bvfS+suDEXm2BN4+TQQ1rpghtWRdj3QEb393+PTHnM/GxETAWP9C+Ce8ulKmi7v7gksGGjn0u7RK
HkYEHxutDGTz3TD6+qxKYvKtuX1TL38H8xQhDi/ejm9r9+Oz+1Np5CvKbq+pj2vXUPRZKyvs4iWw
HuJRWcRbmKHj3muT89Rz68i5N5tlQYa5/uR7xaQ/BlMSljFVn+CaXlLqTJjnM+krvvM2DagRZSkj
U5YSQ7f7V8IibEeWMuRuMuUECOP6hX54CMSQ0f9T2QOaiwRnleQlV3QOjnhN7Br0v+8pXxcukpXm
QgC4uwIE6E6Szw1wA7PUrc69RKjbld7GUxOO4VBpyv1YlXHnSVx80NjZimkYlPKT95w/MN0OFiXn
IPOkIA4viFzcEdOLkZZxcNLuFFi02uG0Ks1Npn7MF2u7MPjs/i762ctSmm8pHSBKuQyOSTzohm+i
IvLUgeFfnCwFs3Mv+Q8GJODcbKc3WK8gOogwNWxH2WAA9U80n0VG9zcbWxjED6feS3hIiT7Ek6Zg
x9swsEGfa+kzxfKa2XZ9N0jQCCpx+R/1JbyXussPBJ0IkfepWx693laG0zopYd2QCC6vykARwNxZ
Kn+HaOl9m+ZXbENLoy1JTzIfZ/5mlU+f8uq0mnd+sXv0CbPjRKYn7kbdqL9DJNsm4qP/ASTWWEe+
8j5y/O1nFdz2z7c6ctzY4ChEQb5DOyH5ct8x1oU1VX9An4nxJuFW2KLmF0PK4KbG8khSylfMLso0
So3zsMRjYNhfq4+UQU5R5ldSzmeMrNBrEWfRf2xOjdeS1fybnsfT0bjG6318YfVMfLAYMd2QHn+g
LUEEfEPG7LnY5mxczq7OZUtszdg5KSXY4pXmYxF8SKCWol7WyVe60El3ybpnaflMWQ+uQHGAFOpU
K7FfJdP+IBy3Rm7ScWG/7bsP88uMSomunyl/zUY0ULlarHQ2tLkvaQKhxfatWZ9wN6KCynY46hV6
Nkl9rHnJM/kXEYAyjpZ9IXFQFrLJPsPMTwZoPtKYM92qXSxrQLO9yOuX2P69enziPJqIIbZIVa+F
b6Zx4sV8h61rw+TjovKS40/ezKYcutezYzCm6Yqxq796eq9en/vZAc6450ZGIyzZZ1d4/ENtuwbC
2d8azUQ2qtUDNoPS/k1MFA4vAg49vt9nndoAuRGiiQEXLJJH00Xil4AvbCF6KPvVA99ZS3F2+b7y
hVp9mqVFWjGiRY80ija8xZtEMFoHCqnk87xId+HOKAj/6lkqavSORTm5tX2ltyUrN2iJ1LuUNGVY
x8ob3UXZYwQzl2rm1XIUYl73V4Uilh7eP4rmuZ2rmg2+KdkWCseHg0K0kToxcXtgkeT5ZL4v55+a
YDnr/nr397BUi3hPQkMUaA8/O3f0l6sgObo1kfJwIKyiUDa/gpiOMCopaIvmnmw0OAbKkN3+aNMa
qd40DqgPkjMMWSdrUrNxaK0QuB+wPrix1KJ67w5m6guxrw7bM7LmzYUYJJZFjHnnCRWBTNdT2yzE
Tuw9FPIteCsmyXLRf1ZcZO4JHx7NR/zOlGG44zvC93fYGznmC7FbRfnOsAku7uGugOm/5r45D77J
OUTUSYNeK5Gl5StGhUlP+tMseKnnkkONmlDZ2kc4iH2RWxl1reH/09wPRPLU0wRnjkhgKiudoBlB
bWTIbKeUcj+CTi0uX2noI6cqtr8ZEjNF2i0dDHR9rYF9gINDELkdi8Q5Etw3ZcMM4e+cmRV2dE+Y
J3Vc9n4JYJvqxZsG0KVH7tL8rqzk1PhBrbpverQfg2f2uzltNKn0PoCtGAvPc0vaWfVc/xc/DsJ2
HdIBawU++X/IumaNuJqmj7TAALarP+wNW2WmX7C/wULctEElHjFNGmn8drIqGvXI+XLdXeMFGatc
PWKK63bIAxvDxKu1oUCm0+9MYyqhVTQl6b9DMPvA26anr9nq01VrD6d6oRyaBvlpvn8s3MM9YCm4
Dj0dMXhhw6d0KfintNvdpa1QDeiPfy69VDM5RCedKfTY3Nu0sLn1OC30jpbmRgVK+jRD+XMk/0ZO
eFrsy+Qfdo/1031zBRFGsJE4vkkPAiRKW1UZB978H/JNn2ZQMl+c7jCjanBL2+M38p1j0rwa74ra
OPKb3ZmCP7gHyNQ21xT56ImVbTJwiuHalHbXnPGbT4/4pYN19rowN65TgWarvMqMdhWO3afZKwVl
CV99hx7TRw3ZmgTHXLahYDSEZfRUKQ2KXR2oRVKxbB3st+ppQ6tYbAfHtnPbiawMIi8HeH/5mU4H
u04SCNQYPUP/1cpHt9S4WEyCcHnxLcUWd+dOD7febsyTULdjJh18sfNTysG0whc5FrPsEHIOe4Cf
SZjgtS+36rBj8BnvL10gFMtBTVHuZIkV5W2eq32EnWpW87gBNba3RaLfJh7V+NO2tEW93Houc/zS
tiXb2NtqN9Id/+sBLt3Nr19qyL2GxiPr1p78hzkTHIQvMFBMlpDAxWjzw/umrk9iffg9NyWR5mXw
xHL1g+P3sBMXy6qAJDXYjTm1qCxMBlEthSgTpkvbbR1btnC1WAPMwrhww+Yij7WbXermcgksWKG1
fpEQehDjOYgmAHkmBFlfVplISOXVsec812pBLMJicuKUW2SYpYEPHtJehU+C10zdQ9lh7FWR+Gn3
XlYZsgqPUpFPPEGZpEMEKsc5dzBz8fevG8Cmlzr51PI8FX87yzLy3q8m3Rwi5PyPnIZBmLNKXoVd
1HdhKZNRONYJNhMdUZsSTi5TDvYsF0IIeXwMDiZDx37bnp1Y2xNVHFCyeytYf8mMUL8HOUC/fOb5
bp267oLzyePDMld6xidVL5hPK9ughjCpiYhN3ijSSTMcrMM5BH3sEIsJ0SJu+vmFFAih10cC1jGO
HB8Yk1jDin16T+IrfcNIdZsjY0qv5zJbpyNkalnJZVdXxJNtpNg+G6wPXyS5bLWpeQj2qQ/yIpsN
8yY5EHPpzvh7qU1wxyrntLWwUuNcKH35QbTNyaDdP5kPOX2TWrSrUVKqJa4HeGsQ2lC2GGC6pyzp
DMblgo1PWdneJpnQglISD+fs91q+Luj7IjaFvX2s2JMMwTwmfMN4+emO/SfitvApYmKn+LWtwwax
eMVVdHgQeGkaaUrF6BnNZwPhlTniZ6C0lRGgy5pStvF4Pe9NZRSDxEHhWCvwcqm9MbYXKIIK/dEt
3JHFma1pgCUYBMvHiUP7vyjQ9Avi/Bz6gQ83BJoA8MNwAl5/QdpSQ3IMXyL5ZLPWXzIrdNEN68mL
vS3Hc5Mudk0tbIK2QDNu0Quu5OpC2EnFMRqBEFXG8aGRQDys9T1jsISacEGRg+335vorLKdPwFRx
/UcxlryK663vfADT/5mweoHq6fJ2TXwbHoyH4M1IUo0Vin7TzLXI8xA+xB28cMSJwbjGaRTTKKZR
MbB7uLYmanas0NCBSNN5aOynRoiwkugXdQmZn1LCa57kQB6it5pkY6C60OPHJiNjeJNy9HrDBWzU
b29j0GQKG6FYco8sM2awIX8rYg4N5SVizTUl3tkCVpfAaILsZPy0tfhDTb8tyiuBMcDbb3Br/17m
v70tBKXYRLAGc4joKqJZekz8BbAl69yVAvaN4s7oLOuAUj00edwAdTN0IpRTf8duz/QRsPsWgtBN
PHZkJJ+hRxanOxOWb+VG8i9KffECQj/e+R1RfTcVhgy4mr7aJ80pMl8jMIcXHYRxQguGBuS+MvP0
EZA91fdSNkHiMjL3x11txyTTmFt2GTRm7yvRcGLt7KHOxTNqbrz7ONu7doo1GKj0nYd9t7mKmINz
qdrRQiRr1iQbKLqJDUL50SHYLJ/elWKpc7MylV66N93P+XVmkfhOjibozSXVd2i2qFORrUNNDlCr
4Bvdpx/xa4DCp3AifnjLyuB2iJARTOV20PMswnRXmMorz3E3ud0B5ZVDWWYEhwAUOX6bS4aKKzIO
jWn8/udU0UEr8d+LOaYBMFQCyGzUzUHbJ6WRImF2d9nApt6huP+X6gQlFYXNECM0ptKasIjNJUO9
+i2Ka4yPA7FA0Ot3nnLUAhFDThxROgDPJhy1E9hD0ml7XjbReMUuiw2jsRzP0N21/Dgus9xsOEwe
XoOe+vfS2i9MODH3opwh2ENkN/lPwxBlgrfwZ5L1zVRSxgxjznb/HRtt5ZunOZ1ifNsTlMH5GdYV
97TLoWRgYR+AhID+PMMOcfOWNc3cZ2ZkogwiFreHnCZB5vbXwhgV41krXZkk5m50k3cp80bwVP1A
d6kkJW2/PDrQR1fREntQWFKlhkQ1fj6yIIxLOWYEFKuk+BGul/CxltkA3UcgLgsBb+Fx3PVs1mFH
iRKbjJuCgSQw7WB0r2lQ6VPQfENuxBf7wZsV95RQcPqOxAETtXxEwXXCQyl6O/CiNvjW+NJXUCaT
cGcMFUR9iwgk4XIBOoGjyRXQ1ML15nOBqAYGmENuHp954DJG8397Rq9si6ulZQh2h48rub0TPWwU
Xi6V7Lv+I5MZqbd+fam17jRpUmtYRB5dJgU6ZXnLXiuShZtzBTKVwqMh2zNk2KSSuPfmy3pN40W+
MhpmsVHqzqnXOI558sss49uQIu9fpZwsKuJo+vfGm0ZhdC7WtpZv0+jgwDLbq8R4P8SbcNHLk5PM
0fy1+9eV6Wjtfcr5KkuSdQAk+azjoT4sqNRCkvsuXe1kxCZ/1kryajO0zSuCaK0kYuEx3KNxO6lC
00XZ4bvLVvHDQqyqv4AYDAHyghDdAISyKl869ir/slAC76hjp6uZ+QoaC4gh0iFshL4BvcbNC9z/
tUozOKDhKef8AT32sXu5+Oujhw5vTXFkcU0orwhCmSVuxcUplx9cU/f+2I3AqremwdxVkEKKEL1I
iVEokuYVEiA+3Iu5eBMV9psCVsaS+g7NX7jCX8BxK92e2gGUhcR3ulHb1bkrdBzvVC6LFRbJ9Hdh
8rz1dahxJelO3lXa9c26vhsrRleCZ9odS50M0hSLS6v8US97kkdFAbqbToQ9m8E4abrCIw+GJ1z8
WpLHw3eA6FzzbIY4qlvlDP4QF9JbxAqqiwKFVbdBRRjTP8KElDOkZcdzNfMTb/KYeHF9S4Oxu/u7
vtNuSup2aeCFzIISH69TNnM3GOyq25UxyjAKVYcc0RCkijOowN/5Td9VYfAUeYBnS7xU91wcmp9/
wV8V/jifV7+Q8CPihwyTkl0KjlVIR4BLGzIGNdSHAusB3TeKW4dtGmknKxTTOTJlZTbKwerTlPsr
vEe8ZWuiaVRLs9ZWKunsLef+M2OLxxRCXLWu6aqCBjHBe5EsbId0aGqx9FEu9yxvNSaLPAZwZ7Sr
EyzsWW4a48Uh9Gf/Rhbj8+6N+NEzY0ba1TA52BU8bPDeca7S1zcecEjhrU2gyfR/vbm10URHHHc3
uhoaeFrwzh2pnOQKx14vrAz+ADwC1nASbMN+ktEg0vS4NQNn5QA9irsxjkjUbQDg2/bIXXrPPW7i
ECrbE4fLZ7Gi8qnvW2/LpB0kFleMJktgd5VUQ7UPBkBRr7k13c25umtMNjV1tImj7v9e22uc5kOC
PCzBcMG9JiMPSZGrZpo2VQJ63YK2W48cAFDEHR5Uh80e1SbcsiWqyJdnEO4lx2bjRiWd2SdZUfI0
t9pk/7wmwFYAS+L6xiaJ60qDegjNMutAICHv5a19HJ7qBZOl42EzdG0kymwlYy3hlapiZLZsjSAA
9ch0c8r/4j/8zlDJD7FESNzJBCSzUJQXmpgL/CzXC3Nwirro0YMFRMuYzoBJGGxMhaghNTFug4QR
K+WSFDnuarISLQdbhLC993D3RoPHzHkLMaYz9Emq33+vOHApFUCT82IJLDfuBotWmCJk3Vbv+I0O
3n34B1NxINkstczx7nfH+foIy7F5pnT5o0qVand61pcJA/suhSE45WJbSfkXKFjyjVbRQrac6I64
vmo5gWewmoe8hG8vEI1UvgmZphraGDgTx612MCTHBS7XpYRQ4Sc9fIcZHmq+emWx5dQtIXUFqq2O
DLXH3ugLPNuKsh1L2pa/jW9VsqZHh36rCegrotOYz0kifUaSjIiXo8xkH5FES7dC5/+dCGNFrnZl
9L0my0JFvScA6awdv1NIarJYNMqFFCDQR/PnInQ6JpFFrcq9mw4LYQKh5ZnCpNFPjLotgLMhtlCs
3pVkQJNYmFKy4rvQJvzx55vCFGqxe0L45SlyA+ffIr5vLCGlchIY4kHHMsbIKlB04lC5yuqjIpUO
bO7dX+l3HT1y36RRBieQJIiQ3qpVt4ye0oBji0NCSBUhXQcac8XEux5IZEjXKuvee7kxfzLZqfoP
panbtBbePHh0PzSmbXG2HQc2/7tBfUVupi/ad7fKA54e9grgabqdnlQGSho06Z+vQkmkw5XRTk7d
1gKN+LtjFd/RapP+vEUpdNqW2SETd6no/sSa4gysZWKU+2LKcO2v/Lff5amzKHzQ+xkDLAAuBgtY
4WpoxCKybrkM6MVR5rH0q+//zbNNnU1G1ihFWW8rmEvoth4yOrhZUzGYL/Qnksp2k3TPBuvXjhR3
K8owdnWHFtoIqA/FioF8fSUUqWrlAwu5itFa0jVbXJCzVZpvK9XlenoD0n/0iZroJXirrnal1CzR
m+WCLdOVX6p62zUanEb7HuhhsyAFYv8g0LFAhgYlsrwoHKYhDdQ6fPu8kvFxTh8YkV8tFlAOFOzY
QyphT41F2uEGybH8PeeI4ymosBGei8bEi0IZld2YY/7W7QwY/24xbGygf8Fa/gvwjx4jv03FNbfg
8RBfn6v3qzTO66ja9OhmxJz/X1FTL/WKSLL2DVY2WDjBkAeVGOi98cHT51qno9K6HFm1xd5i9t/2
czwGKStCWKO1TaYxznDzHjyHvJAU2xoWe75fAV2IPWyp9wYpsG3KSSpE3ei+EV2wqWQeFqMAPknr
NWerqA2h9/WS66A7O/z9UgIZOIhsd5nZnm+q0a4AIvrLOZjrG3uwZ6jZsN54YsllLtaDPakcn2Z7
rO64IquRasC0nTLsCTlpa8AxkrFpsFMDId6C99tw7ezZNFQodoqa2wJ/qNcbbuz0LySi1K8h6q3u
SO1tYmj9H+TydM/gugyIe5noWJrqM2SgtLFf0e1fCbvKAXErVdiCupzkD18MhCyM7Gz7T3ZASbaI
Hx2W0KU1okiASwZcWVHagPN7+65QaC1gBUGzpoQ0WsK8hSK5ctXVPCngqyV4zL46jzO15UtrNWq0
k6YRAENQLjUxLq9CdFH6uj4ziSukpTaSBRbZS/gBwqL1itmNaJ/YWlh587HaBS3bpt24UmsXoemO
sJowvBQNj4r3tHXqh5BadJP29XP7jR0eEAz9G7WLe2phfQsaPQyBB+TP78wCgCaYitWMgrxfiLQ6
d52zDwjf623xZiJ+hFf2f65zTSekTW7bchrKPwvGdBHDLmdQZX0aVGwciL1k9PRmC/fcdC9mhuHR
qeWp/1W782a307vR8zBjKMhkj5l8GU5CtSPoh3lxLFXavOD92FROHoVj0MS21P8x1regl72O8tIT
8xpFcwpln7tvZ6uVI8BB98vXRhXyF6LDEA/oMHnYM/baaeZ3bJY8JmO5ofAsGjGUPv8H8MPXCIks
CpzN6DyPvLLc3l0DxCUIMBH7g/0O1GKRPsTRKQEhyGvQHsE/C8w2kJ/MeajapwEfhoIOyqNZMLlA
WqyFdxkCtxQG4ignlxOyMo2UI49e+BD2xSPnWft8UIUPTuaxbbfGEbqenDkxM5+kG0MroMnpcxrs
C8Z6c+HtyeTW/SihzcfR198C3+nMIiVpn8Rj1CH9ZNH70hg7HI+EsLebBfqKl9XOPLo3Ua06+5Mo
Pfw44/WKu9oORfcDc0KrgZJzSSYIoLXgkhXUALqA/7qACs1aoqkjBVOPUGplUWUwET7dVqkBrMBB
4/LnV487juudC0XwUeKiuhGo+KOXfNC6M/MPYvHigplkGGzicqym+h2oQXrvUzi6Q6khugu95vyO
uwbPWmPRYt6AgDvMLt/Om0GHQgvRY9JqXX+IxdGrzjP2bThav/u0VxJwICOQQyzKG5vj00n5B4qk
Qp75kjC75s2uV5NDtSDt+SV/FIaVZxbr+7JR1/CJoOk/JHOrndp286Qc4MVOiVYbOBs5q4AvM52X
NlX50V34KtyXiDecSljb409PUrIkrzEAd1fawEecT4cXlQNLHgcsxHHr+dt4WNBA3+8rcY7t8Bqv
/83d5L27Rg9c7WBIHizBpKGzIIX6F3DYhTB3H5+smMufJuwJqMiuWg8Uc+yMvWOE2F1J2fr2pcqX
uVdtwOaUkPjLKZ3TX2dz/EjA6x3kouxIvrH4KY9Xz81QRuQ+vVLM4Z9kF9TkKN7MlyNOuMtEHyzm
TJ42oRmEFiZCZG0GvnwpDEJVmEJlbqp9aw5BL3WINThTwn2edWa2iAFjRFqOOkw3BoRMUMGjlrPy
rVlUvM1KrAgdV6nGC+EnvioE7BbrC+gyGq6ttCjaAI6e+LijEccfYVscpDPbA5InzjilXVrverif
iIpt2UlaZzBcuFV++uaZVm6X9weVmjekBKR6Jjnkxv4xi6ZpJXXkVIFHoJpCt0BhMa20+R5VVVSp
jlQNJQsfIL1/JXSyyn2thP/s4x8LHThK4iqIL6SAdNKY8m0AZxhabZlUyq+luyRutBm9ksMXPZEB
u48g5amn3g0Nx6XL2x43iBMYvpKxodhgs/O7xONkUpqdMf2OWetefxa57gr4eIcaw2Pak0Sw5xm+
qY3OBAVBoP/VOcJl+kBGaFgvS78GKiA11uwGDxdDWjWf13MVKQzVWTZ10K0YfTxIwr1LXNnFeymE
VJV4PrdQIEsjI4LogVbR2HaxsFxILPqPkqE7cU4orf/SKgCy6veJFOiNx/cGk/00fDhAeJR80S1R
BVf68iSeXGVueRjrnjkrYQpzVCTlp9LyxIzFiDcqhD6DNJ58PFzLvHxzd9l6zAVed7/JMyVNASy8
03k5MXu3s6s6hieGyL1+PM4UccgsPdkX0hJEVOWWzwQnE+kCb+8d+UJSti1Z1LwBbfM2O4z6zm8V
haz0DdZ/Vd8/k8HxETetQ97KwrBFSCQziUIGCj27J0NKcvyc6Rp4Q8KNA+ARgZnHwnfFB2JqveqR
CAk5ejR+QNSWyYammvkRQy8z+WTr3KGtAtooGZVIpxxCIlUk1GDcBAwRhf3pX4fo9LhSTQdbzh4x
GkHlt6pX51cH6Y2bSifNIPRRjLM88UjBUvBDfYeCf2FSY7j9+qZSjvFTYfn8pqwaH73hsDzONz1c
57/g1oW1LBIe4pR8GVsfl4GFL6r1uEX6iUwdXo8ZOnN6y1N4AIrAwi5IO+FT6rA1ZHaXS69FOQFJ
jC0hxkO/qts4PdSbQjI5MKeKYX3ZAjy86V+DKsmRyOVIxoENZdZRsj8ikJ3XqKxRrIdCFOjt3IGO
2eN5VMH/8m6NBVjnUkLjR7Cgn6gI6SqS900WZD3OUATepBnT5iKfR8LqpA3G8N2PiYZ/8IcSHumk
3ydRYLJ7Ct/yI2/7nv0rKdY/r1ABqAd2KfTtISNGv4eXhYe0xN9IyNT2piN20fI6kHJTzvXHQKs0
aEaMD4aZlYHjXTeBRyP1Uhx5n03HSugrto+kGIPR6rKSy2D3sDnwHRNGsrQe4y0N3AvAopdwA1l3
ugJDCC/htLQlZURDpJ86ie+taMJWXlmRw9PDOQvtzQ5XSrBoca24TrUuHVen8Lm6sbx7kTYRsyF9
ldmJFxqHa06j3KiOtL0rdnfWvDNW/scL7k5O31pgnYgIs5B0PbTNRuQU3ahfk7WTjEzFXpUyvUEx
1sIiLwlUd0TU/CCexqjjIjWKo1DT1C99Wq8aY9jGGgnEvuWAg454dBzVhDrivQdLlkWHZVTmX5+J
iq08htHjDe4VLOz0mOcyZkj1jbx6dE6pdNR1WKaIXXmLaag+4IVrn4cUR6+C4Jrnv32ptnz4ONeN
2eH2oohYbcCELei2/o43hOJqc6FOXNh7Qak0wdkbaiE23ICQMCH6cf5IJIAZjtqYIlRQGvqJF2ot
aAYyNEfehucBxn0WQdkDZPWupzafUJhQbUKbGpYE5DANuEOanTbmHiah/2NVMp+SABD7wQ2KjoCV
y0q8/HuLweb0O4ufCnw8o7Ly0yoV8vR72CI9ZXph+oB6G3skVZMt1cWh7P395MHgxVFYXHgI15NZ
yV/sJP0OIZm4MkpCLzDU/PfVu1odc5tHb4HZnOIzGM7Ab8ZkVsiqXXWFn4eEWcAtnxTmdWy752ct
cDsd706VqRVDIXYqTEpBGnwmwMWTqzcXJ0O+TEUW0yiyESU7ydDGywtjnFFxrInVZwB3uslSz16o
Ddrd3sPr1hEEYow5h5SzMACyMJthYhDtpPPthGQnkNnAzoRRffal4YiGd4/vvZCVqURoRzcuOimq
C1QZK7e7CPTLSWuqYHbSzoMa0B+D9DaDadKyWC4G3p9T4LScHfNIzsd7l7CSe1ZhAI5NHmPcxjSH
PCVdaOjlR/1OLwWUJWgrM0+rVzcyOlSH8EgWtZSdLJeYkXn3k/7DklFRWcA7zr07bP47uju1Tpw6
LB3pTtUtjy/UkKlK+anF83X1SZJhZqnCzBR5eUIC+4VYuTq3XJy0dzUFGd/pQX+yAch/FAOLPXH7
HRRSifCiOKUdiLA4b2eYQ64760jwMZ3yuvWoPZIGjROZ9lXB1HjqURAO6bjwk7Lict7W/QIVUNUf
yCJ6Cx/T7HR99wBg9aOhkh1SLMripwVMLgA857VwSu7QdzPT6+BmmmvUANHi1/dEmHSY80fOpM8F
IsAhJGGRRnvVX2LcYL+SB00rIWgBioXCKMaqyIGt+7u3Ayzv666k6HFUmBI5odz9aggwwUYLiLOI
RTpmD50kdAbO4gVB+O0IYNDrvAHyx+EAoxEV3P8ZVRf7AANkiL1A+I1kz7XT9qlAuLofcvNX1lFS
LN7p5b8tV23EZZyHjBZOixQLuiQB4KA8nWkO/kcwVdhdNRJLr1R1PE4GbFWdQdxbgLUvhTr+LXLL
LT43VY+TEN1ThpU7XtasfLc9pkDzLfYPgqw2NdFaGe32OzdM0kId7n/nKf3zZZ9TccA7KA11HSnI
Y3/fEvdAWOJnH0NBoY49GcZiG2HMZzh2jaZGLkmwAwEiOOxvuu84qUK+hA+cFt9j2z7vjcV+KQ+U
PwnzNSoN6olYUGwQVG8Gf6KJVKhrxRnp69kwy/hHKw+NnkvlLthGqNAQwUuS/Zo9k+LdYdoxcXh1
asHQRjAYHpYDOH7Tnvbo5HzdLjF3Gm7dwVzqQYSxG46U6FcskZW97KCWFfFjPk0WLa6DYTZfB728
6pc/iWwnrTvaGek2TKwqtuzIbeYEprQO7hIRVE/AT9lwCc8hoQDtswOGZLb9jUi1qMP18LI4jV3g
4GWb3JPsUaPMrcMuZZGrxJGrTSvvLZ3TvKpLli8V+iqY8Z8aB4CXB+KxdsTzoszLTYx2X5MQLfg+
ZqcVfPHgGAoyz7i8lw6TJUFHJPEDEFwcgI69ZqqLc5UkNHsRipkUWeautJpbI5M8se3+BONwqPXq
VVSohs64KZBpKnW6YFbUZwnTsI3fMeE7VP2oh+RABjZ9cOhMXzUsVknRfXeyefqrSirosV21AgEA
tBKkE6P/4aCCMG/zt4M88NrmjMOkWf09SjTcvP8PthVGFtEh3seq8go1vO7tJ5n9nYq+H7EAigY6
2Caecwndj/SCyPDgrDcvJ5M75GTzaSpaUFAhuToQmhDC+iqzO1eAOX+jsmsCwDerT9DYFPEVyKd6
LdqVz73a48AngIBGvk6Vh1FVVffm/U8sxsOdIF1+QgnbZBUAHZvEfep3oCbFwlQVmY6BA5iAKh4p
up+RonHyaxQ/XdeMFhTtmqnObd1ERRNo5N+sW+w8p+C5AnJCwqaINrF0031NP8hJPKU3RJ2A6d38
VAvK1AaUZh/jvmKEEOQYLXDrrHXDkAoCC9N+4zRQ8+1MZoX2r4aIZ1ct+Fvdqg2aSVzm7/vHnEbX
pvAMhyFOMy8TdaK40eA7nnH0QrsmKwuEGRC5Sr80wh75LLAkZAhgGu93c34TSjt9m9K+qo0M9bm7
EjMLsFMRfVxRf2OGZvI5I0UETu9ebX71mNqeWAopuBc112pnBC7tCUv1U9EiJbdAoX+RTQiu+lfF
0Dzbu6XFLl9KS+HAP/lV1Pg7p8Jxm0lzurDtipTTA3c5tp1J/uTOvJ0y/pBJS8zPWUAYR3sA8nJj
92lE131C/H5JqxjSGOYrMMsseFT6e1QbrfcpxdAqfSB9jHS5Rfok76hqLNbWaPqgfeheK0D054pC
hUYEAnwwSw0HckKUrUoHHAV5lvQeBvhDYdQATBV6IxOsJl7OL5cacFomEGAx1W0maeYzkHzNOSG8
VQJaU8dfpgxJOVRct6M8Z1lviZpQlZCjzyXqM2KIvklzx5bpKo+xWCx2IpqGeEcHFB3l26ze3wsl
+EpQAzm0hRkv0VJrno0KzkgTXnmuGJJV/+DF9G1h2Amu5YRLoNABXHHL/JYkxg0ewUatFMcxiAw8
8yblf8b8lOgOs79MoupGIeLw7d5essx+tnmO+6EfB4HOa2WgXPOUF9mHlM40FCFT4Cw2YUaxMLBm
07Fl/De0F13Tm/L1vv9LqnaPGKZ9pHgTwinUiYAZRRgoXSBxCqqWmJV0Qn5uvzzWu/0qbIz5QQms
nYfuZ9SRCEKveIvf8GYw8OJnFsslqiFH5GTGKhKkW91Lkm8UySS9yoFMWexRsYNH/UMQiHRUItYb
S82Uxj24W/zJ2/jLsYmfO1a3zxKJfkuqfJnRb7Bzp/bSGX0YTLyoAS7aipwS5YGwezN3cG/jevlU
xJYyTLiODwXjLeIVXKX8u04s6707kQQZBs8whMWGj9f79g5NdeKegNBKFrKwLQoO+JfUfMNJRgNE
K7AjIcma0LaEH6Tm7kblvCXq5T0Lpd+i4O+fQxZ1UmiCARYgbR5idEGRs1Ub6Ke96m9WSqaim4q2
o7fwLHcUKh/4N9dSX5poJmAH49JOW8mgQW+lFD/D83wdQMgi7mnLUJaVGGYFUhlnssFFhZ19zF4v
linF5Hrjaw1DmMFE0He++R+3gjI5dYlKQaCHeRYjTnZ5GWn0Mer2tYk93xWk9sTwKXgbTJ2buRQo
Vvtr8WHXm1VBcT0xmGWgyXaGpPNudRjhuC+fSt0B3Ql3IsEcZ53RZXgyznZpxO6wSsmphNnjZT58
xmiVp9sBgd/KtHvJrcJbNqra+TFft/80ly3L9RoUgAeTBnHSfaINNSeZP0+qHvU3vxItKYdo4fyG
D4pa5Im1ForPaAhHJKfjKC64Yv4jnuWpgq/7gwnd67/fGI41u0O5KbGS6ElNCRnetFggOS+AjMdW
Ps3JXwjI5RwAjmGtqXI8LOmPCqlG3Bl3SDdjzZP3NWcRGuX/T5xcbi2P92rOE4Wf4r7JAdYMXV5f
L8EUDxu9zUEIheOWVp0NO+opeC4Q4jpu4NxRh4dfuc7CaxnaR6p9kCmVPWLJ+9oP2mWLXBZm4gwB
KwOjMbf2OnIHx5AQMCxbHIX4Xwtb/Qi45KQy2ggGlP/vejo9OkRi8EoSKgIwMaPu8lwXr5e0bgJ/
SkUxDxzjdrrHIGYyjWh4nDy5VHzJLBgSos+hARkxKPJiWPzAaZ1i3vcUqPdULAzkyl4haRpiCP4w
O++g2eapFbbowlsjEWa8IPJe6n5lYV+bOZ6acXn1tI+2aAV/Lov6YsSC8D3yJngJJOXNKmCS3lnW
ISo1CZHmAzVG8UWiE7P28xoWLfmb4fiqfbr37vxvDpXLYQXkCZBilvWGQKut2B84g4/Te3loC5kl
ePZQSbG65wS4tj2rGHrJvYALZFXI3CW7DeULBx2TNncWzSPGYwlIvT4BLlgPdr7HrgdK391p+UaH
UjKuRM6qsGXIAP3E253Du5Vfp7a6EPjU+1SzmXK5OHWtStxLARFWp7dkK78ATdOSxe5bniiTXbIN
6zuRbuVprn+9ydPv+TtPTg+cWQq7YSFZLNQ2T++rELju4FHQdkvxTS3OhGhA4xVfUwW+3RpZNRWl
65AN+g/GIuMn98dtsvP0z4VYNrnxMuoiIisBYgHuTCjRfsWtUzs4B+d/XlUTn3CJudP8mkr4vrI8
l+khpaSwaNRnE86wJ4rjxh+Gx+1qH92Hxalsw5GNbYlPuk7/LEwinWhZAxeaTovHFu+DKR91VvkO
Y4Ta4N9WcGf6joFQwRYP8YUcO8gXPRa6ufbfmsjPGU/TM/svP97yHoiH6LaVioChx2ovpG6Ynp6A
tC3tUMCGs6sZWWGFYVIroW+EQYPlhJk9y7BJDlpCgTqpRnMWTrx60WBANra45PF8W0PONjLXH9xh
HTzEdBEnkPfQQcUvQh2IKgdvnT3GqEyskggr3ovFAAdhxslE1nlO0hWd7r7z8QY3+AZnsPbC8CQ9
2nMgnaW+I91qZpO36wz+Ibv9luJ932W7pj0mt4x/jGw1Rrh+phtxhDRhG5AGWpOYDMy7gLV/o1jo
NDypJqMRwhAEeuUF9XZFZDPcnI+8z1BStU14hcmR5rZgYLsztF5LzB5OR4CvlXpRzIUM3w5ZFSV3
j18mhC/1zWKATzllg1fdllw0Z6wrsBrlcucJWeipgW8NJksBH5vT3qi67cXZyHOuTZ1SQQ22MRuL
JFy+/GKc89bynMT+PuguXEX5JfJ40cC+X4OwpsXOstDBbEUAIPW8Tif8EoMAsBqIJuraRjmw/urt
hkmL/Js2ZmFmPrevBDe46GX0DDH9vv8SaOc+DToGam8FY95bBWF7bXGjdUPYcyOy8H0R42/e8oiw
mpQARJ566QLdFq4sPXzhkVe8fHkJ2wWeQNw62XvfbeTZ4C3MJYyqDxWPVfAKq/rjWAroFjJ0cAfb
39rxwelzdLXKaB5YQzoDu1NJ5HQpDDbd7kaVJEvyQ38fuggzudv2VoaBuIGiQBi5XKZrvsPpkC9o
LpCJTxUaQKOokoXoUS4Gh33CQjiZtZn0Y2wSweElb35M4eZRTjR8q0EfoM2tlohrxbLzD1PT05ba
LVXtJl/T/ZlIyY9XeHkj7a7UL0B5OCvgEEw+MuHWFa7uuiIQP4Cd7L4BOMf1Y2189Ylx1q0ekbcT
aVHoZFcdGBUsR8kGE+BVfGnKD5zGePxYQFrdf3E9cepBj9gOClY9Qelm8Lxlq1vQ7HU3gAaYaRK8
PTuFVq7/lKbAquJaB+qa1d0/XatPF1YWjjBGe6GApn8PrsVauGSrwUdHXdqVZB50iGM0xf21MFSq
AIrHLuc2hfkbGGfYJQR074WGDgUV+Nypl/WQWsBYuA1U0t6unOBNu1yeJ/E/zpyrqARrUPGOI+Q3
ELwauYqkeUwRcrrcRFrluzlRczibaDkgNaDdFKBeXCberCHjVFOvtGHqe9C+EhNuu4G1WtiwVJPU
TIOOafUNsOZP6+j1OLhzQW7MMyCgKMC3EjXKa2rYkjZQSrRawa5PxsaiwZkYPHPR+ObTJ9G2KZu/
lrS4PnM+TRUiPXV6As7YkX3+LC8+XcYIWukwerGPx7w6qKIUt2Wfg2prBw/JAhF3Bbe4Thy0Tkhb
LbKVxBq7ewfMk6YiNQKWGHuyo1bXLfa8NaWPnDV+3Ml/wH/EXBctS7+YEK2QUErJ4aECX+k3CEAa
PCmvaZDu1xaw9q8NDdjxu/XimwaGQ2CtAQEewx2UlP85l6UKd96XT919ghJtyNEstNYuet3GRQRf
o3ky2qIlj0wVm1mQR0Lg2K4tkz/qn7JLrR41wX7YDWAO78di0gLOq/+GeNGf5YQiIKOVsVgFaiWn
m7A68AllcdREZpSU87EwDJRs4gFp0RArZIvnuIOZY4Z1OaNOBSwMCMYvBlQGloxByE7FzBNUmq00
pCXsYgiSvqNu+UDG1g+fDMoWuseBPx24dhbP1TBE0XItvFCKYLfryqiS5DrGwVXWpiGBW+glwM8I
V0M1oTrqEZaD0IRBM7GEWJa7vbrKxNK0gHMAOU0EUgAJsc7ZYfXSkZ0WUY+w0WsE5yAoSF4Fj+cH
VPKkfPukjgGC66rYPNiEcYE9WEhhcnlxDn4e13e0lr4pMjQz1NW+IG+kcin5y49zARPaSGe+7h8Y
A2ShMGV72NUyZexrsEuLFzO67tfYe5yXYYELXD1KWSdDKmzeoiop7a/6pyhGVI1lxRKkQNeuYdXh
a6XPOzUio74KBoNJeRUUP7IE+EX1wfRPLAKMQ6gEd9rHbgOcmQ9FokvnzPZMvHIh85fxQa+53rtk
/D7MEH96g2+vgUSVx66N02jaxs6264V1aR1ygf5aTZTFp/vDhie893IFjMngjSs26ZZpcIhnnlqN
I/HHE6RAVJGMtWHV4b/W8KTotmjp1wyRx8ClcVamkx/6MkYO5YJ+qioJPY3LPIloJpd0Xm+bBHBx
EOWpMycyYPd81w7FUBOE74yCkON5ZkQOIZqOtALgRGf4dFj9rCOOpaOlEfdzwpEQRf/iTZVgjCbv
QysirJtXEu44YggtaQ8bihE80g2Xp6XobWligT0gmFSgGBnNaJpTorCv88Uk1uKJ3bSo/BDEzC5p
A16sJZDtijvSYR/gBRcQlW1N9J6nVn5Fu7u2ISroGH9OVHwCOmp7RqqooA4z1i98WBsGEcOramxG
kl2EQj/vwGOma7BRqiSBDWm6r5SMLsAuZsVBOHG+lsqZaDZaVg6SRyz56iRminqaUco8pUUEdslB
5h8DETbHpTN6+653Ee3DgCo0VKxzq/7bmvaeanr65+QTUN29XIMUOUqXdUUhrYqc5vXnf5O7YySS
smg1sBaMgiVx0I3QtpDApADbF6OuQbWaBgCJICs6xnVfFcWozdzshyZ9vPikwExjTj4rMWaz4643
yjkjRA/zEdJV4JESDubOa9915Kg+PjcaoUXNo3CMoJ2vVrA4RKn/Y298JQCb57Z93EFbwFrDtCiR
HKNHud1O5ErpjheE4AwFVhYn+BBHtYPZgAmqcuc0OYuN0sDcXv5XhV7Oo2D01bu169RpYFgGmic4
A97DEHd+fy4gp+XhGEuSIRQ6yuVw0Xo94CUSQZ+T2/pkzurEWkwOLw0JGyA2yBFlMn8/apVzfRvh
8kgXhFinWgYO9KdN+xaRCe+QCapMsbEx5VuzTnNR+xuT6qn5xENz8N53mmMfn+F66R4ykpaj7wWv
0bWmebrsRi1ZihNiQrCs0/KtK0M9OXRUSSegTXkvrBcmEOuW+9F0PI3PGny08gLGHVygzy/J8xgg
sX7xTNs3XAH9SIKWXy1rsQaKL7Xy54nQ9RR4M0WZh51pB/UUKyGze7FiihohhiySnFPfKi0a4k/R
gAa9C7PkhEtkRrhEq6+uEjTK5vC6Ww2sHKQixEtYtqlrqbjodmiCRQXUF2AgqeGGIpMi9I3rdPR9
Ci592Q3EgNtlESRQVf1t99Ptr5M7v4pyObPT8sQAM4u0bGLwkdpZjtk6Ya3vfXZHv3yMaJ6/5EpK
ht0sp9jireE+5e74DelbNJXTMSM2VCoSBCuAJn3pPCIHAfVfvhyFzutMQqsAFdic9NcBvpwu6V7C
SOOGhrSO/wK43AFVgdhoiCsIgY+2mvJV1yqwD7CTD3ESgrAaudgB2SUp8kuQ+r8QixZl0AUsoVTn
xY14mWFMoEhVwrfzpkjqlGWVx8Q7nc9WrO3pqNmuN3hsntonUPSXc5YbId0bhgUORk0UWVuRtCnx
+XscnD7H/1+VUOyvJ5GXTVgU+ID9HOu8gyByWhRHbI46C+i7A7r46I2k/viTYeQxAClCLaHZI4do
15iFQwf6WiiUvsgOWjoEfrN/p8+ZFE3ciBz3P1b5lEEvrlkLARMJblQ2vqHf5ne9RzcwqnM2pLkx
O+ak9dyyjaBJerPJC6oGN2nXMIHzOjBMNxgT4+XfaWC6n8LpWEPWl3Vffo9zeJmkTF1caxh4M2+U
9+FFCXTDLZSUyaAlvCcUwDI4bnNxelKDuAFXbe6yr9DyioePC53K7Q1plHWKfJRNJSPFijGCVQAq
YPMdD02RbqqFYr/DyqftYINetxRyDzVSIQ7xxT9pyoezwVf5vR5bcbWTr6bG0RhVj/f3v5HPkuP6
Nn/GOrDd2m1quOSkYKcdvM6pSoliL2YNKpTH9H4iY18pJHkELjtXWDkaYwV6VptkayHCaEvA5ZcM
1PR7cLX+whd8PgVK4SRmyu1xZ5GYiFXvlhvjZrMdmhp2osO9hTSpco3vsjiDDixIgtmzxpB/AEzU
1IPeMeqmmU7jdqcWSi2kMauyXSj1TsrzNrN60EvT8x7GfJ5x1CWFs0mSQwLUTiqBdsFZDuoQIvm8
RHKjmZ9ZyNVk4ZpvWQPm8zbXoBHQ3r1GDX3EaUOG5+Xfsm/tkMB7CdidzbBooe8w7z5SlgDgBap5
vJKcQX9hc3Qag6LvD5kQCj2lXe53+BWGGnxPj3peXZ9Y6pz5RayB7YNWczD8xH+2xUctE0wZK0vH
bmkiD8AUukbu7rgPkUwuhr4DujwvD9FCFcgPDfFzgfW0SPYxFHa/OXi5/IMKVmYqe/ZATn9Rjeb4
bB044CSHOmrJUHamKTZ2V3mc76jVKJjDV8ieaaaZTvPiXnqmBAYgc6um3iBbX/fMs2Ku4T81Dixz
psPb5zy8xkevL7tqlx/wWchY2Gn+6VXkXhw6kuGiR/ou+Vb/3BhJANF7oxt9o9i32Jn1ix2g9dsF
TqajW/YPZa4kVUf07oXqYZPQ1zQwp8S2PMFs0B9RG+MTt+LigGRsNwPyC3/QrS6cN4f1sM8o3mrG
K6O4wGfexHUzaEocUd+DqWAKcEoY0JRyxCWhHqv2R9aYAZSJaytcD2HlJH3yyp7rzq6y/ydBJLsz
KCxLGfQlVE4gKjHgTvaXuiog6SyV2MCKIm0P6DIG5XspVNVxu04MkJ5zNCbhFs7Qn1znTOO9q4uH
2pmUEOeaovKEABPww+IChwLdfkysgb8TH7rXj2EZXVORJehIhPLp0KMnCipW+2AgYffBGprfZ5wh
i3MbBqXFtToLDvLsuHh9kqNUy2qex9n1n465ZDJKDviJ9VInSlb2zZqxSGrSnrGErI/kSVdUgZyR
NXDXK6xJ0HqEHiOpwV35r/Vn8H7N5y59ObJ2edI04MRWbHYT2qoOinOSphCP62dJT7HSEZha4hcN
SqEBcMtkD9QMM+oA4MQWchPuuU2nrWi2FQJu/CZMeC03NTIN1bhwCY6d1Y3i/C02c3UU13Dp9CJE
BsTng8WqkC9wG4LyW4t5C+j2u2a8ZiUi04T632cEW+iqpQ48mtZWcH4PMpESyhFOupgkKtlVMyRo
B8F+HsgJusE96Vu6H1K0b4OWywhGqa9MZ7V67GtgmxZmqdZACzaZnALEeO9broRuJSg58zj17pyc
8xiWU9nE52Y12kTa93VXHGv4whq9u13m9jm3K054Xm/wYESbA2bH6gTMNQtv0AyBBTRkZD+QA3we
XM5VpBGJrTfCnmAu8VXgirAcUP1bLgKvVnNR/CcTVuRmTfQnJ9gVJmeNBQ690lr+RTeJJtfhwhYQ
oobtRIcZu/UosH8LbxNHtOlKr/1dQtHARmILpUifmKC/A+LrFeDLbEI4M/gM0B3nBxJgjMQqTZLb
sup+C5tB6lsqSLqutKBIONKG5w6tp7/GkWeA45YM7GW8JExFHkTWFUWmKTw6D/prqe9nI9GDkpMm
eO4DadT+qw5dH7vTyIWyRfaMNGm3NkGp/JxZVp3Q7TrUdIJe7oO88Wd/6OibxyC4h39mdtbsgkRO
RU2zk2I3BrOwaX0RbqIr/31USqBS/YA6+at3V7C5+YGhMmakp6nR1VFqOW0roj9GCh9J32DIaoGV
WgiRCge/bVTMJ/L2OTB6C5nFCTf9PQZcg03xhBXASKcnYR9T63KrWRYx58ppc8cqjR8YZHh/87tW
6efL71+zaj/lxEvy077LlwgeFE1VlNx6k6amcfUcaF01s7linrM3iLqmQXJWMf5uO9PdnB5oYtDg
7p7nNAXmMwO64qC3BlwCTHu4IhhRSBhJ7ycw6DwCLEOzIezaOzm8ywrYT0e0pcZiJAkpaQJBla/a
XX0wydhI2KKUv37NSm0hm34imAPy85JQh91Oq9NMCRuDguaZMM9hbrIVaUIS7lA7NbCoSnM/XN3u
j/18xAicy4ZAn6eMMxNFhNACkB86QUTA76vt2IyEcaXyqp5T2G+BE1hTOW+2K4Pv4clHuy6m79p+
5bIOjFm3Aqy+3b/w8mFDaME9fgriPYPk1xUEVlGraUXA/8mS5R43q1IlZjvpK5PHFUtnwzxHfEU8
hkBqlU5A18lfqs0v1xBMHVJa4KhDuoiVvXl04oxWUlZQSllZaZ4vedKpPVnnyn+q+CbYiKw2jAK7
a+FcKDqv+mwpro4WuZUdQ/r8+DKMVg0H45gnYNM/ZanY14T/YRtWfGwoLqAOcYGKX6gcoxkb8hTn
a2DjOw9FnCJlwvsMbQFy5T6Z3pDJaPUbM9gSZZYgb1OCoqVdt4pLieum7FZKYHwFN4hpAsd8n4lO
eT140l9bm4HgvumZgrmGeOSd04YlsbI5yZDpSLsObFEOfnl5XIJcV2BlRKyUn8C9bt4+8VysPW1s
2qK+0mF3rwbhgauvhb/8B2keDPkwFokpGO43C+74mFKAmN1sHy6boLTnkfA7w19KkyqBn0uHM2Lg
b/HZs/KV6B6ICSoBqPiyzCoF1ifHcCSXLSnCnYRSWfgYDzjQDAX1+rxr2QnsE7fcQNFrGggY4oBB
aetceCb54lDpzKxClB3/32gggcNvI9NUhZ7ueGl+SkIz0oetwM0G52QKYxMS9WVBzYqfRx4/pKEj
HWlg2T0S7Frg3nbjIcwRlgDlGple8HswdIljN5C5ih+U6QtZMze9nHMFSxH9d8VPmA9dXpSLhVi8
SZ36g6xYSlqrdBJ/GeDJcWdgVbDm3YwH24m8ps2XXLXP8yTte/K8YMti7oqr9QvaoLstlCNT2Erd
SRuTgd8nG5Y8cL/owAnURHLlpgAcX/R4sF1h9vmmMnP3T6taoe/AVeV8PWDjHrj+xg2hm+WlVv0i
cKt4QA+cG8rNsP7BMDtMHoFg8E68F0heuxzI5u0DpUpGaypBK4izZOlCUiUNwA7cSvhVRresjWhS
ba6fFVt0uYZlkeS6oTtGEoh3BPvvhMFYwPUw+4LjgJzvo0JAhnJEjwVTiYQztwy944PzyTZFTF+C
RfHXds2PPdD9hK+6fnGoPfdyyncVU3Ezti6r5ls3tPTHY12v3mnja6qRheXVLIQXeD2TXGqg+B2o
0T7HbV0rEMFX8ypMoLqXzvxX/HHFnxA8uDeMT67C62zBeMb6pXilZI0rMI7jxQyDoywd2eNT3W8P
ctLd/iN2cmPceLQDUo+/2+nhLWQUFx0tV6/fE075B5+6QMADk8BjNmnwnFx8yeD2ZErVpm4P3H3C
BSRdv8O87OH/yBk5/vEFjSitFy6+rCS+flxP+nPIlCNdnuumlUta3mktpl+bkSKxCXiniyt9x/xz
1+HqGgp91oeSwpTsdPYL4Ig3h8GVOYn+0IdA4+IErXQKjHo7r/Avr+jnbCKCln1DYamxOw2E6W0O
J76c5MaFIYXa7anvNHIBhacBrIP5ZVRIeY305ZFpz1ndHY6xTc4L+z/CwVEyzEKiqGH72WevisqL
emE7J5ATiJJzTpF92raOPFsiNkyIwJMzoADFd58/9HNShAFqVzaDusITUfrFrWMo9qs7p/LQh+6R
dfC47BLEJFOIYZBXSyyNCZc+DebWixTuYLMErauVzNC+/ahMNDWj/9o6iiJiqP1QHnxPf/7t0zVA
NBNy+C4KkfUydusKzUtqbbPMAhaMfFuMuTuqz7ggGvAgH8EAS9ziNX1JsD8dJjRPYDSM+OrgjwK/
bK8P3en4xymRJvJdrwEuBQIpOp4KIQl5IrC8m51SSnw2fBnBWj8cbCXspzaBvp2sP3IqTdALBFIm
yE71jwHbIgA2TKk6aG95jgKf8H4/96y00qWWS83uo9xmoRrp9EK8pJ7+jlZ6CyXmZuWZut9fQ/qe
0+pspxIVgaOi3FpCvSrR93s1/buga8YuF48AAwA1nU+a/YyfMhVXrkcXFmV/UiUUwP9R460dfs5C
fL2xFvqn4W8jMVsRnXaPeTpu3+HabJoIfmC+pTZ8A2okQ/8AYmUKTVFGZWGQHv+FzTXyojhpWRxN
D7zvPJjDVapoYI3TVohBaTxOMJWn5+F3peDfa7wimlKdJ8+yirhRVOOJ2Dmjo6PfpMcud12aUDf1
mIIne8dssDnN+Lc8jQpOEybO+lu+5x58SWocPAN3IgBt6DSoiZKm6sPtMLin609xsbIRVM7VMds9
KvpbjEYZ+yPWhsrOkO/FsJZ/DDn82p/giry1IWQ7EhmVqL3lXSTJluLMFwrzef6o/qcHKJniDsIv
OpqiD01roYwTXpD0D+Ku0JRuGmeT2UcC0wyRNYL+B1NAMRrtalol3JCaF+FhzvBC69/jb994gKyA
OIkgbUMfGT3UPGZi7qvW/a43avF5Dw6FAq46JY74TQM/0+gjXmc87R0F54vKcoMN6IFPLfyiDwEB
mPDwtHVZt0RUfiSBx0YFWKqUio4UiC71XjGfNWzK/ZsXj7nxXU9KqvZWTqWC8aE9y9P+03ap/8FF
F+h1u97+sLmwqoQMyvIpuYNKTB5bToNmWPx1iDvJdOTcb2UWV0NKigtYv+MfYZ6nOVbGBn+2jkS8
JYTxye92cMdn7kGqf6unIR4GTq/9IR1rcyMzU0GFi+8rbFT0da20e1WyUim2p/4LONyLAKbM2+S4
gq47DWkC4JLKTEC8mwpmmQHRy18iYDQzUmunQ4eTWnn0goba27sD31mww0oc7gNGXQAZVWVsRQdQ
MYQ21AKzKgG9KuG5SlxhxCLyBTsFVZpdvqC7mXDkdxQB/BF5QQKTzQK08/bqlxx3DFf9x92M+Wgm
GNLdTAucTRO8bR4DBdjBf3SQzZnp87LvO9hKESpLIT0YpDTIzqfl9fSTqclqsyGdXBEBcwSzmZP3
Fwvw7mPAg69UFF68/xOA/hKaf9h/IXTEUKPxzjNsT+DplR7MVD0VBW1QE65Otmq60I/cT3U5rcmb
h+ni7zDzB6EW16b69Wr/q49OmecA5c4zFTyCMF64k8kH+DHf8tmFASKsnIu4L66WDSQ8+dbcvo70
LGUiLRL9rGYBwu+8mOtVUv/VhqAq/rl4nZ/+OFQPzqaBzsQ5ykspapsS6vh3+6uWz895i1KdkNxf
fBYpzGnqPTw3yl/Eq7kfV7T2c4bVnUOUGGWwlgpvl8JaJ5bjn5eg3AcZ8n5ZLp9dWDcDVI7s5yGX
yaCAByu38xs2+TZW7e3DLoKKOztF85cfGK+ZSRvN8iB12AJrfN6/d6ak7V4vQPrJdiYTx5zasr0h
ag7UwQyKTft0r4xhWyZbUsZ7hUMmgDuR6pEvNkqKWil//ndISnpn1BTC67KTpHddIfNGPchjhAEe
TRSuu3sJIShCk1sfZrjfSNVWVFouJbYEGFOgZI4QnLX+0FPbqWsRPeHfSB8SPUVaN1vKbdbvESX7
7zfGIjfnJKhSw5F4FDFzUrlptn2M4DUy841P5Wp1f83Bp3Mf9dEAhz/ix+50kO8uTwnvj54pGyDy
BUiwntM7tbuhc/7kvNQSl/791FUTK9EPZoDnnKnnMNu7/Uh/DkyaEJCxbwQL2bMUnWMj8IGlrh0e
Xmduno6j4RqmizfH/tsz7YI3p5lFcoKIzhyIW/ZJIP30YsLASKb3EUj6Y7+gD3boGYbldkz6Dj8y
dj6zpgKiEPAwZPWKIPiVuqxuopdEoeUiejVTARzoYjgVZ6lM5ysppD704ZgRdbYYcu7Z3NAHGr8t
dDfTpN/UHNgv1zWw7uuwB5OU22pbpOHq5/VST+P6WjU/pmTSt4yDQKz95TcCA4vwP2q+UozJ7ok6
yTR8hc7cqh2DJZgaxSI817TJP7stFOHHaIwu21faQKnPRrMZ9IiX78B1RJ6MWsFKSbqniCwp5LP8
IBOnAGoQEjKVrAU4kSA7dFYOmSsMFy1ah4pr8LAIn+HdLvAiA+KET1kFJ8hRhcoZM3uDzlABlAqV
FHgkXI5XABk5zmPm7jOL/7YwtCqqEZEKle1a87Liz3zS9drBvgm0tdBI/aFH04pNrqoT/yKTl372
30FLZbsmX615YQ5qi/3OfOBPEwNrLuj4jeGNAVNv0tj+WXirQTsOLImmHVy0ciesDU+5dbMLigI9
khAjHk9sKdqfO+uAZYRtx7bOYCqMubp+J3UnFKLnCldZbtorigxzoPEcErFvEwSUIhff+ZvZlvDT
Yw9xKiiUqn7t05U3sx8tnBIdPLsLvdE3bXGmDTkun23rpI4MUsDkk2tbOwcdGXdfXGC+f5mbjhu4
SLxbOZtLQNy5oIzwH61iIIoh0qUK00R970JGW7t5hVGPu2kMlyTHulyMmRnlH2E9vKh0fd8zlldM
GOFJYzTZDfiHtJWyKJ6qAvxTqYDU2EVYhOSSB0VD9vZdNmfTyGgK4SMeth991Lw+UlkYtVwZ3sS3
96TvpN3AJIZ4L7HoV0LbPKL0UptNkaTMQjMpx3HYKFQ+NZJQN2/8iCTqYl3TyE8DJiLBZysHKNQW
couWpsyR3J89mZ+Sk/drLvZbyA4+gR/dE17vzNZ6zdnHwC9XigrCWEZE8KBCntpScNsWWv5XMqns
PiPvcwOfDxWwVPZNuFZJqwThgVKtMT5sUHCEqaHbwQwcrWlWiLuLogGAxYDYjcjrpGao4qcXc9xe
UNtjxOFrJhlyXnzZSXPDTsWuAYq4grfefp2MK3YnFKswPdQWqF3KfWM/JgQ39Uo/KmlQAmt/Zmu6
qzyerdjFSB2UGIz6r15+6bJLwnpaD4NZjqf4tEFgLIoAWDIo7d/I92VT2QfuDSd7zKEn3g66lNA5
DgdwaWOeOzZHs/As0zKb7d66wO/UBWNUW+jZpirPUEsfEbs71B7bhYprb0YD4dbiWm1xpeEGgYby
Z8gYdDGa0ae9oERcvEvC4bB5mF01d043nzeDH8uR7n9rZ6COPM2bSyxB7Vt2ffCcWEISMTRbijBU
ciHVtHOWJkgUZhsPuoKHTtFNNhvP5kyszClDoso4zqWUTN66F08zcqAWGCvW//VhPOGYVbONs9jK
he/EyxYHwvITILs0nWiE5KtuvfRJkwg5t22QmXq9y/ekfPGQ7SpnbwoQSp+x527/hUCABm8B+2Ya
qMFR0tQFtB8TcIavzmQTPQRxIiiFqAxT2S1goUjUpdgG8HcV8shjEpXEY5pn/mB/TY2V1rBhINCa
guNx+vqCnp29Zk1pc67yLKApNdfiPgwlnTxODUONqeNYA/yLdEi4e5cOVScq98XXMjn0Vx3HEFQz
QoJ4Aayuj0ey8jlsp+cHTUUI6wM6prPNCjrQKsAwSjrp+TzQmBkVc23npuxtPoRGNYF6SMK2xe7E
8l873DnCZ0WqIxbAsZhX8kbFh1a86exaihwJym8m83ZJkdNCUB+lNGMeTvOTaxNE0wkqP+sCPOsU
vAhkGiUUHsYXBPtFb9b5LU+ErRjykvJ2TXwjHJLjcZOX2ho4qz5pR6AfC8xB2yzSaH2ezwAeQyQA
L7sXG+3tIH57OUr5KcloNB2RRp//2eEqyg8kFCkAD4W3F6lrATZVt6ASUQtd1tgRHzYHU6uTLOHa
kRq8xM223ARDZtY+y08QiRDbI7jaW9frV7hM1s6F78aTClU+0vLbLpndH7J5J99XoMIPHdATN1bz
ZaX9gDjHKiXX1RvWQ8WLgOPm5X7F77Pm3ueJoaoICgIvYpv5YBVtC6Ozjt2m+GMX7LSZn+RoGWEy
QP8JnqSROhvRASiyWmj4rH6u6VzMewjt8Dxpj6Kjjv/AX6UlnILGpLsAQMYTEORYlcwVR+X+r+FE
jzzVRdcWaRII9R59XkdwqzoimnhD8EaVUyhQxeczl+AqlpvrY8wJnzlhzK7TORYTQ0ES68cRmlRn
GMfavKW2e3fTdhuO95mDHCaCmNOH2Xp2TXg2JytdXGgZ/1Z3MBXdDsdqzcTA4OPgEQGbILPSrtkx
aK8ZkUJYF4qixzQ5M4MJnWGT6uRXiEfgwEDFNeRLsGkI0ymLCt8I1zxT8SjpE/h68T6/gg4QRz2K
R+I2KA/UtfKtj3vuRGCp6gcuoc20SK2nOrE4VRQFj5nKoR5C8TeMZrEeDmLReeSwCtPTQguTLz3T
nE9gUIi3YKPTlExUhfITzPwfO1QCoFuP4bx5SzKWidXbFg9IKDjwq8HrUWTCPdptkHeib6WT4+bB
0UjKqudCUcsjKD3mrtHKcEAWkOgpxoCG0XCB64ZgKmvOkp/kh2heHY24HatNQsvRJ18QQlCvip70
UWNYMP1ptRcqhwmoA8LI8EgpOtv9jLtYcelao6dtjPcNx7o4rPR6QJPL8L1UphWr5u/Vomk2OgQ9
xe63g6FW8PDXVNCVpkaXEdWc+xLtJTDmU5poggJ3CkGn6EYtXPtUh6AtTewS8nODUlkJx1Lsg3FY
6TBiYMMFXNkJ1w5qwK9RVfSfkmLU4RwmuSICAGdwyj0tYpqQKfbJDfbpylyzclORpX3VpjQk5CrV
mcPYdH91qtZRencb3g/4fLKLb4AcPU0Zo/d16O4Se28f67nic+82advqwSU5mj9b2Z5/RJoSbZbf
lIx9BuXP8YRseWyY3Szi9dMkMgCnkTKHyVkS0xHBZX/dpTeVY/VDqgf9/1orhjR1ym2TCdmn6q7f
Tvb4WVEj8fw3Aa2Ev2wn3tXjCNIFW/WVjfwOM2tWMkVQQM5u3qy2x+ND1+jmlrEXO8n6Abk/WbpI
Km9HkdmARpUCqCyPkk02OK0qmmqqb1GvAvYSHGiutP+YxPQQPF2jUMVbgu2QQYYSmUdpsKMX13r1
rwrY5jqT9TlZeDPPtIo3uKMaXl4nuzzKHy3Px8AwbXj0BExcmEqJ1EUsgqKyuPZwZqKBnPqbJtH3
tr1VKoXs4ilQgkLx8vtotiHwuOkzc32eIdZk0BbAPAGhhivqZcWWjehaRFPSVsXxbHekQRuqQSxY
mDL7ipt8V7URqAkpb+Mp5UGPFGBL3INc8G98yshAKEUcPQc7Fwcr+Iivoz2yDmbWkn4WgmgYE53s
aSpp87DTROMyJjYpBs9mebiVYd2MxBAUO6RkG+myi964bmULooLdQTJ7v1UrQZcMyBCo7yjheSQp
BPLf82d0bvUaOLaWQigrn1NalRVhS61Cnw2wiDhKzLzVw0Lq8M4Ctml/hDs1CeA4XaEtyIs6KJcX
2h6BETkU+7V2aDSKYu7WiT07myRrxmB3VPNcPysLWr8vOtexuGjfrFRmBVlJyqm9YoLl8A2SBfOl
53klGLsA3A4cDqS4SFcUoAY9wjWeF0JwfZuOq1Gcm1uo6Ys6R9CTDLZb4yaK8yeZpBpDDLNm8Cms
MLb8NhT6LyR2JLcFdOhXKaMILitWrHABGWmss2inzzvG2eEJlP0iHqLMbpwhLapgWxdtU1KW+fXE
iBKRVUxPuTDcIV+kBh2GunZF6ocJNtNvLxS3SQZzXpib5U0heZjE4Jc21rXByBkfEAAfovRL0ZIc
uyVG3p8hqJJKsp4vZVJJPrpVDYcZEvLWMNi+RDu1Kaem1F9hvYQzGgGtnZmE/UycGZBROzQhxABt
pttEevyyaeEuDweeCa1Ka0c5EBKjYIZ5UHl1HP4m3Ym19MpHMq0/gp88sBegbZD3oMCRPOwJ7otD
5ykAlJ1s1Imb0dfX7z+KmHoRcPI7Sq2UxV5UMd/5hNp8jWMYUPDY6kPMur7gE08Eu690tTCFpXIQ
7zzWY/jg1IuUj/l9mlkg0Mhw+goOF/LWRClLPVLjnvZ1owXgeQ9z6DNtlpbZRQtpQ/5H6PnU04Ic
6YweHKMA7NeYi1CKkPw2lMBg3UylSAFp55AXh+XzV/vbDsH6Hbylphugmp2CVSgPQjOu/cfmhpeH
MJ30xjgnAApR7jsqQ6xkmMWicGYQc57R0wO/Qf0i03p1MR/XimxnubucfjSWjMVR2PGZ2JXEq15f
WrIVAjExz8Zt1D43L/E0+Smuq5/sYMU1+6YcEmlh1LbYDQ1K8NdDTUgVsnqmgRWyYgjaaVY4FJNK
mfr6NR8TfEPNS3PtXM76Z/xy46/bxjzb7uqxIEqLbbJqG0pMYpm/HJMsjzSIQmofJVZ05GNGqbtd
HbDH/f+1b/xh+hYj50ieBzZPXYy3c+mIzDYjaaVAKR0quHqyqJGYHxg5fFrZrS1BOdKrSeZywgSs
SlDKvOeqq/Z57g7fHSZv/rvXdOx/6G15VgW5tsQ22p+LAJQRBuTUCMfSbCs0GROMtP3rBCrJmX8d
vnulOFt1nff79xVtJZYzLmmDXS/DXW6zQ24PrZY/73N/4j/W9z78An1YtAq5u5mk8spDNKPi5hUC
ONEV4NAx91RP9wHo7cz07rTNvdHeaOmcQzW/E0yUk8hGh670E3eCAqWxB0CP3Minf00QiHH5ngXO
krjUWytD24cGxnQ2GhuLAj9kH1LaocZbeX92bog1PhGhfnXOmw6mM9IjQPlo7cflXteNFq5fWPUt
4rV6/37H6ZJV0mAAqs2vdWJPiZUppFy0hDzSIDk8T2GmYG/FxG1CQRICib4nhwVQtQllOItp7IPA
/9/KK96TMd+TDoH3AJ4BbgIbfvisbPp/xvXVjnVQZ01rzNbKhGlJBBGXhsMO6Hy93LsulElki2uT
xcgochvQQ8Gn5UMuHN651hErwYxZ2s4Z+D0VW+wcYl/F3phlCc9BVEfb49mjm3RJpsQJrpd9HSzx
z0qMhXX6Kt5QwarpNx9tCrN9vbGu3o0+E0JR+TxW36Fml7E35rD2rbZm93ET0rjFMKMIAs3K/yPD
FXP7Koeg7zUub+rO7jWqYBmXfHE0Sn/SUV9WrKpni11tPPMCK7L04ADS4vt4+BFud2b88AELlEug
JlAD4FO1ARoOyKbt0E+IDQHTj9mW4/FOkR/1qCYQSBZR1trq06qA9oH+3IvFkU6z7IB2cNLuUTtU
NUN/Nc9f5vKYP/jgimzWHclbezn1ipGDZaknPz8ZXMvNbHiKgs5/LgRJwHKY/S6CqKiWn3FMQCpn
9SOg8C/hUcdgIyX+vrntFGTVxazWLtkdMQBr+TfSq98cAprRzbuYXGSbOaE733BHsia5RIKv9KUE
Qvtzx9+ABP9SfE/Y1a9bA02hGq3own3ck1KcSAQUGVve7cMCs/NAXKb1rPGbZuTdxD0Ml5Q12He1
ZUFQflnPwpP5P5VGH8nPDgzc7TwaEn/ln2wENJ4Yz01JS6Oba9+2RnupQMFMCE0ozbw+YVQLm6XL
4/LT4dNbQX+A6Q03ut3w0BJ6U8rjzNLtQmgu3954M05SZl5mk1sxcu1Oogw4vDptUQwexutjM1ia
pkfMaJIaanrXMeLtG6cnKnJZZsUIUwp1z3gbzl+b1vKRsMwWm54czVDXAB5NZDrqt4qHeEnicHcx
WQ+Eru/E4dUMXNFtpWRK2N9DgntMuQaLq7y9EDH/vCmDnEWGd7sgKjMrX5vCjL95cuXbhS3Pdq0/
k3uBbzZ26pRtjcbuvzzEEs1ABgitBr6s2eyHgMfikQhb2r68jAfbSP7j9ZYL5cDTDAmbmkcM7pv0
56sprZUZlQ2seEn/wb6ypI6DpQ3TLXADUobPdASLQd5vExetOXo9D7juE8bHGkl/psajspBJ6oMU
zXJ7MR/jqWn//uAxKwqk6I+LhcGRSgZOwArBVN5yEdtjfVet5TK/OkhdlQ6MKB+hPRIt4fwkY5JD
i5sg71vnvq/w+RsOkil0fGJITcbbpEBWVJ4kDGBwR52YqEKKqTn4zBAIIkS664j2ELLJSOU2V7Zv
fI0/jEF0HfJ2x8+xN7cWtQmP4xa9lzi3E/54Jpn5prZuiIIQ3OhyYkTNcvyabfuBcrlfHog2LWHX
lMs7/cY/jmAzXsFKxRnF+GWF55r66Sn//0YxwZTmPpfHR6DQ+xoTZdR/Fpmbldb/fWEg/jgJKrB5
YZXH3qgYCNEMxUn/ZIVbEG7lK63OqdSkqiT3wqLXtfCdMZgiSmktsB9UZ3dRv6pzjMbAEV8lhweF
A9wXccKercTdDA8sQ/K579afB/WAZFX4Ir9kzO/658Bbdr76JV7BieeqzdZx/cA2W7kUgbneI8HV
nui/f+iQVeVks0cKL7GAIQTYJdYiqjEwjxHM8Xtc8Fvi2uaLu21MDpvCBvxs5hkFOvdSM6xd6AX7
sfOrMHLkpyfwqPluprO02cwEZD59P7SXrp4RsnQJZ5z/3SLt9i61l+sNqG1OqmrtgyWj1ZT790sG
cdov6zlAmi5waOTfR3cVTv2fI0NNpVRjj8Wk/1qvc5fkfaS0X5R+vQVcV9M7hTvXyc/VAMy2/Jld
dNfmOkFcXFnINv4PUJhRXXWjZctKGOdoUiztG4srytF9CMXB57uW8QJ9hhfUXMlRvIOE06Z3IAB/
3+K1w/GOyhmUwy7s9TPMiJF6u8hPRqiWylBxoj+0FDTOgBjswgJr6bhDGMclS1dePzKPlWK0Hfl2
nN4sxUuIYI8kLRcgBvvMARBa4VQTGu8uvmhH/72WwnrjyyJYYLubp5gwvber/nCQyRG5U08ceqWP
V2mmz7tUAoLVtNW8upDj4p8xpAkQMVEd2DtSs7tNJEo+vJLpHBrlrIJjIK6etAQ6GhbwRLufmdA1
is1u9CWfbyObvxiSvMs4n94EXCLqrsexCkHrCx1ztnfs9mfylkqO/o2R3G9TN9k3GADcAM9XJjyM
0xEXERXPbpwigdOljdAeLaKMgkn5tqqpmxxs6J6/bUQ8c83+XEs+9fJ5Sj59t+L2fmA646JUda04
7F4P8sCPSm7NEhvEdtlnImafcqPDb26Y27AYMXT0019LVILa6GChefmefIoqdEJuVeDIlNaTcNh5
panInFzONPyksKSzo80Cp/DHGoLXnAWxdLVsc0ukw1CRT9vr7QamiDndeOOtxShdQ1c+eFtZcYO4
N1CofaTIm0vS4EnEyKaog5rqhc8VT5LUg1YGVDs5yO21oLuw4t7rsbZvGaRt2M8vk5mMbBNqq3Z4
Phw39JJIkKfDjcpVROzh33ZqoPhmKezFJakBggDRiXqLew/gVUed6L7/VnyzJYRAOij8ikjofuAj
Zdg/RwYe1eR/9qjag270/QmD5nRYzSfPfUZ1Sj3O8g+3+DExgsKULRWkaR22iPPcR9eQDmHj4KCk
uaLppKXDnuEOzNcXTK9gdHMGbMCRt0df+00iF5EierD7k2nYb2z59OZgtRgUR9QRbz7UNm+HHbfX
8ut426y+H48AyPLwu2Dkb4wFWI8PVfzQHCkO4MyIyedvtlPYLmOa92N1JnPzPGWp1mBcqkfBDJ4Q
SdLuBFfzXk3PY1Udclos5E3nRG0lgpY3QMQxPTk84u8mIrDnl19gpeaZFcGj57yWWMZgxCZd/zRl
FNZGtsx/YsysI88ZZNDEajLA++LWlIe5fugW+19+IEnb5ryYmQcNZ4CGRpNMu4oN3RVX7cmSepeP
ES0shRAwhJb8lzNN4VlmOfp8BLutUtSOB6LousMe5UKCDfdHb/tGxG1VEM9JVaS8ENWH8EqIxjeY
M7XYn0Q+AUUqNkyvBS/gB3ulwAnykXleldyi48ArV0MmTiqxQZLzI+IwvFNbfGE/n9TSXJb+82k/
HMaQVCm0gBq/1d3XN0LHlz0nPsIgd77+Fj8F/b7HSx3FMFIelWx0Lgx6FQfqJUnBN4GtV7p2f0KI
XQq1QvDafjeYnlfp7r/u7011Adrq7PRnF80lCDaemAF0+1/U7tuLa6yiT0uQ8ti/neRTvyHi7u8A
d2Yh7plWC2y6w9Zkx/DxJPUkjSY0FBVnyHxfd/iGmpChKtahFtNixeXwnw8oJMElsli7rxUA7G1M
BZdFQI9xykL1l3KnH6q1Wkln8WY2AxXpAakh3/fVAMZWgtIvJ1iEAxldJVqkXacRp90uXDypmesX
/kbelVtm5z5+WWUgmvhkIVfobr5+dxjs5sstBr/2k2RSBsRdW8SuHGrLP4G/gHx+lw8FsJQNKUPZ
4uIiNdIhs3isuljek82VOvsyc+lrLcrS+5+oUC4kgWu0NrVtTby9vryBhUMWWXm2pJry34n0eVvi
OPfYZ2pybaidcBAyHog35EgY3zV3Wkkr2ViZREZb7gVz9+HMtB0LC56vmiFpu96nQCfvEbuv0EtZ
oaLJVzCj3BFWtPNX9VeVUVndfJ+Kvk6e6j3n4HbopwX+szDBRr9zeu28hzb8nfYGLuG0ltmnOX2y
VPlAi9/o4BkWxCRyXIyzRJ6+1Fn/dMg6D+K1zFVDjpHOhKPg7QG/M+/fbWSfwek4JwD77q2HT4+/
6gE3a3EfD83ANUz1tfcyei5jQ2BpSjgoursij29VT3a5gI4f4PRjmesUHxYZDuoXyQTgGjhvUr2s
d6jgxnkUq1EhzUcn1V8DqF6wHta4PPDfLGxmda0HukB9Ww/AmdET7qxGpTLtr4t+eEi0E+qeEhkn
JZFBQRXNzZ9qb0kLr6pGKoKY4K7u/UQorLkDlqf9EOdHU2X5hW+POkkCbIwLKj0WfyxRuI/SbSSK
oFWBKjWJpsycuIJJhkOy2vRCgLLuAGaXVhAOWTk+w3TuaD5vIn9XrTkAnEAERQd3GAbNAMwzLVfe
T1NhJdKp5XWYxqH474UjnbK1l3A5FgCfxch6/U9xLPWl0UOSpIHy5K2ckjgh6fhi0XWhSeXr+qR5
PAZG3I1Ej6w68bDe6xBk0s6WJmPaU30Sv7s/eLANtCK1lMsLIb4C0vg8GWdOI6tzBHyCzz3uDjzR
iEN0in/4Z7Pq8fsp/SckYmH2jpCs47D7MkvQ/df0KGT/z/nMSBaIHv7L4aHy8MlWZAUEdDb8BwY7
RZPyDnIpu14FuVbhK686lmgn7RV4fXK8FzswupyRShDUFYEWLHQow5Y/im2waVLKuPeLXc5PzEdj
1qENdtutPZ5/cEVEV30iYAQrVOOnT6/WTq2QV/3GoMEjqmDytEG8125piLBi6Oe79FqPbQ+51CAB
kzeVwRnOUmrhFxkHSEngz0IRpRgPqP9BoqgWQX1Cwl7BmCG4LMP4k5zPxG3uQO4lqU1073JIVGb6
clRw/Mbwrw5pXm5kxJNvNakht79E3/npYDD8K8kfSH90SjrrF8oKqCTLnWb+IACtZmuAmpmmTitW
5quUpEg/GCKp3QbsJyc8YeBCCeRry90qFQe0f3YV9zDW94qjLlrVwjczJd60JCRu149QEUi0KglO
G2dH21HVbP4I+KyDGskh23f0IvNrVyksY2aZd6YAEFVfGcRk+Cq1dKcyDURTyqXZ5JJ26avB508W
4aVTfp4KeFY/+BRL6//+lEuBEpNf3LWqeoA4uOwOk8M2lTqHnIWwesCXwVIjROVwlspkN8sitMrp
h/SuqC2bh2afYtxIK3hjQmz3bND+IsaxSZPMz+lb4tQiuyiZ122Vvms/yNKnEwP/e1KuAsX5vWlu
SDfNoI0eH2eFJebHxEIL6S+Y5qC2FFgOy5xLfOKhYNcxYtvxd+pbDIJxGnt9udPlrT5bLi1DVy5t
FXcPmY1xve0+E9HcfHW3Ont85cx6OYSR3MMCBON7XTvcgfuw1E0Tl/VJkA4U26bonCidv6y84CWY
vDsdboVjLSsMxaO8q5q7h33EGJuOqXJqwxUanZ+Q16hjXhWSpCT90O07ILIzpdOqly2607O28So+
Q2NEQx/l3zZrv4EGbiuhbA4sU7xmMTcIVVNuSuiskSvKnLO3ipvC4LSclaFMYn4lT+DokXNQSGlV
P0R9nJ1bnmweEzCKQxGG+eHrStvItMQUHxcPFjF5/D85qVh7lwa4kpH9CxhTwK8OLGcununc2zQK
kIDTyK4fWi06tTdkzw20WwwDqsmYc/U/c+VlAy81Bq3L/vHhmtmTAtDiI8ct+YxpwQZ09RxI3wrK
voHiVpYGSW9LReu/klfugmI0i7EcPd4JpZoBoyEX7I+rJnY4HcLFx3lEGo7D32yxAC7bJdrWveAF
bKrXowelJimS1i0lEkrndAHu3qk/Xkxd/1HA2EfryMIPa2aeIWLwEASpIF4axR4em+DhcQdvM49c
PQRDmHu0noKqU8smd1bwp9AlnITXwzvtRbDR3hloIPEGykTe/VNoLAVkFGQMvVfTGhNSnXOd7Oj9
EPpiHgXEsGeZsKau0EbSiq/Vby4PKupfqep/hdMRsDI048iyWWpUyTKGum+0X/0D/0kNt27kFKXR
lS3kIOXJTb4HbIWLhlyqzSlpzPatz6v1I3ljOgttIsBSCYWRhJ8IfFPm1bIjHIf4sdqJgOzsd5eH
kvQevn7DfbT0UFK5GSPOqjLZ7GPUTHzYJXw905JIbf4c18ogv9NaSEjEzxNmQbdnmfDGqJ28tQq/
cDj2YBMhpo3bGbPsEhe9V0m9InLJSdNgvdjUwM0YbJWG09Z4KFUJ5gAxsrHMNaWiBK9/llKXGbwK
eRM0ZIQCcFAHNcuFLsM2gWy5iwX5Jph/nA4FVxxz2NWHwQFd3XFPsTeC7VUlccOvqmlOEhjRNc3w
YK6sqyK5Fl+tJA97yuwzGuaNMp4cTwCgfuG1cDiha0hVJV/SlxR9uhXxIR9evugWkXGGpNeSq6Ax
oFVSpPtTUoS2XF+MfiLCam5GKWt8ohV1Pw9E/kUIcIgiwCy+vb5gcTyVKY8Q6aZTHQJtkfrhAXaM
vFKPl9JJSQQr08tf0XIuYwcP+iLcSvswvPCJZtp4ghUGvVW+pDvLmP1gxTaKQRUHM+TpvNbC4OBm
1P3NoJ+8K3ptR/uPwoqo1GndYe9E0deU9isXo/HmA9PO5pE5oJz0sTx6EhvDcGIDCK3SwsbVPUR+
jDPmDGt2lgZNwxsB7GZsnFSjaCWm6ovOX8yo24mjL3Sahp73l8JzZuwn9bi0hsehTGJLb2ctH1Jk
jP2lYtkvhpqFkVKJOq5Rpp0Odk8vVuJoWZ+e5Vk9RQ/rLno4GasIGDfuN8ph+JunSljx2PkrtSNo
AHSIgYQg5mO4dcsnOM233WvPFyGGxkJldDYxqK4w8RaENe3EKGxfmb+gZqt3vEntHb3ntGTdrV7W
xti8+yHphcIzGmhtUD1fA3pWCti+vRDvHxNJp5GzhfGcJNYEvcjDLx/IAhaWA1avggpvDdLq73cy
hFe5yG+qgrHmgdXXfxvpHLgbAGe6st8/8Te3qk7JwORh7nj4fcJhrJo512oqeZ62KRyHpK7JBFcB
bP5bd2VbEYECDeZAg3JzREdHVkVmhGBgCc+szSBSrgD6Dc5xfNzAOshTE1E7gVQR4IQaaVFdVyO/
4z2yDq8ZIkK6wwCB5VwEPOPYi/Lx/8lGOLN/n5ML1lTPY4S5xY3o5OUr2OyFCL4BLTRtGAvO/RdJ
y3MdaJ/TM3ttS5gcYYv0x/jhjaJtUhBV3Q7/Q8I6eHeDvLSduR6iOXlZWsKwGWXqzH6FrZKOkaWY
fUu9IoKkMfSb970G8q/aTQLminiQIG4S2a7OXzFLqeJGqa+uT8R/wT1XXvPoQ1S6a0LwtAzpi4Ms
lujB0MWO2hHHOqEnihs7N0S5ierE7wbzcwy9PQOSqHejP7dD/rhD2e4T0lp38F3bsniJdVxMo7/Z
Bq8igaDSwRKpcKX/EekhIKfzeU4WIilhzxTdrVIaPH3TRwvwORaQUp+BSb0BOFwWIXjlGrmPoeI9
pZ8Tda4st253GmzSzQvB5JL26Chp2z9HN2YdO6CVhYhj/Sp9FN6vh4NItejPh6wvTaj2FgVH1Zyf
fhU1AXzX6ysktMgM4uY2dc9qShJOGvOwwamApSQ7fCgTjiQ3m0uyrRa0Tebhj3kl332bJwrMqHcG
BO+floLZrG7MegZeS4TQTXHqpGPyt0MSnAl9+C0apuCSlaQlnkU3jbsO6EgDPjxGdy+gRGian4IV
8qnYXMYRannNWn+D7lXDOQLEeSCZqm5qbVTR3yk7UVfiA6ki3LwIQljwKzY6p+iqa/SjcqQtTs2T
5DwJe1iNCgW7XEJVXi5DIpS1Mq9QwMlMFbXBpfdqWZEqNWpVs8SRQosFPhWJiDOq7v6OBDH818ub
gkRTsII4E4qPY+5Wf7muW3CwYzGPHrtEXntXqwxG4ZKN2RYSQw6R4TbFBRnO+NSThJNyJ2zc2CU4
t0JdC8lG3czRp3b4hXBASt/CC3VJcyOHCH/XqwaMk5ufKV4vHFEMhc9XE/1JQMfnYRfmzBCNPrSP
+CNk5ofnaA0eNkI0UkAR28xoJHSDXckHQMp+33oy8wzWTSqChYgHwTXRwqJnKbmpZLx51n+ILCoI
l7NtXKTf2olzV2ioISdQc+ThYJS8NBePhHeyB4DKwyFxOuUnr5ZwmyM8PAT0HRnaHnUYfUBxwGqv
ILVbFTaJTPZtFvWvf2XUyk7TB/JpvGc7PNuyzWtPUT6zYqcC42zVta67dTUMT2vuLRHOCKVrfV9d
5DQef7McSmwXkQcpJuzfCqVi6WFnQ0aO2myRMeqPLH9HCMZeSRgada3WEGQnJhHChV9ZkoSgWCfQ
EOS1Q4OScX2PCKTuhxkLnA7bnxJs06D9ZTyrEO4QJdnoTxsT9F7NSc4z3YGZ3PJdo+CRl1UIuaqU
m08DphJd/Glyq2BywxFzmadPKOxmDje/3tRPUqdqEs+ezvA3UZuU3fuxjHIIdoeZCcHrAjcK7bcC
WfP6OGtZYiwcYV1xBYZ70VLF4lbfFSsq1igoVcK5XiXj9wPduMrW2lhRaF+qyaqY3DeQGerxYvhV
4+fU27x98+uspTaKwB7KLyRnT1cyUYykzPKnhiT0D31pfH8jJjczLt/+CzHmcIXGyq23JJ09yH22
EFm5JsvhRJmMOhAT+IuBwGlvGhMcIuUr7AVLKLEcItDymNQ3xCuQgM0Jd9MTzdKE0i7b91mqkCpy
kbYxjJBbNESqMBbe7LiC7HrctSED+IAw2js6DF/zyq1G1JfSBvJG+WfzTpc0M7laJjqHxhEKFski
5FhAgweKbejZTOWjGoePs6znN+8Qmf71YISGaaYPYmPMn0HUuOTS+2qK6flyXsbhMKi1kbszoouR
HcEKbhKMLnLfY6lMta3zkeXyH0rUDS/th5Rj5B2H9LjdgSlaUSfZ9z/H/4dCmfNxBqQC7SZxioGJ
gJY9NW60pV4vGxvv+q/FbXujERzw9jgAjOSXTxILIH05+vKCZY53koy47WgADQYeOKyg1tW1+zSs
u/o7KTKBUF4ovELr3GeoxlkhBf4/RxOZZl31Sp00m84PQz+qAaLWXAwMcuflMc81rsmYMpNP3k3U
HECTJGv/QTcle6ZQHpERC8dWV3NX8AbC/MdQrVe47lyU7SV5egzdrRZZghWtDKBZ90LL+DXDzfRJ
U8vLjatT9EgtYTKGblI8gI66avjp7pl3Bi4/7907I9wJCUse1CoGRXU8bbSgND6WZXGxZyAeM4Sa
L2wWjWJPr4sxXipV/7GrEcq4mWIASccNAuS1gowxH+2eSzfX3J5ovDKpBFJyZuaSqs6AzV1ROZhJ
oPO1aqeMFscC2s/jPMe/mTSEQQ25wTldICqmF0ApbXvniO42vuib/O7p+dE25udAoaxu5teralOi
ihwYhXkHWc5yeXPWBfpNyZ0ku5J9q4o/V+RpBfokjlDinov7qN7NlfyQ2AJQAscHgOWYsJdlweT/
EvnZzhZx6C6YlB2Y4nAN4G02ShBrYQUC6HUopodY39seb4pdl4BQYzqFQesn+SEib8DLwWACN6gJ
nF24JHjYkt2feS/qN2644GXsTOWytZltUqCTgIGr/Up9OmENiLikvmrqrrHaiGPq0lqEr6XTTQXQ
bbljBcI70ZSqxmIChVlzyQ/hfjqCGrz7FeVwmoTzb2vv+9CkjlJctNVYAUkmTlQowVrrPgZK98Pt
Rtuk1BU+l+SsG1wD843gNzoroQ8VXK1vAL3znwkOH1BGRaPfvzci0gqGAY2rfcK6JlaX052kZk1q
kBAHVBgLSqDkaorcojpFWs18CYCTcpUaQeyj3/mpzn3oemSmBbbPZu+IB7e9vpcV5mqNvw3Da9f4
qlCG5dx3zqFbYhscWwxhr414ws90EayiVrR5VAGcbD01xlSRIjwzCICXB/FWZHHJ48fQAQUGF+D/
F3pEIRQB82/MmrAjVvz7KWqSztQrgHxWo2r7FzO6Ymo6diEBODBF9sOKK8z243Q0g2lQmqN75BwM
nsnsvblsnXpelhSuzz5zHLz+Gh3GlSc/cY4JalYEiFBKG98oYF3CkXa+CrUp0asVSPHmsUEQDSAE
bDPut+A/OrzUzLM0vVo+T01L3sUI18FrRPb2qGUMRMvy204rg02iJJVKf7KiirKVaa4rdjbOcmPf
iQF+nQU9x450CAkmtUs6HOZqxmbzEQYa/49uKM9YWGaePEhGaSS8WR6qANA37qytD42MEzOO5M3y
QevNDuAbMVSNteLJcUXADN6LEX062PmsLNlWVEpgwVri5Hu13fxzpniTGJbl+60JyF3rsUpmy5GL
2E+jbAj4spRIY1t+Lzqe1/HydYq6pXkbfnDseatfk39JQdUnCALbYJGZDjdtBoh9RpJABaAem5oR
HzERiFRSSfu15tfK8kQGG0Cn9Mlh8pT3WRlSsbTl36MC7UGN/l9lZDrU17Ba26ZshcFp3VBWlUbu
/JQmlj9hf+qmsBOHBxo9Xg2a3QOdd8+COVXdFZpTFi9KxDm+VbVY5cW+sbTjMkblLXmcnV/rFkOk
XQaWgLs3iProPatu/nlWCVu0jRs7KATpeB6iWoIwhFpRad5qjyRLm2VC0eZAqUlpQ6TgtkhHlkD2
pAHt+snMK1ZWGo/80sSYh2q08vabU6b/uTdvI4AxRZXMb5Wi+6lIPC8q/vsKUfx0at42NKs1CKC+
Bb0OsAl+sKqm/eiph87GBt4k3Q+hh0wVSppnrq9MlSnnG4BqGmboi+cOEujzvybMod0K94zOFynl
adlFrmv/WtaUtO9Dn5pErr7D80//yhuvHtj7JRn2LDqu505Q7JUpN54OgIVNjombox4j2MOu6dfo
3pGCPf5djgHSUCfjMce/MM5XRdKki2xrWg48RQzuCpidiB7JqQ7NKT/jYUWV0q0M7ZA1MC/YOa1r
ufIy+htMUUANMq76BY9BT8zb10YOfcJDCb14wBhQXQFQS84O7tAyl78HgvdSqajO+IJvLzSAjhkq
AvSiW5kkylXOTag0OANUUoyCfF+D5VSuQ/KYLlbSCMeknEJ7y9mpxoqA39gmxn5FYKR2spmCmrHl
sY/qjerlH4NGtAPeJuz2mrivtkMsyQCOZDWog6Uz3sJySQGV6uGyNJS4ROzfjW3DjB0u1roXqykQ
6oaD2zqh4HaoaZ183a0H9KQ2heyhZfJjR0EiNK5jtcsmM/iMw7fXJYe9XqthMF7+GiwMNGD1rZqK
yJ/ZSVzkUyqud1afeHsyAcWuq7F3Q3XYbxzKSXzAar2yAg1lEn6UflN1fzAKG5R2yCvTdDzD1dcd
5W5vsn56ituPRMSVetWYr+bGxsmgv7DYtKnHJe+aYlnyYowJOnn+e0B+YDqyPJRN/ypDUaHyPgdo
SLQOMW5CVLE88xDpuO25gT7zuIW1wYf2xbGhsWSg6X7y3IsTed24TDzCu0x1Qn5yroGjSd8EBy0Q
GkZNb6bciYkRTw2OGqbE1Esri+J3+AP3sPJ2IAxE8xSGrB2aZxq7enNkG9LWyv0oNEwOTvWkmtLU
30S7EsDpSf8YS9BsOmh22r7vUGsKXyRDtbW2RnI8WsTybbDM+fw+SJF3i8578/sWQsipvDoSsSa6
UdD2asddbEafvXvU9Bxd863Wv2I6Ce9pbPPzKTZAHXBJhCnV6YWUqrWeJoAhKQzvau0i5srMhn5m
wIExugY6igiOKpiqB8WTWQAGgpuIiAO1rEwj9exYNawR/GZQHsB3gBbEibnMcPfVPoiQ3xRwBtRI
0gyCGUntJZmV2+TTBOAJUOCMatgazvDVYjoTo17AqaN4yMYoTushJ3+w662QnnfPM53LuhBIiymj
SG/oDyXjvGk2Kvfd3UpZ7iaOjfbV9YlXpZbzlA77RG/ceEtTs3BnugzOhZNZF54p2kWGWu9XfCe8
07/AMMnxR3fOJvgAiz0VDaz//Fo+YDWa6YhIT3cdzVQiWKkhDgeacy1Yswdw8sORShcr6MK65psb
iSLavkB0+sU6K14WW/U2socUgu1QmJe2AKvjZ/OOgkawe5EJf0VQMCXYpP30U8mK2rt2qhktHE4+
4kGjDLqdfHyajVzNFjvytRg5+OLPuzdJnfQ/jwGdYcV6eHYyZ/dQNQwM0Q2/ZDoZhASl+AlaIAFg
+6wDk8mw7J0ak6MzDAUDRvmuGfyBi1G8SgoL20DnqQLvdruMSiNV/6IeaBNXTENeYomf64ncNJCt
I/uzOgNYp/mDHKUDBsKh0CS301PoStEc+gkSXzSQwjE4Cw1Ej2CdFU13d/6zG0C1IRiewE/SuoB4
ytx1sIqOQB+PfVQ8CPwowyAuGzck4fJgLDJq6bZ0JH9JfpY0zH7t1gDcu1sDkJAq1d/9HqE36v8w
LVF5d211bge8Vu8f6vvLF/aotejVrrk/cOOLTxR0d/9Vw/v8Xp4f4Nyo9/hhiXgh0vSj5V+MgIMT
OgUgz7Oy1MyYVVK5kZuzN03uaKrkVlT/Ax6k1+86PJumdWfFh3YLOzgIqw4KEYhlJ3DtHg0sXB9n
DZrqeK77ir+eq//TuMWfQOvEQC7Wve56FAXtpZUBJ6/2vui9kQtFOf8JgK8y98QkRnc9Wc1Rr2JJ
QMzTeBFusVMCoyx7bdzNAQWNnN4z7G+D5XDZAiCQdD7PhNhslOBL1DNlvrgGsD5iZVKKfz8OrW+b
QcwB9cXx0lMfA6qQFf3UPiMUf6VYaYrnJ4BECZkP59ftacRpUgqIh9BrYv/PDx9LaBVvU3ySJOoH
xSkHwRjfot7xf8p5mNzp47VHGQrxAsdtMf2BpSEhYyY+EAv+gKizJB06gfn8tMs5N4w/vpOhEVOD
7tOSOfn3da+hXT6uXUr+gYhaVry9gXFsPH6vLo22sWJ/aZr/oVwSeP/bxHeh1Zurt9D8OuEMydKu
5JustyiaqnM71eEymAYopy9nUk9fMx3+X/2Hheecm9Kxt06YQLE8bFpHlnhj/vLX76S/b0TBXk4W
+k5Dg1OZbay+Hj4eD3+qJWM5QfVd7588/KwozbtMwW865zzA4KweFtZFSaXUeR8eZUsE8k1ZHQKA
TPBndkt3tiDeFvGi/r6YHTN/DeQEwkH1NA+aC1cmqtzjPd1iN7WIndXDKjfembLNBQu6YG5fE88S
LFqiih6KmRUjvsdqRae0bE14Fa275yLQjL4kXdp/RznMGtOPUrsjuCj0+29wTh8uNnn46j7V5W/x
EAxkaB4XggMcIaT6vcLMDQ6dym0hfiXuETjLWK/izDu4gZnUjgU5en+ek/Ur5Sg7uaMZYhDckPnH
pJK8lDDi33hlfvcMVPjDdlzn1XUbZCH9v1IM14A7GzCb0s/CwZKxrroJFBjqKBLmfKCDx/QGFS95
rbCNLLUgWFYR+Kw5rvmPG4Yc4C4Tn3nmzfu5F4ldRSXc0fuoB5KbXLHgHze6oHrKXCXDiCKKHdmu
Uj0uLbBzOq6sfGD2eVds0oUn+XWn01pMiHGy9Z16f6VXaHW562n9c99AU50hFKdaYCcu2H3YCu15
ddZyGJU0xw2j9FqTRcm5l99ko5sY57z8zSawA8+Gjtccjd27nuhXd1k2xnW9aBCXeMmvcwjaWOQi
BQB7CfAzTPh6oYuQC1O+7hdUvYcAA9Y5OuaeC+TH7QqxSsGGCPFik4Eo/yalDVuTuLGPthepRguF
qpket2sJ5gfN5xwV1FzFNyBA6LFfXeey+r8RuWJOD0zsZc/ESiJcPmW0riJs90jCDsLJQz7OK/m3
n021uJ2dl1yvvikXuKDV5n0lrgJoBeUOXkrhhodKuxCoWVYjcD5qkmAUf597xH/74W5MsPsk5ocn
uoTHIQDGd8fg5QTaQW4N1aWdl4Ph45P226flWECyHgD4VzqXB7Wvf9U/Q12iVOcmzJYBL+00u6u6
+M+lYbZcpTmhkkt3ZgXET5ttNXDU6MCH25YHjnac2HUap80JFkwH0mWDodHxqVFoEmu1sYzjqsBv
n4tKABcuiZPHSSGQxQXZnSyhFbOqP+dWjp/2hQtzoL/hVg7c9GWb5aWNzCcFRfTSJgiM11qaLzc/
3Lr56xulrPk3rBx86MKWhc+4QOrYHV12Xf+hxMsSsH5p2GLqbOxJdqKe4DXZ/u5CV6mGKTiak85q
GPGkVlFpsEfEqAtvrbSzQWvy3BggKBeIWym1v/X5VKo3Y/iwuUmrtEXlUz7hVusMHaLS3m/qsLr2
EVXu+rfFjTaYVa7DnOnEjNsd+XJyp9YVirwt6LTB4hmVROiXGtFpnOVg/WJgE480QHGpAA+OCvhm
+jG5+/2ZbU1UvOvxgLtXVDTUsG/tpf1bMItY5Ag8h0xCiXkGyP+CEADrkEI7JvfiGz4jZcRR+y4P
gcsdY1DLbGL8bCsMYmHrHWUJ+qHUAceawZ/LxhKXuiG9QOJgiT08V34gDtR08A6MhO9z0T8HcxkU
UVDK1MDnNY8udwjzxvRxRRqFRLc8Mysj/VS1cNiAS0v1avzxKPghfZtiLGCoqiWkn1QDfhhu6Tew
jDlIBpAb5kCR1a9ENIjNSvtJ2uvnRlCOVJhG0pHDLf6i4jo5ItNZygXSWrarI+6IzYfYdwqCnPqI
Np2hHVzT3ueHPA2hbEiqZeYs0Zsl+QntcHtCrWXnA6reERP1XVNu+WrM2bLcYQNeKsdtNgn7WPlh
gc36ECvCe/fxYD574Ejz0+LH36u8Glr7IqwPW/pmvy5WWITvBODaFjaWrCu8yqulFPh2P59ryocI
b/ep/alx+9L7lhlGmfpE5DkEpKc+irAsGwpdmF+k824y0H25WPQHqCXogUOd271Vzimdp5/+zE7b
jDJoJo4WcdVeu5ZAb0Sp4jPNGjvw3mmnzs6e/Jtfw21kVUbDDcNShV566QD35gxowrl8CSsRUnBX
miTEJK81htfKh8HI6ORjQ4rMIEyNs399AwN4SZP6jYkB36FsLL/oE+kKKa4LWtHJ8S6UsZGBbTOr
JfSXTOkTMS8P3n+Cte01TZQwna45IBfXCEwPIDy+np4b7KcRpfvMa8bQSN3SqpSQjn+wKNo5EM24
RSC62bIEiO7L0CLnwCdZnmsgsoVdX2fyXFVF0wd+yNnRcjSqICf48KQGAxTzdCrxLbHH8Z7Fb4ht
2ysxvvhTg0z0+NbIQrvFA5YFn91DsF3m8ybE4HSj8XsL+vRnNaNCXE8zvYijlg/tFUXbc6FNTto4
+O6ZPEnvkL8q4802HVzZYeJGNiSov34Bi6/XYja+XperPd2hy2uTndtbbhSjwQY7Dr7k/mraTaZ7
ACqscEaENwCJXLArLMxcahhBB0udpbS9pMtIkTCTw0zkJivJ1GmUCYeJV/xiE799C93kRTqVCXNl
hgfr7xMiSmyKxWMCFJepZHPRFAJtApZgj++gQJCcJi2M0qEb79RbZgDRRrUSB2qtEYTn9tK7t/lc
rWc+ntbcY6AP9Gey6C4g8NMfXEh5kyevYyuue3WVDeqhl8ECHDi1qoCTJD0fyZWgzDfLmBjZCKKF
MSDaQ7jTrAINvh3YScUhHZPz77cKGNyZHqNTH9drQfkx7OTmQkZkpj92tQZZbEbdh7RoCS5Y9VSD
hw65FeXcdVuRjKU58H8YwcWH6nHTWKur8W1zKUZZMcVTBS/5WGdLCvikex+FRUK9SnphBJ8nXX9x
gV30gV1QSHCMTnR+GurvC6m3StCQRtGlXv7uvjkE62ve+hlEcxbWEU6AkwWBCANHwZw7vO7tmp5K
Z6mHfkBW76zzFgEwQum5t74T6oD+vGPOGu6Qd2lfuGSgcDQiivNIoS+NDO+KsdooyxR0XB1SHM6t
bkoyWwLBPcNiKjBxYzajOEan9PUVx9AwhyZS4EkCIRvudqEJLHoNbhLhAz3w3ZsO/r3s2Ar9Apzi
FY1J+sUO/0b3LrEoagWcfMmIH0CP0EKuXZga4z2YHIzA4R6+DL1LBczz91ueUNBXetxzqI+uEXPy
9ClyvHdI5MRjHXY06JbXSmWUhplVNlsoDYQfRO82clpIFmByL6MT1w8knfF1uDkLF8iNQtDanFlh
beapi1vVK/BoDeeBPVBw8sR5Rih0unJCW55ZGqF6EzpG/HOABlUOun4qBfIcLR2uQbg5+BkOLXq1
ESmerRqo1PBuUtdO7qooGGn0AiD4c1YQyC1cOpPXUFmXg9hMLlxw/VxFlMuRKCsrm8v7uUlSGMY3
NpjDU04SamM2jWNPIzmFRuWe8ivuIyUdPVIuWq2KMbZ6GWhWOPDTTjEDmGbQAk7FEY5X64cOizyH
x9FQVOl6tDNPvzdqVVsdastxvwnoXoOTJzLN+o19vn5Lj3Xm3sT8uZQX+pKZhncazvP01zwXMK8n
C9BPelLCGIrlFUGiBw+u8v7AoSLpPQoQCcDfR6kgDouh2ZvEYiKnw9iJr+ktHAAryP3kAVymO3Iy
057r2zj0y0w98rl5DlQiugSEjsqvNMk79XVoPz5sn/0lv+RYJO57ROV2lFJDY0f5agpMsAdyDISJ
oEXOeT0GVMPZwsEGuACY6hP+pOa3ZSMIrjDiedVO6OU3z5+IzS1LfqZPk0fOO4Ik7UGdL8vxpcnX
Bql/cYb6XLD5/m7z9akzUw9k9SfOfr5sH2KjlclCD3lx0lf4pDWeSJ8nYQ99CtRDIWeEi/1RG8I6
xGL4EhHpXdbPm3xAbVOy1UaJNBCMh2AIglucGwW5VnbZTLeIHexkA65l6jW4YV8BJLs6hMCwGI98
8bxtzcqV7dAhoZGISbW80N/L2HGAIJq5jrvATgLGtZ9GAht4wAPn6ZipDMA+AZSI734zPeu23nVm
q/05vjCqNTknelIX4FLmPPTFSyzMXxDf4C1XlZMUbveTVM9fA0XH7alKxA383FR+QrnU8myfLLFN
GTTu/T5SGtv4E3AyySCV2qa4mCQMhcGJXggcW0ogPRA9SLNMJb3SJyzkUPq5JEVQ2yIUAEgquFwT
W+9Cpd0P08JK0ChhEKPydCsbDJci1Ibx71V/TMMqnsMN/Hynw45wphL5SKfMms0o2LuQbc0Ba5jY
SbOLQrzDSfM2pZZYdyKg+oWpYOQVi5jI3nTAKLqKerFAy2OpqYUkxMA7NIkTrNW2l2kiJcrnRXG+
pig21I9os632BAXtRauPfIgf1Z9HHtDw8mbgBKdNretr66dz3GmnMVOUwc1CON/mLqIDPwA834Ur
YfUVNOultcz+8LCvklRa6+sgYwelacZ04WaDAAMAQSGryDIC2if/HKj6/5ogroF3VBteP09Dnh+o
OeHunHp4mIOCRkInD52kdqxODE4ipgq1owQrnvuY9D2+gjzRcZJLx8rexPkgcb8AtUbMLCwVxxec
grtEuQYg/qb8bUnIFBHjI/OYv5gS4P3h1FZuulFWwEF5tAPGNnIH4Z0SjTpYKWTtiUTySaDK2Nde
b2OYC4MGs0/JhBfXsmL2SLeurjuvYKYopK/xnM49Nu8zCxvD1C0CpL+jAsCPFGpNcFKefxuEURBZ
O1erb+lmOa9Qji+XVTlIDlO3D5GNTlMwDBicsR75NrOCpIdQcu+HTNGV4LEBN5eqbxw8DBqnmU4w
YH6ixJBZl+luFaF8/xYGxD8zCQGSShMs+0FXo8IU2Es+gsx5t9clpUqCkjBgypLYpAHl+ta8iQ33
uk1k9AfxI1Ckzhi2xmtS0IdXxw2ut3P9HgSXtEcI83DgOs7fsPlR6Xmgw3yph0Mu+fFpMikooPDW
SYLEWoDn5LzWEgClCUzVLSpiECNDoe982gseMd/Gdfi60xkmjd5Mz4jpTtFvnT37epcvdjrch+jg
Jcsa/UoPuJDzlH9QCE6pS0OuI+bW4VMnLs1GXZOh+k6GUnQkgRDXZCql1LvgOb/CvkYcCc6JPzVJ
MtV8u0OBzYHQ7kr+adiQL+TItzU6Ihb1ITGKPyVEmLQ7BHok2De8fy62aH2DI17HvcTkEP+YJNjB
Zies9AA5gTbVlEesm+gZMwfU8adV0wmoo3lEeF2u5mOeahvqmAW3F3NWgyiA5PlH4USaVKR7ODZc
V75Cl3iOjz8ebl8mws7yYL7R6cAGQBubF3JRAZ8vmyMh844FJBMSB9Q9XQ/BSlzCkCj/fAJeViO0
yggGBA4rcGWZrG8lu3VjtlOSJ+bhsDsIybPDOyBVz9FnU7iB4PwEjfCWKNKYt8i0ijO5X71RtOKb
3s+kXuJPrB3rn53bJQMU9G/dO0I7lp+1VDX9hwADJYElQXXQXpOwf6FFVNVU0egOvxOWbQj5jBPJ
1tqLMjygZoysGrUmJONjfnIwpHDSfpo6OBI8xGS8Bsb5VcW5VYdPf/gFqyZfrj9Tj9xtNuAXtMdo
TviA9tQ79bZUsf7HCvnLuYqmKqIZf0BujzBljeA+dTmsMvXxi0ZpCHqyCadZV+yJhJbeEPA7P0R2
9gmepAqfJFFu0wzdaONKGz4CmR92tEeutk0UaPjvaXyK3vjszlYihklPjG/ZOg6tX2cAgh3u3zM7
rbB1+jfmySbjTPjSIfJm0nAgum0wnOFNluDvJcqrRTiUhh8TRYtdvctuYixsIHmGPh+VfOP9i4XD
IGvCtw/h+LV5aPotMK79Mkh/o9vphuI5V0USicrCpuw6+gIvcTvtAHJYJWqk1521WztEupcebbH8
VTsGk2Hca6XaKObQ5mAu/NzfQYd3B5OKfguwuqE+Vzm/ySv7heQoZBXQQoVUOSrRt+DsnGnZjS7p
RJzfJX+9dAnXy/XR9tubkkzXbcH8gZ4ZJV0A2bGudSllNpMi3yhtWF8sVP55vPUyULcrpJ/AcGuU
QuVHDvpPerE0VnEU+bdeRBB+ZdyK6D7GThVmbJNIaLMjnT0uxzkA9hzGcsrCqy4Io4zlffcoihGC
9QpgZemUVtqa0i4cQJ3Qe+vPKlzsuX66HCLw+lBuSWNaJBwXgDZVCxmC+jsBunq+8dsKBEVdnx3j
dEDrcH4qWitWKU/OVTid5/ZxzdcXLT7bzMsad+RNW0pbI14/Ww5DxLMHa31gp+UdqsUP7z4bJRAM
1i4AXLVrDqTbBp5yfKxTJuykzp4laN5U6Amk9GxcyUfJ3XbgwLv1SZxXAiQAR9uBuGFSP2MAqclT
R51kFwmu16u7TJWgzshjmBxAduzhtWrSzGWTfMTVOVssW4APlPU7V08F+0GnkMwEqC/+0aUy97eH
5cp1bn3zqfhb+eBu4nQA6+Ikeut0HYtS1QVTFvYqchG+FHpLMF4ImSGGh7jmrSvnepY3yZZ3EBuv
9oIfYhKbUH0ftKRUXh3OGK66SQWSdXvxYUn2cwzeBQUHPeiqEfBX3s+gtEbl1nHFTMQirkVfbmwE
+unBxCXWUMtpa7txgCPP5lTWD+3SdPe6ehUGmHr7b3bS5lS4u2RavOY+BgW5YIjuZqU4GR0imkDs
apm4keCKwEudZ6+9yGlP8yzZN+poZJ9Z/F8turWNJmHftGL6dHW1KJ9UgPjPua6TyMIBW2jv+a5W
MGmYEHtsGT+TemAyd/qevgWR/HdoWyfc90t2JZI0cB3BY4Xy1Agw/3zyukejN/ntST84TM/7gQz1
4qSKwd4rSEJemjs6FhFYxLrOPXGnQrwjqNl0ts57E6irADv7/IHaNcQmWUVWsP0nV3WB2tJn1wxR
GB+T5QpXtv837GMmpLct8+X2MkdOlJpzEJ5a7rtP2V+y7/85/J4WZNFdQhl13F/iMT0gOimW6j/k
VviQrcSuSZcDxXSkBNfuIWveZiymjzWNQmMvUYnmk+lq7lVghcM91GeokYC9Bzat8ErrQe12kmLL
imEYnz5fbuIBk7QIrxocYlnK8MX9CdelaenScgwz/keheZSs1vIJVzy1JKhHvokJeEhxu7tyC5hP
Lwwh5IpQjDC5T4qQrg9JGyaSy8OQwhYm8YG1HHiUZdqkoLbhf9oQhDvACEonMITfzo1YsJXgOS43
54RXrFjlu73RNIqqW/hOKy7LwasU7CMptW5YQLKr0CyGPUcz6Xgj23+ktk2xD2Df5zSr04U6dMxy
jrB8/v0m5bKvTqLQdEwr+BbPcImpzph2ijROqtPZxIgK6ny8giz6hVSlVrhPtuV+hK5qbcdCTM3C
AFiUsl04ApqFduD7od8zrsCoqp7Eo0NYuNa5VuzBP5AlSPGiUZlUQp/OqKH5Z38RuC1GqSSO0HVD
K1gg+I8WMFy3FsJW1RlVdwP2/WAgncWtJgNs56fTDjXt5d19fKsAalUAlcb7DqHv5LozLWD3GuyM
2Wbz5Y4vPL3tVfyW2d+EdaktNZB/+hKjCNgTqO2bACaPnIu6uWpMEFDOLIx9smTJ8aK2TGDIjxgg
86zdE0s1QHf4dCNXnWY/Y2c8CH+47Nvnz9B9V0bPM2xqd9JmBBfEieZGQhSIY+KtPg8hHst0ws0f
qDyJaqsimHJWmUSg9xwEYH4JdaWbXtSiFl0zbtfx2X2zsvoJqB8i0aonazPmgDq74QhWH+qocCDF
vTqhkI9jQKDclnTNpI4MDQCYQzu4Ohd32JRvoFlHQ6sWzxtwfkIp6zBxBgdScUQUk7Qo5smUfJR/
lOVsAmwChJv34YK95+fkccayWU5PG5gwGmqY1EU+pvFPhw7Othkoj8wMzoLdx2qar68rEFJkv32F
fbUIxlx4tGbHoIbcvvl0kaqxWkkaJCVusc6iXREpEJRPJFWwJj7QAt7Zc9gtiQgyBYp+BFjD7oLQ
JJC/ebb75mBGhwZw/ymUphu0iPq1FTp8nm4Km+uRHyMv2IcRfPnFxAChAXFPRG2NRVc/QI8AualC
K4wJ7EfqEUwY8IgH217sSrDMsyhjqApbxpIVgsFHLTC2yXLriFnYtIrbKmfGtTNop9GP7YYDgEaa
UT0n1h9236rWj7/0aMbiaFXce9fpRPV9rp/EqRpmwcObR7YN+wI3u6bBIzx/AMo0LOUrcrZaJqcv
qBVR1yh4rXHdmUPBWIQ0CQUw4K+gQOSxu4WJw04Xx2Ge/pYyCeuwZHauWGlgsYE/9lUEmHY7VDm4
VS/bC10eFUVftG0fp98LxqrQOtS3MUZQ+oTAf1GUNInLXx8rAAOqTb0uXmI/dmzFp4QyWhA7NHqm
xooz5/BfCIelNsEluIN4FcdQKDRm2X9LxG3yICSMKjpNQcCINeAqXSoLJbGfMIR8qz1e0ANihHqL
t73s4pVW7hOaHTxcfPn2cd6OUf8UH6iwAmCkUFPA9QULD1IZ29zAtNlYKw1wIrTHnpNY4HWoiIoM
bus7i9jQR8B4NQLaHd8xWeX1YGIjCtVlvEnV/EcIMx5JddSJM4S6hxyjMUq+neRBjYrNtsQUHNWy
CC9IKCFlTGwz0RC0u+ZAh6nCd0GieN5fEvDLKx4r6INTGOdcy1jQ39pCGmbh1LKmwOZf6xNOoZgw
pFXfj/cdPKQPRrX558Kj70OEdIp4uJ5d5M7VpOb0Y/e0Q+/48zwnqgrzlAGc5QRuxEF4b3+aWqgU
QiN1yw6jQ4hCBUmndN1qXBO57EZd0qG+/94BQ8dPab21ocAMZSFNgErtS/soLnZUFzeYsMFtUaY8
hL1abvb7cZhQzc1euXlZqIaTvxZvMCxXz0QxljhaHtgb76Odj+vG92001KHoWyLKZODWEAz4Y02J
c6lFK2zVL8L8/qYcEpTXkeL00MddyUJPcWt6nGfzhw5E2nJS3AB9YWs18ocIQGU4eUvgO5m1jvzk
rjiOYaWU9ML1l12kwvhGsr8BIchpaRjnGpwrNRoj1/BEB4kl77l5aPhzkvLxgKipdUh7VJETS50f
i8VEVuFsACeT7hRf1Pq4itKrHCQ+jnhCADZkjDgo6ImJRdSzFyMObqm1ISZGOuYNhTfxuzm+97u6
McSGIGyXinPsCRE53KSoEzakFfL4GUj1RVTzLF5q5HO7bbCVsaqTpWPhpp09rlCqYYFEaiac9O4f
zebPke5WSQeGvCNqrSLbIaF5oVKvGXOgjQF/+5+J+5HU6ooT3B2K8iUQI0yxz3CZa3VZ19SwHcEI
DdVDX2KrRXYuw77M+Jq+8p5J0b4pbmHSosDpVfF0ENIia3akzwJvYM4dwclF4XX5ax2lgIC0XRCD
+X180rO+AhGSExeplOHFYoqkBvM6+PC9aDHdktUkpixzQ/XMmaL3aj00hwy7DHilM1yOxx2jyDwa
GQo9Q8m2ReJ/2WpeXdzqvmNSBVFVJLq4lo/qg85R4F3g9RwjfpwMyk90sAy+FfZB/pVAWvN1bd6l
w7lowbLSukjBJ2eXXdPx5yvuRSJLLxXMgC5zNQjVieq5rl0QV8jy6/xIzSlCZaTAYd2+eG4srp2s
G2oZIcoHs9eBMAC1sGSevF8d0Pv4xcVV02aDZ6TtkHMgROB1bagWUkgIfZYkDLPB+3jdyLPBFVca
oIZrR1U6RmvYeX0a+gOMkp3Oa76Ic/VSSpcg1/TLpqQTUBBSH2q+Y+GH2Q8/KxFGIQzSwkhPT7lk
+zSkXNaUDjvWRLl5EubNu2WxJIIYs54UUJwwR1q0yq7mACfouE/7sQug1h0xvT4ZzGjZPtxT/v0e
hrMxK5H2zjBxaMKaS5PRfH0cc1t4EXi3gq1ISyYB7j5oFvFepro3ikREh5iNo+0b7J3Pruye6DAR
+L0aSD5PFnk47X4RPtek2wkbvowlIwZfXHimuSUxU9SFnbWBlRBHHMWrsLpNBGFwHFlt7EaRWZyA
7SPxTi9cTTi4P2yYt2dsXIgo4GgLx0GfmQDBXVysEOUB6at+4mcRopjw7gbQ/gymSYUvr9YoTUMi
QZuh3o2uoeWOKoWTg7cH6scqafOchYIduHsLanP7T2JvV7/RypJp+UFS8wTmJEzkyxlHFD5w5/zK
NQ24WGrOhrJGPKsYXpk4oBEAm4H9VErpuxpxflg7JtJ7U/Wc6H9b+q0n21uaMxLqjOsdNrfYMgwv
thfSk50gJZ/Blw2eFC0BlDo9y2SmeqHZGAJgcTxIgIB4u8oJkjX2VYGonsXOW4FOgn1MvnZbRnV1
Wg3uaCaOohyCacMTGg3OV4UNpag/lD4dIzb51SQvx3Iw2Fq01WZeLgcz2o5lj0iIiweibpoRezS9
lv9/gm2Fk1YrQf0kf8GU/4N3kM8Pe+ULRfvyI7VpVp8vGCTf6lGwCaSEErkkr1rwBlssRIq8lVnH
uMLvRT0Xrq/rcKrO0G+xUVgXmlHPTEvfaMsjCz/mNNu1P5vPrA0BWUGZHYOJCfZVNzVXv6LME8ek
xQOMw5DJykgoJxqK3ng8mVtSCrspUqPbXRzc4Cy+BpEzxklcg0derqUwaX2zR8gqJYVUgA8V5f3K
AGopiEE3quoh7igm3CvTmbpOXJqnzRtPoRe3dW4sijzTEzB3EAe/OkbsDVQd7CfZP1vEAxRBNMoL
ingNvTa0LpoH2SFm5kHHDOfp6Qkfeu+Xa6mhewJkwGAI0Gd6wfne9Aum4GD1+xJJS2NK4MmljLWW
E9m7bA2P+GLcrasITYbHSJa/KN7t/8ekTPzTYhCSFU7FZA5yIF1VT1Pdc7kDpmoBCgB0Ae1dBQBg
YhNoKXPI+Yy5rnBywmxODkYmbZGusHotCIOKHhIm1vMHuet+v4F5LmD5vMCUhIPe1AvRJ2em9m/A
7+Ni8XJxtcPGM/EiYfWuw7zal8uuFv2ilpxd+y+5EDZuobayb1YNZ4R9iJaQxidFuYOWjy5Fzwp8
hPkVGUPCia8PYfoPLWEMdWagAQo4+ZD0NF6HOH/vzT9GNGfd6NvCPTOrhRydsd8TxUY4qQ5055Hy
aEFTNL7hgSt8/F6BabfHsPMU5Mfd8T21BwxZF0cs7cudkoNhc7XYmUkcMFzv7wEtEKJDs8FlHtNt
JL5DXTKc+XFjhLC8xYBlvE2UaIuLDjFrXrJ81cykWCJkVqXR3wxnWAvNSVpjdror6SBobAhdr4B6
DuFWTGpngRyeZVn31IsWJan2JZEK+xpWQ1rfZnv9RPsmhXaOGYnhmhhGKUk+F3XPtEwcD7vHSdPD
Wc0Itkmx+TUYKdlE53kGujYijj7lyOKOZgFAt2/0Mts3v1qrDFr2zzz9ZPjivCfoaGKx49xuw1OV
0T1PRq3FdAYaqOr6d1IHHs2rC2nJIys98CGuO04YZoslOR+L9aSZzc+Rs5cYEorIPDcHG9OEUZgj
hil1sOs1b4a60l+N35UIKvlaB92zwrdWmoVY9/PJsOU2EGbw2+5kb1qeYjY3xUzHoFvi0hY5irSp
T0PKJfMoksnvsqUq+rrNlBi51BkqKciSJod+q18dDRSMEC9un2tkNE/Xzq5YiFFuQppI1sIuJSm2
2vtKAIg8yZl1xse72Nz6vtdZqKP/dL1jdMWzbEJU9ci9+lwOTN57U4LU79GpzD6Mhuwif0kR5Udx
HRFphUgiOLEhvtjqVYle9jdbCKsrDsa6vUIKNmuEngf5iyzndchqav/N1prVGmAzMkYVipktY+/l
4AMs2jPaTh+vDFufNAxerR3a2WrAMqE4aidCarel1H5iHX30sOpuqvkPmYIaOAdmk1JxL0TQkUfc
9eZZ8Br8IwaBKNHVAYpDJn0bbhnH7SoJm+INnz+G/+SCcyl3EzCOVkNVarKfRqgf+IS5to5SB1e3
uDa0RiQNoU3GxhXFvUuzHk+3UuJT8ZKF0ERmje2J88cwzTSEfiK82hYpL7+lJV7dLpeOEza6/xzK
dxIb3qsKJTtZ9yFH1l16S2L01D2wsYimiOu9p3aRL4zEE8nGzii5Yw/BndpXa3Vn1eA4BRpJ3gKL
GpQ4Fwipf5J8/YPQcdzSuEGNu3QxV5gqXt35P1ziwgA5Yw7esK4zMAxsc/r6uChgFq4Cxym/xTJG
Stw4wcXqBtm/60kHJw+f9yxUoOjUqGhZEoMVW2KdpKO7ZQQvLrwBe3AcMOSIfdKmhNzM7Cl/PiqR
aJ1CwtRBZO2nPxsWsyPPvos25lsqBTMPm2513cyZtuWg1VuhhcIkA1qfXCpAaJnZ78mEebUhoVJu
JKGEU3M6wU08DMidmD2BoQjFthiOdYH9xjdCTaEO8+HtnoDg3Uol9XRcTDOqPgd3P94ZpOcbRUX5
N3R6DTTdUpXDK7hAnMqQxxyXO332Ydk1lTLEXfXZfCS2IBvZYbNlaf7L8yJV6/ZqJDU8P0f/RQ1G
kDnvZQEp9tihvw/ijkM5u4NVpVFeU4BQsIrIElQpat7g7cOy9G0W+OY9Xp9V0M7YN4m0+yBnzq/R
uNbLh8EU03N5G74wv44IIFkgjNHruOiYs1jH0Lyxr9E9AI6ImOZn33xhnAcrTo0pcaicCDZt6ktD
RZutODN+ZRUagRCvYnFO1z4Ja2DWQFl0kKo3xD5B/5WdtHffMnwW3DbtLSkNJCD09Ie18maW6tqY
m8DK/DGQ2Dtg6/Z6DUAucQ6CkmNpDru0EgKhrWbsfXbZ5BhHZ4gdZBCIDvYGTNp0pB79R3tsAE9f
GkHcFkOh8E/Q2DBn2ES7BFDIhNB1U2AI3FIb9tufiYoG3jeF3briML8lrVqRTDDVOLqw7QRz2HA5
NDOlny1w2V30/N8ykmaegrlqvSs7SabUkYbvQ4CblqvmLa1/JKVQft11lh1Tw3mVrEo6ysS6fYJI
l0SaSItbalSNv4ytK+l9WeU7+Kly/Y72lkjKFdojn/DjBSlgBs54EY8JjlpGWPlu/9eYoQHgpLMA
61kryZpob2JtmMfbV7AWRbvW/XVSX9yUqEaCRLCLEdOZqfr26yC33DGbQQP32A35lTl9nir+m7AL
8sOsqSB3hHj0xy449n7wJTS19tArFOjGJdxQh/Dg0vs2czNB5+KlDFcPwnWxGB/JHzMuFSXVTmcb
x7eNNijMebtrnz71gmm+jHvPA4GoomhTQhqk/8ssnKECejBpwVPdEOCR+E7hMqdqmzrNMNu7IurG
5zGZkxNTJaGYHDIx3BVohXHW8F2H8+9uwZXDho7eVcuG+Q58H+Uvv0os+n8jx57VH5g/b5BELwaL
Avmuc9pNKvCFefy8m9qYhZxtrnY/Eyc8dbIB2rlpaakg4aRkRVokmPsJpRB2gUqaXH6hLpZh0S6c
nFDO3jn4IxxfkU3OLCeL5Hery4urCtd/PVG76MXvrKzwHr5BZSBMcbFZ1mNNgjOLMmr4hBoKKU0E
o08NUcaKKHZcV4NtHcwjEk7rkshZaMgaw7hfqf4AMDb4a0jEzj/SMaUSfz4CQHHRabQSGsECF+iz
lmb+GZCJae6jRzFWPgZlvETBwezmIE493ckgFIWLnOOs7+ls1m0N9mw939qGTKO/SlhUSDbZIZt7
X1x3PhAQaTXVQX5m4P6xpMBMqgejkHuJGQeTtUIIBif1MTMqQR/b6W+dQPlN5ageKytY+r8PYmDw
QN0vrdsBXUEAV19vo9PAk1HSqYg+0JjpQCKJB7kHn6InZhX157OvXSyH4aBmF4oAZO8N8Qi1Sk8o
Cj8K12v3INBLcor/ttUhGwqrcg9XkmZzz7oazZ4fmYat/+vhoiXk1As7jOcg0PR1hhjKoUYL6tza
HfZbHj6oh9uV5AZ68fYdqKfaruiBe6iN4QNHhdEsOK++dwrUiD/6AQU+8j3Qakza0HU/ADXX1p72
fN87gBLZqlQNkFmJ30r8wfb+rPJ6syjeWgX2aF68bOCsikMFiysMIv/snrVIIwJpF/W4j/L4H0Jv
DrbtkPvY52K584j64+2QKGSk56SxGydBsmpeJW/61NYdcv9xhdpJANyxO9n/DR3vRm9DcgG8J8QI
NB34ju3puHf/GHcanFAxH4RCeSrtoe2/bBLLgo2rqqC4jrEOZHMB8dPcQaJ7ryfaPYzKIk6HpY7X
ewPN5OQ+lnl07eVC6jZjhZdPl5RwSwEzZ2+0Wbbvg/Bc8TlpH/V45/muovgKpl7EsONf32R9/1DB
1LTWeF1n5Lz1cnGzPK2d4k3zxuyG17zYyJB7/KsYaxJkqmpgY47B23dlvW/RTvl4qkzhNgt6+1Vr
Gw0nO0AgcGS3G61cblvv7b+PsgDhrVkKXnCxQmkBTWKaP1tAYROW29gvE35IrJtjh9vXilIhuZOs
H7BouMe/9T4x7nhhIvgiodVOHXuyJx8U5qZLTIHRKGADKoqNUAl7qOqagkX1Qh6ajEfoZsQCiZBg
4n4pHcBgQSVjTuNPtYa4H9bpDmkjvTc7G3oqHyz0yjFaOUph1n64Y9E/kRKKj24Iyv9aG4ohnoya
f2wW4Y44f+dtiC4MPW7DDPilpxyV01t88gmm12wl4z7ITqYsWFvq/oIlUv/aeR7U/C+ZxYSp2JWe
6MAvuA5O7bvxOBHe/UkLCdB+IhaDN529oYrPbuPRnGFGIaQ7Ko+0cfzOahk03TtuvNF89Z5ylEuk
wSqxoZdEbp+gL2RFO1mU+MZnC2o0/E2NnupvG1oIU0owWHjKRxyYlSw4PmaeVhCRHprLMaSQyeXc
pJadEp/tR5VciklQHaZSkJchurlQmBDfgk4Y9lxMEQGqZ+xFSeAZjl4cg38N4qLpN0htA5IdSjB6
XCJ91BqjfK9vgg+XqfiXrQlmVmvfC+azp5+LmmMckWc36SOQPx+VO7UtAq8hFivjYPqohfBFgQle
IZtYbVI289FLD/9+uVo3pGBBBIYKaDzrK2H2rsH3YQCKjtopH73aewqErju3QtN3tJrPNmvHX0Dy
yDBzdM/RGYnOx5IrMGxSbbrnBBXocVOkOFM/iIkvStce7HWREwn2Q/9F6BTXmrso/+Aku/jS/W5H
E1oRGniTF9bE3cqO1vpyhh+YaaVPHwo29B/83G62Vao3pSIipu4xFMMyB6PMeStGYIEKbTBlqEcs
8MVvYNZKGBbDpPYwXy03izJAz4ofQidhCHDkz8t9+gRevUaXagCvHqVAoPDBXw75D3S/xQ1ByttD
O1Kir0VEnmh+nRNcZQ8vVAr7bpTzYOaiehhGI1gNxgqwaDOIrhz+0O48TT0/K8QPMAdSQEIhU4l+
FPxEZYBlkMMmWtY8ytvrU8ayiwK3Uyquk8pji4wT3FrLRWznrZOz1VfoGAytU4CnTz05VcHB38EW
M9u74xULgPX7Oy0CxndpGFLwQ1rlKYEEycsFBir11l7Ai36GqajTL/j12ufCyXbA7+42KR9ZTLq5
4VnIEqH42Mea3COd6OtW8dmminKQZjTKovRll9/apFu1aw1zUj2Gxj0Dp/e2iX134kFlmknI67tr
r4BdaaDUPGI6OdChnMxNT2PyXYHU/lZ2B4JQvIqsDtnI/7QFjhL3frWJQIC0aLlfcsikM+AVm+ab
1mqsYwi+/Uq+uUysPmXXjvQ83DbGP3SosoS76jNJ/lXl70b2MKEjrD+sSAC/O/0TF9P2LPP/1Ef8
Sd9Vbv+d4ooACxi5R5td6gq59LqDsglcdlH8EdlcoCdr/ApcgR1gkXr0jrOMpFNyjViYiEU8kVe9
XRwnwl/p+/iI6IhCnoM2nLseJ7mvdVaM1qKasiOKthLnPo6A6AM5U8xRvrxgg86YzZ6ZCkqMSNzw
Q5T9wkVcmBUz3GTTifUqz5M8HDAl4r0wLvNDZhkOGJTWAfC23EdXtseRV/VKEgFcUsXgFfb52pZv
FHoS48BFEQm/MCJQWwoMogQqQDWOil7LeueHnEknkNNh+8+EfU0PLsi8uyrzPYk6lS57UP/Gu7G7
MA/fYou1jG86egeu9OVOeLOnWRCLanu0G2a405QxYWaYr+bnrJ0NI/bjkWRpTC5uhZp5Z9MQX10Z
VDFeppT1t/Uac18Cu5Bth/jtFiwrdD4IUg5QcAI6BhZf6pLz4PzUp6TXugPFCATY7q0vGkNepIDc
61kDneZPwJVzsJ1IkEwE+jZBDWlyrA2OfrfCqlzMqOC2aI8Yq1In2DJyzupB7YkRvOdvlBtBSvoH
zOJIgyhhMp+/4AbgxINHwmu47GgwGOMjXU5FzCoLEoMRHdEBmwVu653W53cweecMBbWEBC2YWTh0
sKex6tv3APSXV+ihoO1BY3i9Q7qVm3gpISLCYANIctaav6CNy+ez78H41Aq3kYqo6ugBfRV8JB3L
LnTe7nIvOcsM9qVNMPrh9VAR09bJXxt8aZsqkHZ/SLZkUCOokNh322oNZLmsiC1H1+qB2vxkwey6
myOURBUrHruCR/In6+/FaC4vYCT8lLNmENTDZ5OTgPyFubELmbljHZJjxjlxmTBFQzY+m5bOtQZh
W71G7JbO8F3tuRCzanUlOP+P3idNBrrTcCHfNnY6AqgNo/ZTL9btsWGKet+MrOvR8tWEoPg3T8nB
OFqZSXe4ZuxvXfju1Jrki0SnbgC0/0sTrGarjoc8akhGZIXTI0kUaJx48qONGC/+F/dPMwmF5QzA
1J7LKbRmgSsQuPvddloJpBWxJVaxMbVPfn5pUtKHw3dPwNbhapqoYShzcKIeujjN8G3mAhYMwYbE
zxSD5IHr69gw/61sBgI2Dq6VrKTeSVDiOieznlkcvEpRDR1NJINxStyFhT/wMVJOo/oTptJMQvig
chPveObJi7wXHNafKK8w29uVFpwn5eEUSXJ4pQu+ZTcpEPeap9q8qk8ChlcghCzfHjazkTihHurh
Okb7YmjQi0xrcojpXvaWdoE8fQ4awaa9xPR2UjdekCZtuQfQ/9N90uF0CN2bEth6+lQnlWQcTfBj
oi2P3j191DW8FVZ913tN/arZaxFJk3nPLdpVFP67lUGWY8yy6jp37/7jJ3jG6HuzXRa+sJr0GaAh
2iCLHwU645d7Uh93/v1haqqo8tj5rsHiJULcgaRlqSrZ+eghZA0wbYQw6BGkt4Q49ZHTIj9jWHoN
OGJPsYW1FLgmRTBjbG1P+Q/9oeNgRORLkph5j8OorE0BZIfcLHNOeOinXIdUJWkTrdrVdgTmcIVV
4906HPGyvApDbND24BJjrw+mWneLuogHY6mklHd7JW+3fOajZI1c/blAh9Yv8lI/4ZisWsiNEeyy
4HEuEk6VNLrB+z0v8eGTMegyFAbqPMj1+Q2dXmUhDDU2EALN00m1s4yEt4y5AcdgSgDQLerO9M3x
8hTOZUk8iMRSeyXmh6mqcSwGNwNZERFZoccUgFfcb3dNdNs6vkPfHnCXZIVqGEF3+PC0IuYG6itM
6euKkSHQAd0mpISL8sJ+d/lyliaa+6F2sE7rzxmq/ArcqreMpiLfg1ai9sLJ4xohUVMmNCoMdXrV
QAmfrk0lkgdnH2HXMMF6CnDcl6OIjfHbQj/WNIUs/Ds8+9B0THQ7tPKBeiyYlyyBWM90PK3TrpbB
NG+Wx3Z3aO/lYhdwp47nItc+a7JIfA7baexq37Cw/7RqsVICZkbCKYWpZAjeJTtflYaVRdQ/zm17
3lb7HQO1PGtuUyAtCSl1pAJ8THFgm5FpnW/LzhPljEXUVTtGq2/NsRERYvyYU1/xoGM/y5xeTFJP
pn9yw0b/cHv1mxr7zllwta5HC5N8Zlm/9STzm+vPpg+mE2WQYDx4zclSNCrB53HYqnYQo5LJaR3G
3fHCpTQPEqV0qOFqe7u5zwLgH1ZbqNu4/O+H8gTzp/cMs0+3IVsfIrQ+shs9zRW0r7XHTxOSaqQG
vSYbRb6GcCW+q4KeoX49Oor5CMVSM059rg63AVvI9U+lFYrcGLCqKsT+f3Wo3aAAw9Xy3Er7symj
Ne4yA7zGrqhdGd63GN25VDDW3MxjU9APiBbZ5sg2Mv7hxYjTC1yV/vYmroNt1RlPZA5CHCQaUy1w
E2Hp+LjAgl4os1IhzeNz4qDs2FwEwav413RroZOaEc8Ss3Bue99E+zAIzWDJyucCbnCIHDpA366G
xEC7/PzXoI7vSrf49F+h4m2zQv/KJuXrB6UG8s5lF9YSXTAUOUfJlAPT0zX3CSrVDbKDEFR8L872
UUCEtFlJmfXus5ghCZce92ydXVYzjBgVSgPRa/GVTt7irp7C/3VqsKHyXXlcVI+Ck72UyCK4kDWn
+TCURBg6TdEhGOXvi2Nx7Leah94GwbNXfUIrET6qebWFM9/SbNUWiQAhI1CfhqiBcv5I7FHSagNC
OW3BzhrYVJHGGM6S11fZvLnLxhICqNv2kRt/aNl1yJVx3ZBpe4+yFSTLNNVMUiiqVc+oaOljx7cA
oeN45zDPJYIVsuOdrvs2l8G1IPgfPySpC6JnY9XFZudt8fSi6zp/WR4Krd+5StKNwlCk/XoTYJpV
c5I84fxizypaXbxrWlzMD3KGalrJehhdKe/Vg7J6w5z3CeLXd1d8NtT5uSJyzFPtDFsl9s5SIWoV
VS0G/h0H4/d0xT5VEAgrP5Bve4MSsuL+volsfPm8REQyRu1ooykVEI9sHy3ZXaFMj6OQfCFMPz8Y
4SDW1FcOTWQ7JlifqsRWDNupCV9tzzvZGRX9CopOr638d4x/wV6X5cYzHuS8W4Ao6YVKrF5w0mAw
EF2uMY2IyzKavEE/+fC/pP6BJXrpA955KsJJAwe/Wk7+swA5uJ2/HY0kSP5RlG3hXPKu19JYBiTL
fYWsxdQ1Mm8jxDAtvmOec4l6+uLTzIfwpZ7G43aB9IBLEXlYB8gn1fUsHahV/dCmi1/CL+V53YYf
7iaf3oOSciMiQh2kw5dCNbrdl5FhWRpnq4TtCCknS1OVevLUSn83FEdh6JN7G4EXKYCfL0j82+am
UKL3xDdScbjHoM2Uz8Zb/jKYW8vw0XQhsMB6AwMIDeVkWYjMPZSiMBdihvppe3yBq4PJJvyEVyp4
gkOWu/AYBPL/y5OMnhT2rCvzcpFNq7st1EeeAjm3Ueg1iLPoSTRg/su2rfsj5GzZnuepSUZgVeJA
lQdddRVLkQi+6LzICCP9B3xxFNlHRkK/aAzGnWtFd3zStAt2CzoAiBSc2qkmS5ZsefP4ug7sbZCY
X/9DsKlRaJw4Wh05/qOrLpFppx+AKLbeP1jGKX5gSZUV8x6xp4X90q0aL8puns6lW0T/ruqJXyNm
NZyX05o5ILm14df2XEuAwu2jImTbOlE1ZC6byZm5/TEU8k26nIgO8xh+lkZFbxLW/6F1G1lHNs8m
WrjPE4r+zi8dS9uT082XWloGwp9hCrBSsjRzVukHfdm/Cxl4MYZfOmE88kLCp3Bc0tZYOBew7gS2
x/zVnHLVsHOTfWfAQ4uAR1WuYGG9oZaLpLc24LsBEvQLnYTFgsp3jtqlsU3O+8uozRjEn9taYMnA
elSRUNedHp3u6ZWFVwcyjVlisRBcqfKzFANi2054FUqHrlgTFYIRw4rS4gOh7Q80IDZ6H9IPwGwc
W3lqsxHjKq52XqR7IGOJ6TQjTwFepBne4uB8nMWYSVfQy1uZ1A29K/4M4xrVJSw3q9DoKGDY9UbC
4ulTl3/S0PhfPRMy6jga7pLQx+DgawdKDT2kWzpAC25FVaoSSzOfKMhBoeqaFUxxUecz/7ucLQWv
S1OtnOT4qRuZ7FgqLut58wX+sjpXqf20cyatqgFpd1VdQUTNun1eABUblfi7Vb6NCTIS8jKzhx1z
4oEyoR5UhlczQ+jHA5K+F3NHN1vCeU3lTP9MlWc+xgW37AyjsJkRFCZIl4cSzMs/rjuHM2f81xSq
MaKGYYFdrqkKpInqCBI7WYYz8y/FGXea14X98/uJ9DukL66dZ4PeOBfm9dKlZyB1ALfHDlfEpUuJ
2XZVbLzyyoQfGugPrEdf9l5QfjQedc8JdYcQAHE0z8O2E1tX7WBPFc0SyxAj551+K6CCulOWdbIW
OM8anxhPd9waWN5gp3g5j4iFztnktwdEqtv4/B6BLyu3CXMPd5XD9F6zxnDJorrveYS5t2mq90Ng
fKh+12/xoX5j6g7MEZxtuupIx45UzuLTH9MMq80nyAuYF5gQkXmAyU6W+CTLkNqjsTL4HEhqjSZN
giBVRYds7vhT7m6Uia0xrHwwyrYz2P3pSB0nxflFTJWbR3dRdytgmAuiNNPNHY/4JWymhOIEkzUv
3GOeK2QjRm6kW2roPYFGrQO0j0Rl4Ot9/fbcmxs2ya/OsT9nsIAl4CIFzoQtksNA62ku10z4YQ5V
7NxnYPdebgup2Ij3Z3Q/LHWfo7wPWwm9BVfZV0svyTaPFE4sxtXUYhd7VLlRVy+2PyKZnTBMSIU/
xfxCWCgwQdbdlJ19zqC/ax5uei+iWWbaBOqzWJ7hCrPxBFGrEFCxgJKaHdouxOBS6jBMt/u3adTm
ORqsCelDGAgweuw2FAX2vHh1ofB2WQhxKRwruk1yBnxAngSK/68aOEBC1phYJPT0EgkCNUs4oWHk
SmxndDUZZgFj1GlHjZa1cV/RYSqfiG8Zdf3wuQfMZ2rI1NEfKVU1BQPPXoMeKBBMHIacGaWcOGWO
V+SLeHq6RunRPDPSfU6CzMEekovoM5jLLCMtsw4MbJS8nMAP1uumz+FmPGyKYgK+JsSSb3oTwSly
UsHdVZd7kLyGZ+JRLuSKopYMeeUKYv4riSYPj4F6tc/qpk05e6Xn5GldC9Id+oWxQIit4ReIQTZU
NpLpQwy6JSou8NcC/qZcmburGfgMmHlbSOV93irvhQNnJQ1BbvJBhjEAAV8VghthN+o8vTOvUEIU
3eDukf5c+ALu/b3fn/iuVUlDRWau/FgjmjqNwOgnMVZ37QDpUY4uGaElh91TTz7Y8fE24BxmSZiv
cLYNb43HGfhtRsEpcEAdcTFhWDjCn1shgxbdYc9dQLPqNog0RXlyI736Gk8HiWjReCDQ8nx87sCt
yKqRetmiq4ocrwQHc6ow7nwY6OijRxah+PAxcRFaBf3c/DbBlIqsy6DO6/KIBsiAnXZzeJZ4v1sG
nIV5/1U5kPTn3rOeMmBwKWNdn6J3WIniZjXRnll4MKL9OyJqhBX98lbniYUNHLiBdsX+EOXF1BDR
i+gddBxEiwwEowldNscKpZod0TQPI4TMWAaGDl+qOMNV21kD7wRRIO2VnplMPvdHyjcuU/jBalXA
ocqHGdcnrm0fq73XGh0WvQqVpbr/MXTThfgo8agi8wZ1XNo6gJVq5DMeaZ7lgqAjg4B826Fv+GSc
cLTrKXs6u/t1enAYT7WB6MAK/6t/FhNTUkDDV7wp6OTu9gCzvfoTrPxQcEbdPrxPjxJFgbpQDOkt
Nn/BeGSaabegkVv7BuQl6zg5ioO3WSMYWF6bbyNGa/F/qfdYYl8JafYnOsC25e2vM2ffbq+L9NhI
yzEbkBCCTObuLhrOztwclA54jawAJhjavlisrnV5Mv216wEY9dPuFTjdOlPqRzeahqRlhMobBXze
Jdye1kAePvDe14zBvkJwwATJ4cGjzKCsxqZbdAwtwxFQKiZNY2zplxO8GoGIWRRYsZs/4AKfB1Le
YhmR47VuGD0VyrZgrgGVakSpRQ1EiNsKVU4Rk+f1HE3kyzSeR7Spggn3f0hGXp43DuRqOpW+fLCD
bhlRej4E5SoCDtkiYLB5rIIBhEXReKaxCnQ6JbLrHD108euUZeFw2IgE3bqajBYVMmU/zyjli3io
IQV45FlUoau2rmkADMnw6E9AQvOL/AJCzTxnWXm0Bm24ySwJoJjVf3BTXQBtDQxQMk/22naCc71d
hG+NRgJXdJa0SY3QQN+3nZ3gFwr03QQZMsc1cubv0Ec1js+tJXoljBDsZvwdKQyv0RL18/RU0Z7k
YUghL3Wf6da2H2uLvHlqxxWs8nUy6nIlCj49x3xVYbQR4DPDeQXO1NttcHD9gzdo3ciJ8iDiDlS1
Djmu0vTiSLGcPRnjduqpEbpgJ3JRnUfOpSx94yyGmj9wXD70pVbfc/2qig3OmtkqXIppUbHorTNy
gor6BmZWps+OrI4NnMw0kvsgO0xbBteHLle3HQbq3JqpdtwHnxYYQ7v94rhJQuE34HtZ4tsMajuy
/H/CKT9hv7VXaB7AUE6vUawb2vq1xy7Y9U+i35lwClRmAOwaBhb4TmZYCZf4dZgRRg/B1f0iHsC9
kFEVmimgrmTT+g32RGecKW2+XCz1Hwp//2jIBE2fpv/VYKU4B3MAA8IQaMlJPaX6HtaCICzcxGoP
TtnR1+LBvHQadsj0W7FobayRrj2k8L3ACHyV9TFOO0DwbLCSYz5X7P08zuILA7WLkwM+RymCNFii
EvuipqfK7x9b8qKqUMpT58GaYD1pl5LMVigeH8ZrbiO/t0EgizMP+unJGJdiidyLvLFM2S0FkhEf
lT8YQb/cR7qUciE8PLoUQCsjUul+LR+DbEZer85naKTIGDyygaEOdD9gtbv0Gj/Bg9yVRgW7qGbC
lS+olnxq1VhiRtoYPeMX/Pw7BTGy70Env/E8r7Z6VsEeqV1CjNdt+lvxpQG/zY43qJObngIBGplp
B39ntSqKCav1j2i1GHQeTwmXwsn8UZO5NULbHaxspV4tfwMC0tVD19UOdp+dK07TEkwyXHvuT8KI
ckHqsL0i0KS19tRG0up8XwbNc+srlhtpcHV1AyusnAKPR5M7n2N8aCWc8K/TzP4RWcO5uvK26JJp
njaC3fabPEugtzyP+hxEvENwXm2kOASPn8gnqjLykN4RkSlE3Ylkkxhoc3I3C5E5wGbNZGHkqOpJ
Fil3hg7uQD6vQhQRYNCBEGaJww/2rl7Jm7N2CoO6iAyynUASN8rJ0QjROK1W9dxBZDRHh941RqA2
p8NmuqbtIn5Tb709Zg5CS+QPxDLde4RTLH4FqnNxSvWe8Ic6drzJvDNP/hdf4cwP/IgOsIb/Lis8
O6gPK/T5dn5wn7kNWy4o4bRdKotEDtdZotXpk2HJcc3+uXThyYSWTwAuifOoyPaUu6I+XDAmQm8N
eblFAUoc84zQZEz3Sj2gXPFhkzLbGFiJIFSvQwA74xrMatqcJNcvgIHZlXZS8HdC157Cd93806l3
+7pmq3C5DYh0GLDqwdV5XK5uSNaUa/dCjr/s5+ygjYq1DgH/DeZ04u3en0RmE+C+EFGHZCvrHT9E
Eg1AphD9foOs88wWTJz8pjpmpH7TDSzrqL8O+71AD8k5JGp8/pxqz5btZbuBFpG+FbCy7N6ef9Tu
proo7aM51SKyyDDZJs+rMaldqFQysfUh4XMPsXMRoaFrzIzlvAYKX+mXjHLTJUKqJ+Q7S9Yyr7Tf
iZIa6BDTi1nJO2eYpzGbzEdA33fVvgsMduotx8g3U0qWgqEzU7btvJfF+YPHRHqv0E69KET9ON6a
GcIOaXZQktPhes3a6fMA6tamnbvPJmpghfaodIOWaxExEPx7NjUviqsHJlqlecjZz0p/tNhIbAYc
o6iEqyNumm+9TNOh4TBp+z5Z2bUn4LlXdfTY3zGGqX2XhxBBIWVRbRNkEXSnwmDVUJv4u7wA0fAY
PrtjZHW20+fVlbShhCHrQdah3LbFbx2I0DBF/e34/IXETv2EBuBZxCpX04QZTslWiXjQo0Tc7ccA
luqMiByTIyVHXx4+WVzs++kgqsR3plk6o0OAYhfJ12iOfEuno7GgnNIeqBF0okpBMnm7y4Bn00FW
fOsuF0pVXLJEfYSC3UcdXAz/ZLBDRxPO4fG9knl1qWyOFP7FcToSDgR3Zp+tG6Glt7ijpVMkIF6T
p8y770Wnbg8rdqxd/Gqh/aRaOpqU+JdF3hVpZSpLYDLYvFjpHKCk77VMlfbfZpKIebrk/9Jy8BcA
onJsbM7QnXW5Gf61CDG+Ci3dLOoZyBjOqm/ogGg7orwYS5HnoR+3mGIzhokfEo9zoVW+sRn7li9J
zNQE5r4la+e5j3CB+hY6biEKSw9aiV8GnWOvTFZTk0cTYVPmzAXwHfKo3+24WZP8mSM4zCqLFBHP
3eVF9xdE+QtRuZvl0keLjGoe9ba9UzHN0Dz0GOxHxUi58kh5tg7nCkqlmqw7hY7bYjP+qsxXUTLj
T+V/1dglR+lqK011UWAsO3HCxyAFW3rudjwaxbe98erVJDEGMBeMZEzo2DbJmbh5cyGkrzBIGA1M
kAyzfYKobcKOjesw7bt5nL/yL/MdcZn/18Xyy79Ksb3AAAcTTKw4ewOzV92DXqH1oEka2HzraJWg
o4Q8nxytaW/PzT/rb5y88TnQS6Akluk5mLEUGRSGXf4GKAyCWPiT/aHxohmbNxqrBHGtl1/abRMP
RbMupRIwW1x66M9EFzLcyFNuvTCd4/srtemFt5uJiowFWa8Mt/WSaOOIwixXDziZ0IAwbrMz97/g
3v6MZ4vyirAieVpJXLIa9PjXtH4FZSDisKTzMATQ9463IC2fYh20FTUTvwEAEB3GarmWMidWyIg4
hfS9+vDYp0RIj5+j/cnoF3xq2pnOIYuQS8U8bgpDVUitz6nMmsDcrmnNxFBpnKKbmUEzJ8c8OGOy
MKyfI6hU+1/jqHFf1QcISQelYPrX/HzeksU+s+oGwDmJmNlp8kIXUCvX6MFH+NJLjUxFuxbAmMsF
a8cl56wbp9VsXgj3d3ZDqgW1uKaqju5Het5GqQ4e46/9W0WVMnB/0bRAwMgwySXwXX7zEYMer9iB
EuHoKmKIiHjYwbCcAEmnka3/Vw2RzpL3+uCd8GMQ3FG7btNr7qs7HoBUeEvVl+BsNJ6Hv/T50wsg
Qudy2CT1Fz631P6FAxzqnhHthSy2hf+ynDhsQ3S8dJaqQQJckrdpqsvMuUZgH+9ze1VnldkJ9v0j
C93rtI41QTXZolRB35rLg8oln/f74ZQScpHnfvFUfytp8XBlpwHB/kPz7hQzwIW4FeuPFBeJFpgV
MzOPqj/0L4jH0mBWoq8s7TidTOU+eM7ld1di8E40EvToF2jsGpXTDSCf9eHDPYC4IPxpM5rtTwcz
qct8Vxo4mKXgaiZoVWmIBtYXFrzn3b0268a9oUbw0w2PGVQeMsjV1kSR4WeRd+oDqDzVdcgvz9OT
yzBQ7M6Fa6RSGf4IPGsbCpsnPEC4dky5vRKChzLSEUOBc2s0ghpVzK+t2j+TDevfn0QNRKJiYaBb
DPsH3BELuh+y1C8amyzrj7iIYJthHT42AZ3CScTniAQMrxA3p2RaeU5UA1XXXbHeQYnD6uJPw1lI
heNqFFAU11BZpZq4d+XnDqP0Y8e7r+Alxn70uXQI1Z5bCMIvAhAKVFpC+bCo+2sCVKEvLNUAMora
MwgdFI1hwPE3KGXs/GfjXMUzYWeiWBhhZp8EnqSV0dJku1Fb97dgNS3ArS3Ply681z9Ey0hcFr4Y
AIQTDQU7Wm7sjnk2m49IT7VwZOBcpms5mJuSU2uBUqb0CrhtbsvDTORC1BNfGt+8wJbeQMzilb1I
oQa7tizijXqtCaDVCCJOD6HKNVQizUexfyKucUtl8FA851ew9oh9Lu0QxLbqQOzTdW/by9MrYg6F
N19O6I0iIMVhIMrcUgSWxqswGrqwDCLSOjzGabFzEoeffp2Mt8A3JARTHt+slTKp1GntiwWHUX0C
u9+eCgHtbEuYVbAXmXRaFXtSWOR1irl6e1SX+koGAnJ/+3bVvckqmCn+X5ZEhqg3tnb1PoOTTMp+
S7caWd/ok631hhR0DbRRCkyJr9FvDHq6tJCpjCv8VMsVCOuZ1aMXlw3kyNn7/4+6tZdDR/9KyLvd
2uAIhk1LDOs5/YTGrNRcOZZ/fU0CT4BlhE0cVnUodvRHIjJUeONEcohxTsi1qYaIptZV8ALwm7Pn
f4Rt0N5c0E0sBE6g5n6fJg2mkYLU+JI5s2yYrL99yjZVBIvv6E9/mPeDdBDSnlmSFMQ85EwdRzyw
DVsW0jKFF9x34DBMLdVitfJNlEkJKg41xQhDsg0OcwBGe2rvVFKnHLTDAi8odrjK/ae6CSWrJqPv
a+JNrzLMfii2uyl7WvesDuMQBv4BTGKejojbnHIfOAEi4Ph011t/fbbUxxHCEE6zIky4rbxuk/Yp
L/+Oho7x+1Rl8HKSKQQ/Q+kYTm5jCIu/Zc8Llsftar15PqVdpNSrhelOnxf7abyEMkrG/jgkanqD
wXJaeRo1lHXiqGwHIbhAqOOd4kG8e7bLy/oSasoLK0y+Z3XAhSl9EJb/pQGQVrasLpPSShx+L/1O
L7lydC+DpRDEz//5SOuctd4uFy5lqpBipgRGeu7Y7GugYiu9hYkfhogJcfmeAn9gVODdh0jLMtKN
dy31R1L9rGO5/MPJvx5l072eCjFifpuTNZvfMaHg/xraANOcXsDXGTuJYY2XytBfzZXsrS+ehA0R
QozD01SCwQXydO13/kobQmXVu5E2RpJM5i+BGFoU2snr+S0AJWg+8OtfA4SBqY9aUTofubjEHVbv
qO/AAXAdy99YIJXk0aiUdbBMf89TFenStahrnc1Mn2FDDIpzmz1uv31Uc8Fd41SDQ2Y+hJIQ5+dU
VYbglsQcPRI/iEo3tTfmRpLKDiJVlKexi0rkApuMZIDCXwwrABiqR6b1Q8EoDgejf/7j5WFtgHNK
qjeR9gw60t5LldvErn9evByZYX2ouCB3OBqg/cVw1nB5/IlyPDAgMoNtVn8alRLkUdadf1v2edhg
YAF882M/Vxufs+ahapqWPZfMRovW7iBl4TBsNFBn+K3phyk0C5HxH4kzEOf59EJf41rxPD2l31u2
0eye5+rY30UsaqwB8NpHryueIOqotFwILaxYyC7UL5VxdIlKFQaCcW7zGRO/p7Sh53fvSSkY8JFA
IcY8Tfuloovi3VpqowgsMQCZ+iaOEuTFIHVfbxYtlzj7OHsB4R15WfJbDD4NudT2KuRF4ALRO7rS
h66xBqiqGpidBH+nHy22Atk8pdG5DHYrws7k684L+sOA2OhYMah4E5TCxpq/TNss0KUGOWC5MOAv
HS7YZk4nVeKA+7SWHX0oSeKNRGackdWGfheSrn5K5xBAbSEj62u+AOxGEhqPTibfocufGUbGg6cq
TANBphUeZREoUgvhvJAoFpoyIVN485qgPW6OQQeYnV75K7x5DOyYHyJ1cyUVne2ocRnJ3m6iIS3I
bbWzK4ilzf6sor8Nt5Iw11IU1DDIuc/Z4kvqBJ9MiBI+nphlBTEUtssUHUDIcjVpEb3+mdpd9Ir4
6ocymRrep44PqsewFgqefGFvTErTLPXM/Gmi3J77OeS7dfRR9mXf8+UKp0eBCIpJun+4mJIEaufn
6iAYsf67h58mXvR5+YbHkMHMQfjEvI//S+FE1vWxxnMe4g1EGN5hJRkQECMxALN7+vj7WqhHpGgA
HEgurrBWSZB2LGmfVs3ZLN4tv86TflI40DB207q6jRaqxV3HXYeOWi4Dp5ndWiVj8MkKx2PKnTYB
wVkNcUPhzjTbKOjPLbZMikAl/zMlHKvrtRI7Mas8frXMfsHAMs5rvGvRrxxZNpE7CbuzND42pTUZ
OKvHDNBETc2Q6QCZiu6dUG5fow103HwKc7px4rj/PhCgNbS0jQ5Ha8RgA3/hpGJ+c2YIYuB2VddP
sh5pV7QKHG4d1EZ+SdjlgJidmWHsltIk5qrVR9uokRQlWgeyIKLddTC+VHphsKJzll1CxqFhDRwI
kEeCT1WudViQeT88N/bFZSZH/37UF5+iqK6Grx8Mfa+gChdvbABGfyPHR3ppnmJykvO1v+u6vZ9Q
hcMBgG0GQtnrCa7t6RoR3kUw94q2blPQPfAvY9OvelbFUsIeGnFE78b6Qz+AleXZJnwgc3YaKtkl
9AkNAgC+R/76zL2gSP0333yjI7Vz/w4gVertVqCf0Lka5x9wKBqedlKrlLS0i/ovA6g5cJV6JXe/
/JlSuuxr8ziIkmTzwbkomFvz32FXugp9D+Ci1j6jxR0ozHEJEFwB86PKTXN59tRVIJZ0CXMjGZjO
W3dFzSkcyVHo3TqCr7kDPj3Bp4Ocsmxkywc4sXk5NmH0bl4NZKrZZmknMc7gj+wT0J91Ar40Ijp7
/bC9jWO8jwqhc/q3QHmz6GlrqfbvqkvKkwNhu2H6fuZf1aYCI5BRU1RYUc5Z9Wd33gIdrw+ZBZ8k
aJSnPASKb9uKHvlNOOXBZSJOQjOnWHs3a7XuoOmRsO9mD2WwQkAOS/sdCZwr7tD+DKDOdfu2Za9s
7EufX9eVlDNkFgwL6SeEd6msQ64YoHfaNKKFie/2SCXyETPkNFA5Bd/a7SNOf0S4DeB1/4J8LhUB
a4BV//zfu3EaNQ0AGZP0FxTM4fNlbU8rZHfSDfsNUcdORoe9EK673VAqt9XN84JcN5Fn0pkgIYbH
86ifM6yS8Q8QuVP0u/GxVWc6MzMeuFsNhD7AqaSiH/HvMuiHLr2rVQVunqpWCKH9mnjMpYQ0bYkB
6qUMKSF8HVqPEfR+r1IvqW7iUTdN567U5mcfSJdGQKlUgpATLhmkQefInPo5II7I1E1LLrmOc3ot
ABWHqtsh6J5fw5gH8fqAxt56B3fDkWBCPHIRWfBtfnomGK4l7Domkf84CTvlvN4O8X3AHVsuI7gy
dwd+soyMMwFr8n8+/t+ImIZYdz3XL1coqeywsjFk/ybnxGe3iK2pckG/WUZchMcgzjuiyJHQ0RMd
9uhoYfDJkHqKoUeQmDyBIzbbBG3htBl0Sw54IrxLAWDZDW8M1DhhlapRnOaUbkh9FKzuzRKP7J6l
4++/wg3Z/MsB44tlWlLifPVolR/xufacwMX4HC6nNAIZu3xkNYV4/Awss5GBydqGkblPepafjlc7
96p3U5TTrgeOWjFvz2HANtfEIxGnyTsZ9uoXvPB0lFAZ6lZEooqtV8uf/Z0qHKnjbMDann9WCaJB
k7GzXNr6/vmiPnkx2VG0XepAKtFG3Gy/o3+gDPXGmIwkQgqslPJt0FxL2Xzj03buytdvN5PXFKAX
IjO+NqaVy4SoiZNn9OOyAsF6H4CFVXAvPngAbbtnCbIlQiZEtZq/wvTGoIVtKFaOCcTjl8yk7rEe
5LdQS4/G+uXBlElQHEci4bs7tnHTdYEL/dY7uIc1X+ZJgaalFPdRjI7mTCXPhg6EJ1ITNGGZsO87
Qk+pL7yOzZm3f4+Vpzpux1jpxEJ4Jg2K8t4oE7MpZMUabl+JGyxXlvf7BvVRBHFSNJXDw2Lh3krO
a+ZVZaNgyOkViDzpHlr5TmQE1POwEsKbs2viTla+9TQcXjpWv4iN9PzAzzeN09qgMb7aOTw7FPhV
05QNocMhnmhai0Ifi8B/zfA9MvLt8diIQsewrajBHyf3nw7PNLag4pr31YEks06rnZSbvDL4rE4x
2CaoqlGWr9FCRuuD7Kd6EXJS+3RibOSq6pj08ebBbOT2ctfljzFaxKbHP0+IRmEFtaxnkwZIE3g7
3RJUevIL+3d/ZiN5MnGpdCU9Scq0ibv0jwkNlYVAuSP+wQXKi0ZySbwbnj1lX4gSDWdYaTV+oEtn
vgjb2dBkLAhEs3wurfLF0TwW/7vkJjii/5YeYwgvxDVLaDfkXYzHSuxT5nnZuCbznHBV60WiNa6o
0U8AQVd92/dml74nZR5/WkgwmZ9y2XzPg8LJ1GJjCyR+I74m7VbAz9qGp3bC2TxUCImn6FB1DRwZ
GvEpCQoIOHhXu2u1QSQIsGRNPGDV9ZCgPGnRX6xspJO5TKbhcr/nv//EgzOhEiN37l8qewAp+2J2
HOTRuDToJ8EYkKFuN+pyKD7wH9zuobsFzjoLKQLGM9LtoGSdytR1m1WF/IhT31isRkclvAB1UzWW
W+SRHAeN0r0m/13nv0aSp2lB76ngZri2d+4lR/H93RmS9JoSWwyVl+2QmaEKyyC2esdRTzhwvWAw
QnWbwWZcsom+oFCXpEPURwz6jz2bF9QsePWi1yBKQ/HmoSsyVb6LEJ6ya/NXywCHOp0Y8gzc10Ug
AwuNJ1EHWXFTE5neRMuvnA+Ya9AfO5DpqhqniJaUOq6wfBw19WPRR5yJNcyL17r16QTmbSKprHUc
6OLtRhUz/tXkVpcBNxg1a7TXC+W1Ly7MgsseVhD1jSqutW+L0tJav2x7XKMtOyGcXYCdePMXr2gA
F2lYOSv4jklvf11AhbZQKJ5NolEG9qtBKgnHedTlvvMtediVebCQriuoD/y4cWgWaSbgucBvYk+E
SBX7iYN4IyDpx8psc5+mKq0Zg1VRs2badCGGTy2BVcOib+P6bJ72a1ufCLpmdmBwTyB8o/Nwncaj
kHEDPJnMdAWZmQoZECq0n2MFSjJYJjK/JOdba5FOKDaVew6gpqdEr0jV5qWHpk8X5xmcM+ZFT3zA
+64R+46gnnWSKKRCBpx0kMuV+S7tvcFztBbGf72HYzhFabu5Lwu0nzgWOJrP1ZNtk/tXuiyFzgoe
cLRSsWUrgkoAAjTYDDMmN0O6pBIjxt5P7YbaEtFRUdD/SY0AapEmkBEO86Ik4EtkdbTAD0dZYO+A
g8Oca6GLnRs2Y3LaH0/aB4slvg05XI0r+83z+RVwWOiYa9JDIA5dP+6W+o10yhHtpVwZCQspiuZ1
uDgu7DolLSByR9GnabVHdjI9adrWT3Jh8Em9u/jOh2TlDx2ZZxiPkLckej6sHBHdIDMPfo1C3esj
+2XwJt/+uOGw432XVppV6xKdIEql/+U4pwyHdfr6phFUW0NpwVrsqY/UlOOTPTVZeJh7Nf7H5KLp
KWcs6jkmd+Eb26RJUCjVkH9iwLDL73a9EsPomBSB0ZA/00Qm0QuUOR6bVX+B6r/Euri4RtiMyEae
OXlNh9MtSsEOUWQ+j8ChXQaUGvnfn3raHSFQNDluTGofpoFgNRWAbAo/nT+svKoBKEeYpV+8PlPJ
AtIuu47M9u6yFYpZFlI5weJtFKFrHZNQwEp7wJk2esfz4gn7ckcqnkT+79zbFJYXqGSCPnRz7O3F
elGfSZC1+yYmEdZQu/Uou3VSq+TFclmwvsZgAZA86xnZ4hEinIu2rdwvucyCuRHDNFp4AJCX+aEY
8ztT93WyE1oi3HxpDzRqFi59/GxEY1D3efDOHUb2t3LPPes2iRHow2Ndq2IjFHbSMkbUSKrfQ5HU
072oENkUFaFBt1pNE43vLLyrDl2w7y2aGNxq3ArTT+ZkL6U/rwFk7OUk/JeZv3o1l1So6zSHiO54
n9AITlipvJLj4cg/BAsj/lEW9HYgqz/ksGYN9td8G383dFhz1zfnCZd9wmfWGJWUFog22LphDups
iRibxpFPyqkcp0zf66mJgEVqXdNUdjcnOgm3/5AKvWBT9itfTRtN96L+wDYJEikEeUbWPTfXOSKU
LBMvufwG0VRF8ud6OI0DJjL+o1m6Vboa70DWW58jXZspZHu20kJgWf7T0HEZLCNVYNoKQBnEfNy0
VUiMNWfXPFg5/zTcgUF5ZmfDx4KplkSmkOhly93XEKpKfmhweGdwEYvEZurTCKjVzPRIEjYu3STa
gr9UndhZGvqg6bWCe+DdaoQzhPKJLcsCu908GK+2jXLvJ2FErideZcCJ1mOkzzHjR6hNvxonPLxY
0D3wnDTm0WHZMawG9Unphq2Qjyf2FlM+/994HptK+LKVb5JUXzkacbHuWoYkUuK6CYsjzussA3+u
xCdX5PWLf8Q3IrwCDJq3RkDVUAztvobzDOKO6c+wSYGDGuUmM/nRRTeroKagE0XfEf40Q3vlgSz1
pvUMBdn7lWjE1odmJIge7OYBZI0pJemAOOkVHYHkTeu56fvUvsVv+tJN/M02+1N2EwdeJkzwsecx
JhWyLAW6RNSer8LR1Afrfw9+EeCOlR36ASKBtx+e/3BgUVuu8if0uVicamMivvX1Avg7ccMidqt0
eylBCzyO4ou329f5RHZczhzOEbXhL9DTw0WSMLgYy8/a18+f2kimgCLdSGCM9r5qlKbic+sBgwcO
XpFjybNrAfb/7EgbV2oBXXnETE5JaEy2AtWDPDwI5B+JZtCm9Tb+jTHqn8K/CaCO9PbSo67wY09e
fKH46coNjz7/YGBkYdzkjmBG5fgXQmoivwazrwl3w4Jd92sSl2cBnr+HnB28O8RuDT+tMqNbz2y8
WzwiqB7+KYPwj7mBCllRnZCt0rsJt/4J78cLeZZUwCImbIrE+LaMg/0Jltx4wQzvdAFCKLa2l4sj
ubWmzbFaxuRW0wz6H9VvQPy5Yu5/AiWBsVYxO6Bu7ZjomJtoEP75RchNaevmZ9LuxyjhsIFUKCIV
4uOc3LANUzV1123w60RKvG98C2wUCGEhacs8i+u/j1xNBpGwAtsMGjESAsuGqu25UzcUAzbbI3iK
Eh0r1SDG+alDIyF0/FRYokW7fAFxInacXge/wmT39BDpVePS8jPlEu17hfy6brW3y1bgiRGL0j92
UzaS1sUVQdnY3SPfhLhbWa4c7+Yl984C/F8lLn207tK7QMAphOtuJJOyD9cHSERVY7brXWcxPFyk
yZ4ZRL4zzubuw/Vxx6twaAzWD0k7oXpai2wi8ZM81YjNKn+GUuSBV9eLxz/azZNEw3eF9DkvCoc0
uN+YUSEw0GuKm1jBPhXi3qLkrsMAtXxlmm1UWHOXAJHdcv93ki65FymHY/yMhn+AQ2y/nHIC4tBZ
JixDtsmG01BMxIexVXkFQWLgwXAll1CDB3DERvxbaFOa/VRIVjfZx0Fyjyy6Pntntqj7DWnE9FmI
LZmn8E3GwAOKnOeV4ug2+nhty27p95kjr4+PlYEAMUItHpQVFHVBhms6wHiYPNOpdd3KAYfnFT8a
kVe8WOTmTonaD9tq10HQPlFBq2J31MzqXdHsSuMl+mCHBEI0Yvq81Qq2T7bHeg1m2KaBVrBzS6Fl
1sUdlsp6riNfinzunTgiowns19gq4gOLv8CbPKbqHBJVRkVslRRdWoWwBlRF9zurG4wSbYuNpsFW
bVS5djUuUSWM8RY8HEfs3i4JyANXi89TAjhSUe6mOCC6/9jkxLm7Su03yvH1Z17lUa588gxFX5Xh
qjEmj9APTfmkXrO85+AmPqDLtcA2Gj4sNwo4FBRq1o13negiYlDS7rLrt1Rrsdgt06dCeNVL0C1N
RpFp4pOl4ferdCUyXRfhttWgWZ34roUX06OJRHlX/j/eVZkJxMSJkB8ZeeGxri5b4STGmGW8zlSM
xAaeUUxlcH+P4UNjZRCZ/JY+jfBd07Rl3XFOU85C4D4vvjFDOSJ9OngJDIegOhqFdkZaXZbcNl4k
y5BU/UwR12EN7SEPoGdYc2dedHYUExBmCqGRt87jes9fppC8jQ6/I8kcoKXUAxJF8vcijfUD4I5L
C8NGPzw2RbbWflivNRrfy1T3VVhHcDwzIpXmMeehQsDmXqeLU2yFulGSzJuEH/wGeoRm6/FD44gl
2ff8h3wsyCaPtwQ3ArOcV0bx7f1qQA43vyxVBPzE64fclOfqd1oaSDFPsyaCAh378LLF+ddOMqpB
dtAMvqauNgXn62tWrLs2zr90oYoGFLH7mU9zp8/1qDu6ltKDNcq8/5KXxX007aA51wJC080nZedr
5REfQ8jvTdaQ4DhziU/+yH/3/KhoAoOG9BvU8u5MD7BoiVFsUxE4SEM6DFU2bSBVlnwJefuDIBE4
5xvHyge4C16m2o7oX8iYH13wYb7qnTyX5JLO+GRWdHu+kpD+I3m9KJNpOV4b8wje7WHpOg+Tnam/
EKXM7ArX1S1J4Hcvif00Y1FJr057gzSLFzidjh6NQ72AlmT0FRF7q7TZSelCZ0nUl6YXrwiPTIK1
TzvuA59Z9bWFBIuBYsOpwMWYjt+IDnHNAa7i+r1iRshwQezMaz0tousr0DwDGSDixY9WoAx6Xf7D
HdNjjM/Eu2lVtPgWcJo5TGxKU1UiIz3n7fu8CPXhqMMA/X9DOQ7rdOYK9lbwooQoqoU0cd9YrDps
ORHC8aDjYFUOyBg/SoWXjZjcYROTNb09FkIJsA6ucDo6OI9Q8Sl1XdnZeDVTkgkf2J3ZANROk6VO
KxP19TwOLGFjoI11yF3FHhb8Hrm1fYn8WlKCSoV+HFKJKt+RRYMkXYHroMpJloCVubjILKhYXTCn
X09z4A+8TlGMzrWxLO8YeP32m8PNF7Ti/eCx7UZOMmNP4MNQGJPbOER8hEsDt/fDaqdaTbDKcgCG
DMHzNerJwAw3Cu43jw0QkQDDuD8k0yBUmTI583/e0HrjXgGf6WuUnYOTSK522IO0+k82bHDiU5B0
fizev6/xKQ/SgueqHx5h8t2TCu4c3/12+rZQY4t1u5VqEGbYvXSd7ai/vnU1yeXdxgF1xC8weN2+
bUPoL6BOiTB3BGsu9ykhji4z740MqSRsNsif7/qDdEoIj7FWla2I39WYNG4vcNJKoI/xkDk2BLJl
TDgVKL6Mc35bsxMhQrzKC/ma9Tmbx5bvRL2mtFhjYVIC1GR0XmFgMpR03Y0o18mIpyyBqhAl3LSN
JNvCNkrAHD1ksx12rJe2s/OT3w0P+sXC5fOfj4e3Ts7dEnkHnsszVWICBT61KNZ5w1jre6Cf2SsW
j7/ox0D2G2dc5Nw6KuhTnn9GMTm4hXe0S7c7JDfv9DzXStghSlNe2nMr7Ffm8+LGg/i20X8sozRI
LiSOjPJgU8IXTduj5UDi/Abp4JpI1vYRw7RcjdnAy0m7BP2Qygl8gD3Majd7siu/T2ZXg8DxN9Ay
BsqbUpnvWcW+2zztN632h3BtOGygFbdByhKGHrfBLEOSGYdfFNlKgWhLCCwUXR7NKvttHqrpG27M
Je0e7qg0dbVZ3zUyMY3I/Hjmf4ZTeIQqVZDtbedOqPx99z6OLtxK9oqWXOvCTFbx39/oxOdeIpqq
uMuQ3AdJKWdpxQdOXSKabgvpQvWu4FiRJDBclPN9hyNQ5ZY/3Mev+eySyGlTD7e1FW+Uu7A5R4mv
j3g0QqVch3cPLJlAQnUhCSjQME5CViV5wBg2wvy6IdCsNytkfizgvV6x1aDDKdVYjcIJ3DBx0qeO
xp4DlC2V/z112prQYyidvNHwKVD1htnY4lsOtzTEsxirjUf6Kskm45bp05T4f3eJjQdTRDpEGg2R
SExBc9LEMa/hzTTMwWaN9fAeDVdd9aAdE+BZKVTvXjE7TvrBDvJwaZr45ECkp2p3lNTJA1j7YN56
xtNinowVr+RTmsW0Um54tQkyaRkDj6i4Lvp/fE+S9qJtXP/lf4N6vpEk1SVrR6AxRZFmUT/PBthJ
J9pCrAHYaNR1eYCQFZnKzmOK52AOJTjUjGM9/N9M6/wWioMc+2BwOHuLBIN9nFCGG1y+NwgEFkXN
xXg/wvD7YbgmExSqykvq+MVdCkz8Htnew5fxnCQ3d2KaTuPE9/fu9IAaLr/AnVUAJQks88HHGEah
NhUz9nTYEZod/mXMiP07EfBBukIG5sfBxbK1hvVGkfvWxgtMGHLEGIPHctuDckx6Sg6es6mpp/eo
Qq7C+9HJeMzN+VnQAaTzyhMOYaKPL6AxIGrqUg7nZyIENAw1+AI/8AlO02joNoBM1OjJhWwE/2zC
ZcQwcKGn86hR60jN7jjijMN0ib4Z5RLFrjpoOi8OYonlM+eXHnipdFJL/YTQIe9WTfeplm2nwDbW
DGI5E2RCpEqgNY+XWlI3fk0hUNv8BmN2nXTC8eKgBrxl0ft4O9hBLDZIwKcAyaw4Mw6qAQERlTeY
RVS47HoXVm2UxiggXcZv5zaDU4L3TgQM1spDauS17vI5U9efM6m8rvXDhBGBz2++5NdYu8sHLHYO
xLo0Hubqd6o626tqoyctF+Y3FB8pwa+5flS6WjGgfNKH0GznNRIVoKzHGGiv1w+exyQO3HARvz7N
6FKwr7a4hV/9SFdviDozSndnZ/8V3mc6zXVvRuU4B572uVz2mQY3SKP/VlyhafaVYNy5Gkhs7h0W
G/JKBuo2RAINOiLYrt+ECcd8k+bSe7utvE86LDPtemS95/m5prx5Ujo7xEIDtD7jsF4XUjnoNEVL
h+85SC4dHSKzGLmGTXrUOUk5eT8FTK1x2DmdxnZjQ4RmegumTZ6ohVEk9IGqidY6EdLQwqT1JbL/
d8zmLlXZamT5rLQXKURc6nE7NPmX0w727IyMK1TPAnWDFoAMkhUStR7ng8bG85GgOttGVClFRpaj
w4f5zXErw523K2vU1JiboUlzi7OYeqogz9tNZ+HCh5dG6QDfxR+phElLV6Bg/thIVgyE4qFeW0xH
UYIdpmav4wq15p+/DuNjBseKeSXBywNE6Ed+oJpKj0/dEoyX3Jsvg9ZsyAYcSpk9vLQAKhaVyFg6
bzb7/XIDdGFyAfDLitXn9TslUW8hArYBG/9CBU9hE7jLajp0wFrASQuANt+XCIkXx+oR0fVmA3H3
rTByOfPpU6bhpdsv+/QYbYJNdTaaioizgSHK1bNPAT5ebMKVikkjxYMQzMv+aIZ4eS/5dmSgWy55
xPr2w5agmVRBR5vnNI2+WSkXlZtJDyN74OHw3vJzhNt2h4rNZS0yp2U5vVtT82Im4xQCjOTQBGgu
byVctrXxRbduxig7hGgloBcJXW8mbNRukEQv7sH28P0p4MytUufK5R1ZqaTkbiEeQe4TqX+E2EcP
QAhC2SpH0HffnMAaaQ7KeUmCHe/jUonavm4shhExewl13u/m1TWLX2LshAsZuA1MEfBs/n9n8nA1
Z2oz5n6tucbLQKtxoelwnQQsmFkE4qlu/tEUBwN1oPzEzAQ+Ch4tw39dwqkktmBgA4IorM7zb8Y7
aGhkpC4a5VdN2zdx+NWGCs+rcFhyIFVXbfdsHwL5iOEBeA0Wyidt9KHpXJQf5fghKi4ehQv5S/Ep
jc4/IdFHp2Bmgn2rU+n/QQmGeE5TVh6nVM88w2CDh6PJo+O2zyPrAoowpb/btBCQlWi02QtuthYa
gVLNpQ6+6VMteoy7RE7WlNJniL5vPcxfdOKuG4Fj1JSUq30z+o//qdz/rkRLadbMKTDX4RMcxrEQ
3WnsY8Vn7Q21TwcfaJ/UFI8SVMVtBFcsDwsYbPXBU7TsiFOQfyY1D6TRhzx+BZgayFvasfIaBwOW
6AV+4w8P6m0y1JHJ7XWjGM4suyWXZNPYqV/k7ac9BaW6hJkKzfI9ZcNFK9QGF9y7yFBWKxDmhi71
wJZ1+CdIIAXCWrTa98q6z4aAf0DejbQpDnqkfdsx9tbE2T6hJGTKCNvSs9fTAHI/7lOYDCFjxxHa
Mi+eaeHZgfq6ZiiDrEmND6ybDXcSg+oqhUAp8D/OGN/JwvSZhxp6UdOtssuIQ+ejrofxCyG4DZQT
m2yJbjMTLX65JKivrrMli6/cmX/6bVB0EHfBLi/6oSBHVM5pW2rvex1586SJ6WW2oj9VKTOp6n7L
wQNO+1OKxde/382DQQoNsVynmatEPshxGqlh9ScEU9JvteM1mUQPFD0qC1hLSu2SCrFBv/dC7wm6
mc4ihEVCiAF9yqSVgJsE7HGvHk4PrNSU2I+g2l2Pa84fpiyyc8rhtEHKCODAzdReJZrlEBgiRtrN
2etmRYGwWj0hzqWPqYOjitcByrpVd4u/q28JIekY+2eDyksnOfOtOewUAfXExpqem4oqJarazCAE
IcgR0l7jy6JgpXGAR4u3yOx3k1BQDGJMU758cKKaH6yeWjFGHq2U+djHnvy/nv6M9bCPz45OKc+d
ahTgALSZKaDGubTSfpb2Bw9GOhzfKAdc9Fz/jpM16VSJRXEXhqeO7m1oBPSVvdyTM1e1MGPzU1l4
WOsYd8KGuiiuFJvQgYFjiDOaA0EkJwiT/xzDSLby2V/oqAzX0ghL176R5nlJ7LhHD8sjwMAGdu9I
yVIXoC63tc3oGEJHWMF9sPCa6OlRCEcpgqEgymjLhi4PqQNrV0WByg60c4mrqlwXY7eIn2NfO1Nh
oKubWsuA8Urwwk4m+zVjQ+E+P6tCquP8Q6iaVZUHc/x9971bo5gsYiFXiqmM2sgGqL5vdiisbtCy
ftg9mZCBNWqR1J6zfQc7gz7OoZrCpeAfc+y3Hp/JlRQBiIc8slIEFYS1+wGXHZJLEby2t4ycJ9qW
fSiN7Uw3bxYjvpClAskRNWKb7LKOG5warWawVAmE6JSWbg5cTVUmktCeEF1AUCl6MYfnRN0kv7+x
yxpAzzRvY4JXpjgOd82IZmb8QTxg8QRc3FP0zoZxf8szB/VKzAm3EEnfzhSAVYkvuuS2CCCSHVwC
oS2mo/WxW3c7M6YJtNR3KSvDYdAUA/lVVv5yHR0vJf/NROHSwWaQ+G6+9eFyCtsOkWGa5yNiHunk
66XFlgJVNgBFOFtaDhD3mlJBIGZkPN2TzAcgKn4uMerLkr920n6ZS6XIVtqUQJe/Vs8KnUC2RCFo
ZgCuFjNvajrBNbAJ4Hpcff/Bu+7ktI3aMI7MbsDJGRjA5BBTzybYovWxRU2ZaKzgNonFkfBVbawH
f2ZdyQck32jAjq2xpXYKqLnUZh+1qah5ibx3WApQb/o9yUFczcc6/OfrBet2ZAy1eYorQ7+/2Ue0
2J9tz5jhOUg9NnRz5W1g+ad0Ph5wP4Caf7Dmk0bO4n0C0P23cpi8gaY0L6uqV2f10tFyGZlz6jjQ
IOLXC5M+ivUWerlUz2Mk+YbBblfrDAwZfUMaxbVc4FGgAuLdvynybKF5paPk+O31iO9rAJRYva/v
Jwh6v/L0+V9hobPSgMYHfTRgbIwbfzKyY+1XUkwVFEJW7eiqucdPcG49OF+GdHFu4ohGkltvhBbd
R0yIVsoGDQS7YSjPmG5anWTj5x7QW8ZrO3JEAlclkbQcC2Qr4F9Dbq3fc+Rlsm3aCbX2sYJLzfCd
kNcXTERhnqWVnLYyVx0u/uUgjyTfGSkW7pTHg/qQMSM2+Fy0H/CIFukI+zRJh0l8xCJ14JXR314v
a6QQijfU4mH+LZ0NaWMbZmPCLrDBy7Oj22MqZwmIh4OM1VX8HuYUaXDE0cGoba2nHn8WNuHO/MzO
8z1Jb/y9AKd4SFNfm+HYMHuZb+kR6XuHuJvRGJWImLRkZGzJJB2tx5LzGkCfRMJz5M98XPn0ciyx
pFdz5sC+51sCx1xTYZObLcJSWLqC0QIMvIFWlmcsLh8LQTl3Uw7/ybQoZLBZCnmlgS2dXfZiC5uU
gHgTNnCWi5vXAslXu0Gw1AutOXXpy4CI3bQbxl5MYg5SPGzL/pHmLwqBB15stihxQ+MviVuOjGrM
UXcx7GKhKnocHT9lF2n6HP9sA6iRrOso7Zuis7aIrsvp81V/N3T/GydlCQ6F7J+TKrrFYl7zufor
YzOIlyh+JcztnYvBvY/6tSUeQ6NzR2jvt3u8OW6ZRfvuFFHT4Ory7A0xPJHVxJkjNL3J9r1PUQOK
bnwHsDqzPMxbjKD1SNLO0HADHOwM6xK/eAiNiPG3aKuYwv9hXqRLigSTPRyL0eyWNFyDHVwXvAG5
Y9nxNfmGHMPKf6sX7GPJu/BzAZNN8IHmCzIgZSpz1I7+sQatK35VjeXrtXBetMXBjPTk1A5gHAsf
qJIqSLGBZmVYNIIHwoyokgLJCclyEBPt5kX/otT34kZHoFh6qQKX9jbl7B9gZFDpndpIjnR/ZU8L
e0OmIHInIuJdbKWJ++LDASC8tGHQSsIvddEfFVdslC+yNY6Svsoh6HbfZpJVI0LSLLnDKbCn04Sp
G7ZSlAOuUwicbFAkFuudq1G8ZzrYiEEYV2Y2rUKbaaCXDDit4gT5kHDM3xM9kIXblGZAk/QjtfN0
+VO4Z4iexUfu3ClffTNz9SktmL4x5XrxibkR2SNAmlG300k8KnJGKz82jIWEh0PDORAgeqy+l/wW
+61ahf+a2aCFJq0A7aVuSFd176yjbWsaSWsXUURlJuoJFwLCxkAw3MhkV1dWxzkxVVVNAEG9vfTh
Slu8L5R7iLmx/xQdmAp1RY81U5GUbrGP4HNqaEbW3Xz3V6iAomKdNBvhJkqXiPk8RXtgq8INjwDj
1Ut7t8pTFj6+hQRIW2WLXYe3C0Mk9+fzzRZuMBu1D0OhUP0lxTcacqdWM87KsoUMTnwyijAuINwS
wHy/DAWh1DmEUVXxIBe71FEK3ZJqQbGvrCs4dprRZI56sVJjKfe1KHyWLJRj0FSiBFYc7asqMG5l
8M/VuqzAxrigWoJPpDci4Ydm2odEPfRigZ+NVKRsrLWUSnigUdSliQxRZD16L3JVsYnA+bssMezb
+YIUAOz0YL3N7vkAOPWiaBUpvBT/AOg80lA41rHgs3xxprcNilP+5VXP7+7LI8gnPj4Y16lByxIZ
r56PpRPkM7IHR+W2m+9qG+Mf1mpECyEMokQJ1qu/rdGR0ZzqBRXqnFGv6Me4a27YJi3ZxfFmOyr7
Osj1AKAnWZerxRKvWq5zm9Si21MOat4y++iZFAjnKrgAoIlr+hhjJHyGgC3Up4nh5CzkUcerCaQe
O5x44mMQNbNqEL11FQOvlaGZiVae19O0XgjPajJ9rhqnG6f0dGRlcau554D/1hs8EOJqObeY5W1P
/J3z9f6t3/8ODAcxuBtkKPW2QzMSkCbvQ/pmLcGySyzuaHSADScDo9RbrRoazP826Hd9xLn3HJS+
Q3LK4CUFSqP6xXoks4vWbOBu/iVt+XA9I3sdQMVrigyO1APL6OfjYLZ1rTFoGjyvFkv9ygYy6ndx
GGA6bqaKnYRZLct+lcVc2hptR75R73hDpW1OPpfTIDu3xFWLedQMZ0CSA02QjlhGmqih5EN3neAv
omkB4D5c3PFLeSs5WvJbdAFmPoPLhr2fjjusSYc8SK7LBIu4I9M1R19tdW5L86LRghHLK6TUPo66
HC3TqR6Iim3kjBQrBfTDTbB2Cm6LDm2l/ZkvD179OPPF7FT9tMwlRfmk5Q6bDcILDXXBfBPn9z9p
UmeR/NzAtMfMcjw8yv9LhnZ77I56/sAxFPYxcciuxH/SzOYqWsZAz+/MA2erCxWWPLFmSvh5Pet2
KVzkchegSVJKGIKuYByI3JnEQczWL1NdviH/ZsMtAGt5HDCpKyox91arn0jwXMpWR2L16+QCNuW7
vhaWQnnHq6GnH7xSwBw8H/JY0Zjw2fZng5jLVOgM5DW2Rq96b27WnGE5JxbPzxQ8hR1S3XQZf+8t
VktTNIHSevhkm+3N7QF5Jb5UxuAVtOrghub6lKsTg9ylDssI6NdtVW7Bz205WUVAmC2Q44Q2x7HT
lqTUUpdsQL/XLfB3q9/YVexs8+oVV081i71RjbqA1yyLZB4h7DQ8401/m45IXtHyGRhLg9ksbuXK
TO9jj69J7Lsb2fRZmAAwE/iGYsGLmSmFBv/e80UXOoJQSMYrbT96eozJKuiMd5X5eZjBC+PfckUv
jnmuG5xyK4NalwMsGKkCMBCB83gz46M/+maz1Zx/BuAn+er5b0+RSnF22jci+QY+gIDH9/tevKzK
Oy4i9ZulSZfwfwZpmfwUOz51Dqblkk0LSGIutCtTPtG5Qjy6kY5x5iOnVZ689f+iFhWcEusHiZ6A
/biWRTfnO92Zr+EMfHU6Rcz7YW3SHUjEfYuH1rHwddGLIpFnemcCqZR8P+A/VUyiwJjSHkMV4D55
lWawZrkm1S33sbhcuDEtPpUuEBEWwnUlo3JuckZqME7QunLt1fD6feB8yz5IU+zMQr7vcHkM8zFj
fICz9QXBph6z/9F+m914NZRhG31NXvqo5xk87H4Lpb1WI5Opa3Y24bKY+T79GsgT+cH5TeLoh8g2
CnxhJA2Lj0uwZO3RWG3o9SeFqRqTwX9dtQ+NZ++qgwJkX6et6aPeu+yjeCeUgapVqO108lngoXUc
3aD5Cu7PCzwfo2wPd6ydVtSb+30PDFc5fUxuX0TdtfAH3/+EyDDYi6+OQGcaiUahgIESt2FRbayR
Ccf9DsAaIx/iftJ0sUayyJaKLyPmtMFZJghyEnhEblOaRC20PxmzsGulmdqWVzkWrObCSlCtKwXE
a9HEPXFmL1JX7lvAmkYCqPcN6S7lNapIAJ18Xz2pBiQkWBcTGM/AKcTmXzFOJ13ELy6f4t/sggeQ
77blaf1qPK0KdJK0s6e8dQZTh12LCkotFhoTU4U8r75DWLmvqrQzKP3yGB1Mm9wRElowCDUMbKfp
GQtGqm+0kgIuxfNBGDPzJQjwu85mfJMFH14jdbI8J00LxhMohn/nHm4zLtDrnhTNKxClmV5dlcP/
B6P7IoXT7lSHm1Dz5cN+BWXDSEvKBUMjwqB+fWyaH4Cn0Z0jIG97yZtqelszkEjSgy0JsGEaQtvM
CPhBJiY4glhC3Ta2PLm0CiA9kk4MvQG4yym7rHkqZEtd3MK7pg7cirFMw+Grqrp2nhxwC9/gz8Ep
i9BDCcfRfVXHPRdjwIHZe/8XeDZBP+izb9tv10KAn3232MCeGa8UJtpJfTKpek0HYWdN4ZpnY7AO
Yd4I+KqBd7lWoyWHFPSxpBoPhFQepcG64gjKvLo/JBz+0kuIzGjVvBJHbX6lN2Q9TfVsAL+sRVjE
+v72fPMO7KPp49Uf7BviPUSQHfJIyMehBEOx7gQwOe5Dia9UehiVRfFabuUyK+HknK8f6/fgegyx
GjqpetIZSfxn9BHQ2gMCLd0piDwMLkjoq8U9q/DRZ/EZJv3vc5sLDY4nWZBndy8GC1je28G7ohvV
qoYp6PhJbKMLbY3LFGyoMvfQqESL0udNkFjOV2uQ2cT4yFTZ3m4Ua0B3PYuEeESAUO0+NAvwzCjt
YeQ9zou/8NC7iSE6I7SoKqbfmOrAzcMevtIgQkrMFiQW6mHP8Hk19mOhK72RhXMK9XnYD2lNphji
fzov20zHyuTwBLmTibTB85sSn7firS/ph2PI4MI1WyIMcLtChuU0IeUrsQXluawFHixLPs+L6upO
Op0/OHdXtvqF/R/m/2wsl22US1HPvR9tshNKCp2gkDK0BvAgaoJD6GXx0ZAIWCT9D2HpOkR0EWiS
fnGeCoJsV3zZqcjjLI9YtfCpE51kx5utMbA6/To7GTVE8EKO4mVaadbM1wh2zTEhBvdabCA3z17j
eOlNKub88dpeKQUR0VHlI7aMlkSiCVs+hr1HyLrAbwe2rdXKbRTrud4Ddu0NBeyGuoox6HUFAIJr
y4PjbSpsdAMw5+ryMyRKqdmcKf7+i+9JwiO9fLGBKng3sMPvTXN2rW/cde9KZHBj3iH6nUbGNex1
1PCdpcylPq+agmBPpWXKGZl8VxvmnXepPGvoMbXUWuLTBDvb4HXLQgviFd3Cs3ScWtgzTNmajr+t
Jzc3rKNlS3sX0g3irww5RopJ3V++gBEx9U/RHuRYaWHSSF10gNnVZ37Xy37BtxZ2bCLHDI+H7X5+
DMgZ+k/4MgHe4U6uO5Jpa7jW2Z1QKS0YD+TmI+6E+DQTnO1+j5+E8+hLBpWeDGkVIQx/mzjy9Csn
2DPaUwgNh6pqKJIVusIg8Nh6hBZgw76Nq6GJM2BNBTZPrywzJCUAU3m/mpdYwxWYL2fnL0bPJinl
JjA+6dhZPnsEyK2b/gfiycYTbAg14i6KegOL0zPqN/0gt2olj7YkjIWOyq3aJpFap/kZ9KKjHeN/
5f6jUSquesd3ME+z8dBsztf4RKhVmorJcddQMmyi6fqbOkFf1yLPjvvde8b93wf/3I9IP3tpOtyf
KMizsv1jl9QaJcM6tcNM3rRmwuOAZDfZLcy06KuoLunHp5ZhWXG06ke/XOuKzRwOFTXMwNJY2G1W
csWSvHCrfBFBgs2jAYABulN+BE0TzwqW15BYTz7EO0CB7uZtUfCZ+kQ5XEGCD13lAL+lr5jSX8VD
/k4pKmwmmskhBm29FwYlmM50MNqYt7j5GmGBV8rRAt/wcY4mMV9mlABhK5+kcBlmoYzSQ86GGINY
v+cz8z9HYpjRLgPs/Uveg5JHV3kImsrWjln7Rs1I8nVePpetAeOir3jcslaEEj0jRMbyKO5QBURx
yxxWene7TjGC6IaLwKlojrEAgyovaLvA1AtDowij7GDFvkevxybL7gn/GZX7p0ZH/MCo1yt7v+nG
Yvi4o4Crxk36byvV/bSsIeXTnwVUEXnaZIn5gIAlpFx+skFppH0tD7lzTXExrVIcoj/cS5inuwXf
GyElaj9gYiwiQXutHGy9Q7WUTNKxJl2mFY3x+j9S2Ki9FE/4FoHOZQ/OXXqqj+CTi1hTQRpF8Jdl
68IUAfXlmKijdbap+Q1VE0DiYiaxOMxbX+sqD+++cxY3N8qZ4UtcVryyhU2+BQURkHCmHRPcv2bJ
pSw3bUZET7mBkJqHqiHlUDJuQKuH7QlfVMPTbXKWdKeGtrPM7pBa0Xy7suTnalozmsFg6eZEnebA
gU2s1Ob0iXQNrwnIos8dWi5R+1lnC29V5CVYRoM0JgYOJuuWHNma9y9/DTU7gh04RoT32JW/rTwg
5L0GqX/Wv2jPccWuVV6pFtT6KZSkAi+67aRAXMfhHgRJq9wGhRVs+4uBE5M9z21tGhLGQZgKsPKl
/7mNkGG2EKXyqi2q4o/mTNQY+xZQvGm88vg/5vGjkWpG6DPomQXY2+iE1+qoqkgzhmpe4qfqNIVH
OkFf+JqvCp5GK0K4Nm2hQIfan0/9+Q2SHqVj6HRUXLeyG47ycyP4N++dg98NXbN9r5VAfBaRQv/P
kE88FG4YS+H76x8+ha1khP8X9sAgZnYrzUrblkGbS6XCFtlqNyMiVUavU6M8Hypl39inZTxtkpnB
UDSEs4CW30UwwRbKmK5mUqqp5C3b+5qYftRP3WWR9nLjX9u19TmQkkxd5iF/5y6Dcuo2xVW0vfbW
juVXC6MhcMhhdh6hFpLvMIwRVzQXPt6LfDvqNJ/pFEZMUgcDSyuUt/pjOqGZkDYZgzbHAb6UAzS9
9frS/RrhNMux2V5RxOJppIj10Iic0ATz6lC1A0iVpep0bBrKDPz0JEhhNOfOpp37APCFHQv1okiu
fHo9fX4UoYy1FVd0BbCz4Qel5jpgjoCfHLxhXO22L6lS7pmCP0pkYymNLlK8nt72bndLgLo6j1Cc
VdjxhBK6+2rs3hSiNHuVmF5VSgGtIQl1bs/pVxDH4CZbPuAReXbXurBFbbgsfONs7Sefu2SdqGqz
SolpyxL9N3VSB7h8GRHg+e1x4s3BqZ2Sl+h3AOZuNxw55BtsjzORA0OZtSlOgZYADkWzCTgxT89a
5DBjIL8/9OI3ZGr3tZqQINUeci1Vt6ip1yylayW7+Du5J3lX/XVPyKwkjFLngAysEgk918PKZi2O
fggjuv9kqyLmoCwu9ZD2CKyGs+P/Ik5K+tiR0nIzheiJ4Ml/QJ2tN56VrU4UseoFs29U1KBUMn3f
il9NLW4kvqoGIEDOZQVLzO8ePDNocbJ+ThwidlNvtAZyuDkjM0PkH8HZ4X9DQm1CKetK+3VhM7xl
rZJL+OAuF5GptZ+qMWiBjZMAKJwN39EZtEmIx+RSTVDwXK3bcGSAi44roILBcwbFwUAUW//aJcF3
ETdpTLRcL8Je9n6eq9KHc2LFk+LoQ7784ISNUiMvtSG1JejRgSIvMI9EV4kJAQaCLiozIfIkiZxn
WrUMl+wBhEfEKLz35lA4NjqPKwDYmJAr+vzt0cXo1amxaY1vk4hmtWxw7pfceTPpMf4js23kbZ+w
9qNQRvK8HjUzlq2X0Q2JYND3DNJDJHsFTmug5N/LfdfPQAez02nKKhfJuRaMCVhVc4TsFDmJy0g4
TZp08g2V3/0pttvVansfC9Afoi2tzJg0JvxPpqVkL4CWMYycoG+hDteu2VtOmhw+2EVm9OLEm0ki
a5nfcP2MLIRRt17qY9PQm4wbQ5LmSjs/qesn5LJihX9P5WcOuJ+zM8JD1mTwcunfMffIBejfZOzg
jZv0LAWLEJTzMWreboyokKNWCYAKymDjiETyNC8QJLwHatOe2DI0ujnBXHZvsEr4PMvAzW0nfOhi
M33BE17QIwEvtrHq8c3p9PgxlWRnDVSSVteAwD9GSGbqTiN2JPvXpBs62RE/ukqWl5PJEsY+QUvJ
ZXwoKqSA5/ClHh8H+XycpQA4AfpTTEqhmOdy4Ndh9STWe+JYE4AvEL1NcfUrHZnwI+1/C6gTe6ef
85RtwuDrop43ANHXe9PGjLFEaha6Ifa+FqMLPzrUbpsB/7zXDUBQR42w9FBZLNZW1SQYuS8vlqok
aFqrCS+ei36e1CN/O1q92McI+P2KI5EnUcRrN6JzXb+H2IEAwprpNZw9AymIaOUT9t9PUIDDMLc2
/iFwgfVVyZO8AyiboSIjANn6Goh6SunJYkoWlIud7a0FMddP+RvvyLAX0JCesQOsHc6YJbToE2QE
H47z79Mg4hfFUFLNO/Gl1/2b34w823+mtcL08Oq6YoyP4wMxTLZrLbE7UI0RpJeBYzbs2z/NJcN+
BtlY26Otrt3V2o8Rtx3RQSvlD9u6SdAIctouAr+ZDkilsYbz42r+1r+EN+7CcHLwmjRp1DCvke8O
5jlIt7Hbr7fejSInXLWh2kb/aoXLPdggQFdZaNAga9MT7fDbiQJryLqow6oZCFz1ow9WOjhqeTvz
yyR7tJM64D/CZ5ru8S2XE5SfzgJMYtaGvMvcaQ8fyIspZTRSNmV5gkXEN2C0yUtluSkb+PJbfaWp
6KAOJvPyidl543+yJnyDQV+STEmdCGXXACDxhVuup8CQIgEod/7v4rkVvG1OjUsohfE96kSALSbM
G1NKZ6hU4ZvqAxIFYH7qAweq+S5tQhj0LHqvSEBKWyQ1sevmCV8sHX/Y/sVkZi2tW1Dd3cmtI4Pg
DQ7rxmVO58fJtVsh9MIn5b6axFuL8fHsuWd50aK2GX0xwBO0LF3k0VHLuMK3tj60IkkqhRWLw70K
Jx6weTFS4DODdD76i/RcEJIODQW+dy5yGG0G7rWyk73Xzk1OSx6m18KGIADJm7FWnsBjcdU2KiHl
7NUWzAIfWWbvg4mFxGrBkkQ66QqL59OHDIznPPvkMST5+IeziRg8XeBoZxrf9H9qsGffk3kYueba
zqZhHPVSfFrSwk9+jc/r1cSYsPRBW+Ls4WJw6uR1jG1yGUI0zC85Eu7aPi4u27ALXwEp3A2Uv4yp
9PjnGcxij9+KVdbdL07LbIAyv58WVKCrbxVJsPvvl98SdIQuAZ8XaGA+Ut2dQlocv4TYOezwjn//
x7+Hl9LTXwEdHaZLwMu+51L7sbgwFWCbUkWJN/gK+WNBYK2VAfsK1X58fASg4aFOrdBIHw8tvLR/
OFToj2WOOPDFIHVRIJME1lrrYFN/NyU7rY5wvdEOZ1y374/ihtEHw+Tx0AzdOPvuHYu1IUcrOMBa
xQdbTcUei6df/CFJgzy66l/sWqbuU2j8fmUY9eDanKs4jJqHu/y2f1wNsakMe5wWpnAiMDaOJedu
lwBRlZu9RrornpJZIZ5QgKYFQaBYJKJBErXul8M7lvabNnNjPZFJ55Ak2Onb2c603YqFBQGEd4LJ
+WRV+G+8CMPNcu90wax/xPkZgU9e6wXugX7gEFaS18sdWmYXwBKRtmsm28ou8FRFLIjfSrHOHsyZ
22+txfN3vS7XBNw0VQ+aTfFoRxIqSk+v0M52ch/WuxVWW46sqAhdTq5iFdljK6i32ptivPkMNzB0
ZSAoTQeVWcTLcO9fc0wJFLQPgDfNbISnoRoejX0cGeq6BKjR7t3jhKl9N+0vumYxLhwkL5qaP/Ws
rey4d7iRlmGFR3x4YbiemddV1zMlggkr3DQkUMncQhyNOCyzDPZfKzN2CKV8ftgr+UMZt1vO7g9/
bxfpbahyh7799SqyncTIKmHiS/mAkCrAaPMxLKPOh+6IToJHI0ZAw3VebWnfsHRlyD7JvCm6b9Jt
+ziBg8XVlp65QkHnDj+ngdF8j94kUpBEADcqQ103o3ENu/IYufABVN0w470PzN8nbwt6PXOuDJvR
dJTq1yxyeu0cg4dxeyKcG+RrYQWQ/W+dJn27EpMw1rFM1ldrZroTBmV7/3Jzn8JzGGtv896L0CJu
USkvhZAcDZqlLtH8dkzMYAf06KGfrUl2R4o2J1aHZLLUJR71f4XOnlqFAeuSUsVDNU3dnX4vXT5l
r3Ehy+5ssEQczUFpUQOKFR3nO1BQZXiSMKMUucNyIkjBOLvj7PURXekDIWCnmvO7C7O+I2C3GOf7
HBHIjNX5mom9PBNGk/ndoe0wQmPscFmZiwJxZ8Xq2jNzjX+egE27XSAtuXVcRp88Y38qIBiCBtLv
amNgKBu62twI2TLVQv81YlwiDYGXtGjqF4DO7AYPZCLVbMICcGixxeykVnoOHkTmE1LektZAlWNW
MEh+5whHwKJdxo4U0XL2i1pq8RwWdZCjrvi7pKaqdJWtRHQh18y6n4znnwGMGzLi/gfeuAjaVSs1
6cFVSwsRd4ESkzS0hLJkJqUkHMGFilpd9b4HnJdjQUjdubfK5ALnJ07WmboZrhij1oNttcz4cNCD
ZILQalQponDelyNEcNNIElE+l+7UALFcYDH0Caf9YZLmScZFNOLoYoDvZ4dvF88ykiGp67EbztHt
f8k7HhXpcxCU5Z4Ulm7l23ME85GZ/amEyaI36RZgXrW/6mF8zwc6XD1B3U8aFx6eWQ04hUOL9jw9
i5zowuypYWc9SSObNI/r9foFXF4xQNrWga/VjUSm2HQI+cvcQ/w5DWZQqmXt5DrvOCUXu+a2D7BZ
uKRUWqG2rElOHeYFhhfDs/3je6nX0IjenWVpkV3xxklXDIPCA4jwTgGLEo7+AM8Bf5FLG+k4El8K
+O0SF9I/XcsKR9vWaN+LSLFNwp6RnPwsxa11PR0drjDobdFpQm3ibrnQr5Ids/TXpe+57nRNqfzh
Uy8U8/Nvvg+vrmm6V80/RRbr3ZedOy8D5600GZKFKnIO3YfSHR9OwSrATYggYr8b0dlLJmTt/1hb
y4/OGsedhGeY3ek1Fj46aAX9dfeTlM864n706EtJARXavsSrXeKE4YpSQ2dl00/il5ZEt8CvM0gf
8hbN/KWRHhH2TmB00ewtH3UTw5lbj0QIQpJyzmn1vNR1bEYfem9XvSPGnL48Cf5wv0gODAaM+y6s
aZUtovk/E9Xw2PTo8hKK2MKK+jO0sAvp3CNgzH4kB+byWfG4L7Gfttbx9LF3bc114nor8dLVEClQ
cDT3dHvx349Nh6INkCVWg0lBj7e830rurgENiHdJspzibR3NThVPSffnlcHVcdUMhat59WjNpJdv
SCuHLRWoB257MZe5cC7IDuNL7/HYD3WHwZykdjbezkxnzVOkf/rW2xzLTbC44EqUVAI+aoV6mMa+
8Bl6BRwAb53QLaomwobepfeIT0LJck67N5J5Rqr9Z/NDOLgBmz4hZxQdS3IsEUImvAfmba8YntGr
hyp/+vkBDGZdrREh4SynF4xa9ICK+ORqath7Cv45FUG90gKWLj3rQExHbQv/c6OTNGu+/jgnb4N7
h/PitYtN0OgTWlVNevTYoUIg5kGSogPMk7r4upn4ojbxL56YaRH/8ucDInKSVblLKbqzoUAok6Wq
G06a87pJ0ao+CjYDU0R3bH1aw8LSzQQ3O5vdAaNXE4usmIA1hFn8MXrfvBV4/Y8ZedjI7JH6ek2m
crlvH6pBoRGL+p6g+srBSv6se4UqXzgddejvea1aVQ0SwGlkj4DL+lTrU6gqeu/X8/0Nnv8ENPqb
ktZNR3t3Hh7Vo70NYj+2pE6UkfPKNSlLxHP3nRg5l2j9YDRXGmMIMT4BHX4T0ZDRTvPEWlRklxcB
RYXUrRNYGRcqED9waherFKNCTeFQ9+29O4nJeVfWXJInOSr2GeE7dW+Eal30LkfaCaqExTKCZJer
ik73ygf1ZXV1mw+dKDNYL6o5Cw4w28fU9zrpEvmDtCCt0mglQC1SXpgbu8Y69vgX5U6y9xpnhJ1g
bU4m1ffsZdOiQYOxpz7h7O5yDVITJxvcBXkz7PiCaZQrTPxPCb6Aq8llIxcZ2zwHp43KNoU6N5ZL
4md/IHGIEIto2tY1WRg8xiYcPhOKA1FRfBKQcPN0PLpGkEMGjtmEJ7atdxhqFsW6B+WLZ2i5SrNL
3C08fIfpXSrGu/PvIZwQiM4QF1BXia55GuO6KqwUNFKbXJd5JW8WNgBwS6bON5y17MK8U+hUem4w
e2kCGMPOXjb2BmY4JOaE/2Jr98wrcnpAE+KJ5eMmzvCi5Bqtkf7vLdqJZGOCqtY8719U1rx960RQ
7sZ4Yc3UXck/BE/a0bZdCReJLhZ6PCQHPOjmY8vBKQoxckgiEFAofrKyzfy/MQDYqmf0hC6Izclk
I5ddp3nwTsEQnGeZjFAmdLSSlx1z//2ZtC8838pR+aOxRHirjkMH2Ac8WkCSRKl1syXCSHkRZgBN
aaKeDBqGjHheRpnrzJlygJP48h3MqFc0B4+psxJJuh1moXGJO1IK9VQ3mq/RhZaOQqBNVQ2fA43l
zXK64E5Z4IuaWEV1vIB184Grq3Lq4zXHt12ez+j+FoRTKLcwMq/qM9fchn/dgaz9wlLszwSbLGPj
a2v/RV83WBQasgMCrAdTaC03j2rbKuYLkkYxzdteHZL8oBd6FpWbamMgKkKDagOCK836ave0tg3J
jnAJ1LZpieMGAiMId1ZlYXuwufX1UcseEMgxil/WHZs1A92agBLy0hPu9GdATbzMqAuV+aaAQZPd
B+PyYWvVLGLdrRH7mqen99pcjta7/wYFbCLWLoEqZXbRxgmSyZgLyHpFyOQIVfvafbXvxd67c4jc
TVn+AWIrrLsutPleN30OwI1Ww1Pp4urwfkTiB0RBJZzpKnFslaITq9MrTknwlEETzVtyHijgQ4RG
VVyJpa2wRexj2A5bcB7zvrGgFRuG4v824M02HiMAALyEblk0Iaynuba7ohmsIceADVGGRlDzzhFj
Pk8JUTmhxnB+uafG06mC3RxoLbPRLzprOX22DRNx15JJQ0/+x1HfV0KX+NLddpdjFGrHlyda+tdI
zwdrqpGY6K0w/+m6lmghucEaCGaJcMtk4rfqC9uGhkvqCcDqC7CpE0yjWE2ff6zgoqV0sGGdm8L8
OlCtHOg7d7/Y9XieAMZF+MTOChhYdqOTNpVN1By/rKAZGGnUgwaSUmXZ/GZifcoRyJZia4VAYUfH
OXCILCHklwo9avfd+A5BG98HARDHHZyFlfICFajPF6H+GmtqwLnFiNbvqD5cXaqfQ/z2ejJYCb/4
AYAdRKcXLp/DZ7bzJz3ENuuH3Tklw4zPJmmGSQ547/H9nIwkcjs12nGDduQ2BEW40CawQFVCGf7j
IE6HFEr1Jpd47w1HPcViFwKpjJd+PqudzxLLJDIYoBAkWCcm2LGFUkg570w9K4DTMBgr8NTzzY71
gkZJ8OkO/7f2AjDe1HAHVowLKqBgItgz5Yul4En59PBwt3CJ9sWw+JhX3vuFIdeBwJwpq3Sfe+fl
bL6sAdgselaemx7FzIGhUEjbwHitnVYr3NvPrtJdQGNj472+SsJcYUViVOYoJhl0ZcDi4Svi283o
0sXpUAeeB3lD14yjyiCBYAVRtR/jZtEW1yP5Z7X5YXk3KZfXkRUnd+PsLkDn8agukLqvGdxxNPXs
7LJG2FTsxqG34PihinPjMRBoar1DHJB0IGutvYnx6U6nZO5bF+rlww8uKZ6xnrI8rkkfu6lXl1Ym
nIl7PE5vp3GRI1JCNJm5Zo9BlDSlMv3mWPwFcI4rmyQVVlauD+0Fl4ZH2pRNqMWcaIMMP7IYoSC4
bao8NuIkfNYmDWsCF0mpTLnqwQi/9DQ92sSW/Sy4PogRJ+UcWOFj7lbhkbj9/Z3iN/2JbQYPFuKQ
9wDUiwymEKs0BZfnSGkNnJWhvAzvj/GdsRAjc7rj4wGM1ftiyCck00EA6I35tYHXOO482pijpPIf
KR4t73C1XqNIZ4bUBq7QE3YG3KEBSpBvh8NMqXEDk4xuJIF4gKj9Wkc3+pGV9WsqCdpHgFW/+rmW
nAR/qUWBQDwKur28VaX4Ia9x0oa1YgEIanCqVFMS3EVntB8xwH2diSDa5S8vmGgVmFJFmcdgyRl2
/XGx8lVYVEo6p1KWixmdSIRTvo2t6YZTzkGhwr/rtPCVGIyXsYsKiIbik5h9oAWPDTl0ayLble9Y
ucSfMwpc81P0KzIjvscfxSw5yHcXsY5x0DDV7VqZjMnuxqIzxKY6PBCwBiNIJZm5Hxjb07aFPZho
GYHvqJv2Eohzu9rTZX4pki8aGZ6GrUIdmFlS7CGx1l0jQEr6s7ugl2l8r6DC4H0zbjFmHipmwdnI
Jei2mk/dcMZhfKPF7WFRD6OjxSfzPPVWi5v58Ogklyv/a9QGtV5CCrzg1lkRuED+Z9L0vndZUXAZ
J4VdKvrHryQB5LXGeYnuwMBqJER6U1p/lU75mgE52TwS+LAu8D7L2/9b4QtbofG8ocn8piD+0HGb
3tE6B7RdSGxZ03xGrN5Q4GXs6OzWEjR4YJjZ0uyD9hIaU3VieMfgUKZtOfSNruuPxjfhWBsNMgk9
1zkkFckjjmboK7iM0gtwQyFhxg8vo8EVe3ZAsSwB55V62rbxvcePeBvP+dj2TQFV08muIAiH1GGs
t6JMvWZxKO6S8TxV4wnHEPGM5pcBEXLUPXuyKCgUACHZtZGfsF0Pc6ENJR1BHLGohfJCq2nBnpDW
VFjvQi2xY2Zkvw3b0xv89hsTHUj0kv+lfcjwBB6zusFcIpkoVdDYZcV7ZcIY/w4FHkQZZyE6pPA/
7zzs2D7x6lcsOaeMb2NqFKdwP8oIPwl1kKW3q89kbjDbjzATYGcVpzaPDWOY83a6xE5n+pEuvz9A
Q6koluMeTSKRje5vrbG2JfnLwheqbR6k256o82yzCwk8WgMT8LFz/3fIblfhYnTONuYcj1ATl/DQ
E1z/aO0Jm5J0vdwrSRLQNIBYLu+NJI+ZfP8Xwx3SDJ0P+P9m0cGInX/m1dMG9T4qpHR3tSyrrugp
5JihaaHaXtiPBy+kYHPwu0ERoc4RbrgPa/Z407pxnx53qalTFpxdvRNV4HwLynUmVsV86ex5WTtO
wi3D+rAtld8tyYRnioDLAk86dMalnDoHA4JYSbMjwtcbbao5Nq/9Ps6BnTOJ02t5ZQD7g5u1t0fr
wIC/4iFzmIfjIY7Iww3UTHqvlUBlr0la3BeDFxXgO10lvVfjQWVZkrQgk3R/XP4grwMUDP22ZdpD
2KPiV3RmLxmUKbZnjzSChXV95nq15okj2cpUWXkW+EZ4LoQyQ8A8gCIXEt9Zds65vdcZ8bM+swnK
Nx250Mh9tf4GBX9UWYU4JH7nGndh9bcrUVBf0T7GduQFCG6wOjaIwlNtwveeSdCcL8QtT5MGhdth
oYF53kINzAvAFgxsb2Wz++ulUHzNOd2dKJ9S9iGcUuI6AGVT8aXNhRlVqh3K2pf+6lMQee1KTmg2
qzLqSEIoCCgtA9no/d/451a0w2fRlGkXxOYs+vhrdCcQ0TXCFZpY6vL4uzrVeyKmFUPzsxa43QKo
XuFVTlavqHjhFlFoxN82JDFiic+FOdanVJdvWX+jnK7khaN8S7+/9DEIr1Qe2hguizut5knCZjqM
Jsa1+3m3vA926H9oVxwzSzoWWVkA2wRbEy9Q3nFyzlOKGz9/PueDx4M0TaIytK8SZ2lN26mJQN64
TRsdI9j/nKOMFA1+8cKHzUK7zVNDWpPdipF/5761ZKCoBmUP1iojv60gU9Bm5QbaBlpFdt2aoRvH
6XRsloDAOcvCqC3IdiSmdeM4zms/turoOzHpnvl5GxE7AOE3bsiTRJGs2x8zuebBQjcRHSaUaMZb
mlB+uWA4G4fYOzROfTLNHM99PBSnYz9xX5h18jB+Gq9W21yN9UoIL22bWTex1eZAFbc8/vNc957l
cLSzuMM6LWmJl5p5CAUzh6xbNWzc/TMkhJO51zPb0/jOwRAOaS01X4my0mC8Jdl78B74oC99Pg8Q
PBqcUsWItF5CkaoTkiwU6L7zY71kNf8iL64gSeYBHlQSqLW4DtMb6bYIDvPfkH6ADCDyO51KQSEa
qqe8ZaqOlbPdgtoo9+2Gkja7n8J4zioSqjeYjmT30hayga9oYqMIY6p0S5bEuaelz1ljv6Q11zUu
5uSjgXYWKsnhZLPk04X1yZbzQ6+/P4+HlwmImLOSfjkpIDtHOEDbEI22OJMms/OeMsEHHk4PLjad
EOZppsvcP+j1jzc12t3JRUrPX4Wh/PoaCGaf7/mWA5JfoHuVN8SIiyn+IU9oOBfYzyj/e6LY2BOx
UeItFeQMXfDYCJ7+jmHpBiS+fbIHWcYztcBt5PifoqsJj69BNM70W8BffLF0+jYhelRhUbYOE20Z
er7w+k6CXDaj/ZMn9ormtAJv55GIp7uMtZ14siSefbHP2vneKYjzUWL8SVY1qqNyhALvH7BcI9oA
5MjPs7OzCpCKbURj1xqk98dDLT95mepBJg7Vjyp5MFbrX+Zky4LEuOlfhGP00AMO6LbP+U100FUg
uG1NNVrQs0UV/yLnZoLUoddW79/BimhVjuurcP4rfYpstyOJdbYpkqmopl/ff70xdrFDIMquLFBu
C1fs0siueyIvnB2SXfiQoddJyKICqTcHv8HGVA1yJSzTaS8AjpM2LX3iCzpIopRIu9uRw8RlynMS
zRTA/TEwRl0V1bl/qZouKx+Sjs3VFeo43dPW3Wyeho8gzkj03mfaUKwYt2LbNhCFcjbaJ7mGt/2A
SpaO9g9ZhcTyHHfFEZGNSmORzyrhJrWLSXJDlq8F4N80stvg7ppD0gIhrpQb0Atji4oTHxwTfzuJ
2BnsdFSL3B8cdaJoFFpcaGobS/TsUZQ0VleBdQhCatJhmDEpFJaZkcPsuPyRH3PBtSZLJWgw0tPN
dlILA2SsMo6oM2FIg9OSlyHzgnrBzkbiTcc4syGTDdFMAfbl6iMUF3U4yK+46gD63y9k6f5S60Y8
WjdpMovhQPEQVdA3bEzY+xPT8dZL8aQqGyAjcHPoIK+zXmu9iWghxTmkmJb3hlw/6Ud/2ihnZ9GS
p4l4dX+D5kQV3skikZanDTlukfRRDPFs39lnYdIocweY0j93QtrOMmL1Cwvj+kumD4ZEWPKA5dOh
wdcDpay8pu+6yRj/giPZMhB9KpUtqR7cBNeX6MfUXiFcU5izdV9x1eFemJ4QyEGAN6PSmGq5J4x3
OkSGWDffHv2JIaTJlBTikpCSVkcxpn7qPpYs5p8ytCcXNZSecokeSVe9Eq3anep8O0umYDU9mGhA
clIF46c/TKQPFMV3Clsc/NiYqLLH9wugw6sU1uXjxYUKU1p4g/dTToNNWS7yZ3kShYOfgVrHyF91
0FspRhrFn85AilF8Ypn5u6yJ4Y/IZbiFHlG51Up/8KOIdfpdqQRX82UH4ZxmN68PFw1DIS8jWDfW
OqnqwxAw2qwSDJiCNR+Vfu5Z3IxWuPGH35dNggbcK7kmkbd5NuHCuysrsa0AiClqXlcbNhvL0zT+
682t7jfUodAbn8j5w7xEoeoUKKo5VZLyjanXLBRIHo/YdGuT+VtpXmXJQ2z4KHl/Qdopz27gYv2j
AoQ5EpO45sC606BZAW5NsF+ju0+f4u2PzWW3wjHN1Mr3QCsk15BKj/KrYI5vwdp9yz6D/EVXxLq5
p2K1FlSbE2e7070i74E0uRjO5TZTy4GqrMfeIWtqbQCTN2l8th5jlCZ2KDY9cCo+mx3qY+oiFcn2
ifbJj/IB/8ZPfDevRZRKCd6UR0Z/PuA5RVnnzzmgqQG8DC34YSvo5rJKMDvmikUtB8TIqbaHJJKb
SJETI2deNo8uza4wQBKhn4KRKBEl2Su8Xh4+RT3UTmOnRmHzJScaUoZxcCwDpFEuk6wxalqIvY21
l/4gqlIGxZFcOJ2Xw+6Aclz0K9PnpKmn2ZKoWMH8yiD8VObXgI6FvC5uAa85l30zS5ybaUECOaCx
1ZtWH0iksii5XpQysqK7VhiFJDXuy4AhT9Ds4ARve+u7SxrVqb2DKaPoQF23eAhf7mIUtISnB1KK
nDCm6plcEpEtT/iTgvoZ+NKoKXdPWgyxPUxHjuiSGH8QDsjod9zBoVuQP25wUtlcszYMBuKe101h
j+RxPBJoeSoJ0T5wMxD/sylgyjzWMq2JUHxgYlukd/5CVoYPvBAtsqF/Yx8JAcF/QsAekC1/Cksy
z65fZb3p9GR8Ka5RB4PM5JpqnKjVusNnBhydpyV24SAyfpv+76e4VXcZ3LIWPYOneIFfQGjlLQhR
cXQtsbyIMGWStg46tRLY8l270IAC9GPWJAbWAE9cRs8257HWxU998K0H7Y7U2vkLRwP8ZwWti2+q
Nh6Tgn9NOrpJp4ivua666Yyk+kTcXl7QP82F3+9bEtFUa0Si2QLuJdzZdYexu/9wpQdlMBPp0K7i
8yL4Q/Gqw8sbaQG7tzkfpXVClQ/W8mRGDeh/7RYqF0twXnAbAq/FKaOopE2soxrjpFk/szo62dWm
uE+xmFAskCy4dPmXNZCsjPzf10sqhlRelkID1A9ZZQZ8ikUMyIEG/RkmIgCN22gHWcGkuDbIAkK8
k+pBRXngujzE7Al+QVhe7P8G9/q8h7HeHgIbNdzn6gAb63+ZvHihIkaGW+3l9uDZHWdtfZ7Ndmo1
puR7rwvw6OSqBu63sYxjjNehcwpSCPSPKWO/Q18k73OE/+LpMvjAc9WG+ebZxxt2lq+Abti9Kl1i
di//+5UCS9UJOk+Id/jya+tpiumt2dXYhdlUzDwyRLfL24m2wOxF7BhPDk5rhW7FKT5odPo+Yqe7
3PQAl90Zx7k7600NRCzXkT6pj8A81CsN5hii3TaTpses0qcDgwXSa+YlRCqVtsRUeYEeVLb31h3g
CTfbrvgxNT34DnVK/t9NJtiuNRUcQiFRijse/UeR0ki8wmW2BadWuBDsuihApahjK1H2mk0Lk7pk
wMsePg5eh7atAh2sMBPL1J5DFe5hoclHK7RR8pULhY38ksx1WOfucNiDlA+ScHI4oDaFqJr6mIkJ
HAuGkc41nU/s0zLJffFpJcNyEYvtcdBwPJPBQ/lN2EtYHSMV5nIdslYfy8n2fKFmPxtSsdzI5uGz
yTckyhFLmbDOzndV41W4j+4cAO8cgCiPOrU7tQ5g2qe2oCI8Q/IuhzCb9eDtX8iRCPhDc0KnfXEh
9vKbDfJECZQqZCTs4N4jGIXhvqtky0e3E6cFNV5y7wMe56eGt45OStxyo5/aFRIjK9VNYSBQATTr
zJmeP2LyYVsS3AG1eHf9Iad4KbAyddfAcuGkZlcQuuAKen9mYsjDz6atppS/BTRlRXv8CGe4pX/Q
nLw1edLexNgxmx1aYXKF7xg+q+cVSX927obhPeo+Shu6LVDiD9AKJb6mZcCfkqjzqNmByqro75hA
5t+4GF/C9mlJTK28KZLlFYNUyGs7Hmo4658oUIxzfjRZkD/vbjMiOZ8LT0mbvEExAmYCYLIClZCn
ggGa2A8ar2zxdorggHHJ3ZI351VxrmSZx/H1oPold2PC3ZUNfoCVJhYSmG+p+7kfa6TZrdFQmsZo
SzGLMsuEiAgmDY9deNbL0SbOlhwU/wVkw0YpMX4p7pk04HIn2pOHRMEzPQvayswdckjmqyeEdtOI
UPdIXlOl392jkAVlPpY7ss2Jgq9CbvkwJKlgdTU2ynvFNXa2NB0cFsJtOsVvccNFRboQH6U5oL5F
B/sWIRtlc6QM4dOsRI+2F6fGk7EE6tRpNoA1eSBP//ZG2IZscfiGZz8yIh3o3amn1Dj8GDxm7j8Z
aGitQItWkYNM91PIPuUeRXSVAypgeikFlbuz5FJnlRkgCHXC81Km91aeMmr4w0rp8J35BOruWoHp
7OevGBbrnSKVMbUYkkALqw+QtYluQyjyIYTyNIww9HUchFgDNE2wrSpDPupgTtixFBMtpp5KTcAW
qVt8jSuLwfQvbrF3evSHGyMbm6/Og9dnz0AX1+UAt0z6DgOGr1g+8600b82oMWsZA3aHi2xbEs8C
mWbndflPj31QdXYbCROuqg5zqXhlgh4tIGXvN8w+wTfmtmGHX9qXU49HfL49SXjwzV8dxMNai8he
rtzPGbFysiTrOAoyVsVS2mbcwveHZxZZ8Mtt/FXcwAmUvwP697vEttrcinYU5gKc+rxrVM4+Omkr
Rxripbuw/eqSlvMaDjL0/GylYga/zFyajK9vVj1RRC5uxO8H/YqJrfYYBKBdbvS2IPJe2H+2pyj3
196NWdZ1dM8erp02VGlXJGsJ33GQmnGy60JTJcNNiuz4RWRbxy2+SwCF3cA7cgoLyvvEEc73H/fV
4t4p2KFpZTRqXaGomCWqVeKju0eKF+T6MFBRuuISVnWlkxHjJH35Zn5F1FhuXjV81zkhm8hLUkoS
3G4++c1aPuxmWOypVOvaY5Lgvo33AyyvgLKVg1WaeLJXVsIBq269clsGx8vsrb90KWBhUzP5JSB3
zGXe4d2QR4YI6N/AKYN4Gda3Isw4tVegDCSCCJAwnbLeb+WF/XRQtzazPibRQnk4uosNYj3OMT34
gj8dDUhzYc9oLQiZhIHFtB2LBus3pHzWoAW88cX1Ydn52OBX1BK2Fcj3fIC40odSAb20lg5pIMGd
Vjr3ArJdbptnYyn3LzKk64SOFaHyozvP3ZzpRtmHKNMrtJPSCe7N9pABC+lalma426UQL8ROLjnz
0VhKiVEHzW4uqDY8X7hJVWdqWV3f1SvIZPomoYTn2xrkhssklM9uk7hRnQp4V9zZwacJ/1peCti4
kzszSTmqp6Zy9qQ3l1aRTCrkcsR5oUJhBqQQufLt4UOqIjKe9phbONxC442lFHlRBae7hAovMicd
QhNylh6M0CSDch6fYUYxsdJXaaup9dPwmONrhn9550/Lv0td6lSg7bGJu9GVoHoYY0qARQfCluiP
PmiOeAPiEM+MfR+EEgmtlPCDQOxjY80VvZib9KhYzoi5zftxDcnehDQBSfiaHR96/T7CzKi63sK3
dxXZZONMWVm1J/3ATKhsEukUCWmg7ekqDBYfrruf8SRfkbdmhR1tSctce8iJyjlyfCGDHC7Cz38Y
vHXK9aFxXVrtxRuYrZDGP39jksQ3VmyT4fnXpSqu3HNIBCmTiwYU64h2wy5zzx9Y6naYCP7xSHzO
oMUL3j6twlgBSLO2WK7pbXVICtcApC7ztY0rO5XgwkjtSwdW3BOVeQ5337IF87JSMey78/GjHVdB
O5K/QMwcHoX4dLS28nIjv9roZxXtGNG/f7pzDtodi/xQesoflF/5Gl1k1p6QPJQSwZ7Rq7sfRYYX
vO6ifcpMIjoiMYHW9l+rh/UoF4pYQS0Dhwnvm8nfpIaOe+5ScojEXMdY4mBGkWSazHLo9PtdumJv
hW7Af5S4XkZESZ3GAEBiv8HTozgwU4LMD1jeTwquSD5QcK0KYs8NaCCj3Io1ES6/QroAox9KmYTd
eYxrgYLfIHpMwE11TJXCPMGAkNOwLepZFJCfj5KnfHVC7GdCKUfoSsWIJvrI/JLYlSzbciZRqsoQ
q0KFM1I0yZSns91MXesKuh8sSjIeJ7B7HBHFJ8zM17FrzdJv1SdfDhqaMBS/i+yYK8l+pSz3NCPS
klVXjRKQBgtoNEq4T+PD15p8ueM8JUkl5S6WUN+RiqoYXi95/fJysDDsjh6jHDBTYWCWfwR1Oy2/
9jqBzvc7o/MClKdPBCQvcO+xQavXtl3jopWQgtPgEB3fpz2n+kCHlbl3vrhxpFoEuY9B77D6N6AF
OUweSa8ciEiT20ytdXGTT0lEaUobPKelWbdiMk7gHkCwTIMKiZxBJdifXtRQoSj+s7WqzzTzRY4/
b7hq2PgUB8V5EczdmG1t0Ry7fXRSJGn0bLp7nE6a2YIv5ToNnTCOCn719my8bYJbhgZCgbNVKlhG
N8mt696GX8F0dMU/FkRdDgCU/ThaiFHcVTKsHh0BRSaBtFHglAVnvjE4/Jhpl2hkU709Var7PUYr
lk22E0V5j40nI+DgVag5hGJsDFYxC+mSduXoB8lJEfXo1rYc5KmG0Vl0HkKQPOAYI8JDpcttSLBA
Kwc8ZisVojyT0kHbeUD3Vx35Oa7QtfL1Rpe4JFKIaMjx7EaiO8WnGKjXZH/g9YPASWfCsdvRz+CH
EjXfXXIgJwujk8ULkaAw7T+0YuDehHR1W82/HP7E0MbUk/5u3XB6JgpdHFJagPrJgqESFzkXUcFf
2hNWOdYHq0h0hnJWXyBNzLHKKVjHED5ek3kK6Td4n0aBC+S+rtUwaTCPWIdtT/UDzaw0zYBGVVaz
Frgd7IYYya3OteHIO03RXkGFVQI4yc62KlcmCWpoqoQrfWawRJ03paYSH8pzXOISpIE2VDkYA9ND
0Cn2VHSfrzHqg4oxzjeGVms+d1B90tePpZ8pL4dd6wlQxdLZ4Fv19LH/ITRn3Hch2biy6+wnNiZX
3X5TPs5r7JoDjdREZb/bonOIIe+VIzyT6ysVKZrR2J5GHIsBHtq3J1itfOmOm7BpLlBYi+xXxI2u
I/xdnsYbto68TiEJxIuBCf06Vh7nJTnJ1URx+3f3AVzmzy98DGYzbpwyKDyDpmpiztvdT6qLzTSl
SApMMhtYAvAHlOK9z2L1E5FWXFlVGQO0mqTB4yD1XntFaYQleq3e3PPujl7ZyrMiBWr+tsMI19wW
K23usRD3QCk+mJKntIVarpCTzUhNG0d9Ha3el50To0EvMrPpl7z3j/qKUG4yS3nevDVZK19ppZcL
79DNNQ38uORbq9YqFstnYiDKPbqZrg4WxE+w8ii3HgYTBXvNxabIzrtEp/0T9OtECZNt2DXH5OLl
LC9ynDFq7wuQdm3++a68q/5Wm2Y2j1b17d7KOVTSrJW98DfSZarVbVdcA+xAKTOPRyrmHiLEQjQx
BC0tMvtgDdtxI9Cx95f9+NbMWQnqherhEUj9E7th7xE9vKJ8N5T0IIAXosh6VCv6GSm5th4IOub7
Z5hIkyzYjqh/degh08Y/L5xt7HPr4RKBRgYu964G98lduhwTCGz0VZ0WlJqYC54wqs8aeoRZN5zH
Iz6rtFL/629a3wm+poEMoxLEBxbGn8n0T1xWGfZUvQvy5si/B8L0Wm05v+nI2qKXCO/3gSPgP+jT
6qZbI6PtEHPOzDDOUPMhYZmQre29Pc93iRjYeaMI4n2RBlKs8jTG7cPBX8GoaIAypUeZGJ7PprSy
5oGpUY0BPapDQBpcrfvUMZvuoSt0Xc1Q3cWAEaPULA9yw2iukw3fmB2nF5g5beKSFJ9F3iMNXFEZ
DE6LKqB/9Fu7igdwXSywXKwo20ZRaD7a+8M2TIse1Afwe6V7MpVZsXmbDb1d4bQ3TupmLKYT5HA/
yVeZeUrgTXinLFxHhV6cDMRMgASS2hFZ+79OEI5HBz5SYm5T0KI65kRk7aC/wWgWZTlReMVOYKIe
oaXHy4J1Knr0Z6q2K96+L8Pg5yB7mUg6MqmBDqCd+vx5Zlk2OThSAuENy/ItouMmivyg3xW2BVod
Lp6ftMjHeFaO53gKTymKbdA6/Bsi5/rMa9++2O0dVOD8qZ7a1uEQppYZFArhEjIHQynrPA6G4P4/
k60+juui5g2UcHnNN9BnJzKX8aXg77MxKm3nTJyxY0NFroLH50x3nmQ9awZ3xIqise5giZt09+4O
DTFGRSs0q4LEYGvOYgFm/xX88tXZx9V6YB8q4vxrqdZ/RkQf+lHrvTf0+vU83Q9xsu4o8KdbkQfW
P68zD82cw0HVo5p+7/+Hy5rd1tHkvrajAJuF3VTLd2NnBpbU7VfZMxzcL7QiIFULAgDYhbRox+3V
nG22xLuT7QTOELU5ZQRG44zoq96jeTsl80Ytxj+uFC4C1p1vbnl6DREj3bMSf+EUrohnLM1qKEtO
mGLCCL5yI6ofETfkVIF5as4pYAKFC4qmFzBesJC7qDxPMukrjwI1dtpA5dgTUgGxbGF/tSJnXbHw
XtYXuJMtRh6YxhAKeAXc0UWIODKcrAoUYaRDvUZPG+R9g7YNCdBrESLzaEE47CJjibNvrfjNCXsL
edYwLVQ6/MwoV3DAEhY7MFH9oqbYZ18Ac+kUnsbyq1RYVDqB2rX5z06vMLxHGv7Xiej7zDApPpX+
mdzkLkyLCrxYU1Qu9jCkj7hXR24WQdcHCS/v6AjG7sYFzhyOwUUPSIXsaoJ2vuvDaIWXVwUwpUJi
WfUnwjWHmzkztCNKr90uKu8iDWjBVBssWnphQ4nddoUBiX5GURZ3wiWyTZeraBtAFf11OCDhXoIi
J2ti2tgpf7kFkkj7/ogJEUHU8xAxCpRFPcUZONKfJsspTOBPSpb5vwpzMTBPgEgi0DO7W5FLkm75
yUu5YXuSlM9M2EPKmToav1nO0XTi+bhHLslV7E5F6pWRmkWnkaKDq5uPQUBEHyuIaO49mmw/FNPH
fUwk8U3UjlHtOKqg5Fe5/021Inx5VChX17i9Xi5ytaWkMZpGjnSqQSoum4OvtqDwRpiPRNgBNzyR
wGKNFu/D5mQmeTOnlfazR2kV+fZx3h/TuKfVjHJHwlDyux+XLUoZqrC6YJYFd/QzS4tgaZ52+i7d
DS9b7cvPh6AEsRZLXQ+IImZD/uezxItfS8o8aqnnLmoOFawLSLIed6PMmVa/D5iEB/DwE550uZR5
HsOawZzmwxAkoVY0Ef/eMW4l2LIh7CVv+UVaqTC9UJHjsLmKTFGtzLMtFv49NqMbl8EYh/vmdfKI
W4aZjLEmQmvJVKXIXxp19f8VR1hbwI07JTDQknUzYuQNvflNISVa0D68LOmCcsBzlpfYc+hRfPge
u2G57iAhDebXofaj0ImBYfAgoy/g3IRMey2xQrRApxhmsaogrnS/YR2uP6bqSLWrcn/YrP1iostJ
HOOzS4KTEMF3KKPCOURuw2jqe1VirbnKany6JZn5G92g8Q5Pc1PD9365lBdwu8HuFCesdkMxJvDG
MdJ++m6O4ZzOKqSB3GUAZkecD2rSNjF6fKZfs7YNCnaqvfOO01Z+/Lf9rU+7SsYSUP5T3kfPG6/+
qTHabKtAvc3ocatcg3MCMubnY6tPDdEGN6yM5ZDoqovWzCvkG0XipZtscIVQjke7UZ1nM2llO7zf
halkmI8ydPqit049vNZpgUypAZL6ZDwy5cg95BlpSVjPttaC3WnO4KGh5t6DqzAcDpAHBBU5FLun
yYEvz36YnDHFkoMV14YdE1whcDhta8X8SETsYzyYrkmb4VsvGDFJIZudwQ2RG1zUG5daomu07EXj
cV6Ca62iosH0JCW5x/AKH2x4fB0QNuj6vOa/kTUDm/8G3/lmBgxJPAPOJwO6L2e1+GKkpM9rmRiB
eDJwitCRc8cTLjnTRp0yW0sL4bdp+WVKZJcMMJO/rNdQrtdgKWFCNM+MAKvOq7/xebXXr9EuRzs6
YE24qTeN7Ib1a+9RXE6OmV1JBo4UgA0INpcBaYBV17Ob8OFY9p2tR5GAhjT893STa1FaKBBUtKpz
ncFFeKNvRu4m+9vEy800UJKuWC+dW8B60c73s4Wf2a5XdP+WH2Ket8c0Rh2kL3SxsvE5P4y4A/eG
Aek4naUrOYZjGXhs5KE9onGroAQhjHMs11w17M/onNT2qrmkbYXchbj8eYtotRaZCovIgMJl5XOz
X3dY3h74qxj2hQIebOjbGbOp8qCGni3U/vnQNluTquqt+a/p+57N4tYHvweMq6bEC5VR4LtROXY6
UFYI/3HZquDSr8xAH7JmIEL4TlUm1p1QSnJJZCywtzk8uuIL0FCVIBxzO+3NPBtra4asVkz7vo3N
mvuRzjQ16e80C0z0M5toPC6ezQcnJFKvPlnzCb1jKo38FCRPka1BqIVrSDducTTFi52hgxIdH2Pl
psdWtOvQSWHmGy/8NzK/wy+8MmH/zU/xcg5G8r1o9lCTUIQsPOgMarMCSDlADXz+rXxno26y5r/x
JG1ARhlREjliBK5lrkFs+0+kMMUecjVCVmKNQayes0MnhaKakQxU2/O+lGuRrORauAmIBm2DTfXT
LPSf4RnlSXzqAbD//jtVMysp3b1/DI6XTQ83t+qlCrLdeIU8B+klZOQ7la3lhHwfJi2urKHmJIw9
e+XPBSqXeQPfgrFir3ZXhFuoql1B2qo3tmLqLZycfkBMG/H1nL/WE8XklkRI4Z2829azIBp++RG+
PQP6KqNNsyQj0xBJ9gcXPYHP4wSXfjM0Qs4iwrSFknKorzl3S/9TaYIzjq0ozBjujsJEuraBhVfv
aCaX7wa9eZRosIxRgxM6NQO9AmT4xvIUpw60ro5IvTloC7pePiaLqBwCVmc5TTjY2P3C24ckBPPs
W4aZ6BRzL9RGyEOYWOJo9ePMf8Ly2KGSlkLDu9FfIaZjjX2nWdE5RDcuSOKAhgI3LRqGzy/OFOUm
aTV1/p4WWGeRHlL8l+EzhmfbrPU1lWVSRSlnja8elBHfxf9T6sxr18vwkk2vVqsAmjcOijqa8MO0
SUUPISHbKisTq1vtKVxwBKwiZi4PxbQow4Wh1jafkj1WxjAyThIX3c9KFqGz2YaKz563GLmrjNgS
tZ6UOZIczoGNZRgG2zTd40od2yozOSTu3/K9ZCIxTVkIRkmR8eih5wPizcSBuc8aBrY0vhpH61vi
9/myfqGgb6yc/9mNbywuDpmT980xsu2Smu4bfC8O1U4UOV3n+0dVlW/ABtlOSsvbg7P3Ew66NlRH
iv7BfO0aHpstZOGTz6dnAVxmdFtKEbPlk4UknmjZmLZh/7MBS4t4ORvWnqIjnE4g2DdLj/qOK5ja
JKPTrU5sCa2ZxXZGCO5pnRK+F3c2g1dm4u+Hlj4rYk1obPh2peDkNzMHrcHRW9kapqtNx5weq/nE
bTe9hEfLhCv/exfcLqQ+D6QoYpYf+NC4Ybn0p2PgvyMNfcCcFzC3ZN6UKK3wr/obnq8HlWZBAhry
TomjKFl/7zmP6HxXnA0fjChNrMKzjzRmfLh3fa6XPNBkpoA6CRuos4T4tUmI23lxhwYTTWlHpv5k
n+XBdYyU1AaPirn8gOTa77wml3wOFRaTOi4dJq6xLprm3sLZmSx2/FfWiUsWccF40c4KYZepIKBn
P64TinTN/UecEejhT4lnhZGeBHL+O6irGMWFpA2h2jM1nCDDMI3mgxqBrx44afbXUTvjY+AFYoCQ
4Zjh6oGHDqELZvPV7Vo3PA72k7HTrSZOTuxgN+KTcutykzYsVP1X/dVYSE1NNubATjXFXiFWH2G/
ghQytqmd+vSlw6siUpZom21Z/occtF2sWmqo3Q/fAXWHG+WhvDFt9/HNVALUfkE94rzGjBo0lCo0
6IGF8UfGTBpM4VDtItpDKBkXKqjy3+1MoY0Dgd/ahnVc43ahdQqRat4tD6E7yTHL+tA9LLhfTiIV
4yjsAOPrsIjA08GX4YvqtGsDArJr6FAFj1rFoKj3dINWuvh35IPpAOyZct0ceZP0rDsawSsEN0Zv
1kLm9i9itcG/+9tN0YGDO6lB+O7RBn6OzEpOVTaK8KEw1uq1slQjf69X3TlsTnal0FjJTrBWh8V7
XBhw5U767i2CUrE1hKT/wEEz2nZ/b8UlRywPBfdLhzcMzoOsXFYETfohIW8CCwnQkYwCxDBbJbDC
VBkmTAJMekPbY+92dpHOgM1kGi9WevoG3xY7m3Y6p2hze5fDwTAk7U6UYNDvQU3ElkXNjz2Mn8kQ
qdpslKKL02YN4Lrna8mh4vlisNBaUJvMEJ/3JFf9EdkG0+IizpWNILzvC41G5N4oIFgfREKHoAUY
MsRL6MnqjcAAi2jVif7SfOj4FhU6Mkg6idhAmlmQ/sw2ij5RD8pmGRVlddphE1nESNwwQ25bR2ww
U5372YoWoYLHojUbu2Fb4YB1nAws4ASbgHctHJOIN5IB5IcuZuUSRJ+W/oLLlrZbLVz6sI3SbyYa
lMvjcvAiExS/y2/OcUjsLmLSsmg/fvrq9PmUtml7eQY9Z+ECF5G1CD5vU7JRytwg/x3ooeo1Bq9Q
y7sPI81UuDnALp/HeYruaLlzSneTgfgiuOwNwOxjHZ2G5ADS7s1FeJp7tF+iF7fAExWgJFhA44ZO
8RW5OjKzLIJ7jTGtSYGXIgWrM7E2jjq5pfZmvgBZpNDsTnf5VlM0R3/54YshtssV+YhieeeK+ixd
IvL2XkdQ3ac1PL+FF0Ass7BJvRJ5MmD2XotH/ONWEqLtINgZ8R3WlqXpeS1nzLuHvZl1JjRWPNOg
sPdXhhvyueRURAoWuqcuKUF1aGtPahSBJyaQtHx9WEKM72XDV6fSZnXmu6YhpPguwcwwe53CJfpZ
ldnSQwPj2IAVx0f2dV/FP06386y0Xf+O4P4YobaEqXwW206n/v6dMNLX0Yzc9B7iCdi1TQQaIyiu
BShdzuosJpJWvzyjNShRESDe2uo0UK04QaONLmfktgCPvaXWFS0CX0YtoKa2h3YSPfqU0n5Y9vr4
bvEzxvimOgWFZzjwxoTKkPLqKCky2v9RF7lzjz4sfTdU0ljvomcgMymjJliLEW1T9PijGrmtDpJ2
LoLJ/6NYn2VOqJKaGQSPHJbCKB9teouzi75TLE6CkT5vcEdH7RnyYqYn2ftikZ4UInKor1A+hF70
+YmtrUUd25Jx5jU4eNamEcJQDrHUbH8XVr4XH9R1wpjmezjBrquk0XwYQUCSE7duotrbk087HiEf
YL2qPZO7fksw6S3w2aFEhpVQleN+LeuTeBU6F1Tgb4mcIj6v4xL2l4V+9oUjyUDgjLORCJgRQ4e/
ygvfXHHv6KHpmw88Sw08dCKlmKsbxbFtVT8zrfUFFnoBM6lU912k4lWi4aWqJwTInAb5E51GlQcM
2a7Li2MkUOTs/k+ANjANqxq3p4h/Z6zz34NPa916WKHie0+JxXMgsPmcg5t+r0mQHJYWDI6yL9a5
hwgv/Ny+1vpk1rtCZr9hInGJYllphQNiJpturP8ITtRHM2yC0sXjek/0wwjmhc0UqqRqCUxtfLTX
iW0LAPglmqlYI/pvmVQn374ijyxfmEG36S1zg4zksuBkdOwqE0VX1ZYk7lmF0wJ2aXSwdyhJTh+q
Uwuaq4pH8UAxtHMxxhz1zx3P719IY7X1hgymWJkXMx3caIHlVEcQbKazjhbL0LuAAgfHbOLcjsGy
rRCb+yrMosHPQpbUjaICHqV/lxor95WkveOKLNAjAvy7QYPi/DwYk52ytEAEyNYkv7KiSMENT2oi
JESdtrnsZByIFeERh2ALAeyeoJgFGp6YlJlwfQegjy6WLa46RRituPhcSttSD0XkeAxi98pv4BbL
DWMxD+HRz4nXg4JibHFmBw8uhRcf3h8MRjMlYk/LsBQxKXJQSPNLkVBztljsX/axgcFH4ckP2Lbe
41S4VXvzeTm88i11IhMryYvc3gGIoT+kUu+u/rfGwTNp6QDDikvZx2WK/qW0WueiuOsHRVwOZlD7
VkRvMh0Lrot7MwReTYPGFNh5TTLrWVOahcJ/cRDawXlHWhDKq5Kp2YXSwduta4mcimLTfntk9TTn
bispTydDY6HOTszMfloqN74RV6JRxMLee4ss2vt88jaZo0l2bXDsq/+In2MbI5TKhm6R0jigU7Dv
HvEIpw8GHg9CjIKKOaiOKywAjhfC0m1fzT/R3jrpiOvcQsaSSRXuUukjk/O3LZCjzawkCu4P9Tre
l/tfKsQcM/m22IW3MPZ7vfdU6cDM6rImJDZAUXjNJ3mvArVDfePYO9BUD142UIc/NXFSMlHIx5ye
BsywO9WH5kIOyV+gJnVYfXttXvmRenzjjXgV4/OABul8swZ8iwLTq5cU0M2kVKd9ImHqsu1lCcwh
htuX56eK9B0uuQEHyIm5qodlLF1/ELeMTFFWhO/l8O2snuD4kLL8srtARz5waT+zwJI6inRLJ652
dD8cYkCoRx6Ard7T88DY8g3kIhPdKHcr61xBblrl8NR72rwaLCKQ0NO+CibH3Z0nOJrCbx+8pngX
mEmW+CC4l/MHdCSpVp22yhisfB+zt5BfBqXTnHQ3dPMF3T0paSyB334U851MalTKo6mniChO1sGQ
pnaGssT5MuyDuoZhOBDhoJcZEa3uqyohx5f3/VrCI+VXWA4VXWIoWUKcR4GjSQUBGrReF1DjE5Op
DvRpMnZZEMLZEDW5cllq+ktULqlXu27gIShAZtACS2Q43YBhD7LWK0CFqx6teX/UdcHh9T+Vk8Bg
03LW5Zn+JTGDJwJml61ZIcSrL7isyU1a3tZOEyp46uNkfLmERgAB8T75gIE7AokBvYsVviatm0IB
CwBp/LQq0vyDljkaKD3MBMs/WMVCBN5Ip38tHOiqaNAlrXMAtLHYXTDrpoIDeXuPHGLyZGYnRJH7
WvhvRQ5YhO72FPOaDgiRaYalxmm5xbGQfg2TG4QMHzBsgEQH8kq4PSE8xHMnIXLIfzzLQ2Ukvcm3
slerN255aNPdJvWMjT0D+j5EVK9q5sseh3ORQMfsaTZewtG0qgo6f2G6IEccjswKijl8Plm22Xmf
g4aVyO9zqLE0XeBeDYL5l3o56fBxGwxu42gTIHTYxaGFHjIlNafA9gpKNrF4IQBrIzMw5TML1YgB
U8qO7+30xaJl4fuzwKyWyZbgYlFUGp6XtdFEw9anaPUrswebxaqDHRweE0C/ndE/6XtbGF/qoG9b
Xwxf/LVrrK74gF/IFNg2CDh7vId0ZSw6aU4nG7ZDCt9cR2bQGlrYa8MM36gG8UDSXC02/UD0o2uP
jtopmC/Ufo3QBO6lmot6mbUVpLtKjvCTRU0Bsv5VuqHkq7wDyvExKjNzZvpO/4YJDH3Hrv+gYX2M
6jC/K6nbe7jDbbZVnNlFdjEevcOwMeBFlLa2dyRhLqh2ACpqKabTm7EvXYtiNSI3PsIAgk1WrWHT
NEJ+ZRB5TvGHLhBz7Ll5NZsnFKP2NqSgluXM/li+WC4gd04FCl13QHftD7fd6zVeYCQArMSVrWTT
cwO2DXgZvya4gbdGZG646Ob4FvBNhzwbS6Thf0JDIE3d+59C61W31W/86WpEgdRAvNQKPkQHJJ5/
Vju+RhoGgnfwAJr39j7td+iQ2A95zgABgXubUcUv5XK93vCJImS/4HkI2qJ5fyPDk9cXcYl0O4sv
hWCxzVL6g3Uc/fQprcORV87tRnSmsqq3cL3yEoxKoYteRgg/GSMzSaKMwmO5BzdTODvm+zvVgSbl
AAOu7V3y4NH77fpgdH+Szw9sSJEOsyor1aXl9f5N8qrqpxgwaYPYwdbCUrd9Uxs1ThLu+3hsmT66
epH75do02qPwYOsMzkw7QgtwWJSbGTj9ZAvdxk7uSNIf+4tqY6YBnF5rZiPAeVKLlxQZNpU26CSF
GhhfM1cmhLpcHDvm6+0obGH8ZcSlIA/+ZkQxFzar5UZaiiLPvLjmjU91NgdkJAz3aBhTjIFOJkQ5
jQFhfnTJJvyb2km3ef+YD13zEbPY8IkBsOGsSsbOctpa59RyxNf24/9qGo/lF3ef01adhWEJS0Qf
yE14pRhKBArp2xxBOYNignCLmrr+jwekWDKpduA9BS9nwL+mQ0DecvB2yFpzUn218CSf8kAW/h0y
4OuGoQrFB4dDLYJCtTlaSwtMrFs0MTLY1ujJLHJNfD6fq76jrxAshjQgSS1ybegpGhH3CLC3JVbE
45Z0Ihq3voGI0A5MhIW3hqfeh5oyhYoGWb5Dq/jJdestwsMQwasRiJv9XGCyEqqlsJkJs5HWKF7p
XYyNpm6skaRQPNwgSp/P5zsCGdUT1AYUcKyeCdTk77OGEQKZ/obIQ9mBwCudTfvHFAGD70Rxqi+R
+3tVPaLGgsvYuKZ+3iGJzkgkez+w02xHcI/1ki1WDV8qIcgpDXJdKGuBlFegogByOy3cl2I/q9lr
1gFy6qQMMpIFuIsEQetcJgelpUw8o3wI19EIk1Qwv5CoqTmDeUkPJnyPVhCDlqKj1GTSHZXzbCw5
5aDY13tn7ThEMCt5aRP2s+yEKi3RQ+p1Rns3ZPeFVAshc7LBvUcNCCE2rrQvUcAQovvRLR+tAjfy
nHe/JNxkvwgfSEqbi+iCmpVS2yBVGQs3BXdgp4J2Si45ZfjjEdQlQ09yHwCOBSwet6nGSi/LbIy0
NGLLyHxmJUW45fsW1PUxgONv/kiqmR6QtS5kTtYGAzkQgDnowkfU/ReEpcF330wxIGLnb0s4auaf
cydL4J7fu85bwUsbnuMze7LEygSixxVlMHJFjel+Zx9JE1FZ7SAZWi8oIq12Sze4gfKJG7yR24s+
uRW6C2aTNZChu3+VdKtF8Syn3jnZh5X0ASP2UPKbo0STuLeakgyXN2271NCPM7aMSBvgU9fDvjsk
QbKQ2927F175kXnXDfUz+QatX2Bn0creZSK8Pid3kJdJE6iONdp2lLrSIPKtdz+t3IezpS6/PoHD
r4FFX29ktY1yuWDl70SlGvG1Ipcfb9Fg/ntPjWOkru035m4gtsxRMNdROiCldd/fcTkaZy3fIj8/
/whnjefUomnu7z6p0elJ9iZ85AFiPbufQQO/wpjbYt6WVxJwJEd113sExyOK+k5I62artLM7DLyk
Y/G4QFiB5C5GfQ0opHodB6AkEYlOXl6e519rePpg21qEeNhdsgIA6fvibEr9Rui4AYzuzopSko5s
brik4WlQbrZPQNvGN89ahRChm4ZN/3MqrE/+bxtcOSkts5GdjQm+5dM8ejRTQUe5nBwHoZ/OZrRT
Dk4oCRf/bIFerbdoRFKPIK91L0DBEPydlbtHDT2S/qgGKTXm83KvP2++oCK9CS6EH83hAKkTBwze
6wtdoKM9PeV8K14sJ18UzCODFYcz4HjMk6dz84uhYD4458vzD+33PoHNkVwWUxZFt35Coymm3yW3
eszw2u8Pe3noMU073hhZyPdqGs2h3UUYtIuzaPm8R+Fpwc1ZsTAjYizPlHOvy3ZtgRxBY91uRate
3OX3f9C6/W1BIn6wAaPCO1Z7BHQHeA5TiwZ6ij7gB53VrqXZEmvCyPchM/v/AUEcHj3NELZQ51t2
AR+9Ww1j78TqvwBvytlca4BYwTJvoTV+BQcaVQjX+NxsnOOpobUrazDGCdW/ml2P5z28ydLgIvZ1
LVX8+SCnk3MY1H2PkSF/Y+ttpkIreGdxqZv55NSBbNFDfb9EYgLTbb2zzTBVe8MXTgXkephty4q4
XBgLSCGQoIjSzI8xmjOy5MtpoGPcPf0mGBvO0KRiyzYVDdco9Kfd3Oi/kUboFRK+n4lWkZvxVKQD
zoO0R0C/CVfyng6Rwz+xxzuyWz4ui8u0JiExClCdZ6kdhpDRhTpGfx4pb+NNQW/Bp4iWdmhcnpXA
M6r3l1tKDslSpa3ok1qP3kLpk4mf6J1QjjukFo5dQBFEPbO3lJEOBZVPgHwjGhOynlV/3FR9W6AY
Qhd7usbTRnltx3lzirWwWGNXGvQpDYTvztWAN6mS9Y6LG31I3yb2ZcgvQc5RCRzboPyJaK8W7Gy1
qRO94lHLf0Ci8yd+TKHjESeSevsE9JeiNPsE5i92t1DqG1sBBSX1A9huYNU8/5GMrs18jcEQYLNL
gNPfbPYX4ez5NHxyQDjpcnbjjwrtABNRxZhOZZTjgeWTkEeqrhKfAAcXs2uAXknMuip6kCmYd8C4
WlpYEjBtN0E7N5P021xC8q2lzi/JLQr9FeIIAHgjfGc5XGUGe8zoKzuQyeUKemiO6sHvR7EPHgDi
2pFIILumZXI9CfLE3zFiMjHLjzSIFm9ydm5mXKALja4SneS4o9HjyoA+pJrBI/DTYXcEbY91pVtB
gxr4gcrzdW1FdNdzXwNdQ6Sjtbj5CnCV3AYMx1b33HI/vuQwcDjgf47RoZAyv0F785ycZ8ngjINU
l4K7SspgMGrre+F5890BXneaXzLN39/QIfCCUabRiYUxlbXnKufDv2e9NX5lRXhp8UfpVVoZPce+
tqo2vTMXN/Jn0D++QxLPFK6Vx2/qTvW1w1mbVl46GLBJ/8BIcI67CbWISIVgu1cHIOMR2B9D1uG9
D4XiW/ISrJn0b/vYVIOFwaZ4GCaMnLfBvk+e7uhtngy860l0YueQOcHWqlWAn0pu0P8QLsMEz7V0
aDPlqPpk0qNqTOelPPNbp/aAgWWMp9XF8M4PvwxhuXzN1qwfhYy71FilRIl8UU4rxsDYlRPfPk0+
szSO2d8neYoGiAYtxLjlanSzhI8wN1LKqp8u69axrM4Ulh7y7SPPK/iy2Ajh4A5p6UviFXEaCCzg
WXPQfkl8oOWf7J8iCIGYNflgiRBH6j4IMZrElrl3H5SRp8zp0zQGfp7ai85RgdOH5tVp+TcbgOLN
CI7YffPseANLaKkkgxQfh1bEEQKtx67yjyOOD9zPCNvUyX3bwbdG+QOziTiREz73EtqBaihliZeQ
QVOWZyEvOjGv/hdi7rlEsWnwsBL23sJ+MdrCJPfbF/t7yOw6jwaTPUoLHq/FpC3VknSCK4ANhkI/
tD5C2w9VL1i/RDFX9DOcwRkAtGpt0pI6Mb0CJg/GUvJ6wjWP8Jk4cIP8pjWRJIftJuxh26N5cBSQ
Uvvx8QAYyYI6KKdkDyBgQUXkLNpiyH9921aQ0NdRQ+Ux+Nd3yPgHdAOgm15JmcVJJYVwbHUYRT2y
Bxl8afb8fFVQ3IypDmvQzVBF3W8K+J3S+Wf6Jx82b3q8xcxM4b6coKgdXW0BP0pvMZXgxhMNcxyw
PmzZHMgxrh0B4noWyg09KywmtZXrCO36Np4fT1bomURDW6p5t2kTnG2zQ8kOijKEfSKDSAR4Ny0A
SErdrTfpcaVu29t3hnr/fV5UdX5vp27N7TeECex5PPKZRtRnG7R1w0MK8HHRGkZJFMfFGSVkD4nF
5NFInInEKrlOhlqovpzKrQHGxhbW/VCiAw/zouUL/B6zOTUNdrgYTnEG86QERmEe0FKxJQ8kw0WI
4jCd39n30J6iaqAy6hUy356KmljjZw9MUQaSd8cZsMPIy08XtwclCGvlFKhiEb3FYgFn7X5yHTYz
OKGwH14QNfRbBBQ37ShVU2jw3fN+QzlX4vhTzwTxsrTXgSsaDqsm4BMT2OCxOkRZVU/daa5TJeWb
qY2T/ZlAojfk1NDz8OSV6ccOmi5UOLPMSCf+8mbp6NenbaOOAnB1QogohkwsmdpLikx3FMl8uQZG
KUA43kaNta8PTAqh9CfYfub790bpWvaHPULjdMn8jSUr2hfksgIrgSW20EBJQ+47iZHkepjr7fKA
Ya7X9ldv1YFV7fqSHkSXk67o6bHJA41/nyP7/a97YpR+8WUiEksWlKeWjE4R11leGMNnGxqN8Xfp
5UwrUEvUYXY+rskJaF0s5v4UIbT8EjGMYSQDJO4sNRBcoO2JSzcp1FwsKPyLh46BkRVhukXQCCwu
4ISGzdBOtpFT9re57Ih4NeMty2z2kSnUYsGsqzoDD8fqLPXujiFf25tYPzFwbEeulXrzza98b4iE
tMMwOPvZoWIyrjBoJu3SJ3qI37wMyvO2AZroUlihj0Y+WNDSvEjvGeT7BWU/rHWj3Sut4NW6BKGs
GXpHOolC0umhrWwV2YxtgjwaCE+pvifE9ZbO5+8k3DZS0fNAWTSsmZSjYJFGCUFPFqYpgUQDC+Ol
YtcarsZ92Kn7Lpd7EzQ+rZDNWUTvYvjUfV2Pe9LnWCG5+xdGyNRVQ49wr5Hird9VPfaNdoqG4wtR
ngk7lf8CCKUzETv3hm4LBakA6ZCveyfeiXDU4HJgp+wjtH6pOz4cPC2bA+3AQ/Qul5iLFaOz7RQn
xsl2hxitb6SjX0p4wyajPn1i7t1MMoCJiCczA4nTUkZ2G3ifXnxkDbeaNDtTO306QfKrA+6liBEa
XcS3VmgYxHXU11EPZgv6MZxrxQc5e7bstEiNfRaSpdNvrSJTCoLri3xrlZVuy7ZeA8lVPRuTfOEk
TtczFrrWf01RzvQrkW5z5ItY2HAY+nIiEmmNXyr5YFZxn8bRAy1RJBazF0ABuUtkhS7eH6i6O9eE
d2VijQL5P5ZX+SFjN9FO2ztl8+IpyyPlo8Ss+jCf8KjcqTS7uIgdKtMfdkepVE4R7HdFg0Bv/87G
lheWt5mjpkZXFrKVNoMm+iDxEhDieKDAf3SBG8V2UdrUPRO9syPjkXAt2+FZo7i0scunoptFLGiM
4TKMFKsKqh7Wmi5BdplTnEsk4ThNBUk1VBM7Lh2F1qirMQx9VKefXjLECZNBfLKLHb8YbN+vZ43a
4ahK5cpB/7/W96PIqkkV5/e2sJgzUifNSN+WjQ5jgKS5ATO7iy5oeScXEe+3HXgXAnhsPj0ZzRpt
9fX5yD5YpGhBn1UrVywe1Tf1Fl3YvPZNCLMuzFP7Pde0HJy3f91K4hv1tN5tqTgi/zTw6DBiiGAn
dhgwB9IvjD0A0sVGRpfDmnU4v0FhxIDWK/J4mVJfQZmO3Kn7/rDsVYWaFxSq8eyXSrgyDtKkQnXG
8UrhBmwkyHzTNFNgmGuSkV8JQiCQ6GNqdY+sUDhdZwEAjVrVQDF3JQ/OUfh7sGu8n2pivCh/IQxW
MVhrwMJjrEocYAcPtuEnIK89ZHRgEhpsuGUpL1VkPJhM1lcxK/KAbx+thwasomrjDV6w4HMk/fNd
z9aQHIbsevb0HLOFF3Veu7VEZoljh5UNVsew+cVk4PBIag2m4AxDiQp0j5yK5f1HI31lQPz2eUMD
qqBkcfO05md8i9SF6sfMC82s6I+pf2h0KbSeMEt0Q8J1Gjc+qKylgl4oJn/NwvkwkZvpsiN9avdX
DgC/S6taDqzbMD2rEsXmObys3RsdVk85R/7TfmuvC5IA7u5m3b+Oj0vtKoo+J4VZ6x6UBcE7rgCP
cblnK9gHIHk81Htgr3g4xVHlA2zPn4bLYQo1tTFnYP95usGcfzfxLv4bC3LwvTAQL+v5Q7crFMAW
Eqphj0dv6SOUMrDkG2lewCBUnRQ+wCiTji230Un1bx7Q3E1j+6RarY6X4tWZoN0AwFyyQKmbyP/I
KpEtD9eZdL2mGaNWgJF6u5rizrhQSGMHc1depcnUGvi5UGS9MKi0hpPJHFoyccuDlrCTL2orhAmm
0IFLcdPu1ViyJTOAWRqI1IWjVFZyLhBed+i8N0toFoxtvGjVrVsaKn2GvLeJLk8ztuNaaDjg4rrq
XSaXIkb2VMirZ62UlKBJGFH/TQe5wJ8DFQLtZM8a918BPW7b17Y7bMOQ+nw0h4cPcViuwqCuJzOL
WYLpsoFt8bngNjhw1Qo55+YaPDAtSv+tiOYNArzHftxr32XZ2cEr05Eyb67RhUCNoiNUMbyU56mP
IPFkBj1DZq0AQwj0edTpS5QZfSfz9Bikd1tN/89ixN9rTxjd2pu9J7eD9TWF5ajLRzuRIE9mFJNm
yh2Tb4YcoZNtCIzYH6ISr4Mm+SxyuWtazdskzu+ZO2QE1ViI9lCBCtydzcoz7dRIEZ1KLRPfAZwF
6KV2YKweob8rDls1lVPwumWzPNyBdMufVE1WPFJZcm7E37KXnaArd9t5WIYhp96mK2iVjl1aiEPh
sfUNiSsG9yBKKycLuxb831e5waxFR5dv9A3n/Ef9JXgGRfnyFnWBNYOF08F4aOj3lBwoVhPIcEOG
ctXwVFUnSJVR8IdEZrbZonL8tzGtDbJRRjvLoZkuT3beqCY+kE9+zNSnFG0FhZbRu3Z/6c838+xq
ikez4PnvyED6xaHMLkqRfynAElLkgDlE+vFfwCnwoboFkZidqSC0KEAdfhW2W5HAIYKZ8w61lzrd
gD2wOyA2a/XFfU0t1qicv/Y/UNshtBIPdgJBcG/kP8XRG1jpcF62HNpNcQ59SeH+1bBDVEtHKjmw
WaXeLHfvCmsmkO3BScob193z6W/NkpO2hhJFd+dxsLGliGI+qfiCiO72Ve4/aoJaEXVkG9DGlkY6
WGn6dt1XUC+xxDS63QcOY4NkbvHXPob2wg5tTnEfDVtdA1W65LSB4W6YPRzMx5u3CucZ0UdMmP3d
1MF+q/jUg14YIFfzJd9Iq947fSl1ET+mBra/R5Hf7+QtdwN88ZOs+UMMkLxxe0Lv38nOHazbMQbw
cRJ/fzV+q/1zBBSYqMxnuFcEXw2v4XSzCfFrrD2ZLefp0rku3VwroBSjVocIiekz964iw7IkaGrj
GzC8byRv9UvgL1G/BTZsgqiAvGCpvOV+fOem9qdyxSbPXlI9/zjrf6S7Hbg0SYLu7GSskqoi5X5P
yYnCKxJL9IAf+oyD89KMpnlX7IzbQ576CtiQ1gCSar0bnHbB8BoFiShR/KEirC7sy5nKxeMSEaW9
fHc0zVOWVgeFXkHCTG2u5JV6D4qhmlZOnj+zQJt01bWax6uuLDxRTcfIi9ksOukmsELJl/w9l0OL
LypHq58lWOzhmB/vbGNoFbS2mSaignMTmwlRqARBbGqnbsqcXKdGq9lRRVlrAfrrfrh2/P4k6D2x
qt16PZIrEkfgkejYJ/4unpaXVTH4R0vFN7h/CkC+cVn5/bxSFwgO2boGso6TSgv84aIAbSsVHXCf
teRSZTZJnVxiaNlDNvLiCvv69D9GaUHu707NT6aR3P842ZN+vmBpU3NhmF9+FyrJAIFXVxZD9B/Q
/cyAefOqUVRFmV8n0gTO1UN6hFHmxMmzTUFbR0BWwsR5Ua0RfOQ0li5/a7KNPxfaVd8NO6m8yucK
qcU8mJKDfDBTi2WsI6XfoyYV8VBdABsmHDNNlWtCf6wcWzceBdWFHdNFCbqPCZpU/lpWIPy7oVp9
H2aJ74u0nuucDilI5O8mV4qsTFg7cngbzig4UsBuT9F8JthNlzXez0lLI7ctPB305ztetN2QtsXM
lTLbNZNvWjis+ht5nrPq1eY8YSyg1pPgLwPQIffAHSxd4qHOLiQDDw6KJfnlYIW+aNopz9KN0BZO
spOrCu5WkcebDkToih3ib2GRTSGid0cZMGsSCTAnksNuGwvv7dVlTqLTeCBRF033kFVMl4PQ1vgg
d7+b+JoB88LKDvQw4GvW2b3OCO7l4WPq77LiNM+KmAEHC5gvl1DfQrEOH3WxrFksAl4NyOcsodxt
ZpfNRsZMMKN2lOxtks2HphNAlTGHyCTmze8jqJytqjMs6if7Eh41NCh8Ivpx1+6g1pKPJ3B3ojVO
XM+J82wmdeIvn7oE4lkaj9RiSIb7WTajZdebcddiIrgduN84oJPkn5L1zYzbQYEOLpzF7pCnBMDd
KWkScWWDGSNyLAiHGAzKXsbDEJaFm4jtsl+GBq2gJwyct5pGmzHWzGxBj3JwWQnwN1fMShJ8QN1n
jPZzyudMP/CARAyc8U1oI6G+Z00yX4ZBkrmIX3BAJlGty85vo0cSPZqcyEpV5tlLc+etSXHyRpwK
l3zSR6Nf+LQ37MY1T8Ub7Qu3KhtDYNWDweOwvBNJajTnIhZ9CFqn5RqxQIAFPFe4KViEmIu+aZ27
Icwsuw2/nKN/WRUYVJprnA2LywxTAE6tKew14zUFcLepZjVQ9joU1KA8+ZqN5tKIWir0FS2Jm4ZB
DGDkRxVNPODS5CDpOokopSCJCgHuvroMV19CQ5UOmGrAasbcJmN6gfwzygL5gE+mTgJq1A/UAzto
S0p64bQ+QYtpkCpKWfHI2peznqq+fl5iEfdopx/nWoJsg3JlUSBakVQ2vKiPwirnLMM1uqC7eP0U
uoRlLRoffys4j6k79wWIGcGIDodTPoXnayHRP4UYL+p85QXPeNjguST8mY1na03RwVtzzUMGUDAf
XF+MbdBNd/9eZOO/XdaB6fLsCBuUkleZvRrV5Sf339FYcSGXcX1DX7UXapEE4F9pbAmCSyCH1QPp
E5vLTTxaPwRmheYeYluxS2jygjdYbNJw1TKxBP+xYBsvTun6iN+1V8NiDoJqDlKiE/ba/1n4jxlZ
HP+ANTd9mjJbt3sflQjSjpMYpi4pxQVbOSoIGkcFGLBxbBjfVA5ZSHaYNmp0wH2eGwTRIcf8sCWm
rzlNk7qqLPG447YaqQpxgEnv6hr2e9XhLFKvqvs1yJU0ZuZv35c8vknUj96OAP8yfVV4DA9MC6PX
187qLWAy5wYyaMvdcSqIIITi/teYVnN8QW+3IXTa9pflUcGdJrXZTYMkN1lXjysUS4b4mmr7orvn
EHBhTNcwQ6ELAOZUMyzHVJqWz2YDsTVyC7HDGCNe8bFWgNBGkYO5DZvECEoCGWYyrMSVeK2deL0m
wJlKPHv53g9d8mSwVcvL7e796oJFrmz9u3ly4GXH9/7n4BQnk8E4iB6K04ul/fl4ikF6nXutsFx3
EFcqA30ST2bdSFsbCOoV47RbiS4E1g+OI/Z0mJTkBm17h2OyEJYyKJXUgWwEsj8Hi2hIy8jWytw1
OqAl9qSVEcGvs2eA6Fl17Z+1j0qTZ9PMVDVMH7P5l1nt6gFMmE5v6Z8fivlx3zItHKuI0VOFrpik
xUmEHcDUhk+SProtEegF1besBOnUbcZPA9xVbMTTOso32d5p5aIV1hdqyko/o2nB33Uv0QAqJYFz
EyB85sfk9tAb0yKcOAYnFgcyj9hnNTaveJoK6FI+AvLpVUpYs+hREZXp3i4TEU/I8vcQPI2DOhtu
aQT56SzBB2/quJUViDlaOY0lbN6NGyQbAc4mYxIWym9aaQuWpMUWjs5Oux3+cpIIIoHpOAD6Gn3Q
76PpLfM71WpPcs4dRX/6R/eYhMfrEtmOn2zYL8Jdc6ltOtKUMHTIzJmcxp6+fWhS2/0kgkYOm2ke
q3dpuc3ZrbdDfR5r9UfcNgFHeqrZssI7aItVzDwnkkKB5sLOuE3qUt+AijNXdo6bFsJT7hsTxh0N
FrWu+8wIowDKa+xVybMwc/NIRZL3IEKnQispl+QTAyEZBhNee2IR3YbABUCn9n0EOfkua+YSrNLA
5nTu/II0yGgwWdqF47YH3HPfuaGankpzLnZ1E2VkVen9cr3yoVKK9FuOnxs1GcPovodndg4Ee+3z
tAvQ2FuRqsDn4Lieh3hUSl2S+vvAzU/TUKfUwUo29ipfdNDNxbkOWqB2x2FdUxMIM3irQV1gPD4J
npYZxi9IO9hx/QIZZmcydSRCFLBAZsahAL0qZiBNHDTnbzx8MLUYWAPe5Q152epDgGi6AtQiK1FP
Yfb6Az49wN+b2yoRv5TXfZ1nin0GaYSHb3ts50al0dADZWu1ZlaKOHi3grcoNb/z3RXKLHUXhsmV
zedaouC5a5KnfVpkGpp143I4Au19wP9Q5ZMHEw0HD8/w7zawV6bqTw8iQ1dQ622YQRoTPerRCK14
oTDNqTkK8aoPlBndjUWa2h8RKQmL8t6RsYqvh1JjECe4vV9Nu/H4JbN7FvTCcAhSx6UA1aD8XFDt
vRiP82vv6mVlkOByHJ1rC2V2iie9n21oJXr6bOmQ2/8EEJIgtyyLXkWxaZs3+R1+PT03Wmq9bu29
Dv0Nj4RxujmthNH+MGWZeULf27beQoGaU5EUNKr4E/XkjjlhkYi4UYSdTehLXnI1/KKqI72J24rE
vknnA4woR0VcQ+d008+AjbDgIGpZ/TwQZohiJLrXc62GzvGowCpfG1FBULAIm2VIsAzNvV8zIq+q
A1HnzjZp4Luj64HLz7H58C/0mh710zWXkt67S5PLTZRwMvwNQbdstLj4fKKfjGMN2WR0CxxSQ/8j
Or22KLgvCiWkvWwMr6XmzeExMU3w3BImOVFjlcWKIVfzUdm14Vh1RFSARkeD+czuYsM/BAZQYvnh
7Evj5hpECINoSJrTwuWxnAw6a4ZiU9EzvZVGpXjGM1ZrdDuOFOsEMzFMbppKVWpFmsLRgc0pSWtO
P+IXPeuYgvTtMsexQ+eAkNPnjWKQsS19bgABDpS9Fwu7nDgFxNQS+y2yykozesMcq79TBDR4/HyX
XxF3jxBblP1tmqaNabNfJ3kyktcBGMfKSzF9GdPMLKN0TDnHsR27s37lODJGHaHe4YWypH79lnyv
zqVPuVEjh99KHE1XOJ9q4EsKBy3Xuo6ahqJnVox9DcA2MGWVDyuwmFyPwp0C7bpO/ed7Tpm/ASp5
2PZ1jVn5z0R/3LnqmRASJSNGm1BDQnQXRYlaooU0aMAzhbtlNWksuojbUSxP2Bjy+hk45kPdCCoG
RgZtDfnZXma9E8x8iQ1oIMIkxEBhrvjahbtWVfJf+SoFxEX7Vv4lofOrYi1pE2P3mqOvUVK9X0eL
CygbMZGVQ0c4wW0Kt68CkiBkWccVBc14DOtP6BKJXDaETCCYe6fSQPmmm7RayGOdiOatvuVEo6OY
p3yXksfxazZTgPB++JWxvOL92oO9Z53Bj6p4FFjvWsfcikXMIrRYbTb2cJjX+SX1RrBmdqwahBjK
NPJqp/Kpkb3i7r5c20nhmZSemS8l5c4tP/oogHxFzZYtVC3ZqQLONUdoinz4AZ1xTgmSHiSMUeM6
tHtXLuZfXVxe4fcdVI7OyAkXYqGGyafUc4N+WQ9LwQXkdfNUAx7Z/edhrssgI4548mBmk3KUPcsS
jBd4RvUusxRkNoWh/w42WeATkbhBYy7i93REiuuFxXR5kedGLPB4YOZKa0C9gVcOkVRVun7RZMwh
S553vdzjZq9ejisyAjDRgjOmTMS/UACW58kOC7snXaDQ9KCyOHx2/WIuTMjIr+diuxkxb7kSYTFF
i7SXMZHzso3wGWOd34crWgb3cs7e2m3B4JC95LQpSJ8kdYRzqD0N32Tuf9Xm0nZ5OXF3renMLAAP
iF6fNnFdshTg7VrWdx59DDviPokCvoocuLZzO4wa68tfs5Jd9os3JcBPMR/Us/IQnX2crPv+slm/
h30H9zWtCVSne4eExUI2vaQTRL0DRgVkGeLVreOacdy7RM5gTCg/qNR6bs9P2EE7fi+DId0n55xx
MaY0xoKjH8SBTugPx0hVaVOaL1WYknqPnIR1tdkZYa/gx5ZoMNuojpK+KffDfkChGaI/uTyEYoM3
p8AjEtTC5mkPGf/4IGt4U4Wt5NKlBS8amvjouKHmIjERJHqvB8rg0VuyvxEGiX0H5dZ0e2kEEa0Q
/EWZEeugqFlaqmoiw3aDsUDjEJnzU8TM9kVyfVGHtdK6b6+EXPjcJqNWt6LHEEr637G+s2BCjqBB
ewgt+FAJ0YmhtVKPTJ/11YTNjMWlyzH4Dg1j1b4gYYW/CmE/cgI/Ghw/pjXlfWYnGA1FohedTjKg
Umx0Jjz2+wLQEU2NIbDcIlIbOrRw2cOzHsw9aUYts2GDK95ujmHrKlAIQVaG33YEu9GeuAp7MwXJ
DKosMjmV1PtPIUinOnPndBgK/ijOG0S+VRIRpKdXn2UbX5k9YhvV9fjQ94iMVEh4oedxZzkb7T2R
jcoV6tXh/q9GUD61ykqoDP/r88AI+OlrbRYu23/i5Gkj11r7/J0/NcQ41/UYRlSiugStPslscqV7
dyilZzccEtqfmP0fECmTekq3xBcrHG8crNzlOfgVzkqvQ+XbBs/fkbNGYlSZsMtN+IIf0ZQDgSQf
rtMUWxYGEAm6ryHAEQWjqMmSbBRnrqhSZ38iSE0cELU0j5idl9jWMLLXfvLgHiHeaDdTn07yE+Z+
K6PGYU0wbTR3sQoAD52gpNzNhtnMt36Qj1oYqhDtz2wNuseHlsYphH3tF8iG6RShddI6HVDNKBWz
A22LL4vCdMsAklSzrwYbH18xop9TNWQlDIfBC/yFLnX06EHNrjaCubG+Hq82ZKY//Hp4ZAOkyG0F
S7RsHcYY4dhAcqfyfzKvL7zXcIUs7m0PleLg0SspjL067MWHG4bhv+68ik0Ud3Kkn1jVwPx+FpZj
/bwZj0Jw2FrbgjcPhEwOcuYnWFX5dgxxDk6QM2JM61O7kzscT2eR7Y0SUYCoFPxmUfic5JbNW/i0
e95pt16laH4hu3mOxABn9q6SyK5n+P+UP5jBaBpO7F8aISdcqN9BzACvkL7gwIQJsZnuFp3itTqX
WtkM25ouOqLqfCgd/Yx/REfWxgFPRJjwYS4Wk4vodjgN5ON7ek/i+W21Yz3xVIkaEs9wE9grSnLA
RdJ/FeGU6DSUVHeGyGz2A7BFWDW+uBRVBz2x9qNmIUvdaAa0I5Mrz4Tyra/Tr5c8ybx/FnW4+LZQ
nvlCieq9rcXAtOPS6PCLuLEsjC82qObYpQ0zGBDo0KvIaR1Sl0FbNFErWrKWI5YwQSR8pu+HpsOL
nUOZUypT8MwHtLpiAgEICPevq2d6TdRRx5Syw7uvbyQVjpm/RWLYleDAAQMmbPDBM88tocwk14OO
ZqYO2dH0JYGzyRVNjAmbPN/10ptFftmpCN6RZ/JEoeJO9+qNdf+2w6DnInB3uKm/JANs4hVV2Zz1
UrjSvCzb9gFP5b+v0p1OHIGYG5UigJLrmO40a+dDZtKddNG0EkjSIz4RqvRAmFzr5PjRCJdnr8ch
KpF2RLgHtjjwAexsp7sGqe4VUCwwMX2uUHacKKERRD4razuGwEBz9wxvTH+wWI1Nbo0qenZNPUuH
u+BTrQAvGId2VcaV/jPpjjs9IKbehwMtfobSQueb/ilNWwJIK7PwHBbHBQnj/mrZ+z0UntcFQuNL
jHx+FVxCv43kRK+Mft3180Mk6OhpmGD6ay3cJ8L9w78Ny5tC63AA7RunksDSBMhOgnrRCbXwfCbL
1wHxu4Jzi/MPN1b3KOywjDqL3q5gi2VxuE15bBz32dft/KDhtdjpJ9F4sqCIwyw8qtkud7ny+JaM
xBD3vDEOoqGFSdwZ5WXOk+dTbKU9THfFslni2IwhvPYFErb7tz0FLjJ94mKLoxYy3If0WPDyQ99D
Hf/PDdAZVoqXLdfDltBvvErfz/g0VlqGoCJE4eRVOvRCVfvZ6esGGAHp79c7/rqphhFuPmMvuECj
TgXDyKfGvtQp4OnX8Xn9aflGAwP+rQzJUVmHvdKyS9HbjOGYJrWZNPJ6GERNt7y+BTrvd05bHiRC
6nxvbWpyVnQ3xGAE1C7mFClTHXTu8KdfZUMTMI7sUZq0+FOXy+7tkgC2fSr8t0D1/pEGCnF+uBU/
9JJMYFcCbkUHG+AfX6JLApx+C0qZSQJRibXJpKXUIhXBE+g03SePM9J66+9m1hCb644LiAQOTW/b
ksMVJBUziIUw9I0Pet1bKL2divXCaGm91osJ1tuOiW0y/ccm0XzQG6F3YbEsQC+6MgKJ8ujSioOk
1isHF0KDg4Z7y0efDftZCuD4glsKjpRFHkNYF7TS4uBCkIne/faMXLbOmhFPujBE6o5p2miZC4uy
hxl/codIoZO1sO3deqkG3cDdY6Y//c8W7MJrsWFPPUXak1n/wcQN8qWl6PePLFkXczD2r9t5bQQZ
N8qQq3H6L1vrWL7BCGAYOIkm/WX82rJ0wIEV+sK0FSXfWydhOBsGuJfDIvXNRWWB/fQ+SpwnbAfo
yT/UeFIJM7Xgb7J3TG80S118Lkawhm8D2CAfcvDYQDES9SQE91pWPBpylQQbRspGHi3KQDeSz+8p
hoKiSQVmHpGaDF2A84SJJT7mw/0SOX5CsnRkfeHyHv3cVWRTqcqeO0csrGHHLurTXurxeelvjZ+O
RIHkqlJroNgCd+LwaJqdnn41Q1Z3FUV4hgYSgMZlx4PCdMpljj3N1whMwTs85K19DTJupXHWBbQQ
xDRxPpD9LBy/aHijagYALylvKJF5/JHMRe90byedayrjK5pkn5lQNxPsUqIn7nK37VuDqePnsXTr
Iam0r47DBnrd3MOHh40U2xEjrhfgtm7M7o716K6ErBm78q3PrGqcfujpf01TynrP6Qkzdq4xa4tu
DcoupBSRyTyNYvHcbbyXtUMcHfTTl902jRCqfFJoqJzAEB2t6akdQw3j1QtgAqZK6wjNmopdURYK
0U8rfjE6zEq0IiRNQMdQBpIkWr7eUBOEgEW3GNncHHD9o/T6AeiDIBrdaix9YBREo108eM6HF9t3
0jLuOrnQRsilbIODCeCxixTsvvmeNs8OVkDrKpP2dNxUr5YO6y589xbRHNz6pS7rggwYT+opFvgD
yx5mYw/6C9oVVrKe2s2ZEL3h7LswYYDz478j4gvD9yTGmqFeucIv10IGQkBDVO2YCDjFljd9tjZm
ivW6yafkdroXGD0wYc5i4FKZjewhUbEbBhxB0dLyHvNiid5coRn0/yMDKZc15b9BHt/2+8FmAIVt
RGDBEStCjXkZtSVQ55+Hezmpd6QBTc4hn8JJHt3Hd1EfCVj+Hw+G6SVIV2RYvEE0etjtjJH5ZU2P
z/Ll3/UPAJLJBW2N9SCcAZIy1DuCU9WXxWVcYSTGGC0srF9jg28lxv6VmvJFMGDSUCzqqT0B/Dhe
gfNeIwczPmrpobh4xveWnOVUwuwzFNDdOVCYfDtsOO9T/MYzGfKbA8CQRsnM8UTrgAieagy2YCXs
33mj/1eetTNpCXuJ0OQAGsuPHB4JXH7x37ESxhRFiu9ttsIeaMnQbKPmbQu8+DST8CBCVTMpjPtJ
c6KKisbQbb40nckTt3fiHg8Vt/sUgtHc6M7dlP+d7hjNOc4vfluC8M9yED19IPLaGf3IAJNLTXik
0Tgq5/2Zo+npbBTNEDggnUcOeqg/RCDbyCs9mSyGSxWBcIrbMxES+hSfqXxocUI9+V2Tf1dzgSVC
C816wutaRyBQLKmDQgMbmf2LhMGn8qn8xuPZWo7VnlYutcpSGCR7yv6pdviZRL1Inu7mNVBXm55e
t4HsvII3HWECB3J4NZVHyRVssR0oZJr+sa3iaCTfACN+g/YakuN2NQasDne8EEfOIybYvUJde7kf
dPOQstbr8tzxxwQ5gsDNOMZ0Toy2ILRckHA7y152xChThUexYJmYBUhPjaONgc2d6amR04me/k7y
0VJe+pr71xtdhiHPge35jWsw8RbsqIgPq4gi0P99KbHuq16KCFun2R3SEbIrLiVXxDYqmaxYiPiX
TEjDl3Wt50n0JaMOTuQAstMoTQ+MiLQd5ku9dcGRaXieI2zFsVCte3UqTQb+dDPelhpNYylwajDx
n1nFMnELGvb26gc8G1fLmYkyEZaZUPhaHNuWZi2FDzWXbdlVXocTef4vp3kPbNGD/aARrjiW7BL7
CAkphJcDaz8DVQjPdTJ5Jfi4CtSsQee4Ol7lABBYA2Pq9l5PX3VRKb8zzAC2oQSzwQ98sbNC360m
UbLQtQojz4Pmxo2KhEVEs9Zb2gJCJ0/0c/NWYk0mGpW2B//KLxG2mZGCfnNO1ib+GJvW39kqKHOL
I+GG4z9FG/FzfB0XihOYn0gjFDD4mLgBZj+/9ak7ZFE5QsyXdUBZArO+fuoH9WJbQQ1M+NttDu7L
0Rb/nXKrUQB87qX2nz6hn/yv0R9fVeCHvvKw5/L6Pl0BPnl9cGgO9oHUHvugeg3hdEF9PTKnVkct
/zceamocPDBuqlmNlnOkks5y6rtESFvYoINLSZlcaVU9TXE7EmM+Gy4ZfgU9TJF0B6Dn/0UxBnV+
PvcuGAdS40H3RHeJl3sKGOfKc30KEimCiDBW/otV1ePf6dndUpu7R7jLlmg7dpMpKY8eI3XRFBDK
Wgvmx2X7cmRrTfhoh+gKcxfHlGmHMlUpBKq5/MUF6lu8h16DQdFklxdw9KHo7WIGh+szHmqCpPpp
3U/J0v5svJ18L2OhvfEM9X8os0pVY6a2unOH9M2VTRwQUve/+gY4v4+MCXKFja7YE7qdvlh3b8JS
xe2Z7sItsCZiu3L9jihsI6KSwyps/7kQ4YKcmOEQHQqx2SYXqgldH3Jwni+xE8XjEYT/p/63NKpK
9HMEk/XoLIhRDTwT4IxvMJIvmuPXqZzyX/E0LlqdTbenl6Eh1yFvcLEjfDW706v//p4HR8N309BE
L54l6OsZxRtFpVdVc7epT/9gMNPmmelAdKt3ZzzoQucmtL1SfYcx3yIO7bT+Rfw5hOZKL0M1w/Rt
7bc+e95+kDg/FPCjCCkysDTNJtnkT7IGWdHy7hbXdZMuMXFvH0qaG/xwYgSj4dEpkxGRKDberKGt
FjNzJFGEzvGFrC7HMbf4WG+7EYzsHi7ro+DgU3EBre79fOKnbzcbort112mPeo+CKblMqiD6nlUb
z+T8JSG4zVSwGUofIiIwwuTDVA0aU4IdwBg2KPhFZCWDmU8TKhAb25hAJ1+6SGXGswcojEfHNPQ8
PVEEpD58pp8jh8C0MDFU1HKHyHn7mIxZcxsvIBHRThXi4bZ1GYvvEhGmCObpA/w1XJpU3B+jLBiX
W8FFgqvOl1dBDT867BGespiC6Detkmy41oNNUbPm8Adv1IVnbkBx0Pd73DgQX6NiPMVSvsv0CbFb
dOWze3KBDntRuw77Sq3OGar+F9LxyWUZl/5f2vohJboCbstBQCAOnSo+DEyjexeFVxrB7oE8ygHm
GH/l0WKo2CXbv9omNxE2qV/bP0ygNG8htKm3BeXMi7siLHD+bLJ/gB+XdpmFCq8x4Rm0lskLriO0
Eu++bjmkzoceer/oGDb6Ux9JKg/IBljNxCVUqjFfd5JN32eb2GGveehNgzVWHRtyE143afwuxSlr
WzqxOEZoZOp1mqrLO9+bCODxVlBay94F7bJa+waDPGUfCrw+3BL+rayqNmWJSge9dsiNT93ZlAzR
Nd3onycGgaryqXFdpSxurBqIDcE1XJaQNEkxTB2YI5JyYQWV/7Fl2Ur/A/LLzPlZf3OOnfpqnUoI
QUVcF0RlNpOxLHORDfGuW4BjgzebxdsIgWg5/s/K9sY7z6cVQqjwPpzFmT6Q7sCbvgOIihcpKJP1
hrCqlAV37zc9RnhdHcOHUVxabmz6m/hZDKfw1yWDJq6ULn9uMl+GRshF4/Mu6gBfPCyFhD959P/Y
S/0UEWB3/6FWv9KbbJJ5KtSeC5lt9FYxxkzuR4r9IKTgNr2f3itCb5owXrdxE3nIOnezozMG6mhR
mYESFpbcTk7Vpr50cXEC9k3U7EsJnFW//JLv3kO7Btu4SpFn9xgRqzjnWJZhXvCYkNNIFQfreE0n
A6RzqfCopDUjjQkDEvaBqwcymF6qPGUpf9m1L14AR2K2Dx5WT6RV3/litDyAMTeFdaXjeYFZcaZV
UBULxbFAI/2de13sQjC8bZZY3EWb2uH3gBZb331FdiMkh0PmWbhec6GSoML9zNSnHxEaZCfhN6lQ
5xg0kmMHJOvIxOi7oPcf4sGMS21ndBEhWXyDijdoqsz9HbWnZgAbAfyqb3a0vd5p7gS2dWuxOa3E
fFD2ktelCLTmQOjwLCWgRM5OmDF8He0ALo6aLTt+SIFPAOaiBg8eGDaKcNjeTsJdEruBvDxCx74d
X2WpOaTx/cMPlYhifwDLfBsVYyNoczHT1S8INs26O1JQM16bRiSw8i7v7WnztcIkrpAUxkZYy95o
aL4rM4wmhJ36Ag4sNcXzSAer4Zjs1y6MWsXIaglXr/ChTfRLbXygMQ9qOl17Ft5P7w+idE8zrYFp
YazNFkQ54hDc6/3jqssZup0YeO65BX74tN/SVNb3qNBpGIbXIbDaSe4WzPD/UzxJNsXPI1OqPTmA
eQm5vNe8JkImypxmvDy7pm7WLCcQvxZfqMziLDw595xoYDh4ekVRowgaildvhVc+f+RHh4F8I01s
lxZvbQNBM2z7V8m+ajlR1zuAbHXMynzjTMNr+2M5bkqoBf/1sW+3CtNR/XLOzHtp7T4SOK7ETcEd
sK9g+oUcEB5faJ16W1SbdrL3Z5awLC8hELMQQ7nq8JWS+8VvOZutiuL8jS4zc+RjzC/ysUTW5vj/
9JfNfZQtStGZhMEQ5uOMFqF/kv/UD1bDf7/Xfhz6UPEs7Rn41JBIn9RiHquKseg4JI8wzdXt8u+0
CfJKOPFhJnmSukd7r3iCFn1yypxfzvDSIpt0JRcJfMVUcaqyJ5+kwZ0uXBy7UOu4qraGERDkZHcb
DzYBBaspLzEmKFCwYSXG1pZKERChXSxWOUm3TBvxG0IsbqDv3NGemwIpwIUS4AV+290NXIJDEHVe
t85nHgxR3f3fGh/Rc3IyVck2EYINK1o5o0FoQN38P+k9STY5r7jnupC8bOhWaDRH6dRI5xkUF0DA
4yzumbSAm1zHKE7tuuzqs9kv7qmeE4s+odBkX+jrxX6mAwSEQKXRT+EuQq3W5QrQWrnr5xbBZV7c
KkjaNoGG9wn9SEjCYVzpvy4ZLXJe5woSehZYEbgMUxvFT5o9gimNDI+CauYcQP7LWCX9pTEvxz2q
M3aItGX24H78Zhnl/WzDpjTJbWxLXZ/+sHmo8JDc7VvMdaf+VfYWBFhs8FxZMb3GCrhfXY7cnA6w
qCD/5YXRpLbyTEDKLHBFlCx6s5MKZoqlNNvFPKxNI1xmK8fqDAHEZ25SyY4xC77RGY0r7MucEb1L
xSSyXVESHiEvqhjBty0yMMsa0LCSQQU+VJN0RWFlSIRH+iyPqD08lLyfbLHbVqL50vp8qiWoto00
wtesSsw1kj9015acpEAR53S6TbpYoLP2MvME1gMOu4GLE6vxrAB4KCzxIwT2gb4OrQLF7yR15OOz
f1qv90AnewdTozeEsVOkTVFhVb2qv3eN37RWubulcp5wqvb646465Uq0Azva0jVCXCkCm/C+PS9b
DEaZQMC4nEofsP93IKkdtDDOC+TGXt+kmOQy0PGUeePuDQC3HzM8kHZA164fXZRAwVxTVX3nJCI8
eB5waqXpuc+foUA6qtmSKG1XNWUfTT3YJSERPcj3zxymoxbWOYbtNONs9wVM6yFoFKhKs8UXIaBm
fCbASsqyFeNoHIwcckGEpMn+z7q6rIPKGVNvSGb5CpNJpzaoSNZiC7EIC6ljyi4Jec8W1copgXVs
F7d5MPsNgMM62lCUDRBa9e/IC6aI3Agt30+aWbw8WMU9tRyg3uSXM7o2JmodhmPX1WopA1cw/wlF
x0g8gr7J9+vjiKdfQl8lg3ruZDEZU0JaD5q3rcp/z2J6EIje0kX7iPtEObAAqoonR57EEdHVq6yi
Fe301Rdw7a0LFPmKkyGQOojc0kMqcQ5UF9OZVE+Jr2ZrgfnTp/zl1tI0N5GYUqFhe9916zh2B+58
3RWaj2TuixoBfveoCpTrIDPjwkheJnkUAI4fjUzVNYOju0A+xgHKc58dfi8DF5yuk9xw4wzzVeet
ZhchtL4jBvJsKqBGLRQhhvvm90DXiWkVOs+23FowliHE7cfx2NfxM4GOACE4RO4mGTpdfTMVr+Ey
XllL8oFtfEu4ztAd62dNRgSoiZCOwICn+HqX5iEdWmZTHY9+meo52NJllF9LNXrlPbiMdmxeNuw4
I+6vioGOeAiRFeRkFQ0zMKEJTi8wL2msqH1LnyMf8UX3H9kXOkpa5hTXGFABZ1MmJ0swO2FDhxc/
aS6t61xpKiFzhFdlfKBJAmbAzy3x4yuI1Ga1tP0nOXz0ZCAmd18KH2u6kgzoUlWx7m4JG6nukj5U
GCC4NCH5G6YBwy74wEaWOVdcVoa3k9cKgeHjtF36QkP/HdwsDRtY9FxEfCwgfSZ4FOlT9eYN4bmq
2rCXe/cPBetsomDzNMceGe8T+YmkMNEPjxjo9zbp0ZLHcPAc0rVL/vsokKtIjguRb3W6759k5v/i
3cAeoe81WsCiP3MDTF+M8k5FBzkJ41URJ2v9HdyvUJioHfduYQcRbuFptzpajqw4sDoIRKPc6EeO
ehHo5zNIbeZevO5/vxI8dEMPfYOUj0+PLKZZA+nZxL/K50kfm5hCsdSmmpXSKfrObdILRsMcHux/
qXWS5IDv+LwQGkXGFkvEQSZ5kuw+FAjl1U4FMEQ0tta68+bMJ0XJ4JjmEL5cMNOmPTWKUNRpdOnc
CjInDQkwCFMagXg7UWX22Vl2mRTP+f456Ps9nKXxnWQKq6ks+5EpI/AADnZGNas3xcdUnK8d3dvd
KlU9/czgsUPr4tyI6DPNkVWMhKBkdQjQkxRyhCQldrEmFtw5D7AJYuFU40sCWLNvvUYj1s3/T23M
tUlrg5kODeCzF7qKNoDeunLwikJ5gfPXQv0H4PmbkPmv3tXXedVGt8W+mVspkpR/nzqj4D3iCmBv
RX5ysGZyaGziG5hfR+wzsKDtrK4QkzfodjB0MPP8hxIWnq1FUocskPlKl0e6PvyoNPgPElgm7i5z
C2mhMb/ibQZV7l6keegyhbKkaqGY99vCZoajg/fz5hD0XS9NfnGuQ7+s6mu+4j69iMsI4ejt4SdS
tcK4hk5Mokr3sKFu+8ogM6SlY9gWsUaMuAUK4GeTuiBPbNjBtiLG/oxN2pN/CpgOt4tfpdwfc9FT
wEBEefbmTjscvw07wBQAZbQA1mJRdZEyPLzGgEJHMpfAjqOGysNxSsdNZxjhU+RhgxzmAdVoEOus
9UP4NhBGbcOkn+JqNa8jqTm4Ji+br9hASyXmOTefkatP39nEp1HhPXlM7hTb3veDu2DENpxGuDUu
xqaWVD41z3DffKMQH3CGv/YIZClA3CZ2+HSzGvdx/HY6XIZaOJptzLSExxDFoYGea+zVNh/fYcEd
f18kK6uTGo3FLVo5gJvAJf82oNbtbenIa7MGLLJ8nyKlpohCDITpgbN74ice6vFN1rWiF0KHCJbO
euqI9Oi3UcM8CkU/kf10ex9rKkNdndtXix5GGzIo18Ik5PPxyKLkHHMq8z+TlPg8ra4LpuEdTshJ
evQZbGei23wdRKpXgUpvpAdLo8Pynk60b46RF3eAvCCnNLhEecXXh8bpUJIlzz0nS5MXeQU/gCEt
MYaVrmVJ/K4WzVos79U/yS5LognFNsZlkee2sLHdPFl7j7x58A52IcvRoCYUB/xTwMqF0Bwsu/5X
kfy3v0cpwxsWwsNJsJLaP/mqi7jBBM9M5p0E3DhpnXwAZ6Ell8i95OZSl8w4FJEFErJae6qgWxPo
15FvaRD+01Yl7NFNgw8d3hGv2EXJl7QRZ1Y+rl5aeUpcraN6RjH7dwNahqoV+OJHI8UcAFjVoznT
PNvstCTBOaGsK7sVtS1qy0eFydpYcwr9Ru1INlbWf7jlIy0ISD/zY+gN8pu5DkoC4nCf+RPs9Cd6
x7yM62Vr88tc6fRIHv0JH77aochrr8W5zxzmS0g7DFtX/gvC2Lq9kjbHv/t7iHAbEZqqH6kKIspp
gFsoU+zJkW8pdJbFKeQ5hGoVIOBgRcaQq84SJPFHE+pQjW6GMibZjyDCZaEJKWPtsNrTPr3QvaAN
YE1vELtZuZsEDgbqByA1hgguhd1Ssadlbou6pfaFLtsj9xM7dgkEWplq6A++MlaOn0qlcmhPP/Oi
esHyeas4iztBEnXvQoGfnXshKpCMGpJuzTb8DdSeZTO4jBn9OE253sr7vYbxtumyzEKpbjootfIz
nVv+5ZJqU84c1rune5ibMAkrVSWiKeHZDi+rbPoYpDOFkIrSt/RcD5kPhQY8WJhO8ajDIfgy/S5p
dl/JCpVwQ9jU/8uXbil7uUMXKeo90IQvXeCblgnOOsew8UhCEe1mwXVDyvkLAwfxgjaToAZfB+5O
h81nM2p+RxQM7Qr3yIFNZ6Bi3tFu6XWUGEP0mYkvoK+25mWxeYGtEIC1uHe038NTeAU6FXVXu/ax
bsyspqyh/tP80ESx/CKpsTSJdiEJ6ftj90rYBjgo7gk7cLM6Trq3i9Qlrzv7cNSiAGPr/bnS5m2r
xS7o748M9hLvThfzDhgQM7pMpEi3HwXLVxFYBehIFf3HkTqip4VokEo7R8Fs8yqeMEYe/zaVwxyR
xyp8KdNNPPBlNeojF49ebMycQ+3HqCQa5O+EwsjmB5uKrHMQxmkjmIyg82zm8i8Zvp/gqxnDBIfd
PFTS792bOtdTPPIDzcph5pWBqC3Nqf4R78IK0JhKDJ1a4JgnrVywaGO7URa3c1zwMW80Sd6U0f5V
KWIn4tFB6D+/o3TwwVkYHVQ/F4JX5sFcNxyXdsgctVJ2N3ayixzJnfI+RpEsFTLJNBMB0RneH5FD
cj9m97WPUxUqjLlkULfKzzm60p2B7qaY3IJHG4JTmXrRXj+5rQkz4FclRYvL5VHlau87vICudVSR
KJJcQepvm6VpcF9BGMOSwA6s100YQ7QfKlSAd6ntWPse03t2hN51s2u/vhSSocQpl4akTVO4tQXQ
6N3l+f2oViVHAxa+wyK2QS3Q2wboapQU4OgMQInhXNofW//jw1wjrJAf8PhHdma827Ue8u8WGKK/
lLdqaOjtwSId6unvr+vy/mqMrjnZ6gCpDq3vOQH/VOqrsgZk+e48RFPSsLHAthrm9a/UZKJbwSie
YZfHJQWtVamj2OwnbE6dYt2wBWD3lCQUTvV9YNMBNLpZyTZQJ5ss0eBaKgqhv9L+yGhmzQWLSOsr
JX9l5Z2DSINYCVRD70DTQFzoi66lQJBmOWXBpU3xHcbe2G5G7qyyqOGU3YO9AtI+dqovymWhSW5/
CBWo/8HOdt9cAb1Kt/ugE5pp2kUZqUywZIoqTYualHF+uoQnxecJ74Fa4WwN2T4osVYzdJTFc/Uz
stuPWoLb548rWQcr0GehVDdaFo+i25fPmzu26q42sjaITJMZDlUmI4cYrM8mlThixqmr8Z6ukrx8
9DpOwERS+s7sWNLUkeWI9kFNgoTcr520zgcXNg8Wz71CAf/7qTgzrRZGjhoFCGb3/ncjUFrbRVV7
4p2Ezdv5amOAM9uYYWJm8tDG0ROqyH3M4boBZXddcYt+ZQNTHxYD4uLgBCyo2r6CG+t+GCc6y7OO
1YFnKdEwT5Q6we/0nzA3X2dvqG/03479na+lPYEpnyJtXmMSswsZpN+3FIu6JrRQrq94zSPPPOn0
TWrHAqv0qnmRn9oOOBqr0KWS/0dwQiaFxwQ9QcLdYUOk4ujoYXt9JMHsnGk97eab1IuNr5+SKIpR
LeXWZnotmaEY7fSmBD/zGaOee+jjSzY8sa92KpKvr8IZt99vHX2deqgG+cgfvqnKVR+GCXnW3d/v
VYm1Bf+fF2I7f65iNcPFlnP0qHjTG4HShLb3p23r6qTOMmSwQDX5ZGeI34gwqLRA59CozpgQljyo
xONUBjANDs70flSfCTf1wofJTwUuR/dXUTCFYIjl/SBoBnb+7oyOlO+UOPFPiYF3CZI5w0Nuiywo
uRclBtvNR+0aXFhGut20xo24meDHQEr+V7yJJYTDpvJjtFUIcCGG61upET2YAqoaFbHw/rmF+2Kb
qgoccGbChRY913RrvtdP5jTjrVDjsQgXSgSW90mEiH+PpJ0B+R1GN07pHmT13zaR7/H2H0JYPh2U
EQX4YhfRyDg4GAJ+1NvZ/XjMJw8n5nXk8Cb3hVTue1L2ULokUs3GdBeBt53OvUFBURAtSK4AxDEo
l/rR88w9AOz78XEyWuM3VJrA5sAJGcKPTWo/D78erw1UkhBPpGbiHEHCsUcpaXmd9UhpaLM122Kg
dpncRlwZ8uzupqyFUdpdkNqUXUCEr/edqEOI5nsosVInlGsh2uj397JYgtJ9MFtAbgaPh13hUMcy
nU+OgYV6RnWKiplvwkZZZz5UVbsgBj9/KrEFK1OQF+5lqBZMX37qvRNglNRoR7djT8VCu9zTaRG8
1aYVGJKOQyG10rny4Z025+wZX0xGRtp68TG2NmOI8JQO8BRR+M9VYsbQPVz15vBlyX4qVfQwDyEo
BytOb/YLre2VwyB189oqBFfQgQsmR3d2yxMStRgPRgCmT+1OjvwHIR1NzCRGXAqP3EMgyrdSJgOG
v4lGebBi9BWaTl6AtutRnL4twnpHFI8WC6waP/13UlbN1kYELNACVF0eW4ikqzjLT3yCXTO/j0gV
lgVzYje93GzVMS3YcWvqj4z2wMIREXgB5vxfrLCVcFxtVX3ReTip4D1JnBrJOd5CYJlopNPT8eFd
n1eKCruIbbS1RoF1L1JQEpQdD/5fK+MSWjg/xd6NPBwmdq9YGNhi8RgHiUhq6rgQ9Mx1EyDzEBG7
x/fiPOtNXjjWyHzdFAZY/K2xoWvAzAx9a230lNJgf0cHFAbyaXtVjNM91vp+TPrYTgRtgP5qnMeL
HclVyHiX4Df2Wjhu1nA+cypkvuNs/sCVS18/1ls4QTLl4Xbm6K45UHZnYe6hnR8QxbbaDfTa8Jtu
K4mx2vimQ/fKyiMjy5NTY3ZljDIC97Z3e7nWbe4Sq+eAEJMMn55km6i/5DdhqjGPbP4nnTk4YLdq
oM4K+7X5p8YnFnDGrstnAMeqmt2n+xzloLKMf7e/+WmxRqWbZ4oUOJzMM+PR9zq/1Eq0ODO27vBo
oUGH2RXjoTbS5EhRasJux1fQrVNIuzABd8qga/+pucn5EV8CvkBTAvHSNQE5G3sFlzUt3yo9t9TP
0nlSl900VXNiM42/pxyjns99t0Kmsqk5193T+jeIMGIu94p9St6shmYIrlnU1YdxY0IpVK43KDWy
ErdBsNjKdDeJ3rK9L3I5LqqQutFfKwQKXzFjzdgdS2M4RsQP/ZPcCSo59mjHdqdNtAickc9q60BU
wpFGqlOurbTeppWAf5v3UhLJ4bVhhP0i2vQmvDlXXLb+ABq7V5dLiGryRpGZfNE73dIaudKQFmpe
mM7N98vlucUx4bywL7mLgrcOh2YwQMQp0YTnWSDD/nxW5cLbt3B4T2j5bhBwp+UnHQm5uTtb08hs
9PDxwFq9wIWEyytmBJsxmw2ajk2KA65O0hQseY+U6xS2B9hPmx2MVGXuQa3FR+GkNx3KN+vDlrVY
EcdGCkpT93GlZHf0kORCOMZQOR0SsJRuf9ro+Ef1AN27XLQ4S7H8kV41iX4cD4H/qB/ABxoiuZ1L
KPs3dL9FplmLxy3KGYWGwt06L6sqZ7pEmO3ui8rQezkDwplqzriBglR9gE/AUB5mHYy+OIZoXIeH
+y0dkM7r5JzFkmbuEk5JQC7loiz9O2Nd7u7i00YW/1wNpdX30056DBGfFHig3oausT4znzoiys9Q
kKCRmx1LtgEKRy1fITLVrAiDuKTMBxC5XSoKrwmE6+VisZj9bsOSsh/zhlS5e2Vofv0aBG2git2N
KmkYcpu9GRUSZK51hbwipshhDOfylTailxzgeVFOsLLpDio4pW87YvmlZJFwFT2YIMKj2oi7BBxA
5zHhkx021kvEy0ONuDPtgBtR8UV2s4meTvQIYxOUBvtW8rFpjLeu5ZQABeuiKmJq8fGKejaa8Tsx
EpjxRC9TtKnB7m+N5WJwgquCbdBYZMiuTRBot2fv0g2pcQqO2bMpG7eykzLr3qOXlIwsbB7VR+am
lwwMqaB9ReUtKPW4ajLT5FTqmsckjBX1+YMVLrqSWNcZUKG1Ars2K6JVud2niX9W10GtTKpysFhB
fsCh91UnyL/fPx7XaMNCe8vxmKAaT5RvvliI3pwA6rQuOxmzA8UQGb0Bob38RD5qgiHt4op8gxbu
j1oxfKfnj8yw9uXcfD3JlyZ7AcKmI2cFqhF9GyEhAaH8x2Ldfur+jPqAgb8H2HMSymtvJalYo4mC
CBIYFHvPxyKe6bRvscq6ZpfI0TiXrSFQRMfW9FT5a4ltAsRtpoC+QdLOtqyq1n+5jbC5WYX9zd7Z
bge7GxQ5VdJnMEtVXbIiGCg1gNllIribmbjrLoVlza2vOr21n1tlyZ9FRzmUB/ah3gAT1DkfEhm4
g3oY7/6/SCAYLzHf+Pz4b5ciqgJBb44BzXm37RGAsivz2PCwFPGWP/6f5crafcIo/GreOpvw0cSd
v7Jvln+c24awhsu99gHgh7oOU422p6VAMWZdP4sBChpPo/LF1ndVcLW/JtnWAxFb4EVcDhZJI5UY
ShJ4O11PFbXp4gUuKgDz4GYDd6Ztyg6v3v3fFldCvF+E2FErQ970ZTciQrHb0MdOpkcuyxMPXFO6
Bl1s8+pze+C5FXNVXqRtmsA7AVo6U9BaWFI/ug2H3NsKsUnqFvFqPNRuv69XzaBwlXj+LySsIIad
qQKA3Yfm/iUqC93A9fOGD+EFK4MvcXIwDisCSl8EhHDoHluu3dHdrdVsH2HM+uevjPYobGJIN4JL
UQKqX8Tdg58z2h/xu4ppCK8HPQgRMTtT5XsVHKND8U1xsOMPA8QFWs0cXTL3OqME0VdTnwdA/JX3
w/D6VyjcWtsYW6iV5TY6QSK4FyhpV14JqgCd4m+drQ+ARB4Y+w7zIqfqEfd0Gg8t5X4gMNBwWx+F
tWUbN4HwEhWjOEAvCoo53g4BCtsTsoQwAIdS/YfdB9QRIh4yr8c5H2PxRHhTmXPx5n9KSc+F3o6E
I+NT79/LJpbyEj04Ao1GikaPmy8Jgqj/Hc5ibxXvahu+it9K9AY8XJ8iPO3hhkm4dk+FgyiKyTdh
69tuuRjqjVmMh0POCIIagve156Gow1ld5nvmdMVwm8nBh8ADa0zLDy7AsXF7Wqq0NVXpgz7q/QVS
dR7qqh1tWHkpUYm1BIGOnS6HyMylEOEasTtv/hVrqjXR47OrLg9JlnAmGznAtieasg41XU/m7kO2
qlV18vDTiq/7ZvhdrN0e14zJaT3OjQPm1HyzfEFGylaEjYuIQNM1d9d+/MK0ek0bvpXE5S2r2M1C
ZvB0uXr9XRyaSW7qd5uxFgY66zyV3j4vHMknFSu0ZD40dFKOLsQ863imksSZAO2CHTAw+YbBxUBQ
ECTV16SMNcvXu6VRVD920iSmBD28286DgxuMPjL0kZqdoX+qWbvp0pFi9eTiBqOEqsZKZ+/MIid4
i3G5l5Rcu8hfR1DmfDfqmbHLZDtf/uKUdKXV52YFkE+ww23EHPDa7wDpMcTnyVqdzq2sUceXItgd
Z2L7q+B266QK8UFr1a3DShXanfupDp2UXfh/1tqRbSrEJgjQyfM3FrnwJOYoZqLSXFZ+pwM1MlWE
osw1LsI/qgkYkLiY2S2MynQUJEBmSLQ2uYt2tHCjuTPR7ZM4BucVBApTBOGAh/HuDp1Kgn8c/znb
rITMFpbDWQO7psVsUeW2bvOaYlluC7hWEdIMro4WOmzcfKIWFhgDkHc4HgaJwe+LgDwC27ho5PGc
SOPF4d2GyfyuU2S1W5rQzB/pLchwH3YkpudR6m1kRuy8pikz16H9eqaLSqbP7QFRIWRzmlFTno0a
4c07ehSzQ5fte60Kotm2DvxJ3rpng7GicIOz7CUiytihttA/Ls0kNek+xiwADjSgd/VcrMJb9MKq
RMFvV5rCh2U7paKd4g8AK9lmPJDHB3aQSmieXIW4zFEQ9dp8seCags8IcorDBK5W6Ym80uAXs4bc
P9Hn9od3sNk9Apg8eXyzCj/gcnEKq7gHxRMheNqLTdyLhXrk7+u9UEcBEjw6k4S4xEbg65hSTJZn
E0Eu7vRT0miK382/jVHkdHF7nuJwo94/0bhCuuLF1ylFjmVAcF+B6bMz6U/zZ8TAfh6+A5ZgcyUg
SWgvAgO/SFH0N77LVwWdfiQDJaFWm4ZD/4wtIDIJ7uauxSNmg97iKBXEDXrsxqnJMZW08SyUI0oS
ep75L9dNfXMjHdZSte5heJxWY1nshR5IicqmHij+UL2wEdBMIFMYh/5LDUzM5tMIHqyEVJYk2xiC
iw9qJph260PyG0g7wTDPV3RKeFSHQEPsFtNl4npUI3ag2Xu/zDll5QyDPLizV+zcZeRT4uMN24O7
MxJQmiFzRCmuyQmjkrCq/wztk3sfMEY4dlKcsfAYM0oy++7kzPTE6VmxdX/E3auJnLJBs1XuIKH7
M/W5lVNZmPW8u8cKZ4oe2yqhmmwPCBt4HApcqspTkMnsKzq9W/AGkhJmocVw1TaBxlmFgZ8kfpkE
/sQ2Eo0QkFIpisf97u7RsSYzsHlfSOIZmptGbmjjr8RE/XchW9/x6cGS4gy1oW0JYD7EQg/CBHBt
eq9r6sz7Ch8sXxSmgKTMgip5bR7dczVK1k0I7adIWtTYFVtD95+SsoEp6njYSVk4aTd0zsApBynR
1qVbhZbEXs+i1K8NjDqso1/C1TzmUHW5/7c1RxDXEop4MbiMgSAqgTtv/MMS/JBOw+/TpQpFXvmt
iQxeIGdKfUKPdighslqA0b82W0ieCl+75Ie6Eajk/PxFJAjpv8L1hUY4eoZBEAtGpJdb/bzHIfHw
wPHhG/RNjfGqUcUvhzImzwM8INopS4uRVKvKDD36Htth1kqZpypHB56tj1AOnhgwV2UYzxBz5382
NHoPgmrKAQ8PYqcGqt2BfQJ734tXuecqVf8ByyevnPKRIXy5aANkne0Uxp86F2VU5wPysJm4T5lT
viIHOt7ZOUR5QvZ9i9z4kpDsCvo3kdB3zm+aoIH5MEcnaZdJiICOhFp/J0WIJI59H7pkOOJi52xZ
WkeEWvno11YiU1E359FY4VrL5O0ilbTiKtS1N98myiMcJh85mpl+sNPajw9/3wnnE7qwRoldSEbf
Kb3fx/Nc7iFJkM+8/LAj5tcb7EWw5C8w6J6uut5GsEhm2Jgg+HbqD/yVw4oc94GdkeV5H/EmJKat
U11yHXYUBPY3PrUREjsxCumUQrz9WweFF3Fv3IxwwtjMrX3GOKP8mSPlW7lvWP0eGt6mhap4SKHL
a+3UobZnqWKQlZILkuYHk6JkdrcpTlQYxJRTdY9wHNVJ1FaxYdG3IRO0ybELnaId9EHf7iI4frGA
HDM2r2JjPAEm/9rgAwEZ+eb/NbW/qJOb/UaQANAZ5qr6h+K8Oph9wiP59gIAkJKvQhkrQhQz6OpX
HcJq7Er9gMtkbT1nSHYx7ENFRmF+ejuXdG7hpmALRkgwO68vgGzRxmVa5xJTzHOPGxd3tJKZCcVw
Ig9A/k64I5CxtgU61Kyge766RJQXw3B5HoedPqTcDpexmPDNrdH/7e8pYpC4LS/zFQ/AYSev9i4K
VH8hvoS15D0pq3UlCbbQbyDOVFXy8xNCNtlst/l9S5jjiOIibXmUXtUEdgsGEgaYZ++NrWODqwxg
WL6m/yeQApduiypP5mE6jM7+Lh+ZgdeFHyrYxDbDInENlyXV/fjuFfp06zwUHJByQ9gLu65UMDQY
XYNHToiOthpaeoRyFMBpPEN9xBc8pqAp57SKT6JyDZVsBYZWmGZrcW75UBqrfGJsHCHkuyzf28HM
YY/jIT4BzYqwVes9Dz/E6trCuiCbLOdMAyhwltc46/zP46Eyak5ci3ovmKrM3seFBUehzeDmNjsS
FA8kZEB32TqV7ZBbvXeCYJSyV2CRFQDZRDSbxicOaHaDokeBDk+T0DDkfaGVq26CglxV0oRDEZj8
Y5YtxO9IbenrcDX2BCZ0SZ0F4dRS6TMp5sZlgf0qxIGEfFgmXPGp929ITvulkhPxmiYmh182+nXv
kZIWj0737Qaa2bn7RwTdbrqRRq3xV5IfKSUmfgcdBpQTkxM57f25eUzNfZKc2gK7uXzvFX9crePv
upGDxm44qOlWy/kdjQZWNZX7QS5gSeYeqz4JpW1JRbCO4pIGPHi79tlODWqhayehM987ZUsfwIf1
zD2bQCMBaYBOAMLq+IQRhB27jnvK0YzI6/RAGzdyqsd5Yd/MN5pzRbdaojouaX7lcIuyvZWWAYFr
2b62+bYaj5iardpOHueOtoUpQ/tuhvMlaMjgLH47jZO2JBqJt+/Gq3pqqd3gY3eqNwSlYpDMegoE
cphv7F9OCrFuPtz9GgrsTTJWnhkVm7/28+3I28AS4BME0bL5KUzsUU0cMmGXOKWf3Z7mWDt1OTnx
xGYvdHeN88XU4zChrPtmzljk1xtMkrT2r1ImLKAWm2qxjLgmaIOW28w+K3cz3wqunmV4fTqWypBT
Hb7kgmoC0v8IlqTlPsb88meqD315j88w2AFFaPYGaOegt6pBofNU5G4kWqE1QsdisTVEm0K51EGg
kL9FVlY5w1Q2cXrUTW7ThQg4yIcO9KA+FEm6Px95UXF7xwwynqHEhlPtFv6qS2t6n1eBzdL3eZkh
XA6QKbzaAlBp21OKtCogP921dMPMODu7Izptv4VcUyF8HB1TlMr159eTJAb6WIVbaMPTNqCFi49w
Tm3qDona4BCv4U8WbP/1J7l0Us+86RYOJokoVMjn9trZjDOan2LP6FynAo5vlRVvIdr0znc3r2nY
jecqRvigfpANIVtHkhknPk6Jkmh9AGrRSFbXcvNyrFzyo2ojzIq0GB4ft132QG36UArC4+WD/6YJ
AaoHuuDQ8NM4m3APKTDwxlLdGk1pkzKuCWFLhuHjcIPc+mcxGSTC8D2njzYpy8WI9rcepGv7U1K/
rSNq7Dk50KMwV75rPi9xH16A49DVujmg6T35FDOn1aDiSLtjf0I+kclPNLWtOtkL9LdXlWf9aLpH
IO4f48mUc5yc0NFJpahbb0QQBh8gXhjcetpf9NoQXMsQ2VxGsEjT1LfUU6am/HwKjW+TmGRmzPac
2P+XZfRGFoCb4XLwywvtYdKgQ+xZLBmxZ7Zds1NNfnLZmOGM53zUboHDQTACw10a5++SiVGbU5qw
HcVB0US9K5FoV/fHAqRHO1JsREM4rZ/NheNNrark8u/yk4gUaeO1fxzVQoTUly+QW+cyqreKiJrt
M9FH7AFlKwReap2lVLS+6xjXHopBIleV3LiNjzDUOIsdSI8PeiECViYv76bouXz4T3TK/MVRtpJX
P42xHTT1XDePk4wBA7Zg/xeaYm4zlNff4rqPJ8S7O3JNJ/C2TCyP4piA25lJ/1RCdG4gQdvsHi/X
64V/3aQFNTv+Tjzq8jrxKaFWeuiwMVDJis/SPnoJkReRu8hjDA0Djeu9ppQd3kmtvD+rA/i+OBOf
zb/pmQTLSqDMpXMYYa+upJgT7qpgaL9Sn5Nq/QwAjg7X39fhu3nau0evh6XuRFjxZvSYu30Y3wnC
ppJPOZyNNlD3Wcn8OEHjclps8Gw/oAQVaG5DKWNTSiNhfkyFFgw2xbQYIkaV75ifhLwrb18wbuEp
2+sLLp1KtLjm8wUXV5oEvSS95pB9A+uMqeOF0Yn2SOMdFcFn3RA8zD7xnaUGWQWcKIf0fmTrU1Nc
3u4ipxvELadV/9NacPff7b28GkdYyxzdtIn+08AUD/rtXoLXcjPX/iG46bucSBj64LFsqaqzGTV8
Vis17Irra+9wcOBpQjBc+KrHrh0MEADKbFStgAJx2XMxatZd3TD0M1oKNXUfvrwrQEHlSHUhKeAR
Na+RnrIPO2L1CG5k84038XN17ANd/4zF43TeabuqvwlCYCBdoiT5ZVGlZ1aHAzauTE0uOGl0RdEj
rBFCIBdg/FPQpC2QW7+JelHqxKy6n/yoU9tKCza8BL1SBVlFcLJFL0/r2mYGh3T5BhCg9InaoZoT
dn1x78cLscl7Y0EcgCCQYBNm8PkKpbcvUczgFXZOQYxR7TFJ8F9Zws0rgCA5ZUgH7TJUUG5NL7Ue
9nVie3ShizZbUJwYg9tilawGRGaQX4m7+XswU6Pw+Kp7Z/IWIONimWQkaAPep4seBUYPULmXOREr
657LMutaFR2eXbzZazvfsVdeZkEFCy2qm9FIQj8M7rlRW6L0xo0bNdxleXRYyq6bbTeUtJxhkV9Q
9s8meY+Bj2WZJqp10lmXOYZNV6M+uCukYcboBx6RE3Yni6GFj8qX+UTDc4IN+EJHpe1AMY1uOB85
h9lO+rJmyT09a/0Gq4iPP1js1Nf04u5ipW0DynM0lDfRrFMZkzKzgXIXXNhMmbB4C9w4sajo+ooN
eib+B4cFEaptImIytdA1mGbri3uPz4dk1bRhwOdmRvujhvFSsUtgcfaXbsdrZ2Rt+KiSv2Kj/GpE
NVmbfIlFGeiCUInodewMkQtgTirxDjZT0Xr2+/Hgezn1ReGBgBIXJEDEkkqAdhLtzDjaAoPbFP9O
wzro570+lbmQoOPIBT8tfU7edvB3Mp7EoiYY5zLTES/UflZWWLoXNk2vDspZ/9KnV2HMrhVu8LVe
sGNXws9LoBr/905ODoDQOdNMJ76q7tdmn/sJ6jr1G91N9/F+Sgzn1XerqnP/r5MSRVvAa3mAn6Yc
O3pswP7/OAP/+YQ2NxXlFC89B192Iw2p4i/9HaqT6K3qWL5Y0ZfycR6U1QdbmRCRVyQUBAmolDsr
aZfwIMSZtuuC9WbzGoJNXnHlZwkpfJm5urVkET2KgegN6K7lGTKIukG2ZjNUicXkBZ/XS4/ca+Q2
8biTyk2Kr8zquxT6ijdgG8hs9+hT3I9BoYefoqcYbvbJJjZWVqk59WjxpWOVVTq5JdTJsB0hm/m3
GkFhruZlCm9BXLWUwgYnzAMb5qGSlfOWL1Fc0hnrf22LqGx0F9sLj1QuJYxwaPGimgsYANqfxhVp
NtoRPe9AYSLwJSGP0mB34WN+e7QgT/7mFqcMLuaq+atqIIOB9l15tkAVf84Rv4zF1x1WOCwMWIfS
RpjIhF+jrSpWYeCYri+30kA7jaqlsl0KEH9I5lgns+qN5xqi6qlcwzV8Pt922CVmaAe/EeeiemU+
2WJPPfJu2wbSuR1OnPPGv8Z2QWnrvdZWdQgI9aB3liwRkx6GBZ1QnaBZzKd2q0VDz4kOWiVX2UdA
RhwlVhFsN0W/+ggus1iY78xMR7IGD/No20hCObC/QVov09ZRiJnBljuC/miw/fksbw5GLR4BTB3v
KIR7S5aAKAECW/l8c2gtweGt4LfxxChIFmDkbURvJC2Vh4PQN3fWpsavTgMoDXBs0YYYw6RSwzLw
gbCbU+t/4du6k2cjWO42pJk12YHCmZaOawwH+eeEVo9stBVQk+yUS+4FJCxXv6sC1XZu8Vx4Wn5a
hfXxJds3cRTnZqmtcFTl7WK/0oSbreLCjS1egNeYw2MedMwvuiWctaQ29dhXvYHeuSobJyBPkJb5
fthrypF39WfMB4arb8pl8kKyownq5vN+yxWJXXzp8nXVU8kjCXW5ly8vZ3BownTqtXLgUCPH4LZ6
xwIHrpLhF7Rep+L+8s4PLxRH77Wn+LK5x9IEqAQDl+0eAQeHmaRl2VrXz3kr0eNT+Rcxjpy5NW3I
mE5WOmokUxEe0xXb9T2PKEy7/PUfya4A/NaC/uZq+451ieDGj9r9CEbnFU8W4T0pCUBciI/6zcdI
R33BwC6BN7awO1p8eBByQiXIMH1xFEGpz8l4Cm2EIcH+eDZKUtStP1jieGvrZnuZhGmQ8at0VXEF
Lcq3zsYNsLc+CQqF84N3lwueyH/ip0WEfc6/STISouLIV1bwDTgKPBwW22/GMRHjwIXE3HyV/uYX
eo5S0aERraECIpTZVp+WqFmHs62OE49GoqEYjijjdUtEhIdALIQ1UyW0YljA4coLyRI2TuMyRXO0
dVBGKkHDIstvEkZnZ2rP/uYml4LXBSgM2AxieAj5mBq/IXTrWdNnzjvq8Q0sdA+ijE0L6hHHf5aA
ECyn0Rp6wkY//BElRjOUXh/e0fOV6X1oqTb4tUw6a57J5EbYcligzvCSsg1rEjVZYK0i+A46slA7
4wH8RqTHxJxuSMfPu6fsURjMNSsX3Ul0AGf9gZK0tGgRKDwmGF+mjxIx0oqS29OEyOP59fRzufGv
yyaDvb0nhDLd1JqPn7FmdxaTZm5BpyKlYtAC6w2Lucxsz3J6mgw3180yHynytOgazY5z0Ji+58HV
Iakq4NJcONvpfGBxGNmK3BgVbdrwzivHR9Pk4zKorZhZpNJ6ZN5antPPoFBQqoOpc/8XNPiknhLI
jeO7UmZwEhKtIcW95G1dE/vPSc641c+SNRCPl9cOv6dxs6qRdI5qg5tPWuD2/L3mWMFGbGf3lwwV
BRPv0kkJdbtFLVxR5zN+s2l7Jb1h3z5wNzbQ8qV5la3pJrH08BS8RAgB5jgJb9fXmatfrRSl1wT3
o17dLvTYY5x546/qN0ZT/yw4YKPM5BZuxDXAo/eDuYBSQF/Rg8DQlRyY58Lt7jI8v51anaCOU1Yt
kbd9BaGoY/Umo0A6xZQ5XLvtt5YJxKn+3R6gmFXkX296bVfdlntrpOINlxs1+ss8eeES2J3JkzhN
aqOCuaG8cF3qrxgv+Ac8UpEN1s5dQ5cnCqnOBA8EPR0xQQRUdfTFCZUi+Rz5FnigglNnJRj8Gf/T
6f6aQLkHkJVZ18OQqHzH1WvA58nfGzSs6eaWm5n+/XnSGOfME4VNtAlOyvzhGy5fZClLUhzxGPz6
yUhAqkZYmbgy21vcCEbwUjuq1d2K4z6Vr5ngNKqcBII+alpEHjsbrhL5WntWVPOJ1Tj8YCwkDGH1
OItlGl6lqmiRe2t/nmrTh8nnsBnKthCmsWHx6R/nPqDZzEH2CIxsmTF2RDdcpw7oMUqCzPH+973m
L1BqYaXcbEDuqWIGSlTQbFNbZKE0suHMCl6yAmdceIE/6W48945f7+Jqsfn89CJUP9mPtpBNqNcz
8024Fxl+Z17Kbfd2ydXKw5jXsdy+xqkU9rz8bgjT3FbFYaXlnFNlgWsKnEnwHh4ICfsjz035dr7y
YTcL2npjpnQiaTdKyiv4Fyw/yK8tLo5pIx6SHgD68ehIEifyv2npJem7l+dbafh1N/gx31RtMdHa
7Co/VLgsZo7r6Z3B6zK9YPdZsUVN2sa19SXRIz5UJfd/B4QstWJhzMimLNQ9/yUUruVkg4Y3gHJt
JMtujdt4ITvcDVv6j28GgrgDl8h0U8XfD5xUnrqgzZivCeYLpQxEI3h9nSmfM5ewTVADf1yKTWPI
r2VyELCfL2AV9ShzsBdiY4IFjb86F/aUaqh48LZRQ+XCt4mBxO5LPPMYzpgNluxJzPe0PHtyd520
nv/0fG8otvc8rbb9ikiT5XSjMOO+Ib1aLQRRHC1WbrLGmhz8Db0hcSXCyNYtDohw/+JJ6WFJaH0j
31VuK8o3n5Bn0YxvdHsRpzEDnI/tS23CmyMpiWqaTDNPuDTUi4iKQwj7wQSfYLSXWmziqI9AY6Q5
tdj2IAySkHH9//YF79OdE4VJzkw0Yi7FBeUnupS7GFhbuZF4Lfu/ZcEXpTwqBdQ7PBTx0jhgZ9U4
xOkNNjbZcroTXD6OHv5k74FXiIcuIFMkqKO2aVebHEb5hEYP77HKjAKOiX9ArrIm+EQ2HodpJKf8
/7dkK3HpoAXilyA7KMOkUMOMFuH2UsI4T7n2bEqh50AA4mLLjNRi9IcDX01zDHQ+I/EhIMwu+tKO
4oDFMVu9+eXafi7UHAudTzKOv7Syvz4n5RTZVvbT2f7QO2YS7o/cvhS5bS8X64ZyIKzwADS4WVKr
vw0Pr5CPkE1J60dOXOHQ0BoCG0OCl6N/fclSv6PxX+VANwFG37rNWTdbHPd+sGP6CUoUQHU2fSGq
JZrcVpQvOSptJ+N8ts43nlhSz4D3rHUCX3F2LELWxtIpNxpG8lU/Lq2MFlwpf7qLrq82QW0+bsB6
tb9Ya8tIiv4oegfUcU81okaEmhEmSqU9Kr3ue/DSmQkXEVczOx7e/WjGWzCnn75/vQqYeMeCDpdZ
agV0ShjXKu3XJHQ5b0jZHzgKetD1Wi7KIjpExvCoQBL4qwcmiBVUrPb8dM7xlKv9RWRSo1hbAc4B
krwRlEoOivqwfap/B18XM8rHrSoqXb9pdhNJKgdTtUzJ5j6pse+atOmMBgxO9w0l60+GpUGdzD34
sIiSL6bzdhpNS5hlnze3n7cGUqa2xnb47xnBv2XqQOKFetNHesodCr4a/pThHO9yjJcHL7OsbwNh
buIcap+xZyqfutwZ4UbeHRuEnTR8/O0u2oTb3NoECucwsv4DxadQ2q2xnAqjN7e1BJoYilEEaO3S
RGlkYiKeA6BbJ9e5zknZuMp6chcnAUp07aq3gEsz+kMOj5NWFCOoM6Bh5RIFTW4g1szf2cC4j+/7
VlGZPOQ6jD1DdBiQ1SHWwwH17CB7giN/Qy64FH3wp8WlvUxwn4SK6/Sg8yQEef3J3nswHViJeRu0
0HSqNzYHPj6MKZw4I3PHTFxlCzMZrPDZuMWkquhXbX+72fpjcTC0U1/5FXABTxoUVZnjVSFYaOxF
sQXf6OBYxVI+Lo10ok664x2KI2wFz6wk997TtGrOHK1hOpwScYM66MjccLaFUG1FnuPZnCKRcqSy
443AyLn4RZOn4lNnOg7zPIRU2ziJxNt76SQqfPMbe00LI3J1tq1Iv969d+T+C98QW6Co4Qrt6v8E
MptWCBf124bM5oQgOKdPPjzVx7gZAipohSGP6hxnaYioTzz3NCHZLCjKf44S2OfxBkA5iH7R7dxL
iPA+7yCaDjplSnMsTOQVhwrbMLsQ4AT6S7/2bhqv+dU3ZWrPMaXClXqH0to7LZJIKjD76ZugFwtc
0GHqaBlGl54V931kAOfj8B1zhVKLtyY8hJe3OlEEWTsltYIZCRcY/VpZRsizKSbnF/YVd7niU7k3
p8YWB4CcBdvmHCYpdSTq4PPYuQn0CtpUKD+pY3tUsVDulunVcXzE+Kg57vC758SHrepmjro5UY1B
Zzy1ho5Rl97KzAV4+vdoJKj5Jtv/iGivwGXfDCOFzdfocgyaeGjNzH/ZO0AB0lIb455N4/qP6o64
hfwScg4me1Fa9tsO0URtDm3oG1T/H/xPqjMaaXmtTdz2HJx5V3n7yrQcoFzgSwFR6LkL7UfraiRk
6PWkLiZpW1SZokg9U+UOrtJeePU4Z3kbDsk//Ym8IU6lFOSXInThVeRVIxtmBJq9fLf2X/Aq5Hg1
WOHYJNSmsGVRRDPSNsGIjOlxvpW+Dl1XXW6vvK0jn0AQ+Q4ZcwYSLGMwPaRm782pOWbETdtmnMqz
97OAGJFSWmphlNOQ6B+iWAnfHxqSDcm6hf5rFfZmh+lKsejkisKMkBFoV0NaP76yLMNQZ0UDZktd
eFGR+i38Cn1lxL5EutIufA87SDPYGnjZeglbtwbw6QlDcoNyM+SFLt1Aw/F2XP0tRm4T1SEb11EN
5HFkZuKreuDkOVyso4lB56OGuPH3J++zW12SxxWwt+a8D6oca3clwbLLHxoLIpofgIyZU2KRqqJh
+hNmNJkIfs8a4eOZ6iBsxuS6Mm2EHQDDShdcYOnjoTMk4uzAytXDYvXpuDO3AnW3hdPDe+UFgU1Y
SucasRJ1N51fgzepA7nDNkh4lc+mDHk7gx7krd2srY0KGHiVvO7vU7TTJxw0dysYruEbGv7L6XoE
+6rauwzyIbEtMw2NUoDDJwPZzHXCdkyJgZaI6oyUImIihZBnchW907Gl2gPs2szYAosG/qqWC7qm
5JPZUVU3JON9/OY6OOOEIYFJDzpX66L+swEgzTpTtYmrpz3RhzuPQC5E1if/wRcaT3Hi/3JzsTAE
jiEETyjeSiwmhb/HwDel7d5x7kA0Syw19XqWeQNzHzIVM96IV3FGarjeAa707eIWhpHX3on+dAd3
iRHcOzThXUpiwKO9DPoDg6kfvhmbmXDvt1yb2X4sUqUyoisvVbQ4Wal5Lz/tlEhe/5PkkIUN816U
QgSqZM6NugPTTOHu/SzkQ+1k1/cBMS+PXq6OQ8lHWHhIXaQe6NOxIhf0tdhNTuOCcv9OSA0pyJpX
oEa2saynX2TqOIAX6eQsG4TjDZ/eDtWZhrT+YBmdD+8MVbSf985fwczykal3U+nN+Xk1fvTyuwIN
uJ09Q76Q+CGO0E55/GG6iXnJr1/QKLgLM2O6BJIPhL+pMHbA+2WEIHAAnE5dplfw8P0vY48MkJBF
7n7neOZpNrcizXoqtb/tN7WwFNKefD8Qg/8oLWZlcQOgfanFVzUAgP6HmhuLq2uoS0yrQmxASK0n
KUpPRTo26F1GDbtOmpmiOP7/IqnNgLbTzpwD+6npziScWDSitRvrIFWa2/sbOumvl01g8b55kgP+
DJjPDWSNPAUQWdSIIXUY98y/yEnfFxUfL4TFRTgokLY65c1OLTOcbU02boMrio8ImVj1009lEPW0
1EvByfXsNJLK1KIYcYR9fUqTr7vnx83bGqDd1h3fUdz6FHX/9PDb+w12Tje7SM2Kpd9HzU+Gi29t
ScDCO62cv5uYywK9AxbfaUpkEM1SEqmVOF/S4P4buGmZ+K2UQ+2YFThhaod3oFSw5WmDci/O6xCS
gUqgsrCzv0uYkoV1eBFrH0DSA72VEZU9Ss0U2ea5WHcYGocQzHQLKr5CJw1e4U+yJU2JA5s9vw/Z
5hlou0zlfwoTAL5bmDwLJd6r4snJewHNiUGz0l7lRCX1oSoDDwfMvl/VhBWBcFr9GuEZ6Sxu0orZ
xhtigAP+rUAtOaOhXcGGgvFn00MMmynmN4lHlr5zdjv52ri1fCI8tKVXBqulG8OIFhhnLEvi7FmD
Gbit73V/Oq+tErpCbI5SSAgqxeHkFHz+oY99csNpgWG425Xk5eaRV+DBsBJrAmlcq3BYUXOm2FRu
51W77jWXe1GdQ9+RpIBWn5o3l3OviE1Hq2Wyp8ASHLFfaOyyiCv9hISqpEYHzrgdA2RTLezO9ZZR
Iybv3L5z1XifcCqF1AWvghM+9A8jphqm0lbbB7M9TL4JNU/oFTUnH0vfQdcj3+T6IYSqfekV4z7/
ymIswgK3Dhri0UKYwJDbOcr7ShsJX2JxkBC3sMQWMTp8TnSQfkRg0kvGDwJy5kUOxNT2aiaLT0f0
lmN+H4phJU7iZePBcPf3Mm+ZHbwSSN6n0le4bOnw5CgYBiB53ZNOHohXb6fcJ9x3600oBRphAGM3
QyUMtgU0+Pukc9R9bF7HssLEOqvnfyA88jgA7603B6XoutLktglzGKVmWtreZ0AehCwD7EJybVIS
gvau0JjLTTipzx8gVSOq2C63jrTH+rYxA/gcs3GTmmgwHQxNjt5XjQlPtBKUurtvb0JsX3dnBzkB
AjEgZoBctQeJrY+3qMf6bRUyXfcU8V784FH8Iv0xM9ttJxwVpHpWH6AwxO3IxVAmI+bhfvf8x2by
YWEXxJ+0Mo3BDTXvGdUgp2zPDDlrzy5OD24ALV7gROHA3pGU+46bgb92lmMgtTmZUj3g+NSlVuiG
uPhl/AO6GqvfCkaTXoHYWg+reUcEMV6kESvLV1qXln0vsSqVhg3tZtDraoFFr8Mw3lj4ehlup9Dq
WXE0jgooltHCrLCecvDNbcxp2abg7MyEttnvbMadYWfUUPgiNxIvkvDT3om32Ao59DyS+unsKDqO
VpMSGIpr3ZFnmdRo/52Ui6zrX04S5a26OooSEzVvixvzUqrwwwFiMyTnSYeLqZb6AcMrwbsah2Ta
fKR8vLNiY2dHkcpbDk/2xUTOTJd8makmtTDSFwTeiN4cpF5xzl/WUUfxAreT2bWOMohTadCVs7yd
5oo8y+cDTEYs7h4+esFaDkepg549kDfHI9/cO1rTBiJYwOd63/4r7m+Tbb98ABJaGsoFwbjI0MM2
osA7rhMRIiwexD/mgXN2h0B2yVD5kWy2wtDAO0cAef2RfAr7kphDOmNWmCLAYortUJO5BxzrfX4W
kNiIpv/McwaS/6Qx3eIJzf85b8fzxvTrEZGmf7hjcOGowQ3j93EX5KkQZmdorogtWWLcNJpCKx16
gM/LX7KMh6JQ7Ffqp8/peXh+juUFU4HBDWw7BB0IqAsCbmhgc4QQEbHxRUwjcBf3OjHpTnMuMmIC
1/XwZVXr0rFk0bnVrZE2+4qNidQSqNehgp2Bwt9tOaZB8XsTDKmpH/j3Z3P7OYC5hhuAtpHZ19kD
g6rAQEx/8PpHMzuR2Ggzq7zXlJ+uTZmueLlxTYS0ouw0Dv7c4q5u9VYJm1HyVBse8gpKVRCblPWw
/dPEf3zCiuGX5iPGn9yEglJw9GfrP4RkEA5bBkLGg1aICLExCfpkeUB+a7c+8zGJ4YjVNDBHvSSy
jCYBfZ/RjSg7a1eVmjPJO7VqU5p4alFmNn5Y3BMNDL+dqVMET7/dNV03p+dspXCkuCVU0EUFqGwP
m0qIoWKgmA9OxXlhDoGC8YjHFziK5kBXIN920HXzkXbvSPLFeoipO72auFVncd61jD9gUBimLiX6
C1wRYiomnPYjh/fpqN1dRQVd0OnfMHb4ieMQFW0Qgmtx00nvjf6qJyI0UOG8pOr7rCriEEWl8s5e
I6PLaLvXuaCw0V0ROutTUToCCLfIjq+2hIJYiC66+zoFqA0CwTILk1gZhHBwRLpYC6nbFbmp/Tjn
HDJ2BpdVLgiSmxyMEVlvw2qhcaY8Dy6sKrjuRRi1H9Lr6LG0zAdRI9PQaFJKj6l6d+T2hqwQkutX
LIQ/NR80G8NwMp4wgSOAGMfCx8+uDIETqBAfXZ/f3nRNlGj0ThWMhAEImBS18R84aqT74rHUqSu1
VAVnZgsUcaoCTTFLNi1HMpTJXgOMUyHcWqSaRaf+yjGqJBDk23e61Pi+1D+30vPo/u4fdH9f+sUG
3yN/LLMm0cKXrYyGINopm6BdA0D33YIlr083E7ECm2300M8O6GVkEAZZMfPOC5j+9VRi6nGTO1UQ
DCW3cNc/ogCyfrejzhPL5nuab0knYx61fkiolaBlVfgKKyv6W+RHU3WiIjgFMwIS98/uYSatgrbN
hTOJOzko7QftiX5wHYOBuTaM7oh8hPWRbO+2WFm+kEUN/Lcnj9Ia476LKQBbSjJPssSW0Adqse8O
st1/r0M9gVNCShQ/oNlXlyEuj9fc9V5nFPF2Exm9YiOoiNPRcGeXiXjOxtsUBd2FDISuZimYsKHB
HKldiFq6/8BuLQ/zUe4ax8rZ0/A5LprDX7ZiPuStrzx4zuHF347lYhZz6djPhx1eHyaiE4jxuPhS
Tqly7L8HaHFM//XxBUIvz+wbRhiOhYw1kgsoua0wAReOXmphYGf5alk3Y3A7T/SMy2/Y1D75qKHE
mzIM5hMXEjoOTM1r2XLfyvtYu//4Q9sChHycmuD8arTIPvWwn2gZAr+pFTc4HMPu7WPxJaE+uMfZ
s1Pklr9y+Mm00GvwVVbpvwg/cpq3Fxqzl9JK+zp4WmN3xxLsNhTxMEi5IDz3okXXugqZ+oATIaRq
RMge2BGulooZJStN3Hmuz4Ar9oy40Q6vk97JVAJmOQUiD0uV94I2Qt+D47gTrVQhXiETwjFZA1vZ
HW8PXDkbcBoZc+AO32fQy2tLYzwQXYcbodnbMLB+FmIuZBJaF4HA8AOLmR4YA52A5ARScK/JmrOo
hC56hFzd2rSdULWc4eAaXWH7T1k7VfYyZBpkzERnh5KhBTfYMrtxj/48LREFRPlCL1xScFDFtZSZ
sYkXuiq5Ec5ErEBl+snqLHqDFLFqLOIE8LJcpiJoSO+8RX5L6H17FrfY4V39z8gMKBCdizCHYWwm
qQxRGS1OE6nyVSgyPoTQvYRFSS5fWCftQ+9YyXfm1J1vHa7w5v+fFojdIvyYtk8gaEabxcQ85Ump
cge9ht5tjlLH0mYnxwLr/PUqg0ef875C7+3rXhtpP6ikkZUDMkZh8F3kFOGPsHST4kMkvV2YqWkY
huxqTQv5Ri/18CubfQq3KGlsnIQlWgwqUsV3LKHGjHCoSWDovFUuJPii3QAl0e0cWs+CsIBDb1+e
qgr1Q9mgk+R6cnzx2RiWET3ett3OGTxiFY4LYbYdQeJBQ0Ga+tULYae8GLyjsvEFvEr1MXQxyxop
ZHdntMMV5/Fy3UzNr8TES01E7hmTXEcEUt2f2Bv3xlsfxoI+XK4p+3IoKG+bJURY1GZ9BcidsShx
4qC5o5pLcx4zMK354bdl26cmMwducyQY55L2rUX6u9FebBhSmos4bP7uvQMtvzvNtGATP2YHU84O
UbVc4UK1ejlMteeDH5UHOejATG2GSG6IXqD4SiEMZrjIXr5jLQXgZW79p7byT6tlS10f7WOXdlZ5
TyNbE8BFo+gWMhZzNbU/TIQrZQx41eRGx59I4T08NaavDDHnrNdsVx9i2e/XRs4kzhSO1sxikJFd
rmeDZKv49dIKHQPFcs2ZXC9BOzyvzsp/q3qCSGX9zNzDCGKnRO36GMrqrtfgU9c7ubPqatT6xP1F
Z9vypCSBZOdhnrcsQMqGBmYZmnRrF/+N/Aq07SeVCI6qXaxYYILY7JtSIdBKN+Hj1bMCrBhL8gdB
I4ClRxOigMYuQXguq3A5A8S1CFXeuI9Fd46jTcuzaodz9t0pE08V9ZQktrmMg5ug6MtlDfWyPk+L
Wl50NQmYA+o2J/Ir0OI5kx5tfybP7ZNqeC0RTfv7xFdGl15aAId8WFp0o04kcMN8I2JQy8zhiyuC
yx2zsqN8S3jfrFogWWJOce9xY3dyt6nsV5kMaAzUNWOiJFjNmSxSixnms2iDwNrfKP0kmz3wDJJL
DXy3kvXu4aTOeWzi/cBGVQITW7iOnFzso9rC3JjDc0ariw0R3ROOcQmzsruXjShkwYVItuyp3+lE
JNIfHZI6O0p6Kqs9vAPmRjO6iKFBiWv4+SKQXrQPjLifngcRqj0rljtrLcIjm8tTEFNL0Jxq9txa
CwdJHKPa5yAPlW4G61OksuPLFK2UmMutN94ovsZKijRagc2BDoNh8tPpShMxgLCUlKLJA8TUdK58
TfXuUT0s0FOTuu+4bX72MY4Jgm0tDfqc3qz/034ZzqHQiouDrmBmyzbex8Ivrlha2My/ACN4vKzh
u42kNTm4LlKyWlbvbmMO3EzK/BoTupXug10n6K9ZXO6Bp+6DmNk2mECQ6+HP8FpTGPkYieJ9gp9s
B/v8bo2AK7C3xnDb/WNOAyyeS4pUfKf8uFhT62mcOBN48aVnNM2Qx4KE1LOb0v55sct3TJVzYOLt
SzBq1ENaBc9nmfY6cZD/u6VuGGq2Y5UGu5Fy2oWOztuCIJdND89j6IdvFqGsWyObMwRzswzuN3wx
6oQIKq1JaagBEvSRGFyE932HgPZ7iDqAIwpRBBd+ExB6Lty4UnBGLbPscHpybe/+deiWCdw93uFZ
mQ/cIpcr6AkAy87Wn61OdjaUYub69P+hPEc8cEl23Dpr3pRPmENq+L3BWNQtznmyKaaNIlbwB0Tb
gh8JzuOkHyvQB7MfyJtz5ST0M+32bq/4uBrOMM1cEy0QsMYxzH6g/pGlrAv1Z5U6vIVVUlZ+rXnu
QA/N5CtBOk5fF2bn6dQoULR0ydcYgF99vBH+oNmy/S67ntp2jz8xiR/Cn9Rhtkv5/09RnQV/pubc
u1x8YomxwdlP8lK34RazL1EDJtj1G9y0lUArrFPEtXj+ZI0H1IkzcDMZrQWe7VGuECOTYJXuJBbd
N+pvSuBkEXVFc69OAGGZ5TmgGvl37Ggvo5U8etKx1ieBPs+GXsViFy6hFlHT9WTkYVC8BqnddUoS
CmtRB2ZraZJCCXoyJ2vpY9as8wjVo+v28X2SJ+p8fdBy8hx/ogahIW2K2x2WAn0UBgo6O2Hxlxrn
unznG/x7qfZT6yK+fs3BM9VVsOZvHlEkTc06GnfjMLSRoqG5KijsqCpqI7Hk74nZVjFxVFJJaBhl
wjikfvU9CmEDn3Aam5cs2LJHptbq5IV9IqquXxm+qVThnNwsK1imVCMcEFqeonivdKlsVXIXqHB7
dyRuBlx1lTEiploOdfkflAdVtInE0TVKfH0Fwxw3M/ViEA8hp1WjQX2wMHslxYBMsTUjW+Re3KgA
sqgxd6V9X1cQ0iXxcCTnYMa/XgydmwjeV3wS5pXIvqjAlFj4oAHrpq0NWLPuLt74QwUzvXsshTA5
a/Ul04QJdwzwEmsVVrCQKLZnG6XbdPInb39kcF2cgHbg34xDA3SOJvaR1P/yMFpK02alWt15Z/SG
XjVVzSV7TNOqAc5LaFKtXXnWloB7t2SeK+rsjjqSC+Z6JaDzMZw2U3npbw+o90Ushw9YlgRWO+Kl
6Wv6HulQUVFn5ylKaECb2SiRjLWAmn7lWHgC9zYOxMYnHeDLcEguwUSF5neU76HUMlT7opQTZITv
fGOQvNYk5VSX48JWyGx2stcZczSoouhsII8UH1Hk59RFY8E2g1F3wCiGdDPo+sSJFxipHaJOh5PS
Am74UZbKedb+PMCM+JA+Bnfq+cZkxFYg0mG1PDDVdYY7uZvEwUUDmU7hg12XsdQlP5a6gchUtSfh
jwF8d2DJQGt//ImSWD3g8RN5ZeweqPMHDHlRAwX6N3HA0BmADi5Z7VZ+5gnrVBaefCAZ65gEH9VX
y9eglm6FksbCJhpB1CL0mY4VN7VftZLJqSO1CWjLJZkQ1YAYeFpYnts1yUh0nLGPht19S2CovwcA
O5XrEEYKPTqZaY61Lech4IR7rxNWfIISQg7oG0d6Scon4S51TsHYd9XgC1Majczfrk/huGTcUxi7
aA7l21rRWd84ftduCoKm3CotXq6YsJYpyL3TuZoWktCnFtA19J72Pfjv6UoQfEsVxGVwozJCyz1y
Z5Orh0PyRToEU/FCVeaRci4akHY91JtSDnsnJcV0JNpn6GelkOEzw7QkEXxg8LBD5dYIjjkvzKUP
O2cr2+6LQOkI2F1cgz623BzcVgPjTsCyeVBHWKIgE3qUwpsFoDTxkC+30P6P0mxkM952kCSjdqfb
86qQ3MFIqep2MtcaFg0vDc9Eswm1iZs9jYUmSbBmBYG4X2qD/mtQZUjFYgHrSUQht/s147Owdah3
PMNI9FsjCL5FVOfNuoO7blRIV/vlcV1Y9Cp2UJyxKwZ1rUa4t42VkD8AQAZXapowJLxtzxTMRdcW
Oc5Jwiv6eD6v+rL8dbUtt8RMkYnVVLolm35ykruZHEwOAWBbxvhuMOIGGFSEiVcj7Xd7S/Gr/z4R
5iskKGYLHm39hr15u6mm4pFvdw4uIkTWVYbsKjbu3o0HggGfE1p0WufIfUkK3RHP6kB9eB9gCkYH
V+GB05w0V/y6UhXPYan1sKYdPV5hsdY9ElNvb4h5SPZ7pJyVY7glKNcOQMNjjtVptaBPQobbrA0K
OIWO2cF1FEZ+PXLDoTx4FTTuT8W1c/Idzjq5Tn24AFhGRDhggu6x8N3ZvJNdebeNocT/2eye9HM0
plTQpAksjkfxmUqlWdoGAxcBri1bPxcB+0NC4Z2Vljxj8xJcK+7ULN+CfO4kZzivK13Vyot5kv+X
/ia/yoz9yXwA5/TQu2bUPwpBJ1Jhd4KsGB3KXk0E645TKvpQiOmZJecA7aHlxUzPviulpGiAd0Ie
8C+Hkur+knHlxqfHomgC6uzDttt3rGoVSZJgdZfhTjbNhTpnksEX9H4xZwECZQ4l3SalTM0sPKzB
eoOnjwDahlRCrABsUis+IydBORqNQkMIY1aSoAEq7jVultjYcHpccBDnTvVgmmxwehebLj2Ygf/y
IMcxWtmQ9Sfbf7/nJ1CHs6pGxjcYQBsMpLaLX+cL+OBiOlasOoyOfImlk83ZhebCAKRz3MNGqu6o
+y2NIWmqhLEMI5yi7hczvJs/zDBm5JKXLuBebq1ByY/cPekxeAkP/ZLk2L0aW3qxGN2ircmjqjwr
m0zb96mdr8alOlSn45lzQe3TLQf9BWAy7/AVyzHXVopYQdnuBKBlwg94emnxKnTTyT3iWlG1nkmk
Ud7wtGjMPLJKzjL5EquSBA3BE0JldyRZynbjoHGAu9OD44oo013iLWGhqG0Jf9lnQ7lpU7hEqX/H
G8JtyfWq4Z85WyFfMUntq+GKrNTHDHfQR5UpcNjwM6x7Tge3O15Ns0CSctCtGy+S2527NEl4pT2M
s1s6WuYttlwxQ0uuSckxD8O/KSsDwZbBmiH8eBjIx3G2vYSKAxcHH3rq/dwnb9Nq2ezI3TVIME4h
tjYySWPT0AexR7gnYhM5qyZwrKvltqx5C+Xk+Cdepe8pjRMS6VWXVWYD/gWSBkU3kInPJBSnHNlv
YVfecnAAh7ypCBgcofOV9h/fR7z2aTv9mrtjaBVpSplXy+t3wrfHM4MVh4bnC1QBcfvgNaXgC7rh
zan3RIK6/DqZX+ajLY6r4NYswIHeqyvZa9b6ZExZJm6Xwd/X6iYXxsQ9OM+sUMYTOuk8WHREqbeg
eT+spNvZySuRicKRde7dVZXWhA8FQIe0b6RyhRqhHAdYOy6GFjuAdn8mfKA833YU4NMS7jKRDGEe
hzkcHkIzA2Uns4V9KasaFO7rL4OOEcsnX8l2TtgyXLvqVf4E86+ccz6p+RsT7qi28hjEwVqRykgn
tpeewiQiONvbCip55AT9c5P1sg/c71n1xI6XpIpaloa1M+nPT0dPdhPdiT00BmdRjVYwm5o9M+cx
Ms4ShVpY7+prrtzeb4+cD42spgcx2Ft0GaoQAMV/dG90VuVYvGVh/j2tGlHMe/ERNFGLWtJMZkbj
LPULaW12YFyQtnB2OxLFbECnHf1W6lHzUj9myzOWGMc3063pWfzvw+I2Rz9Rd2x2T1LLIY7r8PHq
U1FIc546/oN0W+AsPwC0muhDZiHrYco2fa/1ogsIc9QUhFAakmRp1DRIQf7lqBmPNBaTlDeSQa00
oibeaV0S0kdnvxl945AteeKBv8o9NZsFKRl8+U7Rq+VpIaYe8T6t7j3Yr32GeP2E1wOmSQR8IoCq
uViBYA/l6SvF/XqvYkTuZ59mnZdcuhHSyUlmtyGrp0KGYQArZN9wblYtto/EzzYtjlm2yHOGyrM0
EO50cX+yuOOFCEisbIOdvKBRXn8lLN0waJ3qYfKXE4POWOfo8KFZIF4GYp7ZinnDNa3aDRQQ8YLU
n6JQEQVByUlQmYIkCF56hOviStVu/Yt34nqjNvg3SghczZ1jg5XPwNT/zSeG3JuBYFzrLdkX6NBP
o//qmzEPyKwo7jxPLZcyYYZLae4OQi2GkAKcDQISZzNf8guxz5CSIAIAhevTdFcQa3UgX1QNuX0O
tOiQGsmwNfW2Ax2ethNMHmCie0vpRq33j4HcLizt/NQrKa1OOrbglMC2AQ2p3uem48RdoUEdJ6UD
UUQHRQ7PAjydZ8zE8S5Y3JY3cyqP39svM5tk90L9JCvgH2giUbKbEDzcFlctTJbRtuVeDvXl3z1U
acSLHk1PiOjggNbu76n47z8dfieqm/9xnPcD4oY4R1HGkdYA7MZlvg0W1BJhlwcoWhTRq+6wQjP1
BMl56OzqHIeBUkuGwKbRSL0frGcGDBk9NyjGb6pVgMkvpRX9UB0jXs/WbzeQf3fu9jaPVe+nRJdY
Ci7Fk+4hbqhpSWTjoB0DAAUvKIQJpzshqKVwUuBvbev2ymkqKZkrCbahyGULn9QCjse0YNWgAJyo
E5z1rJfmLuG6Su7tlQwoQG5RD8VmsSNu1gMOpjDW0fGEGrZLQv670GZvAcPfRPiGJ2359+V95KgY
Yc99E6ENR7ll9z0D1j848kV+n/GfArzsbmyiTXPuHOqFbYhlcIF6I6xEl2i78U+240tvpYxtV+XU
7kHJH/9+FtVu+QPgJEWsc1pIhDjNY7ICOwVtZ3Hq4YJlO3J/hhOPbbF9Fp4ouZQH5Z3I0518s/80
hRm6tUghsjQqpdsvvgGuUZGxyNPBSMEF6Lp4J7Tu67E2ZlhNPzo1PLSktHXybVMsLZ/VVSG7xwFb
WGwfAsFp+RYcx0fKI0rOyL80fgew0rXxp+/LvonTyn1NNAdl9aTBY4Ohue+Vlp6jkzZYMg7cav2H
u7431hapxMDzZ9Zqm60f/NOvf6EH1B9QnghIn3xJeX6TLEE81XAY7hEdWgFOmd8fT6EW9Q9KsIuu
fsOydmnO1P0w4l0/RhQr2hMc9O78/okwfnGZ03kenV3EYP0x7Az9OWq15WCUxCigqp4Dw7PzhMCR
YCctkoPKZsJlcPa2TUhefTTkwRCtC7/bhTEhBhEXqv/QRwVAHXRmQ4A533WzzSMW1aElIk3kNV05
esfdlB2SO6dmsxjfP7hFTU5T+B3oimp2/QFbA4t2APjVVcwAmAEwVlIYkRSsQ9GxjTdnZXqnk9As
+371XC6v3NzXKop7uOMd4w5meXi+7kvHr/TuJP0KlatFqYFuhdwvh49L9BiFUwIivX2Xgg/6xTPF
njy/rFMNxvoZReju3MaSq7fY1PhRM0ZerRI64498iQEA/1BLeNngeDn2i2zJ0feOkR5micbyhBV/
LrxXro0O6UmlyJ2f7tGKU8SJpW/S1f0Dt47nn1QX5wTKcp5Ywm1rbURTfolL0BsdAp4vu//11+Ls
dW7k3FjmrYLfyODQe2TSwlJHaDVBdGMWC3i/wYg+hKD4Bv7/6AiUaFYVvxBV+/bz/XzclwGOxrXL
RZFfms7WPAt945J5/sir+HcbfgiMaDuB8ZH2LUG9xUNa0qwjoepNiCoPb0cd+uqhfoO5IrMGk6aU
wFA+RaBlDHgq3p7p7CdNePUuk1buyuXAzUd06XwLRZimuZ3cEpw24RSzPsbn7nNC+NqqY4F+nj0p
s0C/aKatFIFuGLLe+HKDJZL1yxrUFo84iXDghmJkBrV3VVb8FPBdSmCnJCyWrX6JuIpqTIOBSRvI
p70IhK0jiRqqr2VDurKMQWePjjUCe5FBULVKHehW051ucXD2hth+dQaoR80Ixp1UYQRcXgHE3mjU
TEEzQ8t7lb0/4mhP4hdNiRQEyj6tlLnEM0l5PWhULrxlnMfotG3oDxEGYeblMvEzO/pjAP9ODEAD
0dX+ZpscTboYQTFD2tEqqxBvv8A5fdAnHEVCVnMMnvR9sPJ+wy2Ky5vG3cJgALfWLHzsIdGzAU79
l9KIkr/tKRvOCNw2cZZ2ARmwBak4d+Tbg2TAlsX5YqMvrHmYLZwy2hX8pgKM5DomOiMfWz744AVO
gjUX1dS9mjAYKr4lyScQO0zVUwDBdoKuGR5WnYyByAXr88KXoSIOtXpLpEvLipzTkYznNcsysDwu
SzUcbn+HfR5gSgZK5kYdTtaUSo+zktlsJDk6iugFfFU/h04hyebLfF/bBVH8SrDbK6R0qTfEPxcG
Tp9tcws5BoWUrajWKISjxOeAqmUgZCs5wSWC7QrI4VGod8mE63QgqL3LQip0+QLhPV4qFG054/Da
ueyRYW/CnOw63OUTHx/r85ram4Bkr54AFj8i6sD9QgJSKwzvq4aOQSFa2mGSWIn0+DyO34j3YgoB
K7xX0UQ1f/hox2aYzTVUxeiumxVYqw/eLY3A2CKZ0hkS4VBGwii8VVjM9zA9qwKISKjp26VkmMS7
CQac+dkrr9JpPtYApojiIxNYWUGjRgerN3/rlUoeoRtpbOu6hCaOuCXj/StBxzoV+YM3Kb1JjQ0c
R94zhOh2LqNoPzkx72U1ONF8cVXTtQ6nEQVZl3+rgQmHgMqOabBAqFis+FrThwTqhGUiZEtbG3ng
E70FTS6Cqec8dkUX9crDjbCoay7dHX8C2KOUqXn55w3CGIfzi9cYt8G/yRDJIXDLXdbyHYg2WXCk
fxlEIa37WmSTsQL4KTvJlrQ5FOF6Sghi3F6fwolqK9qdzs70ap0tAxzzWK4TZa0du4+jn3rAHriR
20fYCWUPRGpO1oOJoU66Z6btVdq913DtvxU0rDe0puZk59y0YxvbIzjX4/hXSp68mCC8rl+UsQdf
arxGD2+XGUiPuG1UvzFIhdr712VXcsu2zrBLr7fYM2PXYbDgoZhDPJj2xKLb3I1i6ZiPoRwcwVjA
0c13TpVtPq+X6qru15q4RUoRBGx40vxuYOj09+NLhUm29mEfcSu65TddOrzD/OJIx8hDNNfZQB8A
HtKLSW1lVfZWVDRONGqkMwMvgeCLfvbFQ4tv8XTogrQ9XID1zw31VC3xAR1/wDsoVTC5QZQWV1+5
3g5y8PVa5xqpMIsFufu4wHKlaT1tZ+XfTXDOFlJ3xn92jb2UD5PRM/vEHBfR1943TBH02ujJIxWD
iLBPT0LxfhoIj1tLjH9vvlY0SX1lDi1sST0bWpcoxMY7F8DWpgDsyD1szVQa1aLQ4zAYMc0fDcq9
srhzwx5vkBPDFrQ3brpJ8zvcGG9VRFRC73foyABnw1DVMZ5qCKmBtsUX7/OQIryfhmBedd2BbeyR
gC30lR5s/pDweQKIfUD+7k/HMOJXKowEpgs1jKXNGV6K77cZyxenAKjRzOyKHXqT/KFoomRo96VT
W4litQ51D5cep9W0nl7YfnNCY7c0ByQKXuvY3tVKRh3+F6FgbZhuYvXG5jSPL/EYBtVhZKSXPgLS
55VfDmkfBwQfEDqoXKmN0MHl3XIXYYrTeFcDZlTxJtWecH0SK5/o2TGmOnvPMFkArhcANhG4jYGy
jhXCoP2jtIJr3k7wRrwBhzhdHTWJOanucdweI9xcXqkKa5W848AqvHeraVNHJqHFWYapDhvtywcG
14WJDstrX50eZTUyGEj2yRDh1QjRDyGWpywEhd095EtfAqUZYdX72FjbgCdqa3iAUci4Z26Djf4U
1tnPkbXSLBA8CG0hhOfk1ycenkagCaW+6bjmiBZPlN2sSRH2eiG9xywLsx91o+IpDzKU296dp8Ty
6JJtDxsJIePOWjcoeGmwEQW2kDS6XwB7+omg02TKj34974FYo/I+EyB6x78GogcbiesUH/JrEgSQ
tBoIS0X+Jc0W7beMTdx+7efJPnxPPBhZMyqLyHlLbrIxI96KAodlJ6+ouYF5KatOBZQuZApkxF4s
pAoos2h7ajDBIBZYejlcGWOCbILEhvck/1kBn+cNHJW2Bp2ylaE1a4VKq1RvvuyGJeWNE1OUJfzx
G374qmMFtftlYzVuKApNVzVIDXwto7/+VHZU5RqZjCS8rIOfFv+vonE3+3ZsSTIXoXDd/yxKdowi
8kVnw17oTjVs/696YWJm7rWjtgNFC/RXaGFvl3vhW3308v2c10JZWgYTFuWqjvS3kO8pyytS+Xfk
PEuzfBg8WT+Y1Rs3JljHdJMYcbmE50RmE2+Y/u0/d1VN5s0hjA4PQ2ztLknn8iJAkw6nc0DkFcSu
FldoaZDE6sppoHkoSS/DxDhc63m67InobDN105G8zo09npvSB3vPoahZt0p0o2WkSopgLdyr7+f1
guAI4FtN3IJrv7W2TCIbzWUHgVL/MbWp1mmTCIwb4ICXqsakCdNjBXV5DTNbkF4pmEpRUG2NGunA
VXMbvoemipoqVxcs5IKmMiNi4rLEAsk5+yUp/CWI3IaU2f9nngMBoLF8JeH3TLoqWKNEvZ5ZC+41
U9X/L7Z0w061r8jLWmLRuVIbyTKGPEzgIgC/od3CM6GqR1q9YNwOGvKOXVQA6LzXihlGJb+e9cF1
eoNauMQ2icUMJRv9+flxJf7zIzdgTsrpB82xxulPkCa/eOg5koVzdt6E/iJuDa41gzco/ulqBWiZ
hpQjPtzDHMkcvS/jAApMMNROOhyqajuBcr3wQZKO3d/e4y09va/j5K4JlxmLY4IfbzdgG4RjPjJm
OP5aK4hkYQ/5kuxtUfokVDF0080J5E3wF0TgUKY1hmoCIKKG2Pif3IoR8zaJsbuVhKSgt/tNJ74v
V925zOVYduxUbc9FR1fdE5gTzBiklE7RSFe2OQofoXG9bNnz6kdNEIyV8wpD4BxxUMecsSQVsp0n
Wg1Fw0Uri47Erjozh2kq7aV7kvPjWOZF0jHIPWxRpeStATc5+1DvQ9j6bDX6+zpmY+W3mQPO+KvW
T+/T6awWzqUAiXBrXPWwaIXCN3hdgpc6R/cTCaXzyadQeMRdPe7LAwN27dml/qp91MM6GwSL7YRJ
T7XIOPYSaBt45k1VALEWThlvkCBvOsuajVCHyka/pktkAesOs4b6vAVSp97mGIafgV6W7GODi3nA
q3rW/qu72Z08cuBs2clkiQf+Q45t3dL+536gJnZn5u7ygVsko0t8SJWEwKshA5i7ASdn1TjqXu2W
3Effi6YqhnJqayEYVxoHo/VjDb9q60n0oy6oirWHM//V50KTHLP/tft0vWT4NIIJ3NQwyc9kWEzH
JDYOtTuNWCBfB4SIcck+cN1qYSnkVS4PClFtTmcr+qy9kpBDq/4dguWMMUPt/ue1e+gxyQQ1b46s
TAtVuf+3DzH7+M62jhCn4CfhwPC1a4XWrR6hjp0Cnq+yy/fjkPRfFkYOWw+Zc1ZfgF0smlxzRK1Q
Fy+0hFGG80jkgek72JBkWqRuFKppGTIGC13FtOTTsV+hN9k5zA/EnqwCuDRnlHjljMOQ34VyQWpT
tEz0qXBpOMR/cEBeV+jH7QSjDDcTlj5vXplj3qWP8iNZLIIrphvJdf1feuWlna9ojVa/vs7VfFCL
Wv3/fPpxldniVvj76D2/L3Rmgtm7xslLVrReFEKFyChiB0WUK28H8ijzXrZGQdyNMiYZQe0ODTX7
z5APr8fP3eEIzVGSpXAp1QruyLBqPra2WeK1JH7L74yf4utmhZbGzKegp/cBQqYb+sPEW66U0RQl
t5wfB2haZLGV3b3LvLX+8dD6FoEaaEmdSAS72QCeVsV/HD0PE3zMlzlxvSe3EIfiL0ZnPun8nO37
I53eK6AQJaq36YUszY8zvVmuqeM4W6csr9jJYAiJ/3N51oT1YHbVbgzDw3Uhb57jldZYGJYPLim9
lMhu4m+EATaUnixToKgVhv4gRHy4a1KP5GuYYnU2+jO9ePHj6FpP3Lh/0FiEN8bCa0oxkNN5oPP5
j4QZgrP2iCj8MSqltb4y6EJer7bkOEHXegJPpxn5V02Ne5et2jGZGqJMfFU9Qt84kPr1DNP845z1
caUSAjGbbDnni+EyXkwsDyHuqdOkKDedgiN3Qe/f96NuEtpbYrXSyyuzdpvY/HSnJJmAjeHaiLGG
kE+vBpqj4fQT1ffGtjd9n7rG4KR4DgeVLfiiAA1JJzDK7bzsVUaxDz7OqUrEwKVdYVTTBVfCs8i6
hWujgjh3KzvfD9Sj6WioOskPfMrOucH3chO/RKqSNF66oOUlbv8vOMsYT1E1GejIyQ9Jigy5nbmP
Gdj6U4hUJKfrn9ekCgyCPXZx3AEhzJy9FyLInvLYw4awIVEiDoj3LjahuI5Yb2CyzNZpVpPG3f+C
PKDvDl17hkQN6UzBAqKpyTpqe7OF7inoigZj32vpMU/wqej7Synm/PrUWCq7E4eHE4uM8ypDtgQg
trhOEMxxsK2nkqdQGJCva8TqEyjLRIEBnNGVso+TRqYAgCX712SmISIImKHtWo3OL54sMFkfzG1k
HcB6YsAavqD7hR4t6zaA+K6pk9r8xI1SuIPghgsftl5m1pptZFiKXd8tnWH7Af2Y7BtdNZ8YwBmY
lQBmFJW+kYhr3ul2bG5y1LLabn3KlWYFahrpm2xvMnV7S/b6nRQVHnMur1hjMhSgAxys+sn28fOU
44kBiHyYIWWAjmA5FFabTuU2Lj+a7RzrsFIkvOfOMLYyF/+8SySA3C81qGzUOxnEdo4LnS5op78D
7c4Errn7FYA4T7W11F3IEcV/d+yUVtjnFeO3Fekpxcb+D40xJOAfRLRkNer161QHLGMxlPiKkIeD
q1jYmYPKvzExizBbF3WY0P7r7vUJhN9zA4+7iOmbvGhBzs91JGbz30rKUBchggR6Bq5Fnzv73P+F
WBr3J9QXA1nlGYqUY/VHuel8IRmJ3LExYGYo6M+zFF4OJMEVR1tyU716ZXVKrE3EhBvDkTs9X8Z2
BeXyAsCihheYK4Xihs+nv0Y+2qUWbPSHb7+om7ukEjELWQWhZctOV3Fm6nVv7UM8qQ6u7AQR3iLt
pjw7OrGpKiETsJ5XVSaFgU8FQO+G1v5ZjA+tRutStAtsSxF4P47z+Eyi82LJ/O6h2uOmtKb4Kh2I
Cq0fXa/MVn379Z60r7y5CHzVqshN0o+QhFGn0Y51RsvfuQg3evJaaoiT9cdmINX4rYanYg5qHtev
vvj3OGxoZvHR9hIqZroQPynwAHrr2buOCvVpk37N2UoQ051FoI37KHTT7f8zhVt/DeVAZWbVoNBA
GsdDMQCRd40zDxpNXEgvwr8ylpwfuUh9hMrwD5SJ/SB2qQySJMVqN+CyiKKpMd7ZBFAelpGEUIuz
LRk1bvjfJvTAItxOVdRwiW6TPFNB7NlEwwsyN5zXlwMVj77EbC/DX34TF/yAr3PEmRS/1FNKQ2/m
U5wf+2vT8KMt+PMeZ5lF5loCzxJ5Q6kpYC3SQi7qg32VxWZHzO3UqBe2Y7q6wKSP4/3bcY9ksevs
oov9kN8z7zgFTccDPLcn8EVP8qbiK/FuLhM2HqZ/R87aSSVdyObL0sKdLUSfADvHBQy2uKooCai6
9/yjzeKyplogXNjc4v+qYv5mceB5uG54sNyLuZxJe/D0SCk1EgsCyxgfoUEB/udhLHmbrEDMvkOc
ucPabqVADiD7sRil9j2i9NaDqB3lVgWIxzgzmlgf/6gaqJ+BOm72wRLPGIu4S/rZGUR4XEy2dNZ1
hQadjPjwc30B5CXZBq5LHOQofiAuk4au8zwgpKP47+FoBTTyKdfVfQLfNrj3+e0toxAQTDUyDFQ/
8ebvjLivtWURLUqiNDPc4vBn7/EEJy3KDHvxt81H4YH1mz9R/Br3hmyZL+cixC9s+X0o5CMMAtaN
rbWDSTANkcPgw3VnEWHwMLOGmxAGKmReWJPutOlZNV0aVgqwzePz9ntli6gpzxjiwQ9+vGBAg0hE
dy1Vnm1mcXDfojvg+BpbRrGvDBOi6lOuOHSbe9x1harP0atjHd4ZCC/uHpSlQAZ1I9LxJAISPHLh
e8XYzAaxzC8pzpYUvSpJeymVCGMMB8XhxLKzBJ5M5rDCg4V6hy9XI3XqBLMSmKI4OcCbdCnNQCiz
ComCjQPc8BGkWiWN6IYkGyYdfO1cq2k6KFAOnYxN32uYDNoZi9calh9WXNXgx3tOp+6HX2etuTmM
FBZNR2wRtUlRD5QBtnZMoeqNdnawhk7Hn8b7XjobAXB2Ez6syJmaeErnwLEbYPFx6VrUAlOT+SLM
KGoO4t1sG4BcNwpLpJvzFfUmJFyOWcU4t/gb/xWUuaoEYhZdaaOCEaDYe7WMagBpHtaSDWw3ujeo
lgvjxLwhxOBJak/n9CjA/sNNeoWjk4wcGrvDhWrkmm5IXYrglAZE1Cc1ziq/+3ggzNv31op7DAXN
P1Uc5l1X8MVlgAo4I0zFiqVdDILJSL40S3KpK/vCk+qYcYqloqGf1t6/hvtzd4hOyONzwnm35bvQ
v1MByDHTEJwVClPo+R99VMxrDdlu7SA56eiLkMm6jsk0hBRentxuSxvLatlmoWyO8AXEJHiHOIIP
c1p7q25el5jzTBt5/23BrA9gwV+egr+z/irfDLVpjxTBA18Kbxc5b0SBSvUZ8YsUiuAlYiMM6+M5
ZUh73KvUd97npV+XYOcGPGJhwXYUVEAtnVRRS1cioSlzjbR9XJTxxHm3++NuzplHi333bLDYMD6U
bLR5702VtBspNMAqn2SkRZmphOfdCtQpZvCSQv5AXSXSmfS59skcMU84yIe9ywhkD8ODp2cruCTs
ctAqHkMZZw4mbDEz2YvFg7RCQs+89dw3cMhKcFVF7jYlmsnv1HXobuK/1hms4QfZ+fVSDw0p9lRW
8Iq+7Wb3QcxnpKPc02NOp7CwyCfU53ehTEYm5x9YiXt7eMox5PxQHJPV7Yn2By9nrxVtz89K0rvS
So4DQuR+oJJw9nhkK8lm2X88vJgY1zRzAHv+PXXK4vM8jIdCRQ9dCRJV41GMoOKooNcymUXwmzM2
+z1D67HmFdPamoIVsFg6+PO08xGWuLAWTGSgB9YmzWalgO5Juqna0jEUaLL96120XJJTstm5ylTL
HhK2Bturmp58E8PBRSMWDEhM+5ff91z7klMa0QgpFQqyCPG4yob1L/k5xqCLAyIyFC7tbtlIliO5
X6sn/MzOvQl6GJ3F3TUJ4TQD2yAZgEw65WvIiSJQvMNTR/GN9iJjXGltrGq+mMOOEjC8c2ex0P2x
9fv46048QK9/gY3U78L6iuY95mWOxBWZ1hA17BnRrKQuD3im57Obuw269WNOrzrGJX6ApKKdAcOR
TZr5wmudr3/ZQon7BhnVzbIdrkJe8Nx0RJfLujcM4vLl2PSR8+ErzDH2aX8/dsEGs8d9ec34ym+b
LcxfDLCCud4RH0j2p+kdUBdc4zBJO8AKzal4JOxYUZz1GZYxKwZ4vxyHhxD0Z/1wz0NrUTItLM4v
BOcjdqVP9I5EFDxG370Af20Zlu9d8foOIztJ1X7WRv1qrYocMMhWRhfcj5+KlD3NnBl8HkGiuq1r
4YDRLD/zDbWRqa8FhHQFGiRqcN+HI6RbPLx3SrJ7pj0Zq8uI1e4k76Hr9FxezT6dub/Yv0hPXdAz
KEtZfF+F70ysYejxQq+OFNFoqKXw8IckWLjVvEppLia6saJlmttI69ujL7nHE6wXgPYUzDR+/K8B
vgB5S9GS/Rxpa+tSVl5UumShuHlDCvJ1HhLuuLYtFSZzQ8voAzecqLZPw1ZrvELLPOdEfYMJFXmm
SahzRY40jkOzaFi7YoPtHOqnVi/fKWCde8Hy85vXLje/ikWsqJxl6qlzC9/5uY6J2J0hlsN+QPef
BITbs5iduhz6eFu1pIqavvw/arKy2lc0MDLUllNWeKP3/LzAjumnilj2+WvaJ3LPdSt/78ndW5Mh
jTtCsExBJP8jJk+tQ65lPwomDl4zifX1kLOJRcsbj0xxEXOGkVejLlWKWfOVApFX2YCBl4XIb2Rk
Euy7ZKfw8WLjsWnUcrdPpT6n0P4JBo4NoXQgbv8DeqgCVKLexGqXHfAUo3Pbs/WLR51/1IRukGGf
ZdxW/c4HWEYTqke1kUUY0ceo0RgrFqZJUeQSTauFKj17S5shUMSEg+h6VMM72PFAkMzpd6HiSEJS
9KyWKhiadZlsUKjo/1ksBY/q20xEck7E5MUfra/AzrX5Oh3p1Gl/cjtFjRmscB3/zBZ9cqOsNzcu
2m/g8QQSfGHR2uStAnQgk0e3r9SVD5qpp8t/pYfiaQPx6NyeogbvzwwQjW56kK2nNloO3wlvyeJL
emI9DOAZ07t/LEBzbneLeu0pnZq24pcVii0m3OYReXBr/epVg/PDUXqxaZesV8EF3pn1j9Cj6cLp
PfTz4j90CktyURNE8isacPZGk4lo+fTYbM0cmVqkxI/7qnpRkNtvjX0JjFkFv44v9L6NYFJ+3yjS
EQxt7x4+a9x3GM0k9iT++0GrNyxi/XIv7Nf7Oqdm88w7Wj1UmDUEmx++BZOWhnDPhojlJZO4e1Eu
VQuoDha9OX8xYClyAZkTGA1z0TrnytnB0EoAKhW2zZoaC0mxwqTLrdnwOw1PLeIVO2z9rPwpsoJo
HBozYB5KDrXSSrfz6qnrsoYO89A/5i2TTYP6/BCS6wX4ilycGSs0tXfW3NkKi5zWk6pTNmVPp9W1
XK9XNe448kw1wxRzCytiqsUwHFnNY6VjiA9IsLMnbpJ+ogahsbp40VGq1IB0q6aEer+C7xTxkFpc
KrVu0RQT60aTgsaT93vViWrl1jOI4fgB7UfmCUvz7Cvo3aaw+bRSHBkfPZ4Ik4QWWzFbAbOqmTpz
mIWrb4PAq/i+iD+ThucsW8BPJ07kRTm5s+dEz4XXcpOd9tXExrQUdBhT3XiiZousjQYg00avl7ng
soIe/7NKSsaMJSpx5YfIqoOl/nEXQAHfMgfuU5YLJ1kpXfh0oJ+LsEkxEPq2tje3lsMqzdQpVZot
+obZPgNWVcgdHVWpqyIW+ltcgCTbIiYDZuWnrpEtZg3//PSqOjz5tA3/2fgQwczIJFdAoNbEIt1w
LxawhgL0ziEoy4NbeVvpF4795SXl9GGqVV2vp9QPsDp72J+mw/+9KrcM+MC2L5y3hRjA04aH5k1z
LcSP/heuUyLXRP1dwk21Q7HwYjPNBUEOsLkmqZX4oad5qu/sb/QGT51WVeHB9x1rYasp6xI+IL7e
2wg/ROJawLCdLqRBff6ya/DYdtOWxd9NOog7zLCK1iB5Wfu1Pda6865WJNBi1HzY5OPn7C1szXW6
A0irii4DPoa9WnAIW4GO4VoehBp0AHoUtqBFeLhabM8KajqhKecGb9F+fOUhWC6GWcxyJDmTem1b
KSx25FZuUiHztOiKCSckuJAWKkpKy0wlondVIhg8vx821A1zdxZNNeNJ4pxvnQhl6StFD2NLIzQy
unnlkrYh0kFHixl0ZgrXJXTMEKTpJQYkujfUFZfrk4QGPIkmBxgSMx/hBJIlSS6BkRQihvK/KEeL
O43+ZB87AXvJ0EOtgDCBGAV5+l0v0BQ3nfd9FF32KbJniTGvlM0cqam+gODIXCgRhdbFqZBgWMRU
dYKfmRcJ166QYVB0XIA0MheslyXmAM16kRyEI/sXzo2164ZQ8oMs4HfODsLBavBaNwXjNXzHm6z7
SuMqjgNsEXueHgDMjh0oDNRNmQcbbQMlvJ8RuINR4+ZxlHSbpb32N6gq39seJ8kgyDEDyMI7mYDZ
tX9yg5JX8Dst5NvOt994lxYsJKyLgvnPy+cqg8Kv5MTwjFRwDp4ihofNlIuDkEBD3B1ycHlGrxd3
ysPyrpiNpLyBLHLIOP3hftHnvZxfisvs64pLnskkHJKJp1aY7+CuuXBlscTU3thJnvyqYabke1NC
19dDZqwFIGsX9zKepXsZXeFmnJPAxbRtOMiyyaom4DI/RStMqeBisnByh+n+HQoFznt5jLOCZuze
R4aU5M/URiFLb/1+RAVcEV4JQB3VfWjsoqaHYY76IXuDJeax+ONqj+o1nsTniZbhX4GUXKxbCWwd
rSA6xF2d03EIVpwdcE8LNmoZGyd83kMLofVz3u4FZea/7kbtOoR53/zWMzz41asTjQvDz7LFT7JL
8dU7KRcvheSu/sp0+2V/rnA2kTU3v7IsTeynLkgxBoAJqsORMXo6JikXX22Ioarc94EtXh1eJKjU
knJA+o58dJAIKcjr8BHFumVNEztuJNEjyuapX0y4aHxpdfrAf9uHC4OF5jBSA+gB3t8j2Ouw4GMj
Uf48F9BmP6xpFXGp6jJJ8co3acYE1ehPH4qvB9YIrwSM4tfKYkbLQy3vDFt/X8jyVvEM9huf23k/
XiRTXdtb5kXMGzZ2A5cwp0/vEXudoTbrA5EFkL8iOz4lc/ig2J7WWNWKuTpSJkVsuU9IxORx2pAT
/UpdDJHjIREAwiFdqRwLXlKlH/pOKIWAnwJ82zBWhpTXGYXs8R7lsC8/KPdhBPGZ58jJPrCpBtMo
7zjtoj8Ue4nF1y2t068GkQo5EkPPVC/7RzDQ9bxt/qGK1VHrOJdK5Ycw/ThBH3A8FBf/KPpN46hq
AW+0bgmKVnPuMVlon59MmXHfSfsT9wBuRAjDwiS/WAVL7tsKO5crGXq59iQeHvQh1g5dCX2qukoI
mdaYu/DXshNekM/W2ylxJ96h759CKEaIgNS4bbFCFhtqPxyBbk0GBh6mxvvW4eu2GJ9m96PjCAYs
07dKpD4+L3bFUB7NaTMc2NvM6RgaVenieyX+gH+tS/6dBOUqTdeb4qn0cMMOewLSjNfaJA85jrX7
CjoWnanOWVIP7vqya+6F7uT0o5d8PjFbJIPyvvdEXHFAeVN+LLJI4Nuo7K843cfews4mGzEYu9es
0yOa78QVYrfIfD2+oNVdXS/hXDRrw6ArAkhCKNke7LysBssgd6zf840hIR3As+oe5l9OlcNuDoy4
rIXNO25uEYorTc7SmnvN6cYzZKZyt/5A7O0pPGUSV9Cc0FO/q8q2hr69UgfWo0BvoFiLYI/1ytIt
uemfmEZgsPAxNwvZEm6lWqGg7Worx3NCrskiHIFkhSH8H3Epd3wnMsDFg4SX3wwRqfiua1gSVLue
lsTJgSucBECP/J1xYkWGcJwPM0CHWuykD2LjBryY+uomg1iaJst+vtFT4Z+ziWmczsrLUGkSRuOF
cX4sNkE4u/GqxlTWvpy9XdAztV406ZbqO1rM9hVJl/kakstCBc4zSA+tOSbeQxelTSodpYQ9a+FW
FBxlMjOxrhJjZ3n3ws+sQsNIO8CJ4nPi7ZDXt3hYVTM1jPcz5ud0MGiRzuDNIkpQx2/IjHYDGFRU
InuHRT+iTrNjGCFbyRWZZFXQ1T2ExKosDlJxBo8+wYK9Nby0dcROhSQ7RxMDRVFemcR+vZj0FRsj
2JpY4evy498q+Jravo6QgU2RdQHih4sV+3Eb296gpDbOft5cVBZwMPAf43Q6vdq2Kw9FbCZb5EKr
J31R4LmPjp0DJmYMJZyx3WDLcuQp2Vh3ItcfG+BE7qDHYmayzoCAP+0laC9YCVR9/b85lDEMDLOM
DAkhEL4n3qv2AQRKEGOofr21hfKXqhbQWgsa7E2+dS6W3/uN3smy6878kMQmqbmN63L1xoo+A8ge
KSQnFILDbZvRgaTnN0GR1wRtDySnCeb+Ct0OJATqRzzde4O64Xf2TePobJHNJ02e/caMe5/Nqtv2
V2ts8Y5VmgvZMJq7JgxiHRb+26RMEb2D5ekGyK758abF54s+8H6rAPw38KbTnneKVFQV3qVfS/6m
CZzODsKtBzuR+pO+35gU74jbSwnYAwl03trbw5h43lO5DF3fLJ0WXUBMvozuK2yU8k+K/WfyhRuN
caO0Bl+EIZB8JQxJqULlEhPUqNoFQdBttsOLTCC4U1E5zqojHIn92wBuj8wXLDN2s/TU05/25hGY
eNqrtI4tRCwof6cWjZoY0dYct2vsaq5+h5L2RuuGPPhyZtz8E0g4FsE4eRcxK/2CkrfQhPiHXBBf
IRHH/HAz/NBEdkvo438JuJ05yf/9p6ZPl5feWxiDHT1JWnEuTh+SMHV+raPVHpGNWfioeqfbdXWg
gEsvwOLnLivqSwmcg85L7JaCm6bkCYGBgyoguc9CmsVLXWWF8t13NNF4G6zzN2Fw1LM3et0SpgmO
RjlaExG9Lfk5O2XDAPezNgDu9PgUBav/NUcfORuRdgFq8wZK2I0NoEQuYgUUZOWLJFRjhXSGlNrk
JmDJs+xp/DaInrQpKRrsAftd13j3xr0KP1sa7AcZqzqXIFcAfsvJngChf13Hm7P6vpHT76WqKnc/
ceUuS6GfEIiD7CJsPTZqjjawZovb3UgF9njIRZyakFcDorLSJPnf1eVOg3Pb37xLEeTw2mkbI/AZ
bzKGbk7vyz8zHXxrqvEfIMz0NeTWtrmz4yEOI3LPFQFuvj5wI7+oJYvhle8Fe3vHPjOmK4gW6o0W
atN6sc6tCr+0b+DsJyoDlQUvifRQoHnTjtaMqdDvz7UZFBSJLGy9dVK4PnSdE0naSQhtczEuS6DQ
Sd+EJZdIk7BYk03YWM9KjGgebmvwShhF2kRW7svQy5d8GJRr99V3DzCnSSlnSfaNcs2oy5wBmGcC
Ww9RYd+prwPHenhfEl2ANC749SfZa8DDARS/4qJQgmVLaQ0OeV0QoVEA5mwQEj96QuTJjYq5yYYt
hmirDVxjdZ8kLyyVQkDvqRLKjgllX+/A7OnqvzaUfM+9QS/aMEJdU219tigsYjQa0wHFVpgo1dy+
hezf5SOS7h+W6lijO9+wPuebPN3EtT+b/Wi4Dx73Fce1+lNxR6GrqWu+hoVfRRMIV1vB9sMbumGE
7FCo6qbfYc2WOtPmkJ5ywAntyAfFTwqMvY4vnETWAj46GR4731N3RQC1M2Q1RoUEKO/HDaY2rdB+
lGp83AoEzcqimM+ZiM3A+1Bfsmoh8GpnaEwJrSKo22zPJLwg1ulnR6YYAw6d8apSk74KeWr+Rv6/
CQtBtOMLqkX5z+WvPr2frmsnVyCUigAYLSAMJC7x3FQMKcD1I9npVD0ahlzPVhaX3mEzw49ZEmNK
lLLJhSTsqWamtJoawUSitutSnHgbUDFshAvNkcQU5jK4aN/MHUglswywJ2423Gc4Nkv4jkZObNxJ
xXAK3rkiFpH5jDnlWGBgo0KTWuPDmvvt4FVQgBGbYlNARbb3lFAm6/uy47DfQZ8DLnwX5ixMEVU3
0WfsGsKO1goYlBVA/UZcYTboUHHMuw/vWwcKFEYpUnjUg+9O1Q/I6tIsaMEQs8jgNK4BGX60B9Dt
FRxBiMJ9GGQ8gyWhnc845KobC/jL1Qr8GPyFgxWPanC/7vd6J2skvXZk20F5ANfK6+iUY2jhBV62
ak+dO2n8fiKrxsZT7PrWDnnGfYLLh7bCQL15VzVynf7jCuDCEiqMXUo1sUOfwfc4INIwH1dL+y6Q
n81VR0Wqcdn5G5xg/z743skI69wwu+b/QQHiu5UnGDs5n5BcfDGuUFRUD1hRPzWdlRF4VqYG/kv8
32I8lOzedXwQjdOdsxv0V3Xw9U4TTyPMrKiXEhuGGdYF9pJCyv+zrcxvUCNvncsJ7aUH3c/QnxIh
0u3XEJ+PluSxv9kLSncGiW2YLw6wc9wFK/nKdWHDTsVZanSzxEB0JSDv+oX3/MgAJSspRZzJ890r
RCoAEjwPOBt05y9o7Kh1tO0XqP4qidvfr8076SFWrsvArg6UuwbKkbAb+Oy6d0Rd5jQVtLRMmGwy
xy4EfgYppi8xHNR6BwRBsCWZl2lIGp7D/LYCU8YYoUe6UpmlnJjXvf0f/WvL2LlgHXlwpHHGo0PF
KiKoHUGYKymI7/NWYNTflkDbWyWYCBCOBF47Egxmb+TYmg3acs+4hly7KHwGcuvxv/0+rAD683qg
yxkZfMYDD2Vbu+WKt1EgJS/Ca1unyIE2cviDex5J/5Jhhr6UYCnGN472oSfDcD9NtHlrSxWjHR7W
/iRkqQd/WrwFadie0glHlHTfELlabl3hMdFuEMW1UaB0dJfq1TwT1TICPdGrk7bhlPHjs02waDKs
ctuKHXybGqvTIqbeQLucupgQLKIzHRwI2P53EY0DfGCTkQHzSCckZg1P6m8sM2xWFKo95LoqcUyy
ZFtzEOjXGujPUxa8MdMMzYXMJQTN1ufUD2lyckpXwRAP5FurbQG+Xd0KLVHnYItbwiegIVA1Gdnm
ykIb4Qq5jDV+NplShnUFM7SW5oi+kI2u+ylsb4tjl/U9YkXcsiuMB+Boq0MoaYNOYuht7b9XVfiW
XWqttYh7q8GIi7h/W6qxBAFfdG6U5UpeR0/WZHTWg+q32J3kKMWqcYBa0+nmyv3Ydg3p0WtKL2Ju
r+FNg0xZEO3trA57rZcadiEHKO0l/pcHHlYOTqJA3rIcwt4nTyyL3+MxTZ2lVDAwcapZL/MPS3NC
zCUu3evKtmvgSoc/0kG83ld+gu5pAfjvcFjWbwtOBvhDmUr0YCehJpU6Ce+4cceFxkxRUnG5WyxB
nSmpdUP5q6WtUvBfRQzNAlVcyCVpllWgRxWSX9VoqSzwwzwKUYDc70uStHXsQZ6c48RwnikkWkRp
+2qI2aky9bFycUGSX6rs85VbYsyKK0ImNc9alECD5vq1DpaHc+me9QMnQjzA3jC2cVmByHoub+FL
fviWz7ci9s0HJECk8ltBoElo9xG3crtYAkm1JeU+ufSdqTSTXtVT7BR2sX8H0wG2IbDi2iIvf0L4
UtaiKEFys6eo9TE1JwGMhfmKI4LwVOwBIPR5WH1+P8T4SL5NWJOeeSkxfEqoE0oZlCN3QBNiA0oq
TbgiXF03E9SiJWhzinVOzPOQP5X/8HSP5DF48xeTt2Hkyyy/GfRu6DSD3hCQ4K8XkAtsuhPYrAvt
0AcNdysqHJYJ50g7uuuGgBp6IyvnXKzzJDMFVP6TIAUWtJoRv7J3EZIpFfiN9MCeb8JqXI2Ru07A
w82bcrZ6uKnsLxR93XB9uwpTWJ+H2y5XrYOGWf6QRegns3kf2VQR99wpp5SBI5WEfsqZvw3zwlZP
IrJM16K4hNvXp5NdnVldrokYTFuBDPFn1seaSgSLqwVJwK5QevKdipIboQ2hhdloNGyWRCNucUs7
M/m0LKTneHw8l/G2Qg4xJ8wocOtof2sArBQ+qZpdfPDO3tB0Zdps8qBww9eoWQhRzLyCWOtWo7yY
PCPI3iFMofo+P7mRm0+fwRhiX1lCCgbPwqE6q6jqRN+VLuadS+Y6YkdHZJMvxrMCVFQglKBzcKjO
JEqZ49d6A9qsGcR/dOnp2tAk1PxGP+vVluGvXsb1i26G8kO8OcKBSX24uKJx//c/EVrT4iqA8ztC
LoF83Y16HZrsAmyFbWAWNI93nOB8XxNHdyXm1g0Qn8N/gfgQXgLphZIdMbJvUcDEvpG7oPAlGPzX
bSAV4o2SKqrywqBjixlJntZXX/Q+6xAzgKbGzQbfWsCgktqQM60N8cTUg8e3ViUZ/Y1TjuI9Q33f
otouJvcTXw4szK257Q+dypUwh8ti3lWA8hFprchmOGrkhqC+R/M3rWTBNMV8FaL0r0GL7EZePMZ1
NYj/hf9HdGKQwhuApgWXtfMmPa4Raf1RefNE8h2+HmJIzjuQq/8xWEKlJRORZKBPn/eaC/S/Ivhi
y/dncttGtS9HEvFUp7K8hhT2wuemmFh+4koPZ+YZ59kcloXsVjZ5R3rYVKCaKqXvDNQ63glVDH3d
yixBdronxQ0GyQQOrVEz50j3/AYCWhM5dLrOr9NfAIkYY+PZSHQBNADkbuVHBSHcQtZbpj/xwH6E
byIEzM5nmfLtsajZP4lnTu4de5ielvM81L+IElIErOfuU63yC52gG5H9A3AJV9gE+cYDDawGlnix
3Qne1hrcafpFH4cRCqbaCCdIa0cGvAh/bwyv+sxiI7NlTYjwV7fbF78WoUUQR9W+dY1z46Y6ID9j
4NbIxsmhtEF1HLdsgFwBPTwPpkakJJlrrL8o/RQrngTPgGpFcv7WwtN0eoOFuE1qenz66qTvEBzO
vXTeKoJxbQYoWignN1uyBgeVl+yOB/3zpwRNMhvUz47CI2TJiv8QA1RzwPnNjOKWxpC5jLEQkokA
D4L6v5eagwmTXHaCj7g/MXFPkJFZAGZOc+B7bkKaFbhCnN3DvUwDGRiXMkReuC1fcybgd8uSFEwF
BVZ6i24ePhPjCBw3YKLb5qUnq/tTeacF7bHnjtDzvA+D6G5Gbk/f+wkEHrGfizO4pfl70MqsuAQW
d7xRK1FFV/Ht/xyCM+LN+fxoXjkmgUvF6gzmg3iiS6EZ4s9iqzLyuCZC8aUG/mc+ah/tapPsArkW
wm2D+ew1EhWEs0BM31hqXm6gZa+GCLut1cZsYlkFQ2WfQhzdO+TI+q0XNAIZHsj/u2kjvUb/R4vi
xCtukCBqr1tU9qK0wrzMhTXrH0XUC/5RdBG3FPx/Ng9/Y8ayo3x70yVoCtUFHYqAOSRuKw1/4euc
nmOfkOyP/kOH3mT12cKIXV7PzWnAwxsHilyi5GFofEsyv1DCML6hCwQczbMX6FcD9U+cEhibdDgh
9L1eBRnwouL+LcpaQXBgoudatYQ1XJ7U32FYX8kPIdPC2z8FJiOnq8Zv+knwSgQNrIhkU4Fz07xW
BFzcDfzXnrhQMAjhkTLOycBDBXSCQe/P4uJUUyyd05Olk+LFDFXx3jNFtOUzML7gVKxxeZnAoOm0
2RhCfZiLfce2lz+NDskqbtaTebSi5p1mbQVBhZ/VEaHL0OMSIHNxTHlMBf9wGj0Opu9mg/MNUUaq
XZx9/2y1dy2AQvddrcO3V+HB3lmO9wnCCqvcj+T1hIqaWFUEjIHWj5WvYzkLvFqi+QMiiJgJbLWt
7NsENv1tW+35XpS98q4TtkaeyUfspkXB/J/5ENrzWfMUxVIyGOOWejtwmxlhLP0E482vAkSK2cji
2oXfYpzh4MA1LnrVtOZFaoEP71k0PBLFiznQ6dCJpzLtr7cuHUIsnxHnFIyZq1ZBZqKZyaxR/UFy
UXBxE7MvD98hFCa5GBZaPtiZ1bZKtMg4QPfe49vMKMIifRtVtfg4zxRx7s/xR6giqsi1wCdem0WZ
GSYMwy+OwGkXIAaTvBXHL3Akpcwsxi9RaDWRnkMpjIAKBANDcxAnS23q2wohU51KJWLfSMNSm0GD
apMMDbEdDGGDmTrD015kBhQVk29jpsf9Tuds17uKQ2vuZLtNlY3tziP6jwBtEwYcPan7dPEORfaO
Z5MPfMSrnCBE54yjQq1P7aAoiYVt2kOQmMVhNEIqhNY2frQLba9sR2xPNmytcwEXZoh8qpWOnVPJ
IUA/5CesytYCNNRby7fCShB8k2xB9z3GITq0aZLzmhL90eA0HX/khKFhUsfRoSGSRjKpouken+Gb
9ePTbVxHxGpZtX1+aNgHwTzivWKqE47p8kNReq/bIv/obUL23yjCIIu13p8lTGe03Fxw1/hrq2Kw
5A/t3Velbj3xa3Rwmxvd/Buf9mLC/eYBljcG2sm+r2ld2U9efRDB9Dt5soC1g/azV20WqEr1vFFq
1YUPJ3VlcOigG75sL3k54WpDJLSVjWVP/12luxccU207CwKPqVblVyqCuVbaROXDCgiN0k3spvpk
kLUGWqj1vMc9F3Nk66IN+0dy2XoA6WZfM7QKN6WHUH/5sf84Oebw7BKYYMtpxGoDK1T4MQzkagPv
Yo5E+Rn806W8blEV7VlIEpbEShl2UqRIHJGr1z0SWBZM8KKCquI0xF6jLFL1OmTnYjvoIr5H0DXT
DYoBhIjXMl/N/7dQA30z6oXf/3knCMDeVZx9s50G2XxgvdzzKW/2dPDbLIMLdwZrAvqrqOH1BPZj
fROA+kC3dncuUJ6lJNkGcm1Y+pk/O+5AUkF2HmsaBWZdG9qbyxI0uIJ2VOBe6zuWIqHh7oCwgXN8
9mMJDnjDzwOsDFwT57jj5SIxuqLSr4sFceaPehXO625h1+iqrNPBW6LShV/Ece1+t9dlk6VOfxQ3
ATQmnlgLorkMYzy0+Fcnk92p/SAhMG31a8VA5RETqzy4apj2bPsnlEI64p/9dtEqmbxb+ezkOiHC
2LmiycmzUKbADveRAuWBc2YgNZNfXXS8L4pugd1qM6gwD2gPGjj9UIOsa3ujQe89a0Ri174jS/st
272m1Ay8DPOPk3pfyqEOH2t8TH5nFIPk0FNB9Kxtc8aXZyAbat5usMBHQf/blRHNYphq/R20bFpH
Da5stE7XTooax5r/+Ivn6FJZ8nYw5XZ88uEhz9nTUkTwmj4itTeG4xVfM1drKRCh4FvN9pFS/l6F
uE+YFY3i1nbNjoxeleoTF0HFRxUu2bk1TnsLBwwkroX8uNldsgtjVoOVlQkICqk7REXMDlFV7Fiq
niUcUxCkDw75gp98BRmgO3aR3UdhegZCTNaPOkvZ7DCzDWPtQ6ow9FD7HBNKQiNpTSFsN97yh7Km
kY0UEC45QDh44tjNVxZbsY9ftjPcNyR5bTwuZr17ApetgAas07hA+BmqKiNKG7ECDCj9E2ykA2Wf
LR94WyOvQgNzfGIenJmqt96xpZFVKYcpjLkee3CaTcVP03Vkt+mHbFNL6F38vHZMnTJ9sRh1JlX2
CPKRSuHtanBmpHSHVOPIAsVrGHVFKJkzvYvXQTdqsufXjsiw53eOSws4ZZ7nbdpbX9LftxBk3xdJ
BtUoOQ1+0H/geDpr+7YbaGK4WqjdEU/Gs/dmexM/PJ5RuEQZ+mpvncvxD3GTLAHa/3LPX2pwsI1U
lvvKzP2FtTj2S8FDJy0dqPvfPZcTfepMOzvjM8KJO8+JBwV77wbE2TJk6At4JQc8YeUB/kbJbdoO
iKKP5EAwB9q+aVyDNml3Ptig+A4z961arpnhJNAhpTKMs6ErJbxHAFbPdLNZSXECBmE1EE3VNv5g
XnRZxqX37Yf/pNxpxtetlX8rGFK4Z72EKEFrP4iTERVa19YhQ29VTM3B5Lk0tcldNre9kaywkXfQ
ewCmn9Bvm0/x1nua0V/p/pRKc7Mw77i/Ns+CmWPW4k0XY5SqFkAF73SIT3fF97vZtJChIZT++LmO
SToNR+XANRBecJ6jOR9MR8QAbepWxOC52SIiztLnRwKItvciha3TZcK8/KqYw+/TUQfgbFkK/gIn
0/vNGow6vH5iL7buK97doR9Zcy2REw2jdeNh+q/8FlkTAzszr4xEGQ+CF8BLRFU7R5WYQbwDctbU
lSxTTeYvkRJHY53qE+ya3TMnLPhUKuJZJMHAAyp1As7gr2YbKEaMunWebJZTlNKABBz/9eOib7PB
7okxbEszZUZfO82jBdF2ZoDQCMIb+LFjrK8NyFR+cWLyD+w1PKz8u3kJybRa4AZnIIf5C3Y82vZ7
qSkNSQ74Wf3u3zdH4yySMo4TILJbzqJHhFs6G11nISsfjR5bFYrXuVCiCR8fyxaH3o1f+9VljDf4
2LjQiblPU5WkP89Quh81caFyYOVQ304oU1LKE9wesxhCwGJ3wftSof9cHDXVvkK7RlJdSXdDiwYE
BQJKKrs3/lC/z395+vYABlrjhQOH8yXtkMxz2xz+GycMAMXWASMQevHZjOrZ4FYuBbrv/KiZ1/I3
86xWD+Vvce1reEi9kt1GdbAdmhOHsik17OggI1BjbqczNCiZHyV2lFHZQ9et+VZCWKTuMR5Ge8Gb
qiWcKEEicYrJSJUbJ2ZYFFulqkapT3A2ZYFYhuZHuXAO8nUt6RyPGFWWF1PGEIx+7YQqb+1r+4Xq
ehv1yzO31oegnr99lISBlmW6KEAKENDMdcSxQ+nrDk83qIKc7lyGDNkJpuMT4SUehEBHtifV1Lib
RqRGd6B9b0cu2WHD/6IiHCo5OS/68DSP9mkoDsVLCEiP/MisiiaKB0a3k2DVs2rWYfQXg32EgZHp
Fw6Als7ZtFiCxdmldBgAMiX9frAkCXZ6ndxwGHdADQXIAlRXDoAhJhCYGDTVMyEA2+j2VxYZvxNL
i5roFVnHQ8ohB0eghAZBWp7QWr3EXdCYoYUHrGTpWboAzu33Cp/xqaUQcdAc4TDUGYjvIMOqYv3X
x9lOeRxeJ7/x8TQVyADBiUXgvJ0l22QzA2Y1yJRMHfNswYTot0gwldhQxVShztfFCZ3g1USJ8aJu
8qQuCTtkc+OQqaV6yobVrtCeXrNO0N546tDk/8R22EXMw/wQs5oHX3n+bpmqXSkPtfCXqkjwfbwt
GKDwTWJ8L7RMV9bE6Vls5ejoQv+WKVdBOAnMCJwMrg55vIWS3cVRyi0jCeZ4Cro9QE62Zd/WqrvM
0f/WNwZnm9YTq1iwsF5wCkku4x9YDs07T4efkxW6P2fp31osoS0oAckxQdh4KKuLB1JTJYCHrsZg
epmClVH3B78GJ1y+yl51prE7+ejCbHCX4rZqCWjXBm5K8zSGx7waTrJTZFdZNFa0gjYieUe7fpiq
3bnmzq/OwBcySqOAbgmHdaGJIrHo1HFKvtnzEIiFzTVefAC/LYFHxXe+t0iHyuWiFU2CkW8xUmeN
KxgrPTvKp+AoCXZmZ3HhHOqyf78RK14IOKPxJ0gy0MuSkyF4r/7dhEArA5chZK3fC0kQmjwai+xl
MveiOQutv9AoZzZgh9bdKqc9hbwHdYvUpdHx3ek6+i9HExOFmYC2YuHApn8W1paOT+bIY+PnDUJM
p7cY+4yQSLKJx2wx4F86anLZfVBnDHF4erxNiAtzL15QdDjgR6+agJwTWL3cATI9WqW6Giiy04b/
+LfGMbNYeDMrhicuePEiUN0u+Yp15DioCq0NBsxRynlcm6XN9d6lJjrYc9JTdArEOSG9N5i59JN6
FQgp2lX82dUyS1nSu2CSDWI9OE4uZ0gTrdlePQ3HF0TNqnFA3qvbWUI3jsLNwwwk6l/zsaMe+Jc2
vDSMYJ0aF0V2k/0mILt2UULoIl69J3VRb0wjWJRmZ9RIxzw9ysfG3Vpth4Fx9/mmUDLp6JOhlJin
+vxEOaYEypOC6HurtbQhFkHjC9eZ9Cb+SxUjXGRDff6sn9nHn36ZziqL02DPE0DFSVX0n38NP86T
+0g+RymPcG9ZhBbWvFNyGTal8vYZ0cxvf4EOkioZG/Gx4uCQ+Yqhq//+W3+NXzCXLczwfg8XluSL
kT6w95gQYFLZMYr9NJ0EmjXmkdmWM2DOBW8gdxcCsEUJIaF2oVb25uyAwt1SpoH5BxV2VnSfrQ3R
Lggve9DuJ2R/hyl7TG5ekHwSuVTg1xZZ93Wssc6Oa221SRr74no+Cnl6rX5IqbsOoACA8qBcc8BQ
fs+FM4dBsoiTAog8kNbuVnZuLf28yyW+tz93YBMi/bCIbDhejl6ETbtOK+sdMmW3TjduzGDiIDBR
COATlxrmfDkzoi+0Wki/Ef/+gikAASCE1fDaOCbx3p0cPVlc6lbgB4ZPA7lDdXtFebFKsJlhzV7G
aNAq8WnCAOMSu0QB+kf3Cu46nVrmf/LVTIVP8quRLTDpIh9LVVHhFb9IcEnHjfAbMv3jVNIvQHG8
0KmVEMn7oKDt0EpoHcKScDbXv+dWgsnA2da8hVIqPofDWd2K0wFtdJQtLpQHbhZHYojdlRZedEjU
GIab/ek6nfQ4pQTOcPBmdc22jBERoaRRunDmHIHfRRkKPBFrDBrG83EJFGVKuP1lL81ER1ishJ8/
XHEejTdOK0Ko/Q6g9i+U4UYIzhNv2TYDA3HY4xvyIhRPz2SnUs0E+qHac6wY8npligtPUV//BLv2
xq6sMQRFOnZt1YrrakGzCIM/cF7xTes33+M7UdXDhetl+YQ17Dw32ETs/fMrZ/WeE9Rsnho+T9x8
Ft8I6uF2TkkGJnVKwp9PUpGd1o/QsUpZYgIy4apLY//ScFA+Hzl6SUc3nuXL3NKyBTbpkSFUAM6E
+id1LMN8ohdl2xNOoyLsQ6fUELMqOy6cCtaHHwPvcm+IvFLhWQ77fp8xgSlpZ8WcriIwPzeu2k6W
1xEHGC97XtgpNj5819biYcst8shpIsS2c2QeHy9jUjjm9I5H7ghzLWzbcnrOJQNMdVNFuPf/SB6H
5lw70IF7fuZMLza66RQ+kId79G6nd0bkWlV+9EC2hs28V4UjPVhLD8XhLI889qSCdIh0fRAyDcVV
EN3MxGZqIjP+5IUhNfFqQVhz50xBO1LBKWi610lfKJuSbNTOfKMYScQwxxKBaWZSzQVD6q/Xjc/p
uZrp7CURsEx3/HkXaK8xZFtoxZk20Iz8eGGjCXHyFAfol+xmkJo0jzBvbTg0WtKEEXiSGTBsGzt/
N24COAUsBZjCNvhPJtoJk4y7Egk5iql7VrLs8ZF81qCRhExz3F74uoeLxxdb7k7B61OYuO9V3qop
uEIV0nR4se+S7peNWbAJfQdYSV3lFRqTpCZkMXC4SkrGvo3JcRcTgAL7pCRghBeW+bGOnswD1vIF
CmE5CtgzOERU0q+XO2P+2y5gw2G9Y0O99gPbyrs5KgG9FfaHVaDxxj9sJArY3p3M30xd1SZtgMj4
3amvt83n6MopYqQqPxxE9X18o+NfFiyY35gpwPFGNcPp4mOdoel0AcDO9Q1lBdAAxTCgG3/iwSbE
Ns3p2XEy3TbwJCjeJZ5H8SwFskCyzbpqcGaCxCyUnZRdYn/7iJs15OGsXLX0LdzJLHxc1dX7Iz16
nUJshCV8+8jEC8i30fOXxg7Men9WIrFqR38OF327wV81xPgoyBVr4NHm1u3MulPQNKHzlXu0N7vY
F2xgsnMNriPCnXzYOquXclaS4dOFcI3A2LKQ2Bc1x2/2sXCgnVm37vVdaMl+eZm0fQYb5t46B3il
FVcba8HHJhIXTazqCfXC//wqLdHA7F7n/p9GYNorVft4H5Vjl6VJHRfdhf3Ng3YEvv8e8Lpif2a7
6JQ+Ets/6PDuQSyRb+No5wFfr/07U5BY44YF0dN2xx2tVFddVYZPb/1TPrSL+V/ZZH5fM0kD8IzR
D9YdsG6iUCqsCI7nNsmPBv1IKfgmBEUakfjo7vNQfv0ak9N9/rk2jG8bKN0JlS+cq2hwEh/XzviD
hWY4+jg+Y4FM232TicAjmIJQa6t2T+H+WcM+b3mpZTHyIoUm4am1VmGgFFOzO5yEq2v6EmaLvwb9
MTkDh3K/agynGcsweqsmMvFrtCQ0rUnjcXOzGf539p/T94txOp5whe74Gsi68XpQEQ4ftFfQVcK0
QAHGFT0rmzQTa4b9GuE2PBEqBGNOp0Nt9FZebJkjYsYxprUkzMUFh8M8EZ2dLMCfYe+ZygWIEVI4
dSJlTChRafuJJcjAr/oEkFizoegq6rXDjBRg7CWTgLfLDfGQYGWWwLOrVwWhsyRchQK4INgQEk6L
rHUN+7g+70YDRdsvvemS0oM4wwL+HvHC8qu9W8ZF5CQZsmA3LBH00RMtuLVjCXtZrhlZNhuxif/3
VEwcpkyqwGiZUWJyvQ1alNptP5ottn8K30UgARQr894W8+bgCO5RlOQEUTNTkCUUel4PfAKZwi/N
sDxOeftC1q3LElC0PWHKh1sVBnVMJaqfhpynKKgohpgXRMcbltI7nzUymjOTHWfJXJdKSGgHExKi
OrrtUS18ZQSF6VRRz7FQWGATsKw/axSCFtYVlI8YSAzjXcP67fG8DE/sYkj80LeqLqw0/+Kb5SuN
pO1ZaIyyrOly2ObTKQBkrkqYD0U6VSOJfZn9DS6GblZz6hVHi5UvHfn1vxGCeGB+J6Ff9P7JzZLZ
pWGobs0M5ivcf7VKR4fUiKBB4/03tj/9JX3EiUGAoGZheZeNz/HjPBgsvoBFSw2WkL3V+D0zipBE
1YW5iab7M2BonbBUP1wh/W3U8TZjqzuGkV8OsVZJjkWNZ7Ki+oeh0P0WHnZ1L0wp8w/9pCw/q0Rv
BLpyIXRlES8pNP8I7sZQ0TKwr8f2MxWn/ydO29MymbOVyRDCOclSfCwwAiTnIgYBSHRUacX8fkij
oGwaCzmwCtlTm0Sdmj/Z+WRufZoMEFqTnURJRGtJ/gpFhjfut8unDS0F7jmKsAQNp7iwb2ef0Cdf
Wamkuiq6FXdKQK6yV+pGA9RTghtsSufD9QrxXoitfDZTLDvz4qtzxZOqWBR88uxAlqb5E8QklUfp
M8GEx+8D5MFTSzxlHcvlqgXxkcFbyLAnGYo3Hjn8zoZZaXCHO7NT+2CuaKNipulusDaaGbv4uo+F
ojIi5vc84nimmk4bZaP15crRT+b0TQRPlJl4dhq9TWDM5W5ag6WwTXB1ptfYAzXeOkLVA8A6LyV5
XOOt/bpVRaAEnwMt5+H5oRb0nHB3ArzmB98Hxdjz9yF1NtZWxBeNhFo+qWrzhg+iFisr8DGDpn4I
/yhbrDG59L47Djin0R1n1UJo6uE/O2XmEKeYT02YJTFxfPoxAIiQBgxpdNvOmOlOE0f5RlVbOCTe
HKhNI+Te0hq2V/OwYUDFmCzSuWRF1o/xpk09wYOglU9ygbPJvKNb0gRo9lGK2bjNOvtySTYcnJA5
lne5AmJriCFWV3+BgUGqRjvEaNX9WE0qtv+NbRuheKdoYv9coZBECJrxZS/Uag0LVEpsWSY/bpkT
26ajR4eRpeBOEvieQUtLVAgG/Ba0EHidap10EWFiUhjdIFK4YVExg5s+j8gYYfkArcueuB5yGA3d
/Kh3B4hD7ok3w3tfsS89gcCW9dhjwGG0jSpcxQ3f3AVT1JXe/qV9iIaQx36mx22DNd+ZkwTJeaS2
3Kr92RtaxoO2GXpBB56k50AVqah+i51gF7T4aXHXIMzY9WXxBdf+cttL9JAhYy5hrrbHWhpAVci2
wCW70DjGtqRuEO7xHkK9oECKc1/D1/q5I0Y9a371FEHkqi8ElIRQ7CNgxA4ClhB2BNxDsjp1pgxr
C+d2FHN2dXkf4N2BGWtpQ9hwUUAoXZs+Kqx0+bqBpZahvdgu1AZDAHIr9Of+Qvk+B9F+QIoC8bro
zmbA+VY9tMlmDASQyCmf0RXbDlhUXK/7H/zOLw5OdXc0QnfQYM/JjYqRKMF9BVtQ8QHaH4YnBbbP
/DyAkGlBfZv65iiEE3XBcDsDh1sgyU6YNdbLE8LOS96f8VoZLHFsl+X/PrUfNt9WISE9XzdX9C5B
DpKNFROtKEr9Cg5utTVOicPBvaYklWHQoYdA7RK3Z9PgnrU44jnOITP+e79jUCdazF+M8Xu0+GaF
dws5ZvQczC0E5vULWhrYkrfGDW9Sro5iQLxiszofh0AObG4zlg24/7avY2Y8O0VRmH5V4rIcujQm
DxRRZm2dpfTwXSDIgLwkoyVCieiiwYiSBBgu9wS0h4aRRezDEJiGKloU2NlHngv+5NCFL0xoKPhm
dRiozMZC9PGfsOrGJQHVpKBLXFToHaPKb4Wo4vVkerRC0bJOCdTrlttK4rHb6vM9J3BhLEHMp15K
tSFdlJJYRHih8LEGL60D5DYnCLW6ody/s1h9PAAs841E3G30A75WWmTL8IC7zh5yKqMWc38jrB0i
vkVOSaHR6HdzI1JCZP9zBvSY3bn82ePvnG3odZOtUQLAoByMA2TsBfCOM9uWb5/QqN5RnQbPN2+y
AAcT2JubUE0qeF4xhJgVaZ8kwxS9yGl24kdg6w15j6kcitERw/fLsxa6M702CRN6GOlYQcMLr/oI
ustBpFu/8or41JH4579QIq4xV6kZxwmQXrqkeeWTsN8jixPXHj5DygeXbryg837+zGqXIOWUW+3R
UQfwaf5aOAqDwilF8/ZBi4SQ0tYJLXkmbIKBQ4lhC2WASkkazLNVzPFwZm4iEaSROBfnkWWVCnSD
L8THi40tl3oXkkUIY3xAiAbklau03W50Whh8rTgqUc/xP1OyeNtT5kIqI3qoayb5yheWLpZ0mr6g
8YYk1KjWZev/FsLxSo3A6sn1UvvmmqXyzl7mcxzH6eQsNIxzgDdOFkuUvcF2RZC7eC0u7HGo+pS8
onqSr1L+ciMXVWY//O06JdkAK4m7xF9fmj8C2MZkoi4jXpQV9cidIjotG+3I51VADQFZ2jheTOql
T+LfqFMv1tZX+QqeltXqIKtkd2QFvo0u8piEBDqV05vK4Dlzz3u0EgbrjBfZsQDfY9HR39ZI+lDO
bPxJ8+AdRCiwxI2G9/ZSR5gSUkqo80s37/9xWTHHOpaCMcQOrFUVAxJQ5XFsLhMmr5+xLysnTvUV
md8UlUl94R6bONbdQbuopkrv0mXqFMz6RJaVATrCWzohN/CruNP1Z+/YeqxPABf8DWwXrKkDiMtU
RjkLmDr5K4hRqErSAH86GjyHuhSjd/cfhi8ncJMeNbel9VyGCpVciSLOqbhebKDtGjlBNc/npYRE
YBgM6rJvh+PM4xMEAgT3lbUlAX0W6Cqx0uX2qVEMUCga5h1DYWeBt1nb8PdNYc0+bN7IxU03X424
XofoSy9S3E9YYje/jZY7WRK+l4ZvI7NCo4t8q4Q/4Poucgb9cQfnPDU0t6xFm9IAcXcf4Ha45kaX
GIfEyGOTmk2xXW0M2gUd2NoAE1Ge19e2aCOIqPM/qipjxnJ9V+QCqCU/pROhsUwwO2xGi3Yy4pdu
DXYd2GgE3aK6WlnJvdCzKYKXOfLoAVhjm2FerLjDUPsEOnai4ktRosTt3K5ULYtSh+HuIYsQF5tn
s4yM5kMYxijdhS55y/1ICdPla3W2YGFNWKGKJZT3LQsbmtcKxnkJSZ9ddBXNyX51hi+3qWIdjN9A
AqxrysC0M5D0qCbjM4SZJ015YT++/4UmaTyfUDp6jYReqM8M5tAee/g0gDPZW6r82it0utVXF/pJ
rrJahc9K38HHWcEjuKLXeEWpPLOmReEks6whHywhRlvT5nRVoEjmDNAac7weIT+5CcoyGRtLAJw3
AIIawIpJH2a8fuvOdmvS9o+NXFeYE4H/23AedneGxJJI9i2TEovdJpJkYHDy+s8t8uwscjl1qAPe
76kHEsaPlFbw8O2GYeY9Jk/fTlIP/Tri3W3Ml0n6B4Wi2biiqw7xjbbr2QziPkNByuEuHzvERmU1
OcIWlZJnIcb7MiTAPPhlN/8+xZ/X4UYiOik5YnGIwlYlRp3diKrNUX/HjKvB/I919hdb/IXpRAda
790gF1fjVlA3VYRspZMQUhYdX/OYbwqXxGHRiY76YR368epnAUOXqIFyZrIxmd29AyHLhdESjglJ
iCEbgrTkztjRhDYKekgkmFzjm1vyX56k2m5Zvnu0c6bj5MKVGnp1t2BPdRAyFbbKpCrXtfDXHdSr
JGFWJMq9dAEM91CRvNVCrg6liqSyl/8JyA2QprRw74Zb7VHL2L+9wLabFz2uR2oNwr34GUTxuUbG
XNDQ+zEHmpCmb+klY1JnpqxOUgm042OwcugUWCwL7g2WTwdyo/1gF2w//NoqmOjI6qInH0z4rWcO
UZNneH50E5Q4xdwj/jNiv3ShDaQDIvopmbuxUJwtWBlquM5bAJVtp0I/wOxlsnRixf/3Gfz8/CUV
2c620o7OpH9lWEiWv4TVjstFw0MrkdkK1tknySwzdO90vg9rKhQ/HVFZTnxOFqVzqCqWBF3bsqjv
bP7P5Y65tbYt1eJqrtsqXu9MKiqSIDRFJOgjG6AzsRwrUp21XhracFrSmCCB81kQd/PR3SV+Vasx
rWoVk34RJQjSP/u4/lxjRqOWxMVzVDICKGh+LAMjrSDE81fbdTtBV6a0IEaaXYAy1dcS6Uv5ETym
0TTznuI9+Mxz+/QgjLMe5id54zCS8oxpwkQfVIz0AxCh4x22bOljtoGSCrRL5UJUJInhAMpLN3vl
VRks0WENNnoRXmPteufQS6ggDkzxbdSwjE2zpJTV5GBrgSbyssRumd4u/xyxuc/TusPLhlprCeIZ
+yyAuCTMQFwudCJBD7dye0xraw+npoPlp4KYoVjHAOjBgwOG+yFPIFQoMLh4VMaygU1MNx1CB4uz
2ooXmmzQMTm1aJ2g61ZcOrloP1odITiX93neqI+7JNv9eZubNT11ET51Wdz7IxOUou1b3GECSHGy
mrVlPgGyHj2EzogI0GKBRlZ7Qr/yKfBktMcLCwLTyt5dDrVbAol8esCy9DsrxigHSC3ALhE7eETM
+lk4CGYoJFoYeuncICP+6dZUYG+d4uiZgXeOMU8EGxF4R/vHVA7P4bq3W7FyzKw9gElcjCRETcVk
sZlAXxHfsXVZLZ7aRbHXRlsABe64jv3wyzIn6NM4HS+dlhhpBCDgyLx73oviZzveGOKZAoKMEUeQ
RpCDIVKIT4fm/TU3zlM423qzeRyr7x+qQ/gyJ52GFgKGMB8JtY5jQRW3OTELoDvKZnU3P7FUI8if
e9RcJ9Qz7VNs5Yk+chteSnvaYivXGyOZB8+j8JGqe1rGBMaA+s0PqiNYo0bKompz0av15lfO+q8x
ufX3whDFdAfM32+VcDKbodGCKgIDb3s73caJ0NK7NQNOlDujK2hBfDW2Li/7X7WCsv6OqyNAka5K
7lSfGM98PFcrN7/AzwzAQ4z2T23ABMF9UtCPjrQIn+m7OC3XaDUdzf0k1WajnPPklDUqGLWY7Wy4
F/usnwWScNCvFXNmkL5/R/yWxoqmTH+sjxCUC3A7hA6uymNNum9jjKUNxtF6lbFYDpCiD1doOW1A
SA0630jnwSHEDAahO0+Xfb0/6zSX6KVkeskipw8xl350h3Q9yA7hYvLIiJDr75Gmfrv0Hxk2U1Be
Jdnzx2sOl/YsUz4ySks24Txu2PzBSQ5clBzm13OifyXFCjTv6UzSsb81Pt9UZA/Kq0nbEpiruCTN
Y1gNAHfhebOTj2G//NmD8RydzjdMKA1hLBqVzKWsdVzi0IpMw67MkpN+fGadlZZFBfttIvnnk4gL
THrRLZnhcYQBTtIeFBjLWuiPAeA1EkfN3UbfTQz/efDdOq0z8YwlCYFLN6/vNpR8A5BPTovYd3Ng
3MVioPKUV5y0IVi8IjWOYeuV1r5SgIK46Xp0l9j4fpF1E7W4hbzc6vMPMwQAUB7RytY7oSfRkX2o
RdP4/rFeCQ8IiEdhOUZkIugt7YAhDg+WT4eb0e50NZR05fknBtmgDMn0wk78VlPfkoTLM18/TjCq
S8sqI+1TbMUv6h0+GSsZ7OLhi7tZBVIC/jitKt/C9mskgUh2m2vqkkr61z5OroYkFGcpOhmT+d9X
JIfwJJo2o3jDMgomFyGOJjlStbiP9PwvE7g5PBJLXAdOtcd+ClWXLcLocxoYHnUr+MgTL9OQT2R1
V1I2qSNhUZpYjSmnwU1Q1ooi1MYJejoPTu50AugvtpSUxcu244nhOvjXWXto99YDv2fWTaoshcmS
b000lMhyX4ANEz0lPCMD6ds6IOtJlhLmJFYSPVvbRIiCLu2XjXXvBRgW+DQryACH4OCrQjmjZLMx
D9NwercuGq21w8aUDfdd8BAKsNuXpzNZXmma1EiWuzeLDW8qbWYCbR0QLUempJCf+DX/ephjdueA
sUzTjOYFXFmAAd6OaucOea8OMXtwutt8KQo7EMJBkl0ElB6ha03Npo5mMwJ5chfQ1E5mBspiI8UE
Jdfwi4zP5nszloTt6a+5Edu+2GsbJ9VJzYA6iNRQE70L7vGamPX7OtF3FAyCkoEb/lU7hrySpEFH
ZH7DJbKCa4g3T095FxDLgBDDstSCs5hRjOz+QasNuASwkYMGMY6AfXBw9J2H/lIgJqLzdy//7DLx
bzQyhVrKHpQUjPEOTexE/Wp6Y8Fg1I2YfKQU2SclQ+K/6wExolWb0r/178e/9APpJ2FPeEmCQ6SU
WZnjjwFNZyDyvQVs4n4Xji0XvDFk6cDxsL4srsUGh5OgP8SGCA/asmPXpqls/PTx7VxATkNYN5RS
PZixJhhJ+4ANMfbzk7nCygV5jRdaQg4wlZADNqnOa7theYJw9PND8GnUeOOPAli2EShQqDMLxXyd
VWeKxZx6PLRgvTT7W8mXP2iscuZfEWvVCOy3iT1wTbg4RwApVx0sFcuJsPEDt5UNXFurNiOQ9/wS
GaZtIjJRch5YNuAzS8tdCHeWcAudj2O3QlLW/pssxU/J70lwI7VymSSgW978+MF6bodNrHex+tCa
VW7v1kdxDEhYL+yUlmAxISIMWGcjqFWh52uRM2vjYdDwE3tLH7OqoemoDhVTy7J/aj5qOQ5O9Bef
2AMntWS3L4P94toHZBFg41QdP5bwHTFiItOGzHNy3JxLmourmwmuvL2i7sUBPC9SzxPlXxJpb9r4
STRaFUbFybTR/I8qqvZT66y0URlqxXtcjnuFXVDm6eg8kDtgp7ScHNvOXlTXlw0A7K6in8xLWO2M
lTmEr0UcW1I4h1po7XurXM2SkdITiTB0wx5ofnZz7/oA7ZBpk3RtIeF7kiL0qU4a6CicVyw+74Bl
+hV1RwaucaqLV7fa9GMQbpfbixmtD+iLQ/PLt/5sbc0beoD7+zDzpkHbJ7awfZGhrea+/dvjNl6x
JDLIuO2AIVr9ob01NGSRIMpgsD+94HuFnwY8B5WF47CpxWHUJnYCArv+Grl7ffTsTJhE7pLlpfu0
eKEUYvZpL8ietYV9FgR5MomFvVJNlwOBeDguMTIMYnP/o8zhzWUUvwc7/t0Lkxik25WbhYm3fv7R
DOL1kLiWvqY8c1NxTcqXijWazoEGRhO2idRSalxN99LimrW3On+DlgAJR35FyUubmxAm9ivRBh8i
7RTRHnKPBpYN8Ow1dYtGJSfGf+fBOFioO9SoC1zP+N3CcUmDKFZaF9umgYscx3iD5xi7YSc23E87
8/CXn7qxFWkf9A69ECAWDsCQxe3+23dnFbll9Xdf1ijU8WJjLW6u7QgSYHqYec53OkzKAKpbtM+e
XTFDUV9VPP1xiLfwp162EpIdZh3XM/CL4QD2m6RxpSUcXK3PbaKJVmEzMk+Zd+97NXM0KpcHfbV8
0hnW5jsyRllWfivduI7n57S2k64E1Gka+Th/3so6uF58QZTEyNL+ktRrcMScaOUW7RC/fDgo94An
D+5yJa++FXNYVhx3FUXfhwtAFL+FIInrY/mdvau1LG0bPWBaqoLWxPzC23c6ysiMhmXfFRyWFCxT
xxFwakTDaZO+TweO+JUW8IGhHEAnAnOCWIsJ9dlRXKQgnsPQX4iUAJj1/7H4XxSuMGXOPsJa3O+E
7U78BgAdleyFOvSAiDbQWt2b+3FH0rURGkNIAu+w5VrbN4eqj05M/KxRDJsrJygTB2F2Ja3qk22v
9lrYJRb6W9g6bfgHzMwIzkwQZpHG5i9lDiupIlXfQzStbhniCt/IRMolB79/Z98K2SUjpn00jTb+
+jZHdY9Zy0lmjY39JwCqd9lxpBpAMi64/Gxx+WjJe3O6708KLh3Dxc3bdVtDIiMJtHIU5BxKuCMR
pvOl8Ulpn/mkTjK5BV20g4Ne/8MxyvKKO8HhM1BeMeK7HAjdoTYnGGmOfmOWHGVE3mJ3bVBjEgxg
VsiBJLDzB5gmqz7z0W/m1BsgvcrO/OVB0fGoXzFR0RWYQYn2gqGN9mwNwukwbYd8J7WPSKi8ifqe
+74EuLBnIuqidFWNsvKunwk/ugbWabV8NjVz38QHRgl7ORVOuntNVW/F4Ttbq6xxIXipS4VWDbLI
SFF8pR1TYl6Mx7JOlzGETmPqzgd4B7kRjFa43gnD5Npsp01c/dm2C8r2W8G/+DO6f/uM2NzFoLxY
C0zD4kYVqDNEnllWPQOyWFRfjspsgxfL9KfuuDOsUUmr+WDM2g5TvsmXRFUkE1mXb4QcZLS+5R63
AlRNULKKJ5+4CvaV14KzmZiCKDBJhhguzUWO6K4DoOkr6tHkz/14oeVcKRFt1M0WohZSZMfGuyO4
4NYsfnTFWOk1cBf7e0MYvZPgPvpi4Voe9zjRjITRv5VQEQHRxEJif352KvluYr3qpvXjvuOdXpYu
cMAoaxQx9XEC92HVQ8bFNf0icvHpuTTe9rtwUdYVVRNOFbEp/QxReHJt6zDcaC0W2Oyd7m3ZIJO8
Q2bZIFX6LihJwGzfWvur0tpBbqhkMb2ZXMS6O4qLiLl4+6olUmvaJiAYk0tz5W9pnWyTAUXFxIKe
/W/THpMMJpYRKyuevc0OVgP+nBW9BxZscPsqV0Dw3PWyqe8Ud2HBiFB8M32Il0LtxsG4xsFlTYPX
uJFgke5fa1xa4D6PqtYWrqh+jRk2aITG4LopEQx+EDis1RGDaE+Kn2MSrxSYCNMml/yl9MTkDZgH
OMwdf9i94ohFsyeU46I37N9ptXjiTSU4Pk5RFeSJFF//lPhNCThnDA9TNfNAs3S+D0KYDXOp37IS
u/UgVx/Tuz6sVssI6zu3XJ7qqAadrsRJHa0tASvm++3eUcH07sbCk/uRf9KVMDTWnOvAfIPCbGQH
zoPtuTaFDDN/H6muZy1K85qlGbgkb0EUEKvuvUBZJISTv6uszrg2bXKqbOSQKT6Ql5iNaCQd4WEF
/Bz0TY7ZKDhCXXZ53Ljx5B1qUfBOwCyClLzBYCbzD0whka+IFJ04tuYGpAwIlTBIMG344w1EXXcI
QSgt0h5snPsvaBKXlX1IlvB7Nl5k2HNnyL4LRuPoWpmcS0zA8FCn8POaxz1uJUSW9LYp7lNbcp6f
Nw361XQ3m8xjMTl9sz5E8Z9r728kagrP2YgkZg1a6T2SjJBFbEjUlwlFXQNXkhKpQ1Y9VrVxVxqW
tbRoph0Y8vuqm9qZx+jkrWWBGkABQgoCTO95U9KPzaSPSlJcz7d5lnjZOd9yUXKao4Hs8+aM5F8l
1N0WDcFdkN5sRKFWTDEETIaDE0Av6U/IYuP6iVExHnmXXDtAhRuQQxNl/+9yMgXJdZtN7htPaywc
r7H7i8GXleq5jCU421tFO8YE/JxkZJ8boCEm2od0f7+NRN8zmVrECHmtTScXfuRY+PEiLwpliSMg
UEr485VrUi9TE5HvkCDuektsPqkmPyTNYu+ElW4hMwYlsM0XYub/rtgECjprbooKkYaiakllHExL
2MiVpgdIfmkoqAOKWXTC64GEhj0OeOlerlQx5xhcayLDkrIRlWZEuc2FAR23k9kf8ScMPGsSknS7
bfAUoTGcjk651SfuJDEnLrfpPFNHnxOULdZNZ2DYa4Qacmc8y8GzA3dfSE/qooX7VlFqZicBXNai
0YBqszkDNtulgJoBXTtHJJVs+p+Y4U2UDnrL8jsmyPghnohAwDyVuxmF2guLQBauPkkC+Mb2/QUa
7DUX6gokOAq2sqbSJEzi44+pO8fyYlWGhYH5w0ybHcdrYi8vE2/HlzXjPRInCnlgnXFC6FzW7I22
2dDy+v3KTOW5PxkA8bw2DLpgkij42aa8Osh0pkkasdVh2/K+tM2ISbT4ucgXY70n2Oy8R8Y398dx
vgP5We8SdaZbCTxk4dWL5oMtBQBEmdHaKpuW0mTKCg0YbPZAucCkYivqG9qgzeqD0zzIKoK94rTP
YobE+6JbKFHcw2DXd4uuC0ktRfT8sdtsikfKZsSZajcFm4aW6Y1B2Rr9qGH2LXsbLr4WHC3j0I7O
Sx2H5jAP4TUN90FinujVLVxyMOmTOj56aIEVBijYtK+2yqEm7Wc6m+wnwtS73KlvQjT4wzFeE7uW
zzl65YglE/gay3lD7z6sGMk8SQ762UkaVjaI325VfPxEBhLoGYoXoPqBhIla7JWQ2Js+ru4TS8xl
Kp4RJiamcUIbW6CiHkfVYGeLTk0b8PeMXHzbxIVWYUIPagdW9n/r/dHzo6FaMxjg/iUhu2DvzaeP
Wk6N4xkycfGq87QfE6VYAAJ9ebJqb6lAFacvi69MrEagbLXp9ocleFSw8/1EETwwqawSvIsiWZGO
IMV00Q85Es259+qNED6etm3NkoKLAD1R4miE7qTna8zD+5jEW8qW9l7ZyX1cgpuFFB7pjvfVxzdO
lJxnaeIDMy1VkqIHbIBsQEHtUlkBueRgcIdrJMKP/SHKr/c8Ho3eDkkEc+7HLItyZ3EnVAC6nD4b
AJMZ4pTDck+aYoiU8D+Qn+G24LOtpyeHk6I95JXZEX8nq6eTP+45LYNOjPgOCbDWVNDdWKgzl0uH
PbOa0rsf/OYYaPODVl0PZi2CCqVpyaJyJ+uldFxU9eu+FrqM/4l7ylQXEfYCYZi3VqIMtTuTMh55
hPft7ajmgZm0F+yfZ6BBA4LOEsZ4ZWPHuLS9AWSwrc+qaysezeCEx8z5cb743RgyufNiujmv7jFC
tpMJ7epSeE4AHmMko9ekMnYu+txCalQhxEuN/eEAm45S5PjXk+wK0eVlgeqaWZ8Ykrw/EF2ZgsmF
C/eK57TUaZcb/eGrngy2XxkeRTjlOW0p1rskCzQEH/mgJh2zQFX7pXNOX6YvYLq/jv9Csa/E4T8P
3r20tLNAkLqtSWJ1ud6kO1f2FmD2Cl+aExRqAdo8ie5rxhj2tSKpuJLpXagDGrDY2bJXpP4zg+fO
F+CYusD0QJGRCQsUAnuNHOu44TXBE+OfYJ6QdgtN4XJgPvRMFpOjbYbO+Yg7kO7j0Hhx3VrBeB5b
rOzwr3Oq7auf5NmV2ZtzjEBof88d694eV2FtHurJhX5odbQ2eitaKyd7fVhY10EOpg3R8qdZH8X0
2gmFAiTNTtZqdYre0LElgjwanVU7gtf5P2/UOG7qXniXftbhLSrfoyKIazORtqelD/hjiIAQ7LJz
HwlO+HlqVkn2vohT2uovZEImR/OUWr09V3aB7SC8/UsZUPOyjqW+HiA2ZImN0Y6dEa/8loiAG5wZ
TqxGX8Q2jbfXss7XWI+9cpxLMaLYngewbZVTVhTKBjXGO4j6M2pWztUpQ+CDLGcc2VF1rBRNwuKl
KNpqry+imwSd3uda978eVmv2yLpH2D0C9I+PzpnCuxXOhRWmCi5cL7qI3nC0LBGcODtdSy9J4EPv
bvv0KE25bljFZvV3sbXtBHsqaL0cGUNKK1QnV7YuBl6DimJVn2xaCxOqOV0DCIG2Ocl8dTm+zEj+
MBCAc3NzEv1Hzjd9Rg9GL3elkCqjYdVHQCNIWd9cWhEeQ8WPkNbzuFjXorkpZu2kovTOC0E7YRRY
+/oQleBVEXXnCVwg8JKPKDx3DwDJZdkAZrdm/IWY6+Ilc4exqt1UQg9o7oR9ompVZYSXakKK6Snm
FmgxAFHGyuntRN1NGQzmY2kJ72R29fObuNONrjQMsDR1DR6hHTWOC/JH1/jbyCIz+eCrjElIteAU
7OttETOaL/hDn/88TYo0bq8g07wyp1N61VvIsnlNtodBOlUBBVXvhMoZo3Zf+IlxSa01GclYFePK
51367okr722swg1XhgYztlbpNzmv+hrHdDW+5kJzRp5/GHQQM9Qz+2ZcjWtCs4pa71rinqZGA4SL
k8Lu80e7+1EHIUTooQFpXH/0IEcznkBDa1v08f8rvWGEIdSn6YYo4/cotsKuqiz6sVh/F5XJuKmm
oJEyeVpYYhim0QuKUYj88COljQcnSXbUZv6Y8jJraY6kjYKXqX0yzHGfYu9e2ThMlVhNDAMqJRNW
6S6JxwNcA/K3MW7+pSAY7Qk9kAl3Ta2N6EFdmoXDOkA8scJfRpdL9srxy1mnTUmO3BAXmPtL+A19
DfUG5hXlMbYj57BD07vOqJlD+XSQm7xI0HSprQTEoVZLeXEHr2Un0U5+44iXnq2oxHWpc3D7Cv+Z
OSaxtbFYC6kTfMrda3weGU6+cHZMCDgA1OGwA91PP7qpceeFr1HzJqh+W6EhzIejuGcH41dFn8Ny
kp1M8g0xUM4fucQvSSiTXU91wtJb1rX9TuTjGS2TOSpPGmLNIl3WD3KFC/s66R5LOKo1PRd/NLoo
NGIQmsFwyLRw5p/TvKKcDuJspQXdx8uLKVIfKcD0An+PQUDUDgRQ/E3ZwtME5eCz4Wool5oPSAVc
RL1Cuee/Zt7v5H8bswfQgUkUGt1itKyQmofjCNePQNSeXTjKSmiEMCm/vZ09N+fLh3rgrP1ZOoSc
QaewFH9JR6f5AohHc9TaE5mWdFg4Dd63JMEWNMDXRUqqK6JERc9oioThiFKxyGRup/6l+HX5DZE5
Y2tC63XrdHdhbY/UAOQSIjkYZxVXKE88Tl4ikITAyS09cZUvuvcw2fmNX8caTCNFkksZrW4ymLFv
44dFZrDGNZ2cXvxVI9aUktbwSWxUAoegoK0gMWeAjdmA9z4E70ZCR4hwC0ox5X5xYrsEelVxzpY8
BBIV3+cCe+lQOzmOtAJc7H5sRWegH0pA36I6CDAMK4LsDQlHI8HlFMZ1TpZHduwkRv+fXD1SrZVO
2PqVA1knC1aE0hU/ojV2AbyynLKjZgf9jakn2x0vzcYLd1YiF+gU0SIRYS6f+glpxwDlaSFWZZNm
zI09qS7d/X7Mp4+XCI2t1Q0pTDvbYsQSrH0Oh5iLSdMIV7TYmXx7XPkNPPi3CDjyDUe3MeaaGt2i
WiGeO+H+Ks07qlUPbUr9loTzboV3I5w501rSKMULZMtTa83JnaPbSVWYqjqU8vMoqPaf9gLNct/l
a6Cg3e6MpbsC3jkJZR9raJx/fCb0TArR9h5QthkKihr+z/o71ZCSfJ+55afO6mD1YD8Ku+Sgfucj
4YiT0c/tx6tvWoWh/CEnWtC3evvP4MIkv22/jesx7XDqp47FX+zEbyHMdGNr590qzqMwEBEPJ4tJ
ebqon7e/Fm6mr3tjls3Sh3EcSXETfMGNa7njaZ6OgW54UNftf2Qg9k9+FH7Dg2gRR/WM4ZmAoyEi
lJ/Ki2BsxTaQvfBbrguIDQzOhrPwhFG9MwD371lnKpGQmj4/1XEmTkpVearVgp/FG5/u/4C1sqEV
WIWkkGNuILMTvT++z687B/WcnEZrdLMTgSa3V8DcEB/Ou4aNkdhwGWWj0XJ26vC+Fr71hR1aichJ
VYzMWXlTrZstDCb/ki0R6Ag9tqehjbyhFIkXeOtT6BH7W1IquOADk/vcyxDR0CYfa6iWtSvpX2lu
oe90wrlsq0bY8uXBafNekDfgYwTYH+iII5uCfieaIrDRHlWDG7OEdvDCXOGI0CN8eA4fFJx+ak61
7xu3vwi/gZE9r89usjh5TkyTL47GU9vPhxho2cgHq1szpd0Cd1SxjR2j8Zw18W36LAXpAHcPAzIR
8ckLDljOF4ouJ8vzzOkbd2J47ah385MPvsRa3efPOn2Yj+cQtOrAyucRn4etlePohDIn3CqcDD8O
kDpeuvCeXW1CUCCSRfn5LkB3OSdGisCNsEwiOVdAm7Rqmf/cA1Ja75XUpB0dbwO8ZulB93bKjGJb
yBkZ77zi2ieP6z4LIVEYfgigJ/tBJFlLggDHztn9KsMC0u+oYLZ1APST1K/dCDY9Ken0Xp4cf+wB
Q4RADnfyubOZlXTsGfKanJiSGfSnKIXeziJh2D9ib4B0XmGtfi6wzdTpLQq8d8WMn2b0nreSC6Gc
26t/XDiRxkHbHQt2SIfJsOl/OEOnTW+n7Zv+aFjLXOY19CkX8Xn7QuD52Z+AwwGBKLgSQPQN0Y+u
7RfATTpAqn4JVqsjPrnwoVk1bLWy0FXgBkJueNTUtKvKf6DhQXv/+RC8JxJskU7uZrf/cGh3AtDE
eB43bGfF/eyQy3BFr654qc+AonHd8kbJkmPlvece5aLhXxOZOxISUiRY99/qU4XXlS3dpOAytC0C
OVDEf5yLH7Ugcyue0obtp4OIpRVrJVGBfTfYT8t08cjo6DjD0wMeVBrQywsOt7l0AIBKoYa49CXC
05u+i2Yh4Z8iSUbUzwpkaQen/oktSXH9L24Gq+gymYsh+6OC8tiYQk9R9ylt1emqjt/+4eYxoCTu
+nWL0Y+0n/+G/ZXZ0n4CoowkSLzgZkzoURarf30tdTBRNzwndRgdQ3xMT/dCU7Q17xiNzOwbCigq
MwoM3AU12rWyp5GD86odRTj/qkd7B/y7/EdndfhA15QgxvQFombG2OmfGX1Wz3GuzN1vn5Azq7rN
wsLHpHBt/2+iochwrQFIKppGOzIXM4Jy+2h/MCXFPnGaKzoghcQWcZlWxom7rJ3kPj/jCtErWF3H
LJ1nUXT2LYSwdBhA30IVWzLrntQtS/tofusAQ6ykHFPyaouLbzq12lya69AcfGUKWI1Myd0bRd33
1+U/aTvy/onlVvYh0vNYotieFy80Ho+hD13Xm1wCWpiMSiBKZvmHS35Ki8m4KV9FuuUOPyJto3Gq
sGasgaQgBrydEWLqTxdetkKNapea/pEUWtp4HnkvnvwEzrTa7dyw2cyF/alB6+oCkL9uIrUknpzh
2gNGtUQOht/GxgRlBxVekwu0h1NDtcARbqmfkupZTy7w2WJih67775z8SRSDfHiQDE3FONiaf3R9
FdI6eq3Lq/412ooEMTKSVd6whoKHoDX0AS/jpszb0SBvTfSN+u3sbAsWFhRXkVhuJc7U6XVewuYG
mIqdqqDpLtKtdKfCdZGQ+ErIZScyOvSOlmACY/4rFd3qfxQbt36q6eeEM+IlpYkuE4vxnnT/2yxz
Mz2qLPGb4ZjFBWgtqcQ91PQc4jyLOnYyQ0E6RowYYDiINb1CE8oAZzeACESw7Qg12qSlrmPfCFfB
+cTvHKBTNDI0wrY5zPbA9Rp8Xt+c+vFiMub2vzGP11itxoKTQuTfU3HY/CX3qY+/pNMbZfO4ma1I
S3keuGvARPqPGr+S3rUYREwGbSfYK7LGSmyPWAvgZoJ/7STUv/a1qJpfl2zabRt6GAUaEHXvwn0X
S/uwR57BG4sy6pyGQ8ztsxZqAW0ruERdBGVUg24wSgQ/rq3mqNCKXJor7k1ba97iKNSPVYV+vrAO
TSsSfks+OrNqe0M0k9hdseAi7YGp1asRP95MOjUoauMke+gXrjMYiQjC3ay16iqX2q84jJNF5sCC
FTHADLxg7GezJgthdZsSpC7/Zfc8a0AkRvYGW/GVcvQeO/Mqvp6Hcdgy48QUyy5FL36YwVnOZDta
tHYQdDsGDc9qM07LnkdbzNArHnNZkiozey9sf8dyDn72SuuUvCUWq6SKgaoufBs/tLIetQpKuJVv
r9kLbZTE0JAD6VwT/yVBdlksC48USD4OE3eU+DNzMnUsIXM0bnqGigIT9t+ctb57PITfflAVyNh6
N/pU7KNWeVCo3ha3eFseg/1SLb9vOCHMqdUplHpvYKCiylgQksxiQiKempyH3H5PoDKlLih5Dnh3
efxAQmJR3f3EHuJ1dAKFSSIU+VtmZ+R56vOqhSj0eCKlFkCDEHAxb6HXwrB7+CBeDOSq/OGGwVj1
HcazJ0HEBJIVTIbXA62xd2wgq974EzIifnmL7I4kyhm2v6EJ4ev1BpqVXCvUyKUm8El/XPcISPaB
NZfUknffaP8BN/ZcztPhTT9ipaZpFRUS0y5S8ROjp9cXdWDxjlYFpS+AGk+s2dECLULV8Ba41N8w
9BmcKup3xZV2WwxqfjQBsliisPXSGU5kparWV4CTJHcWGTF3nsjSumVwRQSP/KaHGMy/SHwFB4VH
KOLElscgP5z1GuEN5oY8IQWaWHETzjymOnwvFeUvJAaguJlMUSPN1tFA+zzR6xQVU/Po7TljmuA2
1+aRcLHnwuuw3LfcOeEovl3OLDXb77UmP1YNx37SlMUZ3YJeWvakTCmFp9rqXySvxTt7JnEbDj2t
cxdYjx5ZwRaprb9Myc37CjgH6KD+x7lnzqXjBs3I1400l7ktRTo1Vre3RsIPmkSUJbOhBfv09Hr3
1LGK2Z48px5mkMJZF/LRDZXI+cVZlZ0md7OmMLkboCh2En086aV7w/tT9Zagt729Ud4CJ+0XIZvG
cLZKTDGQyVpZneddOmvmL3nM/MsBYvblAiOVkHTZv7vtW8W5zN8yJ764AaArew5w/e/1geip7kuO
w5404ky5QGpYGmRUrdxWP4oek3pu5oYbrsLdLl1r3lSMPKEcEGLO/PnKAb3Kb9rHuc4irEJ85Mgt
L8zTQQxITtKf+kZCAXdOttxknCNkh6tmc4LGvffeuqMBNHh5zUo3B80o1uAEbcftYl6cBbPENKyk
ZP61cPnwDp2rnz2oUXd1w/8zbsOxz24PoJ/dBDW5NlUOgwbtb99gvTuae0/rPX+PF8rhwnU2F7Wn
mY2p3rcgJE6vsL/3mIjKU4JNhZ6ND4akguO5LJxUW/MNQlbq9UOqHQpDvhawH8BANrZNZ8ANMoAP
m0yCF7MdXYwbaEsb7PjxEVHMruRezaGh0g0xNGtBwBoJD4T9znKTvMgo8CLjXJKPjP/3xbvXY8BE
Nv2bIj8zhaPD7iBPS/vSlykF9R0WRCt6c8e2AIrwE93MMqnDsd0UoE5WAYz0F29NXi1ZeJmzoh8n
73nWgs+VScdA//PoEHDLZZ7XPKA3AfrlQ5figaSlujp++awH2mIcMCXvy5Xdh1c7+5xK1kViNFFf
0TqlMmWjvrJtt5hxfAioCFrTBHQFkOa+vFOLbOcu6aB7uURAvnV5zuV2YaNlR/KbvS9THu7xFiw4
Ktilad7UlYnjMcLVq1w0kSrVIz8TjfIqT+YQ9s1/cpTwMmq5JB1wlZC0HLOObAENzNgUTajr9WhC
qVQhvI6znnBNtpg1F2lEETmVXmxTnivQXT0uhYoWKVLWwMS4IRqoU8zWjhhkw0udzm4zxRBYoabs
LSfJ2Z2wmuTyB+G7jGbdnnp+LCdG6UbCMhEOhhKdsDulwmMOjRL4pcnjJTv9LdZXkhUVC8fUH1XD
+y3QCpcrQc6fOL0gkw7qMSWuOVAz4NDGEFZEyTop2o2t67buyoB5+sPClDZDv45j/dxCVPbnIboa
KuEheujCo/eW4c/Op77lgXZGIU+l54wjusltHEnRbuEnbM1O3FnmMPGcCXxqsGsgLd/m84efV0lE
sWaCtZDEQsUJZUux9WvfJTUw+HIlI1tmNiwWTXzAiPEkzNYL2Zm4QeMXzQAKQPRj5fMDzd+levpc
P+p1x0x/haQl+LC48Og2zq+6xT7XLo5/aJ+7cr3/YW6KBXrINcokbb4UyJfpEhqqElHcDzCnNywm
lzObBIGaJsroGAz/lyRcQa5ay3SZW2WZ//UwoMfEOvDxFItsVnAl8IQK1hxrL9MCvT1/VwF5/2ih
QkoMsxOZKrtJI8b8ylZBKA18nOQwHyJLbx/pYO3Ps0kgIyOcLO/OsCkYxpJyD97X4oZqVSh0I5Uj
xUsywFQI4HnELKPWFND0qiOI8eq3SR10vpgiPxWACgAnEUW3NJAlyzYhOPoUuGfndjjtYL+TRvWE
rhxKfVEI35V2dBxql8sWnIPU20qkQ4r89Aa2+1+ysnRWJFy6lRdNDbsOIgS5IEMMT5GDQy89uBSg
4WmVGJk7ONKn7usZk+Rxxc9vS2YtVaSITmgSbnw/sVS7vhAhRmHUZCTkT/BJKj2IPbJVcauk/AC0
gS6EE/b7hoSniSOGL4xqJJ4+2L2KL4fcz4xeC07axPtp4omoI7ydfn43OlZy6yRQgBfiOhSSmA7a
ZC/G5rS5DgQLOzwmuWUvoxlAKq5bICSXXDwNugQp+XkIpPOF4o32TbbPygEgtQkAZg/Mk68dn785
/dwThh4vJOJZ0NXkxc503LyDoH1Kcbw1ZrFgVG7DeXQVTLW9N6xkiXooE++AgI6ScAho1FqZwpb4
hZI5ClHDUe9pggegSZi+JpVZ/VrY11uJIaaDQqWcVW1LUYRPmbE7HMEN2F3fa1NdFHUI0RYcoKxI
e+/ejIAj+E30eGJlsuwZ7eJRFMhFdFPs8hZWmsoVdIDyKACHCHFY6sL4P98rSS9dfK4xc7E15diq
3+rFBKnxCRv50hXhNAFGyne9xuREvcNHNh2cXJrD9AlmBHPClyGKxmgUThTWQiGk7+c2hsDZ6yaz
UuCyGM7yr/V2Nbh3xeBU8ULbz7KwJ1XEAv5aEGI65zgcJRuEXnP+Ialrpu22xt61i0K0Hlj2xWq/
1xyUWU6WFR6uje6a+MuTct0rHTy4E7hMnyaaxX90gyeAQaWpQY38wfUzGYOis2jNc6ECnhqeJFzV
4hGSJ/Hlx546kepahJc2QFhacAPqrlyeNi4Y6mwiMdC+buPiRa48fxKUr6v1B/PX2q7qTX42y2Cb
Psg+MFTJ86grLPKFFSFAbCJ1SQzooNx0jHTX0h2mXlKEBjhPDAuEj7TNIxumR9nSDeN8qCc+ipUk
FV6m3PFiA7QWz49B6RFrVcROnoFbVTHkA+zgW5yTfPs1Ir7qSyDxZWuu1FveFR3MGtqDiTLmE737
oFf2PcA7OW+hkRWZxawkPnW8RrOHMG9wtu/Qs9D0W23+KetOZeqHPRMW9cHmSyMulYUndmcsIi9g
I7bKDXgRglHbeGmbaetoU57J5P7bj88CfutLM35BW645r5qN4w3h0XEAAJCrKK5LmM0wLR3SnaL1
Fm0AbUo/QGeTcAf3Ihpnrp111LNUmFDK33t63KTlqp750RlkCcb472A57/SkvapjaG/RkXfl6hOh
ZKx/6EbjyytFugWE+xoNcVjbqHh5x099cFQwHpYwyUMiCb0hT1xCZJBguVHXe2QlffvBXVYIUtc3
hqw3M9CHD/lHV4C8JOFnV+v8kdJ7vj7a5qxKBx0dXo0BBUpu9/H6nsQXMqDcKv1ftTAkxQ4VIydm
bGWZ2rhfRe68JYFhSTiopc+GpBs+jvUuCb2Vex+FB/xkxzdcLu3JdLbhZenhrHj0d+kX4LKTckGS
tvWa6wk7NShZ4yRWmx0rz5MSniFETZschXCsGCyOTbK7s5FD1SD8i4E7eUZMazbH2Pbap8tTCtp0
4/aR9KXh3YUdXuKsCHJlSECxQ58/Soab9s/VwwQC7lHy3fr5KGXKKfT2QaUSWAzpiN58dLlDd5IN
8H2X/eoIjdUchaWOPV885E6nGtCCqHyit+TnwMReTTPwhK/tWcpsy8RGuP9MghfDKHJ3sKxC1Gs4
TG7WzyZplQI57ZoscHI4LlhCzpR2d2BvR31CM+dz7ArINqsoWvjrEv4zn7wHfT1EMsixi+u6IcP7
L+vvhh9m3ex09vJQPWOaybkKTUsPuTJfBlBeiMqvLCwLoSyZOCU6uvv6dbELdxuby9fKtePcy0ku
VX7lKreM86+9R0yMkBjp8DTjIVtqvosb3AZ4aw6Xq27ZV7m4qE2LJtOSpkDCrhQmlVlslxKF5vgG
I+Vgb+ORqW+CVLQ5rHDqMtmXZUsMpvYgNsc+zqh4h1dHhvAwC9X5xpkg6pJxhpkmTCGIToURP6j3
skM3Oshj1X+4DVq5Tk6Mcme7cZid2WZWTzkoQLj3axyXl4OPXGJ3Z1ZRRoXm5adaWdekC06dLK5z
gaj0OvgdavQBxF7bUbOVKqh818CjYdFJ5brpFviz+hydmxPvhU+vJGdtmIU5it9b8ySlR5/6W7TO
FMCOAb8Gl8+N/Ba2Xi8RiLOtNDeGlbSIw6vb2mU4BLr4gmmdMBlQ55UYwPaJ9/57EK0cDGdF1H4o
wWf9SZml3yHh0ddib0SdPZ2a7BvOsSUNeNv1oS1OqzZF9NnYUoPbRnnhBnBZHnOIUV3+LCrKtITg
s21MzZiD6ekk6kB622GlEfn6Ajr5DeBr+B8OvjGaiaHS2m19kGMcMQy31EVbH+yPkf0AXr7PEWdc
m433PPrn05GcHwh4XZ3DLTXdN9vrDNAdhTq2/cDmObZkiQp+m168DP/2sxGbDwqCH1vRvPtAKHab
87lOsHN70ZsfDn1cqHqLEsotP0rEge61zK3LxRdhhvhDBOXVvP5wsHuOtrMLbZYzBEiNWBiU6y8h
TrSXEkQAbUyAe6zgvq8h2A3ZlHKqMhxkR0LSog/SAPDuP/hdcelgydJxLh0UC7+YpkTfXbO8HCC4
JznygZgeI/4inkGRhNxf5FpqdDZzjDaura9zJffMAVpjVM5RUvfeXpIUWCYcfdKToIuE/l8USmmy
t6aufdnb2VGLkrbQyc6VgtjiXQI0Bb25h6CkMjIBB9zxCG8O8K07096Lc28qBUIPXmIb16ngbb7e
o82sCw9KS7maoO1RCrR2paIM8sXTykkNU+G++BVVxg/HGDaO8rsCTfIa2ZtVPQStRxAQ1Mg1aKYQ
y7zfhdQke55EpC35Gv1jmANIJ4/lMtdDFxCBEEaF/I3GcEDm7CeaXyMBZ/ItEfrN1EGYYhX9KUng
63nfoFpiXExlP3RTyEf+d70PEftcZNHGKwAHRp+DgjddDISe5cxfjCYUWOakla9YLxxF5Qcyjbrr
tNANHFt5fxzNTUmttkjzFUHwIEXQh3v7fbbjeeMw3pAhIcGnP0FpaL2j1sw1IvnVhQzNFh/+Xlwh
1z/7zmHmC3F3vcguaJsldKJIB2lLjmaRl2YZJy1fSUoPPPfLCT9rV1FGqEJXv5ezPUYvpaGrVQCI
HjBmLLRFxD24VeRWgD1MllY0xARvVqqJSRZG7/6RziTfix6MelVRlU3C/gFicFzzFG/b9cvkvbRP
0Cp+y7Z0sqxR79i1eqzoCU16rGpQSVV37ZEvm7P6jHcLw+67rXpYc6vz+sZWLg4bSWEEmjydlLrc
z1aLXgKWaVjTHyFiBGkHMnodbfsGtvMtcV0/2fHbCXU7TSLGgSkBcKneyieC9twXyO8LG+IAUwey
87rJnycUytYO/QhAxCUtqJNB6BB+xpMFAEdsTQK3yelPuZc9GeztbxZZ5b3fDIxjiImr5FojOyr6
y3XGZoPIL6QHeUDV8Z4Rb4TMEuVI9BAcxKgcH7srMhw/0mjT5qxdHae3xcMichhLKPo+io2Iual8
ylU+wA9ZvH70k9tjlib6Upb544AeRaK/aWz7p0nrpwASs+nFPaPHmkD3ypagf3kIW6HQGNteP2Wp
ZhWPJhYL67V7SMq7pi4coT+MlyxjlpzJQZjsrAJ5zmNIuQCTS+RZAA/ojcGj957X+B/ykLqp7T4x
LqsMkHttJAHnU9BEcnAhKzHrAFwMMw8rFJslA6VsQ96NbhmlWPGzKfIeyC/qvjL4y4ucoeMDh/jR
Aj/VkuqeFb/uHcL0onII0I7zYMPUPHvSnlmLyCerEd9vRxnWPZqPlXUC49Hsthc5+TduKcNdlt7k
+1++bClaNMBIkPlbAUFkM547goNOkrnt/DPUL6BqNNHizG+9SDbuqPL9VpDNj/NL+F42Xa74ipVN
tP13KlsKW3J0P8DxJJlQk6YLATA2xtreOHqTTUDXGtL7KA80yqVovnvPIc3Gk04tVrlRfhkym3+5
4sYUemHBNxkztcWFnrMQaiCkSzA3/JPs/ml6xgujLQbXXq23ILT6PxCdwLe4Gzl/t4YXk38uL8q1
AkxbWoO12x+wAFU602AMmACoRcvv1ElcLqPDUrSjyQFlMknI1b9w24EmdpE+W1ZAedb//bdgY+D0
1rfCfdWQQad8W5AmduZSAVajCA5s8qMpqjHVXDEj6R4O0pRW+eiWz2zJfbT6WOxYK7t3mTMGUHnv
Mmv8TTFIiFKAZDLnIaKd7IakJTlU9XW4zmm0yvpZeeIUyPv1QoxF4WDSRvupLEk0Ico1xKNMws/i
kW5SL4KGB8CAvzKK4gUUMc21DBmSIF0Koit6/IC3QNax2zR6exY5pw/wZKOX/Q4GnucPgH4RtMvi
k9qzadxqyWgMxFpXbZMcHIglZVMh+16LJXYtnqzHFuUy5Ei9/hNSItO+FyXIFEYI9Wf4KtXH3kJ2
2zGRwpEx8wRTtjptWkhviPkU5wknJbkVLZYD8Z2TnRmRCaOQAHmGAcb0En4iKf7cWxjhPhb8tJ2A
/UF+AOsEgWfj/W81FWWWLBc4kr9Qmd9ltzbJxZPIra0S6BPllfX/MtSnS3TP1FoDZNRp5oy8hEac
rqz7UQD6V1sbD6RqdiEZPXKRpYxuac+1k6gVV6uK5dwR9I4XDynV/vTrXduYqPCcsFaV7Ql2H6TQ
A85b8dPm87E7+CZ+4A63ye21jebqZCI7j9UvEFvFVcSaJSfj0rUmLgfhno6xZm8Q5UOGDg4EiRzS
GU9dNiCe8RNgh+sZvn1WTgbr39a00CTCKZ9XSMd4iRQADgIz8BjmJ6TeI6uIS2kZVvLuy0s+foeE
7/MpndQwW0BpiAFM788lETk7rCBGNOdM8URNSkSJmmURy9EnUpBnk+5ZQ8tQLi6WvOtJFm6TIjvu
FVeiS0MX23CNr3PCLxoP9mvxQM4Lo4a7Lco0rvsU5VxWNy638tZbknp8IpRaJoaCJ/vfoNMzVOz0
ip2wV7/eGQsuh/+/7PSB0iUtpDZ1RJyvgN0M3l3DhthXHQRhe4m3B7dyTO3ScmGEN1w7Dw2aN98l
oVhzojSWpgpw7rgexVW1tLt7mFMElA73hu5HlN7CO10KWPoDJpkvcl1/TAbxV+JZj9elXdCQpAMe
UXky68+NH53vPyEFyuEANfmAHz60irAVqi2D79pqeUDTkW2Aauk4/tRd93+sZJi1FwF4MuirpFpw
TGRJxTvgcWR5YurR5e8vPGrGQdBt3t5B+GcufyQVqMV8q/P4sL953KtJ0XIWwBFBu/KcVWaMIQc9
gaB1h4hfOpfqPJV7Zeif+M24D/4eHNaY4qjohCQ3tXFU+7WFTZzZMjS9yhe/8YKEnQnMF7Z8Hq5u
kr8I6vGvLezF4d9Q3SuFaEtYTwsfRa835nZnGxHtR6140ro4Cr/tg1JyBcZQk5WqVbmZBBmUfHSk
aZ++Rp1Z5+am9MqjIDTdyie7EtoXaOjKeKYrDA1zkLHtMLnO1TgCxfk3a29D6md+st/rX0afoGHz
hk8hJ8mrQtEQ7lr1a1kyRyWQJI9vgOkEpcIIgvQznki5j4gmfSDqtPWxlRydmu7wC9CctQ9/+pW/
OxH3gDqFszbhgusWUv45bAvuh5BbCrLLDqSQJRpHZ6e95oGB+FRXa8DHtXHOqw+spCCgsyxfW+5e
QiSjO5Ll+Y0ZjlW9R0x+d2L8vEAJvAW1au9FiVBo8ECHvUooDyBaHimEzeujiz1N75ZyVTIn7Wst
DJWQH1oyjznLx5Ky4joGFyYm/GeG4UwFgHyiYulyXSsp1ckcZjFCbsPbzoXc1ePO4X0BpCLoqwz4
6cxO3v7iU/DODDMIa8HkCwf6U00KYSUinSFOtcXf0ln9bbOpSaV5sRu8G1B4eh/WdAbO12vt6Qex
JBGfjG+XUzPGRD2UPiGF7E1Lrg7uuv1HcqZVK3Zm4LPG0QgTHqnsSyW210kLqoig/gUATuD/LF5/
JdsjzvWxG8oc8ix8ouVYBghMdi3YR1wzHiNOHAH6uc4hpApCge0j2rITD953ZIkTh+pg3/Y3wioz
+PXy7KTQ2IKS8nGkhI6+F52hbxiBEMYnDcTfpc7Ib5aC+TxzYQd4/4FVA8cvb7MCAf8MRy63YsNz
/VcitcmM8A7Wlc/ZNwWu2vnSl80Xx7zmduLZH1+LZoLp3vjv0cgSHuzuscaxwjvNPzGdReVtvYOo
KHifLRj02S4AUwvxNQZQo3HhbF1BjDDni9cotgeF+mBdjnJmfsmkZg9VQbVJDLTctB1NGVM5y0/y
BybvEJKoM3CNNtRv/ePgmF3zIpwBiQ758n/wWGMwAasI6e4AjN9+TgFLmwza0m5qxZt3dWnMykU0
S439hCsb65YY0wMFOZV2HSmnD0gtoRFzvFP/BDdxbshd4OyMMGDv8CuUCLz3st3ML3KyWMpPazxq
fXeK1d+Yr1LN1kFBMzVWQFtpjjM1y+2MfuxHUYhXg5fikCxUqjTbCeid3A74vrFjdmcdK81SU3Bx
mVPAu0uyYgYVVTLpu5hD5DPM0eGx5Z9QZzT5hAI6nRLzYKH7lCGcwE57UWRRSxU+kMh85ATnp+UI
1Qcb9wh0sksHtO6b5fQ3rfb2s5xHWKhioWLlzK/blyuzeXd6DDB2tKNO7Xu1CSLyaIKFY2GTdqJf
FR1gh38gouAkivijRmaQGWAN4thXol7pJFu0V/yeHXl2k5CPved8Bzl3Qr3ywuCI/bo9YYkThhe0
gFCCnx/rfuZjOjE/b3I9T6XD/+E/1ccdhTPAGMLeTaLWk6Xjp+Q1L8D6IagNTjY7OFGdiADDSthd
7338ohuRqm/TlQ6MXXywzhdbIyZED7p+iAmaO3HFgLf4RUnapNgVEn9KGdV9/79d4I1LNgGRAveu
1XKUolCEKY1AL+S1kUWul+D6ybEAZ3a3cMdQA3AswZUV2/TIAB7EIUdSL0JRmnyr4kAKWvx83W7a
MNnhxElYc87R4WKKkC+xXhAu8EjY6DrpXKtcNhODna1/W/vilaoJFUPlHOyQUUmgoH4Loljy40hL
0yIRjup7CK+q+yJhLnxl5PoXW2CV/70Jhymsm5G4IHlXeczSh/EqErsW3taK0A/zBtpW4S9jeQxy
gsraM5M4YdNuBDNELvVte6g9EaRhPMutTLDgMc+d8gl5UoAdY67RoczOrHxLsNl7kMWTyY9Dmap8
6s8NNVQkxEqgSNz+9H96AaQGT11M90fjUcoEa2gfgDJkjHOIVTi8rEPuvBrsWpu8dvv40LbifTGg
OqxghUClTkxSYcUKU6Oscf82uXrUa139QMLnSGkjenHfuMQCcsCUtCL/NiPuf6rWCsK9TbN8X+8V
In2bnleReaGy7Osl+GSV7tac66M3NNRYR+DPBMfYsSeJ8nPf18OHDxs4CAuGJejyN3FBQrI1CGbP
dQ4hVPzZRmEgfDpZZBkZolKSHsAN+56aAEPR72wQqiDfv/yyJ8jePa6TyuCBOpvqUFv3SJOnf9DX
xVvvSJ9bEU/Igb/XRVd4UeyhyRxJetMSfMHSJLmGbsGfolGYzYhuP62qTDF2NlH0ccF/YmevPJuK
/q9TmPw9pIM5jRqvtNOCocVsB7gpOatfiYeGeMb7hwxhNBkAX5e00t1DZyDXGO9RzHeRb5kycjAt
99TeYu29S4XnSNUJFB2m9QNcFjzRMZKOBPaz07Abd4y3BwRNWLS5SFAml754iH66q5QBshzCgpDN
tc/heW8wP0hwvIo5m3NyMUnSmLA/9PXwY+4xMeRPgF6RaBflNDFwOIwf7QM41cejuv5Nleb1UzZ/
SYE5tw5GCEZX/Kw2nRQRvm/H8AXjIm5n2LmaZ5SpD81B2niTp58esyLkNbEhohdcugZbbW7KZJkG
b2Pimx86BTVmLYyIM6EdbqSBDvSS8ld6QbyzXa4ephyZ09GBbfJdb1QlNSB8FZmOfBcvNOn9KPbZ
7yyJgnj+z8RDPj8P/CzLJoynI+x2MZ6ku9EZn9IdScknt++f+Uori+FZZEhtd6REh0tahaKFyp23
ipTk0HjDP53oqLdVfKREGPKT1Q+EuB47Vc/VUx4uK6bD9ncggvioY7VaQJEou7G6c5DKmNT6qWv+
hjfJ96wAYsz3M+uy2A7PHrkcgJmwNgMqar9tWoCR7oimWNjnyOg29SLceekkL0wnOfOEWCQMmekJ
Ney2B/i4QHtmYSVgMQJijvs9eIVqK7g+NkUhhjMn9sm9sa+y1hmu1ja+kuWgpF5Lyux6Jx26QwZQ
H/Ts8p0HDMIU4cAqXGZm2F6ozo2z28DWWJnlz89RJulvSHiDLvOF8M6jo5jlt1XW6axuNHAf5do3
FUfpKrrDDejSienR/b/OTQqRYVmz8H12mALxHsdmSyBDvjGDYScX9Rv76Di/4fkuqH9RFi2nWxHI
9Ut4tjtYsvS2EInXLxUQ9c9NCFYEBzBXMaMJBTNiv1sfeFKKqJjYFNVg07sLusZPnSoCuPF6hQIA
Gj/Sw8cKKf3e0jqT+ocCk/iyPpE07bLNo5QK1WTTV18AVZt++ywwqd1jYSWLnsitP4yfSTEU8j+X
kJKsi74cpfYzk8M4cMl7roV7QNPgMH/UARkgyreH75eBqmUh6iYAs42DDjIiiRsfiTv9mL2huR44
+6jNGxlQZW8je7YK915Lv9Z8ryENtiY0knZ8NMYvuwxL882mkCn7q2qAkAyfKqnVoRhhjwE1fFMe
NwtuW0YO9AYyEnrKijXFvOvKCo0scEx9Ltc3jWC6T7uPl9MKNt0Mm0lR5qQty3+mNG1LQu8N0QG0
JTFkZaYq+G2AncqTmBvFWhz0jLVtBJvLKv+Q2hZECFFonSGbXemjoJnTEpNRorMp2rBcseE6ddxG
NeYFTX3TI+LXHo9BFTymBEjnT+NbELNS/hu4U/6NowNpyDZaqyOMssiraJOO93ttP6FJQDiLYcha
6Rn29RXGwCEuBpuFRnevsuLSxSvQelgl7EB15ko7mcFbb0xcwiJawlZrS7UtZCLXb2bW4yTEG8b7
IFW/edCnQISrydVkV7ZBGlJWNFAO8C4huqC2PFaF7WWDG/5jRn2XcXQTVGgOZ7rHGFRGVnoYzE5O
mTSIIXzirxk8GOfXszuscuFsymSx9YrkSebNUzXVOsoCzdWSvbmX1Gv+6bgrourM3ayNPsl7nI1f
mfCI89BX9akqwieNLqpKA80231tla1w1pdFnBcpLXeE3rVBpIMCILbOu6BGxcEtNTBqmyjLDs5Lx
xrQ4lpAH5NkWyo4eEixHxbwSD9NHjPphkQeQeHr2kktNfN8qgQaihi0ZtM9bz+uGLgu3fWjnE7xK
3hoKFtGYPs/MPJwFAFu7PdqpmiWST0mHnZHtbp45o75DIjYBzcaGTEUMHefSDwrEeFNrhNtsJNd8
/zKfymBUmz8I/nMVlaG8FsUmEsOE81sZ4pEps+89QataZiseotJf+dx8ZIKWQ0Fq+ejPlThaTZdZ
pAadjvXPeni1v5LtrsWjWpDErwnwztTlMoTKdZs/wmLwxt5oF6EeamFtV6M7JVM2rP/YmwhlH6mU
Yfl3IWZ8HoQzKf/C1SRZVmqk2wcp2y3q0E0Heufn65X1b6f+iewZn7fPatLe55NNY6JPsVkCxk5T
cq7FerzTv/qycFvNX8fLSjUCiFChMzP4R2BYUX0222N/Cx0Or7Ara/HISzF8pamBqPMAejixnzBt
qCZG3FNyStmgxf+Ft4y+WQiZVvE0+xWp8jzlmIedXdD4DX3wyZELx77c8+UcsMMBiOJb//uTps4J
6VnQdIJCBVjjIOUkfxI/w5Q83WXtvsOa7w17ehG4WMYFYcyZINSJJZSb2+EMIIkYV5Vge/FQM/XJ
QzzJboK1U+P+VySES2dZaGOlEEWdX/Qiv5OzJb1ypDIVcwU6NHV1CWxzVVz0iH4j42SoxIOvOXcn
E1TkSkhPklJtQrPP0I/Ne+aKu8mPL+Y7fDEjIOF7RsubxTPoqMcIPzJ0A37DEqTYvvZALBauKVZr
+OWEcL/PBheKvh+15SzPDsasSSdA8e6/IbkTl7NgdlGXAInv3cLNrWEyzFZhIW6CtT4+YFVA+EcX
O9rA1fV2OCJjeEyARYClA9jy4CCthUF3M5IgYHXOq3EJQo9PbHFLbtngiJtgAZ8yKVWfGr7GZJry
N66NXi0HL1rY4PxFOfXG3OuSgRc3yy/A5MhGfLqZt7Ofao93vVpZPGlRpfIQBIf2xLGP2O69F+pL
jnkWP0fQkuj4d9yreHFeDaZPIegoDG3Wa9ZiKUBpgUhU99hHm2DgSN37hGrpjIHVq+vJeUE29LEo
u0yz4nkEu+OiEpVZH44B6ejkwOA7wlEk/2OdBBSbPuDXN7jGdb8WIVnWNMIYmX8EhKyi3rZqN+MU
SOPEL8Tr2s7j/+yeEIAeqtHQThHnmLVWJb6E/zXZynQSvFEPDRXPG4E76nvHOpK/J+GGpCQPPntO
rfBaDEqhUlTxtM6nwdhq22lgXZYGUh0wehXrVTbArF/9HKtAg1rs1dmM1GTW8VnAzse/kg8HiI6N
2xRT8QTJVsRPYg1hJAhf8I3fo/0oOwase5eaDotvOqt/012pvYftIWiUCtUwhjOndtkwBUKjbD0s
eBaLDXbFYA/QmxjZmmWmKsiUY95Ha4FgzB/qaQQHBXztxR1YjXvHxytiG1CZVt1aKKhC6bz+tko1
1RmbMz2PafIm3d4wQqLP5fmjRiJzMnHn6NoTO2zs+H73Cu0J1LZUWx/ft+5cZm99uo4tvudHKCmF
FWVZVyzpwkLGXBzwgprWpkWjEg/Q83axUzm5aaSBI5dQz9AmslvF2PZ0aMETXhjNyUpL3d5A0Ii2
7+BrCge2fdIL6oj/8129y9M6XbKwtiHWypaP3vHIKRAF85WeRccd87RJBAg3pgWk3Tac8U0NCBm1
5PPaCZXTOmYO+NGhpMfXTLzjgsRiXUmIWl54DVvC8vBn4GVvZOrrlUDEHC3++z7NvmITld1xsX2J
QWzCWJ7NN3JxKhPr17cBmt2NJ81cd0rZARCNaXKEAlNw4AlYGLZTZzkupyNTeoVCqCMYe8TpNAx2
tydaEEHhlL4QTRPH4PURNUOfLwCkSFiYhxp89FN1K7925f437xCSbxBeJMBRm8HtTp+FIpDGeu/Q
Lh2ylTLDMDmJMF4ObDgmRs2uW8srQa+kvFk1qgqOuCfQL6gFGU8+MtfwTo1lqVYT+GA2+hYrMgxe
vP3c8NJBADPLudCWNJHpfI9gyxuICFfkVwoiso4Od18nlHLuOECw4GPFolNk+SE4SXErGMHdZAYv
fcDli0aT5pLHr09VJKKICNFTEY3/uMt01oMjd5b5NMlAFiqm/InxGUhokYhMG0yZwK5Oz+djleHl
jBVVYdXDVFaHHy8CuKqQuawPcBrG6uPbNLGD0TDpjeATfVdpyATp6aqCMli7TTZrSnGYdynLo3od
7IgUTVoWu31p0HfMWJDMgAb4xGTfnQO+ptP2AwFF2MW3GWYFxHyBv4bPKRk/tVBkxIdR2bWbnZK/
a2cyipChASGnp99nlwSBtDGiER4k86i5KYyynEptpBaf3KwlcHeLHkn9P20FCV+wIEN556w5yTaR
OxSjMLT1UC+NHaqDncqqTBiibf48ar2Bvr7ZmDFRcF7jwdl4I4L2MXu+U0zRGVPSC8vdg+jAs7eC
3egd8+rMCzHAh78KW/+5XODRFavCUpSmTLvH35yKA6MkRzShEds0PkkT4LBQcVDrlsAEIcnrqWoz
GgQcIx6XQaoLIX/3KUIDr2TsHf2HukDQPU8ZBqCNAvd13DHwRHPJVJUw88cR1mGXbpjex0H1t1t+
NYYc8j3ixCfhS8bp357dNMnggyeWHwKDZcX1Bw/GqGoyUmBMvX/AgCqOlRSmOuutxSUVKlGUdWO2
b0eroApUM3URnVl93MqoZx4ZONNreMEdVEyL9eWW14+awMxtHnO6bo7/CRVbsnbWmVX8w5jHHptP
gzEWIfZmzcRQronXOtZI32NcDw4PIYl3J4pemR1+WkQmMu2buVrismL0GcfGCoCWxEEwqh3HjWEQ
zGDAwbuuku7S3/5VVMNCm61042NHc3paYBBTAmnLTql3UNtIp3bIVw3MPEd/PMCNq8xK9xejYrvs
maccCT3eWTSeHF7t97PuyHRt7xexJmeqiPuNGvmVbp9cIuuCRCBwlDqfkNNeFP9z0JA+a7s3mbPb
ip+DygBc6a/5V2IczOgdkYilIDwwJseQ9IOcPt+UY0649bjlKlk6aTLuGdBJA5vrBCJSYK+RO71d
XtkAOxlltAGFA0xP+n1JEKtZRftlKYsC845a7kIBiGssCEjtJnsOw+7a/XMJQdKmF6abJp5mbm0p
fSEtSObu7WZ8cRLMPJOKEyC7dCS2nqmUDhkndxk1Y8VBB+Id6xcRjJPbCaa6YOAMuEu2uDAcr00b
ATXbV6TI2PqsxESxBO4/d8U2X/9d1zSthsFSuENNUdj0tbiiEOGXG7Eo6Dv44vn4/C6NRdd3o2uc
PAnDNM1Yt/QjdJBS24uWyaEf5jCeVGvXzkc34Cy+fvZ0yle9hodVq0+lUmJtQAzGrCXOJa8KGp2r
wyCls0yxi1kNN8OLEXCQeaamtge1qimWlKh8Dzgh6tT5GoX4FqNcl1KNJVxDbWFL+8Kzxm6/M2dU
k0iTcMznuDpvQuywxMvVZXD0fj1aFZslzZltyh0j4dritwFtafi6zRyqimpyx5uLtbvp2q9kbPAT
Q+Q11PMi/JG64S2aROZCsFa2/QVgxebNE2U+s/QGCLkGkMFqETgW5aKFlBBvrpo6VPEaWMbmCCtd
5ioEv+3RvMUM8hAdv7umqALKR7uIiefJM/HNBW9soC1U6CVTYloZsMwKT30dzeKjjHVfFbp1015x
bGXA5KZ+aDwjSFaVXygjU/9uuEj7ypPnOxa7tX+nDNczXqh48WrE0YlPxJ1kfQSVN71SIdW1VVXD
GUO4/4RUJ1ywZL/CWw0DJtUvjIVF26bHlFMf8zhtMq8MqEDynv4MqsIsUEI7MdjJfA8mrmFzS75P
PqSuQK9G1jau0ZtXYxb1Ht346pRdL/pHqdvHaS0U9t8eaQ7tZf5gbHHwi7o1JuRFn42IPI7JO2IP
IcH32JCbxCAjqs0x8YCE8a4z0b7pSZhYhDYPJkNJR5RYZ1B/X5CxaJhkT7HtGChcBZTNzADmDlC0
VJDs5WnXWtf535k72lQRlRiFgVqBYyMmFqdevzq39mpw631ZrzSrho50GKP39vOgcQRw57sWl2V7
+4ven4JrxdcUiFVWbItSy8j9zNuyHq2nFh9+Jk/Vclurg1zt2npiPPU5Yy66ITsG9lWjrLZm3c2W
LQ8L84aPjR2dNd2tRrIKmvYXTUspQhq3EWzlgIJg4WPYtyLcLrsY8AZLs9VZJBgCcawaOKFRd++j
g+5jEEKhahCzYMZFNY0rqnQJRLoSgPIT1NmLQOezxIiX+8aQoa94i21DDB9mPdjmHJMJZnW8QLdx
d96IikmjdVuTU6krPviCYAIj6OTyzcHpZ/OkccVQEtuvrSprIqStXzHviH93nmftk2kcJf+astRR
PHaMYw1l8Fwv17NibALxSeluSDx4VjM6uFaurbnZFKvo+F7KKWHlTmo2aPTViy7bl+Aisc7Khf4j
y4+zoLEk4tslGaalhQUp+wb6JPr3PLGbumAfZSQVqvb7mk2gNjI6HlodQqlGiDfoLw16RQeuxlPx
dUzfhaTOkkQMvfqL7J2XOWQ0FZoHibNFzeAsndO9GbKGdaqHmqJaXAkpFrBeE4iYmki6F7DzIcuZ
KfuH/jMKeYt0YHbeu6ezmnwJkwPqPgsNM1UIW9aqjrrLEt4t5pAsU4vjN8hc0pd3oqzN4c3wJMYX
z927jXdX5fnkfMKBWYl/0ZctZ6i/XeyxUD/5v/8yjT5SNb826LhLbjtGs32Y3/dGjrMt6yhUAXEo
NfJKdvSoY12jkTopL/E+drVL4RbpqSiihdN6Bhw+MNRwEomrMzY2OPWc+Tp4L4LmpevX2SM4q3Zp
6J4pWiVML9NIY6E1A9q4oy8bIGQFI2bFowUQuz6XRQDC8VhgZ/Pvtc7DgbSdcyPDXPsu1DrMeD2P
HRrhrNxYQz0XLFTTAUXN1STx246D6H5P3Kxc0efuCTHi5YZpHusS1vou6StqbP5IITTQAs/tLNY3
G/seQyfBAsYgUwbYJ5/QOEnnmoTZuam43tNjSbxsJ3qh7GDUupoLeI7R+dcSSsN/ioBccqWbC70h
/1r3QfcqSoJ5ocIiA0rMcABmtdcOkIuUAn36ro4+4NS3ET6QY/p/zL/GkN/N0ti3F9P8DXc8N88h
cufTLqGfNZeJxmhlnkbXInc8Q9u7o2Nzds73vDOevsoSA9k6h0r1pGVuDGPHlJfgaNzFGs1vobY+
1GZnukoFvuDZ/7vPP6tQ7VV7nrxe7GaYscVPxeLqk/JmWRJkmsa/baDVocoMFZMbRhSygZYEzSIf
3FYomv0QzLQPhbf2Q6oc8SgLhaxR+1jR/HlLjCxr5bLyWU+Wi+ADfsVFJWHt9qRnj8QMAKhtITZJ
gVP2oB3cyCehpUElDa3BZPmwqZKwjOSOue7cxUU0ljVRdUewFeHqcFyVH9Zx43Bi3QBMkCfkJ+18
9iHUKv8OBhP5w++4/7qL2GvJ7Kqb8jtGAtQldePEw6XsTxLwb3nt00i+YgK34TLPe9O0BvLvCiOm
TMLhT1o6bGTSCiDjvyAz44Qmd4TIU45Hk/B2QeDcNGGGFCixRPRiHIcGVuinyHqh4SETwRAM7MRI
3OPTQDkNJXS+6t2aPthisPaTxAjeU11iBd2iRikXglcr4LnY2JAoXD+iKRLo2SVba2mGt8v7uW1J
rbzOwLhnwIl/6lGH3LICZjex6JNdcFCSao83AcyhCwb62PQCTAkDtfSANlSsM3HTdLcYzlD8awpf
j0X9NdaSgU2Mpq9ON8kVI94PkiKVOTTv27040/S39E/eWmog/ghUn3h1+/dXZZIHR3t5UuvrXmqS
JVavRX5ScfP+JUWi0WH5yP+SZX+nkjdDtafi1YJfpiGrFZl1Cg8F5y7QwRqyXhydjWY2GuZRNowO
oet1Nd8+dYN5Jv1p30ItwA/iPZdD0aTQ+RSuvLyqMfQl+ClwfE/KR9ZT8LhEvTsU9iREOBIDVvhw
ERWUd+QBxbDlEfTL8RkxjX6jp1FeUyfswJ7ZXjnJFm3Kxu9888gWpCKLlgoV2Xf0p32fRDUUqlpM
FDb3mdI69eVtodAH29W+b49bIMU6msmsjKdr5opUiEW9zutX95TPGPhugg32OVWZbY5RYZ5O3f4T
48IASDjoj9Ft1f3A8ynXKmFOBdgToupEup9+K57ezMUqyxk2CQBXuBrLreyTMj+11ZTwgamdo6u/
r1eFbsT4l1fZfNOvwLnGvMSswp7TX8cg0NvlzFrjrrChBMd7FT/X31iUySDuw2h6Kw8Z71NOOle/
3UYzm1buJxMFMNez3/uBT4hgvH2cEbtL1NMZyO3Qigi6HS18YrE1UpCQW1Id6DUfvjqqpX1g+165
R7IdnCLw4FRd/zqop5/9+xN/9umHDhqd6/SWfjaOUFdR4OVMxTMN2W3f+PBvf/c22m8bD+0Lpac8
zxDmqQBrDFThTutPUoAyABtxeakRYuwsgVG/Np87gsY0UNpVxB6UuG9cEPBTV1CCzKx+Uz2rAmnx
oM28pVPAQWawTlOa1hRFvv8EBl7GWNczgCZoKiTuiuDns6P4YU0nGVTRnHYq12jG8QVjNhe1Wgf6
go++ebCQZmZwATqxOggaN0islnnarRiEuoXy8a6ruCDVqgqREFamgDbevzC5NJJeLykQgBu1l72R
bfK+ZZavbp8AUIX4lTjgWDMvhldN15kKdjTGMFDOSMoThcTU9p5AWZCY28z7yaYq00vgHYXbFFb8
jwcw4YDP3M+debJAUOuQRJ7BOU7FV0A1Mlb7DX3WMf0GPPF3WSrDPxOiVrL5K6KM1zbeeWpTxnLd
ydOwqLrA3XruVreo7gvDiP77NshlBRDHOcUWtAld4sGCIRnug4EJ8wfVXs2TO2sZTShLjWCnUmgx
Hez822C+BrTrx70hnNPtXaRS28rDaCEeeik8iBJ2xSpuQ9egJ35J0FL+xbseA89B6w7fjfV9zTw4
SfKTFPEwabA0n26vQcRiSgT+s7vZ2tN/HzmISSmWwCTEO359q9qGB2LRXMg0IfyuYjhIwlaNxPP5
Up3hcQPXG1JktqghEm0QDMcSdfZiFQU6/NaCFXN2vcjAI46XEBV5QgFWUlarV4gHZuD13T8hEMss
PLJ9NAFhZ/w2dddZcPweDGk6QBw/BLr/wMqemMiyB/V1dV/QaAGC3gulJTdEyrBGY+eZp4kmeXsv
8kzkw1zkQANY85u0GAn3j1lQa43pHZd0tXDATnJ9ctn3k8c2IK4lDPQwVwF4nyeNJgkTPHOfYFuV
V7DqtqeoODIdSwJb3E6jKF8ilQggX3laH0pipKqDZzz9RJIuKgzuAD9GT0E4ulRYjxVCgQWz4Oqr
D3zM1IJWUZKEJiHpfxgg9XyXji2H/5y5nVUTTCRju/GyVKCzxXSXDOiiU0w+xwTWFroNF9/dTebt
iBBC9rgokErAW+qoY8Iv/grYVvEOpej7pk7ONT1BJb9r7S4EeSq1OWtbZfVok0xVZ8jdBJfKFiPi
NhEdZXFsAbFgmswCtQzWtaKezPSQX9zNDgtwFk1fvncpSsFMKCpks2o+GE97puUKxSa9orUMZvXs
TM+7k8iRsUp6ej0zQjB219vJ87dv8yw3PyCV8c+YIKxvpTe4JbyLjmSxgFdHufOO5qlhlqsEgfmS
qbLOeCyN27ThQlpQUGZTvrzH9AJXFe+sv6rQxnQcNGHvXVG+L1evy4EEuryWKv+kXck1Djioqp7i
Eb9euasISPxnTvRhtcRZa6Iv2SsBlTI5bpYqxNIA+110sQWxMibFd/g3a+kuBxf40rMtjk5ID598
5+aW0pQQ4KeWsC/UIQ7DE9b1S02cCwjQpSNdyt0v9+CWAQv39GT5+EKsUOoiluX8K6WpWWQiXA2J
Ury7n/WtVizAte6qXsCbbVNDq9vz9GuoZCx4LcS0JiZRqIykSHHRp2sx+IevjbwdH1bDWlj1HGEp
stJH/XAcm4qjseH30ba6INnHOyCkimW2GjzJYb+f7Byw83EZGQ0Vo5S53Q86FY8+encv3qgc131s
oFJV68UxqEq5knzcLnCYOPZhU8GlZCt4Ibd40qWl/Nv9x6s5n8n/Izo06vRGj1ut0C2mLZ6nBPwI
Pv+wSCXOpBF5TyW6rohhtW4Yh+8F/iVUf7ENZjgybBG4AIVYE08bf6xH+i1Dw4tWSGkVvvIuCHjY
EyM6SrCrnwnmX3cH7T65Uk093GtBsYo4xmH2uq+xX4jCGdILerFsiA5zYCBUYc4486nDN1k1tlmN
+WP29Diid+MxbEeJNNNPeNS1uNbnQBcC6i74lJ4JUWIkemu7AwVeHTpVnaGwSlsEHi5oWW2Hy3DM
ew7BIl4RVgQNcbaPnyapnANaX8cJlCEByxWCtyBXHyJ6dA6ubsjTnJLbdhTBxuDcTjvuC1c0tLkA
/bxMIWCD6Oiiz+ohFs+V86sxdbXNltsynqMXI354wymjLYEq0CPQpz4siojAT72iXJDKjSPwj5Dr
/ftHpbN05agsgCRz2yIBTVqHvx/Y31EWRCQnmr5GEErihNXgXRNceYLN1S+EXevoaqmBBUsML4Ag
VBO8kRO6DG8++3CUl0Fl87q95gc7Q5L8AnUC5FGPTmM3R0uOfZ+f59LyFhgcvUy6uLE+zRHhVDd/
YIKEnMF6csLgAgdL9KRqoSnREryAybN6w4CApgQEgpbAOi7JItEpkOcMD4df7gyJ0Fn5fh5mP1Lq
Z3sowTYGYgbE1UJR5jxNgQq/NSabJxGTvZn4ozlUgY1Wz9/C2Dz4DDysWTqoMMZ/1+qyE1BWJTyC
MKQetfzNf8K4zSgJFRShUQAppzQD9Uks7Jm1lSBrTTU1RrIkbjoFYaRGWuu8qgPXmGK1sjlQbVIr
u0pN16ZH0Gk/+kE2W0+9AIsvkmKsbpW0t54iEx1Q6wBAMjBwJ+drwz1BEdpHtN4e5QP0TN2tTKQe
oalS9qou3gKDZd0aP3BdDuPAhtXBreopCSx2rhzkomUnqWdM8wVQkycpElV9v6Z4Sj1OLlqzUmd+
wGVCMIh75WeLFEMAqbCBtulu1apMd7neojbMt4cJRoXo352oqQAz2bFQnTltNsoE8+X1j/mA8mmJ
DuEAmd4n4x5PDajGmad256b1ds4ItMhx2SyMuI6xOp1AXSezaPVxI5dbTwt3jIsKfF//UjsfQeCo
HHhNyiHLTVUv6axeUkqbASP1J8diowqH8o6Dhv11L3wx6oIn9MynQrFUuX8nVqbcE92hu+Y4ITaZ
r/iXc5tnJDZ9fXqHcUX6YX0c1iztT75A8gvYXYevSQlzEMuyqiYcyqBMKPCgm/QelhV9euqfcFOi
ePZ1mXvgaJseYfjBAj1JNrUTRy0MkVnZWayDPAdR0RlXDdMxjR4jjM2djOFCFkGsOFDHYufLY3Fa
rGz/QDYvh/+c6EF7bk86PPUYYJ7NiBhCkb7E7Ge4bimjS6/B+hRNj/Kxzob6azYs6GHXptJN4LEx
Rz5Yre7iGTkYEV1DhMyduQp80PbrLm4XfVbeXNob41QpfkIlxoCdwkSfp9Kpi38f3Lz9Mdq+r/1O
w6bzcvJZOdHXR2i9ozIi+XBBcK3HyEVjeZWzrhgVVBTkbzV64k8v0ICCKm57wNExQMl5qWpljGcU
SWVPQ9/TBjlDadl2vM8X1nqcWMzK20xIeAVtxXVF+PM2kfGgnlKsQ1Ejz3Qu6raHWfy0mWNpvrSt
P7YyWB3lfjDDO+kmhskUYP+0/r6tnX+LK6mtzs9quRqu1/0FLRZ6ji1OpGDACAEc4emaXdx9ot3d
I3qTTHzQGoYpwx29rEopkPeMGs9LDiSnky1DA2rRCmSc9ncbP49FiE7gyRlqgI0kUscA22DVxN+/
gZfZXr1caygJPnpU+T6qZNKmmrKwjELftVhbjoDdX6J+icLcLXkeVk3fWiQ2FrEAGeTe8wB9qiWn
Yp5LhygZnkZFyZBQ5U45rmI4zRwYN7hdk4RxETdrr0oQpyUj4cL4ud7PKTGZ7gGhjUuueWGIvQC7
rn+HltQyHzGtdwC8njESGICykY0krmB4rivgKCVb7vr+FyqhUKW1VYGamxB2ni66+w5ZI2FXjBDL
BxeZjWc/ktgJjG3wRYrQ+b03zY+F8OKJQtkr7gGGRVv+/tk5iHCu36APbJa+kiSnZEIvylEK4UmE
G1NQ9PCoktvlvn5rvP7HHtBZF36NtSLgk3WhZO5fPrSpk+SWrxiL+c8OT+wK7/8q6P6tzMc+24cH
EELGRYrg8mJxK/kuKtXuC25VOYptQiLqVXZ3AukYma7KuZdtxAy+u1+CMf+C9LOcDTBjo6xmp3h8
911uyN/ZxSJmpN4Zvf91lehzblb4BSaV16WBSJuPl0rxk0SoKgyV8s1l8cjS1uSst2UcH+V/ZMkk
RI9u7qO8nvK3WOpG4TRIx4TpIm3Bk8qNNBHr6Yb69oS0RT5VihOXRGIgJWnOqbEzCXXWYU3c9pSa
Te4Z9jUwXcACvaFYvPir0gO0NFIunlsf5IYacup/ZYFcGq7PsxAqz3qqwZT+QYbr7/yBu+ILwBRV
F8bC137ur7p9hvGANK3vunye+lZXvENZ5wYL6QgrZuWLO/Y7ndRCJvha7U7Nhh2xsMIWS2YGpgzz
+dHKrp5a0iEQf8I6r/kyEUPru0+U/jUnEzNNz+wj+u65RT0o2c8yUR49QscrPxpTV1EcuFa/s2LC
nEMw5jGu6VvOxP7RbioH21xUpN39Hz5ozlkwHQrsBwfiWpMAEBROHsQiadGjhTKyZnFb163KnEI1
VRHTakKNQLr2669EQ5gaHZWoVm23jwLX8HTwkzpo0OxHQaPxssCUw6gYt+GDpI3zi7jFM96iyuqA
epj16YT72lLQnGxOQy4sbybtW3OCqqiWxXCLRiElD36uT5XDriF0EYaGOZMp/CrYrfWsgbwhQGyW
cc644ocCyM30qbdT/sQNYz2qzRd3K+JxUL3Kafl+v3qzNgVEdxeQkod8h9f3srVf/HyZdbMeHfXt
2Fhe9typwevlghhMI8gZV03vB8OPMx8Ea1xcMkDt+vlXdVnfAtIHti6WoKe/oikfH+t+NzrcyIOi
ewGEmkE/dQCSfPRzW11r8UU/v9s10USFTCDsuTxREDUdM+DhHMHcQSQmJ5vcZbmWn83gnh0Y+NVX
w6bVQea6mjQqkciFxMM/C4qFyJPV3gJ4dZBpZIv3OBz1UVooFj5fbcBS5Q+9eBXFV621snKPTpz8
yhzFSzNids+XcPxtoINSBqTe0613GwSwaWWv1eweSy6E2BLXPWkjf4oga3SwZY3MSyLYkiVHKBfn
CKkdFzo+uESyHicgwLOIFfNAznTg7hxUAZ2GhYav6pohz20W44RHWeLLb/xI0rzCqnXAtGABZrSy
TmickF23BxzJ93dUUQIHJ/WuHJOiBg4STGP2cWP3Rbz+HcDxLvY+1aY30How3hYBSDaVi/VsZADc
Q/3Nu2kqgtUY+r9P5/wu8tIywoO25rJeXMmWPJn7GuOwEzdqGJJnqX99DI8SX5jqKpxuYmQ/jj5O
H1a7Pqal7kXXj6VeVOf2aqjUWfSaIg45f3Rl/XvvSF8Xvw8AGDatYjh7Wzc0baqvF9LC54Wr2vrf
1EuqTDE9ZvDI5bmVwnoK2IOq+Ck5jAYmzRDBMO+T6fQxlx7WuJFhLwUsr89ktX6PHhKmGNIoc+a0
gK1pYTkOiM8DplIbLt/pU8Imkzdvzmy46vukt89sNtxzlgYHsPbdfnPSJOa6nbCgTTiTksit5c7v
1A8fB2m10DHokRti3nfwRfkl97o5ISei7UiIo95ttS0XoeiNxgZAyw+/+ivj0RZvSZUpti1BZJkQ
lTIYxkvBu0VZjEuKJ9W+qrcdCPpf9L4fsVTa1TVt0d916rZhsuq2uyDiDySpJCTAa15Z0/Fx96a9
5SGFhmTCtXhIbhb4Lioj4tnYOMw2f7hWimPTQmfyjnbA+zLdaGXZQ7G8duBWN5In9YiYbKIxuX+a
F1unPVNSoM9320wvmNGO5liERnuF9F5eWqYLfip143vOp/n3+uDhiPOOIOEG2N3WARGDKmFtshbk
TL8ZKxaNTkWtb/WAVKWNvKSr8nR4F785Z/Q2dhyb/QUtf5ekcs/NZdHI6RhMrBRETz3yQe/R66YF
R8Pvss59hXmE5uLIdmrJiuLbeaSlpv7lNvHItUUvqVTsXyu1trGhEa5Z+CMTqtosCKE/H9jR4vQJ
p7+YSpxYL+uAXvb+kmOGG+onOn3XrccB1beHZ3AOEmWFkIMIBtSlt0jrweTPorsckJ990bmPBR0l
VyoLpQFXuYAtqzLaEZTjundJDU/DssyF4sLJNv3lkDv5wblXqp54+XDHe8NRSTcP9V7NbEZMVoA1
TNGAb7EE4NLFMsjKLQIY8AHfNf3P/jEg1eqydpFtvvCetlZdjIprD3O8vGyG4CWtebWEASUoN4yR
8vdwg0P38Rj6MG6OxEYEHwTcU5fq1f4NITy++Wytqzu2DomWhSkB0mfI+/pfrGILzOVcCynt9O/V
FL9fPKisXhOFoWBT9UEkNWfBqB34ziDTojIr746+9igCjB72AMi6cKmw82fwOn/p55WdizU7pf0r
0LrUktw/MiFP5mXww1ijAgxzjP3yEX72LNdOC7v5ixGfAb/vL+2NG1H8b0u+Ju1a4r+FyCtepTI/
0U6q9+WSmZMEMz4GaT8bc+k44y+ZSGzUOxwPIgg8GB8o+/qeiEIpCNAbm4MDR/OESpgN+om4vCHn
tX3eYunIc0VR+5WPTG8xoEsdQhN4fPA895s57oi/98qNQinO219SuDpQTKnXg3crSzGDLgRcOAsZ
UMXizH8SeAVAfyAK4Aq3Em7LlWp1JWZDWVA7ZuWgVVkaZBL4XYYgKf2OUY3/QUistOBL3Bo0wrtW
53/AO6Nwcu1g9LgEEoySByTmDNUpB8mYamJ2DYqMG4i3HI66MgkXGdVdydLkipSTZgV+uhyq7we9
6NR92LJlXzss2cAVcmv5tMdPiDKN+0o1Lcg0V3Q2oeWB50Xcau2AvmQKTx0bCnR4ycaCxm1Pfu1v
YlomqVHv0mZJL3WtCpGRJ4qRQ2judi3L4GdlH0RDm9bQLLf/8z6LF0kABEw1og7IljkyDmygoPsV
ac4c6AUmCuEeCJk7A/K0ZO0Y2/3Oi3pdYRGVB/igz2u3eXCVyp0nMnNBVmko33Ft5Tb4Xlq5zdK6
pOU5XW90Nn6X25kCrZfBcF0DRNmuyzVqOk+svb3GU4VshlrOzt3w2m9DGd0d6Wor0UYW0LG+U5GB
7Z7Pts169dLLLT4+PdKwTFh/rAUPilqDWuchefM/hi8fXeF5iZrEp37MJLXFtBNhgitx9M+qbRyB
mTHuTqt6AKQ9kDjB6BG+q5+TW4eAyH2iXcaFCszR1s8NWUlK4tlI6rIJ0Py2Jp/AiP852J7VXmnV
0bIRzlNxHj+KndvlqDdv1j6MBF2JqnN8SrdbXxhRVqy5V9Nt13/r0Y1CNglCCLGl6B3lma8sI5ZX
EitF09C9us889S5U0lCU1WUJVyGN0Ysbvy6UPbC5lgHEiP14X5IWzQ+J0KMSAk32WxQiAoYxPTZy
Y1aGjo+yKqvFuTOhlHAoDse6RRNusNYTglZGqxa6y6YZ0iAqYgVHeFl9E/45mpB9FFrvCXEc7xGX
hOOST5J/GrJ2+Ycn7DvgXzkjZISY5yBk3bbt5f21NUctYgWaiOjWbuCHEVKlTpQrq++jMsfy7ING
R6rUarPrHV/sWIMfpLX8UPZUaX3MU4HaX7QnWxSXRvOjvUm0NS6wuFXm+a+KvCToZeiU/015mAf2
r0Q0HgXu66IuCcU4empje0qzwc9HfskPSr7zOZpcLpl4nEeZEEdLf231esYnElwSLrP/s+rNLsnX
DGP/mQSJfmtJacHeJBceVOYfdO38on3xU/Q2CsabPgulho002tIzRAiSrh/A4QTQuYyC56jKcbii
2iWxPlVp1kbGRcr/9AYKhlgmO9/zvXCn2dJLR3vb8Pwc+IsPTguzYRmZqvbm1Lzm2EDCsGSfaG+Y
T7lU15rRx/HgqGG4HPpZFnoWpwPFjDBhhOXxkyDWJxPnex9iP8y1ExA9N1w9aJ83P0R9tKQFJzdg
BOKc/zy3TG11qVIlCJ57u+J28dgeteorjv3topVL+5KqYIAFldFqrLJsXydc96KsQhIhQD/mS4rJ
a6KZijw33vcDPK99glJVjIpUuGYryWu9xjjY/qWhGYDfVhbevwxILu8get8Q/I9k0ebc2nh0PHvq
upM/qjNxFjlbYYWt1/aXj4CaQpc+gz/2/bSntUHRX2KYvovB77auRlQ/3Qizya5u7fasucgpeqbr
Hbc0yFDDy7znlwmBymjjmS+j2fwzAEDkEulOW4iMiWWiWbIBnWCP4wFtrgYuC3ovUrAhkCiKRGov
TstKPdnWD7MC1iEW4OjermT097w2AJNpd2eoDtw1oC8rL2ZwmbwoB4S9lUdng9alBzSSC3UP8Z4P
bvUOTNF0StkHGvfk5G1HcMPsxYYBJKvVfmn/OnI6LfORcthoW9z5/jyuu83D84NS88mE1v5T6CRR
jpUtkxD34O7kQA+xVDuu8TaFG6Ta8MrNu175ylbEMjtQVYaH5dbUs3bfchLwwwAUHRDI0DRsoqgr
AJIO2DEkRTeWvJO5fQDMgZEyTa2470+gicNLTqcee2sz/Kwhr32NBst1+mTFsZgerpyovonfxxGX
kMIOC8Fau+U99rzsi0dqXI1Bt5i6u9ovISXTN8X0nAPL6rnHg4i8sf+CC7CxQSZ7wor+soWoVAXu
TAP1EcMiJVGDOOs4BHtuLA0buZvrc83tZtbZbdXB/YffmIaLYCE/Fxxi9BP6JL3C55eMs51N8brc
GDPaOc3PnKMMgRyquMMkm/4Y0wazvKr7JR0RnEb3526LvEn0mDnAtHbiY4+18KrUafQ4tFDZvxe3
Blp9ZyFLR1SJ6ius2ad8dTgbK+HgcDh5V/pIxkf3rY87WCBawOoTg0tzJIzyOfRyBCEiHzu9y37M
PKgMJC3LQunOCm7pGCvP5sqPXw1Zxr4oHxA+YOXzI2XrPwxjObqu5qw+sNNzitCV7PWu4fRkiaIO
YHVC//8gSMehM/YICe/KxZn5qlG0lFj3rW65jCq07qhECh1eYWSCaH5aDme1G7ULcS5HT9i7oPc4
+e8VN8f8CCwJFOGZFb2Mu/i42a7sLiNrOPh5zboYNX4ExOfsM7FQXEVwlRDGihQ//8TKL0KZ6En2
gqg2zkiuxCaGyH64Hz3pl4pmHXn3Rrt97rj5eFC2rDTPY9QSRijWLO48fZDLeCLzvq7y1mbGQ65N
i1cRysEjEeI1cZgj1sJ4rpKyhQY1kntIeuNYfvVuiHNsBiJhAI1hJ8mSMJeYDqRDkm+pD23AuVYs
Iqf4mYB8x1n9Qpn2qb/K2VVcSDVA2vMG0bX5aDHyJnIPKk1FnIGUmveQMxsvfj3vHyvUmktCZHOk
fG9vsbID5oVgnCRdNolN7hv7GqXtqh0RrBZcuXhctnkxrkXMcdCxPO+ZFJ34W2TB/xT44JgCy6Ns
G/cIiFyMJBj2CnPqLmy3ki440ba7ucRIIIf5ITr0Taek1tSoWEL+0vI8g/hoLu0bLL5u8OOGZIMK
WE8gxOknlFmNnAFm/taiouR5mnhNwgnCmC9mFMZ8RvQoa11SWCVG4HhO4ZULa8ZwzCaoIz32rima
uW7+HbTCmx9hfjWyJL7c7ByeEhkQ1A/ILvMIVtrwGYxvfnFDsk5zcHIuUNj48XWuQtjJlaHBu4Ib
3wp/ETxqgjQAIeB3yqaPhhl1P+9cyjHWMWcdlsrNnUIB3+/AwgFovNyd5xYea54qGmeSojtyU1VV
kvIfjqKgBnUXyezWUMnnTSKX16Aa8UmRZOJ9r8YzSe8fXIXpLgRpy584K2pNu69DIpONV8ZCvp5i
emV7eIbP7EKf3KwPCtOREDPbHfkqT4WIepRsE0QAKusv86HJU0DwbC2U1remRFwSl/iHtaYd22HH
GBlK0yR3XQb0EmPZgtDntGq0A8NLiCBbeUiubskzSyP1VP7gOa9wqiOfSobDbGZmqJLb2myBsRSl
8x354XpXwvrHfepovtcahbFo6bjJ7mkSk1+1qr4/oxjK1pjLaqn6jCyLmkSikXyBU7hU3RE9tUtv
mJpEErPMhZE536FUO6pVuodZ9KK+M23kAZHDNbyR65Y12qzMKrTXKfWkZskWLlxx80IBXQLzZL/1
QQ/NQv5mITf2tgZKzwYtZnHWdY9b4jWRbibrU98QCLZvbsRmbzauraNVrQNuGP1N6i7O9euuO4sh
lMesUGYLTGdwxNgGLeGwvtLLVzD/nUilFSDq93dcb8rSZHI9r8EUSna1vXoeV+nAojP/fc57tHIe
r7ScONQO1VqRTBHY6YJl24MjL+zd6dMZhAwNwCorl08oJ67BO28AtZtskLFIEdOJYwZLSCbPyEcC
ilF9xcOGoZV1Ja8JkQqx2cOGnmP4iesILTjZGcNfPIQhEbbBXDVu8qPNs+uO0NCYz3WuK7Phpv3Z
KmGmyqNPDc/lTxHFMFIgUXnQkR5KjnJZBdHzf9AZBls8PTT9LUC1bwa2jWPQJBMRHOL3T4hBydvl
v7PABGzA+r0YoVRzaXtuHqMiDhiDkJ7N60U9kjFVf2zCFCovOtC1OFF8+qAiQyVElsShFEe+4vH8
GGDFG5/A6xVACgwHy+DCnOnlIujdSBLc3TpzDt+gUQHkx4u9dGsBgDxFyE8Ijkqw6stHV3fSj/qh
ET1ohg2lIlNuK5Dta1pUnayxuCduTvJrLSKcqRwdYgAJF4+g78OnvovjFdwNtMv5nTtAkx42JeqH
2iFk+F+hNqhooxqpFz90L3BXPEWzwE+i9rP9Xxsp8dUrBFXT6SYaYB+JT2CWQ2tD63orii9w+Q2l
fTFBYchiqexx0yz2chfuh0BZi3+3suxKw4Yc3mLZzsSOD1Rr6XADZcJ0qNXYyOUn8Qfwy5BdXlXl
0twq9ogI6DQzhhSe2g1Nj77obHQ+Nd/gxJdTcpFHyDhVj6nDXhfndEJbNtPd6EbzGtgiIlt9vVWO
v06uW4z+SMpqW8nquiUG/o14JpS3qZGZil70H6f2xGtlsH7PqVWLD4Jhz+ECo3x1hIBjMDTfzdNd
sb3TwwjWL+7MJJINlCEx2gqBFRo4ByG46HR/bXFXkHYeOaEJHoeqj9KwHg4nIPxD1haqN6aAJDWc
eFc5cL6h4fk+3oK+nFn2gvFOzWH7SevAmJVgLefYe0eSKdQtEUmx7ZDuPsy9xgXbYzPjKHG/crA9
RJvuQ5HbXX5QGpEVeniFzCEJclV23Knl+zj5ThMCIbUSkiRpWTlhHIcCxCGCR5ANSDOMghYO3ki6
mW70p5vOzUBN4Tel/8pQ8jpPkQuC2Cjao3fL1/GHKO5flgUJuAsCT0FZLBM4YDNovjhy3VF07EJt
Xha65eBOyj/hYHPLA1K0BIW2FOIlnOrPDbvIUBs2gB5ewm+uF4aPkNCgjrX1CGsBTkl1SdEqkFyq
SpGEq7LHJ6xKstFJDoKcUydC6nWHpEvvz80w/qojAKxzxDnrxhKZAf23AKgA4ilKJhhz2W9LpPDo
m6Z/XfEdrmsbyihZzWFWQu/Fcj+8nmqAkIUXPEL3lcxPh6AonC4fwiE/BzmKRg61pFKothD9I0tQ
PaU/bLBlbmNgowt+E5uDnlw8gjAddImr5FgRqVzNrlT00MaYKN4HH3bjBuhznnhEpIMtadWXpo2o
piSURbe8DuUCx85FGFREv+zTtKtWtvz4ptKGaYZqY9Q6jfnLK/05JDlUiFoxvfbUqMrZabIyaPd0
N+KkJ7sLY5uLj04f0lKHENtvWHFXx1B5NcOOSe59sTN1rXFtGH0GddiSeoAHhAuA9hkosq7LjKvM
Kns+GyKNg58ZaTRUfAMkTP/LdFQ6TxP3QPc8a0PJ1v4x/YycKlMqREm+L4ALhSZsJjRZTwMglLNJ
hKHC6UEwVFjAmTCoNShw11CSVCoLR5HNj7joON4B3BZSiR8SOWrU2goo/z53hg9haXcPMBsotad2
lNFHV6UDAyvsXjvAwLx2mPEI2p5Fc1xnCOPMgLWEYwOqmqxslEX41MH6bhoovj1uX13YqRzjot+L
b/f0ob5BQI5SoQaTPqKki4l3EHc81Y8lk0v3DcXWUjRYGPrQtSzpEMyYh+Gi7qQhBXorgByTqKF6
NLsCK+hMCeVk8cbIfbbJ0SxGFfL9Hh5S0M/e00iASIFL/k9cuuglMNzdfQPgWA0qDwE8gTr6zjTk
trjJ9gFs31qOrP4yjiu2QGroj8J9P/se79UhhWNSNa71io2eaFF7wvsy55hIeT+1Ie88LRfyiLUV
pL64iyY7RRyM+RUDTbvcfEbeJaFOQ3CN6fvBq1XOH1ukkYGbHuuWP5KIelG36J2CReKF7B3Lwq8N
q7PKcU0o+I3ty3wKwg/c9jC2AwwczQLKERpwDj9zPJ0+jQQjIJdeDC6YxZZZuokQHepst9CWiNOu
bJhfBs+7gc0AkL1zKsEj9dnVBwv0RhZjCgn1ES6k98PiBX1JEqDOINAXheLGrxuTzlcSf6z4A1nS
nPIasEZ3B8hARjGFIMEHrxmtNtinLT+7YWAviTwG2eylICGfbB+EDIjH9GNkv2TGKoVczy4u+C1P
PrVZWFaGwgbdtWkxIaAhCQTiF5O3lMZMDEqnYSKG0vlwP9LnKaGlDRr1rh7XPRsylKF7ENiyrTVJ
yIOLCa9CPo6Il+lJ17DNMk/yCFuHAbk6YaCsRpjL9Hf0DnDmGcrFb/jKg2uCd8dnugj+EmjESSjc
fKMF7Jax0UU79UPyR8hHr7WRbLGfBky27xxAvDXgyBspQucjyU0IpXAt7l7SVzd4+YxcyoVGArBN
FoSMgAe8BsfmNigiTPWOW+Pw1F+nxdsQ/1jgScZwK3a2mSMkYrL9Iir4hYnecql71ckdHE12Xmnm
DsrJcP/HfFasYsnBlP5KQnJWjmJG/zCDTIQEJXhiwRZB9VX8w62rADRpY5EwtnsVxo6FZrLYlusT
8XCp6q/hrkPSqOqnX33c2/UUXArg/nMdaik8JfX34Oh4hGYBW36UNfShxYElpQox3mjyvCJFIkXi
z3nvjQkTl3ElwYMn8IPvDcyYz8iBoMU+BJNMRQQ99PoUZzWL+ob25Pj6ysr++g0osv/G7ZJQKT9g
3myF3BuSYksVNyjpeOYyzQBqi0zSbRrgZUr3dKDYhccSGXc/2Edc8fxvencw0LC+4ja7t6Q8dhZi
jph076ejqvHlLL1IBhnOAtaEz/4eoeG2IWf3EPEfj+1LVFHtukPY9Iu/+j3xOaDKP18LWig+LHRf
fLNKCwcC9PYpZl9VEStq6FFRnVzs9OJ0EH9Rvboc+QbVrUfB6XoCgCuBh3azyk7NEacL8wTtad8T
vMaJjxHNrl8Pigeveb+vleAfAVtzODOxVfYffwCc1LLcVQsE7XkUY6HfsQDorfGiR5veU2kpqiQS
g7aF6uN/9/eBz8XlAN7mXAjwCDY47iZq9U/FbTBV9Iyuv6NFufneePCftKGJIGbF/LQ49XxuJ5kY
+OgvOl733oI1VM70X1Hmwdii/osCTqisPtTSigK94yyREelDlU1GvNyGOMRv+PNsx1hUEylH2vUe
sNWuxuUFWiTATHyj+Odwkm4LgY3arWSitrPYRxRGHmssM440rqGOd6kHfJYvU4jNzHObAT/D340p
UFkHvbnkvI+fSQlUWNsnC2B7wnEo7YDBmMawxexe9aEXdYq8UiENje2OQI1Ew81+mMu4jEFPVyT2
0s3MJ+QBHSBv9AkwxEXSsyaTUdCjNphtyysmBYbE2aUwa++bbE/6SpQnHOt+SF8TJGUirPyyH9nW
lGREDEfWPtuZ9AQr+Gh3KSkb9h7JbuX7e4gCDMC1wiazihri1bpbdn0qoeqJ5zrPycc/32I7gOWi
EOL7EOS2SMZ3Oh/C1JETWgZY7Yai80MSP2ZBVd1dCF5LeZ/7sfD7hNP3zJO4qlwR4i1DHgR4oRjo
dLFBYq/FOfRFDPsxHQIyBegQWW5tiB+OUM6vYVgNSQGjxbet39NSdF3sOFry16LWUewcq9hVAx+I
9zdC715yj7evmtTgzDpyhOqobeliN2y4U/VFPRlttiHkUmEVN6854Rn+ZV3ZhWUPkZj6NLD8ZIVA
E5GiV0AsPzfvxfoTsE0iSw3opr1971yAUZttow2LWGkHFixuaLJzzkNtHNSq0aJxoXmDRnN5rSan
/Mm8V5X5+h/rZjoP6emwzIRdImpRg+3B0D1dBx347v2rlPr+UvY1UlFpNnpkU7RtL4DF0ivtm2PO
wXWTsIDSJX2F/HC3jg7t7A+fYIfRF3yRrN3tXd8i8Oq8/DNepqcMIQC9VotBmCn7zVl4jBUtTxVF
2tV5J8sETk5KLYLQ1hIh+82k+J9lIeW4y0NGIGaPuiVu8DWu5+iBP+/uDPVnk02wpfmbFI4vuDos
PkO7m+pH15Y5tgGqJgVLEhBLz54By3CeDoDJcMcKAzeQKSCizKtnkzM4rjI47sTEoncYJxQL6/tI
nO+e4DxwSRP4JPOvEfcFmVfJhPLDDfh8QnSZZ3A8335wWI41OSRTBo/rpA+/cNIMeZVCQ9TTAbE1
oEYulmrAlrrJJymePh4CBdi4elb2TLpfczXwrVH3gjjYsymlSg8qoitmJXf9URqiFPahgOUzAV6U
ysO32iuSIYmC6+FsQSMOj8G95A/A7DfSk4Zw/xLDTqbxnla3dqCNo3HPobASlse4V5MoCSaQdJEu
+etj9m314EhZ7Rp+kHvgtR1Fo7YMm+y/QsW1pjxYgqhG2WNOQAtINxAAMLL58rRrkuZbdjEPlu52
EM27WBfTZmvHw5OdZfUoICltNdF1/Aeg3DPIuH5GVarUKT5UVRqfSJ8VPRKAPm1GdVSNhg2B9CHE
OYaDSteywWXYigOiIdYrNoEsh7buRicv+bVI/lGj735hCnaoHXvDKUeuttpykM4VQc/KUt2XQQ/8
7UlMwkxwxsK1EMAR5qAZi9APDjzbggZkiUp8lP8gw8TsshLC31OMJpqFW/xa3G7vxeIijx60Hoyb
/g3v30BJ5LAklMzTbiwpLrdN31I1xWPn++XBYr6R21qvLsifa579vH+o1sDEn+M7s3HhYGphSAAN
HNl2qE4dCH50Nua/UTfC1hv7/CEGxyywUmL36DZUfgKl532SQjh3dNwCV5w1JfyySGlGpMHnOc9s
bpB5kpdgdZ/XfbTqt/lgjSCIyHY7U4VqR+pmMHmrw611YHzx/zA2a3reCJTpUUqCJ+xS4TV8SA1w
9XFwhzQqz7k9a7siPmOFtyCxlrmmiv6aVkccUQqfRIRTguip8XKi8h5rNvV6l6ZE8NrXIyh3I8QZ
BWpIknvhJ9fzpV462Sgv40+jZQVeWMj1lXLHkbBB1/j4mI36gA5rIdn8hIKhXB+AQ9sL9yaaV6/9
CUO21OwU4QMe9PWHPwLy1IUiZ6k1lhs+/cM2ZdRnve7ojHmt1loo0Mebf6UmoUzUGLf/UZB59s1I
+fQsF0zh6rVLlKPqNAnlq20uUjXhafWX402LQ73pyxODn07ZXUEjLPm1T4U3awgmTcuHy1+GwCpw
Y0IEwHnPT42hnAPmj3olDb3Sot0bnd4Nz6Cw7Z0ejVq1newXWyGzOzei6ZEiL29KDRbnsuiC1HOq
0XLymUggLbXvKBTrpDP6DmbXuqREfO+BUufdj4qm6WpQ+I0eoDXDtCHHKEy+jRnLxu8oqgBjO8rc
fanwsQ4E4M76Epy19yGEPv1PDKvHg5KR1wr8fTdlomKgcmCcPT5ehVjiRy8XtGzjdABDXpV8N77c
Ck9PmT3NnHe93kyvNqIyESTEqjTFgVZEMTJ8SinkAGG+T5hdNra7dh+bl3PmDxNMIcIjQ2EMNHk+
L0HRcvJMLsj6sQf6YqWeNwuaaz3tsg2Hql85b/dOAnNQKa+1hI3QL6Dp0wsifaqanScy5yCfOQtJ
lLKQjuTydhedxsc5HgOAwymitv5pW7JwiWSSFk0chVExHkx5IMAbucxgDiCC9g4NzGFvRIb8zSri
9cOo5LEM0ANGyhT3jQTT+jhnzJoEfuQUuqKXs4KyTewAePdendu6gw1h2rYt95IkCfT6AjKUve/q
CfVckovxYJQGltb/O/h39zHx8qMyujzMYYmX4R0hBxw4b+ZEs154Rp1aOlVzYAWGc3iG/TmO6YWe
to/4vOac+WSbb/cUD1L+R54FEuVtLJAD671bUr0IknSG0knNp2gUdkHZdFj+cOzF8GWBVyhC5QRv
FhsW6PW2zP8NRZPHzi5XQ4PvzM7G22r/goRwk5JWHl1Fc/rKHStsalbUiOLdBJw1Q+NjpA4SRQPE
rNdYMB6ObuZNjGxnxSn7ySeSKEYN9xui4OGI3A+WWBbaRsTL4wvInBTdD61bqaz2fHfE7xRMJi1s
KT5giR48KMk+aNTKXbEdzaq2TkTHxk617lSdffRPZTb0K3APxYaoEzW/C7PoojynXd/hv37XloJK
aT+KdAoTdZYz6en1kVtVGp0dv9evyxtA37MNxTvxQmQvLHhHuXH1ZqWroLMgMIH9Qp9nasIXAXTv
XM0TpRdNwdO8PJLHHZ9MOxi2eCBOWinhS2OVkYyPJan/rD/KHy0pc3FfAnTBwnKsvcnofjGQOKm1
p2Z+gS90nhfJQ26viERGpyGcNL01/q9Cc+OMN1DwfDM59ErRxCItL4xA4fW+WAbLs53HIimXrZju
LTOiFHm8N6DMMFa4LdPg1zDINzVk2dfBBPYNsJRpf5chveLDcF8bjz6W4m6iQmqhu8XUwYdCIwGD
1P+LdykVdEF8AQBKbfY5F8klm3Nt+n94OdeNy2WbHMBpfSHCoqtWJ3NdKQfo1vyMNmVKa2YZ3P5f
btyMnSIPBqnJfJKGKgvHC9Fd2UOtunu4Oj6vPAAKYsBNs1g66H+ta391WLOlpxE+6LSs7UUlAsqR
s9g2RiyDTWNo7Q0m+UQtlBRYDzf7xX6kabT2gDnsvhayfzljuQEEdsrfNPa1mUFljU+cWY+tz7Y+
g42bsn4+WY5VueKMirrYzPQhYnmIuivFz3Xo0SlwgIdna5wkUc5c7m9nBFv9KMv46UqRf0CA85bz
TbyYU/19QDOeNyh1Oi4hKk/1mv2jHh75vlFLE3A7f0RfF4bIM3InOm6WyF8Mf6Xr34phoqLuHiT3
CVVOGwVdTycLG5oR2ebRuSYkB/IZ6RkQ3LrEA6XvUspB5xvKKJ8MJ1ZbGbT5UYdMCebD8n7Ape+S
nd9LKh3RRjYxWRugNDQ+RZu0ppFJSLjB7KsI4WAthIe6hLPEYiFj6bjTq6aCx+5sQztUfgpFlAR8
VGqzFNJM6kLuM0GchNT58Lv9QA1ZX108dkBa1O9zh5W1CHm7TgwjAzDy080B
`protect end_protected
