`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
K6MLXsHy1mE/e+BDKQWWCf+4ivx+zNnJ8O6cBeb3pUw6btsYq6X7MtHOz2Oz8HDGPA6q9x8lkpvp
HcdJOMY+HA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
P6xTgR8Sldnm8Q2SDl0KldP8Mxalhk+FQ8DKI5wS3in+vTjwT+0Qnq+F+NLFFYSjCVLQsvICID2y
uDTWUrzC2hBYfXhSogTyPkvWjKOEUhadOtQFmXVRiaRRmDsmYIP0VfzBDciE/+KgDZ8IlUPPc2cU
WqlOcJ/eLogYE6zQYMI=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
QdKj0eSWfm5SMookhXL5Mfkv6ZPZaxlVqSnBQx6Zt0SW9kTejDuRAfDQp4EiCm9dC8Y0Q5g8DAto
xJWkPZTunorz0KoMjqzfZLgIPVA5PGWbf1yF86jDL7ftFfK1/8E+/7kecMymdPwvYYkrdFLOrl83
j0kjqGJFjwWrjZ8CVV09XjFElDr4v/W+DOpUjCphuOH5LKetNJs0j1z+JTO6XyruGaCJzAbl5xfA
R3li4pGfWu8XeN8gITkQImYGrrJF42U+3XtYru5NbH2wQlg+/uqFprJWP947IwURkztN7oj5DsqW
VGP0FCt12yKYCT2AceNJcCSCSfsK4Pc0HB0raw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
mPUaOpmvmhBtVYCiUSfFBnEWc/b/39RU8W3MPTyFNUhf8hLULjpBea+PhKmrbx+gPsC6jLfNd/Xy
itAaLl+gJoHCpcTd0fHd0QVx5zBysFQ96p8lvwTAzlgiIf3KJfmwt8iSojdq84xPq65iSh5WwHu/
tEAPVBe9eTqEsegw5OQ=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
jrmiVyp7fll8pzeg0coNDePx3gVSGIxJxJB6Bfv2T7tlCbnb88FAvJzHLMoMUWGpWm5r2zw8eCKa
Re0+GzIsqFVL4pR1zaSSapK4xk4ypME+FriinPALL2yVdhs/1J+jPO4gjFoISVOsvns5g2dSuY3P
GJVpKqvQHiraQr52fdpU9xAyUKpykZT8l/DaSAGnjzaVdxVj+HEfd2wVvaJm2IxmKgnNA1zzVFzv
P08LRfOwoyCo4MCVekMYpFXSZriE/BwYHLhQ0uJrHSez7UD9w9riANFGHIoCRiRg998RhA8HIHyB
SviozKjzIIihOUGyb/M6tsh5Yc/fya86iklPYQ==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
KLs19GN1d72xAG6XSs7/+R2FVv4B0ae56gDUM2+UPaYIMAruFbPejUIaZmGcPW74627oECmrLsqv
yMhGuqy2Y0ZAH3mvlDb2l/KsIFLZJZNfnjHfIqdh2ln71HiLa9iLYqMfDqFpjbsNmlibkeIK6Ye1
6tjFbBzcYUfGzxxN86GVKIyqUC32+XUgV9CY07BtadF/xu9ANU8romdQ3zqjalL6iPbVHMGpO+ri
zswv6sMOd1tX74Na1ibUuhZG1Pyqcpbo+mRkfRQN/QptsqOS9K+PrfdE7Vhte7nW2/xYzDgGdjP0
IIGZJzDtIH+iqkAC+Hw6/elB7pBRqkRDetaGzA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1472240)
`protect data_block
m32k8HPm27Xy1sF3XgmUlhhdaxULN0v3NgSTxzON+3Z2mASsM4BptcgjLMnB5DQ88KbAh8F7Yafu
+YhW91jC7WTZf+DScWwFcR4dc85nCfeK77QuMp5btNH2/ZOzYXKYLBcFRh98o7+UDA8Gd4uXc1DD
NVjJzk3Y3WnRWUgA0HcroV35L5CtIVrxBOITIqOxwiJaqn6QpVbj90Mh5HUx2MYQmHemwLRWqINZ
1ygnpjummT9ak4WcJ/ihKPW/Yk/hX2kFC0E+jpPLJ4pGlHyO5KKSc4DnjEEW//hDsz8C+XxAeBA9
yZyl9UMji64VFpR/PQ/V8zZ/VmfIziP7IAPtigZc9ADvG1ZZ4rpaKK6R7BeOcEfXYYVaRh+sDXNt
/q6XWccAlM6VHsy6F+OGIGlEPvtdHkm+IKeiyh6e+F9tc406hVOA4u/4tHmmma2VUdCHCcl/T0ch
hW/rhKbarAXSNr4EfvBOVQwnGnq21gO1OxNKB/odM6DUk+Vc86RnVXeQR7owYKKLkk+QBMJaaQM9
3yXDg1oCzLqc9o/uS0WRKxPrDd/CvrWioA4BClkkBPXQNEX61KWYd08abDCSiUJbaAUxxa1JGqPs
BRx0F6LQtBnSZdopFIhl6aBxz0/zVEunEDQXdQP5zYBnTWGCK4X3XFYasR7EQXhMhQLizsbqKwGX
NMOW+sJ5cXYhMVlx7wuFKoCJUqPDm4C9QfuIoBRZGvDPJQzqsbwC0BcNfB14acwqT/vSXXZf+zDe
36uSoD29y6nlV2btY03j06Cye8NacFwZ7Vyl6izcvB9xcS9yzBGLA08OIXskV+Lc8QYJCa38SyZ5
IySFizxGZLuivM3cKbc1XanMH4c6+vl7R716ySsHIPkStDeqrVrnggCw97ecYalgakxcWaxJzhD3
pQFebis63xkqNj175DDhGflCZ+xmjI2uwPsif5fg1DBcALb8pv2las4cOA5OwKsX4BuY5iSVyuDm
Gn1gQGpq9mnZJOom6EcpJ+7S5ZCRAvi8lk9rkQQGD3m+F5fczpu59NuStUSxjfjKvfdyuXxipTkd
SLpXAnqkthcXJ1SfxyyInf0luzIG8RmocWJ85z0rWswbJSUe/tVIwAoEe/0VCp6dpC4KShfV2xIA
SIhWVpjdPxRAmqfql5X2DU3Jj6YSOMR9uHI7c3xdvqjSo6k1QJ0QJiOF71+GvjNPHQTkY4H1tYnQ
9Rtge11bByvapJ1UgWGn199u0Vl3uuJeC3/dfhTdmi2oPo93y4WkG13bdhE5pfxarYdKwiO8IKR3
mQdYsFh519XpHvy6IxSRqzdBsmSTl5mGfP0m0DdEvGtmmDWHeV7uMOpfX87HADJdPY1yqwsmhq2M
pYdjZnn3aLVYqbffv2GrYx46Au0AIU6oXHchw3YIpb19zmO+b8T7MYyMPvT1qPmj7HuoG8HUpYSh
37feP24Y6ZKoAjtleOUlFrZLfwip5DiEq/x9wMSXvbc4PoNGFeudmqEjJYTK7Jgyv4p7/2vPuWOR
8TUYwoiDeVH7ZNBuufR5rUACGCZYC2wZHE1S5Ks7DJVvV/4YUr7tKp8uQvkngTRKKvJYR/GX/YpE
SUdhYtU4gOi+iLFov/L2mBbhWPqXB8rMa47EpN7eSPXm3Z7z/+LltNIO1xq+Dt6Xn61uouahEtiW
xv+idnmfConFKDtlBwb6eP/bPgWKsE4L6ossUJbjx05POYE6Heltch6LABtkquyVQEagA4riQXQZ
EzMgrr9Ty4WxyjUnGjG+FCCx4K17HxSLEZoGJGVbGdCGSDTkO3TrJXaWpR4sTo+c2v8RPO5W7D/B
MoP3Os8GTO7KobuFkLyFRoZTdt5x49+kuRKMfSv9rqPDY9eu/floEcd4IhB52w5eDgyh5fhJulji
vxH+Fm54MRntOExZ1XJczxjfEi9hV367vaaQHyfT2mMf+PRGkYlOuHYOSAWNoxz4Bd0fwBF8MaU1
wUBVDHI8MsTJBGyu0ibfCkI9xVlh/IFZKyXP08SOmPuMM0x6aI804Z3Roqj2+bt9ZgfvmdTHl0UC
fgZT+xtHh5uHfp81pqPts+gHR1ixVmn1WalqBCt9V7pk9SIbRp/gbS3RMQFP+PwbVPxifF3XxN70
we9KQ6z41VMXLWXZE8QGuZWVd+63GhL2ZpP+6uzo1gtLimQQbxHzVW29U2OaU5ARSdFt8t+lTHXo
d+0kNroiTbqTaBncaMGebcdP8cVASyi+TzR+XN7gMHZ0HgS4TBtHG+PBk12zAlsKuhThxAXlBoMY
P/Gcf/ca42m2Rlgc36cZC1wtsQlUB1avo7DpD/e39I+bprXHS1GuUsZmX7m4yjEe9Ium+5/YfXbX
Re+RelJlbGOTNEvkVf4YVjAQl4J59LAwUhm3eIj55tLdvTeXdrxHtGWiTStaz1zdnZ1tKfi6SOvi
s6ocpy2VlvykpjvbFCoSGvlVSyLGBh16zlGOdmDJ4QDgjUrK0TbTLSVrNOAJzaisLTwkpER0kfiF
l51CPaEddyOI7SruN6Yj8jfomtP9qm67tcd4G/fh2+bM4dFWM1D4tj1HyQfSr5HGO0mBrVqw/1mK
ig7uND5xxk/HrakQwDNVIj/wbSIIcTQK+uUGVzoDhx/rsxabzjudMz1K26rH3oiuoWwBLtNQ2ILL
enTY+0kyzrTuXfYylpXJzUNF8L4IqMYyrcV5CZKPoWYQzEN2Yu7JM/PhcodTml2+jXxKpYIn6Qwt
X1C/V1OZCu/Zmxan/oVzeWIxOkKMvwzC9sCmDyi0dcO7SKKRh75cVIKDUnuRLWdI46S3TEaQOXsU
8bR8c+ZPP0/S8y8HP8JLcp+CHPNGvxDaaDvtiADMk5MUicMwcj/RAryfGCtFEVbimIpcGAokSaM5
oOTBp+SBHd6a16CxTyVvUHTn/Xi7RkKJLJgubPCE87T8/o/vSOvQJJVkc0XUf/x9P9H4Y/iQEj7G
2G/51qMjjqRaMex1n1xPOHGWLbhyfYifWjoBtY5H7Y9l06CFJc+ItbIU0GevjlJpjn8GPpKcBHVA
Ut3Ue/uR2DoTh8VICnN0ojBvi+WUjAgH4Ri+0bDSyZqRshwbqfxo5zl8M0lOEY2GWVYnI+M6Aj4z
J5zcYpTnQmAlMx2S+lAG1PtafbPRZZ3+FUAXBS9eEvclqO6OMV2Jvk+EnAzhMQQhjyAExBTXUpO0
pBfpo/t97nDOMnPorHXqrWnIKTUZ1/8CJBFUYy2/hu3l3gVvuQD22z6XoWzIvPXSczk8T+i+i2aZ
Mm8aQOj1LPFjf8mq+jwoapcF+jRiHcmIHtcD218e/KA6zUjVlhiqYoFW737B7XxSJNQZKlPcABpO
S+olnKPR2PAIOHKDgbrvP/JS6KYEO9j99HC8shXEQxc9YooMT5fVRpPfrNwGR+dFDKs/f+CuMz2R
Awv+v9J4lOL0ZG9ZYWVyW+bDRecaxwHHLlZ5JCysBb1Xd28bbp69jHcOfvgZVclgZoxcsDxFO2JD
jAPkq+n96oGo6rLYx5nXtHPAKCauvSJC203Jkg5RwlBc4Q7c75xCKNjoi4mENXmqYBvF4PEL1+Qr
l5bW4RroU6cI4drhNwMpcT8AdaA5MKZPHtFkzNv0EhVdP4oWv/Ozix/d6fHw2uvvCouAMZFPmduZ
6L3vQSmyLo6DwOsZPpdR7YEMF049ZeAaE2GaKoLpc7zYe1HdAzDfRneuzljGChvpreD5a2IB1f64
vMNcZgwV0ikEn33tn5LUf7iBUDgPodnn83WtqUjNTa6g6oFXcLHhegJzgXYBj3ABCHBLofidjuwX
ALX54dCrJV9S4ZDCbKnaikZW3Q7CLelFikycgqP7PwPWdS6Y8/IeuF5iJZot+ebMhhYIniX+yFas
dntdKuLTZhhDafNh2UKBkZWQZNN/n5O7GqUd4SifpcsvUQG1q5o7guUFRCYDgtJeeJgEJiDEHNoZ
cA8LxYlZ2sD+awcTCYuKM4AloQMW2k1cm/Ri0s/7uWf54q9QaZRDwCve3sZw09O0+SLxFUwfhk8n
q9Sy0d8A6y3FKt5yPa5/EwPuVkQ1W/lomj/w6eMjBf3T+qC3fPhw+GdThnVhaflWDCFt4nR5f4Bx
yeEKamd+RIt1alfUjINMMSJRHjzT5FySay9nutAXeErQN9vh0WrziwZD5/39/C9xaX3kEdRBue+X
oFRpR260GPXvggUqNRSMBzsrz2sWxnSSrxc159GatL/I7DFf4QQ/EQuxEPNq4euqMLMgXWUhNtLE
4kTQMeRSAu9JCgzYcm0nmPKzCnGLWYxjC88xURXk8ABN2J4yx7t5lKsKVxQdXI0Yo66amelc94An
M+PBSgmVsNK2HyaZ9hVftdbvhV1tjzKtIrBLEKqjZNuTM5rV5XgSyL2bH+IMIyap7AYuo+qtEi5W
Eaz+TpA5TOti7eVMxvmNpoezS4kFR0yc0ZHirK3zleoDbrATQiDJ9kSCZoA0XO6rAMsypmbyL/k8
ltyry+eLiQ+iJRAcNoNqKKuVbRM2q+ZXep3vUHu4Z5KV/GQql8k9teKnp/MwFnU7Y8BwAvQBlzfN
t92Z77pV+JGKIlEruPSNbUCqGV7yzuk328ExUZ9MqRgXh3/o2L6P7yA7J2p6ZT7w5WR2Af3ONhg4
JJV6Wkbq+TgWbgnFENQ2v5Vi2SjsnNSn4CVtSq5fofjRBWArjfljuKHRRyHzuJ5ZULhyRMUufCbK
s4KeWJ0ilW+eDUuT3q1sdPAQO7OjY7eJANmZo1ED//H89RcOqcsANJ2Gww/np+fcb39vPWmMjL41
e+RK1Cnnu4Y1yPR7zms7U9PX9rFodnAvWn/M/mkwqI5VpO1uKbZ0YljyKHLKSxUQQ1DZJN5Xa5Sy
XklBrYV87sVFvIFV48jC8KZrqZdmAADAFcuEh2xlTAfC5QvxiKvJ4sPnoGN4jvu7WmHuyPUcXwR4
gmZq7Fm6Ycm18DFUITqDzGnit0Mi9+0tkCljznLJ8B2PkFs5MRDsOIplRrlVgtr6DzpmPbbzMFlu
ep5qhd6TVdFBV8jPjoVazdtylERLOUx7F1FDk6T8RTSzOhfVwYeV8cUtpPuGdIPo/qZ562Qj67/7
8kQK9lybXOYs9CPQQzNuloo62XkdG+SSbllHq2m5zVwsUMgAEyyU9uwlWvjJaQH5xvUd9cvScBL8
oFBYx8BUTAMoEzIZNK55WyiLfpSh6r4garq6ZtmpnqpkNkovL6rNDZSWpukY0lXd72GuCj4AwUTw
PmqJd7p+bsc1HNQkwDLViLUUeGpOzFBkD36ujpxxANUxTSPISBluVcH10wkyHInNoE2+ntVH6tZg
ocN/QIeHC88Apqa/ZLmIkTx5LCYndLIl23AaFAuhN38k9f8zhbz1Y8/tF0rpy2qQD71ef6jW2kpz
Z7ASirJJeCgvQMo6WE0EJD2sFUCheci1bd1qrcSIUrxLSUhOqCmc83RM+WZShQQG+nsPvMp1Bimf
3KsnXcmyI4NzWLtacvsV1lPCx66Va9wByGYmgp+hHWkKMdTDn3VNax//JP0KIiw6fW2EyMB4hEuY
Zd/EMqtRYlp0ZRvRb3qCKsS/3jWud7girHnUB55EFV9UDD6edvUnIM0JOqyCGETehTXhNYqxK2Z8
6+s5DM0s+9eS/2K9JlOIlqmcIRnu7NkvLqq7W+tehMLd5yG4IBzqiyySI48KvVhbeSK7QoN/4MgS
n7QRPx+ZzSJFAtOIlMcN62BStGLph5VtuWdw4/4rvRX2dw2SYxqr3f8p3fa1rYCQqTQVaFHYK1xK
XrXtDGFUnVDPwEnJDg/OQO9g7tQvNx33qlZ6D7uTFcZlMK08mMQe6fSaS5avzJpsrDnATFZsTRVX
4NSRVSnZesObydyWb844O+dSAnGqQUiCV+RTayTiTEprALYu7U8RMcEarCT5ZFbJvA5kmglqOccf
ZCezyaEjjHZ3vwR4VoszrKBjVoKmxVas2FWo1umzZT4lUiEMa/DIKzju0WhewA/WmUO/2XuskZk0
KoEnr+Nz1uc3z+BbWc8aHFZKF/rIiRF6bErKFNrbjNPV8tdUwEJdRj1OOSJ+v+ZGZcSfe8xEM/9n
UjKAvX1ZSYWzvOCu4bGKpV7ZDVtblY5RjyN0DBWJzdzcBYOe4bjJ1mBeJvM/pTCSiwFcXzWblEDi
WDk3V8wzW4d8FXJOk/CUlBavu906VOTvbqbpDrvxBn9DN4W04J9kSiQ90mW7pio4mfRuAchphwkb
fJPYAOziWenImGznH3/6J+qbTGMeOP8lkgdWRlLVeuaSXqvyYagA6+vtv4ceS92gbakj9QtSr0F5
EMuAoM0cMWWY01mu+cyYdCwT24H0k+fZWe7LqDHPgOs8JIuJvyaWERZGeBllYCXJPQs1gDcTdJOk
QpsiKYb4S1Uti+7ChTHEuQFWcy7n7RzzZFWqw01DMus8iYPx3/UnTTOlw3B3bgyy/rpm2pD7+ESx
tUZGPXUArFZFF1gbGdlWLeX9Oc6AboUdWJnKNiFykaW5hrKZbsm2z4GWZIJLzQoa09zC0dZMFTk2
DvG/RPXYRoe8td/YvtSFKQk+3ULP8vP4laXfbtvCqXiwByvrRtbelfOF1/lNfnpUGFki6xr58Tmx
IjggIK02dflhpc0640721lsPzFF/gTiycHf6EgJzrjqEV8qderRl7RuOTG8j37bl7paZI1E3rdOg
Xw9+N66nfv5zN6IdW6vKzs5hCCV3MxY6Kq9D1NP95yZmwAyeuxYjl+9ZlMTMDzTVajc58vNmY6SS
8lYPLxE7Kn1xOLY0lPKZZsGyOJDQKdize6YGqe7nNiegzozBu+HkdNs3pxuJZS8McjcgKq3xLybR
qxoAzxxeX5NRV3zrPyakR5ReSkEfAAXSZbyqZmrw5FT3VDMPjzJjJEaQslrwjPxNCEFEnOo+Qi6w
pNiXCrXs7FI+Q/TPEzXkSD66Q8J6QMvU2n8L90jD1vkmPeRpfzGTjV0MQ5Zqr7+bJJ4MsTVd8G2q
3J+to04B/xd7TWAbRuaHWWYaruvJXksc2BZ/svqPtlOVNimX36CHtY/cdGNDaYuc76iFvCFFENr/
pHXWlWv0EdevGJhvcokDkjit6+DDdwSox6q0V4o6MnjOGkqinJlfjUYfWwjujaokbxEMAEfwGuwN
ErdMKqiaRM8u2Sj3hKttFBYEptiTbhgbuwdUMR7nLsol7rbE8mk0YMEE5muPvaTU2D15Zs2izm/Q
4pdZ/kEOlEnN0cKz/DY8yqPi39SstMKQ+ID6fqtvPHlUdtwaquCGd8Kpa9iXhFzlvAiWFfB5c4vH
mseZXNLhee0RERDALhUPMVAoE9NtH4zlgcm11/juSTMychhMP3UapzHo7Jbu4vZuXwjqzk7WVU7R
OdjBCpsQlGQ4dbzoKh2vHgMkz3GkAiKPo8+q6OZJyoWyvmgjnWAYx2xWrkTLwRYZwa2aJnINVH6c
OkZ0KN6b2uVXpd4C9ssW0b4wUTlvOk1PFiSz16xyksWuXbEF9G5GtYDb6KMD/PyfpCZuvIP3pWTd
+Ot8kppZR58LZFTTueCkSBAHdLXVFkWLhW23L6NrFFOSR3X2yLES/6wQjXDIWVee5EehyMCdrwwB
mMunN8gqqjCSG3TDLoWaNJk4n9/+kSGsFBMb+Itqyoowtqaf775w8smHaKoEEqjRBYAvX/kQJNG8
3nfO39NDM9xEbop4hyYCqSfSAkEJ7URfsHAwlES7usW/cgVARuVvRnNz6jw2Ehdo4NHRASPJDGEw
oKOgfUjIDglhv6DmgZ848Qvy4VXF+kdQHBH5+mnmjT8JL3vNApuwlk6rfarWeq4GqvRcnlpYusJ6
68R62Vfgdp+ujNLINop5VmXywzeaOEtXFqg8sQfA4KZqABe9bJ1htfEyuviX6PY+aXUxhxE7lZMQ
SGJU2fREeBvyL22b8UMO46ThhtJU3AbxcU+MxbwjTXtJ/mzKTlXKMl7ps5+F6FJdY0ARK4KGCfU9
X2t0yVdStm7Cn+m7F/IzOvTDssJnjmZMKTJzZYvAGM279zCtK5YB4THbrjlPSvoeQ8qXmQaq/yMJ
TsN0KArZH7ujjDV9Bhchy81W6wZ1ypauUUXxnFhB/WoB7IK0ADRBz3ZuM/ZaMMfaiu6Wcffd3FaP
1CJs/okGszbJAa7CyiI3gAY8kQW+65lRlGaJ4odi8EylTdG49qt8SzyOIcJOGkQiPYK2J0XW1OIn
g35c+u/DMjXtXKhYdDiKkcQR6KxJLZvr1w/vaUtv3WUE3zx2S41wEmwjAGcO3NoaIzAU38DXAUt1
RJrOimi6fkZQGvBk5esko80wKJoz0+D/8M+Kp+zfX0SyiCuCTh5cw1tLpS4PebjwNQBtpwmsoMlA
UpcYoPgaPvvrmCJ/weFxvIe3XJkIwX0YtyM4ZeCrTbzmabkQPEFG/S/g0LjdmuFCT08PcfJ52PsA
djLLPcVYnKy00YVoBZjNcdQbD00xff5XUDHoUNpCL+5i6SKNR8Ju0UkuwOfyUVwQjzYcOpDninxF
jE/iGgADM75c+gVvV0ND32wq5ehCg7/k9tT0s80+yQbdjdSZ6NMjaZGgM7GtD/Xw2IB8tCyXrdz+
A6+0YfKLrXcvLm+Dpe/tSyGfPO4+O+FQH9jTFDtxXg/cWv0S1r3LJDXZYVVqKV527WGV+kR8RPPs
urCqwAMh76QPTXCnc+D+SUtbJZVVsVYz8I7j5ZYAfpcY+Pk1AoNTsI7cwvgyHvh782dvkg1PN5Wg
CoW8tCDsl5Ih4fPubEI74cZdTSelcdeOeafh1UocgI50QCF3oQyXazE+O9bM/1E1ZtkFPkBrqcQl
n9flzEp/qPxJwaJjAtT6nqNbfeWaL1gvD5Zg80L77WHbdGdRmxSXzVbDrA2s53NEtH4Xiziwadhu
KR/5n9sg0nhPkq/zyQO5wOdgUc3yMIt6hVy3d9k7UF+eOxkA1iBDIwqalv3en9fubPhdDjcJGJz4
GD9uXrykfumORGHn8RujrD+ctP2MZj1ojlFv2EeJtV6XRme7R6+0/Q23GMdplEllenXoQrmHoKyd
ATnzhUiYn3eFc58qgX99vOw1PboQqbnOc+Ri/pF1STlFC66+Q5feU+LFNP2jmL1NVrr7JtuL/pVG
BXF4XdrgZQuN3V80SRXu2TBwKTbuvpdNCJBDH9Ao35dcBeWncUOb0YQtgyy4wGOX96EPKXnuzUDF
gWL029nEPDYvgUt/kn19Zv0mcHN5WcgzsBiq3RaBly46aoBrTiVO/WCGdsjHeLkGRnlQurnG3QsX
OLNr0Y2wVefjV167jDDisJgd2q4ZchaGqWxVeYmdWc97r3qfp/Gt9UCcF2svkjsmyGFzlE4EeEou
wzcgtLhWo8rcNxYw6iSSQcHnIe5en9lpV2Vvv/+ZXmkrfwujP4I+zXk2PP2ETY/qcgaSvrj/hnjM
gczte/Ci94MqPW97Zmxv7J0P6kRWk/md0OGG9OOA4HnhH9qjhFZMz9iDGXb/yB8z2zJ2576dCtTj
kKWPKrYcU/3J9BiWawoUtHisGptczVlsWja9gHmudxRs9Lq6OL+YrSDyYvLtaag2GVJBTb7ZJKHL
obPyxSbe4DjnbgjWd0g2p7PdkX43xCAxNB+g+SUQkbtQ7PJWqybpK/LTDAzW9NxSYuHBIpywuF6X
rKhLIq3IPeuBy/IG3vN+KKpb9xR4n0LS9pk50hMW+phQo1LnQ2P3UZxe63RsU3F8opBxWQCiHKBw
uI97iLGOWmCBgtG+O0FxE1ey5um1rftNfjobrXIelJRttBcGi2rYnDjNSx8V5LAuRdFvaBo7MvA7
+Tw4oGufUqFNZx+uOS29UFoaZO4jkG1AxB1e76Ugz/Svy3zMtKJzSon72OVezxcnDEGV9r1Gy2gw
C1hz7cYl9AZdU033c0wJWkNub4x+jZ+0+PqUz1egK9fajJoeYZjxOVKahqUCHVb9ysyyR42nOeiB
BxNCfgtd75ZQ0W5qWAheQDMsJLHAifYCMpQrslhs0j7nfrcLxKTjz3zH4MiVxb/ZKX3TVwxSBZpx
Qn1zvVDGFOaXX2MhuEnHpIEBVto2a+uPtTlZELR88kB294xaTzPiYQxwqod1dzKPvu7A1ti+QmtJ
KxveHmsR+pjM+fw+HesA59VP4Gdg9z8o1gtuRBk5GDGhjVcOue9Tf7d7zIso2l45JGLFm5DaeRyb
uBHeFfBEPu1w46ueLz0XcCCPyF34tAghcjst+DRPmnChz5Ux7shZ3og/FLpP0u5rFv14S9VkCmqo
7920apDXYM+DNq15uigkhQnB0wc/soO/+xk4M04nFMPsHkbvgh/xCIgLKeJPZPmV/6qLguEIkGi9
Eae6rKMq8kLudzqIXaXukjs5oAgws0gdTBVftYJB43oDr5d/fWdb8QYLORlTDnTx2Kl/SmHLQ+BS
NLSqnJHnAmv/0aHnxyC4g/FSHtfxtT0BXrcuvUJxHzX9dj+gyBOwmayuxLjXcTgXL3RzNqiGk+Ij
oCVsTS/H4HgtWQ8unPKF2yIHF2JNgWLLqZ3SjtRZv11K7v5eUscR83e72vxQfH5DBA7DyP0930a/
19dIpTmec5fohnUTDVD+qQIf3cQdtrhDdm2hEic3+W1M1qmyNl+PY0o6ldwAPHDFuzjTSfN+l/sV
yISowVj9xdWal9MLrFdCKr+ZEBuqwHE63ORA5ztZmkPosmsr5HRxkQ4V7ZSGUlZHWcZTPK+sCXH3
UiJBU9odOIy+QfNGCM8LtTTtdEi/E1rrOF0yAMHz6AFPeq9l5d3tkR+09JIydS5H7gfMVw3/IIbz
9oChn4Q3Pny+fFpVqX3UMPpYM/m0GsJZQZd7PCxG7+YN0GHnbEftOuY1X/E6OUuZX3wmNO2jGvLZ
POFW3ah1AgjFWYKm64VTwQMKAlPIo/WOVAP4hpGTZoCXGqF0te8HOtDvv13QHlyFWoMcfG4WL8UH
dZyvT69GMtKJB52qD5DVC4BuWoTo6RwF8jN0Jn5UWbQASTjutBpnpAq5Cpb66bSZxVlT1EzbawFC
u/6TT9BNZxrDB0JEKj0CjmRJIWWpRVDgo5HgUumOfDRzAkJ5Kc2OEKeYR/nZ4hZtBQQ3EIrQqjni
D+QMB0WYDdoxW5hSSXo4x2Pr8T4VnTiE1XT1BqKY6hCEwNq1O77gtmSY5d02yKS4GCToS8O+lwKC
7yKk8EgtB3L17M0IOZ9YgaXgSQ5yha66uc1LoYBMprtej18yP3/XOJHxrjCmhNvb4PMdU5bwFPh5
wF9BkdIzGuEL6/HjZEEAZZTu1RwXrYjpgJBTBgaLApv//mnD4v5nCanCO13yMo33dwRcyD21hIyp
kbklysRrrkW3YCy0OXgpGKDxRmr2A9OGkcXTSuv3+G9gcJh841ErlTshzV59Xn9Q2bN2uSW86CWT
4VIHZvN1BIy7/4lWRqz8giuHKaPZv1Emm4H0f2pgKVyiYc0z365arEeW3KXBMqN3qekEsOElPkSc
NOxO/lLQOmPApP5TOmaEKstihc+8ujjAH9J2no41Nr+s2QdTYNzaatN6HoiqbgBzuf4CR7sSGzAW
ZP7iD0Y6i2sQPdIrdkyZTgAp1kI1b5Vg/49sUC/m3BqAljUOsKUVvaHnOazQ1mpX6RPgoKHchTVY
b8uEdDfqUjWCu2p/svV/hP/BLung5sPaXdgdBewJY4xgEgDh1bODGwuYrB3MpqDxWVczx1+yfCG5
n6yuEVxfsl0snMXh6wj5+6rCKWWR9DIVsGtWs++ZrxAcqBgn5L2eRD6svtK76ekUYX3NKno2l9GU
UNYX5xdmnlxGOl3V2tGwsavW2YZV28G4GdtgUmxfYDm1BYW7OOOlPiynQCjyFscgZH0WqO2V+eHm
bRZNwteLyJsleyXW60cICASyK9G9x5x7tcaX1PGppDQqxzFn9Gxru8fmD2AmXvlwCGKNQSzDT3VK
CWA64zejOhyv1indys2pfIZPE37pkAhoCaUbu3Xm7zlwSzclErCcniK3w3QEmj9qwexhLggfpobk
JqRRKQpDoGfV5SuJxwpgiSXH6dQA44JYEgNo2JcVZDVAnaOiDTMYGgMz0kL2Uso/yE0Ef4MlUy0t
EJTK86HD/gQaMk/v9KTdoFvcqLDj2M0OiBdlpcjLgg/bz1yx30n4sZX5e6ZRPG2tcP7bKvqpzIUM
NxamYwK5qQGk1pvBfyZKibg3ESWltsuLNR6VNN3QQZUL4hVviKn/mehqB6U7pBfp+QtIIDhUn/Qq
pa9clJD9y3hCxOlzwsd0pogOGvguGn8Wzi/2uhlII6uqPBnkvr1O0j4eJz+ZnVYWjmWp9VbOUzxW
cn7WqD0XBgNaaktkPFsYtFrSeqWY/Yx9P9BqUA74iOCO6uE9wMJ8bjtITFvWNsTdJ+aT+UcHf70P
jx16CEz5lRLkTT5lAg+KCtqmK6Ms5N5I/JXvJ5ehBMq2CPDsGn1J/6LYXoHlWGuaB8aMpdreon/a
HFoZz6tx36AonmDmBgifsFQYAsbaaf0Mv35MFfZiO0wMhkHC6/or0IV6vtYUkwhOuFb1vTPwEr/a
wp0Pph8x/mEa5emKbAELSabL3oL7jDGCEARpcsU/LrfmTZRepFlVmq2UgYKH59PCz461rGlHw5Ma
+f7ZSR189kYX1vvN+bsbK7qXoK3IYx+6dOueaYtH7gLxsZq5J2IqDrn/WZOk0Ngcqsn+8S/LbZfC
CSUxm8yHUq1BO6lrxsbWz9InWnu1CZ6QZ0l0KVYji8G7bxasCyC6rd3GOVdqwOezuyXRvmf11S8m
LRIlIDpES0FfZqXfNxesA+D7UJo5U59MKsLN7eBT3EM1+OKyJ7iEvKT1x7lzYCY4Kl7BGQ1fNP/G
z28+y9lxgWAC56pSuXbE1xbtrOV20t9oJWBEBDO5aBUsYYG+e8Myxx+ckcPpqyIrsj+P13Q+MYf+
d43DSfYX8cWrauBG0+D4SNKOzZ6Y2NByD4dsnc9h8xJ//z4aEWKQGSSvjj4JdSaV59rXlU0T1c1T
3nqCEdHODrMRmkFuH/hp+fspVqfOEonZgYfBG78pUaPSCXhYqEqOslfP116T2dCRWfnz+0/6lABS
CxlW1nuhawP2Bqv21RpklfiYtbMkgeiBst189GSmPUqV0IehfeYtAQS013LbVj81yFpl4hSfjL2b
8k4nNpbkKMAhIdwdegtcjLs0nzhPdhQeOp7sBt9XUcbv9PTTMCqo2ra8ihtrxsgmw7IIhd/BlkVk
mVyFb7w4l5eDvH6KUUuvAR90y72EZvAopHhRefHs+HNwrnfwV1ny6/0BznSHjc+bTGYZ+Kw217Tu
m32ndIEgolovnuAlA5Rt4U9a2BWDwoWMIrGNgRjz56GXgb7Mu6hzWdlXzvfh4MWfAZjasvlTwVPX
y8ZH2z5bGceomqcwM0GNcPBhZpJ1NkMdp2dFZYiK68SdHHGXkhX4l4BSQ7N+22T5+5Pssehggn65
MXFaQPuCLF+LwB3ThufrwQxnBtw3NZynsgJNu4jfBepfP2yn70yiGotgUhXVq4FkqASv7HqhpVPx
tHuZAXdBmomqbuAmIeY7dzOpSbEBX7zmOKjsvGM1U54rMfIB874Reyzq6dYLs0E4+KkTaJEb77n3
lVatUD15RbPrRaE/NcwrUMzpLTS3TWr1xQBEPzBEh/szjtlbjhUTZmVNQEEEMnsU/dA5Zyf2KZd1
lFvA7IHo0Pof9aeUq+K84CJ+29dK2fobOSEVNaWNR88p1GcAhPqlDFd6uQH5F7IN+/LXlJTQ3M2e
Hd6MDiyoRq1M5jJhnDV0CUPyI4/iS7CBoaPct430WttjU1EfqZloUPGcuykQXEuzgQbNyUAlcblz
aRxPu5w2yvyzLohpRD6gSZemwqwWLCXLRWUEiHd6L5Sg253dppYw233bigXL6qHVRf27XxOKIc0Z
T1reHVOHd0/ZBvsdz4sbLKXLxZHhHwB+uv3eBFjiKtMYoSXfozw8JY68rx6+y3tl/7K8UMabhuQb
sttQesfocklgAOO1hvgZ98doGzjcMBq95SYPbFNPo3KYvuuPkMHCMotEINI8LmMMyKXzSv9nMk73
sD91lNWASiSiSQD1NXrh2oMeLygZsL2lVgMiskKBGPhqnNTKSJe8ophPaqtj6IIv5oN1mP9+sSdD
j5NJ4nqjrK5rSIMLlptbzTVBVMluLldLOiGXZcKDxHvGUEzelRwiqpjyLlTzyL4urSFvkYWJJvK3
Xp8sw3LIyhv7GTYKbLiVTs2VBwyikl7bMvODJhbwMYtbc+ROCc3rzDU/YNqZp/SlqzC8rGuNRx8l
UDwDnJYrDGOLeBZfNhuta6xSJVwhrtADVQ2E0OMqu/XkVJlveo+m2lfdxsZajB5EusgncMfffRoG
ehYp2pS3ggoLmYB2UBbY6l6cZSgSCdsp3RSr3TeBO8KkYn30AMI61GI4ctVMo6Tpt0Q272plLLEk
u0+RmKBvXUTQnq6TP9Q50SSr/KJWC79wlsgwg8eHm8GQsUj5yueF6T0vpUy3+jNB6tvGPrIjNDio
qteOKj06+C7JRIhg7JDDCez50jQ88cynYFeasqb6e2tiH8YxQNkAan5Iqz+kDd7vyuScawwPbAFI
XEB8DCTYvyV7ymsAQemkVAIKKnnTahbA2RvGTFo0jVwx9D/nhrRUMZD8BHiZ+6MMruI12zUkmopR
MLL3bD3jqWw59IcEirgT7E5BrU90yMC1CxRqorpUImSabffUekM0ZO90XUIA6azfXJgzWITU1eHA
crsS1Xr+W/pPbEmrKhuW4J2ITf/pTejmKIwT7vsWsqeI3RPZskyttdRYH6V6YZNAO02RHG3lAQlK
cWlwQKtqwd83yMW1A2N7wKdy84lIP0QjYHnT+NfehULjS4Org2P4ay1t96F5+vFaUWo7epD2Lbok
++CdhzE4pU4XBVZJrsrYnMiu/9IIcjx9iSHWYQ0xDJYJAuzkba5d8XCfszwInMTPRfS43D1p2E7w
liAetyOEucdlk5mPGjeJIWuUXpgSHfLzNxfe3JTaK9J2aDiU7P5+QOrBwvVfdTdlVOKa1sy5+A0R
5UzAHJgG7ZdGZcgpzBoQQrIOdx+0Ei7Vuh/mX4lHIjQes6WuFv1Znh8uBlWySdZBpM9yPlgAHFkd
HUXgw4At8NaNPu7F3iJqxindO1weDUrPpj1bxudiCCe6XlSQmOCkiFRcD0yGIkN45BjxwV2AJzOv
oM27F3wPUHj7hmAGZubx2yX9Qki23h8ff+eiBmoWa+JMjmTZYL7Y1ARx0nIXf2eFJlEeqReYGQ1p
tHsYvETKvAJadi9x2iwd9wkHaPZCN5Yg5R822jJoZNLr/g9XBZVAVFYEdAzpM8xS1cg2CZHdSdt8
1NCxfLK3aLIYHaoq7MPEIKtbfl0p6hTfZ4s3lQVFlz4WFkVg9vDoZHTnfkp8Cta7zcztLtxumPOU
esSFz5O4bBGtQk4WQs4tTd6xhjpsNDH0MV6rqb6Ma4eaglkyZIy32zTOUq3jH31bai4aVJHvtREN
EbBGahLrmM3EpEu1mPmoa17Ikl+Ri7UF3iesQsvVsz5XQO4b6qYV3EA42F/JYLxIJtBWmhduprF2
bG6a6RipaAeb4UBhF6IPhQHnhy7wI8FGCYmdfrtosODzrZZOH09j4jXNaDIhTnSp56BCrnP0kIJP
k6QhvyPralWRqJO7mbkFAyKL5UFyqVxrWOKCufFieAaD4dz9TvGumUmYbniOBfWODx98u95Yne3z
uukNZTi5Md4Vp4dcxgu8W1osHIpvInolARdi2cg5ptnGTBlh+WRvD9h14UK/5LLEuxe4I0GN+XZ9
m5JII/chEnFs6Cxa8dKs5iSH7CqEGG5j295h+LBuFjA4YzVTcd8Oz6TOAtmNB5+kO2iWpHMYgp8m
YwFtAL0nQdG0yx6PzSZEhuuWtRPaA5cbSvNeHSw9SGUGYfvBfkSGb21EX0HBeA4MuLn5GwSucY6b
bzaDWhOsviu7l2BVpNDPSk8oVGqE3aOIvoPGfasWXFypaRoiSrMTM+ERjWPp5rx4EYSqRDxy0xew
ZCilsfs4bgXPaMnHVFOIqhL7871nkjmc6Kpxaqlt8ZYTjOx90YGTm2JWIRDrXBCbiZNFMWkKaqYY
vHrHFPFR8ogV3137blrsST/tys2oqgq1Lh6R/viS2j6ZWND0d7jxC/7er/Bvy6c0lKitbZld+eeM
jm4qHioxJwwhkn46je53MaiVJ6sW3VEiYTHDfuAHq48U/LtTnVa+wvJYO+OF+LRKZAywii3eItCv
uUNsobjb081R8rmekxP85pHN0HYJsS2iwREwvJFmpHyHw2T5bYhjeUpQtyC2EBXSw7el4G/BkNfc
PRMOjoCvMXzHrIBrG7/UB0MxPKAZQ9QhZyqXqp1df7rOAplxw35Djig7Fl9MNm2uOuPqiVTRJyEs
qJWeT+b+77yVzbM40HcgTIJTStTcKtMF+Onnyge4DkkQ91rIBweOLDLRXLzzdmS+ctY5IWK+fyN3
zjOLkGu9D/o+p+DtKjTUbHPzDlq2ejlZgpxRT9t/VwSa4wPH9lAF7dN6cNQ7NxFybefq/Zyq7yM/
vC9n3RKJbXlbXEqPhvUziZlsd7xN8YBKUzQGhbctUgUMfcFJdSAoyHW3i5aNBRDSbkcOtSGvrltS
clqyx7A9oCPAlIuZh156+iHoX+3aOjvE7mdEr3DCfhAVWw9CXtl8UtYTjHMo9q37AfXHofRT4S0x
Zd639ooJ77fVgJQ1mz1dfah39Z6iP/CU61Sszi2TTfuZe1VbNlWkE2GrdEwCM1jQ4GhIcEVNIAgP
MtV2BZsSOAS1cAkuvnOu6KFub6usONtEe39ebSf2wQn5K3v2lm42uTq3/0djP5yPETeGQvjgcPW7
vYctsQP6JVhTMWSHZXYFy991W0jGoU61oGbF5v5uqXfg4Y/Q9jbWPaAs/LiBea2k8Ube2fUotCeg
W6s0/pgj/vMcl6HgSp8IovIlPDb0+9bAZ5S0EeGXSq59Wdyqqe9NDE7xsaN2dwrD4NbmomnZNL3B
3WdpCrKvsEWEpKWmQyWk2XaAuy9ATyYJGCbCLdPxx9LzLYQiN+ypkuRjgWnHb4Z5aKUkisw23pgT
rreQbAucV6LyT65CXyjtDzKNmWvnhgIDV+xXqTdiX0I7EJSCUvxdrEhKCR3pbQyt4VQPbgd1gLDh
Gm377t50wOvCmUeZlx2SKPjNn/wCetYxZ6jMFPLzPzOewAyy+LzG1eDl3VqUiqR9GZSV3Yd7bFZq
a1TqUJG/WzE9+RzUhV63u3Hf67S/2xjh3uFangRrUV9B0GSKhuRt6IVLTiImmC48Lc+s34ppNCOo
J9gRmz4VpAxbX1V/5D5Y5horGAIUJ8zTrjK3X9zyLA8/TVzK3yRKFTRNHCln3S+kGzkd7R6oKis5
SMz+VH3+UUYPsyqtQpCWLQLuDmConPQznSAu1SoF5qGY5oZ9OA3Z3LXUmUiL60aCduYCv0sX10Ec
eto+eXJMAsZCFUyZA7Rb6FHqHk6xCO3PrLHnEFu0p0GrycmjqFRJeP5zJsFKEpgqYXgpELpUNwgR
dfpqzjKdx/0kB21PA0Dv5KFKePy38tFl9QKIFjDjEtxPhrRv/rUozEW+YHDhOJbTNgs2Ua7MnS7L
VW1zHDLlbZPaLh/lfwmnflGHqGvGH8eevIeVvyZfalH7G8kWQ4MGYhDdOb8PGyb5OwU1g28yG2ny
xZyph4uY2fr6VeiC6ghZQTIw8z2cLSPyEFz+Hy31B0e/VZULAsFsRbUriIVJBMan3IiBZwl6IjMz
s1xMZRvOcOW1C5dF3Q1KU/1HQjHElF36mMjGAums0irfxu8vM2Swd/amJx9OjUGhqbHL82I2rDJN
bX//Xa2hcQutFGFnlrt8S9Ag//rnqV/pF37RR9VGmfz9Ob1KYQxOcvH3XVR1CYtsvNiHG0kfF+nu
h4iR6lmiG7UwO3p3BWq1zkANCenCnbVMz1bMan14LQVaf8PdjHGX8Lpt+ItAOaJhoKqui/rUhkwO
UwNJpLxzb/Rg9qx5HvU3zwgWmHt19aSE1F9AK2qdv4O9ATEZ7WnIQLfyY5v3MD/jCom9az/LeE39
DwpfIUw1A+auYhQ8CYF35EXGIOjXrFsmtcEseZhwirNL0dXsgBKaNcnlMM2WBnKPTf+yu7PdWeL2
0iVbsrKiqCMgUpufNyWy8HZAPPfpKGBBmtJU8N3BAFUgLICH4IWeMIy1CxUglcdd5dUY75AfgizS
89jHVdRXF+mzr1CW+h+ce3JFzW1qGv7ayM8S1kyS7Bz4QXm8Tb1UB8uHEe1c5wXu+jBctkQl0Taw
62Hi2Uzx8kapKJI8hQDjlr4OXIV6krfPFvDvVE8sRgkH4Zuc0LPL75fA1Gh/MOU2lKOEHXx0EV2E
zGnESvouQDUi+VH8W7yJInm+Y1mGz3LX3ZvJWgDrdjsfT5azknNzu34lrt+CEQBD5joS4o86Txqb
so/E+lksoGin1zDrmh5JsZG7ReRNQ+rnAfE6DpyDbkVUCYSFhA9lwtMJ2wn2VzFP8+5rNiassLAZ
/12chOqHjuyMDB8QZotL8ZHkW7Inax/wTlvG4I7Xn3C3MM2CCFKEW/xDNM8TNgE4FlB50REEa6Es
SUwW7EE5wsEJK/0bF5pHqtJUZDMsgG2DIxeeFxrcR8Mx7rdt71k8R7aZ19BbDStEv4004j6w/gJY
3p4txm1h4/qurQjtWLWBxcsntMYViF0dTz/Nxs9O6sSaqvg1Kpfk9fqxIF0reqAO2oLodPKDvJKz
7LAg9qioyZz967XrSIk7xv7nCp6HeUfli/kc2b74bpZ/2jp0nH2gf1gJMVND1YGVXZldZEvVq8mx
N44adZ/jLXd6PLn5G5mo4j/UrlNoiCpSqMpjVgNqhERYy/MF1vjXibJLpKL3u0xY5cLqox2LEPbp
zVL/DsOZKo5lBoa9U3Te/ZbV3XFl0hK3th8R7AjAr5B58gNTDWXD2Lcq6xoTBiSl/K5mZobCoJrG
9ulqG95pQNfTxSNmHxY0Sgvo+Nj9XcHl/enN0hAJnrdNURZ7xoH2idbahMRGI/k1aqyxqefxFKAO
bszS2Zx1xqN/UGU02CrzV4UwspylzllMtPEKfJHOu9red1nxhNs7I+8ETulgvemL0zNR4GA6OSM8
gOeca1qtaJ2f01hiKknrKKxiSZm+NmVRgb0E6lRpMlVw7KzrIxKNqn6goyCw7WAnemyLGT1v1Ejp
Q69O61usp3DK/SgNC+P+ebdrxfBUy53hXdKFukpXUo3H97du17ykRR29jn0lAjxnaxMfBMP4mFUk
B8EBODqCYOy6BynPIG21e6QC4E7HZhWsBoIIxTp1kd0cjomU9nTlEWU79iIQ8Z9MSkWy3BkBab1X
DJaZbTjBmmhMaca5a6TB4g9OPA2fh72eIYGXN9YAp/XHLxqCNbrByfnTk/NuL85ooxLSRpp3vzIu
rJqLVHP8AR5hzLCSUNNeVGq/TlR/aOnxEDnZFkn8h1ZaUv5X2TxK7duv7FxsVebfnVPeDWIwQ/3h
wfek6LH0mARHHQASkrqh0eU6Ml/e7us+hBN12WQ41JJcLat22TGeADr4johLZwwmLM4p1xd0rrja
F0omUxLlakY3B4RSHKK3A4UsnxJCj5mCZB8d8rbN0X04pU5bZk0CaNYXLY4IjqKeU0LnPnqvfU0x
RnvmvpD+mFsSIYFDMe8jPgs3mZrXKG0rPSuZo+KyYFV1s0mS7NlXDIzZd+PzpPoz6Y/lN4iIvnpj
bGi7QF7wsVZx3adWF0nHcAMBuIxXL5p4etpiTaqrM7L/50uHzGmv5dMG5HByYxC1eXL5ht8012gU
7fJsp+wzCJmdiyUf70Ss+VuuQq4mtotXx7n/MLhJMrli/EqrXkSMhM1uLb29k/zJMUYZtyVbxNhW
sfSESu6Sykv1c97LqbRxR0XUBnwqEOurfDZlI6YaDJSndOuyR1GarYsfr/hu9i3njUkKLQ9/3KvH
L+WIUfkYgbibh512FBaIzSsBQ0SCy9r9aDd3sC4xHEQ8y8vBTN2pnENNJy6BhFuBT8VQsQwOpFs2
P3HM2oKCGvus36Sr8y3+LSbUCKns5mPS/iBhxWXGbPuqthXE69+G1TaqQowLXaX2lUJC9Q2MgE8M
AdQMkpMCmriWyh5lDvYC4GcHugFQYohj9UeJ2PmOoZg4IOteI4aNQD6bmFoyyi23PXJwfYai3GIL
fAUeiWu8t/I5eTmpIy5bV0V8CnX6o04RwXBjYxkqmZWaRCBx1u6aymXDp6heTOX+y4sg91UcCW0d
XX1iHmmyIW7Ol0shhXzCX/r8+K4+03fbO8YRfAlh8EwAt0MC81oAYlaz0CNU5fgiOwR9AciI9RpD
QLsFNVbpZ9D/XanJaaV8bEybyt8oH6U3K+g1rbNnUOjtmGjdWZeWauHgYbVIBL2/yDM+oWOJy5qN
OmDj5ZqqR2JFYO03PAKQx+V9xO+6mrdfYhuF1fXVOf7iuJq93iMXZ3n0fyBzm42lrxV8Jz/+5zUq
5ZlawVwq9/inOE8yDnQ/k5GMrzl+1FGlUMA5PpQu4r5PSOON6pm4SnemM6MlmQSq2bEjzlAOvwh3
B4ODl54hJ+bybxMGYN1BQVEpiA0gNeWo4sUpX2m7e129D/NDefTauMw9WWZbHAlbPxxTqi7S+wlI
g6nhFJp0kdXjOJLq/b4Gwk7roIhsDpEtA3WWTCAJgmHOd3TVeuO56wvbdsVg2+d/yfL0g0OCLNoj
ZI5uyQsAfps0cV2G3XXquY0t0vlFTN/fLD/6pwx9jmeN5C8IHQ8HG8IQwP1TIoY3yg0sFpsl63qb
eWeXkrDr8mh4KIcUz+UhQhGV1cD5ErS+mF5q4QWh8kECIinGbs+uZpKt5/vccIHl8msMKu4uDj9h
Q5W6yWvVZ53Gn7jEuvbezi0Nmj30XZXnGaz0492OfAisseTOrh+Z8bYcsX5Z1bM8op5BtGFCeSnk
QEbRVXbe+FOH5bdCCSrN50/nwG6iFOUuSE1YPXnsfDTBw9+7mwp1mUOqxZ7zXghD1Pt7oq84XP4j
Cf1aNZ/s9fLbhRO3QpQijdmJd/DxSVM7QjhY5WWNDMb7C5y36kDkkU4KrpaXqhoyz3RqtdVQTfAI
KwPEscP/XRY/ccRquwg3AkzSeC2OUPjKLjDA6cJSCH0ZuExPnQlO31cIP12v9LqkcDC7RS9daOlV
/8oJm00tpjTIWo+tgTOqa85LMO/6HXdnUZQWJ5C8/nzEGRlrSdWMtkYGwAo3pPnDMvJEUucit2Yg
4+BFdUslBp9ZWThgInnZ5vtFq3lI6B0gJHPJ/ZFKldKgyxzSV4yFQg7bvz5Bcq3hzSiA9jIpBSQb
I529QG0tcJQ2QBGpibuEGbsijRvgqNoBiPZR6wq+s7mU3fglBxqOuq3+u342kVpzK2vWaFJb5izk
belm0YQyyQWlKOjOO3MlhO9zVCdL3EQNfpJPfd+kD6xp8+2v8W2vGWa44WpDuvDGH8tEefJ65p+2
BCe7gr5DrxNQPaDLU+T4Rq+zN3KM8yAkIylzCyTBMuwCAfy500dLaSGi3R3x+KnLW3gYcR6dVS1O
uHB4mWZ3Bw51x1Jh8mp+XIh2kHqcveyxs9yGos4/E9ZyimKWWgXt7D+3mp3oa2QCzPMo7dEggGiA
LGWRYoMv1AQty5RLCE+S/UyDyy+xY6jUoHNr8wO692X7XHHHNFdGe+sg629tDXrn8ICkRakhhFji
Pvx1OHOnRyVOleMWw11cLQ1D+qsXWv8qYjSvMT9/jIYyc8lhDelGZYgYV42rlC2E2Uwi2qNY98wJ
i796QgnMYDN7sJn7QgNGLW7ERE8d3+f+zkXaNs1IB5RyOpGUIQHW+tAGFtYQFxLfifTZEbKDy7Nw
d4mYnWE2+yVYilU78UdHKqsJhAFHXZ5HMbFZBzRyFtnlcF4BA6eZzZgmilTP/F3X+joFdaF6kr3o
K4Q4u1PwtPJ8l+aV5Sw2Tpw2QwETn9INljBIZE9jFObDxEz8okWMVs5dB89tqAOgSTWgYUbVOdQ+
oDNYQs5o332u/wf20WcM6nqbXTPd4eRna476clQEUkSH6gVXR/fLucuQperGO4f8ExoC401DVXjN
Ska252bTz8sjVCqWXswRzKCbKu7QVEI23yJpzOeRxZ5ImxgVQkKan5W8aMLZh4cCn1p8/ka3tNQT
pJvI/hg8SIPeMrqecOnJS3wynrasqcZsrdgUdjyMON/dSkNjpR/2dHgK0kKsswwGbnbratTeOe1U
fNrXR3FL+c4ZgXzWi33ilGeaXiDWtfX+KjEn+xIL+ByqfelNPIoYf6xkJcRl57O25R/ftCuT+fYz
9sSBFOlYhEY0/XgNlxoLRC7rdQSG9cCVFLtmm91YE86tSTOXi2oaN/pk78Mky7evgpzXee1QpBd7
+K1L7BNRi5nxf4QhnIRcf0zWhCG7ycwnLHG5O3Xd7KwwLIW05m9QEmXb0qIlE52bawoLShwIU+33
e3SumODpzbwgyWFsglIg+d3lYNoKQ2yRSgViRhwHR/ia2l1w0mawHH5NzK8a/FlK4fLLl7YwXhGY
9I68wFFvtQmWE8XtbdKn6kB11WMdo9PkytgFOlM7YZHYumqMfmYrGq9usjcj3BqOPs353rJuQpNq
tx1Z84e1JX50SXJEe3l8UQG497Vzr2tsB04FWp3+gfLyYdRTDYXcwe6kSVOJcRxCm8/X5imnjS4x
pY9DMctpfTdFs4uLN7bDtccrITuE7Eh1knYbaWl23814Z3ThtdlNvwhOH8qaLur3qQjoTOwAysHB
DpwWjGldT5bm8BnAeoDHJg2VW7mh5+0+bNNtvRKT5zGMz3JDHB+0jkAEKlsgw2Z1Om5gsU5ad0HW
5VyIOn3s3du0yv/rxxwVfyvrhqkMXuoQ76pkWFrXdQBO9KQC8Aj3eVcxMl0/kg1VVO9jx1L/C9r4
kHPilNchnvcJeZttkYqth3bXr9h9ZFzFP9tU2+K48Q+w2f7pNrhUsvGxk7p50mgAC8iCQ02KwkdV
Zf9ikW0Lw7bW6GHIpJRq8XiDky+sJWhq9rNI217l1uOQLWqPWnSmPho5KOkYMWCgHSS8uKw8hpMV
qu/yOPKr6pVj4wPOQfnSeSteGBQyoQoC1/di7RDFEltExRe0rqHqwv3btv6F22yxicRGaxV10w7W
Zp+1JsV5i33d9Oh/lTTYx6fxok6jrduZTs7ZuPCb+avTmtZwA6alCdkwSwkTnRP8YA+fP3Or1Q5r
Egco88NWLm+her3pdrMoMc1jG7MRpR4bGYyRhNoAbT8U7VauTg8HIsWlpVg747F3BSGeQkPfiFGe
X0ZSSlZypWfsjx4h0qW0CGzH9VNXKCS8FajcD49l970R6SdnPEI1GZ2FQvHwg2uyleRk44nCoIE1
aRMnPUjbhwz1tm46EIfyooTbmrfrXV0w3shNcgui1BPDDfWQUqH08olJMMiOtgBvc4bEiUQyMt6l
oaUNXibum+yXdNU0+vBkFPvJEV8Y39k2EYEWWs4Yki6odnNiTlKn0bymcLAH1d/zJsCeQMDJZusV
r+NR31E99NWsQch64tk68zDS892JavsGreOtKq3kbZiol09+2lqdZyn5b/jl8bvqEcxhITyB40wi
BY2tKQFWpE2/BRPXhHgjmAlsCA+onqw+gwcHPQ6h/qHSlkcZvySdQcFU8JYX3HFQ0QSF+Y0sybje
lxawOEx58nUyzSUJ/RwKm5DxSCZY7HWKO1Mckkbesfyrw3hhuw/I4UoAdxrRdjmoBjB9NFQ9SJiE
Kyf6kuf0CnKY56h+lpWPm7n1aqHMHjdr4TbEYyK/D1r4VxYPW+RNMnUh7Yfm1GwHNxtg9ikeAW/l
L7sGwvzd60j6XxIJRMP7wqmpslX/WkS1zeFr+uCtk9Pu5lqaoBMKHUx+9UsqPAfDfyN+//Mpo1EF
WdBgEcyMCRyyh5DxaumwyakiCeBcoZ4pypdlifUDNOZTrbgG3MITi8L6zZlsy3vn1GCpS9sOY6lg
QoDbNk6q/M7XDPL2MGpH713ogHJIwk4rTpy0L6xCiZNrhYJQP3Br/1ZevAlm0+8hZJ0mxyHHp7u6
EQPv5nofqCtzQR1WlyDqr+ceD/h/m8kjm1NeW/PiCR0c0QBY31Pv2LbYKWHpn910xMpGKmPWMjkz
yeHdVw3w1fs3y7vvAm1gRi95vpOTmAX8XsQwWnwR7kgW8ruudylj5xOHkOTkIl8SpxdXdZSlUEx2
V25tpZLjN1m3NZKL+gP2MZGqlH6V/or5zooxOw/UkLgnjzyDkSyfvwdxZCOkQLkradsWk00LK3x2
PMRTm27vjuWA2+ZsBYXbKjU5Zs5++R9Zl6jM3aBDPXnRSNHKB1eNmTMth1Jjtwv/tIazWn1q6pL9
eUJjRDmrXbScMBgBIE5YavFdQRziaQWbbwqk2Y5NywopUufjP/xRwZzC8CeGH4TPymsdbRVcWx9p
tZ44+eS5nZwZRxefrGjcrFd7KPyLrHwycerMXhkPd52yuYHdqA8N3+IJ8ki0lMsY0ndE/EyQvlzd
W34Y97YJ816aRQ9l1PreLjk0xVWb54xM7u7XhsYmuUrFKXRoULJVYeTJoEIGj81q291knRlpUfGG
4jhK3bxt5O5iRQ5QUVZbIqb2XLQ9lcXln4QxW/Q7dOq1+HpwEQ2+19jBm3I+BdcyuF5pujBlcToD
KqdO9xkxiAmSUoiiGlx/37FzfkMzGGm9qOAdNI7Tu4YQEslkxLYKUIfLMq64llfSMs1V52q2zubF
dfuJ+eoS4shfCi2eA9m0BP72iG9UtDuJiuihQNuWrCaN/R/QxR6pHr86fE3SlTUjpUEJpR0AIzmC
tcaRfUfhi5ULZYW8dhb60D6iefe6+T5TIe9bK6UwCrdaxRpTXanq9dagZBKveh2RPkDxUIOCbLjo
DZ9Gn4UENgU2L6KAHRFCZt1egiPcD9Wm3pAT5SZePZTC1GSTLdhw6VRab2Xwq0CWmBgVTjDDc+JR
IboYIuIpCnq8KUdenyuHJUf+VHjiFes2SLOctlBio8z3NsnblqVcFQfDCXFTCgpjuIXptX4HtSXz
jGj0AldNS5WNlvNuVwMcEVk9S9/ImE94kZV5dD0SPIOrGMSZ0A1pYEp75ZmQvNnyvXpLExVH56ew
eaXwU+tOLUbCPtbrF85N3hH6EQwRaZMVjsTvZADHm0P8ntKfoiTlGaRwkKl721mPwEs3QGj1r6wY
0J4duyVpAudIqcYaO1miTn3IMlCY25bCJiNFukI23HBBi5SH2csq2uwnYVbxIsFdl23drQsxobwG
r4kiZS42DH0qXMm5FlCcD+Ivq81orUj6/qcV7EUBOrslfVcBsdIKVO8ILFYl/MhSRrPvmAtr6mKa
jXaw4wmPxpT5FjdaSVBOdQpxoGYEELx6Zw0/RJQB1MCBJewJJweRLzVzUZdnkMV77A0N6D+KI+Hf
A0HEbPVgEnpKdnwJhvmdm2zRV6ZY9baqE56RkQAQkN0/jBQZBG6qkh6D+wXOUSK9nsiUrbJb2uRA
G88UsO7q32b88s/lEQiLRaz3lNDdcm1AO+6bwxYZ1FetuwWCmHQP28QZj2ZFxu7WYtoaKS6cb7ha
ckeh9zqUCELk/Fyvyx8HFxh4GSNhu3mWttdCSBSRN71kbX1MFKJw97ujKB8k7cfd99OvnqVjoIbD
EQhY2FtdTNCLqeMQt2ffBJflYu88n7rxy8MBQiVJWuRn62Wmi0pvIrcMI85fOTZD3+oOWmhC136E
EYvYPW91Cmn9rwoH8WfJLSHDLMjj2CDqbkkOBbCcZPvUGIpzCSW44BcHTQB1f4lrXdTWpS6jJTCt
ZlfcihvGtGC6rSxfEC5gp7mbYshxQ4CajNHdlqmbrruf3qKDgx8AWXkfjG9ZkU6e2Jee37sXk10x
pYV+RpesHe/PCGlnkF/rOJTa7+klydgCqM7caCytgNcJGy+puxAXLU8ov6FybGZHFoCePeFu6TNM
nINZGY2VYhZ3ZRiaxyV6wgAsPzEyzeeIQLsnpwzOfv6EOYDHeUuVwyeYRkt7VwVinAgX63N8EDjT
gcVfuHXUQtVVnMdCRWIepuMe/U1ka/dEYtiPnSNmFgtSHrUX39xis7VFPociAUQmSx/VBOCc9sqe
EOasCQvHqt/ZVKOv57kYBvhBrUVo98CMRo4NPWxhCdFVUQptgQDSybqKCEshPnWEhWA08IpvcuLC
WlKLe/4+bOcfsnhpg/ATkghJpNB227VrGngaO9yzE53osJDmLqJCKCiTvjwcExMAbteivG28NaT/
5egL3/mqjCgE9O1KWonfKyzltZSGAx8u3YydZwjPQvxFOGiYgUeOZZmXmPnmNxfVHb+6V2ystJfb
IplK7vZwgCLRX/17fMIH1gGFCkmZWFaQR8uZ11H2t85HcKMU8UJHxMUZZEy3Wt9E1JYa/FS3G6at
w8sMrAd8aB5pAfSLR8qop8afQzN+LZL8JkTGvLNzpuArUf8r/AfzQkJQQfqLfvScOR2gcj86sjjR
pg0aGSFERZhpTTBdPH8K5J8vSFsh3Gg20Xy4GcBlVhL7CGp+dHXSuIw2sDbaD2mpJ2gnlEPM0ih+
EUdoWScgOtbSkYAJZD9CKx718MpnrYEdP9tsV8oT6pJMd1ABaBwf+qc52xBPbBOPyimQ2GEuPY0d
fZBq5Q1eoXLK4fYVo/LT800E/2trUlkX3D8EmvWz1meHZYdxvHOg3IlEZK3yUK95qRlWUywmwd1S
IuPaQ7FSty5BF/YumbpH52qsF7zCwFMsBQ3XxyE9gBPY8P/A6D95hFFeL2fF2frivEC38J2iRAyB
Wr0mGQX0HJ6D39KRV+KHrxXl8hLoKnrWT8iOvr9MTl+Z7lnqTRMeTeriy50l+dAY7Cl03mysme4N
4QXbTiaTvYbzCzvdqxzKWja6ZhfpQsH1zmAu+s16eFn5SWabKM/IEX51vdStI2hjOmN8lGE5jRbs
0mCdi2jsbJTI0JpwQwcRj281plfzsLKZX5I2cF30dw3ElRN3uDqna/4K5VbBZ5D0E2BnRFpZ334w
Yk4dmys+AQ63KWyPfooE0Y9MpjP46Fo0lqTbeFdSZARlSVDl0K7V9wqCrEiH2Tz1fh75qzetlWu/
LWzpFA0ESFkwf9fvg61NXu7LBisTaEhryZRGOkWoUtH6Hbwj7GM5Tl41Vk87JPJK9BrpAg+Qu8Tj
QqhfvKAtVDMAAR/4WwumEHoWvOhVGvXbY9QHaJDZzEy/+XUe/DhSxY0dmOkFGIH9wZgzUe0CrBqV
Bm+vwDD3fpBCgVZt0d+XqKH7AvuqtgWyOscyu/EmKD+xVmH3wEH60egZPDj7ypgG2+guuKTLh/3M
3lfPhVUGHAys4Cj9Km046NJhDQ8xYEa9GtXRsCt/TeJLja/u9UTk4L3CNmhpaUJUcvN0iROAxamg
VUtFtaU+fZoG0njHjS8e6u+RowE2+HabWYJJ7z/+361ahYqnunEDXvorIpR740YYKz+/eNGmjpeJ
p2XF+p1I3v/p6QYR7mwj3tZknzv77mdRwjzjpPZ1EeObSVTX1gkZbwZOwi4NPufB+WEaH5A3WeHf
I4b3gVWikr01gJW5AocYpspRA8RBFglpAVZ65Tqsni6sGnzsAvNQIkMS84FU2Gj/6SGapxW0trpE
RqxEl6VH+G3dZpfMQ5inUXJ/hHxsa/tb5gghKoDOgOjFPeazJ4r9N6ABj6ecjS1uJY4BCTIcBiVw
KKTeoJyz4rONZNvDWRtj68oNxspadH8koX2FzdZ3aB6kUtpNBgN8dwwA1Ql7Aujt9+7OdUE0fgzH
vUP1D15ECuozJKOVO75J2c1WJO7qZNBS818jiHx+WoKWRa36nEznKj0gF8MoKS/2bynrA4ohNZJo
evO0vQvAOpRtYHY+AV+idSLRORCK/4fokwW3x5vbmDpZJfBXrhe7l56B1P9GR5AFn8OZXXikkZzp
gMWmSdnzYh40g9YOdXaqWdqCuzjYOyiLw9CvVsrhZMJ/djC5Ebj4ir75T18xaFJf+dFaO39alD+M
2n/ZZ752xNlaSalwxwzCvrXCHX4M/plgyinqCG0TyDBQJyqhD6NBm3oY0q5C/IU0mYImwfWHeXJX
IphxuoOAeUU/Rxm9gdjVm2m3tXd3f1yOqv6M3hHguhVBCPljEtK/QtgHxqBE5TTccQpEWgsAAQab
Zi/UZGAdFeXj8Soh8V+WN3WDKknj9nSGujf74cYygyleyt0xp/O+flncH8COL2N8uBPQCcQ/gEAe
5/pUS/LYkaTVoQsvv1k50hUQEblEkw2220xJHQFwa/mlnktUvDoQmzvIvUaKxBdfoeBi+qXKiShm
aXS2EBbM/mZAqDsT6G0q6oUR1DiguzlCVHZvqKulQKwQzzhAUe+d5D/rj8R+wQE6C/uRZf4cyZyW
vrXV3jreXUxoyNjmap/ruWDA5yXrLGSjl927uRuqxCRD2lfSPR5MMjjwkMGFGL2xjtEUzSmZkwNj
42QgrvokF5RArJcQeyNq7GCvUj7dbYwHKTcQV9DTBkh0/yItQczTwHt2AwB+lUpXqiaz10m2419x
Emj58k5wZ0hb9HDnbp1KGa433hehWqGSBIdyW+JVnCZl95sKs+7kTiBZNSe6DWoXvcTZ0VQlvTZm
xK7ltaTscYaFts3plZM4qVP4HwnluNWMVZNtrq7Wo8vqDz73Q0UXaKtnPH8ZKlO0f97UD4ZgxDNW
/us8+fzdLqb6P+pJOZBWol5YK/hsumEe13EhHav48df5jFoA2IjOKh6spMD+hQmgRjzJwB2cYyFO
sX1E0AQV09iwWXL2EHjEjYMc/WUHYk7YqzGhF1OQmA72HLOLx5coNLqrrEOhRcGV2G996zh3UKi1
igIM6l6+tLShmaJccBKqNqK+fdCJIuRsk+Mke3r2LeUjhss0xySbjlxTsTa43m8CHNGV3L2PEbYT
bioqijTNSC1BL+etescGtBLKLDNVYxeWhnrM3gtJe1jf1cTznDneP5H4qux3II+YubgCx58Ccwx6
tuGLta1OYrKWbkzibIszzOcFqvHcuohaZqZsgrgtL9FhBaR3H/QCP5pJErb0jFDesSm2g0K6D1s8
dynU8+IyoTHCXrxw30zySZcKj8cTO9ckmMi7JKGB5q5PuSsqGiepLSODvvz638RPLvbuFNWcv9sc
SDhWxw9UasknVsArTIT8FGy4WAfNjZUayiNc5x3MmGTh12/k0nv8kjQe+aBPzrv5kWJhkA8jrvlh
Sp48jtaZRWT/1DLDpFkM66sZ6SARlOo6tc/r0p8JPqLodnWjABcsPp1MiodtGV8TE9F1+l41DIwW
vHsnJNCscNF1m1K7uZYonQOi2yFaxvoo8E9M45nfntw/ZYjp8mbSVJpfzx9n/qv01b66PXKDu0VK
ylHtUlLmF0wNJBsnfiNiV/UCQVfbIZTWXc90BLN8Le41jYZMB2fzb1u7A188j9LhdYHpEqeu5g+w
kjwQ+MmZ/CxK9Zknbdv8y8ACFAQEEivJtp59hNjVnoIB/jxTnD17eupU7oXzfh+7FflCUq+ZPh1n
0f0Tof8L7E8Hjoz9RbFdgdim+MtnPSlJSPF/lZAqBK2jhabSErIfxjkQQLadw7JO22m4jXhkVy/V
39MCcRVeJeGOvsE7H+as8bV/ghvnAMn2TUFkZQgYeJkm9DbVtdmmn4zuRUMTNNQad+LRQUVwSTxb
U7Jco4wgHupmOoFil/Uxuz4DbArvW6vwV0IsxQ+TFjWaH1LIolZsvPlXzAGGwoA1Xlk0niWyfAZZ
JwIgX+wBWaQSmhDVppTLTdMJ++1BLY19uqlFP7W1rPel88/IRiPeyVSesQQ/Ijxw2NInRVcileU3
hh7aIHX189KGjnRxt73+Q/bBcj/Yl7lxxZ2Q8wKIsTH6uuNVC20rYZXyZFDyy4Fw5SBAYiiam8gg
b2SsQIdiJg6p/Cwr7XqWKTvGOjsvFihqkxsMykIN5XpTEeBKhcm0V+SbeyQu0hX7hU4GNlYD05id
Ey5U6TFXjOp9PCJ/mx8pm9xD1gqZpq7RU7gXuhuZQbAxFJSYRoH14GJUzyMBi9ErV1gmJNv8Npdt
c4JRzlRE53e7uuF7FuDMixTR4aOoG2SOE2OyMUivbsqq0KrcWjHzGsJs7GuV5fbQkh+/hOCN0U3Q
vXp8gYWd+mFbMWPS9uQeHu1tfOcG9z4+Ld/Cn82p+ULGrQeNbUDMqFShMleg+qbMA0mg8GenT/O6
Ocd0Td03aDZhRLYUiJ25N1LiS5wiwBtHeuf5ouLTOlwKL4WOVQYKc7vmJ2ydL/JR0sr/XAB9H+1v
eGD3WRFKn/QjkFgafRKGlN/Y70ffDRyGW5p48Wn5cLUq3KRcQxV86mzmidPcxOSYzqEK55A5CIqm
6noDGYoJQNCQPXM8AfJK4cOld7iLsZZxIHliAy7KOIvHyEUcKLBXpZbmWLvzr+lihX3CI9XBc1Nv
eQTxkSJcs1bdQjZ+X//Sf1pZ5ivvpLYjGsPONcugQ81/GwhviNW8RQm/alT+ifEk09xA60NlFnjo
P/ZhtfkNo0guOUv+PK/wcyr/a/EzWhL11I54Y651PZ9MD7E8wZwssVCBA1cx9oEMICpkRHBdPBi8
8NxHuSD/X8Zb4BANzzlukIz5zzDEHfws05LHLOXb/EAqpPahdBWtMcQkC/jNCtVjJtz4e1onEL4A
Xm34G9P1skB5gHzzNyqCjxs7+9isbg1ykRPIaQDkYZzpTGTWdjKl359xW1nw6gFyjQYMW4yKAWpN
NkPfD7c4YkqsM7ohlvTy4boEVLDD7zo79ebX3L+R9xei+eYdEnrbvIu9IMrV7/0I31DawdGjogMG
hQIzPSv9hRRUcGImQWuZBYyhWZx9j48g6r9DXoe3tqerp+JC+zkRXOucHGl+pKgsiVZjEVd6pEHR
MMvDrdfDc3FJPG/LNYWTjiTNOHt6gpUXQpz/vqJZiaAXeP5/HE5ZmX8PM0o7H+9WDedlOdMVGlZc
VGmXPhBqrYFZQleUgr6QR94FgmBYtfVfUcNz7zp3mGIHsGZy5QvKAyo53lbKzymYIOdPvAs1+lHw
Mz+3eUp1OOGWV7muRt6RcoFfjXtT3dNa4RxTMvxmP0bsvP/keW7QbLFZacsuE8XWQ0yVu6JynMp8
OHgvJvryabZc2UoryYyzKBDetF1bBHTZMWbyoeZYZcgzApkm71HR+GPcaBVOHuc1kxYDxYomrh5g
ndWsEPWyxYur7R2/W3ek44e4Z2jywvigxcmBq2rISAg6bfuO4lQuxmrCI/nVkXFAfJGViEonvt9b
+/nDQe4amol4MG4jjNYH4TRHrBTfYK+HuYtGBEdljWB8OKV17ex2bdHdb8hfIZUqKS8TvH9kcVzF
PmqzYij1kP25pZzZmvtf0stkkEY6jzpQvTmWv1ruKrZjeTWIv7k2wnojEd+ya5j8Ye9xT+fRFstw
RF4AqSEojZiagk+h1YqQbFCC9kRO26SMra9zfYGdS07uhBh/eaechHke2mwjqV61gmLuuE+wXRyt
eTPdtKvxYiN/JBMB6Dt4NAY5OjyWGFkZUhyErS1sgrh2yvBbTBcH1cEyZrXg9HZyHkZFfxo56Nly
wGFPDOUaB5xACv9LC2VX4DpBc09UzTKgauGetMK6dj0JlGclgH2Wzksg53LRSw+I7Qd4dXW43ZIs
TxqGIUCzsIUIXEjeJ2Tet3BinNmdYrwSySeCACog5Wgg2QdnMVezaWCwxmpTOyRaDgut0kvL9hYZ
9wLZib7q89UzHpRSPx5Rj4eoxAyvydaV8X/nR1/7EsVBSET7d4SykLb+/22wtJVcOHtWVI9udc9V
AKlQ3wuii+Rs7ZbDKGO22S6i8ZSe85dDUSuou9PuFDeDYvWzpEBhSiSl79aRq4AmqwsTQXEpWIfG
u7Jg9tXEts7sC76Xs/AZTh1ITPLaHMGokwnQqORUyIAnbjSTNrlotrDMcmgf7ums/C3fABxDN7od
qx0vUUAM7nWTvvzWfUDNs6u/RVZy0y2esAy80jxn+xKeGz7IJeHBPLSgZcWsjYKOYWW1JsIMQdxk
9itWyplYVmyj/wRydftI0p2Qcu5+DxFYtM7Yz/LwCHNZmhtZu9dUavIZJ1aFBkpTIC2Y3kE8dGuI
tKKpXzAVr4CvvFq+yInuS9MhY5Vg86LF3u5G5ljX0aLwn0uJQMLMr5GMNEIEbgHJVWyxVa8duDKO
OnfEh2PD9uXy3p97Axh1BjtFIDoV4r9la08iH8tphzuXux/2H5n7vgdvzwQxYWSMoooQPvKli71D
cRWCivy4hAfbL0CuJ0XKqWLKh4Q1wD3Po86BqYac9Ip57cjtWYkFlQ/s35YJFwaiBPa6UsJKjTTg
5BtB4GyJJvZMTYjlBa4heuOEyP5DIFP/SZ9NfSc7j44GozzHFp5lp3ZDz0q7FG/ByN9RHbWm7rxZ
Sj77bbZZ9FOxgpheYrO2OM0BZMrOCE4GDulTroDLORmy6/3fBCtVcl62DcEl8F+shsAHVzUoD+ma
K8lga0Xd5mVAVERx0ykGeTyUuj7DscCWDqDEAnUDYn33t7Qqerk3Qd4wWnmgiIADXxxKXGTU9dbR
96g+WHySxY3dZuuHCHXQufIJIRrKHCsCbzDKpct/IarGubQpPHUuoRJ2rOnd3If8vlZIghhGYdLc
s1C7Bkltw7IIrxMuRyfYotKloXVVpEr7E6NwzWpeA1dswaDjdHm1aOvwwDwx2dDs8f0Te+aN39b6
+XRXRgl0FATMJGmyeaM1MGtJuvdl0pae6yW7dnusn+wHlCzqJAoKFLeDq5Zb+CKsqM04jC2ASD1M
HJoOpTI4aC8AG8aYk2H+WmrWR2F9fG3PMfkMVUUEs5vJZpIeQk21JgTO4uNjyNWNihmUQeT1yUvL
6b4fpPiCETzYkABkc2aO6VJ/iTFn/Ec1N2+6PVyvBvwwGhMP2vJwsb2UsA5QPoCP1ihSWvA22r05
Z+N5c0KMNXalhkwKsgJTiVl7E+Xf/LfJCK7G3U0bZu1GodcKPUlAxz58gOqd9ZjIZth+2cE9GQbd
zp9aNWx4PH6GSAspODCuSm9eHdaXdZ5nezBU88ji27EG5cbqvH6l902gU+zmBppb2tLxb24na5RB
B0UF8npSEPitPwPYRU6VWkZhgKkWhO1lhslq2AcGlgQGEKWZzVT+Derwu6NamiXAVu3LHtYxIF3a
oQykKYUs6hb+3R0i8bzp+XvrEwOsU91bmjRPCOAmHaNo+MFpndDqqeeWCKnn7W49vavhHxHVRp0T
NPtVqSnEOe3mP1cxy1VINDp9zYR8gCejs+IFHCjX9ohndQKR6gzRsWlB0eX81huItKMvuayO99I0
1/Vfx8ahGo1fAELJbGiBMWY9AQFGmxacWxl2/kKzPnpQz0QrWJe8msekKh4kNqfDl+eFZvD80HmR
Te94Ts0rwbeXmkIiBMHFjQj+055jXZRhr4cJuqa5+vntJRpLiHOdZUSukm4ztoHwRUyUeAnkvSwQ
c7hlMgH/3LWURex6vGdz0Rn7D3nlVtRW9PIW097RAoA5y4DFatyaMeKFUBMoDSyvNlxr4+qaxEx0
LTv+HqEpAm7evLEFA9oDto5XuYUfbLwdGYWFP9q1E+2P0DjKCHRl2Hm66buLwmglZg3nSAGZ1m3k
uA6JVyGUq+1a7cXB2cXqPB4WeNvHMX/k+m4sBOV/0ETCyzGGOD6ZiZqTac2t3BZMqaU+EkTsoc3H
MZdjNsu6lTk579C2TW+8aCap0Ru7rzXt2eXxzc0e0z4+vFONa8Rx1+DviI/VqqrgEhAIM4r6MZD3
hDq5m7LVApkn7gYIT5oYIS1/5sXVy/4OD6K6Kc8ZbG+hzhTcPlQdOlxr34yK+UBrvhx/A/4CL2Mu
gOGL4YFQRGPrxDSlreSjThTd0dAEjodMW4Ocx8RymzJZ+OgG5b2TchJgUuOVrRY5nRJSfzLelbIb
pX8vJYU7ngqxTyk5zPudyf645Dmq0dCAgcl4rLhEBizntC6YJJZhV/+s4Dvs45rRFQRqFTXlfndI
6D0PH8tP48rMdb/Ad0AjEWigKqrx6rAkvOSirUxE7qfkWQbuh09JK1FjVh5egTUroreU4OMfP5HZ
lA1GFCSfanolPO2ZDtwpepM6ZwEysJ34+/7bCjOIufV3IQhCK18x0kvyXkRr/r8vHdgrMvZrZUm8
CWasM2qbrhO2sbyKlOD1oGJfYGe+BRZEbu2DmB2B0pedDrzjF1evmztBwHWgcajhpchvGkE7eqoL
gYWrpcL22ymMuzkzvAfDN4DOjAivUUamf9v3+oHBe/R/uJbzsPBnGlRdAeTjSdXLnqFsHtvlX/oC
q07dc1z5V0fUqnSnuSr86UMKK1JjaXDb+0QNeHA2PUE5gfdNjZxKib99S08p8TKWEcqeHWYQr/N/
MjCNDO/usinAnueetGpNRBwF/2Rf/5FuRoeQRfv71tK6UBGavDwAdxDrBxsErhz/xVl2vUQG36g1
PG7UWX48BunHB0GxJJGlXTPQy8cMkSQF0ZqBGRKOQsJOG8bL28VHRXErUeq9oy8LpBrFqwPIiZEg
1qkJFjnCi3SVupZHJsEgASm8E6OfKekSdBz3G5MODErWV8sIZfOnXfbm4oLnKTdlWjTXarNY0Il5
fqOjw8JaGEgMjNjCcCKPTn3X5R9M3HbVsQ5vDj+z+gGXp8W4G5EaVoBQPxTk6rGYmB4Mhax9sII7
uod39MsBoZ4Qc/1oQTfZu8Tc9gYWHNzTHuWGPTKGev/34+K4UrEGO1KdEhYkSojbV3ooDCYW0vpj
m66ePv0MRixnTa/GEpsdFfIKHdZIbvcaAqDEjLlRrcJKZPHcAzKRuhjQbhks2Xf6Wnb8RL8Fc0KQ
wvf9vQExbJ7QWfxxBL45K3aw5l5WuR98Cr9ZPhuPvMaLEZIIHR68XE/gu7jl1ScIOQKW4vOuvjpO
CIvgZT04dKDff3lc+9XwY275Mq7qPxkboKeVzu1tFgNtfp5KXMcEktGmmxtDrhiT7F27FdlbiZzn
i9uaWEB8WRM3nQR40d4hmAOJjdBTPZsh8rHsWvGG98cWc9b6hXgnbVmaTTskTXBr7ct2cKMEWe/r
H1PtBkSdj3rewx8ruUSS9aGObAIXbrc1LtoOj2O6+lsjJYSheTSZYiTo9TRlo3fuUpoB4OhP4oZc
wwNcxDEBytd7crjTanzmfRkRoiwLZxQz0C6reCsdR/uRILfc+i08lUdjxCIlxUFYIWrKGTRJSdTj
2d+ZUZaR4q2oaMSYTBWUgcs3no6Dc31ujnGBmYBON9dohX2jSu7BrfAxP2nbf7HrBWJEbgT6X4HW
2NS/VL1RqzXawrheHCo34NKLRniMeXfIDd3Gjfm0XS2eJnnBes8xw1x/IcTprxIotJfdozDGxxYC
T7idMqVEryO+GqIbZZ7GV4+AeYTqpl2ShpB6Bresp2QMsXrYh4MyEc/1JScPwPbjWpWCzuP5ywwF
/fI16ZeKU9f5Qy7/nxvqEk9pVVfvmwFbLszgKMhM55fruLLdqE9CiYUU71fLrU/SFmkqMCW3Sciy
fA+xuImNhxvAzBnRUJAxZnhKLfAn0+XdD29yBPSR+h5YwrTcIHKhLeBqKDdLatg7cLdATaek4fD0
4MW3zGPQ0I6oFy76OvuofKoKR4T95cH2MTVYSVSxSRHg4mmJY9JT89f3xMYMg3c/V12AUDDjbJnK
c9tte3KgFGlskc3118K1rHiSuDPmeSSjRbJgJsjtR5hm6zxgi6Shm+cTMVkiPHyzRfgR6Bsjk30t
KTk/DjlsM9E1utYMt5tR9jfhdavfpFyhVUgEW+bRP3CQVVpT7snZBKhMB+LuJsxca/OUevsQMF4J
HAqI0PiMetSoUa2+yPdGD3JM+h5U7d3fA9iyTZq9bHugV0MZkTxwE4RdYc0Dhyi15jsdV75RbRT1
S1evKgrwmzqtJ93utMmfd2aUIn3mzq0sn9rI9LJ0t1BvzawxpsNiBX//nXIGwWz5ROhUGkJYI2Tn
MuJcOzxRZU2YzQ/0id2omTxWS2JJ9vTBiPbG1Cl7nnkZUcD8TfGGyiOKgTDcvaABIhFAW1C5lj2M
9BjmaRJ0i6ixPsVYURevQuHfF0sJToLnPRlevmRxOpL5nKeUSsKIz9jPdu2nvrv/L4jXhjAcx6b7
QOZNXrwIIIZVEe6+Qx6V76ux/ffeu5C3QfEDC8Ydd5Y0DzlrcvhfUKuBfn6e8ci9CGxzrxBnfMQM
kxrf6xPH5AAj2+3FHyt8DlJZPBcx8yTNJsDjNgYGhuwvWWaiCprP8RkUzoTAyHHDwEDbaNjlNhhM
KWoVmZy35D+kszzr1w4bfR1mNru9mRepY1wTj/aTGgffNd/pjR2oGCKfD9Ndia76BAK71bjYowIs
axoK9J3UjCoTxEiGCWziB8B6S+FnUW0qMVAJna1UzUVjZ3IcAUAL6FWphVVEhajqZqqjM9XBhCY9
5BINGxdwTgU/6zDTffW951J0D59B+4EQy9/98bzNnYN59pThN2W68JckeU50Jwa7ywuUNdjKawSM
QqP4AXZH80lTCHayRLvyVf8Vmm8jvsqQANjQ0Xr+v0dePVVZS71KE+wlrK6LcdSr7ZyqUNDff9HF
l4mgtKLsDamotBwzT3fSpp8lapePagbC0twWM7hiKavR/YyEc/xkWqAso8eL16Kdu8oKDAPQG/3w
Ds1yGMcTW7eM9HpFyo770jR6XpyCHicRO02KfKK/40a0AXzGPOJRnjIODscH/QlxSntplaWxhD5E
b59XqujiL3fk575OGozP7+61F2CAhge7tPa2MVhRxhUFdK4XjgolUWHu2FIS4/12KGAShIESIX4w
sje/OHpM45idqkMTQYQA/Tp1BtBCXPbc81Alsruwx66agFgEX9qh4rjlqBkx33YDYlstNMrIXkBD
MpgO+2C/atjNyxOcNDgrDtMmSwkjUkW9wNO/VJ/1nXC6CQewXWqPN8uWYab/3c6vSZVv7t/WtGcj
WG1BG+r22qyge8yuPNYifT7MeB9ewHalGAHx339ZaS9EmZ8rJjhcRUaQrQZH4ssu71SN+t8gKxZE
VvB2ARcByzPXez2+MY+UvcSPV3sek1w7jlu+UnDjrF41sh5/tdWWg1K2JcWCmTuqQkm+OsIgD21c
7MYHoa0POJwViZQtVp6y5S+RPXMw7otxIybvhpBjbSCFJ6Y1nMT2iDsFcZmXt9u76d3Yg+RZtTMq
X9Wd4bOmzI7f71F7Fltk+G9x7Du1TVAdwwMZ4nV0pzwn3ONXqlbmeiKpDyLB8KJMvHPJQxbOVdck
juyhzavLJRHNzQt47SVqagy1TCdHatC+ioMYo5PA50t4n+jutCXefzC6AWfqWekiGf+GR0mLwxNm
BL8gt77Wo5v/ZsB4zIo9GVu/jMKTYE1qdKhsOq/IlWdRT5P/hRsAesXPUrqNB9F9VUgZWEl9auR8
dKUo71/NVLLpDtOfI6J7p4fNoiCAiPL4TYExEu1ORGnhWIpk+x4xSswIbqQWFgPk2/ZymO9SxmZl
qzk8AMZJLcrpQtrCosycFVpgdWWVW1TcsC5eRzP6ren4eE8aP6nFEQ56AhvYevjn2HhS/BUtqaGN
nkpek1UOMTG5guK5XZjpIou0t5KQuevLmSabiu31wmSIaTPHUssjz43x6BPvCbzWG6M94Hha0l4N
4R6Hd6AdMjAufozPmlYbA/bXi+nLyXPNuonD4BRoF4J05INhm9RyPWnlo0rz4Iwv3i4xUoIDLIaN
nJlczUDOJABYSq7iY7rA8Gv2HxB78bav2zzbZvu9w5thmc6MBnAlxf02cPnvQJCxFQz93EMjta4n
9deYY7xB/yumefGx0HRFs2FJ836Gwu1uCqTyDIPuMXOS6LYJwcyHG18AUH2FK3D/CtVkRkJMsEEO
h8FuqnGzAWZnvPzvQ+vrnzD+ff30zkg2OlPYlxCImbyYP2Ob+cdls/z7hHN9f1mCQSoJeAtDQNuY
j0wrejRa4DZZzHi70XaBHlvB+Kbd0ICXHUQq2tpTo2bfhz/f4r80aT9+93Zos0DnJSCMUTsObipR
/SafWj71eu8gbpht62jPyTPvELL4k0igswl7176++bQfOQ15CuefkJNzh1cEqFtDF3O08aSMWHic
kbrDilc0AIi2Z+fCbBIXRY1yDGg9GJXLQdXZgQ3RoIx32QWNpbKvCyFRPYsNfFe9fOHTSXgFDzvR
lc9g1KUHdHawCdGv/YyO6xp1dGY0GYlalJI3DlNtRP48gtvsjOSm9Z23XiVoCqs49hhrvr1Szfbu
5Q35qs3y/A7CKgiO65DPZfhMOQsiXomnl0972afJQ0W6ZJgr4AQZA8LSxtvfDz87woqNI2qzclj5
NJ+fOTl0gOvvpQbdV7bVglBSvy7PqKnX9ZGu5tr2QnAdFTdyAWAaKIhDGaYsszkY4Rj9esxc8MkP
Bck/bZA3sPYkGODnk6cJ+qIu3dQapGtO27dzXgI0p5FB2+2rm9kGatIxbHzM8CKpWXkV3PmO+GNx
2j+LsHGqlpyaDZFW3b0N8bXLPhfmsnGAVOLuZysMT4/5JryXwptySoSiKT/uzZ3EJmMhBH/ey/Ht
v2u47TN/VFQgky+gZTxsQc9lR0wnpL1YMr+cI3YzX+hlP8yh27KbgHzzG0e5BRGHEOx7vpJvmD2G
Y2p7/Q5v2c3ofPznp1XvJCvywdTstX3la4VWHw4y6jI8UhN0OdB6b9DM68InbouU3MLz1O6yS8TG
bNk9cZtzp1yGYbDuM4aQ08jl93m4MEd8XKcGq6mrqu1Aiwo+NLj/4DgylVVvpRsMUMK/wPEwZk5A
gZG2TxP7V+aSN1zLk0SWHSN7VxAeNNi8adZzUgyw3DmbtQFJ7oDg9uoDJR+kAtk28eITcowc2YLw
YAG3oi5rqI8OC/fPmj+gJk1A8QTGxLd5KjVV7zeZj+0qFFil/eF1HeipYDbckvWKFBC0nPaIVTbP
kFOlyz2nFzhpDNiNA5DQjctnt88Bz6Te9A1bDO0ppXYgtLcnKq4Bx7yE4M7Z4M1wt5KQRPI0d1SJ
/RA5kwx1vAj9ytUqOAl2TrWN1Rs1hfJ+cJi9QHWMxNP5UFL67BT/hH6feXCI9TULWCXrPsrUFQV6
Wv9cNBhIBekHjhnuT4AFE3fPFzbftVaZ6uqqMB/LhU0gzeEP77daCWJPTYYJVaUF6+214DgMlS0j
gy3lb0Z8354Z6xUsBZGSu/60CszD/51t5eqkfkkmGeNFchoU4auaZPGr4OuVfCxgD234h936CChh
TSiQKnW+f3oTapTIQDXMsZvONt1f1MQs7PHo7/RTQXYdgPi2S/4oVhkZFvFJ1O/hAiWWmaM3fOKN
5H4nLZFzJnmUf9G/xWZM3lThzc99ugO/ziK5dVyOl2SCO8gcefziNQG9YEJo5O0pVAi5xQdyw/gI
3Ce322cImPZmCbEJtH+mBg9jpbrecNbkWWJ1MhLtz+aX//FIi370nGyMawsqUREqTGiXeQZOHkgx
FlOVaKZTsf5O4nIwUlHd27ILsbVcLc7tGRziXZjG1uWSakiSvwItYiqK09TBeKvyKAS6+/+DtAt1
x82gMsgHgYJQPxE0TxBh14RYHQIPtw5InkguF+mw54UtDwJ4EXiFCaMCitkljt4l8KeXq444JxT+
SLI1wo3Tt7JtVQPtL19+G3AsmtQVIjXeSz9aLdN7mquyoBC5DYsEm2cM6+RIgDexqgAz1ncmla6r
a6rVuBbtOdCmBTLRn3YWQnNjMhHgNeXMrVHDfzw0/PQoFxfNmpxUYVKuy/tNjco5+Y+Uw1e3SKWS
Oj4QHJ5nI7O3E+8fL2HEK/xcHPRcrIp81AFvQxaP3mscmSbjpvpRXxK/06KvpiDSs/8vArvWpOnd
8t1Ruf43niCcNqdNeiIGgu6mxko2mBVelrnKppI5L8yapxNM3Evk+EO/t7Zu0FZMZOD1cVLTYN/o
6qnheXZUA1PbvvVQKIl/oA902EdC7Pa0J2zuEwStqnmDmohHvxVJpek/UKUE3nDbgZIDspGw8Fuc
ErF9PiL/gwdQbJ5CEIKHbE76joPBAPp/hPUVGhJE+SDgRypmUu8FGsBSnSy+JnNadiE//U4koK6y
MKrf09ZlDQLYUzoTf0EdDOSxGXzuu6ejD9OK9vLu1kIUDmehBuybkMsRLmpWncetg3XXAcrQJu5c
ssAxCUmRoC6P3/4QyItUMBihx7aur2oVciqyhBGd2QZuR8pk87Faa+MhdbUPzuq3LA85x9KDqqYZ
y+YXQ9fk4WKugbUZGSiQKeCb3E6MMBCllbeR4qFi3enoFbgMTacrH5/N+JMEoZqw3lNv78cqZx04
J8ym9UBrZdwkN3HWmlFncL8Px+gQz7nGL2cKtsaDvYzPU/svyqbFEjdJ4Q8IKN/h1V+mco4oTJGU
hsHCp2++zXa/cTWAqS+tgrnb4Fzrzo64PdCTaQtLVqmFow71bNL5/hLKJbLb2vfQo6Gk6gZkON4T
MKBXFnm3jn1jh4v771idu02ZXkvnqkoNZlsQmmmhc1WNLltze1tRkCxXdjOEJm1MYQCBWW0vgLAb
1f3FJRzbw1oPLy8gvyjCAG7th+nxEiVqqtPAMzqqvgrOzh4u6+YNeTvw/TjCfQ+7rLjay6Q90/Nn
doQy0nhMJKWMkw2zzzMIPfNy2m5rJYdexo5eDnhH9HmWIgYTfOJNPhu7a+nETJsDnzOViQvMEKkc
0b5OC+ler72mni1yjMZgqBk6APmt88rnjS2T5lRKbsP9ZINMttd7MOS2ZHQQDxACPahSSuBMRtWN
cxfolo78uyNBHqt9p2g6KxtUGrW7fGAX46UTPgkSIuTirl2xvuwPIrdvu3TlW5TemMLdvn57NluB
DI7s6qe+dnPayKmxucEJWtixCwbuSVkmQ9lRM8F7ol/72XiAz7DoF1AYq5k1DDL3pbQFJ2fHM/UJ
Ogc7TVX1AZzw0BFznBCHPvAAJBf3sziDuTUzqyx6yA0HmLxcZqLoA3NUdS65P8xY/vfepGy64TO/
Gxc9tqLUuDPoHQDdpAguGT2rUCHezsQ5nSiDFyuJ5426U/rh1SwIx6EuVeo2YI1xir+zEAt4UGky
fcXSe4zNCz3oNz9Gdx1FMrDU3i7Wiva6pX/Eh5qHGzKF0YpQLYccM085RS0VS3HcJJldeV1dWwXG
EjuX7vhHSCS8L8jA820tnaQm1E8YswEFHgwoYDHGDSBsFB/eInf71aURoyWgY001TOgOA9jz7qTl
hCCuiTfNXsAEFMiMBoLkc1DXXtKNWrePJLYFlyG1QDu9GXZEWkgRmMOfMs3jvctvtZ2GqQVy07lz
yQbT1ROAuKVz1P1mL/CUy1FroiOeK6hVmdvM28GgCbknITIAGt9iEbnVq7qyXV1CEhkBod97mnpi
cOrAhYlCbcbtDIE+9UeCrcWSIbQKUL0Xe1PXUUFQJDEC8weG+pmTmcpak3xAv8btEliXt9xnlBr3
cDgmWyg1muzgSw7Dr7wzkkTTjHpyxiQqbYtPlhEWBMnnygKh5vwwBulWw/9W3Fe470cVa7bUkUNw
1BVbfUC8A6+dlszsDli+jPJCQ1zEqBUSNobonpSktDmZ6JxdVGmTvXQS9kxcPqHGjslWtmRxsIAA
ErdtXy7FdwjYBAsQsEsiDR22iunFlql/0zfskD4frq/A1sKbDyDwMLkwqzKfzeYO9WCfA2tEIlHd
IpxKiYky25+uiabqHP/tYX0tzwWqHOr6a6TjTrCYAND7+OriPCnjpMXvYefpIK/LLlyqkDNXsfyU
zZ3cIx/ph+DS2Wvm4UI6BkaBW6lgK0R+mDSWCymIApddhHnU62K3FfLD1siH+TBJIILp2ZnS28FP
7EASHW+TkEXq5jDpNK0Iu5OikPdvzK4NBhTpnOP4NVFyi9ZaY2MF2da2abMKdPhJd7gdBjs94E7v
/g5/T9o+qnPTrM60H3pE8fsiCwOX80gFdRh1qcxUTAs5dvIMQ26v8iq8KV2ohZTI82x0KZm2LPxo
upIr13vDYknVPGoFTsdB3/BS+mbpX+EI9YRUl0dD4TEZSX4wc0/F4KfbXL4ke/w7PT6xQG9UVgz8
cxv7iHxyXYFpzDaIynzazUR2s0KD0eMKppu3lqWNWiFzDo5g3LxnLg2/gQiC8QI6n+8BS7XjQC/8
00UTvmRIfOD4Dz04gHUsLV3rRbdV+g/ebryrN4Th4zw1Ph6c2Zceu7k+3fy+7y54cop9Nakz4N0D
aQxIovvYihcAMstiuNi75eqdl7BzMtVzlRNQIUO9mLTcl0HCEo2JcdFRx1I8rE/4wdsj6/2waB+b
s+DGeGIF0gy0f2jfKfHtL9m0cqf1okfhQIiZ67LXe47kSgvLrbFjRW8SCmj4s20jjEC8hX34DUva
p2IjOtPVlolfgotIR5uZnwdjH0hrg3p33b8G098WUCXiNHuFn4UWAbeNvjFfLAz3ypty/qaqPPmf
VY4z8xq/hnB1y2PCI26VXqH/YptHciLXEtN13fPJ1g+NXhbqA8M3KY4niep4NwubCR6ea8p+8U8k
iPKGHhJgcM2puto9hILjeG+KAHIH07k7j0Pb7uPRn4vfdEL9gAWCDIxsa6EYIaWZrIbI4Z00KCmg
uUz7XQIXmWXJwBMeAQojYV3OVHb5DwC8jQ0AjSCQVJZzvB1f/CCqs1Go3gpOE+6Za4V2/EtXPA46
T/4tG8P6ePs4bP7rQmJ1tbWqeGV9tMlwDlAfvmPNxetCoxhuxa3Q2Wvm0mm7/YgSadZZo2z81D6k
5I0K6FSuHhUwEPAfx37FuncBE0ni4KrQictNqzLEY6U4MozoLdS8JZ0CP03qgzb5GALdQC+lO14D
cHeRNzsuEMrpNewiRhQtHGhLkhNl4bav7ys5/FHk0bkfYpP8V/tN5SDqPRQOqojii+kueICxDdUA
nAb0Fb26dKWnR7H0y+oJGStv6QE4jgYLoxDujjTE/ArDQlZJxevEurGjXN+Fr/rrerd5lYNRGeoU
kkeng4N45mSPBLa6YIm6EYgkXF2YOWGMMnH+os7MFSKDlrcFRLSjNQIipzHeozbBqMFAltaSIBHv
OUwMkRaDSB6l4F2JlLo0g0AqaI3S65HQxFmNoGnbKOuJsz5R9ZpDCnd0OdFq2v9O/EPHL4Q84rK7
L2IXKWQDqipourJvtVHNa+ya9ZktWFw3U/S8Hke+TJeup/E1Sj1Kn3/oxnJ/m2ceL8F1F2QyBzqk
hl2cGvXxdriqyPGnu9/dpAKZpbphAjVZjCFYEJLts6goh8Umtu7+FR99szCJ9/biyw/iC8N2mfgs
hMCfQMxPjh27b0RuD0j/WkPHGrOv8v+8iMvGmKl42waQJE3f5QDk+4NRJ+5BSrNO/yFSJdOgseKA
IvkIodDkf72DgVgc7QU2HlwLlcmvqSyydb+Iixvg4bXNRczIFLGspMYKIU7FOuPAVhpQ5UN+EGJ6
4aTLeBa9bj7Acv2dRLUiAPwBQwYQ5N3aQAKouMpw4cPsVTl+JRlhYvy5hjYfCQ/9Y46arbBHhAW2
0LBTxF5wcwUu1+os6B1fBYa0PG0yZjOaZmWGkskPSmkREv70uEOlTmdoeJcHNgJjpKYEOyoSyzjs
jbVcWs2QFHAtsI05M8Xl6/AoeyJldNKFdNnD/wjgto1y58Toc9UtCotB1z8ZmeFj+oeqy6Mog9kW
NpzEia6mkOaeUuRLuApHc3xlYKw7AH+iapxLNv4JkPbqJ+gyB+Hsa2wkxsXZUt7C2JW/0GORk20Y
V9QvIllL3z7q5i0q5u6Af33S2A3oqm6C6kwKT3Z3AEd0VP2d2db5pr7ubMw0rQzArsbphQopcXwn
e4dJmnMtafdgmUApHLjqbMbP54AhN9OEOUzEqp1rrHPtvS6a8JqkiAudrRumCGyrZZ/Eemz+RMz5
BlUUxff/SzUko/WbKt7wiw+Za3xc50c8Ci6+0MQzWOPAnW1rIfvaW8zWnQMOTIzs0Y8BYE36mEZR
aLoCjkKalt449m1cCV71dGdihhYh8FCZsCSlEoaYmWZFCOeWXjd3s+Jt/AcH78/hr7YnK0ioSL7g
Y/I9LuGmCTPiPRJ1Hznpme22o51t3I50MjQE4XVCuxugYpUl9Fx2F5sP8UQeUdWMNyTx0xon0RSB
BcJ2JzrAKfOCnj3+iwQ8AbiyGnNfUGxlpbN7VsOfC7We6NdJkS/h7NHkBAL41IVegvyQQTDdVJKl
7Pu989ql0os9GYoBvm8EBpQEUVUjSXdR2gdtOI+Fi4gaj2+NYPiix6GdJc57yR/LV0zYPRnZ7RKZ
mM58dWvdNGs3ctopchKzks5KltjRMU1klUog/0QX+cVs+lbjkSgbhHMd/4aBIndRI4HAuqLGmT+s
w51G6SbpI0wrt38xKAos86MdPwD2ZNpGRoKykInO8ZFpeRIoIev7PiSByYagoTBz/aeZy2ZvUCz0
sshVdGk1i0z7f5LTYTG5TkhElHYX6UmVvaSo37zk6TC03/IeMRrKNPu3AG1Io/RjI8Jc77UdXgNw
p0hPSuBRPsEt35F0tgTswLA9o16QPtzqiINorpxt1GmCM7OElwxBwrAA9uHkEshNacZsE6ckhTpm
PuheBV89BqCE0/IaOnBWXtkdlsdeDn/hTframa6pOHxNiDcgVnYVJlwkIPnSkoZuwUDT5xV/239A
4O/j+w/sExfxY4ppUqGxIn5ywucFwGtdR16xB3K95WUffH/8yC30fWUWNK0daRVNZcBs9+NacNbO
R28twkfaNeeuc7acv/GBXoZZ65op4S7vvDomflXWZOczyCAJmukev6q1K9XeV7sEsrhn3o0UfW/9
FSbFuDkShb1sv0wtb4p0bqjDmHDIRcmPU8jqvePvgQb3Y6Ae6mNwoTIoWDiX88qXK8fWPZHxtwFa
SmtAfc4JvvVp11Ktmz9d6TpFOFbJ83ZjCRTBcTkWNoEnXtc1ZyzOEf7uYn7u8m2bRxJNVlHcQwpq
yCjXxD1+XDHg2B8Yzyn8aFmnsVnQa/lysI5YhEKW2KC86NbzCQbVkj+jx4KIVc8fQFeGGZctiWyl
aLEQJTDcskQCwSWG2D1Uv6BeHiUxcvymvpbL5+BtwOIyhCc/7MyNVC98I8DUSNV2HbcMOyH0Ro2e
rk8v0naARD64uAC27yChfTwT66AoAQkORsbfvHXd59H8dvtjdJ10EAjt/60qeGqMd9T+Gs7u9rcD
ZZ1C1zLoCYfrDLCdkg+JbWArpKp2N4TmDhCae2U+xDtzWaYOq1wwmVSM/L7/QLOcFDg7mht6aW+D
5VZi8BIa9Vau//4qi2lWhAGLOWPkUlM8QF6/5M+B72Bw/645cQ6NU89/Y1txhdqIbpwpAEnAiRsr
AetRCLX9cmYQ40lNXlnknqQCoqm3PSxmm91lZB/HUI7s1VtCuHvghLc19Nd6230A818m4zz8JjKX
KgXznTjLn2pruWNN+A8htz8nInx0bngXz1uGambeymHGkWXZxOdwDvypxZa3dMaDmCexilMhLFOz
auc7YqpNUT7l7PmkfI8IWf6hABz0RdHt6KpocAfD4z8Or/FXdtULTJuqNrn6UV/laGAfBJ4HpcID
qn0MWdhZVR6TOkk2W+q4jeMgULThwOrMAqhCjhbWPwDISTYo+podzj+ZrVMUBk58UhxDNt6y6IPD
eO7D09BofmekiAtk9C2dBjizqsFtlqMfWW4g+N0tDw/Y28G/8hUZjOA6vmGV4Er+DSe6ppsiRryi
aCOqqAmnAjGsVL+nz1PHrmitzgOOi15eMk5ay71ST6ahOlHw/aDtM3t7w2+SWI0Kqab3YVV+3tBk
/pRdhTvX/soPFAq3VcnfD3pBqQrscvGZDOaeaE4+UsTeeCDPiTnenX9YFEdO+0RwoN4BIMC57LVy
jxXMjci8rBuUcH6wkZNaXq6ecIwaHo1BpJDm8P5cvtP8aC4e0KZSA432YQQ/ksvHKCvduVCTvMet
Dxpx868X63+CkgdA1LYNu9B5J0Gi9xa68JazU100fU7VQBPa9magxOwdmv3CX9k99CgfUZrz0sDF
Q1TjpjtiwBO+INmwpvvfjVHor6NQg7H9hy2cmhRqZbBuDvkI/09ycqIob49syKzLeBwbvq2Ea9rm
TOBXZYNwTIHpBv9p3USB/e2tAoEHjRGxE//PIOS3EKULyV6Da0IAKAcnPMmvGpy5BOZbdwCSr+PG
vkNgW072VTij2ype9OVpiFvhDIhU76IZwOa5vsiJ1v5jn06K9edFl2VRamGLAPYdFQ+7eWVazXzj
M6hGaLCNTIuN/S4x9RxytF6riE1Z8+kJRPGL6pqxCAXIAMdAEMymZAsQFEjFFlRKJPJY5bMj5slk
nhIGBbpcsLqnh68Bl10MProK31w/YN71bD493E7eszJwaykM6ZEO3HvEqjm50sYz8MK6p5hNRWVU
E/r/I9WG/U0T/tGfCg0UrfYFMBfQfqmyMwQPZeZETMAcLbg+U43cWUWU1o4A7Kt5m4wzx12ON/vV
vr7PsIQxmuvPM4VEUAwAV8OXyBJKxW1fsp+Z9C/Cp84CkkC+veN3kkByROx2IG9jDYMR55tPDNcL
LeL71SW0kLeyUIrLA3NZb+62augT7xrWND+i15RMJ2z/kd8uJRs0RdOorjPzrdsKBxrt0Mb0LPRc
fDL2xy6ozOCNkvMT+6NoniypVrJ8pxR7n2n9bgPcf6PupJNVQKrrIrYmfkm0uOR16/UJJJeAQfx0
+foY4pHuwiy+41m7TuobBHRDZm7/mCgPbY+xrUw1fY91Iw8PCQKPpBSWytHaDDQDY/SMOE32Iain
W7F/xET/tJMCLBto5v710ZdonDml2muEk2aSDBBAauAaEHqA2dTUQjTMqIhA6bwJH0f1QIW/fo/Y
HkiUBxAAGhlkmP84gPGa+fbTkbnviTo6U/YiGmZLb82tL+ytHJUs513QyZo0gMbDeDp5zlAw4Mkn
yljV2JsTT4Q9fXX+VKz3+7K5Zm9gFSQP39apWoJl+hWaISDr0GTaQtheRZrTkXFX9/c7B1l9RomZ
CYHygZVHEOKpOARoJgIMkCBCMUWUN68GN8Fylb0CKRNTUqCMt42w3pO1hy9WkefCYyhgTTCVssNt
H1hgvEuZ74IgBeoXPvo2DXNzsf9/FAeYFZ8etYJhGmh1f+k0eRL2zN6rPKDrfhWcn30HLUNhEX+G
S3IXI5h5nSnsOk5gBAcJiRuQS/RngWk5WLFdhcPlYvqFYjTmoOFwMHwdWHefqOAM7YQgJudr62r4
6fhLDZnztdocwyrs9co9BnN5r7LRZ6oJkP380IlKmd7AQcdCMo7wkwY6zVJMprtfgwS3q70ozcx3
2RGQI6cvzJaytLxJro3RYRKGcMznXDNgiwwEZa2bXWgKDhocg2i2YLkjAE1YSbIQisUnY0o4HnWE
sBdrUuJpPUWOpJZYJeTLfO5bnr+0tAWaKaMC4/xg19Kenj9L3EZUJ0wnGdUCnmzWO7jXSyHa+Ste
vFr57k//IveHgCgsS+MHu6SqbzD0DmyI3qi4tYqgur3kAgtmIxIvRheLUA3ztmCTOS+Dsnd0tvW5
KTW7cp0CIyEZmqo8TbYjvnIg3+3fUDwV3aBnjAkWYmiv4MAQo/xyJ7f0pK+BTIRU9K6W2DJ38U/u
kFE9/a7B+jzdxjJag8Hi+HHGThatQCzZ7skH92QdrJRk3RD1PSqNCUOCoBWW5d7p2fOSL/XqLwTU
do08PxVF1rvLnKRP+OXYcccP6owN1Ep3k+gePA3NzDDWfkYf33uKiLYm7iqqJtqoBdGwXD42qrGe
7K3+rllgEEj/s+ddCrb+ctZvZZsa1ZVBu1qUf9ZKJzYRABLbteTFZpsieF4rWzXLbQy4kK/LDulI
BNNWrvqZM5e2puNLNrI1MGbqP+KeCxeCpaXslGkJt/Pa7BPGViYSSNxETQA0yLfZqUt7xn6qIBrK
RFDVFs9x5ngdk0DCGPDsCixmAf4oU2LgI+8JXFFD5nEG5C9EQ/0fqUchARYOGKXeh9QuXALDA98q
kLOabbwlqdpK9w+y0UGx97jEUblPvIriqYwEAFdmTRuNN0FZyufYrGv2ayPj/EX8LVelmhoP9gln
W5jTnPvIbHgQfG4ElmfuNHFmFgYVCRRN0M+4h4rM3AnLZHBX/enTNRmRL2euvinHpU1vdcXawAcI
BgwChqOL+VG3RR9ITlV3O2rFc6M4etZ2H/hA2f+oHOwgNJ2KREm1WVjCwqxovaoJc7dVA9lDRUge
5E4s8eRfLTwQ8/6ua5pLUN1/OAVVKnuxMatfb0KJb2RbiWY0YHU5TPt5eht4n8D63rFz+OkOTTnX
sblZAFp0K+mBU2jO3brvGpYdrDymle8owIzEIsvZbVJ/KhxCN5QfFJvMnG0g8i4dv/uhBrVbgV1F
FgSD6ZWZ0Xd20LESjlTuFVF5OaoLYtsGbRhZS8sbuyQ4TFBa4sytCJ7gDfrLC8deaT+ezntFwF8f
3h72yN/j3QYR60qiWHbI7/hmsx1U4Nf69PVLLohZYwAKuP4z5ZhLcnxAaG9rOS/XH+XphMvREIoy
ngEn09V0Sq86LmWSVGsBydow7wpw5BmJU5BGTVVwBrzUnIlA0+kj5DUHbynMf6LKJ92ZwyvGUeo6
/nFG+2h91q+BOomYnHS4rpBecAoOtuOX7foxQ8Y4ouiAm2jLoH3Y3KrLmF/16F6hvdmMRt+2vV0+
f1a0z5SD7j+oSr8EidKRn7ES7Vi85iVSodkq5iiyaLHkxp52uufHzY1iYJki66eIAJLDVITATBiN
JISPyEOoMaTCsgwjFdQDYbYrgan9DPsO5Ty+3QfAh/PhjvW0uMgiKBWogR8TIfg/Y5z0UxYutKVw
+9OW59vE0ZFmIbExHx5hKW1JkjfFdeAn4bqfSusEKudlFUf3+2XGMA7qtxl/7BF9zIceYUHBtAib
cxr/fZUeRntqL0KjsFcTgH+ZIZ9GA6u7q/iJBgiwQbqLCzHPXTvzKgjXnpBBcWUHMt99kFee7isc
Oh60GNsqc4tQnNOJtYzqCyf0qs/G/MMXT7mugjd9nPh3wPIL9AwuirIFE79XyLzvcP0CrEhbL8zm
7Sj3dAG139EmwHijwzoYS4OVKlvpGOPnneTM/q55gmJ81aFwN+R79HszGyhDXVWprZcS/SH1fAvW
CeI+huB4K1hnEBpYYGp9S30rk+SAM5fGk5SjX5kyDt1i0H6xEPZFlhTos7HRusZJjKJy3l7F8eCs
cXVC/FxGmPJfeTGFCMQXR9gtneKnMTX1sc4TqzTvEZ+NYq2RU1rCBed7gbEFgeWyXjcSMIlP8OnJ
jiiUeadvBjWo5l+sJ/FEhJ9dS/0R6VwmjH1KptsKjk2tG+xIEERRWUTbINEkLbac9IB5tOZuc2M5
PkA8dSkPIijW/MYdIvl3JQaiuAzAUFyWid8OG+ya+gSI9kGrg/lRkILR6ALOwnqH/+sz+dy3tyo+
zB1gP+MV39ilzk3eAH7s+OruJZ4Z8fSwA34UVAIwNR9FV+m853tepNtMJoLBTotR4HDOs6e+7hBN
Zpuprc7brNzLbMiftedifU7q5z9C7fPY0OWFv5rdGMkt6zUuhQo/hlybCWKO8pe5xeF0DZGWi31N
EncXJMTa1ibsUSOLWOD+MJLYbkZk5HuO3wM2vvnTuHek7hGMBJUpo/d232qogIYodxkjD+xMt8/L
PAFMmiiKYefC3XnxPFXuDmSPMZuEkG4vLYTpAJSgvdbyk+TUdhGk2A/L+w5sqPZ28ZvVEXLwXz+6
1cIjPjGUV4K1Ipx2jOJzdMin+XAQSSd9s1chSGkSkjiwNMqsqgc8F2z6C6I20b82CiiBUwEWW6+5
iHg6LXnYN67zTYstkEvXDo8pRSZ0adeqMlPqRNfTkVOI3mYKVtcht9YsBrCQOKsFr/bsy5Kf/uTj
S9YZrcpoxT/BgHDFgDHLQ7R3LE8V3pLRjhHiOD9N3H0q8kwC7Fgt8eqn0mKaMw24/nupBzi/WAXW
T/UreyBV6n6ZKHruoYn8Yd0skKNZ252sMo50cUU+Qe6ls2CB1+YRqoElzAHlGi6O5SDyQKIjgMrQ
eAGGnVxk8FDmv9PIOt488HyAhol6lssg7hSSudpyz6/3KkdQNDliazFPK+IlrHKJmzJQhVINXlU5
J8IL7mhY6LPGIBaQBkc+fqrS0njGlqlrmi2/SJDtlXl5i+lXhudMVeW68kjeTBM5boATHquJGyU/
ypSFRH/SM1G7IhZdtLSKIWxiq4gM+me70rMFyzRh9dpCnnIBxIogmIY/hXwgZaQ1rpy3WPJrX4DO
ft/supYbxtmsM4W++ilX+zPELnKO7T6A3GSMDVnmlzp1ANwgSXgOFWXcQD3lg1gN4cVh07gGavPX
PEYbGp0wf9A3DOlsduYv1tJnATDHvesyU6/w2wgbYsVvuvICn5Vt5KpYj06Y3z8RPri7/1YBEfv1
gJOF+T0SgQMeL6GrSaMkVi+GC8Il2eZRqPyONQ9VD3XwVCS6voZ1qyQYtkx559Gj83QUhxiwSPRv
rceMIN93295/BxWrlbBqOQSmDsmEluqkL3bova6DaAZhQyGIGTGgqbOBlb3qSMbSV/hKJCz05KlQ
R32dJeUh06kCuWqiRKF5lckuRyiIn3hwS69w4F/SMP5ljt9xMNdr17NeKQVWGb+MARytV3a2AK11
t2TmoCDZASjDkCB646fvoPsZMSGxllEzefAt9KdG5izoBEkzSkdro4Tbkyt+NRaSowhPWseUIMFW
p8EW86kaywlgFT5qYRRFfcyodbdRJqxsU9Znz1Crke5p2z/AYrdC/x9EFaS4+3IySiXfoEgV//QN
QB2B47/n9aP0jUlnjIlLwzCRzXjzbKMvJ9FWeBf/ECKFu2FboFS1W0ZrikS/aI5zqvpsRXwzfKE5
cpLuyQqaYNt3BcoG3HeJGIRpEXEaNIKruM+8oo8G5pDSCNakEOxdES+Z8dm+Bav5yraNMTtpX+pP
UZ3BF9NcwLXaoBpT1NKizbYMPT1gZ/zpgruragvRuzaZ5UAnihAeS9n/qk01rjZgDja/fCbpxdNW
I6qgQpxDUKHUx2LTRrw3MjaJkjvLE3vlPAQ4BsoHyFIfoqAU3j7/B2y28aoWCN4vQE41QC5OTsc8
C9CI+wmcvQP4cN+ei38m3Ij8swBJcdfdlI1rGdX41nH5Uy0OGMHvZyqrBVLNGln0jPwq2pmoLxUm
ZD+oYNNs2ywtsXjEA42f6dT3vvtKJouuM5s+QC8pZmzNnwqytcWGvScEVYa5bKiQCnl4CFhM73MI
SLeIGwpCQjtZ1ZQbNFuWE8kRqkiPHvRYDb4BE/S8c15tJlt6aqHMXb+9GplI9j8DZJlFuXd0VSEO
/27WDm3f9DNtHDP/QAjYXOVES87ck9RDG5+WweXq6BHMqnSmMB9j3EuvPAUBhqiTmOmJiPPvI8TG
lYp2hsS0bYXEaMbhJDnWqUQ/1AG8CsRGqLL38cgsDzJcUhjv5Sx9v4l1fPgzdwl8wNXn1q/HC3rD
Yx8++VeyY2D3ccC+qv/K7hZXEoYRhv7Q+AeaBCTwvM/hfs4Ab6oUzNKRkqUppI8yWkgDr6TGS33g
xXQLLyVFIUGuyoZ8vxaLD8nPMk86lMX6RzFTKuaG5PjbB2DOqud+fqpoxXd95+BvuyS33oyFrP2K
0w2NTgzVMmYkci/lxSrP7MnDHAaKszkTRDZU0KdJ06krvGRtfuJez25LVOUctdLjtXzV/vjhfFnK
+hN0B16KrAWRn/M91cDHRcfwx88IPtlUCEO+VJ4eQCk9z55q9GAUuoFZ2hGKvXRpYtmYQ1/Oxsc/
exoZMe4pArLxtQP498haDSFheNkKoiHaBAS6xYoIJoa5bXmpcoC/ktoC/cWdZTC5dFDShAYStjzA
3r1FDxYwUQUUtyLpC3RGCj5ljGTBIwsZARS+GVQHNXfqZRrDtRBCdggENg/S7Hz3Qy0ZJJgYMYKL
rkGMVkTc3zYZvhCXdN/SDPZQRIFXMibqHCS1BCcwS9k2r2fTawIRYfEt7QyqUfMUSmJ1TWURGq03
fSrOQ6e9uuti6uFnRhOmyna8lign8wlaR97TU4WvdS1m8edRDuOX8cQOdi4GLooHiR7d3IXI9J0D
zyZHbW6ZRpzp5ao122QbxTDRZxF4kIH3pUCcBYmmsxkCHzK0Hp1NbyS1DMIh4CZ//bAPo1Qk5Gs4
UqWIwJeyk0aUsGc8GdASkocoYtmTVUIm3z/mmG1Nx4xRNp/jR2eYJ0JLuVW3MgfoblEFXs9tkk99
YK9/3t2w5yJnr4Q/yEClELfG1kApeuZSB5IQBnRLwQM1dXCh5ro+d4J1VmFv29sC2X91PuBJ4mYk
3Nqf5Tboi0lFjP88m4Qecp7oP8NIrQyXUugDjkdIqk0EmeQbQX2beb1TV/Gu+VaCypmOZzw7iZyC
ScExywnCeVJl5FN5FD6MbTSl/WhU+KnvoB0Opovp7IDVRffTV+npTNpsZ/mABqqma/U9DDfAH71k
U5NCn/JzkRKgUzQEPQmv7OjEhwCQKHjMie++mbpFKynPKIWOsgosEbPQO1i5Z4PDEHUkw56xwTSt
IoBjvPvUnfKuc2BQsNfiEvYmFXZ8BZEx5H7eK8kwih2KTZrg6xUFf8uzmHbN2xkBl2S+byHIAN25
aMQZL2czSjzzhRYAu8gcJvlPp9WoeDTCd3/V+GNg3ru+n9zEF/iibHnrENccVnwRwFtxhjqFcN68
jbPTBYE7hknWtaFI3fx5mj6/vm/DxL5RjGbGweazfhABvCxkMtZoFb/qVlsP0SteKs7Be6XyJu3N
lZ8y+I6TWdARglDqOMh8tcPibw3KGlV8Xhi8CUGPrzrHBWy2iwsspdX3fgYKwxFu0TkvSlocQe/j
l1Ymc3ODA2jl8dFYCN8xSOjUX2gfygbAiPxFFJ63IwGhUaiWiqahG125DyIv0rryU0wJyYy7eS8Q
HVplJCeGo1jMSi4XAbMFyg+4vZvKYpohS0YqSsVPFRCG75tYjFZKIm4w4J44725oHwdpRBL4ZJ2n
ApUZpp5bY1bLb+8bPer289F1Agmf9Rh5ZSHsx+Lvvsm9Apg5q6ijK1g6XDPt39Qkz0SA5NHkFeF0
s6O8HxmbYhmEptxcluZb4GqALY0sIxXQUmqhgEz2hKTXQHVS5QbXDYOyl9LOnWPZnDxs4w46aMCN
/EUdsakQD1tEa2GUfu1aMoI09NF/AgX/tC5DwByWedbi/U5SK9R+1HEGBJVsC6A0pNSntTtZjBwR
10SX9QLtt/o0yor9cgVSSpH3edUAepDY0yHlGIiHEPT2VkUvLaU08Xa2px7dqgwJFyDCt0cozN2v
HZQQoaeSLP5BIJ8HxaDERGy6Si4ok9VJJzkGiDtykEgQ6ycpa6T/FhA1AadNrIezziliKTTNA109
4ofj7p02wLbIRCF5mvMWDIi2EZKcViBjQreonazJbP6Pqm6h20sUaRUjz4WTpgM9SLE6YuW6g+az
fH+xAFehadrgWRiLCvl559nKX6U5DI0HNzs+OQn7es0PtHAIqoF4PhhtW556K6M4HXmhcbVGRbWo
gPvXZ4PuVYNiLFc51m2bEtcNn7mejx0XEPSwuQcCN3cC+z2Y8XciPSEZEdXPh8otD4XO3OG5GKLG
kzW2VGGu64RKEnuCDbNxaxVbgngAm6249B0JCbxMnI22rYvL94VKe9fxKU7n9YES7fECvKWfM9Xo
x4L4WZRkP08HWrCGBxTsmZdM11FrFweiYuB4YOHwZFWqIBokjiA5O1iW1z5QtGFKqxvyoEsFi2v2
fN0WyrXHSxM8EYI0cKfjT1/7jt8cA2qUXUFupTmT+MBwuNXWpy1VT8OGw97y+1UIlg3ns0xLBKHV
jyuERIvINPTxDCGqK9eeWfBKBiCSx46B9pS+e/WD7YeU5ORSfEay2B7/6HtyOYHPu/2gzqsiGj9B
hgi4hJ3NzHLU9Wdn0Unb2Kf2aEeLcMYoxrldfyLTii8ItInSZQ0uAKuFD4If3Hb4QgVZSE/TiDET
l/1RbvJgjcNLvsUoGYwDdhtg8dcnXrgPaZ7ePAyhkwEAzmZqF2QjidYvgNzF5WNesVjUSPWPuVXW
XRR2ENH7zSoJmwReVF6W+qfkUvM5W66iAcbfWFu/hSUYIdfjkzcvjegLmjs/4TStgpCFoK60iXxR
hitCwGXnDnhPwczzOwAkhgSr90DQtANzkIaScMVJYkHRd440diZ9HzrFD70ib7XsJfcyOjyrjK3k
/D7lgIdwuIPiNVKMwIsE5rMty8mPgoFNcncwAx9p3UngGU5veWw9KsrlViTL8DvyEWbOD20w6pCM
+YwGLXx3gsqo/4bUkn+3BP8TTWIL464k0fKGa3kLQA31Z47vksq1P5b0b9zCQeGBsBGabNSo75xc
Pi63Gg6+pfZ1C4AfWSXD3qpdU1ii+hXJVA1LsQocGIcfJRTCS5ecFAEekSgUEFtE2vm8kss0C4TH
3D9OT5MLPAaLSydhKO3xf7HSzf/r/0dxkjxXB3qgXQZG4NTcysWNJVieUDxHHuvs5UJnM26M97b3
OqgwfTHKjZ07YMhNETlmWzdxczq/LbaIGYHNTHA+yU0HhgXdZ2ocrsYEheEjlDwLEk7WRf8xYyAt
acVCoD2KP8IBmIYdjG5eLogFb+UctpsSXeE8uExJoEAndvBOMe4FcMHijzSyzFyBp/uV4w3mnla/
/kFKS+gBrGVfoanGSdEVrLr094xMvLQE8eaEkE0OLkfICf0oEQV16F6LPlGf2X/A4Ak4EhltRgAS
qZbMir7XBIbSpM3k7kRP0dCaUIAHOPbB4P/Vq2Cr/U/ERhOPkuS6BsJbClHUYa+CwfnAl74JGoTb
FLDxeII5GWjm4sM4N4N8FqPo6WZE8FjgH4UUZYm0r0oekGpwqZwvP29IDmvAIqHfm3YOTl5qvRHf
Kixz4eB/8NZkdXWzKf7Gfre1i6+OwrAn31dBoittGP6z0YU73OtgMB8Ilp3uQfiRIPsaDDX7r5CM
z3NhuNV0zVi1VPI3YIJ3elB2aBkj+MpwGCs8AVCXJpjmzV3XmZPF1znkc6iGjNoMOlvn6HZcfXsc
Ro+Splyej1tL7KadgysAzblVslInDkyf4juBvbcx7b4NhElgT2XyTLu04EK9NxtWb1fzB3tvk0HI
naQuO5AwiqNelqLslv7Th6YVnH/IYTgGFEn4LVIijHONdGUZWYQrraYzg/SoRJ6N94lQWYNDPDOk
KX0ecUVjhJ76069fDqe0FBKVswyBe/QhhretQzcRxfThX54pdB+ftHmXLmP55eAlScVY65thrBrl
9vs/7l6rqYznOZ6nS1AulgLicIU8tmbm/GDu+VS09ydLVOkda8E25IRZhitfxcN8Q4e9GXi0Zh2E
sbJ9Q5igpgGCVi5vclTt7g1TbdY+vgwPE4tNlDEj+waEQXU13nFfVjk7FHovzg/2lgXR8JJx8GZa
OxymQIDfhB0mfZQ/l8DdU16z0k/1oZiDDvZaNURDjOK8ieGTphUcxA3apZXOUOUrpWIj3NGiL9R7
lo4TN4HSHvG5zCynXLTkKg8MPQCoV7KyOnEaCbov9Tle9VjPw+xTfB4IKPnQOtpOE5FFZwuboROq
gm1NcxRXpV1HafvSX7p6lkF/Akg4Ap3X4AlpQnq+GozLg8e5fkcgzZvMCsShsPAIh856WSw1e2N6
RoXPea4XX0Q8owdQFjcG8nJ6cWSZ6Sqmd5u3P9PilYqC2pmMy8dq/bRs1lbCeKzZTv3GoOrq/nna
t37oF1Q4G443vJw3rgI4/qGX9jJLZygfF18Sb9zS5W29WyNQ0Dimqpn3svf+V4vJqiTfn7MrJnzy
Lo73t6zjK7BYKENcbCBmjAi86PTPuTT8PThoEVztSYP0OHgXpTZgVDMtFnIMdwbTfx+F3CTlsaIn
bJgLyG1DloUBFNAfrmJaUtcP6WJo/x6KY8KSUf87LVaI8Wb4wFVSRuVafz8dxx84aroa5eaCAeKE
MwZONiteC2oOq2RIeBuQMwiOLaNzuqskKn5+NuUU4+BOORudm/gymlkt49fNi/gmOGvuBilkLPBS
but04v5CTql0iVWonMCEjhf48dOqpL55II1g4niN3uw3vQfMmI/nwyzzBt439l4QIGRbwVkK/xGj
+fumZKp7DmVLNKDMBp6ap9/73VlhJuAnHifHyzQaq0GscuK81p3mfthpOrTjyhO+lL3j5wfInisD
4O2ieZA1iALw4yF6PJFu+g3sz3VoBD44CePB3xzPz1haiqXLWz52YSEQG3LaegYTwQA/wHVJZT/X
a/bLPltcpIDOM2URemd6ZGuKiugzQSfbni4Qf/wGpgwKTs5VmsUi/3y5IpTv6+n/FJ862MHIDGCh
nMMwup7+rXs50+lD/OUyNJwfZW+f7TUMjAdOd9fo0b7R5AlOPFTWItsbUhvGKOvRM5hhiV/Q0k3O
JEKa5YPIJNWdPX5rnFVd3l/GXuVxMKZ/8t+Ood5PGA8J0oatP+xef0AJrh5hhAk3/JpC8L5M1BD4
SU7p0kiiMzb3iOgiB1b9jyCz+KqJgQDDMZIFevxd9yYDCHeGX+dcRVYV7tvlNZIoEBnEAT21Iixc
nqQ/vN3DXZEod8Pdbi3U53nrvhIx08Wu0YT501ggIRFtFR4ppbinFgsc7/ufMTX99RmprSe3EuBZ
kOuAfTnCEAyKXv+K5BCVReONlEUEGtDsX/honX1NmgV2CsVwdXaG0cOj+C9EsceGsKweogq2slh4
buLw9jJHNBI0xFebiIruQKtSuJrPApFr1W3uzxzBqjwBeIU5BAGl2xCuMlVU5k7rszm8eIIYdo+5
oY9aCCtoLfhJVnm6s99jh+f6gPkghUP/oKVaA2mW2MF9CRC0DW0dl77gKRBAv4bzFvlSDUwfjVcp
YCwQ+JGEwqZ5eXxsDcKzdcxbR3s6MLLDbFChP9ie2EJY1/qOD4Ie6TGhapVE+I6OVxG7Qyl5k4k6
rHvBZ5rSISIRnX8eQGPwNhOQ62GHjARZCxnPUEZobJ8Z7S1pOtlv9g6kOkY+pthH3pPXvJQiKt+g
NwIEqyfi4oMOmux2/SK0kG78sCIlPDkv1BSKI4WdX4HHY5jDZgPrDed8sfREsGS9zYWWwSY0hrGu
15I2LV6a01QkQO2DLSxewpFvO+dw3CJcyfawq2TDZSicxOTff2qOjLpKMkKSmppDmpY/6ijSSVi6
11OSh3FD/iy7V1QBkJNcbJr5v0o4oeuNxRjrhpzHTh+zTdh3wAc7cbN01ESqX2+mfDBqGuzagUgH
j2NPiSepIBQDxAUI+JGPolWLEiHHvAM+3nZnkBPuqAbrg9hIZv3nMMfuGnKO5zvkAeJD/m8Cv3Id
DUnVITau+iMD5WlWOVwZ/YrkKxKUQFroT2pKVBaJl8berAMLi1+zFMZVI3MO5mI/lizHMZ94NKQN
WWhNFwaD8g3KwJsACeIP9Bcet3MN/Pzwl0GlZitDkR5uQJoDUfWtNhrCTHYkNlcrI491CJMF6Pox
iqm83zrTtH6JaMBffaSTCuf+PmRHUbxlMlzqeXyIA/UlTOyWh8xdLAUpPhdzrA2MtJbftCTKBD1E
LS+ADa+vtrpsCmPWbdhqgvhCrWL6sj8+4VX0OsJn3VKGJ95soakCFXrsFUzMBOYhI5vldunzA9ue
fZPOp0U5oSBwKDySr0C5jCPtWoxlqfcvpigNVBgGwCmQgK2uI86/dGGiebMnQR+zmS3q7nb78oXF
2Y48S61E4qEdNHsCHWL8HMLYBUrz9RszkbOSLxKVL+EegzzputW5O6KfmNIAJaX1NAqQkl2OaI9C
pYUShqSiiLfoMZmGHa07U0DzICK4pQqWl0TMGhX/OFzGyVUyFDHl4qQ44H6dlUOc5s10ILZwSCA/
dqeKZG1sfPsRb4mPoOH3e4YNHyzCQL648bDCqNMHQQTs4RAEHCNs2aEM1XozJpZ67Pl6L78SyGRS
U0EQsQZ1qAbcnWtBQriUnPx19x3o2qs0nIOnJKtJjbDpGYXWTwvURZqOl1AoQlkjd0Va74mAMBpW
KmuE6HKLvUDfbhLCdq/OuWcrIJcjGM1xITpqMx+ioZEbzXInICRRgDHFj1McOf7CNOSZKo7UdM6V
t2f6QD569W/Taq32C4rvwmJIqiynTnRoNDzCkoemToJapctOCzE0Q1HpIrVtujzlTloibCEt3blq
if6P85AJ+LAkq/Gm0/P685OqLiyYotMrMelvdLO2kQRfIlwjJkbJmjKHVgWNVXtUMlJ2iFUE1mWN
/GdDTd/pdfFhhCALkCqkX9zWgyXNntWd/rnRnzTlicwBbZuKkiPDYfBHvAX3VVesWKF3epzEtLZS
quURPYRfHC21G9cJMKmHLoXc2L7QNT0h8pn4dYPodnvTEykMVb2EtK8Rufst6yMLI/9zGMcbBIm4
N3wYZaISdOckMYescaTNMImtatDoP0Vyhf8CeuBnrHORONxCA5LNOHgA54Fr8pUouwTc7uT55eYO
KEi/YTIOboM0qNK+OTUSX61UCaJpkbf4tNsGNJn0lyNapSZnEQW0T886vdgSq3uUhLNTqaMmFofn
RKeONIT/wfqvEp1uOJAMheS+O47eBuHt2AgbiWhNemVmlO1nnAlMQ1Jlao6hmfds1AcUkEaEtfTm
oLAyubNPah37kPUZyS0a9uN9pBwWPbw5lGWU0TR5hyek9jDe6UfT9v/0v3Tg3SVeKvEn0P3oIPu3
USqmrhmJfhbbdJ7eU02qq1pDNgTJdcc1Jj2m5jLp7GqfDADJB99Yw+9E08wBvthvphITAA/ihNzy
Odt64MLDNmJEA0/MID+5xTL7iiKFWaK+O9tD+syIu/jbL/bZ/7gb1nVSeH4LA35L2KDdaJd1/E7W
/zfaO0FiBvwOX5snuw2ywndMZKUIyBfn4tT9uvI10AU73wL1KH+4TFWnPDqNHFofvjIBIWW18er9
ozMTDFJeffR3h7ora70vMGSFF5x0xAL/cY0crQNjn7f1sGOsoSMxZDqaUVeKpUnEp+rrbsF7Vn3c
l5CVsYFyv7RAIz+5/oF5CSOIGvKPTbas0sSn4CKIuMQmnUHiTMNCd7lwqVoJXZ7hYE38/LExjtz/
d/PD762zhqvY6kt3/lM9pQCQdwWGvBmiooeqmALB5BQLiZgPPKjMUGDriqiYzKujs0Nc0xIpQIFQ
Kdn6FhFTx9pYi0Pm9ikSzzecumL8vgTptIUrNX8uYmSRz7tscQ+Xw0FWewm9GsjXTQq9KtWHsCeX
RWZ+E0Om3N0qZPtD+PHCYa9hNEYYMl3P/AzM3eG8boEDgX/7vBl2W2qsKKLagfOcIfinxLW9XpB/
gjTsMeskmmTHbaBt/iFRx4NqNWMF6lmnWjOXhXimliFMmO/Nf6If2pUXlcvOsr/kal2kLBcNmSbL
Dz6LH7XKGSy2wUmAl4JCxPUENdkTVWQfJsccTGGNv3FzLcJF20PjRYKn+zlNvl/0WKxKed9Ssz4p
KTAIOM5DUpxmriixg5jsb6iqkMYF4vOZxGs2jo9Jsz2wfJ0kzKWT87pTGx/GyMnIZ3dJ29NXZ1WU
qCf2abeeaAjl7Vyaf2Orr9GSXTfwUz9/A2JvGFPpjgCA+LF6nhM+9RbkgG+7Rl7PKfD+HmaPnLbD
TgmlskBeAdFp/D9q2WDrtfosbE5iPE0hGeRYSwRXA6YF+vl+eu/tQaw6LYoU8MUcsUXkTHGBjCdQ
RM8CNI1J7Ocd5dO2A/NmmGSO7tMTTdujoveYsFuH5Jsoe7JyW/TPeFsQPxQuDBE1F1T9RBxJHfW6
T5ljoh6Xhrd3pi0FnmAdcKtK+ShuR5ZGn4yC7JmXNsbQMoVB/Pk3I9vYFEdEU9yWxf5gKm+f77xi
2Pm+8lR/Tx6quE7W3qPHvcZTpHhk+D7D+8CLhaHQEaDpFrmxkGXmIHRnGzBTTjOEUschlRkfKx1Y
+QajIip0j41te1BNhJcDHPrNrbicAYfnB7Atrl1ffdNM6iafoKqG/hmUPf7NnOAJ42kmbpaZ4vno
USwHkRlWCmavhhCUHxzOmghYHU2mNXvZbVvZFsYeo0lpKY0uZgJUQiwAn4AP8SWSJoaY8PIUJ2bg
lZF1ZeCdJUpK7ZWMMNpIze5/YLIKvxxFWxXK813bmVTFDy38S2h5NnB1bfQwsDBQ+bnKWD0wzp3i
pydKJ5YAKeLALC17DGEIBUC+dtAajD73puLvURiKVAwnFBTwFICGhEShwQ9tEqzcaTOww37gE6Ft
m/TjQJUh5cdKzlgNabiP4dx1JDZ5CgVQyQKNM6AcFpwJEOtN90vJFGIP6sMS/RnGOB/O98SHdfjg
ndzpCRIJIdafFF/2vjgbFUARy+v5JYUPbDGLalycpIWGYmVmOWsMw71rp9yL9paLxEHENdMAa6UD
1NweVNn88Q+kJubJcCrYYcCOiOG5UEOXW/a2uMZi43VF1GpCiX/j2eMkFmvwbGVsWONzmjzEnBdh
4yMZ9SljJ2gtOxqDVXyZX5j7CXBSofXrEboMnS17srScA1E/w143VMaeQKLB678uW1Z++HPFrqZu
u1heL/SfqQYUcqgdRbW6yB2klyn2NUjCWD1iiGZnt+74TPi5miBrzBEtcugwOYDIEO9PUeeTgDlF
IgsZbk6wKYqQVmhoU6CiyPHVJa1epYkvBbVRRPHSOoK6PWth84ALjOK0n7vfSW9ca/rEXZ8I7YW/
mFHKTb4kvaGt9PXFdJsZuF9FgxoMmA2AZiT7AxG/U6HOcLSq4zIDtjXfOKco5B9zv4wIC3dVeY4g
wzrU37bImpVS/V/wJlJVJ5rgI4K/yX8hgI5DLj9tjqMWuxml1i8gW3IzsxsCl4NBhnWtUVlP62qu
twwVw/ypy/0M03flT1HM6dWAXrPyC4i5P5tARhQML6pTZv1VPG4cvXOaZsEs8QILfcfb1djqZypd
VKzh6w9fVWtlkrCpG6zIIgfl4dqwV91QFlbJtj9Zxqpgb8KXIOpxMElTjrfUBgDpHj7wU4MI89TU
mjHMhPVaGxYUH/92IBNIrVtvsWEJJKiJI+Almr6i8YMMmiXNsZUjTg4HU4C5OxfqYMtYlCF4ngi5
RQmF9Jo08yWW8ncxbslL83JhDMojvV6Pt7gMU+kU3rxnMDo1rRL4SEMUJKaghLZlD2/yFlMIkVnL
dV38AX+jeIbluzbiLz2Rp44a5+ZfXinoF3n8c1u2aGtJwu7bMhPzft2NuTkT5KoymbBWaKHcS3zW
n0qIQWf1u2F37QETgpnyasJQVQ1d31plACFS55FaBIdkcq7QLiYNn4BZ967U1KID4thmruiPi/nQ
5i+9Buy/eFAg9L9e/YGHekkkVWY/rNDEAwNlklLYnMVfQzTQ1CSGKA/itSn2x2h4qND7niSikgBI
dwpLx6358l1A4KWLBjmOXy7Q0AHALCafVPrQxVfK7UYYsMR0LJI3N3mLC3Ite+VDTeN9pYBwHOHk
GS/PgbXgUucll5ctaWV5GDMp8dqK3xFPGVviuSbT7NtU6LQLRVHaeIZsTSwDM3icN0qQGtLi9l64
YaT6vWxkMA9pzyQgLGvycwgHAl0AQEjnp6T/8d5ILR2cGTK9sJr99wQzMXYTqyWs2SNE2xEJIpnD
DbXCFAC0kFqbZTfGPWQ+DOEfFFq37Brw4PeC7ttm5QVZZ45rXqlQFgS6PgX4zOIBPBAcy+tRNxyi
mWlG6VioQecjrTyZJreowIKkXop/0IXd7XUctCjDZkcxSoMijT1uwx8f/WRHmVVQk4ZZGEq+5s6O
5AMwdkAJ8qbc8bneqPRtnzhLlQKUo5vNCmIZSLt02d8SEvu5ZyY1SE8Si7ibpF15fe0oTmInIbz0
iBbinAzQpf6uZr4iNouAO6SXPx7Kfzu+REL86I7gTpR3u0Bva9UUIwu3Mn2fLnW6PJfLwO5720Ih
AEZcdu9k0BLUU9iKLifGlst/ZoTrPQ5uuMPQgdwudQg/5MrJ8D+RiIMJVOS1Ex6g5sQJuYqjv+nK
fbGJ6nS/fx+NotsTo8Hc9zOGNHrMcFdDh0oYrWnRFYOTm27HLvMygsjtliCKqjUGDsyHqiaHhwN3
qNfaTGxs49OCBtknoYUXXXx5ERbblFwh2lR9GaKhupRssoGeyXxXPDu5Tg0LQJ3YAiucoyGCJxts
aiSLtpjIcrP1p1Px0kPuT0i4xgap4IMMAoG2xnwYQMLqASGSpycU9Y+6H65BN/WN3VrmBE+iYwmi
IibBMifZARwSnoqNLfUP1GnrKWRXmQNCDVZP/W5IIOtrKJzB8iwhDXTn3xI56LNr/jq0mJltcZGP
UGS7+BH6tjwkur/BQcqcbqrF/I80UU6BsIAMtB8HI9wKu1KmnNiV3vCJDP7zsW3arIeNpBfC6xJ+
+DBz6/YfMVEyjG5nqPnt/i5YZvPYHny9P5u+4PEg1GZy9yR8t0KPqJnv0la1x2buNDNljPo9ZGWR
IpfwWQOWMs5mFlNpDgaVoqqWW8Ltl1fATPPe4icVIfxghHziynRoOtGns7AkviPvHPw4WwFcpqpc
5rJY6VVmI4CV67+4JYrrzawzmGZT45wB1wQGxUmvJwmaY6NVcou+VAmNbla+Hnq4vlorgQGEHApT
AtYhk4uoBkvVrC406TbgKy/J9V53mrZoF9ZcE6vluS+XnafeG/9LXFPHnTgO2eNOOVL8JlkNsDIv
Vna42RPtIr8BiUwDvJMkJ6n2uFOxuDBHWq0JKlCOYau9ur6rYkpfzMs0ARSieya76sHK/gh0iO1w
/hUnwvDqF4rUPbVielTa4fkLOpiaX9gNmzkpe2fVRmvoQNMvOXGTCry5TcdNMDIKzTI3k4UEhNtJ
UDyA8Xoxb2v6ZljWy5lZcYqwhugGHt6cL1Uihgv6HTdLAgnvQ/uTJAWE0it8DGjVt+FzdsgaQiTl
EsmxPNa5TvMIucCmJSBGaUaRp7zLtaSlnjA29+fzddwQ5AsnxxfnlBnKS5BBUyKWE4MDkoi0Bh54
b8D5QXhkdaqj/cOKn00l9lXW4g7YKpX3t9ThS6U+nK6UK1G2axW8u7/CVzX6I5J/CsTxkXorbKdb
Ain2+2k6w+F+YBd3AIELsqNnwTg/33rptjIuerfP0bZZJB9jnB5XI6+Nw4Y98KsALiaEbcM0EVZw
Y7wB9To4ZOmHcl6p4STU8PtjacjgsBP43SiGNEDV2xn7Ujo9NtHLh/0zOhIHoq09Ma231Slnbqhu
kmG76Bud0K2r8KQZ3/84WT0KmsxtZHLpvPR+WiWn5wdkBE6JM1w6Dcy1PbuOC3xTT0gsrfiH3kr5
ckNBHFQX3XbsrjTHMZF/dUih0OQjorDlyxEg9ck9R7wTFDL9qVdMN4xZ95gaAybUmUWxJ5YVCsc3
qpDXQB18yGifMxJfxnB6WljRf0Nkui/Fwp/5W1AkqVNnNYHFDsjIm3mFM4pt8TqdYe3qu6WFbXok
NHaNoyS4Ms+p9w16CdakhXECt27Wdm1ayzdFOwAIUvH+0KT5sljqCSEb5Rhm3UK7H43i6sWN+Frl
Si7ljRlyT+F20/sUKu+PtYLipw7ji6+2ub1wVOtNFaWnIe0+BHlPwbERVjWVpF4QHvg4xS3NmYUG
2ul/PVO4KqDRGrBjC+CEq9ojQLiqfsxcQEHCY47qLtPXRt5/bE7zBqo92ajv/ee+T5wl3p6IanaO
xHzXaHbWta/lSJ70ASLwv0OBa5wjDbHzz0UInmg5abbV4luQAF2g4tN3PfF451YSr+DfV7JF3Tla
gFXf6Uu7WmZ0f/qV4X5cBLgg/q9TeG/6XXtcZIWg9y9BLmEegVKZDNPDZN7TlyaWAnU0JVD2UXTO
qII3+sRdaPG66gIdFmaHmVuaJO0Ixh/uZkkt0PGzpzREoQWN3UEJLsKtS72C/gmxKbGWSmMrr1m1
+4eyCKgUTAa4Ejxkf0v3Kh0+FhvAbNy1/n3hOc69D9HbU28XvnQkWnBRRumYakThu+dO+6DDhXwg
YQvUch9d3uPOMttTlBI8Y190NKfPo51IuiunEcMCVZkQiETxws+9MRLUlA4c6TWoXiDluDNxe1Yy
fod7tY1+mDRzS7D+3yAcdqDF2KY/jT/OiIP2IaKIRyn8FP3H7UVKNp+Jln8kOlep6StXJ0G6uUQX
1lNtVIRMWzE1LljPlNjiOpvjuHNRdGVEHDgIvIG0m9uvLYXCSTE1KD2ovXSw9cLGK2OWlfNqEsI3
YSTXnKHlFMrjBbVTphsOqHnzPCgEx9TOaW36IQbWsWHGJ4Gsr4sK/uIfBk3ZBZxaGzb/MSzl/U5b
1w7DdcmHyUNWNZmDw5f3yYhSlLku8mH90uNm9D3aI7mIIPEr7V8CV2q5rFu0Uogap33n1rUQVFEy
MXOfcM7jnJvj1qcGxJuFkyYuLM31uwVEoYuGSz1sosiRFWBd/GiAu7iwJYv5xjgp1UGdM1evUyNO
ljYCjPcqYpm93z5KuP+EngHphnELidVuh4DA+DsFeda492wrbTSCTP/qG8WBuyI9bVZFBBgBT3w2
L6X9S1CtJZc4DxZe9jrL0ucKh3sAM1YjYsBD36Ij6UaKL2oZYyPatMNyx4SJ2Iz+/D5j+Umqa/dt
Uod3iw8o4kc4AuVEnGip5rkkAVhMWESXMLIEIWB2Q1of4wJ17bd8dPpqv9En4UFiyxRrF0puTU0K
mJJTOwSdDbTtIO5hMLLXumfYnT20zkca0yi4CgsP+mSZQ/NaveSSmBeYMoLpvkxyTJEwSWr/EHHp
vjO6ouujr1muQ2x0Jn540SejVJk5RySD514zYwyPlKL0AeQOpaFQXFup+Gc1lLErJMRLCYM5CcaB
f/uy48EPPoxg/NYrtmaPOl6Sh/Cqv2oAN9Wh2Oi009TOwEJ6ni6b4ImVi73FhzdrFN00AZ5GELbe
uxd9uc2p3p1diSsXlP24PnDTOrewjkC6sKjRchNCq10dPgac3DXkX5eBQ7Cwh7FQJnTdDa3Z4ysZ
rg3QOORgD8XmPP6k9uE/Lj/D9SdvCBQ+lLiG/nclQt+pZ5DstYQwLgWo/dS4nhjUf8lkZxAJnd9L
qiTO4iGvN/933kBrqqZc8NnD4xIfn1JB+tPBZKEzuBFFSTICbS+OKzFALktXFCUKgqTYLzo/rhIl
fPIeWx3Ao+fZU8ouf44udX4ASJ/dC9yS4HZ5arB2qv2YfeKvCovpulyyRjJF1JeWVk6grfOapRi8
z6WVslxiortmhLbiRUholzouEl166uSVoeYolcch/DGSQv0UPTE2Yd1fXB5klZTXJMjLBy1/wPS1
JNvnDZhhN48kbI5hM3Jm1RYxqFWEJTpXukyHT4MZQej6ht+LtuQfmAw9Se2D6DZsAsfeErUI/Yuh
uNO0e5eO/c2FHFYHJc7OOpVOVS2QXX6PTrYeGB7xk1y6r0xXKniYxazas4K90RFP4pbiEVsBkYuv
b7S6hQBJkDpJEYd6Dr9/PqoJfbNuqMAySUlKYP7Vm2tzIRyo3QTNbDRCwE17RmmU9FilZd7Lgexl
XJ4Gqbo8uVKAEUQYcgVJJTIxD9YxUPcbVzGrQAfHrUGcTNv3KUAQaYGk9MTHabsFsnFJwlbEIvW7
SYFwDpSTA+VbF3wbJCHPl5PGAeY7BJ/L4p8NjJWPVHZn7QAhb/PdFU2EsFgOfv3OSb9w2G6GXOVl
2Kejdjc+ycgMGjJXggi5zsma//8/sYNKbDadb9JGnLrp2AaE5YfScMUBM/wJyN2pSjKlSx8VgTzh
llD9hGX2eLnIiyoXIwXCSJ6qaMbm7r4G5hd4JwknU9v6w57z8SSHhgOX3JkQo6oGCmJaDw/Pt3FZ
YvJUWI+7pTYV5D2uPvc/4CY7i7VDkbgrFDu2xT9Zi/WORX+XZ8C67VvqoUpdOsDKRfH/b9S+UN8r
6avYyeUxt1rN78cqDb/GfYtsvP3ZNErdo1HjqzzFTgl6jqeTwB83YuWJnSnvotdhG1PJQgFnlN9P
Z4DrL9mthAdKEs7e3Q0uewSgFrG8JuOUjDXqw+V81AEvRJnyFILWtjwbuwrbQAzFzmP1xZhy8bRz
ayjM+nVf5YT5wO7Jn2ekOeqzx7MlZ5MbKkdPAZ6UIdqp1xwrmz2HSlFcr2xWW0sZKnA9EEDSpR+A
4BYpQnf79MEkmpXfDUf/Yk+PjMtecC+ckFDJlrGG0+XL0YiKeHySRyWCsXgQ2ue1wKWDxcLKYQ3C
lxpKBofQpSSP5fDLvTyXMk4wejI0DOiwHSV+e2vQYpg+JGh7ge3D/rCtfkV4zgvtB3pJeGXJ8DtK
aUywIaXQqR8NEVHTJbfAgtxGAAwQnb2PeK9zxyGU5SHBtWcksPBOBD+r6WCiL1aAh7F0ZbvFNRce
0+I4D5C8KxXruHFNADauT2SXpFVHFiQFcadzk4tXGjIlixtBcgCEJTVCk/u+AuxQ0/9HJtDYKEDE
Jsdf1ymktA0dEhPRU9NUmZi45aqoUynpKf0QPysYz7v6BRm85pffMjiyz50yUNMCiabC8KlXJ3if
c6OCWattUvm2LIduR33Rz2+WZqipjXk6zjg2ZJ3AzUBtIk/f+Hc4KE+MWn1MdqWOvVURnLkwrgm+
PEFesw+ikxN0rFC6cIp/1IZYvs2m5/s+5fQAT375+0FcvCalp1Xp4Ja1PTj2xqeU/s0UHouSCYGM
5LlyCMIRO7qi+YN7oKR6gDprXsPmjWJ0p0HclGHcbnZGoC9N81YCDL50MZzn/FrHXh+bRI5ZcEF7
8qTlFDtE0dp31rVBHuem8oiHpDAeQO1ztCiSlfmB/9YVVVFWAKQENwxOx78B+R6LRqAUzrD+xR/c
u1uIPi8xnTOCoZHzu41CD0Oqv+JPSK0ygrHYnXvTDi6W+37VT9L5akxIHl3Vlxl+MjMNi/OngGgh
ncjo0nNOmIsQ7iRhUDbZpSm9+oet+rYdKh7ICekwR11GEwvNRYalIvn63zFvgkZ03QaRm5OiBKhO
ozPkoKMrQfzY9JtISnQF76qkDe6g+OVOKWId/cgZla8KoMHdXBcLaP3JIa7hlyqeQsl+YtQpNuek
ahlbSarV/BnaiGHmNB6VuVKHjp7LLUCu/BCq7IpRTHPXSGG/XTDdaOK9QIbxBfEjqt5HrSKvyhK7
i0l6bUuuMWeY8ZeEa3+CZiGMAXgiEhCkPqynzQg1H9IT0S7qzaC+cCdJvS7P0nz5XOwlpQtPg20a
dGzes0BFVA+cx+RrlFABJ+BM230ZxFHVap4bkYmDgJ87k20pASLB2CzCjRdFyESoBpwUz9i9qjxH
AWV8HpJE+NcVQT0Ld2NaLTYfJu2vgxXRBEAFqiKE/TaXPM6NynPbL+429mJW7mQK8906z3ZZ8Z9u
to+WP8z2+SNYYfzibleHIIaoljyompd0jC577VGI3aGIR9BlYH6t0LSQBVwIELxb9Dt1AGftWm+y
p11lnAdOt701VZdkjIQio/jbksdz7H1KDNLxOHrQevwLqwfPEz3pEyMTxIxPvrpXyGzqTBSy7p7j
WBcaZUGk+o2jKFjMCoJT2h3fSXwWUI07iiwugNfDFbGgbk4/9Uz6HuBDT3CWbQnCA5OY0qn9drwB
p5ZDoA3cH3EbkY1ilGCcudnkbIqTF1MEjbThUZTnFYcSKN2+Z2LKxcRNB8kpTr6q334PVKe8yU/j
anXTgJIvGPP9TkqEn+9ZWH3UApOtZpTOP/T0TaidU7oK9wd6k5s48We1IwMC96Ep233yLlwv22Z0
Qoc25gtHd1U/rCRfuUytcNc9dCz9+dQYtDSm8/Z63rJY8xrt9UTVRLL8cBt8O6ON/a7iKLGNQRog
nXgXE+WG3vgor6OX/4eJp626Aa3WhDpdAqphZsVjWxBKyYcjoqRr1i9iHugZ9OtbmbMMf3I95PtY
d0eAo+EesIGFmzcVH3FYKwE6pMkLcw/XX8TMnjPbneCYGkqecyKkU/F6wULS0Gn2oWITJvxOgE1G
gr2RrpngqhJGGs68UjnPEkIE1hQxD8mggQMm8AWluJ0hJ4G6Ol9xzjf9LFkPThyevMUmv76ihECN
E/3k3Aa7OvE88mJnfSqYVhT903vITgr0lDln3LXEl5AS61rK/ISFWagUnxXNfVmSlYIUS87/5j7K
9u4NbWnkixq+uD5Hyrk5Ypw5AUUndVaiC2LhTB1qk76PLouB2yYoqeyl3a8M2B9vN79TUZzbJKFD
XBQq7/YM4Q+UypglyPPqhFUXrTL4OwUsdTCcriXkFk4hE2CI+nB8rOK7HxtXL+Vh/wZTuFaeyuS5
7W7zZI5FKzZWiBpVUHUQ7/tYuW8TWq6HM3kp+gatC5QElKGaHNL/H09gQHA11xZhGuayeOoxXfEq
1SijKn7Br4LuRXpMeBv+8w7lWgib7KxjLOgpZp1gIWWOARsSo4adHSsysFZH8q6GhQqlrloGnI+X
UVqIVCmM7uzgRMZcVC81pKhtnT7TlAJIOYflAUstOuBLMzIzuYtvxzRxr4gLR++LCoBRKnTEFHGq
1a/P/CNwHhruG86+BLWJP1bbvQQVlEQGyWgSfae31L7J5naGL6yHAhOLt1ON9uXfqr1i92IyK/mS
kp8Kzg6zAdog6l9xBcdOEboFD/QdwhSsOBqTlxFJ+88dEnMFSRET9ijd2iXccRQEYzj+ihG0gCnx
ZBq7F2jAByEfw1kIEUZcYFVpWOpH0Y1qXQSsbh8+uZVAfmIECO1/svdGf8P3IFqHpR8PULaO34ht
HqAjQGO/ohWf5ZwtDie2e6WI57diMVX+ZCpCHg4Zws9TiHwOfKfcT6mGL3eQ61hIOs7DHIVhaTK7
QX8/lbu6TyNzvQK5kFxawVLVCRlJ6zeBYuyKtTXM1BKf3LtlysRkQl4qLvZgIu0f6kkzBZ7o+zF8
G6Pm5xxWBCUhgferfxNV9iqLYP3grlt5bNFBg29Jp30EF2rrlosPvSkXiddQUcddR0ey3dhAyx3P
tvgSJb4Ylm66CsOIrPKEY5aQP5YB4cTfXaE0v7j1rX9IGfce2ayRQiafdb/cEnaoJ+CNOnVkSg68
F0JeKDp8p/yFUSbWTxHUEFf1dtnXY22MkhP6kzKq0qFvPht/Ir7FBG64qyBNtCkNCvw0Z0JoQufj
eDpB3kJKiiJlxSut2kBwTydY/9ivGQs8LNWDMHjTV75+3SgOc9/SJV0ek8KWXCKCzfTuDgLfiHXy
Drkn2Qxe8BfXuOeCFvLaaJmwXb71eIuefz7D8AD4iLzrgEmYmvenpu+OAcnJoKHCnYOGh5h0Oj53
9whh4JNf3KfveY+rzoqRh0e+ZEBDKPHNUVK5/c7Jb1Tmf4lB/6ettGKf2ZBhtRfQdOBd7fuhJtxk
ws6RZXrx53zJvGtJ6V7zZm671L7AuMqPreoK/I/uOoi/MOhh7yt2IM6twtkoD3eBEf15z9h8nz49
vW4IxMoBXkCpwUnZEPYjPQr7BZvJGunbnF7skGRhXv9TZevuekqtpoe2eiOYowaqtq7QXdWqTZzN
ACuSDTS9Je6rljpTSE+U/oKBkT6tMV56UWbIRuGsDH1QOQvoY1cRDxQg4rnrK6Z+08OZK73QiLoc
C3qXZwvDTXP1UAXXIN/mMKTlUYoAC5yAKiOOmNN5W57z4xRiB7fL1Aoac//Zy6C18/ZCpIk90g+j
Y4PLYMNW4iNC3hLyX7YIGwFIwgjuVdaKG7cgzBZCr0KPJJ1Z42VG2iE9vepN7tTDJJXEWP2CDZFL
Zh/015qjrwd8tAbiHztRjpHevYY/TPslJ2aFjHIXtuNuDe5INAKS5MqS4vZcO+EM8zx8bbUZruNm
ZrWb6OrpDdZblk/k3vYzDysCmJDFDBredY4ViffREIJVlP/8riBvMKM7Y6SOpG5b27Np9PFWolau
fyN6B3QqHmDyd/fIfi8+aGk75tJSNfLXMpZ8z0C/hVhoJ4U0QZlWDlj4JVkeOrtvXymxLE2rFQjk
8eyOAaG2wrme7cg83pxtFP+rSSyk4l7yH4Mwew1RMcbbopu3YNmdEprw0Rkks4FiJZdVT6bJGqT/
rx5eH/D6vAe3+LD4B7+U5YSUg93mQjBDIywxQ8HnqebRNfyQeaOzYTJvPbjWucw7DltR26WV1rLV
sAvashx5D7y5dyiSlS7RueppcqYHsT6OrHdNU157dPwNXLzupWamDLcnsDZc52tN15hHannrlg/S
aULV+GqDqFzG/4AAkFAAd2szDH5QF7sbp7+Qdi19DP9bL1ZN8C6Zvbx/mcenM2qpyFmGX6mD+4Aj
Om5yQsMi2aMnWrFQjJU/0PUiKhW1oaZu63qQUpiMT/soxdO+4SwmcgMsyNVuNknfvYELC0ozhV/q
S9jP7GTo+41DRVi8RGRj3qSRq/1zTru95brxiDRKuew9f33cv1qRyAwy33po+ERGNwBWElOoO43e
UayJrEmwQSj+2cCXLT6OKOljMYDwkV3NM4vTg0vn/YL3xpWCwz6+qM0/DUUZYMpUE2xlFWHWH15J
hi/AsTdttn2yoeEZfcRnHY2dHla+kB6Uh1DbPBL/u3raB2BASzflavsksX4kNiJsgCJZBftyA7Gb
G9YcvDJUkPSWcDC4i5dDyLjBLETw79I6+pB1pPSz4bdAJvBANkBlTkyoK7VBnuE1gPJgoNm/3WzZ
nMCMCU9qLrG018KcDYgnOPNX9ctVV7eryz7cysOp7JQl/YR2mxqx6Y2fJEqWWgwgwc2S1Ar1Iis1
tM1kEz1oyaTzcGDOdczh8JH0Hv4UHzchB6qZItyvSeh65M5cyBq/JIj21/AFDc7rJP6rsBXch04O
2o30WBtHDm9fQ7ysQJoJ5PsLnymB1Jod2yYLEbgC1QbLMsmL44h9gOG++wPqhpStRUJMSUFrlwLD
1DloTWzuk6ObX3fzTo/4UQKnhO7ZL2o6RnJNFckXzh6tgoeiB6ws1y9mDgF4FMEqXOaHASC932mC
MsDnme1G4Aqq5kf7m2/8M3E15dKAv4qWyduoFau6BPGJ5s7T6JF9gO1vzSdMNV04CiDqszyxvkuC
BD3YZzQVIt11pUO7zdnjDzXvt75ZsQsxxAn5r5i6X55k+5mKPd6DJl1JM5aVg6nu+IFA+qPY7Wzj
PNwFdT4+xCj05/LQovV13Mmfk/UT9KFcFcREcmElzb7qqGl5ebdJg+NvaXJLciaOFy4beriCPHyz
XnuMevy9OcZkx+BTKsVP86vGR9I704i/exYqrRswLmGs2Bb+JDdMECKU97qPHnln9kSqhxuL78ww
DLwMGISMR7n7lg3l8U/VRsRiV+scVDconRYjYlPkX9M2ruZwUHNOdHWVp7Cp9kN+Phmp6AbKlkX0
ltleL/AHKTleV59mZeYtlH1EiA0OPNfl/FF9lCvWXlh+nKl2WOVn65hBGRY800bI9KyPKPCqMW9y
kDSv14Vihf6FYESKWiJ7qDUddvZbcCvkv0DpaQ6x8mRaziKvp/zyo0cagw5HUvWDJxfS2fsR9p5K
5Rx3Ks6uiCDVodV++QVkgqwbW6XJPgIVBRhJ+E9Wy9T5y6zThgnrhmR9+PDCZ8Qetiyah7bE6g97
AY1j2QYljOojHAUTnp8rEHKDVRSiwKyD+UjvDVmSWGCxSV77SiBxm1lIkVfMhZLLbM5qlfbYj4o2
Ynwes21cz0zEynpnz29uut+G0JgLvpd68bOc39YUErLQjN6s5he1OHm++Pni5jsTaUwcgBS7u5M4
rrEjKmZuiyt/yBKMOgLUey8hSCZ0oLuljHwA6aDIKTwudYRxDZvHi76gVwSsTszLh8ruwecfBG/r
IMwsrzN1cJ6ysiBbMGUm6Sam5T+Kwl1U0/g6qvBjaMPRsTwglKe0INaw+zlWNmuOSSj0zJ0JEsCZ
DW9Ne5FFLetNR6zU2L9IqtAhxOUnE3CnHTP5L6WG7BaRSJCpy+hvX4OyqfuVwZL+4FT2CZHdnb9k
vXLcFyHveGGw8LS3wD/jhlVn6fG+uX4lzSDHzSU8pO39fpq0KXxZukrcTr4Hieqm9ijonrb4Fk5w
mu87LT2d41A38Xl0dZFBGL+l5wKaeCp7I5fRJmoRDIT1/9ZHwxlwiMkcsqhxhAlUWgfmydSpxBot
xvSCPzhTdAAzzd8JRDQLc+MrZef9p5gmfaBY5TWdoxiBWjR0kst8aXCU1odUi7aeS/lix7fsAlNI
GuXfqKGcunBedU16R+Mac3AvA0jbcT0UWBAONECTYniNRyCnnhB3kTFrIyaKBxhF3fZ/54ZtqZ3i
HVZLtp3wwzNsh3fBrdLWfbQIdeTNG3urKnYDprieMqeYRg+y/yTMtgA1gLZk7ZyVXENjwdc0LLuD
GW8zU6VM/9SPT6GiexqK4r7c4NLP9Y9Z+KzD+g92NdjUD9NPje7Mvcc5DC52cdbODCTh1nesIhKn
MEyufF8UBAT25UBzSFB6YFqz7BX8ap6vNiyn3tWRU5BjXvBhXZYEeXCy09+5CDGO2t0xn78VgpQf
i/5US6LcNCEgXd39232nVf8KrR/w2YK9Fsg+pR1ca22miXr+9ClR3lbu82uixNWcIkxI8redwvFy
+EbNj6u8FSgZzvRmbHhzvf7PzIUMC9PSqtcV1YM4QC5ffGmBXwrqmPKB0gIsE167GG3tbmOV1wEf
u80F2QFiBc8WX7ZhWAfMFufdkeUetiNzi+cfTbtqUyq6RJMkY21o847e5eyHljw7colCtx9pamOb
Y4Wc/1+6uDzQ5dxdXctBlHb8bPGfVT6qdMNCtCXaXbzr96C/dy6U7YAHSYnKP/tsOyx74GIyhg21
MFknHIlMF6OVYXA0Ueorn0Uw6G4kqcGtIRmgsCFX4Fg6tqPGojJjwcBzObwiG0lH+0ivNDRkRFlv
5IJa5sUimnGnPs6jn7/iQ/OPT0Ild3T+r699S5oDRCGzHrNY2LYLHSNGTnu27DF2X/3P0lM9JcCq
k4odtZQbpPzhe3UfvP/ukVTqk+WsDdHFLG49cyQLIAnYv7ZBTjHCqTm3asVou1X789U/wCk6RLJb
ojzeN1edHsA29eht+RGKX3Bgzn1BdxpW24xhicV2AQ1YHxkyIS1fJV6GAg3wXf/5lBogER2VE1in
fzYkRcqBFtqTchQWVtqil/dkr+glH7h9QmrF/b+m89+a08OXBVWJ6pMGnN2LKiKtp7cqauKNUTD4
0DRG46MuT6u50U68HR62v5n8/u1Ab/LHa/ozl7Y9meyR2V/M9Ss9EfGb3j6WKcpJUI5vacaryW/T
y6emJKITXH0wSLkQ7jmt52lL4I9TfbjELgs12/kqj85NVYt8ANRHV+omzwzzSms4tP+jzUL4SsNX
1Nok87ARUQZhbLaOiAM/2W6B7adu6du8QI2AhbbJhSFpK8HjyqGTgtw5Kjfuhh2bJHguokNkGad0
2luxs+moBAGVygsgyQ7IrnzUw/PcbCUS5OTVxqQPqUvBk+sXYRC5bddiPQeveiZdivUNayvg3Xzx
mq8lRpaQ2VQNodfpzcrZ/dmhbJ18NmVB3sIRum7sGk1FnzJ49kILH9cTpbH4u7Tdrqe1x+x+yKDY
IJ70+4ZLx4HBXt/Bpdw04XjXfCg6Eqf5R/Ofczj/sz9WLuwvG+qki+3h5PPHdQlMHb93LM4BPjtW
1IPsq9wik7Nz+WBeOP2IZFCwg+lr3wO/AIPG98yUc9G9nSoMo+ogOpoXExTE9bFMVtOZIQuNBANr
oI6gtLdsiuhhePudJIR4RwQqEW6HWm9FRucRqHU+6NEsMuPBPXhXY37hKvHufgciC1wbQOdygYwP
AKLARc2vahbBYDnVOjDFSVpyi7MbwAHLlPl2Q5xG+d5Mz/GZVWX6QRcaO6992rokseSj+Z08GXWL
IUDDQxaY/2oW43ti/F//dhooF7a8q+fFypcA6XsDE9UUA0ZF8T6IOUs63LHZmDZ8XOlypzgmgz5K
4cAg6iRkO9snOOAmdIhJQY94jaMp7R0XI3HBuhN7ZIPPMJgSP6SnbYe6xFclgVXqjWgZ2V6QUHZk
mwHEMPeAYG4ti3AbntW46D3/6pTpBFSrpmiDV0A/JQwhAeknwZ+7pMPKt+naXxwr+3TNOM2HcCVX
vEd63XpozBQDmo+3s+6ei458orfWb2WO9FE6s3TTwbDGeaqQr0Nf0J8OkCk2Ypg9hImAfXRxPMV4
wA0Tozpy6wL1ZMtPYzIZ5EleUSoVBN0OufXeq7HpHHsHQmQuSzsCyIoDe8lPjx5YfvhGsfEJT1yK
5Yh30dnchzOJSWj0J4FFyyTqVdLrmXL1OC/RFgAurscxkova/CAW+y1ukk2TtKGaWCl9ePN0XPPe
lNIVyHsdMutSKzcSpDtqRlvo6iE4yyU0iu0aJxTMpelSDQl4mgnK+rQxhhdnZ+curNKnRjt2taEE
fKWT64jCprXhcoYdz9VTc0rppYIE22ePbuzpQtqf5KFw2vystXTrhSM8AD4XZdpQLutvC3i/DqvY
6CN7kYM8+zPZ6SnojUs70+F8pAwLbGOMrHRuHb2YqiI3gIy7WiCi2E/Oq/ugVGAtlwrMwaSEZrx+
z7hegJzuAyFnC9EshcL/+azXG+alRj7UcB40n4aR86NSjCSBgllpTc8NU2eP9JGSGopmvxuboVwn
Z/x90q6Q15sBVFRI5Ohbhzkj7SaeiSOnXA/K52WhXuDaBu3Skr9UrbfzY/CvDuyKKrgRliBcs0lV
O3/WRgGLZoRvGZjLnd78Q+lJuAfxtWedUTaroLinFDz4KUNPCyZLTi2Ml/TS9hysrehhsObm9bYF
NGZlptacDLrj7cyCJ2CTzPD5uCLfKvfb1pbGtVxrJxESnGjXxchbL+bY2tgyCqvfbgGuHO8SRVi2
oh/yHWlz//JvaCwR/Krn8Y5A702BzQ9R3DYxjQsZNzb2rg6kCXI96kVOXLKdR2mSJqnwyfNpEpuP
uT2Q6AWZixB3EnjCSWQJ6u/kfB9lSIWJnRcLBxCfjuspl6/jb3iaTfJyQJmRAuLpwLkqoRrmlB5Y
vthYmBWv/+/K6yEom0HT/n3swYbgYBx2i32cSiakBnBCqGdXMhZBbpdSaJkaRcueTsAUSjgeJOt+
sZHLRlq6hrKCYen4cEHButrKw4IS1BvUyk7hFg5V6X5GQBOWzrtZjMaltuYywUK9vR7sOqaQCqnS
c/nesQVKXLqcVVJkB/CqhbUjQAbMnIouObh0WYbnegXsb+OqMKefPZGN+7aM7ott+c6gfL1TwQaD
nM9eh7yzGedonxIOM2p+UKIaZl0wDrQ7VHmh2Q8wj62DQvHbl8TjOyQBvYh4IDL0Jc/7uKvJsj6s
KxSps2DOFNi7cysY1TmtM+roGrJ9K6/42TVMlkpnupZXpmdqFUpSfR1VrVGcXB5+zu3ClWC0mquN
+hCHnNQL9paY3ODPBjlhvPNCxCBUoqYE8PZw2a+P0ij3LOJDU7vGY4N1emkINSYeHY18LtCgFmug
nSRlNctn3kOeB7Z3rbALHgJAjksK9yMCoQ1gtKPe6SWR8p25wdtiRAPP7XE70SMYT6nDHLl0Oj9A
JhA9JnlrbSEWQgY5GMKz+cY/T5ZZNW1Qm4NNLoUfbCY0fc69OjOQRrTQDPukr+YeG/Kf1un2x2AY
J9/fywYZ9DrKrUMNWoLYbTVVV4Lke1r0TwX2dMcRX8WxDy8VwvjJFgDA+92quRrfgNL10wl8jnKO
szth8ggfPFqLOR9joF1bVLWGFnXCL1GwXJENKDA/aZBHbFpTesSx16OemfRFJghq6JOY2xQaHR8+
/dRXYzDOOPxthaghKy5gJm90WYzB8+Mm6LLn4XJ/rsInEW1cunnxprWl5n7iXi05Njuzr84WFVHM
o4mTKDht/FVKMQRtgURRghquqejnloHIgvmgvE+XlFKZsZgIRI71YgFm397rKS2OQBCdBRGtI5Mg
pxMaAQF4tbqP8i5nurbNMWJHTOCnGLvjBYk6YadtK56t8vPdvveOpPpRP0rUociprKW5YI2NaF5p
PV/30+r9HP0TlWZOPchhspQOGB5fGi8dt8Rf6iHNjnlh9xA7zcXAXaGINsfGFzL+zqJSyZ8/SRJB
DMS8UafVHm/VptS9mssCHNAkw5495+avqeQhV5Vsi1+80QyywCs0pfUAnbLIW8Ah/XRzhDvBtBc+
G7C8TuHZ9TzS/pvLinidle5e3WlvSv7Gy5dHj9+Ea2ni8/O6B3X+wma1fkuD1dG3lZjYeTbBI0CP
QCmHdlLGlwACLSk9aL+FRRQJG+SH2O4PKJJeRZuUEWUFFoRLQ+UUiU0tgTYKuEFnd7c99Y5tJ+zZ
/8oBhW3REEkw6kG4TzV9mWLKdNNHmTpauMnbTV+4KaTKgwXi4rC5Nto31VBekqiumKN3vLP1wLKR
iiJxWrPrK4t+jZUbZ1+Bz2FWYvNbeUUgCjLNP3m1SPnMWwwH0Qwkm8ZbLGQpXexcGeBkiBEnBTuJ
KlYbdO2ZHeD++V9FeQsQUgTLF3nDF1SkW4CgbM1vdB6Vbt63jeQR9l+fO+EZ7xQHLPDGbLMy9pU+
ecl2EbxWDkhpReqi0xGg304rlNRZUoOcZGBb2iSMIh2uZMxIntIiTcgs0pxdsoAYMPtZZfvA598M
UlxBK4Ky5Azu0P0dkYinSMiAud+kclmTqJ16tVq0lPew9K/bQEJJp7l5ieu8ulePx8QGPymm3Sgo
OId6lVr/fKIA1GJwwtWHpUE3CjqmMfh6No0gGih22G8ezgK8Tt3kQmXvam7U3x7919jrT3EqoKsQ
A6NfXtXu3ESLG945I0Ogz55oBqHcNVeeEm1ggmIxZju2cJRbyAnxrlnBDoCSJY6LdppA4rpW5V8h
lc+YukK4PwsHJNsEjYWwAbyxQ1lbgQdytZ2oM6w3rJNTmXAsTiFlqgSl08ZMgP2/NQ+j7YoYEEut
nsgi5bThKZIBJpPCmRrXVzp88YwakTjRo7Ewh93gB4Mo7BSB1fA5RelxhSXTI4iy0fGyT356tXII
B16XddBl0tbBQKmoEftci19Nt+yOtYLQXwuhOOrMVZkFL1h/q2r6rq/4A1LP18rSU736G5fW6Q8I
BfdOmEFg1a+mj+2gEDvfC0BiVMzIt8qGyIpXslexS5rq1TdjNcX1VBCEuQN6L0DqMoUgDrQ1VWK0
scsNSK7ZC03CGdJ2C2xcR5uYQCj2c2dauUJ+nEcpx/yOk7ofiYlY/b1N+M4pUeJmHd/9oKm6JkCn
v5gPD0Iv4SjMwRLVnNil+VailNmEun1UvGEk/vmNXVzJe3+gR/GR9nsuhC08h42yFwLSpSfuCatc
Dm6UPAFO0IKq4FlWCFebUfkNVQmoTMEMCoaeV6SdAyft/CCI6KmsrB/P+jqxVBwBxFP8zVLc4hpV
Rn0SOSesv+ThVZnwGbml+tAB7/uUrUaoEnsICa0ilermezXJwgGaEA66EKnH1A3aZ0O5yKVWUu4q
5uw021Oe1m3bgyLuYkVqbzEb73htwB8o6TpTlXS6iGs4lStmFzYcl8DNAWWP9lJyTHvLOr9mFidM
iB6b/J/ih2X6GQiQxWkZUx06V2lt+KbPtpZzUz5jngCd8p0h7Pn9W27d61/5/QMjgSmjY37VAYJQ
7suaoI+QyMp8KH1gkNxUYayVbttS+gpTODhlKzYxhsVX+QSfCiOH1cnG4fJrBz6F/W34xxaUXcDt
jUYedTT20Y5KCdbhzuULvP6uCk5kOqjRiLgyednvNWJ30f6x3/vQNQZPzfUTsQmRLfP7VzxIj+ju
RabBTXVs+gVK1J1Zn816/DE3FVnb2KYyRR4IhZ21PMcwn1mhOtrc2Rwn35lT2irywH+T2NCaXcxS
SRACe2YzfaiXuQAM+Yi53Qv7VfI8CmfLXXFuAhsa+W6VoZxRn3cnksKb+7MleWD6Xrb/n5tf+eqO
UilQbgRvVVmaebwItTbYBBb72wLifjduXIrkeUuZzFzR2o5/b/IbnWR5ImvYQDPInRObtzT1iWiO
2SroJGDi1SpwiuOa/jPqZTgSS6Zc2FaOYq/X7n+KgpURjIGxIMnhqUBeALNo4KTGOkml2bfJZW4/
HVqWzprX+HPpvLZN59AIv3xciOyjIBav8N4fzttyGbNWx39XVnJRROixl26Q5sdFcEGdkhAmud/H
nbpqs5njVszGOFqECaUdJtvcbj5aFYD/Y3K/0KHaxVX9Q/JlBdMQQM2chS+5zGAUQq1WObkZ9seb
BFiJT2x+e12UY1xcCe8Ycu/tYLed5F89P1IRZJLTF/lhXPa4rZJO2WzlRb0JD2RJkyVVGJy0BSXB
3m4UoOAGfc6uqkrJGlgLhyWYdVeeQacYyfdUkNPfPS609zCflMWu/QXItWzsAobOksvn9Ybjema6
neZQE2g+nTIIsers2HT5pIRDs999ieypv7oZhw1m3XCza9uGeHmopMMdhtgS3wu68V4mYIA2coMN
iiMvM+F6DE0o3013nfvrnfqScYXcviXGcE/UwzjlNnzheFe3NEmxtvl+ADss5zbQh3rl0OHp8VUN
wWp40UbU/4OlZlmZneDxBg+t41h3pWUQZcA9a7PCse1hG9AIx7Ky3VGOGetFqoaVYQjP4QhOy3Kn
eC+VjL6bmLIX7ZwyKvFfp1j+TTlgNyOigwcGxiY0PkQZkSnlpoEWz8VL4PpgxS9c3spOnBc+BOvL
Xgb/PLejwkxbVXjBMqkD0BYr2FYJ/dVkskim3vCIBhHLWGTKRDHPPb0VcHO7Ao2iKoMqUkXc+Owd
lkhW94lVCAuShh/3uJbvjCuxwT3s67sT/rAfN0gXc+7/GfSwEmVVN7NTdGDUqRzd1EjLeyb84NXK
gRPeX9nUbXQrbLMKUz9OIjFcoSRjh5YEzMJYSxsAwMeYtBuuffQuszqcQRphe2YgG81ZUc9zEVPU
/EkpjrJDQUnb14YA5NRFD+BAwMKbr/pKtu7AebkllFVxWjCeXXjaiR7uh7yrCibHvKY7uDEDpBrw
DcagQp48j8ztmYyT+9Md6Rd6P77Vpqvvm12Ou+I3Kl5CnePdF5KFLI0YZjOf6ntMfTN1wOXx4T2B
qCWU5IEaphmoyz4Ck7VTB2P8tdH5bgvN8C/Mx/zPvsb+LkSaWSxNqwYWh9Vs9Ziqnl1PryKIaAAb
KcPqfeyE8MvXsE2pyih4sL7pt3/gE9bs6camzxngGvFzpjELmBHAiNGRq6bsvvcleVxCGsAScvCO
Te41aqZGbogpLmDVjsDBio17CyThkDkp8fJfiYZXciqVshhMM2jY+BYnuZUAaUFH4J7N3tMAC8Kx
VOZm9TytSf7bxt5+z8WuNkzxhWCQJy/rMZ9aNjOkjasMdbgCe3QHA37bJT3l70WHQuebE+3b0boc
Vn3K+PAlTj3lD1MYn8dv6LvcPjNjTTh7szvDw+E1jWTXa8TrzVhMKrxexLIfQl3znNzVa1hj5ZsD
+knLHSdD9SW8U76Zc0q6CwjKjg1Lu/2p71Fn4sdC/nEJJac9OnoO8TFkX4HMFW8HxtZzwjvI0Is3
f+v+6G4A+3T4WYzxirp2hnkCp3aNjhR760ldDnWbE73E5iKgwpq+J96rx2jdPgo+ZNrvAxAtcB63
WNDnU54LJ2yRlhFpWCQhqafBtG47tqlo/xTmbLfQuJi2rEv1z3pUvw0fj/VtUqoHvl1B/f4EN4mp
4/274WlfQ7LYLbZy++yN61RjDF/Bwh8QVBBAuqhMSyTxobHrxclin4k3ejmMWeo8tUMSL5sY9N4s
jLpCqQ36SViQCSB5LVfC3wJ35LpsMCbYHGlyYK7dJJv8aVWXI0TOi4Ht0mtUkeodp3y+og2/HvQo
o/DXjf5K6LopP4GLuhC4uS9mvRG0gHva7qRe71b2IM1IgAFWJj6zezWQ8xa7Db6hP49ObMgwwr7+
wIqOtD9H12GykjhDzZlfa9X+OQQVcLF+nV/Nu4567uX2r0BY+5B/2fUkC3tNDlY5kzV60tNrGWCK
jVmgTuXfOee3cjeHTRGTmwPwKtIFVm0C605UQSVU0s/taqSEi2Kh6czZd4BtUVx7JJexG3k0Yv7/
+cvYJUkBbBp2lsw8v11+GLz5LIedw/8k3qEBSp1aE2IS/GEgewt+JzmJvQYbSuLgEUy1XsIUw/K8
IhpJ9Xa0vGtsAfif3FQFfCTtNIWXsEFyiIKeNbQitIGgpXJYj1jNl2MKWgGxTNIPjdw4VBkz2Gg1
wg2b8pqXW+6CHMVfyOESfzYOlvHjkwQH0dfbypasKSbbdEicKeZo3VjoDAaoXBLknVsoD5ex+yJf
AUVB32MAA6neuWfGoTC9XaQVvRwwFSxO6Krx3ePMkRvu7r2DyLJJPEDTW3N8xktckIxuLxA6FIhs
WJKOtox8mAeYRSsVaabCADXgRsOvm4c4o5rWM/Cqh+myAAWOQ4H3Vs8KXHrTcI4z4LbCpfn0MM9U
UL0eq5wW7Ktx25nCWx7J/WxJctiw+Af08tVoGt0x7yKb1Mpn5JzIAy/esRCPCTb3crruoOZZFAPv
pfssY8CR5AOEg0HkM7OQjoGKMgU7Badn3V1ILTemvJnsvON7evT8uUMJpOoXxv61U/h1v2eOLVRH
AwTi+Y7Djg+R6KblaIaWmc9Vj0LPIT/rmouig8yu9LI5UeiVIZLkQnttNE0ri2pxK1MGq/BKwXwR
5kS8XUMwviuQMyDE1vaO2kYFk70RmM03onTYD4+RlCSmroOyeXT+fxRiEsF4ui+quBb9f3omOVAa
djbtrTWAzUnji00/Rd+UtH9fyv6syTlSzVsGBavU7pZxxZ5uk+2aUYP8dhj/eH7OY5q9ucboVt2o
eSrVHn9OMNVr9UiU2E1ahwsgMu/zmBsNf2RGiuolYIip7ZtiPweVJg1CYgrLfcRJe2a89jcSUQpy
lg3aeqjw8az7b6Z4RfYpP3Z6K7uD4mz+bD+FsW4ItV71jsO+itPtrYCMJ2gkB8tuGnMreJPdyBVz
F9R6rqVqpu9shY8oXzgaRomfqsO6+yqeE5ymLL04BGDb1do08ss5Kb25U4faMM4R99ot1X2vHvPf
yqFCvlx7U/is7x05/vZ8F/fMG99m9GCjbS38dPmcYDkHXzf2XmpjwG1EW41kLiTxKDnie2fSDt4q
I5R6glokWIqwEXYg1R7MesR1LJW+CKIEXjLZUDA6sNb3Sxjbw6TTGJ5xI+fXMLz2T1FJhuf/jf5o
N5maaoiFRt3Jc2f4tx/lOyfsSTYBJiNerC5DnBOvgV7O0mA/TVVgGVpxscAvz/mMRARqVXT19v4a
pSfEejLR41R1rKFY3rjjJVKRp3EEyGOp9TwAAF+k4cmbFuTaE4CKvhlR5cEDfojnfB/MX+QzbXWS
0D1Dc1MTal8uvWKI9JyGV2cJrwwwi4q79FrofxR+l3HeYvXJwQtLUb1WlHIVJ5RWn5UD74tUBFTK
O34fRVS1dysEELhVNElMDvC4GkVENVKwuKvtB9Tn1Qtl468nN+wt4rUjvOMJwidUIV8hb/UfxzDl
S3YL0X7aqBtvntzym2vB7pzCnOLr2ejaLsCOMW4dpyd2Fbedm9s/7NhRiqPShmKYE4S8xaWxXDyq
5xB1hFEAW5s4/Xrryo7kMMnKVQwJ6NKnHOONGQI2uuD+DFgyNeHP9Ddle3eSWfyAsZIPGbLV+C6x
xxewOeDBB/9f5dd26plNlgCsoHLi3KAT2qmThR7v1NevfYtbPw25QgRto5rK0yD2vItmKb6KBc5N
TBH/eutZl8VyxPGapxVJIMlYNiWwweRvXVLyaFbUC0go6x1YwW79NBdbGC/BrRCBARhbEeIEelcQ
FbXS2RkG+8i6381P4P8iXC/5TZqgRJgyvvGymPp939f+YktZh/ooj6TPo6Odz9VrmH/d9D6fyMhT
Kl5blaRSwPXQxO8eT0X1DnYc127BSB+o4GrJjwt3fS5a+xHPAGYPNr077X1+/7atSNPmFDjhelxY
W5S0GhmJCiDXhL7FfjCMj224QynAVP8U1c1DMzrJ+WmycBs++FNg9bv4tWUKIy/79D2UXkywaoxV
TYn4Uha8k/Py86+qABP9EQQRqejyWfvyMkFeHkB5vwSDilLBR/T/k6srE+X6PfQikh4LLfzM7jZP
LnsfKiXjDcmr8jDhP/2LucnOe8zzWbnUgw9oN8FuWhEgClgcI5vdqmAZ0pIcWaNoZzi/6AF82PBm
du/ye+kjYImluxZhx7ZumYhpxJewThptvCSUr7B0QD0djof7IkdkjYNH4cH/G0ZkirrGLUjssi7k
96xHMneHBBjT84swxFSlmtvgZNMPKTz+MTzAK7XvZ6dshzatJOVrGXTQDhYTudrbuYhxRHS5N1Pj
3LBwUo073+7rWbFctZWnSzWMGUJ1lwikJZFYePfGM6RjMQ3XUGkOA4YhYn/J3RUwcGqVEFdFLw0E
teJgXtG7ml3IdqFq32ZVSzGbjOzA5uFHL+/BxmoP4SBDzKNtpqqZpnRkFaYp0sKqwEmJDIfJkQLV
VEQ52rpOFVZoFKBFCZZxb+Rf87CmKHnRxN9eCJxfeADQ6T2i2VCjDOEWEU7R03W0towP1T40C/RJ
l9rlTMn6/2l4rD6My5vauw2YX7VOqZuMX6I+oGwOEDJEfckcgoRbWcSqyI0A1PcE3mYM4yzIgHVr
tIlZROxKg2wAiJh1n2+COh/URbwwo1YmRm/NrldD+IlhW/Gfy1FjrL8cUyF+tk+p6cipcccJsgNi
xhMtlrFGj7FB55DyBSKInhRlEJiGd1XZGHf3WblfM5z7LmB3AU5xzw67UJr+q+yPb2EaqLhcIQDJ
+D3siFN6lZrFBAQ6pASyjwTFMW9rmhXE5ilqXjJPAh0iusmog6rjMV5mr12tXXHKyTtnuuocM2qh
v+Q1rxzp4jpxaf6LDyux796E/9oxyS7YrZIxGXJ2hB7IBJKPmzzQsMw6qw1Owki0yI0/BJB9ofDm
jFRHWItEPZX3ml2LjaqxigVJOw2UC0i+tw6hJyXu25YEzN613fj9Sh/DtSQoj2+CbY6U4JXc8Uxk
ET2gJED86QQBK7g3B5FofyfV7u9gywmfa3pZmekmGO4cwpsLmytKEOI88+ZwhTaVckrbI0naMfto
Xl4P9BJt5Di7T8lz9c0cofqDYE5wiC7ddRy1h5TF3Pk7ZRB7oRGyQIp+aQPHPDvVHg31vCUAXwkW
Nh5GaE6fNA4n+V29oQ1/6aQ0e/M1amzuBkiLF8HXnXifGo70xZlHXYFecK6z3jpqG+S8imqkwYQW
WyAMm4whR8RV8rbGFceS9B59GfW7fzAXBv9cPgJarm45ABYMkd4G3nuzVzDsSInvefrVJrhPNZfs
Lvnk9OAR3pLn+mQBQxm0tE87/3PchFCHtqEF2hNxGpNHJY+6U3dzfc6tQQaYbHS5WlG+WoulMB8g
EVMdvEUOCDFaJGCoUtpftM7UQOeUXiMEJ/BelNa5q6K2NvwWZJKWMxGqhRdMTTIt8SvObD3MhWoH
HXxHury/eoaTFmEQinMYXWRl7yRP+tG34kHhGTG10dBL1nhXqbbT4guqDiatO0SCxZ8tvwx1Y14j
qWP5ft0ohruJ3RMBmFki+t2l7VzbKV71o2lmO5VxuQXgj+HFC5S6+5UqD7VokS7quoEv/lpIJV83
yLb/kyLrdXVW7HIuivYQ1jZZSuvkEgiXfAPH2Gu7T7hHsQvVMcHz75C3f+Z9su066oMS0e0OwC7+
07Ts7pAY3IKWb0gXACFRD9zk0zRGQS9RVo9eGGzeG0/JlkmEG0BT7FBTSq4EygAAI4DT6YK1TDj/
q11qOUU+JSLJ+i9qBCPsmvNpxog1mG0MJoUmlsfmMAnkPnf6X+WbZPu6zPr2HCLXayhg/qsEd8OF
dAaXSBMULPNIVMLkEJq6SHJcYifx9M683EPRTvXG5CV9koM/SpJGpnbQV0Lib7UPfeh+YmjkIpNK
UfxuqZWSNtPOnrWc8Mr3Ck7BPnSUnT9SAdYDzqDMWe+0Cqo+FYbLPTgBnBrM8K0Y3GM7Rw+pSXNp
qjcp2cclSED/6NzLFf59lSdwLR7quNzIApLxRr6mnkuWhndgTew3VfmQR8LAmU/t0cenNociXzR9
aEVCWco/maEJcdlI2GShDKZEX1c53o/Ca+XNab5eUT8YevQA/uAFl3fMv6fN0Ay2/eLUHI979ye/
FwHPgjYsg7AnXedZKFAigZWhenVP6dwuu2s+eOFjzEIrm1XBiTFurLiN0Mu8K6EAymG73SgHZ9ne
46baqClp+NsK2dNS2+xCpLLHjw+EuPfATchYipmByQAcNJ7kAKo2u8mZCJEEu3wH0B24i2qssQwx
zNluU1YrP5wCWZ9oTiP5YPaqm8/OKzrkkVNPJ3z6zVewj/t4HiXZ65LrAMi4Z21kVlJ+zyz+xwnV
XsNS3KCXdaoU9l6lOMHR8J8/fiJ88RS32p0nJkd2NBrba64iPfCTtlswESuROVlVJnSDfGtWfWhj
Of4eQnJsCVUOdFciMKwzMuduM6CmOgGumWTYUbwaDiHD7BFVHATVMKIc51TyqGOLvgv+jVxybnMK
gMZS9BSB4ZPM/spvL7Cq0oDsgP4aYFGLSnWUNy9d7SaeGUAKLkGgLPL2tOD9rZEHN1n4lZsF6aAs
n0TC53e5yrTQis+gcx/OYkKjqz5RR9uL+/1ne4+lWO6bglE6uEnV3QBsQ/LD29Yv7xtMXWNZXBPf
CAlMKJ+gw2Ylpg7jm6mVkJ3WyZa7Dtpnp3lP+Iae4Yvm1PkhPvm/Dh7ICnYl5B9vDrEnIH9KItQg
2hi4+YFRlgupFeVfb7EBS/xvd3hNnNjonygPvvKO0UOMyJyq+FkNXQkXA6tBohOF3MWFbnTmj+P9
LiwoPSorLrnM7iLQRSaM1dKD+PTTgUBDRSyqyxrgvWLZD21dy1kPBQFZ+28MukmD284AjZMwL6Zh
YNMakLSgR2DN6LgQ3iyqlZjBF91HtopCpigv9SWE5FDx2G1W6hmGhRZKzBJ+zhKXl6P+9/DBNDpt
C2lvVYp1Pnof/yQpD8fjLN4bXCtRgfYzonh7Wy8TO2yH3D4cfdSbe2EBrY/8KfKyvjKT8RDn9yTh
ccypHgf99YZAuez2RDl03A64hv5emyiXMUzhTkJQXIE65EgiDFG+Ii44O1GiJmjtGwm2oUMkQzRC
NvkVBXTXXEOmPf24EUDN6GgQ2wxADnfWouykf6N4CCNKdzRr14iS1Qx81hgIl8CLDu5s1HytLZVY
Gbty5V4iLzZF8k38OsXF69DlGCYacQGFzj5+66B8TnPoqhU88jKJc7C0bAVbLt7iSE+4NWDxxQA6
51UhTwGJkvRiOU4jC+X5N9eQXYYd774VjlNPPnb0He5mYiWGf2KV1sTKIrONdJ7UM5EuD8GbEOS0
V5ROA9Pp/Gbd2iIqUwMku866KeeeJEZXj50m8DQFzn9/7ApQOPvvayzCoW/wNQLeAJXLlr0IrqBu
0JtDBzMkqwxKxux8YA97zTxmV4Ftf1btj4ugRmjehPb8kWaIumus3N6+YxFhX/tHQEhtTMk62use
tI+KLxnhZ0xA2v5k2oYcqFkx3HdhXeGgo+7Izp4cvDEOzncmeQB12sYAp1bXJxUHQjzyOjzLlryn
omKEE350THMbiicGpq66N/uyQjKnsjq19FR6hVm8Aze73b/8EaA12Gk016nuNZnwHp9zgiV2e2z7
P8JqNe4HF2abBuPrxFfZIsrDhBzoGdjC53BUPoVyXbDofC21EHVYMdo1b0GsxgxcEdKKwx2Hhq+g
aaeEdoOL9WraXjQjK7lNzb+cxjdIrycATYLqFdx61AOA2wOmrQukVV5wJZXWfM7HF24hUcrYPwky
hEMldMloIF86maxY/Q0JInPTRPP2DQDz4jMGCHWnraDlGFJS0WKK9utmiM3S+DA0q826efYnx3z6
lHlLILMMZrN2JODTR0esJ6eVWchsB1Bk1MH4au190jsbQpemHIhe19vN3h40NrtqTBKAhouTM9AL
KdpeOYcFxjX8Acjb2XzameZHQDloss0H0LSvWIc/v5E75SCyFiDUyj9xd+NViu54phrO36sso+wB
wxWNzFN1ODiJCoURGUVvdo7TJwNhrSsl7W0EBQFUlZtmxgVaoihs8Uyiy2vOaY8MGdjekAePTbIV
7V/5d3lCESIT3xdRZJly95+y28tzYEcec33AqZqDw6pem4DHXYt6NT1KI80JjrOZLTKYI3I5lLDu
mERhpx0h4rp4WgqDjYeewzbdQcFayyl9YVuILMFDXWW+WDHBam6aDGHWDmTu7AaC6Cxzn6dnky68
bz+KqWODPO8I9OE/L66QDJoSwE/IHgAgaaQdzUKZj3vyGF/7pXgn5CiFroqd/G6FZSrg4pERaPQI
AT8qD6Tah9oF3l/x9KUGBrIONeZdIYlNwLLZ3wUnhZP6oZ5obv/kK08fjsE4PTWqVqfL+BC0/4od
/nVwmTFwWtdQLEtIkggeetjSZ2MgSSQAvwdtsOnA0hgnLSsD7UTndWGOiyy72Gv11c97B8WvEBr8
zT93lN28nazcdCze67vfbKJMGwFpguFqHHQSL0aQmgplYI7PlIPxq+TREw/pgfmtWQFW547QXrGl
G+EzFnRejJJ7GNff2N8ghRFNDRj0wkDrQG0vC/bt1BGacvgx4DaAgIqOhWaO8fFcWR+Ip5fUOoKE
wB0vQk2aGQ2tqbKM+U48SGVGHgy2zd+3XzY7xA/7g27LHpW9QDoXiOdKo3nb2uLhZBgmRAocp8O3
0d5D3JcI0noDrukHxfhIahdjH5QTK7zKhBjN/KyTvKeB/5sajIyzzJIIP87Y6Kh8SjUehXI374c3
YG0Xp7Li19yq7VYnbqG0TpynY3ixT4vWchawzVaiVFaZS6NMSgunxndXdRhgNC7X3Nxr6aL6eN4g
GA5Lh2EPW0DJV85FFjuCu2H6AlbaanjEdWo49acBrw5A0MQr3tkSOVy/cIPp4K8G2cYE5kvm5V/4
uQyBrdags67T4oXR7TvwRqKTS1FK5750t5DoLufrVJhM86C1Wats4CfZTfpzpjBXnH6dFHLUdbiu
zBgfCr7C85TKjnPRSzIT2t2EZOWj3TKILd4b43MN/pmzG1lwPz26b/4xH6vi6KHf4/MwFf1uHv9t
LYdJh7YN2G0QmPq9o3iumRsSW5M8GJzdghmtQHEKZ43d7Fd3I+6+la8srbxhtOr5KI5c85BvYs2x
5TIwAQopD2P8u401BLaiEiUf6SkR8oGisISQW9WC6FH/OlCE2i769NWscO5GmDen+5bexgdhdu6I
F+94DbVIiPZ8NU6YluEnoc+czdLJQUR+lwan1YYZn2l9HOgcuFu6i8RMYhsD2tpqAjyZPmIZQRMG
vspHDcl0M0R0F5OSg0ggesrzqKnROfMh0+V6BteRl9MczQG6Z4FC1K5mdGMiZ8VElcHqs1HZFW9p
G0OAEmcJ3HVlqO4GQuTyFdyoZF9/G/1AQHeswmk6cReYgBkz+VHRKbS/70bA2iJAfFUtDywaPdyp
a9EWy5eWVbFghRxosYPxepnd9DtCryCwwyXIHD3JeODGm7yYVAHa5DbuGTYHLygIsf//UbbQb9i2
JRPDzEvkDElRmNwEWzEjDv6jwRlpR9WUarIjWU5lE1n5t8AAaWii+4hljODRlVpukNeFkX/5eJPl
ZQhTFwIULDzeQ7KuHSiU36VDMOnmRUVU7icM+p35gJQ6U74dwVmc4UA8rs3HCDHC8HUX9QTuCskg
e6Z0shgpzAc3LK+6aYNamA0aBRKrWtedgmj9Ji43pS/UbisvmDrNcxE/HXYcETqFUOiaZhkpyjka
wpyTRI6Xz1UjmtyDQdhs+HDGAS5SlWLzFGxCMSW6EE6Y8lvkIGBBxxsaeYT0PClCldS5v/0nClvl
TWbxcNNvnvJWdM0R6RPfjEYjfcJGBd6PaSVF5T4qCVgbXg9pa0pSoPWWc5cLDlK6EMYmjG+rQYFq
bWP4aLB0OxC2AGKrT4BuLNtPtBq+DPTujuQFf1D/0AHSKm1X/Bg+pIuoeRs2S64ko/OBxqUA9mHA
gEzSS9nGrhWG227ga4zmhHRranaUq5F5YrKp9bS+NoKVVScjOgqYVvQ49lqCvlAw5LTjSmLkyFSQ
EykQ5P5o9BSsYr1yzOjRtthTTwpeatNc5MYo29axvP3TDyLIPfJ7/OxXW7cQ3YE+yR5vXFV/ZyeN
ewul4p+QfMuvMmHX7bqnIbyh/AT9FxQoASOr+TjHxLQDUzqAk1g6mcIeXlSq1h2hcG3DWmDwdI5G
Rs6HXojXolPhLK1ryHxrQuQZG+NV6JqiArp9dW8nwkk2Oims7z3N1rWoqBQm0BvIEezM4ZMRTSok
dKkwPUHmWFbRwseghJ5j6vJEffDtnCpyNaMyL3UFz2Fh21DByX1RApdaN4UEDhAtY2PXiAkdhoV9
qhUiwZxVrdXAcU5AysjwNNASDKcNkTU+tXNwIxnoV893P/NHXfMkmjPRqYgXDlqNM28zdCgHv01P
i7SLf/um5zU3Z/nTrgq6jWLw2Q6s1BLCvGaBxF2cW9RZAVj0i0kL5XSqtv5bC4zmc/3cBJuqqway
S3SgQhUEx21/cXzQeUCZcDa93dvIJVwdEdVa8pynX+a4Oh699PJIcVJOPFWGrE0DajPWIKD0n37e
H0VFjUqif/FHRivtcd50wbk88U4qodBqcP6VzohqmorFaPYtAzgAu3ramY/kOEBniDG+jckFcDYb
eW5mlzft0tbzgoUaG2Wj+vv9fEMy8hXPBpCSi001EeUrFpPt+XNaIQVrhoiqWHu8MQDzWYTcJ2wJ
jviifqG++QjMpJsxlRznsiBAM7P9Hh02e1R4bSqvTImeGLVnEq83sdEaSEvl3cQw8uZt+9JHSrd5
Uc6u8guIT8NvewgKsjQCULnJMnd9vO100dnulEn36ukPCftBsCmcf7ko3Q/bS/v0QsXJGjo8wGQn
klzG2SRj2dNcXm5/ayvq7zYaUXbtJ70fmOwuJuQfWq/HXRCYdIh8sObxPv/vNXNAn8dwGh4GUXGr
4RacWx/VmdvvAVNHv7m802qyNR8AOepelJW5VDT7ocwm/8nHEQMeSnlxjLQLHbCHDkkMmtn6fdbB
ocEuh68dH6NW+QVmx3010Gup45BKu2cux++3jv319esyEuk3DoF9DZhGPV8dn/npA4adXqlye2gr
9M/yww6GH2PwXDDxOMG1Gre9+IGQMvkP0FuQ71PcXjdNAH5i2A9Hd8zZ9rdy0Ft6dW/TCMqOE4xH
VwykV8FwciulVycaM1NLft5bb66Anbvqqs4Htokqbl2laNahe5NFQXn6gcgFR2NXc2YgqIc4DXq/
wR+7TdLOmeW5twNOu2PWa8pxtRoaGVBr4+XFpvWOMWKr+FCEBXH7jvKOOqkXgiqWT4uM7kHnZ62E
jM1wzpTxvx1c7NA21ka+9g7c1jWuS3r394HH5PdgNhXkTMaQ0OYjR+CqUE3aeMdVKpv9gwI+bVn4
b+5Gefxb7bgh/5Plr0Jyqoj63da2Gtkjt6fL6fQkVDkdd/+7p/omlHYJTyVihIkZjrUeyvjvZpa5
4P6/7ZY7a5hdjbO3C1tFfsZwLr18Giq36htI7CE1siMJF2g/usvYhWt7so36iQyZk0I8ndSTsPXz
HhS1degq+J3nTaoRCOBxz2DvqT276Fy/bfzUC6TEJiTzHfDxfMd+vS/t9qLqiNubez3ubwG9Q6bw
P/0Xd3TRMbykZweeVKwPEldSAB03Vrcbm1KznJGFnLqVyP+des155gaUT9XSmEDYb+g5DrsVTQSd
jzRU4yYxemPe7wOfA5u7VHW1nFuGUTfPg3iD/YWvVZDObpIsCe+rMFDxH34xPAyK1lbBTZPZpbXA
k1FLnvXc6ix7o8BMGMa/jrIj8XXUk87MsMX4W+j8vNiy0XIoBJ/blJdIDNCBEiJPKaTEuNS7Aruu
MNsLzT5Ubj1z5DPB78JYeOyfrlDXql+M/X3Xk/wLpXWdMmqTJeJLIFtT0Fv4vvIqSh9SQsRGK3TP
/OO328AFERmwpUjqqY98HUMnAQFBEJnwGtJY9j+oPLJNqZLCaaRsk3kQiy9ApOeLlKVHmK0hxvTa
MABCf2IjkgQko2AdLiV/BBKK2J5ccpe+nyuyBX8i88oxQmhOKF9ocD3r0stM44q+4q7rt02xxbLZ
FVwJktXbXG6i67QQpykmOxJesaZGTJWwwKUefc1E/S346BwvGyZnP44rPPf6T8yx+Rg+PoC6xHM4
inGM32gCGKSvJUMHO5pcsHt3TcvZEgbSKuMeG6Qv7dSIrRNJRdjYqPkUi7JChusEvkTQR2U/uSLt
5lckq+MjJ1XIzEgN/rb91oIy1hh9U0FdI4YhiWO9CH8lbRzqQORl0QRhIRylid9/gWiN0pZDlOlq
QCPV+gOUJL68iIk2F9UOvnTdAMAsJ5pYRsg5Ee+6YPayIRCN34OfRt7HOdxkMwbtmo3NyUbLzswz
ejdkyQ8b++0aTg7+W9UqXIfmVmJbGRRfrpL1+4ICK9ROZiUhZ1WwnWBwZNuw/Ulet1rGASbmyMu1
6iN6FH+MFvA8dZvcggbuWtYwnlwLHX7uxqRsTXQzQ+ztu7A2OjLTyOXptm4JYGfT0Faw5tamh25z
3sy5KiIda4aUlJh/SJmT16e9fuhDrdt0PSzsM7f/wIQOmChUMaz2LDJTsOeb5d7ITTc7DMfR2Mv+
E9CwMh63uSRqnfoLQysbqm23DxMFI+pdX5VD9TruF9SAEh+hRigC1dO2plimXBWUoO8iaE7XAqGb
zsMgfGfY7j3uBOe5R/F1mLOl32Z+IWV0jvsjQy9rBfOQJOZXS7GFzfqw2LE4twkkl+JjL+lgCXqt
JZwJmYscpOW1iIaw8jt3dNrfQyBTMdavk7YWGFTXUPC/miTm7XkpxtOoDcMmQx1b9ccJKIR2BNi0
tIqAFFhE+0H7C1KHTqf0zV2ASB6Y75+MX9jwYT1bUYqg2Xdse/O4IN6H5h1/BHJYHMXySpvFVrbm
yFkiJcMrJeccl59KsPA+MCj6WOBZsDcuX5W4C/SpZGYOBwtIqWXhAGm6vmBrKD/tySionq8oRCQ1
9FL1wOLCqyMWgzGxI19fVUUsCYrHjWYLn7zvSo3cZqno1/aEnmUahzAwUw04fhQ5JrpdavVkd27X
mIUMUl6wvr9oJUJL3bHMgfVcN5aNzg5dCU6fX1ERHUWwXIfj6e7PlLtcRJnVkdjEtQP4ZHdQZcdn
/q1VFduR8qgYbHT3KA0MpUIFo9NiKNHtj9Wn1Nyx6/imwl83WsfSBT4AhScuroMZjV2MpP67yTEi
K7SJbqSm1JffFQ2WEMwJPKwjUU9eAO6BGuEbTpkJWyWjX5U7pDWVXwousdf5JSQHp/Yi3KNa6Yb6
U01xu631LXHDCT+ndJCCFkwrevP+hN4gTBv45opO/r9TKiKggjTcl9v98mIwGSTqoGy3NWMSnRr0
Jn3TfJtC0eZJZ3KQDK4J9OvCPkkmNo7uFmBcjcB8OlczknmQPeFFvDT9auKPrv5mAXXOWOt/m88Q
+7iK4u5JZWKC5bzPwBCU2kMuFkaEbunNHKsNjydCS1WUF20ekbPmvdMqG1WOZ71lFGKQt2jnjpIw
hHBHyZVEleblpCNFmE9aTq9pROFKr6aKre17FVBW2huq/D0nK8NHCNYC2eTXmGs3MLsNUs7q5nSL
F/MWO3WF25M/A2QN+INmEkPb/2EN2WJgze9FueDZ+iJ6ss+leqKgxvTxJnSsmyH3MGbm517picW/
oU+Yn8A8xqUiueoAERvWk+NmOJ9O4hTI0LacR2Xj5M7SRxBhgVAe8gAgHuDTnv2PAlI90fYLfiUE
R6f/wETjjLQ+qtAi/kXmPcT9AqYnw26bu60yM1KINUFCapuFbmAsyU9ootl2zaNDQ0hFpZpbQPL7
SyGmYPsdlPY5ImWwIk9EsjZu6lgHDGrUqmh+hzD06Zp8gShpxDMeGPflLwqrL0VafojajX68VN0b
t+XWB+AQsclsBa63kq5JrjyAxWOL0Dsph6LifNUI5nvimiV0i4SfIFMhpT032LObACPatnOq+WoD
CJgNZHSD5UcP5QkjhzkR/hk/URVWHd3PRsnTpdJde/lKQilrdnp2Qr717mPVDg4ECELzUobmtk5L
h8+SWO9fRbGkHLkpqRUtUKZSbbvB6N7CWXV/iY/UElV+Bt0ebuBYGJLaVfZ2JHD5hd5DxkH7CI0b
yeLyop82RfjDr4QuhaN4UlwL2pmxrG0P7b6ly0JLMZkrNiZvm9lUjkK3SQLHZDca2NV/RGSdu1JI
4utuZrjGX/7EbcUMPBXVDGOEghITZscQMQrIuMsoNf7V6mSZzubBD18fyodpxy0tAmOO6CO39Kyn
eMuIl1Ew1+lmrb57hosqfVBYFlGOzHgybKQOEZXZqS/Ik7YxbpCzwKaQWOHLy2NfTBVQXHLhqQnA
DzPd6efSOluLJOO+7Mxphj6Nm7I6JhFEuMlRvf5Qg1AHMdEtOarQBiiD5aOaRbpcc+QwJdr8wWpB
xkw9nifpFdENiHUK0reFxBZMbx0pq5bDQ1olDTofN28wq1gRen7SFvI563KwMML2LdDhhxK438h5
ZEkquLfByJDpcwj/A5aQ4elXRHS1zBKgep8V4dVzREp4z265Ffn3+/DdsfOPBVOuEqOaR7rkptwy
UQo2cwq1ZPIkhe5H+e0P2t+1G43TYojRwMqQo2Sph0T65L1UoZ0eNJKQAZEfQOmSKStF8JfP3tV0
CS8n87oH2qieOIibTFPgq7zSKWjYLy4EJdmnAlT5h6JAphF+epi/h845PNzOrsucCsx6tpgo/h+d
ASsYnvPnXJhwhzIc2YJNP2nr2o7L/8Eb51jOUfJTbWlM27WHeXQVyutzUH1ZMUC1PcPsN2CkrBtE
RZzyYpOScXv75qY+Q7mAMRvP4IKf+wjim+SqUnEYJofJqkB1O6nmM/EzDIZDa+ccmzjiXnyzrN5Q
yZ8gc5sIPtS3Yw1AxsRWCuNCB2x8ZhHXNDuMgrsnOaqTtfbUBcYmGV7Kfutg/xQ1NUDf9oMujpCh
Gk5Iqtn0rnXYcAd4mIPmJpF5H6rs9ujGdbXsTu8fdzCC/9gOqZ4Yp0f8rjQSiW1DbY3WagGlwmhr
rIyIx9qNlgKhO23pD+0HwBPUe32Vv6gFCxbl07lcBT6stVRY6ip8Lkuc9xFXfQCy4mpECPMKTRI6
a54efXdeS49NwnkYdfA4r3mIy7KMzOnIAYptnFPQIA1sFZx7rvLPUhut461FMjCAHDTG36GnpbLg
B6UwZckufsqC0YBj+d3IfcAuU6ZNmE85YbGnnprlZKhETpqSAnyC4HIHkhykIhh6BGv/pa5iqB/S
UVyd5zBabu6fETLzV/ViUkHt5EKx07XLWV5Ir9OysEI6touSkUP6Fc7eez3RN2U8rh/CpbWlXZJO
Ys/IbCpWL30JdfxWGXhVam+9UZFPLwnfOedtQFIyLHp+/Xc1sfCPQnk8INraRzZUFSc1HI16WmgK
d1iQehUQIlBcPvO6Y0nZ5dkl4uacLVMUSfT9Np6w9XzgyL090kURnyOsPFELmjOMsw5PBR1Td85k
1Qq5pbLrwr61cG+vNK5RTPSbX6INL3ZUfF+mxZ98sNJU/0MbhY4yZhj2ckutNx6xrbEhZDKzeohd
ocyE8PJ7sTI9PcskLn9Zgxe0ETfDNrZu5mNwIUSFTNCswnkpC94tcKsFoAUUfsw472WYnV1xaAqx
y1GKGtKkSmAuQcEsaSgE7+zyxdoakZLZXJ0+ZgxGs5QsM8J8+Sy3XC8v0qw1d/FjWbfWJAIoK/cj
Rflq2SlxaRRGJxqW5235oBI0oCfTFGHs7SVW+ewLBtDOTbOzEJN19faMEx+fOwu2PwPlYGnm3mnS
qJDqxVfzCt7i9puqT15+Vk3IRR4GhaMP/Qu5BtJj7TOKm5GJAhVTmDGvzeJnYM2kpAgTLc1ZKuFr
t8EokTlxs+mEyAvWLB4nCp3SH2Kr1HB3vpBVPVIg4aCqQTjB8VNVbyX3sQtqLoSphs5nS0n2xD5Y
SAspsTVQ+KHBW9jMQudryUbc0btVM2jd6sz4Uwm2WnFGlWYHUWoLD4V2BAI+Hu0wEs2JRb7VjWc9
KwuvHjjvm4CGBblVntg63a4gL7e4q0HF+8spX3E/Xy76AKal9hTLIBfRWgV1XhpvY60GLpwOyCYp
voxzfuV4BqZUsC4RLkulsT1U6F4ylmTBS+VzcNv1qdnYH26hrrZeWIVESQOzXKQoxARhj0auNCgq
MIxr2r52eGMMpFP8wQIXXEn8wRPm5jkZ9FXUyii1wcMirWQMOJZyabmgWkuFqIZIyi6++wckHByG
2ZueIwIPBTnUkhz5t+Nk7yGbPs89qqRKFXUT/arr2LhiL0H1MxCKA/0VIFX6GmWpeE3pMgk59hp2
k8qgQshhaeLDGzX5Qf84VkinVRQgACQLUW1WtYrH+oYEA9W40rQnZ5+Ocb5Gmrlbn67SBR4Y5eDb
0h6QQ/1rjqxTrapdUn85PZ+7fXHYmJTyCKizNVus9xkAuIx5OMbszB0BmFrrj6rSd5Kq7tqABdk8
Gk9j4YwFJ47YlwnOYiiXaYdIlM2jwfhVCsl733ktMIPOdx/+935+sZJ1s2m6Cbzci2LCe4PhfOij
oqSEkN8k0QwcUEcYDo1S7imD1D7+gwZ/TtDRbKrQ1PjtEUEnOoJ7aascROLJ+ODsxYbDe/EGcaa8
ISuLoJ4w7TbSwg5MIRyaPw3cmQd0e6ajKVWsHewVDKzdSWYNzIzU2RMvSSk7690FDQjMHBQ1QhEm
M/yf2X9HdENagFnSyFHMHkOY2Q5F3o5Ehklky0TYf615zwtEu1zOHAGW0f+ztuUzk66ehz4Lfk0q
Oz5bwYfErjgNtqbAjR9Kj3d8DdKXyYqzoDHYE0aUJsExnKEqGz9xwDh2xpk0E4rRwthwVogTQSV5
v1mIDHFDTBNyeePOiyuiOSAWht9aZFGkmBIkGwDPqsSd/A/PwJjN2t4oTfIlkfF+N32r/zkSZVr7
6yRrjCdbjtuJ6ZiVrbJCxCKHbsdvSNeAUEEb2Hcn2BGxjk3Yn22s2t0bO3uBCVNduq3eovc0hi7m
aJGYneOlo3NI5uBMSqPYZgMrWyj20Cs70ckkc05j8ks62kaEAWm1OanjPRvKuHZMznal673Qonot
ftJkYaWf8AWj+3YvYX8sjY5N4ASjALfk28Bwt38roDG4vhMLAaWTP0IOF3ngN+6Ob204ULOPchOr
LoWPhsO3u0n/veaj6EBFNEjw2ifnlFMEdNWiIEnPSmTHC1p0mlSMSuNQ7WZqkDsUuimQIBYgrWio
iT/1zx6NuAruRssJ8PmuhfXJNsFnuCDJPXQ51ukwpWgiJcioaYIVWuvtlBu2KcOppte6lBk3lThe
Wr6238J2lzF6ebXuAKh8NhN/VWqsCFP08ZfeIhl6z1xnMQ02ZPbMNm+dpKNJbX1Me6DvjK0m21M7
RoPba/wvuAKJGlZlD5MBah/SiJwOhksm7QhS5twsSu2qEKuX8t2rX3jQDbFY1Dv2OPIuxXlqnho/
86EfTdOEMZQVl4nHwnkHACB533Q36S6oztyTBkPBjGDt/Oa4hz+88Veex/UCCnwiVfKzdab8z11Y
xqZzyfKQ6ezOAM17HRux9Za2yM9isPXX7yFETDon6YHXBqd8fiQNSukno+XyFE+dzqzcQRMFwhQ6
ypRS7x4/nRT/24j/W/ClsBG4KvPySCnYpx2MBNhkSai7nh/1Y4V2dT+mbyifwNhu9J0bAqIrSsXY
Uuy0UIoiIqx+bGGC0+9FF4I96epdl5zdVfPJflwiWy657CKkNBei+k5u+dAsGALxn2Imdm396pyR
hxPxlEcNPXdz/yff+rG7z0qlPQ3Cx3ywSFsP3FRzFoG7ndeCLjMGICCD4tc1aCk2y3MVYEvMacVi
2KLJa9v/E/fkxd4BgkhIBVKyCTBf9aUcq2cbvGV10+KlQ80k2/jOOgVN39zr691SheYPW/Zo/hsZ
kS+lS0igCQRYUs2/2PelWuJWLEgvHTL5C0F26KzlJwsr8DveSvQ1Te1to3dOjN4/dHEWmf8wwydJ
GQXmzRjvl7kW0vOkp5hwz0eSXGYsCYcvWmPG8FPfwqlSfSDh51nBgsUdUcI0H7s0zRLzUOYl9o6p
DPkwxZtmmzfsqCuePrJ/YMeJQQNW//UrnxaktU4ksr+XSJtb6Vj+jSazL15K82ZuVYkVzdAuGDaa
Hn9yKQWURVRMjTUvLYFLzzfXRdhR6H366IbGCmMz2eG74bMsqMA6GrujWAA+8Nw7iLNsc0yji8Bi
gmC8RUAoKdXntxSF9GzsZ29BBp7mEtyrQhQD0kgRDkNfZ48e6KGQPYAK5YPSc0w6GrBhTWi33os7
Qu0RFMoGexUnpr9oNiFaxCYYjnlP5hoWDJdM4mpps3YP1xK5D01C6sn6S5mXWNq07aktkwrZgBdw
6wMnEMHL3xXOJtSBrAlwWGWxeQyaqrXvZx/7YQxofPLHHZFYwkn1kExtc2DF4vPNpVz6MneonD32
gC8dnxvfkV0cSDWXKjorMwAEfIWFW7M0r7Lq+0sNC45lkBk9beyC6n7FM2M0ntUNVdS9FNHYiuk5
EU97fuI2HScpwUKoNynPklY/tOcERa6plTHGHoTiv82RiecZ/jDPNsU55B5jGDbU1LEoZZYlOey3
3JZfC4lohI53HeP+zn8W6QmCBjpg9fWUZufIAqZUBPHIbn4zZhSaiPqNZTFSYNzkatIFY6gQQ0wR
IWJtVW3++0IPTYyXBe7vPhJIPBG4u6RQrjwv3bDzhFNmPDD8Yfxv/lxae/aMpO0c2F0OO1uBD12z
gn08FbK4wjNGdb9Sxd4fxZgm0DcWaqJfOPPcPnN42FytpS2qniglrU+AzU4hN13d3oIMnfWLhYPp
fBmDy6lBubClsqu0S1fOjY7x+Zci+kZjp3bFslda/J3VNb8CkkukuPHlvOG8ehnyiJv+FvbkjW7B
7RuNHPUwm4rWd2eIWUgnJlICQ+dzuY5A3Kshdx+ikMbfdD8tUSjDOOs7VSVLzcAJCHVeJKpKTdtJ
/UKRtfAKl5WDGBxEaUH2BBJX8gsMK5kN8rOaBuMsw67BcPxgi7pGFtMI96/p793i9esVNujQUwin
0bnfoFv/Tb6g8CajJOBCokpk1BhmTANG8CRhv2FIzj0HFWffqbjB0ZKO2+G4tVx3cbTuuALNLwsR
7wZFEInPO+mcwK4acqsZj8KuF3pb8GHdN5mpwyyETCDwnyGEadC7VOmkSBUYB4KHGZCW1bnW7L9l
vJ6cFT7yjkXnZ/sJsPgi8QHJrEbomOweclKYb4nzWnO+ktUuibvBTK+FTPoAEpPn4KkxXgSriPbG
ZhhUN3tjcvSEF1fhn9KHMFNF0+k8QM/o7cqw/d1WNfzeVJ190BUKinDzpO3yGn5Hs82Lu8x2pgdU
/0L8fGGvHlxDAzupYWu7/pG6MKYCmWuf9cichuGJFxu+7aZCkzJU8NYxkuewsrCL2CredG/2d9m+
BfJZm8gDM3ph6hamRELcjXh2OBAZaH9X2nHtvJH85JFlAt+ZLl5V81ZeX90VjDfiA9t0C7evCAXT
azGzrAWziGFFYBXsbuigc8p8TKZeb9j91xjVGzjityolrmzBlEyYbIFBvI2KVJRT1SkiWo7+payp
kVh5/hnqzuyUK6w+qrPjPUOp9xfEPGcIuM028v8sNd9n6JhbkycGD8h0+Xa2iFwYjAF1g6YBFWLW
DLFN6nR6/K/TKH+3DBfn8oD08fqng8VdrAnhMAn+RvhjEhOYt+lbwyjGKl6lbQ6JMLJMMWQqThs3
Oe0xyIFzRllVvkM/Oj1pDZAWKmXJbt5+pz30kCr536kDILX3IrJ1moQZ2sLWx7YiawNCyEbq6IpF
hGk4Sy7IpBcQ+Uc9P2ZhlWykLG2YH1/blElAkQkhgPdzHLqATauyX9FG49mqIlYNzDy1pQEbiEi+
Ewc3fcNm7m3Y+GbIfkb5VjBzexRInJ24Jyr57JuCe93trWTdQyTfdhWQsQ+5T/j7dz56K8nmr2fd
Wqj4WT5VVV/M+nSr9X9i2K2WXHvRgt9PtmGeIVGJ/j7ZbobgztHqvTgqtvxM5bA59e8J3op0fZWo
xSNUE77QaCSnCbLgCZCPM30nEslb0GTVUYdQWOPRTTmJYnuxoKvnaJ7XDqPAp3x0ZkcP4aO4w1a4
yYkODXH721cJ5/B/bdbvE7VsuJil2gi6ZUsIwsAhwAyrhEZVv+sUN/qhF2boSVVRFYJ1fZFsDgw2
PJsxuOcqFUVospPq3K1ZtmDxLUr6+uURekELfP/v8VlvPoPY5QEmSjXeoqVuBu6fte/pLMI0XdPb
PqWoUxre5+HcaRWNyLc+DkDcyERBBxke5e4S794kJtwVB3rDs8RmtOYIR3NMnQh7DtB6DYWmPTnD
xzD7AsH4OoWHKkvaAQc0KnIapFZ7KhqdsgFWk5lYdlDGs3BCe4mDrouFViNZ5jO2kDCfoPPNRfHO
aMPZbKL5MWa1SehDBFMBe42fM/nd35ud0eEoWJ974CPycca2j9+RqBNi2fhII7Bykl43MtwvCPa/
5QEzodnnScjfRmMSxzlQ3DJRGSvuf/vWwmnJq0nGJQunrsopth1txxy9ENBvAnyIkWbhiDoRWhRC
Fj700NS8hhLfe7q4p7BkZUrJVsaqnmOjZhxiEaVUQp+AWKslj6cEF6dJU8kD/vxoL8Qncv6apQOM
9sszgCIUpZtngLj/RIyxAho3Cio2BggAQSnraSgD/8sIGuK6XueRlleFsKbnMTKtphqvmwzLA2zH
FFZyxfa5732x4oMF+01j3/ULbQAovUb3t79OqJWPG1ePKO8LbMw+p8+laoBwyGukhMEmmKvmWl6O
ZOJj1VgmvV3z8xEwNqfXPz/6TNWlWo76wmivwj18fYlwEdqGIMd3OhWqNNHoBqRSSo4XdMY4iX7f
6U5l4zs459Kkxz7kG9fDy7SvzYNqlNRrb8RSMJfZbqBLWYGyzI0sR12NE6sx/AeRCCLYGdcBN82C
SC7APCUlnJpGFAHHvNFkuQdFaHA0mZb336cuyAalh0ORIgpjYbnyZjYLk5mrqA9BI3HzNLBlkSna
RS0CAtPZRRRUFv/6yhQ2zJRipTAGaUZguiBIbiz6t6pSjNWN07uaV43KezXp+yZ7rOt56amtVVNY
VadmUwcKoCGCeNC++pBLHQveT3wj9oXndQuTFSeujUaCnVjbY8f3cM7363lRIfFK8MBI8OgE2bcQ
MSG+AXm6c81Ym8SgnzsgijU+0PiVHZnt3UjlJmbiIQ6EvLyCWciBSns8868fdB3ZN8FKQn7yQtEi
Rd7+6kyGZXGVaPhOr+Iexa3Goxsw2iZ7mkgHnby1Dgk1Mgww1r3fyOmUrTtToq9nF30HWAAonsZ8
WYcJ39tEC1TESam6AxbInkj+dwJCMX9bfERKElbMkXtzTZAiBX0Wze4QB/eWRjUk2MIyaGzxMk0v
138u+IwEboRJUhZ3Rf7jRpGj7aZmiFUwwheD80EXiwTB6HcA1z7HKryID3HhlQxFT8QyC36okSSH
FHyZez1pQwpn8B+BzU5WrQlW5SEM85q674xPFcL3hR6+8OhLQouNjTIzVhwz0VPsGqROMx/pN52q
sp5HQS/Hb2WNNm7mBCOAQeUUJHKE2/yQ4qJCKJe61Qmd/ohezWdkIimpOrd4b81X5gefQVsFqcb3
DU7bc95KTmZ+EyeiYMpF3iKPQaQNmgYHo4apzLBoKKzHpIZ35YM1ltGcFxYpF3ZkCEQ1rGeEcQhN
O85HHzOGblr4MJhqSgkZx0/i5GUEyKl2QEofPGyMYXb8/pPP5mPHfxx4LhfN+q6wH1NOkz2+gCJX
vgRYt9J0hkJ3dWdk2Ds5uLtvcT6DU+dPXVuL7C9nJjleR7hXqRl9NnppvVg+Lhhyl8mmqGj7Ww5K
yj9/mO6o/cLB+B82IvfkdAPlWpwvA7s7QZR/Yuxgsh4JrR6hUA8zPGiT0RfTKC9TXjq1JRtksyXx
hTqPYjwShPr2LBCeTGjNrot1D4YKTqAfE8UCz7gl4tIxwCZG03Uv8IQHUSf6oeOaPa5h5gjvecQV
QwjBcmfxfpvGjsUtGm6dEIkJePYZhANiP32k+pUb0Ky9cijoFbJ4jphOAZjcIOxfYK0LOWi7OxQs
s4LgYT3oY78CrOW+gkSDmXzIud/GFnozGw9YLX07Y2eb7DBkFwIvYyeJQcwNl+DZBMcqU2BU7TLu
FX5aynIzwBByVpbKEwS4d9XhN/kUtSDqa04PEIT9Pgr5bAv5RoPHf5mFxv2Xe3WBJb9pzdxw/fV0
3ai5kf3UQHLJqFtfHcRNvR8GmK1CTIvjUvT78gdBk8vIiMe7lwDa19c6jS1l7wbkmIeIs52MAL1T
2110U9kQL0kNTGCghs7elDGnJVrMS+ZFzO6PKr2YfKgCjYS16dMy8n4hmb0nGQS8h9ms9i9B/ItE
22ZW72Q2spOrPQVk1MDZGlcbE6GN1u2qfxF5ytEvb9CJUfv0uRBKh1NpLurZcN7Yx53eEd+GXME8
Sfqsvh9YOPsqPjFjqMzAP+NNiH2i7dhAdxBVb5GphEQSXaSfdLMRE/RyiwxSWbCNhNn6nEXR1S1K
dstZVoaTz+P4l4skv3o9axkCzgmx95xNkrlYS7a6qGKEc9kjRPiT9wtIb8R1vMk/EAf0HkLYZfhQ
wX6GdzhHLxOrjFVRQhOFlByEbxtA3GbUXxDww0fMYG5+5r8YM94oVtWhZNA+xPsqxnXjmD7X/Hxq
l6Gs+BUT4wWatY7u22y66HjbmXTIdzw/gpcsmhK7c6DJ68fIfLv4lApinUP1dJB0mQxqnshwl8ZS
A0ap0/Ff4Rorpj8IVRH5OVO57Q1JMpNmAqWFM/Vr5hrQf/oNd6jAUJc/YXVqj2KDqqrg/dsYv66c
PnF20Eop81jFcgZDx36/DhHiWl4/iALosrp+yh9kvnphxXbVk22zUN5olzGbX3ANOw/z5zYlwix5
Ci8ZqIWsRGqXWAKj4CeK5npcO1jEf42O+TAPf+aptTmsnyT2hiyYtuUUbmMq2JFPmkd0yE9Me0xp
vHs8OpwwZFbdJ0QOBsUTl5ROw1fkdY+ITj29q8kK8vf64Ks/xfLsqQ8W1QVw5NmtVJQ4LfxXXmVK
EkhMK4lHRk893qte4phQ+c6jmf7qzikqzTjRMBtvFjdt0M0vNPdujFTEa1ydYrh0jqB0F5Z0T+iY
1it6+Cz6z9Ndo6oBwlgAFnFAlZwg+/mfY93yDq2dMTpdGqWqMoenm8kmHN8WlVIYaI0mkyotDNGC
J31sZDuTTpluHPgHdn8/eA+6Q7y8XFelM8QmOt86Ad25WUWOEsNZDIJcIV1F+C1nHcer5sB2Hc1k
VLpHv7bgA8x63vb7GTZGWFhcgM+O752DagEx7222Qw/oQPhAg5JMSyqJk7lP/QhJgqyeIFvKUkVk
9PG4H9l4UV0oJqmRDwWd2Ba8YkfmvHqP+By+YcAqHYuZY2ga5iOkgqMGIQZK0LTzlELC2hzX+XUL
3fNS74hmQGyus8DCSf4nk9VVQ/FjXbVAeJZ9/pNJEFWRJOsD1eyXGTA89CKAN7bT/UdKa1R/3oq3
Jf/BpC3em0crFAjiHHMdkUyV3PcHKS2X4+MkEGazP7/oXg80d+f6EHby3Z8HTtuYJAzyyHRAP8GI
rq+lTv5cYPZhkXXPT1pw/X7cx9epxZOIeD5mQeQlZbvofnB0wx89C2b4a+ko73O/cCW7+p8A2F7z
e80qQEzTeZf438Ae3Nh3tUV9O7zRPNQFgQY7T+uE7llac2Us7YiVgoG2ayX2N5Kd34jSBw7Xn5Bi
wBkGgR1YJmOM9V7ufnh/D1EoG7KTYHee1kA5UsD4Yuc3FHjSxDZMiXPW8jlhXCXP8xgVaWn7/44y
DWZbOJ7Y8v5APu1cjCamk3lWOvlZPtssgHM+nmDN7msOjsQoZ6YZ2qQjDRLq680Zy68T2nINg9q0
e0/cfrIyRG0J1UsCw1brxIvZrFdZMoA21SFDoERSSXydyh8quU1OES+sPm85MOQLu3cDYWqa1NmB
nFIdUJzzsmR8sQ7n+hMMPbEOnN5Wl6CJUCr3mpN11hwfN1iOJTPAueFMyIX/jLv7XkF9AXMwUdkr
RsnGB/oyHa9JH6nlz0vaANKG8vsCTkHlXDw9M5Yzabala23ij70yTavJl4U4RX11pqGxLK3YgOnG
AVwAawIcswXVz5CfrddxCOi0JVZNClh4VeYCrWZcNY2zWwZ85OIF3ndQAcCUQpvraJ48KdW1HoLG
aHkATDEk6KoDITIFffXrMQHWIMBlJPPxksQxvJ0ivYtbFheM0xrO/g7cVF2tQA8J1HPrmtHA/w+X
7MPg0GmGtcWGFwTAkQODNEGh+1/+vuPilepcLIRnWWUTFsgbyV+2sYnqUp0KttCPcM9jsAuztj/F
D4/cOdOi03f72AOnpQUhuZbpXDvrhqSSM3yomuCeonbU5PTTxXxZE9saZ7Xfdj51bWWlAs8WSQeP
74Y3Br583ENYtp6nO+XOY2TmyWss7zutSWGBTX3ElUMIj/lbG1yHJ1js4c0R3xOZoLiB9nDU9vkr
NgRccwKglLZ/RmJPjNV4Ipts3CniX89SffBL7Y2F2ISrO6UMFYBQp4t1LbWPibjyrL+v9DmmX2vm
mq/7g1POj7uCH+vHEWB0FAzN/42m1ESr5Nt88dwZdyQ7RatO7BVl/yTW/IWmRDe7JX7DdeaKVbOv
VwQotTJp6xHKHc5rIooDjTZZ7LFcvPzuPd+oBWazwc+HHpJAwnGrQgAqGGmn8aOxLDf7ysZQ9rYd
6nzFewWJtam+8BROQLNfPvXtySLZBKeahYVjmaeQuBumStB0Ndnid/XRyIYwAdMsq0qKacv97EhK
HbjLNFr28O4E+YwY9+tLaAkDuslBPjjr5bOYpPkrLoDrmGpiExOmejamCn0dmFXlm7HbOvfsqbCi
KG3iT7gtIjk6Ppwt2w/UKbIQCovGXYPG4QSxSD1lKBiksdWuyoqlf14OC63fI7/9PIOlt6nUzPDo
Yj9lbxq3G8SdAVSV0AUXRqR/ywVmdrtDWYrlSyr/gd+/FqnSpn0qGA0ybLl1LzIn8vyIgeSRdwMI
zTSFODohcnJJLpmlxscEGDwv6Oo8UPc5zTphmOOTWSM8OjsCNnjy9XHsF6E2Cquu2Ezx7HmkKTcN
obE67zvu+6/jEDQXn5tA4meV3E0041BjXWcni++KKrcolnVSdTLsHOAqqUJaDzDJUZoMEqGbTFZu
L4M/muWUiHYi4OQYTZJkPTKCHNC0BwNQ7Hwgf0HrAHdvPmvVOxv002l86dsb1394JTr6imcU00Pb
BXLeHtaV0f+cRdMukMMwU3NuDTK4tJn3haAjBSDBgxLddzmgdWQHU9BlcIt7Nf1I0Pb65jRkJv/s
NnuAw3YmyJsJ+rlJCINOWzsm58Cji95GmBM0MaIsS4MKYMTAvpuzm77xn3S2Xk7CgWQT82cpYtvj
KelytE04LnEL+C36cgyfq+SpUONKe64aoC1eRKyB6M8R88NEgAhdx1zaGagkDhNu2SdDGuZkj80e
YJha64SxsWr2c09TmuaKJrwm/94H8XfVFT4HUYvvRihaqP2jD80DDNY+pdmhTJTpkvXrfcwwKeZp
dYIRXQhNH5n05Gko1j+WFe/LCQw/iJX3C7WcqlBjQuv+SWInPsWXuvBOxE3ThlFyk3QW36bP3lJn
5xUaJW8FKI3ektxM0ffvAlbGD9UUm+QW9jveALZsTra6AFNlMX087w2UMOm1LaTEDy2CcquM6aJV
MQ5dz3obpMvF1w1NFjrOItSMktc+qw7z0XMQxhmhRA7g1J+raEXXy9EZSaNAuQwcEpdk7GdzrsEC
4CEyu0rUM8yC3PJJbuTIF+cqr9PHLozwHdjtu8Uogvk02P92k8ntzSIYYCy6DN9gzxcStoJ3kvSx
P53nqGgm2yzl4D1o/fJM7T8chvabbcrvalPiKI7MRTN4tl8nBn+QUGLPZgBqTnhYvL0cN9bNASqg
7RGa/eYKshNGIPxDf5+uzGSAqb16r0Y/ReTSafJfdD6mv81WHoEWqGuobwrCXKZdUtLBIVTt19ra
pDNgkFqxl0Bk3gYKIxsCn6QuwGCi2tY6U8HKPit1wgAC006jn6yfNYivzfQ2waOaux/BSk4aU/rD
C/0ykx69Z4hEovOmO70j9ObsFY63dBnW/EvI7qHzkcqyzsKNO+4ayn937aD/dBsgIdiv+HI0Voqn
VzWGL81ZaqbArcDwpMWurTaicoIfP52YfLK3gIkmYfOXQM0WEx0P/EzqRQn6xEuQRfOBKakypKmQ
Xl0RGzAF/bdcyAtwHIOi724nzKK28oUudn72f1BLgFU60Knrwi5Le98Ooy0ZdYgJbSg1W+70In3m
82i33DP3og2lbSaYxf0Y+4IYDmoL4E49yqVLX7DIbb2fknBNQhl4H8IzSMi8nILoHYsSQzjaDZPl
BkpDdyZu5hVFNRu4ficWdqgJ0mc/0cfMLqcDaSnqTEFnKuH+j5hMyrILiZGrQXj03AaNdU4vlUGs
JqcaNBdjkgvUPeb9EvuN5VV6IoyIYxC/jAABkTy/MmGaDbE/50qmkDmDpzFzUNylr6+lAwT0b8sg
elphuHKrZneZ3Y+5tW8KI0Jun7OUHUz3HpeFQAQJXCR/qBdbcptr33EpsHIVBQGx7LU/7V+ZwiCy
/98XfwOxl9by1BGEuFlLZJAG6sFhEM1z0rjqnd6g7cvkkBq1h+SqA1tgMDjmashclpWZLhX5O1za
2jC2YXLEvlVqgl2zrZWLDVIsIn2SrjnK0d52pY0QPuPjW3E0jismLEhUVU6GICJsVqJuVtdMJkx4
KXHqKtH4NKdByj4rSiVZJNDtUr9FHB6/sqK7cZza8eefeGEuXn0S/4dLCJKsYsg2cln7Xr8XLBO2
wGBq7PNsyi/OWdxhmJd6oQUnF6WpIPP3JrxSe74ZmUnOxT/U7cWkVLdHTlEg11Muqz5fWnUSswnB
LvFyMRygSuJn63LwaNOMnkWChmIE6tCljblSTGFBW7NR34IG9wYIBNMAD9P+nDTH6II2qA4112BO
l3iwztaO4WYrpuUHugbG8T8H+LAGR8WvyH0W9KegtYDrg2ZuvP9IQSup38UXOoFc7e4WSM3W/VYJ
DqkeDT0Mif3FvEsyoEeyAE26rZpN/y+C2Y2EPCQ9YqzeSRYY0V+xJa0q90S0FDdnzqlEZ8qwFj8F
n5nV6J8QyisqQGvisG1OYMBk0bi8RBfUyziEbtT9UGzUaFgi5fpjqmSbGT+oofZMRrRhmBCh4eKH
XsK39gGEl07dtNs/ye2Dj3/B+viFLL1gAn7tOFAKaXihlKSN8SrEn+RT59e/e1C5Plnc57jB58Od
WEllTIEHgjJhpunowWAwH6EytFRAlmgCAzUIdfbUU4FtnKk4ZoGbWgU9V5NNpta11Z6N+7ume/hc
qXqhESI92+R6NMYfOGBGhMnoRbXJmTZxuqZ4XG5lMNdBOQPgcyEnamealk4sWs+7+1BGgcN7CkOZ
l2pjNG6EDQJnjH26ZnNRiI0sFdkw8ltPsHjI1jWhVWi93tK7O5srwTijQn3BCpD5I6QQyXx0Pq02
UdrZv74zZ+mnT3bZRRL2XciYVNChDIo7/ARlgQhjwr4w7zFYGW9GngRN6HDdmf8sXn0iMB0RvrPv
EcgfIQIKmNKUbl24nN35Lvwy5/isKoCHaJE4C1Y1NP1233cf7EwkXxiy+Qic77nLXHlZ5Fk7mZwL
wqycdogOmxjKbfayVeOvOk2PasghDZZ2Oi0+Y8j0zV6c++62Xa95ulvz3UV2leexNFB1jB7JwI53
Cul6cKX1MN24cyYDTpjCdWkScR6X7xzLyUz+sA524oETxog/y36oVGLACzHeSRt4JFNnbp1sLbJX
cXZQeDWlpZF2yJEr7nNwp2ZshSSDafTJwd/MQS4QlTBFCYb5J3YXDl+JI1CvhpXB8E2Hkvj0cQ1l
r8xnSmHNxSrJC8fJpPnDjM+E9ZyHkAIjJg0PGaDGF80lEA1t88Bs/+DewIJE0+C74iTiLlJhpfc4
oVewHME9j/1ITgMoxkMMgSHxlR+jJqJTVowCI9a4wBU069An6RW9z96n++eM4wUDS0cYOFGG1S75
Ec0pppK6x/KoTFzF6cXWSoiPzOLk4vMzC37rQhhlo4qPd2P4LgMIInWNK0YJjaKWDsahbszAmD5G
x5lwQ67esGCP7Ya5mdR6lNUC5PsSEXycgCzko5iJlZbEPa151LhdSesXyf+mgK9nqADTGZnlkNHn
yEIxH4PTuLsXugOZ4+i8B5WhhodkpXxzGWwo4fcvBT5W958aCnYXNZFVfZKcoG+wjpkijYiuBNbN
lv5kxhpxx7h3fmfa4/Vd69J7j+DoQCMawP4yoh2/4TDaoW0rjFaSFQmeknFea1vzLzZjlzjGeKzl
Jl+IO3j2t7xR2kAr7Jz2H4HicC8nhJHyC+PY3+T7RvCS+AhQPvFbyYrImU51XQDfdkYIT1zh8DW3
F3TII68jmtwDWEhTtRXcI1121rSihCE5apzUkXKvOa6p4CRvx8KejzZNrkQahbyfU1+ceecZQj6T
ZOKuqShdCwIwPQ+cQNAdImuIVlXzUngUdUXxrjZb7tksWHEikjdg6erI3q+VPst66E43W/rgtt6O
k3IuGM7CbOeNIT6CmvXosEmSeh1G/AklqEv8/NblCW7enKRSA+oal2lXOPdXFY04iFH20dZ32AZx
0XD+O2+2EVtRuUFwDATBWbIPiBcMSsMMnI1RLyOFDXja2ADONdj1b0xudgG3zMU8uz+1klVrA8jc
Uj4CBqU9ZTXorGwB34xmHRe0RuL9sTf5UWb7Smff6ambvbGyh+p5KvJ+C1y66c30SSNXncg0F+gY
1Pz4MAjJvD7g9YrW+P0ktcfxBnOl9EQ5XQnDfmIIvCOMp3vCmjV/2J2Glx4YlUs8AhihtbqUiZlJ
xHxcCRu1sz2yP5g9bkIjPnvB7J2S1wPa4Rzm2Xl1fB3HYgDvpeLckMsCtIise2fj+gRoN5MCxnU2
5MWelfw4xb3qYJFYw5pUJ58PA43LdN4SWV56vWQ7rejJS8HTgsLn6/dIwkufFK4NOX4TDXvOyU6g
ZZRjTw/odBT2QrRyuiJeOB+zcAh2AXVRbFrIbnQ3KB9rkoMLRKfTU57KzSJu6TZ1B6h+8FmMRsM8
Rj2naBbH91k7wVg3bmHOADPHpsQtRB4JfJVUEXPVKxpi9ZwlISC7iPvE8xmBLo6rBFIdyosT0hC3
DOghXLI5QVAYys5p9yY0OFlmxaxKTyFrzvXTpci1JeRqKWd9LSy1xvLkxhZ4yp8fFJfCr7IL1qGa
GdVArFs3XN+TqSzXtPTZljTi5jAW4WyaXBjK9MUwgZ1/OzmAKxwlGgtjZEkMTjlVUJlEWTtP8qKh
BnArFVr1EVG6afkrpCPL3PuH7tw1m78t9dcVZUzUaIj4acjUXtF9ZSuzQIn+BUwTQhFr9q0L8lZy
288iwC3EgKbZL0b99YDSz69hMF5POujJoAjPY/vm4WVWdrAO4g9EJAG3OvVGXu8qaoosw9LykU6y
NZeyvjBJLEtdAKb/7pKe5D0IqyJUBkZRF5Ff9yg5GGIVvMswB65RuOuLMt1HTmv/wPtUU1amESlk
VozH7INa0Qzm2ZpR/+dojlNS0sHS+zmHnJLPdxmuKlxTD6E/66gZ+XGVPJcZ/kec5QjLd5CxeysB
UZahrk4OQRTyQkiWUm+FAS0DM0Wx1EsW5U4wRh3H0kvIFlGpt1C8sVyNitNDDjcNq5j/DuCfx/se
LmItl39tpdQe6iudIXSaPyISrhL1zCD/TIp5llri68ufR0IGxuGWKClYFq7Acy0yptqaxJi34mU2
fOuT6b0G5novdpDUHdWofd/CLCFlBfeTLd0zeRycyG3c3XwPfsLSx2dmvAeKopkl98Ceegnu6jq+
WBBKRmFFj2AOECzulM+Yg5Vp/rAmbRDkk9hTpI/OlHcEDY0DBkT49TvD3nLkUkZrD/RYP2K2jxzu
ph/3wVMmiAgyr1l8GRD+F+4CPHuJBVBn8n5z6nYJco3g8CzI0W1PfWnZ2GbPIwCMMqGNvkYHFTpm
eVoHorB2uCjLNpdHoDq6TwsoX7PsfzQ2LKoGtGiX4rkim0S7CAVW4xKU9rddn4ZGMs4iY8re5Fyd
l50FFAXZ9cW6oURdLN1dWIsYIMHoOFWyTLy2vOkNjo3ldAoVilKqKsgQbInQKNRTG5Exs/gttE6P
wqmhd0nMPGYrmp6a7SOtYJY8Z0FUBgfwQCVxNJwGYp4ofOUaGXMWcjW6n6Hz/clkb+CcCt5GKZvr
KIzsRPLwbBkLhKIvDYEnFrJGgqBgxGQBGI01eCjuSri19jVemR2+gutbwIBCzWuXZwMfDe+6sY7f
DAj1tDuL5pPgdeVeSxYKM2wS5+qG8K8n7d+oyrhTDWMDU5vxvUbfTkeZqXnzhI7LaALoKUx7slNy
inWJv+HFoq9+NjnNfcu2SY4CJlXMEmKikckgze7HTV5wS4lBLaWjlhpBbMFSEBgq6tUxVULAQ9xE
+7A3gaoKXJk9+8tEWlqCYkGTLNd+tXiMIBlH4ND8NgyUPXfjedYkUQVPbpbjxpikrs2aiwon7wsc
pIBV3lY4DFqGE3JS1aBZE4C3lm4yYXRfVhtzixP1EueD1yRtn3vC5nj2R+AqSIUV1hzGRjrr7I4Y
0VdDsFSTfrRB3LKljp/sglfD+SsTVraqW8L9GHlvzsaNfjhGF6B1Y9FOOxC1Bk2MwWePjqPgHuvc
BhQB9AeEPNMiJZDPPYSMa/7hbo2D0XD+nVHrImWm/5t863NUq8mEq5QCLEUAS8vZ8u4Pq0bZuU0r
yM41QNro4QP8HpQtUe5H0KRr1m58o/pMi17O7FTsmqwY2R6W+LL42ndWWujQFpTvuMIJX3t4mKv4
R2wlQqMoVk4+hQo7FdphQpLSjNO+DRZJ8F7e2NKQ/JM5mUm/yNHdbeIdslW5XaLpmuGlPgSLtOLY
oTn8mn/eqLZ5HXJK1aBAvNm5KRDfARx0tvsHOkk2mRkkSmon9pYzwdDskL1+rm6llmGOdtAWeqB1
GJ5i6AaqzUvE9M+nJmMsg3NyRwxACwI/yt77m+Ot2suVHXVPzVTYOHODOeDjSFr1628EYLGct+VC
aF7s29GlXZCfpTni0Q0XbGot4FLjsXgpded0ZvzSy+Qatv9psN9T/h5G+/I3qPTISyS/DfUmqoXl
v2q6oiRyKZ3Ci606wxbe+wATWlxej6WZU5Qb3FyJgp0EELupi4D+dLxSoYF1T/9l8V6LjeiJL2GT
ot5LfPOpsdny7ELZZYPV9vnvsmIFXu049Cq7oJbi0xngXUqMInCkixUvR1KWJIsCc2O6pHhlXO8B
aqLuM85QIqmWzuta9mSTnrS2sz0/sDlYfRs56T0OByUEB3Z/GpCZTAcP/hYcFSqg0jLvPuV9A6ja
lx4wqtcxmX/KS6b33GmwwJBHPTovTM0SNTW4j8buJFfZ/5TcKVunxfmf6VQrc10qOHAtdK8zunA/
ixlvL0Z4B3DlzDefWlMaerHum6qBPvN4WVB94hfynYijrz34jAUrUVSd3sp3ZazF5wF7ozDKhthg
3DHpnFqMHos5k51WD28IBaVyKSit0Xt2g/qtypchgsj4yWagRTbHT3QP2Iu86q+D3rDvkvkSU59Q
nIvdwbUG4IZB85joqmlwLwN6EOFA1ZyJbytMgVMdroDGJjtBGBVlwHV/gbXbIH9U7fwJGhFw7Vii
kKpZBaQbYAieCEc2lr0/k8b0ffep/OrNGgXsgQFCLR3qBbR/qQDPB6GSlr1Zm8AHeyEe0T3BjF9B
TKhUtdFCBph7wRjzNFTPOMr81ON4cNsTHsf4r3LW2Zgn5Jza4ZzjoY3MlkFViFKkbHciRjueOKC8
NYZfMeJdc3/N39Pf8SakRM7XIgsVUxCuG7oEA9E97kTwo555Ohv3QFQr7LCRAOgbwd5g/OzMoar8
o61MDmXbdoUerWKO8MShnuGZqRoDH+QEtR8pu2dCwi33iCuUHaCGm6bz3HeF8G5Jq/00n/mowd+n
5BNDP+1FFZ0rajU/7oKEdByydrt7iA79I60Yh1EzPJui0sBbwXoL09u+oOb9lKv/wM8kNIKkEKyv
VKbin/yHMtpDqEdK3RG5zNAR1/TYF86/mCvfAF58Q1uhNVmObk1lsGPVR61J5MGTRtyLdgfrROPU
JDLWopuud1ahmwkLo0BWO4fI5mAF7IEZSxljGCSTUMet0zG/yEepRuTjjdaW38Yi6clmzAy5NEmE
a9RS7FKw27J6TjAnmP+DWbxMoSyrXOUe37vV0mwqRs87ocMePLxy/Ezty2N7aqrTyweNz8rUwrft
B2pRt/8o/OfG38b1EEbd+QWfKqnZNOLiWcd7ODvCKlwz7qPVCerbHWkmSFIs3J54DYiRkdJ324/j
C6wG+hAn/gy5J1MIVP+tWLUSOfUgpE/3PYvFuvH3ABvu0hy+ptH8jQfImWFdXr+NFvI0gAHL2bbp
OBURQbl7Xc4MmZCLQP67+icFsaFEYdVfT9Nm+CYyb5MgiKHtns7+zhVM08zLwZnmuxBQzWG1pqhg
PTvUtqmYCIxTntEPIY8zC8WsJ/XnFmGeIqMv0gr/dZ/4ZOfS5kJoVQwojYtkaYlKLHIOuNcLawpW
uHp+KquHhH4DrKqMeWfuv39vhLSaXlS55pGH+SDglu7n79ahecx0fnDxxU//LMtUxnoEQ/i8LeFV
g5bp6FStq2obsAPHK8UXvyhPdGf5LLRVkDr3Qzt9IeLUBNnie4SJ/3Qm55Rk/nDOvEdvcB3iDy5O
jJ0SNOIzSXG10S/Jp7suHuishEeAVRseC1zszuG8rCNGdJq20OZC0Rphs7zA4gwvriM3sG+SZVXC
UJk3PA3Am49GwAWg7QRhaEILJ376LnebF3konRoessSMXJzH0hEra88QZtTsY0R84UnYfR0XCCVE
m9KdEeBWmMpMTFL82fNG+AGXt6cMQj73xsFwhkKzsH2cI9ahCXOqRhUtpuKS1NXqxRzr/8lWyqmR
B8t6vC1CewRWM8aLZWnvqN18hp+A9A/eQ+VyZI28pmyZnYvX17uNf5LqKh3FVqJPiyCtgjrUNvf2
03Vm0pERRw3mPcYK+W6qXJaZuASQu4uFbUYfZQHNMyfNqMsYp2A9SnI9eC95UHw7h42CTBIB/Qb5
HVTAFgGnu/8O5mFrqc8ysotY2r4qurWC82PzcWk2/AEuMkelc1y2NwZzeW12c03AaFjU/qAait9h
aRojiJ442tBvxItKcqDzpkXfpJxM2kGnT8LMvkuQdsBG1eMXQh4cWFpHd/TvxpwpSW/MkZFvnUrH
Y4aejPidtQRyhNcJqIU58HngU+GUGbMrphG2VvgJOEAJuoM9mKLZZc8JngxiIEzZzE7kaWwJn8YN
Z/uywcztyq99OIuEd3iR9+Tu/Z3J7Rt/lAGbrjxsXqoNowEXvRCuIGWbfR4y1GX1LBYtl2VsUTwg
mZOuzVDU0Oo5yDSCLehea7zWZQI8Bic4YNiPuVXAhQSryqcxdvlO+J1q0NkCJ956GCOOEfYsVKqF
jJibwBFfAQWJL2PjMf/PHp42fv7rb6K3jE6voJ8o6WzWd7TpEycT57bd3QqQvCUhuV/t/N/4W/zD
qSIkFQt7hRPaZPL7X5ATbCPJ2CQAfe65+iPfEMSWXCyqoWNXN0K9Tpd2a1HQeRpQWPppC3OB9Ypq
c4hgoOzf2JBfCgONqPmDzh6iEVMJe+lXLJI6ZEg0ZGYnw4FNvnKz7MlQQNa+Umi4HjiKbDSDAl8D
2FLdB5o1fqVBjYJ2P6pgJ1kZgjgS7Z4H6pdF6w3gQPWC0FXs6qe76EtWJBnKbCj9z9/SmYbbaf3C
c50BOEmfUE7wZMSYsfdGulnF3Dj118yTdaNut7Db2lAYwkIbcA1oxcwyu3Tn9OpnNB1bSGnM5LbK
k5j/RaF4wtTo/KywlUMRQjYhJNOVc2pvt2QEKav7C5iMCHHPw2mzlds0WxPRiB+yx/ht/lQQlrt+
wCzzhvyAfv0RYhuTluEnSyub5kHw2hGlH97uMDMTh0Tij0yaRl2HWNKk/ll2OadTQxvy/b3INxcJ
ai688f4OT5JSniWBk8dV3s7NOmOb8bThb8DS05HOtWjyRNpbH1kRnG+aG/1rgkzSnQfGoATyND1E
Qc0KiFCXNZAE735kGjnh7WBYwAESh9FQ3zkP5m1hNOlTlg0h7yTIH9Nrbmcc8TlvSc6X1VFIXJw5
uwDz72MojPn/17/m2Tb0CkAgUhTxxpjRBYfEiyXjCxhbldgNmMe/rXc5V/eUY5iDrEQ5zRDJhv3O
x2JiWgk7uA2IWqFLNTnkR+F1kvPP7icB+BQelcHZ7OIvfmiH4M8GZUJbCv1jGgYnD6VyPOSInqVm
A4i6f1aT8oyUqYu0SGDgozlyso4XBJihYoizsIm45+XEQDwwtgm9Uh2hr2DJVsZJqmD6HZdwGE0x
0d/8Ui+cUSSXSHYqtoEt/nhD87+0Ia6F97hbrFFP0RSTAUaER5zy054vPWWbTw9dRBLO91UPdMGv
5wYGTjWsAtfp4pBYKhV7SbZusHSb4PmrSnRG9Ourmhk3sFSLjpfmEoAP24svaVnNQWpxISoeDF/2
YGFgVbbtF/JcBVLmDK6wQfRUpZ/cW6dP+W8cv4UOb2byF9mACMqtxlBFAUcJtWmqXtautCtkRna5
q5jUj5XnT9zO34ZXSh8nD8gc+F797M811AonTEj3iGbieCidaeD3bkvAoaucBMIoGrsClnFi7R31
3LSRw+sFISmpk2EUfTMCVD5Uw39CnQpavsrXaqf2vWtIf77Ixn6KU43lVR/d3nrgTrlrSb0/GVrn
qbA5OWuAql2cf2E5hJVmRSaZdrt/EpgiopNjsKVi0/H8kF17JqpGHKTthPP4RRdSryv8K1VJYxvB
1pUZiRchOtRMB1jVa3UgunsEJ45D0aau9NR38NvZi7aGnQsjmHHcDCdiDFfmdKb+wv6QEN86+efj
4mOtx0MuxQkAnaV8b6nilZb+zJq/v092qcg9t1F4rhm9IdrW+IAcUnc7NxZIsLjTt5WoN15hGuF2
vXe1ha3tIL48Mn3I5rkoRIkNE34WV1oMztxESfiTdalCZvTVIYF0H2xBj3hE0FExOOoDFtRxUjz3
3D9bbgkCx8h77QFsHNKZQuyoYrya21224bPpPGSmLGjfWQdM18NVLOuhaLKOTd4lv2HDQj7cG8x+
3v+YfEM884f4AtU36b/WHK0qAptCFTIQV6MtR3npbDs139DOArxT9FcbC4hLr7UXHAizucJ6UfwN
qFUFICW8f7WaazY8ZTcdgTm80nXNUMA+wtvHGt3fhsVF0K4NkraUfC6kJskM0Wpg5hmCZppq/BWv
tM1jOBz75HHwRf0yvIhcQmrzSjQTo+cv6azKjZZ2PIHnfKNOl0UnWHh6sTS/qGAmwQEnrkKGVEYU
va1veDmArogAKBdRtYlPNNTrbkZEKnZZ1eUcr0K6I9Sq8m7WUF4uTPHOpdaTZCXl1aeEGmXXgvV9
U/waXDmzUNWrjza5XRT2F0Oo2DN1iOaTnb14Ccff9kUrfG4eY0ZufDGsXLATbc0nZJAZACidy+Q7
FWTRdfCwD89OoPYeTRgZfSVrhSsqklWu4AYUsiTGc81pcJUi91RQNnxg84Et4qvLtrNwufTy9Rqe
CilBJb7lzIYluRqpkJvxUuKDeYdhA/XXF9SV7W/tJCYO5Os0t0sJK0kuL2UCfa7CZFWg2yoZWHIx
vAOBUdm50iu6JLuihY4J5g7Q9pjJ49WrRiF7RNk7NBjpkUQDV+xvSTiXP3W+8eqyRI8lc8oIdYHZ
A+62KgWzgL0VdBrfpNwYCh0wshoLU14y8Fp2Y+Nku41WBOdoCqDIYl1cmbIOISgjcm6X+B/jeDkK
EXqxoRnkbcomwN2ztoJRdzGIOpIllCR7Gqch8ZhBT7qavf9y3LB+hM/KrgXTQ74KGu4KMvwcKvR0
j1wCZ3No5dSFUeEphOIQHIRrPU4EeLldINo/aXJzT62XGQU98VCEfc6fyUcVU7huTT4/H7ufu3pQ
RVWqSpmu2zZSALzkd1beNQT29RAiq7kLFTwO/8fhR22MfYyQcCwcWz2tD+qfKXLYvmLwmGggvDXf
oCs7yhsvVJqdbkpecYJd+lWSvUbOal2uJwfjJP492JK/vXoLepyLnCsLmNrLiRsoBKbS578HWLJM
Zoi4Shmj5ShOK0L469jZ3z1oSfIeHd9Rlzi/qoU+kKH/eahvAWkWz92EUsGGmGV2cHvJO7ORnxzy
ASKdpvwQImDHckh+xx1TXvNlgGzIsFlMZ9nInat3TtqiL4BbjJfPjcJeDjtB4IDJuR5FeBl/sf4e
fU2GyZh3KwiBFaLx6N0GUFlWLJ9nd+MT9aC3vW6kRrZuXmgMdenuRSfn/dXlbFmyEmlj/Mntbuj5
t7jioqRh69e3Lm2/1ut6sG5NFBVmekIOH1CxZpF1Yu5RAgJ8PjN3QvOVGNeC2Z9DWz7hYxB5WVIx
Su/8vyLldz89wUifqlbYk1ls3mRzumzYNup7JDHRUinnsmvAehkNV5Ge2YTyEi6ZAKVKOwRRz7tf
K9IYnA+wkGkC4I5igvpmB1oADmKWBjmzVRxDzNl30rhOoZuzGX8SEKTIZbAGnTk3cBYIsgK+P7o9
/FkAPuumwlNBTh7yynXOYmf+3W7A5FqBrP1aidBX8GooqODMc8T1ggKEXNdsOC6QCIqt6WMGqaSr
JgZ46gp77oYtSnEdnqAqt+yOLeG2QtpN+7NALsxP1ks0tVPkkptL93t4TWHczy5vKEuVcb8faSUg
DSJQizgADA/BATyprqWZHGaRsHiUfFGkahXAxFbT9swXQe0+BYdCNW+rdwt5gmzpMG1TWgx4hokF
ATxzSvHzGHh4VpipDuXEbGt9IUSXzx1mBmIpeHVERWYFs2C+jSP9VxfHHCq52G32juMLwIft7R3n
4aS3mtdF0b/rGR5XAXonS9aqFePpGrNmX0vlJnua/dzYq+eZDrjZWBhWVq0QsMdxwwtlgG4a9q3o
PHXCE+oOzPpfon9RjZRK27+PmjMSK2zuKGjFAT6cJkwFTqB63Sjxt2pMtCOkGl4Lb2tg32YoIMYH
i4JXZCNPfDd30LURjvKsxll4B9Hj+dYIF1EVkM+PaZNYBwv9UlImTU5zZE8hoVaQmKCWltR+ww6/
KzbBirVku8p8/tDX2nGciv20AT9+Obg+HrrtZ+Se3FJwzDOEM/HtZ/fiySnZU33XIV/VueOvLsyp
hLNvdpnZj4EiQ55xpNi87XNd5tLP+3PhU4NW2H72uqfqObdkhK52FkQyzaruxskFX0LeIw5o3FOW
OBxtGVd3nFXd98Ivc7Vu00Q2g7wlwL0ADN84ofFPIE9IdskKpuUnngFAxQstBJcLEOoXTzGDPC/6
9mLa0bC9vWM6t80z641L3OY5pazpevaa9rL9834LBXN1/t13M5tAtMirAbPOBlH36uzjGuMADY5d
0Oi0WNdetIBLaqC8yg/6cDK6JSEIA4uyDqBsr06Nr70+1keuKgmabngCAb4DQJfwVKPIsYoGhBH4
jsBy/4YHA7lTzu9zDfp8NbN3qiee2QE28Zs+H26kQPHTpqtAPQRCV01ofdV+ZCzd48fmiZZvAgfc
aAmLfe9n63rvQffsk0gkhfn64buW5clp83dgDEyrM91dz9peqv4RjupDyTtzuVVdO7PkMDaiXioK
ggmlQ2zl8NRYxQ72CvaVjXeO4XWSyYw3LHfqi8mG+w5rfvMIV++LDT05BHo/8WZGTFOy9sZxbEDl
146LlFp/qXDloFjVnJ2zUq2KNeQKCIaeS9fnnnR8w5OLD5ualdASFMa+3SfcNb5RFWeAKl7mjuhM
nnvlFOGB1iEQe5AjBydq/b8ceFlY0d8/leDyt7DKzE/HM7LB0vN0lEfW3DjPzXS9DjRWUN78Rcm2
+a6D0iyN0Mo5StKV+zdHl/7xIA7humZdpbFX5OoCGvu4R9EJsPfXcxjC7NtUalUYdXjILc0THOrg
rPW/lPiWiSH4ZFK+FoDfpyZKbC6IamHpkWhZUEuno/1enSXcMSysNbYumxKtJ4HJWT1ge1nNBQQe
vrxtdYa2D5nTL6u5J07FLwvNiwU14wQohCIIRheSEW/bcUhhy9Hh7jTMofUbeK0fKy4Vm7mMRSAS
TmCT4OWm7Zo5xZ604Dm0mbc75bJ/xrVhIEHFFEbDwL8AfyaUzqWcG9gpe9py4xygid+4+CrISgqv
8gvSeQ+M7Li1A99VHVLG0PJzPTNt2O4fgqHfAPl6r9ZMjuUG3JoofY+axmS8ngMP7p2V45ZBGmy6
0V1OYTU2pu9tA7/VBap+VB7Hed+WEmhgIvs48ktkW6D2pGEOSEmeaysOjUYctwqTu36myZzkHIY3
lAfyMn+ULB5d2tnPb2GuTuSCYWi/g8qBGnzTXWPHHRicZCh9CSILBf/06B+bawKjYWrFAw7nX2Ff
hECWF29YfW9diE7w+aCdotmyrYaUMLZf5eRYZT6EBvBg8DcpiPIM8RJru3PoNK2aBdcBgLwpqDNy
2M/6r7YyBMZJ6z9H8yFk6Vea1OnKTzUAeMJbz13/qcuMwGJzeSPuEWwlDWMDVuM+Wy9ZafkCOmJ7
fT9bT3ieNhhsuOcsJmcNyYCsrBxhWnsd8pxO52LF2hpru8cgbjWuckVERozC3oKD4jwJ636JLr11
FKUjhncAsQTST92pAxD9oF4DAkfGcibVCo4573reKso6cxJLq15jPoQRdm/AReWfS7XcvgmLJYj3
GaARh5lh/aCbItDCzuVKy+qMXF/cVjWXdHkAmj9j/dY8C6Ii9PfbJbVRMq/56rPWwUYkKSa08ClE
ohqVcBvX/WGt2NgOojYG31cpy47RTF/DHOqKtk1pdXRPmuMgCruTCtXUws8DwX/YAnmymDCDak4e
G/ZsBZ/q23Ata/X6VrwET44YT6P2p+Vp+47U73R9hJszFiXM7zlSKhrjgiQBHApIER7xeF2PvZnY
5Uc+SsZ6Rn5VHIz03exxRhXBi4eYUj5UkeycoINuXdWpWcTU+9uRsYvDVOKK8NET5Lpwm5vHqckL
vbXlgQJqNHWjmVeEuY2PGTmuJLMgLTteIIBztRuCzdH6nbb0wO3jhPSErjBHGuPOuVJlXGmsXqc3
CtHzoXf8pUBVSpbM7p2BYhYKykNkP0uk1ebgS1erwelzjlF0f1DqscQdxA/WS5aQ5Y37dISXtlb9
vx5yE+t9wc5ZHZs79Kr/Bh+atNe5F00F9FCmXnJqg28w/lRe0UX537iRMcQq/c3XjYAQeBPQutvu
JbuccDSWef0hyhuHigDddnE5PFsltf0WG4hFASPWG1Xp67q4aT5qMs0nsytnYWdGDqH7ZPmMIP4y
NMcUgVTPZYybwj95AykS+4b0gZks8OyofxJ50YTtQrywenIkk/Raj4a3CmCFFh2OzwDqNIR846YK
QYIfBZ4qGdCU1fzKrCasal6ZyEVe99eqOzDXK7xHWFb4Dkt9T8mra99r8wy/IrKKDRayoQWbfaww
tFZr1Jx0cS1LDEN5I6dBE7rHionoPxVWPyLLlA1I3/n4fjEpvupmJd2jhK0flG0ThIAE+IVUnmZO
4praMbtlnnIo+CfQG6tX8w/RSsmhBF1jltRia+e0BDI4n6JMQNaYqYPpt8TDL7irnYnT7H9fjqaE
5VUYIWryK70ohiEFYj9u2LaVTSLRB/AHe6f/9hhf7AdWNtCEa3Ohcn64wPfv/u5VLG+GNlCoqt8a
T+FX12yChatRn8SqCOG9QYtInTmLXQY/obYZkAYZJPVBqmY2ufl3hOYmhrLFCBKNWB1DqquzcyDp
yoDz0dqReJmLQdWxoBJ/UNHM+/anD4wfdObsdplmjI4GC1bVhmWD+kyFfEG/7alsSEO5muixFmOV
MEmlWFTukM1u1OZXzuSDYBXYsirT1E/j33/jWdVUGhs3TWn47x3IPn5CtlPT6hhwZvKNH2Ti9pDM
/7daIV67AcJSsZWTXCCvD8LUuCx2NUA07JsRwaKjexgR+OS0FGIXQ+OjTC61vXr+s6hVZRJOWsnf
WzFecaofrUgk/EzSaPOg2WDAu90B3vceeDsTNPPMD6vyk5/i/WGZZMDKecQACs5ouKF6bIyvgPAE
gWCtLWpWwEx/GeED/VsE58C//hDrFHgxT4lo72q7TQvYLZVl+mdQths2xfHXgzB+81ATsDQNqcr7
dznMRjfd68t+jM0Upa53rqktgwrc2yYvYd0nOewMFsz7SOB7vZnTXq6Qn1LqQwLhPl7/hEsZ+bqY
WB2zvCMjBkAZ/33V/CRNRfoUImloNhDoOTeKc8fiZg4bwBTbC8a5HsXB+1ABROHKCBQoTWcRkHWW
ftHI3HyOXhlAJ7C4lPiIXXzEqolgvGsL4qigygshF2tsuiqf6ryJAZ/NTBWMGwH0CO8Kevifn5/A
rJOtiU2ENIsg28RSu2XVHnhK3ZlGUEXq3nKFBvyIHloPolv6QdnGfT+Sz+pcfu8EKgpkDSMJbK2N
jbzRuDo20o4leGEGHvzghV5AasUKAbmdsLSYxfZ9NwEq/x7lAcTxA6bzz3psbT3MLbUJgBlJUOQB
VWRlqKCw4nu+AJPp139wduTspWGw9mcG2TSnJv1oQB/HW5klakJIE7v2dh91n0uNq8e1MiF1aniX
QfvEBLCJUUnceJy6oVjVLXfbUt5zTVUO08zeaK3z+Jk/wX16QOVc2+ykqcuHn8uWxiQr4v9W8Exz
2zljZ9bhVvHLfk2Umt7Qq2eR24JeB4PvBqoPO9l7JLJrKJo+WHDggnQzJ5atum+o2OwwqwjgJTNX
KwcGR1/1987DVuumf55TQzHRqX/SnBtkd0e5bf0+BW5W3Rgutjmwg/tpfg1rATBxWx6H7Ovg4QVj
AQxIj2qPUQU11L294iik7rKB5/suVWkAcUDvapUTH8rEpgyqzx29GNAW7viSaeuIPbcsPXfO4Ong
2ftqpJ5DA5Hyd/72tqsQpvypyIRyyR7DM9A6PmSfrmFeRPF+VHhhZxp/rPS6nnk0HvQlp5HRG9cK
2h/mDk6mRnL2GHDaFTfyx3CYc8XI/vOlXRVQWvWyldGOptOKFzKnYbqnuIXlG/rJTJwpq5LaZ10b
i9f0qv/sqp+sObDLPbaIOM4Vn75aE5p1RWoMJGHAnQKYbJuKLkjrvLVL8fw0oO5iR98eVtAG6yg8
PG26RojLKUsXXsx4IadDjpgSebEVSRsF13Yl2DZFNxg6gnOvuC/JICCKGyVpva19kYWvOVnRQKeB
AhH426115sDDOaDY4Onj3jeklSIqvE/hiRdpL23swHjS0zWpmteHVgW8rM2nyNoaNH/Odc5paRQ1
S8QgbdXdtMJNCndcrmP9bap0Cm4ZTFaGc3j0qf2qEkeYltbgELMndW6TM9A33bsijT+Er6hNA/XZ
pZDCrlgCTSOulcDPVj9E9Soa/RXkEfkptCIRvii47QNUGZpKRQaJlzvZcmoYh89t1TapzoN6DJjU
Vbx6rrSaR6HnggOd4jCU/c5VAlfOQblsgPNmu/ITpg/tyrAki4MX/MmjtlhbCUzFbwhhNsvR/psI
RBfIARS3utNA3kzty/zpt6lxSE/ogMZHfXh33GyA4xxTopZgNf6JezGJFddnjIwBiQE5jcExiGpA
51e5BMZsNqwHoDQqZ8HDAJH4lkufGSBSrFc/kgleW3i4zvXKYu5TjesdVSNwBZkckfx96Hp6saFM
kDsEmWy3aHLOUskBO0VVkKGfT6H2CEa2MelmVhm6zy+f26KTQxK8l+15he2opGzxyz2s2Ii/LrFt
oDL/uoJwN9cqxP1EEie/koKzTbvujKngELFq5cLpYiuO9dUCzYXpOEabn183Lu4q1akG0WvYwPSk
6aHzGXP+KxamMIHxGAw+6mbrlqLKpmxGHwdgX1f54b5lJvWMV9fZE4R9o/FucK2GcHDcsC8DDNe5
JQ+eNt192EpnVV/hGXPhsL/sI12ZczyOGXqYRDneXgcdwBQXkED7KbnKkA/VC9+L33iKzhqS9O78
BdrpbSaDhKMVOn9sqhBLhwYLWxps6+1JLt2HjfzGw9kKEkySMWd1Y/uUwFHakgLlxoBrfCk/pgsA
a77gAGw1lfyPbGQC/zPWjn2lTuj6RkTgbznWtsjIHraWIF1v6VKyuPmreqdkuWuMSMRA/TLs5L1t
uwjxoFG3UM6rBP9BV/y6LEuy2EG7s88aL2A7FWA23kvdqMEMeRaW/9jHK0hQc33TJF7pZOMEI7aG
04wmmCnvkumAovBrMc82aoWRMx81FtK6UlVSFyZGpGlf8QICtDm71YS5aGkVvwfUzDvqZvzbzpWi
l2lmcT5AyOEr4tbVfMC1PBN8V6dSWooSLqgiQu0RZ7Izgixw0hoyTHZkHZKBLVAkx3xlXzVXfY6U
L5frTKPyrJZ7GCDMd4MVK3r/jq6kTKsnW3Fpelfw448Z96AxYAM6ICKz6pqyVRawyUX+GXoK6uqT
j9lmbYoUBQwU4boeu3oXPXycNx1dBlu7jUUz6lSvAs/dUeA3+I74oizco4rLsR4LnDyDeRkdvaGN
WLc3483pGRKcQr4LjVj21s2FpH9PVGhJknQXn1G9q8xwWilgxQ7G3g+KgaiIWogc8Q+ut4Dous8V
sYxGtaJ/oM1zjOgBfn9IMxUU7HnFwP8aUqgYI77dWWqveT3LteUn2dY9DtMx7gRZnW8KmwJ7VfVj
JM+BK4ZB++sF82eKkFY+MI/3tBqZNI819uLIyt1eUqlmbu+ujdRUAAOTMbIog2ifzMpTiG+5NCJN
Ph1/kRTS97xIgs08DoEshVAT1hxzUqetDz4kdtvfUguY4dl5AG0vao9BOvThAY7LO4UINPvub4Xq
UogBZvUcpR4uh+0+sn98bRY/sNppeqEF8waHdoPQaM1gnZcM6HwyO4GN48Nuk66SGFdCGHyWWbWe
zUoh1Bbz5brELEmaWd25Pgu/d5sNNaB329+Df4ISWgeSG3F9X3KeARCNl0nEYRgHvPEsPsl8YMfg
l0iy/xIfAi24egDRK+XvwSiIufhcKV/pdDxSBDpi0WsQMRWzjGkOx8UU4fWFoRj/4s/zMB8PDlJR
bbzuRmbtBXN+fdM9PxGPve4WyrIqmyctiVn913EgW9qccXjfuZE1WeRVvG26bKQpSMAOxNO+Hais
y6RCk9VoAuw7p4bnYx6TT1JVVfQuajR4fJWp0EDnaPtP8GAleU2ncSoTOtmdfQb6voIVTHGfBuFt
dMZznu6VZ62vvuelb2SB4aLqFCCPddP3wk0uGqVY/hDN19Q1+j68BTcOctACWjyXZ2FbtlPgXU3v
UCA5uaHmrYHSJyi94UWLD9HYh3LTRzBDbIp7kE9HwDFjoeBP+vyncNRbfMv3WyGpIzD6S9PtywwE
I0ANb0NyZzgx0EvpE/1ZrQe5HXUw0LU/wvBx0bS13Irj6gqdN23UtDPTi1Y7s5m9IxI03d8xevQ4
SNeI2aiEopz3H3rf6JLowKlb3NM9RJT950OuZgtIoOVmDVd5U9cWTnBAEhuGdY7v6jlJTfKN4Zrk
Uh45Vjj5F8+w/sU/UosSloBEze8i1vUyvKW3xEr6N6KXJhjGL73YUKuvzT0RO/bgTrmczJ3mbQ7p
0Jh4jWktQvRP3dbWdSAX/2dcTl5K07oNdyjZTPw2KSjXrHXoaCRUqQtB9K+/iB5iLk9fO+CKdCXL
XNiNTK4jiV52/KxQr6dQGgyfs79mRAJ2eRS2lmiGhq/CRT7mDUZPyMlI1AAochhgbliGf/ZID/g2
oLCSu5yG4+0yZ61aoNJiRsggB+1eW8nB6eFF/vbcmFlVHXX2sY5JWvC3FZzyuOgNpXmIjhG2OSqA
0m0jrm9n76n6C7TuuYULGIWaf04/135cLQzz5/g6fjoV1UNlxZoYLmfg3o7BoiX7qtTg3miwDidR
AUmc7NN5Y+CnBgcGtdZ/F4+/DWRzEZToOAoCNYbFpePGVBy/iqDRtoFfaM9/ScY9XvNcQF4naYtf
hXsw79ydFpIHTYx8fPazBzZtuuA1jeyG8qttaZj7G8dQPBpmQ/SFLYkARIojNXcwwEACUHnwSLBt
AoYxHo2Ee+Ht6MaGqTaDXlZzruLAQJjFRxoikV5uAIYDXkqxLi1TwwQ2pniXWBLe9sKQp2SL0nIz
VyTv8Tk2Gcivl3fE2GtLqBMJpGLLYkGWCE+/QNNerNk5JhQBQFLj7whP6AUt5HPi6PIa/S0YPI9Z
S/msbCbVGkq4u/xPIllfzO5/pol+dyVW7xU9XNdGWaWh80aFnJ/t9ETkEwlQI6q2FjwD3fptEXeC
K9GirWQHHy44ziv7BBEvOri7LQo051bKleCY2k7lFJexNVdpSojOGefWvgMBqEGT3mVlYCYPDfGp
PK4ULW1TPO/MiojyMnU2Ji5vmvwS/yKys2LdRNts5dcAs9m/Do1fcepS9YFOo4cRakIZ+u3wDhcx
mrGHg7n6BXDdSACfDWN3HsBA72G8r58Np3cLAUAKQj+VZmNlRdXWA8oKc72MblkAMFCrhFn4JKbH
pMZTrq1J9G4GfIPL3jLRhSLoSz10iTOvKOxyN2FvPqmsqvMrtKazZYBsDEPWs4OOSsVd6B+LQF/I
nbjefF+421n6BsnSB68FHc9NhXNgwLovPz++oLuGxc8fAPq4RJNGxxs91fkw67+oRnDq08MIFOea
vGgRfyBWhrIBwwhHRlrTs/KO6UfeUULXxm7JuHr7KeiHNX8J9+1UlATyQdCZ8PaQL05+D36oyZGH
EXbk+z8TDJeYa2YHpgizu/L8mm/YaVxoc1F9Fj+d2oYrXhut/j/SjfROsGG230U57Oexh6NJeipc
ENFKDGz4sM/Ly73HIVwB141M6ixAsVp2jO/ChXpe2n5B3mK9XdpcOvanBrb7cfebx1zfNgoxJIWg
wQBmMbkI7y8sbKQWkhcI2yg4/bRKUo+5IT9xF1rjRWKoK/zE4XrtsGco3hP7/MX/DG0Vf1TLkVhU
BBtteYIk0GaNz0thsXWstgUjx4ceROWChAYSA/46c4l+e1x3stdmw90+CEM0wqMze1uCokBSpdZD
ulvdBJDqGRNVcAnr5eD0eFiqgDGRONdxQ0JH2g8xopQNOx7VBR7UGVgbNQgvQcH2EdTWocMlLx+D
ocOmoJm2t90RYI/T91JzV+7TH71agsUEg6hk2uZEI3Re+7VZzhW4vqJlCQrf+skMBInecExT8vZL
xnC1bA5/7lYZUNwCi3CxG6juBedX4NfRMpY90jjfOsogO0/589mIGSoELj33cdqMszM9LEJGx3uz
Chbd3Vm2Ec71hE4AAa7mc2xJlbUdfGjKnhcOF4C3LcBKQjP1OnxAPCYX+ZTScUoWa11EiX8RW+Ob
P672TnoiNSdNiqCxOZyFTXHi9+cZQJmX10J+Mde0AV7oLgjWN6lqS3ljR/bj7baFrk1WkhGtwSQh
NEXtUOi9DZVkZJJCl0CS1zuiFLq96XNJIy4fVzHJ84RPZc3ABX9eQTniejOrJHtu0PR/1IyoWjZE
DTqpH8tbgWbb9vByRCG9L1T2iYwfRywgdlMrDlg3aAXz09w8Z+rP0xpvBtmWF8GfO2B/JwZi7DjJ
XZVaGCaegNDMR0P89BUhAw2I+8ZDUfUICtA7I9xe/hPHdqAhgHewwmpQ3hc/oCwGszinEFTHvb9a
4Cs+slys9u+u+TDuJVSY3I98Q6v1tNg76TzKivD60+6pGUJHhU5+SgwGq/fi+6l7hAC8cI7HKaVT
gVE3QdmAqHzcmF5uQsrV+kTjbCHpByI5MMTrkeEZ4SjVEj1w3j9YbRZEcAzrJ8yjFy1qeCtYb123
FZBN+erZKM9GrqvU35B+OTogmCFusGD0+giTxNLSQ4jep7etHoKUITiJJbWmkDzcuzE9ACL2XOvv
DPRmyaBYsGxrMg10f7CFpf37lBck9lvp1vfWxgZAjt2U+7of97T0/scfNXqXwKo03iQkAnXWt0p3
3c8cQsEf8W22gwUpzFZ2e5MxgYeb5xWcrsloxxqf5Y1zqIlrf+0pcxLtdeEQYXZLwBGYYGyc6g4w
k4S8wWs/udYLvlHgOf6LIKjdINZ/GSzAdzyPMo+l/kjp+Lop+yVYGJLyNuPTX3wXQogNvbkRJJvD
62iuq5lNP7R5XNHxWNKDyPYD+1ziepjlA90mjR+UQB1uwo4DGGP76y4vjpY8/d9WBH4hCjFo0gC1
FDmqJzq6FgD18vPb7dgZ7aGQq1aWd+dx8Z8+Pd+81cHymLTj9HmEdNoqGNG/2HA6EL+VwRSLZMXa
L/CddsSRDJ9c0c57gpAD/7kbYvFV9sfN9toUPmz16XzO6K/V9glPolPJQiaGJ3Uhf6nuGAsCexFf
mJPvI9Pzo1mhXR6jyhTKYE67a1NwhiMmZtTlMINHKaGfyPRCXauFxbXoqhblKUIWMuDs08TVdjKb
/kUcBqIIWWz6rbuRj56fzxpJ8e9HVnY+zJ6SdplO3pEpE9ATnt5VpwkZ+yWwrH7cKW+Vpt/ksIeJ
pb4Oq0pFg9jGiHTyH9rZnCfFVQqza0V5kNiKkGtQY2Md8J8YczUXdzUygQw5kzqc/nnGc0ZUz6VD
lAyO3NoapTBLKQMckLcEeipOy9vZwu069FOWhOFlcVVErYtbfIip2e2QzctBBppF5TfJiKjzqbm0
tyXez/sMXGbDQENh+l3tN4qnDI6/azyq7kfkyatP91kj1NYSGs1ZoSHRH9Y2Moij/e3yIB1+HjIk
2PaIl0/ZM1LxoZ6aPJnmiy9bNcm0ZYGpqnShitXCSJm/o1KNlT9AiStwQ6fxL7dzNMTe5VMX3AlA
qtgHA9oNjZXx2u1fma1mBJJe2gXPJ2ZAXG3kknXHJgHUHzBCsHdumx7GdxkGKGMmZ2VXYLmcIqHS
89eUemLntaY0jo8ROC4pbpyWPmGTsLtWc1wRpwHFpRHBI5Cdm59YY+cfUbz7E30jAJx6utrM9Ae0
HKiSB7Q6REkHtyGKEkrvOpHCdbs29EZcdROXtNqZPwOFA5E2obctnbit93V6Ubd6uwRnDpPzY4Cm
Hpor30RVXBgnT3wNaT0jtqOoWim+e/A3HQYULwGrzuxncgo3ZIdDAThK+EPl14tUEUJX/tAdvBIm
D0KA/rVEPe46s3t7CeQf9SHmMIu91M5XuVkgfJPi3LkT5zaX4JRkH/cZ9G9IyHz7eJZtA+jgTpS3
sTUXS2MDKxPV/tYfxFB4Y9OVOUStLOxD1wNuBbGQ5le0UnMJ9AMgQA2bWBkBDKXOtv3qILaIxAm4
iMRtmAko5xjtjxzH2id4gXrcDsiE83bScxmisx7jEcu/sVY2KzDEuBJMlcUhAHR7EnFXbXuzGl9W
wXTqCLbdko266ylNuWoKl2FCIpUZZ3DjXVPBOdvuGbjOpRKxBoe2f/G36IDSVH9C6xGbepKXh8sG
cicbCPnG2eC7ZsCiFCqGx4ti5gM2xr1TzuutiMRR7mh1qcLheXXpX0T+QjES5/nco3ywEDg5kcu9
f2d+5ZGBZIxLmajIJdQ/O2QENanSLc5jirdklMLW8hdLLIGCCQ3d1OclE/qQJ/rAp6SdVdV7Zrrf
pxbR9RdoTSme0wg4vAeJA4kD/Yidr1vu0tHEwnL25Z6SQ9XMw8QSwZbmPR3DwKyTI050i45OAouV
vnoWQZjYVOeoTXsreGXa60rncWtvr9Jk2weW00Cx/ZttA+ZG2t5WexrSJ8uGnjV9cr+Eq98QJDdj
o0RGaGAb7cH/eTulxXI85KMMmy8n9kNedxVWtrvQJKOGGP6HLrrA7SMbigr/zWYOFRUaWdxOfiIT
8kLDvjbC/K4Fi48Qd+3o+e/0uga0+KwlMtV7Mz3Y8HHhjAmAPjmsToekRCXc8SKtmBQE0KibC9+A
1a2FsHnusn482G7KKUwwINKQtIuf470EW1mTnKUpomH3wpx2Xkg2CqDqMchxjQHZJDKbgzj8hyy3
75A0+x3PiLf3gSbjvHF8nYEGmquH5lYE8x0T+RvUP6yHmGmKGj/rAvYp6U1ala0Xqtmw0ld7vcTk
q+PGPRtD4kvEq8Qix1turTC+83Rsrp/bLq7XZdMw+AkkX3OT6iaCvbu6ZpK8aCJEJhvTzt1YusK0
uk7wpZQFJM4RsUndo7BLtLnphNYYicxf3NJqnPLONWbZglwo3Q0E0nCAr5nBX9FrYPrLjJN89+gW
8huqmsede7P1FWXtiCoAAkhuGLIx+i8mmIwj49rGWTlq2P5xOMYEFTcDp2U6YZL/HMgQB8nP2Hj5
AsyEUKlWyFHEF5nV/1Cbk/FN6uOgmnZSMxw6HAmyZBWNI5xHqp0lNm4k2fAsjPSWjazGUbkdOdxv
nIxE37T8ensm9yEXXrOtvIjxpBddDzMTToqCQ4nvmcYfVKGGyLjegIEoioO9p5wjv/2U1ruBgq/D
/ubq0k2esPiUzBqoyhwDSi08CANBUoGkD0Ug4VzccYA2qApmFuiITCUSiNc470Hfxn6C8ZnFBMC7
c62aPhXZTb+a5de4uOkSK/nWb1jRfFKg8m+t2UtDEXXj4ygvl4n93A1LjAvfIEZAsdm6V9flaS++
l+GsGYG8fWMIBXxR00g2ySNjk9rLlSc1BBHjW2kQnCAb1fkwA9Ly1iHlgXesB9uZenh9rjOX/ZLH
AoDXr2rS0KinyXjnE9i9NZvZplMfcV3f8EL2bFFd6Mb/7gsEs8RDCtHyeK12Y68Qk4MQCKneN+sR
xyy+QPLa+bW734x6PV5UsF1pXzZg9H54JS1DjSZo0Y7NzuCYIq5CMBbY4xuhm+WpsR/Wvylnc2QS
Jpyr6BkmBJTbTL3ynH+XRxV3CuJwOAL1UqIObk5d/7R0qDibd0U++BpxOl0VaQKswrKjUT0GcROO
Y5V6Huex85M9aSkVODPcrN0aZEc8YCY1k/yEDVh2Sr4jiL8//h/QfmY25BuGCbhXsYSVM+SKrlV+
H/7AkCQVxkvrV0NGhtSatQ4N3nbBclv1aiEALZGT9aUMBAgYU08pyKhxLstBGTf8QwB+BwCzsrtx
88FqCQQwjIQa/HMISRr8Hbu09q1GtMDgMSQ5ZoTbLFnxasirUF89pzWxEqEM39mA+FWC630r2W7U
plWEPSHdme7pjFQUAUsqC+f9Sx/PYO4IGVIzoV5P/vMHCtrFixhLTV4zQQy8cqXyGPQRexZXEaMP
L3pdJejGrJ3/I86CUdVPUAjwzz02/rDtrom6n+GQU50BIR8inPsDA7Ia36YLIVAnBCwdRue9eGxF
gCWcE0GA2xXLUtTdcoxr31Dw3KYmgHFMQRtYXPsIAyOcX1POKNlYxroACnM7Chc8XMsKrMGAX7mv
oh6Br/YJ3hB22AdFC7fFrwjiHFx05YSWhSliy35ZexC0u8xgCoivYo7Qrc8/rZhR57RIAFWMD/aj
jLJy1Qyn5Rpb2u4E7262ETb8C46oChNzt3HCGKqUNqbM1mSm4fICfQMVN6qOqAOzUKhZDp0a9ccw
iJBaY3fnoB+GyuJ2jSYBZkeiDE9dWoZ6hmoxVgeMe2RZ9dPccQGOPANi6g2zgZFOhqp3kMMc6hnt
z3EjZK/UrkLxfYfzqH4LZI1dZIdplJtV65JKDnLr0cm3j4P8DklQxPOz8Kql16gTod3fO1rFk02w
HtD0EJqVeUdy4pM0GW5Hndvks4hPI6+e3WKm+AptPNKVntP+ozfTlqLjgvRRz4U5FeIRjn3ef82V
+zVHwlgLlNOZw6T9yLSsNDtmDvG6puvXFPNddgEuxN1M6iPBetFMzlDTYhlFFHdY08pCr4tCgMni
UuHGDBNzbFgD0RqkIe5OGRj14ZZw3k1/eN5uWkhv+/fzKRQFbn9RRcpCS4bJce8xk8b7QlNS7SFz
0cvItg4t6c1pwNFKhZmnKZG+XpI+UoNgG/fXAEzlwtmb9I/dVKPPoCrhvp9U4leP5L/tm6/6SLvj
pMwQFRZXnzMwSRNS9UcV7pGIYCiXuzgjiHeVoyJ5mQ2UWg37GJFHR2j6wrWEx7VvpmHYCCf5VMeY
bGcHOiSRMO1FUkNuiX9djTb4Fx4Jn+WWMu80UqO0W+Zns3blQhvv9oaM/qhwBd/aTbh/bphbfX3F
a/SeJDuQ4X4ow62JEMaGD9WXm/aEbW1MbY0CEu3nIjQp5yfhKskC8NEgKK5583Ip0AGRrE2kauvz
IvUSNMDSj63K+0/jQRKB1GghVhUmBMV9LAtDAbYwtZYkQigil0G1jd1meaHEIKOq/8tWRU8cuJrS
9ohsA73DG9Oow3nsQFy17Cpyntphdc7cjj8MERiRoZOnTo44ulsQtQT3K1LK6U1c0n37EOBeOq7W
HhQA3mcFgzrCJiDrMTbuomuF8Ifql1mVpzxq8tzhkkqpMMoaFDsf5Qdl6bGD0rCxdCXuJj9jqmS2
8NsdsTkey/3hyUtFYTnYJ00WU/ps10RbBjQcZsBn9eEW85cJj9QkYHcigR5VBszKyoK+ERiG3LQJ
YfwamJp6LR3Sbm2G0pqkaq8RKNeLXsSRTwx703OMH+vGJpTMx/glCg+SN+RGQzFhK57vQY88f7P7
6Tx6JF8oanBYdOa42Pan8NAtOdbSwxDiSilAv6ctLo7eyXAWoyxRpGC660HL+dqI5SSeyW7pHymX
GVK0MTEd+Wl6L/BZxUb4ZYuHBVdeIQ1jinvZtTcHnjdHA/1BQlk+4t5YXdjzyvMpRdybXWi8TnO7
pEwu1UqYO6zzyibmW0lh1BmzgRLS1eOAHujV5mtGowa1sxv4gWuXjvnXaZtvfG8Ez0I5W8WWtkiD
XMUY+pFOKxD3LaL04V9KxztXGRr7W34jh8yUydZeCmZUL4nWBghHdcGLfgLr0a22v0lRfvHgCK87
9Lb+kndwugA6lEQxoFRloOwSIGOibAB+Q5hK10s54CiRtpi1kTNlgrtMbDU2A6OERRdeAkWlO7fF
22PbXFStvJeDDS383Jy/8ltddLGPfCrwX/FE5cj4/MPIgE73WGxExcBzwPCwpiqBUw38sq/MN9kk
PaMocJYV2ImazGWVWIts7xVgoFZQAKAxJUB2396EKkylTLmjodwHUPMIO0vboFvGhuzLycv+CKyG
h6JrEMo+zZZsiWpi6Kup6Z/y2SFr7ThC4D5mGH1yzN2nw7kSpj+luXxeuLq/JNM5Hwz+/1qrTkiM
Jvcf+ALHJRJHOPKW3y86qFW5wYKZumsE/gxIeLxhwWV5jkqQNBEdavu0KxsSv09qwK+0HyR8LkH8
AMzD9K3GIwufL1uVCp4WsiMQejJvraqL8d83EgpFCTEbBcZRF9TjSGJSDkUO7OaDly2u+HLPwLoX
ntCbhBn7qikxKEMDsfsdCG1U5wySJFfWiiiCmMEUaioruZJT53UCAB258Jaqn2yMcGFAKPUlmIdY
YcpLCBUoBYADKoZlVVnou2ZsXmordwhTBKhAy4XD9a/UlPrZx1VBzYof6ngLKVFUQ3l6YCrtM/gG
N1Gh57c7Yz8Uc4ZfS19CVRO2ilfVoajILEBaUEnI1xqcJcGfxD1I3kJSVBW4W5PXHsSoakcPjc+M
U+p8g5mHRrzjgHPoAGDWxfAIDt27KfeQu0ryplL3coR/oXNeVGfpAcPM3Dk0FBFHLuPsffMuPAEh
Ng/aD9wzkyfZjVc5lWYOSCoVPMcCoISMXA/WMTSrJ0T3nGUadDqleJxDRqhcFdR1XszGtJhPLqO7
knbsQBvemn6Cj4t0up9/ydIBH7D69VRpBnqDJ9tGNBEvulD2xuLElbCzInkZ5TC0jMnfDAz9g3iH
emWyGCTGuwx9/Kx8gNNaKhJtw1SQ+kgaxCPpBPBawImqHkH8mlZN6OlXO/85UvFKfMIoUXnSy0dL
JTdUuLvpw4ZDn2UPTzyKroVjwdcVTaSOcwx/tnh8kPLtqWtANy0UGfjzdwbYxmdCqNYXqBuhyc/w
oUL/Z2SMxbk4rAgC+ibwQ8W9ohY8DM1TNeUDPaHK0681iHQ9Eb6IgyjqB0q1YT4gXnfcTiYWvmy7
upCq0x7cofjEbZ1bAwzEJpA+gGS/N47PEUcFLPmK3sq3vSv71elpdbTnDyR4vNu+PUNgpPr2/4Ql
0MGBdPtPs6yxPqYu2DEb03D/lEEYSZCRo33o99xTk6embzyOeGe4NMc8E6bwbBOOjoq3ZDHCF6Nt
dkGbX7TNzuhmY/jX745OlXnPALEbXflYUqgR2Ds0lyWbOma362Qv0xBUkI6F0EgDWcdE/0/wVi3O
9P4UN96FbyweOFprGBMr4Hu3X+lDSyY409Vf+xx4rJr2B7zjNHi3ETbwz08edAkPCa+vcwfDs4Jp
YYrz4C9Z1uPDcOhdbMMczkhSz5ZuNKGhSkXnGmmH0+QqihN7XEPgBGxyZQJfJLebheYQq0yJiCq6
g1oQPEWVDWbxxeE6KcMj9k9R9m7aqR6FdeQuEBVgfCaead0+MmEo2aK5W2xInImDFNzHH07QPswF
R1uV2T3irvPlZ3SCD/VMvm8BL2vWoNeiHGvJoG40GvS/CKKJTU5Qc20hfLNxf3kqCVmqqK9Uq2Gp
E3+e2xzzX//CZY/2BwbOZX7PmczUmBEHJ5WXjylAJEQiKJG1r1BKWnz7UxfkMNeSpHRk7mxZCS7Z
0dBicvIiFwMX+cN9tpkyIKUf/weMv9nMKDDLLZMR9/7yy9p9mSAF85KiOVfmk2F3e9PIZxnelcjO
xaUIHJ0WwT0lRRSQ0um6pv+T5WRfLZzvYHUbCnUbFG9JLT2NJmji6Y1zyaT0bCArRLWmART5db3j
PmqZkxcHkIMBS0xDo9hM+s7WKXRofLsZKOFqgWzs6bFVxHdiD18XLhjWFl9Ed8kjP5duKwi1Yjlr
jOAdVGhdfUWlU0mcZDFOJ9dtv57tf981n4q7KwWTDEjcmk9qw8qV2nVLOgIpcqO8tA8aMUSXdQTe
GvzfXo4osEB8GQA24IaQwddr01Klm9pMx/wU8qkyhTPiCNFpDRuegEXt+vp+m9wZZzsIOgwdXK8z
t+0uLktwE0knzoij72Mv8dwCkkbHrDjN2/TMVLhW7s78062CJfLjt7sxMeAN29+8YB5uFuLmfynn
SEbRIkA4WQJwDSHyjXGa4yWFFgkwCDPyG8lYEwpxeT5synIvu+JGTr+8GjwUaPD/AMz+7mBmUiHA
2t+7USAugPmx/7Ol6W3N3PHtotWJfkbJYqgOl5/qGrcA0zSzw1xnNk5CepuwjEh1pOLoKICmgxoY
CZ2z/g7ZpgVa96nrZ5RaK3Trlouotz3//P4b8uOS573Ve2X5uvsx8ePkRmgylwQaIm0/A450Kk/i
zxoplUqhRIpDpkhjEl27IbStOc32vG2ymkD8s4OMZLbABFB4oNS8NyKP8N+wmwEgCJXkp4qtj2zt
YuO7qjPX4V9i5k19kdPktViT1mSYFdrcYDRyiufuw5hldrqWdNqAdON7CiwHWnLv531grzVinXaJ
UkqLROjpcOha97QTr05nevt5N6BzUua7jzNAx+br0M1yN/O9PGShK++d9qWWJ2kvOpVTm/SMqKiV
KTatqzk7dBqMQuS8SPAUHCnCvXPKgXb1kckyE3KNbh+x1OW4P1FUBw0IRQmwjOVUm+mJFVVQDNO3
/1bT47OV84zxMhJPSQnU5pj8b6m9r1ykpY12LFKAtuV5aFeruhnOXwE9/0EN4ZH6I44N1HshYIrx
LmJNSX4HhKSOFJy0FJ0oS6ZmKnSQXK9/gNJQNOZkDb/6L4mEGRrTUo335WAO+zjDF5EoccIfw55+
Ga89u7DzQIMB2z/Hjofszww13+BtoqY3nwLomuwaXQ6Y+pr18a5Si32gowTrbKL9ZW/WI2hUoTfw
gQWarGbV1LCxO+sf/LtP/ORBxXKDAZjcN5e6eEG58xVR4IDwPGcLYks7VFfpixXVmynaCkZtKqCf
8nBp+1LFGuPlRvgxeBZEQC3rMZwnsZvPJk08+mtuze9mHEtTt+2fvQAeFaGpQs0wtkXt90Z9g5r5
4Mx/+P3fS9u+mRBVmfmyna3QLDAuLlkGE/Jjs3lm315U0lJtmxutVEx9//ccp1KY90YO9Dr9Mbbj
/PVF5HsL5AdETT2JHD/kY5bHLWcyD9ATxq0YafgCF+Ux3JMA+C/vibtUYxPlq5nRklCUa8VWF/Fz
vu2tWfUj9WQcQtOBvY0dHnolrUmfwq0OPxPPfNUXcp7vW4q557faIZnSV+ZaCKm3EoU3Zd8Cd7Jo
w15lRfRDZtam+IljYNDoGbAIEmy1zYegUpsxHhf+aZIHdVbM4PKgCtKekkE+etBoWeADfqbyOuE/
DsJkQIyBwfbuONwHPAcqHG1n/Vff/LDbq0hZgwb0amjPcIU3HO8JGWYVB1pjlebZ9VMRfH+Djap9
YGKJ+zuXAGo5DdCAkZlr6B0sK+1GKaKQ9x2kD5BciMk+3tEtz4XpZ4jA2oEP4lNXTdPct7wxihzR
CvfUXMGn/XxURT9kraal05N1zIH61dNamVLhPoewBTV8FuzFQKCXG4QrCmO5yZuwr/2AEAMKsOEi
Fuq5GbjDVGGZjxl2UGgqVesPGhxa3JWsyvUYZ+1wyyBF94E+hiNDGgueSb8MG78jJ9i/8XGXL1eR
raSctiuHGbBQXGlJLbhHokbkyFXFs8UtBAxNsw3gtuz/d3vXMjyc0YWP6t4hr81Y4E/c3UoMVlDD
JKOzv4T4DSoE53lmDRQ9W60dqaW4byHuyxDbVvQVWAPhkya6Z1K7PvWFuzE+PTQWDnJKZR81PIOY
Mq+aSEmlCLRZyb/GQEe7H31sZYLZosAWfAxtAhpSLOu6tSgK2wH2+V46kRfyiOySlsH3cEjCsmZc
Fv4a0UH/7qf49b/1+z9p6cgoLzSYaP4Du1pbcJRaXPRkXBs1E+18rmlcAysjC8yRiY15vzqZ+PJY
GwFtqKB4qVA+ZzYcEpp0hQceF2O8RPcFu9+PZ9G8giFWu2REDkkyCrJdD02YGnRsWajx+pvgdyxB
naqiYrqNF20Gl+ia5DRWba3mgqWnqgkNzWf5l0DQMezTAud/t12pKmB/4fu8pvy4q1+Qn7KKl98e
80V8+8Coer1cgDmM7aHv9ky7rFZ2L4Yb/TQPNBDBI8wPzxz8I7Ym6pKxgdv7Ahjxk0tYKIStYhwB
LgqIpO0ZYLzeZDXVWjfMG2elvYnlh+LN6243xVibt2UaLgg+27aHL5ICNaCSqHv/wtHSNneZCeCT
rH+PtiV6SubVrbuffBVw/I8KiGT9ZtidaJJIIZO03S666f6jMClYzR1+j29B96oqlCOwqkXOy0Ut
Oi4Q2rVvVPi4QmzEljbpjeqOrcLapnWVqdKew5G/ZsAC6AzNJVoWcY13LCXbaH2Dju6KjFY4Ax+h
lgfCpn8G8FV9TFvh2WCFHRGghn4TSIf/n+dkOFcsFgTXXk1GZqgdiqS9XMCGgiwV0YhvgVChqBKR
byDU7QuC2gYCgQ9M2v6nYkzrhPYzD65vVxWg59fDNV4tMQsAx023BEXP2Xinp5kFmB74jI5OuGCx
8/xGNXnUf72xx9izuiq7mRKXVK5plFLyVwuXlai/z68JEmXi0mrZmoKeVzqAIf6WPA2GKtKJgqiu
Xdz/5IxPlOvH4n0R76/xPfpAPJQK6mTo9WfFi6RfuJ+MpEjc2khXOiwdcxG1DzJHkYkaYP7hqMr0
gOeiAEJy+FIXydWyPQsysxQNlf3saXUXrYX/xKSZF2qU3OcHvsaqPEoQ1rnk9LsoC2lpskIytx3H
Xz2k2IKwf1Js1tmqtBCPrzH9VbHffXaxQ9TNmYA+yCHfzd49A4lxlcSCbYe/mvCW97yHt3rsKMTi
UxCzinWUy1xM86S0/vCXn4UIjAL3jQ0p92KmtrjjoLcB1dAx+pbm+sIqFN3oL+BFITABve9i1dUV
R77JpmMgqnQg2uaVQO8MwYcprZ+uPaZ7MwvmqCWvRun+jNgo2FoPprU694OORy+mt1jky8FWFkQl
I5jRXsut8V2l8ehuCJE5HKzNaQNB9EQljs3YvwuEcwvtoFGqXr2ttuZotY//KdexIu0xX4frRNlw
wHeihiFw+NuKCH3owtivScyXPIhv5EDA4xwibRmKopwet64JU9ADtj6KqtvDKjgNGSv0SUCUZ+Lp
N0PFXc6Uro/Jo4iY7xuz7FWrREsyGVhhPXsA/3rlCOQSjdlg8LRza+wuPFMK+tmknTJJnLfpHgx+
817DraeTLlHY1j3iZ+nqp6fh65omeMWSZ0S11CgMZsx40XcyEJDzljDSXofXpGxMjWFG8Vm1Mb/r
2W7c67iVh39Yxr2euc+9d4rjf54bnlhx/MzbIWpAQaA4a1ZFn9bprIIyJc/AwyzepU/Jq3dLZ1Cd
IrUqtxF3Rs42bHlPSEX/n23ZSeNCLOKOnL9j5Li3zrXwbz2+iIEa/LEELN9L7flnKDXn0hrojFCj
CgFGLsUt+3IY2hQuMPt6gFgQy7m6MQt+fm5X+oWo2MxhEynTaSW1V0uTR51EgK9ZXgd6h3sNIzi4
MZecoGWd4mNFNmpUFeGxOUJwmOo43l1SaddKst5EzxnaQAqlR5Iqs6Y3vH9NE+L6hk2BoYBBQfSy
863C/1tct6otJPrhtrEawbCW5ln6voYSfubeTLEHoyFDmW55CP85BS0PrP9/DIv2Q9wrRTtSRNvY
ZGrqe4Y2777lNF3S0oeHSuMZlEGfkwCaq0Gm4vY46N6M/lytUxVqLR8NIVZ6ZN6IxPVNYVUecRgo
fHyTgf4t7/T5xWhOMohlOCgtLARqhFyngyJqzxOFR+qhy+R5a01y3I1DObNfl24MdBksX5W6CEXb
twbWd8JGOrhaKbE5hM09+O7QMdc2gY+KnwDbd77XEByO8+6pH0lCtmJ7JEhuc8TQJWDrgv9e/22J
d4aadbu7kum4Al+p3Rl78MScqZYyAllU0tZ/7gitMAXlMNIFzKqatFjTjE8ZZZkkmMhsgYGE5am/
uEmtVF0+pBajHepDy4+/czcAhljpXin6XI+/28oQKqkPB5UoLBlkx6jejIZy1NV2Uk8DsOTwAOKB
8vmE4gAKKZ+8NSkQzSlnFbLua4R7A8tU3x+Q2irAEXeCl62nPVqTnOVNZ55bxtpg604OvLqWOZXX
XQiT4mAVJbC5ZYnRZOeh+6GMRJepnIZw7fDdRxKgMMfW+xwkiwDruFQPXEQOJSu5EhWslOgPpgg0
GFgsfoYHKiRrXoOVy1uvK2h/oBloxxNGRedYdrhSCg3/CJZFV1RxtmgauvS+z8agtXmMFwSUlDJr
F80Qw4NiCRTihGxx1sgZ4ws1YQpUulgjsLrGIvb3NplekDPjFjnyQUzA/qVHRDX9z1/vTvOWLIUb
R8C7tEucUgJ8n0e7xB0ImUSuc6WYXOxl7OwLuf6ilc/zcIk3XGJmU5ZYD05b3XXHid2/ffmAkQbI
As2DHJ1iS9Mza8EVHkL7Z5mTzB0W8AwjfG+ojgjM5cmwg3Y9q1sVjcG/KBwQpXIphvo1oRvmRiEt
pN8L9LjPr2ZcKYCRO0UPKC+GCdGdBTzv0CsOqFFCJ2KlElvlD4Znk37dCmGH0ciDkZ4jpte0HqQN
NVa6HSRTXhm3vkqLZRYEmdo1TynofWWskhj3Zsrr6gazeRru7gj24eHoPjnlJ2kNEQS2OEGYF8oP
kNqa/kyHsAqQAuQ5BiNR2dudktrMDEn0lcD10tsIaDUaliUhbovT3/RVd7qihc9eMf3JkGYO1EiN
y0pqeWP26aPisI+KIN1izlu7hKLrAepX7j1OS9y9wfZTF/vINDN0noxxc7lMUj0pl71iLiy22Mq/
Mgly6bZf57TpieZhUTYxDyr+ba+TtpS8I5Vyxfni6RbKfS5EB8jJ/t/+mc89AJmA4JWZnRb/jVQ+
kJ71OJO4HwD8DIHbSieEH48RLtr65Wh0lGL2xTbbfFHMIjR369G1uIXmCZSnHH0eqq7H1e9/x5qJ
WKrJBVVISMb9tQ+bP6Z0WjbPCFnIAQgsJSex3q7CG9nMU7Q/cFHGmAlh6ILD7I+oDSZr0VLwP61Q
E70UWD0yX7SCPDhFa04X9RDZTW5ETOz6Kx75ULob2wOkKjpE4SHAToV3UyBUCCaR7VrGPggKYRhW
zQxRdR7SDmihoFqZij1KNCHylK6aPQ1qr1fqrWUPrUb2zakrbjIg1A0Jrqh8JQMJ7TtSX1C7uicg
yA2oEleYH/C0Jacf3lK4mt8c6+7RZt2w1IobXe8Oc8ibDLDzEmYxq031V4k33KuTWuHOplf/ZN+c
SuPAQqK9Zc1ag+Dx6aBMUxfig1oM3zlaD2RewPg/quWjMrUEosD/fXLDoavCDP9zVRYZ/WjR99JA
jwpnKxMFJUwkGrmplGo+mkr+TVoHJ24gZQF7MKxmYKzd/ggNZ+7LqWAPXBiyFT/DQ5Jxn2gVfIln
lQ/l6ZX1+nbP+VFabq0mkXTKsYhslvIC3qKH+9ktuClpXO6kpG11q53iMy3rBV9d+Yl4QzYna8pG
Cr8XEtuqv1iMX8nujLnjSTZkwLskCVVBDR5RD5uqJ4nhRy7weeztuSFtAiyTs1Ug9WtG6V45DuJf
fYH3EqBC6tLb1Pr27N5GHGABjhUJXkvsVANNFVAjrNbti+k81doPyo7KmzdaBS+LXhMx7lPHxwCr
Loz3MwdSO8YsODmKPqUvt/0LbhuVv+wHJD0lViEfshzfbb/VYZSjjHXznDe134DnYkcOvxUi8DMb
qPicLMDDJkl2mdhGU5AIqznw9r/rgM9LkOIcJhUU8/D2HZeAeYiPduc1pR2l2has4X6VpKD4/sUi
myqRw+4WQHjmsZlLmXrFec0KsD8zroOtih4KX4TKcp63mJFf71PuHrH2stQWLkpIDoeDIIaJb/Dg
2A5ed/veb5m4YjAHwWCLnmnxERpp1m6msfcpdHbusYopwlTJy1NUNM7uA1tRdXbUjz3TY/rn+Pfm
YMdMlrSTSK7w9qDo07wy9RBFJArXKHRLEVEJQUu/raZeZd6kmZRsVpnyrfl1LgjZUCeukHRjt1Ru
3wNvVy02JEc2o3Fgb6UKLmTEjfzCrXq3XQAmlpbZJas2ztJIh6L65AeZWbule8XcLZQHopA4iLcW
CCyR6zNd4e/NgpmwjFGipb8w7CvdP4xxrKXF6SoUHFHdwfUYzFeTvPzBUqoxEcrORLXqKqxVFPzS
sUHvhIb2OqgLW3A3v+7YkwhD2pVOXFWb7mEAYCkpeyblKRdQsWHRPJnxBBkvMuzJ27Tybw/0Zvbm
dizIM27a5cgAi+vC4wmst38ZcCbGpbqUQotKeMKDvGRl6Vj7WrOTHkQhZtl4OSBZBRT1P+WItLgt
P+XnKKlhV2lRYu0GnqfsVX7u0A2ulG7jcfhuIGQ1rz5fysFC5iXV+dGE6iPmeWU5NxLAt2qfAT69
2w7rDAA/aGMOtrjaUOoGwqLwRDnARca4U7+5jFWB9/z5M9UaLE/IUKh6lDxDG1cJbOfzRUrTzxSX
t3iVeKC0qJEGDwYpVmlpPy58eEsakTVPmq//Jt5pRICvaqmvZKa2t/BuuGK1LHypnVZkkTHZfFD6
lCCRBaWdKYV3POzs2lrDjE60vGWpOoOL8BIqN9tpIZqQIIKnSeYz+b8zVGcsSewSlUVj4Trf4a3H
12ZsjladPvmDrbrACeWjYCj/0tIzhM1LYlXBbSIyoT4iFZ9dLbdHKTkFSyo/hTot9QVyQYbFNkXQ
9gFzNDtUqwY4IwnQHGdMI7Pmc0UMgVDhHfspc60+PRTa3qCo5TWyOgRz8xUuiffTYncwB3vOtg00
mdA6nqaU6S5BceT77eCZmqLEAP9hg2dl3pte7EB4XLDFA2zxfeUnm2jaIISCFqVh18vH6taIIPLr
MLa7gkNzNYtVd05Djo6mlO+3pDpFJF19YzCPVtY0d3zLs4SH3QTselLuK3j95C62D19hgy+KzXsF
tBB50gUasYp+MgtBIeTzy8+41doAeXgkNpYrjJy2WNiFr1xHI0U1RFR5/EEuDuZPXJa0fdRNlcL2
F6tNN33TPikA7SxJ4Y3XwPYPRBunk9+bJNWBeyJkAS+Xo7N7iX1PNErUfTnmjw293JDdeXaklwXL
EXC52Oachv3+ufDR2MZ46Qj/ojmYtEvcI4ewhFzgqBNHLv9fwrVNmRJj0qRlhXK4pZNMKPlWfjit
aYJWPj/MPLJSnlsdHXLy8IaQykgwwWkZRAQxYQYiVB0tEvQFMCV0EnDA7nzQSsD47YmJ4PQ+ic7L
iYCFNVZ0AKamOCI2BdfcuHJJum//XV5zQvMM8tLB2m1Rpc54e3jP4LU17PTlJ+9n2OHJFkGroLSp
8q/arCvsM5i88/clNxI/oRdaHhg2jwJft9pjd6rj5IJbhj8rljwg8BoJMFplMiERTUf37My/svUH
XLHTs6kqwewObQ6asK2feJLcmkAENHNEEbrgJIb2W/yyH0o8MNTTS082q6R0LQH/sb1n2mdRil/n
pEwx9LhNpj9UDqp0ELCmdKQesfCED4oXi2SqFKJG6RMSVO+WAndO1jzQ/3b3E4VoEipK6pZUySFo
EUTcpglgS8ltDbGGsklKEPdKcSyfeZakvtZI2GDCywjvIU/MwWc3LBEVvoLW03tJbEmdjXGeQF3r
5xs6m1gOfBWCeEVUkYdQOWgQBVraZIizZLAsa7lWKm/pv3hqAJCNUQMpqsprcA3uscEmGZdj3fKZ
TVhHEeA3WJ7Lw+lVz5sGdeoGcaJrR00msmnEvcixETC7mEaiuriSy3betkWolOlR642rcz2HJUkl
fW0YDEwN1/svgAGVI2DRdWlbBSmCgcYv8yGxMWdbImo/jxxOKzkhTnB20iH/oIzPVcFmLF0tmASZ
wSZd+Y4bGDNDYseiiS3kRQhlhBp/kkhQ4y6pGXNCaVismjige9lZNmm/BsL7jsKkVzBs0eg5GkFx
iVNSNVgJ9OUXkK/5UrwWISntxebkziMf7TFdE1UnwDUznDFwrsBHobyDrPiCHr5mAp3591+SPymx
AfkOb9ReLZ/HJfE8HEPlXHp4wCdq5LugMz1OpYyvR7PUEitIK9Epr/Ax7Us0IomQXwHJZvd1FaS9
CqJ3kbtu6f21hgsF9DGAPlZ68EyjPMvtZLLZgS283BKf6v8aaFc70n4xyxHhKMa6zdk+iPHVsI6j
TW3YKQ5Qk04hlLm8HmLmdnzOOJdwgEsIXZbs5nyRFXCDfbLx5+XgG413vJq11lfDxI+ovKwkgQVd
i+uPrvMe5qAzJQzdWfWKQBQVHKlKfLN3T6hCCIZEKYrL7/Kzc7ToDEO/Z/hSjcRB4IS0ZsH1FKRj
NAkOF3LXlfUWtDvmv6cTDP49Vmx1LqCvpAJ3wPBm0eY3WHR4cXZiY8bPHM7cxEU/nbGJUi7UYgS9
YF+kp7/BpL1XJEYbDckTjzcRBrQPX7iaJoOrkmL/kGmdfszKrlfkCmrhpVY199ufuqSQa+RnFLAp
h7IDhI2zINjMJ2tL9oHH6+ij1Xd+RyVRShhPXqlu69t2MhwqFKnYe4AVvlya1IF6fniYTx9JKn73
kvd/rJh9I6QKNgAONca58UW71ZEUnNJpz7+40T+vcZCdUrSzWnhR7rY5zKR1tePpBRSUPHjALaEr
bj+jKsrUZk+RRH8YISMM0b4n1GrLu6233bHgGZxRR78Yy7He7UeLenetVxCvVK+ltKOA2RUKK20j
wVkd95UaWzPYJuTsSna0xSLEcgDdNPhf0mL/CZjR9/k34i5gc57SnB4LJ+Gm4miA+UV2xxko3K9L
SFtgjUefc9NGrt0qXjGq4a3iZBHLK4a1z8N32X3tP3hmcU02ca8heOS9xxkRCoXc2CN5Y0ye2kBg
mbN/PwP4NA+anoJ0iiTnRIWpr/62/VzDkaI/uFyFlPyT6Tlu5ThfYl0BAwrY/2scV4NPWObp4kd7
pNuFvDiIGOwLnGepyyWxIuvxNVMez/Pu+FFwFGLpFvCLtm745F3MuYNfWhZkFzq0NM8T2J+NZRDf
2UGVVWBIhfHCHic0zawB0CP9RyD8wtJVa8yy5IM85LRXU1s3JNvqsi6qVcFclbhQ4SUOrmYygy+F
le3jupqLDoijspSluX19pGqg06gydsSo66ksHahQ3M8Gt3T9mSzQIzUMtgRFN37TUFOve/9GmZnF
kePPtIT76PXabWQIFM1iYbML3UeCWeeN5DElV4+47G1FkM/n8NUrfl8FtHTK9+TqZDYfiHsVh6SB
IzWQUAW99gLKtMfeMYDhr5nLzhv3QEGVFOwq1Np5CsYGH2PhghufhWTo2Ff2befLzPnNlRxwU3hi
/PNcumUYalFNyCgptV0OofuPQWmhWRC8BqmfeOh1ZyvnILKD5fJxWinPR7BnG4jdyJJClfL+uWOF
5b7Tp+4Cb+A/bbx5uj2uKTanTGRB1qDmUWcp8+n/l+JWragRhkQQNyJJbjNJFxdebjRb3hg7egJm
/op45FD9rjn4y9sanrKiWItUvPoe+seBYlfYhgX+8QM/b0KikCBT1ibqhU5fks9Wb3CLH5NJlS0N
Kh1Ia0/R8a11/R2aV1FcmdAONx4LXQNQUgDdRPh5iwctnxHiU7hSOczhlDJsQfcITvE0z+t3P7m9
kaE7b8gp2if1UgoRHDZqcGuprACHgt6jaoibrw2O83A+Z2Jz5X0RZxrwQ+yKDF3HWs5iMlgsfjvT
mzGfXXOCrEcPTKgWAMuTNrL2OsNrxEASMN+SUvosJUPakBceXssSlx5w9NqAFZZuDF86TSqaOtWT
AewtajIYE31c+1C4HFo407FCQaGv6LtBbiycEqIt2j65SlzaH8zgiRAWT5e6hYfa2+zL5NTBExuj
k9jmrTn6U2YK/qY7/4ltXKekvRwUbucSWOVxI/FaaypgSgXWj9jD9IvfJuS4KxHjH9TV8AUPFPbq
qXaYeIiXGGcxOune5RrinZQj1Pd/TrvDR5p9QYQ/KxxAFW2Xpyg3UMIOTgu4zSLo8tmaNOg7YyvX
lhD+2OC5P4mGwLGV0bGlTOS74oalRe+rQam2H3PbkNtgTdulxCKmZNd99VkUmfTJKToFAHMPffo4
UChq1L6yLVEA02NXcZgOu8xS23xxsGhemXX4w00bgJ9mtJPXkWm91DHA5TEYwfEE4BRP5BfJ0nx3
nwLsNoC4SXO3IxRs7rG3Bp62rmDDyR09f5HC2ZRNN77f5AWPA1yXSRlgttsW6f8DMxRkskSpnHjr
CRmhvWA5cDUtPJDcImEbpwgzaWNQcrq5K51h0uvFYqoXUh7qToMV/YGy2P1tSviAxaZjD4DWWwS3
hJq4mlbVuSV0HXfg7kSy1ihtU0w8GyWYlKsYGfZpF0PRQY2JQLD9RVg+Gm8TrcdWRCGcYiVGBo9s
LtuUcJTMJnLjkjLnfuriMuNrXbJ4blbjwGSz+jWw3NEvBG+yGvsdrRaT2C7feRvBZEzrB4qHtcva
GWBD4tz1yLw5YwxoImGgFmbPtyDEoDQJGUZ9bMiO/B14QN33gkBWlLrGicKdqUps2GHux+2mUve1
BvoXq9V1oZB3HYUUFzeT+gQWvKTLrio5WCuO9ssZYgOcWSe+nUF0hlCISisrPSSzGNdt+VLdtTkW
ckyhM9MbZmij4I785cG2uY4xow6xvqxV9/WNKG5KvoHqKyfHkYaV9y0nArMac25t9+i8zy1Wy4dh
mSMlgb+1wI28On3xTuoJ9TZtT6FZQwlcZje3iW2zOJQBJMlzlZpFV0xZjGO0dWnIr1695NHzvH27
isnKYqFxqn/AOQe6zGSaixnVxNBZPB5u9R7veCx2y+NmYVAJuMlkBlLAGZY+nuvW1mOnnQe9tZNZ
KSK60D/nZYfVr1ZqZ7SUTz/bIkcdHPR36oh5jZeH8mjTR47VwLuYZUGckdoBsf7lbzs9Inn8FlKr
1n+s+vmf2BbqhdV/qp7rHaiN4Ignipn2gKjI7YTcR/h+LQGCVe7fD0ZWizks3qE6y4plESVTNq+O
r1AFGeBkFUksEmwcmxyWISl3aPJafKrsgPByLn7wK+n7uGX3CtdXOc3xdavhSQ2ar4cwaAOT3JMD
IYaDvrkw6gMB1flnM9amgVVQJCx3OR8cFZIS1mMaJjKaH9g/B32wVEFJniFnlEW1kuLkwpTXfEMQ
bSyezIX9d/84xWTu139fjhoHRnVOJdIthNqxNvs28UTlU9f3+1qAS715uCK5OOYHn3eXt5t7balN
wnfCbX8O+CV76FxcQM0ocNKbpdnzsKPRDDDxKbxEWOvQlcTHDJGWH1JEO6f0mDdJr0alRsfEMBpF
gQ85+8AYrYNbmy5JrtndrVc+wgAok4kbRaHR3ajPuCK1ysP2yN5COtumLFqvi6ek9QIGjXl46tLd
Ry2gWJJ5CbWLSczlpvNcRSDCmd/SdjDODEX8vdhGakUqXGy46T4Ri6jmxQaGLBowR+HzIW7F7/vp
NgEMSqAozQ+QhJxOTRwO1EY3QzfgdVWTvGLGp94Gz8M84OtZIGPWWoxke1shvNQKbokBnL7tQhR2
6nwp0XYeDb81y4fuxFfGQe/gF8iO64xBggjDKGExwjDsyBP213d8Wj/6WspFpc9EmQ2nf9wsF9TH
LFfHCeFGILzjEO82l29T1R6zRCbIgfW8VwXRM4E/wVtf+HwMhEWwL1FeD4WH2svwm4Xb211M3/ct
k8hEja8hguPITAktCvQkdUkPjLvjVZYbpyFRhjdlt7WQB9q6Mw2xuzrQxWQEHc2ZY0LdygpRoEee
LRog7nnGMRnwnN5u9suRR75C6QY+h/br6KbRWAMknVvu9JScbc0ipVKOBZHQTtUwTrAu3+CMbOIx
NDP60c7o7NORMUDL1BvLCPzHVx5h/rPSk//uXoQO7MXKci+hT7lntjhBd4mCVdpT2NQWzQuH5wev
DjtmuCiiKe1oeF+7QrPKT5z3wfn0lIH39i06lAghLL4e5WNvJqwCYjAWION7HsMylmK0ZMXtzNwu
eVxsJXgomcgeytZKINTON5kmq1KjyZeHyA5yqfrV4NV1Cb0i1J844fpFtjIO6HAfLSqv7waM8DaS
nGv43kmDy+5tCUMRYRnnCs9nyseSsMJsfQ6l6TBWDFD3SX5OLvWGOa6kZ0WgheGf7plf0BpaIBoR
o1SQwIyuKzDtoGdF06T/esqrt1ceDX77t61L4AgbkFyA305skjooihL/iBWlvv1R6Ue1WW+Ws9QP
d6eEZKr+E4vDkQPq2pJjLCHqvQKMf0SXZJN9l0TT1Dp3VvaEDzJwBl5KMY9BvqtaeT8mdBfdqLii
CZRFwjNzz00hepKWQTm7eLd4q9hy2hVyAfH5+R/X1RHiXxpZc6FdW2HzqTb3f5ypV+W3TkvLU+SV
dC6QT1owtU2PcuDyakRu1VXQOvGRowCWe5oc/Bni6cXyRldUnaWNuEub4916Hz41s4Wne22Kfn9u
KmGnbr/FsngdOTyKh/2ruaTjANZnWG7OJuS2BbWeWoxNuncrYapYq2M7iet0rfdG6IQzaXLmgdzG
q+TnYf/i9P9ty5FPub2FEZ4z0wKVSuHoFiV/oGJiv2snadv0I2QmUg/CSGdI0ohXtYyCkUH4JE8w
xr0mgOWJfDWEIxrVFQQEq7lUs06Qw2PLS80dYFyPvvUdd38Xj/oDGB5AhShlmTn1LG39ck7RidDr
yMM3Ppi74Z8+1pY9YTzCtmom5Znsmy3bKcgD2qA9zyGG2b+pDF+TNwwhRxCigq16Or6We+EETd/F
wfrNRPZ/EI55KkI0GiUpozWk/Yw4lnh6HTxo8jVb3EdEhwC5h+YV8smer3lSKNMmUFsYGI9rSU7q
hm1Se+uJ7zF05O9De4PKJzZuaGY9HFsECEkT3Jg6qC24ign9p6MKuOCbODf8XZFGXRRJSxRMAKi0
/cS1Akz+1ZbdsQX0ht9vLNZgCxf6YKNTLleZo3hgg2KlHd+UCtVgq6O+PvaWYsgUuIul9XZTJtiN
0H60wKuzsv9DBn1fb+bxS/JVJB+HNDBXa35cvkcNaotbRwMqaJ0RkqibiUuiSpyL3RZ6qgC3SCvM
xuz0b8nnC8EzuadTusPL1tabIwNskziATtJASVi0UTpcPPVwYWm4zfObEn2e2APv6a/UdkO6E1IL
G5UQM9OVL7Ak5yR+pmkERvtkQJgSLDTmWXQPXtg8ShVeiPsllA6d4U/S1iP06SaLYl5mmatnh+2t
BahBUiRdgVkOj6LqLRS1cKKm3HKK5E1aa/ScEpCbGcUQ5ZcddNDg+J9djO1ZvDqIGS2inqYKw5JE
U+7V/LtD8Tpg0KrcJ3nxCN9WkzKcAyJ/smvuWrNcpJNjHSiydUzgvBSXTx1uigfFhq4Cps7qrZ/N
usqC4eImPq87OilZo+jasSN+28AyoKG7LVL27RNN6SC4/LRhqGf4gyj8+wInVOCIdRvSz+zZ8yLa
gFsag6C9wxt/Gh4e35ScX4h0S3X3VVJq5f9IBl1DAa27kuFMu3451vAHvWMFVzayppgf7aqOlSd1
J425a2HFRPNivWRG3EAVP7QYoQ/sBgLObwkYiDR95Due2xi00vN6MycglKBTV+BtsavRalcMGJlJ
89GGdMNFLLlob1+Rt4kBuz5E9ViYG478MD6Z/Z2fRtOoAvFbgMekMz7I23XtVlYTtswh1CqPbDN/
kNpXEgE3ndNRzGN1enZPpPJdrm5AtCo7MSkRxfZQWJV3Da8dMdqBccmDaSas8VrCDkdU1zzX3Rue
NPHcDLwwpCXvK3QhHdkSZB1owkBk+k5HnP7C88tmpaXb42X5sb203Lu5ihnQEI2id048edyQxyBh
WZuU09SSrTDqPo3Bp7bL8CQeIKPhnatNjh33UBG/va/kQlGrV9xqHd11m7HKTVekQdVEHzK09TqO
UYK6RjkO3/ZiWbYhMrJKIjqmJqI5oOXYslPwGKkgYh+G7cLXXJzh/1G0FJu3A2RDdSF9kAIeDUlh
P6sYnar3CxrBOR/DyUnZBKqc2ktyXwNjkzcMCVMxrcpjIz0nwDJosEfrzjxBw8bFJUUQf5D9Fr/G
spbW0KryX1hEPE4IKJwrtldqMinBVBzVxnLFNVXJqiWt/Altd/7+pDb7NXF/fIzQEPGOnsQbzy2Q
gsD/K/EvUI6jHGQrY9pu2YwtyWqK2nr7nDjk6OfGBNLYyQAtpzoleUuoUCcrzeFK2MfJ6NMhkaYE
cjqoPkKJTCXcVCtAuxNQq+CjQyBkPjQ3zkGhX8F6UodGk8IDlNzPp97gt9QViPOD0CVxNBbwfJTe
X434yMZ3ZZprN27SiKBRzj31AbH2nq4VPQay+5mfmhbNTkznfHOLORwVhxPFY8pqFr4Mt+sNKtHo
gXXNnw+pJ3svTiwhcMwexdKaVr4NocPlX4wvKWzS7Q0XhDmt50T6TdyFU1D8rbWN4NCIzmAXce3Y
HRFiwcoCd4z9HnWTMdjrbA/t8XWfUFo9qmSfYya5TJM5TG7EMtpk36K5VB7rLS8WOD8ID9QM4O8E
cl5JivvRFLp5Z5irvHBpHrmNUY9uul+2873NP95GASfcsjh7H/XUpIFbS1x0LbFnYJ7RGwpUXCAo
6xsWfnNUJUWelgNzSkHny4fvqQB/I4yEMngxnfz90An0ilnto34oixmVuQfjoobQQ6SdJfkP8L1I
akCVjJ+oiOaKjDZ2Rk4gUKchMToxzVDCZi9mMgu/6gqdyXtbTnypvosjpBTuOZcmGFiyFKA2Cci9
2BPh+HCBk9UXkFHysBbi0dKEOyF8UKrt+ttVvu8G6cVdd6TnXNNp7I2fEVsM0V+WCtLArOFW9hPI
NyWAq/1gA5uKzYv440Rc9VdusV5q7dRuUA2+JrkqMEQ7VyR1uylO4zJ6qPdFQJI76cSO20Un4JSE
aQJ6kjl7vKaRxWTN5PaRW2vcA3I1IvIkS6V5Mbu+zJ+HA1BfqMz0P1VVDu3bOQJV+AfW5Vm9YG4F
ZKR/wtPgt/VLXpq0Jcy+BjROguhTSWTGNRKKFBpTNP/lWyJskQsl3NWbqTKK8q82tZpF5FOBqOwU
716I4VK/BeiSAwS45nKVzV7Jeo/k4N/Q9VFXUT+iqszIxN/XdkSd4gkdaqpqKnp3IQ0zt9B+7Nb2
6mIRN+LNi4kV/75w7fbZ7RocMp+Xkfop/Peotf3japES7kDvQE3qxA18PT2u51KnJk/jAklDrGuS
0DOP1vAJ+Vg7U15u5NnnEYkVgrgfA3Md/fot0s6pqhaooL22b90PIU31S1xZXzf3m+uQrVfrDUlV
8DBVHX1CdPxTAwtf4lvUsOlqivpdi+YVWfKAmsGCOCmxQIWqMsYsldTd9FIATO8opkcdVwteSK0Q
ydHvMFdhYpmY+WU0rjMM9EheH0lwO0zGQlOuPnHDBMRYMW18ZZ9a8R0LF2TAbecu6aNSH9k/Tsaw
eOBV447CKBfmymmPg0WnNajHA911HvLBVwJSjAPC/300N2Lg/U5zN7aca9Onsgwr471te6yTl994
sJDFbGfUzqQGqlDDo8orQ3z+ZfAyE0Fu79MN7Hkp/FKlCZcgeWcHnxIhWRgjFRxB4naWx8nV3Abw
gV7w3N+BXZKKSLg5faSgGl9dtlwHgeIUGZUK8w4JF3OkfYfytpBRQi1FbMoI1ZbA6XLRR+SKeN7B
73sLIOaOKRTC/F/bp5cfaHs8/Mfl0/22eP+BRpx8io/JyUPNpNCk5vUZXcQLfJNXRIEhj8VM8bOv
/s8uYDxqms6SKKCrBzSvHcHbBjoWP5YLzi3WOGs9z0o8py2f1Sw4/r7JdAuHO1Le4/G2A+2dPyI9
q0fU6wWwFgrQ2YckuwrV/Pi4gCDjFLmfAATjNcgfrpYFx93M/0X5yBtUr+N42CdJUTO4DSF/uKTX
7xTtXjHtt/SYQWtW4Tq2cwke2IQkegc6jSPp4evC70vYnTQqpWk0ERyQ0dt+ttb8AFlCi70G2OG8
jHOO/xD7BdZHqgExqiTAzvexHhSfOTBeBcYYTYEyRZ0H02lhOwWOOyBc1xXyDnxCf9j7YbkkDGM7
2gHsO1Jt7flFgMmMQBEqLIY8ca0D6D5mzLg9veCB2ClUkgBBJHFhfYEf1HhHSt3MjxklHXuNtmls
flFrvUW50nBv/8OQegsiFGpy94SHNR1xsZwaTSwXRBzys2RwoumCuoi9ngxVIK1ft+A2B8hikFFb
btWgH4Pl8WYWN4CKpdDUiufjjE4biKXRs2WUIQ0cJBvviTGJfhi5d4nkZbkKezhO0XuuYa06/vKy
vO9kDpVWlnYnDe/96g1Sr18puWrgQtC4C7ZaMMJ05kpjwRboQX0wp69UyLJV5yg4kE8CNcGkyMZ1
kbxF2AfVjidbkQ/QZMZmOPXrG3oqOaIIRd1eIp7c2LF9Dn66/6UMDTS7TuPJO12mI6r7TtYKdAYp
nVraAqw5lK5xdVnSuIQLXZNsvSPnaDD9umrOdjzn7RaGEeY0SGackbUXp2MhXvIqFjL0yKV9GFFn
t32A9I0OofcHd8izm8b/mZlYiya3aR8r9NNzyPyAHLYniZR0b+nk86oJcDsA5onCd48f2A86+ijN
2mZ9ICCm1SCJJmbxoAjBvCXVnOXppmp2abXheuPC3lmdH8BhDBB32aE5CUci+BvK22z/V66wW8gp
TNuJ59VMJNchyAhClnc35Vr+3IH7SA+uQ/5QX/ouBf3KGNP65nECoO11AU+O68X8MD9Ad3LFnZuU
SW4FCmnu/FcvZWhFin8ReZp0gAIv2Ela3ftPo1we+OfHcdaQqsx2oe96TgjMy/zzDqWPifwmxh3y
sxYzeQ162zR9VKiW5Xjmo+2RCGIa0jf/VQoAPZN9dclfSi+tBS4gIlDWhPJQvwGu9oCjmoFitVQQ
BjZ9roxLq08RmIFrUfQRzTxB2vcYRWhYCm5/Xhm9yCURhVbQfmcib11ZzDshu9KAnribzJqGhl3/
2MPU0+RQ5WRbijLy68h0kDkLmCA3pvvApJT0kamsSebbalsdXn9C0GuPgQk3SUY8gHCjl+h0ZvqI
B3QlCCpcXSDk3nIm20lHU/0OVuMtOEfTZvVHxh2g1pS1H6xoxt7kV6phS/ny+OUm7CSe3tRmURZF
Qu6Uoq2q/86D6MrMgIGdwMyDtxCyJgecQOhyiGLgtVy9QpfOH8OemI5fWLCS7ZUK9uDAEhaeB4J6
xGLeU0IVnWbaS+R2Ipip3q1MwpFGoAAahsygkFmnVw5o0+ROf1p1l64neDfiK6uwjUTpq2QimeGV
6zymYuqqszIOsf0aaCVg9Rdn72YonYB2DQwSGttq/4wq3Ljqtyxg2B0TufjHw5WTp/xVjQJrWdGj
BScv9mVUSZy8dAPDvhR6LfS3fMuU56NnExz7I02NHLqix5g1fqPx6pPjaepGn4obxDqRaY46SIcG
a/PApilkurFSrNIPH3og9e0BrDnmZJcT6VKxFySf2H7rWpamkqfvnxCY+ukF78z9VVLoCjqhyhx6
1CTA7bXti7edS0JuKH+t12ZHS7OFqZe7LZah1brjH0lXObw9iZj7gs7722kvQPAhidMGbCYaWkBQ
1W5a1WguEGNq2o7vgjERunMTfMwyMlYcwEq9ZrG2ZS7fGNGz3wQxyE7TwZxoenK0nMx+S9l4lQSq
SiTTZ15gfUINFNsUhFxQjN/JyJWryfhWcKTEl7bSNwcPsfL6PUGI9s0Vo8z2XWSSe9viISo8BZ5V
L409biblH7UWqiO5L36L0DZ94/goSwRcq8oiT6DokIbL+eFb/FajMay8oZpg9+imbyZ6dDtsz7Jh
SGxqR1+xfJKE0Zx8D1+iUY51z1Q6HFbyzn50q4YpMep81qiO8v5SXX4VInvE8HkEEIqy6V6iwAk7
ZxFkkIeR0TONLOIlmcub0ezfMcm0sQk+781YXANXcBnrP1Km4EZf91E1V1/eK5gChJrsmApt6ZJt
OqKEli+z3rJN5YdXdhl5NMy/Xab4W9AAF2ImcWmk7I2VQWgYUaHfT1tF9ZNaqYvRrvxhNC4s0XbO
bxIr7ev+M3YfX8SidkIYRmNBoYTwFSUHF+WFIu6eFRZ0xIFoDFwMtGO1kK5c3VevO79uA2T2D8BK
9+wJ41UryXeqQeVdY/IK/J/isXwboZOWSm7GxcGMLZQ+xisgJp2UKKzqlWEb91OiC5MU8uAr/bPc
QnpDi9wBc2hGsBu+G/euzFJW9OAOKg5eWvO6T1vOa0TlZeRhwWL76xeRUmLcU+2BsJXW2Kqrb+hX
RxQLqkJaofb3OTciwo+a0oRe4j+e7bkJKFy+xPHsZXHnV+uIMhdbWv/K838cH0SldU9xXuSAy58O
19slUeuTkTeuNgRNQHq1VgUC4PJFpSmsAg60vZ32DVbQBxpW5Ufc9xUz98ypitsi5aJ6jHwxMLYu
OSCq69mN1NxVUUDMEtLC6AJ1QD66vYYaKZLggFyrmnx/7xD6d0kGfCw2Z3RcjKYT8v3Ir1zNcQEi
QmewUL5gUNS5VZOaS9L/VUnCKBz6b+FtNqV2kc+nISqq5jYqOtdUkOHxUGO3igldTmY2cEZwFpto
WjSSbsRNlhC82JEyTkgbEoBinSPrqp0MT44g8tU4FYyeeWgHbX/MVgrn3ZTOZnmOLaRxR3Zg+Seq
mJixaBrPrq+sZpKfEZFo694QvU16Uf87YYxZphDasiiDsgsZguypXJWAZ38oyLCIgCfPpF7vjHWo
LBoSQXCyl8VIhcd9DqVgLQru05JngGiVwYSF55OOuPbGXwaWDNbl0mA6U8VqMI7rtUVz4HGB+oX/
7gb4j9qBM3S2uUWPyCg/FRJsOoLiWQFZUdKXGd+li3KZX4++U+28j6G8IssaEj5EyRl9NqNzeL85
p5lb8ZV+X/qtTjvsyXge+uVDzLk9byrItC4sl+EAata87H2uQV18VqwRWRInhMMkkY9UNqxoeY92
tynHxhkrXqC+OH4QqKYvk8o9K0RzkeSwvo0DT+SaGYVKp2rDxfT755FEiIErk5yisom2dyn9WAh7
2N7G17AOhs1A6bvR2CWNA8nDStywYrn+ys3gprBmKXWcf0avWrP9uYUIWgVurJqj533snfkO+jkt
EfH1Hg1NiOolB6P+rcRH495LH6kp//cZPEQF2UAUOAABO+SwQbCcfasvPud1BFGg61u+gF1Q3e5C
b0fQVFGU/7TWBaFK8UgfFODTa18x66Z+Cy3wQF7r6qwIKM4eg/TudHqu+msbThpd6vrICoAWsuFb
a0BRyg3UUSTm8a4t29pYlqFrWYmFAygelzOLzW6/0iPcMBtkhAxvCIFm0GAsfQlw62a9cMpnG5ev
TUR7pcPAKt1lZV0W1iHecPnZsweZP275+F7MJds4WERQFOWEHJZiUtJ0q3c/XABGMb8mTUvuJpo2
ykvf94OGBsEGmCIcwQnmArcI97ovmOmLbIjitrnyHV1CtSMGeUVLLBLumggMGgIEbZ4VNzM/ejNe
ke4H4HHtLskmuxwsv4BcdjVBTjyarWO3jutozKP6yG6XpEgpKJy7trYdiXEWXGix5d9NDx/kEw+Y
lEnbO7Zdb9CNRXfjCH4HCFgvsn9ImYwrHNEwfrx7agwKYtZR1S7+syzQ11jKInaXjOiicA+ABvPq
2zVPNBQgd6nUAYkJxh+S59woG5E2Nnd9iWsEo3STZGVwvpwYjNbFRXMJLzixPavLSnVzJFQGR8Z7
MrcYFoA8QFXeUBWEhbbly5TtM46pcIkSL+h28TT68DFIOIfeQplNUkaA5VkqrtPxHfdWi23fg6ly
lpGFE4NmaZg3BcL8T3BJyZ+THXUjvKbuhrKvLwaIZD+02MObl7iZICAz2gDaobrt3r4ZWSobmSu0
gAfDuKEIacjHctWogsKXS/53ISkb6IIiLr8vJQlITgI/LPRR3nj2DDI8H6GkGrCKCbqOCvGV6nVj
bPvwMvaizXqE5EaEOfoRmmN+CIoVt70T88eogNGrTyYPfwuvHLleJtYolYVv87UkFHkJlOXLWDYe
4Rwg7L95ayRwGf5A78MT7cUd5FlrVgeZKotBkMPmkDMYlAHEN+0OWI1lgOTLiC5ClKqX1Ij09/9m
8Gk/vtEVAzzEpLTV63dACvjqatMVdtjn5A0GH4fZqYkdlcuM05JGkNC5YgA4nhNlAP7lAphj2T9f
yT4G1kBGGeo7CuMNVL5ui5itSaxw3YYQxCXVAVHT/WYY8TAAmAxGpiskueiD+QtbVrHMaT+0Y+VW
c/TCyUh4xDEiiZEZNe28ZInNqtFHvV3an9Rt9XVCdl1yMGndL+wuYMNHphyJmnS8rv3EcWX/eLl2
WnPjylEBXYM9D9yQMkjUwjzQER4eYQ1v8oANVwWICKQyZBmRWesy04VLKrUQsBEmsyO2BU1tlH1s
U85WTJS5fqLPg7QN1s0z44+4LWE+yFd2CxWMvuWdPHb7OBxrUIzDNsINK1z6M6wR6c9ykBwSNkwV
HGm8EdJbC20x1SHZrKQd3aX6p6Y4fhHy5XOg+BVOPfajL5IiqvkLSZALIlMykWmVNRvO5ArNx2IK
ywXqf0t83+sqpKidKDLexPNQrtcAwbWGqmci8ZCLs+oaWu+RwGa0c6ODkRoMTxm8KilSldxVaJlU
7dARK/UlqgK7pPN9sJq5tHGsPTYR616SNdMUE4ewZw4YOTbwe7Exqe5Ai7M4BrkYck/3N8m2/3Ph
a/BBH66ZDwqYtJSYoF6i8uB6znoTZSMnfls8omho+y2FSg73K+TpTXNAtgm3OgeAc1CgIbGHh5HE
7hYinEdxd2y7Gd41VoLwNK0UZNXAH+AwPo1kK14la8Zz/g4KqwtIDx6GUIdE3lXeabkTxQaJ9kPd
/MZ/BaKtm6m+sNZY7vTwbd/PkDdw20xXpJFPSS6VCjQBCn3R/4V79063rTYM+IWnSkLOWIBD30IT
JsAvJcb5iwjs1zWXISTi2tXM0qcgbWeduXRUSDGRdxFu2XuW5bCyGVZm6qSNOo+NXxBvVFBFT/jm
H+JM0hOvKw5kRwh9+ws4y/DTrPPqGbpBwwGMlPCNNzqGtjk64EEn/ztwBXYH45W0nfbLTdViLhyF
qX1HvWwoLMtC3I1XXu2S1J5rVnx7PkuL6cBHNT9IsYFlhKwTeCywgDDtGg8a9GGbGR+rgQME9Xzw
cjeIXMRvb2M0DXo6PpS31npor5yVrDPqewqn5hHCNnnpkZeTGOoGtC8kmkeqIEdGgPu3BucKNbpF
IDx2XJ+0g+t67bx6tWH5FJeYPwjsmwonYEu2NXElRDUJDVqA2G3crI0686JUYJsp3REGm/MbUAr5
IEGMT5LuK7a2aI/9iC4ThapW1EpZMwj/+jvxc/fsE+ZzUEh1LNWb/VHVYcdYitiqbl3kTU9MbrfB
FnD1/K7SfpIaln58jLdg5xiHrup+qPE3EDcDbCOXNkpxl8uDCmYMJ3Y5aZHoSc30pyL3sNWHM6mo
LgRgUNMTTSkHL7ZKo6psydYZfTrWYE9/MdnFLtM5DhnGPlzKhLO2UryEAu38+5+PMQw0Zx1f9WEY
NCKYHSQKPmV0FVwdnu3DC2YQzzXDCCqnU/RZGCtSQVgAixvUrSwfGfOSNNjtBReuVr6IMCv/KJoh
vizxkVq7HkNZaaQoijnhBPG31gXAvej6kM0wCv1ZmU0PxSmHHUmTIvMjScdUHI3hCn6fkthLhmDp
CloOUHxAJbhGJ1g6ItOSgLRGszdUDHPZYbVl8yyuNsI2RK0R+dODoGRpBTKYKY927O/31M/w8gFH
89o/ILVg259FCkrF+oQSC4CItrPOalMfh1JNeg9Nz3+H5stdwP6KRme9EOmPLLFIwoUd5WfKbvB6
HLYosGd6wsqyDKHUU04wYUXzzRcYHFYXlFwYrdUs0CP9MbRFxIZFCb0valXjICEtdeOrk4/YVcYU
zNFLOjuo5f72WMRZ1x2aCicjfVcDu4IFaQFLnBk1tQl1XXoDWiwmuSwfJISm0RvZ/ouF1ksAfmXU
I0zc4IpkvRhVCRMQhBk/fg5RXEs/U8ROITlWUQEpdZCFECLlNZpJggs1NQji/O+Lb6MJcKI6ip0a
8g1BPahxE9b1eDjt49yqEHdfPuMr1jq+U8R5sxy+MqSzDVJzf3/3cpbmheZ56lH+qoXJ7az2Ca0N
uTOmqNXoLXnH+nS5OJFC7WBJKyNJZ7JcPR2E2qTNRXKNPJi8QtzieRkzY24F5Rr/uiOAPqnD4gf+
yBfdz4xL5l4+kWl9csJ4p0JU14VqKVeD5Zxjh1ceFpoHzyJxLsqV8azgth/QnblH8oc8lvEAjPzT
UsvqD+D8PLRfIIZzsqNEkmaHdiQCL9r5+NDyRJ3OhLZKMoapQZWDmCsje9DVOKY5ngiQ03406p9W
i3TbapBut+hZC5AvwW3h8bc1AhlJVd9dbi2GJ0vYIDGtEDVKfbC6TsXVUHvc1rhFvfcyTOGcmRp5
YoNiEDZsDqRqxKADsmhpyIuphN0kn5sIh0Su5HELHZfdKXYaUKddSG2xSYEgHVRqvlucCQ2CY5ip
PKa8S3nwNWCKMpDChqWJP5hOHTSbrz/0f5K/nbvgcd/Voi5SkAf2xxU6NxrTzOdvcVMjOQY8zXf+
MT8mfQcIEeGYFLKqtPa4Y7g79Uy9bverrozfTbewOZt4GeWVr4PAng1093AqVsWca/y767r8RYFE
ybdI8595Lwv2sZs2Cf3hhM57O23VvcNBZGVvfv9ZrXoxC+b4T6sD27YkrM7/f//xpAusE7fDiktl
hrpBaTR/SGAJCiRDbnsbDTpQygPjkmdGEQUcMJg0ZwS6EehrSx8zx7qQx+EZIcGdEfjMSyj3gjjX
nqMmf0E91dvnwz0aPJTQyTDDTrnPJlVA4CnJPe5r3ls8AMxZhBbMi0ucSx5+12TsS/Gz2zRnvG+h
2xJZIQKBzQeY8OwtkSLLNi3ThEGWaYMx16EC7pbvMacLzm+KLeVLyY62iZXic/feXj1ndMFW0KmU
kBsJJ+KBNzzgKhH7cXyfWO6x9ZQoXaijgQ1Srgmpub2mhHv88ZbUu/jLfvyv2YzwJOE97aJPEg4i
G0lAvWYkppcBfL3n0PDEuCncbSYqv5kc3hm7uTqw15uZDhz8ou5/iZn2XASs8XWh9nPFQTXXttRY
vZ1odOt13tmKcQ8K7yCDDTgx39oSHrYLxFg6uP5jMRvrccq1T65gIyzyeKLp5iV+cQWpCj8E2ryL
wSotKmBz6x8QhbsKoHu+QgroUB/aKm3rKX8lHQ1PgYQ+ZmefcSeQJu8nx7urm84BqoBH7torOkc9
g1HgyTNc0viqcPO8qX0xEWzWIRv3iCsUPJcEwN5abs7m1w9VGhBPNB1WZf6hTkRFKJrOmmrYCvGI
NgdFN4HbAt/XyZHreX05TfFJC6CHduA3wSr75wbgwCYVVATZbVVEJKM8AELCnpBx2BoB73LbNIs2
PYdnY4wizFpHiIF1hEgzz4t1J7wuxnA4Kb0CC/WtdK0HnGMZgA8w1igf73eQEln43hawh0mZrWpT
ltyE/W2cHxz31drJyq9WQr5+RgH2L/UxcSLLj9g6NxXmmqWrhEEks4kY1lnMKnK8sU/ZPr/m8WLh
qXkt/doM07zPA1yJWpKHcoEvdLDCtdS8Gt8b9VZGkoC0pMnmwopY/r5lNSGY9gO4G9+nXL4fS/Of
cPFbXKHV4fKj/HogSCXxLjKnWgO2CGgNpdkcfh0nl3rihR7ht/0KQYn24o45cIcf1Wjg71FYwr8l
fJv7L/whcPDsf2lg1VEkf1hS6PlaU2kusIA2ahDyPpHTHxvdtRFod0cGtskRGguujFcyZ9gUGmeN
hJ+GuWSWDON2X6bg+L6UhMD+jwfr6q9VP5qpiPsITyWdu9uiVjyScODxWNngL2UW7KzluKKATEUl
DsHQnirpwKNBmug67a9h3B15Vx2gqdih8vYgDmiwQ0JM6mVW/NhamtWRvAV2jFM+rODcWO0ByRkv
3B4aVrsNzKXcLOXw2zs2zh/XIMnvS82tH0aYJyAuKPPezZNkOONcABIhF72Jj0cIbTITtjXec4ZG
UlvcZ8mHZolXQiDzEQYleaKLlVC/XrNrfakS7zO6zAb9fVSrGDf+xiHhtLpEYW4IpAHS4/j0ygaQ
kK0MeuEGQ4vsxSnGcC19kRikqjX+yM/BRdcBJaBwxPIG99+HTVyBF/CgxoSbM7miLQqDYjEay5Ob
70JgkSAXu5LfK1Qt7uM9wXAGVJ5/0sSum8BKHt5UdNNVflwZM23z7rGKEJRXMRez0QD8f7/ETgPH
CYvlpXatEQYyN0pGM1OgcMgcTEPP/I+RPi3BmApOOooir+EDYhSPV9GCHvHqjTLrdaFYXCG3XsbI
kog6hftPynJbtMSFqjZ4zRPzqLcBAG07cwlN/b+eB5z2/2za+zMlMqnuHTWqj6wqk3nXAJ2rdtrE
1GH1xqe9Nbk/cm9R7EESztvjoT29oAQxqBsiWONlxD+Pi8B7OxNhJXvKiuuto82PE4Ls8kKkJBbB
C00wIfDuQQDSQRnelZzGvm9I36kjVfjB1e0hylVlBKBaavAdh1BAwE92J+YY0ZhP6YqNNO3e23Kz
H/6gbCEkGLo+FmJILTnwmqTMRbQdP3a8c1lb5xfFyKD1HgBuMy8pU7NPVZ5mM6545Wdix3WN+tBj
KuJjFLFa8bKNkZ7RLR8wFqrR7OVwz2bo1vKXGAIcc0rZIzS4/3dh/iSHs67kB6+fjrX1bwghvbyW
dLXnK/URMfLX0FLaiit0VLtzLOsDdeGgyQoLbJHA/XiOB4b5Lanmv6zDMMQPXePgwlOSbq5wK+zU
s705EBmbtP9L6Yt2lI5V8MbaQS0akqkuseRXLFsFCkMgx1MH5/OaQyy/eyOH1kcqrodn3THxdTZe
X+93mDnuIu5gk95fnMWKIq5Pe30lBGTkkChicIa1hwMPyztrBV145JZV2A2RgGC+qU+j/47SKqSJ
X1/VgB5IozwUVbxKODI2J7NCA3PIxPYwJClKda4IwTPcDe+G1wL8DGUiz6h2nnRAS0aKnNxHOdIn
1Op5j03cPUKMdgy6tRvh4Oi61YgzdyobzsSfTxYW0PX7ktVZF8ZjIbrp4+pxaO4JLC5/oeknksdD
mdHqmBE/YrCs+lQtWYn82r0NwPM+pPcAoVlfpbLGmFAaljjHZ+yyHlF8J4wIQN7RoUJChbNQGcYH
CeoVUC/UocNDWo+78iRXTmC46ic1CjUmpTdrN9Dv+ev4/EVaIZybG7ztnHHeP2VuDtLcnkAnaeE2
MvjBwZhDPN4LpbIp2kH6QluRKhQosghb/wjSEml17ABtQvBqUtb475y84d1eT+6uT57gfdYeqBUg
7eIekSANrKbaphr5ZW9hhB350iw8m2ePiycOgvEWnKoPkJMCrWdinKlars3qw0lvVOtCX4OxxfJ9
4OhQKS83pa0er2zhf5LFNTqV+wLMsj9r9LukReD2HeZxC7+ruu8LTHODQ0GNigewDN93AI3Jyo3r
KH5kj3+UyAp3wjoLsY3AgFqiRU2ovXnNjLseVoKYEXgGStSVJQVcSPXdRcDtlBxTMXbWOP/B9nEG
Zu6oUB9EodxLf5BUBYUJGJu05cBW1BToD9dUWe0UJWNTdPlntPpHX0gGAYZCsDnWRcf010+udOlM
+1+z5OIAKHaH/eKvfvYGTZq0RkRWTAX1GBULE1wyzlp3DtEtvSM8dVsVtbCZ6RqVM/FakI8SM8Vo
AWkVY6LSkE3SZo74kCcDKxjjUFlZRJ8FwowO+k0QuKQfFBWiHdva57gZ8tlCMQ0cBXoHVbJFqZxB
o02j/gs8DO5E9mqYiIMK9Jvvb9qLaHPz4ShMjaBEE0Km4K9jl1Y5dlJp+tXLMDUPUwscDspeOkP7
swtaFbrzYTbHcL+0Qx3gJRYy8AvjEI+lrG5w4TteK1wReX65/Py7LjGd909RARuijc6ffiutQ20Z
zMUZ4+zmd6EArbrU1qWtejDzBZGQRFCILUmG6uw0zq4kY8RFYQ6TlfL1aoc73/sev2+GCAoXU4H5
jTPKuYPf9sawvU1NGFoMDsTh4a7Di0hpIMJfHj8OuZYUmtzhuanOwbvaeQbGAC6+UwCxUKxtc5Dl
d9NzKOP6k+e3chbIiQPey0vVN3M0LH57YGMPORHHfyBpVLf6CO9kwlHLpDXZcyAqUqzxUaa/Jmrz
hTis7Smgp4Z3ctr/9+FdKBaKPCusRioOcVFrELP05RhnpG0NaKeA5E/PRhybqVSfNo3xxbBt/qhy
vU2w+HyUsZ3kOJ3GUcnAu70T5qhT4W2B6m0xtNL4Z+VOB+RvRwIS6niQZmxaImXqL1UUlYEOCDpM
ambSTbl+lfDyG3Ua3NJoeKsGquJmWrkyk4RsbGLAmku82+idIGgaf8LWctET5Ep0BfL28IMWmama
LvUVa2QpE+KoLSyx1PgtyXVNggI0cTPnMcMxp3Cjkz7naBq4h2LHk/ByfQ34Ko6LOpWnG0gJNs6y
sSX8QIKi0AMDiCioZnhV8iwdnKFpn5KWOlQdN9a8pI9LupLcstfWinuEBomLDfkRmK3LVHZobpMy
H2N4E8fTq82ZpuVdjIB6jcsgkP6s/z4xE0UWulvqTLYsDNC658SbXCArL9OcWIUViWn+lFKRDg40
M7lFOME2jiM1CTRdiAHwgZgmTHjNGf0z6osuzJqq4ANfYVgJoHV8Z6tn5smzvNBi0i7Grw+csijC
VcNxRNDZghVUhFowBJr3aP3GKJgfEFGh1KuSdgwjt3JA1ttJuH39tBLoMOSxNSS4XcEISuzP4La/
4YGi4BUAppQBaAtvJJtScbYTFJODSiqiNrcxUJdZvK7HRB2d7H7tXgMdqlf3YFlcI8YFvG2dvbOJ
0rZvSERHzIAyPOKieH7AjRKKw80pSK5/pz6lds9lrqPLDULCUxuuVnNLmqXQiwmGAGQNzDmlCN97
TmMVyOr0Fc9B6CFP6Ff5NWZi6ZXaOKMQ4TbQi72ZMPydD3cr8+e0U/9fM4J2eCwowfsoC7RDIVKI
rqZg4EsQSJhNEkyXr7N+hzEiwwUxgi6utekfwc7XGTBjodxn5UncrV/V7jJ3WoqrIwT8BLu/oCrk
ZZqC6qelRWjsKnqDXioymfl+cT7GJAyD01v2Yt++/sqsQgkx5S7cKz98TWz33oLJq1zORedh4PLa
HqkuqwzLPeq/wx4mvnhsJv3ULLZ6TAGhu4KX1ezRejizljtvdZwpRapY5+bDEZlIE1llB7tqIIL6
0XmOjmsbZ8mB7Q9FgAvNoMq6ZcQF7MaOmqHEQjM9/ggxbfu2g5my1k1p8dtVgnyO5ON4Waw1tm5B
r64hzmyTv24cHZYJems+cBX6hsq191EVWMBzCG8c1FXqitSDkUm8LBsO57kDEBFGRbOl0TT69lfE
IOGwjxOqysvtdQXSLgAoYt9feNvpYgXhXGSJK2w8ru2BRWkWLN8S/m9VwJs+m6GBa94ud93eKPh3
tJherYiuK44bDQTztle8HndygmEdE83rscGqPEpV4VH+CySsIRf4kQBqV5lGw6M0QLCxri9ObSp5
bE7ecQ51qXqcX9lHHTQi/nBaZCK/gcXoSyWQWJ15XLs9zmBbUF/f1tH8Vwszyfe53P3ia0rPR05D
oeedud9nRZfzEvlfL5KbQo+8t1mJ74LfCKCM4ONrYi4amXWhOA92gDkvwDNG5tORlN/HRRWJ7Zd3
Hj80T6QyKGBOeWX5x8+MtN0N+bqwUtoJj3X/NPcqzo+LJZw2eihXKCbVT9kCyx2GSvlpTV+F/7A/
+6/SD2uSndU03URMZkZ2SgxNhp8NB33nFRb5s8V2+SDKndexvwGVErSrbN/eNnRcxStK9QcFnRpO
IL05j0RK0yrGqjeOiJ9+Tde25OseboPTLSPy1zTS4nfcBYbMxCiFUwYzwV+FDypQoXzgUzUUfQA6
Qd1A+vIOFh5tF1jkcfJV5XtOxf3gKJou+aGrmPo1EmVrblUcgYksd7IyYkEhSLqbawXvbaPmTNYe
OGtzpuaPK0CyWXYHOwXdbA5ZaZ7WNW0YE2P4whNIDiJlPmiKlPHBRpokgNEkVOD6yJ8VL225wBSL
+dx31340cVlaP398bUZkKe/TKsGEijn15spQb1b4EEe52Wxv63qu0ftXGII7rBYBLLzPde3YOD8z
K1wFkC3VEJNmQg0AyBAnME2Smb1o0LGMG5NgLbayC6x2TmNdlbSAKoY0UCFUBb1Y9aPerocRzjU1
uoc0+zOOcpoFlRm3Wwl+tqEC0XWqpObHRKRODv5fp/4idGk/ROn4Sz9xVJqBbCU6eLzY8gGRWSOw
QS+pgrqxLpdJqEEgYKEy/xxnaWn7ucYuqeigdE9rOzEkKlOvN/Vr/ZcCPDi273yLbn8MK6MdEkuT
4cdDKhzADAq39cB+tmbR1xvYZfLGxqqQuUWW3Eo81IsYevgCM0bIPQUdt8AJhTT6qBxgq+wKGDR9
Q5iR9U8rUUuLvqkp4ma7mlhNc8gqwMYq4u+LViYzAIVmwN2b264Z4o7chy1J6pHMwM9TnL4PVYD9
dNVPJyAav0bd5n1Gm8nBooguke/FcimsClQ7sa+nbCzFEkgt/sb11LDbT8c2D0zL9qiroDUZ+2sl
+gYCjKkIPDMfwnZiRrFNy8e8F4zaHKedq81WY/Apd4lPEJDj+UgUi2fTtl9C9CAUFTrpv/9bCBdD
zw0g3vsrs5ONHN5YCHCxrLW797sYpTUTp+vblC5v6XHGKyuLJbUSsONgO5gQFPOyDG1h71rUMpyW
4aq0e7iU8bXjzRGD16DVEpsXsI4xymGZNoYmH3lVLsAq8tuTm2+r0PJCKq5PBmKjzFhQFHfgEV9M
nBs9yxmcN0ze58uOmwH2ID92GcwIu9Ur2M/JVAfc/QOXETPk5jLAmoFqRWfD79x5kw2WlsgveILJ
YGq1yz+CZj1Y08eePMsu6g9Qhilrl46j7/Mg7rXVbdXoL4pyiIt8gxJZYmITYxuhFkdU6mhxnrHZ
x+74GxR2/wIfhTGBC0ojS+f3fE9LE04J0CWvxNvm4/9plh3TDE09X7cqtwfJnH3d+UNdyK8WXMuH
/QcGQ8u33k4WqbETmWY23pHEZwCyaoNGTNj6OgLiBJ+LMfyTVhi215/7cS2Zi15nTVlYY3zcveEM
RKfIRZL2YunE0F76WbZ2CjEkuF8bUqxX1zkbjCOwrBf2mU4Pz4ACFbtIA0KYZ9AP0lxd3ZdO5PvH
POpd7b+eHmTcoJBqiL0I4L1lGGC9zQBVrMYnnL2FEsOLUMXZRHaP3K51xZywrOM0547n7xgyObOP
wo8TDWsHXeryREzhnoajbOdc7EpBLEY37mx+Mjz15b/X7P2zc7jIJ8cTnnZ68cKQ23DMYsCUmU6P
d3rCzb4AHhncXAfYnsLYAGB+Dzp2pw3KYnVRH6TMblEvs7rnS0LqB93rrdlBPoAlbyx/RXAOBX54
Gye+QDposp1257ZrIZiZvznYOfBISGbYI259Na2+6g+pWaCMB/sSkhMWXqrbVYuqC+u4eqrb/5pM
uGOFWrI+ne9ve3YrdjTu5Y0isvZ3YJHMz5VWeugo+h9EMTXUlFPCLNh3cNDL1yD+5g1dKOi7fo/7
RsPnNetvGluL1D/+LoZbKx2hpF/F/wLpzUMSHRGlL39xAlHeRg2s7PjCoKO6xBeV7ASjMm3rr0O1
gXI1FUTqFKU+wtGdDWSm+S5p/usXLL1L4WUjj6RpCsoxwtb8UR3JUjaWIFc2jSLtE4gUKd2bYwvp
4RzK8b3u40bwxTQkw3SwbfQn2GKhLUA2gtJT8+4p1xWnY/2SjqL0N/Tgok+iZXS2XwUPSMD8r1OU
pHpFjSBBxTPM6h5cuce33Jz7q18fJOhXmkuvY61bCyqJzjfNmDfIe0sC8kIeU6Vlfy8yIdDNs4IM
eCJxklDRqPKeXdTCLoXrTRbsnLyHwzE80oQY0ZAg+OCAUABg2zFZTxmoQpRgu3ItkHlci2pGBW2h
o8xX+YOS0EgfSstfJKi06b3O3HKXrppa1C/QYTvrDzhdUVwjKid5a2Bh/Rf+A0Q1iwcDSeHj62Vn
W+nUpBaZyeFi+1c2Voq/xf/hV3247ZEJyRQ1hODoqsaH7qtck6KpnsGNjkgZksJ+e4Qa4/sUHwnW
rwZfhlso7aAxhM8PD32Qlo2w5xVP65IcMkAsjGR34e4juEqJgJgnawe5nr5GKyQBdxLTQrGUU5+m
KkvxWvPLCWJrhnQ/StarkLMLc4YvMvHMZ2zmf5HFOq/wZf7S9E3j2UzNElqr60MxVS42iirdEaMs
1y/vib7C9yr0Ando0Btv0sCeyyJbUJopMNt6uuWKHCgXvohjkdZUBqoOECW/xb4/heJ6s5u7hmbO
CouhopC5UhR5VG+xuv/QRoWVJ8+WInu43v/7hWrMCkwlUDgWhyqoCrLbnLR0l0mHr0VtzqmFt/Jz
OdNB6nAJnkBmxIv7X8g3Fwh4BW6ZrYynuNBvrQPyIctAJMTgxHF28l9Sgro8eS9glYdhG5M5xC41
TSchs9mtRNC7M9fRmrpzOeaIgUUU4/Bm1TetrpQZvitATcQZ+Mq8Oo3N1kM+KWXHI42+vbgeIpj3
Dyd0kpvPVBNBsvHTfd46K93cRt9yr/KCWWXQ0CKX3XDaF9GlLT570BVnPkCLZj702tijT1Tx+LPF
LJp819UV3uv6GzYVqtg5qFYMsMsSgSMG9ukB/VaKRM/0qoYTiqKJ65+bzZsTlRyddqjsy2h8xRgo
G454oTkdbP/n+lqckBNK3XXSjMgj5QdBoG9Dla2VsVAcMsWsFVin+Qa4V+Do9GCJA7uy0MMSqPfp
wo4xZjEXAR4EDMH7Z+rO0c4sTwEVOvrLs4iB7dkRaolJYZuWhziX+ed0W/CQZ33L0QmTWYLOJRFu
McXACHWDPS+GUmMk7chM+ogNbQ2gN2CFN4KIDRDBNiglcSJpE2KnpgvFelMW7FB/lF0hYes3B97Y
RMGlio3oSBpa/579m0SLoLHAL6RAwK+TPLSyWCPdMEsxlyeRb5cyciAoNoraXd/BfBPylrRfsSJ7
+lgzfEFS5dmaV4nNgDCFL3e5HDhU5lrFT1mYtKla0BeEBO3TpSVbd5clupT8EssVT580mNVNSQik
DZSiYKQ7ELSorWYwnuUSwpijqapBjw3L5wzrpljnrKj8SRUw/EuryR8gG09P4h5DmRDB/ccO3Kjb
4xWoLLXx81dtXx/3Hdfhoz2mR0xMXZetfmB3aqncsT+jsnJ0WASOMIXFI9YAkihhl1J1HXzmJ/5J
xQOIhy9fGhhs5NCid+ALLd3OWPAR2FSCzUOSP0KcSfa8+SHIF4FbMV9kqeLbbrC1+lxNB49RP/rQ
FaxIA6HUN43+33ITRSwPQ7QbZply+chGOMFaGx0wO5XB//GKxkfWzTajWsGWoOu+VnAbiccSOSJ/
5bBLSfZQco7mrNt56YB1Cc1xU/YCGgyRfROfurTxpfIj05m8qJvLLaPGihte7MmWbP/7FhymnW0w
GEmvCEY8U4H4hTZ+/26jGXxMmVILj++72x5Swqzkqt5nJDxUweXuLU8c5RLUZx8c84prCwbtQ/mz
KQ3R6TPfXJyCTrQfK4yGFFvFl6DSSVHwpKf4B/LJESjgfODZ/ZYWZgCc3aXeLCCSDCOSEjCsR+iQ
5PSe25G/0bc/blAf5ShfACSUxhlNmGsW4B9ytVGjCglT9nv3qvO+2/dJty+gAAljIVCFa+Sc7LW2
viQ+W/c6mvBZ/fM2fJiE2Oae7cdLO8dlk14cG7CWvyPHBDCs28J5gew/oPW3rxc2VJ1LO8Yw8TAz
GaNoHDjC1z5VZdlDuART7FMryHKLnblfq/i3sBooges0LOH1DX4ox7umURoDPznKc4SrxhWJ5tsc
Kp/Z1bzRR2h5ch5YzliRNLTc8kp0ZVxtC5JAgrSmFDZVeYuQb+IE/HoOMJizsK8Hc/7zSBgw8BCQ
q6MnjQipv5eI6D4UjeSzSKIpQpW76hUW8OuYM/GJpuRoQeJEjnSl2qjMTYBYf0CbL5oJ7WZCGYc2
xtZ3tyyYxnebV8GzrC8bnWM5djo0NgO6FSB0I0GKMeOVsxETO812BSpClbxNLYc8w6z1rCgcY3H3
vd7mEx+hNqH7QRv680ZXQ1ignpuAz3mYQ2l00PBaaWj9vrNqZJD+/WljiVjc4MeFm7XH4FZy5KQB
5kihCOu1nEMSfg73hFSyvlg7EahxjOpGiGMvPyHF5NFmipgEluLxOMtnbYdkX+bCMdumT8pVVNl/
lLvH8iV4gkMbqk88RggPpXjY+X02nfz+FmB8tMb+v/o7H6RwlnYVr3j8FnTg/WWwQ6xZlbL9YEWu
e5oBXCNBgUFDebPumsEMzDPBEGIcDbVnZl4x8bqr9Q7cw85gwL1BGJb0p0CUOZg/8a+hDLEclsjZ
5DfnPKjPs+u9oYx5HevDlxv7yfktGZDDbdcW00SN7Zt/hvnB0gxAsSffEMOFEHdRWwhUw+OiAUjg
IiNCyYm/V6nxJ8qZ4r3qRROLavs+A99uJCko5+Z3gcrNSBSCr/GDtuucBCCxHVhFchBD9h0LZHCL
V9tqV82nMY1i2EeYpcAhNIyelIzzCC+/NKF9jhWHRKPsL6vxeNzY2lEl8tHI2m+xeWSGtJ1Gs409
nGQXSt3RU3JSmzVlNF147g18cadIqFkB4vCxwXzJhek4nv5tr75ThArL+mnpUy/jBeUMF1UOMqBm
4wDgSfsyV13719p83n854N715g3//hyMIzTQJfrx7G6GZDZEdFy3L9s5NPb4zboMIoRP9H5Es4UL
pOofL10vOQONjp+lGTFniSuzgZUxs8x5jAjEtDr6q7SWnc4X/E8RiOVyF9N4YINdrvyuQxlp2b3T
Dr2jcw2W9QiYGWHCI7zsy6l6+gggUrwOmr3Vp5hr6rU+DcFWwcaEO4ZBKRu0p8CN2HyLnG/xHFfe
kSzDsYr7zWrBtAjQWaXTrGPN3Kywo+jConhdBqS8s5xgfRy4iAVGqmbseaP31Ak1MOzLlva5q1Ar
mNwBCtLQIYnrQP+x75Fh50rAg+WPGqOKVL9jfVP0fVy10wzDJk6JehPnXUG04vaY3dpAGGwOGzI7
gpNWhrqwrDjOpoL/nO5Q6InVLQO0gvfmdjbuYqeVYNAhoH8kTgC3web0dIfq8sadA10gNi9uy2G/
J1jXWTUEIWtebLjDJ7PY7sw853xWBty9AkuP0zPHv58tcNJ/He2tHSYg1qwhyMMebru4znnEbJk3
yvGtGvvgWeUXEGYaw7WBmzYhtqfBwYylBrgovHf3IuL2oX3pUqO5Q2XgajTEUuNBrOxkKvXkAXLa
EHm+H6TPod+dJJ96CPKXsubBKOOHWeqyMH95FUSAQyopaqeH/C3vG2wfa25UX2wcoQalWm71AxtU
ItPqYyqSI9bqI50lZfMY0HA7hFYv+cU2ARfOh4pULKNMch/Pipxak4C2vKuS0TiHZLLeZ9x0EhXe
qWGmMm4opSgDHFrHGt1XcGyKMQSgyHtMWz6Msv1RlQBTtL6siByLpYR5AkghJRB0G7GFJqmc6W7r
dPAi0XfUKCCiI2LY5okQVaUqIbp/sRaaf3CCr33V+BSq8zvOqBQ7EvCDHwWr9BjpU44LIXp3rJx1
AbXOC8S9hDYqYVXDNtM3LnFnRs09xSCZcSBV6e9/RZWtbImUbr0jCq9QXEdxJ/mBSF8Y3W4migBU
tvOqn4q3hnQIPfvtM0iV+9uk6fPfH5VnTXWZRJQxTcl+XYD2K8G2khf68CRGhOL6Pra59uUP5yt6
iKP4slLQcPVRQoca5MFRuiWoL9nZcgPaOQ3S9p04OK16E8y/6Za+JOCUSlwOsWWi8GysIWr2CZpP
UZArvAohPnDueV1LnDLDchoUxLeHrNjs6UoPs6nwpYaVCypKCblEgNjw10ViLEEKYixX+7szd6NW
RFyoHg18SDi8sZKzdoyZ8Q1CodmzMiLTFui0iJXLlh+1qNo1LGTATT6uzenNFPsJihwADWReshnd
gVVLemMltROGkfY+IFhThYTnEar3teO0jNdKQzAVCJehNuq4RbXCwCgCWzAF+QiMrwaUUc5d2OCS
toPvZ6iqKwwJ+WbvVM631+OKFLN3m7ueDmXgVjCN75BduW0xTNBu2keECDshzEzOOd4/EYMVpQ1L
MfO3Lds11lynrMeN9QxdEICQ+ilmMBcOfsShFXE9hiM+l+hxnDclq6F6BwBXOd6O/JImHF8iPacd
zclcRTXG4lA8dpGZ3OgSnHy06bs69tZBdzrTW9oRz411x8yVdP5bISthbamQXsPQ+L+xFO37nUqi
jmxRHleULDTdeVDKkHZC096AzEzDTOzZ7dw2FEYZssTy7onxVzNrikw8FbZJiPQxsPMWGY2rezdo
mnSfsvGXB7lTcMwJr88iZroSWFXtchaaT7jPbU7dV1hxDnQmB6vP/hT4/Dbo7nkGHuzvCQrjyKA1
kAep6GvVUT8tDMXktrKYssA5pjymiunq4HbvsQdJRPu900cmbbvy7l9wx3pchLW/a+FvioQedIt1
WpsJqB+Zkbs3NfjWQ5oJ7zfO8Qb39+XpTNP3imZz5M3CZ7NPjP6CXkFA4stjZHF8SlmVyfv7zPZ+
5GqUua2JQafPXBVPr/uWCHAAobAncYQ7TOoS7KHWYFmv+9ff/NlNiUhyPOBdwDg9C4Y5dz78ZZLx
GhEygHs9BwU03d6wBsU3F1ojjj3YN/SQMTZtP1RQLkE9D6OsJdTA/yOSo0PnXMwIjuZlTRzar4nn
cENF2oEk2l7Bf5c9UIUReyo9aAu5I9RUvnuvP98zayN2ZEEyjSIUG0uLDOWt1WEY/z2ivgAOojN5
gqypV45Xe00D/jEydVuxzZWgj7zBpWjMTMqiLvLHGb1jntDirbxml1D7nH7cckRFhUCr8DsGR/q6
r5MYQeZ0BEDbNDQadU5QIPDBqyEr9viqfFOTPIqVF571On/Vi38pratiFaf34/vpOyWFK24mc5JW
oOfSS6OtzeiGNHCC0WX7Ccd0GH+vzwWMMlkXDDB4M/Y2oPi2xANYFTzy4Jabotm6uE+6cIpWUn2a
NTzrWit2MJ8J2bL93QQTzyGzi8fYq8yMVcZuJ9iSx8MmlclaqM0wjCsnzFxtxQUQCi5uww7LTpZt
L8yZAMdwZTvPejjwBkXmpcgA80RoybH8VbhP/jK7pk7riLALTPP0MLCRZHY+2KN3rIUhTg8Vyz59
iQUUMgFecOgMMheUgVX7GS6HSJCVa/jIv3O1t38Rp/tnnBbGXnnzbXKJISzNEF1Np6NpYqzZJxHq
1kA16ms8bcZSU9wr7s55ya5l2OHLY0AKNlpcWLk9VPQ12NPc5Oj+3eeOwM1ucjqfrGe3AR6hDTDX
BHcZ/ChRNhKrEEGZFWD+6nSJU5nkLbU411LyDPvdsk8Wok+uHBJWcjsbSUuelFvl8uLQgaEXteLI
Hi5hol0AekA/gjsosaizqR5FWzuIbOWY3rAhsKC06ywOMRKXi3IQakzwrqLMJV3VGbGlm3WPLXiH
L1qwDBvAx475/FzmnzOHOltZ91KrGJ3Ems22CA0/TB5JG/z5sbu833odi3aHhVCpyekkIEIaKle1
6Im1q+tDV7VgchCv3tT/+k/FWbkoJ5rTl2zCWkhK/Psem3LrvUPKZBbYzqEoeWCf5+mb1fN9HTyZ
IhU1Anx6ufiyo00g5VZWhNUpV1EupivwU+pIUGPmop97P42shEgNkOG7rVbv/XTIB9InhVOMmMEg
BELCvJ7IxuIk+zXJ0zt7t51Xj/8V/ob8oia7pUwGwIYGu/Dc+Yf+3jUGo0NoA6ms7ZbbeJHhTObP
wYSKdHTBmcqlMisOz/3tvNEBV0FCUMRSxyTbWmC5fvm9bg6rwx+exxgv25xgDJwmrCmn49aqVU/o
4Rop7MdvVs0ykkY9N62gDpzmmWE6aJZ2EPwjAcapnQBxdZyqqwBlHs1x547wcUFzXSwteZCcuG+I
jDQQII6BrUazAJGeVw+r3YAD9e464dkY7A+mybiu63uU/F6d/eLq5MlArNjqQ5owEY5jiir1RTXP
Jtvgyf3ubuCd2DvxMJvz8xVlQ2wRYQ7C5MXwn0EuykPYcAsYaMy5QEvgHYfWfcoU/RGz1oykcm7T
qOrRB7Kvc1GjrGfhqezb6qS3cW9svPACu7fDIoxQz68nss6Nl8nPs7lF5651qkh35ve+FjTNsfGb
m724OITx+ibccqxXmR2SEj5wfsoNGiwZGJID+xHqg5/J4a+yNzsDwqUOM19vyPGJccJ5s4vOdxH4
ARdUDvBJKkUcD3M5zyA6N06w/ztq5ZH8fu6Iz97RIfp4oRYXVltSAm+zzh5xtTbAQSOG0gy3Nb9n
GUV4lelHAf96T+ikxjAv/Y2D0fGRQ5tcuRmWoMxwj7Gtkl72w+iZwFrCENKc9M3afC4h+PBCM0Yf
tgQqF3b/L3aK8/Mr3jp9lKCzZ4VRiGmv1qEF8wby9jGd8P5hh5WwncN3dLPgdLc4WtVvqXUHePem
rUACNTjyhW1k51KwXhhdDPNh96b0aDqFmbH3TgUgTq2HHSyLnVg9vhxYwVGbfYR4RG39ERjzZR87
Q3ekkalSvLON2o62b4AgzA9jYEKMbWVCKGnZyZo+vupdW6FVGN/TTHyXKlD3AxulwMzXqRMjwxvn
5pTKkLAQNe71+Mtvt8FnwggHysGrpGXNoIHU3xc4q7x4SlnVAGC9z9xUtlvyJWGxttIuUd3SPeRX
tQAnHj58t80kbg4TOoAiCfsjMJ+mzYbMpQO4VenXo/euI/5de3yMUCXGYCdNVI52dCt0BQk2ZO2D
7sXR7/L1k4469XVBNEKVGa8GRrxfNkAHsIScvVaIWWeXu7+/McJw0wrX88TigpOaeHlL02v5q9uI
PvkkVN1rtyn99yz6Ea4AJjkPxsJSQsNoIzlFM2SOTSXfJMD9I3vHXuxEvnX39fjakSuxecdNnxaU
JxS33hqo8nG0OZjsMoRpLlvOh/JoQpxyh123fCV8nbxEqOWwYM5y/+72SbkYJSLmPD8HZeUPcAJV
qsXztSrJyp4BuXlHopWhfTieOfjZwYzdk27Px52yMOWvlOjhaVcg1a5bSUqTYONzRof0ycQED1/E
13UZWbi6OfyLNJb27U/CN6pw2f0bTHu45wDjCEPD9+7nOJ4IpmDU3yD/oQPO2brjkPCaxsmo2zz+
TZy86+qI2oUhj57jaObj4qCfg/L5WIU9YQyr2YLfeJNPrC6ouTnyNqOtVbY2+dXjZjwh8SE+H0pt
x/x+l+QllTYil1haLyFraAWaNXa0/yyte6XRW6HGsFTWB/rb3LUlpYO7y696nwUo15Yjt1I66JvY
W7hQavylOY44Y7ufu75BD2J1iYUh2zFWjCYipDu3PMPrzFlzqJ0PELX0R2GHC4PFTJH4pGY3Kq8k
DSBOGl6fuFiQXx1GG+l88fx85EUwaeZfFD3m7isOyLpzDuRqFULgzogpWuZ+OzYeA9cAiV7gQNZO
5thoLypyieycJnWi3lgxu/O15hELQIIYFeIDH12MSe57PyHwC9kCFj5vBNFMJQMO12aNc7DlTGSd
SAZ4YLU+MP8s9EmJQxPtuBGmiZPNYjLqBRcRJ15hSQzO9DmSJ4EAu4uv2LNs5O3fTAMdkiefAGhN
JdNRVg31ihZY5QCGDmujr5OTcM5FjY0NCQxzKmsICkof8JwaWKIBUvxtXQGidkLHcp3WuI+w5xQK
oz16cnaMyaThMxPXwF9vbo8n+szbVxaE0flWkyJFdTphw05zsTBZ7WtUyLwstjlgjtmlxBKaxJZM
ITwdIyYrwJzsLtrL6IAlKbXWOgfGUR0KJ8UOcvcQhfqq+fJ6bdgQV8nC2jUL3wzB1+QLS2yur33b
NkVtPyT6WkeerLqDxAUglm1RXcl0zRzDcgjLOIZybUwnfj0vCI//q9xHDA9Z5z7VFSjxtg3mM3hS
HKjGjMHKq/sErYfjJDpGSfHiZ4rV0A5rstbYbeC8fWiyvAWWyD0oZhjTdSu3wl+6nCBGvh0gT5Ni
N4hw0G71H92j/qvMLFXgPmWcilLrsFgEX5yW+Nk1k+7NTFP+tl3fWxLXmS4ChDWRKT+KhouHcrWd
SDkyQ1M562cG7BseSLSwlj4znQQGonLTLSUMeZJKeQgbunb4/G/R+zOHzpitxwF/GzCi7CdaD+Go
KGKOIzS1NCR+UsUxUY8tYOZ0iOr/7n2krd9yfTUPdvzMl4S3QCKGW4u21T+6xvmO3+Q9rB+qeE3I
ABSz3T4Zz5EESjw4gvxYXDB+OuzMdCZ+qoc5zJRw7DMo73lEb8dlvrJp8A8v5YL0fhjlrfXTAvU7
XH/ha6m2niYkgK66c1Q7LNJGB2JqnsY7EwpsvFxOciK0mO95wTDqhj/27vbS42RmH5dh994p6kSF
xd+BnFlz0kAtVPEIrreESzlbqsP4x37pB8T0gL4LppABb01ch5OPYCpiqqEJOITC6JEzTx4h7vMu
e+7FEIW1n5OKOGhHm1VJlK1+yTp4nf0W9tnNwg6wOFd7VfKQdUC1ed5+E+htFx27oXBddXcNa4iJ
4D6Xh8MT07PtBbky7DpBEwtq4irFwMGuVrjPj1wNjzwoAGbCTxBAbQnKYzstLhIdqe1thw2DZ2S7
wlfH5W9By+QQYk67jkuzGTZwvgOavVEBIncWCStxm6aCSX7L7kPLgtqDrbwNx7nGCbjCtSWQWG2A
ZQ3Qvq+BlQktBY71brjCkePo61MbIlpk6PQpatGyz2XghctF4sXc15tTJW9Jea4xkL9FIUhXAqiv
1/UE6xx/1xCSr2lkv9QN92QYTrISB4/3U+6hkDTQruWmLLaqdBkCr5SA6XmOKhI8yeLnUcPn9ciU
v91tS0mKI1vWRU5AFuEDkk3FnBUEexGixvkL0307GLL2tBKf5wczCKSCYnpNWmi5Fa6ioxWP094v
+fPnjeZkuSzan9iA2VRvS6A/IQsqrNLJOfPS3WCGtJt6XqUae7Pha6/Aykok/mPJ/ux/GGHngEi4
C5V5/m+gr2JRjXKkl3t8YtiubfwOv1t84ovNpsEFXzgCA5X7ROx77tBgifH5kJ60hEu3CYc4uuLY
o1bwNANakqvo5JHXn+HNChtrv5IzU3XUxaCna6y+PsScKySQrGTGt8ZsDMZ8r369pLSdZlPLcUOr
4cAOAx8cPEDX0ttNnemdy5j3oRXwYQj+1RNxoNLzj7K0SW4HPaKxjSW+UAM/vjyWwoIohQGFV1KJ
pcsRmzetBicpNAy3bgzK1FbvFPihG9LDVwnXv0Xr/hR2wcXoPwJvySq87ocN+t6VUb7audV0rklC
icxRYiyfzzFbH//iW7YwtfpxgbkX1Kx2yMGQZoiFTisAs8LjTK/GwremZGT0Vg/7ZXgXLJCVUfb3
MALgCjpaNCoa31SyGPRVNfMONiVh4XtZoj/phHAmxyr33PkyQE34Ko6KteoUj7URb1Hqpx2wXBVE
tuWiqqAcEhMXGsNIszafIp5KQs3LeouYZS36d9ZggB/JcNE86pPGXKqd+pXb0NJy1pUMjAGt7hMb
5Ee5laHr4dJ7V0r7wNc7/WI4JyAt2OI5xvl5WFdmvfzJ8alkCxIwgkMP1ymJzgHIkqciMxQNlzWc
R2Rz2W5czV57fG5wj1e91/NOHSI4ioFkTPr2Wltyju5N93q7DuBuTj0jtfr8GA5oS1+WSUhQDpDL
+HWBwMcVabtCRbP4rZyoQoSA3MKW9u9RN06/BiKn6vrwdJgMwp+DAzgDG3+buGIjTBYFJcFaIEHf
HpDDugaApBkgV/+nJHmb/CHLEH0YCCmNK43SITfHyghzUr5NFsPVxzyxCF58tc0zkMP8PyNKwBqD
1wKXrjGQD8x7b5bq03WP2Mx1OAVn0gRHRBidVfzZrHxzxx7du2G0eH4FDNbYh5uOfbp5CkstkYbj
4ZN5Q35IIGCQwnwBfKWAH24OmzP8shtWc/NXnGEZQJO4NgQ3czBlnugzVZVgwu8W2aeUN4P53dKA
BGiduvS7mvIyUL8vDuBqF0Gvl1dWf0wTmwC9aTs7Q/3TnjwtSIcCuGxdS4udMKlXWdW2WSBl0lLa
Q64ZX9lkIF8ZNIIxXePWuVyanLnmxoVsSHq1SpMRJCLz5SCJDQ4brJ11j54g+wrUUuk82hzVn2g5
Gc/VsiRJBVg8pBo6WAbceCHZsyNYrokI1P2B/nQvwX0LIZlZMHul/XEm30DeD3yeUMZY/usdbX0Z
jDC7b6eXi0XXfSLQqwSMWVoAbAE4ri6nJG8mn83N+fcdP9rlAY31u8rRZZ+ga6Qvrw6r+DDrQAEo
8WPGYcA0lmz3WPr99LoBOaBoBrd1cWngciIDLM352cgC1OpGPuR76zSy4e8AyNOAjxH2kLgDvb9J
+pO/lN2HS+8xqHMuFJ2qpsBa19udIgX0vglhsO7erqw/NanUn+jZBRG/pZTzDlt4hvAc/ALWicFT
mYA5NisMtHqRt/6EzAlSMAniPidZIqQV0RJGcvW14gJUUGllTejrsgbo5BQcxhu0GE7V1QaEbgVM
R/VA0LCy1ikPRhvv1jWf88KihLuvhlcJ7jdC0gw4LJ6LxWM00fBazTtMqTB/aXR8i4ynFFh04NYS
NTSO4hq+eLeMeLFN6b/cG0/W/UqcXPgvFqvog1KqrrtmMWkrW8MnPl3lCg5/oAThrOU0CW9qNfz+
FMc1lC6So1aFBdN3+VLcAkVGXarSgniTyq8st2WG5/i9zEAO960Q3EoNJmHRSNTjOKVtLkcp8xs/
qJld1Y7q9BKkMllgKPan4rF9CcNH9iW3h1Hgbj/vEh2fwGrocaFSJMNyYDw++avT1Oeu07gQCLaP
wkmTT3eoM33ZA8B64+gUB+dVrJ9/QQllY+in3iz5ROv15gkEjG0QyyCXPG3r4z8z1OXqhZxL++ON
dDu+oomoDdhM5lJQaRxPMePIUOCXE1SHoJVRCrexy5TdESCIoVl2TzOqTV65ofbw/DcPj4cc4Uam
GyAV4JULSVnHXxlETVIVMHifnKdPJ1sR0KmsSOp1MAo9CA/9Sbv9s5atD2J/kJdy3Bqy9Dem6EtQ
AOl1/yyvNTKxhxZalACafAxk0OVZYDklnJYcMLGn+0yy5sN4i+HNeQmrY9kzcD8uepCiWa9azW/h
2HjlZzUrvFjOnShJLyr8D7TsJifCzK1fhHZOM45sAD38oFss+IRxRECiHQJ7gZ3eWDdiqNwzz9OR
s0P5jmN1pfvc3sNXyWd78qUFnd+UbDJ4AGgoNWBCTJ1KtwGo8CvCHKSOGHw8Q2OpeMJKJcxP0GuT
uyFm0C44EARI9q52hy0TyQF7s/KIdjjNB/vpD++L0pSTYFg/yFgGyUW7rp1KTIo6UbEu5vm7j0k9
t5V0SAEnskgao3g7fgxosZWXWd2nhxtcIlv2JjBiqejAzTNIMkbCguWUNpbfGbKrgPUGcnsRkWlD
0MwTET1RLdpMVCE52XHFXe9tO3J9jcDOiVKoamABTADJxLSTsBB1c8J1iEbmhN90TiQF2X9+tjoR
kcxce1HLEnenRXhTcT77cY3RByqTY3kFs6/NCiQjqO2QcmsuobD8XntluPvxRJ3PdMkO8GU8ihzc
UvLHfDhumGIkUwVvFrqghS6iJ0fNzvAQX0B2k4Eku33QPuPnJm7F98W9efPpUGYwbkZKNtvJl0wi
cOnEJGO0SW3Q9QMs9VFtglU9fimArgrt/gZQhd79xDehq/f5h4WgBaLVsdTtS3i/fSdWQ95EYLDb
3X3o1UmyIAJAasHj+H7CHXl8Kl1sQOhcJ57VnBS9WaEBZS19j6MhYlAU3HEIsO+4AlsDkMyPvw2e
aDFrz0qAwlQnbl9qzw8BbzkwroWz8OKNeSOmwK2WoLG0EaB5Dw4VHxb4Li9S4U96DuJtPpw2SBTA
y7dLwpngOCGeWqXM6ikY96iWD9p2ISl5EA02FA7PgUZYXuOEwK46Cwn5iMRCgzrDlXxavFHlxczP
m/Kaw51QK9It5299dwrfar0P9Q5acrwZpHXcVsOSWIqFh4lm5MlIhBAmDLBrD53YyCYq6kWglUfG
U/dB0/3F9778gwNogsysrI+PtRPxzJ8XCigrjN3nBnI0Y4dkS19EoI9ZMh1LxZXFyu4929zQv6G3
kbZDXLYcBUuvBXjVcFkhbuzpBB07FY44TFaTYVhj1Kpy21CyMrj1LO5+Mgu0hyZTBP1TdbZSDUYQ
fVfj0pJkjFBwD8rVorAq2tu3CBWCdVKM1xRNm9kXQAfji5RX8ely8e7D1MSZ8WsSxQumEMhRviyb
plZ8y4yzWtXrkt3Svl7TqaObxRV1cqLGyVz/wbl6n/UYwmHIqnubPeB5Dp+LZ4WuahHc5DeUUWcE
/MnF4CaXjd4rCoRBlv3bjPo7qHftrR1rO09O/FQDMBg33OPlGvk4LNXTlrWNXpRStJlmLWbRGvKv
7DQ8v4sqryUteY+b8r2s5/HK7NxwSFDTkiNgt19Zc+gOvk9bIMeNqLVOclekfjCsC5jcA3qYp79F
lKVOZVxm3rfPwY+FSonT/VXufxPHFX9zkJaW6ReeSTd7bA7wkBmGneA7fmwoZD7dZpRNNihtLe8c
oPi6gkWylOLjonXgk/R2cr9lHnwAmaJxEPSMthU5JAHp/KTecqb8g/LJefDV2XKXHDt5Oi/bLu/v
RcsBK/BJmiqQqd+ZNmCXTrQm+U2enblt+yb5K48nn6nVkpSPvqXCG0Hfj62bSoV3LykZPrUK7a4C
5BaD5bfLbGpfBEglVad7Pw5bi5MS6mgvGRiPUgPppI/8d5GKT1XDd8dMGkh/E3BdBmz5Xjr2FPdp
gao+cNGmRiIOL37V54US4Rh+wRFUrT3UPI3VmPIZDAwTTkY/thuRFhvB/TRLffUxdy6tMeiqzNy6
A1q6eKS/U5R3u5vkeq9MJubvyk8VN/1RYtDq+8QMcobRfm+upR4VHt5hG4/BzkcPlT8EbuKSbr0Y
VC1An8UqaVPfgx0fYd9/gCurUDf8AFAAKY/lGNUcS1DH9UqFj7LuOsXLMxztGq53mXWccaPlhkHb
ZupgBysuU4qLcbr1DPwHwnyAz1C5ZvbeQ0BwMf3ANG+GOoccgyxjqJrqol3Mv5jhlWEBJEJq6oDG
4qAZmf1CxejC+HkF6Rj9cUk88YCd7xo766rV6wmtw2O5Ri3OdXY3Ma27rDEfkgzYR+v96qKwSFYS
nwl9yHYW4eAqYkJtiYCn0sqIg4KLr3zwZkkQH071FbMibPmaeavMGRQxgKrLQXBU+DFMo84x78pV
b4uPma9rAsaf9ZaSp/liRfxgsTi+8nNXwSi/uFUT+H5CKsWch0+m+4DaWFPP47mWxUjn4NvW4dc7
dOstywkdtNokzd1e67qfknxKs7XwHO7vpblOMnwrwNExjjvt54fmzvmYniRnDwu74m96zK4R716N
ln5Jry46SQxtGDp+g3ClT2UkAebvzy74VOXlAJ/RXhxBhNW/cZJhZ6cDm15nwAmNk9u/UQPhLy+B
YNx/JZX1yFZodHO+0avv2eauGKFIcYqoX9/nHx9oelM9RkUr6o8AJbVbOCJWewJ/PSUeMBfnIop1
hkaKgYbsSQY1RlaoZNYTqWbSR9B3A4aR08Sk8P20+nzpdQuUYuXR9nS8rDKgVbLtbs6Ycwzd34Lb
JgN+gmcs1hMg/HyYS3qsOivgBHJIQa59/II+I1RHJbjxadb4UY+HgOBCJsrshTpUiXHWKH168sZP
XaTsvMwqQUs5/RnGrwAB9KBzjnAtkTV/voeheqSWaNZqsnwDsi+yuxF+Ykp/eFRk/dQWrtihHVY6
Mu2dB3E7AMg0sxULYU0UgyF7ESets9xN9hUuqB21l61wyLsqDjBtMC+aGt0OKVWXnjei+pVOQKEU
6Hselcoziy1PN2ERS8dZ2Q9OkXZC6fPZ6lKHjdHipc5hL/5xK65/ERYYNOROGXuifGwkw7MqnyJe
OARkXfWGiR6iyIs7PoxxxwF0tAYMVx3Qtsr4S/1VdVXnKUOvYvQ/u13lD9c5/5oAuPn5eNJPtJYb
Ad4MHYvSG2AlDMerpiUhjc8OXCQZan69dYIM0HhQe9FHAB6W7RQVQXPEXvi1jfcaCDbgB1aLP/ur
0yubQkItAOCU6Z4+HngRvJ1zWAjtxCR79ixo4rJJiMCYn/M0WzOD9A1pLH2VZKMnM95aEMrD47dE
fjroAB1p0/IF6DQ2i40MCZTa+uLnfZF+Wzqpq9iDvP583Bl0icV5dGqRTtwr+8Z2kqIJKYwDMcVy
fVraDIVUnmgZkPKI3D0OndSFlMxZ2D54TPHTTN9OgXjm4b5mNIJqLoutmbYvjT0GNcThDMY9lO3m
NCtIQYnJhhERB7LtceXwMhK2QstwUuPSQHIZCpb4hbALbimPxeud4eQeUmC8p94nS35Jm9or+2RD
uVTG155KEqu2xLhaeYB0rdYXGw20i5CDjmd769mYD7x+FbJUheCKhXhBPF/CC3Zx6iLhIk3WWiwD
IwBqweL3ohCFkQxcWEsmZ7PHSYevpLHeRRQBxo/B7BMkKkUOu8yJw1yQLZZ2hKkj4QOlU/JNx8fU
6oCvgUyZNuWbbHS9WzkywsD8l4AI4QJPKMUB3qrZgn9FP8QTMFVC7Q8EpqcQNDaomfT6D6TscDUx
pTrZl3II5uZZyZ09Q5mjIAfyFJPUGxTCW06yYsSd0rcWc6JYpm9/nDCGMH0G2L/jcF4bvKiIwTAA
JWGfWHZazu+PAYcyt8f5uD0xr4d+g9CsPPV7foxq4EcIzN3Mc9H1PpLo4AkWMdzA0BRF9jWd53T3
XeQtva+MzKOxIQQdjLjO03Nw0GfCNa8oXeTHRqTQSCC+GC0D5waDCN6Mrs4yrNrywAkGKlaF4tMw
fr0w6No/izqFV8f5GwkjLEHBXfCXT0Dhe74muXx7B5OT1hNyUa1Z2rnH2gh4LHumzq/1J/xY2120
Vu+rgO5SxwVaIKgKZ2CsH47ZcxukeBtuKb6AKktFOW9koLUQeRtuV/1jFtCfFyakxz/GDxjP336Z
ibE4NlXX4FL42LMr6NSIbefJtyUTN9UO6EhpiR+0jkkr1/Cu8n3RK2PlgF4OmYvEJPhJGDHyibJ7
Qz0tD/6v8W4ORXQVVJBuMxN06Vfv59HvVw+HzETiGz73oi4vZlnRjpH2xP6E/yR2hC4ym9j1NbSI
/RF+/HTmQ8CG8qoblmB6hHRg/uknHNB87ICofHN5VAWwkWea/Ig2c211K43Twzo1tXmbpO68/uQ4
FtGN+AN34Q+9MIO3Wt6N5QKdiTS+6+YCvaeoyD+F2pwyJXNsKZFYI1vFt4R9/nkKSwlE39gpePoW
7xaycKccpVhdy9CfuWbCL+Q8rPxKyI/mmtqvlxF7hiWU6SrQBEvoD8POHDepy9bRcl5hAXqqaM/B
r+EXs+sAlouk0FT1uHpZHkSYZGspdeMe2Qpib50Ln8JH036iKr4i9ZOUvJ55kdqNE3mihGnFCHAj
7GiRV+wELBJFYcZ6O3bNGkBaKUePcuMK2DctdrIXAUQj9TJ6w5FW+asp23VriDaqDknnSF/GGTrq
aamG+KOCXebcYY6GZfCtKXuk3snB5O4m2P25li0KMJcQXkp2S7qRzI0xTG1aA0GxrjTZIzbf2aFA
sJiBvK5RBkkOfGsMPgYiIlOCPx12XuMxCxh4VIk2g02rXNGSvwIRcT5eZY5aecBB3zl1LvIAT9R2
+aylMZ2Ph6rvBOkNZk35kXG61mJGp+RjH35IaJIvUNVsak/BBEe2zrp2KOtDEVPHvAxHjr2Esg+r
jMphTq63Ljztg0VYmoqymTvevu6XXLOtmm2Rhff4MJCdT54xeeshM16iQad3RCZYC5URMkYLq7mp
Z6Mhazv1P9hlUjHQNE/AmELiEVGShQszjOzLiG3wAPhbE8AC2z7xglCZz6FiDE6C1w5zEuKlVkYG
VpzuRFDGROnTnTq6lhHZT3k+8D0wqpXFRlYOYLlR1QwyKYpeD9QS4s+SWeNJBo6Xs+kMeditdTYh
/qBZvLFk/1SS/2iBapVyQq8NOqHVEwPj4l9Uoxdi8BuARt7mxs35RxHfhSdsQ6ai8HErHJCIzaYZ
lWtAlHJh1x/1KwiF0nAXRFBIy12ZBTOXmzEBLSE3hXNHG031OCAz48qOLhGAvU3ZvI6kZvrPbP8u
63o+rehAaOEDlrEgnVi0JZ0+FEGR4RyQhsCv2eoxKBfpPZibvLHztm+Yq7iJdWR5X/Wv6DjBfwgu
insleNYYLuX1lAOj1YO1+vVQr99K63AopkYNE+TRdStpXpo/vu7FVkYprie00Ae3Vtf/AecgGFy4
RdWpgY8brS8zIi1UPhK1yw2x/T1ho0d1tLOeNvvmadtc62/wdCgdvAUhMjr4cX14OCrQ5fNT4J4U
bS0PqZZpW4b68nwckZcormKjtwfMHGn1l1QKIOxVOhj5R5WX/zmtLVOW05Y1uAnTJhBMpYBqJAEX
RNjtyL9JZK3BAfR+LEByJBvWELc6Uj0SiIGWFgf1UFn7FpxYB1gM97TNsxN32MYBT2lGWpX1Yb2a
V32XqH/RR41m7TrAILLu633n1bHQEzIn8OtXlD5eNoKxn8LT+eIgZdvNFl/33vD+INK5FYFCiBhG
L426rn8talbL1zW52MjyXlOra9BMtVsnFjEuQizS3rpsqaXfnZm4nCiCEurqWtVJpgh7J9fltVHI
RAXOg8H3aFlRSZ0VNkqiLvaUNTmMxpZWbjRh+dHNY3MmwUsnGK4y+w9WEEq7mnMhBQ7rBy+AKxhm
KrknrD2GNAgL2GPVUyb+dhTAGaEbWLHTa0HxV314NOzHO5dGfRIlBz4TQMCuuyik98+lcgoKTadw
5pvcsBBv5HYM9Ekde+p6837cH0u2YY0e1yX0SL9v+4IYXDkyLpHxo//7k2TSUcwnMi8ZcG64mrsZ
FmumOkX5m4PAbohD1JrG//WbnFmukXOYVr+WqtJOkkc5+S2DYY2+M70poA+DakUbNAQcnOdqZhOD
Axy4AzPeBlW/N3WNGESj67nJKM4F5LNC66g/lvnd4gHWIs0TuorUehSTRwDlYLQ5aNpguC0FcYmr
4bBuqFvEZuuSo93nw+3997ryTmpVbcBUvzCq4/X0b068K0GKdr5WiMJtY3aWNo7UDa5fiQvWAlrh
NObnZs/T3WeNBC8fIP2ToI9UDldi4D6H1Q6klHFtPJCb66IXTFjCrprpG+HPQ2dXVIeniMlEjOBX
lL/GriejWlfWS3+xeOEq8Sn1gwpzjjKi87uG0+clN8P8wIH2FTTqzAZTIESZQOrozYAKoCtrKXXW
IAwcfx4uhaJRfas8OyBsTbxxYqvnwG1wuxCiQcFva5fDtgUJNmQhFFXwup4M5MwYgRxWdU9qFkyv
IIswyoKoGEu3aRSQdAUH4Bt+34cd3BxZJyP5tkHuNvbrSF81L2UuJ5NTqRt9Nwtlq5o5JW4zRsmU
3E5lKOn8tX8HfgJ8H3hi9rPS6NV1z+T5p4RJ115ejCzDamSKAG8Z3XrNXl2orYrpo/1BoX1MsoON
UGeuuW2Kzlnwg6+AUnDPOjuniPsf8aO14FpqGcB7/wGOJhrtUCidWYAXFSHDjUivGip/ojtkNPX6
RSTc4LxRt1WCB/V78HgoFGpdcGX77r6m3UG3XBKs6qt/LvmbhgbOHIOL/ZvcRR/O//iHFJLwuXFh
p6GNXxzS7TGROtzcxTackO0mEzZ5bwYLo4Yr/dudn6K0yQrSQugacd7ek0AAyqZtuHFbIQ8auR1S
RSDqeDTpjgkaz6Xc2lCjNV1ZLRHGt1/E8GUJaRLVC4nhtnHujZTiu7hEk+jziSda8cKIs1mg2Zm/
q95Ll8yrUa+cFTNbc6ZFsy4SvxogVxvx5bE+JGfPYxpjHgjAS8OQ/Zed14EYXA30V0X7sa/jR8zZ
YaPwEYAiPrBNQ3Q61ZeI/XPYZG1iXJ4lWAfnFLR6ZFWeuubi0ltk8yLfpdbRdI2I7sFrUsKHIz//
FRMWPDXaUAvICd7XBHjnjJZzr9gdTWla3Sq5SXIz/xnrD9TXcWK07eYQgocWxiyGoPirYD5914L3
g27+bZkBOj73aRGNTzRsWfH0ehoa/d0B1+oU95uLOQUdcqjzB9JEU2OPuXiemNJ8SoTGRc405o2J
7cmhCMyERP1GOZblUjCh+nzSBrB8eclAL/mqVa9N1mQQgTvE8obgiXhh9SMVD0f1022fx1CZi4oo
f5dbjMxqU6hxi0tX28ZM7utCVwpLOUSFseSONlOeqyKkDpF4LomumKbpBFlw9eHAi4FpljccVpi/
Xz2luqf4+f9MMswY/49ESl0QXm76FHxceqxtX8co2DD+iE1plGZAc7/hUTuhm36Fl78vXO5zbNLK
LRctFAk3ygFgtOx3pQCVI4fkDelDUyH9FFdO/i/edrNp/hhSgxC+YFMCeIu5UoJqFQCebhIEQjpP
YRGkR/qygGL7PglySkHMkIpI1HL7iwDLsftwkeAsIkzPAR/jxHh+KloCg+L70B2iFFvURNKVxqcX
pRhASNZkOHijrknNJ2BvTx7khq7+683KaJ7oEiG0sh2L5oh2z1165N5FT8AbyV/eNEioaDPeZmEW
Q9LoelRsOgFE06ZcHjmhobFlIBXHjQj3dghFzM3T3ZlVwVpdQQhXid0uZm+vJXcSVhNVzWEU4unm
IorD2KWMHqe7pti/6tT+mtTRKTlnmUTXj2eHbdYFUqg8NlolycvrVCUy8rqUzahzG/R2OGihT7K7
U02WnvvZfsMu2S07Q4x7r4PADs1XajQo/9fdUn3RvM+GhuIHFEizfqor+lK/p/pnGspZqjGNQSyH
cRnczJ9+ggQstfLuT938vuvnc7lzgqo9trm4nz1tJsbVJgN70vay2iIDn9SFsRLVR7MAC3zvFoUr
h42PQ+DEqAEoJEHlDoczFtAghkJNl6KqqICRTznMr42VgSVtqI/vK/ZAFTFRI2sC7bQflQeGkicY
wmDcdvs3XoQYtcG6pZ2xhjwij+k88RqHaRGw/LkR61aM/hGDW356CWPBsXH0kkr2VJ30saarASgO
fMeie+T3kOBVHXj3v6DoQ735+6qVnve0qQt6OiMJyVXVTUltgihE384sMiaX1jIQhCfB3KfZweH9
G4V2gpwE0gk+ir6bRunir2KtNKf8P0Vqqad6vQBWQdUTF/ww7mOU0e0WwkdYEtYohqfjjvQPStJ5
dMh8Sw/CsSutFY8LBgv8E0k+t4l/jij1jzQvhla62VZeJWTROOj+bzzMhfPC91Pd3VhId/60BsWH
GcwMQHWnx80DljQjPJRRfddia0Qp4OHpbUVAVvH35cvp9BKGyf8CzEPg+h0PzVAb0qt5LwbrdQ+c
CmbhkgnEpmMoBouObA7SMBHnB5iNZjbo0d/QYC7kXlH8JtSPoco1qRhjLm/xJXeDrkx+fWcFNDHN
0S1FhHlAXkcTSpdjst7op1I10VCDAQpOwjj+HKKiMoJVvz+mlwvIOOtSFSC8/3+NQeu4jqrzX0tS
q9apV0KRjJR+n7NBvDal0GC/UR6My6UV6IfWRs5p5yuBwQYYnXC0z7FfYfzaKtx59XBHzGTF0Y78
FXDYOMuAteHbrf0oAjDkHMb95gUilKJlMC0pQ3PkHDT0sIbbTwX5shAvwv8NWn6Yes7RwVsJ7a0Y
tx6QfwY2D/+FF5TjOpvelUYkbXT/m7yycH+DrSVOHqkZ/8pgC/8xrmuk31iffUW2+DULskhlEkBI
GYSjuHuelRNoUe0tE7mH0i8DE894aJo5xlMLCChwFbfEAUF9DVG+HC5ioGHdQvmPV8863jI+oO4v
WlK+5LGl5KZiJfIHu+V92VH5cJkR7ir/nxCnOjCAIi+2vwoWze2WfJtdbn5rsj72uBC/2azVmh8B
2wBo7bB6uWQdixwMXTa3Mo4t/yaeCuJbKmeDmbLrYCvqmnNzxtJTELAzUjwrk64pV9h4T1A6E9WL
vG0f9C0xA2Yr1A6sXVvRQNgpQsQCbPd9s1Eq1N9uwHmWh0h1zUTeIMunJ15ugm3rswh3nhT6Uwk/
qMzMb29zO9QHf0dhPt9jWd1FkJ+lQ4Qp10rx49Y8pJcOymFLqj/WRebQIYVVYNep580iGnTvYKvI
hhksGM54lYHSBC6ATZaEdJnq5vzRcHqvl8ayk0JkO7aj+LC7x5oqBQLtakRpdejCuvmREmZImQeL
MRoTN0CXc7f856HcmQvMQIi0uaaXjfWYCfLy06KaXSyQ80UERRYJJiqHeBj8f7nDJ6f8XTF5tmO+
knZVFGr5A9EhNlJXBFXtCQFh9lEOuCuZEuSQUg0eyg65q+YyybZ+I48+3jC1a4Ao+llMeCcm5z1/
uBJc4D8GIdHiGR4jqd3dV2k4dK/G0McTkefFOfMWoO98NzZOMNyyKYZCMdOkTVBGBYSHCOJZBCBM
MBwfyY7V2IbyhdbuvHascJqt3OWBqDiJ0Hplwl8w8uED07z2SGTOpj6RNc4MAJPOhyYeJfVEzrDI
5IO2N0SvVxjQ0OA0U37d+I01QNxUxTCAT2wnk3xPwmNxmarvSy3i9bvV6YuZh+GbHuYASfHib52q
vm3QvWyioGuutZ1gzyJXxxx4CmcUTHToB1451NEwN8kjIB/aaXkYpWMwTd8GJwpZhE0WmBChwWNS
CU3msu9MJSFtkrYvnp67BTkg39dQTKDCZQYObbE/8QTf/fhJsMCZiOFwoLv/YWVKr6aZlenNhJRn
28qdLJxWiomacu057bFZt+xQWfvaq0tzYDDBG0DQY+YZoATNGAOdS/UWqZqBIwcpFfvycHxgHzs7
eXh36ZuOH9JeWlt0S8XpH8rF/s0cEojlYCdnZqHeHQGY3PbKIMCPW9u+ZOaxvzBWrmavIXEqgpHD
xTsIyZ3/vitW7j2cdtg5KS8h7zvxGOTtEDIzhVQZli0GOh8DUza/Hw2IQ/BqiFKuNWSJ8kQg4gTw
xbQL/zlWn7EKcKKNIW52UKan5o8Er7eZ7bw/wfC6+j1F8F+JFSusd+vxHuviu5cVJMC6reMVNQhh
GWWNss2tHIFkkeNgsy4Eyb0prdQr/RkKFtx/MnVePAoZ3dZ++zKa5LaBLJ187HacNmhiw7GV1ltf
4/PsU+10Z5E68kKJeedinQ6msrPABn879WXfpT5bA61XdhU3OSjhvSnkl705d1uelw0cUakA+H8M
qujTLOc3t6uMv4TUMHAV0Tej31rEVEbkgnfTQM10S59lduWwtur/WlWBJvZG7CzQP6gHz4ZrgV11
OiTXbknS5/mroyO2dlE875yJliRUWxEeU1f+IQ86vkf6V/Zhvcs6BMC8PNKOxiMt3yDkwYWnmCZa
0MWTFuOONlDAa9i07m5p3IFo4l6d+nYn1dacHY3o1e8kcClh0+lnONkUqdlltW6vzZHMWJbd9A5L
k5d6BrLnHZPZHW5Yl/U/mxEgsyvj+xdrgh86lSc+5nT0XDH64YxA20WUOzhgS84roL1NoAj9eZNH
qd0UNvTJD/4ROk23T15vs7IBs7ABTIupZiYjY/Mb2BkKcWnOxX/Sh4ab1ZAZvxPLPG5GKUBYxDV2
4GKQsNpL9zbXlBce5gQSv9jQzjVD4MTdzk3dFW+TOotNycGrOyatINixVpqjLOmIiRqyGrajRE3K
rhriZTp7aj11x2eZNuL1C2kpyEFEYz3x2162ZW0DmrQ2XuFwLL+G8/De//fgOYmfijA7CfKXx/Kk
pRzvQH52A5Gm1kH/xJK792BwlbGyfChAby2q5C0laV0cvTPNafWkAognorLimq8s/Qn9e02VVPaE
QGzX3hTumb8ZPjuCI+VTJTOOoXfdgRgNL81SQe6FQdhOuk4qB/SB3bF3lIpgZGvfxUMSc9h4p1t2
gKNoCvDZoPNS6FiKdmAcHiy/wmPdqWK5K8sZN1rYijm61XRQqzo0upgvwamoIvFqAfAylTOMPcyk
qgF6gqfy0thqzHUpvtZM6/ZxxwOBRQC5UpWxYuVCDaBVWmjviminFBLDRDmGMAivY+A9wo09GmPs
cMx1ddwz9PBT4vruT9xixqiYihguNg2/ZPhogcCpulf0fjYoOVpdIHHiDBiKY8rfZkHSfpEISA7B
8idhjGLOMUc+8y4r2z1OlfsDlJ1w56FCo3ZDvUOaQPotpvl5dp9eYX2VSHMdoZirVsWpZ6rWFKmS
AyqdCQtwY/ANI8mTzY481gmGPgyVcf9EvKyjdSuNh218uXYrfY8T3NMi781WuHJ/p7Dz/3j82ggj
jUeJnCIYXj9rtgKaSpCAo+xUvkUFGQnEHkiHJHATIqMFB+Cxev18CUZjzmrRMwck4/ptro+3L98L
9uBPFPZyuDfnIgQUd7I3Kp8COWspcaXMFt9Zem7I6HQljsVFTzz+qqPFKdo2+Tv0NDwskMvRDjBJ
milSPA2+lfwVs+hozl1vfXIS0DkzGhsa3AH8jGAcYJfYRVGVOLUgTju/oRfEyYijKFX991OYcRIp
/v+iqjdcvvestEeRyDPCdoQW1l4T0SKoC15cYATjr6T3pjRAvGcEh6d/tf7iT8e5rXZ/MrHu1Wlv
RXJFRz/iBdSSeoiQEQYJKTzhxD8oPoPU0MxgM6uOu//79/LvQ+PxWNDFWRrHrPKqXp/JJLs/msWP
ZfLM6W8B5gtjq26h35C+ribt/PIS01RJTt1Nk40g8AfSvqDuh0+8FeNxV/I27HjIrCYxybEdJo/M
RdLwKRloufJrTBR5mQ16vrg4hMNTJig6HgrAUAZjl6KQ6541MaAUOA0XKp/4v843Pwe6R2LTuBtQ
hJAmbvftjHcNBymemhenzax8YGq7/yHrmoGwdbTut0xsDcllRCOlS7SWyNb6pD/6fAoI39mlWW0H
/XoqgfpeQMRtnk/nZ2amb21BNKIlLFWgoobBSzV3vq9qmPEhSwE5J16Od1JI7mXzBXOonqw8/zBA
/ojWPondl+CtTprOTLl0kdp5I4KIieo0EokYDRK4648VBMduxVlgYNnKF7q83dWbDsPXCZ4JU+L0
ZJxLvNC/i56ngR0bNP49ptnncOhwCrzYsT5NzFCzLHviXcMdGNLQqlyiALjAXwL2j87EF5CukfDU
NyvgFUAnSvi+iNSemxjH4gYFDw1LKYtuAdIYA2auSNRNiBWNf9U9db2hwNHAkLR50KLiB1yUw+Vq
poF7cJ38LWsySPGKZyjHiX6/8e73HWoHHF6LoTH5CHeptkY1RS0wxyim3mazvVC11YY5RpynjOMn
03aiLUdTOXNBd9sI/REeyuFxeWb2e+YDK7nkOkL8WpeK43HsZyWt01W3mkUN6XXnjbaonYCLHB6D
vPBxBXx+otLHbmtEamxcE9CHVXL0O+6++sLeoQYsFnJ7nnX3wONSSJGwOnSRVqKW0C3ARo6klJiO
yx8t6rBMX/zkU/T1DWxkq/TdVQM0x6ocm+zKOoLpggJxvD5L/GSh9ZajoSqj7giNXYzrtwys5YGI
dQgRU7W8het2l0zm3jNRfwuwyzFnvr6hEDl6kTMsuJRraZBuGrL57HXmJNzYeErrYrwQFhSk3qZm
Q0PK65P1tkEqyutuwsu02VN7eanx+AeALTSqGmWE23chIq7dlSsAKMRxQ/D/xrZ7xiZu1V2Y3qzU
pZ7WeH/vsy4mbt7XOusX/0OkonBHXdiStfAf8M3hpN6o/QPLBbQl6DYNG0JOuOH9aMOHmAOhcz5K
C8jhUjeAmSI+lodY6T2Z1y2nC/SriMFhVyyaC2xjFv3PVmcgrPFxPGMUgGPHwFKTWvYs5ZEZqdxm
6a+GyWgiFTGbRVkhaj0ik5nY0cGWIB5D+x9y9xL+qOsNfs1hekOLCuygMLKh+Yujy82977zykJfm
tH9Ie7L3na1GdQJnJ0upX2QE6WKuAbr68Z5mlSLlEzrUOOFyV//Y2MVhvvj8zxu21TPY4gy6uQNS
AzJFGHEGPOZ9GQN4JYgzob31o0HfEbDIe2KNE27IL87PzeJNUuuqh5yC83ddvGj2ZKKlpDzPhzvn
x8wuRa6bJyTs7l7JMlIZ55fg9qByuAjCfw6wHPlzW2xFP3wMtGIObJaJ7zzJcwqMss5PjYBlNI8n
pLffPS22/gyrYRv31b9nOK+p7yExBwS7gg6H+c49y/LzfgoEMldMSbenJypWAM+83dL0sI8dT/+4
lcSbYoNiMFnIwFAd2C05KPAPzjbgHDsjBW1lTBplm4/I5AwWfrxfzXwegHcPluvwBpr9b0gG7zFT
udhPFlYCCiVY8RE78ef3xelytPB6078/ZWW9qPc6x/MCb9zayUbJOApNTlmMALI60irFtsmP5k6N
aSUU5b4qY8HnEHLWQlaQdENd7EmWCiwGndlRhyYxVSUUHuEBGjmhLPOO4o8jdrN1LT74Ukp527EF
pfCNqWXqwyu//BKzHf0VFX3BPLkKi1OR5S4w3c85gYkS3xvZpO+xrrO2DFcrodb8cpFjwZRvOkKP
KiAEZJc87gJeBREf/OtdONCOkq/OJ7ITMc2a/3QuZK1fc18WWYpEwTcf7QS7NgOKaIqHdUvCvfsU
ytLGKXSg6ubgmyblQ5p8ctNNno6Dc1Z6aUt2ftn2r6vNcfpZxhH4sXXoq4PASZxXuYfgH4wA2Hus
/Zcdf0zqR0FXSVC4JlJgDZL/vxkY1bWeRKkwKXxHrV3OxgjenC6UFCWn3eu4RFyW6rXkPg11+m1B
fXYcIIdd5IBsLx49pdKiILv5ZQoZ9Qgx/lPvYgNbUrnWy0W+jyyj17HgHXKDT0SuB5RfVnSVxryb
TwlzWeZPbGPdXuLoiNT2Na1LUYGNFQWxVnOAifBFGtzOJez3huLu7n6IJbaaMNc+9PNCrNGqzh+j
ueztXMEGaj4Nfj4PGMtWRlQeWEJ8XmlAqNgOuaF/sRdr2VlusCFWh1O0t3SNqWm1/IChaxxCUk3L
tPRn/jCA3Y0luwcyvv3WInTn7FA/Bjy8dChYg/kEncLr8R7j49sIi03+zLKeU9i+HWhJ65jBjsCH
PRh00hlmF5tgJVQ68+g5Biz4pUD1pWuWi5lBgpuEVw0kfjho9rwcyXkNx+luGUfPCd6fCz0k5Mc3
c4lXdVHfrIlsfnLkFmDf2v0i8kGRrMKmKrWCRwWYiSQt8SUScmNp8WCPldN2BK1x1oOahHQGVu9w
j7qk32iWtjVLXNVDzIA4GpGppk3K8zmj9ZiSoZkR5zsmS05I/UvowTn7SNoRkotRibyf58cV552e
WmtbY8u7S3aBRmVZOT/ZTnOQxatc3WFJCWvFXWobVEAVMaFdw1ucb91G6qobNirYxSkmOPCGeyyx
7XOXEZfRiTg6g6rp4WURl5W6L+Ukmc+TkAkBWdEIm0XPuHbT18j7XaniC+lLx5hnT92G0VbvJvb9
unQBAl2X/j5MY+SSIRJFO8W7y182a/lkfV8loDLAipHo2l1XcHxQ5aCaKR7IPgbfW2SKcWJYVGQ/
R+V2+oJOpaTkCBk14baGs/phcmbjFL/OosLiRTKhzVprjPO2PGgf5P+Oc+ht+5vqXHKp+jA3w7ZV
YG04CeWgCIdjNA+tmZj0SQ+UY1O1cSR+Wz92Cp7OqkNSlaFQLLbIOdTvTpKZwLoEgklKrGlKqm+G
wWqBHGZUxaXe1wCRQk70x18ZVHDpmdS/qPoL2Mb63fJ2uGIqxNNxbrTdGZlG9lA8BLDyW+mjKftK
zk3LIcQKvEfMjopBAz6Hr2BK+0zXQuIf9NEC6oT3MkrsqPXEB3jnb5AepO+JBlY9ZFxKDyAb24Cv
0d/tFgi7JBV6F7lXylOD0ybCiy59vFjU3Qzj6IxefRYs/kVgZ21N+i6LBPvP5ETMyldGk4n9CxUg
AdfJWQ3nhj6ku/N+3fJ7FZwWaEgnm3Ru0Qkj5WazTLW3D7f4pitG44l6nOG4fGHEiPala9Jazq05
bQ1QxTqp9f+xgF0ERDR2KbcsjTAUGhESNvto3IsGEqq1tkK6hiaWO5FrwFM2JXXRxW+CrvS68b2/
QRFQydpfhevdeMkPRg4/6g+T0MHLxkeMkICz7X8Riln8KKRWkSNA6S+SEFqvaRRh/aXnQIfKgLz9
czBwc2EGDxTWaTY6k3hQbkM1o3ZIft4t3gWtcIHspxkxcGlQN8P63QlUNSrf9UWckU6g90xrl9sR
I/tEUI6wuWDB2tz5zd7A2ybFy8pHREDM4dw/f80BBFb0jJL9xHz1wrl/mEC6RRAsRIccbXFiQMSZ
5bJaejbpcsRpzi6cjmyMDIGC/c9kCz82EeYq+Ska1ObqwFRkTS6LA5QK0KaltsaQEoeHuHajvXwb
fGb6koO29J/gwXAU1nPkyc0RKYP7XHRr3bo5W16gnDy7yAaouQqJVlDFgNM1cTmLQY0dGxWyFGtv
DFM8OKOBIorjssjZjBqoGb/UwCVr81UB+FEqg9TEGRKMWMzSJfVekVScqzU4R8lLO1GCBwhxJKLm
9RpHhMMw5u/9LLet3gE7rmXVfxM67mNSD68quKUBweIlAY2vzc/FeUqSH3Sg6LPCC7OyrjuvNyXR
mEFAqhllZ8XBl+uPVqrad3lzONkgPfh7a2VHZnbB8jGE03LRV2B1lAiZ2aosipGivzZayLm/7XSf
nOlhijGWAxQ9tI19PScOu4GaD5gVzuE4LIFSC0rAWZtlTpmQ+fAyn6oclk0+cMM5LVCsICYFTSoo
6gvcksHo7+nNR094F0IY+tKgHcvorw2bs2nAGqyI3BaKOgF9Mv4B4pELdFkAnXAJWHB6os2XFsJS
ujdqrcPgH9q8k3utLSIJJdcdhJPJBiLKkWiNIawG+TkM8QpaYJqnQ4FDtO8r0Wgl7IBdWiS36mEs
z5LaTuCzrEud/cU0YbXiarZELDxh4N5Qedy1FmSDPpWZ5oTITq6wu16HQQJBKAEjxaSyMBRQnkog
PmgVIQsPm2ga3ouZVS8nJH1NEA0V63MkkTvFCW2rt8pfexxWAbp2+9sMXqXbrnUfbu9dvqXs9mCK
ioKaYejAhQbBIx+ulW0Bo/KuPNj8TnFaKyNsz8orEhDjeInqMg8Z8dgKCPAURJXnS+2PnPzIvfM6
WzB39dA8qtv6B5jV2Ely3L/q0HoCYQMYgDQEEIhBdRRK1qcbYKZiWmfz3lxTODvgJ4S4FjKSvgKi
25pgaRHS9JiYamV2pFEoybHq6+QnLvkQwnlP7sixYuzDE1wHwBB+jy31AOMJljYVGQ8js3LACF4B
LYnNDteSSk0H1QXVyAiVHMwzo1o/UvVN6AeNrnx6i5cm9aXbgv2L8paVumbGVabpoDKAjBqJ8AEN
L/D+H5/vW9TVGqHE6QDiMb+YvavaBSxoaPbNkdN1i+Sg0YbDbyd3SIvYaL2de5K1T2dVgvajWeGw
MFRBfN2fy/xKr1Xbx7s02CqYF5wMCzJrX4yGBFtHiIKlDCw4WD9+4hK0lz1NPFTv378+t7Fvob92
xm9f6Hlk5/AjU39LwZMu0PLWnAZ0XkQ6iwRA1HfjUJLWW565Uyzj6Ccxix3728gh1usaq6lFD+6K
lmh8oP0foL1PBpePKWGPcOnLr1mPChbCYcyOc4+qtDsizBB+x/EGcwERnyNpkivndFnT+mWAt26S
7cCCNv6HNmpVtOw5htTrH0GVzXEpthIm+FXux5KCC3UtLzgQcXhGKivdc1rGb6DpuhsD8bRvJT+r
VFBpRthXfLc5S8JdiWiP7YqasK4Y0zzSaQYUvqB5P0AAbeBhLEMJ+HaW56WNqApCGDNwWhXyDlSL
227cCr2ezSDC8HKoxvzrlJ91NabU2hW7NbbipoUJlMrxBy4UVmmtk2t2C09eSBZNGb4Z9atK6/Py
Qre6ZgpIfzrxQZXPiDmtoDM5a/MeZWtoavTloX19T9TR652uKRfDPNo3N3z9w9DLsmDu7eLk6Kvj
l2vPO3jMrXvbXjBpsEOrTLtP5sSys1GmYlRjgrlbENtRcgNqtqisOv/ysmE3cLGFQKMc0YXL8aJw
jdM4Gv1Wl8+gl7QMCSaWEYE7RWJ0PXus+da2me4AKfb3FAwrgOyAfJ1PABLYig3KOHR594jX9sZm
WSaSCVze1Z/hyI/TFcBPVUS76hupeun4tjILh06AXtw9qoFob8vTd3+0Qk3VCMt+C5LRy+5LHHz5
9xNoL4zzxgvQuV2wGLp5ngCMm4j/BRUIFv60wm9D6uZn3GN0zxTdkdSjoVmOCxlNi+1+6WEkMjmH
U7nFZdPvBset4YPgyMXMqZYsSf+YwQjESr0ay+9ZRfD7mg+l7dXbMKQjLqyRhbV+5KpvJXfVyIL2
dzT5odFvz8BF6J84P1bpKELNAt2V0KTP1byFARiFl3C1KS813R6BpjCH4r9wy+AxL8CPJjNhPE7x
Pb/XZH48q3hDVJ8Gql4J8KHLykyfuz6lpVWst3pK5y2Rg5VDz+Z1Ne52ZDWnqdR29tvAtQyrVW3E
5YdgUuRtsjvLKIujQRZsbn61WpI6Lb6bkD4rVs8B8HLRA1lw2U+y1OA01C2+y92VakCq5ZvDnD2u
vQBSrMnoRV6PK6pcL3yCBHD//o2WhhLJwJo1sU9/8ZFJhLrPEa2bmXz5V1jbV7QtZLof2jIeyKxN
9fVm4dZ4GoYDPyl+aw++62MHcLfoJCGyZOyD1S9lr9Ws42UB5JAOIpRqTlLZzDUtEtsgp8vgqLoY
CI8SfBUv6UVU9eeaiSiAH2SLoI4LWbZ+Q08uY0lnhRidYxP8WpxdYZIgPDlMlb5ThZdWtDf82Inb
o3hCEzWrtL6IIC/gtAlhZayeCeVqox9ec3NsQNQ4VrdJNF1nVJcpgO8+UQMV+OsvsDeleCoeUWdt
orwFNyatNKMS2YGGlxKUXCwHbTBNnMq2ZXUyAKsEWb4mwNNju0J7kM7hwzbwSWpvSyg++U7/6gYo
pLavoG5WIXmngk/0md+5nxSKkRaXt+6RfSA35d0YyTHd5tBS24kz+L5BfaxtEMrfVnx0aXPEVt5i
u8pd23DUsM8zfzWVeWGeGZWENn6eNunn+gUsj5z6YwEOKCDIPwydjSacMqZ8IFGx1jV5wnF8IA3Z
7sYJa06np3yzcXthxQp2d7pxiWJkLtTIXWGbCIdh8fN6B4sd+pDludfb7JqU+mkJ76bvjEy0Uf8o
fgDDypecaV/1bCaJQTggd888U3h++q9TxyB1cQiMW+3pVEo5LAOtQiLVDji5o9g3UjAstsxO0/kM
0zvbzrKiPGNa0Ba/gQql8tktE47zP3iEhbl4Vfb9ajiYiczQlLpLwTIQNxB3T+aUDqol43SDgIzk
WvdGnZQed8j7mm8wWQdyQqdci6iKjqPxNtCDt6/bmwWhUuHt6kd96Ffev4i9ka4Bgi4GgUAE7P67
ugn6Odg866+bndEuOUM/rQVI6Ro/IgNKg9IfMp7HGkpB3RGwJWLJFxGpdqkLjrzcVkTcDOyrDmiq
21F+YsqMiYINoNyhQglkbnfpGbS8TbSRFH7WeTZvWxtlBIrEF4q2iCdo41TF2sUl5Rs24Jduckqu
cv5DObaUJdciEehU+nfhZeC6LdTA8b0CwNeaB6lwtE9hjst3ZBC2mHNVk9LA5Cklxj80NnXJfmtc
wnpTlVTL5/nG3rziRSqKiLpUsVOc6vU3Ax1FSK9ZYfWkEZdgPJ2KHV7awuXGQCku06ODY59tezUp
fLheod1/wl7Nh9jXQga08L2hlUPNEKj1cSfZEZzTyzkIv49G8O/z8nT0iMn6PuBoiJRa0SLGzpXL
KjgZl7/3l7nJ3XORXRQvu5f1MxJuaznGQdBf2atVMhWNo7fpJqYkgjnC0a9mhca43GnE7i5gC0Cw
dNW4Dl0rU2R/p5Z7Fwyeems7PJG1YciaET6f9ap4aPyaPdUCfWhLSSAyF78qsRpPhZoBHmjYBsGK
K+OM0PDUs/XOpkAhVrMNwKTPGTbDwy/NQD/SUt1HdoK75T1P4waMEdWS2FX2wpY88xZzt/TTOalG
geO2v9eFJQ7cYtYr9jU4UBry7k0upbmDtWv6C0V6U6XJbhBvX35SjgYBBomgJOY3CppLS0W9WM+8
vOEMrUqdEpGbMZgHqLh4W8he740cDoKbCfL4sebK1Yze6s2nGUQ5DQxW4gKx6Ot8TT443tcCFDkT
lGFRXdm1mnEgAVWKdVveeY8XO7hGlZQmTdE4RTILMoMLf1DVTr1XGtxtFceso27d4Ran7atemDUB
9Din9/kc1XdMnQiQKSB1Nc03hlJOsY1t4eyA/h3z6yW5gs5Whyp4GEO7CuGgAG1d2LI8mVUHNyGY
Yprxj7Dxuj8LpzOXrh+mM9GKuXpj69xOqoflkhc+PSnBxGkPg/qyaQBSF3NrQlGkH+VJklnHt9O3
TV39zIQPm4LydD1+D4lEHk7ZIKdapcJXGhV/ukTgkMOqXKRleKUN2GVXf32zUMDnkKPyWMd60J7J
Uj32v9ld2hI0oEn3DQNmbMzwOUmbBLfbPwN9xDoCleebL9qh/spDzy4q7EJAzmYg/dZWvCG99niT
8Rjk6Epk6nJ16FWy3Z2j56IygMVlVO5oIED2+wKmbsKPvnfzY/1+Zhsbpe/BN7fkuV0CHMs4Tcja
c3nzleT/TvJl8VZlZlIXUIejJer0jogOuOqpb4UD9gaZ7lQugxB9fqWhfmjDhGYWXMsX+jj2U0TO
tUO7AAMm+YHQcm18QX6S9sRImRyBNieVMCM6lKVMgLJZEa1nc25v6Jf4KSzqW50fXEahckRsv3xA
o2LYBtWEJbnDMX5SJR+8uibXkP4hPMucFQF0bh2YCRt6zezUlBs6Q+DzjJveeTGpvauxbQmd3uMu
l3389KeAoVeGOEvCM66nKh5SZA24hF6FZgSYyTYrIuiZT8WGr9F30FE6i3/QpbZ6o5WvRVKKcRao
zbHy+ENuU7RlxWR3/XI7AwXRVgRP1KmkRGtemDMtTdh20/IJqFk/DQA1pZNXL6zmqUYrF8342uzy
vRSZMew+Yy4iDCiRkDTJqU0QQYIT9XFeB1hk9cmPbICis0lWYPCqcVJkauR48p2qn7yE0thb74oB
/54w0liYgNs/r+ra49qlfR1V0oPoskEgsoqsRd4jxHajFDGa/cYyh9SM2k9HWFwgLIbdSViOI1Go
3u7NYa4gtocfmWOfdTIEZJxmaUtrcHplOSlnjs/APmLhDgOnSRHmxn61xiTGzh4aXYe5v1tQNMJP
BrJmh3Cz6nivmypIsjUvWSP2sqp9TFXHFch5jF8AlhgHyc2hzhiEiKHEBm2EeZEL6SDH2sMO2LBl
pN4zaXfQrJk4ihqPVftoHZOedUBvNH6oOXx0rASL1YeIh2DNdqxKZMI33SwBo5YLcYPfiyEVxSBK
pZHAZ0qztMG5KEOb/KXQjXGbNomzh/wYlgQjPRay9ctAx/47aLvGRid6YUH3SYMWlG6Fqe4ZSd9C
PgKJQZ/iAmO+Lx9a0Ra1E1UlN25qJ0itqYOeCC5OeRkzZLJBluGiCAXLf1qTPCwzqXV1+vLeOGLb
0yGd9wo2UjcER0Owbwfq17Xgui8refeu7G6vamVAqFN+2dGCKXd5sXt6x0j3oAl4X2rNXH+5PSQ+
jAhr+2JvOgnubm/a28DApb+WJBTlt7Xyt9Yr8rU4XDBoNDUyu6vtlpPgFE090X7vY6uGMTfU9rMD
0yvh0wjH5dmKW3I4SKgDnriGC9BAmPKzbYjCbWDOcClmZps82foJni0ZO4gwa5RWp0Dt5skVBo4K
bztAeQRzk5p2SmC7gRYi8ApxaivYRn0MqxFf0tD5Pjp2Lxe6emEzBP8x/GUXbM8eBGpxfEvLI5qH
0BkVN+xUKBqwDA975dYVk+CJ9q4Hu67aMcoD2LmTLCsrSx4pKsaCLq5DTOa48JCi+ch55GZBk4ZF
eEApvnQDp2FZpo8zM3OoXgA/yOODnMvc1eolieGgzIqy/Jz1dDG8Jx0DuH0AY0Ov4OF1VzsMI9n+
906eiZV7PT+KapSqJSy04ZhD8JtHoEM+/fgsZrbpfFcaqY84qcyCAKQedh4YtLba35nnFla5588g
agR7WWc82voTJHacAEjm/snByUHXGcv2ZuaDAUqT5e9NpREOcTb/CJhn46u7R2tqTMkjQrNDoKVD
XLg0mlba5Pr9qGW4FGDAVS3ry6s/HJw0QZ//UMOow+nQf+6+5GYpeiwWeWtTRQ5YtcsLEwFHiDrh
adr8YAE3IT+oWjpbwx5R6bRqwHgHBPDnmMGSbWqimy9SMa3LI/5ZRsLKRWr0sejxA9HU21mXSJw0
pQu202vSztc5cY2IeOmEy16l1xixkgWPfsF+6O+kYHb759WqTjt9r6eJbf7+FjOm7ZLN82iPoffF
tytZH3hv6egHSHqFk2gvv7eY3sYfetRqO7+HTAKoTgG4tZ3Mo7npp4+Rr7/iKHnDBJW7Z5n6IbeE
ia9P88yABG6EGQkmc5Wxxib7kVXhmtEA5o4h1hAr4GDZ6V2VkBTUT7eC3wnZQsuedCioOKEMaLPd
UrvdeeX0/nqsALaMNnfAXcLQBYX9LQdXin33NSq024AZqX20XZ6bY6VMUKnARN9DYva/EEWakUjh
RJl+O8BGK7W1wdzci0vHIe3LTxx8CnHJ2NBIvf65TKfS993GYD5fUzc4fQTs+Ev5tXtG9NshzTkW
L2MiqNS2l0aKvHEYNvOnAu4mGE7eb7+DzMfNS8dunBUFnQdLVZOZa2m5mYoZDT6ggIJ58TPrkAqw
InloR+dyNQJDPfIH+oS/tSFcaqXmfgi23RbESJRFg4luOHI1MlcgJK8q9caJqVhALleR4sDkIc3+
gaHCVUQ3b2tUUoYx5EMC/CzPynIKP8SRZA++oICOfbe3SkLmu/8YHxmezTJH6uWj/Rr6aH15ea+5
uIAimRl5wFsQoRu+tRn9Bc2Tsn9HDgxS54KiDdCbR6wC4AnvcimxMpoyt3Fi2SNn7D0f9n3ZS82x
VnJiKblPdhGbjZaySBsvaJjZ11KzWcvoCEwoC8R3KqAaLct2T96L1nZXkBDtkueyT60Nmbrfp+ad
o/euIICxFowQidGUBls0HwmAV0Z4quqI0CFG8croK+B4JsvYswpYpZ1K9pT8XQsRtBgPW8uN7y9b
WQdOVOeAJ0RaplxF+sZO59Fo5NLeosxXSqzv75ux+bRuNM5ajseF3MBdD/noQJjROosg5oS1lWvk
QZGb3Glu0qsfvNa4TFQUEM7SJC/qw7V2LBTzvomSYiRhAMbxOOvn1y37KGO7b4xHt90ln0fX74/9
wrWF6019s16fBkRltfOXEAw0mzPq/g0ystbrUfQMrQwKF4aNDPtOWIj3BxZNFI96K8JCU+tLoKhE
U66nWs3apnaBO0O5EG1ZzBpUESZfW3AwggjV4GhBnx8nR0DghloOv5nXY/+NhKN/Htzru9ECiLkJ
zSsqFIto7Y832Mb4ZEv/6vKXUTaLkl0DK+4B5SfJjtXDQfmaLW3SiwXqf2UYyOlTkREDjKRqE+aC
QQXVCtzj+uREZxuWVGhc3Ezepp4+XdkOBlO4Leh6EFmWV1YWiikZVsoqyctJplcgR7pfthIRuTWR
FDun4Zb+bg4+wU8FU7Q+jaZtQCGazHhkEvCQi3I+eLZTY4MUOY66qGlTcQPgzhRsE1ZPPdrlSYbC
KVkNEH8wvme4qQdvKbIcXl6V89rLawYSkknLJwpeuV3pDiv+YExBwjz3IGg5c2Vi3YuEkI7wZuGy
Qjk9cHd7Ll5axkRRxKoPzDS3rJ3CdZwBlVb8yyqZ3y2KwAJh5XXm8/UXB32C3Bail4xmIy/nItEC
ySd1qPdiKHdvuyEEpek5nb2kfl+wxOEYkdPmHHC4u2HfOHjPQRTeVd+/iHrdmybfMlXQGl3TfFhT
ufNBZz8LajJMaatliC3KAzCNRbE6tbeeBSlkayu2BsFWj1SeVXCEbpefRRdRr3lJ1P4up5STifT3
u3P9hkeuwlheC7Si5LKfgmth3zAOXsaonnq1YAWbSgLymVhxsn8gRrf963FjRVRMSS8KvImfq4j/
qrPWsUaQbLG00fohmFZk5kxQGZ84OGhCxzJE34JjqXGzpb1pvGZaqn63xK8UVTUlMhGTz7CO/cq8
q14W9guafQRb0MoL2U3OAF1Yvp00EnrCpFmm+4QTtvFp23h/QkbJ/PqCTI0njbnPBJmSm3rTyAOC
aiPCVj60XoP3WKy76lofzmoCcyzr6YFqY5NDvckRWyYc1uom/VWxWl1n40IAb6anbbBJU9Rfz1I8
L2AoQhB441q4v/Jpre08gLYRSf40UWtIvxscmLLfzKr57HSf+q7VOtZbB8165DYmbDlPb1C3qI32
DC8A9QYqZEgOD2jBOgDRbWGeoUzRiBT7Dn4Pi3jKvt9XNS/YDSUO45nhz6lND0MnxDKgjWO0KfhW
Uq+Au1kvJ/PeOaFvirx0cpNsinEwi7wd8IKAibyr6uTCSMuPRpOWX2rDZujmg98uWsHub/y5wq4P
vpPFXwE4FWGV6MBTND172bUUdqzY7UdDp3Y4G4ELHpjLz4e+wQKfr2IS3bqJrtm2xg02mXzl9sKi
y/leo+01ztsLglkk1Q17tq8kSi5hEdRVFyAt7MhfcB0+9yK6aMkgECWvx/CGtGYD2WyIMuPIdBpx
icCnrUDJiA1/L2fvKv1NVEfVppbvKStRMr+UByGK1nCta33zSISl4ff52TB0/ZlV01o4VmHtZ8DU
p0R3XPuuzdcTVsQc98mb0iHmLw62HeU6oq4XHQIVh9l5Tbm2xy5hBBCTy09Ksrib4SOQf+oI11zM
IrDMHEZ+e3CFNtjCmd+QpmZWeyumelRrq0soAIM+lzYXWF6Qh6itP9/OZH8vxcq4Nzogn7/UagHr
JabKhM8lxORfQoyPXG9UyqHJzzqIpixDffjXh7uE4OMkJt/F3MKvBJc1wQkzBrwewfUcQWXSQYr5
CODvQ22G+UZyDKfVLI9nt4FRO7Ru/xoCxhPR4jVLWvoagc3xYndkQQha6Ey1+bXCUNfFIh4lWi87
QLF8HVzngrRaMztRx2lSD44URG0UbI2O788GMwEOTKspPOWoyLycNA876tVMZD/Vy7yAqq+t3rlB
wIi4DnZwhyENQS2aLTtvaJTk6YNn5uxY2MW9rxnYCPH+oNs5gC4H8efcwSh98wmVzCEE22NE6NN3
nDEYr7qtkQQEU1ZXoc0R8hyXxmyKZKXtfGzEzul3SitxDogsSeb7HrgtLnTCbwRnj0+BetNNK0mc
PQNPKn/NGmNkNA59r07DMSflya+WX+HDxh9DzHBoGcOn8rNl4w5cBXspiskYMgFGj+s7eX0DcQXS
zF6wcQYPeT//p/JhlDbfZ0Pa8NfWcYD2QsXfzp85olRJuil8Wz3HRvgpuIxS8ZBc/lNi0ZiFvW7u
MoN7it+HlC/fRCgjWI57RH0c3lRAz+4Y6WK+MdFjfj7k87SKID1P6UfyNIsAjb5IoKh7rrol9hMb
ZZ/qgbXH/61hd8K3MoMBLSiOR/mhkzCUcwmxWFUePWSL1eFwS6UW9I4paL1xFTYMwshUP8fc1wwI
B/gEF/XYb7ik6s1ycX/Nla3/pXntYspJWRtQJoL7+vo+h2jT8Uh9iKYLYy/b90v/DMeEWR/UAr8E
6JBAK321RyzNXr4UiSfrPAVuYfFmuPDmbgy5u/iT3XPk9yKA/IriWkTVHsnQ4nj1VNJqa2WZU9Ul
VuIMO811HdqNOLzNMH/PPNQv4snqPkxnO6aFSjiVx+fp8qbkvu6qh+FXThw65u1F3Zg/nM4gmaZP
diCC6SxQhaBaSPexwvTXL2FmjAY9o/RzyDj1IIwZJ6ipdzVVpH2O4qmz9Dcp36EhNJ608VNac/sJ
a0eqpDXghvKHr99OzHo+QosXBFI3XHxeVBzqRNjOstf3cHbaSPWyghIG38sg0Mf+b9OXjLmvUyMR
8nFj980ehjJWwpjm4PhFe6QwiBCYBfkiALe/i5wm4kHLV9r2QuSEUdHhnoS/aBFMbwh3NKpFvGYP
oOnYe2w0JVaEdU1D4avUK29z19pvWH3B7dH0KSFt9eEDfIH9aYC/Sn0Oq+XE6FvBwqcTEOXBbW9L
Hs3KXhmJk05KhEOAKpHiTA0WntnXfQpoU3ptt2sg8tSRH56f/yXkEQ1UBJUiEI3Ff1yHvlArN2Rk
G786oZmLHxiaUhfJfyqY9xP0diUYXunLuUh6jgpmw+7jxn9M2RuwkNyKeZfRyrC0TqhRhyiOxQXu
+MvTwndbzEoxP9hT2YwRC9ssIa7IsgW5APzo0g/bhfoRmx/J4IeWyhhu2YUqwX90RCr8GHG819Qw
pWjkrXyvWX9zMas5Hmt9qxorS5BhghrEtHfu/v/s07AbMKzUAKGwQ7kbZ8IrxE/nQvrDUyb0cU+x
dNUAiLCxAZ2PpdsAup0i3UlM+zjDBUkqhvF4vvg9QNFi+K0v7+5MkXXRUJd02DqgtXe6u4O/rose
ubJwz+ggxsWt4gNc/sjVNctx8l13h6QGX1loAHCC52YYBZkCYm0IkAe3jg5eFG1O5XrEOz3lcwXx
HIsszVjpmLVAxcuMHW+gn6uwPDKJd9rcncc8Q33DvQEcyn1/cyPtRb8GnivCL4V04qcxgcnExd+h
yaRMbImN0bJGovrD4tcbtBhIE6RqkTUJ9eucIrYQm5KBOKySV6BiJYvqjtIJ2bZdCQgQJMKE1KOX
APBd1hZ+Zt/+E016zuco/8GGCdQtiPJQ1TfBhXy0F9kkZeK4tugHtrw1c/0cCkUEGJP/UinZfmfU
l42DxaDZBCeb30s6CtsKJUWFIsPpuDy3LZ5knQPU7fa+lTF/S0EZk1ODApt1sg4CM+qBMxBpKfZB
WMMjIuABbxdFNla7OLigmPg1sOdANFr3LQLri8nkgNzX2VaEB+2dryjj/00XXDqZ22zxWPFzRquU
4jKweL574x9jDvmWZy0ZBqViqAKimGH1S4ixYj4gTCalSG/mMyywcadd7u6+j4SmTOSc0RJb6f+g
Rkim26HZ9j3VrdoNt3sStEtapcm7nL17AwOd9f6/zHviBoiL9611w+bchu5X70g8KZ7icVCvT5kG
WmqPTUwD8RAS2WsrGMh82ZoUkqzq0jlpx8FeMoxODgG3aFjPIKcSIjP/PDHGoYtxs84ku79ng+kJ
Li5STIADlqcM/lMaKN2YngyHe27OdHh7EDUS4Tbev05/TKSuq/XTuRU7qYWz8mJFWLKwSFYqWhvT
SSPuE3v/22RdFeHBbdu6f4o5DIZzyAgIy0vqBN8Us3P3sKiZb8ChRuvZ4P+7/3kTziZR5NsfKUgH
OpsByxs4ZIRcjA4kPLMgwI4W/84PvEx7XshSrE+4huaHf2p8T/VfScs4pYWOpL9BrbxeK2hZU9ty
HPBhN5Eih6Y7EwWwU9rS/h2FZMXEfqp+KChBjCDPs1QcqPvDe7wNv9DWBeJrDXaInTLytKsQ03fs
qj4n7c4XidbUjaltvS9KpyGULUzhvndnzOqnNHdZAITO/KNwDoDf2Da/5O7DlA0b//TIOK1uAqOB
ZRYLyr9ajZOc2diNUEj0w6LOagiMBpaByheWlKCROb4ekpLiZdvS3YsT3HNL7ccyEaVTxMtjveUH
/iwevSrymoFrLaB7Mya8hPiI2+oFDR6HdLV+47uxRIKXJ6ioZXe7ykv3fgMGLnkhb96YWvDV7sH7
VgGFjEhrj16POb/L9J10Z0vpkT8/upJFH608O/uPiP2E0sShVhgqY0YmOVVv0GnrPI2b5LyIPx7v
V520akM/JYJMmvjlQsOHkkA1NcpkkpOAK1q42mGkzzKiOIHRYehxiWmIyMXQHYn9GpDZDL1YMiZi
Xee6kOb45vmF3YTaFNqW+oK5FUmk7kbG7FbeSn4yuFBtGr0aPXzAx13JBKJyWl8e2aL5JLZkyuK4
UudKgeTSI1lHEU911OOKMHk9ATamUCckkeekas1TSjEsSj9iC9tQO3Lx/2s/VaURfdnTO51nM8mx
HQI7q4dsawhvxXIOKBiaULkR1h3OT7j1J/abh/hQWMJ3jNrWcIa+2gB70VKAyGH0x+VtEEggAHlo
Jnk3xZ1QdyeWY5a+hOojKFY+BIAV+ll1L1YKGTyPzmJR46dcgb+hG49ShgYx9ByADuJ2q99PpAIf
hDFm73E3yy4GnsmRte3ruEF8+RJDuzsKgeNOEbivZrdufHn2K9hgEFG4fNxanIFZDbWWd8pqORYW
Ki18DltazfQVczPj3iz1WZeJiNOZKNyWugmd4cCPLQP6V4/0j0E0ITv36Nq2920lOYQqmUL77eIC
LPgunBfvnPVPm71T4Y63eRDRWQgVJyb+TpQfvMMzNPlQxiIL0kF7CK94Us7dCztBl5fyh9D2o1fM
u3tiwv8wzb3SxBQz32qwTnMS5scyLnIzGeraUmVlQUMqD8RRt9ygMxIPQtncrduCD2n4lVuljFFf
ug/R9lTa/7h12EWtIBd7K+ucICe3KoPpClrr15ZkUmYlqeaMZR2rMujU/SWwPHZPh0EjXV8C6SsJ
PxpfIqZQLtcjbffhPYFQGny2jD9hgLAKD+O+YEA7r4LMgUwElq+nSBf2yCGubWpwgaa2Eycnhe1x
KzMPTCYSkqwTrLL4XV2Qn4Fsqncf6Z0UwhgEjHK7X3fbJ/K0AxiYtjMpzlzLo4uSLiD8il1ZTNbn
Rj9RnXR+xXx3SKuYv3D+nZ8JHrFl0gH5H/QSkA9JT7SOLY8OFNrhdYtOXLtdYaCSgQr0fphdj7du
hHmVhc3P4M09U5DBgnDiCSHXHoyEUsqOCJ1SchVQ4spfPPaXVFg37ZDKd6S+bBVc+TGZwilmZ0Fy
fIdo7aRtXuxEzi5wDM1aU4iPGeeBWvU2iW4mAW20ZkQTQtidpjaiMglVTBHBsh4vbQ94ocq6s2XM
dlluE9TV0zknViWL3Zsr06u3HuRXZwjKkk63NSMrcrXnwXEiiYonXVuxFHoYlXMTsOQmzbHUdR2z
CvWqr7Ucwcs8fxqFV1XCHT1OzDYD3OPxPoTcZLcAoaIdmOesqQ8efdkhSRVIEoO3t9NT2SpSykpE
ex+chCwvXIuzG+R/s35Dtqiz8mE8fP1/bI0rumeU70iUaJmE65HZW8Rb3qZEeqnDv0WLaanGNqaT
0YmK8Tdk0l7k+jtvJ74vVorpl4s3yCjuZYmkdvMkKiWLQ8RyN1zjtBxvUqoqvJe4sFk8XowCt5B7
x3mYVbjX+pEvXV74ro/NFeZNrJy2DwP7HhBwftl8+yt4pSS67gSwvE9r1sjgyRtLye3vJK136eOH
v2kMoP89Z45qxZd5X2ZiP7frkSsLPojJ09XybSRPA1cltZhY8uRUnCC8qbNZ+0TtLnPd2CQGdcVh
mdaIg4Y84x1AQfEhbraHxoUCcHrw5yk3DOGehStbTSOXNzhji7K/MgwJbx55i0SxrugoHKCyVC0Y
44+kuMKSObrxTjQy6B2MBAZYrdUQRpoBJMC/ktG6FVaoFO/lD0Afl5gEOPXwIpNFrZAt9zPkDcRw
S/rRsyI0zlvoX8OrwdHNc/LDtgVf/714YH7r6+uySmzStgrCAYqvqttXFJLMVEbiqC8+bfeekrk3
+zPpUouAonWLr74ppGR+htwULluqVFl6VV5NQ2IcYDmGpRp+yfQFO7HM6RWT7JI5G2TGtyDwEFlw
wFrEcQC3NosQx3XMUkYquLEdjtnsxuR4zij13vrltb1B12rM28GHs5rvYGUmXNpAd7vEh9YsTHPQ
kJpuWkDatsSeohpkC79IXwaSrfFeYD4o6yh2e2qbF4h40RMMkPq2H918bOupZM41W8z8/Pegr2kL
JXI7JZaQ89uXdQuvlTzR3q3mtDqq1FgiCNlmRjhWDX9tSqwEsN7iNwra/5zOMCmxqs2qyEY5Y/iu
bfUENzjbrYRVSi0Oy6My0mzQ9GPjS9DQd4IlA3HHpIncaGUv+BZV7rbP9rU+SXXbSRydBv+d+rMe
LG1q0CCqI3re7sIMwPe7GLhPYwk6JUnyXzLLEOF82GXz0XB0DehRysUpT20TysYTlSvluj0j0/KH
prwOR6pm2jI0qFCPiK1HwXdJinUJOEDsAIzgihfLn2KRszpqpnLmzpliug6xkZvMcCXwJjBxKuQV
sU3tLiMFv+fNLI3Q3ulZbcyhkNZjIzFbp5YGf2/DWAYay44tZ85dD96UXkD/7dj7dcEy+nlsuTMk
pJNFSFtLkcOtMjWtmUeIBsbCojI+bmqO12qi1ydwKMvPtRWU14SOoFYPtd+70wc5oZhrygAFEloN
w/CIeu2EeNUAz3MW0zApFqnqhWZhTJt0UdlYXECbgvV4qjbNInXoX11WzXSh1VgdwInGxjhv73hS
IxmwOSuWwGl5ryzST/FcG5EKKNUEswJolGxQ4WEVZVmUTV5W1/VIXFIlcK6B6GtTws+MDGrXHE+r
O5ZA9MrbMIoLwjGwX7BB9k2lkb3FYMt1ePvJn1rfuJuMGE9dklnaXaGJR/Qf5z0lAfx1hovITKmr
udY6QPbjNHvo+XV+fjGAkv/Zy+fWaMXPmZFlGFaWqF+Y7kcjvSKNzbUJzJ4mpf/cbexFWG5/mRS9
8b2D1med8V8T9cT0Mg80kDwNiiIvKwoCgTHrj4yfoIwnSt7NVZ665EHCpMptTdPu/h3IRcTBhj1e
EGBcvoMvslbkfqVt2uRQE5MZuMBGfsuPIu5ks/otuwEnoLqSSpQGHl8eLdCXNHTT1Bbi2clrEpWl
Ao4ikRrsoE41qJ7hW0/KQTVLYCNNjt9EX5YAHcdl98AamqeHn5DVv3tl3RopaoxXyAeHg15dMPGl
c99ppJVf3Pj8r0Dx42PanGkQ1BwzBTcS0cl9YtC4cYgpS97UbayeVAPHjCwooPNC8AnRM2qD+Cx5
UedA3wTxR21ic1ElqET6AEx492Rk8xkOCNTMjsgo7e95MAyoJhip8LzO7i53Cv7UI74QDE6b+l3i
pwrBlEH/7C3WtR0ESDk6LI5hb/fWgxTjnJX/NHZeIft3J/tFGzuUMSHE3Wg+skal4VvBMRGZajbR
6eqgztDseCVj+QgRUwJxjjRB7pefWOK8B52hphk8CBBIfBsjARNDDMwc+a17Lzofnhh+ayVAfPGh
MdAkgjg64XWZO0FvxevfbjQcimIYatORd85C1sdW3EOP8QcgT7GfqlDMnF0s+7tEj851lBbDzRiJ
ORUuQyc4/VxQT+wf9XfYHv37D8TuQ9XZeNmDXKj/GqUfvdS0/Y43hDSErk7UEUm2fR/dFdDxAoK4
m5oJlu2SchsjOopyIiubw//STyNlh7OYr6bKvPf4QxqxvRol/B8RoSnD/7mVGtiDz5z5ap6CUTdm
amm7grGcrzL+DsjHI9wemUrkqJXxODU8wAFNJtl70mxwJw+xA2XxNrn9OzpxTsm45zdvCci6Zcew
w5VPi4TMiiTqNzMNOPly4z0UkbIoFr1YiAn/nKyOEye4dKJK811Ve2zYsIVywFVVVukri2n3gXSC
AUoA/IWAuf1GkL/myO6u23nYV00W8EvveHkCYb1dy/Gdc1xlcE1l8h5ehoGJiMBFh/7D36JErJwr
yGMVSoP/kdaZERCAdI1mJUNYoj0trZyOESAotwdtzFGt3PyXhtwP1v0JnLNZpXsSs67Nhl/KK+uT
LuwjgBnf2L07RmH+G54NfigCQ0LQofnfZSaaAhrN3PIPDh4Zmf326Q0JXppbwxqjYIHvF6gpuFrx
jGpe3ntJkB6tOaSYTfisRGMzEdQknGySO3SZWquIV3cZ9/S+xPAsPeqs92oFcUwPffFaCxOKVCrk
T2eOovW8hFLqOYIzQzKnf7x9U1z8HuF88r2lS1+QNfkWA8swfx/V971SQa1z3wi3e+391EUyHBiL
UP1LJQlXX/Spdwi26qnRmnRIHtZNr7wU+KU43iUPDiU1ftkqzPTzNPX9LZYlyM3ACeVwotchDUd7
uF3VvB44s4D/kmpsS4OSRug/IIwMtSCit3/blC0PaD0PU0HXU4nIAQELAIaAgEUTOYvi7oXA3elz
MkZKvpMqKWXAWzsf0EwIGBxRvswtEQOcKSS0ZizNWISwwVheGZKZ4J+eOerM7sIj8Zgn/oVVoOTR
IyxQwet3NuKLulDoNuSAAG3p+Y5jdwYyXCM9fdrjPvYz51uMGEqbltfMGbIQSmDEPja8mBQfFe7T
GlInN7zI88AGyz4d2byudFPouWfq19/U1EYwZ1gKNwZk9+cCBr6+L6q9RTkbhQemFy0XeC8ITJbr
K7xxg1ZAy8PFL0ZCv/xjQl78oCmUzmOV8tKB7um2YIHWUdkZHSzA0qgmPJmYnrgyF2TMLzE9V7eT
lQ95l4UmdQETREAWHzxbPzo880DGWijUVvurCFziltIbrVsC6qucX8+8lDGPB9yWyChwDCLEAX4R
jcDlbfMvFm3/0Fk+lPiqRzYVSe38z08OxjWdJNOn45lESE+sT4Qta9P12KbqA9bNud8VMKdPwxtR
Pv7CB0KaBdF2QFQKa+9u9clwETmJvrScgROt/gFlMZh88IOBHyiCKhYyvAZ8LzR5HL9EbPcTgPbp
mF8J9ov8EoSDE1PVi0HDUgHfTwUegct4HSt+PYHsSwErlDANN+P89+H6kv5lIqTVn7tlWmTDUaSP
V+u2v9WPDAn9ZUVzXuFgk9FJ1dVD9JfhjFxbJr2uAgsEf2GECQuR1oibyGdUHpgyI6uyRXTvfRBG
seaT4FjnFJ54s3VwIJ1V33FsqshZ8AUUJs4fVdkQsx4nZdzbLhVaCwE12BSEV+E3U/dkr2YKNNLv
jTp5BD3dD9xF7hdi+9PHCbM0tvhvVjlEMVOpI5mpBrv2w4V2TlAxzGo+5R3DxMq1mO63cs0WLugd
6fffFSb9p/WX9092bND0tnnoAV7rm0p66eXR250PbaCuc1tGNEdC3OnWNlGiZ14k15s41UCklqgK
F/r1UhOzhrfFpNFJ3zRovBtHGUyfBlmc0ZzyITsShXssocdiepIjtbzqtLDsZhqjYf7vTnmO/t14
+lEmC+2gh4ppHbsME1OENOnLShOTIxMdyFsQGzGPqirIcrI7MKkNJCics/0mZMSQJ+OHOXO/6SEv
X1pXsIiLGxFyCw6Mb0R42U6CrDYuYYnfMy9ZRYvHuM39m/yCftg//wyyqk6aMjYaxpx8Qe9nv8L/
lfOagfgtSY5VkaYZcZVGDPUDtQPdDTDqVYBiKqnBEP/X34I7gl/RcIiZg4N5QixbbjFNru9LCZ/d
Rr2NFkPz5WSy8s5wEgZBjQm4OgRRdvN9HEj3BMa4CMmygiAB3RpZAL6oBSY9bUYrBlUuOp69Gymk
4kSzHiaUhRAW3dcnnF13x80D8EBKoO5WVAYONfKPm/CV7lU8wH2ijiCVF55TS6qTs+4xb5dGLa9z
sJGFrgo+zhvO/V9O1IW+Rho2U8o90oEFC4oDRPFrgDt6ALDHtLEq8jr1Qx1htlw1Uu4IKdnlcbv/
BT7momlg5vVNO0rKjBal9DwaYj1WPyytMz2Kfve475eHMsA4WJFI4dx8u47KRjbIUANI6D/ephYb
apDRakiBRslcrc2YxP7Rb3Ft8dWCLw6+aP6aC3ehmYjNfd89LnHpWolhT4k9AqqjcstwoGb5T3Ts
TBnykCmXUi16Z0vISbOoCJwqAkUWvWLKLWqFpwm0erjw5g02SnypCeXaAAqTlPfa8Cxmw0cSzvgF
t31+uPo/tsA4ZfRZvvwEShoDpecOgqGSVYpqfZ8D05y7hus7VDYQk+42ZI79KhgOJH789KzNnD9w
SZsw4h/uZA0TkCwMqR1uJYbbI3IBNz/Cw97GGQvOTHNWkXsGghLjHYDW/1YfHZui3KZ1v6ZukZ1w
yd9GrJ59bO6XpKUHjwC4B3TKIBpl9oIa8H1XbyCk85obTAcCRzoh2UdFVrl1RRTmURaGWjA0qf+h
DxdnpdvgCD7+EzYwKpHO4jdC2loCxbSanItIPmX4scqy6LcCUZwcUQFMUL2Q3lV1Y6O+gTxR/ZN0
0n/qDTW9SmS9iLqNdYYaoyvAmTrKpAvBorPVgYkxgQ5p2k/QdmoraPlyzp6jDXmGJ6jEs8VyUsXe
5mntDxuY02Yfg2wVwf/aIh97rXGNZsZMRDNjSi/qqXdTfNs5uaDJIwijYh1Y6H6CrADg+djVBJmF
TH8DzuGEhkVlAgjwzyo6REhwhNpJxXnHc4ZiW+hqV8noQuHEG+mxADzstb0fX5slxAxukHr4nJe8
s0FJKI3CNMUMfaYRdYUN9uia7RgisiGpWXXGZrHCFb92GZyhVYR9nQAuZG5sX4gCtLtfVezMAWqW
KvYI0kIikU7jpD6sMMHLEq0pzArMjnEWg5pHp8sQhjo2VFFIAr6AEmt/dJmdzSo4kXpnprDQSVt4
Rlh+R5Mi8fx174IjkCwfkgMWjk5DjYKO/yt//wkHLdHYlIcwB8e3XcKwud6oamqnLqD/f3pcQTjG
2uE6Qcl86I4ViXaaseMlV7KQRZUc12Xprdxr7z32/TTpoqlee0nzYSmIP+0w1twDMOpWwrxcJ/85
YThkEkq0TPjzHGXSj+cSWCmg+raSgKITbGu+tvNuM/VIFmZLRZ+lwhTdTyH50GPOw1r//mKaw+0v
U0aNpA1Wx3r8WXoda5G+l11Ys2w2A6lI1sRkK4Iz8Gzp1ZM4ap9i2XDpJkuUDtaCETfFPbzyrl/y
H0M1jok77qsDaUb7NDDHfC4xRqPBbnrzuQVuyWYQfxCKsnNusuf3hcdGbSi19WqnOGts/qdBOUoI
83dsbYsO/CzW5RhIXP82bGaIlhBJAS83VyfSGBjYkOi7OVefjpD60QpN4f96MgTfAquFVfPBQp9L
vqgH1E0Y8DiCD4uiRJqu7bLe5wLzBBK69oZQdBQh+l0eEDwzB9NH4yHNWek5mpcmedpUJnCoujpB
tlcwbAOL8p3NNIVIQf/5b2cEe4CnL7cxm+FpeYMj8r7enxFiMNdmeVLbrx/FE+6HxvAx0P9sfeWb
PXIJeWMtjO1Nqpza6RqoHVOcVw+MLfWfo8Nc+pkPvg1/GdJB7nZnkPH9FOoVMIdhkeZLfeoLLcCW
Z7uwmmyCkvJM/4WS1Tg4+dJtgERDVi0bm/hjYzwQqA4o6r2V3HrFIEJYRY/g9X5O4syOxSZ3hMWE
tWfGSyQZ/5agVxeGAOOC5M2ayNbDhFZt5RK+c8rR7Ql514rL5yvaTER02pdZ6JrkXSTiP47xYOxK
tMvyLJ5I6Mv/bH8NLEgWbzRfpc1Efsy5pfbc26GaWpxfC7JQht5FBsbr74jmrxn6Zwf6W/PayrOY
0U8UxDdhhWiXoo2zqze7S1qoNcwLYdDzdUDe/Pwu5WHyIgrMl3cAiNt+SzFjI8lWWauoJO2BS6al
NS2PrtE8U+y3fr3/NocSgf8OPMyDepejhhCPMvbK7ODBw5s287/hH98Cbs1VdJK4w/VXRo6wi3Sv
hn9TaHCzqwJYuMHiDAtGhmhfofzHFt3y7pwItDNWgtD2O74H9OIMmzG1e6gasUpIA6lyNYthV+jh
IdpibFAuL16vQyexJf0UoiKFvotRuzQz6wnHwmzI4piviXzliOfmms/TyBwnqnrieC1bl4Qh0O9y
ZrVn56MqvqZIbpEY6xZpHpAF8yr/vmFNMq5pWD2ElYxU+/ei2h9EoE3Ad/fBcv4OXT9E25UqSLph
EmwuUhH+qteJOc6WUc5wbCk5CEF2Lb6uekRpEObPcwPXUUYCSJD8xdqHg1ZmWdgsgeubVbQcXqxW
69vOyiCfIndl2IJNjJ5WXY/dr+oiJnjhmlQm3GoqnwchpicMGqUWqtEshV/oGvhIUlofd2tt1gol
L1lFjjt60Y53up8l2DcKsN1c5zs4T6KdI9x1t8GzsJaJjPNy4fz+71B5fjUjDyBQdBUnLZoHmT91
wN0+aExpZvgOoFDy/7WSv/36wscNvnN95/+p6ppCvVT6+NVxa7JW8dPQyT8vMrAAQ10kbGvz1gt6
U3CjlUuVt3sNe0ZVji4aRnpFlE2mP41ei9XJ7v0Ok19OtJ2UmViF6sNLt9ppU9m7Muw6jJg9eTBm
yftsc8/Qa4ZnZNQUHCcI9k5zG3ymYdtnLVl4X2VSAiigiHkNfso5Rfef9Da6iP6A5Y9PVxtKrUT+
lbIMCvf2ZJklQU9QpCxgViQVD9pXkLvPGb7g0PfX3DLeje2kKX0GsbgpNTbtTLpdFnR1rTh/5W6z
yo9ldCfvB3tk/d1wLOjdd37Uaa+yYRM+AYG3eBUJ8sEya1J2NLpCMU1hpP+WeF0qnqzFITrI4E1Q
nzwgu3XghuNTUHLa7odQOxW213EfDqGQZflyHkM7Std8kdzBqB4Nj1wAlOEDefxUdXkorpqvUzPw
SpeHY5KmP/dCnjt1Y/Mp2ODP/gvkdrkotNpY5JTPAmo78Hx9YJfm9PL0bwacM5lGLaOjmDic3pRN
eTrJm9fCs6OmAvzStzghLtQL18aNLyEw0/dsbpgOimEsbLC04FoBv221o84BNcHO/lJoQFuCOWh5
cVUdh19NnXEHRVpSUUrcVwio/KwJwEAkc9S99JnzOxCesNljqVtRDK5RQqIwvU8EOBtHdK61Lqkj
T6+T5MGGmXs+gvAYBuh/Zw4m2hH0zp8c55EKZRzwAztTpUcWOjjPpjAwO71aZPIxUVg9rEn1INg0
zTbAAqzR+suq5lLMwyYDOcPU6tD5pbBsYRJSwW2PuEZUQ4ydKzif5sFvsJO7KhmrFIEriYVIekEs
p73qrFTLg6zXzqjLvFHLqZ8RFvqCfom+51Cx/Vr/NknH6BuX2SmJ6pBX64Tip48GV1kdOIDWup6s
0z1/zc38V7TYVXtqqglpXPCuaz1DNxxAGxR8q6v4Osd+nIzXI01kt2WxAWDwZ1nSQM50ioTomjui
fhf5UrYkmR6HaU5GmpCIp/HIaRTILdaoynsABelydPUCaWukuI+iNL+xcNZnWAuMana68/vG8lSs
ia1oBiMIDcNCEwcKhGRcqcQFdj5hYBCS7KJFqf68p2ZH+R2fMk/4N5H9x6XttdBazdN0PN3VWMfZ
0/KQs6N1VxOQYwHglX9FKW/F7TsOJEhLp9oK/XYBpNc292rdMg0bz1X1duJ+wa7hYn46f5OsvtOy
X7BppWqNxkRTdr0nLjkwr02l1LcZGNzdX2m+kHuolImPEaNK9v6cCOEKszLb0uAeKTykORKfyfcv
yEIfFXj8BKro4R7i6h5TOzIgGkVRvKAt10SjjQf3W8lyMfKBq5m+t5UeKUocMETFb7kWfd6uPjat
Yeg20Y/h03k7/IsMRjywj4GdaJ0MBVZpf6c2t27gqHZ1PSyu4sqD2lr++7dVd6SO9LOxViDz9b7F
wL/KeScaueLzm6w1w0eKye5SieX+AjmPAuDMxgpnvjx0kGdIfprYPaBwZWPMkQrAjEwJa1F5bxAE
rKpvg8telB0ZopwodfIW35PTjawZ8iKgUc/H/gPbZpwxBb6917TrzU196aj3qcRYSjjD3chkPaCe
4L5FRLnlwazLWZzQsIo831lggo01ZGLE2+j2GXKdnQ5F4ZiteJw8zYBNx4dfbcA+hfCwYn+pMCZV
6k0Nz/TTVtXIeTeDBGWCefuRGaRv9R/lL9gvaG6i3vCDPbB4YpmUm8OGYgOYURJoHaaHyR+7/8Ep
ziUObLeru/ZPIinT/9kOoPEewtrHD/KatbMWPc2UlfAF4+ryPZOhcpzo4yVXyk9e2kSnHycD8kR4
L8G056cF8HqLn99PV5NZ/ZWVU+dulj3d3FbM7Ryk2U9W5xfyeUCBBbnt6h7R54SCxKhPau6raZi7
KBQk2A+6PwvUzlsWF43U95bsasS0ZyCnaGxNx7eqpMJFDtc/qoe0Rn0FuNr6j9B/Jh8LHTlnKdZd
f6uRYhe3W41n+hxXXGt1jxMpxzYD19CEJjBjV22OsFO/qVWz8ugAAMopRiNi454jERpPyIKbpvpl
uMmEHdSA641XXHWXVgsVfuh+RnBPS4eSsuPif5oJUGZejNWYS19FgNJT4BistY/GXOL7RBBliwH8
sgx3quu0hY3MtIKvidctz8qDR4+papY012XS9xy2Nds04DZWEJx89FmFgX3cUjiegHck67Q6yr/R
Wb0RKvu7LivPNTwmrNYweCdkCPw53oqJGtJldjj+6GQXYr6ro1axie0uPRL3hrx42LavoaN8pqpM
p4gZbFJeYmm7IU6Js1DNT2Q+Sg9Zn+xZ+AVD68oiFuekl7n+rcQFnt/J6eZKGIVcyjtZ6X5xO1xK
yfBGQPk1a/fne74J8QOGe3PzLI8uezzSJQkbY8+sAhlpvlwt0y/eMRrGealOXd3Gd6dr4KsM05tP
76wczKbRlJkKTO/9en2bebZR7WWdpeRn8pWKRmfYvRoEsoo1j9PbxUjlfDVoAQ8nFuGjfq1eMee3
atzvrFdtIwMijTeC1IKDbZ/EItqvHy7MBq9JNjmZ8tJ/Ob0KgMCeIDiw9gsg/bCVXV7fpfujPNMh
WRxIHOXEdUYmrAbUYcE/clZKKJWLcqEZNCZqfXOp+RPEtuTSjkhqPIRNLaeZZLwtBWeFH1S+IU7U
3NRPktEw45G5ZPzpCuYCkgTpP14nuEl/B5HOkfhsyRpvwmxm5BgZ200IcvfqhF1ZQ6YwSBPDPZDz
RQWYums+U8P3gmFJQ/YZwj20aj66WcSaLcgEZC8et0dZW5VtfTb2MVaPsCZZrWH3+fCkTlhMr+qT
wtpAFHuD3By4K6g6fkp9h0m0XUkJvx0N3fjy1VLdUEKAeVh4nDIxNeD339SFlqVgTAdCFz3+Q4am
cFRSZ9UseTCiPF+gr/IsKgHHKXvwoIu98zWUPmkmi/EOKGo/jA7NjdFrUE4iyXIcuUSiTjh8jYB1
zTG/y6RvwYT9fiyVkAdQltApW64KTGiQfnNuLB5mf6F48cLuqsIaEbP5lrbBl1RfGW10nESCR49U
vgEl7cpFnOzCsTMLqisuYqAifeBs5rEpWoijiwORJe3gIIS/JonLQPRwbiVGRaqfmP2KElAW1qc2
5vOnvNKoIr0KSNzaOhU76kcayyDfL3CRkEJ5ADxL3KMeEKkifeXKd/7KZXlujOROeKKfmYbumAkb
X77q5buultdkznRc3T6b5mm6n6JiVBOdAtmqoZtQnQFJJs7SD5EgQkBnJ6hK3dew0pu7NIrulGsN
uxoLqJ0Nk+nXRPNPI0hx5M5wdLZWSllUjvMasdCOZsuroRdfFdVZJE4iAhkOF7eUBb3xngbPtjTq
PSUpRH+S/0KVvMd1nWIWErG0dvr92xwxn8seYPGEk+C1SplG5rJqkqjgHQBj8+UUeLYd+ahFMSF1
c38hi2WCc3fLP4B/T69LyHlVmmi6N4EPwd03yTSVLe4+h5maRAU+7B+BTrXio2UARPioiyzCNOyF
NFNUjZy2wumjUkVtkocIDF98KAqy+qLBtqeRyiTmkoXQkB2tF2VxXf6N9Tzv7ePnOMh/MQuTARZl
UfBTW6NJqRWJ9wk+k5QhyznrWweeII1GbQDavw1jGKKC8SdWXyG6iursgmNSvzYVKGixbhIh3MGY
3Y4IgwxDE7BWES7e3fHvgb09yRhUTXEtcjVHmDxsq7FublxGqFQBInH352DKM/fEqcf+cyjFw8lx
Rn2C7niameEeXvJTeQp0Ju3Hzn0QHEP78aVXlysU8R4Ma0AOWKRRDaOwnBVJ3G+R5GYvJnw3zKvQ
hzlZGhWjQ65VQL420QZd8vcBb5hUjBEiwC5qjsXoo3ZSrvIAAZyyY3+o+C3zVRh/BnfwSWHzTNNj
wD/YaheB2AHR5MuGMHMwZZeRc63okIIhs2Pu3F73UQb9CjEWewQ+fjSAbtAPr0WPHNsWURgIe4H+
SZlN9bjN4axeusQawRv273MWdabEouBKWafrVzz21QRKHnDkzV3IRwRCDYIfHr92onxGJB35gnv+
TSUfZJcRGFTU5zMWbFVSnE5xZ6TwHsQ3poOKf/s0VBTFklvrd2XBp6T5e3aYWxvtHPdzqyQ2yXum
wsqn15cnAeRXG9OKn6K0P6bCgdZ4uLPtQnKny+Pd81DDV8tQ5jad2R3m+AlnmjLDEDRMb7R7G3EI
E+SfmNkWSFDdqOmfjAZ/NHYxghyU3cG+hWPak41nm7tzmrpB8V9x3STcAxBRJMNIfzSe/Z8O+4L+
M3v0Wh8nSV51bsQ4OpYGdUqAcEor6f4O9b5UNS9oqKyZADxV1eFYB8OL1lJsEaoienAOkZs67Yb/
14YDJ39itItIPZIgUwzTE7nYs+aK9PrbcTReVK9TCKs+8XyzmlTP+VIJ/lQkBZ0iQjqN4Cstn2eI
TK/CegL2VA8jzgPa3ikK1BmHtOjwfrkTwkSjiVUZhf6f/yh4BbDVLdrRixqXceCPQLjVFuD16DiA
UxnGbH/+rkEU3feGB32iL3Jan9u8niAlF7eHYCOPUc9g5DmdUDS5V3DSQc7DSy8sZTwhmbJ536P/
6MbVfEhZmPqA2mnTudKjG8CF9bLhgu3czX8TXrIQ6CZU8ghyuAw+ljzgPv5sot78yvGlAkcVmXsp
Z2UNuwXxRZPzavBnwjX48tdTPUesT70RsA8Xsx1iXjw+io4E6l0F+mpY00POt/IyT2Zx1omnrRrB
7BUX7d1ArGpFkQJlGpBiBP2AClPJixGKe8VWYyEK9CvoXd5EPWA5c+FZOVySLsjv4P2femzcuefo
300HPugIFEIA4/Kn66CCfPC/kkPNveeYoUfKnQVSNiDZEfmTFCC82A5/7PGCxAqgmN1V44c+7wjc
8xAtd3zQxvYcky02Ty95ybMvN/MniVbJ6PV135Fr76fE//IyZmPRuoSzUDlrHovnevz+7Mop/LuF
3oQjHJmH8MPSjkzUoqJ9EM+NNZarC96VioEu7677R4D3J82M3DtAf4lR0Y52jbR1J4aQ8fVm83e3
H0fVIT6Y9ASr1gowtnZYFsVBKeLYBG8jy6RM5WkuZIJ0fRDuq50fwWd9rSGs4l3B9olQP2p2Tuum
NUM5O5YFUc4zuVO/7w9cSYgR4wQ6Oz30HiaL1VsHdX7KBa2tn/7m8vMsYLpyykLkj7qvRxUysOpg
lJbC98hY27esJ23AN/afJXx7DzSwZSyl1vQ1c8lpXd16tejC5UlFY9HB7476jIVLsDDrvfwkHN7/
aoJfHEyaaMmUCHOfkImoAJD1v4uXTgW5F3++pQnzHqnl+pTWV6XJNYHUZz8ffI0LQWh5aAqG67lG
blZePugyZL18xVkVoz2Uwei9JzxX9hSDxrtz+hPJl8EtxKlxRWUgui2RWtttakIw5jTFNeIv0XZ7
OdmkWPTUhhu3oPHtJMB0GB4cHvcj94Hd8wQXGDk2mTqNsfgicPDD9fTh+rFfUHdRTMttYfPQGUed
yC1GW0SiDCunhLJf6/2xnwG+Wyee2k+tSXR1KC5Y54ioOe6z+Gh46gAwWh8AzbaPBF8vLEM0CwOI
iJbSuLnwhuN0WRvJ3SgN+SsKaI2+rpF92CMNI7Uyu72hEjwB1VgiqdALdmS8f3GSyvUMd0HXg1Hx
j0lXdGwzJORB3/elxa2qFzTenPFGzRqS4AJZGS+Cuq8nWassRI13rMTldnOJtACQicro5ufxni8O
bnon7qsFo4WW4sCDqJPBJzg/Ja4dbBgfuIIqxr2Xi585/TNuvsV642FBqxsQPskUbL7TZo3lcJN1
AFliUXKW0Tjzg76nL8WXiQXL77Ol8GxWv/eudTk+FZIH0FSZolH7dAwpuFnTApjc04ztaWWJZGnM
AFJwj7vAR8u4TWqI0vi4YnKXEoe2wjDX6BZ6IttjZr4/KtpgNhYlzEXJxXkYM8Kq2syRcZTowGxc
zCy4xpcpsPe0NDXs9m37IeLqVeI3EV3ChLt4uWZ6YDkOdQpGX2jZMRlpZS/jx9hIAmYQn6g3J+EE
HYF0ixeZlmf/5adhO5TidP0G/fAxPe770w+9MMvGZqOChN1YxZX0U59Uck6cwxykqYQ84dKQu+DD
k5ywNF0v9wGJVyatg+jiUJiMOwwJNiyjdRqGQFHJRO1ka1h83YviNoEW4oXNQqx1E3NOdth1fYwY
vP9/b684ynDl7A8KlzmBQ3RFvWmEwEVcKg9XMzXGskkMoWetqL4woD9bOYNI82IyAVcv5lNt+6Kq
+UYzW9y4kFkCY/0Ar8DXFk8OqoK3Y9cgU8ZuhNUYuvqmkKYC5+kDZi/DL1/5k0DUja7rMS0U5fxc
er8i4FmfSHOFAC47jJUqL0ehqwhGAKGe93oU7UGrC6SNzXcAFFFm2qKQHxuzEhoQ9tAGygi1ggUZ
p7tw/8Gn6cU/GC1ysKqiRjLZiLii0gjWxntHul4oPaQbvDqugrp3njU3l/era9WL6e7znlT2e71Q
LmfKkpqNmPDcKe+7rqTbdKtqWNw0FYC9Xycor+u/N9EpQyRHTJgKhmff0cnhWGHCpnLpU0XZtLa2
102Uwx1rZNa3sSVAR/0Qovg0oDAT/0HlZ1eDZZ1syZVVLkJWFvPAlsGMghytjJGnGMhMrM8HBJOu
sCmRJ+x9RhTc/cr0Wvy61ExPdScahSoJvkNoZQiGm4izYvNTmuktBu1OzRlLpkCV6ej64h2ohAOB
wNH1DIRT0pykuqbF2TCGB7kvkVCTaG1odsTr/R4/7Us3eFuQr3z7GcNNq9HeCWnBpljqeMyfo2PE
UKI+gOukOzF/EMeh0ZtzObr1LBDq6RQCypcW5L7EGfNY6Dyy3hkAKvAp0mC4t77dimGdHzsvy0TX
jmioNa6HQPE1ZlkUO53oxlFxoSSSefLbjVQ73DdaG1y7aPQN80Fxdx2M9WFYPezDUISumR1wq5QQ
/RpsrvxZLO1n++7yRp82ny20Arh6rzXq4ji43pBMkgSnMRyyTl7GWo/zWjEzDSIRs22mJEY+zpMT
KE2xZ3cz0zqdSeGeJdJYLncsMbIs+XZ7R/MEHcZXTWAFFkACt85uohj/f8PB+rLxOqi/lm4adb+K
azdyOxUO93DxFAlGNz2mMRZarlVaOdBKZPMgCsBDvbBi0tuMeO851+nk/zJtIC74YkdUdh2WpYLT
zy30JDWzzZxqJ4KNOLE6sjQvZeVIZDa5snB4DoDuXx65/qPB7kd53nrRUA1JSO49GEGx+ziK2wfS
E1ucvYheJK10V/SETqtB6uiXWQtJcbRVuHN3p3JyojL2Uk1f/ifLC825a9eUrswSU2zAVnY4hSSi
p2cW4+20tD+L9fJv4SSvXDRwhOQKQ5Q8O3rGUeAkGrRT/U8n4qV8P092HjEDVVaCBQO40NDNXh4y
+lH7Pa5ZrBZ06GV9ttqn8soCMeAGCxJYSwEazMfehuodar+3GvzcK3Hg8y7jQWSBkSiEE0xYKvTy
ZOeGIAcSK0W9odjgV0T1j+eX2/JBp0UDCR6/6u4dJubB8ykcI/MOT1vYzPEI0xYN6mEc/5mSyq1v
htz/5FDcTF4R8I1DQZ/nH0SSX3IzmWMtdl19diWljqXv4ibtaGD9RM/7DThJWk747Hfn7pCaKmnH
CRcnDhJ2AzJIdGLBBnuWl0/moykkrXbuVuY7jUCc8V4haEGR6fu2y+B+0dK78LFTjkEPIgtvlQao
ZANbGTC+N+iklHeqoKGpwDwSHxwD3aiJ12s9EHnxTbqySRXh43y8LbhSeycF3y6QegqFr1OEQJn2
7qcWNM+qC6AUxs0vOK9drmWbDpQe8fNYvpslsxQqfOr7SctYyboCPoDcIk1KHmmRaKrlppS0v7NA
f6wzbb5Dq9g/isqlyCD9e1fikwaITwlLL63cdVhMwDalAGF191Xl1DnzP0UdVpeURug4GzPWhPcn
xaeLM7isKQvdP/ohpI0OwNu9ZrwIvEyXctdXf/j6cRFQ1lQa0BQLmwtDY7vRfIg9vzG8y5/QB1aF
mSMRJz/YyRq9h8akjEdHe5RWS7zcjgNXUO8QTNFzA1EB1hWIevrAqBL5kbRaKsdpkCU9JH5bHTZj
Zi4UyJpLW3Z7+Z36vJtcF+F7isk4aHWYwVJVn9ywwkGoz1rVSE/WQ6HSHEEtpZsvz/LAMpmxNLut
Qpc1r2aUaFI5Y3x7XeYKcumbpN0BTHvm9048s1zQR/BCNR1j717K4i8Ok5/md/H2PBdqpbXTeiQn
wJOxxp+y2gClIqXv90O3/DN553rYj29s8XTO/qH1o3bsMqhgbZCxexNteGTA4mTVbmIU2Wt6D6ja
EoIFr2Pa8xZTZCruYrTX3AZruAiY83q1em95SO8cGHEUsyFmnLVOA+Nl8rD0+JHCbZjLWw/gPDBM
LkSaHccw8rRyX65gwiBVWcjglKeqJLb4egvETn5hgR7TAvuaqhATWQ+UAA2TtheOsNh6nvbZJ8ka
M4abrUbh2/FwkWpkPWvSt85sQpY/NdJUBuq9VCJR0c0P08Ht7POxaHl1cx2QcFflArOwxQE22+VP
GYpeypRt+Q539gLdWXFbPCvI32B0UMaS7+IyTRB59ovNb+hwDhp8Bpys4TmaHgDXXI5S7MWSicT3
CpGhXDSvyXCONzRmtP5LRgBzz09coMOjD93xd6yD9xZFxI7z5Q6SkLkZKcy8bORPKc4qHy+DDOlx
4pmT/fp1qUijxd2GrdIPmkwKD2d/Zm6o7yvMyz4u/LqQCkitR96wUoLdZr8GzHqdiYivVULElIFR
5K5HblQQHowD7zUztftzA0jqvrdOzZS3ymwuVa82fEfmkjg0BBQS7RLm7l/M5mq7foUTkeS2svYg
t+OD8FOlVndtUHcOkofXK5uYjqcy+TjXrxH17wAgzYTal0WPmPnnRor0Mtt4s/81miJhDcIW6Kn2
44FdEYB38KoZw0M9R10qbDVzLstJSWwR2XGWPERnzaF0kWEIYbRauAyGLaN5NpuJ97+ePF6kC56g
MfdwUchxpmqFQfbR8wcJOUsQ0Gv26D6OSoA59rqFtCDOWKNhnXHIHMZZNH8AXinOigV6h1zlz9KW
SJrpFjMd7+CtnkB4HIksdTiu6+x3dZzasXGoIuyUGybXWZzTxgbx6oxYeghJXo1fA8s2OkO4Vw3X
AtkcnPhtSpmLJU+ZdI0+URfbgFgSE6+flMCZrLoKNT2fEPl38LO6tRu+fghjXSgYQ1xvCbLVVmR0
ZmlEG422lqCflxuXCWrRnrUCZqHu4Vos2q+ECQJUfWnPf1cMNb2Vabz7GpHPZbS/qb3dJxslm2By
OWUD2QfWPU2Bll7Qc9xL7O2y8NM3zMafQ7uftqNJPiNrZ0wYYICNUsHTGYMr7bbmlHkrKf9DYrpw
qpXGg/6yLZUaRrPFABknKUXXNgFZIJDoN4e7jIcEjF363qXcFt1fFVl3f7NqWJGjSbnY3G/XfCd+
oJwwHi5Tp3Ch6umwW/N7VZLmuTa+3kAWtpS62OygQ2DijL4bY5nU/grQaoeU38yvNllBf+se+8Z7
E6OG0okl/uBq9qwR0u+PRqq069vZaCgsft32Q7yJBnw/qN5y8xmxOO2Hebr1uWgBCtg9l7H4ZaXI
MWIEv1o1hQfbHqrCI8UWZcilCeJQL/iXXBJNEOAi4rf4xO30EYCvoajs9vRlzJ4Q4VHUexaojB2T
Jlra896SAY4WSab8xwZGSCPd9ko6YldP/zziBjiPrr4sCytx2+8Lh2TNgknGu+MAXwKGM+9wV6hd
pC3yTaBBiPCbidhtLIQrWEgRR1Nu2R3MRKkoyoOdfisJck8aHzQmji9AXc7l+QwC4RFJbP0uxDHp
XJy5k+fDJxrnKuIvZk/+RBMpTq/kNwN/unpOel9H3eHpB2rJaZOlqB7BMCkiDSGKx9jVrrXb1/u/
En0rw7owFRczDbTpUDKVVWNmMtQIfccSky0jFXZdCt8hhyP2k4wxhvAJ5fMNX4UwuDkubslecuZq
tvAnVyDR8iJ948Llhaq0NNooPcVIRgjIMUYxq5MZeSMqZycGV3XqLHxL6tOzgB8/9I/UgYHDQKr/
WJuPoZWCTvc5Bn+gkC8BVSFxum3vBlrkxXdD+eAaOmRyijK1llcGqjZo81YUrbRuS7fl73RoMXYz
9zvLhywAjOfsnLneRtcrpzEugU+o60KPtva87aIQFdnoCJlvdw7ZjLKOu7356WBNTOzEnxAmzw6G
GfgCExaB0I/T49PR1/5BLj3uNSycGEe0AaQPqhVLAg1EP5xVOp/3LIUdMqHcYsymvQaJGk8rE0pp
aOZJznaEqxNM6ULxr3g+9gVXbA/4tn2A0mrnwamJ6/6KR7YjSQl6D0H8pNxPJO4uIaX+PfkPsBkP
gzqU0HkOYqGVHY+i0s4ji7boRC2+y/GrwnhSz6LcBkzl/fm6cI+XHslC1kPPcLfZA30a0kjLA4o9
mhePH6MJdcg3sOF8RRbuTq8nLrh+EhgjJK8t5QTsfZ2jEjTwldwcx9DEQXdhPNPnw1lZtoz5MB5E
qQiFFO22qw3lxWxAYPlQ87gXeFSr3VqhTrzYlaDbkVGJS276oT1xlkawMri5KPD1i+DZYBRf4xFX
mlm3IE1sI21gUy/lMTRvOck9jh28EcknNTy1uWXbrMGm0mgHOGUE3jcYeq2xdAolz5lPlZDVbiDc
o1LpNTEgYUHmig7Pp9LdKijNWkSzfZ7TwMsNXqjoYhoUWwL1PPVKcUsgiAHJetKzkYkBpCW/pZ/9
3qBQ6Id6PVohyrLoA3gAFP8f0zxPxO9mnfQ6bl5M8Mhg+9LDSkt+qSftWQ/CUxlehpdKZBgRICFC
S1GohY1KoMhGqDVAs5DLCOKlH2Apd9L09xDMV9ybv4608scMPC4EvgRP3oNoeDUj7zbmOipuPMSM
wfba2ymt4fhDagAOaXa3C87kqyv2aXNY1BG9n7nPJmSNoBCR3QFRe3kI9FPfd2xXb/ANKnTl8s3f
jx4LhN7Qa+JfkCms0TB+kwB4V9oET1e7LNrEXV/0HL414FNTo72o0qBKjf/s1wwmQNdxUtAcRcOQ
RGvQ5mUXGx76D8ADIq1QpPanDZzpN1YrmAJ6BBVr1MNSmDDcWGeC1RMAr6ZYzcyp9HaJN/m0DSxl
GSqxaXi018Ra9U2WLQMlkQjOJdpIHxSQT33B51A5rIQ9T0EXmPt4fS6NhU8pBp/Ky6XvwzFtgitq
8LBBhTF4ArwH55HOxWo4BLQFylbraAr1FBwlAClx4DDqk26qU3lvCBxswIvGruSjzs/G3kqxlHcE
i1JONOP2kje4wJJcpI+uQ9UIib/9Ft/WT1XunCr6TkPQhDQ2u1ZlolE7+ojgue9byHCq73mGzzEy
Y/I3NKuBOHZeQVvT51+AeSuTTEKc4VzxEouUYh6H6uCSwZgfqbyrp19biQJXt/IwH36+yrzMx7dp
ovrQZ0h3oOSHfVK4zJH1SIu9UtLvFNVbbRPYjZbnE87dl2MFEZyZpmWz/W2b+4NsKTu3fpHicTLx
z/83dKVi8ReNX6/TvKCgzkGVomhPjKCxDI3oPEmuJCvwMGIv/uRb0Gsr8P6E7nDBkBG4OiixVDVS
bDZupab7BEdH5WhmB8f4MWWbME/7yEf32HYO1yh6NUFqLOzQGVEIKtbFtR5UuUuLPiu0x7yolCMh
wQrFqYVFZ+QW0Vp6p0ByjoAxImcFewdbkmhNPBzZ+1k9P/QoaDdps1W8Y21WD/0+VinVeKFlOnKv
57pmcmVkDuc/xy45hjLl5g0B1erAVByR2dUyaR8uOgRduft4xwX3WQkGbenjKcAIP56YsAZqI20N
ujMKRzCI6D+//QkK956Z7NEmhdRxg1Yb1RsVPCuN69lYX0ZFTlVcKm+erSBZkaQUmu8FyE3tImVs
C+rZV2/xAVlL90raUN+GbL+o741FdfldqWLeUO3hsNBPTCBV/UQXecNUj8skDF8zuYPttDEhpd22
85tfMP/IyvEwjRxo8GJCrDKZbZ+eFulEdJSCMTVSnE9DKBzfYZcji47KqX8oQdtL2rozk1XQlJqH
VzvxaGm36IDpIAOQrVMeT+6tpDIG2/Z+MtaKysqyeUdpsNrOfQMgH9L5Ac1qAh3+7Cz8PhXgOsmq
PzCrNZ09f4AygxpZBznx9B2zPXXl9+qWpgwuRgB+K1yNFmsVFq3KEwrP0rKX80B1u5kcQ/GsrZ7q
iwIVhOXe2vXsGm8KVAHiTPh3VySSnOSzqDsoA31xYI5DAEImcfDHxKLBxzQKVj7ADThYNrpKeA07
vEfHjNKfmzttJTy78iTTtO3Ino8xpbC5RMnFIICPxoxz87EmRR9evijCItTjGaRuXRJVi4NFIUSx
yNDrW7L9K5AJmuCSVeS+N234DlxSO89oAZIRpkjWy7QrBeRcaNWPrvUGYHuR8e8BYXIElaSPT6U3
zliExMiCr8WI93mwugnx2lpO5WvEtaW727S/l06ow+NEz5v4GoAUo/CwXAkXxJNpFfItrcKY4XCQ
yaMa7ekClWzw+GbkqLg7b3XKWqK7d3ejVLehs6JXq3N14rGRPt63SHyrrV6+swNf9O9Nynb4pXf9
HGSMGKG5F0bBlFdbrzeepZ5Fo5eILy4AldqYBpp7wM33325RctkozMvmscTFiitFszFImCnpAOXL
KkleA7iEBWVH7MpFrDEhyhcLB9T5LVutbt8XEG6qGB/2m/iEO37NiCH6hNT3WQ1yVguE9+DAjMGg
TDahttBp+1V7ku/81U7v6nhL98BOmnQMcl25VD6M2uPlhnIA7p3OOo7gOftKY/GEZE1k8FOzec5V
xFP094UIiyQlYi48EX+STqg2UU8OonnqkXReo0DGi69cv+4L1NcW2u0JLE0vcsrMq+sKcrfwyoqN
zj6iK0v1L9bKus8TfIZhC9ycEzi+EU2iVDo/Mxljtk/tuugnrYqmHaZM371AXRLc3dUE9h7MPvCE
MJfEgrQ6r4gLyFkOy1glSC8a9o+IsfmO1X5UUejGUM/opibgxBRQoGwv4bPMk8OIOvbOE5rXewRz
nx1x2olxFdBBEIWukIBAC8NKA0llaYwcf17ZcvPL5/zRH+VkM+/P1z+QMZ+S32KCJzKzS8fP+Dxp
QSJSy/8SvbecJDdreq8q/QmYRQC/2M6br5rL8dFQh+FPAqmDuHhV5yA4v38p6sPQz7Zx7K5YKGqr
ZhJM9oMErmWreB+lJvb7jd39WL8oPTKvemnFrnncxNadOS9EeRB1OeKmBTdGh8JzSrXp4anZNTaH
xaWEc1UIoXh4IUqqbStG/F1b8V3LbAWD+erfL4F5fa1nXRMCd0olC3BIpj8Q/IqfTXHHzqd1JILj
nT9UqPcsOqfAnf2xT8eKnzzZSOTWkhedM3JTGdxbJosMCnLmTYwaJUCqpzrjPayirwQnvijrA47u
jdVpLyOvhK3/x7B3XhXj7+n2UdquzfmhelzO2PLA8lm1BWaUkvgrmuWLj0CSo7sgE3uylKcwUR7p
VDADYQAn3eH3Nxv8bWasoU+IU3/R0s7k4qkAIadoEshH+2CPW7R9SQ3497DJTrieT8wC/y2WK8Ou
C9UteE6GBP9/xj8pmO5HkaP3extX+SCmRQiVtGxeq0uMyM37CEPRwTEkhe+yqnRXcST60JPRYYxA
94DGFxWIRvRk3GhKajEmmSAPM+opPMgmw4rYeadPcYDiKvVsbFLh1xIMbEWlY8rPEaZzKGbRkdmV
zL2ENXZqmyMK6wpqQReben9ILO8yjL6qsJaNpoJplaV5WjqfIqcYRLP63cHbd/7uUQa+YVHlpsy+
5STHaM67seSJTHVCRq0opCsTEeMzlAH/4ca+/AW5phnZUYybIwRz5wCxicJq0xt06GYCb8ohG2fa
T86hd3x35KkWTTSmKrlGXlEUsyV19MswRqQEhC7zlB7lRmbkAbS2h1TH3LVvFzHA+lQfP3ZdP6YI
MXI4oRZAlKcaWT/2dX36oWnVsxc9qSrGLqhjMt+fDM/gHwt+zDqjKsgED7+1EraCrqqAwiFks2yy
SghIst8ByHh13yy5VfW0LdJBiFibpNEJQEzzn1jEnPIfpGHiZb1oZfE2uh404YmbqZ4XjfWSUV+S
i6RuqpkI7eGGqsfruUgNpa0GnKQRENHvLuBAHo/9NL9QdrC5c52L1gEaKEb4p9dhw4B2X4WpJ78m
/H9/aKCqemIKQNtNCY5+si6acTHYaKPFiHqbQ5n/3iMsUfzTF+fWI5o3rlHvnIqyaHk1CgCm/BgJ
ZPMXpFDxbkd8rZQH7qmvn5VRDUiYeLjbWI0uA6RaO1K2ta2NaoFhzjf4YoO7gkN6aKyhE7wP5kvr
dBSyZot2pJ/X7OY6qEPMb2DyjtRn279lI6V/TCF0kr7CZ7isvxBHu2b70TExhLk7Nkuo2/Gv9XCd
xo4AD5iJZaXzg9Ud+UBWiUTfAl9FJQg+Is6vtIYqLmak4ByO8ORvdVEcpf1xYGHObvLMFyXd0BMw
RmGfDydUa+W62nsLjL029jspRDq9ZDpiSC5i3m4aIJiJxQzf6LPKamMj4TUm+j+1D/o7HPxQMBcL
yQdz+fqTpylaOhHjPCKi94bLHYfDyMxKKMwVuJBXm4nDAFnKicyWjSynfYHMcr4paFqqA3Cp68Zb
kP63qY+zlGzW7j6cmC4BISicWeHeuCMBmiKEL0o2/gTH1pgu7dsTuy8Y3Mem7iK1jchopmmmcGfC
Da2EP2dVR0I/WoMPrzEPwMq/H5Cg3YRXFsKrCcCTckwsWbGiSRSvLnYgAnADb+yx9Qp6T3B2loS7
mBU/sD/uXRDTYI4rZuKSFPBmN+/YJMzeBw0maBp8PRsKEyyBtaPtPejCVEMxhPpoXMlD2WJj7m7A
Jr5KAsOX29OEltbeG1naINCxWgMMA4ELj3WbOE/F8fZmUVkkPn3zvkGQmCJmDYMyUSwY8rAMe7Oc
PoUrAlmsYs4VaWclFvYEebAtBaRsrhE1wVWaqnodap+Fspg0LIle+MxR6xYou5IVg3x4AueovR41
7mgkpNJWGYMaS2DEMdRJZ+rRuych+fxcHzYmp4SU84SXCjiXzm6nPMHa8Edo0fhxbrp5o6Xd6euq
kL+l63UFtULVMRV6TQyBgNtsk9egCuDXO+2XmwU2SDmwv1BxmqkarvPvIKzDkeSFO9tuq1iZZbvk
0KW16SstTO6tFF9SlRtsjcQurvVtKsXjpXfZ3kXbwngBHvERcXLVadQqTKbxJUcUz02MhDOxIxpO
5opV1ejPE6DTe3wwrdkSqykE0BaJaKHJphjuD5IMAOR53C82Jgry2l7RNHJ2Smad8L9THCv/mHfd
qU8v7ShuNzmCnHZ1dVaOlUJMEtcbm9vtcB91hZTg676SXcMBurqJXTgZpGe451/ab3k9TXxlPApz
mrblYc1MKTGaMXGfL1B4bhVe6x+Y6fHhmKcSfJ3ZnqkpsWvjZ7xXKhi2OXKNQNpWsYZ2OZ3qDnmc
DQzK4szC7ExS7Q0qEid/UkU7MjHsIn+olK85QWSNbmyiWAGYMMoyseIwKHf5l+beyEuxB5/8/Paj
CXh1YIRdHT47tb5mk3FnDW2YLATRmiD8Kb4jPCQFFRmS8W/qCa4bQpVTW+KBRnENmk39jM94RChA
4ayN872SQEUcjGWXN1IX/GHdXplQX7hnjjFWsRh7Njhg9unmTEFgWfyfczCz06qJjC6pk6d3qFau
fGv10CAMzQmbwFQytTC2g9Y3SFZbDhvpmI6UkXH3vFQqvAVtQwdmwtrKU6/akrzSBXMPeW+caDON
Epp8Ye4hhJ5Z3Aj8j3oTiomUlCxgUQzr2uB6RUQQBw/sHm8IqH4x04gQzbtThBC8rWZFX96WSFye
tWSItfYvGTb9/vRh2SDgje0zh4RZiE8eS7EutAmiFr1Zu7sjIsHyiFNiWx7xPyQ3/OP2kz9/l8WF
c+hHtq2IHTrXtQju0YHJufG7xsaOLN72Bvi+xU02t1v4p10kNjv3U01Jb/B0WzJRaR63plG17rX6
p4j8dMtLqtE9NdT5HmZ14VM/KL77YgIOxpc3ngw4sRA5VuPuLFfd3uRw9C5hJpbTFYRy+tX7o+ju
32g3c83hGzZ7WfrJINiwNfoZfG60WPhniJjBV++vRQFi3QQWXdp7m5/N4UC8HCa7PzSPjlImRzF3
urPzVCds8J9Cz+LCSd08OfyupIXRNXQNq8UBX9kwTZgrElZS+WS+TBTDQHOlGJ4d++Vdo4PsxCzC
CT3hnblpF0T2PhweUwM44go9SAROEIVtSxBfpiUpDpkum+CcyphFbCzhOC9ctZxqTsGJe3sMlDsC
HdrkGBsbsDkCdjbcuKuW36E3ejuOZjwTDnOKrASmymNeXPEXWJ5gCfzUwdIfVKduOZG5TICHww/R
dxS9XNFSKVeG+BhTE5p9BL6Vs3/4O1DL1LYCXaurVmqxbODaN5uwhJFUw6DYtMb/0ItdMmtM1UI5
gM+ahO1aAkJmOU2BirAqb4IXWI6QAfDjQAP+KP4H47touMp5Nc/wZSU/kwRn5tujOzIl1nugt81F
fE9LIRk4GXMhaU0wkQ/ITRaVtt+MRErg2jj4oEq+DRQqEqnQcUVXoanil63Fknw08wfHe0+X5eO1
Ntw/3YGvRz49ekF9EcU68t2Iq0OjJ4mfvAVP8gwhs/EfTHRokEzlzCDjmxVr79mWS/kI2XPsc2vp
y+AQ6POXD/Pc34hHRVoAT7ruh4KjYl6TdmQ6AY9hANhk7CtAhV0h7DpCDtSeimboqEE3ijPMw7ds
HGPomGPPvTVUgW6n54ByHDUEZpP3QUe89rSZ1e6enDMacdhrSpnziRKNHVmM0haiaHH7qm360AK3
ZhzvN65jfe7t9Iv4BvtmrkbQqq4Kihrzox+JnoaBJgdZzI01ncu65bXF+FRI3t1crxDVSShXy3TF
mCMRURg9grOly1lSpx3kG6cvaGNogFedBNTjQ9haaYRZocdXITETxvfwhsxvqFE1M/SLVnP1tgU/
PRKgbuNhJL5nkDu87T3I1INSvyUWRN/5DJ3P7zdC5xY/t4GN5I4Sg0JqW+n6qWYFp7nhmst07CyY
yKy+ngRTTn02IVOP/+NX/CbS9TWEZ5hYtcWcnbPyV9P6uN/ANYUXBCymg45rVJuFkSpmNmgC07g0
Ir3jCbfn/iwEG9/lHVQ/R0h00bjU6zXkAOr/DTw+6PQ2t51AWNnC+M35pxPVut4heT1mZrLSceIT
0pcJm7+lQe0DhAC0yK+Ke81Yfn30HQ9EVyF60GWfpQ5p46hAJdHlxYIO1tvZkVg3KXaVZj+ICy8X
ziTyaQK6X0MFXbdi0t/F/FqfWekLLhGC2NO+Ak9Ad9IC5vAmHOqWBez3ET1QUqScpHDSrof/2tq0
aZ0/Vd65UWTmn2mg2FV6oeqe7Jzm0w/tmoCoeHsOl2JyrzOBfCUxJTAAyimjGBQnTDtUrD0wM/kj
A7i//1MwxM1+FAUyCb1j83Jzqg7rTLY0c/XNe/LY8b7Mq5HTgldOswysqHJndhzejBElNRjy9GbE
6fWSjolQBTeVyE04WLqBQ95CLB0RUXzEu8uJPjFiIkYbQBJWYmgg/RWeQKI2x35Vz7JddiBHQvwS
FGJ7RokAnMDHA3VZrtcbyl5vYiMjYMozijU26IvTe1WdqyfxfchLCmDL1ApjdJIzlXkt70NPn71l
UjAudBnkAxwXBIAVVlO3mIE4zJSH1ZNzbHIMtn7e2fO1goAtgGOo0FPmfugamlYFykiEImhLVvsw
j4nJ2Rc12S2Dwr7CpDtEhXuK+FUoxbgk5/KVRtB2pW5qe15HHEBLH/EO6LxCUTfpQl7G5qSAlFHt
dAbTldAQ6DTLphCUMyO7fvztpPAONFjNN8ZNDOnshxUzOGMxtvdwrcNmkUMsMsE8+JBzcs6f+0UX
/sfTMG4JY2y4yEjKYPvHy2vUtKWwB5lv8f/aS+Y3DborzgMQO0vQqpwJQ2AUNT3qvK8pFMit8m4d
VnyRvkDdaBEqEpM7LfYLCnk9NXoheogn/gK5PBJZiuqI61T+t4XrwUp2Y76/f9lErUPPIEzzPLdn
EYCEdaTwiRCdswWJcUBlJXFUcC8eGMtaVx7BxlJVHye+XvdkGGeRNrQSLbPq0FCfwJ/or5tUmHqU
07VhJtQ2+cDxw3cH/uaN68ID0h6ZYSwi1GgPPmzRqvjbOxxfdWy4DrIGW9MJG+uop+YRa5nbi49q
5s0UFnV2XrpiRcM2gb6uZYguXmG9zxmfAc/ckc9aXOh2+BX0Mnfp8iAeQSMX4HTz8mg9hm9s18oX
0qMpwqwP1QupiyuYVvPSz7uQLgATbziTDoBkjx+cog1azx4sRJQM6EUnwfKbvErOEmdQut8u0M8J
kvxOERsPn3ugAnEVBDVFmp11q+n82s3EE/YB5t6Hlhlb8oMRtmB0889uyFlnN9kb6RB7Y3uackug
N67uIhQqSBFXMoLceKHOZOy5GVrbH+RcMrlGGxDsdmpelARTAKxa3CXJNbOd8AsAk+q0FZnLSqvF
eCuU8P/RcmDZMMajQkNBWH8W/5NH31XVvU7Q/8DZ176DaOl7ry4ZPEpiBpdqMkH/MXcwY8UKmXKU
ARZTIK49L0nYa+92JCDLt0dePnTMLEb87+gghdR7HYM8yNYV/PcOOAHQHhmCjMBNgn/NWxk3+XxE
z6/EEWit+eXxqx9woq+RNyNv/m1pIUaSTmgfQ0O5BxYTAslGppDz9yezKrwK+98uTkcPOvc9UtkT
5lp4dsTXkgOYrmIr7wltz8OjQJ7VA7h3HVpsSwd/v4gfOc4R0isaFvhJK4lxj1d8k4t1KHCT84yu
G6wFOPZGE+yp9rWPvCcKwHbImKCrpS3c7MsftuAoKh+RJ0gdCRtiH1CcS7KEWX035PcjuA7t2m/C
m4vczNNn4jHppkJ0N8rjtysnqsSYKqEeC6arSeOdGL7sw2f6j+Lwf/Qm8xVt/T45Aq6LPS5AQ29g
XJVdINE4stwE65PKB4iuCU2bPfiWO/3RqvgLgz4BUIcFi6ed5J9iyagd+18Ob1B6Mnm/pfrbfaxt
rAqCIj2LHr+vJN1gfSgiENfPQKKi6FB7sI05KqL0Mz2NOuuNJT0Hy1Vmb4GQyXnaiRKWJ5mjVv/9
QX2jVF6HhjQPAGsDbY3yv4B2W6GmnWmS+f3ljXAlR8iaA3ldkNd/hpKSHxm6k3dv64wO0Sn4vr9y
aYP89Q3Hz7oLRUIZ/h6VAVLe+Ye3aRr12qTvaPgpJ9XRurJqlE3bOWgAOgU5jObDDaEic2uPhjeF
XmkjrVc4pzyskEHaXha+xFDec8TibUsqv+0Kd9ovJ4kQwGp022N7ppFnNN4vZXHWqzwhPtB8ruM2
LytHKCAugOkVYkZb+VqRgA3Kw8WLibLwj0eoLtQEzk0gixZGgmmGY4pWGG+9U/mEHbFepkQAchv3
m/K6XKQllBJ6ama9rUMUfF2+/Y8Yx9cvrNyrRNCdT3kPeSAX9ZUqj0SG1tZnh6veTssf5BKHsdFV
pInzd52oBjN5AiVF30FqImUOdbDqsiCujhBARcilFWb+Xv+6X2hG8yr4wGkPM/uulkLupsxqregZ
hveLkVGd9GZ0qpg/JWJAPv4+VTG9EdKMPuRSnotMmt6oyGe2zwjXMv9XQub2Vlc6kCUP7n1RvSvy
xfzICJjU1k9vdrF3lTwv5U68UvTpEWNTa2rLFuJ6X91l7wT/E5ddg8Jt4bF3FbtrFTbJ9/oc6zLX
wOET2I3UNw0yrrYv1RcVAPg2xVQwYzL9Ddx2KIuqqFHZXscizFIihFVTY7GozLjIegUj+Fiiyilf
UrLRN/AXhXh2hEAeidqZE8jjBX19o1oAxreITQh//5Qo26cYqaxTDdBvOlJgzWhjVsgJqUjyYyD/
ETDiT17VWhp0oMjhF42WMpl2rDZ1qneKrXnvWGVfQx4gIacM6EVDxtRE0tqSqDiKnTUhrZvlY7Kz
GZhU7eJMd12ZPhInLGTi7frY1Q9NjU6lvbszpwo+HLkvOAQx5Dnn9azeSkYCYjZECdvZCEPgMBuX
qFaZeugsot1ndPHeAmbp+Nkq6gLSf6l45HDQ5zYGr7ChRREaPH2SjseItRD045Z0nlaf0oHp9cUi
TDVYrnurXBpQjhZVx/PaTZio4C7xRbheo1ACGPIlXWTGYZN7Von9yb89oobKq8sA/2sYE1Es1xie
22x21Gkne5Na3OEh93ycXnLQu6F0YLEhhJwX+pEW7QjiCqYtQmon/ovbtAIjdP6WyIwIQWLTxFIj
fynweW7QKatT8iMani67zzKPMd+0L2ay7/MUaKxyAv3hqWiPq8ypMZM7K4EngmNBiUcrs8+4DrHh
BsbjQtQTeiUO/OaPOPDuef8G8wY4ekV9sOtJ7tmmDz8ffTE+FZhZlWaGzNdf+HiSDS7MKFEN1mNT
t1OXyYeTgND2K69UrYAjoeRQIMNFpQg5O968L/+07aiK9phq5IC9yyw47Am7cYwrMBYUGoVYxPhY
m5WivsUKDkSB4TczIAMGNXMlgJtRFQx1V9QS3PgX/2GrKprdqaQ6I1vDJA8u+b1YJa+5brmqkzNn
Da8cAc1BVBxJnkkcS9yfJZYFmKTpOoKXa3my0kagHJ9I+tXf4F5dMU+W1VgwjHkXWhcvnzDZPxQf
z19oXl6T5TwgMuxul8ozjQ8/SdsaU1XNE1j2V5ikvYecvH9EYSfPi8EO8+EuNCv2EKIyS4GSAC2d
QmAPTwnPjXUHbGePIEhbQZ3thfrkvi6yVMFofiM+tx4iCR9nna8GK6d+fzDlJesiwirDP1o3Q/u7
URP9OKD80isSik7y2Vg2dgaiOBpLXyGN8ZklVKo5TfOboZ4tYVrxrRYukccQnkV568bFQRGKEJf1
EOABjJokQahRlrMhYvx2pHsQmG4rNLvDo2qp7TLpOU45uxNslZUQjCE1jtq3GRk/1Ha+gNKv254O
h59Yz5EFD1rvTVNbH9bUKZPDfw8XvVH+z+L+FgeW+XiVv2eyCln5Xk068tnty2O4WhZQRtGsVomu
jTL8D1n6sMIrUV34poypXdja4Cc8Ch6KshDuqmVMLFpbIQXNX7AJuzxB3TFM0NNa1b+Zpx8kE8ob
CiTm3C+e8Q9KAKubw2ugE2OegwOdWpF71M8QiuXy3P3oByPF7VVgKZqvLa2xgK0eo4wrZsaontKN
8xCauoc4NTcgPq/mX0Uq/oJ6QgTPDF3B5IhOHP4cGzzV0gRJVqPU6Yii5PCmNfIBIn78VpI+blVh
eA5yR3F0TIOKJsiL/y5CAAklUVy/YmPfu5Oqaokcz8q5hj7+e45jSAzNxtvIOxPci274p4KHlsZa
XUAoXz/+6poSpTPMBG0TUcIC8l5PFrGp6ffxbfrq63/xWthv3XDjd8STwXjikRY0XIYtmn9fyfpU
AQSOHeUMiOSTfICfJVDl6gI7i5nNBekhdkLpl/lrqLtZfdf1qpZF+6DdxQMf2WSX9n2v7thHGwuT
DrV7QSjTaqMjrSPfAJi6EMKF3g1ufcbo8lQlIWznFQI1wSbZaxrQ1KMmHe/DRgICFh9nevL/f1PF
XJM8qpJgIXQEtJTdSGEV3oyrelIuJ4uwfGs0Z/k2wBHw4cg5W0rM3x5HpXXblT6pGC98SlSCq+Tu
IhKTtfF22cvRbnck0BmueJO8yREYVZU1mZ4d6MKt4WbIGExVM5Bmp5Z9ivJdU6GWdztzpvannlzR
dAl2EL0mFgc7U4oAW3ywxcTFPrj9cLBJF24BgAsYmiQLBS3Q4i/cnkOFULMNbvfRcyaf8VWi0BBq
vAHfnjuDpG9R6XJf7n2Kto01U6SWttSN5Pe4NiEDhk9tgxuSCOnZw9L2NYWjHnUrHX+Y7mHQQ+Jj
X1YSgjwZQoEtFVMmeddWzwgWmpMSwvzr0VlDV2lgJ+OzAp+jdo/QSDr1yDfx/IlNtm0fJZvMLf+i
9jq4soYXTOcpKwTQLdB+/pkE/izF19WyM4lNTOjJ8r7O3kx9XjcM+CNIAigxvCRUwxnpJcWgzm5r
IFkvuC8aemOlzKwNs/gk25aSEySv2Whla/Iy9hoyzAwczeFsqUw7H1hrGLJgSKWkxpwsgUAbB6Tn
uE8GFYbWVWgyVILQa5DJ8fhcBEo24rQXmIEwIAZM1kFyaNl18fTmf7zbU8UCmtKVmDYTsT3RfkDe
3XHCsKjo/XAeeXk0ZD9Ow+cj8LL7ncpWYSDkAalUAvVV0gryJSDPQcZwpGQZIShXyFizxZZJLyIx
bQ84chV3063rcHd+phk2f5JaTwIc7b9BeHz9ycmE2nRuYDDFO7wmFN3x9ad4u7aUoxeNT390mQIu
YBSE3ei1uKjcZfqoq8v2GvAVub2VHs4EexkvlCI9QbJ7b8SNGhbsPAtHath+lMFBIkbLMv0hr82p
LFdShP1y0m2bDITLacYxoDmpwJ0EXAquOyXC0FqtDIpHLyogshfFJLQPvsEWouS4OWZfjUMnzpUZ
exT6Lt3EOhvJvmXYi/n80V+sp6Ys0TIrlUqftNQjLc14a8ymZphpwH4YKI/JZoIApWYlC4X0PwD3
rY0onwNjUrHfduQcXDgPUQ6BrCtmKS+7VAChbB+ZsOAyeGzZlABWzC6d+dPrzrzXhpCWb5pYn0G4
LGjGIF7cyoupmOT4bOqyPYpx7UwgjaqdoBmrUgwI+Of1+5Z50FyFC2LIRkbyfkLGxkRKNEVDfFau
orketJ87rN9qEViznf43MIY9w2+xDBqCC9s9ZDbiadp9iSKIIuwtGnOgB0sDd6RtbDRe9opCiymX
S50p6BG7dSNI8BRHxuC+D+l1pwgvzYZX0N8lAj3/WpR7wjpui845ldkXoT4f/zrDmK3OD97dOegG
bFIL1hAgbmLN319+3EtM7UHlDmLuE1P04jZjOt4GI98EoJX29bCsAjO3C1m7LU8soAcl4XxCG3BT
qRLvG+XA0j6iv09/1uqDna6a4g0fBrwLhAwXUOZ+auzl1eVYZxIOr/LddKBDVivQ2TLzFzEal6ZH
IKqulMs19q9BhxKnWdpXBdF9pQ3+rniQHKid+1EiHHk3bxyexCMnxXkIOuwZ5MXnYvoc14yIqprN
hE4NZFNKufOYg3lHEA7bYeayVFItuXdpKfzGbwx/QmzpGaZXO3J38sH6xJTaZRolD9cfzNBILRt+
df1JinND3N84YlD0ANSgGKLMLow0tPQJFFL7B0MaT+IDvb5uifIyTK0EFIrRyg+0SI3HCSHUt5Cp
r3MP7X2r/CSvUP8TtPHFK8BJ2sQDGAJl02d0SCVZcRzelKEni6KpjxxgWdFL1Rdk1ZXBQ758pYFx
g8sxCEiFqyaYsERyuRJp9ZbuVeFLCdxXDHapbzFatoKj2roytBz7o7aWLT8goFuMMuJMPIDEk16F
hAEQArHh5kyD6tJkI+KLeQY+z+COHzh0eCkVcJmfzo8l3/FCdMhqtIB6RDA+8G+eLX0HnN9iLQgz
4pdWXkEtUnMMFSTnHc4o9smsMgz/tUypnoCyylY1fHOk8r/WAE0jQ4P1qj9eEaSFH5dkJRUHqiXT
Vq3/AgCytTEJzYYJ06BcZV1ls4qWQvGGY26KFw8TDBfINeDuMJ5c0jzT6EmnykPG653e11b9eqqZ
N0suzCH/OJXFUYp64UsD3bAddxCdfziRffJXKn6Dkb8HMS40P/NSjrhAVs2EfFiA9m/57nERcR2j
R73BQBqaUYwYhctasT7O0ydDlI/i6PUEjK/IoJZyl9imGQKbM+fwTaF8FtRV8B6S2HAFUW3nHxn8
2n8XLzMgpEuBxDVTW5ivZdqnr4RdpoxQ67faRX80Erz3rJFGFkPESiSX1KubGwf7DNtJ99UP8YYn
nfiT+j8Oic8ZFb4nB4Almq6ApnOUUj7F599aJIjZbV1Zd3BvOFS64fnWpE3lnRQLKaFTVxkvvizN
DfpjbTMEXRTRhtLFVbpvjQ/CKcthnovvdB6xJPV7cppoh5SvfeDLMwBxK/pEAXXGgQRLs+OTWdtc
hWAaPsjx1Bgjzs/QFdzQY+m2x8umz+0IIUdlGHzK2PbCaMSQZPOLE7lcFdsFOPWxs/0wrSiyx5Lc
eREYy/llouZPuNP6ZImfjvIyt1qBZp/ZT3MbVc7RDsUYWp/NbkzGoLB0bA7Yk7ds8ExU7qnhdyY/
Uw5brIZvsqRBpwoj7k86XyJTT2XoaLd8kMBkocaG0WoNT+eFIJxOBiLUCw4xRnnQlQ8AaXw+uwy/
y+vFI/u+0C+diHRlWkEByP4pGrG2Jn5NvYVJQ9y3DQkIH+C4S2ATfW8llqRnnMFAbPGiK6lIWC7q
Bw/Ng6wSyY5ChBhxCgWxLWZ6quXv1MRsHK8yEt7G0vEHIbH+bsAfeXT0b6phOK4dA8HaiOlbT2jY
RPiuuoTvoAT5rgJeAvNZu+eTeYJYRepKkkd11gCpXWTteeqZmbjKfV2FMbXmhns2O+YNRt8mdQif
4g4hUDdtSsfrVxKB/VveC+3dZud4DNJ/Q0Sg3sikcZeQAd386LXMTphYTpo4bVXpFdcbPFlUUFs7
VQyPNU8e7SSqnh6YwGsJEsrwxyJg7Ua7kr3Gj75HL6t0KldZ6HkY/oYzgbJzmlc2QxWvoK+r7d4U
zOybNWeJzi0WO9JY0ldSWXcKBhFqgZsCxXy2gPYqQ+QH5tqM7UNkQCoKtd+CQwfP/1unydULBldT
pB5DrD6KNqrtnjRgMzQIUBTKC9513uYd+zf3Yf5XJV5HOPA1Jgdzlnq+5n98qD+bMTd1dyzXyKjf
1WMBAhcyq/tdNLcdOdIQcs3mjggG08R90gjzFXE/oUcV670/mzE30TC1UMJmh8dYg7Yjpc7gES3R
Xoz/HZ3LRLeHPmYXAZUUL4QUzJe1rJbE5TrpTo+KDLJl/ps++bGBDpnt6LfQMA9U1sInhhXAMwcU
F7Ai2NooYVK4SflndjeiHQ87yCFsBOkEo5UuWKThFyv3a6XXKFYgmyL9S0j7oz1yv16de9vbBCWS
pCT4vKxaNcbEjxuJ0xblo07en2vKzOm+BjJqWJCzHFgN5Aol2GV7FtnHZMtgWVYjUoBG0aTylyZq
Lkr8Yy2L16rOPRlzufSQgU/8Dt73URzvQso7RKq29f4XLaBAPEjpIBVNszNC/BVO4h0xxq5aekk8
9/r0TFtF8DCBvT1eU7Bijg5L3jFtYM4X9iRaNRGJTU58el+FZ+aVudxFAIX3EvPmUsAsMw1HLRS9
7R6U5enOvGufnCsuJFpFqdZbiPRsYO2IrS7z/HffvpaFkbeNMubwzeZXIk8RUY88pZ+g5rMv5qem
ssGl14UIgdhbyxt6g0QJ0Eo6GzchdqwTYOxn0LxScgG4LkTp42XfBHbpN9j4gY6yRso8FDqjwO41
twd+TWFBVshRlYn5z7C85DpHdeAHRqomOJLqAub0FSQIIJ6A7ufKWGxUBCl1f45hxN/aK8Swbkf7
2805PDvpOT5UMpNqFASZkmnsQvvK1P9cVa1YsDKAsQztKfh57MW5C8JKcbQPPJltD7GHqKXZS0BD
sPNPUqbwViTsMbkySGJxHIliC9PkogI6LBkEnPxXKFJo4Ih7iGsQTLJFjTyTzccVA5Ijxwguxo4E
zuWJNtpVpOU7IpDDcR18aVY/Ak+Z+K/x1Sz90Kw7tL9AcGxeVeeccZJk6TpSWN46OdunVvHbP2ok
oz7HgQ7lEL087SichjYBVEtYXb1kd9VSkSgXFAlBbZb3FvxujJ5q/k9GqVt4bvNHuRwqn5z+UixV
iA+ubobzeEiK0uUe6rz7pkcY3naPvr65Pidmzo0BSWXZXjmKnxLTEGcK8jsjK8KEiOwzq+mU9W/W
QOpCUBg3HMIdOdXSWrU9c9tqZ0lVYx6yzeNKzr/+Xt2ZBD31o2ZoGchMLTonEXonBsHXyTgFM2Ng
U7NffvfSwGdil0VQo3qjBNLdJHths8myo1cL4KOvI6C69nbX3AU1grAHDpCk6QubDhNB4wI8le75
uL1pn+u/rCnZcg3ZLDzlddWnTyT2FhnCIt1gfdySWLV+kUgQVHVMeURNTTo0AVb2IPpQ/0Zj8SWK
ld1tvzoXHnuxCj68PMtql6rSpJoc/g1NKPoMAftMvekHNmwffCPfWT7HYl8I2BXZlVGc0Wv3Cwfg
K6R7NVMr3XhxODV0Pcb26RTSP/xoyghrrdzRY48k/t8/gHxSrEbMmWm58DOJEXlbFYt+f79Rr2VM
Rej625EoLTNzoPxz3lG1kMKEaIH+rn0Uh4kg9S2Zb+d3YCNq0X08u/uFQt7E1ZSOOLRL3NN3chK7
DjYiDmJXdo/tiYFqrZOpDEMJ9Hiqi61eB47WeZhh6dOYbdVoBtEraitRXeXDVv855r0Bi5BAZQ2a
2re74UjPIj8H+VKbjV3LOCUiBQE+xvhb2aFCWDZaclXGIoniNQjX8NFJKR1Qs0q8VsmJOTCtTsg8
rbf3PwtFDbGyWxvLDQZ3LqsbzHjsY0Yh4IQbA9AgX5hrmTCnktNkfPcYbM14Kco8RWPCYh1fHezA
w/do6G6VM8Hqf0vdUQXopg5qpXMYskp1abTkiZgECUENFJN5gm6kZg7LBWgGxXeHSwoqXN0qL3Y4
N5SuZvs9+oGthWHtqPw8hN2i3ONSO+kIW4oGOESRd26TSxBIdaojI0CxRzSwOwyjxly6SjZEpSAj
LyNxwSifTzgDZVJ5lrKZvToACX8ccEEZ/UEEiNPXKk0QC0Ui1635vozyc1aBMZ6VMQ/vF32lI7Ud
KOu1Tq3r/d01aQJz1FUnay6a/EoiiOFd94/lRbVor0PZffBgd/fOAyB1TtPvk/6lDrgMj6ceeiCN
SRPUrEf6AUx6pvNKGPN2iJQeqzrjhzeIEkXNl+8Fkolb6Bm+4CdNJSXGFAWDYTcYlGaQHe81otpF
uoauKGDkcb1BhdxLS4f8apeByaLdlsE5lWalY2/CYX7s2CSA0HDq/FU3UUrnTjGXaFIYmN69OeY/
z3LbrIHimrRlgsnDChJgelx5nvHiUT/lt9+FFckIvb4bo0L9lewl+UHEOq8YqIjq2QRo6acHim9D
TlNIxPTi5xuD+p0UUEstXCmwIXo5QSSVZm1c6rHNs5HECipISO68xwbfhDCKKGVZrVREgtxsDgPS
jjMPHdIfiiK8gjv8HavHI98Ix9Emwi/nvcgiU3NhgNjmZhxfKnjrNz2kSFY3RihFvEBC7rnjms2e
o0eaGzxRmpbdp04y1otTNr7+RDw63MEyl9mpTQJWtQe3DTFs2/dQ5ztDgicPgNbgeXeNsB7STkHw
QPtj+a9TM3QNJFlLYjzrF85mdHGruJo+POUxm0pdYOexlDGvMrLEwq38kksXF4s6hvSD81Er+jYy
ljiu5dSCXalMvNzLVEXktIisPpFLBrvCb26SPQiwt/rgAF9QMCli9Gm/rr1HdYv8ZPUmjx05CNXt
tZPOoAJV+nWitFXDD0u2I91xMyMbp24YO/1CFxBX88y2lKzZiMlXpZpHYT5fSZSag089KMlUtLiY
BfWdEtFTh4xAt2SerFZcfHhG1+QMbooo0EvDd9u6meF+T/M31oLqzBHZTNkfdHFSPlIyZ3Fgwfrc
OErasOPM81EeDJLsxR3GFawZldqOYY5y4OLSpVeMx4m5IZkNPN0upOOGzO1TEc6ZlBLy7oLcN+vo
kSJ++/nBc8UreARndOoUE4AAok3/kvypY/fwlnAD0T3IQxPx2R3GgGc6egDWWEw/1HRWg21HED0c
nENOrtDy1NoWJucHq3DguGAXKkNhe4LpkXBY/eohACy+rueSD5tZBx2uiTchmIw2k22pQb5dBZsI
LdsUJz4MdaPloMoY9AKDJahcdAn0BfZc3uRSxPQuog2SZt3Fi5i+bPamTNSOS/F7MtvUKw49hjim
uK6owijO1Ljg33QMTqmr0kT9r2oaRQW4nBTNtAbPTvsTmkCXbyNlM8GTPaTociqXP7vdAkBHbDJX
4O8oADov5eQ0t8T7RsW2zDE37h+I1ANA+fnkWwzi3GInPRZjAdboheBK7cHLfCKGCwFN64BV3hhJ
Hb5VVqfZmepVGHCyz9ZT8bWmrKbw7Oz20X6izBJ7CupiGu88aF59Sl0hgyG9IclrJpBJW4cAtpPM
FCZfJrHx+eDXUBLSBaWVvuIrbDyeYQj65KNiga2SFeYq/b6fZv1nUZygxYHgCK1214vY7j+pswdQ
7zOlvzljaCAj3X42CttgdiVkZfJM/DsmwJliPWVynwExt+RodvycuyWAADqzv9MQaz0Dqe+22pX8
TU9iWQJTNk31S8If1TObb1ApMls2RGSB5K1b2QcgMoFaleGuI86UJfrr09Nus1p2LxmrJZJ9AzKD
AeUkbcLCkTbgpvnwvtmTYJeDthQphE/Qo0cLUOGA3RimetAA9r+EJ+uxQ4J9Q0Svqh/uCRkrZw4E
6fmrs4L9m9DxYfVhbt7kMY4Hv6Nq8YuLlH8QdOQ0v/+E/ZFVVbTC7FhrT6pWGUIcukm96uR7hXy3
rxmOoU2qBinCjTOcsUIYajFYMZ8j+D0NpsdIZn1aRzLrmJ7MXEEwzcVDxl/t9gRb/cuG49xtXpdl
FATB9PiT/s+NBAyY4BuJDetQ7rCptju03yZYd43ij8ZzOVwmZNEq5q+69gVSgl1/cE4KlyVpg/uT
KvEkjtyJmncjY9irunO6xRktBJm7WMmiJnKwt41bdijJkirBVZcBikibSvjmfzWDamclf94BOPPr
ca9k6ZDVBY1m9vv5e53LxVysYF6MGIrJmsaVhZ365C6SGcPnsdg/mSzF2+hn7WOzgVRW7qt8kPhb
rsRNfbzrulZphM4jHgmCxO7EqnZ4eXixDbHhJ7c1NW9TFW+BVUGLGLXLJbROvTLJzNUmI8BZWJ/s
P3Zo+IKo1+cX/AXvFB/+XhYRMm5Btd4uC4rkAMqAfC9njXZd9ZfCCsX/MnjNuw4DhWrhBah97/cw
SZi0pdwIUmwpKCw3aa2AxF0+KlMksxdaUZWVREQFIakDLxBhv+klhb/K3eh7+k7TLaiF6ctlWWKV
EO8FLARA2t2bluB+LANCtFdGiL+PpVNuDDMeNcZ70ndd1LpQ6tnv3ICKFUWIxwhrtzuveHhUa16m
G6i7zZ9TdxdPvARwBx+upk92Tt2d6hgiqVTrucxMmiFiGiAFL6mdHSTOBYdfLXG2Shy57p6K9Ruf
881cxNMPfJIYV5hK+n4pzQWDzFrLRqChcT05tNPSaNmAFt5/0/t6ONJ3YYfhJZQbR82g8j3m5+4z
ftAyaXf3uKTQ9z05PlzaZ3sODVN4z+pdWTAqMTjslJRx31TORmkw0G6OuHu2o+35LC47QnAJt8VN
rjeoGWkz6zcb1M9aqe6GCtZlQqLuhxwUG8SgsCLyta5dcF2SmsQBR8tMelYtENedfiRo8n9rIHib
nGfyyp7m0BXUJQb9sobaPnQzm+y3ZDPlnnxG6q4VCbNHTeN+cONi5Opx28IwVfgnXRMzVi9UdDUN
PnlXEnvIfcEcYYft9U78y6zGRcmO/az2GE3wgaHSO/VzgpHI8Vok9EX+/xePQ7yDh2sis2dcG6gE
wppvHSJaK9lqmG8JIFT3tZBzoBDfL7aaqbzlpHrGrh2epeSBZEPCAh/+4Y6p5sxFzLbN5SoOGnTX
ntEtrX+FDdgCRniM7/f0aeSsIpL+2oJykWAok7aH8J72sxw+Gewfge1zNDcBgZcDzz+lPlYFyyBw
zeLO2cqx+ZgOC7OaLruW4TJNeuHUHVmoxBaEvs5iu/MtnM1TV0+jg/WvDhI1xJFCidXfZQUbKfDB
qflJF2OrHMYG/5Wu6syzx93MEJeExgOif0pESicQOEpg6V2Bontsf14SmXuGyCxzdLno+26DIKHG
MIexDQMocUrBXFX3vy0glbSSPScTiU9tn6tJdjiBPLp71att/6ghFnlsHLSY16XQJkZ0pAMox87o
bunjZp23fDKgy7rz/6Fk9/JFneyxTsDmMpYF+lPiGOGOa5mxpXcwMRfNu3jpF9aTCSt02tjgecuR
N8GeQwswjIwUVbk25yzkqh5R40HqG70csJaYP8U6HIRY8suX30a6I689uNLUsKep5vP87uOm0qKt
ZN1HLDjbVMxZK4rqoUqE6THDoHPczL9dqQHdWv3qpyAHwdpJoITrVkl/iVufFbEk6HEtKhzMatzw
bPQaJNIvFqCxSWS2X38zn6H14ZtrKjsuQ8BmWZaha664WYsHAdGmGmvLdDCIwI80jSGCBgIJiFvo
nGqo+KgaXshM3AynswnQlDTXybjmyhr1ihTiLHSsIeILGq/+lGWIizkBj61dw4h2PLiqtBNBvnbZ
qiL7z27g7kKZghuSAMlxybdk5qMCz88AAKB67UZ3CeNYJ8+DBzGLo0YK1LRSfFyY1aE3VrAA57Fo
n01PuX6SzRsd++IbAv0yQ2T7ch7uZ31aokLkCjO3UNdG5YWEr9eYH5sdrOS+095cb2lFMwXRCRoX
yMSCFtujNHus8+RiUUOz9GNYxRPe3YeR0XVmVCIBVPN4PShiH3USWUn5p1ON00yjHD3lgFv4oKx7
nuboK8jHTFmropjBvX3LXsipJhVtOwOPDGcuafVjj/DAE5uVBpyZG4k0e7upgRM9A0ctg3Js83T+
mJyMzcx4b6Ey6+angWEgyKZOy1e8GMzoDXNCIQcRr2TSzYwTwqOcguSAW1ha79HwDQ3uaSLrgDDe
u86SCbxyf9rLcAq3AHjZ3Nx0MuWfJWtpzOHNNWu7Z3YfoB+4HJXI70LCFqVFsu1Lnapkd9Qs9+0F
xBohengJrp06VbeeM19SFTomLlAtXaARS3DAvaa+jP+8xfWOiREYiavh9I6eC8yOjX9jT3yGpY0F
rwAxpgKu9gp1YlOOMmlEcqvN+UczMG3SfR4a0Lmn0OAa4J2ckatLrqlu/ebcnkeqWpsE2RZI8SPW
wbDvabPoj4+C/K2pqskI04GOqrHwnJJIwbm/k8AEte73d21YzBw1PdTrCj4aJwooKETXysaus9bW
SLyV6gauK5YAzCpdEBEJVaDUtkVFFsTn6s2ScUYiiYdtBX/QgzjNYbO110caMdwZV7LLr0nCufZ9
vtm2mUsm/9lt9yrv4GfV1TK2nL3sJ8RHW3dUE2363rq/XtKeXkDiHHM2kZgRCrpOd2breBpfhnSo
vmiEJDAL/+pnjRgVV5Va+5ZMMTw6p4CSc12fUZn6NJPWtKpOOTEQi/xxk2fKThAaKSqfPnXUY3ZU
m74/d3us0qbS7fmOL+Q8CFMels0+dTH4Ocv5aQYD6PiZBnYZ1ogJE1BU/4J2k13qB7j0tNZrmpcH
271tpWKC2X502yBalbZ6/GakZDJ1hQGwbw+03oT7yH3R/5tKqfaSnsjwYZ8BUFDpMCuTUKO6eOJ2
Oq0RUD4/J9NSEG53b8pQAxfM3f617a+m35S302VhD2MhN2EtDgRIWUGQoDagCbKCU4J7axGOexa7
RiW88ccMVqOdMP58nwVS57jVVgsfowHqmZZZNnbIVLTPAZC83Zm/KYPl5RAFafB5FcQ0aC3HW8PX
IVcSu34KtxXJ2Mgti7h/MCMSHKBe6hSSTRyz+Owkw2Ya8L48IMOyscKsGK0F4Iso/CqGnWMGOHjR
0C/sh/l/Ogxx/RH2OTrFJEsCuu6NBekX2+B/1eFpDlsgvn4jkp2iSHxzsJ0kJ6wxPW3ngmPfV07X
N6Ks/WNesCaIi2mPNv5enrDeusu0VZhr1H5bgEXSBdb8FBunqGSPaW2jao7ihuZxo+9xb7mmWZnN
57GSyQPzUdAwoVj2k3lWP8iwi8VXGc9XDvhwCFroi5y/UDnOVok8aEao7XrhPOYpirNxCYvXFSE8
oruMzIlX30CWk2k0X/02FWXggIIwuv3jbcBLOt+GePZgeZstmi9zyblECeB2TOmXLYNtFUgX1qUK
NDJdeJeDV7DJI79f6SVY6u/JPa1ISMcL4+fRMDg4p1fFtctxQis1gS63Za93Jlrx87TwfV1OeeSO
17afpW6iCmbTVOCm75IHRE1PwJdk0yynlaUQzI9Rva3G+jMEdBSUtakUG6z+tvgr1c8OWLTLG1dq
LoluPrF8Ve5ZhtxA7akNp4LmFoQj9v+2myg/vMAiGDSpDoZGs7moPFE5dfkmjcof1aV/mq4pq/t3
rjoNNTvVdY/A77Wx0WVa7qxoWeS3edBd1HxdiN4uruHsjNmJ39wDULlvdVEVFPQ5uupaRMasFYGP
cIeyLN8VzvtJ2sQEBF00u2YKi77XD7AsqfoPimv1klDtKR1x3DRYGZAgrcLwaaexRs+y+3Mu3jAT
HCJ+L5ksIRtByTMRngBcftDbSmX8JURJset85wY8kt/MASPILvcucG4Dp4AXcxscUI3mQl1ebYOC
riOdpC1YA9ZqH62QZAI+o4BaqBkPR5JCn7pL0/SWNddtZA2qLRPe/zgM6pF6v9LIY0UKTvwVUP9D
mYPPpwwf48/2ps+T9zzQYp3O2qFwziutIU7XAWDL5T93z5Yfdazbrke9H7e6D5qSytTO6YR6yGNS
9CRNr8m0Pt1caHp5Q6J7VGC0ErggjZyFLpNzW+sMz8eCeUwN+R4yXfUdaWhss9qkyJr+2nSBFJtt
z6TdcodTX2z6oo7z/dq65QZK3e0JoCoLUK7kQsftreDzdI4o+RUUYpllxB7YKZDR32jotoMtd/I8
bPWdDrHkvZUFmPB1gF+xMnPb26xvseisovek+f6YSmoRXAby3jNokV+NlZh4o4SB4wBpCkxGHo3s
givLB6RnBjyEZljh+7Q0vjYTHXHNkbdh+6aEr5wxfZHpPWjPJTpKPEzIbdBi1dOY7M3iYqbfxXxg
WmSpof5nS6Rh2+Ri0UwSB1By3S8R8yR8v7WI1ASkrnyZ9/B/jtzZa38FfWxWv12m4jQZNITsasEn
sJUnrB8zlSBwGXo/K+uAd7cqaSr/EmFwGEO6m0gCxc8adImNbWqpAmf/q2VNtIACUF5q4TQcwl1T
JSYwoNahNKe91gtGax7t40VdSBDR8EFZmAiVNsKo04kBpGdMx3hAJan0IOj/iUbbC//Zl3WKTxUV
70x/VPBhuTGeE2qfjnb1RevibJCVVc7D33MKzz0njJsqqBUswCTRfVVvdvjkzwT/16j2HlM4YANJ
q4KO2A8PC4tuOPrEKdRGZPj3Ix2QqHKVhO2yqVxvH8RrRMDDdwT78Hm5S/wMlB66kEcNJW2fPNV/
VrepANWzvydQ39C7owQPdgy+2KX1s6hPy1NjEVLj0HuwwNB9HNMy5lzNdLdYkpLGwh3xLDGPs+dD
YWqALRtl0CSRKfc1W+Be5HTqKw1LO3VB7ejOewXN3dsdQJqio+LwzPGQtIbZ9Q2OCRj0GkfAZmkK
S5v0kIeYyrTHAUbCrHv5evuXZdJZqglEjScX6JX53UbC9d79dv769qtai8xOs6vyMo+4bR4892KG
4/3Ny7mOGl2pZBHT8rAOxDphWhEUWmYpHwysnC0UpBuknLD61STOKXXNO8jY/CYRwZdj2HH7Iyhr
d5n1yBH3i01cnsvNLwQlxc6E7j+Y+fyEy27YZlj6a8JHYGuuilB8fUf8mjMCzxJxUrEtwsTlWdpE
Kcp11WuW2rB8wJR53k6RSGqGK7TLYvRkQ0lqrxARUeoFi+pMB949qY/ZF/Lme50+VIshv0Aewlhn
JoxICIyrw2K0tbm6Vgqrn7SYZB7oJ/Vz1Z1Rhuj2O2MLco8JcqlKD12YeQ5UaP3hemWzYUMOpzXb
zuO5is2lJmjXyjk6zUy3hSwmNxrTgnu8P+6oioyfxyIBVvHfM661xa2qp0lTujKcYE1vTkPKTAm6
V+KsJex0VqCxf//M7zNsGlP02cRS1ekvlP/ucO9SGMhupC+7N/pVw+HPj4yaWvzPZeo9zFbcO+Zo
qO3MjbvU6AciOgCp4IDlfPtxHf7ifhuGCbjSyneqVn0zhWpc2FjqjVKCTRRGI/APSBQZj2Z82T9U
f/Iv7i4nBugrv26DI6qHWb8qCSxxNQt47+zZCxW5+rZEAr10clDpcmh88XXsSAlrdqCNT9Z9dhew
AyVKQtoG1E6t7bo84wntjiQC89QytNhviEhMIYZEzxo3K7LDbiO8wbmxGOyfZyoNeyhpf4nh6Drf
D1B2hzPJkHqYkmxEA/J1NM2alVDMq5dNwfSJXi6RgdECK1b4KdqNnV6LjOp+We8mf+nwHDsoBpMz
n8BmVoHJdJscmXRoLltwGKy8lLkmqC2DqlvFR6e///ND5IYRa/7rop7JvuUVK5pmvhMeeyPhjnKf
DjUGdjvJEqpmM6P/+F6JwCxhmCP1zA9D+JbJPMT3eEzihgo6eSNsARo1W2umW/B0Yvigf/OBGeAF
zwXLEdtxMTbOxak47nNuQvnoYzn8ardrzDTBu2YTHHKDTjN6Ea+rwy2fn76nDDxtlV2Qutzc+Alz
qqAwemUT6ChX0Zq5747KhhrafPPqk8ypvaJn3P6fNSRTVkbL+nWQ5wXqDrPRizMw6auBJJxbAhmG
VlpYgbyevMm5IAPM5inDDcFW9Rio94seQtWFDCrfyue8X2N4MRe0wG3YfldrOz4jEe9AhXcdvCD7
sl9RD2f6HRasO4CUkFnIdZ/FkcIb5+wtz99/WAgCzabyw0610li2F9zOzmVq9j3QVxgLCj5lzpDV
15rTHeErUQQR9Se1BZu8WrJah2jMgJgwITRWR8KMimaYme3L/gA2TTsm4sgtCqKvQO33Zzim1GCB
oettr8u6aohdDwsz9zUco92ZR+nzW3hom2wgINnvf8G8/THwp2vpWwaLDvpgAThlGdgW5VlXznwf
Dgo5aTJSmWgIlMTCGYSDvmJoxWCUAl2coAnZ8k0seQ7AuPG3r13K8QTlYMHdOro8rzQXhv2ardrv
S1Se4brFaW2v4Qz1CgABWCXcsmfMNuSSgKnfuL0ebR9qRvM20EG/h0rj37c5wSBRaa46PNe76lfv
8YDYixL4uSnGvLiZaEVqotkQt1JzQFrGJs3dsv3jnC+QnW0QXdBpsBP8Hm79VRYkuxqekg2Y/ndo
xtIPhXgbm7gcXyRIkQduvO7z/1JSHZgEaS1+exJXNhhEImgJCklyjHkiyB2BXRNGy3mRtjQwoN7K
Ahy+rWp3G3E2GWJc6+hAp3FnYQnxTkmuDEjd5iq54ZGQlRvvKeT86FC9myoyt+3W7I5C3jn7Pfwj
vbGLnaP/laLun73iBGQu0EB62wJ4DOaHOy3jmYrK8/3vk+YFyzSUf8eKtA/2sdQ6n9SYHVJGm+kk
FovyHCPKcMMZrAAC9PWTMiLuNtPdn2Bc2qZ4+BttY1S68JfvvjjQd1t3iTKHTuj58yfve1YOHUcd
us+3gj3dC5WacL1oUgn4oFrLwcMJZ+NgQFkO0FKTGhZu3P+5QFeFfl3bsKFYJ+P9dud3Y3zRAa97
K1MhRMRdqSmOA8aH+NfUiaEEb/EGZWu0SHjvMiFJ3aUpSz0SOI7ci2bhEDhUA+tqGacnZlMPUv4D
A0MqXmDn3it6t7o7vCmlVLXZlj5vVtOAEz6z/YkbUyTchxKauPGsdd6BJHKMLPQ/LSvNySSKsk5e
SVuMRA2znuB5MpKheYknQ4piy81Cyr5CwjglHqRTyXe/08MElPZO3xGOGpuTTyBpm0a8s4fMwxC3
qCSaAf9sWmxv8R1WYBkCQAVRno2Bqio4zWKcf3b4XdZrnvYZtreSxWnQ0c1kIXXZQVekk3jzxwca
CrTg8eWvEJ9NqjWks6r8P2z9IPEPfWkY6ckUSgaproqaLoGgdYRoAwyUvn6fuIJfiEw4AeCDSxcZ
zM0FIK+d+rWmfjyhQnvNAbuN0bQyKv2cwlaJdvMcLaDuWMKrVIiK199x0lKm04nx1HfYO5HzKQG1
UGNlR5ODhzQT7gCs5H1Dn5vEazslGGoMh+5Aqf0RqcDb4Q/SkP2wBGetHHulOGa9321TjAWsP5k4
M09k9ZYRbX9de4dlhqmeBW8cdvGvO6SDHOyOT8rWT2yuPbAtJcqG0pnrlkENeuIJeiCHWHoDbJMG
HKy7Pi14rTliHINF8LCkyoeSwCKxrr/R1WS2vNV+h8PFG14DtkM2wE1yd1hbh3pJ0PstN3ibXO/H
rviNqGmUI3lhnW+pZ2Uxvv+3y8jVC3+Xdf3zx7sa6lXXhezNn8rad0BGx8uULYSHSRr95xfkrLnS
6Uahxhh3hMZD/GqarTd5MmEb90LQSbgVHk1/JUYACG6HuBkzipI250XjuJnL/eXe23IffBWd/2rz
zUxPivbXnOzSCYLC7d3dhWoRc8ZlY/lj3c+/TzZhIEHgVL18xqk1yh5SEa2HbyTuHXGcPHX96kAa
crVRK7AooA6rcOjbjICJMsN/hIIpH61rINOnOF89kGq1Zbh8Vxf3Uo8IR/3gH0z0ws+TwyhYiZo7
VvBY39ygKoXVTvK4JZX2TIIZwFhhhOcenc+kmU9O2a7pgA8v0DwgSu7ENMgYU+PLeamFhL/OaRaJ
tqC175rdIjMlOuLlt2xLjTl9KU2XbioOWBY8gx/FTUojNEeq1lvynAmcRKeTEQ5taKn5jt9inOU1
pLIOSdFAPHxowLCoe2icVKEC/dzEziY9w7Z/vRY2Qcrt+egVA983ye7YyPYJr9+LYF84oYD0+ZDD
Mjeb99zIVRx0ZDUYwvOdQZjsyaqXcATAdc2pNJsA0JNnjgSBRLeJdQ8B4vFofEBJ5mPtIc2E8K5P
4vXOHPvXhtKLWY2cl50GoqITF86SHVg/BPslXCLyRwWepoBJZyNm+jU4TYvD4b67wuuNhQiLY+Oe
+TZn8A6hdsWqQ8/xxvX8pTWHvh1rioKAvA+FwNK98QHQwHUl7z0jHUsyBc3P8dW9jqT8b9B6Abpr
QdOJCKGrKy0fg21GB58+F/8YlvklHqh4BpMfXutif+vCWGumtiyJuiQt+ljZqV8bQTvmVdEeTTF9
Fq/uSC8cYeBLFJgXkSZITsMk/L8AdC5N2uaija9/RMFam+MuWSAO4hHMCBFlkZlNzAZEdqwOfhYJ
Rdm8KDBeAILvRG2Ou0mnO0P9efsU8AhBbdOXzivhlHKzCbV5dWJiWjTaQjsguY5tRE6fnhZeeUNu
d9GiEzWhL7CIy+xX0m1qYkGrkTSj8SGmXZuBcK5rXk6IgWCiwr08giL85QvFY6oPl9V6V1PNdTHo
XDtrHJgnITUMDas/QCbVoQnsnSwWXI4jkfpvASAUWL5gmp041/pGIkjlJDTD6FB6rXJuVAm/T+UG
kS8bG+DpW/N42GEIcczrgQeHkeNZJkxrh0kp4nRdtrAZmZZeMnK4+EZNZsO0mvOZbtlEnFbC5cFn
uvDBHGTIrCjXTvokRjzp7fHvLrA/iGgshaovhqkLbc1s94zTjUagkwTKTOFw9E5pQJ9vlfOcEjeg
xH9GQa+TZZDhGz+mFQq4E48YzpTMMivklI1AxZ3b9yDuFTnF8KJim1VgudM0ZUI1mE/VvYN0BLzJ
sgkLRhh9niodyn3y/NArHaeftjNgJW3JvaAzXq6AONlWRhN+bSw6kgQ8/KPggpoKudxbMPiavGEb
R0rP1Aa3d+AT9cqHPcYDC6t1zSSpHuMTZwsULWTgC7IpoGQGNRGFjJI8zEiauit9mIHwxNIJw+GO
KzOmGptzcy91Jk/0qGR4W/usUOu1zTFqIGCdj0cWcM9aYIhr6SdhqIdOpfK0V2phpvfphqqsr3pU
JWxAW/nllEEDpe5m9O1kUCa1tbK5q8gWClvmI7c5NiTybe+a11LC66sjKhxjIPtAN07bOfINkhl7
Ks715slPq8HZJQLvVMaAvz+otvg5KxApMV4KcQEZcZGDfQtGoiH/ycfD8cQABW7k/ZMllVerDs8f
wpOgjv3PBvbIjUGM7suKHAMxzQ8QlUgec/ySVZXLvAHn3+8V2+Q/WofqjQii8sylq750S+nTp0wd
eFsnGfHaaGR9OuLX70Y/VaHOHo3EGbe9Mi2nIl9MRODtquz0nOE+jvDMc2r3n1Y1li4nPATXRkZW
RSbGxVjTeODEv0RZuw8kg7AdR71JFc22X2674l+S2cWJTWq7zU6ILJm6ztkLPMcAk7vjakNMeod0
yZ4F6wVwi9S7koDsGIxqVkeJC5VMgEEPOy9lEWSWGOHfVDWXA3ujEY4p+a7RmQdAGTNQPE+mQd3l
TcYcmdGaXu27GXS9QL/uc8lFL6QeoH4rgGxLopjRqcll2F3/JcpaXbaqo9nZo5IQjgi+0EI9FWeb
ew5ECJYJaE1s7uGHOfKtqU2qn5hUQ46abvm3eM4MgKvy15bHPn/Y3FuN4EsJS+NP/IjTe+NEVMqF
40FxlKLh4cBE0sEkJJH/3eN92Qb2AjcNENhpUeB3qgUxGDt3OHKD5uaE9K0hMYwMMsOcfHzR9q0y
46qS5eMZiCjXCI+mFvE3jhvFawZ2Jc9fHE8QYP07FVHypPeMhGKLm7v3yP2jnPWJ+JaCFjxmadrD
1kcGAdM+oUEL614ChLw50GFB4pkrTF6nh26EL9lBLWang0IshWoa6C2EJsPEKHcIv4aa6/K8YwRL
uz9/IGtr5nWKx+Uym7qKXB+hFWx3tw/a25BDcbB6g7NqWxv1pQBanIEy/e8FAnWqRhOK7qzbZ0M6
pA9o8jq+RoB6dtfMpwxwIs4JuAfjgF/MsVCoRS+wlojqsIJcVUJXBj33N/tsJSwqc+kD4yrrTjT7
LfKZz3nksCefi5YscJj7xsyJL2xnKU6DBWDzGs/8U4ZJ1MJ8O5nB1tpXfrSLIUfdta58l0/3qc4A
CQt829FYE5tKa0KncdacTFHkB14LnZFaFr5sFuFyYDcnl32uxax0+t6/Pf+IDOj5Y2sO4Wl8DIHS
qCHiKoPjT4+BnKTm/pzk5Q+n0kRHQ+CAUETQlBmi/V5nMtpxHXbVC+1dR9rGG06neC52FqpCvC/5
sKR+nH3B29nYq87PAmBBZ20PFlx7OsNq9bGUhD04Bw4iK/oNFgH2nur02OIAahUVASsP92etUbkM
b5V6n6J4RYhfLXTC8yD05XFsBli4tAyAehFzCfJ8VF8sjZU09W+lsP3ufsjBomHNA3YWUPpaJftr
4QLilhwbn6lNvry8XRily3+52Chb9rZ3H4OUhXODqyQ7MQ6mSCuHdPC/11+WY19lVkAC1bsPjNPC
GWWFXDqWF06fdxcnNu12hSkhFtbBmNACK7l6kkg7CRt74Mxoh2ODioPnZnzGHPIoAiYr31cKQFzA
MS7JOIiAdy1fMCKDbjdKIXBWbWwm7aM7LktKUPx9fH6aQG6cVgWF23wc8YrhHK0hWyUKRHQ8egQh
4JljE8JIMlGGsvjqask4J4br/sScwCZ8v3ze7JBM8lJaWuqyaxEdLomPEA4NrJ4E6UoShnw3n1Ck
v/Ip/7rmu0PwlWCLiMtNt2eX4sl/hXtPoEVnXm3Hj1ALRwHMWVihbWq80jRK2naAWLvPNhKhLLPL
WbUSMpxgSVSOzrIHD/9Kf1y/MNhlulBvmhJCVwFyG88khIT0clZU+b7Kh1przE9yG90nXDEwmowJ
+Sp8iZnOh1pwSgzO/uc3vRm7azYmAM8HHh7qw5DDnf3P2QwgpyKu2pxdK9RoNs0LQIpAdMa/Sj7N
oLk8S4x5ewa05OltHZwN+29m98ts0Mz29CTaMgz9MzoTxgT5bDcCb3sY8GvvnxzPCYec1DMUgnRq
CjPSDACUXE+OvLGfCjAvwFvKuxkPXg+PKu2KqG7xWgpCpCjzHBkinKmyAXFbG7cMHaqn9Kr4ODaj
jZe6LR44EJCXEjMqxnUhXfVFL5+25GgwNykGd2D/x69X433O+cH7pt3QyA0kaIKf4gKH3LjJajTH
ciLLRplPmlvaEPgUKQFTQamHK9B13LuD1Fqc6Oe6VdFzTxAEs0BNpSLo//V48UxNXcHZzl5/LBb1
xHvGAClOEJj2cneBPxX4wVrk7s7wiROK4b9DvrPr7JBZ3PfuNqEs5qncWMyWbYIGhHQc5aBfulst
ZOpfTG190pz9psqWyCDAxbH1nK6kz1PuwfUgVWiX3ybIkiS8AYj2RnYr8la4VqPjSeX2aFD4EuNE
TXyC7aSyz+9CyHiF+g2ZYcu5iMkl1qNN9B2L4Bhnpr975sAqkBdyBHFR7+SFoitiU/iSmRhXK0Eb
R9V8fbuiFvMOwBOdZMKctDRGP4rl956WzNcF9CzhYLA5cuEWrJdIO9qmgRdqIAIJfvo0oPs67H3c
bMqX3MxL/EJvktQIypBq+2DlioePuEcnXIpUxCPyl1QMD7L0Fqp0Ai94FTeCh24yE+eE3xq5tdKP
t1FIAvmJ/c6/7xpgCvZOjPocwedTOMlaeeia6x6fOW82jbuSO4p80eL1Wr1swhyTLU6zbHc2ppAY
QD6TKBhR8Et1FIFRurbl7FemCodoQlT/FdiWmMr9it82QWaSMeu7AzdtJP0OeMFkQNjmXdXpvjnp
9i014hiWnuSa4zmk7ngzkZ/ZXzk+vQ6JGYaYyaZziu8JJjf/s9u4+6wwVHzEvkmO/ZK+Zed0F/N0
bpAFxz4Pk1vMnlv3bwGUsv9d2GRmOWgEEK1d9YJNbH4WcoF/Olq6ymEc5piMSIM2JiYLuGvpvv+R
0vrqAPsMQE3PIlzdqCuimMXLKg6RgoR8BQHy2PxcIBEyVLU8+uSBkjTK2nqDdilpdUsuv0GCWsLH
lJ4wfsRevbgLuBRrPinXO2elwBpDaHhjUwpxRba/VI7Gev8AITVufJ2oRGjwuGf3Gacw4ZMOkZxo
0aXhsLgfZk1ankQTZLDPQC1+hthle12OPZuk0TwtYneSCqGOgNCuPp+ATAFNpa2NNwFUT0K+9pdQ
9TB4qCMz+ceWF1ZoFGr6Ht9BVTum00rLZocNyfYqaK83S2g+6q2m3TzP7ENJghHl1Sd5jq9xmbvt
H/Ky+y/BazAmjK72oEE4+vJRjJQUBqAkN3svXhz0Qs24Yeg1KlC77bfyJheOn35mLNf8/FpCJYJv
7Rr8lPgQVTDmLoXTMzzZiKlOMWAkkMcY7yHdu6ggsZJ+RvhrkWgRXmLqockTrAZ+jn81qlktgKjY
rShrL+ZYp0JpqQr6D59HIup165Wb/5dfdJX5sJGf65zSUOmcg46bIhLVQi7Ef20CccQ8KZC5tihq
DUgdW8wfeIuGr3M3QqKRA06UNdjItL1QkiTOpF8sfkOLzSyR8+8bYvMW/hWOeCHz0ZvF2zaZmkhz
GrxCWsbvTG7H/2aBlYJuhDrUo4tjdU6ApxxX4pRDkur++8str4DyU7S7vMYWrDmbeU+pc/aM9dmR
J+kn3/PgBvvlhlbt7IvUsWT8v5rXYEyCJkh/SiVC4tyq0FQ90BIFseX0/e7m3qxNUTgVwXFX8XTD
+v5DbJqrK1F+ugES6EfqK3pYTtw9C/PRSQ3ES/oyLlNZJqTmoHdL9CJXYU/2DUoSeql7Fszfu99J
33tWy7LXhTWxYtGuQ+TRmhTjUCqPMCtkDcCaAZTY+xaOOZ0AIMiEtBBWSuOWJg9F48oCIss96mEW
wREFd4aqPWWAcVFuWzUXq/jsLYfra5y9Fa2SdSxUiyAGRDsYBgCPz4qHpWNVRVtBUPeEXuQ102cE
IetL2Ov2+J9qKnH2yNbPqBHqKFbjbrDJgZz1B0lxcxi7laErf94QQOVzvoEnvajX8e0JpkTneHBH
oC3t/es91gXtCnsNZ/c1N0XDLG+RMR4pKeHby0i95j5PM2VVAxv6FnpgtG3TkoXpUxcU6Uf172H9
2nTckd/ky3KqA+tw1HrHdRG99+YeBSIUT6Xrhm6xiQn0zsRp6oQenw1w/tyCiwmxlwVvOei08akm
/qDA2wahM8cl4dSRbFfUTlu4sx/ZiJuWxDz9u6KEy+ByaqtWO8iw3u5loBXxaO5bMbZgHrppj+Pe
SofaqWz7+lxqiLcFHIafMDaz9j0VIs1d+s6QRDaaA5Q+D/Kuo8RduCNY5AqBDLaDllk2CZwPGxS/
NQf85bzC3fBBCRuq6I430HPew/Q03ffFsFGEjzh7tvGT/Ms+EuuEUOfMSj3liJfqJGBYAUyviKmr
H8XFy7wgHHgXSYXQQeR1j4jf1SqUM5Y8++vGcfyBK34+y+UAWWfFRi11JpRTp8icL7RHrI+4ZEke
BkKdFJgEpeqEwA7fdQdyBE5kBpFHwUsnBjPyKpBW87AMsVzLvm9zo/3ncM0uwumiWyi5lGnHEMKc
Z6BrhpGNMBXBtG2pLbA9CGQVw9Su2x+4rcUEFY8QN9m/vjr3j6cy2bVuB2r+OaB3i8eTqgZex52O
qGzLp9cph2yEU5RgYJaFWO3o/nZ3ZccBJHKlqpTDI6dIU7LC3UDk7CUKsRCpik1kLIa0WHkm7Hql
q/UtrIrOw0jhy98rS1oKyWLsbzzJ5yttNKDJ8+eFCr8qlWIjIXAHJ9WjAPS+axlbL5Gv+LhoCS9o
WmjEkrblgrwfx8vN8xmb/t4sY39SUn9EXZXmhLhEwoyaaopSWjJxnevVloYx8qVyj/bgb2jk3hms
QUIbszMeaXhY3o/1LnDYJevB4azHinum3sHlsiwkEjP24XVIEr6mrpXwdu/rGCOE2pKjzUVnACHn
6Yiqu8nOPgWJFkQys3nLAGZq3WFJ7wii+7BAui0vb0n5kuZxRtoAtXntvwvYEmWO6GvItB4FhQKN
tOoL04fCASdt9dgDw7h8b+X6k9Kr/hsfzLocUDtjAAvEgM4e9zihlVvYnaAiDw1D9a579UD6SEJ1
o+/2p1YNp4D3noE6nnCZCg1msvdozxC+VhkMNe/BVwU8EM4d6PLO/Zbm5PLRAEoPPzzUmhrguCx7
IsGJeX5c+rpGY41l0b1/oH0HnCyDYgVeUgqN7leb/cy8wnHRqbXJCr454MFEjMqo8fSSvh+k5xwY
nEezIkW2PhlIKAABQrCTvhQiJ/4BWATBsry4E9bZiZnRedqNWPvzCdlIiU8cOd3nYBBe52EOGk2h
0qsOA+o0FH4oOg9gWiqzXuSnYO4nmY4ytihN2VbE1a5arnKCpV5mT7UrOjzg++I54v7kezwjzuo5
t8AnXQ5eM/5H6lHpPSbJ0Wp2ZyDXveifXNSorPF0KHckTBTiqb1oLZMEbdPeU7oJr27s54IQTK0c
f7Qmn3/w7jmzmlunY05SbgVPsPBt/HPGPmMOo0RhRP0BV097I+8nZzFADwue8TxM+G3gApSfDYkS
/LcoPd7KL2NWgWeTWAo2ql95BENPfx6wkVUy/X4stYi2ZwiZIuMcPTU2QrkDxDEKmo0Ys4rLqrLe
f77lyww2+3acb4eufOVzWMqZt+ZbyphiBO/yzgKjJ9ZRWa9Y1R2Minyhqtjwkx8NB8F700nDgIFt
db2N2DC5l9AerNBFcGIYGMHKqJt/BDbCRPu7bRHq3sE3f73xZQ6WWm8Ql/M5G5ft60NReSspSwH1
mQDNt2Ezuqj/HtJqFDSD1TODzdb2+9KfswXgCWc/Ifzk/4QTNJCr/IvVOrKAZOLIGZpChSzhakOi
dy7OLTKdXw2xbkG7uLx1oUjlY4u9HJ1hUxKPGs7TWqHkbEj8oq9vhOxp5M2szk1mLtJZDNw+ZHbu
N42GIR1xrdL9LxELLw8xoNaGe6GEKfdfXwe1wS0vGeb2M85yYVFPo1WhcVrr+0R14kAwmIboVAJA
fGzGGZxIYrRVu1QJOcS+aBFOtT30PwTLWv8wk/08GnJKiSF7lZT4WyXp2jXUA1WO0gsF9z1GdA8i
7xl26h0GT1s+hYrErLjz/APvH+8hQ1U4KEMWD7YUrd1ZWMdIoXEUIdQqvIwYiGLpjJA0AQAifvWv
Eg2BrP4aV8Z6kaExDsCJahTBLTkrB2I94jBpAd4TS6uHjFzu/nWPu2so9PYCwlCstG/XaFzupB+9
xD6S8C8wTE/RctURHRy1ZGdaMnc/r2Y6BleIA6YnUadt2oSS4S2UGdC4wa86Je4oHVIN+Tzn8Psk
hgk/T8tF4vuWX0OaiumSCIQExMvqCBK2J/dnVeI1lfcvylbnMq1oQa9TImgzN4oGMtHVqKWJo9DM
7XPjO7vCGHjK4KYka5MZajgCgT+jWQ3xqJePSauRVaR3GGn/PCWsr8dIvETZL+v8/Tf1AbqgXfml
ByF5PRADnKp3nNuyg3GZMdRjA/l3hTKn1rJFT++7TOVxdtLXZkTvD0cguDGCUN0tKkj1EKDhOK/l
OJMSUDlCTc6ArLrpkXfd/1yNeV6M8K5u8ZRmW0uRZvknFNMjMQoR8GVz7bO3BDXKkDZaq5XASDkf
VxCmhWSEAQi+QUCPCo50qocrFzJGKyQl3m2xcMwCXVO4w5qxlemZENS1aHTcR5nZkaX9NTLKBe4Q
a0m7PB1/stsaRpos7zDibRmK1zHdZemapUkNoXjEqIVTxZhtRZtlrhegpFXfIGxxMonasSYs001W
fnKVoLk4XyrWXoqUJwNRNJNrsJkfqg9wzb9WZUoT1z3I9EUDAZTFofv9r/0uNRqw4HLjaTRo0AGJ
LnPPW+KxmKOmwuw4OXDc7ixHntk4jz69fLcWuiWZTVKMIwzaE0gxsy2y69eNKSoF0IM5S1tLUkSt
uT26Sw4Vq5Fy1bn2obgTH/tpYTi7Szb+0+L+11R1dWqYEFs2pqSVF+D9PRW0YEaEDiN3/wO2qygd
prgjdGlNJUgH4P37CCcddAbPeHIThH1St1OM0BWwmvJaQ1l4z2xFooUTYhQSJI+Sb2VNL1MvqDCg
+KbmHO5jmiINQpeNzKiHGn6TgPS+qV5EEtSXpzDwV4/phrP+dXyvywNY+TKFDvrmqrpivCg/NOj6
nQB4CTdQQvJZ8ObQn0nXwS4uqGVZ5m8hE+4qdGlX7NzLXSWdNuV/PTqo2UCWki6/Cy3+wTiJAy7a
3bvMREYjal3q62uyMAgpR7mylm7Vjs4y5iJNMU04Ztb6txDuf80AG9RJnUjd4Ru9BIghPL8SbEsL
u5j1jMqwv/KInQf+fAQjtQbnJeQmjoQq7UVDvenHP4qLpmJAR9Ye1feCBDRt1lY4ynR6rrDMJ+ND
sRefmrW5sSMuueAuZqmL2krjpTIU9q5+hOVYGgm4qoMF015KD1W9Wvl7l3cwjxFjHzxRxFTJ9FHH
MHAi/mLhck/uIbcggrxXAZFkBFWDUnbrsTutA9XoNX8t+AaHtirrqqtvQBtazlS7iW8F3kjHKIO8
3wYbJsCdoxY15IFFZIRe80hwIe8BStW1gFPIflH0/3IsS7fvRj2UG1ShoX3XAJ8I7J2Z/IuNz7Ou
muyKL5UQtcACifMjluK12n+8heLgzkXArJBsHbKRqb3vkd4CjvADKCbFafYnyK5TYUCF88QGWjlN
nPExaGvAF+GQ7p9O/0nwOmZQCTuRGARoQDXsNMu1Tq1K95VksrVBigywy2pGehfnrCnXtM1mPnH0
0wthfE5IqOJ3T94xfpf8KCCyNVa+w2OjQ0M+JztrMD37CcCL/hhvDSfJwSMDKyopXiL2WpnBqYsB
pvyj+92pedWySXGDE7f7UGkvI1aIdE/qmoUOZedh5hf0yRuqkUEYtqfDbzkJkYYB5zB2O1rtff7J
UYGCUjtGwN1/q+qaYKmSQqtd2z9Hc1Lp3/K/CiQM6wMFPRBmkG2K8ZMsDyynmm+t4KWj7J9iEQrR
eKerJ3rIYuIoFdBBvZhrjgYsugSr15tZ9AAWwipB5MKluBRSFXhyU3sRtnfy1lSJ/D6gW5GX9eXN
fcpW8ZqnDZsxncEyoVZdgohwwv9Ow4gBNn3BjgejRMb+YO460PjJaZTdwzUO22cN9SOJ1PHTNyBx
ByibuEuYCKY7WLpWuL/Afbh2WzcaQELu3ExYZ/Q5BwtaJ/Xr9WrwDaNqOG/+dv/qTDXYJgmOASRl
R8oxZYvlsvkZi56R/vm7aaYdNn0CfFkXD6RPwQp3mablgljIROxlb1ZjhuNctZKdZQ83cRQMqdi8
xlTkVVsPuJARCveHS9sIoMPGCAAlf9HB8a6AOfoXmzCgBXigG38ogLvu3bu0Rt6BDEU/JQRjoSWe
eaAerS/LiSfWZ2yh2doXf/Xi5PQxwklI6gMr6w5UmhgSr8UcncSJ3XeDo1KyPKquUCs0PzjlrYWd
CrLb1O/pcgStHHrSNhI5JBPi9sIOigopm1Fv6cm25ormXI7MUkVQJSNyVFb9Jt3uhe4iamc+Lwmx
czL8Aid3r0xSAqG4yAm8BMlJ329LtwRtgnkPpgNzEb+S1mD+yOK3nW7+c+i5RsZv1v7tEjeinSV5
bHSEtMmHpA+5oZMjVjOk2o/Q2N0ZWR8kiWqXuPFzkdAe0aDtDCTqUWNL+s5H0Q6Et03LxZSQ2spB
+DYZoJ6a9vusiWeG8hp3gN5ZQPzc+ME0cZU69Z4fhuWLAe2R03qno3/5hXv0eiPkAP/dbWmpS4q5
VKd5bwtpc46sItsgD/NrBZkkpJTV/92SOCpK0/aZIjPZqpsPmOsAMrJJGz83tIlNpwZ+PhcfHHsN
JJUgTon/F+4UHnybTa43T3uJJTQ+DAFycch/H2GTnS2irn8/c9JmE6+6SpXAGG3u76ygsOtAx5Ky
WpOjdBnU9Xu3OvST9tp0FuEcwhdKxEheC7hUqzD7i5BkG2BUzCVDfzgCupMUVwqDMDF8ujZaQnKp
e4Xe81YAzor1FMdDllO2NRrTPE6r3y3pk7s6EjP30oXLG+ubNhFTDZtRBBKF65wQt8aXpxr8w81O
BCpfCifSNy3gsTC2StVBdKLtHCMtTrCKPjUdP/M6X8UPcki9wTHlo/XAiSpVXcqFkzDJdxRZHVXp
Lu5DZmn1hex5kCvFHA4DoplEVJ9OSkR5nYC/z0OWl3Wfx+AIQeyGXDzeMTDdAiYQL09wNi62QY5r
CqgAg/p9yNGK2jkqgZT3KVaOUwGsOdJQRxJsUhhkGRVw2WLw0dOQ8ZEegMnwGh8N3+pNhziFCuQz
5S3hMuIbqFVQcOf0g1NFsLbIAkxABRQa/ErPWZZcHdtYS9USxJ/WQNU/Cd1ayUl1ACNgVniU75eV
YQFzgtHjioaHJbKR2qUESv4j+tWQaJbr/phshL1TgeNIOLyLwC57LnYgEhihY2rU1Uyvr4dlf1Fk
r6Mzlx4WTJxEglK15Zz+/ucrRZlWHhVcRngvvCI/8guVsGz9HfRQizCVO9BScZM6vl+B5zEsVUnj
kgdEJsgdKjo8zAPPviDNi0sibcCX+mOAIMt3V25awhYUf581NQWS3Z5NpObBPTuzyiJMvsWTPUQY
Kla88vxH6f8sLI2KZzxOAn0NCRRY6C+Log+hfXPfYDfim62pBvYdKChme/O8g7FhHxsOEboHoN6A
MlfmSdljtwQvgXSqly3W3mclc1o8KD0ITcGdRSq4qD0FBoYT5nPPqYQmpWJilSrM/6i6hsKI5kHX
yu/+MLKjA0dGgYcFvcryGereIoKj1GvQl3bpMGUJimqfjTHVwsMcIjpTFgunwfk8NWSsJ1RbAWiL
lsN8qWVWUSIA4JXQfOe5vr1FcdcldDgun7v2aAtm6IugGBlyGYr/rbnn15U2kuTmxhN0zhT/MwoE
jl2ma7TTjQDEW7ihEDMRFXDEFBoCrU2DAMsvrcDZpfNCpjg+AdrMEPkWoLUWCx7JuZ7bDZch5W9r
Q/TeUaWXJQ558DKvcQwmgw+J4xoj4yFWfyt2o4t+zwIrXWbIlTdNmt0IuHLTyp1tD4yBnzq2UW4W
lMZhArL8RBkNl7bZI7uliFZD+nZgvQOP7lUnSHlRt9P8zHEtni83tCUIT3Z1fCVpvAW6NM76CoEk
2eMENnTGMkLA0bZwfOQJkRzvhyKLpoWM4L5ifrjksSZeZ5/gMp3yDGIdC/JrvLOpZhLVdhRCpMUq
RtTppf3LJmI/EKI8MOvB0Kx+G5iFoC7IBZw9MqDc2eYp7fzzyNX1B8uiYMOuEgLeaVtOa5f1GTlf
YlVIOXMfDDwrywVRCF03IW8P63fNqM2WwJpXPmzKfPjtNzDfkY2W4xfByms4RKKcuyhVOBPam4uv
YF6YeL3mvI5Z+/qVN7bF6LtLTiHe7YBfJe/l4yka1nlbPGbyxTwCWtmmcM+4fVrxOXoa19O9YkCo
ODCKYm6YjCtBuqhcSvOr/gVYMkOOTSOQ5Tuj1t+8idzhyQXGaQvz3gp055ZOU+/6SNg4yBC0Hsg/
bgDDKWonkjTi7skizKlU/ESxQXPD5l1xIsmnUdyTHs0ouQmgjtmtJVLITz8n269G0PU+ETR8ZT3t
VZU+MAS8Z6GJAl0sCe65fOrAev2ym4dlIQblWHdQZwMqWUXo60wwGqgQziK+GBJkqUvAdf2399tV
LzjRDYMIC6Mk2lNOlocvZ9Mdxfswfry556D3R/elvpWQ5HxK8zjVATzlC/OwExW/nY4lOrPSs6b6
w4DQkSscbF2R5EzhVnr09cJ3kcc9M8p/Ksqf/6nPsfEuSFb9rF8ZLKYUAc1jUXzRN0kVNEUgFvv9
fwbwB2Ck2jzK5T7MCOozTf/NT/KbIifVV0rDWCwT+SYO56ChvsR/hhFgOwOgAjwJjd12fButAY3h
gAQccdC/yYXzTkd9Bjq1jnqamGhyGK1yFkOtpTH8z32Qr4uvGbHjoWYwXYyg1yCsMQWiuZYXxfAk
NDPxIxYF18L1nAF/GvRQ3T+UTK/thRp5dL5ow8CgcPBLAxzh/v+DRKmCMNDBMNRoFbjl3l352nZO
GOHLdhcj4/N2ZhFBFlSR++TUSK12cFk5chlsy3tjW6tRTmTAJeFlfaO4pTuThppP3Qk7EgKj9ph5
sQyT3418791ZFV0hoAMVoqnxB2c9pX/W1QZS7tQmDlHwFEC+C6phoixo6O6BzofhopuuL47wjPsh
bOMHA69jgRL0IgMUUxpfPPn2hqs+kNkvNKeGryFUwT/YNgR5g2ZFOo6Z26Jcm4o8DXQxohyYPTDD
Tp312qpdqLY5B2UJltG+sfum4FGEVWXen9hCaoByrJMWM+UzfQ8hy5ujFULaHcrenLUajg1wlL0t
XTZoKNNgIRezKHyfqhj5Z+uq68bzfv/z88TMk8lOl9y5dKva7uT8Dv5jAm3BvB9qnVP13ts0+xJ7
9r5a2K6V6pMPBpg6wtOCSCQNJd+GXbCs7YWCnwB/kjEs8NmVPEtIEpDPdkXJimZCqU5W9Hq8Z/kC
6036H2XdXe6P3FTgOlO5cEMWm/2+jQpiAb33sFO1J6TPdiiUC9TpYKue+xMEkiFTGbJci+oVWkVD
9CAepjGuM7Sljpz179LLhVWdXeXryNT+P025gfy1ByWc/q3Oyv+Z83U36xq7w9YntUkTvGyjetq5
3Jl4AyXBEXvSbNni6s8MTlxO5EITATjNcrYrvhU/r2ziPxkh2az9rgqzexupXYRVfM+uKfIiN9VU
MLytspJVVuZF/Teoun+IfrG0laHNV7RIXJKlyp3UbhOrzA0IbTd1OcRSJ2+75AW1yVGe5QSsjYNM
QNy0cz9JJM6UrG7Be54an7GvFSv8+uiv4nZDzS2uMwUoGwZ1VHpOyTgy6GK+I/YCH+q8QVMas1OY
ZF5gp9hQjmgQGfyS9EiWon2mwIC3+3rJlm4aDy51KpE+JgOABoeVjGDlUAk1gzWH01ATa6bmPA8c
byk6mzwIgj1wqlexJIg3bEjIhECm8ZYInNrkpkgcrFok7WV3c2/rPN1Y7OWAIAOlaAEonB9IQmY1
lLMEO5VMfW97tnucktR2BQ6Cu08fjYdz9jzMv0bEb3VDugAp2KCrbEuUzX5NF6ON1PF5MXCZ3NOk
pwCasFNgQC2eQ+J+f1dWhYj6CwDeoOVkvFGoYEI1WPV8Gtch4wa3CopXl8ffaWSwdA0Lhu9mxxz5
LZXSBIQcMUjqCbe1/N8stZticT67/ArYhzdqSzjn5ofC1U0fuEakAU45aYOirRlSDN02R6+qfUQr
VjUJay/TNcpfsksIrislcVyH+1JvhXRXFv4FtKBCa8zxFHenVY+CvG6yOJRJ6Zpq2By7muL7G3f6
rK0GzX7QXXVNEaFqDjpoecV9ogSNHY69VmHwKx5/3gyypIZ9jBXECuUG7NZbBUoTvbUs/VgV/fCH
0DDt7CoK0jxu33mpkTvlNWabdoK4c8USdS/fbI1NTpuKYCwYTPUnwtEbFaBId21lJ0679yXo5I6D
cgzVVxeYXkuCIiQZ2OGiVLcl9h9ev3EzVUNvUvEjX4FQX9lKn34oDeV1gWQj5VmMdxTC7k05H/CU
y30H4PzpZ7qXzEjfsXzg2V8F33AT48fJxdaOu9NBHvAPPTzs44VaKT0FqnywosJUVpWqWj1i2rnQ
vk9o+/ofVSjU/hx9BtIANQetz0ODostUgZscEYpFBpLvcbV/B/TXZ+HhVbkK+IYNsP8wDQGg1dm0
dhs7Nmx3zP59qUcal24LrAaAkkNqg8U45jv+k+HiYiBLCiwdrUHNskFdhLsqW3q0nAKa4ZorvPcZ
XI6dH3vs0Hv4pyRlE2L2UqGjQFxRAectJwZMjXQABxtDoLWv3ngEZzmWYp5VsoKx/L1V+Ug4JtvI
0eVwrJlsCUYqnzzguPUacEOTUWFeKdVgsU9r8yArgN+9R3ksSGQYalIub607tYCZ4XzWgAeI0sB/
ZPOPAXeL2vb9deD4DeaQdpIwIrbc55cvCLK9LXosLiWP3pzvxPw4sggdV7YW2Ay7HfjGq+pTv3WO
r+0L2quz5HztDvNlXb8saeVzxjVdvneYD8WQcu3w+e4nKHEGLe+2rn0rOkRZLj7K6M13PtF6m3me
GrfF8914VdAiaT4/hw+erWNce3+FjEj2EWFIyVmeokSESg7YERIgHfyxEo0f0PzmzsMcGiw74OLz
CfJ15z/34tAGT15Pq5dhiEf8JJsBdHD47f9RQ7jbgOmEG6eI8Zk+LzHhfAd1vB/v2L/ocTabyAl5
vydLiMF45LFqbwtODGNhKRDGl81Gx5QnWxAOQBz/3BQIL31H/P3n5OUE3N7k7BZTpzePFrj7yz17
ITC+LUc5frR1Rjk/c/yqj1fFsE1sl9RI5WJELUqLOYKmuqEyUYefZuuu+ROmQXzKcxL+YXh7K2I+
i5RuLHTG7CXmrNZIrjmJj8ZcclvqeLl5wiH4TSi3YBTwOz5X7W7jLwmiwmgM1K85z09MicBXvUlk
nRrvRCED3Fs4fwFi5yYARQjP5BNC0nFZfW3ekuOnoMw9muIEbssFa46mMpAGZA1ZzQ3+/MOiuQfH
qnjWIZmfD3ojFYqHm9z3HYWFJ3eLLj2yOLf2wWctIbkHiWbde8u0PW9QXzbCWsVTM7YmONgwr6bm
/tp8KaQUyZMG3K/t0dM95yQp7Om1ji7iMSzHGekX+fjSxi8bbSONrBR3GmjOIgzA11ceb5l7/iRP
oBwmFYhAp2xNoujMVBAfAaQhLYX7BIKDzNNN5Y5pqWTlLPliknb893+xcvF8CS1jLOcTE8g16wKD
6pRLBZlOMH4oPkfKau5y7g1j9hxfdbZpWbc5MqEkJdWiFCTsMxB+1aPk9pCrZVgIl42YKef7Lzyf
kpH8VzK6fY3JO2WIIcMEF3PDtwsybt4hAEFuOQv+GxSFZnqGVsIpmtHvaH22b9YK0EqVTtwiEaAA
hfw2DAbbPAce/SlaNrc5iVlxbJNpizrXUDEBeDrOWOhTC+lD5ZkhRXpai7RPQFMZOFWTDw/9zcEb
Ed//KBD0VG3W1uaJQpVzn6eSgDGtbmei6Xl835NIzLz6wYCQpRg6TaVJlKY51WsY5D9WUHNcsFvV
JunDfW8/M+2B/t0c3lKBTUuRbaFBo9s7KLfrJ68y0ZpoO6yjP7oefb8CoeJufHNStZkwhzKsWAF6
9mXbyBtvVm9R9Rks9u6FTeHPQBPwxjvGlU2JYR0e9ut0ZIske2UGGHRzibCGwehXL1v5klyOmfQH
8s2QQX0Jmzzbi3IsWOpl/wvWPS+oJuXuoLZAPSt4OIeq0PSjJ8vNoTFcHclAaBp2zHOFh/vPblx7
zx8QoRPLpUgBh8XVIzPdA+0topyhD6lt/0kNMVCL8GfCyOxASwpScNRPfeoF2quBJVMnJlba3kFJ
0q/9hyw2EKZ/UGJmuuImEbcJZfONcEJUX3o3IKSvrR+j6X+Owyg28VnU89yx4XrJGPCgU+JYXPrM
7MBu8oqaVn/1/mOYd+rGAh0sXTLvSd5V07680lcGu1uF6TwYQBwWmn90ejJ/X4KBok8oWx5YFHQE
QSZzYjMq6sjO5L+oCMrLhfOewtOcPYwD2VcMTk0ekbtYNd/LYz/gHQwon1hj39xuswAnqkzDMdMu
75J64ytDZHLDbGpYg7jg3dFBcjFG/qkdVqk+pTzxK3yN1PYm73EN0xALEHRiF/9aEP2sC86TIeMU
OQFmVd0cpnnsODfX7s5qnjCBaEfBQvEIDBjdNpcBGJc0uiDhUXYdfqBkqhONfNOoVbunQ6MD+HGJ
2VVW6pKb20gDc3l5BXXnAm7A5+P/jjStKCKzEyFDWwYYU1dX4gajXzzzaEVMxp91WZSvEYiauslT
qM93tP+3/Yuswiv2QCSVyOFexW8Lhb+VH9bMIreC/hM6jRWVyWb3pQQNGN2vIfqkFCN7MZ8j+Xj2
/YOQn9DJxcdGYCycsWdwu+e5QiR8uX5pDDAQs3LUy+b7vkz9Ni6GvMr9up2r0uJfV7ty8sxOOZWm
yQuN0qPd1c83TXHGQHkcF1JAk1e/30rQ2yqbK8jHOvolSq8RQ8RTatKJZJkR/5bvsmlaMB2waWDV
CRmaX6CI6TAgjmV7xtPx6B6XnRvUgMFqF8U8JaFUqn/nA8oyaWWiCjCJDaROTXcIw/AzPSpjiT+f
JgufriFh702sFIFq2JzeqFozkfF2ekpH+2xil14HtndJzL/6tOThURu3GTL2dWXPhoVu+YdKqRoD
T5mtzbBlENl7kkR9JTlqNmOkghEqC6hLwS6BFLNxwL847KfuLtG4/JFY37cvqyt6Gj5PBZ7HNyeG
Rq+zzaPIgvN0pJINXvbnpwm5kfjQGuKJltPX2HTGqx2UacaaWQPWVAjzJEFJpuux3d6g5X2yzO9T
uW8aDOLj5cCt+kyG3XR41G9t7F9sNNIrcYwwL9pt+xpbe4YGmrw3jl1QtMPSbhwRUeNZ+qBOtJEe
XHWntnw06IzOMPAABUMi4YnsTngTxNOeRLReJ+FvWLoXyFLqORgOjUHicYp7R/QRpM4HWt/Rs5g8
dKXto/02I4qq0EINK9uyHWHWrM1vuPbfeIQRRpGtkLS+3MVLKQL7PGdWZUFcMzhbl24pM7br6opv
66XSaGrnr49bU2fPQhPhmoYc+ByjaA4qhvSeuhmxkxtptW+DiIggXg0C5TkcW3QA4+uTi3HfRfrz
Zt0JE5p53qMJimxpX4TmkL2TwyA//2VnOXd2d5i19Nw0ig1JUWOMDVxQEPNUyWPOh8MEKwDlnDs3
WAmU+ErHbbI2YoYsngWlOpLfr4aG4R6ZlmvR5HY/d063+F1iwG7ifDXoUr8NVG0mMM2Dn1WhY8n7
jEe5CBovSSE8GYV8Psh/ui+mTgqCkr3ZWsxm2/RBJMYFc7DloFLyJVTARbVwnd8tMgHePTzHptZ2
gsyKtAeUzOaYJqIf5QbG6lvxB65C9AkWvKCuIPmJR0EcGkc6xcxOxc4KLy8F5tTPX41v1HGKoY+5
GDygDSAY+LUYOvJkjNI2d7NpTjkMYu2XMJoIKQVsMKC5zRRUtzcsp4dDVVET3ud2TJJj5e67SZOg
QCGCYIcLqZxe04B3Dm4Ml+kmvnb369doWAtFxB+wOcQI4xWaOPLxLPFfDme+97X//+ToTJe0EUZ5
+X/2ihHT340TLoFqQjCR1rM1yWjzeI4tsJuTla3tve1wUB8Sx1mhiM/PLEDjxpEGnMPOtFz2lYHR
rVmqI8w3pZ8wWBwbDuz0X2RrZcHE2nvDM4ctvq/Jl7D7L6OBPliRZQhsYuo7WSRbWGGickGc7Il1
hmau1y9rAiiQwtKG/gCs434dkV0Ecl0eOly9PBWefvEZyftllC0T8kdwpf08O9rW+psxWmev5Qg1
uySGFU4xWCVXzutcFCtOWXZjJiCaXPEJDt9MPTddO9QlBQTjKLE9zR8eEPf2CJNycLuyST2Cg6CK
jKEQLkjbQdVYnPBoq/CUwAq6a4OwZv9yCQld61pWS9HR/w6S01+aK3VBwqVOEfl3shdThpJEhrid
sx309aaG/W1Za+pve031wIulgDQ8Ir5SE3gzcFSKlYZNPUyh60bKtqyE0N2NRwYfeju+uO2Vg24c
pvGFpMALkh0exhdbZqcTvRmuz4OKOXuNDbHAyTLYnW8fEPgQJYNIJYDroqzzxW8HZ2Gtmb97ty51
H3+W/yQATM0LdfZxMYNklJznv7pu77DRcAnfKo3s2I2q0qamdZcKExoy1QpgDclWwzYYf67njtdW
NaqRRkt9Am1/R8YniVZ8COPJVvWvyR66SpMBWeEMwrdtgkRd6lHtGuF0LW4IE5B0gl/tTaIOFfW3
fu/lrNQJm+8PzELqW9KvwoCnhs7UxS5HZI+0c1ebAqQtOxloE199yTAtcuPGjFyU2hlDJ6APr6Ja
RiWWXA4dIAfhFbKWzETQl87UvS3tY5UhH/qQSPkKPZ8DPhrDcQ4bO8+3XAHx0NhpkeimwRjMj+Dr
wvUBV9dgVkRqP4Qm1k9ueS4eyx7Cqrb61bJJKHi9tjLHth42nA+ge+gOMHRQ32YjhvDTaJDLBsIo
VOwRo569y2SIks/7uP/k7LiOFrnbWJ0INFMG+A3IkiDR9w46/pjTCkBtCx7ToGRKu1eN23bLmT/Q
VjTYeRAATOxkTAnwZzdEysL0+dPBS+GhFiyhCZTz1XIDMavMlUvo1nJPZr5KWjz71IkdyZ4QZ9C/
F+ZfDLjMZCVaR2bBxPE8p22D0xxsLqQEstNhx+RllIrBwSd3uUvmCwp+dzQkJOvbO3BJOs9edMeG
vMxrHRX3nKdD5QFkg4QrwvatEL5PZdwvgJ2OZh6OZhOLQ4KzmoV3BTLpSBeyeJVU/sySVVWsdW5W
z902bSoVcnuBRObcG0+koEo/aNtkmrK3V/oYq4lLZHc26kiG/wAmKEHhUbHuWA4qbDYueFmkiniE
pZhV6z9tYYBpZPvIQi30i5+h3RT97ulgdawnqqaVNXgyeUKbGuedqmvAWi84JEpGRwAWaTT4uRnb
v88mZ+A/z3UKkxE8GiazzvXgghRQzion9p9XE1WsmoCKwNENzgkVcJIbWJnDPxTIL3saYbNbTMNQ
kuDHMFGvXmwkuNgCpqQ60SRjbVSiBksAr7dPssKoZ1wDcvGosLZ0c0C9iZNBMi+uao4EIatLfPX9
+hgtYBapKU3Ucg4DolijJOlZYY6l0VRBMRYHGtaToMf7mzQ0kqJWhuaizx6iqESxs//X0aRkYUkg
bepNPjW0UbJ6HFrcL6s6abvBnIzmU1bMyeOwIDTrTlRIxmE1J+QKh36pM3bd8wDapqQO58F47rLW
I3guc8FL8DPSM37GCpN/W2UvIOSUFDuuZc/i/aolyJ5kageEQSXGjVnZeXicG6a8FShdpatE9RbW
fnRbj6q+aZTsWzQ67Y5ayDXkYGwizN3EvERQydEIPwhcgSWopCbSK4dGtgeU5O4Suj0kVJaAMqIN
HjMWTzDMwT5mfOdEsQy2jpGwlMZOnRHPnvzDPVa6lzbj2Tu2z9Zt6oKl0dKFFtCdL7eFfOxzih2Z
Y1Vtqa62TTcN/SyUVNwS1ujU2tEBgKCoTsvSzZfNPwfbm/iSv50So9UQ5st5GIwxW6mn5m4Ovm94
50rsSRHXTruh9VUYsBikpLo9Ms8pxNWyk2Vna4fsduigr2MEm2lRlcbEyLUkdZO+HSbGiHdnt0bo
2fy+gLSysKVR7Re46+LHi9u3BCcUAsvhyeDoyXA132mIjF/CoEGgfj1DvSly79JbmbsyilWRFnXv
h8W1gjGiCpRMVYnaMca0V7b7UROOTvzrFWo4jAuhcwBFTRATKQ+SzW/jdhgsmzewu6rCXJNFekL6
dl76LPStcDFr8AN23yJDShpWxzvGHiCDTANpn/t4QqjSrcxUKKQ6LLVlf1yopToNKduvn4w1XhWC
Y7zpNuXwomusdZI9eM0FmOY/JhKXnAvIdkScorfFIFIjQPKw76JS8hGj9F/4TmA/HGJg/3JnWuhP
ejmjvhZu+/DtizOiko84Zz7H5fLc/YFEbMvZUwL3Wxvj1N70bgA6uP7TrtZW43kjkBYgs3ku4S4f
VZM8MFrvNsL0kEOxzDo3DbgCjXsfWuP4sXsXAVtZ/bu69uEkF0Y+G7Jmy7WXsdBa6mLoMVa/qanh
T49G50f9YjIkllFfin+VSRkldcu7RyOcNe7sS2EVN3dfnXru/hCsUyZQACupkS7o45LQ/O16RkMi
NTI1DvMDOkSaEMqckA4XG0S1DqZSKidA1AUu15eYpquqQ6MTnrl3X2hOzB/aYaVrruvtFcSG1QN8
PE1AbhPk2r1Tk7NbZ/CGyiLAyod+pa6ypkjaqa2Gkru0vrof/iEm9HCZSPM7wOCrh95dHEPK2p5u
QrZtTfErmhPbclsdz4SuuJeBa1rdYSpw3Ct0Tw1tuolKn3PQyebxUSHB3qhlZzGNSYkTUTIjIpyp
hPzp72xmZ4UZ/TFu5RqL5BcmWqmXMFvyFTbMXZQz6Gr9rqjGQGMuuGsvTIUGXAKOuL6d3/XNCwtL
DmXLjGPpVjELdtJdFVaP+RbCnYrvmdevmQ3Izm+rGHvYPZyJsXehXdmv77Oc4S0lELeKKBEzzHSm
46OKbTvqoyw7F1IJv44+otcp3CdbsEkD68264vPyKXQrVjzoqZmORnba+sFrAmlx8Wx+sc2ktTRo
GDe8In+BamXalphobbMJJ0W2Le0CrFLEXkDEjatknUa4z12ErNFSOjZJL3kJu7W3TYySlxZNUsJ2
wWCkQslOnBJHfxTqzfuDjxVYL4jq4kQXmph0i2sf2Nw57aCdfoV7KKGjFKuHMka48wqIQh8PzXGY
Mu54v6JwimkwYGTc3aMEc91gbUwPqsxYm9wn+N4BYtO3kKxOLmWtlgnoC5QmAQXdwsOfFLzhU5Mm
2ftNOYdt6vkSoTY1FdUDNRbc1EsA0ln6C7PitmBJ6FOKN/n8EX/5iTL3K+TsCkGqcuy/oH3aIwOF
GYIMo1LTIlNdNhGjWF2jAsXjVOIXqb2mVM7EpnTKClaSz9CHOJZiubnapHVbsp2J7P8e58aXCrGI
6DI0H46n/CXo7SW1trME2Mx76NqKLFtPAvwAUA3Fnwv2Pfc5XWoFGFUvwVuZr2+4zoOQmLwFikpP
eDd0kmr+2SiulLAFpEKwXrZ6bOXJq4fJRjmBxGDBHNRMRRQ5L/jl7sMDlGrO0G/qP0onrdAeyySA
/CcWGd/k6FZZLVHgJVkXT1TzogcQhEzXJRftIGzTKhM8pVZxpfVm5HnER/a98Am3osGY+GhftvBT
5D1s206S9MDpQRcevTVIRAZRRHTzzB5DCAnS3NvnOSz0aD6gZMJMlou0oW7fStRYrzVGXwYgYhb0
Z/SzL4veIo6APHuEdLkLZq/l69BNXlDGLPVMyp4XN31GxofbLKokXBrsNk/kjfhLQFr8Qj5ZCF6N
+RxuUZvoKaqdzk86D5IrPJEMzpyeJdXmMYmfBtOLbVJgrHeo4JuP6PutK4SYajCd0PsbakX/sBgT
Cpx8gbtKvqA6aBAh90rPdm491r4ZOPv9OaQooqlJNx0IR7uRuxLIRmjEE661swKdqfkkmfIPc3N1
heHjDjtYt3Wx3kq33PtprEtguHoC6Ad1cXcxpvcL/Pr8xgaJTb1tIRk+e1eWl6/kPkPZXJcluC0k
2yR2Jf1ks7J4XilghHC6v7Td+/KHDp/82bs7Ye6/Zn9qoj4iDivveC0gNiOPeql5v822onumWNZS
VLrOn2GNI44ATSDTYTJTzD6lspMtAG97Ki3nF34gTFKjnWvhuQ/RJoWrfgxAmSF05FCfC54YETMl
UfZkCBmiPZZaa3+vFjtvOpzcYgxQhVU39AAxf7G+y9dCUYciKoiQs9jHtjrjVhpcyA4q9X2iGj2P
6rIG0zGnA2G+1WWN0pjhBp1+ThnJDB9cSkc9wFVlX7tll8YTRcDisAs/+QgWU/82nG/4XBLSMuT6
3s7YZy6iXHjrMKgShiH1HwkKVfFbHII625l9FJ4rzJQQshYf3wkW2s9Wvat/oiK7nYw+q8ch8wHK
HQAgzrWfDF4kGDr7swuXj9jfAwcvI6uVDkl5qxwp5OXdr2T4XrHIPXpckRCFkaRfwsidwgqEQjBM
6InNOItiQd7KXmTjXdEhkWjvCLd/MDufIwsKe1aLggP11DqlCWAqXJMZMMUQxggLeYwyItxdcKlk
bkVbnZB3Z2wp8jUJ0iPuVuU5zwvbXQ6ZoADU0nUZ2Cng2ZLhOv8hR+16VRpyn9VgbxQgdJngADdK
pFjVydcxOa6b9w0wYYJgI+B3LI7Fr3/04VBk3jSbf3rAXekzj02v7i5TSbnoF8MIVa/Gjehm5bUe
+/wl+u62TVxxPNnh45ezvqSVH6I6/4Ljwa2aRQyy3gebd2iNmbOLkrJxdA61yNTMwOfXiPhpwY+Z
AGDFMqxUdVpxsyoC+h5tOYrv8pnGE5HSE4nYsrpgMVyDMj2VUQjPVUY++HIZwY+ufe/KaDjiYvSY
B2E8p62aqBc3kC5Fl4yFl+N2Zrtliam74gnBkUjCyceFyan04xrMNogEiLQypKjdQWbAAeyxzq6l
q6107b9S7CIfKsxknvRpuiOt/evH/t3rZ+LiEoUbkNaqhlXjdOToCpN7cYGh1NOa4mwB8dSN1YgP
pLVB41bh6p94v2S1E6Yovr2xnrdNxhW5HAgWuMjEJf9oCpCpfZz7Ab+9zS38CyW9AuThdtGNvEa1
usi5yD4uXmEXzbUiB3/gxFf7dYjS/vMIYn4oBwSrTNwe4iK2U1YH9oxQGiUDCFIuKEBeieKh152y
Cbz3Rcx5Hb7eOIzgzzc2cynEbbItZYyiW/PWTl0aF/3maGSiQxuLav7OLy1dBLeW2TOZpY89slcQ
cj8fQasHz9/s697jeh+SStdL/MfhJubURLBAp2go8e9dmnvHSBOO2oQIruugbiKnoLDNWA5pC2SV
1Qta3E18Jf6iUvBNRbuuU5aTGByTjXVFkQOkXQE/020anp92hXtg3YYESQ5lyWcHIHfjTOcPQwkx
04pnKvIeZjxPiPAGaA+Xr6q6ze+Xe9BB/ghSnhnCp/OAKk7zPkSFPFyhh6rNYtCxun6ynCqq1AmL
bmLF/D62Wki+UZgD91sByZE7ZM9E+gkZYnBnIhjarfClHTrK9goHu1lB9dmcXAoYYynSRHth+vVR
HVtyIaA1woGGIDZrZXxJhvpP75zbM5AP3E0tK+OqvcJel6lfRhUNIS7lqT+uKtlVXmktdPBx3hQD
ySOh25oo0QJ9p7d0FKiNH1hhmuhwGm7T//60ZTJmkD1ot9m9plYXOxnp/ghvM6WiacAFG0yqR8dV
4v2pHM3r/GjSSiL7zAqxZwMQydAYy7J/d7B/Im/5mcP1BXhSaEEPN0CfpJN36JAOKPoWMQTT1ZVB
4HLhEhuCBnlGu0Xot3UMEL3z6q04UnMKsH5poc5EW54Zgjw26RE4WeVN3VwQydUo3beIyGr0S+2V
dDH9lv27rSOGBqFSHUXjwgYsFE9TYQ/Z81enyKHD6cCRe/Wb9kjXiZGMfgpQkB7cq2pCf2fRjfTK
4MKPXvHhBHKjWrHFOw/jGbkEtV/AinMB4dtnZADU8ew6ryREpmOgA5mJ8R4zSVhHq9JNgSlHVF3D
uCQ6tZ4C28YT0e8lIUnXkhfVePFATsNlNX88TZXT62LGuTDWcaZVld12pNN+vgaxmHY2pt8/vAsS
oE/3l+FQoIwvZs6KCIwsvLdMqWr9CElruniIevFyO0rclOsnEU8oGmTi/bCkmESA4+ZusCJPDirM
AjMpVWCv/1DnWLdez8MLykT0sBdVTUYCBnlwqcEMOazFBJjvrz0ol0Jaw5x6XUBsW6Cjd2Ch+sGV
Pbx7kYLxaRo+YfDoMhPJ7vrRK87uT/5pI9rkkovT2hRRR8RKNOAoxYaGwi9t/ic0uAY5i76duCaz
vN8JDWv7LH9GKLKU5StB7JTNjByMeLWZGdQuL8TKVBHM/xNLNdF9hxjYovaTkAdB0j65hKomESQZ
/ZuOeFgvk8h6+irD2ys1WTJApKZjj8eeCobLi0u6sjk0AWO/VFV7VqPYjR0v+4RoZ+V6MBDtJp+X
hKFK0sVpB4GWYQT7AkoiHHRMRphrmnrTn4K12N62CTA03N2aX5wN1tCxvRc72SKG4beFqbhXrORX
rkja6l5v6AjEcnSXtn16rWbFrllAjvLdFTXaGkaKZvdNtyq4zQc7n9SnVvp/5xCzHNajoJGVQhMN
Blom+P5ApCMauzz0Ob1b00ckEjZ347OU1NcRKCdtLLNInvrqw1i2hWIClPhfxZO+uABC7fBhrAoG
Vrh/Ymc1tcdzQcTF/KuNLwbmc2fN1M5v6C0QksUtWeKiCH35i8Z2O94uQLOg0hwa7+gizucBimS9
D6oV9oJzSE7/N7PbypPEyx6O+QGmRE0zlcacjGnW7VwjTNaxF9Hrw90CoQg6FxDT6qPvFNk5ot/P
VPvUmwM2VmmgfRPukkTcxZvJF5Rz6Iv+AqJaTShNs0KCpkU5JsJBUwWrXYJs2QPga/YPPvtFfjmX
HkrLIcNeMfXoqjPK242388r72iYsRPkFlM5LbCnP9yTC/lF9+99X1jyNHANiP69k2DnODQWRh4GP
w5Yfp48c/vhxE57OLanyWXxyhug3YyOjmO2q9HXQqICSFbI3e1De9E9vvSnoZ73T+k1dodAIHWW5
C+a9SLYvqLaxLFbJc8puRCERmBNWdy89qzBEGt+X/JMQYpvAGQ8zpos9ikOSRfXgWgHBc6+Qg/Mi
NMjFXoPcFAdafQ648GSm7YFiWI0F0sCqsw3GS4B/I1vHXnTY/TwPVunlqwQuRDk+q8VNZ/S8y2lO
l0rucXRdCe9LMynQFa+csweNVYmII3nHJC7rTM33TTZEj4Xj+nKFv73J66DeANUkdNd72mL8hh3+
Bii23Y1xkIiUfp8OrOQ6oaNxZgJlV76+l4Sz7p/JvCTvhiiWF3pd33F04SUJvxptXOzmLWDT6fnv
fVtsU+vd2Dotr06QxCh/9fQW3azovQ1CLZ/Z6TSq7OEpQb2+UkOhKL94woghCCy0Kf3l4ucOUjmf
PbkXqr5y4bFu6sWafaC+I/E4WuItJvHiaDxggdhYA2TLdi1pZen+VOUHWS95I7W1q5MFJ6G7ApUE
f6cN2q+bW2j7AIuh/Q7KLRqio0+mQqihY33cU7mslwA9ePHxGYgReV1ai3M47uTDFe0S1VSnUhU2
oO7hwtP9QL6ugw0FWBJgBggmOypc7za0HdQtq425sDF6F8quRItsn9Ur0gpGG0NFkvymyidEJdZm
WJyvzMPKYCN5pFbX8ian7DQ40nz4Jxr86Bo9XOO4x6mtZH/Nrjf2dN7tCZOnzjuBZ6smE3ImqvvD
Bt3Wdj1iFd6SbVUD2Am4XRo3zI/3D1md5raZB+WqgqxjWX+qYAFbLAXF/kyDrQ86bXG6UXfirUCe
b3eCC2CSXHyorpqD39Lthl1zT0FXzgEL1MHo2x2YTcRcJC4d5/+qBg4P5+iu+krQGzFBq70iOgH5
69cTFrYdixvEWojCmUBHWvqV0wLxgLEId2+GRGW3mjwmpfaVplyXVmkiSImbipVnlB7u3z6SRJoK
8gdQv/jqZQFiRYS/SNnX3Bc6WyKM39CgSv2hx5mgNXgAK+koxQa0wcEXjOat7YpFH5dxdfoFQwrP
agWwfjzsEPhrZrci3bLC6qBK0i9IB2mwy81HgSFNZDeyr8KcTpeIUJWnz/K0WsG5jCIKeIKmYdbf
0oKTJmnxc8YNlMpOLTDCB4thrinzvD0I3YU6n8iew9ymNOuLYI4B5SWP5u9l9l/8D3XXg/5Tv/te
WHQ8H7Tfq8GbG95IDuG3V0mfk4mumC3fA1Sgh2plxJvIqbKHvIrqaarPXn8S5g8Vvr2DIWsdoTUl
nFUD3ugVVGUzGi45hTpULLFeGEmtxsIxqdMHhVpw4Q1WqmMm+Ot3EO+/q8xPn6AuDeeMl44KPH/v
fzzLr3+cv+PQ+uDX2m54I4BNjRHuGxYWHqzjkSUYnw6bMLecINm0rk3jnHWXRSnfGNK04GWky5bH
yAeL19NCtDD/gzBab17twIi3shKPdILjDQylYxNBh2ElU8iWhnwWEzpm+LLjMb+qBSXzxFZk4Yof
q6lf48iRLUker+NADaXlezoK2sWhVUh8K150gGUya1HiEKP85DXMBlH/k/2Z14gQRePScpkAeRdk
bb3OKjC2IVSfR77Ryxzqofn+55vLSIO8u6VCtsISB1OAgz9KqkCEiChy4LkvPdB+0X83YQ65s37T
p7IG8S1fEvciWej6YoV4E/KfAb/Qkk1ozOj40mrhvuDv2CRmZ6CammfB5ub5qPRpd+B8dfog7Fn4
aduQhF4foJAuyLurA7XI/fczYHxiDrKi0jEFYFyYlMxV1absnnjbbt0eYOWEwkIGuWaiYXL9xRf9
b/LcCyqapY+NrZ29z3EHoPsGX8CaRj/8fq3rF7cFOFnu0NyYD8NtEilpqcEBhV+ZvV25uGdlbWsl
8t1YU48uFH9tceycYWTxgLtBIZTkUkWDFE/i0jBOIvEa/2QKL0OYEvavD0HxgajDJpm7Arqk9RgH
0Z1F9RfFMMLUAc3+6Jr1dCn1iznVaLy73KNWyaKsmtGggc/fMtbGZwuY4Z1+2lBX9FEKXj0m+6v2
xIFY7Uhb2WlLdajFsQhMuvgu7YSQHjyQbFmcf0M2HISXjltq8CMTXxSSunqBjCwQmUR+5vn2GIdw
Rf1Zp06MmgWuslRQEFR2Ump35zLctHdu+bvlaEIdF+egf9J0tnbxBgFBTxlQ9jD++QZH7332jEDd
QvstJn7nveRGLKtt+C+hWDNVPdBFH3fwhHo1BJsn3Q74zfB62Qf1ndWbECjeg9G2/UBcuvH2rNuE
JxI1vTXel0yWUrwXsQ5tmuj599h9yBxzvmbBUmrjK3zbcsq12sSl8Y0678FkFUeRlNQaL2h/SYtA
hKkr+8576ITnAtJlu7veltrywpehAeD7Hf6Eq6CV5KOUwBfxeuWNzY5pZzsQHgw5r/dkIfRNrNXy
usc8eykdY2PP2mgrGxbwTOwQsB2pSLk/lgavmwHQhbBw4rah+2QrFKYnLSXnUstJgBEUjzWFtjGb
IXM3obLztgvvw919ETsf7yO8qyZRaIsjZoMZ3HPJoKYAeaKkf742D/DGBGZ13FheEekNheN/upsx
YhRwwhP3OdusGwYsoQkAwkz4y4AqHHX98IHh8auzmtMBQOlmcBbqtyQMrHKuzgPi+JBLa0zOLf5R
vO1f7Q6xaPNdTgzfPlDAaWidLW/BRYB93CWJbgCRq+KGEoyh90+iwLIqjjrmubA0IHJ1QY4CSaJH
6Rcdt1TZfFOnKdtIFivdkpyQZd+UQA7wij+XQV/AFCB4E4TayEe9SKOwaocV+fHaxgCPBNndTBEL
hkiK/w6gPzEF5vYLxVYOC7RJb8+npX6ZlsvHdwzZ0FgL5faKAPNY8Zaxohe84pidA/G7I0jn0Tpv
z7FWmqeeTJbJEQjpD+eYaY5FwKrGesTBWYtsow4H3RdvG/r2KsVJpCO1ts6lTDCS/6Ed9ivPYwq0
5Px95lZCa3sZlQ5YWKCCsDhq/ZV3DszMRNEp4qFjqfv62lR/Gdj7F5FXxht7C0oxZ14h7/YntetV
NxpTcO0U0WnHDo+Gmf/f7KS+0gZP+qCwUqaV7+7vAHTaZO3axVh3ZLgzM7DMsL/OzbTu1u0hx9OD
oXlOx1KHQ8ByRjE2eQF1ODkChbhNhujsILuqr744EftDxcOzenYpIzJ/tlcSV1b7H7u9jA1nnwnZ
96F0KC59LnjGHw1s0jspgiUyqkPDgYt0kuXZfyS6Gn5bwrHhkxjv/pW3XNgFkTFBCqHxyLkEJwT4
PlwedZAsUg+Ud1Do1xsk2hTEjxSALnpsIsslDN9QcFknU1+tgQWhTzmkwP1gFWO2FZniV45eSNcw
dseRSq9lqEIiIKlds0wHl/QyBpw36I5jaJ7gD+9E8OijeGu6Nx52y0Btg60dasA4dFrNhGbkiY0P
oXciObJV/cQmesSHycwCUuagBCrjNIdtUizOsXbzQbLsUHTJqxZL6UWmkMLZfNPeRUXz0KcuIJYn
69BzCUGibChAV7hik/eylD8RIRJ0kX3Ij+NaXoXcLOtmBcsgQCpjXIbDrV1QgZ8pcGRgKjF04okt
SEvKmUKpvWQjzAc00n7V8RyhGM7vQvIs76bD6wRLCR6Yl3HZzR2Hp1Xav0ALBK3bv8eizuyWB9C2
wMJjDZd4L3yOrSbawUfYA9uBwRvOLFCkCu7MWuOowiTLaG96sbwhqQHH7npJm7Nwecdwil1ZPWlz
H5vnXxH6X0nFWseoPmvthx3qEikbOFzGb4yDjmB0AL1rd7jUI8h0QkCu/2XkaUYMn9HV81RrITGm
YTYqm6saEiWdFeVQ22TyNtceGl3X2yjnshgncYw0Zzx6kZglOyyESiNw28+jNrRruhbda0vqZ8/w
LOtynJyeJTtWFBJ9d7fJ/ZYIhqO2qoKO7cjW6psyCpVwz/9I33KfcwUwkMxxyJ2CmqLFILvPt6SW
9hgVw7fGhOvmjnDBCPaGwkMBj3T0s93pF6/7biQaiOTAt/LZ1etf+1rqgreOzYQwtlETo6eszfRe
x0nNrkpwa2qAp6yEUsyIr+S28ud53JU5itSTVNo/SR0R6dnJyWEBHiOszk4RaKkjZFlzRDMCcMLZ
6XrE8nVJ5bR/ESMCTlGzIk6cxBp65IzQSp1IKSTnUF7d6XBmJUCuwskKZ1I4bK/mGX2jVCA3Wg+B
SM8RGVtkTQ40jCw3+dvkArYkc6FFH4wr0VrdoxnnAjXwPDkNYx1buLCjn01dO13uG2hJgj/ZXZyo
YF+Wrb662fnc4cwgJ9mr3Z5q+n39yF9vxixtr6VqK8kwulA35vfyRJKHlPiG2UUsRCzPkmHNfeku
XSt8v8uT7bdKoWlQ4bVJ6QVcMhcSyF/z2w1xYQB2Uv0R0l6dFp8XCZe1M8HoBzVgxOvf3pLBJkQW
mynCYxqcvFZ/Og1Y1M7n4QRNI4ZFS6oRLLZrOFefbLGWkqSrhig9X4RqHqWXikVva8hhpzKBBQKD
WBWnmmDPr3axu2q6zPjvg/pKkzUvh/n4toU0xzT6+CPWfWfyQIJWruzoJTz44QsQNYjMMV5XmXgQ
QYzkMBw8xdpBBuWYS3iEen+iX4TXFuUfsJosYumgZMl6aysyD6jcG2UgPjn5lfYy4gTmE6RbhaMB
sRCwy+HfqlHcxwhDNzgUmIXZYok/KGUJ03kd4dzvJuocmY3LhYdRE+o4M49/LQ82x2GsbPf7/83J
wzMaNNmoQc5ej+Kr5FJoXWz6PI4UCA5JLaut8SAv9JXVhboQ2fLfjUAh4M6KEwxh3D0xJl4k2MZ6
RqP0MRSdk4DO/EDfpmJWawhjaEN1km4Kxv4I0bFTCbq6FPGoLYZD8ogh3IzizbZi/nKwGA2Hgzyc
boS13qFYFYy5fmJDdxScvN12Uu4JDtzklEM0bab2+foFa91wwlyTC+dpEWqkGw2sMlVqs6Q9c6eH
hj3TqEAsRsynpHYnyxn9YYGN1cODzax8o+GveiIIKNK2uPkqnEaPHbTdmCT3DQcgZevr3FstAgXm
plZtkZvFQtdHK63UjOIKIR9S9zaLJ7JqpXQBHbZpA1biDavX3GETyWXXUqRfrwgArB8PIlpghQQS
hUFpXM8FeXGnuHFu9h2lDuQEDhU6VyxxXGfTP4vwALPYffzXC6mdM3UaQRPrwmQz1VM3tIgC4rDY
6/5rE8y1SI/I2DkEajgIo93qIbAEt8GtL2rbNy/68VTUdhuKmyE+eP/JNm9gObUkgdMlTkGx/AiP
AgYRF38tkRvyJIjYLQxvkE8IY91r8+LPsycBXXUrcpzp1FUkk8s9RIxewbO8NZ2psq1Tv9WqerfM
3DLCZOh4Io+3ck7fADSlTMtIn/3me5GnHq3KtLhSVP+mxuN+vkwuaszzJIxiyf6V7hiQn65fzIjn
BPJMFOVC4klyej0Y+0ToIwKHRA5PKcLVL+fszEMR4yZ0FR034WLs3mscDdQ676AOrmYuZiDHTpMc
HRmhLDxAY9GKMT/6n1vCu/jTWHFercElciFq2/YDrdQOfpmGz4IUuy1FJs9K525DT4hNXcDDOcCi
+aY7wFhZSMch6bJqaqc0qmU1uK7QVgoHLcN0d6kxRGcZzIEaSCjZyEdkZUXTchvHm92c6Fx9jZPQ
sw6e1qNWCpVOmf4/hflwEnKS2BeslGkDI2ht9ohky0b20UCTTnzOlP04K+6ZzWBL5WxPBOAiRd7f
GXmyWIIECoWgNCKLwCCytfutp8G92LCCxe3Vq4uvkLUF5ePPtZ4xOF6Y08FaY2q7v8EqlFQntedx
oGiiow/B8SAGnPd9qnpi4XaOM+gbH+Z9A2iwEcdw7Yd8a63HsfmMNeUHfO+DkMG0mxqG8f1U9uYw
ExCnPVSYN0vjWB2sSCml1Q3ilH3HQKUFic6ZdY3ARmUlDHc3JeHuVkxznI1almOprdTwyLj2UZsA
fMGOd7HSouD+RF57KmzoQbK+PMV70RTskzZmPte5cpgqPCi1IG44FttJCDrgmwNvbTFdwlv6n9Zl
VAJzM1CxcqyXaWBiDPXdU0b9K2ph30QSViN5uEGME733ynCP7gJuh3siFet6R4gtvLkAp+MxACYN
SAz/ePvQHNTq1vhIigQL9NFp6HjExkVOZNR2M67LpOU5aSryuNKTtQ1Pjdj09D1TjIKGOB/TXuWg
dq3iSN6uFgFcSj7SbgEwZgVTffjCDS1hPQlvegIqksSQfiG/6G5MD+YZFl6FMRUIXDMZ0AjoPXFs
D8rEMfZfMZFCvsrtpZ0yrNJG4q0fkqMg1k7x5/pswjC//9R1+FWTOLE+v/NVuDZ5VxS1CW0jPFbj
KiXwK7T/vbpkwtd+cOU4+t5QmlXdhZXB2gCqB80DEfJxpf4OIxydeqwaJ1IjdzaCg/lEZG8FVD19
OMnufE+TJniaoSG5gX4KYdf1jY84ZCr0J85HZxYPYM5GmRD30wwm/3iB4CIVvNStwQFFJBhi8N5R
vRwOxOhTr0X+5M+lr8/IL2sEXTiwObbr6kz+rygR1pZoHoe7Ifxjm3DnwuwNfPmx9D1S7SkRpsnO
0rgOuJZmhoemWQpKkY4L95ZUEOl8/hWKbr46w8nPukzJghpDQ21ufbpXCwBoaKN38m5/NIo6a1B1
7WmP1xkBHafiI3tj+zTCjocnrQSYsZPyYrllC/ANR9EJuGeTglB6UOb8jAUqqhMvS9phL5cFTxYJ
RkOvCxvmVqaYw4p/kq1OhLeYfwB8CCOCt95+bFa9L7VLlVhd+CfgBdJkNQIRcHUhTUgY9rnbHKM9
wmuG7gUFB0nqMFLtab0g5gpg3gIcDCPHMU01Mj7XHr1hslSaZ5VDaKRq2rTPbv971hVt32Gu7/FH
75Ll/ht3XaXeSYZ0MO5uFuGfK8B66pOC9xCxxl6qTmT2uBLZ0dMryzRDokkcnBJswV6xki5gqE2j
k8CpJ5sCtybwiG9XjSyhPt2klH39cfUE2ZOfn43uYzxkL8dg0HBfmDadRec2GNTak2p7feuYBPcx
q4dKKpLZQnzIJh2qePoVMCFEF27Po+Ye6Fse3Fk5C/frFi7LjKyq3+Mpix4ghbHxisKc5n11P1iH
BeCzcyVzu+bc5ihAXoZDbCQDDvfUxOSAiigTsK+kUekG+/WlNiT6mHyj/Jtr4xwGCH7ivqOV7tPq
igegobLwc9GE6dmCh3aGfKh6rZifnl5YsgPaiiJ4cTIUk2o0BHbX/X9ApsVwBeCE3CqE/EMfqb6f
T8vMIkdueodWrMKHdqp6iaN45xVuZ6Y6NcQUVsW0FQnvKDPl6bVKOPqCvCLqUO5SBdC+Dft50qJB
ijXsv+pgPRI/Z8lROeCoN9O13emNqDjaolA4SDKTBLO596IWlDvnJrM9EDx9PM8guMc5BMow0mBd
aY0k+ozdCgwGwbfn4VfNwyDnF/MNLuWlPevbpx9nlEvQDgKkGRgV2qgqPayseDacl1vPaG9fNkVt
KWKEQmBmk35379YbFjyxWz1vyVWPQTheLrT3FQayIZyvYbSuVy+rJKh8iPj7fFX605x46Nwa7+L7
DBUc3Mpo1vrsKZ1jXfXSp8MHVvqKa41YJ2iG052+mbG1SCqUmm5wSKGlKu2+FwQs3UIreIkNjdvW
ClhmeCYN6qjiKxMW5nnQD/jc5WuhPRBIhCwPw9v2Z27yaAisnqKcva6AXc6LzQZT7IlZRP1mKtXM
BmqeQ3lMyhbjUqiD5Z0XAR2r9g2P3VJw06/n9Vh+k9Iwjzz184VHN3CaWncmUoqK2pGtoU3Dmv8t
zWbr6XdMNUySZBzJjknoe6hCD/ynzYGusBEKHbRSfAZ1dAV+mk2RTApYNirEnFOYJxegtzRp9+vr
XkdO9AHm8MQRfHqROiMbltmZv+oVaiBbUCKOzlTO058nG5fcYM+LaNo3vcLI0oDB1jaHrrPB9Ipy
cufXhRFUZc0itu00bymm17ISWHfXR8/HshLfx0N58Kd2HliXj6HSONuZG2gtqAJvZxPw9MtRzSPF
lvbofG8Vvwg8ke4M+vU+Aw/CxcynxOojAHqTd7Uj2mPiYocbwAC/UwlQ7SzchD0XIjoQjH6cz9fe
nyEbasT2wIk/x3MGA3tbNQjKZ36ifyrB5wBVYEhwqRYCbEe8I+O7uGQMQ4DnBEMAvEhKAYMVknPe
JLhJSZflV5pYvnHzfZX8gpRDlqs35P+JNoGN3aZflFublX1k3d9zAAzWhOwgCrT3zklh5V9mmHfk
eLZ6MlgM5E8O6vWgBCGv0wuQCHqNpZYeWCAtmjar+LhrKhtW3lt3+n6mQ0We2BYlZBlrypDEwBzm
FBqQ/sFGPaMhR3Gx+9tTxK0WtpgrfvyjjMzE4YUzPoatZs7JGGRN1Ig5vxbNO7P9xXj4PGGmLnQ1
GxF5kGcp5CVhYqvLlsun0MFUHTGVJqBEFev7LT3NA5FAyUH7Z2VQZL/swx8mldNN7hP5o1cnRyVH
RBOmxcpjihW+9/Pn0BQEFz09W6eQE43kmW7+K3SF8O4f9RSy7QuiA2+LWfCi42O7N5VIAnKSZ8aN
f89trIbPCso+C0zspHscraR2HENvNL6gKgS+XSFAR51bB8o0+DpKP+Pm9EizjuCOU+yMuESzJ1cB
a32+xNjCx/QjNnYNXaUaOyHgEgRX3i2IbYMinhtcAb1oOUuMIJsQFSRvjA1Yr56+eX1xDgwcI3wJ
4PqrffoQlAy5vmThTaWAbgfpR3Ke3gkOqLuulqJG7Qi8F0Q4dAc/aBZkE9VZkdQPdXdjdVCt7xng
woyfZwX/osVcVvCixq3Btyw1cHSUQBDWfiM1hbpHdPxD+oKSWpDZZi0/6kEojVD97tpMVpz8gY30
RSJmYRhO63QIF5YMZ5/JuXgVft+GV2XJSsCj8YVGcQ4hUkFkCnfgwIOZPACy2JJJ2gGNM40eAtbk
j/MPv08kvY01yfFTDolAdhjF2lWa5BdbNoVDsVz01MTsqOYy4AUj0A/5xAIy35+9+0Z/1foFGsG9
PjpAiNOUUhXt08LSCWm4vQ60ZTYQwv3hAjMSARZIl8/Natv9WBNkPkkHaa61RAOprBJh44VCu1Av
pSzWJXtIN8dyDEivdq4ZBAVhzCW5b7n+wfPePyDeCSc9UAny+QkViEMuwdZWe/zpSosoauIvt79Y
PVM2aRAdeu7ntqyvv3i14/25XljmuQQcubkgyMHLbvVrZ/RW1vB1Mxm98r0zGWgxJSQmiAtBEGZO
1UcehRRbPY/7j5tHD0ma67Jd6TXB3WkPYEoMKkxL37v0pW+HY5qa1vH8to2uJ6WPdrjQliBg50/N
oB5v71NIAWvPVgoQreYc1/hHW8RCHpVXAX5SICOBoo6UJ/Y2lSgBZlUl34Liw2YSVyYfH6AXjZJ2
3EJyEsjNFHmeW5pTQTdaMg+gbFxMwN3F/l7bFZD3WPcxtvGvBJXdm/9rB6D37jkx57VCBNW4fuY/
wAURLzjV+SbU5xoF3sNEHQOJ3b7nKzgQRyAxepF35cOgwiX9kWursU1alLUlh582Y3otJ9eITwQl
/aBhFuI/EXC6DrK9Znvdj/WrnMm8PI4W7vG2kz7k89u1+qfIrwFOs3uIHvPi51+0pkeU9Qhcv27q
MajH0IfkqvM+2IgmYiIe8roFHnPCm2zstHEzr7nOMUCP4cXICJKTRqkMF419/BnBZUQI8iQe1bzd
ifze2jK22MBw+RHihtHI9YPg2L030tXjQuDOWHwTrVq2WOX2jKfZyHuIlqXo/IZ0woPtpLZ6t9eA
4GJ0XLYepQWiMOboE+oRbOPt+gXU2D+WLa7Tmq9yLFK7wT9ea0m+/NGDEDt6xqNoJ+KfMRC5jUsa
303Qrc3Ns4KzZUzx/TM0PGbucOG4IUZJVFXZq0xn7tjY6SLeUy2Iv79xoZbiQfLeeaWDD/bmH0ze
JWt6q6WWUP905N+QzMO1f+UrgnzqIuu1YlCe8S9rCPWHKcUhpC78wem/rCYkXyRu8Qho1tUxC6GK
Bq0FlG8vPyTmjy5l9d8NAxRenCWs7Zvt177bEKvcInUZ10LvARm1kZgOeFtdZtLLxNFbxQfupzuf
BN/llxFwcM0PuQ5jWdrqo1EyjY2GSl6eIDovvfICMANhwufMVYkrSThrJ2YDsaleHnmdchhZCwsz
XJ32vuLEzvrraFnq3Qs8Dc3F6coTFXDszjHsYDNKrPPH5xWECs2HlEIjWrtRpJZWRFeWShUo1vqO
5HB/wD7Q8YkvTY02f1xj5CWh5gKjn6l/5hRuKQNh0O7OMi5CkFI2Ayy2MOZu7AS1o2n+2oPRZodA
2Qqi0OmzxjTqozTVlmzJQrNEkNU3sLTYvkE7Cu8X2sQ1C6wSEqtMlVcmze++IH97cKXDa9IYK9Ol
xUVjmWyLIwRtyfDyi710/Up+N3BCM2VLTNX0uipiyu6jN7E3ULVGEqSCnjjEVN4MTLnRIRFXpehT
Ob7Bh8P2rCTbFjj4CWYL9sLw7G2DPtk3RnDp/RuJsw7M01fKWsvKR1gdaRnkFRYwoslk7rDqFyD3
RsIhjNFWPf7HU0JLthIIakt+E40z+TC6mtDw0KTlbiNUgRgnZ7mRT0tnjSrbJS+9BfX8v/p5IA29
KJDGlU98wV9OxBzhi843U31egTPnUTddCYznjAcbH9BR7LPV3rb5UpZXRFvjpxZweL9Gbz7OtdRK
4PLwBZ6XpeirVglS/w5IAvDAy9MzVo1s73rLZohFTm8nVZns6gP/9kQzlmR2Zyih4VTVZUPhFlam
PlwsPYQqaaBwDcBQDZ70idCR+/u1vAetUXdngzf4lfvCJNKZy/laaRLz78sG+wZFbq2i7KqDd3Xd
+fhgyubGWf/Ki5Rcjoby0gpectvGZPFrLNklwU6SrE634eitgwR/JBQJjAP5AAXqZvXAOgMeraBe
jQptd04ZxK6Ie4ZM1U4RgwwX6ELX/krvB5cWkCWKkeroq0k5V0wpp3ARcwcErCZeQLWAZlHBVV5P
p2cA5Y8OMYayb3+FbL3EVnBoRFpV56g7Rsdf9NqI6R3KhHGyzrfDjJ0wMHpg1T3UnqUaIfWTBjtB
yoOTdrb579C91UTXLOviE1tQFMUa9IyAlzYZJ2fqOXKGSP0W6oN4MgW1cLTV9jGY2PxP3ngQ+dlW
xCLfQRqYjtVUZPe8FFAf+8K07BAwU9VaEr4B0hu19/iitSAIHlCZU5Yw4gAQ1oH+tq97Dd1vB0NK
SapC8PuMtzkmXJZksPRDgyOVny9LRTC/phapl4L4JJClRWblHw2fDW7PhQ/7OtxcwUiHDYe1pa2G
LV9s4Fh+1IhYchHGRW7prsFhhA+n+DgUYl969U/h0XGSZ1tgKU4ZgukYQ+b/LSXw9vADUjDR4bhI
ZeoDh5UpJmDY30JqFSQj31i7xFmzcH/Z5GOHVgHI1/GcLORAKQZWAbGEERXxxH5kvJr8dOdOPRSd
B+HJhAP9Fjl0+zZkTKbIPheml4tgxEeWWuDvhKiD1Ks9z2AgPgr+olraNf/JJCt11BPAvfJkMMha
rl/964AH2Jb1Fefd0qZUneTSjxExh5DsC9ko9IPbFBlYo3hbfaeQWxDFNUO/Lng0KiXxFVZcuPda
GeyO1AOA7+72A+sjG7RfwWJbB/RME15oc4cjbnXtwA+BGcsgjLqarT9mqNaEV2kkaup+DiRk08s8
OG4s0ZKYc+L4RJGQTwPaCrRj3pQFtOTVZMLHhBeq2HQLihPYDDqqW0ecT/+ZyAyOWhnfyFfa5ZxH
ZuebucKRxQWUvjMX5zU0IiB6aToF4VoUV8n50cn5652cytD7LrooCUDHHXx7k2aFiTc/lTkjjgNp
iynxAPiRzQy3SBIHl/ravR3aGrcjtzFXNtH31jU1Na/c1EatA2mxO3bH86wosrV16PCF8puxY8tg
TlYTIpblCFULwkGO2rtAo4yZRyqhNTTWqCrEzdppvO3IwFa3NHwMCC9fW5SKIrfXtiiHG7pvZr95
Gi3MQM/C9f7qimjNDlno8SM0NyfrYKnDhK815WPbLaD37iBj7YkFziPIMjrGwazbWf6KgmV5kxdv
WFr93jCZOI7DstdlAPOgmO2D6xu+5FL/lKi7+EjpBIkIEW0X08yi8LK2nAWsGxuiBfdzbNjxruOb
XPhiAtHCoizqQbO/fcI29Rv1ZP21JEZMgGxxsEqguOWHsZeLj1GUtTxzwbCvxSJ01w8igtMb2KfL
IvHU8hdWwCxx2cxaOqYTWbpuU0Lt75oJZFs9DNvihJ7bla8AU66HsHb2d6TXYTH5GWJ6XOB/kvOx
ReFPX9SDO4A6ax34dAmGC54BF1uixL81TtXM+meukRTA8q1AM+VIF4r3t1jylcf0jNPOO1PmQXuK
uyhucSFruBUOx8cnmGBWpT/om3iAVJDknRXchCVXJejv3fk3pqapYfnokobBAASpdubQ0vrDG1sK
2ReExMgAzT+Q8DrWzcuDoTh0K5813o6Hb6h2pxdQ66uQU9+cPLXcv3HyM9vMv9ttBzgG+m3oxP1Y
9eQ6XT6DqLPPO+/DYvihcVDtJ32UynsE2giVCLFBc4fC240Bb77lKRJy8pe3+rR4v7cTe7E7wzoR
jURJVWGBarPHe03rC7FwyZIZ5B/MHY7/CJcdVjMUhe70AwQjwQIg4qFE31MvejsiH/l/8zkuTG4I
FkXa5o5WC1JmPqWYp0EV7ojyCDL6mxLsacfNr2ig868HQswpO+Du3Ii7559dw67pDsZhYaTx+akI
iQoBStKhZqJweyUvJtx88ww5atLuEGwOBXVjiD933t84gQj7hmxpvZMOK1X6BJ7q/MC5dzavaxsR
uuMQvn0IfTYmRXNZogESfUYnu3T0YFeLBAcv/REsco1n+hhZg6tgLhRJCSaiWWl1ckygA/zFj6T4
R/IwtHcOFZP4pPFRC146mNVwWS6aQ93SiviPV+P7Vr3yv+bYRpfqrFss7VwaeKsFE4Rob+KYXkBv
1qOkynbIdj9bdt0uNRJ7Lh3dcMRg+4lvYDUnKZCVrK9OF70KpMW1irfdUbEafgAYzbHZ6H3SSgBu
hA1EzrCHuTaW0WkPkB2bZBxtVfUeQl1c4Bidge00ChsNIIxuJqbOPmLDcOhVgs0s7URk7mhMy+2N
dflC1kCHVfPGgby3oiKEaNUlJ8TJk3B0PRFxo/PLosjQdJSHBdiZ08du4W/fS2/OtoS6JdRY4Be+
2Wigg0FxOoh9ZqP/fYSyKZnPfkV2lQ23pTS1nXgf0REHlBL0iGKpl3VI87PxOWeFVOJaLo87htxP
iafbGes1T5y+8ZujpFeI8zga8ys/ShJBLeA4scUT1g3N3t5U2ffrlZMTNTt/HBW8XZJlmAS6o8F9
YWmtoLQl10LLuf+u2TNZuAYmhVVU5J/1xSV8Xgkjunad1bJkBF82sUeqCFmFiKbybkyekNkWU4d+
AmmVKGK1B+OeKlzFQ0jMVXIudumnhzL7ziAI7Jst9pyI3AYjw7pRZDWm/nLgUeiqDvLqjXeW9C5b
ehsX27Z/06fafFAMJrppgbY3bFLCM6p+OzUPbmyP+LTWzborRYqdqTj8aMmiH/Ai81W38AvjFxoR
c2+BNRCrSoaMg0mAp3hg9Jqtn6v5hTsFioiAzKt/GUvlyTaZ5pOMhFIAmNps9vH/RZhIjyfL2HhA
AoZ426k92DuNFD413daZHrpgqQ6jjeUwDVGU6EViDcyHDn64kaF5azdLqjNr7/tejdeF9rWkECK5
CqJTqivbSqMv3kqcT+dxhM0+jejP5NoPAsekpKYjjQ9JepT6+UrvNpex4jgFPD5EmsJqN5g2injk
FOJfERGBuhUyEo3W931+XtPBw1SVUO9kGnZX5lxEr+9DfcF5RsKJuIC2KPiGoKoj0CANEoyM0XNN
Po6ZxS6hczuMePXkCm4DekzYTSc9RqxvSCLGbOVIwtj0slmn4WCpZUcZFHhefB+9htHVxI4qurO6
HIJ5RsB2/cUevh6V92SxxD2LPXMNPBjUn6Og034tyq9X8mpN09D7rSQWzI+7D2vSQRbHScq89ds8
jxHsnkgBvPc5GA1ReEF+mxJlL641z4xLuFsumTF2gSnKZaLnUiH8nMbdDa0xL3Fns1DyRR6ArEiA
ZsCktCUvot5cYry8W3HDCKyJoPAZpIali/lofQQbFaAFG4yudO8s8L8u8ORQ0q4dfS+V1m+aV5KJ
uw5kyRqWxl8by5qrtMozTVECujoQaGDZopoZ9dN6sRZsuQKOqRSKKdGZh3k8bMZI4dOw8d1wTCaJ
MGMwj8qCZuHegkts5E/3exenl+G7KFx9voXnbDEaoFpxo4LdoCJm2FGW+TocQBGtFAuz2CSVPVK2
okbZ8nFYl8WeTcwAbpkGaQsPjbpNjRQnGbXFG5zISZXlcY3YZAFSNU6tSW4nhB76rrYd/oholI+I
O6a2fvYEU+sALTNxJaO5rT+yK10ikBFkpzn332sRNyFUV7Fu+41XiEm1bu/3Suj789cikB3IZ4tk
Lq2q+cpgLNbcZzZUP2RFP1HCZMoHweJTN0igbHA3CTNi7iUE3YK87UHu97XPXYox2owr3mjpL1qO
cw/TtnJ9Puyfokvs0t6GAjWi/j0GU680jpH3oaDajzc3zSdE30ei7S4gQ2NvGb2PlPxDCjCVVsEw
ukBNt2PC7+pi4xWdcnIbuD9eXKpU71NntQrgULF6TtzZryP2J7EYP8UESE3B0llhVeXGuWkLzd9c
F/JTcpIlkjpWwHgtcL5qSwtzCCWPsisd/1MisV5SdeoH8IwU6qk9IrpxfZ8ATpqYzp0HDm6r0NJS
TSJizxYwIf61nhQrG6vGd+JgEwL+sVdYcGGGrpkXkZmFzT5L9569q+SmrJ59QUlWj0H90hxDiiaT
ozDRR1XgeH4iP60W1dxAFPlVy5bj49JK2Wn2nMCJsDz64gcCsxAAC8bc6SURvngEYuY0wtjuQ2vM
mNRuD/NbT9U98F1cwhKWpw8FCNaN20yEjFeE0xy4KGA2L/E+/6q206puRiDGstXRmwo4QacAynIR
FaePu3TAmoaFIDFB/qM7svNXEaS7KaX30yKvWAC4GQoQy5WMDYvR98gXqM0EPL4lM0SbpA7Oxgs5
BN3XoFkWLbu5Wt2sgWHUfmmc6+y6eJnR+2nhiv6pMsmjChXwAtbubA6KccC690ARDFqq0TWIqxud
D8/zC67ekqkZiv7nQAvv/KOoCRW/7c/ggWWDxk3CBklF2PHPacX2cuocVvbRUUmZKJMB7pWnbTAn
gL2VrGcisUlQmF0UaVGkPq2gQQ1HsKJTasYOppYVEBhyNu9b7GtDnPjQkIdX7UgqmuIGxrOtCLty
RdrF/hpSxKLCeUZVcQX+PbtZCxQfuijJgf2ox22jXLAcEP16kx5CN9r4BzDkSe77gHhzfC+0jTNN
gAr2rmulpfb32HiGyXRCtaoVWSk16/FrO5KWGEuAlOMXf8qvkPGMukvjf2nMFVDv4Ebm24DoKxhQ
23t0XBJPZCVnxm4B9GKlB98XI+n3bVSC6CXkXDXs8F+iD5+sdlSqKrtXCEL5ir2W3rPXuDyugOw/
QJBJcHQcOZUL/NgU+R7r9bo+IVV3NS0HxD3kGVV7RVds7tAoz57WRX8944tAMSvMBimmpD33+Jiz
AbFWaUhaEWJmmt+mTjVEOuB9UA6LPfflqFjdHCHMkxvrPP00sguGNUbiT99ZHbVmFtK3cGKNuDVh
9U2B/ym5Rjc5QzyPDXoiqjVo+WGOxslHpOWmBfgoBEaaYkICfgsXy2TZnpHjItziRyn8ftSKw3Eu
414fQGNMWims7mytwprXvqmvQ1HqOpwQVmm4tiaG2grcg7f01/hfrkoL3R439HTMwut8Q9ZeQq7o
R5AnBEpcwnG40TsskTOuor9yREeXBfKbBxg2DL2f8rI7Tra2uPu0S48Zoq1yM1eXxXUVtYl+q1+O
Lae6o5TFSj2S3KHHZGgr2YP/g9PeaHzzUmOgz6LrDDB8ENHXFPRs82mn2WCfX2LjyitjyN1IDJd2
f89l8UdgXU1W/W5zqqZ34Ei8MpMsI7skrGQAWaMIRRQYKYzU7/KJGU5f+LM9JIl7U+f8r5yLqLhI
fF1wny9yjDhWEWcQdPdCmkX6igMAC9WcJxR9jhhFvojctv99NqL/Ggnxk2VQ7cL+5P1cHykZPuI4
xAJn3T+frFBAu9r2I3GFPshaY69Q7IdmpX2VmAyxx51eCL5opYFIiR2Ih9BeMwm7y0FfIk1lLAVK
xZzFxSLRxHPq7piXn48Ihr1EW3B49YAmdNjkelStUseNDyXJ7k4ay8t1dIB2wNMZEq6m1dIHJv04
g3V6pphhQcAVc+5c4WbWv1OklmeHzb8NcJr9ZpdIamvp/Lmv52uqP7h6T2zOQLl8mCmC25FoxI8i
t8AT1vHM3D4OO7UF2cgYi4KiMTd5xGNVJgOx4xDg00VYr2K7nMuvh29SoZk/BNX/IyR5k4N6CHzI
G1p813exjj4r7Gq60m0i8AHuyQDBMsUyvfY7YGNs2mawHAnJDXHb8yQ6gnFxlMhQ1KQS6OJbXVaP
cDT+4khVQ+EPoXMgrs7l/CXMhTrWoxsns0NssLCmd6Mc1+54PeJGENWjAnEc7uQWVHGrzl8VoVOL
HN9x4LCQmZcbSSYMFwyIOgkcfKwnVJ3C3ye7au0xcXm9YJrHoekYAhnja2w+68MeRexKkmreEsXV
Qjs8b05Pk33EtJKQzfpkJMpm9UDQwXB1uNC7ZkL/qNCiGhwpVS7UCBOxlQoBiPq+z1DvfXN+1ugm
w3FGzP7VQYXyRXwQfGYHUgGdEYOND9EIXj1Vm1+w8+6wpKPi9fw/a5RMaVJnKortzTCvjBcxlfFv
QmG67Ay8DUTlzfIqPebFm4JOZFHLoBZ5/2Z+ymTO41ZvgbmTHot/sh7S8293vRdMzzYH4k0m+2QL
j6k7nLtk5lpPGgzBCRC8Nx3WokPa5kqb0almsEq3Mvhis7ZDpxuK1Z4SChe8rT9bFcYBA8IZnnV6
61UXZcJbneGv9sWa4tccNccH+ey+kQzENt4SRB9W+6ljkTxPql6LES+1LUSps2LwzxQdZbcnCb8p
r5QBKMnVGkcj2t71HLtThlBSy7+F7i5+vH0qqPUAfXBmZOl+OBp48XtLeAE75tWCeZ51vkeSI6GW
cwTGrtkN/VUy2tdxDP6mCP2whM5fa3L7zQqUGgO54fJs1/wfEpKHz89qlq+6YSZKfqrQu1azKOFE
m56mvKx3sA33R9JoXOL3P1wu83kJljfm7KsgfJAs9Zwwix30B4Bh9v8uMEFr/sjfogpoBYjeD8Do
4sQe/oDdmIZfvNZBpoYgQ57BC/D4avXJMY2BWoxDoNqHA8YRg6cN31gUEBc5fdjmEGbVETwpoPPB
nufW6Mso3V9OIYF3ew70jbGCYR99QAbXVr7hnMeF1MkqX3SNDgOgy2lvfX9fzFNcLT7icCp7vWso
9Zmbo48Cs0sTD18nr/4DXsf/qsI+5ORn5xCqajqp1VNINtKhynFjO8h5GlJJnrPCAhfSO9ZoQV4L
DPM02+2Gk1ux5ybKNrnORRp/5IKWQ2t70GyPx6IZWgI9N5lQBrR6Igy698u9dH90IewrqWBifiFN
Yotuxq7Y6xoceOKZpp35M+GgOJl2Ye5Z1YXYObZQ9jjsk9ZnL+a3xuRyr98hSLqtE88A0inG24FM
kOSILusQYIFBOlPOiFjgk7xMpmv2jl2IWfS2pGIeihdjBw4pfX9neuk6q0YUVOvm3Yi4tbQ8a6MJ
62NnxgIK6HroI0FjPnEy/xx8vOm6v6I1hM4iQTepvyuVnDlpkByUmGD4MjbH0AotGtnl/jPoSprL
bKhi3zHYZi07rW7o1GtAuj3r+Ofnj6hsfETEf4LBK3yeFn4BTp+SOqYZ9qcJg6qQc+zSPHo/FoB4
XJHWH2ttLLO1CaUpZOnnh0X/1Ow8lyrf50pvLD1f29W7UTiYE+Fl3+UZlfvcgg6FHa13cSREe2Uu
abIbS+kUm47XrQKxnKi6c9fbDU+AqL/pRQkwwbN5mzcJQ6eeof9Q8VoYX9Z6btUF9P9mabJIeuAX
nvCfDirJGEkEdBZ490vUn67OWfFaAD1Ws/NJlcy9BdQzft5/3eET4t4CgXMYGm8/VnLXIurmUb1u
7PiQsSgebN+pEO+1ttB5+8+hULGSjPI+b8iG8nxTIeyMog7gweKdw5SW/buf0yjuhj4VMxENdNDC
TI8uOUgABBbyA0I8hOKYrU3pUGYuo/HzVozH5+NNIM8bk7HMeSdyFDs1w67xotlKVHiKfDGnb20Q
vpxLRfjOb7NGI7QhhofQK+n0teYQipm+VyrJrUnt8c2/7v8vP+/tKU7NKww0tbEBaM9OPpOzwNPR
1MDUutrIv6cJ8daX6Sx/XGgR+u6YsHhyZTxa5zKNo9+cvA5+QIU2Ibx7qR/4mxcUKHJBb4Kf/2WS
XaIS+klPmoxQXZY7symONZ1jvta+/fyBuQeSTBEGpXyhSLobVkEQs5pElVAWElaBkm4pETlfKPxg
DfyO3IwSJRfxeWN42LyeQVoDGCIq3hZ6zkyU37BuatQYAnrqhtrZv9+bsWRP3Iu6AA4tEybGtig+
rxqV1T8otDdd71Gn8em7+6m3DLeyNLoITLSGDO1tH3lU2hxenFt7uV98qLYCkJ9oUJHNIM0ZRdsJ
rlWKMYqpyro+zKHuYrejKJfTALZv1YKMH0EJIWSt4WJTb8WtfmlWZmMzBidEU9ZLKrmtQX6yAslm
1YvjTX61y5p9pVSdVY3moSdMjQlDnMzacvIRAMxcIhrSyebAjMy0h3XAIWFCw75VoqPfPxYIkHYM
wvh33q6//tAOqc4k3ko0d2w16CkeLZs3vmT0peBr2cfKYJJrUQHGyDztxmpSse/EfcgyVITgwQ/U
GmxKRmbNy9ErcpMuIIQL6g0zYAdxjaW9BZdsvoeD8UWPeWQmpMvQpnJH4bT59nM3jzHOxOyAzpHC
cKCxSmY8RCVgV/CV/To8yh9yav0kXyrZXa/Ckyf7gT6KS8OBZwDbA7F1a+UVHrrGG6Luv1bcAO5w
j7Is2+mmH6GONMpHO+QK+Pi7Z3Kg2vPlvrdpComyx9XarPhhTjJRga8vYto63EbBCtSZjFIYoXDE
89OVHlQ5fqN2SRQZbbxj7GlPI2DSmheTUG3yYvYn+XqDT10pephkf7dP41NY2siGodb9xge8Guj0
G4VD0sa3hNtT71Cd4h3AmuBctWRqto50+pOnR+jBfWKFHhylCb8/CaqL7qlCWt1wXrBhYud9GYVw
b4fm/tEOVTqIhoZ5rdxeB2GSvlZcAkZYgyecnLuRKpRyBOXRiEdOdjRp6fqZyIWIwc3Co8mzokA+
D6FSrJK6dydv/ARF4l/rZ2l/+xbCk0JLGhxZjlczKQrAbHCS40f1wu7QanjzsuXwIVyI1sjcnKEo
OuLg87lLC0QovdIFO4DCGwbmrWCs9Tt/Fz+7eCgf6dq3PrVlcoMskCr9/x6BVthHfjo8lKdDXFIl
2Eg6rEGacy2ETiN7Dnq4/+XRf4szsTYeDRSkqMEbbRcH9+fbrEPZTXbG93siWDc2vOVM7h9OMjVA
hiCyESjHXu8Gx0Ox6+kxzZSwo3ub7vxSkZ5pgX4ldKYqwAZXfG27QPAQ0XsUKxnbIQwtGzCYsjXg
GjEpSPZ7ZqgcuYJVoghJ92v1psmgR4XKke0eS80v51+UKWo9j60J7xT26quQrBc5SxbpXmzvN9cg
TTpqXZCY2mhBCYoAbpwlFAQBswLJ8KZB7v2Np8hCMh8H+RG1Em1yUkhwRCeKAMnQQGi8X60/Y233
cuxjpJGWpmjpDG2rt9L2qYTz68EydUS7YGb2sfluzccgdFn9F5YglQe+oPvm5TbHRGOgh4cLTsML
fBfwg92JmJFBdeylcq1H5DKxExbznEcEt+Bz3jCAFcFnwvQ1l9gpwEmean8zKcYq/OMeu0HRnpmh
L0P1fCA7IcqXnqMwGMxYUyATsfjgXN6Ij9tx675BTaRk619CAi36mQItdrmo/57rTaaMneq/T6Qp
I4zUTz94pln/CcjeTT0GtfFCUkeiIYfXQY5bUY22jaJV6z7kHtMNWOaege+yJxTlWrYWHmxaWmTc
eJSHOZ6fjHAoJBUIpktr288XJ+byNoE6V6hnf8DiK+oXqBSao/Kn3V03YJr4kSMx3rLzTXJQTSgS
ajzt6FuxwR0ahdWTEoTu/mOiHPr58V4i3G+oVWdZj5Xccu1fGdlOtHJ27EyzvqxOr0gm+EDW+sOx
llUH71hUerjeu7vD81OE6lW5ZWt+n/mh/CS34tnS8sIDfR3aHZmOFWOuAIcx5Q9WlFaP6sd28D9G
9wWaKenGN6yQiI3AncMrO3VsWFIEdtQTtvI1eyKvSRrEr1Egy4iqc0hlpdNDARtQ7xNcBw6aZHjj
sFTNg2Lz53c58M0w72D+U9DCyw+jThgvrGwM+BGXeOg4PJgbnZTPB5qBrRA1aFpGhwcU0qjVp+zh
YPcuXTB/FIabL/1Yv4soo+t64O0VwXgbk/oXVhumtfcivMRG9AQeD4hxVBXZ7H6F3WN1x+iIiIcR
BvD8EnTt0GfGo3f7gUjOFSfp2VoNWMefWXBndE5AKXRJ7yXge5F7ULDKE+wOX9BGvGGcEqL+wqWQ
rZ2IdXHbSnfkbXqH2OFlGXChwQFIvQli84TY4osshT2KWbZZQx9udVE2iiClk2CldWjD/yrnf/oB
d4AoO758SSFsaQEu1qnFxQh2/MzwMkXxpB9aOFLasJOh31nG742apKMSZU4JpAsGhjZzw2/wc8Tp
IByw3d3j6aEDmRBF7MLRGDsY6AGYHFyMR+bZXMjSZtPtQKmHGeprlq9W8y8wkfqZ8FDoV5/dwSnv
k96x+cWrgO+5d4Nnhm+oyb4pw+kv2lg+j3B8rI/w/PfTsJn+s83tqm+Ui2eQ1V8ZrO9Gt+sBQUhU
FW+BXMvcfh/aQSfMsQeXqciZFBO3HuKyLUWywjOSma1Q+8LsjQx44aD3/YQnoRHUcOoknemBWjUG
i5ZK5QM0ZGnPOCDsC68bByYzPkKAKEZVx2/XUCsbhnicAXNaBu6IVvrY2+LpHTR42+Buf+/8C+T7
SJdtBDjeBHN4lkwpGWx8cdmb/wx3nEQlnpiPvZvCIr4mTidCsvuBFKT+ma2QH4JpjUU8OCRewP7k
NCjwRDy79rkkOe03hC8ELQTQkKLHBNaYK9AIJfdynaRqRWajXqh3llNP89bdt7Ji5jF0m3kI6KaW
gnmFzJPgNMS8AFYnMl2yMWxvZpITFxq3JHVPtH+NOUzVcdPHKyNrgDQFNXtgtNpkWDE2U76FZcTB
7BZItne2KmsadTY4MfyROo0vQp33CcPlzLA7ofA1c2mmdRAfVGhKaO3WCR9Tp7myjt6ixNxqakLy
5DwBQ5KnaMZajUiUZo6ZsCyjA+6Tleb0aeLOT+3Fw1WDp+zlBFPa/MEcTNKqIZH0ukTErBGX+WzE
1HPn1DaOpsh/qIut0HfSFK0L+6GuQyv4cvHtmTmbwGerLbrTAJyvWCkvOmxjJ4Q9u+ulqvBDmM2J
PT6YHK0gjB6XWuvS+tfrnQBYr4Jii/xcCTd5llwMcxcpyKLHfpydz3x5K8mQb/A+cNIpBYvW5N4T
loe24gm4bVRA9/2CyypVu//mdpeWy7n1kuRZPUopGYkqBYlnViNZn7Ucwo5B5wUAOjWbDdrC7PSc
AsF9Oxeh963np962SWf63cp+IrZ5BXXcVqsRuRmlaULttRhVkLlEeONxLytzKXxEOzh1to4cVrX/
3Ze1PmTkaZvf8xgBqFFBFzd+7aeB9JRmgnyisqd4F86YpCmCYXt3LvdHC44kgOdxNbdI9R+uHdQD
gczLjOTFEN75Tnumb4gvFsFDy0xLI6IpXrnTQEPphs8LKQM7Fjnk8GFJ4ydCkbXjxzpDP3DWhKIy
afPjJtOVmxS7WUt/MxMIEdTVda/FuwuUiq453oOkWrIAxz2yTnRWoXDUtiF28I3YxhJWWOpx4BHZ
r5aS6JmYOGa61XMZzFTWL38x5s/eQ6nqGO7VDVDCiWUwn50JfW1tJwIA9xctRNaNJId7+PXba10w
1TaMGyDIUA4P2neft0P1hAvv9+pUtvQmUAY+CXjcmIr02TkR0bJia0wa1faZyj3PLoBYO8l6E2H6
5VqwYsNBw1oM1JrnSfBXkmbRK4wUOsAt6WW5CL5pcfAh7HE7bWGDzIFn1V9V5xidHrTOdrYRzTCB
kffakEasjuQmXaTKsYIQ0d3dOyvvMZQniwQv/z9u3q9yw2M1umm1nuDjhVKN0LCf+BcyX8uYng/h
8R9IOEn+fcf6pouxVNJSkvGk9d67I2UGzFDWaLBVy/wcmV4ekYEG70+AENJ+/vMm29IIXe+MEIoM
7QcuLtlBQIePdR1hg0qiNgHL3TsHCHqxIref0QtGtWIo8Uk81QXaqjbn/56B+X5kE01fcoB0Xmr/
q0KBI38xaQw2CH98v74Ur4GQprFnOYcMMZwR9AXtDYgED4aYTxZUhV+CQ5kv8HYU4cf9avMjHR+I
SLGWZDbInbJ8qeeYlF48eE2elKZ+buIH88/wUTrNQPpSrGutR2OmNDg3f2pbPBuRv8CbJ9oD0FLY
YL7NUc8AdfeiuytOc5oIcERZArkK/CraAoTDkXB95ahWa2YHh+R7o2gOGdQSGy5T/bvRzHWKdNn2
zdsBSSuYJPyX3fxrc/3uJAPXbYr5m4kFRz7MbRWl6kj3Hclq0NS35WVQ1Ak2peYr7dV6QcdvmHL6
RxKes/Xo/V7qF5XiapaOa1v7QBNaWr+9ziSeQ4sZe3Xvtc/dlzNXZVsBUEdm9Hi5DtjVNu/BRfjC
FHuwFwbtWYNMVICbZtkmBP801XXsF6QCMFrF6nn9izO+vWGnMLkW2o8DSyOz6buQP+zHH8ei1f1J
mPWHJgar5AQfbe8v0OGIOUbJrkY/GxmKeoXb/uvo7bhVv6JFeAm6uZRsIU4xMZTk6cQzQ7ZRRhEG
CRG8wNhJGCvWxICs42WlyeK1otnjWbN+BHAyrXYGM39q6WIbwilAOJcUHxdwzYeB+MINORTjTu+W
QLMoZufMGJiETQKLWt3JdamAI3SXGjFG1xZ/GjJ/z/hMbrJP4q5Y+qAhaZ44m71vVpBSwnYgvutG
uxLxlONXYZhBz1d2+sN+eQsup2f3H0j6Wd0mu3Hp5/A+FmJFteQ68z/P1UjxbnsWfJM6DEiVPSjc
RvfaiScB3/MEfd7C5qqqc9G1c8jRZr2suC2HnSteZuZJepjsL9TEnWGTOD9XLPmHGm8CTFXp/Gym
FO+jv4Jgf8BNc+hqayh3g8uc3KChEET9a809QOphVtz4AKuYLPq+qa/GzJHpCRjQCI+FNHUrbhmU
AfkrO0l7bxRP3Y0wzZtsZVvbuZlzqlNYIn6oGmF8PX4KAihIHsat/vw2oVVodfWCGwPFRjLc8r36
+TLsaFqNnlnnXZdwZYz/CUoAvQAXn9dNvghOZvKrf/AfnvF3O2d/0f7m8CiVb5SDO2aFV6mF7cXA
8LA859EMhvy6cCOt8zOBpUqnWP+dW9DHE1bFe1p/klLupmlwit0Ws8wrH4N6n4b/yBc8x+qp6Ojy
voVisHa5PUUbPWc9Z0xaByXd7zFdGlAYHarrO44+U2hv+EroZlnGx62M0fe+mts3QRhcerHcgfTn
x6t1zArKveBpBFVZWu/Y4TAHCEERA6GZHbYCd3vyClFS/9UGpWta9ghsE2ww2Ak4GZMERQxq8+UY
hBLom2AV57Ck8kwhCyeSK5YAzx5kS0fJ48f93HtRQIBxBMuf8QfmfB8VZdlqvuOU0/bJEz+P983k
jEi5TMirF425265Hg4HM8QjUZM/9PlNS3B6+7yI3Z67hj2QYPQJZgGSW/qjrO9v9Emvw6yErgMOU
alhs0O6ktTuvgT4G0EnG/wiSwQAgzIR+mamDMOzT1NQfmRQjZSS27gNEk/4qyi9DPmJnA7fkEmd5
ZuKpGroCuVv6lB6IAEB1RqiXYAEcvGZY1Lf7dlQql+VOurhRehAqPu1RqMfjxOOD9MerOgAZ0WmX
okT/WDxVaL7dAFq6xHSaiofUwG/CXNino9PWDkYvcfOab2S5VjObqOoJJbrPLbMzQclGG5IIgswl
HW+RLGHvUp2TZz2qYY0kjm3grncMBdVSBgEegdCToJxypySetIfbUT0QBaEzUCfw4SXANtKVzF22
jd09ITTMfdkdnN854WKSBzEZu76ZzXXQ388ddECfrbov/8Tl+MACgdl/9h8RcCNyapLekP7MKikj
ErkGBFSHCJtVHBN7X2c8TVp0WgwGWPDhC0ku6H48w+HAmDwRRLFs3cHzGREAXm1QI9cY1GwqqAD/
IUpVLzZuVcHHdbb1F45zTKOZUmiHpCdxCwfQmDpW+VgfOIAF/oteij7nVQPP8AHItPfDZ8iiVwsn
cUxDkbRC8lvKVGAn0iFKOEWAVQy7txU9Z2AyHdcDY3W5lRiSNbtZomjEb4hPOe5DEOF+16D9O7ud
56OIfYEgJF2qsHnV68xuw8XMPpObmOOlt1xCtu1PXSB4T7EyduehLRsClbFNlxeLXm7n8gOGimSh
zEy4zQ0vl02KpCbdl+Zvhzag52pq0Ip5miwjL7rUDyJr9Fbo1m+JAPQyaJQsgnIhjHQnyt1sB/if
1QPv1WgxtAVuuF1d2j7QYmaGIqNvovgzWl8zslkSj8W3yJIBKy70l+kP7zXmUZ13vW1K4+bK3jPX
5FPs81V9dnQ59/Bm5R+G9TvHS4hPRih1nqreg7UOD21JQo6LXahd0c5s/3NYK2fXYyVEkimTMq5c
jNlVL17ShCDokheCGn0bvpZUBC3cP53uhpl1ifOVUfo10e1rVbkWCUHjOWwjp7c9q2GNaXiEZ5kE
cDdqoaRqEd0LfBvggWauetudku6T4gUeW6R+bzhcAdzUz2ufGhMbWZD5ZMDjno0ZktG/pVaG7VHq
bLnL3nVXasqPutJY88XZiZZEjAlZ5p0NV4kTaLSZuUq08S0zI7vgVBdxLaREhQCNk64iSnl4Vxmh
5B3smuAaUJ8DB1++6SVZuRFsq67pRLBv4IqgOC3FOThW65Ir67xDKiHi/FVlvNzJu29Gu+fSj22J
6LQyidLUX+ctsf6aRHMK+vT3y1Opu29VerpXtuoQiVEHODUoaEf0E7OtTMvfIb+YO3pO6ep7SrjA
YqBG0lD4ThRjWpPGuNkVbOur3O3iZIuLr9QxkUdG7Wo432DOCyRxV4OnZ+LzYAD6Ad/l+71yC7jq
/IS5vlvErOGt2EGtLYs1MhL4YAlEtYVMDtkt5z0JOfxF4fTNCOVOxMfDUcfvN78+4cIqwwCwP+pQ
xSg7sbLi7ES5q/R5B3s6/+82RRH4dQ94s8ZKbZQk0gTAv4HtMwehmtwign0Ob6LAOIImaNzW0jDm
db7ANljI2KlPz5S0cbXAw9SrvVhuHTsJi5iKDq+MY07/tN4BnEX0Dr9EzMAby9ZIiUWFxu7U4xje
qywDGs9qPN9GDdayb3+9Xttpx52atF9bbZTeoV/CYAeraNIBQ/B/EHH6UUOx+LZhaZDvHgfE+9UY
ZWncutXTjQkYbP1Fafhvzs5Dj9GAgEL62XAqs3rrYqlCyTF/k7D47/SztGrIKTwiENy0Wcyq6rAY
PF5ZBGF4vGaWVcN0wrurBiN5BH3ed3fKvxl+PqwBQASRSnKB3ThY08CLp/16k+dBUWh/GZl3op4r
iYh8VK1D6mG1FBCeAxZjR7zbcyvCCXhn2yGCVdxIr+5KWTAqTtJr6OOt55V4oATUc+se4BiIfE3/
lY+m87sFcbIngYRAZzo6/0hE/D0YbG2ziQz6hl0T54pvdqiQosIDE8q/OAvzM6X8XhjiN0/xrppq
AmfLUL3Z+8/RWZCFH1szmwsIIPjkTDiumXo1v2LPKGVF1PkeVsdB+3cVM76wTWEDG3MXDx0/f9/P
wqK2HJtFXPnkpcM7tpiLCN4VbMDzO2vc7PxQTZoz5bACLosfM8ay9XvZQuD1z1Qhr3m13YLkIQL0
DrsDgsaBQ2UKFRGmZ/I9E/rx6Bhw0xphGYugjQLxI4QM463u+Xz7GQO5YzFmabd9K8l5Z2dgV8Nf
f0M6Rlb92UlhxCcAqjykjzbL1Vz+zKMNYTQc7hRvrQ8G53Fjn6sN5sZrIbmVfzvWQPZYxUddTfSk
6AvZWIK92daP2AvrInQi01+vXwAKwIrAkdzDjlPzo9fGTMjU5Fc14wGkt7qICIWUi1KYnDx1TiGG
Jmvv4ULWarQtiM6e2uwqFbrCLErJ0dGd+LNu/1wu06jgFHx4vcEKpGrv7aVLWmKqEwOsfNyGrfLc
GQ5B2LRbUBIL9pyBTui6Qgs1sXfuQSJ/I5Ug6d0PRJSk8JaT4HORKpKHgKLh2ilCFdNNSG4gNWiT
33sJVr78e3AukFv0TQT/L8XUrsU7FNkpVZ4IfKfRfaor7tzTCz93cTfWBz5ajpoRfkc1kc0ihKZ8
yFsIYUp05UYqOgk9SSondtkJj2vyQZum6FoNpE7vrCJ4Mu4pEtXhwBJIBWVL1K/lWaoz+NsClXm4
qwsE3OxypPDqL/DRL3fCiIzOqxlmp7n0D5etycL4BpNUPqJ8XCyDmreXiqpdHhVaxiceZOwr56+W
nkQ2vMj+0uyFhzPLTuXASUKhR96FAMm4IhEk7brlTaKBymGQi3QYHBRLVwNrmpxygB5T+0vdZQhW
/ynKgcsEg5jrRIVST5m1axkes6qPid6R43nR7Qe/wf8ySeEFoTixnvESTa7cf/QiRFrhkeyG1/lW
rWj4s3TmwfbbuUUD1oi0MdcH/iBHrMfDN9KBXZcbOT3C4B31PPdhed6Pjlg+hUNTXMjiWydbn0pq
oiCTL8KMGQJUlbVBKZyoxqpg3LS2Hq8HAcACmseYbflel9aAoINuWeCMJ3iHONSZW7CULLyNLYEk
1yjrfYckl8oif2y3jCV8ex16b3tTHM+F3JuFqnlnyf4RhVD7+U81Aca8ErubPmAgjLAC5Mxk9Cth
do+NzQl423uNo+fOjRNUP2oi2wTS1OdwR4feajMwe7YxP6bg2ReEbFvRTntsMSAf9EKfLJs3ngHL
ZzNqQlgrXEAUuyZWko1fgiVDrfyhceq2vUrt64xGs5NXOQWk0UUKLJQ3aGQK/B87sS7nPu7nIFlM
6Y3NEoqu1ma63W2x7lScwCEeFGi+gM2xs6r6CczrHeoXyj1cga9acNlofZ/vfQCAXpw5QSe/ri/Z
WzusITZQ4igYrcIWXOfDxu6VpIyBCs9yKEBMttMZLGhj6i4aL+xYp6AoI+hPNFzLaKkm+3OLvBVz
7yTEOpZHmO4o7yaSXRDVQwDd6PgyRtCc9RLAqSJCbqqqiC+MF64UwOfLoCK0P2cVCd7aKmNL4Pcn
xriQG/qKNMgsir9AVuGrUC4F7cJX4Nc1UVJ0q5Im3oB0+3Nhq9pg3t5o75H834GD76lemhjgrd87
cdHMLizX822G16+JehuQd4t13KPbGqZ0sHKYgC/OPkAo5j4XcxuqBK+hYOm2OjkIZg2JlFq6ijDk
BxaK6FQ5i7GUkVck2QnXqIr3nxM2yS0nSRmh+yEvYCW+Jczd/EyHMCx5893Arf7E/I5kqn6Y8mxm
rpA4IovZGVo4dUMuIKXPgLOLGBcR0lk3wgukR7/hPMQ0DHg8idtCFNMqfe0ClsKQbpnoZVQaHPla
Nmg3GXgsctfV7JzzzbEtSAQM/q9l2lwrzIzr+OSbhh2PbrW12ke9sttU9gc5GbGIQfNLsIawcCCv
Vkj+rri8htMCNamTKw5c5yr6kQUwUJv1K05pmtZfJo2vNTF+XflbStPdOMw3hR64Ro1cQz4zLChS
9Xx03frzVwSSJ6D3CsxsOgj/f6co0L4neuRWkRRpcZJvWPA4QrGLwUWqDdzg9TCYDHQKIPOikLqx
qARk4JcoWjws/PW5Sf/ZC/+5TQAXrm0VQ0GT/UUWFqa5BTFG8XKWf0CS6MAjf5SbgEAi5WaSC24F
Av+NzCJXjA+ZDbbt2iw6lPDkbnN+szAEeyXoRKrvLuFnb0FmmKVksT1Vz7bAyF0f/lywjs97bNhw
GzxH+v424VmYj90+lqvuZTBiYxL1HSFowQjUzSJiZCKYF3QePzgjRn2OqhGijds0RJoKWhjgqwz+
KCLJnL+0A3FBKyFA9P1N4c60p9/AWpmHkjd448yye6S+16zhYzQ/ml/5Sl9dETpk1IBytU6UW5Z0
UkN1U08Jwi7v4WwXW8SPgTzyhN4v0jHVrNTesi5bomcDRIctWhnsOX1ogK9sVD/j42R8KOTeGnUU
o12m5SY7TNjh3dU7fL/nk9aqEbkn17ibnAS1O4sNNVonUVowoFwSquZ4hxZZOjUPHLAyw4MW7vRJ
/EF6Aoj0B2/8Q7/WmC7m9GLtBCC/ELYNDIfagMD3aEKsvgXGlhqL6uP9RnphqBByqEAQIgWb4G8R
TR2TYZF0A3CY8lUUSCw3EErDYHZroyaqMlVRN2c3FrjCsTHfQJ8gTRa/HosEfSF9jdoq6k21Qauj
yKjuKmEO2r46+UUZMbJsD0aowfXZObEEGnSm9A5wulM+OUQ+kyuGXvP6nodMoHsWIGv+38+sEUWM
ACu6sYrP7uPti3KUHL3/CHXUPTYr48uZGKZpEQ7nMeygNxJfb/rvH8s41f4X+pNSDnH5Jgqj2eIC
kBUWthThg5gwt6Pn2ddxL8XaFF227LgI4eTc21WZYnDWttsEY4vaUnOBZXyd/bcajoI/gGEGSM0s
+qWBrkBmkxA3NRf+z6RM1EHeLhhbPwQh8ruz900PIgmFRXkEFmC/wpIjOpIzYWiT4hclPutr8u8T
AGOWosKWnpvw2aoylkFz/Is5OKywlYfThXo8NtMgdkekycS7fSWYAUnvSIdkDVqMgfhniyystP7D
7z6BJJ/dr+8Qn6wUtDjIkQwkRhfCJm/qQ+qV7983XB9JiyLWRlWx40kNXqxFvNlucmx7uN6toaJN
sLO4H7TMI5y05NkvDVeRVn5VxZH/Ph30uB50oeIwnBt6NgsxMUzkauTSuhjQ6euhBOFHCKuFuxq8
d2Ds72VUFKejKibysrLzdiCwWaC2zPbeAZx8S6uR3Xj4XJ//Ox2dfYRPBkXh25hQa2wy8ykWoAfC
GxErDZWky454Zi/HA6yypJyUuNMhenFIZvqwSE6lIH+DOmcDQ6b78S303RgTse8oMOe/4TmQf+xW
27/W9w97HeKtgZMrKFUDmiZqRVAatG28BjNSxK46qa3l3IxyCvDjElZO1yDFEYEaXlF8cuaE2Lrh
7WsF5i6tjBIrSqz+ysIFaCFh2JSPx+GntAEMBH2P1yd+bVE+pxy2kpDVYO9zx5X6tSezDCdwsa5f
BX/Ll07lmb4wJFaWNceoA6TSAcodEgZCpz7Y/CwFCren8oLx95NjV5urg6WUnukiVT8gI5niyvtW
BX+ZiKxwVGTFwkQGwBAkJ2Ilvteq0A3ZaMk2H/qhSp5blf1NuRXGnLdNHJlmksd8Tiuelsq75dMa
DyeiaAfoGPaW7GFJ9k3J7DQiQlvDrkj4Qt+I9bJogVCCfVFn9IVWkr/N5T3R038wWq+Ow2VUao6G
WFs2aLTa53YE+SfZd0ohExhQ1hkDtqBEbBB2vYlba9RhfEDyIHO8RQfnuHCe9NTdtxZH439GCZyw
VQPJcQCppSJEvk9wKK+ZK9c6aW4ysBQX0DcvxT89vpVSLeix0Kpmcf7yRlXBUB6iCIS0DFxRiQbI
3xwUkj9HoVmbwEfWIc2vgQbGVWLoT/u8MV6C0VvUDIwc6zRASjFgDz0DZ3ICIurTRiSbr1G+sH/C
55ip8vYwOFAQz7gmnwsOYh1WGoKNeWm1UxmjEqajv95v9bVtFDtUn8UtXwXO5SxHZmylTjXQSPAu
9olHJje0AYIAt6moFgFqfj0Ei86MzTjfJHb8mh0ElljmFoQaRTiDZcgnlKbNSyUKVfXwntORi1Lv
AQlwv5tPudwzTwcBiti2Ye7hcBfiPTDHOBF9j6qWBl4Hrr5Se6nMFLvjru5GvUEnfEFT3Yhu4iVW
WC5Hhl8Dwe/VHlYBfP4B8irawhNKzB2rbr9oduY5Z/5oTvwkUl5q1AgW328YrLzOK5WXUXpWFgzZ
P491GGi9JKCw9ocnTaGPchXY6N3VqjvTlz4TxuZK2lI5WCKpi9NlYvKbvW3xV8xngr1tc1LN+O/a
o/0Yro4J9caamyo5dpeOfAqhjhLuw94uixiltgMhEFHKg9UTbqC09dkelJJg15lyFyMFhi9ZJrc0
n74BKyGN/S9IBPfbifUCC6eL9ZQrs0iL7aUF7670cXaCEZRLtxgzBJMpzmK3JvZnJEMloSKuWE2p
UH8wDbj0O+4643QkaCNf+wDqtuB40zGu1+eWGPY4TpBkYyBhX2dkOS13GuU2zfSUjuVCy7Uhl9IQ
i/GXxUVFhdied4YXbgc2ExD82zDZInwkvJvmzSsQj5Sy3D02DL1OIG0IBrEfx66Pjm8rJlhIbL0d
PpF5uBWEZ6XHwootjsSXu/l2sC9gQ1KL4uDKRLqjFbcQELu3toADDEsST7egNYkJ8zMSWtzskF7v
Xf9GWI+Ps9i+9LNY2cWNbLqcJX6HvdMREgiCx3xEzVaYBaO+2cnXlmOSF6PlmqNBIZjzifnnit0l
/2D6HsivOCEz/GEHUdv9ojMnk3jPTLAGaaO3dcriUNpAteELMBL9kRLRN7t+6QsS5BXstpRLA5xW
h6YXfy4hUeSBTysKHCYTEamytGeXyhAd5OR1fg/GaBd0qyni/6gjxYOgLSrL52C2FlqMq0HynfkM
FFv/JB7BGifBERWCWhGaqPRGFSpB2bSD1G75V3XmhV+omtmDl8GRLGuHp8GfgW6O/2UJMAgIee/n
6e64HePV7yBTruan+tllo/4JytwqZJc4r1UXw6ewBpiN+F7aYqMELIGZ3lDkai+RLmYJ+eT0vkJB
+6syJrHnOJ1Hz9nxgUeEPJZZ+gWbDsSDHsoAKG1dvLXjx50D375uK1ovEWKJGhIZV65CF2iPgojc
o+Q4soXC1THbiomk9ISKz1x9o7DsHvEhEOLXdDM0LcifRfOyr+Rzgqq9ezsVRs2V3y4p0MjSnLQP
fVBcu5XMJP/pfdvszvgHSnSFYoTBDqBtRcW1R1Cvb/q6BJiEu1Wq9kNysuRVeS0EmWMdgyHBe3h1
8vznl1RpujVl90BRTiXE9tmPFCsIfnhgxHKFu8s+QOtUlk7ckUcigiRjyRmqArDUzePLHub8x5hs
x5q3px1luI0q13zX04NluLa+KfChm8JQW17Rki1cwTFCycQ2clOg+47shzkkOQlXUzhgOkzOWCJ2
cw4p2W9O4b7nXwPvloa/z3OCMc53S9dZafIJXuAgA59e/I0irOEJTLwIV3fc6Y/qcO3GFgY/oy2m
FdhocLzN39QuPhP0H3UoHYteJxz7EFr04A2Q+fnYoTUkLVFqxzVR7pyke+jd9cYx6uC4N8JJSG9C
mRfzK48wHTElcDDq9chbbCa7mu9QXCOMbn76Xpgm5w5QzZOAeql+pitXBwmHXJmDtAIfkYIRBd4w
I97sWMp6aKX3J3cUHuqnRSlzJUYZmDe8zwIbBTsrNc+70zJwgdeqoj23o8ChMT3qpligo8xidBY+
GMsRQ9WuBaGPSlRvPBiDNnqdjlpHD1sr6AXH+g49obYt2GokKgfb5Co7Qe72dTNu+VlCsvZIGG7z
G/zhbqByv1u7+E5VbdU/UJ1/5hNtAZmLHYTAJ9Trwo8sdHz8PdKo654y2QAW9Dxz5HA254tLGikk
gCFW1bx0rlLgXd4Qewj88bYRPMUVxn4pl1oUJxfa8xlFr/csnuuj9ZXzNp00F7G7rsak/iE2+5b+
2QWSO36uaAJ13/vWMvRVPvcEH7R9OVFvLHH3GYWhyTkGFWVMQGqthvlk7kLbSkW85zAlJ+O+JPU2
xx+wbPDdkGfEyEOgTK8pYHSA9wSqdBCgVi/wCb1OiwAY2YV7NMS5HOKYkRYPwF3IJYlrwWEWDy53
q0JpNdRsVYCTHzqEGmDN/3Mc1NmyWCaOXr5OZp6a8tpW5cNGcL+kVRnkeXXjWtdKu1PXhtohTTE/
CTKmJmfYNxDW6cwto2WgekUs6nPRY+MWf6cg5gRemJ7AumAOiso8OnF+1fUPozI8MAAK+m9oIMOR
byDAqJigvJSCyXjuxiXJqWp6Y7fNnSKwwldf1tHsWIuD1Rtui0vs8G5exY5TVNM9biUNZTh53qXz
9eFaGqRjKphtu+SCL/+q6pGaST40KwK3gVROcN9KLkgXRFwGX5OoTO1KiAd7/XNE0lzYkvTy7tBV
vAmRKb6U9cdXOFgBkSZnSR0su4gdHALofD/a4mqSlVzJXu8qQhQwTZ3yyj9xNxhTvj9CnzAsS3dH
gkBTCFSthQ6jjxnqQveozaeWpseG7snv6BxVBpGTzRayo+Hpc0nAJ/H6B0Q4pTKTKWcu/b7ZCWvE
mEeChnPD5UJ4xbbmH9iZP83M6zAmRCB2Iip0zAOSXQWxou9jvCw2oC0oPLLJ7oUDMbVxU314fi/H
Q7O5WOXyaYv+5KgqPsDr4tiWm9LFR428g5iIRMdtoNHCSEhr1rASm5znoBxe00Twa8ot9S6Zh9O7
cCVn4pSbI4mDtMwmYiZJG9pyuFHlNzsloVviSFdZe/ht5zuolD25/sBX6RXTtrcWolfhAp24nDwP
eTr8i19LMiFvY/uMC8MsP/nUkt29AfBOeae/+j6uMnx6FQqd8bHAu8Ms3IrLJkQgBgvj14aF1Kkz
Z4wAYJuHfiIkFsV/igZFMVqZunvDwHEKZNPSBZkdmiAdLHne7AnYTk8zx7J/7tQSCgMIONkcSe6z
8M1j0xQx5YgQr9jmZy3SaY5sRYwBxrr1NXr2B8Zk0nheozV2+Zyv2V9tarKac+RmjfxkfTAuyT8z
+QehB7fTnAyeR7KW5vXNcY6EpL9ZCKHYj10xbtkXdmdIsnAuV4B6O85kwd7eIzSehBhS+iOYytfr
IDIi49JRQY/WLNMaYrNe1q4i7dJBLabR+unsEZPVpV1bC0yk1HPuLiSBazvPyfRNLFU4U6y80gxc
PerEVKTDdWxXdmW8JNYRsUXHxRYiITpHccbCr7vYp0ym67b5+K2o/j5A3HbgLZRyV9v6ElWYKsNx
VcHfx0TABa7VYVKKbdeBpeokDLJ14TAYR4Dp+Ixk+QyrC4hE6oiiHIg29BgGt11AwoSUGyyM2VPF
Td9et8gr4pgk3urHpB29w+Usxhk9cZOyHqwu733fWHFJh4MO1Bk4sTAbuUi6+TxT/1f8UUiFjpgD
vJWdnJPWLX1PrtiCI14AfeN3W5v/fnrbHZ8WqMTDQX3trkEz2Uerjl6JjdrXu/HTFsw4ZhNl6EyT
PlZBf1bGInkAmhJjQvzVammkp7zdlHXQcYBZDRu+lAkIrPYHJsvRS3eMo9/HudbNoJQMkUIr5lFU
O71SIbr1UtVCpmTKyZI2qLGogQT/SSqh50yE6t0YMCnnlZZVE5YOPi269aCQbb/oz58DilSkEF+3
SofrlbvVw//iZKQWf+rObticDQnBFb4vl1wL91Wx8kEoVDxMxxnV/G183TZ62N76g7zaxILLKK21
+lLZYzwExUXZarySIrC1VBA//z/0CrweyUFyz/vXjOCu8tCb0pxF8dvgGwe1kEwH+YZw4UO+yePq
qqk7v1+3YzDOSl2Dvr9+Ci9Rn9eW8dqlfcJhhKdHx9L8TEF48n373mw0sLx19SskSotFgQvSot6g
ylzsKxwswu1YjXT5qt9X0615HMBSLpi599fpLEL+7OLHp1+oQPtFLQ60xdy4xM3KAHv+KYy87He7
tWkO4Vk1jou0GnP652KJKMuO4/y1xvTU3OiFlRhlHhm2fljEpZ/ZuYk3bzmR5YQtHyVIQef8unMb
h9KyHtfxKTVr4+mpb3URxYzfLOuRg+UGuinNlgaTGEdwX5MBbBRxpoRg6Zch00Eupq649KrVKZSd
mg3ztAA47p0IogpSAijGtS8fsVrblPL/Qe2iRG6yl0T1U91Fiwp1NJEZ4MND36uhKQT0xIiprzmr
xncXqTUgASlcpFjubj67v6sRiBC2pu6e1tggYadVqyUhnKb1DmDHjfjEFgmTGWWQhlWbNRAVMRu2
HlTe5x79ToshKxQQkTInAmYeAsJ8xDrV5RSuEdCc2Micnpaole5VKYwTJp8LwnxVjHBejABMc4aT
EBdE4SDp17HdJjti6furxncI3jymLeLfniSJubE2ICba3FmDywPuvZ42yXM33QEwSDQAZhiYIsn9
XjL7GbwTEdChpfI/ZpPg0bzd1leOpYSb7i1txjVdCzqSYGcU1lN+bJwhtQfN8WDusfYbGCVUPEj+
zVcIhY9R/2/2G5EI8pTz+tl8DS8V2ZcvTunkMu+3tDg2PRwSo+aX8NlIw1DtTotr9Cl/GpYOo5XJ
zIpT7WSI8XAAh81CBsMVswB41mRg7KEbYZNDDldUHFg36nrVC1HwF3WLaEbCTfe8wRz6mB95evcH
SIUM5/q89rpDr4Gi3knDQ5OYB3jB8+VLHCv5jkYHG9kanG2UnAEU339t/DrsBpc0L+9ceiXKS56f
DXHIddL3CiBmJtKYTFpdFwPRFifkaATLPHIYb35dGQNEgXfca+Voiq5pPCelRW7Ut215v9OtqSFj
zY9gBHGjyTDChTM2AFybupPTKdqhuGVvl/Bnbd8ezJiLTqTQDFYYVBAEOfQ1Jm+l27B42QGIUb2m
FUrm5a7LDC/+c9AoY4A3V5NvUS7ljXvo4GeHlPu6xzCC6TZ4F6cRpJj5K7TwXWJQWpaZFpt3wGC1
GzBBJbJUihzS622evNf9uTqFqWHYKejLOxISDEa4Zeb1QtucZI5u6aCHoVodXxCt52OUtWtYKa5b
5PLyyepP88hITW8F4oEOUx5A0fcBLUUOpdXitpKFuekYop1dqTltkAc80gP9MTwfLrqfxhwC9Ypg
5TYBejlHLWsiE1M0OeWIBf+vbdt/TBQ7Ob7GmBIaID1LOry6Z+fn5KMWya8jy68yqUDZ1SYYNono
Al6Clnst45H/sgFwXmA+PFBgqudeM8Q8rHz7NCJowEHvEGEfSRNenvfNfiVyvsnHqvSfHN2pdU9a
Jp5tPDOIZEaT1GhDqf7Z3SfW75rSWsjNHOmOaWFS1Cd/pZ5j71b2Ia4zcNlk+4N48SZLHps0eZjB
ugcUqPjcl92pa8b3GgnS2exap5j5v58nSSwChY/7/cYrlV2u/+5yA/bExN6QiO6qIpoiDeHKFjNW
sdj0CUjR6zr//Xojva7BRBhc22EfQ1NW4qY4dxhh6hIAmzGAT9j0HJ2P8vEVk62b3Rruq7RZqa1+
VAs0cpzRCUQaXHQ41d8F3fxQ2nih95CAIJBZ7Cu0BxuHBbdQIm9Mb7sHwDugEIqUOgnE8itS6hgG
/kImHx5KSX+YGkMl45ia5dXXVFXcFoJJ0DmWoWScV3tmKFmNm10MCJsaXnQ3SiWEqzzoUZURJSLL
LKzsio8rD+Ik61v4xEJa1KLh+1sMeR6wSj3Z7S8FGywmErVsgzJy6xIg589TWYuQxr8npeAPidO6
osSHNbxeKZuS/yL8Uej/Vxnh1EIbE8AjSlP1VGQMlS+DfRJaY8IyDIUOvDq++Uzer7tcLyO8MvMi
abGpoV8cTI/v8+4zJ8GESyLWECscUDr2t11kq8Eu5szdsGRdjgPahNqysGU6ihIUJCD7MfFAr6nn
7GVXlqRs2mrQqUi1bFFbkKgc3emPUCYUdbMYvBYvYhZIqa6Hi5TtB7u1+ih3K7ZPf6Q3B7q1Qq5d
NzR2da1LGEy+5cPJvjEpjkI1zZriGOvgBKMrpa1xM3iW7bdM+lBsK8pQK4pmohEiUQ50y8ql3Dzj
kVWIPNnliV/8a6PTOvR6X/4GICv09CLmRaBcACP/lwDE9hSKN/WaM9KdlLZfxs2mdUpyre9xItez
spRzQUny+P0wgHvB/v2N3/WYD2p+RMJVpPAeDub5FWd/p6VAg7Z2W2ivpgaC8TQbDWb4HXw27cYz
u/lYKjzv+ZNAzFLSud/GhhB7zMdNuAVf1AXu8xMq71WCb7L0WJ0Xn0uEOnwdbuyKAmGoJjUyyQnJ
c2+MZihgAQovh5WoBCDNTz/vnlpLA2XSBLq3BqEaftWLjazcQpwILMqYmIzNbjdnlxnmCpJmeBaS
Ea3kaGF1nzuPaHMKO1mp42zgZUe4p5noplN6lCtvd5y39pUx1luarpD1uLVpYwsaLzAGFfrGLrax
Wfy/gMYfVOfyNFz6whyjpiZjx/TAgO0HxI4mf+H81ViDds3Z/I7rlHuG9lnJU5k6eYOglt9V7O6J
Aje5DcjDPmx/aH3uEtIBubjPd17I8OD3IXQRXfQje7NLWBYTJU4Blrag5YUjqdS0G3lcjZ92LZN4
Li0CrvcTd1DN2zUWaidlz7MqIQ91RLSn+OVbptOOnj4wQayVsglskVtmIucSbMjIIYf+ULf2cnFG
RSIZYwKKhh+upiCiYC2nR6YWsrj4iMaLR9eFeaIdsSoaDdICcrEyrIUAhM7rUmtlnvJrpdm8bPcc
hgTcw6fR9hfkAClgQvAWKGukS0IPsCIb5pokWGAsiDNibF4Ef5e9APEbTf0TrLeIp/Ndv4zTk+Lm
TrKCpK4EFSszgZjXWL46sP6SXcOQf6ja8Xb+4WkbfkQcy6XU351rwGbmKvRc0lidOCj1wnhcGTlF
a9RPwWXEfE0nfZXYn1JOLqCCxT52o+f0NZk2E2ZAw0d9ZkuBsLlh+exjcbv4KJGfARnpXeomkzEY
sVTluvwSOhrz20dVD/K28dfUPinM4fZ/Pt4UR3O0xmBiCV6oxX9TVQTzIuFoRuDz2SbwlX4OF45a
T6F4+FswSvcK1CvFXB3hhiZ6wj02pKcqW6qkmtz/WyWQSmDzmm1o2AZq+0AZaVIlW1HWNcHMVPhS
f9ckLVFPk0UguGqjpaVmeEaF1if4LqoLw9V0oeAtjCTZpI1MiyS2yid/Y98WuS07lZDeI3dSnke9
f6U67tM5c0NEP2ntJDQ1ta8r+VlSbB5/6cvkZWgRFAu81zwRYYAOuffI57VxvgjDTwb5bttYtFVd
5uVMJF1VqOApT7wwuTX6qskAich1mxSHqnX6FwSBEpDWUQQLzNLCoIXbOoYc+Se1G0Rh70BwOHCn
dRs6E09JDsmZQMUzFyABaDjLVaGN6vixhdaj57MjMxywsXPhf8jVmXwqbB1pqNgg5p4RCEItbbK4
SLX42pNeCl0lOVeCrVl/I5ij1D5nzaj9qrz2lBruhW2Ow7wdNyjq0124IwM7mqmPLl6h39D140dE
GeevrOfmivNaWjxvkOVqEF2l08OJbswQ6qPvQLYIim6jIgG1CNTzS4JEqW0Vm6HpP52XjqdXGwKp
vNq3OEmfk65fxU2R1oLQT3NEDi5G5GIYVHvH+XdLDkhal6NNbr6TsDPDQ4GjlJknRQ0C87N/RpqZ
mTC382EZ8mqHT/UHsittag4mGeSltxzHZ+NSKGYYa3FZlmnEKrd0jRgw+94WdxPizH3U8I9Rsbwy
zvV682QFjmRo02yxQBY+59p0X+0xjuxFFX3ZCWrLhWGZrtDTo/+H20dxu3zbMcrstEaED8KTzCi3
T4YI7PwvG0p3TOFYHmfy/FYchawY+vOZTqCy+HJ/f3Q+QSJnSVHJIilg6RMJjJ25mEX9d0/MqIZz
7daHM9aZjRauamNuQgEa6+npgJ3t9eFgke7as4WZa5UKP5jb7jVbtUCdcbHxaA48D5KcJVdDwSrx
DIU02kEOyw48z/XnSHMLYf4Q2pAXyfEIWWiGSir0qmlbVBWWnssXp81bZ1P1+eFVKIssQWhqYu3X
9qVIaJ6kenXnaBCTq4qHVXaH39V9ijRXgX6/Y5lWwWCAQdO571OW0vFgKWi9XrqrMvFRunsBG66c
ETB6E+yU6ijGZsIM3iEJvb70QS7NJkP/ybve9J7cPfYqDRcnstHoUbhAJQcoDpokKgdGFjNvq3VL
efB7p4u2BTluKGsAH33V2SP0UdxDUX2HPWhyGLWC3U62F+qSLPn8+Ytqb4HeVC/mBI9dkToRagZ0
q6IO7JzicwB4IGP/S8qexaaa1dKOvm7RUx/UFId7QdMIK+zO4yuFET97MR3KScNxQAicXelqF7iD
ZKVr/Lcm578Pxx0qzy0Czz6l/V05fHLSzvAMcWSE9/lA14ueUDtlXEZb9YfaJMB5CENU6b0MwYwK
s65h9EWLrXbsGknA0ytibVDOpsRmifJVVhhxzXz2XsXzvcEGt4cLELUlQ4uGcGKdsHZihALAoZ7X
cwaw3tyBd64E56vbuMrjvl/abTsH9mhi1NLMvi7b+3v5YKEV26YW8GQDdf2BPv/0WmYh1SvAa3ge
ltZt2dUNkLps0Eb8ji33EmX7ocbHb0YvCXjUzhZoaeozSCGHWUWeqzz7NMUsYfRUnId6Z9ZteYJN
KIuyJloeZ67lPdQYEl6qpL/yocEc9C0489W/UgolhKJPJUYaqB4Kws4LES9R2B2SZrf537q69vyX
ENsGJa0P7pBUNDrahxUDpo2xD4GhfboK84AarptKt3LbW8poSZxL3FMRzxVFTuad/YeQoHnhgC8g
A4FZG8kn2fj59ACsOriHTJ+khaGlc8AJGXH9+H11qlSoCsvZLW4kICNAvrPvawVKbmW/d1/b976f
xPN4BGwYE0eX9Xk3TpHsOTt4Vr1zKhlTsW0EhYgmuIUomAn66N3uOP6aq8UQyaMY8Zr4K1tAFWm8
PvbwV90aHgZUm9+fuWCpCJuL/6mmbICCDopTKJlIGaDE0y04a6GIbyWC0u1lXHJwHNZ+OWZvPINX
hEp/Wt63OmCOtiVzrULz7blNZFbPwTErMbCxGsD5xwqKMCZYCbYtQBXqnn3eSw6Qu6rZ/TAZ/ZfE
6cQewxRb4RxIhFa8UpeF4nKp8L7cQircWkphkLHTOM82WEoWUOMLwXDQ962/61uj48M8ujdZUBJ2
T2hAtUoUquOWrtAtEecCyDYUz4G3zxjVkYyNw/IWrZvhpcKMNJ0mTjkvZ5FvAaJS25IRItIVD3CA
PPdLpB33z2XQ/v5T74rwJnNPLH+aLXAd5FvNJGCmb4VfSbjAJW9b6uaPS44eICSWuN6EqVl+m7o+
lKMRiwYi9W5a+IZaywq2AG1h2y5LECYuJ1sWmZgQ+yzEVvZg/hMgtcUTZfDLhjgnE6CkX1eChVSG
IFQnPoYfyzUsZ4mBR6RCOBhIhWJFlJulx4glH42K1T2KaGbq6S0TUui7atdGZYj4X0hnN0+fXXDM
w4rsaY64t3WdVUBjzV18ASBPCSN2vJhIA7NOlGZEcTWyo8YvrfV1aL5TFGQZd+N2s3oVx74c8TNR
bvEj63roWgfFO6nwmtn8VyUC41PGClMj5aDxWZousiTMBcgNoMjE92grNYIRflpODRWqoI5/C2An
iaVMFcislKrrtN6vozW+hMknmUmTKzFxrl8Ij9uJvaUA+n+JheY/+gxKRuMBNlYppOtTZ6aon6EW
ayIBvW+rbLFdsZeC8enAbGhymSYB05a6jvWMdAbTo7mDtT1heP2PVmFC5rJ9g6v5jHltbmVV4Ihm
l/L5X5LGcsPDDIKVvABvPJnDv6hmaoSQzXuGtZbR7IXY8MkUZLOSoBOqnnZAQEearcQkEpMCNi+q
sRsC3uchjUuvz3OQ8QcLTr679xuQZ7ZB0lkHTYpO8qfduYjAvTqc9A/4YNeU9DqmfZyU1pElchMj
vWuENrBDoSZw+E1fFbHdy5E9CeK5Au/EL5DsFtLPXz14vHFWEeFWjU+ytpoY5n8t1aTT7A1acpfO
Cw6Ea4Xu/cR6RvQY4fPXG6WhywSQk2wXfHVfhVJtJgIfT5/eZTf5F/ya1hjW1FQYn5CSC2Gh4Oz1
CDYKWLwAocVNPyJIkei0PAnb2X4zWWKlFRYrS6NQdvGSmdTE8ajTl9uUFuLEDKkezoRwqDM8F+O1
oVGb1NJFAXTrOVC3bk3hu0PAIpYEcOcWGB+/wFzlUKrjDhosIOhk+s7h0BgYbQdg3/0EJaQh163/
ShqXDanElJEsTc6dEnrq1E4N1nKNJbPkq/bsvBp+Sr7g5Jd1CkGwMcIelaleGLbwRHLeJ80+I1XF
H33lPtPy3jIYkjG9TH4hMtvIrzOIle/jV99I0dcL3QyjcFIqXQoBwz7sJMFSamEieAfz4yHq58Ul
XiV8Am17GOsjHeYdSk3xiPJQwMisehz9HLBMigG/hYQzUo4rlEpzp9DjTESJ+rmenh/kKjaT2yIu
6XQEJ4BtO0o6q4wsm7HVB13JisQZLK+5uQVXR3QjS2eoB2gh3MgswVk6wZg0PcmbPUrsB8zalO9b
7iavfpQOYpSQ9P3VCkD7JaDAx/zMpwn17Lf0NoSm64Q0tbhbLg8DQmG1oNP5Vi4f1Mh5k2m/DFh8
aPzLTk2duOn+lQahTfBsIOXyAiaAvD1M+/Yx1Pl2rqrLBnySWdw2HPRKFw3oFFVWDRVt/2w9gra8
QQOnTVh4H/iy77rdQ+jYkFbjzHL0zm0vcQzyDKaTutiemvNQ6X5bNoFTe2OtqWFIE/ZjTo3uOfDj
o0yrXdWkGO6s1UsXKHHC9BqxDw3FymmX8foPj4nxDpWjmRuGI6ubH0YY3KETbaqSNTcZvanKtotb
QC4PpRJN1TE7IQdItrsAkfn6JVV+LKJ9NYym5+UWjxERYRyCA3GK6sZ/Ge7lED+NVgqzcNA+wDHL
4YgyFqEb3D2RzHLGKWaK/oa1XGcaHSdeph7Xa99L4Yc4lsB//oJ0ql2OkU7/1qYYh7MqNBXmx97A
CAxPwVQ9oAm66OdIRx1KTVXUkiVlqjMAj2LwqbUTnvNiClwhFHB6OTBBFqMAEVIkVMp/lhCRWrQY
akJP/xQHsUEkpkiYRkVBKvgbCTQ+tcclY7G0zco69c0E7HRckK+k4TsjdHB9EuHIlgJOo06/TDrx
WQ2G+CuXXt0gAikmQ4Qcsz/JyPWke/HuntLHdSIsPlTWXGnmh9axjhjAV5cYSOt9BBnbsUIsnDVv
9OThZCZuW0ddpmEvd4yASmrQ+liIP8VHP1JBXLsjqpJVWpeDvH6V1ot8ySq0T94V6XuENRfWa6nk
yUwdG+bBITGH4h1F4icxKvOCnIHzizLr6sKwK4I29gSoIYUeMIXhkZKE2zgFDtyboBDi8E688pJd
2m3+or05nCRqdIG/y4ifWUeeetH2ztZnURvybf56bfkZLz/fsQfLPiHLAySGich5iMbxfYOemADk
CqVHJbWVC0E+eUcJVMcbGd0xkXaBUD/OQRRGi/SG/hpQAzTQ9YlJpRpfFH6KQZxyd5CWCjrZhzPw
h0ONh+SLScz0DWHvOD33Vlqufa9M58EBCoIx7cyxQ9AjgemGGP3IQfSxB73f0HMnyJU6LeUSRlPc
W6TfPZxLYOOfo+eil75kVo5SzFFwBcWNtb563DsOnM3oPYIQKQ2d+odAwy9aTZOjGXowRGjWlw23
7pMeaeVp6y2gKSXwJma55ugL/C5fMkzqMc4mYEpd2xUxtD52C7TRSEjjynfX2e5vcSGBUbP6bxeX
Q/wlfpNXvqKwY+HhzquW7hdbXKxNQweqRgrbUuLYDXJRWTScsbx9mWBBpnDW0m5Xdk2/yrGd3BAY
MCTrplLEBoC8YGjdJmrjkpeKeLwoU+39DGh328Tpto3WR7aPKKd+a6SmJBJ8kmyF4tfsWt6Rp4ru
QLxWZfbLzUoJwJIENmOSjcA3+B4v72nru0sv6HMQV4RCfUhfxbK1CMNB0aWcDFBiWdgmYkQYcgVi
AyvU+eDWBu+OrqULgOFYZKltwclR8xUphz3gTvS/0ZB+Jb/lfrkJ2mEHZ4oIOdXaC4mkxRenZm6y
73c+D8Ln887lKzcZA0qRE/BwPc4cVMppvMbQbQes5/SU0SkmMeDthDDfsBjnYZlY84PhxHleqqXl
GdGh9rra3UFeYcrAB4D9uSq8+/HlGORknOZTalMiT4AXMoWMdCbxd0uSdnO7k9uTpwTB9KqRGRha
gwwsluaNY5et2bQtmvJFWwRB1FduP2HU75JcB36lWvY2idEuxLp1OjrTMtQiOhm+JK9pXvhLutkW
RJ6XiqfOfQa4a9gh5atz4jgrp8fS+HC8WeROMAXIWqsmswnj7i29neb4rC5Xat+7G0KzRKWyN//N
l96HocsGEeMcYcoTLefvS2T0LazKPspm1nyRQguroPJHBp4XkEcnJ21KSh6UJFLwzsfnZ6qWbkJl
zpazOUs9ncb2T4Wln7WZiRJidu2YvDCUh0NQUZOAoHeDPPDG3mq1Idg+fuixbgVgEUbjZVrscATJ
6Z1Jh0Dr6b57ssXs50jxkwUaFcIIgSMjrplWr/2TDFJpmEZUErmAkfRTj8U1IWweUhqNWx1vCMzg
d0uQvwP3xkl7o5dzmqGYogooWf7tcJAlD8NZFT6Kpp6ZJqVmgshGr4FZlQbY+qzuoosFZGvT2qCP
/iiuoOst7f2FwO+nY5+u3L/FyFxSRiEoby9xixUAJWajfMzyiGw1w5f27thnJz68kvKRs6sXoaej
84Pmgv9I7dGcsSjBdhfqVpTIATSCIRtt5gsvqOBPQ8bZUE/q+Zei/WQU0sCfjHHcXMG9P2+V6HdT
5ly0MTswdSlFtHl3/yjwzaVvuQvcMmlamYFKCXyKRbx3w6y7QYeINbpIVE9zew1hPp41mN0A62Pg
xHXgDsB/YgdVUdOtRzf4VOzifNjcNIH48BGeTOkc1GVP4ItJIwGHfmk/aOgtyKkhzg8tU5uMXZgD
tmKcfMeX8uyKdyUgdC7HY5UBU7RW29/Yk6ShMWbw46f3xIOYbVw2nkm7jeNt18HEyvqD1wei7j+Z
FHZiAUahsxHT22BQor4H7L0rzsZKbyPj4prFjBhS2GlxE8pKoAry8s7rJrOfYYiE84iEARRoBFus
dDkptMhZj++ncydmCN71ec+yPuodjdI0Jjak5PzMpAYjulu49WSvUEOYyug/nhwPVLelDGvNFQHZ
kROQogmVo1UjWHrUOQr73vxz2bdYRqc3zSp+iVXyo7rg977YH1jFYoeEUaKaFhMN58+OfWdLK58l
gYEy12hpq4pP8u+62sA+nRqsqpbSo9nzyZi6U6JF3Uy/Euv5WjnS3hdVAXkNixPSZgJj4QV6v4Uo
lHqBb6b9P/tUtS6AJQ1wiEVqX6IcamDp1YuEqCJbHvSAaX86KZGqZQ3fYg7bgwJqAaLo7HEdTh5c
5iQ9i5mpdK7zTlLaMAFA4bnaT9BEP8Bt2T3XWa4O1XvW3b82vENfSg6k5d9S5SszcYk1pTmA39WI
EBfdjwpwUGrLgdBM+C94ghhRdNmtHqkMrR+npzrsHWLqkg+YN1nSiZQVVKcd+6rip2Q3oJ3aZmig
v74Q18Qm8f0m8dpENKZ6vQnj8ZXXE4115HBC7ZDU9FYcAb61uprmkmT+BJf3mLKIBuwlVssYwtki
hCpNuxoebOSpur0T5npMd98qNoQJ/pjfbE3JuRH6DtiLvdvoQPvlDHzI4mTRLM8DZws6K5yChK09
6YHJZEx1lMU10sbLdD+2qxbkZjvKJGItdjczXQ5Y4Ddh3lVx0/t+oeIvAm97QOWV/dBA716pFHq0
u0f9KsPvze1FJb2hhmgSgdY2BInpDdkrKKavvVWAucJKNb8zhpuhmivcgkLlneH1ujZY7DNIZk59
DY9saTNKKNjG/tmJitCHL0HsM54RxGtpfBbo5PuxIPCJDzKn1rzukxrzDf3tKcPoQ5ANmjZSk7VV
mcZ+ORlB4H5zjbzAmUjSnfkSKiD6w0BYVtQgLEbwXpY9AB5ulM3a8+WJz8MD/y5SoTiQJW9eepfP
n+mMX98JZSZsRIaRDr+L9PjJSVRrUr90DKOZNKxKxJUFwO4rOi7dByDBNzbv7zqJTYrvgn+ZnVEC
4Wz3gkbosmBS19XkyL+ReDMuozf7aAhgsZpbAeNU38Y0UbVYZtMxZdJveV/VJk0d2qDAiA6DW2NJ
JWo55XlWm5Mb+Ft7l7FqRbjL4dOwwxP5Ry04vnox3L/fPuzuLDefBJua6sNmw2v+UKU2VFFySeE+
gNLoCDfaj9dwXNQVsR53qUh4w+68xmvnWF6qiNFhuO5lQQVizhsFvYw8LK0GvyuqQ2Ot9sDNYk9q
KMUwpf/wmLmKN8pm40vsIfTa9LbZzNTO20PRNyXOF+u01axPzRv1pJm+gGe7uoBNSiYzq3WZh9Tg
3fPpnjCuorSFKWpWvDkhafNrU8HxxhglUUEtfezvToZS3F26owiiZXiUWizxRxcIY74bEocAD/5g
z9ZizDLuj9FzmIScxniUiBryHVhQnE5lqaiBdQC9NT/7NGfS2g6fZizeHurO/XwG4Z/1XCSiv5HR
HVx8llOLmJFQuaBGPDRKkbVMaq2dfKBaZJ2LS1ozbv97eXbp+8l7F9aP6Sz3Raoi2bw/OXgSg9is
Vt6B1lngb3ZoXZyjT0pTC90lE7nTt06SYQsgRA/qxlyWMQoZvsGwtP/80ThMWMVaMRV2NWZwd+Ej
0LWcvR2jyZdUbEJ1DsMxq12aXPeAkQ7lgetDRHBORBt8A8cwllYq0bbxeDmIMxqjfaOq72z2SVLT
ZpHX0V9wnJvNjZQY64UFek2bKZMOkyu0aBj6JS5C/DyxTBVEzncv02eABzKGj1PDsHZE/AmpsUtV
SQhL2BdrGkFyR+6XCP7un8QdIsFxn4S8D/DSoc1gxxJ6PsmOOSA8wTuralG32Rs5mkSxRTWlQMW+
AeExI30haxDmm7Ojv1rtl2wMIJ+Kbe7R5sqXHpFd94w1BERtoY2ynyXoL0LzNpxccbPQB0608MxI
H2SOsMPmzgZnX5hLkS7YQbFp9j9hSaDr6edjUVb8GqNIALrz2LU6poj4/njkWGCLykMiX//PF6ob
S+GOAy+8JZoq5q/alFEX+HnvR3+AXq8Ua2OnBxoE7EH+D/M5StF6mRshtlLyBGXwEyIQrviItNbi
1ju+faDX5JCfIHvkBxMO0086ueVuds5gp25fXxqTbk2uICYpUp79aVw8ocu3WU87x9Hv0ydFdMTP
esAwyc/wD2e7ugJrohokZGCf30zYFegXa1dRx4+vQyt13Xl9GcPgSC8jbah/qPr/x6n0XfxFLUOH
5lxWnYJbePupKpZv4tWdaxoh6BLZlnHf++2wcgk2+SJYcjQ964GcJK837zBFdUmysdBsfSnIH4t8
iDf2bai7wB5wuD0siRAxexMnpx4va4n/rNfmo/rZhARo3+u/O0fJKyb5ps6ziA3Iu6G/SmiMCtom
iwpUwb5pVh6i+N3S86j6Wb124BWzHY54ssr2EotetqNMk0cIQ/nBzi15wU/kjpAbusbExqQro8IX
17WyFxydCpai6IWjwUdYwauIKQdVWaUUhvUnJOSaRogbFca9N9hbaq8Lv0c5bAhxHCkENSop/J8X
pUtTUPq9ajpWmbxpfVjJhvalwm4RbWhOtk+r2zS+MHkUJ+djNTkjSLOJgeZXJAh1d66RMGNex1P0
FPtQ8bmXRQ9IBDytmp3WAC0DzYmsd7uZCk5I2Yc1cI7ZNEJeJedWnHyVZ6xBe4S/+5psSFKVLg+u
3g4eyeKFq0qVCd8borcoURqBJC6d+E39jQM9qnqikSL5pCECODre8O4xhhMqS6xz/0cVvRptLj41
Do0s+vZ90qBVc99cWpFA9klVv/ssbZ0ovfLyRImrYlR9s7I2lNVZ3izGKB6mgpBGWKtK7ZAIbUDD
wLnkWv5EzWo5jRt081CuG9miE78FEcK4u5F2DBiaJUHB+kEfLYk+GyvTBhqO6sVAqhFyqQSrVszU
sAgC5+E5Ekr+vB1MxMARGjgipFa5RoS0YvQyM5adTKIS0S0pF4YUCGLG+lLtPyRmWDLaR1qWnu9h
WEHO1MY5OqcT2V9lXN/9mwuurjRVL5Jtej7iZTQR0trxtNd7Q9N5WXVdurlOp4u/46L9AhcMeIRj
NEfTaA8rj744qog0VWi17iVHlPYkrUDmbFttJDZaHKP9N8IvSM3HNNKwcB/3ScbfY3Xmj7UjO3r3
a6XENFNNqsqEn33ZCqjNiL7yYN1m2Qdvj/Re6irsc4W2IQg2R/HOc5zlIssffPh7oMoBsCBdVWPg
pN7iFT69PEN3mwrmeJL5tK7V7/Xga1WPPllX2dhIqg7GzBauw8mMxkl03V6f12hMO2fEEyZ0BzCr
k9eZG8HN+OccYFTvKmIdgwONkhgfMXIwE4Lo3JZqT1vHd69gnzbiwFwqujSwu9zRuq1KyOg1mS92
DHY9LZXJYzb8hijhqZR048nKrU3TudOdcJUmjBmeJyy7sEGICQ9+RToRFf0RiLYS5oVM9UaGvw7i
EzuVoPED2yHG/3J27eFyQBW5GWjoYjAlfZ61eXs3U+RDAdcQRPLkNjU6HyyE4M2g7ltw6X7VffPX
LZpXzLF+c7myitxe3Ke2w7MTgKuNm/ifgYGmrszfuhv+BzqKCgO+92z20bfIsWKJHpkISlfiyA/w
prN283LJADFu4NMo/fH0lfgcXpQ+Y/8wxT+y2qWgInUvDsKly/JFC/yiSnz39KwMUhfrURPeE4Uf
C11Vr9saNoyk/yQkKznykNNaGqCZp+jrBNFPsfxp3KxdCaK4vepR4quI3Q5EKjnRInaoISWcTcpv
Prr1dWHB8pSjchlGw47sIiE8qxXNl2jXfEZWXWcKnx01Z7OpQprNGtshxc7iLjARYslbXC7gx8Hc
vqIj5vrf1COm4bN3WKJa7M772jYY5UZcLBQnZsWO/+bCKL94b+7v96SmzBxWsbwWBhhOiqalAmMQ
mpivElQVY8sOgvn9iHKVOVXgrjgfLsUUTtDD//3kcQcwdnQIZpHN2tHsN8331rue/xQkNbKNbc/y
PhK/gHHP2KBgLYgCvmag7u+F1NM8zfjT84bkIYtkWQF0KP9Qv/iv5wCULrTQ1/8inbXn3Q0y0iNk
EHnXjx0eNhx9ad0gtl5ttnqOR0rIF23Tl9u/z3diUg9nUPg3kg0b+2229e/RK5KpgweU5lBl9s7l
eBTtoxP8xYEznldgSnZRK/ZEp/rd4M2HcqllUJ0I7PwJmkH25F2Dg0K2DVt+QfJ0P6a1YvI0R79g
pu/slHAXrAHMy6eHwezM9w4IxcH/11wHQuHKuxdqZR3eCockVBMaKXrYPtAxt6db9ebsbbsBaR58
YXe+mfZPfEDBKAGxJVtlPyXlzuZWjx/kMEPzjXk5YMBGbtfBMjcocx8Q8/Sn+/uXYQWyuLvB4/gu
J5Ubds1TfN2V5Fs15oPHRTG9RC0bAeXTeqkhQG0eh2r6b7g74qs5EGp308rVxPn9jnvFLwfk6iDj
n/csoZaaFJUo1f0nGoKESWwX4ehjrtKJhhPJhdeSKFB9FdDvHMV0sPp8VslU7DXDcp/Ap/ebXHRp
EH/J2GAO2qbz+ysyVmrxsy60v5HJ9ar3X5WuC449l9G1Ut9UPEuojdZddC7Sm+NOTcfIeIzuLpSR
hi+8mbIU9nDhniqotlj+fkNO+wnK/1YE5d578ywbWHI9DlQcPFkYybPmsTH16MEdYzt/bzDBZ6gs
Ad17mVxc2jG7fHoY2aIjoXjSmuChP1juk3Lu2tgV92ldCjWn1U6WIxj6WvwsTvuFYY1a0PGL8soR
lPEuBRDLZoDja+YcxhbNs8HgRn5GZOTkBeR0PDRgubkBgbymrI+z9K+hu5nCFhnfKPiZjyhTo02w
QpzA1OADmxtl+DcmuHpzCEGQgzdwqlpAtdqUrVjOZ9zmEIoJd92nwOaF7qcHEfiL76izLRHgi2pz
7Bv3M3s4Mnlg/DR9owAPjpHreqFjcCipowtU/gLnD+mQf58tfcA3JguP+D53I6kbUDQmkJDAmgZ/
Td44iQhAeJPxt4CdDlvoO83eODfPRz4TgLR9VYbkGiPhMUfiO794p8X20vbeonhw4exxJexUg17R
HYx5GwezN7WWgsRE16a17cMPZJTNsqdYfHq74LjCcPDHb0TPmVTlltIeTlE99MVeVSZYFA1vNSJg
WruqqPHAZv97X069/rbr/A3rexybsUFjW5FPBCVSxB5QJYRcS4TNWCDnzkAolqQT5hugUACaXaWj
PEOjqKkKznM14lo3nzJfdvhqiuf3qtiOEsisssKWuWHPCnp1xvwoazZxCPxIyZ8pk5RFkM0+XSVl
omfBzF+Uqb1oTJDzehy3a6p1x2HpivDEOQv0uPgJP69aJcbS2u12w5aSXs3N02W1el+waIoC/st3
ZH6wo50JrwzAf6Mysyhib+HTo/caCTWDBbPqStP3d6iSYG+7GA3EwhrYDihgK1BinhilpVcQ+kL0
ja1eg/mGv6PG1Ks4eHxkWMzdmxuUhigESFff4R1xx8g0NFrFc04KUVbsXQV8Du06ZZkubwXAJ9VY
hnTgdEosGSvs7vqHPAxOt4mA9V3WNrntTXi/kewpJvBfIDfPhEvIE5X48fB1qnOIl1HjECn4yKxn
n3daN1MsM2lKRZppKEflDi7mOo58bOb+y53k9Kn+3MBKg486EzabFtha7dyvdEGUJHdSqF6UWlNg
ubns4JIDA6GfGtqlA0aW6TMhPG8ZUNBqhYfxI8fL444OySN1+4NggLby+DHqchX4wsC4xeOuv0dK
YCUB118AmXn9Z7MyUUZdMkkDxRFzgn3p1rk3nsL4ub4zwYpGhWoytpKMH2o9kVn8tWa8IkG8+4QM
j6lfS/nG1Yfy0mAwTCjb4HWfM6ToHDUmzw2v3nNdsWxY7h8Sc2lrr12rUvTjN1lbQ2cM4O1MUwJn
K64A+uWJFFV7owenEurmvqHsYrHScvbCPNekJ0qZLc72agDp89QAnjC45qcxlRVS6fBwC0QggOLT
JxNMaSXEb2ClzetfYs1j3o9LFZ6dGlVIK1iHnFbLhk7C7yJYU0ZA+kr0SQQL69hzViB4Zr85wEsn
sYNxES5DlofZt8Kf78xdbR9Ux2fn5C6qpz2yjNb4IaIXzbADKBlzcI8cHOOavfk+KQJzjdtm4U/Q
veSdJGDuMNIA9eNrK+VAN3MM9xN5WvotcjvlwHM7JEEAKVqTdZLhXK9IG0f7sFbrVnyoQYrvq8aC
GtYN0Esc0ULNm4SxhMX28LIHbqq+Fq7BL75vmjx8kbe3iFANGrAXGuKyI6UtH61ZaxaS70SMxhQv
IFcjBiyjSBEpCdelZuymNXDTTFrzva3K8F5bN9Il8471AVNTnAqHctNsFiRA1UNdbdZ6zyKwlJ+K
CjaVFThQ30YJL8uRBh9bW00zQ4BqkH2ip5WvV/phvmMrN5UHMDw6sP0T4K0HUh902QlH0D3csKSE
pZr2gbkhrlT4HbbROf85fV0L5ROWaZHLLQ5nRgoavk5Djy6trLI2jDsEL5cIuz57gmZiEEIlW8WO
xmzSkfFgROijcRNqHLu6eGz7pwJ9d4PaY3i2fZPrnI1wkBMlCAqPBnMyuLcc4/xzN9NWAZV6u7VN
QAJvTEQ9vZ8MVcVTfBN+cGPooikfNgoDJMpEmkFj7GGote+4SE7LTjRHJhyhYersHOGP0WkIxe/y
YQxdC7U2rfrLPTZmXCEqpoGFHBEP8Gb+wt7QwQ8iezZNTAkhlZ93Ip+hsvBikUhDfRBmEpyNKPzr
hZoZIlRPF3HYHxMoByn+ZWtFJ9AhhFJm5LbkjEYRkPAwq9t5lvjatxIsFQqpgRXbVY7vBiCEKveI
z4ZBC0rvXz0bVh1gKCUlAM0MCbDbxsKxMImvEHJa2o1O5YV28w4GCovFbckRfq815pUV2H1l1DNF
qp1lcl4U5YPewXwqK2jtgH62f7JgczglXMpsIyBFLaS+W9SJf39R6cS2Ty3ivMmAd1L5uveiYjIi
3JMTI9miZTqxhKBNOzK+rhdk3wAWWJZMGPJ3RQdI/29anwsIQqG6ojIMZLigWpxwlc8u0hSjcXgs
B5mnAFgoWTRMyJOtrveDRJFzq26qi5MJ0mxUU0TtLJJURBjK7fferm59jqmfaOh7j5Id5qQbW6QN
wUsXDQC1odgScK3oA6DRAlOiflpt0Rrb24UXquV4/cJAt6CCK4PF1ZRNbVNwBvzArgynqzPMwy/1
0yHoN2aTXQPwClf8H9/obB3/Urmm19ztBGvjpkZiZJDz5klAv6MFqEKMN0VNBIko604o7GA5Px5b
65dMgRFG3+q0zX4/4JvrXWl3tpJqqMHixk91h8SyP2tbJEfMft/CiNY9eIrkR86ENo9eToHZOaUq
dfwUscSovRjr7WoZNbx665SEHjfl6+RtR30FcPPTmM/m55YXt3XMHRNfz/wlHkAbaSxmTSYEo5ni
xYZSLJtx8VU+UAYx1ij+XC9iKvTwHgkdHa0nqN2KxhH5mLzoctziPe5Wfbo8vQnMU2V/riDcQ2z0
IlSYjta2Wb/rztkIqBGMMF1jMbfqZuYR4hdPxCiWfXti8p3nAJO8q0t6I05mnlIIfqyr7Z8ZMDDR
r84p6yk5JIcjg9IS4UhyAZldEcvmIEtFwc+bbJTdC9M2u4Mr8r+fihbjflHi3y4ZSHdnP3J3U+HC
goESeM3N1JqaWYTn3rhFt/C1Gpz0/P5zYD5gaYPNcUsnkytuQk4K2ySR2ypuMviVumsnY3mDB1mx
xDjmqMHTYg7BKnNKTMkexKjVUDWQ5VfKJBxiiZnoU9iZzLxtTxzBTGVU4DisCZb0XModn5Nyb3sk
+M7PH4oFh+XO2JA2TWrX1CGvaT6Im4evxF8zEEnsvAbjzW+qloa56UtHvXc8+5daC7woG7hisTew
W8cUWhsF1jI6xH+R9jy4CgzTnfkMgTeMcgW5EETVEHNfQ7+FC+tGIAbSViBCdZ6LbIa7vx9Hbe1v
zcwYLVmIu3VVBBZgJxVvFISk9A2a/a4iEzz61WLffRgoGadJ+/uevqeJv02h6aQ6tyNuvdDBemR4
l1WxjQMwGKT+TdjxTVLf4X0rgE0XxEiBR8qW2qFfNnZDtogf/uae1JYuPw4UgI9y7fMcLJfoGbeD
Dn5nsjzDMZwtnFT9Kxpb3zw0ByR5bRpraJsu3DRKLWsuMIK7h5yuhaQ+IlF/GYPTA2DzoAVGq+pf
UBOQ/Q/KvbGyyFesz8QmImDMsz6eec3N+G0pJP6/ujFHLfm5EDbQErG5bAfJ8yjObDCKbZXY6oI1
Jm75iEpLIe18XQn6cJYIzkQ9cOEA4ePzD+qS6aX2f3jU2BT1jEeV/flvUePfkQ3NvhtDYBNkycpc
TbKeLeBDDCTggYp5VYeqWGJS8cLWLruT8/hgTw4xZzoWIhfcuMws4ka+FALGnv2plIAMae/AP0IX
qXoc0HfucWitwYzzY3ys9RdnbYAm3papWKnq/gRX7BE7vghyOPYxizgnA+3Fkfv6SnRKo7zXOvHm
GQPqCuKHQ8H1uCrQqCbKxrQXfGhjW4UuupzWAM0fmW5GUi6CLXrUqnVAGX94P59b4HuBBO5R7Lbu
DAJCDr0Er7jd6tJdoqhCSwDuRWn3k5c5/aSuMM6UnYE4maxYp4xZgPCcKAhV63GjcWJbt6NC8G4Q
gMQjlOpMmfys8sDWA0jfYEaGnkjpyMadaKnoeyGT6rKpcS3vmDLZOadhOkww0kKngiezHSHko27n
KJ+xWfCqXlrcX7+jsh44VcFHHlvXvXkqXC0Ip6/hEz6BZVNck7LFEQrggdhHpq7vHD67fM30XROV
9JQZlniiwwdNyNjv88UHviWYUHYefFoRTSvlRKIWngwcNqv0t6qjVSl92p2URK1OplyIcVQr3m8X
0W+guK1CbbRxSUcG5Prs+4bfjbEmkSWnAKlm9N7CDdIcbtytfGn5kv4TNSDVnmN2jsLTvs3Ak2aL
0mgKYweYgqmRyxzWFdhK5J7uXnlVuxnVxeZHjnYufljphmQ9JWw403ce6Y0qg2uuXXRCS0Gqw4S/
O5YgzuIUypCn1dS2vT2dzUY0/XS/qfNP2V5TC5bgf8Z/GpYGsze/gSJo5VMZPCw8mfSVp8XAjSIj
U0m4DI0NZVTzu6REbOohlCyWxxq2C+XQiRfSjzaB3adDeWdB9Hwr1Ug6fmEQmBB7giwXg3ArpUsK
bDQnUBY3ny/Z/pkm9kT/GEULiEgwlZOacmxzG/XoQn7stc9mD5jSBcomj9L/eRVT9Mngjv17b5Kh
GY8RQ8wd/EMQUxnuf8svcpV3WdtMmIIH13plteYgTe9rqIqgjRwie6itVHTGG9aoFPp64SH/BD1m
xlHC0cnOegS66KW4RkWXhTBUSlZJtnXNwWvJz0+aaVYn6jEPMajRP5fo+j2PXS9dJY4SzIznOvbD
ZycnqTIj9VSIxBjKyFF0DUhEwMpmPlni+uitA1RCnVRMty+NoQWTjgdS9zbalepRTMEfLLZDzbjZ
QmG7j72wklT34c7869gDBu8HF+YDLeLY+qpABVWdaE+NDSaQSUkQwAlrZcpdAxRd+wb7+5x5dQLh
lMUqqSGjkRE9fDD1Smtvk3EbruRY651/dGCZFzCRZdRneVD61hN64ZdYgR8M9eao/x0IG+DNjjXU
Fjf1d7zq8aR5gZeKhBrw07a8PAtQPFmIxyDQybxtg7pSWCPDNinYzfoILVqMoXft1ru3HxFozqA1
oervnnI3wMSoB8AvBSxJgI2Kr2mlTsgrVSX4lDKBoqCreL74Ogdc/fzwvib7NMht7bt0TbMBL8Zl
OcuOk83bduQt10O4NdCeieR7WGlhkC/62h0oEMBu1Ol89o2nkB67gRPil3nUBndWxgbCOlG/9N7b
W+MeJ+HGYC7ajHeem1jCE7R9zU869wUsXB7prIkSDXleVlVwtt4IDcpv999QTC8rkJuOT04zfe3K
M9tpnq5PfFL3WmG/RKN+FgqRn6p++RDryGuyHsJYwQgftqhLVoHtxH+lr7vfezCcrPLDtpMbfmn3
HhBU/y7JOgqA3BeL10CPxYMz8VAw8Xax125lEZU9uoGOI80aUGsZDTzTt23hvvM4WLfumVXmj1X7
Skwt0jow3VPWXT9lBaZDDWiDNwAC/fEg0uxpa0ICQ76BTXaKKfJxddqpgAhvoTxOgzkR83Q0f8Vy
G0VXa2llhNjgYDXMnRO/jayRGRv6Aiwwm1ChhE6jxUX4rXwWS2e64dRp6KyYrlbi2I/3i0FlHoxj
uVGzzMDdvSPuuPz7rP2CC8AyelnViBH1Jx2kY7EEXFhZWXCEcZfvD7NjnpkuVev1LKhps+vqBRTh
FEB/ARVOjK435Y1F3B9fDccZj8vMY5zHNpH4chsjT0WXtMervePKlEZBMb+f5InU0lHaB+2aQ6tq
LsUpLR7wAxXV0fwY+ke7iXRP4EO37mCe7kjN8X1N8cgZDd1WV1kaEWS82nvvNc2C8mayARWrSfqm
lFdrB2N5XANfZFbVC9VY4k33Z5Op8s87gT1rHdYDHRQqJyvXGJy1cc1W9LDwsdUzwBthN3vnXqzZ
3iRPYtIGuApNzkpkhHbXrbtJdvIyjznIxoZf4QcYHcB8ARGrPsdXll79C1ft8S8xRYIYAqKgw/1M
J0dmqI81vy4E8GRuWjt0KeqMpc37zhbuVIYO5NGfEVjyF7IbZEhwKlNl4MTJAKh2hnf3XKmNflUG
kgmEOOHKumY0JgQdylhh/YE3eVSYP+sGzRUVXILsyBXeRZrs16k0PZRoVtUUSLOkQkNTqDQvvCll
2wbzszzeXWxAiqQ44GXFNQgCs+ZMNF8GA11yKAFFOPTlr7Jt7XJchUhaU9pumDMuMVdN4P7RVK+j
Hk51qxGM1Yg0m1VygvgA93Ip43wliP96PwpIRAADoQcNb4ho14tkdEYunfx0wk9L9ZG9+anxfrtS
tgTLD8TgVlvalYVoLyV1tyTd9h2cS/mv/hG4DdDa+quzbZYG9RjduqVI7CGruG+foSDy7FoIvOsu
BembP8V2+01Y3SQ1esws357zb7DaXd9x36jXim4KHnuUmiMt2qj9N4hy+YESsr9NmWjlbR/+ICOn
UCks9Y4cD2JWeLjn17XXwEIXKjliQyLjgukq0HoIal/PXXwkJYGN7EQE+D1ZNuXflbhwzAzg9U0N
FEMLJyjgdiI7iAy0SyqyOuVtVUdMNPBfE1kXIXGvBAdJPFf2kjaUUu+DZlrahEqRZZuSxrRGI2nk
bih1uWx9oSo7cnmc/PyJvQRRZ9tUhg1XbpWViAmD4Iwdh+HiKDJTdrdX8cOrx1T9SfoeWaGVAVVv
8Klv3oxlpV86i1U+Eg+oKuOG2pdpbRVJ/Htl5NxNMeYReNRXP2PKXZnZE4XQnv/txbc2JBvQ95G6
AQtukiiy17MlRZBPlRKdA0MhbqdCzhLSjhCT1d5R2Ah7x3i887q0QtZgY6wuh3geM2l3SqCtDSyB
Bnb32DHJEogZutKqnca+GV3Yt2Mnvzzxg4zV4udCRZy3u6St+AOcIUXPcNaclHQwG2kX3cdmrSCJ
ypz6tD3hpiQq/1s5nLBaVeZa+2OS8RpGD2fwp3SVqnNahMgPcuhv04fwuB/FIPQrJdK8eJcuIo3d
2YiaHVrglMc1AfpXWSrSZEbtIHPT9+sO2tXEZ6vjDfXGSkorm5ivcusbm07V60p0shcQ08f9ctc0
WvffPi/W1gP2nWEYIkz2nI3Ys83gEk+nJzOp/AihsLPMNmweFbw9QwDadHteBxpMnt+kg3HO/0NH
rdlZRTuRYbaxxSC5CFhpYQdMiSYfhfCpgfF2tVUMw+Ex3+TY2xcfL28xT+7h7oU5MrBzM+rAyJai
APKESKQdA4saKq1pj0ZlaRs96DFpS+YYRZ37qpbmK4BeNfZzAWSBSkcl5jQ+pZP3HfKGwoVXCGu6
pMvqoDNpUWuACFXFiDYQHYWNTaccGLl64MXj+IZ2Dd6NnKtuQvl/HY6uPaWZAFDIcRr5GRGnOsmc
OOQvt3wzL13d7ZSwHgQDt8MlWIz+pU2b190W5D7sDrjZrzB6tFjcG12cbMGdjfyw+kNiVzx/LJPu
NM//2M4U8TgTKB29suzR6NyommQ3MrA9AoetBawzjwGbGGWetDRqw3Qs2WHGvzi/59xXTCVbQuVl
oTb17PTk/4e0YpiAfV4QBo6slZrN7Vmmj46ZycMcaCjfqc1jmez9a932BxOfn9AB63HhlvARDs9R
rUBN6T8DIl3uIv2R8lPStfWNopKgkaiSsEmFhzHTGuwARc1BWvPzx2OpeqgebErTVVo8X6Ea71L0
gNgjsLhTHTkfKU0lbeHT+5/SSHxMUfI7W7hMuQz+g0PhTADNqyTYkePYMrFm67w4iDjIV3dy9arw
prAD66z6hipke//cy8SQjs9cZgSLuxc11gaqf60a3Qhy3Oduy5iftXCTkrK/DB63NLNb9VjGArBN
qshkA9DrbNGhsZJTwQ4CyHaZbiwhOMOFCeSc19RiuavXEWOxVp1SHd3FKvp11z8mM8w9Hubfpk4F
RQ/bmbwO9j/Uyfxb9UyIwV9AmNllloUYpcTBF6akOFpUVWSg939CYfXSfI3zxhl0vOY6A8eVAByC
NIaxKS8BrHzC7CH2/ZhEOJj/1elhUmLvrWZPjLSMriuzrHasvxQVG7+ybe9vf6VDz8V5nvdIYCKB
0KPEO8m7ooi5Nuf25OCU2hjCMOuR8wd0HFukqSLyGKbyPjIq3VYE97koGqAdIBK3Od6TQCqwCZLx
Z6oEl3cKS1wdLZ0iLoe2hdmXgngvYuBS+yrlyqOr/eDCp0GdIo9pY5On6pMJwgLmKOa1eNJokvt4
JZhKqg2yEBOi4g8VmMz9VVliKfzenePVsY6rcodanKhXM5ZpweFph866rfmtVKDy1oZLdX66Ug+L
OZyNUaaG7dKQq62XJ6edUZlV/Po7qY2y229AHRQrE4Oa8hCzGiUYxfj4oeinJ3OtfugHS6bwcBPu
1Grl5Wwzy2YkNbJ+9aI2lBfIk9jIdYzIFz5g1q2YVSBz/OcQvdD01IqeLIhlJH1hoyqq+W1aemqv
LmBeFCpxJl0+04tV27IbKqvigoFkgYWHwCQiawr65igs0fMKb1S8JaebZZdFvkFmFiKo40xGHZ5v
aGuZDkExvshWd5RRrBTl1pap/LujuaPUofHg9GDr+u0dvh2VNq3EC2wzPDgV+6gCtFawzl3BBrRZ
NfYucoz49k3nAmFmej1c91p5Fi0yq2j0RNbMbjxMQl6ZVuS68mhtCG6kynkqgUO8lRMuPBLDSrUJ
RuCqoYWX0s/AEJVJQhwf48OYkxnkclF08gqEac5LPJYUYRoqIlnrC5yiPeg75qX0OyYMsBTocCJM
FkzcXZQoflNvapUUPeymYufSh2q88RucMs2yXSIHfKvI+KZttOVEOhInvQkWB26JdxPkdqoQWeBY
1f8s+zJO0GpP+FZesDm1EoLGBuRn0aVYjEuGEa9FoFO0G5hW5jCp/PdXn98F2T5u1ssV77ImrjOu
lngvrk1hgpgYyzVdmP5gFt1eB71LSGxN0aSq3ZzIHIzHZjfEvCTBySCODa7xRcUYgkXNmrNcM6BX
8LLIdOpSnRKOCzmIce517sIv4lOn5zE2Zy7wJkwtSMCGges0Nn3CYeyR6rDbnHeMAf2zBDpUumF0
ZZaD9b2IEfCIGvqvSmusSbuKg+IX1vC3GlAn0LTm/kARVh7lux7nEj7IIEEqdGnzv+F0CNXLbEjn
Cu7A4LMaiY9YBSoLrZJdgYNiJfZzD5XvMp7qSSAWO92471fb3SYvpvzWmXMpTwD3dEHQEkqpkmv0
R+/xPTA/PfMcCkbHQiv2G2VrFAiY24uN/1uZeBe17Ld3HFrRJAOJqWTGOwQWbqmTnCEWIqDJx+XW
JMAuZKhHU9nc/6k2YNHnssNWtWxOXKAkzsJc/F3sftUjl7bgOYD9Bibd/s/vWVY/d4qVwGiQ7mbB
1o0XxDTAahPU1+tbSgixNO7Gq6Ynxxv2hxvIaArx9ZMPyEHCj+d06ttwy3gnLPia8BCajyp/FR+r
mt1YWzR4AWvp4fotfc0LLkjPql/CKHvrq4FkwBKj+NSv68ZOpxjqJjUYT9EWSit0LAm7AGQneysX
qa2yNJ3Gqc213UFpghbc/ot1/MShzfar44JJ6vzLxDmE2W00GQeSXsZ7f/3FtEEEnsRDGoh8hPL/
M+e34Kr/7gyGUQp8oPjjYU+DnZLdeXp9Cq4RK5yyGFsxUAjJ+JTUqb5CuQSjgwaYIbis+ZJ/TYTT
o178Hm0cudnaEeDNaBD6gL5kweM3FxRsUBQDS/wr3y1eFYFvbEEzjbPVCOMZ7o2eR6P18J54j+Rd
qvjfDHgRQKDeLOG9GDjGXELcGqc+woPCNEJUP4X6R/EGH6qPPAii/67zjp3Edfprt0dF9S7FJKjH
0GxljsAlCBvMXILi+lZK4M04A42jwzzB7sXXA+YgekoegxHrQMELt6GF4tNUV9kY/94edaAbw8O+
DsCUXmHSfJywfprnVLFx9bqJo6gFJztK1KtWKJKtfh5/AkQK/6VQHqz9iNJujwCa8auogLOVkxug
IJuX+LTeVYh5RZrhwdv+SmU28VAWYPiqKuZo1tig9rlplIz/ZntEzoWSHG6WNBUVv1WHbz7I7vnZ
OECAi0ejivIiCmjoFlq6vGEzhMx1ha1ekgtb/jQ/qv03SpR9GZ2GeKp7CBNsKTrcNnWBPQ6v/7xD
0wAys+MeMZRlXnolWfKlGDvOdU4CCOQZ5b8L+g/dmGTG5hwQYZZERmMenVixYJfxUXsQqvBgyNTb
wcvQG7nTTmLN1QsINEonpL0Hwmixo+ZXgwSy0vHj4vL5VZtl3UW/JhRnKE7IVfAqZ1+ib9N4lwT/
IiBp2A3jDRnmye5xG6C2wkEwSQFE+Or3cM2Veyad2OeTa58PT4GpK0diqC7J8hRydsHKkGqErqos
56TusZJ02F7SQMq06kZRDVCVl8UzHae8xfjDFWkAJe6ODY8lX7p0oXqWODfdKkdxe9C+uOc97/9l
fri8E0rzHMhOaGnuTWTry8Qnb3wsfyP13h70LkLDbYHQUb2wr/RIatxYoJWwI1WqG/j8ZYHi3bao
zBFO/i3kAjjeotCHv89Ok/FpMTN571N3mfQw18/idgg6QBhdyH9q8G/Lx2NhTmOePQe9hhlcA3/N
aWXnHfWx/diaLARBN2nXDYcNLgaUk96N+jZaOU8l8nzbwUdMdAPL5apryGXoAOYlmJDCf+eVa3Oo
2NrvpG3SHmcmuOEjc9bA741A3UY4NKCBZW1eGYrC/Iv//Am67eAdpvz6qCd2GtSoxmmMwhpwyO/c
/oePY5f4elLHtr37GM8UD5nhUILkAV2X1yUA2pwxWivsNL6ZxJnvgKFdRO9it/7fZ+NmQRDzmBjQ
jCsLZO3juKVkJV7qzVE9s69uJZdu71SKH4bjR6W7FmaSuG7ZNLqz+N5JG2O47HwgDu4TDit4uyEB
WKKjTiB92jfJ+Dw4xXFc6TT1znUeJ5/ul7EBi/PAgTSgIOPsTJM9uK7ak9FDDiaO3KlcjfFE7doh
AmAC2cTt/pJBnv7dz+Cgf340JDdi5FDveWAzygXvMuIWPVzvEZAY34FXX44EHWNOK0lnqRL+mg8w
hcGyJwHhRRZC94qYEQh28YSYG77dXoFebcJsp7/k95TEuoZZGkZ0ZTk+mKacW+owFDjnpLbB/dMI
P7W/x0WjR4E2HgTltGYbQi9sBlCZRRdBsw1pFwfQKWUhN9+D4xeGiogyIZWFc/o+Wav7RCDyyeYB
Q+K+DcxywZgy0eD/fFe+r8/cJiY45pCxpcxepD4Qbp9aQ56vpRL1/+8k6FQBOvdWzropjnj9XuQ4
9OSaUsvaC10rzKqmG1qtixdP5E6TK+7jGJewso/C7QV0/iV+1G+EZtagkW6n61cW7mR8FdBQN8RB
9m97C/704Pe5E2pNXChes6s3W9mpNTrqINQ4qQYbpJ6Ru38bt7zrWtNNiaceVS11CVlfjvHHclsD
XEbbQKPenzmUZC1rJJkNcqCIpGiLWCxbHDgjbrJKzSW7IqHMjF4HnlKXEjjjywqhy5boNeHJJ/Vs
8TNGt8c6dKrqot0/PUW5uJW+6QdtRP+8wq0etIswpVNvgvIHImjemhIeS/g8xjRHP/BK9uC+MDEh
bLs1cmxx4o2La4Fauw90D8VBuXGN7VKykEawpa6wNV2eNKjcbYWd57rTI+hvyobaCUFHNLI8cK4K
DgHDbmlbduJ5aw1Sn18IXdZvarEQ28hQ+JPg9Z/wvsFnkliaMOeKImg4y7oylwaX8DIT1kkU0xJa
u7xreg6CUUKy1nQf8QlwBrOEX5DG9eiNqoOKzzODeAA/ceqv0uN3O6oNpFgLbzRVxxwTaOxTifuQ
BnLA06rqYU9H6j9mY67034ZUOkfHQaAcp2790Hbwp2vKCGtx19cj6OGYIUDLVKnwYmLX0jnvsvEx
6tlSyMtPQPVVtQSlxONo1sGlTlPDV2co97+qy7hyksBB7y22AU7XVNt0wLThU/JMdzaewyT2X5ln
W1OJ6McGs3L4pW0zxNvDhHJpNSS/y1v05em7pV0FjEVvFhP8nZDxywnKNp0DP9Jh6SacICv3BgDr
dLmxMwYSehwCUYzKKE1cvdxR/f20mdXm1iOOeDWrOfxtFkGTyR50Samre+0gmDCkiLT9qb82qcNn
PJfgllrg2HWCrK9Iwu7wOMY7d7zxR4lpXD1MEFK0FsaQ+VY9evWpd6H7HjtBI8rIjKdrvJ7/WFkt
y0xgeUe5IEidTfDnRDX8ZquieY46dBY613IS9+2ATKYoTOiPNxsn50dfNDSeOOdX9jQTipjPIgwu
4S00LXp/rNz1amSb3kP+Tj84Xq5bjmg5Vqr9wS/FF3zIlQZBfMwsVdiSYgimwXkMABNGbaw8rjin
nji3qF5z5Vjn9eU28r17cxaC2hyjvRVNyjAjCbqZa5JHaVV1gyD8ZSmXr5D4Xbgcy5CWJgGLKoIN
VYqEaHh0VkT97M4dQYNx6HiqnDyI7SQg1qaosHlGJNF+I0ivtxVfwMlHMIRF36KPSs1bFIEnryDx
leaWdsq5+iv7bCplccc6zeyO9vpbVudbQoC4iB631U+NYUaamBjNMU9ioLiVcPYHtWhzfOChUciG
eNuI55J2JfZrq2BSSabFi67+eLE51PVPF3bRrW99EiUKZ/yrbXR1d2y5udyvwmmtm6WTTSvTF1tm
I4jvnDaoI88fWS9j8W+vK9vP0q3q1PsCua5Z9txpKhPsGL9kPDB8TuLb3LP8ShbG0gX/pap/b7PN
wZvSL6+8SEkKHlZ5+y/YvBN10iDu7YKs3CSC66jD/4Fha+88s0tJrZqfMkEwFDL7K8P8rT3eOTDB
ldS/MxM8kh/XxM8t3zEuCZ+Tg+b9qrKg1yBYxlXas7TPa3uQntJbJsGcpdV7vwpblCrw2lGEwRE+
TVjFvHZ5GhG2NUCTFGQTjqh7eCe/CNcRN6Dy9f3bAtLEOknCLR03CzJE4j20lmAw1zOP3YSKQwBo
DsrVW+30sEJK6/jjXH8Pv4qmgnC+KfE1j5Q7mDgzirwqX9Ee9nEti64NhBdQkAHL1Ql1DKz/Vp+m
8BEWVMhKYxRHuH2ZLhVHCW52swNW7lrNBu1W/TcML+GqOLB6SukavlMTWA2aTe/LRqfWqRIGDjFY
8pXs4911RxCnjaxL+i5DyrRPitTeKf40ptk6PM9v+ow9BZiDdlihdp/VfjpuiMqHtu7+ApmXB9uF
tnTeNiOfmYpZSl7Ot0wDrdMzajPPIKY9/jQ6eVIJqwJoOxhqqbw6Fp8B9I1XiVy80y/La6lNY5Cv
mUzeG1vf5KEMeQTLDoAKcVItaVIPWql4pDEow2bF6m57bW1/EcFNY5lKZpD3qz7KOhoUy65MHeCA
YupZWjunhgJhxVszUuRO1Q5r8ksqJrofNnGLL+yX3fgp7f9RtS2dF84ak0bs77EOH02rtW7x4MjI
X3OSdy19W172mUOiujcrDsqDM84qjBGTvt7Puv6XdY4b1l/zYnuRxMvmgQiIomDIdxqhfy+0VZna
oxBMywI7lgojuAq+oEOIJmyi8cSu/qxbYdvZQQfCwvWO/5SeBeirOVQR1/7SStENs73aetNGTqAS
QN6swL/HXC7B6yCX8mE1eqpURx4rX3HrcatNhVJM35/057zuWOrUIxGQCx0+oEoALUQJ1WDosgJv
F39yMRH+XBYRJUTPrHafnBuuh/taQdM2fPiX4AdFBKKXSAr5itIsGWgHxsKrduFaoJz9SmffbtDO
gp+7QTn0uN/yIpcPRgQl3SKwKOl5WneVwz9+NbWuIufdhe458u5I+TEXAV+Rg5Ns6FsLjHCdEZV9
pihqAVd+pnQbU/jZOFAXh0xWa4611TPW0Oi1dV2CNqmgilVaGgTMr+0IEM1iq46zdB/yrHvlSeml
V3bvt7znIJF+A2hEjCEManQAo2lSe3FoykAT5awwEEtHtZ2pdp5ZGH/ZDEPA2bS3zDI06uxEbOmQ
tPSkMW40zB7z0jbAAp6H1NEA2E8FB2KFQb0AccT0HiIkHq0TrTQs9QDX58WrdlqhjjFLW/uspx7r
tR6z4pXs6czJB4ifWYgjlb1IClX1PYh+ujuI26B6VDSEKfUBHPTjFlSkPhJPbE5sv2Qerl2y+nDU
Hzz8qYCGCRNnU5dW3T6XDolpuaV8VrEQldH/0q0BEcsrEdfef0LcMge1LDysC97h4JT2Fr7KCrlH
YTIa/I8WAk+G3ydy6DnThP8BzJFVDN9Q8CpqsC9Dsk5e2ZaW6LEzwJO3LXONfhTUL6WFH6557Kpq
6XFqGTDh3hm/i/GWErUjWXGvGRmePPayO1nDX1v2JT5tzBVrwepEbGSSvbCAqDgmvDy7H6XnzoFi
fe3f8QBUtT+AdKUlL7aigZKpIewVMcNVCZz1Yv2iF64SmMqUR2mjOmY1HJRc/HNp3WS8Pv2AMj2+
AtJONvQ8nmiwS5YcVbvF0bZkMbKiaEIzkm/Ywz3H6AxxJJ19Mu9zcwJXfBIgG8LEy+9/fD3LN1WK
JzNIe55Iq0FEi9/mfE5jVdPTWgswldl+50OPhqKyNrjTwsxRg/FPwVVIeR/9e9ZPLW76gsjnoOZY
Tve7R5KGJz7pYLa5lDq9+EoMfha7EoZU2+PBxqn18RNp3FIl3QxzmfSgZS7O8CdgxLrzycpyUGVx
GTbKYTpJ4QqtDGCYnSfap/OR3AxD6qqTCa165IfClXjLqXcFVnD7Zi/8/YaMZ6PcZE89egTKhE76
ZCk1/v9sAWNwZV3J0aTb96DbDjlVRYDE/1CLytfu/H2HEVTvCUxjQ1p3vqc3CK9K+5Kr98bBEBdv
NLLYBeYf1WzxUFX8jPyDws2iFdZILSw/22BsVe9qitAH2nfdFoZBHf90PaP0XDIp+Fo/zGsdYSvR
89p63mcxnX1f+dj4l3syXkW5Cz3iBm+IA+sBocYNcxIoFsAVP5ragHboWm8C+NWcvXV830b1dtuN
s/gYMMHy8v4reM87lWU6h3HBnvRyzszuVEu5zECx9fWYG5cfPNkXn2REAVPcl1DBkyU4lnXxhf27
14ATwkyGpmvl8vPG1VqJHz7Xmx23h0cuAMcv3EwHaSasvXbsSnBD8f8/T0Mu/L9RsPkvjQlnoqo1
mPA7hmLEytTLCIlRtS3BPWAELVF0A3HymqT98yiE3O9abHMdFjaEDgPYK3VC1wAg3ewMg33pG8u9
3aKrUizQumOu+gH6Hodq2RF2RrqrX+dvukLDZRJw3Du0U8Hh/9WLg4TW1hui+uHVvLwb0VfY/RtQ
LDjQehhnSq/zil+kgAJAxnfNhLAxJMtyqkcxdlAPo8dozFx5q60zmlJNnsTzlkr0IjFSG243cycN
7/fRfNFfSaQRVGI4Vl5HixHhOczmooTQPGypGl1Ol4a2h55OiOCq7LDjPw8UJ2S7xuvdIu4GsyED
xer1BaPkjlfm0BkBa71WTx+J5IzInrQeqEqW6i9r9xTIB9WcQ7Ei/wuFmygr6VaQeqsyG1Xh5sBy
8iDYioMP4+G4ws7remMQy1lIx0uS5Bnhsu2YsJVBidBIowzDM1ftkZhR8fW07p2GlZhVRxEZWlZn
KCd6CmDxSkSIxJPjx76axnjvVTV4jR+/T9jJdeg2NZ5kwpZ43xoVg9nurhvTVwyT2731+IWx5dyw
KviHFiv2b+qWXqbTiwA34O53UZYLqeMJeGVXTJpOZ6ejZ0geYP6EIyT88eocWbHYl3bkMoERro99
xAr9LMTr4uptbEUUQL3Ji3uTLRKj1ICIl0AOxh0HDgAq2Q+JgQIptpBc6OTgnwbQBb93jN8Jal//
nYctvsEdZTYtjHjoCLHPajy22yiNd4AaXpKpAauEs0xF2jUEQksZCA4OarK1/zO67HuNW9gsT14W
A1d6/f++1aARs1vAQyko7Nrp5ArCgMgQSUNNEhfajoWoAGRkvPWdh5DYxNhnH2awJ1RlUrGTlqfS
qNf4cg3Fhy4rOdxjxXaE6ZWCTJnVjS+z07gHkFd77+tP05OCSDq5K1RCs809CuVOk8CgYOOh+piH
AhzxNe1BW8wzUUFWf5gB8K1HIan+576Bp8Fw7IiyaQMD2F3C4rEvP2NyALJPAKc/GLQcyNpyR/Ij
ES9lXAa56MbgBQ8tGCm/tb+gIic8yz+FJXTzZ5VMmkquhoUsLuMi4tq5uYJFoy/ADh5wHTu9yoY5
4drCeVyrDSKv1CJJyeM1lsRQXvWRBiOBDnijzR2fMwejxxi9KwR9Mr/MJsNKnp7XY/AoWfOXPIVi
bZbPE+LkqMi9Tu98g9a+pScukOKdbZBJxcp3Xa5e7ksMBObbvBhCae63TFm+S0pOJ99heBfPozD0
/wzeFbD4IDKHnchRiEHQ9iDz5lxKRrjUJZYS2dbaH63TU8HV0NUpL+mjCbbvh2hQADogk/C2J3l0
gGYESN6J6v6ttGwBObWabkZKyo7Ey6v50FpKnHBmNlrwFBEKwcZyFwgMGdndyIXsM0mx8RXhtSAY
b7PWv4yaKIXr7N4puQ+pggaFdvIKWy0EoN6anRGTgFiTXfmGx+LOUCHCSlU6SYEKNGlPXAc8eDNk
MstRQdzPxpXTMsKYcjNcbzo/60I8mFc6fXexdXj8n6R1bIWfHSeDGY18eQxeQQ25hc5ZzaYrzCuZ
/ye6unsrbbyqY/PqspOFkGzhWDsFhiyjwh6UwCciaZEkZzNWVG9tP/bLNWuvOKg5QS6Vb6J0jPU0
lITnRcj7xdGkAvpZ469/BvrCIB0U4ZiiNHj1LhCbOG03dm3gU/pvs9dcRBIBHVqpM7qCUhe+x44r
SBC4TyeT++hNGvc2wddSCWATp6c4gpuTdRaMt/h+NaYp6RCY0pHhUYU34aWZ3Xkmd3EFOeKDBvAl
E05MSDLAoGVonUpXdj1Fo6bDtQMkRlc1/avcgH1HP0Ib4JmRzmh99Ec1Cg3dooCOSy0af0hFsNVe
bt0VYoFmtsAK0R3NDp4k6MgSRJYI6G2TN9WF/Mxy895rBEZ4H6SsXQfSe3dOp/eRUDkHeS9MlItx
gtHtoT8Rary0p7yyGwt9AkhUwqC3o4M7DTugWjVq3Z5JVrLFVreJfAeBg3ksjDEeYJ/qgtrx1rRK
ximVvk/f56Pz4gENsQSV6/xIcfn+LcfA1Yn7cjHz5AHRHQ38h4ve9sPniOBdbidepBmut4gc0Vxi
g5FJEY+F7vtTfiK6plsbJofJ8E43ptNskTDuYfBJmI/ofzrStmipoordDu6ezeAkF7WUVqb5BuM+
w+iNE/gEsbDCUhWMPYAaErtiUzFYKrcB7Bb45oSuvMpfesFIddr08cacTa8WlV1JiDzimqfEa179
f3MTGGvIeRj3Da2uWVl9rRcVQCRzM9kzPJAY2sxbHkxNrvGlK7jOc5lpPtCVDVPNYrodBIJtu4tD
tetowmudWKWWfYj0OftcaqvTln4P7rXVJ0lBjJT4HYrVImsFBM2Zg7VM8gKdqcDRTBr35XS5jH5M
FzU7tqRQKGJ1ZcQhOxvCC26i0eHNFEo8l1SmYLuI32JAprXx5MWruPP09h/eNXlCIChf3uJFlUui
HhPiidiYP7OY9C3Igkcbg4deiW3n7x8aKOww0tmN4nNH1trOteZDDbYR7hCbYYT+nBLapDQVXseH
x2kG4BIya3mKpX23pvcspK4m17UBXhRh934elLOCQUC7Wyom3XZRqSTRLhYh/t52lpL00Iv7U2ft
CUKtLcqjr/VmU8qoPUC55N/c6CoRBHm/C4rGlMBnVf/z4WA7jTNb1RK5EYtAC1l/gMz8//W1J0h9
oURgwDJNJCdJw6uRc9ujPuXogAy9sYmq2cutq04PkSDlXrkgQKTzye/hdUn0oRxjBMfvao3senni
7PdD60DzClOzynoKzFth5X66jhtdrfpG+iSbV38SrWxwdxuW6uSg/qb8M30YMDrsf/kVYiveHVhN
Q4VElZzhvcRm35i4PVb/kyOYRYc+4wV9/Sx6UHFbkrWpmNhK7tzaNT633U3YFtVNiqlL8kCK5dKB
8VAatxW56pKkHCODJC/YijfGmOG5NhE3pnKwbkVJ4nvTPGrFhB5B9sjw0NzXawvMnN5zou8GHOIG
ZmfQ52sqrk3rm+2YV5MNo4amZeJRj7CfjdjM6QVFId+NGhBkipBXCwBC1lFKkYjwdqTTz0xAiSNN
/JSGfv65/hDbnm1wAhn7OE7xEiZKiX8gqY/MfQRxGmxZxgh7opyVSC7mJK0jrjw6qvVDz1I5elXY
5u0Fgyh7qFYWWX6o9bcV/C2B6fFXOolihnnRi/2oN1WhzSt9hI5QbW6ld9hQx5OiKED86irX4i98
GI1hUk2etEVffXwa0WNm8rGAJ8FYpliMl3M0lWlYcnCH5ubwdxJwQ9tdmgOmYcAhQNpVnR0uDRHM
00NSJVVOBz3hdCP09dBkaAT1c/lfM2vfmX++6qoLv0kgYxs88XOaSiumstmOWxL/ZT+cN63brhq3
UPqsI1xm2K9mc9V+hAfkQS3R9or2qDCTCrk7y79TUhVn1WaM874O/5Owb/3vpmqRUPhJbW1vyY0w
WyibL6vmL/2wH++gXmTBt+tLQQZ2yejYWGNl5sGUYDp6azTo6Rlcdd12bxNyu31jIJGQrsFX1egf
XoycrzGIejuBkPj9BKc4f2sfkQh8q3C0ui0jEk0kkc0RZ1fk6pBgI9xNx0oU/o/bgxTDWwuwRb2A
GXGkIJzJwTQU1cUrXKRWGi/tAvoMCNn3edvXpWjOrnpn50ijHeqk3/EDwxKh5EPD4cIpJrdeknUe
Q85+F2qHJbiimlG3+4Ib2lhHXOQvb2gV8vfTzuwrn5zSzmNeilnuoPLRqBoBKYBruV1IwncWWufT
ZKFtx1OltHW6y3ir5GkB75+45/aReldqPjMxiFO9sf91GfnHxIBHjt35y2MrjCwpUqTvU6hrybNS
jLZ2WBpgafPnNUmUby1wmCk5UC0LeiOaYGl/wIYXi0BXEFDEdAhcdBXOt+zkYmHN/pKl1bSJuybe
86bDf5lLx1+6BnOKM0BZwAQ9TLw6MjNS5qAki7qFl3S08FqfmtI2eevD+A9ED9GV+uSJENPDu2Tb
+twoM+UkJ/HfgTMrjClJ4dxDXUfQehQaA1bsT3dnmq6t1L+MQTHzr0ffIb0+apyPAoBUgNqaWgcK
VhxuVZ3Em9PQN7ShhMUrOMtt1B9F0qzo1obqp8N8Y71rIl1krHFu/cohDahBLlaq0IP1KS2p8Z7G
yED4DmVwhliDKbjA0RxB5RauO/mfISjhJZCeVeD/G1wYS4xZa40wR6nGtaihKpDVolK+NqipG7Jb
m74/gQfF6ifQkF5XMwPBjkiP7phNNlAt32PrJBjePnr7wQNpkAThsZKC5oXoAVPqzn9MigjnJTGm
F5VjaeCX5c3oatSQk+D7uD5RUWu78VVhjjSM/T7cMpvuXdSizFswx1d2+Lt46WZ5EhLPp8eJplee
BkYSQZNhwm5BbjZ5kXMwybLVOPeN34GBRQ5hPbweBBFOffqrdlfbQGGOhBKDceHwmAm8ZvSJoIpV
Vg98TBu6mP6GUkCy/z0HLX/rpPrUDiv/Pak43XMCmpij81I/Xu6ABeyX0F+ultr1EhuXBHaK0Ns3
5SZ3yYC/3hfTfZAmMG+PaakvzNv4OKT2WP69654V2DWopn1mqGVooWwuWPnewYwhUaOBB9JlXT5B
0LWhqAESDPa1IO27IUyckTgJWXJAT1XA7PWQUxP4E7qwV85apl9PiIbw0iPJNkCIIbGv9m1QDS6w
W4PAbmFj/9ErxWCNVO4DfQ+OzRGH0+HMDStMiO2X2wo1VvlIOfi7zhG+zCuI5jltWoI+0jLlGq78
KppoeNldUeESwIDPO7Ec7dI7nlVkE79UapJRM9ASn/lQ4+Ipz5acxcEHBR6J3MPVrpn2+XlTJrrP
1t1wlJQeQ2TGbvVWadJ8VgsApCRgbf+OBznMt7gZKz2EYgJF93b07ITT8x8scT8WIlanGILBqcWS
nVShUluXbyFeIMnpem/TsrftO9iFIG+/C1g2nsFIQUh27g8JutW/hZLRaK293P+m3mZK24Q0fPzC
otIM/gzIfgqyNlXj0NwwEbkiJARnXt1n/KxUgnsBuwBubOC/4xE0vrrXScdjyhaUUanDiOrySM5G
XLGuHctIUC3/RN+UOQDYppJ7XXdLcth6+ih9cgvJO4cx3igcNHBVHQpcTixdDQVUOfkAfBatm/Ai
bfCkrp1TR+xHJwEIq3dJgL2YIy4W6PMnPu/mcicPmFg7y2VWtv3truU1uKOwDEHcNy9hAlgweYLj
u+Ie2WhCUfBqGf5GeD0Ujy2JmBi11CGUIGyiH3Yd+f3XolZafy2RF7dYM/ZfmEWIaxRWvZjs2Mce
camBHE5ra3rhBvy1Pq2S4zczbAXFzhBS+Xzjm93FxTk68zAqLJgge9eE8XIqUbJGkuOez5rYeCDv
f6f4THJwRsfjI6in1eZaN1sO+KdVuUFCAYg264faASDGZpETaRkZhOCAAZsrY9IZfIQtl2jtN6ab
vhM5JZrc9G7lCdOh8741A0uMqe2ZjYtz4sSEAcwmd+FVgdp7HrY6E0N9mVB/eyKsW5WT5My4st40
9psfg4FQbXwxVeIoKCAd5tgXn2vSxvxY2VzW/ZBxQJPwxDru64SfbfAA1mj2p4cfs+T3aM+zdwwV
pd2IuJuvPmCXIh2xI9Bis7MwXkD5b7UgmUn4mIg+Q8TvGixGyRVPwYvzIPJvVaK4dChLByYfkX1l
rNYEvtO9drVhd0myq5EuYush3TYWa1jruif6kjgE+iax+yh2TzVNSJ081cVPM6WT2w/6+TTeCdbf
cAr3ZLwqv2Lb+9G7qnnAXJP15xozSM37rGuMOakv0+xKZ5DV7Um8bvWGA+acVr580o3n/KzTeFV6
H5vMAQCod0N0z69seJSldwtV5bt48QRebE6bl/SO5bG+3IRQ20gFvl7UZ2W10YNIMB53qiee9SqR
wSEppMjklfvshZspZOWe4BXQLtL2SIlfXyV6q/PVanQRpltHCL0Od3BGvZqb/sy/z+2ZEvk1hIKF
zq2iWsn1tW9Yx1g6GdQxJSXk7BYps/ZrTVAcQ2VeSlvCCxtSbrfLZ/KA0LAEm047qV6XaQO4zLQW
5eapreSMvBjvUHU8ukvhT4h5bBct6ULfN6GJFzrq1a5gPFgIFeIIBW6sfEAVqKTfSaFvmb85/7oJ
sjuZsttcKU/UR+7pBLkmcsP01bvpJmctMxDA+MTPyw8Gk2ZEFXBk1xmwODwcWpVEGEJEGFcZFrgF
Ncxg0rVKzYluxZNqBAbpB6tfoiJ57ELNEOaCPzNbA55LUhef66ZfQbugAVvg4g/ZQ/VsRVg1iQYk
xAU6kpKIZx75keC+/wtPn16yr9bCXNDNd8yWR6jlX4WWC1MU2C0uB/nWS1AZQjbwxa+ikztitqbR
+3DADG6+Sc7swb4ZjdjxNXPFcALppc5GpJ6z8zMeeCHiev8Pc13Wk1YX7eAkRVdw9ubiFtjAgonG
tDhIIVBUFjqE4TC48BBdActA6Rw9LVY2o9tKfRYLtei2VOUuN26ausgKL05lWlZewylmgmaokEkC
2+n+BwkvbKSCbf7iA9DaudvkF3vDAT2VQIKu0ELjiV2syWh0HaDbDkHsD80TG0rDrI7pe146vRrJ
lF1OaKD2NaZAWeAl1BQ0hmPoRXiMcrSO0ZQFjZ09gFAU5u53TfyjmQuRcHfQJLeiqbY6lRxnjUcn
lDd6uCvMAEF2MPAHEGle9mpaeReuyNswvOQWszu6lyfFS/Dqvp28mpgAuPbYFT0PSU9Cb43DI9IF
4DGxhXtiN99ZjQMLbp7TVIqG8gIZY78F2+5ibbn6DeWJJ8wfQK4eQBr5Pp/NfRzHh4fMixafwxiW
gMvlMylEPU1ZJxMmNqOWYum6Clb0ibMjjZgQKTAWRtOK0/OAov0DLm+WEXVUtIWT/M+eI8hYOsJU
w5T1yRQYmj8RBvCjLxYOBqbTT330p/B/XV4MCTLYWHB6nHVXMffJfkXAG/jBw1KtnTNCePnL3eqv
C1KgxnimAfaxHbAfkGw0imJzGilTzem1hNpbGgn9CMHlDTIFrtwuqvOZdOky3qendOomSUjJD/k1
mvQaUeGMYuJdVYYqSZ/5RJdeZz9IZllVrnWv3vFj8bMafuREAYxBry0mYX3KXbmsbLtJX1piqtit
XTUeiYYJ/QeYvlvLIS5ZTf4czO6Oe8yvbKEWXaekZx7hRrI9jXJ0evjxP8Br0nScnzjD7S+cH0qZ
tcsuUqnGKWoOj2OVYMiH36aT0mTpFieqExUYWRfxby654QNuWP1Onh3D8dj/sTS++I65tpnXgEcn
W1rpatB5UvyAbdTRiqcjvFiX+fD5pbPZUG7O5EAh7C75MkWzIIM3hwHvBzCTn47b5jmQzL10y6Y1
h4PMTUCKEvB+IagMpxjkYk1FYU3USIfQB1rhN1W3zH8U8N48Caq2ONmwII1q158oHPHus/PMfWTJ
UARHvQMCCJ+MQI8f8uZa2ncLWK02/nEsh07ih3RIy6/IQRz2OkNSY1xzTMVmRCR0hRMpCqH6AvoV
xVRVxEond9sRu+grF2wOfh4NHfDNvVVjX2iZWaCMvlCIqRXXPwvjetzbfTlzYhHxSUG0ddtdo//i
pbJtACvGmrnbhFm7kIlUwen7xWLcGfaMNp6mFlmXgUbL/cq7JtPO7STCqEX00uoRZ8SapZh2yk+V
zIhww+7dA1uggVZR996mt4nKdZyOHSSsVgNiMBWW9l6L4nkYgPHYQ5hm/1VNip5xKoC5q6H1LKuG
5MOBErJcMMWniOcNnpKS/BLBEb7/LQRk7JN+en7r3ekKuzvRYAl1eGB2yd6SyNR4jkEZfLp6SbNA
urqQvA6f2o4Onwyy3zvSeOudxnuSLl0a/yohKODkCydpXCV6glcKkN/yCQmvbex+yfBapa0nUra3
CGhIGSbE5TuXNSgdHBEpLCnv7gnEai9R9/oeRksxS0oGZdB4JWoGAW13LjuIC7dYP1ndtHop/oJ1
UssWQG9us+/hHs4P9/m3B7uG/w0c8Lyu2tt00a06EjP9KZkPPzYSVNu5pI5Vv5uOg4n6E/jdZYNr
YxkmxFfOQsBbsrCxOIQx2wFnDXRvBwDK9lVXZG1mdLeOMTgWLVWmttSV/HPXWww8C8B3tjqvW7Rj
PA6HFj2hA9SyX0+wQ/CIv0Py5dHUg1KnDM7OYIsvRGEOjlY5bVgR5J9hlpiWBlPKHQnx6n3HQ3MN
6XKD/sZg2Fhutu8TRfBanh0q23aKHu74XrZ2WR6hRCOJn0UEG7vcMsgaVNvHss3eMKgP9IcK7QwD
Ytw0BJ9Jc6qUJLghMygIeXTbBOpd5skTuM3hYrKQet0d40B7CPBjhX9s3410EcTvspotNuosaclw
80FC9itve52rgx6tnHpfGDy+KVUYz5VtmNzIosdYS/wKzUPslrL0WzizIrU5oWl3KxWDUxObiEVm
61TVJH8fY1fjpkOQGHWfA9xVyEyEIfrOTJU1FCViJ7fe/UQDJoP6ZK8FqRvjvKZBZLzACXRE1/c3
rWz3DtgyL/co22ep4ugHNaMPQ5JOw5/Psl6FMf0yT76+vwdEiUNPMMg1FbAiNitRXgBM7R/TLxkI
9EKjBDAZneOCjkDE7G9WQoufBahjRhg51NWW39DwXN3neZkP8KCRkdzv39PpQh6hRw7CIaCG8NTg
Md3dQx0V3bl3k77HcdsMPgRtX8imacIvqaD+5p15I+Q1j9HoLI4J3KBpMNNKPgprH9pVdu0vo8f4
ij2/saKsRwDPi2jCM6t+iAOIFMxuKc8tbjJR786gGmMrQKXNtyI1P8EDesT2yE2Bv72jjFd0Ffk4
XTk2t2hFkQRPRw4gM+DoGwCTIdbB8epOI3JpdNTnOqTgL8HCKMkGLnKfRhlDkvZtrijYYKBSQWiZ
AGy2OV0tT0y6zWEbKRss96LSAUveOONyvkhBBTxcBEdPALHrMS8Sm+WRAPSASbvyKDEzEvTMWeo8
RAoRFBgRHILvUUX/NzTYvES8fVYIjsHGStqvwp7ZXYkgDJRvUI+RFa5IE4jBUsFc0EIMTzXvKstU
PeYf8g553eV+WBEGJI2anUrykBdnud+ZN+j5JZvOdLj9FXRrVn4+eoGN+YKmJ/hL812/JIDMyH+/
rYGYhVlGQF/0YTRJ+yt9MGX89PM6T47Ul3WwSgP22FEhj5Uv8AWoU3wRijBj7B6XEOC6l0dl9qXh
LFgps7mOS53PXl2KP5ZhrKwgEae/RUUizIOR7fjhvTzS5WPaEAjTQRY4U/HxQLm4TrMVj5vCdIFw
2ZzmerFXCkxsmN8yqZPU8S35pMkP5H3qI+coifqD2vzD3DTFOyhAjSlBciGI59AJdiQuAe+b8r8Y
O13far4UOcKyBqP+t6ZwpDt5GHgeceWozNUAQcoUT9fXc6XqUAGXvsSneCrsKTy9TgIY8+gs3rh7
4ettHzb4BHtz3jZGI7gGRxHPpGRCm2r87FgEpWmDQvauxXKgnkibNd+EzWZ4qMUGCidMgAbNB5Tv
7nH5qjeLg3wqwHSA4YUMGAWofLwmexHEkv6lKh2UFWCEAjW2HDMg5Fox27u1apnPPpIs/SjzsDYn
GpoXf84MIiVLNgfgNf+cpFrys3KRJWN2Vn2YySXKe/4JcrzrDN0Z4e8d5oIH4g8JmiC9dVMmKYS7
7ganL9NRVVhGbKx4z5s9lkSZ6riXdwWXGYWKHgox7vckoZT0qlX+n5x+nZCjf2tUko8tJg9YkUh6
I/asAW9EDBceyHUCeXcW/TDcMykfi9LaPKX3Pw7dYvA69SflWoiRB1IO2cgGgd7XfNjDQtBAp+2Z
QGZzBN4+kBRIBgqzCYRv04chu1FSsVgy6u2XGAmrXnkpp57Q8FkihWyk1rzIixZaEn/RjaYFs/kr
+e19MyXlrsw7NVnAlB1tqrddFBjkgPHw9UbUdWqSU5tIY3o27O8n0TDnklOv6eVAszTm3kyW4Fry
jTVJSdqeCv7mBn8zkQLuYPQTqrlNjU1mwuZbGvGEOSTm8OO7HJx8AgrBtcVShWT4SkmhSvZyHll2
FpX1cBh+DWssenZHSVD7Ya/HIsuTYqPS19Vp22kUtqWDQR1SKWaB2RRHRK7QlmGBp5bTuCLtilTl
fhdIMBu4z+LC3wZzEJiAEc/2+rZGCnjDBqzh2poVIeIWnbOSVLcRTkEp3m8N2Uu+1AAx11wG8uQ6
egb5J+8IGLykcea9Ul/BibxmL5o9uNDrg7oMqc3wNdKghhQLPFOeMfb5gXkgnMvdqlj1nNfLbPTY
5IFvvC2mHH4idaYIhZ+6s1gWl7FjHDzdbSPfkS1E52NW/5w+kTedj/CeYNX8u5N2zUi4v+HZDSXk
tApEhR32JbwpQcn183/azzQAdVjpOroUdJrDAEFFDiS+9d3GAm9AHEJ6MyLkfaKt5J7jEFr2kaqx
S9PkPe2bqFWJky3Ht2A64eW79o4kWT5an46j3X2Jl+8AvPYxqCs20aH/e61kx05M3+Dh03yHgiQ3
LOSFoMvs/GmCT6AeMwGhxEnoO50cO/vsCLpBkDa2ofcYhCwNtIy8/gBt6sHxhI/EnZ1YsxKC91YD
GS8XH+bXWJAvSyOJ0g79Ek6xngXVV54Yir1KA3E4ReYAuRPHoetYBQx/hCMLFjCqhJG3dve6Lc1n
O9dO5G7//utrAzmlOawGcmUS2oLT5Ko6GeRioCKxCnZlgVd7t1kmeSfya0MDSFdfIOCLUAMGJg1B
n+P9t1UtfGC8wfPODdcZh4RReUp+8uvxErLuS+OfOJEe5+8zYKilppikNbfh3BlaNceztsj8++36
FeKE7VbCiPIg2bglGyTfgV6cjqbu9+BMqr3n0WNAd8WAUbA5fOb55z5/5AtmQweSbYlRE6oHv0Ra
o0kvkSio0A4zBobn0WhkeB1vBdNlZvpvEleYSQYW9TZvfqA/mJKuUfdjemdwkEkzGDHLBmNg4gQO
lKwvoLQRzhKzKaZZXcOTmheW7fY5wOucazK4+g7DdlrgIY6v/seVQOeRHuTTtXtwB19hNeyEVVxo
vzJE1rYfkA3FlukvaDbvHzPIeeUoS7517DikuylY4Nx7Syp8ahqqN0Qn7Ve6J7EMT6jcC//Vu4UQ
QSXZaUvDis6jve12pb04Y7AW2LpAjlO9cFoWnd0QU5htSHcYBHPRBvj2SkJ3YYswGA5/dfip0QVa
v5jWeETcVJTvfK/xy17yej5/SjAhNtfCzSaWWc8OBsVsW+xTiG/MZAYgKfJrUCERfgBsOxtXKwPZ
60WnOLHg/DGboKaG5Vxnn5ThIddohkegkETTzEkxR54N7aiqAoL5XbUZqwXsqVLS1V5YHNAJjQSn
3OPKWYMENPZD+/NiwpHSEA0bDRi8jDyvjb9ZqnSVraE5jxH2wk/rQXIY+CoTlgL+t+a/RDwbdYok
empCvOGjPnxop4hyQJfD25YaQVbUnmH9us10w9Zp9VjOir5f1ommuvQ7n1GGyiaaqQapp72+u5Vo
smaamcp1Nzvu6ryUSU/M/ze2eGgQ9efaqr7Q1woHLn2raC0zkBhd9tp109n47K/ZyiGeLarsw8v7
LsAS7NSFyFK+jFORFM8va2bicG/Ai4KVklyDaC0beoaske+uY+5zvz2GVOOA2T0PcYtH5t3DJm9E
vWDGDzNvGSHit5PhSg764OCMfmlpwINpllilyrBzUmavYcln1SMmxAjK8w5xuWq02URdY94Ap4XB
SEm5M6ydZoJmUmp/SYWQ1Jl5ODD6NN07vKnPY+6G8fmb6JQSgcWQwaR4OCMnrcyznTNgS6gcXKxM
mILkFSdKpXrTTRTFZt9Cowi9jnSS95Pdi+5YbMqT0Ip8yOBHv23XFh1gTiZWfsUlj477yN+Yjp/S
9l8WcHzB7iDW9CqYvJSzOu26vLZTbM2xKyeLr56Ue4futGZK6ytdWsWLX1A4Nn6U+sRjDUIzQpzg
QN5CLK/WNolmycGTVcuE4ieJiBXThChhB+D1aMfBcCQziWRJW8HvnEvwCrhOcdY0JTrmxOB6GxzD
+VaIiCqenGLKb35LJ+buhnupye1hDrPFOZKvZN/5gQRbYwPJ+2XSJ509D3C2nUMalA5Fs6U4+bU0
taAVYETY29dhNRmPQOReXMep6p1bUX+VMBs5eB/AuU3axmZyluiWBeOPClPvjYWNTe84q+NYleFS
+6YD4Gr93tfa0mACDEVNhCuSiCUSSa44IVnufVLUMR8hsXERJ6yDLULiTOTlfjjsEz7QqVS/Qmwx
sg1t+4OxHT/aUQJd3P3m4v4lkMBlEhCE1kdSnvGEWliU8xkKCN0IZMhA1wCmuwLz86OHzI2mcww2
za5HZf95b+OY0D8CliNvK9Ieu+rnT6D7R4PrjCj6iix+TBEHr96+0HIKQwJIV43+mxdGonEUptLK
ZlW4IQ/pQ6dZxM5+fRueMSt8rfZByyF/LfG6udZ9ay0v+qQxHyNSy2tlJd4m90VVfG6VbsN2UTbR
fS3RzVcSefP/x1C+PtuIvFP04BDe+WtpkimffdE/3ZAn4FvyDj+3PkR1tdn9OVASRdk9qAitgV1F
vgwyk2lY+k8ZmHSk0bxQ8lnx3xtLynGFelP8LBuv8tWj4QTQTFAIxtJmAD+BXct9HPYKj7/7ePMH
KbopT1SI7d8a9ILQ8SU1rKwie8bUmea31OZsQFsLpdAvBkOyjpG5DTRU5JY6dE7X632AhCFOaDRC
wvWpxhhAdWdUYtSYnGOfgxW5FmwKBT2kYanFbhyd+SHchEOLiG/HxGAVcJg7iNOS/yHnJFCuDLEB
hJmjpMHEQJS2BxnQgoLIUrsimJ/RC7ngAr+E9X8Dh5YG1B0NHRzKxJjQjCRiKLapN2mehR/YzQsi
QxkP2Wf/6RNWAKPV4JJimbU1VqPuuAaZWwPDNGXLBhrCztjcvW1PmcrG5fj9dPkk9w8vXfD4h/Ym
+qhzuORZhfoKsT2IUvUY9MGVMc0EIq8WrDNTtaWPCtJn34IJUF4VrMUZvwKWcV5EymYwnFY/u1a8
i30nPP6+9iBY9eYaHgCd1aRcabixr9ip6KV+yyEn5TNS6hU3znUf59YH3YRm//qZ2M8vTyGt3Qfh
Q3yrq3wliQ1Q2tmAXBy74gldPcN8yFN+HrYdw5j8JahrgJDUyDfNvLZR4cllT5sMLOZVuLTq59gI
+9rv9fXdFJILLldcyz/cXnqe8pQBaOb/+IOfd/Robb0jtmFWmZ0CU7GpXhCog/75XD+KP26k71zQ
xFcjU5LuDNwkBD+YerI5+EGTwEoyiGW0nakBiLS0hvm+doeAiGE8gW8hC0NwBBWCXaZB5qFfg5y0
vDnUQkn1yuc27lEaXt5eH6pye8L+zdg08xcXgE1NNv78P1XFTm+L2EId8aZM5//bb7Q8G5olte3a
8amOQ1SALUW65saLZrqcP+Jq2FtwyPDzMQXMUfJ67mViY0RDzwQ8hg3Ca6g3IovzynQ1vdy5vu9k
sXUWWXoztTGDNlqSOKTOKG7ubG9m18SP0+U1gSG4672A9PVC1e6KR/QPEKrVXjjKrpSlvjEkjdLb
bwZ26q3jJ6HFejJE8fqkPWcn5BevyHrNsPAApjQWVp8ISnueKGcuGlRGZif0JFQGWiJ+7qnA+nWm
0DhVqclkPh8SjYCSsnbjU7Q8AQSr2yKKk7lH/3Rrb74AyhU2+qZLCYqDpEncp2rGixRweZfCLOHD
seJqWcSfKBirb7csTQZOCtnbUsy1aUhm50dWLPGZNuDl8bI3cOK6ZLQjeolvi8aAjCMBhme7g0sS
ka3s4V9VupyO4jO1J+UrzRTZZVcscZqR5I04JO0RUSUhtv50xf9ZDHkANPHl7OU8KOvMkyrR6gVe
YP9sb7ghoBc+CKlNa+O9i21/NZtCIeD5Yl3B9ym5V7ETFeibZRE0FLQ41e2aQfpD6li39UgjYgKT
WdTHFkPF6EeMEuIscp1tB5zymp59jeWeJPrPrXqeZlduWS+x4+gykKI6NZ7P/0kodtyqvUh/rJRX
wi5S+Z+/8FgsujRzkdIAShMiJyIvZwd2tpwJopWfoNj0F0yGL/KOGJ5NuNbZyNBS67olQaUAWonZ
OXfGtVKZnplBQGVBYkP+TidIUhXoosHf8YKctowwrqWXKITuArrOBCGsSLyvtOBa5iX0qF+BsonH
hQQlpNq7oORFmEGeC8dn3Y7NW6YEYDupDfTQQPBRn/8qDjWPhtxWg+qqRmN025G+QD0U0XkOARly
fX7nGWNLfMfhUqbbSSElXJ01d2EmNhUgrHXYVT/IM38p/vUxQeDjerKs0g4Y8xSJd5UraKula2ZX
ZMuc7aey+HZXMDPxVfSKvUYEMyg12SC7PkKjc+8MySH/nUjwqFfhuJx4+rEqztFx2ho6s70rdsER
wt2tzca7FiTIsebQZ0DS6eah/FOazvSXy43JD3usaxA/5WKVxdNUJBikkhhOa6SsRonmj6SbbPGG
aZOJxT+JrSL6A5L7/V+RwcuVjPW3naslPR4iwNT/qBRphsCggy62myfVAauRGu+35X2UXMbS7U7H
Pai1DQVO7HPdgKklSNsSMNlc0loOP0HtdmJBpaBsGIGN6Dt6WXo0TMDTBGDab9WK9rF/qUnaTizj
wv33LNvOP0VRX8w9innup1QXIedRnYMkCxTm2MEMM9NUWUFRqz9w7cAk4nh7UNXwy0kBU7k8VGMH
e2vMFXKf2gHBf+vqk3VUXgCdC2rX4+pPFpLkWM3ionF/wEZGaflyitQpb2xW/tm3JClEDcgGmAeF
88mlQopYwHhLSlq7YHu6sGWeWsvDVS0ssFAfxyVONc5kVG6K58c0N0u7WSWdRJKAsrfVSAI+YSYh
PZLhMqXrlioKgGYkT41IG6z21oqOyXqksK7u9RHt40ujEip9gkFTcVlEGahIObNoFusaFFibweXs
cjW/uGJfpouHt5WaZ6yz9Pr3ffTvK9jHnFxlW0SgcCIo+SdMufuaDjjy0E0b5ZzdRMRtacHrZFBt
BbRbyVWCxrXBgpe2rlBG1qIB/sd/ngff5nwoq54hUC5PNpCYsev2Z87+sZy0rufC0MzA4St51juS
FPgVPDlYIPuIUKrkEqKeum474usCIKMAkGGK1uD1wIjo9u5oeeoOtt1ElbnaeuN+xrDOASquNneY
Tko2DfVsXcuCaULH1ZPju0mBP6eYpj/x5oJTk3iKOCfIB9969ps4wB4Nhx0YUNNIYrKPdrByDWOQ
as5CLL9WIshxIIlsedgIZKxSkCxwBxfvXyRmcKS8QEsEOTui9lL3vegkP9+XWAx+XMKHUVaFVGPN
kj9b/tfyzeXZx7/DsHaq84OvJVZaksILL+dTdPLS9fK/idBtzFkbY9NoYH9Fbge19rWNXjazSash
AuVObuwVBmHA69QQAw+Fcosa1fZADpZFaSf3NHP7ZJFKQX/eLRfpfYVyuzflJH9ZuH3BZrSNHakm
bRv9Rb6bKk+nhopn3MHuVpdwjyF106ZtnRUAbIA266e/5Ww3aB3RQkybs3rL2qcsNLmYZHrSygZX
8HFSTWeA1XFaxcxbKZNmG3LNWDvR5AKd/QTfYaUVI4TwNn7g3NNPPkW2sigRgv9+kwXpcBhXlClR
CY4eXVzsp9GIm/J4Kq463w4aFuJkQn+qAI2QVx42OK8b0gQZ60HbYq3KEohqPdgo2lETAmEPLWhW
kbaQIPFgsPDe8vkCNOSNyRDc+crE8hKZuQUiMyLE70isSXjDzweQ6xJTFJkd3ldF8dZcssRLq4Es
Lyzu1GDDsQJ95jnzy/yX0e5vSNZxDmSwgdpMXlQMHtu0W5Nk0CnFC0pAR0EfZEAXbODc4jxJRbCb
NtI8kvVc2kEuD6pFjHkXgEgiCrZi71hhrBJ/9Tt7WRpfjRgIiST5JXnY1GAG9r39k2ZxgcF9Rw/M
+eFe0aobMaz6jOpJr55rCxT/ttR+F55BhJT9TicHTrGeEUnv15quMS/yS4jZUosk35SWJM99L0R3
o+XnMn/Zpsm7mPsrHWPyC4pNzPlt2dxxdH8MSFXXNSgZRN+iFUcr3ccUtkMy5w7QOv/PiIN53TR5
Yp6oKc+kjXpSx1TACCrYvtBlRH045TIgmQdTgOF4AcDjbnvKnLsVL2T66Tbryab5/iEMFF5jS+gW
9aHmqLVyExoE8LLtSCvEO3drOKQZdiozcUZd8iCrf0BvfWAEVS85/t8OeZqaXqklG6Hz8tupL28x
eJLE/z7eJU6wwY4LgCxfAnyJDhEp1V3u4Nl/v9ISchprv8a9PSquMCCjHBho8FnxvN4HE9HYprmE
ZZof5K0C2vjTqCulrC+duQTzM5JNp0KZBaaCE8WxDLiIpMmXcTjrjP9zZx50F3Wu0AXl2sOaAOBw
STKPxl4VknNRtJI8HmvD2eR5h4l3TMDmPd7i9S5nqKAyd91GNqrjgWP20LkSAG5xPBF4lAevSlet
DGogWjKntDw8tEFDSvXQ2Bnt8OeWH/rbAdBoiNk+EmxecS+5wFQuVXYfWfhZJPgZYaoh3B5tfJyB
2nJymPevtwE8O4YPAcl/19JQCb4j6DOzvbAgWlIQlwPnyI4tCPY4pu00QoI6NgTyIok4JtLXo6U5
BcUX5koeYXErwT2mp0gqQxViXhxECRVL/btpgFkcTCVEesNZ+vRq+XhkZ1dSWOQBTy2VvzbDyzj3
E88ISrWYCWe7O6d3NnTzP/jItlj0/ivF4cx3dJMPyAnrvYQzSIOH35hUTY6j9jx7yYSFQMM/42hG
+uwN2IKwlD/pLTp8T3KbMNCHSfQdeN+CrAucViropsZxMLbRINMzacFnBMVr+OBWCp9dGmuePpjW
ZGfJhQdh1wmB085FLRfKdXB6iF1yXV7uO2AFWVUeekBTWyjRB/zLLUJXbJSKxYOf6P/KG+H+IWUU
78AzJ4raywDHyZnTfiEA7hUGKaz4061tBcvzOAvm8VJvdMnxLdTpdIFP6sTjEO36AbF/AJw43Wgv
am2ApWdACXm8UphUpvfoiX1NLCveWOLOXLFX15KNiOsmHEwR+VIwNTQyY5ehz+E5VvTeQ5quJkz6
ITS35FO/DzmwjpGd1TWzuDI12fYFP6/nRdo/lPIBxRoh/oB2g+CFFRHq/wRjWW2GlSquRvPUqGlj
ZvdQrwm/pRmWd407Mdl4u0pphVei+RV6QPJocS69fVGHS79XwnXq0ueArO+GmDkMb+VBTB52NuiJ
0cm+MNYSq+UL01ot8wQHJaM7v1cxHiKCokBHqUSE9w/AMWOoYelYjWC7F459VCmNmiuhWkQdfmGb
ZVSxPmn065TwoSmGnNOBNnYTP0K9VsG8/zMIhUjKQ51ZHEVLGsVwiLjMEtxLJ+S16h0R77HTdB/s
PjOLNK164XomBFrt0Hqg0alv9TAnS5aw62mREy+m80HAhYN3X6XN+RhRk1g+XHmkJTaORFDeMecW
NfB10hfCB/Rsc8pWWorD0CQtQPOZtq5txx6pMIZ3CzvN/ZZlEj3J0POKw3SWVS9KZwrOUp44vzj8
KOqA2bI2PYPGZ5/K9R3LjXTrWUhO0Mn0LQwpxAMNVLWVHCaU7EZ2TQOWaYnPZY4BFIrl6NyOFZ9U
iIabZvw5/JSWF0xmIBE0z/nGZZom1i4iKbXodUkF3DGC3bNvXNfvkaV9+3K7R/uOXRyZ5dFnc6Xv
Dr+yjEPBrerl9JyJE5y0xWHBhAk6PSjE1pTOrAlTbMtzyEeXcfCQh9ojP31EGN6lIqMvwrXFZ1uK
WsascOhsnjkEEHT6gKVL+/K9wMnggW1AJG9VRHE6Xopu6U1qrxNS4QK3PfD0VsSp4FVZ6oErAbKG
yj69TxsCcXCQgrP4AKvJgF0eTdV23ASd/98jU7kbIifRrmoqMMGPmJT/n/MVOyH4Kossqil47hKt
JK2YBgmr/vXmqwIAp+dNd5AUGtdzKH2fsTeOgmLcMkQIQE5NxdwwSpUA1IpfRj2m1kSV/xL+vLOB
IVkVF0g9OU0chfbRrdX44LeaK0HJnPbmlXxzOdvSV+ZRxRLrQzOfskw8UWg7IpP/PjiX1ngAh0XD
FJtigqjfk+HHrvHeHzdlCLfAux7X7ZtSgVwkA24F44KcnhbPCQ/chxsjEFwHQE6lnghSfy3qBnED
/WSK7K3E5pu7yCY0s1ZAWnwaT5yewP2j07P6ocf4rd8C5a9GnpWT90SKuh4EUHVXKxweIFlGOSxl
5xA8NBINUaMVUYUzyyZFqjQl7qVn9Q7PMIzf0GYrjTx/DG+GTlgqV9weWju3anMH+pRPqBocOV0/
xCfxJr8ddZQB2iK6GjSq3cc6gHN8sQeJcWp0y96io9OHLpbqJicMBTrv3joN2v16UrieYKM22tNn
TdOOwxBvKIOZ4yGfhGSpkRw9sHehcX1OHrBux+gBgyW1mLkPWPwvw7rebiZuti6l1x13G+DP/s1y
vCYKnPM0seW52w9oRoshGZnXm4ty3XX8iSwyuwcBrxhBkdgJEcjR09XdKhj8y0ZChtgVl+ryNEZj
XTvY9bxB7lCM27HROameMcMxBvXk2Ed6/ZSLKaHdlqfFXVkufORNZdIBxLTAYOXug2DuYDALHKPc
679xUd6FSbiCY16M+eLwQRU9qwePy0Ez9kM/ERbxpVNQrUuUGY/Wr87i7Sjjy01ltFH+UjLMXH+K
KRDopYrqT1BlBRQ2/zcWea5gSIt6yDmYd1T1MjxNfuknd0Pkchq7+bdA7weqOzkUElFUKaPGDNXp
CRQnw9cBEfgPyNHdhHZ3Mernt4qxFa3EFz4gzEv1g29wUKOvmNcH5fQh8zJQkJX6IbiryVo2RrtH
UKdKmIzRIpC5usMoysfQcFl90aqBVA8Og62LNkP9Iz9jYAU8gtHk/J2esunewESPrumpF46Ag6d1
TYue1uLQIf8pbOz1wn7xM/N6C2JQhZr2U7oAzi/SAqjnATns37+Yl7/IzO0isaVU0K/gPD45113X
Kf6BfpohV0YICPSCKDFlvvTChsbS4XyThE3ADkCqyhP19ZwyQNraWowA6oAj9XbwoullkiUb7TpY
lE4OeaOcqJADRf9Kh8MR4NJv7Ku3t/wmVuiw5aNSXJAsePu0VzpCvjOwWzhktJRGszjWUEQJc87Z
r5TQ5BMvUpQimeXE11a/e2BBabdf0j/LnlL/mc76fbYhJk5aZVw6a4vmLiplqqmkEaomdPTfx2Cm
ZFR8p2xyKwYZwDYaZJr+Axa0OaBZcUosyD+UvN8jv/UmTcIhhWWWFk2viXHM18es8hxiU2xV/BrT
ViDS1WmQQr8IAQpvFNU2TUVDqU1EnyTQSy/a+tezTOI/Rmyscx3fgBhe3+oD6EnNhU0YH5hqbM8u
BPlo7iXAQtSm3M1Yp7qU4v8fi87YzCV1WBcOCiLDMYDLt+fXaFuPWkoA+29RdocowMBnYy6Gwxr5
pfvKZxmDwxIye77Xwf4yYC9hmVgBVVftIwsObaI1gONMljwfnVLJqlgC3S1QJSaCpbjMGWH/yJ0Y
6TxtMJ5zcZ3zhhBuT9JXQ8ajFLFbV1ueEgQCxP2NzgcQyLdHkIz4l94RVI1ynnvM93dTBWsABOEm
3w0DeYTYk1Zc1Ux+EZa24lMIPS4G7BXJr7i2x/7T5JUPbWMpS81lNN7LDVJTH+Gytniz1QeDAxOV
Xser3dxkfva879W5HDTFasqOZqV1DsQa5nUdHH0MMX6O4PEbGw+diX0ZF4UfjG55a9yzoqAZYY3R
Fh5sAShB4My0oG5Yl2CqFgFo6UDCrSMLtRTMAPilP2FAWmoDwaFqNJW9W+OoCwKOwxmrsAd0i4dk
LZh3XwhZYMFxs222Xxkcr/1t09wwjWsSP7cLjsQrgALjEkrkApa0lvQNEXHf6JQ9lDgQN1161mQ6
NxsDTG18liUhK5dpGDarlOv3K7qO/lt7UXedBfxH2SPcrpoXh6b5gzw6J0EMdLkrYqQDXxZ23uLf
L8wBGFDCDsZiSMR3Jg8gws5YbSr/6LWDHEPiG+Puk57CK0wksdZFhFkUv27WzKcJ7gFRrqtNZz8g
oVUUfcvPrJuvwJRXiMPCJFb3agwBFq1Xoynb66qdWdk1NzamOVSFVed29HQ/jOGGelnv4zAQHeKQ
4Sz1vayOEYN54sgdeSkZBXCvf3HV8Xj0sQD/S3FAguvTvJ6Lw2lYOjhJxvfrII7Xd7QmYgLFQoHG
ijIFZusAsZ9aNs7Q/T48b04Qi46TMpBeEPLPSr7oaIDg2QmDGAloMPfNKtE6/du64sMDTVksoea7
GFn7JK+OOnvCqFN5JncvMgq85jCYm59Jeajm2G8cy5yxYHj79q+OYB/tGWFQziQbkOzV72tcRz++
qznVDY0zqtb76lah2pkv0HPlJzvcIhCi+LfeP4RA6NhhYbmUonyqoOeNqTveex3cn9s/yXNGxLTL
jxZV0cGiRMBtvrqTsv6SzeO4iEBoDwNCl1vuD0+Y9AGNtEE1GHObVw2TkK0iLARU7YRSZ7zWKSUu
SzWI3IzRs/MXCji7CCRSq1sHdOxDAXQKzrbOFqw2fABuMo788eZqiFeTyH8kKwS4mVP34OY3DrZc
+ctAIZCCuZjcWhRD30PYe7HF2Ee0cioecXFxt5CtIwaR2W1zO/rcHOYvEyAhPSCP1OE6Q2ILWelh
44jLk0IugQ97RZxHZ1kxuotXDx1ILjA17FoTno1XG3LvCiN6SMvTSNEuSSszBnvMIt3OafUcvhYv
k86+7v3BCtBybREP7O3ZrrUj2+wKBG0L1uE+gS0iKW7m5CXsGwziLEHMMguyGbJjw3ZuGGyn3/Ah
h1wL+9Apoob+S/5IJrS4954CP77Q4wadWlr3leJVomFFe7N3wS8fJscaCnGimVYQcEKBUIeuUZL4
ippgPJXtc6Ih+lgeIlPlvYcowOofl9+ebQq4kuPUjQFWweBM9v3Loyi018jIuLO3btCzM3euvoWX
Wr4nsX4e5bjnKUx1HBRaIYdWRnmvA8jn27ujr+TRn15OX0n7v+euSy5BrK5EyePvryK8xI+gDLAI
zjF0ryZ9tgvYBfC1lT0vsX/IQoOPhAF2pMGnCwFbWzYJifOq9G6oOsb+j21tHd1BSz3Tzqlp8XLg
AuIohknr4OmmDjWKFAAzlElSoEsgxa5ZWmhqC8JBat4PazeHk2b0X8WuvksJX50OxsigMG5Ae8Nt
maDanPyKS8lN7obrNxKaMfw4jq6k+ccrnWpA/CQfAJOO16gDfImpyhMwXHd7IicIZCmjrY7vGBWH
A2Y+aCFsQkV9PahtyQqg24yg3RONPsAPJidXM4xGDtfeTLMf1EidtWNsG2MYh8IzpCTX9QyPedc6
y52vghRkK9juG40xmAtRz1gr7tQ4Ow+kAe5h0pUEhOyXa7DBQyQQQp+8TKo+PF35w8aKk4YYupz7
YtDD4RYNGGIBKPb3KhGJy4+hRlbOBW4ajyaLQMzQVM+8MhoV6eUNulmoZsdP4L5cPzpXFC+fW9JC
BFO06aK7y3u9hAIRQOtjZpYSxXIT9plVTeuek29f9MwzZtxhbXxiZhuPMuxb21413fL3FiVAVE5B
3vMAcnimsUC3GDKdgSNN+4MLs/B6j59YJEXHfvNakBqusWhcxqq8B+vAvKniJadNRlWbKeqdFuCP
raiPk0x7JvV9u8GmqXd+z7jdq12UAgF7JWxLe5IAQs0t9cnhEumWcSDVTkuDUqoevFMMPnd3+MJ6
aT4BbXbg2a7EFWEb+UMTElc4CsdjpccUS7F4Dd3+JnEPvoIIyW1ZOr0mXDeonKxGxaUdlSkAhMgA
gTYZManTvAbjRoLVceZrteiwlEOlLtvvpnWods5BFRT/UNc3uJvJ8Lrp28HSa3QE+IXRODd6Ox0n
7aPaGoXxYkLo+PpzIErqpwW7oBmtGMTmB7ku5F0xHtiiQH1STR3jmDj4bLnjBwJanjaX9MzCuVAw
hK+p2UiGBrNpZoshg78mbQfZsfNMPtBMCr0SUOmV34irqrbkPxGAA82po9FNQ/4KVZbRsYJhXhD7
Rzg8sqVlEZKKXSmO9oXbOLna5/ow/4gs9DbkYyFxFn9q2ktEhE1qPzNwq9ubz0DMO6ZBP5mZEC6I
v3wgzeEshUDBnICLjRc4QnE2fRhFXHS9yhiB/d3BkXDudpbFQmluuuWR8v4w/4T1rqyqPZdEdMpw
LV7kfC5eVnGy0JriZLJqaQoA/iRBZGmeCs8AXD0+9Vs2qN5gIM6J8UZ925GoNr4byuJkFeWR+2kc
EuqAcNHi8AwZHPUU7y2zI5e/XAbLXQAzzkbsY2gXavMpjCnGDe7PWJwhDUQ+jYNh6P97LjxUwd/b
THaQSwR33UR4tDVzUCnhU1I32YL8Tnf02soLiZN4bpqcLpF6WEJ2K0bLIsG+dBzBMCoNEw7oArfq
tWxW3kyQqqOGbyEfin2x2RkA+jk+Bdl/tihpW06ti2NAO1Tqao9gxg5l66L0Pw3RewCpioqPlALT
i06pF4xir6aKa5JVfMeK6Gi6S1NjX2n4StGXp2U4aVhIZ+OYJKh3PvfxI8cwCZGqf6+6CgAFeEin
IPumfu2Y6mjXnI0K4v8Zj/tLJOkAtXpA2oOj9gXi50xKR6RliqdAFet2kEW/I5iIi6h9wlVcnQSf
6ETWVZAGrvcKRgo3OmqoNp7OvHKUfrzpi6ID2QwTxl5uvZkOddT00x/+Hd7SNLTafrniezM6g/LH
7ST70M1V2uBvT6QZZd37WdFhhdIrW53FsRaFF6pjv0HgroCSzIfZovE0CjHJQIIw36qVz4GWoxnM
NZLRyVNA8wYBxmmpdzX7dfI2wXZj8bLSMgiNk+VNJ2PKgttNlIcBqa5B2SipGrrckL14/lFp0K/7
N+yR1hTp6jueZnQZMVeiaK/fBroyDyrKAbeGlhxoWL79woVXTUl93yTWNDihIoMYv5V20j7ktpEf
T3H7c6jzISuv/BSOlKIAbL3cle5CddW8dH1OT7YeuIaf3ZMk5tSTcv5I+v7c6pG3SNjsq2NsNejN
YGUtfb2KB1MumvIPtHGEBe0TzxmBJs+pJK0zIqNWqbCg73XbWu9jKkYS4fXWZxk+0n5+p9jRIcPc
gF/kwQL8rDxCBsQyrWosAVO/vF4jChVoiyTOWkq1N42K9br6XhgNt+wRLBaUFmXZ7K6ZXUNd+XnD
NOx957MjUmFC13gaG7cL6vcNhWEHVWnY3EQhnX0SAJEO/2Coqq6ibfwakpXgsSCvAjHhSnSTARei
lYHSb81dX/XPXbZnBjtQyYzh2Y3aM07o8NtQdALOgRk/IDnjDwDEczDKWBWC0e/MzcgJ+/xxfef+
gOZkUy2WVbeceDLFCDkJv/+4TF+fnvjmwt6QSFNthHYh6NIVK4wxSp0upkYvAlyk6qz0W6Ibf+g7
1i3gNvuZvUPyBjGl6UF6xsZVdyzwcIAkdotG5vLzuSTPRSDxPkJglErfaoAJAMhuPcnu28ZDBabN
Sq9jXiOEG4gcTOVBPG4ImOksSvDsAROaFxk2nM7nvIf7BzNvPH1pCcZfECvyDpPTYUeCwGefbf9r
DcPuSXtqsF8yy/+3uCQwe4fRVyfgC7AQE/fC4qMOdjNVKUm/wXZCPD6TrEoNG9QuTwi5fBuTo1EW
Oh3lawwXBfDySikqM0xKs7lMIylKQ3hAWyjYOceuZaxnqi+3rWWg76uvL2T2vb+1peOa5bv1KFvB
0BU03pNXi8JnqvS7/3K/38h6g5DXKdj3QxXdpdmiiAv+znDNgHkakTc+OxqfIQz8d2h67NDA2+Sl
uLCCa7NSd1nmgo/bQcH9q/dbJDngEBzozYL/Ineg7aSoVRl7upC9CfP8qnF65oHve8nrQocj8I+W
u6Gyj6LVwDN6UjEMn4kB/5/cBmM6Oi/53NLoAHdhoA5ct55t8zEwygFfA9rY2WBgydJfn+8/uycU
ZML3V0TLfXUs2R/pWDhiB7LSEUP9WJAXJbELIkqZ5G8GdtCKff+Z0NH+wxVVIjhc1O/6sweCZyIz
oB6CjSJKssSuNzKzB/XaEwv7lMAI+jQ6MKPHwdEV9ilSaea4Xy52a7tyeqW2V70NoNLMrzSQY14X
fZ4/8VyJQeoQ7SRDQJTZoJcosoKe4uQufvPs7flxZ5Eo/RGfkQveaKVQKAn9m51kHR/aVQuvwk32
n6+zWGTtdRWLSeW25F+Fj3b9Kb6pQ0WOwWjbWWFu8iZjqU/8E0L7JG1YQu6BcmFg9LLqXG6ysJCg
qXhGGwm03kM4o23GSknY3O7TdKrAMgG02FWdcxkPnx3pLJ9gYGkD6Ej3wfK6P5YW/5uAzLgouiHw
uu4L05mCDtPlbu+QzJdMOdDP9/Fhyh0cspKlhiUZITG1/CCMa6tpNMXoxHEm/48DIvM1qrajJGHa
VI7q4VG+ePETSbHS7dXPDQalKcch778yLCFOT/4rSZzpxXh6qTfVVWTK5gMCPb99t0zHqXNz42ZN
2eMJtnXaIRSjshxQtw1TMq3O5R0pTlwgaW1bZeKU4Sk+5B2pfan3DzyQrnUTYjt41SfQSmzUVag4
j69DkgfIwgc37cjv5gMD9I01SqXQKJ23lW3pvUD3YK5u+vDucNnBA6NSCoImAl26i4dkyBS2GxZx
YlUz8eOhmRRV837xkQ/wk/bXlRUKO+koC7SQsiAN3wOwdv7J+iSZ/DHQ0QLIGrT5OyZNwA00AGtx
uqBn4SaztAKT8412PGvkUd1GdAhJeu/SV5GEj7KDBmzzEjvqz0vzNsA43Kj57NHriKrDxJQfwP7s
6oqHPbhLtU99aIrW591+/SFzUr2hpuhKKbcUcTY7bgVAkeMDN79DCwPXcsIf7nrFMb8bP7CAxhL4
7/hnhrfQZV5x42z3jfYajmy3/8B+/XWTh8Thx1YwUGNnFYcBkhecz6Azu+BTEgJjsJZRX9R8v34B
Bs8GMXK+Hf9UITEj0k9LKcjlHE5G6TEL0BhqO5v0E2kvWAZe7RI09CDtdS8ZZQue0JihpUtYyq/a
ASyFe5q21X5k4R/GVOHN/WTpxZbfKJ+XYQCpsNifD5g5f7Updnyq527FKVO4tGcIVXOZ+TVkI5Ik
TK6j/QvlO4FXKwOmUIsPcbMJH23etJ6wunH58RQ6kL8/Ss7Z30oKmYtooUXoWvXWjT/FQ0yIOexT
nH4WTDKBDVrazQsbEpgp3Mi86+2gTAlnY6NscterKVxMWkz+6bu2p5JhxbnaZQ08m9y7x8Knuo29
mu5BBhZXDDys0ItInThlF4M7hxAuvkOXItRNWNIpwxZCv4THvTKx79JkcnQy7UZMaMJ3PjeSKgLk
bpsHd+px5BNwpLtiLd0Bb9J4KIzEsnzyFr4uv6hebRsYcmFGXawwqtr8THBR9vKrF3CirDHZiMxe
26sy+hlvrwiEhUoGkkhugF/QO63wNpdaRkoseDILO6bV1tGXCeU6Ao98TM20QkoYSdD7atH8WDSH
hr8SsO55uaNd34rJSWGpQtidj9YvN+ASedvyvljhMvYzl9EUpNgedMWunn0gWba9YDmh0qU2a8Yy
mh928lKTgg53xlbV+TksrJZT1eY7Rwhwa+/xjIFW5Avqa9wja61tosMgZD+oHcSuT7KXqQ2TOsAM
4wSwNXwL4BzHh+a+FiW1qMHaRCqQ8puTQn/wW8/W+XZTWzjTSYZSTpjmUXGUYWpyH1bB3/wP8Bxx
DaUBGlTWYqhZ3lt28TWJ+Z+A/JnwGnsMsS4V2MQNPVEzcrUpQlStgWhQLedrVq6vVZaSEWCmNYVX
w9jCN0k2MQZ6cCjk0Gl2DyW36xqiN84v/ttZtVZj2j7R9OfaHCKvGi0sCAmlgfOCr62IO1JAxI8e
l7FSzzHYMXirReZTWTHoeBkfHY/VxW8SzrBZOeZa0DA7pUYZ0YsiUlOD1gVAcKvxo1lHQhEnyLpk
EtJjW/tdTkhIX+BoQyogRg19UPx8K3aZDC8zdkCxI4/UcOXF7QDADbLKqrn0MpKPtwaAzEyDYW8J
9bm0Oj9uXIOuzVMAqXhGeCI/CpHONnlNsfswS2/B6pTC+NxDXvChpAOXdXl8M8Qb8GbmE4EYslZA
Bw80JGMYlIBYndPBuIFian6dUrWENM7rjuOTJR+OWVQaAVSMl9oTf52qKbgVtf+LhpNwTmC+DotV
IoyIL2a5c7k0liML7FKFdzjFK2hfO+x9UOkQt0Vq6k86ZpD7Rv75z8voDFa0638ogFqJxVOehf68
GUGZePObFcmaufr3arlWDhaM+dY5ROqyzwiIklyp45/YQr5mmN+SDc5FD45tb+NvePXBmnOcjnqw
wZRzTMFXCgvz3P/TGegBPFIDjjxKESCTAQogRwUsbdi0yKpCn9fVJ3EYTC8DI29xJ+OxCpdqOMv0
CfHm0ye+1PJbapzEncLPUMurtmmYNzZNwqZbxwzv4g55JzM7Uy6QCBT4WlAejH9Zmk7id98eXHhV
K9ASHycb7TL1B3wvAiKf8ykgluToS/dBmZWnCzOUwZjps7aMLeDuUPoKeNfTfrl+BBBXXUieODwg
ldhkyclv12cJZP1fuXTJWfHrbl7dBw98fSJqnxYXF70TQj/HjozoCDfrZ8C8W3lAhXi05JUfzlQn
KEanX9xNzzt727SF+EJyT6FxAE7dl7CgbZuyzjPpdMO+wfMk/oA4oUR57BY+z5C9iMpcDU0tV0Mm
LgzV/ZAJUx+h1I/D0QT+8drG6ioSySFITBbLhA23ayhsCLOLyeZwQtoO33MyN/J4l9M3eYLuyhRM
oTA4rpYPRqY8OqJ/ydqRyDkZ/0s6gXIIUo/pI/LkrSSy9KDi/54SB0JOM9sodJkAPES9EeXPXCwj
9btmEy0BIa1V2nazB/bSsv9GUyojMZMTTyopg/r/oMJ2aroeu+UPQh7d/25o2VVmhioXq9+XDIkZ
drx9nywiQ3IGc3VelK9LSQkOIKvP0PrQzZiSRFprjIWZbM3Gmn81PXk1nhMK4T4CAaWEcp08MmSR
Bj2UJ4RQjTx8yzTU+xo2geA39ImngfUNzt1nKDz44oamVhUVwgumMFs7HXPtLkrXviYeyQbls+yh
Uux+WL8F++6Qc0Zbqxg63YPnitBs3mte+/DuR78C14W8i/x1f3q5wNj56dOoeWeQdoX+4fy6IPLw
xYLT7x1P4EQtmmOYS9Ln+w905dK5D4l90nJj3ETEJ4o0l0LJO9p4O+Y8ZUl+DzGUpIl/+9KHjvD2
E2ly7ZX6d7LAp2tKp27ePfekc+jj1tqJ8e0B2JQlFC1Y+h/Tb4NmFGQPe/vXug6t9hhYPlzQ68uR
hbI3A7yIFm5UT4ldROqUj3/VesNGfDLwrem0eudKqBGNCewJLYVQnoqYsidQYl+uA/bDBeb4k1bt
MYun36lavMMWVa1HY2w84IP/cIQnrzuDT3P81RYU40PNsrN+WItjr1njGzABavYJPTUVSNh9H8CY
69INDWuvSUeaDm107absOEytLMWQHvOigH03HGhq63fKrWuqSrqp6VeQ8ER13J6XoIKrEpJ1Lhro
kyvrA3KOOyU+wUSK4CNySFJed822Qo5b1ALSZXaBXp2uxhSTYlscvOjjIIwAXySw/cXVTbuOaYLE
oIrNAod+evSvdrFK3t+q+vRUi4UFbT9yzdl0OvK3EPCuphlkbotqXEYRnCct08kTWxzEalapHmny
XUiW7GW5ZeT+Nhh2djL5QZh8wpParxuhSIzjBVi/t5M71ol2UK6r2oyIY5/qxzAt+p003U6Bnecn
gONYLdUKROHD6ypaKcjcBVdKNohJ06uPCbg/8+oH4LNRZnh7MhGPRQ7vTlFFVeYahdGlq+NgC9ad
U/bMZgp/eEYEs4UV0yzFpwy98scy5+0E3L1qN5pBa33gSaNUDndQJJJ5AbnxL4hPaQxVyEXpES3V
DvPU0wp6sk1tbvXyOpbv6/2sTvU4DeIABG7/aGLzFGgDwc0dGcP8SXV/XH6pL2aSITk5+9z/smsY
xFwaTO64IAE7xRySLZR6P5t05mHOccMkAxBTpXVnrr2NdqDl7AbidcXqyRiU6bNS11+2syn52R+A
cmlv+fGHVHAg4mZET5kEfgMt/CwLiMBujxf1KOL0o2wUApe0q3o6erCmZm26jdIOHUabUBqU/rIp
B1669USd9UJexXotZh8XLYkTwendBE8NOeUtyWxMZcSmXK3SE7LdvVgzzENAkoBAt38UH+uvzXw4
2oagTjYWIQb2wSdtFg+Siv0SMacm8B7A7QLr7uAPso2qvejqEfSavt+rCu5CRlk4cCJN0vid+ZxQ
qrPsVKM7ARU437qu6ujbs7GAV/G3e4nC9wGvoGA5cYaR+8tKf5TzFRh5eYFoKmeT1yaj1RbSvPCS
5r2/eeQyKYHhYUw5mBQPMx7cYNH7WqtdwYzbORUQD1YAs951kFocaIdVTtr68RdWvdGh574Uej6X
Ji82nQly7mqYtEQXXmEz2EIyOSKnP6uT7PBsW6TES8iR1bQqHFQFSdl+VFl+1TXloncgO6IuSl7W
sp4ZEFT/Y1rSZUN2Ql1dYjRm/womZNmR8Fisu15jTaTUULHQI2Ntc6+Cm9kAP8yzUpcyti/fi8C/
h/zYXTCwmBowQlK3DSyqNWBSDXgNRGCD111sDJ7SGb53DNigk+AffACBJLSxEj+u6ikiNvcujBF4
WXcUhMdYekU9FY67CaiQ/3F1YhSgRt8BwjJKNm24TK+8z5LSR7Ya1kKZ2grPSe8XnMQ9SUfVk5XA
ucoMyiJGtgJ2DeWB8UOTMF6Gbp+T/yRTwx7sp7KNNAk00zvo+/knaIcjbQdO2na+lvyMkEJM34Yg
l1caZY+OSSMG4ASEctQVFvt586StNFagFWesI/6ViCw3axbhHp8m0xIFb/mrZcfJ8KW7RWAIn6m6
zbksEEKln02Jvi1SxBDBNukRg+kDhHvryQ2lV+yqOnfOyrggHpXXVDFdvjzvxq3pu7aj0QdhZ7vV
lKCQ03hl5h6u7Qqv1ivP2a+7Uzm3niaPwuUvsrEVlXtR3qXswsWqGAxsjlHTjAQclGN5SJxF6B+Y
Amt97rmp5ilETGZDtV12nvHdYVqyBh2gUuJ4k+Q/HEglv5SuPl3IbbFIUzTKPhCYXBts9JWoy0f/
3eB8BN+h44fn5Lt3VJ0CQqS9rfZi38cangI2jrm9RsjAwU/r/mhX90Qum2gBy0FFlZD6J95KsKd1
Xs5Jegtagf4Jro7sF+wRV20zBG2v81r7vSHvIUd/puQZuXtf3izxSlxy5nyWv5zf31hAIB0/E97A
E5P58v5OjLzfCV7dcfSkLU2GZjqCd3f953G6fX+Q1vb2Z6qc5AhRmm+f77gEwPN/wPo61veF95uq
O10H7eNlTqCFnPzPFk2Y19ChriA8xrZG+PIvVbAYEEpHsUqdhOzdr5v9ZSTkdV5GrpyMpQOv13zA
x56aVdGNe30F//wm6gpGFSRXC76wJorK+DD1ZexX5Xdimbkdp2HQXpgjHoWuqLkJ8fmO0fNNZB5r
/TtcAqcUAdcJkGgFZZS79hWyu0V/eez9yDgYS2vakLK7P4VcFefb9XwpEu360xn4hKgSQzWqayN5
ek/04j52NOOiQKqQty1q7z/iSPdb58f58ji5JGaDtj4oGGDbVK/HTJfcSPLyFLUEewVjyGZuUojc
oE8KZrfyxQFjcCU89mHQHxOo9vloQLfvcyFfY3RINpJMcQJxH2xo05kZzMHMAGaLDrMaWd6Z1bDE
jhiWKIIVfS8qmnHy5LRMgfYtfCKWpm86VhxcMyt5bpLRC0SogsrbVl+LONQtw2ZwORY3KeGylntB
cnG2UN9zNcKIJWVIfs4Dwenn4rpvs4vSdaKRoY60z5kf2Adh5KRCiUaOpOZd+G5v0mx4UQ2fzG0a
Ig0s5/QeWABYBuEKKVpIlivWmXjQ1/zPVSwIafB+JAYXxlPdGEphDrVfpX6QtTDo441WgZfwT4FP
G4mADfCIeoRvihU2qXWMF13bsUf77vLpDaxL/NJ/ZHHAwMdvxe2UG2uzhHQqdLrsvBeN60pVEDED
ygHvVatNHww7xXUohDREKgB85Ph9z8hUhQUv9h50kJ0rcGi1RztyfmYTeuS5dNmrQPMTsTP/ppHt
aFvJNMdQ+rDN1vTzf4Gv0a2iw8Qe/rMd+E0jUc5YU/CR6U8u+SdAnVnTEUiPVRWay6Zddu578jL8
n01dO4zZjuRufOsxHHQ8XZN/vy/I0cGK5XZasIPN3++T7UoMCvrJC9oKuKYNFCO360W2xPVkLAFH
7zBeP4qxaFj1Hr1uLtak4T4ha3z/X9RY6h0SENOTTLwleG4iK19TL5SrnAjwk3PG+nM0lqxQRzPT
23erMaD3STBvJ8wd2CsSHlc7prfx8YpzKyh7gGNcr6fL4TBFlcFkyx8/LCFPSfmTKzzTcZCqzXpf
6m4OvjDfDapcAa3pD9ZbiU/SecyThgDmASjG/MeEBRTsJRKMBWmtOc4cCmM2Yp0hUuAWAVsmS3/Z
daElh9+MMgcjSvyYdS0jHAYQnl2Mip67hcVIRvLACzbqXNzYl/2HE1EYimM8oVk0yrCvdCySyTKr
qNty+/4aMGcINRJmZdn9ZjyNX8RDAnu5oayX/b0XBUxlJ7IdZUH/Kpsidvmc3Q7CqlDls+KbbZrh
J3OiMLM2iwJHOcn/LDGqLWwi7Sl++bmy1tDY4lVMWSqo54SbDmJLOmXMEM4Sad1qjBQQRO3bnwSm
FJIIyDgG4RgXk18zJEwlNCoFrPdEwFoKf2qhsyb2Ba9MmqcsnOjVWlHeuXtKxiJeoSDdHgIDdMjj
R1M5fWRMqHdCyAwiLLguIHRSczSE6AjbQ5WwBzY3/8N3+CRIDUge7TJg8xTw9t3ooMCHUazvtRT6
fX1flwEh2MLVdLTuYoKJ3X/IGjnkFop0AxeOVL+NeuG5WBx/5JI3Fwf4XAugcHB22+0HiMCyLOix
2eAIulYky5nVfykxHpc46lbB3KHmvsCCsj1pfLIHptgs9sjEgpismF1h0ssGGAVg92A3xGP+eMU7
9uls1K/0OmcveaNFVfQXeeitIy4K3e/ASfgd7KA93ZhJZ64e//2+VLlBc85WwIZAhZCNxP5Ydtzd
tubxxDkjb6FOnrWYN661bH08Fdq4rVBlBAVMH5AU7tBiFUJfQg+rkJzHGNWw/U4UquZ/guxXr/79
VBHagsyTSJfZrvUNv7gi11G0YaJTlqy8yCFF3ijLO/1e1atr/xg0kVg7bSI8w9UPTciaFe7ytYqN
8gD3wj4kfBfPOSZdbHPr+dbi/27/ZM75GBqDpKZassdHFEF4rcmSAA6K4Wq5mgY5FqYp3K8ZFmha
KGtPMAL34uQgojsqxnc2oxDc3jJwW60eLVR2dTfQ2pnGXtHP37+f5c2DaoBmGV4u/DJg97o0MsZd
KPSC7dNCOBthMSgJb94XK60V2jUnZSglc8af/ZJPmw7k3YhWKUbfeK+sebttcXMA9jKajmdL9Xmm
lvgtlFc4+gyQNrTsHI8H1js2xt9lBEcCLnUH+lWF1xxDBbYlquMKBlz5V9pMpP/IB6vrCyvXiYey
DvvC4XwzL16MjlRbPrJVi49c+G7v/DX7MUujQvnhQtgigo9OO9xBzZS0PXeN/3OvOzIJT5gDwZlI
D7irFHiXK7Zp/gfzOUU5OwuNl1m1XGpzvViFVU8oiVQQEBhSrMlf7E0eYQcjhaeJi9FjX2A1Lp57
2k8McSIrXBAo+JYeIJxElsFJwsswHCUTP4Mgwh1p9VzT/OO7XnBooU+KkrGm6k7GwtbVc5RTddWp
ZCMCH4mmneZdnr76lNIckig6w6lerLnu+pLeNJqkJQ6dEm3Cgmi+Adxpq270CmErQC2lfjQkEnFd
j4ExzYHlPNqv1TqdHGwZxsI/e76YlT51z0R5raudBlQ3t5D7c6YgJSSjCYsprlwM760LI5YaH3wo
FsqnWugvN3p0weTbjggkxHJswU5rDiaXoldlgmErhLCulVY5Rt91c2eI8h6nktDkPa4bgfOZ6XXL
n440VdZiO5hpubGBeWiMekeul7MrA4kdWjBUbzCpe02Oi+OuYFJnIDiitu4FHIyJetVP+uvKkVHV
yQY+VXuzpp+ObTcu6OtaIYhluzQp7MvFMJThNZvfbHwD0cK8AOMXpUQHYB8HOt1ATUIrP3pSFh1W
Pwklbwb/pciTDrAPRaa0BE0knpY9GOWk/QjAHXlDjvAP6iewgcMob5bfh9HHtmskWldmdRa9AVoo
JDxsJ2D9ujqXyBvzRBli91cyA42wCPwaRI209bQVeMUBzxopvZ2Z/pKsmSdqwjlkhvWHdJ6KZve+
MoFtid5MT39fGhaov4Mr510sr708iRx769v5nAHmBsl69OnS0FbmQJmmiDc5Zn9DHuzZ9ci/hL/O
Ywnb5NYk4ta211ih80+Du7aNnFktfuccrvcZwsKA+obBG2ZRmoW2GCd9A3FWOb4AVGtW4i1FhcLd
aFPkqKzrPQDcONFFnCUjoZ7iiTBLAXGmZa0kW83MLEcN4kpfJAFSl4T/2JC2xYlq8do5WZSNF27A
Swlnkep4gmSLrHSZkYVUY/sTJXSh8sUeBg7SIJm+i3cR/HX3+tjPx0jes2sQLiS+40XIQY5Ekr1h
dy0gbHiOLnpZHMdSjYS5xrt0LyTA2qZdfhJ+AruJFFcp16+qAjIraR+fFottmk5+/v4/0w5wCGxc
BFYhc9RFsPevfJVxsjNoT0/P4+//VAprwtCtEch7Q+B9cELYHHy6xzXLukSDeorK3Dth+DoqTzEN
kWnqWq57Yv/nTAjBIvcYAiE02LwtnLRAGm3xVhjxQDItGi215BuHyI1OUSM7hO1GikJVbu+VbT3W
In21xfuH37hc2itstM/3sZl8tRvevJmgWx0K/PHIijrtQ51svtWjLK0KPEKlOFywAed7xUwreSCM
+Gslv0HKgkSwnkmc3cgoijsBrgOMQrO7hGJt+JE1uHZnTF7ynvEkrEoHs0vFxoJFZP/MHKw3mmZi
18PGNS7bg0L6WZB9mk//VlDFtYiGpRAXvKoFnUAb4JYRb4+fIg70Zvux8P03HgjLLgwE5HcFMtcg
lfRIUyXiyhDvS+nkGO5FoTARMW9cF+6pZjMYyP9/AFtVvSuzaYiq4ow4NR26BB533ByJra1ey2/S
mC9oRjS+gjthuUvxlMaRMcLr6TLWTkoDMfz+AJJBcdkDDnLkpgTHyPgZX+ky+JHrXeOK23CYjmhB
UQ6jIfGguaewC1xsi/fZzu6v5AUf7stIly5OOFAHho3liXgD0s9broEKXgjvAYaHM71R7runiiFC
vDWflawx0JPrc/ATT3Pm6dzRkBwh8TFh6CeGkAnRpj9TO6kNG3uTbIhp6LMSMpkKDXxErlNJZN+v
BreAYZq/R2ITwcqHrRCKv/M8Fm7OJU+WJUOPEP2XrOdBpsJdhOCeu7E7687DVbexBliMsC+ewNYT
m+fQmpN4cn7gekLJDK6N7KI/nz13o2xM9FO2uLIIa8/FQdpfURcb4Ssafa+JUXUz9uDf7slvhlov
dPgH0F4/EBXheZh4s3doU+J5btPm1nn45FZWQm4ZFPjznMuttbGQii7qrk/pD0IEbTnlfZfLImDC
P6uBLnHrqoj0V5Aj9NyHiiCQW7rfHUwujVxG17Kc0PJtKq7g2ed25yUo1IwpQlxe86oz1M7HCDmV
NmG1oc7VRd95HMq35JeIN5vS1AYdtSF3Z/9/GfWC4ju5lapZ+8LNgDZXgVc56E56GLReYpkMbd1M
4urpHjLLzMaBj5Mu7PFgDbU4KPLZ5As69vI0ijWRIxNrwV7vryGZA2r8dqJOIIA/Dwz/V4xQW6yl
Qt55ySwA7iE1wjSbbezyYo3r7o5+OhGIN8uk+fon6VeboXTX1TZnnWGr406tBhpx7tf+jatM50Oq
a0ncby4LHB3oKjM8IPUdm428/91V5fPguOsC86qDtkDHOzjeDawKnlhXVGLxMWQAsEDWYAOVw9qc
jXGYF+uHJ45dnWoGTj+1xwB2jF3t0OjGXTZEzqr74pZ2INmHDbvb1dPCHaVOi190d8FFsvJz4SJk
TWls6w2wirdkEnocaw4czLpPfDq7/eP0cPFenF1C6vqnesb335/595RRZSPb+h5UaOyh9shD44/b
tT/b1vxMYLXtnSv+H6w8lOkByq8ErG6Da5DD3GMEaTsHabfpIZfaJXvBWiuEr3WgE4KOWKwHOPkX
UbGP/mjECpPQSCpfXM+ReEv/uVE3WXB8FKoxYPPNr9hmOHTUBh9UfC7R+GnerNC+Cfoudz1R8fck
11eKj7xMkZ0mE8/43rCeq3xhKPAMrx1fgBwMMU/P5TsLVLqNm5MlBm40h1wMj2V6XZWSaF4C0dxN
zJJN3wwKnAEO4HAa9uxksFoGFIJzIh1tWdRIXWayUQmXO4txdvsiEQO+Oe4+hnnHa2EwoiDEO7pL
W70oovin2ogVjAtO2bEjiyKKqtmUZUYGC8CdVWOdIvEWUZiwW7XToceylmwZglYq3tRrJqocajRx
5UtggifEpFAlnFwEojfbRc1l/8HVO1PGc3p+EL8y4UFcaZOfV5SimA5a1PuxVhyI/oD3qYaZ0Rvn
xnzjoggDbxIXgAsKJQelbXOpV5QEMP1IMqXN7R/RriGnMzfdVMWtK7uPz4UfibjSosluTRBcr5gA
izTRAX95elg5Xb44lQ4KxOwoHFqIhtNlDOCSaIdd6S/VuvC4ZLwcXA4x0DFL2Ens113Ix8KsDn+G
MzSuwIOCafkzKR8CsaTMsUkVgwqnUbwW+fPIjn2p+LdVw6ERHccexuh1imLfGwT/vA/uIG6IwlpE
620VazKLq6fFw6fLOoepB7aedeGUT+Ab/2s875dJ7N3mBbOgIxi87BYhQu+PT74AM51PQkOuKcQY
Qgyxxg1gc58/rPij1EGXqEJ/VCYSUnS2al8uVNuOBXf1I8F3DiiEGQMMG36b6xbGtaLRlT8BPApY
rgU2S81wzYoF9QVWeUJmUmhnN0Yt0uVOrnr3GcMdt+KMe37cQy2LBaRICeNS/gMjg63CQw7y76dx
7TyO4ud0i7tZsSCtmk/l6DYCSVCw06Aij4W9xCQE59ybVV9eRQ4JxwDqYsqk3hg3aIq/9XZoKlHw
im++zCSS2OA/ITXDWEtjWWQYZX4AaIO8ajZYpBwMHELNiDPWUFXdzPSeT6spMoIEeH8Nd9KUNxS/
6Me/nehgXhAJgwqlu11/6IgALlTEsxppZ6tVbXYfESmGGZv6c3yJg1Xa8xKF0EO551GpeOJOJol3
O8dJ113PjEE8FbIORiZ7AlTlBs9N6aF8f0vBYCPmTlvXqh+safi3Qae2OrFRrUqaQ0AvGneK+OCE
G9oIwjeIzNkKxpusXEsL66204H/szY2Q9STxdLhVfe8DBclU1uP3WQOO+0lUzuplEhJ8pzaJogXd
UQ2s8sNUrbSQ7nV5DceaZGA4kG/28hGQB1mXa4InsG8jwGlzz/cOfm7FaVX+K/AitRzFAKmbpOKV
vdR9GYUwW9l7nh9HvzudRC9pln0nzkuZ4AucPrT+6I9SB54gbMrQQ4AtcCQyVcHtwuVbYVfFxIDV
svOYG3KWSft8NcmJYnH1CBOeDlk+qORm9KtukEg+1pdq4PTAeJpFLSXRyaD1hLiLb7aPikOII6J8
zdZQ8dUURwFmXCeQFaF99icHdo2DHuxC+wLrqSrjG5eCwNmTbP5VqD2x4XkIvWmp11gOYXoq4dIm
gAJxqXgRbag0m6poVGMRVx0D0dPXogvDZgTMH49L+voAqaLhrXgaPZ3e4Ng6izkJkd4bHYKbUwqu
X5Ylt6oezmPcHT2XYY4EELJNG/dtR44R1eh2EpN6P1VbiTP0N/hrZcITqd9tHluWrUTp//j+ub3Q
+FOCQnxkwmIwa38UaNeKkZEDvoutwtzy39Uf+UamKJ43Ie9ytVM7vYTBFOXZR9EDni4lhh5RoluT
ZGAtYGxs4977aMh1RoIKhofcHoNFhiK2GoB9oVi/5cqUaWY0bOzYri7TxZbor3qQx2O+HTLLZ1o6
35KHK8IQobubbH5+X7POwdhicrSkUp8IwWfdaXL36jL0x/szOmamxF70C7JeYPh6DgCDHZ23XU91
GDqJf05naIfTqme7nvbw3v0clphwQCKa43j25L6bR4gRN546o4+ih+81wfM9riEHCp96aY+CEi0n
xi9QdM43xPThDFGa8t0WiUH7hCK92Da2rHK5TKCXSxIvwsW8LrWXwt6DKvv+YXzBU58y/PlHJU0v
04dlgocZ84V/EvjLSTwc+SqNh0byBoxZHOliEpnDuTgRpeTYRh8W+nc4zbVntZ43ZoGpRHQQCVW9
Wyxd5hV5lyw9BKzCG5czLgbc4iF2r6MjYDHnQJasE6VfBSCo2uya9AlVRy0mHA/aMxi7PtAFTGGk
rhMb0i+kgm5sElEw+0LitXbpZEd5KWs50AnrAJo58OSPnd0tdMKXlMmSxRwnexRButANVLR9aACu
NS88ZskykaRU0oxaOMo/JR3ntUnAWc8nz3f1mSPuhz7gHCo8cVaqpvoIcalH3JSYjA1Ioy0B/j62
2p1Be6/XJHMC6XFqlDpGEObmkQ3rIMf3EmL83EKA2pBYBcLvqVJpXILUMgobDpi6foIbd6ZQFQaL
tvJHMoi0FeNgxcEPXBv7/KONyDUzag/Om48P0gJwuGDCqLT6anLO6VlUJwNooYa4PXFHizRn5Q2v
Hp3jOmGvJU4ry9Igu+OSAVXrzGdGkfp4Pzz2OxmXXKG91+GI02KYkcskM8VQ6jxyTjGOPgnFNIIe
gmrILa6UiYYdMAhV4ig6urODqPWPzITO26TnPPcQ9vhAobIC4bDYh454EZswWNjmkNqPjeDvUEtM
pkzQwUfetw/f44vJzj9sSolrSzvHOh5pKhS/Vps+d2FHGNQDDkr1x1S9H6VvX190bC+iIT1sWch8
t1b9OjekL7bTLcCBYkJgI+pipCui2/8UzT04/ul9ZL1JrD/wx445WpoN21iIAPt9ck+5E1avQNQI
uf9OcERggahkJJFI/czlE3pP+8JoBeuUQAD8LCUYK0EfpiCbhmW7P1MNRwt4cEXVa651DVvNdDRc
zp21qyRBba+MRW1hJG9PbmGFKeWTlNnmwp0PEfBeNCWUYMHMvNGOGfA5Kd7Pii00w9dcb2Gm/eY7
u4DmqfoZI/T0rjODK73IQyGVfyu61TGpz9x1Su1ruvYOyTOcqjWrsgeoh6hbJXwzZ2rG2L/CORi+
GP9sQUyV5J/tW5FQmAWBn2wanAs478rUcsatJuG4MyQWodaiFAb+jgwVKPKrESra189pZ31+YC+c
e1eUAeZX4y2GJUfvkjUHR67MP4PgML8vUd1c2+8zy3lTBUhJ/QMDG3sq8exzcQKiffkno9Ud2XRd
qaLyJFDiOQOX+bmCVjbqWGQvy1xeB67KpEgCM36hRGtaRVREsPS5MTonYXL24QHEHH2Ie/yBnBkM
i8Ex/2HYhgBn81kVfgN30+jHmE40oSGMxo4uOxlYHp9C2yzFX9zf3et9Rz9gc6QCOD1xnrlkGk+y
rQPqkOnw1PBti3hCH3ptT5Aq2s7mGK1f8mBh0F8JGFUgzG8jSQfL9UL0W+W6MNIV23vVgf+o0sub
uAMuwCuIk2GlxgfOYyF2L/URbhh0JEcVq78iABaWv4drBr7061ULy6vgkvm3AnHrEZh/YbQDhTze
heuzMWReyqr1RmEageshZlZEVIGJjDsjqZEd/45YdhYOJBOy588fiSzxYw/U97rgGK42FYYmJkKY
+TyIu+2ogAHs319tfnp7lGAQqCxPICV5OLvsPZ8ajhanYiUSLqOu/jWNOpBiVBcEvwBsN+WimGCe
k10JzTK9FgjqwAzT00kMfP6HKNcrnctZ0GH2IPn1SnsWlRr1lexqOH4rdy6RE+nZXz83pIwhOiMW
81+rwri4C5PF/fgpmwg3FeAHXCtKuo+wswQaNuUTLlomZ1jZL1ll/uJcMvoCV73tqrkK1RQ59jv7
vJzbC0ME/Xp9u4ql4q/7vyaam56xZikEbFoaPAiEb/QLS4iu9IZiNiBGBooUn1IUaPRDL71P1OZp
kaFoN6KjYAE9gk82yXL/wo/1Px5VLXhueEziFYlHwXIgE/2iGBMK1kbB0wZYSh97Ym3OnasFfRzX
V5s4dt+XhQmksD0QmXiFEHZsU1ImdBq9wfOwWKeqObSor+oiBRVYgkj2+1jVGYN9Reemr5Vlv0KL
wJ6XCbDqUB7guEnqK8bI32w06bpgB1E+bBVOc7nVnqjSpIXk44sRnGvtQ6TvEuKqwzhqX/7OZfuO
u+tjhPV2IQXzR5OKMN5AiK86oI6hHMnB2IeJIL4xF2YNuvi0+5yH80ZVTo3bUZc+GnqD6eUChT81
5OucTkjfvLGVAJMxuQ8wshDk7Coed1+0zp/orX1bnx9OojK/8NmaamfUv5Jvd4Caazfcs1TwvzJ8
wr4xt0yO4gHVj4FHwhQpcappq1bP2gnriMZcdg323SlaVRAR9zMwwyMZfxJl2iIy5f/+lvjwjpyK
wta2Kku7qYuDE2SzQEM3DQyqXJeoo1M507hV4TCvCxrrZzJ9ognkmCV0ISd0ca/nqiQJxrgRhqcp
pZLcGzaekDi1bgtHs8LxeJi+IsEu+cTOrfa5Fw/r3GzXjtm6plzl6DXQ7ObT0PUcCs3j/tEY9z+T
cbo1hCT7vbdtQerIRlEQE+zDnfL9dboR02vrglXNUoE9GY2kJJ7TCwpUa13yQEPtLaJzr5gCN8XE
8lzPppPb4MxiKVcYxOIRCTMsTu93+CrRkBRHdprMi5ZWOvyowsZaV7vSY0avgaxsN4J0melaOdxA
KuqDu21mt2pgHZ0WvVGKHZiX5T+xQ8zAiD7sZ7RcwMPM4YhBV4iKL7mFAwvr+rqYKBh4GBV2gZSx
TwUE3epYtI04wphtI/yRnQfIviImSgLYK5hnkTn5NJ2LUYZEhPH3S0iaDJVJXVpVzq/AjML0i2xK
lOyNiNJ17U/G+Gp8ScGuxxbYQ77Q7zhKJ6UEpyo1Igx0gweS+ULPa5uKwQ2K67llZ4VDpTGWbaUG
W4uqOAI1t3hl/v7EuBdbx455xN7x1S78Il6Rcnk+K27yabs2k8mw64rJuja/aRCAR0OnJBarX1Go
ZlFd/XYx4Lz5cYZ7FTTS0Zmmdrny2VpHKZXUwq8hHxivS+ra0h1ILzxioiVYgQH3CK3uKYurwSke
xemAJbgvcsSK3qMIYtOirHIgp8K5GElwB9NHISO9zkcu5FCoWFN5GQsgnmV6rgk5uRiybuPlBPuz
nWP/0mjZjcmBNgz3uVAC2q9hU3ANvonTQFjamH4ijOjiKYAiVPx9ty/sKI9WNFAbs0rA39JZ+ies
aiIOHycDe2uhu7VtRQkhCoB157pVkT+7E7DgmmH96vgYNqoxbGboH0cyLCMUAYXzIbYzxsnWPLfy
k8+QpvxK8DL3hBszY5145Y7GsmcfNcuc2K0ymTdKEa8YsDeG+GC1elwPB1NmW9dKrIA+c+RyHt4X
yeD9kUYDKZxk7iDFi3KbXG0/BREuCa1WsU73Gf4nAbLJiIQrRyCiCoDeIPYTx65fRJWLx6sDIEEc
HjHAZTGL6xos1PwnFQgC3OcToKr7oDN3uwwWdkS3+f+Ic35CGE0ADSrefs/7MLPOk/l9CwCD4doy
WEAlgjKHJ8Eecn9ltbJnhnw86cYo44QECAKUwGHiXXLRMZGzx670mgDKKuYhdyblwHb+cfgWcGhC
O77AtRJaUVOsqbi4ZVLPn6g3LESlGeme42z55Fy85NcwLFhMiNAK8GtwpVWTZZPFUsZ+qKKi/K93
oRSPG6MgRzrQjC8OBXEtH6L34BN4u6BKioAc4iz42KAQs0BxbkUCq59FwEAH3u0PhQ2fFnT1osp0
ZC0Jj+7JmOl/FdeVpIYk0rMBhk3pck0kG+rz0D3yPJCAmLBLkFO/CwTY/NLuXAjM5zU+Xon6ujOc
65Ir6iRPEx26yUN3JqDxmIZjGyFfV3dmjlVTeyy1VFTH1KV/leiYZAr0DlOgdbtcMo8k4ulSCC9H
cuzG91WvYCByq6N5+DP7V21fo/biPtCpPAak/dbUmg1R7XUO0uf4fw/n5ElYU8Umw3v+ThxkLcw+
DwL2sGOCvln8vBbolAi3VmGIW4ibboCekcIN85k5p8mDrsUXKJDfveniATUDAKfMOK6oNUc8nW9e
1J4V0y9qM/ZRuX0buOE958WzQI2azaZdSGmWoIROmaeIXHVpi9OBVNhx3lM4NPLIprIY8jAd6jvy
5XCm60xcKMX0vcacAS1V94TCWHyp49OeYmV3l7u955IcS8hUyYa6wb/1oB4WgoaIQrpem/AoUGp9
jUwFyQ5ICBVBVTQo0zRtqOEy+uap65Jt0xgCEWKF3WZWLIn2kFBfLI0nkDohJ2oXkMOfMUqu+d9n
+n1hQgH6Algysk5hj/ahiCc1RH2M7SY/HCFnAEmanjE8CcaQY5Qgz7r8TayWdm8wWj8Kw8rFWNWC
fw2iNjga0baNsz7IoYMNJ0at4Rn9aY2/nJWdOKugBGkJj1tyvaL1PBZP8JIdxQISdbLnrSwJvfS6
k4RTRP9kQ4C0+TCBo6DyxUTULSg8irSsuNkHPtxR51cFY0XRwszJCek2qdDFksXIUZFR1frXrOnY
ywWthFwP5lvY/xvb74VYuKOBjocYs6A6bejyCVxGmcV3P5Zc4yoWc8q8+hnV6IOxORE/f8iFsW9q
CNiq0w7ylfMEEYejX+6hGhXqdNY083U3EIKESzRHpNRm8Hwxxc1Gux8Ky3jKjVS6OcctfRjG9rce
8Q64hbl28V90JY9A7g5S2lnuuPCxI7FQbi7zsNKh5oEIwU3TfVBYZqGgNfeQ02zoBvvC1hHGDW9N
wHQ+QnaujbuFg5X7zkOKuELPWq2xqks6uYdzoeszdukhOGuNXbEqsOPDLefoBWKfz3ywYQoHOZa0
/awC1HNkFrfnU7CH908PvnnSm4bZgW7vAUcoaCLpnf/NAX5Pb1i5040gagICjXgSDOJpn96yTybD
VFCT+6hMDXC366EMgUv6oLm0sFzKXOuN/v1AzMYa86qwyP+X2TUmAhz9U/o2FjSNO8A5gC7aJeUD
+al5MKCkilk6KD14RaA0nmZz0ekhoSBrVLeiM1AXCv8Ya7dZStkdNIic9oNPmdtE963T1piXOesg
8rbJzWONI+JATv7fAkvAqrVVEtm8fRwrHFGJ6bt8OQ7GtE4KlBxCXQ5/KyPvnh7dNmuPmZRkMkbC
LT/nnr2dw20U0jdBg7rSN+dNhWqSzoAEVE6mnB76Vn2pv6idpx8eo3BxGMftv2CosRqDfOGJ8GOJ
W2SVG3uXvQWMzAeDb2czgpcjBpTWnpl2lB/TRqkFUjfJd5ha0zVUD23zoxsqiOJlB0SqhEj+lF7l
Q20gSQh1EmiZB+c4rZVgOHnxGY6Pvm3nxISFqyF8lQ2D1mf4DCEJZULiE0y4JtgQPooD7SfCwoxd
RGNCcSoMprOFU11OsHwQaW02uSnWry4fgSuR0Tu5kZYu5KZHkHaUsS36kBvdPImrlJ8z5HMZom8F
EsR9lzxQ/P4F3Oyi1VIAiCAaoXdPDxvL/e169jEPVqXlvAkIege+UJOZtusketjQ0mmYyJLVGe94
Q1my6wpKFnA5RBZVNsXtmkmFtB6gj0MZLhix9BtBIsqD6AqCW6So4Sg9cxv0sXeSdCOz0liDzKgf
uXY+Y4wIqH3hydDTy1Wtq4K3oQViU0mIeV1+rAmdK3BKCQAbe5+UEutBS2XZxbuj7AfGBvojBapP
kgvnIjK3ZmLrbSRmvQouckLwd8Ov26izk901/OiVmkLkBk2aakLfX5qWFiGLYUdwFz4JCXEaJLBR
O2WUeKR0asvN/WcYhMhJO0+BdnqTF5nwDoTNlr/lTGUDeF3Y1FSyBo8H1LyC5v9apjZ0Da1x6o75
6xYOTpSdy4GC9dnVmwjcJonMuQb46Kmn1uYiWluQHOBE3U/0DO6bjikqhPm/cuwm4CLvjoodw0K9
Du6MOC8BwLio6AeXifq/v0Wd69gzijXpwKyRWQxZDgwWHoEVJqc9oYdciobnEJMiUIwkRBBBi2mr
u7OGLLbhR0oX6oCIrZY0TOehguYmEKJkTAWdRdlWpavDXhGXVpXSJP1uwF0HQERXEJExKMQY0sWr
ooDpvd4lD31ySuJwi8aPk1DhaiR6XS1BQShf2XQREEuC8c1DEp2RtGZfbZb9ZV++hLErg+LhDKtx
RQ57Q3TIZ0yfW/bXOcsInP4JiJXqg9JLNcMfAOoX0HVfsu6zImQ/MyePY61IgHtrF3LeOv4J4+v2
N0pOLwyzmY3rOFJuSG5gF4hB7OggwMt1dM4J7saSUf4/8HU7JktqOAMf1pGj7Ftb4dMq4guxe5E3
t+PnMzItWKr+MNcF5fAkD57tND2dBRPSktTZamAYiEp/p2Yz/XCzirK83ckjo22bMrKVVOqLYSIt
G1Qm9PK5rmo5UJk5pnUy9aeWUjySgzyDebN0W4DplI90kGAAK8cKtIVmWz+G7GlYc6AC69Z9erOf
gffjshiUE0Fp4b8WHB+5o6QQdye1B+jgn1yefgxWf88YGUfwwPB2XY58nTJloOKqjssLWyrLNaEv
G7F/vazMfABd/lXDFpWDN2BE6hkYh9S/bFLVNCJhVw4RFSMUc+zuNaOrRFXesQ+DrCiPpfS1kaEW
+pfzly4GsSPEcCzbLhWxiyDcuJ28cCc5QQE3DIGHHDvY6ldaIlCey0udSgl66Iw+sp8rVYLobFmQ
4B3iD9xpi8XIAUnhdU0/0h5YOxqH/GgMNGF5zP7WvtIsFoEVyHu2SjKER7FpwfRB9hZEHA96JrLe
Xgq+AhL3nhU3p4+tES6C7e1z9Fuvsv9RWLEfiaIXTHy9z1gWy/+ZBTAQXuN0fS/yN5OdPs0lj5/t
mmScSDkIlS4kyNNwV6XNkPRfrgnYbhJqGqw9nXyHRvGAYw37kpKuC8B9K9+3NQpi44BwJLyfHklv
+ZxX8+rkrxXR07eVpXnd7nx16Q4mqZfr/1k6ClrknE66DQ3YiqaXeNe41vdM7JaBVi74XexK5I7c
PsYsLTpKufE6NqVWBDu5RbcB/FDaSKDS0Qkf5cq0U/lHcLtVnXkk4VdsHt8Wi+/CbQC67RsJPmoN
XW8j6i7O2We0Rp0S4LOja46r2UI+1QlvCeBJs1fRtBKO2fcZnDBxEOjJzQjTrAFBCcZuXb/Vtqb1
gjPAVvCb5ev+M2XZYnVjTbumUi4KVyUjOHivhZaZCLWPGWc27fVMFoVYM0BHULDPlCT9SvHzsAHX
BOe+dDVqut785bfDzIy0L4hHIBTUbzPwSEdJcexnJFTiz8L3GHs8Yhw+ZcJJYobGdNbt2lzyGdyd
gQphgkK7POp+vax4IXxKipfeovL0bYKaAcOzp5sP01ySB2efG1ZoxBop4f6OFB8RKldpqkyJigdv
BSh+5IFxRqu5sJmr36h//UUQiPUfSWBTnfBC9bWU6u1h4ZIn4eQdRAR0+EvaG7jyNS2r2mzqRkh3
Gh4s5RN3SOtjL13h3LaVLG1y3wq4TnWqjlaiOfpQgV9H8ngK45PTVAAlCgsvCZtFjadsVcoO7rrr
nrEnVkh0LHC6n11MWaPqARrEyNO0+ULxFDIYX6sbW8laJFgmLnhaJKc8zKamKp5duCW8TCujFvVB
sR78ROzGBPjm4FJ4HC8NB2vTjLJp9N8C7Y6Ih24KsJUSGnEyqZ5WwzG/dEC/sjAbMRXimJFV0B5h
UIQom0qiPSZ8PobDB2faJC6cb8LXabPHf5SdWR19HMuz28CJnWfjV70KH5e2Dw5bGWN1QJ+wCEFP
Vbx/B1HnT5cLjuWPVc7P8huvAjTYkPdYZ19jyYfKslep47I9Ce7g4rcnttHp6R3fLu5vRH9ibCDl
Me44HtZNohcoOoFUlHUkRq/QrrgStLWqJLq8Rh7WY+n0J7tdKpFiuT6NFjV0IPjdPp9toefRVHPe
PH1CgF+1BBHuNNQiwor8IYTNhDIGSSYeOuj7k6BCc8lzVa3buWHlj1xuzrhf2JWxxa4JC+lKD8QY
TaJV15JRiBpKwTIoehl2/GP6N8w1TrMjluH/xdG4IEUOPJ2HiiUgRAS8zbSBH4E1Nzz3encjESnu
+Iqyd9twAP1oo6gO/7pwsFi9UjpsgHU+lYqWot67Lkc+LF35ynZxGGqOcp6lMyfL00t+Mamm6M9g
tOAWRJv9LidAIW1+QybiecewbKB/ShGeNBVWvvpToci3xcXrvWVncvEg+Rz8AoCPFUMOCg4KN1g/
BO/HKLZP4q28lvDcxZ7zQOcn1JYxh5B7ikWJSEj0rQafwFNrlFkx9Qq9uhWkIncQkbLxXY/T6v2H
zXGCozGDeiVB9InN64AmnOT0as4xT647qmX6jXRBjkAX+A4kXd+iOFAFqZWGReumHOr4+KWKy80m
x0BQDZPuAvNvYL6LZfGHltAxTk0MMfQlvjfRzl02wQRUpiRbeqJcvaN0NCEGU5s1Ztfn4X2jXrOT
UEi6s+3nQQe1WNcf2Cshg7mhUuY9nREWWaHFoBYfLdUVzTPaFETA4rneY2kGP+PWWnMJnG6rOGdm
PAzONsP1to1Ub9G6PXCSGbJlciXEOm6F5HltgC3F6yO5n03ixNsk9N2b18TCqdDmHGHX69wP/j67
aDgT4fK0ofurAVYm/S7bc2AWdFWkRDqd8KfmnpnlYvq+OkPl7HhU1m9xZrJ0EEq82BY++6LODXGc
WX8Rh8+ZV5X+KQzS7sR0zgDu+SOANzJgTu1JXRVtOmxNuUtsW44l6GMno8Sh4WoUj6YFfvQBgIsw
qjwOTYWZ9v8k8BNMzQDMzdBfB5L1/4KOafeIvdjPVEpT8J4nFpUIIPKWuDq6eNB39MkRIAN8a9I+
SDtbWneErfRF5wZR9WJ8uidl6CnmAULM48VYs+M0FIxv/28DibMorQpWCYbxRu0axmKxBOuv/OI7
TU7BV/sPV4jDz5kSwIDi2rvq6ccr02DMHjaeDokngXz800lfmR/ociAZuxtb9hKjHevTFAZnda1X
UBHKMKk00MJfIa2akNS7Dv7aDLAhpKzmFTFCM/LgQcu1m4lIVIJoJaXzDuAAPvq35mMXyffOIOqj
voVZiu4bBHNwQ16rbD0ELQ2EWYcNx35Q+vV1glOz+9XsopC10kuhqZVpktaDdmkVKE0ulHh/7qDe
sGppwZSMGW5ClX/lSa5KRNc9rZUjgXg9S7rqthnuWwme0K0Udty0a62NluC+hKhw/KTrZGfpN77t
u7ytW9vzX+0qAUFMs/xVXI8J3ximECeWozotAD40L1iuSt65IUYm06JsSzfSKXyQRQ7uyi8ZqpgI
ujuTdc+KwDeWM/rvqnYI7l/Ht/b+nQWP05Iyc8i1INl3TipaoTjAbrwHUFV71Jzoa7Ghzue0+J94
mbLYfO8zzpjJR2PDap3sXd/Dm69+cCTUMtuKUIDTrSwyAFO/cosmC+r/w5gR91BCJKjxms6jCRh1
Nbi2RTvC2dJ3W/i9SgPVdorQ5Yn29Gyo6MFmpVXpUTUfflnR3MuzSGQe7wPLu+50BZk6jDCUUjd0
6pm8nSD4zw2IjGpUsJ4cghlqtZD6xTeSK/xL3deGgLi9/zttf5cEOVZUP5tjmBFVrC6S4P2bqlxG
QsJseFNa4J7c7RIWiJRUoGzqYt29igkQk9tlIF09+LR2zBrovEz4c1JQRiP56c9GPqxnS39oJ41z
m7uC9tqsFaMBNy8YbO9Yqr0kz1tsz6TkivfWXmy/uobGfCO4p5sPjmZ1Taxhzz08kh5zima1bt/l
U7+VgX+Qz4bhIk59O0zzzNuZXzq+c+IKaVug/In5YMHaSSm7wzuRIl/QhKZ7ueWUn10qtC8hZ8V/
+dssStH4fZdz/GsfhXqhY+RUbVWHwl2tHoOpP6z63S8koT/koI+ZatxKNRwPhicAMpsmYqBrBpR5
kpXnkg1vtJBtnH3+XDy9rURpjC66q5BAlhmza6fIhvh0rbGWEpgNgMxeYQvZE+pT7EDsJrzLuD4u
xPMUgxCebcXaDehiEj2Fx8zGyc3zXvHmN5+3GLTe0sJcImts3daxwXhmNIv2wSbQUhrbKfPJdFyd
QXCgmf1fBZNxHdhWdT5pVmWtgF3VH94IUzT75/kEYYTgEAnfm4XvcCpwgK5RL45j6tqa8wHUCGC1
+qO1wPSB8Jgv+qqw2dSLR6mTKP9p4TTtPtlkUvxj7BnJcn9fO9H5d1EQPGsBswvqth2XN0qzHYLi
O6dxpH5KZ09ZBCmXQ9iP0bHOwLdqlA1FGDRqmAtts/5QMuXSDkUIX6K1bQoUhOI2J11cOlxUthmg
sJvCfMQjtEMJuIGm55aWa4u5VyRcs6pF3kUi9y8mUD6Ck9uRBcyTEJ/26CKvR9hIOGAF6RKpAN+E
HLMFftXLhobgMIYgjQXZRwS5JrIxn5RZFf5b+S8Q+orebJ0PSfguSeXKgaVDHq7HMJb5elXl9dhy
3KWFneDmLiETuLYyhCo0S4IsES/uudzfRJELDM/seZM0z4asUqpQb9CPFqvIT/9kOjexy8bB1KYC
whH+pnBa7lgDHGrNCPNW5vomgrR0ajQQ50EraSuSWUoFI4E0hS1Y+KqLH+ePR6fLaum5fnyEaUyA
XKtp25Pmqo66sNP6X6XWAmySe3bJEd2U09ahPVWYW4htrGX6E3ZoqpYdrAgrHpgah+lysD12XT/Z
0wtwlcjei49Nw8DAGjWDE7/SHxjZNyqpQZKeTRmI+SrO3LelYCOHMgpiX07lzL0dmmqtI3+vBUMg
vJFTz84P/uEzNvk1NNKqzxX/2Xm1djFSMbvQqwFhHb/mvp3+xcbKwSAbju4ztmpUXQ3cOTZM41R3
KJRxBjULzHQc5b2BLUmAdfixd0GCC+jEr4Efal7DPUMrHjejpENdEHJAgr1/wSgtZyOF8y661XlA
3QzX9iR7x40arHXRK+9I3B9RRSc8GnFmYXNrYlBWTjdafGH1PSeeLzCssfTSz3oJ33x3hvuJCpZD
NcUn8YxWI4VvHCEI6Zbxc4eRT11nplLW1WOQa1RoyA2fJalhKC6XG+YajRFJzXUZSJ1ssSTPKh21
jhKsdoM3f2N2y8XRmCorUkniS9xeJw5dm5cm9Q9p0sVLxzJm1jT1jceYsnX7/B7YW5bhxrYahF3J
m+idC2jH+5/9nSWPtbnLkAw88m/Jml7HaWMMzFHHU5WdotIzbl7id8Wv+wduL9h7Zd/oR7CIpDfb
BIF1okrkOE9kME7LigN7u/GSG6nkX7riPofCoz3oHB1c993cdtevooPT1X7frTFSQY1QvVpyE9tw
46kyYlMJHr6m0rMrwEgHmhikB1LrhzfyGyzR5KraHKL4/gpiR9MMry2Brnly6oYf9tKLDd9DOd2n
wBW7/AsIQJdNSSbHvAuZCL2E3s/gWJMvmlCVRpzRHVOWaowLUAVw1u20xqg3rIaPfgkYHHOkKsld
CVI2/XYj4pZ/oQzrziwU3SECeYt7uFTrsbsL+BP1ozPwKDPySf7LggDDWvZRN3G10EWjA7LuF3pN
vtQoIo9zGhz95oTCs6ofkyn4oMzR5YMUBiLqwZ7RpotKMAKmSxs3Q4keDZLwCoeUuuY7CNf2YFNY
3IRBkRemBnv2bojSAC7esNDCjwmNTC5PCblTFTT4+E3dFplQeTlIF9UQgCalWD9rJBDiiZtusqtd
hBVIbBq9tUM2JKIM+4jcV5dEpksQgJoVS9uhCtgXKmDjzl994x+gelqX/wumWyLpHy/CcHaSD96j
LfpMlrzKnA5KkiNM6yU3+6LakHK8xocyI329yp26SLaD1Hle7J659vxrms9uCK9Tq8TJJWjm1rVe
iOhBocCTVfMkjZQdjaRGVW0p6vvg7jc9ALSWeYSHnzAfXzpkii4EIAOsrJXNJfvxD3NZL6RqPnZn
DQN/Z4z/br3X0kpBlYRfmvo2HELuCyoh1W1rJPEgCzsKaXDQk1K3VDxjTSk2do5x+4tmiU77nVhQ
hbxFg9CoPZ/wgRadZPlcPIyiLY2svfwb21R45J+OB2/pKmS4lmT5zfhY+7BTZxONE4Hc6xVPrVWN
PaXk6/mLPaXK4r3RWu2pPXW8OO6hxMfnWukMwUDBSD06vaVKi3GUN/x4KCw1yXNA0DeX2qKKDfyy
5P/FZBWIdEsafyBKsd+dPtspIxJJ3h7TRnWLIUugIAZAsIUnukukzzopttwGmQrSgicD2cFlaDNw
R4YqWMV1nG/ufRkG1pcBMT/cNEwDpjp0SnLR3ah8p07g1ElLurwhWBmHpE0HlXigCnLXLIqBfTR6
DeC4l4+MpqqVXOwm/a7Exqv/wStfVXS8EyOgM7auPai03lWo8tnAOOLTtTH0aDC9iANWvSkZYOtM
LZDwwbak+OsdTwRLU3mdlCxqtRuHgibvguiiRteUnH9sie5fxcY3S8Rpu8r1aLGrNiQWi8DrludQ
ZLBmfRmvPLvwUZ82+xIfKrzcZQc5KBe184+PiB1vabWrls3nwwn20xV3dwa6Xs1mLOXeqh1V6Edv
5+4nMY+SiqXt+ni+Sn+ehvsG5N4DYD0X3D9BIJDF7U7Sk6c93SOnihw1VzfBoEm+0qAK9J+XXm0a
ADOxRv9JXxX9u8eHrvmIjA9I6rV3rI/f1pxrDhsFIlPQRMejKNxlXSpUJY595bLBd7npkd0bSvNF
9Diq6LoaR8sjLtZ0sVviPh2dW3K/DPmHA9KvfG+8RDm+rzYiLlukaftABKajl3ZDkcouCbm4iJba
AydI4zBtbI0KSSwtskEYZVKRQEJdQPZ22b32JQUw6z9sUONlnUrZ22g5rCz/4GFTMUxxBI+3tgSI
UMWLyR72L5v4fgmWxOt9dSeOsb70EMzWp6YavwrOXPbpSYa3XmPAyEE1HeN2stheaBHXSXI/6rvK
dykxusz0Fu9pUoSrEb7ak75Y6nagXHJX2ZKmeEtPEZUzx6LcnWWpsRPl1IN5n4+nh9Q86k63GLiv
q3TID1j4gy/gxbUxTpEEaBRBXwj6JLhMbtxGdgqpwDvC+YK3IYwr75zCegBZiv4+nVGURRGNrGQE
x5EEUvC4KZ7QO8a3YiSB0yQtRYcsa0aCZfBd1bAhyB+HRjf1CjtqvkRmK6VBm7W9NJ1mqhLhrDyr
xSV6YTLMvc3na31FS0zazQBHSQjy8+a4VSiemIbADrGNqpGmGuF7yneGRfcG1NtV0RdxsTVVzKjj
Zr7VrP9ivu88CHv4Gwsl7cMxYgxks0o2IQ3TG77Zrw+Z3I1eiPfa6GDzJotEURFOLIGGbwIJD4ix
Ye2W6nqHI4CloiuEKK2923ZdSBFo2CTZVkvSakIDs5SdUAFbZ1oJ5IrjzlTzGUu9q6Xz6UlpPu+9
JkCjwd5iUkeZA1M9GRLeqkd6Go8yYxU/xdPkyOwHkdd0+d+M2lfygMoa4has+F6I1olvu3JLTyPA
HhyFUpFm4pAulIGjHlJSMZqQTSE8a5C2wAS069/IXnuc+8AfdwAcIXVK50wunpMvpS3XpoZoE0Xk
7nASHJ3CKmbXHC8AgVdmSzQBitniS594es6/yhT9bP8rKW7JWWuunt0imnZJMpX2/MQOIg7PuR6H
cMyWhE3si5WTPO4UbXUlpAEsxIVBjmM3Ku+2wq3QAZeo5p8KMSXXyNrAyw4OfiNvKdpm/rWMZQKw
ebwwlAr/ZWM5LYPYtLL5pR8PQCeTDIITeZZvPvRcIjKEGlUKA95xS7Y4eA/ojta5sva5AW2xMBz8
4jwO2XZ8+C7YhM+WPrQQffdbeB5zPDfC+fgawMpeH/fwkeZssesyYAtXfxPXDOuM4jRKq4YVPcFx
HcZhh1u5ZrTHWHi/lEBzC49xSPeydQ6BhBdeO4/cYbVQz/bgShMwrn6qUSxxnbywkaPG3CIrlgjy
wXmtXSUn7ORD3XLqhIzbBZBvVwH3xKxVieivXmLg0mWtchX0olTDAZpowuJ6hh/VSp462OxrP0kX
/+H3wFPNDTkmHUmMxAJ1FTaJkMnqifEDqOKKa+fmEiwhRYtVwOYSO6oAe5/NSJ/FZK1vEmwJeNRt
Z9GtrLuo9noPm6eSkF0dN9cEwKShFPiNNbbjiGoNg+0bJS3EWRhCbGkXZWfrg+FRRRFxCMCFO09X
TjmZOS8Hk0wfPNXPRRi+XXuD2UlAi2GJBIkln7fM4nB7Fr1/ribMTgo5ryqI3MhV2qZWf17fYHlC
R0ovbio63bPQmg26BpSg5OvCTXEOQLaODjtIll8E1vRBkmUSjk/ZitRCqX+cf9dyfv6gszWOGa+s
0gW3zI1CiSl9u0EyGu6gLrz/hs3Kp0NPbdngctMF1j/coUXGSW11xxcrxyUAHL2SpFgnQoUDeaUR
Awduws1DMye5yfDNYdmFHop0NPv2oWlXvkKcytsJv0WEoSXVwkJxDQ3WcrXcBEX3Br7VeUuWmqF+
0t/UhfFJXSyPZDyglo8veXVxgksTUT7P8hCzQ+K31r3RljaNhWJQqtuwnqgKDsYyv/ebPlxOEAji
Om1Ye+7BB7KTDL0OqMAdksKeOWGSV7vMWGQnw8v9R5KN3FsXFSlAeUUccBy0+dsTEDYDvgQoX1Rg
1UlHwTzOX8WejQlj//chhLCgjQeAeOvNbGNrILOWZGiTJwQO/K5uhsjqH2CrjdMPZZRzlBcqYiky
Dzynj5aVEHyJoxbYU0UZrz0o1tEzhiqXGZhrSp3i28FO5qxrlm/rRhyVaVKBcDFHgcAHnfBURto6
Rs+9aVLf2HSijJqsA9EMH6OI8wCXy5PZ5Z4oXtoKzDDv4m47C9H6RJAp6wkbbcHp9lG7aVtmSUfe
f0rWSsAAXDeXYDjeX3oTRg8wc8clQ+y9zxyuAyx08GreU26a494H0EN72QvohC67KNB11ulX1Mqb
J6SZE4dFsgXvmZCDorkQiuULGDiCZ9YG4F/ZcxwmOPiPfiOO9flcSP0sqPgDu3CTDawFrp1HlTQv
E1L0EVYLDMvpAT4KmgF0zPMWg4e4M7tVYKok5uJYMaXZpziaLrnJmkrmKoOK52zGsKa8yvjyXUUA
0griaNZzOlnMiQKALWogJzEUfA31RROZPFteoi5hMq60Omgxx4KwZB2aERo+y8orEdHnwQDO8Jbi
EppOA//YLWlKBk3CzoWPqnon8tVvuC0Xy7Y2xNzW5GAvvkE6ztRcUfR4jGQxXeEvs0GR0kwaPbpB
azcF/lmHsVpANjqnogtThT26otI8Hghcm74EVRUQ4/f5qFNsI7zJVxaQR+DdydgT+XoV/54Aeaw6
MKGiMxsYeGAULk5l8InRNyn7WmY2MAocn2I7E7c2dfyYTxqqznkn3IbgUyU+vln81SSsfbL44jIr
R3loowpB1JmpD6X6WsfxQk5cC6MFdlIF1KsAg6o51V1b1M6c//DJToNG1mq5X4gTU3xDdA7wS+6E
r/4f0hfgQJwI8CRGH6XERV0tftdDUSjWUgowS5aYiglG8kU2DoTLdSkzV4+eGNAXVwPjEIv5YmWF
LKUp4adePmO1315tFPOC97zZIOkzB61F7mE3blzm7a+4gHmsn1tkZIL6Eh/aQWKkXkLWo1M51TFb
HBeDhMmMhf6/D2omQPTRmJ/L8+9E3PglOlB2tFKH9ExuKpD/x9ajF+pE0LAoHkXxPbCYgdPBbjx2
RKk9J0ocYfz11Is6hgVmTOiCkQQiCgvI/6D+ukebPTxBjuHTO0sNl/dQWYlRTqCgVhLICVg870w1
M3UskQs/046LrnkICiE2KZRjQfkAaZNkGD65mBss9//WJLWQ5khT1yWfwjF+nw+CWlHNxcxLnKBC
9nYDZbgevWCST2ApEeo7IQcGjC+BFXSgvZq3hIssSiNgo/IEKiEUP0liJJWNqQ7rHu0m3esW6V0D
ZQr0klaF4FaoSZrynlaxxSAmnLUoPgC0VWH3vCZboDrCdLBO6UgBDepS4JYdIljhXUTfX+K0i6FZ
3cosnP0GnBadZCAOnRi2CBtSOHjwoTpHY9T7210C8CcA69Lg3Bqlewk6LbD3e5nTliG4fEOV4VdR
43ok6J450jPLNlfwcIoBLx8jaxwlDPHeTujx0Rk+dp2zO60tRVDKS7YRsLOJcHhJsSUpxTRzzBRk
Ru+iPxk5fGU3uuIVDEu6tcW63XKSRt3B7hkPuSKuNF8RDO55XZpQ2Fu9vrXfgw43P46520Ta5FVd
9HP8/CAVF3oawcu1WVetGTw2y35Sm/YxUalOOCnq4xFFFquO0ExbvyXmZGL9M7dupSHki6kL+dBu
ORDoZdyfN0gF+LVWnHeOh+ydZmypr6Wry/bAdWZPslxBpPshJpx10VR5nQN5+IZYZWkfRhvXX/xy
jlLv7wiCPhD+kKHLjJVQxOyX5wQKHIsQ2/38FHgz1UXGHziqtq+9Y5IkgBuQREc5xoyivkXsSVs+
/NLkbG0GvLhaOpOrPBHxIzp7Ego8pz6/swDq3m5CmyJbTsL7PiUgPVhMGkLD5ra966Iy/Cn3eEDi
qMpA0nvoksxNMs3NSWOT4wJRiGqcgxK23da9FNMwX5jO2UhRxszWUzpynfs2FZe1uxaTIOp4veEq
+SzXHTlxbnl+Ovrvus8YtAxm2lnwloz6UIrXBcEL4f8Xv/xsm4pOGxnKEKdxlK+PnUDOVN/hzTLN
SB8DIY4KHEx/omFHjpkZkjpBwiXggu0yBGj+4czf64+jviqwb9HY/5dCvYyR0vZRCJCu+dM5Ohmo
dMeflI1/JbYPMFGVBjR2oLnetJikJx+Z9kQBAIPehUjTZTp2TT9QmBCCWC2U5kd4ueZqhMmNH3yG
3LKzJS+3dnI2eqOLIfn5vE7r3hkBwB/Q3DRMYi+T6rt+TK1y9xjCTQhPVIjLSd6WsCEBlD0Hut13
5KhVpMALStKYD0maEzW8iMNX1/TLFM/vqDD8oAU43A2xwiP0Xbs0m3hRa710XhYaMWRMKvilasKP
EpkkMHxM4duIJV2zMGkjmqN/f3YoicCUbknBAifO4S6r5wYTQ+MXdzSp4xR1WMo5QAEwE4IygX5+
gmU3t4tWLdIGNmcHGoUT73BMRIunbKL2MpGDggRQcSkhSHibSednTfe+koSKSi3Un0aAlDSdezNP
4DQBzmpLBMeHNT8z7+KSWG0vVwYrv7T75K2BAwajS6vOq6FLr4HiJ4lEHooXW9N7Mxby000sruLi
RAw7VwBflk9zONIdIuh6bbnpEeixHl+Hu7ChA8dVql2fbPcvm2RIGPKTTXwgIf+WYdxjvd6eCyOH
HdW2bZTvCDaG57x8BkWoFKLIgmNmOab3Nkpor6vx2jLrJ1wNqr7PF+yR9eVYziHXnc0b3J7rt3Hs
pdRKi944ya4Jxj/EYR96c/bV/C0TBQ5Y9SvzUCppiMsLfew6RqLj/HTSuncdcE97anp5ZSGAcoU8
cHlJkAE3rLwld7/zI5ODtfO3VmM2gfbXyYwdMqRGcFt57O8/bZvx9wGfyWHE5n8Vl8KdFH1RGxHR
dDzNZqzShXTIFDdUEp3k6XPJZBCbht3KeNcfAJoq4cokms3ZUxqbYVE4GfOI8YSn8TYz+JptYvGZ
fYiO3owtzuGmycfJbk+01w+DksoqYTCQKZXMFqmkG1V5/H2HBYAxu9HssKXAPhXPvXFA/lcqrt6i
WdLJqkAsP4PRBExlZ4zSoWrMGlUEz/6WtzLEjgmGvI8RGkLoEe5VA886X3IxXvMHmE9Uj6sMcTgy
lggfObignwlfr2c4ofQxAIvwyfEI8dTrVdDFPIsVs6iTRwjp/nrerQsHnwg9dn8JGcAekPLtZgrA
LBbB80fEg0oduhcA/hPoLbZfzA2rwiZJCnPPNoy3kIkv6uTj4litBWL7Ek2Ut0zy8Q6nKD4WZpcw
2V2QTfHZljvsSMgeuYlnfP6yr7sQOYxDuoD2MKlSyvM4lyGxOaTOk82Gk74sXRLxsiJ0RF4lkM3z
++YWZw2ALLhwHTwK9esJ9LIZhRYBHG3kHz4UkmMKcPv+QCrd7nkcUu7EbX55i6ZdrtxLalBrpLO+
wXd3RHvLd1vHxprooGa21yOyAv7pdRVxVKy4vHeUiC80/8vpnbJ7xxB650hmaUJsLI2E6L3YLc5Y
3fa8b7OVzBoUXgFxTNyxWO7+Ly75ykVpV5zKkVSEE8xKSyruRcgxWJnT3bvbGFjX7aulLa+0GqCl
wjksiU/Fp9tANkLH1rHjPBDl6zO5Va08gigPkxUNLGqfqJN0+JalhOlb3VmJRmdGOiOkHtQ0rxoP
Z0RMf5M60ITrC6oMWSS/8DOOfPZI3hXR3//vZBH/pkhFdwDp5iUK82jtWqksOj6iZox76oOj9TsS
st4RR+qx4ehkvqNzyEGOj6n6sffyTEWderPbuXw1X/68xjRrAbwP6oDbX7FcB+o7FLL9i7pKNmJZ
2zXX0Zi/oD6E4EKhqa/DXyiOvcTIO8X0ZUQnFilzIEsf/XJrwgSPJLu9q2pzoJZ2yOIwwKnmzjDk
GgcPPlXwLZ8CB/kmn8l3MVybcRVL493DzXJ1SlOlO+fZarNFmbcBkhdcL41kqy4Lkpm+ESIgXnrl
TnnDgqclx1o4SJ3pzunc+929iDG/x1byRhEq5D6jHBIS6QNk/x/jbpJKMZcskGlL2lsjUTa4GjTP
D+Mt8Q8T5OkoXqG5L6uHw4ZaoN3XLOdxpmE23apCLPnXgfHDRITz0IwHW9fA+Eu6aFY6YcWDV4IH
DKDrazckwZlxStgRfO8jSECdMVC6ZgrxmFZXltc0hAFKlY7Ke3ruaa7+RZPnl+QpaM4roNKXI4t4
EAY7H7tVAOzp3A5sUb+6uTtoz0PI9cNTLWh7R/DoSBQaAtZbfX1gOr/UaQa9MxRHTmLxfAs1r2wO
PKXagQ+VGBxERJju4zkdGYArMtpkEMjCyxucgr4RUXq/Ki82VKLcAuz0a8Et0JMxzXwkb7SljV/h
iKeN1zhGJeSdAyGqkyA7sc3Kw537GRlJ2eGELAMaTSAV6HqM93WLsXxBYEl+dEMA0MtfXSHsRsnS
svoutwDx+FDQX37YqCyj83XXUXKXuc3yiY7FswFGUjzaAjhc+iY3Ug7k47247Y2+lLDSD9q1otWS
vm0oiZiYPlM05JPIcwsm86kPgPwXumsxW0TZB72alFZ9JmLkq5TUTJ2DdD/F2ynfcHfIEMEl+VeA
5rf611Zn0iJPXGcR1Vsv0ZGMDWFhn6eSIAzImS7vOSBud72UBBfsYs567LdC0HReqD46fuWRRjzE
QmWIkxU67HeiewG73gi3dkPDcD+RrnsJhWlUCMvAs+JfTS5j3hQS3Znmx0ktaIf0sRj78YS/M3Cc
BufIlwUhqlTxR8BRmzCOBq74hlVRFAy3rjvQ4dBmLIUvNVjtge6DWKHzXvTHCvEx2cfzPVzQ+JI6
2b5rZLGX4yTGdVWZ9eHdq9dCNdxa2DycwTjk7H57tAWwnsS9/MAahOkWyUupGnkCxPwKU/+glqzO
6jhNvuiRU0NC2KyxrTmQCJorkYNoyCyeY5bF1ch64iZg6bN4T0fvCnV9iqLOlyBxjiJkMy50+Gix
jUMZXNEqP/mlF5SGTqWuOX0FE5CQXg3Vo4oLLoxkWTWFHvhvtA2whyp3Ws8WPnRNs/StW7NJKXm3
ZBqWxv85FqLF0PUdmn+qofAS8Kvq+E0rhe2qBtPXOrV6EiWiZNfo6qRbUJm/eEKfIw1qnxRGmEAm
kKzAc0QPd1CHLM8uD6lhT5KFt1in0/KPdkKmTbPUGoIWs7E9PkcrASaEtZ63AJ8r8HE4FZuY13ij
jVD29Nl7h3VWUwvdoIrYAMZ0/Fkp3902jad8QASaBpBUqG4TIg03tCUnwWpvnxbf4l42tXkMHYVv
dZStn8hPyOR/3dCX0gFxN0ey/5eKy3Ar0Ji5bfIHVGh5bCC4OYPR59msgR/F8fuu8imrFGFbplhM
25lNjvs68I2SUOG4kSOfbCDtv9BISGVxhMK4Ch3oA5p+tXfJlCcdCTGldredNmMmIHnKXSnXrTsr
q2MqQINMUGjW7s5XlgPuhA0BAEQJskQ7k3ZsRsdBwN4AFNe0Ge7iIleziR8XrpBqiwAqhcxy8Z2v
mf3w11QB9TbsYxy4GJAD1hV3SJpko9j8YRn1Rf/HEYQXz7zp583OdkyRpWA5pnXxltUD5uRDR9Lq
l0Nf5LdR5j08orgiW8Gi4MQjzSccdfPmBpDnQAvRuIG8LI1wWPQ/GsolTwYHKAlSwnxcA0Qe+BEt
NFIf+WtTeHVm6pSG7iT8+uegn59MxdvVKSaVeSd2Wv3KL1RvcYCtUTskhTgSGuIj/2maoOnel+U7
1NCbG32nhcQBrM71PfyPaGxm1O9LR9aXO80K71AiytszHFjzZ6aczK3GiZI5TWfTq37SMDHjUZja
gTJCsbuzMncQLt772Bn5TjIXO+u1pCete1GtHHoWMW2j3+F3xjaFdX9xJ1qoBV8gZlpM5OTlplwP
QvUWHQV0nceZxs62A0mn3W3yA2/PROGi2jKS/ofsgY5Tswq1mmY/BSciZ4j8UZJK8CvBWV/02e0g
BWCNszX4wn8m3eq8HyBJFirpfGPU+tuupvr7xJIWwdeDe3QWXT7WhxG+smwfBbawOGzKVq5TcujF
dXwqTylrDc4qrRXTiPWlBRXlGNgI0ILSTebf8JsuR6VhdMo1W9UrZrbHQEwL+FlAJIp8MOhoTUMF
laWe2vIcx7MEr7FH+lsNFZzhRXj5PfcsHoLSdAV4oSa9NuGfSL0vyGBykRX8Jo8NQ+XKF4WmOhzT
tqA+FvjHIggYW45r6GTGO2kxs5TwistWjnAp0U0Be1J/l3b/cx88hYYw5UTl1pxECnFSrR2xFoE6
7gVb99OJEN5+8vt0CedJHJHAbIoKQc7X5kl4PksrkQdhbQNhN6unfYLMUmfXGZmTeTdpUd2KP6Cs
aZP63/KBbCYrcDGfV7qp2JNteVJ2CijW8xGlzJYSMs+H7X0M9lKMldnTabCBA6TzAZacezDjPV5J
UpYgIQNF6gq/Syz68LGIOhJrAVzdr3pIh6jHHgDfQuZVsJHotIKhvzrAGNsHqGSgSFnGiZBZ1Prw
T84KmiS8p/Ptq7wZn3U9OBT4dBYEPqJYlbkT3Kr6PwFeJ0vaHm956LO9cwqndTN1bNet7+N621VT
yS6fF5vUAo+GkbBNUyHNiCoE6UDB4J2GsgsNiOGgxWDR9h+9JtBHvDROYqSJ4tfhoS1lgZmpwQlB
VK0UPutwxM48MKR2mieK977WjxFXpqY48dMO/QyMti/B3KwWark4mV0dbDmq8j21sIRcfwhrInJI
8dkuO/blKvFBfPVlB5py5YpVWrzhonMx/ERPMfJK/WZXpRwfwOmCuSFqVOG9QyxWyR8Ufm/7pvnj
7Y7Dxs8YRTVGtUPH/6jftR4Udg9HTx+q3eJDFEwL9+vFMSP+A856/rxeCtpoJqvxDdBrFpNM0iQ8
TkN3QM34mw7rYTGV0mTynVPGzwTh0onVVwp4se9U/NXQ1oxZp9V9S65a+nXvkrSVu2A+9q4isP3W
CjmK+edLBx/lZ56bMieYkyJv0c+vhhORW9qnrUeYxaaGt69yfGBNcooLOSbHy12iXUtCeslT7KHM
IGfgEGMJxSkSCXYK8hg09pH8QPbWpCsSjRoww4O4WfTradaLK+tzszwDTcUBDrn6Lx56wm1GU5z8
k096/SasgTdstjDd4u5EB38XvKeUwRRIfTXFNc5oYl1tjGWinHC2K/ZyOl+Fwr4UJY2zvuhft5v6
+FawHJ8p6N36aZZrz+bl8JSIv7PJ3NJq7Go/EXY2N/C2tImLnfihhiMgEVBulGUACs/LZDhnp52C
j4wVxGN95MD3+aTOTb9Efb/WqMb8Kel13iOMxAkR+CX9dxuHnRLidix/4znP91ToMisFXf8izM/D
ApJSmb9yKzxjII8U2/mO7s7IhQ0ceBuAtHZEkcZza41D0VOpClWrLdMeQ8Jb1pwIYW+btQSG7nJQ
V1qfcBKB8Ik5W2+hj/bValmSkxtqRy8bPrRyh2YN81UyM3LEpbLLCysjDdAKuS2u9YAo1G6iNXk0
NxOONhy65trvqJAsjD2345VnJUAwGeWwOqOo8HNTu4/Cws1QHRZownhHI9mQMD1xge4YOgAvN3fk
FNO0Efvy3ZIHMnhraCLJLHN4d7+i++fKXylgpcFIcBeCuBnj016k806BMjrR/SGk84mlUir2WxrM
KsTKhDsLyAqMwmN4IdxuiPeMuqKUAZTkixYEFn2CLiEv+9t1YqcN2Ul8QoLJnPeUoq89wXr9S7ri
tbo0JRWI8L7ouggicfqAJEYB4QJTPRuiSA7Kp7wXtaYbqfzo97FzVF8GWTT7BwfXZqt47kZ/dF9m
Mcl3/B6bMSgHfI8MHF5BWjWkw42zgVqfNnlSOz9krildsklAHAP1CSguWr4S0e+uCVRi+52GLpdu
+svn0DpfVhW7tMlGGEVuqbiChKlofhYztYYTz3m6jiOPtsSxmEcoB2sXXvWBRUyvT8PHpNbWoMNs
yCb0aQNiSiYzCwKO0TXeKF09GaEuwFRYauaAIbgcryDoMRDYwMVv7omToLiIzC35U274sQ4kebA7
gO2z1hIAK4cuSahCJYYPWPOcOXpA/Je0tR9aRUtqQvzc4oA9cmUWXp0Q1cn2TAxstkKj0Ru2K05c
a+iEdJVfZuvZJmN7MZtPbghjhEZIsCoLfTcxZ/tylqpW+UeCuepgV0vxFM9tqrz8gzvdgdEiqwP8
SVXBwzspcvwi9vw8D75hR804RYvvo4ecp3kWU6yyx0QegIw+Mn+aQmZPSb+PEFzNacfoUK8GEw5A
OmoMtkQm2tcFNWmRJVOVOIVCHKcHARs8UuQSdX9nDyoV6rmRTmu5R6WQrQ1RIvv8T1y3/sO2k0Sj
vMNpMgF2Fl7eScWaXoFT89w76b9yDk5D/tCWQvz1QOaUYhvEQUWyckt78R3yfsVWHzkl1w43M6sh
Qih27hovOndQJirGWfcJUTjqhWpKtOXDAhp/ZPzOiIwAp4ErQGShe5fFOogOYt0xzJ5ca5gDD/S6
O0524cuSRWjP4BetxQIT0eU73jYWLmaMghJ6yKd+Yw3/psCzPoAFFAuOB7Yh/HP0I1y8MkOtna6C
U7fXum3wRAYlF/pEE5w9TBzbw3ammIwvRcaIwjCk/H6VcADHQz6cytWww4IDseROjv+VUH6s9FWy
Jjmlqj430qiJDyNmzHYB3yXjJWyDZIyQyBV8FM2nRdARF6+SpEQvCa2PJMSeqZtHo9/25Njs7YZ+
/sTLYut6HeG2sUg2eRE95tFGZMK+jB+uqkCIMp/c1h8G4xv41MH6HM7sUhnLpmgJ610HgTaTSLAa
cN9GJqEVlsCMwYlcGStvKy7ocRPKxfLyt09TbYHQhprlpl75dKxak6CXEub0OshNINyFBe+Qk6kj
xSRKKhRCwvzzU90SFi0L3IjZbHiVeq+fa9LoyZDCtz9MoNea+YRmw/yLMnQW/Kjmxhi+qPJgNDX1
sDRJsB9t8RBGL5O5sjHIbmjV/IAy6DqD2Pua/mNgr9pWMpGv3A1ihAMtajVJm7jbpMkFvsbMjEzo
lspTLxZwfXSqw4Ttvw9uaih9WpOkAIzl7E3LrlQfeIVY1J4+RDNwt45Qnw8x7KoOJVL4MAONFHCc
pq+gsIuVTyW7v1NLKrLGrwjIClb7zAeX5iFWX0rccA9BQMsLFH0+vQvq78ADb8DM1yRIwsVnGPxY
Pe0Qz4/RdtI+kcAzuCmguRo1L+X1NPuep/JQsemeaya1Vp38ueErojz5QcEREO3Xk0uhNt4N4Lc0
YeClUQiL8uMa8WLfS8OihhfyiFY8Ez1IMajJUIM19w4dC322ZlQNL8bwmlDo6YvjPj/p93ROhw7T
pAsw8goucjmd0nbEtGQEore403aJWdQPNg5GfSELHl/r88eVtT5b+X5rXzFqhEDQaLtkEuG+ZuPp
SmXygF9+Yq1Bm4F7fEfo4dNzGkQMbCNfd6awFu5J3kjpv3D937MHXrfttjnK+5k1LmPEIgooJH1Q
ZxtYQGqhX4bsFOYDAJ8g4nDawZdFfPsKGE4ouYEljMCglbGbQA0TgJ/YwjCcQOmugflnUDBDeavV
sxe/xe55a2u5ZQ4m2iC6X5ZIMPXGtCI7xrzmU41rT0MwK6hC8D0CvW26BNGgIRomAQep2CDLsBnq
jNQe51W35Gtr1NnCpVBwkkbua57l9IegyjSGJbWYsCV1B3WOmTxDoGvJ/QKOSBsNkee8g6/co1fl
Pzvt28/Ms0ss22PsYcRaPCqa3OvMrW87zkloCHatLDiWuw9mRR3pBRwh1G7Y78kwZ/66yAyTaMBp
drQfdvdxfsRagAQiP8jMGLGidzSDqACzXwLbQhn5WcZ1fESgt7C/5nzPWYpwz2SWt6BNIH+1ycqI
88UeJhtbmNZLP+Hx8weG9yrYx0f50uE3FGnNaMTj68dmGLf1Ef8OnZz+KM6lvu2NMpfLBwZv/Z/G
pFz/FGs51/GtIy4muADz+fOsw+3fc+6i/EF2oQAE/N3XeKDId8qBPMIRFiz+97Wbt0lLsnMj5xuq
d1/fx2NWn9qiIuDNn+yNiKMD1C7ay9iBQH05oW+QczEXgj7JHD8POFZziG4Ago1UJeG+VAjwHke4
iPxu0cTApF909bsVRBtWTw8Ibzp3QUQGTZ84T3Ch1NaNSqFfbOYUsZGC2MuG4dgwuuzf2nY/61Kp
N+CrDukj+cdTQPNc1/wWAvBts5wXliM1O77f3txUsrY6Ok65V38+oAR7GDoXl8yrKn9Ow9uLrzzx
sCkiEX37M7IaDuAaGUEWrKoTco5BodI22ofHfFSpBXqT2jE90KWjtauFw+ZrzKQ2ItT209vi5C4X
LK5P07IpAu8iWxUpOSxWWYArjmlXOpDtlrzgsFCgZlssuWe+eOXdbegBqBkciEowiNmnUkhf3R2/
FZTWejZjiAm94hROIk6GCpBNKyduYpJdR8cBGg7buYWh5bGGTvGTzWbfBGiqoYQ+mgaUh4HjkZkz
yhrVUK13fYgq7VxtH8OgXXY6+YmpMfzBl5tIWjKtQ27x4D1wQBXOb/3GwM2VqbqsUQXbCrdHcOeI
3uBd+eyagvcFQIOaoMftvfjPd2D166yvPHx/xp5Sbmbcq1eJ3fJIWDL59mGTsWVoLUW7lcZ/GvFO
q5gxJFprSAM2j+7afszFqeLHupShf99FLShKmtlGenMS1Cw/M4+CZMM/c0o7WKmgMmOIS0BY1Fyt
Euix2tPzBrB2UF9i9KL0zQhXTmvuvfJxftTCxu6YvMtMmKN9lCVUN3l/K5BBUR8q2Zo07yaGAHJi
Uq28sXXo/W+HdpYLNmCLjjme5wpqkrsCKA6T4AuFdTKp4LxbIhNDnmMMeTFBA1QWYCwtrBllZ7hy
0749or65/Muvwb40OnPIR4UzOdrCMvm7kd1WRa0h22nu+iOJpg+GFUuDBwrE6B0F4oEkCeImqMGE
HuNj8n6KzgG7/JdPwVOmVxTZ8vmTVJrssyVzy6+npqHE+vBKyJCjSxHw/z1RopVpf/KXMXvtELCU
HT+/KWCcwDal1dg28aBYEuq6L+F+wWWKYeOlOS9SlVt41OwTx9479yAfzsQpCx8mNUde24Wbhl9z
qYWxEOxKTuIhm5efh3F+D0kkl4nFYb01harDKQW12WW7qGpUVMk4Zy3a71JxyjTPtowK7i0JJwTY
+kU3UZSwbInt2MH+yvb9tE0uyVcNUqXukzZY5Cn8ZKAczmPvPXl/NNeriY3a9dd0+FL/ZuD9ZJU0
qKaHbGoJvpOIJDTZkriUlexmbKY8qfb6Qh5vt1oESpeKWhVEEQE61hOeKVDyUa/dU0R7nluAvQDG
my9lchgPwpN58jFH7k0FtEDqM3xylGSDvwb7OyRQEBqCxAyg6kPc+VIk4vKocqnf5/uKuQLjThh5
LFSbWwPTHkGanO2y2XsMs9NMu5FAn8vorzFUM6tYq9BlgQz8gysbLQgAnz9r60vWw6XrrmFPprTZ
tL4dEOFFFGJhX/4sUTtPWrbESW80w6L1fU0yb54ZWLxa09GnUth9I8dv/hetMrZdFwDE8XieyThc
h7P9L5qf5AfWlUinWrciYnd+Sm4f7CrUxA0j2zzi/NR+UxS9IArcY2+PEdPaTuOLL5hMOvi9GmLM
E5Cgvgd93WKNMgvxukVGL6VDqlt79TyA5uBDJD+MrnrFLrRZ8G9ap7rBHe5KBdsB/mlmLpsUZTIE
mird3Z9ql75q3cCmNBA2ImchtB1NhSavmGK4VBzmhScYV/vfXN2IW/cOzTuLLWEcq2pJlKzKnj/5
YdGdwy5CoyTZX2YZ1uZVLtcFHofhDn+L5fyWpfSVgxoQ6w4iq/n7ZShdr1v2QlT2zNROdHbfzT1h
aXdj9/dB3PGIY+scwBxgDUwIKGihpuoeutApfIN/Z7GrBQoT3a1gvyRx4JlXwMMhz47bwQLIpW1G
7+gEE1dZ+CmlzhEjIpcuGIkvyLA+I3Tb5o2CehCft3llaCgtMlcKJcJ6Rrb/D98rc1TWPHM2OJl3
x2oHKz4Hzcux2DUUN6xEyDrK4gGIaA/d0XCARE8z+OP+EYCnTyPSZdkgNdI1bMEXpqc/KEmZMGBZ
DVli7Ql58VneW3mqt86hUQ92tBbZdJ8x0AWgIklaxXy9zwkqiSYRm7I9WmMESXMuUank6wD+Pj/N
TVami2ksXripmXKOSeXMWPcBVLzzbuKW7IZfazC9UleT2jUTPr4ZTsAefW7Oou02q34AkdavfdAj
QOJbJiZD6yOgRdKRh+1yu623dQQ2omRSdxvk8fuX+FY3ituCGLUtP5/Sx9SBpFUX5QlkaMrmxE2W
4o1UXUkKClIwRfg21Izw88WEC30VdiWtDhNNLicRNBtiyxCLBlc4bCrwpomFTmr0yjFI/Tj1hbZP
Bb5L86tcGjtJO4TFam/qWkI7QS7jW48ZlgYqH66cgnF8LIUoK1pgbAeseHDCwK+FaZ/EOhKx1Sld
EBcGJ8osnkuAwxBM+XOmQcj91nEPbQgaEisOhjLF2YtRpvSYec/5duig3J8GplXXUm+8ItlD7BQ/
Z2FQ9mZYwiUjNdyrT9Y9ZKQhW21Ix4cg1Tht6Iwqv01Vac9urunWQw/0Vxp3Glwce9VCpO8yOKWk
OUpryvGT7A+HvhZXMZ7q0tqg37DsE2rUe36+Uu5mpft1MTQ3DvuOldvGM19jvJNBshBDiR3UMIB3
0jXs5VfeWF6sIYQV6yyuMZJof49ni9RhDF7DQUY8LW+VrhZ2HgEIh9LrLDr1R/gF3hoNJjDOQAbv
WQB7Slscfq/BbbIdOVsqCg2LZcC0OCCo57VyRRXsXj1JBIAqqg0Axk6YUadZggGdCBvt5JUnm55K
V29ycaX2Afic/TN3rZ3vHw+37HZfXUu8T6wkuGszegQ9cyBwJkgq8xGERq4RWEZQ3nMByJi7QHx1
av6SPoYHu+n1MxG5Ullo5FvCgIWAeEEy09k7xGOKHpEUth1lBsMgI0un7hsIJlVtJYjRw1ihgPCi
CtC9ykZCtmpm9ARGlsrJLhrNd3rBtc+WakGPQNSdXbnx6D9iPY0gLeOVMVpyKPi+tjLwxhWvO4Sb
ZrzIL29hXUQvi2tZg5eB2ePQK4b1x10pTOhGbb+/+BqkbcXXP+b4N8bS2RTmkaBKcxo+5cv2q2xj
tAqZM9AtBJX2cZzvmogpRlilhrY51YxPt++tuVH/QO8i4fqos/ui1D0NR7pv36DtIdcxUYw9c44F
aUKkLvDzpAE/MnLLSutbyK5CGdG6Lk0eSZkmwFdo7YjGRCnbdDgx4PKpCYS3WM/k+vSAlpwL0/QU
ThhKgMfhjWcGiiqfK55LEare8X4SawNMBLaiOz+8dGnSKPfFrP4ouPHKmM72RhkSV+UtTjlZPhNq
x8UbfWCT82BHcpRtJAJY89IdlC/yrFDTR3cOj2bTG/fF4fhj0FIAtoXXWVuEiTNQQt0PAUjEM/42
LTGalA5UUOPHcLa+XuasWTDDLy7PuVTW8FnJGjWhdsrS1blTQ+sgtAKE2Rydvc9hOFbytmBmLnFR
vBOKePksktalIfG4BexyFrbChSTdL+IqWYp5V2cQwv4o+vQiZ9VZ1PjKReZB7OlsDOVGjbgTOdtp
gZS7WbPDXK2IRzqygeS9zfl20c1Nv4UFz6Ybxm1rQupMrL/Kga9gdccvfMde8AlUIMZbpnUZoy1a
89qxEhMmRemwNlCHeNS4XvMk6zg1jnufqiCLtzo72bQpFyM7W1AXEhjE6m8QEBNv9CbhQgeoMGx3
LphwAlFLOwe3MywyOgatqLt8p8gxG7o2brXHT2VF0M94wLVV6sC/SpshZEXEDCobvJlvuxULyL/t
ny7pzNW0fNKAfM5wG8LG9g/uZ90+eJersnUyTQd5ZxgsjCidzvM0qz3SODg/4ydVxfaJqMfPu/U+
HC0K33Cana1Q+ytIrPGu9hxLhzpJoCRhN/yoWVY5Bro9OYo9LpZLv5r3G0Lh8g6qHOGYJko2Sf+B
c3axxgCv6szOqvRhzBQYLVpLlPdok7gBhrEvQFF1g+lfjh8ndQSzf8RpgpwKYcUvzVXGdA2UFOkk
E9T7QoU/feZLbLn3AnO501Sf4YAu2F+5KDjNmE5m/NBwH6AUqSoOLF/ezSuHdz29o+JtSxl3XC97
CLe22xDvKz0P7z+fLl6F+PAq5rFA0oFeBNlakFYNdXqPRBrbDxyQ/89XpoXFnHgJcJ6s9slgPiTE
VZXqBb0ZsJV5vTGKbslqIfsE2ZHdzmAoKXdvkGFKHGpyniy3WY6Akb0HuopU72uqHW9T7m0VNCqq
rmixB3I/uxRzJ63Mbra1rnQ9avSnPHnXp3H0tces1A8VAvU13cn61LlSgtqzp1z9EWT+A3Ik4i5I
TSc+N/03Efw+Im7AO6S7QamLzIidw6DsAQ4nrseCbK7BdCmxJHjHqTK4POq8YEqRjXK6O/c5YhHU
i1TcMTgZQV80bu5WuD/kVJei07CNeghr8GThOb+RVWKwPEox6QT4C4QgctMfS5a7kRj62iEf1RqC
P8IqiVqqOyBYsqox5bmfdk/CSyGBRJ3h1VrOnj1t7jE7pM60TN1v8DcLqQGDooQmSopj/4tYz0rQ
bniXO2goYwukpxIamMkrmFrpisKp7gH92zPqWFa7shgL2Wy1FyujeA5v7UhRiU0aohbXmKaJgFau
5v4JYw81Clclu/yrB+2wG33PHDWyyrLkcY3zZSPK5l6T6/R6gj1q88OmotLUZq46r0G/EdLxtRUy
rwWTCb8TdDg6ZuZLm9p5dUVBFM2dci30DHEweloMz//EJlGIJ5NtaEiaRU+Co3Nj1xtJBWqsWl8g
zoFscfyN4+y63209GADlrfcYS/HNihNOcJBqgYNJ3VJA0KYaWeaHhTBJ0TVxbxRJNhBdYmPdftsG
ffRrt35JJ/auMtzDxLl3ajk8XLs+2hLmlcZO2IMMLwV7DV/P4KNfTQwY4FVyMtFvC4NFQ+PGodOD
1Hsc0sdZlXEjTM5pBOLW3GsaCfnpd6hz9xTjmI/W7niNn4XtMvVruLHbEwYxBqODXBDIhCafWWUA
co7dYxz8EJQGQ/6TXNPaEaRABFRBLN0emFQtQ1Ne56hpjl7xFdJEjTe6GibMnOm2GsCiHs5Vpxkg
cqKJPGYRXSIEJ9NmqNrqGKdroo9A0NQjfo+a5UfNpjDV+ATQFUewOsreAR8s7Xw0VCKmyHviOsIS
QiywUPp8CKdxRu+F6UaAFxM2jvlLLmKhXv3JSkrTYmydztNVzUN6T46pnCz6b19VI3fINe5we8LM
INe4Oxon1SJnFgFVutz5RZhLG/WGOBx8k96ZIkd4rfwlFf425l8bIDie23jl+APVlHvLsQEbTv0q
0AFTvTeS8deAkgurUwVdmLV5AYi9PeWZtwcy7HYn4BwI17l8LFMvNoQnaNGVFnn76KehmPVMFY+3
HJHKGLN0gOVcAWth7enL38ULQiLk5YcqmCzfBcQyBs8Qw9i9SHZ4cZCtqicaMEGDqKE8jvw62sKG
xl6eti1CbKSSou2OaHPBvryPK1Y6jl0qqhNpSxE0NDc4s+s/4cQC4MeTdH3dtowquNW3pBcLtRKs
XGhenf+Xd3aVvYGMCXkyMyztNLFXgnOaA7fC52bXEn1qkcsYNjkcDd3aU9ipWAUWn9Z/6uBVfRPt
+cZvaZKxl4kNFJMbbpa493OBS3BXUVuhYhi3TKtNbOEryicPzMeXVIenjAxZRQH8V4nh7J4SwLBY
/kEXCMYrlReGL4E732McqOoglu4ECnsCrkPAKB2qeeLgxGB08kZdIMj6Eah0mgxN2AdZffD9KvQu
bWF4IQDkGRfVWAvmTEtHjQQURS0Asup/f5X3ypAjumi2lwPA3OUpZzzG/Y8+zG8n+HLVlQIEz8In
qER1mXFHT1Kg0NNbQ54tR1y6copMoFDWSgUsz1M9Fl+xbal/9ji72Tj6JQQnHyu0YgT7BrXYjj9O
uIJvDySdnQNEEogZ6ReET3NzImflhSE9Inln+24VpE5ucVwWhEWzxwXOIZ9LW7a4G3uODM5loByT
S4/37AOSuCOviDsOFmYQXtdPG/9Ni78BjvzVrGbznqyNiPEfg1ecvjVcDPGzFVnw2gFpofRtT22k
+pokx3b/8oSlY0IgfJha+MYU+FWCfvzxGWzSn94L086wbgJpEuePPgf6EGoaFBlDWIwjpsGayqSk
q/DK1tvYxjqA6ckT/WUllIuRgyUXy4GYefThIDpy1hL/Tbx8fbbAry/IQBlo2DnADUhien4A0eIP
5+bZyrU4kk5kaOhP6JD1w6uMsbX6xjwWwcV2TcetRYuQiymIRCl1cN1v0LPehUDMpiijDSp6xae0
rYgSzEBYLBwbqifGVlinSk7liYLn5NARJgyHXiBDNSCP/gIz1kXrZ/ajLCIihHWeUs4i2OBjBsE3
tRs6Mvkn0sIz5j0tJ/XwakjL/7NDEveAdrVsLLz9zEOxCa++IjspXWHj2VkRas3qgaA3nfZZTV1G
6o3j2gXGdziJCGAVR+GyDgTcwjTLMKn8e94ePqIsuxpymgR7gaBB8dOfVFmAfwNEHxP8pCYYd7cr
O12Obwokt/vD9xHmqyjp6vsmh2YoWkbAbkz2j4rQgbbqS6ck2HNKFcTPbQC8nKJPWoP5crtWeJBF
Wv884DHfraZA9YtJcv+cKLgAMPKg2NJbYDjqZ9IOKN6tgwW2M3Akn/lW39MoBmF5IY0zPJ42H4b+
gp4Iba43doFj657glqfAmxlAPpTo8nJIcSuxhiNNC/Xjv+Sv/MnTMMn/7r8XbEqhRXc2Blyr16gc
hKEy0mlLVtvfWR06DwMhIH1PkKYFGaFSzlGbf2whlB+62cyV3D4kYwBjwOyOGauMsfV0FVxsSMpI
RPYMR+Qf80Rud66K60fLlQs4aic+7CcxeXP1zBbC5DUwSevQk3p7V38Irjdak1KhD0C7GTYwlU2r
KT9auJ5NdVv636rJDPAPxVBTyNBv5JdigqqeKVvgMWXOb5hCk3ODWrPf7PnwviXQYyXwUX3hHUUA
LCpFDFmGptXsHoa/ijKu1LeVMFJrc8e0pl1AK92STsDjsaM5wW5+4RhibEoGMy47uXOaYJGoUwXq
8bQ3B3/1vxPM9Or9IekUNCIHRmRRKecZZsgLf4kRBZqJ0fSBc36Nv+8EXYNQrDQ/eca/2Hw9j6wG
+vXzpJ0V3zYZkRXzTzs12ku362S0NmZwQPQc+irkxQI/STVIuJo0LIBjfiNyKhQDqIx9Hhqrl9Sz
B1PRH6F0lnwb/wQoTNR1/HhUzQ5Ezt+uKsE4lJNChvitwRr9wlGcdOlYjrp3IruHVtlaziIkXoKM
nVaingTpcyfY0SNFiZgQUF/DfQGfurcvB4wI4ZyZtkGmdvPLxSnli0FCsD0qZ0p1shP8fIOjMxG7
CVn9OMr7WpRi3kJTdFkBttl7H5mWXb4Z2zy5iR3fYUXmRanZ6iSFvKlCD/WaqzaCeZnZ1hcCFmHk
qDCOIYYBwB5GbG2Bks0hPk5Iz5E77+uonzR1I4TzHOzbrZ0wAKTCScPQ1Z5ZQHOMyl10zuJC3ufG
zv/8jT75vFuqpVAjVL1oqkDaM1znDpqHq+DKcBNJMPisgFCh5t+UmiT2YJyJ0yL2RamZITW3kuPv
hby5xQHjWkRO8CgF+kcmz/qSNFrq9UsuHlBQ3wtgw+3uppVtTVV9+jhQ+Vv8lSv0DXGejyR/xhqx
q5FC+JY30Im+6Cgeu5nHFAm7QnenQLY0NE53jpwOstEIHQtVx7RbCl22dcKm5qCYOpI4anuolA+L
WN1LZbZLZDA6yghiIfVnW3BvZTrDnVFpW59vPL83pc7ZoEmsFHIvWe4kdMm7cQOIomg3S5UaGBsn
Zddo1z/lOIc7kNg4XsE1NnegOGcabyAf+5ZEMCptcyz8EFHLIO7Pd270tiszWD2jqPwQFF7+SsVw
8HuFqbY/WlDORKQ5vvuI+Ht8mGBB+dnpEm/6f67fYHSzAXn+A5SBaeWG7sdRMCYiGl/kC23xs2KP
6vYWZ+T4Nvyu5T5oF74LJvMsdckirqvQr/8bZ/+fZwq9FMJzpLu8Uayq5I9ePEVV6CaVmMC5hFDg
vYrCeax1XOJSFk9yT1/rcm2t+eXS2zrUKYF6sDxDGDKKNYEsnnMRp0ZCpEez4oY0Bx30S62vPHgf
ZBpLK3f/yccoOR6uNny6vlHqd7wb6FLjY/EwXJii+3esux7gIWKBHBOmXG4b5k/9t8rmm6E7yGvi
P/ozweTNErWXQ/f2anHDmmMOedq7KOII9wny4/wzwI9c8PNZmSAWQepM8OFWF4CcIBR2kkPx1ZKE
ITEdWmV401Y/t56w98qKKBWOzjwQyG/h5gDuK0CLQyDOqB1zi8qBjcqj5dDDheRmW+PmS93Lo0fW
AlceDUNuJSIBC5MnEzgCct+vyaJk0HCJQD86XFLerh2XaZ0hiD0R7x24So2mgsrrsg5WC5oFRwHs
HyeJ0H9hiC8L6GaWgKI0UGsVyPnn97BRlEa+pdp11WY90i7OqMWrokdyf29N1skN8pTppmxwB92L
LZZ225Lv64Er1oiTKxgK+PoFSH+9mc1x40uLahCX39ng6C/b5vfnunvUaLOKeidX1WCvB3xFLehA
vdJqUEn7lX4Rm6vnxzBh+PTy24usapfwz+q65hkuVu/A0GEBP1++WREPd8186WpJCx8DHCqKlkve
8x4fSsOt41ZVWJd2ukBNBR9nWpeCkKddXn16cMxMDQ7vrgbzZnoQynMo0zFLKYwbrtvQd377SXYQ
cH/XHjOvAJ9OPvo8S2nbAVPHJ4QOLopjt4zS9M9bkxnw9dVAgOAVQzkCl7xIlDnON1TKXPOAmImC
lNPTZXyv8El8l+xKyEuMW72+pAiLRNHo4lbC850i+i+XKmpc+CDcCgKkjBo0dzSQKUknu2iDiBpA
unN+C8mOChA99pYMKE8cBn/efp8DLpOm8/X7uPd5EOsQSg7TD6pbENTQsgiBtHaQXRhvaKS/pk/u
uKBmDozJM7N1xeynqLygOtWZcz0xghbhfEGfagJw7iFs+JBf3H0Q0V86X0Vxf7NrWO8aB6gjwgG/
kb0rIoNXnHJqY9RlY5H73janHZsVzttK6nulESDvh/fzGYinKT5er4AcFVLQmL4MFXKslGiws34x
yG4Xo6xwam0aW1scR9QGdB67jGpp9DTz4/CxY6JhUd52Y3YtgFp2twCnO1lJtHBvbHiZAc0YwJXN
TnNCusoo6AaiWw3nVULcnC8MHHnxJ+a2/pIS/b4k6mLxJ7L+EKm5H9jtQnPXk/Ujl7fVfNNPaI++
GCXVQ4MR4gKbhc5o7IxTbKg0giRXA9qVtgcHj1AaLYco9peCRefVZaJ6xSm01umXtjZPlEXBN8Mc
fk/sAyOdSDNcryin8PYYODigE5XE2n54l/QXhNBLTOuPypPEsoCCX8Mee7UaWeNWd9PaOqtKo1va
oFYkuVJhzX+j5BD0oNGyoBiIqyvzcZfiLWdJcM82GU+GUrbtf+mKmZjHlvrwEi1JwFVqkDkwxp2N
OmNj0vxNHsuESpNvEKMpc9w4XJdsAE9tyxe4Y0OqT1uhG8yxfZwrFgu3p5DPEBlz+hmZZRPDd2Ve
Uf3bduwAoJRXkWz/VACcYZcSsA3wMn+z/U4b/uMnMuqmvC0quHPj7blml5ljALyiq4NSH8HCTWsv
CmkSLuDaZmURMCBoBvNB0Aa/sp47IRjCpKr9F08hDZGJu5/Li7dkXNMX5UjtM/Wvo+GNhSShcWxq
4qNhOaQ1Zmcq9EBEQYdQjonFkjEUCyhj/KcyqS2HTaiduta74/HNEecr+QuBY/RaNWl1BYaYwm0B
6gUP61OLtk3McF66mt25uOQAtzIhHbjnFb4xwyGbLw9060a9eo1lIHQsTNHfGCfun9gfK6UU1b7T
okXI0dCiJaXnMrONJRDqGPfWiY2GzaU7zNZ6lZm20G56FeEl6gWun0ex8yQA6Vm2SpDHobvoD05J
H+AKGyT/J/qVc1wuhDxKo6YKr6z3hSAPgJvHeSZyGKIrHZNU21tmo8Dmi7vumgSrEkLfiDHQ2zNM
oEwFhW8wTZ5wN6Rqcf5ZGRbyZyWMvO3S0MZE7sZuwyNnx6K8w9hzAnhW2VaEyemFj8dE62TwlFgd
da+A8UjH4/Fk/QhSHeE9U8vwoizJdN7edBSkcr0lajotweelfDch8MKVSE+Ezb/kvmXDfP5/1NIH
7u93PAvrcFkB37bLQdbVtXqPhpPX8vTnDKaGhCgrRwFBg85//pJFgDYd26iaQjUXjgAOsZebRJUE
H4KkzyMfS60IgPlKFqInDrfuoWbKuGFFqwZ3zkdIQO+b2nxxyIxDsfJLrgX9l5GyB7wePIWk1U9V
IfbDFJ6ubCSkG+ODmInE9m5DOOUTkqy7eU8+Gj+SzU2oXR/QMMJMNe865stSvzplTRLnfz8kmVT6
wBE5a0UJ4SwZQfSnvMn3VD5707OwIvp54AuUoKpts36V5sX4vmE3yNPcK4JxHd5K2isoBIqw3YT1
wQYd8bktWdJgaNaHjnpAci/560xbrwMP2zoQfpUOy4zfd8LnIRl5MCWe+rPySwDP/BSOGo8VQKui
+OZTvUSBZNMPDTd88RqfLoOza8NFWiSU9PrK3/R1vc0MYIhktTOkCksJ6u3RUg0ajXKBG7ZGXCPo
y1hb4X/SFwuaaffhTBsaCxinaQw/tek5U9GP2sZT2j4gWbqxSL/akq9+3O+pH0Os1/hJ/XG1kC9O
b/EhNlw18Mc1FZQ7QcJoFS2hwEgSTP9OZG4BjsWd4n7Gpm/y5U4oK8/4O0uzdPn5nzWOB32rsEbL
FlLnJdp0XEZXX3HpIWtUXeCqyG9qaRM/V8dutPjbAVf1lIzOiwRgULtjlZfd4k6Re7IriEarUkOZ
e5BSgzXIllUHszfu2vKr7zJa93uqTXkHARC6xtlW4UqmYcfzbFPBZfx/03WkHnPq/DCpqcUIojlN
llJorUzTnDrhPBST0YtJ+Tp+CS9kA+wFDQUYSKUiADDGx+aVgBZIG64vikqlv5yTt4fztO/YtOBt
0aju3qzYzdPip2b844PoPpkL+U1tF27FNu3wqYFjuyHKgZ2vc3RV4wxqB4Gh/czRz5HbcyaV10AX
00x8gQfDaGrWE3LuHzuC4dDXAHpA6KvtM/KadpnxJQwiFfECrk2TRdfwTGjqcudEn9X48nXsd56m
1GavAyBZkQDEicHTDNtWHD6SFxQhm9zUgrxgnYkntsj55Hllh5t83bvOKFwUGtGC1G/IMJJwSmbM
DAk5hbxo1I5+vNqVVCk5IvmAlV+o2G4J+fZw5i6eFGZQjE6xPZcLyNRuqEIslBikePZ2RA2RGw2y
kNMaFMRCC5rO4MHfS6RobubzEvWlNIzjy74a7wfCVV8D6dusPgG690rP5GCwnGdGtj/b3wqwPUqT
Y5YIh4cPCQskFt6vqj5CLEjutSEO6uIQ3Yrlq+WWEJy9dgu5mGBnbF28IqzK2kQMqOBrf3PJxakE
L5YVMUICFH8C1UqBUvkWxfi+pUAP6PHn1+C7/T2XuMML75DAnf7Dj2LPz/LLmx+Jpz5nuqUSreHB
GUUCmY2HdfxMsFbkxwZggh0jHQnc/igNYmgYECfujRm+5mj1ol88ZECq8GMFHYq7EYtSnvErNXsP
a02DjU2pA+bvGrTo515FN3s9v3gbYpW9gArJqSUkQ4twJZSyP9LT5q97ajxB3SErJXB/pu0TtgEy
PE/WWOGk4bnGXgq2z0DVw5Sh5MG9BgGsTXgUjEaNjE0Ilxc6sjpyD4+jL1J7bPopzwp+NIUsv6QS
unKY7JG/1SyUDjv+TKWuAYIFV4DjyMsZYVE4ykeXGrvYeujg1ZcbdznLuACHP4SWc5kVmyUUJp5f
Ci3YYleuAmnRVbFKwDQXMAqJuG4Xgj1JgBd+vEVonZFWYYx3w7ADqVUB+aPhZ89bimaGxWZ11Qs+
+GVgosizC74x8s/3vbuJ0R8Tcpztto+WjOAwNt/KW3tFO3QNoiYW1QewqCdfUHS500YiMq5utsIw
iyF+9Fy0H0LbB+6hxz57JPrvct8CGdvF4z+Haf0kQJGnRkWu+uZIewLhfp9a9t0AOCHCuzKv7GPN
rgE3mSdOW2sJMjZKRb6HT3lSuMlo0/M77I9y0K48IEKN+fwweVmuzWAiju52CWNCmv7CQHJdDfho
XWJQ1SujGxrELYi+yw92KaHqZmDuAoA+/7Ec/CkoQUGqzNLj1ntQU3Vtn8/GsIOprp8uSEItRmZO
3IapNtdigcsxMm7AzwyO6h+mV8BzxhxKvM64+30r1RSoOMeGAHS2uo3h6agxPzYy/nvBTwJN3Jdi
V6Lqr2CyStXa6td1d/HFmEIlwU4yzFeCoOuoQxTinoWJIvfh/SEDMZtvnN/x1LfSDf4bMHlhRx03
4SHkUJ5pdy4wFXF92u/KM+nX+06ryxtIBTRLjAgIcJPS8+iKv9/D0bm4vP6tNkrMCzor67laTH0U
UkrSIuIRRRwvqr4HxRFaEacJRc7rvOdh+a54w0ULXtlS9micTktWTHQOLfF6fQCTRZD1ny/aLihN
GWbBmcMTGEHjYNwVwPtdR18RHpNI8qXr8y/Vb4CYZn6+xrzltQteLneLI+/Ok9vV1oQaJjULHazT
WikeepgwM3P2zFR5Z26wjILMMj4gW/e9r6iL4Y7F1apRIgK/8nyfZE4+LrZJj2PBtiDmodwEar5V
Uu+GqRpwyMFwvdxMqk7uN4DAypXf5Cok56MHn3D6JEOWtNOUYwloZhjg8Oc6IDkuO0QSFsFYrf4S
TfdkWYbpiDVDtfrwCHvd31lpuX9yp4J2pyXEgzPfIFEOJetERaij9nphbUGOODzWhEUhjNwUZvAL
dI6S88KGnMjSCV2gUdZlmwLBsEhksgXMquGp6XwyWh/6G1a7hWUomnW3y3iYGy2M6tWZr0NIsNu9
Ify7ybjNLzzJwPQnNbVtmZiKmTTk/coxRAympf2gt59E6psokNzlgKJkkp5YF+18SYGOs6i+vxtO
jTrV/pB+gMLi79E3pITw327AjORtNzZXoHqxUC69ekq3Oua2bWPHoiVGnwkhOzmulK+cykwAQRsu
iWcraSTBpH4SLXdBBqc+GTxrkvvj8DaswqxZSy2c7j5mDt+0xa+kKviZKZSknugkHTJH5Y8yY/Pt
RmHQdu1Q88UTyrNaR9Vc33h26lSUSsnNK/Ka/9Sf1XmQf+mTa1oIewVRglSRtFF6P5+nSF0zkhly
ct3FPEuMw34XWu0OtM3Ob2rNQrf7AJnYT4Qmk2002scE9SDGyRoqPDcXfnwZYvAatTXHHxPUTOlj
ArMfqOaky9GXXyA0DRomXI8sbjzRBDWYUktgYh4kzUt79Ftdi9ECDrt7/GrUoAjVHlNxZb3NdlrB
UA46jG1Z/rCxEDH/Q8vSAV44RDA87heyZjC6Rrcw6wpbxAieuRK6E2jGPXLu0OsLyh6TrOP6j3EL
FVSUkxn30Q06dTfFp43hPuQQQUZMgs0NSUr/nI6Kh57/HyI4cFiVWsU81rg1YsEHOSloC7k2cjiH
ccrotIQz8S8/Pch9ACt26nxE+f7syJk0qwP1z67NxKHMiLYCVOEKH5KEIHzS9g4qLsNFueLoebyf
n9N4kKy7LZZCghuVeXN+VfAgRyx609KFHplyvUZ1qi2hJAHGS7X+RZcaoamJsDfBb1kq+gf6rHx1
MFVbyO7EY2OkMEvBPRMqsmmItQhHSRFLw7UGsZHM23+6sAF5LWLOu7w+eS90GygGtgm1LW1BzJXR
m0qyDwDIPSEkFiQJNvCZiTOLE9z6KXcnt9tuhtIsVmPxkQ6xeAaGrX7/0sqQobdgtHf4RHlfEYkk
gwDC1OVbqRcKKo2Vt658c1H9VYiQqHLFLGu+2qmEVGpV/3ph3jhVGxvnhstDCwyrvpOpDU1Ufz+R
Ae6yNCahGssxTiZznSW7BFJUv+faHU+3clO3+5K2jAGEd37kBjQ/RnBgBt62PjM9CwC7pT5Hfy1T
fwm6hq6VZE6GCRuS64o2ZUkGYteOaMVL8muEd+jl+AnC90a13LW57pCrFt+LJK9v0Tt1Zcs0QStv
j8NtPAPrdCyNne2U70BhEZBLn/OsLQ1z8crGtopVjYoC6t5hpGUHwMKJSewxivP2IRDrv29wz/rw
BZYELrSHtLk2VVthjlowKabSkBC0Z4MzZTSnJvaARBRadEPmyI1YZkFlzEPxlKWKMOpoybNmJ5Bi
2l1rSp2wDZAnINyW/w8HAL8kkBvYoROBRs+sMtvprqFsBmc6JsAewH+6vv9VWd8LLms1o9tMV9cy
MuLwd82nLOUUj6Vi1rMCr60qBXXRwkiPmyNI2+NIpynMiPVY0AueeZ5PqlnRPo5GKC0v//+VCosv
wPdT3HaACTIXpLKONtBWfnaXoWd0uPJzqH+nYFK28GPCY7F8ESEEzP0VPY4+qrByNeMXlN6UDMbU
O6uZeisIwXL6/FwhuRstRJlrBlr30hmxIuIWtQrrRny5KpoXB+PcXr4I72Nlr4dyuctqhlL+dfcz
/bI7B/4bJfqem7+7QO9wUhXJLLOU2cWJFV9Og9ccld82tBwaeEOvzrhkAJwTGUck+fYPBYnFPbEc
D0aQPj0EkC6IlpOWKOpmC3f8oB9j5qLN+oTseC036ASXk5mfVjHZlYSjYYfqvIp+Cm/CRo+DXSft
84p2FLmJhnRneA0mfGgKAiTyOrrfFevxr7ttNOGyLxed7Cu9BhsYTF4fTBOlNz9NkfnuaYdYrAAy
mJvhRVc/0k4i7ooeA8y/Uzd4j+j9FP+XTiBD39d8VMyMxqdPAywd8kPUcjQxlTSPmnBrIQhoTyuK
VhvwZvYi3Z8MkYa42ibJxgAzw7OeKXmQr3JJsh0IT0hjAcx18J7EQatIIuouwWL+LXISmvdh7b9r
T+//MK+0oZb6yyeqHOSbJuVhNduF2b8ko1tmC61wsCBd9bCclsavpbL1SySXq+ruGO7e7FX2bz40
0uHd24iJdbMFotKTDw2uT3O8dVZKpFBaUpZ4S57bJRsCPhPDgPoh+GmiidAHNNkNILsILaP0uOrb
HlSD5v9uUMzTdUfrUisS8uJaUlwVX7drie6563qDu/6iP4fd5NJuZlg6VmkITS/q5J8JthjXZwu/
3IAnwa5pSYg+k5H35PIsrG5VZZYPZ5FBeobphN2Fx1TH0tSHhQRbW40cPTqHi1qFWDwWyhwtiBpg
KFME/JwqxPByfuJiHp1taijOsJ0mpdQvzCMyURXK785C9GzGLv+RmrEk1QTN6jHXhmBs3q0rxVce
AbW1jxRXkp3GPeXxssoCHCuSoEoIPm4EP5aXdbHqDZnUlU35PjZdUR7fYGekhrXGBD+T5RRUaJhr
3/lAiavlckW26V8ryEyHO7btKAQpjailefEKznYRsiCvMG8v2FPwQsCS0b1MEZrTUKmZxJh+CcJ5
ENiv+85QqYipTFez6pD7142XgMsIC9jvjn+5eZPrY3tDfLfLAQXI6NJ657ql60Bpx1xgTz1B6yvT
Rlrj+oGxsxftjHuioCIvdCfXV6ZKr5HQYdpF1x7IsqHtuR0jn9kCgiw1kMTzduk4Z8jPdXZWP2VQ
yw/xPZOH8m3BzYWAUxlqFjX1I3UcuYNSJzoTLUAyZSRuUlxbXXTnnY4AvOBaH1MobM8lLJn/uK/+
NpYAhKGv0V+xs1+h7zEIVigNaAacQ1l93MqmxUJGsR+9Jejasb/oN+GhnECF0OvF/j6FqGRcRLfW
7WisIeZNMD8pnMXWHdZl1L8eiRU2sGG+d4Cqh/qqdQh8z/S8XSvuGTsCZ7FzNiIPrU9KkwJZvEV2
TL2EZ0W17zUiBhvY35+SbVaYtr/c7berzMUQkk9424hNb+vKmreR6esaT4mtbuBRGym76o3IF+pB
MqQ0RpRG781jnuGWGIduhHpFAf2Ac8MYtnfTBt3b6XQzdLZsoDumFSEQg98V2OF4IRtIoCca4WKg
pV/KYDTtoL1AG/xCRalVkLmUVr/dW1ttGcjHtThGZIiN//RcbPuYbPGtZI89nZjH/enMnP5Fd1uY
/H0J3exFrqMHX6GELbE6vndDoi/PLaJQNDh46x9UUG99O3F/YxnlFpCYqx4vX26mXlJMlTmB89ji
4wemm+W8PcV/T6gqo7W3d2B/83oInN8ywxN3crabeXybrGa9VYLJwXTZaIq4eFXOu8VtGrK1Ya5A
oEs6u5T2qE5NEjUrX41kzUp7guvhBr676UWONX1lp6N16QKGB+QzL8wmeGXCYOXtAMJCaJ2+w9F8
tLg4vsW6tUiz7Tz0TtL5OzC+r7q+HCTl/YC82qMJsuYw8is1iMFD0nmsf8dy51ROX7y7AhUqY45R
pHQyxe097Gf0H6bkmb+MmUPVd305u82Ec9rvNALusi/0pxSpv/1mpMUQNRZvX4pj4srRQm95hwmI
JEUCqwt2piFQ2Zmiul04Pc2ZmhTEdWFtWAh535AGo7lx7rAmez6wohOPAfOCuZuFYGkEN/Y55fmj
MJDjTRXrg+EnBk3I1U2ex0/rqcRR4ZKZHTE+Em4NcNw1SaTCMlF3a5LnCo+f2jzR7QR+wREa9U5t
y6flcow6CpJQZN1BwIqAeaHXcn37VmR/2i/65KJJhgu3coPpnCoUE+KTR5zKdEXOMv+nzUdS1BR6
gmCKMUijswTX2wOqDXRN8AWgXw5v136eLvpJcyCvBEX9+S09A+p+Q56uEw42ApBo7kKq7Ws6lVyX
Kozf6AR1Djtu8APMU2b2VBnjjBCB+1jFMe34dFBT3pGoaFl7VoVAf7Rgm4C9HAgVmbhLbKny6XYA
9nfl6m64/PT3S07CydiL2wulOOTq6DYnXEHB7xhEgBBV1kKMgGCv41kbzn+ifcGsgfwWDcLhGhVv
s4LgMJJUHtZLr0KqDStI8sx8hV2VVfkTRcyH/K9Y2evcjhxgR0s53GaPsGmT4B515Z8FfMTD3VkV
ydH8+WK7nLP89Ab7oK6rseViwhwWwPJzXw0ZYzcG5fLPvRW+5PoMSpodcq9bnoJ4jKdh+OUiHIMs
gvJE5E/Gyn3oIpuJx0LZL3cvzn5MSTC0t3TB764wc0nJR3lbd3nwZt1K9SRcic9u4ZNCd7cxe8KS
dbJym2uTEODri9keIaBDqKM6QQYbyJDub7Ja66CivADi+WoJvefuJwV4PZSX3Jy+gdwvmW5/+khp
ygN/VIvPungJ/YcOvYCG+lJ/WEo99IwDYJJYLGF0hlPIacX7OkkD4fi6nAQDODqKuU1XnDPF+CDp
Pxip2HWebNO7hVZUE7eyMVjMW5ZhJKefB8RAgYrOfJFf8aoveqMMYpVmPq9oShgHjrRf7u9EKEM6
HMYhzHs/flmMVt31bmON2i9PgdJB3vJpOLhHQSL8gFVsfHLWA/B+r58yus5acBIfYr96+LEQOhtP
7i+K369BH6qwjxY1zoemtlTNckepEFi/3tNu5Wy2gB0WpgkoSgjN/yeLo9/GFBRdkk2Qhrb30ao8
uoNplKUko1oVu9GYkHgECgB6nwRCUU/ehU8DWaohzhE0hWl8j+33jzMLJWcGb8yvkRR1uhubmtCx
SsRPSlII7kxY068EI6mM2Bdx9bXZTTBAWZ0rrEb60odtxq+uLKM2Q/BkYar5XfUBioVT9oH9eyP/
DpB9N02a882+kJLqQoy7Rr56W2MOGQloEXI8wYmX/uRVLxv0EwVhh1SoVvhqfev7Jz7dYnHvhRdd
Gn1cDTIfMVFEB86H8xGLDhHEa5taC4xjnDwdR+I4Z7p8SYCvi8M6o8kZi9e+o/pGX5WirvYe9Yxc
kgAG8LpRimy4ruRhPMRPWIUn+SESpeeC5ZppZzr6xIo4zgyp3GSVPurLOSZ4nUs1yw+vlwSw8kg4
XwbmVyCwjwCnmrHhKcIqPdIDjUduu31coVBB5pWpgnXvaMcT0McAKoDv7f8c4Ny3P3WhXSOSUiDB
b+QV70TK7jG+JenwYmxtabJ8dmCRHeUecIFKyd5+uowJKd/QMctWm9wrEckehKnYTGTSQIyoWaag
qJaOp+CjJbc7CIAeTug6vjWqBdOUbJmrvPmHLd07dgDNEUqAL7FHfhSgjUzfDDpIsi2JJ/RhET2e
F7n1EHzPLFX5NCoRESBYWE0fOWLxKBVK0p5D3njU//nLIs6/2Z94OYMQYmfIEDobLAmurb5ThUZe
gpRI0qA7E/ygNmBTaVDkDkinn+IBb9XYiKujWlABYrCvkNw17+9qP3vVylymr+cxmaDr+ohFkoP/
G1Q0Uu/42zAwwHZd+fUnOyVbprtrpyxH6aVGXeBvtYLl7GcFBRwMXn0zpmhTQYDxaQt5F3LpggzA
dyhUvrWyjIwbauwh3mrbq2btChxbJqAigJoKaif/EM0bz3hdsRBvleSEDdbVjiS0yyA8XSJpEU4U
VOdoIc86pnBUyw+dNzNFJ+ln6HSSOriMyYvvowOVBSxCaTTzfKKaLtfkJLekc2uFm3oxvpYTsZhV
lNob5RaWCALBQOE73zZfuf1659DoICNVOrCLqSa3HVvzVMGxVDtryBs7JSfKCbZmFYWtwvb75VAb
oXIsfWLydfXBuK8p3fdihE2P7DaMhLm1xWRC1nS3HnR7wxOl1N+XYMRHfY2alHIcMJompezvVAgN
Zrm7rz5UyYQ4WitedsY4DGyBYEtZfpvSZkIcQKZtnTekML8Zuj5yOLVtq7ys8MFg9D1mmtoL6FjS
Wx4jdUE4eX11eVqh3OMGR+glh+tXYQgd8hQ5V+MIn5zamr4q+BcPJd9D/6KmnEW4BFmCa1mzdZP6
Nk9iB5DOzRCEXYQ/91zBgPKuaUxCNsJr/4w0sArQ+/exo8tISqSfK9O4aqxnvJl3g17vyXl96SiV
0EsNTWODFNtsrlRtZRG85O2UOcr8PEzNHse9j5xrKT9Yt6zNlrhyZ/MrD/9UBAoAfBY+HGV/poTf
NDSqgVhutmCIxcwso9mDzo/klTooi4tWMuBJIgodp23c8OFTyqA21xKDFH65jt22JUiU7OfEVeDR
mo9Yp11lnhiY2m78SKkMZUn/c2oUguZjst9izGPvni9DcBRD4y5nRmNhLeCa7pAKixn87oyoyrow
OWin1aDZwrdFit8FTs2RKf/tmk7XJMoc0gUgAt/epyLBBXmW0bHdomt5icpsAi1QcgZQABugtG8d
VZ5RC4amtzlKOIEQaKq+ggfYBebjXWqYlEsL32EiUQCenrg/rUspPgngd2yK5QYdSzcUK3uCLWrk
HLRz+/GMhRpYGDgiqGT/7P2NVf54zc1yVmweHVMZe/RIPYqI9Ay+DfJRvzazMgmYrSnkAo+Njp4A
16CeNKp4W1dg3spfwiKarFrvnkJOrsOtBJq+2hH6qcoWSjP1oANCLErsUCWo9AOfvw2/vzSOmsUW
GjXBxmtcJ4SjZ0ax/m+iZLrBA3fcltby8DiYAhVJH41TXjgkwR3kMZ1r+14Q+jN+dSmhwty05xs3
ig3EIWVQ19lWLLKO1Zpd0tpn2J8cz3E8ucdOslb9dIhWJ4yv2u1lh4DherGWQu/kzV4Y8oHZRf7a
LKVC2lVG8D0LCuQkZy7NS12CZQT4AJA72SgGPjDl/SYPxgmCWVSNK+RItUKYJZ19W9deANIe7IOT
w/LOVP7vFnwjgcuHfUH4MKhAJQERKPnsKrruymCOeyzLmi6aNYH5DQPoIDVa/Q+9SCvrFMi5/KXd
DxZqopislDdribYnKsuOxOGH1OyApnHJgEudK71R4BifJv47raU2ooXIQYaIuCefmlPp1MxYqa65
WAOX/2Gd+ZyRtI4b78LbPPoa1MTft+FdiBiNd7LUY/8huERwNrqrquWuBx5dAsOxefjxU+qlCjhv
pZU3BOtoOolyWjXj1/1RElOXUC62EL7kVbmfas0xYKzt+3fSIrD02YiGJsfOuQ8FSmXlIdBdrVP/
zelez/fbG8/DR7PAYXonXGUyrQeGSazwi02cSvb9oUeWNXsIlGTYKXfyeyUCRlEwzdqbchtyrZsg
3rQ/fUJ08dxFsVWrnI9c8hGPsNmFZMm9jxMFPzcKDIjbT7uwdVX3Dwcg+6QPB/lj4hbVjKDAuUQx
bkgPDW9h4AqsPyBEo9KEPvIILU9SaKh+uMthjvsJsV6YaXyvm1KCxQYCQFI14mY/0N7rEIV/9q16
hKV4vJm65jPk4Ltw+klUjFpAGQoMsa1LjfbJNyVdAs6gJJTRVZQlvCfgP6FeKqRsFV0VFtDPsQBA
tAjbGzlBSGIK+i6cF0NW51la3XyM6MGhJON6VH3kgvagyxZHbZ4rYKqAbpoqb4hMsq0yUbWZ+ewD
v3B2Xe1kB+IBm4KTBTsXaCA0gTOZ7gLHFFB9kYaplZBFmaJNX4MLYPUbrVnOtydvEm6iTc49g3me
Yl9hrfDlGmpvy+oCT2+rXn3mPvFjrP/1f/XSWGO46sEX5J56TLt4i6q/+Ec/Bz1hN4Y5iKPKE17o
5Dn7U48KNAlRJpUO7OQKdTO2ru8a3HwtO05w2l6m5+feqQRyeOJbjuTsx1ikbMO7N1no01uyynon
EIpvc2B4xAsDtiKwwza/Ibvm85mZ1YOMEA42wENZ9R38Zu8zDHsw2E4emTJVzM0QMZTIL3lL8wJi
mH5aZ6LPzcH4Knqsxeu0aobxX4NgiL+rJTOfrLWxEiHJ+Um/uYtpUwB1U9o/u99T33Cw8cYmCaK5
qS1EHqLCGQJ6B5knGOpL2jjlnwuz5Vf0wxkrWug/nuFMW39pK8I9HL0Mz/IKrdfB4DrFrBw6kk32
4aFZ3Oi/+C52WoTKZHF81xuBKAXyxqrAvkl7sfLtfjrYPxTzesj7jKyPdyAyVan8QBCx0kpJVOqo
hHMo0mVOI+ay9RMkcUtwKRuxk2ikHWVi5nO2kakcywJw055N4YIU9pSKamqOY6GNsSRRheW68e10
IaPn7CazWVx3ouT0AC/XJbn4bBS0sTzKjzzNGuFIyh1aWFrEHblXh+ndOlVcjgoFv4a4+8EJF8wT
WLOL4McIH+tx6Mi8kWBBJ9TozgqBMVlfhbzNmOyOqhZK6QNplCUCEk6xMYy+lRfcQBEbY/9K+cA0
QomnbFeAZoAGQwuk+mKRdrQw6q1cKdr0pJkPk6jLL5nVkY507+FhavlQzlAquTx1GrWoKGNZNwbK
1E4S73dSniPkYQgvvOcXqrLaGJ6OPsm9fBSUTureDu51f0rAtzxG/SxISHA6COKCg0dWMA65XT1r
KwCF4BeZ5EQkhMY6qLZoB9pr/skLd8pckRXCQr9Vd9y9VLQz5S2nTq0tygBjexAcLdxq7nELNWg4
kDeyPuzZU1mv/dmzS9nieqAPRnnmQWkwz6EVtlMeSJyU4sl0n/ro5aC8uwgDA7BVWlCEpnFx9b3c
jRUX6+Q+iMBh8MNlIH09prnEOKi28RlaCjUUVnzSx6FLHbjU4Z9h5i//6UCQJ8V3vdSF8SImZ3q3
EClImRy4KmdPed2C4Xgn0GvWKi+ZPB7urC0/dgQgFvtbpnWuhWhktH1Py8KfB+oraYgJIKEKoF9B
hWDMyCNN0jkWz8uWgmZrg4FWEK+doQ7W8aFiH37Rdbglknref3QqPvxyZVhNo0VLOajj7qZyhYcU
hEaQD3dgPyn7qJeQQ+wgi2PNsmLe6z0U+g0g0nq/1ZmYQGhiSAMeD7aPXUP+hhFnqutxfpYyzIit
8Stu4XBwY50UsW0wp7QPhIJ47fLNs8McSkRJh/EDuW1+k6e0+FY3yS+kE3OBm38FkvtcNIZHijZU
kq0nUglZ9mOajncTwDEITrV0VER/6sSfwFgCDuoPCUBhxl9pgEqTjRNQRFl9hi/i6qPA/4t9xJTv
AXo1pti5G9OMK9kNAIkBvvoE70aj1nbjRecRN2N79J19JtEhezrCMixUchNZiQzdG1YA1WISZuYu
MtTAzGzdEAwkgBWsZgR40sJqpv6tJCMYfWS29WxrwVFaHmlaSMcwyZgFMPma5LHCQ22O3HqWAdNB
j+ilY2xAjv/sX0MYLVe9N8mtReKXb1MD8dNXvYxDk5xlKiW4/OR9AI3S9WBIUUnw+Z2AxhCf3yYO
dFhH5/cDCQiGi9SzR5zZfJe6rKUZZGGUXf/DWRDm/5mIJ67vUzddjzTFpP1QwOH/EtO7t3nzZUg6
JGkxb8glKDttj4SgjaHHwsUJV7P9jxogFb8E2x8sy9/SlEsWX+cLjaImsGAdsOwE3DKtEmeAR+AI
be9NN3lMPtc1yqXyJsT54jtvInebZWYrrADcK7D7OMYWgu3q7X7Jy5iKVMFdy68jzfqdzI1GMXGy
g/B0sUdhXA6+4DfuarPNbOUtazLb1gKOsiKDyo6McyugSsxsoEjwu1IiAUVo3eFQOyOnO4Gp5Nr8
hOxF2RSj19oXc9oazM5d2OVkU8YJAWrRz8LFBzy2LCz5KlGgxmcaC6MeUKk85zwqhxeJaFrcUbnq
85su7bm3YXccowcJMU38UBxGwFt4bhNM2q5DANzbzeIpgyZQcaIY7rb2K4rCyMb8GiwvOafDVria
0VN3rK6eNxcahjhkMab98Q0Hg17JnQRTNj+o6jpHJzKKyT0Ylhjlus1oym7uQ8+UGmbZ0amO3xQF
nZJLhYmdba46529ydk0E6ZsDGHuHYq3m6bi8WcnMBFAu3j7GDZ6E5MfhkQuyu5Le9lAJtaA554ot
XgqP8GVenA7vrzlDPikpmKQOeeEfF1vFMguHLNqyoffiEyC0CGOqLiRtaf9KI4I64G/1BioNLea9
M0Xj55sA/yPytF2kCdQmy8bL8pWJomIJpnlmZLni3FFl2hHdri4gmewXNfTEBrAWhEZakNR23g7B
fwFtpZEhUoFVmpUXn8s24xLZcQU4LvllBi3KVmVgyti6XfZOMtDGiehHQCFg+lj2mJreDt0iMrKM
EgRRxto/8aQ2SFbxly6DPJB/wUDRI0LUcWPTjcTU0iN3/Lql+f+OFXSPHg6Kv6gSayB31DiCqgeI
NlIKaxp9mt99iz6Tmm02YV4LOMWaTnH2e6flThBjkxujbglsRafBInyPp2zFqDWTCdiEskQAAx3M
5rSfcIF0H375vWdLpJHQ1/RZBtyE3gZXI1T46OF8x8wHD/5pzxg8duvRseS5Bgz2Geq6BcZOFiP2
5Yw2eJC0YtVuH1DsDvx0GC0Zu6KQhs92bo8tBX0TDiOcThUnuTN7HfUSMf+oYApwUfco6Cxu/6dE
TLm+ai7LwsI+iVtuTMBEadaLDJQXToKh3+TbVaNj0oCE+yvisEWPDaWkrJTaQPVneqx87shchqQw
fQ9j1b0NxQNtqh2Rii+/i3WZJnmkg0VfJavVwPFSJnB3z5mYyOHFvyyxssSltDnq3Z8j7SHxRlug
1+n7Avl2HEva7wK0hIN8lsLWKXFNifWxJIpd9DCKVjfK/Ns1wRrQWgIvDBM7nn8N5sL16xW8klpu
qQNBqSAjpBwIwHFQp23MrOJgiaUP5uttp97QPqcVrVnss77nPMsdUcgpYqX8OpUPfZs4PJewx4wH
2D3g3JQ0uuZ87cIQamMl8H4qhweqBfeVPS862/FBGGHFzqf6cd/ZMF5rDtHrRDwVCKzu9/AodvEF
OWAFWz5uUk8ekADRNLKdkuEuknZmKDbPcBMK2wI28AwnZZV2xlUbVVRscUbzSCYEyb7AjBWh66kG
WKxyhwu2/8usc8MUfSmxLaAQn96Iw1oezf7vQJXHwGP9jgk852xvh01oDF6BFJmHSVs4GfqX30x1
j0QdBUMW3dkFEtcc9Dubp8OQTHooRegmuwrbg3pcwItErkotKimnae8OBf+l5itfjpoml917q0bb
x3sU4MfBsPbF+XcA1QPgIp53SqtDCVJSqSs02lEplYPXp2jQneyzv2NgA7hWhAb+JCtN7o62UC+A
6ZdWHWhXIMNwuC7UA+ECe1Ri+NFIQFi8WJIZx4rGh8oyUD2rnHR01vl0lMU37Y6wgz1w8j91V6F8
0XfhJRxtRcIi8wguokWB97Gai5W8CwWgvTmH5NnKDq0IKmcvBYFRkTpdRo0rJuJA3gwfrQ5I26JQ
R3BD1ADKUGO0XrQULDi5QCcWHuJXStLH7Svh0GuJ2X+0D9f39AS1vO296dXx9ajSb5MZihzRRCMp
9ZcBN/o0TLDMJjTMYGhP7JMkQVR/DmsSL7tBHNQY1AQbzM9iwbNPoSTqbscKBT1a2RnOOVzldlaS
DWZiyTS5tp44fUmiex/iDUsXdj9KiBtjuqUS6Rqfieiok1y2TOWgLsxk0YKt1QF5A0CHQX/oIFsX
JJlN4in05Y5ziephOGoL+n8IxgvclK+8ufW55jjP/pFGqVVH0k+eP7DtFTm+pS6ynf5df9rjxHg1
9pxLp8RkrXNFrd7N5ELCwwJ8GsM/ASVS12l3s7v0dihTTmp5RCQBZzv11kdHgD/fE3VkpsPs2Mrd
pz0h+aOvO+/2xc7hzQtMRypCrkdiFUD8uuKxT71DDZIebCEvCPiXmHkUdgsxNRkc7pJd+rCgtY+d
pVf0kWsMyQyo/hUCdi2s/DeQkiQRzZtvFWvLPScOezYHMjXSmRCkleifxvgf2sR32FKfKB2WB/P6
QpHMmCrgZj+k6uW+jbYMw5a81Ce+8HeMhPx8y1g1tSRidAmu4qxB36dKaWe06aSomCqFjUEsBKSv
H89QOEzqB5RkApEVoBE0G/JBVJveHj9FLv1gLNOoH1cfMA6YQtXaCSmcG9gxIZQ1oBkvLpKiywoY
xyLgHMxBIZcwXvBHQ/TmWiGiyP3jxwGk7Zk+Ha/H56MWTi0tua+qi/kRArP4HkYojXShD8T6/C0g
buChOEQz5CUIevlNsVZy3S7n5JIMPmcTAKFvZ05qldciS0DGKGOKWz2jEE1/hwAFrSe7eol7vAj/
u8n8pBohf2m7TI4UduXK8D8Q8VIEm8fxSZrC+VVrrNgq6zKRpndr6VNpoYDFEJBn4yYig8KYl3YN
VIAFvbl2/a0Yl54iyYAdele6nKhaRI3h2gT3SlQ1l5+0Vi6bD1HpqDziBq5m9SUh9kbPl+OYZo3o
k+Unq0Ai2JVowr1RXA73hCmrKdsl2xSGvlUt8k5EZu10c8ZllLt+r8fnxckdqOoPC+jhlGlxRayM
BuzpfK5dkX6DoBGS0vQlu0L3MIWZP15bYnTcDjxYo3zJGsg7Yobqo9XWjMsTdXoVaVlA9tR5dmCK
XFzdVdmVc+s6gK/A+I64SWTyF8KZwvUuxlhVRwH3mWC2l/VeEXsHEe9C3+iUmcvAELcn+lWtL/st
E1AsC9zjIHj0x4g6NW/ou+wwO1C+FgGObo3ud9pgJdbGDCDtf8LsYdGQcKAoT/he2qDzWKCTY6hq
mXterDXWxJTip70U4zcMMeCKw326cCJ8FWUzKxqoINkyCauJeUa40n0mLwmmLSR2HR4E6cxA8UYn
BOqxKELAohMho+QY/ZJCyHtBp2ijVcX6b+gmPx165mI8QptKqh5WuyJfeg/HEyJgdVBUv5U7OUoc
TecOswSocCGRYiQtYpWU/Nx7e8T35a317nXpiKHGwY/b4RshyEJYMjW+X0mM6eKi8B+NUSESYtUh
Iyzb6VMJ9FzWdoTbSuAxh8FnX9vmpJMJJVefs/rpLb31A9jVWfFubtQ5iKEHEAljGC9zZltM3GUx
Fc/RA+7MjmCnb9O40wfJx+z/Ri3Np00Grw23DAyKW0v+ZhSAPJjRWlfzlXKoNo3IsE/P3RIOLueD
T6EYiSTDnY791EOxZ8/+eP8VtF+e+aRXJmyT9u+sYD7v4cOypFgsariaP2A9Zkvqar83TMAyk396
XvUdU6X+9H+XH9rVS8fxLAZTUDKJHCjhWOU+abiEnPornBoPcAbk0tMlEoSHvDefDiwG9XJ2hXNX
YOzMjMbm04qpyGjP7PBa5tDu6sPCh/A4aPAdoxBpapQ+Gab+BtWqSi9P5fHe5BevMFXu+ShgRU+v
thpUefACPfgTgjtUc2WmvyjTo8EMszWenOmhlXdnRZexIbHwD3vm9x6GaVsrOHK3c0FAbdRgMcTU
lWG81mOSA/n/HE2TsvNT50YINC1Ro2dMZNpOXewitaQX0ul5VAeGanL/oJCInT3yP1vieZytmZSc
xtkbx1T3H+Xty7Jj66ozy8Rl2c7Q0DDBrvTqPvG3UfYvHiz5I5h9RrTEgvy+shJ3hk/Dve7KD4v3
kLF57ZIhRcx1xirouGR/JvICxDdzV2+Ej0jsB3TlkHajxoDnuG232vy+PvM5ampCYE2fX5MwESjD
ete34urqjMl1qvvj3vVxK+oJpnZiPfZKlLuSm3y/YgnFcxb1o0OuaoMwdmDrtR/r1m1Ueb39nuWK
r5E4Bg0Gr0udraTdhl30Qpxe3Nn1ion5jgtMDi31pHzZ3mFRVgLZgvnBoaDxS0yt7EgZb+8hv/l4
WJZhcCS/IbiftIX0zPy4Fl+aox5k8EygFdPHgVff3Ls2YhL3ZTkBCvf4SYmIGkGbg+DIj7icCb/x
E48dizDFFSNtqY8YC/V9Hp2mqL7B+/rLdnrUeEPhqQjwOYeFgKWtYZKNKZ/6YIjEHzSZypY/8S4P
gg65t4ipOtc3X5uj/UAHNVzEt1T1UHqj0sbEpk7C8riuTLiGdbSt2RTkCdLFtUOdIeBYSjjTizlr
9Yy7YNX/BoxlJMJdTO0WCx8/TgGRiRS2229qox01op55pAltAIDs3+zuh23UDMGVlQUyVpVfEh6m
PNA2XTmAvsHl+FWLrE7fVzV96madGcvXkEuTU62CvgBS9Ip8PUwozSUxFrU2KJFtAH15hL/Vq4Ys
BJb2+TmOmiDAgPSE671SvIvwhEQkiP38+5UG0dT7+tEYR8PVTQCn7bklDqkgqKDCYpVkJeMpLFvI
l5JGGUXcjVoHrkOqYp2C7QWMGV2ZLfBiOHYsJgBcWIbqjRFAFmtzyYSURitTQX1sOl14VUeFSz4A
GyqJzk0PHbG9oXteRw452EO2lugR/oQN6uZXi4GdSLxfrKrMNjUdSgeevukOpInor7/A3Mh0fYoL
83DBl+LkB/cxolSVpDxuu3Wumu4JMsF4wAZeli+0Y88Z0+pXXmGHY/7XS0yewhYdE4rQnZChEe/M
JhcpmqFlK0bH6ehjtGUbpS1ENcxBVpDzrEXEXpcg07Pz5Tcbt4r14see49b2C76peeyreYzuk3IO
Bn/5k20WkGOhSFllQVG8BdElsnsG0//9qu7pp6Ll1Sc7RQN9ScQxok2dQBhbMlG0wsNwldPfRbwY
hnxoZfTxUmGH53py+4KimcxqqfBPj8wElYoVKovgGcQj3ptoa/p2Nr9uXuutSvxlev+0AAh5sMGz
ZSf3pj5WYKVZBBBbYNAuslKRHR+HPXDgzZYAnXFUike40dr2po/MfEWTqwIIGwB0Z7yCj78bi+cJ
16nWwsCrQPinzwE8ZZlpZ+AI+hky1jZCkwap0uOlU30TP6N2Bkchok/R+BF7dmyhsxdFZwq7994y
2cFu3LYoJ2vgJBGHcdp1F22bssAFCIOYo1exKHvLPQalXr4brDj6nOvlF34R3UHhK+DVBMNjHt7l
BS+cwIAOmr3w5OvhW54hEPgDv3prD8eIZ89VZICQUmW+hmF7imzq+65uC4F7L8g2lbWNtUMZRyKJ
CUxDYQ3Ie6k61ciqMut4botKBxQEQInCD6JxwQAy9vVlpcnQY73K0YLMv2iiri0mq31YETyQqYeT
M5mqLrSg+kZ8SHBZxDlP5cKEUWQrn+UwVEYHD/hzqs6KkRL/sI1x0qCsdqQExWfRs5o92j8GsCR4
EIau7pLNcB88V1uzpZMBjza11TUUOALEV83Sars1Wevqo0fPE2rgcZ3XFR1cyl+p44+epmP5DrYP
B86reeoW2Q89J4RlYqW1JmCkvPQmY09+AeotdUR0DsD4IPXxRNr8DjlZNaPNaISMNWkFzK5KVIGM
eQee8dOziyVIt5OLe4NKZWCb+wUmHKRyYCrd0v7S6pi9dE16czMu6Ge/yVgPbby4SKT/++0PU8js
mniaT3pNeWyJEilAbNgSGR3gXwZfpamEMxJ9o11dHiRg2PeM7n1nKg2llYCMwmnJJupGYZe7V6KQ
JLK6Kb5rz9MjVssHwebH9wdkR3wOPKKA8PIVMpHr2K7CoF+EmjiVdLv/VBxK8OTcp6MVmgOgNGtj
+kwdEo2Z6e/jH9jpgJUHkKxPFdeHbTlfLyi9fEK+Cqc1PI6PXkAQDGmZ8Rn5OGx+KDeFznmAsfrv
nCOJs8K9EvmNppG43YsMFCzu/Kn6Pj7709t8kCqjxvKR33JpoxgtzZ3Lkb0fQnhH8ovXfUuFCJ3M
lbz9ogbpHJ5tRdIz0KcTJ/NLBcVZ8OrM4JqNde/eh79dyf29ALcML+Vn3T8T8LIM4YZMKcjOLiOZ
hjisB4zq+n+Lz+C037rTjWCBcJiwjQZb71Zae8HN2B0xP8u6L7zo8hmZksvtuFvXq3PmKLFt9NE4
cIs7ZOJN1tnAPPo2zeDZy5LQIWi2l8N9ST11lpQoBdoBeB/syiEouItNu6NyObTSEU9hMnaXQLe1
CgPV5aaYHGKhZWpzfpFg1fxU7XcDYsV5L3M56HJbL7K27NFT49YPplpEHfAnXo0vKUtz4zGHa+IP
XlVk2a+IjssoDyTjfGpIXx5Sm6uSZ3o10eVJLnVMmhnRcgZGdYNKcQzaWuET9aP/sXhc9N6908eh
fyFi0yp+aZaeAYUP0CKS76tID7Usfw9/qhH+WQx1cGoG27MsytrNc3Ou4CxDOy8S5gg72rw3tKjm
e9IOHKOixdotkl8z78rquXvG4Yg1RXPIjA5l3sIxVUleAC4zVrfQu0xNHFyU+uv0XRVcPtrPN2Sf
pbaPjx6iL79Q3nEHkIworpqUDt88px9PN4tQw4GiNoaK/mMG5TMmeHfcS4M455YhHlfnvboOQ4Nf
RVUoXzdJNH0rYHFX9BiiCd/77JmXTx66vda4HockRqJUHOHFXx3QQlHkBMzd9lWxsTaKntUIosEH
7qZwH6gNYPOpBNZrXOCrH1vSlweKLSs4CUCfEhCLY9qqBg2ZejL0u4GnA7QDU3M11yPUR234KSP4
pjJc0LCifp51A9ZpsWlD1NCTR+4yXMP4yMvVB1oq7rzFrKKNJxrToxG13OyJsW/4fRZULzNiDWm3
8JNbjkeD1O0WlWx4xZYSv3Yu7WAVlScxsiEZiPyXWAtF+9opy8uOrR06klTow731j5dEzfO76Rq5
LBludAVPpDEhXsE9EEW6u7rtZdE/4YcwuTAArSYLyD9YBMiTRew1aC49BnIHRPahmJxAaI3R939Y
x4ufj8fHdXb4OUdo7QwTg5l/cB9z+MRZdFyllkuocLydUB8UH13g6/xQJ6IqsJX9oR3hEyaOEnck
rhRoVvLwgvu2m/ef6d8In1XwTLjZj7Tap36HQsOEUhirY8zZqKbfiJZ0ksqEvK7AALSghF2ypyY3
wNU0rFWBXm5iCZRD7lPMS2LuGXy9RV2SUeCv9lQNiKG0p8+9RNRAKrXQolQCYpElLb8lE2XH2+9n
JPBsSBX5EjhoatiL3mjG5h0uBSj5qUjW03+yKIFhl/2gCjZkrgSqGtnG/SRj8KACsK9MaoPRQt0j
bdvcbpm5lIso4qce6St4MMjp78OYW7kC2xBXzYsS/jP4hUzdYD4maHu+8NIBmIhBIVkiu3ybhbi4
kB2PBqwU83gKSN+SszTIXGk8BfsEtlQ8n+b+8hOkjRq5dEvmAQ4z6nNoTWSw5aTcbQnpkuT952Uc
II/98KriP+7krxJkBdIlFNPR6QMFnPPUb5MagReSXPjhgx2cdCVF0/8q51OyfY+7LLE5bVuyYoGK
gRNkEKeaohboZI++sRdcT1/G46/c76I7vM3e4LhAzkdVvuyF8VLMONivM9BxeoHwWM5PIG30XKP4
+ImTWS9tXY+3CFtAf6adI8gfRKgB9ViagocQyHkub7FYYkkirXdRwyRUwRPnVAksUI9b66HuZMF0
uHx9sXucAeCP7u3gN823KWNaVAh+dk0zl4JZYdtQK8U8/b0aSCYDbRwuEJ64yGT+s8Ph9oQD1XtP
1a5jpID536Ub/8jC5+HHwUZ8Xa11V90wGxnfOtKWAi9wfMUjfEMVCLWOR5JGHg7kpgraDNxZOEYN
MTqirwXlo2v2VzqASmglsI/bk2G9akl1RZwGaecqYmjEyGPIZB1yi5TV4xJa5De46kvnTr943eL/
TTVci8d4lsJAre6N+Os0NyDFJ5r7SxX71A3vIZcEBN+Rp/jza6VTNALV0m/Dhd8Z4snYAwWFY/Wd
dVgwHSVtXYGoo98gHFW0RKvf6yVNfsDOddLRpX9xiOJfGR7JVSe0Gti+jkj3ERhpBLCpWsTL/Ewt
RDyJfpY3eomCqvmtw34NoP8Hhd+4CggK6N8baWOIR8Yv83nQSSznT+aura35ycDiaAuYUDOKCzNI
qi60l+h7H37gwOB16XSUT7kMxGD7w2gdd7HhUAb76M3eLuQ/ybkJ1OOcW2ivx0bZhPo5t/9zGi/z
chyYs/YzQ9twukfIupxt8+m5+IdDltm1x2c9ZmkZANq1Y/IUdxqywPUPcMJIUNcc55Cle0AFAQqH
USeniXDfU36qEdd8/owb0idS9FBR0ume8QkkC2RGENvFYCF4gEg5xfP4AGcDXbQgZ4VstST7sz80
/BuWcAAccg1byEJgR7Z8ZEJbWNMbEmuxFeWa7TU88gCHhIpFPPm0FlYyIYJ/JVwJdqZm7Z5tOyKT
RpadW6K2oBBsL1LZ8jGaKbeOCUgGyutgeMmht7NdesXbvM0Q1d9PYdsDRl5s1UYht0zhVhTuI1VD
c3YV4k6jWJUHP6Tu1m27EoWHMHYFZUN7/9qaYunfXTJGyKxtKXOuAlsaySVGzHBZdsyT8sUatheo
cPS6rLsmIcLmtPpfbQlv5OgiyW2GT6mcYJeFon/l6h3fAo1WyU95ItZwWUd/o6bw1LqNt32LHGl+
29HOvEjiWQlGiafTyInCPoqxs2BPpW+eQ0X9oDcJ6Tfyjdz0J6p9wq+W70YA1OJgw/KydNWoFI3f
udeXifjY4HCuKKeDqg7cQL7BC57b44TikEvgQcZ7DolZDR2buCsyQE3GWtV/2UCR4555Yi+2AKzn
S1TQAosWaxQ8Tzsy7xQJ2DuFWFTgKIgKA/83Z04LxXWV6JgY+KuqcnbsW5qD2rg2T1G6iKAM6/PV
694ndwbfU5pzW8gSS08GjkzQGUEUXRdXuidV9au7d2SLI6OG3SBQLTfAnRcZ1Ubj70SGXnCLjd8F
TN+EZCt5WO0XbMlwvsID0gPla808Z3qQxwoRhLCfacE36BgZC9npJxzcL6JZ7uBaB/e9sh5k+jVJ
zl3AxI9ppI1Hc8GyCNBSfDnjKdc77Xr8SsiuIxn94uLjVXwKDiaCOms3aSs9qq0h4Ec/SjjjPuEs
zH/MmTXSGhmx20mGv3fiVzkEkHGW5kjU58qVt73eRe3dE54Rq+0w9IGCKylKdCPYJUS6hlFGIeCY
G2IjiTGyZUzb++HKzR/k9eGA+BtL8aAXTB4G0s0ipBQrn52Gx7ozQMsZH5e82j5Rk1HRcddEVaxb
YIS1L3R0bWQdPAjQxHjkEHF//m74LEq+vV0yN1s4dbWA/Mis6U6OhzkjCXOmV5lOW982+JZ4KdlV
k8fL2PGes7u4SJCGdga4NqUOJnur/W38tR93F5GVHTBLgZIUm5OPJgMZdG7gd3z9eNfH6x+Ki5ix
RT9GbXWbuBcitdhu+nMcRSuXUjtRoYJKqGocuPho12/lytRBGvrdOYsxq+VTEZwCr0J91Rj5ye6K
l0IpLIFVUxhRQ7udiDwqUQOgL1dHmbaomWELzSJAw1k7xcGmVIxdOXSqY8Ibqfk1CfJccgqjnYL5
luPR7mNAkaFw8nEx4pocaEUYXa0THRC0WscbPGG82JE/fcSc1HMmROuKzmDdLKma7xT8nK6Duos0
pH7PAQAWsAz/0BHfvp61KNT1/WLLesnsJif0VSffgdBIvAOSUlsqstvt2stgGB3vgEN0rfWxUzwG
ujDe4lF8c4ZUySphOw3t5+O2vPOajbz2vKRo7aCYYf1dxxT5Eu0LFgM+xvV/weNnK54+oNiESsvY
T80yNIcL2q0NJ+EQ+wh0JZTlsWoxZlojoxP91XPMXzNz3NXxW73a7JJQCc0aGzz2LxXurG9BxmrK
HhNRlq874CMr0cA46P/8flI4+uFkA/2NPti/NKEkZAZqftlWjfbIKCQ+RetD2qMvYqBda3nuwwfD
/29nmZVPNoGtIiONS4C0BtW3J0061C4v8hX0n506nUzQ1Tol4GyH+qfnKtKnvijrQ4dCWVsYgkaD
XU/HCgbw02o/c4AWpa0MPLwY7+LSfstX5Fpg5d39fWmB1k17WlpWXqQaxpybOIjTIr2CeNboq5TN
uaK0wgmQjjmMr6AbF0yczZ93BSreqyuKgMQFGM/ZWbRjY5ox29xI2GSlaSANvbt2RJyNvGALxp7B
C6zlb4jRtKukniPEKvA2AFWQ+vclvA9iY5/BK3G56ESrNExgnazMyw5OBtZyXOSqDGES4UVCU6lq
aE3IMNhfdBT/ZQW6rXMmTJaScTUElWabdUBegOUz2LKPJATQkMJBizLpn8iHdU7Ifu6pioKwDTnj
0JM7zjYiaJxSXLDcDceLbTgG2UlXW5ZFNIlPVWqyMtWAmEeypw0zH4SgjSldMF661j64vouHon27
frn/8EKKSW0uFPJGwhkmh15Ey/ahnRxNjWxkUvmbBldDVGLJjRhJQM/5+5NWxsKhmzBTYmqvu4JT
tMyifX6hFDK3ORKpIXpRIAGgL9WRVUPQXpQPyYJ67ZpioGuu1R5xQW9l97bLEd8cHO0reTrDb8Rw
EcVK9lWiPSGODlOvhT/aTAlKNWBn4GG7hRxwfKodmviTOozNmqPoHrBqMWKtDF7KInH8xjJW86mQ
oFNJMAqyWgUgyeJLfec0P9NxAYDvgbQTSvkFEb1VTxKXi78X7HAbs5Y10GsUkSvF6HG1SqGy136P
eQG2CrVGGnemtmqx/h0zEJS0z9Z+zddPZd5FiKSGO+/nFZQXDRhbLbgLAO5j2oVqF6vZNFtJAVv+
F0EhQICFLymkpTiqHk+BkTXFNg628AX8n4ah5hyjS29uMdXJY4ZJB5+FVVsw1gtFuL1hCSY7Dksy
0Bq5grJFlKSpH9vq76QxDnfwLU5R30G4HE+shrMXXnfzMKaLC9EM6VAOdgvKenbLJ0HUv1cTzNy/
oqRlZXImgOo4nlZ09OUqyEBOgg45UWgjOxgqQdTYzzhPirrM+PmpdTkQ82dgwtesJs8iGosinOPl
Z3mP5nFKps4uSxjegzaTyOKK6fu5TN+euz5er4N38nX1k0nNUngF0i1Wv4IfXZueqc6gLXg8fYtJ
nweVqTdTkX+4QHV1jXCsq5/R1B6uXG0Ow85AdlndoZ3n3xZSXpCOMrwLIM06cVQoPVhU0rU/9uSP
bdVJZBfnmLB4L+ccDwwaeS/nMaZ5jhmnMFPxs3wF2QfQPwoC63NvsC01LzbSLGx7xQ3wXuY6MOE8
CfMJo5jB65H8ARwG6f7XbWE5M1C/ntyQ0wE94ESoV5bkpff1ZOs8V/ckS5NuSds3SqNLvZd9zUT4
gCTgha5WPm/l2EhdbnMU4PFWLhVaX2f5Xc1hjq5e+dArHs+JW2azLNZKCgINcD6D/FvM6LkaN1h9
05MO+zFqInWkaWzVpA0KV415aQPbwdujW6pVaRP4bV2RN35DirxFdh9bs6WGhaB0PlYrlMXsTyp4
WnGarXweLYySbJUke/3dXy4EhmQQcqnzdP3/lU1p5BCirk/m8t3RJjjaMvxxgWaDh1WpP5ZjCFGY
bKqHWs5+SImIElGPzJl1QMEcCss2ziPUrMzTJC3zm3xelZevZPaXCO5mf2dN3luGRgXR4vy3tHFD
HXOs7aqGXDnSDyu/R7KjxWl0onqjhn0ESSHKPPhPOoz6i1aQcLRt0m1vnDJhvmeIhcTmHQTik+YY
jo4jFX3eQQWMMdQeKF/2fkgmpfCwnsUu/CXAtqCchn8sD7WwvxrPRUD2YxbQeyuDIsWwMpSjPGra
ep9rsi0Cma5rxOwS4e8T6P897mO09Ojv3BBG8VV+Tht6Y2TIP/QX3dfbch2XrxevH1B+DJym+TDf
3gp6QtbqCa2ZH1nFvDLj9L8Tzb2iLt8w1VRz8qR/EjHPAUc85NhQdcax8RjYzrNB0UKhCNgT+hot
oZzkpoX+FCTOUfUjsbbJzZWhPt1Onqodl8DL1syy3FQRVip2DQMhBxY0nSkDJc7LQHxE+ZMu52PO
CvsG5EHgOD3UYz86/EqRs9Hw9iklGhDXASHBY3fBTQLrKEk0ElvUNMGvuksH3Uft6NlSo8aFRmMd
iYOZKH4XgtcwZ+MGALrHQOxHqlX6Pjswl1nXuGh1UGFbKAU52B3QvuJuB/Tm1KHmfhva8cwatVvp
7VkuzE8CuP7htYxadmOpwgVjSKB+m7Suo5wUzjYbiKK7MrGliAVlxddpBJJmaDfiMK/GbhM535te
jpo8sA5bpsEIrNsUkRw7VJa/kdOPx8xGoOFDStum9bqxnr3RekKlhvMAGNPpBBIL6odoB4UPKTdr
dWphRZjpqfCnKKTOuZ/Lf1jLCICeWmecmuNLQuKYTN+0a0imnLKX8JbeOUHV/c8JpohXS27XSW8H
0zeGZZcZ4jx4+Bcdfg6mLEp+WiINLp+hJcieq6f/RKxOp+MUAL2JYxE+DwODTSYZcgXx11QJvUf2
kIbDfUznyJI0NybGISgLoLGpKK9/aRvsnZMpJQANJGxiU1AN/v9PeEC5dAJr9IaRDrL61Wf/M4hL
Yoy3GXLQJFjYjlW6bogfgOniQmTpk9ook57k382DBr9ZEMOk/wl5S7yH6AYtlvXYG7fCIUZFVvPN
hbiKe7ABpDb5QaEw4ZzM3hJkwLZJXlOWmgzjai2OVeyQoietq8Z02fNtmuYRB9yJ6PnaaSNxd8xx
JfY7hA3tErvjpSRhz6Vxh9QNBtzkXboN/1+rhv1ypHhBM/7gCb/3dzDVaZZD8MDzjX6rYuD2x8DB
TAqHW86Y0Tdy4E3vfXopNxVv8mQakxxjHhDonhhlyZqTWqBFt2+h5MKPbhyS5aNs5sWA54Z4qw5b
EQcSReH03feacURyyUaRfEcpbc/PlyhEjuenwa3dJZ5uM+D1/dDD2jMshuFCrIcuWwOIw8ANbCfd
8YEJ8oOOS5uBonDDhFtvi6lgCDCYPPASTt3BvjCnLF9rQ6gTBN9/l9fVQAph5Xtd2SZb9ybkOSoI
ptifzfN6rKj3efkT1qCrNBehNTWlmPj4DjCxQjycX+JDubYEiPRW5YmbjZ0kwOYMvf91VqatiswZ
8olvelbfadlFmRVpsOrh/Bv3SWXT8ruuwJwFgGEYvuPFcQEobJhmCSo8E53hThLykzf8/pMip//G
lLlB8cTmtmDGv8j/XPtkzP8TogykMcuFNWivTreEvsdVS80dfjy8/w6d+zn7gxutGCgv+63UbG3h
mBqnQvtKEE4m4t+FCcL/rt4j/MmqLK+QgsG9C/CTNx+KtqY8SB/Pz00LoA58ZOKtwn8DjYZGyG/H
dV3F5gL5+K9FJYfq0rkmEa7dmxDiWUwMOlWkdvfmo4zxIJKkYQBgUdWtcaFsS/ePndwCJfFANiBU
tSAex9UVSv1eGVB9kkDhKhXC0eypSMI5TwAJ46hBqGAc2VVPGO3Q9hM7dlCavcmPzkzgIEWRwYaS
QOV38J3xPholibsHC8UlryL4ytKsuNn17lztwzmjY52fCa3mLqogKZ8997KsVN2bas0DbbsQsMGz
3h0Wd37WPjFbyBSC37FtDQUnlYdyKFXWtR2//4SKuVG1CbNRLdrWr76OflRWQxyK6cz+JDfMjyAW
1M0ZLEvZg1CNuvHjPVCgQJqtlv1Tj779vN07cg/HprF60TJodCa1pax83Py777SaDjMPci/+wuXn
mSkeqwBfHBTfr+54xWK/f56VVyMebIZx+nbmoGd1pfI+q3nXvqd6oHKWp0Xf46Rt0n1aclJ6LgJA
Ws4yX4PnPkPi0RvYDJTCsAI035vhQ/aJ1QPSRzEWfgyETwrVUkNb8VHdkpmYf084e0tJ5Ptw5/CR
jhaCoGHVBd2F7tvaWCejOBIl4Gabe45F095pW9Ggo/I1Sm/zj9HNe7VKjq+tOTQEhRyqyUChAEr2
d8wCiVU33+jdHI1Psa0pnpOT0r+B3PflPs57kZMIz9+AJjDZO8VrnrAkFQpr6vX1qwsWxg8pNunF
Q4T3sPksJ8KWNtC8RzpxYdlbu/gopbmb7Pxo0jsw+vklRWsz3MqUmTRkL6BfMBW5LX79uFu038Lr
I+DaD/At6XrwWJslheP4JnUl36v4dZPC1lz8L+MCBY4DeAZwrdv40yWSj3vDjr6dNDFhMn0iWenM
zeVDeSoRfLo8JW7pCRu2vj48tp9hJNGqXj99VYVoR/TK/WAl/GD0Ub46aIsiwJ2adGBjnoe6RDSI
w2BWC96b/M4SPMGOxZ0uKvEN3o8I0LuuUfm7m2ms+ZvPo+sUhK8NqwqyfyDikezYvVV14apz6hDL
2qnPTYkAVbi2hdguUqayEqCOku3t8l89kyAJTMmA24OlsvUySrL63SyivXXSU2g8pAny9Vm+PnB6
olWgWdG7GhYgm3HiVnphRwpd9Q3QZdelmmMtakQN7Efgb+ZdEviThTqhZCbfca21RsLJsqxv0l4P
b8ln+mbkxVGnCE+NloeTNn2OuAOk2YGH8DP+C0DhRKmnt3QNO0kaP2qoccspGUFiMSCUa+EGzlaq
LBAsJfQVu8JTnPSbSznoeVZ2NK4M0lsaVc9hvWqgMQQeRnV8W+SOQ5eEWFcBEcch5W4s2nBNpJ7g
9yaw8nQGNRcd0Jq6l3+I0TVcffQ8vMuhdOYq7kHr3OTJKDjiC1sDIDFwqZJcygD4JDWBW9tyi4K3
enceX8DtcC702WUOfEd9zmM4VHXnk12AI62E26VagHcHZQmYr8tsFSzmzO0s3pANNXhihkTV8aiu
haOBw7wMRuDRJbzQ5Y5dsBNp2rp3YZ7QdNK4FVwy50JebpFQ3IgA+jCQJJxo2279Q8itjBsksFa0
7f5X1vfCdOLPWEnw6WeD5JesKvxoFmbLFbzTLEsyYiR17mARIEDn17eub6ujefiLcAPnlzLAB9cP
MfDGyKEYDrE/gPQA8RlTpuyXOYHBBg7Z9n7FiA3gysqapbvVgIhs7NO+AGu7RIsWgFm1Ipgcv0K8
oiv1Wcg2K1Ok9LY7CU04MwsaYObZz3HsYd7B4qNOs75AVNeFasIIjl9e5lthv5bYgivd+hRUSvg+
1nY4r8VZIuuwJiO5j9v1e7YarvcjC5KsAGXMXsJEerX2/1pNsIZ55+aDc52vnSCRVylFnAwws9JH
oruyBmuKTnWPIlTWb41U47sodaEVruSHr3AXaKyuVDLzYQpvrEVoEhQP5GkpoFAtddLt3WTSiIxs
kuuDCGkv9IZh3E0c+Ek3iBy+oSrJY88NEWi+OF4GZ8svez/3LTO4MfyB4xEhAN+YUky3lI9uonjF
U+lSY+JuOQ84/j2WDMjgv8J+4zVcvnplEl16vj5YSlyzBIe8pdb2FY0IaQRvah3IgZo5URQHNPz1
0BwteRdQvF4uNeS87TqIULYPGEYZQHuM5CedJW/LEO/Ljn1Jy4vy31DlKQN/gLaca/syeb4xgj5v
Pgejaem+LR53fWzmsj28XngIshoBC5q0OgUJ3+H/vEAZHcHr3gtn9Aif3tSq3vNeGEozAqlLR+8i
cNDDnuormr03VouvRv/vRhKJ96EGGNMBxcjeYoxhM6fLqnpO+E30sqFawLa9JJdLmXAqIE364mDQ
lchvJ1I9LBDdkBvXXUBXjbaYdzSby/1FRAzxMzbD8THO9E7ly5BjVR1AblGZMN0d5Nn0qf4FSOyr
xuKxSxEO9J58YEphcMOv7Yvo0UENx3OWHYUQmJSt2ZjlLMziqJKicCIYEYWwxgqKOaYvjodf91Oe
WrQxPqaNKdsNuf1t+6y9hMXNZPqUn2EkbrFTyxEySzyGCQ1C8FTZEXVD7VtMC7dtgbj93Mr/ZvTR
DASMQtB6A9CF4FxHPlKASY/4FAn/2+OWuOkHgfFkN5yIjdxQypC90fEOxcux7pRR/0qjkjqs+vxi
6vn8pIgMuzbhG2uTNXx3PaeKG9t0mX3UVibOSkZEtH39U/okeXCqyNH2UV0K0QW4GGenhrpg51Qn
JmfkhWy4oMtaGTpRyyD4dDINeDdTAKrwPAMphAIKwO/TxIvz1Wlra4fqiQSRaCd0mdbhwvbP/SGf
mu11t4gS0mVKB1fCsGHP9/1F+73QqU9+HF5x6PI3nH5xKHecfcNHj1z1js86ipZ3z7vYjZJwGTsT
ovD8flh+vjspkVkvegaiCZGNhz9/1ho9q+eeM4BfwEHHckV5hW4+YD4SW8LNGuqxFAVN3tThd633
4XJ3tAfia3p7BbBr458T8w6dmUoQXD7aMBLGoGJAg5QyEdHO0eMkwWiHTKXtlCLheDIDuf/1L0/y
itk/pPRSF7OK7SPZY2Zs+SOEcAJ84k32L15nbZSU+kBGpQybCbyPwWjCxu2n4nt3HCzUiXlIlwdY
ADE9jSNzNXSY80NCY+tQYfhHTM1X5Ye9o72kRA6I1/fi+LZqo69TEg2YAWz4zA2Sj/o/SgzL6zfz
BXvzRoLK+bA4AfpX3OynUJ8Z66mz4ybFmOkID8pjGHHWoD7Sd59JkMqLwQrfOrVUwUT76yYi74Zk
4jwYtADg2NL8KRl6FAaRB0SEcgRxY4G9fMff0J8POB4PpCdyLWrkZdc4I0fi2MibiiF7WGu0Wuls
XDv4+dhEtvnnWTOW2QPzdqSXisBxTM/mcA6OnzVBAhcYNdH5kemTfb8Nlpu//HtP1tAcpz/N15SD
KFzfwM4jbZXVLaxCflbzn3fJmXPPh0IlqtbJh+Gr8nQzVZdz/jf8fEdr+0dYGlgjHyy/y+fSYX2m
8ACdGSzuIjSD3Z8usrcR6VCTnxuPIX4i4YAdHF0fMM+3bi7k3leHCIZNnaPVADBJH8wqSo9kXY7R
eQAIEFCzOEyF5X8dQvX1hfc1BljE3bpIZoO351wOehJd2Hb2bSdTzro3jBewIGmoCNeh4JuDge3m
PG7MqjnnRFit0XscAn1SS6Nh3NH7/cpItpoctsD+/b7+kxBreTbfOBxrv5+3rAJZP/rBRe1tLty6
g/pOTUAVqsEkKz+en7Dg8pwEJWN6PICpASub4JS+D+1DWSr1g0elBvWkN/Gfm2gwaxjhk8UQWrbb
DZzJmseXsZv1y7FMh/V0FsGNQHXLoXamIIfDh7qRbOxcPxrCTCP6GBYslwGyL4N/d1/eBBhIQJVe
Q9/E8WW6B6/GPrY3f6KgVyR5scg/mEKmKsAOzdKAn3h6Cy89LTvu3jKvts58oHFMKzfEECluDz1V
NwafSM2R8y1v9s3kAQ4s2Ymnf7/hXaZTLYHT9EwKxoaBR1wkmDc37wKXqXTPSxphXbRwDVEaDwQ6
S9uZUfMQh01Q6EDUOWS39SqAHYZxX92np85IYcnVJSb38xZLCUzTkBLgn0aQFg3EGBrUphqgkXhG
WS4MgkE9cVuKcQHW1B5evWKSqSkp8GY68WEFBfplDiIhKc5uU1SYYST0WtwKCcgBHW+R1HIlOOjD
h1dK7B/3WYgOH03wShyOksOc3ANSUuJUqFp4Bq9n6a/vqHIqOIKm+Gzmbq+6TMODKoPr9hw/PP7v
XWJQDcWwm1ms7eZ9/R6jw/g45OEahC6ZieX+gsQDu+Z2kKl2GjeTMnEEJlKx/WBNAEbzgcWqRgjD
xrBLXoistb6uP3Hr1xz5AtTA6RezQztKeB/qzvkta//WusNZ0vzMjDs77HDnvULWYaf73Rm9bYjV
ey8nUVT4JMIopk/2AXZVGqNdIFnKrOzUiEeGiWWKwln7yYDMgqj7EgegD4Vu2/sbBEDafuzRDZ4r
HEt4+aRRXGNWa6Z1XyvFxzB34b+VryANJmzuDvvJJuxPxdhIQlPNZo31RxmvcRzTx4AoiFB0W5e9
ZmS9MtPRMl3SDyg1JhogbvdcoT8U9+evMsKiL/hqyxwm/8A5zKCEdM2g9OwGPFlPPlSnKSprQ5k8
1OxBvpw/sQQOYymHFVNAJvmxFlINgPpbqxUnl77c9/OXtHKIjfz0qXWN7sxtcZEfbEUP2ya94vwO
mEHzTz+32w1zDhi6MWBUnYOis+3rxkW7YfT8430l/OEM6rf74Hx9ocXBNcLbZqF4A8re3vM4cIlm
AhIawgU5TUsBSTke2R3Z1JC3MjnDlfoZBmvgZxFnwMFGVuMPbvfnfOGwGwhlKhcTsnbMjNK3uixy
8RbkwhHIKUA5mLPWWtHQE6rR0fntKU/BDojLjtdm+DRGm9/rWlzf6Urb1AcNA//CXWP09Aen3X9B
XHgt+SandGMb7Sbg8ZjzJ4RPbsfRkPyQ5Q08s75UJCBgvR27Nx2eNzV45j46Qcta68OccR/n6ezz
W4UMIZZPDtgp7iVY85YpfdnBknyaMPyT1IRx3dWnVm9w8xZwgjAf8VipXlE46dPgZ6LFeZjzpbA4
OcIWB7FjKiisxkBWFX4cMEAlh8UK2ZL8KBQQpr4AZ9RLbUBqXkywz9yHmiTHVVwgu1TcfRl60O3h
TkLKzIrxYe4C7o0j/xHHCp6r7gkk6rl8Rg2CDq0Vlk42DAT5yh/7vur2kvQpr4dAYRv8mzJFEwqo
Nd5JiAil8iI8MxpkgFjx6I8NYhR/or3ejfEWy8x9nDNr7YWFhGA2ik58TMInf3Zl8FldBXk35+cs
YprK9CgZNLvuT6MKINYn2hpwG8s1inhqrzm3bujxsHXWwShlCsZMviYrjb2uDPv5nSJUPJjgEIqt
lzJ2P90mZ1eb7t4yzfF2a4eq2scJWEDCjWR/OylvB+cAxP2RiuuLKsx8UYNSiulhlpo6zMUqhw1f
t3idDi4+cr1PJXhmruJ3M1iiejEMrFceRA2NuzoL4rQQkKey9NsLLczo/TkDZkiFM8yinFrcQW94
ua0QaSD37dUQDvTxbKmmj7o0DtCoX+ngbbT6VIkmMJLiKOHNo/SXg5jLfG/9UciZnzweAyk4wUs/
7jSO4BQei8wksX/mpvjCfZ9uTqroPsPjgtaY9pLWveXGcLPUntiOTKHJCZleBCCGo3x0ZhYUvMz2
/RiWkbo7YZpyi8xF1Pk1bnG6JYQxnq3IaRX+8uL2mpKTVTckUF0c0bjFa35tigMphidmYQOzgOtX
Ui6oNsjYeAnsdq4dS1fAfTPYiKszUQMSiEf/nM/sdaoiXojud6yg1VwZ8icCxmbQ2xEOnQ3gLWnw
Liyzhvev9w+iYCu78H+HfGpSNWOZdWyqrCZ5Cb8UXKA+3Khpo9EPTwF2Ik9VqJOSBJHaN7pg3Jgp
OL+hubsviI8FhZoILNM/iLN0xpiQQEN8WlUDt9aRUwb1xvrM7ZMVWbEX9/fDyNY3Cq2v9OoXHQ2v
ymbVbpFKbphSy85dznDjMY/eTPKsRD+sbmpPOVLq6gGOMVJKXtdBxOJWI0fiENhCzmUbsUJ7I3K5
Q5PGlOkM0B1TD18e/2Z9nkKYuNh/ulSKjqbwQTdqB6rTdnPWD+wk9sN7JGXyX7MuRhuBidy8iP1q
5wqAV8d6ygeSRTuecauKMT5JAJ1Pkiwy7UdD1xP3ZUMVHrgKy2vqwo91dyRTpXwgqXPisNw0AsGs
ix4MoC0MbN95KqeIvX43YoYxp8PR9jQEkBC4y89uYqyefGsd+adoNpttZFh0PSCM+vpc38cyqnR3
CTpULM8STK9lZ60yzsBNqjKCgI/TQZOIGpZo3O2JL1cJNzF+hiPneajj/qcOUoHtWeHv+GCwc5aE
/gwOB9YskPBFiKJz+n1fR22eNkGL0DJaqlDnK5Ux7uFcnk2GPJSCunGVRn9P171oBIPyu0qzwqEo
8HLjvyhWp/gcecXvXIGTrLNUrS1dicHyFjwIuqS34w0RdO12mDEuQPqXHfSy8u1AT8Fkfz36ByVs
BHuqz86d/zxRzEVifaTbTW3Io6Qt+0D2CNLdiezcfgfJgiGeHlyk92CGRTlmbM00VKvVpXDdE7Pk
jbgCTsK1TId0K6B57eEVPR1HEqQLswKe/Qmq/N4hVi4JIj9w+ISc8YYK21ab1LJuNxe1BTRgKIzH
dDZ/1+ghmw+jADkQIrKCLXdsYpHF375sEWWDD/GKFWIwe9+tL0klk0uEOnFvZPskbLL+8gP0rX+T
CwmawRHnfR1nA8yBuXJ79CPQni1qtV/9cSi4tbIMJRNd2NiBYHl5O49Vqcm95LYVpZj45JGCjA2S
hPjl/9SdT1O+TFgd5YY+zb8gws0FbiCzc687GyXcdoWzR/s2YGBcfDWUzZZUt9xPLOw8Q8y9QYdO
+P6dcWwcs9TkQ4baswe9EfSP7bRGqUaV6W1PRawPo4l22sZeLPjTFOf0XFvANb3teaP67hGdgsRQ
dUk+o5Mw4C8dmqyFZbsmBYz8sZU7JqNhqUcfJ1e4Gp/3NOOIX/GWx8j0zMWHl7zQJOhR5qhK+Pgo
eSqV8wyYHCe4KHMrR/akQQoJS3tR6Qwh4hz+iQGNC5FSpvpKOQfr8XwgFI/d/CFVfu2uL12IOgnj
2V/M6+ahPBZPd7IrQwN2Ujwb1jjQNKz+Dsu0NVJ5U4ewLpRs4QTTpVwC5wybtzJqpZMBY+E7bsVS
PthP/jzW7WMjPc8bxFGOxb0rwlstENrrqjuTlKqUy/hz8hrGBYWT4wBZAHh1vk78wBVxBoAZM99V
MciU+XH/5EN6XZMzDLAj1rlJNdZkUgaHWIefvCMTJd02b2+OMXG4b2xrifKoWLd0dUYQhqTRZucs
Gn0MRk4wRUR/xqWYDLmmo7QIccjJKWp+Vt9bU7jwOPqzeA5x2rC4br/ie2BpQeAByQtmuFnhIaMd
6Zb5iL3/8Fk5L73d3GGaPbQXHK2H94AOVzytCc6/43PLOGr21m/hXwmqyU/UA1Lp/WGsi7EUdrrs
tQYQCWFLNBHdO8p4JzoQExV7iTuWBJbTyIY4mNGk4ZdcAIyMKoJ8L6lYLoAsZGSmTINAtnmwoX95
I2/iwcoebVQCCoqwcYCJiWMg0MW0bgHGOU/CLgA5jBZi2K7H1o1qQ2wq1lkRLkZyYRq37puUzbK/
P9achJ9U5etSa7IQGCeL3P1sayXQPaaA5mHLSt0/yAe7PzucYYkNKduJQB4gg7FZKNLyt2py+K4n
GxbjuiM7DyU4FaTTi1NmHa0zGUPfmfznNADpwzdbv0Uar5ucGz7fjPyGiQE90ck6Zd0+aVnEvWPK
zUvyzQbe1X74/gidXjWU5+OZ6mRf1zP0GgQteSK1Y/z7vXfdPpIga7RUAArme3RSmdBy4tsk5UYR
uWEP2X68mo1//fbVzM3aosYl74mP4Myw0wsxvUpUoDgYzD1/l781BgypFCmL7aMzaGcwaHsZodei
v3bNahcywO8u/yVNcxrdfKMX16ZyrSf5n4XACErNSAHwPYX5PliXvtlLZpyWt0ik6Z8rGsJInwZQ
wIyu5uAvp4pQ3HPLG6iIcsiF1oX3R85Na8iYaKCgy13fUd9JK8iBXRRL8RUyyueKH9hS9NP1SILu
curtb2bUMSics5nKJguKIbRzbag+YnbNkwVoyM17f82oFsEXdxDUCpTXmZUqItat2qQDn3rMQ8EH
KL5feZLdGyYYwNrMM6zLn6i22QN4Kw8eKDvE5hK5IrB63nfYGGZlEoegZol0mLxoePW4o4CA4HKu
mGwMaxGAsO9abJOfMGD3F0JtrAMOYvLjKelB83JuLuusxms9JSBTiTWrDbffztE2RJ0tKUH6X1MP
Z/Xcx7SkfWb/kJOKQWpng0fYO68J9RRnDv5fr58GA6fz2n3KxbdcBEzyddP1gbtuKhl72EGkdWUS
qNwMc5PGFEEuDq39lL0tYhtyHbv19+Rb9bmdSEP3ne0ktF6PLP002KmGGkxPnzkKXMfCrV8hcxBD
Olatf3xmY5YCcTdA0pZcWr2PfCVRTClsAW7uxYqIAlyCMhqIREca/0V8SWVcLPQ1NK6ql/4kp5py
xv99lvWqQHVx1rwpiK1kNMwFMx68SdT2NOOdE+dexR1A1VcUthP5vsP9XZZeuGPAUV8P+Wfp3Ggq
VcnPpY8dgzz4t+HRuwZt2/uGZh+Muz8VO01L7iuFWSd1uTlFvFJrOYpTV96WqBsaXYCvaiJzk4V4
5lZs5fq285qMLYCdv6ns3y8D1PkxUzWGkYJjfxBhjll3qNclOIL80fpnH+RtyBO9OfyaDlzYM/Cu
Qyq7lhAAqURhBZMs1du3a+Dmdb9B0F0+BE+cF6Pw01DefeIuj/YfkTySZQsCSakr2ln/WIhaeD+T
Ku09D/58G1/y0g83YVLFTEgHaMroXs6AsUS4mGu81mIQodFhdu2iMQSO70U+PJezcORkvSuwsUG3
iKet68d9PXMSI3PrhNAhIKL1dfUDYVOqX+qP/N0es+KQ2xcHZMJAjWBTTmHeQszVRmwVEIRZVkdH
dHooxZDzCXokZRJt7KfyiGAfQpkfBcG1xpQdHmY7F1CIgtyYKXME3GmDSHZqAF7bkAD1uAbR00c4
Oy4qviGnr1SP8eOAFkyKmDq/cQJy6LVa2yV/sUjLaHEXkyg6dm4DYk8H6lglhEgsCMstKq8I/wiO
aV7ZJUEwoERerfZjkSPwxXpfdPWg9xwvPJ4trenntnnsf2oacuRLl+Dfa+3Pj3l4Tmrq3CTa3Eg+
B99wYRG9nsCh3lRVZxJKS/ZjUycJzk2CJFJ1BI/Q1JhP6VidfKGWy59pqdrox26zyz0ApI5TW5Av
3y1t3UG4neN4MaoN1x84PhbyQx2il3/5VescRyunvCGdp4g1SEDoZsn/ob+Ps85ur0O78LG1vnc1
OIRzzA51brsrgGNpz5sab0Rpob7TgeW3IB3HrNBwa0bOAEegAPNjhqxhp5NHYzOqQBqHp1d1WRVp
n+ybrCpXV4i19eEdSlH3lJdEDlckf3U7FAAyAsVzWDeu4qQPXCRdldC9cpfP98/S6LtwBxPLc6H7
P2+oqug346NmTjNlmF01OT6i+4Ne2IjAM9ATtN5kuhAP/UpRO0pgZKpVh2YhWoDAxPGOXCDOJnVN
XfGEg1lWKnvchzutRkCNJi0XamJUIFKmTXaBXVYKCGDybEr6G3naZFdux5MhnJEXf9quhCphbtkO
ThP6mKFRKtlOJM9x7l3RMkDsZr+5wnQl9Yk9FEYXSf2UAnhnXVWC6uNfxomH5qe2bK6beEmi4GUr
Eppi0J/GOoD2IIPQSgLllB2FuupUCuCOl1/U01T8j6PK0Yt2Qb5V08vNQ5uE2DQPneo0sdr35oDB
hNjUSxSmElT5JUZofEuCbZP7n7SGkV+14WuM5sU0F+UOl8DT+9Ms2Vlh72J7QZzJlrHjbK9s+QKh
9osX2C090mZA+2dbp+b+Ycc1Wzon0/aJdsj982jgxMUnga/iy8yF6MEpUccax87lmd0OUO6C9qLv
BppNXujLIfkvzWxUt+guxxH6QCF4kza7pGOPPGRth0j7P+AWEiWRUZw3WqtFbumX7GLsTWM57QCa
x5AnRU0PMbeYO5iknXyqdJSNHhzig1WpIoPviIpL0mX7by6rGOaCjdlAzVcu43aTlLxrExfP3qfM
E6M+5IyYtHUt8Cae8scGnu56JTd/0akXbrF3C8yQObdLkHnFs5vtl/lxHB91afEN/yvNjq7l3G4V
eBuv+jdsYroByKVxIbGMOMTUG++NA8nOhqNPn+DPPrXpZDUwpwkf7kRCrho6dcXVU4GWZjM8227Z
PrMU60M1hCuU9L6X8ZZSr9ojzmLMoecK4WBnY/Evr5VO9WsGdcety1s5iUO8YYXUBeAreXaBJ2b6
x+HqmoXhBWDe0HHFSzUik/1FSX7F29NwVwo/AuCUxzUXoc7e27OIcLDBLyEWSfJ0A+rYnV+8wFy9
Ejqgx4j6lVfgbKVw0kMi1bY19IFZFhWah5yrSdww/2eZ35+xUJbaYVfxNgNelM5f6KlbSlWiRivM
lmk0hcsOQ/ihSzXo4aTOJvQ8VgpBMapHqTgtTruMNy9hC28nEoKmAOa8XXmwDROU+gjl54WvTbVQ
NqrG2FW8Qrl5MuToeokfmU0KfHW/bX8x10Xz13Gj5yUfwodOPcgV0XUBBlEnxLKvK45tlpZnHAKh
n9gL1/fRVQf7sfZ4Q+Xl+8Szg21zXE+1r3EIwatBoOhB/kghI6MzZMZvAgur3SzUhio64CyTBV3Q
DrLTDS/1sYV0flb9Zv7H+fqLGrx9roU0BL8clGKGU/qXpJJOHKHyvkXiR2IFt6FHyC/P0Is/K1G4
VvFhXo2J0vUVo1xxddUN5PLfa590R53zJFgyNPzE+q5lenYxDpcSoQ7o6vMyfebRd4Wi6luQQElK
c+DYSqEl8fxERhtHl7a+9LwnBJ/INbbl+Z0v4QMfyBx1MG2PXM4TwDlfS3KTwEDj40GuJm9edHbM
MFfDwDbPXFDfJqMZ9sjJ7cTcnsvJ2R/tPcJATs2FEsL7peHpRchdDIcjAc6c7I3W5YDAytpTWxkU
2ugbBRPJ7r8kAI6vExWnh6ZpWi6rwxCDYr8ZrOLHtf6HEQq2zo6YgwKuoRTmDtEmoStVdT2A3udh
58HUQadYFQPmM+v3z6J5dVMSgL6K/ebrdR9yOBevAEfZA1QdDLDPTqWRowHHGUwVNeYgykyFEC1k
2prw3656FuZK+p3EaCPDY8qLjV28nRB7scZUjoVgeqhsBlmHkwYDvq2FV0CR2OPDSn/MifuOfV3K
tb5XATcB/I7QKrJ1CDEBVPQNzNUWrE+zoYeChLqjyMMptkEgOv0eCZ0ROR75Z/72YnIp8SZ74uu7
3TOq+fu412slGxVXTOfwbx3Ht9vGyaWkCrHH+PbTKOnjv9vaoeowDFYXQRXa2M31f4IpswTaBirz
dLTvzxdmQb61zqcWxaTxTvXq7F06sNp/glE3kLuwTgF4Ag1gpXEDoIXVA2h+lw4p1Sf9+kwogD3C
fBF89uYmqmgp8TtBDOWtLzJq3FxL52Pm2ADKdYuabgGELr8CBPuXXiN7C8uXkosyvPMOrRxQaSS0
YNvh2DHc/y0tOdyr7IMc0hQmrkEoU6oQaipW1J5eYL3zvzHdIhkdP/Qfy7VRKoMjp1NpOahpm19c
EsqmTkqi26KQosGDgkxVlLDKWaQ7N0yuCa5RHos1ZyT0wAfBC7xveqWSDf21t2qUxIOHGRiaWryu
4CXAEaRsObT++PnqWNvsrgUhBEa8sxzVBEfvGBDcqNeZ1NHCxorszE6IgXkdLTvGvOuRwMnYDHuB
wbSda0HhKjLxZZ223QJx8GthU/1J+0sYoJgaJ1ydfIeVfaZsB8aAKMS6xlpau3PeskhOzOEmnPU7
TPRMoMo/9DqvNbWrOfqsWjthF1FLaBvw+zU03YNVIqIEcQb3fURny90u064aR53yI0wI+ty2sUci
zvbsK/VC3TcgSyp+1KETZzlv4wiZCZ7XYKfzWOrWCHdIZ1G5fScv2fOHIEjLEQXDXtwvWoRIYHEM
Kxprq0SKHhB7TnuhVN7T40eyLgsgJ+55AKefuFtf08o+0gG+mPY+ZDL1kNZEy13yJ5YEjRxeKh0a
zSbmfVpyTvwaRDYW7u09+sSCHrWWC8mpj2+VuLT7M+Giwy67ScLHdre5bs0Pb1s075FIaP9KtpLh
X7KwekUvBKv+W4ZtkE0tQxGnA6Dlmoi8XUoCINJQGlj6zEbFQ8Sy6rRRBSYS7r8HS95fnxoqH/ux
DwCe6t1e1dbBbmhU4A6s5HnE75Gk1EkRC4u6Pt9sk90Yuiiflype9gZ0rgfX6Sc24IWnf/VKG+4J
4gHVhtNADA4qgelg7rkoPmuenK2FP987/2JLzSwGWWlQU9LXA3QXpLlfoHsrKh3Aue7DzvGCf0nw
0fooSnJ8rcDHwUWwwMWqKRVad/teEcXFuFLKkRXdigkHKX+B0haZ/pxf2z/kqvvEGNPE772lU2ER
OuQfk+DE4xCPyc+IllNgQWCDC10eRIpyoh7WY0KeSUyORkfTGf7LIgH3bJU/fLIuUIm7OxySRIwe
T4/04pis7TYi2fMRjtRoSq4A70ZVPOdCkgnDuw2Fq/+f730CvJtDSBoFusxDvBxpCeEmFoVHo8M7
al0/R1DsPDDRyT1SQxJseh8p7tQ0mPu/yDc6irIspIl18GsFL7mZX9t4Tamxmse3qjP7qU2wDbgZ
+ZhQG+RAOA007jDrIDClmjMgvDdvlpTVrfSy71DoZPf8QJ+BYENFf7mAeubiur/4yv+3O9u2YLB3
6hPC+htOMnC7cbsF5A6r4F3JoymbjgsTKz/hAb814ZnY6AicgxjoGtqOIyKJrsdSkaJrtaXha4uY
EU/5Rl802U/a78D84N5Q9jJj/F7e8xbkstsknpBqOcnS8Ht9GjdQnKd0BElaR05GUMoGE6XlDwxu
o2ertat/IMygvbfn1zuMQCyrIokp+qW0Uo55Cncl6+J/V1OqDOTyS0clbwFks9PwXlsK58tFU8sl
EgTf31Tu4HVGsv0GAWuDCvrBSGpDSQvYzyCBDYXOFET82aQWyo22IxoqdL0Cw9F1r6isnsLN00d6
epS7cNmKLw0SCnkjwYHqtxDO3EUR364z1tG1/gYgG1/G3lUjkXP3Prq5+CS7uDBaMGzFhIKOuAvX
QLXS0bBJxauGw9rCUe1m4CUa1QEXV5gXeilwK2GTSuWjyMuXZonPWHgDOKM8u44W9sxkbRbgw6QC
qYZTq/OQviUhyEJx3DStuk7ZJEa9f+pQKwcqqVIcMqeuWN9HOe8Do9JnNMaTiwZnXGZwI9qWqUql
mL/WCPf20N8w51+/d198UNSfYaT5vMG1rldYQ4jaBD/GWF5c/6l1SI4R/RyJBb6zpcX1s2m67oSt
RA66kQStMoayX+DzmAjB1/KoHQyUGl7Dpb25Sl7CEf0HA0jq2XQZDOaxGRZ4I11xHkAuv1Rvq1wl
8/zfWJLckCdlWJWheAiZnWz0Qr6sRsaeWKG5UFwrIse4AWdN6eEmgxTHMLysVZR3YjD44OLVLftT
aXgIVH4RoPnQSn661HmHZ+6CgqrGcG+mwJv/ETlaHJZ0Ip31Q2lojolnyc4Lojth6ejRkJ4jDXRw
Dc0OWK7o7ocZ+u0jM4tkOP+/2h/TA7Ai7wTP65z28m8b5zUznoA2KWC3Er3r2kbUreBUIlE0WKBA
vwX6DsdTrP/XiGvGLRkLW7v+bLLW7/65j7jakIWh9CTSdQ3xsTDmobGcxCYHw5Yb0yhRqwleo3/r
uff/VOg5DjnnQqFp/hHjqRcI4d6pIFddKvintrDDdaTFxQn+QueczRQFZqmd52Mx6JWfP0nW5LHZ
rJbytIpnraHUk6fxJvgkl7MLOEUt1GWQ5LeQqSsY5vz81l1rfXE0IEEWDyO0fonElrkZX2mnxi5e
NWYVpI0HUiwbML0g43y5WPZxoWteBfztz3h4Yy/GzqRsRUA33DK4cGZNvON5Xo5Yg5jbRBIBmLDk
gAgZHyMZb6i65gxhyqfczJ8f4849moRByKmPcSlhiavLJJ0oBtw/tR5wMKqhGUEcUjdoG12VYsFs
hHrQSHjkJbEbAGGOF3q4Rq8xtc+iJa86N6pAWt3QGxrZe7FyIbAubbx4/jvsyWHf0iQv74zTWFpO
LJYCx9WPnz6cMeAkxfb+b6ENadWozw7woUUu5rXrzId7h53Z6FVaJcBsy5tpA1gMiM2+XrFtihz7
AevIn3Qr1v/iH2NUf+zO7moPMRUFCDHLrk2FRonENjU86aYXxpx/bM5Oeh20GEoswwMabCemybbm
oJK4JPujQwHAh+tbVMby3+RYIXoWVlBvx9OxFY6RaHrfOJw+ssMQgmfoXzwwqbkmjE0DwXDntpuD
dQkIjA+j+eELhkFSfMaZLkYkbaCa03dj3qwxJQ/rzTftJ6bWoKhLKHEMGKXpV3f53AQFhMjv6cnU
vkoiVYpZ0Ut6P1/gSqoZe8dtxRn+KxOkShCiKCqz+vKUjLu2aIpoxj+xyKCfXL7iAza54AsXeVni
dHjJFG/1xzcqtBHPVt6I3v8YL0hKHX5se0+wIPTnyLou5G1jE0k0i9oQQTLv+lfxjZ+uGf+MdEMD
kiav9uCfz9I1X2gv4KE3VdF/giezqJYxaOTKMqEy3Fkh+ZKTYljm0G4MmtIFXXL3mg91J2DLLQmC
7Homb/ODfmMotpkzbirVA7dfKLTDytHPMEpiY1XZyeN93v9Gr5wlNhn0fPq+QaMHEbvogKebTWFM
cDSLCV0f44RrFkkL+V/oL2sY7aH828VFxOQWJaX4uB9NQQK9adlVT9i684oGku1q+oXLUJvvqNyJ
x1IB0U41STlwtbvEfrJZeonII5QetojjkhiNXjzKxXHt6MCnibVIH95uGRYk/83A3GhHyGbG4DBN
qfeSd4jRKzY3cFU8wyxRiORwFwZD36NZ4llhvnVXcqtVP3W0CXmS4W28x0LnwBuO6p9l5aIGIg/s
DmSCiLlRB/e68sbLbIJEaqgu2vtaknTb3ru8rKDqyy6ZAwdHNXDGjvvzq+0/t0qKMdmLLgDKWU1m
neWUxl8CY4XobXw8G/nGcM5Q/ASwhJWIjJrKp+ft3Wc3/l7k2oZaWlni9GIY0q5AK32007j8m09E
zeRkn1BEzZD7jA2Q7PX0MR2QnmEA4C5O8Fi/0kPYxBavqnlTnVqhrQ+AyzFRzDHyVYJOl1vTJ00G
mW0/TtWqzt6sRRfzNJxJ6tBHq/eUwg10YYTcdBD43+AXXTSAkVLawQmQv2e69stFmKvuBUVJYMqw
Ua97E6TN3Bpeaoy/X6uXbq4xqQ2goed7b+3d9yGu4q5b2v8HU9AY7RiDdwhd3DWzqvWEjUSdu5Gl
08GJ5WBMrY41pc836IymPuc+q3NFkVBAFIos6tBnCp6eY6EknrUXyior+CZje1mysFISjfJCiCx5
+WQ4fkny3RWW8qNk9FYsDizX8tHJr6BTba9erbQLKq35z2fAwqlstdkZuO6yE3LubntkRPWqQZSK
nPjBOEG3tXHhVI1ZoQ3UrTxTFo/V5/bpTRcUC8WHvZUQiOeqz3WkyrELMId/FZ365d6TtSx/kdPY
zn+sBGxYi6OLVuQjAfe49Sa42ZHblnTbVEOcBzwol3JXN4vJ+XBMX3lRs4drLboA1XHUPq3/vNb7
R6I+2WnRgpCT9ETdSnAs0pubokbhQ+tiTge7MyaYAZwrVpFrBEEKU15I2zBghCzvoHpm7HjeLshS
B7HGBw/4jkOok98CWzs4tcymCRBtbKp0kMIK/S7W2ZRHO8IA29bVcT677C7G05up5HxLnehqaz7u
fJRffoHAHEgxIMSf7Awvfhw8Xe1V2178JO3fbkWWEurSiO2vvNw9s6aQgCD8qnjlbF/4GwySCk/A
T8hp9pY6V2Y9UhZoUgKTbCOAba2lQzE+8RuqXRaF867wa56iNm/Zgax2+VeO9gEHsCmqk+8LTzjv
/sujtbkzoO9JrZrSmQgXhw57+vPB2atSUWWwYxCMTj9g7FnWbo3LGkPqz9COyEe3UBM75UxEYqAe
uqqVfD6E9v+vbwnsnartJxGdKVIoXDFKeARnyeV+IyuKMb4vM3r0xNpqCib7+qGH8/tgC/+8fEgg
Dv7eWEx1QXwk2aRGm1EmLTO3k8GysaNpOf5B7HItB1J4XqlfpOmYyjsP5iLCeJDrHVP/Nm8F92FQ
FwwG/R94ycl6vL8jCR31oAMa4ck5iFZP5GnmbDox9YpS8VZ5D0ftKY/AsIkAWspBiK0k2U5h3gwU
H+Bj3bgZk+ADNRqN739EswOwpYq+M9ETXce+UKu8X8iJ5hiEymn+MW3s6heRxNJfN8Nr/vvlDm3u
Xbs5kJumXITpDU0oNl1EaLXKYgXuKdMZMi2e09nfoNpRh4dKMFrmPB61ft9A1zG0it39Q1/ubEYg
qQT02Wmea8QdyNWzWYJet+/SAA9pz7GcaCgUrCxIz9at9unrAHSP8Hq/nuJFX1FMcQ+KmQMf1qDh
RGeTUJ+BppmOuZft2Eyf0xjMfbTmwHAVJzpS8HCGf8g2/YNfUoqJRapPijiZ2J0ySaTtFQjarJ3b
xmEHSbWw3p+kJWh1nRG3ayWRc4OA7QsgFFWsAw3Svb/FH/OLflheBmG3Z4HnSlr3KP+6dlRUi3lf
4F73Qs5er6XO8NAQkjWwrCBmsV9C4DdntFwIuOrK10Fq+yb7ESnf4mEvXZPPeopMgUpyIZ0kEd/p
I6kOz68W0/R67ypXv6GzMmQCzQctP/u81Xnjpm0CgSkfNmwOJr6Z5FYriJ8nbtoV1uJzKu5jeQNP
J4bUfjWIe8MANeLVi0aetwO42oekvC52U1ObrK/OOiFA9R7Ro2tJOVaj5ZQgz6D9BRJ7lAbMleyM
MeCLMKZgpQf7M+wrnhd7CB+Bkp4+hTVzW2Dg9TsCXneOJ790Q5Mxi/toDZSjJqZNYq6c3urFEsAD
IP8KPJ5dwthX8QVFL/ToxLL7l7alBsbf9idFNJq7RmNwDff2J6PqltxUhVTy1Ps90GjwXr7B9mC0
L7tZ1V3DaZVl8PJIVJakfv0Uv9iOiLA99+3Y0dppnyWlDIa3O8Jl8JRCMRcqtlVlEUyLm99B5Lz0
QW8s2PpNXF1MSbf5nzZPWTbcpq2vLkrebM+wuku9deH9vBoEh7tao/QuEq60yL+flM/p+yLEh7TT
KLl24oNCpUfFc/XaZCp+9blv6fU4eI40RjCCavveZmxZIGI6mnle8gd3y41bIMh4QSMi7uOwfFOj
q7Qabbz3UqzgtjmLe+MQkMFKar02g9E4aRX9CHFGVeO6N+LBoxsIUGv/y6wSc60kJ0bDwtBz1MM4
6TIkOvNBqE7X5KmZ4z8yrVSnkXoglFlNxoWz3/Chz82U+WYKJgyy0lZHpVAB8o6uH7yWPFdPZ8fg
IzrfyDJ0/EuSuINYD6NVJuGR4LnkYyrUEjo1SZB3oAZFLyyQ4m80qylP8u14sCs1ATv34uUbAlHv
FxqBYWIzne/f6HAClg2Phf4ami18UQ+k7WVUJaWiM0nTbnJ2CJ5LaB+Om4ryHZr+Eee3/hR+lt+S
Q6WURZt4HsWIVzS8qrDWOi4Mtr1QGE4VvYXEucaiG0j9cmDa5teCjYl1ki5xHD5+gSAq7qLduKRw
5yGY6QBpbEcHkOAyDh7f8mLTjuDCaGPfTa2vgfRcJgGE43iufMHN5Pti95UNWoFDquA9qHUSeOhk
a4OOKpDqLxbLJVCTlb5DQ3xd2fhBnOVwJDutUiyydWqiITd8XS7s1JZ6mCQuoCZZk7ti1ZB1Jse+
HvJqSwRKfkdVHhOq7eiKj3D8MeHuKsIlbr2XIh8O/aDIQ7TGSaeqI4xHD6kK2ApjzeQ42ZjswLh1
eqvWBnvA4uW3o9iljWIlMCVl8avwe9+sbhI05r8gcMTDuaoDdt4edTfB7HadmRjiuS34+W4vU/8K
aSgj0VUrrx/8cCGTpwnWpL+8uqTSy2+W6ad1adiyMidaLeMcg4pjy1T1TkiErwFmqYXU0moiEoZx
IWozLlCKEA2sGswFaF+R0ZKZVC2jC6I/0vdzle6HIZDTrEEfJXa/b0iCqH1Yfpy8+YL6UlIclhQ7
GwD+iq8varHq31/Qn1EiGiaKHt+OZSyOckL/Fn/5Pc6jJXW2uJhYrEDIWv9+VE+gV5cJqQhy3+li
PpWIF7LLVNrwAME0rDFKDf+kjIezQRRReZ6oytnxsJN6/Dafokp9E+tqVPpKiKlxgJ43W0o7xhZ3
ZMd2bGn7uoGWUQ9g8G1+Jv6xpVt9MFyUp3uxCVtA2yCNTiuE1jmGfT6Najnqtgob7dne7a8RcoRj
QvbTcBvDo7eBy3ueQ/kD+l53UlXtqCN/wnttZKG2EQKUbUrr802eEYiyYAJMXRzSVodTD4nRn/TQ
C8AgqohqXELXz6HLIRejGhnGV4F201A96opumSl+8tW0HtUsqi6db1m1hpp4jSQVbMyFPU9WcsF1
dszfbG1vscLYD7PTtKoheFvd9vtRGM2JBmaKwAVQrAwCSva4BdSgWlHrMC/s5bZiXWpdUbFP8dYj
dIPtP2hzgwftDteezV8BSvq0sO3fJ3hvfdsNlB8LuFUqcnUel+xz/mpriyj0Q32N34F3bpMGxrFO
YVx9i38X7nLlqkz2HMxLuUZ2fedMEmu5YozgKvwMWydU9mYhlegb/sk1e7ySjEL8DxS+X6WTDBx+
W7Uk6iY1UiL9CgvaMGA/zOC2rJYLxBFXUsijXYYCUNIHYPHiBr08vW1FezCDZkQ8ffQXym9g83w2
pMrG1xoXcweI7azogNfhb+TcMnL0Jf9qHEbXBzKZWWjtAJ73r8VlrSeF3jQyxf9VbOtyT+LPg8tQ
Dm/b8yDmzDPd4nKLqlJmR09cutaeSgZfMCmUuS5RH41F2F2yfxgsq9UiAoPUqBZ8T6SoHWOLPULu
wEk9j77U/NnhFf/cNIJslEQi1bXHfWynXcUPvDWbmrq/N0YLYiupFcU3Qchw6JiteFJ8hC/pU6g7
IAjzv1NW1qjtMjgNLH/s9nJxBL8SXSlpsStvNuL5dEYQxiTo9bVOyav0rTP5Ny9dzpW8PiMYoO8i
puwG+GA7DNbzVHrZL3h7sDs2uubCtAIWR0ahbOO6zOytzgQjUpKtUyBt3d19cSsxQgpcrf4Erthw
th7n41iyxW1v3Qiw9urk8wYvquFVpIWVQckgo0vxfiEJ+X1HvihizNXK+mZLroPsehQcIfLuLde4
4oYiwnailcL3UJzhAaMJ6hmX6GKprGlBeBQYXLhE4Phcn+nxYULidWcIzlOut2sg/rubfXHnvCXm
lhnCP1GrkeSWgXf+qDw0MMUdGCHHGtVGImq4FvZn3ojzhyJiQS7U1OzEKOL7XDutq2xOHEB0iedW
Ep5ZVBaHXUyqOkj+8eP+HVqURnzdtbV++jZKgNMUREq9VLqu6BkUipm+TXPyUsO82cj8aa3GSmah
NeJq13lUD8m37W62JmyDCx2qdli5otZnwY8s3pryDr7X7GcuRbvzMXPNzRz5iqxIEUZ9bQLyL7TN
2wZqptGhHR8/GpNvO2/vsYeVqYblDjopiPGTqZHHtZAgC7OCeCOtoNlbXT51txZdjqaVkfWZZWrN
XoUB1b5zKplIUBLBfb2Wo6ZE4N+a2ir5jJ7m+35K8MnU+xnHTRk2kO91wg5bO+JtELiHr57GW8lM
rWfCAy7mdRoZfmUNIvhFJwTQmSnhkN7w2YKJ4rBJ16xk3A78+aW5nPHVTX3DMmA2GCM7SlI/QXhY
0EN1aDtJ0m6nnrlKEBbXigqxEloYI+CCiM0Cs3OJDjyzB3su6ipFCG1Ht5bv23HhxUzoN273TvWv
s2Guf4Bovp39q7HqliH0fIJbcRdwE8RtvLUuGQT+OXxHjAyWXIeDqp7X96gEkAe2Y82rMWlwUw0u
rgF0vovgUs8B44pERVmXNEM4tgvYVg7791hyM5wxGr7YQPc8LvuFZl8bHj+RRYBjcrD/ygZaPcsA
6xitVJqFvVETj3mehY6Vfq+9Z8K7NfU63dJOyeRvesluaOM13m3nIfkUZcCeHT90rYH37fQlXB32
MsjLyvkbZquJFb6/vpYtCSxXSYvJMRyjrDAtqqQUpprBwJfQojJza+vDSw6k+3MaNmIsH5WnjoWN
37aFBO63/WCpACTp0OeCOEelqNSr5OcnPjXVpDFnIWf0w8VHq909UmbZVVUdTwBthkiqWIidcBYq
HwzqL2j5djzCJUoKNHNr/twLUu8FlmabYdrdASKpPwuoby1QrRSJqpR+vYyMhUBjpLOmtDLel3h0
wQiGQQH0Cy2C0e3cXN1Doyfhxe0aIDxLNs9sXk3MgsCLve8UeBIeBcf1YVNs2iP4l7DoiB5H353y
6b6rdEHRKDeVJei2ilFUSSMPfGnsUSvjb6ts27CVibOGkMVdKrTP8xiBjtOMiB9ZVJJasY0gB/tj
d0A+e3GHEem5MgrB0f0chSGJ8PMrLRwhpswtvUke4lgsdlt0i1NXWfFpXibpPuQlajp/SieVYjBT
Qxv0s1ljLbw5/LC7wxHk8etKP8A0PPt+Qrfuldu4k6w1cO/yGvzly97CvwxNopDicdqiZsj8t0LY
v4lR9fHLvKar55+Vdgpii+HNQhvGVDcAUNctt5QpSZgBcMhVhrf7+dL4gp3R6Tq1DjBbroSbg9fI
Ge9NtyNE/5P4yWurr8eUSd4IA/KLsbIWS8GjhGPFxsedCBKPnsuhPMH0rb/+j5AT3/ijwtvw6kh4
HG1142e1pwzZW24XisdApn7sihXmYUYnIAWsolY6zcfUxUgZWsXXWxE31LZBkAMIahbqyLNeZFz0
EVmI501jUtyJuZgtpuGpCgZEnOdmfTpPy5Sik+/1fuA5XJi2l+pTYYQgePvkjP+osPSkVKLV3xKm
DOSLdWlpGyTBpxmfe8qmzG+qcbfZ7eDovkCHYsoeLEepdgkfWsyj27DeY3UK0hpSRvRxu5ay3XNF
sl4e2VALu8NrGm1NrhGSAFaMRSTOraRqSLI1zmkEx0uWvmc6ncJWbt+e57t/SbwWe65DJE/H4VnQ
oA5SYS1NFNgbUGXTRaqTUPDyvEMvAtAJW3Uthp2Wbt7ZRdMAzXwXL7tlS0OJk8qCbC2bk18RgrL5
GQ0Cd/l+E4hWGZ5A1WNMpnQ4LQNqLjEfgQZyFYXbEVww3Jmbj6JQSLorhEqpi4pdiZyLbfqehIhu
plvjDqjU6XqWqKArbs99EkAfmrA5Imf4NJ84NDTYatuTU3dWHW4G88TmZw7Xw6wXE1x4XdGhHc7N
6oCXrCLyirouYa2gNx8Gc/XyEXfU68Mk6EuRttPuop21G8BCpCC1O3qG19fP1Zho7A8J4EaIWTwU
bKvpm5qXkpZ3x3qbSJGgsTdjl8GN9DKNNe/Uk/KEKJv8uaaY/46LfCwy5/aNHAcweYRbM52oUg0U
JaDL5GajW9MsbKrWu8OtNR7HPMhKhTLhM/Q0La+Lke/xyXSlqMNMnMnt53u08XXJ0X71aixOChII
Qg1BCXRvcSWpjFAPO7GyV9hKQSVgK4JbueuBTy4P6URK9KZNy2bieWvWyK6X1PA5fJAtDmhYj6rY
wxo6sYUlKRLay3P9nXixgPHUchVAAA+F7c/t3DOvrwqZjei40VidT4HK8AAzQCZzkZCVOHXFq+K6
qTNYrr8JqMk7Yqsl9D59pclrdbwtJUSPVkdrzmPTYj/iohpIlpIhVPccXKFAQrSEaenJeB3iuBdx
JylPCn5IirMcOtmnDz3n8heQwnDJ0Q+2cfWVQTEGq6JmQB1e8E+U5j2I/QWwaWoxIl2mvlk8SLYN
NKqxEAc2lTLfkPxiKIStbSUq+2Gql2mKRyGLQCbsAmW5wDg+7COvyYKxBAkY6baPM9FpGIP4S0OS
4jeifsqWu0nDTQ42t9gsF4g6LhVXcMY5BBKH+PtJ9BBQBqy2GGY2NHzOtpHQkHL9J8D4xsTSX4ID
qLfpsfWY5ZEPDIOhBelpdme60JiRD5gdiThekRBcoFyVFWS8BXxjBgpNZoE1m4fHcdpsfkMayWVg
8cOac9BjUnGHzf4bszwID3wjb5MCc7ZO5z6vKeST6JC4hXG42t0qwA3LsCXYJskKeGdPeW9Qteck
clmE0oe3R9edWEE7C+pl862dmBNdB7dWkREZv2hP0Fl7uCm+Dd+34VvYJCVoiqR+GxfGbzD+XEam
/Ulj/L3A1e1Vk6/TBu5Fdbb3qZkN5mVPiA1sHqCJaK499qcAwkY2/BTKj7QYAakrAyu/iAZCHMWG
rMAnG+voMyeagmZt4PlDA6KeoOdJrKXGqoEqjYDxoZYvvIB33kqLEfLDOdKc0e+J97uN+zd0+V0K
QxSOoplzZ6CPiuWi8TggSpuRhuhfYdAzdHeckj/YhZ6fS1W8x1/NVGFHsc3cR4ddSGVFGPI+mPnf
x1jtYd5rc0NEQ8LO4yH+0W6/ZU4R1WQvnLgGdzDyR4zHKq1gIORpVSdCczURfoMQGi9Jrs6u1AIK
ooXsNJpQtdSOkmFIJKsKn4++mguHAjAK+gf1iCVcuAin07E48PlpjqbXSW+ECLmxhjvbipyN/g2C
6mKK0CARypSJDyzx8EOZfOHJKZddJnYUtfh4G0E+um1Dx7FeIXEI/wvB1u9iSxS8akLcjBiuXtF0
l8JVWbLauvvbn9FIZVVxe0+eIBrrH2hLGz7RteLdVAOXnmdzu3bzVgFUoLOQA1Q5LbynqWnT4ddo
bsQqQC6wHWd+D0X6IYMlK047u3l/IUijyK8wrp3hIuszVEeYWiTyDLVHjLm7+ynsd7pPR5TNb+1t
ioyn6vOZ6gDk9TNGJbvGjZS2Ruc1s4WqSQ5dHTXQSQ3owXFsZmn3kZUugYVwLj+7GOPa8GyjTE6O
cXqFwrgfeEEHlv9o1p9mvx2rhCGChSi7rY1wbpUlH6ExyUCwUQpcsLZ2B3PFJ5juzR5TFrLmvo2n
KDvQKHDkMPu3q+lN40F1bi/OeAn3w/ABhV1aVMNMeZpp/eIY/SGhg3YDMclWlvVqsx2yLbDKFRoK
pzowsDAClTqBLl54p/upSkld7kjYLxx3NmWbITVZk1b6BBWjKHxow4SSxe1v5CXYr591bk4IKVGU
JIuXmMhogPkB88YgLVC7PxM+n++hANd+P5P2pWt1D+oTQDNA84cOhWoDb+YTCzDGZuNBbhcKtZjz
T5m/HsyXTKy1jTZXPofmhS5B+hhJh2gu4u7xgcPLiraNWVa9mmZvFEy9wLX0DSekrBUuvs7Jfjfn
J2Q7aEwx587wp2ztuoepcJRJ9oBrrJvKamrk7L9CvibDFc0+3nqyIf4tGJTyZgloQ65BwCEdzgwz
dAp8cHnnbRYpAiamkcp/zs6bZXEOHjxd5kA1rlEmAka+MTBAM3pWn2pVdDZno0HymAHCZwf7Xnw1
38JxYLMPDGpbuDawf4AnHEWbwzWWsAWdMCa6XiFEKRPbKuTZH+6RhXH+9rVEUtLrhF0yQyJHWNic
giYbA/QDYokGpJWVTr7N8J5Yfnp0FvVVH/X45SB8tqOaXhRuWIXbo4YR4FtyZvluHQ6bvzw6kiJH
f46RyxpdLxnI3uf0pu2SguhXBpig3/w1JaTdoiJEUQew9L1qtHFtGjC/X3u+zRMwAdEiLi8vAUKj
TEE8zscWWvLe9irDYfqIlMbniDF+rRYbcjMqopl1gM5Pv1OlyU6zWcTkcplJhzhksgNL1jTgvxpO
Kv6/rUXYvM9tdXf28/7lDzLA0DAVLqRjesfN9S6DJwjeP29XXChrRoBbevoaRX+7smDB3V+CiZJD
zvmxio7sQe8zYZAxw690fOSfDd2PZ+ySl7kG/vrSlb69X3TNyrwFwjZjsJCLHsnQJd4szgNvb4oW
cxyCKMkpd7DnULF/FLgDzWTgaDDgG2+bip2GM5R4nnqqMrxVRdThu/bycoGpmS74vSoW4bnv+/n7
5K9y64ky8fUIuuA8mgUcOtTFNjlv11wa9yt54//mxlzhc4QPeMGCNVCrBHxP9C6hgZqiRbluu5iI
SLArQzkmxIaN2tR6PKScEQJ5H2vRCjaN77G2H0ixjGXzOFWUeKIZH1qcYeEGnLMD7rnSPg3AO9DB
WYohR8WmPG8xXz2CX6tH0/jK6X5EoOgw4Kz+KOZCB0xecKziy/uFD0BoPgvPqlOW3IzNOq9tnOJR
MbY0q2BWqepIbgHwNLA98Uhlx8Scn0mZy5DMZU2GAWdwam6H9jP0+EBFqffjehFTTq7kY0M8wSGQ
SNXB4pL4Y92xPMmwFFCQzQwUna2oy0scdfOf1mn8IPWet8GApofgxORkmd3Ncr45QqRQLjFgzPXL
aWYMepyPVzpJ6MpzJUUItnvBZLsPUygbCV1W0QZ98TF5nhoIezm3sfGvbuFXx3Edc3PtI7iuj1Cl
ekMXJ8hauy3rWvMkEs/2UWPXHG4yKDcB1xe1sLwXmVk9TWKjJylW12iC0RiQlQGWllmvEpjAQEHG
URqFAEPzdOt0GoOTvbG6T1BXugUxtZXyw44bGPPBZC76h7ysYwrLNtihTpv3/6c85MC177V3NQN4
5/iTafwitH96ajB3dUgHOA08RDUPMqN1sJraA65BiPXQQnxBTPOqOtxsQoxSqFvha3/Uyv8p5EKZ
fU2IMg8l5sw3koj4KwifwffhRRze21CPpPzmc3zN9xcLzEBdFfnJxKSK2l5lPl6JlIsXtjb7lLcl
b/qkqXaOnw7eq+E67AM4hYVL3BjuDd78TUwocCeIJ/XesCW5GIqiUnYrO+BwxcWacjqHEipgKbyR
niQQZLkAIrQJzsOA983ZQpWlph8inFDsLL5o4C7cJPRw9IXNc8B/9sU7sC2M7yB/sjZuOTz/iYb7
cjkaVa7tvnq0LKBMQIMFaoLQ5MiOegshhcYDQAIolqsv2lmEkjX+zopmVHev6VWSiaSF18J77ywB
fEZSzppEwlVPGHk87kAOeE2mO5BnM1Ackn/f6EbDNChUhBAJncKysoTTRnY4WiYYBQFVCUJzYlWw
TJHz/PyV+YmuJHOdjC7qA86aT7C545p+yl5mjcIT74P1b65FTQ1m4Tq1fppjuzA3Q/OO7dQGcJT+
w53JKaK6+2SlaZj8I9Ql3Qz63Wns0D0iozaFnIBqN8pOQdmhsX42+hYUebXZsQ8sGFEijfRL9d9o
AGacP6hrSLKS7X92vjk6gX1OXzwCPEmMlxCfUvm9Dc46Dqu1cfBIPDDLTQ635VorCLQS/nFxW2hI
5yh+CMEsnoq52CXW5ly0fepYNu0KtMMvHB0meobHqit4Ou+nkPFR2i94pOtj7q4lMjsFx79z00h4
9vLeXNt1yYsG7zkIYC8NobJxtLSiZ7PUr/PuiG/wT/0UnYFXgRRV9rtD4FnovrqNOwAieDiT1u4H
2EavtacXxH7GFUnfsUSeN1OD4ibjrexmGPZaUuGIt5tIMyWfr5ciLMDOy9fmgIosqok/GxE7Nu8t
kuA8iZnWZqlavoTSRUn2W3+0fU/RJWeSg7bGlqihCScosz/Y+nAq7o3e54g/b0wxzEw27FNAodR7
TAlDsABdSQyNUdWIsP9/zaVj5d5I9pVx0CUToc3PwnOxDKm+omE8mV9c40MKeYM+XvahYkQAxExZ
qkdfKw3MLVYyQn2T7VxlDmc/qMT1D5ERHMnR5WzdHg63cgdV1EfsydYMJ9xuAbgN+b4SkFOoRs6d
vguWR9LQc42WfCgjF53B7zqdI8Vu5BoJoQbBPostHnmFytihFWtfqd8qSDHsoukS+XgL9hw1r4yK
Gd8YNb9LoE3yLjiffamkaxXc9Fo3d5/ix3u7ZAvTddeBslLz/ycDlOSLP4O0h3PtT9jnfAPgzyL1
Dh0eGwWQniLguEvDdY5jUa2RpJlloM8dV7DugyUG0y8ADGZER6sU8cDrfvwwNbPd2rp7uYyA29pb
TLRfGg8Fd16yGpCKCURJCf9EFzIfj22Z79sv9fCkqu/mCyJc1uuTRrH3MwzrEFJjF06iqPXXYXgv
uLcoPvdHBvXPX3glnee9arwks/RorRbXNG9rYr+Q5Hd/UZh+ritbHXB/oB6wJwjZfjADhp0ksW/M
gBhRWOqJFWC2KtAFgS0z2Ul67rBxUJBSk2TzsbR2Gq8HrhmueYo/jiecd5Ig4X5CdONoe/V7QBTW
eIBhSO/TXj6IuUtTH4BKPHig0q9/McKNGfoMRvoknu3u0F5+9Gr8hm78F1/3oT+35YbKWgBrNOcO
DjGPSe4Vs87xGwvWnm18fnV4Dtbub3fhLUpxXyjM2tEJUQJZXP5D6CgXwZtTS3+wnc97U6w9+A6p
gtX4ghqYWox397rRVVXv0BTMjkm8nouwY2lD0M53lfRS9yA1J6VlWOhYm/Djr7v46wPv4+Fe1GUG
zx1tEHgHcje9esWaQwhy1ucegWggKnd89yjwXXJE/JjIi4MvOdfi9sH9J3qBBromaxlYLQMdvvOt
b6VPSzVNVQkDWA6S3mkdpM/fV0LjLmxCQAX3ACYBZkZJe2ultA9PvUc9xxiVRUEOGSNEpKQ4SlNr
to65ZKU2BPA0ptJoZgyyyu8/FyO7XvuVpVo204L2cv9mpkiik19BmP8L98rACEYpt43Wo3+Ix40u
KIawWdQf9QUfc3KRIcazVaj1f6QLQ1sUWS01vCCF765qnI+cAK/qh1eGAy9FlKr4EOKh9k8AQ82n
pCBVt/JCm8tRJulKAUKo0hiBW1ca9BFhCeFYwsLqfV4ikGLD7NBB4tno5K2UobgGanFw0kWsLYDA
DcyDl6wSjBBUuz/SgzDn2y5WyADtM7aXmDirTq9O+dt2C/wBDaPXCvim/uuzcYyy4rvZxvLhSm+f
j7nhaXMKcm/FnEgDyMfU+vJSntmBtUS6aOvO1Jp4+SN2C6TD3lGN2Tc537KKJ2I/ohlq28qF9Df7
VrUddo50p43jSoVyKM+WujfNOShgKl5Wk8zxE8FUkS4pBYtsumhO4ybASzQC70mOB2MHfKqg5n71
SFwagdrqDiTob/++1FbVuxKRx2IlmVjchgy+S6iFtrvAAeOcPYRYkFmE4B+k4xZIQuJVAo2MAryz
2iRrgMeqBcb1PR2J+ukCuZrquYykGyWLicBUljOnClbN3mTYqxlrricPvqtZG6CbNvoN8CuAfuPV
E6Ro7QSKwlW9YLQ0NldKu9uKTi6X8h1B3x/JhndMBrPUyqDHVwLLR6MRA9JzG/BV0VfVWGKVg0cd
izt3abs9Q4TiXUAA6sNNzNt73xI0F3+hI0K26zARwT4cP/NZCr1i7Xwh6Pna3WmeMNT5FxMQfn2d
XX6MTvvmlJXGmUV0MFLwiGvYz2u7L2V/9CPeuXLsha+ME1Ki3LkMOzvRqtHD1fG9e4VOQEdGLTeR
9Xwzww+TU4ql2VqcKlUfJO8CEO/bpwZ7BU5FObsUSNS1cAsfkJwtSZ+csYSnzxGoDWV+YrnBqBQw
GiN/CYmJKLirpX5zLBYa6CKF4cZCcUFFCXw5Sg/PJUsf6TVCrFlqQLvBQWQ8Dblx+o1VpXSa5lGY
WsYtWLxnnNwu3QDHDMfeZ/gKy5s5+xrH1OESBlU7e/4BnfjpMGlsaOdFd4d0XTXdc4rK44juNLOI
rbwH+7sXIoT74QhAWsBQ75LvcTj+gosKCbHiMwLaFK0l//uHKsHDuydrIf70ICdIc6Lu1ZvMWsyF
Txgm05pht7h4fOp5hZoUaQFZNLM1ynK/fyWzBNymEtpz72OdZBKpJzb+TDTesuHIHd+xAnSxx1Jj
JZbDhSJTYrkJw+HyZt0+vYmfltRmFhPByfY2X9btmRgZx4hD3Ey5aaJA6hpWQtrJ53bsAwdaHmS+
dQ6yz7ZvW3c3SknsK6ewUwzyyxuNqk+b9qfV0m4jKFa34saEgVEfdGMsYY5+Y7WW2FlqfNcZd/Ox
FroOokOkqdWuS7nKpXy01lrJmiXNW7IseV2wze7UbJLM4KJ/N29vIhal46QBvU/Y7+u6Sl8CCvct
Jm+yF5xiAfuZ/qo5AbYC6lsgreYCJIBYFg1z28TSkAH61Nx0QOM0xKr7xqQiIk9d/mn68Ls9UASv
M21FSIDfs0Ssv7w5+BSzJ9SUV5G8pUJWJiLhqL0csGhlyoyd6ohDzGZuIE9neQIfub2EaZyRy/Yl
Jbbaal8Iwrg1SKvwRjyTAS8jrhIlqidO7llyNfB3LktVzTPow/TKI0Mz0M6yZouUFpYE3moeHUdT
987Lymj6veY02J7yV23jcK1O+pqeWVnVPBpXiQ/XSDzCGzQgBfqKXgVl61CE1lTyr6ZGzpSVQ8Pn
/JpGQ5Y+WSiggk+RThl06Tz8ekx6Yq1RpI4MP1Z9fpNQ6/HiWu+s66hDiAtl+psfzdtwwYV6O2sM
45jj5oNYzpIodlg1cP8OcLdIPaXSSx0NdWuLXQpIztPBEJPrfUHDv1etfV3cjhnYOv6ZdTg/4vsQ
tGneqwzn9PY9ejOasL4Z7HKHEV1TzBpdmjzUv7gNTgA6eZtrMBZEbgtWQdi/p0/DMTQdg570hjw/
f5RRLN7L+EPcQzn/DDoS49FwKm/wjX7QKumHOb5z++2puSF33TmSJ23SwYj2r2lgf8+Oi1P6QXsC
SO30fP6a0XGsgcv+OSpHXDzC2gm22600377GyVSvCzPR5oYS51Bg35hjGz8I0m4gpWGuRhoM4LMA
CTIkPYo9LjAjnAQGMCDTN5WsxAOCsu1lXfjzwNOzat0kulRalgwBhK/y7iSxz3YBlvRmbljfX4Vk
mgq4sMk115X9ubH7M8cKIZltztTm+kJ5jsOcbAVPIwCIGWtl9jLgrS2z16kydfy5ZgT4N4byh0+O
QPVkBni+J0OyEegqSnowG0NNgO5vap4EQNabf91kJzHcfDBPMhjD4Atn/ssNpMrZ2l7YcotPnhDG
5PrY7/vGxiZSooW90lUMhkYtJkVAGv6ngDR3EY4SjH+RxBO77uPbN5kPB6Qg85tODGLOrrOe+WiB
FXeaLMYvzdKsR7MR3EaLYLfDAkyGku2p2kL/Fel7pp1mM6ehxClIefe998TO8MNW/28CFDtfKI3q
9Vcfm04N0EwUNv2mTLENBEftGszu7Qre95CzfwRX38wRGVjsS3FzfkBXhxrdjtTI4ixGTSgTzQaE
97Pk4DsThw/Tf9sg5ntQTXrTKbgtF2AwT2KgPg6Xwka6XIHmEdMj8JLItvjpeAGPYJmL2KmVE7sU
LkQUloJhf8SCBclLyD3/hxikQGJP24841L5J1cqIp2YHBCsAIrtyYPBl8cQwLXvuZP/0RTO3K8Zq
UvsIlAM3uLNtVC+v2nh9GJ2uslJ68+UJo7b/m6eEcb/Ig+1jm4TDNyqBJ5eFs+NwQcDw/+4nn2Zg
y+dSGe9SYLDV26WAjIApVKDTDdOvfTi436C0wYAboPa3t7dwjmA3C7sJZFNFPffvKCXrbyQRzp/I
PSW/IWbIJLCWMx8jc5P0jkEXiN6G7g1O9vJ8HYH755d+TcWF5v+W9a7EdjGBjVSQ8o0SCkLLQ+1B
cvALi6+vWjFcgnwPJsZfF54E9WAs5FyiOvl+rbcOgIP4VGcuY92tEe8fj0AHdBT+W1/rxCsdzwld
EDcmkqT1VXCyIbVgfEd/2H6GWlL86RgUpBytPidN6XVrPNiD4uI+KogINAmXkbVP0TkwpQx8U1eC
PeWMiRjLCwbBmewryOgX2w5o9KSDKh2BtLlMQVSSFophATeeAuG5rtla9Qierkuif1HxlKaWVhOS
n93juCaHuqP0KEKF2l1IgmQ/p4oQH/tt7Q6IIwJhDdTj4MYNai+xdPRAhWIII/Ohhp1kFy5IBzi0
5tXA/xRNFCVFIQOfmtkt+jMkDhQ7bnYsMdz42WBPYf9Qioer1IFdLvSBq4WihjkNyqLwu68Cm2dB
D8YGTPtpk18eD/en/S5XHBbAlD/rEnaYoKfmkCN/gtw4sc6rh/i0Jd859h5LPnCg3P1pK5oZ6Aki
iI4p8zHQySyYlXq7/KBXZALEt8TNop6seir3nAhm5nN3E36ZWKkcC/NkQJMLBP0v7PsnyKH07IRg
d6+8vmx0/7c67jNHFqfeOIHoE5eOQlzBP4wx4ca5aSXpANXkIwf+HjNU34cKa7INIOk4cxSMdo52
6xaG4xQbPIav/+j8IPUZvTodyQaPqHASy6DdQRBixRtKHb/OvALQWakqIAXOoq/fuyK79rv17VVQ
iFnBP9LlkViUoldo5f0an8UMqklw4FZkL7JR6MX+PkztJLt/TtmoHRdzmL4uZT0t7RQqTIgq/JMS
B/py2cBdREP5gqa/1x/VMhZiKNI5k0SNlllJSbWI3Y0BhNI0SYBy28QhV0RrqNlmTzFtksRu7xub
hU7Ye0fGyJBMFBZNvbt+skgoQ4K29AB+a9EJzu/Z0FaWTs//9+7JPC83Ip6InsD/r4jHFsoITFtp
KkuHyZdnGOfq64n6OWIIbNxfCMcirvyW9OQaNasYvC+Zqdg9Mgjg+kyV7QZHVHA01e5BycNObvDE
gl6DUQJNooV7/kwAjTU+Po2IQRi8frrXs5SAyIrVeVZkZh/meTCYJV1G5SJKg3pDEU+GVP4CNCDG
j+ulsFf9agemiDDVEYhF94ImR2BRW5zF8DlRAWqWoeUWbWvcvsjvD7uTzd+NYE/LmnydjO1NSFkz
E+tXPWjZIy7Z9PRNvRThMP6gQu20xWl5EQvF2BJ6CLJH9b7SCFArhk8Asj1iwZ8a0DfGiszBpdSA
OpS0b9OWcnNZ9tv5t3cmCdKzEAf9mfvh5mHqzB4KZVvrSzSZqHR5daANAQhXlQkvyrTqoyX5CD5m
LBokx9YscTxDvCYvkcc/wu2SLULAQ+A6qGzVuSTgrWpSWuCxd1ev+/Eaj0VOVpkcjK70uG7hJA1D
mmVxvy7I+ZyieQZTXiMYt9Ij6huJwh4BfPLoRApnrpo0Dje/CeXxFX3FVl0qZJkPrLrcJU+GL4FC
cRtqxHvZbCLdCGttvs9ZHfpViKfCnwk3/EYFoy4wOrFeGzG0OxalNrRjkz7Sw2obmfgmOjdP2Mig
V9g+JldG+JeLk22Dk/9GawEV2QFRpWGeYIMB+k1WIzgyctl6GXJwZwzTQmbzPe5buXL3Fd4tXXiS
nz3w5hKZham+OYrmjbBuu45nvZmjYTjkTS2nB2PlckCtcBadiefcNuftq28d8WDxh1+S2fKjiIV4
dF1Tc7ox5UbMO+Afd1x8xlqpFgEx9Wuh0/0vPVII8Axo52JuC1nzKSH5BpkAUsGHu+i0TflfrdX7
4kpMM50hVjNiyB+cCfFvG2OOxbxRB9h3rdFMnqyLOD7/hWBz3lQ5bDiVFjDam2RFvqis7LZ6ipEr
K6xfblv7aYjllrHnw9HoVDFuPojRK4oGlpJa4jhgBNbBwJKl8PZyBumCKRLS14XtzFZDqEXP4Ysv
1JrIZ1BkZf05svDbIW7qrHcym2YLf/dElCq/6xcCVkli4RKE5/JSG2iVel8uRKS3sMAu2+Kh4Y//
E5BZCmxYtJ5QCjnBQ+Q7ba8+05I9XCXpGe6nn51+LfFVEHwAXy5JFLYX5bvGc3I0r7IaMuSUI74r
CLG1MIhsV19ZPemDZip23IFgy9zhq8wBCJG+6uqh1noSSHUG/KeRzZX+7co4w+0ySAnt+G5Z/Y4h
CyB8E6pqOQIFp8Jne1Dvu7nHn4bK57BDUB3XvM2ps19cl31t/d3EQqJH9AokanmOHk6FmgoFCVEI
teN7eB9ERswgRvexsEnauZQluPzP8J2ylIwBnmfnBmxAnAzl0+N7486YXd7wERw5jtCrDo0avM0R
/Ri7amj4/je31m+namcCQakUQKDdJ6lChruToBS18/k6pWW+O5hMgewl6NxZDXhW6pVAFfhWQ9Hc
MUn3ZdJtubieXlBGgvo2bnGTcDPfHgLgn/oq6gEzD2cjY5MfKnxkD4P8mPwHPPHxqjEf4VvFTcxy
Q02m6qr0H/zJzzYwQgwOMKbnGClhF9HFYDSr0Jax+VBHIamm3VX7uQLZzdYaUNmTvsvkDalJ+HyN
hjLk7S2wN0latvI/jRkfqq/89wJsYzbWCz6r7IY2RC5EvOUclb/6MGPPA2mWxe/L4oQiFfyx6KqM
9C3JSuW3xtfawBVJCsT368CJD50YN6xTxj9WqWGhAG1GnDRpvGNX+8i2oZrITect4hfFE/aH68IQ
lG0YLlXdfdlC57FiW7IfecTOI3tJDP2ri2+p6OyIee2Gb4Qa2CJBXV+fmD5YoQK8sR0piOLU9ItK
CCac/hrRpLRL0Bqj5wnmXegVGBcnTECTT5eoyIrXBoA5Eym3Rgch5QFDV3c6WcycTnM1OQb7EO/V
dXmjZDZM8hFBO6gRAq7OhMkFZfbqc1ctRYbWs43PFv0gNaVNewbk8KCIh2u7qPtFnqda47TN+uuX
pmK80aF6YGZIunyjXuUQTug+nBd9jEP07NhyOSCVxyF3cv+YDUIHNHjVEWSvSUdqYRITpo7+Blcv
NTrgwtX0NlVbP/EXo0RwfV2UyALHDFOrbGmPGp59p+y83THjT3IUUSVqhRbNJARqMAkAEyw7vUti
7o8yr11Hh2TRTpxKV8gFfvnU1NHGRVw/osGe4eQnzVFz95+J4ZotQj/U5HKtndsMEuw+wc5fCCx3
dZzX0aZl60cKtddJjkmHliQQnBDxUB4X0KgaLlLxxwfhawGjJD8XIyeKRSGbtuQlMeumDRNx8dCq
jTXzQYRHesZp4kKT5aQL9rKs3wHCJcxe46c7l4YeUglLHX7/TezXEx0e1WJcXyctMVaSA6sme3v2
9WkpT8qz5z10CCqidPe5ByZSxnrDbOUYaHCTftzLGVirWOuTfOMhluGJ4hCj7uJC3MSu2fX5aFSo
2riVRBTptRejt2QYD2jiiZ1qAoZXJKVNikaKOcbKH+bWfYpEQl8LaCndloLOxUxBJz9f44CJl5sd
1Cij6QelOka2v0lRQuDQmQ8jTiuQHcrn28c9dRYtD0Y/P/zojGrnmei78erpvRz2fHTuGkfvIzfR
S+5rabMUktXoT/fW340DM7/edAoe5WBWBvpwe8mPAFr7Xw2iuJvegUz/uDJYIU+UhQwW5n1luObJ
QL8BEp7wJg8TxjG2ZrJeMyTNxFcVWvAc58XZ+9+DAJQgGzqI5vtmyb6hpBVIzan+f8Ic7MXb1w8A
jcZwUoBg8LOQD5iWkO+xfqgrww+ju5JJuAK0Oo3UmHeWpuuFIaCQqgnuYwaGN4BM3Gdrjxbfq5Kz
33hjv8y30UMcIK05AYWRSlfDZKMy/YaaVpeKwzlxxinmnD+20Vc5fcbUiSlhKg9kafUdUY+qWUp3
tJhkE9y4zQ7JPu6O+KLSV1BaU9RKvMyMzgf3hNMdGkiLytGtE1MM/hjumoDFofoJ9YPOOkpTNqtA
/2GVev4j9b265Qk6QVQTNqkdojpl0Y1vQcrmq36NbFZSntBPeBUaRk9engnH5jKJvgYKV6NKf8+v
5az1UaJc/i7kenZ63emikZgP7I874tg7EOXLJT/a2uDEnWZ0EGnsAaEQraDn8+kyzQymi6NcPo69
2EyKVJEWPXGECjxXxY6MMHrCIXoRRgetbh3vc/bvOLlMxyGvBbxSD0KcbySzHyrdSjNO+paNxgLB
KEe7rC7mr4OSbuZv+OUzdEIY8WTG3WTKj0+gh3fbN6Op6iMXwe3dtxxHPBWDOVcmv8WQxlPQJOkN
a0mEioD+YHX24XYAeEuxmpTuVI3sXw2N1LFRUrG2Jeyer0eJsS1K4ZiqKzqcOt+VKLd2iXA+DRRN
evKh8ZmKeJDENk005Qrzhx8IXp1dquzU0FRThZHor6Bizjh3jAxdOjhTE9ubcq/bu1yq61ptRCiF
4HmKbHwSoxdlPmAVwIzoIMLf2/gP0XnXd2Khhmanma0kWmfx+Vsu+sJ/WJTnrSAWKdQJQmiNRnpP
Pwb22CTpq7fjwo6qP142oEeudmksKilOcMp2Vlapq5oBjRq8wXUXoJXgMalx4peb81sbpQfR3ZVZ
fVn5Q7doP2xfH3TYAawFKagAu0P0izWrxPsTJDr98FXuPRKRFWrHZ2sKg/tPkflpXEKGuEB/kU9W
yC7XUS4seFsqu+eySqfRK4B3AbwApyRvz7c6c9IO/lNE5sMM7xDkWonmjPCoRk6kllQBwZ6NDfUN
TsPiyhOplCaHMylSgkknTd5ulsV99dss3Y28f+zbWCRbYhJqau2ZnpZDBKUemXqukiZTidAZACkp
7EImJZ8AG1gWdwr24dTfNEOfwo9ogpVcf88Q0DkDxh8uY6WA54xgo2CPLS1s+XWxFZbGkVbyIC3q
6kMpyZEhm5dgbGhrImxnOaYr7zzYbmmBlHQoZwcYN/B3Z8rrY+O7aNqsy/+QC3YZLmp/4pHN3mou
pTCgV+zzi2NgfIKpkHeTVaRY7g4koPjFdZvCklpXAGFNz4osfLosTC5QSE5gqb6ykHbyASf2eAYH
DgDbPYCq3aGOiGcQgoajxo3dZ1NtgCWog4+QlphljSm8H1w7hdeNyhCAOIfZlBbRY9ITl1JG0VWG
MV6s6HWbXX+XbVbFAeidHsDdQDXuY46sKiZMI6Uj1GN4Sy3zA5pTjo68cmNS/uwN98hZn753FSzV
MD8eBkgMFZ8wUa58Pz1PvYZpQbHfm8PsjnXpi7WdO0WktfifZPykfM0kAuUNcPl7z3r2nwDJL9Yf
bhsNHiIQUuM875ajfHa0NfhbL5c8sIp5jg41p+jXcwz0p222pxTZnycK8D/PRM/aXIeNWbasvDEE
aExiEqDD+RNefMy4sqLvrvHVWLrOqmGr7AW1YTbv88oAjSuVLE+HLQ+APZRjsk6UcBtvUh3JkBbo
W13eMduoVEzQ2clOzRfQWRJQC4wZtXxUlCKaucMMJZdGVx7pMPFoZLWhavZKQkEwyVG5orARp0/+
wy+wyttxy5CY4tmPs5pQKv8N3KFKv36rbfXbCbM7iw0/0B9B7slRRITX1rLz505H/ANjVVSHbobz
zwNsa364UtLunmDSGE8CthQaZ6zHRBidJQ3mzKqHZXpfn3rUMDO4XOre6LLQ1nJYqO6tJ9qbiZqk
t2tGAKkMKX2sLLil+kfci9cJ8G9QIEqDROab8toS+PKV5QsuGs7pH9IXUJs7Vn4OZ6FnCACDlyQH
TxE3kUe63wWtUkC/sJxK6l9j/4qj2tN2DoDTyY8OktCt3p236aLNGcKPouiRHc5lfjEtDzlRm3ks
ynN3CCyWCohuCR24q9lSMhoerePZVYfqWLt3+YLyMOmYVkIaiyst9Hko6uEPvbWTAxO0tugHQOV1
Uf6JeEDvcrGACOkSP/spXOEivieIX1HzzOwNN+9TZWz+LI4++SxTxmKPcOVyTQTBOICPWqsbmHvK
dAtCqu9St3mnb+fYpvtbjgPzDR0c7kyb/HGQ/LC2yQHp7/+1Z/Xd6/zlmXDISKU1bBtzYk8UF4es
Z16cBpNfHWFbVfYxHBJ3XdXU7jlThpPOKTMsKBrjmJOc/YwyTN+nuWf2QMcnoRopZpJvcoOfFyHu
rxeTcQm4YdqptfgZBmEEtuk9qoatcOdYkDChB1xq/qoc3+RYUEuX+zJV9AIhYuqp6mUWFZqiGytZ
rgOwn4ceo96VsRDA7nb9+CBpTtuclOoEbOOR2tPy4flBwoqq/ACA+Gt0EoOoUlaaE3qwoJf594Lx
/S7nqNYxwfKlRE6CBgp0n8/YsHQ2CYBM5vUUVO9M99P08x+tZSNr/g0G+jF9mji/1mmM/pAgeBiF
xz1BDdQgQKhxnlfeZdfE5sfSDwjdHcs4JH6tkn1PPm//IaLH1pcKXcKEuG89EbnS/zivXplPO/Pi
NtoqS6ZU48pntz1kwbSyDVgyqUbSoIuZax6Hvmv/qJ2i4GyFbZIa38sVosyyuXXNGyoos48HziX/
JPZJrfrclxh0ozg+jUukZm/OWnSfHEc05BB1EDSgC9+zr1RMXZI6K2JuL/0aQ3E0kQqgV8RFGi7t
KixIl/Eraz4vJ59M6joNK/o6OOD6ljyKcSv6MkpVArZj3YWYWGj5KW2ggfV5TvE9hOXZOkc+u4WY
DRxzZo04Niiv0CQX2FibyctZ2QrUbKIS2Q7CikdcJ0j7bof+fukvwZBdpFtzXRCg/OJUKNWSOP/X
7PHti0DQvoCgzWeuPnc1vfrqr7QZm2BUq+WgMlLHKnsSc8ELR1UmPgVPmykEs7o7AxHnojvUapXl
NBL5R3yH+5e2uzX8CNT2RuAAHd7QVukLa1CnrY7oZ28VwwE3zlYXaN3ba9Uj63kUPly/XhJC61YN
1veU/+PyC5duXia0GpEr1Og6HXCWTGfdkzk+Y/+DTnzn7wYbpy/IVhpztwLE0s6cCyVczqJl0mep
PHwSCwUtd47ZuTzHUFKMV/m0CgLvnwnLOxmHQb/hF6d/4JqGT/VwMauvXKTFcUfVfCDVVMH2ASgi
yh+8PVl5bBC8bawk5AzQJ7kejTpDwvIA5DY9vxAazkENVrdZ6e5sb7BKoJOWGeLvaz4J9d5/ROFV
O6tVRzA0nPaZk3J86srzFHa28QAqHh8A3NdLuHQ/KfWaIS2uSsv2lCOBnSZJjlDMtUNoFwKsdanV
XnS4Il+ZPY/YVOYqQYpVF/DMhcNbMGbMgD8VDiDmzPr+PGp+y7OioY0L0y4K5dEv6zrGCFGuB617
ijX/LMU1y/2GqLv0yyduB6zuixHG/pKIjyZpRviPLmpw9psMAd4bzp/tx7P7sfVczDPYzd8wWMXO
V9ZHeyhR82vb9hlMDiHwSzeb1PQ2g1iX7mW1KCEggJBEh2DszO6b+D7sibi4MyLD1cd2dRtmf+sT
foGw/NFVDJyA1rbqiPvNM7N+yUhcXD13jD3vj4QaG9zjy0ua9O+t2Wb431gTaulxPFRYoZCSChLI
PXq+CBmq2PWMe47W6ZGG1NTP9JSWyPftAvbRHf5EWzGT2Crp0SlMaqB8SkHiSQ15Yxecu5mvPZ7c
QORNUEfPe+fTICqxTE+P0e8DsjxubQKPJHzSr57Ahz2cI6+NzMipIdEShm2Y/O8lZErbzYp3c3ho
r+4/+RufCdesPpqPn061CHYfB3om5FV1FZU/z+me4TOAUIBuBYcMvGzdzaUsXpNihyYHSKW24748
FdjM7Dlkib6HJ83dxOgukrfTPCSSwCsJRKsmul8gsxdPwSdJWocOpZRzhbJgoL5yI82fGvVK4TgU
9BpiPOMBAE/F1mOtR838cvWUL+VEEZJ6Yisb0fUf4/WZunNNssXtU7C3SVoPTkjG9jTo/61CessZ
AzmfyzYBNFkKH5AfkW0kKJKGqsll+g5tJCmIGsI6prdAT6FVvluYyWkEID2WaX+zCBW8Hx9N2e2M
rZuJcF3FsbeMrtCZNdm5gar/wR0w53bOf4tEQCwygOw8NedZJ+BZIfTRdfF5ZezP9DMjU6OkpEVg
QC/+/KG8H9oJ2xnBc+HqrN33NNJTh7zRiEwQpETfDoEohg3e1TvBFGNTcUYuSY0ShDEzX9NBWjcF
YPkypT4hN80ss/EEj4fXh+Crw9LVu+VNvXi0h8DrRreVquunKEbZYCdPRFxo5jXY1owN81P6Ky03
in69uOrEs5LOXMo1V2QodY8BtNRAQfbgLF0uf/oNVYEsb3Lf19Fn+AZEQDCxxg+4dcnbHBbD7Eam
8NsN7ABBPnqOEvePywnjS3kSm2EsyzvH00XIvU6HDGQnX/KaJSUMx4vIHEYN6K7Lm3NtUQYZqPlT
BelhI56PCYKT8GJjwjiVew/cjZgGhCYbGiNsK3obGYgVDz0iwMhn/56xrjRxZJU2xbMDHTcGlFld
IixR1/OvwhkFUlQCSCBoGrt9A8S2JPG79v3Ux9vC5s+JlSBpqjr4T6l9M4DCi5+U0ma2EBzfKFSo
tLlS6LhAtOmdKE0JGxN6wKsitGSeW92a1Vig5wHwZ0TzHb1zaw058bG6g9HjVB0H+odph9mMd35T
0ewllFJJaXWoHRR+6OmALbq5B2iZcI8ZqA5kQQbTUykEHISJhk84JkK4TIZ4HLsTNXgzPNfMx6b5
QXY4auQ1ekTJ7DcJ86JyfxCrW3kNZThqyfqu6dr0f+gdW2vVsv+F1j+pEWGlZQscZMMoPtB2D4oy
4YgACmMPq/CgaGoM+wuZl7zUq1lAT/yCP6RvsN7RZvf5XiGgPg06IlOaWr+mRPsV8uHV6sxQcLby
V4CQshWRcs5iYT4+YA7tSROGbQ5EW4CLlAJuKYk1wZnYVHCGtRShMqcuszsg1DRzRskEKppfKCCl
tkb1yIxnW5r4v00amQisAo0DzPzTXNuOIlQkGPRr1Ln974zzLzLW+JvsMXBSbhhg4PhQeVq2FM3H
pv2h1tUiXX39P0bGklvBzbOilYHa8e2tFQ1Wm0fveAHh3qzlJfw+EHNXv8hxu6O9Jire96gMxPZ3
8cz4XLK9YC0p5ofpmHkQ9+gZux2ZpYNynvNu9h17zKKO/M5oU4/tnfRkh4uS9uE+My+T9cHN10JS
iVlpGV/jFbACIPG7+xPY9f0uPKEoz+WGE5UrIG1HwcXmDU5oJwxmzGiLrHEAnSL+XmIyo6eaWkvt
c++iqojlLgQW5Txj0beodFdRbqgA3H8XhcXVME/Wp4FM/lI4J3Hm5CHVqtgxy+n78s+2qBhQ1XTa
XnguuUbMDB4lmdEFtyIH78wKve4EqvX6K/Mu5DwY+xL1y27jKdrywKMDZQrDym9QjpsxaT7x+pek
zNDvrNsXeMpvFcG6MDF21Tr+UUwX5KB8dmqwwzrw58L01KCqwX21E+nZDE8ZYqC8OO45MlBGc1CT
dVz7xd2bJYI8AmPvGst67Mq4TtSsdyfZeD5oFWO53B0MOuOnerW76LKosXgBCKT5u9l6ADMt0WQv
cy5pkXlnarGGOhN104wY1rEhv0qYBR8wPsfe9y/ZjaW2luhJqLX4f0JYEoJy1rFXV+M4uhFH3K3l
M9WnoPyXIVU7FAGtjOSfSIurmF87ZIc2O/VouGkBrzNg9Wa0Rf6+oEO7oQj9EflIfCVTlyr3cTP8
i1q0hUgZmL3VWhaxoMQEzy9HWs1t4Ek/DSqdS5HMh9PASenu6YUs4NS21Y/JkNqmkg9VD9ng71/J
3Otv5ZT/o8xSssO7NJT5JoOUkLA8dwxI7u5x2xVtdVPnTgZP3xsmM0OCyk9qhqZ5iuZos616xIcR
xOaLaKIuBI6SZKQJApMjSHjA2p6mr5p8i9iJcnVKuM8b3JGKC+fS/8LQoBRCv/FmITcbuFA52yps
VkL6Dmx2UlsdHsMJbBn1DE0CRS2e7a9W9Ci+Pbi4Zobox9lXE8rGnd8XQ+5wwyexaUfRaA8lopWc
ThOx09KXl/beIMBGT5fLaGw2OjYlWW043LwSxaphxG49VaeiESUw4MbwOSIAitNJFP44eSGdMQJ1
TSEjZuCTVwGFa1vEAxMQRXzegJKoJpv4hWAKcxHPm36MTyme42nD8lzFIQQip3aTTt+jxODkrol/
5MTNjvnsUuXtfekaYYQoiLjx5wnYx1+eCKQYONRRBWVThPBQyXo+2YmpgdSYu2F5cbPOizbV0zMC
ZH/1FGqsbpjoFfkafENOjYiZl9cvLm3gR0ib+46l8V8p5a1iO8zmz1rkAmlTrLegCV+WuDtregSS
+q+XBFBpo+cv5Y/ooFe9liojOJxRCiXhKAMyoKtxwdj/sXzc3XjS1yO8IXMd+kmfQRN53zgdC7td
5u96QWYIJ6tyWRf6lB7nSXebEGckVyXsXSf7l7S31vMJIEVFbMiEdoN2go2lfnS23NiVgn3k3Vxf
CRjS7nrS24onJABMMqLIKBl/r/WFmIdTTTebUa/mrer8zdEblUkaIXXvqjVGSV0C59nchLVlC6qj
m0kJz3xnhcpi/WKd1Pareg+lYDn4hNKepCvHtPZvKWoQ3g3JePpyKMoCkXnJIe8UNIKBUK3kTdva
Tz/pMfVLyY63Djsup9OEXGWhn3h/UD8VhoPCcEaHDwBONP4MID6Q6gtQLVNdpQFTIyPvw9IvZQr9
r28Rt4x3aT/S6NMfTVWU+weNKdj4E9xX/oBJRPcTTCKIuItsZLa/PZwd3cw1TUwccFYfrbSD2VRo
pcAQLIRpTjidDxTQZfDuQypcit7ERWDoQJaqP6retOW4iNngYKEBCYFC3qYtcKOdEVV2plyGK4xR
Rs1Vln5FlCefR+g1H6K0umFBF3IQzZL6jIRRyjhcthPsTyHxAiABBoyfqafi65XInuZDMfg6YKcH
y0GnV2yslk6McC4yTloSOJFjDPtkoobcVsCR5Ux+b6J9vNmxc/fhS5/dvbfCqHsIID2/9Z+VDNJA
cnmFyjli7XAfZBCcsmOGPPp18r77ZRYIErGIkuZs5LI+ekGL19a4vcoPsIsfGEXXhv8ZW4S/yBJ5
cUvZPvIbyo9MLG6bvOcFoHxWPJbBdjXD9gAzpuVl7je3leM+EyI5rA/QsgFmHPeh6kbmIU588qTd
g9CVDoaQR5yxTL3e8Ui2SfHDZhSvEGfsArCLzNf6sZPW1NxIhJwqzM//1vEb7PU/7ylEWDPJ+M0H
mlN0VJXCJYDaIirkhlNzNNwvaY1tj0eUjOmiKT4aG/R5w+2T8oPask8N2+zJCCG+2xzTDTBD/iSm
b/qo6d3uQKxutPB638KEHZkbLpgNfUQAasFOLvPAjsALyjNRpH9UmqBHBw84ZTEolijd79n/yjhG
+B+s/DG7H6+BPTs/9zqTFC5B2xBEcUZeWphn93Nqi6aKkzD4yTFIW27g6RO7z2OtXrdKcAMIh/ly
VK++CZRIODhtCBq3D5n/z97qrts0KJHzsGePgIDobBSBdJUgqfyZNZEZq7DMkl6T8A402fedWQVC
WPmmZR19rT1wx9MNDlmUhPjn276pxLuf2g4sPaX+ydyps/ZjvSSPfgV+aErA3WKuJs5B9bc2vjD1
HZr2C4XE2nYMruECWtvRQddpfq4nJZBghqhm14eteTDZjw2C8vUmR0ZUx5maPO5J8+26sAEC4LUY
Cfb/VJldAUk2kYFfVj0i4eKg8+h+xTb6+q8jkvxsvgWZ6PnjCwnSRm7y+k2pYpgJHoBhnEb2wPpZ
Iax8u1AzK5BSPTo6+sgVTFUrSKFYlIFnojpuMrt3fVUD+f9c0otW2UZMTa+UB7R2AN2hbYNads1W
uDooWVycQYI7oJV9AvmaLNf3jGnJ85s+Rcoc5O1ZxRPn9AgHV7QnUzh3Uc3vt5zhkp6fA/fix+1+
Dckip7gC+dB7Q4IWEJ21dXtFQTzpYssrZ9lJb+Pn42SK3TKrZPocMgf7OBuv42GQOpUoJ+M+2bWD
1OYjVPpurqgSg126r9RsGwmflU8rNmJXZnyfODrGjQr/meDPqE1RR1378li30iJS9gjQTquyTj/Z
fEhhWAMXQF65I35VWF5TRH8+4EAOhYbf09hdChCWJS3gMGr2RjPKagb8U9+oIK0QlC8o9u2cY5x/
3xqppfxpdBZa0UoAkm8xK8QlNTPgUzpmO/dfgGaK19gcntGrYBYfs63qdMahmq7X3xRnQzsbK41H
ZUXWgk19cHAsrG+tHqLLCQhvT8Z864wbT7jRhSNpy4aKMtouhfx9MiM/T0UDUNMRk4gsDs+5Quvq
kz/nUAQIp5eMmfoKlEFrwyT4QK+8rm4U45OZSlVdDc/mMwlb2cCCZNt/9WtPpWtKYGqshaEYFSv1
3Fc9v9d5R5ZJFMbSbNNbEm0VOHKNMbxutdU0SjtShWAO49FXXMdklc04fUBGJAOSvPltlJoyxw0E
KnJtH5Atpy3cHL1oRkOeh9ofr1MYLN2yPeA+zoww1/MtETpGgIoWM6zYKFarRjEhTF75P6yoGPhn
/Lb75+QG19hnfZfofDwFp2iMVgDYeBpg7KcDYKxqM3tXNQK/8eyFyj//Br7zIJ5pCj6694x2n7uq
XSgCsDyuX7uO5ObyDf5EpXN7DwLPlVv1R8gxT5wxjN+o7pbBzimB85zDWShIKg6WPvkp12jHBQ0R
5uaZ/aOKpBeaTFbCTFfafRVh2SHocOLOV6L+8wUOeq7vJvbeON1N9nrpQCgq0zuzJHcvj02e+12u
DnTTCKJdN0zqM3vHCYVGjpyqk86c6TbKkT3XEy/9f8LN7g4eeCziFoZKUwF3GemFKaM2gomL9bxz
hO5W801cAysLYr7HXeA2yObUdNnm1Nudt0heCZvS7wIkFps5o3YPvwpyEUIFNQLzhgvYJ3QKm42u
gxOZUhufhWmbd92q2jLLMWww8UFXaQ9gCrSpGsF7ntb5lZoknVWSnrJChLqHYdcjoCY7vkb/M+hM
KiBKdyrAVQMA2hIA0A5cc7Y1tdbLvvfltsVQHyIIqfT0eEGCTUi1pbwDQQMwXf1Sz5GtF4/n7Uuw
ANp0x1HgWyCMAPns5JN3Vy/dsrtqvXEXQlOyaPDAfjGMqMr2P65EB2adrxyo8EKDleK5vsJK8oVO
BXvfpO6kGgmxCGO2btH5Efwr9R/QiyDBT94ykYfdRJwAoyFdnuZqPWG9ubDGGKd9BH9NB/Hrpgzm
ANvEET/jXxm8NPX037sNFMVGkNDlL+FRpgQjyLAXOXbdgF47YyiqvhyVFwc4n5FizQSwp/bZx7jk
a3Jnu6dqdIjqk51K4++vP9VK9VDxZqsZiX7+7lsGByx9nJhBgGb187gzqqZ27oevUU2Nu1ngvvvq
Tj3ltCgEpgpistOiZP5hq2VrTcHZrnkoVdg7hX5G2I5yapMMBWL99YlmoWNhiUvaEZ2dlw3oDq1F
8m8Qvd3YY4/hrR+faWtjmoHOh4/SVXP9hY5FDAjWaFQymjB8+10DSDxRTob0nXNkhgai4aGtwV6U
2Ao/K2cqGGdZchkTKk/Pmhtc9DdcgtCJt64u1dqUgsSS+9SLSXvR2vLur8pOcWzvYQEFN3drPKgh
u1+/+9O4B/8NEzDyyZmPpalhfkjOLUjfz8XDBFUm8n43ZZiQAIrRWDvzGMttCp0SCCe2aasMXXof
fVMQnjWzfCpdwVsZ+kER8Auffs4Ix7Plw3Yif0zkzufCT//F/3wEo7URHeE+UK7R8d/GPg1894zI
70HkGqSczF0Hjy6BcHz+P0Kb+XcRfTHsMgG/sddNe/Hj7FdxnSmMfnxMoSzplkk47pWf/a4YDsPH
n0jEPmUXZWjOOuB1OWsMtg9sMSE06yvQxucWAQreOwr3lzZ2PrmCszdnunChy4rW8GLs4FI6m6/1
ORvuLXC+zmrdxC1QNnJm4SOz8bDXSRb5uCUu6ONhAeq8qZZX5cHKYBq5Gy9RQmAI0scdXwHd5pIe
LCb2vRkcv7mvvp7jHYjGLl0bHnVq55097iwO8beWGzUy46sJgIDE5YIzgWEMIFR79ot0z+8OFC1F
yPqGmnBU0qbd/U8AsrE/ys0VIN+iJnZaeLygelHZBbxFAsG8nNvoh8KD4XR0RdGp3xRdVgKGX4Yj
2HcCHHVDZwJWXkTbFIEFr5pJpdToV6cBIlw7BnM9UNqkpoxhirU1d6qP4vDO4iwPMJO1d0A4xHjl
benjxD+9mV23VjvpwMKPW4Gxqfy/kbKiWsXauNI6I5EVGwbGlKFcg7T+xy2HPMR1jzjkjDLfIUZ2
/ymBQ/PoXkshQeHrkDaqWzLUI0CgDHJ0kun/h5+GwTiQW8Krk+gA9c0HFUt6RwgxbETAjazrB3nG
92GsUmjkmm6cvWnBa6nZPcZYbCd0cGfKoenD6hMeqLYgNwHe9AEDihn3q5uOdXgYSM6d784UuMiH
4oJQpTpW8wiD2xiRPOfY/puOzF3y99hDoA2pVLw1KYXyIOZr3y5gXSUjnK91kHvm2JZPrD4UTv5Y
tloEl37E513wtTRo53Qp+GzByLSNLrnmz34xlBzB4vi+BCMCmEDHYI14TX/xOMyu7Lze37lYmZs9
7IyKXrOpwxWt+5HPTnDAscuTExCPAaxQ5PD8rFi/0e1Tm2Ojk0MLZkZ9vHdGFuW3wmsoLNk0IiG4
M36gM43mFZzWh9EXAdBV1JBS8AB9rg6rsOshpDIpfyJQmCjdCOWbX6TKl3ag0KHHXDkoYqBisoWp
C2Sq5tUhOJ9dm0mnQ+KkZo5l3/OZOzf2J5uzmxJhoXwia9cSI94mU9c6EExsfS8RFHJC7wvVgBbm
eER3/SXFg+h/PXCC4MxfzRti4xqcgbBFg9tsDiyVwg4wF+0UB97B/9/OLgJ/GDU1O25k7Ijn3dc6
0Btf6A4ysESYLQ9pemrtzum1z/v+PSGiHGuicPbtUf34LO4KVIh7hZAZuC7tWN6zs/tL343msuz4
EhgR3/g2r/LuEDj2FrOyx4mxeDZDOAJIDENANqKBsxbaphh2Il46Mp1Y2t+vf9mD0jnSyZpVtV6q
hxibv/u/J4cUKvMRXkmSnqbR0g3FMvsmL7KSIk+/4Vb7STkE97i6vyjGZ+iNDvVXpRThj7cKPqdc
AL3blJZa/zqTyj8oV8ttQplZb6JPgw7/oR72HXm0H/HdU6s6ibO6/CAGfVut6bBmT0EDaxVpG06V
5eHE9qXxj0zJSw+TCEOXRXtWWvKmWVvptWSv0a7jOUUiEzjzN3kaQ5KoHHieBnG33FQ5Ep1eaxrG
uPZwEOXdIpPKVShCGjZ4ie8cJx3ewXvt7S8lsc6dLLSU6y9GjYhEkUKLAms8QZrzyP9W3BSbeb33
WnbbDXylEayAdXhkNEqChpxvD9WjsnwxFbG3Qfx9viLUUT7Ra5QAF8UlWSOByky5bNzVvcs+zlUb
ITGUYM5+T/Bv/MIzKMFjFFXIuI5ux5JPxYmThExydoHZbfSNS09ROPFZuj7kDy4hfiHlKsfU9m/C
wm+/XX4hYlMh8FZk7VeiiqpyJIutyFmc91JM4RGU0hMKnsoPwg4gI6jUbgBBppjtQ7mVQbxYDLFv
SsX0F+llLHRGEuNgB0iHHSEFONf7+AdapuMEw2VPYb5Rj8/oPz0mbbuKr94IUtbBO2DMAjC1hRzd
/66vMBXJCsU8emc9xwRn4VnaAUyKXCKlsE0kSZyHv5gaTZvvh45Q2ZTDdNO/MWGaw7gjebAxOz6w
Bm1SVIV6Jxcz6GqHuxXTVwgZpuqHWKOumprq6ingRexCrhmRwZKt+I/3hPyGevjaagaCmFXvdcdY
P7Kxzzm83FxN7s8GBrRV4U73u6yGtta02lBm9ncDQQEe2ljoeyB+bYL1HIgY1147HcJxj1x/PcgV
jvsn3054IOE6mv7XSD9Y2BBCR060zUXiyq3VnYaMZRiEcgTxaJzGjQFlL5YPp+hj9BE0ai9l8v9K
/r9GVR1JpByNmK1ZCAb29M8gj87XWPs05VcwOdHFgKOzcIkrwp0dt9223EQoxJJnLraAv9/lvv+N
MzTYvsPNrutQgnypnruq3o8wRyMP5ztWGtgISZ+sUn2PuZlao4zbgiIseFQ1sIKYo7+Wy6zJ8g36
yOywxJNRX0YQ6y9cpxOxgIYLWtDzUn4alkv2upwy0rCzIdh5zlqs5UrLVor3sHVSetT4Yv+cldSp
Vm45Pv4ppLIXEp7/zpsT/UP3qb8VGcE4tz78cWBaC2bQJBQPSAHntaKxwDy4s79CYDxj9vHoFET6
509jx5IytPjpu3WLYhvgqx6tflgoUtSJZJDpjJc1F1TN+7iSgHK3vS/OVc5w/5h7LrlLeNwYAUtL
9SmzOnIfFEhYcbcbLvvNoJ9FK22XrEjef5z5o1xb1yvc4Kx3i6x/X2zJYffnhzA/7TMEJImhLhK6
N2KBScLQpBWTYBEp0I0feeNOztl+jEA3Y66ZILYKxDtN3PmN2SkPdXciNGHlK8Qbc2csBLQMvNW5
ntQhl8QPOv7MZxq9sUDoUcmFDM2HiyT4p+ZMOiZa5FQ7S/hpdo6J0TVOgbxhuelY22DvU0CD8/Kv
mm60UtO71b+jIzDl5gBcfDvNLWdRsJoK5Bf9vN/nx9VpQJQvQg59Qg8/sJB+m0i531aAW6nFPp77
wgqYBJh9Zi98wPfOUgUnEz/cJFTdGEvW2IXWKExED/NspihN9FxGFdRir8HlojFj2a7NR0G30GXh
Khw4z+NNY22cmgd4neusdq0FnVn4ufFpOqpTYAdgF09+gJ1ukY9YsRuSNQDVetUVel/Ocx8oxF+D
s+2lOobGNlXAFhYJyNgxbA9L8+8CumiJAlgdrlZyR6hC9WbMHXA3H3385CL+RsWnuyQ4JdR0+rKq
ibsTLoe1IpNkeMcb/dZWHdy5Wo6lpgALHKAmCJOHhckIEGPhs/CCVhp6q25rBESSnhdZj/lw2uAm
CtjE5Xzbd4EB9/ARWSsU+IAKnhpDGqOyOLsD9G+TOF0B4h2RPJoHXNMfnVHi2dlWdi6bedw/Q52d
9JYCJukdGcH2muJRg0KtkEttYyJpC2kcINj+lv5+pHCYAUuETDZrxE/DuS2ySPNpnBX1ectCyZai
ETN35yTZShhduQ22bA2VjXz4cy0cMmiRyoOeYuAY3GQ4lPSwMrTGWaqz/j/5WceR0nqgeXAAajqX
GIRqSpxGqzW+LarBFnNKij6Fc/mqGASpIZgunU7cYfIbaVaFExF7dQurzVbXQ2+mHEkwHf82NvMw
sNTvKzQqoyeBZbRLbMGn3IMAUUM1OfYqsLv8i93L7/eTZqu5Fyu0ee4VWPQuiaL334uqF9KBjEc1
GKRwonFj9LBx3J5QUivJGWp1ipRK0JnIn10q3zBiEWTi1yqbkKIlVWg5cj/VQAyZqGgCbwV8Up81
ra4FmLeZb6LeUBz3klS3qGSCQJxMpNiBiFn2lLbVwxIXPD/wMR2vLT49lQ1BQBThJfs29qYkXCDu
C0EQb2oAItku4OOtRo5MwH4c88SOHsumjqVh3E91T6ZEal0SCtapxrEQLjh4z38HK0bkpgI/ldHU
f8uMT0SqR76EELikxTwV16yAIfzMLsVuPWi171Mbtb8ML5ZxPvFP/US6NSSOkVgIpL2JSLZRA4Mw
8mpudZqQptO5OAgPYLmfoO52brwHSRk86UXDJPmdFqFRExw6SGNu0aycUGYLIJ1UH19S7mu3HosM
Gj4oyIMiyZTZ2qJL9nSlaBGw3NwzCOkFv2SyE9cO4iQ7TmmUtnNcuNSFuOQAgTSAXoRHsWVzumhv
fRmlfBzw2nq4V4qFyyxWqPBe6y6Q5XcoZj6MjeI5JaQE+w1FEcutYDLyCspgDkTcOeedaKuVqTek
U2+SPl6IJXLZCtlJmw5jptWcF/BUGW95IsDJ/b8QkVSsiGxoaem2jGa2YNqY7a9fY+GXt/fZxviB
bxmKB6yYWDB6Pxn5TdnyJD1exiQoO9URyYUTlG3E4sNPZGUlGfvw6YPVbbv/9KZlRgyqzBA3iNjs
nGrhCuUKSOLzehTJbq3Vo9azRM6xBMW5qvn1/EKfMbiKh6fwmUIY943L2LM8htO6NP7IN7vviBW5
CR/Bpy7DU5YKL+1m7GTktQi3D9ODSh455dpXDoIs33Usx4j+4PTaJdMSDEPHIq5KjHCLn9G5Ka8c
2lolqiA5J2tlGE3fFu+wKBKMCN++oblqY5MBnf8NDyilHsHvVIAUv06F8klgT0HbMXniAJee9RDn
bsetcgNuvN8v3Q+CppskppR+aZ8/Tix/fFa3ABrO6TeOBTU+cJ7fJdn10b+PFcPEpYLUDMQeZLbE
8uJG0p3N4bBYEnYDQbpGOf5iHg4rTHPB1qfp9nErnF+zfFQkKGMUZSVAVc4Inij0g67Pr8OjT6vn
j/aC+QxPcvy10l2+2C5do+LdY+Z6BW7HwkfN6vewedQWzySkcsjIQjfO52jjKX+LvW7xfA+AZrBV
RrgkzCGYwWRyr1GjziHZrtWk/HdkvbdQ8kN6JChkUwutLYPXld7yDmsIhUEALz+NWyTRtRQOluEm
Sy6g1L/BQuAJNRbON+sUyR+u/4czdc0cHrSemTenk4kwrc3Tz6lOnzXD/YaSSCpCOh/WHXlyLZzz
IC67f8hBqURrsKAG+2usLc4jqecJfnZn43Nfo/Zbr1gfSv2+DPD/rHvJJglk2ZPjCCsFH1dMLyLG
bHleglxsrzJdPg9/5gjCyHyIGazgFs/87KI1DMSk5BvMznSVGPCX6U/Ed3hHobArWMUbFnN24NYr
HCZKVLzAZnIIhZYuhwUgayk6sGZVgma63+K4NOhrQ5TrLMogAB+t0/czCT0iclUpQiWwvNcIXjP4
KZ1RT/1W+4YhNMF0slNFQdJGk/AXPLqg6UtjXwNDX0io+bhqajQQbokHb0PrU2UjF7nH+8GK53T5
gCSnH32EBFR6esOlsZN1NagzSSK7OkQ1gbAdsNzRRuXEZvBZeXap1vqfMwLG+/aepqJIo1oB78RT
P5oy5vHqdDxBmTTIXpAmTMbacrTLymDTipY5o0yRhjLhttT1BLCLdXMEroM4wUjER82oiaSvl0AZ
RuOjmD+eG0BtdeksyncZXu8rmx51R9vKBWfPVTExsdkwVQTEKX/sDD3F8Yy871ggyhTl8/8t2RH5
tharyY0pZTr1mkWX19+gMtLDs6SBXJSbPhACFGyiO+YydOYwhfJjDPDaehyK1J525LjgAhKtVy3w
M6KWDvmeUQm1k2WtKbTKhScupdKQO8EVDXEhopWLs2SsDQU/Cy+UaCJsF4fQZKUvvAIMUD2YEj5z
qkG4c/4x6ZsK+MwFK3tUhWTfNRN6RZmgITNS5yL9mtqsWM/8kYLS3FxuNufI9fES8cNssdkhxbfS
E9sTkqYQNoxqx7SbmiRAL/VSKW4dU9hIV9ea3SFMceMC86mq6lLZwMzbF3w6ufAfJV1U1ONO93mu
3olaFc+tB2B+Z267rmbvKoUN/S9/fxjBCFWEQddlm48GV11y1aVfRkP3Gw8qQ5LALFEGsV5iVPOB
ppmWwKIEueD/SuyUn+tK8P94DbN6E3amazd0KijH4iuiaFe4WKaKyR5vbf+xwgx4S3io0hFZnYad
n0/JAMvoTngzHNotuiaaIScSAxiXCe1REzFRsu0/i4qZZsxDygyjaKhSUYijn4pMuqBjB8+3C119
T5/a1n5K9N1zQZST5tbv6F3Xm6iP8ZEVD2SXE0tDevF1M5k2LpfaPjq5bWkuwTyBD+sC8iIihc6e
/D8sNt+Ri5gkSaLJWoT66sL0A/m/nF452PfKjMn9PDF2mYlI47q4h8DDybK39gkFeA/BNMUpVPI7
S+kzjVOshbK6uG1gAcxhEhlYGrFAPiMYNADPm9apQ1CaELRZGsNbwNDhpUA96X1JBZv/IWfEUye4
MfjS+6vfp7s//SB8hLrI5PTSwmsklqxeEicGh+53syGZ0y4wnMu2gqlb5JR8DjNGvZGAP4xWqk8z
p2DpozWp//2pfU6nUX818Y7CQkkT3YCbbtVwA232z9PwGoninciT5bNU5MQ2BS4rA7ZBSNRv1/M2
cv6yWGCzsiwExTvFFuu2aFTE5+E50kcj4v66b0EePisb8DVAkoQhB+vXw6RdXzOMxuHWwj3wJ7HI
+KwXrAyQVDwPkKRD9WrHhbIOrXWCwYSCsWj9oen4TaxVuQSEWw/uPmQ3a14yJvjOvrMYAzOOmO3b
W2+lDL0FlwJE8pteJit22r/C9jsAD/n9BYjWGulGb6l1m1apHmAh2J/JgnmXynIte8ZaOhT7KMv4
rnxP3I9tiNmv1Ez3ybRn04+TXtDYpz+Y3hLut4rKHowgK1veKKM0JxBckOTk+KyVfiakrKjScA6B
XHgsdCov+oGPaykTlJJ/8LCMhjon5Ib6DeNAaN3EpQ3Cvg8GzGMv4Lf7XFworZ0YdvT8pkscHkOn
wjEGt0DMnxAYBQOEfOaAR5VSyWCjIYfJw1tCC2OhAnhfqpNP08URQ3iV3a/6+6VeWcRFMffxMjIJ
cmdeQCjYCdgfHiDw0jNGFC/tm8gtVX3dwrR33shNF/73xNqWY1aQYivqBfc1naEZFScBo1u95C+V
LndHbmf4CmrvIWhEXkn41rLJqpc+PJpvtVRDoospo970wzsVLZz+/im3go5YkHpgVCXogE4H4jXT
N6ehpfuOQKphXHju7LLx4JvslP8c+z+Jw3lgh9LKwjAqLcbeFNYV915Beea8h6TX8+H5g2QZ7CFh
NXx8tRVhdJa7dFo97e3dSFX/pV24H43Ws4NFfykx/KlVTQBWpSQsAjXPWz0168exCGRIdUBLZy6F
uaQWBejl6nWRoip9sAcB2J2sVSEHJxuKdkQzLJnsdbUs9Ha5RuWxMw2tb7LntkGuriCA9KxHwWPd
ktf7waVRNxXwpzbfeVv/ZqGku52UGQo2ARdxjjxaAzJnWBdoz2Pa/SS6j+OMGUkVxxR4nDgKak5z
m9UWZij8stWCQzhXcQBM006I57g3hdXdGl/Hiet1vTl6toP4wdVwOktkxoP4qun0eYMcECEcf9X+
82wqH0tzdDFd9oPiGFsi8PVAoSPZYcWdT6Y2ZkaT6BCJb4Jve6GvAq2SHLlY+eOEtFd2YlAi+HEt
SwF0H9SQb3T0UxoGjmfgmSRwwcIYew11uOm+FF2Y9SL6Nf4y5WsYlWxkTfYPhpaVClpkG/r6uEsT
istEVDIAolrL/HT2dtkBoFq8jVZ/18n4nvXVXFi2/HCYpG8bfP98xIVtcEnhm1Z6MGAJE+oR19i8
FmdZ2Jw5UUcLuPh0oTkTCejMqyc52puAdgfV+vZ5ArXkz7rFutH0zmTogRXXdElbsm5JOGgSGlpM
HfM5rEXYGskdJft7eDPJQF+uTJGskv1fnKtG7pPxx3bVwTN5ewbfJr2WSXwh5kcuB8InHQIU5Q1O
hF7RSbX7Zq09Nyw17/VdbyaRF3HExECyULbE6BLUHxmbgpZzONP6s3E7hz9g7qaUFsNVjo6+e32O
AX4wdRzndGf4DJAcsjifKVWJck1La5Ee8a0DTrO8q5fQxFt81sBA5lMMiqOwnltpHZmwi3pUpTfE
wsZLN99p9TzNcnfP1TyspEc+oKWbJZTFSisskbluPgYsO89jvRtuEQDSz6TpD5AcQhWFR39BB/cA
ZUUqyiEVOJ9wHKGHQuFFnCjMJ17s20acCIZWndUUAKOIkh85UF3mgx963NhMhEeUt1XMwmGwAg8K
JhVf8PtsHXy9XJDVu2/OjEGoITmEEp5dpuAX75ouuyxhsnZ/NNkW2DHuI7IFye6MDgR+dI63Eho1
xhNnFH3QHMFh5uwS96WBvixcZri69ha2qHIlVQa9V6v7tHjuYNPVgZk/Nkl3yVbOKET+6M/nNOOf
nDix/nm4F3qgHpSWMuCRkoIm+SYmY7Wl+FYuIKbfOB/SZiX8EswFAcVb8o0qWRXKLbUBQ7cFXdFc
t7pWLNgQWnpKJ771026jlmbKUqBKVDDchxzIRAQuWlpTO2lH4EHepgjTPfee3YZvXZgOzEc30EN3
adqRsbaD9AGfALLMQ3i5lRlkVaJqlMPSAVIXFpHdGzpw4o6rH/WRgsYl5gx4vY8HcY9FW54xbtAk
/dvcavJmzETX+nlocvq0ywSu6DpV3jesbxyqsiQmoats7k/o5dhhBaqVf86Ie5lr+j63DxWu8d5m
iQ5Q7HbAHCFcpWkoZoe/jAMtgbRFgf1Pe9+uHGILCRSepB6p0TZMRNMt+iIkqhVqB0JUOp4twkCF
fC2iJYVTcbmP/kMbTjC89x0e7SHjTudl1B5+RiSW2+1Ebl7kzrZEvViUc2ELnRcihHTWL2Mf8mVf
PjCJKvVQs58tNDBD9ttMVcr/CvslsEHNDdMS7l8Lq1hjVICBozet7Dd8vIlo43JZeD8z1ggkrZFR
axz7MmzKmQj0yFJEWyRKVAA8ANlLTD6jDW1OuA8oNVO3PWGX6mZ70cxZRnAgoVeU2XAuiMVoEkRB
8/9d+b4I4Cf5HVJ54j7YGjPLp2p4U0/6Kct2IkljnpwqYdezm3Jdu4InXBs/CicNZSHwF8DMsGaB
f9AZzbABkDxMRvs9DveMHZvKXR01AYaN3puyLe3Rz2DuLhVYMGKqE1J0/PT3dfSE/Wd5Q7zRLz9T
2xLsC7b/dg2r4Gb8J8l7grt+hnrSN0gkkUKFcASfnWGneJIYLCJRFlT5rglksjRGHFXOKHEtYvwE
7xqThagBRT8+p3AUCQ4BKbGpPip9Lo/+XCHL+JmAQltFQBXfcNRTF/Phv/HPz32YiHFRcW+2UfcD
bjLtiBtwhRwoV0gLVh4l+Me0HHlQ6bUGro/s1B/ib4c0GZlxObx2qsWj9geIrJUjOaZ1yTQ2jX7R
d6rAKceu96ZJxtwoCqY8Hp5gM2B3fQP4B/ZHoeko/xky7FJDHmQCQv8hfaXhx9jb3axEL3zxM5oa
nwUlw0xStFUezwRhuSPE3NZ0WBnmsfLZScqElyeJvVeWjjZD7OOuW3VoIfnpdCV7ZAM4WK2jUQfX
D0aWCsVm48x13O7dDZlI36IH/TtKq99oYDr4keaET1O0ozC1i0MgnL3YqJjE9q9XkmXc+IlGqCHl
1UbIv+gdpS7vvuoIYG50GShuOY2U2eyOJsjjiLFdf8WjDFRfwbGezfJOyaxfJst/T9pJduaeAnFF
Rt2vfygbWB4GWCZqbzKzaaSpWdKbH1RWWEjE5A/0HDOfwobQpKHTRCJ1Q98uxugKICaF+poAGFP4
1kAhi0uWQ1Q8F9ke9gLXH5Y9SbdR/Ib+k7meQHqB6phAVVlPFAs6Cu9fraMRhtMqon+Tmem295in
8hPPcigVS4CzSCFZedsU5PovgtAnyI+WmCWtK5i7ZOR+ZwWLwC1aoV9m3wbn+RzbvbJ4uwvBOZso
SLJgxT9sdMolPim15KmWzEAXimpF2ayYc8MHMD/t93EoK45QcQ0sECrft8OvRYfCvtJ9rbZYzVI+
SfYyVIELW+4SwcASzO1Q6VholCjsHu/N9fNWIewHvmfLUSil5bnPDjKnHUyKNAMAAGIDkLW0WIV5
C0jI0l2p6fDBxAPKV9jbTtp+GUi4tI4uU4LpGHCO0NomvfTljPMe8y/jLPptD9TI7UVNeDRd+5YC
7WGLHsQZjMvCE41UdcfAyG/aEGRxbtXKnc+OOjKGm5WHwjiYhLk/YGrGkUCN88y8lNpAuX7oAza0
tlNx5NPesuu55kYZSHweZhfOL0ecOAhvx6joDqFhb5YRhHEs3fjqaOdqqOA4URvihnxLJRGhRHpR
cN0ANSr2zUgAMtRxU84G7oNEIXuGEOnygZ4U4wvzBWLXrNyITM2YYdKbQqSx76Ambvx/Vbgsyp3X
D5eRYqA0/qQCbZfThjS5GnEcr+ld4inzB+GG8zUpPT05+/J9M+EQBW6TgUzZV6nR5Kxb5KkG67vu
iUugR0XrX6e/5eiDe3ibw5077jq8/FNC4VejnmxqOZwZZ57LH+Px4wFgGUzl43UL/QprD4ITco6i
YGVcq5DTwzrDgePx1sufM8/P6tdAaeKT63roFT3uLQAvhAUNsc5cSQVJBsjEgL07g2yCoc5hzWxs
92/759bSEqAs9imRE2JtAjnh6IJ+KmVn0L0ofYOj3WE8Q44oqfgfyPTu93iHCG1qMDActJrBdR23
na6yCqeVeIVwa/UH81ue5A0KVPWgz4p90yH5OAnTUuFWbEyAlXBhfostTe7zgf0mfVZINpcpN/vi
QQeipBnb5azp+QMBGPhUJs/IFL7FIqNhDS8i0E1SOh5siMT7TFmXRP4wvK0lzT6f2xg7R6GZf49v
3Zbz0dzM9L0UkpZfSlfp2GK0BEcOZzVFzBCAgka+0uWZlUhPHGXFqMNV2wrYh8FKlOyDMvUryLZa
RKmjycqapE1910X7ZWY++AxUs4NmJZgaWklhNNpLipUuXZC1xk66jwTjC6JI7YTiKXF8axnAMQqj
01ZbrBbIB5AiDivEPYPz4lUL53QiZRbyochSiR5NowI5jmM0QtZwE2kLyK/pcQoleqzygZLh3813
V83+Mq/+lko8hWLatNu2GMKc9LTqjvQYI4djqqCU9jXAWboiiVJxa2MeNti+n6ovYzxkaSiZ71NR
2XQfFPH63jb0jF9LKNCTe7qbhP9Dc8IJ8KPGT5/sx+FgNU0Iy2cl2ppqsmNtrybsmpuTv3L6v/bj
O/cEE9lc601YvrBaBjjK13UpfXVjSGE2lub1T5Vz6x26glFXXdl+0vifdbyfO0Vgg7l5xc/ox04n
DFtuCDBZi9ZRmRONDIDjXvccysXWAv9vkgzxejrVxGaLQd0UtHDXSZd+Ynrs5Z+x8pLlWUNcr3d/
OuMlm2BvPGWlVs1IeStzgUhXvvdqcMo8NQEGxWmkp8nYep0ORgo8XeyiNpPNrMM2LuNXQ+dgFt+S
jf69zPlYyxAA22EauyoWIJQ1p+wqfraHXF7Y9l4UhOr0WGeM79zsD0pcx+s2WD0HTTuAYPi22idb
+xD97ubctVt1aiz5C/LlBHrwe33HftPfOXUI9uAxz65S4cWpd4BdXgmVgNw8nz355hxDvP9PT8Jq
fV2+sXa4ADQZTs85de+C67xU22Z+PPkB25R6jmFxd/PC6oZzkniz+j4ajxRCT16MQzCczXieIjVU
QvGrS+KLLNTgB8VDG+hWtLOkAmBRk69oRoxOA5hwdBjbKPJIkKBGBaMfykQVP80CMA3ApEUXO687
Fi//TrnjqjdRLkdKlObVDg519jjPRbkaAis3clBa0eqGFmD25a1zIfxuOrMvG90jknr5GkVWr8Pk
9yn60j1Zar7uAxKkW8OD8EhQWDkNTXda8Rbv4W4WvyNhPJI5VmXtgfAXdh6bTaS7ObtPi1mK7HHX
alu6rTpSuaP862uR4rW+ek5Ff1Qztwy79SE3RFwoAQqakau0gNnEtQDYObDa7GTMW6jT0QSGzZDR
GMXb3MtBNgKrxCiOYWmzvSc5dIZZvYE9bcxkYYwFsrMnQghmj913WUHw5kr+72Beq+Kbvwr6qIP/
oH1+nXIopuunKwpzQr7zdvNOhNcGKNZxWPM8KIXBiWESr7MgHj2Jn/bk3vgInZB6csFAr4lnziyl
UQKcufz8veU+tdI+yH1DoJV9G3QRNWx3kQYiji4oilBH4Punmp/9QNRG4t0To+3wiTgdrhj40eR4
zDVg8twDf4H04qDc20XISQT5dm93CU24pdPWiIcihIlipb0X9eylOaBdZcuBXOdQnPbW1Gz+duq8
uS8Vw0AsLpfU63I68PpHB9njgp8V3WNk0BOKq4607e7Peg86peOxDx4LGkrKcA2ud0ItQKwoAIrk
tlxHvdDeAVFk7W3lRjoT7sKK1BsttUuyh4OlCi0dhcizRSQXxRebUwi26MV536eo3ff+4QceelON
02+SY8iicdL0xO6zerM9mM3pLOCD4WI6PZK9Vmipz3+DdtizFmz9wwtNwIlgu0A4cvJf7Hw0nezg
zefhrluBCAN0gsxHRfhepXWtAFtIl3utKIYdl6n5i8TOiVdEVoghY9gl8TzuoRkE+zmukmc6W9gm
y9uHQm62jl2RTThgrT741LliG+eXkosNDIjNXQ7P8bn/QP6GX7QQGEDA4dPltPFrQJ5Ys1QtFKrh
JR3fDL7f4x6X3HsARm+k3AtfzmwjrTv2uBXPwNWcoazc4VQgEdP0mLVmkI6mEg26aH3ujZPyDPfe
HV17tSkpylZZsaB+QAx/i0b8ZfYbpS7eZex2nlHwoF6B6Eu8xcc+aqXs8M89kW7EgZEtXXJD9G+5
NnXoGfAoAGc+OU611/inE49HnUfPqH73idtP81vi9gKirb+LNZqX+Gv+d5dbDOPzkYIsD41ORxcH
weUKVQ6gRGKxb6cGrkGswGQgGHRPkFsI2GcPXxnLX15IgLTk9Jejj+T+1RK7DSE8sYjKR+Fditos
mO1bgigOO0TdpuIiDZRq4niiHJKuryzKjMTw0oYFBvWGn68XPA8Odir8tsnJK10RybnnPdeQ0wxP
4YmwJHzFclCc/LWVM2PkR3Qd+pdjEOyxAh/GKonYOHC8gWNI5cHjB+/IcsNtIplpCYo4YIFJWG78
1/iH0WoDZKsTZCLXXE2dRpm9lwAPXn8as7tqK62oHB+8KKeoua0e2e1IDzdUT8pKl4szxbcG6QdR
XTkRh/mRZ+3kL3E6Sz7MRpB/d5hRU2VKAx9pXued/g53BS10qCdi9ynwdICKIMBtB/EGiolnY7ke
EQ8AudLD5zT5oBZy9uOLYf13B7/2rnCv5ysNhBz3RiN9oZPHnosck4a7wka0O98vdJiCLiP9VHa9
qEnCpjqFFzXWiqi8Vt53HGB9TMy1YItBe6xl/IR+85ab/Ctd83B3hLYuMD7ztQMrcSgHzTE5iW27
mV+tLpBpi1B2Knbclu2sZGAnv3s0PAbFxhL/fu8SlkEaP9Bpd94g4E/pvyoysfneQTJ4rZt8FGHB
fSlZUvxit5jlaQE2aDxRGCEq+Zclc/2aeZAsjgDSD0/9i3vnnZYGEortTWGtVvf4frlBQmIzCIuR
+epJTtctksSfXVXQTSYywoCK7OlWHvLargNFoSrlGJA0tZ2FuTtE6rWvClbo9KOPTqdBUZWQgzkN
IPDXr1xh3xG+dSGS1cWmjokXrY/nMil5KTGd9eB/vPAEV3t0Y0kfl4Yu0bGPQWwWwEVxPd/UXhjw
5gPy/hAXRZHV8dDUNLvhMv+yS1VA6NzWZuOEhMCkyAqFK+yV8HM9btChjTLoJVbWuYNi54zSIFuT
zV/t34AOTY0nKsCvMUGwb6d+nM9MqGP6mu8tr+ZDoqa1ZAbf5fhnO1Z5QPpWrX5Co5ngA88XT3gw
L+YVzR1x0n0oizReL/WGviRsO4TWNI7I141MnoEgr4lonNLM+r7/w2ZGG1HFdjuMsUA2qYT1Elxb
456zp6eXyOPcuCTN7eWtf0R03BWiUCjhmmVsbs9FKl3b5wR4GCx8P2rYIqalLDVCWjw6mFSJkDml
5ya2zyC+KuafYyWxQTZMq9SGHB9cwKftNRiUrJ+CRjWwLXh81XJ7v0AjhvoHVnUsSaGTo7qPJogk
oyy3mncSVBw6ZiTUCl6ZfStkQvUTDuWIMR8XSm5tnq6YwUw4oXQl3NOCstqxpEcsN9t3tWItOg+e
2u9dSeG9YpYySoChRAeVhRQmD2e4A0Ea63ZrSAbUXh3dNFImUSs6mfKbCcIOhCJhPNA42gYcK3+y
LevfGB44/jUlHu8vx6+Bp/9lkcu3JNSLygTg5bi17sqeGklRl8/wPS2KBWe2p099ZRFq17IqELUw
3Oan8pBh86D3eW5s0LZGfSOq2yOS7OTx/aSbpEGMR/qw0MZWtpl6WbDcUlOpUAzbZOk8qVOQ7LLZ
zcLX2S9pbkKfL+fmhrYHhm5gOJkVSuEyPBee/CwCupdszTnpimnq3KzmvibNZqDLKn2GmCU/alwl
tB4lDrSGkTDfIUo6cYZiow/MgwYo2bQGHIMHKDdIVLg3twoRgVUCmJe9Y2nZHkG5aZSizlmDWoN0
g7QHS3X/10G2xLxQbwdXJKr3iL5Rf7NciUHc68463m6yu2VSLep6XBOsqInzP9MtlrQjt6EQ3GsN
jeHTfOEtTycL1VR9mcpTIJxLCscWrPCQZZGhG0C4pzZktS3UjlmgQd3ltPBR/UBONybq9EF6VY35
eycBeLvEHj8XHVe13XG9KelxvOIJcMxayP31MJV7eRFBwFpVy3CwY4nW1PDZclc7mi/vzvVSUqPl
SUOrIoCmUYczHuHLAcc0hP9Uq4QPPKJp2f8l0X+rumeNqoHC8J6TCSx9DgMH+QG9Ha+xWUDvLNEi
b1THG55GzGDHOzBa3yqDFTZ7T80EXU//WeJftZR4oIzo89jVCl9PnfzpTz+2AK8Qmz2dcSP6DVNi
Ron8xkaDfd+4E6EhY9UF9BH1ouuQWYiLmkNpSTn3G9bK2L2WNdmUrA0YL4cnoH9H2Jm8ZU9uWGVt
G6sHSqecjQHKo+uw1WwMa9P5lnV78cNsjM3uHMw7zpWpkDvMbuL0b//C0AYF58Hd1n+TKENDX/E2
/hpA0jFuXtgenycJn0FEs8XetcsspXFGHiQYdCclMjlGUGXRRwr2LC/CjYEr1rcpst76BL7rvMt8
gomUi+Y+4/1VOhJX2eT8ztxDbSB5h0cX6O+ONdy7l4FVP6vtw7HWKsJnKB1sPycckxbJL/yjD79t
heMUGWCMTltld1sp8861x9kvzKng3wCYB0bAmeUy/jnj2Kab73d1I16Q2NwJVoIi6lI7XrXva2kz
bXtaRJCqfupGceRHNUGMb/IygGMl4txLueVV9aSZ2V5m2iBM0FTvSb9pHG7nbpjDJxoTWJQBbn55
qXDqNkq7FQQcZK/C2JhuzyO32HLU7l3kItSM6wXrvLpp9v6ErTfWFYNfQUjv6vlHHwIxgwUI0WnW
aUWYssaUhGGI5wEescuFW5RcU02zYZOWTq5pE2rUioCx1YLlDwQP6+EnHacfNzgMwy1Ooh2QiKfN
vC3JYJAfyIIIXM9d2S8Mi4IflAVjJ+4IomMwk1xanNexjkMNDEKAzZbbfH3fosR7je+uf6oTiLfu
D2eiqdoCDQF/elsF/Fi+0qORpSnrnjOjLranRYo3USRTb4U7ddUAolB2diAAal1WVR+6Si2+RRvQ
2k68GmiljbwGCYMr9GXfLGfm8whLqauNSwsbdACeetc10jldQCMQBXbjGTPHc2rdSYCbEzoEVgCz
Bnn7bVNLEzL9kpoqfJJj3EZaCWOWjRS5KfvU0t7DY/M52oOUZ/iNxI8ziyUBiJzxpFZTfqt+xGyV
chiYgBiaRZQSRXIVG65kcvjBUzwpI2HYt0yDaSAMI8dIFlLga2WczU7ZCND4VOUyU/be0/XycGR/
+1pTaNM017x8zbykcgXwnNN3BrGj84WsRbdjUZw0GgEiJ5nxtWR+6FoZI92kpLGZ1nE0b+S7KIgT
3PgmqXlIwdbTjXjfx5OoRReqITd8cPbCNkNosJecg7D3l+ZR97f0iSrCy1Yt99Xm85Hz1bPF1pSi
/c+XXBTuMkQKbJLXEdX0pvbUb32NCqvYYwc6cuSAwzv3as2zRGDvIp5T8HV+7ToMp5za1J2Vq3ea
WuBmCQHiwfNIQWNoZewTchJY690SLAdg/xx1sZX68rA0wCfd50PdzfDngnBjN2ZeyCX8Vq4Vbf4Q
Yg7Q3C6v0Wh5Vn53l1WrrF9LExg/hns7R4V3wseP95hSZTm90GYqFhZ3vuunqN14LZeAxJXJHgEI
SiVrG9wMvNKKgcxmavNfZWPzR44+H/Snaoqp13p/3wa2sR/PLgf0EP5ZyjCnjwLCCd+K4T5Fj/GU
liWVfzzhDb6aZL852b1FHLZRwTWTYWht2D7qcskQLwpoG/8Qprai1AAJ5F4cFHLj7uQm1jjVc0bV
0Xm4tj4iVhrhJWGvgtvhiotAHgswXKy9Fb1+z/A4pnLrvce6U1MEtD8yXfqEFDqW15VeMHuFTO2E
em/PaZPFqqWhfHBxelZj936O7sFsVrCkYkzBdNAugstZ95aqN9eJ/PuO1cB0kbOgWnpYsqLcwqGB
Y51XVHABHvxF/1U5WTTlA5/a/D11g6IqEbgEY2X2xn2dlRft41nPk6r4KwkxKp47CcAyLXi+FKNE
AMOn+ffYR4xX8qnPWPqrJ2GNSaju8iIGWEz1oLTs89W4W5LL98heWCEXQMRfjJ/RvVIMmOUi3Ue7
FmIjivC5r6/qjNPGQaOV8jFXhqttyT5mnqoX/cqFAV4iD3BuVG6q1gtOjqOGp9C5VJQ8KcUCOf0n
L9hPRzDjdk/+dUWCfIahCr/15DZ5OgeOG2xElG3QsL18C/eBJnBB95m3LMu++O90h2991daHMaDi
HKY+DRX024GVh8vW/1FedvksKE+0G9Wdaztl7N5Db1NHkISFx/qyBbZyq8nzJWhVvchfX2173GIe
VXiUQzViejeARUkAokP41HN3xife/aoD+ss4v9+qACftvWU4r+x4TJkyAU56ptmg3ibozXYU3o3e
B4pBn28eSVrEbaZi0vE8sXarmKOF7WAngK9+dYjM2z3Zxri6imQCHcLRWKhCo7H1PrQsDtrpvCrE
ZzIWeA8CRbfG34Ou6Zxk/jQhjICqR+sxNRaadZ+N65MLN7lAOt1MpBkb56Iu5jMRB/HIWvyGguPa
NTtZuOuHX7d+SHxNu8WrRSSCGKbjDIHEC7CFGj3gF1MIzUU32EfnBw36YDILhZB3sJi7+iQWBfEn
LPPgO8L8TREj2mrx6q0+XGTTrvNK0dLcGpTXQ+TetE7rd9RSwAvSSjSphrR1KUwJ9O3ZdnCVio8J
8QhCUI9jNuvK5UZaXvZrt5jwpU3DsjEGNhODi0yFTPwYhSGA3aMpvErFQ98NntYMshcgNkCAdSCR
6hZLPQ8hN9NFXKE1PcceHlMWqs2z9uB5s3S8NvYwOXswPoStqZRiXc/Mmpktx0LCMHyoXD6dOHIX
0xc1KMwgIpQ+rx0yiWeKhCTCSs7ZwvrVHXTaZQLbBaniZRY2BrfMxkS6vsg6rKzxATl6G2alwMm5
ztHAC9KxJQwuOOQng41f3rI5yRy27m9PWvPivBbr/QSSDqqSwGGi8GQaQupD5IC2Bsw7/5YrLeta
QneNxiutQYWsEbcdIKtjgp1+raJzR476wssRnLrResxx5r3h6TZGMhnwdKRGKsFpiE+pYzgFK39Z
lE9zpsxwfcEpbpkNzpXotpWBXqxvzwckZCGJtwHmQWBWThN+xm212pQJzHeFw4Kgp91nOlrWD0l9
AbaJ7sseYywhLwvE899wLd3tufWo+6GBAIJKP9U3nbvO6XjaB9Q5mZBZ599XV439dsORkKYvdIYE
3qnS0ezJGntCndG/GfpHwolGBzmWgmhO+b+Ut1pVkYcDRfy8J2GK1pYPIFFGRhhs8iP+koLyzVju
5c5PWV8ZPhcph8EywcGOK9v7HXZkzPKE+Z21sc9KLdbhQ1MYGS+8WFwqkOj2m0PTLZj5+RFQH6ok
mNna1/PysTwWeObvQnx/8omnVjwqWIr3nQLhCHVcoChihoMBZPulxVjhPbjB/kbYybPdw4oxpb0M
Brs0t/1qesVd72KG5/QtZFxhMSWbRrcyGxc16wuy8MXjnBymgShcQ4aB1ZFyiEcvQ7SqKnWjZ4lV
7c9l0S/nlQxOmeqXXFFL4vkDfdBDx6CIiVlxeIlq8u5SQu/PezMfMWtL9ALazprqjPdhBewQf+B0
gC6HxU05TOFr3YQFdkDRIFDbdchMqUU2XgQOFticEXMTHAbHbDTj/nGtCW9t08U37UrJffGG/mYC
We7rr8cYSbs3U0CUykBhUW+juqBmNajYoKerSfH9sK6EzK1x/u7J4QjlO4UBEcOpoSzFuIdRzso8
7+Le6bkoVWTjRbFMcJQiO7m0KVUpUCn7krHuDXa5DqfWgJD+bMVrbdcDV5VjxoAiQ54dFL6fsDLw
eibRU7tgLTufXfMK2dtTW+HKr5V5nXg7XNWPpuE4XFuzqlsMKBGpCL6E64clmVV1UUR4oPlSgrT3
jKa9pL59zoG/4vAsrTzFYlrUBx3BFW2Av5HBX+YNvDcvxGakq5ZmwstwKdmJzqmvDLDARehN0cMn
r2EYFCBle4HW0L7O0/0ZWzLJ+G8wsMOH1GoDbWxDV7Gb0HI2bXnbtp5DKmxt+L2pbC22MT2R1qq4
NiC/7gy3M+jzdTZfY4oRt/AeMANKMdt/sqbOIJc1m+5Ezrzz8kZJZr1doafFWNM0pot1saGQHAZz
IgHqOKKX5MgIOGwR1aKohesI3Js0HPtFGn5oEAupMRJZdciU/d8kq/hltF4TdkSdfWLxgfefnKzv
s4beEmMgEbC1zed6iAPBVjFO4X+sNSNNtkX/rOt+mnWq7XG3Al36pnndMENHLCv7ZrlEc7PbnS3I
Q6Q8M0+OmtNNwUNcMoz7yqNfuIeGhIzvH5glgPVcqOTE0t3b8PQjPqWoNCO/ko5aXXeRAXccFdZK
q3bXJR3ab64yZtz6RFwriKrzN+NTEcHNuqzD6S5XjhchQcB8AiZ1rPy0R6OUfXV8PDIK4AwdSm8d
Meqkxl8OPNPhd9cTaCNAhq5VLjAQTSN5g0vbxt90q/c+xverzzlOjspEmDgeYVLrmPsCqzEELBZp
tP1sm59cffaP6PiP4isrf0PhkUMv6VuWpT3kydSHKS5cqmuT0IbF3oyw192+BDPh9kTX+lKQmj+Y
cXDKaLGxhX9aPt9jvqbvJjacOpv9xcT1CeWc6WHu1HcNAhdKCuZvZBA2/17izErlPdgCfrKiAtBq
K6ZX2b8bAT/6hPms6pIjkhtdMpw8fi8fatmoNAReZadd+dmRZeaCE/6g/T1b4KOqzGv/DdB/6Enu
TdK/LfigG16AIwCMz5GxrQF2NLi0PqKEFDOsvbNb54siG2gWXGjam9Z0mUxf42cPhxzsFya4UDst
hPUZI4LhRo4ZOK+bDR0xE7eHsgYrU0szG9xLOXyDUGA4ZTrb7Xs3xQfUg7kf0f92vGGU4zHsxFNH
aUOHscE8eqKHWmqlRkBdpXwrrKHUpi45fQspk5d/D5o+WOllmHGUf/S6zB7WAu9ta6ZxSUvDpEM/
5Q+3KNKGxTPJ/tyVY2Qwmn1n9InzInu6+8F6MipFpc0QIQ1cmAjZtu1Ot55lzqdpP8iwEGbXlOIp
5h0tx0ysqykbocmaX77/qluABKOG1pzeYiZVGiFWOkl7Go0XKPo0Ykoa6ddyjbgl2/F0bwiW4fgl
xvWiBAz+Wbv4ar5mgXc38dN5GmwJk8l8c+C8jP2Z1mcU+A8L5eyDpgn5CXIvpiKws4rUjL5CI0a8
nOFJpTttejwJBksf193KiaA3KY4yARebjvVnnZgqQPBNP80qLaijZ6vSup+evqGwx9UCzeNfCTbU
96vzi49IZoBWnR1Y6AjCgAva5hi/MLIMINlGHbFv1bf3AAMfo8F+anQTwXbPpGzv2u68Mzsa9OvE
CelsOEhWwyjVAJL1qsxCVZFUEKAtEudHccskmdHlyQwVqeljk2SYp5ecwUE6zDM1unPaq3cBBZU7
C+RfmMdJ3S7mKIE2HqnyF2SNLxculge/BohciBUhjK6a/YYKQz0p0f80dlgIpV5Cy4cHOOk3AVxU
sB2HupMxDji990l73AV/PIBGtraygnKkdnjA/LdbJyxyygihpSdggSe1jfuZvqX9gaIVs4hY0xwK
w9VLNG13JkT7iTsQHpcWQ02BkL/o6kQMCd2dMPQbQqNRVEECwhk40x4nYheaHXNYnmiXJzOUd5kQ
gPo9Lyx2z9+8jmolb6WQcHKo9sXiFeQU2uPEk1NH365QTu5lOnYr6uB8tzGnu0/P7UZh0N1ALEVP
Lj0zIugYMrZNbbJcqRs39O/yVoGsd93qSCo5EysnRxaHSvH6DaOs+PFqB/oB/flpCJMafsjXS98h
H3pAodJcSbE50M1L+GJGyHg2pR8RdfwQRykZ12lZfkEgLTjVjU7VTzsyj2L5qGVzjmVWDBv+jGDX
FgPSQhIahMDANhbfYYytJE3eY0SjtoRMxJ3dKZggqxiLA9oU5HaMmQOI+I9HPW3CYIpN3sz9bV7w
EWVJKZp7sYrXhh5eqMJpWznO78sCQLqDolQIn8EeK59BEVdTidBilN2Y1S+ALsdUhZQAxVhDGdZP
GJZDhNZklzFQExsqNiJKAEnBkVmNN1NN4TM+e6SOsmp5HLlU3JyAIzWyHlA6BEXPi64HHXNPNwVR
tGKhA3Pm+lUU86/YmbFfVrsCnJ1v+p/39nqzWKFywPrThFjz9XHPwrSf45ERSP1UFj8b8wuTmZPm
DUqHUCwoqjpKLDf8LwABcZUobiGk9kN7IgCs71rKphscvyvWEqefzWJvQ9tVT2JRHfTCScETwBjH
0gWJn0yEIL+cn1TfaLqK28AMtJZZNvle1kL2RGJGW59csfAcukNA0WnEuBhPp2Pm0ElFHlTvbua8
DKCA8/1klXd4QtWl4+i4vBmnsGkJMvmRV7rf02bEt4pREc7Hx3Ke80bFQFNVCTRvY4kDl5OBo1rD
9En+20x+IkkNv66fki+Zrmh+0sWdSrPG7ENoNvEYP5oTiDXUQMrJNvcwBWdlcpWmNZ7N13/sx4gC
qv9aRYTT3ov/k/cgXpifigCB2x0APkwri8FPor5uddaVKO7zWz/LaQRZKPU+ZroLMDM+XOwGiGjh
R/AdBgaUqGRa05AVAaDwLpLwPpn150UtRWKREGtHNNr5bfU4GtB8a5zOy/az3m7ZdJz2lgS4f4D2
ESif6Nwh8urE6jnab7Mqtl3nUFQwwyBbcIaRvwrVsU5jAx4g50kIe4dMFxxwlLiKCM4N6Dgz3sSs
GnZ56yWLs1dNDOqGdafIhR2iiuVF91uUvN9/lGvfvNdCjDhBirKa1ZJbzJlFwyMLCKpp6jw75Hrj
bAp/TYaimN6P7BQW5iqGt2nl/tH1oppqchu9TRvf2XpPNoqOQ7dFxDPHwk/ayI1J+MhX2FYdH7j+
lpUgZlPNyWlmjFK7oNnPtERCm1KyakCv6BjsqWP0Gq9s1GVuqHMdq3qHTV7tucP5sedfiOXQl1fs
+H2YeNbxLuJjHSn8ymd72Hvml8QtGs2YpH7h2wmtD+yk6Mu0rMABRxDnfuNFfrmGWptkR5ansnwl
4TF/ZGeT9ROGKXEFPmaI32/7J6XMvhvq+/dASUWJxCmxtraoMroNiPUzDYy4L/Hfa8ZAEAq771Fq
lvi0S6V8qenACe1DVmS2+o+/ilvCwuniuzJjbALLU1kwsWXkWh0fOXqSLZTO0OSwzVmTatZkBlxp
/NdFT5Q39uMlLw55VeTbv3uRwKlcqeTJg3MGWT7hsX8nXwXI6gyShz+JKMXSIZgO7yRTqM7dZn6M
Cj1YC+GB6COgIRKaO2Dq82njyxO0LQcZlAsPzWG972RzG6P8wh8oZMreODwCSx+6/l/2wELTPDIB
XVcF/JpzQJ/S2L4JsC82zR+Vk12spmqdgmOpi5OhBK7m6Z3Xyv4spcBATOMIq+95NLZdSXAzuKQ0
8a/4RTcGZMUqDrAnIUgTkbG0IcHD1iUmszZWiphtjgJG4WvH1Szf7Zd6uJ8TjDM8juo5MnSFbClq
sbJu1F8WVxwNGcrquBE4pvqwwii4zWW3Sdrx+iYvTgczxhUyYoyk5CB82L6SQfrZ2JvFIA6L8xBI
3wlc7kD8ZQBN6PIm8ateGcQen6ZW9jUz4FYb9eSaDXJ/5Z5kXHCX0vGqDyP1QtcgPbiJcGZhA7v/
F+5OePrhdJjJpdDzBQSX/ohDv5q11iqyXf9BPkVcojZc/u3Gt3kQzFseU44bNo0pNoK3Uu+PRgh5
9T8QpTxkNAhYp0NBeWmpO6eY/VEnUm/qeQ/2lRVfFYkr7AD82I7A0fjQwnRZ1J2YiY4xbJ4U+tQF
XIJHK+pE1DtSLA+oLyBHkLJT1FIezDReCyqjAtQYs67cNMUqGdF7v/QoWoxZgFe2IGva+hPsEjYd
WyvqZHHdHgerZFh9UvWJVBnJ3iIlnkZ1hFmaPhsqwRQ6P05+pTDuAQynxzIri2ZOLzYsCZ+CXDkj
U26+HfCrXdFIvRIzCBYN0ixkbEQi7z+p9Ca/trRZjmsCIxAU4OvlYLbLf/Idreui6kxaqMYyWnE1
eswYIRUaxCZVCziOO0qw7n4aIuM4g5jXaKOskJR0rkyNADldOAwjDCs4eQbe+5qrT7GeCoa7xT2E
HUWG2u2Z4pJtK0bgwlXuiqAYfCAjEFvfA8rGfHLtbSKTAxfO6+8r9FO6Bc/NFDVkt7tRNBeKII8b
jO0KmCzBDNN9TSyAJidHHK5jXAE+5WNYgKKpxtw3MroqH06p1lKHKGIK2drq2Y0vspFjVyfE4DG0
KAD0jO+ia3p3U7HpgovhpsULC1MIFbAsE7RYSe2kYyplrx3XKmFzYMDjiqSAUooOiOyVP7PXcACB
0Ta4FjvNgyZqTiYvxxfTGvQwHPwX8ezX5eB3lIaDQOIiHvkhHHviMN1371vaO4DENXZ4rgODIUfh
0zgYd9nvJ3OJH3MuuEd52Lv2MiFEzceuyDNR04arugzjMJMdhd0cVopg2J9GTpPrY+Kf86OqhKCW
mAlG21RPn7PthA7+IkD3yarZq94fcFYkoQOA4lKlAh8KHVz+iwgumIOCoToJJhll27r97eDASsG8
p7gvmpR8YMdW1kd4l4gA2sVMF0JrghhLjItjuH+EQdJka7tBEADdz7NlkIehRtgQTmprlWcmqQMC
9RslkqMwHVhGl+K3hrY8FRZigBp+i+9aY8FH8UJ5fbCm2nq9cFF/F2fNYV5VJY7R+ISWBtrergY9
AuBAaGE1+YAdiYHCFxNNqPAUFnmbD86DuE0gbFV9xIUKHOBeXA8cP/3rpgZciE7L9h+8TJkbsKwW
QjaL59umIet7v3rEiHEO2oYc1Zd+4RiZEYoHT6ZdZsFU8JBmh0lLgZ9wkog6xVc5G6iWldZfWM/S
7fd5u3KPRt7ReIIx1JJPHqS8I1PxAwVQ3JQDmaNbRVauY+8c/QQC2E5QBAddxKMG583qnLqCmNIp
31Q9K8Dj/SCkbdporDvmGod/1Nr0ytvOiOxEnBtR4DGW4X+vg4kYrihgCvge5tzfWCxZhgpvreGb
Hl8zm+S97cCb4dcFRbn6GjAgjbaYGRUmcDjX0NtK8yFcWIalijX4Kx8AeqzWZ7OfVzHjRCwsKQ5M
ERX6YgkGWvDFMXZoANsMYRDjlalJRvcG3pZVqt8rjgEZh7E3f9NFqLnDgiW6HIaOuVA0P1bBMmCV
nvQVBGp3ztaB8K5hGx4mO/qQMisINew5ho8lm3Puy8W4fOr986VAPNWh2IspCcLdZfcTe/cihi1V
viCp5E9chpyI6UYIJJJJ2OOTHIPh9EviyEs3WWLYN412eV5BuqeXoIe4is4ymhSbsEYO2OvujaOg
f/ptV8cU2uqPZ1r8mQfeADnpOU/64TacE/te1YKdABwJMsKrVttBo8e1DrQ4I5wWSg6xUkSnaPvA
IqDkjkKCoaUI+ioo2LwZL9ZpLRrKR/7MfmOS5yn4CN0+QuLUZTHZffuiDl0LyHMIkbK8ZxK5YCE2
Bu+EEIFiWGJ9tpb9eYmD0YA16ZSwE9NvEQ6TgXwSkOt3EKs5T9BTKTeDSTEGKw0Dl6G0SKnZ3rbw
n8tOQrgXUmzNZkfs8IZhAK7R8ry9mlSmBQmjO0vhit982EY8b9nUrUCNHU0CYc1RU8QtUczui2Ty
c2OncLa9m5AXp+7YYc6juMMd7vBbgfDqa0LajrT4kiqWeRi9SAq2AfcxkPObxp/c3tZ3c9yoEHsx
Eg2fxeLaQtMa0q+23LrqjFS1QQK2F6uznczdvOofJALIkAyAA/xXVxb8AxXZBobGQKPb0SESCBvC
6YvFf5zcWYGkEcsgpX4kc5gvbANIq/nJYjjp71lZO/5SEk1oMznaEojyVFvQhAjYYbmqkB6IL8+V
DqCNmssmznAMw0QjzpaAajy+rW91qfsuCuALNHBzr5DipnJX6F4p+4NmJpqwEJzm0d9+kDP5lDvG
pLMw4de2+gkvnM7Ebxm1fkSXnyeiS2f4Q79AjxPy/DM0BVTeTwESQES+NM8otrNNZPd8ZYS+Ruu8
/K28HY/nkiPIYiJufBCjp6Pwll0fnQ2URjXMRAXutoPaXzyn66gvUb59pdFa3/1rAgHs3n8g2Fti
z3wcggGKYQdaHhw3tl4GFLeqRjqpviy7mU9SSf9rlxd27wEMQdZZZ+IGWhHwyFCqQQx6C3ocxTMz
C9ibcnIpolrcArnZP1Z+SXWjdt4dmansh5QBCePwEbfQC5/NrB6BHTxbFJ6GCzW0FetwcgXnkIu3
qrr609e9+kIbaJULLSlHdxbIThErGVjI+gq22+7Vrw6TPkYa4kzxYZNGkKzz32eY+KIUDwVMFf/S
G74GdHhIk7ib9MIiyoUO3Snf/tbV/WfZsSlq4SpJGXnw3OLNh2TZcJ2FVftxTBTUQSDvLtf0DMkP
WSDNQScpEFop/8llWkXA3JyRl1G2jRs1o2Qr7DE1FsLzPi+K6+TFayeoCOBb7KEqjgNmYUt2p4tj
tl/ZlWftbBFouk8Qkb5QNqwGtzYoUtOXz5vKflx5L+1vtkSqZvpJQqJ9RFgpyLSlIRuZy15ogPvz
5/ktnz5DFVEoC4qOLlOQoU6wxWG/AEtoe9D/x3tAfTIjpoUSAWzVRSC5USpoMAhM9C5HfFfy7nl8
bebx4XS58nW6A88AonZRi6D8RwJdC58cjpbAgtufinGHMzzRQp43fqwcVT2BpSHRrfB5cTSaHa5s
AYfg7inRF0hkVcRyDXOFS2HAvAb4eRoRYMJST+yrwN2zWaZub01tOzoyz+jr35EI1KyVPtPIUMbX
W0r4JdTdIocJHFwwrMja22Wn7q4AxePo4SIVZ1qlueMLHr1Fo7Zw/u7HlddFr0KYGU4lhfEMPVly
KnTkWYILaXY5L1LbzvLKxaJwwsb5P0vqlxCodG4EDhoStVkETRbSRWXk+vU1IIQwqYoZ6L2oI+t2
8tVdWcsFQhIWnPDN28/6FemHJ2kAopMLr/CHnq+utNh3QH3rZM+Q0/7S9XFNrhB3reZDQSZIp6+e
jzeN6Ltrc//nQGILw7maHVAqixXxGt4LfqkS1N/4Z2ElnHp78xE4z/Tiamod5DpWZZWhME3dbHP2
1beJZpejWms7ZrY0OhUDHoxJbyNkzozKUzeZD49+RW8yI8wobvUgKP+J4atRxlsYFrtIlEfYEa52
h4SdMZgto1f2oMLJP6uQZGA62yFzTyk1yFMitVM8wFzBiw3hRYKKLW/FLSNZnUpol5Wrxr1y4WFs
fZp23khig127Ld3Y/JK2hlzzAQ78y0ZOCofgIjBXF8mpgAy8JbXqnYG6s+F5mDEdAp8LxY1ebnr4
zTADeWsycP8hPXO4LeuqZ2owj2wMJ0oO7r+k6C+aidLRV/YT0t/mbwPW4J9vxxaJCNeT5AHukg4w
gS8UuorK9de5gHmHcVxypuMXdLYLkGzJPuBpiXRm9LzBc3p9Y/QtfHsHAHZm6Kcn1Z98tSHSzdWM
lFpRN8d6w2u6krW5cF49ExDIkWmtupXNs2iCmri+Wm+8RNExgohgQ9c+PQNDT9bo4K17HSqAqma1
G48MkZmbGyxS7RF9+6Ow8+PUblIZMHsj9srkqpwRjRD9taC1EIGYH4IPSQ4SNtVNJYFBU+0b6t2w
m7TVTLw/TuBp9uPsnkwCAnbIgSuf5WCXJdmHinK34KsL1LGXrmhaoqSl46F1qbKPMc9VTKEcAUzN
hbOfwMGqNHPtteCUvnWjuSf+Du961BgXW9LmI8nmoRCV5bBmsutDg5WVzyQOplVXccQhsgysn9Pg
d/tUVPhrxVEzQOPewJjvqjvvNnalNbCBF5P6lrhbRL/cD2tZMGO4S1NiLxVmYCC8FFHlpqrbfz8t
y+BfmpndlhJNoHkUG2eoIBxLmUl49fLLSEqWJFa2b00zoywFBo01DAmRFXNKleeewwwUgds0c3lh
7a5RM5QAjgSvEWniI8oqSQxxegnwqf3tL94cVzzfmod+o6eQ9s2GY5DaSfs7C/2hO0bEc0KEpvOg
+XKwJCN2UsAMEDTtSisIFf3uiiuG6c0m3wEBEpi28EAuHENHUIS97oocr2N1ZBhot857SMIhLcnP
XNGk5/4joKnIcl6Rh5dUhJA6IT630sabgiiOvXf5vnf8hCJxnnM51b6AxYVjy4L4lCUrMvZtWAZN
f6TStZEOwrNG0ZNmM29YCPsY2bE16sTcC09u7kksO9cT9hztFYcXIjPIbybz5j2Byjs/GXNmQ7Or
rJfhyOgq3zJxRAJKesmDk1TyF+ikn3yEueJJn/m+WlLnUi0Oh70qKuHwtegas5zcau4C1rlOyKCU
MPePPe6xhEbdbwrw1JM0mpla2PZ5svh5lJkt/WI1BR0vTSibbpx02nW+OViWzF+ZtemniueR1EFs
ZO3CNS+c8J2JeaA85Ra8JyUbN3+Ab9ReIh1LCZzrB2q0JWSqIoFIGXs4z5e5ch35zRLkvlLRkDVO
R9ummed89OwqbtV3HaFys/8JGimnRHN6IhXTaMYKnDYPGpuqUw5tTWbqRTdu3KOtCRRrDf5Raeib
bFGvdCK9EYCCX6BJh/ynGyC4VrmI7K0GmQBzTzGVspXNDdbzJrdJiBKXhxPC6Tq/5ENeB6as0eZk
4YhlmQeQC8lTHXPeKXV9A/hj+Hl2FUJrzFYmsJyCjxT3mHb4ENw8gkurtRnYKOCcLUeRH01LW5uN
p15yw81WVQ/KGfUq9D+e27VnMNQ87CBaFg9eTSHJentDpL36IocNqlUe8SjdDcUc2IVl5NwXPMl9
HMDUrhCnVV6zZYTvooueafC/54ErFaY5LLa/L3PwxEs0THeeKgMDkFYWRfkxw6Fu8kD51LcAmtlc
MOsx1JTLfMcaQaW1ebU4Hbt2URVIZmFhq/zI0oX6OTOsnoWffabSu/6GHNW8ufkRa0HaNyyLD6EC
nYbl2oejK2Fd91NOYKY/eWv1sF5iFU7O+KFkpGfWiKEpXieUvlO7aHYGvwPlGca8mSi3oLjOa+EA
F8vC3i9kg0YX7R+MU0l4e2TcPV7thE/8G2HV+78U8nq2Whw0hoboa8GayToWE+agvMyuKBOZYAh2
oFD7f5+6bfZUiPdAH9Hsl5INt5SUPAmeyNO0+Sc43ELepITwbj+VMXQbh9nKhHy9RJpnSjlu4OLE
nmKAACVmDpvijXaRGpxHqAofcn5MbqxBee1APegS/yt8g8VPIV0pVv/6V7lJz1Fux+CeHhKhlo3p
3AizlrhY4U+n68ixQROFWrkN2pBdDCZMPHcRs+t1pUOdoBT/g+MpsIiQt67pXrajgrKxzMjnsiwn
T4oyBTauVwlqbRxNKpOIZRvPBG4qo19BX7IcCp9kUey8ltARILZFSzGUsYgh0Qt9cV0BkyvpFptA
hy1D0mviQTqzG8bCD9y9W1YF4Jryk1j/l5SxEUFGQuv70aE6veI+UrFyqAt/Cwe9352uXSs+vKgF
dZHRSIDIH/wvezgXxCX4r/wbAWcbXjPjZhgJiXUKa+HBhIFYIzLg1aSKhvRCZrunmYdUgfl1O+oB
RHVUJaVpBlk/816t2VDhFNzrrwnMKAHpeQ/JeSKqVbTEYPaEB0hLy8X4/BChdTDaN59bG55rPnSH
U6WmIgz3FjUOnS7duK+TynlKTqwHfm8cCtLUgS0gOPxaIDSilPxhz7K+aRUEpSZHxcQAz8U1STva
gMrnAGqjz4hT+37sdSqQxUjoHtHaDJ8Oty8x3JlBUmebH2qN1ET5D7AZ+t0I6mJoVESCz3ha19tL
U1DZk8E801nkMYgU1XjXgAkZXGcjbncyeF/rQ5cRZQY/qEeQs3DN7TAhWJZpPaL8Wb8btAyXNqny
IBnaQ3AMbdTk+A3hgpKUn7YUncUEglv9Ik8YPF5KJLgswBWHrYd6esahSfFDyvAqPI+R969Z2Wry
/0wDOf4YIPP5XGjtPYA74ouv+Oo/H1JoiPkz6gIhuhr/80/GpTTTqnx4aaBU8ieGRFkQcbF2aLez
MbMl5PNwAAvzO31FApOgQ7Ci8XmNTZ25FDlhdHYhIKo68CZ177zkvnWj0rwICLKiK+OhOSWhGlpt
8FTGp/5bNQGYgCCYo8tTX/Qj1R24sVQ5Hw1DT77IMK300jOGHV0wh5OAPgVswtdultVu3B5rJZc/
GsHkq+tzfJ0YFDJ9qHdDK39uvw6yANqotO7bJNfCfm5HvzjwgF2G03AHwkrCLXFS/JrGTj9Zm/UZ
7jPjCdYkgV8qn5/aN2UN9KKPpJaMuC6p/aiT1/mS8KsgvjxW6O4pnixugIjYK0bb1Nuos38lFdIP
CkIHBFv0o0rCsx7WxUdjrZ2ebc/Ur3MP4EcFdrmHR1DsjkKjbFougQ8WdA1JeRWo7Q/cvmyBFyYa
5sIMk/0cYKdAi+Q+BSkaDbOMS0JsE0r50HSP/qNRAvabOfW1jG+ZWcf8PuICsbGXiyOKEgVEZdtL
RScMithhD6Pjhkt7XFgquk+ZQicsS7n+pv+N/keqh+Jaa3H7Sj4Q9FmWS7U4F/WPm64vZdMJH2mq
xAEgp3GV8Z6nFUFnxpj0UCxXvfIzC9P5AzcO5gz5YTVipfFEXXnAQvCOyhEGOge95LtJRvBfw8dT
ush8bMZTsL3ANiL1KOPXRRb9V53EsM+jUIQFFfgiSkAIahtX7ROUhF9wKDmoA/hrsE0jznKmYpuY
37FZMUjGctQbKQfXtnUqKDOdqkE2iUwtUnOl6mVBTbyfCzBpbfTo2c9quLRBm7kbzVEkIfE9KlDx
iqlTOHS16+Dmw9HYFYhbdL8seGOA6jHM1KmvVVx+R3tuNVHF46NFQt8udJEuyDt+XAR7duc26OWR
rb3rug7Pi2z2S5ow9DUlLVExStFBdHQFvcP5RiD6Hkm1ZXqicuxLItCoN3iViRm/B+ow+U/pGABp
JL7SqXGk2I0tvOciNAJIxsxhqt/wGUZs7rYZzg6j0/OFIYb/3Bn4tlIFGTHGWDZ7I+AcC3chDRGb
t6TNlGHjVdKQaw3byGyZTMdzJkWs8Eqlh/5CrHhWdPk4vhevvc8q1Gidn9meTL/bDkD8DhbKFPfe
AiXPy/mCc1b6mW1Gh1xKB5FLbLumJEaqKQ00Ac+DvPw5rHsRl83UHFnPQGM90O3RIYs38rFmSm9M
oiH7jZRgiei5SkAt6IBUsu2uBFWrpaAm+AZyOJhNyXRyyX2RscT8XiDrcxBB+oKfeWvbUluqtKX7
Taq+xHdN0nIsMu8KmCjA1IvysWF96dG9kM1O7kBwt3FlSdSwej8AG0PlsN4Echivn6bcO4kJwvxq
4akPJIGJQNvzVzymQv+BhdBH8ldJOWnAuSOK1nPHKJsKp90tZI4nKxaOAS9TLp4LyaILhZQYpjX5
jFZ3v1gi49Qc0z2O/0GwpJnpNqfwlZi4/N3nMUcj770W1D90bRRuzE4MeI1fZVYM97cYsTiZph3P
mAILobxqMEo1PT0XwK9yUubZZZ5uOuyjNt3czXO2CckSe0qR700O3T7OHw2CBNLSx9JNe2UqJQUo
RHzY/6QaW98WwRUz2P/OPqZtKCiNcSKerYHlihmtL9yZ6Nj/Vdog/AC3qAACNSx7WjvU1FRwswtS
LkJjY6yqVFBiVyb4LiMd9OJYfs8TWm/VBDXO2GEnm745bMceYIrSv/roEBCX1EGWHwjWfw68tGQb
HmehLEs37pZBL+uOwJOqgrTk+xj3/TrhUe1jbDIdWkJsbVC97XJMfT1h78OcnKzbLFmImPM08OgM
q/mu2fQckrFp3GaNMnW6C4ywGUfIMPC9iuIDUIu8hd3NIS9Ro+bhStURHqD05gfdTgHxc1GzJWiw
mwxT7VSoBTUfusBKbH6Wc+LnVved0FVQcBzgY8iNdAmC+hTUlwk91leX9ttOmsmt1yDa5goNUDdC
SWy/7PwAprSsXafujaEBK+tW9s1RaC7iv16Oaag8xfuTPynJgGz03bopALnhxnxk9twp0Tp6gwPS
hVSbAn+jlxdKvGzSoQrXZ2XNrnu+1GL6741QKhhcpN7Ikp2wTWfqwFV31PKlSRNVcwmbMngPlkUE
V0wMkft12cn4yQ3HCuZIgyuYrJeWTryh59fxuTRGuy0Sg2pocGP2S00UUFm8W2F6EYC1d2KLa5Y0
2V5zP+zBCiU9CTQy6qoT53wpuHknXEnQQRyATqd7fV3CY4JW6QR5tN07mq+GtZPFVXoiEHMgVtC6
k0tA+CvSdaPzgVsfpNLQLH4J42AViz6H/ARJ1INh7Vv813575QHUaXDVzPYg2AxTfcenQ03GgDb1
kqFRwFcQzPj3dLb9XX1pO/EUHTTXrweD+sissIUmhDK5KdckFWG/vh3c38GbIqUlwwX4aTOY6vHo
YgyAUvkFAV60ZEmg3DW/bU9Qo33Zl6BZUg0ihUqUZ+EIwi9CquiC4YrRMtYVxtj92UupvuXqc27V
iOI0HmqhJo4ap1KbFBF7xQPmyiiVntjayN8zPcmSCPi2/aJWzldXBmdNrMCCobsoWKde8RYKFUuA
ymi7IOa/Axq0isWid1e0DYc8NJphHasfLyvH+yQ2LeBNsTo4USoQJxhLw68xE+QtKgmtHSAZttu8
83ThbkaoKWlbonI/uT9lhL4KoMfXQ1GxjK1752hp/RmoFvjv0DbNxl6ZAWef3CnzbpH106y9C5tS
PB+p6Ez7FCfZdOkZgakiptMwSWuwE3qqvvzSXN3Mt8H4exD9q0X1i+uECskeuN6oO4AjaXT6NYZi
j7YwRWdK2Y7g6Ugs99y0cYzPDi9R9qj0ufztz9IjsR4ObqQo4uSA3K8QZiaY09t1fUxUXpOM98Mp
DCdNlCUjrBFPjR2zRpNg8z3kFJ+ZW6eOj97xF5RCYOJJhCnVGdTLi1k59O9j3wTfTzG8xY8Fi0fT
y2qNeJG1bR3VSTcCUqstD/bU3zg9TMF8oIT5B95PW2psqqJdEKuBD30mFfJsreXg1Qqk3IzsL6iC
rKTkknd2INvb5z7jfS77NOl4s6gala+amtnUzffbt9S6yGf0XeE1FOsZBS+j6EGZRrnbt2Zfg9rc
bfo0mLnoJdslb8NrYuuuILy64M2BIMIWsIGFH/gW8LPipou0fJWBEQdD3xS7nwA8jfdcwGASmu/O
aEPt+gGelrIwCzSsDs4bJ/pWUXYu/31Xs5Bvs/imzpjPA+SULSrWfV1dpwfhlNR4JVPQAJXTy40G
xm8WCL+NrqN//6cQ4p3bGHvBL6zJqnZwTwFZoCApGwW1zu2LwfXlL24GVaEDeJSMMwC1fPCYhGvH
CWz4h49J6e4AdqcARVnUUDEL19jcTGPbE4rnn4DPE0oD68fYdPfDuUZEsXJDst8+e32bnZZJUqTk
t8i/d7GVJm0DD0BUErBgJ4Kj7P27MMSTNq983Ma54nIT0vOOFt7gEZ2MDfPhOeLK6KsMzYrpCaub
3P54P3CaOmiv+Iv6PumsbtEDm8tCfJScAHa+iXetB+l4NTWnsbb+YIXpdqhNVuxbEhYd4MuP08MX
F1l18SAJ2aeDr/oVmiNT9r0UK/Ic2j++8FOgVsAIV3ejT2Y7cOoRryARMwDB0lSXCl2ZJmr+88NU
PeF9x4dh+gg9tKUg+xlq75//toMVhF7jkFSimHuZn4TRCG1Y9aRDoNRpxgwocBLWJW5ZWcVf2p4a
fgwn+RYZNsA0f8pSW6Fu669F0svUXRQq2hjyApKFqyXqDTimnGBDBFCwXawhqFexEODrMTG6lEQZ
qZaubO0uoHKGKlWxyBG7PSAEnY5EiWLn7DY6QGenIztWllbUcoQSr7PrKtLXb+myob69WG6y97RW
cK7LnJJJ88yHX11Qj/rJYzoBug7AdrrlDaSMpnGJKTWAJde12Zxuz0H0qHcWaLQKiQOHwJKebO8F
LM66gPTji+6KZioBiGKml9twFKoylqaNb/M6CmUO6kIcGsYV6h5FFNaJHbkwULWTh9bf8nT8O3YU
Q6w9kdyCgUxRuDoAX4akZiymxkZVR1a7j+iW8DIeYy8YmnJ0GJX53ZKvr/Pp6FBwWzbaZhh7i1rJ
IUSz5talUD61PivO5ZUfjuXDjf/b6UcXqy1F8L0YunfeS9KLoHSXnMYgCMcpfGW976VHRj6kffBw
khGam3GMLKG55GqPzj1isgxQXfh979iT33KnT8qZNDZlE/0NwLmjG2im7bB3Abuyv51lG6Wtvmox
tlrlW+WVTUpsFPhQk3FbmoZ1wmbGCgmS1X6g1X3omHEW5lmarnZgwC8sbAaB2FLiwuCzhTdDuNX2
BmkuKCed71hzc3bEv/0Msg4WDhtDCe+ZcDVaZgiTRiJlkvMxTezpHvVp/aSyItp4GDwhnwo+KYdA
heXF2wWrg/qXlRCbPWaryHCNQMyO8Yvw3tiO2Fug89p1O/I47Fhcx35nX97XHqv1yQKOxhGnlobA
MzPJHATxlUPnHsyYWyxtl2kgNZZV4UtS/9zLCCyq3CkJJnt8JgoKa88uZXt8Jkf6bV15gRlLzV93
xi2QkL+4Acw/ZuHn+kgbpnt63OCZ/IqrFoXI09B9ZFqm4oHPONA3C2Qc7Vf9VWu42g/f3+ZwCCFC
sDqDQ6T6WXn6wEuc4dSPXmD9sKKL2hNd5QOPnsGHPwpGUCqn6daJby6G+Dyl0mFxh2qPVyH+rH55
sjml/jGlRkTcNphxa1+Glm7qVCjiuYQ8/GxO3VzATKc8XTKDKM1zozOMPTmRpAzvvIUeztTKhDTU
8mxRco/ZyvTy7NgW/hYsBsG1yjLM15hmgnvD2lEhwxbmwG1tjaco8e555KSWjJOFA7YJS95WQBtO
c4xYEbtN1HCMiZkmwAWlwE+q45Y4c+1Ef2OGW3KqbxhVHA0+Lj3hsB4qY5P5PCE4Ea31lfrRiciF
K2XGhO2bLknRztWFRMWIc182F2983VyEIzlw1WUO4X2IaEEcUgokb3Xnlk8oncK/haxwZp8hyRhC
h6hrRpBaGOhAOfQ56/JfMHUo4hNk0xzNnDkvAQWdq+1wwtBXLV/EMbg9OK1JeZjZ7c9rgK313wia
z3mFH6eiM1uc7VezHzP/TOCkAmVaOnP66AnRwBisyYJIFi/zQNehTmbq4bJbb1V8/gnF2XwCnPRN
B88XliXQUwSrvzntjrbPZ0cfvTpi1YTt6H0FBpyRzudHxf8HsEjJ6xIzLldIa1MjAUOTogA+f6ea
mMVtWJjdTFPgRxsZoiYI7gP99yO0uYWdUHQFi+PXq57R6+EoM7WL+LoS5kOwmL+2dv+VTvIa2fP7
szSFzZsKZt5/eVLgqtP+HXqv5KV9SWSYzlqZnVBuyD4MAcOQOxWWT1ubgl6dVqs64A+w+EH23NJ2
oXHbYfD1kL9oPoqkgpmgsJbBpiaP5QEu/zczWo7h+ZYKr9z2FRH0d2gQPXUhGYt3geGCfqj5Szgz
YiNMWxLvAvFK5dXaTG4nC3NDHQcOlc9f9v6qVcMB4HefKJMGdoEtFkVLTbEAPQ+IyCExrtiA4niS
jrzHKPK1QTJkeJ755uDRo/kOVdpBtQ2m2y7l7pYRUadPOkpi1jnu/d6jo5VlUbczJDOndC2+aUns
KpL0Cfpse8fLa80W6nHuOrl7BgCNJy6x5/qj51cbRw4H1QF/iV0k4GxI981Oj+4xwm0iH+1KUDEJ
8XVCDvN7uo4kAz7iuVacwBE6iXz9gf2T6CmeZiiKjFFraCCJF2R2BWsYll0tHmQNiKDvPXIHNawx
oRHU/+nJCFmnLwpDA5R5Yd5gUo393dSdtbVv1PEbAJinmPfohOn2UGu5zND9XP4c0MEdRaUIVQlL
EOPU+IXFWDwkBAXLtDOoPdR884E/C4vkDzWBUEj6i7wq/sbRxkwzImeUORLHj//4iJ4UyZdQXboa
MzFsRDKGBtmzOHiPaxVGnJyaAaE0NbHO6GhflzzDzQmAUyFx2wqV5AXpuMqMpv68+2mf8HQGMqo0
76N8DnvtJtHACk/0WysVD8TG5uZuBmlW3t6zafWmXg6wqvHy49DzrCQ1LJkV1qxazSsOzvDZMbhL
aF+kdM31d+BInz0NxxjUxAuglBt2Vs+suSLikmforeAdX22qtcfSYufw3ZEO2AZEZsyB3JhgggYd
AvL2j6EM1LwjojPivpIcEGMcRtsngxM56KnuzO0bqVyJi40+wVN0ypakHDKlQ7VT7LwNnTXCqk18
56twCDmb3g3Q0Yg3fAhMy7YCPMa3MsvjFNcvzgbVvNYXyYEMTqtUgLhwCDY1jFZoB6Ch/GI437sz
ByfA5neJ7pklxVKyngLh8RBdU2ZS7b6KkRSqDLssTTUtUOXrdH9vsFAYxl3zapwFY2yw7vh5rYOx
0EG9co/Tw8dYyeWabuqpeN4yofIRRPqFLr6M/TzOVihi1CCqcrm/d4psJmZNyWLuSbUOmxUP5sgQ
+JYMXfN01EIwwZ8bRKBKmBZypB1iOoymi/OecP6d36TG3vfOXgALt+OO2w4UjK9GSIP8UT2zL8n2
9IBqA8BvlZywDTSVJb+Td1X8MAB4M0J0qZ8S4CQE6B2G1yZI8keXh0vlAABQaWL3/K3DJZRjT31P
2vXRi/ZpkwEaa7rKu94tXxqdsfLyR7f8lsMuKcmCnvgG4qhZi311qd12HeiOFYaj70esDIU16Ge3
m7cLyL5f0nIOcPerWC23CWWUt6rbn6d/rGyAUi9RajWU2dng3ADNLqPvxoNGiC/niQsmRtfq5fMo
dK2qkVvqjBOb2tYgorUNsiUtjO18/q6N64BG+s+PfVE0mhS0pEO+62hYMYjW6cQaRugJfJlqAF5v
2cbdBJOUxKV5Nr12KHfcABlPBylbnI+fQVYdgMik9BypUYiIxaWn1CaFpN/FQL3CLZJAI9GV/pSh
q0J1H0TcpAE5riKZNs9fdlM/xjFZcH+NpO2qRyw1Tka5+0UAIbp6BRcp3Kw52F7ZCfCSgAdPlXT1
XvkwHyl7dWmBLS6Tl0lE/MlXHaXr1O9OAuEOSEZGaPeEUMPXngnotBZ3FWCQK6LWBW0CDL6WDa3O
dBr1wxENb425+igHge/cnUe/GoHY+G8mJB6NEPOcsCISMsCYxfrVwuefRVj/Ff2ZTD7Lv3SGmFcx
dcoSGuRjjp3ncJieyP/AK1NMH+tQaaVzQZ1OowrMfH1+0VOTMGs5mmauxtyeK/V6tEUxnDA2nm62
E88u6Idd2BkGICFVf1+4uO0HIAv1P3jvRGNoZ+p+oagQqxpvwKvykSEQFyQUklBnJnyd4ANC0Bht
7+4VCLKMS2q0CxXmhblNJ6gcOTFcfgpe8iLgD4BW9lWcBOFJOlzJp1ipfzSqUFxHDd63B8vdDePp
Se3xjOuhYoAeW1zsY0t4GPss9XjBr+5UqlzHQf7lGWR4ZAHZLfXA49C+ux/p2NUulKvo2+VWYL8w
ZuImQUECNsD3WAT78vThVUMzrSTT+BTtruvoBrmGad0/zAMFMbXYYwa3SqwY2mor9xs9IrfhpLPY
VJd9npQsR+9CDCqrZ1m67+Lbz7B+zn7doqVv/80iNNEH+tC2If+wphzctu4il0O085gMFAIlO4Ft
XPFgRzFsqAlzkXCoYs7ic+t5UcS8sM13bylwylsO2WFy65qKnVPjKN4e0PfEm15lAcr+pOt9KLSq
auaJh8K7o4n4irYsIi4JxEPIkQLrvXRcX/cpWXZoVbyzFr/qmxpCX1u5rJxfxtxFP4ujPVC+PqRi
0ouDhXwsSQEtiSh2XGmJTDqfMuFYdcA0SvFOT9zLiuEBepLWe7iYNt8MkKXxoTG7HjDuhzTCuSiu
7lkINpCBL4FHu1Y89nH99pdW4HYfVPPu/o6dw2motr70kcvchimttwgN9QTlWI2luiqT/7YX0Hm3
1CDkw4COOATJ8Hww8+LyiCx0QnwGaNPTcZ3Ox6i5sE83dxekMB4CIZppr4vv6BN833m+K7R5xUlr
xDFJetxSNXZ2dwFuul59YrFIHVFb+qCTALCZm20YIlCU34GT/OrHmxiSF91BWTgMQgl11CJpiXbJ
rNhh2/fNV4nXgUztMl8F/ppbu8RTccqhJTPNypq1cJqyZlEcSNZwhFd2+q7cxoa18YxHfQRe6Gei
ks/GJwcK1XaeSIqe/LskFqeXyUc4CARMm7uyJgvlS5kERiuJOQgkZTzesjdTkRd8ampS3QzPEumq
wfDYElgxSom476YtrAfYHEB5zdXcwfJ5Q2fBxtEftsHYOLCCpRCnGu+rgtaO+60LfdqOIn3dI2dh
dVMKA0laPfOPWSi2uibRMip0opIbL63ACgDE01VQgVyhn57loMLmDUKxjbcKu8fYwEb6+cYJiKiS
oF5wFpjt3Jr2MdJfTnXSKgp6PlvyZbF+lSgRckSBCKVcfHWWSAvcY7nY8IuDePo8/AL4IFVNDpDC
kkbPg2zOYr9NG4u7QmfXB79wnGm5FOGJJQqfvIgd4QluiXMSIxxOxe76C4t4dQazJ/rnlFlyUUmV
1s7gaGn3nUtjTlHNUTYiKyOsXo5wkz/JacwihdClvwae5HfOkpLdHCIQwcpMIcCPTRaGOrl1kU4a
aI2o7g3431mGF1cc6mG17msyqG6G8BUAyNPpJ24UQSoM/FOb+XTJjH9nyFRcHro4Saq6n3hrAEno
v9jWyAQgcqdhRi2+E7qrC1QkjHQFB+bhOgMdRgTYXhSqqSml5lw5k9vci0n+Oh/wnrkwZQ9Hy/eV
sYIKhJSjosGQhdUiH5RZjnNLH8ORiJmBUS+2tmbaLQ4STONo+MRcI2s9MDSclxQyThYLJoiGsgmi
JS9geu4qZ+hHUNhS2j9ohWjypHjQ6GdtxSfJ3PmD1bzOdalMXkawhgmzpb6tB4H1f4sMl7J9vnwE
+zqhgSuV80VIV46pjD10mSDysJnv9az8udSdHaRXMP/4KW+0WhoPkmp+9wzJd86NHXGiZ/gcwPo+
ZFwDSK3RwdrPGfaBeJo+EP58dBrR/8osG17cLA8ozJP/72APzcVDBg1tB9PB2ahRdUumu84dbkZW
GJkaF95FqjiUvea4MdstIjY1CMfOdn8Sek/3PJgod0eNR4Rlr5zp2Lcljj+St3KYeALQiJPVfQDQ
c0b3bbHoYbkoAShXGD4mpAWrD3cC4klrgaLnj6QFwg+HpxvHxcvxC+KzXuIB2WFOIR5cByVJLIRb
oDEG9rL9LYUIkNCufWXHldmvld2ruxsxgoda6EwE0DTKwFbiSXxJAbbFTH7PM+Q7tFsB1NdD8m1t
ngY7XeWXrPRF1GPO3IwlIlpjCWCxqNNoc+OQdUGpHD7geJz0fvJmTBIoTM0zjatq+Z12v6O9/C0B
vrpdfwNWcMS+7tJemBR9h0YUHCGwBArXBPwbFne/FC0SoWd3wahkygeaKlRVR7HPECqcbtmmByQn
QkCVI9Lab2XWRZIXW2HBfyx5PYdjUuHz2sNGEh/7H8qFlFMSdO30mBAk+Aa6+p3yRhJqMxYAMa+p
eU9dpKSMx/7p7sH9SNt3URIvU9vSoyWqmbAGZYhJ4EeOHwxQujzfNGD2m9Hl7XnPiMRuxuCOWTsL
t/dzwwgnsrnA0Iff+hPkY8KqGebq2fB2hhhHLfyGj9Pft2j7UH1msH4KgTt6IxQ8qzSEQsy/J9Ld
ke3Kii8MsQgUi3Qn4VGdqLcu+Mbs6KJOrkwX/+i43RbH0+JlY0FSmcEeSn5PJl997sLVeeyeOYNJ
0Tk5Z5Cn4g+3JM7Y52rtIyBoVGwISYfyV4KpCeTVlge3rCd0PKgwWX7gLqSyn2iZviVkzpHYS0x1
DB62DVwPA46LCNSmbRTr+ptWMagYCyJikypOWBmT/YjBG1SoBmOTYfcyMHtxnMImXobdL0gNO86u
Gw/I/6GA534/XQAIEGiDjc1G8KBPrKXgQOoycydyHpbODB8GYW+fRGcWjR75ym7iD57iZNP+MTQo
Sw7phe66iqsh9Jpj1fYAT9fWomJV7zp3x/hyCSxi5xEadheTeL0b2IFI+AW4h7K5Us6XbCONhRE6
ouJvo+OQfnf6yG7WJ/Bs0YWUVZL+8rSYjkZ2l+ZuByskjdZ2+iqJQ0mckZAif87GST5uMCps6Es8
P0u5HPQIVc8J4IDvk9PaqnOpq5qnRA1xw7y9yCvmKEaoNZkx6yt/B8gGrhaybTAfFttDo+meglyw
xcGFcXWAVEphRt9UqrQAKB7Bc4DNh3zJesKBqfasmGe2YsvbpINDlo4uFiCP3hC33ft48HD4fOL3
n5YPXhcVY93uv09uUUYR97Fq6IyRB3mEOY4dGYd74/JNaK/Hm16aoJM9PM7qGgw5EgIgVO7jQvbR
D3hBAYl/MosZ6BrUanOCAa/viOtMlt2nl5ZCrZ4fAwliKichjjPmFNGUq2BS5Q6yQvG8sDzbPyVF
cSQRZlmc553GtRWvr5GKo2i//Nufrp7CSzrzWioGi5T/K+KihIwWmFxVMR8Q1YFty7iL7LuHlsMW
4BMLt1vWCxb4PpYQLpXz5yquudkCd9NPom0pL7/M5dctw1Drdhc7qafDkNcwzaZuwvNtNy8D1qrO
JXXQIWEevz7MM0oJWJ73Wtp2CkA7jmLhLRMPVju1bPnPZhLh7HuyeP8yxANkCeGaHh6mQLoUm9R1
4Dg/9IfiBE8HCzw2xV9q1D6+8mOwd3T1AHOaDGOhABOYvY7l7jLacp0adIS3Pyv2pue6QKHzOH9b
iHzssYT08mmiuUH1wKWvfjXhlWYSvyboj/N36059AI/Lr2yDhaNoCEYw33BYrhg3t9JkQezGIx+L
VCbbEwoxMLMXhFLGGqkGPnf5MSC/WGkKnr5DpyU8H5sfJmESyXUGLsPpwh/620MhsuJdICjN/po7
PthtdHw3YRXy3hmBTAgs9XnTysUmX0K6rCPPx/08PLOQM3oVeNiUbhXTixgslnhPWK7qSAtHtAd8
0+O/1Ru6/wIgDFSVt54Ixpz+Xn5srPsaBVbVEAiD8TkYfogw23n96hUk8f5SRKkMG7cTO7MPtK0j
ZTSoFFIWTPpXEUa/ucQ7Te29SZcMEQMSg9Z8TacQOt5/gSecWBN7W6reOG6uEpwqx43yhieMaurx
mUlCEB9T5CsFJVcHoFuTWORC4uaY3pjvRWf1WvOLNmzwyZgDgrv7CUdnuRc2MPFR8d0Dwu4d0Psl
hqg9yODz428gXspqDkHrsYmNlL9s3+zZaWcIQVFxeigCDybGt9UPFUU4X0nEWpDIsukd9opJTmFv
Ns9W8LaX0aoQDC8UoF/uBWDam2x5IdKuyvvaml1XAduReNEs9wJxQbT9tBJIkWCqouXPOAcsBrb6
wJrA7d/mXmmSD9rmOGxotMsf1iWIHxoHwDJHStXCaX1REW16vVijgapyI36LKU57qY+7c6oxIETi
U/Lcubyojs+Kygs7Rcln7JpjSaBBZLSa+d1y2zKCTPvDcQRkzVwYjoDiz5igS9hmSmzEPGphu9Fx
peXJQAz4yBKm0YKgbrh6SxizMWd8XERiHDrfhNh25TUFs63rvcD9QADnC+T4G424vGD3dPB1QB/e
tknZ6WC6cmyZ0KNrfR28koshqYV8hAKLm4u/r1SBugdiS38Iku74Nfw4GAccY9GpNEOkfmTy5kIB
5JTLytsf5ZqoBunSprVUY6STJsIFfdJ+4l0s5cvNliTt7XyAi3iH3jlXgxoAkHO0GR9nGcY5tTpL
mPGYEin+Wr0iR+npt8PLYXLnTbbiszjZRxnTHv3JF6HawjjqOhEhz9g7VGLcmSsxIBL4pgfvGvVL
e9+nkjFHghFBlI5aHApiGrvC5nNvuAx9R+W7xzgIyz/Kgvv32YeKjZeLMQtfAvWflR1QAlDgt1ki
KNyYgEivymPX7SPIev3Pk6BKMRZ3Y3z7TjiXSzgRQd/JsAnOgiTAfFglFF1I6vQ9MQbMoL7e4X6V
yfvBOvqw/nm6uPmPRrf3PKOfOz1BvgZ2MZZnoT+6+09oVKyZoPHVPfx8CmlHco6h/xGOyE/44LYN
tpRugrec5sIbNra6S/ogda++OrQVZmBKFYGD/qWVnZbopCXDkADCCwwKng9fX3uyQACuRb0TSmgx
AuiWV0tw825Z6MqmvktQifWCuMU0JoPbhX7/w1z1tF8NvDGJxC48JQ+qa1UEgoruTg1bPJnR7sj7
Q6d76Z3cCVqAnQqm0Hmo7fEky0X1+8ggGeHLlHHgpxqtFiwSTAE8jPIFXSz6+zq+tDcpQy2DTQN3
QOD0wotaZ4fSDiL1wrXRrVw11EBC8iyYoPyNvmpDV7bIGNPhla5L8FDAfg3Lu0s/6F6m/ZATXTlE
Rs9SSoiLkQmNSAqxK/J8i8z7fCSpP13Z4U3AWH9IWltBK1NcWWLQuNiJ8Rs5BxeYFyo32MV5b3s2
/ykRv1oaVxos8H3/Yk9YhwKPKvMjr7yWXd4ZX09aHC0qkV1nM9y/fuZhSfykEI+kb6k5bQke099J
qt7v49IWPupUImr3vEvOBQW2P+VKsr0xEaACcxiNEdzaR41uYZWSCKSO/mjA1aeOJo2/OTB0f7Df
AoFL5tV5HNrclZHwz0rpEfzkD5FgJpzmRe3yjSo3QKh3cYJCT+VCFoaXtS9Q9oiydIO99Frg3bBe
Ca0C0uw2ReSyuisjrXGtBQVzj1ehlh4jtnRcEahTMbHkVgoGjXRXM4bTvuClN8szMPivkwJE4XFM
1Aq+Sl3W4Xwf20vCw2pfdy+aIYGJjFcB5slt7cocA+yWDTbalEFcw7qRLywfXTFjHQNeyCbGCa/2
hcK07vFB95c+cxD8NX0thIc6t9Xgv45IwpR+haSWbZ3uWnfqvsq6uxa9mUO0aKmmYcCvw+MOfbTu
FnlGOfm9lMYR7NtCtdRGIZ96ksHk3FwoWhqkyFM72tNy+G79Hu/HozmM4m2l3kQwGWHyvZi7sI4Z
wge2VYwWv0cB8d1gu3LfDbqkWOErccXgEzg/1sF6ZSHFhU8MjLqE8BGf7F1oC3n5Vdyiy1ksP78S
ochgfaRmM/DnvMOkO3F50oLBJtOK1uKEI5SWw+i7K6pMreQfuab8NHSmELxgqtFZtbGTq7cUVVty
GoAOgQHADGF8VGjgnfAZA3BsJ6Yawqu+4VpSE9nGHtPkQ+PKtT2cuQQMnW4ML2x3vx82fLtcucHC
zh8eP4Kr35ujiFf1mFt59KnifEVV21xXPq7HiJD3gaVRkM/swbdRm7cncJyjsNyJrP6cthuU49Tw
wE+tCZy1T3zIPDIb9pYc9FeFAA6tKkh18fLtmP1JmN/lPETlKON842y3W0dIGbn0sG+Zkr/nmaTV
zhz/+667/SsYrlWIXKd+zau69SXCtqwjGKsLbUGogf2oqHHzVuG5/QlWzdyUkvh7gtyD0aBAx90Y
Ktj1xWjcawIkEr3cVkNMUXz1+vlrQSL0ZFaWPAM7Td5nFPia5al6+GUB+OIxdhb4UjrzH6a7grt+
lAGn+llYxq0/4t9zbYD8giAy4N1eDpl+waBRZBvYuY/nRqvga5W4XdD4ha8UwFA6jexLvtlxghKs
Z1+o+NDz9SsTzNdOsFx8pIaZiJRvRZn0CKNsS3gPeW8JU5VgA4Mj9G0JXzWeWHdAQOs3UMFuZyIN
pbrKtcitAqHA3YitpS7F0lughYyU4DS+ASmybwb5DI45zZOxvna0NrM/935NrhExbzRuIlty9MGz
VqJjYs2Oiqk2ovywuOytGhvYJaU70uuBMDeM7TPXSCHGLpOr77ACDXfNh30xRh2Poneza+5fJveU
tKtb60bT39zNA6mbbfY4fpBnQVVFyR7xv6sKL/KH1SsRR726Fs83G2LkCeEaXvBNXbhXBSnBXEAs
arM7WysKRAV5mVdGloLIoF5hD447+v1Bmo2unzCg8TZRtUttkj27uqF22mU0eT0dIrW5ik96h2DN
q42268v2nN1RoHOYlIsS0+pfRfQ4RQw4nsqh5ToNLylK1sPeUQG2X4IUWp6IOw0IUNxtR2/4q+iD
zQsCYy8Yc4B2jxkXll7oS1zIeB39pcTGmrgK02MpK1UY3FDeQCLcxm23grPs0RAw6bSTXqzf2B4Q
I0RD1sA8+3NaUjo5nhfD8HaPvWtpqpQW2BgwSoqwk6m2je2PU77i2ArSXGoCE7ACf3y+EMODObPf
sk4hm2WavUnJBKKY7fa5XpXrxp+RtRR0yLgrRbelH4QhwCY2fuRma/WlNFcYFJc8bJsIyt3GDSRy
2mvtVvhs7qzNB1i3/BkjIrKBGr0UQKYX/3Y0Rzp5qs1+wg+0iesVOihrfmHshX4uHbrxxmk5Ltg6
Hg6LcNPBbL0u2CZnzVBFORkKCOeQct1cfqsQASTXJYQqSwDFLC8+t7RegS1HSKXvv2uTGmlt2fEv
uLzT06i4eDMHMQeHK2yWwZkUPt0AelnPjY6rMCTVukuroHfLzqTltDn/lIwgbss4M2rZjn29nufG
OEn/sriQYWQpYCdi0RHmmuMRZVCBMX+ZixKeeHOYXmbFV950l0or0jgyZ+R2wyhOR6Rs49PYykcP
Crbu4/ONk18vY+nB5MoMy0sIkL5SuJHJRysDly5YcSOV1nkfqPp0NGDSUlg0QyjOwEjTJDb7q/Pv
Gj+tKXl2UuDlpFkT6BAdfQwe0/go/WT0d/lc0hnZ5NuufhfFwyN9UdLrLR91Pef+UpvW0C4GiTum
AdPUFm3Ew9eh7Fou1O/2eJBuee3kJe6bplXodXzmFE9nCFCLgJwoCyoI6YbUvpg2TaNkLmOZfWYJ
1443LJESPTGRUGcrXfAPlcu0Zy9v7Azm8ansSilrwZbT+s4dCC86CwjSPL6H4smL8Jx9X0AJVFtJ
hTL+8hG8B7Kjjg9TImV223EaAPZgiy71uW+ai642m8pnBMwRnj+ljIrVac2M1G3rQXlrxKjA77E1
Gm3bZV/Ho2BZEXAYpElqoJifArm6KA/+Uiw1TGs5letwwSQfQb7Rd+DnMQLCj0qm5LT5jtz8GLJA
Axq6+7YJoVeOzJWQuDHV/2dH8GNTLsRp7PEakbFCBOZ8++WhhdCzvfDEdElfiIGaGTFjCsFhnM6E
DPdOZ1oIUPyQntHExpaTRLMc/qRsNtjzpHKT4fFXiZiwhediHPbrYJQe0tJC9qbVlTaP5gt/a3pl
q07za9ylCOthV3xRYfvgRf10qM18DGTFis04s6uR8fgNZUaO67kw1wVUh1Ra4hz6BLNyQPtY49c5
+Bbt91Gbk0yE3sNWuwOXqJi2y9fDWGzHwZmWbEyM8RrOvms0AE/Oc5PWiHBuH6P4gY++oGbMNaRT
pvSAE6tlQPp0+z2V1tkCoVsCPkJN3jSjQPYzlRZAjpuNGxlPT4tS8TrrcDrNr32CG3ieAs7KGvAQ
TxBwE2Flq97PtXndvs/GgcuBb7eqXz1/hz2yTBKPjXgokmVhAD2QTZZeHlBjvxcsO0aMv1/F/D+S
EeLyPNQ7r88aKwYg7L1aOvfsnByzFdSkmUEp6tFRABJLFgKjUp0yI7DMG7GJZ/5gtas6auHWlls/
mTM0yPJOW8rFjwKqb0Id4fQR4hI5p9uHboeWRmkT+oB+mpRTdiE10AeXLanP2h/0Ruel2W2cO8RP
93OwDpWP1ADk6DO5cYN+aUosDYXwbgRoqgDIECiqP0weQuAdoraTgQ+HnA8ETojHtVYJx0g/2Va6
0AKF8k/8+CfIZktDMTqxR41xnCQNXfb8RURfGGSRNXe2UNS7jlgPYHM0eP4zB5jOGqwc62tuU03L
0Ht0tm7ym54v/75iqVf2ZCkjIROzKk2XOZGFuIRdnxeRTimdFMxZke71JGrtQ+dZKNZUTv3pWTH6
bRYi3CEZWMVpxxFmwxs1lumrLM1GyGQbzXeUD593bfMsrAJ/kl3R4O9ps9mZKeKaL1lxg5thlWnJ
V65LiRaDvIrb7TgRvWkZNlHW7X6Y7uDDpAgENHCHcRIkwTJ9At9bjOP8w4pczNWoFN+iVKsg2Qhg
iTiNcVwhRAWqjHzWyf1dOyQd0f9bO0eXyZ88Ieb4tyGKPhGP1HNZD0VuqXcLljXVIQgM/MsNsBW0
PHCzu26gsVlAj4mp1y3HQBCTTXxk0co6koMAnCxEu9eKR/aVagWz3WUUb+Aiuv7JyjkQ/S9ABTyL
6z5RBfUG/w0wJfPMVXXhXLH6iJZf2aw/78ipsfu0dh1E6yEXYs5aBwJYqHBzl3X3xLH4LyZsOzDb
mkADbCMp8K6yMF3MkOBJBoZbbf+PiIPepfCn/zjermHNm1eFkqLbejR4GHLMqNDVMtSZxfWtClEF
+RcFMyz6gfoplYz07Iy2QfPy2HrSRv2Re5cBRloU7m5hgBLv1+2rlpcVUilYebdE63kbqHi/9d87
/efrWLBPIBig1JtPk45MqJUhvBVSfcQVXU/+bdCVFGiKBNgILiPtg/sOQr1nUFEt0gjejTuccCxT
TCthoQPwNBKWKGZ0uWE8y7ITDi4b2pTz2sThsrsCWpeAjhC3xoRJhJU3oEmQ/F5Bz9NzTi2i7BK/
WcHIHodb8nO2ydlrRzZfW3Ff4jdt15OuIpLjpwX51GZW+SVL6hicOmam7qBdCHLHiFqjxt5XiD+h
ZcdB/NJP/50OM7AaHb/OOKzJuWDwSPEqW1j/khg9bCHl5tPRuLLKmGp+YJ3o9HKD0jH8nUJ8hnrt
vaIE62+JGlHiSTV0BR3S1UhDQUk42Gh6qPf/izVc9N8P/F0x4Nx2RMiwVmXa1RixsjUadCvQx/jM
i9kYNaC2X7zEndTFxyg7Gc6jnYRNN5IwQs/iBY7rd9vZgei6ixu3bEjvgVLoTjbICQm+S/RCyItF
/xuUuVFQQNIpLwCsKuT3DZxGd0eFIG38VH+qId8EcGbwOkAGfeRHTLYuedx5Czmol2z59g7/AomZ
VzgVCeo8pYynd/MFrj5TZo7FYBNMJC+iLLN9413ew7Ob8zj5VTXsqqY5NVPklK6p7q7++dtv0V67
+g2UUsfyeKLzW7NvpGKh5XKGUYgrvtJXYVpJyXmPyix1h2jS65afEhKOe7YWXZJgCWbVWDXsD+Mg
K5bY3f7zHty/uDZNyC31cbRmBTYquh4mF5WguhjnvQ0+S2AkX6XLDfkwn8OcnSNDXFLB8BJenGTz
kbl/0Od7AXIy6ikw6PcNjKd5xG5wse35KSGFSjFI8BIGY0bASXHtVJmyjDlcSzGHVeQJ9ez2XtgG
9DFB58zIxAdk90MC0awdzFST6jH2PqJcKmWvnGziVxaC4xV+/UI1T4eC96IXYwZEvGjgRtV+24P2
yVGiKG+ASwHdBjfdVR50hLjVP7iVGhkoUuM3KdzCo3axewippe545PJoQyb4FT8Yh/0GM5ijqkqB
1H3ttyIvjeqfhtNXqUT180zgGeUHRiC8jafooZ+vkJeUTpSwl8vxEIp5WdKyYVt2vli4pWxIEPHE
X3hENAE9EtjQHNz5dsDRlE3HpYDs2hU3V2gA/3lGhk3QrmNal9AUWI38GzNYuhlFP67unrpV9zSi
QVvjVQLXKUmj8gtm6apdTA8OZDCqmJ+biNvGt6P+KFcFdXbie4L8OFb4myi8YKjwLv4ad7ZTp1sZ
/Hn/EEdqBOlwYviWs2r3A8oUZ86dZxsRTmQN6CQZyRYH5Rtv5vWz+B3ZVEF3iPrQi2YD878iR2zy
NwH7wgad7+VH75+R6E62JtJ/w127niKgPwQ2p8TJreta2lqSgUXbJa3KHMnsOuT6W2hXkKNWLSR4
h7rNt2TEW3CKz0eMpwyFtWKnwxVjxLxwrnxbRF9HtsMbdrI/ojeIYTZ8cmsMxxObRbmIvaw6/+5W
xm9nm6X2i0F7c/pjByFKPtObPmbwsoceGXUxhVIcuuaL6DdXEDylMnpSNfb19HCddjkA5L8OfcKE
T6U2uLBug34STaZCqxFaeYETG5tKaUtTc2ODDI+VfgxXJrk1/8ouPXujWNr+pZk2/bCblostkJJv
PckThfgxt4mvTzgnYIAsKdH0bsNftD0RMlLHZRFI9jnvXILxrlscdWZ7Hv77UeZenbE2xnc9sRVr
hX3lFGjw/x2zaCqbv6UN9Oy7EidiQrhg9ZRGDsaGmkwyxMy+uSHQvsqQKPBOy3sFih8x6BEbraqJ
VnXOwKg4gKPZgy7hu+5x8/D6ug2JOgmoTw4Syf0XfaYFbfvSbhEprhrdVIKi1vtiy6shQmEp/DIO
4jYlGBTGHy+PlavdXVYiVmafZ8sig08fgjYrY8svdYxlsLrY5q4ACs3Vh5hGJur0Gkis6cjTKfCf
L4k5UgaljKFq2AmUPYvtSzAPR040r679z2GlUE1V5E8Wfpkmuhjv70UFN1frWBgEAsuGu5SPqP2Q
biK+0wtqSsu/dfNKBUzblKQUtHLk1PCTiVO6eu4mo/dgV5jcP4QII+H2tDA8HRRX1pEs/qm/pXe/
0UnyEutpUsv2BJMI4Dr81rR+AtNkxuKkX+mcwcANZM2DznafGqPjMrT+zir6Rji23TcuztsZPHpy
mUfBraeKsZjzPo4Y9N77vC1QKanSBtgdp2K9N1CmRM4FbanIr5sbRZ1RdMEpXTt5IMLYr1w8ou2m
HPIJEbeok8ZtDFBf7BiGz3Be+zKpbnoOVL5t6dPZE6veUqOYywePUK8aPrk4Azk4KtNWKFpttZTN
rwvBy0dpL64isdnULf8eHNjSlLCF/mapiH+ryrFxzMlDYkoxayfA9vnCAp/C9najkLAP22J10N86
D1m7dmm5oEobxFe5UawP5AvDpaOB6/AaWTJSQxllgDASrSvn38mo9xVAMgoNaBdJMEpbGr+gw8S2
faMcOGRq7fRRtfyB6EfaIoi3EbgtLZILuGZTTsheuLAe8Q7+Gvr0pjdEJh3ew0YI8qTLTHswPNyW
JHzK/sTwrg4gh5mx/TaEcn8iAx/waGTt+SUxHfVGWbfeGpXcUaqyRdKz56Sc/tlF8svGIUDcplzb
FtWTO4Vw+u/9ozkO/1mtLelHeRAFt7pWEnHNtMGi8h04aDYSOhSZegaY7HmK81T9HGnHOj45mker
vJBfhjwTZ/c+yWOABThoKRsVJz3v8YwUUFyWnc5s9OjAPP59hf0djfzq38J9PpjuAEpATXucOJRJ
EIThmAozLQ5EeAnNSlaih3fEtB9QoPHahI4IDVlQlDFDleQK8zO5ZXoGMxLBt1xxmM/VTv/1iyun
IGioj9l8RFw0nlriFzVrh0oORSn7TWlzVBboc2L2V8UNk/qkSLlJb/cHLuKmTVcBDqeWmeDz+Emn
h9IjLKX1ln7gxSQBQmbCMFolkyBimZKgVcDmqrSOioR9oiETX2IImQorVhpj66NWxavyrFkASKl0
cKlCVwNPpEpg8+lFGMpmX2Es2RLeyhcgZ6kZaHjbahEwNujESm0bQUV7Q0Hmi6a6HEHjDn3Wrapj
o0sd79eEbGA13PVNHqkLYhtlJf4ZlcaYbKLa36RuHx+mTYaaA9+IKLy85rCU8PAXSwzVa5F0Q/ad
QS8zb9TdjamklxmgkmzwznD/wE57N9lpP//6xAK5Ttpe7ScaaIj7ocZmCJ8y5kJOJXh55aetzXhw
mvAnxTGxU+dgtPd7eyBSiHGyXNlqWBNOpgwU9cbfsKUne8gfYQydWzrO39LtVVtEMV330HNgGMn0
ZZEXFApbzwuGmca0p1apAfyehfZqzCc5iaacaM1CHO5ZhsE9zFZYw/swgCJSt+kRfIZssDze0vLg
/6+EBZZWSI+OYwwkp24u2ViMc8ssxPld/tDg1GIEqk764zVKzexCWnw3Rx6eBQQTj1J8rspN482W
M06n8RbJ10NCnIJ05Gk/O5lV6nYy7+ipGqZ0vY4WU21Mkoj8mcBjRWcnMCWnlPCTx8cJTYxzLAx7
2+5VShbafcxG0NS6TNPUrnouT18uXeFEkuEROd+eRKhhhxep6HQ4tUvJEkzvKUSrU5dY0pst7bD3
XLY4uLdH/rjhz/SlBk8BB4F/Y4U/gONuI9SJWnoq51e9R39/BYHSS3GC9NY5sUS6jypU1vxHawgV
9cOcnh+ghoIztxySH2J9I1epNMO4UR0xrzwldF+e4MmOLPC+fhhfYNWXS636YmSPIRmHSYc0LDrc
za2F2FAv8KMIFesB0oCWRs8gkDodMewhhdobkGPZJ71jDVvr4sz7bW4gvHt6ocyBmZpukO8vpVNu
DnfjshatknCfo6gC/mC4PK6azzKZaqkRzmNFdocfFqE+/lU8skIIm9HBp07C4z1Vrv24tNkCbeJ5
R2jJ4G4oUKnQZ7M4y6GtHL2ynDdaFCBKV3uV2mlDDQTU3pGqh4mnqu2iAN3jLf5ndEorb+0N2YEs
LCQUqwc3OBQFN7QPrw2TCWNbS+AzSMK6zMeXdGHTf1sL0YzRXznUXBm+xqAPbOnVksFhgDh4jQZe
omdpnSPvqg2VY2a64AYrHUpBfpitlkIREOQuuhMI/Cz951mdYNSbqoVuTltQ0afgkbKK7pa2C8Hg
iY0WCgajJhYfZVMeGR9/LWIc78ieIRBUQKUA7X/pO86l1p7Jb9fjH6F2PFMxkjWNk0JSF1Kr3fRG
ESpjKlnfDjxkjSQYq/3xW4/id3veQ99lVzDMFwSx/+TwK78d7WNLuMSOuT1bFk1YVhDnLm6j0O6L
rbKnuF5Wyol/wu/EyLP2eCP0tFGDm3Upr2aXwrdNlnVysxzl87wsQ19Jc66N/caMuMCcQNW8qD7/
8Fc2NmwNIGk+ttftW3/bfLt0gEoI4oJrqgt83fBox5+0OHQwMQSkih+YkM1FqiML8x2ry8AzfHte
Mg23BqLl317RsPEA/siWBxUsILRej78kXfFfSGouVgDJ6V+pHd50V2BeQ95wkX+LT/LbA8ljMALf
tUHmljpjcTTrmLTdPQfTB0NFSp/6cqb8jigYGORm2BA9YNqvVIOJCtMEoDfJi92BUghIAcYWnSRF
n9wjY1a0rIBpKgMCKVJHppKKHxNYtO/2LeEUTjqYLn8Fp6LeQNNi0braQW9VNnWiUn0BBsCajvKi
oQCQgEcz+xmhZs5rEVVsYp+ltXqScLDadLzjG+tAPCayLptyPi99AKpl0rRSHnPowyZfx3K7RHMQ
rBEEjZKJsX16xzQ7gQ6czMf7YrMTL76ZJ9QcQCL5PEqfyFREW0+dxynuOlwaIk2X3amm2tMrRlV5
D0Q1CeqqDfZ1Qkd4l1ew+MAY/9liaMx8hJ0cPbaRUxIrkrrIcj9iVYRmoGrUVIJfXLyKY26bVA42
QfHID1qbqLklgvB6UexG9XMFjjS5J4AMnQKSZ4371BUgnwHU0eB5A1sE411eRMTPDf+KHzWBK/tY
L6cbjWdSKiTOUiV06bxf5OFri5pTXknUimwb0NOjwGu3HhTiBTHqUL8t3NNg6Y3N3UMWOc2BYwcW
mjxiFigsFy+jEy47jDzxRI0HZYpmiNCKqb6LH5Z9uc8czYiXeqWCPHXXtb3boOSKHIdVDvGtARTy
glmWHkTiFU3KmPAPOh3MnPnPAnxQDjG5oK3b3kzxAUb1KaMjVssCyjITykWkYBUh5T7WxmRbR0b9
GGy3YUz66n5bl3QnsWB2Fzu4XzM6E60Ske9wlm8Y1fU0FXZBKTetF5K2GQWZoBHjbZvHdMxJB9Yf
EqjA7cmkZgw42BZvRiFAEFcLWRXapvITunjPNlhSDhecqmCQwH/ryk9Pqwe0luNx4mA/wHBnfN9D
qXxG253HZtZ/OxiSkFxFl7VXG+AJBcrEXqAnCvDohLDnlmEg10UhYNzJHpcD6cybEK95GouPRIEF
WtN2ifJZype6dmtXFsiBfSDIXzexO/WeQ4rgXDoP1flGDvHF4ixBbmcM0lG078XiNUxEg1zntIDY
rFvTrPloixYRB/+shkoqRpeNoasVfItVwm1QzHxYJKqB1u9kNur2xqd/EXIIDBuhQ7ZOBDURdaK4
XPg9aiIlCFm7DakiCxo3Jbyd+j34yN9/5HLuQGTbcSjoonmnPdnNnwvXJQROdPzPoqzIQGzcX3au
g39h6/gWHtoYuT9UXS6kF8WxX1iPHUETTG27EcgQVaYJfZK2dhun84NtXNgzOQhD/EWyty6Exlrk
hQoy8MMGsOScuyI4glhX3AXhvezQHKWhPQwWWaA8IXB1IpGHxUG5eVZ2gsyR7eUXBqrjjBHJTRRL
bkcpu/rfoYTDsdTCUE+5hWTrLNGZQJ3e1GGwnKZB5G1vldsnOhv25KGb5dC7WED2KzheNoWYt4tv
ikAY44njHOHNpisjbfu15OnLfdSPqPGfV/BOEdUxMi8sD1/JAiVubS1HxXI863q1OnSH9/lS/6aW
OGLCIZmFud9TfQ5SL+OwUjkN2HXxsUEue86pz/g3R8/INA1GG3d0qxbRwgbvRZTDUCYhQu15hxhq
yGFH29bmyN/hxs9qliS7m2UjfgjQRDQ64ixPcSBTMl+izzAezv8i2NePzYtXgpoHZPHKKM3JTCQK
NRlcRk1+I376r8eFUHaxER3tEJ+n/ojOedH9OfRO3jhTWgSjPa9rTDyxbpP6QRr7WCdRYnIFHxJL
Oh++x3Pu1W9VakswGDqaHu9DnMfsxcT73QBE2Ftys9AInNTUW2BvRfwgMEK6w0M3WWdyLDdbbYmh
IXPzkg8f+NrrVcvUju40oh26pMp1RphGlbIOug7h3xO7pkDzIbzPJdxdVWTh+8fUExk68tQILEh7
LLGZSDuLtADYcu6+kUVyYVXNNUHMIfG3/TGJtGMof+vbc0b1yst/QfcXwCT6gwFFXynWKgv4dd7/
YlWGHfH8tNCZOd4oCEYjKLcsD5cZt6THbXq8Uke7Wf40+O+KaUsSBqkYMBm85vacVYqZT2bHdAct
tTjYhz5JKHs8FV1EQUhd3Wx+v75mcGrt+59ny0FLcILGV+ZFmcCxRXuzkLa4NcGY8posExga7Wi2
JECXnbuGlAkJtqjbnvYiS4tt22muVSTX3ZbhCTWODNlm8bblYEKPJOlIq+9lTDJ8kUDro1wOdo05
/SW+G5zTRrL4qC9kRirefQ++iZzaF9xFhzPpkQ10pihGgcA+w4uQ9KyizmA+KNZv29vAPk5ylLIf
58RA6I3X36HkpJ5FduWO0RfRMV1S/PrU8B/uXg/XmW6IFg7BQn62LwevO8UUEYMSKud0hsLR0bFm
PseGZKSSKoIcaF246utfeJDvfi9b9ACnvCD8AjB7r2zpbmFG8zrgvrER10cy1v+sktxCuAjdJoLp
rQ0GDdYh0wkC0xAcekFeO7l6iscHqUkW5p1qKrVO5WRgS0BNYlKyrLtkUpBiODylcWeyuEEmzMQK
5JHfYUWT2v5L+DUpSRd8FvbNzmodMK7ILx5+409xiYB8R75JlNhYfNDX3s2CbYZzewcsZ0Il32vl
LY2O5LDRiRMK2FWRPR9xB31pyYUoFCNcOycXwm5SS1OdHF3cBu0RYjXyAT9Ew4y4yRlzMTUcTurs
1LDg5/vt5+NCNNRlsoicmBzgsjV8ypwqimYLAWRtnsXwCmEZDgkQCMFF1AvANONnd+63Olpzfzed
PAk/S+JK4AR6gNJxZ42PLlyujC7ITOagQPQReb99qs141Ut5PTU+jJlBvGtTpy/Y41hx00kDoiB3
oMjh5fMDv7G0Tr4AJdasGQmC/xn84v1kJxoeo48pnXCoVCoHtxFqb2CngoNZlPGLYbANm9ichCf4
h1UDJknW/LWo06iKL/jAsSLb92Mb4lIJmKb+lvO1jsBzIV5sA3+1GL/xbQPkSZqGDI14U+lrgGBk
N+ysBLNZErztGSI/gnATwnHlv3lzuSUr/5C+AVx+4Y6xJXxrVMz+8ENRqYq60XRpXgONqClIFXuE
/syKpgDX2nhzkCEE1X0P1odCJN144AQ8I/vco8xj3tzYtwWst1Gz+AKMd7ROBLLa3dFk91BEOr7/
IKymSBF2FvOvSekLdpo35qInPrJPp+1A1GjorU7FUuBwoVGCZ8rAcL7fkPGBS7dvyWfo6hVGQxFr
ohlTUnhonQN6+A4GBgwkAi46TBIdib2Dirxq7N+SFQWWHKejx3uSN52Wn42rA4KpJtTOG3xqwgJX
ZbnDpOn+Fkrm/ZbbsZtwyxrcEqOLWrh9QZSjZTGupVdo8vE6VIFu09t82io91+exkmpyK6j7ozYn
dHiTlSVoBTOXi7SC44XPJHif5aAhPLef6s631PRbAbC4fbu2PysD8Yp3hN4yyEaqodBfow36SiTe
ay4ckLjJ8QYOdXoKirbgEDftWpYxe9scIMSaTObnxt4aO2pnOpjMm8sEdmetgwUjobebNJpUbUz9
HJjnOeNl3EROU0rj+bXwMa8LFItCxOXoSGK5zS43qqz+13+oeB+9gaUxpd2mSFY4/BzVxrs/fW1u
wISjLhx0wrffDj3PojM7TZ/PmNySoNHOpKmRnavRPx2PWviVSpDStohDwp/F+P/UoIXgQy9FSZFM
syI2fVocdphOLCK9l0JNGVFE1kYx8KlOST8mJYHPDMj+ap56ECRlk8N1/pTW7f7jOwcQ5IIVHssu
bLGTbn2ldr1yjtGyIWQXzN5oT62HnqiEmaEwMArw+uJj5Huk7x5pqNXSup6o/HZWcaUBulw1uguF
qay1LkFXh7LNlFDfto9JINnxg5t1vn0sz4S+f9Siio+iM1+54z+49SFWsUdqKx+6CGTX0QD6/uuC
8N6OZvcfhiMj9yBSJWbmjntiOhI7wno3L/dojBYbd+W7NuFqN9RbyR5/bETSMgk9+B+zoNdg9KTz
3cL9iRPj9HWF2k5iPlgMme+NwCapqa/pF0GZ98+GnCsFibxAJXrQA3sPLuslWhytOZJsv34l+UOV
N3fplvszGznjkyceNETJzaAUbsmVLhcCbCdJkWri/sNzCOckmH/njLNASqjU6iBa8kEBBxpp0t0p
JC6aU7wktjcg6AHofc3QiSTGGo3yU9ABw/ZU++cKeBrZgw1A8oLfzjOPqUbtkN3KR7P7If6lthSz
8gKaUbqzO6yuQrVxVuYHGUJX9XGDeAffG7I4iCa99bGkYR4TsjVHHJrAN5KgxbtHVJVQUMlBqDc7
aASCuo8ylw/Esqvhhz1K+cot9Obwr0XIEXhew4d/Bl5XdgPwzutvzLiqeVz7iKX4i4YyY6YmrtfG
WahsRviJiQ2V7lpgK9DZ55g7creKFuoJpDpZDbUA9qYJXlFHNScNNH/O7BCAaiU5a1UH2V2lf7OK
RWhIO1k0u0TuFu+5SuT7M6E0HNfDGuTtX3LM13kG1W5N9p7xGAiUayYQul526MfK1uQQvX40cSWy
31INCZCGsOvODa883S01yDrDaYaiQggVI1oIxcHOu4Kptbov+rIg6TJD1mT7hoLoY5iWKZXDaJAs
OLoMC1IpmQvvM0r1/nklP0Gz8+e33QUiVA8ujDjr3xJso+nVXHc8Vqw/eavtCYEOxWPP9AckYCf2
enDaMCxy7C/szNm0r6qx6D2IazKFUf531vt1y79eQuclb/EfCF81xLUDTL1UXA9KZuge/Dq60bgh
RJn0T0JEO+AvKfWTq/I8JV1Oo0t03gRiiBGBupwBqDm3d1+YVF+G+75zm6UzGRVf5Cr+W7SkxUMw
+Aur5A62wNzuRf8dNybDOLxRi4JJ9PoLS86BCDbB5lIsk7D9Ua9h3D3hQNTwXb0FVAQnU061y5ua
ExnOs7/ebzNg3vlrmoIEon/KouqfX7WjNcHYfs6PWkFfdgQNI1TaQPOAVLF9j4a8jo6xsjNU+J80
80W56yTjzFPHes5JPzmpwlc4bVA/Ubs/5DssmIwPj8S5IOhi8r1dvNj23ZxE30tu9OdfVfEukg4c
dd365QX8j+/VefsJAowquqHKOzZY2CDGiSUS35JkwZQpzq2Kq2ybhxmBJhGD9Qrtw9wYZbUmEhfk
k0bOxiOBRZIGbojlMWKW52aNJiY2vF6+Eig89lOLyS6FrG0yiXaVkgVVBcbFlpT21SzkFDZ+qG0k
LucBow19S+nYqj7UgA5ynTieJYpd+CdpTXqivy46u/ktwk23l8RrB7VGxPgFKO1PVQtQrM+WMAQe
7HiBYzzNs3X11KUlTD5svL10/t0RQZ4mH5N1SfpDoXuN4r7vsDGE2ZeMIdEcFxIovnQOULNqt/19
7U1IMugmAkVq73WbIolSE9qe1iQndc+r+vMQEJhAJc3ifeH4EsJbQcv7rkcNafPPYiIqLhlY2qCi
bLl6bMNQ98R14ghwuop0pIrG2QriGFOkbVBmJkfoufwRHoJ4NfgFtBqXGppmr9XX37NIKrN30bgx
OB+srVZIYBUTb40Lfll7j7H+t99oZLRNX+1fz8uBUC2L1smB1nRfz1ASSHPiN77a7FQhwhdSvC0O
IK20gB0+3X8iETXNKvtVgFR/TgqtBrgPNTf7mmkOBFLgEs3daLUCSil/KKbNZLgBj2HHSUKMJpxn
eMIsUv1z0s1k6izIIh78SQBnGUUs6OhmZHu00aODP9j7th8iGJrP/gK/wvFln0DRpnS/W2Fr+TyU
OpWjcPqA/mPoSwDMlB4K7IijAnYYkZjbNz9UPB0mxDXomGSIQ7frNlxMQUfN5bOpioi/UUyXjjWd
6cG2enuemkfFrlJG550oosDa9VG3LLocTsmFgQORKv3POA4FFvZWB1RwUrSATXJulOlV7lgRow8C
6+owHdfZkClNYgXxaXzkuxZ8+LPD+3v2cM0YJ2jvJ4wNSNQ3Yr6X4tiyB07lw/4w9KdgLEvm2MzG
kAbQFCCZdYtz+tULnDEWFYMxyw+VgmRqNDw9ds5Gjw1hFrtqyPDs27acloz76ZMU/Zq20WbNvlNF
xYGckISWrniaAyAtSl4cP0zHMHz3+uRmiZWIzbTP1Gk/+Vs1PzxwXgbRBYj8ifHdJ5EzNtx8MVcL
JkdXRmGFy6ElNptjPve1k9JC6XSbq+/QSkM5Rtdr2qadi4wlOzi0P2RHzi2VGWTWELKPJJwtPyf+
NaGluqc8fwumyT3BQ/RQ7e4e3TAAj6nIrK1eYNbTMP9eO9jBSGb4okUJQNnnfrnQPL9xS1Dnj6ls
2QvgsWONLecoGs167zE4ydvkdCRSwyJqLg1b+arj2FpIaaNuUoIvRtMCMm/u1Sw5waYWnXX8d+sY
XVlzylmT/jB1AZlo5xHiBTcu1/eRSXsCCK0QBtm0aOk5tu8R+Q1F1/rfv4xqL93IR37ckP2XRmDz
ezlWAp/l7gLTqzdYYx+1VNc7ZbzoT28e39L7dUHF+Ar5mZBNKsz69e/cJli2a4nEQ1GMqnnniNml
VzSSiP1eRvxXNZBLdFNitj8tZcWWMq9pa42US4LyhmzUjChkx2PhuqlYh6zER3XNb60qOemxDhwm
uw7y/XhbQFBS6MvD6shMFizZRQ1RLr56Xrmw3mqTOE8yaTFu79sQsCLGY1NsTVBy1tmcB5lWrq7W
J6XBOuE5BqPLgIAiwwHyQD9xknnk91+6sq77zEARDRqXUCrBJzzwaxlQKmk28QHymtJaBBhTeL+u
0LU+oF+wzar4h/RYKqvwbOHj2oYfBnRpLI951iRdtf8rZEx+bzRanvYG6uhlTWZDNovF2IH6wTxh
pbPLdLNVlTaqBLmNHeXQ3UE84E7ONwNPFkJR1f5MEdkPNEMTl2uxK9DSWkZcYpLr9cGbqZTwXtK8
uNRLX5MQNoMkM5CmItkjuvPyHRJQ0gBunpYPzZTZEbN1r03QU4C0EFOijxSHfvn21KNTcLy9vjnZ
SKMeMb+Tcolk7WGLE6ZC1x9t3gTm9ivbhGaRvugg/acu+fvf77AhH189rrS+L3KkKMRvztIGzyts
0/VUhc3RpLGtbwCfWoh/m24tRbwy4nPu46DG5UpC2OV/oNSCED+XZov3iUyk4f0tLqvWj2EpRELp
q6zpaLMDPJ+QO58QKDsSjrIS/rYd1QvC2gkyXxYOxB8xFOAkO2TWlznjqhnzRHlXOWQuzhxUyeYT
XII8MB3yDPGRHXkIItJUEjgdPTcILzo6aJeyWP1psZHA288mA8hvUC5AjgV6M9axLAHhTqud91tw
U2FE730OWm1i3wDDkV35xkcoIOrhJwdq9t5AexU9iMLVoao1Uz5ZDRSX5PEdDhRhX15VQSHwInJd
ekQBeojJi5kloB6FQy5dMoJ3AajTeQoiYVezA6IpOjZ2UmQETu80RoiSgfbMCRLkK9G++x5+a/T7
4lWuE/mEsnjdlEsZb+8Gz4buklnMmkWSJk4whbiZOyoGyz1cqjPDM+VkeYvBxiJnDYL0VsYlCcjU
oPs7YL7T/rKBbCgDukUPvG/gVPCbZ2hg/KOr4QbIFGg8cCaDrAJUnu0bQdftdE9SWYNsV1KUtRp7
HM6akqtpjuT1e/wxKtoX9A1Aom68DhiGtDWWZ0Qr82wDb0FidLCk4MmMBWGFNsZPhN9qyNd0L4oW
wCpxyf3GbABIkHnt+dXqz7QsJpeCNrlwhJUfo9JOKtxjYvaUy2TXDC0QU/qLB/8xHUJRe0dDQXkH
PDH+KRGGo4fJXUUa65GyDpQCYtVkL4SkBay4jX+C9xQ9UISYgfeuZS5is7YMVjlPjXFLayIJA/Xv
kNvAsnfnhZ1Xl1JqgIjIzQwIeB7kibTHzYK1I2Unw3Bvz+It3sXq4Kn3Y50qY+KkY7Wwh4/KbGrL
XwTnr2KPfSUs/aJuhSbFZX4Dl0gGPEShmTxfrhEFqzKydO7fXXHbAV4nIcu/GSjPAYIs2gVsaBKb
h/2dSCdbN9ghUyqJbuzpKt+jZk4tsLMFgk4JS5LwIe8jAevkgdNU9knKs1TleaDAWz3ZL3rxQU+J
Dx843TL199MkGgdTms3lmBofN14QeysB3rrniW+pdP0a2h3GxqIFvJEf39k1mUVGoiJ2OUlFc5GA
kCI/uQHt9nQM+kM1+vYaJ7T/oMRx1oHK+TMPnTPmQg1OsUmcwUhz8n/75jL8HVmSWtw1Joih9Se2
vbdttK6pgd0O6zeIpDLTRz+gLLwlJOdu+eJmO517wcRvqCZdgIlbbsVHAZzyZNWEuKS2c11PzUVF
gAaZxupxwCLW+f7SAqlZ7CEKE6z4d/I1DgVpQzrhyDGrUkKU9y/uzb6ADbndUXloPg+hlqsT1gol
kEQTNcGbAPY1u2dG8/oU5ZyR/fchM79eupqENsMUn6saEplrn3tJBvlUpTFg+sU0aEk9FFGVU965
h95KkGrxW03SYJkhOB+rKjJZPr8otkjEHI4NyKoHL3bE3dmqE7+mPy0dcCg/zvd7n6W7L7BVpsd6
l6PuJtZSIlHtJZWsaPJu2J8Zh+QMh2/dxpztgNdPz6/SDSBSHnnm2IieVkw/aN9ccNgV1WGD4/VK
+SNioap4Sx+/P+B8pkClLhHJBdgiL06mhk4p2ZzZCF3KK2NrEPeY/Gnr2CRjPRBLcKxwoT/xpqRa
ikh9MmW0nInGkPALMkuoMuG8UonWlXR21yo8a7RYDqv99NVfDqBPeRe8+7XoXsqpeeElSjcBuiK1
vUbYffvKLrE16yBCz9UdZKE506973k0cgwv2oE6j8lQmAx/4KgDw3QNfyjhO79eVqbpiM325/JI8
HTDAMwp/WmubGPiRUeRPWho326+4pY9wMDjCK2gVrufRPnmAMWSajaEio+N0C8ePOrkCuStv/LV5
yOKpF7CyoxHtI6KHfHGtcIPNv31lCZ46X0rxIa/pKiiWysZUxnPpgFetFsC0Vd1Vhs/XHijhqMbi
9RXLzzgBYHawvIx5vggTRtGTqCLsO1gc5ZwyyhE0JOFKWVbOupdInk3Yz3q6hzot3gY4ZLyErEFR
hqVkUNgYiU0EVKqXaGKOEAOyDWwTOAe4xohvOe8zZqk5Re7saetcLAos/ainfL8c3AJ/WmHhbgKt
XBt3EKnzYQhabgbIdajqgDRaG1RNYpAL5UjQkZw+Nn49Ei14vnqmFKaF3BXYocakePGxkDgN+owt
ql3mpfJGUoAZEXu2Ucw2KDgZqK7O/bPVsuLghTsfUeZ6HAhVRMJC9nhGJnomjgBsB048Hlb8e3qA
L0aMeHYovXoKq7psitEKmV0MBD86CeMyQFRn66domPocwD/wLojS+e66obhi3sq+W1iDL/uQ9XFl
lMTace4R+JEF5qNPrn6IYl3kiyy/31gMOyEHiVL8657ZegykWjRbVWdCoF7gBBFsSu9e/HAXXfLU
imVznzOshW+NjU8Bj182ZfDW8NF1AXl4rwxUNFe2CTdFM0MxzVnf9y0NYgdpzA5HkpoxIinPY2bP
kPD13x8dcClVoxhamLJzLoRSEHCKkeQJSchE+/OZ/1yY2FcBr5zQLB2p0+NcmHcHbQpHUUuyFMzh
pd+OABOjD5vWmt1TOMobyvbiYlUY6YjsILwMJKXcb3BmK0GYAkDHlclx4SFyJ9gKsVUhvITQv1H+
MJFNRyZDbLDqZX7rPwc1RQMDCmTOHjkbvpKC40t1yanu3J0Gw3aOP5EaYHG+a/Vb6TglJyPVelJL
aK2Kao2iOhcAZcQLdf99+NcNjIJydwvkctegQV9V6S7RpJldWURnkNU8iJ59597uGgSUX4VXJUY7
SrQyo6C52i0YqJpU2Kov6KryayF+hqxFTgxGD9rM0goixY74GZZWE52zb38T8nMqr9wnp5dEhKB6
NW3ti58wEG+GRWnV9uX8S6QBmeHR55blCgmnYzlPZdUSjcA06WVcQi2fJRgD/6/4ZWSMKmo93Pys
Ro3bfSCKh2Dt5JcyX5A5AR2b1xmo64ELqu3n2H9iT4yt6FgRUnz61Jlp3hWFknqPi3OnJ+yT5kKZ
hnq+zkDARIp7TxNCLLme1T5REFO60wOMIYxkRRAC6zlH/peqi3DC2nIwXp46AvGwX3WzI/OacAkQ
i3QhpAEkqtqEXD1aXy6M4I2CYOYGR2QY3jBSiin9r+h5n77CdXBr21UCLVNx5yC08lHVCmDcusf9
qvT3cYJpck8eNT7iuwzkPPKB1Rg55Z3aaWWZIpDj2Ff6lBu4mIGT+fGiksekQEDvrYQCxdnQZYho
mxYjicnz78CmRcAOWoZQko8b1Ls6VjDJk0EtV8tbV3XgH/7Z5r3JYYtKOywlLXWd34BAlgbidgMx
FJTuUgwI3wJtJ3PhsMXdOMNQspx2eROatCUT472txMfotlhsLX+NIDNy+ZTG7r9CO1hX5Ke83tca
ynm5goGKdrO6SfsFn0pkxzTQAUeDEMtyEDLy+SKyW+v1utHb/dC9YO6RPrvrbUFN+xeUuCFr6eHX
vkdnyDppxZ24sz599rYhV7e1bL+GVwPP+09ZNXtFXFZhUKE3ZaR/7I0qmOAUppe3H6jSHT4cdrek
OmVaL8UGGDU0XezFohLn0ulLuPFPk7u6YFlCZLPqytJPNv/d3CDbR6D6a9wxIHz77t0f7Gz6Qb+Q
mSBly/wHPPnBfdCfh502LKtFO7CydDaZmo3/5AnwN/eKS8IIguWzvPokhBokw55PoxeTouB5xWRp
R5McBAEcgAFu3kf+LB+zANAIA/5TN3DBpA8Qklw2HEd33/tsnZwOZstjGUziZPA44NQLTWpNgoVb
6pNQQBFIiKm3LWTmEpP6fhSGeooXBL7KGDD80HrDD+yctiR882B1dhgbeVAPMPcqOi1JEzz9QtGT
/YR/fvO81eC3sVGs4iiY/jUaqYj2DeQSQXnLsZ4vrDb9YtDs4dvcCDt2WApcw5lJyyL/Epwp5Pjz
yFpIi615ZkofullPsMqE3XTBolk0pSlPgtwi/JXQAgAyrbxgESYvXL+KjlqFn4CI0jS+W4ol5J9o
f7UCfUwUY9IhkY0QjI16XdnmKus7SLnIr6mB67Pmm8lT/Uv8Podnw5NQqiYb9xfBPOVc1EYs9ql1
fqN+fENcD71ZIGfFBcTaGlQ/H6NPJWwmHGx7MzlkCoN+ckwNN3Ed4Doj6dOpOUKJeNydcFURQgCp
UfeYC5sjvPEqu/44eqKxPccJWwvFGXWMoEImw83VEtn2SaPygVGA5rifx7difSJJpmy24kRTqLYx
jmlXa14cJmF8wMaRjw5zpQ3IPyK07KTkrIcYT2sgQkixDCnwYPPhSTB02dpCW9yQ1ilrlaeu1xmA
2GbtUzCZHrh30y1KB/PoiWO8EoHfkuW1w2EAiVZ1aCu48FJSmvGq0bCTxLvYUjoMJdZSlVFaAbJv
Q+z/TUYEijzJ1/jdHC+FVIZbinCSu9XrWO0qRQRYnfkFpmQStZ73YOBjj1NndMlssReBMtkhVlgX
rExPi0wSkTbDrS3kfeuNN6AH5sJGpBmKe1pslUDJuLMjazPD5yuFHNW1GpJEQ3tVEr5tk9mTtYMI
jcVovGVZMe9z2pq25Y6QB0iHvbb5/6FKew4hH1Y+bEUmmETGD4HWalt2UndQw/P8U+RQoYRKeOZo
rQTYCfb1Dcbpl4ea1nt1VMNdaZZV+XNFBK0sBCqiN9KBTAtC+Igj0TmCpSxokBaObs7714mANJDQ
44QN74ZQnKPilREIEcEhYFcbn8QFQcP+3O5CjFyUDsC0c3fxjJjgGraFkajNMZNDxjg4cIa+QaRS
5v/UE80s7ZnYc971UPa+fmrPZE5r/fofBSJKO0FLxv6atI2zK1cUwYLFKaEbBKZ6WgZCriXuhFlu
UcBeinW846e7tig5AWTH6qYao5vE33KjMZIuQxkl5tS2thWaAxfcnoGqZAAxuqRd3rPY9RuPYOVV
YpdG++Eln2AgUqFNo47HMLtmwFbQySolXfIrl/jkC6swkDZoNynj4GxY5V4nJbSLHvDC0h163Rlv
12FVXKlmhIny41oYjHwNgibKa+c6qpQIZpZlbUyRPs7KGA7ymvsWPzIe6sX6oA8kw85XwhZKnFKy
gJ578/tTbJMGrDG6vQaGkL0D0UEgVOUyWKBEZ7ecYD62FQTbrpXzdD/Fad65EVaR91WYUmL8QCT8
Qh8cU94NIectg+ZLzkBUGk/SJLOYdGTiLEvfK0b18a+1Uk6HMcZLD+SiYZkr94zl/k74VTtPRFiw
AG5gWKcsHP/6ar2JRZOcSokL4nuAno/F+CdoV1PlO2MzS5Aux2Zx/ArvWFPiNcVJ5MgHEG/bJCa2
MLZflh8dILmxodtlzMv6oWtf0+oHWT5nbHF0MeKvaC3A1q/baxbSFuu6W7O8eiIJBvvREGh35Img
WTHhSUxYzaV+xrkbxMWf6Eob+fnY/X84azSpBZ+LkfEVogY/2C38AakaxaIoM/vpIHfOKOFpbqbI
izSOuv6EvjTlR2eZqWn8JbcMKp96Kcp/ap0hbYj0jlSFHu4LcdlD/kGeab2QJQEqQepwj9WfRJFb
Sxqvf30xOH2FIcfzNEodO2WwaxFEtcyhhUTUAFp3ONHXilvejBmtbY6Bk7EeuhQ1qQzky1NLDjUg
fKBDUw6dByr5RotxcMpLYxkQ87n+W9yg6Gp/dPnORHvns2CO8S7Yshbng5rd8ZXlqAZTHyNmtixu
e0slcz96TcUVcTuQXEHSTPF3heKDF0XDLBMgSwYZDTplqXyp1Nqj1GpDb4zc0GK1eb3kp8XKbNXs
vgdLvgaVmN0chcV3EprmiLzp2OPknMvUw4cEWPersPAhmHRDbh7PyUWl1zD7tP5sSf3v/ysv5LHZ
fke5dqzO52fNZ7eSPkMM2miIVKiIesh47KMyC5/Y6pQna3Geo9+29YJ9nj8FyTCaKP/F3VOQAZpK
t11GWTAACbifIaIF6P8eaZeoiS37Y0LJffaHmJxuhC+Fc5nllLPQFeMbEZSM9gY2gWz6z5IQvzc9
Nai2DXrqhpoUMPhfuUOXgs4NHaOcRjIKPcjDGkTeYsw7kMbgrNPy4fj+NKBuuGFZCJ1ynLcB3ii5
0AR/ltGfE1H7fBSWVZU8GoyqaBOzLDH3ktc3x6t3e0O8oFvLn5xa2yo7BepClTKLJ9ia82OGCcvD
eeqgILaZkvgqCFk2jyQ/4zDTVLkscHw33Xz3I8kWQlB0wYE7it/sUTZIQbYdTEi1zE2HtUyqS3vD
6oBsFpzSyDxKRZBuu95URnuGGaHvOrfoehatwNO6s0Qcy3fK807plZW3jV6ZcE+5y4mWcgVzVawx
1BdsUiN4jX5+G19UAQcF6XtmKtQQC+x0Z6TPE3iZzY+YCkpMAMfbpQ4U4UUl0pSYDg/4WDs7p9l6
1QRIoZl2w+cgTZrhzBAMLNhtE9e5AkOb9nk1XCHV5Jxs3/AWO13xFxaP0hZUR/xNZg/P56ESrHMK
O9ctUfeRJdfbsfgCOY3d3cGlaMiOLPqT3SwCZhrnrKaATWyTpsblqdxIbyNAOwDwyWpQy40FBDFp
5nZWD6i1s0JxUyAJNd7eBgi/nIFdOJhSOYFcLOJllUWZkUXewveFxR4flybxtUxy6BxawnT7D3mj
affyG8aSu3BYZMNq3zkX0hDBD5T70KcJe9fOQ1rplCSfTiaAqQgwfQHFsUOHRGwPwbb8r2/ohdYs
HA8vvLw8IYdzICVM4/IgQJshNQ0YJ2SCqLrcTjZqwjwaaQJM+MIwl/2MR5PEEJp7bDMThRz+lJWn
HRvp87hvXFkya1WRsghT90+McpJS3PH/y+mzXSE3TQF5rDjw66qpxe+Rw8NPvxCOsLes/nBsSYmy
VLmwcKe+gLCMti/8NQDdw2tScsJ9DfazT5QvgMtkETdA/xZ8yW6Zi3enL6KAo38BNXxtEqmn4ti0
zHU+eS6vn5e1DEaNGphyUXNfKzivwi5aoz19buowaMNTcYmSuuLenvwVtWrnNEJVPfqEaaeMtNnn
QbMVq8/n9kwvY/vK5oETMYJRUeJ19NRR2h61g/d2cTu4MLtGv45LtFFwUAn6CMNHI8whDQ65VrsA
vDxM7Mpd9Rr6K5CuMI6XTXAH8pFUhbrI45eZmVqOMXbD35pqMyTgcrn0h0BgGgYwNpJlB/XP68G+
TlG0pQOmXoONrEjZcjHPm+lTPWv0k8DkfTcLG9ILrX07tWu/ujkO9TGtoehbP1DZoJJ46Eao+oJ3
Hih2TKH7OyJBFe4R+Kmw3WWQhkYuAhP2CKI3aqdKtkIKCFNmd8Fb2q0NafBQErgVqTEcsGZac2yu
XTfFu9Pjx0Zm3qM9y3sOxcUAMpjX9GYs+xwS2G8vXWrlhQ4Nu4GUPTeFTXuowdw4Q5cesLQcrqJF
uQMlQU4rLSF4qwD2dDzDWKwp63oTHXf2kqyBu+qzaaSRLLw/d3GFdtPiKePf2OAXWv6huxGvxgmB
Rpr5EM+z2F/CDKLtAyvKMoWvJCvsoMGT9cEodzQKaFbUbM0jyYpp89NQLYN5kkDQZUQh70F463SV
j1RzWEs2j02l1Le285TqqkuOcbmMjNT+eCAeWMafNndBrLGvHV5XVZndgFb87Nrfg3k0le9SpD+6
ZncAPyUxhgAQ+u/JYatZYUnOftLAxfip6BcMvZR3KeKw2LphKGBIjfGEBbPSNHWJ/yYtvdzShnl8
BQDqDK2VoQOntp9dP7vJ4qXHTW+XsnlDmh63HGVB+A7nu4JNJYdPm0YMEoJ1z9aiWMOvohRR3Qm8
VC8VoBz90oM5sEQMTKPZtKyv/yjmGfPBpPj1YVDhdA0J5ZvgWoU0rPezf3WklxcG7NW/aW7AHO34
m5uKoRbWbWiJvRbd1WS1aDFSfDcVLaL37bBMYFixuDSLnDv/53mz2N4yiwtPp8AO//lWdXAgXZJq
FE2Ie/25VPS5r+f2DlAy7uIBj/8wTNCB/oddnl2iB2a15Ri8rglsEi0U66xeKPfpebItZeOeVx9w
xtlGFyUo7DijbIk3ZpipK/1ray/3lXevIqit7FPjtezt3kK4gzpmfOJsPbaEIa4cvztXgiAczP6A
hUtT45wzj81NktuNjPb6zuqiQp55/024yDaductadsp+g5jvqfQd20Xt8gzS1QCiAKwY1TjYiO2V
AZp6Pailt0pOkNCMw2Ts7Re+mOE4PNdYuO2F2/IRBHFp0+ydI6I0Bag4TaF6JbZkm+BtsZAWgbz8
vQSyvZx9CF4Xpv5b9UuhS1cF/lJzQktrZ8qoOJYFuOGAeClr46Bu95M6IhIFTSnxKeHB0G9z9/lz
mLqfscYsQGObPtTmkJQQY2sblkfiuyAqWXw1WB1m1o6x+nRCh0VNCiJQ3j2UW5wZ/3mdih/o5jir
usePaq9RxLfD+ZD8nyj3X50iIkozzEeQoZ/A5Z2PS/S5YVyDkmXM2rrobRKkbWSnabZ4PQJEy9Ub
cKLz4njrOMunmG+yGXJgp3clmwZxGDpdnqT25QSPEEl7mwzrL+eJIauJuUR0Q79uFg8JLCgTozmp
fG5SZrRN/J/lZIQm3tHzpV5Vi46M+xvOp9sCqRqXca6Tbwxc7grcRvQozunpioNP6DImKeYsirzB
VnbrBxgidTYLo8Dd3hn2qtY/ach7UEP4wLwE7O6d3WR/Cwnt71yz+4jick4Y8g5z0laxhat0Bw/0
eJ6cLuDEZuoLILTK5vxCiTq3/FoWu/o9tY+E1UMfh9gREecm6aIUDVXt529BK0rdidmOsQNoL3nB
Nw1uVobFQxyfYEVtrfqoJqTVPwhB7nuk5GAqiV3n7mUI4l7Z0wyCu0Ukncjm7VNyxSAEJePFGt6E
MdBZ6LhBbSyC040Qtls+6yCXne7kRwYzgTqiAwiihQ+yoH8kXNjqjutfs7wDWtVCSP/UdMXAoJ+J
KBeRMTpZXMZ3HArnuxDZaH304FT7OEF2wjS8Qee4hnTEuT2PAKa0HQ1pi9KiZBzu9XGoBjyBPUa/
gWqGOuZXpAVVYdx8nSM4B/gapgO0mrthzzfMgpT+Bte4HDIJxmfmmNWRNmQsesFI5LvQ2PIUNjQd
F06zzeizi3wPHpUR8i827YckIC2pq0Fh2YLEs0Pi37uVgYpyL57HBB7ISKdSHWP3LzhWckDBOVhe
b565iEYxUR1w0hV5gbl3ssPV67fVyX0xaOwleSzhcUR6Geq396my8QPkl3faldLugWG4azP6FY73
UIv2p7LInmmA++yekG5T4DoTpRUoSQoZ36o8uYkUhqdKt7KiYdgU2EtRgX+jIt9zIUz/Iiqb7QK4
tSUMyKh5vmM+wQKbpqN6YWA+977gVdqZ/s2ruy7isgmTQ6k7P0Rehw+QJo2J3/9/ERCdP+jltSqH
vYaW6u5+5G1QwZkNqzDD0zKM0GD1NfOW27pLJqphLmdrWLmVOpqy1Nh4Z1zuRq4OuP5OdEF2QUha
+Ax8D6CCQ6yB1PoNZS99odJRW8nh1TtQzgf/Y+1S4VqbxLdFBN/sogOgMeAwtSp816pYNuKfng6w
2w4lk00EONykyHuTb0SKZMPk25ldzjK4rXz8TrBMkvaMX9immbsXpjSbLmFIw1ZYUajdDqZK/3Yl
RTZrusBgmy177r22nC5P27RLPg2jhTy+X1CokJpCQO8OVT4XCUohZrqQyfsx++CIzBpH/axUFgJs
m5Cy8C4hmDVf4jvqW1qG94asTyNT4HzGjjK205CLnsddD30D4irujycm+TUcQwNqZ1jIgsT3H+WI
xfwB0AgfFjWWZOLApGIFq/amzLFCnF9fVIIOm7uJwq5evDz+JDcvyv9WAJaLg4KqALnolU1pztxq
Y/mPfoNrYgb+yNYqM1wH37B/ILFPK/k1hl4TCPMA99FWSzayMiHTVacSCtQd2rx/HYL9NENzHjV3
WeHElk5IbS5Ca9UIqSiBqeucexTwRWNWPxI6bQp6yp0n2PrSgsqjNdOCU1djf9tQLvF8/218zbu6
UhvHa3G8NEEb5T5YC5x0L7MXcrmsl+gqN6SXltmUSkIWnpREOScxRdW7G/1hJRL9mJGPrvDsUAWw
Z4oOaOK/ZEz5W8NDN2pMe34/G+wEzBf2PLV77HfX7EFlZy34b74HPQJe1QkfAwCA1QEwMs9kKCKp
wFF1UkyQf4Tg8iKAgrwyk1SgoyaZW/J/aehYJbiBlwISgDrn1fb+TEpYfXKv5jvGu/8haxdHE1UL
rx2n6y2ZzRVMlLSM76ncFMDqlg0wfnh124cMG+gho7gtrGCJx3DOx7MlgguhLJ7WzDRnWJPgyOIZ
EyfCEUKK6nME/co9JSN1Xe9Q7PW5NB0TsiPMpjJOcYADpOHwlIfbOGJlsqde0GGhyIMQCnPcEEUX
XNRxTS06FbusD6GZg4bzNaqD31GggJt6uO6EM+5Uqwm4NTAeyreprv0ipCi5jfIfOtldfk+0MtHR
Be7enauADTHw002NuuYrYh9RwjrA8gaeDTLV6lnKx32Fnjf/NcCpSzMtRG2tvWrKuKS90vkYe0pV
NfXg4NsNroyRowv1EfiyRz9FPPPp7YtBRa3A0A/YeAzrN7JsLcA5T4v/3MQ588/gJEgs+ash5YlX
4dS8dWJNEwb3/ROxnf/j8xE6QSEo8qGGY0D6URse7f/PcH5iDGpLzykkLiohT9X+/ox3/DbZVRjQ
8ltDYuV5CJ441lXZ+SWgpV6EtASNbDb5OkcNmSKsrT4GgLNseN2fTsXbIU8EUbwOYctFpzUv5+pn
vGmYkkB78G1ajFI0LhxvJgHIHh/kvY3bY63TuI5mQ5+TjvxHFvidGSk57hoqPiDP+qX42nGw3tZH
7TU8t+FyVI/QUPmBL6IEwmohQlxZ7/JziFjdvhLCGl84dMWUwSHEH4IZwKmFPWv0pTKi7tnzcHQ/
lSZj5e6WZKJmXJnlXtzJ8b6402G3QNN8HpwWvc92LWnnPRNh4X+m4/+NxIBFtC7NgQWTDwKkMBE1
HPYkzlPC7sZWeAAUfKnTLOUpUPSPT8uVLhAN9eXu5jFrfqSNjGeKY/i3OsOdJRl2fWk7bZNcug4h
mOOLFMkO6BQDsRIWaR4uW7RD5T0eXHysod1BLLP9yAiiWTsj4n6vFcS990CLoVsCpoqrJP2eRpm6
L1FWclRaq9x1xjwAyEwjFtNGmR5GMCQx9V2loIytMqJBKCdrdl9s0sgQ4X6iF4DgjnIDxNgUeE5l
erPPnkQEqiP0wDrBFcNysVmyQtAT/B3tObudqHK72oksb2dXGNKMlaBzvo4F5T7C9R0+p1DjssB+
+Eb4n0OprgAh0ws/JcaHHs4YCiY7ELzMVS/oyt5CMFOvn9acALNtat0eD8MT/pM0X2dTwsiDbT3Q
SPuoy0/YQ6lx+gRGcKRYrqG/ezX8m9T30WO9cv2zsW17gS34oD8aZwhZmiPhKdWtdTRBWkJmIotF
vxWyX+oKRhzAloTip1AmWduaUzrxCq/k2bl0roWKkXSmAEZiOoRnLl0EODEVav4Mz4kDiVS1IUmF
fb2NgBHRU/hHq9p/v59Wf7T79l0pmMI058Zl9/DZjEOytLcKpIzrjcM5l8RlRzKNIAfEdqPQ3A6S
TC/5k8JpS1fohYVD0f026P3H5vrKd7dh453Z7zwNnynt7aYaDF6SXxgWt/5jXLUskXQW+u3rhZog
+VkeL3fgOh0bpouQfjiRqhVMxf29xBrO6kOe/2k4KlR2wpNWr0Yy6U/OwBd0LyFzchKYSCA8dLFq
aBZcKU/jDNPVwN/Ge7mzKhqtTmRxQPX/MU7+LMVYWa6iUyKIYr7YcqVDHWiWLc0FbD3OQago3gdP
76GkNsAWp831sFlDBN+GHQquCOWgX4ySQ3dnGz20M9ulJMF0ItxQpicba+OPv8VRDHVvKkxZ7nSU
0uckjrYXUvSzxy5/72zpbJCVELr84BvAak2QDRxZ0CnJGvXnLjDViW7crl+eFL+78NQ6L9/I27iC
u0KHLCVUoAsE98rSeLuRhhOhJP1IkCdTfVHVKBoTuQiuMDKqzuYdVjvUUcs4A76EMq+MKorLC1Lx
8NyQGfAntpKsbdRvWYB42pi5d7yH+Bg8CNVCOV9n5gkNm1zMO19REKISmzXI62ZhFDn+/u73t+/o
L34mEpwdt+z8xwqYBD8D7GGM/MBAsuUPtg8cVnENZ/QGIl2J+pFgfsVeAEZ9o7iYkcv4RWRTMxEu
Ra4JLDr0YN19SnQ8/u5wCOqqgRmi+6ZluhNOHvtb999cHk7/UvLiC81ptrGhqn/6OsPdk0YxQX/8
rKpM2Bqptn8xnEIRR00RUtLC8UfWfayJr1kTK8zTxDKOgu6GGeidoWrWJtpuYxrOjgj++pX1/Qqk
z1EBB3UB2BQwecz1k2elSHOYextVuGnR9zLsqVgPo3CuID/NtApXebndusUwED/B98Kf7jj1he39
W1joQuVEjJvKcKpz0AhWYzvgKluWkHluU45KnF87RN3BrvU7eAQWbTOXx3TFbDM+ka1qa5cvUIa8
fJyTTyqCBHyhufgkrlMks7Nu+Fp3qcNOv3KlzTm//N4AAqievdNRvA8J2sSpI4JgFIRGVvVn74NM
WcDEZoIPq2wMYbKL53lFLI0Z5q/TnZ4807yOnSnlHJgoNN91Z/GNOXiZVD0AQeuTzihYFdafTlSY
sfy13b6S2zDugTEqgBmmtK8Ie6PqMQD5emnVz8YaTuEggwgrroPohonRrRhKwoH/fv0+En8a6WD5
HUytTAxJBrPk9KWpdKOkjvRMfgfIVwW1rBeWxSs4/mRq8WQWBu2p+VM//9ZRckflztxPr2VMjZo+
upx9VZn6BGobhwwuj1gDaLhjruVIYmZys2fUYJXlQVytJGk3w9kUkpwEWojMxWQMWYl/3vOY+YkN
PgyrCiwshHsThSLcKPpEPzUKEDhb3yL203oWCX41eTf3vOcJ/Sv/Am9BGcQPX9qGCIVXUzVDpVXY
eEUh81fIOhUbVbiTi1TvX+AY8s1sB2alEAhMspfJ2w4SJdRI372ulAcYyfIkUVQWZOAFgzIncWGd
zbaNUb48snwT5WgL+FLBGuVfWuuZYgpcs/u9zKhXb8wL9I9GPBgQQvQWVrv1SgMYqCARDcHun28g
3OSb8vvDk5JDmD7tSU7lQMOa8Bydqsj9UqGpm49rG6P/T+Yo5IPCZrnWYkFkPpuY26GNUjZprMCy
MnJhc1uyIiah8Ps6hDUIZ30DCPVd7OqQ5LC/PszO98GrX4idydW5R9B2992muurlkLpnYq29VBJX
OhJ1Fy5tuMn1W7LWrZM5tNp/4DQQbrT6vZGDqT2sznpng8sCxXg/uPIcU09SnSj1ksDR3wnOn756
kaQ5NuBzeI66DLInN8DaNlRcBEIJbavc6MKl9L3XLQGyvdUvVcqHL9ZEHEwLGHwTL56U8i5acvxz
jVtKeb9rD3zxqgDWxM5dWkTlcFkZ6wKTWkg4zW30ryx5tgI+JrpYTPbcDcIgQwAppTYhxG/PSMus
TkQtQhkZ3/rzhN4eqHiZmddjk75+n5Siq4VW3MX/sUwCuodY24vQNaV3eqilRbx8mK2NVpMJYSiJ
JXXPZ2Q3CUoPRkeaQ9kKil1og9IR+QqWRpgxWkxwWPKBQ7pknA68yamTd8WSzjdm8Njjby2l/yzM
W779UMzp+9BsfbAGuOuBCfMdeArFphAADKsta7Lz3PQYtukxjIt0lZZh43+CU77sbI/G/O/dSuzx
D2HDPlXKjlHDRbi79Wr2PZfBZNmPcT80adSFLo+0l6fiSIIsR9FdeImudQ8pNAljY/+prO6WR2Tb
S3+wtgvdqxpghfi+Qz0DTZ2ocoOyWFbC7cerBeNmblB15d8CNE59xVhC69Cvnenf2+guBEAeRKcL
W8KoEoyEHJHMRPtXap2pan7sOUqEJUPUc6vH/gUA3M3EVJwKfeYvLP2Hs7FRtkrmdF5KFRcUK7Ku
GjhuUZV8P3EsCZrwQtfMPcmNWlIvFeHxYESy2aW8aBHNgTveTJ5R6T1EmOAfJqhLHnCMmRPBebwQ
OnFejCo+EMm9VOLFdlNstmdeVoHv69c9XHBjtrSnM9OJo7EVWH2KoVmfPbkbBkIPGL2pl25EYAUd
fw578BBaKOvSXGKOAccCU4kP+O/p49zloBoRegNhvz3co5lC2Q7sz0SGt3LLeDdJzMCb5SYQhBnE
nIEloeTLUmOusl0/Z8vTS1cN535EdLwxWUSZBNqbdSqPdKTdMtgrxguHnBFd6uJx+EV7JiBs/Ogm
U3F6Lg0eHru/wPY6WMWHiCMAkML+jyBmolUTlUA0WtNiukWRhskmEU4mtHfp6XgyoJzQCUBI7DZw
GsJHfxpTKFowUaD9q52H+0RGAJX/7iNeceiY6n3lcdi5VGmEmtWCvqLu5a8QfjNVaqgBz4kyuVbx
RfZNr31CLwp7pl1jShdoHAehO70xVLySdNR3Q/UzxQVShjGQtXaAGvSrksfHnv22PmFN3wi5+n9H
34kVNqOCX3fGbKqFZZdxLFMdBuIVwtIn9LzknTesJz3oFfcwaP7UZd/tneH7fg9XAJyj3NnLAYLN
a0QOTR2enPMdceDqDZeJ994B4Y9jEniU/NLTIAn8Q1Kk5xo5WDJ3gI3oWgRw3yHDEjO0MWUPCbMk
7JTNohgyXmYqn06guwXo7k/NnG1tHg55MBMMIqpHscmYyhWG98XFs8lWkRLnHEi58sX2S1II2WYJ
dd30ys/rf9aeOZihsCO1jU5TQONABW7WvNI5HRs01xOESfcHA4KA25Y6AisNgDS+fH25Syt3XbL/
SfFREq85mDGgheQyybq1j3axoRUDiJArVtT/M62MMewFG2PN35MmEsG4fdae2YV1A/e48GLnyHSR
wUraywrzvHP4XP4/CauDcuY76j3WC+OH6mzG5+tI9NxKnzO4M8boE+UnNJn0QEFR0ijXc67l3lHQ
q7d/dc6jsjxe3I1NjFxTmrBEjPLUuxBs9srPoU4xVvi1IjHbJA2SEiWUmW7vr15vflAHLEW6WbF7
23BbEW300xFpcoHAZVxpUhLErcmwtIvQY8pGV5cR6rpwHIUUgDMfsPkx48B8b9hRej+A2y6VPakF
uPApa/fca0RgVMOLEaCC7ZRB8dX+9Lx1Z90MBGh6MPwi/b8rFEy1gAeysH4c97VNRmUssFHD3HHk
hzlaQ/2J+PLVejYCgYs42KT/4/rhxLfvy/5VFoYEr5ngGyu1lq2XVKHQhhuS3aZ0KZShHHo+HvQ2
qfkIMe2sJqQ0rJ6a0+sBaJOYR3CRoNUmAtcV6KEakgQxDVd4pOfO9MU8Ty9g3igKaXBHs0p6E0o+
Q5BgkaMcnJNo01X5K3nnX7LKfmjNNsgERG7XH0+zNsmNbdHQwmCZEVwVrCLjmm63xfz256tkmP5v
kqE2ZhLswR5L6CKMnQc9xLsvztDsOp0qkdwRpsjXD54aJSaC39Jz4hQX48D+DW+zoUqIheTif0eR
Jm5ehX/EiuQ0wtKWJxL6VGNBg4urOVWxMSH2rArkvTm4PEipEVmRz3nQ7KLoeVbHJ5YXadQyYs64
HPuUHxTMiWxoDvj9VS+wP+1T4sMnS9pWB/Gw1nq0ZdDQrgNrLKV7S9D+poOQ5P7JfmX6XOT9s7YT
odUE+/CsGXqx/T1NajhyRa6KnfWax73HESgNK8Lo+uIN7JHR4BoO+Sn2z5iE3aVnPXOAQi8dgE+i
HlsMAvuK8LT+afHlv4V2ffG53C3B7PMqDfJN44cNyGFlXz+M2xOt8fAwLdImbqjZbKo4PWfWvC8L
YlA6zH+FqRMTvwSlP1+GLLWGhJxmg2XtSjUzsaQJ2awzNFQ8IUGLLHO5P8SEVF4Nq+wcH8QJYjdj
ZiT6P+htqnwifRoVGBHS64vL0gSW6unYOtbUzdYwNoD3+ae/hip2OjDOf/DFH+YsPQcBOrmNe2JZ
ramkjDMljXyC9pG9/sg1p+Y3JVvBKMvMyKPBnw8wi0JevaY8SxqCnfLHyWAI6oxGgwlTTO9BHnuU
hr2S9KX2uU1NslD7lyg8tHo/Sd0XXxfUbB7Wlh88Ck1MUCEFBJdG5V5cRFog4ABq46XYiIBrIO8W
pU6+ZnE61IOz56CcPqeS6Qrtu82W7IVkd5oeazb1uI0f2swAn39bjxTn6qcDdXUvH7rAyb8DXrzE
goMLfzwB9vEhQz3pr/bMRxnZFmuSp/R5nh7jjHceQmex6da2g0tfJaCj50tuU7ZQHfYZ+coGHYnU
QggBA54O6/pWSmATxOQ3+iQkTQf99o4aQg+y48Q8FmF/+FAM9O98OpOOVIdSMv+Ag90Gqg+UtLud
xjCloM67sGNBWj563Bx+qcq2koKzdF0VqI7+k4Upmyf2V/of608IY8yhsG3fA1zTtNenJgrvISTx
2Ig0Ty88lEj7MJm/lc2DERY0oO9ruO2UvZqCzHXFfmY3ka4+YJZOvyVmLJGL8o8Q5pnIYcVstvIe
BOq/0oaelKJapr1V6xeDracZW3VvoQeSG9i0bcxfnVD9ppE1lBWCPoqu1oL1ISOcmzNxkiKahOyZ
06UIH87H0fjP3K9xoED+j9/O+EcW6foQsQDFOJARkpZYnKCuFfJOFliANbzUSQy6VBU+3B5kkw5F
eB7c6nEzmJhWIEVb4RWzJBZKZYMjH7ykQEZjW72jIIj14RCuqyGi8JauTDvC6L3Genmn7cJMo1Vl
0qN7mFO4hGU3nPs+ODMTaZ7eYpFvj5JC73suY9HOEnS5Tlf++hRhZzDCGQj7i4AIHM5afhUZhqpm
XlBVnEAvvo4XFIv9z6AsXerpvF/u+BnvkNVigBSbYTuMj/wWT8VfgtNvkBD5QSlmCjoWDtygGmjU
Bh79oJszXkwuSqgbIaYOePm93NmVzXvEJ3TKO5ynbt3ntYo0jeCKFTGy3RqlWKGCxcv1RZvbQ9SL
LdwXfPUyk3mZzaeujbHdjOmwbo0nYWzcqXadwmYMkAf8fwzMNZXzlHVO0c/QVUfDyYwIfDOTRPjY
L+T8Mpv2nTmLWbC6K0VueKSiLAtBsFoWZk4rcGmTzVxVA203AEok/RXFw1vHTBWEvpVyQ0thGqm9
/1s1gier0Qp3xUHq1zSSvZ8H54H29mDazGbuj/GuqAyRA5ae4D/4s/vXkOrPFtu0sImU3ARCPax6
Pj8eP21bRRbp3hPtYPELpPqOWIdyIHHOIrJ7fflgKb8QlYYovul8jX+FV0NvrhGI0tCJkupboQIv
CCRxoC0GK6JSDCLAfnz+cc5Sq7WeHZcIpt0yP14H/G5EbU8oJenD7mqf2NQ547a7SYUiLU5XZBL5
NZTWx1siIlLlqvaJdy8l+LPRfcxgVeSyeuX4ehQEvflpxXHzccJbAiFc1So6fsTH2nXLrS6i7Zmm
mN2fBJznVHChTLVg5zaQqU3LT8/ke8fFdj87QNKRJNKvH5GM29pSq9uRC/MBwQdIgh5C82ppuVLj
T4ILOTohJtXpSdqbiv15rXE8/VguzxRKtcrDBBP1pjJXOx5uaTz+af1zOmBhRpbnrF33jRQ/r1vp
HP/VuJQsWVj78qW3AJe3AOsIjmv4hoJDgJ6sFmfX1nNJrtbL35veM2SxSv4dcA0XG12WtDvewIZa
qeJONtUNthHsqZ0F0cX+ig5ag5agXTduDn833HOX+VnX2I0X2NhCQzg/FwPeAj3E4NP5jV4XlTmW
MtA3EKIfWRioGj+IHlDyW+x+C+hrUKvgp3gHlkQn5dECstG0GxuOvIslWdTOaVAS2v/5jYLCNDQa
jXUEn5x0moLn/9OtStNc+/re5rHoEBv6qyqszw8XAUVYWEeSZ8qBYHRQ6U1C2gALvA4mzCj7UqAu
98xnov3W95yD5zRineQiyKe3MFBmBDjzj8yBmiqROB2MAriYJftNAjUAF0ucBcBF0dfe7gJ9X7EK
/R/BVQmaHjNgAL572HT8ALKFn7T6YTSxBDrZ/pZyAMnvXVC/x17MK6/883gBo1TXe9IsDNVNh81t
wrsLDxZ/IzAn5mFNlhMKKMSPOPqooj6wVhjAyZicWzB2mbvCvaWqqWKfl+m7wA2yukCpIR1yPW5M
Lyuig3De/8kZcpuxvUVBqj+QVUS4Yc/zRdrQRmmiGE6NPeM5nNSKbv3ta8GErrn9cQQWqTJ6Vgwn
GdCioceTlyMGpaxRIwL9qqRXpOKg8Ji8BTAv3CTxr8hhb7SN6afVOqAWIT0U03S0vEhQtp5rj9vo
fOTjbcU0qx1GDU/QmcXaoeVrMozSWkPbQlA7uG56Hm0ji7ZL065SohH/Pcbb3p+puZ2l0GfkGjz/
zLnwmEGjcqQRzXP28wNipUK0ZQONTpRrn9NRhiFHzQ54/4YFaNO9QxaLCuI+fFH0laSWUJZefNW3
9EF7nc7PxPDyUczppruZX8q4gLssMDWH2nHheemj35oKpL4U3UQgHmzgcPZUG3KYOE/nIJdf+R+H
horCrBEZuL3DiXA1buRWdYF/oC1hcjebrUW7Yy4fFucy9Couxul1q3CliPsgpIYJyeTPLrxBR5xW
m1w6JkFZQ1L5qdQKHIEOuHIFdaf2nlwDSEeJaNHyKJMWTsOXonQrza/WLyz8i6VVjmKB2QMy7yeE
Ypon9KNDYv1As+PNRNxXIgyOgCD+mG+SmUuZMGKeaI46K7VKADXGxwzRZvbGLkDAxdcBhoTI1KX1
nyMhS0g/pLljPPEcNZZDigETl4Wx0k5EfYMDtH9amtBHNK3NC+M2eMPT6gjON91ONihqOtRZ03H8
mFo2S4Ujm7eSb3ckw4CjEosweFDt3/L35TilrO3sOtdZX4DnI1gv5kwlLYgNzgxnrOjcJMSZFnud
8yaJW2EQ9WDh8XBEqquZ69PmxuN3GlUc0cJv3jJQ/cEZ8c9S2jgvGEQ4RmsX23rzLKSDtT5KKX3E
DKS9BwV1CnrhA8O9/gcfwvovKo6sKagNm5eQDNDqiQLN7M1nlrPdoqFCddtxiiygcorJCw320DoA
hR10kLVqPD8UCX2BBpJyxPV/922dc23y4SF8nQr9RWAG7m1SnmQDpAsrWn7GtITq7XiWmafx/boS
BckBGelBV2fD++vbWisAgp7ZNNOS/nJxgjmXOdQHnWGo5B6isNOVSGel986O6sAbHzCTeLZ8QqHl
SvGhKcHJMjM+gbCmh1coEfxORqrAU2A3AFMn/+EPxYEE5t8exOftvoSUCaqRwOEskrhhxBe72Acu
8pb1atw7Y+06QE/tLBLQniGqnFOoN2tFQ22qj4ll6pZQZC1A6xwev5ycBshcZ5ehnWzAl/GdJvKf
TS+UbL0zVLf9eOh0LGgTHPUFPa6VHw6qK+UlDHA7GTvqmEyYxZDK1wNyNBh2zlCuUOSmeLfjwvNM
UM4vUYS/pA7jjFRRz3gUH9joQkiUsAKI8t/ibqeMjcCLpUL8jIuzz16gCoq3FUL/k087DuGPwbWP
oABJKxgdJZScO+IjHNTxjQCL3n92sBu+0rgPj1BM6+FERUKFfWvSBZwxQSDfFQUP4QPoUujgIbP1
x9c8WBCk7LGS9Kkv+nKIndY3LeZLfaOiv4I8OnmsHYSDlPK4Covt8zEBEDUrA+Jt5uMxdX0lgJh8
dcj82abVqniCgyXm3DD9ropCBbPvgVhbYiluj1GMvZaq76xrLvf3T2PAniO+q2Q0Tps/gW6JwMTw
Bd/PNVZXR5jqJYowMMF2M+9AeCvSBHEb7sYDlx3Lq4ucUWygtvIzQm2GiUibvGiK2xCiuFXKtsqN
VHpbscyAeXRep6Cw0VeAm6ZvuaUisFIAGu8+GZsFkg0/JA+naWMAvG+sDB4Rbh4yQIdgFgZtxkuU
58ZdptChK7GUi2AGLD6mG2jTcQcRddkL1v72nZn34BTpepIm4du/hdzRFJz6BiVLAyKn66X/DfMZ
lwEa6X96Qac5+MTQYeHZUdQDPCjg1yF+EapcNXSRUFRq4hJBrK87zgs6viEuNI+5p9C/kvUUZkGZ
Lhqe+Hsw9f2YGe7vHPuTSTv4kuQwVK4P4IaOUM223sbgZJ/GxbjukeIaY48oxwKlErxlpmytfear
GN05ImhDu09/kt6wfmEpeVk1wHfNzZczGHlEvGo4/N4YkTa7GVWonsJtA86XhfsLjdtkX0Af+kj/
wVlbzTJDGvBfZoihzCcBU0PvsbpkNPMV+5PCanarL2z17Eq6KVw1+qSV3r24rgj/61Br+ReczHGQ
jF0oRlHuN1vbRyOZc2v5cphbxfTY4TAIjvl3lnMn/JNteD94ZBnpTqRaKFySAikUfp5kcaWvq7Ke
hA7oxAb/QtaVxxhRG15PKf61DWHxh1cE98RPJinyvbWnv2iln/pJyE5e06BN5Mbd61GHDTjLCVkx
E8b1yIoBbby9BgyPhkoZg5FFUXuqB4ip7sYorJ6DXXi1zs7mk3s3rSwZ0PLHntyPm8iCPLc8AoNY
GqK2fGpt5Qmhrmzsb5hAO24p//GfO+vAZqvKINM76CWGwq3bULSFJDMktF4fc0XC7GWrAfzqXMQN
TbmeDgX/rGLkpMKnevlz2+0Yv7HpPZiZE4A9Vol9iKCvjBWElMhVmtR3xbJzZfL43EnFxFnRCuBI
aiI/vuRBHQaP24OK3FuniIu/aFd2ELLLTblLoh/+Gj8DQ1qe1NOjs3eqkB3h4HRq2056Kk4geSmI
X5E1huRI5Bc8opZ2bHpePPdgt5fpusOMi/d4L+5qT1ZwBTSua0/lB4vDlCIwQCWUqWT0tEkn3glv
yJW9rDrRvDMqHDRRulx96Xqk01C/rVGRM01PupdJdQSiSMB+IzUhESFaf7SpewuOxZoDfHDZ6Wx0
AUL3RqzmQ4ZRSdAF08gQ5SgNRbRStm3SMgwEdk9eMOljDRwTO6Robf/j1P7nsj8xFUUZ1hpgJ8V2
i3GoCOc+WDaMEJ/3clnLEpa3uvuYbjt8CBMGqrKdFQGPyPXYgGt7h28blR2cNcAuA40bPWPKYFFB
46+H88KtC8S8F0BasxHeuBwEe6q8/uuxNtbpBd77KDdL4cnE2H4thX6ejbjuKm/KfQdnEu7GEbdM
80GaWGyRM12aDNw6QOS0AETPyU4SUo6MWNTLl9yAOeB2llm/jnMR7MomplZw2ut63tABqrH0gbK8
pQMeZAeKmRqNsIwE3cCd+lWJoHmg6pFW2akw/aFbGP3giGglrQRhOGJdMtbE9szIEUbVPE0sQv2p
U1LhRvYMSGzZ+mpXEwsDYFO0KHfiWYyofrbo5tTH82reGva7Y87zewbBFs3KgTMq0vHbLESmJ8CM
G+WA55m3mWxr4Z2Yrmlz2NVQDdrRF2DmfVYBiPlgwE8GHgaHHok7+u2eiyNGtxYFRxR/XSn9Xrwe
t3lh4qMUTSr/bMzX2xAuKsalpYrR8vsmEKT8jvj6uFtfI8RFXQ0p5Zhly7Gph5KgxRhNg+YhabAL
X/gNv0YLmiI04uv93NheSvdKdZeDYSj+c/wJB17v/ItvxOGJ9uOac5WTf8UEcBM0zgXWEaV36la1
tXdufDUSkB6htwMIYA9Gth4oHjlRJXkbGe91eDV7ourr0g9bObzsv/eOKqQYhsNcmylt9j6j48Hd
jPritiS310LpaWSeHEVu73bGfOQVC6ngqSmxsnr0QxGNoLFcV35c2yDjZLtSPsil5tXsf0wzv2Ce
X8Gl/QcYz116UUJmKsgVVQ2EB09x/PssW1sWlsJyQD6tu8hqlowu8DjuLz+ln/uWco6+CsD2S9AA
cGeVNe3QpZRHPwieydBTJvxt5c958N9YVZHe1Bqem2wPTn0IjQw6Trbbqr4yTxMPw99FYoqcZEPw
36sqYYMPRE+XoDA6xHrDOip6mgDnKnQ0Hlf+EYGhCYJhFaTfBR3M4Tg6AWfdt5ZYb3NE48nore4Q
iECi143xSYycgxBWlJrCVpaml0cW5eNiCxnZobVNSOtTPdPbOHi4S2raNg1u6Gn7YBeHLhz1Miwq
6BoHyf4qxnAZXWISAxHL2wBHeCRe4rixyLQsYSFCdjfZzSN/SjlWFrp5Rue3AnZGo4tPXuacVKiJ
mNR/Uf0le/uoHL/FAnpH/YuRTi68J9dLVJ6f5wP1hhS3UC/jM57neUbOaLupjqBqHzfjf7BY3vQ4
YC95U425lrmd/DFIZKC9jVxZYVvtLSI7yGbNjTZOBIzgFMSaGixOygpLslxpiZ4ItZmOS95J/NKM
cbiftqmC/lG/Ey9nYfCcLUQeL6CQZiv0IAZeiIQcnqzXHIQWalJsTO38swmunaBp2XxQ2m5TPw50
Npth+lwFdcFi+c8m9A6LQdGq+pB3E7ccpyUFU2W0C/LqUFt+HGwBYP2cEF6Xk5SnItvTMBabC6fm
wRbLzTeURaclxZ6Q1H7MJwdQUEQeZshjT8nHeJDTc3Qi+4smq0A6rInxmDHI0bV9wwaXVcaNS/CE
dSqq4KhJDUm5AL3ouvsdIgzX/KH4QT1vtvmHQXM5e5Yt9FUqrmh9XK+hnhqeDL/P1EBUuvVuy/Ja
GumyBOgNQJ/wgRHOgHduqdGAwyup6Nf/7TJBHRhu6spCNVwKdlmbVNuuOIdsaeH5tt2vs/h/evE5
Pc0h0DBKBr5+AudgwJ+06Z45O9aQhXJWub7IHn8hcB+dFQOkQU/aflTWYa9wne52X0DMrY1lgLdK
hLer7i0QifcfNv0FjsQsi/e2FJsgwQ3Ab7OIRiSvayejVLpzCAoHUEqyblEH2WDnvjXmMSh9+/NX
acl6U1qzR+7cEjhs4LHpjl4re7yKC7zsVlge0mt7X7j5L3xXM56OeALZU0Rjn+pyYYV8XitMbjhi
bdl/uUENdMJcpd2odkRTBvyqRG663c3NyT10wwGMy85RLNk7Ro2aN8lD0uvLAM2wu6mewoZtZsGm
NvxKgvGLpYPFEAtN6rx9n9YuyAEbg+6QwZQcs80ITOA0k7Lk3wfNUc4JtEthQXQ70OWjzd0YHPqc
NLROsBtwHxcfbcHvG12dCeT8K9ZXS7QMDHkRmyRc48VatJPGQDMmKGY6ydKtgkQpXq4l2U1t0WSl
7B8QeePpDT0d8uoESAfD5UZhm3Ah1mgCsCH2wy14nY44yc2ckt8udV3pal98z1WgCGJXYHGV+T6R
lyICOSiE0R7TcU5URqiSjktber9oPODjwm5VGpSqqkoB1jmQjRlsMQYFKPmCs6vrKxUv3rYaUK+o
3pA9exCIsX0lLHFuN2gcz1EQGv+fA0kW1lKzdv9WcJwiCZ6aSjmFHmzfE6BVqSj0b2TkZ5WTlbUq
hTksz2mK9BL2zN46dNWO1/8J4LE5lHP5/6/lypBrDbV/a8ZTCugxadV4nGztn4N+VSJy/sWQFL5i
I4zmMwqhobWIx/LL8qeX4NazMrH0DC5dMOyU/xNjE1b/aJCTOTHoZyKFdVHUfn2hLz3JcYK2Pk88
vOYUkTMoW4bb4ydR/xbnZm7gS796X9C4KeKhpCADU1Zz7tJsjFaMHIfLaJ/9KKeTSbuN4zmdGB7e
ki1Rn1wNsdSIYkaNT/5+0U91udFs0/pUFSA5Kd4Fj5/JAv6rx8qd+oj3P3RcDcT7X/rEWPKSTYkD
o/eiMPd482vAgCBaKVlQi6XoovLxAVD+rHp4SoQ4HbJLzRcNRgxTUTYuOm8lumpBhE/DzyV/yx60
1DeVVRrZZjMp14D52iIGAKtNGNYxcOl8WgnNFIVnR0TAKhWNU0dU/I9GdB1qxI77dl14zIDccLvf
UYJxQDdyAVFzv4rpkRzeofelzfSzzrsM2Euyuwqyl9LBwFDTgawDKMbI4YLEcIyCxQz6OK2w7BgL
c6iOyJFFQxolLn4oOuTPAhHR505akK3UvRWHWuqkb771ZBd4odZ0Yw3jNvqX3KDp/OSJImLOczAi
UxeyNCWkpSjhK+/YR/Uk3WG9e2jsKDdmtrmd9zNefhN1lgW5NtzZaYwPDKeWPVDjTPcOEwmomANB
7INzt4FOTtzH1UNl1gV+p1XLAhp8fWYOvZXYpvJrwgVjThBhjHP6qSDcPLLtZArCBdN4/3ji5Ke6
hpFWg99SUteYlMF6J5VBlV87TfNr9OaGTeNXSpgHaXU7dEc4qTzvg/wM6Th3sboG9i4CarPldtKl
8yGeosPWRPPhSXjlKxQZ+1s8jf3U5q7Ab8tT/fbwoiQQUnLz1fIFURYk9sHl6hhe19AK7pldG4op
vehGhhrwRo/14SY07tw6l+ybApoGQdL38l0UKOleFQIrvJZ/GdD2v2MiVhmbLEJ59S5El9+RpB0t
ei7BUp9UPFWe8rP7UccSYHvXPc3op2eNdrk3IZ2mSGN/xgywQh5ywZj69qmdexHElN0AIVKOakpD
domBMwLFQySYG+cpHZe8TLhAQ8jxFYad8HaY4kSu448hhUBqlBouCjrDibFDRDNaBmvL4fWhEq9v
L9Ic3cbd1+7YLZiCtvi46KF5PsLCP8JM1v/XxKw6nV1jcdlNoIu5ldTUaJwGpBdoskLjYsh8dJCO
PgGXR8W3TnzbjHlwCqcpi5ozr/zjQOVxHekawc4gy2SjUv/+PDdF2d9Riw+SSa8BKRp6kTQzOVOi
U76yHGSwixrNTORe9wZZxxg9iJHjtdp6a//m7ml871otJcqmgf022Qvhb+fH2Cum+MC4pThmKpY2
lV/pq/TpV00ZYxgmmDa4VJ7BLhWaHEHShaxc5DEZeB8cgKVzqJvIlruKRZ7bFYlFbxlxn3W41zHH
Cr+MGVg7du/+cCbojXdpbrJqeCP6x8AyYyGjEySHa3FkkX6MJ/ywpOPvaoERqprxi61qZTyUVw8c
4zd2wuw2oKONS2x2JnLQthJpJtZp9NRXgTviuOedS+q/wvcACzPVAmErPLlHhMDGLCxhzzlwltxY
eyhbVx2sjQnTrn6RYc9kAz1xkiFO++eOwcvktdVHTCw7fD5kLiAVA2fly0/YLr4wbJbmXccN4iGU
jE+0kPKNx9ku8xxOtW4QL5bQwC5Ch1ZNaGARFXqkyyACu6cYvL1s2aoPq21cUz76bMAFVDxY/C2/
G+npLh0oQdCrBId7ynl2m8iTcftmt5gmXKQilrZKRDXtpLv6VbhalDK0h8kGdr+a2JEnWdQ6r7sQ
fuKJLvCRcYushrV4diJ6LnDmYbmuxWdY2WS8MFQ+CtHEZSGVjKpTpGMWc/rB7gKTs2Z8KXngy1Ab
CHddx78Gk0xMloKK84cuk9Le8HOMGItQjuqY+yF83JYqTaEb6iX6QavjmOmRoYKZ9Z0eCNybzP7H
l4QFXcaToXmCONI4IlBs39jRGSwUavjpXsw0Q5CnTA3CjnDfGimejYFonZLJ+0A1p8J6N8uwUBWr
3Yhka9K00T3i/y9D6NFIEZwEpepl5GlcDs2/l3SzQVep7AKIW8Z9AEvWlIMLXaHpN7ermaHXFQK/
+pSMi/1m+tLQr3b76k+kGj7NSg1kHpLj+wT+lfeXTKiLDyukTCPomdJIOiu/ALLPolA+xbwlbwav
3lDqjCIRKpMC/7PsjoLrsR7UDGkoPImlDMS9hcyq64na3Iu6IVt4mjFQY1jdtVWIc7Cd4tGCZUQI
uNcZeHplcW6LuWyxcVzt2rASddPrtj5K+zjOCH7lwPFbm4Z9/RLnywQjP5oh9mFjcIDhnObMc3xs
xqMX4Nc1K+SkiZISuJvTmGwvLwnjiLQUnlFpThz+OA1BpEVT8xNBLAnxd6+QY1yOzCOZQsYyIyaW
TEWYYbdNTt82+uF3DKrLtgHT5+UKXkynvoJzsKbkKOJjK9UlOU2ORV7wgATk/QnzrS96UrHiJexR
gH/WXluhKkf7O05+u2Dg2N0aMj2afiMI6It3JA8C67ENC7FYDjpwxwwg1ZVBAYaUENf79dgPIKiO
tKbhw5u0rFYJYgO1JDpaAaik8rgL9z9DUsyZHjp/jC3Rqh0mBA6Y/HZqwYkBnVkgMjmVIbwPOTjv
rR4QYfvP20Ohye1lmhGMcdsKhtDtw9PN5Z2OgWvS2ZHUrUBlp1WFsLudrRQi/CN7G9KYr6Q1wZqf
RVp99ZPtCWtFIVDpjqgfzcRTuHyNFYHQlAJ1V+8PQw3IBw/UpG3oLoLgQ78hjWgwoIlmnKmpMmd/
A9ZUKolL3GMwAMFr+pF8ZfYrBqg6KnI5Ho/HchKhM0gMNq2znQ/ro40QuWbkonUfgqvghgjZPhTc
kSmwIX0Nhr7REl+dkXt6xPXv7bunFbFmff8MQbp2m0te5tkhSLvB59JLobKeQwXCA+gJP+3yJ0Pc
d/VsMpU8k8v1FLU3clTNip7yKS3rRJZ6+pRngiHR0sXV4ufUe5nTaNxML13HwBWhh+fjknLnMbZP
Fc6nirz/DmsrmF731OZRxj2IixrebHm8cBE9rIO4jRU/RkNpX7DSguOO9PjoFWoJc1jOM6Uershn
wvBIgud8/5GMfBeH6DcXcuae8MvsGLcDIHnXYTxmuONvLddyRH178AFW5LlTUsZW9R3aUZhBmlPQ
Yz8eECDeqcXZtlj+c5eQeelMiSQUlN/F8/lxdq20cR5ZTR0lSyQTxxjjDkxZP4oyLksrNe0v4HgG
U0VcXrwrGYhe2+iJ6rGtrclGuxg6WdP3Qs4FJ1gjvOmnmGV2SN/9mngzhtRTJiD+WFhOVHyppOnQ
z4uOgC4ZsRg5/jahco6cTjQugaHBhIYm978qQXLs9k3lT6gP7LXTSKN5YF1pg3Y+df3cWvCCx4Ll
67ohyg4ftgtWeJPnZXe06WHDno1OxjrrcdeDRZkeVDdBwyo68iPOaLsh2lYD5nRxI7ORj88wpp5X
ZKVzfvWEg0FboO55pOh+zLlEirJNmcrR6SwbkDqvyzss/XodKNBZDrIY2c7Pb7/Ch0J3lfhaKMar
oMmhNWZYBRXll/jMQitszPOvVWktXLVwj0sfns7CZfeX69IE77DnI2szmOAhhPBTlw6OlJ8c97m9
LfBydxdTU1n3xrdPyHmCX7ldv8Mr58lTEuow89LBpZyRW0bMg2+OeDWwDKvWtPIJvIw6hrehk9LB
AXn+0n5PiWxIGVS6DS5q9rSZc69XBhB+0dtXy5rXCGST7JQKnlYMYgJR6E5KY8amItg8HboZ13AE
Enbk7zbTlkk+cWbjEOxKUHzOwjKY8Z1EYFRrK+UqUNzJ3TdbhVB4jBQQ5lL7vyY9zXBhUdKorym8
g1AaHvOGfR+Kj/SjITJre8+q34hLLRGLPXrrJO5Cs1UG2PbagcOprFXUShiwbr2MfnF5MFGh/x+O
dqEz5FVajtc39siuJrjDmWCuuoNVppbZw3VeS0LkpG2j/N+R+EQ7XHgc9LWhNAIk01EeMri21mcc
dGZic2Kl/ruhjTODP37IkfTRBTLkJ/iYa2JA94GxQc3IJ8V40J87ybLtpNfcW945MGdtZ8PHhDZW
427BMPgmKs91saJwJ0/ZoOJQzbUMQ4FKgy3bFdG/6+juLomoZeCKT8V11zYpcufaLvWMlylHOhvY
GHHflTb0oLvcT+M1lFu3XAvC94IEttDg82WrkzlIVnxkTzpMQP7xcomJ9MZ+wyWbwO6+rcoG3rmA
cKfz9HThJ91FTPzWDJs/DHbkPnJXG7keWgXGxJrY6papg3sUhBDwanx5nWKTEo13SIzRGaa4P5Ge
MSktdIpDBkS/Ng3RdLolYWu4RK84sEGZQJM2NgdoQhOSIlyDolcOI82koh+KLr/E0pggj1+j5zSQ
KaTrFqwRvT7JlYU/g4BPxKpUJhnFiaQjunZuErvHn6bx2rUOHngADluoS8+ja3lnzPRC221YMVKl
cN2mOM1ivFoZhiotekUjkRrWZ6sznokQglsnVmQ7I/s/inulG8DKWP2cZOvu2hsz+ixUNeVhAdhj
S2Xh6orplusRMRLnvbdyCr7m4e3loD8JFlK5fItMO6EQ3mElju63aWX2wxqT5Xd00RNPjUgcUiuE
W0pp4XKnxzZY8aH9d0+zEPs1Y0acsf6AEZjl7aYlU5w4VivhX1yHY9nlMZ0vN9WJIGJ2N1cCW1lu
XJ3PMq4wfUeeL9cOZ3VYTXPgmwqlA7Gz7WtIs6zy9k7nvXdWKDbXrzNDgCNPv3kHgrGTdNLWamQ5
445qHEndrE8Ae+hoFLeOibhlVvz9+pJKOBX+XwlME8YLKWYcYw2lTtSPZ+ogq2CxsJeT4neuwN6c
OpLBODSzOjYuKZ+scCQEu6v2WbvXPGdcOx6RFvLvZQUxo6/TSxTRuSG+ATb2e4TZZlcFo1HMCdtw
pN7WCW4eEk8dOh/rCX0bXhCQek/OusQNMYbEB5WPa0xcw0UD+M/hlsZ5FWbcl9wJrq3CLeAKEIdb
a0K4G+3sFGqlNh9LJn/canmW+35uMnZD+9On851lS5A7r3MJxYZ8pTJX4J30ui84tjk6adnyg1HS
MFUNkmPuvZ87zVUTTgTtmpUX4t3JsibGlmk0EQB+YPeL400VlXWnfNqQj+ePFhOQ75KwESD7O95g
Qg+hg3H/CmQ5AnxIi0TkKGcr26sjx4/nAlKkGKcHA4OVvfhdXeH6jnp3Db0PxjPK/s37Uwyty7iX
zuuNhskC0Faqt/rvCupZ9eKKlS8dYkKZ7f5A/G3IlfF68j7yZwciX1FvJNO2o3L0A2Nqeu9JyfuB
1YQHPwum+5uLrhmA3SAkuCMRI5ouTILQFGgX5F0mGi4XcqfQ824PuoXZ/jH6HNwmchisPrbgN91K
sfabqGwRBPq/T5CZHfIAA1RzSbTdmVcjqfKfEhaxeNJbpmrDT74grOnM6aLrdn1wxfAHj/7jnp8B
McWgNW4zi4BBq3j7mSGaY1V2V4BMj9vN6pTHlDjpNU+AQ1SZ6cDwM5WMM3nZ0XYhQsHezKYlmbJ1
a50TZGSgIDnLsmyou3DizgS4M/p9XUbaVU35yFqQ9RVY6FXR0+4TPP4H8/L3Xig/xtgZwIzZyADD
pooGjPfVnJYu3M1a8GrOYHnqe3xBcw1M+wK5E7O7btAfMcvt4Bua+ksmIM0PeKOIZe7FciyPO9CC
VvU7v0CPC7nJKfYEVHHl62V6IAsV9SO6/K+P0vpPD5FZNBjt8DluqSpEnVeBubaEQfy3mRs0mR4N
p8Ntw5yPgbcUoDuHNL4Og4bJjXKkE8H9srejKGG/dSJadr5uUqcTYmd2jY6w4cDJjDHnurr/saKd
BriKKxWpx7GgA4YF/aCVSUTRQdP3mSHCXSURXbVCkreoTZ/PafdVPZORNWLNpZba4LhxkpEhPBxB
w5yldU6k2BsW+kzDJuuAEfPjCuJmQ7+/tEISZPchbu2xOwq8hnUMyYGtElL6SLqEbKMKohauDZ6h
Q0wQtyoExhyKKut0Fu9SfkWUips6cSM/n2UQNI5oUdLkFLbOG6T7qTiFsVoWoLgEKZb79XKJbkw5
waVwwLG+CJG8VPx4Re+d4ZpIU0KzFdfqL/f7AuJwi/VUdOl6AX6tDfFgi5XusI5/gctFWJPUmQYn
TO7A1N0VKqF/H87VwoGGgL585gq1I3cCU54RxPvMbUm+xN60GvBbYUadgNmCyrXzH+tFdvC2wQzv
fZ8G0GZMYY4J7FbTaNWHayu6/ycx91fZ9q6yNtoEvLRMFkGHG9Y1yzyBJlOLG0vBVNeVaSkENeSs
g5cx+e7eCCyTVJgOZPJ40WfFL7M4t5Z7F3nPsa00gc8WRP0Gg0K3K+yCuyOvvnT/AEc7LIfTB2VN
Gns5etqvIB59gNHF3Ld0a5lIdCfnufgASXhCi36znHPSQpMQgZPSkXybZvLjS1opNH/dg9cbDs+V
KCAqAU21P59CsCcTSevjglSRN4UOnbcW7R3/VQE+MOAxGibKl4LDdd7X7cLecJcfaHQdZyI0uBb6
zZsh8DQh7KvC+LWAATvdpJvMnfoiuORmgDOZMM5t0qGoRss1SR/Yf81qMXNldAsp4L5AOAQCoEhN
UUuaZvlFrZX6lLq25Xx6pVjr1+aYLISSd7a+5AxliRrmygLvu3LP0bPQG4N/Uq4lLnRasII++K0T
H7L1kqV3Vz4cdm26yykyCEP8oOVKUS32SD8nMuky032QybxCm9GdyeuXH70tqMJ63sc0o/A4mHT4
qsMJuk6g7i2eA9ZhegZCkITDg8f6Xgj9L5kZbTQ0CTttvCMvTTVfH31U0xWk+Gj03SIJ9aGRS9va
nvlewwqeuF+eFxUiU3xLDhO2ddF8VfgGUqaUoKVB+5zEQ4Y/yPn/6DsleG9gSyJnJHa7qY8EZPfP
cKE68eXNkQ76YDhKibN3KfL0PiwC9U3ldoDF/r4wsGTvwVSlL9zS2kaEf08S5qWVWZpsrDtEbJBN
89kx8Ed3ZN8+lybsTMov4LhGbnay3ZwsOjqbfqYvocU70jQnesBpigC4kOW8z1qZErli1pEfcJH8
r2U7cL1N7tP4LDXSyjiB/NzfH9JQcQ3KrU96/6UX3Ibhbny+SWfqkmR9PZKQ9YDStbSZQZ/oFRth
5C2n9wh1p+3mc2Lq6QIHJx8HvMCjq9PYr6kJemkrnNeKB1RW8SVuEcDP6cE7uUW2XQ0XCAjXRCZd
3iMnTH1xfTvZR9AcdDvptXX30D4hNaGW0agLwlUomRbmwlU9gXybusDIBJD8QQR1ppdqRDe4GMiG
bKgnuvoge4L8WQmAV4kIsrZS+r5kZDqegYvbmiqZlc1fdnk82Hui/yWgNat3VKFwtX6fZ8buQ3Br
WwJDuzEjyTMjBaztTVi7cYShDnzy9PZEjcdXTQyKacaQLiP3KhZEMNTnAgxhlM01EdZyjvC4RTgC
C7ioLy+dF/4yxfTgUkTQrGASAB12VHRrDlug5cSotsYrZQwJZogRq2TF7ckpmsr4GTGsArC3QDth
wGjXO3fY6RRsST0SW4H1ndDkg5NNw0srxQskLjW1iXLJJO1reTjei0Hyb/ef0CDv+lcsiX1OjmB2
7R7qUqNPslgtoeUyLxSe2BcSvJlbDIAHRI+cZIiWPM6OkiEE0opNtzs2GJ44b3f84uMDbqzehM0t
wV0nlni0r7XoXnmTyffmJrCDi5u0YY7bAvJz9NvRp/TpfVk05uk11xDN9qR5vn+1ocXCy3ESaUhW
oXa7l6Zm3zOR3PTcJEEvfpbGDpUiffyiP1F52q040TtZQxPpzIk83jwDShWgGYgywrQVzJEREOzg
zv2Z/ildrW5PJe1Gfd5JFB3X5HJZpOXz+AKEJagDNpN5Tn75PVzFXempwM4+r2dhrVmUZXN43iJw
4Y2cIsbGSSDWgbemnqmOR04hB13eMGkk88qyWL+V5TP+rB7AZzwELN5BNR9qnPStX9vgzXeJP5R+
7nEty8NfXThUVHjHEQsTXFMHWlU/HIkKplfWN+OmA7X1wExsID//pGxf025016CKz1NtcW11O0Vs
meZPJcEY45Wi2f8GpWryXkABJN8TagreB9+fsf2kheamxHzROw3SKVQAioGnCeh8jExu+3ktsAsC
fkyPVZP3ehmRrXePhC9yWkwLC4DExofwRUtr0OkM/PvJE+Xkl0eG+gJ3jKZiPHZ85hht6Tkws6v/
Ieb1cojRXWZBELGxf8WzhKz2In9ushIaFZz1+ZaR6u1K8eHSYl64jQF26f1ijBCsGZFkmYjucMwi
lp1xCIOpDD7SIpE45KCSfhfYfGfxSaGb5RdplPKOIImeJ4hZn1aVvvooOgmON7Pc5IjOb/BBuO9T
QokuFc/ZpzZ/DsWxy59fmnjPgTCjuPhfNbQ9qngfDKkEKzK66TzhH6lLfA89ExHSFYK2Bw/Bx0n6
+ojyvnoD7ax6HRL+rMTIR2WrI1korytrkvNmP97LqSgCL+KRd4RXuh3jojd908/jvGCxK4CPZPMI
szIdSAGVsy+DU08NHEyRBBjfCxpCazoRpT3WOv7mbCnsFEYjaVosLjrSbHfGUQM+yZMqHFeoRj8I
eo4ObtKKs+B1G0nDIFTnEgSvI/QrCcMoliwFkE4msYGYq25kga3bxFmFehuX3qRXfYS15buR8XWb
csgu1l+cZskOWcjBopDrxPcwKZU0WJ5H8C+2MU+8kWgXw3qcuK2G0XX4iZv9/35Zi10E5EwR6wUS
OPKKqfSiXarI7NklqLkcZ127hAF870vFjHrCqOaRDi1udkWh5NTXchVrDqdvDAn85TRTI5CqnQTK
Cvxj+r9Jf35gm1iwRV/3RM8xKz2zpx/a57sLJDUeyxNVX2B+ByiQVxpaq9Gx1fWlWfPHgoK1Etr9
jVq0reQ0YVOiqQUqPPogDnK6TCeJiqroSW6hPU2w/JCr9JGKdDPjqiFWiRzkFgUwziaKo0YxZg42
nNzIHBrnEQX/v5nwZpjhtx9k9bR/6XqiTPcWUn50VH6aFAI59jnazX+DI+z/dtL2yqB+0fN6/weO
A4/YjeFIlcEmMXSS16qTcR8E6vBofpUDjyCdlDU+KwGPPzsZbGfGpJvZ6kwcfDqgJYRF/XsJ53Zc
9J6yVjXohTzlwkTgx0P6bzR0lJBZhhlB+ttFaoPw0ofKaCrDfEiM+FlnIPSTV6+SdTvErqjTXtn7
DOh9mp9rAYdV8PxCjbs17D42tJLkRjG9h+eB896P1hIRfL9qaOfjlVI9cvttQ9hJ2KR+i5/8DKgd
NSLV3xxqk5XsSZp8ji/nKg9byodgEVgRdyqv+2r1GVuOw7Q+cmyauneNK5rQ9IhUmPEM3TMqrR4b
8dQ79DjttyZr2qjsTf7K9LwMtxQLeDWcQehK/RtHrUjNbHtHu2Oxc4cDQx+DjzKv+HmI6QfbepKH
BViWHFKdHBXdY9DcGQUV8rLCp7Eqe6hC9AEh2j3uKTG+LBNSOpAVrnhb8+on3/6LVWuKhKlRa/0f
cg4Y+QSa6lugLkydNbEv0vDkLGA2RkonVCu6HeRewLDSIVMQ+FklxA99h2MNHGAJpNttwld/TGbv
LkX1PHYaA3fIiyJKM7BBHmIqbcDq3RsWZllW8CeupiOmO/jD8OogA0LoEYMamW1eM4ptze9xyx68
3fAjBvhhF79TmhEglhMUjkK7YZOE3G0ImP4YgA67/8oDifoAFiS8LOJ/7FCjXJOQHLTnTga8Kl70
Jpr/m1xc+pSDIIY5JiIRr9Z7LUOcpCixhHFwTNkTDeD7YUXoDEgpNlrJCMNfBp8RCfULOO4Efk4v
LzwzoRfnt2LTw156w5ISwmgR9vQGuba0NFb83xzYRKiNGwP+B1NDI1CD5U1/Jj2EcqF5ZsigxZlv
QLeTfwtAImw7lHfNrVfc3IKBTHq3R2VM0n/T1VrGWLDMJGq8kK3wXxM2QMpg1bP/2dD0l7CySiZk
RRFSQgm76dkQCNhd1cS2e2M8p5628RIsbVbyVL+9MROE0tJgev1z2xe9bEc3+BP3TlKlqr9gbsFj
dVBl/GfllXYDIzQXl/1EyU4CVbMeakY05QSdrpiQ8TPWJD9eHVBfB4/yAo1dl2KuUgSXx8Bg3wws
UE+dcEPtZ4z7/FeLgsv/gmAB01XzeZSJzw+9zmwdRwSKuDGIshxcSXA0HMgOVsJpc1tImCVbChQT
ka6mQ25RB177BLd8PHVoYWs8CIyHXn9qhCvLa22Kb/R156sC3Z1Wqtgt9t3XIMuk6pFC/1hmX/g1
hvaFzhT6Vuq5zbO6wQphvHsx38616kpS1XqvxFLcXqyHnh39ser9+Gby9CDWxD9+I33wdCe5HRAO
wu8JphMpoXcR899cw7D1bPd9Ubp1jY+VLK9E2KrmvrNl9DwrweULW+ghmKBvSxe/6j6mlRwZB03g
eO3Fj5HahoUdKAeiLDrFerpQQ/We+iAAKuBWJZ5WRroDrdwYLRtu7d9k8libLSmGevQL95ZOfeEc
VMaC7jtQEbn4sTI2x9nH5H5lB6Xryfk5GkJFuHQ8nKz0W7E4dA1j6hofZArT2xNuhHE96T1klNhY
4zgjCIM7tsNl6pwgXGeoLf+0rsyRiCUbweyvnkwVGCQhjtlwuAI3vC+Z+c1VlekwImzMaw+/KMlE
uhgvVLgTA4WvgmZExa2GfGhPFGvJWjZto4N1eL328MSGksdiDb2XxqdbPEkM+0oGTnmFz7Qk2SaY
ZIT5ThBrZTdNcv2GMazsfutp/Dk3IFS0Nwfv+wnCnYTMU4Lacdy4rb98ePVj3OWpOWRLDNwmXdCy
o/LxeU7lgd7oPpIl6KXOshjOGqFgwrt6eQztMEWtbHFgsPP5u/xCDPvy3dUXwdj+EvDXlwK5x9ey
Pvh/zmsCbpCxf3lLn5iRWwJaBa1camQRFaujWEsKS8YBaCuq49g92tYXMMSPssJwe77dWn+tAWVk
KWrxnHjzI7zEJD9FWBwiQk2KwLRX93Vh1fRCd/ZoG3lB4zyRvZSi3qpl4IqyVvrvGYnte5rgxdEI
hWr5ZwA+t6arZ01zI2f2bmGBTuIyTpNrTo5M94T1w4ZV0nokmZUSU0sAR2dYPK8/xdaZqMiocS53
0B936nhifU/hJ0NKoBsUU1KjX3fRN76VCZ89C5GnIwBwJCauROzCoFkoV6G4bu+co8ifNhmc5ysR
QxRHk+vyhpv0d32Wc3VR8Ndog2YkCuek0JG7+Pr3NoHdSpfB71criD0IAUA7nPP+5n94neZig9Gk
F5khjr446V4aNeN9J2FY1hACNA45m0RfPTXDAnUS+XvprHpsYFLtwSzNTD+rpR1lPXQXerPMYgR9
dl6N3ofFFTv9eAi2tn2ON5dHv0dKMXxDNnSGqBF0knHWI08AEOcay7kX5qpuO42G+1EEXQIgWXWk
LEFVWUPrR7KG2bCiC/Cd8xkWTgsSCvsbHwkOtccEwgPP4/VDS/kGK1zK6FKUkZTfXN/pDqU7OMlg
x31Qt7xjV/pc/7wij2Gf+ijAij3BguwG2clHi6VjtHfNDnZUKJBJJWMb0Q3JpMM8lwnrJQx/eQGG
10tGjI1Liy/wVmROljPJe1Abu28YJuiokVckXTsKYjG7ZGKsaetbPrJaXVbUq+aYQyyfiyR1EpH6
6ddqvECf8Zi9G7WvSjegKxyK87Cf//aHNGWr4rJ2qXibcAk1AXfZyOwd3MX8VvDRlBEahrzR/mwG
zwxF2viNBK4Lo0TG6l/0QKJcVXFOGQ0vqA4QYH3dDYi2h3EFWirk9TYt2viunpA5F7IQu8MO2KBh
5HRvFZDsIh9LFZoSWzB35Puo/ujeXiMgQmDwrsfopq1Eo7TXF8VUfwGsBnnp0B5DzoT3Ud2zbtmc
D6OHwzylHrckZ/smHcVehnz/smxfSuq7SbetPW/QHYnMECHxIBtpg6OHjZR9/OArXSy5Npgncgg/
XhLO6nNeIzNaIFArfY//LbmaB9NMc4HuaTzy0UHp1eZp5iT+LbmaNAqo/HrdqepOUmMgB6BAd4eO
r02m7poSUYcuQnAZyxhTFU1xmnEzXTb66T6q7B2Mba3zqUVJ4dOqd7OFXcRiibDavZFvwznYMPzZ
o8TmCcYxTJhkp73fjQkgLDHcYa55qtIIAlJUR09avfRiNKwyUkt04Z5GUAtpiXQ7gCbKQPetdXT2
nSwgdD93hxskTkXvIsEjlr2GRzzG4M1a2O45kqhYaYbpHMHFoDXX1ZzzkJzfw7hmOMiK5O3oP4ki
cpWlRa3Vnq/2v6wcZ9PU817rw3JoPVX7iV2itVgxDGozE5GqvF8tOQZlIKshheGEC+1QTA0cuZkC
/8U57Zo4Ay7XgtnUVTMLun/UCw10KIPEwtGcj7WtjgNIrJw0IDZuxFXY9CjSZXzM14CNslo7eHiF
gm819XqRnjZuVrbnkO1oc4HNkPSugv1qw1s3OpIdxuiMO+zcHd2CCFmFmQ+ouT9uuZIOnPcrVWhB
Qyb80U/IqtSMfDVbGbAqSDYtV55FMXyBqN8/ovCB/H3nMunBmKITbyYP3jfwDgbRAVC+yHiHNC5q
hbtby5XEoYDXWrDPkx/mRx6ybl5TUWMSlgcWP47M28nJ/hlkydVVhpGGRcjJcMFE4ik5UHFnE8Ca
7/VLxfde4PHuJaPYUt2NbgbCoMvkvEldsfew+ICmw4pcOWskcuxM1MLJs/ne7vkHFatwrWgBn0FH
7UJyBTucMchYfMwRdCsgbUEMpmjZnm+8W6GGhZQ4oi5BkQ/jcjyW5M3GbtVB3UvyJFeoBSCYMzhd
RLPgRFTwYnliGNpl1WLYshgpu/Fbdc2wHq4kPH/CktAM0WVYtGcCMHur0TSb3ZK4uiOvArLC7lvd
LPhBD6EH0oUWJGB6dh/7VXRJgErAsIjTWVklmKLvPSWZY3Et0IQtzQqUOkbMsbie7sGxxg9IydLc
9KXIhER0TAFEGw8v1kTohRVH92w/hOHj/QvHdFtE5WmootK4IbIpIcxJiLwgxJyW8r3RQt/AhnSW
S4hSpEvKB6QhQIm/5awB92BscFhHoDugHYH7nAW5BnOQjHJW3H2BbFsit/1i2Ac03zm5qTtsaRZX
qsjYK28KPv+CJS6t05jlrmqMngnebMc+FhWzeWYnvqOkIs7LP/2x1Ws3m+11WBlt5YtTjdqIy/Tk
WjAmMStnQcpc7u1bWcyHOoacu/5EF2fraSobwerhngBhGwywvNgMD9h21S5rur8Nyv1ylWVILD2d
2zgWF7RgK9r9shO/TgNTJNEyBUs8QGJrsCSMVuz6nd53RnMdXCvo1egX5AUEIeF2SKIX3EuPaUlj
MNbt8jKdCVmZCDqWvBDn51E69FZOXMK6LB1qEfnn023OqM7F34QpCyBkdY5P203+RlQUt9eu41cL
mmdpjUvXkpndYdd2xjvP7BNqDR6s0KiN+GUjHVaJtMklRRmcIAMpFY3hvysS6vOSMBPtUbNP4EUO
mbo6fKwkm5mBqjFP/iCbBIhWtAp1HZNufP4Duh2ZgihbjT3qquxvYFzx2ckQM60dNTZTKk8wXDBC
spj3lJRH9MM7v7hFCTAkBS+pW2cBKkV08Y0v8GSK0QpoGB26j0eZKchv6P5+49rEKAGtfuOGJAxl
f4ObM+nd2VprQiTA5JGhjgSFOP+dSLe1NGUiqA1a5PAAE2YWghuK0FdSZLkjAmfYBUHN/Mkr1rer
FKJpAViE7QDLt5kQehDCY11Q6Xrhl3RAuoZAxVa6GGjj+Goos4K4f1BrP6XuG5yeoTW2wK0lpi+8
OfpvF0mzNKETbhUjNLt2NCopvay5Z4glzbp2sJ/jeONSVnb4g+EHr/QzzesYR9Jb7wmSrPcRFLXN
8xCtIOG5Jl5uj3OFuBdgetfDS4/8VyYIJQui7sE5XAOI+UPaQ2GL9zWeHOv2Pcj9mloQmoanFtnf
mGgrA0omeXNZ9NvXL8efIst9wcrt1tfs461n1EAvegkijjA+HfwMDflvg12iXQeqrpbTMuyQQtdj
vXrMGsPy+SkWaTM+k/zGg5Px/67hMo1X370DE4JtrJS8uvEiK7vsER0TkhV+q4gWXcp9r0cf18DS
UC0FL6NYQ2DPAYdkRu2CVdOhrj6ZwoG1h8T8Drey7Z3EnIcAPhIqngLUoLURycQT24N0kzHAZz0b
Lw8Fd1kinH2BsM/Xr9QrIeqRpqtX+V+e7+xL8IWIU3NcLLGKcgfMAnZi4T7lhaldZTs59zeeuUqq
gRhKpxIFbU2MErG5bxarzW2YXyeccKo6n7gMPnOWS7yfZfjryhpOlfoKXHxjjMqRe2ogALfucwq2
OMtpec4WGTJ1ZYxJK9+vEFzGTjj1yNOpOOBYxCwEgoHrR1Lv46VPVzUVk50YWlt1Np3fSc7GQSKn
bIHXqojpNaLD4nZO0ufXPanmGCKJ+yWzgQ1bv6WBjj3uYSsh7nD3mIka6/pPo1wtPSBxcIS0iMH2
SOkUCbH4RbjFmam7h7KrRd9zidd2sS/utRD/n8pJYcOqhzIR5kRc4tJSFuYtEyzK9FOuK5MsK27J
UCo+6j05mVb7Pxn2KgRfE7fUGylRKHH2Wc1/cOYp1p5CSjM0QGMvrobJsmzkhzRprmM40ec8+gOo
NbgtOHCdd4eLX/1otn/bzK9dASVopcqWDCv5IBMA/h/y9jjrXaHUuyYrEV8cTauHwJZEukvVcNSQ
/+F62fsckCBOhRXQm/aXRARBDGeewKw4gABIef2683HCjYjNaFliQBsig9JwjLG09ffWYfMuSKIE
xH3kGclerDZOvahJnyWFcITYQe1P3C8UOqLjcTlr1rxletWnCtEMeadua/HwUVAPpwWA6Bgk047U
Wu1Ah4AzpLi117ytY4ZUp85UO4yuHfeitM2fL3EFfrKV6eBvh4m30x0jTuFLRrevtLeDk1k2kx9u
slu5NiRhQyXa5RFlr0+4PtvFyweWXLK/W3N61udamC0s2XJVUIbwkO2qv4i7ccNJXJnj94jXc9V+
KYUWCUqFT+AofLoOJwwzLxggivBT7XN+06SkfMuEwp9b9r5Y9m6SaFUqHzAmZhOm71G1T4HNRIcX
BS3BrgdAj58+fXsu8JJy4APmPQ8ZRgxLNGP0vix7pVTle4FSv0LRMmoH73IOhQQ7R9SnIxnkIgfL
XcnCTffoPYyQ0CMzINu1SNciZoVGicztC8VyJEzcFabJTxQ9g52M+LdW9XmBDgAhbLwH9cLKLb5f
AfUU8HwWEyhjrRejGlSL5cj6Ni2BTPqEIvVfSQsu5xrNmMvfbVFxI9jhX1tJyzSwEtKyFgsNDSPi
aEgxHOyAWdFtdRmyFs9GRgXjLXgDPlcDHwI96t6AzyWZRhfHFVqttkgSSEGpe5FRGkY6ZwPO9Fc0
3NCF3L05v68I780WjOvxQ4omckU+Xw+VeziEZ1OCXiCHWfgZzANJ20n36x+u40JBrQ4lEEk4hCpt
c0YXA2QG+Gcd4YXF3/vgSSwBuwO75RSl758v6+3LgV5iHC26aQwFZXJsgJachy4fFxJdon8BVuby
I+pHwT0c5oTZNxWVWS66Z9ZIoR2AKsI2M5Z3s4n7w4NWmLGdTyg+M1EsXI/63332jp25W72sYrB7
Mx5Li7CmFGNpjNHt1rziY/DXbAibVtdJ6NTCUC4attIduwS47XgRRqGx4ou/nEvcKnSqfK0xQjjZ
j2GdbxToroQqcy3J6SyppSnmi2myJHoThwVmeYh+58TBpmEFKcDPIjfBHRX2aOlliFidFjtonIr0
IjpGO85L1fWOUr9ZuQIlXlO1Z3MySJMs27i7z1zJwaB89twiy6sArcSrsvXcfNopoa6YrSoZcoQm
6c8Ww8B+gZ16LjKqHy7q1vh/rSS7L6VDgDB7jzjGEQnrF7R7Yr0TyC6MAnYb034SH+VHDxA0kaRO
IViVZcxeP4qvGHsNQ2arLoIzSQIFOGGFpynrJqjMk/bdRDufgAomiRCahKfO18YDnciBlLTeLrH0
t4PycW0oyeC22h/w0vT8Hyga6MoGfNJNaTIERRtF9oXch5gqbK+JDziZsHVXUgulXzzFU/UCIiBK
tRz+fka4LFjHqy20BlUXTOHbgGlBE1+1BVybldNro6uFl/ndK1IFkc7WXIk3H0mOHtgwn2McEn+Q
SXSNCDiZQ9Tro13Tr/mKGKY9CnRGQJL6iKPzpF30FPJX7R1lWQrUwT0SDAS+lUdX4MqllPHVJ92r
kupzzyPzBctIW9GNfhkC+VGbGL1/lVAgIpYEpXL/o/uQmY77iLztf6q3IyulAtBskgHgS6VydTxt
qMLzWEmVyEH8khoGWL8r+KJMf2B4j+HuqDvZQ1DMQicYCl3AeqG0ns4fZjYQzml8007pLgmEclz0
klKnJP5O52KrXvdVMJEcV0xV3QRbt9o2aJg/GlOb6nK+y+mY13Tw2KKUJm/0iwfSEPv98uTed5Ob
sO0WRpK1SKSg+WU2Ku9JPsVQKqmYNB3TZ+O7nIcTV7T/XptmaOnMBhdYMAhY91Rg9KOhTO0X7N3v
tJqVjNtilDPpFrYmF5JdLXcf4EqI/ZpSS5lVH7lembA6wLPdBI8Jth+hF5vytj0nxEva9XGKXzO8
b2oSOCMFyWL8RAOIswr+0Cs9i0VsGSsiEdOR6HcO3Vny980fA5w24k1u7Hn0m4esbBC6FvPqX14I
51DJnpX8T95YpnIYX/C7lLz0RgUl7akCaMwNjmIVgCEHLZSHkoLFPrd6c98mM5gG55o0/xbXT+N4
AZhSD8xc+F2pAY5YGt3XyIEgLlLLk3oSVAHSSInat4PNOpAUJpzHS8b/gHoNUkBMigcqDxruF+Ra
YQsfE6yATud0ZqwEWBrs2JncW8FvTEzFZANJ2qXi+fd3qU5wPEs9u2T+ZQLjrod9sPH8oxr+Kqv3
5MXZ3DYbRviNE24A4v3N9kd78x8EBkHBegECHzGtoNGSSp2Bf9EwXtL0oBhnRLmygVYS7btJIvpy
LghuwO2JH5T2dvqmc05NaWmyN9GOTgkKlAADlxLqs1jOYk1OAqOTB1VVHcXyj6SQaMEijYA+XzNd
ZHke2UQr5IqA8VKzFlKVAxXs+DNGUmpefFt6GD9eaThEA4EfRkjqSCnODtm+ji5IdWKQi6pONmoY
wLny6yh6Oa0oGe2PxECKMW5/c1iQSZFRrIsathXqFdJkL7glkvb99NC9OtN9LQtrNc6aOANm1eyb
RjjZ83pL7Xfv5Les0AjRvPzdJ/LXkJJqeDN0Y028cFT5BNE8SmIvaje3C1yDJWwfxP/o/MV4vCbQ
ehcshRUTMOVw/1y6F2Gdt3rJxQa3phs4G+aE0uPPiSBuTz8JzWIXsYP149pITeZknleOfuHP4z7p
oUyuf9ZAc2yZWrb/XipzoqB10duk11dd0QsrjmiJUB6aqiX5KSFVWtae/f5eAD1OCRiwe0giOz8N
frvTnkv4puOw5JQhh3nzMfcUDAMecSkmKB+uiwgrlVq7pfuC/Zx6lI4O0iceKAZ+VsQMCLcSKVoY
RdSfxoSIgBv4aAT2TG3jqCKdHZ1CBgeGabt13Bvoj+bWADgEPc/luIynCd/rRFTsUnmAGSTDmUgT
ZjIoDo3uWWDPAGIqJWLuXDx4FCwNTeddoU4XuKTkUV/Dh3BjQNESKp5orYonrTGtBxHBSwtLQ1WA
MnUBi7ur4LXIwnmIyR6k+PJtCQlYyVRjfvT4Tjx7sLfXwHkirKy8M9F/b2bW2YNJlOL4HtOIilFk
tnOb9sseAsCtK5bm6lRA40q2l7cCvMJqKtTGmSRTR7XTYa2EnJAehIwxgvTT9b6wMGszI+01Up5W
w96Ji+AhagaKu+fBOdSrbTIRxoRnaE/hbXGXVfONqUuO28Wbz/UitojQNsr9Osn113CpER+7ot5m
5keSI7rcmJ5ijGBun+RGO2qH4G5EBhwoSyhzOKHVW3brwr0QShC8+AM/P7DbYujDvdcQnc+kLdMV
3jChzaSosAdVqEr9ZLgZVGzEzb+e8+UY/D4VWquGIw0kdMlmFN6/AfjTh8urxjKKcs7ixGEqEctc
9sgkVHyIvDx4mGwFM1vuhsMJoEzK5v4BNCSSqfX6ifgikh8s4s/orAt6hPtcjpD81FC82Bzduruj
L5DFny9EnL89NctWHbcA236Lwfs/izYgV8Oeno8RQQGKeKQH15Pwy/I2qaZNeexL5BCq9618g1U4
TKF5TQtWLMK0PODW0NHHuEFRMZu6JszDEVKh65EBFy60lkYf+0YidnfGowy1HricOmdhwvz8vpcv
/WLb5iriw/ldPzy2ZGwOcLbgMSKEw1kAQBfAf7hLmsa+OeXfXcCQMK9dkOD2mfRgaIaBJoVHsObM
RDT5Bmj3Lmka7qMwsmQJ38YK29PcnYdfZvtJAFmiVlF1Zp1T3cN3Ds1LAGH//L1fjrW06nUkl5sK
6F04UpmnSL4D5KI0zWdijDBo+dAyi+8ZYZmTB6g5IF7xPQx/OSl6oUQtPM0ULzqou8CzclNn7pBS
HxAMuyIb+IyWOEmQmpX/Lcr5DaZOwEiYY7cNfvz/mmc1QUHKANdc6Hfas1FdLxafTM7oI6dkNKWB
pwQyTqhXo8rpduLHYNNxzQyUp0iXHcZPGT1BYLQ63o7DzS7Mb+LfPR0shpY6oOPnhbWnjfK2TjIX
GKK7fDsK/yzLyNMhjUHncJCzv9c3gH0CZ9I7HZxUv2GiNTWWw6ILSW744YelG3Ka0NbGNEYpPeaA
ZrtriBnbTzZjuoPX8BYSS3q8bmRJxbVCea8qJuO75x7wVKY8Q2wZMZEIulePgTpvFqXgf8rZQqzj
JSvd/7jW/HZY6bamdeQYeRACUORi2TpXciHW6Tkd133p7Fkzy6jevIxQi09NCunUMj7oBQHZR2Yb
Pto2XE+7kZziMRJ8O9PS/nHZB7ujLk0yEjWHDgWqbyqkkW1/0hcKBW94S6PZ5OPELL4KpMheKh18
rbcPnd2DUjy1xJxLL1o8S/f4HSuNI79+EOG+sFSGJtFIcYBwYPzL1pVCS5DfHyvM86oU0OwyTJKs
n8p0Qr3Ma6Q+wmIXHi8IaOU9THVvFhavlC+NjWhuFem7cE2ft8emsx3iM735o3bONihlLZLhwgIK
sv/ngNXykfp08nTmoPznAXiDndk9C6B4YcNES+y5ZseC87dQdln1KATJ/KuRAGb15cnWmyLaUJaJ
DFIfeEgqOAKwHCKzOdA/XXQxhriVaNwBUS9NRufvZAgSDEnETTVgbJ/WgSa7Ck+O9r2p5sEZ9/Ud
+Eg55eADgZXYW3pNJSRS4NuUMR3stN5Bj8bHKcu1LHI9idtvcLo1Lf7hiYl+PuAyO6i4SgJ90wxN
TrFHldSP/S9X4mC9Nm+X7OJW9yWuritS/68s7qyxrBMFdn1cvQnPsdAqiQtixxrjskg2EmHg5Ehy
XO+6C3j6kYvffwmv9HXpqzx0DnHn2YMWm2RhLPyvzr50JOUo9ws5K8TMbM5En9VFlD/RPZVOUvJo
bX2pbjc2DkYAfrStV9dNRUqeIdEtTruycuho72IMJMLWWRypafnWR5KzZ0bB2W+LLH0LKrOeR95M
lDLzAow8QZdUe2Iv4ZsVMyHEgNufLvT484RYXKws+cMIIMm7JnoaVXnipLXimLXSNZSM2g+BQ49+
i55IeUcWRT6/lCUHrwIZikrJBz6+20KxBc+wqKH6YSYjgipgMZYGPOhxAUtzUzMVYqms5V0LuLno
3fXMbVWsAPBT2MBUSy/pcedkM08i0t+7crXTPvnbrADaFN6/KtXtv3x7tsUVE3yHYQUp1EtuhKAK
eLTMssXDm+C0r4izPYGsM2fIHVlzjWM1QVikrzNDbw2e9opzkF2vmn4+19NsmJYcM7ls7FmqT+tu
ecP456xYvXCESIfzw220W412svWKoV+VUmVLpNvSjjM4PhYyVDn3Vp1EdxSzX/VL6EvmF+15rQlv
UBrilIdkIA6CN5oQmC1Bi/h0nT1NfYb78gcOCchVdDjGMnsl1Jpn4CPr+iypS6sB6mzc9x9oRZ0Y
ZErehnD2t1gBCKDHz3ZkpRGiblJl1a/NIbUiW0G8Xd3DY86c6gvpTRmDiR8waVZlyBvtbNrWS98J
JuxaCoNv/svithHhimTsCDtV/1QMubb/GJ+ZKuIxeDy5sX1HHVEEwsKAx1I5AFAh+TX4iwX7gKii
uvZgqaN0v43MN/4IigOHGkW1XnR/DEBoHyRZxeKso2e2/vV8EUvsn747DhHdFJPaS197rHg0Sari
gjvqSGQKOh6ZD8h3RPO+xMG8bViEonDV4xFPyzlKOi1nm2GqUrven0W0Uq0nS/vAdmhzczoyDgUa
MZB3I7AU73w7dqkjHDPkpKh5LnJuF0eRTvuNiodaT4Gtwplad/2PdFGjdKSDeC8FwACaBd8eK9uC
xR4ac0pkd/joZE0N9VOOKUz40fvnFiRAw/eulutd4SMZxB0d09noJsip8Fgp8Z4e7Z7PWdSPZ38j
w2eOJo5eS4lKSmm66ftXfuDXBehhoOLJC/pjKxVz4z+50Cl7X4xrrJ2QUq+2n1SZeRh8C798Uek1
2FMaX3xypBxBAXuzn9Mmbbp1zwBU284TgWErwFawj0WYXKdfuSlCxejcxUl4g1/l/y6Wd04nTqFJ
MDJGUAtJTcsDbB+DY6+EBNYvMXOsdjAgpiiyeQqvb1wUoe6hQEGgEIlfMqw/bYk83tcoMSFGN97A
2D45/iTwAzCouAeFr68QgrlHEuuDwuihl/rtWT9wNeSSvZYaYm+NlJ8EJD6fJNdCoE4jzlO8x/EL
aH40SdOXukTG4J/CtDPo/8hj1j1hVfE+CM/07QbUcoM+EPlcgaRDIqWH1MVpuqe0oof2cwwIBQIE
PwUsjl7RYc6p8b17nTwQJgPMptCs8QFkS3nZ0Qrf103TzffCgxkdR9Zs0K9OUIqcOVgLBQiF/HDr
gzRBSHlG+oYz1YHPZwZ29g4zPG4amCck/+zJ1m4Gj2bGgUNE78p+VM+nT2yTr4/QkiRMXOBaV81q
UeZClZ8sUHpLc0wfmhlpIOzNo9NjvM26iDXL6HkvJGreFbACTtjlI5a3BiWGrHBFBk/jFiH0M2Di
JtWzGntjkqUGb7nZJMqPX023ZUjEch9wvAjq0Yhn4UbEfSG6Mow6hf8iG/ic5OYg648o1E/Hl/XD
HLwdOOqVQJLF8HNKN8XU7N26YgE/IHFR4cMvUc80zlreIBehwVjXmHGRU+uTCq5vCclBMrqJDilC
UFT70CIAJJ9jo+rxCrC9h0UeBieD/mEkyhLMGIceS29rhydh/LqnXb0kqPX0l0us5ZM40jekhq+y
arc9gUHQqJSn6c7m/pgWn80u7sX1oHUxX5q3QEdke/iFizVgyvf4bpy3uHMGEnqVw42svcgRhfGj
7HkDvydXzCjV2YTaSlqr7ShVS/Uabw9DudgTCYTW+iff9/mYNEwA2zl3/RDkUbahUugEVMSa090G
TcSdOjhil21vLPtyC4aIcvFFPZkLWag/EsHUZN8YFofoh4Pf+KG1gf4RXRUJcxDTeATtMOrJ4R/C
sZWJcUeXeJy4rGHY8w2pbesIxQS42vYU6JXWk60aCDCtQK4ABaMJgSUFnhW5unhd/C3HFGc0LDcA
i5PXl3djgoBLPhDAbP/1hjsega7uT3aA4UgObrV2iNxwl/+L30pk9S5C626yJLloJqaA3jqDzmW+
37MWZieFZKOLOB6o3ezqQi5LdpMMrDCKZUlofUYzJCY/KFAsWuOiEBUE8rFGimg/cUVi9M8dXRA1
z0lezFyl4e5a1HfHroQAsGn9nfcLrhDSoHpwsuwkev0Conx0haWjFvOwOxgoZls0PAaDGRl0t7Ln
16cbP0xkPdN3ym9ZdR8PIOGc5f/jFgPihnoOVwY7wARSEVmyi0zsL/k4BAU5BWfUedF8VmVBYi98
UJ8dkaCEWFMiUsDWWnM3G5Cm9tpNAChXAbAX/OuxE5BvRfbJEOMhiB3Ad+TkpO9kVnYwsAam+JoL
/jD2jA0BOtUeiTOJ2PF6aZTMgu7AJBlQIaFz3LFkXRvmqtB0jlVYaC2mRairBggrk7RlrxzB3pHj
aFoHDn39DSV/iKo9WkU9wPz5GY4KYE+L4aygw0zRDQnim5jydP9EVEco1GcXVDOrdKoYgcSoF2FK
LB1xJWJQSuGirJVzLnxtxOo2/dK3C5N32c9cm+mExftW/Gc0o6SFKVmOFNcT4+23C7++e6LCUQYb
ITPbUWLh7+7HmHc+lFOQ3zhJuPJV/pD24Vyo6jEN67eR1taMDa8DsTMI9rzYcDaWZHhc2fEmiaVh
8dOBf0r4mxgBCcxyT8VAMgcXL/O2HcggJ3jvg6dlFUTSHXw+trGpU9Pnq2xP1rVLE/kxuI6Iz7c0
WolH8T7Q2ABxTrcRHfx7YFLOUXxp1OtdvEHNCrF2tGd4YM9owDeWZ+qNuzZF9+Z2JU5MRP+nN7Vi
ZiaSptYHI82RicQ/3yQQ+m7qRfKWlvtmTUDlatb49nU2L7RBZFKdlmd+ZCC0Sy2bp4lneuWuWksP
zq1Zp7J0/Ue/3A1RIL3d3TLKxvv0eM2kLhIfK9kPcZ5HxsDXmWM7lePaTMRYmV9g1Fc8S2BAyh6f
kiU/nVoJkC/Qje1NyvYWlwAlxvTM5nQNl4XB9neNDkaan7GabpFT6EHR4x8l9P4rhRoA0/yQ4sR5
ajb6vaaPKWEVRGYwWt10ZMoVVcbqF+3aIIC/bbhcRD5UVmEfrQHOOJ8HUPKqEpVd7ERgfBwJy8iP
C9TIHOx3BX8/sGoUuVbYe5rkc4t200iahtxxv8Slo2oq9/hyylnAdwz42ZwLeNoUcGSnLXZC28qq
3rVKRPpvvBY5WSGeCwQv8wpSismnuTOIDxmdFexA/kIumeCiQnHF5ZL1CKUw9FvfREp3OBhFSzRW
+fCbmeYWQ8JOhI5pNQbhUygzZBAOSpXAjB3nWIA4B12o0xVdBJZyUwV/fXkbFZdg2dVbzNVOTV0Y
YafkVmCp4NgfO9d33kcnXS/P9oxDqre3/+ttKC8NZn7IWdA9010qz2GWDDwA8qMVWxsbp3iwumnS
KzcRLZ1IAeqJEkgUqh4AhshfBIOsePCrN6TDDrens2m+KiC9OMLi7y1gFzsCOhkr+/506ulTdcn3
fpkJsj+yCtH6Oxu2SeW9iDJj0ZXSZG9U+d1q5DzOL+LxXARr1yjyncDYyTeLe7nRPgOLxA45Jnah
oszD4tdMhYBld3CZG3mpVI9zTIcd+ZzGm7T9R1ug7RbII2QZnW2FzP77yOgAlfgpwg5aCOuf+awh
kNGtELjoIQMnHsnV1A7yHFc/qAOcuYwfOj3DimK9mAy8E68HqaO/JETbzenqwz7cJ6E5P0yaoSPj
4ZuKW563HxM+T5fyuKp5g4Y0nSCS/ITR8Q/4kC4XkSEUKdKs6Owec4lgJoiaEpSVz77rsS9q20ad
1oGjCaRptkOkDKKgefz7b9sfEYq3xM7zSvoFErX6Sv0X7IFYky9+LU7btIo5KfuRgc2r9xdc/pLU
vTWJ0D1TXsU4IcvsXwDxNFt4vlOsekgJm+VorvM/zd+i7vJGteYrO/AZVRSP4PlYXlj9tkFTfQyO
3cikSsyXN1O5hvX0H6x3XgxnYFBGZrLHRsvPy6tbS1cLv47ugk3EhHRNUbmyN+UTu/0hxeb7VpmC
+iXT0RNZC97mX11IYea9uVH/TE4Blqdbm6eiu9ehQliYMnIwTcWozES5DLRiM+GTO0jwPHfCbQq2
XFFl6D7rfEUGsktAE5eBc2TcPyMQddhVmW3ZknwbddFPbD4HIyzM37k+d/2JbBv7yTXx+PG50Nei
CxB45mzf0AvGmUEXGFfwvAg7131VIryOc4TPnsKOt5P1C7yuqWcMiErxMKMTgIBPZhyDG2HwWgeD
CCZeyiRiELUykmxaJZ1+3Bhka8EBfkDvEJ9pp0z48PfGfBwHY1DwDOnbFKpOl89faxv5xbRAd+p9
Rt5jdJ5NxipmN4E/ker+Z0Cpc4mctOvC2LGCPIfRRsgV7dF5LO0l9mZxBPDnZ//leIbHtz+M9mO4
V+tsLjNacCpQEHLrHBkEMRGThBjhjAFg7Yuy/Vl7YmhYlusnz4oDKAEF/lU36ENqrkYWFmYaL64F
HgRdz1r9h/gN9JN3lAqOKe4cNGeR5QDWjmv8yI4e6fL02j+AydKqgF2zwcWOjoGQF2vV9srsvUEp
3CPXPX0wUqD5lFMQpjrhRPHBUVTdgCmNUBeskanEC9PW6y4qxnBRyUYaCBaV5AzeJ007j3MNVPHD
5jnNJ30B2or7fwqFNW8nWbdljkFHrbaEO8ZgOp2nhjArGkUy0YGhIPg4ikJmgPf8ObyEGClMSLQe
TsG6+4JWzAH8lwX39fKtSXTNe/hScwZVVlIfUcOcSybJCInxFao+raGd4F3HubxOwlda5eFR40rX
23/y9Vb+csLhpfxokrA81VuLP1gavZ8vOFBQJlpfBnmbrneeiImqRc7ADNWABtrUXe2z7o0ZblVd
m+KVOieaS94k2QMC0DJMhPWU4uqeOSCPuiH4wr1/6ixdGvdOsYoVWX5pXFMtW6A4XAiDAmF2H5NO
PrHJvFhrZngqVFiRIrugrCxo85BPFtsZkRTz4lYnwHJbva7sxwsGY+/cJV5TNo/mds4NMlaY0Myo
71h2V0DhXmlzmsAUDJECK7GtlBOCZsLRh24N47KlWD78qM/HleXWgykZhTz0gGLYMxN5C8BTQXBa
EGjfwOCVtac9Wd9su2sz7GaGaRBOv9iTR6NDNfevNKmSRAfMmvnxg6PYPK1ESRxGlfnqF0av6nvz
4llNJrCISdnzjkkarrY+eNRAw/mDUm3OnmSKOrVKJw8vVF/r0XOzfPRPhGA22E+CKNzxEHLYkgvd
aW7+/RAmTLsxSY6ZrOHVnSDsGoO6S1s+s1isEwN71bVsi/wOQZB2gT8zDaoHSmNgtPrLc5qbyNGG
NLhS/a//3pOJ2YW133CxN37+yVKp7mKwxHTXJRM+285a9D+s4Q93zmZFT2VMHwP57ZQkjx/qFHKq
dvPak/nAKRDXw7Iqa0fLVgR1Ng4bKAKLPikTGFWq+2/ake2sD6ykFODSP4uDBOm7dKq3GvcrG82m
pqyvh+LM+YgGAVpkuz/dVTrj3r5NMqIYEV23cr5LFXqO7mJf/91HZTW4+QWaTcTEE7VI48A+GgmX
GgsL4vbIUSxryh3lyMxzqMW1wMABiqhNJiGbUdsxP+hfEva2w8z+6wQSX8oM4vkMIFdBX5Tz1beJ
+0/CStMX+aS/5uZfh9TLmlQR83+62+rNWIi9nH8KELmY+MLUn8uvEPCeE19/q/NrD3wDJ3pbIPvE
XERr17XF5CGXaPHtSl9S0rx32YRC6ATLLZZ0NgmjL++4lZ0t9yqYERWip26B4ynSGF7fr8jpbaOp
0JgR7zD/O1s1pVZ4Nt9+S8LjT5aHZmw/u3FIzSptZynC8c3i1pfeiJI6z3/ynRqft579rQdZqHZY
5Ywgz67z2mFNsYmFnqGwUW1UP8eEy+bP3s0ob2HPFg8BoZlE+tK+VsP2h7qB4tP3K4FsunUmnZmj
1OsQefhGoldnKfQ0fUWhOzWmgx44J5f1OUthDHClAW0mZE85NwjKhBZ/JKmn5aeyl1AzeBCUTQif
uFGek3aZ8iZkw5ElDI+2m3Jcu/XZrXL4vHleK2ABU9lBZ2L7HAgW8Ol8yjjj3/kvuFL7IUcK3Tzy
Bfjd4IuDpxSrN6anf0oQkZD8yfR8DN/8dDhWjWjwgRHS0o9TO5P5sR3zNYBkPmN8YVQj7WXhbGkc
dLn9UdDrr7uYkPe6AN9usyH0gBbwmMdxplXqb5zyeNouHmzGCA9MHatNYUUrggsFpxGU7zojvEdw
pqQK8nK5uvdv5rwM1Tl2acyGS1AZoWjXNsvSwKew8Z2vpCeLNtKy1/tsGFnHY4wu4xU4EOw20I0o
+L+PP7fdzO2E2T5sZoIa+D8dKorZmJQJaLMsStDiYvtx3Yw1a67Dwo0KcucNXqYzV/v1+FRE7RMU
umFJIPYfjJrENESlTDdL6PBkt3nRAInULtRAbZmbersGpyi6BWpmhC4ug2t0SX/4373l3Tq9hEAl
QmOp07cTaB9OlYK1dN+1gjRYpPNRCLjBYEFU2J68k8SOwyQwdDSvqwbjCrWJABPlOOnF+lGBknbw
jgcUxjBBRFznrq9Ha4ICbqbFH/lndZr1dOBgLpiLPKVsAP7fWHw0TWzWtBxIXCpuUx4i2Z3Bpl+x
ODvxc8lvrJ86om7l0sbPVnl0JBeh9ORLs4/tWWa2I+Vv+WzOpa+k+IEycdw0UvhYz+dsVIscchIR
SdLb6Gty8ebmcfg6q46OnwPqaQMJ/jpLA7A+SVla/xyyh75nA7jdJjq0LRmw2Ohce/0DL7geL1Ew
hMPxVCzKGVLAaPVjQCe2C7dv7ecsAkBKPUuF99NsA6F/XZNGoY4r/4W93AxlslBE4PSn38Md81/J
q8L3/+JcxlKRp7EZ46Lnx4QklYVYzNBqTn67L4+XNoNP5kj8amxfgiJb9icJQJ/NcaKktIhW4g6I
cfk/UuUeC3r9x0TcRYuP+9sgwHhxK6pW6C8qhtafc/kyo6QoGIoPpBZg9vnvHM8cZupidK5LmOMS
fStnsMUYK3tFM5VZiUFDPL+poorGZT8lSrVbLi1Bxfg/VJRbcLLReuupqkkvKrTMDMFqw1lyCAkq
dY9+X3rWpQn+Q79aN54P7qo0cdyVaqgMIK08Uov9snKCv0MB1kWfCZzyLL/Ty+owAPThtf8nEkzB
H87JC2VpNUDxDEj7P2uyaVLFiykOGDo+m37BStmWHeNhw92/ztfa0SWcPSexAcEiWrpfN6CB5YYz
/KZ2KkRNCIeSG5GI0TPT6wXieXNt51wFPuA2EXn6R6qwBgBmqJpCms3cyZPboQ/fjcCqQUIt65Dx
oLQ8Kj04SX15xPRCI9FXywv6TP4I2rwX4NAR4qiM9juR/lIYr2H609Z8O4uSloG7JsUoBuAu4c62
VPN6x5w0KYFOMi3Am9YXAG1N0QA6ZW80jdKVc4HbYf7vG09Fu+kvJoBmbg9BBTA7R7hn2/dtBiLn
gBeCQsJKpOwdOHgf+W4HgjTHD7ZB6L5bdZvIFhwFeRPRpyOPXn0qgJpzJqysrN9I5nE3hGsKbO6P
hAyaRCiQ15SyxgWNfZ4TuDU1tTP9gjW7yTSNkL0PIwBgNMbhAOc38ydvPoaFkdRVGilXQyDiL/wA
yzGzvQsJoW9urrJD/DnAwkdPmNvIxSIouMFyPJLcuo7MK0J320Hcz9pLGXbwiUzODcJVpy3pHcYE
NTnyy8jGZSZ6iCnMwMgNujbgTHcd4xZV5Ix0yRA6go4N121h1OmT+GI1qKStfOlmMWxKQZOEbpCq
DfHrFVRxMFus03G/HsTHLPxpjCZYLnH/jQZ+JJW/kB2pfbj00KyQnellIEX6yjc//Jltehk4s3Z/
XdRYU7OKyZWHvQvxKEGCvPFAApo9eMBrwInK5qWqkm+Fxeps73BQEWHzWAhKrPz3r+e8zSLOAbhi
0sTviE7zaY4dP9CUZyoPp2ng3h9ok2cBqadkA21tGEZC8QeVj6Fcw991WKW19E1I51eLXQ0ZaXog
EgDxKP4SslD11B9CcgqHbeJ+tbrqruWpqfC8anNhTNuBYW5BIu8n8QfJRMfWpF9Sa8WCLQwGZzhJ
mDun+ah6APlYgX2P29xcFXF8JDn8neUaIttN8ylPzvnnLeG09ifURuo+MIIM2fMOLTb3Otrcs05r
Y3xzmMoT+EZzBmiWCOTTv99Jem10qZJY7i/NNqM46PiGIK9LCtKzWb+E97spZDGAssQxpo6HFNjX
atu74npklrfptSI2F6+xs2m4a3/YqOyhhAcbAYwuu1VTk377vK8Abz9iqtskgqQ8qQ6MbY6zK3Kc
cNcLhnZWDX7gO5J0m0zN0whry558X/kqTXJ8xsUjikhhp7OWcqkLJRIcFwbaXHTaz2ARCHzMwpqk
ygtVDfQUXimWe1P77//BLawQS/oWOVY2feFTxZ0sZH6YeA5IiLY1N4FyHx/OloE0eIEFD8xwwVif
JkL+8tjAlmnKMYNWRPf8qKxDdqgIy53nphTxsN1NYkprbWl6f0MwcQ8NuzbPWwzEN3jT7qYgiDL4
1HbhH/M6vWRBsmHFFXF0eWW1bgzGy3g0BAu85CDt8Ntb1aeRtHsEOUviuRo54VXIS6DS9FxyilNt
FzLKMnB/279yIKT3XngeLjkaVOpmE9vmKwSGTY8UcEs3Qr6GggYA4SRU5SYu4rCR8ngVKVPWvbHG
j647LfGc7Am0D0rTHFrQkmhCJ1Kaxr85WSSFBeHk+0QULCaMOaYUbVmnXh/7ZGbLWqJdqdJW7myw
/zjhyt1ABovgvd3JYVLCYTq7q7BGVSMuzFqTqp7Jzb1FWWWlgDtUyiKzC06Elzz1RPlJC0h1bVU+
rBFSuv4wLFyQrW4aqxX+F80vx+PiaH2HIkP5aD4bWXLlcgoThf4IF6ihGigmz3jiH4OYmeKs+OWA
0B5pxybgyczBi2aNkQdsh1mqpvA/aTOzfEXh1c/oWs1pxC1laXQEWTK2lOXsiopQcwPg1AmEDmkb
fveJddgBkqtezWiySg8W62TLqDOXG5uusXtvncXGxlCoBApsvPCKuUmaOAFUGyWyDSqW2JXCv+hi
ZDmCUIiak9eMV+w80SrmfUp3cPo1H43C9c/qEzDizQZ2bSJot+sF+hwKs73mdIcm2eqB+MELRnSp
BRxKoMeMg8wlU3ncgxOU8TMrF/c5EzGrMEiS6l+sR/NzeBs01NnV+ju8GJwj4KuVeqo4hZXw2cPN
8U5ptCqECvkvQBgF3NF+l3QD56GMy1QauUPOrPpHAAv2ONBzcz3sN851uro4DexuFvc+RG5pgQxd
0Dm9FfEPvRq2w6DfOE5IWP4qedDavkJBahDvtuMA/88Be0k4qcK3ijQTc993wjrUHLDNOZhp2wTC
uVawWFP9EE0EMN7LJSOnFqj01r2afzXNf37AD81lLVURbx8UECyMid2O2y1uAzKMVhRWxRDzoBFA
imSY2jxilmk8DJIOvt1yWZUq8fAd+D49bLatq0qXuJmi0SkQL5ca0K7jS0QeIpRy1fghDXeLTFOR
Y+C0wthqtXuJqpH/CNym99uSwfgX8jHnXiSdi0LWEPrrw4EWcDgPRNJ+fYhPMIfZNu0nDha5KRpj
ZaffZiUTeDinuA5ToemDlJXh/CXyrd8MF8Ybl8y6pVVx+ehYA2ocBDOdDQXKW1Lc65y2l04ZKgCQ
hB+7Vg7+63sFFxnFpirgUr5GuzFqFcGIs7q7GhzA/XkyAM+WP3pSVchiIIBSbegXRu7naS80MfzF
BRND4v1O+CmXHBlZLJjUzNlq8POWegKw1CPQCWQtTfGwppEV17hz07peDFw8+r5SseUAWisBxCQ7
UzhUflzpFUIN0RIMzWL0xTwys2fUz5VRaaLd88kv5O2EuUMlkZ2CuPdztz9788p2f33dvsCDVWD0
w21a94/qjFxn+zD5cMtka+bm5mRo8PaCEcwG3JnZ82mg3aFF73wGS9PNwxOeing5P1UX89r/FyxI
1ZcNuHTer3LzIoGIpaFLE5LQSuVKbGOVdnaSP1jBB0OlLOt/s3vZz4UCjJJdEK6xUhOuOsMDLr8D
Ji7ZcS7uhjR4xlFSWA6pJ+WUlpC1oQPM4RHC/RROnvdd9eW9fjGWwZ7nB3TooZcQVp9vOmkAsnZV
TekS7lsb4V2hLYNJ7tHArSi6vKjssL+hq7J3xuTQsrkrwVyZvvCuWgAImE0qTVq2tay9JTCmyKWW
TOWH8d7xw8TBJpDvhBHMxnoXvngEfBg9XjmIy79NqdEjrW4fr7UvBXG8xs+PkfS589eQMO7XKgUt
tUSu0GKTWc0tausUJ/BRkYl/3m1njYhf8PWYKlfvRc9vnrrrXWfYVgxjmjVP4eF6Pu6/8c9rHFHw
spXDH0dOj2aqwRVroJl+fZyuG9bB4ewZgd8bGhru9AuX14gqWozIn+nF7ipT4g8oxp1SHSRuwdG8
orpd20YWDFpUeSiZCTEdWoEPsBSx2OozpkujqrT6OUhheloDAERHagu2SrY23/0QdUYfhFkrAN6H
66XfSUoATYbCcR2tO7MIPNOznicGwu29tteamDAum5S19MzwQGE8cDahSUYyDrZ2nlK9E5kLnxwJ
+dXIV2QZBca5oQMFsNmi4D2gBgfFkAcVHwxuQA/KuFBbEgF9Teaj5lcJlP7Q4p0TKMNUR/zOllpN
3wkd1NeFnAB7lzNoxi4hF8PH+LEsDM3a3kHgqoW2WBn37NuLuLFcvcTiUq0EKgEavWBSatykypid
nE9GYswYTmcy5ru5roldF/7QHGBd2XdCp4sCcWavTlyu1D08uqy7EBu/90+lv+vzvAOchZ500Dxr
i5oR3SaQod94YZ1leqTsK9FX+URE3tSYN9faNZQLPB0vQxN2hHkCVZ/BhreGLAh3fdV0If8t5G4U
h4zBtEw6P+BIXjnWQPmpmnOTKn/Bxj8RChD/CUzRGXFtcX2ynbcW6YLM5jU+tFGr0xjWjbEpxysq
YqSlVxuM78d/c98niwtVYEon6Toots3L2VN53jR9pMZ57Fij4Q0ZFFRwYNzPE41ki5XI56ngJGIr
RvPxAUYmVZvaug9fah0GzRjrQeD2Bvu/0ITUKJ/vgKP60ZQYMXz3uX/sy/FJs+i63VV9QjmZKEG8
tNHdyHEaEtgqiTHZaDEAPyof2Fpz2/h7hr18LogcGMBPwXecJHJu7ZtQjMJuKXw/Tho6ldNT+KAn
YY/ur67bnOv6QshvqA6hLpyTuDq2LD4zsDZzYFWmfgU0FZmhp+XgEmtVVNk9rec20zd1hwpPKIVA
hV6kY0PxNMJ9sCeO2bKi5ePLPTTgVV/QXHxF22JuqvVClKt7dx0Orj3rZOswNeX39cL4zWIYWmE0
jS7QBM9qOGMYPiONIap1gIC3H+srOB5RyK0ETsLdA4ngvcLKZjkfnDZ+l6qIBXamjdAp36EoiCgm
TKqtqEctVf4ttzbnY+YqycudaHB+4WrNv8kB1ACMe3uX7Bxo4EsgBBs+ekJfKsbZoJGj0bDK4kJJ
ERZmtd6K/xjB3u42Wr3AL1hsnKpGhuhr3c0P1nJ2flxXs6HhLfEl00tRdHuQjT+v3slyJnTaKBqh
rPevvtZDE2rN8mTiDRGmQ5OJVHf+0wXPjqdUHcZNhBc0SkqDNWGRoPIIPSqIGCpLi0qdTA8twA9c
LA50tP3ewb0n1v7IstXYOkyoPd9+3u80spqXcNagc2wvq9lhITeTO3WIpEKpEihPb9AGuO3/BHrA
e/DIK03ubEM+QfQV2zZqzCInUuL42cFsGlRCOg78r4Bx6Zs4HfjNO99fXL56ExRoIJEE9mZUmiZo
sI4zdfHpg5e6BHaQ1I0Htzhse8J7kzi2sAxIdXlJrowD9xFJ9N2hshuddPDwLi3VNZF+gDwC+ia+
K0I8DGwKqXph37iGNj0uB5+4i3zyvzrcV0ppW9qY6h8XzdUn0egwTmKFjoEdKpf3IoHdifctF+La
w2Og2K9hpOqjZ5A14HXtJLw1pWBu4SwRBqDOWSxZ40RleZhl9z/FGgkTVxJXNOP1DbDzz6VRrNle
Nq+l/IAMFb+46NwwjOa+cb/xTxOG4cuyTdtVz09V0E1Hf80gBYFFsacGy4mLVgDtinXU3CS9P9mJ
I5A/mOABZ+9Kiqq014JZCST2AyEZSqW4rXTI818TZ2R1EzcdMRRMgFj7FpY4GPsHWQnF5Pz7SJxR
SQwTCYwVrYrJQfuXl+zEwXB66BYAhhaIG5Rtshz6glO7u9PTxXdslv0KJJvb7zcecrv7sTZyyknD
TzMvzOproixkHKcoFJRA3tSOeMsqa0AeCgeJQYx3z6BOrZW22KOVrI8xbGVIijmdxCjfnC8dEOng
Sh9DQCOSMjme4mDVaBsb67g/ytcuuXyJQVIlklPfaVChNvLDxUdXMi/F0Ijy78kL0JkkUXzhyyS0
xhBQ/Q95c04wwu5XYFSYLyeWTtWNRfzZPqsmaNcr4TNa+O2G5VJlPIgEoA4yvPvAxuU2VTfbIFgr
SOgpjw+N1G++r0vXowLqsZ8mkKf8m4Dj1NTkjtSV0nrjrtCiW/zVn9TpZRyXSQ2FNJcE1wZffp3I
2VqUi+MiPSt8pYgYbTnzdhSOEkvwZMDwfDpOCXgleACyD8GsDhxQ8pgB//dRmx2uREd3+it9/XW/
8Zz1zCsnb5A0Typnby34YPKQ7TudpNy6HrF0ulEw2bhxn4HnVYdJ6Q7FrguE6mzn0tcEDdiaovXh
2Mya2TKK23irZUkVeTSkAlbNCcwSDub1hw04Zxrk3C4wicZJDZcFqgIgPZKtQniICkiR8Hu6xUNJ
14aGw8LaRFlOtq7ajUX7pSBce30ua5mrOAb6++4Dk+QSlsBM7UYKXH/p48sdH9s5aQOGB4W7U9Ld
NR77eeaYQ6dLc8N7P6wSqzhoAk/KsmpnJvsyIxyqucaHca2iuq/SN1tAhZvDoc9XrXy0yqZhwgMb
9MMsUNm1zt6UUgHPPQebDZc2WyXoSmNhPVTW5E+EGpW3CtTDgVfh5NIsFFBSMiKmley1xqkAIsUv
msr3Ysd9lz9gNAlZXfCGc0Dp5cDlzWLVeHrSEXY8fQmEfrT0c6uAmMM7/pqNp8ipUBvdTYpooqn2
E1Hb1sSkfEcbTqcHbwP2wkP3kqw3lHkP46vvneFiwZ/c3zjvj0dF3H4bNDBx80necx4hkxES4x1/
nVuVUuhZnzO0rVKj435Qg3ccYPVL1elCzV9vnhb+mUhlLAi0wtAE1iIm/+OHvKauDQ8ovXS2u54w
F7VqBI3e+qRZ+BQVWBFsRd+qw+sPIH9pm4D/FPqHQ/4kSC4WICGI+ki9SAEoF6Qtn+G4nLLVxAii
FM6l4Zkg2AmOmgK+dGR17nmy2Q6OLgl+71ShnM+n3wX1eVQfLP/BLotyM4Lwbj6lGI22GSTx/g/I
HoO1gcervIpYVuYN0F+VMLen/t9zf6mFV9vAUUZiU8dJFv8vEDBlkEFCJUNbNFuIM7myqkF4I5Qw
Q6L8QrZzYw0ajqSsGbS+oQ4uV2MAZ+rCHDTTIW55/Wv+QMJvNlfjYN1dAVEbBt1XmNJs7y3v3AE/
soQaZrhD7hArMa6P+0g6kvKd12ViXvDBQx2Vczu7xmzaeigk3AexsDchxdql5N3gkOHcv+9Y6HKJ
234sRpErC1JO4SaRX1BsSoTs9d0qvtuFDYqBtXrWogki/wJtgHreOFBMWLC4/9dTIaOBKSBmJTp/
SXFRsDGitOYrpG4cBZ22U8A3iptucNubMlxgDykhmg6acXjNe3FnCARFO48z72b5ajYpXJtqPAnF
AvfDG2bOLgl6OJG3I00cOi2sY5WHVmhTMTYZe9Ds97smdIFqGuhf7zQgXJfgBzqe0orJJxwdPy6E
0g8e735s2IJvRJVYpOt6X3FGTUits5YuCS+L6Y7rvhEl5FxUXSG8bRD9Y+8SPU3zF4ioaQvD2Yo+
z+g70q6MDvsiVfWhvoVLYuMIE+T8OsFdX5RB8fl2hBS0Jl3krN5C26UHgT888qow12lbqhfZiGyD
nQqSPid9YCNIq4iBRzFVk7gs8KMUES1w5FeiumMAx2iq9Ni3le8QYZ4/iaVvp9CIfTJdm2r3JJ/i
oqIK/SDo+KUk5f5Xqv8LopqllOvGfE/ooCu1DUA2EO774c7Cr3KqzxwD5+lb1E0BETBAD+yKVT48
mhH5QOf4XEvIlkH95fZ0Ps2l2YUXellXRLTrziz4HM8jXYs78Wsi+GXFJCLFM+l/q2gPAXfVeTCG
SAxogu86Z6RSrHEUD/SNUzmoee8gQjhtH5gR2mwkpo7Y6fl4dsk6s9/T2kbykFSzbI/pZdQa7neF
yv+lJGWKB7q4DOxNLe4TEcB2mgPPZ1zm4KEzVk/zCOHzRHvg/0AWorAwEkJZ+ooz89pKCxgD9uTe
KKG3ehcFEWMw5O74SLcaujYdMd4ujtLX7mF9ntzr4HWoHbHn/1oeVCf8bHihA+AAH7K+bn7UNVS4
tYmm93caXa81YOSt8AUF6DuLIOBAosBPaTQnz4MHW9uhlMVi6tImCSixFJ/wBM+2RG1qRr44WFbs
+aiLZ9aZ72WV7+EIRZlEVf6M5g6b1KMXxA3zsfzqH5W6aAHdOabdQvDx1lhNrr23rKAEF2rPq9jk
KsORUW1L6vM5yCKqUhRq0/RkIVP50UtlBBAPWLoyur4DrH5xYgO9yt1YnYd+vbz23f7LoOJxNCJ2
g81RLzm9jc5mAg+h0himy/pzK5wTqM85Shln1lUobI9nMECezvrtj1k4Ib0Cs5jGf0fgEeOAry+1
ez75JO1+aJsu2MzCUdGiLtPwwPwvkZ9tUwJSFXEMphHV91ZdvElLtoQkwfzScuCd4sRuCdikCgrB
4VIFOZipWNEbgeFS9PQXa05BjsL2LrmPRckoFO3CAMazO6LwD7erZshxvgC05fNsK8NSaFOfGiKc
svZhUYE/iq5MlOrRRD4npvEEZLF8WDc3YsWtd3WACY29OGH6erRrUu5B6OX/hSI2DBuHALo6QEGw
AkRAbujqz+WwsWBwdq8En6EJvRBe+4WuIPepO9nB+TDgUxebrWnfHebm7yFbuKuAzb+9hUMIfwfY
BPxeLIGtU64cpmBxjSc4E4yRgQbKdfaF/XJ2d2HbqE2L1hSPmyd9Psk7a5YMAUdP3SRwu6ZMXS48
3VaKvG0MJbu+Mmdo5I1JRuScpwdZxzxBlFm+AppUyHDc0EoOM4aKw6hQwu/glOGbXQrNiDMSqPoy
iCEP9mesMTAi6UKYD4F9Zsl/AOstTeHzddKHLGPMtGvm5AIZ2da4k+ZZnnyyl0YjVjgHPBUOymHm
qwFUAuaeuNxaIVhNxEDI+1SMtxQsCOCfp+xABFrEgT5jNPy1xzlHcKo4IGifxgb+zG4Bp2+4v/B0
c9Jdj4fIuFZvV7h0XYgWtIjMhpqv3/pT/0ICPUwSU6IlA0W970W5tBj7Awp/SHrWXSF9qXqZgm1B
Z2WKPtliFo+7lKewe8Al4amf+GhSd/0Cg7RECk7XghuOZJ6wf01dKvLSCd7ClIKYtuF83G6JhI0I
qfYEaYxRTLPH8eClea9EPAaenDjbOaoSjI1NoPrIyGXA+ZCz6fCi/EMyxnYejApImMHkfDTsSVyG
Niv9Ul2uy4t8+/or42vvK/ZUc2h+6XfLusSgXckw5x8G4bXQUJSvTWTJ4c3UTgfDTsYELogt76GC
aCFWN1CdOWBW4grflVTfoj8CJu9w7Xn9fv1emwOW+oXGFhCroy/Cl92YBzZdKSfi96NaD3oIJacU
AH4WStCnpVbOuTqHoXjV/ofsUsh9Tqitp7YRJAZLji14kDCfeR/BWKuulZHhfaQ8kyIq30VWKJNA
+DW99fHTJWD+Dai9Rlgo12CPFOzUxel3XV/7GVNZNiAKep9h4+voi2ISpUWz0I+2UEESyLpmISvY
+i7YHSo30/lpqbcTMy6Ngj6jqHxwn+Xhh6f95Q9uHiwGBfXOVxEmEhzaKpldMjxLOScfzYVFESCi
5jSv7w+ZDIRFZcmw9lg1Zij1UPK7n0ta8HyKBbR6He9Vl1O6fYXGE/0Odn1jE/9AMVycMsM9WLOR
uyTYC1iBh0ArCPYfUrRH7ag7svidGs0wB91ohNhDWx1wczMrwfH7Wob1Ew6D2o5zWRGDgf/gtUfw
jksMfmYfiGB9QCwPW/jVwxBqi73utWrQkFMtt1pZnsr3SOoUPyFy+RNJOrwZZ4Uq5OAOLKScmrDf
3B8BfI0uvoYJgawRi5rNC2sLUeyxsSGmN0kk4//AqX4Bnbz2C8EKZV+AKzryjR1XtTi493MDEDtU
QTCsFXbNhPX2iSG43NheYreQ8KYYSIfYnN+CnhMxJO+ayqln8l9MLBiWIoJYSoydGrc4ftNRh+TF
gJzBZ7Eep3NRS9Klc6RL+lmfrwwQ6jXrvNzUQV13wPDRrCplsIv7oV5lF5fshIH1NX8N6lPkichw
5OpslHm8+sfhKtrzEhqZOgvnHXjHa6gR98oe7ABbwuoLW5bJvvY7we1inh6MIAA89F75baa0BQDr
697kpt1F7wU4hgOAV1YNUjl+vIAfWm/EaMKneeZGOsex2FAqrPA63Gx3ikz3+jbUKvqxYg16ZBZU
cV2wMALJ506atGeJFet4Rn94e46KlCMCxdQfn3HbM29c26bIZ6xaUd/dE4Uhwj59jpRB6Az1DD/5
jxj/4C0Y9mMLzjjjqNO5OGPUzGUFSGp6a1r4emjZvMdZY9Ns0JmFVVEQIvskmEyoH5I9kS5szdIl
ZFT/7SMOMjx8xFxcoX5dKXmzNJ3RIBfTW5w0ylF8bOlDsLadkhC6gUyx6hwRskp/bZaWcIwfp2Ui
vMrcv7v0UdkDrgOfBDPVY2FF+J6uaKH2hrJsdUqU/5wtoxY48ybgMjm3n3gpAqBUXnkRW/HmVah6
FJGdWOiz35/omot+hjdttPePTmeYWjKWeYfEyOP4xkf10B9b6czfGPSZxeD0yAe3L/VJ+53UN6bW
KHVMrkz2xZbH+WnHpsm8YpABRWWIPUf9HH7JyebIvGu1Wqjuyn56E6IGRBwp0dg54p1t/mRBf7Bc
Ojw25Uo91KpCaM0MnVyMLUOVHn9TMishG2psRcKfZTNCMu23KrbzzozEhrrLXElRmq3MEJBiJttV
B3OfNt2qM93kUBd/eAfTi1eRyLIEKbFZa8XKcug4ZoRQyDjoNMnr8z35jc8rQys2UWp/zVqsjwgG
gavAFcQcYdw9sv0rgy3ll+YQIym2aEBDx8Thc5Cf0VFURLBeFwP1UjoktNW98NLP/UxE7pY3JqKg
q63MObTEH4EvHFUiWcpeMvSsNfOqEaW0DdP+MmxLXgXfTzAXZALPNNIH1II8eJwshC1xh94nTqZ5
mtz4N6uphvddUgt1ebsDexpoeIS6wLgNr/B7rVoO98EvnK7Mdxd9R5vdfGayVglK1YzXqwFHCmOO
yMSMRgXbtHy/TLqt/C2yOZRIXqAHFVAcXi26FoSavA9cfFfS7gpy4bnA7FZ1EbwopXkRFGPdsAVr
biQunYUj4uQfwfUMTTLbbGmW1C+TL25Z9Zt3jIpng1wfEbYVNJOkiK9TtPtJE26psMuPTb0CiWGo
NXidiqhirsglqTthDzUDGnV2kst/4JxjBItOCwfhs75s8HaKnHdYLnfWU8zFXZ6wOR90vYepGcdf
wIJMu07rgScz0X4Z9jwkNzkIUhYYxuKj+HogK1QxZ9op6kzJD6wtaAQ18UfkyAFkKSHRFGgJrlD3
eJBpleh+Wc46p0V5TePp2CN4Kqzt2f4gajzUSiKC/35Ocg5FdGslMo+LR2L78c4DsyC7HZucQTrK
HvivgP1/RSHTCJbTgpreSXZ0kloxj18cSKe+UnDtS3/Lx7oZXqurQUvdzfV1yfe/LwniAUqkNEtG
WmLXWt5LnMNUTCgIZg17qrkdQtG2Za99FqpE54hLeSLsdLVPKFXJDlPgsRS6xmBD/1V84wV2HxZa
iK2RVdsS2ig9HT3EZniDNhFhFVtL0v73RKEgM40fLVTWM1whYh6YpLF6PsLoSaalFJ9M33GmeR0y
1QAVJCqcpCcJXnCTgceub7/VyCnEcc/LjXwExYvp8Q5kOC5nSA5gBh2Q8JTVQvLjQ1gJhFn3Wuhq
Y24uDaXwovxi996lr9HnInJZDwdMqHfB5dZgCXzrcpAe1lO3gQBYUlXVKb0kFGsoE4H26V33Os/U
jjN4j2xa3CTI0g1YoUNzOqzy9m81bIulmd6GkPC8z/COkP6pXY4FHz/lYqgxfflJmmRY35tJMDxZ
yArtUwyOQZMHtdJd1ji2kvedfZsoSiOWW1j93+MCExYe6BOm6xabKwE4Xq8RCw0cJn0avxArxk5W
pazN4BohasmgDyS+1Zx2RNaCqCjb9DSVEgj6dm3wSgx9d5K6uQ1/jUWC/Cd3SaD5ktiuvSIdtMzg
G5KgKhEwSc2QqbL0rNmqgK9M5WosmD8fIecfJSlsQVCWZxTXp/vfsDCyKJpAEneJSCGER3OSEgFN
xlogYS7bmqYhLf2xVZGGQwf9Rm2z1TMknKXhbLENqJ3QCb+LxhHPmafZ3R48LqBKq+hhOmnHe0Jj
3dUj4YmFGhGc4QTy+p066Hz9/RbxoBo2HbPexEhiEoDhzydUnRY7UfTHpLkVEM18pxCcruPMqvcl
aRErrixmPGbwuuabTl+d5ulyumpCZ8L/wKHQBPx0oYhIqsOcSYqjFaCrAl2X/s+gdtV06qv6xPtn
u1j6WX0kOzso7DqsHizT9027/PAXYEpHFXp44Hfv6KgtiZInFfhYc2ZTcc0iWhz7BQWs81dK8DCC
UHhXwG028szpGsRbBB6TTvmwvqsgYCFdiuBnj9MWnexo23HH51bGqx30SR+TVyXhPcM3hfD7kBYu
aQuKzfmG9lbBE0aWcw3+DzYkItZwgoNSew2DWQnU0TWOeDXp4EBUTZ7U1/9gKzdIA2dJD63b8ATj
hv9ITB5rt5rWfUnoeB2CMBz2qGUCSfOEoa4j3iJOype12oScG5OtOwmoo4SozvLeZYwmvKXGVmeN
YT9wfemUfUoCOoDOvfw4HFxLQcOuR0X3x+3ER4ZEYcJjf0VmEvMIKyPjsYdeLO6oXsGYLyKJdNWt
RCO/AptVTuBx5dtzkbEnKWfx8icnb+C191NIoQXYXBzmiTPw1818b1eyiGh2YDRLiyM05CsxRWhs
aG0dd+etg1sl1UZwP22KDtmVdxfuex7m+9pdGTVdSqgTDuFtuxSDg0auHjGxGuO1FuF2TxGtPQ0X
1t5O612LVqTEcuvsXt6wwWCX+X/NJHvxaaxhLpQEAgP1YOal1KtNR2Bt7C0y9FU99G1R3QwSLt84
WcPqbilquvGgN++fgU7J3DTXffzN0JrMnetztW2uJ+/fef2Z8ODX8QtH4i1KFQi8SK03WTwf7zs5
1ie0tp9Y/kcFCIgYWh/MEobfj4YBG2qBBPSjolwcvhilsxHaR4uWc4a8O8ItNkfIe2NeLBCBHoc3
38uiUd1uC9PmQjOXLWTDF4TGMaM7VJofIo6Rg0x4XRFM0b2D2Q96H2BFO6NBa2nGcgDJSQLDddnm
yl2sTjbBNuBXCuQZwf6ODo6ziC/aao5C67GA30tmTQQq/oIBr2ZrKVZjdl6xrfgYdbF0r3+MCq3X
2IXvxekD37wqhc4DjWiyQozLLskwheqB78omdEoWjGtYTmwbpnvleky6+CpxyXTlrDJqHZUHsj0H
8YHeW087j2PUtm1I5LMqjRpiD0gdTZ0FoZSQCXzio1AKsB6v1lCUoB8zcTzSX9OhKJ/xZ9reKd4f
QnYT8yGiG1a0MtGj4SFh3r0vUyLwhm0HxHB/Fkck+zdzsqrEWdqKbQ2DQs4Brsy693ID82LkN0w5
OIx5ZGmBIpdXux1ALHWmflTk2FIaXmWg5qS92VBKhRByV/+N7gBz/2sZGjA10RgHDgK3ohGKHVCB
R0QAbgiDGp7FHXit0kLkDU3L/qd027vq/9h0632MfAvQop6u2Q3vLAjswliGprRBZbsL/AjXwWrS
tkr5CDFgrdqt54rnHhxPN2sPveOPXhUan1L+QM4A7+W7lnSa75V0WKc9rowIUhubujZB8pScRBEy
b0YUdfCBqQ6z+uWXNwJWm7WLe3vskQMOOKsfwnCYIRlsv4omeUbjvJZU76BkzGK5TbX2MCrSj/gq
YDeDo0TfZbYJitNUyjRYADc8czsxMitgZLDicyjO26+jLRLLe5XwZ/NCq/CBF7r09E7Zgq5rHgeV
qBBGOfSvXHi5QnvEhl51C9dBlVT/VXhG+jKEgGQj+Hr18zXS+wSmjrRPO8FwCQwBPHapbe05mgVM
OxDy0sOrDEiVjlIlcKn0e+iagIV0jmjYMEJdHG97axoT10Jh9SkiYjL4NxwSsG4qG3DjutVqC3Mr
rz1lst9otdqTsOImpsz6by2pSoREnQd+buGH6B1WxQdL48T0E1hdBMIEDbwDf12wiv4qirL5pSVi
ZCXvgjS3LOtLTHpzR8AZGNwn2BbdNaJ+uljhJCwZpdhqMfLnC+n/PiWsrU9FxSIhOyohzO7ZQq04
bINYRNZ4+rjSJ1wYtL9xpa7H8EzAUKWD5bUhzsGdAcUo1g+yPQnGDdNPNca2Yty4ZcFbdou23OC6
TRdFAqC0GPoJCW8FXSCJQD0T4qTChqODKVIliSaJjcOzzbJNEBCJy27TONpOJ4jFHRjFKgeI+teD
5L/fsoPANdbCaLtmuLxhe8PRhyxTgixH62LHn489wy7GtbW7rvuskLjn54pxM9WVLdAIqeKMZgLY
73DUN9RyrvBct0hPyV19uolCyCsMa+uFnOtmZuOlGLJkGnAf3rOjU8wb/GYvtoXKz6ii0oMFIQA9
o0AVobpA14PpQS89fUPiMRvKY+0dEfKz9Dg7OESRxswDTAMv+wkf6gvgg31HiMetTbmwPjHTsUHN
TmGs2XZby6gbhyh2riRTr40lYo4AXXIfkL3phiFA9/wj4ByfVcnBPyNI9lKDASCpGbEJJQpgSefa
01DdVoC3SuuzYuYq78/kRqXkxXPqm8fPbrOJYgbmkA0eEvrvSclp0h8gNyv41gFhDblxWQEKBjnK
hY32kgN0Eqgo3ke6TCYLIS6l4yBX2G8wcWRWkjV/rguwmz8jNPR/zCHrEzO1JS6Ng8mKkQ/6v1ub
rB0RVZb7O7yP94N0iBgRJfkM7UerfCsh2cOb+E0iY4Em8TUdY3E2vzVuJ85T0I5Zc0VxDPyI8YAR
Dw5aSYdhDzclxF+klnK0Obyi76l/A/yqw+2N3hCzZ2DJvqx97XLoLWDR39bm56k2Qx8EZnOOezfN
UeXL5O2Xq3SjmOiOsZvL4W+q261w6651mAb6K28uGVZH6ZF9Mo23tDRJFCBegAqLczExTwaCFLQh
eUtjq/bj2AncXlqlRT/KsUh6e50fLzlpdzRJ+MxaoJV02k0v8F6oa/Uda0hQiGN6G0r7F14TQKdh
lOwwgUxLSLNSeuPz8hkABoPSfzM7id+j8a64l5GE9rAYkSXdxc71P2uG8DbS1T4bj+3kfmU2TqQ8
pHxOnXpbQBAFFrLpnT49BF7LBQZYMEeV9RkjBKIgBCp/A9LMHP+nw/v6kQgyduXzgLwkUdR6tfMD
zszfW9YAlqjMV1rBB4lkcZhLi8/a5Oku159EnvZIf4kAJ0a0yiXr/wweSD5uVZlH4PwNaJlguFWo
e8V/wYgCsAIKQdz/MxbiSjhC78fxss+NmZ8i//Sdm61hFplfAtm+I41sFR3JxGMLP+ssPEVj0RNc
fJnkAx2C7ZJXVSKqRTjsLTqdszOFkyyJdHcoL6peZg4jPAzsrQuga7A0DdEl+csT/+jIDoiqPK4E
r3AymNK7WIzu3MU/dQAhqlXSpNWB+2ac4fWr7AvnJ7GSE73xUCTnzgcDgLc2hLUAi2xIjWXpbDBf
To7QB83tT+YQ9xwj3pVI17chiAhh3OFjVau9dwbd+WZbiRmTMhN7iNOccFctmcMcrOS8VhN9EgI0
6O3jOb8kN9gHfKjdruyCg572rkn7i4/YMOcowAdbPmGQpazWbRmRMQdGCADc4SD5UbWW/6GlJPTV
k6uFLARehZTPaDDWn4d5witwTQQuwfpK+m0cA6UIyR/DutvEmlEGFzur5bvLUnY8FVWn1TKh8jRF
H26oMnJ9LHSTYuMJ0I6t35MoWu+w9XekV8W7nElJLCecOCEYsW+PydmqpLN6tAsuaNpeSADWRGDI
DiPaqiE+3IwhLgEhYipwmTHDbchAVAkT+5gpe6JyqAhSlhzgcqiXwAYlpn/Av+r+ENfEOJaG2Vg5
iGuSlY7vLWs6E9c5QB76O8ss4ybdY94UegAEmldW4gd5WyElsHvBPCEEUye7PHHjS1tRIC+qaIq/
uA3n3xzcapNVI7dz8Hk9ki8LOcPNv02caJwBNM3RAKOZf4ClkbXK2BgAlsfaXfs5mvyPesK6eC6t
DOwQe1DjPSeNdmnMGIKDLKz9QLydD0InmH6rJ9d7WGrqPUlfU363MGS3B62VaCwdz9eYZey3yKW/
KdTItm86pUNYMGlEJ6NfVgeviE1CRvSwRj4bfGDBq26fl5ghTE1dFU4tPIGlFkU/W19ZgULYDuXu
5RXzfaB0sLjLR+aGXAL07l/TgTcU0nGtmcemHIeL2LSKya3sjY6dNadpkjJ+z3oVSrAWMeGlUh5Z
AYbezb1Y8zz2pvCzY9w/QuPIBQbJbiVIg478JJLrxNhfqnjrWOFPUAoHaaBknu7RA2pBZfe4JEqf
tSdUCNzmyq06FTho02GNnbzKKjWt0NsFsR8zei3LcXnU+rLRPqnTg6NEZluFCqsORsbZKE8sRqOF
7+k5fPhBdKBMaEvRHhoa9+ERvBpjDc5c/h5md5Qo4ETO/se2+Y0DC8zTdGWhS8DYiTgghJq0dG1/
L27aPNO7/7Lpy5YumN1y79H+Ev1YIJOf0WH23UAZsbD6HCJF8zUwoWjpw1K0xtchGBE0SZziCpHV
13WIfhSy1mVQQ7RIggIdo1Ju9dU4SC8/npSsqcYYCIjtUvEiHCbS/yx8jNtHW9k7opGyUFB3iy6x
p7BHYYYZuVKQzqgBR+1RW/Jhkc13+9Q4cwFyx5Fw+Me9+sJoVvfPTM1fK2Y8k6ZUPJLRq4p8zGIy
xH4hLNBvB73BMKvsN4aSixeW5QXu7KI+03mdajWcfJJ6aMGJqA+Z0ZIXZf57OE4+6Wj6sFyuVyPY
2oR3ax4GNTvl6UyLG0akp5/AkncA2IDjDK0zgUZ6C+4oIqoKnOuQYI+gi1w9UFmZrk6cMC4gn/DI
fa6CbOjCs8vsBhl238cekJaY+5489XUmJZ77ORdur3wTrBKwpBVbZ5y4s/7cDVCfXhW/uCDRH5ja
QkY0IIfmwg6VTZPTQ2Po5S3r9HntpweoBKmtsf4bVhMbrLdYKNV4AzIzoOpDihb2EkQrkX7ONOQc
DshQ5KP3eKzbrVSU8H4vWrZ4rP/XZxRMkQfd5Argzip+OytgiZv8unMDe8C/89zXABeSYbquXEwc
uN8SnElEE3ccfXjG0WuGq8Pb4cwf7ghuiLN6bAIGukMMMCzKJS+Pyi4ppsqkRSfzIJ6ghBTdLMtl
m9BvAZ2TV0XZ/1pmN2yMDPwMw9NFhotHznnaStPKJ+f1/P/yXeExSDqru4yWX+PsUTgIKvThjVjT
FfAOLWVzvnumR+/pZsgngx6ZcVRi1ldeqWzIoq8FwTcqLiqCpW6KxgaGCcryhjEG+Oz1AuH5yhj2
INy822tgIKovU2t2inuQcxLIHtdlFlFs1OFUM6bYtBAKMfhGz3knZFiDPNnGmwjct9nZ7j84zEcG
xA0/zl5TevukRj2IDcCy9PMsuBlIufi1MEaLO1MPcRvLLjtffV9yf/w8t9IVmh9Ck3QFPrrcRmgO
/bqinpaBbsPACEdbdKA/M0SohYpjcAeJSTYb/vIHe3Mw2DcUW6MPgMYgo2UG2NUn6ODv/7keYGdT
4W8DRSU7HpqRioMmNoXCnrFSTPpwoKBw/t7Ee1sN6Xd5E17gbtNXHoUyFmL0JmQNmFMhvb5vhlwH
4TFjv0GMw1Twj1avglOEXRd3VKa2VC50DGkm6w/DrT2FfraG5VjxGwJ8Iiqy1ym1Pr17c8SSQE3X
EsCdpKvPtxig7O1OK1MXrNHAqmHFmvUYfikCzTsuvPUH4iSFx43ydT2SLbXTrJ8agSukBRCNYvFF
dU6vyfD3TlSEV2pt1dtBnGWiXLP7Keb60Owo5UGLhEdk2uEBoPw7OOkbiAZFIejjv3Oe0OijTtTF
wecoGSsXM/Jryl3eFb8DT4iLTgvxM1Jp4ibKlhLt7/dZlk9b1ksw24ZVvvH3Y9idVMX3+Aa2QM2J
3Om1J4Sj5P0F/Kc71AWjpyFzTx9GT7eFDWCGJ7sa/MBn+tjE3PqDAQ8UgR5q5UQ6FZ28zAAtfbQt
dUBgI/HYekGWJx8TY0r+9pY/S5YQvqlpJ6QLkcJ96yqo3WG+UBssYUjjf2U+bywB2yfwrN2yIzuV
lFe982x1qfjlWNjxQQnm4hNLUHH0vQQ25vLnOnWEdt1nxzTcbcoCD3hHa5YOdjwoNV1qUNH2ZdjM
HEEDlVfO3TPVyk7qi7dUXTboTOmlwmQ15Ot7/QJZ6FV2/BMgqE3BlB7TazBhSnnlN2Y5PNtSdMz4
zglq8D/lazdE5ixF5g5mE8RuFtOh/IvXuHCxLLLvaiO8gFvuQ8a3L24FlHX1KzpB9PIQlQeKj9Qd
DoUiFUkJ9aKcOSJmVtmZe8K/70Py4hyUuvhVqIRHANl0bjlBVg/0BOugjHscUjj0io29IRqSUebN
hp+wQQI/G1xFNhaMWufjng0SkGQk3CF60JWOGMHyG7YKwizTyNI6PSTd40YAdgR9n1nQBMIbWD2w
u0/nS9oJUKxVVohcWoUd1nk9FIsOPvyhLjKCXR4zhUTw0zURb7/zITtRMYv+tzDepK61Ilpr43mu
9CdEWyz/8D9xknLVV2ALMom/0FfLNYXydO9k7uim85vsgjjc/NWxHXrUPnx52I+4vrWdu7GK8aPt
UY4LiMTUIgJfhrqWWA2UshuJ8ujfQhGSMGdyq2iWn6Vb+bpoKu/MhucWYESzk75+5JlsZV4S55IC
meTjx6j8dI9q9dmi2kZVJhMwvEJeGUlD7vtJ1UAlMKotJFGJtVBg78ukQ6lXfI53iP0txm4Fi4u9
a47l1Num5/7Vvv5UK7Yv0ez6RZjS91zEuvhjBZlrFcvmTip4lbRRSZ7dtCWquWHKtsY5ghpmef+f
WMwvYG17SnrL+4A+H9GyqCfcQPxYknzAtnhHpbkeJhaDo7LDlbKGa4O96raE5W/pAnitUJ5eCZ72
pMa5GfdraBuTWH9aAFznMIcDsou74Z/Qe0ErmR4kDJk2skfKU0RrCTmPxw9g9xe5OV6o3n42LZrl
78LKZFEPmxXpak8SxxLHIKnXVZDWGAI2nXn/qobMIywuLWIos+DLQ9CAE+BGmskOFj8Be9u9l1aM
ek4R06KrcFpRIi85+cyTFOiLG3m1u4wI6w0NpF+vs5DXUe9aSi8pUshdRM5VARTkfIVO29SpN6f7
NU3KvNZ82CGaiCwMSF3RjskWEg0i5qEQtVSsz1yfXoBs/L0mVWVxv4zHgonz+miXNTWOaoraX/8p
C4s89P2JR3n7efmwg2joiRRhztg+1kfvh9dNvnkARHy4dpis+Cj3iN2O7Y+HXGf3SfmABkSgwVj8
DlcktBHZOb9tKaMNiaC8QL4NNc8TtdH6fncCIT/ng3AbwNYQHlOwnIvXf9akT5/F9oLxgIRVcqts
00sTTcAX0VF6xuR9g+anuza3yarNE0RKj9bLNFdTXdFhHHSad0ztHAY64LhH+zqBuOsKBzhkDGHv
hkgyFNiHTmsjl+r1W0VuCHEy4rXjjbnPhbrI/9ciKL0ZAPoU+cacGzwwMfDfRnlzVyyFYX3eNFs6
tAoBeNGymu/ZEQsebCfs+eKm1YJb5urWwCG9vZrP8fOgpcOcEB9ZIVcRvQa++eeZajGoH3bOz8an
5Wz3Fp/QwOXwAt7UipISBROaH9zPXXAQrLKL+9kHBcQc/RzgtCgO3KpOMGvi8G4qA/DNax4ytz++
qWpDgE5UPI0nhroUG42Fiqj9flt6UkXTUNsaDcjZXhofWroLNES2TKPzQahd947hfVPnr0/R5aqC
hjlZJ6JEl7GbzRT0FOR77gEYKIbykryx5ohiklPBrePVPvqwT5VteIGsfJoBJaxRvO4rpiRkWHCL
xNsifIm2S23FN6StGlGLUfhbRQr1eVjB+F871Wvyag8Y6OBoHv27NJoEwDnVqlMtUnaZOKvhekEe
vE9RBd8zbVz/6F0CRvqxfiyaQh+YHimbsd31TNc0QLUkk0GBRNP+6+IkcO9A2oYAPWCZQpqX59EQ
oHYsjEwN4B00CYnhwp+dcRrUzNAoBxgY+TLiVZ3fKK7QGSp0rY+HrV+BHn2fEVVx4ld0HkTYtg6r
7k+mlnw/JY1pRBtdMWQZ1WjdEIsxfcJUH2/rFGDE1IrP2ie5ngHCe1vIiM/uk+aT8tucXCOx1enb
KQF0IR6aw/Gz8hkYAyDc5TAmw4Zt2W5jjt5PWEKbilSD+hJhGt5YWR/Gjw8uIje7WvvDKHmme+8H
cqDELxKNGbZxoBpveB3fbmzaAVeBO8B6UKTs2OWbuMnnbdCw4Lvedclv/kl2HjklKnwSVpIu2g2y
E0bJtFU1JZoRsuWka+9+yMTacSxBlLzLYC4stsqickBe/D2io44ow1GkFt+X5Rbz6X3fmojZrYWL
OJUEQZ7Zatm6tXQKoNad1kN5UwdY72aAQqT5eADmNItNmBg1BGNRVzkKxBNespHee0jFsAe++L/g
nxB6zup0KNzC65mDkzFFmcWMrfy3HUmyKqjMTUTXA/gH0j8TS/dhjy8mUF63z89EEx4hEOpxYrUj
qXnYF18TGEqjXBbCOiYP7n62Rp58Acz/5iAxqhA9+Yi4oLqyoxLW+zzO2G3LU0Iy17Fnsn8KuDsh
SrzeNUGkn3HbubxiHK5dpsoDv8qCVVstCxzFNiRIhFQa9nQ5cX6ZPMEkvIj7Hi3a7lXG22nA/dOr
4Ux7I4NrX1eWYHSRTLhuzBOIpZ6RnvXQCDP0IzEF73GSn2baKBBg/JP1BcDdahE0qbwMccqBEUS1
YZE1KTl5bxfxQKKHlb6FFpwIfJ+YoejJb6hp+zxeI3jPkluTJc5yx4P4UWlglYPeuFmjNiw4aTFT
iGtcCdq9q16EAQWC7XAEYUv2d4+i95NhjzF8VUV8ND7C1teXpQ/LPZqvK+6Ra2R0w2qO0lufST12
6QkZttBEYj3NjggETiFdA93NDncu/c1aiwUSof3wpYCY3bTIbr9hOfPr3E73Wr8UQd1OMPDJ0ni3
seHVDV4Kw/dM5KbHpWqlA98X8yOnzubZCQXq3sG8JLU8h26jZRMg7MU+zBwx0pgJMgEfiYWFOutA
jIkdDzp1R3x2fGovRJ6L48PFmotnn2TO86nNq+20jHhXlb9KAFGjW5rFR/jWmzbv4hOtqQRQzGV/
odm+szWYdrmECI5IQGGUMy/21WPHHgg6zBH54ujHZdHqww+wApx398lgLX+/VT2EC20rC3RilV1k
jVcduVJ0srMaKHWjpz9uQs2bOGw7u0KtWuQ2iXTRCyZIgy4GUC84CwJOB8WhshmO02CcgepULHJz
E89ivfZz4ZnGAbvra8RjLXdD5rm61mExJuAKowlsQ1PXMiMhRXBK2OcyYtTQtLOJRyoh/Ic2n1en
r1/12TCMady5thp0OlByZm7pZkS81q/Vt1HLvWtEygT0KkPyNYe664cauoe4O+z19XjHhOZW82dP
fobeZ5pa41OwxIakJUP5KVvDwErms15t9SJTQRA64lXLpsUgBsc/mgsY3kwUM9C5IJON6e8I+phN
tKpPesHRcfmCUMRB6BPlQD5uJ4XnFtOrZXHL8OnQPa/QIf5XnCQLywvF6dECoBN8UCiuUL0Gwt0/
1fe4WrcCY/hNxWTmcI8jAAERvrL/zPiwf3M9zjBl3hsNtgBt0TscWTmViSjiO1GUe+ESwJjbxR1p
cxXkqwwDCKtTyTSFnbrPE0IPl1Ho3xG7j58UQ4rEU1KmmuSriyZr0WggRQhquU0OP+kcy8adCFX2
xqMcMP8wjB0+0zUmFh+DrtyJ5bIGGXGtrywwdfEqSEqAX+Q3ZSYcFnRQrrWwQlLy6LHsAyFSazrR
BCUWX6fu2c+SDYDQjDOStMpBdHWyVnISp2bEkk6wOnBVc7Yb+g76kVC9qQRuWCDcK0iVlJBDUFN5
R0fSi6xvoue6/IxMBmoxj/nrf7VrCS6yB41bpqZZnP1mRgQy6e1Sx6e5/VXw5qPc1yZh5/zM+4JG
vh6A9Q+bgqYZAclpo3SL0xFQ4KMo2PpnAur1lxyX6cJgAidh65ZnOz2VnxaitWN69x1rOZjN/pYk
d6pN9qrikc7BQ8/AomhYHmoGrSq6ePjsTzOub23k74gWJGHcLkq28TpbF+OWUqZ5xHTmX3wY4H92
w9hNSbmaK+NFgS2sBFmWZTogv7gHMd8BOkq09axH8uYg3suQfpkWwkLyCncXLupQhbrqUN5tuP3Q
Ko+uvMKqY+blD/4DsJk9MKeSPMUQ9ilfHlkjXH0p9Ftn96M9JAsY4mGWd/oTzhwXwNWws9eg0hMm
J5aVRfsXVs28KGW+zlapYloaXOymIvtAx8VTkgu7IgdvHp2ZtleNKCISWmcTOg0byMSCqdFG+JdJ
7V2+KiQHVqxGVEK8In45Taokm0l6s/6pRGOoUWwAYA5dpjVfLGlz1JFdYjy7nuKZZJ2jxdsyGD61
DDum1WeAYhWdJc3ORivjxlgR7wdqWMOUvUOk8T0ISEYTpunCuHjHJURFgM8sIH8rAzqUdRsdk8pd
PVdb5AAi70X8lcmQcnP4IH6dtfzSl+lU2kce1eNzx2KwNBKSoJB5sbqNirEzJ72HWfVQiM/5CmSE
t9sdtWZW5KPb20omwsbDgpszMpeqJTOOXRHqT/ufHbnKxIlPxrFHAmT+mYEu3IQBtqFiBa2Cuhq7
21hGSAaXSBsM7MS+QP2d2flKy1UbTp3lA0gzJZb93wNLAI5vVZ0STTJiBzlVWgGsQATppv1DvZ2T
2OV+59eVBKfyCNEKQ9nY2LeATQissFZ6V2KJ6xBLjeCtn9tHQ7zvcx1MoW4F+stsVIXyjX0Ejd64
EfGldYQ8+s/EYRMeqeEcZiJpKVw4VUeLz57wDVHvM0rauysWOReHFXLvlVS2erCSFCsjQn+Iv4Q0
yK/wJ9kaaPJ6DFKV3yG9PCQ/rDbxYIlacsWMwsul4/b3I6WgTXscUxpyB/i39THHmi3TFzTOhTZG
CZ4oe0NLkQrLTDOOrEsIFuzEvgJ/fqMWi1vkeQNJguPNel97abpVFQBI8UMsc6oEsEqA9WhvDPhO
lL+OGmfULPKZJEnbMYWfV/2xpEd6Da97CIWZPbdrswnVXSsbks1w07ZTyLN52uUI1nCBiHFsIL4J
zS7IokMAv59XqnXcpi3hV9GMxTJW5oz0SsTQyi/yAISTo4N/+CUZT43eSb4mRs+hBSmwGqlIUvQm
itxi4UL4IN0XcBzdMuclAYHZjcKcJAEyK5l3bZjWRRTkZgKXtnf3amIwsHmgnowEA0Tdgnox4n6t
4q34wMAq1BRwVQtWVa+fWOoh4u0P5c9fPpX46wMSD6ny8FwG6kBhwnp+K9ODM3JcHEQsoIHS+hUj
/OJP1FJD/vNcfJEQb8S7Tc0Ol30460a8Br27bp2gz/enYactZ9PiZH8L6YXiQcO6Odna8T7S4bHi
4DPGMX4xub3Wp8UGMR/9Yik8XNEfFcxzLvxD1Lk2J9gzvEu9GeoKA1+CMIoQ8Io5mKlKUAtBKkrD
D1Pw2Wc4HcS5Bs1NVmj9s138+euLMr4SG+4VU66/9szBTbPQk2F5I2qy4GGRY5yTz7h1VoYwg8bO
e8mnxi6S0xAdzIVVoMXNHDFbzz5aA6SIdybFcs3M7jqIqmA3MA50Xk2wYv0YY0w0FOfm3Nhksg51
S7Secm5U3BRD0I4XFCY28H5/FHWvISFajVnD3q7HmVgWNcESS129u4I1MK1AOx0yMpOAPfUh26Uj
t1aatD73uvSSXnNKUpDRLiijDBAteBzzAtfJe5W616YmclTCUhLdlvrt8XV5sUFCOKu5oLwwhpru
hTLIDcsdvrYVip62IlBSNmTHG+t4ZCwRD34KF/nzWYocloHwlEj3kcOkppmqP0Q59G/YF0foeQAm
QZ1ZSje82o8sZez+tazE5o/INqvcglhh5EJ7pry8kX4T2JfyY818qc3fddqIZMaQWJdzisGZh6k2
BFK3wmz99r57H5RLLexJUXVKJsDRkMYDb6GImC7iuOhGKDagXLAj7H95rez9Sct8dGMASmH8//2Y
ehzKhnZU3vJSN8Z497rigyJQ1Ti434KWJP87M9vSUXP9xBYClCbjLPwAuQnudJd8SwJpzNbXz0wb
fT5W9F9mpzjaqUn96cFO9DkrcCnazANnuv/aHgAy4241GISslKw3KjVqGAYLXLawbCuuvr2SODHQ
OVLXbs44reYg7NKcHkFqA3rYSprFNMzEgM65PrqOYld0HzbazN1U0UKlaEwpdbqf2WTUY9PDdZTd
7pt0qnLhl43ABHW8SM+VTdN2EFO7I3yp7EaLP/tKhYkFhqt/+RUCB3W7Ta4VTRIvTqHXGXdBemKO
jD4tRif4xnF/ZnGVGGfm6S846ekbrJ9HJloC4fyVv7aQhPmK5jERaLUAMsZjpgaR3AUZZniKu4C+
kg0Iz3c/KrzB96a/Ra+VNQIrIda2A18JaSaprIyQbQQNRw4W0EY2bnHeujgrGcoPLkFNkR2hdnRf
SD1fgr1GlyK5DhjBIX3Utr9AjgFwgOqUozsmwWcMXtuvz/uG34ZbzATbwZoUyDCg7W6mIkMZLwMM
zXHCdt9Pxv6PD8J0apHPDZeTDywbXGdy2LleGNnO63MrpiBSFvjqyrbDwDPALBxfuL06FJiMwF3Q
6qWFzY8ujxTtvLLuq93qUMFORypDAw1QhX08+wjsrJKLmh9R5o9d+z9yI6zYyoza+geLmFukx8I8
Cvn0hZKLnLLmvtLPA9+R4e0sb90n8jfTI9NYejiTDJHJOjC3Mbzm+Yq96n/UBLGags6spHIJnpp6
huWGC1VFiwElgYCFXvx3R2W34dULktfPbds3+WWJRprMleqo86vimqbfp2cC/RepeNksdP5+vHty
MPmCI2A9kO6YWvSEA93OtTLuZqC36YVa8qwb5awL3BrQwWmahLdit2aysi2NsTnwB5wKB7DAstF4
Nh7pBTMUwU01uSAdpCTMLG4cJPENbINQFhWb5f8rQGzwtBRLZUte5xvT9S8wtuUydzw5pjwxz5hn
W3crRI/ygzJLTn2oClEyn5bnpKjeKY1Li+UEgrvSU4jfiPl9/EclfzPTbsBMQeYpYhB+Q8QZRNOX
TckAGANlsbxobImpCNll3rdPtTDMClYg94EoE1/Ug4Yo1ZJYfJo2ahuUd238hoeD3usM4XIIqglo
LdaESMKbHeSLNm8jstVcmuggKMjEJqL8WLMorbzjUxJRz7aQS/EYIl6iBEsF0WjC4g7PVljV8hro
ypR82yOz4Zro3QAyPh8bBOPOBMV2ijJffLChUtCqSe5Lpojf+yMvP9yoVzNkn9k/bBnF0ggbJfjA
m0znXClrnuCUen4xUujAVnz790lY4uxEkLEDMAHgkzFjIuvDJmu12Xwv8/zL+gzpr+B7KZvhA6jR
Nc712Pq+yVIqqyVusdOY2q8DrXRL7L3pfUdKOsVyaOmkyzJXrX645gKDZHBQXB2vV2w3aIaTfowF
hoUTHUhasD5qsYT03idmLZhh3ZNWVC5LETa7VBlA9s3fTCBzEe9ZnNcTUkXuYKJPw2ak9ddjW336
yKEjHml8fTOcblxKy5XJZhwL1vj4DNjuTT1wzALnZmWNn2uYSaKWPiIKtbwaWGBM8J/UfLWdtQNu
TAJIt4CVm5Bh7qFqSpSJ+VeKEL6MBiilUqD5qQ4vKUYbtpzgyviAbqkZJRVOPdOLJBmR8BMU+Z+s
MthjeAqi8e7RLU5qnIJoIXUIFmg4eVfEYTJtJwJHqr/isF7aZJwffK67TPjEvW9GG9qKg3zd7/56
pbPz2CRAHXOCkMfLYOZrJ6YvEaowqVatmwNx41oRH9mUKmItwcmmltBj7dt96FYtB/L5Dl0TjdLb
YxJBZw3PjTFcY6r8e30tnra+7xD4cYG/IFWr1A6ImCgm7et4rt6Fg9UIIppF5yFZIR5KfAOL7S2h
v2P6H8apyQI12gJNZ/oqW//MmpJt13N00vN8Ogwajaae6ty6NswUaOKZR0WiLxA/RYCYHlcWUE51
wbv3BQ77nfCtJ87JSPEisP/c3+EQuuTJSzY37c52NxPkPGmEwaif6VBEC8pCGc/pfdFC/zPGZ/AN
XuzOLH9dFg0Vb+XK9e4kinGoIK/xy8AJ4RWaEqgTuucopDJa1UL4EXWWU5vZcQf51vFtn9bj4n10
EaZMS66u9hfBKLUZzovY2Q9KY19a7yvhpR3vqxADT18ElGYvj9lj727jubXmzTLzwejUgTB4Iwye
3Q34yx7fNuU12hu1MgPWQU5hMU2/hvqgMzohpuk/tZhMBzWodj3rLorzWU7biqfaeFLIFRdYDOWB
1MLUFEl6pVZlGLHRRcpYuzlrUltspJN91uXHlF0Q9Pc1VOWhuKj8y5/364ChgnIKOpOVdN1ayHlP
dpV/Kz7RFjOEMpN9OuMwOVlBHimPU0dEoKQ4iCo1bqsOp886ggmhw+uoghza5MtSHe8O8N5ef4/H
Vt1BiY1T4DauReI/+L60sGV4SSsDz0keToUMcYbaQRCLjN9VDznY1iAh7s62DtCeYVNRwD5gUZvB
NrmEWrjxBaCAyFWgHfzxR8oLk+y/Q7GXcmv9ER8bfO7KGiEEl44wYWCRRdWXNt3tiHXuUSRA/Lp3
r4Oc+G9AK6x6iaQDhv1+ovG3pP0biniD1fpSAr5WbbtelLKFJNQsehYT6w4C6hJnmnUZeylj6p5A
ByOUTnto8nV3bwQCpVlSNCl8Cmdjkc5Nt5tPAPKtGFgeldoOiKTv9PXJ0nEtVIYZqXXOyO700TkV
06GABcynP6yg2ELiYCdNLiMpDLEGZ7L5yc5Ga0SIDJdUuIy41bVHwWv/LttyvCm9376sCqC5AsXM
+hQxex42ycXcI9iDGK0fdLQpnbkPB9JosFckJ+qmOe/RS+y95v2bAA3WaNO/y3E1rq9t083XYKXw
K8AeCNXfYfdXrwJ5bgFtNjPq6mxfKOaVlH3DPwIbmuofIPYZD6zBp983HnB5n+jcJMAXHxd9pQe7
+Ox73dlkT6QSEdv/cUHo+MOnH9nRI24XNLwYoipiF+OHX7oXzvCm71Ratf2Uj8WGGH+Ld+vCZO/u
zW/xSYENORNerPh6M4tG1DUeI0BxuDwiCkUmEN3C3ekHG4m3mnT3hAAJroLkraO9gwWHLyKJo9um
RMptmJ90vy5WEM24ONQmstUBe9oErZ2iNXFIxBufRuo5Z2+rbkrFPyiuYV4TnMxwHbtSWU8LHmfa
fqAmCA78uFx7P7391NmPk4++q0qHCZvtL1Sgy/TRGlTzn5IU3fUbJAE3GkLz61LLrJs2mjDh4q9J
/8MaeSLl30KL0kNV69Wy14H7Vekf6fSlbUTUK/P947EVYiM3aQEbwePXKrlu06MFTZHh1o/N2ICR
xxMz2sYMuz37UJjbbeirTNRQQ6XC1s07b/KWjLc5pGO9GOUl4ShIu5i1eau9iSarjNRnxvFCl5v8
KgmO0PkJgVgv9O/+AboO2D5WrdYtSAGI+cpT4f8je/IHh+GD5C8Lm5hBqJ+HRjKJZqRZSSlmhlC2
GaOYx8kSXrHpmLNcZy0jGtFPGmWuxgda2zRhQJD/pv0zum8z25og1PHr1SDEI5EO3+6oTLX21MGM
867TwV4L7xRo6HccwzGLl9M0pO5bKg3v3lhMC1Fru8ywMMz9QjVk+oarc/cy5z3tEFRpWPrcGV/P
+KcKqJ1iQgiN9T+Pz/LeQcpUhmun99O80f4Nx9vmxVQ80mm8Wb1ImSWspDu0t9Al9nCH2n6sg+2b
7YBjpO0PL+QdMG1Zb5qRSjsW0gEHH/Rx9+LOsjts1sk9lpPyNAjkswOoQirJ3Y6JK5fF6ZanY21b
ppx5EhPbqBDZrmvLRdyqw2bSR8y0A7IBKU6uKV/EH1QPMl9yhi2dSFfEwzCs6/JhL4KmqfVAFsdy
hcLmW/Vqh3TheQXMLvNftuFPQcECCCh35gwdMNYfDfYq/ekS/KjyNMigib/6LC9dcAXbCiIf9Np0
xt5QJp463N0VOQZJCG5uJeCLS8ztOyGunnc4/Z3MzsFFodAfSlI1uH81+x71ixPDgbDaIZYs2jrR
2rzf53YRSoarcWmPiEADMYuf5a2mqAEiRNhvk8g9O1GQoOOFugIe7OEKJbmRTVSnq8QwjdIBwZOL
jjBnIgMgvGyboTSTBSWIkVkLU93ocRvmU0kjSLJN2z4+9mhlgTVc3J/uz/eoom548oXxm+MInEUp
rijPlGd397AolkEOZe/61L10blghWLj9b7maKhuIZl3s8aKCJRMT71dBSHXgQUEYjx//BJQuT0f1
FT8WiSFhGaJu+GCS0Pigh7FqR1AaZAlqQaCKsUXihdekxxeKy6yAGAWPs7p/qCybu+sd5jV0i+06
1xTRpa5ck/KEvclNzsMpdWC2Lezlzqes5po7nfyebDJNz0IY2yLQVx9LPUvmK5w0Q8zVWxa4o/gD
URtQJGcL0Ig2z90PZDBVeon9v1G7zeW3Rso+rOSiFNVdR5cZBXDaZunyhtzf6RBWE/bKRT0tSmCe
XBQDWr8c+7GujsI5LMy9xVJK4+q3qJszCAenfBWDHpNX3twdqFsnONr3+VJVoaYANpd8zl2wRIz+
x6p1yQtCB9tCTOowD2FXpOVV723PyyvaCndLpA4yWWnWZ2K2tdQvvOhwuJ7vDmRgi9izNXIiLIkg
u7OXyB4fXVzdhKbuApzxbMOg33CBtyTTQBtqDGZV29ObsgsyIaKlKJ35NLaDuJ9WVMaav3Iu8ckV
+IYmrmYVJupfqwfTjumxXBbBGA1HHq9NMN1ruQGFMb0pgoqP4jZ5XOkuRPZ4TarZI9BOQuqOsfvn
Pqq5YQJih8VjM+JmlA/7hB0l6NVfwUIZeIBs7ROZw6HDCuiQAtJzzfHtmNdpbxgw6GIwDBbsusYV
lVFpr6jnHxRqZY9vFN3Fe+1n7wH7r1j5IQ6AFGao1rtPQofwthlAgOSeFvYxbZBr5oXCVs5i6tJB
9YLwfY76Lyvk1NctXOxA8bQAJJYIEPCc2lYWDuGZADtHMGNlqGx0MkRcNh4b26IKLuxTJWx2FghG
NfP2E9PSQNK00FS0r30g8qIRbok5RUBdzVlCUnFdBpLSC0pQHZh92Bjw5y18EQYzd5hsQlQBbN5f
2c4fXrwZHwMy7ShEV0ed3oiVjA5q76appeWoRjjfk6kJ0ljrHvq52m/1ENbleNlY8Um0gVme53Ec
1Htr4KTg02xzdYJuqXSsT+JDGVWCvUYHLRCqkjwZpqkkZy84mojz4H4ldEC9cf1h5/HxLQTpAKwp
JV01JSWENxW8Lm3sGB6WtY1Z1NZzT6gVKGKwnct3AqFVup6iJmkT3p7NFI6Nkd4ISXouvpGf688n
LT32LwB/C5q8ZTAse82v28hTQ3O7bKwEvdB2D32Q8qXw2/4PbbLEIIjEK7h6frLfa4kSlVsR7nQT
+fj4ti6jiKY/NItQgmUNXXC7mcGg2/QHtI3KJEE7Mwl1AZN7mNRGI2ZTbd+8r9CRd9A2qwiuFWG/
Oj2xNNYNqjHrd2kLP7E2F6WpqHnEPB6H1F9xijhtD5ft68VsHXT8by1Vl5D4CGIdqV9eZ9Zg3Fep
bSC8Mczt5ooq6li0BzRAg6xe0wsZWtBdylODx88vGVLu7X6o/lcuKZrlSbqeguS+CyWYD+VbzWbz
1jYqkFKqujAS6BNUTpJUHPwAaqKvu+EUI5YG4QQ6iEIh11mx1MGPSl36vXjPTcDc50rIBfPtH6Ff
Q3zxTke20e3ygJbB9aVKMV3dsiTztOrr4XI3P3qy2uW1pG7zEXMNwB5dGUBa/K+3Zy4g6dPKfxVM
uo4wZ7FNq+Edlpp/0LA5y9DnDvvtInBWhPJ8DjDxw0mtrtbxjLmMUx6iOUXi6Sc7RAZv2fiPmsLR
9a5v7cPGeFGbIly3j0dCV7gMi3Rv6z0+QaCVX+fUEV3RE9BOJTG2/OF4GKK26UPQ3QJs0CHKB9QC
BKsZpdVhQkWDwPcRjBJ0SHWALm9mBHS1PZEgycJxch5sdOlxraIPuYhm8vrh4L5k6GPKeeCHkjtz
PmLkd7aEGWvHy8K5Cv9KKYdFlrDuLagJcXByqKaoorTMr2gJt7sJugEGfDebdErNqQ6D/S8y+oM7
xE2qzQnBQyBR05cJCv2/LuPnZ2KIaZc/lsvHeC20MDSfSC9ooNGQCJ4s40NSSthaPQ4EgDWhbGpx
Q24DfkYBo2vhzKGVXeZ3VGGweCSL6uuvfb+XhRD6uHgZB5nGEnWhr0iu/HON7RPbcqiQvbcK8zDv
Xurzte1kom0xsgUNDQ9W+Fb41TivZGyo4aO+6fhgLgSt9VmO+rhmFrGI7T65us4UyaPmvjQW2i0F
YRhXyPcJDKitZ5iiet5mkn6wq+E5DtdTVTVVD2ahxAvk74Jmwe5PWf3UK6hF4JXr5lbG/xqTclBb
iGSqAqbYq8oWB3ivbQDx52yt7gHD4JrYcl4UogvFkt0cIlyPHDIaYnTqGE5EdRVdt8dNAZDJsg2G
fajzlUYUoZzKXGA4fqOWkeM7gF60cntgdFYDnSDR5DaJtwGekwblEpt0AXFfjDnLQC28iAwGipA1
oDKBKvNr5dTWAfkrhEANMSgQkxQIdJqfwT92MlTDckL+SLkS17Sf8Kel6POiJtevM37n8ZwUDlHf
FRlNQ4Y7XH6wDiyuwr9k1OpbksKb2QH4j3CmpZyXj1WnXo9iDY8Taa9nbw4EY9bjKPqD+4ubgkM5
9mEMwDW15rjBF5j3X1npoCm1OZ2GIn3WEUC7Ux10Q6zrHtsnG8UViuDivtBx0R938X3I5SqNCK5e
JnBPIED2F/BnDdvSFnK95XYjh0D3QGUgv1dBjgaLAIcI9GjrXp02xOekk/HB5q91r2edgtySJqGD
Rgcr7C8jYun5jkQTVWYzOzygXMkESRxyTagSSLEPmuAX14lO1t9Ik9Jz3FOe4CMBbzKq6Ol7HEtV
s+NncYDiujT5QWaVc2mvanRJHKrrusbT/MDrQShLqDk3fi9N5Faa9c4CMXEFw4y2rZXqQT9c4Tbk
d/c1oeSF8Qwy6Squ5u8zN4UE8mzgm3TO5IYb+FPbzCpge2v4njrH6E2r2XP8L/CSoG3x8QQpnEiK
2nAy3futZOSye9GxBiL457In85yvhLFpUTPw9WrIc9Kl1i4PygGilQJ93s3DQH12Huya8JpaAoSx
hfem+jeN5EFsJalZ4OuCy06e3rsSA18H3u2TvFK7PAv0uoZXzK8GXkq8gqftTjCXXdHOWgisD2+Y
ZBYlmaxIcec69/A0xQpE4hzZPNJnZoPDHhRS/pn4eeZ0su1zfax0jEo/yNNg11plFubjrcovyxiZ
K/nRjsWqZzrfv7NGw/pVfXgICQdQcyCbZcezm2OAwI8OXXJJS1qffxIu96fRA8fcnKq/f3BxF30g
g4G5Qi2/UODyDxzrgL51I9ICmTZyKZDvwxc87a8zg9UBO3pDYuVWUHedbRC8QOr0ojAYOlVdFPXL
sXN0PSj2bsHFKbPCjaXR+7QZPoBLZB4ReMh4J6B+4hX8+DWPv/16evZxByIpHnk1/82P7Kp/uO0W
vWObxwg6ucWJIAFz+KrbOffCj1CAr1Rli5nHfv23KzgimqYjwsbbrnJwuYcEg42IyhXQukQSoSt+
umeawOUMyAajbn57pPQFWm7k/1kSMuoiP2jdruNoQJ1lpK2bMWuOuhamNcnhgj5t6M3kgVMVUTjk
+12fKn71voNytAuR9024hWrWDzx+MKdJ1aoWIQ7Nwzb47yr88wKB1wB79dsNLTeCYObCZ/HRcrFr
NSHCD7Y7gLJX2ARJS34SKkyaou4W0wn2tet7EPYPy3X6f1TNgyJEhV9pvQkSYTqQFl46g0s6QamN
spRFRYeT2VAYgIwG2XJf6pdI8d2kPllxMS1D34d3NdneJY1u+amn7hG+E4xFwHE9KN4MIcB8BR2k
HECe7Kv3nBDM9HxyYmFltFCWPowepCykoL02okbQsR3s69j5PQmC4iGKd4cyQOs0q13T8VJke0Zj
ryjmvAhWUIUTyJ1+9YD406KrIrm/hDMI5NyypZOpR11iT8XZUQ+tL8lhkiy3t6YLgTpR7CAzH9Nr
TSqK82xZGVRpzRp6Can8Op89qwE0lUEUBNIDH3FxjT08TPrUx1Hx59bDhRbtaiDrHsCklFhYF8ZK
ULobzKqLE5phAHmaxO0EZw+25HPG7lP4aigB7a7enXy7/C/Z20qKn2G+POv1dY20qQE/c/2RLs9T
w/S1dLGMw+ezIJtVKEgvBghTcUXG556Uj7dE40RocyNjDYOWEaRXYdFBxeeQGxXGhdBmHg/8YhrA
pN3TtsbCDZyLTyxDM62K3gd65Kz1Da/bUb3QctnSI/YIy+viPOJC7Rs1u7v4TPbrWd6LrTbyS5Ar
8uSQ7BYXOboZ6yCvm0nqbt5zFmBkgMkjo49Dh84pzn94cHEeMVE89pax16foPayjwoWdMa4dOdVT
kepWV/BXNpaVMDFGTliPnbQsygYXEcsHVAoYeC/1yTpsA5gDLvGyLff1963JcJUTcCC4VRVolGSB
DvDS0S32FQLsLqhJwmSYYbV/3FDhfctL4XagAvM9mnfMYCMrkHL7SaiqDliNdZzAZcMV+HdfR6J8
SpN8hIrqo/xxq5nn28rbQaiFjDPc91hGHjwM25JWzQuuHirMtd8eXI29Gao+uoSX+GMTB3E7dLoZ
1eFRx37w1qqfRDlP1hl+eH0AoCRtDsIyiO7M6EUds/oYxCumiQR1ufC9u8U3OWY8sKQuZULUn5Jq
iizNhThNR2QbBET2OyEH7zNFOaSovv/hi4L0sRmFcnFh+ms4mHeJNWXmGFKiF7QOvmeRtMDDzXvN
DkyUa10z3/mOmcekAc4pTcJdMIniPsqOnsGe6d7aT4Q1MVEdTg9jyIAngyCQV8jcjBB2/cTLtOwR
thRqk1uiHaHVctSu3BwHXOO7Ead7XhFMbkUpTGyShDfrc9g7+dl2cDxczIa0DpNCAUP3qM81jR/N
+9sxnRk31u6nUfVlCa9adQkEW/k3yo0MFdn/NOyqK1JkH0i8anSjusv2foRPEbvElgVc++1bmEKy
SlbwNhdyaJ4tL8IU882BXjYrji9vBIRgmAnvOkPPeYEtnhVHjf9Vzq7po8XoBiOKnhu+u4eacklC
P3gX0KOXDZ9GW3gHcBiUF4JGrtHfWdIQYpSK/oXpy/t7SwQXKir7KN/FBEyr+kwdw0ydfZXtywd8
jwaLZu2+eBB5guRR16n92F0CGjf3YgNw8yiA/VcozkmePmHc6yzztDwB8UIWkuX0I2hetDtyj1MP
bPyHFDwn8HuTX2mOlw7AIUfCQB9z2TMPv7mz7kGJrNazQECes9Ui5vRQ0AQG5i4AGxEka9TfGiXV
N0/qEb1QFvXgvv2Trvm18YBWKQdXCfsozVZLLzaLZELAUFRjlnesOW6ol3+vzDRR7ZSnrrzNnBSQ
sdqwsGLkPffanLNgWaLXDltRbvagxLYQ3fsLVLg10Far0rdqS5NWkdcJGXwXGE+ecJ4yE3Evr4kA
zv3CjUhg0ncqEsSzg6JoDDlfkRMjhK/tCfmx6lQlG/vJnkA8joVpfLnzFYdCO3hyGhZBdaSEb6ED
Zu1xhZpc6ejBYNN/7pSFnUrEEBCIfLK/ASrP4py4oxwWDHdjt9X/R0pessAufhm+MXmiAwXMSWi/
XQsKqq+YkUh0P2dI1a1njo9ey4/IIs+aysh9lpqH3IJlelAGTe/K1Sa4ALAQx3Ly4VG1Pce69Lfl
mAGf7YrMHAOuQT+lNJ7jaKfEcHepZ+ha4QvC+FGtNAiMup1VDBKDJ096x7NBG0IY/EEMt3VgSYcQ
U/Kd2SnEAsha/4DhEZ16+euXiOLANgDICTfjYNFrsIzT7gYiwZRHTxVptlLKW1lS+9wG6ME715z5
StRrjxa7HaoBCAaqcS8YnwACpFSVr63MI66KuxydNlnCys87Z3J0K5fXNsqsUoFIhxWuOldQvP2c
t2Fc9UcM5sw7kZvwbuUKJe4R+zEp6u64rMrWn7HUQMZzBskeRAPtN4U7noGz9fbO4p+ESELAwjiJ
/sDDm+2QTNGP+TdKBx6uO88A+9sL6ZIJhFbSj/tyAx+R4U6rFLog0i4IuMdiYbGP7yxze1vnUxr1
mMsqwccu1L7z9vpk35nJD76skGny/ifNWbVoJiHEJmvN5y/mCAnBVZGfJ4HSASgyt0XNvMfxL2s9
58hBLcT9n+yt/oL7T1cr+dbuOl6v2SXjZgZDoSiE9P+bTVubgxyyw39fuHLp+sTGqEP4TTyOas22
omOSTl+zYvZyaXyaBeNy7ICGFg9rc4H7K4ra8+8zyvj8ktI4TVnKyqQo+gzAm8p8YKLJCSaSBoFJ
XUHXRDseG1vkQvhMQNO3vnHyOai+yel9FL/0vSWlCHna0hau7VcMaQsf/KGQs8JnwBEAuiUvhpdz
ADO96/ZCvHHLHnDDUklpPauDdI1CGvrFJNfen9Vp/g5vwKLelI04Ux/Y9PwjrLYEHM8lMaQuhDG4
vxorvFZG/Ho2dxQ1tOeRHe69nmytqCHLDKBpDdDVvI1DMHnDaAD8opETzSZjafhyytFlNuoJtsxy
G509+mjxKP2flDUwdYauUD4fDa5VJvqDXIex7Y6yJr2NdBV0XOE3xab29TMWwhgaETwRudCcQT+w
E17GglbCjEEY01alm4J88jvBm8MsK6PC3ErjnaP4hiQzj60kburfg361V3ty56iSTqlpl4ZSHjQn
A3dMdcxS8LKbeLj7g9rEzsCF4XZcDJVPnFN1dtzgY1Pi6Ue1oBBXAzaARYqOyu8Qf5i3udZx0ACB
8Eq4xkWGPzjDZpolj01e3/i+rVdnMPns3XQD5k+W0xG86+J1JBcTAU/uZJNvSLwGZlmewZjaLmKU
ZsRYf2BVBCSuzCknchv9uhwT1BNLgix9tJLfxBAvojBkJ05ZiBsGj0pWIKgfw9mE8te0RDCgT3Yu
MNQjhTjkjLvwRW9n++ERShep6hajnQy1Doj2v7FrkNs9wwnfIp4KCOxmHCXXpB0G8HkwIj3x8zrf
6ZKEuQ9bIHaEPvCcreeOlnf5E/fHfsjXwC1dc7gR6OUHJsbTMyHJTZ+h2S2KNm5bTKC3uN3Cm93H
D1MT3saZCErvAIoxT+4lGAnBM8mkYqUw6huGRTJD52qnaVBwqe2Pk0lmXjrBM1KZJXVu68IeQ2w6
ZIOBlJS9P3xuBCvUoQwlKxXP5U06al9aglqspdDI3OiM/5KB7FFsPah70Rt8il5RUXKxq74O+TKX
3RJs1ROLzse+Y2/a+pvxwg3fsi9qiPnsPywgLNRh0AgkrjOmbxx9b5IWoLltz49Gtsfb135nvowX
Val4ySGOXoLR6lNQd/hZoTwLdh0GS/k1hS9AhI5WrEc8I1rYvjljSvepw4xtiWdOCnRLFmhYVCQW
iAHuaUs6WB0jzOo45GLHuGNaTrxnlvKdac7xYpmG0z2wLHnZ3S1pCRIyLHbUv4BMwg9CZMafulq8
bILh8jjNcT7j6t7F6m+RB8OyIwsdCYkccrsmZquDWCmkIVxYhfAwjUrm4LX9YPv9/vuCSICRAl4L
JHtMF8OWcv1zXL8a5z7IbzjliZvj+G2BLp1YiLVS/go9bWg4AMleHytviNy9Be/B9urrRWd2GQG4
T1LBmczJJg+ncslc7uXak6N4+mGIPqBzCqujyqAuHuINcwGKhDJAdLTUTEWcDFBEV0lXUtW7tAKw
TqLR8XAnBXgPfvCSa7vVksurqOWMGiOR1zJCbODWOUpfEGGW7vX22im7BcVhhMT1Rcu0IlOvRSDT
ENcD7XC1z3o34z8JDQF1G1NCK6lWVTAIHLhW2m4gg6JMJ9Sj2SJjZgODqKT0HJIilOrdI4UFtDFt
gTDqjS5zAJswHT3VydGhboF4abc9VKiDTqBVvO+2mE7DSaObOP1LlO0JrvFpHgQFEWtq9+78iB24
k3wDd0Sbug8w16nHXmaVR+FwV50a9jj3JY55u3TeJoYC8m9XIK2/egPXBWw4X5ijAR+z4MQW5120
1EPYSZbeyw2nNHiE8Bl6u0q4bEhSfnmItdmA7meO0wn8TkX73rPtfYaRJAzKby2i4JoKcJEUSiXk
mNY2gUoh7fVQ8CY8AtUWLn9ixH6xgGpRq03v0H3kM2KY23x2/rtSBXzaV2SBTi5i+vhn6udnp1OL
XqMR8ANJSLHOV0dp/2XKuGvbGHw12S47zobWyxPGfjycdLuO7fhL02NoDgFxfCibhvbLbDKPQKlR
OeZX7hoT2+04cFKarurdqWzOLKTL3zkPVEKUbYBdNoJz0QeBt4i25rvjo+uxhwSZYL03mff0TYkA
73KPbHMjLwhC94BT8u2hO/tNSH+iyJ7Q1Fjbwpr4i4W5DfxnIaqxcqOvlzMjdE+4HWTq+EEHvsBv
LeDb1gzyP9Jua9Tw3DlmXhNK6mGn2eZr8kSHHl9A+yZHjIS2YcI7HgGuLP+hgJK8K2CgMA9C+RrH
rEIa/TcY7cIhyrVmf1DGvUkCOhKCleUC5pWeVByU++iauJ3RRXVXzD4qZrBFsfe5N0MS9Yrg6H+e
SY2TvvP2/XgVgoLK4/qMbCoTwTCHJKgyecfGSeZExHbxkgD77menuS+FOQJ0r/bFKVdMe95yPt/x
KDuCHJ7EgFoA3Q2n6sK/zI9IQZ+m0XeftHruDOlRb+xSgLE2I0nghBpp2cNc87wBUpwQxcgcUddQ
Lq00jIWapBx2ln8gJG1ct/4aYucJfWEmA384pgm6pmwad3/ZG5Dg+c8gROfAHhe1YrYQ2+XsPmA8
XIJE4fViXM3ydC/eHMBiKq0lZw4T1+uXbQcLz+yCGkOJUYEl5Qu6ciPs8t3rqbnzc3ZA2/IcBxso
5vqClZny6hZU7DZLJjlthu3fG+RDjY5828nSzitfMrsgnlRdBJZYhO+KByBH6aI3uow8lmPb6e0S
yNv/QigHmOHzhf1350czemdkQ7ZDu5DLWFvN5BE9WUhF66vGUVTlaD7r63D3CuyteFTEX73PIjyG
7n3w9pBxGvw7MoejZEn06Vn6bbhW/Mi7kGn8YyTHGQYDFwF51B0CIIvyA0O+3FPhnUMgsJwHyfjJ
HzqAF4WWUgBBVUrPjowJCJybpX9o7GDZxl/4515Q6pBq8cExgk7f81ZULw54TJv3icFuTqPx8k28
/gAxGX6GpgHMcJWrZ4TUP/Jext2kF8zdcanr94Fl7owbBDVFH+KBo3MkUimBUn6ZKagp3DSRTOAl
hofOzcB6YKcmxOGWPUnuo7KhqJQBwq6YJWJ/AYOJ86Qj33qc4WUkPk3H0dv6Yc5M8qOwA1ccFQL6
q+nJAsKvb6qb+K8KFMBqNnrL2HAdetGqf640gP33xDykrzKQgb6cep41geKjKtZQeEx+fnKz44cq
iZs+Dz+dm516EGLcz2fOWwYmiL4aabhe6dPfGKOa9gxksC1WNfdsjReU6B6Lncz9EGSQI8yhyTU2
UZiVMYZzQWHW/OiKIduM0cI9pVfiNZmRErt9891uiL4Yi2aT4nn5DeBL5FWqYyQYZkm2l9svUKtP
9J8RdTkGcYSji8VFGQFO/ARmBMsaZ0OxZPrFVpnqM7OfP4cMDiboDw+AO7J9T31YAVpKOGm9hmv9
Kbdz1JzePxyuPBlunwHrQ5Zomiu/ZPcxnbMjR4gk08Xfa1Z2SoJ6qulIJV7E1Fg0Aq9tdMHu85ty
3vtOXjBO8VJR3tIuumRSzzxNmteuRclr01rgcW9yQOztHC6gR4PkEwErtLbUfMwhLswWZt1wUji4
qp5JuYvMHKVWz64NUiwFq9IijsOjaB3eNlLPNEVOXRYXIJbQAEXzovwKGQ9t4CbuaMgF80OiE+lw
79wwSpJEi5FYkufEfL05o8n8ZTbyMhFKdBZjVWN6AumtUVvY1Gi7yi3U52wMGZ1yPfWFQsabULmj
qNWma/iJ9M+yzxjhmLpDMKgLXBm3SB6FGvb5wiZgLsmPV6mQ/pOuwhPhAq1KN50r7WwP9TL4XA2O
qJDx3Wnsyih6SSfIudTRMwSEesTQVytaD4Nm7wdlX45Vd/0KgQf5PDoOE5Gx1GvYFlKZ/6S8GPVJ
yt/ntBqz+S3M4eSqOHHWFZCTdnZ1+r2x1UJO5QhSOJEmnn9KHUYn9CSYeH8JqkeNkI2k69lHUvLP
7giwJpBQICmkPYtheMqiCYhsUeRQY/ptMrCkosY/M6dg260rUChbrcn4X/5UyQFD385/KZeblmgG
aFNJgVW+rOFN0yv1gDe66TYLEAYXzauIVezU9LMtnH1mRFIKq7hhSde3USITBaM2VzWLDTokB/ag
fFeLQGyLHSL5jR4gl2kxmsZxFg69+hRtgMEipRhbmC18Oha5Dr1jZo/hg80+O+R3PU+Xb+y728Az
sEhTO2KIRulZ0PGEuYR8xON9yMeOdhs8VqZReM7T+HPImATJ1sDIpcVoSQlxB2Zfw/KiS1Nv4wsk
Ct5WjzPk4XrHmcWZDDj17BJFjCxJGDadyUoBtftJ6fR2AK0ue+fD+cCQ6mCVY/gQdY9kWFXCTuzv
I+DO2rkd4JbY86PzY9Cqznp+e962ujRpZYyDOne1ICHtgpKDrrjf6b+S1/ROigC1nJB8wIrv/0+n
KIlcAfyZFtY0fvwTR5J+JXyvRuy7DHZ+7qO9T3hBOR3Pr+OwawYGIJcpPsmS6bNE2IgefhEx4hf3
EfdqLnXpzc2mtjJXkpPoY/s13GgsqRH2X0dCjWFHVeuJXj7Q5pswtBwui5LxGJR/Ivekv7ZuhGvg
NCbLNnn1DltFObnAvaykYhkeNtcSzB1I1LTKteDv3Gcpg6gj4uR9WoyQ/uQr3kwf6B7biQJpflYU
q3NhWTsZF6YZhC9N7/T3PsE/6CsKz5tjBbaKUEmrC6TkHNkFQSWWmq0Dx6hQU6YMxOWeV4j16cQI
IX+VLVI0GpFI3V/hjjb5hO5YChMyiqqVF9+2Nug0m1PU1RwkhOoXj/micioZMGEfwfm91DmU/jLS
CWwFZBVK6Egjjn7/D9ph5HpRiAPjEVY5qVvaPN28hRcxXkB6bmsDUzQZveTo0MfCzgp1Td/y1kwh
912elXVxAaN/mSg31cFDAL5mKBuOoPp7oakVlbTM5mkbg+q3XKI9hHDR/L06fP+YP4ixzAT3AjOy
nzp8zrTNa7UxEnYobPwQm4uLg3IRAedSzQTkVzqO1gY5Y5yp30PfsbupCBKLiWCRK9QV3RtCS7S7
16c8x9xxIvMHQBma/yT0Rjiyedmdvm0bLrgerwFaaIjHY1I/2qSygzmbu754XvLT531jCfKrsATQ
dfvtgerrOSeFmhqY9/WX63avD+9+6qBjElxU6t+tyjciPS3t9l8WenonEEg6NrXUnWcxoGoDEKVU
Fr8G0Jhp7LMmx+9V/eV06AquqFH+b05Ieko+jejNz/6ZahJEdZ8hU7A6DSM5aUshn+sKq3Kvm117
hD4MTlNCAvtPvt7wo/CTmckgfYQCChi7uwaybsHCEsGzFuYKVp0cTF87WSjsDoq67ZRWQWkS8Jd8
Ie/Bdkr8XaHL+1R7d6Men97GvVKUEC/Yr4cm7e+4ncni+Sc6dFaYsinJDsRjWvxbQV7+w3C79GEq
P1D2Y2kaGxwqz/kvQBaysiNZ8BDDhh/rBWIaHv0rlmWZ4sTkRuN1wn8s7XYoU2tLFDLARnczSIjm
8wesz/oh1kugqxArJA90Iwk79Zlc1UiejpgfvHCtY/sR5eeXIxv+X4w8vR4c0hDaCuCbg5/k4uyX
izkkmcyhw2csbnzZ6+Yh0Q8GO191jZVuGxNVFgT8yreG7c0Gh+EghJ81s1oEJEwPD9sAznqc3kDn
L5sufh+FJdnkoWgR24AosuvNCLn762Pbu74/jD7a//tzhwYoT4d2VNVX8NqTikwwxEmW8gpyTd8B
m5pQuycsGz9Zo1yWUwf2TOPAXLGdcPoNB8yGBGkdkd3hvtXtVS8NeFST4g36WSGJ/3lX+Ocidpr0
lxBvveMHlVIpbVtzvFgnrDVu6LtNjE4yxJp3KHd/8/DmWFYYq+S2F3ddhkArOsc7rKAbLtpgaMV5
aNQWqPaqv8DXHZae9mpl/djJcWfqERHhvCgIMquYnTNO47jrLmFEqdDnCD9YK1Zr2PV3/fnqvBnq
5iTtFOGcRbc5Q43DC2Xty4rKgWJs4Zw9D26URF02lEMyWWuggB66gkMBT8nPMFuyC9SuuR4a9Jey
dmZReg0fb7Ix7Mm6/oNsOUiCDGMtbhq07lUQ7/4kKP7/omm/qJ5jYydUtgvlJXJS76ghLWVjRJnu
ZwJ6VyaoXR4tY7boJDVPyUic+WPYgbjQ4FikJmyC/y8/AtKB0ra536x46fvL4a343lObfogCyxDf
DhPf+fXHmA5DoIOGtgX307iAV5o0ArOC3Q80601TGeXVibONGUkh00Dqn8SK9xJxSOvx2KYbCoIW
kfl7Ts7E73/qZmqHkyZ9ynUHFCQJKRY7tcpNguJCDfcZ/V40v0H+dC7VyvP7U4goYjyOk65VSU+8
8C9f87Yprd42P+fzaO8qaiWBk2NCzEpP1mUJgoJ4R7XC5+39wNWCGwzmJ1x/OHPw+7UvpWL0vmT4
P3lhstWlx7DG/R5GzP7vEzVhpynW227bKXAEkhpBL+Dd1gTyzgxhyDPH/UM26LcBV6LQJCDAypXd
lL4KZZJ6ghMLKKm+Zo/fHKXekUr6ZhD+b/SO45umRLumLF69i/ICSrcuLGIfYrq1iH0vfcJaou7h
fKPmupyho/XWyEy/mUlfPA46NFIQusMLB/++aI8d98zFcLuX/mgsnzsBfui9QP8kdjC03V2MzOsN
6olxzJg5fnP46tGa6cHktjrxIQrc1Hu/y6+pkBsMXY/gX3ELCafDGOmerS0nbGfQ8YThU12KOEWI
S+jFnMN/gPO7shq7iwkdq21HpO5kIVE5pe9AOt/kd87Ta/HvG5c3eCl05olz0MmZ0RJR/JUiz4Tg
zpA3+JV+vXTkW2WJ3n9FpmInTT1Ep7YwGRim8zU0QP+LLWbP37wJl9VWyyTGZKZWk473232t7Oxv
LKlckUsmLYX6/0xYu4gdI2wv1XuNle1Sif85yeXcpzbKwIAcgZwoCNd1xgWAKdHwKjjOGWl35MMw
fmB1lXuQI01m5JUv0FJTIj/Fn3E9VIryvoI5gfXP5ktfuxhPqvgtYDn98oWfy08iGQ0gWUvbC7Ti
TylBSM+GvwSKsFr0b4b3bbTVV6+VfdEVC+I49kyoC4Ny/mVB7X52m344smHs/7oiUfCpBlQVdNm9
+1iWO8/+v10VlhkDJgGUEcSmy8Ybt3yaep/ASChBGYeOhHjAbq13qzCWGOhnGCCSTMjSh0AlnT2a
XRQNfIXpxQ2Y/R78g862z+m+X0qD9cYVuYdLLRMrc2tf7q5kFS1LsY8BUKGac+qgdeB2mifImKNS
Ftmb5hdV4iDnbhJKpUxr8whQXnyHeiKC5GZxh8a0Do1QlIYqPFnDKsR7158YuMm5Y7WHuG88pTAt
dc5gfupFWwCGY0c/ZsQoO0VSSnAKWGI2CLCO9FSNsfCe10oEq+oUTULLT+BFzOIF5X87pTr1DHou
lGvmUifBTT+2dL14m2s6ZMVawXHm+QDH935o0b0NBcr4NV4Ib8o6YNWG7lRUMlFmW08DvIYkAGq3
ysJE2jWOif0f3TFAmHSS0T2i/nw1GGn0tEJDDmBnKaw9h9CT+dtFU7JzPfi7Lipt/BqwT2/WTBy9
Y0pd+3nAyKYqF43MP80ne8iLbhlYDgrti1DKIzL6yHOo0BUpK5mYgG1kd98NHagJUogs1HOsLK/0
sreH103bxScdOLU+t1nI6Xfc3U0Ndfus1ylf5Hq4ByRTd9uvmoAx0tYYgngC8/fMKL3Chn8FKqS0
qgNDKt0jcfBrOMRXKSVb42mjnEez9rs3bozKkm/AlX+jtznp5IVsZ30PnHsH8/IKcfpp0WNGGvZW
PtsKd8zLL1Zb/n5eYZ9hWSLF95Z3IcCGnpgN8xnkURiAMf3Gft5AUu1AY5GOujGANoWwJ9B1SiQy
EPDEaTGwN6uRf/KMhB8x4G7nU5jZBY2CkZqif0iS3h69wPUOrxoSTOQmMUF1gHWn/KBCjt7zXHeh
PJ+jC22qDhU2deR0r+5emceEHi2Ew42FHMZr2ZwVm+FEKm1NszowgE0g7E6Y2xp35tWlI4A2Y+CS
9J2+G7Spc61NRv8kYuqWkfRrbYqwYSmJKQlaRX9dUdwn46u8hWjKUfUf3kxhoBKTRi6nnuBiDoWz
EVnc4noKDtugMt/110YsdVfBKhel25s+iKZdhXnUvpy5fQ9uuHX5TQUV1DzQc+JHH4SnSjXJTjoB
qJppWKUVeiaTE7BF4HwxAlwPEmgH1pmYO8utXfVEVZpg9io3yJU/u+mZl7PAnVxvJM0SLC8pHzwR
RQTt0I4zknvg0Xed3NLNIev1rSd4XoWu98pMHw2L2TCm4TvoJUtpqXrizOG1QRfwd1ZQzpFvt9SK
rHoiZmaIp6IQ0VbaEpxJdoICJyNNIZWcpkrRNP6XGqwCOt4u36Xq8MxcJytm4GR1KaIY7eMh0a9S
tVFk+f2Ak1Rnaz2HsI1PcwbMuz9EkHlJfR3OtjtNySg+eWkilzvMtNSSzbLm7b0kpSj2UZS3vjoH
OMZ9liK1G2/B3I9WJOihUC/sIore8MpTKDNJGxfBEP8tv49dU08SfOxQR4dgtH95SRlkCi1OtEUF
obiGvRzsZik16APW3y+tzwFmsYmfU2m1Ixdvlu7xFXXYMvlb/tuf8K5Rn5YiFPZ72AbTVANVl7VI
dOZq4zqtZoq1WbkI9TWz8LSG4CNcQgpEkDCqIbkxnarvGBBN6ANxbxKWwDb/IJDc3OV5SVZ9FQKs
Hzf3dU+vPxCnMcgyn/UFGLg0lU9xtC067I12pLjKn+WNVJsXMuRC2SGolNZeLSxH89YLHdFOklcZ
9M+qyxCXiwrKQYvwRceg552JHNYW0fXcmY3Ab6cfZmSxeOzu+fhRx/itGgIwT+eXbDbXdSKCBeZL
8vGJFM+Dh8eICNhtlIH5TmSAJJfvWclPHJCcwnszA1iMhv3ouJ5sn5cyog5IKgZpweKmrYLaY39V
N5JD2gvbtnTjBmo8SUZ0hsw2LMXS6gpRfTpgoMYs5D8OT022UVFaqFlAq9m1uIF8MeYUBzVyi1B9
SjAeUY8JfdhAjIbCtgw1NFCPwXo6Qe6W5l/1JwO3S0FnoaRG8zYw8y3kJalBAXdphSdpCEBXd5NY
dRzdSXsxo4PGzSqBM0SpQmZz27uE1NaZM3ltHlrcJ0FD+nnYtF5blOsLnwJu8+aReD+o0KzyPi5J
5QRF5X7t/Cagzp/FTVwqNiLs4SksrhrziHdUEJAboHiiQO2JWzqhIo5TLcC25vmjOu7qaiJiqeus
46oQfkaierSymdJQRLX3scXMnPuRAyBmRFelw2MsSFPbMkbiHDTlnFjgjpvwv5PenOCk4QVxL72h
y5W2pNuryGP3geMm+JNpxLb0t1HdqEwjUqEiIRYy5iLOd3sNmaPH4WqSJnzUugwUr0TV7UM+e2+A
PZrCtU/C74QK2/vXXviPUDlMvNeCNnuAU+LzVDTR6jMzssomTlw3eswf+xufM1AAPyJfTp3+iMN0
LfMEQlvpwfxkhcggeByCkqH8fQoOqkgNzbgk5VAHeLVtLbOyOeYkzM7Zf5pf2VzzaYPUtQqs5ZZB
6ahvyazrLodJW0Mt0s8yghJFUphOpjY3yRWnNOCXx3RSnEzqCfIT5Hq+9AQQ9BhBZzIbHZZ5ALCC
7QUYq75GvJFNxyxH82s4r8npfknglGnKyihgf3Hocs4CyPAFGabqu5hLVIlgDBoIwKKSPtankVbT
IZFduhcuQRl1iys4Oq+Tzx4HZERK6QRUHkLA8ImEmABqwIXC6L66/130ecZFpDrR1aJ2+svbktno
1zFE7OGTDBiItap/uosGC+j+GYEgzqUioa1v87E28SzpF8wNsHDiEh82f3K+/u081QmnbsY2QlKl
yCxYPPZyRZow2FG4bOXphIid7pd0OM9fPl1ceAq2/enJ++8HyT1kdypSWmnB+5rcwZofh04Dpoh9
7/ot2qntfFufEMc7HEqlL8LzJ+5bJoouuBq36xlAaKUolfwIzHcOWbd4OMkKcB/kUY3bvBC/P4NZ
+qW0zkWM/KJqkyd/kzdCPbRoqeFo9xCx+sawfCM3lOdqeR4oYs/yJ+W28WBwsL63sY3/qfNpWMIG
oyxhFaK5dmvt2RTijZ1xmezBeuYcJzSh7ES2V6Dy4EOgU4yiM5h95KoBujRhf1AZWHNUwSRcCOB7
qQTpaCXolQirTKUAZWgGB7HbpVIx7fY15oKhJ+xZs3SsFnv6jHtLQ+DP6r5nVbYKAD8oomj6MabD
ZX/Rml/3/6Amw6bwyt+libwofPL8Jst15wmt8HZdhMuTdckWxA95V0wlkqC3IGJARGcOTruOaGcz
CGQa5A5T56/kUb9Z5UqdSThPA9f/oW0gRMzc9+Az3a8lXSC8jq9dddMJF5OWMaSa8jrrq1461fLw
2PV4Wx5gCnsLk36Cvc8stiLjASreDnHzvJt5GKrrTlafsBu0dFTvnUn3/ykQItdb0PX2rlpkHLUP
RQnaJRDNLtd6AbiRoGhG0alItpogj5n1imsxCdHPhC8qmEQiAexAzNxa3TuFq0mEiM+nJgUCD4M7
4SkVnShkhFHLygALeuUjYy3E8r9pC1X10RSMiQNHQyift1pvRziX28E7j8o9aHa4CnwfJQxVat78
XIORbQxXaOK/4ULsPtJ+w2PhhpzlBFy8i6B4GG9dpUJ3Du+4gVuFGXl5TJZbQv3x+djQjsIfbyT8
q0yvceSLBz+DHkaY4RoHQkXKkgrm6p3D+6ECHg+A/AQQMINjnrople7HGjT6oQhboLAh20fpv4U8
TrDoJV/khgCDJNbB2KxkAwgJZR+7elCfp885NpoSHexFAswVPTCt6MRa+1O1FuhwL+QKwLnasfVu
QauDmXcWIkVbMcgaw1oO3RpNTmcbQuAzejTn207nSoM0oS/MqAcYN+Yq5XQR1Ljlef/o4WbLv6dc
nWR5x/qVasWe4zwlQXtoc8bdmc+xeKex/KRoIMNjuApRiNPKog5f5uX1+W+rbX9LK+Hf28f5TIvz
OjUz019CemrDSs8kUessgTAsreNKiZzIHqca2uQxkV+UlKTZU9+OHWC0zBC20Cok4/NzxpdinrW+
EJgK5GumxN1niVrV5nyRo3Uylz47GoAuYAcUAwocJDl7E6UT1bFmkY+f6Ky6ArNkYJKZo0Hy4HfB
QBiW28zAC9W1419vMsaXFMfcDUPd56pi/9WXFJa/v176zta3np3O8zsuyy3iL4TWquoUlvr4c8VB
Kb3FduBrk28t4HRHhdr/DBKx1Rh5Ht6jn0F8euIHORIjbFO/hT8ZCAmZBhOC8t66Ld8qU6OUrwV6
RAUoZtyf4EuggBYiAowiKAG1sWvXtmNbdTPRPOOPKZHx1UnM/leCZGf3mS/ZgUpSD9hAWi9831qW
KUHB9PipqRYoQ3oaT2ZpmDDmb+Cj9HtvwBpAhZz2ZJPVi4bj7oHfG7suurgBd0NHkPlZtGLkDCxS
PtifjsYqWw5mD0PetnCzChFKqQ1JmTdua0HxoGJAIlUO4mCxfM+eZOibsiVHizyyrnb+p5Fuf8oQ
3aUwWBUeU+5c/IkZrJ7HtvWlLkDhxV90/kuXUrYDtbS+pPC7/3jWS2gcRzGNvS0UYt8CR3cPGbX+
Hbh2LqyH4O6IwZ/k5d2Sqa61Q2Zfi1rM40/PNF/0mmf1AaGwAB9v3uQ1kQbnWzrTHJXC6I68HXzW
qgoKftk4WvwQdWUmCY/ZzLqHIfytA3aFeD6iYn/E73Z+CsH05dGNWmjtXDzKoOryFzynzo+EpYuW
y9NzdwqO4R6aHxUEbbNCH7ky5iGARQcFjOhWNo4+PZtbPKwWBhIxuG/dCO/0FZCh6kJJVIcTUuZ0
oFiz8yiWuGxsMKoPxkP7cXVfkf2oSv1W2DRuhi7nDSv3Tzb9UDvYTGS3Ies4Y32vooqygKVs8DhV
XBokB7MVGhV3sa7YzAlADOEBukZtdpaXC3H1lMjnD+XnjhX3UQnqO+fYrH5+QNPk6R8qbYcuDOIk
MSCo97sAJ/d2okwwttUF1ut7dx53JVTTnVVuPgJZvS0z9dLYcaRNgLB/UGvuogpB7bCD6YJcLcnc
1Di6pmUk99nuZJYWjurlpLdhN7s08a4j9xngt1vNH1NgimT8rRv8xxzOzUrqVm72E3Xmqfbyjb7Z
2zoT+37Ri8wNta1ltm5LlFmGs8ZKGUfXjnTh0PBEwRN1EyURd/ICuzJ4UoqE4t8nmyGLT/9YsZGx
aoxofvKybkH7ORQ/3b9AM/7cb+Bj/j9Ru8gY9XKueQ0k/Uuu3HhSSrwVHlMIx6LNiseA8JkI+3qa
HDqFSF/UQdvNKPvkdSkKqZ22c8CVXgZt3Q+j9SxEBZ1iwwJ/nZzgRrD38nlt8CzWn2SqES1qOhVA
1zn5rR3D1WPeP6ULjSrqehEiOjTwFnERtSKkucf4bgFnoFkFUSL8jl794P61dAU5nF5byDL9Uc6R
y5laotHI+o/M3TeluRzpIoh6DAYemUIKwXrQ7pMQ37pNrZZCCC0+CO6SuNBMZRlFo3dK5FkZ59nM
63kONgGHPR0vLC46hnyDsoIpV8olHrIbpnxQwuBVylciiRWBkPtEcbZrM+oiBdFbS2qTLOXxg03J
pGyAD1wOgBoKcRRbLwYftXEO2tkaXEZQcfsT+lXV550cmd31Y2aoQWYhrrAgQsvjiDwTWXbv57ky
WwGNJZb7bJkrTWNZ4zslnJGOtgHawH3PYcZQ3iMuOSyJ5cRIa7jjhoY07Ln+inV04nfeLKHxpY+V
9dkrrXP4jCeHKc1jY28CHKyqEiW58liGbBuo1EYqRcjohtnIH73PMqzcvOTxzgjbWUyzNghBPQkQ
KRo6VQFNdOewtDZC1Rd7Ug13TprWEnQGsVuCZ1/eFC7HI9NPXQWMPlJgRAvvuc39gyY+2O7/If24
flYvWEuYGDFI3jktmmNveRWOQ82X8SIO7mR7qMiG/FLEYz4LH/j8nWj02B9qSaNmARTMZCtmy0ab
f31znuYwl5cMMGNS4ApEtU522wFfqEGX6eAecQ/EEjts7g+RU0SrFfJevaHm0IE+8zXD3zd3lti5
jqDwoy3AXn4dpTb4DaGNfH9zHeNxdUeKaRyn3e3Rn+cxh7AQC/uAbEeiYdlqBpbNKrvFlngV8OlZ
0sqjo1ARzA3IsuFL+LewYE5BfFwfbNpLF3MUbUWvHD8+jie93PTIFbYr6Il36/Yy9R/CcBW21kX4
j/QY7m4t/O/NDnwonxBEvc0BgOPPMBlINyMof38meLKiNY/AJ3dRT2jcWqVMeUjmR4dFi8yu3H6U
EJgbUp8eCSGoS1sOjZ30GZ+64HF3ioNZg4q17kAknScvkg0Py+xt4QEM4/D6dhgXTq63Rdm29zk7
FHcZvS5j78oTkB28LyQVdx6dIdklIDnT5Rp3tblFLxYbbdFg+sthpYCGpXGp9QY/MOZ5ULMxnb+o
TJCCT6WFhMpHdedGHzMG5ADd+y6rwfHj1X1kktm/f9Innnyn/mjN711N+0gkc3zw9az+v6Pfz3VL
SeutK3CcnVhiYBzfuIR+qVLdd6Gako9Le4u1/YPmxP1sUCWuAyZtn0/LoWegX2N4mn1Sy0AQcfg7
VGQiPOje9daEidcYTbz4fwrWxewbbHeYqxyGk89EHYUZpGNSKjOSx85KgxQ/VO4bIfHyUi9yRvKb
v317q4qLaE36lKxyjftOnLGOQDB5oQOz/SasWJm//mqV7eq3SLqBHhhhVUw12JJolMTljnX4PD1q
YYw42mxgG32gJ+kr3nzmUwegoi2K635OC+SZHQHwje4Y2uiw314qTO2tiG65IptnKpb/3Yh/1hF4
V5EAsBfL14/KgvHvBZo9WvFFtZEr8fdN446nEfdI5h8Hm6hiM8EPOgMZ42n5rGUoC+4VTPZ9dN/S
8BjPDf0+tv0YiedIhLBqUUxdsrozYSsHp8WM8ExgosT71DePoHRzEpNufDlAo4Gx0IfbIg2K3/M5
EkSlQcTyF+2WdPykKgcGxMVIE9e0OjLJOdpvGuG1NtUImt1nxv8+9iJUWCZ6/3w+bwOSYywWU/Hw
GHlSjHkWfcf1aqgD7rEyuvCRGU3MXVMyO+ey0psPJpODHTlWOZq6HDf/TGIccpPh3Z9a0nMxjyLQ
lUs5YEIPbAKhHspH/H/k6ZTnMevXOT2eL6KRn0XIH7zmm0SIw2rkcgR2SKF4mVCPGhzLmjf0t2Qz
Xce+52Wf18FdEId2GtYS4rPgJUe7fcQc6afRRLkaslt9WFTLWDuIt/A9tBOwKSAGbAXdf/LeH4+a
YmCiXaeLJqxcbccUqeA2rpzOVatHh5ApthLPhyrN6UKP/1zHoptCtjy4uzMk9eoOr3PSnaN1oL0q
8PRvLuCBcuo77+z1KT+QR6mjw8Xv1RAWbfCoUXqjlwgJ6GIuP15o4Y1BUMqJIDvfUEJS6DCVbUmQ
Bx63e1xwYIwGR3mgZp4kAtLj4ltZZVlaunKS1ywpv6MuS1u/9p3fNOGdGqptfJ6klXaFIc4u5j23
NZTEN9/x4I96xwGQCMxStT6Sm+shn7Hcs4VRKCUOIO4RdXsk8kBLa4KV4Y34zibXFsx3TRQu96Ak
cgSiszNaXnL4afNkZHJEXiCX/hgJguelhKcvJQ3BNPAlWZUnJ2qRgPchLmzLhDhdSqESkeSLqa31
zS4rrwlRCCHpWvXnZXz2uwgXUBWZCVIG3NkLgSEExktGStxnTNWorgwReN8ea+gJLQvY1AV2U7xI
eis/2LKx3b6xcZcoC/EjR1puHIG05Xuu/nJZWq88nPNys46Y5d3s5js5oW5UvKK4mnM3cavE3EIg
K8Ci6GiwL58EMxar5NkwCjGSEv6FTvzIfE7PE8s+qExVdwBQhim6lsxORHF1WiQKqwmcPPmIAo8x
R5ck++5e6MJABWXOfHDwfR9KxxaQVb7RSiqh+WjbmU4NeLkJ11Gu3PCkxmeYYFFVFZ78iIPFFsH/
CtVT4KD2b7Ba3jk6uQ2OpUhOp1QOVG3HFDAXfYgXb3FQ7jpDryWT6l3EUCtf3MgZa2xG+YErP9p+
D8j9TWz6Xop1+lFqmArTog2wTDBY+Oy/zHNh1bg4ChRSGmg1PLmJNF9HX//8cuF5BZYDkcqU0WDo
YIt1yNQuc8KYmLl04RpVuDnVVB77E14kq5uTTswWGYVf3MPGD+258914wBLvcLXxGXtyB8Cokt+v
KW2lC7ZgnYLpfmtae0b1RXbU8yGZp+6fRnUlHoNqvm3IWsEgLShh9VN3ShV8TMbGHA/5P6q2z+iV
3mpI8H7XH5s8OjHpesWPCAOX356+tJrHbx944gzg9BVysXEUXbicXWQc3bPuAiEdD4Om4bWTLDlH
AupkXYnKt+RuLWXDh0JYBZJyqtByu2+q+y1bBgaicU9gq5DIuGULrGBqWLmepq1NyH9HHqQomoKi
zf1FFaf3EJvIwu2NvJts8mcBkXUtpXW9iPNovyBpRMJNTTE4+JHDwNZ8mE2TX9FlTTd9muUgmNh2
34t+9QCtEJ7tDn/wCi0V4kc84vs6N9nighiWGddvbx+sM0STIBPZrr3/k0LU/UH9BPy+fnsYcMTf
xzaFQRFmIurflRQZ82qz7cjYhZQ42Mti1wj518TfPHMqJki8sBFKoA4WtK8Igp0lnpm0ZvI0Dc5m
ktTJlGSf3azyjw8DgBo1ou8Vi5/BM7ifRbTckrUp6LRAWhIZlfh3kWV8E7xvt25euAyTy/WZhSqJ
pdpojzAzWR+kX+K79BJcFeZUwgcKv+qb1ptf/97e+N2HXMXnXDkb/SK/URKX/MF3leFEXYSsaGyH
KQnUw/27A5D8PwClCfnymuOfFltuwWKz+NVuf9UL+liJjADVkGCpt+PfhVZfmXer5Y1lA05Ckvsm
b3T8ya3dpxdwwHRu3glBBKd6fpOIIMwZ8rJvztzLO5TG1w0K1G+IcbQrIBSDpcMG6rftTCmm0aJv
kGKhzdfKtESpsdUSAgNFcV4tOetllv4Jgk91BZJXDvn5diwiaelt+KcUU+7KyrTSzYhdyhGkuO+W
MJtj9CHhLWbyEuJ0HQ14lUoJZSEqWHa6wpHwddCbYX1OovZqjzeykIWAEMbPbpn/Y8aycboXRQGD
DMXC1PXelAG+jN33iRtRAJbBDCMuzS8r1o1SH5hIQT+l0h/VJKRwMmI7roLvPpYvCSJvsx5UvcFa
hfCG1QfLkIVe7ekQEmwT1g8KFaLnCppMviHYhavVFToj3ty9QvMeaw/7fsIg+Voq+nxhcaosY5xu
kyaRLFh/Ic1dRikljSUTg2o7zD5zmuFEY0XRollvtQNd7/SMAdWwPr6GtRrSSmDhlhC+YBdpBtlW
zp0uxMrcXP+mYSL1F6YG2sJ5VqDc1zNv+YYm8XsgcNAzvJdjFZZ46gKacuWGSjkl3eVL34dkytJ0
bcSrdtccro2DHUdPwXguo93Whdmd/YbC635iljCn0aalSj/JvsTP/ke/zDWC/cWXalVE2KW8suFK
wrBbKi5ZJIGKDIbZAI+p3hV+YKUVYUGnEpKiVbvsVSDz+puZvYwMlrWbid474UJXnC4fmr0ICrS0
hyL5nfVjCnGbBKDTrnalzv6F6TU0PlUQZFNnQ2CLHO72vmse/40HzSemSOEX/ULGVKfJ0/lFKDeP
0ICa5atED4+X6Fmzp+aFrrXSAA71ToV5f+okl9IzxR/Qtq40nYkkFAmULCB33bz4295fIiFS0k+K
7nv5pncTYIWKirZQB7EBxD+e1Lw3ltPsZs2AWIVXesG2AwrrYl4FhuoEudkat7ljkYswwKX2GJqh
2JnMnBZiWd1lzE9BWhjBt2XT51u7tv4dxXAwDbMEIFUn4E76AFMWA5p2oU1IjmYCEHdEKkft4nZl
Cgr2VrSk8dTV1AwIc7U/pIhrZ/rdX6rOhXDLGPgqOUpRWibJX8qO2LhZhBWM/x/zYYOy/ZK+6SQL
nDrO9qliJVnbC9cK/N1j9JiozuVBwSmxynhjYEb++xGay8SWhbHhLRWSMJHHviouiM0LOH4Ojr06
zQYkiyx3C72Cvn3EVCrfBOhklGi59eSvXjaJyFQtpxXnDEs+NEFhRfKi5Au8/FZPXnaE6XCL2p95
Cexhhj1gUnxzsdRgz630sdOSHhIb54dUrNWHW2mfqREaVqNIlUMMowVeKWk6Tr8Fao9UjQKoEdkJ
fSgC0FN6IpYsSeD00UrDpQCV0vHwOdhkGN0zPLXr/11PC8vnBAEenxdSSQLKed1Spm4KchoJ1k2M
HTbozu/gAtqYKUk1DN+lRg6IlLCIeei05R2xo9zVvbDVo52xFcrJfWPHL2v9vGdc4oGS7r7K5PxP
eUFUAL1F4ApnWrxFLuvS69xLAT8nwcMTmxzRze0r98T88vm47S7RMSOcAKDTM3G8+mZovqW9vZZ0
gDtnoja2W+I2JpFtTLfO+eT9BPRaCqPH+XUisTjw7+bccTHMvGnanPTvFUOwSQnI92pV3fxjOZkT
dovzKJH+mEwab8iCrkcI3yo4v1sxuApIxLK2lA2CuZwvpuS4z0JstU6cB8HJUyHQdaX4FKIF1TDh
KozUSDLc7cpRD05BJK+80KPvuGUsTAtCtwd29T+iB2iXG6xo/IQBkvHLLrCYU9gPfc0ahgLfqLip
WsgrxnnpBh8CaCh7RYOvdU829dK3E+6cc7PS7k7fx9Tpfc5lbY8Bp5MOCkJPLRv2yoCgHyMIDjxc
pg//oBfRx9CvcjyaAeVLAHa8pzAXWs//JUgCCzZZ1U82suh5HRD0bG2MdFGbRbrskiirt9UkwhUN
31TslzIN4jO8NH83t6OEOKAy5aP1Qv8FRoZQgWFRZhZ70mTVHbgsaxfxPwjAbmG4gwrnyawQ/iki
c7msw/DNG/pyDIBS2v3jMr7u9WRQoQgfJaaKLL0pzkz8UfZAM/5/72drCjtr6uZ1UcJLfWLyWirm
cQL0Q+QbzLRPA7vFn2oforA/CscJhuhRJb3hVV51SKt/4Vd2uvAFBrUVvCbLCgVIlKycr+BlTom8
4a4jOYTJeSAvtQ25+NV1CW9gE+w1dcrhFVuozYz2m+uoy4Ge3WzHrpxS5y4NdgoOLblbD+PFqVtj
WfAEgh9LrER1Bj2oYitXjO3wYud9ERTV0QGvFJZ9JsaTAhMOVRCfixTV4uSznOd7tlN+PHRa98NT
FFpjjOq6sMtHzr+Bf57SiFHQhWQLGIioEG5SxjVZ7AhaWu2ZVyXR41jGeINK9bJl0lGM1DwxsEws
o6wMQxKZJAlN/jtpUwszH8mbu1DceC12I8rqi2qC4Ss0RLXJXkAL/8YLbOugzbC9i4NdoYO4tpvh
Jpe+CvoPIHW9dGwkXySYeauLu3E9ePyAmauxy9vP4qkKOCMu8z8aTZJVD5gVggCcSTaSnXsLuRhI
WAb1tXSZDcTUpkQCX82c9Uq6ejWzeY49Q5a2smqUf8mc0uZOKMEc+xA5tIhMPdibNVgsOiLxUKl3
HadTjGOtnx5DDBIm5+HmYPIn201XHoc7jcIPW59rii7g1h5xszhekqh78wFfoSZl1aCyYlXtV/G4
rO2hnJa+A4U3ZnfnIqmLqzVHnJ0x83UjcCOE3tj3IunGJuzMQGv5JU4S/Pj7eYbF5LLu4OvDIuAG
zT6Ks9Jk/NjToBaOVJTZ90yrSgqPsLRyRjEAOqOwy0q2AoFgj9OtuMAINLmMsGN8poLCO3Mhb9yQ
9PUo6cSHBTc+QIRNwofyBE8mMSilLLXFIy05nv2rGE2s8yYfVpV01rFNJi1DFegvqkmK7sQ2dket
cp66Tf2ycck/n858WgmNj3p18M+PYFqbofp2lRlpLSevCFPyu2QTteW9F2uH7b6fRcTMyt18PemZ
NFo8E06Yl/O6/PyD6XEhJ7mp/dZxaK2EAp6QyhrGVLyo3JDjBWv+p8c2khUMxkaD+oDrDOK4V30q
GfqKvc/mn0Tnzuqd+Vphni1AmFM1QNby6VFYXkuMwi48gPpOpuDoeB5+YQkXXEwwMUjLQnM9v431
AYStfPlvVLu2JvqPEmY48r+9YyRhstN1ApGBY/3g7buvZ9eV1VMRTqppDqZHkzM9bI/wJD7M/w1t
rwsQJZparXJQqxmFPmtwXlrwFB1cf0Ajg/ZYrxIuGtdDN1DEiQgvkcZG6meU6iZiAqVyt7fdoKfD
sBR50jm3aq8+uDF+0EjV/YG+OvHeI6afCpkTUZraRXbb/7zOc9laTG0eE1ra5GyRTMFxd+p2BGJB
bHohoIzVOukxxZHPwFLQKTbPF4F+PtOXbA+NS8W68FxBnfxGC0iHR6IjJOibbbLp+3VH0E2jqexb
pqUM/fQDLEERqMEyWE/UrtauiY3QCrD3B4BlwaTNTFBlzsXjEVWOwKeYlJJzj7NIU4IS5BX+awAT
Aa3WpAKnDjUXiCW6bhQpcBxMi9NAHNiEWjBqQTZaXsT3/zFpSmxLnFazhQv3edv4qHK2N2AZJ2Oe
Z3iSXosDVCghVXh8eF0oCAEQjGkO8n05lsvyOtrboA3oxSdPx6ADK6i3lcRVyJVQy2y13Ex/LgjH
o2wSw4PPHiiZgOCR2o/tmM38fzj5F5RTyJ75mJwVEUrL8ux5mQRCSU81D3+wkil2CLxDTS0+Y6to
VlGwuzt774RHDSpKMvRK1xhtjQlJWEhb1ONesQ4FxePKrZiXFl/qLMCDRdfSVQUJwLrZj+PVO00c
0omSUbrcYnSgE19CVqHtNmM8GTInsGKtopUC18CWp8lVWT/6GcdYFar5AL8i8WK3mz0YUZzwXYQ3
a16czmhXNR3kUVJnH1yr4ya03b3/KluBNHUgCK/TnpFGUdXof0yTTBXMyBeWVJp+a7hs7FHupi7r
CBwUfvnp1nq+QUKtloTWI15G5yi7vD83Qppta8GmUrxgdxiErNzMgzQpEFxtcCJYpBvvK/qa0z08
ptCgM8zaL4quEL+Q9B7XtwDTWYiuzkKohyPrFNWHfj6+/0vgwoI7t3wfdlscKBAoAfkc64fBsa7t
oDmapjC499Up39u+j3hB6GvqTw+Is88XO606tAutnFmYpac6xgKdy3HkBAvrxUoXVo+49/XWiVRW
wjCgfr12UIv6LZekdMgTddKd0Rx6lsNnK+ibzQNPvkWkKdxKDlS58gH11HW+PiccfplIdYDPhXmA
K331kF3G+1s/k8GWF/ntTFRvmDD3A/W/cvLEJlHQU0CKsoQ7pIdSQRMnwyAuVWfyEPAA12stm8wA
1/GOIF6Y1ii9MrRhNVG5TYZUduW2/WDPw33H6ka4XdrrUwqHr0Q6pS5cxEXUAlYoCwFLf/pm79lC
8sv6FKkTO1vDLMVjN4lDnK09AZpA7Te6I2KXsdVcxiNU4RMDmWHxmNAU4GEVJznUO9mK9aYMRBNp
WfWLfkg2Ql+2ZRy9XzqPrhdhKOq3oXkkIkCEWCRx+zvsCunewmvtl/YGtFXuV8qtxaBx8YKX6MhH
drF7c6yn4SORjIL/+cPf0gReN+2xX4BKrULDyRlGxspKwgGBQUDLjjT1y+ejYdSZpgMlET2gTyCa
3iTGP6Mw1V2dySS8ay58a9esxY3Vq8HwrcBk8IrRP2xtg5hsqUMGKtjHm6JqHTrZyAEye9GtWJH2
B7QgQP/VVwqJqscBdXyq0VbocYAT9Zwasifdb3AoBC5ZW9gd0pz+QTi2aY+R2MGma8k7EtaARUuC
qTpoVdE2MgGYOoOTjiaEPTsmuEziGdE7e47dGUHRg1Kjd0dSzoHtU72A9ql+a4yjeGV6RORiDuCk
FOwCX/QpxgL19WNKGr8DMMbTdfAQM0MOk70nsDmdr7BietdI0CygGexAU/Dl3YWISV0AKXbHTBgo
aU/3tWWoRciwF6kO1wQvEkUsX05Q/GdE376F/tCJydqZGGsWeemXFGNYZQS09dxo7NPnubX71eSz
cBIqvPJFcMsGjPsxMSbKpP4uTnyzBE7ImPSMcrKFqRSayzixmi7Aw04EoNgMu/vjjcQIjcvtdW7s
P4MSwyv+xTFucCRdKow1csycuFiwysqQJPm3F3vGclYez+x0szSoX9yjXs6Xmusg6RvFzPrUHETM
wF1ImygMX5STjlIv57JHOfDTg0wA5lA1A898SyHaNXMoZPMqlrbic/8GIkd96zjJaHIP126KODjf
bhe5nGDDqQnU4DpP40yXuykdfndxkCdcI+MOZ+YjwthjfMe1GRlrV+xZZ0phnZn79I/EkT0rWWKm
FsC6LcbX5iiY6G1G31F8ouhuyPqcu7wcsoeb+I8kKJAf7k8FCFGLahQQyfRfbM5bBQQ9x8JRuTt0
6vpgi6rJl33OIExkvmMqFi8bjVhWzJA14I/Fa1OkUWvffYZflK3EKUkQXb53e5HHwO8mxTKbXhjW
fdsgyeXW9vP5aHVuK1RFbDVlxiYnD9JkUJe7xwN7One7QDQIClYcNdHIrWi2HRTAPA6+exZKjRM1
f+jnVAgsx+mSZGYcQ4u41u5vnOa3RsfirmMNMc+L4lpxATsCjvfnjXmcnLG+YYPEDwzddBerm3Zl
taFX4oBkJ0ihxWUATiDlAV3rDbEb3Vi9ZXEUFDsR+fdFt00srWkZCuIYfiIsOHgaIqo8oPnNfix0
hFR7Ajti7uBRrv+zQB3k4yAjzWTqPLvHYRfLGLFx8p8AjDtHKah7mIVJBWh6qbjNoZ1WBLGInMH8
Se3zYWHfP216ENgvBIoX4Ltu1oHx1UOCDAh8Eqg8Cjx/Jucgl0ibV7fwZKQLpinVar0u63sS69A/
TL/Nw5XgNceKm/dveXxk2xw2kd/F5KZtJ8q81Tq48jP4twpF+LL2VURUfk/X43B/ZVmU3c8Iar4S
Z6FGxKGDEAvjzbIubTyJaOunrFfw59USiJFhPvskW9h3TRs5x3FtNy6h9z3URFOh0pxqRq+GH3Zw
8Cn9RGmXVAJYAgtpzm8O8u9vdPJ5u7EQuvYIRzqMxRjuqLIvza4Iih/JDgX07xVMe6Ad7I5f1o+x
84WJLv5mChqJPA/FwqGxxq/1UDZcLLoVXSRBu9H+9IMhWoYiG4JmU69deHcuAZOoqQzOriLLMDy7
9AWzKSeW5tdwi3bpREZTesrJ8xCqRkuzYM9bWuLUDK3MYbDPb7L5Tbhz0B2S+wnLk/qVbj1zgLh6
wEqPmi/veRiv0dW7yd/yGOAixjJR7IrIw49/QtE/WHzHDDjQ1HVfWZya26wrN662lkZiC5XG1pbs
wGHOkj1QtUMjs+gvHOAcULOorIWHVpBS9+ubkBSS/dvdJL57AYe5eqHeyFVtYP7fMQCf3mwHi7EB
Xi5/SlO786JiBGa+8v6XUjf3rrkYrS+QFragY87RYsXnhJGzzR/MTjHPntkfgb2fqr3+Dx3d5hyy
dlr5jSV8grnx6HZOD1ohL17V1A/yXAmO50Iq/T1w6Kd2QtJCcWf4H8g8t4q48Jwu2t0H8LtJfwpk
5/25Gj8kq4pMvdbpJDwN3YfcgnJihz18Z4VoavAABrD1zEU31PpjTM3c5d+kH5NdzHw7/Tv+KQme
/JL879fLgV5nk01sUh6JfwrQetSUMmabnijn0XJHrlWQCoodk1vK9kIRxPLF7tmcn6H9DnofKny/
BdA7W0VlJvuOCpt8woMkm8XJRu2b59LD8fuzK4ImFbJ8+U+Z0CUKCmZvDAII4wY5WhIS4VDLYRY2
9CuC+RUWlED4y7VWaVhHZc+4h3w4RIvUDVMgEcfvnPB6wFwnzYn4LOn/vjHBrEY7Rz//Bs8OWyD9
ckkgZVxTmOWyMG2x1ubd3dapasEqJ5baCIGMkO1di9UtpECdDZ37oPaj+SQSgHYhYEdDsROhIBg+
HlBzeEDZjak2viZbk9qEh0aUbAo4qB+346JBZ6kt6RHWBVdTeo0O+QDH2YpGG8/SAR+u1rcJ/n2A
/rqOEdLCzdJhTiVFjvp8MI/sf8GLJ38Llg7ITkLJpW2wWv4l4WFPNFWk4CJ2V9iQpt9llv8rZ/DK
v3Afc8Vefp09c3IT0Tghbk2g8uzX2SBgjhLPtd+oRpxGr2O6pGe3KeA1YcCSNrdgAFbiknUbO3Oj
Tatc6WhK/YYDQDC/yU+xaaqplzpt4FXMNKG6kPqeJFOPQ6sJd/X96haFBJuYrqySE3Wxq1NKwiJs
qd6HWLkbBA/ZvTNy/t3RXBamJSQLvR2TewJz7/z3lHQqxSMiE7QlRM10KsfnME/MCCqirHzvKwxT
B115NHxrIRn00xawGpiHUZIHoeppEQt/sN0MtTrRqp4rNDXzgiEBrhykdWj8ue3IfA8mvDAfl2Y5
x+QCJfo35s6X7Can/nhBvmy/EvSDXVLDVDU/tSWfMSibYPWLHLqNOFcHcP8o4pr0BFf93NYrBXHW
mqOIWG5egpKIqPcu1hsggHni9/yY5tfrJiHJAp8cKU0024XfA9i4md6hBW15r2FiWlzFyf9++fou
hOKSBVmXiJa/mhPzXY3WpV1cziuWzAfFJ4oyAnA3PsefGjXz5k5iBBCZlAfEMjWppi8GBReiUmGB
ag9flDtxmAM+kRbLlYxeRUKCQts3IrwkNw+5CkcpwC8tbzLoIDYxm7z6SKNgg5PCuhLSBsb2ffmQ
CdtSuwmCInqnAnNFKN7+EEn/YWX45ANbyKmF3lgYCpKGjKHfIEUwH1GSkrWE1BPjVPVQxdJ2H1MP
N8cMaE5MMtue4u5KaZw6P//cOzpXADrdR/0vPQmYYKF4rTXwz0nBe92sEh3vQ4LimPU5O84vvirW
TMHzy32ARot82BRpCaOuHS5HcRBxuey3r5HZr3zO6eTOd/5mYeVr18Ozi7oWPV4b+Ik37gQ+kbwh
5+vP/z/fjdlETGdWCzT4pxV3RWAeOtxW2kuoF9ukNRCiUNxLHg5e0GS6Hc75jN243htW2XzCk3zq
s0pumsxyRXgPuffKOAit/G+EAS7A8SzmwXwu025g12liilIkpNRfrvOWsBFHbb06izjbRrU8ZueV
ifmYIoB7Iu7k1r25j3kFvVTOM4HUZxftbSCWPKmZitABsA2ShtLub8ekPTFOt92m4kgWHVFsZiJH
TLPcvyz1tRqPIHNmRBIStK+2YcoNt/+2FwgNb3ZQrlRo4sgHC6Z1m/tbKWcMas4pZ3+j5EEi2OvE
BG57vJ/bNmWPtYCUGz+s/AZUggoLj5W2gxmKxQ0sRkKa1IwtDXRTY67UIEX2dnAdFATqqkSmSWxH
uGK7ZoRVBkvOFrcoD0hPvfwivpODDUXIltvCZRUOjeZ0gFaCg5cSLUADTMcWLXWEhIlNhBgEm54O
AuWhgnFK1Xq8yv9ZwA+xPYfTf43KKx+MYqazUhfkrrtWPT/nIEg8eTjsFD94tlL6VpTJRHskVmNN
VrlvlHoVXe4A/GyeugsUR4SB1C+7q+iisZoc06hLHrYhS/XiCuTlCXMg1Eu7iE+EuK3g1iTRDFG7
+gP7whsYnABvAcYvXnbM+HTWpXzSGZMZV4JY7QX2NPJDaoWCgKIMLlekbbredyzGfQcLxbmlxUH5
YULLwTni2JrpjH+Kqsl7V0CUUvMLlNX//1WpG2SAHR1f/FgQkj35qRSW7ZIRUVFCZpANYi26j6RN
ia6PrFTbq1TOUBAQJpVwCWzN0YCMhtDPHZkJaZxloTxh4Vy4opqwc3eRLi6NNTraDCktCLyyMHXs
nwwOcUeAB8p3gGjHerao88i5yt8WA74uuOI+buWbtH7Iw/Mry5+YyWQIDrGSigHq1o2DMaZ6NY4C
etO4Nfg/z/0nKmPvuF35M5x7f8fzb4OU1y+iySFhOg8vnUjJKDR/Ch3zcVULh67uvgT7JVOP97eK
eGXc0XJeTu90BL8QGq1wdXfPBg7krliP3fjnW5IkPEYtpf8W1HskJt3UG/KbJ5fLIsgGPuluB9VA
Ycy0AGReFP1TT4iu3y7Awi1PskkG0fOymEASUCsm466ft4vcYCRbRXwwHMi2kPmg0j5C/49rplY5
gM5zzgsJs8TXsAE00FLC4qne0XLqL6pgB1q8Uy80GsGSf1bB3yH0cGl7GtC6Zgm2NADJmYfr9sBM
qgm0w68aKrNIVkPCKw39nFKZFPYKOkK7fKDy0y3TkwagzEEZ9BCCUYd+2WeNRhwI0qovVgmL+u/P
LhMEax/tRSo9QUQ2BD2LvZP7sxZbPX/dl7VKk80YNGIhVBJ1xsEwalJMpzsp8IXxT6xVAzL7sYN1
jnBRsnokcpQ1z/wECQC5OCwOvJYf4eiPnY01x+HCzf/kVf8zJyhiCq0+UtY8WOVzXt/RP8wK0l0y
gmXKWut59hXRCA63VEiuNP5+1nL+tosxSIjD+1Kun/soPF7zIdScgMroG+Cuuoi+OxPYCaWSQUp4
427Y2s8EJn1t8de/7W5/yZCAxiLp4mnSIaffEJKREeSvi6j6DklVU0UqqpJjoRG/ZjWNw95jeOgS
xej4YsD2EJ7/zG0cQhpZ0SslegWgvMLDugAsFTnsGuDayDypRJyKrolZRXNXAFO6bBeNEj1K0OiW
DrK/BhA9/22yLIlk66wfUD/rybC+MAhbAP0NznLCNr0cWgFxdTXgkliPB5U2zV3G25JPleg7QUOy
AIOi+XbCdIpiHU10qjUOzay378N/4FrERAFB6PoB01XH8nvbQpxu3aYiTPtkPJkeglhzKC3tU9jk
ktbhBKr8VGlDWL1rM/q44YV7PtwAK31vrCGAdQvN9xqof9WbW9/sjjnqgvUEopPtir8UDlbxl+eV
xBF7rLfB/iLbqmKykYhiInaSOlLlePkhxXs7FtJCUwSG4ZQ8KR+bmrKL6DCkSYEchn/x+6OoAmpu
7UP7BDdHtRhR058heAWzTRaXsudR3T1ajSTxm/aqcI7SPdrHy1seTYcHy7U1a0DCf/6yl+0RTYHt
//7bz913MO3W5ntoDH+QRln13cS179OIyTttyHRwcK1+mgKnJEwk5od2H+lOgQ5IJQQVg+nAqXFu
okGGxIwag5IJszdbkTkUgm+cEgeQT9nT5UhgtF4OayyqkZVPXnwr/MzCiXMJG6hAkjXCYlY+zHFy
Qc5WuV/PYCAnE9nFRLq8puL40Nf3/gAKWYAhkvlvV9prRNDP3uezcqxO1vlWR41JSEdowV88ixLF
DQyG2IirEmpp9w2ACy1Yjb45xdsTzrmTxM9kcO6n90b2ys+pk8V7l9MHxsFIxmVUNBBDqNfypmZX
B+gUKkGSe4MnWaa+sxhWltI+ECSLej/pYhGTQD1kBkd9gFRMRwcFoWGYxd+YRtBdGfmfzkUegv7Z
QgG6WvKy6b0EVq3kQoZhRNIlVHsgziIkOV1AWwCLLUo6uvuYmWP80k/f4Vpf95tDerjOnKg/f5CJ
xjAJms7fWjaF3nj22YAeTTMqg6yS/iuqwl6Yw6OOMHZheGFsqwYbXQtGkWlD0vhJZFPhlVBvnjfV
UjetFNwfA+NbQNZEjtHOUKhNQpt+usjv/2PhYL9fvuM+7ipA+OMR0VtlchoYpnlWKCuPm3M658e+
tjowG+jIuA1GbdjXwPabxzM+N2tsQWy+MR0IyzdfpmEU7o+djSInRE4swjV+fT40C7sQfcuwpxiV
ibrVZGoADPvD5CVHZERDMxe0reoffkPfe+d/1ds9XhPgxNYdL5Lvc6ka3tfdZAWomoB9/pwtOrQP
iDvi31ebX7wyjKwANeAoZH+I1FvUU1LdlmlI4SnQEzENR4vLQZOJH3mzE8BmCF6NRPISclFISWMV
NEVseOJ3/ksK0Bp21CX64cWyXAR/a+0iM5Oc9Mmy3WHDmH8ZP2U0dXE4ZKymBL1Hjvki28xd7IyF
uedRD7noIIPTJ5fqHlBdV7lBJqcipU0U/EizhOr3HMQ78Fbe1LKz4zkF0Hc+nqTtuJhxKyzedTrN
w3czuiJ72k3DAAA9tRrUeu0V8dDRo/aZI1SWHJmTgUIOzNdTADdsPnKlydgwnmKEp0ueN64cPwXn
m0k8646ooOCHfO9rut82lVbi/YJYRRxjViy9PAiJWbAXYXtbe7DDmfQY+9DfCTorfM35v41SLqer
6cKD5yXpFq7gGmTfTnMM2cV9NJRNVSk4onaKE7zQ9v/ffBxstetRXruwowT6LAYaeP07lcleDFOU
Z28MXVMvCi6x9M4+6L/93SsVqqtjqw+jIqfW5A+nf3LUHGA6iuDvsY+vd44Xb3kDbp8Zu34C44rc
r4y2nVPxsZIVpvthhTqME/0HjhBtBpoFN3SlOeXAp3og9Wtp/3oDPNOJ2ZNHA/oq/PlyNA/oUG+D
KIeB5B+ykbyt1Ap5kdPLddA5b7gHmHNAU/s1TXcXxtuDdA4/wdV4d8ILOQNMaTYaQaXvXi1klM29
K0DJOAZlryQGMu8g22WZtFA9yAprDj+VxVl3L3jvvB3tnRQfOy942zblxqPaKj1sGF507s5owlK/
z2yrr29WztsRgUGGy9uK1XmfPQ5G/JW4VPIddw6sb30Vej/yNTWae1XfC0yog9O43w6vNlhjc4p1
ZmGPgFVp0szEN5Tw/anh+vJAc4uhHY+ok5eYOl5qdy64DsIL2ymz8GZ6Da7wq8csP4q0XEOKD/BK
P7wIQILPza7ZeHBm8I6IaVNkZxuBi4eEsmC1nihgK5dpH6FOdpPY8oXeHTNRJYqsjFucExE7CJKb
U7cz8QL71KUyCruoZPaZob8/8ORR6bbjzCXZ9l48CK0zQW3lMYv1wh9aLlLbZCL2/3xj9y9pTa+y
GucuFihd3Ed9tP14DHo0hSqJ+jFf/CtIbzhMef9cjQpPA1lzHLj0GTJCDRUn7kNPa65S7i2bLfD1
d5lG73BkMRC5s8yfx4vtNE+IFYUvNYr4aL7NaLSk8yOsyXnweMag4vucXQ52iP35KWmI0jKAiLO4
MnKsLwsflczz9gKsycVqya5GttslXnS6zyrYmms6h22dPLsUh56kY88xFZsY1ElAJn3ITUO40GA8
dgz9ycJ5dAaKIBf8l+Js31C1czc4+83BSSEGIGOArV/x/ndSwBsdNgm5aZyTmeFPdYohfUK9/h5J
mqNUKEND9UUI7/VFlvI7PbkeJuB568pApOqjojWn76B6Y8Tod5HLKepE/kuq30NI0VfkqiqKg5md
ffzvInY9PBAQenftZ/2bjrBnSaZQ/7RHQ/xn4yM8c1VvvL53Ll7RnsY35FJraSTAoOKGekegNC95
D/v8TchBqKrLq3hodkq1jY1h1dBtVby0JtSswzhfamLWsxnEyNQwFgPdl12wLtGBE+viJj0nnDA0
Yboc4l0l6O3aDKcpi5alZbqUhea3QJSXA3l35WwnNSoxayK3GcYUgfQLHfBStjKrjrBeIFigsPMv
6cO50BykCM+XNPtTK+yeabbmX94PNCfk7WPBgCeBi/w+DIL6nOp+FDRYcR8DndR7xZzaqLa1k5Pp
YsrlM5ljfjjyGW8lLaf00Me2X7EPA6xrUiyT1a5ep/KnocDHNXfG1cVpuem0DxD8mXIU/F4bFHPn
hiBqn3ysaqLCvB+pJJ6/bxs2urEzEx23OOwNGCjjGODIIOLvM+1dh0Yo6Jc5Qpvf7fg3o0uVNXOl
LvG2DABJLLx53yBb5G4OGxowxW1OYvzYewc+BPSOGX/I34qRdk4ibrOhKR3lFaxM05jGvU8OtqBk
i1ppct03epoHzaGUY+L8F0nlDx7ktVDaM8YaUbeB+iUlki2R1Nyy9XiDaAfqLES/KjXdEHGXA+rq
eoZHHEAm1ajtKtkXD2ZzZxYS2TI6ixLzCd2Dx/ZpkB/8xeo1dc5ZH7YiKckoy+ntgiIFI5dl24zv
QjAacvFbmJaW+SAqlEo5jdIfoLFA4AlENrYqFHf0oMW3yAFOuU+mVNWzdeiKx6QOA7PWPPil0ADH
oheLWJhY0z1E9JGf2VQIvdtlXDRH1UoHnCkebrEvhOSVeNeC9ejaAo1i+RvxR6DpXG2RTICbteyo
4WGW3xjSi9eCCRZUW9iwFl+64Jb2CNRUSE0ddRj7krD8XOWBnIN/gsS3lCLRvWlHjHb75Tmz43qN
P2yJtYrRI/DXJPm7ZQdcnfxQEMUWdnf1buDe34RJJXoGJqMQpMwWh+gdvN9KZeAK1jURY0RC01K3
QkLB0cCe1t4brYlNti/NYeJQzfttWNiuP7BsUZWNKS7U7WpMvfWfl8xFL4OzcUBEZJhmvhCqyeDj
SIHpDn97r7j+S3TDB/j8YRbSu9Pl2JkGB4Spj82SxvngtbkLrmEkUSzoLIWpyvxuG++Th441pFnL
B1mx/G8uOTl5MCW8KQCHlLRKXTW+bgdvv91cfw5C2akrJx/mw5B8yAEeFYEVz1Rzzj/StiLTnWbF
weEiAPPY01UmKU2wSM6+NmYXPpl/tIzw3b1r41a9NqCa5+GcgrKEIV3IS51YwqTcETCQy3lfT4uU
3f8oVcyMMAbeJ34jRgUZYtuJo1w84NqkAeh6sPA131HmxALcKORuvF2PSHWAxRVn5AsfZr5s+s0b
QJzucxctWXleBnyIwprvmhAe9Y+D/hIkZY+XMI9vDmJoeDCvAUjuvPDzu7aZ2tJ7KVQXCtmt4l3j
h1K4063nZ3E072+IDAX9u6D50WrwQQv5JbsScLqokUE6akgN+0MtuizWZbWLWi2R+ElP/3XhFmsf
Z/nSCTp0SmgWF7nrTxyFZklQaxw3X/5K+n1O+imG1fP02+ANcwPHF3PVA2XjSgV7pUhXY9xsTHnk
rD2MJSHlswhJ37VbuAFOsZQ7qibJmvPgJiNvRSBkp+XVLlOFlNcOrdWkfvVy039zw6l1UnKBbOWI
cYEr+dKgAF1VMnebDmxW6m3OFf2Qs+opcwwTtbfLkJlg4xu1rCV3Pi3RbbW9PJBnI3L5Cu8zG0yM
zNdSnHRfFgyHhVApH+4PIpkl7NEMFyivqObrcrULVRf4fbivN/sc8+x4rXYCTYnEKanisMqOClLW
hG2IQu9KKFnwnfZKS5j2jR8RSDc/1xK+Yk136AIn6QO1WB0FRU9P0n2HikWv8dUEeZVheLIgNWKc
aflCQMu0XQ8gia8Fzl/lBl5l8Q/FX6bKwN3/W4MdVKFkDjrT8Ipk/qQzBb+VhurONEzQN5DkPrIZ
WIMIVmIwGYyVsobgEHmNsDGLQxbum4j6bVIaMKK7GcbWA4tNI32YP37dA+57XNgvNsQP5ksUE576
RlkxH8W44ybiYezaggyaBK3/wBM0evRa+b4Wd3MdqPAg6sccOhEDGmJ/vcI8nrQELHIuywsAwMHX
O7XQXU4yxnEAr1mhPdeXi2cfJJOxDOQiGJcHQ4Qrr2+KAn01SIe1If7Eu6v1HdvGMPgqG+05OKwn
zi6kYtYwvTD+00+sDlJZgnQMlYnZs4/Kh4y4x0FJktM1Y3XEBg1yQcvvpuAhL7aSwxXWFJ8pYBdK
bzcbiFmALxzFeHuHnaadqYDNlEEIJpRmWnFmlL5qTIrh9SHP8qazg20tXScpZSXw07pFrb2CR/8V
dSg+gt/t+u9QTmO33/oymzZ5hRHDeS7bzSlCqejyp6erLyUCOab2NP9KQ80iRoCwMmLK94b1iltr
2o65W3F+JU9Sq1ly1rkyXHGSbmrM34a4jWq1UvZkpymcY0iQ0tlbA6nh+GLa54luC6v7lLrblxh8
g6ROewCRvlqIZfrmfrIrP7Xl5Emf3s3PP2PX6l/zvCQFINfMprGjbMDq9QUcelZ4XCrPn0Cgl3vZ
FWUWuRj+12fmasoBtAoQHvNtl13XRnyCGy+QxSNcpKT1ZlkxAJeuT/WbLbsyYVNChXJURBUOzZqq
RVcTG/i8/g5IH6E0VG8/jo7xBlRAMBcgpHHUqDkK0wpYcQc4hcle7zXal+PmPNwAgZmGAu85+OOv
Iy6vJlkaRjZKbqt2S+Eh4Qj4VEHXL+kgEXJxFVbSwvYLIkLkl7cUVNFQjC01WSGckpyNdxOvwnof
0FqOaq5SurN9Ow4Y7mC8bk+asy7EcgNasQAQMQLqHu6hyKSpnYFSQC9Ne3JLEIv4tYbwwwap4GTs
2oG6h9FeXvTuRsJ6KzOVgnF5mhiNZFazlRGXL06ls4mmruKymbIv3sMMZjzhBaG/kKQPHrR1Vdwh
uhLPCSeYTP0c9Es1Q6k4Vo+qd4C6utJbx9gn8FRqR8uAiIYOYc1ifljHvrYRw4MWvX90mAVR7UWT
nftU7ExtjzK3awD0fkMjW3epllnaLAtSlzHr0uIE97Lhq9lXhw9YZZm3IjbERgO71fhRRAQgjYXl
enpTt1FRRD63DkklPMz+QZ2VPZfYKG+hoCEFU8lV+Xkccyy3Xp4MhrwEk7Xp8ieRTVowbFcysg3s
7BPWSw4VUwsxE5mrus4Mt3oA6g5/L20xqQ3QjHEZRtbpm76/UGORNvyIPqero7qm5I8dSKi4BiFK
TS4Hw8PGgdX56QnBG2rVLRDwFt+Zyswt2hfsgqgRPMO/tOv8lWyM1BGGdQ3R7mzE0/ABdyG8aI3G
nn670l+FVBSb8o7Q9dP6PM8vW37za0OYdSKCJ1O4m+dx7UxzQWTod7RCS9Mt9WGtmiN3zI0bOgl5
bBdbv0AzppKda08xWiGF7byM5hKE4idtKTlInnIp7BXT8EFP61V08jKdFv6C47aQFleNFj6pZDu3
/ev4lHgaekrMobklljQQI42F8W5pb+loSczLpzrxupDzJ06A94E7rKgDPHcPeSxG+8a5ncz91t+Y
w4sOplG7C+kpRG7PNB8TuPFhdXG3/cvUhSK18wodDscfIGUGg2/vBdco+wOIEV2TBQm00mbtJjW8
zsJ9wwfpI1l6TkfT+giF5p3y64AAN3K4I0ukHqXbbuP4SEG79/THCy1D2zqCR9bXFhQ3+mbeufhR
O8YPIPfID9hW/6f/IBUgn17HiXS9G6SUQFOXGP8fLZ+Z10aNwqQM+jdVxqmdGlGpj/uMSnd1Sb3e
eXVi27qvS5TlVtB6SLhyU0GTWSX7OD0K299mPVrIRg6EohqKYzzNDxPEr7fh3URhyhVTItTReMvL
8eS1hB2JH9YtD8JKGUYq+japR8AFz/psu+ev6c328kC9oztBH0Ym1GxE9E4g1B5y6YxOWtPEtuFO
mELm4xx2CVklGWW6MMB8A6mPRso0pEj4KMksogY+67TZf2IM08dA9baz5xz/iYM0+JhXeJE+0V3S
ZsnHCCdc38efDUPB3SeoxdjRgqFKAmYd/bAzkxFMQMvqMJpSB8UgYd6lCg93DTsQMB0uWh/x9HaF
WIrfkG41atz7A30lgcCAC6c4gnGv/z9HYuR7niMlGI63T570TO5rP6NK29hCKq+cW12xkKPUBedl
AaWmz4EH/lASkPcTpPA+F+msIN/wqNm9qD4kTn+CPgiZntQLyoEBZmFkCAlhhBSpJO/Y0fAn8odn
+5uDtP9wOSZCo5+qkWFW1Z5m6yLQgPL7Vz50EgR0+JZLaoaB3ndbfpwhjF9KMdiIXPVH+Ay3rH/O
ib7T5U6JGyPP4fjt/Q0lXzVwPJv8nOTwEQvVlJGAHeNk7YxWBTXhrNlVwQ/8Hynuuv88RcDEz3ZH
3edCWF+IaGpcq94mP9KPpvMtt2e0TXgIiCVm8jc8l1clFw4A+W97IFp6Yyl1N81Jth5Jd2N6LZzD
kUFf9WWP9XUmh+nyh7jerQvOcNGn5lDkXL/tM7FYxCbZx6LU9gUAb9YatGVni4SzOg1XkMfStmVT
s+NBiZzYb8SdVKupiwhNsv4ssCgbnsb4cHBtaN6qXmB2cRHynE7wEL/TSnSjZuyqK+tqeaneKTmw
Y+A4ShT231ycmkDrFeE02nOCrTXaPRqGdhg3bKnTI2mhV33G3KoRAkxRhpZKqKHAtW4abpB59k0U
wAN1cW5rczf4NE8y23co+ma9L+dS2GvKQmhvP/v59wAVSNeGH1eNBMOBxEkXKblILraLmBFQcZQQ
uEI8y57k9XP0vLYJbVimqgaxPZFgdATONL6RLZR/M3sK2eeQUw0cM/9a+oIWBBADjpa9aaq0xZI3
HlJOGq6rrqSk2Uy3V1QfquqI/QorjngpjcLmZfnElIlqTfb7XvlT8DB+eqBz79gActW0tSLArUSu
hMLchq8X9c/VmV3UMHMEmr/R9ZhoZpSPhig7IyBDB/Gw0hhM6+I9ieg1bnvU0XIABlyGPUoJvngz
9cApiH0aJAuGt+vM+Uyy1wygaX5GzNBFdPm52dZl0w62CR6p1IF86xjjIJd2FEN/icbCTJBnzAr2
5KOZXoDY8m+rIQ9YWcJYSkH6ThfsVF4Xfis6Ooi8LMhcVsQQMOB3eRBqa4GxBVYnBly8nOq5HYF+
ktU7uKrt5umUV4NaPkDX4lDOhyIFhak6jFCkU64ONJoc+CWvzgWtHmuDO/VCj22igEA9RXu0aiPE
tVQRFREYTMbyFpwsakt5XoHJuOIeYrceQKuB78lN4J2XmtBglMHNz7kygau9rm2hTj/FZ9rOC1EN
wNTj1OYSnOiH/fI8sWwGOoSkoE1+EpNih7cIDQdEuKtEar2YI0BY+xrL2yzU/DMmNIomRHCV68PI
lzOwqyki+CoS/HNNQMnYuHNpKXaDAQmjfnbDnHpStTC1UnJaiCLPM4SawfG6PCMbh54ReTIkA09+
4hUK8bzAljbSSn0lbO6HTz6+TcKUU9orQUg1GtdS9I10Zo/LtpFUazp9bm6WrrtqZRKXCHb94xIL
L0zXEsca1bYBRAyPnU3EQtnQKjxdU4W3uM9JWFLCHeej1grVHhs71scHioIc5m2CJ0lH93WDYufa
TxY/1OB3UmxSOudUkEOfXMQ74SqzV0r4DSjs/uiTdBXqt4kKXYVFagErqj7xpuvb6s/GsORPuuLD
iHavbXY/50gfRF+66RPmd7HEXcIuv6Er5RrFbQqvaKbvqELVTe5+QZjjAuBC77wrwr77zL+biY+E
AIgZMjiRyqwf2F6ybWAmCyTM5kGp10oNj0h1YtMeiCT0o0gB1yzgwxUWnNCIqq3SoKhhfk8/TMSi
L+nQyRI+yPjKwhjRReuLr/RDfpjGV3Kqz5cq0U393NNyLHPPmZv8Qo9g3F3lyN07CVBt/2zr6FsT
8PAcieeEJRRkULpczizXCUxjrFLBYqtRa/3HarNTcjGi5uWf8MUeX0cVeloLHr/JDEpI8+PZWRQv
0DnPWRmcnCSFYJ8qC+iNM+BDDsv8lL3Y6USaYjzg/d7EJaBUYKjIx/3kPcfZfiINvRk5wD4Ys0aZ
VNU3/+Hg2IeHltY1Td2VNLTcKZDUO3faHcJ5l8tXIme+zzr0/tyn1nMUPquO8wmnMkO4/AP0iMw3
NW0YPKVFYf0sGlkp6yzBwT4Z8etToTEN+YTgC/8hrGULTwoK8LhajUx1JMO7PDP8zGxGQdzB1lYq
kO9Nko2cpsRT0ovIIhMGDAlCTA39faxxxXhWkG7yWKh2Qv9T3G/Egzxta8vK4uuTQgSDzFI5eYGl
kIIbobX3DKBp44kdoLma5uasexp+kowkquGnfZCVRMite+KZfy92zn3OmC1SoVoyeN34UeQHmm5+
doHG4euZI7AQtz9IB0pUQU0g9fjK45Y85558E8OyeqW9Xx4lqUObJg/yu4Ttg1VAvl2BnMHCnXXL
b9Cms4w0CFxVFfuWfeiAeHnlkv4as2M5FsJ+z4/2gjW1v6YM3Rlz9lWCBnQx6/nQL9tSa4VChrSD
4mul6tJ0wDVh3gntNMsk/yQK2W0JYvtX6dawngUvMVe7uZGCCA0k4AZR3l/IGB5mLGpL5VyrNGNY
eb2vtN7kUI+rVeoSAVoh6awqBk6/n1U8t5g+8QNmKWS572vn29kmkJeSBo84mrhqZXU6vo227ylz
HBz00x1g7HcIv3uRuO1K+cjADi8UZdPM+3YRf5y1u/04db2IrjU6xmWI33JJK9kIyncs0xXyq7nl
spF80ijXZI+ZHsmEMw/O9I0Af4wvY06D4GUSCj0eLaHjzCArHUTgQeQtLsjCa/n6s+8Eq4So/tBG
OxtzB+BOC08NRisHimrpG1rnQYDG1q05NTaKj8zQIM5dL8wXaR+SKOoXpJxPW4l1Os2R3pAEZKwV
+J004NByfgZML6zdtGQ6XLxtt1ilatLWqD4g/HurhbHM6y0nIgMVx2j8D5aA3ytfdiDZjwEQChOV
6nnP4raHUtDU+D81eWtw63M2DC1lQyrLwxuK/e9MjoyhNiHOe1A40OQc/Awe1Sc26cDph6+4W67A
ea1PELW63LHYAdnyRnqCkR7lX1b7gdP97OZzT/zpoxvBd0mHeZa07+LT6uWBu1+VO9isylMOhpzX
FiQrlvEToD5mA5IpTOCWtxrXk9s/fxvZjtVNZV/yAvg4lyCNPe9vN2usNbnD96cX3GaA1U5tMrAV
Mr31ycB9f4G6Hi9xgcmLjqYwcFY9GBlu19MCoV6WC8RaEDy2SRTR7u010RSuVHYI8lIx4kp1kjT3
hJ7PRmqpR3dDffBULkbnjF40TRV7D2VYLjRGw6kLVTmWVtDbH67d3YQaeIimhA5uEHHXSvi7brIb
eRdcxS0bFneydSbnv/v84CCK9yU6fbu1O9co9S6XSUOfxBOk9vBR66Mvx9zSG6RWBI4CVRrGqPAW
rFaSx2yZmEV3RlT0i9LHv47YasIhx/MfJ2x+6he1mnQxdw6xkcWZ1V//VAO3TmExELbz1zDv0LDi
4miCkstEfL6smpQVV8Vp7gCb3CBSub0LYowzzsCD31NiPn4pUIFiA5L3cWh56atRMEjVwTffDcLW
mkra5b3x+DQImhyBjrQwzzin5Y1qCOKi5IQTzwC7RlVjQwEma+t75xyeO5sbVEH6YLeMkwZTDKpJ
/M9IYbjI5X7QbutfjmvXKTR09URC9jtcmyErsAaWitE0+zncEjDMZ5yuSMLQ3if5PnxxLRkhAV1i
2z7JZGW780trgNvBMKOpCkUqYcunotzskkwhE7EWQOvv9mGvptMq57gUuCTKRWzyWW19PTbI4AqI
n1SL0IVlXA3Ij4HHZEGkkOr1DSJfbymHVAEkrGrP/IGdIvCCxZFRknJF6G6ncnA9zCNO8yzdXUrB
VUMeKXf0h3ztRGwE3LjBlEJyivG5Ac1/be3OcdH9WrTD7YOA77R5LtTCRBxrOxZKA6g52lH8txJM
1t4BnmLxeUbrzPDDc11ype/C3DfsLZi87EnXRPKyWZATXg0B+Igp98p6xSsvG5xx5+PRLNLSoPXF
1Zyvh6qwwfuVViP1o1xX0UIZTX3uDB+LKZ7TBJdqOewsC5gBJKu6tZBPM+iqW/3A4n/RxdHWVjZl
oxpVYaildoZ5Ln3WRlsJDSgfVZCpy9pcEPXV2fy1Eft6KSJLcbOOFclWNtlsghAoh+Gz1ZvcBiDa
3s19yK/CXim4EeJ03tubC2S4YrYJ9uSa7aSc/wcxD5iEA4uHU4F2Y9lOokSW8O/e/b/AtvKpEyqd
x/kSoze/wZYDRwsujyu+izybwdaOZIQltTEYbRujUcHNyjCJ8uo5Lh3um4ivjsH6Fkozd2jfJab2
6Syz22WDOcAXEOboTQeQyidBphVVr9+rPtW7cja7lJlQutBZQIAzuGxid914RCG/Jzb6HA6JdgdL
JNT08WpFC9fSWw3MktXuMpl4MnLJsHuqgmvSQ3JSIIk08xrz6LrcpLM4UOdD6aT2YVUM/fkMGJgj
KEumBGFehTS/mCsuZAdf8NVohqLyyhajqxqgTC8301xrUjuXNyeTjA8ocva5/Lvcxf8SoYmTTMXb
tVJYDfaFPN7iBwmFaOYKQ9gRLkH7grmGKSb5Fubd1lT2VswIuF/JX9gcNPavV1nKUiWGnEcAp6zP
AuENHiCtBGkON2vckjj7TQBSS3XcR8vPSQcHL5ac9dc+Mb01gF0LjsPyqg0ThO+5Rpn7UBGXLFOO
qtOJrzTNXwrUL5H3GQSC0oe0dLY36FWDTaiLvoYkD+oJKag5AUO9gjWzy8u0p7YTqWt4BdaeGaNc
moB0Rw/m9jq2DWf+6Ojyo0l1P0P5BHlFH5TbfFil+W3suElpegcYhufd4/3GvMs2noSIeQQYdF9x
Qy31kZ/Bptkdcx8MxcFV6kswr0b7Ct5nh2WA/L5PsEfrbUKLQfxS3CxvkSFgVs0p2qbOygd0ZtNq
Lx5BSrxcgYfFpL2a1W4r6e9WDz/7Zg7SGsBCkvPdN+mTb77mq8893fUDLSZucVzTpPGNsy91j/uN
K0o6rU8dFe/nRAb7OLTsdaS5PtjAek3+mtUCtArP1gLHBnCVzY3pmL1pXF+ptx/KbE5DuPt0ghH2
lrPQdZwBTfyR7sYEVFrTyq4FVbYeufRXacVv7Gsmgtzef/GiUezBRudlFpv6NU/juQaYEgmoykU/
iQH6ienFIbiDy1fZcoLvuTQOvTlgndk6CHLSPzBMYy9ullh17NkLVHqdAVtOTgYxOPfTCXt4L9zA
V0L6NKP1fglYHiakZCPdqtn9Ay2rFG/yTh9sBjM1eXOZvtHOs+ad70SjgE/Uovst9trc0HtIGJPE
Ir16BThtkSM3L5R5J/vdFIz8jVQxYBgtgWwN8xx6PHgLClNzjCwxfTkYLkFJFf5+1QnaYMhD6Dhd
aDDerwKqK6+i2TxLqLYkW7dOVr/wtF22PO9IcgRD4NuKEgmZVVYNPO5s1qcBoPQCsVS7uklmt/b4
HSpjCCvK2bJQKBEtncEbRnpDdVMdrXgggB5gv+RZNHviRNgGqYKp9RhzrmW7riKx5cYujH/fHhtZ
XclutfOT99N5tXHqX9BVW7T2Cszzykkp5LnV9C2hKTfr3iJzL3q2xZateNK3jOFoGYGLzVXbySIV
9EhYcoGHaz78e0+vtVDX3dJFEFq2pymaRX+VpA8ph74P8VuMf1QPnfew4YnX5UhLlvDZxXYv7uaY
lioUO88Hn5TYZ1w+yD5mT/m8yoa49IkMTH2p3HKtdRMizU23PQ8DQCFymAjs/J3C8u9C1f1T+JG5
N5Iy7fQBu44y8UcjeWWAVq4jBIK+puF/SGMxqXTs8yteJzsK48NROuweovIG9+MWvSHwNyKXDDTe
fKyS99YvUH5MnbXdeXhfmoX/x3RnRI/6kdJX/DO0mVkuGFtoD+txPJVb+0LNL+3UZCeX8VgkXFRY
v578oVfqrQgpVMNC5FgkGVa4eTMm3q9f5uwfm3gBvpDFpUUtV99rF2XugitpDc0qdty17t5gXI9/
QUcEttGuday38hvawXkmqc5dVi+8ujLBjShNov+iclxhKwgFRT6fMOMJzZN2IwdJRk2cCrNNGkkr
YLys3uPldaXMkuAkP3R8up2Angb+ysWiaBqGtx1K55EGB8pKijPT1gNhQoivacQDYwpI9ZxWpt0t
s6y8XSdlyrse9XRnL0MF8HsAYLbSdZTDfrX8plCWK4kt6pePgmx33A30UIK0NvCyNrSN0WghEtTM
BbfRDD8YOBoSq7fUBA2Q979GSz9yEC5qjx9kldcinB92L//5R5YgNYDYBou3Go4BYDhySdV3C2l8
9u7qe5qr6MmD4ykLH9kajh9eYUr+etDdunDGTannz1dSaAfGJCs7N8VyvsqzcOHXyn+sEvqaPGAW
JU519s9TDDmBMkO/iixycuF1uq696L0NPE84iygUvnJr0sTRRGqw+qzJqxVsmWLFOcJ9qZw4YBD2
qRkpXaj/ltMlODih9ufNNCFZFH1P9aKNqSNf29bwzhDxRRIi46w63rgjMa/a5GAbCIK2cHcu82Pp
IM5MUHzS6QzTzplXJ5b+/47RhrmNUNg8jLTWS5Z76LTZrXhJPmvDS7EJ/HoEVzprtWEhIdgyxBH0
5nDnu23ueHJNAx9wIYym6Hy+nhAkDEBG25vK9eRu47vGhebtArJPTghJNhErIgtfUfnHxtHY05dU
dzHJF0+MRN7fFPLfYb8JKTdf726s0llruLnl4t/ZrFQ4i/CB2C/9NU6goU3hAVPkfBYeOFo6h8vJ
/b5D+3nOWXMs0mHm0QWCWpi5iUH1Yfi34ZH6mPs0JDETqglwuTEgnjOaazEiyzn3SBhEuBd8qPCp
BU590Z4GX0Ar1AkL8h4r8ga6umeK3gQ40hIamrbxcTsmPQwM9ERyRlwBI0uLlZal6C+62fej71RY
5oGvrIXb+W9EeXzjE7qYNPVFkDY6cg6vm0iO30nrEW6MGq9phs+G2+uXBOqtfVdq+ufgXYv1U339
6hS5rQxd4xendKLQBFSDLWMoBWNVCt8NCbdAZa9szcI3A1vtDykKBjQ6PigSTqzjH6f43Q7IwEB+
032am0JG4ynNyZugiiyXXNccdUEvbiX+fd9m5M18+bgooQKYaKYll8h4j2YPQrmojQU2yZt2Yg9q
GRi01F0j034+YLHOavv73J5jNXRYLuOcapLTK98+I3CkrnOZf4UAo1mxYU7DOKrXp/LkCRQkY9qP
a/yXLWPrrOq6hFZZBZI60tAXuUQwBrr+xOXGF69mp0MJ/gEgEGV8M8EN/BoTB9iYJKspU05MOrUF
S1pPafRQtj8WSv4yAiazWJGW6DrfSmQDp1Pt+20goI1CLBKKylWUmX0FH6a6tVfCXoVnlvRZm5Qi
vNAzHChB5mpPbeUcOK3ybXuWLMsJWoqR12iYpQqF9CXZP8eyqrdLEuW7R9YjRRF3pRTaDs3BkSes
8lfD6VaPxeT2ViTnEvns0NXyYqAS/e3q8X0vDYn6zMI9Qf0KAQyrM6rqkYk4L1XZwMjUWWGAlk5m
Eqo7UhW6tt/cN6gUM2QT4BPPw4Re3mtoywy/7eaddJIxvc4o3JQ0Hx88WXswBUEJUHX7wl7vnClr
RHrcJw9ZgUYnia43G04BKvSC3TyJsteb2//RRnHIJ6QPEbeEtmk9orSlwu18AAgvHMUofPhLLJSx
YVvoZA4ffO/AVCLov18dUFHtib46bgnFmPsIWSTXxx37eAWIOx+OAKeAzLUCTMcftQUvHeaNeqi/
bLrej/Y/eLeQ05LYciMOIQEt26tp6HPg6tIMFUKwg7eNuK42CRlqHny8s12L4VKA2aKompqRq1/i
SUObqpSOTrXBBCtIbn9AaZ9N97n4sOb8FWHV/QdIBXMspvB5hY+89uoBsUwT2qyyVxcyLOwIetIB
57+YlHFbajFasxC8CReHKT88EIj4amAd8f/4JFRGN9q7V0ftdt1o4JSHJ6Hv6HKdKW6bfGy0XHAf
I0fytMqOHFAq3Y42tVFItRbmqVrqHGb/etDbRESapFLRvGyr1J12+K9kpAKtUdMZsSGDT1R9D78z
GxWcJlwUrSGApc1+A7x72+VFWyWb4e0GrCg94uk9yBfJdsSK7mjHZ+iN/FMx09PsItoZLFyEZROl
uv0O9snkyyXo6uy5JuiBfF4kznF9JCjjTiSgJUYWh41bp80ZIXa7lCOYqqdvk3P05jhFgcYHbwsR
3LSISKQaNsaVq9A4La60dFNFkXHsx7dQuZrQc3xXZnHF/5dx882vc4V7xJ2b04WYhi5Gj7c2lmA1
6kyWMbdBLUeDQJ4COx/2dYgheloN5UqeAi1cBDWJpIcdwS4XTr2fOGUuPVSVO5gDUa0nCPwclREo
+cMa4VijjJLJHz3dJUFcjFoK0S4P4yoh2M97Lzs2tvPwYNQE7RY9iTpEoFFrlSiKkHUDtTeQKaNu
1572VWBsU+7YuWD1/WdXtPkmCmL/dXbi8zsnii3EgYkCYO1NfO/V+8Xh687YwAOeHSwre6WijjqP
8c0ai1No8PaSeYxFyftz4B3zKyAFlbCcc7lIXRtHqf5X/Dtk7495utZG2gfsPrl42/Ovjt3kH8ML
76uTRfF/PcQdOSk9wMZaON2Cnsd8p3OC6mOZjAeyNJxs3X1Z3sniJxCpaZnNX8KCZNyDQWYn6yO5
LpG003wmt7iEN4Cezo0jQyCyDkxUDDaj7yzJQ+md6LnTmRUwcKi/SKVE05gKfSlbxNQlcWTb734z
eoyq7x0487MnJ9C2l6g4uD1pvl5Wn+8FBZ1ITd2VQ/JGyKq8KQypD5VmL2XSapjV7q7W/2OrB6YA
G4yZK2ZKyt66sWP4SorSxLcn91sG0unRiUNDySutWaidj2sOnZvfzNXuhkev3yeZPCIjIJw3Ontv
gzMSmetLGv8TtiKZ4/HTIGFiAkMnsqxKv+ZG/BDm57W+3iTpgMRAmDMumP1P685S+6pi3rl5etgd
0ml5KAD6KOY8Ztwa/euM1p+DQovz3NclTfGu9bYT/plFQ/hrs9qcKRtOU50j15MRUjgbFL0P3yo+
JiYHtwFyZshnvAe15X0iQzmF0Mh2YtkBO7T6k0RCSt+HmAy07AuDKj/3ke1X85xB+ILaz7RvK9ap
BDZdPW6SmXcn1Fo89rX73rIdTZHgQoav5TZCEOBEIWiZrfpgQyzDrmcsoYclENpxG9uGcFA5PIx6
ahP4reXLTeAB37RKzrdInGbS+pKAlfYEYnsY6crNR9XNQ19KodVwTfphscvJ7KsFFYc84Cql8YL6
4BiZFxVU+4+qTFIxpnCRVz24Q/Gybr/xs11M+D6vsHzkckBvbuk0XcN1SHWLosXKzkpm8kDLJ+zm
ovhls2DyPHFplNkj9+wSyHrzNbVXtxb4ZJuXyr9lUgToh4sD9J2kPsL15FxHv4QyL9jUPJTCGy59
sz/SFbEDuVU04ws1UlF1Q/tAIuRfGn0FLOmtZpWgHhPRzrCeqIfat+/5V29xBRqyIKv9MUWXtY+t
dhMsQtQH1y5gJFXXDFhXdHgQovHUrhvvPTZOVDIYpHykKk5nhCmZST3+F4/k9avPDQB9zOwaMg3y
RlunijZEaeNFos0olKfm+Jd1LHoMkU7Hizx+Ak0Jozw7a17kmTf3UH3dA/n/2WYq/Y3UUa7EsNlb
WWr3O45Gl6D8rdCGg0cUOsRdw1vK20GLuna91HGQTKXRsLVY+YZkfjjKcwuk4nYu9GX9DnA9x//Z
D3Hs80AbhGgkD51hHgnCx+33jAWipuPFvpRmrbvlWTVEkWhar4Wh9CeSAQrSKqo/eUzqQ0GDKibm
A7bIwnrkfbT+YKNHPVjppH7KAh6jPFVf/eOEWxjvQlnS2CcVf95CiQEcmakXkyLPEDVn46aag22h
2Tgk0qVEg20X8J8XUyCiyYopWSmZdHlYGYJfzyGRzZ2g7Q3zTXmtsC3qwG9w/+d2FxstA9sN4XVg
Si39J47jHE/fQ/ywBYhCMuKdNMObzu5K22E1Szl6Mma2t/IDRv1eElq3E4WlhEKSLPrHi2bIUmh7
0rZ/4EWesvViJdrvM1W5Su8mzNWR+kCYlZ1EZv48l28odQda4fvg8e8AlQ1pmcXW5t0VpySvUczB
mdbSnJ+3W9hvtrCbg1ir08Ui9PT8zIIGIH0ldmZGowDxUVXMVjg7DbD66xW8KojcyXc1s3ElKKsL
tjRPxPYMI+RXHnbGr+GJ7SdO1zRv81nv0dsMCaSqVrLg2WDBRN1uzpjCgx3KNwYMECit7KNcr+zT
P+5kEOPsj3vx6o0J+KOIXwzUBdgnGvjnoRlJyOdZ8r1y1w4/OeYSjNBRz9KC79jIkKu4vu6dUTW3
xYfBN4xmm41VFlxEwWI5Gu/9GwwVfb8PCSwRLsRkpEKkxpXuiG1gmOuiMcCPjn2X9RcPxLOSW1lh
LtjBeQVLiGES+Co8VAjipuKpF6G347clAZNt56IWvjPvSY6ODWvFqN4ANcJnUWPKb/N5EIg4BXi+
Ft/IE5w/zFMnwY+qRn0wUithCQ9HXCpKQv37qZcS8dnpEZb/H++B2ZJvxS+vaTaiVsEu1KdClbRk
1H3GSi9/YOA17VX1pTwMwrTmlnofgLTr3+je0VwgWEiEVTbaOi07r1p0Q/wIJkwPDCdkfCF+nE0H
tfHSE7kd9ZNaC/V/eWCZTbLYutXkkzPJFBpMaT9t8DQg6ETpXRN9Zqe6yQ8s6azI2/eMYAassLGL
6vcu8BK0ti5aqcEuaQW5Dn80tS6R3rb6uB4xO7kGDDNuXjHnwXAhy2SrckICuBhublKh/2R8d8Kf
139yKZj97aH8q9W17ewMOwMDPhQbW70iRI26AszgHsBEJZRo9ETqvm1Nt/fbMXbFBocvYlGausdB
AiUsRFXTZn+IeOZ6QB4NDKuQCDnYvWkbKoBJR8m9uEVS2ApnivnIUk+14XGVjzZZrkzbNGigzAi7
S9CjVPwcnm4UYQFjRg02WaU74EjGz+CjBaxWILg129mc45fylTyjR+ZZJ43y7Ho+b2QP3zLq912w
r/yzyw4m6wz27P9SPiBUcmy1dWzxmqn7tiLQShay4Xu88N4CnPlDugzxfD/kaxJePWnnD/L+bG2m
bdlTztG4ahW7s59piV0IGYzvqmxd4YIRV0yLEY+7UXxXGLIGTtUy6MjXctXcbYhYj+Cq7MDltX+c
p0CRrShkknuaXHhm+/CFEyQ1QgjTHIEO5QQDrstnjMhdAp0DVvhyeq8jmVPlRMr5jpog+LYQnUxh
E8AWA3QZl+MK388r9QloikL5v1bDsA1npTze58OiyPpRh+sNnfAnHdI/h/ECcGvMHhANhrw92jIv
RMEPqT6dhbJTf3jHTZ5HXP5gQADSy4UIOnJu5iuSui+EBv+cTQonjW4qM/xivmNhDWVvKOCVUS//
49+e+pEZt1KUixlCCUbRk1fp0r37Frb3s07ptQneKV1zb2VElzFsHg8NhVYJEbAveV1P2uqjMvT/
fXtWtjNmk82v/6WXJWJTlXPezGHA42v8565kHZnYoL4k+QwY0y7JT+9iCskaan2CUu/g5MoBCWN6
vhmYfrb3Xqp/ZdrkqQa0t364BW8cUzFP1HvtJDJZ90uHDa8zZPHMZ23mJeEpOVQ5gXxsU0d38mI0
oxWey9g9GnnLZmKc9EyizkX3Ug+yKTA60EYQnduW4UxdPyRu9vmw1aNoy988yFptwiP98xe+cM/4
VRiKduMNSu/FlP6il98ZfK4Xc0AdRPb3PsDUUZ+836tBAWirPGKOOrzDsMyRpRqzigaaG7Dpj6+c
h/4J3dfcb++cgsB2bDhhn0HbK6rKKkTXqAMjQuoG+wd4wVuR3ZdNKMq4HprOaPF137sRaEIfSo3a
yyj3GWJ4O2jaybtwtOYe6ptqECtnyKlm2WwrclOrB0JH8BLDOioFomCFChWGYup0p/o7xJgyc/qp
gU43TmupjMgdocNNgc0voAzMQGuPd7+Py4EqWXLvTU+ijmVtVAbqDb4bXoOUyufg1H1P4LnYVa17
znQRH2kqwla/HhHXsCjYS+vdw6DTKqgZ/YXSWnHDY0D1nwRfNpE+RFEdLJXkGmFc+K6aN8w3Lsoi
5VtnOlnYqsHTyG9zSuZ9RGgqzZgdeEdjbz0x7Q7fe8DsaPPE2Hi/FE7rNMT5T1vtccpIVL0kMn4W
ZMUDKtQ5KlSlHbHR/6BRZNY/9Is+VRnNf3nTlX8bucccdGxIrfQQ9vPQ3Mxwjq3tg5o9o7OOR169
fQl+LQGoX5gRJU+tkx/1XQPxoze0n9e3oNVIAyyiQMHrwfkvfD7JUpeHEEO5DTmHiks9t6GDXfaB
BkmSRIl6OB/YgjjN2gQy3wZ7IeGoklj2ig+ZFA/qOg56+6CLLrOmqaFDW8o4zrrtO3SPSth2jIoS
240ph6sNawoptOkwuu8AwdqzRbsZjzVj/jF7OFR+MWrLVFztZOL9SI3XF74xQDuqt3QZh8GghOhp
RecCH6ZwP94KBlpKaXipfbW/eJp3QTTJJ7WK6aUb0utsvcB28rsSvt9YVRE16Xw/2W7P0EZqsDg2
+7JLj7n+2OVrfZiwaynBUtuX5zABrg+wXku0jMMIA6hJKjdW4eymWnNXqOoq/r+ekgiNVcvNlOmX
5FXId8C9dCOZoppKe5GLeHP/HLxUsJ0H6B3F9oazC+V8QXZsz6wFX5ZqzTAHNTQCQ8QTErB8SCxk
u5mNqDefODyny0GtmdUOiyhyjz8aOi4NuOv6OnF6t24KZGpD6Ld9mmu4XHvfOLuT/oFeAh2jMUUm
s8uMJ0YwiElVDx/nduwfJ5w+9GsRXbbt1tLy/aVXUuQpEWNigcbzGu+UFKr4e0XHXIBmKurfxWs0
soC5zCIfc6WLTc+Ll07C5TlnmpgRdteENJtID6jqKp7OvVAkW+FseXySmvVQXkSYnN7lMJ/b+OQO
xk/ddIK7KieX7+QpjbmumS45wLfCog8pvpSnN7/yB0ihVdBXfCDOl5VWQnvfuHkaaJxUAdx/BNW2
NtLBRQpaswgEtKHxb0JAIQ7ms8q7oFk6RnAofirYL2Oeq4m8L4n7VAEAEOcbC4GvEKZ5JXbiQvie
PNGFB4aTXHB/8iMDumELjXNxph2GKjL6J/WtGLZRRu48oOiwpR8eLwxXHF82LIzWxo+3Fg3Lh8OQ
dg5w5Hg0rzbolE8O3GQhHvHUdEmGf3JfegEuVK5DRkN2VMLQ7H/is5I0YihtUferZFm0fnHMOFqV
x9bs/1arpyNZbacsz+cLK+OBwO32gK6VJ1gWCjfLNFZS3IUXFUUIzNgOP3oOWQParZQpH4RuQNt3
TkqGwR+jeMmq6b2v65EpxRJfYMOM4WhZe3I7GC9U89Bczs6wgcXvbp8payEiuNt7EembfffVP42o
R0qDeucIeTRGM+e6kF3Gy5m1QWm6KrWmTJ5W4WXsJhfsEBHJVguKKRqZvL+85LOvzk+FCrfuKrHd
M42npTBho0VGNRN6iZG6NKbjoecwWkTOcODkxfOUkAUlfZvVzJ6myvAWXCGLHUQVgojaQCGluVJw
7yL3jps2PEeUw3VpPh6OQ6TqYRnlODWiNSWIRcuSaTYHNUKo9QUYil05BwrdL02/zwQXn9cn79Lv
77nV7MV5fv3W8XVKrNcwFGnjtshxCdwIuYBNwYUL5dZ6BDTDpYTeAgjpKCFX9eXDU1s7gJrEqhuW
sL48Zu5NeC+Pa3nkiA0EpXYJsD4+w2MSZKXKKnBZ11HWE/t67nuLsPVb/UfYZLqITAoIO3qb+OFF
Fz2gCYt427TKj7iFC+I9EkkQj6mPOVkn9rL3Mcat1JHe6TeE+xd+hUdNlb+RkpwSDGi4x44xbxgf
aOXmf597eENaDRnnScgmzLClalO/jIiZmf8DWI62OYCp5dSCYyYZtC8F4DL1+N0XXLwUIGyvY1Lf
kD43j+gph4w5z8O5e02rOnS6hb6puH6fEQxd+tyNHCI5e4NLXdxz8ouUYMsHRlp38ML1ipu/4zxX
e/Gxae6pisVJBh2HjEd+3HrlSc3lfO+d0pGkgg83AG+IiJSFTyor+Xr/xOM6SCOq7zjO6QWeOziu
hdVZftxCo987uHBqrhSi0lhYKL2/l5IvG8JKoe9u0Z/rs9zhRjV9IacG9bU+Ot++LidXbPzQTFPW
9YM7a8zCNcFxEFe8BVzyID5IEQ+s6hswRI/RyEfutZBEy8uJa8A5sMZ8qriGPgk2HO9JdvuThxO+
XVQqgaHn8Icf+K0e3xah1tryFkXu+KqLygEKWTyFq8y7KPlmSqZmFJdmSeSsiL4GUXmlT/4F0BU/
YblRMBCIWMli4PuEmMvb16a8W6klWjUbcIgbGWNOt6fdxrVIpI42WXA9v7e+Us5HW4TYV4MIi0Iw
QVQJd4klgvPSh2n5CNc5X9M1rEHuXFEAr2wsUplNS+o4FwqPTqU/S1dwx6UMbxEHw5de368bv5P1
7D6h5H1VLOzZvSHpstCRlGRtbKZE7nXRKpAlWD2XU+5LFeHxZZBeiPDGk3hZL5tZrKOD7/YfAcWb
/fBBzzU3pBJUf3g4gTVmNShBW0DpX8cGelQZE0NlUEbsDrxdo8DcbgSQVnQU6nGZ8/Bo6u/MAh4f
m1kBuszw8ueIY3pi/27bnggw/5PejDk5XjdMPizZsF0W7PGxFgGBydmLUaMpDhbQcJuTvlsPKrGq
Pg/qzkWlLIOkaV9oZ+HI3l5cNTFsI9edkXPmPrKUO8gTi8TuhJdt59fpPMBMCAOu6GAGYdxkB+n4
5PLuF3LLKEV1e63+DqUJnlnUiael6RZzUPFQzKRHDRkQ6LldRtGr8L3UBuFAgdyMnF05sbv4xkBl
19Q8KIzsRz4QoWQN9mrnGLbpxSm8KTDVKaMlip5EvAjmAOvsbFaNNZ6huf6Nlz8T7PcR84056oEd
uW0mg5DDZX1DOeeK9Sb1CvP86R3wnnHm0xHZCWWD66PhaHeD3ra9dWTbS8LEJ3w+OJmVWM5lB0VP
HyfOp8/DIr4Tp/6bvmcUa8EelHDoWMPWtleQNk3DNIDDZK5mVWRxracTj5Ti/+8nrST7ME+naQ1Z
NDeNhmiKvnWodlpSsqKt1tUXY61q49SWGanj+9vzj7wxB0Z6pEeCMUQez6nWoJztnwzE6DYW+1mT
rjvT5wOtn2l1/K0yfmBGFJLdQ7+00AokJO0f0C34oc5fgMeJ62stJoQM2kFiwMeH9dAYKudOO6L+
yrtvDx4eff8PuWseCl1iNhjGQPbHMxHQnWr3gGeKCE+zPlgmw6vjVAQZSj94kLsjYudw6MCS77IQ
Dy3bwyNv5w8qDwSHrnXqKgSe1ueF4H2D7z+FeSCoVJwpjvbZ8EfIKuF8SvxWBPx+LH4L54o9fk/2
6Rw8XLOOAfFGyFaRVrok/As/CR1BDvv833nlhX4dnHbCivAh7ste9oEBITXmozFulKy9IYtpON44
EX9NQ3VRFCIIZcGPrGVvIY5oK82wdCf3DL5rcWkDr98am0hjRZI0Zhx+hZ/EQcC8S0IeQJwdmLBr
AbDRelX08yxKppAS4eqE1mxuztli4LAVH6wYNzVufxMznutkPtyaY1WKYnOc0d8i8By7VUSR4/qx
frlq1QtAzncQMBm+fBcDKPtwU4Rj93DLp3/jf2Qun+r+KLLwEgV5PMPMRJJMEzg62Wh4fbjV82TI
Ox5B8eZVsJom9WsBZDBxK94aP+ok6FYwWSxD8BB/aF8dwuIG58RwOJcAhTghmnAcjvrGCFguWi0O
AbpQ5Ado/2JkLlh+kXMXArvdJNGE/aIPvz3P8qMAIO8dRrfRCHHvadnEUXOsUfwA2zosGejoVQ9D
clnxAIKG5EQxFE7E5gVQobOSC/3eFtPN9ydix3t9aMRDgvaHmvKgR6yixmewHoaie9B0wYjmjcpe
cH8G0zTcnQ7Z+hAkO30pkIiFMZp7z6iyAgBnJfrAbeYC1gxUyDQtS4YbeUn2KXtqSPE8ioqN4fQD
aKcMOdnmYV6M3GwTloGNTjAN24Z3ZzwiicmdIcZZwu8CGcd+DgKhTxigFZ5VKLVFKFyPdluChWdt
PiZLAt441rowTIxDJVDfbgP6rs82OpRogLjSYgsXKM256J73QqOu7T97CWAzqoKTXyV4Gn331MA3
TN6hJsORXdfZ5IhAg7N+j7B53c2ACJ0qYfSMXLEKvS4gwHr7fKGHBVeOFzdzHNJgSI4/+SX/MZwA
WGCbinplos2wvnWeZgIy9w5yRfKlLAOoQ3RZOel3w1HgoeURwt1wCcbrLABrZJf15zv+UcAnuxcf
QZP5h+e+I/2JPLTM0Zwrcx++MYT9lc8GJXeTlznKTUIoyfrznJaxFnd0+eteFZSbWLhuqW9bSDiU
oLp2gcdfKXeEW9xthyDn4CKFw4+CicIr6pDbacX3+qe8KAcnZuZRPa1dZ0HhEZZohhMJjPHyMdEN
a8U2yQwmco/TzD8GPHGWNRbq73mO4YnqXv26wEaAFDme1kx5wrOh42TUTVrEixslXsE+PthRZ8OU
Gm9crl6Hd8ySthJJsWBqJ1XOGZJz2xT737CbXsTXOumzyQ07bXNX9GbqYenDaFzrDa9STd6dU1HQ
mXVOsqd2aHA3GP7f8H/sHzpaCKjg0Bv1SUiTdL4IlCtYAEHPd8KXUbZRFKgvDwZmvAVIMQ1SgCbA
0HjEzx7+gU5HiwLNZXIG+YrKnQ2KE5KOmcqbP3n9EKZ6cprNAvVnK1vIFVBtuptGoZxzxd0LVsUN
t2gLb8JDkIWy7nrD1w6nQfLCCcPniCP7ka4ia7cZL4wm0/uNVDFgx4FP6szsk295zBxJAnEqbB9m
VPNj/Gb5lyfdiwMZYGWadG5ZixYH5VCzEghBPguxIJEgKzsM6ywRgv/+1yZ6e5BiT1xNQp4C2oPc
3IMMjxj6Uj73PWv/zechAgj2rXn7s6ieZ95HGJC4uV6g406ru0strj+kHLm+pOaIUnlz2wCpkl4U
AC42JMrILGN0zLjb0DaVZkl8cFSI3uAxnAFq4p1+i8KHt7U01U6lgP/JAa5+s+FTBOYvb/m76DbI
yhL5ufxwn/rlpuld8sgzKmAa3wjMr0C8hT9IynNhW6xN16p/NEYk6YD6BaVl9FZIgG9KsY3nl1Qm
tifJp36c+ZD4HU3FQROiccgnD5iMWawK/3rP0+tQ7NBQz3S2LMX8sNsxk3Tyj+TRxk4FPJB64UQl
cuAfB0OHGkL9UVhG5F0y0VPxlx5InP8kexih69AyklbRyJYn0D2QnDaqYrQ8HzVR3780HUEcx/Jq
8F/0mKdIbQrboz+8eNBtfKSeL8nHQe0W7hSbLnJBm4QtsCXZXZAA/jAq9xtnvg0kXqMXj4zvJlT0
fG6uISpOpzm4I872s3dFEVtKj6dghQsvumiFi4TLE7Wb12ltMIKCt90Jg6iobpUVorbgUzhH1nUA
xHErdn4ijQmlKW+Ax+H9D7VfIj1hF90SqRXpcyWymRcJYbBMmCFNbqxwKCYMuJIeJsIjxmkpJWpP
tBWfscsOI9C4Ta/kHSJcJGE/Q5MI0KJQ+PVm8qiogci2k93jix0bMfhrhXFEnqN64Ysxe+Xw4pxd
H519wcGsBcwCFL+vv0RukBdN+Hhvud62ZHermj1v5sxW8Kfa9AWj+hZ1zjRGTRziYNxnQw9XxAgW
iqf0xw3qAGizvu+VgYtsH6ETrn/fRb+bN79P3woLfrRSwesajUXj4Jz5lKWcvP7Jg7r2PABCbEGG
OTA1yHZ5/OvlrKHrYFtRPtWUuhVMJ2sE++b/bA2hTOtSMSd7Gg4KdJt3BfDoMposgcedpwz2G5sX
vQ2dpKVWavOHCKdavQr5TQ5Fhtl0Vnx01dSnab5oOqYfmVKK8oy7kVU2x+K5NSn5SCRpExo6HhYN
D86o4VieJogEoErpu5xNOULphPYWZQ4a7Kx2tIRTUB+cjXiMnWEOU1Jtkgaca4g2buUiXquUpvoM
jWNuV0SR88mu2yuIBiCBo2/Kc2VuaPE+q7YA0OxwXTlFp9+AAaoiYlWHr0BMKYsredUwKXFORJQ4
N5XtIHheeXldH0yqaoLgx5SocNGjXKDCzLq+1vNwETg/NL7f1dOBgWW81poHKVSc8Gv9u2vceC5R
XlJcAsu1h8Vn+S1nMkI2Ei2aktX3Sevl3mFqvXxOR51jvrvdXQF2L3i703oHZSp1HHUvx3Mdssce
O1CoLqqfzH1W5tnxGdKm3j1zm9WTemcDHTIERbjdFmPP4Fs4WENNfn46mm3k/gYobcWAdbxlwo62
6KArtWgonKtlKAY5yjqTjk1kSCec0d/K8TFkVwnR0M+vKhVCxoyn+cE7ogbTfFJQkyHz4ViZOjni
qDbb1tEel9ANScsHmgqgL/BhsmoJmaDS5g0u4bsWF29qRYTgn+K6+YI6j+UxViv1aC70843/WR+T
+02Yh1WyB8Bus9GyKIr2mlleNCD6LtrfUa3GP5FndZLEEYzkGFMOC7Ha1wxH9uGkchuYFKHeFGip
rZZMe8444U9+s/wvcxeNPavt6b3mf4EM7v2P+BVj0XUSPuaRWUTGoiaMKZ7wx8dbCo2+uAMwwLZe
0XwOWYIqckiVA4JAxI8aXvTnV7PvenHmBBd7Bj6FXOK+scbTh4IrWyhgZVm8nvJJaMYieSHy+L+Q
fZXd/FiuWFGF7OLu65QX87wlb5oK9pntU/juanvex0JP4wAu18Gzt8KfU87WWS8KN/LXU2T0JB2F
yh+tcP4W1hLPL/8TX3oTUyfWL9vV028DfiIhxKfURnAUtWld2NRCDYFytRYTJkdQmWx1dnh+jhy1
J1ktvd1oJhK7rQVHVa3lTjuIenbYUjzRaRAytirJ8Km0p3+/kr7LODLG14JcXxPX72tdQ771+og0
S/SHZtpteSWe1YeEivfefjvAtLUXOiOrsqd6FGgh8gXY3IQ42MblJoqDUz6W2gojZTKt4MIGqVEZ
1ZcyAB2M1gYzjG0IHdemSaF2tijvjN/qfgN1Cw3W9qx2tEydsDiYWYRYZ3+3RQT7gNlB4zm2a41m
quriXCPza4PGQrtO5WzMrlPp0/D9QTufUmDc313uFIbH9btKlbkLyHNO+0mYxGxI+txSr9UT7abL
F1paqGlHOzpFnIpQ9ffEnqlnoIJz98NEWxBIgGtpCCcfsJCyeLlvg/JkoacI6dr1Lm2jnKfcFD8S
X0qVwgjvdOv7HH4zu3dFv+ZD79Hw5uu1SzsiyurDkdXIsMJMH1Q0woiRiXKfdP4gS0r/yf3pAHK3
fMqXoqHByG3TOKpYdmLtmOQHJgFphWMbT72PQlHZbZrYDJE62eyyrTrLZyg9NNgxJ1UkFABXZSCh
hk6xcQBA5eN0Tb/aIdz5d7BEvc9ob2VPS0PnZmRZ8sKlOSIbvcEkHCn7QySlFMaKGpHe75p0e/wu
tVUoQTP5lYtkx7jXpRvCqG/jfkyzIacrOAqHiJI4tW8xedyTjqSHA3fiuR2FX8a+B/PLPj0VAv+G
VWjb4oyXvnV5EVrzAFp2R3GmjCKLOW7zAo+Qxnp4KHaFJ1/CMhCf/UDxEaPNYPEui6KL6kF2R9Ka
XqTkBfjPfZ+DRDWleNWSfB6A7OEPefcV1Li+OBRj/gnaen2cStuEt68IaQBMgwEEppkIPii4HPZ7
Qagy37oQbPtJ7UoUUKn/nTt/9f+psABMVKVmjME8EERdElm4yLCqUh0K2dVr0Pbay/v1h7D/szDj
YjTxrg464Q9CCsygRiSYPMznSsRjnCt/afkKzfa4KOh6GdHbYjYeQAchfyw4I8NPGPAbeYt8Dtvy
vHlpCFmRLT2f3d8oi8NFJTBMVUXhfk48SKXeVNt4UXD+xIdNWakNtnn8CxpkoPNHwc1Sz3klqS5W
bD2gvoa7DujFmfe+TwQIL+pkAwj7s3AK5NAQ6e07I3VgfWSHFFg2UVMpCTCznynOQbKV6SelhMs3
2bNe7i7AnDDZt7A0Y8Wg34HKZ8nVJbblgg54FhxIkxmhJaKbXxsSbE+sMBvyQsrk3jjHx8siN+eL
rPSLLrhLTYEUr7mcBuczQWYV55IpTzoSiIPqUEcTdx1EQyUtq8IsKLsZmqIPpC1uWhu1OeHTZjnY
a7oGGv+hMEdvibr+mTxBiK0z+kgj5KtB+qGhu5s7KXXZCw2VtrDZdAF07LJSUVxzUTX473BWxtjX
emT2Qj87Jxd5X+TZ/0caElHYyYLwLqMEGp0mZulFYh36QM4dTGYhhE75TCauZAGOj+ZXWdJmvnTl
NSM3njECqL9K+k8OEqcahkdOQGeYm5U1o8oHtRyokGAjg8BJQVPhjC1Nr8X34Sc0pbpyUeqLs9r8
n5vgOtqxzB/DCatTrvSHcf223rYd6b/jZO6sWLuOOH2fk4W2y7wGic7TfN19olx1LjctYWERCbTV
cTA/YOBeqvpECW8b3dUurZTPzc0qo0kwV55ICbFl3vLO4cYe2jDULz4caz1UiKHOnDhVw8G2F5sV
nBJumwY5GG/fNlb7J1KwmfW1GhOck1/Bb7sZXAlHWe91THmcIHz4IrCyUgJ/T3308ZifzM+rhFCk
F0MDn3ICSn/w6jS6bWg9Rcfg9ISw41biHOoJHApbnjvfs9Nl+X9QeC0QbYbERJ2Y3226V96NHFRB
yGQqAZqDap9+E2xpoXe+PGLmJpUzT3cBZkEwgSe8a46oKuaAl952vPmu5Ob1nNe9ACopF2FYcojE
Zq4vMglhtPyD9OZ32E1b36CZorsPH9BQh5Zq0/KI+RLavHARQQP+zJ64R95Gy89KzXAkeI5EDVX6
T4mOvxSS5QcPpu+YMRHSiwellyETI54oE/bMsghFqLfo40Y1ff0ZNWUeme9BTegJKpyf61ZBqAeQ
8SmRPFYTU4J8oT0AJk9jWJ+hUteuRe+BLXKua8Vl9RtJ3T3lOYcecqUhOXfDBHp69LljL9rW+bGi
pxmZttjXX2LqepF09ft5GYYriAzwnnRQm48HfaPxgPS9FyJ93hRhXCfJ/tL3UKIFOxVAO1CYiuc4
AsHHofVAvbPqi03OlLqJeZJFiDKVfWz3PYgmxvc7bZ3pzSZ474sURRo1CxyXwPcDxiLu2mxx8kxO
kzu9goY8rdzEJeuQskXQrorrOkdtY1SNmRvbiKiYHPTa2A42OU9YqQz5icBNWtSCK571u0G33IVq
cCJkkcEvyj7d8lvLZfYWRFEF7NCqKG9m9YO2UAbP7eskx0GdQE7yeGM/YO16Y+kIPVtKf9SebZTs
p8QOoRfakOtARJspvwd676fmUW0oXvrr3dDwOoAv46YN1qSfoVSaKlUqdJNjSWcRcNw2poe94Wk3
ARtlviXaLSIkUY45TlcmPLOnxDazrsAm1kcHRkxAZOPvjouLVx+0L0w3PqMbE4lEBF8P7fUU6dlT
Kx9vfekA5XdzDWwYCwzkmDinSd9KUlm9CJ+lQkX7CXZCsQMym1uIOjrHvlbzOVL6wW4Afce6qBsV
zmpm07mqT32A4bkn04h+371tdJudWdUFWVzJP7VGJnHuZN7tOPiE9m/AKwBm+IKBvE3RQ/O6Axk5
pIdaqXb71q6XgYWPcdVwHRuSzQb3E/AVj0wLUAneJDNzAA+OiZFB6FiAxHX5zu43r3EPQuoAhqBW
629gIUovm/oYH2GV+oLuM+T3ZMEL4T83ra82o/JIvvjUqHj/kyOiU4JIJd56UBJN/hzCqwjHFIaf
2mi+YHepXbMDQm/unJFh0k+p27voQieaY9yiamsLkIU2JCcpH0NtIIVuJPm+lmBXRE7+c9MwhSQe
t2kruFL2NoKvoQiOwMjpXHTu7tFUDT7NgFRuO8THxvhIsUXHYGQNJEN2Dw3LIMW50eX17m+b3Igo
2VHf+6dpOx40Z4tFAuv7KZd9dxgf1BckFhOVUZXseeO2jsnok1b463FJO4gjCAELkbcwo0dGCo9R
xehYmURDXRfzHUCSb7zU0LLvwHhONjiaxudbh/D3VVCdlFuq5mpl73msQ+kpTgCLgmoPd7qqmoGd
/3FeJh7nnhVmCnxO/q2L/xFtwz8TOQXJSYodoo/21YcKNEmX6ePLdZ/47Yv+umqT6FiNe9uYE2bl
nnu4rJP8r31hLL2Dhsp8meQTt7uNU9LPoyRPo9QGk7vMGC50FInnbou4ZECSa7hStlQqFFALQIoC
ZEEyiFc566KqZnw/u0VTe58hDbRnbh5jGMqu2UMcvTy/11hwglQwsHHKKbGmjsGUwxgUrJT2xEwa
I9c8ra1X76Kcb28yDTzjplXu5c/Iks8lOZELaian+fRMiT4GksUjJukw88oaNrR8BbVKLdAl8oZA
+weuNDhS6TuEYS6cifbeSnFEqlijuMsdvvXvCi4ZlKLzKCQa2gZvAP4Bj8iViZGFpJq2FgjDh1Uq
kcshMM0aQJJ0Oe5X49z3JVJmaLG2B5t+3Hl/6l5Gn76q7raVYTPkqJDLmfUjRpUnP4GPrUuPNN+l
qpqFGX/Z4GMZI/IZryGX7gIJxtzSsV6LL2eLN2msWTs6cJWZG0iABP+qyYqmOI6oNEHVDk30yZrD
wFSa+U4NTlb0kDwNVlyRbi0B9t+5k7CO0cE3nP2p12G5V1di+l6ISYEw1c4ZZmwKFDWRkGdsSGeR
Sh8hE64yZHyhWqYoqLny5HyL5n637I7dh1F3SNlYP67U5kV/FAf411Wg+6t6hHGEuCW8v2qvbCP+
Y1W4KWLCOPk9KPPel5RJfQTVeisV0zLTZB0ZHQBTZG//os13wx1+2/v/CrNTSYgNuj62+IFbnvZZ
VnND7nybyna2sslj3kMGoGs5B/wwE7aTpAHXJ5qm2N2lRSxQcTJpe36OFFg63mgptaKuo3YMkUKn
d8qgDzETobDTRWsDMCVYyUV2EMAQ37orB5EAA21esZlGocMb73Tdsolho6M2wild7UU0ymiQUPIT
meY1hTUhpaqxh1RclJ1aR/byEoiN4soMpZ7IdKdYmp6gSXgWh8MVzsUOBEyTiNnJOCAFW9rXmcu/
4yzlLfTv5bBYG6sqnEjibxN99++kKA5CaCrLeYtdyxBhPrxpOjxSZJfmAFfe+HHXyU8eThFd2pJB
KsLaqH4TLilBp9zWwIJJSeSEIa1jFGShf+SIYNik00gaKI0uBj9O/TcX0B4KYQVPOB+Acq4ysOzX
cZ3GY0JMtUd3M7JIzASCH3Fqjtd0svpOF4HLNuMlWX2usZB87UW2zGeLMoZcnxl5WZdQ6s3N6iUX
gwf6sVDcT2VS8QnUjti0nhjwI6HLZnCLo93Ko5ZCQqHs85EmMpNbpmEMI2oyFWlg7Nb2K47qR7p6
l90AoZ4cZUOlDmT9MwCiZ0Dya+J27R7cXycFT3T0HSkw/vDHGYaaBa4GO/cjkXtx1RHVvxZE71Bk
Sj5Fv6lfFR44kvG9uA6fUbJt3NqL9qSci6dBI8xUpvIAQDFqmn1tQ+PA32K2FVZe5OKy6cz+8ng7
BQZJlCMTiaOUDOuKzSqpATwRlQuIDa+r3oyD6QSw7JhBIkmaSSSh0f/vXgIjJM1Hfng8YKgCNuox
3Y/Hjr/0nifz8ipdbrodkZSSQl85JR2uXJT1y19gActsyroLM4hoGkTT0NinC2r3WD67m6DjKAvo
kB1qW4Q0FQx9FvVCTqqtAEy237bOSMFEyIoCQ2hjRiULOxx6GKPhZwjLIF2cHJzBVc7mf8L+NOqA
4sNHk1/jRgiZB/Pmf9Cfq7qCt/Ak6Rh6INv9AO1vgakcVu4Tk0SSJhLGA8w+ivZZg7U/+MZFPUY3
7H+2u/Sl+IAMK0UUsLzPCJM7LvXTfRXt0Hp8iZi3auPBA340LLL99NFpkoWAiK8ZhF82L/dwMvBF
pNMBQBjZy7UjIggTwh6orL/7jvfatZ8C3tKxIr1DF/LrbGGZbVF1xf6XrGzWU4jMUIDflBaQoDZH
QRkAVkS9TqVgBxGRk6AKggihABESs1YHDub8D36ctYO+JBSS4NkS5jgub7nQfV6zcN5+mQ5zomcB
6vtXDrMSXhfh4eyaBFSTygKwkgPgOw265gS2u2z9S43R3OvPoSWjK296jNn1fPn3R0iFHNyM6laT
3E9GsHhwCsO85N3FNl/eO31lE0oTW5c0ye23LKfpQm+tF4sz0AJt6sXNZua4P9VD8yWww6cavWtF
h4z81dJIrezHX06vh+B1F6AaVPpngaSINw4VXoHkvMMQFLkqgyEPWVmXkT8id6Gy1HW62vHWJfts
lvMNcE7cX7GUtULVFW9C7NgBWlyKduYYFsUPI6sV/teB9rS9iCMOUM0PKB0l4n7kwWLzkOWmwWhB
6K+/jAdic9+bSLzUurZp5ZKkEups1xREpB6Y7EIuADltD/j8MIafm08jxYkwwZLfw/d6PMrCknpn
J0kbrpp34W+EeOvP6M5VS2NMe2x0kW9zZxIe8Y92bcr0AKeLRPOjwNLKAUm1QTIOWrPAHfb8H4dH
lOHGZZe/6q4yDxvrnogaBITdczHZUMSwnPFimUE6xwqA04CBOL30xzoUytDvuTLuvWWZ2qHbelDC
hIisUD4VLXq5Sh2KPQEUQGuzs4xTTTFbu8H6oF/AA6y1HJg2czu7Aas6ws3PabJN7VRntroDvd5Z
4LxhZU8j6whXa77u+K2mNZuzvceQ4fjXvHBzIqAHFq2OHi5I5wDeOZYl8TVbuZMskHasOn0Rw/IW
+lhDc5O6zcHb9u79eCoSIkEdlyCUo7HLeGsBai7K1fgfp6OgJCIZi/zTxX9/4533R8eL0AWr4P7S
b1gOQjDvekISkGx60s+H4V7J1gnQoq3GQ9q5EeE3HosaFja1zNv0yDht2p1LjqEEEkvFzIjZlv4J
ma/Aul7roidTvSk0p/L9MWNI8UWGJ1Ru9pA+Ey0YYSMP1eGZnqhAaC3YFjJKUKrcWxDZxWYsHA36
+xHqofhRXZeYoea70r+sQDWJpxKj8djhTEDFWM/0F1Z81SY3XVGlrlqJDamOZkz01F2gyaOrh9rF
5bbBUzj7Ul1/48liFbepE1jbr6NjsbhCnLTdsaVamk2sj0N0zPQIqZ2lpYqfQRVlbAYVKPqWlDgQ
HK9vltGlnIsXkUpjAmRj1L219PQn6iXLN68PItHNpOqccvyu6ZkF0UX6NzOCRWXVkbIgF9OaHzeN
54MM8ckWa5xPnjondaaeHbLQt3ys8U145hsEaQwNUNNpendoHBuVkoXAexQSPUIPop88SwJfaV/L
AlWfWkIvgHvdQfvmL64HM/VzMR7O2jd8947A5SawjGI5iaQ5ui2CAOWCopBQGgsY0EmscOXOd5pH
jB0/8FlFtk3t4ibqIC1FbsWvfCeCsyHfEG/XIXASMdEbMLhcLQHedFyAl9qk/upLQshjnPbIYKqp
8qlx6PEBUUTVTsxI2A2Ghq0yBgxxydL2TNhI5gUTdTAnVnoHXkxtWQ81xuQz4RC2W7E1SvjBLrfh
QPX3jbJPRDbzNrXSOGfs/Oq2HyjP+aX/uJxnRRwHGaHZN9CqBpdyWLfcUgkrLnQhj4RMqY29r75h
vvJczC7EoWIEB3Uva4sV0+fR26IEXb+p4uVK2WJv9YEDESoy4YWYW5LZcPvJfWR5qCBpXFF25+n2
r630KqFnBKmMYv8zwQ133N29//vb5fv4X4a1aBr6uCQBGiUJd0De/GQTivFlYJ2KBgWcDjmtD9hD
ArYLQN5tOUe2/Q+8nIYKn+ysU3MFTci/TAi7g/9vytaDC2ayzPMg/v3xieqHEJAQNxmmw0vewtfd
kNvSuHUEQWjpBFuih4Sg2XuPgcy/U1a9UpKt9MubRYOIC058RWzM6Sp+NcoMruqs1y6FsiWTH6Dk
dQEs8ZlM90t9Q3/CUhpUVUuanxNxYluDsdLmUPch4Y7hA2hrLrcyTZ+nwMJvvL+8/KZIVkY5Skza
Chp01QP/WS8O4h6J/vNXEctArQcYMeTqlJcB4xiB7JeV1R1YDph/lWePJedlEVbU2NZ1GDz7Zswm
4RUwofrtrdtuXnYOASo1sPa5EwnMKHQrO60jnn/CyB8s3hJPmJbL81NX95977BpJq+qABqaBwDqt
hzpWAfuYj16VY5NxVfYkZBMrnw9OIi804BpJTSZDhRJ95Vrfv5MGobIIzlWurBs67Q5yHMMvga7r
I+ZqpefA7raCLciTXSyFR1LzNPlO8xLIE8J+oShYEA/o5PA+PP/zwEPNn0UAcxH7eP5dIdLtkPUK
7KN7uXQUe29CxRHcv2lL77ihZRpiPKgBPVUE4Bn1bNDCWSKnZhdLDTMnzmuVJj0sBPQD+uMhZy+7
IRAZvOIRXpcJYIQTg1b/Sz8eAh16yANGXAOC/2IQ1vNHty15H6GViVkoyTHlvmk/qk9vTtvdb2Nm
sZzGxgJxrErodhYivPsF5U2shxDrAa8Q+0X81BnN13L4A/msjlBKBheNrT+kM49AQhpA2ZBemKo7
79j8U7w6W1c1VEoow+m2nIQ45psllwDVdmj7zgf/o/vICqlUs4u/jRG3IsWMhmb6zrBLwH2lFhDR
TjtEVrOZYJulEXjVdvs9RkzXQV52srUJ3YA6i9zj+AZISkT8k0l4ZvkWR1c/jdpa2s57JanW4/Fd
66GByfINoDJm27LdAbalZZCInVrWt3wQ7OTTilPHDL9ur5pu3Kv0GZAhB4fMTl5ULGr+ZySkiNc0
OLOWC++GwMd1g+kiMgm/65QsOQ6MWTCS8RJ9QfgTLtgd4ykFE7nt08sJJZyBV5TWhLmF6y6RqF+L
Q8mBHJASyMCqIp8sRGIJ+QdNH1V4pdfZbCHcInQuBpLbSlRR6q91MIeKGU7b7UwkraIIk52Pwprz
AP9OvVYpTHbezIp4rf7WGYmN39WvNQdCWF0mhzODz3dNrGsE5dwER1wb+jCA5Wp1alTEQHHy/aHl
WL7YUFnEK+sdwoilCxzh0hNpL8LBgdGFEMRXkS5vtR446nvgqOg5sUwHSG4Un2ZigKd2YCqF+4bR
fB+wYbG8w/edOG46TXeeL9gZ7k9JhasZ7wEBQKLnhTDMEqJA9XICeT9PClus/xftPGN3Hu5CkF9R
vt3VtvRwQOKyfF6dt5PVvty58EJnkBzCtkJYtiycd7cNlyRrZQ+o012b1s4vbEXSTKznohO+S34L
HM9ZtORoRxzFlNWbgP5mmXZ250s7k/cMJxtI2qZjWE4aoxDMUIf7r5DZQRi8levfIVIwLcEFzHtN
K58cjGqtV/qfmRDmVdGkVmDtYSujHho+8vrDCsU6GtaBmv/cHlwClzMm/BpJ01y3PNpDlE/stYMV
4/KJCKLFEawM/wXVgQiZeXzDoEUuZzf/KJ/RgEBemf5OIgtQMx9WwVEtypURI1Mbu96OhOOYQJIl
IkOwcw3CNV/KZ091MeMmDjXICW3GKhoh+tQpJzvD4xJqCMFGf0T6EWEpOTMTjJdbY8hAiDcJxTQk
T5x1q1xfoFkpPt1tByCkRSa9J6HHfgEEbCC/9iu0fv9VOOi4WfcynZP9yOfw8S1pEpM6Qyy2PX/S
m6+jN55UDKGXAkYPCtCw1vyV5b3PWjHs/t7mE2hCgSamq6tZara2SiSfnufvv1bpT1GCNs9T6ZXR
TUR86151XgHJMMg00kTWCB3S7r1NqJ1XX1CcOzTdRia7AjNGeGyAHy4aHayJO03jALwi9UUu0hvs
LU2wbblUFjhWIyA3lT60UuMxDjUv6Hex3HHsuSSiuSRYM/52+3e6T1Ou5OduKuCsh1XzFVEGcKQg
bRwNAiAo1yf/mYl8BFJy1OtFvu+toOZHf+LP3qQy+rv0wwywuzuR96ndI0o5jM5tx2GMp65MWELO
Cm/Q+yT5PzlGH7W98A/EGnm86VRu0c7ul0E86yNzFaDlYfjcsz2519YJ9f7Xtjsu7k/mYYRH2t9/
Qa1apdzTkXrrrtJUjehEUlJsoFVIBhBft4pvSA4UsvEEtvQaYkyZYTtYpErLSSCxFpVLUdylyfiY
IzQlpVDEmZoCX6+pZKfn0kejlD+UHdjMUzfkCBlL1xUwSRh8aDgq7c+2PC47A6NGe7bF0fMlSVAS
KncFsiv9I9Nw69b1amLIIpdOCJ+E8iyvRv2c8hjSGD9k3nlQQHj7hj/KwaY3jQ83ij1aQaM5va+b
O8UCOKb1U3v0emdfAWzWm42wp4B2e7Ym7khctcxmOsTuI9QHSMqA5EJwESJOgt4+tlnvfP/KSt7/
HXJ1kzvhdhbgqhG3qUFUNMG02kN5SK1o9AiPJhDh/E1a+tFfw7O4tB8b8kFIhmo5oHLkyLEu9lIY
D/SNol+prdzj49+TIJuJAsTHmF+jznEVumdxiWMnoeYZBXUHOPZKs8hUTzo3zNdKWUnSR92OnhQc
C2FceV9e8u2aL2T5FRjODNcBEuN6PjZeCOPBx7KLPKAscgozZsH9z8coMQ2zgRAvfKOITtO5SVfW
eAabIuz/RUSiiI4camJvkb8fJU+ZGgFi3oXcNs7ZZXPYkNry4CiA0lLXh1dJHcCB2b+ktwCLs309
Hwj9C9/nKBDF7vURp7eYFeoB6B93XmVyeL/cmqb29yaGBVAViFsGyoo3Ydna0vYSgaLE+7H1aCnk
D00H2Vxzb3Lxak+kHUp9UdxKvV6zw4vWRM4fNtDse8GWudljNM5HudTpbChgegsElALMYiQp9j1t
akv5fOoYEjxByxk0jh75TWsA8EUcJQEFRs15I2eS6jhkLF6a4t8xWOX34HJ04AzPniE5lRstj1jW
8Rv1xoEkNzOROJhh1Thx3hKxR4k5BWv4N4hWPE9CBokkt/X8XJsiII8tyrzzB3dfy7bydU8rFA9d
PgHd0ArzRNTZnnHTjqjEUIwX9/koTJ42M31kRuugN7AJXdZKg1ObDTM+coXxYL3k9O2mcw/CYmlz
F1NOQUNW12p2ijto9oVGWg8Wv3Elv2kSs7fIfqLv3Vw1ohK8fSxXOJ9epDxyXTsTAzuRp0j4lytw
kDMryKeQDpv2q9EtFMKWrfKCwa3a7z87nhJmYWku+QoP0KG88OkoAT17GJkM4BlTd1Y14zXE79tw
30rqbE0CPcJQCRpa3P4i+hvsOtM4SjaQIboEUbGko+RH6+y60uNmjGNBd4m2dVRiCroCP5MxBfcT
9KSeF1xPZlQmZZ2RxnR3LhH5CKt8tlJK5xKqFwI+x6h1qn3lZIUl93bqG7U1UBNLH2LI/rHvm3/x
5pmsrvbdwrVEmT0BdweGyf+Q2bEqlmjll/4mvGSy3IAamAdlBly81Ry9IU4IRzw1A/ik3BOVCEPt
eU+wvWybzR19368rA2Vk57elr+ZT9q2E4AURIVoVq3tZGsE4E3T4qcPKrBQDoUAz5ZbAt3syIyyb
ybSlJ/pk58zMyIM80oZ0s2AAn8UHKAiLDqb6fdC54BvBw6120lwXP+KYcEF5vbOfBMbWjzg0rRuR
ipSbENCatOX9P1GbhfXNSGO39wXOulfP7ERsJBTMu3XOoFEeULLdVUBZzeuoq556qNFnJByUWnDE
VzNqwGHopw48oB3V+BEKXq05k+0uOB7bhlLfI8A0LfwTIm6ykzEudbc2m4hXsw35sKvGIdI519L9
7fQgomDRM5DlCC04mJ4L5DWilRJEghyoShZQHTc40ss5t3GOjb6e3z1XUryxWrLUGtDtflDkdjho
46boqveLy3hk62nydqneGiDx4KNym/QAPSvn5DkFMkwLq660/tvKfSzuMwg/BRKphEHmey2YWTKd
OYXXYcXdOyiG6qH5Le5mA9iHWcsMZx5sXWKXQ+sRZU/Zu2E8iQD3IWqH62Uaz86mJJKWssn8asBn
cEWZd6FVQRqzIJvyYAuKNnnHCAFMI5jcpK/8YgsW+XPUdFoXcYb58qTcVDs4swlffN3xoSxOaTlH
LgivyfnRnN5gZo31me58eRDdSLBHwbJ9XR7J3Sb3OVLo/3amImzWwawGze81c1l5DSvOJ4cuzIYx
nYYaAmJL3J55I3pSFMMfl8v/G4Qr8VIva2RiniLnEL66r7+uWJIfEVgQWdjXA2GOkrYtwV+lqHgE
LRcTVY7RqlkohJT2T+btYunO9mcpHhAzPw+412wRimJ81nJw3TRlpP5NygC+wQMyIft2ETMr+n0Z
IqVdputO9e3qMPQRfHZUAGSqQZ6NuaL8BqZS5awkBcUdAXawkUkFxfbzAaOjdk+VujSq2DjZkgmg
+9Q3lFFbASdJt7PFYJ/iGoowyrSKDPclPPUW4SOv40y072yC8XNHhMIo7YsYaYi9zeHYv1Tf4nCg
TSDXs7GQuRLT1/2Kwex+Hu68ybxt5KV68gahbvMGsloA5yGKE16N2eHSmGfX2rS2439bDMsfzODQ
MrhSV/6svQlW2s0fng+F8TPt5BGJdOPLVCoaLdu/FcLWAadH0hcGz69VKxC6jR2+jrKuR5l+1jpA
1BnkN6GwwJlPWj7EPtosSN0ptCQUeqYOqB4bSCaJBYCApWzL2bnkLuCiRbVcOAJObncf5fIrP3mI
PZ+N/gd8Z/L8IU9Eu11Cwoxwm+n6rOP0MOU3qaZxhVQKYFkr7QTbb7TuYoE8TAc546GUTzRDeoqG
ONVRWfyoCJchYNoEXK8Rcd/1GQ7A+qO1bONE/+/0hfOJK0APvxvdETSVCtwLinm2bluxBuOoZk/d
nT1OZzTabokmlrUnnYbpeeJjecet3Z6bPS82Voi3dnXSjnkppICIiYsW6Mve6rGLCEt0ZHNnY9js
hN/5EJDVHE5hVcp/BXDIFrI3ZHvfuuuxKbef4/KmMuNk6wMRRaHfEaAtjzF73tMNuhx1r2o7dQs+
DnSlsCiYplFD8et6MRmhdsRN3iRJnIxWoPZuZgq3r2z53j263K8062xSJuT4ssc/7Cf79U8YsazN
OIdxNPaf4VMY7vzM6cbcijP4SpamxumlsiDTxIAu97Avvy/YtJbV5HfvGQESqXaDNV/AuZBluFuS
ZyFF0StZt0nuiDpw/b4CNP9d3yr8isXptR+o7LBiuCG62e6VCX3tsFq5+8JCYvEE7eiVWjHvgD3l
YhGrnNLNTHUCZFYzZ2Eo5flCZ7lusffPInhp4VOC1JhnrpAwH4FXQ+hsCPAbIOgbqqm8+gc2pR9v
sA2gVVvbh7nKxBhsNN4blM9XRbEkIkGutRFbw1rckHJUwNXj677b421z/XZSGW6XWTexAEJAde88
P/4bky+8X4S3s+S4bUVllmbo1UG8aOd1dlB1AWYmlNforN97F1kiGCyur3IARZav6Lhmzk5oWqd/
c1Ucn1gjp2GxPIwVnj3ZZS4Nv6QrppGJHg1c2pdD0J9jZqEvTKtqvu56DlF6aSf/uo+/uspYZMpb
8gWK5GDT8WLu2lnCvQ77fIpHNQQ1jbuiATYn56D0v768lFGJNaAe7gpdyacdbBfmZeS3STwRt0Fr
37m0ryc8fMOLEPTocKR77OlHTdBCbZD62gIQrpmZqrHuXqnosK75abLuDHXneSiCTemzZgYFbrH7
Zno/bnLdXdoEpfFwOI3JXGByB6xWQbPVZnpFXxi/yy3SKRZsC4hMlLiGEHm8MxrbGxIVjXDa/U7Z
od6FNOcS+epVE+cXTteAu0wrFyJwStZPMPjCHCJx90QN5G3AtbBNJ5ktwJ0IYv/Mf5AboBoQKjt4
ATQ2y8/rqqaAA+/CP1eDtxrue3ss2X6F2teuyTI3+io1uGHbpeJo7Dj11U9MZVA+jIaz/4ReTfAQ
f6g2OAbBvymGuUtxoEJteF+nPEjipj81BH94CvIt3XRwDtiQjcsrEKumQNY3skCVmfGMKkdBcnaZ
w4I2pujBBaNKw1uj4gbmnEwquXQYuaOd5saXFAhtjILxRT0cEHINF7OUVoUofTdwFiWgoZma/BFo
6yd0D+RlNpBEx8IOepawCTFc9ornhv+/nqEm8+Gcj83lycRyCZNxIPXuvodPdYew4HTJXg2UfsTE
NFrWV9TWMpKXvWEjuAk1TAbJiY+dNvfPWes5rta0/VKYxt6r9Ymj9Ad7YuuaeXj8gc5nmFNfdm6W
yjeP9ZpZUldXP/eL+FBjwzvqBvgPWjaSZDhD4igX6azX5WG2qmX2ntOA6U3Uni3T5UfvubZIczdZ
2Nho9Qu2GoLMDyzkvRRrqU9rdP5qn2oUgq74iSZK9xXBiz0CntPhr/TlnNJlIn6URMWJbhIbVhdW
rkx64sk+37Yt9AqYsYryopTbGz/i2z39SfdffErdsBCbw/AW8ZOiEenJgGcGiGkLlJk3CNaaLE+l
1NUVasYZ0BugDWGm0kcQgmho65OeGui+L/HFqN192z1ruIrcfO8KyvLyP4Dr1nRnUr6Qd3yOeLhw
fyaWJepEWtjO1bGRSBdWHt2oLE9YzGevp6NeAl9H08elYN5tn6Kvk1DsAtvka1c16jeS7vvSUPuV
hM8JxKz4NiqE3ub+JBsggd9rcZ9Fwmgj/ROKF97vhJFhtfbTuEf0y4ZrfwgYf/YpwVDU4jVbiLiw
O32GxBAsjzd9YDJm1PUib3qC2GakKkEbtCfrPGfet8NUgh5Y+xXRBDKQI/01xW96sUeMKxSofpnX
LULYfOJQUjGR1OS9ffW2ZAXlJTKcMTc1jSweJgoTINuh0/ek6M/JRUUOZk6kAJqgwwEsy3dvBBNb
3VuaLyIjDWpXir5AO4u1hAToJhNjJlwss2xweDy5WA3nJj11zpcg/tV0pjkoJX71igQ7Zf2WlAN6
8Kb8aOVYWv7Zr35ls6JN6ymK6rh402PmGbnUrfrJotxN+C5M+t3CLNHlvghp7+dr4uBqOAHToSou
up/pkIKg2wJ3wI6WHGXU5e51LBtRTHnKCBw8FD8HIOJp37d+zQc1N0pSg0m2DAlAitkEPejDDxXO
IC29kOZuYHX74kDv4Q7sdMukxkPXe8FMWyoCbEb5N0bZf10tlhWHcf2T0Aob3ucpMCNnJ9Wx4seR
nru9sdWbFm9l7xV349o0zC4AQpANMRysMB5eRswat7MI0NJ97q17UCf+qBZ3mh2VoaRAE8OBZkcU
Qrll8JVIhQ7UnAL83Zw9zZVE0aOdI/S6S3JT1tPdN7vaTLoMVfoUk//YRkNfW5IqwQ/iLxMGlEiJ
JjAggiqZmldJvw67yH+ViFC8ylaRSzOp8fmEApiRjvI1uive8PaFgKXiIUN0g/nVHz3pCC59V89W
w77j0JHeOXW2PXM/0aWYODz8pH/W8e+oiI/W9Nd+RGgyISrgXM+ZSn12oppNiWRIOnbsiCDF2AuT
hyrGfXAOL5TEAOO9HgI2NayXfZ6o6Qyf3mg4NDSVH1SG5kwSvl4Ivo42GDADikIyGyCP61PRAngk
4jg5/ZZERfGMRyvP9V9uDc9E+8f0HSrPjldKDV+rHqGe/29lwSWxoQrQMSlXP+hR+dGbcwlZP8kt
n33PrXj+qdp+KgOjfsJ64YccjrQdIvVobjUIHgLapW/48JnXcK7QBZZUkeZfj87B7/8xUdzDAfah
KaJ3wa/nr+f1fS76q4r5vjsFh8XInyG2SNLUAxyc/1sCUDllRVQTPzxU+6SFKJd8aXeYzfHyYE92
6Jwa9rGssg5gvhD7RcdVO4MHYjfAaVUl8gviksEyM0dpV2vNdW7V7EQLcfGci7An/FTirFh7cBC8
DYg41jqIggIaYgAFPMBz3B7sEEQdtB+fxR7wKuHr67UM+KjHjt/VVPn9blATTYUyMLEUxhcWBinU
pTd787c7pBLDhoAwVVZrQthJV4pH9OSUJ5Utk8zDbHW1AFoUvNeLDa6C0j42dqQehDbfa6455Gyt
gjG+hvSJZ22DTpBDRUlemIKHCHStksMx2tW2Rpob2pPkdsXEuscsHm25KH7122jgta93yOhD6jnT
AptxLOuUzCPnrFKT2gtOP/OWVF9/DxW/cWF9SIYrmvgeRgpzgIs34xuczgbH6wHBZEYrmj0wfJVv
Qb9YPiE0CictQic4jz7BPYnUl6DOetSQttPJhm61rWSTMSjztr722E9hEqPBMxEJI74M+25rCFZL
lqlf0QIWjoHC7y2D20lizhOjriBh9NBGHJvNP/8uYy9fvaUpo3Ni3wWa0hFMMZ4GbVOc6W82+TVU
y3/izPivjZxNitDe6NIQjiwxwD7S4muob/3wPSgWFSmDF+GFqMAPEsBKlaJw4M8XFkNEp/6wLIiS
yqDp5hzAjbqm/kGqWz3V2xVZoyONwWOBiuzi8l85RV57pDiFeWCx8FfYPCfXGWTt2GcCfkBI0xKM
vL3eZB7utz9P6MwEJ4x3e8tjIAwUAjttl2tGUqErNrs/CcCOEzl1bSOSwSZwg7ghlTcPtRZkpeNW
vnMm0f7ExNVZbOx9ncHjHDYRO96ToTjWERjXh1GTl/ETFpNg+YTLFeLr+MtzNI9DCPhqFq7Y74Z3
km4hyAe9L7B9NCIqSYQLu5/vhY/pxmUaCqky0c7h2wk0dzWJIC9jdD3jkU05VA+FJYhye7qQW0E7
6sRYyCw7HLzSMCyG+tF/SDt0XZAKhrwsYuHJnr0J8zk4jgFkBFncjBIaNVmBCCpsH6XV5NHyRN0Y
FSlgWr2/rvRqXoLD9BiVia+5/lZ1w5bN34ViAN40LPVSk7CudVHF9upKGEjTho7MZqUFfl1gvEXt
eLENIuctt15cm5dY63+PKIKNLsDYJ9RE7qiTJEpI0pepQ0DEZC4COnTtAZP/H25LsSrb8lwsAnp0
ng08yWaEnpoAoobxaVL8+skjGr+RMBMtY2OSaYg6VIKskaYJfiHga/5lNom17SJgpezMGzfGPgwz
7Y5Ddiee7XEHx6qDVi7bQujsgbz+14prOhL5UsInZxBCScqva5OOWUpkXb/47c/Uzn/MoaSybaK5
4ZfYT3VktRWFaGd9l2lBaEBFTRGrdB0Nkw7nHo7YSixyP+UVr+z7IpcUlCUz0N0P9LonCMSJAfN9
guKB+LAVlx8I2erq5JFBwg2Wj2oeCGJ8/aqOJggUKRnjcd72PtUvRp+iVhw5Rrzmi+GtdDIg+D5R
HgQydVlMr7A2mWhCSNxcQ3PyUOqVazGkDVvIakjsTpZjJoKt76JG8i7+NmF1b8T927LLh3B3KVb3
3RJNkgfh8LCiusAiPjaHzJK/vGK0fnpqAq9j/lRXUN8Ziw8SbcbtDCqNvCna8I6dQld6ns1escWO
BlvV/AjKAvEKKll+TIW95xk1e3hQiCG/vj6X/V17rAfPkoz+v9/D8aROcpz35knvv9eFTCb3OY24
/M8Db6bv2XHPiPZ4Twv/MX9+tmBQNUEqAxf1OqjBbXjMn/bD31+nsco98qKg+z21CzWhNq+d3tHy
2frt19OqNBGR8aBnyfu6cK1RC5ZVLfKmQYJGVZllHyY8KyRLh333MsifTOUiiPsDaKyOurnjEHM/
natac78NZLK+0D+egQ+LpCuaRHf9HgFuaCsQR2uXq4Kj7/xh7g813k9aKjV8wUDZdLouiwI7KDI6
dO5YwvjM0hORbAP6RGdjvEXy23dE2LfMk99HRwRZqT9+7WfufU2Q6+r4IYja2CjvIUjEDnx4VbNQ
tGNO/GAIfiRxBaCXfeh8ihT+QbCsUYMcAkwYGKKPJY+UpEGeHCygkTKR5Dy7XJPEhhix4kc4ayu/
71Gb9xP9O7vzBkQlhwDUXnR0KUoH5y+kx8s0L5tDEiJKxcpfhk8Uf/BRAGtbMTZC/Q3jnfUpkJma
xwmgRFlEXceyW2wP0DyOQ/nFOFNoP41mNQKgWFS05v9YB633yv25zZtFpmQVgcMI2RdOzxy1gM/t
/MNqtveKky6iOvmXHjgJ6u4QQWw32AQ1UR4382TjHGq3VM6QF0qlNwxTnfjTmP9sjEI8ogt0a1sk
gbXPesVXyNPZCbixpnaYXQRFHnwslyyMjp6me1wYj+ubW/MTOFrZorRhvC0OGugDkOIGT+ghHpro
Q0Zu4uk/ZsDfWy577Ta3Ad//Db3C6T2QMl0EGCTNSi5iE1C10mj+1W4PDALlZNLbFIvXhGobjVUO
NLQDCnSvlqdWOs8gJe8adz6mSI0fAUtOCfTMrZEXj1brdptE+YJq/3AC/RUevkX+P6pNt13fv6LB
haADH7WyHzK1zB/ciLXbDdVJ952WI15ZJ61PMkRfCrzSAluRk+/P7pbtGonHOd1ecVQSHi0Ctu90
8kRNAx+kpjZcqmkmV3mOlrpZeXrEDNM7LcQXBeYQht4d+tIENfTuicilAhTiu1sxysCbV7RUR+Yd
VlpNARncX4oh/evmlxeY3PPdGHej72SPrJ9nKYb7wrao9BS1KqnyAMyfdqWyBPRQjdrlOQW4FW4a
wq7IBMqgqrxB5fXwd9L7ZMX2BkgddF2KluYVsdMvJhgDSCU6diZJewYdCe1TjlBL/Vni6lacAbSC
ojPn3Ehzzqt9cmgSG3OO2oklRvVRtsq5Vb0lcBunTIS7q1wA9tSo4XOIUEtEJGWqR+5cBGXsz5WZ
9hRrcKEi2EV3UQTescQo1uvfVtgkmCe0Cx4fCm4RU8BZ+hR8wWJr37BgTTCOJnZYgm6FGiOmeWz9
ZHe0O1x1DUFhHqMQu5X4tnwl+2/5tdfU3U5Czonx0yyK7YFUzKSgHaWDwlsyHQjWKYNGfHqGEP+I
g3pfvhVME8zRE03X+SJiFh0h3Q5UQdRIv+ybqpxRNre6u/17hUsX2g4SPSLGFNWUr2ynoRN5U2Y7
FXqgt4/hVqJJyvSs4BiBKuLxkK5n4jdGe4I9+IkPKPq1qz9aJ19Mir3UU2mCqb5tkwCC9zOHnpwO
CRCOFbs0qZOMZfKpmi9gygEhub2m3hKNlFispq2eypA4A1w27obraPhuaHOdKDat2oiZdw9iTtZ1
xzUykijdc4YUIggz1nosN+IU3UWwYDJjLCeoZ7yOM0w1E4GT8cKHlDHPi5DtesgkeFvQwdmhkf17
7ZjhhrWBas3XsbpexWw5L0BGvwYqmoIwgn1Xfk+B3SAnlyHI2lfaRO3+ncx8WfzZB1ZoTme8uwhm
S4DlifIbSLse27kvEI14MEYOS8nTfBXq6RIEDTZRLvsd74vYAMwes+J8moFBvK3+Fmz883EjDlS4
CgoH/p6t4XicBEFe8/beT4blOYiY4AdhEoyj8NkJPsJiD8Eog0hDdQHwgqL/wls0bkAE98YMdjqe
fkGsdB+8c4rBqz+AN9LlquVmdZIOHOWL2ZUHNAj0WzMGn/8Gw4EF+jBJ1cPXZ47sDxuGPKyA2oee
6UjV5pt4AtEV/wHinAYMCAZonzqBp8duhl9ir1ej4oi0NgWdavzzWkEDJ29SlVNQxlgeTc+ihB6j
Z56PkSOQGqg6cYQaluDneb+08h9jh/ethqg6Je/Q+7l2q2WB8FqvpBu+Q538jW4ujJDvqHArJ8pK
dcfNU+uMr29zaL/b40qGEMi/5XA0IJKqmLMVww7Uw+z34QXEgZGjQ5OsXFyNwvfChOQjbGtUuhKh
EUj1MTzj/7s692yxzWLaq00MV3j+HuuUuJdm+yaM3ThQ5s2WMN25ho2Qo9s4Eh4up9zGCbIPISxW
jPF++VZX6UpqZGVRjZrz0mqAfgRrPeyJ4In+CUeQqP4EQBz/QLSyhfE8ukOS+hhZszYUsrTr7nmX
HJ+zqd3/8CzgsMYvPadr863u6eupchIdAYUZDCuDQdQAiSFQ4EMtXMq/2HPQYrwsjhAExMZllIHJ
CxjY8jUGN9ZXZycxqT3ELX9VNAq3CMcdVef0Ds93xRgJHBviTg/0KqsejuSHyrYCMRANutdfv+X1
dA0PG8bOIKnknY6QiuZBPwYqYZ5zu/+3wIP3M+C7z+eeMRhjcoFKnu1+wy0Wt3ij7DOUaDCwUcek
s3Y/AyEzN3QOVgK7ocyMyqACfrL+lPlQ5HVixx1bObGkHRel1+Ue6pkuCvbBw7X9N7Cz55deF1Dz
lN0nUTX2D8YV7ulf+loQw/DgVjlL15vxgA7QuJjgEmomsFWn7RPA1TSdmZDSdF0EY0yJ2j8c/lNG
3nycGLeyxLgScw1TAQAYcg9lg+X5X8ig/+qdjOJfeY72fTioiBdgqJM7lmXlqVn2vvu82j0Yy95o
/yhRPc2XS4OS+y3Q6+r/WGWhpGpm4+ZjcIP6uPy7bHgGQ83bJ7Ih9Bb1nqGPSEgQHDIgJ2FqCo1D
kfDJQ9ublxdIE/n2Qhd/V1sxLtDdkKdKqhnRG/QO6a6UuOAFxaf6GBm7aHlqggHJfFVYp690rPyy
qz1bpP+B9g5NpHdQYtjz8sBQbeFmZLHtwiQaLfciTMNlU76wZ9Pc4YWS+PAbUP1ORidHMJTMB0XO
gVIMXz6bZtaEDP0FSYNJ2Tem0ZXiM9giJ0gvFx3feUsNzGKU6XQ6yeZr9EqLv+jbg5Wf94TUQmOI
dVcYjGCQ5YtNegqa4iApZmQRWk5IXWUkIgxxxWFbQv1ehy36ICdVdL4UBeAv0gajlZF2g0li/DV9
Zg7gLdKTkS38eNgnxysXRIUIx4XSZc9SAcbYsgzM1XqjU4yJiQeNMm3M8D1Oah5fUVHwHoEnk7rz
CeHnuvjwLJi07FydwKjyWUczNiWIoFbTWfaEdivu6wA7Hljyd6PrwrIiB49VxY7b72vJ798pLkon
kXLg+Le+T2OzUN9130xfZmRIQ6VZLCOq9EVyz6K+TQHrpgo6paDRLfUBlTbSU9slHJF6gR9BC/5J
6BpbQSej+NcLhxjZc5LKSgRQWK7aLU44XpOg8Txyf8Kjsbh8Q6d5qLSpF+1McHd+EKOqDrmfQPcT
VeM2+FO4dd78qSsy9sYxsg3BSAVyAJz5t37ptdRYYVhvDSvmEJu1cScyorVum0f0r2QFslLxDPEo
0myUCb2Pwwgo1V9ZFgkcuPnUMBNeLwY4nsjgZNl95Rbq4BIfHfgSaUybMLdsmbPh2qZ9rPsrfwVf
P11ywK15OCSnUNLsNrV9Lmf+7hzGAg31QUBnODt9WfIhQ8sNjcEy45mRxdzJPkzdxwo9C56ZUY7H
L29WGfmBWOO1NxDpyl1aX4vHqjKeU00suTImffzQa0l7uOn7O1lqs5KXyOd/qaKhvj/Ew6+qA5G4
rDYdO0P2pH80WBp4Js1/p7cgwYMuwsXl4oBoA/86Iq4t7rZJl+SqzVLl52F6b0OVGjI6TIfk6bKC
WpstVhwB/eHW9IunfBXkUm1PxlmDAQ3iLEplDaUVCCySd89I7l0E2zLaV8f2h2Xxzs69lY6oNNVW
fy59Q0u0zk9HtcvNrY2vCaAC/OkRf6yStULrVwW+mcPgRHFYrHQRMTEYRIbRx8o8ZYMyTlZ9+8aH
oLk32gZhxq7p4tMtW/pVTmjOEkwxMHIAtY8LlogGsJ+vvH5D0qyU+L78YXC2pl5s0qeZLk5xuoww
pZWBudXrwEXgiBTi38uTyArL0Sut8bcat9+2WtBm+pzdT9lknspP2kI+Zk7IS7czeGOaecQ6FUvG
sJYoQJzmhJ2enY6K0LM5i9ZS10OKzzntURkwSJ5srir+2c8ix1rmP0fTkVFeBv4wbqQu4XsUFjNR
g/BP3ESYyAjFj+mPdNK7cOSQJjBzrx3XPdf8ZgYOaDnvuy9L9HtQUwTAEND82eXJTax8fOlCSfWZ
3mUxd3g4xIn8D8ofmDgBMOwiSwXoeOAtVHag3inxug4ddqx14+2u2cSv9mfbtHd7Xqv4uly3WMyI
rQXjrLGgmjanpiplMXPcC3pETi03ZqqR089Am96va/wYIDtqmTMkUUhGKVddMTnPp+mDai+uDwRX
1GY0kWiwtO9DWasoed75Q/EdRY8f8ckyJx9kBE8o9c6gLqgwWqIvIFPo1409E98QrGh/2V7KDtHw
ufQMPSzh7fvQTuDCVNQ/R04sey93ZwFor0ZqZ68lMn38q/pd3pzVhHsLQj21KdqEa2YS1Zf85IEs
M6t+/nkqGY2XycCFvtjc1w/L3LZUDjqgku8ipzdBgJ3lbyW5pr1LfIqlnmurmxKTFYRD8jJZH6Gy
WB+dGdFdqhE84dlqJVmNJDP5i9YwoSG97sGwq3JSmJjq2qY17TOloMb5yfZjabq6eua629LVOx2X
JBZoJIxNbcKFCiQ1hMeqWECWYt9Ll4Xgaeqmg/bdG/puIkbmysKMk6rRN72sqYfwYupzVmgWdwIr
FrA62aKxTjLqATlc8/LC2oED0qO9zipkC62xgbkDWsQxa8uTOBDb91BZ1AXw7dJoJLnX3CF/PMSu
GYJRfWxvzvvzUZgSCrg93Rg/LD4nXJwwwLYSAAntx+dSu8t7+ysX+DldiFI8i6eBOSMiSbB+TSM0
OroisHGndu9DJpHJqMwdG59imHUNHog3WG94quYHFlHzf0voxVjArbVMLCIdJCRV239TLL+inp0U
Sd/f8n513hGWyooD1zIKETIS+YL5+6Nx4wfIfyuQ//g4fulgywD2KXhXnD6u8822cVMt1x968BPF
HpQx2wKc6trp+k/8qTHuw8h+4x4DFAW08cBcVDzswLidNqa/opCsdtetaJBdnRuXzphl4AVrC03h
QkXIM0AKZZaxyzlVWuVmS9CK7uY1qlc4HIccWEh4eOE+U4Qm9MivwNMkUkgjAzp9Ff6ZCWxwnDCc
fChfhA9GtDRVOT1TvReyaOsSdEZEgAwOn8nPQ/OKSlhtYYpc8fzmZdUs8ZVdH3biRz1pOiREPUyY
8jyYR6CbtUXHvcdnMt7Vy154h+H+sg2ggLXnm/WmmGv980tyI1wmlrG6eaD11JIB3/RmB/E8lLjP
P9jdoZPXKdvhV2tYJ+YfP7Pb/uXEw3z6Rir1ZiyEwmmlTrzc79FtY5kVr6TPAY9SM5Z+Wz9N+xFc
1qMOJwG4rk6g8QY/AAseEFGYSXWBlnYi8d/oZSi0Q2DVZWe9BIFgZ3l95tCW6pGRzQodKn/NUjAV
zzWb6C23gYnmjWHu6FAJAqA+Rta6j62eEFUqPUnaEz9r2Wo/2XAdAS7WU2BYWl8Z4OhcQwnJ/FmA
yYroGUGOa1ZEoU/GTOHE0cg6vXo3qJvS+WwHXRelswtqClJtHIVLBKVLPtjpwfOJXPraztLnDLi9
/6Bfp8YqxM0mugIzoW24elLSqjj8KEcdf+5TNR3ja2f2aBFUbBfP6mzOr9UIXEDiaj/Ws/Hh4DuB
2fHfS8ilJBd0ZSiB1Vf70xbK8y+b5+BVqKsB/OhrfCPEHSEm8panxVltwzsv93q1H6YTThR99HcE
2IZ+w2TeVRBDh4XOPOZDhLXCr0j7KxoYlvELw8dAwwI9GC+RjUDZ3883Dq7h00MF84tSkuzIHHJO
VrqQQK5uOQys5XD6GV1FAaygcQEXAAaYTSC+CX0mz8qH2GGTnO+UrlFoZUX+di4FImzjxFJyTN3J
YWZcBSMRanBQMO85fJ7MPghkoW9zzaOhETTjC9DOCuxSU0oOYg5EwJprpXP+4EO7728LNi1U2xbD
DaU1eIcRcvU5sEOold4pKU/7i2claESiyF/8ihkbf9quv1bmDDksVQRTqyCpW8LNtSmxVlNtrpQS
y0GAFTgG+HplYOGhs4h/ZY+/HnAmvZUP07sBf55zf6zcZ+5khBOnFVdJAhs6yHHxd9JIV0YpH2Di
a9o0Lbyd0517RBhSa6DRLX1otVwIhDY8xElxSzASPtjQp/Vnl7k3NFQEjEKvBCy7tdgNdJLYbKFC
3axd1G2UgLsaNj3UO4MbQtD1dEyn9fGAxWi4rPrNahnaLn+YnSbfy/uEQRuI6/VIX2E/dUsZBpdG
Cf6rdFP8VIY6dZA5RzGDp9suGlUZqd9blAYkF6gGGvs9MSIkLyT3oGUYcu8tiJJlnqafT3ZFfXaP
udgqDBbQIa8LN4VIupcv/ziFWFtVLba+ZTr0ISC980Cu3Qt1v5IgNp2U9F6g8jJymBIZOUNx7HBf
yS89tDvc/LE+ko2GlbLMblgDvsgMnR0IsTpQzKYeJmtq8aLSxuZmBVS8aR9CzU95VEH06Dm5ycZw
VX744mD8Gsxn0TM1a6LlMncTUpm0CObeHgQ3fTCHhTk17iAFZGFTn+MO/wyIoIBlyO+F7zo2gLYB
GBDXAWrjNWxlfMjP+jOBcKfRz7Ufo+tknjHwKRQ9Pqgmf3EIaa8SK3kAqoEmvVw1cgRCBNwbKW2T
r6LUTMnJv+4p1DxBFZPHooOBjG5L4rM8B98vAnQL4HOfi6qIFny4bGZfTe+5Pa8bpjpa3Y80a3BB
uOw3rLta6/L3Gi45g6SLMwRlA1J+W70iEAnQLtvDvBmnqob//b7DAJA6rZWtGO/YLBNkkKIVf8VO
HzqGhpgK4rcjkL98X+R56+8AwTXOEMBCwNnpG1DgTfNvG8O3b/HWPtki80TzYBIUXuCe11FF0EQD
C0dJvpT7m8EH+TDxIFSqk2ZHNHyKh+02jeKCCt0ROPfEUZqoK22kYEftckVxcq/i3yZOgXxThgjC
ZZSkmOULy0cCskJ311fvbbr5tCFB/qwABTexoNgq23u/wRW7wrGyiZEvL8XthYjrNfJjrvjkd+/2
CK/dU6sb+mNqlKC6ec4NhFjwZ658poIqX59fPGUfQWVCKvNOXyYJ8i1/UE9I6/X4ynuWJMld3cvP
HNY/cYdmBnyHXDjY/i/CbeSWXa65KQvT9Dwlu12Gt9NOZtIHnBkXijm+EzMBUZkjaqc450Ah1lMw
2BJiuhP0tHVLG9wGmbDp57CbbfFvaO9h5t13JyZAluUzoTRDFXiWQj60DwSTySEoRjXUHO1h5OzT
5lTlomokaFucqDKzHdvUrMZmMlEUOhBgI/TZB6OOv+xk/p4t+sqASbKnPFkN49LCyLaaGyuJReJs
j7E8ZzuZYAA4bgJtMds1hQn7htTrqurC3OSGSK6Nz2VgL0nF57v17MaoGF2eDOkQw4zZwvEc5J4u
tSI0p35gbB3zHENreFMi7BW4bdYkNgbLFJ2kfzVhnzUpuKHGI+7DfRj6e6wMDkFFA7Gpvj/RMmbD
fHKZzcYnftruDCTJ8emUwyXmsOibCI0f9OHH5NfQDlLlsn5hCBDVXY3vEY+b7kj5UH6jr/EPHDLc
Vkc5lumyPkbi9zRVxNyn00XlTu+RXFMcmYgqgKWKqIs0pxFvwCsk3K06mDqPSzFpnLibKvZbTloa
sBSzrunDJyI4RRjUcRoJm9fFuVrJKHr2AZ+7gZ0Qhf5c8O+rhArt4RY8rNvzkR0DgUl3hWrTnRW4
UaSgvXzitItDCE7IEx7+1Nybc/ddnfeQU/6F+NUbFpfykSXfzJqwfjjxc/I/kGhyJN+pBdlg+Obi
UeTR4QzAlFDyiKknT+KbZcweKaCEao7cZtfSlTK8Ynd48uYXQ1ku2ZdtXuhifWjzKJWidnwmhvDa
WViR+DgkU3ndF0Kx739xI78z63mEXgCWxLXGOjGkTj6FkdQXKjccnz0C9fExArKLokBzVd7BS8iv
X7zMNfjd/X6bus3xrGfKUGPlzalhUvzv5W690qmxcNRjBGNOqEU2NetaSOTPYmGipOtnLNH87yMN
/Nz4B34TlSMQaRXhCH7XbnSUWkc7CH9q77c8l37PUS0j9Cdg0TnrwA96vpsH6NhdH00t2CVl0xcA
MfzXggT5DvbXGvz0tDxvB+KIrv3Hz0G68c8Q86Ii+JDcgb84ktl20nDy5Jg4nyd7Gcf84N8E9wrP
cv5uyjSxQ3k0IKMZd4XNnYlI1zoLYeBA9WzxLPUc8hoTLVFV3qhSb5GDL1F3AVTAZyxFg0J7cGdh
3A6ycu/udLlnUaiza6sVb887jrBhLSlJ/WGTeBQV8XkNpLOAmklNAKBUaklbCx3Il84f3VtEb9vp
H5uT+0IFUBpK50f7MDM44Lq0nBZz78R9bCo7Vwb0qKCMGuwgMIA1MqiKt6WecCjq0dEeWVolOAqP
ZO5tQ/4O+7ZEj/nJcWH9XTfewr3SblNKovSb+Dmgqj/XkqDOEgjDST91vuwRO6G2TgaQhEzdFVtb
CI1axvW5QMuZvuxUw0vyT+VSNI7ENTaMz8WWE0g68zXJxXQ6jK4GyOy34YhCM/aCaBP7Suy2wP50
oCWpbDQ/uOdm3eW4WfqAHxdBppFBHJZLUzh6OGfhH6o4R2ZZfgikGq+hkid6PFJYPbDjpl3FvdIc
LLfPHMREkeJKc9gtiOXRg4f5zLgxo52dyrMOOog0YgZZEhhYbWEnjruZBznIk3+B8x7kQjWaZ+Bq
AkGJlCXqpBQyPtk2f+PHdamgyaRsBsJFlChMQGUzr2KbBjHxy09cvlsJyaHAGIly6hbejUm0YdH3
DD5piv/3hdTxGZyJ2IrFedQoZ+wxIOaJNC50hpeAens/WBEHqpRd1ZF/oNQMrz96w/Htw3bGe3bx
1YeoA8gcPtgFgp8Q8Cb/OkKTFWBICsEZcQmDrVVZi+kDS6ZvxMXomsrLy+3wP7bCRwQBn24FLdSL
2b/tDK0Nisjxg06ZaFkHaHj+lnApbOhv8cDv0xmUo7YWrGwwfg16bnZa4VbLia2qUPNXBjhVtbU9
GHU9w2kn3/y+pcPB3lSqCYYouyvbTiyrs36kuv1Q2qW+ZHqJfGPOxDhJ9xu56wZyoKQ/3GtR3L1C
hFKcvaaOVnt303GyWSvFRyi0oxvXjBFVIPTBTDaataAhkyMQVDnChrD58SwCQMl73QYcFydJMoa+
qTZW9vHv7LqvWINtURvAR55N3hIPIhbJhS2wZ0WZyfznxj6J3PiY9FNq1+fbUiIdNM2ZGOmLP3LH
NgmdXW8LpiOjynoRWus+/Ik3O+56cmstn7GftN34S/ktT6L9DbsN//6KsZmDDSpCjOjshcF6GGbV
LfOFKbEkU5lg5jCN36k/o9WPxQAHN2+noQl8VQwJSjGLH1WsCPmA4gY9ldxZneubbJoy4f705pev
6iqOnYeq3aCGr0dB4MTTLq/+yUroapSpTbuYtxR6h2qGETXCo+4WDO4rAuNnEmtOvetXQZK8pI9d
NGi76WGfYByqBWX6vbvwyux2jmS70ngEcTidUpxm96KxJekCa0mo12wPYkUUZ4k+GIw3wDcZ2FmR
Me2eyFpUYY/5gHkCGiJSTvmocc8qoT3K8iFIFyMDoge2aio5AdM+V4dUPEEpop/stLF9M5vS2lQg
ENoB4VbD0qY/MURjW0xlQH8FPSE+mubDyd+e2dklKC7AVIEUgpGqW58dky6CPkugivtgI63E7/j7
G4sTpmV3KJMzYxQ4DoiLOSMSGveQ+1Bzrc6bwlaYxYopg4ydd0JznNyJoFd26HSPEPXfDv632CQ7
53qiCbf8xePvnFVbh3UuTj6roY9B9hu9uubOveTDI2QNi/w3SoyRdX7rgJXWAFRZgKIRwNMQR5pE
Q/XuT20zyfGyGkF38P+7T4aFeA65Q4kZaD/36gWrtO/n2IIX2J535ckg7XHJdVouyFrQpDh7yD6Q
W//J3YX6zyTKZhy2FIq3u2JM3FtTJcAqBWX0LUwCuSF1Sg3R76kT7m4TGaaM4+zx3mIJ8cUMeUWK
VJ6Q3z68asY6RCXe+5NVz12fUJssVE5EkUfnyjTzGse1bCPW8s2/hqHN3s95rVMRsuYGdTeyI8jW
BKmYZIWTnxAzR/FNpRxyISX8cmmfcmtqENMI8eHBr9IZp0QZx6Tiut533bxTQOpQf4d23fj1v7wQ
em9ZhvY3U+Rbgo5zKHYx62ZG7Cln1OXkdoH5Oxto2jL/UTP3603qYPRRf13RLuzAbVGgjybmI8P6
eEwA79XvuaFQsHGdj0OjGXzCh0BiMeF4FM+KHxhvvrN2OH9RL5Q3qATfjTh48ISz3qs0Ahl4JZBf
zs988l2nuFkbQpToda+aOs3MbhQ91rXebBG/wABRHOb5h2UqGNqoW+kufbRlk0WJ3Pvda0QzUdsP
/VgSjgjbQEHE4Z93rS6YYGjxSImGjARjAN1jwK2Ec0QRWvGnhtOrjZWn24r7xMnNmh4N3Nh+0+N6
smw2Ki/sJX7N/xf/DSo1VPX+Uq9HinG4AhjFMP7sQXOjKfN0PvLruW31ewZhrANZYpGu+bZ6gsUu
lB1ILI9P3qZ6U8oUHOAWRgsvCApPtCs4VtW2Of9qGkC3CE/DENcewDDOOzt0O4+fFAoViNWHIABS
sM2mZ0BBvXZToTOmcUMAlORrvf/9KsygkHo7E7r91n9NdU3ARTfvaJRFpJdFQ3nrXGBEeBc3F3my
YTat41eCs5x31m4mXr/WqH05pdFm0l5Wz5OWOWr+2EYJzdNYhatIn2LuP3ZfzVBe31DP8JG71/Iu
qWCVqfDWrumD63ASsjQco7CbeBcStvY2YQEc7qd3uu6w8Ec4mDGNqzQHuHpc7wBzdi9t+qCqhf6M
IhVtLKVx/xU5Zx/yjapEBJ9kLLsjIW6Di0aR6bzxLTYcovDQgJ38EusJABDoS/ogxKnKJDvL42Td
Jg7wfptO/aIKjRSirEGxPq/CMQtGMNEmtgDUptvVT536apdV918ucrbDiLjqn7EInG1Ci80ffq7o
nrB01SLnOOroMED93bsErDITfhN0YPehFKIDE/clQy1aBd7vvTpN/KmMDeQw8vRJ79NWG5WVAL/x
lcp3tmK+HYhHRcnxzJmaJPVhcRUGWq6vea5P5F7jttBmd23qs/ZiISRPdDpx+9EekFgDH5R6s0ZV
nesAs1HTRguruDV0wne79KiVc4GNQG10N09BcckyG7WHXlRIIeUuOrExeM+NA1oiZtOqbhFSxlXO
kRSRaW7WOgLSlMUCCNMNfvbbyKVwU2M0LwHg58f+T/7KdofWTq9Hn9kuXreskHsSW55/sc79fouh
gzTbzI7i7dTk9oIu3YI1lT32QcvMPY4CsrKX2LsMEZ1/i3QUASf+FoJ4p0SWSUJ0ULwg8wpBs41P
Wt9gr9hbI9sm2tLxezjWD8t7sWoLPzeMPMmmBUxU0vkPmr3QUZNnCS5zdyZeTtIN8AbvQew1eVO6
udbLEPOqfwB8xGoRQcembRLp4Vad8XdH3w5sIXm2PK/vD5wMBofjNLhbUESwhmo2bZ+ybHN85BX4
mT/Fw2fvruh7OYyUZZM6gR1v9x/ePp3aK1LqN7Gp56NuU43NCx/QDjOrBEpFC/fpJB6d+UyrdJ+E
f5GWsJG7HZcDnBB7top7vLQcr8/8DNfpuLuhNEKe/YoFH0veZ863yalPiom4s+Guuh5q/KHWlx+f
wOH8fETz6ZVbQxdyMFCROhW+1bqTzTk/+c1rQNVoFbvN+g+v36p2wDK6YSLMLG2MNjKV0XXhGkj7
hpA306TAAboHT86WCw3ccqew2QvsXgnyErSILXpcmYgOaSHipIqp1330HTci30GqNJQw4dCc5JFp
OoahA6hBaOqQ1tLFRcd2Jui/VeGkR9jJcREjU6e0H7wd5m+gU+cCGTLv8F+xS/P2gils5IeXDnED
ZFbKXkl4vE/dXdHwBIsZZGKzNNsaV27j3UfKIseqijuhrj/Mhsc/+lyJ3JBtj6S8y6rOZBnF35bY
KMW6RGAZXT222PgpiYJCFb9KDmT1Xj8rZ7Lo/L2HDftAEyyqKt2fCi2JMxjufxn+OAGVYcUqmTLW
JyIa9HjT62gxxomrEndsq4UL1GlqZ0wyZdRyj6b2/F7jmUWRpN4d6qM8GLgSsPl6kSsAs8sH1HeK
H64ng/1hs8Bpdnq9cwj+UwTwhDAMcp3oaZVIg9YFBw0MjKgWVnabOWJ46z4Kpp7rOVMldE7salCU
ql+XOw0p5aPq8plyQrVERAjWM0F6Nkpe14VtCbVFeOaFSp52tzTD0Ab203shT8k1A1680Truv+W8
uFOzqh++n0RrldPAuuuywYOE84y+f9p975sGyW80i3Ixur7adEkETRDTtL78z/YhbTCMGPyVCXIt
Zl4Dk7pRr9rZVhyPveQoqYAIqekpX5Og4+ZF3nlYpHRhrSo9+k3oyT/kSUUofqT+XOHUY4E2yVqX
Vp2ht3KuVahGf/w2q1OL25be6xuXWzY1vS/fTdRCpxDsWc1NHjb3UhONwZy8OqGrUUMz40IBvd7z
B+4k/5xA20HXThapdn14N0KH0cjhVf1psVXEwtUBeV2F2W293ieBEzuAgoBQybf4ARbBCFOpBA9x
6f8zTo1yZOozi0Zopszb85JOl6ZyQKLI4rXhBoR5yHbokUr04Van3XKfGxQLGw60plByNkJijDxE
LN1wwZm0dmCUs5C9QHi5n5cyv/Li7V9edWS2bgOmSe0jV5wITTU5nQlAd5M6wLDcT4cDXQSbU9sH
01n6F5qRFnsHgU9l1NgG7DlPRwY78A380XdDIKrZAIWnSaAfhbhmeZrbr327Px7gk4uiLPHMPuZo
MjhMrcOMAhOOzQZo8YqDO4tIvVTakBWF8P5jtnwg+wTODNIuRrJMr7C0qpi/chDXq+Nvs8XO/xEK
ui7AmxE6kgXD8DdzLRRzhTZZlUd67vjxII1OUctUuR4HQDY6EbLqJ2BDH9ZxiKsa6bdD1v6Vj0YT
+X+Jdbj9yDzxBEmdn1IgseG9vs29yfmZJSOERzWKgjiPR0Xr/+WHKupT5SwHxprn3BEzQLsTEF56
2rX6+aRsP273r3vzC83mb8mUpdJDRVzkjOlHQrZ6zNXT44ybFnI11om/J5fO7xn57fYZ6HPvSRXE
q6pzc+7nfj5yRwBy61eSME0xUThnaOeaIeOLtvSg2SZ28d9zImaB7AHnbJg8oez5JprbQyUPUtcu
N1flpCWuXnv/wFoVLIt157be5CGVDW9I3idzAxOP8C2zm1EGSxThd1gI/toGdGfWrUJU5dd9xcco
tR2IK3bgP/pjCgzzjenU8hNNS64k/SzPWKhdZ7mzFI2RqJ2mQSK/1OxfVFGtsyBNfSeYwAFESQ+e
8XB6O9VOejVsB6ZiPBemqwMfkS6GVNd2DrlJxmgX5JsOfxZ8rVfv22k3kbogOE2uYY4XWellfNRQ
y1AGg2yvMlDXhgZOicoQNfLjKT9cCv0wQVi7ky2gjCogM2syHu5R/AM9IaSAfvsYsZqWFZ5dXltm
hhdNVrLkOm1I3ojzvSQFLmqbIf6HU/z6QKr9VgsNeYbw8FtgsOKG9jpgQGfxl8DH/tsbM9OeET7o
UqZO1iQiRvBpxHbsH8S+b58dKogz83Tsvcyqx0XCZxEWst9sDHQ+VWmSOAMZvSMoS+971wWSZcII
s2Ey3wsulEg9Bv9jKZb6GbQWtlxYbKmH+qBbxlvZWHG3dAdkcbWPpyo4zKSuyPc9sibg7Ox+DpPQ
gNZbiGrQ9ogASydd1Z1FOs4Berwwn+3eFisRtKDJHsX653Wf3x5+R7O+CLtPrbl40foT/XE+rf49
/ij8tA51vXkabu0AzyoKH0/ATdHbb6cLMFmAag+dPtswtakoFBPr6tktZNgVm9q4aLsrBFwmAxrZ
GpyPp0I/qsd9SGcQm4kLAXqm316jbQsUoR/iO4k9ddzb3YCg3lFzeNffu38clWZRinwGL/9XiFkZ
aCp2GQGG9TJmwdyQIio4GcT8L1c+0gSzrM2c6Er8HunBZbYW5am2HNdksWi5TFIFTPW1yYs7bK6A
TxcnXtjY6MCv41/JjhHQCvPBydARIPRCk89myfaOz2xgZZyqE+Z6os07rttSzyl1tYmL9nr/LbPg
SD/aqw4AAKOrmJB9ddignp9Y6hK/B+W3lOCW4nzL6suBrO2k8MKJvLpdRuKWkFkKJ7pOCKdMnaub
hKrwM50Wownmp6JITh6y2AhhcKFs6BveXm1EdSsnKOwbSd9GPD66ht9Vx8yaC5q9bCaaHp4zP6cC
4pybxYYOT5wOFBlxfESfmsm0onfeP9JuwJ1GSV6xeUy1/LP6Ej5ndDZ6pyIdxPxtHRuzs1g7LvEc
ZrXDkxgUJykKvzxnIQ2agYMwS/ysDH8P0x2aHuELlgN7qvRn9Mtr1PnY6MKFgqpy93zeerjKEPCh
PfqqxyKjGPNpsfXVsj/H7aW0gavbljIyiu4IZSEL5Sp90GJtIa2abajlcGgShKZcNm3kUkZ3H4Jo
EAIIzTJhtc6GxV1g2VJioocYDxiUotrvjqvCO4g8yk7wB6AxttxM7NzjDKcLSWBzLfFwshPYtYH3
jyLUe8dFw6y7FeuI7anAjoWGHw0pNuV4uSSmdFFBqrhCCFwYnaAQbLz5Tk12wDOytBPXTkLoGz+t
Z0KP35/S/T9l9PqUZCdComC4+P8XH22N05TrqImIGL14NQGrMp2lnyp9khBVvgraQCdW1MsJlKjf
gUytN0pCbu+EhASRn49cMMUg3iV7RqCmIM1nQSWBWsvEYSKZtK6gCKuJJxDeGi9RvoxhEk0Iubs4
tnd5IeE7aOx+xY7jqoxhmADJBAfqZ7AxiWCf+xX5lmSb7N+2dg43hE/f4yvp5FGBJdJ0giFLBXcO
V966/rXsr5x4ARDJuQ6omAKUQVgGnz4+SkNeM75bqm4UqNuUrrCoBN6p8ND/1VSsarFXXgwtFQJg
B7hsvjSUQBLe4yPnQz5x+MA6uiDIewDM2ouuh2qOzFr7FLBYGX6rdokwchL0d9wH6Qx2OOa7eW1v
IgvL1uRmRQGTKhtztqg0ZCzphfYW/kHETpxwoT8VKkUwxd9YvFtvzAD8MdAY4yvBkgA5f4Byv8zl
NTF5KoVGMK+9la/V9TpbLqEkceY57IiBzVjFVzgoNFSOiCrLRo7EsmfcNWvC1xV0Sc8AvlDufQOo
3T18LTF/In30hUmZ8Xr0SVn0EdiWspGWOV58NNFvjwNuqtLlVSRD29SsYreziUvTxehd8NzNvFov
b2iAiV2zfJuceW+z8L1pMUNlCl3/Kg60fpuL0cMJNNUqh28NFZhvx6ZVmRFmfUbpNRY7Fhgv3JZi
CL1veMEWvXpspQkKcCGuKrrPZHknh8TxJZ/3tjUDr/WZR03TmaScglwPr4GZsi3fwRcoecLEZKlS
IDwt3CdEq6biiHfc/6NhcHkL4Eri5ZXPwenesRyeaM0vzuc84QHKNIm6L0kxMiVnct+rjrT7oq0F
Dxaxw30XjKZL2OQ01PMf3uWDayz4+rmcJcFwaBTJyv5pNQah8lw9s4lbSndIe58pSbd5S5NNZjY1
oO0i1FhnpRgpoVRoSHnB5BTndptyZLGJv2a8vKtYdsDgkITCCKh5rIVledy2a+PypEzC7EbHgG6k
eizw2enayd1mfrTjd0iuvw40gHcSLP9TKVzlyHynxUrwmAL5h+pK4iTuCvd6Sz2ck4Ghl0nm0t8B
eKfCjYs27WgyVWmnBvWhqloDIzE/gTQvFpiOZ6Y2ddx5Hhgt5ZFnG2XD8LDJP2OpSz6c59fGh0Nt
+sx/QFVLptkd0XERbgLzf+VLWwCfpFRMwc2Hg4bUmHm+1kSPHUmtZy5dibiRgiIZY8wrj8p7Ux5G
Wm493m0xfUWufrFwEgCQNR1uy4zu5B9gPGR7Ben7GS6Zkno2BjLIzhhbb9CFnp/A9578omnceoJZ
6nwT0fasUt3BSEydiyknc3I/kiepbik8nyUudS0Ggcd6RQPM+tfqOXHzpcYPqnnsi2Nhyjebm+y5
1n1YNsRh/dtuQKMNy8Zqqm48appvAu2sGDE2FlrMOy7sECsgFro3ZgT2lDIvLDnE0ghkAIveSRxC
+EzxOZF70uPrvtmrCxQkN/Ds+/Q6zznddUZK4fk18zr3UsFQHgYamGf+I4MUwjnhaza0Vmbrf+F+
XuFoHMXlOX/1anzFS2jdse8VUmEdv0F0cssXK4SgQqy3K6MM7rqJnjCYV9zkSMX0O5GacCWqx2YW
oO0Xgb9zh/rvuNnLSw0RkpZXeT0j56A32ml9AJuQG3G2OH2wGNNmUkvOjh3QFKoJaHMfCr4VgDlm
3hJLeE9NLW/Xj4USIh0qCc+myWeEq3V5BREK6NE4LejxkAbREsIkZ+UWtjhcG9a+YOnaJo5/eKas
OgmK7aDnwwvCzcmrp/ZJOymCDyuWSD+L490VHXlZcQ6fUAzuawzJLBeRBOqxgrDkfjj5WN5WhX/T
cx6a5t1vtyw4QYkWwCTwgIpeaVD9oYYv7HxxqGv5oIyghKxvzX/6fn9HILJt8wEs9CrbioJAFHWC
o5gAMBY3GTSB/neLbH6mB7RMN5ktUkcPK/c/lJaSnloMDQRH4IFqdjgx10au4XuNZ4s3pIGc8mQe
9p6RfqYteh5muQYPIFxvPnl2MgvpAE9dM57jvcbRBpQNDosh92lCAorOVvQXwKf/XubD2FdAPKJZ
rmgTParU76fnqeWdHMwaP3pbyUWtObZKXKZzkoT+1waDoOOQ3pYZkpvHzp9x1AZNNDhqptYGPDFK
90twq9Q3VloexnTUxbpjXUd5o4W2630/rfc7rtckddfEuzR3dOQYeGj/GpkGLDS88wjkwFLUqut7
aQ6sOhqYyDOiwimd3r0G1bxH3cKS/7rrf/CHKUI0FKeNBpz6ZySd1RwhdVn36nlmgU9IxLlBQ7c0
xcNk91gI3IYcuTnz5dhmTVTE7BUzF1fklv/7JrOHBXASvwPyIGRILdzSb4ppKg5POyQEPWyIWl+v
EWPVHT9FInOxBNDu9i53vYcb+bUCmxW4MnpQl8O4+tw5Z/ysKAtzg7UU6FISxT58JKedgMIvnKn/
/xrDnwm5Wa7XbQ9rIzwegp43bfQVc2tEUapT2CstomfntjNG2mJ0PvxOuryQYZXdxqdlm+MxzOw0
nnWakXxSNmTnbUuLJI0338LFbCXfE5WXC+YfkBYXANb4yoznVAS3RLOsbyIm3sh7MRRYGdwBaAAm
3YTLZN2iuHfUlyqKMqvuYguHvsMtGUc4dlDylwMTSkUQh3wsIBLAFQCgErHt4f7egSxpohk2s+bm
AMwMknzGd1L4dPSbr/st/skOfC2R9SLGftwAdmJX1yrzzyK1YS0ZB+4W5f5/Sx/kfD/Go1odHKfQ
jRHlttaiUZihtntv8MKNWslluCgEQnXUYvsLLWaaBUiU1OROzEuMPgQFmafMZDuOa+9b7c+FBDPe
rE+B+Z+o4ECqGMk7JwG7Z28/88QLPd0aBRFgwjXVhebpXd0eZWb3qQeJFGpdb9fMVyMylgs00G0A
oP76p4eFWLo9WGclq4ngFQN5fe6GFK9ZW3gG7Q63Ta8geEn//9P8X3s/kRCORjpQp4BtC2nDnANL
KCmc/SY4Zt5NgnlGpYpldfDl0HTJzXSlHpAIpFglqLvRWZ1LMD721UqjGxc8dXqtsDSDUvbnB7sd
SWTdPmI/9eyO7t2cPglDAyXl8Lb1O0LXYCA/JwPdtoawCKhl9qo7eU6JcF4YPvRWF3So8HSM71H8
0YkRv7v0ZXEbccs0snpN23UIhZOsJVO8UFfYQK0q+5jZEm0z4uIjWQGRXs9KlgvZkFjub+ShqRe0
FA7yz+ot8NR1l/sMW3jFSvVds2zPa4hRZxH1RymNoEA5GTRNR9nzP/KTmu1DfsmX8wruDXf4Zni5
lFCZ67Dv1PRATQAq2Fnmgk8BJQlhr6PgGpG1vXzNPcHGS7AqOCU/2YZwwrphlAwkDDwR5LzZCOGY
x9Awkd5/6IxtRHfbm6EMLcVvXE6sDBYvto0PSf8jOoxrmqM7jCO0OS9mTaVDj5OCSocheemdiHvJ
VTH4miAJCMmo9St2hZn5MAQY0utcGWL9QjbY3PC7aMWAPS+2AwHcL75n8vrQ8C2ZkdXlcul5NwRM
6QADFqE28skW68bS87Le4K7+kwEFXNDfe6+BP+we0Hs+/kPGRSdTeDKH98B8yg/5bZlx6UboukYS
TmZMXPsbOYQtipLS6276lhcteDppjUDgZLRL89xWOT3xnQrLqeLH2etATLV4GqAZZudz9u4HIY2e
CqadTiSmLleYQAfVI83vsqMqqWmwgHxSeNDQT2/cy/10Uss+JFd3eNwWBZ44qOSy26s5TFz98Fhx
k/UqByuPuj01IPrQb6UCvKgPkh8EvzCJTG+KQe0q0WahD4U9D6dJOIKqMTjmMR0G8uE6MGnMnXyt
chQLNjg8S8RodeYwYNOex60F1mW5XNlUWKqew++OExcIgztA2ycdKriChiqcpj7D9hEsmlD+3Hfa
54F8Mutl6Kl297oNj89LqYPzYRm1IzNBfGYSoFpuFHOjAi3U2W9IybKYiFZBAg/ngYgf05LV870p
1u2XQvTRCIV10HuEqK3KmnMD6uDMNGqbqnN0fS7j/cbF9TzuT0jvNSQ36l2Z7iLS8BYQRqRi3fi3
MW7YZ+fzmJFHijwMV5oboB2r43OjmkRmARwxHh1fAJbW9pJboQmT0We0OC54qsLgtNxJIClBED7O
7HqebAMRW1P1Fu1Pg9HlhwdEcqlfLbM3QJX6I4+Ase4tl8FATsdz0Vc9wMsk/6wkUjgMCwUe6dvQ
loPB5GqLAn+DlZ+tRpob+fwWY7QS9Vew0GuOUy8Q9+lU7g0oHePi+vVIWvwcPRv9dzRxGtNLkRlO
/l086SfjmZ69t/Y0+T3KweUGE8sVpldg7o2AvCzyqF/CZXT6f8nzzm/PIjTA/b4erRrLiF9gYfxs
JEG3g5gM2AUMs0ob6ssHiQviswG6KKdt2o9VCqWnrbBJKZXhPzFXL9Jdu+Uy6EwgZCSjA3OxLq55
a4cElq9P42V+VbXZMYL76jkrXUX3kay/UeZ56uT8tw/RYfb2isxwU2LwGT2BcPppzGS2fdbxX+ws
twXbo8XgI3YTAh3AMcLiC9hUDxW7/1aB+mMcw2qCH5NVJo+nXhJEc6UnX3qALlDy9mDFjiqrFd1T
ifXEv1zZ9dY+5r2AMfdpEC2Fge/vGW5q9/c8oyRyux7WaZ9h7BE6c1PRUjatulIzMB4zHAfbgi/n
BNIWRH2UEGdejQYoxKiCqejR18WEEsdIlm/PGtFYM/uE/R09w4KWwvtrXnvNe4OrkTjgV2latt/T
mFuKSdgAfBPntX7DYIMmHLwDpIoDt8Mnj5GZkU9U7j2k4fAZD80FzGtvA5otl5ZOQhIluwmLH/o7
pWV3R6yhv6o7wjRcBt/UUewt9uGtj5W+JxBWiDZxiV9ojaILUEbtGUibZhE4HybFG5OVAV4dd2YH
sI0OW/mmkzPzH6h6V+5Dny68jT+Sux4Q8w8/BAlVnbdgfHHfObUrLfYl7mBeH6JMQt1JPKR5o1cE
qxNYTjFHuwp72asq1dak8LZkInX5ICfgXVzsT/1HAVOkQbjxjeN/w+sHYhrmOTZNaogWYiR7Zgtf
77TKWZOSwZWhrcJyyvOKSmYVHP+ZCCYusk0baPVa9SYdKz+0tb1bjZHHp4v6JTluq01ZBxctd57T
Xu63ByZMQZuj7cy6nJ4qihTVRKK8S3qeOYYfvpWhkfVw5znxpk+hPWZq9Px1ox7eqzq3Tmf7f5M+
QFKvtEHZDH95LLAi13pVCBXjMM/gBqng7iWZ1LiQ4tn0oBeMcCgcWf7+qLNS2oR9JePljh/NGesp
xEWrylHk21feb3OQAF0oSqyCopDa9a5lCwDqGvdE3pP5Hzp8073SqlLGoUmra5QRxPalemLPDGsN
4//mQQfllfcPK3h7JPVPQxAtklZYQvVU3gb3WtNnmmR4neKW8ohnsz1Pz+YQPYVv/ee340Rx/Aid
g5Rx2v7TnVUcnXSM/B4dX5535yW0ebk3UCUnA56pJfmjm0h1w8dxHjy40cjOJhOghEVv8NfMnN37
XIUdyYxgD0u2MHhkoln7l1DGt5Y3Yl3ppxACI9sLyi6gJidyWhjKO4/5XpgCWimkCOszQye6oJ3h
dXrinG4H5LhcmjlPCXoQOp9ZJ1dW3yjViJIT7X5P+TQID5xRGeEMeoWJJpsHsx6YbwPemoleyU4y
j+VfnG0RRx4SYOS95dA5mC2IQFVAzAEm1pd/AlPy5+kGVClx63odzSui8i+Vg1q/7nTM1iUXwtC9
Qw11IohGg7kroZFK4XYFxehsk49Kx5rzUVE95dlN8+JA0XngASyFQnKgci/pw/EkH5T5C0Q8w2en
cHzGqYsfI/k2EXXcANHI59MJx0KR2xUR4wplXWrB1fdDE7c4g6OOWjt2jL0tspf62kDHjTPJavYt
XtX1PgzHk7kmo4IyK8Y3ZDAMKNR9xmc0mn1aDmfV4QrTC2X4CnvsurGKN2XjutFIbARAICOMG8dA
m5WpUG6fbV8BvQtUHa+bN/EcxqY3TJR9ihHt+b9Xknd51Z/JW6m1VSRINvrmeUb2LxgegCtAY7za
usK0CNsxny4oPg73SVeICnaDnqkME053QO3dfSEtPK7lNPEsgoCtVwTV2SmNDY0HeJWJk+pV6AUM
iG0CcPcyy8tR//hCrRgCHnML9wn1rsEgBLJ6bHUF46lOmxzVDwY0FBeryKtdCmrEiuN/jT0r3Iy5
fI++L4Cls0UUaBBskp3crPwmERcNGE0unr4wv+OfooZF9aUDcMN+jbaKeAjKG3t2yMuCilVUnBPy
227popgdxqd4GGv2Etd3aoYYo4qoc5SJYdfDtLCt9MyY+7Zdbtf6a+Trwbp8yoxqN8TU2iKM08cS
tfue7+NJgb4Lcil4hsO5quVWqGjy+r8VXeQfRGqhEuYSEAtbtl+ubxIFDsxLOLq1fO6SVZ80o0yH
OPJ5khhYDyR4jpI3MaHEbjmL0MCVhV+O/JV5VvVlCMVIV4v3T6hwbV5X51mTKJO8VpT06zsuPTtD
lZuMEU6ZmGuK4rCnkAdvzs2/qZPBcJWe25HiGcZrCm7rO+dq2LbnXLOLiOgLBSMc03wgtQH7wQfq
G2/Lyehk1NM3wWARwj6GzriLCtOyDf7ZxOyQrS1upL2wUvO1qT4smrLEWqnFrQt8ZEb7Q5eCJQOM
DTKZvUWhqmtvQGbHPhjsEZxDiAHka+EvTxlxV4IVHsur49zbgHoIWG5Yp4BUnOAIrQHJ7Qs7uotg
iLNLdGryzAgDs4lOe0hkbZz+/IrciTvi8mC0JleUe0GlWlyztqn2eF95DaKbi3dyj15uVZCX1zvN
DP8pbLXkfw232Qegqk5FLwJyupBNShgHR8QXAZybMc/nIJYDcBfEwgKFcogqLeO0+OzXi12kOtOP
Ia/Gb8GBNhlk0GiL3uE/gN1wJAXz7CVwq8f+TLeHDpX05dL0v9LgepWT2cPoPwfhNnJvO/6uSQzN
4WhzZKuZD6a7FF6i5YMHV9xs8POtz8SaYCU6bn7SjmtQDrhDF76XyynuUPzGGIWiCkheUwZHASr5
ibCKbF7Vr5Z5xNkEguP/sHF0dtCMZ/I9oRZ/lmastedoSI+cO6U01IbIoG32AvmZ/mf9jjDsYGNX
iQ9ZZsHpyJrw3yLJlr63XOeDcNVCZcfTsioIH5lSdml/jA5DCVrWvfzL78u7RnefoC61Bw6mYM2H
QyxQ5q/tVyWqCutwkB4CCb3BIkSI+y9zOstCiafI4FgGPz3g4IxgE/iJeolQcnZott4rW6Icf2QM
gt56cUYTizkrrPd3jzAGozdM/Lxa+Ds1xB1obDFG9IZFA1ftkJ1eDCJlgEgjteBj/a9fr6uHxxve
yHPNMS5UbNueOGDRhTquYLYd5d1ffLsQ3u7AntbnWwRmaAUBjhuuXOn2w0UcaHEkH6oN3MeP0nuw
VHWMshJ6bOr4QE1vYc4iFyJqvY6pER+v3/WsXAiYmWr1lY7HZsSEJLkzwg5j57KRrw1/8fiasmmz
EutPN4fOcMLFnSp0TUhVqscA7Xwq4acbxuJ0WL5ZKzHO7lcSFgyc6iBqUJXCO4ZSsnAV5KDq/XUg
knXT7AOGX8O99D97+F96gMOH2tfqkiuzIQbMk0bNxJbykTv8cA/2EwYbGOD25sbOkC3MhfZdDBJX
AjzYIS+ycsYzYOLrp43dobINq/vzKdU9dnI58oPglUtsbK5pRRnarYOVTLqPGUJQ1kFq5AXWE/o4
KHxcG3i9n09L2YH37/mhBwHrA9r5KuL614j3edD9ylMO1/KL1Pv3NqIcXOYMeg1G682LBRG49sSV
V5XhtopEmf7x9ciw9fFxNKZ+tf74EAFioekHBcqzDSZSSp7nFjCatfmAHip1C2Mp1nBlSluW1azx
OrcnGDpO+faXn6Hg4Uq+QdXjYxMOvjv+sEzUVbUlmEjviAgUixhVv0AnZP3r3Q2E8fpTjPfMw5+o
3YzKYk13wtq2S1JcCU4d3B3ahQ2dux3AuDCPyp857rs6ooNoVDECsNRu4zMFOEfinuWk+95DN/xG
iUAystYhI9RSeCyZLH6WwPV+60E3NNB5dfPP1bvQoYJvx0E8G3jm9ZQVuLCCG7zOc7gkd4EsiyFs
v4wP/f5yHwyR4g03IvliVSQcnb+32UvG3IjQnNaIQXPv6rX+DJ8BbJ6j30KqvCZ5rlKslRgubwMc
yH0O9NpyLH+1u9HA+9KjX1bfcXkPiG4bpiLS3RUjvFK4UjgYbTpsay8cwpAMJ67yRcufexTD7q0m
COJMBPobTgDdvxmn/9Ip3nOn0Hne8raSHIAJ4tNjkKinV+2TLvwmKn3b5Q7djPhzi6DDWG6U5nQo
QALlNoUmlXJ5jZk4c0BupdG3cOFBN4rW2GpKfpGHKR0SAwGYhR5FXovB4uzHoXWhs4REf+NT2dpI
lPtUBM+EcULBX/LQk0hryGSfgXSlSZ+O3UvhpWwV6MYZdGzIM8JJh/q8ERw/An0N9xSvSTIxtxvO
1jiTFn1JIRDZaBFkcI9E6cFPELYJ1o5drO10ZDtuVs8GwdHpINzld8oTDzeMofR1ztcex8zpV0XG
t7RXESRkrExPmJ1hjacJGp5mrMPXxE6g6W29+Nnkp/IJOSlFKjnJQNUEW+re/iMrQpWeQ0V9E7ov
d/Mm6StDz3Oohm1DEseozxYxLeFKuoQ+hDe2oE9lC8ABZYcZUiJDHoQrt55yUTHGwPBWm3Ajv6lv
uBVylejntrBqUfkT5fsRM2kHKtaIlPskA1Z6SjMrW7rhI5J7amvITCnNBD8nWd0wOd/A5m8wUssE
4xOp6EmYUNJqiT6mWCuR0Pm3we0TCiWhaiHIK/7tasV4AwUnRevb86XW/WRtv7G5wsDn1HMHqNEf
jZ33YyxrRhWvd+rSMn/QuKWX49L1aSGv7SgQLRY6Teg/9PDGteLDIMw5+pzaMT2GLGXEdnH6iylE
kbGHl/9m2o1swPOLDq9bHC5jQtv9ZUIVzugj2jG8MKe54p9AjnK+AGXgQpmaP1GqUdAWZ08LVqzh
xLel6WWQOvx3hZxWz+9HqLTKx/l8B1hG7uXQ4MLmqUyfdSXqGFEmEpk3VskCjnNZ3hScDbw6Iras
MiURmXG8bkiAaXmAZ1iZlapHy3hIXyMILNrLjcB6NRuadMGgvOpHpi6+K7Fw0LSwN0rtJxEcp+Dn
fY2hKm05o6c4VnXF48GChdcmdeLg9LdFSKH98SRyIpbnwyKEr8+NXnhRg8sQIpgci7cpo4pKSr9n
3vCVecyh74zsel96gZ0U2in6RNCNIoI7yOy6Cc1NiFPMO6LdLebosO1lYps9gZmGSp4fHigfdPKc
xsDaaPy9SUqR1CRxFs/t9KwQBNmkGxbHZf+f9D4icxCy9o2nhA56CEwzBA/J5ohi6hekACuJ7exO
zmHyNs9ZFnJHBK9j23+OnuIJvKmdegnWlrtKzTNDW3Ps60q6ShtXHXW78haRx5rA1OZ92Yp73oXl
neP4uR+Qx00vQixJPx2DTXCIKU1/mEcLn3P/toR+pGjYfNVOjCYy+P2iarD9t3iecajZB6K2u/WP
RcDyXDZ3jOlW1nR8TUKOF0bnIEIRkD0Iy3m2OkS9invCmaobFjq6+1wyaZNocnOc+8KTzuMeCS5L
kmV9RugxGOnSMmuycL0A2lJjGphYXcQLAz//nOzhxn0sHUw4ZMAU4TwoF63vjCwok6SGemDOy1vS
vRqGmvkiffUeQqqGcanc4odLSjcIXGV5DmXZEuQVSy2htL7fyahD77ECvHUk0+ahpTqPBnv0Ip2G
jnB8TWZ+9iEwhnovt+38Lb0Kn+ddrVUGe9SezvXomFOFsUEW6kXmAJj473Uo5ATfAuzNEHrRN/PO
haL37EEySNWSzNEdBCzh/2wg/OQsL4LYNS/mnsPm7bzOj6yKyhoLQUSj3dwcGFny1k1mi9vehf8b
RQrixzi+JIe6hQETRpmrkqQf+75WTluZVl8lpJzTR0cjOPrKdfwPh/g+X0ueN51e0eAfbdu9EYun
1NDSAKGHAQwZALos3OQi3Y8n1TBFoRM87zNy/A9uotvfo55cqt/hpkil8lKPghAoRawOjMewoFaf
d5HqbStwh+o4sso6aneLxJBL83obXJ3sHd1sktqdtH65yWfdYP52VhWj3733jgwni58HuBGLhjsU
Fl3LDRIJKosfUipimgsIebJsAF7dFrXOUaaKdH7bggQWReIY/UoXo3K+DiQ0pukSaaeCdcP1mrUA
0ZkwFjgdPQ7d8D+/SwspHhc9pVWX6CCrXROzY9ABByT304lO4CiayHiplQbTEkU712o3DKeeV/0P
ygiliUtgV69WFHrpY+VKExqtci0kNOdpTskkI5LSQLDKaYraFTKzt1QCVGBygW0gcc+agupsNM9k
I/GosC51ZZ9CTWwtbs6QS/oC1l7LvEHtwa60CYONTrcQRlo3fGKJSRTo5jVgSaINVYDjRdSKIoqA
eKEsuELgdXLu7kaQF7zWSdvu2c+7jB1rKErbUdVen844J3J/9r/7WGFf3bIxGmGy5NmdFxGj3s/y
tknFSVKinaHqsC4rZ9BXTVOE4UJUkp0HwEJZJuswazQCfZ70Q+flxXoir0PgyJSbdNX647ophLjf
/mFcuvU7eiMqSeABqJ5sGLOP9bw62vWDJ2uiJ3SGGfnkFfPhsRS7plJcMS7lkgVR8wYsd9HqUPHu
IIcNitfc2cc0sottYGAImOPU5yxZ1RPSD4/hnHT3BzjzxKOlIJ5YW1AymlbPzZzXSLSVCCyKmwLR
vqP2wz1nTzVlmCcMG2x+URg0r8I0k01EjnKcQkyWkNC5iyBLor7YlSBw82eNpRIZXsLgGj4MY604
/v35oOIsy/YroMr+EeY39jSQCWb+X8i7NtENRxOuCuoZ13lKnnVerS6jffliKqDfNTXsiGSTjwwR
Lrk3SMIO6Qrb9vJ/DtqB00wRzNPSOp0ijtxceNaQB+L0519rHEnHlK+tDvVV5BGo53zx79HAfFy/
Kl/C+obuVsb1oqfQaXrbZ+xUk9VD0dznxEzegL5J2DQGSYfMQkvW7OWVZS4KWbZqEwK5AeUALFZp
3GTOd0pEM2CpSI6U3W38jf+94sEQjxlfBZsnRBUPk20egXfQVXQb73uOIe88xMcsEkJqHlkP+Fb4
f2tpuDpj/x7ET5DsvXHVaG6/bDYdghG0ySKyw3lQPRf0dtaOGQvqQKvyPNA7kFtIQLaidF0TGSbT
ZdV5qFdzmbxQbh8PA3Ddx2dC7n8ClGAvcOi0ZCrime/jJYlnqMTvTQaQi1YW4nd2fpERavHfv54O
XlN7SFEhxI4W71hDohM1mnkzTPnY2AriPbZR6yXH9sbfsy0k7ukI39OchCSsgrhZlK4vLdr3busb
p6dEJvsnEXPvPKdjzmfWHgrRw9lM+MkH0e8G9q0nFvdtwCpsLx520ExFnnBkSUTZoEhqTanJZzOJ
rFFheIQ9mhp6Ii4nwoJqz1NK3u4SMeRnW7rw8qI93JDs86Jcz/4LJaw6ENXGIb1tkLYANef4ZNxJ
h4In7cVyzPXygoS+oKxpbDXi5z/+FDpmyRKJU7VzbMH96x8/JcCdFRzxHKslGS6OvMajWxxw6wb8
CewKCYWJ/cH61pzdjq6SvOzdHNpDaB7p0s20rvYhxqjJJcAr69rSPOXtoU8mK7SCoEevLkSYqamg
e+31db/wPq/opnaDkFkKEgLUJ499aUBacCjY/sbjslWIl77PDrgydNiWb8nJKPurfWH4SVIDBhwM
I6RgvQpiL8tMVaF6lphguO9e/U+n/hyUJnImo/YuZExBGXaykNKafQHoy0SIIL3JOOJW9i3uG+Y3
nlznTPtu+m+cBYxr/mgJW6DDYyydWFPHP7aoev4YxSWA3ggHl7LWC6TqMBPPxiQKscwA27ulpgQv
f2BaoI0cRK0Iaq/r++PYEDcxXl8X26Jpnr080+Aigr+LlovWN4cvennKvI5BVfOLUjf/R9RJ4ibO
Q0ShZz7Ao93Ap1jOCJG//zCNXQJbIL/mzsTfA6nV1OQVGRYq2eJZoc7/vK77MKOjLKyrStDtNTdl
05EycNIR86c61pry8nFVQEW8gTHUcSSMyvfx3xSNr3+RY+zGy6lRBlo5SeHBNGvkvsL1PnSyqN2o
Gu5ZmoydxbzTcr7px2q1TiLBD5keuNuc4YJCNUEH/KHIMo5hMfcsj6r5JVf47febL43hJIRTp+pq
bmw+KdjtKknUQHTSLwks2Kc7k3I2gcKVtamnygDLYjb+cPK9Pv2/uHjcULybiLKJNV8NUcG552Qe
d5wfSVscAVLOpx1X6ZljiJmmgJLNWqw9SdX6Y3PIbkM1is+J/oZmfkmEhBE8GOgsFIKzpCIJOpcu
fs1V/GqmZwomKdvIQxVcMrtiD0dK03PuEhYBJJRCuyU0EGk6G33GVef4UmMXr9fTRNjwJSTi6ZNl
8bXt141XMTRcKk3ji7if0G8CD3L5desV75b7pp5orcUjouqCreo27jUlMCHH99WGpZcFKYEL4BK+
5AIHb1burteHg5/LBNnbMgEMIdLyEPPCMGZ3MpfXXjPI70eeYqyuBfh6yx/dbM6jEyP5KhC7Kzme
dWbKSBFx2s1EEErEOAcOmEP2olvar9UDHzN2uPVnhC3HetJq7cBV3AihdRk3gQ1KN3gJVVTYDh45
e4dajzSMYcsVAfLvHnVdwU6yWhXWEldBU7ATvtBt33HlXl7eaaiaCEgRokq1fB8TV2ESgK8PHzwy
KS25r+gSZ3gEgZs9vAlczPR3PeltnNuIlT0kdiu73Idu1d04RB8ZjwXcawwrcJpw6INwoCb7YZrV
Mzai1Qy08srbrsLydHgR8Ttpx/YY7K69v6s3iGoXSUvR90HcR7o8M0eXKRTmteHj3oCIqL4TGkrU
sXmY75kXUfVaamsYyinnZhL8tevAbitwLaY7cz1w6Lt/uItoKbXKJB1OrrJvd2mAuiyOsnMtZwMx
69tLDBxczg+kJtGipdk8BO+cxdRBz7A5mFfACJC6kpFt7D/Q/Fou/ka6lIDjamz3cj95XY5Gyp7x
MEFmH1zuFkQ8HLVywwzXKEtzhWuANOXoVf7gWm4ffx8AumTF5qUUaBeP/r5OKApL+oh3zE79PWfM
jcs0h0T94BJgtgertNQysHp7J1xhF2/zwfjoUoig2K9EFyBJuNttektCioTHEGDBYejrU4naefQ9
8gi3SVqYrn4BbWU9FrpTsSGQLZiIA2AZZriz/eJzyyudV7seRQh0NVtvsHEXzrhgcUKaPvtWYJVN
oc4XacYlOo+ivjZXVv3RClFr51r7wYD3kfGO3Zx2LwLOcO69Dh+2UH4OiTYvqhSs7D9OGf7N2Fwo
7ryecf/vVXDViNsQlfij6XPgzgJ1FRu5YDRczPfuQ65/XTXSsSYZaLIQxb5hxKRihlUcSL/ixoRg
/CqyFzv/P3aU9zcMPrsOnCENGhjWx4UPD0KvGprF7DjnPe5dNUQV5LDA1FLgfE1fBJXkeq6j3xuE
Ckiz7fawp6h8Wo/0G+SL95u84zM81kLbuGCoYoDwHclW0KdAFH0Iiu0oFwzgsT+FR6IQykvC9324
pwPjnRH2vmzgVHJouY+qW33Mjq9xeqIsUqRVjKvH3FxPZ5uISJncbDAR/A9PvG1qy4i84aEc6y2i
9LiJN80/AI4U/uvvAvmcDVqekiSkgebQ+1g3pPzsNLPOCDvqBxeJBE+wS7JMAtqD7+Pu343+HnRa
Pj2+PZcgo+Ombq7Bd6jOZ2wgQuwDSXByvYdxFoXm5Zkgc9fZlFbP9MgYNX9eLzwoKwpjcEh6mUdy
0kZ4HQsG4lRvIji0heEiBcaHxukXzVzvBrzVQaCS3offM+i0PLHlvPu+WbG+q2ax+W2k1Gt1NcVb
E0chcapCcgUn3UwkWQJ+aSOeYBUUUyAOw7yBhMoOa2pQ0Cy7dHGTMc19ou1ck67lCuuyGcU0LTnL
x3RBpTdx8zKfzW+3owk8bWjWqRvslyJGLL+Y9m/FsLPD4fTiS9VmXBIYu7wynzu/LtMFn9MqxFtT
LtEXCHIQ9CvZCmE0dZwX4+Es+awfgB16qyzDDToVVBBUmp89K0FMQeMdje4c00dQB36SIPKbAKQS
L38JW2uQaysNHa2jqZmQWvXnkgUemmuRasl6BmU3A8LvyltXEEjqW7FKXczLX76CQ1gcVeg0V5jT
Iz9cL7qEINZgCaIWiUX1hvlK/Xwlkh0PHajMR9uW5NpwqEv/PZaK3BWOsv8g0Uar3KyyTJvyHxsW
f83ZskfF1WAeyB4zGDv2x0Av1ozMKH640QBmlR/Pdq0pFzQLBWyVH7UN3hInxLep4WNeMNVw722+
JnzmqQbrkXxPRpuWGmvWV8XmiDXL0dCNBXXLdGz+wMXAFMSdLnMwpEMPAUAsV03pfjUAV8Doz9Bc
LuWt0svdQufpiL6ayhYneLfgdGUnI2dTZpN3YExNcQJ9uzbOOUTd88Kcaec+3kNupqw2UaiquFNh
GQjwTNm7WkFqvaXcE3QPi5M8mkAEHI3Sxg4ZexIXhe3w+mjL6E7Hb6IeEPKIlLp7i8G6ibr+XE1y
p7YexwC5nhhxGKiL1x5xSmx/QHSjdj6ZK2OwEySUunLSblCnaeMeGjNQznev8ngo+7AWhCfeg5Yi
QgWsv1EfA3WYCTcEl8tRv5COFLjwgYNpJikmJoX0uA74cEcMC3tTSo3GOtQwCKaFU/cIo/ncOSem
o5IHOgudR7G3RaiMy1yJqJmGaHs3jNqrUQJnTiI9E6rSo0crJK+SSf9vt7KSinhVS1riYAcFoogC
AatiaA1OQ2ukbKfXbjGu5IFcvx8hSyok2CXPUX/CinuE3blqpzujGYYJgd2FSOIvkelKjeA1T3aH
Z6bkvKwEFjjb668gy3TupmOnAKc+Fufqr41LR5WRc1Na5UpmlI9cygwcIwYte/+HGRhqUhZ2hSaY
F4OiRQEqfFiFVkJi6OvXN+DQ4M0/20RF7CekICnsN//vMXkMpTC+6mbqmh5mrqj19eTHXf+Yfpjf
2n69D2geTgp9ZURYpGiN6zVaXfa2r+J1P+tsB2KXy/i+lbYKylYeG0KSYsj+F0mDgCbEez9FRrA6
Fq7Prz+do+kWpRPxtVi1NySF149Ul3m8Az8ddU/Q7K9lI0+KTPyEIDdWSf8KNnf0VLaD6OhlGLId
+YrAR1KcnilE+j9dtFZIYQXg/+2u82lkR3eBilVOOygvza49LUzjsS8sMw0b/l35JO4HPzYYbxuH
eEPJjh+Wy3Q4EUvmlhxWAlBGwMoWAzi4/DllRTz+poqd/iX5tbGbALUmWHY8CeVla0iYnDBY66fw
gWV+/Qr7BLbqZBRg0zgqNxx4Lclzfxkp6K/QWcWX+y/zV9pMgjihd4IukhyTFauJHgYupB+epdOx
cxZk7OJF/VD8kFO23Mp1UPEnKVLljX1mORTjEqtvL247xv6wR0jTVYD9azgI63UZDCbyozndZk8B
zAUHQtfyRz78sPbIMIHwDiMaB4PLt19Seh2c8Mp35Ar6wpybeKJ7W9ro4BCU4g1zKqqWAQ57NEYI
hOmUknnfRi4/VGL1wV3ng/Uruzbu8p9dhI/Gjtt7LQxi990wi+A27SGEQwI3JmhloxDzhrQ6SzLV
1Gf4OvRZyNiUPMlOFJAwkl1BdMXKsM+kopGuLBNwlEvxlssmxwIHF7TAohCK5/1dk6LGf2Bqwq6v
utN2UnVfrmfEakyHyuunVkO9MIW6nvXOjaoZ7XTYy5RtmgMFAvRZ+RxeoHjt8lWHXOIFI3KZdRuo
b4wrRR63y6q3e78yxtNtuGKD3IqmGIWNZJFCT6RaIZntm3SlQWVx/pyjI3o5gm8w5GzdSZzK0zWp
xrWpC6v0PWj+ytzBGK9WHthvPckaKl8j0anOkdZbTIrFPBpDW+mTAsficyfseCf1w5JAkMlcVgrO
X4ehCYhvfDQnsDMZ4NP/3r1cw3JTr53RsFwEY9aSuVyD6pOLOQpnGRQyRk1ejTo/EFMGE28/J/6a
vloff5bIQzO1r6TQQW7ZL88kOcSjJMsyeUqa7iC5EfC4lG9VV3HuoGYpmRHQUTaxtcrtwOz5i6Ih
x+XbjWQO/cSOBM1484XZcAd5Qii70Kwn+xe42bpB6TFYW3tDE5srCAvwo2gquXQyZoUpnsGD64XQ
aW26tQwCcZMxXSgZj/G/Qff3RQXkCaLtJ0A4GYXvIdDPWL1qN+p5nxSsx1pBwyDsX8GMYyutusEG
OhnVzz0ukTeIeUwLZNz1v1a8Mjs1T22i3hJJZn6Db7WRFBwNb7LgctvfjOY5daONm/e4IvGrxfwe
E+hPOCjRE9f+tCeSD8xOQO4QI2ECbDNw3Ds9IiTXkwm6MSYuvYon+G1mrVLR0bUMixp5lm4+gmLT
J6fBHR9PAO3wGRnFEjvJ/wmgVO+E5akXbAL3t/aQ52s0eSm9nFhhtNHgq1mcDa0q/igoZvHZracv
zaRfuzWWqOKuwsCmEo8P466+e6R8oBEUBx11qCSiiu98gVjCSiCbBMrCP/g/RHORv2HuAKgH0c+t
CnAhACfvmsduISP0fCFZTIGZcwe9P81fspTbQu958hqVFX2w+c2Zkcm574+vkoyu2Cils3831V8i
m5tWoERu88UGpZUTMAvY8sSwfzRtuywBQao5p5ZR4X+0i54B0ot/YCCWY5QaQpoXBecNk+B/4L9A
AVsbC0CrKXEocgTOMhCgPwY2shy1LV2Jg5zzt1OJ+igOcfJLbIoxzgDaUBKinzcbatzRtfnMFvFu
QVWzG5jZKsm80ij73yVCxZJT9MNap6F/2dFiDgwP5h6x/wzBPG5grvuAj2LreV/+wGBkrq5D80nL
rtGB3XEdHCG5KI3vQVlF0X1iJKIHIGJbJD436De02lRdH1P4Bo2OhuutioGPF/kTxPW8GeLoud2X
s1RGCg6yshU1vMhBBfgFfvOu1n2SvQz6zYUgavvCoMDxQ0b4/gGC8/QAdVQkVhfuFtcyq3+Kgsmj
fiY7R46SDpj8Xlk2ilW5oaNV4TWMJmNAlRKFxHPGQTxjbgOlzjjKn8YZkNiVDe4YHFLljyPNKiib
rQknKsAwfmqNWD/f/h1+iV2jQKozI4QGPDhLvHIBNsOIJslSFe8Pa49a+NGgQkkwJmrXNH0O3BC1
eLXyGcGukWj88gDxSUzVEI+J+L1NZhBCQVx0mv+HE3iK5NiRLkf+w+YG0O4BWZfglehmQTo5xJwI
FzEZEtrjq6w995php409bH1wfaGvgOIJ5ruZGJfQPyvpiy2YZjKiCTBcFhF15CvX08878Ao5WCuW
Bg3L8eHWRWDvPtCDVZ8QCpzqjsG0gPkFqUvEkNtO5PnAq9C9r4798cN//zPqq+RB1WdqYmIZy6rA
XDHN4VxFaIC3LlWQckNH1DuvighzipCBK0qKpKnIs2UM/KhYRdUFtX97d1zV5UlZJCeqkPA3P8fQ
EL7Ekn/sSvJLfg9hda+TKgHAmkD9RMSeQTT060FAjdGXMwRzLkuhnsa47WTZwY8rCtKfKiyNMdmT
vkeBUAVxofScPAtLj5VBFp7OSTv3T8GRgpLQgBCDI5Zpv32IYQqtWtIiKu7b+91xVMCJgLa/T5Z8
iyC2mWLC6La1sLPNBeSCVTB326Uw/NIvpHeVDlsPm609EcFT1cjjCHh6i+XdR2ZKyjTLlGexxn5M
blvB3KqrKCd0WFjCwAfkJMWJEpKR/8W/AOPR9bbByvzKruG4wHRe5346x/OTqgaj0WhK5ACrntFZ
iui/THw4JITSN3AZhTFrmXuR4CeW6oEdJ1mUlrt2FxVzacncNOIc9RtbGsEvGk0CU1zBi1plv/zf
f+hj/jJ1vhcd5I3jXqms6oEsKfTiwJaQR1m8CDrmepc28/gD7W3eOJDT3O69QTB29GpcmLwWVUQ/
TVgQ3TOzVEp/14OcMlvglhwvxqDpq2ax5ccru1/3vKDYYtMI/BOvKHrYRt7ONXU0ouE6uV01aSxl
1I+OH9lMLYFsVvIjKe37xNiOTifUQv4eGHgQiZupE/0EPlxgCoCU4cVlAyDXdo3wDA7H91s9i/l2
Kds8oNN7/xwywZJFp7ry0B65nhfK3wt5vXe5pyGtsy5yxgEKbsv7A6Ii+k2wHYl2Lcu3FnYf0bRR
b/xu0GX/eGhWv5rNiFtHUlA3s1c2jOIjD5iPojms1LEOSd2HwaGDt1MEWM80UT25JUr2rUJ75LHQ
NnMcnTdPPRHqZs0WKxTtvu3omEWSl9IDIzxJ4m7H3Qv/q28o7nX6gLZ+x+vEgMu/or2Vjmm+01Uo
I7QCOiQnk9feUTFMHDs14W6NoFdWZQkMuF8QxjWq3i9+5TLyEdZMJI3uhKv9qacbL/lc9MZJgU9c
EawmRaSZOWNB21oluIftMz7GQdwFUy6z0ZyxHfxigRSeNHR2deyJJiWFC6qMD8CggTPdHjMwoBUd
miPBP3X9DGMXYx0VPubedX5HlhcD1OWZRZXyzCpqNuJsD8hD24gYsolKz/AUdM/9T7lZleD5+CVe
p0F9W7jDd9In9Cbjan5KEhMX6xSJKCzPQZz8o0q33RYDZ/RLcqQAdwZkF412dilqv3osqjyBfiVv
jMXxWMvw7Es9CK9yQR+4kdPTrDM+JuD2euDnketCqJr0+KIHhPNG9eqdUrlNY8mvtLRF1nOjLdg4
I1UI2Ir/tfLnHH3hq1x5L9baomUhqUiP/I7MxfyzhnEG45HLZuzqBnbGiIikI6hZhBA1h7gtk/++
ciEsQjGFggiYLFpOI/PUegSqOplzKuU8QxD0dSZ2QjMBpTRwUXAvIs7HgK1Fj8PcL1rTkxueZB5a
IjeQwMEeJiJcWrT65/O2qg+6tpXODj28coxF6RWZu4/TnuHXWX+i/zwa7d0uxqTfnK9nCa2bAfda
AU5ng9Wa9Jj7OAC125TGu8PJGBDbaGNUvTG1/PEdKZUaWxAo2MJugqA8vlhSh0vGXzaqcrXIbVa2
MfcoqnLOr107gCpPswj88wY0lQs2ZYrO2RrkdQ9l/V5rcti9s8Mafs1CYG8TYDs4X6INAsIAqHVL
BYPEdr/Q2issAjaAtmnUhE80AwM+91H2yx5UHWjboc3/vdszk1UUQ10W7OhDr6691I92ce5LcuR5
BlKKQd5COEe8siFpCSR4dTQ/gyeFR/GxYutG9VliPOYVynfKGc8Qk37xvnEvs5QA2iNud6GBHO8+
mfJZzY5ob/a6VUzw4+fhhFFnyWJRcLPuldNpnzcR5OgqzCkDGXqakq73K2ZfuI+Tt7hlfSXG/Yvr
Wf2sQiWuTr1FPQwgAT3oj7tjk5WRLBumkoBjB2v1QbRGiKq3+hMGCIuJsXOWsM/OjMQHy82mKQFd
rg4lHo0RymUovnjcgoVlUC1ODwYH2RXJeuS/Lg70O3UvMMcXF/ICp0IgFkqqftXQrdsaOuIEevdf
v7VIjhUnGC/QlSx+YaDrVZahvHLOpfn2rCmTTsKVKhAtBpidIJQ/fuSkL8kxIl5PODPdlGBlJlT3
4yQfjEmOAwjIYoEonsFlnBVl4/G2e1GRaMmVrg4G3n5p5m/ndCwa82Ep1ohKXdRsaY5befjDkjMN
utwieFAIEHX8xwJJmoN3gAlEWuWLKVpfLCuTupa1i/4DLu4y9di/mcg9esSzUvlzLbhlL/q18uVe
hO+19MPQUgMZdRX0zOU++NfFYziSzQYruL4kaVRKsFvLnwC62B9djYAQR0TDf+NRHNK6ckY8yWdx
AKuLiCJmWQIxgVjvhPF1kgHU4IbJSjzN0g0atqxAsgN/U5CSzipDZy6+EiwYfBUOeXcuzTTFZ93W
Q/fHcX5dFvamD1JaRfMKlSDMX3pd3dn1LsAtaL41mIAnBG9/4AEmLD/V4mApgpZaM+TW56w+KgYu
pjdhSfTvh7R7t2P8frf7fDhN7wkH0dcv1CRFFd/N4Ay21lissuqw8Tq5OUIdxsGL5W7NoJPnMp2E
HypN6jVZ+NQYzoT/GQWU6gvCHhLFL48B/OZ0/5aQHttrySmJ9ifVJ6DolC9UL63g+ZH2LPd07eKu
VJdr5fhjKbPHVnoZ560PglskcsMoahMWASL38iQS9MmOHoN5gaA29z4nIOZt1O1ieXJ47+hnPgqh
LdF9yqXrsX/cxxCNRBbj1t50PefTQAM7UlB78KweBYzVBsKpD5rA9nmJu1XyceIVGIZ3CqSqlEhg
0aqDtyvhUyy68ek7fr8b63EN73ipgltrqo/qt7JEC9qDl2wNBZqnxsOeG6z8J6zBEyJPRdX+pBks
9SK5+BEzz8i7EQPH0PYc41XD8JR1ejKKK+y/RPBCCPq2OjkLE+w67/h6PYQ7CBp6JEBEKBSW5i/d
Rg0mBBGAmtJNN6MQMM38Sz2MOeoJF1VivUaqeDK4tgzCrfieBBn8BxefjaozFbJP2g0AoWUIoa2N
ytM1HQcZ0lmyNIP6ggL4QjPV+Nv5UaaXOk+S31fySJUtTFtgYOvt/gvRcEV5CH8XPbRGWLpX43Fe
hUwbvb6pWeJkx70UlkGwv4b8/bxsl9XmdMSiX/MTDF5XjZgkCxN5iZ4oH1/bxeqQmDhwEF2j8+dP
wLw5/abdXEjxt0WrgQOqM9MwYObKv2waRuz4PkkQcowIy3mNRBurejLHuu5/LRR5OpWYxjyylpwb
fWu0Mb5NG6NXsaiDxJksgG3n+BYW7AjrDF7ayLNm0P+uUT/4IkwwVkkAROWNBLuVBtuWyd66YZHM
Ix41ZuoUmlEg1GCpsN4Vve3T8YmGWeAlmifclZZJWfm9tR1aQwA8j0g7Erd+cX42getF9+vA2s8+
dUUz83WtpfQ/oKWL3lBN02o20TSeaJI75EjnY5KrgvDoIZFx81bAlO4fjaRqcO6nVvwilh9KgBAD
eNOfRqqQ4ZOgkSfibtvA/cAOGGS/+lCW8Hvw+CgUmOp1drrimLas3pK7oThQKNGV1+KkkviPXKJw
s4a/Ntuqs7wh9PzfRy3XKL1NxoHwl/9u4jwUdTk621yKlfBLXFbK+SEZEL3vjiFsUkEwZG+ry5Dp
TXAlzTHaXmWVCOJP67gI+5J7KQE0/PvNseV2W6Jnp0a66ihrTUYTjQ61Gd2U64ybANI4SaFCNlm/
1oT+hO4Vt5BRrOpWXryj74woQNITjRXoi4/yUZqKrO07MIN79X8UYrjpntEg6BABuC+sMdmqFbGV
dxMiGY2MMSV6Tx8+HQe5pFD4ryT4ClqC8aOcloZs+TL9faGBN2pQ/PyJesytz0WrOcBVrE30twuO
Qj5EGuc7E736U5cHRc6PKvtPB47WH9kp9Jm9Pc54ha4xY6nN2ku6UN+2PFAWJxfeiFlp1BKio/bx
m2rJlLYgRbm7oofmifOVYpebXZ9mHtGhGGTeygdIkY8X1stkLzFqIHdxeJfw9t7SUb+HPns1ip9O
fRL2kVIE6/LeAPH5NZkHGMeSgnTeeag6DlnidHf/HZmpQ3EReWB06bVQtUpURc90qZt+sQ88BQHI
tWjxz5/CQzPjjn+FcOUkoNH7V1ru5SgFsViL0XW4xIBDvkZjXDGbor9aBaD+okPOPbLb+PGB33z7
GhRM0yIu3LcdyAFGFFrDNzKzdpkaCKiXLNWPqseOEdIn70cM0K13cPGfn9M+CXAcu/o/4j+VzT91
HKQe2SQbjkGVzWoumePeaNb9t/lYrFs1zcU3DFfBu7ffEV1ycgGh9LqQrKfU91K9/gfxW/eAUxaq
SascBMue3Buj1RQhfeIOOzG35bJft+booX6D0Hgaa0utQVxPysvxBro7awFOfzE/h3d8iwXm0mkY
tLmzt8quLgjQPpz50g8eqaHkAjvnNZR+OMjQG47+y951UVC8smPD3WdI5WHZaWlWBvcY2k0q2BVr
fkeREhcu8qA87CXAiDTW49cpCR2NUqu/R3fAwVjSqIJFWo1JhTx8JXDOPyoHqaerDJDp6v6Zq/OS
OnnRF/VEXuga5b5r2fcjzz5FxW4aesMg+nt43BlR5xKkkaH/Z4ZA+F/nrFT1O4mOkTid4GlT2CTE
NWfkSsPkJeWoeyq9P+a9By2fQuHgBsTRvJqT8UvMG4pgvhAB9JQ0YuFh+wUeFoRisMruu6t+gkWe
WOn5F85z7VL6NW6KRmPHxT2m9xi9pIZ+fFmwHkb6iT3+Wv92XiRc8Q2TfBrY/zpG4dnaiq0m8DSH
6NFyIY2yt+5wjG/e3TH4frJvzv6aQdrvJkRwMANdURXwwWta2kkPiEXCbLI6wleLfcxe/ohWniby
sPPHKyO906a+NWl3kv9S071o80xICKgUtXyQREXEuzkiu6cizyDAs14lOFZRhEXvjHT+Mh7a29ZD
tiFwjSx7RnoYn08ldsZWP8jCt8hzy3DZbvGQBrLTEpqLUb6AmYl9ZRrltY6eYfCG6m72sQzidPTx
Cd/dXVf5qaCFttCzjA17WV6B7XZ5ht+slzOsJ711i7wOmzfQYyV6TRzkkpGjMpjcgKKyefQDYGjm
/1mLIy4ngoQ6XJZ/EHDpe7/Fb4zGkn2cc/BnZS1PbQ7ORT4YrctJ7XDhvNceY7F1Ch4W3tXL7xly
0R+3loyyPkVceHe9tE1J56zg9aSdtMsiXZVs8mcemZkxUquZ+OnXJoKpy5zuNOiUdCLR3CkDw20t
8WOmj6ySBHD4mx6c0tbOzC5qEfLOgaMcgumvc5IGjVwI9lLpcJCjjGgmzg6k6ADWcXY6lJ5gVSX0
cjPb01E+cI8YPmU37i3/PesGozkytcDzK4QJP7Mi/Q04u61DfpHZ9+nG5GVlbw3ZzjqAcopkFgOY
FlpVpTNRT4VLH83O9LnnBYIu2+0HN60mFP7hH7V37VcjgXGzu4BtvBAD2Xe7DIw9vRCZAXxi4Uhe
AXT8BrC1al0UN1c8qg9Vx3XdSCWwo9V0m8k/1OpntFnKL19bdIuS17EgPmgidSNLDVwdQJLW+ghm
q2A0TNaIp/weVORjk08erNfi3YPEYF8V9vVLl0eDc0N5KyRmTb6ZyGl+h07IYAH0QPzA8N+ZovSU
RBCOclKC8mMLXqEEiSZGhv7Av77wkwOwPs6jNmfx0QYaT4408R7vakXfaDHb2PF9J1A1jn0QCKqi
49fkmjc0u7HE1XzCBJFGjKoNarDqmnoDpC7E5F/17LGPQRvX26vkWMbpuGr1kNEr4i9oNIyHxndO
kKzhKZXIxoldVtrz1wZ19uIJF7meq4j9b71MBNgs5FxJb+hiM24JNAY0OQDmc+Mz391Os2yPxl6p
H+RgmMOauZHbat42Pqfa6WWjmfeepg/mceuZpQsF0XAI3SWlTvk/YsJTMmIfBrm4g2LKf+ZeIzeE
t0gRaNPTrhS/8jfsYl8NBGa/MSgmo5y2D3+m1Fi/D86YaO2eQINnTpoqQiR/ReX1YoMMaXBTXJ3r
y/uxZDkyUClUp5XiiDkV6O7efgNC90FmvWJxATMLDIcTAt4xif64Q6p29z3HVzLHmUxDadyNkD37
vbuCI5bp7Cr5L58gxd6bq237eTfFR3/smRS9w3ShVZY7fCim66/2mCXfc024prwIYbeUoUCx7DG3
tAIOspaq5hLbw3YNe4mOTv91C6lBAr5E5qKj48yBDB54zaVb3pWMlvLys3XKSG4AmwqTEEgk1ymQ
23xJBKZ5UVX7FF2Hos2O0O/CK1NWNiTgzFMWRoaKNJ3P9zIkEOIo6IBAG5r294ru5Uybg+TKnS54
eT/9Z9zsMdcJcnx/RK1EWeluceTGzYTMSO4xmwC4+TRUR6T0R+CVfcFzGdoVgdfe9AB0wjwaNSlu
omoNjnUmskjNuvbLB2P2EbuOIPe5d3mS37OgO93lv1Yc1FJEoYhAz5SkXUT3WmyAvb/BzA3L+2AO
Xpg+plzHs4ZzoaBD+sGBGW5BEGCjXv9Ig09F90rHIQ5nz20DomJCi6HziS43/P9DrOsiqUKJ1PCJ
OoBt09BpPd0MYwu/4Uv9I/wfOjf61y/v7XzbgW7q39nVr5ajbs9V5C8k97qq1T2TM7mPP+yCG7ft
VXIc8jYFNfbQcBiIwLxrcOpZQ14WdeIbzWjapxRCHVxrw6r1yFbs/5/qM1lj7e/f9cIleWeroxU5
gKBBnx5fNtpjsNHvpxyKuTfhWjADC5YqHI+cdrIaWo7jM5r+feCfo/qXLVlDKnDB04fOlchtgab3
PJYfPs8KnH2LSQMCqmQqigv8+cXn2NV7bHJmcPli5MQE+ESP0mqP6sHGbrCoYHX9ROJXNgXLvR5h
3362dzuatZUgC0Gzvsr4G2MIWnjxtbtGbca4ir9/A13a/lsRzmetw5x9E3r83VXmfQs0uL4drmm9
vKlGruDOb2IzYQgHDUiEwk3xsJBRPm00u5fNMKaN7S3rDspveyZrJLrmNgOkCmr8ulyHLycZPrfF
Hg5j0Jt28urTxYn+YiofKG02Bibaqpa/5+Tn4Wcns9UAhdll/HYmpnVZtZrLyaYzOIWTVa/CyWMV
a2QEJZWIpaYfzF88ek/Lii/OwSGevk8GuSW7ntAeu3O3h9iZC13t+oW/xMB1u3xJ7OPef8RfoN0K
t4YYJjhhPlhKaNFZ6JpmsKivq4lB2GZpofWHUd0mFOESLA4tG1aKCnMMjMl+uIi+Csn8rL6UNr9X
llUwLoF9l2T0bbkU2wk9LtoXLUlcoBczouniOhh6QXGkP8O/U9cCuSyjhaY+Uf2wxK2ksNEFoBPk
n7RNlVWjarQ6kMWlhmM3mUFTe0V9H80RkQjnX1rwPP19fgLAytuYZbcvhBfqzJV2tZhd+l+CDGJM
5L2wP97FejmezYp0oxHji+goJhgh7R8tksqd0SZWw33dfLG0o3YoIgL7TcR8LU8T1Su1syEtV+Iu
k/dqVR/BSyJmL3lkpMRMTLWMe6I1cdtiY/we9cpbxp3lAh4r4oYBDeXK0xDyn7T0EsTxkVoCZjIG
zuGZSX5hSkSoZzdSGQ8h2/Lw/XzEmhjBTWbtB3Om8tlCiyhrnV2CILo6PiUdfVf2xSPLMiqI2Wr7
EvoWS5/bpI8BGXMLEghdBJdCVV3ImDmnaPDJuvAC2KRqN0GrVNnDUMb9aQVuRXQdUv0g2Iivo9WR
wsMN8butXxrNxR9w3NzH4W5XKAqRxCWYFpVgO95cJNkczk7ojtEUrmwmsyy0Jl9PlkL2IVqCKyYG
ODGMjdE3xNCC7zm0yRTq7yLSOmKUb/HCDRTeH7SKdTxZVljBN6MMgFcQH/3z1nCk1sEeoQzd1Imo
sLsrdxyymaSHJx3bOjd7UJDe6wc8+aE+9TVchJ1w93KfRhIlqZY2W9ipnYJgLvVcY8hftCGJ8qn8
SCqDc0tddxdDKlsV/SwWPrHtVNXuoT7vlTRdjuLLHr+cOD2b4UR2t5Dt5w2KsFiDxKN0ZKnvZ+KZ
AJlqwvUulgZ5ubl4JWuhoDTNnoWbgi6IbjbdrKrKvY7he9JYl7bRYZQJEkAdeVbMoVQiibsxTkR6
XPzc4GX13sDJ35nSfgyDIQjKkQAhlFyJdPgLmK3q76wGdexT4m5t+QwScz/BiG48zCiI/oLbZm+M
gJxouIv+poCup8q1mReVgvFgOl2GVD2DGUuOzdRfwsrs6Q8eQYy3BaRcxUwDrWUwEOLGPVPdTPEg
Jg0k6RvP0cuPjL/Jty23xm0/Bxow1poUfJr107qX3zzF84nYxEthwipgtG15VQYvOwciffgryG2T
jfiYl0DwZV5KOGx7Bf0IkY63w6qY1cA2hMqOLEVzwP4uBFvPfGLwTy88SxBxcsUtCkIQh4hvD1ae
37YGAReypxl8fMgzTLYmymxvOpvDEb8tHQ2z9IjRExlzoq95gTJEtJlotElj/e5SJibGPtPtsf7C
rbvAQJsylaYS8Q2fIjOVA4emPzH516oKJg33/2GBjC8zMKuvhmPNWcMNdIR7/tlj1KS/ng/JY7oB
8IHi1aFHZGo7ZV9Ystj/Xzj4CrfL8C4RSPltMVH7b8T98i4yCmJHMXAQXxabx+1VZ6KcaA2ziXSg
Drf1WmaZDyujUilFAryi12dUAs1vzvN60vxZBipd866jgUXDfEXa2nGt0potvbwNNx8Nsgzn50NQ
az7CpCM+ot0tylJHZdnUXnXmLM1t/3P6q2fI6VqXbKvdkAoRgIZhQcq66mHy9WKI362Nbg9WYJQc
/TkEmgeZLbTISx6jpaR1yNof6Q5HNZtBJ3TKYKE19wajshhJWbMcw2UWsYkdIkJIZgxjVyFLbEnf
hbW6K9Xb6gdw/V0eyQCetYMtZfl6bw+KYyJhWPjxgV7CAF5sf/xyEN9QDd/Gb/32nnKA3AMyNag4
QcS4MD9v1UnDILTxBRj6eiZRmNbuisZmBgNVTH/I8nEqH/OHuCr9ms63Zt+/uOm4p9LZJ/HIpRJ2
PeB8RO5+pcoEhWbJkd5SONeyQXEpmgIhDCgikCErKAV7v0jfFuvCBVnV925C6T0BDwKQ2OxT8EOw
mKt0tO1bRCtkP1YzbeC/Lb1mQCQIlMYeTYYq5dkGQoolepjENamrT0gleOj6m9XQKpZhhO64Q1+2
NBlVoHeCAWfhulfPG+/T6XKix9w35O3FY2mw1xhR3V/+FJTLuh0ozFjjfbsrer1lL19B3v2Wok4E
V0edfYvPkrcx9dG/rknZnS9HKD2dtQDZpqAxu8Ju/XpswjxdGNMKF4IrSqGVdgkJBZ96/I6mTkh9
vO0TYkCVPmlIvVlyt/TO+sqaO1TScnGUZ95jGPfHtJItYeDA8wvC8gLS0kb+oRUXFJUvQvUnPYFX
UzdR249gbjJ6wBKoo7CJWzQMmKo2+ipSm1Soz8fIWmKYOnpN/UcnfycQZBA0q0kFlAnYRbmeU0wG
g/V/78fAJvo1ReL49F0XUmPkZUDb44EDnG5sUMrtpwObASBm3sQAWKqxYuOVrwZVAgrAFTG78gfN
Z9OYWVZLz5N8q3NZqEcEajqe1hyOvB2CN/2OhJ5sUKBI5Y0yiNbCh4bkEcdDbZEF0CDCA7WLhspo
rU5Ofhf2PYIkRHNwDDGRSAeQyY8zsde6hdCrIt0zOZsqkFFYNfiOwlr0xVo6B2yn1ZKVK+RT7HKj
gPCBefjv5Y5A5+cN6KOmADWzDTwJMhz08nWOmaOZfoHZAasA500BOmf/2VMO75990IUPjVZkVk5w
3e3lf9+lGoKJneNppcbQV2z3oMybU5s56cwzFKk4LVzDZieY+z+RF/3RXLDsipTmFzY5uBnIDbSU
FjhCr6zuaBk98yKXdtP+xEP1C0wgfx4GoBAMSB+lGIzbscTSDliuVqN0ghvTSwhwWVWSFKAfKxly
1euII2brcDjKZ3WLrcI89NniURpx4YUeLX3IgkAI3GWX3PZlYY1vG1hbTde86ZUcVrfxe3mqdSNZ
fo6BjWwkKhJUSR78u+Xv8tQNeMlDA64O+EdAinJwzKWHHKoSbFvU77BaVQ9rw5ioY5GXwWPO2vrZ
LQBb/nrhFjaw2YEjp4gVRoRGAYgApIrfMmKCMi3kv0px6jvoEbuWY0HQGzqYSv6R9Su5vzkh8JEY
3jXD/q37BxthF+Rrf4jEH7lisCHVIPV4i1PSmtp7eYj/KVes0YEkqQgw8dXK4E1boRDz5gMEoYyC
wSZNmsXALZDloM+MjQJXe8dT+6GevuiSE+6DezrqXFamf//A3eyEmKJDFTPgaNvJmqAVoz6CxXXt
pKpV/IEfMe4q+9WiVtHa0CP4yxLxT3fIQNH/SCW3vT9o3Aiq3DWMHz2p6Ebru61Z6BIvyP8DVOHL
dkn/43LQNSDQiin31cyqGFSzgJjdkXT4G95UA8kog8BZnJMxmntmgmb9eqCaUTmXf+JKWUQ/XQPI
iaabg+CEbjALuu7kKJ1d3n5NfcJz4wVg3bVzSH7QXhu2Kbp822f6FW1pN5kHrtNtqXJxe6cIoTSB
KtlFjb7HsdCD6Wh1SaZg0r4+p1fSzDv6F9aIgoHE7aT8J7gAcjcoJLa4byqjXM0i9swBLhLeqcrc
HamZy/opJAulfIEwoYvx3WRmgW2T6q1+lglHckU+e8RxKlWVeWKsjZINcMu6rIqOK3XjT2nUNs9r
W/U9OBLlIqKLD0UIJR98T+GmKW/Ns6UrIiB9/gfJz75CVf9P8RVH9RnMM2nerlhIPcT1ehLwMtS6
4564CNd1WIYBAHdyJokMytSQGWlS4bjHzo1R2xoKrEF3gKFxGVCqiBwiKMW2lVpJHk5JnTSOElbg
duHRtbgeVzQver+LgHQI4DU1vUVYQ2AuOpSnp3jljQxChk26jApGaLFzDYQpWaN3DbGzpODh6dM3
eVDOYxCNcrJaXqPfBSeAaeCcShFofo0zWetgnEf3mNOWEx8r5b+793dXkpu183ZZyySGleaZ4iKE
liKPvNqhZUHSZ81UTZHjFZPa5ii4tYr300/zfEOtZvUqbQ3PLX7c3dEJYu1LmSmanTs21FLa8dFX
1jZR9k3c72NAwGTcmb+XMowMKWjtgMaw5JasVol89N2w5m6PEOVwEe4AvNrjQDuk+dHGZam6tgCY
VbKCYS7/0So7w9FHwGfA6LvyjRU42ASjE63C62fhzfd4WVyHrMom+xn6C1mltllfR7ydqD+Z00hK
zeWuomHgYnCUe0krjU+ZmnzRl5UFU38yZoIDKl3FJygIwh1Z0847E9jJCsm5TvO374WPZ2ZSVjgq
RUYWzfH8xhGVL5X2nl9T8jXy/oxxxcWGYdQPF+WQ2Yg1JBzyEH8Pnbn9o0jm7Cg3FsGkZtCS2gtt
detRLnyjN2dL0TGHentSbL/LeDjcZo1dJcKVwn4pX1VdPKFA1S24wG/6H38QcsYp6fCkCb1jz8Ml
laA+MNj8HlKS8noXMjK/eY89M/tdt2xE+ly7GzU/F+peZpDSSygfjhHSdp28yNNSGE8UcFKSA25C
Ukq1K5nL7q5JX6H8BDYQ2Ot3GOGSdKu2TQKvdDPMvG7q6JN1Unlc+Y2Kfjil0hU5hlKfREzLRYz8
11iGsH4XsUqHiSFzo+1j9KXBYlDGktwWRxKIHJwM4f7swIe6loApEbXqH5C6hRPQ/e/YJMfdzLQ4
fCtAN/Q8/znqetjEuhGQeuhccaPPqkQeRlZNuPWcIcmndcvRjQVdYwH5oZalSNofSDVE/+CEO+y/
wNTrXVuKLSy804whWXnRNh2G5XDU5XLEAxijhAQ1UTw0ZbbJtXAtQpU50YjNPbPcCVh0j5AIIJyh
6BClLM51ApxcL4eX3Sn1kNvFwna4f8/igdWyQlUKJM5FQzfcsuZIWtZo60JpeIBPgXcCmylNg3DE
r/W1Xk2ECPKhxT3BpRdUlbj3er8uZnZwQjpVHy0I/sjSy0vT+nLa75l/Hp8SfxTfU+cKNTT7FfRz
jENs6w5oqMU45/lPHei1xVa4IM0bZqcxC9FLH30UMcBSPrqN552tdkUXGJdoghnWd+2jf5LhqDDq
wOzQYquW5QCvACdb/N6hXZEA2V2woK9a71fAwVifL/Ynvovhhsccj8XohdGEZaB0olVDflColDDl
idkY3Q+XMSLZf27N9v2ryaMrFb10z5tPSIsS9VwCAN7NWwFBnd6ArJYdTCdjY4FrODZbbKNAAttB
BINIkg4MiDq6s95cvADmsb8kg5ZpLejtb3Uc4GSpxtCavg7lKePlYJEloy0B+Own7ZspJUnN068o
00nxfhTQX4ZYQ7aKW6CVIsI8oGhvJAIKwf0drZol64bvtQgsxFj82/ctg4ApfrAVUBLOG3VXogC3
V53WnF6H7nyG6C4ckQ12fmxrbsX0lhpazjcFLcxX5tfE+p4gt2BqHPRZE2zY/nEtTMF/vRXLBZzg
R+3Rqi2Z2kUxv3Q8vBhSMaRh/9kHZEFeKA/FR18wojnijpVEe27ew497Dz1m5dfZTGUZNUs6bqxE
k16167zzH7Xo102SV+2Jt3oHh9h7XriPjkh/mM/GcRR3lUTaYBt+lF2FFMh/qruzrhUxXcfRHbRg
E1j1DpPlo0azhC2KSz81CPerA3NvitVP3yihANCPSxJINRQvKn16KOKZpSilmegtVknch2Z+F78y
mPPQi7Ejc+ZtdvZ0YthnG2yULTNqbU1S+F6Zsp5JadTzeIIBXWM/oDhLkbUXWTda7Rjb5RFjx07w
6JlG+gwuBkzH0eG1sjRAYV4Iu29W+03CexF+S+1/dU87W4UH1MYNzq5rjvmIg/omQwWsbsXHAGMg
uuMzTQA6GO91jx6xphS2Kwqj/WfGY5OoA7wc0a8ZnI8hvyNP3wJS2qMR9EUmumkwntX9+8rYpLlL
AC30c7oXZrZEeKD66X2eN4PzxO8mFeKP3TwiKZ6cmy+FJ2gOOXF45duld6ix1Q35AASLsR80jHnK
8lnxpMu/3Kor1uf/s+usuzcZT9lwcqPjw1emmZjAvDextLi3eTIiDJHxd8qFhk5k7uj2pI38rEV0
OPVNZx6N9NR61GfVej41QqBdLiMRFDTWf3TyndUarb7qY7hsoH6rXiThnEtgj4/1TkbGK39DuRBH
XqForcrf+pI1iaoM3plRsHfe1kGLgUCBNVqZyHLvxdsJQ3nk5ML6PLwjVTCrCz8/Amz8Gf9Td5rc
BZNzPwHVh4Lu9+Osq1Eq28kec4pBdg4IVkvpbqScDXSgV0MQ92hE6m4BxclrDqMyFKC8Dh5oZ8xU
mMBdlBOg/NJ+5NU91eN9QQOdG9NUexwKGlXOSCj3xm0htViKhYQJO0/q3JvtKFf+/94k5ilXFx+u
CaKTnS8LwpojCQIBot2xnuwf7XqLwjY716HGEJJSajszKTbNkrkpx+0xCh5jPUCXP+Exco58r6Cz
rRWVY0gi0aQoDpinlcIMem0beSxaqqSMd/pUiCoAzCHt+G4P6ulM90TOvvBKZFy8aAXoyQ0gNaH8
fa+urYwQkpUHuBVg1U3DLxi3aI8zVgCKxe2HQc9sY87UaO+pUyPq0srp7LA0x5yLtqeahKHrAdF/
NM9KQfcgZ6PSakOQ7LzypgiNzqIqGEDdoNIWJMlX/OjKz62HHp4idQIpGsEKjHRNMaeG3mr4D2Xa
sLHReE6Z6+gHEIBFrgoVEhs8GxiZOe5nXxsv2DMpzfIwEI3+sCmBwq5sH8+t4mx+anInx04pIxu0
ZtcGydkxDmomU8RnQ78rOlAE+jqA9Al9d44+sqvYkEkvw9lGUKXwS2cX73MWWUdD8+01yQb/mu4A
aDLhw/XgoW4uUAWr9XCK0S/WfFqkDn71tMXK+XeQNkraSQKni0lLfUBXO8BHabqM2O8buhGU93/A
VmiYLQGiYemINS+EoRonbvOafd+doSHb2iGJhCCIwWl7seFCwdRpiSqivGn1jWjyirioB38ffMKX
nVqdHULl5DE5Y5PkJ1ZL1bguWkihwRdHc/2s45mmJmARUS2u2hEOsetNgrvJN4zAx94EZcPNCvW7
rDhpIJ7q2K9/dcKJViDbrqaDmnGja0O4aRdZLBi+08d22qILlIsmYBZdqK5hMVzicnOo5EVVSvA9
0MWsHptr05FJ0U3qW+yNovPcvw7fsC+yzrOQ7XzvWt//bpcmjKUWKXqEtKhzRZlT/HEjBX4nxWYA
qThqn1djbuk0uJBMHMQUeluLuDzUo6tEb15hsqsGPr8GWJkfB1Nm71Mszvd2OHKkzkosyqFgLj9t
3K1FaTA0c0T43hUVVrodZPHfWE7bXFF+xlHsDWM+46dBAmKek/5fgWiXR5EjGUN0HQd2Jx3RRwWj
+5qHViTdBPhhAyRvowXoW6fdIKoWjfIK2CZwLc1LZEnUV2IKTyHdQZoiXUIJlsuHDSs+EfiPybW6
2BxTQQl/VhbDmYYYSI6VrzHEHVlMe1tEQOD7KaKyhDhStXaUaKCgRIRrmOtq9/wgBEXijZ9JX+OP
0yNHOnP9d5Vt8hYD2lrehg6GkcZX6oWnVdZWM038EPAY6m8w2Kfv4ABTbsTQo3joA4+AVSbrsHU6
ewu+IV8kBnm5ZaFEjABs9tgroEk8+6oA0lfAgFh47gTnAcHMFS3WzeJpN/neiun3kmt6pZpDyJxc
MVpq8fIek5WBnuPVrT8tEe0h4Of0ZEn7feKmcCNLtNXSiSwo4TSZC7BaXNTXRj+iUc8a0hQ/c4yz
xK6lE22RitpKfrDtz/MmLaZbijFaabXMTuZxfkfNvHUzdN6V974b0oDt0yuvQ/AusjEdEbScO2+6
ET1xDw+0+PCjWugPlehCyNKox/aPXWepXxTAgc/a/A3iB60HS9qiD9/hm1BNYuKEUJdcEWK8yqOK
VFQDycTOkaf7nKAk/lBcC2iXc4yEeGD0HSTvuf6OCb0F0fGCtEBgJsYj7NZBq/BvcmDj238q+MBG
Ac7w7Konzv+KmAEb05DDjjK6oQeVgJ5VOp6/TgPGcYhyCHV1hMmAwQcgQJmA95CuQUAKTiNruk1f
gu1gmgRHftHM/uOdWp3iD6AB4Zfimj1NLG7OobA9ibfY215XQSHASc3XACXnmRAZk+xqVxP+8F2I
l2kHfUuDmx3MTKH6pqFcHtS8il86md3wNn7eFqssSv7KFpcaBA4a/aiBWRnhGlRnNps6Cbiu/jxM
lskO0c2WducJPmq7pdz+wmeYX0qdqwXnHrt2FawQM1O5wN+ERicNNrN9D4tTIIwukoMIQf2NHZgg
mo+/5PYbGqy41USrWSY097Bsril6kWNc5oHJYYy4JHGU1x3mc5wLFUWe4JjuSduD1AUHc9Ok+JYa
xRWhom45QXYkSd3/swMBdShKcvww0kAT4pIITVgqryikgsFH7/B0ueLkGOi2DZxHtdAwJRGsN7DL
6Gb0KweyOgVHZQYUHgDhY7jImHslhREIeTgYLvtQTD+jtgRRISji/kPNqMx8w0apIDPt8Dv67MSK
1NFAgL4OBcQAr2/YPQMfYVWKlNoh10gssfPH1amVfvb1TaJU7IexN5qYcHzXDCrKEcqqU7o6FgGl
uIen4iSC1kqS8r5P4Ig02DZcIkqQngcwzJ4uEUcpaE8kRyAhz2fa/SNBWOCmERrODfs7h8+UpL3f
rE6QwOiJajqH+ISVKUzZnFI+m3B4XaaxIvP9BynjRoNfkqXUjrUc+UO7zWAd9dGq9LekaIfmJz2c
+vwcrYfDoScmliLUf1tvilDGW71k+N6rVdkXsVJdSmkXP3GBxOFYKsVeKM+M4V5IXCKDcnaiqVHG
GlCxVgIJEmhZqs3E/0yGyKUIECYitsUmG3vzvRVNaRcVJlb5QVWcnpRmNn/abVKkYYRga17mA8zV
8wwyPsESybvgMHNTExhjwdhluq614mSMxNA9/MaIwPcevP4X3oS/F2m0+XbsWVrOfNGC9H/iOdaW
NrnSZB5wVmpb+2muJY0Kbd3SRC1JRUGlSJTWjIIfLpgnsS1kVYJZCLBApNHG2cIN9GHzBUAJqdhs
MZPOU3J8WKBDAEBdpdhel0GvqZof2WaBn6ef+iHqpuejcO8fBkVZBxjpExvf151i87EJm60Gqfh7
hbFjk1c5qON3vWJNJWMd0HipVs0z/YFspTqTb6ssvOL3WFy7Lyvq7BHJceIFcmZGjzcWITQyEzkg
/MWyp2LVLAtzunGw1J6OvzfD7fwaGShbRVhBJI6Mcue0qZia5Vj230WVLtiiopX+ECBjyT9nNZcW
DB+0cOpG2oNTSw+nsYMDWa1ULLb+TBHrqH9U4zSLvRj/uaYEZT5ag0eDUc2Mmvai4jcdM/g+fhl6
2BXNmwe9IWEIn44i9dhoeSHxjUmESTIGjko4LB9qkF/LAc3XymjOmkJgKFV4BGlxPUxYJxdN+FQV
rQsVV7nUCZIHdLw37Sk3zFXbuAc+2ubK3+TXESQFQL2pyAvX60Qb084GKdvoQeVmNGOgv8vAONmt
pFuU7VcmEffRLQ3lcl71fnjAziXRuemqM1gxBk13BJ0ezzxeL60R1Thc6l8lWJvpmhWwdI9XG/lk
tWebz1SFHKMfSTwQitwtF/KgIcA4PGJ/HXfuYJPDFG9uqitYXLqK9zgLIxu3t315y3lqF27Y1UrE
4bNZRsmUYv+T8AG4v8tE7IlbPTPBPC0qqFrZPkJsOOzOncgUwN5gBxiDbKdpsrtmVJGgRwGcTCDo
S/MqzO5Kvl1LtQV5DqeJQV7Al0c3GI1a60m4eeJFGiz0IdOTpmSsA3od0NaaZulszHC1h6jqVIcT
hVA5Upl+aiVZ0Ap6Ie1UXagfCF/e56mInIic+B36TlekU5PaFISfZx5bGDLxwBQhvfHLulogxjFk
43hfPTaOTtvr9aqGYU08Wo6li3NpbBocSMQWohKfR/mwR+4hBvGj/JBm7MpJOsptZ+L57JyL5guX
RQ9nKwOPpNlEEJEHKWYUDzJDLzsdtA2UnolfNwl9hRRr0lUYehi8QXB3zexWmh9k0P5fBCNtIzSC
nVSuhS4iQwuvo/kJjtj/5IpTKrGOoCxIPh4KMCooA0wWLjNW1VgYxp7GtJJDBtI861WENR7Oopxq
obVDOCdi+GYG8k8vzmBvPQezE9cA4T+3fqHUyaK6j+kCKB23eSW0A9DriMtR/UmkG4q3AXKCZYIs
TjDBoEhMiATK74Eud2t1CujjyEaFZ8KnBlGcR4XEB93l7h/ket5AWkDrN8D7v42PjKidsrIpIeRD
W3lw+aHQjOfRWDFD4iVgaL1vkq+ShiL7zTOk6yS5EcbspxhLpwWZEvnaEZszHY6xdjcE9w/dDcak
JwA2UI2oy3+18SCpSLanpOPpTnDFbjkdHPnVn7l2gboHxQ93hr2OkiBfXreci/hoe+Qq3B+GVhGa
07clQzX6pjJsstIY5uvpkdXygvIIWE91skV0O43ualpZB2bwm2MeZ6UOEU5O3h6vxc/OXM9X7lcc
KqpnzpV6IewLYQxP/pJxIGkq4yUCrflahgiS/iavcuXjvCEp563lhdSecCz7usba4tDecIRWqJwF
2esaPBlQSkxY4o0v/kWqCJc3ghO0FCYVTg5WN4PCEk3CGyp2Zychtp9ZQI4wFN+TzVL2Ner22Y83
24vLwqXOj3/Wtnj9gA/1Os9UgkjkpK/YmcMnc+uyf8j6tBVm8i7KjGS3verZYdbLS5rujszOG6h/
3CxticT99FlQBqDnJjStX7Y8I2AXFncn0Prf5f3jwOIBa21FnkHPXf7HOdEv2cUpaKZ0I4jQrUOD
e/47RCufsj55saE0hz/pjPd7vYnT0jh4MAcJITm5ZrPWvlNXgfNwi7gPD45RIdLxLjjwI9OYwNfF
eWogEWPIPUJbh7tsm5GrKyIdULIwM9+J5c73TGoh0SObWf2F4jvbgKG7vOoisHquKj73Bkq5CoJH
zjAUZR+5DCF+nNl9r2iH8vZ0IuKf0Blnn1bg/S2nUcWnWQXaMhtCKNeM5pHC4xE+3Zzon39dTLYE
cqG5lHrhnv0SxGmslihVZE1smzp65ATbMRTtQrSK5j/TD/Sju9xcxCuCGabdQmZDfT9A+LURHCPs
RdkDrt4Q3hyFAb9YQNYsKrNiIKtPVwJ2yc0mDoUBVYM2FofOHNosekiZe/zFEOY2z4xaVYCr1PDx
TrzOOgHX143dCamsWbfDdR+8c42J6viORO3zjS/qYEzudkmF5D5lC+nXkejPEvdK1yt0I5BtAOHo
Hcg2FwFLh5d1inQ4XDuyadtDG9H38h4m3VZMOGpiW/NfO42doV+x4FpiUC4Kg6eUzeO7Uipmm+CM
BRSbWKSIRCy5DC70pPgex2RKXhtE37GwirqcMswD/kTj+0cJN4ppHXJdTO7FRV4Ps+Dpq7TldHZZ
pWOpwiszgSJH394LjTIX3PID9GSFryeUUClGj2gsEY6bnDQJ38XI20Qio6aZ1OFWek4oiRfopfD7
8dsySqPmtT+mPYfHNZ2dIHTt85atLWKHXKassYiKSYH+hZ5Kzogxz+he4aoEN7bsr5UxS6Nwy0B+
lt8AYw2DS3TAnh/uQdVGTByjngWWtogn/aem0mZJHzi8027pK/T04lF1ShfAtqVCR37BOg6Bz7Yp
GuZ7keAVXh/Nu7gwJz1N27wQt8rxBTq3dSUjBRMZfFTHqz3vBSghIdAe+Yp5dSKKAOgIuXJ0smYQ
8zUSnKkCiLb9TASnllsl8EuKjqa93UaCTayx5JPihJPKbVdQ44CzUcMvsgBhfyQpVx0J6Pb2CyEI
Xp3uiQ6qJoXUPFQpLvFBwOIGz5iqGatflMx40REliQN2zreHOPh4DdO+QDtSoWO6nGUrf4jOUzDA
qZo6H/ktRzXDlZRq3AdoUPfKSLnwerEL7wTjv9ah9iC5hC5oO90JxJsq5kJ5rVqduE81MZ7tfyFW
PTurndNTaNnzukbFIVK74rBKYTtTNDtaN2LQG+h8QE9yTJmprnQWhpVaVicNdsImK9eCIhCyihKg
yZ5fl4Q1URWZZwDbYoLMJPqlVjhgwYOpOqbfR/agODmAONLStL8Y2u0+pyUPM7hwlU1EreFqZD1j
24uk9YPA4yfrqm2F+een5bd2bv6PaZcn1O+z4bH79KJU98b2aAVTrON1uJq9BS/IhObqNO89Sxj7
Y6AFOX+fPlotYtJDGokBgwxdJYi5VZpqsvmMFzZStgn7Ft78Rmo56kKmXFoeCN1hNMrEjGwvfWdS
DNAh+C2WO66+I49oFMK52pbotcD80T+W325GBCAUDjblG3Bv8vnBxBDCXYs/AiiHNEuvcJQo/2Hl
0vgAiLMuT0/sOFx/5nvpWVlZ7qla7vCvuXDlxbojJGzXzeURt3TNtJxIFVYdjdWkiKqoehUqPULm
QA1VsJoKq9gtjSrplgREkzAncT5VNv4JT103f5lEp9wOKAdmUmqsCGOmLq0cYpZ3HfidpJLvyuzO
PxK0V1J0i1iGgs/lt9Wo4Bcs+RpVRxh/rwbvCZEvWaLYR2YdAFhphSaVxuUs/r5byIR8p6EJRoZa
PaM+5agB3itLVwVESMXLZQz+Z6Zki9ew0UmeIHjOrZCNReKD+uoObFfbxxbxiD9zU2gNSM7XO0oj
QU2NuML/AMSQC36MHAfeU11HOUcBg0obLl2nrGI6LaIIww9k97h4tEloLGmKpM1lus0kMydKXXOx
e4XACNQnuz1F69h2yxYrsuH2lZ3uIFf8RydHQZ7vakjP5vZ3r6OfP3Hjm+PFjAK/PMia1VnI3jGw
Ipwc40bBxq+xoqGS9mzKpZ9dv5/ryw2Ze52mpNI1jJ2Ta5tJF2SIC6ne0OsSjI2YCjDmXffTF1OP
5olW24FEzOrSuu6WeslXoNVNQCAcfzVZ37pbnrZymB9z8yj6vMy00Aj5GwPdDvGNf1O32DCxcofz
FQb3KwB3IBfxJMNcNHV6qNBDVdywHye8/mBCHkhGWJTDRjy+ru+tAVlNo9uFqMRuN9drm9Lh5feI
JY+iXFgIoxDgeiVYW6Wp51Mf/K0NwudfUiawRBgSXYiCvaSkLoERX41AIAMqi6RSJ9G8mTsuG5EV
S+zH9SXxzRhWO9MemV9cDCfMgxj3pYATXGPwrrK3gvtbvCWDdwnezrJ0X1+IhNof7PfbH2x+u5dt
FWrhTIZPVslbpgvBeoao0UILR/UUKRT+POJH56X5qB4s6zvSG+frG+fIHubzXfcRdwtcikzeO4UZ
D74Z35zTTGus4C2wk4MT3Z8M+4KSuRWlgIXaulIkoo7QChgkitrVaeX6mzN98RnqRIPfbnYppMxI
E4112VgAtcQeFuaTA/P/QAS+yJaPuFsJKuSyhF3qFB56MrO9GzmZ6MJB40G4oaLkUdQj/6I2ceoc
EecpOz5NyQ4SiLfTWeRhomR2a6ZJhkcNU8lOtgT6HDf+tLyWb1ktR5Wr9GFt/Y5BMNB6Dh7s5Z8o
LmD7tf6VrTRX/K9a/p8BBdY7vSjha9SEJda+q1c+iAquhDTq3hJY8uXThfW9yVMpjLrFg4oLUhZf
FLooxyzxAqmnq5LchS3RcqlfK+Nj9TJuVJ/WcFtAQ6tQoPjIfcQxTZTlZ92gWEg7P3UCxjSSb3tv
6qIraLaCCPmLF16q2MxenGh5mljepnnxAOjJfuwF3nyV3n+Vh547523500Bejt6TA/G/v2zTpQ9Q
RAMog48stVE2USim46QgpAns4lXvwm3oRyZ5oBxPtv1GVMxsvIpATjcO1Com16v9HgWkJYOrtIo0
RrAV6HvpmcYGNXhxU2tKUbcF0UknLRzUEi4awUnthDLFbYi0seOQe+Rxia0hETT6cOiY0CvXR39w
/GNyJ866uj8RByiJ8t85Sf+976tfXD4vHUWE0Kli4C5nL8V6+0pU7PnFb/Pt0iRHY3rnBH7xAFDe
0xI7d8vHUasy+cgUJnSXy0+zMVP2d2XqUmD+ymg1jYYziYLHMBw0F1SYjAxq6Xdvr/VtOWrP0Thk
5+TEF3+X6edIbAEZ1M+Yiwj0Czi7jXHXQBvkLKyEI/e028g479UVBUdcP4YB131F7xmLJiV9E7dG
9o9+Go+oTwb6V3o4l2rZ2F202GyyXKEs8ZkNDueelNXVZ+EddFA7CLa4YQKa6frKIohcYEU5A2pW
kZ23qZvVWLViZqOKXz14e+8sM6riWaont8f/PmpwHY+35o19TAuSyBkPieNnCVII5sjYjGk70dn3
W1bEE4o89edYsXCZlAgnEXFf11a2Jq5ahx4nSbIseuBk+oIqLImirMuejKnU8PtRWPJLwmmBnjOc
qvFhXgXi8cvktQM5xRuFQeLCUfELtr7V6//b+EM6zEr0XR/jAXTcigKoC56Jojg/p770i/hNJ3Xr
wIf2xHKisfJq1x0mn8aA7vjn99ZuRsIu4oz72E6REUIrgCNiE+ya+tniU/BUPE3clyzGbZ3/4b3V
6gTPwD/byKQ5DRglUdE46jkPnHttPq3mF0VDvjSPL1iMEfuxqXJDV7Nls6s+nWtrMKdP7R9PrqUl
qiOmZM95KStw6qrjnByj8eCmC2DeTjesP++Me/U1zDDbS6guQUOXJ8pt7pa69FsHvQOMW9A14Ugf
xGc92vLQ9p6EmIgMBoeiw8X+MB3I1E93U/M8O7Cn23yzzfeB7XLyd7Ciftzoz2sQJRGC5pq6Iclj
BaCvIMvAOu60gA8WgwT/DA0oX621BrDm2+dKdPmBckYicemQMoR4dZuxYj506wIkwD+GihpX74JF
mgXQ1ynd8ZWaCB+c9kna73o40d5nLeRu82uqpdpuQ5jlvmLxH8J25j5SCt/I01nPPoejpphxWKgj
Scd32ugANIOjLvceI6FobGNfinHXbqriIVZqpVvH7CMVD5Pa7NvtrWm7+nVgeUy8U9MhzQ4MJt5X
JxK7WGAIQm7S2V2tJp/eb8GqwDDXyKhmdr4WVkB5RgEqffWCE8LjDo5jNqpdUq8cFYB+VOH158y3
TqMKLPTZPfSvSi7LTfUKdyyr/5UbsTSgg1rrhqgxO6QEKO9PtYaZcCEK0SzGAtrJSZUWIvyy3mJd
hakZ0QkW/tKcTkIWT10EE28HSiHk6emE1y+fsvBT8fsxqFJsAc4mJJ+bDNGaEIzywjvEgXMigFNr
ZV+wEcGkxOiLikH9or5hYl/JlEcoOoXpYNNfnr/F175Ad8PNxqv/sERtsKmeP0/O2ojTMa/kz1OG
KSsPTkvPMYddtyidBaSatZvUHu7llDIx+hpsyItsLgVVW/ZTHb4zcgtNjWBpiwlv1M62f4hA3ZwJ
N0F4nMwWBz/Z9WM3hApbKFQHHcv5kf6AuY0J1JIT/K6n57UtKgWirAtMMqLGZ/PBcCUNAuZtF+iY
XAtOy8qwxp6a5Lj1W3M9f9FE2yRrKYHMxLQM5W45LoDfVxv1CeSB+hsxYUtVAr/fs/iXrKpg/c5z
Evre17Q55ZvZhJlR7D3SAIKDp1hYkc3DQ7TD3P2+txReDKT9jXNBRT8oU/KmZ6ggw6HXGM9i/SDj
0XAzUeok23wJ0xFmSTFQ/7zSRmU8FN0xOGWFpRnXqfaoSQnNptsNY24to3fQPAs/e7Ww6Asymgtp
rMJ/6+5lA6j4WboxzRibUm6R5kxXbNOCTwLdpO3FAIwtp3LXYI44gRgx91npfQT/1La/7MqCTSw/
XBehRgTlhB9Svhp9rYAsfbwh3Q8eSKZ6ARomS8INyKig8VVdJUbEiuJvZSGfNHf93TS0p2/1SXPH
6gmtwVEP6JgI76qX95mM8HaQ18L38poY2Jeo1u2yegqifVrkJc5jNtQHSlsshNUt6tqEDxPtxfKp
pvVWRjM8HCEbDlPstzFmkIa2Ahs1ZJ1411zBXe+f6M85FPbvea0uDSsJ3OOFINLGo/e474KvQNST
0Qc3BfjPsJ47gMSKjlv4nyUHUBG8ckA5Gn1Qb85ATk73gYwGGrtJS4uD4Ar80ykXBUna6vfV93cC
T7zoH0hjprYb8arkKwxmy/HoO7+55GgTBZT463XkLqHjcKij8bNmuwQxRZFWZomXuylTXonx5Z+g
NlzFW3X4XfxpPKcAxNQEs50b5oxx5ugcVw71DTkeApJzv7Bkv0SlFZo4+8xjPIkDdtOT9a4zwpuD
+IbC5kpdqDSwqpAQdqcZlC646kRExoxWYUzunAXnxuIoB5NyJsD8CMmioAnzjxMprzma59NfsqcY
wt+sGG0hqB3b8jG3YnxAl/k9dzF2HgjkG9YFTJOMJFf6ag2FbkVKKjA4u75ga0xZyl9zcYYFz0n6
Vgf1GA4ykbJe7EKuNZe06oVcdGrW9lJihQMZWETByGRC27p8QVz2gM26Gp/daHAtTAr/wkg4RFHr
nNyRl+0Q7OvedCyxMj4r3oLLhSu1VbiLIrHvMdaw4z1QMS1+vknLDW8glGWZDPKks7KQPCNYvbop
mxO6/3Et75TZX84oXKnFl0482fNmChFV06n2Hlq0kP8WsZVrIuAiD9IN7iQLIwDi6YtMCd3vDumR
DcaXjdRgQ/vnNAywGhA3aEvanFl3XILjfNF/chOJ7Vc+/q6EfXnuFAwnEdpQ2/QB7x7pe6mq0BrW
OeXh4jhOBAzq34efSZBv9J7svI7jGZgOSeW3SF/Jq8RucXa0VdSC1fEJlpWvYzH5ubdBJSbBlr1Y
Qv1e7y+9jeIFBM7c1zPyj5B4/P5O0VImS24c8KbXaRaPzhZOabCe+OBhscJKjUQwm0Df0v5Adn4H
qIH4b1XbALxc9W0g7KbFZmKu7GHMC5ubobGRnEzaFLqJkCctcSEoWKKlhrfm36XroXYEfActhCqc
3a1QWWH7uztxzDoiyqf2lQaUvq5rqn+7sJrbRdaZmh/TZQp/DatgogN1OkpozhNsHBGM3jx+XX9l
eZM0WF7SnQmPml+P9Xb+9Ui7Ms0D9z0b28lSTQTzpTgrvdQKZuFlq5ygIZzzRONkxyNusQAVpct0
/rsBKXSIl8vIPZsQiVQuujAB2d5htTS4J+6tohzm8xdmpDM/89RTz84pZpr2cftjzzf5FWf/jejH
WdeCPPGhdCrPrIXLtHIwusNK7Wj6S41x6pG9G4zTUFJ2CRiaDcqIKreciFuoaQGcZkBasW43MtVk
vMNI/GGvYtC+PuKISQ0U6J6JxG1B+dix5xKcWkPrX90Z5AFDvGTCvdIlpUjPt/qZ3gtk9ehdv6wz
jhbrzuMSVYkvTB0Juke3rievSazgAQ+Kg9SM8CUq8lkHh9ErlTduowNzdJGlh99aOaX7Ftc/eF6w
nsu95Iuo3VC7XGLn5a3YthWnz1UmlJ22K3ccEH4wTn0mlkO7MsO2vw0QkQ8YyAzs80OKAF10M90R
EUVgOSTmrwaa3loMSYq4gsyLjSIAKJwaJ6t2PrOnR7uSUtO9octT/Waq9RjUArUvZ92tne0tuRtp
8vcekJWqeBn7YcQcqeC1zivXv/uCFcRCVDl7A3DphXpM9jbcadFQCBzhxoMoIv/K7ZKgrj2RiKnf
T0fT+LiCTYNi6KD0Fv342nleht1Muz1FrNxC0FuxaQ3KwKokGsIGot5yxqCdEeYPVkOeoEF2U0OZ
x14CSwZxXX6rDWOxWVUXxSme3ojfoK/Fb4oRdQ1BLI/RR88Z5m0pGI51XQW+PXehvGrvylgl0764
QIQNy/6Q0zn9lsFNUFX5l79nPBL4mgwN8nFpiDMrrY0+xyqCbxRyzsYxsoOQx0Euczn0d2ypNrgA
mgRdhLROPA658uUajlyQlgAvZXGpN/2ZWffXGRnE4ow3gzp1GGczyR8UKYUZ0+3lBIF1uyRz5peo
L2Hf1178Q4QaQw6sL78drewb7D6YATJAIZ088EqPXQmVMdgdZqyhCFY+93rxdxfHM4cVdqHp7vmA
uG63YkMl//LKHmKVoqScUSXSKvm600uj7KgxWE3hbNvqoelGWOXi0LUtmm3O0FvrPB2agAfTdD1l
Q9eqHEXEWuzroFBa7d0YbGBfMPuRjl4yB/8vMuATo7GVAvFdN5A3glk1wJJKFeYw7TDwJW43w6mf
rLvRSYAJcSlDdtL/arvci98rafmxLOoRe53jh94mxWhOvFK0UtgrZe/RljehR0DzScTMRLBf57+s
XvIqLwjtNGWUcn+jcZG2oQxdX5O1hYlcnFiY7ud4y5a/KkupB9G92NSptS1NHjZd6TCVXwjsyhw5
oZKKp9nkbOkwb/e9pvLza5fWQ+zfW9zMU3/DhZRINipTKG1QZMVJz/yfyRhnKcOia2A0WPh+iVZL
hEwbJFaeelvZftM7Xji8GMqgybpOIgQ0/gRwsfCTJ0H8ElPO3No1Mv3c+QzRfTgg/9euJPU5rkTV
/6+CqT2NzWfv1Gf353gOcy+LhLaD/RgGbD3lsOZA+n3WB+nw3P9plMTVx3Kki0LhBqlgqwStjZI/
guSnOfqA/QZmUlDOSC3eM40LS7abotJIj65tZlOkMJxGdxzVIbjd+fUYTRwuVPr8ADV19bmZykzA
22ICoC25MChF9u9oUIbObXIF3kBaw0D73cQa/B45ndwDxfa67YVGugsy3F3IfDw+YcA7H+ZWy8Pr
pvY6A86ITslPUOM7X3LBItbrRZBn26pfQr750Stuyd1xwyFQwDiocLL/wI0vhmpTYfVFcqPNGEzS
CzOkaOZ2+g27yQE95Yp8aUk0gEBHEwn5EAe6jHizS/3yd/worLqpcQfr6aBpdEATPg9mxbPTIlnK
Zv999KZv1rL/Se+03kuDQdS+TbK6OVrE396JUMWBdlelz5+4W+KTf1hl+2I29cGWboskqimUipnV
6O6HT9YzwQ/uZLkDbH5SRYqliHd7eEpAHVmYNlmbe5sysjI+JJUZLoVCuRQtPAkNNjrauWsFXiCi
hQjxDsK/P3yqKKxvWdP0BwcyTDsrpU6wWv6+mUALGEuAkJi7ipFXMPDADs7I03jMJy31a7rYTP+a
YivVd0hjjuY+iuvkmaCVfyrOioArUCVUEl4CnHHUnzBB6+PkgOBmOTfw/eMxGQw8LG+Alzfa7lrE
tE6KaAvdsadEMpZztJwp6KI3RVYjKr35mweuScR7/wgzCrr445/Ga8O9BOk5D8Ex77JsKzYDy8w9
NSQcKhDSeXE75uIki/7jGpl2PHH1lb0+UIHPXbI1jHRsZYYKiYaqoTWGsa5dVbuRHCggKW5rrsTr
T2Oj1nWzzIqPpvq2xb7bqGyYeDHTmLyOZ+A22jYjfkVvDGxGeLpktJIrQvg1xhv2vOp4m+XWQihi
Ytplz8EpdGlPV8twBJGaFC9oQXtK+DHow3h3emzyYU8xk9RxSH87zVlAY+1MYre4+aMZePvtuzbJ
tX52rK65KQvZMR8lTyxo9mA9GlmOU5m+TrpR4NjQfoc0+K+EMdrWyaKjaypK2FI4o8wtr2vugd6q
UVHYeDZcL0dJXNX26MrGcBWb5DS13rL/991qWFbdgCSgysjVQI3/1ytb9oogtIhYCTTX9x26mUzB
timSzlbtgSPbvvFg/Xq+N5lHa5gzkp3kQr/uDHz1SEtzhYYe83W+hmYifPijh3nPiVwoXfDikIct
vns3KRC69nRA0AKCzHQ6jfI9/TNp0EzS2UlEAbQwe+7T38yT40IKIhmEkE3OgLwSBin6OohtfcFP
MWyRQsXMvPXfA50G+C0OnXVq0acikg4ywR+3/cU6LsYIOx0Bpb9htteijTCOvWSVM1VxPcZV2QWY
sZph/j6OrYnXEgZibxfcABOqb/u5YsO5+NwsBqAXGrq1AllmdIl4SQRImNwlFKAPf9d9Ddh9pYTa
v9BxoPq/7lviMgjdYHze6YgPdKKjDBCcGlUXkjclvk3Km7a/kaLtsQDZ0IFB4Vcam30p3VDJPtQb
TIOWym46+JlfHAENPE+W8zm+3aNf6ssxWzZc1jZyouZOgJFVASqG1jASjooTyRmXEEWnaO7S6emS
IpC6S/83UULsgPexsGLGNGSIvr6OKFdHBETQspedDNUDYuUvszQG6StdhfKr8SFzFSRAfAyfqeaB
zdKBHBZmsakq5lxO/4TuUfVqO3TpGWH9LrwmafYhWGNYU+q1V6FISgv9kjKF6OxWkTlzyYi5T4l8
s2XBVJcRJdgYE0pEeZmWkJ78Opcu1gNQ0IMJKctcDVAT50IM4kqhtDgPNJTBHwR+TTtby1WGlvwC
c0TpLpqLefvRfh9TkfIJdD6NWTyqIGTYqj3zCh1Z8HZFN0cmGZUud4k+o4ulhaluLGWSH9wzVapW
ItNhjevx8WU1NiPtD++BVWQ80LaOTS62eJAbjIVe765h9EfdjZpJaVUxOeA29DdOstps6m2KNwSg
3jz7mYLqJ3uWh/zBDh0BXTfwwYwhsEOsaetweJlIh2KLnMjoQPIWMcRw5j9sKIF5jhsYbssTrPT+
lMJTK8PeHPId3Mohjn4b3xQ9SJtVSSuuiLSAleWA2cm2MeqsDN2KmuzIVobZyRf/gBzkTEkihyNY
V56VHtAe95Zabb1iQNlZmQagyJwuEqRXt115o6cdRFmHUOyky52QYSL3SSW7Ccbofo8SpF9g4B5j
tZrGdzdywzzcwC1J7rUaD99tje33dTotlCTOq6Jr5GPxDA9Rnv7/CzFXOKI0SVkJwXjPWxNNEWbZ
nsTvgQaDDRWlOm2PUPDlWcsO4nQSPhiNB/8wB9jYo9vBVGobRfcUHtKT9FM9nDj+6Df4vtCRnwKm
DeMrnm33j1rvdvhQwPxslXYhK4QGFZ1oQntJ96gN4OKfnbWCfMVnkK95wPDnfCo4rGeR7dQYHTCO
5YAALZF7snGzI7faioVH8kCmZomLn/YFr0ZfRFxm1E2fWj4waRpeu3UFVBUSJHr8i8wSAtLKUsiv
+4BRFPkuz9gipyS/H/gUUNR9OzpRFPtcicgkx8DROfMH/LROfV2tyLyuiueQctq4J4Uz3ZZ9Bd1D
dj6NETc26L1kMbC/ITb5frSrsF1F2VCX6Iz7BskpIZjtcv6IWcbkCSMInReFDNMlQetuy4azCMp0
Af4R98r17Xbi3jy1DRFvsERu0vwKZFqg9g1UePMI7fg18sGrE0Dg6TckwTd/Ngkn57ncHBAblLgE
RgF7yqvQvFVFWuVwti8YrF/zy/LzrMTJFKWVYAGn6z4ujqHjCYxCtysNCa1J6krul4orvyB+OBAR
idaHgX3sTzWCCsGH+fvL7ShXSweeqovdujipNLHVp6OeWZwPBsCwXcuMF8HEmorja3mIKv5UzOEU
wSEtHp+zGabaQsKFkjq3xjv6dkGyMr94rtHl3+rhpYQm10RG5PLaIM8rl8G2Ekr43OyTQxOlwIwt
yWVxOg8fKJExJTPh2ZXtlMxN/+7cPig5IUsF4SY4DRvAS/xBXm3rcnJTIjr1dcsL+4/BYU/UEW4N
8GQmXCerj4ErGJkDhLJd3xdQtINS4jQtst1eDVUuiZtg6txvGrcMg4+DmTUKl/okD/XPVxGwzMLd
5CkC2avdOQAZnBY4g/tGSQxjVGGKoOlK+1rMWYIHkix5jXqcX9eU85VkXaqpqTC2LL+kOA2Bw8aD
8KA6niWIALpSAMaN058Oif+9qUgx3pcPaO6wx7Ro1lprjtvnAZ3cbsqtoT5/MErojHWtcaX9s7in
v5MBdLLvx6i7Gb2VgrOqswK+JLWwVLUkKqp2mwgsgGzYv1lRjsLbifN6DgtoR/dxeUe1NsYs6Pgv
9eCeunemIpEkoTfR/Vh8/yt13i0yWqvfPtaFOwa03cWDKNq967l96FoC3KUE9UZpMP6/Q1NA827h
kBV6vmS7SFCJw46n62jPgS3Z0F4hdQVvIIgXKXIG3J6TzX9bw0n/pJvYcr2ogLiwDMV0GgxjwIO4
zds2ibNwc+idC1IhhKTmUfmsaxwAQfz+pf/UOjBheWbXDDyLnPJT2bkEefWravrQiMfEtwuxY2l+
FneD2YIf5UtDJzZKiYjEpJ5plibo4DN5Np6be2k0TB65RgQH7DuDx1MWBTsKIPG+nrZaVV+G0jwy
/zqBOYAtDQnjO/QJ/Rfz/CD4/rO47jI7OG6V/exycfX+tnd4Q3hHfCBZXK64/jYWSzoGS3Af2uCI
heuKyv1ZEg1L4IsO5jHLERsivaDiKqbKpsXjxJqAxg+bJZS6E5rwvdz9Afkepma9ReKHgxR1qqIL
r55lzAkLUAU19hvU+OD86fXycrXqrLfPdE6IQkNVp70uSs3Py4iNgoR5h3XxA16U3S/KgHYt4r7E
lKRtLm3pYOl6kld05mUarDpbqGp57ORj1F91sOjN5ANHJ1uUniirpQ0hyyG9lCxe6QKwt13wJbhJ
R3BAsCUqz2Lfq4F4ZVyl/buINUoK1vQJbNlp+3HmuauNII6t3DD0g/9j5P2t5tKORd2Cd//4TmwI
wELfsjcqnGiDgKuSQvRNMOYKN3aZJgd4ot4vF9AcBVtbK/DMlrEG4pHCDU2WfIfX0jfZYuFAN8Ht
b3+z088zRUx2V4Y3d3T5rh47gbiQoUrj68z89qkzW/IsLvKvgQ2CM2d29mYeB21as7g/8o1PxYlt
aIFygpX0esqbTW1OLOlxFarrQOR3swz5fzkByUDhi2WxT+8yqrFg3ZevGjvat/hZX6grCfZDLVIF
TrpurzRvHKYwVQWtBOw3n7WYWCDEdku6gppbA73OYIpLp9cyHSce7F9hdWdPq5Mqil4TkIwr3izd
atM8E/ZPTkHQWhkpMrm6FOeBvZxQIMUibrgv8WMLw/5kBnPWM493H8mJJrmmIv7oEAW7nWBSkH3t
gqhHbZzEuEYEWNOu6/cUi/IDIfgjreiISqr31NhOebcfCJGzEnZxdtklxPn95CML2oOpGIRBSWTU
z67OfNn4OFVWMr+LWsaurem0f9tFV7aCu6dzYa5scsc/Sbg8Tul/zjUV85sjVywuIwrxmZSv9OUC
+XCotKdVUuPC2DtGh2B+ykMpG1jpHD9zF+M8yH59CF7n+UExgdmh514q74nIVuwvx4yo+U2cwW3V
AJ8pIFEP6p69UPCv3ARnn+eZRJnM+gROBxJFEqWKI6BXcLVC+gH/ilUJAf8SmBcX3QAlzH0LdX/s
49+ZdhXUX2fTEa+nkK0IuP5i7T4r4pLUhyRjRDYO0Cr/FtdV6zm+I3jRSCVF8w/NMtJjrtfRAJbV
DCk6C+C9C0sRprE5VF18JuA9QPUyNjbEBmHbYlQPQFPedakndTe/h+LCV29iOebqDcZA5OZ9IcaU
yUooFBejaHv4jZJw0RLLTT9v8TVeSkZoJyWyWthsU0BQMgAwagcHUCHYwIswVnvpZVmClbR+qgP5
8lRQ+5spxgqG8Mg9F+BUWlWuZJEB11+9Bc/+esMROG0uRuwh9m+KvmS32dvySjS+yFJwPnBYoZc0
Colm3o14JplF44LmMQZyDOIamQAWkr4DIA7EXe5s6DpwY83eyjnZm/QzmuPRJo/h+QnPVIxuvBCR
TZEz9zu544Ah61WMeGvA+E2k/V8gcgEwhnL/44y7GLzCPq3Jtc/faSno0Tzj2EXQ7jlHt/TSb0D1
6ozTSQyWehgmoRVFlpZRy1BUVnad+3oR3/85UeEH+rAYktTeDmnC0G3iu2GFKleFVoUjE+c0n9bn
iVEp10jfbjjQtwVmTGmo5otvjTogOvLszNow4F5QvRRFvNxskkrVP0apeUohtrA8QiIIewvbJhs3
0Nm1mTBggW1v49xxOyhIGHHxhwj5TH3MtEEfWx4TaSl3lut4cxygDWJnCOwaMi95RdTEy7yH/Az1
KT0SaxU11QDfygwbPBuRaZJLhfDubZKK8crbkGvUY5ggZ+zq6aB4Kuc82IiNOQoAtbG6IHdzt5JW
dT9So9pgQ6wNWMgjEd995gIvHG1eEHVDOToBTCbLI853n8mz7BEfHo2o8nx3aN+0kj4t7NFu7eAd
4FFx/CBamMfZpetes+Y9x8F8Cub3qwmGINdJ8zqCcityXnZI7gpCFyN83zS004wbQ6xOk5f//F4m
qCLbNCBs9kNnK9CVZcapfgBjT/6HIQ0E9lq4kqafu98QntWeW3o2MEPz6DF/az7+duxbfPfLGLoZ
eTnJuWxqFPktYroyUhthNHUk3XCTarqphZ53b3yF75z5wcfzOLx23B8evzpVr602+fS07EGO5xGe
hW1Ca9RTmOE/VDNz/8xPageO3vSceWDYyF0bMx2OccAnw1YpxFBOLC29n2lgXObDXwqxsSRZ0Zo5
5dB2PyPmFmv7FLScO9S0UeToZ+FEIuwXl5hFo5a7n4ySWD5NV8k/G+t+6KB2MmehnjNSOep1gQ+T
depGJIrKfD4Ph1YIr4btclYVEDhyCctTytl3DO6ZWcxbWgXLy5jGIG0LIMK5FRz0Lw4lmaM8vXW8
ZllG6o2rTkp75WBdgVcgqQtHg2PfhWPGPSrI+CW5gM6R8RVaNnAtGi9W/sUHwE2LNXQIUXJ4Nr04
WZ3qabsIrvy/PMJdsyB90zMhYllQTTS558U/TSYwEAVic8McNeDxYQPFqwX9/sOtzKt97cxv0PJO
5uZIo3PAC8Gh241p8uJPYqGav22Ds6kl9wI7yGivWOInXCPHgQmyW542BYgGm6nWoxuXReiW1pke
AsLJqPAwOyTuZ9yl/SFUrF6GXGN0cOj16RKiB+c7FkeuHlU3aYWn0d89NLG720azZsZcvKfjE1Q3
PUJp1lQ5a4QlayEctOyQ1zoymmzUcjk+2swObnay+rr+Sq8iybcGbuVoGmwSyFzgpV+7/dw2ONwJ
UzC7RdVqhUKsvPoxRLrt8Yn4Q21gLBnZU3VwMyyQEbOowsAwoEzz3nMFhqG9ePLZGKu718aCmzjJ
uGtCzzHGSectzlBOaHMt8Hrgf1Pm/hUJhlY2CVvpTE2SVacqZ4JR3b/Mxs3wXbwa5VAlGQ6KTeDB
EOcVacmUy18OPQrgQcO3BEDGKdHJbH0GeAHtSkXRGVIPbaSyguAFjZZZJl8ZDxKXZYoTUVuvkm9B
WxldkNWi0skudjOqQqPBITbONYzeBPng0H0UFxgtynV1cpdbRr+BBp1Z2l15geVWuHav+0aK+0JH
B2xGxj0NM+o3LoRh+CDWIGxOV3oQFQowSwpv+lvy9I5ZOrOLN+tHNmDZOYRSjQBNXvHjTAffEoMu
j/KLGgf+BSCzLC+8YfBkX7jg0tsSZHrp/JqggNLf0I08TpwmBhyk0KJ5rRxfF659yayLGHRmwMLQ
sKjHopjTzOTrz4I3ptHOIMLOStdh3C8r3ZYfiaJJGEgs2IWL7KXRnXAqvJEpEaOF10S0ReUmiCyh
2RbYxga8dwlhVGoxeUXeQ7hNFaLLB66h2bir1CXrh1a0d+K0SNpitcMbt3nxZOxclebXjsGhPR+n
kDdD1IETclVnH/MUrTDEGh82VfIwSRIOTaPyys9nDNSTquzVPzyvW8WaUHPZ8zq6kULYwfeaSVon
f5F6ZuDwkrHBriLgcYuf73q0OF8nIIarApewQ53tDi8A9jQJY8lXl1B2xvYM3JnAgB2SKZxdt4OR
zIqH7g3tKhleXSBbnsgghu0val476LV5BBzFyYjdrEsRazLCGro0CT9cBAD0oL5H1cRhPp1QEOjD
HzpVdoyfW7c47PWKv/OLnlIa6kwbEdcFUa/FIAQoYVYS1c0pwBIEX5KAcwdonBdjzn4FLjBO95fe
Ue3Et6sO7HsU4DxpEoV53vOqdYmARGtXYC49bPhMnXnVefRylT1dEUgvwh/HHkhxXv0lEH+ZvuXm
sNtNLn6jZp+2c/K3dhJsP259S4rci3qxcwFCQw0DvZdUV619z6+cS06ffGV9xPCjaE9B35HIQsLh
L5WDWjSE1RIu/Y+u882Db+VIW9ruOecWGcWvmU2K9ApU/xQZyDOpTsFulqnxSL7noqeSy/kmLyez
wI9wyUM4BS2h83YBuAMJQ+s9O1ckuHM8eUlug7+hTv3PYMdXwIwvIbbV/b6lIuWmonuZ2+UdP0yI
tYqtv57QMNI9vcVp8oSS/4HQ9lqvgSxTdER69BtHXzMOId+WYO+cMLTGFJ1RJzck5jGy8J+s0sbO
v7ST8Czeb1O2FSCOhcyHwmnS3+t+8vpI/vuYyGS4LGKir8vHjEX4VXXuY6YyOZGXfwTax9ENfzjy
1RHYtK+33g1DBdFeejx70UokdRhVqTZB/uz6uBYaIkbSky+d6MxHpYARJIU7oTvEbVyW/W2zmhh4
mlPczzZ7I1dRgzVtdp589xtyhvW+O5x3JvREfqaMJ0N8wh/qiNl8MJojvPlqqKAMeuQuzUZziDJ2
O9h/KWjPxOlSA79ri0CFDyCTJZKngErRs47Fef8769ziG6ETdVhvSkBmLw5S6dq9vgctBw/6BNI7
b3IvFIKwfxXV9LB3ViM4Jiw0Mzt4nWQ+fMRgP/URL52Q6bL/vZ8vP89eYHXoy6Azjz+yL8hz3mmv
ak18aHbP3XYIdiU+ZTRzPvEBZ2jrhOXFafpxIoKrEyhw32UAsoYDbJGmgB7y60Guqyt1Yd2dSc/3
XFiKukEKklc0tHGrMtq+zklSlxkoHx820JjsvYVxkfaAk+/tG+mWLFsCgS9wsp/T1FxDbdRkIMDr
rLYIZH+uAmAlsDLbxm8UzzqnxrkhJ66s3ATaEtfO7UBvrwKs3AwNE8NCoVrMFor/vF5jfvya/8xc
mwrtFjz+jB1i9t9LyjgDiOsnDyYw+4v8DLSfCntzwHA2W6kjrSO1R4bGR8CU0liznyu9T2JL1DUg
oiQgVUHY6oqU6bH2MXNw7FKRL9GQynnPRFH3GJq4LIzDGp2vEUs/Ee9/1NdZ35AWfF+PBPWUyMdF
abIRYeMxdQFDMqG7HyP+3EYi12RtM5hA5JANXl+NpU4yWlCpFzv4zn4Oj4citV2HK4aWi7uMAB43
iB/vHfQ9hbk+0sDOPwNXGwlZHTbgLsLrV8gbRPDtCEQden5a0GR6FPC3YMR2ggnPpnpLTO4jH3xK
zPjtdLzi+zyuDy7PASFNjVsoKwdhZFizfP9621kBaA+tXWppdWio7vYAN12vGkgOfUv0tSoSaUnN
P3bxgRI8uUXLKw6ejSTdTzDd/xsCu9akpdV97T2qeYUFDz/wJ9qhDsGt348VMG4XMUeoI+vsdwbZ
e2KGWVqWoTAPokUHn5NQouo4tbOr5m7PUgWkfNkGSdEWjrfs6mUfOlWZsxTarp8iGrbuyaetzZUm
YwOpuRpyNVSgSVHaSHp0fzx9VSX+krVGiVPVQPpXLDd79BVJbqFd57VO60ploXQ4BF3BB1+hD0xJ
5spYH/IHdFRzhQf+UmqrrTeq/ER7S76DBa/MwBYHOb69XBJ4aHs4gYDEwaua61yHTjYNqb31IFJ/
eVrWdRXvwtZAA8kKxDXxOkTdXuIgHFWw2S1Wdt42P9v4BL0INuPB7EcANDaI/IkuRMsBCMQ2r0uz
RKFLKI2kvn+J1Flq0/mzj1LaXfM6UcYeGeObV0y/qfFxC04H+MA7lmleHfibCsXpa9hWyRZeXM6f
dzOZI0tkxdZy/hMF4SdU1fY8/euY782DoE1eCwiaT/ojE1NjZHXfV1x3dS0iaKtE1czFc4i5hcZF
2JB8xucrM7M8nIP2BMyM5Q3U7K2HOh/Sg5sYrtfEqx6uunggN5D04+MLzRgOcpQ3N8L/KO5Muhcu
iX9B/kDa9Rp+aKNruJZfLC74uYQ4+rV9nNqYtuHc5rDLEmanXeJ03QjRDqqwlEl39YP0VV6oH/2U
RazO2BVgggATMz8z6k5Dfw0lWUa0dxaTNWb24JXDvijpcCpkhV7dJY8LWUZTfKaTvQ7s6khNieZC
D5kNDkCm0BMkh1pUI9zW7+Sq9c3axZ2GKmuwtsGs95RCZS9GBkKbJ58A2bRMV1nZgP2TjLDZWAlX
PRkChkOSEKrnEIhZWFiXVBKQbK0h0ERmOLWiG/3sfThdtxJlKvDg/9qUYQfFA2djW5Is02UKPXCP
LzJZVX9BCIdKiPG8JirEkFPFUuUHi73ZgEWjqXjxcU62005Egi9zYFXLK/zuwqOI+pNzYs3xFb/b
xpWrE35AEv5X/stMEZ9aIXiT38JNfOzyXHGnwVGLnAcIJKEOD1UVKmwaieSvQxuAupRB8KB1gy/v
I3IWnUnblKwFmHID7AwDEHahfqd7Flb7QTm5BPsemSJkZnBuRKQKXle4uDXBj2ysRw2sFYShD5gs
9NSyjepwECfAchns+iBP2XraXANtO8y9d80AOYERzdKsk+dsc9anjmXi8kmX4w1M4LzjsPRLgZtd
p9MC7Mjjca00hoqT2C6nj1sjRL2KyiR9DfrPOGaJ1/yM5OajULSQVrccmzXo8uRKKAdC1eVac+n8
qBJ548daLWB6sTznfcZ0oejxz8x6MOqcjieVMYLPuMPxqSLprmFAyACNrX0RHDoqliTA1nrS0JzX
BXUtmN8AP7r3PWBXDTmoMYns55wv4c+pf0vqxZkQt51mB76iVU3uFo55o6WXzhSBdh/UTqal6gb+
5DvRABkAex2qqJ5w3XNZ9D/Z6z63g1qUkjPokgoNoptdHGMrKA/EmHV14BAPjqXqZpyk1sOyojNY
MrhSiZBEEHvfdNH7SvCYDvcbPhMxfPiXJJNCKjM03qHhZYKZefhwcIz7zoPSszcy7v1FPxyrhROo
7mWww47WJIe7HomH6F/NL7lAQLijijq6fbShuqFPVU5EfQhYU/McYAaWxZ3Z8YRUi3bkoeOFgzzg
8ihSZ4yg9sWI1cXlvzlNjcKRwmd+juwgtt8bTB1GAp0u0n2r7Nsj3vDT6VAu5tw0cR1rC31oW4Tt
BM1IvpbeJbtC62efB3BO5X0GbXXPaB93JtwGFt+j4fUfZ+u7h7h4ZHmKLhrgGZUQnti4MvS38Xkx
a3TDy2TyuwauL2+G1qxjEhMW6pZmFXxNih/S56F6JawBYxZIbFq6i5DcT/GctQzaGuwrT7oyvAY9
8ykPC4mS9ov2A+aeLFUPS89w4eAXGF2cEOMEpdsB5i3BKF2gQibzVikJrsEjlUe2rvNHAozTsqm5
wbAMvb1c8hqRFChKZKMjv5vkpgqi/EoVYQSDsAWVMdCAPSVGwt1Cs1dEKakZ5J9xxmh2LMRHdqox
Exbpv/ieSboDLMs90WZ/vHRbysziLeIt5TYKp4qubT+sadH4Fp2AN2BV75X3CoE00ci1VCMwOjv2
v5yQhZYHuOUPO9aUl5ilApORY8VtFeA0tuvrw6N7oU4nSNHXJbC1dKvhOxoGzsO0pvfl1Ttd4Beq
GwIlvWZQrxIZopO3pNNC+H3DXTZ/X/MiA6YTYKxoDonAv1RgZzaKRr9I/PBF6YRr9zCOIAo+/M7H
47ojEIFRejfW6ZbZfRif790tnEW0N2D8CMCY6plESkr7TaFj2H0hLvMGbYqqz4mkz/1VLNRd5DPX
GIsRWJBPF2Vr7BN7hzm3DDq6v71sMsYBJcyHc1JDCxeeiQJHbbjXUgFk1LxC0mS3bzfl7wIJIIOR
nyUBqUU01jWmD5ICtaYMRsqOLl5QQWtL3JmpkAi/cddCKmBMzH2Kjv3ohlr4zM1JAz8Ka1HW9bTF
Kvys9xWj5k92nkXbpQt5lOwtfVvtyLpmjUWUoWVoboaRJT43W4zirOB4b5l5UNkHxMxZPLpm3CuT
n05oClPC9OUUFwztnC6Frd6yeu+Fl5vQuD36rg4wbHjBAefbI5j2Y+6MdqtnkURLPytAyUHE9Gq6
0szU9J4a4OGjLQwuI/mdpufJzT2My1JJdgQ0wGrGTq4VmUJW+R7mAaRzfIYg+aYLNLOwW393BYDb
wE/0jBY//XEWjexS0qqcbsYbJD3qNvuSQhgSRq18b//ZH49AwnJ7UBcG8NSE+qJyBC/MWHZTGZ8d
3IOclL65wltwDpXZ5sC+sApzmHvgkhambI608KnYsDzw3Hpp7uVjoxckSPwZUVry5mjoJo5UyX5F
yrzldmdGIcGoTUZm5jhxFUKarAuKeZ7SOJICxCpJJ0GQ/65SJCkyIzLzFRFMmCRxpUExf1XkxEl7
0hCsS6w7Y7QpR2cP4dDJbK9otQdlFNkx085trPCdidonzGdMn6q2UogyHlMFRBxKnq5Uy1iAlZ1I
TZtCQiS2H10V//JocGlPUERro4yzxECUgz+r4FoF9lhlSBemXdYFfO4xAyEIuDAOnW2mc20Mkmwc
lpsRu6R0XsUBhHOPvA0FbWcONgE4yPhSkkcdMaKP7EYG/r7G6+48A5t7ABKlw1v9xAsFi2psO59N
1fOgz0vwsadMN5CWNIwAUV1M+2BRXa2QRlHmZEJGj3Ktvla3LN4YOxqBIaGm7FkjsrApmhv0lF3K
MQf3C3Nx5c2mrrA//VDxrewQkcRwSosX0j/U5ThUyHz9Kc2qisARMksuVbJ2iT8qM1W9pDmPH9Kq
bNz4WhHHGcISGd013BGAfURo7HJA4iiXwDJ8tISGlWOAHdipIKsKVwyoRRNUY88feY6Ld2Nydv9q
sfhO1HuHb+OS0laYbn6DA9NLMCAqdCb7cv31Ze5UW4CeteTrn2PdeothFZaEJfnHvpgLcjBv9oDH
QHfgU05QlUacPQcxUkJiQ5+uYFWPCzXle6o7Ag87YRUCdmnDA+7Y8MO0eVMvCFhDsP27dW4+j2xC
5tcBYO6wSRdpoR7mnHon955OU4EXQxnB39CadDBgjQzPDZWX+wXH/0MaqEzxPXOvMb/TJPzPPCQx
ymiVoXfKv6d4VIU6y4FcV0qIpg5VlkNaJP+b5EwPR79Pi3RjSaTUmoWPNMSQAXN0x3d9OOjRAii9
80WxdWaiD0w1Q/SDnxoNFzzILBOijubYmswqmF/1N11kWlKCyL2qjhyesnp3GFv0chGXhyuIucka
x8L8OgqN6k9bey8tUmnTc88t6QuJgci1P5TaEztWK0hGx8LnM+7Ya0E/9rwX4q+YKsgpQV/7MGXV
d2BidT83tKmoIhKvzXlaehIlrSLSoNEtbsEh2+RH8KbduFgKFWcn2zgYo3GbK4OyDXGX8afo0yZ8
2NszcqwCwFOVM5D3l3J7QAnu2cGQn8R0jPPMj7N6487YzYi8+1vjQeoFUzWBOJXghAfWgicBnnSY
ZJkk1gmchAGTVb3qPLFfwGnRtP0qrKuBn/uCzP1oUVr5B9xWs1jzHhXa5q4DdJBV9OJTd4/t1yyG
l22cDA5nNTVdKzA4mQ87OkVPFZJdqdwNzEn19yb/sz5LNUowC8Ksrwt70PGBIub9yE1O6IT4NJQu
HeOnxOD+OpYGZ6fIyaIvI5gD3eTJGEImVrcVGhp0yePX0mi/MIJUfO1ZFK8OtXk6KpjuILccKeMY
IuI/vosN5pK6jR/Yr2L5bOZ4D6194C6eC+KZVUMGGAO5X3YHnDzL5pj+07WCFKui1rhOKuRm9qum
Po6T8e5roj90OU3KYHrqQ8GaNPkklTTiiqsWBdfBfPVO29lXh2bmaaGWk4nsY3AZWHrCsgF7/sWW
y4wILc1lXQVTdIzE7jBosTwEJZ3b14MH4HdQXhIQ6z7U9bePCIZ9rDLT9VZanuWXhhVB3bv03PSE
Q4PRxf2qcsYB7Jaw2b0MxBpMMlcs48gNuAMPdrU83HYJaSK/OzQDZaHNQ5m4t0lB8RorxeAqCekL
L7VyYb+vN0Sw4wJV1b+xT7o85le3fWTb9UlSVXfG3OutAat1vvHg2ZukLb1G+7L78VUWkN2vXxsu
p4VFQqcKkscnz+CUMaITSLq9SBNbqIhflKXzFX08rItLhB5apSdRXDoGEJyiUdOYV2oqmNrxbqNR
ws/7DbMuvCBC2UrO6yyJL7WqT4hYjC26HnDLXW7Z3sojqip99pkBfuZcj1Ix69ctsiiLBJmgVkMT
8c/8/TXSTuUrU5n981QOXrAV+MTd1WnZmlrDQwmnmp9JjdUOgipAtCt6D8Aobrqgm6WV6ze6Aycb
tPDgduzNd5s918uW+sM6wkIrEyckYPNC3trNaBnpsNkATfYWcXiiGjF7NLVjvQ0ZGEzdI+jnFN+P
DZ0hk89lMmrhrtfnhrGiyTTRnm/14XoDh3f2rKHLp1RTRnPdYa2NFpzzBSwsM9/GPwkFqcGPYq2g
9CZqB1EbP7echOWwPZOsXfmfJGho+PBe3AbP0Q9RrgogR+ahiO37i5Mm4xkrT/L8EJ0RdSREnRVV
9mRWnOclxVALQDU8Bs87l+MfIq6fpEO6DeEiEXe5oTUuShzmxKcya0gaopzUxp63/hTzpzLizaKn
qklpARgCXio0opmSY/gDWzv+dtyoy1C9HetzrAzXK56uIOgDON1gsUlSh7SbZdkkzpHRvxxlrRRJ
o87LXX6jzsM7+nurTp1/4vDhpcoexPNnBVn8xcAIEXMx6S7t/RmYDJOwB+5GtcXcskr0ZtXRkvfW
s2UAPlWJWJ4W4DoBNutcdY51vLvG2fgKCKByfu4bgXiQhoKxapOkpsgF9bHG02tewKUzKTZI4DRl
cG5osd19Yra2D3Q3HgASQAVS+6BOa9RNILUGB4/wdRWEsgwdbrENUGK957Ha5boTBo9dg55tjRFd
L5B+dLt2S690NrzOQPHt1bqQG2CA4sMkSKgR+yHkEdSIirgnI9X4U1PnfOoRFBGk9dZoAW4xHXBn
9tnYumspkhT8Usj2RNLXMG6fXubEM12ppruQbU/X4yLHe0tPOw1o/AYnhYkG4oVg+L0gXkRkY4xO
RLoZDbvwz4+LoP4LlNT/t2nAoYk4Xi1OSOUnqd9p3mF0TF7rXn/I4IfLPThumqgxILr2PSHe1DtV
YCqFlNM/pp4X+hsKMlKKjSHUW9Xy4u8gWdxRFPZ2dL59NUJNbrHloRGP2UfP4tC4uGYHmjLfMlCZ
C/kDGxEQqHiiUx7l3UMhWpEo7LgOw2zU/ZyWvobUYOuEELeOoDNSJO+OnSguMvCvldtgvuzf/qZx
xAGI5nELOPvMBVlV1KBWsbJmZx5AAhPJcsOCVZXJuw1yrzsdK/KI04+A80RZMSwbsgDDBZFiYghi
s8D5Bw+EjS25dZfCc1/rpfI+AmWWwwYHhBwrC2hwHisMWVL4K7GGYFy7CHYcyCuxU/Q4iKRunmc3
9R547/gmKfwV7cdG7JHM75woDB38T5y/E6ueyxpXVacNOS3ziXnSec85aywrmjhodFQlukFEK8cS
mB9MJrrbcc6Qa0y3xl4WSwJfobZBgMpFgUvCF0PvKt/pqltOchtxx1rwqWysoCgFKSyy+vjOPxuA
CV2UirXpECVIdUoPB4/S3Je45myjdhWugXj1Ck+qh0NrAIOaOOqD8UAZrCV0j9Akdj7VXaGKcUWZ
D2vf2RyHCq/7qXpRFJ8z1YmTIzUVefWZYn60lbXCJD694GoNIw7c0xuK9XY8AcHiOx4gu/0qz15v
4nkpIYzsBJxInQkkEsivEFturNVZ4pPZ4xpPBbbUJWRmlpogdt6JGo/f0dZkZPfxLTZc+DqEkQmb
UYmNGlt49yNiiOCTcqaf+hmyD2cs9IiBIDydhmc5vlIsZSBIWVfyDsL2B48xUz20XB84N0ctKvez
u8p8fYkyvpAlht7/CgCbnvcxirTuHB+4Qxxs7TMTYSFGPnPvvORAYHpPHJOnHcnb4w2EVtbbKvpk
oc30G2CT3Wpo6Aof9PYO4Q+rwMNNrZ6mEFMd00p2c9roVts1Mr1EBfF1w5CbDGI4kDDN9y/Wjvwt
SjNh8tPimYrwd6p7Xx91qiOovNXIMB0GQ0Z+eeXnyzo6dLdCOnexVYWFUyCGHcTGKET+OnoNkhT5
TRKbAmxygtHT41/HZ2+p/3KzyBCoBFokCVBqY35rv/Xkc3vMXJ0Rk+Fhxk68jdEiirpdBMkHbZXH
cItdEapK877kxOo9UWvPNU71Qbyuz2O6QyOlbAJaD4GQJwGk9pJIr0OHhAONyNzoJFBNzC16BP2t
irHX/GzEMpPEsitJknMmM4tYomFEyW+joU5rsMybkrA/20uRv4B62FonL8f13PLRdxSEFP1f8F2k
fKIzkBA0chBFExqXjvmzdFFw2ba0kVQR1Q9AS/71d6UWo7PI732yfsCFbFkjje8kK6nmuYYc/JEi
V1dtEg/9e1Ka0p/3zClVoB8aAJuP/O0F8P0Ev4x6oo/FfXdip+AOrPh8Zyyy0/ij4stmbUeXjXU8
q25oLbhITjzoXB2uiH/gleFTPWGwsHzOLMTEEWu5l0Ff8RBdhM70SJ+AgtruOtXyIIjZIBwW5a8c
VkQCvTVSbDYEgZJ7n9icLpEsjU5drN+d1ka2LignjCWwOKOk3MCwk6k8/r2N2m1Nt4KdFJ8cV6gk
ClIzeO8G3oKcT1MoLJ50VacjpzDOnnE540dyT1A1j5bi1xwWInng5TPVxftlt9/eP1QrQpeT+TbN
7f+j0GFtvxjiGP39kukl4jWFEge1cSezUfkgirn2X53JmuiqQkB/boMdId1R4HDJy/4SrBhOT0di
SFKiX5svpx0K4Uxoxx+4MuBjJei4n4m4AFRFU/ftUWBBWLRpaBfGnaB8lbJVaq/fVEp+xziU6cTC
UQrd4okWToFeyvyXtD9372s6cBImHYA1/cj9eti5xdoUDRDzSAsgrPmn/BEFptHdokOuNuRNnjQE
rmwhsROrJGP9OidtiBkiOo5URAsBe2NdpCazEgceoCPE1fRv8rGjPyJGx+TJ/Du9FHYZkhVderem
k7RIJMwfi1MVhpNygEe8f0QqCK+Crl2QwybYCErXjc+ZvjiKhIyJp2gtNDslvt6iEg4nt1MGY04a
ty0kRlfKap+Lj/YIg6UTE09iNXEmoR6Q/Rl8pnrCuiB36fQIujPGUeJsxERBngpKJwwVmDtNXS+d
eT6+MGayUrDMzx7cqPDU4HemYCdjlXsWLX34+y6VhWf4Pua8tExEZoFOsXWlv5fCRcw3qKOeaQrK
5dI2CwU4Y48m1c/F0ZTg84o/3mPnBkRnT+HzJLSzLsBZ2UUTdo1qp5MIAs0BY8ZhGnH+tbJgV5O5
n8QL6MByEH4COFQc9hhWihInNxCxYEhwjZn8Ci/e+uxLKQaARm5BG7mn38o+qNDzbdvD8AqVVxPI
GTfFzTMdESdkw+3K6wUk6KxPR4KbwDm4JLzGIirKpXQJSuk4bnTV2ETKo99wTQSguavk6zeh/C8F
Tu+o5ciOASb3533QE50IO0JMw/e3aywye3M8EU5HI5Zi+FEmduohEV84UYscXWzX/PeEWGHDlWjT
7kUo6Z8LbByQUwA8ggBgt9YIgYfz71LtS0V+0VHvTaunVnpfYSuKYzrXWmVFwfC5BVAMxlBoEYhG
xV+u5bsN4mf5+XmZLJvfMBR1DT+ZI9lNBwfhp39W0quexSuZo4HIp3mmO0fi1TzP6WxXmr6vWHx1
Z2WeqfAEqZldcihpfSwza7ay13JzKk2nfcFVMKFl1dTlX4hQh+DIwAGM+zTpj8+TLh6xKQ20p4Rf
WOfLwMBqwkot6CB9/vRKrzrd3UbTEcqs7/21kOAgvEDukLh4ZmTMTtG8vf4Y6dnrzw7535NMuuds
VAPNj+Wj6rseDSRP+i4sgLkzE4Iob8bR4YcfT1axmsuqvrSzLkT6DDrPD7RIiYonNu8GDitdQ2Mu
tlZd2Z5vcJMbdkO7AZU/Zn9ZhkOei3Iah6eZrUy3bYksVLyb0aQtqvhG2i8mBK/zYoBEctVnQlB6
8XH2amRkO9tuJ3FY0mJ1fK7idQKzUVUywtXjm9oKK9C5xV4ALolyyLePqiXDZaGxRnaXcVNzx1he
GOhe69jEzDkA+egkndLX+AvkLZiYRi75siPns9xKsPp9WGEil1dzMhUUvUEbPS9ork4Td2/Y6+6G
ITvDwdqT4ZHdRtcjFJCiUsDorqCIoVga8PSE+2wcWpIXJ/uRNTYmQSnfJ2b9Wyg4KwU+/WSMQLNh
On3YDZ2OkElHPVhcX1IrTwU9213HuJyUdb2U/6XKyRKZIzTBkl5og0kyvIZwKHi6XgfPvzvzzVek
lFfMqlUibF1/0CRWGIL8GzEiRKZ4SRCdtAmuh+zmca9Hc45xgnA97TiK6EuNzAwvvxW3BS1QW/h7
J4XVORQEgGkg0oBtN4H7IRUMNv+BYEcpixzbOvvNa+9zGCzM8/oTpach2DIlJqyt8YPMvaoRloYh
rm09if4HBErOR+aldblOckp644vwaiZ0n4/5pTqfyxSQlmjIQbaHKczbYAntI/VubsLkSuWKEz1R
VcSvLqbRUbWtd5bGlBe2ET4sYtnY5L7i0a/AbkjYGW1LAiGiBwA0cPLn0QcZ0Oadcx+HQw1Q+ryT
TubUCDy/PvMuJBVGE9dnYHF1Aeer38d2yn8Ns95UbHo/PXdadf+x3v3dKmfXNiUtzBFN/QFrDBkD
gwYmOlye/4W0ft7/4xumzLCchKsy9aP7iyDcHk8bV3BvCzmGHBtqUYu4wpzbnEK4svX/jXAWgQ8+
q7ex4UiyQEnv5nT0JdTxp5URH24G9B3o6CQ68xJWwNHCBPIHQ/zTjh09Bi1RtVABzqVl4p4AEQWu
Ug1gtC93MoJDXjx+1Ppp4aO+Woqo4rKLlYJNoPVasSdbiDMI9m0zvv+qzXFhnlm6G5gBgK2kCZ9D
vNf11wEkgFUzqSnJNhcrvYLXu94gfgV7YPH7Z/BvC6d04iUWIsrh4Dlx/ICOCjQlruaH3Z3Jk5/p
TehPAfouasI08weXxz4w65L6YrpOOJy0s1WOO4uo3ZPQckSVa2rIAJKEWNdTThZ4Ut+zrAXTq5BE
V2LTbl6WndFWys34xYDCa4ZXM3Q2zvXTnkO53wleZ9TmwopcWhhjLtV73MAcNMWBjYUfhsGE3fst
nER23gKvElPK6Maud2BrqNQz1lvHHlzvNCgl/qpEniB3+5nqMozU51yxkJn61lQ2qUpw+WpJsSsf
vLCky3AW7++jNDTN2qnudjLjVUGrulEASYkJxagg9WNY+66eNbnB1XTZLVk8879Um84HRxUV/XBh
KU7EQ6/BJMIEEXo4Kyti8nL2VRn3JrUAp1mdETAWMxkTICmEjvXRyc6MxwldTNrdk8Vu4v+74N8g
P8aPieaqYXpZEdiEFCnVUukQsnZ2zcvNMcIpF1w46/j670fdOW5/v12MxdGnpwKjXIYeFktCoSeO
ehR26aC3OfcppxwpHnaxRu/YXa+IuYtME42DiXf1GQAeJ8YLOgfo55QjP9m3OYvxf/iQ4a8P2Yxk
42OIhW2dVG6WUnfWvVDqaf8H2Ia1lgAYvV40Mghu07PGfX298zLXtxwWiXCVQnlcKxClBoy0jLGC
+Uu1JzMY/fR+sY1VFuBzvwjMmFnOhXj3JlaADgnklirkoi6+r1S1lkJQarmbb7NJeHKL+Qdm0S+b
J4uRS8rplvP4AJj8EQxGIzFRRsC07yv+49sZAZAi1nWBRp07M8McYXVWvsPDAavq4CahddwqR/xW
6WL+B8EoKukSd2JhDNgRKI3uzDeEq11SYA3iuYozFfFG1Xzb4R/Q2UdjmG0foAcNc2tPHaPGtYrE
7IZFSset+4UL5JnnAL5+uNxckAGWV6V7jwZ21hV4TiidFeBWd06Ve5Ry4IbEwvYPa9pZI+oR+lI7
LCWx0Sxvr9gINQrBawZgK6HaoGATJuiq6RDnzMFmPO19wX8v3bF5Ww4w4BTuWJXEnW3HCBFqL3W2
vnANY0syNWwy6RzMyKOd9vNg9XJX+mn2MPpyfIVfij7BFA9x1ydcEkekdCIDVYaDCavi9iU9/2tD
tfj/l4Nr7TOuEIsH+ADiKuUf8Yj3th+L832K8cAx7YWrFZSwr2wGIMpJ3gNBIz8uWXLf9QhFgslE
8AAr+nJ4n5mO5dUL1XNqzQXLPKInzwcftsI0OM5pIYPZUMz08UXqeU5n3NplTqVPcP/XgIwwaBGk
zKB84Pm6dugGTIWp2w90VxGqWvcjMdsY0r/2euOg30c3wogSqgYWywthDjFhz7s0O+M7l3WmVrvH
JzM/1LZM/HwbwkRmf2606Fr9Nz1S5xaEsr2g3n5EZJUkdiPJ3maPyvPLQX3fnqhhUtF85Gzev2hc
0BQP3LvccGkcRyx0xVQ4MHa5AmcZVCzGnnse1nku9xJfjmTeF6O31emNGnFaquv5ZN3+7g3yKz/X
WbjqrdTFByRF1ytV+pJ09pfqm5nF+6nU97GMg3WvCudW8GBgQSi3IJW09iLdvSyS3Gok72QB68bX
y5wNakTZ/Q1qa06KT0ypNFV/9+4y0MBxzfxlxDrYDxjd60heqzrPHxCUioDo1ztee087jmzeditH
gG6xPt8yp+8u6MeyeYQ9SMFNdKXqJyKX9WW2J83A9IKwVdnsOpO8IqY/rRfZmrAehb/9PsUiXka6
Zi/d1kU+IwajSnLrHuE4Njtf7LIj+24HpjovnxNbFZedooHWYLXLf4WhDQz0a56PlUEuboGzPuOb
hwD8TN79jFqSOci7HYK/utko9JIMTyQd2k49Covv1Ti13+5uGinw4u2Vdm9XIO9TV7d6UE/k23sb
G92NKKsf02PgV3molMlD8czh32HcvyRaVkQyp6aUkbb3z/JwXWpzdp0M6/ehtT3S2Y1xOjYeo77M
Gety+RLfV/lsID+1hdX6JKYQvNyxZEbTClTuqmqn+6GA9jd3cLWQZiL3iwkeB0TwQXiNEYbkGtr4
/6mc1bWYkyD2S8aI/ffCFqe0A2DHmW6VX84CkgBCEEJjkDi8vla8Zfj97khdc/N8lW7hxzczCrd6
NoqyKUEhB8gYin1grHe1kDTEyoOg6ZtTAPnKS1QgIF+LuF52YBG8uduQBMg4QBboiB4juEevqAae
BBwsewD09jGEZppIXepBaN9RcU0ZahQ3q1fp10LtyNjS5SZYW9gA/pml10rBJuzEP6P+pM0F4oxh
CvmvF635xPtahrUPHxz0avt1DpyUrBmQ5pyNYnx7aEpq/A4oD9fsXQAclaKjbVjc+e2ctBUmL9+U
cWkyeRGEmCw0lZPRtDsRVZLfYInLo1mNq8h/qrPoLXSWBSXkfts8CD7fGlxtW8oLmgUTAyavpkcr
hxZSYO9H3rCtTxIYWRWootOoAkP/LgNUzhrvq/wIchCSOGbZOyEVSek72vnXU1o8gM7js4CnC7XM
ZHJdnsFs3fpbu6WHJ4ueLNEWdZSz6A+36R9m6j6zI1OiFgmz7Z8JFPaI91aCqZMnfaiFP/O8nTV9
P7RyTng30cIG+/GcDtDFHttiZeJ/2NLdLMfHt5+FKBwpcLp1qPiCXCXboSMWV024XnAczFobXVVN
jukg+kcN+E2mtHg1V02ra60jUkPIvCHD/HO3QwtWLbQIT7KbaQieQS6CIA8JT5r6Q5W9KelEDAPT
zQs91eJW2SRoX3OaUdInSE59/AfUQY8G1WVHxOxRWSIOhzF/hdq5hfe5k7nk+PjiHM6hMjyA8wE5
plGGd8ivWbjZXJ8pjsizbc72vlUpOSexVOp7VbALaGeYg98ybhetxDyM3RNkA6gpN45DaVPNdAjM
5IQrR4TSC6t99/EvsjUWW/+KdkxV6CUJwm8+cJ4wy/qfeDlk4OIYwMSLYmw3cUdSAkUIppTmkHJU
4mqGqeeLL72uqM/S69pdwaj7LcoNNPzWxtZb1rQ8Dza64xry6hFfsbYtaEaRuyAcsR9QNXaBPUhG
dKIcwzyAv3VQFFXbI7l7sx7KysKchICvo4uZW1MMzimfXds6OnrW465FkeHYUPk16fg2Ulp1X3Sb
84zn4HQQ/zYsx403ehoJzK+WvuYJNf8FH1Tmzs9UXslwHRh8QZTDkEhaDm1XF5fPZIBZnvEljken
V1BtU/+T3PGwm38LWiUr6zMaSxdVMAdXQZki239ALGBxVy0ft+BdKPA2hLOw8sKHyK+eykErG0Ch
lKgtGMAQwXrEKq0u5EoiMYvCHTwlufXhTzJq3410fhtktNcwjPiBQpFPaNuFcHshh/yuMvyBb1lv
U73NEG8hHXAWheAZxA/+6P3czBM2SrVlajSpTTeKQL23BW7N0IkXih40n//G5kQTVFLzkKk3VPcd
s5zjDshGDHgN01df9Kf/ADXxMnDO6VC74rcHtD1Ga5CLFl4GyZ7t75b4BQa+H4IvnTGZGReafuW5
V00Ji7jiAzCIyxHH7Vj1ioXhGab8403fuhowTTGXh9aThrx7ukm3M0FhT7zHfGlVWygrmEQup+Mx
6R+9PddbPFQWngWz5xgDvV8PBy7EpCcoI3pxUQuZmUdtpMMnhKou51of266jMBcNWo7K2Z1Wzl/p
31CELiYwNzP88ryHRbYGifRmu0IvoT+gi5J2EHFW4Zgmhsc/Yo7UFTbzTGq1uVa0nCXkImBzod+f
s7e+9Io4PJO4sXZD4GwyLnkZVVfAyQHby5sphrNXSNkuDp+gDxXVOw9YKVltPzJj4YOrDKtjUzRf
k9v3vy+4flGeokTOV3HJmEzw7z6Cz2e9uU1z9c2XoGystx2nijMtN3/xU0MgyRqE/cf0ZeEMnJWd
MFooysFl4kYTEo2mltFI0BGR2dRgWeA5VrGga3gIFy815ngcMgl7nHchJIJ7YsyzV7EoBue/Sfh/
RLOXmatV1S/MvmxlaaozZLgkK4SstzevYrpQNdjnrt0UKUKPGkkHepQDnUZ3LcA53d0XhL6XQ9zf
tM68p0KBz863IWGjy03bDw4vZ2L3kLBJ2NYhjfKRGKo2NNWhh28Rk8Jq92r3uPWGbzN0/H8jopzD
ZbwwLvQzb3lNCaCtyD9mSY5S3nQ7bP/lbfjJEVImoe+6C+7Cf+7i0AyVd3Y6ScAModtGklaDtQOr
EZ2xeBMdn4Oj9INgG0mJ6B2YstQP9KEfLPdSy8x6daKwX4WcpN0DYd4bSyiCDmBeRNx7Xcqqp7vB
7OvAIaAhwz9IEORZ5vQm76Bhag0i1QomY6s//T3rdxO0BZEdHN8QuL2OO3c+ypplxkkIO2lGkqYd
egtv070TOYFhMvlkxGX9MOJu3C5XUkDNPXMfcVzAa1veNIeITpKR/9F9WOlSwOWA7c07RXW0xqCq
s3hXssIAAKLnu1dL67X49pyBFzKFT4dPD8Z91/nGAA2GQBzqNjWHX4El1QLOos49n73Pe/qvHMmh
8HgM8/iSnvwiOWTUULATGfShj4NgCY0iM5Oe2s16iAaKdHiQDlguH8TJcElA6hPl9ZgHNxm3UxSz
XEeR7F1QDFxKbzQmyVRPfZaJ3Ek4d76EKCrd3NkYePu0KfjDE/20TWfWfCzjYIQsfAvAkXXKCcSP
RuYc5yUxm8QiZYRojFc8dedbPKo1bf9aTRbhaHCHVbAdBrib2EjhpRdYcKJ2UITzBhNJ1ug4gRvR
Ne82MjfoUHY8WiA8UEkcEzLDfn7oToL3C++A7N4F5Is3K0jMMuS+K8Fvq631xw6IZc2tKn9UttaM
7u7lHBR6Fo+HEB/S1d3yWKk/Yy7O5CWNkGOuaimCK7FiyGV+0/w5SSvgFp5OCqBx6SYCN17DTHOE
JUb7ts+hR8T8Ov+1OH0Kbo4oqtkuZJcsYodSU8r/6UsZZF6Cwm94CEiPngOfWoiAxgDbS5mnaX1o
yVJLBiHnENlhTDL529/Ye4ji5pdD+zSgxpBFV33IooOAOE3Do+XxWr/ELkFweaBHPAg/mSPWo+F8
90hX1DGbYj5VJduyy6TvHYyXMm//H6Eq1r7VdH8rusbroM52ADDolu+4Nt2+OsxKHdM2SnhTqIfp
WfF1j0CwAne5oj10BIcOepRe+tuFS9fXJ5OyAIwF9za5VVs9SmHGy7Pq0vXFdtR2LT7lnfNDSt/0
bTjwbWey8HCMHLDVs+KH+HKINT69aSnc8uxJfSFQkEpox+zg4qAwZe0c83z6Ijq/hcpJwVyVwyQL
amQ1/706ZcnRoqAwDFfSohMSi25/Zn97Qd4v3rRX9vb3y5wJhM5wh+MN4i4P/RD7G54WmaqrFVma
os6iAVhLY2oHn6frgA+Io3Ossoo/yaq0Hlirc06AmYgPKpqtJqdaWp5hXiyUUUYABv5Sqw9+nq8y
FFip7yqh+PG4haFt3T8zfrsBURxwmgy1/oDG81BPJ3Ol+yDPwWvupX9myOQ9m+GnLbd2rMyLCKgc
l7PpxRnOZ8ePXsjRIQicksgwADWK4K8WF8uj/09TTGWu989OGxDqsBhVzi7LWeOgEsM0O3otBVlj
oFv2WC7zL68gId4ATm5luauli6DgGFKOX4kCiWX5cct9q1jf5cIu3iQH7UnfR8COk0wlfqPntE1n
K8HRxTiDKBeh6BUxOWK7T518dXvf/MtUVQIJSZTnTVthED5GNcj815l0iIPGpk3XiUEtF4Moy2q3
/QHiBH+EFhjdT2M7BTjdnklkMuLBoQeRWT7hBRauGNdsIbFCGDiUxp2uIAoHYwdDHd6IVm9hOgYX
UTMS3DyudefbaLr43u0vUnK86dyALKq5IoCK//Z7GchUXElNxPHU95MMWGwSm9pdvsrv/F4lHMwE
vBIrcjEjhEM1omoSTviYkKHm8tRoDdbNgx3L6NhJIg/q2TzQ/4DLHf0nCJammBrXo8JIxpHYf35W
hMi6Xv7gaMKoUEtiCbZsVpf9IcG9Kb0XuV9PTcIjSOj1j6SEEbbXNim3vRr9PAma0VgIHZixvzLc
0MEHJ5rtfa9T0EBigBeUMbiYwkqsZ5HMs1e7MTYaFe3c4uT+eMewMVwpt9MlXG5E2WgBQlBEBJlz
arweu0obCsq2OX4kNrJctH7ynyvuCDwFgGWgK/F5T7no4u/B4r+uv5nB4gBfwmd+rsNNcQjV08o+
5GK0L2Z74lhGHZ9yBukghKTzorh/QLm0fWYU8e33ITDYEMPkYhGij6u4DNtcftT2UAP+ST5k2PMs
wEaXmd0YXHg6HKTMwFHP5CPiMkXdqp9lTSdIWN12ZFuM5NsrEGul0hzIUPD9j2GtqZ7EPh7X/DgW
WFi08y7kmxAz3PHLmpBNmt1U3Tg0P9hNRwgpN+nVFI2smvR9q2suwy2JQsdO3pgVxiGsrzVi2Q7o
SOgoBwpTJFqllZxHbXjf791SkVp3Fc7QUQWWKLZXYeSFA4GFudLJ5O95OtxcSRNpR8V4E3Ib4q+x
sdu20UW3eESpQxpesN0cuFRcnwwzB0xmxMu89Pxc8QovKoFneYB6Th5djNstl+xlKc5QBQ80DZh/
09xnNDvL7f5e6VbYSZo+ZWQWo5cW48ecyEfPTXe9OUBT2cb7LKLuKEU6TgjlpgfzXYL2d6nwyEMF
Lk9+Wru+oIb7qFlxaJgRT+/mRhNLGCKfPeDXc3Ye+0RUhkj9D0TVfpEnPZGdwXXhXe4uDi30FcCm
AdZwn/Ct94RFX0aLChMnaiM3XF+fmxz5uUFLNYnPBxoyckoKXAR5UElWWPnITth0+owU0+08awei
Nba/yDAatGhL+inWuLG7pPKY3p9SGZA4gDdjr5acCL7jkuAliwazebZqTOyD9Uqcc90iwQaw+TJ3
F9hXWKryMVVrFnMGbSTUSF6dlnvH5hf6D1c6LC47i5iYach6Uttk1nkEghcztLVoHNXjMFhg/nQg
NX0jOSw9fvaRXbpGUxwwrs2t3BFJ8JCBKgSTHnvQqJuhK8GfBHF2W6oOZUCF5UdhfsTmbi3feq4U
S0P/ESS7p5qIOU5d7THSfl6BZNERMhStasZibeXsDJ09db9ieB4xB4cOd+zs4sRp6qYofmoUXe/Z
S3qf3iXxJCkrgAhrok69aHWmnMOlA4Mmel7D7YbkG6iZmEpMkcsZcwjeiABDd+neLFqN3jYPqn1D
oQBe1o663xuRU0xm8F7ugQKuDWg3ZXeVBlXMgVYtKlE6Q3IuKhRNwJXmL+SFH1Hpk6AtTLAxYotR
rAt2RG0ThY+MnckaNK4cLhDaZ0+1TdNcse5fhR6rm8WRj9nIjMr2xcXKfL5QuJtADPz+qcomZW+v
lJkj4u9lVk5uTEFzv1L4jgipHsM6Fd7sPCclmfdeFy8ogrorw4Yck5rI2cGXMLr92ODwnAtAbbLO
QpL+Tjy6rtGvx38TNUY9YT+5OtFWg4w402tZ8pUWFxblJSTuekHYWz/3IOy3LPVyOJsoqKT7+5TF
/jsdEQ6J+QEINuXFv1DKKjLRESH+8305eYjOtB2coDaU4UY/6/0wJmTb4eS1V16zsTe0l3m400vT
3BKR5hT9jpJswNQJdvHxsP4RSuEyK9oHHQhNbX92sxPS0BivjJNyTyOBbWg3ib2TqlPLOECDRuiY
5sJqAMHHHzxRMNSmiCfx7zfW78JpmbxjApqOlOReavC7RWdNAqcupCbjWu0rFXhUjehbMk0+CUSI
oREWvprBjTyGDlqWlBvvgvG/LRSdtkVrshnEK2D+8NuFufMT7ced+sc6jV3cKWaeJuP5l4kQJ+uM
isP1xVveN7JDMaNIqzoO5nsSLZWCg7meg7QHUnUPa278KIRw4DiTnZ2NCeSaYjaHhViZ2SBvDKsV
JiSpTE1nqHsIq4GktQR7Vw5BktHDhdBRbCilw9/1Drl/Cx7Wsm8Bal3uU8EIdaVr4ffC30oQYZRI
0h0otQzxR/sDO4Hd0/WUiFnHNt4vRo4VAhfW8V06q1E5xYbT4irF7Ddsn6f1h4MWnzysl1ApJkFy
MZiO/WA8Bp2BntPncaHaUDBoM+T+xACuUKKRaSDeDRXRsSv7Ur7GHg2uXgKu5OdDR6ws4eGdmEYT
5W65EsSAPsxER0a8PWJLgZJnp/LEeUY63LOjIZ24E2U+nkRHzcFyrR4Jmz2p1E2Jp/2+XbWMxj+U
8udHz7dXMmaSbjdzjiOQogU+aUjjywq8l3LrUQXhSMl6ZsFa8XnyGrLQxpaBtPuL8p//12DAcQSN
TBLzpNpYA+pPlHrUn+Op6I22fq3ldgXD5s819djLEYIJ46UFQkcKJE7YIJFuPaAgxIfyJgdCZNKT
dH/HeEi3Ere62tzXsvzBxfPzePnz/yvFcwCsN2y3bi6jJTvzD9m5Gi+1tEon4UPK8pUfuwI7ZU8c
BiKqh1dwpUBuUaQsYuaAOq23JmmOIxNMzv8EnkGFMo8Y4GbrnggkWXntw1HUsPiA77CE0tYEpUF5
McAObhlk8M8caGBowYmk/6CjgVwuygpvQgzMLPF0DqBF90C3cPr9Z2V8m13UF/QU0bV09OmuoBKx
EJ06Ex86bva+U2908MllzudoRITjBPtC3yGobhRe/QaMFdoGnq5UR1itCoAjGZ0eXA2heMJMjCaI
SNRmz9yT0QpE+JbykUY2dRW6LVCByYo+to+HkaLxJ4494wVKOqxSMopMO8XACBsjtp3UOQabrX4U
oGx9xBx8irAoo3N3rmE5BXxB5tjuT6hbt/bWr2Lq7IQ9KIAZyPrES5fMkCec6/VKegY0pylPOFmk
OAsTBdnnoQZcfN1denrcXFxBUX3zhoQvm5kfRxK/R4e4vfN28CDupqNN8sYYy3zp4sdJAq2VvxSj
mjKJGcl2juCPrtgs2GjnhOy1c2WC3c93Debg3in9YOjJIamdS8X7JLFFS7nE6VeOJUWRuvHelcea
mwDrM4BvyGkiVHhNBRNu6maKnHKqOrpXbbbwM617bzKrxLDILsfskL2R0kP9/NboRAVKAL4HaFQi
h/cyPY6JNaznJzLcBKfpz9i0VZdESnDwTvONk8DZYUWPY26TdEWsYA6DnX9gBGsoxmWHnfDik9Uy
EIFp2CMQW1po31w+8wuSoAWqbLOuqMoKg8NDPthi603mGqC6hu93csdnCguhKf5Y/KRafFwka5gz
OMUBco6QiA5JmvgZsm9TXuYmG/UNx51ayf43wJfYmIHvQkd0hmo9GGsgcUglZHqPM1BmylURF2m2
3BKe4LkSk2RvdbUJA+f1MFTp0u0GEqBvALqKkdLXs31peYGMu0XYfsmc6nwRfZoaNC0EvhVQ/NQT
0XD8WSWihdUnw84XI+vcUdIE/y8ZBNoBrlsJpDqzTebo1ZE4Oj4BWSoxQ448xtquFDRP48it6fHP
VLCHStVd6a8vfIZCNTolTg4uI1DEgBio9nWnwNkz7g2RbpEu54EW2y0/cPPdkeRQIy2D0tEwvd5r
xx2OYTcODxecUzl4VgGpTFVtBA0bKo462BEjtZPIX6xn5eoHJuwoVHQiZBy1qtIcwY6QX2FnBKEJ
wbLqGp4JydPfj6IRWPejvSpTMpXyNpBMvcZrzB9QRUczwvGfHYUTRq7kx73CmpZxLCxnVUGzUVK1
8CEtttsKHT51rlr/4ZXbhM6aeiZ8y4bEa967hQnW2a/kf754X2TXGUS9enEyhvmp/hXkTXmApgJB
QBEf1QOGoCxsACCopzfLYVZLFwLwAgri8LWDtU6vKej6QYFe4amH0oFLj3bh5zNKWWIMcuo61y3n
MISzOCJIvsPRj4EiecK/pJI4zo3oWmUkUqAbMKLxKkB0t2qYzyB+r078yklwkW116eFfZfI24PnT
V9PMuh+zRjGt9n/xJ+/+WkQ2aaZfNXhUtVOxBsGHcZVHrMKXyBW4qqHQH4D5QUZs6/6BsDOELBNd
sFbUxWygYcChXVl3V+5BDIF74df4Ad+UZ7Ccu23nUen8CtqNSgGrH7hdyIdDyB6Cs6fFkS+EY/iL
Na8gLmsjKLv+gODcf7MT/3Q0kOHBXfpkptVGhKBix5l/6Su3mYewpQFPmQTe0ZKQ+LXdLoadYzyW
k/tKqmGm/XfKj6hZQNDwmLIgOiAdKKdvFUQh6yQXdwBEb9ZlWHadMOHrl7zouqPS+bdMPtuD+ON2
UNDAQp69qvVRfOEB+XAMo7Az074hlXL52gR6Q3wVaoue4FIQNH/NNVsN/AEDytr1W7VX6Drv1iCP
5Rd84gMPrmX6fZRN2NtYmNIBUzUHJEDbB2iKNN8UjaSWQPknq5sr4y14rMyLwSQs8hj16ITg8ZVo
3YY8ZYsbY5NAMm/eKOb7KhDkb7uCvxFgEHlMm56OcEm0dL9TLmZkaBElwkRWv9MNOIGFrrmWU2uM
1J+Z6dq5QDv+Ljn+iI2yFsTF71SoGSGkpH5fBHGevROjb3AuwZPjN4GMZS1r0kzFkHQks6jG7US/
2/3K2pCCfYu/gr6SpJEiY4IcWKa1+f3wmAfsVcHun2BlUwnP04bX4fgUN2zllzKEVJCaFREtyVQr
MlKhRzkgHNZK9H9+pwp1O3uGkxYDdpQTJ3H2LvsFe0ogkJkoev8gabIbJQ6w831Yzxtd3aoNvZbH
N4ZWudJ1glq04OipLOBp7L3B2UTuvBA8cWwo5vIv8WuQCBE13pmrZxRKEFnNnzFlyX5OpL82JEdV
76/OfSmO/YPZXp1iXGOP0evmuDz9dY+pHMjQWk/bjlSzgaGQ927+cobC6iK17U0FX4ggyPjStjgr
v5U474nwwNMobhuaJLLZvpr36pFpH6Fygm52TJbgeaL+qgnwhjgqMHs4I3Vgg0PTt7J3sCVFpof6
euR6LYqPpIb2y5nk3Q7YUJVptZd8GK5enPsajN8cAok8NVxA2CSvQI7r6nsw7ARvL94+pFCR1/he
N0ffgxXbmMh7mggQFrMMobsEfGxUJdgIOT+Xtydfxjv2Jxnmn432h3aEhqgJVSoLVvTdubqY0Xjb
N1/+NjFJvWwGBGbBJ1doJN2gqEl3tBAEjC1e3vZzCLsI9Rekqc58K8plO+PoiuqK5K4P4fZqrTil
p+rVa4bH0gylpfwBU54JcrDqPbuiE3vg2XsRiM7gR0d9OpeITcTQ02t43DCPc/X+NztnrXGy8oDV
A49sa9+K8Dvj4sG5+d8WH7i1M1praxAZSxeSNrEJ9VvyTEDa77ERwkVV8xVGHtw9mHj/HQd6VTzC
GxftQ7uyGxT6d+EUeYrtprvGoHDOfgOvx06jhXNp11Cut3LyHZT2+vbjctJTQxpXJH+ho5421CLF
q+VVct7l/huJRmEGXhAenk/C+x8OiQzcw+1a0BFuBnZB5TdEcZmaq+bQkQ2JoXBjaadCHPXieLay
Ps8dDFNn8OJJp7GSaslOeVdalN/xd2XuBtTnktQDs1WbOFLGSKXEKGVsbnkMaJL0hAdWTym2rZPX
pn0X96ZJ6biyRPKDwTpQoXNealjbESDee+gpBOpkTc1IIbumbotUVsfSMsi6dQ/SJztS4LPZUnss
xt3jJqK18vM9/26I9/8DZ1mhdv3DUDjLihTpvx+3ilBdaip2DJH4yCAgwxjVLAdHIz3wtWgdB4s6
pyVtniTB3NtH2r9DiFUqLq9qn3vXgfEqaKgALHLVKzV+Cqe1bEjAaDqL2/A3Yh5uEga1td9bhouA
PO+RiO4kHzZixJ3bausOqhfKVdnNXj+DLaVHtW3Kd7J0mtKe7wZHd5CMGMcwf8rq/FxyHa0WE3QC
EJktqQ8NB7rUp3ex+w890IXLbCyVJkU6Z8U/FhtfWSSy5fmSgbHhBnmUGzL+Hexu1nFzLFj3hnqq
Dk4jokM3Yjs/ZN+s8MaDLZg65q3S2qBNrxL7FyfB81VBKgpjEUUOfcgWrWT3+Q+Kdq9L964FgWLF
mu7mhKmPjjwJu7d9n9CmkZ5MuXPz24XuhbPbWkPGoIHBk7ycGT5x7exfMwxgSekbLgrcTZcLFown
AVLc2lPbM66EcR6YwBetUx8b1xw83lkVPTEQ9lJdneGDzJNiFHv5ZTID7fOgcvFY4diz8sCrLxdv
z/JRxknwzbzsYip7NyJIM4gJUlqdLTTNCxHqBovI5xSj2+0g2p6itFuCDmd/T9bO0IETE6LWr9N7
1ux+m0WH6zieiSK1iGUfq0GYFL/PQh8nX5QUrL/mzKycjfzB3srpE3+N0BZUXUOp2Hy3irH3YiSJ
3KaCOTb+66y3eBToo4xzyzF0RpeuHQG3+imeFJEe3z8mJeZyUv/VnOoGmdwBzNaHhNrU/wUkSg1k
BBxLcRmkGed7Q7dPevxEhi6FllCqzPD2nm9mvjY6MeFxjJ5YO8ETaybeHFpX6lllGkr7vdOQ9+8z
h1s3Tfp4YhUJtyjf9pX+5J9NZHUDqqnpnnlHNxR7b+uyDBK3+PsVldLtZ7MzoYIu3sc7haZiQkkz
33F1xbStsnfj/IWM+wxK+hPNhuxI2Pdl3RaOz5q9ibZpWe2O+xDsJIe24MkQsx6RzyYXvk64dxLU
3EL4IolvcwwXL5DCdnNCrTM+rmdoKEVUaXzUF2In/lQMsuJGG0HrxoBbdATW8S0+dlre0uaTXrAi
EiPqW0eiZ33/ct1DN7zsT7KAVApTmxha7K/x9fII3obo04/Nz9gSIeq5Gc25kYnpdQJusBBt0DE+
hg7SovwzjKks4b6GlLNu6esTmG6MjQFT8NLJ2Z7Om8jsTuITit4uoEPLXkEqwWw5Edqw+IGwEamv
45S1OP3HcwJsNdl9fYE9DcGeLYeO/Hg1EUJ8JAlxdr1+E8liMjuu/TMhx5IdcHwTCd0+iGKRUhUI
8sPoesc8iOHMm58Ph6j82gf0EBduY55O6HZtVKAi49yEuA9TCPUdnJq75C2kKWb2AttAd+jS02m0
5VbFUrWiELsROsIMlSxCq73BgqwfHfbz256L7DM0jHzoEJw1C+sv9eGxxJA0sfTZhy5ShPaNezJA
mQfegQyihIJAfu7bD7qWIMVcp3O26UO42BYaY4xccBfrufo2BzPeKhrPXE9feRtKU+aojajDZI74
1z3v3fEYh+K8fNpfdN84GxkDxkvHn6StYouA0pG2Y02lOq0LsWMEBI1RfNob1JbIFZTkxd9H42Ho
174QFIi6ND/KMLqEGru6tp5oRBeRh7QtsXalcXOXAQmm0MhOqp4RtG1vI7r3GGy/1zX1JyTkTkBd
YMX+7x8cSJy3u9MJbdMmnsdT2jUZ6WGtgnQ3zf5tABz6fNk0nvXQmlWhpqgXMPxNCVzI7j0UzRzc
OmrJa6BCOeFizenM3BVgEokWbT63vSzprXq4hefKUStHuOGXV7UYH+/2b3eIjCZpJ04I1bXJFqFg
0ibo5kBYmXhA2YR18vt/u1AlmuqshdoO7BANbIx+ILhl9t6lciYsOXod91B+1ukn+OaT3KloCv+Q
ebM4mrp7KrItqy90bGqo+yfGJy0hCKycsqN3OC05SBiLrNBItUqoMwTN8hr5YswAIC6+1u2rFz+y
oL57ALcDIBYXcih8BEMg8Ird5LIbzq6y0yd93wBPes6+n53aH09e4BO9xnuHGqndWpOue5nllDY+
zR2i6LtiC+QZ+KqG7VjGccy/9btmMz51q0Li7AWcrHWDqXqJ8VgUzd1qvaoEDgtcHfO4RiV6PG3/
tZwvDEj3bFWDFHEOVH4F6AFDzdPIVs5kEvh6vPVKx+W3UbKm0ywP0eY5jVVcDCYX6rBvH07yrspm
WVqxSH1w33BZq6jzxTWGklH+0ovMloG/4yfgOPM9ypowqB7eB6sIus3RvWJozMLdHlnQKoDjzs1k
YR9FUjcBq0muPQ/076MRt8Va59AvR6RvERa5lwuqYOvmRgZgFtqYRLWtNh/NT4sv8fk4seVirHPt
dRUuUMXhtD5axws/1lkcCtnCmrnaeC1XJCrefAuq6/issuO6Q2N5TvKVgCgkEsLefA4qdJHGQOhu
9nNNhltVEnZDWFPn/+VdGoRBUfNvckwE2TKj9flkL1nRny1ayYVMl4NtBMnlFc6/btyuzd5Bekyl
GjY7yWxpOKY2Ol6t96cx7XWgNOuADUdRdnJvfOCwEozug0xflQz+3Ykz1Dh9wzSGfQLiNH0tjPR3
OiYgphH8CWRg1bqhKou7d2G5+4N1GSamspLhjlHO4jfy4PZSErX10H+O9dtNLRPbcbcTFK8xo/LX
dmkWrK7gV+BALanj0VtLyuzKclLa+XXAOI4aMtrW0zkd86eTXBs6F7wkU0Te+NZK9HDZjpJmvlg8
7H0fX9u57Xe6+rtJbhxrx8WkkfaY2UbDg2RLhW1r66QxZ2ZgiQpDQWvg1IUd6W/efY0VRiZPgR0E
gySyoLfu+nTAo7BsykpxqJVIyROMfiay34dHLRx2yXpWcrrbvv+TQ49zdRWzeKTQYITZIRIUGuk4
I5qHpJZ0/tZ5h145uVXzkr/qEg2V+bz+0gXLHj1LeBWE4+ZOyhREKiO92cGkG7uBJqo9cihBVhA8
LZdRQuSOEj/mOGy5wmnSYFMgE5qQFf4NQSgr06Aq2+/m/YePptydUv+/l86uohFFFhVA4YUVS+ev
lB4bxsAIW/F/AG4UVyxHSRwK+80yZNDtRLjqKBSsSXQHe8AAxNYm6B/V+cK5t/X9QCtr+T5kqqlB
zW7utSGqKW1uB3UhEzgRBaJFXvPQGQxrceYQxcLUe6nFJfZ+Yph82Z3/ouOPC1hxaF53H30pkndJ
q92ZNeJ5ud8tb+dmjGMqIa20FNU2Ec0OTf301ifoCXYjNjI0qXE/KRlyAAu8AR3nhnoCzJ9JCejQ
fWepoVLh90vTinAAGW3VwKV3cRwsWIgv9hD6VzS7cgJ8KGKy+6EwST7DLi2fIt9QYIS+sL51EIbk
IdIWD1PYXjGqw1CPjV6Xtla58YeXyIGhFncBXdxFsE5cti+lV/YWtPYmPpm57TNvMJogC66fHC7y
OvX6GCKkWN2WQBFNo6QWarYs0u4wgmF/AIC4zqBoYkAwuGRm/h6tt+2syM/DQ/gUiUZuqCOxrFBU
OODM2IwhyOC6xoOYyic/8eWB8FNDfxLoiW7jKHrbEkn1/6sUwx/RkQzM7ZMhCRnLlg47DnYaf9XW
C3WG8C41iGdWNSOtxlcqI6fLyAqgB718M78117CwU2dlvDwZI2tgQKg6LEIwkzcg8VZwtaBgQb9I
4MSC/f8POh6pgMM7uo79S99XMaamOT4+PUpjUzTFTXEYyBb20nw6viGWG7knDTr1Be+4rUr73534
PmO0Zf2RRxdn+qgSjXH3JDR7+zZEJcldJBERACYQphMl+yv8cbFs/WlS6+w+XcrKCT0NsvkotgL5
RWc0G7/DFWGx0YdNYnL5nIiwNzuY7AYZPIKmSlYIeWw0DqTSTdf2aH4MCgNY25SSJaiTl/BWN/x/
YpycasF1X/koJ9TcZ1dvWLBOlGxmdut7//LRqPZTm+ZyD6Ggzum7C9OeXpL2nh9pd4MbVr6+n0xl
1sNphDqjHJSsh2VIwlDyhsT7pe+mdGbkwKOZ3h3KNyQYoDIlQXNx8ap74Zj0cRBMIqSiaLkxfqnI
kGELp4tynIzPwrViS3D0k5DYTQkZuIMrhUEZEZqtHnMVBwB+wFljV5Ig8jP4LEtDPGrTnZiDrC24
QZNkHL1s4X2su2cooM4ds1CRjQ1+rptD6LwA1UOESqMtr8hrsoh8/uTrHDTFG9GLBD/+xfovjpPI
7lRttes7J5UC4Hs49BIobqhN5maE72mTSLIaGMUf/xnG2Vz7Q367g5fSI6CdlAG78LHpZQ4BmoIy
BfEZehdVdT/yt0EoZwElmzPyz3xdwwbwS8VLevWikUTRFmnERuN8DznGORWtRXzs79hbNANQCj9g
KnkQnL28x8oq0Gx90pXpaQyUAtKo/95dItXHQNJeUsES9DmbKNUKnegdtlNU3JAXgMBdxmMFR1zJ
F7sOzTn9x4L4LQm4pkpGB8jlEx4UYY+5ruTemHcNelm1W0uZay9/pM3aotylaI+LAHOA1i+flRS8
bPWYFjPFEMjAGQlqtFmhNfTgKhA8Zc62pe4ZUDK7elmKxJQ2rB/LSJptruxiWqw6A/zD/hYquCGK
l1nJNtVR1d9d68x++L7X/Ceazjblv8EkMp33sCbVj4dTwSDrHJBggMvNzPMgYwBVzQRCAFe+UjbE
fbrLcrEJ6qoqETT8gaF5Jfe34SCw6Jws4M7ClgJscyXIV6aw/moJrsoz0PYSydGzuCuMZ0YEIVIx
jyKgBiLZBJ2FuAZK5qYPIE7sX0SHyDE0JYt7lPPyAHU+NPFLGJSKpor1Q1wqLr69faxosP9rEnXf
pHKymn5wKW9Fl/hvFbtD8fJ6Z11GoaQpmXhaabfpGjdc8wmq6ld9PiDOilupWVfmvoxidQjQHhPl
WDLeVg/wTv2KulH+xsMHPmdGGeug9wO+hRZn+naeqnuiB8n/obTBLsQQhezsJP3FF492KxA8UUci
gG6xQk2c99S8VRRiNVEn0M/ZRhQEbkcOhjjoGUvrTe73GPW6ROlC45oaVYvL/B1yxxSmSO/qx5Gj
XUJOo+Y9+7W8EbzZ4/fYELWp6cKuyRQhhyjlUGqqf8Q8CWmDPI+uDUs1nzNm5ro1zFJ54gLkn0cR
abUDKoSvHc4vpmayw1dPop31yS/BrfqDffbkJMwFDUt22MOSaDAKAIafDeTkbu5bMHE0ZZ1tqZ4Y
UR50FXqa2APyM8kmwoHJWMxssr/tHOW6QlcGMOkYJua17ttNLU0Iz6/quPEU3UhyA8VKlnN5rXcY
otCWFSP8v2CJL/J9OrHtoTo/+wPClclAFjkMTMj4x9VW6L+BaOO/MDGi1mkzmJAsSKYVdYTjQHRT
CiM/sfzu5L1++KiX80pOI1iEAD8pwEn1BGe0brh+Vd0xb5FBbLwLfnXnYAxCZP5gI52EBvrTWoJi
X93dXJEYMvdA2Ybja8THrSpSiKua8ev4yDfJceWNXfp7TU8yEwrSaUqdgnRVCr05O2FPASr3JSeH
mB3fG5NVqoZJglm2fQgIlgSNgB6za3fWbD/mTcQTL19HgJp+m6sap0G8LPiIAeF6PTzOr5udh5jo
svpYO09EUEZ2cHsRDYRbJ1EWcXMu4tUnzGTMkxokfeiM+6mA4xJLXX0HGR0Cq5PGPOkgQmBg0XSd
LQRlk2BKDyJ42l2/dVpIVypl27NZaiDR5HqBXLTYg54VZQahVq6r8fBPwXFlmyKe3JqVL5ytshx4
PLCloQKTzyMONrq9DxTEwQQNBxld6PfmkLMYDWjDU3fQnl7hwx7Gc+xOoJGwZd4S7m7UNjpNAEyf
ko32I3pxijSOS9oPro2ReVZCGpJqJBjGmH9nj4UxzUHDlp7IZJLhIDWystkJe8FQctry0Q6zxMCm
ZTlUtgHs9ozagkLM1v1thh1U8aS8u2QaocH+CXuyjC/2hvqNDO2DQDJbegyqdEPixxWpjFk7BT2Q
9VseSL+e+9o1zYEt8Rk0jlEPRJSYLA2WBIp/wDoNE//KxvirA0b5FFveW9Pes+Gh9nEL/tMPWgsG
NZYTfDFDH5P/JIZKZLAXf1oqbQJ0KfylH9zDiihfZt+fQ45qhQlcMLFV2UdAvz6BoL51ngBj0Lu8
YU2X+eBNPIISAjTnO/CwCeQ+MLATKUCML9CDvSIC8q9xJV9m4gAL3hNiV3C/ihS4LA7rvFRyktwp
k3be+Et4652qGS97nwgDKbk1N0luMNi9tonob1FHxIOtIMtwZQaus+dgGhwgCsY11xavOQ4DleXn
epWUBxfvKOuYhW/mGeBQmwv5lLDhJX/zfdmvBluRdnCndIWB3qDw/O5mM54vPXjTlgYQUCsqz5Mm
mkW569XGbH6HNyUDXdXEuqrZxQ8JpB8Dt7wKRFn47Evy5x91BelcQ6pd8pZvaRBkLHAMO+mr05yI
lfgzOIm0iiZejh1e5NYgwI8vvqdv03BWA9BgWOI8IQk0iWu8sZzo6+iQdV/2FUXeemXxz04mLepZ
bYCDYLK0+uJ6zdSW8VIRr88yX9x3k9vT+0ZPjPRZM/Cn9wqYeY2LYap/2G5lUjVXKnCR5KMhnBNy
PWtcPoOp4rU8ZYmj2S//dzU2NfIOOOnn8TGher5T/LarLEMiNGHVoeqdJfg5oU1qLKn8t4UsSw2D
tgqDi91YJhsMQ0uJoOkXUl1d0U1Nlm5e4yxDZUQOHA5aShDBTNXBs1ZYjBVoFr0Nv09eNo0GWfwL
vDFQkl65d4edzl4kHMO4OHBHoPEpPTTTsyhseYwVEMG35cvNXell9h4bK9iIN+A4AeU8i6a1vgu2
sMbqlZd3spOeKGVj2qiSYyrwRVamNppsmjmlkzZbo3YcBMEjzBh5rSrik03JZ3mgXfCFljYwe06G
/VB8+TPzlW+Ed6MihhaaSxR0PRm65JLdmP4ComhMv9QgoHdfLCjLTTdvBcp1nNrCzYxcgZz5yEqf
HAofWfSvAAxXymvzeM3s63FNpeF+ez5GYkoLn8jZoUfWnreNKfo1iW9yBQukdGmGpb238zabJ40H
SFZZluHAqjcaRMj8w1lx/CUhM88Vw/RxNnXFVE5EaIaqX145oEaXcZcyRT795nwvZH/ppbdNZPwh
wCAeO0Qa2+1umUZDVpLj8Twoz8bOQQGyL3/cSXZNcQgsRPxLo11iCO+hPtZTis0VHXAxCYBeSEuz
nfii0T1Tg0gPTcZafpdfIgW8Vv80E0JNpx9c530Hki7XdlB5a7OfW8nqq6WgX3F2RNIOzBo0qcxQ
5/nUda8hYb1MYYzdh9/hbFPTPUYJxS5D0R8e6548ht6XKFBVeobLs5qIkk+IxWy+Zu2k2pQGRoCZ
hJJx5Jrb/9IBAlijMxi6sZYxOjXg/szk2Ts1plQlty/3FCDnL2PZmYoBa805mb4rvJf3YhdgyM2x
t9fyOq+D1Buy/vXE3st8u7pfmh3CAvXxkWAeDyazCFifVO2vKBaDj1UgIMO3cluCQ9srYafVezLi
NIp19Ixn4OCmtbPGbiZY1oOGRwzgV67+gGM7KVN3k/+3uicWDHHdPL3E6DgUsDVIFdX0tZJRCqPP
ANh43XmVnUyjCj5aIF+uLP20e5JAOTZTq5fTQ+qLCYZc7halLaVPxquk8foysuL4Jr2Db5yLwce8
vThJaaEgkxxZc25nA5rfjwrVo+0e/skPh9e8IK9CxivcoQTfcVo248sI2oX7AJfelFPU1gnfmq8/
5E3ZlEkaudvLfde5wrMAjoMWHXeWZms8wiobyJZVJnYh5jQOMjrU9aeEdKfrogRg+miY3Ns3qoRO
jdosB6zwpPuD/M6xh2GfOLIWOHjzF2wSUB9ED0wXTTVRsL0+gQdyoZnunwnODDxNhPkRL12Vdl99
CfMSJdwz7pO/UQJHnsrpAE1WDKCRpe7DVW9sdk335Y0QlR3nuiMy3YCIU0R+w8SYCk03wSv/dMJ7
ULF/UMrMcqUpg1wBSlhP9dLw1gTYNiXr9w/Lt6g9t031kZSfUsymfuzlIpiIIPM3Tl3dYtlryCnE
uvK9pQTrCMN5UqXv5En4rZ+BOcRziTujCYg+T5DiDmGxIXkgrzHzFJjRrVq5Kp/irPkANcV6Fbsr
vEAzPWHssxNu5mwjXeKKSBIhlh1CDlQd/cLyiSYYERRLlkAAriFewx51szNxQy4u5gWpyesSzL2P
Cn7dniTuNVvVfFhmSglql6UmJ6qLcS4+KHPbMbkjyyRIDQJAqE/upS6LHx56u8GIGCbT4mob62Ny
43zH/AhSFQVgdYjYwOdJ62tExGHgNKTn/qROY+5NwQXraT1vs9sT69u4VvD64UWaHHqXOBoYy3j0
B9LlgiGYah7XjfXcV9YOAUkuIgVcMUMI9Zdwe/Cy2Q9FLFuf9f9ZjYDabcz4F4RlfbkemcKwaj/Y
AaHCz35eC82PXPWgZGz1tOjUpqzVS9ucRftswmOp//OPtZGC4OWeE7GhM5uFopVuf3K7TzwHN6ED
Ov7qV1VEVE1Qt9YyZk1tOVg1aJsma+btb5CO1S6hXI8A8oyxfEhzGkf+1T+UKv4U8AkLQiy/Hiy1
LSTFbzF0mCyQmlC9hB2InR+xYZKqH2G6V06mDkFFPPxXtVLkeM+G99Y21M6COh8TgUA8kNdyIxM2
JwAptf5X7xvi8jOeBeWUTcGCCZOWzInm4h7XgB4VIR5lEs74hH4llZQ3FoCShvtGJ81kOd2wl7vG
iriCAl9PS4NMdaeDUyFRp6EQZy4eW8EUsa6OKRF19uz2k/nauW+5ESLBjnbY/YDrASfMvLtp9q0R
27T1N5YWXcrQMZmphZoIAyHsJFVuH0S/wap9y2APiRJ2okMfUMW6a2ZsBoFWmczvx0HRLoYY3Hfl
xO0br44OlOSjovLytBsF1YMetOq9ifg1wiMSSZ/RZqSVDl0/32fu/G00z5RmbGsfAPVIjijNrvv9
CfbMB0RzFpn+nXm/MSCkBKiSno8DnG1MnTdk6ARqSn6rLXBSCa7CgMhIx4pw/LDsmWu2yHL608Zp
UcH+VDWQnGm6pl741un/+o1DXKQsRFA5FXovpka3Jsr0QvFFOzQklA8Z5Z7fL2NQxGnJw4Z9YAoy
nEIJ1ATW8dWi7WK+r4rPrDWGlej/yDdKS0B6GQKKXIBLyA6AzQFqb+phS8hUf4kGYvQ0b6md375y
OiXe4z0W07KEPDiWHQKiT14tzmGXmDtELMxXzEefAomh0PYlue4WoFd2xdXsCgFhq4sWfTHpol4w
rnKfB07t2oPjNTI7xwGqqb8uIGTAeHTrcF4zLdkLoDxZZpSMyh66QJTP6cSTy0Z9qy950D6YtRq4
u6xpZVzRp0P7govjPFyid2PU51SYx+2jJgXF/GRML7ch4Y3W5Z/WEKVby3bUifoq6By0TmEBUK7d
VbP6pttwAs3EJDvS9dKtIXhiyHPk1GVOqT0bZ/EOh8FwEvEQlXJgh+TVtrvxlzEWi7KXiNyDKU6s
j+pEPRX8txdIJaHTikcUihoIFdpojsmdhCe40exocqmYpJxNjo44o79asWa3t5Z9UZMYW2bNLBuy
AGezn4hUkDTqmLPfd2ZhzlU2io5pkNjgMcduTs860pa3F5pqU4AC+2LO0uOB99PP6sXc5klxU67l
3/Wij/N1OwFPLluMmjAv1bdT9jesekKQ1wEkQHZoc4+dla+npYGJ1oZ5j+ztapqtFHjM+5H39+xW
7XqfjbKGhhjv69/wkIMz2GcMcNNLm7Y+k6mnJV5EcvD5z+enPMbuKyJ8yykjdB361a663w+bR9BA
hzG3Sl0NvT80mPg6EHg1YswhWyyWKQLxmAnsmSUdqPc/fNDZ+SFjGfiAQuz4UbGSbx1eGboLn/XS
eQ9kuJWiYUZJtccl+ZD2bEzGfx5CkN+EJMEwgCo5uarK4zaObFEAZB+rXTpv6uk3ixT22b6wa+Ah
hi75eTDDr6t7R1n5E5VbA9HvRE8XL4Z+wbVHmnyuZzuhwnuTqegFssIz9PiM9F9Wjn5GOURo+rYN
at9gzfTVAvF3URmM02dLk/wJn07Azt14aVNwpKj1dTHvsszq3LDoULgNq+AOrRnv0KZOgzAdDmd0
PJSZNFsQMv0S9trheAoYYh0jQJ5wRo8/BHy5lvdIKmTLIWp2NiFe0Q5il/ZrPFTHRNXGzMCTNIyp
LWivgMa8VQH9DXvFv8iJi1cPhnVgsAYebDu2nGz8JtxcIo3ClSye85mhSoaWT/pAIurAVqWfLqNQ
JyVd/+vh00u62QeGSp6cX2+uCaMi/USKne7bdYBMylgprmhBo30wiZE8vMOadWaVddCM99lLJZdW
6mbr/lAWDjfRjmOZqwr0/hho7wDKNacVI0TvZj2EElx+ffdUto9Z4W0DZyQw9mHEk5sjT1CC7Nki
D2Qc1LTbIFhy8QIPkK6t/OUchmpXCC2zTxeR+aQKrPF2aCVcbRr3pssMJYNQhaiBr49iSwSgy1Ii
Cxb9Y+IH/7i1SkhZ0dpb54CPAeR9sau7lc26vp64yBBGWMo31X3kQCN6Q6sKEYy+nyFNRPcJTirm
UzPu39mIXoJuyGehbCdW66nYgyH8yWFNZ3vLPTLWFiLgQcSFydGXLoqlLyn75tvQQ86ozibizqMH
nhtMMHL8qjx2y8i/d6xVcn4Jbmjo0obuCAzOLR8OGwORgE2nNCQDoPLDAO3JkZwmblsUriJUdrHw
Sn0190GpugkoujVaPK9AObtqjgqlBs6hsJ55YRH6vm2zhYzLVEbVaVZU/zPF0B8mzUa5lVIcLBkr
G54xAS33putH6rzlb2in05SV8VOiUmNKNshz/VClA18MkGRDoLFVJF4Rd82CPBmQQEclRXKPhAEf
3Dbba1Vmns3C08yNeUoMRFm5ITIDzWUyUcwfVbgSYt5bGNVB72zANjlJ5M8pu5PWevJ7tC4EG/Kv
TNNjvBYDhiUfbvKTmHjCA06zc7kS3IWhLY71RWTPI1n69m4CebL4sR3nUfVYZyEDM5RPpaUjypfc
n/EZy0ipJZaS4/VTiZbds0Q7KYIsMn603LntMRsMIPbmnVo8BedIHQDAGxEXVtLChLCQwa1bB6RB
Jm2vmspUDqMXNDj5cch2cLGcq5aHRiT3HMNLDTQ4WmmyN0mkeYLYJkjPeq1kyok8ky6mwDpQHQm8
24rFLtss6Lwchx8zvjUnqj5kW7QvzUzXthpo0dPsgMYezBJtdVXu5PVG+ZBVaOhGLdNxNH7QRzt2
ndJbDtKnEbFoO3JySSek3cnbF2HdfKhH+8Ux1ecS4h0yB/EOwkHjAPzR2B/6faIa16L+v7TBtvQD
9e2p042FDEn26l3jy2QjflTITPoXMw+8uWqNv1i4AU52WhDNldFwrjJyeE8m8UVRWfrocnLw0c7N
9GGrWbEeBi65PyZnD4fZcURAq2FYt8ny8XudUkxN5adY1QRJNwnwgpO9ma0icflout6zR8DipfxE
XHXeodsxzhHYIY16Bk7ixLZ4lN7ZFRA7cHcgTi7qh6+e9ByNQ6xVrqlfnkYC8WvpalAKEjPbkgKD
sDt7DWp/Ya/q8YTSCHU11lzXa5/HzVxhEozX9TYDnQ7n1Sb7uAIiMJWbjDFPgS1Od5ZaXaFbg0MD
7rX/z3R8bFhFm+knZNylYe4+KHiJ0aYq/yvyr+YHqplnMDxwdjWyF2Ai1PlMeqGYvhf1AkIFttt0
yYfqkB7xXypP9PQQTjQntHQ567J042aEnHCXNY6E1yEQNuJoP0EYthTwNVdPATRaIeylgiwwUZyT
wdJEU4yQcs4Gf1bPbXhqBQ1qf4+cFxLTfJy+wbfSj6EZci8GV/Jokpw3i4C2mojnaUyVGbamTwQl
egtfqUa7yMzMh1ofuSg0jisMLRFIxV0sTCJgN5NDlnTYhI50v+TiVwwgK9Y7sXfSeh7ysk44LWdC
j57FYHoPEfUY5gHCSRCNlwp4cgp2tUrcbv498dEF1CtgQzhtFROaAi3pztFTJlWwlSdwocuyMK0a
1ItOmFNCw/vlVepJRiBsQXdc1QpfvZL20DCjG9fvPSpufloVAI53Ap3uD+raIYHpR322M2WP9hO0
6fepIawtOlWumlOGkm2gP+fQot0n/IaVVv/nWV+burSygY/wCNbPDqDg6CgM/nOB+wTsZBSmBMUq
AaXb+o3AkOEqJrEuxP7yyylfE0mx49vMTaMHCJwMdYhuXzTW5NvW1hJpovJGJnTpoyXrx9MoUy3B
LTNMMTydUx9bgcUTYh7iP8UwkIphkhIVNLbSpPiQXK7EvQ4W/RIDiI464A+PmgRU+xrniLleZRkc
p9reOSpf06zcjTRaEhMb4uCKIwpo3aTd8yWiOAq7y2G1dsZi9QevorvImdmjFHkntyC/y0hDnp3+
hrOi8/2LDpTB/QUgLggGNSJ6VhaVdivv7kSgrZKZz2L9lFwJBCHrq8sp0zl8FcoDNpRgbkNUELb6
cbYz/LDGHYZRXmtO46TM3+cqGmo4/C6f49w1uNAkRkaQ911hYLkmPnPvoYTEluoTAUhuXIPCoHzs
EqZehAjrcKeHyWidRiu8dnpFljqQxUG+uKLNfHHS3MmSXBaoCdojYi5+w/+XIj39EX8fOsbXLmXM
DGihxAlgi3IUhEGdeaWXpMvLBKoyGSKDo2LkxQrMYldTT2+St0JPtvPWUWh29T6GA40F7ZPCUTce
G08DlbpS4+jedbYY2p5yIdCHIY/2xu/JhEZ5s15jDYXKg1Pg5OVD4aWzBWxRtzlxwWy608kokmMP
mKtpY4BcprczNgH3tznOj9gUugfmmRMFAX2ji9o2uN1ku4e33TIawjxR+ssE2rdAdwqCqNl+esKo
9/AuVvatZOIQkGNihYCs/rzFDsoTZl6Aw51E4oP80XC5Rt2oUxwvyym1OQSpLCW0C6sxP4AJhBKu
JigwxS4YLw8fwOuLCY0W+a5yqi2M//7wbtf9SoJqmI1UFVnvdAdNxpzEexaQf0CGI2qF/nPbT8VQ
3TVIS+iejpj3rpU0LGqpOHoPLqDhrr1XZ9IsLYEpgF5/sCm5YfjAgYF9gg/+HKefQqMkcKj99Zil
F3MPYFcQiEPMSulav24KIcecH4Yup3wf82K69gv4m2GwZ6iWBKbCx1YdUv6Rn88Vud8nG4a/vxIw
H95FI+NTUYOzeTAUO6ptm759sf0X11zs4GF8B7Kfwuxz+P96xB1kBVRALPar1VZDJikSRV3ETEe1
Vdoq0Xmr3y6BTvJtXCEf412B7jkRMg0D3kCz8tKroggts0xEg6tI8KZkhd+iobwV7R5jg5cqn0sj
bfhtTsPVNiN6JjsvrldgKZzdo69LcM5qBU44mBZSp2DhUjZngyGzEvX3M6qXkzfHubzwMDMfLIth
NwX23Oslb01SgRHFmJaqskxyOrKWV7W5XzYch0sgHGd7qfUSDJba9sXac0FX+9HJ8YDWBIhTd8a5
595pY5Kur99cw0ZhXQhjZzbvvS0lxC8g57n3hqUdH1BmLRE1wuYDDRTQPUlADIvLjZ9ZHwk8mbz+
kxshYzgzj6KuXGWxPhEdE94Vzzv/dRBjUS+l7kGCyUTsKTLWO++/jlUqmXFjgqXZcWQBMBQGafkh
wFrpEC4L7h0uHAXSYllP7Wx2nJx+OO51GpDjbQO156F4gV4YXQe216HvbKvhjBVdJrSdsjA+DfMA
VXzsUB5YDUvRyR06fCeKe22uf35sUKhILBGDsyUh7nlBsWIP6OGBIhP6a6tAH4osSa5Ws02Cs7Nk
bPF68FnbH6AgcRPduehydnjFOEchetUUeFPxJYJiLjg+8f6W8jEZ7dU9WCiPPLJ4XRWULPi/TtsC
8fz/Wcx+lQ08IyVe+OaLrImaXhRbT9iG2wIeCBllW6druuOjokI7yuXmprXIPzs/CLzKyhgDUxbQ
ao94F5BtfiBPmOhCAfMj+H3W6fiBaCkJHTP6Aq/oRLf4KKn/hzXxlkJWfnN0mib08yjCvZZmRl/w
K0XkzdzcvYyb/EwmlyfTcWK5gqS2hE44QBC0j4LP9PtCXabvhF2v0/gER2Zza4eMfZaG7rMejeqX
9e5IBsZlfHrL4MAgplxdPLRrKQ/pfmMLLlWUUEr/ny7q5kO9uLAYoET7uz2mh6itq3TpO+AFzrwj
gvA3ilBjCIqNlANRUturTuuZ+CYZUzxB5o3Z7sL11LQELpwNObPXBj/f0B5UhGCI4JKm4jGNULF6
AxZWlUVyFdG+fwKaDbjf0k6OyGkPE4MnYZwV+yn1kV6df/UNjgs+NUKNwvoUqieyQh71IuIoK3Hk
4p4T9P7h7+OooPGkTiVCajTB00Z6St2fZU5CVCwUAfcco/jG4XE8kk6ql29MWHNGASLdHTEMVhEr
wCvkJ3/x9hKoyYj0Ur5NzjZuPMKeIyvK4Su3FTsbKXuA/9cMkQoQX2+PKxJGmuPjpfdCALEbMRtj
V2TbuuezON7Bzi707Hm2VlNQlWsDylSkUxq5BQTciYB5gs1kUc4xpoq4YgIToaG/XXhv/HA914tg
bBQU72ewtAvyX0h2lGi0ExVCj4WBAM9MMf29PSDSI9xwiQmIm05AMHEZHHOE+6EDa65NQR2PfEfW
mr8u8zOdYp+xecUYWPcbyH43e6ZBjxYOB8JphOHR9kRM4luY9UiLLn+u9pRhMwTWFE/TQLR2Iju9
uDub60kCd1ZOHSo/TcNSVonaoQk96PFvHRre7nrsA4XAsaRvtu87bgi3T8Vq/DH4ETW12g4eyqYo
tjPp8IRV1669wJrphWBPXmeGA052U8kzNe7rDemH/Xp+YUFqWZbkvAaoruxMeeY+GE5uPHiL76/b
udJotjRiJaIEqPS64U4wchqU59Cvcr4BZT8wR1Z7zKg80Bqwjr4DMH6WxEMlSiNSprTR+vp5UaoN
r0D5f94KxYhoGFryAVb1QdDtgSs8xk6ccahm1Ggt+kYWLYowScnBdv5nr/NdSnaPLoByzOFVzmbZ
U4NzlIXoyFyO2ptWEu2h2/ph59MGU6jtVBE+4Fg55V5tVnTCfRWBNKMkf+lpl88/xk6zZIf8KHHE
Z8fcdTnW2e1l6Ux51vtti3xKMrBlkkio90G4FZXSgFgvzpV/QcgcyioAXSHBiMREjeZyydXT2WF8
ql2HrtsVDv1sC4w6R24BOZ5adW5SxivPtHOy0tdGWNuZsi0/tnBARc4vqtejugKip4RLNFNtH3m2
SBkImQfgSsWPEp7YWmkwNnnBT4uMaX07wgN/lzVmVkEqNUCtd5bPBvqRgj0KQbMG9nE7GrHdDpKk
xhIZIa8IpslyoOc98JDfl7ud+y3SaMQEPlu9jCyBmC8lsuD4/F0nEQQy8t0ZAq+7aW7flDNoLNdF
5ovjY1JQUzHmaN++iMETAwo8f7CtapskXPjHji+qB6sxgDlbSIGoiSynFzKKqlnSbwCGW+oxNEcu
otFjEwWwDYRnkVabnlD7pKDCvvP85uxKEDI93a0rg9IUkQZ1nAHjj55fJH2633LvHFRATfo0iiC4
wQUCjjQ6AftBO2opp+4jK7wGEcujjaTIqvgslJPEOl2nrp6ukmPLi/MYEamtwqDdBrBDUWsZjeCm
PUgir9mApXYN/uWYz29UrcPmVbEHNoSAU5OMeeCV4w0eBhWg8EFwKv0p0kFHZyfKJrwxGdE5AzTP
vgW1D3OMxhqiRVsp2tJKuSGxwoF04juNWHdQ7tgCgHtNLKaXCWn4HiSpSLbWzWjV+xyaGR8rrXrW
H0Fxs+hpcX6RTQgTYkCym89l2J7WO2BJnJHiN6bFzPrcnwaHFHu38sy1RDhg6MoAD2HRZFddzR/y
uZNnOACcsDnTN8n1ny8KvRssm51iZlFPrrrl3wISDx/LYnvwym9kl8zcJ2bSNgWq7C0r6vvHchXy
J803ZZvZQYwtoJ+XqwsQQDWk4eT2Q5o3kdGaSetkMfpdatY31lUFJMidthY7wTs/Rj8Bo4MRAtt0
VVWQ83+GhvLB2NaaUcHof0Hsu4Cs8ZwuKUehRzbuIbTONeXNoPLw7lds65nR3wEHt+bEFeILG4ly
kA1TMSaZy4oZJZbN+1QkWJ4AjE/eWD0PK6F16CpQ8VFaSdTgg6Hi32+iqE2HUGvidb7ACzsdT5kk
OjFAfWWHH/mfNnI4kqYRu+8ZDtN2I3Rcqsc9UQ0qqMPQiLK+L4db597t4UR6kIBj5rKICwP6f/lF
qaBoRrYYFc2EAdyZgVrLSCln8GWnc1fI73yQSTaxhcLj6+t2+aifT95/ndVcnn1k8GBZ2SWrrRG8
1R4ESPmLmbnkzGxt5VzcPheAtQGx0suzV30iRbWICMeG5y0bfZO27lCOEZh7tkxWoAdxYunW4b+8
0rJUIXRgoZSPQSTi1szwn5upiMc5bKK4lZ/jsHpQeKVROlKwXWe87auGw1lmvqEkJIeQvzvpMiPG
KnLlggmyrdItQH4FBQCWILqezBiV4OVuYQn0sfez+wFShRGmtFnF1QX26thNOM0J7PLTY4xRdbNq
HaocrMChGW6JRzw8SXYf6WnMmzhygpsNO5bMr1bk0v4sD770u2nTtyh38kya3oLnSqGushgtvz1x
D/jKGQQXtqgfkp6iec05pdzTyfSaymBsatDM+ZBVrOX7hxzI/wTtYr0Q5BZRtY/T53a4hXFjaJa/
HpJK2G64CItiDuajumxh4wXle6aVD4WEn4+xycg1GO25DLy4gsP4HjLGKQcgtLf9ONXIXWxUpxLs
ZWedjpri0ur+K8S+ZP6jGJHrBHx4HyHpukkFQbVRYIHsal2ZGoCKui+DotL0vGLSUebOmsJH6tpl
RuXGHfHKKBO9WqQ5eORdHM3k+iOqn+At2PICQIAOVJhCV8vbZcCHBCqiY2aft4kgSCr0SaSh5JAT
zZLnjSJc1yg2uduLh8RyCxQshembC9TFM762Erc3mgkcru+vQW67+AvRoQGwuWvH1/7A3YBIBQth
H5DVFfFW8XnQXraa1IBa1HP6tvu0JNLwP7wGa1cEPwrmRvaJRF+Bwn2ylQl+bPFOwKZosbIcgoiv
6okK65k3gfDZfS91AUATplGpk/2+tvnTSUWTc/B5iMQubKAQu6OzkNENpfC/ZT8ydwTh0Gic9T8x
yXMw6bX97rY8MSt3N+A87+GPW6+oTIXLtEqhy5f7AgazY+vnddph7mfNIHLtZaQRYcYokCODRjVa
5Kzhh7Ij9LTi/qmlwVT2Yz6SdN1xvqUS9ZZy38wQGtlHmSiLbaxfM2UU/5iofszEiqK8OHA51beP
8G+aJPUfqOy4sRnMLiXMCSx/5mLJZQi8Nx9PA6147yx0e0VQ34cWdMyz71VHECIKbRt9zGed2eKR
DfQUwbj6Px0k/oUWkTWm9Z0845R29iNPkopnVQSgZSzLG9EyENXL5uOvgDvEZexOVt/uTDXk3wYJ
Pom+DGR21so2gF7TawI10EVJxCnvpHCxn+TQYoE/cyYwiRSUOxvVfNEJccudCzrI4S/TW82SqALr
AEEg4Eqy1Pg/CWnkepNoo5fbCuJir4pypdw1bw0OnVFhq7AYAbYixaB7DPsqSYVkOq2reI8NnEJ6
0RyxuRwBBszS3n7kfkTTxxDoPSBy7vS8/coYKmOJDEjrDwj93g6rQc3e+rqEGfkpCV+wLY0jxU09
77a4k1wgsjRJTIy6HrQTT08szsTl7n6MoAgHi+Ys/AT+bdAQeWQi7eMr9FYpJiUEOgdPpWgAfqF4
V2t+R7Me/RVjIPWg4lGzZONN4YnTb/jk3X6dyAK+pU3CXmVwowm8IS/p8gPzI4AJcTjNxP+g+0Xo
S+QYBbx8YjDAfBZw4uIdPR3a8x/AQW8RVwDIGA5B9B2Ub/7qqbU5BOwrX3ValQKa0eP9gxOyODl9
nUUKKDNeDSfieYEy/IFWRmh1/1EHVDf2GmjmabBbHEfCGhlM9Ruj3hBKLLUjUOMhk6G+ZrmwKlWB
9+4BySGS+zIKlyG89A0LyXj2q1CPOBr3fyLDqzIXePo8juNwzsAGlNU0wSolbrX1+/C8c2BJIeRY
3O6XvEZkrJo+In+2KX742CSPU+hOD0asoksU4/exDdaSbgpqwq3JZilhh5qH75h5Ku1WWk842+7g
Wkp6OqRb3zTFn8Np0e0xu7hZ4JCVwpYaR6FFiY2FvJPhf70Y3Ufzmbgvhe1wEaDzfIo30ZUBja2i
ghTHQv/PY7luYQutWILZ6iQCgJTfwJSOC2IwQlZKdi60ErYqLEft37NcCIKrogYWVXyV9enTwzKr
DNidg6xC3n5IS7Gj3J+3rOU8UmIwo6NO2u5GiJxQHqPYTeCdloYu6h/ZZzyWBmBF57wzEdnYQRSo
LKq6HkvbNGwVaeqAI19LAOJ+f2T+KIIu/hIKzNkUeH7+oWICmd6VmqrLz3MadG4YTX29RWTgiMO8
0yglptiJbi5MmmbcNdcFwQc8ahYOUPBUP1FojsEz1SliR7DkEaiU+k9XTGXignPd8iAU8+85/pn/
/yvJsfA/GDXCrTc4kBfucoUfTR9+l8aWvN6zXXGcxj96RoXayVYVvxMWh9Q2jsQL/Do2D6GyKYA4
/7jR9l/6dqXLlBtBp80ywX32oQvklcZzOmdPlIzUvEN981HK8QvYh28L9WsUxiwQaInWCj6WQ7dF
Rfa4GxWB5ReRHbZxz6AcF0fSTbb0Hyzdqe8Y/40VrT+pO/dYFrV5zrCmhuZjfVeVvjwMZDjxGDbO
zcUvSORNdLRloZjT+el1STMUagHyP6wW+FckaULQwU7zTXpYGwoJoXhGGocnbTxkMucF09oc3rAz
I9+syosj83kMs6KlOkP4CdGHmW0NYlja3NRnA+yOER0qcSDvezmeMpaUwL/vRnu8xJV5vYI3G4Vq
WlewgGyvKDmgn356bVikaJv/ncR7o2Jt1xXUaPE2py7Y/IPle5Jf8BwRbxNVBaDBDjdSDh//cxvO
7TM+rO7wl4amW9xGPjPX4O0Gbepusb8uxP9I30f8feBZlW54W9GLItqIYu1wxkRCSA98LVOPrKPU
9lKdFFSGvctO23QcYxiBQFiCsZ+zIuprKZrdJ2DybaaG4tvpYlTCbY0OIpIhc4yIU1kTwRlS0ZnT
2IQN5zqCKdwUou2f9ZPXcxNfU7pgIgKwzHWfeoN/wuU0Yrlg6nRKv8mwv7VhijFh+vUZW2sQ0wp6
jt2x52x/XiEmxGvNgAt+kas/KPQWBNsbUbuObQl0ytwat4INpTv37xspTP7WhoOYizyBbVEWvWRT
XQbavBeqfiMYz0YrUMNxBOc1Yv9omJiF3HjXYSDj5QxkeTNWjQclUqQXUZ8w5vkEoiggDWpfHAG9
cQsdGMrkdKRQjgT2xVMxIGFYTdcZEHS0uTCWBjnA0/Vtx57V4z1APqjW9TfJ9Pc2UrCtfGydqkdd
YIUyyM2O58yhjp/UE+wkt/4F686BCMK7rIuTR32aWHJJHAXbAFkWwyfjpP+J8VFHgugVO3jXNhSV
gAn4q83adTpsEIxQ84IRt70rI3acJ4wdyVwrF/foVDJ0YlHC6/4h7IyxkrTY0+us3jYVf4uXjEow
uBzxGo33mjS/icFAu1V1PWIs0u/r3xxfLcWyhudEE++CNwSm2DEDpBxcm9qYKap+IS+uZwTn3qE5
8X9qD4WSNfhi8hWfX0pJI5uEyx0V/e5c4RXKc1HdQ1YXEahWqq/CFgh30nCDq5Lm3ZOniwkp//x8
MDYe4ztT5MDYD/jMUGb5v70CUXVJeh65rEUtGxcOj+0xXFhL3SJ12h527QS5RaUvpwUuPB3kRmb5
oJepF7QgdNmzLOt0uwPRn7eI+heoUaCPECreTeNwbr3Ti4AYy50Me3H+ZHLBUPbz9HrQnMhRCm7k
jsttzsEzo7Tzqd9Ldbhq0oyHBDmRaoA9lmFu9+4YMBmqpgOh3KyzrUp/q/9egnb4eQ2YOabzx+cs
0OSMH8q8yt52RoVdVM2dzgcbLLnZo3NclkMCeDhvzyj72ZZTCUTKuIHSGs6ModjFwzq8sFbCACB4
m/egqUQH6w7LPw/Y0O+CDzZXHRpJKhiw3sWHlVD1GzHWWCrAZTqwh7vzAcT4atGpqk9giQU6h6N/
d7ZRUwa4nLRmMtET3veofKDTNBH8FUILkdIJQAg2x0AXqMUbULrMVgSCjo8GOE1QD64F6IGG0zmD
brjPEhAUOl4cRgkNDW1BmtsFyMsvBk8KsiLNRQFv5mOf89qbI1J1VqamFvTbHiWxLdugLJOiSHVg
7qDFgcKHfVkTTuDzlVVi7yaiSAg7XZ2YU1VWvuhXpfVTMSaN0/me423er5B7sTr+JEvHFpBQmQ6s
54RoEaw3f4u/W7m0vy3HzeFw9vBUxsZ7G52K2Z8PzYxpqzk81ET4pIHBpPmV3MJsP68AedvH+ETU
Z2d06dyk3+ho/x64KjQtsoYgGkJu5CHjQrotyE9m9/qvn+y9c/+McvCYePTMtkwhLWTa3F9cIA8o
KQp4ZyALL5Q6zED65b45iYQgMjZj2DPkLps+EQYvC+agPgG+KfPTSx1e+2q9oLuvjQlsSyUTBkur
YV5OudRqtmLYj/e4P99khNkf7C5+0JUPFTixyfq08jKz+q7+pPHtOpzbewEpihx11KuHmAeBUq9w
95cM2tmQWXSOTHnHeEEsqXbMaB+2er27nBN3L1QeikEeegW2WKxBPsHtBhrs1k4CSweW4AWIh992
St7nmg56gd1mjvtgU3ANzKj/ra3kbe+xQ35IQtPUGh0xsfPxbof1SiLoMF///eZf/QwE2NSdsoPp
KKCSSNqnIpviGQp0XGNdFxp4EZVAfSYy8x+yihLPhmvWzVHg3Wd4ys4AM5Kk/pNNC1ZKual3/Y/5
uY1TLu7UzuLk1K4S7Om1IMxDd9fLpBpbwMqUV1+vbjMyO3YNRkP3DhWhBzS2b/oPGVC4JPac5pcx
O8XYAWpsn/Tkm4kwP2/VlvSi7omY/43cM6NUgansRobNJ6I3SdRdUmcaglUMA3RUkU9dU7C9jY3r
bZqwJkMuYOk+ocuVnZxc7C6JdJDbYidKI+seEzCaiZKC9DTuJP0m+f0VpLyci59Eoklp1RV0UdM4
2CtsBcVUKagjogkOtBg1Qw4wwLaRmiWEpc9VfAu+/yiUprY6aN0QCCmaQuGnWTQoIosDFNyQ7ia4
dIq1/1lNL+ZezBh7CBzsKh2F9wj2NsXdyIaojrg2JaXNd8tA2Liy4BOoCuHiEtfdIh4oPY3E2phL
Gb5+Rt4r3y8MOUEoj7SIisBC2J0fG6ijVEARtfCuU2yYCojBSoV/4cCzKEi58mgwjxBtszKyg7mO
2rqT8zjjqhjHNDn3jHKZHWU5OW/ERZGh6+U/7MCVKce7rkkpOmex6cyRTx29cDvA0DvJ87x8Djsz
gp/bvQdV/XDDZ1vcUFu1ox8cSTkffV9RVvnIw0CCpTeQkGfQ9/vRZnNrdY2JrARJ9zrgo6IJY0Kn
Jy6iXbwU4yt+WGbfdlEnr1KRfMiDpAozAWZrhm9cNU0WDg+xUEXyECs7tQsU/ESK/Wx815LLVb/X
xfv5uSrXEHkMCc5WAjhhylctCc99Z2HSux2s6G4ERvd7evo+i8A6f7gUscnDVoZL1w5l+de/dgfj
WqmAtwfukuzm/0fCIXCQGrEwZ+enyW1wmJ1qZZVEBz/YROEMaPwmlFxoYUxuAXLzeKWAG8wXsOI8
Jp3ULe1gqceC+VIHM/JQt4Zo58L8EF9mDKGGiEQ3xhxe8hxfbWmAkjEIETkovEhle5vTGBNIsArR
2CMbFynTlWYJCKUw4FO7VOX9u8k0WfdGgqxqjvZhCN/Ax0CDJ5yrGOejxuIiLhugFYD4RK+8tY9A
P5juWNNEMkmfZDH0//C6J3u1XCwRZXWyFMyjyFVqJTIsZ3wbtkLxMbJNzPseXtsqwqwlt2sZUWpb
9LA7fZWEwYaar2jmCuI4N9KbnpeDfPStWQIl9GolozHtwsH6O4j275HDCKozoov2roIMnY+egPnD
dpKauPJW71X87ecX9TuK2iTWc/0HquyY48ypvbJCAHsanIYkBEwlJvygdCAevUGZi4nYL9VFX1Za
e4tv21LFUbNYl/K55WFysQ+QZfuXTXVlBlTrqvSxaZEYQSvZj2XQ1yM5XaGT3WkW+jZUCY1YTpf+
KfjLWI2humYsb+r1wBbQrfK8gQrXj84cgjV7yt5vdbtk1DXj7HhInG/JWbidu/em06JKaQOSJWhm
Ct4HekHV2F2o8LT6+jqghLu+6zcxye/vaQfdY7cqBWszH1mhd+3grbIHSO7EasYemdtsp3vVRqO+
jPqR5rMeKul5/tDI71ZfqckkjoU89UBepZNMh/izaqYp9raV8ydLhtFSkKIN1RBdRlhv00EZeJ4s
N2rRAFQBiPLo2GHhRgQ5+cnz3YZVr0fDRHryr8smw7NU27JYHRKJns8CzjTCocrcNPDWKtWgvUJ5
LT9Z5fFnO5j1YV+Frd9wmML/9oY3zszeth2VBpOxlfEn1/Po+ZHv2MZwAJaE1fcBLtl6wSOuJh9q
Z2j6YsnTMYv10UQ+CWukKb5pZIaKP8L+gnzNnlnqSYocpaSfyCQD4aPdYWvo0Z+sFDHct8AuSg+w
L/Zj0TnnkCGEGRdrhLoPU3QBcutmwAId2m8Lq5adK40QU8EPlcqz+ZAe3LYgbMgqNXuL3V5c+Mvo
p/kzqIMyvp2jtKhGtqY2WqHW1grpbSmETwn4BTUErB0Ryrwy3rxO/qb4QdGsGjiWC5DhIY5eUROx
u5FEkRtczlQOtdqysXsfZAG/8sn3g4glgnePQIedrd3+lZHeABaGx7jgmcwGzI3nnHQfrDMILL86
y8ogdQ00msiyc34idGbZnxjrP76utCuwo/myuxzryJ5zTAzvF0h0XNwnrv8QjNKl0E5cTpvv8GA3
W34tyncgIaqEynxxKsRjrUlX3GHvMy2GjnBAMf0Uo0ZZGeiJ+yp4EV0n39nezCyZzWZUoG5NrNSO
1l8DKjKEHFGTLIuft0tojoa/F5cnQKXiBIP8LmearNQW0AFHUSRRd3e8105CbERyi8KdYtsdFUBB
YsKaxRZMCyTF9H5csMYh+ee8cmoRix+ncUFz6sKsjH3bPL8ELI9vrMjyjegDOsUNrcGUQI/7NTyr
LE+wp+s4X5cCNIkedFm1SqCUL+BD1sSnefr7Z/Q7zZQkxL/mhgU2tk7qmhQGugahjcRmoLHIhxQu
gXK/+vuL4l5Bh8KneYVEPKTjV7iugq8jUeoTKlq8u7t9cspEp+P4Iknz19yjS0PRzW5Ca1V0tkk4
TYxdPMdrPnnqEICDHvqtZ+whOw99qT7aRK2V+KWWbsxSPs9F6IetVl+ZYQhvog9fI5HTPS8hjL66
nx2G/owsfG8EHAboO35LXJcVdMd2RMhWKRR5clzj3KHZbSihzo9s1P+A3kzGHa6xlhb7AaTbN8YR
fYKENkZkQ3NZaPmA+NFY7dBRUa5m96dpOvSfol2NKX7MvN9ViLLK4e1r4+QsLxTQvO6CvGiIsp3K
paAFLSohg59EV4/ZcP6Wsv7j0a+PLL0+fBMKQfLs9EfS5tWG8b57ntpz5MSOS1ha6oNUAeShDwU4
Y+uTBqxMPwLRDJzWNwJx/1OqexwnpHiBJt7XxQhxfmirzwm9F+dU5U7wVKnukBFhtAd0ffzO2/JB
xJNyOR3U+rL0EYXVPUU5mrTkdWXgmpAkdPcovTLFcHHaV44Tvhwb39BqJzSnLI5MLIp6azEqj+vT
57cLE4gSvw2i8GVispr0NrnTYOEGBCzyGu7S3OHMR4Ismx/saNzvdKgaePgGJqXpFRsCGqqW3DRk
CZzjGbNq80g0/38s9/Wz6XkTBMdcQeGd1UdA1ncO5dI2zA/DdxwOPxhNsbscRMXPa+05meKiYGE4
tMM9lKIx/6ZoXY5BStisPnpLWu7C75kfavrbeyVqa2wMbHlAoW/q8aVJY62apfeMrCpTl7F4m88X
UTZkAiQ1l6+Bpofo2oZKXMqjCkzXwnmXQ3sa8O7yX6yArl3gXPrJBs3i6RLrlLG/9hdw1j0BdH6T
Mz3j0yhfOhlXUXRfeCVD7G1hWfcQjL8BwcV4KX9egvlApPr/5yhc3ATjBfSyD6sWbhtRo6lJPmmh
7B1m9RoC8s89s4HHTpBVuD/Qj1nSdbjh0aNdae6Ztc4zlIztydk6BC1r22Co3L34/XQwww28kbC/
Q9j5Vcvb9KtnLp2kGnpHTzRqMZAOsZYeqUJcqZJal+BIiGVhx1kiiF5hPmaO92FIa5echThww87+
9s1GJG47/kL+8Erdt9bE+h4ZBH9A/oKpc4zaH0y1NZv4emjmE2oFlpZUB42NyrOSyerlxwMRbVJJ
66iVNibr1RazTFZipYtzqRgtURSTEqw/MS3sE1lv/dz1VXoVwghuUXCrQzvdwdSSn5GCqk4Xlfn3
vRpWdBK0CIf0CoaMf9QpHd61C7yZmUGaDz0QVvzA3tP7q9ydSffF6rQsshCU/IuWMzUmgNx1Ph/E
nN0Vojol0Jtm7QDUIZmuBRoktNSdLmHrYqNEJmbMHW2jU9laaV93XCAAFCfluf6KuFciQfYwDEDZ
qlNsgb2XfeC1lgC1VMJ4lZPNJutqiJsojujZIsY7uztioM4cI6IOB2QJsDDBbo5BM0IhXsEpLoga
ck3z6rZWmpC4pZJKUfDxGXZH4OfVuaXbPexGK7ZaraHTt9jnlZtdycGJRCcpII52aqwqWZJZNKNY
tHhUsDFEvQj9UWekiXr9lwXn1WOQmZk8MJiG3WqjTkLiVXPUuOlElpl2Nk+LqUzlc+8Vbw8RCkUN
9IGgHMONzQaMBKMSNwW7+GMG4GljlvhB1Mx8cK+5JXXYAhIbjJVeMPoMpJRmYdMtUu4Z22nG0I/d
HoKPXChyzB21pnMuD0RSUwcNYD2McvzCJilAOcWJw+XRur4eIHD/x2izJMkJ4gMH8Iw2WpLI6hAT
2xzNCVUhrP5oegbdJ35UpYWQ1UoZrtB+VxhFg15LJsqdVp0cLvumhR45WSqQc1ZUAZMZSRVnQjFY
KWhurR1LBl0FAOy7ib4PlRSgjKWY05gypVnVKT3d6tXryfRuJ9O75ILm6bQ+8zZqggmioWLp1phz
CwXoKWbcCwFW8k6pD6rNhRLOd8BQTiTQViPI4goH+lxcccZ3YN01YL428vo7FWzSQpFGcpvUTPf8
dhQqbfjuE+2n32s2Ihze+V5dZKH/e6zelDTuQlSVTrJ08UhPtjaaeZ8yReBOdaKf+IKOt78kwquC
Be7KRiZOhRNGsf72xeZqbfV/QdBe0YclZZ6MS6xxHrm8h9XWdBdcnXmgLhNRPytuwBN4D9xuNzee
d3iS9mNGmKhinppmYDwpcMsnS/Ose14dZvKv82Yp6AxZc7LE55909/qkKIupVjFT68Diaw7FvlMo
HMdV1ZgbsqE6TzQa8KaFTfVWcuxqHEdVhfOPmE8pZlbCm8D6ASduD9lUYOpKEXM9KD6PemUWSLzs
K1EIO7j8zBzezfsFXeCttSw7SVtwcd6ocnD8tiyUOm3piTjbqyhwsw8u4P3FZ8BlQW5iSOPz5quz
1V+cWVTWZ2E8AiRW/yFbS7YoPue+LJYEBTPtljKij3irG1MUO8RKFaFpcIeQCUAEx3mlr/2miFtk
aduoLvjUaQEamqMnOx8oOlwO66QWfyPf+QHmKqyU5YSe4TA5ns/iEhiValpw/+qznzPQITvW3gZQ
3tpQ4E/SWy7WW8MHlGgHMKj/h4V6Ib+vWvc/6Djdogq5q5PB4XzO4i74S4FXpDyg8cTbU9AIydbJ
VTpmiisBbmHq5tJ1yOWcADggJKgVOHP8bAYzjJ7QQZYxqFV1fKdpyaigywyeeUG9iT1Hchi1B1lg
DZPlmOQeKeMPjMyRw+VrwNoReJJ5tbirkva1assrk0JeCivazrznwAyz3micHflz8ZT/+O0EdU/I
GTCS4kf5pTILECysogDyYAI6QR2KT+BVsvX+fQZi2DAlGb/9yZmSKoYOdeLzeKf1NZ7kPvFIXjLO
xIQvcaiOJ+EUwH4iSG71T+UXZc/hkof1mynOv8uDVguVax0iTh0ku+4ajb+Gu/f4xrLK3i9mQebW
mWJrWBRrWNJuGj0FINdu0s6CXUnItdRAWzD20hZxcnMmSCk+ctXtW4alazo0x7ax5Ce4dbuZuL5b
WVf+nfFC+a94nc8YsqXxgNFxl6VcGQ71Dtr5FpLb3azw+r+2uu2PDLZxZet0xNVWSSjiZZAeb77O
YKOwP7hiQtWYXx7/ZM6Kdiwfdv1WNw27a8ejog0v9F8XHimg0s/GWsVwPlZI18hf40vsA4dUDLBU
ThpO6CVCK0yl9ZnsF2Q/9UOfiQzoPyxOK4kQgZS7LOOLmVB5PiEQkT8EVC14jNVhAYkNAiRtPDt/
22zgG6NzeskOs8xikp9MK8bgJZc8VDIW1Pz+Nc6LoX2UHatBJ0GR3KYRAprcs8uYhvDIRbMeGdyC
t6HhGmUMPqh9ykTvlw+Ao+ZbQZHkhhjtjf5+wBHdiH3+NU8SQefSdl4uE8vXJ+M6RPyJZr9ZSvgs
nAWvgUTQmaJjfN2wWPHihftrNhJJm1BlVvr7zoyZQVJRuL0lMSb+AWFOiqPlt7Na3vS1/zBDBkNf
YNo/bS90v954Vv6J662RMt4tW505G64Grvs2lXQNf3ltnICO8ruX1EEqg2ork4AkytodgMajH6fo
KuFB31YhqX/E+ntn4lo3fmPPX+F+vPN28MskMvgMz5FpOIrjMgJqyW0rXd6cJz0V0doK6OxolT+T
yBERy+M05HBJijYyhn0kAvjQslPa79dS9owH4U96wNFVdUo5a75RmFh8ioM5OWtK2DoMc2qWCzXN
UD6LbLNkDiC8mtiAeL01YCwdnQ7e4NogvWjmgDsQ0zGSTTtu+WJjbEwecOxTekFwmEuigleIwBup
Hu7bQM9x9n/UxaNlJFPc9BFUZYKKouuttF0a5V57zMQLfvAknYFOhuMV3a2lxFPSgKyn5+CZwWrB
6N2ageUvXa7fiQb2AbBfeL7BubNk3UEHij3ISgcbeQnQHR9JAA/An9e0JjLXB+AMkRIvGo8Il1jK
qNxyLM+3efkb+9McSHsonsC2uGfNSgyEYGsYg/PF5RD7llRGhGW81PpY8dpuJXVkK0Qb4OQTqiZ9
HFZAKHgL8CoEBXCsAjk3wJWeHHp0gMNndbcPULhfaR6uqlJ4lrtDtX5KsrbVxpmkPWTjPylQGiwd
ppNNcsm+MaR9Wpqy0SvJtSKXeKODS5hVX2EdAVi6v03GPB9cMJmm96Otyr2WaZ5UI84QbbsinWOc
ranYzZhMxGkZM//QpWP7Pt3CokZnWuEcrdUEYj3m/5AlZOCIItIqnkmmac5Kvrsa5wvUmZE/u5VD
D9ZnlZR/KUr30lFej2MCJ3+4aoCJR8Qv09wLJxIWsDucDbx2B84neI8XRKbvRWuU4o2VMaimsEQp
ZyyU7sHlKTLfJnyo+gOiBAmWJ2spdNXsV2+Kh4WL5CSspVX1GScHFly+ILbWfTkN7MEbd/AJAIbD
MjNnh47l+TbRYD+wGMx2BuXGm3BGnZJmmlNvEn/PumFc6D8ku26dwWSb+bf7W5Nbq4YXbJKQpZ6h
DREcMNaVo6XgKT8ytRcCG6OKnwi7xD3u/xn2KDByWuNbc3vJjCCCZExAH3S5viEiWSbEUQgwygqU
1UL2exwzfj/AHQLkszMrHxvV++NZJr/54PL4D0VX9z/AKk9Rd1xaEvpmua0lw7ulCWyEZkim+lNf
9j40NUL1NWXRUm6CW2zH5K6kcAXorVia6HUyKwCj380ZpF8KAeX9iS3r2mRjYR3LsGautEFSnWZd
Iu7woBD1mLKijcxIIt2z5MHOOKSRKPYjvnToXaa+b07D5mq1nSsn/0Z+h2IIOuZ4K+PMlmFzubtu
Lac5VNZUxIwdukym5BTBnXl1rXm/eNr4Gs6IExf9JWSZDCpZWSCRd40jVFJqX+nXsiqiJJpEa/Uf
eU/2gxh9J3k3HCgL2gn29dMDO5yyZQq5sVQu+huhtyOzByOlE8R5GfuezwuqdjF/2f/+zsmS9Y22
Q4zE0upbLxuqkS1xn1Ra4JK3ZGQYkFTBoWQ6cYjXWVkuMtTL01EE6qfJLYfL95opwKXfgFHRKlMh
7u11dAGWg1Nem09JH1abFrMiAWqCsI2knOPs5D80Fmh1YLsZiRDUIqnrMFm4rAf6rd8CuYcieHvR
E18j6wTmh97X9WBtAIwcvGtimftNGA628HPzNgJWDVrga02plfnwGBjXC+JLtHKLuGBy762zBU6j
RpbyA5xt3cssF4LWodQ7g0+XVzK7YhSudLBRqk7x/RBnY4pgR637JEyDAidWAZI/DUJ5BqVQL03A
0YkidsKPFl1q0HXC3qy0EQT8VVyUr+tXZT+Q2RKsWzOrLN0TMh2dadEQPhP0AbKcf2SXPB3S2EpY
Z6oq5Yw5o41rcIrByzwwkEPfcNxlyf3h8fpqURaiYuktU+c0uzsFw9xImdJWPbbDY+qDbQPCIwu+
8W8TYFLV4+gE6t6w1Roe66YQ3TYZFGpi9XTAC2DbutXj8GlXU8o+wzF5bZuKVSKk76SrI4P0yG3y
+lG1VlJfQsuwKOeeu/BM5dfK2DDa21YX9HinywgyAMAsCtxkl0CU+MKldoMqXjkzZSy3aJ58SsYn
fahgTmh/RXQgLJiFm1ce7mERKFzzgU/D5CVLsSleRISvLafj8GNA5rE4VyDxE9q8sEVvaALOubya
jblIjsNEDsaRZzNgx3NkactyHWsOpAe83dlbsWEQsU8hzpc3vwIu+RO4EtrPFEmAA5mzP1X+ukoC
A7/McnZ3idIUnai98sHt/w0cvmQ27GGhSM2j/TM3y3yNYSvSIeq72/x5QuAhlwoYiTEiiBP0Qs2E
ic8fRbEDPeOiKCBmXMvJxDMC0s10rX1XdMDW+KlNYkq8ZMA9jkJ5s9Vt7dV7vNTzIjbrsCfflLsF
fmI0be+ShMyqxloayYJUrKO7S0v8OvM6ZxejtavkOG7qhj+JtgZHjvFns/6ctkiWIqKzvVitDE0C
g/XSaKDJsqNUjd6fVtszF/pVFGsnHP7PIgBmguxSUg8soRD1FkWi6SYX+56p4OQqZs4+CnXeEgF7
rpY37btrFElQ3Bea3qqxY1ZuM2BmD8c+fIdtQSR9qbLnEL001E2ETBHDEqFVgW1+KmjgLGW9qWm/
h2MRJcNtbdJ3kNNlYrYh7d3kgCXrgZZDK/Xcd6SSx2B+BxfQwF09I1C7sgR6jcFu0Wp3I0RtvKO8
ZAcKH080Zq+wLV5TiuharOL5ZD2bhlzSwydOSuGYFEfoMODHQRwNEgq3fH1oEj3yItAHiCciK19E
tAPCZByvzMUuy24ISpsS+h5ovSe219O7uYt0amw1Ee1nU+Y1wK9lr0pqoeTOALbZnErQQy8kasA5
RAk5uwDUNzFoK+cqqAfmmv1G0GUrhaqhpW3DS1BdsEahesTjoY0EiDq9LAT4O6QIJT1rNEO/40bL
W1Os7ykWBR+/o4Bxo9OOrSxxH0sXVv55Js7wVzP0ZtZguYG1Ct72oROzfgPeaE9LiHfMtPQoOFej
d8/39RJxavZ9T2431D0h4TziPT+dzJC5l8IGa+g1SYDWqIMdWj0N3hdMNBsogSi8G/Td7FPRbL+O
KACA9bTLL1rdpVyVo9LHW7Fisb0CvjtP0Yq6HZFQi7NdPcjbXxzpS7Zw6PWULldalWOTee2W/THV
e+g1mvOmOLdkPkQKoXw+//O0/FfKbkMPzJGwO9sq9TzvIO30KgG9sT1ZoLFZIjNIxEa2WRtp63rL
r1SIS3rOhxHBcrCD9biASAPvOAIbSnGxja+zxWNAyFi0sOAADNooHB2ERNFSJXByN8c3peQrjLBh
QeQmcvsalb4KcTNJuWJEE6jd5F5DRQdOL/SlElwj5U/TXKp7raofUO2HP2sNbtnt7u/AgTYirt1F
3qh1lRGQs8weHGiD6DTjCVpsbCxoNbXiKecYlye3Tsrtj3EmbJvCR00gtFcoCxtrm2vDDFhDXsIM
W3/+e2M+Y8HM59JhDGbjycuCano1ftU1gdxxqKKSZD3kjj+qhQRQOnZd0/2I0azsXUcqV/g57A9i
R5ou9ZhXfRe8DZcz4/BDHtvu2K7ax9bl695+UvemCyRd+lvHSjmwbtHpbFtDrOS6Is+FFCBUVTjy
wPLS4QIu7XizBYN1BfoIicGrilz3giVYQfQjEfbIUGJcucJVITcVfN1Thm8yWXfahzTk3y4NU9+5
ilCsNU9SwB7fr8WQUUsGQILJio6oSDQNhwk6I3LI24vC/e59LcuUt91zS5eAmfjd7kolYcpaZTn+
mN1XbFQGa5sNdrhjBGwt3mkrjNGOHGQhXLmKwwAv4erkK0osD7HxGnUjYdU/6LSvrh4+WpgAV2kt
xWb0rnUDjCm33XPf67aahuqh3otoqYdXV6ucV6lwa9Q/8uO5w7akd7578nYQvtt20dvMAvOQF+u3
MZNM5I0q6GHiLyY30xbDRl8aAjmkSCOYvMdTJeXXO9WHlHLg5pP/WWvdeEp9rMKGZZPYMXqboHm0
FiFYu3IrMXTmS5B1/qmM2tp9KhvF1r4ToO2RL/0fzDlirQKJO8iUhM/Vbg3fnuiCJnrDQh/bA5gP
kwQGOUCzVw8V++8T9yvLlC6A7nH5Pmo3uDGUmQrQzXKXP4WuZSIZVlbC5Z8BYEEyNtH3mvkOSlst
rR0RvgKKovV258+5z1/dvfsERQfBYcxTchAJUJs0xpQmmLDt/QJRmcALt9VFUqD8jxm1loPWy/xJ
OHWbOm26zOhYUlAWGGSZsj7M6B05zLTjsS1gY7x9p8QcrGJIpHzXPxrPo8B8gryTX5IDfs/StkMD
MBQF0uekPkCqMHWI1W4yoW3X52CUFDB54LASvo/qn3gQV6OFXazXvX/KmkBnjj25tymqZrf9xFo6
IW2gpAfPKofafewe7BhSxe2cnZn6wkuV1NBatXSfrugCTAHyn7rRnkdd3DkfzYeNVB2qnCvtgKpG
6ZmAtVy8rywdsOgPdOAid9BBD8Pndcn+3B8yfxjkvyI+FY90ZpeObPR4DF3Bzu/BhGUVET/JyCLD
nxX8fqdsAL24YZ1qKc3FsLEE1eF/fG4CzJXw1OPledsDnvlLvMx8WUP+AG8rD4NGeYb7P+UWJwoN
vHlqmxDsjqbsSIn/LEAn9P+XldOkEYL2R+zusRAdVgB7Q9eJQon798rl4QxTpBZNRHH0U8mWdLU4
9ZCJHEWHZbpqye2R11zvapRkhDL1fsslqyJqOmdpX1ToZFQ7PujcRdanONe0C6E/z4Ibz50pSZG6
IAkD7mbP+rMQ6mRzTseQF+eQI/pg3IhZpJvptwVnLsu3JT8qBkl7DMQ2NMm67vEiXxN1Xryvaa9A
33msZGRe2s50qBZRYwMMYPcpNm2Y228WDkyCyY5Gq4nUo4nKfutdF4RhbFt+4c9uH4jkQF5nJkBC
SU2FmSmBnRE+iyxFP6wwzVXekyOMQ/GPnpTzKYbDJvymcbES2Q+NUfM7TDLU0OS8EoaqmmJJ26uc
4R/a06NQH1zcj0qPzH0YYvONLLLyYWPQ/EG31+qyXjZrsSq1GhCFlOcLMJHnsIWVo4JpZHrCZkBI
ip6ps1Wm2A/SOlm7x1Dbr5MbC/v3v3WWTmz8WYa0UJ2t0cQJQ1OmOWq3rwSv4R0n9dN/9v4VDxSX
NrcOuAbE/odQmb9Wt5zoFNlYiwrgAR3/MuF3dzouIhgQkvGe4D+sEtDGkK5hc0TqOtAlVVXnxKrk
CK/OmTQx5Reg6PoV9tQsVX+QCsIoLVZ4yqd0iErC2ltmiEekYnB1fljF9deyNzCF1Dmw5oJwoUL1
3ms0Y+TTEIs1G7LQl7FOE+fyShHjxCzAE70Zf9InsM44Yo0pVkWztPEh7UcCgCgYRMOxCUbCdITr
Q2gdFHL8YNdDeAd2YVGv03+QfF0+tkrL6AFZc/xQjm9j2H7tmam2npiphnog/5jqfhX5YG5QiDdv
OUJv97teUZohiExxRLNSs7VBmV9tcfSGDT9OxfJDDOQg9cCIO2c22WW33JX9nuLr5/knRr8m3LRy
CrJC2px766aohVk+6AKhdu3dDYGR+hOjEzJayZtRfRLUybqyHmOgn+mB52HdnaNO7yxeepFspT/L
K72mnZ6btnfbc58NziBSm/TrZdTFpXk9CeZXXI80g5ums3B8JjIBDNcA35OIeh9vJvknZgjIKdlY
xdGKc2rKSVg4XbUhVcO0DSaBa+4oSzPoZSddKje+HwljKnLWBbKVQYBVMQfCTf1wMT/Rkf74IRkR
fyrOw0NgMlgAWYIMnd76IJ7VYg1OlCJkLjcZPOA90rsPkjrD1Edf2m4PehUvASWJPGcpC8dYgd39
FfAEfdrxyOA2TDpDZg+eR0SdPfVXSizoH//IuR3BRfhItaNXBe+vy8Wuf4KU0Y6e+j1d8nM+z+WA
UGas8I4/JQDc2kFiFi5R3Q9oYkIokL3iS2XGD6IDkWtYrfuI0wKlW47pI8AlEroU7YwzDUSAjOaN
oMw66LXcSWTXFERGZHGTZPhNP/GlnqsYjFX1L+r9W1+nReRleIIotygWe/yYVCY9pqbDhgjbzyev
w4CZw2GBlXSfNgJ3dzJUNXDwV/4OhqVy81lrxcdN/7m/NiINfgXjSca60hB1EQtNy1dPZHeFMWgb
VnWyIuyBpizMMykAd/nPzzX8n/ItXkZKQvdFdLXjfAP76ekvTpI4NrnmPTVcMA9s2husIHl+Q8rp
H/PXAzSMrKoDBUzYUa7Ms0USZAY1e0pdhfyW4Qy48LP0Tzyr2PnMoJUX4OFujH4/SBYZk4VJQRLE
ZZLc2xSvbMtzWviIZa5IIOiQdKFM1zlLQc9Azqp9w/Cgs8+SjIeI9OrsjsEgb31IGLDvHWtSF3y9
KihmIfHuU19jM2m2M6j+TRJEA/Puimznc/PTgQ2pNCFQ25F36AZlmdJvjZVg+Zcy/zeUVmDYCPn8
Y3s3qEwCA0nbuvGFj19NyxxG6d//LQTgDDirCagdAMQtyiB8OPdSokbbSIuKiQEoIiFmRgY2jPLF
GggeY4r8YJn11RgCLEGvqgLfzDwdn5r892pJO55/Drhp/z4Kay+HuZwBWLJaHiq28mMJWf+co88t
oC5jcVKVVQ9stOimRFq/jGxlSZMP3GL2pKe0XfR/VM5Q7Um4l2LT05NcXO9i7+3qDf9T8Qu+gpxU
gOrditodRwFaRn3hmEZlpYSKRIyMJ8lJWsFO0SnTmTPZuhQbnLSqUY5lVW9XuGJ0irnpGJqwtReu
xxCyGTTY5sHrOAOLJf3RQIiDs1cHhd2ZdpYiRR6pFrtjl0hNrJNIHs1WZnT5YS7N9vl99wfRe6Rw
6myc4FEclyU7KJsFzdIKZpLbxZeiKjWBtEbY9uP4IjE/G0caqOlq46lWUxeSes46HYASl9US7HH0
0JNeCmRAMOhd9IOGKeaQlS/8zGovKQ3rLxpQ4wsBJlnBZ1a3epOonF+u5ThUq/7rL3kqHeUFQNDJ
Ynl8Po5EOqP1T8E3uDQTB6AiQkKWS390TeG+cBcVNxM1x8CtCAQtv3Sq5MGQ4A51r2jgVOlE8jhA
7Zka6e3MTfUyK79Fg29jFgEtXx0dWy8i8Nd0Tcbzhqe+Cwqjt/czohcu/pqyw4I+UpPfZWIRJ1O9
+duCwo37v25CKyt21r0Fz4JUyvnEpbPJAqZ+jtxDH/ztY5W61YU0ztMrcKKr8tIoXaBS9ujcew5X
eGLKDbbRESebFKi+SnnAOKuEz1Eu0PDieRsEK5LaFZsahwuY+A562uuR7IjJji2V4zAQ1BCSXvDs
dNz+fYhnYmRicsYEaNmdxzggDelRND32j6kMl1nf9g8FH/hmUPUjy78m80NKz0pUb9r1e9TU1DU2
RLbvILjrpDIlgVIe9ccr2d18gDJzkxUN6pZuAtVTugGT+rPT6emW7XBH451hOTPNtOXbS7zTcYYP
egmu7OzgZEdNbpOLfy0upFXHMvAI//aUxcWHTa55qDd3qnVbHGfCPvw7MCNGoTY5lLu0dJ3qgUWx
dTPOQEzBPrhosBMuNcWFc2IyhhZ+XGQ3eB9ApCZkLnPNg64mLi4RFuoL8w8mM1etm6KDxrm1Tuai
jY3ducKAaIgedH2SumG3VU7Dt0cEEQ7bmOsC/cC3fONZT1yjRdv+yzVqzb+Is6t2vopDM1qL0vHC
+BaIBPo4yqaxb58OUinhvcU58gk7xZqJNTwiHPBH6fcisLYt4vH5+B/nMkAeZZ5eFoSeXBpLwiZj
uAYWqmPxmg9/eFDrG2uDw4/soDf7HfY25biZCYCsQy2TXBZgIltzNgj6frb6VuKzXFnA1CPTFzAD
JHPlo3XbLZKRoLSUQjioQEK7llzgJxLhUHb7i09K+ovS1si+SMCakk95Mj1yNk4n2f9apv+iaxbt
A+Z+kD/w8OF5TvYD6ngV7BXqJJeOawN6L+ITO0vee1oghcQJXJVtlLLeX0ZasJh+fdqMORywqq9s
RBychHHL8MaIME1dhjFbQjSWTfES/ih8v+ow0bNssQBiwMq72NHEotc/xWOBzG2uS4xOFN+bCPQf
zW7TU0ZSpAf75rXmR8EZHBoO48uX/fN7evUnUNKiaGb7ELq1PfSk3eKebHwb7eygH6KdqzpcCxI8
UOWEeousSz//3YQX/ELbhT1b3b2c7iS1w1ROww9ZVWCnPFKblmcHgwxnaoLBZZiYgWQs/IlLCvIH
/ibFtK7zUzEP4ccdy9JFyjFh1wrFmJW/734ZRhq3Jg96CdzESCXsj+KO5SOAhsQ7xO+Z941n2EQY
pVVr94L6eHWvcOWFZ05jbSeibj1ijw5g9GA5xjGLqCX0FKFRDU1qNa2kBF1dzHKd68pU3AwK9+fH
GDJWA32O/JVVBVQgP9ml7F3S0Dwz4qjGLpyOxgbXaWMEcyXhtWhlfjyIcp8/6C6gZHjik6NuO/fv
sJW/oMBju9PRVTUVbxJ3rc5Y6NusTD7deUNnP7OYr3dwqqeRO3bJZ8a4G45uXW6QymuwzAqeOeuZ
TvOmiXNO/jYMiNkKh7Nc90ORExM+tNS4CgNA6NNSivFdEfWy28IsRI+4+49bojaiGQRCPOiTzcrY
I2OO/k7DwHrgm2aMmrdauN3SHpdoVadRYCNy3eAqnR/Yw4SUVNgEaSTh9meAG0yeywCbZdhyQ9x2
69ct9+NLEtq0iLUsJrotMYb5mcDbKvFPsrczQqTnzyDebIL8vjLJWie3ncm9Lup8qkOHa27WEQbS
aXdenliu3fNzmn6gVM8JpkoDk3GI9nBRZoC0+MGm71q7KYWnhS6tOkKBXrFfDUr58rll02eb3wO6
HaO5iNNS6YzQsl0c/4tLW+9Po1ZOmuudUzosQZIvEk+rdFNVHJ3wQkz5b3KGuFT0DIbnpdy5Mx9D
IFoAGbQ+tG0YZBdmZFycE9VuOiFQEB1+D64ej33gUJraYx0DMrQA0Fg5jjBm7BYj6Fb9VNurj12v
ZIPMpB7DkjDsXws3wh3GBMXrzu7aY/0MvjhybyBu9TuDU68iQiVWIN0LXekBeH2btGflGKH8RCJU
7hmW8Qsgt3huw6FJXmmQy4Nibo3ebPoFwNu1TmwcoW1bFhoVqnPsUtvX5EUErH9IylMR2IYR0Bym
0Ia5JVyAqHmb7G+OVud3Lw8dl0/y+RiNvWQMjiMZPumezjjCv/gszAGeU0x7cSVEPAycVU5eRFZR
nVz/lwOSjIjHBPd00Vz+5MZg79rDc+P2ufL7s7uP5vQPGEmAn6UOAw3+whLejvUgczyYb7l2420R
RyX6NY6X+NDOodZbv8f1xjoY+WKWayloWM/GKPPGg5TZ0sDz5Tb/7li2ImcpNkKtTsUHk44jOIa6
h884Cb4ecnCGb+cqSYo17xfb2p3dIUA/fSpF+3zaA+dnVPkHoaraDWfih02W3gKr469Q8t0a4Gtm
HT1AadZpR+8Qz1J+B6O7EgL2PDh0ZUVBPY8CihC8w0YkB3vgOdyd+jdjd6gZcyugyvdshpWJQ9i1
/w4c8T183zRkb5MZy9/ZbfpDISB4cNsBOE3hf8n70u3WLN0EWMl/tcYoLt6ijiNnK3zo0+MGwwGe
HyZTpO+toK4xWgP29hlhN9aYzfIqceHpF0rcqCrizp9BEcSgH4QB+C3C5fpEwgrsN8LPfAOZO1OY
E1rWAQsZwdzGorwIh1hlQUu004vyS3wYv9kQ9ugNogVjKSnNf607gs8NUjo4puj7a8ohuKwGucej
LwAQll7W8W57hCU+Ku79Ksgx5/u4Z/GDqL3Sma9u+IyLXxbMwANMFGhJ4uEg1eTxAlp+Xv58fBN1
Inwcy3kP7F/xJ2xJD8QRXG7JJ6muPxuIL/x+ZokY9lovIaauvkjsYHDIao9EG8xkyR9MXsSnnJUT
Mk09mQa3X82wyISBfiXQwnBFv7fHiLnntzpXAViLS6yt28CLVm7CAGrMyFoM3uBZb26qeh3NATg1
L1roYWp+Ka0H0vZgSUFDqxM8mEOHc5latRObc1aSIuXLiyOWZH4NQhiJRZ6+YY4sUGIshHq0Ffu+
jS/TAGB7v9EjgcEjd7hNeql61qEDFgwqxgHmZ8Tyva4syjITgsgSFTpalbMPsEaIQybt6648avFh
JZ0IH9/X9AREruGRE8+ZaqRlX/kzmesQjwglyzM7GsJgZhzAA/OztjdnnsKnYz5XWkAGj3s4L1H8
UsIwGuai1XA1WVZC/ms2IjZu0ZV/AyKDgDYKBztWeBhtC+LgdDO0Ip7HAD9cH1knOuiBMncTtZfb
RTqWBVIoj6xyoj1IXtJe3xntGsWmfeJgma9TzZRp13SPZfV2ZddgyBiV+veTKc91jt9bVXpGyAo6
CRf+l8izaDoRp1/rvYX40ab9z2KdroUgbtPnasojT2Icv3Jp1XCEYKbE+O/uTb07Clt86GN5mnq7
jZxwTQFEb03C1ljJHMnGYlPZbJT8N328f7SlMBrsz4ZxmTobvaX+TzBMBk3KoHnCH9R+OK0I10lo
htbYvRO9KgD6Mwlc6mM1gJr7yW2FyB1fgHDDShTtz8S+WZZuYgx7Cdb99htUFlwVjs2JunJOA2+c
2GhbIkT13SnN3nmQoREW4Jyp2bgv4a6bGypchm7zy6wm016lYF9E5lUYXXHf2olHw3vo3HwswvAu
Fcugn0xOkm498J+Sci+LcN8dVSJwV2Q9nbfOwVogwSTDXJuEYSKxzTZ6XV0pM/QvpKQBnj7eCL9y
zlvTD9nRNjFF30LGAKaAvK5cp/ms3zSZA8s2jds0jhJv+d8xEJ4IPpdFxh+fSWjpYBvsnUR2C3fC
yilzNHHxUOlLr8l8QFGYoCLatd678F8/0HgUAxuAtY0YBaU+6rAOnpXoDkQ29Ep2Y3/aqCR5nus7
Q1YhHXah0ic1Z9LH/MtqUqggwYKtpyozsdIYYYIC8PQT6cmJedr5q5K/8zi+zgWZ8MSprQt65F9m
6cQupjK1SzOVexmCzz4ueLs4PxLO1r5zQZMka7R/zA1jg2Df0PyXQusfG0fRJHC8GCuTKGS+G3qL
0vPn9o4rCdLS0gRmgQ/JtvpGZOtbWn9wQlp95Jm1IjqsQC7HSbtOX5Fm3zcJEZUtcROgo2HmFkiQ
oNoxisPmo9IMkFMHG2Gckuo0Q2EcVy9d0bD+tbiSGQlUJHzeP2/++uEPlAaBVVFaliHkWqYY5kYL
ERxJ+h3Sp4E3lBDB9pQ9n9IoZyEpretjFjXhe0nXkmNW/rjr/KvFfF5HdsTXgUz+OTC6crRFP2ml
vXmxzJt1Yw9mAQCva5Ec6NJwaoVq+PaFQ/Tr6KpQfpIzgF087txvV/7XCSo9dOrpVEuntySa9diB
KpHE70fGLg+YbEVxYDVV42/UQGpfehRx5RKnDnKVxxAqrQSq9VlUNsqK3gOfRfu8ki5lddqQoh6Z
mO2gndcZng+6qHuwulQb5YmQMBPLlVT/hDY5PDY2WA6VWu6BAmKEo0z/deCejRWbc2U34dkshCsy
0TUeQPKOZL1ZEwgDdxVsUmBbWkfoyzJi9N40goGN7VE2DCVJvbptQMCtLantPt8sjM6lCMIZ28go
JXPjD90UfNnGOp0mfeeRN1IUACOG9pYfJfBJgRNy/RJMFSXWQBXZg7B/sSEmp/i7/a2Rge/KUcIT
YX9Ai3za+Zd/6bcKc71Dn99ojTguGd3CJG+ghTNqEvqjNcgGr9wwCJzPQhMP18eRKxE/1La9angZ
T4Bbol6eKYBGtFaChfuvydNBrZhcMMyvvIyZ4BkA0/karVgRIdNsEGgD9wHybW60PXeH48mR7hUl
q0/vRLYJ3z2qwo4hD1GsasDkrydimX0srBQt2PjiypFzxWBY/rpKa8gSEKuxEfrvauAt0HDlNWkK
Us0GHGdQ+MJLKRu3ygEMLUunrMkORng2K3pTUO5jYqa/GSyYuJm/xlseNRAiD9narYumXy/u91r8
F0k4+mOliB6Wxs+5/JUfDsbxXPFPIlmvwmVTEEDHkKDbOEeVfB7aqtFcVO5lcwFCjxbZybrYhSMC
+QZMnk9dM0tcdijc+i8adhvYFbdlU922S6swjBjUGwYIYmGADSfZ2WASssGkxtIW5kRTgH5OsEnG
J/ltfBq/RV3e0JlhWww5d7hcCvM2YEO2ewtl2eJ/BujKcZKAlHeKMbdNLHKsd+UwxQQ/8tKPMHlY
H2NSyGcIxTnod36YVN4Tfy32WGyZb7e4EPl7svnfHDQWBqPOqs8ssBH1MuIJtWP25kDMF4I0ZuAd
nR3hOwp5Ic/BaOPM+rXjO+hTY/MdV053g9UXbr1RB+7tI6iyIneTunK7f2QKey+043grhaSdJ4oI
mXCscQjK8jam559BgaQ7nMBmJpmfE20ryk4NMu/NssnLOwRQ85yszvJqSwvTYMe3gmzYvIu71liA
o1OEZzAOdu4auz0n+9cuXq5/g+07hjIrTAg4BKPjKkEe/2JbtcrqOxEoi1hAn2TCGkYOiKZiRU5Q
OGYjnXMfiX7XjlxN9k1gPodU+ccWFFfXylE/vVoDkWnlok8OsKIyvHkdLOyCUlDljx7/GibHuwrB
DPkEvQxKYroWTqKC97lAOTTA1t35ok3V2PoaKi0+arzACPndggx5eqlyivFLS1dLd47qdnKzXBX0
1MkazpFZSPeUg8uGbg35Ac4AB2xbuSP0nxTJNB39tfJ48Hr7HCmLwQdrQF+zOgPw6Varjpt/3QMk
lgjWZhhCs2Tt++o01du0fmN720z7VD6jJiVSF5j7xKheBB8A4J616MKMijnMwNvYTPI2TdgOOzhs
Gt+cdEYrmnmqSWsdS5iMll796o8XfOu+84aPipBzbyYOBjx00DCbA6XNU8E6N6HhY1KX3CAa9ZY/
SXHyZx/5qobUPqJZrEvziFYF0S+YOKxikFSCMzq3A6wX8AqiCEmauY/2oY8JiMJvlANr1BIiVO4S
UCfzfXFCgDEJY7qSs4SrA2nz80QUofZAMTVgfjPs1Je8Z3+wt9S3I+BCK+E1aB88NXVaI/hRBM2K
hBg8IGpQJY9PWNuSCpa0HX+KQ+f1vHakp2wyL9b8V8D3HwDuXW8VxQ1G2UH+ELHkRcH7qo/vaLq1
xQAqWz2e13xE6DEx+U/t493R8ksllB9xX7hKTp6R+fNC1dU5FqoxX/bBi9qHxtKb26t98H3+3hJv
KsEfZddepUkFA4AIzUU0522TV8O5md6Lob5tSrso9uO3vNcjcGbAOic+lJSj//qAt9odvr3f4QBA
5xzgxn6Fg8tmEAk4oYvDGnaaz2cxfXUHFZJB2YBmgglLLKmb3B2zaN8iafSiimM2E9pZ9hXeL0M+
SP2b140ISKANY/S5kOSkRvgtgDD23LJVw9+9M3fjhy/yLbBqZqWhA3jxKDfkMskhmhvPwvLtOv8D
zedqqj98lWesfHcQNtMOJdHnP0QGufJ1ejBA4hSMMvQmLJekmiSQSKiydiYK7H8HYBwTfz7naNws
cxUVZDg+DCKPqCcyx5avrGSrb+HzXA8iBC6r2FFZgiqtuPw0O2TCBxMA4mVFWn0YHCvRhuY4MxQg
4fJLnEInSvSoVa2SrM0RyrL4RCNqJxmadrOvgftmuLHFfuwmzWVm5D61W/xUbSK/w4I561WFzDv8
YhDswsPhlMoNJQ2ZKE95S5y72VJQd1YDXvVzz5i6IKX6bupSddYTTptOfYkGeZ4rV8K8GCQGQb83
k5R+sEhsDRpgrZ2OyaJbjcCHo9EUqY1/gF+K5esSXgvLt6SgMBMuC6SFmBMC1d1btIJUtu1EQmqo
iiSkwWav6Fkybcxy8iJoqAnLkWlfT7y6tq9VeJZYuecNnwAUW+5knms6ydnaFP8VD1BWLfQ0fPBx
/MLP+k7/5AgxnkatECWcUK98humvnUhgRMHvodMmy24ibQrf4Bw44GMAIpq0MfVlEFUGKkq+f18c
nRDJ46zZdoJXErx4+vvwpFXH36n+50lOu0LJC7CVIplg1QptifrHf0UjFtyBlFrCR0B3k61m91RW
o+5G/kEayszS4/kN1n0LujTrwUWMZM0EQZD2a7JuNm7JOYl4alX/mqWMOtGBraxIIpRo6bleDFIr
FSy4PgmaY/mgHYMavjT5IQk6ESBncsqGVf19VOrXstnc5zbqL+oWg78uMmi2K/1WY6IEkg36m1Xs
o8mAaGxR7ISRTmWsAlN6sQEXorB2Nn+gld+rPlwG0osHEmfGGMLiToaKQgPzuOII3MRUdSODbmky
izX7OBd8IVeIElxT4Qv5VbF5ypnadvMSU8GuUpjghNALeKvVBpbRfv1r7A8MJyr1WDhkEHp8fRMl
dHWIyGMYo2wds3AomGqPRbAFrWAXV72Gc9wAyhnKlkJ/NiPEYokXIyxzePP0JUli0WCQle8Lt0nw
gOV6ra2r7U1v9bHlH/vPTcG+ctMuRR6VVUTOXT8PhzQ6LMEPUDFSgSrU6fhkMGVson4bLUZ6pZVe
y5NL5OA46UnszA7gLw3pwAISdW7fDRWC/BHMONUrUN8ygbPKvBbniaotXIcN76h9JTL0TtzwA90I
3oDaBBr4p49eX+k327g++2OfnDzd9SyxSGLlhyHXcigd+PBz73KfYufPjoMqjGXofyU5+J5DQS/h
N3ZX+NF/mmnty8TLJJOx/blodu8crjRIbgj+44qEaEYBOR+V5f40RQB5aHrqsn698/fzhYRcorCK
/1HeIMZN9q3T+BP5baxmmc1RrY/do1sMEXCYe1OdZrsPT1iI3JzI4g+SJLK/k2/rQge1WwbM1Gch
PoefGM+E2MPHV40TCXN56l9tKT+VaXV8KU7VvR7c1p+P8kD+An5Wv29JgB1abWecpTrs5vKDvvpD
gJSsm7VhbYm3xzsvdC92MO0iGq4rJrWR+gxd9Pjaxvogs/M4ku1bBrpw2z0rWrerHtqzPmrvaGcp
vtnXbgIZ6j2YX+cfCL/3yRS74BstO6tl9n45ht844XsXQJVd/RiS8B0myvzkCLD/q/8/8DMaTqDK
EJsnb1N/Lzp5Gmo6inN8gpbjpuTmqMl6rkPXpBy27ZvW1NdV50gjp/pMHEaagCvqyft63eMzTEsx
NkDTunzO36LJFuVwyc2EdR7lGLT2vbwYYoeuK37t9Zbho9JBRMd8bI0+mauZ5XWaVoCyfnKNDZDW
nVGWx2D9fwd7qzMUMt5Vun2nAzdA3RA30oBKtIC7iYDijCuTyGxFG1JXlvIJXSgR5MtLdmV601xP
faBt7i/g07+1TlY8lNYpyHuRHbvvbMBmCjXfSejQFWs0kXPP64Gh4ixUwShEGNyu1Mf8rBQ0KiN+
QXD4fiOKfkh+olmNFHPkQX+aOVkLRhFhceS2zxd+ePeIRDiYTidsB7l+fllHx39lrihiyiOe8NuJ
oz7VEjJNXlqrd/ezooUQy6tPmMLhk/60G/7GfMZUtcGPS8cBAFemOrgXCuPbZ79+BJjEXAd52FXX
745up5Khd5CJmAOgMy7N2JcrqVIUgtVQHoKPvzHLopbzfGsxyQjjqNXkXZdbmu/ozrM6LPJaPo4d
z1RIpnFrB8motJDBbnCFq2D0ldFvcVqLXwc1Rak6hs2aMOub/K80ncdlrqP7FTrnazNzZOI+K5cA
EUmj/cCbFnACJ9zkAJEhtnvxuK9OaWR/6WATuzbmqMLmgSDZIsBJUpN2tLQH5V2QhAI5/MTNJnFN
sJGerSqNcW+mfibjxSA2eaFv9LFs94Sh1st7/cZasjkjeg52rPeRElXifKtF9NdlZrDhtgd+cRRv
nwmI0yhiq/h3DDDyVU6gvGoe+njVZ1EokNg9JUVq6xIG/bc4jekzkXFgpPn932iuYlpn0zS/Oxgh
KIF9pXXTBpS6YANBT3gd5AIdZQCUvtISZMRxGVD+38kXB0GLkSZTSOI+GAokDKOScxNbbqKrHUOV
nOJ0zOL41snwaX8uei3cHgkUkLW3SmERKMX1CbxmdoxSRmiju3TQ2hZuwEayyqIdCSu++TnLQnBv
b369R6WavfEeU86whZ4+Nx8KFIb1bt4Pm58yCdrmh8AGSTpyIfffWHcFvV3yO+w3hPy32ckmjnwi
eKKJVze9cW4lhQwHUw6jyEytsc3VdU5OUeFUQQlUF3GB+ZpxY1lpCbKHe14832esDWeP1xBtVA8h
ggyZ1tmF6VtSFkCMV7Wdkd/RdGpW2pzk4+i83VEy/pp1d0CBcJt2ARp+E+YHisTFavo6Sscl1JSs
yZTVoleSJcBufq0+yqOO0J4IEccfiYb3JrbA0fBDaJn4OjBZLkJ3KStIoC4A1750JugZapq+RqKj
OADJT1i9YUkU0c8MDzV3wYTpeyb3sIBj8Es84mB/2/vwIhBV6pc7daULCBYMRUzm5Tc4DkGbRp6w
YAXo/D4zyluuziL9w4zQWe/TMcphK89nAeM/BVjoq8HGuy/hJ0Q7DP+eHLUD3mgyGOGn3FperzoV
QxbAUXocqfCGty8P6ASgJzuo5KUZqOFibIVoroIOzLJvAmcOZcGhqaNJNkzDk0/K3F6U6hEXXWD0
5KrJYpkihaLVb6mDXg47L9S5UpvfflQ+j/9UmUl1PMpByncpkgGL+2+b5Co10JlvVksw8BhSUqgc
8cHfSEQYOrcImYe+obDjkTG8hDhSYqx8UvUxEvSys71RZtMja4Jl46R0uYx0f5hxIpd4djiR8BrN
+fc8SqCaS6Isf+UeXVT0JGa+MX+jbONoEcII7xiNjmKgcv/c2TuVNhJNXyyfoxWrVDDPmuXYq5Zx
4qGJjUovzSAB/pFG6tfpzZsi4SvdMuZfpPYby4MWjEZHLlDkt5lN/LVgpKbUVTe0i8IiYGNnr9Gy
xL0T/XC0RhEDd8t/CxP9hfty3tEqj9eochdiiub3ez++darZXgxaeGG9BZ9M4N5NFdxhKko6iUJE
D7lx84LAn4QGDjvSQlfV/yhTsK6+QiQ0dBwZ/9fQ7mKF3mQgN3EqhRxsGGZPaR2NQ6XQit7kp9NU
A5GIgij0Jf4ck/7UGBZyUApBLAkVSpWPjvkab+YLRVmJZ4o4RZligrDQoJpo4ocPJryF1rmhjALC
GAgXpvRz+y4pL2LAeeNfbj5WR7MmCSs6ufQyex5maSl+oMAaakfSTtmSSuiQ6sT1Km7tgo5SEUCa
HVIhIfNnRipogCpxbxU6jzVfOQyz+cmjirNizW3d6P2YGa80YVM3Bgw51Uia//8rJRoxI3RvjCgi
GP9DPB3UJTzOJBdp2k1fXEZ757i9W9IgP5z4of0ubeUQOq2fP/jEp/bVHJUmIQXYlbsyELU5n7oL
Wi1M6Y3h9u13Led6axfrWSsfr0q7OvBgtmtEp7Iw6ddfKX8s8bsycWjwe3JGfdEzZQh4XSIrBJRA
/1neNA5tN/hcaZvwublXP9Z0dBZv6lQiIyfKcq8uO1Zlx2Rkt2Et7cImM4NgWgHL0EhJ2cRpTTXx
uVeYdOOvfgjBqNBJZIcKh0ozAhwGwu3mK4GURzAYOzNrOSz+S5Uub1PritAdsdsDeTGb6WA03uK1
hjdCjnI5CrRaRg9gAr802MTwl837f1TQZeakb9R0/NowDRBEcAmsp4fIZc7V+Ov/TCshW9FIdhpH
asFXmoRmtBO16Wk7NAVr8J2k0nN1UMoxwPKAwOqso9Y9VIXqZivcppQ+zHxfxXNRa5JDM9Nv/qDV
EqX/NXFIwPyVLtebGzyy+rTi2C4DYzbPNe1E66cDEsnCyfq/uLcVOLSQB8P7d9x5hjwz2RjUnCwU
uKia68rju2x/VMj1VBt1z7AfG147PkF9NiJP9URk6dUwS+ZOTEIcJddf5TfSUX8OWFzp5hJIZpjt
wprMXJrRQA2zXVl+vQhg4SB+5JwnoWsVWt76WxZIyTWqnViuczEaQK4Y9hnOIHFSizv15ByThK6b
WLkmyCABOrlDL0qfRTjJnhDkVqOfCoxNegS1nRPfHlt2nnKIKdYxSQqaQMuj8k2jDXyBsm5NWQhc
7Y5FROPNzEcyXVEG4agqp99LuVShtLvcrXax+ufL2I/VKlGdO1BSBReH/6ZJM0ZAGIDUen0nMXTa
Sb+HYCxqcA4pSqTmBdFTOVR1po8J19Qh+iQttJNwRFcO0ecbo14lM0krZiGVlAlIkGYqwAdxg+vZ
/2J1YHy4vcETRzW9t5GCOfmDQcmwgb0RZS6LTaU+bySWsbC2zOeoruyzQCpmypfrVPNmnq0wgRG2
YqRdI3+5Ojh0jWgRVkww7UwBBciV0/ebcvndccVDE02YjLrdyLEsxef58V+6Q9Y40hG8oGRE8y6p
lZTlyY0wH7GUDnswrLEB1VnD7y5GNUBQKy56ThEi8RyTyQ6pwLSvbfdv8H9ltq1nQQOClIPqyu9p
7tZBnyJC9+QB2v0EhUUzsYpWNpuphAb4mNJiWq4xZEsAcRpSnJVTq4RKdPeU9L5pQZGqscWOzWyy
lulVRfLNb2C0zknYB8UiAuVEOiTeII7Eutl3tesy/XisOFrsEl4YueI8R7EZwsG6b7wgTTntQCcM
qmfWEyAFvi7nzPuZff7UMQjFrQUE1GPpVrim9xbrvBNzg8qPLyoYz+flTXHCdIvYGQMv8uYPYhks
SOcQf7x8mp/W/dzFC+nwg+eN1vfhxsPN+cdieycleWMHXSZPJAn8uaVHCG54kXzKcRzMmFzSsNkS
P4VLkhQ3kUVsN0I1Uu68/p/qCM8JLUwkw+R+PtKDgBqy7sVCkeyrwpN/BK7tgLyLJNL178G+TGB1
OIP77XwO4k7IVMK8xt0icu5URpNiVq5pmx9Ld1g6iyBs2wmMTKjvO4+IOQOig60jfKD8t8jI7KxK
Uk5hDg3shbfkyyO27OfNO+eDI3Nqzt98Cux6+k9h03zOveU/pxvQNQi5IG9vRTriYcofUvg/m1DV
w5naoFQKX/kczBIvauqZhrUVmQQZ4MOqXh7ZsYJdU6FbGzkwISqDkkzlBW2qCuiR8IyDaiw1/HEH
6RjCwGln7LdY+cS4dfQipp9r3jXjjdpim8o0ujq5ABs2+HBIeBq1Df/k3lYPsKKLSFpqoozOnf5Q
FuxeLuKiaFl+wgec50QHepbzj1qUBHWvmh5IXPALeIJw20//lPiJIshyCfT7rK36SiwFRnGONz+c
68Hv7XnMls0AVtm1OmTCpmpizXIFzAv0t3uJUP4w5dP0XtLhmeCb1v5vkcrut9ZlS0nskkRMLGe0
jWVHZC9AFIyu8pk40FZ4kNtDukXw5s88Flo3C5xBvKGvyMUIAu7/NK+tknfSAnYRoAM/ROJY9d8L
9iD+M/sDzQXd6/N9T4MEr4KuS0UqB9xdbgb73KMTiZoVuktbdRZdX3rkI1qNpxVk1bqTN3E8RTzE
A8oRPrbMNwqr2mofGyh7jEfUHGI3JBDiFmYonPjJdqMMViM9Q8K5qHasrfP1zPNG2tUi4zcyBRxe
a8Do4QBThuKxqirvni4KLaABUfAO4EJ7F+ileevQdEy6kcVOcwOkSgnB34Km93gD4h/r+AUBGeBt
4ZPAdqed9f6p3jb67hgXMFwtPb/xof7pDBo+/mZEYnGkdpuybCtUZqAbgWzGa3NDwdtMRqPTxV4H
YGWaCNzQIesOsU43tbEiHadCoKsmMHbea9y85aH79YwrrjUeIzaTX47DKAtnosgZR1+6C3JpIQdI
3/gXllGRg4BoEj2Ss0xGT/fCG+gX5i9fKuoUgs2Na03XP78vlQR7PbsuAaIhjV27Y/d6nguQsSAj
rwqhry8JDCWrFFlgWivzxVUlDjMrl3I54KuL+F+JwRb9gwg3sIYZciZBDTyhRLfV8FUxad/83fBF
15MLgQ4pfHHr8CnBKfr8GfymidHkP2YD8wAj1oXsYTo+rDa7d8s9dG16vTSmxZwdSWf37dUNniI4
tyKQi++NkmQpSp9AIfP7Drqbo3SJk1lza3RSsssZbtxtq1xXbbW2Sqkf5tp2yIN6FLaRn8GIV8k4
nXkOvHW7i9AruhGVpv0tkA3HjxidUfbTRJsEIISQgcsZXGt7zdByD8bT8k6IdmE/v3FFe3n261To
Phg3RdVxc0GFHgvBk2I5VbLt5OZd5JB4HaFVerReWjoUdkCafg8p5EzGel9VhBZhE8a6aZX4fmwS
aNwtCiOB1nhKf3YoQuXR4LKmL0QTw6Ia3tPKiglvZZChrhzxPtbf6nYkJsCAlY8PRTI9Z3gd70TX
VfNQmbmst1JYa9v8A5e65KncyBJP2VcMDtgmFx74lCP5PWF8soSDiwMWBu9GwVRnfCgI6m2vTxvK
247jAoESilZD9l4VB7s2o6z8ysbjJGQg+y+rH/3TtkB9ZxCDa0H6FgXoyt0pI4UfAEKORr8T6p1j
2d0qXcdZt90hOIqBnwIK3W0yYxXS7xS/8mpEc9h13ji8WZEmv83y7dEmHV8wIF3pMGB9graC5EpO
ItEVw4L5d80Ay+VPfGup3zzLZcMq7ko0LJOD3XPbOB4BndYL+Z+88fVap+8XiJLQFgm4xUYbfgwH
iyzrB0ZTrDkjN5JPr6aiBPeCWFZu5Kdm2RQRqfpPu0Y0WAjsj5KltXJfA4a+v89W9We6zUhoMJ0a
Ty1cxakm+v54BJbCTfj0nzyNdC9ZCDNpNxCZbjP+07xgPGNw1N4vCLSevMRgTi6ZJKlLcm4aJwvW
Jy4PkdpxrJDYTBtiY1Kv4wCy/CJyz/3chzvtTWb4+GhVrEjZrfGITke9S3ELw3JyYK+J/b3Nfzeo
Eaa3rcXuqBXgTMQ3GotGtKMjh1heiUwDIBgV0q2LISB3h+qsND9yXZT7GHaHgL/9yF1g8V3eEyB+
l5tPqFmLUgnLXpY4L8Crjb97SDICGxKFguDDC13v4e5tqjY2o6zGqox3KECRpH5r4JGi5Otyf5mB
qJMmHwcV3fD2AAR/tmLcGsCkghfN5/pER3yqvAxBHtY352rFZaHYUKRh+V8IryLFRN2fGaA8Ivjs
+iwjxrJzcBuyLMGI+ft+sc/ZO1c2nC8qTcE7gMTAoPhY0X1g2Q1ZAcX3rhKIoD/c3dXSsXSa21vj
hh/mdihuSP9Xx+VCm+NwcZvwqRahUItgs5hFywaWpj7yPpwa0yV2wlpg2bfRiM4aY2W0mfsfR263
5WJ+hLyWS3O05YoRhW61LnEubIXWauWyVRzqO7VxxlDSvrJIXxakfQ5uwY8Q1YtI7Sch6Wt8+y/q
+nKsXKDcLrX3ekks+DuR6dpQu2el8bAq08TKGHtMR2+tGpCt8MchWnIEg2J4Tl0aqe0ilm5KG87N
4u/f+OuRMq4G3KawC+gsZcKgPqYwHnJH5rVBUqp+YAqaetsGhr6hOJGl+JF8+FiElNXjIU096KAm
nWacCiAODT3FLHc2efLwSbbyNKnnR7zkt0kYGcOrfmrWoASKWlXm1CdjBwHBT+xMPmHjdE9GbeAz
rk9wg46m1BB+9bfAhT1lWCmiiw50tHRN6tocmItCA9PoiSRK2c9AUthg7+UPpumdbd6QCbUECID5
3xNLRMDUs4cubWjqanym9dbr9PObUgwiJRWJHsbA7kFTeGn6sNLvLaOIMWWxBHIHBXWLm89Vgefd
ml2hpfRFAzEZg+M/6i3/ASdrN4WcMvfWMRqt3Z9ZJCIbC4X3GSWIP2i33udpiA3wyVujMGqxIZgH
R1TraMLY4Zg4xEmzgrdKZtbVVofMiSZhr2n1x3VwijJfds5FvlLmGfWv+5pFeObBSN52ycingiBs
TOw2gPZrijniGco6wkdTDiiyajDnwd4K2n6ekRlnWxTSbTYY+ihxontua7Hb/AYMa59XL50Nw9u9
p901VXJ8TbUzBejYRANApgwItIGErCTtaF7YWV7S7dsXDAqBdmxM6UZe5biPlhaJKjxsWveCwbUr
LyIw3CniL/KpiQFi8OF3HKcYxzl3Mshy5k0vtWVNxFdKfDbPU8Ajt3bPztWJF/kdR9XOj+gIPZry
+smQJDK+M3sBDsvZM/NYX5QR73B2Ev2TPYUIW/SihUK5eR2RTzZZ3cFV4E+u7J52knE+etr2W9WN
OgsAp+M5orfStiQrDODwZ0y3pTiRFNkLicoPbPByjFpxwnaTqQzVAWUwTzFq1nN4eAkmQQiVv0IW
/Dr7KCKeNNGJKieWa/P6ehrEy3S0gKlCtqq5zmRZsmZ9sGyLIrSI1DsiLt2jV6GjCKiTLmUqlzjp
v3JbPRjWhVBn3UKff8wFRPgapcOEqwxZgo72cts1xsCTEbl8B01slD3DSlb4DHJE4xZHUcBv+ev9
VRAuHaY6vCoeZvkPxW8sRkpNF+SQRgmy8qx8ZEM54PjAVyz+87rOgnI8TlqJjM9ycKrXV2+VX75z
hXh3YChhlFlfV7Vk6BTvEubT+i6cQ0xw4EdHqVCZJPkQBASZwXjC+VaZQ2hdbHRHxAf2MB49nrG3
dd2iyVAj9Q77H4NJyWcPwHSIBOLUjFSyAKuTXL0hbQIJhytgAeFTyxV185vzvMFyyoWyIVdHQgSG
7H0focxrHZF+sG7Snv5XagjNlRQLyLfRZJkHFv0cTkN+1+Ot/eL0plp4CCpeMX+Nj9UX1mW8KiCB
E8t+fOD/xXU+ut6wf/b2yTNY+/ZnqOLuhZ32LdZLveZU+qYYbHdDNQdxLbeOQB4UyqwHfBThIByu
3lYgD6JQvAxoJFcHBxQyzpvdEdpvnrTyZn0B2Hs2PHdurehs7tS/JkQqd5TQLbWlABRYq0/3XtKb
vFED1IEZqS9NPaEIJ0B7dWG4OCiGcP1nrvezjOKUEXgt7Y7z6KSvGX9HCDI1CAcdH/mb7nsRvQU4
tGrdDvE+wYdAVTfSkAlcjjcw49zZta3b+5cQ+HMs1/1RyPpvNvPTTfCBj45LU/g6uYx4g+19MhY+
LxSAnoLAp+7R5FXhn3m+h1qoqSWZ9V3KXlcyU9iq2jtzGl3Z5zfZnD4iRY9ADPVJmg5Iwtlg5p7E
sutcA4CS4sfRmGFSPNve7YMpeDv8dHB8YxEFYE5ua3cYxtWM4w1+M62bglkeShyETgLEh9nk09HT
+Hqf0t180b+OAZTy0Es3tSQXoA5eSJP+FZoEhQPEFw1csMqegY13NpL49MLtBkm7HO6ht0TWUXWs
+H1UQ7U0GgovCCO013K5LF0HKNJ2YNr1ev7wpJyjsKSpDs2AsReI3kWBf7f6ZI/43mRclruGjn07
jtkTzHQ5TZBmfRUYp0PLpVMwt++dsn8z0K4PT0BYhKwTicGJVbrpZwHYSr6b8rtjNfuTYy+Tam87
7430T04irlBj9G8J2tOh/Xpm8pWgHsCD8wktwvrrNXzvBNIyexROP+2gWNgt2Ih2rik9YwxBpQig
Iuzmxxifyy3pze99Ltd8EBe1t2TLNzTgczo0FZ7ZicxWFjHjhTNXiOBIdM2zkC8NQagd3uqpNS6m
sYKVOWYwBUzryBl/CnaKcOgOXkTVtd2eTCEkRclraIjm9tik8OI/0Yvwo6oh+lDSYOuSoQwVQ/A8
msaTH44hybZoa0oXdtl8S/4Y8oh71UPno/xHCjKWfsYDDRs/dCu5odOKq6025Nj1yyvRTT7Z+8nk
I44AFfZnrkXdgs1YrKKq6x36QiM1P9JULqa+Efg8LdO9R1HP2Wm0p+CiHNuCbz0HDCZZlHCmQhVn
ofbC7Q8E2tT686vjitOrdEBovG/nOb6/fQsFxzoqrahHWfbBMNXuouF/0cVyiw82TnosAcZUv9lO
xQp+BgBQaenDXnwAVlPlXJIX2yA5CO7bCXV4Xqrz6pqReW/cSKOyKsqVlQGkxDyNAN+BOaRx7JdH
DLLOUHmrJshp8Hb71dpaF27tbO6ZsmaSlh8xt6uE0D7SOjq2v4Dry46JfBANAiGLf7wXyudx4B47
BGmTg4dDHh1xsakLj/rkBaUAZsRqBuSohiOzovxhWTmZ+rGnZZcFI8XAXtzdKFIH9roOtHHTvS4u
uQCqdHplfDwS5y8mi0I60ojLV/QyWqjjNFuhmQdlYi8GAwU486diMBWtvm7WysF6mxlVeTFcAuAS
Reqh+rUkv4KpiA9RWCyOKnzqnV/72F6mrvRnrzfdAePRTjuNioRZeC+iKQUnmXm4CxqahLXi7Y9Z
pGU56j+qL9OnOXR8XzBRUjrzvlLIzr7pII4H5xP5ehqyl0qfz6R+IawF3R0ZsCZFTSjQgFiiWuXC
9g5S48GDg0RqJfcP7N6fJRff3RdYFH6UnTR8t3iXStx//8x7fBsUgPcal3z77w1bH3+79eRTROql
cTvPp1vc9fu+bIFClfrhxIDiaZ0/UNZtI4njO+IIALA4e11FjfSl0mPxDgGK1ASUmUCUkHIcKP9p
zrqQa36prgEBuZ4jZK2VeAyKGokrw43JtBz2PcX5uQ0ELeD7LCsWEpNCwU2+uz1TrqhdT1JWvvkr
Xs9I4swjTPbzNUtb4BECPfoesCljoTWJr+Z+s4/U2Hm0tTirl0p1Iu/VaXLuyjiiYXAwxd6T+Zbt
Sua+WQH40rtJ84QfvN+VBsvG7ygv8b1qoWU02BwA1hHcRWltD2CMtUZvX07j3/nLNM4f7Qru6lON
L1cjV8gnrkn8nJs8C9I+FbLEGQHK/IKqGs8/m5xgLOzJPkVKhagmh3/7VbVibK09kXHpQvqkCUOB
fAXQM7pDY2PzfAJhFh+TgPn36dCsNzmw2rOCsG8nGYGPsLpy2bsn4vZG6yUaOKr8/ViM+/3W+yAu
seMsp2axmt8a/yNmzOtveSwWT/i7XOgtOVqHuU2eXGsc/5KxYADNkf4ojACvF2zFEGP1ocUnYeBm
ov4fjBCe3j7DQT2n1rSEZVRmlNO8GMkcKl/bE/5GYSJI5QFPAP/XnOjFJrEWf2xzTTaI5lCvPQDi
Wqt5LazgDHbdcRhr+GeIN10Q9uWhS2Ug4wy01fxos7m3NjRz9LgcnL+ZLw824DMTwoeORUDOZrKk
tJe/QXYIdnF7xzS5EktYP1CGBhGzZswa41bbJaAskOk+JsCppMTkQTOqrkOpPWzgYnKTEuxnqndq
YS70TUdQM2WpTIXEgxrI24hIoCeHEGMrSaNf4f+pvIb6duIFpgYox/T++Ka9X/HFRzrm4bPmuVvz
ajvG5aj2rJ5uBg51fhK6cnLBt4fTJQuLWZwP3pw+KD5VQJXEsHAn5XXIS5oz0kpCKsbDrZ9NnvpR
IFl0eTQBV/eVmwWwVjsQM2iGtyI82fPJNfJ1tuIpTj2pfesLkRchznZmnGRu8XD0zI2c2hl28Qpx
0WzDyvGA/qcmICZcqVxbHPt+7MjpDCBiwBPOTwNE+Rf6k4firS+Zqwg8uIe43SIkiWh24RN+tqq8
aUisqKs1S34yp7Grs5E0D78/eEE6okj7hT2sWZFNabOCrtXIDOG+HkWRwmCTKsK5wWSw376v0mFN
oEO0HQzSYum25H6kIt3AGwUJoUR4xXRuEjUMd/niYxRDt1lh0adzwcN3kIOlVRwPeAEYRjrZuAxq
qcm/f6oVjtjbusLlsAX0wlXrFBhsURk2qVAO8b10GuBoFDr3ghgxLan9/Ja+LWE3SZzIFY3V20dl
e8rKKJG2MXsm0AwdHpvOGO9zoFI56cbIr9JDinMPG5U3j4HFYYbdQT+HPCSSyXV5ZF+cVkQ7vbiJ
c1Fyjk1YGUlPlhNrFa7M9yw1e8y5hxIfJ5I9TXjgy1iPKSVa3XliQdAbJMHDSxqb8hGUAdqs6V8S
KXbVJhFgQMAywXJeqhBZb4nVgjaqOonl2BBS6exL7d1TbIZ/oyUUOcEJLOvCKfmgqoPWu3W8irMB
dPqDa4zfsnWWHK/CUm0s9uH6Ru3vYv/X/aiZjY+w2QYfgXqNFLFoyfCqPIN3Mp2C4BDYglyuBjOl
TW2Tqx2G6OO6LkGblpDgDtXmcQX1Joq+ZmGVQucjqclHpO+dBpraqE/NZmQvVluhcCjHtBI5nvK+
BU70CbiwVp3Llav7Ro1WDLiCy3Fwt0Dv5ZL/W79v8gv4l58H23Gei61bWdYHMo6PSY5wdylUBV2a
2DmCZxfiZNv93htkMQHAQYeuxT16hj8T+M8ijwl92VbsLZAAHoJr7xzVe47q3PWjUND9nkXiGIBZ
uRiPHYryIw3V8mEfwswZnxA+/RFQ5C/o2S7prXViAfPpEzjSiwXk54wFkww5KL96DJchwYtzSZZn
Sd7b1DTj9owO1v3mRtvxAugNwcDtQI069q9t4XrCsL26fGDKBM38JVGdqJ9qw+JpXtDGtATcuXVw
iGylwghz+YF8aSjrhlmwdPW5U03077tmF6tSHfMKnRbzeYIF5nRNrU31gB43Miw3iq2ne0TFg4US
dVfoTZwdgNJqVgSRrt1xjVzxhxQ6QBM/Dx2/PVP1nzIwFntd4ePWZU0BFeKWT+8j1tOwkhahXyUC
dGEAEto3nCE68E6xhCuUit5nHg6qh7CApnBnjCWf59UYg/MQ5YY3n0fqiT3aRQrCtJcvXsw41ron
k3tLP7OtO/xBM7gNwliKHzt2g0q29WsRc/EB65WKLQdKuSz+NIHQ6pcp9j8Iy0vzuozNBHR11sgq
57gc4b38a0uYjXUcPYLFPzgKvlf0I+LD0bB/ztf9mTl0rJWYc5wREV1DJxAhEmNlaY8+2PkAtxaB
G/CEeYk+ultwyU3ppHirMDe+l6gmEbbnI5jVeqdsl+lv2q7nCA3jc3uSZArCnlGPM9FjDfJiu+nl
TSk9n7/sVtDMFUTh1VU0uUF/NV8QhbxETBBCqY0XsyTMuABmB651AfYFTkEA9XoXmw3mO2ANWgWh
fY69060QCHjeGJM7iDKti1GyqbuXIhZ1dhCe/QUJX/klvkMIL9dX2ntPzOVDq/3AGbp735umX9kG
bmEgrNR3GkcQ//XnlPCVcxSXhmf72qxIwhJ1sMUAsLtqoJLb/U4+Yqxb90cZdPA/XyH9YJuN1aQJ
yHrD3U1UJCL9v0+7s0eEG8lAPxAvq3WkZemmF8CEOnMxldI58iynO7zSCTN6QtYfR53PI6FZ6Gyt
8Q8kwK2ZdkL8gfW0eqwV1tEDGbJRWJhiSXH1+AgMFLo93c0lOOK1D8KtxTdJFu4x6ZJ3LAtKkAHH
GzKrkLc9Y5mNOe07eu8L2A1FKBbscoy+hQEoRIKHJykXmL7p+oEsIPswbwdAxQ47e1ZLgEKdsYZc
f1k8WuDs/uYgLdWrPaW5SV/IlDadGz/vupniYNyrQqxaxlnFuQW61R0dZFno9n+I778cBdeCF/J6
cX5hgLRpjJvBEo3k5fo6brgQZaqagcPs5Bx80QFSnx8ncYwtyp24hDMJU+G9Q3Xp/2v7846vyG/d
flBLMujnvI+CnetHyqzzqWkUoktMwFutbzJZ0OBpsqiIRVVxeiwgwmNFvDQhF8dlCRGkeiIkeAL5
j27RBRID933qw2kcLt1KMv7x/Iad6e3lLDYW42hAY1svuKUCAQN2Q5mzcaNj/4A8PGGYZuRZBoHM
sahJN1cCW5YNvnAGOzVyuwTDMmicbj+n5ox2n4Ji6zmOaAL+L5SAakI23ROXX1ODTj3fIhgB7tsk
1fk/B4yHqPird2qyfZsAijzUCAy+1RuevM7wwAkd5x2b2RRlsy0z0ptM2xjb2eumwZ5CylbeYDbD
As2zKCrQHjYDHIWCK5LjKX7jo1xwoOrKOU46iwKjSlIkgp3BfMGcbvmDzbEXZLMJKJo8YG3zFKGN
NOEemrnuLteKoCoALgxdAJOsR3IqDlNemrLqNc6a8J0ExyP2sKMmzEw1aCulfof4i41cCq80tLTG
ORtoalVxnX23e2KmlUiGSO46ZR/Htvr3JI+jeW7YbZkZRBpEgY9GyxihbJYE7HX/mEdB4X6Lq0Ku
ofuPTRxm763AEcaFA94uynHTjznLCgVAGeLm9QaNbEV6E0p8mVplBfEmn6A6DRgp35VT52CeKn4f
ZBC+vCiXytnKh0EDLXd77/RGElQk+A9dBP3tzmN3AekYq1n3LZBkKhx4UbCDrU+m0aylj0Yv2SZK
HUDawXrlk/QrHA/D1rTIsD7rSuCbz9oeo/54QpkrThJlohIvU+5dhr/Y641HsI4TjG458Z5P+2i1
xDgfVdZYYiF5sIlfU931SJytgmlXqCu47mztnNSrPaY558hY1qbDe2J7BHtpWtK0zarDN6n3DFdr
IiX9asnp6uxXAUybb1V1gOAe4tzxv8a/il4kmJhjzPd2PVOc79wHbOP0QzHF7MCEeb+NRGgBjnqe
OcNFl/V5wo/K2+Du8+fPUZxxSx0pKMJg0fXo2czky5aBgBhy90AvbGVDkYuNp3RkOnP3OF2uLet/
FD37RW56lE+nuzzEdLa6ZMu8Sncn5K6PmgCLiZIQhGxhRwEzqAdSTwkSAL0cntuNErwzLYacnM6J
HkHcOjG/fWBVZn6iDXybmxfL+KsVuFbg6vSkDXHF/LWMaGGCb+u+wQQ8LSzqnQayMKFyqaTeVKfM
xNlPSJ+lkWOV9kG1Y6UBdjrU/0XLJ2cxHS8L6tsdSAkl+g9hJwBUXS/k1iZVNbKwCC2giQqq9lCH
WigCDmn82f+mdAdqRuAqp2nQopDJlQxG/4a4sxl0So8AXFFU12ABubZL4rw5XPklcTVkV0HA/OMO
cpdO9Rp7ne8mOdRay54il5N9m5eXt2xHGUEckbhErh0TjK3T1nxqAcV1dsLQF1ufw32xLh71suQ8
vR0sYkXoPRfPY1zb03x1dHFaUnYpVmUKoJtc9CgcgvsGceElKTweMg1ErkXzdNK0Cu6oAbAChRf9
gM56trGxG7Rgy4yPC7tPmbzl+7HHkhHyb0YtECWhZGFuzLIpuRLP0SQOB9Tld5kSgggGlMrW/3Ic
FI3rxHnSUO7lJvbIvlXl7lhLrFSafph6TUpuU7LiHpAn/f57zhSFCeHOonSvovfNl4o7ZxGGTtm7
vnOGjpr3d/TlAnC0q0vBtQiFdxn3yr31MvfEn44EFRkHzUUX1w7rQXrO/lxp0iXp060CqZtigTyk
P0X8YQtoepj1A0/x71nwNTwgXZ9C9q37D7OE45Mk1bod8vIfBWj7/JnanJZVamIpISL8hdbobxUw
+ANSJBQUKiVtUrDNAL4wdUdRkCYAeJrpZ8Bhb1+KuOak716Xuu2OPar0zIBRuv4nVn5VD2zAnrpc
o2ZrYFcerQaZCl+3mJ7ySFysJZYl+8EUkxhDuEnCc3tmLOoM4O+kv+qONmaQxGE7F9lRvV0SQqRb
1qXGzmQdJfdZK+Qh4LurKxUgKSFLku6miQ8HP9CEBamQYUAZHteB707JkktPle51Jt5v9EsjVJmu
WeNfuCI1HlN0ux7cG9dZcegVBxdcQiyyYkjAUS1C4RdxJyR+yTXFqnzOJ1f3bAcMYo8VBV6gaaUX
KivKqb8IfqzhVG/aoJ+AMX6gRmDjMF6iy0FLDnvzTyOSnNcPtr9PBKH9fIzJWUuD8frv3B9SkIE6
wWXI9agVc2Z63oWOVQsQz4juoyyyxqKmyNiApzYmGf2VV/o4cAMl/JcllPCU4P5/cQBakTHc3Mzb
Qpfg2oSRacv6MQKTGXx+NXhUtcHBDS//L8w4LvcbcyYPdQwNKp368zu2HJerZCsLAN7t2FGOj3Av
zosisDzOlmO1LF/UCdbXsM8jTs1uwCxf54QpzCmvVsLfzcUGvl3/hGjAIeU3BAWBZzW3NwUcmXSm
oeNHaHeEcScTxx2MTm2p4wbdRle8wNWhswHj+F/1ctfKqtnBlEOuBQdFEa21KvlvRo4/2P0aPnXB
ts4Ps4flyd7fT8FtetQ4NRxoV3g2HVpKDOgVp+nVDgFfKim7LwDZg6JnLXbX0buzsqRAYTUxRLCf
qQ56BsMv+8c2DRUkU0K48SEmwrxqXT+vFOWyrVdgK2yXufrGhWgelYt+fzO7iYTwmimH5A2d8jyo
a6xwaBd4hlFs/j3ErQ7Gx8mlrg2f5Hs5XFWttAcjyxJQxLqsT2xlenTa9aIxsbuutnJwgo8LU6Nl
dPeic/FgPAJ8o/CLjSN5SFFCt/EQ028ZKu49zFg7NSj+4ts3fMzuLXAFS1pFlpFKcDo9YMbnh7/O
jpHd5PxDbbemkymjcCudm+W2GnN6NfYOUBHJVCjI0pSUZrrPMT9fjebu5Rt4221cILFPrHjUvle4
HfODovblLO9DGIzShchsWXy4TcPRPY3n5jv+m7KCwFFYfMttxBVCy43vacKDS+McaWiKpwbRx0zR
h5+OxwPwKENfjWRL61AAg0kZK/j2V96wtCmQxRolU+V07Xh56EKfuNbkrn7O2HHHuNI/TCjejg/4
Rj8cdJy8HaS4YpXTcUfBrPx1ovRhL38XoDV5e0qHUCOdl8lWC+VWvsgilcAuPc3XcswDOK7fp7SH
CjPGmDvA5TfEpshCNf+dUCQJGiIiQXONK2NkiueJ75hhlEQM9ty3GsaS9fC2XfF/S/8a5rO6bSiL
N1jIcNPhLsSOlHZllnIgATTc2RxuJDz2au9YV/mrtQXF8APqrh1lB40GJRg7M1t/U9uy8sq5J4kP
xEkvAfBhGyXIurtKxaNNDhDkcZ/K5nRvWnmLmqvPBdcEiNvEdkrUO06j3UwxDx1KtX+J4Hf6I4el
5sGP6tBLgtLKS2L+ruNqs3qD4ZjvjqlN5uM4QLWHJ65zpx20NS9tfrvJ2NDCICFlnn77qCNP/5bK
F3cckRAjjygGHBM3SGUnF6nGzuiw94Hx7S4BdAFrGemw+Hj7dSROFYYGFiBPl8xjqqYZ3HLaQKMG
dZkBaIZwt3zELsSHlmCZmINBQHpRE5xTVKIqqjzfHLKTzUe4RSAWZ+W/QnnxDPMcp5FObZ+V86bP
GSNxhoGitkopGPSqAqNn778abQrRz6KVxifa04OReKDxGxDD652R+pqoL/aRxdmWmGCuZ6TbPiyB
SNTAea4X/AOqcC/DMTw6ZA4jvAxBzBZs35y1YCq9UKz3YvPtI88CE+yUQJ5JiJU1rTnDSoKh29HU
NFJCDxmrTJMIuvcP3RSNVcqMtLG2Wcql2VZ+BISwhae+3+7+A1S5fB56zG5tX5sNK5I8fGBeIE4u
vAdGtJJf1UxnO/U5ehpeN8+YV0S0ryVAH132Y2XpEE1JjvGsZZQsGwKVvmU4PHw78sAYChocBn+X
Uxr+am2m/2u9QLhdYJ3Y4l00aD0MdFpx5h3hCqUlCt8w8KpC2mBVIVj2Rq+g9TQLZKI9i2PyKrmT
mXO5amDcsbA45mU0C3LgZVaCDVlvklUwy/ORTy0nmRm4x+bJRZF4+tTmWK/4m/JKzaLEelb+G4Ih
OA/lwJeWPrppJbcmvDxef3gybaJ9hAROQvDg+5K4Dl9rO/VifyWyNACa9qnWDXd9PQF4zikJyiuP
KoFXgrIA1zjHsrBAITmqXq1qfReONnueOWP6g4FYRTQE/zqDx0uznm7KiK5tM9IF1aIJqKBvtia/
K0apHCDqPGjQRoV18lIHsi5M/cg8Q1xgayecJJunWT5Zlmzg40Wp8xaEjWrA4eo2+nhvyJXkko0V
OtvzVYLq2IWH2VdmW74nzGV2T10LhRjNzQ6OOycPO8UeOgJ70u78+wtDtpjeXI46F3efDzaEQ9GJ
SgS3x3HmaSHKWvOTbGqo9/5cIkdUYF5Y3kIp10Uu+SOz18UC4aBAZBTxTHS68B4g59AMNFmAmlxs
+VICqKbNIcelZz32/3YaHlGoXEJiQR65jVA1IOhF5nKI01qweVJcL1+0nYzqZi0jce2LRex27gNE
AJdCTQ8U7tIqGxX8RWZx9DuBANqmZyryI6MEjExFa4ZfFhAIACAU+GoQJKOG+upZhKOh/5z5T8/v
kCkLKHnjbGOQ9Yk4urVSetPrXrMeSt131ZuT1meL4timPdgpmV2yHuS7Rls6U3VACGOQvUwgbWBh
73xQSIRg35whv8jMoqIbZbF+KE2+/ynPDndP8llImkPjRVw9mbX80tZU60eNhqPVNmjPX/4tUi/v
AQ9+ZiJXB/tZSRBNqCe6DDihnNFnS1FtTFYR5NRB2tyzK8JtbE5JiwbXmHW9t9PxBGyTnKxLmR8l
Mg58Q/n/ehkXMrm9pQynH8UL7H8qdT+pKHyhr3DrhcSdVYlZFcmDQjETE+s6g+46l6OgRWYiQLo1
TfDWZebi1GLbJrU0ZCf3Rd0DEzFI+Cn71yOEE2NHGjE4l1Z59unn1r1pW8v3Qr3WzMfFjCQXv2DY
PipswlglRSxD/pgtEiGo6ONauKUUrwoaSuzIfDhEkzx9BW8u330zw3WsWJMBbq7lI6nks0C31Fq4
Y0bQh03/qvHxeMDbtQgCQaloKZfkfggUgLN1RdKJarNLoWhYN7FwwPd7kTsi2hNAvvt1kdb796a5
3d8tQi4MrvnGwvtgLDbEWAcKFe2xOcNCYZkjp4tHf6/JXhWNrW4+dsOfHVl5jCrdzOoifh/pEarl
SqzA8mXt9C3Fnbkdsu/7yjhGeKOfoJHfcbkLVgwap81K9bOmnYNXX+eUHzh2lhgy97cEvDl+YTIX
rM2ViDwwsK2Tw1Itr1uAoBOPNiW/EoEH7EmYqIGCDD8XJYxox37FfSl0kCF6+BXuPu9Ia8t+NGrR
NlphY7CvIzhx/O4WOk6EtSC0B05xz2tAWqM7MYYjWn+Fn6B92f2EBLEcaTpgEIenHP86jg3fyei8
QxyjJN29N4pEAlliQtoNh0TjUAuVh6YbF8moM4gcowjt1QvG/vOGFESl1jhfMhmlc438po8wGniz
AgIvdRptp4b0R3N5ZmDxMWNGWbmwMoS088Lic1ldMbqUHHeLzIFEsfAEo+mIRRSp2H5IK2fxiK38
cdwEvPNkhdz6z+Om2Oi4RT+fBMDE2NvPnHejQJuwwE6mE2oUfYGEvmaRkZNFDS8p6MipUNeCdNX+
Yf/ARA1Xicwg5JIFDEp3aRHzjWdPS7OJL+r/t2UzzZoFA8YpakCz5rXjUcET0q8HJpoJtFwgHwym
uDlfwHWf/+SkysveoA55TTsFLvYmbX0S74K3KbiEyd4Wf3gMPKd0rkDuSEYz2Of1TtYSKljKxEL/
yQc0SJoT/Bww+9uOoGaZ5fNPeZcx0dY297UlZ+aoXw5YbOuH4xbVoCD2g0il3sh61G4Ngb4tU3+8
t98+X34X4W75ZZ8aEqYt0bddrdhHdtOp18a7p7x5Bjto3bb4+JiA5j/AfvkMWWZxmYPP814tZXku
mcW1ur2J6DutCEEAXD3+u5ld40ATSf3MOjUzgeH1DhJyWlGZ/qWeTYPI7X95a0LoVwoH/Z5SD63H
8bUq4jTZT1VFjxhaZEfMd0Wtj6i1ZFY7r5j8hjHb29KoJBPKLbmII1yOoUtdb+5kmA/+9XWo4XUs
E6jt6mC3BRL10T9ZHvru72n2wGpFYLW3p44gvCh8Y6jAKtoMsbj24aeVIK//4rDKDfccsbbxOuf2
DJVjGnAL58wyQjvkPNhv+NgjHeAuUavMEtKUuXxUr3FExruNbyvLH/tbaof7CIyIcSa9r8uWHL14
hE5sGhV4iXJM2Iux4LDqO34Qe/pIARe+//TCEUWWgTrVLoqaBuS6i6ZxQLEgsk1siuSl0afzeJ9y
43IW0cWw3vkYHkdwqJnZ+Q7SVwA+fpywnGNyPpTNAt0lJb9LsPr6triwu5A83E/68AbOXki7RIsO
+bDcsOlAbtv5f5+/OK8YZm16xeBipUNWH478nAGZC0xM4h1PwQPJmcO3+p18XwMuKQpoCBXXbRFB
YRCmbwtXUpcnyWhuAb8YieTmSt0N7J1JL+zWcW2Ph4OmVoMejx1cfN8A28tnTvqsJ7zXD263nzxH
4l+kNv4+eupHo7gfma8deOC7eWZoLk1QEzGy9iQDiqFWj9a2SnEW/OEW7jbli8/Dhm41wikwdoX1
nkAU4jzFV6itdMoPlpoTez9swSbC/LN+dSW6vR79Qud9q9jMZwttBJrFrO+UWS68WBS8rjdXGcu5
DYUNpH8B4AJ3kModwiwJJJ9l4UYeRw3/ZeF0b2h4OqoBJ1GmHsZehOl7w/nswb8QmE4YWF0+vGxx
jmeywUzvzpdkhroYCCN3yppoCGZ16ZV4gjoNCA1qw+RiPKsEK0FDFcxSXv7571JXwN3//OTovDjC
zyf5D7D2sxQiaUqXmHJRVmRJA3M2BQSqeio/WYXeYi31yDZ6ExeUPQi9Dc3VI/YWP3+8sece31f8
oGrZRypjkfSP1hJnRn+OYhilTyxIcXmVHgO7eDmrot5i8kWyONwhg9UTaQ03p61vx/gLiezsNJO0
2dT+eGLBJdjclB5a69I281kdh34PDCTyhf7ePZ5H4sLZqef5vKTQXeLW8riXL6OJjexHd/4w3ZG1
e9VhPsNh+rNVmIPN5OcP5rMzv8Zk2GrSi2jpTF4UFcY9Fesyok7docttcboftVd/abeTBXMSYQts
i5VqURi9ArTPfWv7DRctrXMtiZxbQCGC2GvXcUtlwlmaoF+hCZlJs4F6QkF/nmM1itU1L/eSA5C/
n6jC89FhbvCDf+GwcloVI0YtRiKVi4RL4i8FwmnOv2ctw0Z6ecwg1sb3KmEDBK4rScnv95n38m+T
yulIaAgWr7YC6AHFxvV/6Wpa2a6h/14hx1AmiClh84RJh7qm1RF7qJKv+PKw4hDVdbvaLt53QF+O
qnl6b1jLsNQXvtrtBJdn0NHH16sVwgrxB7iQ9U+XUy96XVBpV6aabFndaIFPN7pExL+LydgsKfNi
uxNCqVn64lEl8qk5qb9ejvUxsmZIA7AOrhpDVqZXy+QlwjrkLWhkN918FGIyie5EX5izKngYlTTr
2YL2iCOrsacae/Bp0xZZDa6pgrGAxcFrZk48LwrXAiUvRJP/iwZFqzl2lt9fv5Z9uNbxRzkQXKmC
hggTdxDoXhB94eztIUWSrxEHnxzS+jPHKBVjx861ZMzNrieehgLi7LSLeohNjuttAMeomuEDDxC9
Tp8HZ2ft7ukA/EBuiIKdVapYgt3PbYcwfnnANvCmlee18sEyuF7obSTp/10z8zdorCuTDhFjdi04
zH3LljFqUD2wt+VlxRJO9GwXQ/NtV9BqL+x8HMw2zyVokeClJVL3BXbXHNjXKMZci+//x5yki5On
gDcX8Fh4JXomxQFVfYF7eLW6kx6460cATsYMuw4JSd9mCgshmZlpRaOh84d66PCzzjEFgthu8koK
oyNXahb0jNjmsFkdcUqPle3LVNIzv4+MawwVJdkkWDLbPxShU48CGFDuD5Q1Fj1TGz94hZCvFBGJ
tdTWFVB+O05lcBME2j1JUPhiqJX2Fb0/E6HuekF6z7SIucIs9MLRqdWjipMnVcz/JuQ/kfDFRxwt
6cxUH07v1qr0++I9XOZGiheb9xVSkFJKdlJ1IrM54FvbXkYWZDfbfN1jcBZqVa7r7DzotlVfXwVs
ormIH8o2oEf/FBrlltGaTNp4HTch/YeDGMiN+YHargbgLr0EzfxJ3NZyfTcOIpv+QCpHhyV6jYsJ
3aDjoCtBJiEDryi3tbHmt9GDwHMMleK3yzw2GnNaA253E9buOyUyp0+6Snyw2WwYqRD+5AnLgBg/
PPnOLC9S/hzJx8Tnl5F23h9h9PQcablioRRbTdARGddLGpxlBWw9UhFPoSf3xWPSsE+U50XWrY2w
wPpfY/Iw46HmCzZz9YkUl7okWRbZgMe8ZpvemtdNeh8dAerlUEg8llo/pNUQadhfSXgEoEZl4L/D
bPF6o+/WuA8wQZNN5pcQHd7n8xI0vNvkZja+R0ubw/Uxce/m9m1U136hdwePoUwEcA4MOBGPPyPx
Dddx5zzgeQxoHSFLk0m1l6lo0popDF8Irblq1uAL2HRpiQo5bE7CFOFmzaitC0zw+D3l8fUXscxQ
6YldaoL62b86huwsOQipKsFOU3TAKhYNVfic4LPWBVxYddMK+ktnY7eFPzpPpAAewgd+dp7//tiI
bKBr0G0pdV4kyjawG3KJIEmFEWGDzVriUoXdWYC0yWXZccftPDK/wQLcSaxnZxPlAwd40v9UYiHP
UE6DGGjzC7fPnjYqk0ZLIdwbEv4haAGVmM+V/+Di1JxAvvl3ZdsB9XJPjNcI3KWEvzU34nY06jw8
q9Xjc5ngOOF3kz3Q7ghj8gG5EZ4AYUfNgEb4O9RQmnpz+IE6OH4siM7scfa+IyUzEy/1YOulHW1R
/hgKN/i9SzF+4U7LeU/HG4R/U4V8NgNA/6ikUnmPEhVdGV4dSfcftwtXOHw4qn8iYk7RUj1JtUyd
i8PkB+zbrD8iFAWrdw2BFjjwa6kOyKPXiR66hTl8HZTQqeVXt83B/4R8wnXo8jrf3YSURdkiSY4j
gqLWM9kRubM06PJd7jVvP6sKspRds6VhOiM0aFx3jK/x26081qrz8Nz7JZe4Op02xcPMMZs0z8wc
66Rxew0RFAiw2eAqfuFL5h/DJazaV3Bu4+KaWQg5iWhtx0J2e7XdvWTLCN0ByX+o4+J/ln6V++tm
Ce+CvCyoi+AIrmpOTKwsATWnc58eTXZVh+O7pIT3jfpiX4Ys3vOQIYTEW4tS67WDwoTWy3Z1MdUK
b1KxvVp8UuNz/TdOmVBOcxex0/ZlvoLSyG5LAljYKOop945sCSxuwPMLnUQktX4+OxnNmgnRyZY1
vAmHUcVHH7TTLkmLkrgmKe2/eMM//v1OogxoN4UPHG5v0wsjZzBlwD83mvWzCUa5gh2ctO1ZZazP
fIJGmeImU7SB0TU78jMIAIckHr2eqzYn/sikgDHVwJPRZw6tvstJrMgJj4kuP/I/yh0lGvWTk0y8
5l+L3sKlL9zrwrfD58PgYn3gZuRV/yg0o4NXWCDSmqMsf0Yz9K6k5Ae8FMEKSorvAc2FDGMVylGr
7MPh8nXAdMXtFRGw8EEzAwmmqCisFgVewgCpUtLd+14mI6pMgLy8PSROo4cCWzwiPQuwYgoV1+/k
s1+xDl4zdB5980dPTIDlF4PTGo2WTxutNI24n/Vcohm7XEiS6p5sMgN4T2XzMekZ8PtswPVxgKRt
y47NMdC68k1CUsnMIasGmfQvLHtkdGZRQpeiA2mv86z+vaNwfxG6uuCgivxH7VmUCG43zUEdMheo
kpnlEBJ/PNAoHjKjrsrt3x2jBdtjYtWNUMJ6t3T3VN2psWFjmkHUOJ0LWe4U1tmGVwbznk6QhuA7
JKs1cgmZJk2vYWxgYi5XnzFSbNPEcGOeC2YtiJg3f7ey0NShf32onSx0J9K79GCfWyuqijNiMass
0o8X5Jf8O7WwaRO1S9mthD4VPddRE5e/TNt9nFtbMUft2yD+8LE4wQHkU7eFoGd1rHsYxdXkayfN
pGSpqkrfYA4Y07EvRz37Kdpdvw78lUqmpxhPjTDbHW33WlIrVSAvVaDiGXZopdiK1xLxTwPOadCw
5NWbWANsQnejRZuCTdyrReTnYJ20Jb6z83Rh1vkyPxi0VqN00NSK0GzTOYqmvbgFx7yaTtzNOuHd
ylDmFhnLJMdX6Qvvylz8520TNa8QJyywtfcjpvDi2xovXzBp1wHlKjaO2p/Q3GlaS2cwNGz9FfHO
rJz09U5ASclu2tb5aArxYPuM8loL4e03PseqEeREVkGVBP+9MhdI0PNGv1Xd4+Ih1/uKJMvg1BgH
b2magXArDbQERZP3al6M+o9my9t8f0ahc3FQSCwDVBg5eUyNGSDO/ezZsPkmm/+EktfipaRSW07Y
KmQFxrMFMDv4XKkXfVq9uwgI/1aY6iQ7srBkNMPhzjxPQ75ky6OpQpBh24iDe//iVIRPBKtomVvq
kH7VfPJHNUa55T+lsYpZ6qcGwSjn6vi3Gs2ST+ltkFwZviHQhczVbgSgS+wF0EivU61Wm4vFciNd
fgz8t556npHJowf4mifF7XUYU7hG5W6bPS0rpWl9YJ6vZ0fLB4PDSsQNoYrEY9OsC48EZDGc024f
618T4nwHS7sYh7IxBo4ONc8QFBP+PHoObDlvLn7qcBFDxvvgwNYokirvv8pga/s8tmKq/MhQA5d7
5nm7tB5PP/LN43HINQqDsi2DVobDHKSKOR/OwWNkus+x+sy123hPKkqvpno7YY9FxefzB0j6Vmg6
CbTte0/eYxbckIK9b7WKmCkbsZ6SRAYcDIDP7OAbsbKnD0vXBd8bu8Y41RDrHeZqJA6N4p2WiytC
gkSP/BCkXNMAvMSNslDxlVArDsAuMEo7Z1i/nOwtWCNxy1M1E9bpKZOu9KbhC9OFbGDsNBoNZDx2
zjn8lE6x8qCANYFoglbvsGh+DUsQ7UF/C/ihhKEJdCxDDY6k4k8idmZT5s+EkxIMJTMeCNmKxBjs
nirqCZODBi/7giZiTlptZ85yJPLDJJULIR4/NdieJGhxKE+Fv8hH3kuT439mIXJssD5RMyrRQaQI
scg835kwdfKykG8WeYtAikUCjl7EeIGxUhtlgXMJJeJJ4weXxfph8y75UXNLt0NgI9pXizkSm+J6
hrPKaQkS0vwNlpU2r5wg7lBfiCB4/jCqsMWhHWfWlBhD5LgIT60JL1siAsvrt1lHOPyYjZg7oDls
T5nIAkrI84J3uWw1S0nb75lp01x31HzpJgmmBAieX9XFkp5knM3MUxzYCP6F5SCsRANtQ0H2FV1+
agxEIdeGOLRM/dVCvyb8EKyapIUcRcIbHB8QjaAE3BR+AD+kW/S+IDT7rkrAsLXVRKKEnLR2dztl
oMt5ua/fa9RtCEKX5THxy3bZ3yq480VvWuPdgjzs7EcZdLJjFd6AgV9A0uS96QEhl1WRq45oZ7Tm
PG1iHlZfHwUDG3ctqO35yyVGDv3NfX/Xa2Whf+6YQMbQOBBRpD0TYrF3OcJPzzzI39jlAar2s9lq
4i0bfPzeufgyLxrA4CeQw8CPszLZev7osM5KJWR99MbG7j6tIMARNuzWHejMvZA8ccyZsqnDC37k
XEKC1VsXI5EYSTCV9EcYn7e7jLTjdaEUjCQ1ogznoQhpmG67/1AUYFdoctzDtLsw4ZzvG74N9zgK
HK7co5q9731PSCo+LPJgWl2qXaUno7/vdGAa32uguulTnDwJxRMXMvnzkJEVgn5AYfSGEmdfJSv5
ZbiiMLdvDdQTvscw1UtkxByQ5WFMkdpG78M4EASg8bvtemDXcFk8zMY+hZsjI1gx6YvWzDPqPfp7
BgHqMtrKOnK0OIwp6Kp5COwrFt4WlekOJSJg7S/lwhpGuZT7sQSaQspxSUyHWF/oz6qh3QMHH5Dh
9cE8ZdypYrAE6vZmbz+6zCwd87eEHL5gtnNLaC8ASvDgLCWuLyjw/UtFDYL0U3A7PSKsV41wBvPi
vmihd6bzlCdW2bKtPS2DcBmn6H+4ByEPTrvsfb1vum/NUH6XwOadmnLnR98qW0ucJaS3ejZDftmf
DihzeKx+vWeeOuawtAc95xAIETXqjneGhwVY8VOKDkGVw7/k2kVG5HCkcIK6Dbz2PBRKX7ye3t3+
pfUiITK6xnQhgF9DNeGWkiJ9A4vxhvQVKaDeBkVS5fbSE+3XosS6AJFvCB6knd4kzRHad9dLvtMZ
zanQ/SEbvkrrVsKiR8tnojSw2kjeyien/WPzksdV75+oOLIZrCbHZYxgLYFKsIBOuPw/C+E3+Rxn
/Z3cUdj6ds+PpWoVFerKeUOpYgbS1p4R1jlQpodIVjxGFsmQsCgJGvBqYg9COYuqmcoyugNiZ1tE
6GNzmsjH4FooBz0LmVzelent54oZqDo97GhBHQTSwAqy3eyjBC/qa/DOL4ha9ADiZhIPwVASDcd3
lZGaWtd14AqWAdUiUUfMTdlYL1dI64kLqmV6bz/IXAIe7prBWzBs4om5hBrLlmo9cOv2sHUVgM1d
13l22SiWb6dSwF0LgUhmAEVtxp49MqkslN2pAVgigb5dD9c+Fv+bAJy0wb2AUvjycu5RPQo7XWYo
zvYD7f8/p6VZLNyMoQ0A8/p3YvSGiGNlS5s4OG+FqYmVhO985N9UmFeFOL2iY4WHeE0paWAoPDgR
UvFGeSXw3AsE4Ddc9iTKyJBkjHujAqjRRM+AZ73kCkkAJOZdPoAsrRVjQcXL9rovDqBOn0bvxNSc
YLAODiAYiFIO8l+8c9LEFY75A+I03wPgpP/Q2lg+N9ygsD52yTG2Jr0vFNa09vOOO1mq8RisPVO5
9KtQWRCiSAamB1c5JKQUuMdHNPg1rQVqCJczFG0hmL4+LmlfdbIB9fIGyaPyY7l4FzHgy6QRDoAl
wFrVh1FJRlsC4ht4Q/xDf9fys5xDj+gg6koLa0RQwfzhzYThTrtgjJmeLL/cmgX5pvDDfv91LomU
8NOlNRV+7tFSa0P6kzNQJhKbwJiH7cSoWE+qOwt7BtVVB4w7oY3U/rp53rYsEj5L7S0RI9bz7ii1
0fSGIgumaw4nCbWSnZFO1Ds442QXPbuAg111q2PWk+LKptF0uPyjTV2TdHvBa+PzS2xoxYkgUOCo
z0qB4/6xOLSYC2z5+ujPtP/AGhZj2XXUEnVJGwQbvEgmeBkDQfdh02xpGC/xeutfGWc92hgEjakN
RbQjkTkH099yjsnTMzFWs4tOg5yhiVSLWu6vAndECU/aRJYLV+6LlsROgkYr5ohSI2iK00Zr9xue
F9FHJe3otyVRqirHiTTcNDy3o4DwGNHktHio/fLIelxPO9pFRun0FuRCceg2trqwUSWRYhW2N+l+
hr2CxBBV80ARe0aJVUi8SvJauc5A/aE+pgUtsB8FARYP5LH4WzpN4e+XhgpBMhbN0Z+Oq+QAiLoe
xN2ju71oEH76FgQjTJ4XsNcYozl4GD+D5btyJcr3i/o8qzJ3+ZoZMnGOhklNuU32h9at9z0DQi0y
ovXeeXPxvA06nk/xohhp5+mxpkInS8a9LSQuqRhm/J4xyuRn6pnm0NQDH9xzHnb+grQB6FSsohNa
ergQhldcf0ZrtQ+F9UWXL+XJeCEfgq+qSWEdf5M9qnZfbBo4XumWpCYr0aWD9oCHAQkri1s0mFtr
paR7lUxJ99WrfolR0zzJKhB+y5aIO/h68Ew+ZPK3dv1bX378BqEDue4rdOnoOaaqAqjw3AkwlSBQ
Z5xRtwif8w4Zj67OKIC0Swu/4qDR9t/oxNQHkvjmvdy84jLQ89pkPXYxlcJpDtASmCtg0hYTVfX3
s/pmcR555R+B89ZPVluc7sJS60Syi41dMKdwkl48PutFOIANt9/nsC/SThgUk6zF/u1Er8FDCfW/
gPQz8roMMQb5PEcCy3JM5L5bKjUn8uX9VaCGJbGzcV5vpR9XFquCizmQxzIHaZM5FC+k3AJ6mD6t
KHKS9rIFBBrOz+EwINS77OIQ+Dv/flmLljEvzAAjuckT+hYV5j4dqPQ4jGSh3XqkeSxyAb4Rlbeu
W/f3maGw57s5oeNMxWUrmMaCglF7v88jGCr3ZL94q2N9Xkm19L7dcjdemMg35YtYMe2uF7nHUnJC
6QO62Xbr+3J9vlw9Ujw8tkH/4yxXIdLv4vm39Az8Ddo8UQpPkJhC4EuB0S+uV0d+E69xpZ198m68
R0pM3dRasjIKGnfuwgLCWgSIkmzYjB6A5YQtmT48vrCq/NMQZmzOYufZp0H820jRNq4H04QGX9mp
Y8mP4P6WkDIqT4afeU9CphMd48XvPP56lhuioqjwcq10nirVZuKcX+/8NVzG8LkUSMxEsgFOUimA
CjzbCqykfj1eDUrJG/5rphhh4yvM858BvGuWx+Y5hYTpUHITaeU/ox2DqQxzSUvltpOK7+2l3Ufg
g2gkRz/g0LXDIYCwZWjm+MJ9P0EjRhB+SRUBuuFQUcR66wqwUt2qjrJmVPu3bWC4TwysFrPKxyDN
ZIjvcm9BRYCmVDUGPwYM2EzZ7W2nOq0GE2Hh9RFE1kf6Tj0uOuWe7w7jYLMM1HhbZmSTdVh8M1/s
Vu5MgXD+a8//bL3PuNDMeGwqGO7dgC+N29PFpC1XhbPLF42UjQ5FcOPeCKbo7z3+uwwR2M7gEg9u
Pda6ZZhtD3+18t/eOembOKZVRg5YaoC6C+y7P+iNH/Qxk7PJbZH9lIMmAdDXORzGhKmrqk9yKwpn
iAYABaHOSAXr6wfrOKs5HEZW/dIKIci+WKLHWHIATuyJxmMCddI04y5FtU5iiy3IM2HP27uP1det
b5w8UgfZSoUjLZU6PUyjg3IegpcYDr/cJX0iMhEX9GzUFxv0c3L3OD/cGnEVmr6OgTSLmv1z2jrF
IBSeGLfzPYg75MnhscrGuk/760x3hSG3llmX6CZpzIkM6hc3XyD3Vcg+2dp9I/Awofr91bJ3aQJZ
E+791kAdTIGRHkOLlHPr+suatAUisSwxmqBo7C+R77DYhNp0mMgvhpmqubZsP4u23zh0ZrUTOdfc
BVwJA0KyyEMgjupZ//FCuD0gmnR+83paYA9W6+SBEm4Eb0rWokanBB0FMlStpPLwaMwJWaBSriGN
cIVHxo3goBoWn7TC+K5QB62KqoiEexhLN4rFEqeY6V7WTgnq3pYpu/X79F3Lq0B/eIWGaQdu7Yas
PP0eJejNZbcqyYGDUoMqbzEj2uZ1d44Z5wyTnMg3//NALuGNUxqNE2WadQvIOh/O3IDobG9m3YKE
IsWS9AklAikXrwqk13zs74hBIudMU+hLA+scJ/ACJ3/PIF+D8a1QZTRy11JQvlFbn5XzblXGUtXO
WdYmbqrUsNuVKUSvwu7aMbxbG+LD040x6IxJG2h/qh/YER6QAc/gwbhWqhADkRDyS40ofhRO+Y9c
2wcCvJcNuGF+6m304MZ0jVbYBJKJckThm7QTW0hj/3xJpzFw62v91ksN8y0r7ZzbqJnxwGZW81SO
ody5v/GB96MI5rkpEbUVwejkE76933U9D3cB8mePYGhwzp5lUsfNWVCEw4d49j8XVNY39x59sjZP
NmFK6To/m1Id8WRGySTxGWuYLmyLHfBtAmvrZITwlK1faEMUmsOJgXMkrbSNhpX70h3kAq/22jgN
O7w3geQDdjjKH44w24mCBbTU+bZHuJ6UOIZMWnaES7i5h8j0HXj6pAqG0KhT2ykFXxQOSLKxKmvK
SdlU6JQ6E0Uzh7zHgziQBpj6A1u76f5p4wFB6EmI1pVyOegmT9VVi9p69s7IETbwNk3HgYQELzL3
Sg/LW40To8YJAzDACz+1+jGB8/6oUfcCGmxg3YMSrP1Cs1iyZBkPgMeod/XghrzEtCA2Pl/hJZM7
tAOQaEc8fP/SYnxj8dEYB4UxPrbvAzt4Hhxdxom69gWqqJxhxzCELei8Ju8zPZ4rL21YkbRFYJqd
pwxSI13YikeR85VeQ0BIWFVgsG/qI/ftCwB7qTdAZsN6ai2vPTlX6R82zWFnK4Ky65guoxDKid5C
9vRN6HWAQCQSB0J1OqfoMq7zI6ooqVqf2WfNLCgJfjJ2ta38VnNZjblUwZue34BxA81H8moG0AR8
1iIkW14QJG1KHIzOPI+UWiA+shMYo2/VDlDQc4D4s2OwQyT4zt+B/7VYBIq4g2JfJ/jbJRYLAH4J
FtMFiODVilmEtpnTJaSpeICz4QmjXomXF962WvBArm4xdiSPddtB7HX0FXHmNilNffSS+Teyj6AC
mVMmVDjXQLXMxSIgtaZsjmdaKbEHN1TNXBP3Ws9ip2DlYMmpAeSuslRK9TD/Btam8V7Uykh5ASrT
oQdZneK8GuuxAQZAcNumQYBZi+bxZRUWng1e9IkoMDHG3H8H77xAA6CuQ4QKwY9oJrEAyN0LmzUj
0GVcjoWnIJe4EbfMtJtQrc4N5GP3mPdAaWxJuD5CXgD0P2HOnIccU1qY0xk22/UMkx+uPEa5G4B7
y3TO+Xrg03tOW63/hc1GVWzpKdXYmZ/4oaGq/AKLxkYkk7OBFPYHIIEu9DOwHY8Z0w9WtL9aKdQl
EUrQ7QtgPaQWS22GLmfa8d+aMWQfiuT3TF5AOU+i6ZzdhP+CKwmz/9XWJFEiwSMelhrmccUAtV1M
WZN4FN/OFThIJXZ7G1UEBaytmfLTOoCQ5Uinlc4nJAIHlYVlF1XxtKTyfnPHf3THeUP0rLelTAsO
GLLRzWjvceHO6TPnizXEl3dL3W5OdtzCqIuRyxZPMi4gT9r8efygAXZViVmg4Rz+03Ra3crxjbR7
5j2VTtFiL0tcoR7szOQqOsEsk0VDHYfnudxQUsNeajs3lqctv4ijpPo8xoHhh39H/P32xmbC1odP
J8yXQZ3jDFeyXmQamcgpmz0q10kHtVWonFA312Ckl0k9oZpIFQva7oXRETu93bRi1aswloz9RVcc
6zmNvUKgmqTpI3u3tac6ShgbLucjsC1BwZ929bwFYRpLLMXWoFcHOndhNSZbTg3B65cE6thcvVGB
VOi6D/KiVCxF0/Qjw85pkNt3km7gmpIcoXgTQSjJ/ycdXTVytWsa7CKHyxAfKVqiIzc4OsVXyC8p
lj1FJog3k3ZAoqZLPBkTNb0zQQPQY6P9C/bSxrse+3KKnvhAMjE55HQdbj+T2KWOrs9iy6Rj5qvq
nTpfhfd/ldU+EWJWrO5e8ifD1VVp+B4X9RUYJAESJydCZWMMaTe3Kv2dhW9JML7LqLLkCbh8YDeB
h2UiZRNTBpfCe2Lslt3DybekQrGMOXwvxmXCt0V0/dF9z1GacPchfsbVCcRTrl7LiVhKxTV9HT4g
qaODWbgHmUWQsRTiqP8xLlIH9Ri9uVoP5NZ7vMgfZP/RB6HnXpW7zrTczWOoHfENXQ45K+dmZt4d
DuUa8Y1TaQQww+EXRMFX7qkEOYYTlcVbNxNsTq/76ysn41L91nyGJej2eOAryNIF+i7GAvNk/Bni
mE5TLomKOS7w9fHDvTojhj7IIUopVENwyeEKooSbhauIUwnQ2n3yiqOOpb6VokwRd8XxkNfs/1/K
lv3vpXJrvF/ckzwxt8W+GhodwRJi8AwnCdVe+lSLDswNQ6qrlu11yKm872qsEVYHi5l+AG457UTb
GHQLM4bTSxVfp9/K8LhIhpod9OORtmM0imn+pEfNlS0/C1tWtto2rrFmOc4J2Xp99UZBdEkmn3i3
dfdFVe19NJSw8wsMT7+d5s1C/17T14Xs/OqritAc29dsoduFXCNi8MrQQQ/9PvqFxHWKo6KodlwI
xbhLHOt/ctykjVxsBUgBF7LVUSu2JqLnEJFZGeJBlxbd3BLi4kHCSTP8eZ4INYw6r5iPcU4+5WBj
oOg71LKkaYIpiq5l6Vj/Td0dQgbfVlRd9p85C0cTLx1OIP0VWMUrJaVoN47irOQdA2ZpQjgARCLq
BYuPohX6xiCllMhrvQ8Zx0JQmboOuTsjIkZR1vJKVd2LkXKAC+CkqSAi7BOG95qCc840XtX0Kyba
/RwH5DZl44VW/whh5iS9Z7cNxmKtaEdA0eOKRUykLFrqHmhjF/EQfkadsYbV+j7yfSiQLR1iA+O4
DQgP2BTnHCN5ONQJkvsDKZfpmJ2vMVGT0BgI60gGrnIE1DDByU3yRgXDAdJqS7CneqFB/9r7aWwe
bx2aHjvJltcJlWkXE2D8pn6UY9qEGKT0kqtNmgRkfni5Xu/2X1gdW7Zt9zl4yZWcLYUfrooGaqGO
GyJ0OQM76wChR3vh5sAPLpXsA7EDXZQ9xOUilVKNiUPM7wr6tCBURlYUkaPs9ZdTBOpy1+LocS9a
DgKLvwsa2Va1/JsYfF46ROJtf/BiOl2Ck3Oq4YeDBd3D/c9OmXoQ9wLJRgfqjCyBVtUutEGhOLcf
wLWSDqRZ+g498hr28lYZtdkP75URBsvcYrOpeyUV0s5xjJC+X2gJvybZ4bugUS1RPE306jMu1NTt
K65IwoL2QoKcOW4MyFRYjtlg3hImbEc+znMUYWUxriik2g609NIeFNokQiCoESJfI9eyB7qmzsFP
+Fq7pDOE0ipRr3lFj1LKFlUlcpO5FIZ7FD2dgm1548zVPvhRBPuxUTnBCFn6+KijStsX35R5wJdy
kWo96kYGnBFQWry5tQYD9qaycIYtID1F7ofbbH0BwQT1T3MM514AO1+diC1xhSwrTxH2cmUQKzQz
oRxg1uK62OBQGgRVsxCCDNK+x6TEcoPBwB+OHXFXhRWUARTmB967uXHcT/Gu+MV++ND4BGvr6Zc9
7sRp6yUorHDtsKng2dIqMLPxAK+yM22g3GEQ7PF6J32wFCvZgCnyNMf6s34HioKWn0perubWIJKm
t69ewpvzJq1n6s05GQ63SLz9oMwP+wwinz1rfpEtj85aeJcSnxIPrUFgTQ69QA/uLTC1LqfYUGOX
xJH1wAJRyrbX4D32I00A+MbsL08YpaCZHLM661GZlLPCPdr0PIRPGSzP5PDjsRwzXQ/EuIyHpICW
pfTY59bv2n+XujQUE2Yg5DxQy2LQRzR6Hp+nrefpySMGac6bu0SiSbsiwMrP3zsfhJtazXkM7PMV
PWaq4T7J84mpLlnkEPvINlrSV6nHbDc8a7uu2cusZzYLdNlfUkfYlBYFahX/RxF25INVE38zhLAS
or9UXZBm8Dll6wcsj83LaDqdk2GqVYzvLtEPWAAAW9hICtUdUL+Wlvg9+vuyNughb057gwMWfJxp
GdGONJcSg7YZgRsry4FyN9ZMNtJsTRm7iW2GZ9bBRl9VsbfCw4wvfgaXdGTzIu8aIHpQfPLwtL9d
bfBLxD5Vl7N4orASmNfQkz6xy0SKVJtkI/eJY5Op2BjSEV0+I8G6ywnl+TN1fa28MDuJ2J06l3QP
EjHX5W1vLvO7Z/YpMrjEh5aXdyPNX+lMRoEBuWkBgRPaXCvZKjFJTugFTl29EXF/fbTVTzkNLF/M
q5GCWoCfsAQKPMPBAl0kMxIjfwyTX+GZJgemUurYx+6SgaNn1Ce/D8WHKuBRJbQfhWGdHnCnbH/p
UbMq3D39CVJm1OcGIJYIzHCiQzIRFNkSveB0LqeUwcmTwPhhAsseuwf0ZhwkZTIZyNB7A2CBAVCA
hHl0ibiOOzBENfZPmVeFmE/0RXF+9bnVSJfrl0eth0khvg4iNrv0SJqJeH6Aniua6DOHhzUvom+Y
9FkHQj/PpgIaM2gGsl8lCfmfabSZCsSXnHvNRM7jhQJZQwoSy9dhafpF1WCrJyhyGI9uEACMgI4/
WnDiNW/uxC5yLUW2re6mRJ/cD2F2kMOsPMYLAcIt+NcgEYXNG9GYbwHPZ0Bz3PI2CY2MxS5hca3c
SEIWnVTmLMzXv47AWVOwxZBhX7dJpvJvcG9lOHO7JFpI39kCxXlVDjZP/FonfgGhkYoMgxeVEdJc
vOLxJ578payQtCBIgwOaPWjcdLyHvhA7L/5sHgxv8Jg+jYGj4iWInP+Rosv6FeTUhvhBHz9iRFOx
/dCJVHwivhxyOw6/nEXADsIWvFtXzI1GfJ9G8RZSyCScGOQoTqF7E9IFnbWsWu+e963DvPBu/JeP
BoLSckC7viwaB5S+BisKvFcpaJNc/Fvy/gQAfI5v4FE2CjNWY4fXvsf2BUfiOu81Xvfiz/i4JHH9
hzRIewrj11aZ73Y/2PqWXrR514y522CtTbEC7XxXXNSuhWJYWvgXzmAvWnchFUsQVAwyF/1fGJw1
KwjbWuwODGElFSVYIx2pYa6uKQz2byK+q5G62ih4NB1tyxB5Ddkv3o2ngqwPV1uTO7exf/z5yiCb
aDCMyek01UDPdVjHjKsbpr7YB+giGmbmkI7X7/oQUNC17B23996mo4hT1/C+CjRaoRqOwHHZvOzh
171yfdCqTzijQT5mwDb7FXo4yUJ8QRXRLD3npayLzd8WaxsYTbgMIpLPsRn8HHht9K00PBt0V3hI
Vpv1BHS0uONbekiDLwqLZY5NSnGZzz2j9Bu2QuhNIWA1shn3Fhg57o4vm52EIT94E6WOIIHAZnUf
HdF4mg0QrSUeiwrDTjfPqDEaHwpQ1+OCjavVV35Cbq8wG96QE5N6jxS3W1d6cGWZaBqroIBX2UFu
Nwm9FtbZIknipbTmMxC4/1uw59CqqkT9Y9XIamMbO+vLGkXgB0nvBtylwPaNBexjlHLxoNAGyNub
5XWj2jbNCzrnYVPOlcuJyyea26vEJxxFdbQ6mRTm00OItzSLTqn5NwUxHw0WkVvh+R1p7o+C9Fds
n068Z4Gnze7UawuJtjx6btQ3nRIJDZt+KN6QWzWZoN3QJqSi/BllU+/CHJqlnppZvh2joHDEQOzh
x0lvYGt+I9fWcXV5bumAcCgTKlBpKjdryfU9qGAyctWlx/tieukt36YYhnRvXz4HcqJ+b8T5ONnB
2+ofn9Noqp8G/ueRD93SC1WNGRUL/HGsQ77mVSXo4t2KZilF+pOC6E4ZrW0da9OfB+REv0DbZsiI
rYummxbcrSlEbBD81gQNlpvoE62uox/3Et6KciofptJOqKieHA5CeBz3WbgIA4WGVJomEP1jdrb6
ztABBVUcUczP9lt7TMfND13GtB0GdDu/XX5NMAAZAK9hrCgbepNXBZFeRdOI4lS+tHtOHijXLPh5
cD1ADEMQsvV+n3K7dGo9tuwI9o4M44QMJonK8tgUj8EpleAdXEBiUm01omdTNB1CcRvzaDG0C5j7
ezGpcfEE5AO3nJU7E3CEfWPK0NnTffB2yy0Tj96Xt0GaCrn/4dq/nRm1CMWBEAw5uULJlUKbAVTi
f4RwsSnFb1diSn/Z+WevMmGt7eG9BxB0zDhtljT8VbJBnhnCktOAn1xt9j3DQNR3+yHzLAhd+qbS
R5nhFKhk3RUuXmPa4LN4PMHYIsDo+Gj6U//rGkcC6Z3VsEZreVteu2o8qn5fpnlt0DMW/wpsZxxi
o90+DbzUPeaGyi8iNAcvow/gxXiNz40w1R4ozbFchCs8qFUgClzzYkgXmElm+Vkj1JhrWGfEBWa+
cr4uuTmRhfzEBeqG1zFAYA+MWkdpTRhWSflgXoisw1RN9CLgaNGx9l/3NmYTo+gsiPxAhV0Nj0v2
JQehPigG75IxKBx4at4xXjYB3eABXuhb00XAXW6JvylIAJnrYDCS8bxGIz4TwhkufY7XdFIdanD/
Bxt+zidWp6beLx1ug/4L5OptXBNDZtSRcbklo9KsxsMBHUbZIzPeQ6R1I/P0xEmJTcdqPNXDGycE
cBPOh7+uM46PlPLSYmASFAbfv9x4ZS6mC7EmQJ3BVMIv+f1cCtzlbNLkTXnayU/zVgvOuGKhz0eK
KSEKop4Ghh172EjgEDkADpW6DRpuE4u59pFB0viXy0Z+O/FbjREdGhqRVWokQu75iJernuuVZjeV
bkI4gFEFnV85YLOvqOS6FcVnqCwisjld3q+Dvvfll5vS8UNUaqyn/pOwN9cDT6eOV9hwdoNSAYMK
dIHNO9UxjScOtkLd5QmJf7x2Gb2+jYL2FQL8NGCF1WJdPlBtnK/or/pz3NusCNxEWNItDblTmL4y
1VxcN+uNLM5aK7I/X+0VwED9I6h4eQqZbK7dCK63qzlu5AeC7kRzz9f05G8BUz9XnvKfceHsBhT/
vE1uNdnLPjOWXKs8AYOycTrhCQeiQvYRFQysib2lVtRsszD9OcwY9AWdmZJn9WLMfxbtHuPL4OgK
NeLaVUU9YHbfWlPHPt7Rt97t5l7sxHfaJNoaBR/46cm06S1Apt7sO+A3tVeGNumyqPaH8F1eNYoS
WdUur9uvLMqxuAOW34kt7Gxj+wJhJiONj/l070t+nN6cOP54RBCuhiLQFiVWozef3ZfZC+u1LJIv
UJ2HbZQ/BVIhB+yFC7DVhqjjOTUgGsfUjJCvs//dt/mHhTKpXdCaZA25m1H3RFJOVlOM0niKMaj1
GS+P4cqvlf6RuKmJYiFjPY/cxG2qKFbsMbSVPyA84dwA0vcCT4MZnF1zVtlz4aKlQDI5k+rX9Y8m
PjIH6KcUvHPZYJDqaT24ZkwZEHZX2vSvE4alLbiSXKASrObpVz16V0Mtaadu3U4m4DiF5V5eWyLG
UunSF0hjIZeO0lz5+XTDaEClTmC7CdVWMiqoau1cmW46dlXRM89Nnai23QJeQzugKN3ymHUjmgqN
UfY2MV5fHZGeK9EP0bqNzrlRc+uOObHWVb1oYxSkfBE81ZaclirVL9mJVm4LuN9E3fZFiIMnElz2
r+oYLi0wYGoMMIBLnyahg6WA7605cc4ifF7Y3YXpkJsnp3u40xgDFBRJO/yGcs6+RyS5mcxfC5cN
/e4ANv+QMJ/9Gx1awrOgIAZseHZkVPURrRFqH7Pi9I4/4kAQoUcwr+W9heqSWBgn/H8YU0rqv0BM
7QPrSFC3Za8DeOshMqJIAMGwzFZsu3193JT5kBWn/1wWu1/gCbJbglG3zvjTGbAFpL78Ox0Nm+uK
Yb3xq7U7a1ozlQx7HhSnSQCiza6eY5U5ZdfdYML5HLl74iPIb08+1Ch94O/zoGlIKebRy/0tSfDZ
OcHicXF1eGOodFgB1v2jwVgiKsbfLW8StjX2COo7bpDG9ypIKapnUnvWbcvjHnxEz4Vb+SNNC/B4
Yn0twToIvogvq0QxVAjWrN3GnNAmsHB5znZ0F1KLIu7lYSdY/gQPGu3Hh1adTUxp6wOJDcBApGDl
JyK1ZdwcV8+k4euhH/EIDikBo2x+vVspbwc/3jK8qX49BRKYVnZOrzPOy5CJ8BUi6oZ64bImb+VU
O3tstbkpa2KyeYXU54WeQgyJ/LkW29fPlsO3hvXIIXPQWMpOaairyHGzrRFk/avyS7iRe74PPAFm
MaKauSMzoJJrrp5/M1JrvOgx3ERHEel96O00kXJpuFnwd2nm1wog11eGvnTOiJ3P8hYZFhLP9XKg
f91jJQ/ApD/xtACu+2dFoPk7rOo2T6Sp5P9B4EZ3tdW1H+jr9Zi2UPHEOGquAoNQjdgmGplWptOR
ajkPVyG6bN4SOQwiJpGxaBX/6lNwxLNz5/JXHJFV8WTWoqyPYd+jfTtY4QNh7NFaO6EciIAb0Hn6
QqRQyqIb1y8N1RRurruzqLvU8+CXjk2vLVM3Dgqra7ykDioQEMJteba6nASm+2o5UuGshfVhOvQ9
Tr0moxFxgmfRIb8hqlSZOONVdlZdtc+vQMMTxAVCzHYo1l1LXdjsMxpnAk5HkakQswWLvnbOyAyV
gJMNklrZ4YUcmlR/Fj7PTdR3NAk2mRoyTWrD9PWlDLV80GpkKjT4fbx7G9tx+vYZbOEcvylwr8zG
AIyBYPg5hCsz8W4PKV9cUlyypVZdTeTwlApPuURdaBxHTBu/6MtGoSk6Ve/7usLEu8zCq6ZrjM9L
ZCpLBQQ2ObgrodBTa8VRq5uiPi7RTptZFF2PP6qHWyESIqnSuV3q3V9aiYrVRaMDZ9clvw5jKXXT
jniZzpdpSSQmHOnMl4YIGi7AtkBtKrO8G1lERM7yn234NykwmIC1HCA12ZlEFwxeSRNM24kXGCuT
jkzltpE/bM5aEE51xluMh1gRCjXRRCdK7uyx712Q4xGZ8ZK7NHLeaRPFUke4HyPaKSvrqj7xbnfg
kU1gdvUNovUmpaLjcxokal4B0W6NCfYPjB/JFHp0tcyWB9G7W0Bd6oX4QPbistjQkHxOB75ElmVc
XSedZidEKF1K1uB0XC2/Bej/MyGnD+XgIzkNU4/TefNWfVB9xQs/7X67yG1dVIKBWzAIY51DPGDK
UuCBHnOumGe4F/Mi3aFS5mdmoqBz9oOEpNQXg/NJJSLeZrOEYYXiiPbJgNdhO3T1glGYt5pubgiL
MCUwJmLksAwBPM0CiMQ3oWp7NVAsH8TgqxJgdxzTW/B2eh6xwdAWOvUuKSGFifOLj2yx+r7/mNEF
KFag/6mkWyC4bkyRUzWC0lVs1B0A+X+ip5Cmps6x6mFJX0iFfb/o2WkvVcCZGC2Bw6nrAB0mZc/f
Z/e3SMGSBZOP5CzFommATEMP1G2yUeX+aGYzj/qRsyx9ttSKSClaCI/ocH5bGn+yUsdC+9Uv36Pb
+QzGGiEjBoO9ljG55WgQGyLhkjKDM4NPP6VyFUJAYX+giPB8TsA/SGN/xOgEhEQpXTVGdNaJnxa2
1C0KOJP7Yz2WfavPn4oowkMecUYS/HBxOmluIUooqsI0P6I/8CV8oHBjI/kv8rIDKZX99nTgLM+S
N9YXPYr5LngwqBJlRp5yR9Z2R/swq86e8FTgde5iVBs8vG5IE4z5KtfiKVtvA8bLt13XEgntT90l
HOLCbSo4+/Rt+gPm8G0XhtJsBwGt4Htjg78jMsy55FKoxzIcuNC+LMY6GGsJ3fzWCPBgSSiP9iqu
HonmzYidwg+T/JFIVwt0uIj4fazI6K5+8lcSOgahaRXHN6hS0v4QpJMwbgEgv3Znn5z+gw/9ifDL
2DhuPW8dX9rZ5qsPDYj+1fc1OkQMyJM7mJGqKDAinD+TCVNuZdXc7/rRGHmqcbmc3otNXs59C9P3
0tdLVWBxfKbh3J4ygN2lBJeA5w/tnubBfA4T4CHfApaUiO+6uyjMDQF1JIgUhYd6MHcWSasmY3KB
uJAAFMoN6xAiHl9QijDw7wXuTDcIEBIPrJJP8XWpcl+KPfmcQ6VBrD5ao5PulbPYnz8xghh7/3vc
iwP7gWior0yNRDOS3lhvlNjMIYD5BFCY84L+kNu7xV3K2K6z1fAMWBHjOhaS9zDw6L8XX95+ZCfV
HJQB5COL6P89/VyFZJY7KFlDMaQZWKeOV+iNgwyGDcnXnnNCuPK+daq5gRK6axtXLTDyZFZtF/gd
8eFeMvs9Iy8iWrxNz9q8nCmPLH3sS8T4fz1R9PJuNE3CPUQ3MMAZTZ+GOJG2Csm7BYblwfYgY9/9
9vng9m1kX+SmFf/eJh1dFyc11IHo7+PmY2XOCP+bzuXlQT+zDhQWyU74AvdJmwZmmhVkZs0G61tF
FHC7oRDyNjJyk8h32hLcDrZySeGDAgxBvpp8M7dc//3PocygPwsXd+qiQkgeMEhlZ6uj4Y2Tv7VT
kf9olStBvYnrdDU1AM5oSeDA2M525zbTXq1MAQdrl4AHorP6mXZWG/JMohaZL5HEecqPSdGD7STo
2HL1ZUIRMGqYcWMXnBIA0P9CsoqqMywWz3cezLZhsuQfo50dlCMrAyTA5yANEa9NShgOnTQtVDta
1DhVm0BEcaJ7r9VuawQgTrFv1GcKeNJIoexhauCcS5Ky9YmxWhaSkjruUNskis2pj4rlLZ3MptYH
zuHILP/XsGa/LRWtHT6oNbv+zggf2OHV6zhTuUpClLMeJDRXamSCgnbuS2rTE1ueJgHmtf2oWhpd
ll4NNme73TAi4KKrjFERbZU+VaCwG14hRVBi94W6CA9rkrucbUKq1yBpo/Pa/eiIMRZ+j17meVxK
zzhWGPwqD6hEjYD8OK777Vcp0G7+qER2YPTddMqBggJGwX3z6pekOM+eKxoR/NNA83df+4lb3lLa
RWKyAvMZasN3A8Gp+9rBWJJSMlJgfizrJPo2RuM0xtgVEs05wpi0eeNRE1qN2QEsGERLmPAtm9VD
BNnWWGBRugPrG7oztdrjWAwml5onTB5ciIhznpvxTqeg/nmrgWF0dhoLHNbSwFIRVNfTg2YQ32uB
0Wt4bHDRXiUTODtp50t5m4D9esyFSpwpPECd7HFkKXgyJAFv3+xGkeGYnBv7kwN1KQGpVSY3x0M7
jwznZf7f/TbQcivGftKosHnnTo9K753obFqjxfww+0z1k40fspsQtmrFVyBTRWD+OMcQYPzx1jok
khmJRDWlszMwAbIZV0VQa/gWnxnrIl6N4nBAriGyEK+qBuNRbeyPaWtIngx2+rgUWceD5I2xgkek
bmSHAArM48gv1uNhcvC4T3rpa7oNWs/0PHrPEanpRVTazc8D/K/N8acWO2YCoWb5q8sNIGZyzIm6
Aj3TiQVt8w+fnq4+E8OD+GMZcjqU9Zlx3de4sgjrZtkJB5m8VezI48h3AvnBC2rS/WjLj8GU3ayv
Why6bTfDi/gWQSxNvl4e2gSMh53FiJvX+hUFUGDsGx8K5B+t2ZTLq1fQNDn+1i1l4RINzAQs8DQi
dWkL+2GopY+MG8OTiBNykEo8Hheg6uMn1Od5g/+nIUC8ihHK/0Oky++Shff5bnzLjfMe6bTQRvli
oMY+r9448LZoHBnUysa/54BxQFCUVzvvPOBkHaLkqoZgjktbh7xE0mDKovW1h9JH8z2y4GR11XXC
FAXMJxgPpH1LOd7d1NcULxCIFH+/1m2B7jW31giV0nPu+XKr3mqc/C0MMWixJFug0CyL50YztIcN
oYHsOiMFu2hDBhtDRNtDPLP6tvVk3MRIcYnVLMWUjUGrd+dyQXdAMDrRISkdCS/9+GoYHgf2UZfw
Nc5aJWaCZ0p2nSdv/qoI25dVLvGvHPp9EEzaSDLKAmX5oopMSA3WmjEuJ6smYtraenBMM2A3LuKS
8bMlmLwgjTTJhy7zvFlDCcg/t3cETBxYs1yt62A6yjJndYhc2ISxguC5YSkXYavPXZFN5Hy6q0AF
HElbFi+Jbhsmog5IkiCwdXqJg0+H+8ZUO4Ev0FQ2AmS3hHhP3EigTpBlIXdn8xFVB4GobknbolR5
1zmYGjR9OqOOFMGnTn1lBeuwd4pJEoRoRNPLUbPM2CQWKP1wx4MW6ayTlWWl4I7/lAi7ZrHSfHAg
z810J/lUPPuSL9QsarEBJYxRW5khlPZRi9p5xxgoo17/3uqgZNvJ35EnfxE5nk7O/ypHInBweNcS
lk4+G2HR2U3sUaY1f1vONSwFMZt1FGzDqNYYl/cA5WAiDkyMb/I/ubtsg5/cSNNtPOswBGTrdBF0
bSLbcAI4RirBdugWQawiLRlxn3hGAcpv5ME0glQ/fy7Au4UJW9Cuc7PJY41DGBu3iRdcv47717zz
NbUQkf0NqZvCvv6l5DrqGb4xO1wxKX6lqJcnp+0Q4pYtMpyAlacsbZUHHAzKCwM7HB98QklXgOmq
D1cIrSxp5xMPBIc8E3AJZit+o9isv7sg8rXvoLb2JUq5Erjk1ceGj7B8OOWyVe+zVjhD9px/T7oa
O4K4c7OWu5MgwQY0HzD8RGKgSKPTlTjbPLk4KtI/MtN92ErLD2wA6GE0zWY0ZBYbPpdv+WJTCtzC
oJXBRkhTg4lwzZbo1go0FOuSSIyyKZmEmNIsTngCaXsBP0xaFLhhBZuRb43kKB4+kCdghI2TA3zk
1KZcI6ypVGtDt91SgkY+EESQc03auPjuECffMNOlB/LZfyags4rGnH9XZ7gKKKL0WEnPLO0njFKA
b3Bd4fVjOtTLez5OvDk25eMflMwNZwLPDa6uIuI9qPkGmPLNyQKlbquYIGuetLHI3xjWqnO++AGr
Z5YMoyHdaC5PgUfsU9F+UoX7j05rbiH8Os/pMr9MJpDtpdcR3c7kPTC8O5oZTID0BYBDrFjJgKdK
cNz1xjUTLd/88+b9UQdx8KT1I+gymQmyrbDrWVp89jJH11dByBXrnnAkM9Lu2OtOT03A+82xT+um
JHDAu1H6RDtXCIR1mvwOjjKdYYRCr5kgv+879r1RHSDIci8+WQLoq9QnMWQpgsOituUTPbtu6/We
dL24oPqUiDMBU4Z1QfKnDBw+v2Z3tGsr7eBXsQ7m7xaeMkjDBfPkivlXeAwu4ALE6oVAzjXn87C4
N/XIR9Vn5PDSp5Sf+R8eakVZvWK9Gzx7ymm10pLOv/9U/bP1UivGGy1ngSSKoZdlIgS0ejgnBkzd
0TGzZP1tv7Un4qjXYR2keIZhd/ItfstWZwxacm42oLLC4AgwBTEjIBEQy8q7mgiM9IpvH5xsehxJ
N2gL3qzlVAdYJCNGl4QuKdf1deQC6FLQKiiVdk8CPToMU47Qsv8XQE8Rde/VMo7tFQeZZfMHgBZm
94mCVvPFekXaKCBOQ0JU2wxAYOS3WTXbIDC0vQrKoJWUgbYpDjI//LmjsbfqG+k6gE1M3Wx3FoPa
PM/ZQKA465tyP5snt6ZUARppttblm2hMA9vHGNKqbCoX18FLry9Rf7zM/2rf5m7TIZjBsgK1KFzs
7k/XWoqnFR2yhT4I8JAtm9kcggXXgh1I+C3UUskq2zmz1YXkLQIVhopyqKRm3aUDK2G0Cc1glfkk
6v5S94Q1De1STMFC3+STgJf3BNLE0f3caeY569RuYRasr8gD4ap7cTlslXZwBurFqWNr1s1iQGFM
8zANOEjS7u/+dKhVpx1AObgq+xoIhOtPDYYnSwfG+ShpfvVZvL/JkHRz5KSXWq4gStwBV6TuJ51T
CJRSLzh64BKC0zG1+QYqMGkz06QTC3dkRyObrxlvjTPJZYefUQplPU5tY52fKfa1+7lT0k3kzLai
/M8CODhih1UuuwlH3HgiGkDAs20oX+UEV4F1LfWN7uyJ2840dKdHC2l6EBvk1mkEwAdIW7U26vca
dc6y7vNIaEWcDr8IFlq6aRZdjK4sQWHZ3zMqWm4cblCWL/D0IZUucKGPZ2rTOzPmP2h0UTUz0m5f
Zv/2Sj0BYSR1XpX01kuz/mbu3/yJW2h5xzxF0ldwUF0rgTEddetYBtEDyakoMy3iB9RhmnKzmGPL
K0TMMGq8jfUxj2HYA0GSOd1TksKuSi2RConixFAXc8ykdCREbV2NwSv0nEYgaqhBUxAL/zwkmpq3
ArHH1/vj0Zr3fulnSciLRDkuZc5fTDaW/bjKkNZvqItjnxuS7XWPnJAmGqBNt4ALoM0wj9iXIfYv
cQBDoUi6aFqqePDm4Pl5wrKCdiJCVJUaXIHeu1cv2Pg1+gpdUxqPl9WQC7+ZA3GMgdxAW+A4p+9M
EotNGVoCVOjxcWguwo/4OMntJjIZY3cxOsn3WMzaIvjIHasnUjBGFwBVlCyNWpDrSeTDEfrSY2xF
qi8jKptfyj6Jn6HHkVZ/DYNxxHR0Zzs1S23ll9qC211LRqkdxa4MKFhodtHqD2nXad10AGcFZID/
kbDXDoSJUZIUu3TbROkFEmybaUTl8FLiAkT9e4l3ywtK+CvZYV0xd8WcME07aNxdMcpXRe0+Wze5
1W9U5CzLTIwjMdc0Atqw2WrzEYk5jXQQO4PDAjrkSH7x6qSLZKrS3dF+AtrzSoAzj1tyAtLFLGjW
gsU7PBOFkPEkauBUq1ewdlaJcUvOPI8qpe14rC7UogFOOLtt9WJ8gjkOo7PFn6u06wtH0DfW4vkY
AlI29yKg/9Gb4QKxkTe1CnaH62eMdp3YUciGERHrP1Y/bHyFENOPKxCEWAW6DnxpWH6Duu5VrP5U
tNn5bgGRgAeztr8aZ1aK9hZdc+7lUadRbTQtDg0RqU7j4t7m2Rlj29PDwylIrOahhvJTcYyRoVA8
nnu22uWUwboHj9JSwcXjh4mz4t7zB0bfKpOVXJdPqcGhOD1BNae7acNmENn+wqNIc8jHf8VEqTYX
MG6trWNJ0r5ohTUxjmC2ijySCQvjbRpVzS3UdV3U974Y6b5RRFUYlFHem4O7uzRYDSMo5sXYBwLJ
DfRuzMH7XfFJm6h/VTWRDrFspQEjpFXDQ86iM9hwbWmRdkEY6WTtHy5h9hIPMymNM3/VqYXwEr8I
JkIreyt/qWbPdWbZ/qmT49K/+ZnNQwfT9G3hrUQlM92yrzGAsgpAYlqTSkTRI1mh56CNeIET2Yhz
nJ05yjSUnWbvTjdqRcrdoAyxRreuE+0ElPSN+I2C62dWVLdIxLg5FhjbtprAiksioW5oVjMgWj8z
1I9yFKy6Nj0HamP6VeFW4GEuGUzJ41mg5uIiFgGkCw6gZoSgkzU3fnCFFlntnZSpBHckpO4B5ncD
EdzmnOdrwXmfdcXtXmw6r7Fgn0P3GjXL78dZLmWt1Wcv3xcZzaT8UxsOHNVpQaELR4BeYYnLtCAT
e3GnVcGzNXWQvbxklAofV/qVbcDr1L/HT6zi7hjFnRcHKA6PI2fuhsMjCsvjKfWSPN5oTOihRU0J
uLuzys5/2sLSzo/aLcgTPZeOUX/K5H058xveRKkyTitVE6TF7Vll5ls1L8jNVA1B5CnLxCZ5ek3t
V4Htfx0ubKeaECFS8n8VZFcICEVYu38joY5gPPpeQCjlWF3WROcn2PxqyeTo0qCwDPpuCa7uNwvm
reZmOBS9Sb0A/W9WDqcKbz58QcP2W/jVanv3DRXwjUBfS8A3Q5tCWBYhiKY2RKkGAvqUEtTzrU+F
hfg40rLHnh21fH4Z8KWPtDhNxWtjGMUXld0brceDFLPRriBfKMZHGPxSpQ1JC8KlVJLTkmmpdwmf
QZBs6VjNwrw/QlolQj6/+KXo23zR4F8FztK9PX2vr/KxD+4FYzQZhpMKZpLz6BLOriGahwCDVEcz
CJuCerYGeh/4Azut+RVJk+35XOmChJJbuJud+7SE6ihbwW4oCN8lfPbPkg94nuieYUajqJp+PRcE
tf1tXxWnrdWxzYP8EVqc9EfC7RiC3EDcIIOOzWrCSm3ZHKaoT2o2J7CaLUb68RMydZZi97YsvU/9
PXfj8hsEXBEerPkS+xPSf011BJfJIleHeMWzl6yXQGthwCDulVp/Tvw+3IJjyFf6u/zVm+3pnlac
+TQUa2ZwBo5myRROA2TmsGq/KmoJaNJHwPoB6f1rmA/FKsJ7Q6JUTrUfG+hh13UzH6q/NjLSIiiB
okiU6VA+r7KejiBcteyDQzV2z9bAuJwnCt7Bf+nyadw9oBous6rR4rDPjho54u/iiZxfE6UinMH6
P868gn9ptAhJjpU0OY33WRPnS8ggxj74fEuWblX4T9UWQxu9MV9Nlgo1hVe8NR0qOV3uhmAvfdIp
w1gxYS9tfHyKXYFmb64jr2J/oseAuvQC8aG2JIPSVApgCKRYeU3MnJ34Mu5o8xWvUbeA/vfkC3zK
f1/+Xy+7dKyzAXqkE0GQj5bAzXXYuIEQu6ZA+VpKUwk3SSq99RR/aDLLoZMPutH58vS9O8UTUaRj
zsmoKsdZv7q/ohLpTxvA89yjao3cvvBJAeqGgY6gs5+moiLMUkxokZJ/SuEm/NbXHu0JDA2LKNi4
wZ23TK4TumL2ybAY+K/VlENVa9+lw+C10Gk2rdGR3LzOHDZV/i+jjFQgUBfU0TLu2IzX6LWSVZrM
0ASt1jrfYq9tNGHFkiZLZuYkrcRkdticdmUoD413FS1OvNzy8pp4mNoEhpfenTcts5LBxzbL2NNQ
DFETUsEk8ynqR5Fj5khmsrtjUyr52y4JUutjK/8EbZxXoQsc5JNWjNBbTv7BhOl3IGqmjxhnkYEt
Vagr0ZwBGiij8OglVEzy4QHmAhXeAvkk4Y2doHNLBg40nG5y4vZPWsbPhQjUfYtyWDEjb1mbSU22
BaaSF2p94PY/wMA2WCrhJ2d2aSKJLZLEPmuyKqBEDyoLJy1yFLHcFHv0lpxp+yu62I7Cmxvcl8tI
wg+ntKlHTp7swIJrm6LH966EiXqNxUR08q8GP/acfigVurbsiOZdCgp8vYSKqfQqmIznzMbodl2y
GcYf5l+LG1m0ygFlLTPihWzWm4NfpDk5ErOOW52zLq69yrmQeh72NldesLRcNpGw29yP8S8gP48/
ojohbUiUJCA0PhSbMAwVqdAb8YZppzuxSjjoglkX7OA60QgQ0v3K9ep4kzJCGH4RXjcS2wjKeMJ+
U4QdoDuXgE6uu2zkAfTaTPrOOHaNb5Lx2mfLDqXSnZcFiyBD+fvosgzXG6SQCZPKajgafGD0olk5
PdIdKzx2HsXaFgijxmoAGQi7uuPBcIliLnt8TlhHACnWppHAc5qVx+cALBvcdo9B02NL+dBT9+0W
ChpCUF6l6h+v4badK73TR36x0nPIwxFIo0SfLhLiGbVx/CIvD/D+UGmtMCccfJe+84+GYkP2Tn5E
aQKZne6XXGIoiJaOBmZWGdiyJrxIqqyLoluhEpzx0AetmvMgu2mOEkXO/+AalTBWyZJXpxYZoQjB
YGF8YLgPvrfk8vXDRZhLnAD6X6AfgkXtn1DoDBt1MBsWd4BqfmTR5O0rmRbfLHtdwiqT1meXM6m4
AQkHbmuIsFT+wM3s4YwRyJQFsmYn9xzhOylTpxcIluBQExbqCzwFUdHKUVBuoM6YyNva5yAKdMqU
RcaFYfANI9dp71GEpNASKA8vaBXgtfu42ToGn0xHnTByiBHiMhHtoR8PMHOzBiDc/VaBdIgi6h3A
ZB7MA7CkERstPyHNG7sLoll2rZcHSBX66OMwOcm4zh5rZPHrb4iOz2bnjaq840NOsIjR+KIixORX
GvxAwhZ8K0GSG20uQEQT9AU5TiKEmxH863hC4cafdUr/RmkRQzkuLHp4dEW/0YzztXkCStFWAgqT
zerFNNKQlxmHT38sDxG0xVHllYco9MSlczcuSxbxAtN99h0Oja5wiMzgHoZz7Ta8F21Bogi0HmqK
L0VjFtWlxUwbb5K8B1oPqsgDrd7ND6aO+asHgKZlfF3BwBqX+59+eDRCF9gK8dG0NJ6snyLrzx+N
x1Z/MZoC1TVT8C+J4VMXcrfQOI+wewZ9LQe/BCxf4+Em2oKKbr+tqnc6p8wkfIc4+Zlfr5z93J9k
PJQ7hQr5l6h9HZYmYyBwlcd60N5GoR6pp7iV1UfHlUHcxo8C3OEosRSq8Aqh5fdkHsKX8oKzZ1JW
PltmrAVOn7hz8BiQjQfSzEdjOrQTUdfBMp6YPtFABuFJKBbBZifaHByOEjjyZsL6cj7//wxgFDZ7
PghRJNB0D8m2+T1BFlcqIUfY7EcYU6fCAwMYKt+DJLOwMNOlGan218ZoX33Dv7XdFrE5BMXbWuUa
+nOo1j+Tv+50Tux1Cr2htJmjWPHoaHq2NX/JYypV0evgkQoUIRriySOFj9XH3yp/+dGe6oFMBhHD
2OJ7CfR6C1Ek7zw0BVVjvXM7kYQ3gVQSSMWsroHcjGidWCnwxbkxKTmCElO16yGs7VAXoanFGtOS
hYcRnBNhHkxpG7tO+S2KE6t0BC1Xc6OBHzMtgobilX/Vang1Xf8WlIir1IpU4PMBkNPvA5eboNJn
Rp1pWHblf1x5w4/C6akqb5c3WOr9Rg9xiaXDIadLNWLiiBeTX9P4ta5nyqtKGTdevlT0Ikt3yvBw
z/V185nVUnr0Z2R8yXp72KS6bWhir9S9VJdVGmn23qtYSLoRO1foVp12W3vgfl7SOB1h0aWeerAA
4l12zaBNz9MW4NXqR64Qq8aB7EBSMO5m2mpFbIgRzHkh4i2Il71ktfL9yJ7Fm2aQW+VybkHi5MV1
LUEliOk/gRS7+O+qiIdu2rAXWGkjBtT2ddftnYam4bjzDYF9haV9b0UlnQoEiQblGNYI+4XZKlWe
Hj7ewJDk/i9UO+BaOLra35Xls4StGA7+cCpwa6gaNJ9QNMqJy2phrd4LUAIZd5+s61upflZPr3/d
kQTcR8ug9J3xOe1cUecxOtdE9UkJiLKsb4Dw12zpHRU28kronAEGd87AaKBe8glYT8zPlB/+tJkM
QnWsdEKzA6zT4wixWaATH018EvHUjaZSeE/RByZqXW34YK+Dn6yHs1VDoIP2DP7P4OLVNTNX/Ye1
ndFiOwootStY2bzD3uTXobTNWQpT1WYIvQZ9NIEOJ/db3P3lRiobvYmedYYgvEJwz3ILhx61Ikm3
Zs3tkfRGny7oNpzFZCHKIFU6exeKVSy3sPZsb5aj+qckQ110qEIOW7T+tQcDjfN/AI9L6WKBA9pn
6e+nQPGaGC6K/pbvimBzLli7hX/yQbHiaQf8qhUZqe1J7qxapag7Gw31yqyNLvAC8oybk4EVPL+5
ffAEaKGUu8Yj48FMyuYZpqyChkctRbUhQeAiaSfVtKvG/cmxYzWNmPSM8+rAVHFMPeJPZabM5jP7
snrkeyFZHob3xtyxe8bgiiADdEfucHqf5k07OEzdCLthjJ2HbFuWIauyUphR/d90tLX1++DGm5Sm
Q70Be9rqpumjgmcmy7UMUIFGd7Dj/0B0GOznu4N6dlhVqH7Tf/g2gDLFmjFbaEdpJ2UA9YgTycgG
BP4O/PVd+OXAVtqFG4xovdA1LYDCFO/kUJHTp/Nm8kxh9fKF7Ciu9jn1izr/t/rh9qdPL/rQZkyO
phMNE2OgD5XMlMttyhbE6vwCXJChKbxqJ7ohrBaEqLUT6bNkAGQ8hceSdfV9La8B9fQT9h0LoDM2
xXrN9x7y8oZkhFmLlmh792NYINncYMndcHCmgzxN6QvAyxIlgBFRcalldir5S2ZXzgsCxq5n/eZi
MHjdtW5dI6msX7zEtfid8qSIUYP8Vbpv0+SNSFag+1T8gHYIwSBW+JS04sOOo6hj02+QZO1oa6E9
ui2+Ptetng2zLjcl5VH/jBuziuNCs/yAUmjyVQeX/iFV4AnxUip7xYHac/gUBRcvmcNF+ukf7WhZ
Ph3RRjoI/s9rE/K7Ol0UNLNiHbR0WQNgD2nX4/n6GRiNQ9BZ3EsrPxDGqhLxy//aUQrzjLVcN+43
6M4PYl4QJYeiOhhigjuvGwuu7BHwPnQRXEvhRQGTwgy/Cew8bRHPXQKsbnj0nUeTlXGhYA0Z+3X6
Efiz0u/OQyBkvpli9SJ/laS0d3og1YKc236hE6dWt2tjGEJihR/2/znb74MKCKaOIKeySCYaSV1v
SMbcgqGfx75pGu2Ud0etkOX3p3oc/LO3THIOzn36Z9L9yIlTKY9r6qQZYeaRfDYlIlV3MCo9zaKY
G0d+9YpSeOhh0fl+QSX8/SZ9px+Ght67CzTuAkiVGoWF2u1/9fnejIwdQgQnEFJjPgTsA31Ny6iY
lZsILkT/Rrnvut5iHZbBjYbJVMfKr97nQrPY3Pz+zvg9puyD9vxHFpyBIjlkPdxTpeRq9IlqrCHp
8gPRF1vC5c4Ecrdpssee/hWYTXjX9rnIX6UqnkgZF4pudKN/cNL6Xmt+nbQboXVnePBIzwQU5nvw
VwA41hSlV9QjOdJPEQQ0g828mbgdYfKU6bWwz2Nqg1BbBvt2ZLPPIsPDHczYbHmYNZXQngj23K/t
nZFvXLa1RnQLHU+qb0/iUjQ5CeSJessm19VM431SILL2knDDUxMwUzKPznoxJs8tqATDEfoxgouc
lC3vxF4hIzjhMccUSy2MHYfKiHwuxX6gOOy2RNZDJOeiRTpmSnCpXqKbpdWygpsFisDsBUeAlbW9
WVJdxWJheEdUI45zUAslaGYPrO6bZqm+/beei3pwe+2P3zIURTYFTVAG1mGY781he3qIfrEvIfqZ
lw7xNnNkLxeYrX0xupMBcQ2IZTfltrmRG0Q/ppJJAVTJV9PAau48aeHHfMYLUX6kr9u477st3SCU
SI7JBXOP3vGwDK4hjmK9fYRuNKvcuqJ4/brpPG/haXd7WpLhBcDAn7HsCbqDzIW4J03tZsIZmhpT
T3OF5xhXpopVWezDVbCKZ6F4T0rD/DUl+Nxvf2vuwGDARA+ZsTuvY0Cs7Mw3YUn1paAdzfcGW7Zu
Z+3D2Kqg5V8TQrhXJNsXt75KG2mSxN4NPjbuy/ZRWkIYQ/c1hD5bERkC0bWRBumwfWq7TCbHG7Vi
2juSdk+IWir+kaF/OA3LhWHV2mMYRoAPfwYNCjxjKVtnKKOVXTy/NiNdbqFa/CY/nxMY8bvXq3lR
TWF04T/7cMs86r3ZzUu4vQ5ue4/HQPwSEiKQA6LCJHHuHa8ivTzheXd2kwbPmITfbqAf967Cftnx
k0jAF+tRo+yZopAjCLzP6W03UIMKXn5rwKapN0L7xa1LWCHCW3o4I3Y+YwmBTZUnR1fGN5TiQgRM
o27q/ayu1CjR9sRhnVdt+FNSVx/TR4JrYx83NgeJj/xCohRScj1tovx3x4QT/zh9UZ9xc/hg5g+/
3VgX3D6ppqwypqqFYPHuLFRtOucOQp8nN4kiU4EhC5ro7m1L1xxyGFZsGB9i8M57MPYwGn/arnLN
PZCgmY8lzfhSJXBJz6116rIolcP56/4P3FJecyew78bcfW4gklcC5A6Vm/GZXs12ukt2fXvDe5xe
oOOFeSVZW20Ja2ZtF6Rqe410DRrLlLBok+caqC2ky8cxN+Ajy5r182Fr8Q2QI8g2kddRyo8oxzEY
BIJ6896w4LxXfsY+eRQdp186hl6wiaCERE49CNYnQoylJpPrkSQsX3VCYukUqVAMx7u2e8ZkSGOn
ymiP2B/bDUcTUtvKwQwUkIz46NpTZYSePjoOKaLN5t0JJ/elqnZFXKVvN+kqOdJwtOIj/q8wWSOk
cIllH2rhP1IM2ZaK95XQfmM9ec5PCIt8m3njvJwmjJqhh2bgEQbc8zLtl7izNv0ZSuTUMhJZqkHj
lNFqntry/NOtKGWBEQvCO1QsmU1nR4uacJSiH6WfsEK/AcFijWEsvGans+96EJ2nmPecabv3FrjT
86UVMf3tpP0I+Y3LGlI5KNlyAIYnBKRyzfITf1+iXDlrSosuTBq5s6vhm3bQwdqwPNIhn/A9BkxR
OKAuQUT5nEGL8DvYBJcnpwGoFfp7QByruSu5d4OsOLpq858QoxvblcTdqyWx2V1OTHbNq7ufgPt4
y8JkiQKk/qI2rGbKkiq+RnnYo/FLfJFFBbspVkTvJ7GSrGXyfnzaho1C02sSG7OnaSC8/Zz+J7Ft
+M9WcuNbH2FI/T2EkGvMaeSbmey4LGS/7p1//7eGUM8s/jty2LkrCgQ8ywVG2tXuOAC7jYvqdBCp
bXXCobc1Ce80+c4P8kNTkwBrI7FO7fKWz04JuDR60E9ifY2ratQTlSidn1j273j3/p6m7fyLcxAn
AhRiLMMsClQ0z+bB9fTeL4dUv6Bt+HOOndiC9a0OVdTJQAORIRJWutALAZQnSsbQyj7vpRIgYSkT
eMpfZbNfpOpf9NGTLC1Mumrhad3xDRp19yongo9yFmZPZLWTFhi80EcshdoNZcsrQAk3T9M8F9mE
IJZGGPPKoTRdp6rr4KRYWVNostV2lrRLKYHmNC2eBNSlUE6UE8Mt3ow+0wOBWoYg+7OgvgXXHrPp
f2miFb5EXUYbUZCBHYltHJWHOMw1VdPcgclu8E0lC31wdzel6lxK99Al1iGV+T9z3jkGIy7ewEyt
gW5LfJa9g8FhtNPrJWk8CaeUoywSyVeNOVSoVJEN1FPsYXfDypg4qUWUk/BEIEc3N5zuuBH1I6Wf
bKegDnGCsT81pJqC5CmNp1/I5RBqYjudONxwvszRSyYKl4MclfKJAcgd7WbqdDZf3nDkm9Mn5PuP
Scpj1RpaCXa8Ocu2ZlUy1xfXn4fZchvxqQQFSfYDoD7ygZhrpmJF+6S2pTTdguwJhdcA1HoerWVK
D1+oBLYPLSKpxFRQHpD1mt82UwHqCWs5ZXUjGhPp4CVAh74O0HngITtFjUJnZ4afedrv9qzTFDLa
bbVZCDrm6G70pLYrdxNiJ3+5/OJuSqeH7Jon5ISYcUn5rvrKyILdhJEluIYOK185HiawNCoPbnmm
MiqXrl3pLEk70B5CF73NsxAEQgnX6PVk9EHyMKVvRwUEYdjXJeuxO1wY7z4cad0AuZqQq9vCFOIo
7z3NX0++AxiG6/q1elKI+9eJdL5pDeMlJoaEG4O9CCovVlTDoUVkABfTxvGnjJ9VX553zM66gZ49
jGTTBRTgwRvDO+7cDq75u2Kz7hjI95AFtP5cFpcLqizWKCL+K53PwXW1hlxxeLMBqfJIXmsJ4lvm
PTkz7kIjAMEwpvYDXEJEs92YbbhgLG8z9gDEe/iAp+IkuGmw7Uxe9p/CZAu874K6MnD3xIJkGZXo
k6VaUTabDfvFN2LlofpjYsfpa2JA8asLpTcMyA0SaT6LlegHaI6SrRgPamtOh7z2ZXDnEtpSZkMP
ryFLqm3RWm8WXByBUO01Ze5A939mfKyCYcJARP2Dk/gW5Z8h6TRr9LSmTxt4NRsZ22CdkM/w9SxD
WP5b8m2qxazzAWMzfsMVLcVHOivn2DnvhPzCHUbVIda0kkeHoLiiA/uB0mz3z07/f3TP1Bq9ht4K
57dlB/wy/sOmC5F6faTxPKhKpK6UjKnDVwXKUTUMBcTz2DQ2TdLlhCt5QsPMUM7glGs9bt0vDPED
EHxpeMgK4a490PNk7RVXiZz7lKU0AEpg4lksEIvACaYVtK4vpFhm2lbiSbRruWoCLYcf95muC8Mw
HuGSZUvvI/94C8O1T/GkKlf4x71Ecd6aZrc0nJbd5oC4Ve8yow8bbTpu8VcbX70eoNib3zZ1DlxT
fYEigEaJ60tXVdzWd4t3kp2poMQZwz3nI0ldoRLs5/jCBO8jx9v6mL7u5UMZK/tuaS4z+OU/cVJ4
nZ2qG/8MCoyD8HDG2qSopV0QZ3sSzECUtry3iD4GETyf1IywVtqARBKGRLPGeGnw9q0+CB3Laumg
tL16VH1Q4MfenW2D+57/AOab/ILHR2hfAQ04jYraImDpqI17m27J5fJhNZz7xNE2u3kFmmDN7rum
0rVOnlud/lNxcVhQdoyMfntOAINywIeHvOPjPwqQkEYbQZE6rxSzjn83gvPLQ78QT6ZTJVqTmR/N
pNartsFn9XH8Gvgo/nfwT3VcFtPp/raIktuaabok6aOkRSmrfBQUFPX7ztpFH2SyRmyauDBWonBY
cvP7nA8ZZNtxi78yLGXeL9tXd0xRETGUVE8P72k+Fg35ksdfj9Dgm1yx3mM5IEieAZQR5eDt7uam
8NE8Vh+33RDOZx2xAtn6q6TsMY2UlVEi+uL7XE2axlupUf67aSv4lkkk9v8Wgb8wbgasrjcjq45d
///P09aeL9W7hbDtatCLRCSj/lLYNv7rnjojS4OID7ou2ljk3Qv3cwgcjT2OCimn8aZf2YEJKHEI
J+IO+5ePyc1jb/vFIHXYvR5H09bIg1KNsDZVB1aGOJRhe2XbXbD4CmbTo0wCFyFCO22L6nxuvufZ
iwNrnjIi7H0NKzIPM4tl4nnL2ifNpS8ipc568zgk2RDv7ZBvAHO1zxFy7nkbRFewmY5Xf914ZA6N
G7yCzCLrNXmohAIYEML45pr6QER8JkRGAPl5Mr+gni9mPshZM/d3SZFIk6sH4nnpWdOLwrgxQHWR
SaqZagRwKWpwwxlcA277dySiWOKGemb60cVlmf7dkZnttH4OTO8Au91px1PVEF354WR7mp6JUpAs
8oxHLOuLHZ0GV8cnlTp3Sf7h9YygOi5f18kpocBjEqqbcrAGGtP4YE9oSi9n4GdCIUuOzIFpbmPJ
+rGbB76BPbRdV/zntmjNKh3Hl/wKV9cW2RtcmG1PyEMeNQNy26XkL95pIah6TLaeFMKz8eUGV1GT
v/OabIqfEMzM6ZKDDOLfng9Uez2RNEZNAogepZsxHIfdPNOwFvKEGiVyAO568DR27PldR2EYHwEd
knS8b0w8vMPKcULVCyqtoA1qMYJmTGg9EVLJE1P+1Bi/86dzdsQm9S0gogNU7sjGtQ0hQuEsjRkU
JmZYMRgR2/7/86kxKA6bwZcLajTt2Atj498ZjL2SJ871TKYLcNs0eWIF9rxL+Aj4tvxTiBWygmUm
z7vJPo+W0JnkWhtf2I9ncOS9QznUGVcVHRCN1loLgRYqT8M9bVR6BVbs8Gvmg5YZlYtvEi7gDaIG
TkQj8ss+ulH7i8KcdoXhCj8DIx3wr9lyws1cUZhHZ50VktVBh2sgbPcmXTR28AmRzQmzdqIGiUNs
AAsg3tkLFEDuwu4W13zROFKaGkTOriLWmJg8StYzeiIMAHn6igX0ANE3f2uUiKBZt9l2sFV2nlNc
/ILAgGsz2EAQXL+IoEzluhKjmdNK1egGvOeLWmseMv1JlDIPdeMg42ViQyzjTNCSsMey7NkjSSvS
sRz1ZQQIVtPGPqMnBOUHFMfPi3zcu0IrTwAeG2m7Fq8sOKrPgvfjYivnxrrVa7oPZWK5R+wMgTVD
2RO+d2n5WcyxVOBJXvCAPW8D02ZFcqUPXbuSfh114qY6UefBxynyH9HdFHymWHTWiWI48nSp1SQe
SMoEtpzXXu3Ql3PI3jbgWh6nceahldyyyLi8wspNLOMKkWZquQRpHJp1aKpyhSxZ/bEEGna3cOHl
mCrSGRSf/WB13jGyCfL6lVaQMpRovvY+vJ9y3Su9NtSQcojvWKtYLo6h32vC6XbQxo4dVq+Ym7HJ
xxdHK3yZdkQxO9hzFN58Sp3cuct754ajwmoFF/ynproZbWQodB4LHAQvqMLuncc78St90kgyLfO6
xdkmDaMfuhOV3Rnp7Ae2yXdSQj3Gef8ECOoDlCUUHZdNDTdBDsyYG3obGCYPmdXmQ19HUVuWiQ63
AKBEt0UlbwZrHL05ScbEUTA/ncG2Sx2X0cd3hJucCaDeNefwDiiUzQCkdEBWeMQZPyx70PgMuuBx
6bERHwTbZtj8onzZEapGEvrRcB0tmfXgNqVB0bZxW7zYM3rjmUyNiCS23FKx7GVf/OUKxLEH0E7X
aaOXstLUj/Ii58YlHoqKDfQ9f6FInuFvlyNDQeUhDuRDiHsRLZjkycQPbKVUSbBH0cy0Vp3RrUmY
dRSkkk684EdD+yn1LwuAbAR/ZMVYOVtQ/DUelLjjycIZc+v9odyLWxO6JZ5ADdeHG+wG5C1ThqFM
nKXt56cXDxXqiIIuqCjbX0Mepxj8QLNHRQYknn9c/4ftDWIJwhOLRgqnnxt71FQpVact0wRoouER
ZstjBFdPHObYDa0OlAQRy5QoxOY/iDzJzIaZx8RRMQx6k2oqx4bqqpB02dLQw3RfiVgPpXFGgBic
J4N3xYcBHxw/1gp6MDiajkuGxf5IkFLIdlqW51E5+4eWc/hbuBX/i+7lBZc4lnM+dY8my67tcMIO
m50+ciAq/7+DonV3XqJwWLg98x7Fx2A5puT7CDTzMe2iqKIRxhA4oS/T8xqc2NFJLb5EvY7C+4Kl
FzdcIBbWPkMpDIT7fBGgkAsgMhzByErZjj27Rivj9D+kS2ue3htWf7ZSLgOcDM+EdQzBIfrvHkqg
7PGQwYJZmWrDmKqEnkJmAw9Fc/Jcr/6rPUJ+rqQy5q8JNr3sRlZ2mqO5/49ypkowwVuIcItuAOG0
wGTlix41MF84xiL+mypQ1ka8k0SmEzbCEtXaT1IQNbnvZk1dM4c6UnEaA2KSaXSclixcuB4mlSRL
DUp/OKrsAavf3cL7qlO5eDTGKhbT+xHmt7w9wtqBqg2HbMDoQPY3Nxwllt14+S3hqR++PEJt59Rq
mkIInbFP3mm9xUjrfNiLi4CGfxFohVKy3EwWui7f7saD34uIlO2CNzxJZHylU9O73DnG7e8PYXCe
6Hfaz6gODkoi+4GNZ8IXo2EYm66FXbRfxXhr+JbGixxKbXaMmYx03bj5JAMeKNrtEJK6jCGQzi2z
lxsWA8RYaYT3XBEkdElUKA16Kzye78++HRBxcLmVQgls9T939MfRwPOhC9NNMLGVAn1bQPxo8t+U
SihsFVf88eE7WzYHCxnEVruCvpI4qeqeJgnfsdkq8eu40nF2GVSgvCRCY4L4wltmUgshQqDJ3aT0
OFRmgbN5IFmkeQm4QL5A2VuICIYzXgb8LFryVRrYDEgl05oBMbBFgUOvYtZATNFwdT/bKG1y8Qba
INA4jSzq3qtW1NDlUhhX/nczoj2iAsEPjB3J1CeixSMe3FL7ZAFjvJihnknjcgnh40OwWWy6WPAJ
JXYhoow47DYyd7H1kkm6ug5Oft8Y6vm9uRwM3dtUhDMbwcK4Hgn3rlYHDxReTvpITd0p0ohzSthh
M94Oo7k2mohizBOde5WGqnlVQtSTeVxT1c/2OJrRuZDQOIlVIaSsIEQbLPUsqpGtZvrOifrIIZvX
S8/e67/GK8+/DVOHHHb1eFhC3rqDf7tIYjwf8YnaFN14Q7btTdvfEgFQQhZ+jAsmmFTfR0jX6rMh
/+UX5Bpap/D785QRmP17o2l7JexKPz1G5I/M+1g8gEz8BVAY0AQarXnfy/y4EACMqCVtq3pSJZRT
KkVVs9MtW64EsoxHnZnKSje9hLGJdmnAzKgZWbfO7sXlnlNMUkBrQRSRL234UNrKhttHJ2A0Oxh7
4mtgjl/r91RqzpfCmZl+0tqCaBHWWfuo1vrePCSvXup6zaDInksyfl12f7JV/MVs5oqnHwQhAhUu
gR4KxASg1HZ95TeECyqygA0r/AMBOhk0Y53Csm1x8LQ+KytTXnOtVWlY8sDiRJau/UOqQOg9C73Y
Q45wjDC8iuntGEuS7/4NAN02BidMWd7Gz1GD4FvckgysFdiFz9O6tFfnD8m29MusYIG+bz62Bglk
a9MQTlX6jlX1D4Qn9pga5zvXYiXv0YKWWeAJ+SvdJ8+TmlzTYbP3CwD5s0CPhRWU03sslmigUCst
/wQNXC1WLVzke+hnx+yllxnJSqUNCaEmvEHPGIVgZnXiKzpVocfZRWLYjbBWlc+gRLQer/+BOanP
grKzwp8KofankakcYkENR5HUdjCIP7jgga2f3YaYh1CDRVy1V+5dNo9UxqAaDADdY6hxE6wv8mIB
424eov+L7gyd/jWanEbYo7BpEGnOO2XraiifG6tXWVLLrgv4ddkBH70gTqy7Jtl1Mlqo1KO+Oi1t
nHjRyDl/Y4/07THsSZd73nhjNu8NNo3czElTW830okgX2Y3ANTuHbto6b5VRdJWZ93/pNeW/tRaa
+Al7MGAjcNhRtXFavKP3KAJ/wkRiT3CCoMQTKX9rZlkFsi8hbBHn0O2v1T/xJXVwEH7jnA8uq/gB
U2kAWR6gQHol06/etfy+6K1P6pdeiAArVJH+/KRmLgErMPQgxxU4OBvqI9sOQgC7mJRX7F4oBMSz
o6tbub3izJVON7p6O3228WzY+NcRmGyagzOccu5tY5Z6OlrkDFZRyC3dirFwp9EKB5yYqXoEYpLl
nikZ5qdjThkZGl1eZRUiQvBgaH+GWDbsW6PDqezushWy4kRo5pgUb1q2/YWyo8+U6eeJ/65qazdd
zSCbgIT8l1zAMRt/tKK9xSZ6iR/Qa8AkMoOhiRaHLUtcEvSQWA8D+HUFygkMhGMM0HQi6zwEbhY8
MEf2mWJSbjHFEjaUAYYj3Pz7xvSjjJWlPzEeDF/4w7GzA18QOyZSgBLoPYjwgxBENm+gsgit8EMV
rbi67hZqueaheMdWdXB5cX1TKMgch4fP9rbIJoW3H6oOdw8d6mM2Qf7Owww/ZilhBWrJDQPNOFca
VRc+ybzq1fyPff0Dhe1MDOnnaohoEhOc4d4mZqs/KcoWYoL9bBJCc9G8CATr6y8hipiO5aMoqIVK
+EZCmKctXJan2a7/SUTuo11bRfoKEEWfNfZpV0X0JI3qoZhHE+klQvPIFkWdExL07kkYORS3UspY
wScGsEQUtt5DZ28bKGIehQu4iYS4Q8oYnDjmhXepk6qa8Y9zuOILgBHCnQ4uQuEBlhcxKUyibnlf
XjeCQBSEMUz3uUwt66laN0asyNoi2Js+/T9EBT+s9P+SOeK5D/vgpUE3aazQueiX8g5/cliNBbSO
/a13PaAYqL2UtP3ejXQn3D1Oj2AF09h6gElxnLT48dNp+QcYyLn9kR/uVsijV9BfQgxSYoYWINP6
4dQtweF9DPnBFuexXMux3FdyAZ++4CyLffCvGUzUU7uappWLRFpfEedDRnHoPBYW7PRiYYKz5bZo
Rzcg5o+BoQFLEnJFbCp4Xtibr/qGMOX48JdThi/4rpmp/L01CSsCZjiAuF1KdpKREuTtgPyrjFg9
cgUn425C2/u+8+ve/lBPaVTn4Fm6we6/IkIGc9LQ2HlZoHBKFrUNK+/qC/kBYiN7xvzKICdWfnyM
LlXApKbUpKfqg0FV7ldqsiolSGdFHdt4Z4Cu+6fa4yT/QEYCNN6tajArKRch5jpvGt6yuHjg8vvh
hKtAPjU/jbRiny4jn9vihR8PjgEOuVwQ2/Dxc7/u0ekrA7k+w3qjzUFf8LWDVCMwPnRNChfPitN+
VyWYH/2K4qB808SpH+iJyS86vhwsDXncUv3txL0z11RIJ7xbrg6ZrE5EvyMCUiT5qOjQDqLG2/Jo
O3Qzqqo6I1TxlsLi9m4/gwRZvqzZj3NsLqoWrSdC4GD0eQh5G94MkgIei3SAVuezxcvvKbQIP0+3
wactlnZ4Nrs7mpmK1F2Gs7S7ZnyyTfuGAoU5nPeEX0W2DlzuXMI8LSX4XQzDz/+CxKbXjrZ7Geqs
yRkG5fQuvVPkWfpYQhwQCwMXugGxfeMESqgon8RFr+ZSFK5oGSF64llEHwqjOJZ8H6eEH4G2JwoG
MDxq7ZIfiKTquB/wtyza0uWYZ1+m8Wb/JuLXJLbovrojmn78NYp1rcy0IMQfCKIHLupSY+/s4X8s
QCX9drn2NsV+z1XXZhf7XzuezS0PjSapEXplhA2tvbvJePAsJbN+Uyx6WwIAzxJXrJTgpleOcWzZ
UsU6vfV6US6VDAK4aP+x+MkXwwfwmbJGtJa67sXYEx5SMQGa1g4N69AcPPkF0FR6D7TyXC4No83D
r7gwcW24KQp3nrfdsfU/kAFDzAIFMw+hKECcZ1WGrFS8EK/faetzih5YxtLsuKH0kPmWE+0J7sZu
KRWqB930j+caNVYtZ2sfTa7D16K1oCK11tVbN5mmHGPR9gws80nmYFMSjAc2zoGBRsYFy6sK55/R
X4B0QkE6BWYZlFQAijj8I8CAIPaxEOOrgrITQIH8ZvZWAW74sWrKnDbIajmCjDXkXPLwgPjJixbP
G4y7gfZ72PZqtqP3TGFpw2SMTeJ1G67LEzBz8EVaLHZtqww1+3fWWauGS/jAsI0Y4hLJ3+5IOt3q
cnv+wuZS64T+iASRoaY4onKdClHCtEI/NC6YktDbYkuyXL1wFStqdXhbcb9sOCb5yS73t9rp+wxF
+gTEIl6gIggSXbecqrfDkzM9Hp8tiNgXtaWzt6lfI4bjP5+dHJ+gtxJjeqZKzLemgJDkesjG4PlW
9Xu2hReYSwYcf2X2rdvZzbHn2oNuJCb649qNGmoEmVvOfAggYjOXvmzfncjBKTCou3RdEz35sjtf
IeOU5MR8KQNGAK1yFP9dvIjQ6QDoitQ1iB5pxbl47H5qyjTWjBSwBweIOVSu5oumJAVFOK39HKuJ
sw3iXf0fScPulXQIa7SkJAdufw68hW06uRAx9fj0CMZmKPTbXEzzXgYX05XHdarg7suSpLcH7hLY
3NMy52sYpnWaD7oSJm9hYPyHNyu6BEpsFKPaRbAGCJAgpi0slhG3VfUp4t7LtEn0Efe743uioVP4
89xnxwNU+FzULrFUe0/Jy8xdUGDC18XaybOK4sT7snd2aNA+isnR2xXsr/9nTgwuGk+o/dcPX0Wk
TLCEKOLdyeQOkCIhEU7803gnekM4LAjqBLvRWX0QA7gWuibx6QWedoBKAOvvZrVs1Wb+uRJex+xE
WgkYsH5GXRcKXhOZa6qqNH4VVm3GDka3PkIiE+E8LXFTlfLTTbwvflv9d4WpvtFO4vU3uDc83nrg
bB1akRTBY9OzCKjZubM3UL1NJAkXVqAvucY3y2lHQc40Sn+n3meZn976DFrfUbFM3i70aroC2rqn
s95N6GgidaRydi8mqeYaL3qZ3MiYloyvGb4SKMYHlJnJfH1csXYttSk7K3F4iQBQj9f41KOCNj8/
sD0h5sCfO9YeChrctgPMfdFQxxW9VSb5ASErbCVatDHFEysXoQiJSMsrGYvTgdJCKwXKKLXu4SJJ
jSSjXNLvbhkgAavqjfETuqh28gXzOvV9/Nbzud3Xrkrl4BptxSvEtM4d+COmKHWWcogAfWBTYSQk
s+nVXqtiuy3FqEgkZdAv1rblE/H16sEBh+p9H0/N4fh1Kzlqz4XC5b5Fw6hr8aP70AfzxUItw37S
OURzJRBjudtY4eIZXagalrDSjSYcTcmMhh5S2R//jQQXvqBpoVifeLADMw2ephewzymwF0Czoas0
AfJAnBz/RZTAexBx4wrdrDOKwzZypRe5QeVXTUJnQrlzBNmEhPFsKY7K3Q2yPyhbY3HWjdkOxU8V
PPm8McchKOHnw1zviTYuRhcSKoiUoDFCNgwMP+uL2AfFjQImBEw5Mf4pSarTlO7OObWaLX6g0Ouv
bFHp0JhctCwgJ2gEZ947asY4h7wmMgC5sjp/5QiL/h6Qy93ZDDfVd4Mka67H/ttHjBdppzILgxN7
QybxA0yOQHkMdD9CFhs36blrkhoTpsUon4yKGOMA24DlF8R1k8bCd7Ob95gVBHUkSxvUpHG/doti
26q+2f2ya7Y7vqhSX0IjXxLIagBJ7ndaH5xMt/nUMLvQ17e5nvKFNL9TJFTeVqAWbQbZApgJZjsL
sl+AphtYMPRNqfx1/3DskkHhhDyjO4Nv3pJ9k/MyLfTTTADi61jdvYu7M0s02wH1ge0ci/8NjIEu
X4I0C9SqTLwxCI+y1Ggzj293dbMrqn4B79f60XZacB1l0o/5cPGYoEV7T4tcbz767qfiwp3ZFyGV
970/VBinb3ynBPO5IDQNS99GxqwtuC5/IHJP6yLHQaTEcH9BUWxcfSgnQ+yGkrSf+bMx4rTRkmXB
wAcUXl7kvgPk/pF/8CUotOdEM/1YyZE+rsZ/O8j9d39Z8Joh2aIHuHflaHMviOWKEbmlbecH9bie
CJi6E0TA4BX28jpq4KFRX2IyYRCvAdsl7z2AfvKQ58MlIRaqrzl+hmyUl5xfi8lYktWyYek387gw
5/d/Rn7SNPe6gF//0xK8J4XIzJ21cxHhgrij+8KaYtcsY7kiajQi+PRq0AsrpjbRAnYnTgOGuK6n
DNjVNLqp7kaoK+tojQtZOq55lL9lm6i30gQZOaqF8BP/Q/FZRcTSjs3mQANivwg/K9M13BzCLJNF
WtUU2lg39yjQG5E43qbReBBq5OG9oZIrQBIpYxo1puxh/avymGbK2HNXcQMlAs7ASf04gszgDt27
93PY12thVQ1z1X2pn9Rx33DyO/RV1vRRQGcNwyR01MIXUVcS8n1wD9B5wUIpvBvTvNhdZTozde3l
sf4AJWZjO1khZvv6diJifg63ZIXGc6Do/74ZMyYpcJyMVYzKKPOQio2Y5zKT9G/wvbSLYOzR0BRK
PsOKAz4MQxF+/1c0wDllnaAMvlfzNFuspEz5i7wfmCb63GEaQpcZnSvUfdQmjH5++wC1uYQv9xyw
PZWW+CHRAeZ31Zt29Q/Xv3RySPtpJiRILUNr2BqmJy6ShrX4qrK2t/Lkdf9Bu3yGPgCNXZ6oLIXg
KO2L73Hga263boLiYZJQIbV1gRJn+ds0lPgT4bQR5ueuOSWgYbdzAX6Wgz7Hjrcm1M4MDmdUat30
LbuuLeTnR+ANRWJNcQ90XOEVQFYkRDi6nUzKeZZCR621Y9gxjdy+OfDdQu54tR8fIMv3HLla+1qT
yPUSZL5gNDtOH4ZpS0Uu3gROhC1iLiUTZvwcO90wTpwPS50B5liy2TciR3rPAPwdBpuxcIPe+M0W
BmFnfOafk12dguyB+680keF3ZmZJBxdLam9hXmzdar5R09ZGCx6md8EtfasF70NkqWGrBsrzWeUT
eQ7MN+KEEjOi+0Ooe1GpqpE18A53dR0yZreXEL7yMeGVDR7HX46Lpr0wi9r/Rh7EeQNQ/mQXrRi2
UrQNxn4IyobXCSEtsB6zoDE1wdACKqTHzHbA9wms5s2jKQftEXCktTquqDTrpc4Uu0nAa7wH0zOf
BObvMxUMPI7LHGfF/M/YCKTuYejLFI6OfGm8FBlyRfstnx4e+Yp6jVOYJ7ja2EBoZLwTIgGhahw4
DjIXmHslxObLrLNznm8GRC7q4VWXTLBJBSa+71OQX/h+SkQzpFepB4aZCI5N1eoFcQTxC/Aq8ny4
cGSXOiizKSH8n2aNIAx4R64BEkTbXV1yldL1J35+/KpQ7AY4Vnlb62iYfFVu/B4RGfyUuNnhhI0c
ZdNB1btumid2oc19BLSq6E0FhWzmzTvx2d4PN1/v9otXsCeggS3XiH+zZR9Ee8s356dzQx+lNm+0
ksdjEZHgQBdPnlP8aJVq0Lx5UPx+R2Byuo67y1i0M49qJ8N7mvTUslw9ci+0rM0K9JxqLr8td3jx
zUeZh7ya9QNkIqAOzOlZdoxI2Qa30aV7wTdrjWC0cJ6CeBUtQX4YgSwx6Db0D9GQOJ3KSm52PDyC
vTbzVm9hFqSnFUMTzMIiOS/juGYn+sldH8TakIfla1oq9HvXcvuVO0d9jhVbYKI0HAmtUSaMNXvB
g/uyDgN0Y4gCgsiy2FLdXHPz6fwcDHVKc1Ja8AfHBaue5DohhzKJZ7aeMUc+WHqPxjXsW8m+MNP/
edKf2JMpQYqrTweVn7uuMfGN7492ZDHtmZrE7isTL1+AVdi/oX/fFkD7LEaJG/4gOW0gumohMEZ7
aXMDVxIQouuzAEsldCXW1KA+tTahPHJ0S+1HdUciXrY22vzleVGL379lADasp2097y6hLOZs3CZ4
/AWxlsCRvk3zvYPuoMlGO8ydW9Ejuj8UCuXAnAr/VkJ3dbaWMuzo1CqAMNQvMYqtI+1G5CSyh9bO
UuqS2/TcfjoPEKlIX0HofQf+vkVP2qFyxTo3xXI4KF84xNH7oKs+nt2esUB0gNcQIKkglhrvWvra
lKtknEuC5rz3N2iFuGrSqWm2zVGwsXWHIJTv8UN9xoubr7jjLk5yZ/Z3Mkmvh0vL5aLATtb5JsnZ
FAmDmXP7ScbsXAH+WVUX3FgdFtjK1cQnlVQ17KluW22xVyQCzhWC709KkLveCnkfXHwt9IJw/DfS
2fOZ3GiR+UUOSH0VcAN5ufylZCzfgytAWYSHQKhWUyYQwitu25PdjDz5YeFYfJM52VVs8vuI0Lz+
LuPZr622769WcQIJs7Bi8yYMWVkPdQjdsy/MYNbI2nL/Y7opoPVvX2WL/aQP8nG0eEf9dadZ26Zk
V0fWSqV9o8As97P3u7LTm3b+JMa1VMZRuuokv3npcJ7uEK5QHXUWNpJ/Wyt0GjTPF6zk1qFXYq+R
KM8dFVO3TjYmLIvEmyKzYm5C5qxjZ4rRRQPCRQM6yaDFg9YrK0t08rfwNHq3kQ5a5b6xtrNTU0aI
JGotpnZkfOANTRSYcbU0pbKaUN3Hu3Gabe2Dnvk5Gowoz2gI9BbGPLrx/tVlvwNSLE++iEPt1Nh9
fUzFAQvvvuGyW2CeCjgqR9VH52PVYSjjxcHNNiBdh04FRmjiMju940Q07y/Zw0c+UzXe2UYrbnoJ
nuJKrVzdRB/iUT/jMEmilKLkdKIXInp9uGk7neh9kdVCwxyFY1YH3cnil9yYxwjdpS/fhFIUUYda
lpa1INa65DS4pYx9LM0aTDAQTqDq7cc2yHQugHUbziaS/yqaY4kOTP+o/hyPe8iAyxr3aDIoaMkQ
9vHy9A9YfCR3DbDIwXuJE4IVjfWzZv28Gqpc1YdOhZ8ajN8rPkxaIpt18UQD9SKgJ3Z77GJ36R5t
0km4o/gB3iuCBz5iqxUlAGtn4BcWNuUv/dU18vWKTkkCLcoKwcjCrzS2vnyP108ONYw7lEnPNqqK
+bIrQQXgbKB4iOqYohQnaFN28HTJj2ANGAn2tACvI9ip8+YCZGOMQZlvE+Iu2rMhYOXAk1rX8Ntu
xqfmITy1Qwt+ybyaOiCLx2G9iZc1uV+jUzae6/L3bSzBJxOP5E1zLitj1oqerChE/XmvqBvPl7kG
7frvpNJVMdTmmB5lWZYUp/4yIa2xK5aectYSSVgpu3QmvbrYG53mIkQEIzDkyC5fFaf4QJC6rHtH
pFGalx7FBxSktw6zpbvlet4y1s/I0h13AiIQLsaRsCQtQB/rkbJh6ZyFZmmnQ7wnYEKGAVEdpGX1
VmPoyPHkALAxSblbVmTUgJ7YiXLjdEOY7dYDHr5A8U88tCASNN5OFrcyormDPOtexibrvmNHPv6X
BhVZntdgG56S9aoQx1bToKk2aZHGZYsaxFkxILdLhFVTt2FNjt33Em5Vmppdi9aw1qFHz8JKJRza
rxggYMOhIkMlki4IEnlk/66IZOa/mo8WtdwUyNa5SpnEng9glXVJmoRKrQkA2vpCgv8jmewbIs7Q
lf64wiuH37p5//U18bEUiyuqTsjySyJrIS9V/MSZw9fxJjpUDJ0MsnJ9kIIj0fdGshnAyazkBrLz
WnCTMVrZpUa0b5itA1tE0P5uGudaL8v9Z+BiasPM0XP50XiilqRYA84lltjPPeq/5OR5aUZeixK5
nOcM+E26TnY6IFY62CckC79WzFXLR9y1yQ482foe2lsHIldCpufontkIDKXBBh5Zry4uOqORS+4M
IZ/Rv4tDPQiCBuVsioZSmfI62TBtG6JsFwyGvXGB/eW5VcoQRHQHz+5JS5leJ87lESIyp110X2Qp
9RMC9P5icsg+Kgp8JhtaLyGGFAoL+sKFnYJrc1iZ9Q/zmfQXRLR8aXOiQR839TMAmAP/4gO+Xfgf
a84z6Nq1Ny7ZgQTaE11M3C/fyv6wERm63B6bc5V/T8+OsCisMvO8L1IXT3YyO27XRH/z0JCtfIMf
4zcGo0KEXM/8QzVA2OYNJijq6UcoxfqXhoypTRJimnK0uVZH9z86CHgoGA1vv1emWi6c4YxofR7s
ZSrnHLDQ/e2yWJU2NrRHGgN2a1pcDcaPusmcPnPJJPlkDqfXrE9lbUk5OIdG4gcEycYghtNvoB9y
C6DJ2eRRbyi4TimTuQH+4KfbGelo+2esbzyDfmfzkpME85rkizMcAu976BcjXyVFa8g6/qEZ+V2t
LotrPc3kCNs6LEOdPtt23OoA/7cN40xKPed6S4jI6E33+pLkXz1MmJLIUiYf38eDtAcRzjTdAdI1
oA0j7Aa/+YNCNVB+Fx/TLaE2VOKnodCAxeewN4sang0CFGkC7fATF9fFdJWxJdBzAN8agByP6OD/
GoIWO+2MSSPLTKKGW1MeWkhjmm0ZIhLynsSfsucMbiOVSdsAw/yDwhDvgVLiip894krLmBCVw882
CUrj7sSwUKgISdHvhKoUABXlVIj9bIW0/ocO/lpcqcvFDXy5uvcXT1OrDjp2VUgaJJW8RJ9V7vG0
uR+sBsnrWrdPoCo4MrB8CXYmc4QDHgpcypkkIKG/y0HeUyzH2asuIpqaospK7jQp1Fjcqk6m5t81
kTTPmjrOixc/K5XKUbSLy90/VHrURw7BxHAxkCcg3q4BGeOl6Ebb0vwcUeotZ0C6PnphfFU2Svgy
2fKk4MgPlEgw2RJ7SRXm9jhExfYnXhWamQcbhF6R9nbA/qARq1RhWB9HKo9FI7iQEdZtbabe4Iue
/gRNFxV/grUofoG7aJMvV8P8ZQQUL8DbotulhHgtV+Vb34I1DLiNIhtof8E20WaSIFjgTFfG00o2
0m9AxjpWTEB7u7uIKlKRJ1hPeGczOXwvnbgMOlR1jTdKjtfJKVd/EvALfURDCm1oNOqn6ukFy7ox
68SywPZD2b8+uX0PXr5yXC0y+ike5EXAn0F1TqIYJqB2B3v0fErRX9N97m5ns/wcmV7Xll7ZAuUo
hawdsQHb9XNPWBxG+FufKaFPM9lALOumwPRmcaHwOUAWTGHBir1XO22mJZcDQSd7M1f9BZre2pij
l8DesjsTwgeCwcm0i4eKK8NpdxC5xtwlNdIL5Es79sZ87pt16bSWOsTz5RGeo8z9MwX8AXkD8Vv4
79lwyVw2NALC+sSqhU+J9TEW12RZ06Le7XEjSZYYCNMlJpXNhHeIgxfhcbkEyt+sXXiQDI/1Mx1a
+OyYq4YdoWHlKYbGuR22VvE3SQwNs3O5o5YFePnw96hrOxOSR09TVE2ea3ENqIbTN8Swh/VP0eye
ZH8GRwLsR/kQcclfY1cRWdOfq/k/L13X0yGrprzFvf6iCVrZ1YrgRHXBbQUV9YbYbbjPsO7g9TFb
90TpAhpL9REUilABw2C5qM5WqGMTRW9AlU0nRTqztGxjbumDHI17+UdXDjthFNxT9fDKhmgQIgjF
ZK50EAlxwHEzlmWarpzPrOM0jvb9X0uLt2Qh9PjXJ6XrdO8R6AEccgk4jTtpoC4TMskiepcpknoB
Iunc5GV+AjcVVIMpCxkFIlaC7RbGDLNY16Lxtov0M+v6VqosLr0VDGSTvMFtEC5+lhSOq53KOylg
c4Lj2FUQtV7caXau5V8NV4t6d51B/FPBAjBkUYOAGUTGb52RQ31bRp6q/cOAwhdi8pXRSda/UrT0
gYubjF9oXhvWrwVvit7bRIXLQ/UKsAznV+B9d82Julb9lqB6ZTMjcnTbSwZc4DJM7p7sYDjx21Jb
pJpjVoup4Ga+31zZxSdP4ppXV7XwsJmPijf5gSXqIpPEg75wsS4fMibisb6MWt7tVkuNSYEDQ0hi
o5gPLG7EESwMIXflZfPxBwjU1WFaHCX+O8e8mZOOskS8fMlMMuPkROqNmuvt/Wfm/LPLWWvmnJN9
lgQ+58Hv56bm/8T5Juzc+QUOAuJeQBC9iPZQxR72bfB4tE11hAt5WdSXg6ahxAavhISsECsfRrnZ
7Ed2Ok+n/dYe5LLkYafWFEnpj9f1UrsKP/ifn2Em88HSBdf9DIZEsgaDKre80rLW4WNovSVmAozH
BiPO34+Po4ZKLy0+w6W7vKFq/lvjJM+w7SEaV7tNhMG3aRGPAeyK24M+DsIVOgWEdckzeHlWtszm
X4nJccHg98540IbJFZhgJJQMWRBh0kZPyuEpuh7+LkodMk5mD8MfLndSSPSvVWX46+M+e04ymR5F
3zJ9UdfPXQi9ZLj1h2yozvbuCExNn/SwooBDMMVyNsGwxMG8cxysjVk/aGvBIwI9oNWeQ05oCcDS
8aWwSZwje+QAlljVNNDr8bulIhAKnytFXha5pyXPsbVKdJ25fQwva2KZEzPRbfy8+ddyoyJ6vcxD
/KeOjRFCRiCVJilRU3ResUlqRuvJQSeiyoMy3MPNeawn1t8xiM/xeUty00JgZzCGkZS65AbVPX+i
HPwWUB4GBltoShrs5XnuzkKq6bFlOoAYwaldtaJI1ODW+frwZi0rS8/Ts4ATuDqETTzvswuk4187
zaRGk+HH85ZwZ6aNqXKJDJJ4Zk0/jIBwBUNMwBssjN83mcwB6a8+bzPwscyI/HmgSmb6/r4wynAn
YwxEFOfKtB6BJCcwkpRXcArWezisMhN9ykPUtSM/h9wmbYwxRQ6eUqA4li0psO1ID0VBV7bCF+xT
E8n1VUk6Af2jeSEJmG3uCajlzmIaXLEjYws9JZD79PO0ZFcfBFrUR0mQzOzgqYHFZ8qZBPs0OuLx
y/q4+CMX7tjfJnDQTOUUFPNLaK8xVgtYKmVeSiNmWI0xenA17RSfeQy57brjEaJEGbkAlaCB2JtT
8hZ+V7blh2Q5zVZ/weamLQcpu4bx4lsbGCG47iWuOsa6Bl+WPq023Kuv+PaYdzCp2OhyNAN7J2r+
v6Shbw3GYvTMSEzBk1N5kQuXEK/5EkFMIMde5sG4fVB6hgXaP6atLGYqymWkKT2jpXRHNdYucxob
kdMPLsPkvj2FfxPO2OLDBA8J1w++kSCyoYPaXCI07ufenV5X8ulRsDxunJ3/foq9lmQFixRh0g5N
g+ETOU2/+KW6D+rKg7tbGmVEbsv3sIJp311UF1DEytPHWu7bh77I4aMHZUj3SJRa1Zz3QcGdozVK
0EurrnJ36074rYolPZbL73bylMlMBn/Oz3kc4/qruNhtua8a/8PbvBFiC+kDJRIL0Z/ws4dlZp2x
cNnLA90i9NYzvsQ9rbv7OB8IvtUaH1mEmX9s8jpTTwRw/RudaTOPAxouvJVypWR7L7qt58AdgsfH
JWYV8lSJyLlVc+84MonoXA5fFbRSe/JFJtOXeAbERlhjusbrMeQkoI/8DDAk1dUg4gkSh9PSS9Px
Q+Nfpa1pnrnU8NgBJKF4Q8OPkvAWv90shRT9O3xNkTxYUl6aPfrH6Wen/U/xFEKt33LOAz1SzXug
gtJ+fAiP8hLqdqHDBujGor+OpLdOb4ZiKws7JPYbYgsC7sgoPaSBK32FrQfvkJqrrIRn+x+MiGTS
r99/g1qfrk+LPV8+swadpUE619BM0pRcGEUA8j4b/iagX45kdlUaTKX1QlOzX2PZHoAY6NkaJBwG
i2nLylZfpTUMxMRcdVthC9Zq6oAAr/U1BixHn3AS8mypAd1qv4EdDAEcnxse+LS30cSZ0GqybrsS
7bdShDjcYuetow12+00hdTnhSbH2DMoI1R6xbOF49ESLzHyF3IGGSiMdo2zgAxGjamMh4mC1kgkx
2uZ0DMyt0ubArSraeMtiugBlApaEtmL7Ooln7qHH8tFX2AfMj2LnXELjCANs18+MxhUzsqotQphW
V/xBghuU5xs0UNYbhodoxIyq2udIhv/QEn+rnrqboStcwXU5NkMkgBFY5+HfZ3TQTEjqEoD8KRK1
R/sfsH6ejZhpB4kGr0geL7gCsnE7fkt8Tie9eYHhHzGLAWrC+y9gUHKc1LeqfHveSrI3UpuWYVNj
KQH7/kNNzA85lzsjK8scfGq9BqTEtOwob/tO1i4car2uKjjH0mV1a5ZWznyzaTda7wUN3mMrC3nw
VoPhb2ZsDU24HJ803PmDTXuKqdT0umK0yk4KF1i3vWJbfm7/PkmatugdW+Ww6JRu5882En6f9j/9
NeNcaaBRT+X3J59bqQZuhR4eXilvPoxXrSqAKzL9B3ikvbK8m0c8ffycyoxHqRfRYICuLKPMUI3p
UH3ipdrbu1nhQJq2dJvC/T7EZzxuM4uhhLuGYsveTDzHsIPzz7hGQm+nBR7zyLzrpBRSkThn3EaF
19or5Z+AW+1eD1VfHfjNco9teJVcleVEdjbNDQrgaD8gjMr8BTRmhV7q6ahu2rBy9gwlQwo3c91G
sFHwPYB2loG+pcZMbtRKCn+kQvD7vT/WAHxOASw7BgVtuq4NiCqwCQ4k1A9+h74bpelD8bj2FU5z
dxNGE3lZ+E1JF39AVkzWmKyyNqI+GIq+WCmHjbea0/+Ph7+X64cbd5mKkL0DNwfwnnEIXhi2ZxpP
1vdPq8LlbfQ52PblBhMVfvl+Csq778EtMhSBbYhV1kYk7NhpHFAaaJk7/CWWQnXmYoFTDZygUdi/
GFvUEAVT50HjnnKbN2MnJMQ0crWrNF8+RF5Uw1a2LIvOfKXpUlX1BeIiAyVCoEWc+CDY35nsvpVW
0+DNNhRP6zuzf1qKzRbh8Vw/ofmcNPwojhJSVvctnMEOv2ASr01/g0AUOVpZy5u7SnZKsNonO272
mtc+wxDxKRLnWzJcVmUMI/k8pVUrm28pHK8fxygeycE7fKB1DAnYtghqHdx9eRLmKnAAnXS2y/Q0
XlbtJMSRiq2Mw5rkZV4NYvo0U2FNJkYbTfGx6FZIS2XoG/VzDWYEu+9pHOwqZ8ndEIAHcqjHCw3U
dQTRl7x2KTlKabj7ZNucmeU8HaRK9PoDKQrkNbKie1d63JhUb29g4cXVYIXIuerh+X40Y+ZIJyMO
acuFYzrTduQ3lEIVY6voSM2boC1JkFbmx0rPeKY09EPW95RN7iNfFIuUw9uQURTt4PXFH51HS749
6iZLEcmfMKxaAkrTBucleS4KOZ13YYd8tOmT9QCnF4TfQL3IEp5d/GkstTbB08Ebw5feIAgpA4xG
vZ0P7H4Rns0DVqJ1IZ7TQp7qfYpUf4wDrokijmopZbTHDV6nAxghZWkIcqZ8EJYRZJwisykHFAVa
174+YxDVkbFvGYP4KJVAllStXsfaL49qBJDpVwgPzyCN0Bm7GdDvqLSeFFPuaQoM9LqlhIUbR5oI
gNC9sc+f3n54ACoNXH4eGUnFjhDXCb+Cpj98f2dNzHJ12C88zxBgqCVk065nfpx8ORCpWcNU3gEW
XW678vWnCMOQK9qTs8/bfSuq4nBXlQrYlCTUfb8F2hfcAER9OUvemxi3/Boqr/Pky70O3Y2IcdbA
30Ud2sbOwqimTGpIGr+0d9mkUE2zrFxBKMpm8bpPT6L/VL+OliU9ONtI+CD5fxXR22tZKJB2gdGG
lJ4jN+WIzPXpKRy6XFuTrIvWv7VvPKHWnkl7ZSphBXWzNz9jCiuqfsjPnox/Cj+irsmD4PjwuJ7V
SmTKkae4aba68FbSocZ3WV8cfQrn/G+hTM9TTNrjlzca4Mojx/vYQlvl9TnMh7XeGaBR/G35Xsyx
Tifdg8sTj1zNAHOW6B5i8AbZaGo++79JzpJIDEYI1CbODPnl8P4z5ch0mvB61jSSyGA3gJqiCdcn
TQlIyDFN2/rNedwXgvicbkPruJzNwFLcww4GyOmfA21jr4YR3Dt5PZyoWWnsKSxQEqYPdy+hAYsz
MoyVxXU4TiFvXyuqI/Qz3w9xXp+TCsa9/daAXSfVwy/NeHTREiLFIUmBlIQp0Ubrnl7S1wPhFUwi
bilFVLh1fnWPyi3GUbDwqxK/6wNFcaYnb9a19tJxc3MFPGt6fBUk81QvhliuF8FLZDNnnYd40S3P
T4RmwRBYKFHwv6f6uiCnK9eHEAWM/Ofl92EyigPnkUifpC2WLOK2Y0NrY476OjyWPsUWzplXrgBN
XmlsK1j2dowd/uvXha2HhS8uCf1R97Bipm/ocE6I1mBpwZF9OfuqJfgoqrAxJAN3Ln3hz7HK704I
z+zIKiBDG79iJZ5NOcqRbdbgvVownPeHt5Ekf588cRUd3CRbtHcBcw8cZXSx8f0cDUk4pnjE6cQD
sJ3IHVz6tdCwB+KtxbtfQlI309ZhzVTZSjB5AMmWEXQgv4BUzxkVo6I6OyUnFlIpwliwIDDvbyYy
pa4t9jK9f+myr/V2xi2ldW7Eqs7xSiH4GZELrZ9th8ZDFpPttyt9YXgpQTu/VECUSuHLvT1dExT7
apUyp/FsVu0wYvjlvS+uRIhZXozU1B76JSTJo1XPd6n19IBIN1wJSl9fjdB16vJhBdO8Y6AL7rOx
+t8ReT8Ek4ugNnK1gq6/D5CjSUIsOsp8vnPaXMcKJ9Z13G78D65DIkYJTkOzp42sDOs2noxJj6uq
qFPcTwKJ7euILisnWkR6lzFI+jOOkrxEv+LcVtGrFE72leCu2V9bj3ow55/OwTK/t5GlR9BCEoM9
e6N80aRF593vutbSY8IXqzJlduKKRGQ6bgHMsNR0wXnDe4gSIer9jcJ1DWNjej867i1PcfPyv0h+
qHZ3I+VvYGfo7sveT+TqGwbHDmf7sWjYSO9x0NvWUvAbbwjprjzciIdofwapDJs+kMxtYoZfGp8o
PIK8SIgFF3DpCYtlwbP/SPI+L5KxKr7FeTnm5iXPiFbvqFSmaQLXbooCyW0Vu5zpYIq7I9Aeii4B
gzadkG11W9egaZHWxuhtJXKaqroeBqu8lIjgCFYvQvLR5g5GqjHkFfhahPtgIgCgPVPcwbbwn+pn
VPvRPNOb0Z7fBL76a9/uBOJYZT6A02tCx8HqNJ5Kt3rLR7uIRPb8HpfHkO/XkDsUFBWIzTOBvFT0
fQMGfP49H8wm18XWUSqwkIKFMj56wEGmbUAQ2IpiP1ME62/byTVYfff+gZDG3xNCdnwMI0kJ6y4X
dy7LvQLLX3EQGJVTO2xlHaz7AK/2FjV0rec2M6Pf6Zgk2avFTyk09d08zSGpVqs8jY3kxcwK7lW2
K4VbcisXXbEeCrm6TpnfaMOOTzRA6e1DubcGw47D0aPX8CcYsSjg1V37bGnLf1o5n2FCk6J3V782
PT1LrXncqBZjx5mf6pOGoN/OHV3fYbfpfP7dDVMnjbBP7tXZPlVJPqlq+mQcOo6siXjcdshiqjOr
zdHXfioFQe9tqpgeDWBi8aUaX67uA2cyrkdkIKDjWY8c7TQ0/+8OnoKrSIrpd8Way6yeHxXgXaPR
mVSQsvT6GxuBFsB5UMoF+nKZfzzBkDqLtFK844Ksh1FfdZ9S0TROp5EX1G8QXtuWnTObL+kDipMH
lsMsz66FG+TOSjx3m3DPbPgwBy9ZQ8Qz1ZI1aYCAduNlbEl5RsW1p7rsnj5GxesJwkRN2ywhjkec
c9j3vF0USViFJu+y7rJaKCqOPLtb0oMXd/q/9Gu/MBvpusHtOcQNeu8iR0aVdmn/TkeTHvLIvBnG
+YJiNMas7KveNhxAsSuXnegnN03taB41Yt9455E/+VjzAKe+bc90R4sFCs1ha2WDeyRc+qxXPp5K
b8GzWsdZ+EGpUMjpwLcdDxlgPob+FZchOdeLLOHR57LOq4k3J6XWQjUJC5AlNznqgd6Cjuivwp9P
hLBoSlBXriquo3anYJef3k+mCSUiGjXK4mGfGZdg1mK1ldBvG8780KdWxbJBAGLNtSxTKsnBWYbG
ob9k1+eXKYcyBpVizWgYNo4XEwSYlHs/oUu2Or1h9/3gtSgZ+ymVvsTCV0c+uyPtKjaFvaNdc8se
GjUvlY3fPl9nInBY+3V9TGe57LcaMPrYhvm6D+kxIjMNXJhfJJdLR22oyeMkhU2CVub/9HA8JIwm
syRks/K759xyLVe2KU0YqI3eXJlyL9VtUoODQ2jugGVvpu3+EIltFHqF//LI1MBcR3phg/DMXhkj
34CGTXQngAt6fD0vHeC1W174NUj8lM9RMqlxHGGEZUh48M/WZFOp9Qvc3gop+iqKYXI/w85I5YuI
rhfwdHHXjEbN3igPLrKjrH07ZRvYw1Ky47aLHhmuCaBO3hDiJcsfJqYgSSsqmrT1/pt/ZsTzM26a
vtfEZAoj6QvdQox5mUFHZ82aRx4LC8amPVGnxgSSG7VDl17GGbQ/BD5cMYup02u0DF1IaO2+SCWU
nYOYTg3Cufcj7IGwz22PVVwEYEx+Tez1TKkq09swNnWDbFWEK6Eg/geeJsmwQPoa7gE/gySLYkZS
28lrCWoHRy8eIv5sUoS75xqzYUVzOt+43OJu6WqJLzgmQZfBD65H7mVdvyScQGlC8odBS0FgcS7/
IueuQCq1S8xvqCez9J2AAYZsfOAv7159priLXLwoTuUtt+hsiJjhMrQ0O8rhKOh4ZJDc1GfYLoOJ
c+uK8MOC2UUUgAQ0r8JTWkjzjGuVJX7ynyFH/j0VWL2cyJaPM0/Z40R88TYv2Cu3Wv3PktalBxh0
FdMRvbEGUWx3ifyFhCeJEoKvoA24RIYgKRfLwfH+17Qwh2uZ2MZQhK59LbA/6EmTNu2GWkYB97DN
iMznoXFZksGhwy1sgzxuNKRjhaQXrer33oUFZeQoe2cY+NcJaUFGfNvtTMDDXYbs11KLBOUXrBfp
mCt2V9gAfhoJz/FDLMpXqU0hyuoKPp1diGNTw7s9NPO88fuCbOsi3guGWgPFzNTzUOd8kvwSFdUQ
adVdCPAy9g5QXgCSG+nIHUHxv3DGAdDCJGrK6tduh55XxTZMBXlwBj587PVaAnGxRvJxirBhlUU1
oyZ55WQjc9zuMArFSE/19v6C6e0ADGFpWaDLFfKiRLUTxtt0kq6BM2vkOC9FcLm2YcaPo/2+tgKI
knX5BF95MOM8uyMy3J7P29yqXm+W/IoWoHGGqPiLW2SxUwuD1FSGMxYMdCMg3aIkfdv17cKFSiv2
JRfTMfO5BFWEYCfBx3ubXhVW/q7nj6AL0rwuXkcQHjcg7gLul8YVcDVIdx8RqtUBgrh/u+wSCQDx
2TBzsFQwT8X42Fqluj7rJxPnkBQqmArM7phXD69603GKsko9CR54oqxd49uZsW1Cgup0ZAT1DzXE
rGVsWlBLg3sx2aPr6c9Vrd7qjI7UgTGR8IX9adLUNS+5n0rV/Zu7wLmB8Qgw0qN+haEZ4uMrtewr
D6Uvz9usmldmifiodyre4N1tSyXAWe+43MBaosnceRF+LFz6Yu/IWRaf+RTyObevvDbLDH+pc7wu
YdYXAVrjqs+XNO6xN0DtC2jBHCAiWrEytl6kQ4w21KzaUOH36OKNZTzCN4BbtYDP7u13xfTI51Qr
jnCjEyhiXREQtFZDT5cPZfZ5hvyuNS99qaVl6TrSj2X1d9N4voonKsGcXDYC993MWTSs5jZrME6y
i9BVvjZ4ixF5pH767K0y8T7Mo254y9Q9RxvMQnN3yPzh/3CLLAYV+7OaerqqcPqeZv2BHOO8Omqs
H0VwiuJSQJ5rNp0ZBWoobKJ+3pwKKhOWFpt0MZwsA0jTiBsolwVWP20JmzNG4qnemv371CQZandZ
Ip5owLpOQixHdJirAN0YCzDQ4h/7wqSfwqy1GTA7p5dnYIIsFWpFnEcY/wfSQEwzhpTJ/tZvll7N
AEW13s2vbXdCegTeSO6AEmlVeGLOX9b5P8R8DpptbRdx6vqi2ukAgSVOrW70IGNjwt2I8Nlgnn6Y
EpFlGYQ2JBA0YZKy3iBumhCdYLvq/wghT/KsPNZVr5BZUwFlM9TFekUvOtaEfXYuIQ3CnKat2Z/J
9XoFPy52Rd9rRmiro39SpKNdOBzA0ug6IS/VNj87J1duJ2QsaiGZ7bs1O3F+tD+rXdyupqfSviRp
TSsfrZX71vi2zlfw7IBJ8t6NVGvcJoe3OVRdTBVSbI7taiAu3w1gnjwq1NVMjxYL6uFO22tITgks
tn8idSuJPUaMZNqXx6riEg3fOdC9LS5lvvWSaGFmfjKfYKRGMz5oGvmQx6tlCSi2+/BCSv93Cyj0
LSGmH1rQFX4x7+QZSTpY1kAGh2mqRW73H3qcSTPaN4E/7/aAPFWCNRlRiLM3YwvUpmyOVjzIE/fy
vHY4TeSB8Ly6TemofCaN339rvWLejM9z7io474P7wY5yHv9HyEcHkZLELZFJTwrpUWyckFlN5/5z
nuRifV1BGr6eyBsfDmAROlnKHk7FcIRIpbcCkrHQPjmbB4RElD8Eg2es50FHKqjueJUL1g6plzqR
+qC/6pft7nvshmMhkrTc8ZFBKpG70HE5KAKYDvMXH4V8QZsC9tLdySkOPuVAq4pThkqs1LPAZquR
M7QnYqGKH92xTfMlpRxlrfL5Zdjm3rSVhw3XEG5+80o1aqx8SpOw/KdRdFTUQFXxGdFY6gqlpYpx
Tq35+WDgvXIXgDi6g98cRbgvooogey6z2xUnnA91z72FhXkJmWJaZn7Js2DtTTU5siFRdRPtTI4w
NwzBFq1XqUoPybZ/JP8rXMPPu76rIIBdjsCJt1KRO1llhGpuwKiUTZ4zPlBy/sD/anAusMxHloFS
ZkAbyC+VRO1nwRlUq/MbPaoSlGPpF3vLKBJ/TiRPTvk4BiPB+vO9lXJnET0dN6O34NVoXLjgH11z
4I6ST7QcSxSDVoDinToU/eWXaeGGOlgp/H3PQj9pd98q5DE7ZsZg15WWg42ur0wdesvUNPuccOZo
BlDJZ/oWPIYbeRWSqyXwG3PzWJyd1Lwn7L9KJBQazsGfjiE14j3AlV3IG5muMTxCc2J1zWrT3elZ
ABFTQVYmaGOZ5dV33GcxdXuVIlcCRveorYZhvK6wVsoNt5+z3qXKLnCo23RpVtBBaxkDDC0SFwfL
bA/vkZJG8MyUV8X5Ij12y7QUWlhDzxa7rmF9NuDtam8JRYJFutB7dtZH01WxeLoZ6ndQmtz+A3G8
xbVPprx4Z8sOZNFEI96NCBBYRmKoTkAKBQZo9VvNFdlBr+8j6QdiePSa41h6dQdR6GKxLW55INx5
rNhxSi29UnyrxAreGrCGo+o6enZRPoL/m/6X7yPeN75E/eFHNDxVzfSvq5q3LSJK0PuC5R4WEyXw
+cTDti5T09ZnMR/KQLKXZ+gQyXvPZPIbmd7/6Dfy2+0CQsvWfgsu9QrzXH3pntsP9xUVEDufHMzR
S1Kcox0YF2uHqojC5AxDKUmK7me+SQUgCk69g6k4StAJeTr04YvVsl9fUoI4TeEDWlenkv+YPCHd
XUw+ys+zUS13j6bZIbuu1AGqEA/kDL9df+YDgW7VT4TuA6pjsuLFYMaTu7QxllnjnYGrP4+pvXj+
ABtGpCpYU1rgmyeMW7X5jX2/zeNL8cYmkJ7fOAFx4O41tRSLJB+4ZUI4En9LMb2VqZrpqGyKdArb
6W1IqINPPSuL7zJpm9MN/ThoUFdpDv+Z3rS7Nfk6338Yn5nzRFEvNKD2KL/Pktkcnz11BzbZHJyi
RPPdmUccM6piQgB1727VziK1hQyfX9PFbK9HZMB/zYN9FBbtKsN/TwshS6lS/Ii8lrLmJFRLhKsz
i+jzURDM8rB2slYVuELeTAI2S/YmLBOAXXwMffL0pfRLThXsD7HqlpSJQRTpOmn05QNX86tL81u8
tO+/e+Q1L7woxNk1JXZxCeoyfHTwG22zD5S0aFlI6cY42zTKHF0D9bV8pkLaMgB8AtHQCGj9U8jj
6EqyLq74APZoHM4KXXzWG3CqDc8ErHT+qmayJQCDZUw5N7Y5elGv8dr+7rhnu7CEhpkwtJ5MHVP8
O4Ur3aEf4hTH1vo41/mPAi0p2b56oPLi3zIJDOLEvSwZL2YI114/Oa3Nw6cBJe51o9lJOuClj5Q6
iv7JBJLrFtJX9G/BIbJ9P3kXmySo5VFxgBtehOCnzmqlBC+Mmylt8cxxjjkv29laHr+9NIQGVPdG
wGB7LBDt0vaIXsfHZPY8Ms+H+oZC6xHY+HvRbfzWsT+pIkVTIS7R4cfyb1yyQ8Qawm6dzqAvmzwj
gqqSz6dQuYV3f1ZE/wFiGUQIARH1TexgVpkC0oghN6mi+0LTBet574JBpdjIP7+4jTa0fthfAl6x
IsMZe50eVrvx4JTc4YylcYWXzEc8nJWSlQBBZUMOyjR0WdQTEsgUJXDBkuPzfHfb8+w86Occ2RHj
ZNlqX1F8h41554vjXriMOCCNM/3kWTtYOh3N4iayXopzIQRLv49E280yJOVYK/w76gidqNi/oiS0
hKhlWgOZGnqGkIE25/wvhmJ8w91sh2Q/XBtv9fzMNv4wnXs+B7ZoT1kUAMDuMqa3V4WFDrcDRiw7
U6oEXzlkOgP9CQpKYHJ+0f0ncYqCvWKXTHcloQ/jz30NBdSFRXUUQ8UNIJE7TIOhuuundMeQpURs
ZvbN+FI9kz5/qwo8YqZ7BPQI/ylZXZF/GdXKY1NB6apwXc/VQP71TzTSQweWALoy+YBtC7YVAhg3
jh6XmKoYmwvgK4g/RheIZ0uPFKZa8oZchlB/lnw20BBYupvynvtHCZcF0mJ2F+6WGqJX/vEYBZmb
OA0cyT5WhPylYbmGBUz/JitX/9emltd0QQrjE+H0qktRsGFpPLMt6XGVuNyF3iz0Cj5nCK2tqpNs
8Oo8WPI/GdGbAyJyW3z70Ovddrs9K1awoclufWB4YzdxcX4+sxi09C+nrHcNyya47s20EgTHtzRw
6vqWJqRisC3lrizmNUSVzJEsODhC+S861fmG05Ae3wHhja56XHv4FlVcmav2KXYwW216GeYNk+vf
bYTZ0vfqSkjc2LzYYAfzj0Lqwiplrza0muwqfWFpdkvxaSlEghIOOZ5WCnusWxPd5o0TQ5leVSyJ
UetryPkA1dTBStxOdoHK0ouwoHfudJi8mO9NFea+rUleokoGAUFmVv1phNwY517aMFwaR6L/TPyu
nlkfdlwpgVqxYfd1tll9L34UELvvyWVqjMZbGbytfysDAxKbUWghi5ZejEdeBD7tApGnvuKEWHVI
AESo3/0c9hmmdwboNd2jnJq6z2KlqWcTYMdTGh5bbqduzvPVA+BhGoTsnzz2gBAGv7teBH55v1hO
KtdCz6wee6D1NWx++Ga5ERmVxAYOzK9QqWLUmG8TO1HT2t/xRunyk9KI4K0WHTeUZBlhJvcncMA/
AOSHyuJ/n/lJnveaWIZOneseoppbHGCLC3mpjKelmuJXo+sqN2efPrhZnaDdptDfuCzetQYtoiDz
T32Eu/2Qj5tc90MmyPKBACnK1hXmr0c5F6HQOBBdJ2TMLMvbwQbIjWcYpDVo5jOa7b/es6+OSgtJ
eD/T+caJJ62g3J9TNXKY9xG09hNKozHpcaRzGa/qsnE7IilPcOL0BIEat304GBuRvBwcWtk5vjuG
UocljnAUDr1eM2wFNzTSAEt2W7ilHw5jLKPHRJAyDZqww/EEQCdjuaWp+OtSXQmYxbJa1XdabyjE
EGYjjpL1Wg5JvaaN9CPJfexxlqulYAHAIvUKwHpgihmTKBH6I0570BAehRWNX8EG3WAxLWQx9cv0
i2hxcnjXtTnNStMQ2bcIXOiIsMvhTlpVo7TEKzZrsVAhFc9ro7qVvJn7Bt+62Lb9Ryq3Jb0nq+Ul
d0/JmOJZ58Iy/Cg0xidemhrP+xon/7JpoetwE5NjXBxAmbjh0GDw8UKJywy0S71BmJX4LJgVR7uy
zXiKd5K5VV0hQ2HgNdyzTcFOlswcwinDW8QgdmkWe2Py0mdBcv0tSQkTp4dD/BXHsfuAPZH0y5Jl
lpM7w/MMzP5wvwIMOOjcpzzX+9kLuqFbkFvRaM9b02R0PsuA9pZ0pyQKvzGRnhOK2o9oEgODvXzJ
vCK8jGwIP9qDcrG3pRSool6+9dbgBtkqID88ntxa/PUHPfb4jxHR4hhSIz2M1s7551cd/xvbwOUB
E3+nIzs0Pxjb5Nwi+/PwooGa5zTnWyQfHZNpCJmVlXK/Mz4x0BNb84ukdsX3djodnmjIONPMBBTj
k2Yv1BiKCCMgl3cRUZVHXPXANgVD2cb+Ci5cUVyqY10MNyKWj7KRJisY/IMKZ5uJdQv5duHyxqp9
EOEC6tKkN5qAG4gxOBMRE3kRbLnxWZumy/Ui8iGTrcGbodgp4alt7+xqH7iJ+8me5HRnMUUr68lc
YnSDAjJul8h6Ku1Xksu86NGwspz0KrBHSFrbg+KUk4Rh40Lr2xFr7tU+FAACUpmi7Wl4Q315KQAC
kax7q6robNeYhjahhWK0W619xLH59C9sWEaFPfW+TbrI3rnQqdYXizrTqN0tJsjkoeW50RzZisO2
gmz1Ka5o0ZcXJ8SX9Ag6MmtT0XbzFpG5BlIY4zyLJOM07N7T0WUpRqMqh1QUXLAdxKLe+oeSLMOG
UYcnhLL6r+2qo6TNkmp0kOA1xQUyYzsnd3ZrYO5gmjqCX64+3RVp+k4Wct68jjz3GPXI7uPUfI2T
x3IxDfwWXWbq9Cvz+TBFc3P8SEw7FcQtcA3lkvZNL6xvFIboIM2zDQqpNl7/qWMqdIwD8Rb6KsgH
XNZ0FdLRvMj3nJhtwjVSLZictHYtEi1k2hOhELpBujUiKVYem5jAaACW1bBFw+/xlUYui9JMu2u8
mrOeZijxdDTJyP9vpVbHwW+bTZh3wBJto2SHp6sFcJ+S6sGx9y9kGcPrelaz3H+lGAzuWRS9r597
aZqEHOLk93YsZMQY0GM0nbLqb9vy5IxjcyX7sUkBCDmHFvZs3FEyiVOz93gF9ljv2Sp6zc5ZW2NG
uBgE8JjO/93shXSNfukSBBLzzuqN8T0/L2cm4OsSK7+YzfGHeaH0pCZ6eyhI628EbufkiETtILlU
6Os8vOCGsMOBsuijh/+yZiVDWt8hkraw/+tZyQVLoHvju/se489/BjmndbP+QF/Jy9mswqa48wMe
3QPG2mhW7njehER4qZB+FZFxSa3YsnHiHIZO6VNWEMDplyzDqhLdJojHwaleyC3zXXOjv4vEBcN/
eIXP55s7Uw1NgGDrz1uMpcAGRlCP4T60+/q/4+DCVVDylEcSVCYcxQOkwZXaBrBV9238HCdJx5Vj
CizQbc5H0fuv+Xm38a9Y0J891Mk2EQ9hOsNnNQ+wctiQfwVDDCuaaKQK5MYCMZDqFQnF0g2QmdTY
cooOKuQJdVJY1yZRhBHZmmd0o5v/sK85OF6/yck3TCrmzxLtUiXEqfO8pemPZuI51yxGqyjQr1dg
8xW2NFNkqrurLdWzjHEqAuSnuJY5n/GqkuHPif0gHaeA+2u4HSOwVlSPaPI12LvKXA6+ogF10UhT
nsJgPrKfKon+hEZ6LbN21X73xSzupBr2+lUGnmReTuIgNg4RIGaYZmJjtRdJg9BivvFlz8xl+KSW
RAjQmCR4wUTrWcXMFhPUBBWTHLm9wCp6VSYIynvq4FJ/w0akrnnhT7oSV1uQAwbGV8jNIc3OBai8
uslsE7Ph5wt5uWCq/Hd9cjRj6KujwxVutKfvyr0wFUf7h38Hvb17U2WoQNYhSisUi/SUfA8oqpR+
y5l1VvLU4qboWWrDQ9gjB0fARkr8X16MkJYH2re/8VG+Bh81Jzw6PJNE6vCUQYheDoknayXK4/qn
TVtbqpDb/axY6j4wlQWbPrgpfkhDblNNlNgQDs/U4C9080YCVlTK7mGmQhv1h/VGB+9lPjxm+oPD
LEwPAr4yjq/9h8sNOLo10F3NqpG2HnZhxloJnROE+Zoji8oZE50wcYYLRkJOzr9o7muJRU/OkVNs
HvPHvqx7SU4h12W+UX5lNxIc/oxApnf1FpatD/jPhvGsUFKn+e2leS8QxTpLtE6S6Bq124DiXgU7
YVMDXyqDFpF6zU1MN65ZqgSEcwrOf0yaER96YKJa88mp9NECelY4+aCQkYWWJFM0zPfc0GMkiayE
2KRfD6QoR3uydM0MUIqs3NFQh6uEHhwbRn1W79IY4pSMJ7UFVVjbyamCpx0ArMs7Fnl7BNxO1Z2x
Yrg31VY2MT8Pggc0XvB1b84SzKZc+JR8OwS3Kujk+ooNChgmiZrGbXxmTMBp7E307i/Ph88Hg93k
w8oM6aIRg3robhgCBcnwcp3r81iNUMzURRAMzJyM779r7rlawpSIWF97JWp1T7Rwue21jSZHrIal
BTNeiuxGwjI72iYCKqFt7hAL1Gby/28PxCjshIodO9MoJoDLYkt8IVXzOuI29PzArOC3Nvl+ObRF
GH/E/gKEPOs0moxsmLszoK27QVzIAft0eb4r5eUOuv5DNCeFycr05w1oVR2M44GZ59g8aXQ7W8yo
TrQ+Ls3pRaQaCpElQxj2jtlDsi2iz3BCCbvnT1++CzyXVpCk21wf6qdkLTRiyV+AFz4rrEsHASFj
m416vpBybeib3SRIwNtiq6abTuke9Ruh2DZzXPkV3OZEIn8PqZUch+6nCMSgawsEPMJCowd+U2eA
637CeIMrEkpLX+/ZnOW3HP7MMAOAU5b+gdVTdmaPcK+weDo9xujOWWrKJ3svz7A1yO/ZEpQ9vsF/
3UxlSNKQ7UPCSCZX7hUs/nlLt9zzdFD2VPPnKqCWg5J2f0b3k2veVnvtiu7IkxP5rz1uxDuAqm//
kOIMw/MFIi7iaBnNdc8gr4Grjsjm6LrmzdWQqw/nqj1ACr1iimeqN5IaYeLMWrobhE0bRwJbx/bE
urRkzf40N3TSvHYdi/xk98OM+0LtTArXxP6roJ3oIUsMPgigLl0X4d37vzZ1stysOIww5PlTaVBx
RsudFSYmNjQ695OE3uPhWBHQg2NprBjT2LxzdoTtlK3SXDmIIpfUj4x5g9VCgV/8OQbMy96Bg1i8
4wcdgxb47+Nmm9ZtlKsxBCOGUIar1mr1AVCKnbC6trwgOGyBrGnsXdS+rDWYl0www85r7Y5NXlyY
4gbcVVFYPQ4wInLWMLb8KqMMWxP23daVT8iWcebRnK1b9krmB1NK4Q2NNoRvhfMEY2f0J7qRNN9w
KXJomPAEHn4WdlN43a1y73aRc98axBXw9xGKis/fiovH3dXur6AYUF7dorrdWNAbxCqus+wD69dd
AgCsuBm3/1jD95et7bWPD3tvkVxlCUhmuyL24ta4WnOC9hi9xnrDicw5ul4dK/FbW/1u+rtdKVlp
MVjZxp1V/+iCrp7b/fYw6BFSr0jfsxMMZgOGG6+uoxl3efUcZTYalLhuoEprX29Lce8V5nTFjaDo
GnQpaTGXE+vqUjuFdjVPwkQDSH6i/SXteppFd350aVX8QNXCQ3VL7tK/txcTP1QM7uaBa+xT7ae6
BxvOdQjPn7He+5WasPgwHwiTYkmlSAkgxPzKEK6PGH47Zd+NSy+BpHyGg8wHXnaals9OfcQzxd87
78DfKF+0fx0Ayt6wjowjO9DgA2pkK3gH+e7cGXGt1+yExf5HXYtFTbGPa1+AyhvxdILLiidf/Js8
4kq+YOOpi9X+IQDeIAayoturrkFAkq7TALbcxUuGCIMoR3gKV1snLI7ncnU+ys4Vg8Mj44ThHVpM
06iYNvbSZRlnNmA//1FgStiB0o2ZE0Gb6svSStz5dJ4umNlxT4r6hJOMtKJRWtsEXUSuYL3Ot4uh
42AMIDeI744JRQUknEbDIVmxcdHuIz91XVkrR7Twl1gadPFX6XI6RH9I9i/OSkh6peG79VBqNvjq
yePOrb+komh05bFemF8v1TCnASxI1XsoqlESp6LLVstAln0SH7tDyaBWanWwjTltC5nEAaBr2NNR
S3T+cK/IDUdyV9h9GPhk5MpEDfydiXFsN8tWkUAmURyRWPQZSkqNw2Q5PPNqy3Mj8G/RQASG8RRC
BHcux2WhAuVRPds6RiR7fZ9pg+M4BJ8NDrfv794gpvgC6QNspFb9nF6zcIb3sY6ocGX34NQ78Ach
6ceWcgKTPOiBIniFl1TjiLN41QFeQHXUzP2QtCCNSdG60m+TTDDp19DR2MApBdSb9hKspRLYSamc
a69eEHn8diR+TcPb2FbKzbNKX8COJN0fPoVjGZbsvdnYH5U8q8EqWSVfQU5gBofVk2wFA1+d19nD
oScRE88Fy8lYCyaHiWWfM+EnEqvfdEdeYe2Eac6VDYyGBAbdupVTactji7W31lKvJthb0dz5+96g
qXR8HsFzLOGnYBbmMDU9OfEeFQqh1/eiHbJM4oknyFQH6naVtIFTwwcJEcAoIyds3NXmT6g85W+o
RnXibFHtrlJjNA8sYww419uswCUCsji26LqBkUSfVc2OXQBOaLd8Z+jOxfa2/otjL8xJ0TcLBNSQ
UMcCx+YBo0/Kp5HTH1P6mHBdvdAdBmH6JAWT+J8dlPn89GOLWKNYNITf5hyAEBeZ9hpAMSllcoyh
+f8AurhlXAqJQ2xglNPx0b82XR8UZam5BEFNcJPqaFWBltrM7H+I7wJGFuTgEwJ2bcDAebUT1JO1
ev8x7fQy/If24rQC2AjWxp3Sz3gEnRy0oL74JNZnGXOR4JHwEi+LmfNF/tv09oW8brqLN0vWFjm7
JfrZR7D6CoXEhwi2pQj7MkHmx2xR2R3X/ig3FhlHDozD1NRhbKDnai1NAGZzwagOV41/GkQmirlr
8+u/5LHNTudBJLvY+iDVC1ZDudfN9/VdnzDEncWuYx4Yt1CskIb4FbS52LJMSmXCAJt6hb3Ofprr
dyF3iKIMpozACMYpz8DgkwmNgXOIXdIRRbhcUXhC24k/Enr5cUx1gaYCg0jtl+FCJSPLYHJQQwMM
4DmulTEkjjVQVcOGR1L4Rhzou4+10G9BX3LQpe1iebLL7yYqaJZZ6P5G/uPTvohDpNzkqThoNGP8
YM5889p+RQinN7igoCfgtG1up9IXEi1hdRlmTQ8rjmqxVS/iuB8C2JM/yH6Vf1aFYc2r7ixCuv4I
RYx+G2Zzr0afELRe6ejXPmyo3KnvUhRGhV6JhNylFrDdFlCD9ymSTHuTZYr5OfEeTm8FEA2H9m+U
MPgQyI6tlsDutqjt2Z40UQrrzySApfv/kUKy72TtxjRET222kTkGFEFNeAwsjtwpDEm+tqW7yjSG
7aNy/MxsWqSs1Y8pac6GzIAYTXsJW8guHgYEMBeRdUngTWRh18SLqh84QoG27lQa6cTwAJcKJmBA
FshbUs0S1qfKgI6Wx6lWh1cmA4CtBGtLqgQE9oAgbRSvKnYeWjAYGPtSh3kkI7eWtsRB1topAXvu
s/9E7mjUk2ab80pqDPTEMejh/lXpnwlW2lIBuHQCz5bX5YvHH6Qcn7Gq2EA/JzC+upzLZ15aNX5q
eA4zET9MF8WcwFBksY7GBpX3TJy2Wk9H6uU6SW6eNOZOKXVdazHwBsn5aq0xafabD/MAoK3ibVtp
7o0VfDs7roV5EBvTNhVo7kWOl1qlLv4tdVJHcgDoZ78ULT61Es5B6vC6mtMmXT4UiXdQrglRg4dl
xsYu4YS4qGjca/O/KMocjmsOsb6ULXLx+f8qELvjpp9Wnr6x5qZb0WPMr7ewH98FQCvp9Gnj2Ux2
1N4uAmEKsOnG48pH7WHKtvjgVFBrl+nUqLSXrBQNnEpzGk2cmROtRZlXt1STMig0BbR6FZAeqIYi
3tp8N/b/dgLE7ou+EXe6Y++D4t+hrJObu8TduPnBRITQtS56/mxNVp+GbrXlEIGyA37vkMsPvZxz
AQ9VdEf+2sHduaMo36ua2+50tAxcg40S88AfOP+cBnwUqTAUI3d+ZR2R+mEz+fvQ46TgKkmMx4Q3
OGzGk4PqMBsCgtviQfkJXbylZOaN/dYVDIr7fk5Bl96k7W+9yT8EUDfk57CkT2uk1xGmWW1wMQct
5NxMrBu+eIgTXXY8QFHsngqDbXrl9H41U856/gqci5bvlqGKNXembZDlgShFscGhAGWfp0w4wGJG
WBQ8gCtLpVWYRUrqZzYTCxQolUh2P/pDzad4f6NlbzGhDGRUWM+WxyTFoBDC0f/fSS3ySOXdiMlq
eCuP5swwJwhaXVw399C0A5hQIfYGGxILdlIOB9PLv0khI2mHhp3rP/pPGFIUufhb8otUw5+Gk7ZI
yF3LY48vRVl1NSlq8a0PByodpEWYWkcoviABklr4ii5hH3bMG+G5jsTU/GV36u1O+z9ddCUCwKYz
tFZBUjiaD1HwhfMRcOOFUcIA18zDv3VKfmBG54McGGTWoE4MaVlg7lRf/jvU19mpl/Kcd14UgBmF
wQ4/vkQDbaPIBAOmmCkVMhEqcm2jf6/ujCrxCSrNyd/ko5eXrrqANGXWnede6P/R5LFVa0rngcRI
bVSfXnLbw7zAgkv+b4R7fuy1mlYouGDyl86Wv0okkhZ+OXMrESUbZ2JNlYSnnEI4v9cnFJJwJ8nn
Fr8Xkably4kXTwzmHQtZu9DYf8DqVwpaT0Rs1iLSovvfLaZvtJsApdODLLZxZCKRRh1LRdP5LEDy
W23AgNvRPC4T9Mwjj3AwnIKPbf/2UiW0q3t/03HOvKaSIPVh+Ms7bdWZoF8WvMcJq0RBfAMpfOH0
MeI+5/NJXHf/SAIO+jo5aEjJz0ZMHvPF5RK/jv6RGupvoekJfA6ZUN+vSHzXgaTN6ghLGOjg32YV
2TmIExJtSshHXQAi9/cn/jOkjjSL7Mb3sC1qrFHIZfFh4imdYNzEurbkf6g1HG+ZsSfTLFdRf4Hf
I4tfD6bLz/1bz0VI/LlLetSkb4qC2kUH+ri0pMH4Yss/FbeXlO46bZZw6r/WR3ILaDI32JzTvpG6
a7pxTVLvsZxE5HFUxiL9vnHgc9xww/Kd8FF8QUEk36jevAsy33rKMUn2kCXRMeNO0o2Eh3dlIttS
DyzleM7nSCuZ3iI1o0ior1AZMURDYpAPKvxs4xUmVNwGzb34afIatSc94e1OHy7iDrsIUdOMtDFy
QzBpPyhwWN45uDqV2JoCjFg8ikrt14219MNQjkiFRgwcbizMcX85JDRbMAyNXiRAbmsN8BhY8WYh
LJur0nmQzDG4bruKixiDanWeAgieg3meCp5v2aHeMOpyrsF/4TMoIjtElG9EygMVxWLD4Q7EdIPh
wOHEUtAZLDCOL4FWtYPU+2ywfUIJBjBiJmLKavsgjL1QNy2osdV0OY4eOIKS1NYUWi2HbcvVz5/a
WBgAJ7k5v1rSRdx6zmpu+in100lykmp8r1evAKJqw+yrCzkQfngs6tHKS1aot4bNBD7Nn7JdUCCP
lzylNUxUeCFJC54xtnsNn4mYl4KZaPycR7c3V7LOsxhODVFE5zd+RqO2K67b30EiAiDaqNr8v9li
vef9G3nB4X88VBsvkyWBm5v7PoVIInhmp5w8rQ8HboxtJHC4wHnZohHct7UCDhL8lnI+I8Ij7Iq+
Z4P0u8KL10bS+dC4w+pCr5wRbfRDsEBee2fLY1Pp4VF77L8D23Ufwat8urkuT0ukEH06lklLgNo5
rggKOe33Fyu+cmTmIPs9LPw8J1YTh1+kQsciJ7KVMhHl11nRtbKvkQT6d8Y+Uiz3mM5k7lqMQ1Aa
nx2xdioUHdfnE0paQQPjcrwIccKUZCLPeb/9131ESo7SSy9KazEr9L8l3F/3+3qXMKVeU6fZnS/+
tT6hS8iI9gn3dLdBW7/FP0P64Y+LdB/wV8CexdHNhEs6jaCe9tDnLuUoQDsN2x4q2eZ2igtlYwGN
OihJQXikYLrQIRaVLvMyEjZBRDsBJXMLlM0iW9yOfb981rNT3CZXXV7h9L3cd3/W0dIaFclfkZtd
fWBQhoW6cQMGK2hyy0aFv9hzyzcdbhvVIm7Dc+d7Q4WRQxMONwF7WAJ/jNric/Wr/dpQdJ7vfYpm
0q4Ou71PIl8DZNQHPRdIBYVNjA7ISlENmP2Ke+HFn7WduOEYYBNDCFqsJTGgB5uAL3kkkeHelI1B
zZXCuw4xGuRRbZBpwoQ06NFfERTFbZyRB1PXj53YC1uI1t2YCaxeBLuSFYnXxVO+E6Af6oVDnV97
n7000aTwwrNb4RWB3dfkBWgVovJIlqazoXFuL6FZ1BnHyCTUfO08ym9S5XhCFJUekl8qOBDHu2xY
zqepx1HGCY98ux/o1e4SspSx+CNSzQo/AfOOdzy33iefSDTarUqa/kGDCJH8gSyGCUEA0e4jkIKJ
11/WXzxvcjrDbhMDMu5NyMRTRWgQhq0HyyQ7nYwCI0N9bI70VqpnKa8FM3KJj2OzpNKU2AUn/GXH
d6zbNbFKqS6DfNeLKcdRimkM9IiNkEE+YrkOMNifJMOpN19pcv5njPKKrrYili3OrwlAqzYV8/FQ
5qHXi+rL0Otbz0jhHOci1LBK8P7Ma0rZaXs/hgwZZTsf6oPA8rLu3s2wi3aFslUX7y2urCFjYzUm
TSPaFb97/MDLjd14ml7odfH6QILwwwpVdBIfkO29cY2NfiQL/utxFgNuK0YODYwhDHYGDhpVeFIt
zLVgnexA8F0AwW9N4pNoAz3iLhvs78j3eaDO3IonOdwmtBCaaFTMQqGRnPjGOy+rx8WQGS1Wyatg
i+9HRUUfB0xrEeimipPDeGtEgHqT+pDRCq3NNut6mL1wDY66b3DaJ13Ev6NRPwyivplwH2BPzgrY
6mX3oaBpbbCIEg5LoXSlLI+W5d12AtrSC71+1ihHDi1UzroXMsx1FfmLinU+b2D7sWa3hZuYpmsa
E2cK4bRIJZLsu5MpraE+n/5d7OYx2GAZ5m3x+d2NWywFYvWRzOcO7b0z0C/hIrMbmip5aExwPjk4
T2GMdjGTXzZuj+cTyyC026MEwwZsLXPB/PUI7GeQwRD6JGo3fU14Clvrqp8LcIVd+4+C/oZSv+36
edlJ5UQD0/4oZ6fHpPU7elx+XyxpLmf5KpJuUcyYYy409w7vVtmu4Q5J+OM/eMg0BENFewR5Vz2R
ix6YmuQjxhDmrV1n15jjnWRXsgUwkQCr7R8oEnPsMPuL+el0z6NYI11yeNAPCV6cB18IFYya3j9A
8hBfE3CY7lvtRrCSHM9ZFTpIxpksC9CSpKYC49zN8QpmdnC2iEFgCv8X+qXG4JMbRmoBBH15ssRM
6hPJZJHLeLImHvWoZWWjoPW0yVGGd6wMuCtUsseIzpkGthjdAAs4unCB7rvEmJUI/1ycyVZvMWk1
mVT9HulBHK1A+ES0vxNd3R0yAtJZ12dvduWgYCQkXAfsNOA/rl0CIAhEAjKeNxRCI+ljkhbCcqwi
/ejGnrqzp/DjSXpGI8nhbb2XbrQ93K9dDO6r0JY1oUbNc1lHOK4YWpWfxH+hn1tpw354RaJtkQV1
ICwEgfySwtBE0G4EWvK3jLIICD0H5O84D5UXu7mjXijETY3H0NM2WApXcmBC/bE8rVbcB+RZU51H
ctg65ICasaYp0cB0T1kyQ96+8KxLmTfm53rzPW+cyFgrz6QcpMaLeUEf99+kUxpNcLQjX49OdCC2
V9Qp14vInAuFipG6oeZINjx3TtOytocI5k2JQH737XqGi3uiRPbY2xmQA9979bFPvg5bf4PoT8UE
D1t25yNxgwIqT7JT3095qU1e9mceP2n6vq1L2CEFAnsws+k2I9lZMhQ5NW1z7uRjtBisKpLHn+db
sC4i7HqVBmNY5xtdxFGioqXRFW0dSW2P8FnJbmo6fe6YjyK94SOJlL+tJSBHHVsQDb4b6DU7RpEC
cdJoLg7eyrbzr+ILCXbJLzj3gDYUaut6vy5cUpODidBgqepHuSaFwpxB2uxoeZ4qkbd9cBuNY2nB
PqNsUefM3VJt7hqSRDXkUGwr/Oh12i6WHEU3QZ49kBL4ETvqgI1vK8iIKzum9sPWwadJw2h2WhhN
Fv75XJSj1g0/Mf0+2VHqyZwnNUfyhPHCo5ZIbE1DFj/cs+T4GT1auSD7AMC241ezvys1fxw/wI4v
fey8CuAQuYgH2tmmDnuZZYTU5Wd1qB5C8O6LaFFEif4ykycnAQGfvFmT6NK2h4sOK/k28Y8BiXpq
cyl1swcSj95CrB8Fm/43Z/J5YRaaK/bQM/Fm/HMD3puyF8KbEcvmAJ3o8VWqG1aryNhqfLwZc+Jn
eJoLY9WtmtO5RJcdOLI8idhlm0eVb2vb2uoKFPCuPpIjWdtHelNlbueOnPIxXJSxdTdA1LiYn6cS
UAXf1pKZw0dohHBmgpKIEuzU+t2xRmSTOTFljmoPnrV2lpPsSPLWcJ1NvkreFhMlcq3TeTWsZB+b
epkl+uS1Fro4UONXcoWwqe73x4YZeW4vN/0pCTWrj8AWuIsKRNKo/zNg657pzRvcVdCsd8mjklUC
5YEICXz8HRbd2P4+s9PsF8FPcXeSSsKz/4otww/h5M/esTIlUb3jF0zXA7o7Xe42VjKK3UzST8WT
ptm+X+MExpoAxpFZufaymmHW02Y78amlBDVFMz5TaOVSEvXtPTfPPIJMEEttGMkWUuwX5rETp7GP
1FIQxkTWts1ifY7vMW5ue6dKeAgGPMLIUg1JDvhMOF8gIyOL/MetyIuWwHxzITRidYEvCh/5PkHi
e7G5NyhMkyqHS8wcw3wW9DUJd5/2kOBI+QH4/LFxtLfvvn+4F37uoWslKtBmkgEYek9ynCFLur4D
5tpKRXaZF90fB5lG+J0+WEezPfb/XntvLPatcuckPF4+/TOr5I4TYxFlx/I+kXik09R6EVLddjSr
x/dsujDKOPLQ1Mkw3FvBFPqB9F8ORe25QSPbesn9/TQ6v0vJck4JBv5N2shZUQVRkNHErlz+/Bam
onCn2M1kBXD6PRzD2YHKyWGQko1MkR8R/W0DHw+LV5obkW2E+bvTQtT9ecJOUYjNMaQe3sP5w5BI
wQr6+CrJshaQVR2f+J1CT1dyNjHZee56PBYK3g1eqtRggGiavzihfIYNEW7/yRUFoEvBnSKsKWIo
plesJYGCaor0Jp6+Wy8f0c/soZWFVUvZp92ZZYOqfcxsjM+tHDtNIYXvw6y403xBmVg4AT6eUtpQ
Go0ho3dpLiYNsmZDUBPh3G+0LH9qGMFepv6S5Ub6GrsZxrVrKTJe/MGN2k+KsCYuEFOTiJPwO3IT
iraqlJCojgA1oPAZJlofHAEX+9aZ2+6E2zfZUtBWgM61QlEWrptW7IAqZHN/5zuGQXxkY7CFabM8
qR72r1CYdPL41oQ5lbnKpU+Rl88xvLSZdPXT8phCum0Tg1eHAp38eNAANmCENZbnxxgZioEUc6y+
25GJMHxicwSkMO0i/LAdOVtMK4a97uvEmEnfh3tTSFXENYMQR9mJ8li+EBzsBaWg1PHeUSMJNRvr
hMhXmpCQJ2d73jCC/rgVk+ICY+uXidS63mDEeyK5rA9OHCLzya1spKScOIRQgSBOv2BXfPi61Ufg
MKN92vw01fHW9g4tDzFAGulV/G4PhdarXyG0GaKVyjWdCs7naofvVMV/ucPJXc8ObC2dcHTUOj1v
IrCym+up4MrwQgMNcw5GHIDL5SefD19tm+opp43Jj1vsFNYhbQPtjiA3iVnmL9WyamFTpiwBmKdb
2HnEbYrETmGflAZJeWJpcKm5IcK+pw0v/hER+/2b67FU23VvtIUov0ykoswT1aOZUX7kUCW0UjnW
/tfcplTMXWCxvqebPWoP+zmCJDefTWHdGnLP9RCsJuyUzoLMYnCeCUacuie1RXKYfp+Spw7ICGe2
FGeWzp3WPGF+f6cwUSnvCXW5JsLuNmwg7Rk/vSAhBzJiWxHM5+W3RSik60iHzE01G3AFny2WcORC
A68JIJY+nVM3YnL3SG3uDXtSWz2ngCyGjDsncw3/O2rNm1TTP3DzLzYa7TxGUATSXD3/du0ndTn1
A2QGFM4qxivnjSR++ujJmsmrVWlULeCbVgbfGoZIwpM8vIefmtT09a67NhD4mC9LqtxJwBbbzZ1i
9r5+353C1i/jq0H22IfF3lfPvSi8f82ZpIazpcvCS+vo5I1NpC8gJeM5ZcjDhtqHZWc1B4f1dp6f
7j1TmdIi9njPZy5cKNterncx2i92VyNqM55FysiO3SqZguCFbIkxPEWRH2Wo60K4BihTyNnL5Y+4
iPtJA5xaXPWwuTtIBn4J69kcWv7k4HYd8GeoXNB3pNPV1ER9R1XjOi6r8gAz91EF2EJVCvXsx5aj
umI25WLHj8qZ4jnuUe8wzp3ttTfwxdjGKA9hmd6FGjF/qAByj5dfZhnGncg0oyOx2gYLslsN+pF4
Jqe9EjTGGO+/d8G5Zs//c7HpX8+uf9JpKfhkd2OO225w0H7fq4VkiTeP8EpO03igQ9XNeINeasCX
dh2XW1st0RKH2bHpypATr42UzcWyIzFDJQ4jcNGCvoWcY92Tcf9NVqojX8mORorD6FneBQHCXSqu
5RLSmXgsg309k+y4+UrwUUzPBoaeB5iuwBc6XB27gVgPzUzmUeLn3NSo+s+d6QmLZ4SD1dsA7eYE
Au05lbmsoPXQW1+z3SlnOq4BErK/7zsXhf9y2hGsUlsmLx0RKlKDGNabGbDijQ+LApHC1f95wlAW
lWNYoSoW+9gZdsvs6SgDE8jZPhKHHWKpxGZfoKxJJPmMdAQvWSQkeqcPKRoFxp0WW8Iz8qgPo7CC
MZBN5mlCwStxgL6TULFb6+B2wIxfPUYaT0SZlijpp0yMhVxbAQCZ6kw6J3OCjtYSp/ykGB71M12k
snsonZjgk1gNt4+/UnwyQpDETZNabtw3R3f88bTO0BtoQiGci9seNa19lfGTMocLtLragAit48v9
Rtbwk/twcw/d2/a3aO1AqGKzOeiY5/12z2VOMEoKKD18x7kroiNIAXWqjP/J6KPQ3z16WFExIf+r
uj1kWJ9ZOiay7+bs+m0gu3OBe2jIEcFiAI9lqqDYhW0rBSdWO9v+FsEXCI6g331APcP1IHygzlPt
kjG2dXE109dZfCbO92pVRUVtmWjX1il9tmUsx7WJIPsnU+5XY+ZZTVjXysfAXmQtJPhdVRV/Gc+i
ylbOhu8seJ3Ym1HCbrgSQJAp9SsN0UIdFfAkn2JRumq5Bm9aHCME7OOrSs2ZyczTHFvfUj/FNIgA
HrQGqQjIm9eiXbn14HdGo0BT/gAhpohcKW/5Sn+EzEc4hSjZoYvXwNVkW337TqdIBbUG4nD1rDTB
pb7iP1so3Gq5BVMA3nm5ncDwpKnT3nWfJ9FT6hKYG+0PeeOqB1SmdgUlWtUJmGX+U7iLEKpIO6t3
0ygr/coQWaoKtwr8OlWq2ZRFKxqWsC9Tio3S/FA8aenO4XYbsQvdHw3Z8/PlpCU3gkNmIDEOjKrg
KTl22vp0BSniRZ9EQ+Q89g3WF4Zb24Zad2i/LV2ofO7ztF4w4Pcw4TOmzYKU4OpMHf/PLf7q1gLH
YQnPSXHb+2MFwDMsvxlNABGgHz5A+7tbQkZc8PsgmuWi3XUbuk3iN/PmMhPkEGa0HuWzmt+Opop9
UWyYND+Ulcplkkuod2UzHBcGKFKcCd3I1Up5gB3eIWvADY+ZyVWiXOOIbluZ2BIH3pqhgO52vK6b
oZJ3EXyp6aLYe/53tei+NYKM9RNB79RbTrtNyC84kGJDS4RDjcvY/nzT3nTgAwoIyhvcDRkR108M
2SHfQ/YVTImrddlwAdUOmyqIftESAPpx4MLTR6NrREPfmpp7dUwBL1u1mv6xes2NrPJtrGhKv4w6
xrrkR245G4Z6FBh1fMZdL3Jymm109qifJ9+ugg+D+WHJkMfm0N8V95mU67jRWrzRZxVkU2o0sMla
FBYDMxoISyXBNUBTqndu76xHnB700fEQWuo455ahzbEJGILMa0j8DzWZipLDHTP5MhI+LzAeOIiF
XukcZ/IE+bbNytDKK3VetsVDDkPOQGrPd2Micd38l4amUPqkyyi8lIcSHN8TJnXajCUYv1TQZ/0d
TTwP1L9bVKJIyp+35S7VYebzrNFXMLFCOI43faNBg0Y96bfPu6Tui3Slp7P5tYd8OB9yOjClexji
TQyKAvC7Ba3Hz4Uk592ufPHR3cp0IW+oYT2wpFftqnuy3DzUX3+YzssYETBEQMrSthlSzgCOROJw
ro4R/FCMX8epXLB83ZNu+ylmterskGqEmzyH5F5T0nbDZnjPwjVIjv0H7b2CKXAbPcZFh6CJmLW9
RXgOVKzg8mSNwtowJLQ8K0XjpzhExjpfLqGmX4c2IVeS41I2wMUFHoGYdWiFDh47LB0M0oLtKloR
aRY3MsC28G/MZwuDFPVUSbsMkCO+999hQsI67O7+a1akGXClzWjKIvuONE7kIMKtfYYYHGOH1Kf8
Rx4oCM130G2SqYlJzMXyJp4Agq8f6UkencX8pDofdt+B0SZc5qPTZzAVptoPwk+FPSg7734OLI5a
v9d6g9IRj/Ija7IEB74uU/Kf/j3q3RB8AOTh+nqRpdC6OI9kaZKELFtk0T32nyvhC1pYqx/Zyke3
nQ3lxPkAv+wkp8J5VHiZmmzWsC+JiyHkJjUT0tgX8axVfMJFpJF8OokxWPmTub5lvls4lhbOEeMP
6ecHWecoG1+44z8g2pC5LiPPeBrxhxzkxtVA/l4asXn+y/EuX0UlkXA5idYPBKLTkV+tFMO6rXoE
kSRcyMWldLdXpOjLlssSr5X12EO5sOFWE69x0RZW8MeIxS6CNO/+mYB8Rpqz5Aq+BjDt/SJXUqQX
6H1Xu1kejf9TEoAmb6GS22Xhb+uN/+74FTXsFqmdBThYLKfd8mXZ6g+cYwwIMkaeTv/rdCHhJo2G
msECmGbLcOuDdquiLEZBMjJOto7IGrxZ9ZJdOYD9hdd4yAe4akFAY2zi14AFTJjH13mnP1kOQ1kL
8/qfcYWZlji6ifGZP+mGdyUkMOzkxZ6Ofk4e3QGa6VYsB3uGLPGqXo0CFO9I3aHkbQSofpNfMSof
4dbERUDNi4us7sqIO+OaF6T+nMHHOwhdmwGReqhsbGg+0T6KJx4zWpdtGdIefTrZjR7OF65Hw6/t
5ncNfFrag48BI0kJoQSmsHxNtUSxxhwigg1BWgP8xyRGjU9qT/Vttsy49aXoVRu5ukl8XFOzyqfx
pSsmbQBbE/H5Zk0x9xLnpgm9uQo5L/wrcbAkEHqcaObgc7ZdzJ7sXenktvrUj70o1w12LOF9pnE2
oVsdOXffLaluwuIlXUrI50IduguqP0yCvJ+o3EoY0h8gNR1roEhbC+6yW6tK8KrQjsjPoGZKCK6L
3vtsfe4a4UHVtQI/4drskp0U1w4vtMje8Q0SnFYnMFxwLbUwGfgadCw+3oVuusezwWxS0tpSHh0X
yf89EkrhzAUWJH2e3a9vcbNvVHFxO3Z5F12eA+BrfPfes9cfytdnDClow4Oi9HPAYYOJayE1tmQT
keo5/Y/Z70lpyJRBudg90Xx1oNHpCJvqNji8ZLenxU+MHjIfnMmaQflTM9pPbjV3stkF+1sV5y+M
+NFdIShTE3CoS3GfT1FYIOptuV1+jqPLgWIa+tHC2IFP1MWwEJumPtrAIsVYYuGqTcMOoMYbJ9/R
TEMxnKgCV4fiygcRPV9gl6dcJR4MzoNN0NfsxM2FZ+QetZJOP1X3JbyCpUpfuEZyld6BY/bu6KM/
yGxjoBODe1AKdX9JUQuHkTLtNalP91XaZ/1je11X4qyjvhd/LuZG9SYP3C58shrKtzlhdwiXSV8C
vhfXIZlDGqCF2ezI/ntkCdthV0J3s9EgcFN3AHEDwL4lYS9k2/8vizLeO1d2FMJo1uruo0jqSUAp
u6ypKWjI6uvpnoLdmXB3vKRF1Wgo/quA+j8PFQCwdE3fVqtwBCQNt1sGCK12eQIIJvahhEtaIRvL
8rH1hFPPv/IQtIL3rD6/PI070Cm6Xc+bGGlzKJPmf0sKSQLbRSIUklojMkRj/dyDBlAwvCfWDO2y
sW0TyRsxp9o9uUCM/LRxx4VKRxV+yaagNjoyYS9YWE82VOTZAzwFr8Emc5wbfn4j65NEcFz1T029
GCBphdi7+Sy0Fv1cGQ6ByWNQ5eYcYLiyMm0e16AWIAqDpnGEU9T7fN9cwB73xWd/e0rvFpJQYZOH
uGoaywspYIIzPAeBswai3Yc5MLnNjyg5PUL1KMJcrduHTZnfESdeofd2+gFYWIwLqpby8iPBmu2F
ncfRf6fHVKhUwdPerS5PSFWtPf5icWYXdhBtlP5WB5xKCwvdj3q3Hd7AhH783ruShjJiC2VJSCc3
D4zP3OrvqQtHupFQ3RkBBrMRk7kTTqCxz+Gis7rM2QViWPniUp6dX8YpeGoaacdIIHe/xXt2nxRm
EPpbUyOCWvOL/ESIeIU032TMbJwTRnD06lvfysC7LpnLmBmaB7l8CFwDmVzkXYtyC5vtoGO2kA1m
1H6bvC/1YyNwvh9nGFC7BoLwOqMsZ0tRw2uETADXfYxfNfx0xwQZNPaoo+oD9QS9KVU1/ErylseM
bawHeevdqkQFYrOZEU7cmG2VrJN8W/i0DNJgav1zDGeiczihWRRat+JTYcqt4rmDphGh5UFvAyPz
Csjba7UmtgtwjQsW/QCe51dJaKuVbiYPxTGRP1vbdTBbshnk8tACrUmXVIsmncr8T1uEB1LjuFqE
kcsbkJto6GpJ+MGM/rCDA5/fJ2FubyxRBgBw9qUwKxjwehSUYiFeI170QUFxhRpeRlxa/R095w1G
Ghri2v15uhKOrzKgIGAOdTuoC6G/JTSOmU26RKCoUfcxW6bIPwfE92sNIYzNkThWI5hkSri3zLQC
QxhERqCtzpyrEHJBo6xncb8FoKkQrCXsD2V4y3qsYk6rUISVzblyLGdC3S3/KokQiB7G2hdwqhuO
54MyLlGA03iKCYViBVggCjPW7dbUeir0MV+quo4hAqteM4VQxsYm7nK36NXYYTmLM4VRnz1gfjtI
ZWpiZBiMUNREAk73zMhjRRfHNaomy2FI/0b/YmxWwdc/3mhaih40gcmMxmnZQ2ZNYAienFTUxl33
K9HE+FGRmi88jHsOa9b64UTitsZHRQGiq46MwXeLcSL7/BQFrFSl6ZB9Nl2pHeljpCSCwHM+Y8XU
WI38ES1LUlkO+vExn5RHT6G0YmHcbwseAgmL55XGDo9nUF3c54hU0UfQIl1pbHXNCNU5LaLPl4+I
op4U4eRSDmeCN5BjxukxoMIK8XV2YiedpBRI1FXFCLZ0YAHUPWRDlK1esQU+jEBh0FbTGUC+bLtd
yLVkYJMa5y76o9pYqp4/khcvnBoIGdysrhiZLBQVaGLxZhJuIZ4RL+7psE0GVYYUNCguipeUbPhq
iMDWJKkplNmb7EIZVrkQDoV8PfJ+i4y985nqB45UuBztYk37e3/8yDAH9Fpu+HD3l8Zv1tE783zZ
WjXcAfQfbfd1+uZQLBspfldXCKJZYX6fsaVihYDgDb2AvXOGtaHJ5eZERY0HZAVynTdG5CV8SFYJ
ZNzsLviuLmkONFFvhlI+NASszlOZ27SOHmtIjEufjBRmuRJFsxeIexfb981YLmSVUZG85kQqNPAw
Of77OZMkU9nDdbQubMFhJGzqATfpZCkE+PIVOjlb2NwHGkhpuBSJ4VclHPeavDdUvUX9TVKiyUsy
SMXevhOiFM9jNKSTGLvFZc3poOqSC1RhSN6V+iE+sYH0RcHPgkXkt6zk8jS9MC1Hr/hdiYp8yC6e
VGW6pNcnGVw+QxbPcpw3mpmkh7Rz5yp0fkAL9DHKNL/fRuBx7kgJhXt86M5CapduHGtgESNf787b
NFYl6XN9y3lcwDHjoJZXuGwpL9PtLxhmu4GXdxiHs3L4t29HB7cUYs53ttWV1S6+xL45rTu2GP1v
iZ60SEysY6NV9yodFK3cGWXGzdGxK5DzA3JCfSrtR/B/Uz8+m6MW0SlKZRsUlyC/1lO1le8JODul
4ZFyu54DzzCm/jvUhF8BrV74v80WGEE7bV/bYGhYMkg0Ik5ZBP8iqmmZ+39rvsJPx/nv4IQvt30v
/UCzaxJdwwsMpNNy4m81oHA2BgpyCQh8Km+d3ItxQMMqDEjMopWnjxRZVbAjZBujB7n01hc3JXzu
1jybje851DashdxLw2hhGtmXykjqez3lEnuknbixUopZ+J7p8pi81bfJE4omKoEstAnND+E8xner
B9hEOlDd3k+K5ZUu45+hqiVll0TL7wTADwvgyHvUcfpCncxkxtJsGO4Oi2NfhKeGfosw/AobJnUw
IzWLlwc7Hb8Vyy8PPiX70XDYrzPCQluq3lJAE51x/yIMRcIAswv7kVO+BhFTbbfu2/qTae3ypl5y
F9GrlGbMeYtvO4n0n8hCJLc4+v7lFP6OVgy91BRkcFyFFzQ6vw6ubRsdFZFErIN4wJY444TAXKdY
algDPYYJmsd7Kk+YqbCN5x88mC1XOVVg82gJnHv0eV+YausM8PEiUpDZ9d6MqvxjF19A3iUu9wOQ
nZNZYRTtU6q4bBh8OM94zhG7JsP3scFbjl/u9bH8kYN55jVgcIa9FXLcNTJCZ15lMZnI61YUOhHY
yFuWBzSHWAh79v2AiyHvZ8pi/Xs6H7BO84Dh+cli/ad5qkB8CZcouHdvvHkPlBYoU1qGf5ew16KX
U3/mGy0BTKRNFraBooPZtW6nBIcr+KpEPFWYS8uI4YFVp5EoRvsMoLzgvrP/FNcS3oniNY+pEp9W
xGWnW+E4YaPEapyoVq/SqFu/84CcB9LKZNK87ZZw4deqh8s3lvJneaFMPK502BcgPbmEe9B0P6pw
VYcFbBfFcR7daHzbBPbXxJdRdOVuJGCyCNa6Dqav979Y8JnjuDFhyJY6eIeKNBTgo3ZWa+o9Oeye
PQ2LZcQYQAOJMXWmvQB1nXWHgHFQrJhha3KJ3m3YNz/Mc5HoGFz/A5M+Mojq0FSUgXbWCcNXOAPf
+OAcx0sgvRDXZ7xEi+A4Z4QevNMNHKGnl9kwc+mQTtRDW4QLRIdjyR57s57gJJXRheo4QNN0GsLJ
K2lyZmQl+Gtg2+7Zw2N0A2f/mVVaQs81HKPOSHPdA2/R2e3gatmlYxMpaJ7xVqfanHkzYwrcc7qm
bONsG8d6qZKv1XgIKe0zEwZz4W7bws1nOVqgkSKaUdW+BABQTHHo9M096/R34j9XnAfIUj1XkkMS
yNX3jj1pdGdB1jW/bhElkiDRrwNvxgUoPHeillqs5K26T/alXXqr6ow6pMnjxq8KodMR2oII/XvR
lgr4bm00KoTDdoiGmiulYeAS54u/8uK5hVnQKneVRuK1yEgbptG1QoTat8kGWs4vrTHDECdgQjWa
M/YzDZ6LHZez8pio1oGK0C57RTx/rcjwTv3SQDMN+ukNuVJq/t+rBqWFVFIAfWY1tG4vgUTnK2k7
gQwNPO/pCHe1doyRJNgJWtXDzfuu1Ihd3yZwfhEOeMb/arbFGnYLwDPPTvC61++/ic41obL2KQ4I
n0wo/QAesr4LhRuKbDg9qYswMjHIwaIBrzmDTOp66yTtTv2qe9QnwNGeLiYuJ7byuXbPcVQN/o8J
kaW3yWqCtlPWjMTuR0M/iL27ip32CJ1ThJXv51IhXORDNGYvlJlA0klkAB/GtEEdr0bmsi43+2un
pztrojiA99AtVBOvKu7sHAiGAplDM5LlPHXAlFjnH+QAfo9kvn3HURsAMtE6voPZ7TrvQHI93ReR
iALmMUWw9d/xDgHrQrBFytxwd+IgAqttbcAxYymJFgv+sl83sufX+Fg2+rwYVbRhtavSwNWc/yhI
sxc2qhIUjvSdNncVBCQqgayCIWace7nyYu/u9ZEUzWyIpmQE0i0a2Ff4EHAjxEkyebrAtMPGk0Dv
pv2NkS3rEteRx6gxdwukepdo5XdsoWHWSjG4UWhTivkudmMpzHeAOwkP3GiWRX6fQ2QGVpwP+fu5
6fuXLtYdQbaJPIIeLpONAv7BPQ/HKzzs3ytGAlLKsvozdPS0xvqpncNDc4IKZ21f347c6Dp97zbS
JY/eAF39dZVRq0MHLFBR00iPVkitZw0dMajj7ICCFcMI/Sei3RZlcZG4lveDpb9i6GN0gFA/jrHv
Q2hihLscA7u5uSicv4mUyxjKhhG5ktj8+zYkiE660iviRE0ivNFWEEpDbPeRNqUBYzWKsZj+OmTZ
LaVwSKnJ1sjQByRdmymyDc17U1QonKNjBRdwHuqpJMY33DVWI0HQVQujIW7Uam5UfsfwmuHEjk1w
wzzpH9PsuQPDLwsN5G3YwdeYurmWJaZY+OIt0nFoDyd5VD9QKvGygenkGyWdRrlLE1BrhfX9IW0I
DfOGNKPxxpr2f3jz4pXdx+3ICfKNOemTMLdpwa0NI7q909ELRyX58g8bVii3G9BPprfDEQp0+QVF
Dof/Ecr7pNTt862h7YkfK4b7AIigJDU3Z4vyaWigqqWFAkAw1LW/J9Qgzwtgyyq8kN1xvQ3u03VX
VN/p97RgMzbTJUBJEw+OxUk9jcP5knfLSz+HXz17SzSCdKFIJo5HvvWbvQGD0g7nhREqTVdbcLLA
MF6agpchiFLnOK7UmeaVduK25Ut61dn/7Sf/avNpNH3usOst/9Psn6/silajext39ksR36VDr0Ji
WiCeFyNHGIKRhDBZSfBO5XTq4l2+GZ6i+YwbO8aGTgsHOedKDIiyv+nunlyW2CaFGYZ/HG2o7FEA
FxvUl3acRxI3N6vK/iX5MPTHC/WcnaLvGQGX+3xDHa627Ypvf4zuJsBIRm7scifOuq7W8+ckTZZt
L+43vcdJDgnJ+UcCY27wLXkuf1liiuVH5vRvNe2xwcrVDPf5mvWtUAejH1l+3628JuDL1C6CwMe9
ERqATILjv8QVS2mHu1sNK9rVA/2dcs5LZxm4x12J/ZuS5F4357WgQCm8sGnD3DqOXwjC3Pz1fO4t
1ad8R1F2CXrKsU0SbURC/RfQ6G9nFzhS7i0RQqe6BJER+m39obBOxOJ3muuYEKiCLfNVs4AOyB2+
pM1GXo0MKk2KpB5oy7C73fsnZIgFifSETOmkJd62i4L8F40SJXzM00LvlYsGn1uEI0UBpNavJ5it
rm43UpBmK+TOnlBA2+k2EpqUBJ5obBCqiY5GjaNzWuqGKhHfPtU7mrlr1z7DN4IdfBv2G5ecVpIm
y7ckbHuGLtibOgfSRE/4ZEQ7ZWkWDxJS/0roGogSLvcsbnWRHe8jIA6r6hBpx7uflFf4pcmZyf2i
v4S7A0Q7yWrPUdkKbAX4O/Ys6cmQ6rdYZCOuoZw+ICXIyWP0Ccl6rABMNVn+7Q5q3i04mcjQO7s2
2MbMll1HyM2ncIfeCNX1Qnvm5m9OknF5LMuGLZokmlKbEoeeE3Tb8EAq3ePlgG4Raia+MwbL7jT8
1fQcdx9jf+eEgCDnU2clFvScMvSe+zbR2lk4GrCehjhJvo/2GttnpxrDZCOZFt8Jpbe86pqh5u0X
iOdHt3vENx+TpX78/iq8EKrYutvQVsAE6W8JufmoYjo/i2BIdYKtSiIX4DFOkUS/7gNXVx/w0n7h
D8pGUL9gpMRSbkgncWqLzoX9/Iur5TZxQge9k7gyGGEl6K348y22iDUQJ5Epi6wwXhZC72/1klsB
ffa86Uj1vB2eBjk87T3l/mGEzzNS0JtxI7y2MOhugEd2L8ub09Zxx7k/5TyViRRvBgArMV025egu
0mz58jeZ4lV/Ss/xnejpwt3YnKtcnFaZX9h0IDHOJV+Vi4JbAy+TWnOOYbpLDw+EDxkhfHMOrxDp
gIpcV2qd4cLrcmBa9irReqAhog/DASM3Q2E2bsaWrf/jL+EfpY1FDJ0jmB9b3vrIUTb4GWBJ+G8X
rMd+vXoTHtcK7GgGs2FHiL1LzbcZfd14He13BgqbGsyueGqdvOweOemWZedEOP0ChvJf7qwWr8VI
qrQpwHGLS8ruCm3rumn7M8zKyjSRBoAx8WSKEgjug8Lcmwfj4CvKVDCBIsi0Jm9nb/Z1TDp7ofoD
2P8wl8BHqIemCv0b+MOvemtqrTxOdRN29tUtMq9D7qgjrqm72yNXpQ+by08iWp5uSX4qK5llQFed
fchwtkk0BvZuFuE7yl2L16CAD4tzAZaJ8vnnm6OBDmnwGcPrg+dJFmSkW/JbVei6zjUb/VNoAwhf
v+TX1DUgXuSE5GNEcQ38QyIcCAv1gVvooFWHmY+uyJjN5JVGb1E1YQ0F9OapdJzsPahrCMLx2xIY
iXbO9yHWv0DwMA/LkDSwfaeuAsFsorGgh1mUTZLoiblGfK9dmAw51RUu+Wn7tOJlXjQ8shZKZknd
+8uw+Wh/X7zWPj/Ycw+lCYlQFw4G6a1I865B2GmgwlsCjhZV4oS42qLmYD1YHlqxc4lDeETjAGaQ
cyameMLllcr6qQf9Kvm2hQGleFCe4z04bPPgga9Xt81HbbdSpHP3cJ0mjm9EqlR27dBir1dVkwXS
RiVHRjYWGOJcfGEHGGAgGKWHsVYaMc5Q8vWL7BPDJa/mrF2XwIl9CSDFmrnEWaZFXaZ5YAGgSriK
g7YDaNKdvvoG4MUry7R6b/1nXpWdcb21uUbmffgUTuDLyph87KHDVrMTMCr6bHQ9BTAaWrao0UYt
wb1Mur1URIA4TQ9kNxd53ECMvCLXtXH20RBneKnEZa3lD5bDEav2X7Q3TWiEbI++VsiMphfUHcDP
xD4foYTmUMpQ2yp+6oTdUco0ZxHYwU0jHar7D/HM/RAjNn29y25FWsxgL/Q2tmV5prrx/Af9t3IK
FtFCg+MDM6F0JaxEot+wk75OVrL8/U0ILnwGVS4fDM/OlVBA1X5uFQoXmhmos6vQqpKBhZgNdMN4
N07T9eE5LnJzJ5zBVHbWmIRAdlJC6p9bxQHsdvHuj8W25R6ac8w/VpJe7c0UWp9M5ozr+vdVkcfd
5UAk+iPllqMS+FTY+u3v4Jr2vJYZTbyl0yiflpQiRtATiChOrI6GAA0HNdx74p0lDs8ZBT8QTmsZ
PYVwZWCE7UxdrnBDN78UuzkLPMOAczjsrwwTZAfr+8DSX5IS7wQM57CxdEd8JDyUCl0eYP0cSrhK
vpOAKLe6YLiUuRLdxYG8mhaHuTYkJ9YkNnMGjD/Fx/IxJ1ORNaFi/TwrooS7bk9D4wHpJd0cgHby
C8Fxr80Ml1aungQ0+NsLFgQD8g80c5ANB9IjxYHXtn6XxvcJItAZJk0a+AplfW5EZSrbs8p7+33c
LsfcgsnEyDcSoOYc47EB+IDV9Z4kmJBsCWwHm/FyT7oiOPZ57MQ7vuWlAdUIA68sjwseHFIrp0o4
ze5JWSt6tI0EMFIbisCYJ/FaMjHiU9w2yy7diiktJhD3Gh8YbZ27kZ5Vz3w2ggQ/i71EXagkymCf
OgJWM7fg91AGc2FK56N6zOCczgphQ8GOGlOvzOfJ/pDDkFTm1JK0IcqjKvpc9b9GWo6nIHk+HlCK
awWXtgpZhHtUJZo6RHBkmneMKTYlRSHgh9JGaWa7bgjfWZ493OXShioPNkmPanpo1nIT4ez0NRS+
v53k0NHWkvlvbRQSqYwg1n1rnG+/nWQbWpOhOq4DjBFSYip5F3lwIlu+ClEIcFWxCNdXphQyn/+y
/RY2NlOsvB67HuRuFzn//179+clACg2yF4U41CVbrecqp18Bj17tv0DY+CvQ3qiTwcDJohsr5OUy
aXBTlLUvrNBlaWCjmOgVXdGpj8rpc6QNmpS5HiXYalQ+SZnAKLgHFXmYzQuJEqZGECqoOX1DFDk4
Ak3E2voUBrgqEZIyiqAx/REsE7j0uCgJBQbUgVhY9CckvDvQhwgyxL6cuVSLTRkoem0DWi2DSEnK
+7EfHRvYZDkkzCNn7MLX9TqbBnqQhCH/ih/h4laBg+S8x+Wc18fgBPpteqi+A3UM3CpJjMJQA4K5
hNYGGOq6C5hLuFkAiqVSAAf9qz8+YmFuBp/2sFNIEi3WDDRyt8ElNNbSG23F16RSzaqjgSzePIYy
g490LMpfujT8J+j7oCKzrTDx+UmfKC5GeH9qJuoAAH9w1y11kymUgkCsTqdH3Y8/Tpk4rvpp4cd+
Wmpy4VSvJKi9ySIz12cGqQuTy/fUS8P0xKo+D8gNGCtpKlMuR6g/RILnhPZg5qxTI2kgME7U/iq/
xlzQ/VS7R8hT3aezpiJhEMZa6p8YGJWmaiaO9+zfp1TswuGfU/9cabe5KlPkRKaRj296IFpUdqXj
WULxbj13iGKmhJz0WspVJ0fUd/Ah8AIzZG1tfDw4MFQ6liTELiQ6F3PUYb9OAwNu79LQKK7rg7E2
YlDSmMiHymD+er8Zuy2b1lvxgV1Z2w7MdAFcGzrYqsptadP9T9Q79j3Y3I84Unz1TTaqAR4zZ/oM
PA9EKmJbhpYv3GpgNHRLJRrGUB4E9fP4Rqo8Rhl79yYUK5yhvw6vWhSvklcVcpi3quoPcn7oqEVM
6zDNUL6ZsYFbW4G5SeCcCMKn0kZv16kfYgCznDwbJUzaKQ8+kWvX3bYj/JSresIRoYZ+oXm+NzcW
ODljqmP0cFlT8MeoW/hyHGY3ZbLVOeVbXtGVLa1DhtD5mj9Fd3bqjVh4JXXiICbItJsGlOig6tcY
uiUl8KJ+01f3bhAA0pL3HeZ1J13vPYQf4APMUaXYHZ8vJklahCFsbsjdFEYUqgslFQuQZkfneSwe
HYkqUtDfZpNESJQc/ptLg3pL9bXdXGqSUi8tJcdWgCzIkFa72px/Z0ybOXq3lAR5QfE4x2A4nbSn
BxFM/dgrlxYaENhL2ccmj9O7buVZkyUkRdv3FRikt9BlA5gQ5eOwarf7YtEmna+TR7K27ju+J1zo
NxGaPEu2BUfVUH6Jz6+eCov8qT5ncxfI1JJbAfHrxDWZsEe+0GxulSSy7kEC24hC62BPqShr2KmL
SVLX8xMTNgg8BrGfrInoEOSio/FY9FxEYOTIb09GSIIvfxwXmeO9/O6yCdAQjYwwViCTJa+e0Rcg
H5rt1KMSwpPSGuF4NSe0KduOp2sdVmu4IBCk2cVMtAVW+YMT8J2k9AEqXUNFiQBg0hCMGWEdv6Fg
JcrecptlhdQRRpYk5bsnA5g5ql+BmoTQszIq0GcCRCizOVknl931RPwonggO3q8J5dOeT30yLiyK
e/Wzr84vWOVSv/H+loq+LOsFuF/+1mbOxOap9kUacHvmLU93OgraBX02vXG4FWx4ePkZkIqhx/h/
Kjn9DC8J+xmpjfmKcG4ealxmQeeAJbVPJPInXs9uhsvAH/13pdbzQrJQGhS4gFXYKy1gBKEuGHzt
u55fu27/0RGtMDc0IiCu++xyiuKwO4PscT7wLiMmaxkokT9sNXSTbJsfIH6oytE1DiTekiQdYM4Q
UjODO06wvxIRgpFu81SdfayE0eDXv2orcp10emtTyhZpjkuMJOwPOSqJ+5AoH+YBNLZ2xNdiypDu
dzfH3FmNp9pk7JMygvUi95CjPEv6s2RwRcOjI6RCGbGA4+Vm1EiONJQvaceKBjwzHySaYHhdCmyH
u8xBW+8TXTFg4mQXvzSek9yUjwQ4hG6gH+Ac/wmx1g5/A9cso3c6w+OmYNJmcuvYs+HG5y1UXV0i
Pt6v45vCWMPCWQBTntvReeYZqeDqOOAD4PL6auWnvcc/cMI+LE4xC/kqK0CJVIfh4nZLyAqUxIUA
8bH/67Vy3Hsp+2b6uHOkW9vA08L98zGyMoYhJGPl4yRKklHPMQUMlKB2Wz4aWK2WQZVsSrdZY39e
or2KRG+mY5c1GWE1801v5+ydx9UPsdc2B4CtVyZKWoe98rVhBv8+Pj272oItgS1OdWWbzl9wE7sG
8YPfYi/yftvrFQfQYuhuSTbHQ0SvNKWkS5b9Wcygwh2mn/dbas+eS7rCF/jwVWcDlrWCjtdeYe4Z
TH/B4I2taFy3XEHwjqo6sH5LPuf8wUtEknoGV+lwIq0nNj7wp8Cfm0q1h8X9FMg/R71rbwaSVcnP
Qj148hD/EtC2JK4ZQcQe8uiBhv79SUuubsyLVcQG0J+TGqn8ouDpebJbfRKKR9EtII5vrRVCZlbb
nfZz9dWb/fhsz3FhPflBVPs1V58T5Q889BvwYOH/Qmeajqnuwi8tFZIZBdVwT7y5zLSGPtSoj6wK
RyLCHhf840HBuZLQ/t0vaTsL614wNGBTKrXJZ8nP3V61+q9MhMVuEhxJT8fvQAiKKYCqBmWGxfOP
BzmRULODG+/wfHnyneaeViNrpFMl12DxrPfFLxAToErFLWLzX9glH/NKiu3QrE3rFthinmR5foiO
5t56IRBYrfrIcfHRPkZnXlJ86s4jZnQ43PfUxZwDwLb4BKInXo3MP6+cS+ntVf3+K26u6dDY0DES
/AH2I2OD4wZPdti0bNPamZh/SRuvaWDnzqXaWWfUcmHD68GXzESqIlC+hZqGCdMkVuThq4gm/Crr
jXgIIjjCjt8gFwxxmwhhWIOeB99WhxXjUdyVMy7DPOFv8YCKPimJroauEvQNenpqWA1TcqZO9nPL
qpXBvmq1MtcYF4Wzrxc5n77lKtTmRvDoxZgeu/FbviL3reCMFmRMDOwdKTxuuEfbxso1L5t+6YDu
7lK+szwyccjHQ2pwZZUo/uAayX4Eh+FEcw/dP0T9BqOMQzSYkIYbVZNZ1N+hq/iFCWRrhFju14Kx
xTTC8P6uElLbi4nWt3e2DKbRUUrd2it9LG/ELHi8tz6ofkrnLGy+W/TDkvAkutY0xk4gYgIkLz5B
uqVyIM2AqIVOAD934t5J2BI/haMecDC9A+ss/pCR3aYJPa93UOxIcKqUWEhhBZ5o+6BavBPB61VD
Y6+4jVHpltCRNKRpeYSsUy0doO/AMHw5mCxmh7kRd1Pi7qyNfeyDkIjeMHAwEWxoQtttIRsUyROB
/h3uBFX+zsGf6YYOqUF6wzQhBqhm0QVhE27oGBpUi5HIZVrDSMirn748Ds/1D/cQXOkuSMCnbS/5
72esDuBjk4eZSmHfWmYV1PT54+PbT4cSZ8zMyQGP62qxlMkp/8gSdNYHiIK5ypuGEi36vI9PekP0
yHcZhOFB4hYJeWgRGStyq7wpnzA0s/YqCZALpmEScPXvk6bq4ze9Gy9XYp4YfRv5ZpgVjhuhsk4I
UQUYxs6YFuS8dmmtlKide3amYPoY2wSJ08WqS22b0nEiVYb7l0AMNBIBbL01WpYAlfQq1h9+40tx
oCAFwj2ozvMS4YBhqf2Ny1LPvkX4hzelzCWgFycTBNu5ysbrhwUabuo8VvK7Y+zzoBPkjDXvSdtE
7F0ReDr4RJMGTId64cd43xy/TBWCZNRkpr3keITkEpPgiF2NImmffgDeI50A1qfuKdIta4Kvgi9v
ssBt6FtI/O0oRJunxzVYm8ubTf6WEmYNa3s54tNSIIiNJT3lrkqk9DHRTbOftx4qAghkOkYG9IE5
luP1zT7+57FHpZ81CDuyEinK4wQXviMa0ouvwzUMUbqm0KSGsM1CfR+8o+pYmwxhUarVM9fVVsRu
x/pURGi7APU2tHSmmrP3pUrFIsmvtAdPmtRwX53dAfmbGcLr25uwtF3IWpjxa3lXog89am9MVpdC
H41mcIBh5FTH7exOg2QdDHLcRBufet+OpAmW2P46yeIGLFBL51CO/OQ3dkiZOl3TkMcIPvVIbk97
Z6wKtao0Ei2EypPhpvuPTE9TMt+wSRUT980/ld5rAA96YB7AHiee0zXRN/nyLBLsr0xb1JCVFu6a
g7o9Q6e6UqVz4PuJ5cKmHQW8z6G/qw3gA+EH9s4DCACpRon6MAppjPQnCnN8u1KTixrs433rzdAz
G6XA0VByKwyLNTGYC6cqFeN42HaFyVZrAfsn6ghs6ioERQB/vLuWhVwMFesXqvWsuumOrxjKsC9O
P64L9sOj2+7rhO27IB0knyh4BWdMooQRrNj6NTA6Pd5TOUgJ72pHAe9I2OUczjzJnN6yxwuSiFaH
5csjqyZFekOLCyy2cZDc9qIR8TB0/0/UHgiGYk4QTDRCXO09ZeNaZIRPL244RLz86X+GV/DlNb2v
IStOq1iQWhZAZq36A5PHvF3ATfLvKewNQl3XiC/KKM+3nIE5BED1VG9Qez2OQ9tSmjVOqgJ172Bm
9HcE2eYKgJEZb1ddaz5OsfUuRSQXo7vWgyp9JGokZtBg6j/5DX2gMYZf2rKIU+xRAiVfXnqGf0YO
3gREYqWT13V8d16hInRaao0Hpr0LOYsqVe/s0dbceZrdZzQpoEGfxNK2Ce4GttrByd1YOmzyc1TF
eOsR2qtlGZKKbGm/b5vnI3ViaeUfVKfhO5LzbDTdE3GjsvTAVqDMwjFvJnfk5zwHer3mLumVmdcD
ZValitzFzDjsGN/XNJkFmKADQHJBZfNaV/1BBR1HRa49cnX0FyuLixUMkk+4MSIggUGln+FtoLVA
d1eAXrrsp0cd1vL7xdqlHqqZLtw/yyd3SdcaV7c600iaDT63bMEBjHAPZxNtMaZBM+iBg4PWVZa4
XMEn69JszUySPn/sHFIBOccjvHPauloXpWY3urOxu8CIPO8bjZHvQR4X6aT3wouvisAfhu7MpGPN
KbWeucXdxu4wH98WJRj9auc1AqzjixN4PnwlC2jSvb+30D0zl1jwm8YbIdg0W1ckN/w1PxTFArgg
2D4Lf7kv35Jycf75UUalSv9oeX4/bq7fhpPQ3f5S3yBVQP6JbQoEcYqCLhHA7xJnwJODF4cY2TUH
6ftp1RgHTD6T0OCFeGWwgkxjgdBITZfHvAREBPy4YPeOyJTtq+nVUUi9tFtFGs3xnu6aIMLzwJHT
eAQSODN8tZ7eMS+zZ2xQwvGp+QXgnI2d/BRV/ogj0xIv6GKrgGZ6vPzgAirh6hYLidqYuw0THOX0
aCbnojDaHwnYvfI4jB2vhrjWNd/3PBXWdLr0dskH8cyodh25FmTOvr8/QvLNcRKElGMr99LGXNKu
wnWfswB0zMtU+rn0UU4vgzyRlYxOmOIXlcWWW8t6vJh3ruZQWakmOxD8aUYaN0Mf4IhH7vf0eWnD
J22npG+UbYlaHF9WST4P5vY4EndSd2/ebgHX/l/RjdVP1zR09WjhgbFo5pxR8pxGYZQxqjyAWy2i
NP7mCxaYt2MPly3UPEGQwKFMWmuNphs6FabzEL4T3wQJujGyAXMKR4WvKtJt9oOaIMJ4ALBvFAT7
6f2st1xyh5plcvL9P0U+cm6BKNJy1J5/8hvAgJ1irJkVZ52ad6+nuSd69lMZpGm3uoIvSsK7V7/i
+EjFS2asmQ7j4RERENZaaVmXdv7r4gtGt++OcBPvhS5UdQOwBFIIVECmTV0sW0htLBHSaEMgtA1v
FLmexTzd6qHC38m1hPQ3aOVee4vrQeSuFkcKzXWjEzsBZXddR8ucGqkOGBK6QuM4SWXEHTFgn2Io
lJN9Z/ElEwoUT6nZPty+mp2pkyPUKLks02ItwN+GcTGqnhU+k//qQc3ULlnoFJH8s9pyfll2p/Zb
KyVdSjDA31XG7ZW0wlqKcKzFwTS46HcOKN3alNt/irMCsMW1xQW5e1RXQNiedrQp0tcStBVntL6m
JGIyyny1PRT9m5o4unh//m+VJCnlcXEJTPM1OMO0HdaKtPnTgH9QfEJVKrxEUQAokxkzPZjmdpaI
jR4K9gN2M4YPALqxHld/8hNmLL5dhnZ+mK7gZlQQ0jQQ1I4bxuZQR0TNed/eIbPE9HgGie/z358t
ou4ysF9k0GmZpbKEmIkP9quXWf8vC0pWIEGAGMVnni7buhGBcbg+zEnF5FpDg8rGl34kOZiEGahK
QIWMOcMdV91Drit2TQUtktdH6Ncjg7vrMRtiL4x3Z4IkKBC+Qyrkdl+33BIcewsYuNrwmXD1IoB6
SggEj+vQhYbMrx//o9XirjYFLiNA1Z0fEZpdmPfm6Qbg81GFURsO2FuAb/ck4EQLq4U/soxMPtX+
RQneqp1Op/d7VH/xxbeYzmDUWCJoxgyJSNj8sit4rBI2DrvITspad8G7AOLkaNhzZ7hW3S4X0MQa
1bVigygd2vhIvwpnpJ6VPITmzJat31YF11hglwH71NrlDL2Ots2GkAxkei855F+RBdQxf6YaPqfa
ADFPnwOrXAthSBgboE3rTmsIyD/yILR2sYTKthclcYt+qD9B4NKw5ggDYWSq3kjAuURh4gkWkHq4
nhsoHyhpOKubZuAVII141La/DcKptlrB+TR3kIdVcCFMYmvxUmnMhU5PgNQSWqsqn8RZrtqHx4Tk
6Ajowm0WYwU3WOcB+fNFeti+KXQ1Y6fYVETsoVA5TAU5zXGQee+HwCokmfuwGCubPMC8zcvsPIoZ
roPhMkGmY3m2cWXXUtal/fGyA9MBfsIQ91wWyOhkNNgSb1FGe+cCVRfHCjcTpyPrfTeg9YVu9hia
rLsOyksc1gRKmwTlOdiBhKVUoF29sBtGFQ2Y+BD837C3tTGFaVbqACA+HOsVJQpghBUZ0wlnsPW5
rMtYKBnnaa5CbfquxmN7OVW6sNdmU6AvpePWmFSKoh3oeOl4FWmKj+WVC+Ly01P7d2xMyuORYF7v
F0zmKQyQYnvNFXl4Qkm9Zwr266ncsKOm32pdpYHbBNN93dza1Q19Xnwy4ffsz8oPe3vIjLCZrO/d
E1h4JRKdlcFlm2kUAm4o1Df9rMXG/NvaRN1zXTu+ZNyMOw22chGTjPaQevr7TUfVb4Kr+o8H+r6o
VZWh93a8CyCluqEJrRe9cCak8hhPXgBFw12THNnCRTqPgIIwkzId7+psgA35/HTMjoaTq/RvXrD6
P8+P38JZ37HPnj4Sq+EmfFeAqPAjeGGCHJNq2p+0MkSrgmUGzUJOOhKtdAnAI+nvedjY163GTqV9
J676VhjHbhs1DMIKvWWKaRbq9J9Sp9elb6rqkR8rroxGzGa+7g7ef1mIIsFa1DWHwC9pnInAiXx1
BxNvhaPg/Q/8BzvL3MIFbVxkmd8twF1I5VirZOx+KT8pnXHuxDmdUXFapvGXU29xzBF5RYUBACsR
KRUrxKSYoskGyI9KJXyXpCSe1n/S8rjcJO0+ZJGPwSYZwRul27eyDmDbvu2nwuoz/myvA3FjTJY4
p7gu1rIwPtVgytvfIzrtfcdJUlLphEhC2AvGvxVuzmTv8oMVYQ64ph0oWuB3f/iQPX1ss//le6m1
Gdu3Ss27sZ1UmptLNnHSjmjXb54ZVMMrkt5CTJNMv6PYNekYA9pO8+hxthSRmVVfO8JyB5FMPjln
UNLt1+Semk7/bHnVlvCvi8nhZUKkpMAT9Pzfi0OdH2qc+z9aPa8bUDW5bCtfBdfvRWzEEz6WfbF4
KbOspmyXJDaAVuT5J6wPcmq0vRRAk6sXrHmnwHH/T7H3Si7Avyk6Rooe9gexUArhZ9O+ifIwPhEA
2ppQ7y3zMz/m5gddEF0rusMbb7uYdxtOR7FAaN+9SdLc3rZZPq8k7W16b+tW7sqH+BTw9nkSEVlo
hLQTHNweMX8JVg7zxo6bPV+zZkCZiKCumSEDjAejCrR8osFJsdpbEXIaPySG83T/pHqjVXTd15BB
oV5WQe3wT/4NEYJkabwHOUAeoKU0QJUw8cNyCshUrh61in6vDjvpBE1LacNOVH3pVJJOxpVnZxEW
rQ9RFuLznpSF2kim5tn1zqJld6sIRuuImdIwzfD2YYRERsZOiyli+KtzZEGhxy48+43zW23h1o2m
ujDl9I28ZoshPQ6RZsIwYCBQV9qT0Q+GSzz7zLYKNO1jIoYRhpvTATw8GGTtLIiBMo6yjgWxI8KJ
xhOSFkStqzADtjlvXx3cqnoYhMt14ImPIvWteKv4FtbE1O92+/HN54Ibv/ZjnGofZ6YDv3KyST+E
3/plpZle76CmuGS6kfaKo16j9p1/WVQUJYriIKzYrcXdixsNNNFDAQmvajRsXBxz/1qLYU5kcZjX
FEZEyWjo3KCT5NdUKeTPqCHqZbOMya4nenJMcxt6nGGKe8itt8Fux31qdtbEBJTfbQI/GUYS0qjN
C45d2Q1nj+AzXaLjRDeNx0PBcBzDpIzA0W/XrvE8X/fHdhq/ILa+LO81EX9GRL33rdPpAIdk8IiA
Q2Gg00f8Ok5PH38AAxfStliSkuhaTPl7ZAAZ1orcQ4naVNK7sjM3I3lwjsl/8KXBNuyHr7sEiSNu
tBDH/RG1PPo7NSpdUl/deXMlbZYpt3Z9zNpsd5ENHV69CII8/Hq4k+aXhTQu6P2dDrGcATsb4isH
4ppQdPMoW/y809otGs3+bTiEYXFI6m7Qm+xR5MCDPxA3IuoPlyLX1xSKUNq0tKi3YvYtoyt8XZPP
wS1K4rlKejYygwnUI9/V+jjv3URryqvdJckhnkiwE9aYI7z7urrSKQpL4csFXg8YvIWCh9DgzLVZ
A0iOQksqD4x5vqXQK59OWIHJLP7fBpZHpgXaDl3ZRFZgsINuS8fv2YwzldBwJioh7bYIcsxULasA
Au3AXMlgu26JSifo22G10zaq8W9KuPh1Nreia3vCCMxJiDaFj2x5nVAbgVE+z3dpPEMCFVue/qQk
SLAktG35He8T/gPV0aLuiyb6cRkXDuSPSZQGtOvu/wVk70hjiIhchfJxBS9vOwpRFU8NZlpywxlV
9WK7YuBkAI2ybdRcNdOo/EP00F+90fEy54jmaHF9RSYDgDOpS2ahUngs88xfqTzo/+sLhkt6HkgS
cxByGv7zmmM+bZKEG9lDNAz5tjAr7bB9JwhakoPeuqCTrfjvvUgGCRkYxHPT0km7zK66YSwMMXPK
UHPuFsHEfGSsx1gx8qxG2gWZGkfoLxhEwKTjvFdvW1Xyiv1R0dhmf7h5JF1eVhWJVol67gQ/Rp1z
BU0LawucPyGYs78+iFJtIpxfyFjc4msgwMS3Kos9HDbNuaSOhK/WlGwk1YOkFDxgmfhXJAuZvMud
nAsH8EoInxUcnc2dKj2AUDQ5rC1/iBMSsLfr/r8wWK66d0nT90U3RHdRt9Hk6fHwVRnoSDWDfUrp
tcSVgNTFadAnwFoxQRGQ9K/82L/ahYWLfmqOqZ5cQWB6x4HkCom4IYxwdqV+ZUxgTGNMeygNdoPg
RGRzY7yYUFKbjYKCk2dNN6o2A4qg6usnaZj7eE3W7o9fisgWjv3UUUgATOBg4m10qjVZKSUwldnN
ZF3Js+M/8aavl0IoK6Wdvq211QJDztSO/YdnY9dRFPq1OsGQGWk2xUA0GJdGcjP74Pv4At0ixQ2o
j2QggSw89kkygNlD1Sneu/SZHt2Uu4ITFcOKS1tPNgAChhvQWndgI4esYsDztLTg8uYD1xK5yBM7
r9sY7SLeHBDfHJAQu+v2YWQOb2jKF4n1PYUmMaw1hHWPioX1tLSUOpQVj1qDTCMPhyFQRc32tnH9
/lsf4qw9q+OqTMamMdnPQFptAzRvWZPr9dEtuG3KXsXOA/TCCO4WUwMoQLtnoRhxprtihtz8sOH9
j1gUELhNa8D4Op06e+BHJrcM5yFACKQJk7Eb7LbP8dfEg+T9OeL0tTkmcFMmFGJyE/3LaRuy5RFQ
xxve2jHWze+qRvpdVO47207iI7MKB6AFQVNWpXzumgBsZFeR4mueIXeg/Jmhox5JtJu6bq5gylvX
7lmZaV7rbRLO1ATsOvgpVhJTRY+ruMqmMmUeM0W8xEX1xqomr27ZwatV0bL+iPf5ycUd8c8JUb1p
NIAQJTUKweleaDqWMVRyCxgNnyAqOJPooq1nkfBQMwDZQAXKJM2Z9yxMbOPNNBddPZNj4aPXG/BV
b1RjXUivdty38U8JBWlxyC7FoflxeUQXp5aek4qkpCpQwa4t4oQslmkMHszTi5sFa4H3vwRL6qFc
SrBZyTwjBHBH76kH9PtAmXNT7P67QUNg70jqhFWZU9mbPFq4PIntljO3+iZCSg9H4eVRa7vx3c02
j06X26EBOSAWCXcmPDujulIPW1QOzoSHvGdHMosphXKfMzS5hHoLgDm0dojwffXgwPcJmOXF12N0
2It5lhaiOOFJ9+OICCHdNy5NsDANqIlZW/ZHCHvnVCsVhPlz6q2wTOwJCKprEnCLBn+MboFjuIT5
/YzizDiuPlROkv8ZGv4UsaAXkW9aG6ox7eGerInW5BcttUMcQ12yMFq8f62x2pq2q3XfnMPUepOe
adDU9kUEApvWvYosg+oNcGVbKfPHKV+Pn7AIiRJo5dlDbsJ0T063RZw2Cfsij/FmgXC4fgh4+Q6C
e5lP/L4yd95qWBr3/PeKiPAiSPyd1Cu1L6OfsLFbERMK19ek/puPgXq36p8v9l5Tc/78K6lwlEMH
A0P3/GiKWiRzv12f04Ao6AV5Wgm+A2QhfZH4JQqFFqU+qmHRPHFlN3RSu3iZZEaH/G3k7oY6s/dH
+y82Mv3/nq4n4woEjE1jztilQnYfabvTc0waW4NaQXnbZHSSOubqAfVxv3HVNWwqZBMHl86nYuh0
rofbz2A+OeYVdGg0CrchoVRZdosqD6S3jNR7g4Z1yRi8pz+VPd6KTEPAd94b6Q4eZWedoDhdX0wu
7XG+1Ebj7aha1j7bz07S8eB5aqDkLmi/XMHwGkZmtFHzTvaDUg0+FO4JJKLdnZNXCMIstPbWcvrj
SEsRBY06JCksPQ3rG2JrN7HnzViXum4VNUlyXIP1W5p5E/lAx6ni4K2Ps2IBebKsA9yjuT/+OgO8
EcP6MBqa6695tfj///nGMyxojizUiq88G9c0OiRpT+ELd01EkkhE80bMUVlIeF0J83I7mMzD2jLl
W5RbcVzWRabSOjsRHmYT0S1ZDGbHJFKZxfs3+xsM7TFkZDtMXP9jUzkk6qhADNro5SW6MOmISaGx
2Z7Uer7LPISOd04ZsAotcLNK4nf5PdBLmyqVOuwsJpf4KGKxnGRCmNJfWheCT3zP8IcPgqyLl5yb
jlaKwPk7VzGHLKOkP0VHaIviRXF96q6ro2ARaGGWj3xK49jheNhOTjhhbj8GYv7j/I6jtuZ3zaVv
psXiHBMf28wvUlfIusy1WuJq1wawBvS99EKdIbwitT65LN+wGu3vljr+2nQmQcesmgGxAGH0qvxT
dzImQCeezNpNyVRKlcHo277Rb1P1frXcMGZa1+A+Y1yi8+F/xelkC9c/UZIAD0wf5l3X8Uv9mEtN
dnILqZQejwz0w9RV7U1DYyoYp+5vcdyxO1DAgaFACIYa/s5/ews2z8Y0CKuzNWlmJnbUqI6QqDd/
8BJj0TyATb1Fuq/P294CvOSqWL3hLIew8XEkVrwmHpuXAlByakAjXHruXYrPPc6yebux//X/rvq5
1tJzAqkpSX+pl9RoXaR/eJgc+xuMlVg9OBfO7WoXc52a/Sqe7KzxcT17VQTYfHtiNLzDdRtrNCeP
Yb37ao0MH4XAOXMMwyJaWEnabEDHb8d2nYeqYxKTTY2wqeWyHyOwRQVwxlhxLwlBtRUr9HkfRlBi
rjV+yUNeQrk3PTym8UFVMXngEWZZPhFeD90uiig7b2l4EJ89sDCXHeng/Fvo+QgEliFyhNDX1X62
sO/CtxuInA6745K9r6nMQOCLqlf01EdABU/7/E2qKtUI0+luvl75GTaKszMWtAYpKQkhmDHFOnpn
9Dd4uhe97mE57vTHEMa+4vKRVmdUmIjHpYjm2o4Mu/zDJdGkFU34Y2T/ukOCQ9+wQ3V+JpbQkj53
a0WeixI1fi5oD88yMdX5CIabHi850j9A1GhJCFmr/Ooh/EVBcgaBEcqU3AXQRIcKi/g4T5wdzu1T
n+oxEYaLf/3/Xq7ZrJLWHiaLibMNUBBid6vFqx4HqVn5G6NSdA388zSm3lWGW/PTxCitjoHhkadB
YDiSGTjZ5iBx96jQTkMHwD1aS4LzzunWNcrTOlVe2KQBwWXqG3xgQucxjQzBVeukTbpgOmxH54Cu
EsKxd18ebOXdcC8NtJ4WWG+iA6H/sOZZIKwxIl2tz2+1SMPgCj4s2i1EET5HTZQLTUyaNgHeM1t3
JGotzNFeXzSHt1f5/+wk0Wdfl+lBa0QZ2AAFeEeQwv1Ah2gMF9mIwKq2LcUWejVh3w6oO++2k97K
Zdz3NArdrPBMBvJW9x8bgFQ35N+j+nrBTpOnZe+FqVWpKSpuNI6mMg/S8ctEbMOlGfEge4ZPSDBe
nzFPVtgR9yRneD9WIggm59zOJmbcKT+MJItUOeJ/AnQwQVYdV70AMV5Y7V7LLZroEOMLf61R7U+4
0jRrq4aAHHcjMge/TZp1gw0lO6bN76+NSlb2rZQfe3cSFl3EHHiqfXKoTdW/QVbabz4UfHhaTCDK
Ev4HNDI7g9G9r0rcZvzooQQnX3fGl2oQdkP0kLd4J66tGBFwsd9KIrmi3DKKuG5XH6tP+QIu1GGw
RHpACn/2P6AHsJmn4KgCpA45QyR29pnmLJZpTwSJkOCAHhjvlE7qQppNl5oKCPOYALsfAjgQ48bI
o82CGgmpOdnUzSR2I2HGKFw4Ihg/beLm/a3jgV1oyikavFnt5Thj/qs8nCzEDhizsPKuY+jFTOIg
FhC3Y7USQ4+3lQaJFtnfTE5jmiVHWKMjl1lJHUKtgxtqVYXlmLNzuUeNqeyLSlb2pNvkIlXYzhQy
YTXkkwHKy03UMazfdqN7KlW8mH3YswNgzbkbuTvnR9Km1p7KFE+aZkgs1Ux2ad0QIAmM3Ijh/aw+
Psniq/nung+F2A2W7nG2f8BG8rBklI9vuZBv8GLo+dFUiKNqhXfF4qRRrUp2tkfAs81cytoVSyyM
umadbWTtyOZ+Vg+0DV2ANxg26xD5rEr+IiXtBQaoz2ilOBrcoa3IAL8lLjrbDWQCVMkfPWbP6vAy
JM3xV6ljor1qVzwvqLTFJEbnufvC0cOAMA4PMcaa7ZgnvS4zR3xD0aUYanoFrgcIRDiiy0PS4I2l
RwkVJ6AFThDSyMm3L7ZCPEq6QIhMsoPdCvQouxDjdDb6uV68gqo2AFQTu5VUDcFf2s8OHEwdb4uv
ZHJ8p2wtdP7/KPryV5Uprsnk+Hm16/OVo+1tjUFMuM+cw5FR8N5vJVKdkBCOSNTt7jXaLH8AqHf/
CfX/X5NpQ+mDsf5no7G7BLBAOXwDJ0ykPfSWiEkqO/n/b/CRJX8xfXb9CosHhA8r2goCCrhy7cwk
vXYDkruO/cwdL9AMlrrV+uABLJD9J0JpIyZ7izSpvjuIhnzEmU8ho1hcSS5F5AIJHijP3D/De6fg
4yjLe6P7E/7i7iZJ5rrRiUowpoMJGDIAVP0+9OHrrsqvRm/4cldncNkevlXlzcAoeB/ecNhhiGDC
e47exNSnTQak5uSU1V5tZhb2jCEuMFFFNlzgOHr/V7CFAj5YofkjVwTuupVgOZoPRmieNWpBgD58
SPj9f3SWdA/rmsgQXHp6yLQJJGdfyI7G6G9rwUKQRexCVcXyfe+J3PuZr0rMGHNrNUCUmePRMIwI
uxstu132amDWuxj8jSwC3pm1+u+o/LlXlhI9NqSwQstnqyRuJcAeO9wUCyFam2Fd3zmkZXupkWRj
3U61VHHor4aD3bZeIJ78wT5pCLKR7FdhL2rYnIEf/wyexdl85d8ATsBu6fisx0LBNzw63zfttkBZ
Oj8GE5+CoHCWKduw0TN8DBJTMB/E6doE2WAGZWMeAsjXWBnLFpWrRxlynU/qVUkJrf5wVQ+Mfkx8
ZrAnw8odR7xfJU3X42C05/QBEyzKzA5+P45dxNWAwpYGg5cSn3LkWqapya457zRmvVBlVHsAInyK
pUBfs9rfNTgD32yxr9kL6cjK0UR2MI2tRuNILoG5LoussfzTGjgRmgizCXjHr/2mWHlztNVv0L20
xb8c46AQCNhU3K5rWubPqJ7Eorhz9DKbVGALqsW2DOuOr4YraJNmYMX1ueqEEND05UZ6o0Q/dIJN
fzM9W/ekSvASRQcgNgj3S60nOiWB6jDGQYui7M3xusPn7w2642vUXh0GCJF5tKv6vrhrGpi2wcXv
WZ1DvexURkr1kNVUwoUEo5vtW8p1LrgspGGX9yGd56msCKU5U7ip88avHH9p5bGdmSTzB9Oj1yEk
QuHeuNGs/xSLcXq2guwruxT+9SBqaCcgL1trT/VgEIknNJ1oXH+NI/l3wv9OAn2ASBEFRwWJVOTL
/Qe0XOWtohih4YBhynFHFgWmm8KeIsxOIcZ/vWyFlR3xBXdZT/G/dd2pWR1KzKGGuY3lOR4yzDh6
t27hO9efYZzu1shO1AQP6dO3S4yHgJhUsPa01RYL272rFE2Bn65UexXFujuLEBs4ULJTCbADQ++0
yYXyen6dCraxW4sbcUofwmxoHn5cV7SBHQs6g7opX/aNqDryP13Tk4TS6Fb+HAwL0hHazxOZ/q+i
negX2yxJ1pakdKSrLlOHvsTH9nsCeESLJ7RVnbBOu7Xmz5Je44DKjsjkvKQ+nw38Fnrs40iyxZyS
QHQlY5m3mo1/oqRdAzlKQVg7iN57340HuKkJIpIGRMg8h4semE61yWVIXBr/hsEsAXlGf4MHSTA8
bh7Hn9knb7jnxRhZeqaaRpwFQ5R3kub1sx/dyWFolbOq+QZwuxNkUHm6/VHhdYMVN2HtnizMrHc+
AgZOmmUqVuil+yYFdbmeWrNABWy1YnYVLXcMgQzSecTz8PcSCFEkCU0UEU79tPp6tM/sMtdF5g2z
CuOuwOp4tYBTj8CN9maTZ4iTMZZVN3wbNE+YTw4evPR/xdi5+lxeFdRED8sY0Ygjgh1fxcnPDKrA
epCgRINKWx/T8Ovd498YOrMvh/+kIP/Dm50+1vcThLiPWBVAArCHCCcsXdA/j3w3fcbGsVGm4XRZ
ac4REOGZpv91VEfzsauE1JuN95a90/qFgufvixGlG58HpJ+/yxYgvjXzhIWQAA3eJH0r1nR6+yLz
weL2Khx4Caqqnd3Idf+rwqUQ7a1ZJWEHByLQruvCBiSuL1pxMNWInssdgIM2sI/mY67+pc1PtTAa
xly9pE1dP0S32w+UiBxZpFoM84RssHbOiRFvEQJMmr7AJO9vTy81x5LWo1/lTlVg2V9zRpURbR/l
L8ChYR2n5zdeNPPjPXPayEW1ygvlMwxoPYINP0KZC3Cid12OaDstYQ9+rPGI98cmpaqRLYb0pmPJ
TFrKGAH36Eq6Vqe5Fibj2BWuXUfGxUdEFw+HUavGkcNlFoLIigCjHDFeOWEV+9zyhDLO2wo1u5Yn
YvxGYRaLeDl1rfv72+kMf48dks1HORI6l0fco80NCVsYbRMcBV85Keidr4Nr9j9Ay/TNtvVOh2WF
4Rhx/8lylAl+gEN008BeXPtpK00P7krFGpW6fdctxsgXQCQeeUWBHXagXr6T6JjAqHmqLGpiPqtI
pRYPfySDCXCQRf4HZwesGD/nT/+KCj6n8cavoVI8dMV9xUBe7dXMJFMe83cfsvEa0HPITLTh1JbP
UUMdskLWrTf1bkARPvsXoFIFm6LEyD/8Uem2w7iONFZoQcPjFRuCNPh78HkGTqBm7sEpOR8lLgM6
z5oF8Fr9s5Ch54se4xBdutzDIKjPTAGUZnOXBC1ovo/8F4RqLFm2RJ99jfJgQJ2L4qVcxvCcTjxv
C1juqJ23Jxq9rDXw21E7EKmE229wQqNDzs70fbem1Z+T+QY53qWenFViXL8okKkSFSDcI8EUos5x
uHhKrKjY2W/6RYgN70Tap9x7ZaHyHbgAa67t6HFdcjIa14Rprk582J+qV7sCu45n4gOInTwIMB0+
Yq/4bvUtfYzRrRMqSUlLKSLb1jdYN6xncF/MKsFU66pK9dc66BeOisjJPfVyx9RNFcR8H9mixNWm
L3y6s92OuBSnw3kaZ2808/8rXQuriIk0UqnUceg2QqrUabpeeFzUYV+UtkNtPnt8PPT1VkuanoOx
NmqL/lrB8dor/5U6q4Fevv+c52UHcrAValMnKPnoxxb15W7tbmWUhWmC9sNmuX5UcNnqKeFA0O7y
EnhdGnL8LrPGJ43fY1FCr+efjaN/VZXMxO4lsh3opucWH7zaVmvprMu3LymfS9xA3p5LdeDpXg7B
Mbil8hfojQwfQrhQV4dU74fsgVRthnb2EJJqxKFWq9Wja6CLbPJI1IsIqKsxdN+p1Q3SwywSw4mZ
bTLUKyHuSuftvjCrfzGbP8/b2AHUMB+3kfLVxQ+Jn1JikKEgYRCgolHfrKn+Mx7p2r7Q8yXrHAeM
oXe11RgdGZCjNGIftbDCnhfbw1DnTz6VLBfX9ltPUFlw/DpFq/m6/RbfpDie0FUOYrRhuof4RvCs
YFgqFtwm9KbPq/Z5MfPgoWdj3v3KY+ktb8TRKQPfh45xh/Y/leVsRGz5d8+1XRlio+sKIM8XWfQB
wHcU1J0QkAJX5/VmEk7CagYOfhQuuIwsrmUCjh5Qw/xvaaG0VKFEHVaMhpUUxlTUDBEy3rIEsxFb
m+QjJJRu5jMtrexuky/RUnwaGusMHDcHuV4KWF6cNzDi8gXyv7lJjqRRzf2oz6v8H8R791oVMsbs
s20GbrRzSKDci8NhoEI++8BHyGxz/4Sb3SpF5Mav/Du4Hx7+jiRjuZdenl/GtjxRHchQb85vK/Ij
Fp+ZsRGWV7bOIzsi2vjwf8IK09mCY5qnlVrSUupA3RkhkV+9Y+3Y3MZAjj/+MX8kiTEZ3Umolo8o
330ukRtOeFtdDKA/XMFdofd2oPiocIjts6TkJQqQR5zXz5K/UbI3r9+0M8jbSalT+g/JSoIncncB
qssTDT8GnYjGQe42vOOri/7kSYdSj9U8kqLhEkact4JHaPGWGPYEdTqrBgdCziYf7wC8Wa1QddP9
KU+Ig7TqMtcdMaqJMLHjp2l4ou1S6DDIoe4mfVVH14NTpOkorFwKxZNn4rWip6bCHW0jXMzTO5Qx
+Kx9oIXGwgPgKqJPgOaASEYXVUQGIVGqkTXvXhsldKxz+VtyJWUk1U5HIEhObZM9OnslYq1Ll/pH
VLEjkAQGUh/FLTZVWsVMZfOkjGBvWREnEgGVmlG9QDN+FtgaAQVf+a1e128/xX+UzUs1N7sUgyuZ
epidi85FIqaorWB1ROWimZFyqLbW/sUVrsqaJprXOa0C3e9VtJXJQZ992NTN5hBHZZk5BNYgqEfd
yFF3DySROP/JMEpMGfi11w/RGEtn2x9QsPQNRVZ+y9ze8Z1LFz4LdwDkds0UxJZ1LO4b6et01cuT
bjH/z7GGoXZ5tCUGVf3dNtaBRaQC31VQXUwISh/UZnq+36v/3dRtFOFkeP/vlua1zKlWkeqI2jW4
h2+ILRr2MXGyYp9VoRbE1g6dCCSFFRle3+dLl+3dw+mcYJCBpgxtszGjrVHAfzMDO2hxP1inVVQG
2yMxqMHBT5tZ97FaBtQ8uJR2a1nM5/saZu0i0n0AGSVZeYn5OVFCNTWlftYtEspX/RJBbkhD6h2d
srf4iaSCQW6TBByixv7CbPpdQjlqmK7bO67e+uejcHVTpZI+gqUhOMkyFIf7i73yUKq0YMSOtu+2
z/lvypyXPr3Mwqg/ykQ3n3R630ZM1Y+dlqSmCG8tceMrihrTXNX5KT9nJRZpsq+lFWTX2eQsMscp
fxGHQk19Zz9T38vL0NNdMqAu7WqcgBJvBOeGIJX3qKhoscV5Q4oGgqMS8JqS2reFAQTGZXq+leNk
RlwTzVTM2ZFX0BftIUTDCodJrkGEZOO7cCNALS0f8GxuvE3tFKldlTNlLAxv8O97hJubdUuaJm5u
rdqbGk/QS8ZuQRHAR9jdXF4BGyQujhFDJ1FnnuPZcIP7h/KnmoPTTNfzVLVAYClD8bZy6ZPfwGj4
3PJtuhWupFFQkJcgbAo0eq8UfUQ/mAT+50jLpsgIgfr4afPnbS4aDp95tKNUk2ukh6ygD8fII0Br
Syo/IMI/chLGORC86xoDYdZZBRnuLCRQDgtXSu63v4QrTAq1HOSvhQkzk8UN8X18YBG70rVVdsSh
BNI3fZVD6wFt08uLCX/gt4uk/p0W3wAvu4OBkoVAiEnnHcJcEBBIneRyWXuYXHR8emxWL68kC8oW
CKLJyTbfIZDWusLECjcdiwoEw4ljIE2YUos/VqQUNHNDK7auw8Jf/CxzCFiDnezzt3qJOGfBMuzJ
WyaPlY9FR2wok+8rca4rd70vrYA1fKnH24nz3KpzT7IAShUXYptvUU+eDo2QSTShz+iu3886PI/D
aLPDFtMq/Tn9v+eOaf3q2dtQkRIy3/YfwTk7yG2QyB588Fa57zn2uTQYuIh7NSC8v4eg+KZd3Z0s
JEUJYq2t9OW86wHhIUANTWFGvczE407f0ctea2cL4RBnwaPG/K2UAqjW+86Kz0r7JB9Ct1QRa4vS
MkuhOa9wuk4Tq9a27fYec0koSWrtsUYHqYnASf105Y1qv3ytoTADV06gNZ1cYx1EueBrLlii62/Q
pb7WleKoepqzWjOkHcqYvNPsaURCY9AmMmIc/RqUGZSOHvYA4AKy8fjXazeXTreLOev6gQEctgb6
4BidNoG1lWvXx1k8GgMHHwu12wAdHKcOH3e0CzVUJFYqsKbO3q0vMhFpNTgP0x+1x/Vj+kLgBZsd
fmsnRMeNRXVO7bPAsyzWoEW7MtUspMPPMWW5Evrb8AkjBjIlX2rOCm4Y+dDXjKsQYULzzx4PCZtq
RVeTavGP1EQ92oY0LN3goQM/eMGIpGkrgyoaurapS+2xdiPFQlQSvcr7TMcq5DB4pfBHQL7AULx3
FXELZGSWxHvBqqcr8FQV1RzIrY3q+VMup/qPX+hsaQ+5hx5f2NDwFW9sZX8MlOuSr/ZN8Fcs3/6V
L4b2f5pc2kGni/TE+I/7IXXJId/VKdv9IxW8Tl0lVc3LKHQ26LPSCPCv2YuFDPrg6itSTV9NfRLX
bdQFIBKP6ox6LXFwTUXSn2BE4NEYZk2f2yW64j7pHky2lmbOwC7ixFBXqOo370Pv3Zz72qGypIgn
1hcZ1oTmFNkjKH9+z9gWXG293ejVXObYAc4OSosF0EWf7Gt14ij0E92zbuRYZgloGq/oFr2Pc7tX
FvsXarT1caVLBnfKMx+UHxdOwDo5/3ynSw4AN1LJDrZbAbEAZcBP3HXmuhg7mUzTPXz82VOY2TgX
laS+RlMnXAKPrFewrGcoUjdsyxyYd9ixLBqJct4WplEhMz1+fe8ujpqfxnUt3xBGP+lhv56e9kwT
t75zh/nkWWmA0f7jpFW8pBp9nfY+ojyiQdx8veL2IshpcdqFR0zNK4gI0A8ascnygBZAPJl3qssn
etY7wmwT5QYBzOLpLZLkkMcl5rN8/kTfVunkKKMwk6STMnRoDO+bM9GEUimOzij7TCKzu93GS8k6
5oa35a4Jnr5WbDagQ+e6cNkh0eOS9ZcRy9qsftXSEIT6Q6ElLoNc5YaG7iJrJu1KwMqCzY336rls
OhKlwV8wpDnYkooaKxsrnV99DnL45EJAHBCDJ+56D+fUUoIXmNObz1JdCqCLkWDBIjBLtOWWNv+H
HHQweGU5ecEF+K5pYy7zY6EfDXJEFHiKEBZvMB7yLVr1lUgHoL7k23xL/xkuqCU05ay1edkTnCSA
grmM89+URDeHyW8VPhQut/iLNxGIX3fUlTHZfqXneFrAkd8PXGIqw4RRag5KTm7dkLOKbcB+LkR/
nT4bzGRuV48y7l3+o97AeSm1gmNrGDKwMb9I2CUO9BqQasS4oPq7pbfsbhFbiGfC3on627wOT5Kc
g7S+muhfFNfAAnrO5vTB5Q7Bah9k+xID0xPQj2lKJvr5I+WXCbhiUDJlUJ1Vr88MAapW2ApnCy5i
V6CRK+N8yjuWKBXHbZ7oj15CklmsuhMEqURTjCJ2sGDjG+xFHRQge++b4KPQ2x6T09MPfLJ30DJi
nyDkZFdfYRrKxhUJa8wHSIqZ0yrgaU0ljGOf0PDoa03U93DPjIM0XgJlZDOXSC3x4xFailpY2Kwa
KPRTzTwRx+epdqeuRFN63DSg6Z/C6wxrrM5I5UDj4O3Dwn0BtNLl77LQ9Y8ISQm9ot9qgHTBmTQ2
4jXscq9vWIIhO8c7BqinF+j0ZFR1ibB1jqAhOF4dSv4Fjgi5KJROmU5R+4Mj92/4LyCPNo/Elk95
uQbpxVRxdyFVtRKv7ayvexdfK9PzWN/s+376YKqKgHjmpdR5f3OXPGqSgwS+y6M5BMM0vA/1YR7o
o4dMXqHZvNEJTlIwhCvES9eOQT7KuBv7OEFYfmnvriqyl1hUH3xrQT/ybzlH5Vqe/SC3I5qZsfV3
ussbjeQEN0cuxGdNUKeywloQrbB27LOoMQwSM6X5vi8+9kGSLaIr2ZqNQAV6gazGOxOn+Uzcmczj
0IspziHqKqagwLweoA0NlMku/r8BetIsR946DBh/Fq4o7AHISFo+6RohL67mm84gg2pKxW4vUiy5
r6Sb94HkO2r5ojPFg7J9ynfQOR2zcYPRB40cpj5Ve+1UDOKvEgK/b4pXh8LvTt6mFHB/VZuIi0Hp
zVgsCd2X0Q/qq+0eKwoJsWj+92GPVqzATr13zqRm5h53lSQd0j3zztkuEYRRMPzsvwJlSrCIZzMs
tLaQOwvGRYpHaQUNd8zbFHHgAWdqCmRTJyPEwEFeo2orpdA7F270jEbqIUO7aszliA7g/fmKDij+
wE4RxElPWwisENrWmny3+yrUF4H6HkjZVGHowlbxYdwXqQ5R0I84/bXemIiJ/2O3Z9rybuKEDIJu
Q1+CSs1Z6afZEw8LQ06LFEELydcrAihLf+OmHcl9GoggXkBDvCeUOiHwnYlAgbKCqtAojmm9rpNQ
ZxE4OfmPiwDL2Um+yxR3qaxpDUGypJleX3/GKwkZyxvaCV/NKRsmvLkMP+XuT/riTWZTjMumYtaQ
gY8Ak7OrQqbW+cTnLPdIjoZiLys4CPIbpj5XNfhbxdhyKIxnAG0yBINCUOw2TFE4rmO6pBt7a5Ic
V5UMY/1DSVVHeNPD8klZZoIDBCPkckCctLVRd9Hi2l/crjVHAfYTzDN54Co81bQEio44bNOKnj6l
wwy6+4XAzAoqC5sdzKzeRMAU8sv719YES7iK5eLsoKO+wcZEup4evhODoDrK+MGu/2pt9n345SEn
VV6F8c+bFDFzHpb/ylQ0HMt5BqbiEZIwfWtn7HT1dzx4KMXSdmJPdaYqXFMZW5mfgnprzX5DvLVN
9F8KKMPWwMqfGnLdiSTqL+fddkx7ijsXyr2Tubona0WKqWnla26G6kssQmZiPdP9RBp72ZkiMFxp
/3jpVogjfY6phlVFMC33xoO4A+4OP+w037BO4QlqHHpg7yWT36r36g1tQmA1R51hJGo9T+cqyy2f
GiVMF63eI0ncwUI+0v4Ou72kgSTHIIPde9AVJQW2fMxtWJqNjB0XNDmaXa30uqUi16U0HV8+lGh6
jcAZ+Z3IkazfkfIG51wa1LD0i1lOnJqSSSTMtlpK/C4+GqscTXm+k70ykUD6AE2mVMmoGfjcqrom
uipAyhmRrxUA8cdtNfQjXGmjT96HsQcirSxdsjaNluOTnMPmiMpmkw0+eWSKvaljyQnRggZ1rTTu
CQ+D5Boo3u+1d/aW73p4QqdNlEp3+dRZ6QVvO5lAcPhd+MdiX3sMDWpxAJcUHvtuC8pDjdWwrs7Y
AElW8Yf4w8dgasGY9QOYn6Wlx1OWXJwvFqWDqnjHuot2iaR5EL6fhMgVQzdRAREFhLm/kv5qNApe
s9r3TVvaluoUEtXI5P8L2xHokDJVC5iPt3ZP9awsBgYwPqLZ9sTq55mzcwlw9ubu/yfYYNSQYuiz
WwHYdVc4wRqkip4USoJ4sfAIsv22WDYH9HGtHaCMAWKByr2pVoEAJSIYm+MOPQlEoQ6val6v1Cnu
fchENHATI58Qy88xWGcVn4bvWzcHAh8In7ALx1lfwHPQJ1HlCnUdqhArAO1mxX/VMvSQd6LdnLDY
DuvV8f+LhjYJbPLYHGQIRJokyEUAlka4BkJzOfP61MSSvoQj+D8Yp5xED5BE0EugWGldJSVmY+wF
ty8SmfWRlPznaNCX2H7zR6YJZFUROK0rW5uIOULIPhtVFPKJTxHnPS7H07niRzd2//XMTXh+pgpK
aBvti0SYA35tM4MBEHHO+U6Lvt/p2wSUvOYvw1S05yN54mUPUdL14GCNs0bXjjDg7OlVoSB+zQtH
tbaKMiVlSKTDmwJ/PmJ7zA7N5KZrd2JpvQaJ6krsQyJHW0TvTwNdxaDPPrpplbvIHQzWm2pOicC/
QcrOmVNVkeI9MKyCWNQpSnCbBl++U4IEjtGmlwb5+cQtND++ulilDfSqLO1wraKsFCn7+mDtmy7h
FzdrdmZlb406M9xFaoKIKkuA0YWlx8akha+YapjxX0Ysf9EBWbMqHi/Fx+dBz5P0/2ifg7ciNygp
c/626C3hVJOCgnPPdd5m43viCyVgNiU8up3TbyeDXcQkqMPDqM6b0SQUnc8eCY/FXAEWOvHy9oIv
CSWn0ftR2/Kwn4CBsw7d/f4BVrAwdKE4BIhIPGRXvoY4cwylgrJQdCOs+8zi4BUoLYzSz0mbCDn5
9WG54suooAq+YatMBfjTCunfPfP1IQ5xRcXxJQtHr8Tmj/zAkNvt/3EYanyuS/a100nEzdEmit3J
QyB57nrOdH3nWV8qFS80Hcw3WW46BIBeMVgVDyC5y2kJ1Hl0GqETHjXMMnffr+K3WlvAO88WLEMN
hv79T/p0ZRUW2xupLkOYKMwgkTw16dRT58I0exujcJht/332nz1DwMqTKMJm8TdZmwlSKXrHFkWk
0IDY8AGD9A146bL1LKVT7iPbhK8kYZpHSDTd8RG2weKvSf2Ko52CImdySvqtBa5t1LX8A2HU76QO
JRNS/8mYnjAcw1iU1E2pR0b4E8d8by98mnajO4w1r8ylEu2rCQNZG/AuppSgsbfOXBBzCP3dqNAK
X4fIfBqkylxE6xpT6XtnGyRqNYrAOHsIiXbqqIawG4awpzNRfFEZ5kI4Fnx9Oeip/GUDmYPDUX/l
R0mWKzrisFIiQCsfvSAeOymegl71VBQfbu+WT8q36DVxoCLs3Ut8NjRfeTI8CEGBVXZGh4aFhWF/
7zqGcS7rC/oq1jwVOeQcY7kulZRTFqnLFISAx5Ysc2Pvm7eFaOoAH7u91sN47PQT22EvFeBS+pFS
OTiJnFvgezNNG0bLBEcUXuw5Vk7q4bS5bQ4Jc6q87jbBc9NChODJyznOwrU1RKH+YZTBWQrhfVs1
zYSwFk5Q4ZZfeLDVRRA7oIebW0ZnW6/PUd8BuLgJ50KesjbZVH/CJ17lVL4acAmf81bG0YabmWWV
UZCipUeblL4Tasr5HmvQ6wYegxFWOCGKrnFF0moUMikFm2MfYXl8bq2bFH2MokJoLWK1KVwvBuu6
81z+eITpzpFU/l/jU+Yfqy5N2E/6ku4Mr8TyAqiPUIE1wNB8vlm4GjiU8l+1JqXif1jQv28LygCx
pj4ssDwEeJDl7qL+F6hW5PjIKGDUwH7wELfxwy/E7WHB9kiHIHgH5q0Qw5FTe5rxs7zC8ECRRYBH
TUrSNHnrCXRNc1paxGdmsRg+xpsp8jJJWT5ciGa1oqp3YKlwrHlUxd1naaESQ9WdqXKF42uYzAKd
Ft7WZl1EeaWPv6hLV7/eOVj/DnmD6N3BA3IYdh46d4fV3x8+kCv0s8Rn5mnQeXIVzqXytQDt0l21
SdwVCmizs4DW9c7nd+528trGkiPAyRzJAI/fCdmiFTrA0lXRkn+skRhW0N7r2Mn9wtG/mQchNXck
cuKqfmuLDUWxU29Ps/ZLxMvGchAimjoia/9MPTDg6mKoi7QJLviSLG1wrsvya8YYgDCqQmm9u+90
S6RRYmvFQrV5JNjrHPO5qFjjEQA3XA39mN/AYFHaCBAVYNytMxfUtI/161bp5TBmnanNdArEA1A5
dxvqq9MWEB8EiZUp4/RmR1r5d9THXcE4WsV0tAF2htjZlXZhtXxyM5CeNRt27Pf6vrUq4/jP6w5G
THJ6WF7jyNF50wArF3wvh/0svAPCYEUdgWzThc8RKLvbeYdm8zkD75FqCEmKQzJL2uvWcGwuf9Xn
pdi1ConUhnPB/u1/NaGBP/hTEDx4IXpws7DxxZ0duEIOs0wdu8T20X+h0qWEFs6yHsfG3AHaBo3L
0UNtEQ3qqqdf4cCaC+qmmRX5XVgRHj3rznkpP3JtOco7kOKw24grvxgdepsdzHSC8Gv8NQ0pm0OC
oqep9u7CP5fvGI4wA46nM0HTnfZQo424TYDuy3amIDo7L/dsXrpvAyetuyF6VXvL4ex8YgTpsnWP
PCuA6jRf/jDRk5ek9z1Ho7Rs3z1Zx1CF9exBOoZjVuF2lR35jjpEqFUdvIzgRl01RN/3mtNakGGx
ioIl0oQEJ7wdBM+eDtGg/7VOgxf7yk9qIDDAGKsiM9vDGsRfyQHLfWiUimY+GnGawnlroNafFVQK
QKkfXdFpY4jTfCubhqLBbO7j4YFYhc4stTTjHO3d87NzS0bhJxxVKvLsssGHu9hh8RuVb++wMjKJ
qUqWyp8jOrhJSQZmqr0GoqO4Q8MwpscAXrW0abNUL392jDAE/aINMme1lwBSwH3mB5A7OBHvHwQI
tN0wl+jx496Gq1/BlAnmQu2YriXcbjSEqE6qQ9h0uDrRv+QV4pwqCdpeqyanx2yba6mQBTbKU1KA
H4kF8/r/It4XNMJ1VpCBGvXcpDqpECvN/e29HVTUeWMPVP82ArKJHHwojpyBMX0R9zF66I4KnD6v
TMfB4AwjffEOa+ZEvG6l4LSLzRWY+46XaXfHHSoNuCg8UPjFMtkC6blDIvmHMjvL6OM0nzJymvpv
VpS+UW4LkQ/0m1kQMD7EKTUN7YFTgpp2+BYpAbfs7Nk1HL2kRaDNt6v8of9LoMoTgTLA/7N49jEI
FTEji8EHs184SYHPmCdTV0ukZuI+CWogNse5GVjRzni80PO2/SmdKLdYfFj89ywOG/bVPlYWxIAH
8sF6+NWXiHrZ+MCYqS9wsqZg4Muh1iaruGYQerdm4U30YuUtgR822BTRZLJDFBUjB8CYkViZ6omA
Dp3Bfuu8n3FwOSGbYWWO+RJxum1gDDydN/HxGXR/rDQTWXjvQrPCcPDQQVsiOsmEl8cWVJiVQxgP
dqb3D0sboyilCIpH4LUOcIlfI9FNwcEPp9eUJnXV4GVzGUPmhC/qhqHH/xspLMnlxqrpQwDBrXeF
F7oNcC/4mbM71zgMSTzmCvM1jZ/8w/5Kbw/P3ZBS4/x3WnyeF9ukAdhUpSPapIDVKbRSRYLc3jzo
JZGqYhTH7cuAW/wxlw3y762Rj2JOyBrUkfvBAmgJDsRQ3TGjQ5Eetu+FseuQTBCQeXVB+rHzip1/
tWZKaMceYWf4NLiIWZLILLqnrOVQftWsqF71Rjpq5I1lzyvnA2lRzrpBQOo85N5A6kyxMXc4M+lF
l04VT8VVjybraelHur0FgnHQ7rv6FzhyEY7ljhrZxRMs7i7mhVK4clL0R/tVi+rmZrNI4uA3wtsE
UxXCRfQYO5N5yelC2Bv9ERZj8iQRweJokKbBEQJ/hTBVRrA3Z8kfQ/VYXJz6VSnfZtz+BhVgNo/C
ORL6ENTejPTJHdFkK/FxIpKjmjRFqEW69HFBeTkUone0w9X+iyDoKUaljNgqYhtiguu695tupdmq
D+Yae+luNHlxbXJiwxCQ8zGze7p+2FnyM7WmKXviFbTF7Mo4ZSYDfvDWEjAXTJfukKpeSGO4S/Ex
jCgVx9GPpST8Jv1mGwFU0LTkRyGhZyCjJbxhI0RG+Q+Ea5KBLWW0u+RfPXRqM9ttwGSbpwwU9f/B
dqqR+oHe4HN4yCyf/bAyctW8YPr/g2s/EH2TPfGnE1BKPytN7DVDL0DQB5Jb0cnmHJ979SimaiS1
4e1kXs8L2f8rNhiB2HR75lV8QWjEVrdk0FTr3ZVlPfv/uTCf3XaaBaTL7ycrMCeTfZlHfYPnrkkF
YPTqQpOXpbFUO5T3nhy7mQxMHLjDqfbkh+zOICvg9zKMYLQAc1gbqVJG7uj4EC/7IryJDtBr3+ja
kiLEj+0OUqhlsKYTjXEPBKccaBsrdFdbDmdQD9vcmycBBn+ICJ7Ds2EFM6KJyhmhtBJZm/o4VAyv
lrHU6epq7Qs9m90tCN96X/ipZfuht2Y3QyQEAkp04mH+7u33+yEhzp/OO5dwMGc9rI94SJPRHj5J
KvVhFIgBaUIMC+oU9Hy8oNC1EOXQ+EUrfFfB7dQYYhRJTIjtZhyY1RsSHTpNHqsa53jCUihiu8sK
QI4h6LocUoabRfykZFUh0lqMoDvsSUz/9yYFblpVtpNl5A8txVcG6LCsOPHEB1t70XPXwpIlS177
UfrzL3gum96grAaOLjPFECAh0YOP+QdoJFrErh5U7s99nyVRimOEtaMJgytIVeRavRg13TREMxLl
zxAEcF3tZ6pPolAAoLRstm/V7OBlgnjH0Mti0bxkCsX6FwB4Ctnht3uAKnJyZdEO91jzk1N1YOx3
x+J56hVE6oYroQOfNW+EASPY56ExOOOrkygoh7nYpwxwKDTQtxpLTsUOCIAIqhFY7jbCPfiZG++L
unjwTLhBMVxZS7ypVErBJGTS8aAK0IXn5lHthdj8Lf4aZy5H+fX0UFN11UThDQ0rLVZ0SmDay4Lu
LazX8NG5TM9TinwVGfvY8cNJpWkLCmGGvDCB5369qDFafY4qQtqMyb/rK+Uscjaa2JoVemagazGp
vTr32wqJt6qQuOulgXvNlJuqoa4g26zvH3cDWxqdSWZOQmlQuADwzochE70F/YCL7Ps4mn/7Fene
2ze+MLfve85KAATWihpxTaS/zhOmXEIugOZ5ZQa4ZTXUEnPp/UXSXKJOJLmNb39W9ua24VW6Abua
0iSe1R0jFFpNRoqZlKWRs2FA5cgJo2uYeVlsYyUppHWzsFHVjTwVPsVwgY0YVbPDWQLAIrDmAgVC
sUs8dbzZUTDmseDtAlKsIQpEJNBWgzchnrhH8tOUlMFyv5oM69O/LWLfZ44nlqhFeKUF2Rwe2D4P
5b/zv+HIRjgm8LVfTCSS9njCULn/d7zx4vBnDIKVDwV3zj2KmOZ8DaUTzeu3Y0vq6RYyOXO+wmva
+WppZN1xqSNPCrc/tS7xty0gA0uMKvreEqmDAnaqI7lvp8yqKXZVRyYgvSCme51oUI92RPZY4Osl
smafFxVsIUoUfHmGUuiGSFFSf+VELf8YDMPsCUe3QjRNA1H30nJSEUTu3QaNI85d+j1wrHSQ3Tm+
gLsSGDHw+YKAnlFPzik/mgjs49R58PZYFlg6Hw1C1x8jCfDK/fmqrACVe4KoANKvLULxwfinZi6j
a/P1NetWGUbrxaZN/nAZ3gucuL22pPj6Vdeg5XS+ulA6U7xhZ05rCck+gPj0bXgbRhGF67eJuudI
NvuNwevsHXKSFpwfe/Ujd1cqPYbLfpvL2XnqoWR4rHbs9dynVsro85y7A/XeLr0FlVnCIo+4T+nx
H2+aqRKNPWvdQIGocA9Vni1JaJccRmSTl+RL1eQf8v04fYVtgfNc0+tmNXIgeiK4HFh6zaaOV9JD
Nd0jDOrMsk/3n23dl3vGlUlqT+BciRs0jsifejYGue9bI1dcM7GtcTXvse2S2NaaKWGTszOcNqQp
XVuKQTSrb7ulzmIkH7TjK2lyJuc8tM+du3cJzNvE72FhujLiLYc1ipfmwrK+BC78AJv9e56OLbQy
T6jMihpqx41RGV1/8INJEFyeJ4MJ5TuDfgZAly7xDRjrACjB6K31XZ+s8g2JiveIrrMuJOU5sBer
DazvhO4o1vCcwiy07Ad9Wojg3ijLBMYob8folsxRXX2mb9jUTcLG+GrUeGiwYN6/skBWJPIZj6CO
uQ9vYKp4PatTHKFu6rZPgVg9DCVEQMWk1+mVaYzky9TSY1hWiGc/WdsG+VBdrlghAX5wHi6FOwIR
1wxdLMQvRgT8/LYeb4PvUyqKxjpyTYEg8cDqdDwVv3O7zoKo2otlGBugqkHU2frsJBkEofQvyjHP
4fWpBVooNoLWRr80Z/2CVtiD83GJXGNgmqeeJn1aJgFdkRSY9wwe/sXFOsCXt/vOp7UELaZlaAk1
1ET7qyjWLPkDBBEsBxE+AzULwYFFpnQGDh6MjKQZctw2PIZlupmGiQPFy8Dtgu6tzKbD0LZHRO5O
LewkDVt81LcF+XGAlQdUlKoikINnL4oIpU7ZLvRfTs0Ly134tatBe5IOLlQEsWhO2+LWDSYp1ZUt
CnJ26llNY6m1YhVD9h0hkIf6URa7hNmsVfaXmqI42inVP74wTCliUppeAwOseIQuCdN69snBDkTr
vM6GHZOelnob35kEMdR5s2HhKIenHjXwQcW4734HOaFg8udPJqUdDaoSJ/rFrH7bUokk8HSXkb80
itIkRotjH8tKa+fCXRtU/JU/6l7ULxoObOFdB2CSWXbKAPFSoH+ertWZyktuDc61zNag0kY+kb5u
umGXXFmbMr/QdftEMarKAbY/QOZ0+MX3FFwTjnM5OX613mFCobW0uBHEZLLrh/0FsTEKDa3o4D5r
v1WGWJFlo0Q0XNGzY9xsfVfOCbM+n+BVNQez36eOlmxhunRHSESXQwmLy8tkSB0AHd8XXsSoRFV+
Zx9CpxHDFdNZ3ylWbXrVDNpTSxRVMgWJsLqzU8WcbXayGTq6OOmV7hmv/iJ/LBFYDxSaGcXxje5O
ojkjb1RCPDP8UHzK0MYEjV150k6E3cQL3G3EN2HqzF2aOsIwxj9T1HROHhFRrexK5e4YgpMPPfIv
/cixS0uF9OkekQWOXoxmbycLu3GZRzPWvD7TNtPjtxt0aAI9Hn9vcN7qpW7Uk7vUvdoFxZ0zjjLn
nlitJEveZgNznWd6J6snamM3P5LLXM3SVrrjzxNK9gLJj8K3kbDM8hdHOsmmIeHdg7A8AXaQBWQ3
pM6Iix2rzyFDKEfxKab6ZmOcXVciHXfjnPJsUSrjmS+eElChFDmLyv6Tjfqc9xVq1Ck+ZzEonenc
LzY/1FtoS1H37ALjKqBdNMidPSt//Vibj3kzGbXUncvBHDkT3h/9NlHcgjMk8qU9nl8TyhryGavv
ZXH4APm5NXj8E4Rp9JKK8EMtNfogUzthvRbn5o6fWek5iH8zIMJ0JOB+wuU2+BEJgnHaes3VZ/YV
HuZka4juyWE1jc+uF7QAW8EEmoxuBzKpoeXjFb/9lSpry2K3l2CRpiyQ5reT4yZ7SsxZyMYv1vM3
Yn+tS6N4qp1yNgQsXpPTUXahQN/0ZXrwFXz/9P93zetR1vtIBHvQfsCbNP8xzBNuxnBRcz+qL/xI
QzbJ1prZZNiLEq7ZjRCg0SFFGmViGNqW32vq2sNnyEy23Ygz7ZWb3/tUutIYl5LqgLOzSKPvJSw3
X8JBwpmnX/BXozXy/h4bwY+UdtPqNDAKIV8aD61s9VFX0TJBzXcxg+NPQBZSPhvTw7O+Vp3Rrw0L
VkvJYcF0+V6RxfYXMhNcxFq8yefWpWDOe1f6Eu1xeKhdtF9LcQ4zJJnFzdpWmh1pK34dhezR0EaT
sqrHl6JVlSg2FPdeQP4XA082tPulo3kyuWxY/R2P3JAVf26gVHocppD2ulWWdhktcOWMqM8pBfVy
OIPNRzumEIhbj7DOu6sSzWyPMLW1RK9BS1zFGoG72TYvx2RUVF1nMTIu7jD5vYWtN+Sg+Ir2nJDa
Nm71yfRiz6YPZ7eNwUidaTYj76SXC/cBbpTiNSTHQcnxtHij5eaUqYTGJd4vVyd5hSxsDdlKo/OX
uk2KSrT579Gyx3snyRwTtOG4r04UonPNhokwnS0eazI145WIJPlDIST3iuMcj18S1GsKeD6DBE+Z
cCZytkemS+uEpZZCQ28TsFs1jrC3VJzR8yjF6YrmY5WXzwWxcvW+uSB5d/QhR+qRFC/5vjNUW28P
Rxe8whfeOTA7EI4Gk38snAxgODnjacg0ZdwRVJztZSZLGq04g2o6fzK8twUj/YyDmavQyBwq2MkP
JGvZGHR9T9LMYqB+CJifxFUsIFNnCDGQamka+FVe1RDjOtr3O9KcyQ70g5omstWf5oPoSsR1McR4
jzHmxeemDLTl6kiKnSFUuYbZST03McWcndMtmqyDTDF0nExxwxHI1XyZdkYYS/h35Jjo7ceOH5cM
WYUhrIBiZA4LQG1tlUS4sHDh4HjJ/53wJI984C+faviD4R6s36/IHcS5KCBsDDH22++3JCLrbszN
GtPfMjavLe/h5BKYaXP4GcxJ3TjXF1xNkNAFaaxAPmPusQuD1d8A9n7DD2nQJ2YGqnUMcDwDl70f
NLFuPYKa7k9IbyNn1Ut5QC/Or50L24T/sPMy7OGwe1ZPP/cbxo1z2SFuVOYpRb8c+L+MJOGkGshZ
79/s+14NNo7Xi7pps5Z7xmksILEkw58pApTZ7qnl3hsBf30ijtxt+MMczOjXGsf2UsvpZGvSQ1zb
oYMkiSai7ehsHMTsGZPg0UJnS1/B3Xu8WZ8ekkE5tIoOtS1QQaggmqVCcbnmdbS18lS7b1buHes/
Mun97S2T9zpAMIXamBpMvdTxTB3DotYvslIKgHlvCNqz9nWW7qKt0u9FbwqpY9dRs8GjPPmGgiiN
GLi0HY/ZhG++tViHR2uDRDrkCuRy0ViJjrYw0Fs38O8bVgE5O3CkSxiFya137XX1GAL04SqIeVBk
l2ZGc+NMcDsv3NeVihjx18Te5skcXiFtNsYc/Zi618FEdjmc7OnwjyvdG+ET+l2oCg664xfd18we
fagwvf68DqKTQLoLd4lgF3ehHc3z7CUoT0lpYxi5QZEseEagueH8k6rBT6dEzmYomVkAKSefzVc0
fuhefNvv/bAY3zKiWY4cWVYR6FULjtRmMQ6ZydR8lVeAfTJ2+RIxfgZVqGB9ju+/SS6ajzXgzjvq
z7LKdxuyEQDDD4wnw9M50l9YZ9B48hZOxfqJ9/x2g831kvNKeefFTBL9pTauyb/YXfn4r7qe+dv2
1uJAo1+RZB62zSBlXhxgCwIr1vTozmPaDdFec6RJjhQCaXlBdy8hq3So+D5AMwi1cJanpz+DTlyR
OeMlmn1aslxG0e50YDIjzKjdbbwhjOk0YIz9wjC62oJRNy+tZjEhUpAT6mUx1jthKYok4FNgMRGd
s1dONQVb0j4uNfTitNTLXv6c65pXo2tMtYnF8A6+OMY7zMIyvR+JAfDFi8C5PSXkkRRXGRyg9o/d
58ps2/Z6SBKyiXzuWaMA/1tWf4O8wAN763lunGuhJrwGNfZCS27y6v9uXhhQuOJG3babc6TsmJSp
a4s4jjOSisfVqzbCsMS+HhA43eeGZlVktT9CGy9ej44TUpi2+u2PTMtXT5DU46XS8cb8vYZS2T8s
mwn/tEX0zdk5YjvJC4wRNl2mmaE0bldbpxLzBL0oTP/EssIQJeHu47JlJKX9TLD5KXWkyZmFch2F
IVyYMVVn7iizlATTHnw0ragXi+nqlwyqgWJ5ecZ/2X7Igr58J5pLShtwHwfjX4auQvB6HxefCvOU
9tKN3M7o/7zq0YKkmROVO5kFMLEyzKHRGjZ9IIELnv/gQ9snXsfJiQX3BEUIdg2etPU6uPlmSIba
68AkMa2SOTKlGJl9PAr83seLY3oOCiL5t1DEmV4hsPX6aVpsGWUNIGxRBKy+E6gKg0f/5r0K7hb1
fARZpoG2LdbTAfJIvYr4UbnyCvvRBSaXNSxfb1+2F2HwwFGApyTX72+hpuwHW60MVLwoTwia6j85
9QaF/jz/hNA4Lq8O6P+C2YdKBchrzFvrU7Y4kL8wkPBZcB/hOf0wTgbrUTk1o5FuIBF19lZztutN
2XfRLBYz5qG7BJYPH5Tp8ARnzeZYzmo0nNAXzjEUfw+8sxYAIBQmTEvKPhFAq9ld4vGGO02BjRru
mBsqZmEZtTNJwUxA19xUC+6eT5m0MF8h6r5s2LrsqCDjxJ+iD8uXcBccZ0Whgmpmxx1I6J18fUIS
iMVnU8pf5VbBMMXZY/39vfLLhJGMiMGFdEliaL4mPijRun9Dg/+OMdAsWuNOmzIWNtZw9MrQfFhT
ECc1xxYGmlFyTVBe0xG2SQ2NlN0vyk91OttNdiZpUF+L+Rh3BrAN729yqD7Q9XDTGqOIFUZGetHE
EPHH+ElzSuvb30sPJDLHKKZrKktPIvY+80dpVh9GuwLQzBUZC+f0jdxin0Yv9812OuG+GxU/yt7F
+dVkuhDhlK6cPyHngB3/crGMtVWrdGP8y8yQ32PMccVNpkp2e9g4SRJhd+3QTOAkJHSjDUN09MfH
JHhlljuE4pBSyZmc5DsaX5rvY4O1zbdkBRg0Zyjj1+MdiKftT9plssK3dbxtO8bVNJt277Sc2j1E
0ecT/yvSF5/58oFELGRXQksu3a2wL/hBvUe/4vZQ57e6+rCt2XzbB1opVtbe7WtmgZwFHT7YeBxG
cfPP4FmvL4HsFo3HOPfWqVQD/tYJy9IqULYF13QBzNOdEkPwd0oqxfXp6N5JPI3sHjf/TBsUoo+S
Yz9SyrQRv4wwqieqQmLzJ1oU4HCClBIMio/vDb6tfjydgC242t5OQVOYR/o+5DM5OH56sT5aLynT
zOoDsJ8dwA5ixTjM1k+44/0HLOw+vn6+MoSAZTApzBrhRxK/eawLcXuiS9JRRAERzITxMlNEV4HN
EAiKHET1q3L7b/vEFNxl5UxiQcBI/6IxJeC4z5EjmjdHKIhu7ekHp7Eh7cYJU8TuPulMYdDeV58R
E2K6+I+6Hvg5M2N9oUPzSfbQMMiMjVPPDUjCtz9HTMDz50eFoNoGAL80gMXp1DjnsDsjWnLW5W/P
BUMWqML5ft/J5pKIJX1RHfWInj7hjzP6FcGS60tXWrwnR4VuH6JRy6/PzSPaGeGG3OeDQc5TowOc
GAnIVqLL9rVudFYlPU1CdYSU8mzmmrVDCRbR1+saculGsVE+qkvp9Zwj1vrDNZiOgLdTmQyFZZbE
smlxPcGSC3HvkllOud1esEvFyQ5RiQZfqfBCtt8l3ea4Ka5T5eCarUx2GPNM838g8KXe81cJWg+a
J/cYh9FSVwGm5BPOvI8XxCg0JZb/WyJVmknkDO+OX4L3qIkKUpvAsgDCImYy1vebhlshOr5PhbXY
eBfH6VdObJG8O1SMq8SMoq9A7VUb/oJsh4medI30XRoQcFl7VDs7GT/RnhmCzEjbb6pWSXIRUYiR
rdg8Qi8RYCZa7hrGpnG7f6fd2jjNhI6eRCM3QF50M3FTgJvsNcSDOp62venOujvR7NPeaKqZicL+
xEjBGX1jBblDa1shJT5eJPEAzMZ0HQ3ecSuWAwLwvMz+xEVEjlPaGKCQtBK1mtviRvO6Wp8sQk9p
oi2alMaYSRlpui9x+Ehf8FFh6lIru8GkXX2WrMRRPDBv2Z8FK/i5jIujmhAcvtomzMXqJVNLhMHV
2KLqrxO78UOUrKTJ+MeqyWwO4iz/MSj8N37Kd14fLTF3oQA0CpTekk5FuZfJ98iAC+UFz4WRIUP6
08U1h9wNPP77eJv6MZonZzk6frpGheamH5fZYuw4y4vXyDmOqSIcHaRrjQg5+olxk/GH/QYNohXv
0WgIIai4olj96m/+XrRi3EM//RqC/BqbhCBJOwBehgf05k1GocxZUC0AfltM0wT0Un5Q5Yc6zKJd
/X5qsRf2vJ7gxRM4S7/i4eG0+1LkAFwRF7a45QISvf3sRaQ1Gekxb4j5rF+O5t5KdrEDz8RB7tGL
6mLM45cq1L/NfAwYPZiPi6zCk6gCOA2lWCwsWC3r5Ql95hT22KfNKDo4ZTJET5YTS0S02z64GzAv
yWL59AmGq18I9CFo+WFO6D18YWrqqNohI3JH/mP5PkT3lRHHW+ni8DcW5RKyE/wM1j1CPVZngUmh
bTRpMB4Is+173o8qFVUOVi2K8gxhXnpgJ7VONKfrVR1LTbflQYLvgJ43XQRGECawlB8IRE4rv0nI
EtNpVnL2emsVWELkY2LVlyoBXniBZiMMmVbGSTJsUOhMOdzNIH3vS9nMluGaeOh8pDqlH28SJl1r
bx3JqaRf6mJ6o+HHANZ2uKimzI+IlB+dEWOIXA/PmQC1lteZrBMCLr9DBWGfmB+k3OaQ5rA86xwn
SDAtV653c00IzXBT3clgJA9qO99VQMTBQd29ZxD5xD5xicsVEb/asdf4gWhULGM3r4GR9ZB4cvye
4Eh57LEqikHeVCio/9jufkIpGiTvapa4AvnfRl7LWgA68sLErolXEK5vXaEY2hUiAqb2o1euEWtB
OerPqdrUhxFA/ef2T8N3saVEFwIzt7wpl+N+gjrNjuYF+TNCKTLMTmaafaCxqz3NwRqUHlSL3igr
QkR4O8Krxk+lWa2fGTOxyDZ20oE3YamvGb+9Ii8cnNtXZE9dDbbdjwhip5q9I8blpUoPs9ntAzoS
+AQOWt/1NtXj18kIOI9WKBof8jI5vnufvAgoMVafSCG78NhR459QP+0Wv6Yy9YdN150DsGc7C8gV
ZF0joh52iYN/3TnKJj4MtoMJrM4IiJ+WfCZpeXXDNolD0Fe+JNZpzh9tWq7hwxwpYwYCPYbj0S+8
qRD/zuhWhlO/WKSnOTsRpK45Gpj3mfAOoL2TEvqfLeNyYkWB3wgkxloX0g1EIDrc3xAUovcuxgRl
Ce6+3FNkxZC40OTNgdTtY3jiwfA85Cm0OiOba9R59im/U0er8zbQlux3exw3umaEfOQLWxd/L+YA
X1YvIuSmToftJQU0/2qZzFH1apK/1ct8+O7d57AkaOz2pta9L/1bsURxZ//JUtECVimHSoki7hRU
EPFd8Dsq+1xFFcFNFbRkCV7/hfx7na4kwebEnVIpYpTMdEBdaomBsC4oIuhcKIXv/YqI/0pkianQ
lX7gp/8pEnPAvDJaw1V7CCCOvvHMryFUjK5rAqqTGFhixg/kRnXTa33SGhyYKaezDWe9rDL3DBDU
E3zhLqt56s9nu8U1687KbxqtisjR1tEMCRLAr/SLSnB8N9PV0TbnTm3v3UxI3EZNoOqzYZ+HuHGC
MXY4lYZzEeGnfRzlDzZyTLF/FgGBUxpUTW/tS/gQIqqms29FtR8y/bXBkIrdniAM6D80cyNzAng1
wLT/HMPd8Ni6fIw5UgpIcqzNVdfMoImIdg8ajf7Bc9ra55pKqsIrR6Nt1sRfPfVuA5aazA3Zms3r
b5t6yPXTrSX/dM6mVQqTllpuTxQcravxHYurbyl5joub3qPULBCJVqF0CfFkEt8LoMh9htSjF5iQ
IGvD4Ti5w485IXgTTpg655+nGk4rnsa16F7ewaQAmQ3ssch/Wt3JsYHcnCVkkxnqJt0Kz24oIune
R6F0fB6DC773fLoQzCfYnmxKlh8+IXFLZsMLxFOhNyWeVwupeEFVM9o9fRKJq5cGaQPId6zntPFN
CuUD1hH2QZsx1L81DeS4iYVBI4AHyKxkKIzzmGrMQMHgf9ihXQSKnv51lkWe4GvtRed2lIgAnTBh
l5wyxO3UiBgpufaNLiKsKOltLaiPREWnZrDKA+0r2BCQ9MbkKiU4gArXFisFECY/QCqiFayXsNJ6
v/YcC0ZpVHz8ZprJVPOHRQb2UIWdXtrUqF2Zbr9/Np2fwsJWUhGss39VO5Wq7lRa3uYWWe+WvE8I
FoeXmz125bRv3GgsNQZqt29v/mHUubyq+wMzrmlYV5QJJk9rXL66qhDFB61yRRg542nsXILS8rdc
AOosWa9ThnZykJ+s6v3WzEcf+6dKWeYVPM24rviREXPJ//hv41H3VKPyn/to51nO466Qh41t9n9i
GKt1W5cnL8I58kwfFF8GGTs2xZi2652cUQDPWzpVwyJCcrQ8KuKo32ZeOZ2sgNi9u4nXoS72kJFl
f++Ik+5q9HA9EMM4iYVDow5tXLZeoGKyCzx+GyhnGWyywigEKIy8u7o3oGOmZ2+fKoHzOnTAJ4y7
BLFbfxrh7LeSTQjVShZClubKFvYK3w3id2Emgob2SEL5G4vWRhyOTHWThTnZV8TS8EL6CXDqw4Pq
7W27aLRS4KNvUTJk8W/2WQfRadcG3XIbTQltkxtYsKYAQWqHCeBsTEPThpavtjdI1vJS2J3klI/A
nCm6WuY+NrHjoLEUn+v5eFhruZzQ3LPTyNHbuiKJeTFEK+cPL/Sgt+gVnyaRHwlT2zf6EBUDYhUa
sBjXwcwpJLMvFt1OvsxWDAmNCPsHU94QlRKMRhmXNiXtS5KSYjvNq52LFPvXQ4OSV/wIwoCS8n2z
Ss0zpu1QUoLKxCuZJiip5N0kEWU+wQ6AXHvoeKj5nligI8+XWF4M2swDSvdhyAmlD1WsPP4bCuba
lmQFQ8dIdQEBXHnckijcX2SdDNsf2pjEdQ5DYGuJ5skSjKBndJUhUH+N1PGm6c7Oc1Te5k6PYizY
YNMLPTbOc8dxci1KA07uYVsfugGe/Cmb9SHH9b8HMKa+Jy7GIqQAhVth2TjwqqIYynDyMhargcek
SjhsmpaVMRFNN8t2p9cMSN+GRVt/dcVG4WFwdnPSrrnPwN/68rJ3xt3RHd8gNzqd6jHa0hbFpwDc
ShYXdNCwgWx2Y7PzSkWuAvUsfCfrHljgOhdSUh8ssLpOFTYPaRgRP4cmEbl6KOHERuPybbk+TPjh
4m4rsBelLgMUlA4AZvQe3TnhU2oh1PZ5WGuuK9F9wgdM0p+pa9ZCTcvge7w4aASEq0c87y24zFxH
lb9krlATfxDYQQu1CyjQSAlj3eCMiFhKo9Ty9uXZGVP+unViYklzwmvzNxIY9zn4kBKIe74IxX3W
xPU0YLCOlrXhOHWIw9WrWopmHnFCGmphZ+2lIz/CDMGNZtxU1sJ/TQcwweOWsiOWuEW5G8ZMh1WE
Dxk0MrxKCcDMnZBCGtdkWMS03e5LTBAHM5IbIpf36mJYUtQeXucXHZJklgehhCmXj2iNK+miG8CJ
4Q4B1P219bUfxASiPuYaR6vLozXv5MSrLwdF8LCaAF7x3UbhXehECovYF3Yi7UE+j+RPcmyNZ8pe
zXQUAiYIqF8S6T0guD0u1E5HrqiMhn9qBW1dflWAzhZrJFRYkTdeTrp4xLJ69rZ/k50QmfkBYHQw
2Q1Hz8bADuyAKrfqcHRvSEDcKEEPaWkaG63VgZ8FHKXPaeFTrVJJqIXt7fX0QV1Gqrn/Ep4bnUT9
x3XgLTTS/6kpxN620JnqlghxrTZmNA9qwF+1yMe7cyc9Q7xwkhDdlmUPiXxJInfqTDLyqMKKzCG+
+KkJ+GITBrQCB9MKQPahSI3DUUYsW5fn9T7qQHiMROF9YJ/8FYUFeCD2oMqhEP6mvOTrSwn7hH4L
x7iECdwSC2MeSpaZZ369bmwm9RYit1mNTCZSUFocitjRLfQRqAvwCAGb9ZBENbnLXt/+yd1wfxy9
qZfqP8FLlswZ+85GgBVkTiuXB8nabet7lUOOGi/IUW/nCbudXHD+KZtM1ssGTcr2cqWVwf+On9zb
pJyYYoZZ1UeJsUk7Gjb12HZfCqI/7y4+BkvHGQhzKWARG3GRj9z6rR9CWwa//SR4rAkAKFRgbazu
mxccc2It3JB4PMixv0IgzDic6p2aUOiOJ0t8jB07kBXKnGJ+7VG+MAOahhXn5zQrXRboWr+Asdkp
UPcCYuM0cDsHtjAz7YbrQLF1iIuLtpuBaUKooyEfQAEYd5Qh4XUd36FoEju8cyAYGTIeUcmjjGkK
V35XoH1rsNpDQzgbM4yELrTvdE7HS9K++M/YMjdzonCAvW86+YGJ3Z2CgAf/5mcI5QQMC2kqQpEd
xreTpOSNSoZtxLIniUMrhFE7RZjqivFjzIB9CxrwK7g3RFBUlyjB75LkOZEwXe0R1nSVco6CzHk/
76NOZZvF4VzU8kWkdF9YGHNaIdfBoTuSM96UyYRxkasEodg8WkjyYR2ja4ufWE3rHynnnLb3iTNz
eO9fSxhBj6A/mVkfT1AgAUhaeqwHR2CAaN+con0OR9kUGYIygD2OQ7w5bEloG/zOoClPvv63nt2J
oyjEZTwdk6/f4qHhDUsIS9hZxnJKjljypvx/6e8JXXq6RegOV3d3ydD+wjiviyFb+PrU4R29BaLD
OtBDZf+wUR6SNZS2R0mAt+2Z1HpAwWDNm1chmEGXsZcI7oIIYtmLFRefWdu144bm6sJ2R5gns/++
s4en97e8HaKguQTtCqb3f1B+tAbZpYX2mxtEnDh5M57N8R6VHtXdPfgVSDCXdubqN/tq3UdUF014
zZPVznOU6pGPO1+chly3N084od+fzsrS6tYZLPJI/L8BWe/UKbbxjM5MAyloKFk/SPpe4nsI3Kca
lCb2CwPViAwQGq6p9K+L1g3wnwfutfq7r/rQX+UclNMNLoJxHiahxOW1uFv0a/FPdbULGmpE9fII
rZS5FkLQNaD9yDbptlFxb/4whxvV0X513sEGclNXYDBBteSflu3tqcqEZs+yihCW6a7rRYos9iYD
a1+TgCGDupfU3Ib7FGd0S6/eZCftsC9kCuX9VL9PnDEizA5XD6gwXmjIRcdxF6qLvQMrgC/yk2MX
uv5+ji34vDdzWLLf7jsqJGunpMu01jLi71q+93LP9NDNFDm38hmKJtoYXL7MnZUhwRK4Xv5lPj5F
K7SBn6X1AoFetrwbr0N61rRUlHYm/9EyRkLczraArN1HSiJ/ZrjqA73LFEKN9ODzip+XaTDNNScN
NuXN7uQsj4UZhxqXbuxxqjm5wjFot3jl+kIeDZTiOe8ybM39EgUW0P768pocfSks1NSkYN0Wit3c
KuGdZuzXOTw9jC7KdWO1M0BbkZtwqbqv2I4Jvbqk1lA4wxt+PCEmVJtv2STxg02bMf9oQ2G/dm0V
Tv2xmSK1vKxFZy38Cn5CKW0faIzy6mgM6ImvuCKGWyd7rcjK/2vTeAwn4twxJZEIq+KgAl+MZKdg
+b3Ma2nkZSU/dHyVIyEajLDjpFTHX4eb/Ff/9DhJPb1gpT99USW4pJGgXkchf4rCrCIJjGcZ98NH
o7U/EtVttwfNiAleHU7g03KlHcOvLlQj/eO7C81wE3PXW5+iskYqyIJE6Jc8CXv8ItjQo5oRN2HP
T5UctgqP6bO5p6+O4DZfbO88U9UDUNHzrTjWoeHKlXF6utH+YazuVP0/DEnKdURNXNrYSZJAqJNy
UDD7ld1aKMSGAR691gbE82Bxe3XA4qta1vrzVqc3nviSjZLJu6O6sxmJF77jqzjf8BPDvVDPfmV7
3fXSrNfKoY7vUe8Xz1ngfaWKF3pB6zyGOlVz3FiywvZzUC5RUdWGAThlrbkhHc9caR+pG1Yt9dED
ejjwSFHmcRKVYslJSuzLv8KCU6FQ7jURPGfCdMTmrEZFYgfAd0H70EDlmsLpUAQqhBKCrHIuJTbA
a9B1kq0xsKFXPptijji7iEuhWdCE7ToTi03KQKSq60JQBH/hCWthOz/Al6826Kww29lig8QMxgQO
Vt5x1lT1FpCRNQKuWB4i4h8KFts4gS+EAk6xWVd1uHZOKeGP/i1wmRI6Dq8ARj+q8iMRB1USQfc3
PZu9MQ69AdaNGLzvOol7UwFhgvEVPGqx8WudY0+Yr+DHE553+Nq/PwMqd2EA2VGQ8Hyucq9Abwcd
Jk38FtYXuz7cu/cMuiu8i2K4gTTjCBe0w2Yk7BPKZDGcviPIEF94frYiFPHWUtBLUU7Fv3bC/wqr
eMZQVjivCQlfE8VSsu8nRLVszCSKvlyt1H8G0F3ueS02Sw3crtzNO+OLvpTcG990KxLOsJyBl9Qo
Q4KYGas32X26sukksLFQsqmBGFYr3qdLV6e4SLsZB68zTQvi+9YJtmS0WlSgEFlSNGaqehIrPtU+
GGbaOLNsh9aW7KTLSxOlpPeeWudFEy4oRytq5UOBAKuKLMTZ75wkCQIA4o9J6ibmE07SILVjjKCg
lL926i8Wjtmz8R9BIQQkB0Brp3O1MzCp0bRPNd+ItoAlXbpEuBHdm7TyKKDidOofRBYCj/TgXfif
wPXtDyfmLAcUkRmGBmlGaS5eXezU9MbbaSBM8xnADH2ILTHUPZgLfVac2E5l+obGOhVaJHvrMMvS
ah4JG2ZGzDyAO3Qe+Xpa+lpTf9dqvVa4Hbk1UxJ1AjXOoFDvwLGzipmWLjF/awVReo4Ko33VxdyQ
C89DqsHJTAcpGa11hEmN76oomUcg2eRF6OUNnVE6UhPg5HadRCwxcrHGvoejTtp4snsME5rKDjhf
0w3LsJPxx3/T/Y1BU9E6Atb95Ajbj4MbBVTKfFjQhzFrrbGWE+mfUKr7H3XnpDMoTMuERX39ZkdL
yI16tHCwzjNZQvbjvHMuv9JBd4zvZ8ifILyJUwZNUxARY0elj+kopLaSIwLfb7eg74c1O+RG+z91
xxhLmDDPdtBbJ6qVivuDO1ZbCa97qK1oWuisMp05qBwT43hOg35czERiznx83NLJipGsvr1jSt45
cyH0/3udeWcKZerkkhk+5zrPXLaL8Apg+DIXcv21usBUk0KVzGRJm33iLxrIhWtZpM9jxi9RcSYj
U6cuHE5camNzDEaQnlbd8OCyhjpCj9+QIwP3/mqisSMPp7Q0MPAqdRCvb3kZFpB6ikdBUCzv5OEl
MegzCkuZAfto7YrMjeJ9U5q24Al0uM1TMkH7v6k1Ndb1SOgSLRX1wbqW1o9y2/EKikW7AdmP3o/K
phq2ibD7gkixDCa1q9OAeEN2lObXLCbSvHyP1PkHCVW+vVNOtuTCIshmkecU2NBASugeLeMHxw/s
eQFYsFUpUrcpBysS6x7zXDEStazZYlb7Q5uVcXcfGp0+8eGukJX8hNKYkT8gMnr79dnMeqVF1Zcp
2Zp8qEzP7Ap+f3qEXBXTCW8xNjaa6hCP9cRTGsXK53HsW9OATN0HtCtP8PraSTdJd/EnN6uvM23X
sHXufM36Xy1OIPABSwKEebbOvYjlCarK9q4u5WrIRpMqSK8YENJGMpkIyXbGWWi16deQArRnrLms
6OnCac74ARbgarfSU6EXwNgQXqCNSNK4xEBmDMM2R0J0aLzQWgQZ+fM54BboW0OplJ98pxd9rqRY
f8qI69jzuDSM5+NJzy2uYfNrRp39mmCVFNESkuFx6nCsuXjd8o096KF9xA5/4W1lrZjK7puDo/yn
bzNj3jn3Q86vMdQCqSofzCiZ6fJN59dKnmfTePVXa80+ihCQP4mgcFXLGGuE7bQ3El9eFmmyBL9c
1FZjff3xrUbT/UIxFcMg9c2CojM0+02Dpb8X14KniV+Y59LYsvAcIQ5+G8FghBfeqYPMpo7xif+h
TsCJJpTFv63/oKK7ldRMpH/zkYQBcObVM2vfVuIf8HWM0WfMCLD9iy08TpB6m5pJul983VGsQ2o+
O4c8Dn2FRYwBdggF4ZDpFFoMRhBELwIrqikXO5+xyDArEaFriUJYmpYX1KAYyWaNbfRI2n5FzP4G
MgM1dbcOI26i9rAngI3UZB4+4nlp6WQG+g2xrp6SnkrhZpNJbYlJ8G3nU2POR7umHTT+9fyac6+E
9DUd+u/ZiWWfe3h2RfO/ujhq0WWpy8fGvAURQ4JVlw8rG1YBVajd1BjC0GqbUQ41QZz1DOZAKnOr
MXg5LvcGESIUzsYPjH/lEzMKTy4AwVN0WM/Fl08wvzTKz1OjGPTYjs14Zvq86a/qbI8zjKKhiV1Z
69fORCB5wiCzILtlnk74j6Nn6jifm8jdp0AChDvZ2Mtmy9/IQ7006/gRnEASHlts5GpGrBzchcom
kN6axJoO9+tSHAlD8jOCGZzRpkzaKZvqEA9jA/L4uZeOwUJsw4p5WyU/wRDY+uN67hjqL69fOdQY
deZ3IntPU1Pjv043JM28d38F0Cw+c1+Vqi/6Ox2IRu8T4oM/9NydVik9s9YmpjAalK4xkch6thTJ
bseH0HNz1UUujgMzEognoT/AnWaVXK1CUF0eHn+jwZNNv2V2dpMUQ5PI1S/4utSpRx59y4db2JKH
klBd/5W1u3CV0uqsevZaiulGBlme1f2LaF6aBzlc91lgQmRTagqS+0xwtBcklBcYG+0/SH/2OVyR
hUV4eE9OfIAAHMisePhCKSpmfRhFGm/csC2SpTZ3SOtAHUHgQeyAqiqS0rD9jKEpMN6GGd1P+BGc
LfS2ueCLoiy9vWg6dLZy80P4kUk+C70kH/+/UEgHFeQ3m4k+GFIfBYxz620FdYBuxQD0pkiAtDUZ
lM5K4QHlqjAe5OYqjZ33TUnYAnp470YoFDUsWztq7BCvrQ5DWxedBK0cdlMl2sLbK7WLxUheFRBD
m2BiH6gHVMcoJuDISihiV8sm/2SkoAp7dbxJ4BNH1FMauo01IHEg5szyqYmJF0bP+MsayZPTbkCX
m/bSv16O9Wrud97MQzemhwD/p72aA5suA4ulwUJQ1n5tHxFp0lCF7xiMtmXt3sMiDh56L0hOx9Cn
3nasFCuOuE02PxhN2HzV/V86TKh4Q/5cQb3mhBlRn9joSh12JWRYoZYUBElC1CMlmWL+ot2nZxJG
lEBg086aLW78AOx1ikSTAsdTCbznMBXW54ICLlrKOm3ANyMcff40TfEvt4T7GyxcVBqJJvwAVhRi
SeUl5VkJro0niFPMkuwIrDt7szpcpbCuDNQsdQfyelH8wq277KMZXrBWcYFRSlyVoEb8a/1SGQqN
tWBIqz+EKmkYgvYJlYcd7kR7ylQh+084oJG4LN5yO6vI6b0s2r0nPZA2+RlpT0QcJoCyDFKHKPwo
5i93yg+FdcsMMs/RQJRdGzi+PexVpXGftEf/QGqCwOYsOKMykyNRphYGM3VnMq7+qKiMm7LjHWdf
wKnpBhTaR1Irfh+BVoFz6tyWCZ1WfHuhjxuoUgFtT+V98xa7Tooj60+uPKxrYPUOhZQlJut5HJBl
j1/AWfZW6csZrmyMtsaUwA4mFmn0KHSefEvZv61OjRrUxSttwR0yJEVEnVRSPa39PVti+70KULks
a4jBcyi1zwHlCnJ9M1jBY2SLZ5HEmfqzTM2v+SfAamWXd4KQpmEB9CSor5NtssZReVHGjwcTxkqm
wDZgrgxkdThhkCh84bnb+duG3lLkUvsheHWuN9PsegcW62lNTIGrekrkwIQ4wS0cgpQ0+S/oQC6P
avxYM4fRq38nZ4vC6E83JZa37VmUmcHHk4Rg1mxjCKWNReN0bTAFQ0jDj766BJNgMTaRPckwnexA
viB0ED4qEYStNODeg0FROsRYmln9RUvHwhJ2gylVVoL1JIoKAfUP64XMJ10euDoBezo7nT1fHw39
uhpQKMaP1o6w+jO1GRMYYfzsqIoOuGw0xgPPp2+MGq+Gr8sHcv3oHNHAVSNlwt1fU3UvktsVJ0ib
1f0lv/K2DDIdmOM4rHOOY6kAWBrV0HCQ7sKlauLB+jPvAT6HuxNYzHm3tCVLZ8rn8tWuiY2weLVM
ng1vKn7jcokVAO3r+arPc0YuyG9cMLp00nFQy+BID58hmY25H+q8T1kppwKGo5q3XHZuGMSEQMWj
Z9dHyzMqpWy5i4qCjOLDnhtUoQlRRZmmOq9Jdd2Una6TKI25cjsn5gVu++lDkZSjThhPs0SAu4u3
8JXdcgSmh2Mov5NUw9fN8RxjgENWVW7CVJEz10R98ttSBIAc7uj80pHO12SSDzesRieThK5Dxoi8
gjroF78Nh5PfsfkigidV72s0z8ixdBv2OKb2e5RY/6Ocfpi13y1dfJHG+v/JOdciyNAHvCD15j58
f19AIspmAvVIbA9M10bHkAbQPX2USMHdYRtu0zs+8gjVdB34dx9bq2UMatFGsZ1VV3ztk0ViAiz0
26SewxKF6YnEZA91nNge2iEhOWYVANDxyd0Cb6C6acVpmoDO0m+59qBNCCUmvTdKojSYaH6ga6Tt
K1fI5NYYcFg8yEtxiDPlMDoODHPLgIjbyxZeP1zl+cQWLrqwQ6r3uxcnpN+wfHFYZ8ffCE/igL/r
wmd6Wp++VvKlBpGYIiN+3veUKHSMWcRS5Yf4HjH7931sDyejC6SgEjEkJI3bKQavwJIzKw6YbQ0n
rS+p9YGUBpdZo7/5x7jB55Xa0Wmuj2pmk/uk6OyAlDY//Cr869dFLdLySMH/IihLgigOwU5IosuC
vVvZ8h2Z0FFVDsYvpOEe8RqdSh7l7HjvIzb/lIKw7JGuHgYi1J1VXOmUYHcd7UTgxO6vyDVNgqwA
IgDaDIo9hJDtGh+vGYBWQ+4MG87oL0zRhPo+0D+wm6Y9y5F+XKwBBvOdFdRQFn6rf9hKxMPEqBpt
+AKjuvWVeP0ccrN1SW8uZqzcCmTqxk9RjBRmK4NzkGFHrjscS9XbK+jHdc5CjkWGaWHZFuYbvHxO
VxbRUMzdyH0VYfxvNWiDx8iaGW0WjU7c3oBxriaE4TyXt5k+RvGsaXP7D3AvnfUffq152EVgggCh
xbv9QUntgG4ywaXDVMWdSG5KYhAQhao+ObwIN2Od5zlc+PgFpYxtMaETdM4ikawvX/jDTLgURfs8
qtbg9AIYOnY49p8lIZlXjFOoHqgwyaY0rl++gAyWLId8wimzyWtXAJ4ev1WU2rtVTymvToSriAUy
LXoh4VxKP/4qi0MSyAFqVzXps70qatluaNk0sQ7dbLTSbThJ9j6aiy/h4zlt9/2kpf5CKuwLfpOI
LYO+hil4Se5c6U7axX4rLQdvbi871S7oKfBkgQW7rMn2q66FymYyjnNe/AwoSTwTOUBLtT/rXN+4
goJYv+mX5j3q+m9f8jIGgYBMizUyUYepHrMNnMskWChthCcyW6Msg7dpgLgBFzBBjvyEeo4KDAFj
b8BYUI5+L3PkMugmQNYNMsXo+Y3oetHbwKUuKVMdqYcuuLs0TM5ebjMa221lwiOomNYuq+l3PcjE
y2Nkrq7D+afpfOiv9scpQ6HAOGhLGGLs14c6OSarRi4FEYzizheNxYs1ODzswT2hTOILnbrQYcjp
PZrOA244PDoGyV/91cvL8RtqevdwMBfQz4G9PzBWLtK589GKo5rvKThMfT7olHm0MjdV3ID94Go2
JueSGzfntf2QWK8TQTSdNN6ThS9E59L4QcsR7jkI/NYRuGbD06dco/6to6jOhVADbZ1sj5T/LKGC
nUvctWpNrRm2tVgm2199rksSx+JY4yKlwzEfcmXzDF1dTB302xx5nWWZ87pJejDufFxd7opBR9Fj
XxVyEARhskYeh2Kxg7tRBvs64OUxXvXFRNm7GQWc/ZAqGKeTIZdOG6+SHLvvTx+CZa8337LN+RtV
wvxIJ45bheXoUl+2VaWFCd4C7PVnGMZYF0nvEglGlNOzW9J2lYXobri54FyiCvcYWG7zFNX+aHeY
yowoCO5/SAEm9cmoJI6NvLN1DlTtuPEYwPf7dlm03P68pidZt7FsyxBtG7aZQE//0Bz531AJdR3D
YqpYIWiHI8PLE21QMcbHmCVAqmV9oLFDPOrGAXn6ehUCJxbUAkwf8JTuPis7Ia6RBofANwXpiABP
DEUapdya1lay5HKx1QBjWrMPf60uanLCW9BW42P/udgHFMGKNk5CTdPKxVwH6D0OSNg0oYr9xslY
D9zTca6piazseBcZcce9eM68DsExMKeMQEsb2FGtopzGSwDF4y/b6cQCw1Hz/SrXu3R3V7LSNryt
oqarOeHkjxMvK6UsVBBEtV7k3Yw5aSYl4dfX8yrOLzkjF3CD2U38vJBiDrTgah6nrnY4cZcVzxqg
pVNvpyc/NyFyTt+/z6JY7LM3g1x7Tk6GLxoPsyZtEEbSnw0pYAjWw+ofjzrsZPHLM1rA8bDL43AD
Bizug8C98Ne+K5+nCVTwJ5YAJ/WAoJw36CGH0EOYF7BkXuVtyITO+RaWIApc+UxcXDOtjeG4BnP2
qW2RL3zBKTVtIWQBOqV5t+cThQYw4FLJcuvTUZG2/H/9a1ZLZaTDTqyDRiPBmp3x9pVjFLiFcGom
IMU45lAGdtOsCmunDivK+RyYXsfcifVHPOq+Ff2MH4QcF6uFhxz1Umaq9qiqiLfFIlDcMNNRxsmp
LRo4gJTufT4QqpsmWxpBG8zMoAQSGnQpUSkWVlxElxHr5t2CZkqEdbPbwPjTXkzS/yWE5vRPZnt0
PWyIZnRV/hPaUMYcIixNGvpdzlpdxhpN8h7/ufc8bDw05w8lN42wPSEN4/7tDEvNgxukDJL5W0cl
VUlEa1VotN58MGed5N3rbaYcSVGc5FdIjPoyMyMyzn562chWxyXZBwrM/Gj71zFSm2k5vW61R+nh
M1YssGRusudZO4/ELD1xRnU2oTrZbtJCu/xMq83RJCS8M4qlPblL3vctWRsXtH0O9vD0mk/+kF7j
dJ/CmzLaMe5QZHrIMHZZxpRHJnw78CdLDfhbKydTG/hB3zqII9c/3Bo730hMOIs9IWwwHP2YTFto
RcfhBgVR4qwsUq97ixPAhElBTZ/VGqON98BtZdHf9h8hilwPuMx+dI2HDFe7i8Alkit4RIep/6Sf
Y56ULJwDgdbf1sRpotC1YQh7ylvTqh69/kUwTHgpOgJiQ1/KCRzaQFqauWLbPeNUdGRkBNvQCXFr
SBM7AnBlle9P1x/0bCC3Y0EKGvyYcLfx/+gsQWAs4kY0W9O+k3faGOZVm1Y2Cxv5MpQHoK0ZZDRk
VkBuIxzn5QPXpRdJnOag1o2cIeO7j6CqzK9BzI8n4EEyxwB6PNc0aAVDYMa9igzBdLf3RVRO2GI/
LF51IdYYrm7JdDykz6Ndl2mBK+ggn15MIXIbwP0CU7acJzUW+DzRBrMubSwsH9+BR5yhk3/zyBxF
tFf61Gl5GrDEaw53YW52M50B+3dD/X6XA5OOcxZJ2bCfWZ47C/jo+FTTONbD/8+OR/k0KJaae3zP
BuL2N+ljX5A9X6M8YPyfBOvxcDcLPyiITYdudbCMi8XgBFChMDFWzhiDnzLKx45QfwLQjykgrps9
Mpl4hovgZWXkliLLdT0kg85V3btgXPEsBiEcBWG8YIU8vLh6DCFiJI4pTFU5XcquWNQcLSOG6KFR
6on0FuM2cxjZQ9Qt6XqU0QhEs23dozuNzngNPvc7hT8IHjSoy8RbUedi3ArD6xGZI5fUHoVWjG+N
R2HjEwXoZYjcRk4eshNWisGMuVM5b++iCDPpvolkRNFMj7qqRqEEpGPvs1cpoEkyJBR6EgoIvfId
DJrNLPquzP6gMdyjwiWf2z/o/GgwZCYk9of0LMMIMEXTwjHsKYIIJD3wGWyFTLWVcTlLFM1l0HQa
/MY5hCFoS9e4gdjyBFfompyZULnuIphW/JsV8hzygcVked6WTH32BXWARQmYrFc4ZT5+JnIg7mkN
OvsoxcKF21S5OAqeCdrLbUkuXv1OeVnjyt9P0gz6o8QplZPoIxs+QoK1roRElyGiwbRyMb0/MGXC
WB1+yTPJ2JY9jS05unp9x9gvgSbKEI+rjm5VI+6+8EOD1FI4QfwP87UZprdTzMYn/bsoCPksIfMD
KxBhDvxsVkl+AaiLIbgTyugIL4d22YxC5uR/v0To6lDHXU5qgHSruNFdjDtgO2ddyIkIiJtbZvpi
vBH9PQNpTeVoI4zwMBTEpm93GXuS1g+U15+AP2dY6uiqsGXPXP5D+Wnv5LE5if4cYc1iBYs2Xe5t
+2HZGBu60uS5/ODE6Me8HvYoK3WH7laSk5ns7XfAUQN+MerMmfUXPPceIoc1PvP4/EzMvRbeW3ZK
rf7O/ZladVcRKJG/yjnCQ5IAhsWbZLq2GtE9kAe84E7jT4y9Jl/BswKq7I47veOoff+KQXEBGW/b
uEYWT8Xw0tVfUBwjqmZsHcHow2etlDfj5+geYXbLSBm9RN4xlVP8ByFfzhExJF3QcnY9jMt3aqcB
4H132U2bVnaESh8rj4WtNVIVDMknVaZdg8Xa5U742wEZfBcdxIkIlu/rBei+v3D/AGowMmxeWD1k
jVADeAWOvK8AJW77kwWC8Hquna4aD9XnNoYpdE+F2gMYCceUSISooAP1UY9CaKMSvCwmpFgy/7sE
X4o2ar4rFutGJXePHlYTUJbI0LStMolh0uHBeoYdHzrKTWxOeS+55r2oVAGqhcKi4XuG+cJSUd44
2/KujYNWLdkge8OECE48rtfcDSFhGZOdmiZMpCZOfkueqhqNOG2pwB1SWLZ6DYuL1/dHDcJ42bne
ZjxFliA0UfINNtlnWPSuLywtKM3H6g/TVH2VC+JcIC5TEkEkWz+arGdDq5q4mrEJfyrd+wWwb7U3
h9MgahMrnnb+VHoTKDM3i/cNUqBf9IZTBZ3wHqfxabecEsyXxHBJZJFPq/RHb91UJUR8DkNF7FZo
25uulRh5xd4Dp9jq/CFF4fzG8ml95CXUqPoe1ymj5fVZ4IA6/4Jg9GZPaS8nlpn/1L4BoC05drc2
YmfrogHa1G2aNHsvXks3N7kciP8sUmoMCGpgxZpMO1wGCKuNSrfOjezMKZV+Pvgc1kx0j/IWeRoV
WuWmTum90HPWxxox68Hkaltm7XnFomNBGzCyekDIF827xweBBjF17SMs8JzciDX3nHfphjuW7StV
dRhpssMQFbL9mL+4Fa5Z8P1GO+7BoMnIqy7YrnfjeamXmho+oxiBqg3rz87RLq8qpeIqZklXtqxg
6pdTgL9YKtN4/HEU9l3acqiTGw7sj6EzjFrdLq9y1UbL4+yeunn+ccrh+V2gHgSPpGKzzv+xUcET
ls4Z1ahRN+OnP17+/SrUdnH2I+5oKIZiKWWvF0NDPmbIFVlzjR4CY2fXx4hPIA+G4sUuTWJ6CStW
xo5j7uC9EJQdS2I0bBIW0w4MS30VRvF8X4Uf0dchpBMGasnNK/nXFLWkOm2uw9nsKCh0M3wLxkEK
ewOU16Aq0xwJ0pGQfM3Iltm7KqqCUH903ZF5SML3Vk6uWk+X89q5U6ZqOgIyuvQu4jGIk/D8HQH0
ZN4FCnwbmY1vvStv4ygIxXnnGRoG8OGv2o0NuCVkSeBV5754A3R+3Qimi4QsgyHCSkHMCPojXCQg
p2pqqqOnkfXOss5Ov91skRBXuzyiX3Il/9HWKFP+B6l4k6V3JWwhTiocUt+3aWUE/2TvXno2+r7k
sVRlv6b/x0buRkwTC5NKnCwSTYFyEfnjlYQyJUCriWAc7gRS82YQyWMHdSeHuK8+sC0aZWi1oGw9
QoYFhX5IaktkgqtPoDg/mfT3MN/gAjRqu72yzc49n5poNA9w1o9AsoS+nqCEXDx29c18r3IvUOCd
rw2+FxwhWLGo8fAf3XAE3YYWI6g4/9AvApe7aWZH0KjXzyf9LtLxf5RNMSCtTCv7Wms3DN4GsOlj
LAsaKdkGKtPOEnu1T5guLiYE+iNd47PJSrJ8DiSmF2AvLQZzZLtQEGB0cjse3I34vMvrDjQyXij8
D4lPJPcSJkhQQZaFXgv7KKp6IjEMsEY7bbE24bETNgKpaKOI2R+QCALL6QuwfCiGNw2boKi8NeAH
r8EZoVH4K6V/2NNxX9I2YSK71W7eT5QgjVLgSSKkE/eA2EW0eJjiP+AgvegUTwxzKW2+1uqIOem3
o7XB6sG8pGfN+i1i5DuNFsng5qAwzFtQtGTDAiuLWmWfMHg8kbj3oyDJcUar6go+jODAY/ZnsM2p
g06Mp+aKhl43H+69JUx1zoQ+JaSaTMMWxivPAmFlAWx3oA4y+TKPv8fbded+oRAwVXB3/RBV5CiV
YoJ5FlWnDETudA3Mshs5ceLHXeNGbhteZS74+vuqwm4+LtONoW3zxuzadyCMtAKqiJ9Cd9oEz6LZ
00DMVZk0Y1W1oH/Ioj+Jv7di98blmVbZkfj8Zccf6c6rDDJe9jyB6O3EJFJ3KjDEKQWzf4pRK9m+
9JBkqP9+YKJuNkShQZZPVVngp2tqXj6EQroffZFbdTxMv49vmT4wJd76QSyt6VFDqvZIButlfDyx
9z4WFrLwEG1m5WxJ9WKwM+NmiTmwb8PWNlD01m8ZFCeI2YCEGTUwnhn/b5CkuYpqYvGvwT+VGeeP
MBWnU7R+t8vJP70fJv14/dU/+DH3BGsr4MoqNGkjmwUceSqpu2Zzrq+6YHN7hNYKpHAPI6t4b5Er
d7liLSYmK9JnIAuhtf/CJmpLk/r5nfK+SE0I0gzCQQpKVyXxT+NLBsdg1Ui8jzigLKZ10giDOsZw
Akpq3hTGL0fI9yqOQpIWFKfH4zJ9rkDvRgXABmV7yciIvjwAejzPAiOH/jS5t6uWoDJhR5p2hOPd
KxZyUQs4uxNQRRSEcrPOqG6oK4yu9EDiUjfczoZt+Rvy8GBWayEbeUlzz54WvB7sTXxFxM7nxSZE
VEqLgqfsRon+l+LgYUYJ9FkX8P9kuVUettGlpgv29oSWtUBDczjAB198xQVYj/i3vjOuVgKVaFrs
8qE/zoMyznhd9qw/HESshMpb5fi+M/UF2fZ7yZNxomWU4/U91+8peCq33XLKdy3qQMc3UyqaXRe3
s1qNjnovT5nKC22d/Sx3/oQkg9ZtnGbA3gDNKXFshgBRQD1gDFK9GkdUMXwHwaMv+Jo1xlCtZ4Qc
fOV+PbFZE0mp25AgPY+67mk0NG3eIrH8XgJakqNWqXAA+GVgOKRh21hjiGGi7D7s7A7NQmIy4oHn
pI4NcxNpcbrxBUeLcW3WiqFK/RG5aSIOPcRkbJvr2uWKaw2AOXStLemvGcZlV1BsDIWUG1Ii+mZs
InlT0d0BRyFUmhEzTxxZul5Xq4wy93aPn7fNdPr60/CnOPtCvNCjh+fMs83iMxmImr03G9/EykTT
dV7vEXmBRrvRYHj8wfj9zUxHcWmjnS9yXUpGit6tmRQIz6g//drCjTlnFaDH/sBNS4dDT3N1Upyf
Y8vu9fVByA1b3rhWe7buJqs68sEPA+rPIwFhfQ8P1lg+sE/TRboTOi97AdfSqqspDEjf1v/vTgYf
nLa1pEmGISeyhEmCT0ZrXpsyp3ENxF6X8HtU8l/SBtwOHWyDA7WjRKT3Hitgvi3qZZAMArPwEXoX
WDAGj2WAcIKyu4V7nxGU2qpvWesdt41dQ+Y1j76r70bi2mLjQPN+jEC1hWmuXQL7ZURZXdOSAm6M
zEdlGeav7ly+ksp1K0+Uh2OznC+Ri+BteQfWkysR13ozSrP5NGeHGyNEiZ+oxunGUGd4Vn4+8KhI
NNwk6YQTaDr10686LttZRuGIbEXT2NaG1FL4jvndYcDzRS9u0yu5vxTCmjXTz6Wzb7gzdXaDpaS6
PpxAnon9NVsxP1PWSJEdYlBPQQYVhS5pV94UrRBFdJFtAR20radrhCzxHAIYUBY0yVDlvjDQTQWS
AlC6Gr0bgyWcJCJ5+15FpypNL5T7jI7c4Hwe9Yt8dc44q6/ngVgoZhvJ6O9XIqWGlrSn5TMj4CgL
dGQXQV2n1HlT18jTKSQkgjmfoC2tRIKo9oqHtiHvCIHrrLdrwSJ+ZPLzKWQHoZnVLNcn3QC17+cv
4f3U5j8Ayf4jO3BMdd+mDBuJV2nWV0cd4/YsHyQFn2KKoRGxKtJZXNQy5Ki9/okGYwJb+xy28I6b
fV97AD01Oa3JTIO42YdgNcBS95myJm6uIHr+WCSssDc1zuNz5cyzGZ4m8UoZrD2bHmuB7/so6aYE
c/pSMAgw89zGcRV+s0bgRj8865YW6IAoagNo00BG+wXgiOG0iYw5nRCwJSinAhvFp0AGAYSdSibT
8jlM+TxlX182Fv8ly3Sz4mZ7sFAkFsddoNESwIbNC8ysLSQWcGv8AQVLZ4d5HjcG56uP0V3xD+xp
7wMVJv6n8EKIAul8ubMx1p5BLQzR0q2F90Y2yjeQQXWqVtRU7PPdEtck5U48lSPXuk/xdgfnleGy
kUbOe2wIJP01J46mmuq3sUyElVgL042JuRVxBBv4dtE7N98JyzdkZfzQciRv/Yv9MC0mKyYDpHat
hHSt0TEjsVGkJRgBDHK7PPjR90A5+VcdMNBFpu1G8Kgp/SVIfW5mcpZEziExN7vYmribXxrbd1Ml
8L++JjVh8n2MnVpzk3j5/Gf3Q3YL0z0u80p17xxW4wyL9pHSw6L0oeqG02k8RWqSp9g0jhHPamgk
GR+CxK6p51BStBbbMtPEPWA/pVVI3gZdCAA7aTx8PX7sLUoabT9QOo70CUWGdKJPdJWB6xP4LYNL
pN7c1OvjcaqvJGlOeGBudYz6HMQDxt8h1TK1NLhunBAGsO3w4g5PWb81UgRFoWnx6vFXT7fKNyLK
cdiM9bm71B9QiS9VMOB5z+fkduBoYflTE08S8mwDLZqeEfahu/2umFOEeAh+zQ4jufkYMkv1Wx56
hNvuDASA2zotyf4Hsh7AJjgEfMKFKEm7yGTJJT5ZX4i9zLaZtCFkCA/rtMxt/eKRrbpCFb3r+zbo
CC64X6adCFLFf8A4Jcm8NEDr0a1BjNyq2189pZyElMPDi/l/W97jrMza/EWXDtotkwzloNwfEv+6
gL6LuF4CWVD+6zy5oKgK6vbf/DowR0jhkY6/ANUEXjbmS9aiaIhsjw0b0SueyoxqI7rQg2OwHB5R
auQvIo3fkOY1Z2X04+reaHd6o+i2XxFNOOIgWYBbge1tN30B26G1vvYQk+LPB9nT6J62ZN3aYwID
dWR7iwJb2i8Ljh8quvHDeOeUGeY6wP8B6JXE7RP9BiX3X9ZQabwqJF/ak6n6Un9H/pj9c92GTmAT
vsOrFw+FfwvTZ61Ekl2RVu6d2T1VMFydlJ3PhC9mAiqmVsHse4wgouNLdJtc3lrpP97KXAgkRNVG
7gD+u6JK/OASln1C1NJAcmOhwSM3/XRc+8lYnZQlgv5g0hDOIsLTclWOuCgXHYHpPYGzrEKh0XwC
C+UTaFQB5RcBR5q3BQ8Db4joZX/j689n2HaP8GNxqSaGiVjzKcZi2NxO6eTXRnCxip2k3rmu6w1i
RQSU+1DA/3Rkca4LVmm6U4gzoEuPgaSlj16dlgkjq15nKn5JufiJH0XLBkxqCAeNPBaeuB6CmiB6
oBGmV+TLoJ8+zpQcI6mg5y1lxoA/Dh6D67UAF9dn3uTJhUSdQZ6bhAkRrgt+9+nrZb/xL1BLPdzu
nIUiIipKILN09yjY8BWTdmg5vYfcgjBjB/Y2z4Ab58ZX/2Vcf2I9xarVgT0QYicwTMmTihiirtlB
jy80S4ORT1857qTYwa70UtqHyQ7LkbY9zZC5IM45HbCLKFNytLf6MoyvE1Y7fJAtFAE8iA+GUOhv
2hPz9X/aOHjOPGGq80D0S55F/8WerrILW5jur7djINXSd2anQGHajwefHcCHfIGiBNDDShSHadoj
VG3vvdIH7YLIypi8AUkzH1zjyIbUBLDFlVaWeq1kLDq1825hGomc09orJo4raN9QrcKEcTK7mXvV
cMSU3xfOt6+UZKZdxOCUB/ct0u6uZdIVRSAXds7+jzvtwADfyo2JpbcyyHZsVk7ce68rR/G6jXBU
+ZdzkB7Vm+qrhlQWUlUIBoX0uWvKEj2a0NUbg7MGGLu3o7EwVWDjzUPupYMVBoNdoqj/QcZmOSkl
jwBeLfaPJq1doBuyocVDlKOJZn5Oy7MSujfDEJv1gCmOheCU3Jmgq4cXl9ScFNcMWfcKYRiUBrjd
OAQBFMX6uYuiFd0GHzTKP8uXJMklVJlUL6q+Ei+JYUUvxFsrYU6qxAJkPyH8HVvBSGZ9ciDwo6eB
DmDaGmsO+0H1RDaJ6uWI5f1xNHU+LntkyNTqum+De2+L20OkinqfgT2H8m4eyxGY43mgY59l67My
mnPsrSF6Yf8yqZPO+8f7vwhmCeq62SA9BefCiF7Rg4LgAiqj2gFaKqHUYlNIWhaYmu4jw3pECZUl
rJpo773nmgiy1NGYlFIrZoyURq/gkK62qvNScuerPXmjtHUWUG9iT+4PbLVUpKkT7kb2WfeANvjT
qY/73SGFQvVlor2c4qyXb8cUUx63SvZn54GLOHZ9YBnltA4cg1Zm/EqRzcXSE95vejIu6gXkYFFG
bE5e6MFCPTiwNmbfglipZEBCde/Yh2xwp9NChG40P534h3PyCdh/biV7ZCbVer39/T58nZU3ZCkd
/PxLG64WOyAHO+5eWgtWEvOuMzX9qHUhlgtypq/28wrF63wxh17K354YdVCUWOI3APESsSVcdES1
lXI8350+XitPqyoCLzVkMewflnGgIq6MsbnqhySwME0xVHJqT53DeWyv3OWn6jfQBCPPTLYiUjF8
dHkfBJ5LtThvkY8Nu5+mDC3rseQ5j8x4ynyO9dHUw+2NDuG9MGVYUuyMH2uBdOOnvOaD66Rh3SAn
P4dkepFvFmkp7SNcn9KvKXES1hnqTUJAVvj6Z8Cg1NMO3Jx+PF+KMA0WGuv7sCYeVfziwgBKTQhP
eLshT1zc6G1T8tkbcP1JoMMBdNYLIrcUYuCKfdzBSUWxoGhoW7T1BassVwJRdKAgVKxau1bIMu6V
l+FXTjaTB46a1V/L9lSCZ9ksY5FNgMuwuV8Ag2wQRDs4vRIP2HQ2Wp6OwobGtfO5Y3LIWgO1AxuR
ToA9yFBRZJ6z3bk/fQRoqvKNGWiShB7DetG/Yciuvh9UmLPMiW/fTSMasRFj0XdNTXIvBLa0RDib
y8q8xlaQ5meyPRzn34yN1/8Vahn8nEZP/mbxekIP5G3993mX7rrB80QvvJ2L7KWMOI+ikzAnlGJS
5iO1cfkTPsIyKGakEV0VcmI+ApCHAdoBk9XhvYTRpdq1BBgO5B4XKjDok6DJwElT1YU+VOXjzq6b
AuFl79yxEjQx6Rr/hfcx8poRpLkw0U/fEOJ7OkC8v+86jvVnDXXtIH6GrFeeU1x8vTpqgtjtb10I
zxbEhmADkEPb6LDzmMcVGgfijrC6m1o6ZsK4R0lK7pzTlZYULiMp8rU5/pNL/bSQ9ITheVNrOD7P
bslFf1j/PCRYVDJDGf/MOghV9FA+4oKKOPjFofynh08XdZEwRYKsM1+SCQk1HXGORlr+KxwtvDX5
DKac6/pOnv6EHg8WtemQf/B2iF+0R338h2EIN/HId+FVxASPFB9rJLgzM0G7KgoXUgBuf8hv+VD/
8BsLlDWFeFtX2bM4TWqxR7QQxknOpQ3lzqG5/GMwAZ0zCBW0mGl9LDq6jfpG/ip+YP9yi2RQxrDK
1OIAKDPAT9DZCj8ctwhUFInv1JgeivuptLQeVKaNqQFc8wvnZ0Pv9KLsiKyCxEXkDjs4Vkm+WKK1
rq3qtWqN2tiY07lrT5mSFat4+kiVlza8HjwejjjX9cfobo86q/5wR29SBnVhMtUI/8ePLgfToS3B
GloKXRX0+tKCWrGlLmWP0YFVBy8NR63N5EHn5mW/yjNcJDSPY95gy6C5vwZ66IN+eHwiK8lHSGgJ
Kx8AnBTuReknjjiveJorPWBywjuZP3gogTiOrfi7eDc/aa9rEYuonQJlEPEmqnd3VahP1iTWSdlo
fD6brPgJ+42B3/w1ApZELUeG8g/xNdzd8euKxhRvPG74g5ewLekq1z3NtlcdGHIRPKjlBHEdMAjV
GWcOnACx+K39GqeqptDp2lx55/ysLXs6Dj9UhYkwIsZS84/70V/2TxshG6AccfUrCX0P3zCHMiYT
k60oGKYFi8COlB3su5nq8+Ieo9GE0gWej7lmx92bLJJlbHGiCNiaIoFBQ7kRktfFcLj0kJLpQMcC
dUcTmJ0/mpL3oLjvSB32a6y5X/5YVKTLoEdrVpPlYYnlrtnbigPLq8VGtA9FNzCDbExBjJuGNhe/
N2zI3zFdAOHpcJk/b0rX1djFkLX0Pp+d/Wqp+oz1UL30/m6/Ye8Cv+9tFIdc0K8lYcoNK4dD8jGV
uGPbjf0/cw29HsFBQB3ipw+tm9h6HmigceKJJus+Ny9tTXx9n/Lf9XBUvT77uH5NmZiGz4+3srmP
7rd2z8NfGVzMR3b303MBdGQxn5B1UusyvK4tM/rKxLAJYoNuxDNxiwVpUeBmHteCmgBE1u4nNvIY
uL2UKLsAY7S9zuChGIcYPhsgoqW97A+L4jm7Ql41SXEfc6bMjGLkZ8BvcdbndTbbfMc3v/YrZEzt
ne9mLvHrCDWxEKbdnWs2zBJoCYL4U74vB/gJXkOJ3RQIGMsjO5aeV7TF5LlXhHQnKY8LnQ3BKShh
z1BcLbInI/0i4252bS9BC9qzKq2/Tn5RUGpC1VxNqj+GAy3ztrP1hqz8n33IDw1Snq6iq62mgq9S
bBRVn5UYoDS8ipcO9hJHbv2JoSagMAKCLpKPmai2yE9GwiSyXyXqP/63snwvPHE+KobxBWrBGPB1
qla/NNzXa6vMGrv72mLYcJT8dyBct4oqzKFzN0eNfYlxjESnqmUmQQ1iu66HK6lvvm2GJMTTxDde
S+9UGc67Uhu3nJnk4gxapHY0bt64iyxWm+osUhQVdfSpGYmpb04g7bkweCKdwaz+CMf/DPm8HoNp
Izhba4RQycWQhkZbU3DPRFGSvpokp4PA4QZc0103CSSY4yYGEfRIiZ0seiqsSvwvvpwLvFyU9dX/
K+dLH8u7xSi/qlPkUYK4pTWvEP4R1RG/tnaGIujIUFlsCXPiEr7bQderEMuhBg9xJSuG9WB1Cnph
b4ihfyi0q9+cyWhECF6BbLO891BthNCB94tFDzVtcfW2WS2U8pFlGHQGOvjxhtRzgGrIHMa+61Oi
9rJugqEW2UL03jHFfNLvcS6bfg3FSjimCNZ+itY4T6LJHanhZDDstxElE8ivCOdIGVHKYLc3pk4Q
VpbsnfAc8xoxudQy/fBEizCZU0joYiNO/WamrttAPWnWMPT+GOFoNsd8MIgz2fVcUKBgY2Frf+RS
+YUrkYPbkkln3Vv97d+j7aK4wLAAr/vqD1VXmfloMIXt7P8r2JZBY3v5wc+kSLJ+ZndgTtSTD2i8
ztVSzu67tiLVZM+5L/ihr4RqFEcw1bpyzyXj4SuFykwmzZVkYrRRMJh2lBhvQfrRUgyI9KkgsIij
NAj32aqcUjsm1V77asq68EGw+PutHlGvRP4hCrHosGiYMNlDMiUTPhwUCiF8WfckFseb1RrHANE1
eUZnrDIj7K4+LTxH7NQZIaFaGOl/fSqRVvzXkFWsJd3yNXxVU2dyoUm/aI+5o5jLsml+fUiSRyeO
iUcvQS7UqEOL/XtTeQBLm4npxR5pMSK/p0TOLVsNnu19xKWrQj3ERk+xYLY8B3JpslpJ0JvdfonU
6J1yrfPlQScP00QIfSdwk2mNJ4AZ8EyR2osLf5QAzUQXUqBue7RygFPUvf0t/Bok1Qbp43E/+x0Z
mk1W3K0HzOIT85DVjh7gBrpApXgUkcnyYr0/8bYQTTbSNUDryQyq21QBHX/4E0eeQFXNIvPM4mIB
39p5qe1k6hEzUUlrdw1OqASBMBJgsBg8xzE75CRler39rgiM13kBfydmJgDGe65dOh3+fjEtwWwx
IyLDBDLefjOYTpCjw0T8ZSNHCAlc+eqQu3oVfTaA/OWcDypBHJr5ze/3r3g+byXpN4XfuP0cFgSm
RvlDEUf/TW5/j6Xbz9Wpi5fVTaP9VyI7DbI9+IfXVMr9O8fdyCyB4yvDWjgAlFThUKARITEKC0z2
MYVfLz0LLmhBYtMpgO98gkiG+qO9kv8Wl/0HEKnqEm9E/oyWDCq74o+axjqwVCdCrOKN2Cci8uc8
zjjulAiwcoaIcgeIT3+QKjs696eb6+Jof5eHPaEplGyhR4Wb5H7DVe6U4Mxnne4Ix/C5GnN2aZ2+
T30grXAbzKhp+QCQsRjf0qUwa6WrCbTMddsD7qIjM37nSioJF9T0H/iQ7I6vwu9Cqon201OvI+M5
nyCM2R4P/8oBPPr6te1M1xwIXOrFDTFBYtkIGIVwninP4vbigsSpOh6cJAnHCsl+HU3nkXZ4IKXe
ubzRxx57B4rhemqidkPAOFg7GQqIkUlg6FWx2sZuHBrFQZ7vGMibGQNd7D8au+D5trbzXQSL0v4D
WcDvpYZ+V78mELojX+k2nzsJHM0RaFMWF8oElzags3OPwBsKbue4Ks6KYG3BNe3N8Cw7Trz53Qmb
V845Z5fzYhlledmDQGiS10dAs0jI+zOkZjovzDQM/3Nj3fLzwD8uip4iZ0Y6ZT+ph9DOYFY/uSOo
TnWSb/rakciMZgcTPtb6uQq7DPL74rufzsVITmX/bKQF+nlmj/g9rqkcojT9cHVEjzohdSO/U8Yn
itY1wqH7iSH74LXByeH/s39CJM49mpPLsBAINCa9bypa+1Zx7fuLrIna59wN75okWurduxZeFqED
4klfcqLV6cON+VICXlxijXkazoXu8GfSQpmgHlc30bz8fPAdK/xfguYcmE1xNNCjm+MqtxYMI2ix
wbH6pyyJFCgY/ILITtqo0HPmVQSgGvA4GZjpJtyzZpeC2R9/SOcsEPoAJQUrHMoavbm2UV0uqnYV
7kmunlaXhwRfdroFrfmVVDcBNpzrRFVxnm1Zeb2hVDe980fTaJ6cG7NvJwPcm+fx6XpbKOzqYxVs
qvCiKTxfubLwsgf20Xr0TxFMy0cpSbzEAvQdWJxTD4ipwR6yDzN0IcutoxUYlsWZcT+LCpLNdnBR
dOlr42pvmQrM3x+wHTO/hjHfDkrgJTkUmSzra/mQLHke7hRmLbRtf5styD1dTN71eg7678AX7+SG
Lyy3+/h/9O8+hkhDkp/08eEmpq9GCH/HlJFbmbN2f3HdVhsWL3RRuh/GP+5zrQwA1qJMIuv26Ihc
C+a7mPcaIaQVmx+AeerDiEAXCWLGXbNh8Gt8o56phcgCdogRIb2sfq6lQyfk++naqLhOdIAR6h/t
9h+ejRIZvAC7JUFHYDZ9KuOL0vfWi3dxm1TVbuoPubWDOtQC4vLLvS4q/M4cFBCyEKTA+EqPdJ8R
O81OB/OUFInI/bP9CPfMwdNqxRFJ0lOGeEmypH/Q/SSfMDtqFSaPSJk43+EO73AYPVsb05+RynWF
Mmqe+aZdy6U7UsBrBBNd7l1G/SGjI08yYrsZ8av/kOceuTFobQvq8GE7bS9dzyHda5sUDN8h7OfR
bSbgqn5d6rdEK0TVQ0OhLBsv/Z/g/TaqSg39pIgNed0A5BFZliy433gr8CsxEQcsRYvChMZ7Yr3V
U3dYUxwdWew8xyuG7HNipaBTEYqTahYeuKTY7cyG1PLPTqIi49Il52bBwr1FnYYdqDKJS+mkUeOe
1CMNayxD3H0w0yYIuVJuSabaTJgeU/70Awodi8C1MTBPKI/zDse2vbLAHZ+sAtJ6x3JFbhlZapjK
TiwNcE5AOTULB55W1u/Ifj+QAXuUGUAmG5q8mw7ogRVmSjyRq31OriLsmLJTrey1+MHxnV+2Ge7y
qQ9mFF9KC9sdCegLjJsCCyR2FBtkoKlmZUeRIPxKjLnvA7NPxdtaVOdevvHIxWeWEl3uDqB0XIH4
cOkQ+Y3h2WgD4KarFMTpR8NGtfjEKFlFzPrJj8VFX89WdxGCyJmukv2gMqmxxces85E7+Nx9Cp0c
vqz6ACZTBYu38H7LbhEVje3j+q2jZ0DYdBe7sT9D+88uTQOewvPR+Zs4BmNUc3hXilT8NR7BsIhs
tMubB7HP91xwZT5cQmeIciSQ2n5ktL94gI+XTBEi/uFbFO4bU+xQo0GicQGfvzC3dHJazyBpedj2
zpL872D/S8HlBUuQoDPOiahJuAWTik9iIzIz1wirMKszi3/gi8clRpoGL/UdhmKLoGLs7woTT0fC
u1fdJEjkLgjJSTKacWPu2+EaVePysPUDqA+oT6cf8fsqJ8uzFjKsi3I4r6qmOCcjy09tngyDiKmd
VoNlYXZqjh5LvFs6GZD+BJHruVgnlsEhoE2OSLNsaaQ7OVdEFiFuw6eWJHbaW1bEjRJQaXgTehdf
CkXBm1/zp8FBrsvEY4iyMotGE4mzO0wUncsYrtVqU4JJdGXodENHWpT1cR5U/AMMI/y4ESXuVe+k
g02PPEsXtxpflNsN3fO/W6UrBW0VzmsNRWaUn7FVgvaGYx6G8AS+eA5rhXkKaAQy8xj/8yESg2Y8
lPxgmsJkXAYdfvphPlTxaLMC0rRwXerBGWJPcjjRFUp0TbYoMcYAnMa9uLmRlUC0IhGjXdCm6BAL
rU+VUwEvSIZFS9Y+yre+2KGC5XlgFSFDlqxjaavjcb5p/hTcn2WZvRLmpdzj+WnZlQS2nnwHCxNr
BYMT8Stta/YQ1hR3DtTlx/4KiKE2htq02U7sLp+GQ0MoyzfJiQ3aHI/ReLQiYsEvypyyHyrsOUno
Yz4kuXrCo6ZGWFbA1tHU9NqFgJ+EWe6PNUr8KSGGyrSK+GwTOEiFMxMRK75uJYqvNBraNEDu84C1
x3tcPv0Qzgfi9RtsPR7nX/JSZDyDBoRHl1AqJWRczBSWybclyTKsEYdo9aCeBBWc0UHVF2ED4Xrt
lHhL8nFJNWmASQTP55aDQj7aDdyntal/Ad0sYzGy/xtNzUIzKzURepRy8jhaLx4BocLjVMC4SqO+
IEfz96qBchNJzyRryVQKzgGrSpgSya5faVMF148IaBkOxpQ2OzxjdNST7lRi1AcBQ0PId4UdK+FZ
HCu6AaTiagKoZgBqrfJ3CMq/bnxqeeVKOOx94nOzJZf+ItEHexrIaZnSmLeHq482Pj2xt+H5Al6l
F7+0JAvtO0TmtjzKLpXpsL66oeyutqbvT5MaRtz+lqy3weeQ42avpUYdLbyJemrCV1XE085cPB7k
zKMYUXjzMolKpMMhTYqzizWSfym4u2bq6njDcGPM/gI4daFSJgP0M6mZdiwa5CmqCTjMf9MSzsOe
WFr5knx800exOgPOk5yy9ckcpcuo6u6jXY3vKXLJ5TVEkl3kou3ZobwYkgSWJRT5Lk0k7ty6ONe0
w8l0WT2ItZLXc0Ck2ImLu6amr4KVqcSBUbuBkkiuIG7khobuSc6+eosGns7WffQfP6tHcRRHT4Kj
uCNyCZPyMtOE0cpZom8w3WD1Ltktapj9QTzhsyUx1PLMZB12hZDqwzutrIPteyPMBclXF8wVIJz0
CmkjSmzSyJ7gVuX1SHdyVwgRInPtfZZr4S+wNqDHewiUy/1E/wkUqWpSuuJm4YVjdD3Hg/dqryLx
Jza1XYLZ/yVZr6e/sU7WUFMjJoTtZxocC+EYc6cWk+XvErfvJ+q9p0L7uMXf2d0ysA4xzBwst93j
GdskGMDMqnkwFTlIvzZu4fuV/N/RWSfQI1X1mWzJozh+qTmq1QvvyF9TwH8tR4ggEHczSiyTCA0p
iMi/izUTuPn5u07iSD0vdiCIJVBcGCRVXowX28+iEPWTmeUDuQ4K0LZn2wCQtv7vMYtx5+5vHBNl
60IdrSfr5LsHIX2sKVsva+s1kUCxzJlGNKnZV79X5FEaFfSa5biMjslzVPzkzajT+ij2WORzNS2d
dtMpVgjyLPYmP6kmaxfMl1bEBZ9dUe0/fe2q9OjkVYW02VKEZzqx57MX8mxQjEco2jx2nfF9Hd3A
b9ks+t8V8SC7I31ilaC8mUhz38fzNz11+iz0F0og4MPYxnRUUJc7cYczqzX9aCIabKSofn/0T9IQ
282pRCEltfVJR6eM+Qjrdx4G3EKQyDJGbqqvt4Lw5a7KcATS7bcW7PjkFCplz29iKkBy10QS1w4u
dkmOnIwfOjeKP+Op8jSnJI5h4GvPnM6hOGT94w11Kku1oxzL9kp7F+NSV1umuOi4kx6IvpjDRbOg
JfG5Jt2/IC1HhA3MECLsmUi2fJ0jsPkciBGCc6s1Jyb8Inn7dmCaIc+vWrF72UzBGWjcuMjDUjQ8
SVQTRQd6sdCxn6b9x4gOA5tmHZyXs5hbqhZUxwPgTaCgFsMlRRwcCvlw8tCaPxthfI3IC4kcPyAW
0UTa/QF9whKQWTtTHgXkNN1cismvg6O38O5JFS/chjHhwUeI/bP7OVJvt8dZy0XDe5V+CfYLMdd+
DxAa4Lrhg6F1nPo9TTcQkUp+u7xIaAMEvKw3RPwW5ghORaWmGbDTjPqZBG8YltvWkHZSWOFMnZLI
ddFgfqoiXXtEBVXzeVav2ebqCOebgnGasV5Jnn0aIh9lrjvm8g7awpFWcFmXCosyrMLYkbeeF90+
loWspsUqH1x7O6Sn5LEsWPtzoGh2Hg4TQNRR8osSR3arc4hWO60sv16t1O2xfU8HU5XuNNvNgDWX
o5nqJItSWNjivtn9s0/9zSi6j51JrnRgP/5ChksxSGpHdCnaqEHmac7J0OS/LuFVOeFFLpjqFVKC
auUVhx+vmR43kcGFi3MpyEkPg9Sl8c96fiARTxw7uTLg9mLzfbzhm2IOld5E9SE145pyx5O/bggH
OwLa9WXe8ZqELDwGX10/CM4d0XGJOzcErm5EItwXCPbRYLeE17yma/SHoXopARumRuumAWwOQprq
Pid2rNuRQKTZU51J6a7Y/jap4ipR/N754fVKGfx2z8Hev88os8OOhfWJcC/ffb2Qyt4rfQEs9RxO
5S2WsUMK6Bm2QrH8rPPmC84Jy6ExNBTaHAkNsrih8uneXynNqWtXXi6i2R2Rh/ULH9UasQmvRyg1
c9+AVQeTQD7NKq+zt0sF1l1ixS6gY+TEzdAZVK94TerPNWpV/iw6JmWZi58Q5WFotuqd/0KHrcOt
ZYNth/0rB5Rgwi/YZSS8L7+kXxTbyq8qmua9RfcwM439vRB8UXle2aJK0all/ccotQ92+ocxbCji
OcOoQdpfqufR/+PRfEoSaxFhhLVV60LDV/BCPd8RZfRdYXfukRob5EMtDmpolee8QLTchXsU0m1+
AyuVHeL6Gm/OF/BGYtgzPyFHrmuEiH4l/2jIOXqKRd+pRHDhSUytfjRsXVv0FKbBVohJo8qFyD0e
MJr12SrThpp8egy4iiwZB+yY5+r3yN/zGt6eN3pZBOGwHxEAzCI8IAKeSCejhtiRhsNp2xNQAhiI
hdmkOqN/U3XAWhyECHhgn8nNi0o8m7evtAoxaXJIlUltdkhz6Jec0zA3jSkgIaUKSm1PSIKKDtK4
G19gJHf8B7PZFlHQsBG8M8Tjc/N0tovUiTU3tus0c1jZcdh3GfDjZkAOP6wMswHqh1l2fyotjj2K
o8WFJ52xl7ZWK646hJS/iDHksSOY65T3AJfX8NvpRvEW+1E1fOB7L1zD6NB9rWZy3OJnz0tcNSlB
N3YgZwi/t5upgDNntcAsoVBx/qx0fqBeKXNDod+1KVQMc0AS/97L+b6f+gXCuqzOt1h/Qgc7SF+v
RG8TnxQW1qItGhzEDNBnbNwf3w9Lvfogomwz/2AT8BSZzBbJE/AW2dR/M9Tx2/A1yqM3Z/9nXxBA
fNnp8MjXKFMT60sOlghU9Dp91fCygrhDruoL/1Lv/rcUcyiWKuwZNFbvhoLO+sHc1MH6sJekdFUS
MCW7cNgFHp6+5xcqYrnzBL3zRWBh0fZ7grXKDaaC09eFsdBxHquhj8en+EJ1Dx6YFwLI+kG1+ify
6K30z+zf75ZAgSOGKq1t7N9u2PJS2WKzu7c4X2DECFNwgAP+8qRLJErls2C9rFELtcNK8m18S/Ej
U+B4bwhyZkEdx1z7wboQAMsiY5jZvcTyQ64XpBqAGkd3s8MtCNoTzahMRw4qYqDje1nBPDoszv/E
wUSTodpjcV0tlmDtDw69RG2wLY4SULBshBQgdXkJN5fIDI1Y39w2jmoZVHVBqMocay9HiY8sTfOq
4ktzQWawB14Ad8PF7huhtqpzwklD6ctgPKHusQfcGzbY1nRAZXh4UIh8zTWHM3dgRtzIcBM2UKwD
TJAwRrewunbcXScnTkwJdMER42E3JzdFLhgg8T8oXrKgKBVlopdQqSkkjiZIXxse0FNlhu3ZI59s
O1L9xeFv36rgRqn+7aBUwXQP7+TG8rzF4/wvgWx1/6Kw5PJLOFlmcoP5MPEw3PKZf+cDnTEVrz+P
qND3DcU6hTC6KocbIuHBUzftBYdEVdfDJaN1dd7vtJeJ3Od2ztbeH2xfBNc9U9J8sPQ7pMg7DWRo
Un0N/gk1NRlEluOv3wwSxiVr5xdsK5g0xUlUbxDxaIF73HvxYNkI/QdBSoKIOHc0ZihfHHNA7560
MUT95UlN5YA451OlUsYK7aRSkke3OqmEchuBv6ANPF68mTFE7BLi/7jDOyt5gQaW/q7dd8hvrLti
BwE8WB9YJGVjzXbcZxxtzha47FSuwwPR5k80oqOd60AEMm6oZ2/CLYwlIuvaP/8+fAVcA5OVrv50
zYXd0E6rvgM4Vi5iCEtptNdXP46FjsPlkilGf79Uk8e/mVTVK6WX+TkJlsh5lgm8pBhJMbYSSkvN
3B9cCL8RshtqCfHzDd2q7uoN9CbzoXAHBzCvG2g9JKuLyEZVpbfeLnVCv9P/o6uYd0UMngb0uJs8
rVkjP7wPW4OHJKROm3/N3NSsimaYsL8sB+gsSGIpnZ55Gbul15OQ2FkAUN3MO+4+td4stbirSvih
DEuLKn5zJvcHJwVgbx9lKXgsmbil9ubXng3DXfr/4ZjxUSDFwFgddkbt14ZHC+olrQuMXNihhbwU
fAopy8G9twZZ2Vg+hh7gUdel0eBXVRsdsqnI8LBnmMJdQb6O2Q0mlfG0xTiRHFFHYXvcwJibV+Zv
J6jFTXlYtQDiEo/yM1HEaEU9ZQ2nL431snnVrjBhbcBzc3Vk79CaOq/zT0ptWhyh/YGgkqV/hbH8
WAoyq2SGyjjvxKYCq2lKGMyLnXrrFnAtvaucZgBaVA0vbyMPtgrsiKAo9SKUgAs8QZV+PmHwI2cI
DGSiJTo9Q+ZBcdEfcldPDk+4B0O9RAPZW7ndItSCjzgrbvwqaZwaW640qb8jYC4gdo/qbiedkDm1
nB9x3VaHuhmiNGEWbABs1JYacLyygrdMDBSkGYt/sq1DHyQgwHAADzU1HpMazi3ImIJZodJYWqA6
4leQA8oASA721r6nk/c78M+S/gzLu8DF0eauxnJiWAWIlOd+KN4teeDl+5FVpsv5pTE6f+oWnsSE
gXD0++XZcYRQWvDoskWPLxp1wdemmjc50LOOktMml9WsQfggCgwoi1jX/jiZhaze0a3U3DiErL4v
94mE32FHexv2raF03S3eaGtPFB14dOaNnpKcWGQuRlqXnkvEwN3eJ139o42oY0gHAnVzmIcF1nBk
UXJ+AbLAZeJn3RBBuD0r9MZn5S9CEkc8R6BnaIMaNP4h+M246zzyKvmU1mY0BvVdBMcgwfeGMAl9
pzQ9h1P6AZVNPhm9/e+uWrRvEBOR1z0DaR+ySlwxuA3HWbtWKD/VMDkiCEf3MkYGcWnC2JuUMGnJ
U1yQX4+60AWAllMJyl6DU44XBooi3U8YYGs8i0xqhojet/8uWR17ostjT87mE3PPG6t17W8s/E70
FpSCmPLzYx2qy3p4DVdXRUogKSJSTDbcPQ8FzAsvxy+FKZsUp/yjFhv9zsGg3mpFM9bsEWCUlUV+
uZdihLuVl647KvUS2X2Q+kBcB/1mteKyqQCRCe3/psaVA+TejTvb4cbQfYNXDjpJEweuw1Uv+/Ez
Ox4Fbni6D1aCxFJqBJfdw6r79n4tJtknr6iTf/JDve2mry3UXTb6TX96r0ib2hfEEurlABM3i7Gv
Ntac18R0AveTZ31LfoPZtUCiah7fKDMyoe3HasnbQto3xX5TdbN+TvY+8X1ElGO3K2GKe/jxbZtP
R03NZOa25ys4jHWx/7trTAvwrzsCukvD5xIqkQwNVdAikvKhVX8tlyKzCXYdYIY1wB8xSd+3tloX
560SguD8CsyYnd+SnWGoTuw26bfHb6qt5akn79TIU0mYURgUcWj3/6jfb3bVlsMoWmlVEqQJ5FdD
4GcBeal7QQ0Ft0a7CB8pO1j6vlywuflJmWhpX5i9Zb85OQ3han79+sLmpu8DtOallBXz5OZzKSyZ
n/frdalsCytqAVPbQgL75iweLZgXDuhCj78J1oSxhOKGhRS9jTZ4tH+saOBEH5EIv/c494GXbbBe
6TslhPrfrSKcejX2fF6tNx2TOtIzxAsIesQtDhwCtad8j6EzxOwmkMdLRKjvUG/khMHN/7Di9efX
yaKpLP0e0iaGOeSlG+mp9bBpgBNLOadqrl27JE6ONLs0VQIEDycErrxOdeJ+FqhiXlSTOn5RSUJG
qJh2ZFJbJiWJtmr3c8C8B+PRUEiT71X0xHjSnnNx92RfRF/WJPBZqok7ZjDuIiWwIHSOuKgRxLOc
Pgfn6wk7oFckjh5ge22dmlONpX+yFA83APLjTocS90qUWHN+HpYIrQVdGQA88bUAsJhJXrWyuQ3/
Y3IVDdTD5tv/DYxbCSJgZAUiCKDiHVi5ejV47N3Qlhcvs5D6G8n/RctfAQ9+i95h5SKnuglySRD/
6Td2FNmlZXxkHNMKpAdXg6wYqunu3yiEVFNO8bNvMKbAtTZ3rc7jNxzhdq/6RKR+uTayjkibZOmk
4UX5ZfOGNP27MvPSbJRu0VdshWnMyKZom2zgxwz6glS4Hd3T+29T5lrX7OgvxoNNUvdXhzjbkvkD
OrEhExxLdlFlT56p1AfRW4U6RpJ5yJV8KGeqeMubx7wnX0rgjCA8UmCPo2Dj4rAvm/hOe6QxVlTB
LwulfgUv01x61DzWoxQ2bdDE/vcxSMOiGXjJBaqVsmuc9wTz1hNgsXswAjnVXI+X80ijVaud4yWM
WsXLJGKqCpZ3tPN1H+ACfBGF7gFf0Z4Z+mPHa5QFILQAmNhXPXMWfmvtrWuh4mQ70x4+KqbMNnUB
UziI1JxGVMcqwTH+/hwrm2Ggy+Q0uePqeLAeGgZkUEKinlwIYGtPGNRlvyEH+41VxQZf9tgc/Mgc
Eo+4xV59uDTX+/UzJW3hjB9Vh6josF/MT8Htsawml/p1NCFObZef+tj0sLSeDzYySHw8Ie4W9tmS
TFdIuqaQh56OqraMBpqz2SQkZuO3ylkBlzaC+vouPL8ncRpnDMSMbCSLAmsoA2AB1Z8thTRPdwXC
0HkSModQaW9cvS4ai7V3oMRoGQtfhM7r/VSyafiZgjNYUqX6+jz3SrJokJUlmWXQjGMsXSS8DO3j
ffHzuHV6Tpzr5xu+GH1vnJPVbTJ2TpNaMecMQ72KPzHR3EYn7IyNgW8TciEggFvFRx0gOPGjoler
vlx6Hp/dyUNhEVCvYYQiJ9OS+dz/kkB/v8YiMl38Zx6Yrbst/8AljGZG40VYO83G1qB1hIl92orx
3FzFWdY2bgkmii1MuWGyc8O2438TLbrdQxsk3Upvte3nmtuAFVcM8joG0Ih8Q/sgCE0W9k0ppQSk
8ws0Jjrps87ZOR67YpqkRDFpINIES8dxuLmsIXFrTMyYkNsNhyVaxftwlyas1EjNUlRl5SN1dFjq
k8KZwVBSFMTW2kXkuWe35A2WDF0+ZK2ybvqbzrLPGAxwK3jnJ+Po4qgHYbvtFcoj0ooMHVq7GIhQ
cO+Xj6hh4HiAMkJ+1fg4xWeBzmYhsD6vJ83x1AtUOFFLE+gtRM2y0rkCL8meQQXIYWTlCObaKP2L
o4UHnFxZF9ENJUtqUdiYrvVDDkKNzWtMDHXFQ1Zw2qL8YO6CaX97QvqJziazPjBxswOfjefXyG9Z
ykItVsCJb8z8lj3nc/LlhJprMWvsIi1w2KKqkyZ8vqKfDJvwS5wLHtrzi0Ll9ywixxD3f5rQSzj+
MYmttZzfXBrUQMpdhH/kOaUmhOxQN0hk8s9wEoe6O4KcABwikBqRP6xLm+0BU5yo8yNA0/FPXyh7
WT7eNQSP9cEvuuxSvWZVFZzWmi8Xuc+T/xXX0Btjp2PbA2LI6+1zaENClyavSFajjE7izWu2xvxe
8gRs8OIFuxG7YWkDq5abEDgjBCqxWnHeqqvPZaY6dRliG0Ki+tWVVQpFZQMexBg8fnzpBLra2cRv
VnkYo8KAvIPQRiq4otCHdWOtUXUCKmuURlzD8Jbdqtiofru8wUtNg2NlB69hZFap46nY7xEvUIxn
FpID41vApNkZ8JOsvZ98Z60jycnV09T1swUMf/3UQJXxogpA5j88/2IClEv0wyo8V1CITCnHQeQ3
q2/Ko9rpcwD9nIJU64k2XvUINvlm/W7mj+hYwyfIyNdN+aFH70SYY8iOTp6J6IdatK+2AixDKs6j
09miZJYCvl3xhgQs4HcRL3qw3GPdTiagLNEjbe17WcT2oUys6eAvbafSf905UMXDy+eOFCndoY3b
NCwfu2BXlMudQOsr7+e6a7FoguoxqqEMHl7a/zMZQbOxn+7vL/37glsx00Ar3ty+1hivaWNov9p/
jQUewDqSL4fXQ/hQd+JXALcPBdgIGxYuh9ziaSEmE/88Gpacb+7HqbatAZxnoPj6gUM6PpxKWaSh
oqzoY8x6cVZyy1REU2cLFZhdreZUujmXkEhSz1BULMD0F7/E+aNiZWeuXfzfDAC1X+Z2Bybf3EZ+
EKWNnJONyDArHI1oRXwLtJcuPiwwQ4o7dmrHy535vM56U4K8tRe5HAaVWWtzDQJFPwe3CExB1H0j
HM48KBxX6/yiuslFc7w0ApmtzEcxkPi38FnEgVNvAcTStWZs/n8Q2JsCM0rngaf7NTIzy5kak+bu
zhv/oeylKHOOCb553L9AT6NUVcvUrIO8olqKGqOW8/piE+DopTDUK9WZjGEAkYkhisPJ3HdkeRfP
qXxNJM3H9Vv8fiSgJEQlVMOU1r0+h1gTl7ZY/T2gaE8HftbqKD2xIvAECCcdDbUrUQVfqf0AkHCO
+ecio4do3Kk9eWIQPPMDdJ0/S0j5mQppNWDmgg98/2Z8pz6VMr+Th6nGzMs7y1DzW390fEzpoDin
aUfGnKmBI+y+IRkjP6oCYribPzf8QSaXOl9vUd4Jy3KBDgc8MUQVPhYDOO7LmGI90g0hTYr+aT9E
KgiD5AP/hHe5J8X8KM04LmQcvIcAipH5Xhg0sShgGMdE9wTPFFpT9/h7FBkvu5CiLGb6XonHntAy
7eVZ113qaWsTOAXyeyHgfezU8wxcbo9sFS3NTKXv2ow5QhGvBrpSC1gqVJ2y6wkWRrfoPv6dvWMM
6zQZ48KY3v+vwJhEYADu6vw9E6Gg8WaM0YnR5QR7A/cCGlKhsilWrIZ3SEknJs/i3HxDUf3pJEBs
/GLOZOLTLlIuN6jvjrdJ7qvi1odI/d0jZ8F9Plbx+jdaM4JMaJgRCqVrG5iOtdQ4Pby6/mx1uJJU
4MWNI8L9VpiLV+h+MgnL4fNhjh7sL6d21bM9b+emRRKJ16ehNVFZUZlJKyhgeOtTL+OZpIi2QYhi
FmYh0swBvUmmJat1w/yvHHaJPpSLGOHSImcAbHG98Fo5DcNztB+30PnUrfS7k0nGBdVZ8jB7vpA/
p0JhceIontonyBb4YH8JW9ntvYlgwdsFFfGZhxY1WBmRlcccIXzAx8elUaPsYx8BSJOQSsMHDbkg
CoUM2M1E+Ln1A4SQ2uA336YoZ4yYda5X8aMl5ixPSctqt/jW0kGpv3fc7Wvk5lCGzPJzkI80P6Mo
N48euir3YEoQW7WdAr3W7WEcCvMYMJZhXXwC+sGBVSnBJmaX74ZdXb8fTXiFKE3zsNXBBmfE4oQX
WBF6aIruX6uFbx9nEkPU68REKlI79QicRu/GXv+P0SzucgoAEE5sXI1uhCgcDTb2+uhxPs8nVAKo
THEwxOp42FvmIKd2ceF9hNI7wAayMVndQ6soNdxtW+USlNkawFZnFIYwbD7CLhKWlXHwW5PHfWrz
6Y5BZCQuV54f4C4lxQXmh8gtRW834SwI6rd01Lh00Voc5io7sKLnUSPTWScXash0EdbRjPtjtVfo
i7OPIpS9LQ3mDAM9WxrlPFZKUqnvCecrMwq1eUkA9Sf5k3IRIkKRCwR2k42Q2kfLcSNwDdhJQ739
Lsu4XYZRY2tTLowruS7AxLrYbbVoRyzBUZioopa2s651nY/oQACHs8sOI7YKCufDiALh+vlXSie9
0myioXmHv+JEt5O2C3rkcP4WDIhybwA212YXoSAQx4EVqfxVLqFPqz2oXvDIqIzfxDFyAqQ2gfKN
3Gd+nOP0X9TvsAw23rNCbWKgiwRo+TjMp4xAFj3dq+lrpCC45JwyRX1qXUhHm7VSHs6yHCeM0Udj
VJjanxf8sWGkAIlFtNS7pWgDkSSoQnNd6oWwj/j3zSqQoWX1JbpRYYSAfVu4fyGEdbWIS3ZPnoEP
WMjfDenDMg3bVx/So9MO9bnEREqh7r7ZhXt6KN/U/By6i07Lwtx6y/o8HEcG1eiedo3OHotOIxvU
t5vy8oAVrPIkGDVw1Th00eO1TQFllwbYiVuTOniVRKtvqOSRsGl5c2bE+zUzBzBtI2Ir+hrtvOgw
3W9eQAchAvrtP+LZWIeJQFRl/+ztTcxX3FShMKPftfg0Y6S14Fvy5drMIGXh0WOOXN2NsDzNENPt
B99MP5/vOATWeecPTVPMHrJwaJJiKmrybVXUnv80TlILm3WmDqXERSz/4Mm6mzi2pz4f4VjMUD1g
RTajGMNYUTFDvAUDJljKQO3iKSp6ItO/aygDMSXQAlSuiSLa8fBqPLWZFcXIHBfrAaDGC3+TNm/I
ZGRh7qOu0f7MeZeLxCpAmapykQjE33u4hpLoJa4ozyUWPYHhjgiHlrlh6vmhKYmjvQ7vWq0Ya4OX
7ESCyBqHJi21SOWWT5Q/i8DUzKeBSsVrJlWKk13qKkJp1P/weP04J1e9Jje1/hFD7iveHTc5bKsv
DGczj1r4qaS20U3+9UDTt6+hAIi3hWFaaCODSOg+rXQsmQeODjmIjk/jaSyHxSgdb+XqonJL2T8w
9jhiIZP/UBhyig/dz+UUnkGJTJdF1MGNfxjhV2NrZ7ET5xTmjDGK8CCdKVzGMcJMwxsQHmJ3JWM/
acOHB4wEU8xNp/CuQyHAlgUtVQ2pDDarSD1viUAPg0/EVPSn5ceO0pXZzH25ihx6vNJafTiImVVZ
CwxxAi1RFkws3DtBRHBIv5AftsQNkZI2urJXpF4JzNYxxoX1qRy2ArMP6ccdkB/jT7l+UwVqjcaT
cncMvXKEYajERGMwxv54uEu3rRe3aydslV6dXqCDjOBahK8AddG/pj0wojkmobgZOT/jg3to09nF
YwwvU+dIzK5sEGE2UuX7rdB1snbqDbT320Gv7cMi26s7fnxDar5yY+IRVkqWblvnJiTzmKDYnz05
zbz7ivt4wRJqOOcEhLxECTXM2+JU7NZOjLmK7+eQFhWYEPGP25f064MQylPES8s8MVYwEFyWwiMI
ks1qki2PQF37sd/XH485uqD2L+4fnoD5tyvu3rYbwef+/awTrj2ngo8FcbNPeyyAmsqylVJEmKdX
HVKMrkC7FJOuFNWrG02dOK07UeZzc13TlbQ1kmrjz8tERqXvFkXL88BGY5LYuhVa0j5+f6lqFbpw
vyyL/1aX0lqP0klYRjSed1ESLQ9UKjCJanmlCDqEj/6xGLvgDKZPcooQERToq0mwk2LdF0eh30NN
1ZQ0NpABX0pyqpHhJzZst0+qFzCMhGd5uiHeJa6LyBM+U1ZVn0qMo05pPdyC0J3G6gHPSpi8AIfN
UGjMVbNYik14bYJ9JLC6XP2GCtRvWfciVltKvevhvtaS3riSBMZcFtLEQl3RF6AZ40V+b3jX0SJj
n4afmNLM+8xs/DZqKc9zTK7sV5R99EptfKNT8uJCZQkF2rguNT1Curt55oqhuMeZyUEdMNSNeu9d
a2kG6YYsrf5B30WJqGOp3gVGWZwYqXpWfz6mwkfLAP2UUlyjHyAPjzIhKQg69GdMkx4TopsDVXpp
hhUkJSPGSIaqYVHPtUbEeWQrkpZUL8SZ+STZreC6wUJNEsQEZL3JTnqBHtUJXtUvl1Uj4OYl02iY
QH/Y/jj3Er66TVe1ChVu8GFJJ8UqYjHIDOiJkOIYniPCRureewBDZhLZWmrYXEb2d0smNhcR8TBt
FQRvaYliKncLcdEFtHJiNtEciucpEAJg2Wru4BuKVShT9KCG7PwQS1PXd7beuBmSlhNULGptFtWB
mFPvkDez479DMXXAM7byLBUM+L4/8E0cr2T2FWrko+mWxgOQ0s86bR94+SpIVUQeDDWLbKJ86VTo
KdfEwFHmdJUr7NR5TFcmG1iVufgNIZa1FAt+WwvrFs/nEGZKazIXOMRMFtN6BEsQuS9gTp3I/EAq
TIlExaULPh5Vbbe7oqA1TjVkYxOKRh8u8iraIRhlr0aAXg40+HR2BPhJM9P82BApFBcj2pVarehe
Yure7nWo8STYRlmvCE8kkFIlaHHYa2bF6BJ+6oenTX4B/fzWqc5rXWwKDq4zp8irSF0jqwwaFA7H
A6BIoxb1Guzb8YaooMLbw8Xv6MxIOBvMUkOkaiKCIo+lBcfqY2A6TCRn7pVyC+vfr39w44C4ICL5
WcuT2uQUMDiZUFI11M4eFZpNCRjZNaiQpNQcKcuIIor80FT2Q2uT4m/CXb6mrgFBvG8NCmde47mx
lCa1K/TYQbT7whnkD9srK/aL2pY694zhXafjOuAZK1n0uWgKaOo517v1vlKV8F9HG85juY/KHFqT
TFm8njJfwwuy39R9OFu8BR67g02Fxb+YjKBSa0Y02kqYfcLwkOhqmttiXrJh99Ep+cREwD4zXHeG
wdq1l03sE/WBGHwA8Zr672o3WTgDUUb8pu2keuHMKgki2MMqbetEpCA/ZJSEn4ticktqZDb9qZev
sD8ZZ/wKd9eKaWlswChLYoLqgZIF8W+RfSi7U8rtMfPchdO6Vnq+xt+lvDQ1d12pZ1QekeBXfeNZ
brl5VmomBImPZrwQK4LNez+W2wvp9klyI5Bfp7RE6BbgnrLuxOiEhLmYEZ2VEc4RLyO7m55mD0BN
7GLxl3coWKpEv8Je9UgCsadBMsHeTBXqVIPFp+m56droHqJ1MzjAVpkBFyeTo/Pu2/Fn7wRyz1Nr
VziKIfKLAyWMJGfE9vKy0m88iHeQekQBCmenWW1urDE+GaneHtyGm8IdNzWjFVio6ofkX/52a68U
nls3XZz1cYFjWU0BzYuZdBpp/pXVnD2zR09ZRrl7BhJzxglYsga+ooBn9W+v2kMMWsvWEVKimrAM
fzHbhUasjM/z5P1jzFIug+cBfVvFYM2mqj9tXUvTEgUAAR2BA/szhJizEEkRdy6+r+3aFxZMQP+a
AFOktkanuFSt4KbOhE9FveN1bfUc6UNBf/+5fO/Bdiwdr3sWvYKHTKUv6XKftKauPsJhIEUgkhjs
rUZ+GInktxVSUSsTYOmrTrI3OThu83un+WQOBGb9kb8UAAvS2GFQs4sC2UbsnqJr8J1Wt7aTgxQG
864mzqw8f9Xa3FY/FXN4V7+X65dZaKQ8No6bmeIsui8REe5Oywlxru+RElVzgE3Pf4NVt6wy1fG1
Nzo2VBrKP29IL6Ntj+70RMfUKJoWWGLWZZf2oWJ4iogtyUZRzXHhws50nIMZ4iIgaFXgd+Rm5H/1
xAeBMjWYnYKTZLZc9EGEle1jtnHUuv/Z88HKyn3p2rlxZzEN7T8jhlBOwmrITrvaqAFX19wkt5us
+rEB3BvzTDrGXeQaCBj24Kr63yT0j0KrCK+X5NoJF0mULDAijceh75O8IbsN+4Kl/mNWzN/3zc0d
0S6M7d1XTJaTh9754fEKYGCmcOukUuijXLgXULqPn1/AcpYOapGWfoGiWuSIM10FmiN44yLXkS3k
x41nn3emMEgndx0fUv2ScubUR/WHQQr8yGGcyjdFoVInOpZxC50QqX22GNfUR4PqI+s0TC2gGvwe
6x4vkGjrFHvjGI8s9cSGCmFv3L4ll4yYO6v312aDrmOpujsP821kmImT9ACWMF7om5rI2eJBW8Nj
YK75jlFXuvfkLSlKrCUs+Y6hI9qasn4t5dB8HOcCvhKZNmrn4XGhM6b736p7sWkOxwtSJFggn5Hj
h6TuidIpXEHGDSFghJWViKTUy05UlGdpSBSZAA5X1ZwO782lh4vORQum590UxwJUiCvGHdkxP+rF
5ATTNG0yJnOX8lUvQIJmetzULJoKJrUve9Qjjxyx+rH2hyuX71bfoGDiaxShSlPUnP1Pwx7iuzyg
FD/xlRieE6UITT+vccB62zJ/prxxR+d2BhL2TkOveex+mqNOLBlAQUo4/S6M180dLzsyQuqeznED
hCPa5ehohVSMlnnXwsGaq1OtnvGSXlzUSUaurgUzdQPqEnU5c5fmEiEGYUTLGyj5XxlGz143SO3b
E8+9p6z3aTYjuS9m2TzowzM6X1WMpuDAV3J0RE2CjMCwILxx+XP/HS44eJOnh+kk73IErFnO1DQk
k9e1CPrIEjjre6zb93LH3d8Bc5HqH/TeS0yRN7cJXNe3wZ1JA/Y9sJE7UefTn9BCZ4a0ZG85U8Ut
hBw9klIbQKAIia4n9hGWc1KfBBIpXa/OpGQ6n82/+5/S15xsRZ0tijvWMc2HisMXZDFYhlWZDn9f
5HDWVSynzD11rBwpT831zirChgX91zA9gUoE/wDNxM8SvrPN5550SEXtgxylC/2gUI5Z/tkz2YzD
SkzxeHY+tio+DNnAie9hhO2pg6Cg4ULEGn/O8nNWVE4cX+yRoQDza+yWiktd28wVlzaO+UXf8I6r
qRbtub/4qFxPsyEbhC00bzbU794AyfBLZig0JnKvdsJ9akZNSPkbaJNoEvsPFOUGcbDSczJQMTRQ
p9KwXoe1Jhiv8vlBFBySMTkBtOVr5qQPR2Z1qeCrCgiNFNJhad9+xC4dwHney1b6IzvMmppMbGJO
WGI9wVFHTxq31eWbbp2sjm8DAuN7xZvkBtFtc+bQrpi1nuonocWlwVXScRCk4ZpRPYA4AV++NwHv
erfB4U12TktC7lcSXXnITd3IDYFSHReCT6tZO3TRbiEEVSRvu/2orqhlcYmBzPrkRKhIzMt84C4Z
t4AC076fffbTRx1hLPPoZWXA/Nc0s1Lo2hHXFp7qZVZyuoytREOMdQkScnovq5WEuKmQ0Xap94G9
6zKwXTIx1qaRaKCTTRjZZZSuTIi/vDmNZC2BXjc7vAyviHyEtc9zcv0Esd1TQD0gIODYOYw7xgNt
no6V8yagl0d3APG/6Lrh4i48Mx+m9hYogDM/POM7BmXIZi0O8bEYB3P7hr1M0EkVUmmswYh9AyQl
Z/A9R1RlRVlsFevL3DlYqkcBiLIQlKLglS4vQxZX9OnwkrxprzOSQt91tB/54b9Ynk9HnWrfTq8+
eon+fTEZZqiK+CtQEhbaiehVHyI4geQrvLibHMMgWEARwD8lYR+mEb/Ssw+4C/N8YIjvugCSd+R1
OWvctrepYlQStUB/Ak4p2K3t8nsIaXQ3G8YqL7umUk68nd3UosIxi29nQjiYYRBo9RV1FGP8XP51
8t09UGpxRcmNoWQzfQCOXr84Khd8PWVk1Gqa2PbiqzJzaB6sC3A9KJef82ykWyYfsNtQo/sLf9iy
REf5xdsVVvztGnD4eTbErW6d4+KWTj5fJcipVmZRpxxJJew7gHiGQ7THHMqEVI9UzeDwzoWwI4rW
ZkATD4qWJrpfNq8ULB2BUtJJ7PyDwDpqL8LBk+Ey+/Fbo1nd4GycT1geDKxxewkLjObGJmTfjscI
6Ikw9ktyLV5v1UDcBkuVGvwZ1aKNgQtRfwar5WA8BRZryOmV6J2n0D/OoPgWnn3mAFDhwph9s0Kt
r6yTefzlapUOQaWamtPjWRi32XQb9TP1LTAByabK0he3t1DIGgi8/BOBzyzd/N6nso72r3FwaoBM
C+Tpk9D+hTue6K1QoOyrNIVgKLzr4wQl1gdI0ZNhckrQV8ewH0JV9YSbGWs64qBkcl+PEg7iYY19
OttNX/FqxyN/c/dbKOFsUvjb8BfudAJXW+AvPiOeByVh4Hsc2SOlWtRUq7liDkJYnqwt0OYikfwW
J/67ut+DTqx7twX2b6AoiMteS8Za/nhsQb60cEgPE/jHnQ3+ENEwz9IBfpG8G/vXgpPZJsRbsktb
4W4TDdpwJp0LVebAeiJyiMCXOdt1etXbekX/Re2GXJdoCBeT5E8l/atS3lOgOA2tPZuRSR835BnZ
9tnKwcPvjcwnMRjllNVbxZ0+ec/DBnhi5vf6XwjGCrqPpsL2+C6rGUIEizEpX+Zhvnb6h0xf8MLL
C8/ERZNB5/Z+sp3hI/Vmja4q8TiHREZ3z6dZ5+1quZOFVT2j2a76hejD4nl6ynRwKoUR1Ubma0wj
6uIVNn8z/2CxJNDb2xMa7X4ucQa4uTUWHCsI5xzKFhz3llQAcdt4x5+0i9h9PXZdcsy7t4Fb2BxF
8QjVZLm3jYFWKo54yNnsVWIyV3GGt47ZGE+CvM+azbQkasTRQQ43T1P6RjfqqLYp1SaP8YVP3hzd
xhF1DTpc3Ku+vQLzT9HIOl7ijllQPqSXkr2M33Ph1q3Qi0cn+rfDiWxO/xHYfqzFSZtMuYie+0eC
qbmDcNVZrp/RSknxBXOTK4f5mGhoux7NJYE7aaXhPplwtDKWmxGXz4qlSOdzqlniXShmzGKowsiy
CWNxIC5vEfF29tROC+GgUhbhEQdECrciGMxx8Em13sMudZWCdOrquai2etBtNRRDDvxk/8xRrr/x
XxJgqj310tnxZmX/4RpZTRs1O3oUbtqAQkcQ8IWYe1XTm9SZL3I4hgwhNF7ZEg/wwEbl97AoGqAD
6loMLrWU1TiVo8iBx1HBWyw6rcI38J8tFB9L2oXtkTgnutD6URdFfCZBcBGWCmV/d2fSZID6YWFb
4CABL6b4T5Lc6BCHJs7hQw2Kfo9/l+HcD1v3IL3fJfjLOMhWs3dKDGkC1aFrUMhZ6KZ7NWl7Fshd
X55ywes08/oj+kHHCs6TQxpY0KVr+UgUi8hOxeSZAuMjbCZ6ixjBHbKHxW8xMUoeqFX4JTlfvcVj
h0l0BZ6q54Nmx79msSFL0+xB1Nfs3PNsvrgkMMJbfFyh35RZ7xgyWbz/tPN0ciLkfv5mf3g8RnGF
GEGNnv0Yb/xdUcwkCwiLGcA/V3PJBc3eSSpMxp3ZYXDcixbi0gJdQaojFdkfTsDZhIKA9LRd8KW5
rZQBJ8ViE68P12rBCrycbF598mZEMH2AXDR0yxoDjdyeqXJ13ja4RueVK6sIKRwcKF1XPDLe/078
3IQAenHvl3tkOrWuLDEsNcAPsf6RBLG/0MALkS7ygSnKf+EueLAyWOznJ0K9TU2zp+uqb4N8XziQ
bfoBJCIiPyWpOaavJEq1bpnefufuDlxZRmgLl47Rap3YbJnaszOs7/pLDdOjmiLD7o+qPz/IReNu
nm6RHtITDl81aZt2KTvfh+Bmo95/+5+OI/4c1xaBs5re51O1rAYC5RqoCsGZwkJzugHlso7Dwyi/
3X3qByZTswwNGmTMcVVVDSmb8nIZtkzle29V2AsW8WtaQlhXI85Xu/RqwJT6Nj/YDGpfYugYMvFg
5ZfUNDfEIwudGZdx4K38aysd1YCSa9BzefCT4+kk+2Vca/zVLfgg1VmztsTFIGl1lIySMO353Vhx
0ohULmysE/P/5e1/KxS5Pc+EIhkHd9+lAJF3gkKkpNXQF1dMglS8fTagYaZJJKxhlwj5x3SDk6Xh
vdj79NCgyJbqInVEQRJ5EII0LQoKsoD4cxGOcOeAXKOhieB0LuoQwAPy6n+vU2I8kLfclnGtJ6Df
A+R9Xfc2TfECVOSFzgCa1VvFFI6qfz7O1jMEwbwEl5ZpfSlKjdXRkkn+sEJYevsyPhOcsyT3sf74
ibdpF1aBeh0IU3x3MzdpoEqBjWLAUUsAlY5nu/qXoLeMFZ/QyWqVtCDuv4+ppvy3uX5EzLMFqQ1S
Dd9X/BjckhwGag4ya1f23Y9Uhvt0yyyXKStuCAQqpGzL8uE7MzekZoQ3IQMOstJ/F++qUlsUkLcB
fmWe9n4KrEBqdU/DZcTiu/uZfJ3061w0UtxM93j5ACsSxJ8MKm4+d/xpTDE7sgj5A9kCvVW54WGP
OpP8/W2DRiiKcKReOt9e+TB/sGv4IE/t3Rf5K/fjwULOS2yQrwgiQ8Z7n+H7zyCEypH1N8ja1kIc
FUUITeTcOKXBb9KSE3TU2/3vyTzZq8C4BK5/xOKg9MfBALBZELgYs99JOSzKhGwFcJl9DBsQtIXA
koADPxZV1l690rI4whJS40WtwIenPnU9qbTHGzi1wB8tq11s8dMrZAA/+GvnmBffVjxLGImxz9KC
zXOc18iP4n3oPJlnCT+lVayLhuS4UQaZWQeT5va0nn5zRGMLUMvM8WRUG0sDwXcFI/7xE1CiymCN
WmmHW9CAfBZhngosyh1Ggt9mxSUT+z7NpMYUu1vo4gAxKIYho4st7tKrAphsYpNgsmF5uhc968To
CbxlH2OuPbLqNRzzIg0sAfXKmUlccND6JzDpzR8jFdpNiuV4gk5HbNO+Uy/Q+cR+YbwkYEtbQVMO
OwqLYhybujIZ5xlyD7E5TzX6nJGPLCJU131FFWR555ZJZlHZ/Y8FWMgfXoTGbBrqlesJiNHLDaEH
ydSIzLVGXsMe1ihmBbblEHQJHgLLFrjWAugoTHgSU7fDsIwuQHSGp+xHgoOC9BROrIkB6B8ybTJw
/n0YEFg1pg3YFV5QX31/7AsiUONJP/d6OKSuEb/lWfsHQtSxxO2jNTvebNcW4c2yt7MRLMKfIlrF
2oX5KutJ7Zy2eCkwOT1BVcDjhf4zgwdUbWSjWe+SG378hrdgENohCtyQK4vmdxi5AmbhZgaHf9jp
UXBBiKmfXXX9Iw0oFb4Dcc6206vHI8MEyfVk5jIs7/xiwJ/X0ecYzVr68iMS8OeViQc9PHKL68d9
+pOQyK7WNeDjGdqk/baZgkcevNhmwKCOrwhT3C4XaXee3JfI+pAUXAaSPlpZmGLfL108zneZ9LWS
h+L5WTZV+QsyBS/7IaDIXCm/WywL0kiKHuYBRqtjT9gtO/q3AR8unOz3HzqYUFtNFyU4A7Vpy7db
oCB0d5WoXfNuuo8wnpk3fVNVn0kI4pS37mIS4H2IIVysxlayOzT2NRIig8+GbysZA23YCcFJqL+L
6Kw8Y6Ys9gDyi1cM4fR9XdQhhI1nqr+5DYEPoxgjDdl4GLXNHrz6YlzJe+70+x5AZOsJP5IKlqnM
mC+LQUoghr29ec+79s+drbUVNXdjuN5q6VCeHcgO/Uf9NQ2qNyyEqyHy7+M8T6WduuH1uXPUPTjB
l5LEXDPIw8ZrZZo57jKbS8oA1U0Cg+ny0rcwUDuZSD4VaIRP2KMIGy34KzClUhiT7SjER8Fh3r5h
Wyz+mIWcSr8RsRMc+15GqCTmOk0JMhgjk/5bLqdv6lEqyOoxnUPchG340x+rTca0jkoslJDNc4DT
8pskRw3IgTTOcQ7L5vWaJPAzRuJVBdfKlhJznz//sf79mJhgLJintiEf5RCBZiSTFTEuRWXU6hAz
uYkHU96CG/WWUg5PvaXvz/U7KUNUQF7P9l3of1gUeDqoDyOrKqEgxXCmVyPjcw9z8w+LedWBe9yY
bwhIycCe2v2ofFJVm/IT7HXmhmOgox49wswKwzQbu9dE1TrshJ99duaaMyUhEcXBS1BSJ/ooQQnk
Mp8zn+kcuBWYVSEXWVJDos+mxLDSvvWicoRgVqR52g2iTs7vbKFRfNQhEvLJ0k3ac0dMNLPI0q1s
peprCaKUI6Wx7LlqSUKh+K1jBygqcEf7dDV6QtKI1sg9tSNlyBjRpXolBrt9xE9e4Bcd2CVeSRWy
W/pIfoRruSCpISiYn68XC3Ppe6FkyB8P0X51UwUlxyTzGEV2iPWwpg8IUnOnXXZbKtMTGV3yKeIh
arstWpr7gSPQmSKPVjmqozpUaV86phG61tuhBdPYbj8YvAKlhynhnL4/5Z7EsTxpjqWCLf273w2e
IT4eQitdM8VPqf2jTxx9zCFuIGfE+1U55aP6V+vfSDsy6ongLK8Osy5Og52/EyGn9gJRKLLRCQDT
SpZrUh/tGRD3FSzO6ZKzVNji6/o9srvHF+OT4X5CmK8nlhTwdYWhorwv1EfTnEQt5gFrJjUPhLbi
AgWRG98Ba9G49P9RibGOH1awhDkYVCAGyIYH34JFjy32O5Tcy9y/B0PrNI2hlcgwH2m5gHxFjcf0
Rr/0IaEIS0D0pGRMMG6kAD1aKPVu6Dp8hu/3xi4OHy75yxhMwJ1m+03OEDU9fygBdhtwFE8PAyCY
xndCuPeIsFx+9RtjqaOsgejnThdW4rCoa7XF74Z2n8vdyRQRZOTZEu0dnlaJsxD2PnDq8jAz1CH4
3PaasybnUpxBF8VoOZ++unVo8DIG2dSWiTUFnAzWwUBXJ5BqQEzj2WHLRV2ZUyj6g8VqCH44A5lI
4JFkPehczQxIjHdh3JfKPAVAstLDaPvxQuTQyjxzczNi/IXOOaPGbBk+CTN5jjixw75SYvqzS9n9
w9ThjPMQ/gb9ww9dTsCxvSvDXyDXo/QTrOJGDxt3VW9yN7b7dLZ6zoXYSnGf+OJ11El8T9vc9Lby
lh+tPDT++jVL4710xmVj5YJ7dygax5i75Jp+P1fgiKQgBIU45FFhFKh+Jim3kJwxCym6KmX6wZWk
6LvLZvnl1T8RUrdD0DtyrODIl+/fuflpJKL0amOfBKb+H6KA/RT4Ru+YwMqc/0o2BUOAWWR5gtyx
6LZ92h95vFY/FQZDrBQnH+BdWuo4Q3yW0bDZVmuZrF5z5Bx9HaZ5mA7G0WQx196NoYkxHK1QnHdE
/gBeGTbUzthAIpFkNWfHVtoTbYXC7nuajj3+/DFGMuHx8wS0IIloWv0wQrNzOo9jJlnnKXKrPktP
UNFggoo1VWMtUGmvKXVPosXKViKlQNVtzUdsmmMU7Hj8ePEryxFoKm7LMAvJAWw+rNzEKpOKsXYa
eHh5uhT4HUg0A3NEcEjwbKljow3/9Z83IhqR4acC3Yja08DO9MsucgBGZxdPLojiA9K11A15VGaU
RHe5iih7pDxC61qZyh1q8Zk6Kyr5quq4HX2xAZp/2gcfuPqESHWi9PSIDy4YQHWiEsU70XsJk/nU
SnoQ7MmbiJdhXXeQ6IAbG9se5Y2VxUxY8HsJx93dE/DIHZbcg6FunRckR9w8Kn+bgLBkpOe4JmCk
34QGcf0sGmqpo5VXCxeeQWTIHjuZOM4PD7OabWCkwPrsUz8S8E1j2QJiR2lMzF7BO+NA30RjUwqm
vYCBRRm+dK8WqDxCnAE4jya5kiYQaYN9qMZ+TbVfao+je2lt1eh4lBtO4dSJ1vW44GBn4TIiClbY
QkiQ7Iv79+q3bd4JdezZsY6H1jMrfSITIFjon1gXfCVPDj7bxsbvMH6zxXgu7Qw3AHXTT9DPSN0M
O+qiZMigWrlHRxflzUY5PJ5QlF40WioRu9RSlamm44WhEoNv5CIEF4tx1OsEjwzHJ292j3hPFc4r
lUbFquP86+4OLq/LgrpcH1w8f6KV8jeLFxn0K4Dy0AqcQrcWY8G7dT2rml2aRtl9/9yXw20hBBLe
RHKWIxhR6vVKg/zyAGLcT+QPKQYJQpvZO08e7sWpq+fkgL2qIOiULdZqyLI1qFAICb2EODJP+g+H
mzQjysHCQqVsu1ri6lZGH65D7RTCEsEU6YJeFMMBROVBVxnaMHSPjYTHFOjhMNcn6bvFZZuvsSEP
5lvw+S9ep7HPnK0trOnjqwRzjjdRJsJtdHULmU1qwiNETpk1yS0jvdOOipQHYXsQ8Tay3I/+tqTd
sYG5J/zUKPnC+kGs2m/SrIHqQpxTgPH+oQEpDS1skRsmceO2WaB52UWU9U3/BrVBseS7jMz/4c+A
Rs1B0G4YZDd47WRvVgCQMlLTzeoew8I+ozsxdpOqvrw11YkSGi0IOtMyUj0tiJ31j/2wKBp9/c/V
me9LOmafq3GI2dZyrkBAM65hv+M6TFwjllFkFKSAW67nUTmRzBY9DhJO84l4JQwUkq7iwnFZWsJN
J/vSwM5wcNAE49VTJrsfd4sO9oJwWp0bFOqXzpSmsvtv2EhHxs89gi5b9PSdB7KUxCiah3IZmk9l
S0Wccx0neOm5PaRuTpmqcEFLgb4ZxE0UBrtnDMUKQzlNebK9EZt8gA98XrNHhTnUC1iIg6NPInwU
bb9615+D9NEFz08TIUct2d516B2RpIpXe9/ul6mCHSTbczCmPSmNqLKReFTU9UPbdwtEa6ICWBiq
8QYe2Vef8h2/TXb+hXJqvrAZGT8ZGjLed5gFaAAtkGybpeGFrTYUPULdqFufasVnX9TbQmHtDlg8
H+0qSumqtGqPgjPFM4PU2diU29YOXBACrd2HR8r+em6JCWMKhJH1bqcnqJiT2jm+KZJ5uyksOvsB
vhX/xQBzyFlgmoo58wSU/MKPUyez1Owb283keimid1YnFTDE9VVUsfHcQfhZ2i0hhoPrXctyL783
gjsUbY2r3WHj54DSAqmCvJMoa5S7PvNm9Gpgt1m0r4mXxTFln6gXzpYdO/COtuxfNX401QnOivot
yqVcjey/5wUANgGDz5spCN0mzqCRCcdjNEEz37rC269zUPumQCamBjIIUuZBuhhJcgbbVeywnq40
3nFDz/l4TmXe2N18NI2sazvpUnXuot3wP53LJ7vrl1AIhFT3uHXGRxKaWK8+689PPLA+OyAOnYxt
iYsUDaVuUmHQQMWUfFOPdU3Ds+/tVev3XsSE2hD+G5aFi3KsxHXVUfHgr77+ZkevqmSW1xZzipxq
40kytuatK3niQOTSw/WdczaQedL0m3X6XdLeGXCfAzQbpDvmG6UkC4zJoRUwXfxCsLp1YVzmegcX
BdjuRm1VfCweJtSEDZZOZ6CdDyc2xJseXz2bcXzwqKbY0nBC6TfwCfm1nU9ps/mu2vdjNvXHcBYN
1USwQOA9JXJx7hiK9xX2kFKdyx58aWJQgBDPE2dB79wyEw2ur1B7vM9yN6oYTQtQysNC58XERlIE
uv3KDkhveSdfU/xK2vbCxx3jKtbbM/mJsu3JaZAHBdHG1nJTRQgovwGTtOkFELWO5UMlnYjKTbAg
oAK9E6sgHYCmQzPTkUPO9FTCkWSjAgdSpYMzRKHdU+yHvgCJ4LgeiOJq47jq2kmdOd9tahsy/fUL
VytDjYvFIvoxtwzAM/7M7m1dE/wxOVvMb3TezByg60GhjR0DXKrOGHMUmpsgESf+2wlPitdfcCF7
0DKjaW28AH4/n/c6MQx78BYvylWWGCKYQmofQKQwxy33UdOTXNoOuPV2yJaoxttRvsruT5uiODtL
e3uSGtjGjNFI3cnriXjZKDdQmg5fTZV0DGGVvB0KhYbPm02AkoW1zi72sLSFJ1DcPMEz8Uutp0Pc
Sqhq0LtFb1g15FddH0qhKBTK0uoxIt4CD8Wu6ZIZWxSCerpOvYFo9QNF4l2iMuJT0jLiDDQkiYUg
jHg8XzRg3aLu3543GNOLIGlKtt7b2uH3JKYYNEVAQWE7Jfq9vgMjuh1T8ml0+sX+SKPzVBqG+1MD
uNaEt0MbiHqQHt2iLpUiVReryUD7JSNTqBCEw68KjF7t8lSHKmxERmEx6u64ctWq4u3uN5pwayfd
1WJ/9+Y6qP2VIp6VWTxRli+0agFhdQoqeeYq/0aJdBpAf685vfOx1bvpmYbC+HFBKx9IdUjSBrKo
aa/f+w+nI5Vqh7PR17Wg2dXfe17eVM8qtuLNTCUdBpsLST+pl6MTlilFjaM37PkvJaLBjcL6L2T6
GYkcKUmWJWJ16Kgf4nL8nEqux63zAts6Fk13/y1WCyh9KkDoOOqDmRiqh9Njj9LWMHFtekv8bqdD
IZVICuamFk754bWA8MLTlcwSqOWDYJWEnbmgPtiojsjtkivTZkdHSM3HLLngbOslhmE6GMsHgPjN
YueWDnk/NJ5nOdiTTohM+6TlRIefnSdmeVaHYQQKImV/kBfmUnlrKmZGINMuqJI5P4p5UhqFGGIV
2oUsxD9g6VwvZnbM9tHvLDUN+VbxIqCXCkXZ+AaVdOoYfMidsFRXKVUCARxESb4XYnAhtc7r9Zcu
5kAjgDgH0P408XUjT3F8oZt6TtpbrXSUWKGFza5/03U0j2H+Gf/MoAB4/Iwm5eiNtCk9pGHNsC2d
C3E1ubi41Dvc4cggcq7PivKIpAO3uVRKuFuDp2kuXW8mkX+B1H0LnkpRgGOhjL8V8sfgRARUAKNq
ivC3YcnoTNCYd0rdoMzcNH8sgmyl43wg+7AozYaU68Cv/bnmG0GfFo1Eequ7IcgUzuSFA14wGP/7
ThA+S3wq+ygdaG9FfuXPhpczDvhFZ78nlhJQnVy2tWlseM8EvQliEzJH2oH6TYYN8E53rJv35XaA
s6EZ8s7/YgNhd1pi10eSLOzX/11dAUCDRfwzYjBckt+fVeoBvuwy4rIAipZ5xSJSaHJI1Cb98VBP
hZtthtrCVv56wdRqkoCY9HRDFRthS/QdrbGU8y5vA4B3uDueJOrnYsM71MMEJRyVfQEU6VK7VGAJ
i9mCuYsMnL/3pl4oXOo8EXPzb/LsLukqvbyvezwU0j5dyuV1gbxB7q/Cmi5U3K6s8H7fylfnHz2W
F5sIzLuxfjg8VKj5LzmerDwb5/8tOpAVVtK+7oE/hsRZ/Paz6GhlNGn3fZ4n6YcM8ex2/IEuFC1d
NfWv0bdayT3ggfxk+bJf2uhDpuSNyPSsstpFcPTgotNPQhYSWEO2Hj8OqDiQ5JbH2eApQhd7zKAG
P6ioQNgf9RT7ioAu9hphZzZG5qvF58bwPbzDQgP9N4ygIhYRyTkcZL5C7FI6l8IkfmOT+tSwbXNg
BBxi4H+TWHAeGtrcxMxvLpjycm3M9DggORF8fepc7IdWW/5SW7ki0yGjN7DiEXnN/M/PuizFKra0
OLEcM+SuDFRdFDWd+qyhNM1a+NxtvH1plxUwd3pA6FA7rQNNuhNwtQ8s16cY8ySkXUNhtLcRkyTS
ZCsitWfmRy2AYGq1qcrhEyfdEJrlO3TuMhhpiSE85JM2v3VmzHOg66+KNmdIM/tTsp0+BH+toPwE
KANuSaDDyq5NWi7pQdMpQPTxlDzZzOQDmY+qRf+3xzEOMT3TsmwxvDJ27qUuXp8hUiRweqJ/f23n
SsOTWGQZXoGDX5wQMUOluQ5GOzvwfaWjV5iZaU2gA8Pey9dCu6QazxaSi2rnBhb4wCMADcyzgqv2
LOJ6ejp/1A2i44d6V765JujbSZM/qYp5egrvpNIFbj3oMZ9yPKzQv8s5TtAKRkTmGs2efuSROLph
hTJRwZPBG39ldlMb9ttkCMomQMIfaaLlD/IJA6Ie0NHxiNt6WG4LktkcIPRorRVSb8PXszKXP+n5
llzMsw/qCxVnSewTE6RfVfZHCZwXC41WK12bxtWXFpax5clZGHMg6LT1lRAt/vcjlKPrXovs8Igh
xHQm0LRzbJ10Eg+D68ISOPo1uPzMvXilyJQmk8qTZzYxZD6exf6WlaID3xAOknQrSS+u23ipZBym
UnSc8+HaETaTOq4OLrlldAnifGmBQIQN1Ke5kTsAC3F4N2N45J4DtfDcq8uQ/VN9TcACpVxVYJZT
lOWne+277laftUTxSAgFjqiy/f8GIxPdLOGL0/vzFZpWNunutHdeVG8KibOaYYe5FC2ahC3jOyIl
h0LXMLH357b7z2b+IGBpIlrpIGb8aW1OpQlUn+L3Dyiz9wz0tlMtFv3jcBxhGsUdsZnCGqtnSUCk
hku657nX1q3kVc11mFGf7poFGEDd6YuNoMClILLnhW293LVICZmQ2OnenwgG6MifBDTKg+sXN80o
C5LFBGA6P+CE8SCDid+Sy9C4eIQ3XDF1/IISacRCUBUI4FVX0jzviRyNf3Q9t3iZ15p1/cTiuRu7
Z5bpfrsC6l9bj7/NuKeANOs+bsJlKdOulm27sKtKoOiN5K4M+bSMVTfzDIw5A5+48r8AkqE0Ue0v
quViFxitTTudw3IwRR4IiU50UQ7QSUJd+RhH/uAAlPzG1Syk7vdsXKpmkM3oywRLfydmHNCrywIC
bJLIhR6lAoLta/7Rf/1MeRj5YMhsgcDP9nKbyTr5Ferc9gEf/9P9bJJ05V2gp3JSFc6Yucs0BoY6
NHWnOK1krjkEIOLkVYZsc0BdrFkYCCVNOZDGtJ7fm5F5mfrWHxjyR9LElLGhKnsVi+9nV7kSmkz4
/+vjZz2YtokEmoUjfTOe7qnVm818EwDM1WiKQF5c0/gDgTkuuFYZTZz5swNu1s1+MUoUOEBeYiro
yHQj7M0kC/pLq8iQel6najUauQCp3xztpJfBhy+eDC8FJRf6EYIdOuUJPFmT0X1BhIdwgtt56ObA
pKCcAi9DP/jrWt7ObO1jwIoU9yR41sUi9q9ZUWVRcFSALyBTXm5iUhpSHX+pi3oa6Ih8JPrfI3rq
HfiQw0rGOuMpjNVBFta7rBv8g4UNjmzVo/AOcckwmPJRAyejZGZYm7gNvYtnl7KAzSuxWtVkQHT6
z4SRQRpn4rAlw0NtszQFXh1hBYaJGo05K1MSm5ZcSfCACdqoTqA3dzNxREhQicKeQ4J5lxeSqYOD
q3pgfhLZyoMuMv7eXyH5wKc0NHJ/XbRe/L24PCbsPO8hmql0iq2/cz8usPiLrYP8zQAni+Cpttve
+sWTGa0NDCFXZr7RUmqz9AWDDRoYhn3T8F0LLuhGiYbHmm5jMo7/Gbl2PFdAUgvM8ATsMTaFgCHG
63nzmbkams7NQEBPjOGrUf0+8BzBD+vmaMpfOdUEWpX2lt7uHwUpBuOkiPl2vPYTyRZw9L6MPS7z
xRQechIPHrPGjdmwZwbAv02SwITC6c4Y/68O0OTyxrvVL1qOFa038j+Dis0OOqgR+b7KjHA4Cn/v
3Or8uOM0ABpkJGB7jaqrjVE60mslhj+W/LH0uoZW1lKuJTJ5Z3P538g8A5RNdjkzLFczgPbMEYbr
+xWu7wiph6+NMAB6vkck/kwkl/kqnSNc7grJAkiqic4LznZ+s4keiiFfiTCJM4+a75kvFVI7bfET
y+QPgORAA5P77yo4sulUvjpkAXN70DWJeQND8E16VLn6IhU9rdiho/n2IfftVgB5LTvzI4k5WZbZ
qbigGKhSSSHSWeBl7ZKTe3xReutFU4J5fLIEP/VB3SJk6ehZ51JzwyvjGlbnKTNcYT3KI2yfPh1I
wlziRY4h+M4+/XQHZZeLZv8tdVbc8N5w7yXmKym6SMhXcgvo8p4mNPuZB6P63DxXZxHScAn/lp3u
PABk1li/ZezmTVuputBAc3moufKL4MrfsQeqPJypYWsuH7tOxAn55uJ7pLNOliwemS5Lb2yo5lfQ
AN0RApWr9imqfTOKQQL5zgY+gUsLMHEfHOYWivx3gWCaZ6mC70FzbC9lIZXIThypZ6ve2ww+/mX9
3CSwOMTDXrOHvCbNfTl1x1lH9CrakhDyez/kuycBax9E9/5ZeZBWf/xB9XQpmLbbVOfH0G7lqktw
6NLEeSGRIo+T+CJc6hhIXj1aC0zfRGxPvtHahq+x27s6cduFBuq1EQ68BimnNJz6vigKG45mZg18
hAAT9YL64PrG83t2IJPk+ESf7J/BLZ+PqSK7y0rRYC3VzZo3pRkHqeqowqPf6RYWENiP4Rg18AzZ
YNLJ7AqbsGO/4OuYa6yQSGreCOokxxsF65/079rgxMq/SFOXBhced9w8J45jr5FQC97zQFvV7Z6V
pwTdY7tqm/6HS5FOb0Io9JE6xLSjBXRkcgwh38QSaHqzdpdqCfYgdKoEg8xqFmyMR4X24bT/vfxf
nyp0MWfma5ygLV2MlvakYdiXYfLZ/fk6aLsLl8tHEBBtD7anL9WYF2LRavMaXy3eZWsFYTD0B/ic
GVQs25bma/9Tbb5JzwXoBMnMl/8dMPAAmY616hQvn9bE/sxDxwlEpwsG4bI6nGxPvHU7+zAJYXgD
D83A6Uef8RszzSQIhZC8ovqgAfM5e2XiODtrppBrhXA22YzgO20pqbyjIHlVQaAIUCKmzwq1iGOz
e+Tua0ezk/3+ozezrpl5DvEzC9PPegW1LI1S7nXs5yHAm+SRPWRS7qa/FLTO0/aav2pAoVBnwADJ
ve8yLiJoEDjjOljQn5r0k6cIujlLPjdlhcqfVy+TpYnzCe8qug1Hd1eJ6CtwwPiAwtRoFwsGiJab
6OgX5uLvzfhK/dxsO1B3hF76EMfzUhW0ZDKNlwKMzC1QZCuD7nC5n4BJDiTvWbq0Zi6MkH/RVMV+
iSlWaU7Q+V29+kmc2yNmQePBKON1+fOUq3gKWEx+u8lC+fChfwuE7jP10KeOAiMUR7qwkZNrjDsS
aQdcEsmAct3Pu6fmMdnYu9NPOTpEf486X8MXV05+bx0pZQrVj6F6mh3Rb2xrZ+/Fs4XsvfwH4pjI
GA/Wjy2GcTD/q2HqNSAl53FL7mCPKLlQBxo//Pj2BpVaMmTR0UTKSnNDAg7tCqHdEkn/SLMrOgcX
X4h2ojXvMQI15zXCKzRXqfF/oQ2brRjRxyfq7xkKMe3ifLfrYJ7VbOXpTmbBjtXoS9IuRM1hI0G9
DWsIEafDISjhriv9efK/LFUS5BuNVrF99/C4QftXxvoQd26wQIOwovQ2iV/2btEUl6d+VX95+VYJ
+m0uz3Jf2tAzuOCjRMz9zYMSSW+NEDqaX582c0hj/Y1FrsMww2vgoJAcdzCjABQHZnBrNojDnmGK
v7xY4K9l7lymglF6PU53ChomxSAk41iA64CMPU+YzMwRlGUI3YSjpnDokKn9kTQfqpG39WiHm8Ak
kdz8kBbJGWQNnh6hA2NKglVWFWoqUU+aB60erz+krTklgP45ltBffncdxYipIcBVCSfvzQfn3Sq2
PY8kcnlCwZipCBaZMK4UfFd+wylUnYy7+V0Icj3dLoaOcFv4Dgm7LqMPZfEsPIshBjt53E4U9HbI
0WglW36tG7OEe+mxSUrfrOCpXadKaGyB3Q3pupzqpr1h9ls8LV3CbH9GXgpGaAJADufYNRc+07Ti
TwfuDOzcONTEfs/Rp11CZ6fty/4wXja26tXORF74bD4RKz08fpj2ELC1XQ1hM1sUupWZLoB9uw+B
Jdx6OuwU3nkWnIoo9hMf/PRcbG71RGvxHPRmtF0n2jVYhcC0JM47xTFirW04DEKPhm6AcfI1YljW
peZqu3qryykTZW7R6ng5FI+xElo3e/uSxZp4/XUGaVKYh86Abl0KxnPsS2efKWJDrXPpm2DhyEVl
ZVUJwCZb/MJlRpVLla4cngUPq2Aio8M476U27rOT69UHGCOhORXX9miS1404L0CcpXylPTCSaKF1
DN2B2/YYlf1c6TJszpQmFiyFqfUbr2eDzEQAcNdG7//759tNwf625fooT0mfOMs3CvxbRLA3kq+0
dfuphM08EMj3tuce+vzmAfqZ6Zs6NEhynZYkgJhBKaTnqF5BrcXKUa/AoeQ1RhjHMse0VM0pzDfT
V6lKhXD25SDIdmTH2A56hsRL66kPFI+Uv4ONr9f/20xMr6dgb9wYd8awY5Ic7NB70fyZ2Y0Y8yfX
aEtbsVxVODSSSOm9NVUUamhxQmsuEnXovv81LNWKKLuxJ3P/0uzzEudFToJWs3RSJe/bhSwsVqIQ
VmsN1Dzu4L+rLD3em5Opwa8SYwr+t4gTHdEKtKOOQy684Tg8AAWCecjDuCGu9/HXWYMtFgbheI/+
YcBkkXbAA8LQpTMMLsKjfoil8RCYOTCDvREd8lUcMcEuLkclMyNmGrjirYybBGB+d25FmDU5AYso
II5Bl/kJHLjEqPg263kEItypZ755SMV1qx0qXw5T294T16WqNqTZUdZAhumMH3tTsddZpnQdq2gn
UNCz32SoQEiuAgvzaXUcjH7y8lUxD9M9Lpjma2tklbD7e3NDUYccmdsnvPrpKjD1+6ylsntWGt7V
B/X2xE1kzYRbTmWUgg/2uSiSZRN1LAVpjYEH8PJJ9Qxss3UHPIFsv9Pu8HsjwhwUbrSQRDJLKZZs
Ro143P4+zp7TgrP0KTDrEJ0VpKqg6O8k/jVc6If3rjVPjs/lhzonnk4VWVfV+5iN9pSgfnq776jl
a6B2vzEejX+B1tW/GAzi2ekmb1SrFtub3J0zDng9vg0fOtvey2coYHuazw6xkilxpObb/cggOKvr
EGdXVdK4GYU1iQnv4m+hR4cgYMLGCzbszwfSJabQvRh9IX+pIDSV5vejkgKP4P8eKcoTxTdfw07u
J7JSD0lJLSXvBxaXD0awX7KqU49KZROTDr4HVXy5ue+Cc24ltay+JH2O/iEcmnhdnrsWmHHJtTr8
9OHbNF7xxB8VodL4uFJXGb3jISXWfriHnsOf69tCMNeV3euVgYuqr6x1flottlCkTAhSrGi3BYNQ
9oKpiqSXBwu/+zjKRYaWIO7prh77JQ2/Gro9VRg7i01mag3PNsc705K4MDZMyXz6jln9kLT9eZz8
2BjYqCGVoKuuFDJmbKm/gEN8CFzJkIoKxYGVl2gM8ZLIHjTyi8aQTlHbE6wc+Fs6iO7Aru8awjDv
AFIUcr6JrXfxZz989D4SvUQF9d+LZZ9PUe47OQR9CkV9XxyyMCJOWlVNK0P/3UuXWux7+9rw8Tr7
+lgKJLX9MfPBjdD9ggvGDE+wlwDGHjksZE25aimccx0vA3ulMsCBi1ArHEHCGebB8MezEbPi2fy9
rI/72k1DwYr5XwfeWxVc2IoBHNf10EPvhmcG3fswNZ2+sV1ZSnPW/ICwoi+gdU6SBpNLkz/acrul
t9YFCmXY/uL95WInNWZwlhrJkDwvUpAvi7Jxke/3iueXe6FVM73hQR2NkyZ7z+5ehRGWn7S2i2NU
PF0ife4fZrkILF+sHzfim56PwUVvgwl914beB/AQKwcye8g4Dgc8gLgdVRXTtKy1nIGJvcVhqLjh
uOq14HeERHPhdxb9SAAaGcV3Y1pAvZPW0c/H9SDoRW0mB+zy6Jm6TvOZuvJcPo6HKIwaCf4S3xh5
j2h4ky/HHWq9jKC+pdk9zFHSprZfSG7BQ3t7FVNy6omFjhGHhqRtoO6ErjdaZZwvwlmuD0v4s7xq
oACFaq89crlYM9cUYky8FnxmoHFK9uYQK3IZBVTyqyzNmrESyAc989LfNctP3UnoVAdERdDyqpvF
iRDNnqSbShCMyrIWWmCew9kaQidOiwypptqv80sfN46Gmlrtexu6IqbDw0+uLe60saVtZ4AB5VfG
PI8s+EB0DgXv29tb6AUgjv+xvCFWLZki4VSOTGlpJDi6SpcUXQz5onI2i1jVfgy9Yw4oTzh5DGBB
v1A79I2MzIso7XZHVPhCxSs29uIxDCkn2TEWtpbaLkunYgiYQ58+xgZIlywnv3yKRvs8UM5PYFds
Wj+MfWaIzSA6mV1H3BeJGO6AwVefqW3+LPIX0D9V0Hs6E1xkWIAR9mgi/Kdy83zhyjpSGb2MKnJV
n48KtfGSYho/xTeJtMh68sSvOkVqB3r0LRD/x1nFXcQWJ56Y01EfpTdNfZ6SYcovx+TzHDDwOlWD
cJfLXx4mUONlkeQFZZAKZ3KPDbUC+pbSVpxsjWEkDBGWPcHrJEVuJPURoBkLVbm2Bu7k10Huz+x5
QqnNt/gwili0pSIgVYhbqi23fzYKVLAXxs3R61gAJ637bC5Q83leu90gui0Ia4gG5xjC+2jHHbsH
JS+BSdHXz16LczvCcYrU67wEBzEEfiM+5NPPdUvf3XDP2WqjlDqs2ONmGMDpHkWZRh9PdxbT5cX0
U7SRieIjKUtXZqy8fbySltQAHQhvNQpkAWixTcTMZa3QTRLhIr1M+MBSg1Lbnp3c2x3vls0EscU+
NZZ030aMATaCUs1xNbKgsRDfBWE1e1OAoy3wAqZIxoBdO488ZDpOSqSdUqZoS6+a2ylsFo4+DK7U
Cobtpirc1n0rg9cON4dc/87u8GyTVJpQeHRx38o0qYOPgEidTvOzJ5qIg6L8Q+3tPlxetHJbOcSi
z5YJ/nXRJe3dEXSwccFPEicu5UKkE7ABgFnONYuRR4oAYUruoyHUFW664+JUZrppaxlQrhNxzD3W
LWjPoVLAoy1JGZ1nuLf4ZERw4zA341C80YMH6i0IiLz7+sjwwpRWhBKaVRdgnOLvr96zKWtaHwHE
Jiubv6Hp+EY5QRPTySsTuivXl38PwJt5UVl46WeqJycd0FkxWPXy0xaSnUDlZai+SxCNYnDsli/g
885V1IK9mkndoZbNUSbt029ie+rvt3k2yrOyFwvyododmD+HlQ85Mc8h27AffYXaJBePzaVC2unB
DSoT4JToB88+2xwVJbxJ5B5/dxSdlGVGqyljFjjd46JwN9GztmVLX1AT3up/Hx4jZLc1cyuZDWyj
ZjAbCBCHzU6c1c0WVn2Iqc4iR+r0pCZjnI22Th1jbDc5wxLHjhgCdiJj2esxyPoM9/GaTeIr2B40
TFNcf5M0D/prbtb8OUCpfEfoqiIqxXLNmSnOqRd0TsFI34qjIcz1/HUuv8Zor2m8OAoPfTlYay6r
oQaqYxzPy+HacOEq2lHp0OkqCf+pUp9QXiWlb92Dmg4uUZsMYC+7kZA6Te7c7L+6OLcbxlhbAgV8
UkyCFOX8p94DyJkJd9WPydhaDIAjAty9+jEohVrZYs+IPF2DKBOAfnyhDIVNFB9C9tkM0FdNE/xv
rxM1htDxhv7ULHhjnrEb53YStIxIj9+imYD8V/RZ4X33g1xrtS8MGEugz/qH0h6RMsvBItc/Afmy
N+KW+O6Zy1UNTsgVveF9hVwwxcUnjhcIIH48LJaTOyPPpjaNmNM65n5pUMEmQGx0ncb7lnGJl6VI
AmBa47zTBKpGK2mTiJRTRiwqElrLokvgdl+9z9Xw8LgET9Te+cuFS3CgOfnDawuVse8WRcuk6nGc
Un3jJ0zTDYCW9QHlwcq1PQDG59cSBSbT1ONbRFfbQFx3O8jh+x1DX2+xWsyMA7mIbLv4LMRqrhcu
uJ/Fbbh19H9vhRvqEp1Mw6vQenhgRuBYg+uYE+KEgy40QmMrJ827Sq9BUhDnRDf3WAr2+qz//ZkH
G9rGVvkze9w6TjVpBKsEi6/xG6i/360CrmDkqu2JuSYIlcMO6/pd2rcOMBHC0wLbhHKaSz4WXdVB
RTIQGeCCNBEJckKqjHCLv0tNOEvP+DmxUXfoH/0ZR4OPk3a1XaDMgKMiILwV9S7Ww3xdKPXhHuDM
g4HNJtkbbGooIPQco9WVumxP/cXYiK56suZJcMpT6oiq0TTyARy7AI0tqGrimQEak5H/XNdr+/Wn
/vyQ4X+AawoqO/OfSYKTMbljgoR6WeD4/sRFdqbH68FIYCkTZUgLjxp1OzXxHDniQzNoLICJbuAc
SjRGDgfajt9WMXyw0vp9JJfeNNWsoLKG3jY5w0xVZO8stGcZ8ztw8yoIt+VXvwvj4LQAVrh+F/8e
W8XbFIKFQh7x7tuTGS/XiyJfN9VxwLDs5Ozks7m6m9FGuaYlkd3gg2AQ0giHUrNWDppN75xGQg7U
RkqrlC6N3DPCcCwaVRXF2OJaenFMNSTroMrFRd0rdra6OgnXgF1e2Jzq67QMxBeuHyMXbHHGeWi8
BopzX8I2MttYukSgaMhb5jtAT9di541tsMJJ7MNclbfr2FNhmKfiW+ndGSSEwPo8n3BRvY2SNWLZ
shPhqBz9Ku28SKCh4xNFoi38KChMqzR1oR7DRvUEVQw1H1Z4pSecp3VdaQrCCRFQKbPLp9Ej5kz3
rXR0WUK18AhuBGZgrRCSS4zhfoloGH9cza1vFOzy2k6F8Ej/dh0Hu4Mi7L5rEThlj9FJMXTUhmjQ
BV8PiSbGo0/hdX1iym/pDT1S9T2UlrQ1FMW3EtP0LTXFfkKDZrga1U4E02oizU3soQ7DpaltAf06
iZjWZRVFxuyraUivH1F9LOoe9hVeLVYQUJKdh1bT21TgIwHnAKMi901WNPbtNVO/UEUK1eTKQBip
g3GpDVxOztkF+3SmX4hX+XoQA0oWcG3kkvRVCEZYE9B47cu6iyYmaOe2nSyP+jVybZhZ2KELhLM3
cr6W80seLnOHfBDGiKBxFH1q5Vzi+csZdKmroNwao0Lcl59ci9W4gLu0aWe/r3mZ/Q1mF3/CZS12
ev+m7hlOJ9epOjHhpXbsUFhwBHK8UGFtoH9HuPn5osfKp8WDJ9BUIO2PdGR6fku9Xb3s8qo+sr34
+qboQVK2Kvj2j4nPggC+kwSCw43XZ0fkmR425t4kOOUB7RDGIek1J2or8cyoSN3QF7Yp+nQlWHKs
Cpw7vrc7Rt/SR7GCT0PpD10HIkxDXcfFc3Y+lIEFMHImnmUjpS2nmXrHgrsR8sYjc+xuwMxADcAj
tBJhdrAntTi1b+buvEkcPAPlvF48r2K/4D2wdha8fg4/D/EoOCTdEaTKtG5SnTqxaQkgvvmj89AK
X426j7PPbmDzZhjelL4m/v2UTulEjlXPfrwxsPL0+I/Caiy+IF8PsPmbhArQ9VTTLRc88VqXCYuV
1ATMwTU/fKkh+JMKFYNoyVbDoRH5gvW1f0r87oBXvvbSusrcK1f50nSr7Vjh5PEviUjBKyL3AEn3
5Zr5/Zp0OAKCdaZLAhZbJ9KtB2Dupall/J3hehfLUto0CjP7u9Q2HPMJivGQXdtS8nVpoBPIS2oC
eYB0CeOz0qA8NHluYAzinN8j+1vg98ibqL8QMSnnFYiFqAPxTIjgOJlPAtuKY+bCcJxOAbkdreqP
/XQyY/TQkcdR5ezVdbNw8/HB4xUsK7161CULLSNw3ueIpfe+36/BXI8iqNGUFqB8CJB1BSkbTVN5
4GRSAOfzHRfFBPJ4AeHYUe4MoZJs0+IkUIrELpMg1cP+cLb0IMhFpi17RLS3Pr909IxdDJ3VLm9/
7w/rsh58cFtFHSucRwDgCaZr197fzwMwXiAr78CL7utRIeNRw6YPslm8sOvIDF1+QoxZp7gZTNUj
RpsKVteKZI3gc6hNUzu+5YnLCVPFSyR4tbE+NHQqnw117yXlU7XisIy6pKPaZKNFyjxoxrdoNrf3
4WsBLliuc2/8jC0BfJn9SuyqK2Qb+Qx7jKhDUcMJ/38vbMNDLzx9HdeaZ65Yc1fVq2OXMYzjkPkL
sqCHrHf2ZbUM//oijU8GO3R1Infsc34h6RSoSA6LZOK97CD3HYsZVOOQPaqacKjWvwlDug3iyvNs
OYRvRaRmeQPjreLOn9yukBqYo9hlOifmYNSg8qgagqyMx8qxLBWuW6pjs5tDHNGLccN/a7mS3DMR
89Jm/dbnR1GaesBTDbm3tce49YE1ok/vqKa7ypnIeLLL6PtQX9shv+0RzP75B3LzOA/thoseNZTS
HjkZywrsckXZYJ6Pgp4lAKIlcNe+Tg/UH/6D7Pgo4kaMuomhYVSTins/0yaMdVDLvNr7JoYgwk+D
7zzq7TUUrzXCXudDTNcNoMggUNRXZyXKAyoPSVY4nDqwkKQynqgbQjHJTSKtr4i868Sl+mSiev9+
kB6/DqqXRz982X954Nh8Ck4Tx3dIDFjiK6e7GPpQt/ScKbcAnuM5J39lUorRJoWqmgSa39POTQzR
z65y6n7KwWrwfKi3NOM1RbscmuXgBEqPuInKiMrWyBR/3gYSkIzQqNjK6j24KOI2W7nr+Da9uvcI
qYit/QrGPBdxkMwoThMnOrpavj4nc7LPFQHSlF7Z8w4fSzHOsg1nmrG4ZGtpwOkuJ4blfngMDbQb
YxUISlQYeUqtF3Hiy/Sk7GzMm9v2Dym/TYc3lqlKsfwnSBsbqjt+obPAQLb5I0TpYycEcFnsw6eq
7dtOkfq9IQCGOgXCXFv4B1vnmWjU/0oU0rUnlBYa8BUebojyEeoZZQRy1Tz+/0VW0tFiYc2l/z0q
Uy4JvgkMnj1/x9Ech9qHNHfHUkHecggSY0/LplHxFoW28T371utsP3PDzsX3eiC0J6t8kjscxIkL
SkFDMeuXF3vwM02A9Ek6FYFc0bqYgza988fXPlLotEQgdFZAqzzWqTDSQrEOefboT5hliO7nFOEj
iRnDcQpnxcDibi7EM6A3x42aQevl6RKB2bQXSpNTuw5yfTRcpjePQpKiF3+n9CgiB/EWVYD8RonA
PrGZp9j7d6WOyB4imJPmh8nNAJHIvsHz7z5+kffNNjtJRqO2mpHZwe1Kp9EbXbOTQYeUFGurEu/R
CPnVw+9WKZOdaRxC+ufL/0FTX5btHaR5NZNIawdNiz0Hy3l8kCSxCfIdlSESw7ZdTJ/pZdAqiteU
uSCj+/Q9XNUOceLNMfHoZB5mn8CjGRiu40LWglrkz4frfMwk3gurEeTPpxQY82sJoVpvoB8PVyjL
E6eAiF5IjlRnOVHufoH7rx7x7bflGmeACYYH1rptIDQ3e2/6aCyC8bovr+RPfhTXMCL3nrSx1aEq
yozXs5cqaDdTwzzgoUglWXQT8nM7D6oTrBAAnrffqJYtCPSh5vJqdXu7xupw6rZAVE8A5j7iYX8O
lC7c+VzVt9ulVVgYXa6XNoi7nOyg8sQsRKaO684jB39JlbNP2Jkev410KTUScGHlpiLZdPvwSHQ8
BOxYs3Jnxdc9fX0uCTfhIrUl9mMTIYJBiV2HY09LehHfvAPQ2sl36S0I/R97jEx32fIMhi9IW3w/
MwoYw8tkgRlsbI0pebomaz8U9HI/Jk8PY5bjmR8h9NyZZ5vT8L486abC2KTki9uzJQiOGQHUamCP
7GuyU3z4oQEuLhis0kxcQJp8Sjn22QycqyKBjZQniXjWSwtHrfEZPuJrjeEdNoxLcZGzY07e9Inu
yK+g+OO3B7wkhDOhoyV3Vq01hSehQjxvO6iwahDmbAdmdofbeISkgocg1luh5xgcQr380HPIhCIO
mLzXejx/2zgywuOGfsEGJekz4i5pBuLUnkJC7oUYtFfDcsFs/ZQhSeFkzYgZISMgd5abG4g47jOs
MwL60aPPNrTNi+0xJ/PapyW2Vc/KUZtUWlSMytJQsHaVPKvoUMUdqlIOgHf56izd/mydORqo+l6+
a1jQaUsmgiG7vrEXzzsxtU3zxd7u7bJFbZCVNPqPqnNokP7iCDwkCTfTf/kxERSY284qF5DMe6TA
JWCji70U3R8hLrvsfb1u2iZpqVYyMLsuhIx2yu/SlQ3V9PJbHTdbr7mLJP+A7kNPpYNG04OxSFTt
WlKUA1N4nPAStI2pPzbXu+eukTlWtmpRdoegfprlxtZYSdlrl3O0I4k2am+4r9J6SBlbK/xO/oCl
6aBv2QmNJlbjiH7ElxBCA0UgeQ2OQZfY0qCknUIO73+eRO3MdBaWtMCcxONwhVAyae7tCD/quHrG
H54t7HChzveSYy/FhUY8qr8gVeZ7t6TC5xQyoDL5PN2vnDpH26v2mCIKmweorrwbVBVEElV3oyUq
Ti9EMESFdvH0cnxFSy8GqWaaC8tlGaSRzOa4qyOtuBQMBQE6y4vZZ2yeo4nc9I4WDt72Y6WdJhKK
0uusnQp/7J8rvbNNmGpdSyNSKD5GioVEF2QSAnMKEOHQI2Z8jRJaHyWgd8A4pC/bM58YW2RP4dy/
CUP8P6sW16CMXpli72KIrrJqufrdGe3oSUAH8RQ9lDELBleE4PcEvA/eYtzJCM/hofHpK7MK2xSj
7aN5tJ5l+WRjRtyozX4dTebzcWNvBJCcq50OaZd8ohLul4FSExDo90X8ctKmTS3iX168QT8IASBo
/HSpOg4MoAxiEKP5Y8cWeLwGiu4Uokw81MXds0AHqk+5MI0YB5oi/J8rHTpIlHIDScM84niysfW/
gZEH5KvMwEiRiM+E7W3Q/zpze9U2NrsbjMr1ik3/Vlec7EKtJb+TYd6C8aLO7H5ralwkTcYQCJwV
0sBw47CFmHsJ0MQCl1BiZ5hzZf4Lm+7WcK6H/wxqMJEDOlhP5b2QCmk39R6obznSdnxHSF/4TMJ2
QWplVbzdDPCeDGlgeoVyzHJgjGGzMUhsfTil2rMPImNfrBPqTOTIBrG+AMTZAy08OnyzjWn3ydqf
B1MEJogCaV8s8peJbyYGRQS70gP/nPH0Sf/WCTRhLqxxmYLQbJbPK29o0peuraBfybk51FaBU6PC
IhEzr07IZwdxayQONpzKhg+qk66saxKLQoB9KtgWXb3aADFw9kOGu/kLKeuX8c+ZrBu8tMEkyl7Z
GklRSSrlTHe1Ih+HrsTrBkvlbaZ/tidwUscU6E8+5sWPZ6V13palZzcuFoThCwjMhrf0ulifZBJs
C5j0Q5trQcVWTAYxcX/ntJAX7uTJBc0Kn5Si1PYdkOZRTJt71iLcGKds2HGuY43GPhgOnvSBhOG3
LbKod/y0U6Jv2G+Lck1GenUl7+ADsv/pfk8YQDh16oELxsVQLv9FOxZV7ASt36GJ8n0oGh9jAzaP
q4N4MMhjxDWAzqXJp9PRllHa8xL3vX8j71lOS/x4AgP2zDSk3p0aYvtuf7nX9CrjP2Di3Itx+87Y
ssOpQsPMQiqUFIypDBWVrc1OAAIkbrCQwgAjjU6wmPsoquPiBks1byW3PS1kVz4rBF/WAm1ggHyA
NBewykUhxopUn0FhyIzEnRiZd3sWslk/NHpqo+WviigBySZskKS9KhlsGmXtga9bg6V49tO/WV3S
UuSexiaUK+zpMVc06NwJyPX5VolGzJsMdqFRB9V7DFn+abarw6ENPEW+owqDexKlESWhbk3IrwoD
KXdpn1PznwKNhjnzY3hgu1FszcJzPNa3LL9XNQnu6wRYhGJBVzYy6fL7F8JCG4ztJDpeNMVHnPsz
fFR4x317PEir+B+aCpQY9F3E94IZKyt1Z3zTd24yAiCzixrUGRUaVVdZjRJI3RIgbW4as1/j6kjt
NjSD5RLVY28q0YkalAqEUUe3nrgs4waHMIRlm2f0ukULQZTRbUfzLiUnBcUp8Scnmfna0NzPefx4
sUXwfHBYARQ9/24egQ5lvtrUq/2IomeSBVbkUYhCsIgXEdczZRHAEEmdQYWrx1SlM3ZLqqSCRPw4
JZsmQ7RNlyVX166NOlJdesegKZJZBzC9PQNMW8fz+TrKM868WkBzrreT24dkHfxkNR6Z5W4NtmBm
ZOFMrNYpcRhhQBmDqS/j53zq0z2Tss6LnJrJQnnYVou8qL7KAE26aCVAjLvfeA3Akg1uS1Emvjx3
fxOxQUeXtRh2WgvKHODsSA6oHRsjY43ByxPkKr8ATe3CR4V1Ij5kuuJds7iei8i1+njtuiWQooHU
utcNLTG2tcuO+0Q5HekdDyUA6H+1cCWo5oxFbhsBZL7wAJJ6v3Fdm+DQMVIKWtHLIrGThnDp+A4r
UfIe4zHecnSW6xfPWuFuW6Bk8AA3JRERdvDEnze98wtIKcjN5Jqd64rNgXBsHFLMNebNh/8Wv2Ua
SXLChOi7959xjMHnoQL/rS1TVpqICy8vvXC+Jjs+earyiAiKUJiYK5QvoCT2L4J2oEQbecZvT7aV
/mYq/V1lL1BX1BgspN424YODvu9I7TJMbZluvptDzA3Q8Cbezv4Z/dwqSMWuFFbSUH3g7Z33uwyz
SkCAR4PsSghD2StainX/DJsiiohF2GDRZkjnLVJdkq2WMjE2tgOPwtPhGEognCkam3LuVfDnIQTo
vhfkCAT2srXlnhQ0RCIDOuP9NkuCiZoVdkSJR//F7jHAlW1sojbc470wYh4m+MibTKjxSXgdnfL7
DGkZ4ylgCe7/Dp9fSlFMvu1xsMJM6v8bY5Ps+rIkS5v0z/zjtbHlUopxpNkhowKhJ0LvJ9odcn5H
MGftrliK4DdAtHasoAGMtK/int29rHH2iNFcAaxFnEelMzMxRYiS5mJLL8oS27czW4r3KlT3LO1e
ssWkMNyXrJa0Sgch0KyxDOLfUcE1MkEJ+iylCV/Se6lNzBjdgmXamKGmgFbK3W5InXKRle2bwN2N
i3V6ziqSPW1EdA8mxWYFKHQpBJOeVq/03c8OPwm6TQH4O3+fRfrNpYDVl8ClCFOuK/vhDNtuoS/7
JPvaeRvqxeU+aOHpKZV05dLFZimW1bk7Yia5UNkUcNhLvDveXky2odff+FKag+v+exuk3OYbod2x
0x6kGlfA2qBCMfajlOK2GUOi7nSZy5LZHNZD2TISoGgGP32SI1KROUW8BeeR+c9s7eNqMDozKKjo
yLUxTqar6aNTOLDe7rGcVbXcxeOvxOBDn/L3qQsFx1HcaApIkE4HhpKToHsdw2pAaWblZfKrgyT3
Ak9FRFnXMKiGBIlUoMfn3KVJEDBmQRS6TwqSrMqQxT9cx4jJm2tu5yVvxBE+3gKaj4jkJV+pMAj1
EuRdgL2QzEG5l+ACk+iUezBv/nvlfoyZtK1DZQWzPnIXn4C1x2yu4hSAMdkYMty7l9HkLhk0vJnX
K3jBd9JFuj4VV88wEALKbwEfT/JRd9As5ZnQqemW792a4/B566Gx7ShTM9XtrPEapLA0kNoLuHjO
xtjLAl9xdnCGPtgkdbsygjt6j+Siwg52pO8p8oU5GxlM6JUr4YTrq3tn2Dw49Pd42xdfMsF4ofB3
gxX1Epj4OfEJiRZ52nnhESXiLutkaMWccmLcVrFumAkDXG3GWLVKFdJVJC2cByjeiYkcD+M9GW7r
FoTEyMPGhAWdVtcrUb0NDQaVqDWcL5HvXFPHl0CccRr9/Y2COMmv61LfkHBat0xNmoMmCpJ/qfdB
uSMT1XlfloVygyLsQ5Lq/n0GGwBM2zGRRN24cFi9fR7z4w5PnUKi2f1svxSxNKd266KeUWuKAw4E
SBkmS7U+phMorLqsdOnuNW+xDIc07FDv0W022MIO9R55JaR/B2B3UHwbekGd48mdToQw8yOlqqsr
MqT9hdFNV5Vg53bve8mra/4/a19+6To/yoY3EGRfHSgCcBUHKMIZbb4FI5oKJu4+uRfMTfbI3LJb
Wab5Yn1XadLMD/k7NqKYmc+qN+HSIGloFG1MTcfWuPpRlBiNV7xusDHtOHRMUKxwR1bL0QU4DVd8
tHhaRTeN/uC27cNkHKef8s7r/2BsupgeO3sTRkYciGe9mEPQ8bkHw/+sB+J7XC/MukDf/h1KP8AQ
aLGUSh3ZUdlVzufk6NlKfi7bOSzSLT6ZxeXO+o0yVk5d8dYR8VNCFZg2+KMDVUQRwZkDGNOBfzGO
SWts5P+Fmjd+ZObVzdTrS5eOMMqU4mk/2ethLfxBkdCKs27020XMA2jJzXJKbOUiizKf0ofIthnZ
kJZXRSx1uivTi9pi++BvAvAaW2brduR+0uJjqpLKyJv7dbxZ+G+bZOX7Jdq05v4nQOoYHoPwwx0d
5zaBrVCuDgXzemfB1BS/L6V7owrSUVvSzgi2C6Kva7outAccUOe4KCtL00PN5obyKkb9VYggN2yx
Qfm50vSGfA4LTDu9qR93+cF4awYX3s7V8NVdg9rA3M/ugMd3bSi+07rCOsEgfwfIqYkA1xpb0CGo
7sXrTlFUcOC68vbPpf+faISid2DxhJghtzZy1UZvnnQnoUfsAMc7VUgeTQEPpAPkqn53T7RNNgT0
QCGyqed2KUdyaH+OuLIYGkGDMYP1RpLk4asU/6z1Fm3Es+JecZdevvY0xEt2uxSEkY42DfTdvTYA
A73dbdGVyqKnDypX4AKRDuW++oeCQtM9VLJIPfLD4klNPWL9LAtUsm2M2nS7uRAvC3LuQmiFvvo2
U7TAWBXvSyzmuIOXtGVButA1ebpddmQXRGCLh2Jbg+YTjGIedDCIQtLpSoXHTDPpMfIiZYtIfWZt
9lvWValJ5MyN5y3scdYlvwFUsoxGlCKhoNFcsasDuNmT5pdC7WEuS3Kik/ijgQazJF8DA952d5kN
iY4Kbynr0WxWGEfyObHuMo5HjKYjWO9gdkbjj5WkjSDPu0SgODAki8wWvMJeh1PdL+kM4MCQvjB+
jpR09FJ4d2O38ytYNRPq5xcFsj38ecbSTszCl2Uj97SJOG2wTb4RcEUQM9kvANUFzJydsmFXEtwD
FuHV/DSk980Sj7rabEeplt559zvGnf+S3PFGxGx4Uap8RYSDlt/nY7RX0Quu93TV6ql3+KKNhqOt
MRCtcvU59KeduhIDJ8r73JctUixSiqhsIfBeeGn94Ok0kDJMvd1A9+5VBb8GEpVDkFdKdNj69ylR
NWIWYrmoFyTfOXe0MR6+JUOzs1BPTf73q1jGOfOVjz3CqjNouPHEL0CfLySS9+zmc4LT1xVcBiZc
O+hY2LOFTwHSAhJcmoFgZ58UAyUnJU30cWCzjQroNmqPKlfRw0svhq1B0fVTE4H09v+sfZnVEGZ+
QiRtqyFQX5RKRbFgjwlkH2PJT5OhrDSVrocz38OS7SEVJsbgOGEujGfjmaKrKo0oV6uwjmM5pzwr
PZmMtFnxYlV4KIe/rKmU5MVf7Ge7tZRL/5lgT7Lng2eSRmMbPpa7JasMqzwalvnLXjO4Bmzm9mgH
LCTHf64OxlttQAaFLqPvIx5W6GYjjMkw75grWp4lUWCywHBTe2k6/J/bSIA7Yno3wA0oIuv8fruN
oRfZFiSkhQD5NMRFkkiz2Y2n20WkiEF0y48+JsHry5x4sbJdcBikEezVsJRhg0Vg0KdZTpB2NVs3
ELpdSVkQa73MBex6bm2VJIG+zxJ6awbTHMCRxpHr220b4NlRC1ET3dUrZ6HSCtqY/eSzg8m4YazA
YW63lZpuJf5tdS/ZETBRnOV9wgMC5c5kmXpl/0yOPzIduYO8ZOv4rYY9cPeyYb0e3/UL4vWNkgHU
quUTuAv6LsnkAtP0aTeV5ggRe34dYOM4h6hpXrosfIypM8qnqZkkjWxn2cLdyOloLWdXlU5Z5npk
KDOMUDr7zYeAM+d2NLAgNZrq/ILr6klax8FSwRvUmnB/PiX8gAvmRqoQ7lK673HUL/ZLI2n9r0pI
6Jc4TCEoO+WenQOKJV3/4ncTWn4DGViyWaOAjsGMXQTbszfxDjrcskGuphm9p0U5iRQ1/b68oVOR
MSwWqe0sukwQuHodlXwzWPe+c0n/lvHOfWal1HLo84llibYOxk34JIWfoByyelSGDxoXZ9xeT7Ya
gAzMQitgeQV1r4u0tsCWNNL2RCfpqal/k/3rjLgav8HPdW/f5MF+qIOZUoXl/sT5fFrVwzjbhSry
kEWWaBYHaUErC/qqlqItTKTJRGLHOGNrN1vpkl0vWXNGtjYxZxhSyrpg4Q1OoK+xryZvIRf978dZ
r0ijgAn2swKWQzOpttSxFsnpODhoa70KQNRFWqBuwzcBPXD8zKX+Zp0dlCBWfUfRs8LH6NLL0anX
ip8i828KLr2sKPxyVs75Rn8nsXlQMPA9qRKO8iq74jJ/VKo5kdkjTVwf/h0SjQbdiDghJ55SW+BO
2wwiQgEZ3NbAOXVC+RPBAFGg6EjtKnGqEDWleOIWu8vSmeInHzxhPw5/8yxc6SXnEGzp5dpgOGdL
TrR58O2MT6XsH1CNdrvsvY5WP2Fct7HiCMNkjBNyfT3U+6y/F6/80wieJqKMSWIDR4Oma81HPPhO
Vsc5upDiAI8hWg9T1vtYCqw4fX4niXPO8hi8KMl1kqPacXbWzCyz6hYdhRRi40CDC9xhZH6OmsY+
Kgmx7W54wNLH5Rcqvx6zD1tSfoll9/RDShRMgG4X0czYDGoRON5Kz9dm939dcjs2BC5KYqlAVhMh
BDOOlQr9xeL54E9EMoa4fshDVj1x0hERy4KESKoLbyOLSSI/Vh6/MqSHogqzFuBiqVuahBx+xyb+
62sZYIBVsroCodhXfwUir5S4GMaWqhLXYJqpRsafXFGBzVcvKeMY8Rn6cV/EhiGR7wvRwhhRBjU7
Wh3llbaJBaXmUDzcXY2pMX1j29YJNWgbiNesQF8EQk7m4AztpcLFQcKLobvG793JpC1iSiH1GqdV
rbRZy4gHnbSl3lJGqCd5qxGFo0SNgHzMUYdJYeVUuIRDNPfHfsHtCPqy9Jpo62Chhn54iwxvfbDE
+mop0Mm3o9KiOBWFY9WWO0/B5MIU5X748Y1o6Hz36eUqwFELwUq0Uk/g7ow3ZRYUUHXl26o+WA3p
+fOYNIiC6wT/qzCaM5dpmdOQcJ/ioiC26bYmzEHxbVGF9/tHhk446GX9NVSWPrrV9dI/IGPEkhDN
bSA0jQg1he9AiC2ysl8T4JtaJXk1Svq9ay5lgvUqKnuaw7JS/XiEsD8cK0RsDxd9+m+3FDrvL3vM
2oqTqlP7h5bRwLfAtrOBrMDwz2L1v4yN5Mf7y1KFLZPCZUfx1upiS5RpvAyTVU5iQmsBDrpgbkDX
TD+EpMi+I2bGxvDREDxyBmIqfTEyhLmY7AmXCYG78F4N2HqQwOLd0Uyf4aHSHBdsIVH5HzYInX+1
cRvCvuFuqmxMUR28fu/5WlEaGr5yFPwXqH75NI4EvwaMdirfY6N5oTOR4ojgmSyEhpsUtAT5Gy20
fNk3p7y2+NTFd6QEbmfAgBNdlP6lnitiprz4NUsPSHjlzVgBxu3vXKt6dPOn0ZVlbQfl5a8v8Ch5
85VXFJtkxe+wZJb1G00Ges6XPbYWUd3kF18HMJv90l3mpFrvNZ7bjNaAOuhCmtcHkZXwPjfEeyJ6
JFANQU6iG4rUJy4X9O1InY/eimICMyCOmkWM6o+wxBwEAqcL17f7ii830uYoGGPn0Zq6zoc7xrLz
1Zi/HVrsuE6dq6ioqgi2m28xOXLgKYMpdjfCqMXoffcxnhnUUIS3UQRSbDypQIptF3KRtPJeQv4O
RZcLH5dveXBe1ed6ncHa4Ia0HkgUoY0Pv2UQZUHpatzoeOlDI0QGXugrpSdot2uVIElmXBWHXPx/
ZackXmN8BNgLob4uiDly/0C73fw498tdSlxFQhEQ0642y+CnXVkc+kpGnIaigOEmzrqKpANjfqmo
dYRs8wma6N4kbKukAH3h64CCh7MEv6vD9mNaYYg8OAr1b6WHJnVgAfEU3bXyblXv0Qp7vxtaHvlV
j5G/JNvD6ULCqychVVe0Isc/spf/l8eWThFLCxIOsj7BUBQmdDKZSBiyy1fjZ0zg9MgeTcYbAIlo
C78fEoxP7xYc7vyomTb3jngIukR80UZ11sJqmxqSJ3mLsTcTYANbJgbyLcbQBODUHGTp6sAltTm0
A8iPAyZJ4+RWmLH1u/IHzrA/R+6LHALtyn0d35xQl3aHHEilv3Hx77enLfb67ZZcrebHRQ6gyD4E
JG/eR/xqQu8ayqJJn63b5QrklTBOqCDi8W83iMCzhJSR3hYJU3CXW9IeSbyZ4VvuFdegfdHg0eu7
JI1tsVMHhCOEaiJAPb8HHU6CptrZuul9RkS1yNfA6mh0UiJZWLDqjtNZZbtExyKWX9BlgZbFDU9W
NxmKIuLl0KCS3aaWXOGRB5ZaKB00dTEuXRTmvv1URkvDE6hEqIcF4akTK7FlOQkctl26qXgJJMil
UQGdzJonfEJHlnYTxKzgEv19ScdVKmEeJ0/qY4hrEEwsyEHkJscoMpScgvWYxLygdleteBLu/Fj8
jlZ5+MrpNEiaiWPMfhY3rRn2AE5PSlV3CjWVmP8UqhfY1tXQEb6VYVk73PFHC+Jcs2teqjHNh08j
ljY+3VYIOnd3L3ShIGKGksV96L5GQQy6ywxTlSCInMVDpkRv1K8eusmJ9DIF3TpYpm2DHnFBBhSq
QInT9IXhoJl2HbxPcZ9YI6dRUQeLrFe0XbrXntKfq0b3I0f3aMEr7rScLQUHjM4X3AWMUBE2R9/L
ReJiiskf9qLizVjoqObnyxxjGjwbv8EgabDpQ9t3ReoN4tHpJ19MKWaPtlY3WKXP7PH417x7Msji
slDMjtF/5gXbimGk48KMdCt8od9tt12KbSeQL4zKlFwIMNgCB1IXv/BEWqrjc+KRxlyguQgRVp9N
Mpl+9C3ZtxRn5iCO+N8mkQ0FuXd4eZnv/sGfqRqA2ifkUVqHwoeFg+xPWdxKoE4P38kYMPt/8YqG
0DOqFbYb9iyJmVlgzPfbRPpn1gLbPU41+8aMyWVjWRBKJNptO4A97bf95mwr1QXzjCAdqcgpFTHn
6DNLyczG9L6yoVYejJkIurJzAeuRLB42A2eCKjGnRDETnpRuyvuhFt+g/zdSvx+cv3xLIwikwiBf
+gpOrA76+zhqByfHL7eH6f0tZQTJ+fQwAWPhXhrMCo23UUYwMwAUkcnS98/hJZ1qJ4yBH3lsCPYq
AHpYQ6xzybNv9cyGO7GBUx8tCQvQYJrJVXBleMVwvvazsq+IT9rB9lB0jp4gI9xWpDgDabuOWRFP
iqpe/jBjP93nyJjqvr+MVaF72i5Q1/JTdWIxu052wl0Ll7PjiE+/Lb1QodbfFJ3RvdZIwBXDpFmQ
gCcH/XYdcYX5n5BM/+qDvjn4AGSmk/9WicETCpPaYfh7bzmeYAxN8Xb0lIM/HEkp4iOdLD51l9a0
787kD0/9odUlxO2K5i2zKyqV97TSYRwrbrTGR45d2OmVqhJ1Eq6sqI6CBtHj2Iy8h/yirIGDwVSC
cDcqp2szDFQuk/TSST5cbfsc/PAWnN1+gwUOUUmutk6as5+N/lFZE4GgrcN74VrYTCVhR8HeR55Q
hLqIfN7eROEpXfmGy0G/RD3SglfDSk/CqZoFaOj1QoD0GXSgfWNMxNj4e9EExZ4MEZBAuri+3HK0
Tc4MyrWu5Cz4jlG+N1/5h6+UXy12d4W1Ci60kJrSoqDKYALEQ8BicTtsTD2tgE5qsAW0uOq5dor/
InzEuu8mBtn8nCiG5zi8iDs17dlPZj7OpxSvE02O+Ub7jA/nywc8TJuHz+0kZlShQyieNPgncm9h
Vw9dYf02ml1Qqk2/8YpnM1bB+0kdSfIV/8NX83NCEpkbVbVJ13n3qX3BBYwg5xr7ig7nQba9cbs6
Uy5BK0hnOehbd9ZYNvdMXOkXZY44JLfYIkCGZOHvznQ+FcIoHq+UT9hqEvh+dndzPVxhGIs2fJ45
l3QNdQe5TZB63hmT/IKuUngVSBC0TPdmu88773jN5ycP1gvK2p0AP9UE7p61vJu+ZezDoLROb/Mw
EMGYKinzrMyLPHngnGpE1lH1vkH+Hh/cl4kOalXvQNCIFaDaxJ6Yb0EpGddIDUwqpXaUJbSsa1tw
a0nDi0KuzTgYzlDgwWf0o7NsWs4f49fBPBgtKoEV/0AqNtoOLcUPDIirKoDbHeqmYGkymkirstfk
k13c6PDrGz0MU7CfzSpmZhfOgDAMLQkatDO/wU8kf5/XtkqQfk+DxGEQH0KdSJjkqYDo3fRxCXJx
OPM9Sho0aD02+x1VC6ybhnkhKOuJ1fVdB7RdV4gZ3MqlcCjgozJqNJtEPiomc4mxRqLKjS+PFSMS
R1GfRTlrC41s9H7XHo7dFBWqfqToJu1AMpLZpduLhy383IcDZ9M7WwTlUG1gz1RnTYDq/n8kMJE/
62KPxZ2FbRV6ZngcMk4egfg4f00uj9QCsShRL7eo9UZ/sWRZFaBkeLEyNINBGfTIEtKq/v7ds2TZ
1MZJjsHRJA4+aUWmLEfC2tBbyNFgUWlTTThV6WmITbx0ddeeNLeQXr9b8MGNt3gCMXrpzChHonyK
gTWCQVqQ4SZ41zjNNEi/LwNvKCfkYr3mHXWuqfKYhVJAlFy9R98zHkQ5AtXirS16V21dY6z9SKrR
ut85UUqhtn+Iytg1rif5mExgt3GJZzBcm7X1qG6nThbbC+rQOLr0rBDDPylDZG7NeSxIH09/v/HQ
MIGnrGEj2wib1pYFBHn5z1B6Ph7KFJwsTqzhQbjAYXDKEyayGhH/c8JBx5DfuP5vg/Obh2ymGrIm
FhwaEn90aOn5Hos3MyMoKf9n93DeTal/oB1jwuoDTJ4iY9QswONldyEZn5iEcnEdJvLhx2Ih3FOP
qA49AEcaDkGiFFRzCCLJbq+IGMVR0UF/zLzTFsiUzeOaKbzTSxw0MeIf7Du0pN4S0xWHWXALBSpx
yJsaKz6pEdl9dgmsN23ZRZRbcjKycgx6qZkbSPYD5xj7DHDfs44L+IfwjjFQVhqK8mw9ycuqVMUs
zQX/7wghpGfHMmmXuqv/bPz6UNRx3+e/8rMBj8HR+Sd545dlQoSPIu4/8w4OI5fKrdVr/9S2r452
LRJ7v5pLnM8hhaJwtuVsU6E/83BPOtSBKvP1raZcw7GrMNg37g4rnYQCMVNEOPIwWgU3t6eWEOQo
6o02k91m8bKNGw98Q5nWNQPeyDrzEo6Q+bPf/nkEmgg5QuDX5A3Aj4oXEXx2LuFlygzpgHdVhqIH
/JyNOW3h2fTWD7YpbtJQ5YRvjHRjsm9vl9iwiSpWD2Ihg4o/GP3aQJU6TxoGCOOrNzfeIzo7vVes
LCYn/54od8OXb/5s7aR3xBIHLxS5jdjUI+gMJJhskLOi+f7uyjrlsbnujP7Uzi7/cUDZUoMOPo9K
ylt9r45nVVvT+ZhNxNqSRZK/KLx8P86jgVNBJLwJ6JAlWkNXUgCO7uK/9XPfOYvILHDGTiQjlfZI
XgB1iC0QvdIsmnr8GNUh8+WLOwCSK3um+8qnvHJCN7l1rmuPzhEzcv3W9MwIJPFHWeGFUr7gJc+X
f37Xm6XP7Gzpuf82Ca+4mm8ZXHPDD/nXpjwogjQTlC20G1SRxjP1RHy4/EDmubbjec/n9OQjVeBB
+iQqlIuFj40JgZClsH2CZ44EuyxEWIDafkSH2rbnj0YJqE6zIRNtgOnxkb/3BdXQnGb4mOj0jJAe
ZGd0dznmvo6joyQ/hy0qhWj4UBN8COV7a//qdzcQRPmCSMFUWokmWhtqFZyFicuG1PEQ85F3n7P3
ZLiMD9xsbMKmAFyGTK3ZaYsbCHmSE6iRlNLt3c7hDhu8b6iWT4T8q8NWbYxcuZcPf32HTUncje5A
qmP3464HmxNK6Pjm0I9SrTexeSt9ZmWjtid5cP+OljKoBvRDZ+pk+cHy4TqbcKApM1PV+Ilui2CF
UEOpWhb1dSjr5PCYNaXboiAsJmEi7/JWOct5fEENFsvEnRPmtaQqdPui6BUKNrr9SCgJxdNYoHMd
ZpdjVDH6XYOfsi/bvv4FLhq5mbcp4dCdYmZpsPPVeoZx0Yl0o+BQ72m6yXPgrx8qoLrmo16lSNJN
/fMCeJLUmHrzXYdF6lbvUSVOSX65Qm0TNgkoPJ3P5tdVRQidw+v4xsrn+iZ1+pn7tV2nuiwbIbUG
hvXgQdU0qygWhJ6DYPJqsHfn6d7CTS+V0oz5/lKY4zUqA379VlUAMorLnOmSUnV6CPY4dbCmvC72
lm1LbB/PyIPp0i4zMF+ycHSD9Gh2Tt5Lermns+StHF509DdMI8En8NwglYujmPTdwraTqxOg7q/S
uzgY/hZUSgYlOeigCfmOExtfd86Lj3SBTu1mAMDsVdyMuaR+b+oobcm8wDFzq5ir1tCkB7Bufukh
R34bEehq9ESVAeFrdl3WyGFKMFAlFHP5MOBiE/Dm88qxslQHwGzgWyQC1MeKSetEMMlEpGPEpzeg
llyeArz6obrpQIzpqAR0m06fO1THbILsPiWnCgqXH1+rPRbOwuP2Ln1CFg2Tc45PQHjugwxYlxR2
o5wHHGDI6qP1sa3bNaJ+5ydUiTe5Kpkb6xDjAV1+KWkFN4htv0T3s3pb92ERuVa7O+Hh/Sb1R97v
DLhBIagioDcRysd9glTaC6IXRKejanIH6u3N7UiMExJquJjprWwlsBaXT5R009PJvsTCPAUWMx/k
hLQv2Xtk7eQJH1ZYTZYFBPSavD2/fduZLEAslCUAcR3pxWOp35IqQAbqOmUna3XMsbxOldXzz6fh
xfXT/WhXESTOxWRUOYln3/TiZyi9t4jVVP9w4MYdKluPo0zyRAW1FVPMowtpY1It1waxUm/hf5fO
ZeOtZWvulwTgvDogB4SLy0ucYyaHHDtM3TNzFFO6nu5ebQ77I+QguNAWh+y/6Y5aWODD+BEaHgWu
VJYfMFHzRw8fsuUqqRL/CvW69qHEt+Pu4M35T4uo4V2Nw1pGiB4pRJhJa0aBi1t0n234RJmW+GKp
lZvUfbmySWzAoWiCwQWANVQb8jfbcly51yboaofQRA6ViaqPZxf+DjESskYMwK642T48Rq6STA3y
zNXrx8pB+1g0mYDXXE+cpFmULQ4PyTYxKIAdeGDgP9W29DBZJCrGJ2OzjOrQ40wR10Z/3nJW6QVm
Y04VZS2TyeskyJoOFicdr77QKEqPH+0E+auoflp4cKJNQ6ffuiOFuDfAL7MRQms32b8yI5hr0XqP
2yEAiglbC2HhxAGmzFNQLkcZm0JdqLOhnU4axVqNnJELBOZUVynjqWFl6V7t4Lx2uuZlI4zOPxyK
OddiFCNe+nT+X68cG3aJA3hcS4DafaUg7GSTVw35JCCK8ONMzDRpPv79NCezZZ+sm0CuNVNKFS1w
J+I7Gp/+TlZsHniP6fpOTysSAVBpDGlk9FVUu1uFnmayRWAFChdn1TTkCrBadrOcHuV6Bv13DGgh
w7d7x2ICtp9rsrRv258jnq8/doJlEpRU3g3ouV1PQFhl6SQDHro8a3e10LTuko9/nQLEElbKAlYC
Zb3MVzjXg9AgT6DOSiTw25lSTGQMERtqcjpU+JWtVsEYSVtwF8WocJ6buBtyvuxMsOPX0LcNAucB
RjeviZGGqm+JzWGeLfrJyrzImv23g5OVZBeilR6Qke71hBfXc8Mt07twuQmftDVZK/Tg6ECYFsDd
8AhLaxTkPvMEsz97E+vGg/q53qhcITJRP/Xu2akC/Rs/RcxOS6ke09WK6igfGJuy2iPy5WLgvdNf
FviXXhnMjgHb66A2BY6m+0koa8EW2jn2htqLZRVI5+raCAm2un2Cr+qGlUxVdjr4jjeadPBa4UuQ
m9jrteCJdwGPey/LXrlJ81IfbeMPDkYv1d7BCBhiNNP0l0tp+ZbWttbYcb5gbNcRCJOMUHv67+PD
Gidg4BgzKZGyJPmHVi/MK9uv/G5lcccMFddxA2vHG8OZq3+lS1nj1ZrEtJqdTOE+wEXuKTUl0d6m
45bkC4Ch9csZhCsY87izXIEqIe0e/Wwu5p/MaG0LVhfaiTzR03+1xgLNQ/ZI4ZiMb0inEagLan5j
frjX4T5oDfmQc28aGguLQv3sZznnXlDzBqLlBV4p6uw0N7+jXui4Vq+PUdt2a4Q3BlrGFhb9i0Qf
ego+zVL85lbjNZlHvgkcXJ4O1sDGRHNdHaQro5HRaNhkPwCWTDeL+iE+kwZgkvOBdxJaoRoAaLTl
+zSr2BFCDuuLQVItjYZGpNrv0vL0x0iwC8AqDLdyohNgjXe+ML8LP8wgUibU1vB0djF7e1zDVa4H
FGZL885h5Dtr+xKbeM/eYEJ5GAy9q7GQIHoDHtxVy8W9DKwceZy6i7w3IqaRbNKiAiqvCmvr2nzX
DKgPbAi7mDyrLY6CSZr7ROZDh+QnzostjGRuJhPHTjLElTOoYpfDjNob7eI2fwacpEwdXZcNjxgC
Uwt2aOCH1Ffhg1pgU9ad+IKfZER80w4RLgitM4ta/+fp/EAW4KEmeR030s+4B0nc6cCNu8keupur
sNj7V5TvMcj3Ypc0a27zrJ4vzjq5t7EgOuHwus+wXnRqEvx/cEtC5GYRQUMc8JTTm/1J9IUkMydF
NoUIW8++6ZYSpybGs5l5QRpf1MtXB8OJM6Z8nlARySRiXt9x/cB7Xp5m+Z2ct74ZH8Rb+i6bQ6Cf
OiVimr/J1VC8IBbvksqP9mN3s59UOIbGO9R2VAqtfNC240+LBF1TFnLbbdXFeQz3N8n9iVh6KgpX
GmJWGobddae9n0av4d0UBjqAyFB9BGO+azTuDM6jGOLlNl0lh4/b8j8VgQ6ucu5kzpfAkYUOepyI
sHwWDrnDbWa2+bGnKAnSEYYozO3OBVpZ/mS8qlI4EW1VM/t6UjGgJMSRODakfVZl9Jw55HRCvHXY
kEMZPh8i72Xnhuk5mVpX9jkyvNey4jtXGd01lcKDoDxvCMrJsJmGXmScqCL69mfFfkt6x+dUPsVO
7NazlLFI0qXWXayFCluoFMQRFakJ/IrQ+KPfDqksUGsFyS1OiTjJVWDdmKrKm4aPZ4h2tWFbtV13
QSIxRMLXn9VQmE4fIIOQYW2VmzbLmaHdITjMJcXXTmveB6jlCa5ltJmf5ngQ70deCnC2/Hv3RgAU
vvo7Xe2NwSmetipYAvADLiFxGYqnPzy3ZId9RnOpl4HK7LRM77vEkeV+bPm0iSeZB3QhBJyTCDCw
TA9IebT17EB1qdjkUuVwMQr5XaZFZiokQ3JuECfUuzVAJ/VxL9R9RXzuHw7UQoEDQZou4gkAXbEw
a8rhzSLTV3CgtSFEmibQNYXfOUTeSYOuuPrcXeybIAmwp+/183sW8gcUOFRZFlyMxSXlFgMhI23W
xixiOLXN/qvVJ2KtzRJOmxi3nGaqiUe8Ffbx9AfZEdZyd0wN/nojN5b8reZGuPIAwuJdx2+kpKM/
OBSjpbhBEcZcNtVWN8PKX9VicnecyqqyWil1SnVGmB2KkSQp4RlWabHpU8cfhSFedGPnYaQJ3g+2
6B3zeTjirSyKUAGsU8rFDrn4HaEtpnXUGbnMhFA/qR80Zb9lu7UVIbd2gDyKY7EitUMKUKLf8Oyx
bv4QmCpWD9UB8KxUqmzO5nVznxxUtU8/C98CIplbQZOaqvoRqoD8/XOZKLoSOdfNFJ3NppQDTSJj
oGvf1TcCFUjrXjgW3wRhbGfNWfr6Mdof3bjts6knQe34k49WG3buKHLnnH92n5+cwie7XRnb96ym
7RoBkBkYFnpoCb16wWotTJG3aN/u3uFfP7p7//UhMBVCDnXR+ywfL7rQUodRovfLOnQOex//Peew
IZciZ/vGUktMMK6BcGiQB1CcRFCHr5Zjg3iZ0if6bIBZqrSZCWjSU+u9SBQNCfAwdbqrHXuizdrP
lgiRAsK5bUVABr3kkFFZEhTdX7DbCO3JgVEu3xhKj28LJQaZN88LtQduffYCUOjDhtxC/aeATzzH
fHwS6RFXHrh1h7ld+mZrwUm4lJmcTw0KjNvVqdikXEAXu/S+t7LnWUCrzdNW7c33GrDdwk7vVYgo
xtSGN90tK8DbJvNewK8NwAFbp4tMq3BaqQdS0U4/iIemAZFbfseiE5zSGqeIJ/aVmGeDNYjGAIX0
kRXYxSE6b2+CK8YOS33fyLEVPAZ9KzOxpCDreG1E1167XPvSCATgLYWqkEmMpA9wB0IO0JZy+beG
ZPP8J3ZiT7z+N/jgLxF9HBXNFHldDPa3oylQ1ZpQlq2CccCQtgsXqVupEATN9+Qrfm8UelegDxbw
QlZsOBk7lycdL0Aa6QF2nxGByjKckrgpXr1N/VR+UpP5TeaODXIYGwlOAEGPGEM5ZMO9XA1PhOHB
UPVP6VskZoxzQl8DuLHsEKahK63Cc4ITF9gG73Oq8wQl25B0pT9moC/fHH7ZayHBR0TPp0X8YLQE
0eRisu3veWr5c+xDEWBZHHSIdUgET4kvkl46lNR6zFbDkPA2VQjTBGQBBgdngTr5WF8XaiSSh/ry
+i4QV0spE3zylnomw706lNvlLCrTMLmlxpM4TmbIHl9oPulV8sWuCDPaAjUcH/zGCs4vS4+UeWk4
BJGzYNmQgQ8Ex7qozeDP80gR5QyeTqF8Bq7vdLz2jMQTxx/SWf7RwJp+b3jn0GQhMNoZ5PeIbnIW
i6fvfov7sX3PqNHqP5+vO9hchpzIvEUB37Cr73ZiXYcNtnm/4gC+cE+AKzbimi8JMHoC9DrWM5pM
FMuuuTArj59ZGEopeNKs8usV36ZV9yv9H0+eTlo4AutjvmmY5qjJjozRvWpY+pGPivyAC5Bhpwbf
4PCKYA8UYY6WtV/aiBuTVLkpY0w/BMMblyunYBIkO97Oj1JuFZ34NUJ/wSLPlTK8ItocD/Ke/mv/
mP6on13DxzIBulsvGO1m8uhyZkioThbYDnwevfm4upXznB8QhPPLVwpCpDsHF8YnLiEt7LKOrjJo
PlfpPlj7qGUKrlavMA+r420IN/BJlLGeJjPmabij6AdKrgxBSYRkmbY/bWmcKjv1YehfEVQTxkNK
wBvVI4/OfHc74YcYQcNoytIfUMZ/jAfXB421rR5MaZ/y5BmwSyHX0deSAPBYer4N4nhk/azwZAIY
pYxcjNqc/paPOlQmmh6hjk1zl6aaeagzHBIVCZop2Ytts/T8cJekmryI5BeFX6hrRSOiJJYvKx5f
7Gd6xSE3VeQkRLxblniaw2iG9QEhtQUiVvYziB1oVi0RQsjjfKI1UDV05DPF9oj83CXtOSOOjv42
MEkvbxavLBZgHCk8IlB3qLrY839EYbqmc6j4EIE2LpqsjMPNQFraq4lrXGSN0RXceZuM8egfWzpn
jPjyWO2I6KiqahHDxTINLFkei6Mb/7bXL6za71Q2XFapx/wsDvkL6kE350Kpqr1FWTQnW0lvUnJc
YCgv8mCN/EzZV2A3XC+D96xpm4Rxzb94upF18eyhYSq8e8PiPLxpVIzRjGkf9ixjirSGUVxjGCDV
V3JbMdq66RvW9OtZ07DlZMB8sTvQ2IAwo8NKLvZO/wPNwRv2FBp5V+g2eRdYleS15YK8CNpcsdr1
EVjWCTPhJ89jSwVQqHTG4xyAGetktrsZ3pTOTcrDi0so0rHgClO2VjvxhtFQYkupxiJw0UZ+RdzB
Wf3Vk0x1yh17BHwMKeXL3PDQOH0JXMKvfes4S5EGhXOuuL8G4GlFNltOaxlRLzISvkDYQsMvopmI
I4EijXUTEgEWBdIUZY3wY9x1Z99+Oy6Edc9irET4fslXIuvRxgIE5glhnKLR5RYVlCrdSY9II/bu
h616qYOj0KmhwyKIg5H9rtIP7bUWTO3TbhwHLbiJnWNC76NqdU4XNaKT5Rt22+lVvpPHQocXK8Pr
4AuBlzSyTJ0zaUpBtjcNm1XeLVjxenWmixkDkZY5/d2EU9A4qvtxNAoa4Dy6mLpM4jXlxWjIYz1s
Xu7Dop+XklE7J7Z/qzdmXi5UgeCS0sL492uvlDt+/I5gv1yWHEILhlaK7RlklE/jqA2LoDS7ckql
JHqBz1ixq7ayn2J2CeKU3uA++Z0QBsDkcom09+t6W6VwNms2NX866RIX7aahVUoBdnPy38Nm9F1C
YY1oA+zxlF7gRZWEccuwzu9kuhns2gez9brYenJ6XfBqYKelBMg4d29K0il2g4oFXsoxly29ZMk3
my4fJ2v3omGaWQyyiI/AFNifNYVw1c5AJ0rWYH1GUQhYY/M1riQwn0EteTtQMBKt6QKixvKECT8R
pu1YHrNYXqskCciUdYjEaooptP5sx1rEnQat7S4LbGSWYVnvUgRRwFjlRp1S4hevKBhDEGh/Vxwf
MUUD3xasur/13lQOfAZWr4YpzhJ8eS8V0x/cK2j3Q48AVvdpobXhB1cZzBxp3Bq393BvzmNqrJF4
85UaccahIuXKunQAzm0L7+DcA1nt1HilUCFyoXEqOaYd+VnM0SeasA3yHmWQpAd3h8IEjlFemACU
7psxtivpi+Jz41nIOtS565AFgFwrIWC83kRWmqJrFEHzy7tI9UrIGXB3USGSfVyg/yQBC8ud4zVp
6qd6lWbGCwao5O4oawwg96nDNAY8YLQkhyG08A8EGtuB0UvEpgRpFIFCug8lYBeXzVPj8EIEdjVL
NXxUplmpi902WsHDTcqkyDux+iKUFMqob75PAOMvMa1GPYJ7kmhxQkZ8x+WllBAtlF/T1SY40Bxq
AZMfh2SfrwYVMnTvvUFUZXZAuT87XPk6HIdVl/KBubxFkEF5DmIBTVViGe+Tnh4ZbpNXadlz/uhg
yv//Ai5YbLwMtoXfbCLH4qUD0rBMa05y/DQ+k8zbytvOZGcor5syjEtkW9Tt/nzxp+seO9WRvQcl
FE7UyYrQeoVAAO3ohpHgsxUae0oLYbl4hj20yi3S2PlvooWeWd9jxO/CWyip7lZxzfITPhxrUpI7
6OpspJmr27w0VXw06F22OuNzo9uWz52syniPxF1pZCNPKxBradeP77m28A6lIcLb2t4btsOANz+D
KVhbyD2g01gtKgRzP4LwM/pCnnPrdVCdvuIoDMwQkl0fR0od15Knh7mCW9u0yLrZF2vzFB78qebj
WzI0atOl32Tw1gcrn6G/FOI+S1myyPjfJNPS5VfPzvkONHUvnaRqtFviN6LFeUGUXnw/C1EIuqu1
UxHKHQXaiqZK+kqK1RmciwMBHPKjLjV16x+oi2+XXw/vK9NQEeX4b9DvzeW/x1a5AuVZI2rQbxWY
EI4Bm5mwtm0Yn2Rr1PEh7nkfaBEMRQ4/X6edtbpnuSFgTs0UdcgkmtdR4Rg1KmiOm3u22GH8kUPm
BMzf7zjXdfkEyGLKvRK+xc4An3rJcWXhKu2uwU4Q1w9jedr9EJOeu6yg5mo0neOUaIYv1GqV+oVj
hP+j9xU/e7gfSd9EdXXgpTUP1nkAVJBjMSpm2q33adA0vOgAyDqHFj5rz/uGY6BwosLkaOJdCDXU
kCO/vJmoQOk25Ce1DDm69PQOBwD3eQFfJ+2dHlw+o3DeZpo+5e8jVjwitoOJWLAk3UoYoETiyBX7
KVED5ma7wVproS4mukHU55DIp14pGoAYPtGvQgtvbfDsb0II0jEVGH9gXbomN0uKZQxrsaBFSrxk
lJJ5E4XPzdF58jTLpGnyUfUqW68k1vTyaYLCahimvD/Zx29hfBLbla3SaZvqyC06KM1mvUyTuXWM
rSvf3lu8JnvI18sKU/g7+jfjT0qAZ03C8aW0b9O1EMsaueR0eNPM4Ir7YYT9nRHLQWZ0UJ51QmT+
NSN9/yMVZkIWDMQKfSE0JFUK4hZeSbIHBzxgIKAnEeWj/zR4w/N/nEiEb+f8DvazdWa3NdWNSFkR
sucAb7DslOyL7sJGjgvkiaDXNoxt0TMzjXje8PliBRh2N/2AUyF5xKWZzmXFLYXU/MOifdubiG39
fcEgidsyqFpS4vI0YOldwzbb8dMQQq92avaoe/f/PCd41speBiH9J5p6c/WXj4SluvG1qsOedCSc
X4rqj8rgC50wR36ruNzfX75S/1RjNcZXoDBlfQaShNe6tdguPqxIUVcbYzGHulV/zwybVClY56HT
a5ROiaaIN3+xYbPUSS3rHbJAHyFpCs7rJ6cCFVFmMgbRjx6CGc3WyyyUOFjgtuum3aadcj2JVXOp
krAoqG8BERrDCarUI5Hub3O5DRZ0CfpRsmlyg667jgme/dWPx0j6oX0jY6JKxT1/rbr2wDdBuhgY
MhizhOVR7FKTy9+yRGpBX9UlpfYvqSGI4pPMqjOVgRBsIIEwpAgQPAWx0rKP8RRH2GK+0bdTvsDo
J9BbQ/ymIwVlgN+8IgRLVdZdRkkrTOVOz4qyyx6FuY1LC9rtvSdCJ9OVqdhbmzG9KpDVrtfKIIBB
2QFcJO2iddzS7lTru19Lw9JEKK2QdK3QIDmtncxJvHgweenUitUmAKixwV3bIMzR+E5on2MKmtls
gyeJevp/jZ+D3o1qwWndkHt82BypmaSqbboCie9YG7Yehlo5+gvrPHHWCC4PmdSQpNC+w6ZIZGdD
edK8vSINp3oN5CAF6iYhq72FLiEdQVEnGoqiagOKc0iX7dkZSkuKm+LW2TglQ2fxqaeuXjRhn4Im
P3Yx8kJ9H0q2X3qbPkNfj1xOqu5MxB7SY9vOoOZ+gO6ikQLX9GqZdZgkN++yYCt1QOQdOTrZGXoT
wTB0zoIhrBZV0r0Je4jP47reHQ+2tGgVQ0D6OknVsCEmbsAEVjWBX7mJB1ELbRUNCBP8C4rwD1QQ
JV5FPkrWy+5KauxkQ7OQ6wHQ54VKOOM19FZ2ou9zKo2P7UHOfJOoRSHRQ75mrjLGfpqbS+tY/C0u
sQHHxBVKFlukXucRa/4b9JbJNjksg273Zum6TYOBsGk6u6A7ZfmoEdmD78AxM6PCMhA39+mXzi9p
NMuW2hNOl91ccLVPr2dzhf2L59NssYFOEutDVICoP4dcnbRnOzXh8cBBgWovxcizi2OZpy0PoWUR
WeyNbGeoxLhYPROl51hFcFYynU/RyIQJCeInbEhdOBYMFwKFMwaKGV1xJfuTEqX4N4+W5ZAXJfhX
4Kub6l18fCr6ZldO+03pAGEhQL5sJoPQPhlIWNam9nvjJOaUhykFD5T/qLuioSYQb81CQhAZyT0L
jZ6Gpa1IYOHuBvY0/GFc56yCW2Y1EHGbSs1nDXkiyneEKyaCVkl6GFIUkTLSb3htNjzNz65Gs+sS
kEHPKpCvbOvbB+36Ib7AKrpKDG2sRCQCG8nOr48LrJ185n7TmpCL4zQ7EsbnHS4OuIQslUtquj0F
hdn+MFirNyG6anfknnknzQlTaQsHs3BRgpLDZEuau3dklfUUPjcss8U4wK4dMg63scCrUHa+PKTx
BwtaM9Wakw7jN/WZtmLsUjDowWksULq59fF81HqN2NkpEiCKo2qC/lgzDqkahwg5Y9EIIMiZSOyz
d1PZixwoht3m48lBRT9k/4On4xIb6WEZSw8MqMr39HQ9qGR3YpcXsvPrqaj3G+ASP6P+cGVB7y/X
OVMN5SiOq95i0VAqDs18qDcRSgwaKmctFAhP5bT5gIPF26ZoFZ/wOinwB6RqqVz0drdCx23joHtf
y0lp2VmXquDAwlC2I2edtYr6wp2Qdw7XD131I+Kov67RzqhDXWN3YIJMKWEKuLCOfyWFrpOQhmwB
nAgjVwvVDVTmesSBZdi/j8vF1Z+pT67NEfN5pNRvqRxPuj8pBWvNYgstCOXC8F9ijlIxGY+B0Cf4
1T1jqg31K14g+8WHW0ierGCgCyFg4ZVdiukFF6oqHJIixJIykUDSjsrsdvbAbsowczSmM2OWjp4Y
ae7qPGGvzFcpdLyWv2ecHQMAfw2gLQyNiUNsvVGB9sOWYvV8BgJSNDfgk245XvdqHCt77+Yd7GmC
ZRcYfwRhviq6jV6wl7R1hix2maLMpFzfjJ36s0xjB3Qi+iNBJ9lKQOzCwuCdFAJ5HvB8dDueK9pn
pSmY6paQuUdBrJSw/1Bq4TGPOC7DjJek/1lX8+OCS7hwVotWnIeAxuzBUxWBUTSg+Xb39qj91ppv
gyk6ZbguAncyx/sIgcpz6YRKobn5/SmvfclesvT+c+zz8ZI9GgrbpyCaIgWRfW2fKcA8jMn8LTHB
vPEXvm7TUe89lHuuq9dOkPBRzECNai8HhtpkUXhN6yCAOPk2RblVXHe+4ZPPXGYTGx81dvXrZhh2
vLTPqJlBv7SKx8NOtLEIkjhsd3TzxMw4vz1PNPHaM67iUQdaLYS4z9LRyiYrkGqfWn2gis5sbt4W
zZUrrWMf0STfu2topSrVLlfsux2Krsc5xNbMONXhnAJAhhzysUDXSSfpfAPskm3+C9gnyCnTaSO6
tivCYJRZjnKsBOSWk5BfPECSY+nQ2tKQG4JlQyAqpuDEbzgdqoXnmQm05pDBj2fdCo3UcAzYfz28
WMJOHOwB2kcvg10DBuZsEPQcuOwgz/EPgxlDm2nC6iS1M9cPc4o6WmNZF9IU8EJfmLKgz+hGhiuJ
VvJKGBiY2mgTJHbmtojDsLNhJ8Tpr7c2flUGXbjvWrcs+UUnRfuYsFiV1mml0KH96/tR56Xuw0e8
dapkj8HzLh4KU21mZvzgRABLVANEtZNnxDHOl7bAiIO9EaOwnIsXq3E0abphDNkKJgWE76fgaWI/
te7xX2/2f753xdFG/K1JuL2p5NX7ORVHPb/oOb0w0tS0u4Ve6nbk6azl33vmqHJDUn6l5vAe+Ljh
ziUSthzbevGUCe+HV5dHuH4ZTqgV6e1azqpvHw2HxAljXQGrWVbOQHz+VaFHDBYEMrB0B8X/Jaam
o33W2aN7gVk9xfuUh5r1JWHMFcCJOf2lEUk9vqkw6IGCXeQb/0KjiuI1c2AWSVaUJV6bnjbWU5vA
ylqWDFiQO23dOz7IgBYvOLPJ0agBGaY+K9jE7HoW2ImnxyutS3roLS8rpSmNViGM/3jFLKqM3k9L
JvP7xtG1P5cXOpBDaZOKv+I5/v+iaj9MNEtVc0s+BVgMWchgqHP9K0WGqYxDbAz2VEgdntxoPnTr
/gQkwd1mX/isQNpOtijgei9ligShytFa39dNJ5lKS5OboAfixfK0SpikEhqMvIoTOTapypH26tih
U68mVfgteFjPn53B2v7SqEASQG+qoiPWFGBnZX2mRFiitile0RK92hOb9/1AxbFUJb5RVhKNbrdU
OJh8SYpkwl1kd0e7ucY7czWU9WMH+cgD8YPiuzeF9TzaH/kLsVqTBEDgLWqx9XEYQeeQTuegXFez
BYiOUd6nRxPTKth4WyKH5VaZHkePyfpPTJPR6EAaoj7CD80Yk0E3iZjvVFuFg8Z6Xr+N++rakb3q
CZVWVJmZeyI/dZTymjEVnBGWC7tY6j7OMzWu25OL/4Ml/S+zGCUFHkt/uyiC01pl9hO0odx3fbg1
xloE5LYh8sBtfWZQrZrSXWGgWk9o6yQvXTd/ZAZC8JEaQPOkHQtQ2BPW35YDlqm/DXABWRBzvF51
fdPhoVbHYFlecpBqfaUgrX3UAGfCQPmwJ8ZB51XuBiznxjBfqTPqhPUqXMG5M6EP1MGKjofyOtPv
usVP1V/QBok7xm88Jy6f/+WwW/tk+8E+x/fRGueJoNDFq7QWg1rhOwn7h9Ob1wsn4e5mxPQ1MREe
WP+80Be1SZ4nQZALC1WSjPvrOsJnLAm+Gbuq8ogr4ZMc/yLb+wKRhBSZpU6oT/ZgbqV51Fv4HnG/
VcJQyN739gwHpWi3YZgHKkN1yXF/pV4TuShJnZSCy1Gqt2obZkgTHijQCaEQmv+f/CYhlAyuxd6I
XtthwhZPKRmJjkMZr0ruTGvX4OwoZBNUCLr2b1aYrpU+yFBBI599NDN8s3K9BXMqGczh5TAdiLnE
7O7KS6zlkaJ1xLhEYVaSGHksf2mX12mEytyc5FyX/Y7d6n6YxpnRXhU21EJKuu0qc70TB7P4qIIY
u74wQrjqvmVJKXcslvoDglhLJv6RGPJacY8bYsaUlQnlR8xm1SEZzoKDc0/u3GUbSSj/gmZ804yM
oDjvP2GzRlhmVTPzuaF2mVLs+tx26pGbvuFdA+T+8pg6p7E+AuNBaWwgFvNFSno7lXi0FhWam2Wo
3uheu14qhVmDAad3wN6J5W6Hb6iAPFon8g7lgXF2H+ui2NrNnA13j0lLeXD9K9CKxZIh+ohWY8Ar
dojOxRrdEXrS7re+lm4pkQpY1rE/489FhguI6+dKZ1M9M3SwUWgltMo9QUen2AwdN+HEidCJafWa
1oYEU2uiE6OsRdyrh5p0zpJNFjW2TCLkyVdij1GhGUyYBW0l0bDEK9ez8qo6btG/uA5bxI+gqUQH
567YosAqhiw+anqNR/swRXEgkOoqXTREkJcHPACvwirBICuVCKPPsGGz4bmUeKcuyYXAW29/PXqP
ZAHrb/GYDWj7ANbdlCdhCGaBLJ+c4zQQjyfYBlgbFRbG5qYy0hunC5VlUq6YsogGLIltMGmeCEdW
XqjEPzkdTJLX90h6FFOkkmuFK7J05PvYLLcQFZ6BzCHEtCdAqC9fqizyHXm1BVEub21FoaxGRU/3
GdiIHxJpLrwO9ZeMMHbnFEEuKCuQggJqYfkFNRmvqEth8y+g2cb4nMtQvEABqSMVnKoNuypF13OE
Hk+CoeQsixVivHSzBFQRYtOgj1n4/WeJXwZ6AqxbopCQ/Z2PeAjeeSyQF8J5jkwmUrSs0ICat7c0
C32LP+ULX2pVh5vTqGDMK+QZNEAserw7mCqNI/40+qUDvLChLbSYKlBXSieogX4pFZlQpIq/33mi
zt81ofeCVYQkaP4qyfptyu910eFXkyPaZnVuoU946wTEnl/iEvIXOcKiX98nrDqcorHMsE3bKHGY
SZIQjdTdpJ6C60gFxJsHxnXAb2I1m0phUsphHuZXFATv5FgshaAre0pgJb5+ZMN7HhkfDtsx8q9J
SyQGqglhd/amYOlzqy/toqNFGVv3pcUTSImddOdyqGe19gwJ97iK2c+9uwQsn+YmOcASUeCD3uQD
MAt03bzakD6uU1ptRCS8MQvKrM5Ufuldy+q1laydjRv89LXbc4IJn8yxWo0DK+Sy5aYngn1qnMdz
VLpHK2KYpPJOkH5WjkYFcD16/iEjZE+6ncdKEZpV5vuvlIlNRHT80HEFIpfD16MDmnUpDt28peWM
PWPpo8sOPMGgAIFg1IlqIs+zW5izjXfl4A33vf97YGdM7DXKhZGZnFlB7SY4ZcT/iIk3OyTq6SfI
iyTL2Pnws/HpLE5v/jwpm6853GFSUto42c80LAyy2vDvnrdcUdkHfoBzgZOR81I9gDKDUqhCyyxc
R9RkDOC0hV5jdwZN4KC13M+INjNozjuGpC0uV0bBa/t3qCx8RSIWo11fZdBiCGGvhQUeXN5hWtrL
Pq3h4bMJsbIhp/Apy872qhfM+Z4CcKU/aBlxiQglohFfN8GlDjyuuPFeWkiWzn3Z8FfnpmD22Djd
Vf8SPe7qv1YnYffu8IzlPnsGX8ZG1NwdVtNQ4sRxPYKa34rISQ6eqszArxXiiR32kib9Ox3KVL0I
1YdoDHXUQohd3SjyTNTDHG+5wO0t5CAKKf4hSoohyf1hUCdwqyrJwYFw5gkaBP1iSctdXi228EuH
Wku20vH0xER0oxhI58iE21f4y82CxZvMwoklH0AlP5BXlncETpoPJOKkYqEm9vU9lnSuoaX/hIh6
IFmc6aqqBQ1FmoAtjjYTZw2ovHLGycS/pLeweQDuirZGpmNK7vm3hOalScYCk1ox7WXT1HgPKqdh
rX1P3SFG2PfyNAnNCop7ftcvmVi1RW3V9e4ZHzj4l2RtXGY81WN2XyBcxUOhIK9L5ghx/kkQUcU7
sJ5Iomr8JXcGTp/Fso79inGw9AifpQ90n9FVfUomQzoegDn3l6Koezy8orJO7ycX5tRViJIdja7T
qpLwvO0tMDx47rquEwOuxeKrtkdSjm2fhKOcp1HQLjjCaEEQqNnCwFrez/2rTSLSCi21kQ+7F0SU
n98k5hIKMr8BQvXS+ZZSSi796PVBX3ylhOWb/ro3kd3fCvO7cnV+JmI1blAhFT7biBJaPyPaOxHA
aJ9dZL91yd2G3ttuRILUKuSRD2fExbNg+rzfxJDTFMU93sCReRnRLrPVF/lWDX63nJyPPdHQX3cb
q1IXYtZYui3lMtrNm1HbbINRWVJJN7OMIjGdnrz3QBwUxiQkG5mB/5VTrmwnLX5e14V1496rrpfR
01F0bGZqhvc8v4dyOq/wxxovWggH0Y2CNK5mFYp+IzIgNYCRi74wRoQEmO8iq28lNZIofIeLWOSX
Qd7vZZtwhah2VzXWAGhW48MChLUxJ6Nk5PcstOuT756yYUe0EUrLEs7/Bob9kOYvr/XXt9uT1Zq4
3oQkK3vczLQS7pkHWK+oxwqIHNbB5ptbeLLQnTwaelInainvJQOIfc2IpfjyqFLKkt6tMJgKUfj5
y841Fq///8eFboMCRCMfG9UQ336TL2aBvtwWzolu92jRKHBaKdqRBAy+evlS8YlvXZ4+IA8av0l3
m1KwSnIvh+b05JQle4s8gVZ55X6xNftwlPIpSVExrAl7pAZ0SXeItMUSTeG33rk/TawvYj4+fBDr
cavola7cVOi1qNwVaVbU7K2l4hX7NStf0ZjT6CNSrPoPu0Lc9K0pOEVZK6zWWs/DETij0u0WnJw5
IejsjvAVFdBXgfZKlxeU/cJeRYtOnt3vgBaHPOU7wMFmSjj+cy9AGZc/3IJp5JvglLZqYVAOWpnI
mT3NtPVndPUflejmeJrbE9+PLT2N4Iz2cuqkv6kzbjQGDHUVUfSt5Nvn20KqM9rKal5U+mFNMQBK
kyB4ypaqAYKf/uIetjHaBJ9rPKVjvi8IIYTyY+8eid2HAHVDem0f0q9xaU4gRyybYRo5mClYXX1D
IgMre3T40OtmjeVMK3gQgueP5phHssVS/11yLOtZz9U9bhe3ZtT5Q8KijXgOvFHV6U4z2enA97b9
qtFkBAdGAMWvavUZtHN9MLgfTvY9eCPfU/8WxMP3OV2efpgjf1fzzG89r9d+kUptgsitb38W5FCC
/PL0mobaWwaoBPF09vbipipkC7bWIIlTCc76PAxYDJxOFb6zZNAJnb8Oetd/OpMuHbMQE/kQBgle
kX6mt3hiIeJalKNb4h4Ryry1vPbdvWQSWGeB5XP/BnpTiwbcAI1P5N70QSmnq55MBKUbbstyYwHd
QrqaRS5xZDTBrLKwWfc2jaU3ucz0YCDaxrxrzPHGouwkF7k+h6ZvP9ihx4fTLOSbNtBTMWZm5g2q
qARhQ0VPvvHBt1gikHGNgGNAWyhBDJy2mpJWvHaZqghFrgoQ1BfPx/Hu0yIR1mQv7SjNuUJObPJC
XbeRMujuDwzGA8vZNx7/dGuGIQjS+VDHzlAXt64qpjmI4bAitgvl5esY+QZH2+qFZ6g46e3HzxPh
WHdNpKWTG0SYQt87e3VlMqYBgoDXh4ODRBVuRB2/qKbhzbEif3VFC11U/KifEJtNP+Nhl3f7ow7V
F/xLzxWRZ5Ck867j/4n/VEJRf0Jjj1p4vasoZbpHKoC2AAXj0vwNwUKfbdyY6BuMBG6NgijiXXWR
Oi+OLvESIkn9PZrc8IKkilBS4U4IEiElWzCLxVSIPBIqOTLhAZNj6HbaLE6Wv0JbScetlTweUsYx
X0LOJSVthS5goJapRgtEqH7mMNR59YhzNqCJQmbvVhoSur8QaVZ3pxLLDYpGMZi/4sLUNIPFNpqP
JqlDDdBFytMOyfEhHwZw28FMPcPs1hfGo0qykBoxWgN4nUB/ynu+aU5G0MzDqEJ+6Cb/IVzawJJE
2Y5l1XI9+LyivfyOKKozwQh1Tt8SVjZsCaC1WvIWDYPGbUlr3WNUqtMt8eP891QyQ1IN22e/b0tw
Wrrkp0sjmhYJRZosKb3FpHMoH3qSTk05I5Lyf9kijndE6mqSBsWqIqcCkWvjVICV+kzFrj5T0WE7
2xsiVLAzNCDmljZ/CH9PlfiTrttXM6v34WXwFAsfHUsVsAnEIiCESXxpUHOkgU3n2UCdPkNxOEZJ
ZkC30jzbnWu98r/xhoXnx1EkFsMn9sj5J7Y8nMcu0/1tYSsX60n//hOI15ft0RmxdjXoT4P1Pk9k
J+2qcoJIenUoagLjRbfdtlO4Zeou7pL0md97kfijaD2pD+OjBsaZmjksnni5WR3wZiAU9KDHmMYt
tQLIsp0CiNgvZP9zifDogWmS+1wInxzH3uPvwLRidCxAUzVi9/gfOoSFKxqmMDpn77UqKE5qs+E3
c/D+kNCn2cjq4CQe+7tMSAk7BlDR7wccyTjE0bKlRbg8DZowaZkp8xVAdyyxb/f44AUY1Dahyto8
/a8uIGPsOTc2+xdNZFusz+52hsllMozYM83olEmGhFH7zAJlqBKun4OWQ0vDsajpNQ987kMsC669
XYwhyxE7xCD4X6rN52ipO+MtIYHdUvT0wDJLaL7Qp3ou9w4UWZLSHc7FEQy2lTW9OlkxN5D8aUTW
XoBQDamYziix5hpPsYwvl+7Fnxy5zOlIGl5v4qPfQZn4RM6zSdOelN73bComuIcrUeeHftkmF+iX
x6mDC/5GioWOLkjlBxhY+KYFMSlhWlHJKXygyUSStjE2EWFlTIPSV0l9o15OTcnZaiUZJdnO60XD
mo9jjoe0d7PYA1l1ZnjPhbHyw5H5WweTG9jgqgHcYMcstxeZ1qIeuUGDGRySv478gojq+1yXjlY5
Tzk4z/X3ViDlCCpbAjtNLLVRHri5cK8bQ6zg6hKKzGZ/36Bqe1JsVY+yxLJGtCwxlnF4pnHHR94i
x1oGSPxLDwXh8T/Gc0dS2t7S70kttZanoIwYLHQFskMjLPX85a+ZonS+FSTj9b+k1lvum71vLej5
vvLSbgKQoWxQ7qeeY0FQXZ9jNGm5qMf86PdR3SlSvFEpgBOCyhxe8pkYqIp0TrigKS1R23XUl4Sw
qUgtG1AGXRL2gjxreF1ALLTZAD9qLzsFcRZxqEFzjYEpN73wGWrz3DxSSVBOsPWltiW9egFJoMSR
Vdo/ixzJW49aoQqjLd6zHABP52f/0/67+oBbEsSmbtFsvA7elBx0iHdlz6fsG57J2TGjwUBsoTzW
mOWSRKGHg2k7kATmXims3nD6gu0otRV/102updYBgOf80yC2RUjoB26iEouwpLOsgLKqXh9IRZaI
UEeSxnHUSnuXqFC4obl+CaloB4IwiVFHeQU67Hgoi54BYMl3fgmqIk29imr1m9pvoPJBdUrBZ1aN
lfcFzauFPmIaBFTHtxvwwTJiPgcsYwnkyp8eDOYJPSZDAO7FjXaUHF1Qm45OKjgg6xO6/nNpI6W9
fC3lWeoAl8awKHI929VFYQ/EExy9w81XGr2lH1X5DpcsfLA+EPPVCtgWnP59mdutXpKd9XDBdEBC
y4zj4sivau2diCuiLUnOvwpkS/fILa814IlEQ2Se2jL4lAOWyCIQxaLYWxSTdW9Jiswe/+zZYVGk
MOpXQzIr3/qIn3ygk0y+6dox5tp2vBswunBA+JA/+pHGuhKwQyRQVgaOjLPrSXr3TFkjejPMnXGK
KseJ/U7P1U1AW6gFmP7CrJ0GiwEnXcQNFqaVDWX1pkWcFKYvR/oBMfRea4YTFdsoX/FZBnVwzh5z
8/Etq0PpvtZSWcc2fZd5NbsK81EApFHVz8/nI4B6uLI9VoT2MGooK3x3mJA+9/6GpexWzLprnvli
rSeM6vlkGKqA8etbaLHhvG53fIYUtFhJtdG7ks6QOjJs9111cOZU2r1w7wEb9mQjnVH0zG7gM+jJ
tdiUTz107pRLRZ/K5birjSEvmDbtIFaYYJee00sTz8m6BOGw+Hvqv/aic65RxAes/gFJxhh9A6S7
Ik9nToQsUprhGtsfDx2L6iY6F6/ES9r/7pqije/wGLpdQN974uLfQ31WnhVNITDHyIVNPgn2/78C
ZSjAIfT+JEZP7fy/Wnq25xA3chyLfhSKB/Z8h9BNcCELM+dHCNlkTxly1DbJSfuzaRhGsFFzo8vB
UytagLX8Wrw+TM2licSCS3Rm0X/seXA5UcMSff/Y/+7ajmov8Mkl1upOVcSOWXFgxEkfYdPsO2Zk
FO8+1Sn2Ci9Dc2B9RS85bfmQrjNAZxFaycA3D2bqOyOVVHWTn2ksvhHO41nDDgK5B5fbF8Hb4cJ+
+wV7IOfaRsiKkqt6PmNo/dz22o/j0Vfiz3stKmEnNuQnQ7uCo4DOzSfouUQH2lY3UdWwTI1GnaEJ
bUvi3aZnw6dstrGB8OgmYry9pIqZp3gAnkYnhydqKVk6GG0HM0DpUXKWvgdYpWWXS3dPNKuxOO4o
POMAO3ZW3BicHUDSemmCWDghBAjw+YLHV/ilL9VQhVxS7XO/8BY5s3/n/EQ/2nkpDB9Po0TGqgLQ
yo1N/Dnwdr3hkD2y+MUwasmJcwIqJjKBYa6GE7jc9FSGkPReeANCDUtxDQvKvKQE6kIrB+F5bk+h
EkH8dPOIQMhLbbXwkFOBieIkuT7U97IVXErWfx6pToz0s+cThvgH33aSzNd3cZtzYu/M7MfHmrv7
SKAs8wfYi9Psld1v6tJJbZv/Q6+C3zer91WVb2mY2ynRmbVvITFIREhhxK1dXNqUDY1c7CTDcqd2
zpldoyg6ip3j7zwtc/AYj8OhvbDlddR+KFDbFmV0PYreubiSUy0r7hch40pRiIk34TkJqVGVKY7o
v8zughJNfRncySKfTvkR1g0cgvKYhOB4ZptF/xj3SRNh/JDu6H3KI02qvkK3xt/G/W2s/chjmKax
wBFkxPfBbaOL1pobFI7s5dGvxewhdd1SNw+MMqa5AhIvtp14psLBEj2lMxCHhasF8LRQJWocoW7X
1znVhmZUFmEGg6ehSVKNqxJvoiA5s2bedjHhdAnhTlw5qN0GiYBj7b2x4Con6MhQ7+Z2lN9ZW9tA
hZq6ZV4vetgyxr494XGHJoorG424mHBSyNXomke6rzu+1mHJHrvlwQbK0ExpSZ8k+GLbq6mk9jBT
duIV/8n0lJYGLhR8Qx1xTJWe3AqLUJAGTDxGo/YVzMOsaYUryrj2EzS7ocugNT2AGvbBMOW7ODZX
u06YuEVVskGwgvXEnEJp0vFv1i/WYTnZd4i2Vein99liyhu4fZERA0dqu08LX7p4iTvmXdTAIT8D
+QxOHHgFjNAVYNkWLTu9O13Q/HGrAmFpdWApOPMOamfiAzTJDSJmjSKIc2LV5BRpfnFLdQM6jETC
/ltETODMsNN0QPCNuSZn0g9d81LaTk9c7w+aDmxF+ZxY4r6MaU8IGlN/fXs/6wDFY63a2gzsWF98
hMEAqvYszTtDbuvqob5WX/jNBvxoPj7akE3BZLZktrSItC8CLG9LKYnP+p3nAO4/lhk+wmEIDpiH
QyER/jfh3Bov0+8Hf6ts4aCQ6WPSCypaEJgPfdPZ52nSpq+AgAjOO8Ie5byUgbGHnMiSZ3LNCfdd
bjR22lJG1Dh5p5Hd4UrWKnkoD1WtKCiqeQL3sf9NwXdPr+W7/MdQQkenCG7PANtIr0eIkh/eJL3S
THsXob3Gu+VSmusVYtg01Yyzex0Z5F60KqgWs0j1CG0Rd6SKxv5/BbXSNbv2FrnozzNuMiQAYvvH
lShatCEUpAf0mBd4DC4V/hBZMWITvMTa/NT1apHO1zXShvixG8IC1c0cMhKQ1/3Qa5QvPbw1MwMN
wqX4gwcjWfh8px3PVa3uFcZeNUBCsXRHhzGTW0PA60o9optihoK9908OOV21htY0+kIyludgwUIV
XLUztMmmk0CFGfj6tsxFzj8CT0pf7ldy03MQuRkyK5UTdsVqjSVZvNzDn3V9j41G9TbD6f6ZR3PS
kTK/ZEipB8WOq/ooNTMOiMzGTOixoIcgC+iT0TX6iy1X0mdZ0lU8+hBcw2G4eqNnp/7Rjx3LIO1a
xff7L7AjyjOfuYk1A1DrYsGwI5kXKZdR73ma8JTuVAxHITK7CBxCjbl6dNt2YKVUJhf88a0+5q6s
EIzNjMiIrIwxBYFd7U42wlIu2C46soe756j5Sqm8upKxB4da0UvjR219/iceW1r7Ha5W5K1YwP03
4eXkl85HZ554C/sDMUMCtwZuLvSLkDiadalfUu4NRnM8UHvWIg9O0VhHy3i6dfy897ud4Bnz2A78
/3tFbH9pZmoXL5zZIFptSu4ni+cCPTXvwCaCLXOm3AMFOffcuuQ9TYtdPOojjGua00tysMVHRyAi
/GSamQSzHUpFHrs8H4Js17rRnGrjDqi0a9O0qzqxyDtelZJypviY856Itgyzzsk58M0mJ8x+LuOY
JY9rNZ3PRn4LXshcTBiI7oQrXF2vFtGdihfp0u83BLhL9WXF/lonAVPzJiVLSAnaCBTh8Cc9hViY
LCk0fG+CIw/PKdwX/+XkyNepWyLA1HNqJ385NmqyodMio2wCitBLhqa3gtn++FPtD/V4DoPyLc+P
o/6o/0NnzUqa3FPmD5wcBbyYUuWEoejS5fV8iIHacNKiaxe80mKTsTsKtVIcoFJOrqnn/KhI7sQu
cBFoZnz9y6dhjIlQzp+N4lCT+jCktYV/6IAZN7CL38q7jR3XZ2nX+y+Mj+kmHDlgOUElBGO2Q9pJ
6Vhj8r5+xfz/p23IYUVDfktPFi8mNir7E2kapXnMl7A5KUTrfL1Vn6u76BxxZiSe4ehHqgdhMEhs
Zc+fhxZfXi4bog3K2t3H0FUFPnGUom+JND8AwQK8+iKYMOOh0BTl4tQntp1WFK3jDjRbI9nIjOwS
FVQKUiTctyw0ai/b7vo5UVEja32JXHWSAa6pTS4BgpgQGkIEjnou2dD2DHWaCqghug2mN47TjMJW
mVbnq0n8+alKy1FZbvkSJFtJvXFlnpHH8L0Sdk3M1zE/TDhI2KoKZ3446GjBq01JQQ6BSQgMXx24
wI8jRxzn0dEYZLpt/PFgGpkSJy3iGwvbmN/Hr7keHL+bfPdxwjkMT86Vm8zBpvgAUwKPfOGdyJrk
5DZ2joOiZzbPWwqXrHqCrtKW+AB9Pn6lD883vuFK11obFmsS/ep8ymY5hOOTrXHIHwOlYEqdhHGe
2Vw9sXYR2K4TxR1iyaAZPZxZLbiVtcJFaAcAc71cci2NPQd19c7EhOzBkx6J0h0vyj2Wo7FtY4ej
wKxCbzLuCN5R94XfWKVHu7BTz+KgI4KwrJ9izxjA2wptmpOhQOkgkfwrqmKuN0SJWXymuzzuJYxz
lfKRf7j5thBDeW9pnfSJSRKNNouVON1BDqAUDnEZeosskZEYLsmkGN8QNP3o0zu0AKZYRiVvyCFJ
OsJZIcnqf4vPwX9mEHK6zaHUq0XzXstNW/5arqOLIWTYs8NAtVATxpRaQIlowCEHMWOZo7C1zJVw
h5A0uliUsVXwCX1Dv6freGS5d4BHUVbsX2fY4DRnKhqAxCLECERPcGTsPViitFkCpOVRB8V/js2J
TJ26VoGTvm9fBXEBNzpfW1arhixZyr6bYmAoJXJEMQU+Xc+mBXWYDMlbT99DNAVqOg+Pk/smRCaR
c46YXq6wWbXEnxXLrFVl99Ei+N3WYf5S4q3KjX6InEXdRr4CbaRHCWZynQ4P6odqHmLnmVIGpxiF
FH7FZkJBqTG5hU6ufW0ktweY/UW3wxGuAm57TYdwk1k1xhwyNuRQOPlBVei7UqEC6vpd3WXjMt/2
l/AQRxOf9mhokSYNFRxqEC3vWjWPAV2oGO7QgT9ffYO7Ug+ISV0u1YlZahINkeqIxciLRfVtWkme
K9rsEWk1+TZSHH4uS4A8Dcu2Yl+l6RHl27dTh+L9umUrkG/HLJt0uXhWH5RgL+i1pPdWMiAjWsh4
Vx+TLCKzQxaMkQR71XExEdsvjMI0jKJjSh1Re5uJe0Q1tEpt526yLe55NHR7ZtYDAJjIaPVH6Eh2
mEJPaBkPsC+KV+Dy7j87hBH3j9ycgVwbRy8QQNp9OwCsc38Fje/WWGWa5wGhiuy4/U+01FO6s8tL
6DbqFE0Fh+jnKb9diF+gNu9I6HmkjMx3FjOyMIXblkvzHForwsS7sRCCClshtRmvLrjS+VuYCdow
Fs9p3Skx2oVI0bQXFkX2VmQ/ldpRlI2fQIHD/HZ8q52MbWWBI9Z1KuE+shdZ0znmLSADEcC2dmHS
aDQsEAwQpXF1wdOa7HiXyKaBCcLxuNohOUhuksKfefyrODWUXnANfFZYYmyWl3Gg0GXzMz41zVof
i5dGrf8e5NiFOsd7b5nZfzdCZjN9fnw0NM6RPuZAd3zmh3UsirIt8hIkpckapQyiVI+6sMcwIE+N
t0esVXkx8emtLQ+2en/YjrrhuhQQNJ3EZR+78a6fv92g2xCOSBL2TqxQNBaKzACIpcPklBk0rk8u
wDnjaUQMecrdmqsU2mTYrLm57vQdnp67Ha5bl3aynoh2QlruWv62vd/IkXY43iwDv6y9cDZvgR78
WlVJgqVMLCF/rOlPF34DVHCRRa0nPUDRt+wgrDWPuzIs9KeTesqwYEgUf+wTJztYwQDDuW1kPZIG
nt/sMZFx/z1g5C/RfhjYmTxYWEz0kDIXttxAWryEHiN3HAffHDH5y4VPQXOyHw8O0sEnZBm3up3x
lJMGUkqMvlF+n8sQCZZUF/1ovr9Y1Okcp+vu5Lnlw4ksJrC9wlbuO/5f3KPk1jhrCvtfZvomFeN3
u/k/P7xB3ksYBd97ZikND7UC7aSOk9jRzz0j02qOYFRrYJvjLrJGgtPasZM5At24rdelOBh8Df0F
8/o6XJGrvWFqIkdT/SlM2NMTR7qigAFux8dW8LAOTjUbcanWU7xrWKtToPXLRAx5UrI4Mg5DtWr+
Ff81wFFmHg22Ns4vQ4u++rWe6KNrYmhZwC3zxJJVKE9vm9VcPSSY3poGQzn2Nz1tA2UpeFw+9MfC
rMe+1hguwVpq0A70AbEK8go9T2JJgPzRPl3ZnjuONLm8bNbk5Fp/OEPRjXlVB5vYO27ZY7htvoVJ
dkOfUG+JI5nobp1/+97vsql7Iyc2ldo2Dqm3YD/q0XmBHyu2NT6OvJ8osknh9ysomAns4C3xrIUW
qpGErzqvSyuKmJlL9n6DBcCBIVG1j7NebrLIWvGhjRfI9G6FlvDEt+mmZ4VrgZ7xyVTn3I8p9aCL
C/NlhRsapygn2YqonF+K9AJhlRuaVjLDmo9bkvvYRhUiMD2dRY2TfE0XoCr6GlxJ/COeci3BtNpB
H+ZBe31epzpAYtav7xzXtU8kT8NFuHPpFnlWrv4XM7WbqzGor3CbtyznhOBij7l6OQp7f1Mk8YZT
D57bTwZQxc6Ln4koWTH+/kcnjvqi5LEe8t+rs/JYVNPSuCgUP9tOYtauZSy1WWM8XA7EWcK/IRuX
AN0hqW1psXsJkuqhVz47AmmVa3Ictjfx3d3OhnGrqn0egTUs5iGDN+Ykflmjs9aTojnL+52SG9jS
FB/R7zvNwWwnXjg3rFmWUP7/ihLmUrgqLX04ANAwZxDqQkNHlTCwep8Otp+rPMb+f3zx7YHVqInV
VokkuPrGb8zKY3j0TFj6uJYbJQimEBWYd+Pj0IGPlkX7cE1Y6JOhWWVAFfoB+FBGSObTIVOqSLIT
NN2FtBEvEBTqrvOtH3GTcEGWPcS83IFAlaykeW6gehbPPVtsIHs7VugHgdIfxZkITeAlyeZeN8Jq
PwcgnnFNjigrtZ3Rb1NEdCBA8xQ2/XgrRHWU9CA0c7jZKaz4T+th0WC4T/1891YZtRZ/NgoZEItG
Jr2TYfuM6Swi4crDOKldxVltBDwSjMIMqbYuaBt5zBRXOoTRaGGeEoI6HgX9vGPuYoRMJBTMy4Ge
MDUA63e+/IitaSuHGGkMWx4UMSGKsu8BCYUl+F/ntn/6R+n9uhbVNgT0mfA+/2msMWcq+nLdm4Js
PdDI2+QswXLAPFHbNKHmKKS7BBHwRO5iww19Bi6RWaZDUPCV6CT/KGe36qxJkLz7n354Fs1e9Uau
TiWztdpKIAwiF3yfXlDQLQ0DFfdTDuticTM7KVMeH4Z4ORBOD3jFVlTka4Z32BhhS0Cb13HjyBmv
RxTsqjQv7LL8IW89BHA4bnFfUm1t7kxYWNYnFjmTvnFpAjfwr6PGqonMf4B89iHy3Lw5YC/Dt86e
AVm7BOQJp3fe+HoG5yq8fLEMS9RDiz5Ui28TMHjMNxMd5CHJqzCuamUcXFW4OiAMLz4mZ2KDYN5f
VhGavBIoIjOsLNePNGAXJKDw7INUjI3iVwujtFR4mKSr5l+CbGndy376Gw2U81x/HtyeiC+/c9u3
4CNnKzwAYWL/ajXmNiRz6m4yVQc3/rClPoecI3elTh3DrVS3IZlnxFlTrv6tWQUL9lTvDXbb7I8Q
VAHKmIdbd+JS8GPZV9N0H2A3h6gS839T2tAAmExpZrSBqG11EZMEMcHfT8LsvLV6gkZPisFz2LmT
xxGE/kn2UxgAr/2KnN88DTsd78m4sDj6I67OqHYpMCj42HktxUKTjSwAOUiQ4NolXF9hfTOAatwH
S4rVJ/tHM3eG+gil/jqLcKE/Il6RS7FcE2WraHcKQMJBKwpFgq7yhCa41CMfk3Up7zcFQnCZN6P4
G/JI9d0DMflaHTnzCc1pJt/ZM6kf59jrGoKLYb0FWQT1e4SOwPqFffgisJXkb/VHwyviciy/1PFv
qAN/L3IrtA8/t1yhJaoyFPCvm44TB2KeO1i1y8/O+dFjLjJ8N/Wzycxnd6SsViy7qkHLB2Zbevzs
Frm6mcakiYlSFeaYaREac/pNQJ8B7TL/bO+sbpBte3TIvwDs99V6Ihz7wtr7PVq6pMJMVVMGTkdv
zz3mENSrXPf7o3avB3utGrFoe5nGy9SSjMc5is09p4PELZtEp1fjh6awLQWl5pBbv+02diQ/EisT
enCqJ//lTslzIuIpuBACabc017zJ4R8tv5s1U8j0SjchMNY69Vf2VTirma8+sPzOjz8TPJRHGOow
blKVClacz/mircjTxduGACtVFV8NZbTijvne7YAMjGLy/MOyTcjoouV6JEDG3kEAQITVfL0Iq/Q7
VXjMputX81TEiNBXpepqwD0JOup+BlaTx4ZahEIVhOw/cuBM6EMKXuotsFxLv1G3TMph9b3btoGe
J3rRz6SzkIvlvRw3B7drr4TVLbptKEA9tIa4q8NHzgsdU1yESORxmaRhX4Skm4ALk4gKk9gEn7o2
F8VruDmlfQAzbz99QWFKKyKpqnE62C7LfGELzzJ+ZVwFRX5JvuGOu6JB8OnlxnVNx2DNBVx01GTE
h8/Ax30/Anu6Qer8JaX2UkAecDEn49racqGQrm4NANpSpcu0f5MmuEuJClYHAacDN2WQUspwzG4D
U+ZRODtqj8yGZkOJl8BagqC77UZJD4vH9axqAqTyWVeBryPtTiA7OuYMgfTdT04vh9qkhbrSo/BR
4n+bF4LbceJrJ/6VlvAe1XC6SnED7dff7WBWU1eN1H2kJEvfRvZ8CpCd0TXJbWigXaILRAP1Eiyv
YjgOVA5m8ZuYEvIIxUfBSZJg4/+IJL/wcjde0Cu6w0pEVdBbeGvjRGfhVi0wL/lXoudebYsxqNnt
yGc60t0fJjwp22754i1qUQmBwETRV19CKo+OF2224t4TWcz8NHB6t+zkxIpc3dQiT/7YozNpGDUm
oymXjEB5gHEkinTBISsyIMfV2zDJKc0NKGhUVMwyuYXAZ7nxPl7TikSaT2bnX5rbGrRV7yzxpVWf
EZg+kLbqVP1sF39pxa++tsnzuL6c8ucY4HGfQA1yhYvZxy4oxyex2Vi640jdBxtDUx9a9FpywTQo
kRLLPnvXRpoxp+tV3o0QYxzqwX9b+ITRjDqVS8nAOCPC1szrT9dTYqWVx5lQRGM5ppxJ1zUW2ZMa
F6al3+Z7bvNwTVpw1aOeD1hZ5QdbzTz+rJslpGl2vNbRQ02GaVdPTJrD8KqGZI38WC+FHnnYCuVb
tfZajxazrdU6OHhaWeV/VlYcHfQQQsGRItH7xJp0UoqNSdVFHTbyWXRTNb5jiPdxycze4wr/Mudu
WhWZJYuHwdGulszRuUnnjZzzdOC9AF9GouCXJ8MueO6h1jbYZBlqMDr3YU6mN4SJLZOVhjVrv/ng
eNf+G79tDJkVP+z6jW9uyeDFacrTpoAcbpngyo+0FLxw9dUEeDmkIedpg1k06HUl9nYeSr/HZiuw
Z7Y5B2mXP0gcOR8HKFQXrSagwb7FmF6USMXrpcsf3ElCkCD/9DqKBxo06eSRyzrUZp1fmyANMp2k
uHtH9V9SqmDgAcGMectCFuodxL2FBt6aUpSsEkSYJ/iX/x8Z8vX5pXBJH6J5e8E6VLv2D4T7WnxI
nF6l+z8aB5/WnnBX8rtrxUeyrDBBGWE4TVo4VKHlPWqfhOqKmWDih1yVrW1gSEwMje7/2BTqQuAE
fRJP8MxKct9FeKUcTnJ8bS8kt3bYsYKGgIQ/Ft3I0/SXYoMutO3vYhmfLqk4mtpFdBu/Or9bkNUY
bs9708aJ/X7tDLtNoT2yOfoF28cGlT1ihE/c7ZMH/lvSEUfOpDgHPcMBVoD/lUrwlddZBSRHqtlU
C57fVjr8Be/Z0ykdtsAorZlGIp2MRN1St90ZSM3m7cDsm52YP+X7zsgw8+6USprkYkI9JrAtn0XW
HfI1zoIuFhr4tbK7dNyc+/E6SAYjzLL1zt4PH4IiEcVwmC9uOQFxZ+TScTj1o4M5uphuM6KRoLNz
RO702qpzUKqV7ViIM04zTOfNXWgz0brWLx+oZv4GEPY+3VbymO1EmZ6xf4qC6joAa33bComKTtE3
045weKRbF+dzzHdZe23rBytwP6xfk6Kg0Egr83LwrgbeJMxehOkJ5VYxMr/Vf+eOhv3Ecdy0CjrO
qDLGokh8gvZy/olyeFox6di3h5SImm7zVb6XkEqRowG6SihpE9i116mpZqHpIwUEQjhHqK7YtJO3
h79OkVG1xzdzxGKZvzHAAXQF8qjBW2h8flmoJJdsTG7T2QkIZuGcqfW1uJxWmHETG+hgqCDCncVJ
Pd72iVDwV2z22IVDHnMOkFLMublCRt+AtkWhCeq9y2nE7HG29e5wvJqQMOxOPWr6hltB6mJ4WbWr
dEGdrTng0sQ7k0/zKt4GeA3SUtx+zJzRuMyJaYgRb7iMBfAVSngAetVAtsJi3P/AYcOK5dZ0Ck6b
kt+m2gdTRWIeZ3piZUlQv7CjwHnIMJxMrfldLxzzFReDmxlc+FcQnAzmmfqaeJmXeMYlDKsTW1C4
v1OM6Zjxrn4yIzOaz3ejgItPfJ6oVQVEsS/C/CcDaUjjIprhurHzDrJVHXyNoHw27JtKWN2yvoYP
zGlfH/KzdEAzVZHtWojVAn+srhnwVYGeVKzNoqCNJ2g3adljZaZfX2H0L8IOa5smAo4Xx6ksjXG4
MAtrJMxLlk5DtBCypzHZyB11MYZN3VDw1R4n51wrrFTRlBcqbIqypkMu86wPKOhzTooGb0tJaxqr
q0nRT5Bt09yJUEB4ne6hmnFr7fu7XUNztVdQGaiahXP6XFLxSdIbk7L5dvQmrWQWtR+1eorUTiAu
FZedXbMmrMqF7C+gsGz50Q2fkbY9QlTcpOOGReSGmJVMDOlRB2g5hjwoK/6yDz/lpLJiNk7azKOZ
g4jC+oO02lZlswXsjMGoaBgemiUCuLfVaqaqGsKKIFot8t+03ij5mxqa9Hnqe1L+V1Z5FeV8bBt7
3Kk5TX7UsJs1jSLpbFET5Vi93Cm5pmv7Xb17Y4TnmbnkDkUHvscLW/VSvYMMrcmZrEawvdV+qpth
SHmDRidAVs8gm025IVgJ46Iqzi0tmeCPXO0vfNfNUrBXvoJ9LFNiW3oAFCg6OYia/qNzZvrrzNiO
GYDlDp5xn9nYr4v0EeWDRH5Enf529ngUhKv1fLJ2kAE54dWvhTDKkcj3wHX8EMGO+JQGucWXnFNw
AIncuj86A99HuJJ4pR2KTFNqIuW5qZ3heTdT0TcOlrJXQBBgZtmz/x8ZF2Pmyiobqn4P1jmJnuM6
anl62D6M3Z/jHngoGKQQGSo7zG/3bA4R24hYnh34tbALbfNGtDf4+JkdNPqjriEO4JDz/xsBq/Bc
y/jZUwjr98woNcHt5IXrP5A4IfjUkngb6JVU/pbSNfHy28D/YeAoqG3kHly2hXtSQ7UNwblrDx8/
qiCOGwDilzEeaIAre2NHCHU2mLYEB+itleXH06t4d+v9h90Q/PTf0fD/clxTJV7tvdOoMjGIPGrF
iuf2CEm7sCQ0wd7QOhCsdCD6jfB21zX6Oxwm60fQQPwlCniH8PWj7R1Q0tBmKH6VPRYkBtmp+w0/
BctgkdbxuDNYDh/i3x4TjVUvfk/1+hiFYMV7IkqvGGweRd/xdcjgLZkufFTbVS8AT2UIMQSMxLwO
SI80Ic0Xwl42q5jcPh6kqSVlRx1yq1J23DExLChBtEVwDCml7gRP8aeEp0uxuA1hQdPrC7fuTtUZ
RKIc742fpdJu5fWt3REzPRYkPi8cyQ+w0spYigfvcVpUvEZRe4elx1/Eg1tkhi8FXcwfwS8Sv5v0
duUbMuWz8h49t739fw5JM2O+Fx490Vl/W5wTep/doBefVkPt0LPFfj5Kkhc8dyKfux/Ij+8L6e08
HvN6vNaEX70r7ipG+L5M+dD1SMWJUHiTJn79oXJLdpwKBhfBC272SjtHWc/KEeuX8XOlmyWTAJSb
XowsG6bcEMceHY3aXrUgoTzygX/fxVIL7C6A2sHYFa67OL9NVNBK/uoqeqIIbbBeUtztNfj8I+YJ
xjKlah6WeuPZL54ENItdBfiSWYIw6LRxlskp482IeW+fajHfnaLF/fbBUb2HvWJXwwbMywYTgIVZ
0B/YgUVQhyuV6Ad3870ub55zYPRaYdW3qTiELi0tKquwj8a348yqg8Q4XJbUypfM1uOu+2TD7Y+L
IULC2nDnlxAwP2JcJ7hZ+FH7291K0bdBa4Smr8fKlFibasN3sDaxmDKrv9jIs15j+P0aLCRPCIAL
8QK+PcgAvnmjg11i/YvYAqZx4FRo/uYKIUQNHrNsE65rOWLElXYSP9mJyGQoBPiL3EJt4I9Brffc
pjeMBP2Y3KSs0LGA/DVD4e6esvpH8GryDzLaR0+3zjIIWMsOGvUm1VgqyVLeVOzRrZp+HA6Daota
S9iQH+rcI9G+9inNsngF+kADH0wmaZXwvvdYNwvKlOUWPLVWqZwEbXnttYtn9JGLA6e6q5IXFTgQ
le4UTThmis1ND9zEsHqAtyqGiwqaXFk9fl2BDOA8pe4r2G5UBiAN/EVzR4cBuB8s/e5QLUd94fuy
7QCY2ilLj9eYtU613TSuFM6zYFJoj5/CTztRti3N4qgTn35j1NOGZICOHebtAQNhpVdp4cI9c06o
W6CNFuFq90/vyNeksgvjmA30xBi/4OwLkLVN8NPtHMQzDEmhoHcMlGryKZZyV2skrHxb6+5nqpKQ
cRfeIpq+OtxnB6Qn9F+KqMfS2F1Riv/1ivAsuzi4cHKQp0WyBennCoxTnZoXgcNTR2yt1nhR07lL
H0+EDk/cP5nOEs/rUdAOywYcQUjQPUMQ5fFvNXjrG+M+tYyUe1FdMBIuAteV6zfRRzIZEMdq51Ph
txzVn+d3iNrEsSsv0jEJso3h+4n3jhZ4pjq3kN49Pgl7AcjJAZWWMnwSS2FYHGeuWENGeiNVt8ET
K8syA7eXD0aAfET5bUMANFAXFffmjY8/Umj+WWfBp1kFcdOjqSSZyW+VtAuo000/m6wExLYKv7bb
KlzN+WmgkoeFEZ7mLxO9V1rj9NSF+W85h+9UNo1tGpQEtdhsdp9KsVUtYlKC5iMtVCOdlWEdycVA
5+nVFd25ZnPDBT29OEy59olh22waNe4bTT9Qprqi5/osVhpmVJ8x71JauG5Fs3n6A9c5Zvqfcoal
kOt3quMyc+tWJGD3rKga0ckgxCGxpbz/je4tRdsPXjW/WvxdZrwxDvp05enQ36ooy+nttG+a7iL+
WviPzKJU98/TwWtcFlSPb21enpgc2/Vm7dBxwkjjjoEq1FC2e0yp4y24Y3yzn0qvcX5b9OkHDRRt
LP8DRWVNfeyTB2U0qrkUNs4zwkKXliLZb/wCr7OXiSwR2BrzXmdHfR6dxy9W9sIGhHPRMpHIOf7Y
PbI0yBabLAXiPeeaGkPuoOPdnlfG2i1YwrRhADbfM32AWjIzmaQXniPrbEeSocQ1OPrnsm61IKZR
v2968ppzqnu/Pforlg0vSu1lipLLjjoUYVdwv8usGd0Xqv+kx1pHEUjYXxYGVQoepGxI7QSXcKSY
SzJb+YRUk2Cie6oxlzpMWeVvqNWYBT0dA7H+HdOMR3mCE1RACB9HXE5P9EqO9XuHwEmjgySHH4jS
hfaDEIS7ZP8GKwJnOD/5SsidCO2K40HqwG1+VlllhwEmEC2HRaeZ4Zosv8ixpSf+0paFAZfIPKmm
IAsPu+nnFE0QhE8VhsMxZsyINJVox4td+hfhrr4wxuvM50RpI/C6ltAsvrzDOU9WxVHrAdw4nO/E
ARMDEw6E0T0QIQjcpJ/3TWUBoIP1kjF6iOsg7RIULI2fTASHhR95Q+T4tKnuVnwM5frF6oj3mW6a
vUmE6cvAinMueUg8w+BM55e+/dmY/9CZaDyGTUb9UINqCmjNnsAM657utFAFH5kqpDDJ1TQSCXoZ
p7KJinVth79nswIzkAk2MKsJck4aKXOMSELMLXzrxHgbGPRmOg8DUD0LM9xeEOVckmMd40sJeK5R
bvrfuRSh5Vy2tuU9hnA9n2RfsH6514gSXymIzxY0UwPziguuZBSoUXE596vz/hIrRc3i7zeIKciV
rwz4PE6HSF7zZLJdTIA12bhNgFg2QFQHmp0WHZrrawfKYUNnFgYw2gTIq0hbHVYSVPZP7zCYdlRs
lwtDI85qZ3Xyx38+C2PlRx/hBHBNqHttYnRq5S+UhncGUZWRdRSjf8RYcmWS16lAhR7DJCXCOFaf
ckoIej0teYe8qfIA13MxLk9uvs7OywxhEYYwLFn4kj27my9NM4YjhJWge9khQECEzdkIB7AVAOcK
hqo4Fvxi+tlNQFKeryCEgHfBFlph95Ddr5zo+X1Mw9g2CJ1Cou+l54XS8xs9Hb+Wjh0r/FXNjZFT
VtrjhY6k9/sUDTJgGGIUynGt21h/t6Ll4GGTY6+XcGd/O3RArke6Vb2QDCKld52yk/W+Mpvp1j5F
uqW7imqHH0+/4tN+yVXukSCh/SxsEjed+DeVDmf8QPdhtweP7JmPq+ZLzpmQ8AjA4EYOsStPr4LT
JEPMVjendKWA3k8FUR2JlOX63MOfOJIG8RPQkp3jYto2HoY5/BwkUVJs6zlGJOnHPaPYhR6nnIv8
wEi+uNBkaQ+1QZzA5wdyDRMoqi/vbR8fpWmpSM3hmJqoQddDrHwg51aW2debKIPX7SCwBW6n0ewD
rPUrhz+qVm8EWpzLaGcvWOrJDGSwP0IoWfFxKrBB2lnxNgyqmHexszdtikq/NuY4HIIa9s8Sap9M
icbIuky+etdW5IhqWcA1lWp6ouzhQXcJp+f6MZiVpAmZ1KxKniqqZxfQYRiE9zvfIzRCQ3UEHHtM
WhAXg7yXkffLD5vH7iM8/j04T5JJNWtRwtSn4UAMsvmVSvkuXukEQh5uboR+mrTQHEEJnavwJMF9
xIXntMhhSEIiz1behRp/ndudncwW5dhfpvHvJhi/w+M+K4yYnDV/Y9OKMI+CPCK3aSZQA52yU4+9
CzOniRDIMxkadF0bKooux1cAPVevLd1GIdlX7VpK3H2AqSul7ZHkTkwOZB2qqyDIKEQpgYp2RMXu
N1pZTgVZzcKbHbtIU/rsh24Oqi7QhH+Nc/6bPDG7gjBk7Nlx2AMYH+qa/CvYb8BB43jiPUUcWjba
Bto6X4Asfse94OE5KTwMKTbsHzDee57iF3kONuOvFGiIFm9KlTz0MNNrlT/H4N6ydZpowttRlnlD
7GHA2WOKmr1046PXcfJiKuZPemwTvN0yMgl/WOnkvPzuKvfrNvnxWFVx62aS3Y7EJb4EVaC0Hi8W
eWFI0WhrcsAo8lYn9e4pwv6VGFt1WqNIhQAGSeDl2BRSaQn+/AnPyJFI1S31mmjQLwmaAv3cz4MJ
UCxcC7BW6Xk/7E5vK/oidbMORq/lByuWswuXj/Jhxek8jo0V5ZZXPKbDr/jGynEEjSUwU3FhyIzV
IovI7HW6GZRoYDk2TD4N4GgtcBTvh7KiH4PfonCFpw3ZMfQej0AXykE2f1oY/Zk+/+ETjaUqJmOF
WX8TEqBm27k8pmKl/aaT0UaEDbLxUQ3t1iiFmYbO3zQuuQCcQH0eGHwja1+aCgpzPllbLPlRF4w8
UYufa1pvZwad+pvZBHIn0V37M2A1anFxY8RlpQzbV6mJLCMpogHg5zaQDPOPdyZK1oZCaNzOf23s
vBrhsZJeOfTUF4f+qDHGrJI7HpT8yq+kvbprPvH5UZyIy5dJGAq1wtf4H2Nhba5J0dR0zhan7AKG
KJpKI4nLLNgPAsZH3j3Gt/45gbn5liH5PLe749Yx5kWohZeNKN3PLVl1Y/vROu1+dvw+i3ZtJ82j
BPcdFR82akMynD0r96r8OoZG3wuCpEKKjE7BenQICV2XOYAb124aOwQwdNF2Xa0ENW/8PgicSI4g
b/UGYR622HpusKaUArxXajxH7HD3n0jOMp2N2+fyGQDgg3ihQ/7/aZGodaQwXHszPfX01SBM85C3
l4kiufnhqdyqS5Rh/pANB8mseGJtRCs2c7hvvd46lC1jb/9Sq+/9tTrYiP/eEdGThOYnkxzKj3cg
YAlN+47PZ2ywW79GyuRVs0ngm1O+Rws/ByVdVwnaNkoOTmTXpr6AdMIRKlOta2FEh5D6M6rZ1AaV
5sFZplHYIK67p81hQ+Hj1bN5ScQMIifzhxcShkoPVmAbcp0oKtOovTE1AdcURntXLlfNnLZeORMt
iLSQMCkUhL2+jzwocNkmR/cCUriCBmfDQV4ZjBhNPbczsWiZPPqrda43mP9QlIAFniV+WETTutwI
qnsocWS8o3LaOrD9t5Xn5GH8TZQ5L+m//Jkvij+u5ZVsihewYgyDUL5kx8e1Y1zBDyi6PJaCaEJY
kKyYDg+nqwRBx+WnkWYJbGgValZMSjka19T+F0eqNUls3Wab4KWmGysvDjgt0NlWXT0E+eDR6o54
iU/NQozCHzkOnXrDSo1gLifac3EJTHHUZrL08broYGTRYIxSxwlJj6nxTjvIqsVrajJ+8VqJSD9A
2A7vrL7aBREmSaa2r/mUsI8aJG7FDpqEJkdaTHW/gdVuVrKF6EEyxub6QPct7Ooklwa7gsidgiTl
CO8wn1Nk2RNHRNMNZzC9bUVoXfdbs1c06tjmZtyiuM1DIhS9yWu2A956RisDaD3pyDz77Qgjsc0X
7IUZ9eaBO+LgEPxRXwLph1tM9ME2WaMgIV26ERU9MVG6wxqsYs1t99eycya+hQPhgc0XPf9f7ywm
us1lUnKwOPi2Nx+7WcXOHzYKTs416xA61Wf31oNN6sWG+5OzrQ7U+25jZcoe1mnfsPNfD8tAxSEE
yriN61VeNbYQrre+qOhl8cnrO4+RWOAYaLSh/dKsJxHoWAVlCG4wTxL/sFZPgeaBOnIebRkQfL0O
iI7SriZm7nU4FQFPQu1SwQKvnvqVu2WA96czdNHr85CJnjc5MT8946PaAdRBeN6V54cljqOZFhen
yXoLWMC+ezXg6HjRjwLKgU2NsafSwcAC0z+JGMvQ0yp1Wm1CzULcgXAENXvJH5sVQW+Ec1Jo4lIM
8wlb5NPbDlnrmytf2r39CAhogOiJ863xgq37ENJWgGBZ6URtnROlh6gszSDXPwjQWzQvTMkLZahC
tb386VvCN8Cf9xa0127C9P0NKZBDkjoNfHHZjOhtKIg9lrh+jZvIEYvh/gNEgf8HPUvC+cDfmkDS
hnYNFz4ZDRUyVgi3HURuTgIdETuABGbZo7jGSPq7lKWjXBmzTPTbLPGJ7TVs5A5NyWsuMkjOGQ+c
OS9hq4VJnB91JP7Z6//yoBmwwSNyA8NgGWdX4TVGPoItNB8C5xa6bt2nBzD78LLTwb1AhGO6aJGM
hHEqembhaq8G3jy28SHKqttPxdZxJIvsKzPr0Px6r2ol8GgYvh8QllRffrSwFj5CD5X2I1ARjMI9
yFuqMbrwmZOKngqZcZop43eB3CBIqxF0kCkBpKN1YsExfdhmkBAEKpoOKZEOUm11C5MULsre0mti
PuqKoonWVQxfIznUoGo/f5/3jjHbBSdh9PtEZUz1mzxvd9Xtofxbtwb3QiMLLj7MQ9mOhTAtIdK1
0e0FeVkPC1VQ5WCbwqGtFZ1d44C8ZLgcq0Ja89/4Rqmw7SWA1/RWd8rJzMo/PxBiot/mZeI3VbrS
HF0IN6WideBlJ248NBZ5qlCmvdoASFmwbWi03z7QU/d892zp7/5yYT2BaIM2jj7acxTaiNzRzZn9
xaY79NWY8BH2Q1oqBAcKnvmk9zLgLbtXfOv27giTwKPj1AB7uFZclm/6YqUqUqLElmCYfi6lDCUY
kEIgvqpyKF1e0TqTEvi3sOXJU7Q0SWmiL1GFy7yCH8QVXIvOU0nx9jawU8P32DwRIvAM3Vf18tdB
96di++9FRdlXN9U12dCmXPdgw7nfrzX4G7wjSUeFI6CgeXmuIxJQiyl2j0c0xZuj0mjOOYDWQZNw
KKSRsHnDy5ea4EcumawZE9rpdm/Y3zHdOyG6e5oPdLOKRyRfnPSzL5CTB2cl9DW3dDSlyeWmQhbL
DxurY4QM6flMeYVhrIZS7yVJ/61P92dOC3zymzX7LT5MXixzwJXFrlEqFnyIUUgD+WKMpoXP7w0x
bGrxGlYPp942qDVl8qzzPFz/JuTAG0I4TbgPwN6eguMiVrh2wgNfX3AvE/3UP6p3/Ua/D7mmLml2
9tMUXjDH3bpR1SrfGK7RxerxVpBNzUkx80ahfDduGlbQq0/1YSRdjt0wq0neEOvZyD5IQoMTHGTs
T7Qsh46C2aVC+uUtP+pyKLcfVhfK9QZLB9MN3H2wnoNt5izqjmRaAnGqJjOu2mZGinUpwyLQy2mg
xo7UekCWFxrSC52B8B14FtYxbykluafaZ416ViWw0Fwo+OL/HCDEH5QMT/NKwYirEESGjKBaXU+b
35JGpq/1jSd5CsazGRrum5xrwWJlwZIz3xpPYqZTFwYY0xXw493+zGv5iAjUVSeUevGcQkwqYz2f
TtMg0JzUW5P0QDGZALqHyIuPZfQ4RMjhDZ7OsYBeU/LM3ac+g8x2c49NYsuUiTsmAr3im3bLsSTG
sCKY0c6tRnJEvzK8i6/lTqMM1BCE0pk+xNEo/nAc8Frh8PECT177hvIeT09g8gCwn15d6cVNbZlh
R0xHeUFs6t6tPBaco0euBarqWKe3y4jeF/lyHDRmaDmN51ijdzTGPYfsZS8cZE6njjgWpIvHAQh6
AS4XXrUKfD61V2mmBvOq+5SYQ7zvUyXYE41MXMRKVXwhuC4y4E9YWjwYDGiOXQyFU/P+SeC+/Es0
JcRxR1W1M2kVJ2FXWcZrpqMS34lANENP1H0nrWRkUNH8X/y5OhCQI2mp2yEn9Xc4XXrFca3AchdB
CvSeR+YtpGJZsc/A7JVUnHU6FrXSonkhq1vlTaAMALY4tPz1h5VEmCaN61P+Y6UhYg0AA4outIne
JJNs4m3KRCpGwhySTAYu/bIyz3gZe2i9RExM/eFtTqA1Y01Yz+1u2wo/RXrKKzOLMdB4YCqtHRwz
cEoEoW/xhcCPoWTnjOAlmqGkVeLWYllR7/bLFcH1nRgGDpjB8QrrVcDCKbKoFyZQIXNk5kfBP++g
yd59/aLoRzaKf0aXiGXKQbjIUd1ZcgqkIxPeuI2Oc6aCWP+KMJc6CBkeKQPtUkvre8fbFlR3NMsm
Rzci2g4XGScLrn1y4GfixcVTO2ok2JUl3zJyDWcL04fFL9k7hMYcN0tZ64DeSMce5qYmOQ0eCujL
HCuZeJsSKn2NFU/M4VMCNlDH0nMgWrAnZ7u0NMLU1sky8GSyjmdMOKuEYcaXAFjYJQj4jiVYwi1g
rBjgpXhd5KH0qPSx0e+4lPTWm/aXAkq1tRNYiu0CayTgGy6cz59iCWpYBcLMtz3S6nHcItO3l6+P
fje0mhirzhPPunzVG1Az8bKNCDHbhoVna3gN3DktkoMQSEjC8veqleAXSL0qI9OKNA4upDOacy/0
usp619ye0Kwwqsts7/OyZrOSHJmq7f4HPuWtxsPocLG32tztBKH5fQY//+84tasHF6nZVCdqdleb
AdeMxZo22Y6FhjuG8JZG3YTMWLgrryaEC8r69s+a4Lwqs9G9qEzfE8dahMwMwj252VS47+v7shIs
jiGyr0FuNkm1pwXOt5XyZX8KRrIKgGEhkaFKniOrSjsWKKnHkQ3LS8eCHL6DoPbCQE9D7oBPXy1K
cMyBbeeEXQqH/olDOUeqLrVjlOdvN6Y16+/w2OkoYk45FhJjKgQluVItIKmtdn6ub4636kCYLVvB
yI1D9Kagn/Csl08OUElxWfPDfPIHRwPl5KF2nafzhblTB7dI34WfCHBDynoOIcAvzMjvDdss3Aoc
xPECSmkzd4auJq0kMgs9k2ZoDMXvFhrpv3Ysn2B138c5EOB8iyJQuGZOuSs4Cf2uZ2uiTBwRmJE4
RJCQriQcStm8blsGuLFeAqUSuakUNW8FKY0BU8ZhzM1E9IV8J6+Rd+EQsbGbGcJGZPfCt4dtrKV+
IOzmfsLMWrSDf+PncmhztX8dzu4vqG6bHtYPVgVLQ4k+Os1mMcYbF0CKRwp91y8249g2y64EPYRb
VcaTrjF691aqILaeSFT8KqPHVVndzIYSRer8XyM6VNjijWgBATbhaISLOfDHvWMUhjNvZ/3ILRBY
Y0mpereYPtwpDpzLAh1ZHUBw7DTjMe814FTRq62Efwdf8+PSLboAGIjIvzAzfqKtwTtbF+g5GHk4
A4uJKfkLoz0aTlx2dau7kujipFLiAtEiOsn6JdYs5zzCn4QIW3lgUJdnAQGTFCefIiWqqfkKhuQM
mZKx8Nr1jXenXBE43IsMuSPonYFoZ/lFsoX43FZDyCOpLR2qkSgrhihBly8aBChX9jxerrC0xHTP
+OJffR1qa1ZXcjuGLZT4LuBHWuAz01eJ6EpP7ZviSIqd90AvSuIg8XTUDqKQVegU4XgbgkFGlwXV
wmsWb4UFCRtIOwoZjR6PIJuaCMXjeIEAlhWQ+6Mu+pymSN3Z7rdHxWbtU45rCabeJaL3FbVFiNHG
871mDskutwLBKnmqe+nvD7W9IF1cz2f94xCyQJ58rB4qSyKzePIv0Jn/TfRxkF3kbUXTEMEDcklw
d6nZLAt1PnjTzE9PL6FEz2WSvsmY0zDQkZV7/IfV39TQz0t+JcJAxXxDZ6AYoufZgIciPjJy51Ee
QSQEIxLAeirEDUtCTNH1D/JABh88p1x8NQvWN9UXEFsxSYYF4H6NkgDql04GJ7Si3f/EkdZbgBtY
IwkCVVwYiVnaf7D6/Y7FlOt7iWmFAX1pyuVJMs5yXU/fS8MhuPn+6bVvc6/Lq5iSFBQ9h9h54lz3
SF/htu/phhkg5BUK7//J/Git3Br6YCxEB6HxXh7XC08NfQkmJ2TV+tf9YxSY752cE1rhVJOTqrKW
pKKRuMJgX2mdgfnx034cw3A7GLKJUapWx/EfyhAJwJJG1wBDhEPIfCQGaL8xAUjjlmyhAZzZLPH5
p/vXroIPr1cWLj8H67KQbzU43ypdTO5+heGmvvNdDc4ZjwH9rOlTVO4sQRnF3vAwzGNtLZSVFMWc
5e95C1W+c4/+Ym4tLNcTv4TShZgHEErsW5vy6shazRpMXsPFEKwUhKklNlchOLvTDi/kZd8GaT2w
A+aRR62aj82bQzsM/ovzhN47/Vkrx6WA5QgypH70RlXYJsFcDKdrdx4kQ/JOuUihpzpehphNOz59
DGcSVixmK/wy6Bc01PyjjEAH6f2lzz98twoQNezU8V6aidyBcTDAmxKxHt09nnAZdURzV+sR7vs0
i4pw0oOQdeG1+CAlXg3wVgz5nYtZ8GZoOHzpQHx92jwnE2eLsoyfm4VllyWM9TnTRFiAqvJhcHjc
5I2CuHlAaBYYgjLy6GP62Wj21wWXgIMaomp4iQztLW2pipw/puPeYgfHSt9/cJStNuJ53t427ENt
+CNY0RuVlez78MIRKZ+pTaVYD/khslBEKdk2dPt8610XY5fCv97p5/AOBQnzhoFocAULXyYY9yCE
BjZdJZCW99FNLn0GGppeFVZxJOXNsrFKPq8G5mCJoBRI9vPyfb1C+V/+A0GB9xKfnBD1bC0jvc7n
N0m2rxeSrUIAthvRqiQZTSRO59U47EW8zWww4Y5vYSKtOxx9OdkxiUgHGVe2ZExwbAyEeG3LINT2
XGvZcbPLpU6Vk9rEWx7uPWI5oRlfP3aLNtOXYmcf9vMksWz2fVhBVdmTClQVMVjeAVgU5a9erPX0
ZwM9oWS2l1NhT1Zik2Xn/ITIlOWY9y0O1o4C9KNw5VfmaA6MOHox5ZyxvzvrIlzrhjcCiTPIjXYe
UgCz6dB8AEf4muURewSLg42LnEfUz5fkQ414Lqz0IpPBvlVumpbKBXSRoKwB75Tz419vgIfWOJAN
xoHcpdp/00/aYBLc1Gs/9WNMaw3I+FrvcIr92KMT4nrFhNVzfBCIM80a12ItdEAteEqFMJb7Km5F
OSluBwYlU1j5t/oyj2Nhhm8RXuzDNQ53I6rMyy+fBHiXbkZDLASSsyXrFIiLOugyGf8Iu71HEyDp
BvXc2z1ZfR6EPeLZpRJkx5D0DXrcRHDpywbjVWt1fgoOGe0PlxEuFsqm1UnZXcIZZBfVaKuObMUj
FQ1PlqFFhsslAq0o5G26ioH2r0XXj171l51cVvsNX1bgOP6OFWFaPjy6nHpW4p/JpOJKkGB6EVtE
ACJKskwR29PvDaJ8uGV412hmJWB4au4DTWgc+Mi0EZ3qRcMaP73b70/tLPDtqcmTysuG1Y3HWdrt
/xHjf830BVzYKYepz7nqtXYoDwNQ2qkoiwHH23EaSmsGOr6Qs6lSoVKt9fANYH6ruyIJagnIJbie
TBOVRVrgurSq6Kni1BHAAVbWhRAHb/P7Ilvpf3DRue680TQkkBTxonfEHJpHRu26Bti1gV1UCJF3
Q50y5Yzmdy9xfkS1jTNVFkCJJmKpXu6DhKtEks6LWF8tCKcr5OeAshy8djB0zXFRVUXv8Q0N7xlF
meDuipgAdwmE/mjO06nKFPEsVrV7Ry2tPGH8EooWaguSrW6/YA7uAFwu7R4WG5CDtCNYXydu/LL+
EAx4HY6BgBMQ2EV5f2NVg4kdcKC13Lm9+OnAeGzAsJ2O3AE+epJDNZLsQIduZqvRB7ssoUZi4TQa
W+8A9Mr7qntvzgHaxaYlOUFQjkIgR6VxM0R6ZxketJiTgY613mglXI4nXh7XDRFbtLxQ5IOXH0/i
dNZgdD6TJd6DwyjH9eAPWrKy/a6tf0MthQ1xiZL16m98JXNQUv/hW+/BWiO7CulcOgfSJhlIqPSY
d//7AcVewbL1yGNyV2C+jqze2TXLxP1vVrHj8TMrLHqZY1qngTE6MgbXlyX8uZ9tT++NtziSbN3P
Lu8i+ktsZfygiWVhNHrzYobRjzKlGU49SgRqGuAXn5kkxDF1lI1lHj7uffLtrcuCaCvbzVMpTQF6
ZdfvkCkOXUXX1X4qRVIKnmMa9imO+JOHOdisn2gTLvyQA+idqSYu3gYj/IQw872W/NPZyiGmPsiP
ecYWZ4u3gWmVtLSKdT0f0fJTIqNvRx1G3jpi4b6CTCl23cN6++8LTHiUwyYsHyvotI1IDK/IO102
BxtNuuysP8VGoqUX9J+7Zd+mP+6M+qTEhs+Zj6cZ+sQtFcdqmBwdiAojlZcWDXb6Xpk9UidCch40
2CTFbaxFfi0AeGGKxGo3EEUP6R4cjmexzjKB4l327+L4xYuKj32unhfz/c6SYdvp8uL0GZkjXuxk
zPTt2pfSTUil6pfiPovZ+9WgL4Cc4cmZrWxaJTJ7SD2XnkLKtFm34IVHwZSi4eEhmFcPoJmfGvzm
A1jmP8cDkRtrW1GjsjSjI9bHuqia9Q2KzpRTz0Kz9zQIIbVMFGeWNP7T2H3kKY9crCVKuqCOZfkL
FE3ahWAt4g26YJInDeTf9LGtpYrUI/X07qsqiqHD+QmRs6tiVrgzut3Bp5JT8EEwJp7ZAfnawXlW
HgjHAWJJadakz7TEobVSk5G0mmjv581BeefCooez5QoIRJ5Jb012KsVA4KKEG5pAibtRd+cNuw1O
g5PM0u0fVcItT9mXKbaOnGEsjuIm9n9mpEXkadzo5jFPJ8I5zXtaDQgWUGSJTcVN44vYILBwU3Ai
HSzz3wWNjcSCq9etKUIcpGRq7AsUvA3a2HVDIXK266SwszMKsghObEOlZhXYxJxiiFNtPwZi0Dc3
zSRkvWwdLAYEUzwIs3YrQzF7WsNhEHJppb6MVDoY0j29ey6rlpieybG8hI7LEohVLM+NftPntLOz
KVky0f3zb5bX3RejyXjJKuzWIps6fp30fzhYoSxg2oBHLRxH8vMd08Pz7tl/LfcUgTt6e83Vh47i
eajGSp+F+6JFmj+askf9ZIq1xiiU8ftxSlsN6miMZKBPAqFgqpaLuZrSNm9L5G+E7odOrlxwBwq2
4DewfAZh7C3rxX0Sr3IfwLipDRrl1nJ8s0c/lXqBa5REruvkDa0gciVwWVZOEgz6dW2Lv6gX/+Jr
WEvawrvoSAH1JE0KenJGUwQVIbW4rTawtY06uqNjCZqfn/zoH9ZFgtUEiE674bLP8vnZo7M7Cygs
xW8Iu6m9m2etjQnmjqUN/izSlWHc9ihSrUUraHKuNiHDDXROePmei+PRiyOW72RgLo/+7vZO+V3A
tig75t4hD2JADiuS0cvgcg4sH4iLWLDL6x5t+Pa6RYgVgH8eAf/qoxOUUwn4a4iE+KO3nA4JbBkb
cuFkK7x0Pm4NNmgS4myVkdHT8dVgSCXenkWGxtzbvdqbDm1Y8ygTNVQyXMmgKoo5HONW14B9beOK
C9DOooHURs8WhL9k2qmgkkg0End0rThxL0dtrY/L5qyGnUrnf9ylKMyXRzDn4KShCQo8uAXvWR5J
3kH14f+jl59Ud8shDI9e61/3+WxgnaoxSCugOCutW28NFc5xNhjqI0YkykjM/yrCwV5OGZ7llTSY
qn4BZzYlKkSBbg7BPiVMAoi3Kx8XLfSdGuJ2XiHsoST/4rmuoxddHBQmBU+PJmzdE1FrdNFDSN9d
CevogOAVnZxsN5Sqe5ApCFPLK9Q8HqODvGTib6+agljha8bCXIHK7sYKIUc1T2TBT8JZ2DxYa9mM
ldvFokWA+p3jwNlHmG9aDAYZiZ+sm9+wTZW8wGAopndcPuatEsiFC/+Ot18P3k2Ce/CVcL/hs/0S
az6p48YiKW0ZRfp7D4s913U/FhuwGOVXci/pNqPYPSqHKsV+lW8TwoHSlpRPSwUPycEisqhweT9o
40CMSxgLECxBaU/OCopbuGyWviOCjTSPsmp3hrdba1EyoQgttXPkrcW4lyhz5qlOVJQq9QK7cehx
JZsUsNqpQqCs6cCWHs12J40Z4K7PvGGqdRv2BM5DFw+7zarcEimG5jFJBhp+nbTTqQq2Z1wM3DpV
m/o2l/Xnnqv/V0fBbN0862Frp66pdn3OGW3y7yr0NxFPpRRBT1fMNjJNS12SX1m94Ns+sQMUnD74
VxWm/2Vc4T8pyGb9aDI8FjrBrgyOHlr/Wk1DDpkIrOyrVm7d/zLoXWjPiFX4ogFbLg2UvQwNzLoV
SaOUGx4y6xEl+n7ApEJ7xzhdqaDYr84xAgISSdK6N828s86j4cP+Xne29Uf1nBF6z1C8rTmnXcTX
32xTQxtpYT9qvf5bfZ3D1bsmMVSp5gM6TYwH0Lq6VaU8bnWEetRuzyxMz2csNZ3tM5+MUT2tw++E
3Ddq5XtAlbeuXHntrdsI8oh7NhTPhZqsw36NxS2cDyRSMdH3bXz3EHJcNGJ9kIogcJzTQBQkqNby
o1XuJZ6zd6bXBL3zPKWEdy6eAFRKMhi3rG/bE5M0O2+wyxwMFPzd+3D7Rjk/40fdQTmsTI67d0xL
4yFI+zCo/KKV/ODV12cFQjrLpE0BQPoE9ZIrCWjnOoEf0OSAg0iGN3JtSksno65wwPe4O1mXQqTv
uq8FYjHzCK4q8vR6MNdN5q3Ap7ptPI9bDyoarHKFJdFik6jGBZneGqRWAjYUlunYR8DjtZzvvtkz
t9ES/GMpc/ZO0qyEyek3EqxpcvtyoOgmqXQd+qFDz+o9bIV6U6VuwHI01KUXSL5tRveHz3aV+scV
CdJcOtjOC+lXzeryT/sM55QdzgvzJbLcigF1LfXyxJOvaRm8MxER51uubhOKdO1JItAjlyVSBT5w
fRrZnANc1v+5hHs9QrETzVo7Kd2bYvTI92MI27fkVZ6F19ojCs7LkA1ZnOzokYKPHce0Ga/jrnHk
e1k//LW2NU3iwuluoPNbPrKQfV1mw36k9P4n0I4u5m2bcG3uOvXKTbvZ7bT8kIP4DHai6ShVAx/h
uMILwPY4VMCp0ltwbGSwJHVfUvsNmvsj6+dlzGLcsxCAm1sKAb3pP8I3jDNbb0flkTMPbm8DHetL
EQZUWHXAFa4VOgD13j6PSkPTccYb6q3M0z4Ep/96k6XRfwqwLXSHyrbGhibciQwIHzwNnhgPmaRe
iVQh3HuAKffzjgTZqGHaHGHQ9BL5zE5N2SOvObfnxXOuOagNt83Grne0EmQ2VQdFsHmeBRK0eHr2
M9yEyMaFDcDLAZJajPeizwZ2JJ/2aUggKPAG8TA8JER8ENdAKwJVbCgZ3rwUuXFocp880cGT0cvy
ahYzHbXDa63MPZ8w68kIlSef06gChwO4z13/pfjraqSSzhpQYuoAw7tScHnQVFauZflv08DJvx+i
w0+DCW7LMLYUYgYOMqQ/YdVzATqBdFc4p/nh2vpjLfmrgXy2BBRNsQS6BYp4xkdvYYMRegsTrSXd
BdI1eTeQwz5mZcQ/hwVYdBYWqjTvsNRtSVol+fitITniHLaOdL64lA3inieHmR4ujprAeeLAjOjq
F5Ul3IvCBBWF9AV6ZMb+CK1s/sYPj3TEkh6vqj/DNLL8+s+erMNyljlrBSajErQRYEPbP4wdds0M
p3lBu5zhnaKoInV2bai/ONnA5J8EYFrqV9FntzvJCjzy0lNxnvZq2vio3/pzr/Tu9qmEqJJgrQEk
PwQeuBkS+mkUM1IjPTq9/C0ZOHyBtQ181sm7i8Eudc4MN4SBskAr1lGinIrj3qa7scqc62uQxx7O
Y/PYAmqG4F+LgX7AYyWkAF30GLMQgTPGNJetq7eDFc+HTlBxxzf6+x8vUQwqIQ+4MmJEVeJXKB6j
FZj8HefS+BhAgbFoNzzkgo9uX569EZpo1kZLfk9BbXT1PVtliZ8Vk0P5YOWlI5R0WzX5xy7GoPnu
riS+Rv29ZWv1duHGDvemXguoKMPp+SWZVcnddItKDDQvUwYtSn3Z1/XykMaoFX93PGgLD/uuR1nj
cytHz47+ewTsS7CD3+3X+UcinC8M3ySuac8MpRMN/6+cYx4aOOu1vDDAdsgVYcZbxMyHTNzimTAT
EG6BJ+LCs9wqtyFN/vt/Q8YtW2bwB4Nk3F2UnwfZfYMv+7MMJ0xEiHDCcQDh6yUm/YHf3KKHe8P2
rIutdRVmw3Nf36JIsHORl9i0YHpLQ/sPuBBryuuNCXvciX4XMmB3pz3rh9OQucs17j+Du4Av2n1/
ePzT/BrXNhjBIcrDHg7eLuS0388QBwKJ5emAuOdyEKmt5MR2dP7o02hF7gVB2wKWNeohZkOEcHA1
C3wE+SrTREPMe2MB5nJzf4gZ18Qfm/KrdWFHBsrZI1VsIntWfgKJnpIHoeWnuNFF9TGk0l55y2Su
dI1qNgk0jMwjqDVFkfm1Hksg+joyXbws9ruhaf8rwjQpHA+yvAKUv1M+XtRCxwtV/t/x7iHMx8nb
JUNqQAM4X9g3tHLg2Ae6TcDL1v3IRmNgBHUiVmq4+ZaoJoaSHVUQdem4TspOlMnNp8MAP2IpenBx
C/JH0wEauq2OXLnpzW9hyIz6bWC9iKlsE/nTHotHXq5jVG9EtargOYCxYRQ8DYMQ0sYS70Hli9o6
HttyQQe4THdhvyPuX75yQ2wEhTKp455Oh2rQjahFO0Xi8px5eJkNnjoo8Ve6xjgrPvqe/CGQk70c
Rbs+bpYUDix663WdyiJmIDuhUeDsOhpkTf1NhIVneZGvviT6kIsK7GPWQHM0YGodxHP9yTeMnOuz
XCIv/l/LNM3Vm9ZAA43CpQ4951LIvnos+0E1gV+tfXno5S4arNdhjRT6uPFOMeouJQT5uoPL6Voo
EmubdPv4p9qGYnGhNcpxYo4CO0sS6rWf6lTNS5Asmpe7zRhk9YcLm65KEVUxWA5R67Fpc7DAN28k
Epx/J4YaWlR9oPUeDHbaUulrPloQ6mnhevVFgq2iHqmEMYcJohl17eLJJn28eRYBLPdXCkkR0z6c
itvvdVd3kmJCGGYB+he2aFwiMhGpZPtUFAjuClJAGdHWJFxpUBQZOpqRoVPgjymsOIvf2s6AsSFo
r9S2w65avYXYBQdUgyTnl+dHn5YqBcHhjce+ObEfnabMA4C6HidFwDr/h9fXvUDgtceQGeIXv5Q7
VzXtVUOvxEHpnS8A6YLQsoFm7i70+SmM4KaiBQmtM/VWdnKJSAJAQ54AcJ7C61+EbI0ThGFVc1aV
PQlcqF2V1qZ6Y3D7n9TFrilCYSaAjM+1z7ZnZzhFFQlUPl4XUY81zyGMqxbqXBXuCrrjDavFT/wy
jgEkIjCA9hgCbmPyApP8tDCAwUnqHEyWoYLXBp7tZ8Slf3lJ0mXX1WIs5zxOl1awk51HNXW9x7u8
uSES9qGK+BMqoxO0g0fFqkn1P9a2OvQ6zMne7CVkl/LnWF7hH/BNtoj0zjxsS1c56ujco8/uugm8
O6bMXL1YE/pPcN1I8kd/UWqLbLFilZcf5UexyDDgfs8TDZJHlrBdsexCSGXrIFUYyCsphV3EP767
wpcNGBeeMas4Nq71AoTag0OK//wF2TCX8b45HO1I0hTIJ1pqPQKp3Pm1Ib0ne8nmkZF7YDcySqqi
duycHVkvmLf8TrYwsqoJpZoIjWg+N4sumXVROShuNqC4goAKixb7FnxaPz4ED0QWWQW0UmzKe6SY
4FxXq2DJPUtyylSizvCbXU1/WBpJiLv2IINO50BPpSmCSZcX1/80M1s9x6xDjODWUsa22jIkDqAg
GJFRX5tlrTJXolcYt2+tQbY5J1aqeIdsjfB69vnb9oQg9SOxbX7nReyVLLq4qiOFks3c0oDPsPmw
dUSmTaCtvXeXvE/uglWOEWlR/wYXTzdcBBy2RqkscRqWip032wBdD7Fv1QrT0PM0QUXiGRqkE2fi
TAGTndofwJPlJ4LhQvJS/tgVeMXL887noSXvnOAwTIwdT1qRcwdVguoXi3a7Gu1YgJlsC5k62b2y
6NJDXsMpuH+JIir8O2cP9fgamxS1eNtx41sxaVQMC/JxGFoYbcyrHaSynSA556mBQy10sn2VjEJK
eqnszd0Ov6bW9BUyf+rcZed12fhgYmnC7kIa3liRf5oj7KJ0uTxRgJYwT3g0ipsx4lasm8sQE9xA
F0dbVlTFwIS+o8C7OtNUjAAM/KDdWEc2Y9g9JRgswhF0uzd/B25ZTTuerokinmiVYq8mcryEN3MU
uq83K3zOFztXjXmUAIDTxDhS68w4wsAdYXSNXB9HI9mSt8Mly0W5PlvExiHN2EXjZEa3tkXGwKc1
atrY1fIZakZxqBXcodVBel8Yu3Q/Me6wevVF7YdqCdjFCoAd4i8Jjfl3PxrvMpwBWRVju9+KCGyy
kFUGHRpRJegfT66LtbMZEOfUUzr8JY45Bk7dji6b2zGYTTn5ExaTmSOKJFAplyfCsmzVW3qVTHo6
DrRYQN47M0oBMzXGjHMcQdHeoxWFPxkmwZp4SdNuL2BieZgHEYypDy+j80KvNQInvDvwlp3mYwVG
zJuIJ/r4Ho+6LPud/6MGCJLZILJn2gsFIlpgr0VLAvQk3l8gr+wnwYEILC7wQXUQWySfaDOlMN+u
DbkvxAVBbqrSA9jNM9sKE1RcGfr72JcdORSYWG/jOkAosKwYH/ZCKmuFQtsE81H8K5DMZHE7jJMb
U9bske2ORtwc7bkHtflfJjqshmu3zJI4UvTmOzz0fpIVVhyNOpvqZfGhBDdBplQQrfso3TauNAsr
jW9DkHEDrRTPnBpugP6EOa6L7jUp6l14LzhRJ7ASlV7tLjrZ90uUi3/lv/NdqCtCb6hVav2i42EX
ISXHMwhYtOhsjHA5g/hBuKGtHm4OCJHtEdKjFmCBOWxeyKXSjoDZ1YO+E3Fs811x/Zvp7DyYOU17
v2ki+KCLv3+DLW5FGnr9zUMe7ablrgA6sLncqeWuVeP09EQpYeOK5OMhael9IzK6nPOTg42nsTFP
d0LB97BaPPyUavu4YqXtwuB2UwRnuLuvN6prh1CAxLA5Wfz+7nnsDBs3cEoHo3PjiocwL2jTkOW9
CtLt5pc0VYVnVCCzU1tgqYToDwPxmyYLzMgR6gHJFwIc9KBH8F70OhgmKM0gM7DmpPufoCthyaYN
tC5rcd4nuEhzPMaN2nRZ5B/ABV7+mxoeOIAWGfEsligZHDVNPnGKkTpu0qVfEVFgQqAGEIExuGYf
HchImzuvUC+U/ZFYA+jQlOJ88lljlspGyjyauX+zJrQZRjlaCIbj6qzWUh1/EBHlvcVHNWbQw7MD
6Ffy5yNivOZdpS5+a8iFcOExfdCpP/MW+HnHZam1SsnuXZHUfiC2luSwDKA7oMTHXGfrV4c7dL44
KLtsZMwTzXD1TEQr1cgaVWKS3vXhBPq7klhswxFCvvQbOJ/0bDD1BpFagt4eBV4uFNUIbmcq/B7+
submVrTs4jtYGsaZF7BYS+Pwq2hucm9SVNGcrfrfIMhn5837y/kulVCZtRC/6EwVmkXij+JXm6jn
Doj/+rGO8RWGG2uXxJrwpX1UDZ1AgU9tvylUyNcUu7DbXcLmOq5/PpEgDR6tTuGfPjzZAEeCynuH
garS0D5g7nq4QjZbiXR3ITGbriIUsq0v58a/mk+Tk7rbvgriZnRHSdnSSl3vyFx9qXgP1aAXX5h6
Hn5E7MIVQ9mIvxTus3fi6w/Df0OqweZjhw1nHksBdoKHNg1rFR6+cwNkVyjWsAZ/m9sTBWtvApW0
1Cb6xNP0rZsNSt26WsXW5nGMm53nTCKBAD15jtSSk8RE2ieVveJoUSLbcvcg/akS2h+CV9GjIDTd
tXwjohB0qH1RJdtNU9X0OtdjxPFouQcgJWrjgL1uOrMX2c+Clp4wHXj8qk65JUSZCDKHlYm6tBrB
5oWAr3lV0pBYVFHYUg/RueBHqsmAiYw+QdnC1KYuZvvRwZMGsebnVQ48zLOLcfXtqF7jUJyqtQ1D
1NO/0tpgRHyeI8QuQDMc3i0f60VQ3v3gr58O7kA5fIAqPMumHTY3nj7blg0ags7b3Zg63cBK8DOQ
VaKmbUVT0qzrLC4x9DIouOVTC1//up3JzFYRsPrnzIshBtwtVF6wtSyFcA1fpcejGeDwt+O65wED
LdpNDFa367VKXCsOnA7pytQGcLGW9EQhxTsjovxNqU1gv/uLVRbOSSYPCKPPuf0eMAyelYdhb0vq
HGFE0ckFepjfA2YLdMv4lEX0ShLssdcVZjf3s8JuznJrX+CMtyLI52PudSsHkYqX24bl9tCYME39
uOa64+H1tKJo2/66hsznm/3NA530gsrVllADfPX0dbzvd/fvVEHLO2XB0G92zvnlzhtwZFk1862Y
MROX006TdKVamSvpE5KlbFQ7DsxqFyfalCk1t7oeQMtrLWC4oA/JRBZE0m7Z94QmgeCsIWP3AVWV
mLF48tHvmUE6ePyWV+zNZWoeByRiv87cFD6su3TL7ErGVGEOlKa+DZ6NHRy4MfKuLLTtHIAcCfs3
nsiEZ340jVk5MSFali4tjlKWpKGPt0+YyJyQ5PpryP4T3HbVDDI5ba+bbKgidjT2wTu8ogFoN0Gc
I6KCe/xFGN2Q4fCZnOojeJs3ngYp/8e0fE8ZP+k327Zl4VSorSnlUmu7sKEbIxljdGy1fFj8WSvd
qQf7XxmINE+d0xOtu4FTzwtJzhA/aFcQy2GqoVid7Ipu0o6nC6nQxeb99wA4DC/6/ty+cCn6Ywtd
oBiClBNPPkXR01vrUIUg2h9wdf8PxK91T9p26EplZ4ViOT4CpDXT6u7uu01gYaxRZlv6Z80WXRwY
FZp6X2LL9ljnB+QuHqz2qCqa9lR7pGggK1OjCuq8lp2Q6q37til46ZJE22GjNTyE1B8gqpUZHTDX
1o7ffKjTBvcF3V2XQqYtPyuTydGyCVvz0GlzgV6UyJbmWPlKAWLI245IdcIvAGWXHu+0bB98+jhV
OGklBTaBQtHw8gA4aT6o/RZUDvxiSHSK8DKgkbrOxNnOegp4Jh49OalP5gounAnx4v5zToP4+/H1
YmlbksJaXim/GQdbLYSqI0RMkS4PZZz0C5hvj10UIeOGZzwdBO4K28tZ0Y29acB2NHQNEarn3vg+
WDhp79fm1mDeBarjfh/yZ9rI6kef6NbSa/u2UjXhQ9vshUm7QadBqrKagNzSVUFFuC+w2mDrdS75
6BO5XcbPEmAfYKq6dsuoD/6gZZib8MkNaG65A7OrYz05lphYOJdo+HCKKMBxMhmbQwRezhT6HmWc
qvnkY8TNb8AQBA2lLgX1s4HizEH88b7DATIZZXaGlJ/wLkJDDMJMaufQZw6ChkFzJ8w0T9kZmTgG
T42AS2KF//MoevLHz+AaH12AdW5mZz1mHfCMoDaMB9ZLXfkL13gtm4f60jHuOheUQ2mSCL0PPt4P
6O+FKCRlvYGJn5TFyuxbROxPKS3UkgkUyFJUbI1tD985K+RoBRd8RME3F9vnYSa7mCx8ThK7JBfQ
JPWTPKHnQTuirj2iOJn2vrkWOJOExd9xHDjzzREQUTsJ9/6C3ud96LStJgZlONQBIo2O6UFBCxWp
TWUo//HLyEK/FX+cdOU/48WN07Vwh6HFmr0wZGhTyHHX369uutiI5O9bmA6LBtpe9QpBBwrpYfVi
NqGYPQ+jCoY0GRtH2tgeaJ2bmON/KzM8LNVJkAGJzJh4XWZPLUP72TLhHMMuDV3Rdi68QJ/BH3bB
BSntsNehJtd2FjX3Gey5uOOrRtFbM/+Fwhq8qJ80FfW6qUv6m+Wft7r3/NSJWUUJy5jMaetIniGz
mTtdCEToKjWiW9tBtyorlaUArqegPaxuLcqOGeTMlniVT1E5i9kQF76ilS+uXNPa/mnvszdS3TDM
rVAJmc+7EmfqKs1S7sfZp0H59v0Td09nlZbSYl11+uNPXaPVX1Owbx2JyrPFdQFsoZtRY7XsC/lg
N3SvDyS0ykxa+0tFnLYf9nOmOWWv+gWp9cRUTREYpp+xndSdyW3swxpJYilVHhR1NKMhgQiGLTsE
bskMILkaywsOD9UbEKVAMK55GVk35TQBSP7d+ymvB5jn9XTavI/eKxAUlSH9oypHDMhRUp4/7YJm
30pqG3DH7iRZgftwehP60glAKyPsupVeLVfEK05guUIbcfUJvUqpQQG5yjxmemRraxqehZvWElA+
e+qThKFnrf1z0Q5+TWjIvmQLO3kSibbXseI6Dz5sZLMebNqHBj5xEMXwccU06XeETkAlNi5MeRRD
BUAqYUpJc12K2xEIvIY5+0vipNVZCo+8oVF7WVGXwgYcGwFd0Ssb1umOr3d938Evys5pa8QCe7gB
2ssXms2+tRnG+Yka9y5ennp/JN04MUVuUAfnYbCo2yBMrCHNhyVQ+lpwrdxr8PQHhOGFoil6/mss
pnp6T+aPRIlTz1H0Fm5lj9rULatqDMYNkYvv8e7Ibt7HNbzGPe7EAu2VhdxXAD0M/y9Bur3iNFza
fPI6ocOJdOiKjv+rBBxAGJuZ6CMiOJBbxK11LoVGVXN70wFONqhrbiZMPm2SY2OT/B/I0v7GGDkr
E8Fc4ydnoEf8e/p96KlCiMUgmNEFSc/TfGiJoRYcmTt17A9mrXVmEkbd2bjHzdyECx9mA8SPMP3M
M4W4af9BYyUxLGzA7e4kaPKvejUv4TjiGTibe/Y1nt7FREKij+0n4MUhnpOwZigOkWsWZ6jK7oZh
n05YE64IB21rTN6Lzy8RYQ7Qz3qAKrLUIgmxTOb5Oq73QOOvrcb5OIfboMh1KXanVK28Q/+ATVdz
nnwLN7Q3DI5w/CMLPoTT1hjYGin8Hg48c31XfjjCVqHqaOnbhj9i7qlV62GGKJ2G00Hbh9wh821X
FXIF1jjcwUfuI1d6NTCmDyPpHp+5oiuYmTUO7f2GLPxiNLII7lgD225ybBv+5SxaSPG4ibVhVCch
TZ51/AT4A8bge7p711YE4aQj/ortQqwmwn/W/vyRE+2zaCaB9x8+rHa4y0ucWQTusfOudxV0kuEd
b2hf5ajsx5tkPwEUUlcuUae0sgtWjDmeC9oVCgXgFBPIQuaq6EK4xd1saASvIDc4kBa40S6o1CFk
2VHidrj2u1dP8wLdG0rCo1qMKXLt5b72iIK4osEhZyf/8z85ozwdxD/mEvkW4Diw5Qkxx1zlz1MN
CMmw5lBUu0JOck25OFoTbcgfI9oTupRMbmDobNQTVVzfqhRxMyrnr9wESlZQYePD6BD1DYiVxPup
s3aRSFRvBBhYg8L9o3byH2yb10O5Klrglhks7nN2o2UNqAJmttcMbJd5ZpYbxbE0F0qf6hfxenU3
rHy2FcILQMApN/V8NSBYLUHEcJTMuBtZcSqK/dHaK3BDrS9MfMWozVhfH210qYsmGwWr8Rn2Kb7d
KjsGK47CzfTwj9NDXrjeTLJKuh6k1jJhDRr5fw8XjCj7QJUhKLueh/n65GKePXV2tE+lgWdegvXX
OHtd61hjgKUgzWCx8RdjXEcpysch1DeyheZ0+Ifh8nZCuzMChZy7XZgKOn2BuT4hUIW8++hX0oZ1
e1rusypER3wrb/3NY49Go9ehiFnyVIV1GWQ5C+f+9JDL2nQ+yOWgUjsalDgwiZTYTuTz02+b4LCE
rGOLnQIhfh6DYdTh/cu+OlwlO+opudlvXrPlHhG4L+ScDmBhLBUxltS0q7CL54z0JmNq9Y0Ib/aN
MbW3OLV1ow7yBtFX5RnAWHwKjC9bFlxuA8TN+eU6bw3eQVPGQRFqqIfL1FABga2pMJn10zCtFmKU
rptOh3jaNgLb9wrHxMMqzHretsMa91yPc/u+n6oVCHc6/4Xi1dbQoAvgOamBQnSCj97hBQk9Qa+s
Lht6EuWPwGEE+vBLsxRt31ks+1ddS692cAF9sDpOv/jT+8INYxKiFn73onfx9yBnyL86+k59YUZM
jxPWD86Z0YQb/vhF6ybg6xgUE5AOEPWIDhu4Ag0U/x9wWctZDW+8asfAgD8HorYhNNk4eTcUS8V1
dPw5cugPux7XJfqKe+06jsSYfhDGvmd+l1Y+RNTAFj1geD87LmRJdv5S1f5Hi0jhF3b4xrtRt7Ci
PTDffUwvoRA3Z3ziCG5OKv1DSJ0ukB4Fk24lgnaxmZhlde9ZmcWqeEtZOLgH3sYQpb36F9wvFwSu
LTYL9qXbY24ugyp+JphI+/tBPwk6Kg7Nqr9cT0p1eZ6HdVWgGLn/aXFpN8NH6ooXecXnvovJ+/3R
wBL2WvUL9FYHcD6DiY6r3qvQKJdvxB/nyivY01N6kcBHg4bHAKKUpyy1H0pW6KL09VSRkeeI0goE
eh6b95mTKjQttdPiURJ8BCMQGTx4FHO6SsRbqlJ6QppItQwuH9i69yl04lZhsjFqicQxOvzGQsth
0Pg4TxIDeUOy+taXHr8jcGfB/KYziL+ScI6jyg1BZaPytlky70107QHTwfmhDdaBxv+swv4gdZxo
EbUJTbEztuNBHZu7HXq6I9pcbEqE6a2hjknFeH7txyYMeV0W/SBgrWxY5TjQ9b2vgHwN22RTKm4r
MWkWN7nnXCjLS8n7Nhw/Xb7srDIf4ZqoA1VJpbKipRY7l04ZS8ZDMOoBNvlbAHSjBjfBVj7HpqB7
Vi+xgN0cxr8jun6sIA3x1qaX8+c21ksRijngND/NpGnD2YRbx6jgLIg0GKJyUi4RTqWigtBAOLu7
+5fYbVRP3DhThIaLf18o9djRtSNYjnw4iYx6+0XVIw7l0le7QBMw1A7im2Ah3sXzFb206/u0KF2V
z9eFGdiQQc1UtmMsqKX1eLgq6yJKmtjNiL2Jgh5sCyG/KPiXwB4a6X2qwmKHhhkIkYGoYJlneLpX
yz2y0PJj+UTgjwMC8q0XNG2z5j7T0p7pJRIDHChvK6EertfwCBOwlhGz93A7m9SkPl+fUBcnTJYD
fViOlR3g3Yhl0G3xX5pYNdNQuFEkNZTyv/PyiFHMI97lvaltsi/cArYcxSKpgUx6AWmffOjNVPxO
06AXRpquve7mZIlEmfQA6AB1pjyoKgxmHSyVR9sNShDG4U1s2O8apiIh2QXu88uczq3ATRHRfV4Z
RAYGsxg2ZGDfjLspgJEH7rBbHFuPdSCzKpAtH/FI4I5ON43gP4yUcSzPo4zkRH4kWuHnE/5kQoEY
huwAMq3rEwAgA0NhZnAXYCpHWs6yv6hpCoyvwQuM/N3G3twdS+FFpCd/D38klkgjYRuzCohG3IOe
q+oPCadh4VkmcSkmjFu8r/7Bpw21XIXGw1eEhBtLP4v1XbMTnNlZ5edO9FUaobFwm4mbCL2raFR0
2IKucBjSNCcPjNlfZSBSzyIVHwi0VSZDRmdOFgz/lVgtHI7KPODjysdXlsTBv5dfMJ50KkOxXrE7
Bi0BcKH+F+hQX88/Qm7h+sfxcAOr80izW2eSXnrcMLwbRD5sY/rK3obprje2OITOjy6kylbmcoWl
twCTMN6GLXdJ+c/hmmHmhcHA9b+y5bf4dVZwiLUSFRjihwu3revBUORnfCLEIYzqo9/DZaYtw2m+
Z2EqjYe66WVz3rjdtWPAi0660NU0C7KYOAIy9l/ppljPwS96hpdn8wCNwC3Sw789NJIfhPbNAxHU
P6xMOhUTLfw9Dw5mcz7WY9Z1qFv572bTx6rPS5ph6NqgGvXxZkeb5Sum0uM29NzxK1UtYoogY2H3
cjllWc4Ms1p9WrsIA4plTjCSkiym8zIFW+HbuqaOjLl4zsF5UrECW53eEZ5rjulMGVYeDNpi/eOo
SBmQgshzmePv5RXSWmslbHNDhPtrrZekMJupJ7Vjwptf76kt+jtVEtrPIg3AxfghnEel1iWTnlDR
rFyJ0So9sMuFvu7C7LL6q1f7jgWdTlDDGxXPv4xKRC56EBUgJ6riTbtfPs3AYn/JOBfJfWBki/eU
GtR6pcZ48t3f74k4dsl9jwFCDeA8ENPoQBf76j2ISfFoyXaFOKRdQfBDrtHJ9sRpzOI96XUfwAg/
gU3dLmMbkVj9VYmdkAH588W4uZsNdGoP9xxuE/kPvqs/d3JcaHqhqU28OwdbezIwzPbY19RH2aUJ
wPmieX1kuzMzdpEFBq0FFMRil3+KujZwTmlWde2nC6iHJDRI6ZYCWDfR/X5qHDi+2s6xQNf0+RsL
yZPvE0THctqiBVrPSqTk11AfMyvxWO4ByMbxWhTPiYxfCBOk6IlUws+T+2XP3ykKwbRFxiOeI1KE
uRew1dnXJ5GwIB6mIpaZzpxb0RLf0mL+NuxpfrwBFjCPEn4JzpMCkOQ3ONCB7IF4DaJKE5o7GvrP
iqGIbKajLTK1nLPtmljhLxBT/ef69kKqbt+stdBg5o3brPpIJlf/+Wp2jaCq9S4kw5eeqQ5p0XEa
l9HfALPu6m4AtR/JjKzVMW5E4hJBI8GudRGOA5zaFKr/APXfGCavj/uUisW4ZH8O0G4xwskG1XKE
xD+QI7kFU50+FfA7uWheCxDE0zxCA9JAdDIocneoVYdVvgaiWzTY4JoFS+jmNkUJqnl9k77V9jAb
EZZ76HmiOP0iaE7SFqrztsl1CvjDD4DoTRwIgXXpl5GOTKfifs+v2x81QS7pHzY/Xo8aGClr/2fu
2AZlL6td6uA8F3soctBPzJQiSAKCxBPu0KKHHvx1LTCgIte/MXA4rn7TT7QNIjg47Y17SsyqoiNT
BJpHb9paOsUDFMrlJyVdZ5Q80lm1/M0rl5UbCpXQcZIo+pPfDbAvUqpGTh9jwOv6IsTHiRcR+QD2
E1KuUf2MPccXVHl2qIXkNByMwCouV6YZY3U49mOo9U5MZWT/RKtCG8DGDxwAAGEvriaoBeTSZtUe
S/M41tvjE7opMN4/PmtYfi5ASBz+71alfblKAsAzdfAGIhRpzmlggcXK1kdmm7s47AhVW8AEbL0K
JUutenirBWtJHAJua3p7Cts059PVOf5xCWkuYbPUCrHVP6i7FJrYcxrcmllxd9WrS7oXs63nw9WG
07sihLZyq90hhI07pNZeL3szZ042Dh/yrTUmkv89m0cvvnRqJRlR+AX6xj8i1QL1ZQBBVPvOCWa6
0FixdyWcC0Kbusvx+wH/au3C6hKNVLdCyD4K/nOk8L4Cuh5UyI158bpQ/UhQJubMITI+4TO5NwtF
AROicZLJrmVECvK2x8ZisIUhKI5vAFkiA2h51tQD8gi6Egw6lc4fAJi1nGUgGXaYhjfpIzZlNdIm
eBmvWhd2GrThkRfvuPwvWqkrtotSgOBFwT1PpGbImXAakLR0+74n/vfYTGARSPu9UfKUStKSCpXw
Abt9lQKa9jhzo8FoFxNXtCmtFuh1stAL5nhU0+J3QF8hbPnZMY6LmP8MLc3SNTzUQCyyPHOIb+xj
KEsuFMNv4ry9wKu/kWVpgCP2H3fFtpYhZItvyQ2QIU/2QWhKhyJiyFTuGXgKAq1kj8UIpKMsnOmr
8GGiS4elvCH6SMB+ZdqlbZh6hKFgsHNC43vgOIjX8bjYKWn/qi9XSn7wLfwA0QRijdRin2oTJrnV
Z+anYwWwwZ9iryBNUxiIMgGka5CVIr7Hi16KZUUnVDWVSA2m+ycKUY18bxa2kOk0i+gJpQO0AZqk
jGWbnAc89eiQcfl+h4MOlZvFzYbu4zuN3MrJIxb3xZKo7Aj4xfMhkfrLGBOEKHGIG0Nw4UT8pzjc
jzr2ARTRn4ZNfvrroEWvqAwCdhTW2tmUmDYXEVVx7FAd5pwKd3CrXvV3obQAxXiP6hoc0iWuFRyj
2Q/H8dObD8vLMAJl0RCwfGBruAmYvKudvhNwvt6UPGc5aahBAIiIsMW3nEx73RVowhaLXZebUBiV
ASMbvj7vhXagrAVyCNkfCCycXj8WaREUW2II4ftDIhHG6xICA8v39jqnkoSL7pcyTwvKYYqy9Jot
ZTlMTsnVMTOr8OkS8V36C3n1jw0K9BRgtgrvYUylOOs0QfYrhr6PribusvGuNIAd7cIZrh0uwMJK
JyDv6zLtE+8RMAs7KUAtNTY/xj/bFWKHf9+Pxn97bFKdEO90ao2VsAUEY6saEEk2xwcXrDgtD7wS
f90XxgV1lAMR5CjcdRvYgvj+gaCBkR9A2iGKEiQ3ajP1h76czh1KRf3V+aYTMJ4krOduyim8Lyrb
1HKPKkgFJL83cU4vXfzqYujRQNRWX5ShzCVkr4+PRaajET6F8DBLBlZwh8lufsIJ6mxVvPGouC0O
16BavUR/NdHOGOkT6esF9r3JueSrn1pBkfvWcveK2Teb4Uc5ClzpGxnDfnKxSOxINEJiArkcNfQv
IEa4azh0eTrb5/ztS59+OiV2RmIdD8mS0brveJgmpaE/Qxc4z6dG0jlBuduFNaL/+zpK/wbXpTN5
86JASHJ1FFK3tA3Eni3BRuyPpdyJcH3JSbTVriIo3DX37QSrmyLPdaVib9GXz/uhjJnVFramZs1G
yYQeEHwAGJA/IC7X9cqgCrB/pBb3cAQkV2UR/+ddtkR02gGmR/VpAODLQH/wkqn/iqKedjL64Ffk
imwJgy8HSAqfClTWl4OT5vIet5UCQKcHkN2qyV9JuYSNp2yKI4jxt2MR4QjiOEaop2bkisKYiikM
19VypcXFtNSMmrP6bUMa3VeaJ4oVj2KRpv0FnlRgNGZd12Y/CtZD6cgIcswe1iU6j4N2UVVyMe7k
0MoG/h80d90lArNXSaR/C12PlWHtAdx2jgMNbNbxsA2UFSOMQYofYLYjB2A5ucRPJkkbHTrg6tG3
SjReeIRRsJgpZqUSlTl6Be25gefO7toN6UAJ2vvrwsPBFuS3h4L8pTmYz6EXWUO6rroYwT4EHOGU
Y+d1cW8F6mjU2ah67k7IkYf8KoPZJC2/xecRQltj5fg5orfuxTJbGqBQgnCLradAx+0AMqjde4gV
ZqIfvdHMkmuxSNnwadumTV8auKkWO6rTYomoGo73XqLzvG6TlmHHLR5v+uunMhinIqAMY8s9j63J
6FU1YrX2Is/avbMl8Kp/1RKvI5GU/dxbpLm/2TRbMmtCzzEuHhZrj4H8JWFf09zVDmJxLMtDtSzi
219ovh0DpmcwHurzaQKJY98QMMmfYNaTT6cNUQnjvM5lbPrbkvETw79Hp93g/FNINDdL75CRSVR1
hiWbkl8ZmY950PvnHMqZ3gGpIaaH7dBeo8V+67qY96nChj4oLbEVJKElKbcuF62Ww8cBSLDL15fb
adNT9IszG9QPqQs9tUi11oBp8PFuDZwCcW3SliUXF354vts0P5BDzZieuJxtynLPB1H5hm4BiN0E
jrrd/yqN1zaDOsXsGZxJ2WypMSePgrrfyvfC+1zacPFOiPKsYLLc5KkD39nExDoiaFdraDCXxh/P
9L4Gyc3eTKHMxs9Stgqgw5+SzJbx7M7uLwX0P4KB5NQ2RcCXtFeL2BZbPMwqU8CEMaxQp3OKCRnH
+dHd51ZyejeD99+sGf86+T7mRntVUqGfq3Mk3DiqufmIZBn2OIHPVkz2nbahW9n65oUfIArOLKo2
QLPBzQaLDPbwnDTFHMGdMONHYXrYIcgUrsrrOWP7p3X4zkD3EcoQ3DCLp0PeMVRLI5baS7+ViEao
u9ZaPK6irxIwqoAxhSgf6P5ahwNHurakuWTca4PVMJKqe9g7wfIWl5sqYM+wcVTG7yrRFRS0EJ27
NDGwxJdJpFZ9LQw44TxjvWgJWG+uG6HbGH9ieYxjpUT1RfBw6nC3u4kSaZJdeLwEVhZVhp1cMhHa
/KjH5tbap6xRNest/cEsmtrtLKaVwqZZYbZF8I0QfGk28TiS/Jd8JMna9caZvXLI+BSO1hxDQaVz
LRN/6bbrnJKbTvuTMJjhbtrwecS/MDHxKCV8s8dbaWNCDhtWhsbv3hVv+iU4SKRGgcsOqVB69qHg
JjPt05y6aTzbgCkCO3vSp5m00fkKCCdwiuoO7sXf640MTBkL07mm4wFwNbrKuuTAJAIID12IlFvn
Q8GRpgkIDLASz37f+Mu0bRIavsyqUi+5ulfxIbSUatiNBDPaEJ7/zc25vvPJMTxc1vKIvftysFuU
HEOUKSA+QhAXdbvSj/s49KraB93+OsjIJerM2hrebTTSkMVRcFUNswLzCld4OtzfzIrSasKTqLGQ
Yew2Mmd7Nl66OQ2xZWRcrFcm1yUokj2oDV0LsqoiV1EP0lt4NTJmD6jpXDFcxOqm+4TFOt2ZrUsE
5XekBN5ayYnpA48dpEdPhbD4UXDnl2I8RNN61NrRyhqPFnRcU3JZ3QOGTR6LNJq/bMLOrxc68Fwy
Whj4Cub0lj8SOvu5ETLHAfSdrNJT+y8jvB8d5HQ/ldgenWbqH3sNr/tGXnJXoddhkXD0LfNLUVNE
6ydZiwCtFNGme8gu029FKPbVbU49jQZekXNerDIM6Yb3Ltu+ncZ+R5Iv4Ax3Ytg5ItS3bxqLf660
Vi8uyjMWDwfTX/SB+VbeUB5FQ9Vh0Z2BYDTXBtzvTmZS9K8y5qj/8YJXpCViaR59MWFQXeb32EQl
3BYf5S6z3XTmgtmyVp93Zimqt7iJxHOFLWygdJPIWBaBjertWfE7RR9B6e/bQwukWINGmYMZyDqR
To8ayqRIkDOpY7wqndmNhZjnvrsgQqjqiA676RIxMjBn7iFsqaDIPpiytH5R84xJ0ZZJORMdUOx5
YASttSGpcDMnCBrNeywMaSDcN80erp5La6IairO0XWfokqtjkBRSVQq+uGQKNt+NxmCDlK5GM8/C
fHCpwz+++icbhkD4CM9eZM2roN02lTk1oDEEoDeqy0pvh5T1oyCnLItpE425Qgf3yNo1cQ7maJNr
vvLjkHoVObzLBYKSeQ48+PpRAw46HVIzPkpSZPe7tjntINHy5x+mnboTEv585sDibMDZfsbptIzL
R0Vw2nP9kcmykiossEu1saTeiPAYhtJ/MiCTzmdp2DiabVNiCVUw+oTxUV21TsTbVW4QB4g9/XJa
9BRKBmz+wWdjEMB16yE01hm8+SXToAJZkDdHgYtG6o5AjzjduqRg+CuuYatj52+Cj+zva1KJiKND
Y5z/XMBdMkW19pRLj6AhNBNfBXIejsuZvXlEKYMy0sIWoLPzFfIeJbV2ANvrLMOpSGkqLxVLSK96
bPVM8OIenN36XC633f5dlfnP20FVkkjENKlaa73VoasFN4htlCjjsWkDcuFMViMexkhLvpeizWVG
RuARjijtOQEQmlgC6ueh+FqvPBkwjSrKlcV9ZX2aTzKAlm+6dyBfBgBo1tSgtTowRTICsgA1mFWg
3fTviQBxYw1NJ0RDm1OE0toCgYKFwA0QVFyF79AqkXjGx9EbWSFGzHMWtOh0RvCLYqBuCr6QWmzj
NOdl8LmTUhGAx5dDmbRDjAAtuuDxRi8j06UUieGcQ5XNJj88wfhFabnN9gOCOJ+RFZpgirDE+xpz
S/WN9dX20qm1bh5k0wP6M1pRJZgvhHhheVN2cKbLPFUIMf73eN2pL1L5yHGySkXACkabQ7Cxtstz
z68KZJXkb97U7ePA0ZgHVxoipj5LdMYy5agPiP5Z8TM2PZqFoaoRATS7j3jJSVXuj16J805I2ZrF
d7ypcouvtCcNFiCgRR9lRtJgxKmJegbL40gg18ZF7ROhjFN7DdRXmyFeCkJwRGs0UnJNXAT4wwaD
wP5AkBGFfArtNggzPDaZm+R1p9+VZ8FeiGts1Vvr/HuaR7jHGiMIP7fbW/6oI76RWbLMQVwg2u2f
EEUvC9/jFiyQm0N+2xGGBrxtOhUnWtBpvbkucVKcSeb5F7/TPtQkc190kpN6ckruq7m6BZe/KHfo
gnnyMYE99HwnTZ/ATsgkybiLLAkH2ugaBdJeDXpJzdm5SBXNtGlEIINChLDD1w+w64HEhWNa8bGc
jfa7n7V2KuSpQJbF1PjGsJy2iy6iX8RCyq4eIZSiWZ9ijjeZ/78UaFSmT7rwI5LZxj0SO5gCt0iJ
spU8uzLtV8QNGPImepvXSIIUQDktMPRgUAMOuzgFwwZssLHI0NhTD6UmZ68W+3q8mv6cdXYHCeUr
VRsGzVt8pD/lQNsvt3rf77tByeDk/R0FvMWAF/NqlulwYGI+aWwnDZzmzpslKlSfXhxfnQHcEUcg
NjIC1mDRhon8WbMZBBoG0/ei/kCnH6V1PhIoA93IS5W6RYrZwSrWxzbn0vRGrVJIRvbWOZxj/xmS
EouKY2Q2JX/BV35hYXm7X7HW1KB8W32bGIUCt8SLm6ojD/0icQmQgwAKB3HYnqQ+SuM+G/ZOXexD
TA912vVzKqe4qqqL8yPeg5e4MpwSa18Rm+jfYfiLsd/LgFJe2YFs6t1+4jDUtEcbXpe3Z3cTgrO0
/Md00654dzqv/PIG5VlQlMPoLo2Ccwt17vQ384y0grZzBtWU+xgvIsiO53fv7I1ln+NzTwCXm5ft
LZd7sTIaTTHuP85xrpUfM2+7MMmD860iyeOHfppZS9YYqBMM67Z20mhihbMdDW5wpOkTsbbz6Kp/
hkLNig/2J4dngQr1hVtzRAnCW3Tf1MlMGZHMdI1gUgd9VlCurhSUf/BcU4GsfM+n0yeLCnh6yykJ
lZb5tAHNM1/r+eXHqAuXuBzK8VSeap0yaS4jwr7g/IpJvM73VMWLhFQfF8C6A4fZzULLfnGoOKvg
yBx0AMhrHURwtakWT4J31qPCzlFY9ZoVMkE/liY7BFYTOMvoPUcoxGkGkuN7zjEpBXFHgLOA/YlQ
u6gL9ExhC8C5BYlpZ08FAw8MP4+VeEvW3LWqniV0soKLPjFe481u6x7LrtTWvgF3q6xJDqsf96qP
QFGTRhd2GVQaJUveI6cNhh7jbeasjdIZbLvl55p+PdjwGMreC0/En0GFyBQeTWyWXw6V0VrsrcH/
mcUi3zf/n2x0s5TWGXwiwEiuFBaoZna3A2bSKzC7D5ct3NB5wnuSwft4EaiJ3mIGL9t/+RAB7ooH
qvpWPoKIIL749ZXI9pxf17lP5Sb2sIDaDzVoqo2g9UBO3ooniAKWZJKT2RHBI88palrV+XOg8Yr5
s/U39m7aZ4FqF4FqhqhBjSK3/KJA+uqhnUeQGlLpFWNJezjyis4bzOHOCdTW/YWgqc+TYBNB23s6
g8G+ARJNUEk1IfQtPebtTYwW4KxBdiU5fTERSi7GDW0sGriKrK8q/hzDzkPHoHMg3suniIr3CNlF
JbLenJgwWr4gXU+kDA5JG4A5QxbHl+9vowobb9r9au8XY93DKMIrSmHPGSky08zk6BL9zhjQW2Ix
V9VKSAS5thyYhfRBlbVITPRgw6RMfuIzyVn2FmlqQ7ZUIqW6CGqv7S4kPx7Tm23kywBKMnSVsgY8
F7kq+Hp2hYCgaFd8wMlDJSor030u1tTqsS+3t3oWMuTa7YHroEodNiM6u2G9wBb1XM9n/N6RGTzH
kGeZhTH+xIB2gH9e7pPm/C73hweNdTqX/izpfFRfUAQaIxmU4iJKcyjM9tnhT0eILhBb2WzBEzFv
vsqZZRwX/ipIwHFwLdksgH2/JJTc4kgaZX9Qif3GDRPRBKoUSk4+KNI00lm82tK47qZ1YFxj8yfT
muW7GC/BHUhYH9M5QrJFytPoAMFFodVfkAvHzAr5E7k4+QgJGKwvhxVVV3Uefdp47EdHvbQqh1hj
veKTPGGgmKw1t8DqfrcIqf+GKNdWRwl49UEIOrkiszgNGGDeMqZxNWdLews4gCmJQWgBp3W1YSHd
aD4tkuh6f+hrl9NPou8AMlrzWs2pCfzJdp1/xEjet0YZq/kBIhR2aA0ml26oOEXe8Ilo3kvjuAtb
BcHhbpZ/8NrjhUtDyyEScjWUIGfaUU66ogBAvTZEZy3cBmLI3cjv7u659LDD4BVKmz/akdHmqu3o
Xr5L1RSDLVclsXW6A04jnAhbwpoDc8vyL61LmR18owWKdaHFAZZ1au0QSuDJUm++56Cf9DTkyLJt
XwhpzEQx5r52pb5xscEhSDPtyrPV9cSU0RKeQfKZ/Q/KEq4lCwYNSdpS8P5mwDLFc9QnfYs67Bz2
maZ49ASkcko9uqLo7JHSlekorsyzLCRyXlGsS/z+Gfv5DvpP8mYx/cUR+rRB8n3pPKgFIOSlHAoZ
AKqFOGS2cOa5kBxc6yyGll2rVKqJzmO1ZiMtlo5zapQRvMMqtHhsgxePXWFDHrWf+Yxe0bP7U325
yHileO2GeSOq5giehJN9VMoRDf64Pw42w+SE8ZPdsXnU4ytMbuUr1Ne1uApM45B/PUNcmQAKf3oU
wQ1hbraUytUq6EQkF+p5eCVDNnyMTlLMKxhHDkIFBY+4KTlPR6sXjX1fiaEW+0I8Nk/8pcJK82P9
DWOoiobN3TBMbJ7FttBy7WORt9uj1+kWzQCXt1LNGfObiCA9kSHWRlQiQg66WAlx/KVNtlm6lHCU
f9mOZTg1qnfUeVdIx0fgOGgxiv0nWCt/OIp7HmjkumkuiQirPTw05vSKwoIEVAY/8ypNNcpZAzrz
UCC65GBqCvF6Xtuw79BdONApLn9QCktBHpdvsaLeDkjNe84tW65llxx2N4MV6vtoq+ftALyTUKMF
g6AV8M6g5kliySVLawo6C9c2/zIj3txMvU49fDsFsWvErDVhvo4NhLhIMUpvimj6CFN4TalMQpsi
FbHV82PThPSbunXTDLhaEbMewkBFXqVSrxSkkE1qTu/qfEEcpYlu3ZhOgZFeamTuhnPsQ+YCtIb9
KVxXQ3yKcQNmwGZZrSzPRGaLkG8ORA9n/z0b28OkVbuA78mF02MmZSnrjmgRCRgT4XYgupORKRP/
Mo7d9JIBBtY9oj+9HprdKdqrkaz5Ptu3HFar6NyHf/hoOxhg+YOOfhpZCdWJKCp/Kf/8WoEUF1zN
kDZ/DCYZezcoPHQB4+TbzZfV/qyjZTMqiD1HGRV0oLOP/Ne/ug0PvhHpywd+QEGU/luPNA1ZQKA7
Vxegidd0m8OmxbOuhZE6qT44lVdEoHy9tKTq8wbga/QrAxRVz/4fyj0iFtLQTwRfwwA+v/lpbRPS
HgYpGWHpGsTFXQR99Ra9IKdKStEc+qCoEZyD1BhSn0wdxvaqu23dg+CaaOIIF9y2AqrNOreaFQ5n
JlLycJzvG/m/f7p7npYlAHzChXMYE17TEYA3PdJXm3omgfQOzYfvFB0YFhvC2VA5vL+tapOovZ2E
NxiUGdOjh/94kWKNtLBMi6qqU6glW4I+QHhtZQ093a13XWqUcL9Esra/MM/UxHv02EDJ5XlGbAkQ
N+sA3AvzbhI5OgYAUqgu/4YfyIZcH94CHrzflZqp6uuLRlYqZe2nA4yZnrQxdHV+3dWaJffJiPir
9+oHQ4zWWI2Fsliba9sdGAUikbQd1FYuUe6CRORCr3/oIYUEB1XTk5f8Oa+6llpTYf7B9Chqp1lB
pmV2719iZdBOROczkOf2X0AidsXyz84OutHWfCJ3R7wb5+hJwYSC7RDn/YMjBF3ympO/i5YvowMc
JIkvNoK356oPqWoS4aEhb7AF5UJj0gnkts1EzT9XpnjCkCTeHm+ia91q8LY3kG/XN3Rew0Op+V3x
t5RCU165j8VBa3ZbqDk/SC5/jG7nXZ/NVRfgvQDHhXugz33Zzu0GvTziPoVdByiUXPF3ceRtPDgz
9kGJHTyNccQ87TA1XWFmPWNvPGddwgQXcls8Rip/m/g4ERl99iTdc+tZuDG6DzuTQl0yCWXrlSk5
wrlatv0qZQSZnF9SOu8iyYKHTFj1BZHGRTYbY7+fYAdcaYM79EJkZXjGDjBE4ZzKMLkH2DijALl9
mX0si6mUPp31cQlqPJT4doxcQK4DOXA4zZi5hHENyz4DQb86nf7h4CBcZklrZLig6/XiBa3Ns+h2
6+Q7BDsBVIUl8+WfEQH46q5M37x/H7E8I6ui2E9VG2luDGvfQUImxCK1Jidz1JeXlzYX84uDNm/8
wbSwkVOYh6B8JegAhBAXabjR/gA9cOkozFIvc0563PxeIqmsEdwV+/+btHBYBhN84M7cICM9xHOo
+btmRjbTrNcrXtcygvxl8yTJfPVnSSGgdaW5LhsfFsSXw/bbUstayr9jUosQx6UaYZ6mkSNMmTjM
4PJDtdUYcMMU138Z4Sw3yPHxaUKbk1/qgywzncSoH/M2Z9EoG+Gum+ZJ5P/MAKADw/+YhkyJn6F8
HCAtlk83g7QkOYpPt/KZSDE4DM19a7B+89Cb3peKBGx9Nu2A3JLjPMa/WbkvJCqYjqtjC1AZTWGA
Lod6rhq35WDmPGwL49U2madxv9i6YvFia3wfsrKMzhEl6cuDlU4Noiua5DbhON+ocITBaWnT2pIr
9ioSUJ6G0T9WA2uX/tHxcB/bi84BhDMWHoB+2y1toeqTL2v0rdVrAtRLPsrE4Sd+1EBjylBP+lwA
OTLeCOIDhD3BcJGK9lLDzWRRdZjG7nccIfbY7OJ6zFMASbbKg22mc11b3rdmGwFCJSGBZI/vJkJv
lQEUAp4th0Qi60KgUcy5AxVB6NvFbOJe+hRjABBAkSsU5XKvXSH0VF8AQeZxfw9Hfh99THHZ+Vbn
6ZiC4Jq1qHVCPujGM/n2nxz0TNzScAE54pwZnUOnOWE3lFRYi/Hi1dpj+NO+6KGgrqaMfDgOUFgF
XOt2fLfh4kAfH5EFclBJVf2nSNtl0Zzh3I2o9c3DaU8GECnt5eDjme4goN36TY8RuKl/kEOkyfUz
FmJ9Z2v5Og5Y1YVImpQCzD7zRZIjPd85Oy6Hi9xNCc1nwez4bU3SOhQXUDFqBorqxz6aMfoT+9PC
CSYhylLLZZfuyzsn5TBDDLS32LYF/ssdGx+2nViW5bwh0Uy49FTPcA1/ZvxzhQueYS+554oZ/6io
+irTp25PiKbOPTdqguxPuNx2cgyJf1CYURW+DQtYs4nW3rL3HVZnFYKhwT8qByljDEvlMm7TSHTv
6Q0IfmfqzdQc5G/HhXN5y9kJQ4/VCdOkYzljdgi/Vi3b7sBpvj8BhERHTriPHB/J/lDgTeSG/+2H
8jn5m0NmJF2SFqeDI4JIONyFLOvJktwwULP6i8k2/yvKNC6ly4JW01erpcVYFQUi61KP8/dserJ7
Symre0R9z7N7lbUWTW/m3OnBCqLOJacQo3L+7ZGAwS/JKMm34Bh/u4+jXLy5x04cG1iqk+gJS9Jj
fc+CKP8s5bs9XhdnH2dbDfewIyXQh7bLJrz+1fRZXmFy3dLi0aHvYMKRaJ1HYpqBl+Jp0iUFJULV
HrDRl5Qe3kRfetUWTyHrID9rEXc7vn32lv6KNhUijddb0uHd4z0V5rXm5zflO2Bn5Y/eJvPLYZRY
RpwWH5DrFTEY+SyaVoS6iYR0fPEAOXXiUqrl6HYI7nbWBntaKl7wlV6P+uAQp9UPmQ5xjSQFFbVE
BNwpD8EFEEhT9fLJw+T0+spycQ0110NmYsp7B0UWgIiWcrECxboGLkp0NKFYYYUr2ilz1IrAJX6d
R21yklhuxMHUfxBz8XKu3K81tuc3X5mIKRbGSPjPkHWGMHU/FuUD/w3Mie+etaI67c20m6ec5H2f
bH6JJO1mLVNBfHDrf1pnq26xPWjnaDYr9CxR2Xk4XrOtGnK1y+FWE2oDM7Z8X+kfl9rGdVlxdyMh
XaLy/CnRn6WhvdGvYT4m8YNad2x00AUKpvkkcDBuboayFcz6vmP5l7mCAFCF/dY6kq4jHE+9odn0
Cyesnz8PB81RJ3jYHFiR1C2rao96LBYIKDpVG2O7dxneRHCMxE1UUOSOhCUZAFmGOlXk9vBv8der
n0ODhX4LhtyrmR0Zd/l/Ta4hjZO0E65GD2/GbOsjcyZbIbCb4AZ/aUvg7kUc5WJSoWEA2a8PLE52
O4He4R83nLeyWA/3rCICESsvbhBU1dZFKATKNTAU7S7YfUuH1sPnqUbwe0TXc7FJmw7pZ9ebnotA
sjTaneDRJiAO8loYfMXdSwWiejIQGtBpDsPGCNGDpVDlDwVkUR0uTpRVdrdT6tejvLV9MHLPAYkv
AIy9/wy8tQzxx04V7JDIjb0mi9JFTrEBiinakmJbJRB1VRtbUKOcAvlYrXMvTRez0sZjhkP/Y/ok
WQ1AfsyFYI+8tvn1E4TNJ/TykIux9Rn5CivlXwDpTVDxgMJlo7yPj09snMzYP8G8MjxJMXAk8E5C
/vF3TP8P4BGPddUqOux0MY82/aKTyQLgOMqJ/M0955XVHmGF7TbdZoBycYnxGTlnxFOp8CnMucal
Iqhxcy8lRqOSUJoUvoATfdebEb7qguhlQ4RjTjmaV26T9d1OZak5IWisea177rTEvEDgIRyKFKPQ
Db/aje12kaQp+kW4SjaySyOFKzv/VNDSDDnM5HB4RauPWPeqhqta7ogl9AOjg5Al9uHwoPMLr0/y
qV9eKd+HtnOz4nsUim/pVdXA8YDnigdhDppNK0/EGbuInN6+ZUQBZnzXHn0pdrrpdQ9LeNsy8Uoj
ip3o1jV9CuSqLjw/w2ooBhbY1CHQyFhjUylcFYwOlG2bA7wipsTsJcXcmbfHcTiCHovfxe8cSybr
hnUWimwuiadPoYDJPXSuFPvybNTqaFLvlY+7ePjFjNHG3V4vqicDwHtuMn91L2N1fqBmD9Z0/n2N
B7676EfjtZ2Xjqeh2qBvewqfQMd2ijFP82RMCUIznYVx24iIR39t0MKtbgDZduzcMcqhvAMp7LoV
sY4uKSA6b3o+eTvPLTSzdpDxxw4bbhf+3xwkx6g/I+xjwz7ayNMiITAREi6I64dlhhkngHeMTUVt
0eHsT0OAB4hgd0kICMbk5FNkukPgeDRQgqQxhL7gxS1g+ABHY1O1/QI2Y/emnsk8JPbUMqugqbvy
dsem14xTS+XIL35OKFZm6cEewMe5I+rPzcSs92sR8UVE9zOkILKyK0FTxR/YJt1ZkVck+kS3ME2p
8o2ruTgLFozZWrm1QSjBX1CtdNFnpTKt+UAPNCY0C848zyx39GFz/qDAMYKoeL2lK6BiF0q935yX
OcRwLWHIBB/n3c4XsXfJ2jCGNjEygJVmPxpNt8012ihS3CIPnYcYALhqubz2zQl1l6Bxphh7GVVH
5YM2rwJ7sp72+6yA2tN4+wvWqwrQQNCT7j7GGaqA/Szhm7jIwlFcCQaCLcQoOVmL/ybagy8MONGy
yoMNL45oRw+1XXcXvwKodE4YP1bSGvvEZ9LPpuy6QHaC2WpWD3bVN2yx+FiwRYzwTeTTpAsvbOjJ
zTT9Ku2gZx5iIJ4UPi3L5OEA5Qw59rUujvZkCIozAM72ZYW6dD7ksFYhg/IaXbZI36uQ3pYkKKc8
miPyL+b2USTJkiCr3gCXJQUyRm0kVuX1Ty7UxQgtWzSo6H/Z4fSatGLeumj3qQsGw5SMCsnhkEJ4
Y8gGEnpNLQ5NLdVAssfHMHgm0eO5IJemvEeZ8aB5ktWQOM/RcIE7cSISGw1bGtUirjSZj1ROJSLf
nDo0v+E3dK6mmQaevw1ZRGr855mhlMji52hgfW4//P4LoRXs/9fGCqYoX5+1szIo/l6CNkv1b/y6
si4kxq8iQeta4f8SU8b1lUV3lNQlHGU1jm5MsKLA+IEdwmLytvd6C6SlcwO9HKreFnzkdNbQAm3l
tont8gRGe2HgKOn5z6kidFvjoLvSclkxI7fkbTvGDfq//yo4JGrj4HJDGJAnovlgTzYUp2ulKsDM
p5zEKws+PBmn5cbRili2E9TI9vC9rG1NLw0kvefBMJteAXXMhUxFotTzGicSFk8Ko8BuI623ltq4
hkWcBgUwpUw1CV2OeUuuUSKTaPf3k58qP7xx/Og7uQIDqAlBa4tsjswsqaCGNtUMxBn/XjdUqzg6
61bVoL94aexz8QJX4vJj9wJb17z8YthXb6z4exhpALcKV9N11G2x2TqugTIy8uvSd7YH7W6yVsEv
AFRUCUF1VQkc4A8P2u/EjOBmkutdif1loH35LtUYsJYGQqd5XGwR+xitduSHjvZr1+K2EWTvlt/y
PJh3M4PsonjMvGcnj/4JJEKtaZcjrxKXYOrypldhpfB7l6NJ8QyGhNA8CzRAahSJKw03bC5n7TuS
38lXwCwpeEl17FEDuN5gUyqpB/yFxJfVNbmnBA56FReT5v6rGHxd0LlmF+9v3pLzwlMU/t0DEy93
t1TmVps3XdLlgNsxvdj1RBL7g0/Bys9eZe5i782MlWPDwWSlEZQqyr1F9uBas62cCkZyE0UzhQnj
6P5BKPzoU69UlzGNxaQppX20rpD+poRB2aq8LJDGE/sN94O7V+4mEKzT8rObEBHyDd+JPZN9mEM8
bumDKhXUyqrqXTsJDWsuIlUxxy48E0R2bFrmzkL+5FiJFC2XeKJfCTYsZ552FItH3ywiwiFIyVi5
4hhM1nY+zFmA6ztLU6paa+NcyJ5qXPAeW6+zXIuaTWcYFVOAPBVvCfY1v9i05HQZlVXZ4ekmSpL0
2g3fplaLLbNqAZNixHMTRilMR/wxeegSBfXrpKAk4ybsc1oAF9TNZWgBMxBjXz1Y7c1yPbiQyOdS
V6Jf405mMI0dy5kmj1KdtMNBOGN4pEsaP0aKNZJHMehoJGAKkFZjbeQqBTbpKeZGb8nzUhdYJp1j
jn17hKoWJezyKfVOWFxa+gVBW33A0ltokz5BfoynFNQAHYTHJJz2tul7hbf0IfOr39QR1JOzleIO
c42bqSF+GrdIpQxpJ7bY7h0H/IBMf7WlhjDj2fjoni/sATaMn3W5inj/54oQ5xfxGwxQIbaRjV5V
qCoYXCXVnybKG9+gB1xuw6bKYnjkrxEWjo9ksxPkGolosczW90vA3FMpbZfIMPMIFGhVd//DCbHK
cWkT4il8zJ1KDNiC5dXgsCR//81ItD1jtXOP4y7qBLODR42O840w1l3ajVcNv3a7JY4bAto5rlaP
/vNZ/ANwy2f0Invo7GGOEYb/6hyk9E9nsw18bVOS7zAgvjwZrK7HBo6e518qnomiF39UumRkwMrN
vimlYGXRQN4MIneU/+ynIhG8sGNVM8art/ECIQeFVHS0YJnNbJ2j4JapIWwOlobpOl5ZPa+PBX7i
/06E//akDRzQEd9LwqU8bE7+Snhx5Lnz7plFAYmLxM8OcE5OpyNcmJycod0Q9rawF6nLP0L5KLte
BuvEXE1SgdCgrfKgee2fcT8lujSvEmce3rf1TsZmJekyz7GbMaihq7wwzEEwr7m0z6jL6s8czSgy
ssoIaX7K5pPBC+5W7DtIrsHL6gNnjaDshbseCq0DtAdglcHi2QDEvXVi29TnI0SQxJtemLoN9X5c
pPWc9tnvMARz6eju4PZyvpj3QtemfFLdPWinsaCt4U7oj9vYCPQOBjvWaLO7cxOKHcr6ocST488m
BA2zslKC/qwouVHdTN6TuEYJcDRCyVnB/nW+8U+Nbn9Sd/+5uIOXoJalXAg08D5tGriZD6/7zC6d
sCAoXMfEUGJT68lUHs5M2UCj1OpUJIFnIap9QAi1KvaCs0fmBtcO1MEbAYumZZZ6lEcJsx1sT9Ps
SHRsn3TgurmSeGo6FZqLj2jHXUKE7mpGudfXe3gak35wkHH2t8XBDNNoHI5D1FFKpvRewfdF56Pc
fjaPPCvktv6s+jLHmwtqQIe7thAf4N9CyaMdy9jXDJwNw0+c1XP6NiM4bDHwmPGw+54lWrPLkArN
CU4wQ4iJHjDlgXfPMOCtAG4Wwzru1asaC5DjcNnT5JnqojwHYVPmmrVEmGlwT8z9UpKSO+ynxmri
Kme2LIijID/J191rCHche1C3u7uuKz0d/LWnNA/P/CgPk/4SnrDfVcWGQjsjjtLKjT6ye5xcdUPS
9QJfFY0KYg515AKYZ4aL8JBM/Lhw+fGUIULDuAZLSE6pvZ0GZiZWPRAW4V8+S4h4geEAxtcAEXnh
SQTnP9zwnddniqPi1xxmhEYcIk3WDiaLG74UtwYZeAqUYHsSEyxnFgeRZV/XInFUNRxvUd6tDusy
ynRm8unZdcAytN/nmhYv9jN3GO0vS2Th//RY3UyGT5xJUSjhG39mi2jxBVO32oco9dmTy0e6pNjY
/wSWj4eNtlwb8W/D+sj2tTfladJ7Y6GQa4yZATCHZoqbjEot2yat4b6TFqP/ruvf5l38VmNWS3gE
r0T54HXwGVnwj0BhP4P4RvECyoks9TNWK+0TZ1Rl6f4zE+4Mvb7Xoy45qknnNSRXo5U6QqgKXWcU
nbyN+IxMoPg2/9mzY7yxwGVjTJPrQnS0GISpeK86NaD8P7kFvaviTIfNmm9f9uyyPVBh7YRgDFtP
IidzmpodxugYlA6J6TjR7GRkbxU1dnVujP2P94cZT5UrymoYdWtM85kE8aP6WXqOD0bD/nk2F6me
vmXvsOOgm5e+iu+6+sNY/76bhp4YnOSkXPKdCN4VszW85QmfVvaE/Wfy8WqLe6O6hOVszjXJIGa3
cDELMqlN7Lc/Qz93/YrSjgs7PTkoOibaDlate5wbC67q1Os17vuvFFdom+rJFLr8JcqTonAviUkH
PSbWGEOJqCqRLNoG2RZyZZy0rlGGbYNiLh0Qbdi8wv6mAIXVVZRmWkS6Xv+CyfNGFTz/P3wtsKYV
ImIBqxEuZGn3SwxCA3/4J1cIfmQVaPG7HHAtAHCvb65zAeoH6p1pyXSl4JAMoFL6gRU6ROx7ahOW
rkltZutU37hcG9ISeJ+P7yLf/0Hx1lxWnqcDB4O46t/mazp094GUQ3iFmx6I8ndpio9b1ip9gFYJ
IoYsRHW0tjFsbG6fsIHVV06wlx79IgClBh0GBWYuTDh5CUs20TKdR4ExyuIL7FK+O4KpFqYMPciE
VxnFfMOAOa3VBPvyNdhKMA4w/Xibuo7UMnACGrHlO6Kw3YeWNMx/o3LEsq8dPbSgdI42UhmLmgUi
uBgn8AjV9BuzrRiAO2DJwtfqBkhPHlDtDMVQc3eLMI07UYCogM1ydOnmAv623NAozcDOEVEIj4pt
TyfMVbsLfV778Mbva1PDNmzHPGuaMp9Imi68Ez/vm1vK9Qcmj9diyhAVass2SJh4HJLCzvGOAJCo
kuh+Pfiag0HSrG0ENef8IzBjP/9d0OtiF4p6qJf0P5PAQftADUTOI98kn81NRD6zv7CxtXqCVYX0
nQwrR/4eeP/k6xpgRhRWnR5GGYEQJnNLAa76jr2AOLCNzMSoL9NY1Y12TiPJvAHgXWmDN70CKbnp
WnQWHd1fAn0zULnJtchaxmbspM8QoPVYdkYCCXZqWYN7dbUQCrUj1FkB6aomZXEdAbPpqXdQuXCg
QFwdutKgZtPpqzwR0+AtU0AurjEa8LJfrqw1aNBMk89IM1AKOTA+PU6fIW0tsrUKYSZ4X8os/aDV
leb/uVqK4QXRWAAGv74cmUIEA3wY73i3G0+rhgFpz5IR+O3R4jnC+smK7vhz+peXgR4E8hLelBMf
vxkpR9dXQU7raPO1lk12C6uLybM3EsSEKvUCHW9Vp2wtVwAmVjuwf3rEE/Dd6E1dZg6pTWVX+MZ9
tvqXJ8MbjvSYr0Im826pdArp1YVl0uEBKC2EtgSGiShrWExvangEebeVnOHpYSJSDOsRc4a5nAtH
K2q0FFGaqVFi2RSnOgdwcgrN7Oqet3IEYnIFv5iTtS4twCZ9/UHSBvqHozANLC1I7CvHyosj3pZz
WhD454IF6pxObUg4vNg4zUfe5GoMgPWyA46kBoQiKE4/X+akwbv3UmoYl/sFkr3akC80JBjyuENC
RNClo08mb+VFosQkmFfDuIAqcXFQLR9GVgd5y2Sim2AXePXJ2CEXorXjV+xHq89VboQDkBmIFLWY
iEsXB86AVTuVucGlqzpWAOq5al/t1e64GRZ1OkIAa1WS1koGuahYKkeSEVIGQ9lRlnQDKrSEaJEh
CCu/JFhSvqFtHEA8uDYvDNhGZqPnmPWWpVUuX8VscV+E030Eg+hvhQU3bxhLVvPwu7cM1eAuUp1E
I63pgq19Tnz453rqrI0xN+XY5veMiHXRCg1PMETuw13qApJfNIBUjaJRY0Ry9CGNLc2BvZpjoVGH
C9BCNld+vrNrgPBtgO8ELxArPK18znJIM8BGSJoXF6/dQ7SMS49v/vicAREh2R6uVc4qk62jMeZY
BmXY1IhuijpbSuQpoEJzO96nk8YmWWdIJnCbKmCHRPTPE3sC1TXWltWMadGllZQj2xTwkywv1y6b
g5zg52rbZdyIf8UXTV+wbnborM8yeDGX36mP4y4U74IxoWoI3BQkgVMm5qQFt5ZYwmIImABVvQYe
q2b8kyDn6mFlzAKl6HegxUfPpsO7s6OO5Xhn/xEBxj927vS+jCj/X/90l5qLJv9qI6o25+1IpDfF
wfAnI0hW9jtZklBEyq1X9znGl1irn8ceM622zuYDlOtiqmgWbmDsQv8Do+10u4dN76Fe/p2M1f4b
KltLWWdR9s+k7CB/o8Q+I6HNQp2FqgfDyC5OwLiOCMw4DAZNv3250HUbk8HgCldD7uvR/peeC2Ds
CMu6uZ5yojg1X/oYZh9vBQF31myAlVTjjVbfGJMFn2LKiSISIrXF2sb65pXGjyDU47vuCrlUNWgz
wq5unaZm59r4yxTauDHkx4unS5dznWRPx1cU0ADvYU1C9wSCwniRo8DE8Uoe+dsf2xagrfCe201E
qGOntHmPqofTshRX7o5hJpshxcHm/grXcsKJBxIN6wNPU5SjCBIkCNR6bNanvn74p2xftfQLJUXR
qsqvjbHODXFE6YasI29es6BS64m/DisZT+i1SkWxEU6k1SPWvZlF4YU1NTbg/6+m4qBCFcUqHFc4
2lmQD9XfBAg4Je79gszBaBmSv+qUJQUdcc1nXlPM2Bw+j0uWfckdQmURNACOU9I3Qa9uFB78AxOv
sV7jQKV0UGCB9cqQbK9JlxtfOKkKsQS6ebs873AF1ArhlqIp0n3/EFZOMkH6ehZU7yL6tu7b/hZs
n1TPhmON1H+soib1cD4fBGj3hm2j7KDl35Lyv7aF54rmV2ZeHtFsPvPxBCI3WbXw3TJCiMBzd53l
tqseo0n0yCIUCD6WWTXVQAP/uHV9wdqdyEDWtwpGRLWfz7YcLF0jN3Qhxh3IMhp5eIZn/wbS2xkr
nRTVu1pCjv36gYrruvDdBduxyWeb8ryvT5jgf2CRNpLdqir+qV2qfCV1TFtEdmeCwIB8Vk+rZAzW
TGReIYUe7+stjQ0K/n3sw7Jjh4SMsbWxLIppGzqPSWn+R6TIcShjRO1xEOrQA24wFH8+Tskd/7jE
26kJj8279RM1axb1Xux6AapSQIOoK7BrOp0g9JkyegaJ0k/ajhTaMyIyfTKAG8Bd2d70WvElXH4Z
AGzjuHEbpAkXR3S2tjJ9MZJebS/8dthkOq2av8IlVkdoKSDXAqN/SWEtxd6UnuSmfIGkHGv+InB0
WGy8JD3T7jdl7/u4prgfllKh9OhHMlMjygTaxkSZs3hm6wTxm2VDF0V3DkuaYqsuots1jMz5T42g
gzC8NTsFEukwpdH2ueicQQVYYR1gNyeXHHzqmmjVCna/xnk/XX6uFqNTs/n3ttWIA3azXqhz2xU4
jHzsPaVOKuiQ+EGptQ0ix2nDSb9gJ2icZZ9C7Vnaa1U9u5uVBr5cCHdQt60wzeysnGsK2y8KfsCr
6HtGyXNA8/jkOcVzy946virf+TH7uZXG+42rHWV7TAUyZp84nFvwNYS17Yx+CmPaJr6G4wH59Rc6
vudD7dAdcc9AaLvcl70nT+O0CEHeB2NwjurT5blIGfrYmhZC4zYh0dgF2kLtdIKVGMkUinOVOB1T
vbehVCFKhL4ZlvlWKElr1ajC85ALyZwzQB+DsSkWBb+/eIfvfG9lJUaF1Dk4xASRtP4fEtZ5LgY/
4ut1NoZIGdXs+FwfIrUtURaQskyWGQ83PlRrPglzgfPH+y4eHConJpD3nxE5m3MHqA2KQicWTFnj
MLb3egcC1x7bjxA6AA6HxnUdOUptv5e64uNOXk1zOvE8IYXieqI2qv2zMvu8tnqGq9Y7RjMFylh9
gHUa2nI4IMwfMeCgJHrwq564oOINmfKO/zH0h5d86s3uhL+87K8kx3bRqsKM2mapAQgrnqv1P34p
KBPK+SrPqtzENSODfZ07uoMdycwjlAHJOGT7a9dUj9s+O8O/pObbsRbNw7QpFD+ukqYZ/uYWYd2E
M8wN8jmzsSEaXOvYYcIZETm+bFUfxlw35c+4JZMRY2XOAo1gCz9vYz+H+vJC8e1NjdyadVzpj5yz
5px1IHbCk4K+PMXpFsfTZlq+TvL/2K4iJNOGwLjdwG+4Qs4Q12C1scuhnDJMyxieMmT2rnMZJomw
l4+48AdMJcQdHF5Gk1ab0Z/+k/cyPxm2k2KRaEMm2AkvlNjpYJSmgyE1+VzabfC0TGEalKaElmhX
TKuejQnNwAxAdA+G/ZH3MC4QEP0VhEPye0NKSFnCILLS9qcfyW/UhHhD5lGaG8jf/+DVddK2qlOr
s5jaE9RKFfsEyjmxfoLWZLBwZ82O7zOwT64alQFQmSIQ2Enfcr8GFjbhHMRr7N4PMhTMN+/sGZ/2
ey7x3k2uKEL7VQW8zKA+Y02kdxtYqYy5fSdLXpSWnjHYeJgBw1mXFtom3X+5u8U7kZ0QTkHSLPAt
1jTSdaiwPgw7+5D58+HDCEHs9Jq55758EQuNDrp9xAx1FxsLZ6WZOgBX6tCNfC5bhg9d3nNs1YcD
kMk1Ne0Pk2BOE8Q7i4E06uEgnsWfwO7BEa9wvUoPhY0j201CWXviizTiK6hFQP31AMyleq2yjCIx
Bpqlw3tULPmPth4dyaI/4cfOKTUvp839+np0gjS+0vkp0tiqfAIvRHdqTOF3YAoGMsdxe3WXxcpL
BLLwbRIzkIjObxwyeA6pW860aPow8CGmLsYEoqj14P5LaXbYr21RYIniEX3gFFcRjaL6TLzA843u
85Gw1SDfkPWK15Qp46eoIJGpi6d6yLwq/8bFzrBclzI89kN713Eu1uo1YBFqTtFlYC9C2Dn7m8k1
1fPkJHoSPXKUi+zDBwtnDbo5p9X0MrRyU4SiDSTi8qcmjGVIv6PF7+uJtAzBxy0AmdfFFcYEl7iW
khaAYrMYOw+kM05hbF4ncuxTRA7O7ZhSCPROdjMlAGU5q5YWBku7ycBJB4Yi/q8F7del1PAo+7IA
iJYTtIRlCEU1UyoTAvyFF+HE8sahtZJX6XiQltTQRkj0OSQKOVWpqUFwouP8YESilW4ve2KRv7/g
vV6LS5XW377tVq7OvD2rojIG3p8cVxdTvWsBhj9AxsD3LgM4vPZd/OxYmRp+ue7ecT06m2bxF10E
DpQByfrinjH15ZhMZTgz7hvdky1bPrRy/KNUPR+8VELsMS/CFFydU0R/gNFMBcnlYEMyLgiZ4aDm
kfos3CjHBwXy2UCGTpzBsGTtQ30ar8NFlwY343aUjj6Q4auWeeKBHIvftH2FDWrImKQY59lMOgoI
5etNeVMjszUEYFpmq90CPdz/IJTbtG5mg0UbSRuWMLHGuO6qmRPiv1f7tTZqMC4yXARJZ2b2Lwcx
FGPhNJS+/TbuYfZhp8yCwBT+Pmd9Ux/WnEhpzztB5E8dPVzQpWf2IGN+LE858D6ZQjT5gWZDZ2w1
lYzOXtgwtKtos8nHZqRioufcHVtB3t3c80wRtRqXIX3Wo3b2Qz3J4Ycu8nsAVssU18Hl2ZyJX7nD
5wwCz6GAbkUgKLWG7DXh++jixPbZtAGUndTCiS/WG6hgTlCD/gKOAfI2NQKFgy5OoLG+HtfnM/IJ
rYXDhAw2eommxxWU8jZ7+SpLYmnB+yWD36QqPJJuV9oliJd5ORIeS13U81Qa5zF5BGzEvcCWauaU
ZFYq0c5S3mBFpowxZuQWjjSyb1RMJ5GqLJJgufvxenCKRR31BtOSgHvES5pUREx4Cti53lv+MEgY
RQbYcaf3Tmk6y4bmZTEAMuE35849TCEvn2R16e3PpILFCF9ScBUUJFL2B350R8558HsrhvZ3Xv+V
eefssfSmeM+rIO2iAEZqmj5QPJiFQ42n8LufWwJK5dwudSdtBBTpL3lrBT/nEgmkL9P5aQl0X5xY
hQT7jRrFpCONmetI33g6E6PCcXiBC81wUQ0L2e0nUE81dK02kMS44xQ0EwGFICk16QIbfIX3Z/+I
2o61arrmOzdmm7FOW76LlBt9S9s2NqbtkzTn6rPtj5JRDQfGm6CzycFAC7U+rQ0RLMI+ryVNjFIM
LfJqgxIxpIxIqVTlVG8on+LDwmO8Jrhp3qOxz7v4A0xoTTexPxWE5GlnWctiUau/Ac8fKetDXJqq
wzfmj5OdI8eXj73DRhigVj/RyxVSZ6aTnnKcy8f5xBdRyLqNag2z2466Knjq1XfPKJSI9iFPp3MR
DnJUzKe/Zqm5Zj5FJdwOoI7BpaRvpooydjzzclrT7e54eu+A6ZAY42v5sJiTDATTP3PvvlKSxmrh
mD8cqfiC97RnUH+Bh+x3LM3IzOwZmYMt8gysG9xooUHsPzVqLQrLBQdMWd19ufRTrOxaLy1CTE3q
h4l63RIxg6M0smjaYQuxaSDUZOQQryWRMZ9P6uMO9bWlR2+81wVgLRap/e7jgHU4ylzWU9IfhZH5
bvD6zKL2sdFWztmd0IPrCuZyEv9AAOopmb0kQc2jrSQnwc2dMZSQsZOlz9EHSNaC09Kf7rKp+ZiE
bVEa51eR9zNAG/KgXGdnSrJH+0QfWS9gH4tmspeiqL9rwQX3Md8HiPg+w/KK1uWeWuBpZWrxJjEm
UfY2xmaH2+4eTxoJecNjwSWqtmFsKwlZdd7kqRwdr7iRNzCROGE7PwUu6G/B9ATG3rDkWOMvi5s9
1vpgnYA2vU6kkcDz5ZGpj+BvNbeAPI2lR0JcFVHeWKRAMINALg0eWg7AjsHoif1pYvjoTGKs5VDp
HMrIWfnQMhGqy8LoshtrS3cpZjFl+8yYkGky71zaloZrIdlKk2/4nGmmM3EGrGraG9/bYB2f6Rfo
MqXTDKV/6sXZKSVWLRN+7HRzSbVV4PwrXQNS44VxAS9/70D8WBPVPaZ6kj4//O+l0Px0lapYfTKL
PX2/cQIb70hjWJUJASxSPYwdIQaxEqo8KluWFHmR7kA3OOnb/haRPLSlpzYCIlYyjODis+HyEekP
C7+CZdDQHTNT7eDSCIVmTJAJKU4eE8hhlXAnf+J2peEQpoWf30KJoc5QYJo5rK0tsLQO1IQWcft7
NRbGoFZPZjs+VYn7GWYs/iYilIfp7FuF814t0CTIoQGH/hYcO4l33t5PD9djgVaykUAl4oFs/H38
QvwMfIZxGVhh/OMH0NT3UgwxmjqaEf1qMhHwZ/lKPuuhRcPEPAzN9ewwbqvhUJhKytM1DiR7c4mI
fxqGXgE91ThbYzdNMDsZP48FnbODzzfyXNBDeQC/hc4/2mr9Xn5PQOHDUY1mDUAFyUebG/bJ2KE0
nn/kzT6XNpJlGQUi09sdbA/I7zWmXAclHccDXyhKVg7saPbs58ogP9DUV+WreAmDTaYEVoB8rBpn
RaQYMN0EJkUAX/G59KqbLBpK/UNwSb9MBSgvtpWs4W5cwR/62lz6ZWlCBouQ9iK81B2dGGJ2wr7q
DO89IJfoTi8G6MI9QuZqX64DQr9w23AfvHoYdSFuAwluouiu2ZJEQMXWpq7SPHnPyhu8pGATwQBr
GE+yYfyG2Cw89Lt2/QT8QzrRwsN7PjvTm7tqG3Q7sEAc8E3gXcBinf10g5enl+Fa6N0zVO0RqECH
Qlc8TPW/d+hcjocE3FKJHD4Zg6n7D0rpiBfsbdcyfVt1moDx4ptTer0Gj/urViI/d/b1oDiGsZ3m
/zmciP0yFdbOq4kPtRaYlXJJt6S0GP9XHD6zb4b5yqj/lw6tDuJLDhi9qeyamtuI9i8PUCcY3c3T
VK9PctA4Iu0z4c9HVBh4ZjL4MWMDft7j7I0SROaZ++qgsiAm74WnoK8xm4bzdmUv+XPaquJdiLbv
U0wJmAhJFQ13tWGWfVzWroXff7DrOE3aQZc2mXyxGO8A+groQq701bxbM8Pa/MRf29SlEOVwQwPJ
4F2NuMQO9UlaGwSV6+JTbouWjtdHCIirBc5AH5anv/lqw6o8KM+G9eM3t8OlJiKuCt82eiOdeQQt
WccRZpJW/v/0g25qJM+73zDeTEv33oZivMcK+mHr1ptfXc0uba2mdI28GY7pDj8CvM+bF4N0/jHa
0bwyT0dLx4T39RtgDczP/2MJcLgdj3B2ztJoLifDG+ZD6de2HeqRWKT1Lbyscntv4GfNNqWI2fm4
BPOpMe43ROzc/q7s1CGM74Q0VJDDEL+1s3WqMNsY9MqBKwTP0bXwUgDxR/OYGtDSTMb1vJ7dILNF
jhVeVKiU1044vyt4syyp+YdRMDJyhTH3x4E2YjDpaRZjkqDYtV7Sni9QMfu/Vu8LW8dgSr+VL4jJ
Ejgi27tp8PsB/Tho5Ox13SISL/uPMR4fSFkVuA2O7WqE1+pC2Bg/YhI0larg3p+YD7h6+cW5hb/n
96p6qOLpYOXU4M2AY5lxQmDoKG6/yAXOFRZvNxr+ez1mbOMBiK4JjHxzxEB6ZJ7hoNnNzlBpXoPF
5WB69mEl9w53rwqqPt37lyZ08y+6bcT5ZYHI+La0Lpc8SCVOfJWNG6hweU6kf/eZgpkVhgi3FHux
ooqBUz+1MgMQAmdLg0C7SdhGFFVnqoQGJX6UOEEh3JT8Zmj4r/nKMMCW/Uw9CJiXJUOL0Eucph61
8tPkkYZiSHD3D3kV7aDBFyn0apNvFX2WMaitfbGjIvEzb9A1l00UyiwyhBWuIt7bxy061mkb9LkY
aI/kq84F0SVPmGuWXdYIZOwufWOYs6HIbt8NxNqpyQ+X5ptxxpGCOH65uKJVIAyl09cSjyFW8gQ7
ihDxxIr2S3MxQrJ6CcOxU+7VyA0Tu5WbLHJkaDlFNPPYSfXD2APj2F2c2wlpoZnr2bfAS1FaRjqf
uVf+pHgnjVdyC+LMIWvhnpXQtlNfVm9i2d6yAyWE84ByLBr8jEAUQ6sPWuC7VUbxNu90KXuazRMU
D1o/oV27UlSBlcyUE0+xrmlfLruig7lou99w3h2KRN5fF3S+sFj+gnEc/jw/yF0peQrJylhzmgVG
sMIufcLdqkAfRDLVZcpoiu/Lta7T1U6pmUjnUuYVA9j11ZPpifhx8ymHJH4jEu61psQeTBoVBPnR
CaIE/c8BVDbvLWwtySMqQa6gikBHlABZ8yhkNGqjeNQqdQmEjmD+WHRegbm0IC7q8B6q6ebYyl0d
3iWFUIPoBzqDls31eF4CQ43ncWWYg2y9YVe9yI0aCG2ylIUWMKCM0QJdmfs1H88V+PMk/BErBul1
97kSuvbUKXjoVwvZ4i64nWdpwclljx23GVu0kzSY2loGXIj13vGKzEWaXb1gOec1aBCcpT4rPPAy
JRz57LjStogvgSX3rzBgERCX29u8vdFvYC9ynZ8RNol06XPCQ426o3ljlRa4kNDN30yUvSnp1pm6
AyKp9kufSup8WQ97s4cFnl3XqqBVwIgUxrQslm+BvFZcesjyv7n7yGSo1B+RXG8MXHgNTSyXwnld
gsY7wR2voPhpj8oX8mt3Q/8asV84lSsRP+Z0OMxzWayplGJedWrkLOUJaNuUPWsnlMQs+3FmxtC4
ZJraVVBgszL5FcrMzn+y81dfi6OgmulXzVoZTdN/Ut3h+i5K3TaHAk0gFCs8i/lWmbKVYnNKQsgX
tsIFPpKWmKuxQpHlnqOp9qmnCr9JI5i0PuhEA/BLvV1iIoDwge99MsiU5xOef2eoMxr0seR4FP1E
jGNTHAV1S84Pm8F3rxk1lmKwyWwutg/GwDwVagUXDGwGdV4pgV3wn+FqiWrmNdG+6tHYvphSqhNZ
8Wlu2J+oFjNVRBavxLOqnBQt/Y3VJg7b1LQCIyYw5PzAG7N9LH7n68tGMqbEqS+BImEWdq9ImcCd
lem/aycZWvNKQvrlr0GezyBfFaAceH+FTwWwg6bvxyHLclmKI6T1U7102XcpcdKGkRTN2IhjnPTt
yps/pjPPz0Dr6ZIVhHiorCC/oHh5987o9siiaKn5btmEe3hAWKFtwwoOYIav8OSkE+58R7hfIpW9
AHFoRfnRx0l/lipmL6OQ5a4jZtdm129tsQUGV0TuATQXctNI+HrmnK5E6ZaDF/GDl+JuGZ2CSTmx
NkFRWWoaVVNB7Y/immvYjgSlg71Q9xkAXCERpUk3GbGCQFdic31W30lTeIdOQSFJF204NyA5DV5Z
wpVTPfyBPs7OXYmVkQ8TuoZya2sCNPDTU3HFzg01ZXe2aF3f/GqIHyW360m8F/O0EpnyNOhJ07EX
fslLLVPxmrpzvdulLagoqLBB/HxpSENUzBY4xoWqg4QHDj5xPQqw2KPtiEdFrdudvwzwOo0DwnNG
0mrOJVgeVcqGiX9llA+n34Re6Ui1bpyHp/4nZ1dPqVW1ubEB0ELKxpGb2JIJLwTbqOy1FEYRXnEG
oqdsZo5ZLDQeF3mXroJ/zeX1Z/qgWgrTdRfWV5VZVmBBSoNu81eUE/99E6wrSWvLp25JFcwEqJH8
OeIshVNPJiahoJvs0+JSdqyf831fzVUA+2Hf0xw0wG9ivI7W45IWibR4j3Y76cwUxJB393RUIJTW
IXJpynaxxuRJiH3Sv24fXtHX7z3qiaHaCiaRGWCW7baOyiIn/sooysd1ohD5ODKFu9oTG/DMroz/
TQB+qeInHiUbVlBkDPN0RGOUI8SLYHcOqAs9Vg3rLeAQBwspAghhCkQlXq4kfXYleixgusfgnXoK
hHUtEBmcS6ZAXKgk04H9DjTY5uJ1KWHWTDAx2veUcs0SloHgxe1JbU2aqw6JFfEupwBvpREt+W0/
aYUo3VjnbE2/M/XUSwPUMelL64JBRT7es2ZdDAFQFx+h71/dL0o7U5C6JZv7sGLxmyKEWs0KqSlA
BDTCP8bKtcuNr7j6w9K5urx6dgQgFaXN7aMnaOnWl7+ouETOel32alDaKb6d4jvzWjxr6VHW01Ke
svFoEPc8DmwQ7jXMyFPvWREM7ietOe1Ec9hcNMNvhn1JFmAIKiuGyW7eSjGUFnKAJT/OZfZpTKz2
tXlptMCxJtf3P4iHXH+zmlbSiEsKpo7k0exRamFaLff5EqrkM5o3HNB984MINLTG2oOu9vMx8wAV
Bm88un2cJw0HYnBi7EI2JeoPGhD5u4aCTFCgjZIkKlDAxXPpwOT/7OU14Tgz5XLCz3bycqbqoKcH
Lsa1gE2U/fzoBF0YiLyv08lkCyz4pKRHz0Ei4CFC/GNpSYlPacu8r3H1/YbPJhHahwzpx7mgtIXX
2MG6hBIQ9FWUEPLI1BN6O4JsTIrFtnL8+Vt7QPK+9wOQ4gfHYUM9GyNgCGOGc0N5urp4yJVPK37d
vpwqWlC580tlWztBs7ReI+5Y5BqHBPeChJB8y7YU/bGECUS+258inFwFEgbbN32e5TnxoExKISnO
8wwUmD5VXlaumwnKiCvV0ZtJcBB9mYvEXGPVWKvfCkVLojYDqgD9irisacyvtrrWQSiuMFVaaZGT
B1NawP6fCO8uPBy/4bpkp6mD66BzHd4aQohO/uEjJvdm0m+yvsDZZzbb3lpd/CLO3oV1T6M1t+sC
FqH3iZ6Ep8Eeq84tSYERPHAbAqwIpE+/h92nWW7AqLFX3ujU33GrTGs4Jmazks8MZxQzZpaVKBr3
x/zv3RrOIQq8kOtpEfikLUvtlJSzjmHKx7c0a072KluSNJsUdXo4N+NNA2G7pOSPFBt79DEPTYcv
wR38h2h6rEyJ6z0lXHfFgNWtxf7Vxd5c9Go5d7F46VpRPKaC4nGMZjFJCuqy07M7BomWvYCuCuv0
H+Vx2O/NnyhfMJFCBirhp+JqeMlM1Aqu8YL25ltAMgngtNJ24Z5LzzS5RbBpHgj0cc0JmV4w8zCo
CekDHA54zyzkwTtI4kcFQtOoNjWU2SSFcmCvfZUGvtIyb8Jy3HawZfFgd2wS4A/ue5dTW/P9Xngx
uYoPQAgW1l/608wUW6WyEBwufjKnVRCx6jWA/sBfO6sAWcSldnEeHR5vhbNx5RZwpaIwWz89Sxdg
HWE2k2f1ljzltnyaUBcSUZEZyf8m8o0X9nb+qK0ULyzXQi0MQkYccutkKfSQcONV8EVAY2VRmvjy
qft+3BVkQ2PCSr4BHnJGfIr1YtykXczcGUAydzQGXkHEHzsFBzjbQmhoNWjxRRX6HcNPrPzGifB7
bpRURcrWvgwV0dA58BBqzxZM3CRTLBkg+7oZNH12hpUgwyiTFEE+1E3dZwlzyPHeaf4JPnVxeI/z
9Ehmwbdp7/Y2GmDpye1xQmoOf51jngfWmyT2Gi87m07jKJaxeiPrtRZfI8thNaEaboHBsKZpTodW
k/7T/hPlE9sOR6ewKMaPD/MEhh5KLfBS10k+6qiCKpg0GuenVPXuSuEx1WVLtxPwHcXScgW9Sdi+
f3KXua9Urui6SO6OCpyH4MjVkLigfIzIp0UzQgAjL1f1HO6q2tEKRkaj1drLhY0DFtFYu1kAATI5
ME+p8J3X0IfDVylyKcmgYgOIFZ+8yhjK7V1248sYmDRmmpnUQHNb3gIcCTWvmW6560EulrYTSrT6
L1jevIYXwx5W7akEHJymmJ5UHNaQ6fiJdxcz62s9yH4lSSmTsrY7Wkp3wjYK5/UZN1yMfCB32pID
WJhLGQ/e/dTAGrYE4xGvQYXjZIpz3Ln/aHJ0l+HqeyEMxgynkoJv+nEr2sUeuK717KD9J6xHrGvC
VLJgXMWry23K4GxIwVOCWzrZQ5QwvF8EdJd3OXLM/2VVvMUi5nHwrfbRZlgVdI3RuS+3j9QtldOb
kw3YC9ygbg1U5MgiyioTJJW5b8RkcsU3BbbHIDl4/3u80exLfQDDxNExBsYBL2MqVJ3/pSDRcK/D
InesLEjOWfrYDCxpaRBtN3JIjXBZ+1LSEZGpG54x/6ecVQzWKjxam1OyNpTv2aiuKfyMPRN5UFnt
lapV/e3YkhmS2ABfyVY95oklhvJrC7awqsJW5wxPEUutM9m5vL6yQ1TFoYof6qDC/sUrfyN/1zg/
ytuhlWMkP2yfyNk2ZuVE7BhyF8sLGT4eYVsfDdOSnGJCjQARzEZvLw/3iWQfZ2dVRjA86mmQnNH5
ZwUa0TN/pl/gSrlGa+pk8cQRPeWW6Bkb9BS53NrXtDCJLG6wdcfIUBQwxkXOYS9RsRkA6vrevLug
iDspML51N3Q3g6Ujh9pzH6HG1PF839s8go/pzdR9YIfd7vd9/YqXhfW/5j9VNybBN9GIiTkliN25
6D/9/dLmEsOaRfU5cL8rL7WMgUFU+Whug9u2B2Xrb/oOQbqKjXx0S8MjdK9urST5veWmxhIcjxIi
Ju7vVfRX5kH8uabYqocneaxvGmbv2b/NuqfFo25KPdEBzmIHi42xY/syUpUooj+c3FzvXW4Yoklv
duHbrmQPDEmBuyt6x5YlHrr/83RLlaNmSHVHfqtOPI5aBN1D/NYD81sG4U22vcAL2jmE7vsqTvzq
+2IHeeI0KI4oDo0XW7Yyt8WMOK4bjzh5gA6cdfSKlOd6GnW55WckiQM4uY4KNyrnXhKWlpQkyen+
ibzTrNwSbp0AgepWsZVHzb4JV2nlHUkz3QSLSmHIfHGLNiRnRKfkMdwRqMRKtId8zRU6JZxqsF/O
DviBFjThLASpHz79yciAnkHt86oZczdHBUG1rb56jMnKdFqgBMB0xrk52dyn8O5sFWi09+M1zxTS
HqNRxXLdh7GB5chrEpCGUieXEHyVyAJdJGDE4HLQ3JSIDQirrUBwECIbSEtrdsx8JCwtO+IwmHeE
jrzBAL9kmLw09vlixBDnMKs59o5sVXja9R4Q0sYvpfE+K31B1eWLIkZO5CHtEn3EdPat6Ly1Vw4a
7I1LwOiFeQo5+/NtE6Jb9uDNO/Lu6gH+lYCM61e1ux19Cp87nCDtG8aHYufm57Mmq4QL7vnT7qPb
uyHdXfQAA9RDtksdFF1cXsHZ/EZP+7jTkNSKuY/wiOD4rXhqXFerBnB5AM6M9ni6wwDsNmkrcqp7
WNIYqW+KCJraortIhe/uM70gFDqR1S1rKPYQMn8XsMr82XifPwg/uLvGuWFEZIKnjiGEHE94Mh1r
MT9vbbkTwxK74EGR+UZhMmTqCYkjcle3SJy3TvH8w3siQNg9GLgjLirRkg8oijYh+cZLUwX8VgJq
EBol8ijYpvaAGntK8/b7l/wkj9qcA5ZZ/cCEv+aCFKGrmRjVr1jrg1ijk0o6Fp8q41BZnIG39564
lFPdJXsceBAxWzO4MHU7lfKkn9TisYLdxo0S33TiTAOA7BQy55BrWYAVWS0ViUa/Oc3bhg/pP0Tc
njuNnc9CCkHZ2N7aeptLm3ezNFmQ2mr42gh9J8+RpdhVxlznLTLj3eKpSQd6+PaxXZs9PgzJrpZ7
bDOViUbh3JPHNfnaaS7T5B86H9cEQZmoYcFoOvDkttDoKK6A8vdVT9qjQpy8FLZ6hdkoYj1CQzGh
57EUMuOkKglibtzko2ySd73dvzsttw4j2FtL/VfdD8lqAumAysOoGNDsci9OgyBB9Jwl6QjRRemZ
JgVlMVmQaCgw8fV/2XEWfZAxAQi19pLDAp47WBeIcl2mLZQm0Mlbt5sD1aXbtlGVccoXJesBQABj
G6qAR28Ru6ch4DwMjatZofMLNSJPlSo7RfpoNp4g4LuGOWbCtUf8e8QqdX8TIfZeibB7HmUxNlCX
RIa2cyrr2inrUv1iyRbxV0zfqosPv+7YZhS2mSCI1Kzh1QI69W2XwXG0aoO8y5h8RNSXRSwTPPtf
Q6gtPbnGEYxbgz3H34Z+ND6o0ejFzKnHMjWpJ36H4DUygPuCQ4VE8QXjr6XMzwEFNBYUo20UUzBr
AecEnmWrOpJnoniKxw9wgKViC2mkWMlcDQmLKc/1KpBMulmRbLhgHvbZS9n9J8cyc73/N3Fkc3JA
TbaYu0ONFc173/D/xwIqWz6fI411+xP/53arsTDeroyURu3kKELZlnz4nSChEG/5KDsr9Rfb7a3t
A0Br4s+BSyNqPRk52QY1OauiQQr7CZjTzNsvpSEjfQS+f7OgthUucIdrYAbsuI97gRJZYu3f7cDd
wJauzDUQkZRYMUAJ7Pjh22jfA98a4y1e65JrRWWUJKn2Ua3C0kNN17W9uT22CSsoTT9iAX8Wg7bA
JwMNFOr4lb2AVwf122SxArI/NYK9GsNaXCEtNjZJKvULGtEB4wuMQgFonru9pKvC/TbB1Hr5vDYW
tdBUMH4c3nKswbsrnk0NEOvqYNx/IN+xiDgY5hP3UATch376rl8gjHtBZo4ZT3pSoiQJgYf4MJ69
1BLB1z5cP7XMbvviogSmc7rDF7f6mh3aTkEvtbJLRrTOUjnkxDxqm1ySoYWktidFWwkOfNecDyQN
g56i7r073D5yWwV6Qmbnaza6hzUvA+puvKzOlVcNHVxQ+vkwO8unAdGMwKusLM5c+R172NO6Whuh
EM23OAG0y/c81WrBiXGpNur8WRECli45PDYFAI8Q4uB6tCqpxOZ2B+bbNQtAyPDYz6cRH+/5oneZ
Shhf0ba8kVRnKA+kMzI6aoHcx6zx72PE7OaC8yIa+/M9v6IAlFrOgdcVraKRmMpwPpZxr3k6VBmc
DJ01d3xkQO3PpSSeCVm1X1V6M1QgAET9k6JLrxwoAWmoPMf89YWyedI3rO5BspsScZD/4M84Shcr
iHlQ+8YDQfUGxvBjbCXgHnSS9lCypuLoAG710r/a3YCtLATyj9Se8hkW41iEFl1q2D9BcXijhw9u
X8rQAJqKjvfjfBlztTll6Kb7LWdxPGAkNST6w8BqpnLSiaFsFtAsZrNQUSiqExbJsx6+BiwnshFk
6J62hE0uftQzszTsFyZj0vXnb9eiElikSYCl7MbU93T1SLILqpfD8s7zNdjim9h4eq8WTVwrvoNn
XVDMfw4UtLgjA7tYd8SMNeP5M4CqLahXPjkOxMQ4z6SiSiKuj3mlUYIQU37hM4RqiXMSLfTHq5K4
9ZLYZTco8rUGwa4XzbuzBL+18qPi4TlIIk3U1E2r/qfftTkxNOd4snrGHaDGjVikf+IvbWfzxwtq
ENbkb4no61CwhEMHplXbxY2Zhpqn4FcfB+zgm9EhW1stXhg/SJK5Np4szERIm3yub74pGCfkwqnP
AN5keEeocCs3JKFN1GCyTEaly29Cvjv5AA68ctgAn9ye1MdcEHVbW1RqC5cA7xL89+htEfFLPjbw
4PKN2baXCpY5kBkBF5WgEzH5iJ7tIamwcbAMnsdNWVo+9/3g0RoSNdhymigfoNGYrDbVQbhs+/Bs
D9gxJh1KT+YbYlLU5v5Ovw6r5NCoFqQAzTWN5ynxixoOPmK0q4taLw75VPRdd8A3XVq59rfG9d5r
RuKkc48sqtiLu8ZUAAM7ap+KizuHewDRCFLMYUXk1LbHOKPe/z/zcaaUTHgS9zV9KAfKAANfh5S3
82LweX6gc9f32pdowjd9i/1kUj61cS/1O/lYnnGoNIqLbuz3qpg7oCdCArnPpkA6x40dCvG7mhnI
UkB5q6VNIti/raQ90a9EwabxCR+p2WxL0zqgy3M8Yl/QLkQ+iWAJZVZR60BWCnQNEDusaf9vNQUj
tcj9v9x2rnknuZF2hOzdD1wZ0nitxwW/jNiwXcZpOuqN5WdxMMj4om23WPr7PxsI103p+4Cz9fDk
8L6CU3DwuUzg9PpJiFRSlbvjqXbFwMdfVQNIGLYRzVZDamL4Sn4vSCAg7fOJaUwVs3TanLR2jKUG
jfvZ0MEmfBujtNNsW57uIFkz2soCOogY0wZMNl4pSkbtMcB4Kkvv/M1rgbPidnHr0pkQgZmVS323
b0mbQKk7MqizWe55hy0rLBRwaCbRD8lXQruTFabSHPI/Vd5Bb42ZoZKfR+SkOR3wMNxQxhtjUAMb
pSQ9/xa5bk6syX7gHdFV6cJx9bvpU0OCa3f3EPXw0l5XwQ2lSEqxwE2JFlLXA8uN47L6rZfQVpZ/
YQ92QwdXI9swMWlZYyWq+fLi7BjXzGA9/MDE3L8Ue5B/DDxKxB+dY2QOMH0906a+euX1CXVTUfzf
JZHTpbt3ClA/TU6HDh+KcZWN3414mwhOZYHvej162sGg5eLsCkPVEvG5HTJAUgosODdpEHoPjaSo
LgPx/NTtwX3bPPdAx6i6KpZshIQWFFKzQXR5VVpEYL8U5tBzzO6qAsrQdUqlWX+1C0m4fqBvSTWV
EgrWc4lk+6Hjw2HfUsMwlPitOsR5rr23i1493HDO0uTn93A01/31HuaS1V9d2d0w9G9QnmoFhKJf
LoS8km16StYiPu44C0GyEu3Up9eoQAuj8Y9jOREGI6xD88TIZGwpJrZnVY0QNHXUO7i+pCD54q1m
4SjBcGrVONZI60D8176+c6jOQq0IgojneHYtLlAxYRe/PZQOqdQ+KU9ifI+/BzvkslYEoBN9Cvqc
6++3V4c1/5KmMj6jEKSGAg1vHMgZZoZCA+HicHBJK3FRDguWsT/rjvw8sC6aYuqqeSLIMemAbij3
9aVtSBGSncHiuuAc4UazeuGtbtWAeMYU3oxZDi0tdhAco26huCu/6Cwx8cJo4qTitVmGTcE8ASSR
Wq1ap5Xo/KuqKGwVrsQzkSRGdDrWwUu0R79XH4LHjYpWETjWUKEeeZQSYNd3gfCxSUq7dNzWljJb
fcgb4UpEffXaroF99FaPgcbKvnUhILW0aQeP31Ak2rJ6tjl+dR9dtNPk7Ay6PMXSO9SHPsbeNFzT
UOZedtxJTDEZKcgDM0Tt5Rvch2/JyNkxZQ1MBbkK1pY4Zg9pMZ6bFTJLOgK4c7bT9mdUR/G8bdIr
b2MCYPgPNGt1a1o2W8BZS/iTQ9lAdfZFyFpqn9WcKyFmtw0M6oCNf4FbChA16huWH55q/OGbpGeY
WQy/Qxu3WnNb8sWgawbOniWHzo20Ug270FUvwgyYps72RJHaonBkaWRV2CfAW0E3IlTtLjBb6JnR
aBnoIrBTpgfxMV/vtuQkh6W0bS6gEJGX+Fk1anfTxyx8ThrTFIJKt1tdNrZEnKr4lEdqsuszv2gP
e8BsFm5THzMqVzWnDShzUgZwFZP+PbE1xNMCFbw/LnaQNHc5w7YRHgI4WYprNlkoZFOgA1qFRAkr
MY/F+/218jS947OYbx3FJoZzN54x0Pqq1JHB6URTrv0NBxwWE7EbhQkOr9hvztMEJBUIjypUa1WX
l6kFf7IDWt+UE2wV2L6w5zAPoNEwFubCXWS6HiMH54Upi2bIfcLC9KCEMq/2C4f8pM8kDSzATFer
fvDHuyF3IuVRdpuZfTLTPO5rs8RUuIgHNahD+1aE+yfTtmKIc1sMS0Vz3aS9cfGwTY+C6ubie/la
1EsCpuZwKF6mNxnF4QoDX5+YYwxdFtAkDri9V3NAd4tgM4mW0JMKDXupVhsxUCboK1rznlixWY8o
A9CN/3v7NnhZgY4xK4qia6wQv/YYJHvTvElZFA9dyN6B6pMfZord4tAT3k9J6i2agYkdzeOoDdLc
DbURKTKkpZdI9zM85j+H8U46c2uug3MWviikGSfy94iy3texOXkDtgd/lsfF6ZnhIVFgExqLS/rR
QSl76Ewpw+GhCsebQhyF3rslW7HTjTytD9Y5caEJCUNlgAmlp2+76+fWMXQ+SQrYw1g5MIhy3pQc
9mRKYHu6lgVwsUSevxzFZIA7joY2a3jUqnDw7GB4yK2IxgfMxM7dL2021FbIrplFxl3My64iwG1U
/80stsmFWet9vFGui7bqpt3H7ztyBxEjYTRN1ymb0uhlmgnG5cUho+XhnRNB3Zn405IDjEJwyysj
+ylKTCQsHo0gHUFzIMjct9WKVlMzgKGb66c2KUv2x5ufdwelUWxYgvn2KJti1Q9WGugEcSq/wzOq
PmZGdDVSZ515PSlF2qkpRE14WSnZnfAhkmZXuhrCmzrM2XMlIQB8cYMfpZ5KgeGKj2ImX3Npx33g
CDh8dzHEMq+0qOJ9EtqNSMhhyIh3NGH56PZw+atLtidqVGVyQ4ZEFLXn87fJpbuHrJk0x8ce276q
tr2VDZvhcKK+dj6MLeveBpdSHo0IgW2LMaPpDjTk0RbroLt4ncQ8iu/P1hHuMu2GvQWedZN0O69C
x48GRlOFVffuTxlW2hu+WKnjr+1XrIyy+YDeWetVQ7U4myBhFW1jfJB/zoyrdhO+lAL4kuQPWN1d
CkgEt3w36g2fm9jXvWC4eEgA1VPJTyamMv0ZxnLN8XQ91rdD2bHVtMeEHHDY8sKwzuWFGspDdpst
x0yWdyMDgt8V+aXXrQ7JxyRfuw2ho14LDWIVCPR2rXUpYWrCC1i0vZEXXDuR3sBNArfi9onfV4k9
EsGjW6O/6dDrvYiX1sD1Xqua2wL4dvpy8U2FFjg3+k4xNXcD3mH7REYstesJGFFjSZ7fAuCbWk+J
2mYMbZDjPAfo3c/z5CCBP0C56Ntp+Ak7P+pWHiHKSHtjvKnEDGRPLf4Nb5oVTYNQCex2Vw83Tgth
DcRhJZvQ8jDrPUnK/MJHq9aX1rTxutEBTU9TMGN/hDLWeb3W68UysPZdiJNN7z8ikQ6wYzVyshod
i3tkRERnBzog+UvMgWqm/bUUZyVJffF4cDUXYvwteAsA1HQFNePTXmvw+GoI1XijLKRDBYoRyu9M
ZJibUDWxJs3LrCTYS+jxy9maAq0JQK2EXXXCMFKeCyNstCQp2SkUYxaj5ggfaosQ81Ph8rdoDaj7
AP6zb59yu9DyvLZTqeWh4/5tce9s81BOIS49Q32m+7JGURX/2LU+ZMyTESxAcDisdy0DZ3z7cuFo
B1kBycPP4uEsVe15sPH1XQFOQOxXXKMHhakAgrWtv1M6/4UwVZfk9TWaEtNBhnPgjRv3akiRd2wJ
KYHHOJuRbvK+I5ciPE8/+Q45K4CcwlRtR5J8VD9k/r1d+urnTLzCJdNhf3wRnMjou9RgrZZY9tjI
mlceOex/LD1kT+jldNUMyZX0y5ve3w9REZTKwbWdppFvs2uqPgcF/7WFFgETzAph9eiYkRYWBSzX
5mdGQb7oJx/w5xWVaU+wu4Vk2ri7zuaBOwpMvFT9oFA/viWqvPrQlaaydhhaaIvabrGKyAJ/ha8U
qNrUyvkgltC8ZBp3MioGQrqQKYOftAuIaTqnZ3QV484d4/F9n+q+ZGtDd4evM1wI1cehy6JEt+Zs
0wrYrAth2A2po5B1wtaVcNpEIIJb9qKxJXCK7bTcDaCBc08Or6GtC1n2URtfkcIfHpDw08LVrV+5
NHRoBA4QwFKby40te5hmZGBUFWt2z25ame+mC0lL2N8btBy33vNooxebM11szygyURfrBF/X2xZh
hBBwhGNYbNLA/DDkP5Atj/efGD33TRqnvEhlZrXgm3oBXdJ8tR1l7CWKtILR6SFXM/gbXugMaY1t
cWjkGspl+Xtc5Na8D9M/XJkdHVnCvx6ywht68UWMKASJOUdgCWFtxPtjgZB/1NxCfamNxsBcMbk8
/qp/xctpDqiL+6a9UYQ7CcGWusTHGEVPPCkEE+1TSZMl81OTdVCOpNIk50+cAEHZ63WcxrMUmNTV
rXQ7mNEHYL+5tGExE9WeG8tOU14rsWvRfFywvgwmmCJyM1eMvkftQHcI2c5J0PVz+5BMRmkBVpLx
/DdfAooq4Emos0D199yYNvU6HPv1l/2MaOshAt0YDJ15HplxiofEh949MuQvwSgpO6P9Y9IYuiyg
7Q6qPeCUvrlddE6MXBxnPiMtpNcrgPvv5AuuL+pQwhndUb5TIUVvWhL2ZZZ4NqiCEcA+8MbxtPAL
8K78Dn1s44cCb9wQKaB5VEIGrb9XKa+8v0YVu583fTqUSBYWGGLhytlei7+bgoYWCWEnQBpV182e
/uZOhq/L5kcWLFI0no5dKt9EtvZ3cFAcBeHG1slCmISVgNrjOi/K7d2ZmjPQ5NOFZXeRPRrBSNQo
GOxHsBIyXv3jAf2Cje3qINaSI3HHrigE53FaKl+zD6NfGRjdA3XoIUY0mqZawtZo+suvwI5FLAbR
Gg6tRTcK+BLIzs5szAIfeyCMjmtqBKqngHx0bRFJOmkpbnpJEyoILGTYodviAW2z6DvT0Xo/A2D3
34TAkvIL7/JF4Qw16IxMMU3IApSxPvNBhkW0JljMTQ6UuP6wh9wfZEfzK18lK3H5KCx7H56tvzKC
uElBsgx4XlCT1ZaUODcVspjOoDbbiSWx7mIwOzlGejpQzGxrWP4Oik8ub80dwfB2EPndS6glRRiu
HeAFH107tOMawwuQNpAlE7hTuZ2gs+dI47lTfIiMgQ7J4lI49/tsMpn3i99tw7X3D2BLMpMXauAh
5E4ltdkhLi38ytThURZv02loH+6J4kfeOjMtJg5U9rDcidMG/k1EptBwSRv+uFATksfgFIBPWHjU
2QWSX3a1VyK6lQOUZ0QxMqUejxJv8vMoMfpINo05SX0ohN2KZPhvUL3a3eb8kqLDaJsHK+LfwkQ4
4Dc1wr5OZx9qUu2fd5uSEo9AlB4tPzwKdMOBzHJrqUO1AD1RdeYhN3fkKicGtzVAFt2YgiFlOgCj
49QVB5mXn7FNAob5MQvuqrP20E3cqQiqaU2Oyrj6MaMm+WtFvw5nwybeIqEdxrB9BEiR3X29Muaj
IRX6K8P/Emiq6VR9hJKC2DBQqtejtN8LZcMH+Xhbm/YJ0NHGuWAPYQ5EiAKNSA9GoB/NJCFA45Hr
ff2e69LncxvOoQYwb8V6wKgCSha73YX4V4M15OmNEYt1RnXU8kL5CT3gyiryTKxcHRdQb9uL3BHE
JuEP+8BiOhDUalCFDcQnOn4KZyy63L/Wd05GAuX3p6/FSPwrStAjNz6EWTA46NiZq8UTAlEWO/hI
+OoXjDFcN0SEKFH7C5n5vOdjxQb5o30F3bOXCVJLcHBGVidEfDVBlVs3qvQ3S2U9uGJ91k2GPnzK
6PNdc1Z8F1QlOYe17dNGDATXSImKwB1TFebXp6+uX9f0FF8/pCAVZdYz/N7Kjk0UcZgjAaemrf/+
sD/5iQZnmr9qt/nol3LvXVQVfqJSWFcltbF1Bqzz/UXvz2F76WXjkOaF3XR8lQadK0FgU64kanYS
/9DKLb9MxO0BpmZwayUi9KGTWwdIWaQK6zQm1/piEpAm0RCBPIsL4I34m0M5HOLo/jXyJv7TSwKV
dFDa2WuNvrDleqe5uUPD9IGW8yFYuK3g+XOeNRQ05zXieDzk7HOheinDejR+Z2IXBc5IUU9+WIVy
q/Yqtt0YgmHc4rqc3PPJK1o0Z8pmguRh8HNh7Vtcm3MdSr6wWKTBSLGj6rmRU/bHJwTbpj4fDl1i
6X3LR+sCRvJTSO0e2Kc+CiPOf58XPsqVlWnUt8DMYNlNBFeqIgV2cTTSJAycq78Q1U5gKzp3E6Ix
lfRvichsmhh3mpxDyCOAFHZqCYHj9I4v0/34TzwUJMm/w3xdc9jljox1cH0szsW4xmKAOQZUZiiF
sw8Sz/zW7/wQ5P3O+ZNA+OY3aKNqLm0vb/Ty1fEuk7G29q0ZDxJVRQBA+MzoAcjWVnCpNfG5ldWL
ojQzi8wvYkNwRDMQVjzGYfw9rxLCy7ejlap2iZtAfz8Ov0rIW7KhsAV4q4DDQGi7KiKDkiB1/+rW
W6yMvFpxJpGHLQFq/3/F4Z4a5AzqEozrAgBleZKAmIgf0lFKiGwWpyRx/K+hTHKmelnx13vBBPN6
/vTDopciSy6J0vZg5Av943cw73R1u54mPgBY2HndivQEujqdkGjIZOp0O2EkArNPeCnRrnfFmvEQ
xFlNvMWj5C2YdfkSi5Ae/vkXjzrgpH/bkmdf+ymvNqmSzEzwi2p/NaSmlULc0gdj9/VsSTAFTOS5
uUPEYqt8raAEjpVgwtYa/YNQaOYtvXNHhzLhBSKnEQV2yR3RUpALL4S88ry5xnggOLCxDVASzLfy
0LVRL9zQsd8iAgop7qbo0+r8QVT8HoyvYhc5XbARwlPLBYw8r0SrkYHJn4uk6rvrCfxoi4jFCi0+
XlYuC9EG7Ydg1KdKeQWMCAYAeC8l8JyqUFsODjaLNQ00JYnCjl4I90hBr2/GXapw9mKO6IC3ultV
QwDgL2ehnIRbzqgdcl+GZS97+/7DgEP+y06ZuJtLfppeoy8QRG+lr3PM5hXGdxx33+gCr3/NOixV
w9MS//5M7Pvsysb04I9tIN0QuxXRdUVGt7qGYnrJB8APtW5L/ZwMoebTbnHspKt3BedsKZFqaJLE
f+j/7h/Ui/xdDvQs0ROXxR+2wx42fWagkSy07xIQHxPOAUGv4hTlG9i0z6+NbR8KF1S7g5For1g/
b+n3or2soBODknU1pCLGnRVu7LpTrMs2P2sGCk2y30dYmJP3VLnofRekePGeYqVK84/Zox+iFlk6
kU8c44H3TUFYXU+wgq03Ab2HNdrvA5R9uQfrnH4K7LEnZvPQckQtnKTLr7J+rvJcipsWhwvIPdsR
heX0x7oZwvdfU5SSXEaWfR7qSuQSeNsYvhBTCF4bkL3fyBhEfqfOnluJ+43du8YCN990Y6K9HT7U
JkZSzOBTGg3KuMjg2kU8XpQaG1A14kwxXWlm7sshrcPXKYji/le39dupJUIDbcw4kv2A1PG+2Tms
lb9y7n0EGTJqyLcmZFTIq8f830UHNJDMDreXa+V6LBBQgQtExhSRFh/J4GbH+trRftAE5onSV8xW
SZ7/KGdYJoS+p4RG4rlBo+ZVQIDJUeG9CYvl2Hvq76XjEHapV3oF4MKCzqdyenXHpvtTIOUEI9TV
z4EtG8d8cJHK1rnApkxxnClC7jg8dQL4exBtgoRu0VfI9KjZQXItnwxjkpxx5tIXlsxU8T8Gzjrm
VYKA7pWd7KpOCacKkdyBTx2JCshQML3FduPkCOGXPboG17rvQg/ezMtNFkk3xZMHg15BxwUCkYJJ
+P5BRkWDMmMG9iQLq2+e/uSlCZDCX5iZIwNrSE3zZipZgDCS3JDAlPYhY3FlzJRDZSPTjNn1TW8c
0OoFkwFJWoBVEJOOfr9+2+Iv2spzOYS4VmrAQtyXeV7BLeLQwBAiPyskiCh4HwGrC559q15jSDdM
GUYbubjrH4xUCDZzBiTxK+DWdFyGx7hSQxPIAaxJl5Z8G4QyG7t/u/EOiWhxwbNTHYzkLYK5RjfN
1slMt25mJ++SUuLzZF5WCGZn69eGwMWCkjDe5ySNXeR80P8PMJDwD+t0Yvptzcuphx8cSI2eS3Ch
/9b5cAy7fIlSEqjNFaRZw9PMghqxCHRV7s+jnNQmwX/cY3hAI+P8umMd6cIxY85i3Xjt5BezDh9w
ZVxu1IFwb51LuaOOyILAteKjNEkcyqOYHBRg0miuBvtRJUef+9yiChxXcTx4omeQR5Uhp5mADzo3
UMTN/QT56x+WGGFKzSN94/k+rWam87qCU+j19zWvQisZBhL7cEp30L/82EcC0ychMhfL3T1ifE6l
50qe1fiaS9OuO0mH8PcjQz97Uy5E7L48HRTCjTPNQzzeJTiOD/SakEE1ev8IyxMgATPDTHvY36fi
B1GbsHkZZH+KxMKPgSc+IPTxOpQMTt30UKrnXSamUMao5ptzyFu9cKnBf21BJm2DEpuGCVDk6Kol
J5PH+rdBM+FzeYoLtaXXWUkLa0FoAk4CVYD+dpfQNa5Y7MWH05bgnDHiqWvo2SfOXNGkS6kY0COC
6XKyAP/8IhqUsSkSjCbDd9CyjsVX+9fOYYozh7lRm+AKpOFcmgX4SappfVDHI7DeKfTJXbnZUNzy
OhY0k8WRQZ9QhM5zel1jEZLBU0LMWS73wYJgCZY3Zsn3c85JAsDL8ZllRuEi9kMN21UntQTZBKoO
XWBcEfNRaPJskf/53xic4YnfO/d3BdtKqLXLL8S6Hh1DR29snqav761cj4AGtILjaViCaFi/jWkX
BPhBkNLQkE13z6ewv+BdmEK7c6gm5ia8ejAj65IombtULMtXgIpgL/6I/Is91zlLRqZYMpAmPP6A
9T+iYN0oyOLWXVL9VJ9MTNiLa8nf3ZqJ7DG1JIu0sgplEB05xCKNWrIvB+7l+3LnIzOoAqkbjYl5
LIpOrtjSNM13dpBFyolg5JcHCe50amY8ERf9zys+XXvqtlnc01VkaSJf74Nb8ThMGnR4/tqLGumo
qkW9nLnBfLZ3VvLjK3DLrMoIQVMHruPiun5lyHs/ZcDZv1uHl/dAaYv3Ifx66ya+sBJflIY9SAso
4pyC85eFB3xTlnByD3Ua8QGLrfVMTI1ok6v5R00ssKn+wMDoQn00XJ1zWloro21TzSGBiF+dRIZj
rQnDW9000t888ELlzvRi8DfhtzG33tWdh27eniZnaQzXJDVvdd1e+JQHSFo8SPmPRCBTz9B0Mw61
Jk2sT6mUNkA8xK4+DNKyUDdWyE4jm1Bk8aHBSdWximQRTxk9r0aVvYlZM6CbJ+VqYxJ1lD1dKMPo
qCufcV37MeyCE9tiV1r7fGX/43YUlshWa3yvf4hoApR/83hvj0sjS2G97rm1SoCZ03S66vqcufEF
lrRsUrKcQLcQKxXtmyNZAszTpNuNQVdChgKoOBtxDNZRM+YwJXmSAyJDQL1TElHfbwb+J6XbBz0s
gxBqtaQCoG7FB2wVSy1LNK9WgkYGFBKDun117FqGrGMUlTyA/VbKrhv+JHb47D2EK/T0AzqVsPqR
8vmWkfeo77ypwwbz/m9QPfw/UqP40QHZ1WM9LyEqQfXhmdGYqQlhVPTyW02Vfa8xfoygXW4T1DOB
QI3RilO6mY0fXKOZH0nm+tTOlJOEj8zfsk4dU2adZAZOmYeEpmejWHc8P4e7QgOE5KVbPz584Djx
CMzflQ3l0m4RpdLO3crUsH2wrSJUti6uXfye3dJs9Pk2Hy4Ha7BhvZeC39ZGEsXrqohCC+skMMxB
nNu0vUpcQZapKPPYRJ64B6PRa+E8AQS0yE3sqWVjaRor18S2ww65jw7ne6ZZfOKuP99crp8oilTN
2T/64wcqoTtXeEz6yFnvmXIwiHZJMI0+zF7/YLCn24d63XrPZtOie131HOb6WsEbRScXEJtE+B/9
9NegFb27607AmLC5Zc8AglYgrixmFp5FKAFpZVAmdWWIdtRpgfce/MNPWnU1bYRvhTif5ZSuj/7w
CkZP1AbQWpSmw/IfUIEM7jKjEn529eoPiVQLws7Pxex9pB+ZDnzIrSs0u2bR5skcFhqjMKFyJQGg
LP0JmX5+DdALUpbOudZ1J2pLbhbBL8QtPwN4AgwyocWx0OoiHyUkbs0O8RXwmJnSFXGfBItUyHCb
toBD6K3XZ7egiwzhuceLnmYEW1KwN5SfRElXBaIMqFyqWYfpEnu8h6fK9AzoxqRPOpD2Q5deviJ8
TzxPo//qMv6mgqIAF1/fur6CPfuvv8mnVM9hWEUFIublMFyFhKUFRphV96c34C39zkNQGPWwsWoO
szQbZC9mvw9EEHUOvyCJnr/uATRizapI3VPgmnSFXRELIcFeVQQk0c2mdjhqVTvHBTcJdpsDffYS
tfLFqvZuo6XpWjF6xlRlHjKqfWxczq6+U4F5UpR2b5fB/gyiq4JO+CXrIb/h5qgQsklnLJtom/JU
btaNj7p2i4phhbSn9c8c2b2/TxFm0CwYaPDwEAP0ISOCKyBbU6bjIK7d6kLWAfpk0f2w1Ih4xIV+
Hd5p1UDm0QVxkM6ju+yaK7gZc1BD0aeA4UvBYV+fGAJ2vf14+BctUr/xnZaBCSN2hKlh/oaYvb7+
Rlxp9Bn/hofCsMdI2oSTKqW7EEsTigUcA87BuKXwU8WmbcPgCPNcH9uF22ruP8Uv/xVlrHmlYP0y
BctzAevCf0fglJ6xIn27dyc37Udh7QrOOmiYM1gkCeNLGJal7gaM4lKq+4uw31CURD/CHZ0cVTyo
/A/MazUl7h1ggJCALeCVBWt1Vcmh2f7sdAo8umOE/9Pd1QYV3yqNT0tZcdU6WA8HUx6q6k+zhi+F
tvCDWhrLjo0JOGxs95hYVshI4NBhJcOnocDP921Gn0+EM7gPdZG9dSuzJfZ1Y5TfrwMKqvgPYQKe
9Z9+w68Hosmk5hCQIUxMU6S0HgOeLmtDqQApiPCt3Tgd+YsTzNokU1ChkrSZTq1k2HI1ViEjrK2s
zFzVFtdYf0mAQuXdwxke+gWxXUbhsK8D09jJ2qX/Tbgo1mYC6vvcIwYGfNl4EjAUP8lqQ0Y4NwzZ
kASc1kl4or24Yr1sn9+f3MQM5+CY6kngs6Jw6RxkOcWWMzsksJMGu2DQfCIzNUl47zgwmrQmBkzy
toJzk+wtjYQ+JxYhZ7fiWA0lXCvyho7ObQQK4IydtKLV4cgSCFen/vSDqDsBLjFaGKe1e5ydU6ak
ptVjR77BX9sNtkU+H8ZYOJaAZc+GogcPaJIkLfFzpC6s4w4z8lgiEefLDmcs8O8et2OKl6CcKOf+
JqOMY9c8lwP+If38xm0aCePlnEqbNMgsRU1lkRhfGFYl1nuAC6FJiu/Za/0kHmUD+8ytIvyExW1c
1OL8OJ2WKK04vqAk/dwqV1Btwf2Vs+XMiXqR7dMe3ZImTRCgB5L71ehPKphQw4bbsyyMCh2qBivY
WruAyyuAeuIMvTHbGWMAZvkK2Xbq8J9YBsfWUWvUlhcPpre5aCGaDjnxQZ5JQSZlkC5cE7TTIhSt
0IkIPwthT9iHHzuKD2Tm5PmAXJ9H+FevsPEcnMubtXCMxhTzJc5O5lwkrN9xxjdMf9mtCudnbMOQ
kjCqJTG8LtFhHhCbgPZZIje+LRxFc3fETzOHJeEJLtfp1jrLZuRrGqE3/98EDOOWfibrFXT90ewQ
xz2EC9fxT+pv9FRwsdTWwuKNJt5N8JQn9ymv1GQ4uPLmgJpGHlvhEVNjS6ZOVIqDBz+UdiRjIEHo
7q7klN7lVLUvQdo5h9OeQLbDC0F0TegCKp1ijrgIm7fS4lBvsmtKxR7sIGINc2dJKyE3sd4AdS9g
mzBVC58x+TAyGqpSJP1fNC5dCL9Y+WDtfHwMa+nCkpo7dQGXBETiih5FllWW9++g1Rr84B2Hdfl9
mPqIoA7jFwz3kQOuDbZBgdG6PlKA4vyvC8OcWwmgrkNuaHfSoU2BVkCTzxFzwQdfsKe0C3IDKCTY
oNdM+EfB64TLtT4uU94NSgn85q5GuV3nReFXbdi6jklzs4g0dFLQg3SoWbv6ywDG/geIiwRUL0VF
dFXlX43sVSwMcKBLXivmo2VbMGrNJ2gP4qzukDlfTqqXvLsdAK3PKOiHjGSFZisEZH8EU1FxPFiZ
msk4PrmdrTO9DXJf4xdc4t6LhqlpMLknxR8GJ1z1B6JekR7ch+OJRIh8EYF8IgXS/ER+TZrKGk+R
A0noO6WeKdRW8Fkg8XNhdM7VOPyIGQkfmckOOVoC3ar/8vXKenP8W/aJRcDvxowhNONPyRmS4J3P
ZwaloTR7FvFATCSjfKzCZMH9pfkKY6hJdt7ZMdYcR0Tpek261MFJyq6hbzfkVXb3daGxPRG7d3AE
ptpm+YqhFQ7mrjp98zmxQVMGNnRBIEBPX/vXRvgfcylyq9g+hq4A0PqSfdFuA6BQb2wuWKSZ0xgE
SVQ8UECXSKG4ZjZxLnpQBHZ4Ikt9fGgajl+1WruAq//aR35+iZjkZAxBPFI+Oe3V8DYz5uG7RaRU
DqOkQ6ccWD4ss/kylcDotNI0FMT7dD5+debPqtdS5xpOKB/ag456fpkOVwaDhHtTgn1qQtadAtOi
yuqhWASor3n6XS8bYorN1SLtil7vOwAG+hnraP2ySKTVVztUWel9t8H4/LA3S1JveUa8EsiT1a0/
q4Gc6dBpnUMdMQEsuFWjXmSziO1yH22vyAw+aNk1G4JJsmslVbaqkqmrIcY8XV966EirtPDGZQnn
7swmYoqiOiTZWSxngxmc9kfZEKtP7NtLDmLlQE6ve92bbk16oXYrd2a6+fddLb7b+fTqrJWcz0xZ
MAZUvUPzL9D3mcqqc4wyGeK8osLVpE7wFkZVVYOxExPZRQmh7poKhJRIZfN5AAzj2RLPG46jJEVp
XdFgZ8Qd9KUf52YwBJq1iRnmvD0Y2QonGbnNS16OAMK9510TE80Q/g0xyf6c83gsQZHf5h8XEPIX
reZdcVBf/qzwsIHtGImV+j3hekIrwoTNseV/cccj6HThwiAO0oUWbt3qV0aibI8dQi0TOys1K3/k
C40GPDsbJZ158e5d7pMVHC3FNvqXFsDf7zA2A9TpbSQkBpdeVACS4vhrUVqNMgcVOd8ltnsYU9cV
U0ul/labOBXSDDv15koff1DM9HWukxpEFovfmJiSBceE5d+mCGvKCOLtI47zfg2SDqdsF7mHHzrA
VbCytIVHPhoc81hJOLDs76rHpQj36m11yeOexlVJCmDIrCn2VQ1pFGwAPQ9vFN1qwnRLX64tqZ3j
pGsCtT3Tcf3POg9VEvE0dFcVV7X5E/KNvB1PaLP4fsijn1R/JyDwgEDJWih3zWjYp8P7/d3+9DAe
Glf+N1JcwJt5wxsVNt/bZCWrkpEwAglesadTuUEJZP2tqrx+5vzdlCcHPOK80wN2ZtM/oQEEi0Ou
AtURY1zOnOPyfkJv2q3nsrHJU6gh6ZhAM0+FsiXuIXqj7AkZRQONYM4oCuOBsrirdnlTyc9Bm6qs
gaP03NzqIVdkPZ5toMwVSSE3Ueq4oO8C9kjlvEjjXIB+tF2GTknpqwoLTaYClZ+DOVFwmhrMGAvh
KBVI+Y4RC3s6WiXGfFlQC6H/kzYaLwDlQ+5dPx+97Lps4T5KwUt2IaDOS00y3crjv6T3H6KMjYe/
pGY9ATR8NvO5KBF9lT9/aydHXul5/bkhrlOneg65RrwOqVOET2CQSS7Sdom1nZHG2cTMgi1/BsBq
Y85L59pZ9r3FitxX7MS2STayxzg9tq8VWla017HNeuB+L8udhuFMYLHUz0N57iyHQfrIJNiC52ZJ
auFg0m5ks6mFun/CpQrPW8sA1gALHVnTSWWMAYSzogkxQRfFT2FkqEJloMmGT+lUEBWrqKE01gi6
UXYvRUSCqKmHmnpxXEDk0jkYff0ntAhj+CstbNE6I2kAJ8Q//Yjgxf/MmaXjbdN4xXouRZZxufy7
3CoiHXJVX5JhPOFu6WRIDfSKfJv/T4Sgo4rTuAc2KDo6bRWArBqHsJVl8EVMOZn2dGUARuN5FeW0
0y4kJKAAeh0aozSOnsDpbx6krq1xy02nS9T3RGBTzHAZb1JnWgRTj/vCjvlegGdUxV2s4z+dj4kF
/81wpx83EhDHOVZwP7GzC8fvgI4FW7SV0gF9EDVkWHH8QNhIfHpzD/Be9mdS/qKwIA0Ra8mOipYk
PPXKG+8zC2wsKyUiep7DE0bRFKRSt9HY/kexCkxfKbwlyaSqt1EuicJ1VvKsGFGsClq/1oMRgQnb
P9g3q3bg+1P/cVroDmSwYcs7ggONbpqgKUaBckrGzLmbkvpN+4OkEtfEKxmasnz9oDfzaAdvOarK
v10/0lqpc8mSuEhb+Z/fMDJz6/1Cd27R6nn3S4quWnURnJi3kjdAApGbZ8RwFmmmcdL6RDGcx7tc
SFGNT33jgbzJfr13QWUutnTEcjXMxJTuqPHCmdiF1ZiszQyEKtSPz0gnSwM1gPckEkFR9hr7qUhg
pxQRNPMqYMs1IoHW5sEtYTPnVFntuJXO07TJIfcUVNVg6en/t1mB23VPc4fEehedJG9MJgfdnCHU
7uAioitw6VlZM8P9c5xOROVgicfVCaXL7Jduxq21s1OtUbu100YAV0W3DB0u308iclKvoCXzz9p7
TSP7qt7BhbLsqsN48ZmB+ftpjtW2FvZPnKv+J7t7spPyaqRWzSimNFjVa7s2OM6PA4fXQOZASxMb
RKmfzR6ylMYcYEqaTTjPATPjp6RLplFnTBy9woZyq3GM94WXQDhzTUyDYrISrtRu7oFxUMi2qo+k
3U/GIVZxwmeZN4EMxQ1jWCrVmt5tT2p8b5cnSKLhIttSiiY1ubnXfpOR7gUr6kOPa4txG9Lm+nYr
zBUJi8ET0ebzqTCIzk2Bru5vaT44/iQ45W/E1NgEUhs+02Qa0IVHAwSokYkQvV4IQjMzG4lhjlRr
QDLRlNfTnQHGG5Ktl8u2Ze5jmy5Qnw44HJY7tX71AAT4MoEU8PYHOM0KGr0A+GPKPgCBW3gqgeP2
URrq2Pegca6v5I8woZNTJNawzjG0gEUbeKiOuQJlbyV9RGlOLn8sQ1cEKQgOAz0l7CoOotYoPvCq
duNgeiNOZgu4+dhH8NDWnJFdxe2A8gMhTYKuKeNjfbiHkAd4FfnG2oyNBxrA1Y7/DhHN4TSfVDfp
g5b1qzPx6QxnXog1f1rB+LI/5PMfsNUq0jJfHx4Gznp3IiHh+W59CyMrxoXQAbgfC1tjU4RMd96+
5CmyjeLdB4N0iM4vI6UFTZNrN8wB12GyXugKLOpRIWOEoI9TqKUW/jVsl5oA6DsbTOZ13bJwkH1s
//RNbaCgsyKUox1V+fy+YZXUPKLy7a2ss4L/F3y/0/DmTSLNqmfYoXp4Gw31LF4ZybVGsFTSJV7L
HgG2exDMOizBoGNfPdiF0OSaFyyzmr6MyTpfHG9AWk3HMmim44C0mpILilSlEgmOyqYfwIx8pLgk
DjzI5GtFfgB+laeDMe6HoZuUnnQpjeVYgRvSE6ku6Iy2j7TR8nSAKSZxGyRY3S8+Zy6+pJ1gM8Wi
w6MsFhh2gEh6+t8ENEIDx85voLdaleUGxTc+/htrYt2ng7U7nMXQgexvvnSKBt1LnvFSX7I3Wz0K
JPu2QHZqpG/3tdBFDfxKMmd2CcXiFKKgNDgSQS1t1SzYlzEzzTHRx92jR+C35ogUXJCGSiyehiO3
wNxIrdUpQKaUk/mOg/tzzVGYtIwO4PJ6AEyZu9j28w4keG7n6emB/a+Wa5ud0dwogjkjCwEnvzP/
yv/REpo2I0wHyWjpse3zQAt6UVT5iTUi0Rlza0T0m93JrYB9e4kF+hUzqO99pSo48/q4Opc8XXQE
wy8GAYgu2N0rb434KfrINERBsYqQCvTGvRkCRwBMl7SLDTYDtJjsYcwxVqBg8VzHSh2AwXeyM809
ORyZn4sU0kyb7cTQjIq7PaxHstR16mxJgXfQqApMdqHaEPZ3Xf1dEfL/HjXBTHoW8d+TsWbu16rU
sVFB1FrctYMc5OHovixVlMqjJMlszT0kulOVs7Py+JtwMh888LLmmaEbPczWmjhv4Upgf9ZAu+5U
X/z+0H+gTzCx2/glHqwccnNee0FZk89rNG1PKV4SzATeuXIjwC/6y3t0SQFRColcVamjse3B6oYR
1ce2ZNnMfJVrSzoLmeLJf5lMsrNxyYfbSRtUtnxAfrxgE9bL9UVbt4aRvlyHUH4M13gVciOgt7WV
Ulq3U15xNfCV2Bv9BmYyL12rDso3s8fhGiMFzX8aJTk9mNuwiK7aoP3WOp4JX4Z7A6lxQiNJzfNx
l+8DNbJ5+MwExgNDhounF7JXrgxzW4Z2o7lfSPQjZEXmGx9RrFZaakzQWxJRLvjf8/jYM5rwC8Tx
UmtXNJHSS9T86pco8wlImNf3/UxKlDZXZUvlh5nhLCgVMz9GiJ6B1i6kZyeOV1snOo2Zk6UuOIBM
lukb/v6jK6K1Yx1WSfcw/t0g+PcAHqLerKA3abI4Zew9UYB5OSe96BYwmxCFzv2fVJEoTVLBxg2R
vAQM7mxzquiJAczxOPKkAwToXRu/ZNZBWxnYtakVdSMZ5R2YcTn1JAfO8qythgZ1zE+Hfz0kzcLq
KfvKaLEh/bLM99CSzRs70IUhZmAGfaFfxY1Wiux3k/55QCYlW3slBqNE0qv8yGam1I5/ms1WDKWT
fAppGgNDfJFFh2ad6KZ5S8TW/qZ5Fl4xLZHnK4/z67CdKWPKBh26GCE6xbrM1YwwT9sUJnSYMN22
DAX9JqYMSOmwLZIUKHxDMYc+yaMOeHZnAWicufRdGmUUNBvGjXKp7vRc0qx0EJeebVQHjooX6lb7
jlFYHvcRF5z9cfbeeFFNFEivVsp90xliD0W2xRhSetuS6eg8f1XTP40NoyFY6JXd8pAqHs6gsRGb
wweSl04O2d1+/NfV1/g7S0e1JEoyJgFh5VM5AAHgV8rjlBYt4BAlfqVjCT7zxbflY4PC0n4CVpRI
di87F23GqQX2Q3Otbc9lyS3hcD1IDSelklNnU7aD5XDnn1E9h10PT9jRaqzArVPgTXcvg2CWh0Si
gqWZwU+1ulGQ5jrgI6/Cv2XPN8l6hEYOFLj63atkYU7uDgOkyiRQ55/iXb/q3SbS9e+SZV4zkO4R
rLVXqE1bKu1TiL19qr9oetW8T2Fs54Q+H2wusTqx6BjVRdWDQXMVZfi+CW8csGNddZgk6F2sPBMc
UXQ5G/jdWce0BAaOCnqMzgoWHNkwLbNNK3kJxmKJPuDti6ixNz6szDmnZTQJIm2Q1ZvGom/jxTc8
lV6Km9z0KW4d7ux05SNgoNOH//JrjDrYJKsgLhXeLpcCtr3T2e/2+kuYNPjebSd1CbuAaOXMy+lg
E9Gj1xampgCg4XDls1yw2uOZXfkoWItCWKnpC+sPBrgATD+MCX1+oTBB+EiIMb1EqJE803CMZz/8
q4oNOEd6tEC+O5Ra0SjPzPZkY//Oe5gjSZV++tkhb2skG0qzGgHTo3sT29IeIdh61TNX7j0jb7pQ
F4Kfogagx/9c4S8iSUJpfAnaEUPY6qEgldTRycXGlWbmjJSUng3kG5Ol49vCdAv8Bq8G16/3MwVE
EQRoPzfchSuIdUTcmMfTa2+aPvoVLwFOs7gB4UoXQqRQ+gY8PiUzmFLcrp9gxMdwXDfRqVYpwyU7
8Q6IXes5RdPsq6p9pux3kaW6SUDneetKXuFAQ34+vT2S0BWv+p7P/fcJo8xxcPWPQR8KjVTUuQtE
Y9NM5g9h44Xqf6sqo3Q4tLTGIy4YUzQcaY2l96Uy8aZZLQ8hhCrgRnmQ4osAQ1QWD2QfFGx2Zody
1mBAKg3O6InbzFi3tiYsiZxvhifMQBGANK3Rd6nyB8GKSYHCU7FNb94LAe+Oy6YNnbJ6wvPLnC4j
152f0SQIQ8FtxG48TxITsW7n6ys9zehLfbZP2+mlQrdbU7sdzWovKv0WLAaKF+vgMPm+Oda1DI5s
QzkONr6QCSkcw04p18PTbCd0ovj8lelKLXdHV+zlj0cPmHOL9MmEbSYs3o7SPvPkI5sUxi0e9a6a
XzmyQq27f08B1QlTP8Us87WT0q47p6Zvuv8xevxkPjO38/OnBV6HLgJHuAzfKNUQ5yTocwcEvNQr
MRp2RAEkQTbWRTBL9+SqyZWaqyQrrNAEdWAtFpe+kFPwucVz3+M8iHFjDqMaj3pEl3voRCAg4cib
3DRZRQM8g+d2W3O0shTnn89TRpLx+2kSw5PZuDK7lA86mLyBRTfuz70nrfBPnf5paN5onukU31PH
rl4HErfIHnnP0mkIYy5cbO90b/gUHwB24AdqH18aE2CN7kCZdlJjFDIiqDRC36tUP/S8h/E27NR7
hmZjkBDXUiA9H0ON13TSn0TmdGkLdclIUnkt0+ey6G0UVeMtk6k1PsIiegBhvBWuZ+g6ORA4vLRb
DNCJ5x/brhTi25K+MGujWM7Gm9njJxCiJ2CqBFPV1N73HKU3FVJEcrkO8KkWCtJ+1huVdcg1wnhG
R+8rBdvcXQUcvxWX+gb8dXp2RD+AktpEF92izRgQZo3uyIZVhcqBrvWsShhnpVW47A4PiU8SGlxn
YqWINxlNVh3FG525k7P8Fj/SuB0CJ7djX+bEZcpKt7me899MrAPag6jC94/qW+rrtA2N/MbFiysD
ybD+Nrdxb+r20FFOgpjKqV393vtwwyX/I7DqkjMgyWuU5VbPHDL+Vw9M1qMQ5uR4vcIVbrlJjeAu
y96Yc2nFWjy3sqNOkLp5GOE3LApyHz7p++FoE0umHMKxzQKQt+57MfSzPWb/sef7PY0e9KMVRzqX
iUkLQ4M5AKHpaL2mfNPwVtou3073PgQwJ/aJ4dewN/Zn4t/A7R2+Y+fDRA9jmknwMijLCYNCrSbQ
lnAWUmY4ScZqtVv+5nld5NxFFLjv0OBygE1f9uuP7Y/dhd6lIxWkyg6LrvgWeAJsoQLYNwQBVdJ0
GaNB/WIgkp4ByShdujZ/tpzZA1f6K1WCv6BdQGpHIkb9szlfOljqQi2zv+G/LY4W08ucMeayrP7H
oL9qH0yZW9eszu4IyJEFikK+cgjupNetzz/FXv2+zN6mbq1uEPwHpK3KzTyvGGB1liE2Yqi+BrM0
sYakVH/aa7i0iPEzWKBS1vGhKNkjjjOTofCcsvg+H+9bBccMrQkBoV/tbycP20l2PCSODtB26amX
M56YnGAx6/Hkq6bTkMJq5AH5ZhwYO51x5CpAAzCDMomBWmoL6Q3FxznZBzeNshEOsVaKYVBDAlLL
L9ZMMN+eR5XAqBPNWpBbdXDPJYGXXi+dtysMSenC+meUHMSnKNZdGlkY/AtWjA7sCvCYjweLfQzR
7X+2SmgMLp+M68UMngy/klLqzHqruZmk3fvpL0yU4Uzr3sRagOar1MGcBv5j82ItIXyx+TZYjzHa
ewHUgCDraCKQzIuqfDdRjqBcFjdE2k1Krix13teO6g5gVZ3Cr47AdBudyinjlPKXbYmEdn3aSUlO
IjRsecu+tNqf4lXFgXn0/KBX6AziBqtVqy7DlvFGerWH7/qRChF0oQcC3JULLGa47G4CWN9hihXu
CCqJbF48KNbotpmEKrnqjFL+mIX+pWCg5oXGQFdvSOfo+UBIZxC8OnXZspTOwIJtYCDtOOCuVaSD
y0/91k4FwxV8nDAV9qPEmD4X7EKT2DLzQO3M0XYLobVGRcHyXYkt+nU4vPfSRsm9q4jXgvVWtJ9K
6Br9tG4ta5UniN6wG8C7emsz2a1sjk7j6S98uPDHC7j0leZTYEFFLYKNEfbYmvBH0st7k1forzRd
WFXxCmJpzVTsoJ0xuD93xicOhsnWe2AH2QOu3Gp9cx1poBXxmo5j/nXG2J/SNZc2DYul/AfFX8tf
qLtDbcYdygPdwd9S8JFP4sDdUat4nbb+LGSewGXjSgKeEIEqplzdwZq2Q6rJVsn/CmUI4iGjEoue
VyFdSR13ikEpMi83XW7xpF9Jp26iDLfBBltOGm8TN8ZhuD4IKs1AXb8hgo7E1ujIwqxvNUVHLEMe
/POGBMmy78g9k+3TMZwUz7vMR/NhR84iitOZd5cRpGBsd8bs+6V7bKGiYe0u1YbK3EUaOD38NYfL
lEUiO2y8w4CNiS4UQypuZu8zHO85SvQ/yXNzr+zt2lR60vfjkd3XqBbYZC3gKTWNmUEYa+JJ3RtC
IWgqFelnh7/nzeqbN151LA2sof/3LtaCDW7d2BnTEl/ycirnbI8KwIAUQ5QlPxtSleBsqb7CyZqp
QJfbeQ9Q+DZCCpMG5mILt9P5p7aCEEEstBPpTlcUMKe0hVAbpXTrE/OA70SfME5bFWLJym13bKOa
TZWotCvlkM2a8vEZ7hA/qC5CCHhBaoXuJSAu/OslPGw1nBambP6kPtRdV43TyeUir97so0jpIFJ6
vJ0m145+UzXSkHjSf5gaPKnG5MsP8BbA1oplU8Q4rzT3O/1BOWN5HG4vgSoI6WG6hZYlAYWj0IAC
h5EPZDuRa71bXBoEJDeVLLvrsHGHsgq6ciuaPIPiQDwEdIz9reWeW6oRqygNWJqGB25t1vnTMH4m
NfW8aBGlNGwvQ5m/FuSjMkqoWmCQYbdh5BsDxUE9Oq+HAiy9T2R9LkZT+t3+zadl0gwl8N1L0k1E
DQu2cTQauCIFAHmOCMmpbGk9jDN1Sb2SgkwvODQHBsFnZp/psUgCb4GOreQ7j1+JNVtJe7i7ZjMj
S2dYbzSwLOQPWp2SKiwdsD+1AI81m5qT6UAHeA7hLR4KDNluUKBFBpYLd6Wa9l4j8QNvr1v9OzLl
l9LZDu54rZDh6hGCrYBcBMwnbD5u4BLXau+yLRBLK7h/q3+Kprxf2dd2AOEwlv5MYVPwUnz+Rzsy
qrz8vPPEnQ7w0ubjWT9usyNPflO99MLOqCI161JtR9ixs2jqYRMcmG9W4qONxTpWiNXLQLgxlaPb
+ydCc67nZkaF5TgBym4c5V4w0V7Bfm20/zfGm1vORNSPqFquxajsJkZ9lCM2sDEw1dNEQ4bUai0d
9JacaDgCdCgYJnGj4SS39E/XjvP2INylxdDfM07ml+1JL8zCKqfPu0/y4NaHuCO0Zj/S8mk7aWY4
EU9AnkeFDLOsnW8x9/QbH8ECNOci2oYekj0UrQusUc4RAAHSeauisL7YAVm8+nZQkvjHPTItAvo9
mTQmcpX8KJsxTaXqQ35fZO0IWaQvsQooYhNJFq4zsZY0mXWC583o5ThEEMUS7c0lL/yosg9TBwXU
SYdnFcELcxfA+P6+ekoXhPRQuUIAXB7ypMbgdbQvH4HPDQotcdMeQgk+r9OP4xnzmG9ur2hNu3wl
ca34J7ELTgeo5JV3bA6EXAj9jMQUgRAigKCmoVD+iSJuPM8DSHcI6mBOdcPUXZX7dCWmvVFobZOg
m3/sgQSpdni6J6ZYvyHT2fFRD3Qx4rp52RNa1OcVd3qEPhE4Dk1Y5dP6bLIP8T03jzm5/xF9Eqov
C2UNy1CXMN3TUAXYz7hQ+LqUMygYVNyiRBFL01JZpQznEyeEOzSiFBJIQwLi2rNQ8CRDCHNT3DGT
R8RH3/LOIrbc50ecYL165XPr9vW9Tf16Bq1u7zHhvhKhPT6Lnbr8txCHfNeTvMpHlngEcaacF2HW
v5nZ/ZM/S6zwESm4lWaIAoi6wdYLUMSuuFIo9Bw8D4FK4eGbDWvZYsZ6d5I+3DRakSsv//T7xxnG
FQArajFLMnZ3wwWSvworY7XoA+WsN7Ysx9nAxOO+i0HlRhjWPP7JqjJPc9kdJk/o5B4YlqOnF3Z/
vBuGjqZ77OFmDjTmhh697WPngGwbeZ5dvdxyfv9JK7vwvasC+5uccwwPabR0X/bB/mstNJG5LkSO
Pg+6ZD7kudaN/huYDWbTwuxwxikOkSwny3+F7e7AAycb9Oy7+FBXEW0Xd8ocQO7khCje0jtKzg0w
1hntM7T+zT85h2J3AHBvpnLjRSLSLtPtpa0AqhskDZr03Qp84TeQuO5K4dPBdLu7NQZYH4BPxepa
hBUCo5Fp4O87NQwpDDY8TzPOotCYewrt/m25c0Vk+m84EOJAdILqXr8SHiR8QXc9I9PAYcPkDcRI
3Uf2uHXeaHr6rIU5oToERo5FExHCg4+Gf8/qD1mAlxXBoYl9qJfxYwociYVxd5nF9Es1P9EbBDad
yK4Oa2uPE5CMtU/Whdxt1QMwOROhi+u0J9RhqGlWScgVgpHupkqi8U2bl5k0+tG6RFJhDxgNtCXy
fWb2sejz7psytSSNElta4JRr8MdmHWYCCS9GdkTh7U7tk9rppo3ICp6WLdODFx6NW2NcuEb/fHNe
Js7TiQG3pL3kGUOQljI2VeLfMxA7OQXyILu8MHP2XtLb0xIOGS0ord2iW9DRqHRQVXwJfqW/Mxnf
hRpvxxTlUpMSZS+BREE4CsiNA6WB0bUomQblj0ZGQJX9yeJsTipggYb8qo1pO6ujZoPDgrf5BcyT
Epr1eTa2lUrma5RcJASwYsLugHLwUDAVw5YqYYbz6EKMgtcMKPupQ8SXkACMpVMuQOkad+xYwHZX
Twl2aF3gH6yxWgAL9ucbJyCKlvlEf/UnRa7fDmWbwxJ89UR2jh9aze3GeJ4GFpOidvbgy77aSXM4
4pgYB3GVFSjSoIICVmNK3qdCPCfFViXDO5HcdIJlS2LuCmnKj74dSwXL9xFKXi1W02oq35Dd5w2Y
SADGJs1ajDyZbuN/zYX5A5EsgaaBD0vyPxark+7Lp9R+m6Kx2T8k3A0zGmgZZbI2n1G/F0XXRrxy
OJIEtARdKXAw0aHB2fVawAM7Yw48bURAj+lGPtJC92QzCggHPLgXB0evcG1eMko+IEJPZ4W7UiI/
k9u73sYKi/McrXW1XZXOhpvh7HjYlPOkPfRHKW0SQbXu/4FdL9nP7JvqR6UbbPrnH3uKEYA+jlwY
TQ9cuxVGAYLSvCjOpbh7DE1tCTfVYj+z09M+JTDxtwcZxBso5edRwuTwPop2d1AYlVFPQSCCVfmI
EtBP4NTGf+SrNqtCXWMhS6d5UBTjijewnKq7FKLI2OKaa3LUvo78l7fhCu9fFTvrtYj3kdHrxjky
/NjDIKH2b88Lcng0OxxXmNelLc3TCRMw2LAAkImpDmAKZdWUwYsD97eqzmVOfoiUtGQsuHv79vUl
aYacVz4kXx3MXCtyXBvIIeJ2rdTAFEvHRXVF1sa3kqJcU9pwz8s3awsR1ycR3/dAFEIIN1quZ1Ow
h6bXnxxL9zwwFsvHalR9+PziYp6H4LMcucqfnWBIxL2vQYSzuc2g+cqVkj0TuK9nI72G2/ogyIDu
lnNL4qUrkmY1e5sf3h/jCZkW1p6eNhC5FgHzWivxRlgYrVwhmGeqCGIqR1l3BXrbcySvU2rydnpd
LSuDLqe+JDmxBWxZE5GfotEbxIIcQ+8d+o73OvQT+aJlVndJ+9hO8gLGuiwNdBmGQzWrT4Lnx/3Z
DcgbuuvUkjuTvmVJv2jg38wCKYCSJefSKIaoBC6FE3jk2XtFyxYqLeYuAwWqABRaa/O/ZgwsHizn
p35ssdIaGdJXqtnBJYi1/5E9ZxyiBLx5i8TzFnljjQpPAkBaMlUpAnfoL/+Wkw9Hz3p0obNK2AHg
EBQsu2dmJ/w7efcESdqbWT6YnQ5bFpkkTKiVpKe1aNZQRMLmkaFhnfGQW/VztOufV8yZWcQ1KoqW
+KlzaiPcMpZA60yUciOQ3ghEZ9bNF+8O4H7RnjVf7UTRlpSFj1vW225mEoCou51xMlK9PnfE+yl3
TOQ0HTn8LoYQFGNqPOSj93GEC0YC9njsf7do5pG4DZk0bBOwolbPrBQrtWl8hueqSBbpOB/D0K4H
O3yCZMY9Nfh7LGmM9Ga/gtLAObQgDTcotLgjKbgWOcH0bpiai7u0ayt9KwazmEUpDDrR3IDU/qmS
2rwqg16Zh+3+ZOyKyoLuz+AM8j2Hi+GWhllmz+pQIkSmIZjzCZBigAXabbEX7Tgmry+4u2aAIqhd
s3OxBMR76sWF96t8qUXxmMBmMDMztCpFLfDzm1NQCXJE7qyov+uHcUNA3tSpJ5oKMD0A4A/GfauD
mFsKDz0sAm01BN6NPliU7wnHd/guTIiI76tC3xDtHinzlRuo5pDQ8bvl8w23FXDJSyCq+DQzXGhr
toVLCXZtblAAlYNDHrxGqTm8S8Yoy9TlqFjeRG01oUbHfc+FOAg5lEfysMiClXMDJALEDyl1KEVc
duqiEUZTzcA/caC/8/07tUGoAduqLecvuRgf3zj4Nu1B8N6owTCpdY7hqnwxBDpSnpalC5qd8TEE
LxKuvaUVNkW2sHbHLt2vLn0jHnFshPT6BmoIEgjV1rztaf5Fmtnvodhz30Fv0Wp7i4BwTkUVckCI
Z+fIeMjwMFqquY3YJfkVEWa5bOga535YFSsC38ffEXNet9iHXXp3AL1F66o7a6CGNFr+sK4qKBOu
lNS6PIFyB7Dl+R1cS/fPwJbhzhgBMea5IRaAOkyOQPyj4E6hiwK8AzJMulf8irOIMJ5I1YK2fJd8
oXdrGvad2xLTM8bPYbruMM1hfdrtMRl8ptDGGPmh5Czg5OoeUYpYFl9lBRsBNRNyy0/Qev1y/5Ma
P9sOkYM6EWuFlHdD1gCTowtWguI65irYrD/0rMC2mlSSwfzc9M9ar08boxpTu6mt6o8Lf9qe7lKT
dt6YtVXgVUo7/IvKVU7bL7UgN2BjS2VqQ7gWLCde68t8trxHNQR1MXwvkJ3XwCCVBYafwThon5HR
5WcKZKI7AN/lUJeSBi/PaKjXe125NdDDh+2/AIKd28JIBsQxvABZbmb6bWcFeFApJBvnuCJtnCJc
/Nxi99xbwQwx20Thzt7JQrxv6u5/y8vjlXMz345oQNleBn2Jijr/HHtoVUELHYVScDa+oIE9StWx
jy7hjSKvv59zLed/DUAdAew2N17YySk6ts/u/VqCQjCUtfAujv7YiVt7ObLWqYQyg6i5p/LO6nkq
Sj7cLcCfSOVlaZ+mVB1vXhVNBTAci5OtsMmsNcvprPHaSI2R8+3sW3GokkryTAfuZD7z8J+oX5Ub
1ynmMpPzBCIpTvQ0yUd1inGA/wPby3ZrpeK2YD7TjmdpMLCzWbHTbqy7vZn4wrgaxI8KTSlbagr9
hdAfzBdWzikO0V6kKvNx4Lta0MXRh7zE+Slq3kSSoLlTObsHWb0EcLyQdsZ7Gz9ZDsEenRHQfVuQ
IAJBPAnScKOJvBTCP/Vks4NpXdteDX4kp6UeH0QZjCNf/MMhuE28S2SmpycBQxG3zvlzTfk6f6fs
vN802xpSQmm2Z7gnZiBXjBOMbsdkouC8X90P0rbhz9bxdmarlgh4PhfNjW0q8+xYwrPovBrOw9s6
OOv8ERrlnpYtz+jC766NyPbETBS9vVy16sIjr4vtIobEa87O5k2poCEOJJ/LsyM9+5lcXuJkigOD
yHwq1UaT5uhws/rUVNcJiORExeSHR0aM7555ycHSNpuIxjdf1FeK9XmMFodTute5RzJiN7MECj98
cnH11f+ud4s399j25Tk28PijcBukVh+Dn6+M4Huz0ScBn1O6OZk6d5YK4DDru0ghP8mQa4SOL15y
HFV8HldAVmcC/xDwvI1QBsJgiS/HAgDvSvyO85KjF7piCpZ5x9he3+7D0SUmLzzvV2DHS3mW/of9
sjYqEjlLFiQcH6mZq0IXZTl1Mq/OxQcuSS232n2tIeuFjZmX6lralSbOBhqAkiec4oI/MvoOMCy/
JA1tnLo2b7YB57thzWLrPjamirC92BQ2bz3HlDSmKGAGcXN250LXisr6hbktqdy3gRPK07nV3D9K
c0XEoxZfjwTLMphuPe/wLFDaUdfCujap1WoaxOjQ7VUIWhFtKkw3BFOcQl72J9/rAAcDiLZD7hyJ
HNHkBpmi1DDtcTtV7uQMoEOQZHZBZxNFczRZ0j8TzZBEEXs6OsM6+nBe/lDzW7p0eWP1KCQ3lgaX
vhCFo03/AsuVTodfhg+6ZGNa05Dj9bCoUc1RcKvtlUsLphR1+X7K4383DvLhlr2vwjFUg7OUBMNw
hJW62ASxek/A788fzsjZ6MZtStWX9pZg5sNYUnWCcbwX9/2ilvFzSxNER/2Oj4gFXcmoo9a9arqo
zyocDYAt+ng/YwN0c1nBa0ppJMQKZspnnKmUslZxpxHePuhSufXn951x+4XmiIGXkIRgSXhrS1tY
7D+EjLYZDpPwfD6/yv4Ke6N16m0fomX25pESz4e+dO2OHVaL8sCIN7pawPzapV+67vNk2uZGGOfA
y267w2TI/ndZAkWKsFWAFax7gCyryYbTnC6TuRABAK8WoW7bPCWBqjz5mrezeKUF4ffNF/bu3adU
bJEfERtw4PXHu7X6ZvRvIovO+OtzIVATivIeX27nlhCf5Mdlc4yrTeAWBTnav+cz9YOUBvgR8qGy
9U+Cw0j/CTdjeiMei5lohWAWU4wQ9zFa3RUXldtP92jSCNS7tthQOZz42R/WWqnZHn9buIf4DZLg
+yiX+K0DXBqS00ds33BHiL38h+fcOkeO2gdbe6lROQjNS5Woq0nDq2dUuAyVfAORsG4GQoIRAop/
SppAs1sfxa7aSBSCjGdxr+AVAyquYx2/cLxgFYccX4RYbHT4PPWSQtxCS2MJ5ge1bliF1hKnPJdB
vdpgu9EcXN99YFP1y2jRPYVpM9slsS1oYFrGLjDC8iueZyOmyN0en1QQu6iXKZLJYXUi5/vQAz8r
WN7iKyt2x48gwthylh+0spaQlmLurVjBVuCzFyCadIQotJ9Dl+AMx5iyMLBsur7XOtr1ppdvtYR3
PtmR/o1kGKiVYSrrS0QPTafVihd6183/Ij/ELF9FdTWk5R6cPgC0f9/X1vDMLo66+w7O3Ofm5GLB
M09bjwrkCwRuPFaIuctWsY2oexrj+ThxCrw43mEkFiJ2Y9oLzmwH3ljfobpjcUeTmuQddbJl8+2M
hJ0FY6TwsiT6h5c5aWeaKonfHTV9NxAAE45LfSsnAiUrdL6YZLR09U/Z9V3dASWwB2aHCqGwDWzq
Eu1eetlycU5U3cmqGEfugi9pA03vAvcfMHEi8FKeGTyU3sAesipawlQ4a4gzuOAK1WyCGFIF5wQq
oLPmdTa1SziOiZCZ/RRg09v+1TxeiXH+feA3ogSWWTcynaYjnuF3EIdlO4BvCStre5DQd3y117Qn
fML6Fx455WSWwHrNeBlN7NCNx5ggLk/qo+jbbjq4AXLwaZaw8OswLzxgf0d0YSX3I620tCuuCGLE
uX+Mr5BH3mpqhNfDywlALLrk865TXb4NeX/9HyThEPAUMXtVgbzmPowmergMRhMcJEVK4xrOHOBq
Ccnk03Ot1hC1yOFrphhcD92YP4YNe4OWhsD/rY4bvTHq/vm+x6F/QuEw3Bw0FMffFNW00fujfpS7
vz1HNkM1VOkPwMV7vY7FZfykgTb8gk3R0zToNq+S0TbgattcDONAr7yrvO643Y5X+8lB/P8QZR2M
Dr4PR0jc1jzLe8lcJYDmaw7mhANQwKyZx0UYTsH4RxeMcjUKR4SCXdsXEJak64T0/TH8mI61GBue
QXX6eg5dT9j7oG0aYm9GlE0xB/GLU3d0cwZbe6rBSjqu5THJ3SA5ot/hvWb9RxqqQK/2UdBc54GX
2YYamCzmSrLFTe6g7nk/dwqcrV3/rHfQnYjV0Dtfek5r2IiYCqaP1Y4omyGY5f1nBXfnJ1N//OiD
lRTj9mPOD+UzSmPffP3xh3EcYAExNgTXBiAY8FQdzxXrlNZt24JDYYIx79By2bNvcHQq8Vw9b334
QWGlaXuTYBY0XJJPIYUkqE4vNW+H9CDkavAOhlmXKkYpy7Iw/Sv9JaDUerepRg3u/2FWIQq5o+ck
l7zN8tPxW1Df/UQ/OLC1TMpLxfgJjYPfnEteELNFufKghynB4ydeqJfwK/uQEVBhVh9gDfEQLVXl
CoXcjON+eFWOdJCXzbZEhPnfUgCVc3funwjRJGxZSKqQZh14JbKU9DR3WQc7uRo7oXiqi1v49e6z
KR+RtGJSnY5ZNBMTaibBx347WTo1b8RkGawLgA0FzQ/xRlNu5QZu7Az4TU83u2vXKS4L5MISaSoA
GGdKWV5ooPrgqKy2/wMJyWk3oyPfmfeuIJpRNX4onW3j3bm4A5l1/lxnYIsFsG7FF4tgCQ2DTiZu
OAxwAVC77ldm2tLpJe8R1iTOMA1evOUQvKdGWWPvP/b3oT3b7L4XQIrPxxFYxhtypZYs7sYETEd6
Q2Zm6ui6VH7CtJfHKKanDibHVyOuVHLpay49sHkJ3x7azrYLmIwL61EVos5S8oS2R+so1GyV85wg
mxGxCUAereF3GtP4OhNSZhUV3B+FWWDG9Y6cYe243X0Q1vJXph1FeUbCnJ1KQbpYiFpy/4UR2lBh
seSXdO/6hSm/eNgWjXk1LFl7afv0/cXgD57n0g4AGq4aHFcV/QvsqylzO5DOk/yZ3lmFeU5NzMDT
0msBQUEIoXPMAGVG3KBsE5xtjhgTqGlUE3tC7LAh7hBx6xsphUzwASVG97mQpVLF13yTfrqTkQLg
khm72g/S6f1odoayHnB+EaKnLDz0z3GE7kbjWniGhZfFPHz/vLUUwVAXoKSEhEzSQAX2l0Rvk7la
MTh1neIzJD/qMOS2vfFRGEf0pxpCMo2BRJu/x4/X8hdg8KhaoCTHwCIXQzFw+6lmHpTmiRUuENd/
8zx3axrWKq/cqE8ExWdnRxhElfIxjaRugytSghijsPKv3OIp7rvEnOWX2kYbg6xn3ogdKYmn09FD
ZPYMHfI1nuAOFNWc5a6pkTO9d3B3qdgmfurMKAHTuray1pIPp6DAPEtTFMHSE7ujgPNVd2c+9egt
Uw5rozixkW7pOToZc6PMuM4yCRn+e22Rv+K9OQDXd1C3X5Lu1T5QB58InSPykfgfB1ZpUfHjXbcD
+TlkiqmlX8wXRnOZB5dT1PReu3tt+w2eOq6ijoVI31rDLk1SLr9mexETHE/4zsw/FlZDrP3yvTgA
cdpTv6S3Blq1tBzuDyZd8cFnFo+cvGupFOUuOrrz+1qbieUneIlWYpT7AVbyPFwl0OoZLajUevrI
ZKoMX3N6kuEjfkBHhdel0Vr03372yuPLI8xhEnwupNvXwXyPPoTlHY77pWmopkZfdkNlM5TtAwRS
KBDbW8xwwpKBQhPN/JpC0GG0KLjBp0JgZs+Wc0qUXaRUdhb50BNF7sm/zkJYUe0ZOFqYn4fadpYh
z8rV1FKdlV/1UP8cz7+u97O+zl8IM8ZCLXZKAYlJ4eJEbc5RZBtxAK6pb9LOk9+4U5qnA9Fi5rkd
klHRDQLIAE2JMlO+i6BaGlA/gJLLKZ40MJfIpddHoMOQWV/8Z3daxmDG+quftfxjRdlaXaOTEZUZ
/2FZugzADdrq7jNUDX1j5yQ47J/W5lEZSwaX2ChzedSJNKrJkwl7vymg4uDflbFK5YT2OObZ4BRc
oa0XbgdSdka1HRIALpH1mFqU/bAwJPonshFMHSz74tyP9IzWkE+7bqhcs5OP8iJtJx9Lls+B7SeJ
/VqrlBhvmibRri2kiegnLW3x4k2y/o7iUjOga+A8mjPp1EnhjEQ9IEEXr4afdizVI+cLCXBQt2IT
fMs6tGmKiAwSsHOD3xObmbtRMgOwog+SDW8g0yy95kLxnZPX/jxaYe2Ae39aP7f6kXAgQ6H9lApv
9rY+W6f0TCDXk7OoKnOuhQ9rLPtegb6Ej3YMAONh3Tq9qrBKBWp5D0yCOKeYtWBHKushkfmcdLpw
Iotf5BWZtthFab/kIrF6YDTc6EgIGRhHKg3vc5ZPsC9rhW9ysFnzgEMQ/4vqWiSvFuJIFRlG8u5x
QS8Na5mtI8ZyHZ8wJf1akRJ8XrYV8zUVKqSIwyzFx5czVWjnvDu/6wrknVLbw2CJr8vejh7F4Hm7
7f+VkV8BeBERVufbP0wTzaUw0wpiyHmnK5pCNkUi49JKSQDcdg8bKNe0KHt4OwUPY28kj4oHkGjW
+SXWKflwOZB1KkST2eMsWJLLqlN6TfT74xNt8EAlU+HD82eLuDyumZvQTKZBDXKfB3xO3zuDq603
+hs7NCJ6XbKB6GaWWnM4ys2tlfMQpSHh1eHcOwkv+Rrr/uTnB7c79xkfAh9rnCXtGnxaK2S96dbC
fYIIPbdW0MIW5LW4YY863kaDdQvdyPNbzomLXeUGl9M8eoEYAxdrjAkuHKHk77fXGECiWuOMJ+LV
ZRyfBd77Dtb0i7oi3e+GC6y86xr2CyIRSk5DUchc8iVMWNCv6xSKs/Fe3IbFynwoLhpo52qWanz0
8ElARoNnRNpveQdY/CCS0BxhVM8FmDl1OO141vLCFkjJI5o83spJZ8Xh/9vvYtqBk34q31HyGfzu
ftML9If9PIakYuLT2GTaTs1PHjJaN/dcoP+I5/9W5WT2WgVKiKi0lfamq/1Tf2Qzhj8gTFvFOiWG
qm71+j0IeG0ogSJz83ZZ4KMmc2WCPiC8Alc6QFclBWlhx0Ll0IhgLdGs2oguaU4DZi+VGnwVnQ0U
mGQeKSGTR6B7aZUBzj/9Oce15Izg07Zbff2swImyrhDKOdQfxo58p7E1JnIdHseqDsmSz03yCYoK
Rh6k2SeECrU3hiqxagMIzum9dBy5vQ0nFmRJ54heRkHEQlPeJN26W6zA4li0q7U+zG3QRYInoIYr
TsjaM2X+zRwt69IKNfzYdEJvVLif3zp/rMucoH9K1MfeRGL4LN/TKOaeOetSVABW66+sg2EhPCrn
p2bnMOe72rqCnrmwKlXce3gA5pgCaIrMMZE3XIRxVUYhiz6TMvHNKAkvP1T7pdZ4zg7DbY2de20C
yetF1UrgC4VeJ3+iOV2x5TxnEcgJ1ebRbarC3+n1hzu5lhxfPj6lEhfRcaDi97s/pPvPIzyIrqLL
qMcwKrWTPz0KmRT0ofdffSWIKNZzlqd7vkqU/rus+WyZnagIkqfW4Nvu5Zf7xsr520QiqharqYxw
3W+/NCmuQIkHoaBiAizzpPX1v5JGC/pXCdPLUmi/UTn9tT/xtyG4f2R8GhiJpXSFPl16zOt6Iz+s
dUlI43ZrmACO857rcUvbosg28kIJMAdH/b63rhrxt00opneUu876xqAnPO6e0p84UpV1NQxdXwfz
uZdLB4QRyxx+Sx4cJR+iGwCVE5QpZGHeo0ZNgHoqYKDqT74yUmrRfQOd/yXNj9fF4RaBZemSUeJf
L3Bnz2Xq7em1Vfyn4cuMYQGrMznJOxCCiijbiHJ6AEstrTBcEhYGY8NNJww3SH52KlmTPhcfA8sp
XkuknJBgLK7rPLOkdq3SjJCGyyeJ8oVpHME/n4aw+cv0xGNhhqIY+A+IPm/1UrTFsWwcs2IAwZ9Z
7KG3KjgeYc8OrhoCNyICsOZzqKSmIp1kSqmmNfAbDAO40yzV97OWtoSMNdBIRHL/tVWaOq5pMFyF
UqNK/16V4jC2yO7xoyJH+aUTxwlMM8X3+5aU8ss8rdTfzUMf56WEQ62VE6oDlGsz1ajJFwl5AhCb
itLpAGdVlwmMMnB7X5VMXEEO+lvv1LIIxEyVTcUCig3vhfh/arfIIGlvF8CXBg2i2/L0JeeH+Q08
pH7MWKcYFuGB4CZcwZDtkxYxvMVxW75vrwxiP+KLJYqoVteHQOxUywODT5H7T/7wXTTrecBnNezR
xzKkGqIc9qXyh/cKzQku2e/FQi1PKE5S7PlVZbIOuuqKSUjD1fm2OchPCD7O/eZPbhomEfGuYjzD
qVqrB6Mu/huL/WpC4KQ5sV4135J1kpNEaNhfHYnOagxBNSPsxs0XHLtJgsziciT+p++PzLHUIWq/
j6PvsIjsNqpshb9y9XE6Wab/yAv5vWRCaHAka585mFFwAiLOCb0zxD+PFJU3D3Fqk+cceX1/ma2y
tuUyL/UDFN0LNKlDF4SyE+83dvWqEmTu/Fq4xJom1SXVfkoGgh5i4LDKzqpcIVTZ4XATJJG0+3v2
31n5BkJifaeecJ3f9utiSb6wlDiMXFN52fX6LgkJYI1rUIRpFHd8IbVxtpn/Y2CVXHxWbG4ijY5Z
9CiFCLFNfL9xSPZ0+YFpUpq4VPRmQGs8E7em503ey1ULzPYoVi+vsWehX9bFSafsz7oB58yGLvB2
HYlyZSqr3nmvd+pRJQ5BNe8/fiKyWkxctb+1iP+L9R+AtUtbTgqLmGClpDBYYVW8Fgx5Vvm73cUY
EGd8TGCZi/IHlaryQislTWv/gmBi9xyAQHT+acX3j5ueR08qnTfl0r5vw1xlj+OTlDNv6sXmo2vO
mCYJ3rPvANXRC03wklAX8N9jLkr4kkmySit3gSxtfjFiTnxxlA191FXmYZF1Xh2weLeB0CL2aa49
0RZGsN0sWP2oD02Fb5LAM2QNPV8CNHWLTUHV8lgMPXkUppz5FOUL7lCjbTgRoIeu7CLbZQY9jn6b
NBaBzCgkewVckGqycM9zzZwii1ERTcK8GeORHJzwqOskPZNGA9kPNKRXpWlRDDhRn3NQ7gfCKKpk
bB5VPK2c0G7rS8zIE27TjKORsgF8VccyilWSUCmZIzcDRSF+bSRVDE0+luNjcEFQzTgjllWyoRp6
yhNOjoSZResSHoQNoeHrg7dXBeslW4RZvf2GJ495p+5tRFTTZMkx3215L2lDHkDL/dF/ZXP9+Hie
A984PkjQOUHNq+UN1rGlxKESldYw69fpWfiFAte0CU949suQSRJte1vIACI/TTvmNinIre02jGB9
FaiadsEyAWKo8YRmk2ufCgT/B4mgjFbyfbFNb6CmXf91knb9gRRRvULVGhhjPejblHD5shcDug/M
fircsz9FoWpjoc6xw4oR0WhJnrowz4pHtMFY3PJEC2bb7rxBgC6WobSY+qCPJDuU4BgYptQCzt44
HtkasngQLrkV++M8Pi8FLsEbMo3W7MA3yt7aC+bhXfeQRGoDir9I2h/FfCnJFjraJkojmWxQ6ntb
Ri1WcXavU0O8m3WstzUDvt5rb/5ziRsfmn2HyRCJtTHxK+eB8GdKeFWJ3XnBItMHtQefTXcL5FTA
QVseL1KbJEPeYF1TXdh4Jj37RMFnq56SuSEidtQ33ZJhZdOafMc2a+PSf22BOjqr75PlawfwbGMO
zQodFnJ5bN+5fLmIMK5zTNLh4f8f6poF46+X2pxlI1Btlt8LwpBerJmVBZ3qcN47M58otqSe+M8K
xw87E5MeTJ+VFiwrAOVAEZ0WQXckGYNcEPmS4zRTE8EnepFohkpk9fuiiJGWRcmTVqnCcYhMQGwI
+ehXmaX+3oNcG1Z6/eRmaWlTvFHQNKCrtQ/gaDMRKvpJGcK2r/28hZNHqn7vbr6J7aMD2LkyJcDv
BPR2dHsCTIv/8d1f41hLhqIwjkluYwhkomwFf1UxcruFjdQ/yYghn8UgzY6knYQJyHoJVBaLkmBh
V3ziXBLYi7JvoJQ256qNnokmqafqVu7WP2XXIkdiytS4kc1O5d3o7o97PNwr1teIWIlN2T2m3Pum
UK+OA1ue21+aEmbmkzI+K+HlwjY0GgVEWSOuYGgwQtnF2BSYnTnAtNU5w59gJByhyeYsLgQPEZEB
sh0MRG5O1Qvlx8W6pjZZMKNt2zaS51pDUFZd6GOH8c5Mj1eEv0Ingh2aDPpmJW1IPz/3x3qDd5Uu
Lq6dw7+vtAP61nOD86T5Fs+oh4nsYuDN04UQ20sxNORRCXGEXS+5Dyu4NSpW8pgv+mQML/MMMo+K
zhVR2cI0pYzJ98/+pApy5CXoeVMXn87Bskr1gd6T4tEb71njK7lwraHznmDsrqDBRPqb2wBTzkIL
na51BOYtCcJaaDQX4/kqAmVIQgBvkeJKyIJIKBVEu9tZJtfQ5fI0wVSo7KyzVoPQtwe1tLXf7hYz
m2rPGcewIW4Zh3JqH+iUqeD3K3KE8vEIV9e1NBgL44lwzAC0Iisk6PZG1rFnxBoNUKuPBnSjdOX7
2J+DsPP1ZFwyXLINAhDphpC1lq6gg6NzAO7S1oN1eZFoK8Qnvy5YftVsIiLlixkZWjOUR0NTH5Mk
AfuQJcKdQCX+g4a4I9+11VVm+C54Rn1u1iko3aoNCDdQuEQzHmPJUyFDq0GQAG6YE5L9+lx9TH70
cOKjxJrJ0g948N3EF/12gCbEyJJn6d1kADg72zqyawqJ69VSi203gkJZqwGYBMwRMgWGCxjlEiXV
u8nYlrj/xtIV19zNTBhSuyv+d8Z9n4XPpU7KL1arxh/jlbrgjCUgk/79qGHwzX81XNi+8l8YUx31
S39ZXjqWLAnBltgJq0p2/KXbcQaYY2+oBja+uyfySwYiLsZ4ibQnzfn84B+uC+iPPJHf4ykOqlr5
H1SguIq2wTvW9vFzXC/2K/RU65Fen1tETUywsmfpQAwiHMwCTZeTJCNeBSVqypNNjzXBQXCDBHcG
2YKltRhfLri0POFNZIAaVbeasoyT2z9WQcnms0qpXwafy6bwRH+/4S7TLBEOuelMtOotnAotic0H
5IikKOGbP/3yAnUzEZwemoHfptrnEmGtIMWHH7i24hPpm3g/5WuyQcVNzM8vAhK0Urq+5HG1S+/L
x3jdr45FZUR3iQ/ajktaBJBwpIdCGaaMSuSqiV2RVlKv9enUYbGuWKjAHIroQ2xHCQPaODoJp+ja
Nc92g1SWb4BKj5hW1jpzqtmDaNHpEAh40EZlCAPZrBfsx/E2s9aSScO4cEH5VEnpov0qsy9EM9tk
OXz6L9pWyvo3cbmDpIXefJdVgIZyOkdo2pD/3fasPKicF/U0uZJrd9JMQDAYyUlX00bEt81aCSBc
JwjqFVc2nsT15V0eCCJATGFFAZrC/eIZ1AwwYmFpNPokVMdM1kvXJQV0XoTkh+dBfsJme5VlAnxG
cVKTHOHMsdNKLSsFEODo+VDHaazk/XbYXjIPefaj3E9LTORGAy2sWrxv2BaJp8SQ2D+usc44ZlY7
4mlYLW3CGvU8JzG9i6erTVvy78hsbmm3Nc/mMpOle7EtRNLoN+BQB6kWzAWQMklq2FUXNkichgQ8
XNpSmlGwEW61Hcka+bL6jW/W1K5Lz84bwoQzxHCy89u5cJ8L9GR/pUY4AwNQvK1L96+ECIXvZ6Gw
csRnl2csQQtx+WbVfCJb+Opjl1fF4EyWQW9QfDLSuSnuCw3bs7z5HT0ISlISdM5DfN7YDFPKhMR+
TXjkNZaGLdCZTGCkMd2P/WlJyHcGDEKUVDF1Br86so03E5ZypuskOSby97Gp3fz37wkarP4rcEyK
+AwkE7sG/NlxAxiyBLXu+E0uctml8f0BHKdzrPtvRvw1wCVZkBnRhgkoXdHVzowPRtFhTTI7DBbG
6RDFA3OJGfdU/7z6gPsKUF+0wwBGCfpy9B0il/pcoaxqGNRttqvBS2u99IAz/2mNUSdb+zj1+PJB
ed/nybAFp/iyo7BDmvg99iYgFJzCgjWpVqHr8jJ8KzqZZiyMroIByIjiqnDXPqz+iQxymvSeFVfq
lh16LBgwaR8Oin4vkD6FlPauj+/23A2SwQQ1eMQFuYfgL7ba4yhsFNIriCDOZ/XnqhQCQYdDvat8
rORhkyDr8mwlxPIjWBzGq1d+MbwQWSBFvRWFcly2g+uI5VXTGlTYBgvf1x9S7Sla7iWrur1Jn/JS
3nALQaXsiUFYUvM3aukw3rH7CSMbv++ncKTrbLXUw6VW8FjqCin9ckwhTwCtNNOGlVk9Xk6rKOrT
BsfeFGzBDvlDD2oc3zfRA/0Gttk4EtLrMXK6LiroV5cMCv4a/setkgAhLYAEK9WydLitZV0aXKUD
gMdGkuE1A5tgcrmZhfjGYa3KnVEkLZGVcdzD8nVbCi8GF6vQP/s1eiix3Jjj1l4FmKh7x8vYFCXS
2gCQBPOOhdULVSx3gmmGoHmJWtH8gXTkcH7LCFMubE24eyqZ/XLzAJGY/xeURAd5p6dZfZmaeFQR
K8GmbHs+rFMvB0VZ5YbuocqdgdfFq/F2Miwv8hpYKWLEQb02SFb/FaTWiJF64MDsdjueIhOWVSs5
9CMA/GoY5EfaVTb1yy+9gQ0TyJiI66q2k3pc3N2FVpmmuL3lbiuJJG5S044CyvtcdUk2c8OoGwzd
eeiutkUJZRZlwFvGUkMCBPdPWkePkx0Ely7gBWvwxgpMvthM2THrKiaiXdikd+S8P/oxs1PitTOH
ZQYGtKkKcI8NQp5ItqDgG40p9omv8VQKmMr/nrPHZMMb0iDkVF8uOsU1bjBZnFUIUkwlVpSfrSdE
DsOvL2LtMPj4QsxAWaanpeZKeW39+g16Lqx3I0Ge2sx2/CEzA6rIkbIf8/7Y3PNuLAQdRU7R7Yph
adT1ttooTYOe2bikahDhT6EmXJl9GP2RFNbfFUAN6Dn/mJrIOH1ztsdSkwAE/39h2Tt9PeHUsvn7
/KApmDm85DQrAgQaxkssJH1zIGZbl/KZfBtYbOisSikSflwvBElyD/gSrPOzv2DJ0c+MWFfjXYtQ
G9oBeADpHR9P7kj3SBOt94XFVTLgi8oS2wBnlaPO0oxzXrUVyqwfgOsxq3J0BtXvDuzQbWGZ61Fb
/BiRzQwJ79eUYGO7/D+dsPQwiTNVy09LMcVdlCm5/ljliIjX95TbN2y9IO+gBoi7mns3JoOeAI3S
B3avK5agJP2gltradTsSf5801k6JHcpBDtzFTaV7jGEci0TSKx0mjMCWwcnVmd9xEuuzkV5Br3wj
lGaMr/RW6kkD/LCV+1F5MZDqkC3BAcViRqIvn5oAeVQt96wTTwtTBpDCVsru6ZJ+pSKquOayykap
7cD7b8NDrcTTI3Dm6G9ZnvaY1b7psCSRmyvcToNTw+DwwTj1EZ/GTw+BleuIL6L/5JH/EGClt7j0
NgBgtWDa+bahQf+NoAXndDgvzxvvDhsL+JANh4dy8vlS3J1dK0bo7b92hFKfQFQBB3D7gX46UAeZ
7XJmAFXhdJ3bXCS2/OgnV99vyyjWLulKr4YOigC3KWjNjJtAh/y9YRrKEKjSeo/64yeK24zkvdzW
N5y+v91js4ZK+/FKjh+Fp0D60CVqvsbqVd11KpK6ISugyJPDKT7RrY3pcMbAGrWt3q3LqovJjDeM
dlhnNR9aaQU1s95qfht6T3jg1tpL+G0r0aOKLyotAD2qONzwmKKRInZFwdfVbWCeIlv+8b4Wpcs9
gVN6LxnXmnOLwEiZTkTmrW+Np/VcupTUj1abGoBuyIoIL2nM+Rmv2UoWzk6OnqUoHLZ9K24ll0qI
Ms4vjbP0YwIJa7dxhHtC95iVJUpm7nMlr+H/E5nA98WIXC0FIk5uyt4VV6aUQqgpAiScIVHOs0Cf
9vHXZF5W40IadcmlySbNxxpAoCl/rAqNaZfqcyLX3DLdUHb/yTseFqDaU1VdpEI+jWSDLiuyWQHp
LKLjjWZgGPMaqKsMRjzQF43vsjMFd4XH87Dpn5XZzJ2HxVp0QYjCG/OPxQJOztmmXyCvWfWzYfbj
X7Wey05RN/A4ctLw2WvZPuokG/Oiwjmm22xfA3HO447Bx0GR1A6CgSwdw4tRPAs2BDTx56Bfdccg
VOLK9SNvP7h+g8n1oYJbmPk3dMTgvNCUHt8yAqa50f55KRmR8LtxFbLjiow89Mbm5viz2zXOvkan
ZaJvnvRq5s5njUg9PM4cjdpDPTGP32o37ZRpMvLvbRWXBhwjWErAwtOcxqY+JpftdxUCfO1D1N1H
tAcsNqjr9R7COec65V+tTgUzqt8wbMSltzH8L4ylRpjVpTRVev7jKmbGPeTADaUEpM0Gsc00Kvpc
nW6XtG0FffoItWwzEmjmhIkZh3F5SSgCB+jfM6xC7x4X/sd1tp+4CjUYj6LYgaE9jsk/sXp4U82l
cZzGNOnYiYQp4gANdVd7jUScDya0XJDpS9q8E0QMq9n1V6qq90NwuhahS8j4opEASdCQc79ZNubI
7VlhGMj99IWz7zfdsmKHEGwmQIRIW4RCrhGPvyps9zPU3HOA+cRXv9N1Ko7404H/qi61pktbajrQ
WdhD0YsqQ8i9lqav4TuTCKviHtVTb9N+kNV32NK6C3avxdggvjyRzU2fnB5DByqlQq5tQLIK8Hqw
yB9OS5eNCQP1GpPdo+oTMT9ISdrRoUz1zPZWGuh/4b7x56CLAnbm9uze3WWYP3r0PbYPBrZYOCFb
HJRAmdnpjpQQKjDshIk/T/VXcKZbgVLCDsDZI0HsShQC3DzDZl/b99QafHBY7aovESv6h+MAWc61
JgmbvYIrfiJyricuzJBy5a1Vc1zkoaEUqtOBaqvLqHsiU4u3jlayeuc1GN8g1RYQDw5XCoCSKxdw
HbBDrk1wYUCPnyU/S59WWxyubqeWQhNI5+aigFsOedRxzTfTa/ejJQ7WcXcgAld0lBBS4bUK89Nq
AARnrnWU3Ifkinir1k9a8m3HpbIRrNEG5rmCXLhOCwn4VqFu1ll6DKdgcsiRBNZx5KT8SLdJEN7J
KS7+GzJl+tpOWy6mVyh/Yqgx6Xsgyz5T8WOKieHRd4BG2XqkvumHL4PillljrqZh4XDa/IkS8Xz2
9MuQi2R85PHAurwN2mAi2ONHnyUcdL2WM/A++Nef3ZBUrs8Qj+XWKipFFAQqAS5juo709nyDh8Kx
FW1KjyifxuAouCkLdSznBioWERp7f1YjXqJ5+Ky1G5Dvcj2wzEfXct9Cz571g7dXDchWSWxj0luz
5DqMCGCREBFGZyz+wpU+aep1LgGDDc8ISpIz7p/A6ll4l4b3CoTJoO29Iw1Um9HUmnDjsmIu5qu3
vqWbbWKcFaBA4P+oIXADNEwNPSJjDcWgGzu5KZGQ14r5i9rIpq6vu/5oPHYV0JIvy2hBtS23Aku2
LOpUpttidk+pNT07z5QgZK6B1Hez2z/586N/UgvUiGv3Bb/KUmpLYsG3el3z1tstxZ7AaISFa3He
IuzEOEHsLGmTBcBP7g7NVbSGiZJCo/WHsZ24hOfbhc/w7D4NQF587jU+AjRKNaE6DhG4+jojsfe0
IPGo6eI3wInr/5EwRadVci+6RHziWBmFTgcLvDXal5C0F9BBKdnzjMVhlouITej/zi+kwW8OEWCL
gMy5BKusWthlRNv2QPy5Bl3hwBfZJhegb8c2QXLT+k4rsuOuqoeRSYBU4cKWHbwh9U3RGH7aUTW/
FFa/3KuGwmgNZqLIa+HZRfBYzuIECaXpk+rsbt5JhfVZIGwCev2ERxm/uWYwV1LFeTmBjPp0Xrv9
poIxtrn76KKprfEnQPXEMN7yj2XF6+WgQatxF8qZ20/sErAMdKh6yj2aChR9k3JJbvVvVxToPr/q
FiJ1GWXDUKOA435j/7N1vF3pJtRSMFt20xpbR1o2XS0qbLh9IM8lBPHz17OEJi3BFSq6H2agc50x
VVDY65gMShm4EHNjBYuEekKjVwSfO0d6DoW1jhpykVyTodE95WtYaaosI7I2GQgZgEGMnE+QiG5C
zCaEZxAptu5K79G1u5QwfIvM+Nb3G1Ug3eK6nrqy9nPtN2HqMdO55G2djNwT35wL0u8DZFxXITCO
bPLorm9wlwkCiEGwkiOQZugnV871UtV/ZnyYR/6aEoSmQrRp14MSUTE/lcAejppm7KLdbwJzz6hu
l9wk3I1KulhUnFkSJn2RoPKjEbQIATFGmIFI1mG3S01AxkOV5qexfG+IqGPEBtR7ftTzEuaMF5B2
HwF+zgWewjoMPejjZEXNrunwdPT/ltaXPPEQU8DL6NW1DZA3OcL6mU/bJ60igtpG2mix3JpqzIW3
kuj1aOz+lnayKdT4dztHsU1yH6X2G3PTZqazpKL45Bx52Jy7XsDOayu6jjUSP43O04xR7XDJ8N6t
iP64a8K8UjVJrbLEmVLA0ciR5IqEDXpXkF9bd0DW3rWpnH56Zj5czzDG0/9z74HxdlqqrdEYzILE
HsvL0cgXruu/DdPCzhn5WHEFPMFjG8N0AXz+ag8lnyP8uVPIRgtCcskI2VcN0gzFJ7tkU2K39BRx
3597690UFMqiTy1QZOEHZgbNK/bhXTr+Sy6ukSrrLP3zxdE/5JCU1kJdzvAo1RAIv15ZTfC4Rw+J
XIRM4sC0urwupV48jlB7VgmQZeijn8M3HRtzFZkfn2P68ilvUjNyVjWuAPStgYOMsV6Fh4lsJAdW
88rPHoimgK0Kjvv7Aa6rLkmf2jVmCDzE5N3zO+MC8rJQAq89wvySJj7dEBR4c5DI3m0Ii8nKKVJG
wgSfciLueEI8FhKTtQllCFRum0j/osS4b6hhWYjdLq9C7Y8uRfQKSzdsxoD00dFcX2uOzA3Trf6t
Lh3NM4GVeugmgSNqpnm4wqRfY7m6gXg9lFaY8RoukfSWRTOnLJ9hSVi5CtAk4m3OUdyoyjf1oiZK
oMLy01XKyLvL4hcBQXAPM7GYJ0eYeOazxnrZE+Nm/NbkZJGTnbFkj6aB9mnDoRpsCP56yo4+t4rJ
4PI1WfpPgHHzc9l9D0YTfvESYS/cK49lkU7SgzkyHbtRY28XeS6iXzLTAWKRuGS0huO1vYQAE3J2
PNGp9JAiQgoQhOfmE3MrYobhoucOggXLMX3DrPfm8zBqSYqonOBmwmt4y9fBF7iB64GvxzOURolp
1h7p13rht7aCFi6bcAo1NCXdLXiQoEat2Gca4tFrrZ04+nf8V+BY4kWZwV/LYlU+3C1LpANDq9iV
xkB6v9bXfGCarjHDKtmeBhfIVUT2MHTwCFkTLeCrxUyfAbejtXNar9yEDTmyE8c+eI58EMdyhvWp
tlrbJ/Ci+x7937hoWzkC7E63OztGHXc+u3RIQEafNVZWgAL3Wz4pxeN0G6EyOQBoQJFcJdmPe2md
ERnT4Og7acAspH5l0v81ZtmWQPMJ4jO8WQIXbRrqyWLrsDpJhLFU1hAtgkqCm5ejzTdBHRO/xXZv
YmY90NuR/0Lw2uq6CxyEeQM+Go6YBXz3GDumsn2IRWghBkcutm+jyUF7x1+IgVfLbt07ouxE+zMP
ELq0qp6ayni1rf6wWJv4QF1PvZPl6GbECngvWR2IKKxNcJnKPxk/hIJWh7IkkNOEbbRrX1R8X1wb
XKsOBhK6k7fUu+2P4VyWdgXcdAb6b+EeBI0u9J03pzVGAbwrV2htqn40wB0RXxhO0t0NfTIxoUJ7
Ko4PtWQaq/FJ2okmPE3+arW8fF4GGAjlT5SQKGdhUACIae0u+xAPX+J3JjxOjEXLt5f7nxXSfNUX
25uhsfaiTp8vRv5nd0Tsdp1zEU5MCsn6xMj/rOfsQVAUOzFjZ7NKrpw7v8NZGXJj70az55sC5Ehy
KtjEUa6pyMJnxLiSgzMCmAZ8yUy3Kk4tLJUEtHDofu7IqmeSLJZcNgkP+BF+VJiHgcIV6DkELEeU
SP9c1Lw208O+1ubKHgLtXKLsw91PBX5MiYJly5y5iyQJpmapN5ExOT916wYiJMVHXcId3rDc3sZZ
+TF36lXy2men77Xbg1qEuctRGhnBHec4kXrFTgY+/ILRPC2OwsV2vLDTOsLXCiCM7lc7hA5BqiyJ
tcvB4nkafPyP3Be7VorSugtvU4xCKRiySS/JflJoZC9a8q87tLrbEbj0T4P0iN4J1HsOzDXmQioi
v4Ipi8yKu93hAQdJnRn5+jPJE2l3esPAyaZAsOs/LeAahDa5oSSgkkmR/th9T7t3XWbOvyDleA8Q
EGaaV+uJqPxpJ6wBaNJvGRDG/RWKoOAXrg5dhtoXNtXAyOwJGiGCnwWxm+iby4cRSozY5OkZqrCz
n9g6jnWhg6d6Gf4Dvo8QImcp6QsjXgsSAtSjzUevEGpiRKIOcCZ0cpnzce2yz0/Hd0GgRoQODqHc
yEJazA26HxWZ0Kpv8MEASoFZYPju66w/05M8maUhN9naOvvG0YvGQfo9jtBy03W+sK2gsvasf2C9
xvP2XMCzOX0vvSqHRe+BB5bKsyEVLXMuYhuzH0NS0a8jrQ/drzTVeDVoBnSFU5F/RFSMZ+RR6I8B
bZJmlrk2mfhPoWbwVMeafwTTwl5ZGZT0eAIPzy1dkV8x/qkQdYgmbO6xOShA5Ck6+UISjuz9pze8
cLE8yLegD/NpjehB+ZA/9cQ/7Fg7mPvl8NbPrUKDEElLGb+y9Qe7FjYxBb7Y44UIE9Eh5b/Tk7tO
lru5XjFDYwinhBGvF/xMrMh319m19V5Z5s/+v9gTI2jrIHEKJfECk9JGV+Rw21H4JV1MiWVHB1y2
k7NaUpVqWdPvuYH9671vdWRzlbcBuJG2rom0vO5aeuy2QEtBcJwyUnPt9WAc8W/Tv7scxRnwLRje
fFBjNUabcy2D8203/Wi0OVvZwj2yzZLPhtFitwteo00zkgzMrUB2+ik1UNgs6BEbe2U1R+2TaemN
+IY7rhZr8iOaIeFes+OyvRoRVedFWP2y/DeazHyekFHaF1zPXt7259/zHR0KG39k6kxlZ7ndTl9F
BmVnAXY9DkleC0cYggjL/NsonXRXlPcKSPtWECjjI2hy2RqDj89akbjG0v0FwqvOtWNNjEbXkRuQ
p9ei4i45CWuTm4EKeVqxCldKKqXPV53jZDj3eLH3vTdt0qEY9x7keHJPysY2G3PWPKFdiMcel+Uu
f10wUOrDif7cJSuFh67N3k4Hxthwc3GJehVpOHr3nhBJul/4yvf3Mzm1w4f+NJ8eaFN07yF5Pbed
I9HrbZmpAUN9DiWqjr6IbStcMzWc2XgBLTVBEEFseJIkIo8NHux14h5e7hZMp068lYSv02B3IwQl
5KEHD5MREU8Xy+yEv/BG47C0iDR7PTV609fFKUNKtdzKre1aK+excujZ3pEuPLa2ehQp62PmYsBj
aLBjypE4GACoVp5ja+wWi3oa3z5RiNevyv/vqsVfuNKY30kKLY3hUR+T89ZtqvgmmsMYSn6xR0QF
I8YFsUm1lgSuari9xPVGF89FdUCVJEbENCiDbeKeNz5+2JQG+MKWWkjqEEXiNS/mSvQ6+HvDZ81U
Wj0laKuFWITuqcjIIAF5KW3u7YsFCyprdaGrtlPQ0L+e+Y28rwLJo0y/kW9UFoMCzqiUTlKqkDli
V+rQPGw4kentsTRjcgFj+BbX6AoEZENy3w1rsD8vQgF3rTFOq6/XGpluOisITA8nmQwKM5wPq7Ew
L+o+OwI2lYGp/fzt5uvFwi7w3DuQwJiNqY6Fo83obpBSk02HbUVQb7y/Un8CRZfUqTVjXq5LHa8A
i/YDMjIKfH5O0klWRLY7lppVNgrNdPSX4bV2HJ1y7kP+JmBBF2fyOmBUBJMr2HU4mPpj1+a6SFUn
pN7tOAv3jdYIV5BBFsG+xUovziYxRbFTxEkzcpL+e2AvSjAoqczXfsTBVlwjHafHrewgR83SEfdg
XHN5+rLQkBBJlpSr1a6DJZlhZlIGa1b7w5Xs7qN4qT1MNwN0hKvxWXXmRl/U1ktJYyWO/aqg4eS0
HgToxC3T+z1xdugCZmn3aEFXIe1IvmJZuQ+DufqrUngvYRG6RDSYHMBVkpsscsytpTL4QOW2eBkt
xUFPn1OFVHzZT8NOfD5gpwiut0Pp0u/a6LwTRm9bfH5+AsM/ZVGsrf1eTgmZK5sT11mNriD9ZZZU
P6mVfWK1zrXkA7MJDGXcsZakwM8HnMy9iYrFwktg4xYLPvpbL2BUhfgVVdyDnTXiTL/zNA9LKn98
kYApImmgikOjSt3gLE6h5BElidzjMKR4PA/abviMm8YVwjLY7u2nhOU765OAjSdgnj+bNto3zjDM
KwhoBITY9gZtYsQ7KC3wIKDi3utVYsOKK9JDyUil5l8KrLRD0VnpiqgSbZ+OQ5biUHKRrrd1bsFn
3gRkrRF8JaBPzLXiUISuxiWu9uJp+hXeQCAf8pitcxVa+CPVNQCJztCKJh2PgyjhzBCMjKLm7uRf
Ml6Cersd9u+YUHLQYNl9u0uJ/bVAdJKmtCAY6To1hu4rADXuM1wBYmWXowrj5hCwyIPEXKVm4eR0
2/5FV0Cg3Ey8hAW1MHfQWmY5+fw8s4wGVZoeosv5TS6iXNYX/R6bRuq9JfauEN6HfLjP1TlDT+0m
rK8ipiZLOrJv3XZd/pbiEu1FX4l/OeVwY82gh8lKsufGwAA1AdVKEIZGMrSXRLc54dy0EhPlmFAB
hWOlztc/lzcmaXUVlouaORSCXBofyUfS6b3Y2v3k00fRo1uJBICwsxjPizMCNVHZC0d4KpL56oF4
SPraAskWpO1akfZQA4b5LZ40vZBnvuNKdONWbZXRHRIgMvmRAuExB9+YDzcnypfj9QF6v9Xvuz6b
Z4UnwnHwU4i0CIZHj1/zF38njeq5GzJt3jQMBo2f76ND6z/xeus29bkiZ/n/7igjRnWmiyKumKKS
VEUS6tUxQ3KaBpuayiaaG+XM/5vj95Z0xLUrd45vkD8OWjjhtf6eMqYkTdOkD/GxuXt+aw2J7G/y
RG1z8Uv26UOfWZ97Y3BGBPREmgQaS+aXJsnCND6buoheLeSRz7mNLHvozN5ENp6Kue1kWmKtjx2z
/S0n88ZbydZrkWHA0HkrZOZ3oQ535Or2FEMp3mQmBPPbWK0oVZxUZu//TywktdFRriSwVyqxzADl
ST8dE894MpQ06ZJEjMh96kCpjTteknE2SIrZrqSzCQHfFbl8Gy4gfQ/fADCtwrY8QdjzTGNSxCsv
sPdd9bkaLNO/xb08cNRRwMzyGsfYHb9e3zHYMIVwDbJ6emdM+rUlmYZ6SkuwvBDZfFi+Tr6aCgc4
2IbJWg1yjBntppl+4GG99Vayuf+NTjEYL2ZlfJIACqlLAg8LcqtDvBV10UHVZuvg0p4FW7xndtYt
6LeGIdWcjtR2IjQxgH1eYmR/Amva1gA3jLA/XZPjrjL0LGQUWomtCbgJxxxHRokvkZ2qBuYH2ztD
+DRMyeDrcTP0rknsxQ06Ufwc33tFfy/eTPlvXEB1vcn1GdsPFPIFAXvbHkH8DtssLD4mdW9oksYt
2pQ6KqFpfv8orDuTCEYDjDFNikfyQJdrDfBCIgWzENDDsbfV+GIV84MXf8WUWMREp2IvAiPCNPZQ
KRuamGGSQ+31h+vMTiw+Kd0HZLNslELJg9/fe0XsW1VkC09cXsMrx4wLB9xvPKx/wXuPnbTNNp5a
ZuCr4PYlJTTCCXbKSQ84DPRIr18wWZkCf28UV1qn487pXe3QZQ/OIifVLAFNh/zG7l39M4juPsEB
np8AHDsTOdptJWiQeX8O6SHg39gAWrFbXtsy4Zz3orDnfI19WY5nCd1dly6kjO8d+aN7BxqkcLgZ
jMvRKi7QgNv2EBeoUoKwj9k0ogxLdxJXPXo0yDqesVqc6dsF8b28el6hBI/pN+0Aj+05r+qAqmSK
yYHYILqMF5JtxTiXrY3/qrrs8iF4jNzpBRuM3AW5h4dsr52t8SGMyemARcMb6QIb/vVfgcDBGrgb
7Np73zNIXCvJcajC1OxycwIHHZ2DuGDTkgnNsLzrad4FMtgV5F9AOU/S6Otiwom9O2EQHgZu6C1w
OrAyG5oTLLgOANVZoVBskWZ1u3zg6gKMOLnNAjIveO1v4n2QlGppZc9a0SQnR3YgTy1MEgk2gFmi
ME9iMxNzvEKm6ZEiYi0UPyiYQaeXOB37V/c1QExi+xN4CAl72/+Qx2Q0gXNLqfJPA0kWZ5bJA3Ww
Q3YKv1E4Xwz5UoSJdkPEZ2NRm38Wg6VlPG/JRYLd/jZaQRz2fZomH5q0hSXyTTC5Sl8t0myDA9Dd
KCyWXa7b/IglE1J5r7Z8HtGaFMA/TPvcMD6frK7UprO/svS/JuOxMw+c29w7IdfVYZlu43m+5Np7
KIjV8EAXZ9TmwqPpPB9+CXRzJHHsWU7jGSI1hY1FJ8CYqArkd1vsYrWZIjxyTeDtWvCPixXrfauM
zzsfEOmyQiSwrxRRz4pC0Q/2ulHeQFP2Qvwd+gv3jvPvX/jb2v67fQov2qFfjqdAl6EzWUsedgbx
qfva0slMyl6NBVZr5O2fse3h6SodJvmFRVdL85EeNJDpBLWKBnjkp//aXcOR6XoUeGG8AbXb546D
GpmQZg5TljVWEjvZnFxSSTlSGkox4AGEVXw7qfbToVXrT3HKZYQ/9ntp0Rg9Lszo3iiXsqTk76v1
4mtz6EfmgLjTw36IT0eiTPCowHvy6Bt7a+YlyEzay86sMUh4/0Yota1gtNIxZ+urcSDeMIsh4LtN
EmzgiM08NPkTFFVF0I4icLuT3MgI7P8WT98geEEnnHha82qgkcN04O78XZBV1iqyP0nT75omAoij
LlIKeOH4SE2D34KZijRf8GViLJUNCFb9r5Kb0HlOraEIPdiIZ3acNdCiG0+OWRiEJ88aobgiGhjH
n8AlDN8VB19snBPIlNN1MxZt2O7xEIUZYCkPiP20BxP01ZhG/Ta3VR99IRhFdmjfbWIlG0GSdy7X
mJvcurgtrocZpvFqwpU110zpn/FIOhoXzuxF7DNghAKRduaWOmzkeT+AbqXvXdF0Nl8nN5y/T/Xa
3QvkiqqqL3o2Qwji2J1ViTVAuxuWbWt30VZfuyFIflf4xXclH70tIfHGX5XoCWVnPtOAgbk8j01r
Fr5rM32mNrQ/g8BSzO3y7AqChTlrqwx6MPOJknHHDL+TFCcSwskEN1lXXgjjCL5LbLJGAfj7yGQw
8EdW4Qhaws9wvZOCTBQum4dmSd9ko/lOszDwt3rur8JMyWbBCLM2BsC2rv9P7LefxYJX3xQTRKca
NbvHhEWTRHaiqyFsh+Fne25UoCkPjHG3uHbooVmEKCCEWgUCe4gwJsrS+iYmbEUiq/6vjXZ0NZUg
UHN5DPwQBZgjB0O3Wa3ZDGmcbDvPHqk4ASKCZ4KA4FAaL0uwrCNoNMpQV2PuyPObqmU6ReqVnpau
BsFwoCjFOwj9PcvWSlSybJUfvTq63wiKI/I5O2U1X9+Tu0K2FWXvjZHvRxHFFwML/ooP/T0/iBU+
1Qj4MOvATaBQi+DIER4JSnyJhe5axzJrRWdFFlOOwAu4O41kq07/eOE6IcwzItlZchVnNQkQ3V+g
JV/X1Ak7+C5Z5DebknF24aPuhvnqMnAih+koHXBhD51026Gra2dt821ZmOxaTmAVtsVIyDl4jjXr
anhGRLF0coI0T7Bk+bYkH2R1Tf0g63p0Cc+Qz1S4WegofrZSCk6PPODU12bS6BNzx0SHEpRAaKc+
c2O4JgD/pywOHMzOgslj8+PBrfFKZ5Xm5ogA7uYlH01b7bUCfMa5H7pOxfoaClFe9czfs0hie943
UqArLwIsZ8fJxW8fCwRNy0sDCk9uZasvq9hGJkxk7+TOfS0g8YkyQecWEqnqwrmzY4ZyDPsVEoTo
eTQ3Av8S6RXPzv2pUn/cnnUpHZWJD3F4SiP3LoA9MKdM9n6nqO804kE1EPAPGlKHF7EtkvtLKXzV
u117wc+IPtNXqa128siRhzFxk7/B1QHVr/P3IG6MsPuURARMdKxyhZbWyswl0VleJx+M8NuwbfJU
SaVBAknUPAHj0l+GS9sF8EovTIU/jZHF1GWfjOobsXWUeT4b3pXXCrksWEgXDcIhKqW2EQcFYhIs
MffCWmTl9KziuiE4yhB3IJfjbjvwcHYD5rGYlYrFsbcCDtQVT5GsarSFqUEK7NOeQjr8r/TJ4+bz
MDJu+N5qTBpFCJrclyMKOPAXeYy1NKzSz6YbNT1tnHnIYYRaS2o44lzVOPNW9tS8sQRINgRIx7Jx
8T0LgpIu6iL4dJH4ISTfg16ZgY7O8tCV/UTAF9XvPZ9s59M9trrQgkdSDuuYNkWwIok147O6wQEU
M5zY5R2A3SnVkLodrP4rKRRWQ0978spJZnbHnmhCr9tJTHOMbQpKHL9Onlv5r89AjEQwIvB2yD2N
mHzIzqdyDe8qPRO6ukcrypAB6gP12zqA2Ir8CQ0ZQCCjIkpCjNR2vLGr3eMk1kumI6cepqzC5+at
SF92ruTZI9VMOXjCPcO7qbvUBIHu+NtRfDoYc7N5HFCwQMeGDcsVyh/uvHWjBgiHE5Bylb3Bv0rs
s9WwGZaliADDfiQdsNTZjygWgzIpeDnSmZa1fPbrKlDnkSoC0iu2K/dUPFlIxzdmEAmwGF1mJcLM
dMJWwHpFTNCnMk9b9kVDLjRJ86xxWqiQzakpPplGJKYv7bAUioCbRqRINf51LXwO6lXJc7F6i5iu
DmV24Vcrk7wd3yaUWJ+k7baz5RSST43/AT+2R11ln0SvOUcbJW+coJKNrRY1fFcEm87YblfaQFJU
x7IY7dclnkUhzRSzRyUiwxOpgwdjfdVBTXuGWr9Z6xZ1N8YUVbdhdhGe4dkpbv8CNfO2ndUoHFpx
+8qJTV3/S6wQUPw6mS4gWi6nW7s5sFCtNwFumjIXGK1Xg6gRh6ZaksdQ08+6I+Wd/qaWgC/kG3VE
0L2s25fUwBXAB7JBp7mB0EKoFmeONdIkzgwQOPQKqO028LBtyDWisCfouMX5m4mEe8wsyqDjaqSg
h4snXSDzPFYjbKnnfYpARKEBg2OGnWhBO8wGlB6/rRvcjt5bwqRDWOK++ndHmNVICU+ifR8kRU1R
htX7NfgRiBp9wqJGOYs+CuXDHnmmyT5wli9dJ1dl/k1gP9Dhl66qogXgiiUEM1GfXibLihi9AkPn
OI+hGEXtiKYQ8kV/2AdiDbEXscUkgLwfqsyq28WSkWzxMQp748im7gsdo88gsRkRU1b3Hd7MIXEU
mlApM1hl687UbM63ZwzN5LbPiyb1AbEKVxhCm111yTjICgZhPPrYMJSv6hvhvVX2RWgSrm8zjBzp
Q3cyTYjWDvkyERP6GNYDnc8IPSJKIcFJXuplxR4JRrK5iFNGWnxv2j7GeH9nkYGifZ1gE7tYbAOK
CWU9l+utDDYfJpq1b/Dblk2NJ+mt4qb5AQb//r+aNjCGPd/0zHb8ZXYi0+H8YGX5FNghA8NmzINp
hy0OY2x5YtHdyT+nAKG/fPRcV6vjGfgyzF6D1PySjsdXtD8Le1CIcm3yrCMH+j3bX+MhP3Y3jMBJ
Fu9oG+j2ppuvag9ZsMH1gVQ18bMNyTKNnlL6c5y+s5S6Y/IR98HTAlMP8Hh+6Rpw4eaVRiYHhFNP
8j9u2/Df9tnMUMyZu3vGl17mK3zlRJMfw/nUeZ3cBxQR9o1uHPHwwF/r491fqndoFX4RqXE8StrE
fI+B1YjAmlCJvCTby7SFbulmz4JFCWXHaNpsQ3NpWZVBSGMRnmbPgQuKEh23BXd5rSoe3lDKtJe5
29i1L4zLzigjcFtXxt5LK6BFUHcUehH3Bg5I85J1WQ7K7oxoi/v5GqGJD4apRlVwF0vTWAEAv6Kw
fhAm9jG0eKJUPMtYHCy22/KjE0FMojM4WZkt4Y/CzlXAVZZMDmGPb137GrY/5yg0k138GuuKuNhT
gJ7bJCLU0/1xjERdWYZalKhBaQKQUdjdBT0AnDG0RoKGto118wJ0YM511PmkIImKDvcj9la+Kcg9
6Zoi/rYqF4Qs/rUu1CN9hPGQO/heCFQIkS+h+busJSLU/Kj2BqG1MFqVRxj2vICWu8tuI/up7mLL
mf5J492lZ0mLXRhvpUG3ReZXhfikq+7xOya6kI5OCpaTEdUAfV1E0IY+XtNdvBN3pP7gl6sYN3H8
n75OfG6aj2rhEPDSNblyf2rEjz1f4QBGhWYknvvZSFToWJb/BTFSOjfo3uOl2PO6eokqVonesRuN
UlP+GQGjBWEGQpu2068CAYNwH0IfmHpnMCDgslv89JZBCvIlYLc21QtpeXLsoRYkuihDkhWEGcH9
wYUeDOWdRIQrJmRl7qzJ9cVUvLtIJmL6PVjQU2/fyG1/pKaSd9pSv+Y9JhRZ4Wds/5aMSw2hM+CP
vTWmkrwbdJQgseCVTc4YvLumTcBfZsxTjQ4n+2wE1Dr3f2selKttXYO2qkKkYrMajV4luxtpNKL1
eZragRUGf8dqYnH9nI52kYpZzPZIEi0bkSNJx0woUfiqjvG+LWCh2siXY76mvsW9cRbjwfvwhxD8
wMEnicx8sLSRH/lDb4N0vSK1ra8KG8Me+iYkresoaC533IC6g7XwypsjFRe+x/tXpn9f5so90rNW
AWdN1D5Sh8XYybrA8W03/49jVYWgbVMMwr8zvTB6WLU+7TBqPhECwlkYwbu/uYD08E7PGDuhyPto
rZ64yLMDxpY/0btw6lvHzDezPAxbLtRy8e0FfwcpUU05OuM8J+ItBPCJyYE+dNGQ9o0NbBxFe8+t
gaKe9O9IRPFwxdHVqM8cgYzHvPaghYam7dccDlttru5UzDuMR+3iEvaqy1KxnB1dTfv62VGNLK3F
urr6Pj95OjIe5QF+f6Z4Ti6D40UWl5iW68wQAOHSKwjN2r8ucdlG4EhUjBUn/sufogMaFx1Lpe4z
1T72y3upQ020d31DR2q8EA2KyOJszOirjpkZD7Cpb8y8HTa3kfmhjk/M6egSIyjG0WMCDRk9so7D
wfUzeYwi9mittmdQQ6pzMghtvibV3Oh0R5hqXtNPDB8yY0Ir+OCtJO0YE8aXunU0eon/dheRjceL
HccmkOwyriYgcmQi8OiLwBfmVzR/ogEU/NHfscsCBFKL9SGyORFEtqJ4eY5IgLhU1gGmwJjR5aFG
6rTtLQUud4Ee3auuE5O0HwgN4eITLBcl3daq/G9vwj0OkAvU/f2xAVmFaFTinP0U1ixxsnyMvIGp
PXQJ1gFK4Sl2MAu+3IBDCbH52zZc/F1XzBw7l6ueb0rB8nirE6uCwGR8Nlxi7M+u3o+BwAwivebB
2G+3/oQt2lRjO8T1Gy8gPsLn9YvQNMgod3VzhxXRJAdvaMqEkTFHDO2CW4bDFMU0YB2l5dYBfwm8
tIS2DjC2tA/ah1onb8aD6hh7RgZehYmVSG10UVQ23W/It3M3Wm/47xR8imMlTI8w9UM+RNbx4+95
MTh6GQvd1lcEWl4IHqcq7vKWAg1ryJ+3RTMQiaLvNRzPk/7/gh3QW1O2PUF76t1Zuw91A7F1NQ/f
x1bKI/Ahp9E/8wY3r+y8ztJsNmXC3pBMCF4XHjuK9i1MspkRjkBjUSE50pRB/S//okI0LZ0mHVKw
HYpJCoCuHguUeERcnSLpfXZ7hEE7GZxmU+qdye0+nvy3FJigJsOVW0XB5lgZR0OazO0PPIy+ycW3
itFxRS6LobZ6isngo8FnnVCwQp/nn4H1m06OycL/ai3ZDX1q8WgjMbfYDH2tvYITk+2Ne67w6kSv
XSIyd+7xzM2fa8PcC3rg3yV4/yB+90EjlWv8Bka4BpDqkWkW+eHPJGqVcmazZwq0p2d/rUhzfyda
VX8lfjxTNhRDONDbqWBDS4xCj7OeeQyKi6+9vn/oZ04wlQl/sqRNOiRJAl2+H1W0eAkfLbiFsSw+
PWjKso7VIo7qK8Bd1A2bhbmss2fgbSAUkxg0aAsB+r42GBbYg1FVT0TJL4CofJrTM/Q0vpCYbzsi
58LzGbROgFwDChNnUvHqA6Y+hOHklrYXKaOmc1kGZUekW9MqRVe9SwGDYNufMRKdufIW3DL+MGOu
yV7zYYQAbhinmzkic53lEkjvJ9bwNA1F95aV/Ovi4MEB040oE4qSWQhTGMI1aqcpvfc7AYndsSJE
Qt8YSidEA4BZ7DMW9beYaivdoom/YS8jpUknh4Vh659QzCVUv7hNTzdhU0TsT3/pwTwbFT2d5E0H
kwX1Pfr46xfaYcw9u604xmanwt+p2tAN/6tXUaOQqAsUBxJzRBMzvHaB7vlvygLGuepH+XSwKq9E
qetYyfEuuR3vnlUkhkiLzBRGEJQ+S8/B+NzvkMiS/6VycMCb7zJWIVOoxXVBtPTSPPWtmW3xGnVY
Zl5vUpDzbtLDqIrI5efFuK4k7GoIiJepxzDNsUUKnjAvyO+NgUg4moFZE8QBLvTN4edjM7BVFhZj
MGssaR9ICfXAFw5/5JbXiZi+DCzAWX/oIvBvUKg6lfmBoV5oFkY4heS1faFvItVHURMfHveJmvXE
UsRowWDfJAZytFXV7tHKrEI4kLUhYXZa3ANn9Ie8y0nsiCtGYKOsLF7ApVCu+ri61cfYhu66flff
HuTc2cM/W5Cqj6lHI7ShgDEWtNXZbvNL5aFFvD4HTF8A7RPpewv7enXhFtVFfF+e8F58mAUc8ioI
30uRqCKd1aXGr1UHhUZN5OakMTlpnYkyKfLRyzIOqRZqnjsiI86gScgifVPCakWrqHCv2wcXn9rc
3jnbnX0vMZg4qJ/xBBJ/Hr+gsdkr/adJ6kQQxoVZNJ4dRk7Hj/YBm+jzxuEU6rr+cU2EA5K0Sd6u
Dg4/P3mKdfX5775uzpJND9YmyY6XArP4L0xHDMkKj0Ld2LSnU1IAoi9xRuWvZeDynGqpZRTO2RpK
x7sOKA3rMg4BsKsSN7hrulfVa8jRBwllli0rZbKtS3DNfqmPDa7qp258Erf3aHThIRqIVEocYpM7
gwkPji/VDv+++sSz2XtO20BlbIv+jRp7bsmZug4d+6X6FoI1hoR37+XaKLX7dQVDtEAPcLoxPula
Kh22s1UW+uUXMeFgmsY3GU2AfgkwmGaJBZ0Ij9MRWss1os6VL4VnhaWDytLdIOkG2JkoxCpbZc4z
j2F1CA0dMZE3J7JBZ3+tC1BnaOFBp1KL5LQ2VOjYOExNeMzp40zY3V+e19aC6YBYUXEezEva0eYr
+pnkda1gQS0aISruMT4vlQjtx4/kdSof58CJcEEFnHrJJpiZ58Hse/hnMZFSu2FuhnpJvTvmDVs3
yY6YSJqi/JXHYMnuchiwx0hxNBxVUHS0DVh2jDJ7I80SDxSCPxma7oWNhCO4pRWDjSf8UrVpD05f
+LqiLwGy9J5kuxbEK5ViDixEzO/SCpLqUQbR4/Ro+y7TQKusWDkFMEpe0bWc0ZROq6CI+9vgU3qO
Ns3JT13wKWXJO2B0XGZmTbzgn7lkY/fwIFd11yVrbbxOcJtZOFQbnSCRP+jibb+C/XaNXVQ2lhPI
qPyWLzVkn2O13xVV+khi+ahvDe7gjj9pMZiBJUHQFZOru30AxyQTpfFie1Hq4R+JQj1Tv8f2jWQ9
/wDz8z7xqCl9OKbquESIpDpeJZrwGcUnsa3SVaXk8m6BpNlMJxzgndzQEIhJE4EhbyIECavy/axf
lNW+ztHFCfGUeF+JSluU6cuKj7UFmr0+yVLUUtac0+VDLyeFpijLXU6SQEWMIzYKECNWmoPNHL5X
lDrH1PPYqm4AItUTFi93bPqLjs3EbvsOBCHepOSQXuul+89cXTUs2gXqoVgzQKQhlfHaU3WOBtOg
v1HugqLdDOY2V4I9aQTpNJsNPW00qoNL3ASGfZGhR5ozS3wYSEA9EEepvkUOiQNCBESvnhbvNz7s
YuwVFAfs5uvkLvmePlBeSPDvgQHRQQv68OrULUJiutzeTDq/dSmSYkqYg0O934LIEZeifJRtpifM
Oy4fP7yqT6ciwvJXlosFiKOXB7PiE8Kou8wHW0t9uECSyjzO+nnzo6mQ3TBy9WEFnhDNVyta1PJU
JuvQoedOSMB4tYwbfc2vELrsm4og+QwQIqmSS5x01KnqhvHwn2EE1hfIO58ut5Lmp9sj/W7+Cu5G
bmcNDD4M9HmJ8zrOcDMEkJnofC53O7+ESEAf4rQeBB+NlaL/+3Jt7VYIrZtHVLNKq99hsaoqxeNd
VkzCQLt+e/wz/TaSutEqtdUEQah991e6WsJORtwQ6nA7TZG69PyH4v938RWmg7C6+mjeff8Iri2J
zY8MCdemZ0iZr74Q3vLFiNDsHT+2alOQMF4JzYZjAxQB6JmW+k+8UdDcqCNHYKg87jI9dLm8OBDE
Bg03o7B6jGilBXyqU1X/oa8nH9JqiHe6Jw0NhZPiQCq7vMxX/vptM0/g8Bpa6HrFZ3/s0xtLgr1y
QpBbbWLXjm8nO8ZpaLOBmFerBjbDeWFI+hcWbzNTN+PvAvWTM/E5Y4njgbNVZgr5KypkBpeIMSvP
/7H28/bltbV9uItefTAYMXgO21+0eHIc3cKX9cyo29kSyPH/f9vaewbm8eT6klXJ9ePSjhggDmdp
RcecdCWbop3bDVcRW7zNM4mJ6MnEHBo+rYvKFXgUISYul3w5RBWh7nZnczejaj6+KbRV8XoEYknZ
axG43/mcaIoNIO1nStLrqWrwa1cx0HdBDFZoc1O0JFXD6EKKWuM1EKjWT6wzbul41aMuIgupNmDU
xegb8EmLMzHSHzFMnaUfesaqm7W5RHmcIzTguEAUi1lwEZSVG8cRj/ZW2jW3nZgMtKnUKyF4qqvU
Ha3exDAAbRCfsqAeV1qYOIbOpK7RzTGdXh3ZApsvD84oJaT3diUaTSGFPfSJN72PtAZp3oASi7YT
PWDzVh4Gnzg+o6PWjno69KmzJv6Jt8NYHREiQ0Z2b0knccKYP2/CvFz6roQDy5tamhnZBalhn2jq
jdO3ESiWN4Wjmd0hsNstcZW4SeVVxJJsAd7ahtHWk959BDp9DtoLzCGVzyIhxjNy5qqmMwms7mS+
IqnHRfLNIvfAbdKUfCllKqyDx0+SFbp6VEHPwzXcv73n7XW+oGGY6e3Gcs6oUF4R9axp9gw4XrDu
u1RLpuKADkpyygCqD4ii+yBqcBWd4kc6ruvmN8XUvGVMrL7TPIlKQtdV+ekqnUD9bCWv0Z1j2X95
iLFRl8+uO6c7A4hVcV5Zhsg6fokLMu6BsfvlqsOAS9vPAm/n1+SGnV+HMD+800Ob1HR/GOGZ2Fb7
SSfGvb5o5+IFOROr5xIVPkD1y0qxVDZOyBaYqgOxQlL6yUY0DcKmxyhl/ygVVZHzj+g+wShB/pYS
pHHyVfYhK5bhursT9Vw8sCsBxExHpR2gkuni9mwopCBtPzxcsd13kH6+6zx7DUKaTqgH3VWBKyte
Paey6zfKPeV4dbUCb6oaT8yKCPlHHsD1KQ+AprkWnBU7z+PqzHtBweZazuCX4hiRTBEr9bOqKsvZ
5NCzbIvw27se0aF4Rr44HUEQYwj/IwQOLibWDvpcrEVYZNA8bwdwZ/qx0JVUdP1zTqGRTyzg/1sg
xO0u3KzTchJn2JaxPYXG9WZFivvNkhnE0LxNeYS9Nh0XK170or5l7QxWYoWabjP6MpBm8cYUmPvX
7uWmEyhQCeZR8BFHkG9ZJv9S6pwo8nsPavyrieq0W7oKzDV/SXooI52DWdPMIYM46BoOg0OkRuLo
wIek7aFyHPJvNEWnD3cNc6Oa3ocrGTn/wopiWlZF99ms0kH97sUhR5/kYoJOdb/pparBhKT0gXc4
wzuxEbOrf8/FYaoQo1OS4QcHAzClx0i+/4wchlxahSQIef+MaArjqVzDSS3LhSZVTkrGZz1cP52L
IZetCUJzxLCvLXMsObiAzuRPTVjyOStTjdSbuR0yJlvgHkxOoeyeODFMrzLVt8Lsxk+kCjf8HSc/
G+SoPDkefx4UwYW2V+Y01MQEBRaGSQ9C86M0nrJsX6Qli4mi7nXYX5lMlBBX5E+/DOMQrFRzS/dD
T12WxgBkRHi6n3kxhm7GFK2mWTr0xNNpCmG9zfJBz6PbM7UqJOFiOUw8eN0/G8yKeHbelCYLueKB
zR/vXTDtew9rhB53qQMNaeVIi6kjEfmi4aBiwyiwOpFbVW2GR4AdRsci3WKIPLZh3ldeeRkNRtyJ
OOC8VXMQsELLNQ5YLcqB52cG9QfcIu6zXYRnydLCYqX+r2GDaqXlIO+TwBybys1KypPcrZFA8ZnG
jcJ+wji2nevQOH0V86eukA9eEUk7AL+ciyOPa1hKti/BGMZj2E7CZotb9robygimiyhBwJTFPzZ4
MCAIS0vMYi9zWDBsnF+G1Opi5hQQUpSBdt1yV6jOTK7C3x/Oe9sxlSrPEtcNhJyhcnOX4PJ33TSa
kDmZwBHpEwtjX53VCtfKDzqU6pwlW+CaQvJTHnV0HQ1GsDhK3/dE2LXjLK9N0PO4iS1vV2x2whhO
rAFHgtLk02UWDskS6Fv5mVhXGKN4J6WpQAt2XklBYwJhwaqLtA74uxQmw2cKORupJQg9MJY/paRX
v/1klIyM+FzgnxQUEmRAydtsvXe+dSLUzbgMvNYw5Nzk9erfMNApMfXVxToMXIMbJOeieAwPXbbg
6gNushQe13/usjjM8xfDaWtpPAmevh5UF3QnDRRMhWs4HJm4wNaVwJFYJKbXzQFWAN/JYx49uurF
064spzCulYbokEXeI+YGMtqx9nSwkARxxUA+GHgC5ybQoT17B+UaYsp+OjMfX+0UWDfXjiUs5/V8
MY2YTrGFsNGJDnhZXuxgDhMb/A1Uo+q42i2Q6iLN7xnWxkd89gDFD7r/Chz9Ja1MiMdk55AU+oFS
+I+0xq3JdrcpFF8xwb8vc4OUbEFR271wJbixvoea+lO7ULBZC4EvtDbGTGJk9PM+KGogZ06JTk6o
AyFMCtgA1B0FqnHE01wQyC5Os5rUFm9SMAB0RBq3017ev5VUMKM6xa73oqItjiLNwwHGDX97akgH
Wke17Z7+tBK+BrnNVFeBF6YnC6UnjpL/acD8tVvbg0fd7Hyz3eGLTZfmEufPrzknKt/kSoQ7HBiW
+nZeJc1bPMsxNUl9+eje2tiVLtPNDNMPXVp44Qlw80RjYChC0u6yurjjUYOR6OMv0rIXDUhQQBr1
PWq8d8KlBv/yTUn6HX4FpmJbVL0kjDFFzwltiDVTUqtdc1HrIMBLrEDEJqCvM0xF873fjWkFZSJc
DrcGswcfijeUcEi+dIwcPDo0zsg+a6upADT9/0AJWeHMz+hlblM71WH0lRTlDrlckWbvRaqXnBt9
17ExE8bhxHxfQ5q9l6uOmOAGtKgjiyk/HDaQjADhjoNvSAWH5kNCUPaj8BmcH4hhVAHUsCRp7R+q
C0A37wdS3osGf2suOUtWUqCz4Mi4uQPMg8/KrNtPT0OfHBNdZjKafZmUnmvMXXpBBckO6z7c7w54
BsPKR5btVfoS9iHKSTKmu+OeBWSt4+3HRrNhdZ6g2YtkHtaCGeopxYy5lkcz03U5nAxL0f3NLak3
zj3Ilb3REma0H4YglDVQPyUtWttimbaIfZIXNOZRtwS/i4eT2j4f+AqqPote5bmWJlT1wr4COStL
ngLpmUh9Atw4+ddKCAv0p7N/HOLA3N+HIULoROvGkUsC99ks/6RDgPbmRWQZwYG+2EKlBr7wqLwO
8R2M57AETHD5hOEpp/emEQABt6G9/iVG3LduXyuiEb9j0JvjNYc/ZoN5pLhlXVgxYDtbHM+6fN3F
J9pdTP1VTcsqEYBAjlenmd4Le5w/qxyZkYZJDrNzf8OBwvCCNLLmaF20mRl4BhBHu7BtWnHpxknY
KARh3GzirB1V0YihjIFrn3kW4dJ40B8G8fzheg9HCfgK7bd+VEV8hrsTClSVxD1xAgLpxYILzjvl
+dWvcehMk1+yMr8c8kBpvgNDfpcAL3DwrvXHoh9ShrtcVfbxkJFrwCAAU4UNf0BU5uUihm85UIRp
XbQsTeoak7MTz8PSTcGumngO2Sre9tkW2aGCd2ioi+ppTT+SJMylxJIv0vOoJyBN/t2cJhGqejip
HMdIK6utVwQEV9Zx/Sl1EH+lbGiai0RewaJi7oTUKCZDsZINSb0087BdrUVB5WPA7X5Ld1KC9SrG
7/cFYEm2xR6isdHAwAAb70aJ92A7FXFij44MsoQjuWfgJ/mB1N9nKJenjn36EF8E8mTh8T8ABaHc
7uC5x8wKgEwWzOXlKtFvy9PdVrIQmxpchqCVcn3n6yMLRF7x6hImePCEvK3lBZ2LRqjq0AQxqCcL
biSYuTjA4/us8EC2o+N52t78h9PG2cjqyCarEd9EmvHMw1HogaYH63fWrH8AvjHRHHv7pWaVVsQH
XnRJw12jSup/TskT0lMaVeY1UQPSuWrNTOB0I621jxF97tIJi3mkLQWiJvLQ7OmN5zP6USSvcF4j
n7VG0xpTt10LVocu64OJY7PD4jP0yEEGOj4kjAe/IJsIIS+hOl7fyh3r+GbjxwHnG8/kO9kcBxIp
+LzFum7CB4AvsK6NWsGBALdk0Qf8AJvn6kcizQjrgWfr8aGIGbrmdvIAU11jY4/6lA6NSo/EMO9P
DjG/WJk3jYavvH1Og9yJUF4ggQN55n2MHqoB10Xsfy2McinUXmbHZymq/fuRoQDy6iiDY5SmKGLH
znMsFvVWO6t55ZJc73W9c9p4gv9yCQ5QLpDhST3V3BdTcEXmxeuHNVF+B7L8i+UFGFb6NfjrucPe
ziipF0x/D905QYCXhGfRcrnfgKLmwxquQKkDTWBGrJinjbD+6ijCtiKL2I06OZYWtYeQ5MY/+GVI
PFrFq3wW+EUwWHeGEwLTO7h9/ZsnyDHXwC+AJuEFElZG/DkdJXNvpbyRssB9AqIHrc0K9tSTQVOd
yZvMV7OJef4n0NguYNCx6JDqqNW4FPEr80q6l7cZgJUI4OiIfuOnwdSnlq/b+DtYEMnMtkExxVd6
QvxKrpgj+eAk2Exfm64eZt6DRJXKghW2JlS/bRXjYC3Dn/ugbLbBdomY79IaJg4HEIVTpkd5aIz2
Nez0rdvlgtMwUGui139HMB2uTYDNJRQZCcQN/i9/0hkBIhf6ONUYfBffD8KffJH0SmfO/rusVQhs
+M8dJocGOxlmuvVOYDiEopLa2xLi3DoMJVS9aabOmiK6/0AifKHT7XZ342ti5/qJ2n2zEgTvmh5S
zkPhXAhGW2+Uur/IkMDiL8AZiBgpfhXThFZWkXC8nVV8tITcpymvmVudBwqzwcpC8fZsBD+bj/hr
GxmRhgUz0sd6IpPSdEtQ6o9mGbErebDDdzBuhpfWCo81jTL59Xes1Wauz9TU9pojWaCItDg2td5a
QpweLeBErV932nmlfgxLJxigM5hIzxB+O951eSKWGTCI07HptZUV1ExPLWjzlnf1ztmJvPjwS0HQ
b9PiZUypz1Dx5FzIPdtI0mmMsjv0PQBKHl2Jqacqz5JFFpxylQDU8BJG68JNXMrbccuBwedoCmFz
VkXi9jPC1T4NtGAoJoC6QNBCT+a3AS1ZADd5OcOJ57zHrsiTHvK3qAo8N4Lv+dsY91nTteEv924s
u3EhG5DaKJOw7egpuE3CJDJRb7GaNCbhPzgwEjH74mng+3kgijaBc48Tq0F0yj88KFZ0fwWaLV52
GoDfkTpUQXc22s8723klcfvKZNY5bakyPIJKD68QsVoo+z/SvIpMdk4fbbK877wgQ8poikakMb41
1+2WA0izUjtpSXawifGpo295kUNk2kDhXzveo3ej13wccWxIqtjiWob16o8ScEUs2tppHxcjzD0I
cJaoV3CsGPyRWPkpFkRMocisYq8Rzg9YGycsrYaPM131t0z7LJk/8QDK9az7HajDZvsmA5jii+si
QlM7Udr9otan7dLDgj/FGAav1NN2SxW7mUp9hbpljZcqyn4V7MAgcUf0hMzoHq1RG0TXXFg+lmcI
a75p+vygeANBYeehpsQS4h7ah+JI7OWqyc8CB8qEj8nqWwSBz1MMUrPDnP2bBl+0umYM5R2rfOXO
1T9vm9jc+5iC1d3xdSBAWb2uN+/fDdjM2Xv8DFO4fwg+QYyZJuHjQOc8rsX2tqNiq1jrp1aFaCuR
8PjPbrlKJ/1SOkebZNBqP+yAI5kTVtXloGiGUxPUeUv4KEvJpBWXlt4i8dArMlxhKDJ/9mT0cRzl
1oRSMeeDUtzTzkTPBt/I0hemBE4sa02Hdn1CjDVOBiZgznsbohozDmT50Bp52qlY3k4i+NslS6DW
oKRu2lzuYmDvdTzBxZPD8Ksoqc82821h0vr4uCcgYp2K/be1UFQpt8O0epy9xkM4/4cbf1EQbGiY
vbg8RiCtYmtIsoxIwgbSvKSc6P0QRrq+cdD1j2sHCufT3Bqrx8kEtCYfe6bh0HypNomAtJljIOMV
jZoqUeLoDBLgztt3lICMI7lRg8jVV3mrd63kLsI/CfH6Hi6UQoHGYoB20lDRnex6H29q4F1CnHDg
G8Lp5sDmktl3QD6XOwm/83N39aJWUu/cXZ0rrvsnmGEk08NXRUUVt4Kkw2jLqo/XvLnXGlv0k48P
EgC6bSsL3adP7zaue26ISaUBXrb9YkzWn527b7YsLhD/OLe9fNztUlFQlMYSm0oNuhnk++NAq7pi
mrR0AwH2ul1TLCBPOqx8Pp6bpu9F5/OTBnFuMGhPDWOwdUWePRw3z/vHhj9pmza0eq5sq2TFfu8P
3p2bHjxJ2/F1+yeHpGql9899iN6+kKM/Sn1H+tM9kUeAthnzY317HgJT5vJuXkoD1qlILHOFJaTC
GjKvKlqb1OMueLb9y3CE8V1XcT0Wu53h6uwKkx57jIc1DvT9sLUeQOfY6PTViXbjjWwP1cvP22Ma
8IEjCklshVkL0rXctIDhkcCH3TKXAP87ZchhV+CshycXnPDNnr6YLhZOEUbdZXL/hl7+jWDQiV1x
MPJg0R11ZIEfEehQqIsmsd6JFJ2w4QoZHwbav+2TPMm16ag+Z9BFJ3P1IcgVRqKNzOdiqHyPVCPe
vZVY9qo4dXbcjNqMd0h5W5Q6aEreFLzp3w8s3HAi1lyIwuqBZDKT4LIxfn/i7vdINdSWL7qSiufm
92KXtQE+8PcW11qSjc4Be8diM9tgEzxSRDTzaXSGO2rUFW5ZFdBaCmqhyu7kS/vgcrV/KGdtOicg
ek2WcNXeBuOLZw/4z758Jr3IMksUdW31jtcNdIQmXPWTsH7OYTTuh5+Hf6HfzQQrFbBcF/JHOs2q
jXdZefFOzWZUxbyjmO+y2+byMhXhDlf+HTK2yRWFlZnZSxiVAdQa3sxFucfxtGyMxWOvlpmaOh47
ZwPDuMdHvpO0pCnRShMUHafRC9S17SeSPbG2P/4H7ZoJDY38kARGMD2spYvV2aDPFWKzbl6SXyCQ
tGq07/JW3BnyWHKETPd1mCSJPumfNjqI7O8fOIttiqGA40CTmoL0ac9Hr35hKtKje2YFKiUZSV3+
JusxxKSEBhNy++WeYdniTu9PO+43TwjFENcAfVWr1yxM2W4cp2dBGdl4gkH8+QI1/yQMVWFhk1uc
M676Vh4s+U5w8LgF0AGi6Yi28ZUspTVnR6WkwqdiHHFAihV02KdZvlckdiH0J/zdRN9ECHZcXBr4
k6c6xg2Lrj+mN+qrwYmMMLhdxw8G+TwSb4vgfasY4huEs1foLipYxF5iAVkfnGN7rfwVIWEGzfag
vxc4TNJD3TPsSuaiRyEcP6BJVKVb9Tg7OAMFvc5EpU7/BOKj1yI3Ft87f2mn+3n+MpChaKDU03j/
yQhgUonHfNw1Nl0flaBvA0T47gR7Hog/pJrEFb8hDpctJDVyUP1NJ99Z1c8kGgWfGMqgYSwhwMiu
tF6ejQcwDJeQ24q8iJz+BBoj+kEm6V2DBXZICY7cFz5LaFV0keYDiITSnMcTyTvjCSDqpQSvhYXM
bJOwGbOOhIobEOlVrEVAZNBPuj8Rbp6zjck3V54pknwF4UEY5Rp8GVFB5pXmD4/jevYkcrubvfxW
hEMnPsYp6BU2Y5TpgX3b0HdPpCMSZqvYG9wwQNDsXkSMDR11ZuuGQNHSroDCeNuKV/kCLhXT2zvG
vikTAExsZbtDdXxk71i9ezsDw9pkb/yzE18tXiiTRT9qxch6uFChhYnKHLRpK5PTD77fy99P96oN
ytO/72ybbHatr3XI2NJKKMJ6L0x+pu0SZWY+QEqXz7aL7IgYJiFgIjKkqOxVpzeYhHavOPPl55+N
aO0r1e7+XKnKIy8ELBJvlX+YRDmWrw72YLBKUVAOCQIlqgwXUqmmcJnmb+S8nhhO9seL+15j+xAm
ZSMcwvJmjWYVXL46UGMBJNy99Qh7MrUcwPQyyWFg2K4SfLPDl3iHmIyrPdV33UNEeW+H1VnWnt+f
n6/VBDj9cBIGocORk+Sp6x+CD0MjNy5tgvOeJn5NE/m9c4rGDatAeRXPYFYtHI9RkqkQdO6mG0tU
UP/rUEIzsBYMwsE36A6FgQA8dqjHhQK1B+6RC85gFHAUBflYUCtkwsrRm0Q5hEJoX0xcFSCjxMY8
dFcKyBn60/RI78RC8g1tf7ic6fp8Uv0mzXwuevw0QmyUOKkuKDO0f8n+H5Im0NNL+NtjVkSfquNt
eCko8mm0d5sH6KxwK442ofdjPqi1/To2yd0lcVh5MpWL7EKPhGb00+uuzTMaAq3DJodE1LMyjEDJ
YwHdhCwi3scdxwYnFxr6UFFRh9KmbrGomdDQLsVXFFfjGO2RSN8biqrObN2YRPVq5uzGi6Xq8c3i
9c4kf2Ywsb7iq6Hg/HbhfRUKNByeKaMRPe7o2VXEAEVi4QvdppNtPE7xsk+1e3ec+l5ySm/6/laW
Q+TjoarEnbsvX3HeR3JmA5u9Z0QeIl46KIAWMFmrNE7xxAK9wqsJsTs2j59/axG7L9IiYFTAlY+F
XbfzE7PvGrcKHhm6hJYNkKqC3X0Puwg8rKrBVhTP107Bw0wK4reF1q2HN1Xlqd9rFvk+me8MIE1/
kDwv3hOeaJ6O6oLC+7uthGjadvAt249SNh7RkuikVqX/W+Ur2aEHZ2VK9NpfRZApQXoFq/0EJhWf
THkLb6fh9ISdcwkdGY/7RntE/lY/y3dm9FcVC+xcDqXadpRZQ4z4othdohyZpQ99XGFyXJ0/3hZY
2PHC7myHzPBZcT/Ng6EFbHhoQzZmYSMfwgaPms3q0MXkzYCt3f1I0wky91cDvRSrceLc5PysfiID
XKPuyIeF1XDRVUCV2O02I4rKu/SQysp/gXsVGpbxjSQQ0ZUlFSmgXRsTNzSLbaLl486zQhP7mr/q
2daJUmfBTrqqQU1/OFpcBjVIMOVcaGuWze4HKcPTcahmlGuI9GndF9fQol80BtiExEqeNHUiHPZE
R37RXI8FIIAHZ+O8iRxCJNWyX/ZrLTE/21krYTyBN4Kp7S3xOiNyCbgHe5PVe03P4C9ohfvQpO69
PoV3HtF5NR3Bxaauh1gU85XPf8XZWYOYJEEl/lel86SLL5KMtQxbXD9iFE5j1AZ7ywOgPmz24U97
FzL2e9Cw7M2IQ2wZUsPD76up8RxTxyJcowabRyD7cSo7bdYhJeuevlVTL8vfgPLQnAQVWjR76lWz
AnZIJrIS4eST6AKumLl/cgJrjhn17jSRpX2bVRn0K9fA3d4yMURbfdnGTUmy0nEu48okSbWyJoNK
Qx8dFFMaXc5YlaxeKgTVCSeacdrdMrb1CsWOVEuxgg9WFPAJSItrLR1eE7GmDwsNropXVVQzeOkT
IUqB43E1/sy/TXND+tHYn04nWMqrQfHQIfE8k4G5qT/+L2V39Qd1NJXvRBe+9UBJvb4lY73Zf8V9
c0uZDLi/VvMk8N9ITfqDQ3G/uEgIQoHwwV10JqiRsE5hGgiMyKs3P5iNQ0Ra423RWb3INJppmABl
UojrtBOLbNbtikaC1binbp/hoF5jCwQ0VAGNhpPBRIk40HdxzKyR0+r0gtfsgLMH06ILx/XSVuhG
ZXcBSWMwpPTbQXuunPh409F40F6O/bHnb8AHtI0PzIsfZ7pVjypOGnkxzC5zOcBi8l7tiGpXU+zY
2EpI71nKM0bGJh24XvrW0aQkBD63AHevgUAGvo9v/vgFWOLUrPNJLiRihR+K2LVi6GU5CEQy8S5U
HfTqRCrkQw1HFMG4Aqq7crT5ats2rtGPZsyQAZqW/0SSxuxoRuw+qTWoUn8zW4mXbofTFS1ewNnT
d4ChjEGfB1wTBSsxhObdgO2HogIS6kAqCBb1Q/HvW4UgY7Qwc7ZY+oc+qwdkcwXsXPn9jMBRPo+I
Zy5yCm+FRe5WP2xNmhYoXDOmXMtEVNeEFOGslSuyIxWVZHCNHGNxGyBRT70FqswyiOkJ9Bgq47O0
z6Qk0d9j7yuK+2pKLB/7Gb2OX30/oTlulBO9kOYWt4UqzK6+q/Tm5XSlCCqRLkKNmdQ6WNZeOq6S
ET3idJ92DnvLMWkM2eY1VmWEWDfCNBBZCgeRGlhVeW+UI5jrax1k10Q/ZiWfoKSsjC5gqG2kdUGb
wGCtyaJKd86ci4d0cW6uFGSJiCExo0xue+hbVqLgTPh47Z8EhWqsI+OFK2l04lQPZue90XnyYlXY
to/N/hoIrThy6JRKkM+HxIgMXd7bNQvJwmfjFPpTqxeyOp4taMMrxX8CL9jpmUB0FZPm9fGIs0BH
Sw2X4xYK8MM34eX7MBJyHExA0Mmj/u7gIixiupf+cyCJOfw4HzzHcH+qX/9mqnm0lvEjT77ii7s/
mOetS/t4339qQJLW6c1mGqCo1hs8qRjh/kRuVP+aWS7DRFo0SKciQX5KK4ubRlN84jbPm8Qfn23U
gYFdIImHbNLcxAw2CwFcwGMKVyuWCJys65d4h00nJEwu3dDrdOcdDWzjNZB/mPD2VhZfR+mAclKf
MYnO4x7Fw09TJuhLXLhq11MEPBOTSI3yPu0zWYzzHd39PtAQ8MDYjYSPL0SKSw48vFQ5Bswodb7M
rDuvGoZMiFp84ONBLVjQXJAS8MOpGafkAynAruZFC4XN1GwIJ3Oy/bxvIAt4m+BH3Bh6/FnH1xxH
wOTK4w/E7ZobsdMYKCHZtTm0jw+0nWyAkspr+cN6+5ti+OeoMUvzi5kn9QRxCsfB6rLzl118EhuA
eCdunV86J9G0cxrpsrj69ewwTccu9kx+sypBJ7dif5K29ERqnFEwHHERrsZJsad4ncAUnCASNS4d
ytP00vU3FdrISCbwO19SIdV52vlZJw+NLVCUdEFcBWod3JbIjcjMtiX3n1HYoYR8THj7wUsnWuKm
CloU/Kx4DNkgwfeX7jBOtX1EQ8Ao7ZTAuzK2XUWF/N/y8v2aYbF/h/5ocHkI+IpS5iMuQZc8zCJa
nx/IVo7o17XYFHBrYaOKsD51WoXTPjRdx+QVx2F8u557teNBOKKHCw2pwGD4QxnYbWEXOeN8/5lj
pNaCweU8QRjTyq90fQ2SUtsqW/MHbY9CDx/hCJWLRYgeFPasDjpMAXq9YJ2gLOerZay3Zt5jYBbO
NLb4WC4pn6PpKttG3fGTXz9x2Cz3SQFFmRz9LjsZPJpelSpggaRfXC5c8XlmRwlrUVVJxvoZF8Cz
YFOmImH1CSKLqgm+KaOaktxeXl5U/fLA0F2a6n9D/R5c+j8S/l0m/Ai1FiRM6p8igmQ4bPajJFoD
61sr8Q6X+2czPms6OY6n+syNS1Awe4+WDDgzYykve6ZTHcLDeJtXhhUewSckksMQG2ziWy42Z83/
xP1hOXSpht+DdFtf13Iyvf+InXotO+wJANncqJxUG0UGvdpQtBH/eR6c0hu2fp8QxKCw+6RS8KJW
hWxKGK0JUI/68/JY9gkgHVI1DlW3lTa+ixJKjASohyXrw9C4pPwbDYS7cvO6p7KmoKLcmhklcYXe
AxCJhuGmr7nfwbBGqxpU+XPnEZnPaSTyMktDuc16FFgjfBFfXYzhg9JFvO+7KYCCYkOAvEDTx3fM
PvzroO/ghH598WkcYLNUv+qbdged+0T7jDfKLCEyDQmPOFOKvqjN99l4J9Uwz3K53OVBxYZPRp8W
vGzDNoEymo/Az1Nl1jaXYfcSVFfW6z5wTNCfNrIxSHJIdkuDxokv9a8Qqyf4MrDJiCU4s+ZI4R49
VRYdlpqCFRN8g1EMXT0+5HtF5l2G9W8yqRugmwR36scJrP7hnvSFJ6/4B9sZsjUClOQYHtdOQDld
LfRh16+l9ANrwPWEfl/YDdP7fAAnpz1u+Yh+9I1F8qbW3sv0OfIJdlzWfWnlHlUGpNPw7SFc1NXe
mXiwkUhg72CNlpHpaxRufqoptnl4dVml6/q5dt8vIFvro3gnfPX40EJJ1sO1YssAhZtDdnmOfb80
hiMQtYYwjHxHmgVmtNlw2guOwOJVc3gm6bnMNrHf9WPjERrfvkbovuGaWt3wEylR2VBqNhDPbjmF
bYi80eKC2Z1RJ1FJSuPpUASuSklbESzZnNfbcOzwIlyIQTGA4cTJ28vT+YiYfQGFnMC++BOgd3bx
604bxwEcAWIAnCnt5qwdMbh2d7dT7pcC2SLhasUKcnO3OT2WPS8bCekuGgF3X/et1nrakoRvujZN
wsPLrY1Vu+iBBk4rHLB1YeHKXNMY5Kx9qAqUHNN0hUdn5THaWI5lovRZSrWiQ3U7opQpHzfcZtjW
D1pU+M81Um+VMIp1xFGSNZlsZP+dX3ShW9PuXvGgH4b1oHEv+iICoNITnpjOlUw60uK/wj8KDUA+
yTUVLEF6b8LZcg2TeoE9cEZa6+yaAmIKmuBw+kaRp1VbOruq/PKMMBxnfG7A1j9CDqffLXi/NqyP
0AquopaPJ4JOK43F1TZX5Mr5Evyzrfdxiczoz8MREL7AJ/MK4A+A9n15gw816nE+M9uEoTUfKsy9
WGxDX4lqhie62zOnsstbJ8L5KfrEfPMylN3K/P4feZlLoAsjko9n7bK5lDUE/rn8n5/BA85+inHo
t98yKFYsvJkHV6Y1LFS6BiQJ+ZpYXSXWJ7IUjyXZmrSj0BQgfZHgg+YNxntjrDtmk6e8hxpFPH2i
xvXV1pIu1mL3oi/LlY7EhH/DXlbNyY2LTRRbA9hwBPydZwXyIpCaNp0A6PKuYAdX7r/OyBuGrI7t
bRlzoG01i907hyo9cQWGQ3Uli6XXqrOcHK0Gsfv3w/DdCdQMFeul8cPqpoQiyYvd6vKoTYDi2T+y
y73cU84mnIr2vSSn6VE1EYy7OuJyPDLMwOFEyPdYCUoDoWgE85HC/aCfZtXp3cAx+mxXBX+KWfWi
F8rpCsbrs4tbcYJHPh9yeuxHewdoXwNrWpllF3ToC+Ov8qMePVnKF6HdLIE7ZJDjoERU/+lKaouo
rPZKGa3Q4/ztgck6rcgLGF1EdsQWBid4fGVyPKJJti46w/BaRan00k5pfjXGFqOKuZxOTGQd+UmP
Iaw18GZ4XQzudlc0vOzDTBNFHsjXzxMiGtx2uDmBpLU/wRqbO9YO+lmnVPoFvifLexgJEbOiKsE9
8AFkvRESPD/rYJH79g8xMr+SWCssxJ2XANFwiy3qWXonnUEOT2/+vBCP+hZ+9h+zmvcW3xP8tLdX
UYowJnIcuULE0yuJg9xcC7e4TolKeCq8KiD+fxctn0EWP61749scJZ7aoW3+dAQ+tKaK6h91J9dz
FQjM2la7DHqquDJYMBCeaZ2MuUu0JdzhLo+/xJxuCVPry5+C9Hvy4SF1cNrYT62vuy/uTy+0T+ka
ToRItSjv/pnyeeWji1uf5AhwlLlbbH6XdCXKnyxxyU72wTUN0JHyrLmrUUt7pja24XLRaxKJthcH
MDPCQyF9sldc7F3uYIbmNSnos/i7hMqm2VH3O8s6Lw3LmiQAO5qT2RbKPcu/QH/AFZl+owtvD0tj
9E8EzeQwEb/wvCJ3eGKYT5EUvADqbXyoyZSnKoe3yFcYMWXooQCtX3amgCcIBHXAuwhEGZBxyTpq
DaUi1tlFw3ngtaPpqAjq/AfKeRSbX4Hi6yYQUVtCiDCdNQF4tT84JBKRn+yH/fKwHX+zzTIjgoWI
OZD4MN4yyFlrI75Ak8No4IiMlTHd5dx8SpTBq5UBx0q2ZwrYK5dy0C/PC3ndYRUAmD0TW/wn22i/
BbSxVyMTgGR6wBdYkNp6KpsqhDQxE3xOYEA2UddCQ2sLi8c0rCaCIlEaXs7Dbw20tFnZuih/yIw2
/aFuoA1VKNw5S1wXpH4vFOncKeoIEAUaQTyIgzjDbFAMpSuFysUk4BHFP/Hd44JTCAVHH0nEMNgX
mI4npUhk3CAla13CrIjrFAxMs5xqmvfUsH2Rw4Q21IQpZfMg8eVCB12Cs+PFMU9W0Oiblt4t6BIH
pfl0lIpv6X2yUryZ1/66Ib9jgzSqW3VE6RdElVX5szMWaiPccex/48gMCGXHhQgzojVUp40mGmCI
FKz2r07304nHSDhCdO9mpwInGzXTHOZ6aobkITTaft0Vn7c/yrhxgrTJ4oj2wnSsMrGRSJoAKNA+
YdRa45Uc/UR9tD/WNGD0kYWSh0TMmwKpLKiruqEAWp+NHuyO4cjTmmUUOFhiw1GIeXpYDM7HGjGe
wL97PD2TtCjXCTrp/vLMTpfxGUXRPkvI6BFwkFxracIda7SFUWkrOFr9/evk0AafSoyAc0+oV6vq
m9f/NDgIGnmI8k1RfNKBtDZ5QYTxapdWV6vBp8O1N2QeUMIL+Sx/TNkVx+vS8MaGTgdSYXOSP5oj
DMA00EuAdzGlPv575lMmn5iIZuIh3GzHhRAOwjI58vnxPV23rWHAPShNlR63OkkY3NAQ5+OcDstK
P2O7isN2AGFPCluIPXiFkfBtCM5MxJ0YQn/GSkx1Yn/T/YkSWw/d/mZwMLbElueLkfuGxJXkFVP9
ZPNHLZh1204e5kEQqM+y8NU/ztTDp6/1KuhEEEX0QY1/RPNBHB8qeLYD/U9pwEP5fBSRmh2JCbvg
9LucM7kaGCop8Nby3svs6Ro9vISE9Jx5shcf5Iu6q8u6fuDrUvQmz7twUVrCL8HnTL8YPTWZ8J+X
rfPF4t7hbrFzZHDCFNpJS9JvFUoPznVMPqmfqZjOBv1Jea6zrFe4mWxTUZnyWT97QjZqHdyhgigF
pB9EKt07HygjvJduuElxVH5e4j64m2cln2mvYywjobdKSp1UXMW5/d8v10fFvhbDn9UZTvPc5fsg
rn9AdPIlsGM+7OS6FU7WNcRv/oqu3U0+5dKf3ZySbbXl9MvRhr2xBFTclkrw7w1wR+lCdynVOJdi
sDLnPpnqjXUMdAd2DU8vzjqaw6yFGwd5mRqDwsVDuG/aPCXMGZmjRT3MWC2apnMjS0CcHDXcm8MV
0wN68AY60W0UxBdgtf3ep5qx2OKA4srgOq7FeBj8hChTBRMEgpS5yxR2ehCAlXF8EZZ/skMgQ8hX
onnEuYhM8O59tI297Ardh2Ihs0ObINKobDLhLIDf6duqKwfNmYnEZzsM9EpAnNoZZ4AC9+YfEHqV
nkE0/3p186TmCuxH5dEssEpnDSyZSkVzKqY/ydXUm496wmF936+6mrU+8dlO3dekInfT7Tp46ZPF
EaUb5OobG49bSrpjbNmhw9X4pmZhC+rELnslvEEuVXUxP1NyryvK3ZcKguhS4ysdaMgoc+UjgWdz
vvqqLCt2roSbgOXKkVbxYhCeSV5r8Zb+BlfLHHnR+LRI9+1MJCMo1a6IpXv9NVenLHkQ8kKmTU5X
x4zssAGGEkVj2PR62k/eXZlVMZG45FmCkV/VXnXIRcBLbp83OP9kUcp6kSn41MnV2uE1EvJlrzgU
BtLusc5N4pt7nPKXfWzObEFjDS7HEEZJ2Z99p+zajs0RTOFgfEzzGPZwpr9qnh8uOkchqwepNcss
/TVVI0g/R65mFLHmYb9majpZvmqtlv7WKlPZvZeBLTxsRqCVcJ5+WjICst+TxNQHrqFDp3S6gbtg
0U6o8kMjcQVhQ0EXRBopfCqAZ4F4ebP83X7AAqI5r9rRCYxrLmFht/2Lk4BLkR2Ug68/TgPSnMO3
rQndGfX6CRXj2rs8jVkZt3FqSmi/FTDmeMqD7c3NEAmH27NGCdBRU3DaKCiZ0O+ulQ1634sRCpdf
yforsES3jBO5tB42J2vy44cPXyPnKyA3FSPk/cCmo04Jn1B/2Jjxg9B0IQyj0R3bJLhNZZQZ1lkt
o4Xbg1QRpYwifkn+ZKaGcwuPmxOXqBuHtv2B2q/zRrscCZr4ARu5FPUuPtQ1s1w0veVJADRkmLi+
cjcBZUWC0Z8nQE2RqdRymyiCGQBpkvIiG+CaY6HISAhUXnrUpmcCFlzpqFpXhwejLb3ii9C0P0tG
/sgMGeVDhsDAnA2geDe3PwJ08sFVlp0o/dHbo/cfUbNfrQTZKTRTfI8RvwXgQUOKYNaSA0kg7CQq
1CN4Bb5w42Cghy5pcVAHDV4OASp8ljRRamSR0rbq0GvqDWhgqG+Qv7stM7bkWykpqwwQxLrNSo/y
nPzDJLPQ2jMbA5isLKTb0hYAZXSCT5cqm3S1EpjNYFhwxji9MJremPTHGYptiMnt4lfxc4mOqfi8
dzEwxkZPffOIxUIg2rY4y11i7qQUHGGLWkeJsE+rApIZ4mQkF7cPHKDCJFAnPLLo4SbNebck3qSP
ths/521UEhEWs26XPGbYxYa7X62T/mEyfqdm9Et+md/gTAm0C0JvexQIUvHXoLfWx3eVpkXIwGfc
O4qamkR+pkfJRaZ+w9tu4IBqz1//RIAhvuoNuuE74vw473DL4qIiNYMwj6rAq1sIjq5pOfdXAO74
8BdBS+wLQzB91NGDxl4NCEc1ugr9otD7IbH8EQKKJq28OtvhhYbNtaIh4TPLCi5Bp94uq71Zdg6x
g0QA2J3ydTROMVemS40FShl/yKY4JEKjQk0rdiyYHW8oh/JXRvRmo9p1Z6/H3fICk+QYSIe1cYbS
OqzgJyQhlfLV+Npw9hp74gqPa8+c5VULf6VT+vZKvB4gyCldKKdXZYIeigLAgSEhnQmTqYOoq3nA
o+g0VWQ62W62musTSdUIjaS+J68Nvr1dd5sTYG4K+yK4OeB+PoWcFrgDn6zk/1iQMHxPkW1eEiNR
PxkP2aObnLFhaES0TkuAfG3kF1oLrKTO+K4cN3g1vMU2Ir9gd/FCPKvRJlJSnxjX9kDeZJrgt5Hy
NaHCgNIAepG4l5KtaL9FOv8MQSxRWH0Nf7ARjIs82Pc+yXUAPygoSGlV65TyMegIC+SXkymGss87
ntSSmGvK4tKd0Nx9oZLWHkYnH6ybzrEto37mbXJYWr03sVRLgd8tPI/RyTlfxBG/xCCxI2JKOy0L
CVOoeQtnrsbVV44MlfRJBaBuffdMFERVgLuoeX6MvRgPMTwKYND0PqtwLBdWavvfcsk7B1lk8oOi
05EcMxkwE99dj0UEs/bISRJlTrblFpqkmMtxEntIXvbkRdPO/+90ixb9aYUVusMFZ90Av5KMZpO6
Gv5QtfVPCs65Xt3CiG1ZiBqfShMnd0HbP+BZizcvCc/X53PS1zIHh0bhc5RbTCml1QeFLCcDVsMy
r5JUBBC2W52890PtEoNzqrCbZjwdnnrKpZzH/PWnYmv0sKiYDbfRaQZqhEODyWVrvajADjjONXKF
/68OeX/SXo8oBXEloTcfY5bMgwTyMRQS4UDQg2EaZigq2A7ClFAQl5imk5Mym0nkt/LILEsEkkOt
Jp2sxdvbY9jcvCsnw2Y5+7zv5++qM+mS1MaWUnU1CAHxFVK3WUq5YIRwvLWyCovCEcUE3QKKjQOv
W1V2Vlh1xhZn8OX1Xe7RQbmZwwHwRLpa5vQCt4KWsE0hEW1SIZbrAojQjstu+Dy3OpuB49pXUuTt
seaiZXlHZ1OhiBgsrYv4qkFwh+CE0s1fYUJ1LhFdcNDBn4THI4jPeRSmj2k3DupbnYq1Gjn+jb7D
N9Z9ftssoY1m5pW4wFCTB9wLRjk63ba/6Di3z3jY9EwEnx5TKYwA8RdUEGiPic/zvaU7sjePvcgM
c+/AGucKEXyoMZfn9HKIVHWNV/swlNPFONyOz6LwXrscNclrT80968Nw9yXiPFwgbzopp2lt42tY
Ly+6NjYNYvR+PopC8R+EyAUyG9QFHrVrNXCzVjfhwlQfzTIup+aMIZEvUGsVypERTehp6z6Fny87
Jw22+En0c+T3DKlUN4Je0h2gxwS31H1mjoLDC5t01BXrCkLiPRUzT159BZSmxsWDYUZpFEjMA9oo
6XQYhz9Tid3H5f/Pi0x2bruzR5DrJO9HHTmQYMLLse+KLZfy+lRt3bh5HZZKrFn5DnmCoBYf+33t
GuXJpuUhC16YcEPz+/F4KqmAehJ/y32DsBrNTZ6ATOZQ/pwXB8QmstoipyiCZvoOG5rFcEnrvkn4
HZ/a2GEg1niEewWYkmntz/XXIDgkXaN1HNJcXKS3zCqFQzG6etbR7iNc94A9JTupm6UOz+ILYl5O
xK8vdqysmajNhvGb2axGbsYvGZWQvExtU61LnU3h9cF/whKGhdlNnvFwtcj1BJmGt2shGUqvWGjE
R5MXwXOTRWhvrp30ODKaBu7TFVEr20rooIaX0+FdZvBOC9OvqE4Q/Rys1t8XA16ncrfaCk6EDBGg
tzzRUfxPbk9tliTVlnKQNVsHYzL5h6i5Hz8ZrYap9p30+0ihXQpB+W9Jigovc9iZ0tDa+8OoTVBG
4mG4ZTnUs7SR/A1rx65VRGalm4B4sqkVZDCFd1VKSoz3gTClqk3V3zVKwEZHZ4UswzkYI8KPa1Qk
9brPq8jRL5iYDOPYFybUAQGcLZ+d7zMpaXEXqcoOdjZtx66dtk2SDVnQxV66VYX862QJyX3OkxHS
MTFb+6FKtzCzj4rXSjFYkuPteWQglI9PI/CA5ijDE9lOjkKqHikTnB7asrZxiZH5CVf7fE9/Wm7B
hj2bGRNNB1xoPnrVhntHoCFEq5Rh7E4+tLKsv3oLAvjiSttZEpUjjXuFfdSueOp23vDfDVMah8hj
WriG2gZfyPtSmY7Uz5GZkpTlmoV0cveEKlYSEKAG28nEtF33WpLZX/cwO60EOFj3nAAM88X/mJgG
YMT/oVDzvnGTlMSEKdDYzPCVAF99n6YPrNdf+aEFo3kC/z37xKIBIl1arignnn+ZHTTH0Ov3je6W
Zq29jlbJe8ch0cjfMTOFW9NoW5wo8UQJP1ErXLftXtAWX3dhAD2RtBFtnAXxRKUf14ckfTpvzkNi
gGcAF2MLbtZAVu4HYzHEH3QZmsC2u/UOJK5PiMMq08xt8pAI2/DZ7Knnsf1XxZ+x8eu/GAEsQ+pS
yEK6h7YIWqEGfDWgoSuRljS0V738n2JOxjEPL0ySyE8YmqkuBxmzvdpuvPIR8ud6cCPUJ+OUKk4S
ZBDuRvstOzDqAJsHIrX5+1JMwx3q1sNGq/FWLXkPY9sRKlQY+ugV5vVV84hP0dVTqoRGvuxFNkhS
nWqcCFEr5k4oMbOY9yj9a0FpEasq68QQWr31MzInmtpxe5Ce4pHpANK5X+Gi8shP2nf9BNbwYHrq
pULbZJRUhz2Iy+m2DXWm5J0MHHdaFsL96UjYm/LGxFkRbJw0epIO02Db5e/Mxi1lVoMetMsJM9Ip
2iT2Sp1oGW7wI3DaTdzcI2OlJsEVQAzVna8qu6YpXkqInROeb0QkuHUzW3H8AdP8S8bv/Lnsianf
+85b1CAJQYJO2NdbLPpjQhRV1JCJySzXmuN0bvox1aXS8bummlfBFE45DOGpDavmpE9SM0mqdmt2
0dw9HSn8WF4vqlGROB96uIIENsVytjiogcQBLKclBgCsjXJqNsU6fem9cSPyTmwoX4Ivu1+2L9bV
K3AT1DXkySPgP9actCKN0WhFvBDSL/5xt/REtz9c9doSuLLsluP7UJzq3VmMvkt5/7ug3ZOxaBr/
epM1L8KKo+s3CbJWcHqcCQWIdiCueRKrssgfYkkkRIPwQtg3m5YZO2uJjGSAmRE7TCNEksdlXOsy
Tfucx8CDbiK+4jXzUD5Wl4W6itQtipBt8OIF6dUW+I+RRoLiDDldwV7UnrgUWGOlgRZs4eQbsOrz
SL3Ad65FNU98EB1zPu+q10IL060LwgKHj0vMIgHrTQtcYUGKe6h0o0jPjNZbAiPa6VdHloD4wiBZ
nnYgdJ16Z9+DXIG12fAuphwyd9LeFbP+ee4yEhiJXNJR0eGVjHO6sFkAoDKa/sWeNsuef0OqYhnc
6FF+pYDKp3jPurW2hjPkOCXehKzeYJlVnkdWIDEXsAFlu8PqvytkzOLWtIAP7N73/5fiLUo7K7Pa
+qHQHpoKR3UhgLSCMOjM523B43EkgntYHuZd0jCv9o3dO2HU81j8QF14LK5O1++fV96qRBwszzDn
O4Jm9QrqEhmYgYkHIq4qZvSgLCwpPShmAmZi8dWSM2Lo1xhuB9FN8CaVVZ0zFKoKs7WaGSQflRtS
VMNDxgzyirvkbJpCPxmzeDZ6/OQr7XDLiSu8XclkXJ6kxjHIWst/I/rHCIX/gncdrv56ogQDcMy7
gqIvKh+EOC64TiUHFf2i7i0gKMHy9DvIaDPiDpqRvPeU3OxCMfNU1nA6HIfTuwFyb8dKeOFeXCGX
hmM4sCtkfjsn27N2IeQ9VcyR0hxsPel/poLyfovOAB5v4qDv4wVogKrfRVMT/n/qHS30T+hECWuT
SMiJRabZ7RqV6LJd1t8pg30r/3jOjHicSwkxQk5dh3z1mH+tcg12A84KJ4sN+JC9YAqdhDCB25vz
YdJxMdiEQdEZjh+yvxXSdP1O2W8uXPmXrxA5Dg5AKYnv+07p2eAR4fTT6O2wBPwxocqsO1ptofGP
Lnmy+pww9OexwCTRogCsyHQp36kv7+QTOagDUpGjthyU0kIXwPvBBdFwL3inyD8K9/PjiHwUwpIW
/aLVXD2WsDRhr+8U4ZPXWYLI1Gv+vbTn/7sHpOLo0sFltFPA4BSm4FPbHoWqkz50zOC7xtF7vMAl
fy0aHUCLJcsqzE01ThL8KPH0PeS7xWZfXV7yavlROruJHmBrzi4JvLkRZBmp/eE8LUbPsGRK9PfR
Okxp2180J0ppqS7U9j91jZnx80VZyzcRabAw8xWdhqOuh6SvNSh3ZB1An2cta84sCa41G9D6jxE8
BVObJH7lQefu2NVOH9Nz5V241+OJQwc+1KkIP0qA3RrLn6Oc+71ohS4dcrqiJezfbPL1gqK/Gm6e
2WsAbmcgeyxt9tFk35BzXTwk0c39eU4njl3SLEUN3YNM35XIUrIrKB3xS7JqfC5DJaE5kaXJQvbH
Ld0NfpFW9x5gdr5LAqi1ASvE51hQzEwJiBUcPmIqsRhS104Ls6ZLJS2EX8zMLX7NdAX2uPUd+hjM
G/ALr4Z5Ceo8JmBkm0z0I7sW7z9I01/CPmEvDK0ou/UpKRSt0BKyZjzmROHmJ4MfHtG+wTUMr17z
3tMNVoEDr6OfLyy19u8anIlTWARgXg6r3L+l2VbPw77G5CIfp2744bE4PYlxKdEd3Ulj3zZcEnql
xq0H0h/RDMztwH+myxy/tksnefZvhT++EtdqZsQfB1mc+2abRiELBJm73D7Cb2tu4zghbHwZlpwy
nwQ45Z6hFDhxbc8zC8y6+uKJPACeBTZsMEdOq2BVZW2DZMHLgBZHNaSMxBhdR0y3DivdmA3eK4dD
mckidbsNcMzMulp82IBCRiUSrB8VwTUozZ+J92y4k3arQjE0gqclYG6M2gdfnRcAPQpxdvhL8L2C
p8kmvyql2AgrHNzYvkp49II6UZf2/tRwBGs7SZfio4cUjFPBsKMXUg6qTmC2im+QxJ3asXBH9bYN
lgKMP8vh4CFITVbI5O1FK0ONWC+2xIDqPNsBzdF4Xkw1klEwrvAn8PLNnsRojQok+MGVSFgoAaYe
cM/e1Lh6AffIUswhRCK3i/JRDU4S1C6hvkNKwQ4H8/WQeq5e9W0TYwaPrrw+iP/PL561kUGWAbwN
kXpINgBjASyTgU+e2kG5cMSfRwEReaixheeCqw9Dly80ESgEZMoO+fTWhd9xJE9Xk+CRVxEQ1evJ
ozgU+NlqEywfdUdVC+Fp8vI0j1L0rT2V22XFji2R/vCLESxBJgKAdApned9AB7xzAOwocZjGj5vh
ykCQSCUhwVcwkTJWNjx8+JSO4TujwcU7rafg5KP9gB6Ocj7rTRhUzOzJPEcHxdiIQ++gTNcpNzp2
dXRmaVrsX2M4bMWPWWw+UPih9PrIwpN/Uj8CGaZqWCO6zaO/MSpH1riTC6MrrMRMW8eKZWFHiw5T
c46JyvrGuGEccOoB5GhD1MfWLxBaYm3PRFFBB6hg9d2EYS/NXeviHe8HkqgzKmSLQ3RysvpFUUT2
RcbshRFKYEtnKM0R708lxNjMD3x3IZ/PLcHBp+FldQdMcL9QrKz8n4Ci1IBN7DM4RCXbQLzZVRfZ
lBBAJ822BSjM2Qebxb/FRMZz2Rihv/S+r/OSk3PkitIelgRl+3DRlFiCc0oKtkp4u814gytAoTw1
UJn+nJ91cfXHwRTDiutclkUJ0ILyLnmPU2WHLEvwpos2QyI0zylUbmwQm3ROBWdpX+JwoCzsPdMw
zqjwzXDg9Mpt5/iwhEi19GQ8FtnsXlXwgx6wEfdo+IALC9vVW95UyidiCEIITSPoIHIn+SvIWxtx
ib1MbhagdnmviV2tfdTkbiSonv8NZKmoiArUWMsNX5LwsCAbDlu93ZU0erHlf3pGqV1I74WoyfcJ
MF6XUOvHSJiqTSK2Se3GXIt/kAYs1pYZ0njdf2yMFh17yniHa4Bw0daW7M/U6Ag94facLr+4m+/3
paeC7V4WkPWXa6Gk/n8cD+wZvBiPR/hSufUzTuA2+O4SU8NweO8tANExnZ4WqqGUshC/8E6/BFo1
4zfKWT+9FrRLqDIuCltVj/gyG0meIKj451fynO4CeeuQtN9gq5eImvjsTwyreU/mg5f12gmrQI0Q
tiljjwEgAKzMXpkkudu60krYgS4nKKm2rkxaSJPJUAnzvPp/8UMS5X31vYHIw4dY3dpUGF/ZRVvs
KJ648pxvn2eeTPIyy/J5M60vq2IBgZXia+vJjdezrxgrcadvx0TNaHo3v+3sXK4/DXCzhnZ8PeSs
IW85VPtHEHN3VjdI2Wmrj8xYRRt0HBnKu34Ek9+Sdoyxs+oEYC+8z1Dv9noeCi5ayPsBs4s0vqux
NbmeTvcYxY/0/ABGhClHuNq3JV6neHynkWV6fWc4b7nfPdjcPg+wRFkUMKOv3/gSS5NU4HqVtA1t
sIyn7ptapmaCLM0kuQa4cbtWqJodSAq5EYnxBwptq5sRnYsc8yRp1TRt65oHH/726+4lAQj1iZ39
vDVPQJDTa7Q/23/ajXNEZYQa9W+uZ5Lmk80mjakJ4rXbDanPwYo+fYDOKzWKmHxjymDRhJ8SF/7+
HmHqc1anrIRjmTZUXxP+n0nACMhCLg0BUNAocIJCbuDL/XE9P8aroGXfgoFweAefCYcKmrZoWgLw
oDbL7ipvG7yjTvTeTeC8yG3q6tEoUeig9Fxl78NnBxMX+Gz/18sRmc4SwrLwcckwEVOeTp1QiIVi
eiciJ2I/IRH/KY9Emx48w9gN99mCElNZAkSqPnrPunlfXNRmELruTrq2E9pV5yZMvz2jbNSmWxRv
BmO6UEAu36qDaHqrBZvm8s/10v3vqY7dbPkJSr8gmRp1QeW4e/5yOEeixrEvXUvxzixFdycfhrqC
Hf00kv3A8I6f+87whONcr1j4eupRZpl0RM7p1hSL2JKo3fI0pOxxjQgNjz50uJGW56YNX40RjeY8
vkzGxNolIb9SLWt7TTwvMnAq6n2OX8rstx1orbvIWzhTI/gFHbBWUwQVIXqUnGsWvsE0Lm3tf/NF
wvpC+IKiYUT3ltqyQSQ7H/pLUWZWircARwusYz9FEH472VlxWej4cXrHNItnYtvWEJpLUDk59G25
HwvNR0BT07KXFPLsO1oXvJJWSRvRbSlHjxWQS0ZxyENFEhWxWzgzd+rmeXAtsLI7/Wk4IzDqZ2en
REEpCCFmQ+AQGztdYUsdLb+tdqmmf5JruTbDhLVJPVNkcrJHOr1E3AOQqH3XYyeLkmq+BJeY8G3v
RG749miFgg6fhyjdfC52F1TFR/MQuHiZlW32fvXeBI1+FHcfc6l7d9LYLF/g+z2RT9Rdv0ul0w+k
PkGMQKfMziLgzXIwjohYoeMvI3WqCwx9YzC43PnnrMdjngMAexjumLmN0S+IAQ0oiIQnYYPk8goY
JRsMp+fAvJOhU5SY5xuWl4kzMAWL1rDQuAzmiR6R1CNAGOqL0uw4cdPZkhLh7sdhHC9g/NdKtuAJ
X2NiHQTTE1xpFYF2Cii4dzYQLyOuds/pHtto1Ck2ru3Z3sVRIDrqqLTeLcB7hpKbv3HFr42cgBZg
tXUUSdBuI+Meou1qcycXor1xP8pcjdrTZvlZhVtdxEFYuFP18rGENVV94CTyVG8+qo0iELJtZzmA
2XqessuEPjjsj2Dc7F9NNUM6zw1D/D6FXOqSBo8syx+fBi/93Hm6F6VQSYRmJ5GAaJdeRM5YL63Q
7oSiJIeOnw85ZFXUsEJQ2lkxh3vplyVoEfu8Tra5BlohM4hIUJ1JyeovhLg8Q3HONOpBt3E6QIfN
3T+GOM94t05zphwBQih+3r/BMYsIPqN6qYP2XyUUrL3WQ0FMxvv5AfgGCdJfpFHXyk088R7pzCm8
Nx4S22hL5cyVi3tOlA+OY0/tfeGrCGI055rRfertF5f/p2M9ndIZ3EgBWzTCYJ/PqNFWmewizYcF
eZdvppRc3GbwqGtPxqlUMtlfNzk2C4yKMroOHYERQEfl6vdB7Z+aVlHxCoBLq1s/wgLkxYtnx5K7
haj/hsEDoGV5Ee0uxEauFCC1c0NDiZ4dP1+qzhezPwTqowpPO/0wbKqfVB1FwFz2KhpyYzxuPKGC
0XBxQSXZnOeBF8hHWFmAh06Z14K1g9lYxk3mCWP/ws5e2vSwsilgFW0LwAmGPNguhNreztg7ibQf
qIzdLBrxOJ56qLZO3alDe3WosREEsTX6DwbIgNydyTnEuLq5ODA8Aw95OhOJ7ty3CyQNp/Jqa1g4
MgTX32Zp781++BcR/GeOepjralJZOLqrAk4JRuzqYGwFYIfljB9WuKlAg2iYkAbuFZjeYTXDG284
5NMDdrGsN5CR2fdGISJNRACyAylgiuycQDVfDl2yKf5ZjNvBIEI+KJNFWSY/lh+54qwFwVHLjfIW
VVNClZtDumWs8U82wtDJ04hfvGM71UBZSAT4qFJrV5ZOmvSjr3eUIFWrtQpvT6TDR26mx8xX5Xf/
i3N3aB/WWVnjAOSAcVhFJfHOy75NwlpQ+j2nH9disRC8IFrPHjx7uOcjHVCpVMm6eQkmCq06pjfu
WmjSdKXu6ffsy7cnK0+TJ2CRBgNWjRlKNrtOzCk1XIr8WoUiBzEw8AXGpm68eelH4W5Znm5AWeUi
sZaDCb1KVi8cuDnjcLdtvJvybSBXia8SP9TNt/mRMpVAkR2hookbvPogV3zQ0+/ivUavU+x6L58I
5jMc6qJr1mJzrFYDAGqUM/B5bRF8Pd6RJha1wLwxxuvCgPzFPPVan79duC+nUroh8pwuMTUQhJ3g
95Ta7Ojy1nFfIjGM8dyrDYbrIGVEYyD2mNGpCTyemp1XZqpelz77uY5N795YuMnWpgkleFvPDkPn
BVMsCerAGlryWLkPBm7j6wLmItOHPiDBGuTuprmZY7PbcljNHVSZI47eEOMiZsExADCBGmgPTSkd
BXL10lX7TJ0ZuV+IF8gmS2lBwbsV/MqBp8MVy2OBE/ilba1JgwiJzvemGejNQR6uLrGt0R9nBCpT
SL7QKA8Asu58l5/CLnC88i5aWHytb4B2TUgUn620FLgBFGXjIuQG1fluvMBJB9layuK1XnW8hG+I
5G0FwyJY7z8UGKfxMTUauFPNcmPScExhURErxFD/qFL8JiQzz6SKN3jYhkeTQtk2Z699VI14QxCG
ADmPgHGE/zyMQrjDDjclnDYcqdLeSib6I/BwxOH+uZjCB9tePHVyqZEh71F2Ao9j8Kz5sl6wbDCn
bkWmdACt6kAe96etaADrgCQDiSSTvvNqM7F2ZThIrAVq7rA4K8RA92cvf4FS+SlEeWSzgbYkp6l4
ETtGeOeF4E0iyqh6gRUSnjw+2DZTV8HlARBfOlQZCtu9DGD8Yh5z6+Dt05I+ja77FxDRNnrOAsnH
mlM3DW8PtyPOLyZp2KwN2zaeUKwnzwLSJ6pnATB1OATy/KTL1oLpi2naefDoJsLaXyMesEclpCbg
30LkxVJ3l9WOBSuLDRiGCTJ0gCb4APCXslRUlypMhKqFqPdXSY1x82AnU1DlsuEkO1HIV2oO6tXv
6+lg2B0/prCCYV/dMcxobkb94XFGmbTspJVUI0sBv4TCMZ6OwWYOoICP373XQZ1dmnpG0vWdzHXM
ROiIbBu85sSQNSNfdUKm/DQbXbDwAtJAiO7wssmmHQSs32F1wf3TLEiOAPYUVgRCH47UXmIJcG4V
VQQLVh+NfLMCHf0Ck6Ks2xhdzsIkYgzwwcSAnEcp/jdZS2rOgs7E5/QWivMSphus42CEbFHk3678
ERjfMRbj9nAHS12qZJ8EOeTsIA0P71ctdNCTKHBDJaorSpTTrsAVlredQfoBIpRwbaZLc+RMgnqI
vtYVlF6vrgzRdbpeTeQUJ/WnRdEpg79HHRUO1aaNhm12shb8UaXWrdrNzAKj7TuEF0ncS4fNjFps
UUkYGBRfjj0WfxpQa4VXyJNnzipol4Amc5y52eYgSl8svoyG2smsKh8mfByiH910W0H/SMsdqpHr
/duPX8XrEZHvlf2rtDNH9b+HI4tkOcf09/p/J8TyGAidHCdaz0pGTgljdvSoQ9/5fFf5EZhOrlqX
Y/MHqcbq1m/BczOcCYnunnEYdkxlluA8veY1S/6cYWAaEJAgK4H1arw/jx+PM3edTrBmjdKSkBxx
yMvP5vPHs+YnDB5cYgbS1zyLyTyYKbDB25X87YSvEwqUTxstp2+Lv3zPp0L23XEK22y03nQt0r4r
1Sjz6Dn1IqZeoRZK+zPZKGkz9vVMh5qKYwJehKpk7rF2PENIGM9K0gMY5o0JIaywpxTB1T98WyLE
WcNnqtnCfVaAoX5hFdTI6zaY1aRX2ZtPEsvhNz6xGWrQQXSgrv75sjZYkVCEUFPGP0YD4A2Awbwm
cPejj0Ko+oOSSKAYv0HGNwV23+gQeaOPZGRXr2Dk7AevSxs6WWMc6UPa5Gpj3TxtdyqBI+EBZcOX
Df2TJD67NZFYVmsFqYnQAl0AwGqUTaHmCLGnLi009Vhfybtp80SNQzCiIdsSKXKYYnqXLfAb3VIl
yV2FNeL6JZVY2V+wDD6/riNf1ha65cjZn9/lYYVC4OWaG3MdQLldvmQEbgTNj/q6x1ltRu2BHKoT
Tc0RsgKk3LvDpBNVcsQx4G3uGDGm/j16rK5F/tcD5LR3JJqicmq49C0iw40NjM9qXxl9rEdLlDws
NhDwMTiwhUUhddWF6qTZGpY5BJP83EnEXgiwJtGgCchMTV147LFYKu3vN3COYqEnPW5z7tC01YMp
uUypDTRoUmbVqNiH729tYVFjGTSxX3Eo7/cnVXmtQpo0qhgmSXKKSZBFQqF3etSGOZGJiQbOD3g7
5j7Ch3UjQTOM9NDdgJ38R98dZifSUzhCAjC0V/0yaZie0Nk5U4BRHgfen9BSuWzAHYD+DiVPpZiV
0onYZqf7x1rLfhuYOjxAGWy63TGQoyorS0i/hrl4/WfBvhsjOVGy+NTcg1ggBL2D2Qg5f/Y/3rPN
jbXYJGAmkmOX/CC+S04X3oVxRwsqFl1cHLZH3i7E9Dlg4Q0OvhKSGEk1JBpjAXK0usT6vwvEJtNg
odOn7bmJ4pi5FCwcZbeC+pnY6w1oN56z0171s+ZHFTpr+NVAtsN0GvO0l0mag4Gu+Udto4khCHxr
I62K+BReyx35E0C8hPzHG+O+j8Ts19gqQ5fkoFqgZpxyhajuB2m44uyEmCG0V8dd0GjBehbDm/f8
bgo+6e2IYPUxUS99suU8h2iYe87iwmE6zwsnfiWdlgX30k8bAXf3bwn3CKMTfnbkZ7IYo5G0qh94
hGxgUVyyEzqgmVhHToELS3MXsa7Ta9vL5pZxaa+gtAqp6CfTaURR55hbzFHyaSl4gG9pzx1/As5w
zi+XcDe7N4MVQaGj01IRHkQTX1amKLcBtU+rVz8k5Y9fIWJwXH3lOmKHaAtPePJpfztBOsIG2hdR
c+VNTBUpjFdgwEvMhYX6/9/cWRY8/eL6dNgfhNJe7sZHK89H+qHVbnWNPQx5bxG2k5Mcse0CzTFE
9F25lYlGFOgi0ipPmKRKkwAqLEzBv1BjRkiGeDQvG0mKFWxxtEhyhonAFHa/5OoRx94kCOOlNnkv
BtkkhLMNQny9zMC+aRsLYnBZYRExYRhmqDwMEpY8Y8e+nAxIJCk6Nx8jt0XF32kjdPh5fQvdLYiL
Uq5+T3qSePDxsEAoC1zuScNFZbVkzMqTW/tI/J3ceDkPzLyN6GMn9JrU0Ke+QbWb6n1leq5pV/SH
5vHdpVrr3TiV0BZ8LbLsBCa3vQfKzMn9Td9P0w4YBpxQlAJF3DfvndnbwRuPW61+Nup0VIyb0uyK
iXKd1sI1zO9LRmY9hbikBBM8dIFEz/1TOZIAeWZaYnXrSdz6cgzapFjlkdBV/PYzsz+4nNqPRckm
Bn7KQJm1BssWnFf4e1iqTP9aajdy5ZAqyIcEJxnuYODn0pjCy+UsDXLunN0p6VPP3sbUARNi7YFq
UdNEXHKnmVpwjJ5t4h7cjeEJzx1PYNLG/U4es40l+MbltIhzhYFU4NX41F1c/beUl25j7gXHqZMU
zdB+lRZSh4b1WpBSGwCTS7nzXdHqU7AGD1kN5XI0DNE71I0k6WApFc4wSCEgvdmPFWf/s4tvuOx5
elIRQ8xj+cL4AR+VdVVHbgNj8ppFvfSdaMxFJkR8Rusy9h0i/+7JmG1GRQAW7Vh2mF6j75KjCbxW
HhHrbxOMcZKLIEV1m2Sjx3CxTbDQ0/idlrvX7Q9u2uUkDLuVEE+FyKRvo4KwbvBkReDLLLFutY0K
AoLmDWGJjgrVSNULt8Ck/D/fHpe5pYZgy9OT2OWd6wp/UzwfXfHa0OK8CPUoOHKGS+z/GB3+dx52
WGcAjnoOs5qfIQhnIQVrOBP9BOAcTuTaVYkv1SyK61ekUl60KCjksFm3Pm7hrm9Wn8mLsJjD0WTy
2kkioFeW6/qQQFhwHrD5RZVEY263iwmJU1nXv2qQ9hw1H+NU+rfs4Ozk31Y6sWdFWb1uzV/RavPj
nxBYBxW5d0O1B0bnGZtzHkcq2P0FWTQO0zntufsq9coGcbCH8pWr+IhgC5GxJ4kUb/xMmEP+FFIl
SDFgVJGfBEju4CXZdoQa+NP4upgKjziwrDCFpLredgthdG0c4xWG2cu2WdHszruLZTZIFiajLVZp
Atf4l6Kjl56LSBpfCiNpSL6ZewCQUuLo5f6MtfK6Klwo8GGdukOyF2fkW+/vhtweUokBceuDII4h
LftAdLUzgxbyD6qAyL7ldlLeVuo+CpjR7AcTb3KBzaFX5AHGa6o0ZDEzgt7MKV1ipoL+6Lx2ikNJ
2nrjDizMh4Ge/A2cNNk4aDFKvuOiO9cojbxAYMmw9a6vDBqeOrI92TpJvqVf/3B/qkBUbXRVJodZ
fQkS0OlPC/xilDEZQjGIayYzw9nyBy0dxD5zggBg9x/z04uy6TjLpedgFTmZbJWIuWgq08lVTrRy
bwBso0F6gNPQYDzG+2Waud3LIuRAemrjmIkfG3GWgpFsCr6fsJzmlhRSZruvv4VmUXJ2RMn/VPiC
hzH5gItuIDA4WX3EYYONb6On1jdRvGdkd5iPHvo2DrvLX46BdEmdpAOWVkK2WuNx3RJpISXn3Caj
zA0iUstS6eSdR61XQ6Z+goTLHLV3ixO0Q6NmSGsGBLfar93uABIJDykUkdqY+Uci2tSda1Zt3vUA
np0ipIO/lJ7YgkklkDGWB4SaaKIPcVL5+TKgewGsjGZOQo78IqollcaWXy2N9v/CakjegeAp3QGu
lmm0EM6oPrr1ayMD2X7Y/k8/VOM73W7V815L8s2d+nUVP9qvFmI0MOo2L8oJmd0dOVASZnR2ssw4
in3QyDI9xU5hlTgOZ+xfzKhVfHILigRHZG5YkMSTe9533vMQ22HvDot1G3xFZCzek+Z2B2upcheX
GtMwwgozfvskNnWnEnDYK7DvvihUrqYPLDhWWLGS16FiT0vORZZWaJzgmmkgopliDpp+ihzpidnU
XddPiMM2wzw51BnhBfX2qAZghD4xhTeQ75sdUKNhuyyqqrm2RRNt82+plXtW5qa5zV0hpjqvn6Gm
zCtxZC1LkE/YHqhW1nYsJXrGp4WfLOMHBFlv2DQuiFzb+dwgh/daR01ipkhZ2lgJjS9nSz0yR9JX
fEO4MMNrEEvrx177l+lEj7Z5PFMglxd3sAVIgcncrM7xWKozE0/FvWZPIo1g6kCmVJ9ewXZ+Gqiv
4A9rXtaz3MYLAFHyANDgHbezFb1UfG9nhXDQ8ZxlPC+xCL3jrn2E7E37ThWVCwFQNzJnwhDklApl
DnEO8Bf4VLylQP2PP7FQx9uDeKpjUNZpQKhwGTKZlEzK1aA2elFj6zjIkUld9OV7T9ywtRRMCutJ
r7wPmbGU/uiPNtgA9KlAXZdWAf9KyDVTmTWlfC6gaB1NHtjoPqLw/1z/Ky3pWa9IK+Nd7i/lTlii
6rkwWOnVlS5B35q/ftVJIAi+19JcMOpF9UrjYrx1Rt/wo7rsrF5WILpJNRdAeMKYpPrBX40NDNbG
WQoTJs6Kj2Z76I5LkXtW4AP5/U+7T26OH++CIEYUbY6fMcD9JlDwh3J1vUAWuBUgsqM5wIVoILTb
4Row9f60N8+QxE8aaFPFj5S2tyQWW47N68V0P+C3ZeBAZVN2oYI5p/e31puqTPN/4QjfIyIMTXJw
Y0DyGD29aJTUaqg8lG/jqemKJ0dzsdIh54U1JfdLC4heT/LLnTVufzp3uyT71wku+ONRFUK6uHk4
vNxrLj1hlLa6b9K0aLFzvt7W+1kvxfeYCXtdotYqDOuMPbBit+JaeVbhHL7ubRYSd7ANHKmJ05r3
80a7q2PK1dq2OLA58RQ5vAgeD5OzyjNKaK7TxlV7aXbVYx7mkAAayFCO9roMj82Wlog/suuZ4zhY
RHZaxlPnqzTJSAvjDKPMLtLjosUVi/DBBktIQ3Kfcn/TK4BsyfvFiAS9X9rOi2xsTFxY1n97XRjK
Owm1r1tclvuctn8D7DDhwJDYmWSs7yBUdEI/uEEatm2gqKusZ2BHDqcrZytSpBkq1b2eKJCbfpPS
P3K+6a34VCPnQmAz3XAgN1C0feHi2qvLCXpeX1UKdAbPoTWzzT1JOzpAmw1ewTJTdr/h1vbQ/Brt
pHpf7hyFZRxBVXK2za0w6mhsu9ei+bVNM4vTL8fLr0mAkL5SCV6ASznH3/FkX2PjOIryQ0r2bRvN
Ctf7ZZsVCYG9ISb3KSIpz5x1GmMF/OZuA2f/wrLn820Nkr4P+q9obxTTAksyEg6YJkVQN9xqSLE6
8Ws43+3Cm2UMZIZHHpNG/cGYWvFvpcy2MD0rfoJEF+bDSnAqzH+6GIqugLYB+rBLfyBnCjcRn1ai
OROqvctN/wLjrmclG2Yka1rk/skJyRz3+w0cG9kH5JKP+7h4EyYiuKulWo7QWNLUfrUNqhDsv70i
7BCQgAOKGFnN6qlRcp9ms8RRt90JaEvxRpl4nPASuPbPvjnuyGs229+3VtyrGBRKF+LjlzLixZXP
lxG8fuX1SlNidY3Pr50XiBYf6yN0UTK/IVOVbJVmuuztUNAVOKuxHp0UyyYAeyGvVulHeUpC0+LF
dp/Pht0VpExv0rhm3CQYs/yEE0dy9NELuVrKgutDaMhHTtFLhpL4QZAy8KAds5mxl28BQBOeuV17
hawg/Pv7UGDayVKM8iKSn0fro25Vjq+5xv40xwWTopXMuUlAQkjiATrWXmNTx5e2fTENThgSTp86
jZfJiATT10UJ1BmINWQ7AbturHGUzti7oPanDyk7BJFnLuLYm35yGB4ONuacjdzmwKn9/1Z/CrCe
vpIYybazQ44dpUOz7Oa8fgxVMmYCIEGK6PRoVVrJWUtexBD7T2soUOWqoOWF8gL77ADXQnu9bwx7
vz2r498s+wlCxGI0cu4FMMnScQDgKU7O94uAcQrLLdQMKpFsd5LwmCITOgHSpZxV9ZlSWM6EH2u/
dlk/jbBeC3kx4UeMNTh9nbQ4YntQNVhwqXGsB3Tn2JAO9B3hyZi3QscZldkpPg4LnMHc91MA0k3c
4Ru/ise23r2xEz55Q9eVf5PhtAiOTYKwh8CNh9iUIlGAzg2jKs4eTK3VBdFRTqC2cxpZMVdBZ6yw
RrsdNYukvAj1QSXE7QgZ2AG4eKfmtviNUFCbTf+OcIFA8hPUOswZ4A7rNt68qvApU7qnbi68L5aM
tbMNpxO9ywDz+aZmXTkJj1LH3tTd6WbJpUyMKeveFIYPipprajq5MbNb1Gji9T9twCWv1dGipZQe
eOlZ0eyI3OOzmBtXIe/vHV7trvTc511TtiP1CaehqV3UzKMhWof/134qNvdTTbqQEABvbvQAYLjU
klAYKhKjktNjJ6JHBdBR01SYkNJhTYYPnb3Gi9r4AxejFLsIE/Fups2HhoFiSUTa2eI7m4Xrsc6w
N/s2leU6doVJzdp8AzHNF9at++omz80rV7XNqxBwdBwwPTJgTrv6ouQwi3isEo7vr4349p9kV4xc
qkkpULuh6qKt9RXtJx09KxvXKzhQxhrw8jR7AU2LqKRRz903BH99WBPS0LVFysswC9K/dAwUz/gL
+GbJRKPXOiLSv/s8HmNlNgrVxydHZC02COq3qmvkIC7ojYsaP7TgcW37uzZbPDFQZx/Sq9kWdUM+
f3pz0Fnz/xD5mbI5ULch+zU0gWhyQ4jDIBPv2BAgWxzfZwwIur33FUWZRbgJAk6UYefJ1wC25Sx5
zXS1/zhbNYsv/5kDvT2JpqB8ZXQsvaxe/ziaUYaap6V9tUqn1gN0URqDrvSP478l8DzE6kn4DtT3
uJxUusptI8Ff5gUY8AemthY5R4I3I11uoBiFQIRYEpx0uH9qpiuIj3hsxfYNX3oQgyAF44hgmvzL
TJOWivFkmebcsTzfAiEmRGPbUmzW9YXfS2Z8F2kTrB2VRBp8v7W1kR6PzmM+3rsTqI31Zlf/t5bf
DR9RhYcFi+M9iSRjxXFfhplzEHiMyOEdO3jCXD6sdH/pRcSh56pn/EgIMI8C/n5fN5oq9C0eHKEZ
M2x/Ti598K9zOLPHxtOXrrjYUC0SmIYat4GKXIepX+SPindcrlin7/BCZYNijJnPka1AS9yEjs9m
sOU+C9dOtxdCiVNSnjzAqwk4DvEN3MWOgQyzotTXf8CB/KbPP2/gnmcNCp6BjwXBmm77erfUYhwT
oikjFIyhWxI9LEMk1wSrgJjgoyssUbE9oX+ovZJnUFHXrULojGdSASQSNK6MJLamaUrPDIPeGJvN
qDt0FcS93THG0C2U5towaDaypZnCMrF29JZ0ce3jJiwWh/MvQ0r07dVMX6l5+JhFqnvd8o6y/ejv
REcB02LZSE+uppzTEn7wi/j8lpWwfZIzdgILjeCOa6Fk5I5IR6AfJtninVzAROKrXAOQB/J8dGEY
WvTG7esH2kI0ErlGs0y3tcWxmCxbkX0bNyc69vaeTHbzQW3JTevguqkjcMrZS4wmVkkx8SOnWkTs
mCTU54g54a+US9UAMUSlF1eR+y8wA/Mm3SBQzPhHFRCOASfeeEuu4M356jx7B/QIoEN8k0u8ccXb
PASiyqzrX2KBNkdcPNJGv+pW70w7JpFSfKRGimojcZQfi84bKXKK5pAX1BcNmbXJRZsftC8lLxIG
O7oK1j+oInHwoW/SOuUydFc2sg/mYaVDx59V/UIvY1zKndnybjDJ9G8xN5aZ6eepZ/hNlK2bqtt/
21bs9DIOKdHYzipM9ObLS+O/+fsO4Xziuwy/0/AauY7Lsq3kIvTjcC9Mi5q2ELLEIAxBoLRnXFgK
S/24xlR5ObjehKZQZ5cYF/C2reBm/j/q0o3dsrPhbsAe81DLp04qwM6t7iA25J5vfc+M7h67oylA
wpWXixjAbanIGjZsSoVZZzyEHxD1JC1oWzcdQfNB8OuUdtUiZvl8tjoCOvait2K9RESaEgN32c2l
arMIdofRlrvVjsiCrUEqMisvv+qAHe88Z6DFY7ccMOuXReJIdbiJ9L0TQ1yMbbfwgmorzcx7Tujd
CwLtXh2SFsqGzFJemJTuT1kfzDYsS/UxP2tfarsMNkomKPYwA2Zuo/AdwpIl6rhKUwojTKk7zJM0
jFw+8SygvqjDpOrM+rGNyl606KlxvZd51+MicZaxR6+rEsjSoVLM5cp/z2LPfZuy9ltCi+7XZ9Za
nNl8eD/UCMnLrdSGzl+mRMyPodQ2IFOC3pO9eMJYZLC5wjSi/Eeul3TWnxdWtsUt1JPsVX0IcCOU
smvbRRmx5moldGYE0kSs/L6Rs58lJWAB0JFh3PGE+O6XQ42v8QfGHehkfQZH7EgCCAmfxwGsKaKs
n04+UaPd6aYp58+V9/CJgeTmasfLX9Bf8FmlDz7SiAVfd1eHWgxRvvNYyzA2VUU0dDjpJ5ZEEY3o
K7BkU0h+E6O7S3Y4meH61CRJ3eP+0I0rFF90aNPO70UbiikDGqUKL9I9c/vUOzfmLBKyMoJ1CCqd
PhAOSM16Dx0fOHCyZxH7DjrpR9X+ry5zF+8F4MkD29aAjEU1XElCnlQVxIAVHPbLwyVwWg7QNHOB
YModQhgf6x/ko9Om+v6rqf5X+QM8LcC559W7qEXzdOVvMjxN81a/dUO1/LtPxfErzMoKfxOReKRJ
VDsso7b/92Orq8j3W5LJJYwbH8M8RRHlK6aLDBCFNRFeNqN9qqnLU0I5i5KtMtRmKGM6zS65pOU1
IJmC3fouZrBcZgK+J3/lumETVav3SRzm97QXzao2G9TN1if6oa5VifEGl2JAZ+5w068Fid9+uYHx
mOe5cM4FDkSOFHMrPwJaiMmo1U3yLlFf/gRWt+4jS7sJt2f3UPez7kwHEU/+o3yUMqQ9UN7BF6Vm
ue9aXouDy1JC53Mp72tsVWggU67JlPFiowQcf/dBYtM5ci4rxf9fRFRqkG2/YZZziLT2FvgR2/dR
D7hZhweSGpuf4djKR3NyNuMaYCTWKPegoQiGLrve5mDoqzKHUWcLE94jmRoCEl0L15z1v2k6WWVf
jlTfALc5Oj/zd0fg46VIjQrz8rfPT561FUHvjNlKKCJvXFsB9pI8i5hYJC7ex8DmnCBqbqL1eo1U
K0JWS25vM40tr1IGgtRuP1rzel6yrinF+hWlCZsgqLlmfiD7PA+ia1wRxpYRCeYpWOV4OTb9TfL/
MRvu9XuEgDCnE9nqRqqqkrpQdN3244o9z0wXCQbRowPfeu2akWVwWbGBTv0aJbHHDy2QmRnxTG9/
p3AezROkeagIavCG8cXZ+raIOee6cz/wYggmxGSYdOoSkAn+s2nOFfDHqGv8fobfBmZ9HQh9hSS1
G+y687Bc4E+0JlROoaZZmpx/ytqF3n+Sc0Udmv94qP8kxl0iMdyj/z+zRyFxOumbMOFGRAmo46BP
5TMih4DOiCgxOihPJOUT2GAa85ojackHv/8USJyh8ryYC7CiItv86gv2Tu2jom123rhe07L05IIs
ttWvFBoAN5OAoT1px7NIATBHCt57sSJ3rCt3oTbyz16CHwpy1y3C4UljfkauHFXL3HD+fmxgJJO7
W+AUJNEsEdhXwU1Qlbb66xOiKgIrxbZqh1JqvI8QVEcLzgyZMWZ+5OE4FfRs+8s3Qs+QcyDdn3YR
u68l7zK7bMqJ7bD5m3hUQ9Cgn5aHJmbHxB6uNEabOmbCG8+bXaBzMvwaXxhauWyQIIhfF18ffMTe
gtQLo7oKgiWIAKkKY1ZNgAvmbQisT9uZKMdYr0eehxJN3/M1PmKyiJ42If+gtnhyl6HatVjFJpbY
9FCl28r4KQzu7N5A3Z6uWsk+a5s9U8q9QusenopCgd+2F9+KZWynN2j1Jur2A1Y/zzaqv91c31AD
ErBPfGdM73uksmzq5ReI0MYR72QGiuON1dUzXsAehXaw3KQL8ScyzfpDevZi9Bs6yTkU4H3ZgUxF
F80O3eyYVCXwbBaQupimkYxtdRMQLdPQSayQpTChUBOjpx4fkqfPGpV2lL0Lx32ewUNIkUkQEItJ
J07Uhs5KeJNJCaiCWWHmgZNgL4ME3BTd9FGD+VggypYPDFgiSCbIK4H3afmiM06o3Jq/wq48XU/w
BD71llYnpZ6vbm1vhFsFb6VMaaz85JZQEXHRm2Rhjpk2tH+iFFXDeBG31rmMQksvx0jNpqOWlPtY
SRcUWQB1u1tUG7q+Aw6tkSbv4hmx2iqRyv9tfVXt2K6JPCRvWdDo/Dq2ntMIlaeA0oRhMjL/NX0h
oNnLn0VXF3UFr7RHxzyEXXLaNa02lIflXJYL3b11/oaHkD6Xf5vtH1k1/IraxLKjMpqD8PXFNSFk
bGRwKapXB9LMphRdORO4aUZoKk5D3UNL7vt1maO/GhjufWFFs683PAQgKgtLJa/rPNtNpsMw3tK5
lqpzzoXiLQ2Gd/ju36ICBA7UKzBr3WrizYUPyY5G4fzoB5OzOo17r6mVeTF96LHuU+awEWZNQR8h
1x+1HoINNYxK6nH7jmWvqAlyHyZ6U0g7QoiRLDYoJur80zLZBOnvGf0hcntzqkd30G4g//jemDe7
tb42jaG4uq1ieJBYJk4/mkvrru41lz8WoETmkscVDux9RGCAs1jiX6ae4ou4sciy9J4J/vJNGWL5
84m6w5MkAm2HBnLTyox5fEZSAqjwmUoxmgaS+D/xIJwz/tcyQE3r6SbvM/yCp0RNojyNZJ3m9LIJ
OUn6Pzr1XPZkT4yAPFUWkJGXVpisJUTMjj3q8zkrbKuMXfMivweHF6cc5lC8wqHa/TYQdVRPa/ql
uBpPdyl1zui1U5ObJQXdIL2ZMeMZvnuUnI/khICwkNi6JxnxlSdGb2JlRFPT0mv7zmnWgC13TH+g
kMt1TxJLKaQ0OQVKwNVicdSZ0E3PowsAQYE6L1O86k7tEmoZ/pvlavOY36LL8GC5TzYN7Uq95r1P
nmLSyn/8YhgJxXhMJ32sMyYfKi3zo+zEisruAQ31vUu1r0iSA5RWh3yH6p3a6ZNUxbTSza8KPPWI
Ykdaji3e+8HShjElHyMNPN4lC8lQylU+yn4RbJ2XsnVv7o6vfvgjar3fcRdfnPs6Ou+jtMeCt9Av
lgraw1tdua7ztbYalmpCH3cd97verUtetnLxews1JJOsMQNVkNawaSXatD1gKu4Sjt+8CM+Qvgwp
P+cXZGDjlbbazTwfCnLs2qK8+S7fms/EIldy6UpIVm2PXu6ZYWoaQmnMkjrGWNm7VnJz9U0Klw/U
RSCh70toQvEA9Gwhab62WjT/GuZMZMNv8tYT2Xay/i3FfwrXGIkdAuWvZpS3toKinfJmi0caVJUs
mnri9ac1+c4HpkNd6PfoTnpn78Mx3XH23dZXWyD8tVpLSQHw4GJc5YVrGmoDG88D+zP2zlyz0DHp
HiGoe5OCbCTCwLWuwVN9O6WkJsfqwApV70CORj6Y499WnmzexRO02cPz1HsgOqldHmc7ZNuIBDww
hdbxOE1jp+28m6q6Du/I1ZUrjbzColFv9HdvaMZjqvBmgSSQcRDWXhZ05fupfkEb/Ndk2IyGJkUp
reqhELe6t8B1CKjHzxUHW39XEE87o7t62XDGzNCcr8vUJ7ghWTQTmtYai6qzZb3OoqbEE93eA1fY
eiMLIa591aEMyEB/yXEg+Ma5Z2H5jl4skPAWpWK7i8Im1klmP7OIcfYlUUwr8mdnGsvhKOKer8UL
qxAAAldel4XMmsFlPbRwLJmUEv0jbFk4fYtWIK7cw28J0ED7hZ1toR1BxDRxs7FgSjgHFXpLracc
LJWrFqwzBb2a29Ta8VvtSETg6OMhWLxGoeYLYVXUyJusPPoWBj+edwXNKEqojetStnX9IIKb8lZ5
/gGaih7TyJfZccC3PBXMqW0Jxr9OfU25Yrsshjcrg2lAlg1yYHp2jX9MVOzwzWb3vDoZJjIOqb7/
GsOm0h2HBxaCEneisBgGeDYseJWtW4NotSrR78MOFMbgd12qlTMj4S03m79Xgxsy8hMkEu2Gxzoc
4GYGH9bpHHX/TRQjcgb+7+LLfZ+7HkHV3ykE0Uuj5XUtH4Dcq5UP/uyY3je2ckLeT5Qvlk+7ZjBS
FidcRI4+FE3wXVovHS0pLKU6vkF8V36z5FDYYjM/qow3s0sc/HnTFD04aE0NP66VFx/p8tpc45F1
KQg/OJ59ZW3Tp9Dv1X1uazwbshnWF/InwcXdbXgYeK8IoEcnueOpIQYmzlcFq83UzqByck00h1yi
GL+0wEAbS57qfAw1VohOTC1u1bNMJdq5Udrn8qrzGCvK/rK0EhcfKAb9UtnP5zZUqPZlfD3ZkdXg
VcdZo9ZdsmsLTzbI8ErI54+hD/aGGPcgjCF1krznpZnkrQFbK/9TlMu7dwr9pSbCTkVBPV+2yOmP
U2Z/4Q8tSE1KZGk0if+KgCXk6MeX4nQDzvFP8dl/yruS9OPwgq2BOw6dcPpKJfPX5XeEBe5pYpcF
Nede2mae5jiclevIwDWxDkw/0RFeRw/czpaPP/w6Zs/Kuj4VdXGjRNeCaAYLR7BzYS6LLfTJ+XUa
uW8KB0ExzWYa4mtTqY3PGMzae1OAquWjIBcJVhQ00ED07v4v4thrbCZ6wYAUJyoih1ORMqmgXLww
JkP6/Xh8bDt21KWjG0mCcuqnL2zn7pX0vetWGOuRLwCSTgMHuCO4jFsqV3Nvn8YndOZBhI3Ea7kl
m/jyUpszZgdfVWVm+7ZVOVPc+Ex7zcfNWdpPbf5OSDAFVhioq4EBTeKm/MTnjP3sinOkA4/LFAUI
63n+8GDpRULNa9mR6MCM23zETpD1IfVojE0z8Gupfiex3C98z8xPBFR98npZNwQEXB7WnYWdN3bs
4ESTsageeIPRSYUWQIzTJsChXFdm8/wS4keU8i4V1Mljc7ZKZwbYuUwJ8n6Is9i5R6oQy43QG1bb
6oUUzn4MJ1DcKpxIh2XmCPOzCZ2sqb8SZufBwZEvuX5Zirtc8Q20GWsI8BFr6BsP3maBl+CobLgT
C4TsIUSAAUpnEmI3mQY/2unP5gM2szvV1ru6k/OCebJcwl/1wiPdByW1XS3D3iHbRNnRjov6tppu
E7RMnrCUeuNtoZepIf2IXDMmLUdr5dv7FSmwkpQjFSJP69BnvAq9+V4oS2EfyHOkqnrEJEDZBn1M
vGA9Z/zeSPeTsbjxhz7YX/9VMJ3loTXJbY0LH7q5zGLKcfmX03txoORTEFoE99tbEWgrdXrNpDRp
Ne7PPcsM/qwg/AVCDA9j/Rvphv7zGt7i9bC+kS080JWei5a1bQ5opKk4N6LE3hgh6jtPFEWEECyv
d73UzVNkH1D0cKuMj0ncuC1zAOPAEI92uaNABkiZNzXtSwpYZUYWPVskj3ua8ly2E5tb7yyvr5TJ
IhVQhbXPS1PsG/ewuMM1gqbX2UqOUm/UNA2Qnp4s9vO4ka4GHGHgHEMh5G61SiNY6hEddGGCIprJ
9h7P3xUXTlM0emstjC1KippJXdRPDyiiqOUFeeu/D4sGTwOV+Ow2kVxvtaLePQzo5I+EQsGkqCwL
DWC7NE368KoixYjjj61Ur1vycFXeF33JTOpRseI2MKQtv1QO+jWnoj2HqtvXBueo7RQVmfW1msxM
OEk7U8qc2vv5ORdGE9+fs6ufdVvsOL8eEIr2oIvqZPiiZgxAsewGd2APxQqXTAIRmPFLRv2G+Vy/
lVmKgRFeyI533HNbddyNKJpJUpD8fn4bBWkd/91OqSoP/cO/G3HrRXnTKuHb4n0PvQd2bTEnlEV6
Mf5TKX9mEX6k661y61DcEz1YcmnTdCE/cmea+a29qG4FJVnDkivC3wWuxU/3xja3+1OyYyDp6loi
xkjkvfsCE+ylW86/KoO8SL1fR+p+CKOAKWgPyYJVclJYBJuZBllBOMePmdYbDy+x+HBU+Lo5R+VC
3jSupuRdIXz0FBOmLdMD4koL5mQDAIa2Jtb0Er3z6q0vJgfzYAC9qqgCmVgMnswcMf9HinOrAvZd
WQCdXcgiWCWit8E295j9a/3Osi+4nFoG1d2BfAoaVD1vzkYEAbwP5USYKE+pVOiGllF8qLKOvVz6
GCW3OB6m0jwIYxmtXmub/pBpYj5wEcWx+H8/BcAFqreCzNOPVAhkc7qGMEpjVEW8p9w5BsRrRm4F
UYesPHaXcDZwLQ5zYjCHp3sa7OjHrWwuKnlm4E7u3fdqSH25ktiYh5on4tLeykaqUylixHSbu60g
Q1A44ut7F7WwPTMGJG9UbQhVKe7pGsU/M05pV+EOknkVUuBELyVWXIXy0hWwjgObZVqrTRS8PjSe
gbwpiLyH2Rabkh1yJZFHAjBoMmsrHQ7HkxfB6fbhsRafcecUnlC+M0yVPro/I0+ra25Fc2etx/Qz
J4LEXe3HXQyHCySHJTtkTlJmTO3A8kVSgUTlnNKR1BFokY66y19iH4VFKutbHNFVddGVvVatgNh2
1uexCb5fSzpUf+QOAQKLAoG28U0IjdhsHzlYuKSrrx5rCpt6GZLh/moFniJR/BIpNo1WZ0nM4bJO
ft65jvWNgBaWpdv2CWR36UixTzws3RmnzIrBlJJ5Q4Si5pzHnAM2lE1ltBnsnGcac2YxoHcfwn04
ylHA7b3yrJ3LA1QxbB9wIBxSVXQTIKezjldb9b9pFIMPTYRm+wvJ3ghLMMANh5vT4OqFEdHJZLOl
1hZ2Jm2FvWMAjA3myxv5H8qN4V9W9hTvxQX60P42MyP/WIsluu/X12g69cAri/93lZuKn4IDFfuO
IBFx23b3znMazM7r3Tu6aLiZ3TaA++lX6jq4INGrtGLlFcLjbE0gKRofA/1a7c+vxfh/C+ZYYem8
76FI6pccogCjHfdUDE4oh7uCAE6ezeijWBYMMT9tkwcex61w+FcieoiYYxbnpUZkqJCADlhUcYbL
Scm8zFuoxDc+GUDiHjRsbJAaQ01Gp0yT5suXBQ4WFy156qhDOvbN4Ih2Z7zgyiWXftTviOcj4jWy
+WuFaq9KBylOFYwtWqsdOpbB8JCLpUMtl7C0X+/liGxuo5YJfeCem88phWORZIszvlJga2bjcS6K
3Rg/swOW+7urVf+aF5vyWHhpRm54touNld5ECB94h4dJ5eAbwuR1Ad+a0lmgt+Eo0bhWPWpF3JrN
K/wcQdeuMFqhJI+JwROnTXM6uZi6WrIc9WI7Xd+fxJbuXf/H01xkadp6GgM4tMwH6gEqnaMihrn4
vJZchvvJr27TK9y0E6CFKnLQ5aZ80CHjczhY4vXW/z0rQjGrfQfW4K/lLvosElGS1nSVWe+0QC5w
yyQsL5/Ww+rrdTsadmuodkZXPWnpDe99cXhHWtjhX69kbBwUKmh4vCOHQzMtFF6Xu0L24S+yMEFa
1D2kEdFOpsTKeVcpyAjWWk9GJned5I6XmKBTGne3SZp5axsgPVMuOLf7wrw+XolH3b/WMOYskfE6
PogJpe/EyuGrR9PNw6Hn4rr6lwQ5OaV1XL2BFJF0EQShnHiOnp+CBJBhCT28D6bXQZEDIoL+D1yn
tTBptPWcidvI3Ll5zPQSpIwx7FcTsfiVDroQ41OBAIjnP00l0yzNYSvxmw8TC5QoxeE0nK8WlfPe
nQw9V8WUZNYM+CySHM7hYAJGxooTH+PvTV40EsTZn2edIHj88JBlFxwmpOh0M7dl9vXoAIaiQASW
xHpfiH6WpMlk19UcfyiA+l0TVNI/LTx9xgayEeVJxyP8/tFYUAVtSmRtd2SpKpENGI8ybDXj4oSo
jJgCktWqbfSefHFm+C4rRgRxxFW64R8lqSJq/HKgEmfYshomMMvkL4NRo9Avpx9LJBj/YdVRo1D1
mkHT2ugI5CRiOhaQkfWmS9KXJqmNNU6f4xdUplaNc8JLsMFt5cfnjF4oovJHhjoEYUo2I+b3IiTK
TggeShOeOj/xuiZWhr3pTIZUuoyS4goB1TqoNcQTNric64+ECeHIyZSN0Wbb/fOuNC4qkebsafmC
Zthw+YnfmhWMTYvK9Iyu8Ws9t2XPQHr3RHJCObT+Ml7+3XRI2JQegaMxEIJk8kTMDVC450crq3m8
xJCkjg+FfyNIouFqVUFLo0QWvmB8Zqk561ZPTMpA1XkZLZ7oXSWYGqlLKpvfEBFmmqms7r6WTnH8
cJnMJoZCMLOjb81DQT1rCQgHPYInWr/S5NA5EE778iJlVF8v2ECn4B2sJay8FOYOHSnD5ffMuXAH
1UspxEjMecXhYolnwr6ho3AixOGwa3H1vpY+BGbGsOjSIbWNyC0vSaePzfUPVqWk2DjJNGoABezd
0Yt3UXoAfLm6V6gHj7XBe/r9VqSac4rEC1cp8tSm6iimph5t7EQFexadNxJQPgGT41ixw76Z+hxN
G8mFC8vyimfGI5b10Ey+grAyipfUzrR/JZ+EoyahbtRiwRXNOsIFPGpDllFEdK3pjtdQPTq/A0Ih
by2paC1r/dOG0r0WfilDYMRDQQAZhfTMF3V9WdzmCGgj+SAvYfkc6lC8dsenDyThGtxDWwXgYb7b
oPV/5IYw0OxE7ZcK/sBf2pT9KOdIKp9s6PEvdAoc00XGA2Y/8+A8LgxeWeJouk334SSLAZMzlVRc
+EQr+vt1IRv498ycnL8OgC+d6kckW3rCSC2yCYrxtBUFNpN1F0vTPPwJm2qkt1Xwfsq45LF+RDLH
kTC5gW/mG8X0K0aOaIyDhYjfBGVqmXhctkDS6ZuTjEAu53J5zh2M7S+uWSuskkxQ+nY0+2zMBpks
kuZVM2ZIvhm1poBBzF5N9W15per3iirAxLkFSJHFSu8sfgyJnFGaMngQ4fcv/x5L1s9+jtowK2U4
paCZDvPKQxxrC3pohBZAN4camKcNuTB8tJu+gBO2AQXgtIK/uuJMCvMqKY1jrx2Q1mCRW1F5j21l
dF2qhCJEGjtisiTe/laqrPJRWVGIg9Y+Asmik1pKe2LMufHC7N9pMmqje8xVBsA0P7AduMYLVqDh
MnlLSUr9EpdO5ex0s8IJZ9vGZZnTMZynm3EqCJzZ81sl6fnRKK8All26wN5zRxMi0Z/45dJdhAXX
EFcZcn14zl+NHAmwwQz6DeVre50uP9QMHMIDBjRzv/pqIZ3OjFEEhbkajPkMheRAyIL79NWPjOKV
3jGpe53Fzgi2TCHVLXRaxB/TcJPA5k+VYa6aonNP3dCX2J6MH3dUy7NK7+fLwohEkVhpfzx5pS1A
oSgsEzdBlFF3Fw2nsLea1Tz2bhkZ0Edck2819epoQglz/Bvj7vaKLBiwrGua1pc8MOLMTn6kdEB4
ZnQIY98cZfo0SDIOoECjBY7Djv2Kvk/YPb+VoUGl3qdKz0LBrCz9hzH7Dc8iBpGJfz4ZwyAw3hRp
nNuD4DxGASZ+pRObcRkNPzBwFkB9DRyaMsgSPRZACK8aW7mv79ew9KC4puT5Va/r5JoFAVUaJmNq
w/EVGiafV2IvaZP1t4EPO9ypvYsoZsTu2YVybFvZvo4Kh+UKdGOtbIMFnebqLX6ldWCTeoH4WItB
GvDtLlQbv320ypWfw+YiDxY1Nb2qewpNzaHHgPEj7Rv0afHPTmrk2o79/lVKueyERqo/NlYqQLKV
5eLr8U6cm7pNAxKPgFsXFCjB5c2EpdWkpEOfj9xJenLW7GF0qgbxITDTpDu1x58DusWMFuNi/bwI
QfPPabrPHVYuCa7UrSOgt9M7r/h/p7ivPhbsAaDXySINueAmsYGLctq0PbEIL2AB2D7PWbsBLrss
8LctcYh4cVeS2pk9ESVxylA7CpCCRWrdbSELT9bv90ZMiDA8axevjDP6uACxRUFf7AA7/x5pjcvp
/qVN/NfclLK98RwlV6RyIGMyO8J1Pu8er8R+fwjkQeMI+1Y2Zo5/1b4vVp6akrtmq4MlTayEpotA
TmUjkZLEI5QcosduqPQIycsgNVBjcoOa10MbOdtN1EjjHzmwXnaMewPUQElTf2XinKY9VgFhioFg
St7V3tiDj9flaB/XEC5Z5IpTUb7ZVJRWSIw0vrWn9RZzejAJo1VJef+J+L19YYKhnhdyO87pCR+s
51fRs6ua/sLGHzkjyvNPAtUcf6f4EA03HP+k2xCAZ+EXNPewQwGOHXL6cP/q7vcbY856Y7jLeVLD
sSDobRrcbSvTPaKv6qwGk75G8gQqb+gcoLpGxLsj+h743b+6PuQpY/6Jv33bHiuJOQBVvEeGCIdX
uKVV0RZqQ6Kd6ANpiID1oDaoDNF2uJLPVL3m8GCiOvVSpm/U6/ywVA7xlA5Dhgz4uF7BBg8KOjmY
sEUqOF/gx3VTbmSshPBSPrNlRYv7qGUImERydgfe+B3zjFgUPIpsKEOs6EmtA33QkAsA7R5a1/7G
bxYCeP4hunCh50Slu754SJq0nrghigZ50mTOtgxklVVtdVObk58cbbthDAvTtscmBTB2rf1WC2je
ZylQyRKKvE8muX/INnp6v22ZwBThAp4F09zrU56dxn37OJhAM2nvxL3egr5lF27Lx5U4TGxUXZNQ
DkO5U8f5yHp1xuw2PSLpVt5rEkwdMYuEE2yFtANQNMWfr8rk6N8kxUmxj9aOORrPMGgg90dKj4Gm
whh8ZJIPO2gGUwZvMFwEvJd7tVaR/ZBiX666Flf46KWPT9+4Zdcjmcku4c/+Hgbne1UsNjE6AqJk
JmMklh5xfGRLRzYBSXhRg9sLOAcMhCLLQJQLB21zhgJUSvROVogtMkVIXBNHkRAztB4EHS0fxVdt
U4d1FnyWYxN8msaDjeR7n3xN3YizFUPxzaMBLRzAP9IfKVqTYvXbpbN5xJrdhGJUMK7sy+tg8ZOz
54JbgZ9/YZ41CvmUMVPFlvB5HXogcf78SUOF4Lu/HayIFVCwv8iJWWzRhvzm2zLnkaSjjZ4tM/V/
0jCc5jNxUEKgpb7D9rHoGnwopIQQhCGtVOkZcIvRjUlVIoTQAvTfmxSD4Gi6z/h6N2h7NDafeTaR
zqXGecZksuadRZU+BQOF5Qyf4VNudc0XklRhSSqFrcFIM/lXpirjcG2mmyH/IjGBKw+H7NHKtgeg
EfQgNlesNBRhiMn5zPIWLsohfGRT1xCIHt0GDlsOWAbFdpfoOieNLLe6So/AiZsIaLzw4xyuFObx
klR+nrJkd6NqqAoDzoMWCGm+EU+bTqKyIU/Tcfx6W4XA4Ju/67J1Wr6M6+jW6wBv6AEwOGcNBpaz
6SeeEWfwhghR+sZgcoAXLY+Em4y4ywJXrOGs/39qunmCzUpL3tHYpVB7qdETYC+ZM8emL5orwxYA
zeuyshZygwb8eNvINRL5qEPKQXfMPUAKhNU+eyYDw1QnZ2eYprX9wMSImz3dXRyBiBn3+yXat0Hn
2eVfrLrn8tnqSFQmCBkynu9SuVydagaOBYZhqfzpxHroKJZLVk06Pi1XOVK0LR537z62DUDVojm6
1huk5iegvYSewgsOsKLNySNwQEz+MpX9DFINeiWS+3G6gzcNAB+Z0Na+ImnZ59mBeqxgvRsorqPG
Q96xkn0tzMcRx2WqubOaO63yaqve7oWSPdq2Bh0W3zpXN58kMM7162diQViCOydD1487x2TQgXZg
SYtiZxg5xYYbpVNJHsTvGTnk06V/BlCiJv9aOYonfppij90QwpRNSZox+91wJeXRPGGWNcKaxcug
TEMvSnuV8PKMJaJcRILhRrVzz5bGYLF67yfjwR3Z/nooUSDbsQ34+HLSvprYRYzwkRgNkJNY/Aoq
rpYzQ3eWjOHZ1j2iHc7A0gazM521TzCGxJyxITSFxdN37CaWVEGXCbwVP184b/fZk7JXVOFYheM0
t17ijsTETbALY49WFFtcqDEmkQcQQ7LF3s/ratPt+fMXpVkImMGiPQecUxi+007EUi2qzqeh2Lkv
XcavraAuBL07ksASGjLNIVA30He/0eozwT8MkubW7kUrQWlmEzMc/bAK33CloBPDKcjbzVDXTaWC
V1oUkfnkF//W63vg00+lny5Svca25NAUX1kt8m8uqItRf2XbjRTx+q12hUZyX50O8shtMIXpnsJJ
rM4n7kul8qJxAlqiLM3YksBM4Aahs6CAtAdNgZXvAZOgO2F3URT0OaqqYcxRhYH6PatZ5/OX0bJk
3vC9H/LjmxVd5zmktvTAGXVIZKMF5eOvpfF1slTJwILMyTKswKUuqggzNEsCSW4xsFBw/YnCVPzN
sPta2ZFJ0RhabxT9SN9tqeiKtnVXHBQGwO6df6z47o9D7sgMZE9CNOuHJjNQLAhdCaGWdY6F7BcV
jCEkJsIb3K6q9nVWMORG90YREsdy0hibP9THarNbDjCMHjxphwSdpnl9rQXSNVqLwf/AquL5C+Vc
BIgS3HzNQ9yuQ8djg0+zmED66/Rdh5q6kqEPqmD9dwto1ZEX37KVur1nIjZ1B52Iyu1FtM9FsG3q
l+6cOxonGQr9rGsYwGGg0McEXGfZeF6RhlSVXLSEuvNheoR1INi1hj2miIHfyvW9RqOJRB12Vy/b
nu6gxOns5AcwpA4AGC0v1rkK54fawNL9LE493A+G2Nf3wRnqZls3v6SdsC4hw1olDpF7FRxzNRNs
fuaQD+bWCxpQOSaG/B6S9pVNtYlULZ5/cxyGEx+fGOsHqUicHYPYVyHJq2zajU4WEFfegsLcOtgV
Dys2SVpu+jbHRCTN7Mvyxgn+OsQiIhLohjSG48+h8hJVCayK22SbyoidMmlhZxyVKL4Qz6ouiF65
WkCFVSspT23O1QCu2+/Pdz71jkdgRz3eUA4qDSQcP/gnzE3l4T4THEK4huSZXRdXP/hFakVhFgXb
SKVaYBENTK+12Ctye2HkMXzGTFZYHAfKknHM3qp0PklmwIxDanPaDmhbBQ/x51HuI8WPB8u1AKVN
KmSw/9lpr8hJ26Z7dzm3VhO5+HAYswqQivcHtJjhRChf92KVFT8yawASOOGBSrwiSg7hj/QXnxo3
olup51soqJL/PeCb9LXph70BQNsIMzFxquYThSZWAk7IjP3U8yHSb3ehwAA6FojaLMjKkkYifJyQ
MzBflLHKnrFtvtPav2s9mPhDzPrFDByuqhhXv28aMMf4AuWNAXMu+/FZZUL6Bn6c9dKk9k3QhiMn
V0nIVeBsEz7g2xfkaHnvgYzxGqWPfkZZkTMIhiVyDphV5tllV1E18/YMeKqupVqyo6c2wu4CYRgJ
fxMtuYJ6F5vlHmPdnn1NjlXLgcJVye0wJE//fc7kNKxLqtPQNBX+gP4W/Hjh4QhikxgllXCNec+e
0z4DG6yox9SiFYO2D+XAsRMMffoH3jtzy03I6lZz7MA+0rbj0M7wKQdsov/aCpUpD/MEVbehGjg/
+jc4Boqz0xyJRJp7F72tajjZGy96feccIHVh9i+3kux2X2d3WcPDmH0R4Z/UcnmWvW/9lJjZ8GLY
1rBYMMgq9hb555h7dqUIGAbt7p/Ge/s3etIi9MrHhJQRKXsMsqBHseXKx4W6oTE6xONn1kTJUXDZ
dA1C2nE9KwxWgjYM0Z7h3DeYPBQOK9yS1YHprZ4SQ45n8GxJDww1PJVvO0MVpG2Fxfw1zLLK3SPk
kcEsbMce8t67ZLqGd7KwhLoSDKMnZWTGoMWljStazLUDkjg6+sfr62IDmXLiDlrlYUn8mzDUbEhw
mOX4JTzroHg8oP1LD1jVCoW+YcXOBQOla+3o4NAfSgh5Vl9ftS0u8VGLswD4Ocop4pK37vKZT28R
CKqhnWtgezqR2XNOYYVqepM3TIzM6SJIJG4aNZiuJzYv3DJTpFxkK75axXU8RSwj5UDrw7ufPr0p
Qbf7+TWtq6M19tmgVZ1FoDCOxxt5rmGGlxNOAE5TBBxXZ/FyOz6IICII46/LTjDfocK7nKr93ZCt
/LRr1OdwV6PBNrZhoVLXVot8nLVr33avSP80qhobiOPU7kwI2wzjGxQnwSONPi9UClNcwFm+2CBY
MQZ0ieNQ0W6cDmSMYA0g4uONbnRTcI4uJY5dPAUwzue+PldYv64K9w0cXrAz//nykfm0S5QqO9W7
Mmc9496oOoPfiuXbWmM2A0SZ2JohsWXtQYKSy7UR+lX+BIJk4q+ohIb8gH4PTi18ZhPK0gJ0L+4y
T7IK5zab7R+Q2Un1/aNwIGi0TXuzKTQIaddADknUkRDcQiZDB4r3v6ffAtMsl5p9Zuf0m4rQRKs2
EPEw6ONfYaQxpoLGn25S3iMTzXSwiR6BbHdnJvNnz4rJsgcdqSZwUmJsmJNSjea3yCKDhbklFxko
Sv2RLckcyI2P9oWCNvjA35D0mpidHVbITqFVAbvIAW4oC0irriZsC/hB5cxhsm4tww1AXF5dUzjH
YjpoGPpTXxu2vEbFgToA4I/hqRP3Yice+3a9bSRoECUogK09t94nAlD8P+88JZ4Fix8F0aWNQOxW
9q5ROahsZ5JF3OqJXVE5XWyBg4bBmFh94bpnsWd86hJBBJ+opEvBh/fImKRz+mGFB1/VbMHJvmdZ
1qDgpIotN+8/b9OlEsVsIVPF9N61V/KIMxD7AiXxi0QO8gWaZhE6JqIVMI97aVQ4+tiU9ZRmVfzu
pXmoAQSkurZIXrf49DW5eNdxA9+5412FqEbTedS46s7q9K3VBnc9B9lWFHMflF1jgex4rHS7mrQn
JLT8h7uzQj5/STKkHeLwStmeczeRK3Z6DV27OsDwExtVVDFX4/hA7yI4eH7yR9rz9mGOa3lsd4HS
Hxu4/2JU6qSPVEmrrD1ejjKVyoRDFZdDX753ozMxyDrZRdLvtSR9ywl4mOJRumWSfJLEr/I1wi9s
+EmishSMcFmRKngWwqEDnsTAvsTtS9L8KLxOiSwCY+tDf7b/nFeHq5B0Kyx2uhWZZ87pPrHPzEr3
gYkeUhHSW0Habx2U1zCfdhg5LJMoBPOXyuhB8hXJJ1sUjjTGJMplRbCnDZA5aFBS+lsKNYiUHpoA
B26LsG6bNnvCimHFZ/1D20yf9lFbHEGI3kQVPr9vLDh4AUi4WF4SSK1JgRILqPSEMoqX2QU5A5jS
dqvArQc/oG+9VS90dNcYoC3GJ6FVuXnpKprB11FqSZ0z16O1K7yVFvASsMjK5mipw7qm8mb0IsgW
4D2ZTDuCoZJ+BNDmAlTPrYcgC/t+xDN4rC5CP36Wmg1oF60LrknKMj58IhWVp6dwCzW7Z19AnTeR
3yirLoTXkO/Q2ImwC3uWTr6vH6Zb1vXusRsoPZHZ+evz+uVYVA9TmZnpM6VJobpAHu7AjJ3uGGij
ZG2WykWMpRPO2uSKLb0uyzclzWQMia/7Y02E6bAV4A0sRIYymYFiIDJDqDmVKuuysbAyZ0VEXu8+
kZH8AeTWUsRToACEJjB0KICIpBESCFtg/fQLvP5OercC+8EJllyny+HmvJshkmxYgY4NRxkd3CQB
0YCmwy2d/g3SwXrLtg6T5HMkS1thWRksKC/W6Qf7TT2tsYuuN6On68JiR+3ZndJ4smHAM1A8qmJN
EvvpxYdBqXLWojMejbWv3vmIQOOmzqZ03mj+WO2c64Hm90AUZeRl4Br07cn9YR0TIuUE44+4yP8m
px3NLeOza8Q7Dfi07h/Wbfe0x/mfPU8+Qv8HSebuddeG4rHer75/6hrr+OwNbZHFKyOfc6rc/9Sq
s8JZaIpUH6m4IBEg4RR8JLPOjeIOEK/K8uy743dNmIdyP6OofMKX/SJa61pl24zepTKDt6KGjTSY
ig6Xuvw/BiK/ndjmx8gDPnYoo19PPNPpssBpYkd2KjV8uNVZbksvS8CrWI/KMb7l3pK0NGh3Dren
6Y26Dc/wU9Plrdyc7eV6bBjqf8xs64OFkc5UPAwtcQ+rnAeV8ZqR5S3a10D/efiWlsWjR9BvKv1a
I3w6L+EpkRJe2KlUsdRqYpnbQnxXJgyG6S3GyAwJuj4xGeNBIAgsWVN6ApQkbDjcRWdDHcN8eA1F
dEImkoZtJeWoywv4LcIB+6cZ57fceAoQalpM3aXJsTKc46ikXcVOAPnSxROV2ZGhtrP/hZ0FXF4N
2PKtalN1V3J+IAKxmXSp0cN4bMS1cCUXaOzDXS290TNMYaN6al49YQAvxey/0kO/aBk9YWKkaWZ8
kuIqhOvfpzi40hXQkqV+KKXclKg5qFUr2qy2d9hv5021Ar4Zs/x29bIQZypW5iS/fW67DXC1t9ED
FPc49+F1wMVuWtYG0ZtfFyJCvIs4omqP7638QHny0+SGpzcPz4YImCkN0U+kNpTpESkmHuVcd8LT
ZBj28tM4nYJicfSu+b6fs1oiJCm/1wZjucskoFK5LL8yerALpXfF+T3BJjsLPCpogIZEXeApHVyM
8izVPKb/Lodw5p2y4H028qDjNjBdp8sjEolNaMicAtSLzS1WOY15zd0ccgwmXHQSoMXzLoq1ohKc
P2fs/UBvi5UCrdd5N6v5mhoTS0Zv59Kr1i+U3i2TgimLtTYCe2m7L4GMEjN3N7TtbD7dRCrEJvY0
dc1LvkN40L0bag/WYT0H91bSkJgrFeqZZgRAVwt4K7pkNa4fs7zMHqi5zgUpEGcgl739nRjbuplk
VJdarSnaIHqOJ4hmdJdJZ4tzezxM9L2huVQgh12NbAm7UgtiquUrfVdVT/koDOBKfuJpjdA7ixip
zG8RgHuqdL6emyrhDLeG6IEtHZWLQgs9ZdBEp7+KcjYM9Wn1s1r+XcjA3QQk+UgOLcjwnlmbS/G6
BnSy46R86Jp/PoUrvy0rDNgNiJ4JE5iaJ3uRspFZOSZI1Hv7VyAe+aEAWA42X62jSl+qJhTgw9al
lLBm3/YElDMFLveg7cT1z1PLCTmjnniqsgd3K4M1mxyP7GG8XEZF3lJq/bQhAcTsfOdvd/+keTkY
Kv5Ng6ASM0RV7066aJafIkYSCgI6R/9DqrYwLqXm7rdHr004Nkjj61UatnyPhcRXqpYLKVZbWU0J
CI+TmT2qnOa79yDQtyy17gQHr85yNA55TmKNh+VqrGCxDCKd6M8e6+6NYpsgoNRhWMi4kZM19frc
Fbvi/nOU6NsOfyIUMnfQazExKenzhn4PY00ZdUUk41mLU1qBA/bL7ebCPCL74OK9h0zk/JlfBepe
LA9IR3W0LdoqclSWb3V0BbZrO5dlJmI6w90EwF/xaTNg9AxZ2kYBnHxgKw0egpN8D66jc6U8fzBa
/FCPqyI6wkxJ10k4/MHXX0S6Ni62Wp1V+9aEsofk3h4L6njNZ5MHKJptsW2aIU60NaBpM6xejEg6
nr6x18GOuK5y9CVvmdpWISe4uMCgMQDbmgfWf+FlWPigACkSAxzJjIRRVeTwQUVdqnwYNIfUoJok
MjuPryM4pq+8+GhUFEwEOkUeQrmgxRIasy/MsVwS3aKsDID/3aRQsZzy7qUfu0TIaCPlx3khXWX3
fRGiPBPVL2QV9m0/u/KG72kw3ayn5NVJ9e3tWQiW+eKJGdriCIeca707Ic8Q0X26Fra8r13fqRb4
AWouREcng6u4hCccRJ/WwCqNaIddwPSIbH+7kVVRcR09XTKEbgxlqzCx5tmzLhTuAUTBxrskHnMv
JsK0L3tzshEdZC+nDMVLIWQVyvmNv6Gq9gB0nUDwFzSADzTBl5G7QUcDspRoBu9p56i+kep6PzTG
FfRiDk+/Kd0wpeTmSaJfXQ8xqxs9AiuI8LVgTVZeTN4mzOnwWsRMMVPKzkmPsLTAark6inpCicns
5CSOLcpb8DzfRBizYhMDqeWqyq6x+ZKOxl5ynlsUM81AtoKX80bcKUZ0S5cncr9ipZxpC2VsOo1x
kaBBoM6tRov+D9fTnEJvyKF/FBuBfcHqOhXDkYLXP4OCunfD6gZQIae78a+hc5nqLexXI6+XctNp
OS22pdMUbvm78+bN/ePxCMRBET93h4KPkyfwlaFXSFoN3h0N+8UtamuH6PH8EgyHCEMEaDdHwvkN
wy+9mo5MmpSvqGEJmb7el01ObtIWQdTCiI/oXVBGtA/odxcmd6JM4NCtaPf3OzUisdnnGHhs0Fdf
f/Lnga4Ym8BQaoelrULfppYDZ7FN0LQ/RocfBYuB9yUd2vljuHtgHYuoddmyvNsKO0CD/ZIUOwfq
Rnf5cFIcccXOKXu5/tuLSdlefw8TAUm2CwwOvvykbqPB5JCSP1KJ1mJZI9ejsqsPsiQjrwis0VK0
dJ2Z1pBZ0XPOV1KDOLAqqayA5wSkcPx5Tf8HQfuK7OyirTtl90FmABW8RTOABNyqDw2Lr5MjLFWg
Pq/CRlqkIfiiny9Hee+PZjjiJhb8YVLuVrCrLpW/TkrO/uPDHTFJ8JJ5TDO/zl3rnLAiV8/K+ppO
2ib8OOio3CCXSv6MDGmMfYVCTjQFQOtP2lkwAxWoR9cjQTKhuor86C4H2uIFcOsb+CE8fVQLNR0l
0pVBKsgFpjT9vc4nrS1gJOEiL8yLexhMtSjRoEVo0Trl/7oAjj1cQh84+mI+pmIfNZFUEcwjzjw1
Lxd6Rw54hGQOq1f3126nl2TWNovZu1Jhomw1YdalcGcdN8ASC41NIVyYjl8AR3HyrYkpCF80IJYK
ul6tjBytwiR/bleCIFbVICHQQhkhM1DSekCGcgth9PN//Qwp4KnhF1U1OojdOhPev2df27Ca1W+m
RlmhQo+8KbC3hUtnYEEB8nocgu7Cbx8agvG6hUzdMjggmWBAHpJy0WWb9BosNOrIayrWh74FQK93
GzaiXb27h7QUOEHPGsKNjObPfDE2k0Vs77l2VPZo9YGbvpdDAk3PIo4DAFlrj/P+eILv5qeJCri8
75GwoUKfLIeE9AvEX/2neZLNnB+uRLY/7gZHAL6XS14bP5FyNpctIAjxkM+RSRKH6HK5PHqG52YL
NXX8HRY1sesFs2otU9NwZg0LYMHWdypMZtTt2NNRUgVA5pmi134HGHG1qVK/ZMOViwhOdsl9ommn
ig8tOc0Wptk4ZRqE9Fu5q0Kr9P12CzxZChldAbEWHtKzyNQplNfUAY3eB2YLTXgeArnGplYZcJwj
xMilxWsQkjjl2iBvSGwIJ3bdSWya8n8m5zRzdb6RH8mFf0rTxRUayC8sMH6eXg9wc+u21PhwcZIu
UvbCbfF2+o9bDf9Prdp7YquMvCuxW3/1l5AONlF4JTitsHvLuyHK/Xi8S3uysHhP1gZqmXaG2Us+
g8aSdlF90ukDsniYNxwJgX24uVB81jE1aFQzuIhqwcrxZ7wPa0+Li2aXWy0j+JiMx7FKygvMJDCs
zXrJEwij5aFt9LLb+hlOayjT0EmDZGWWQh+jRN5E73m/DEZP/MMyGH6sdBtUrnKC0fAc+ejq6ct4
R2VYbx0RQYJ4oEsymcTtUhPSV9tHOwVMi4H8zViSdbXYGD3fL6cz1DHRUMF0D/Tv+hF4AM0oDhdC
ayzZp42lRHXBJkcGzQ+1/M1bKhg9WI4Hw78TsvIouDRPjcVooLCOD1V+Gjv6whvclNhkuP85iYhb
dOyE1hocWWhmbTWTpDFtF469Dtkyz638nLd2WW+AUx1wDr6cCbQVpUrfkOu7k0qvsz6ETjT8BgL6
z5eCCic2cPHei+41Q1E/q955c1FPquvH7tap1Zu0DAdpBaisHC+ahySpDCLnkC//NfVltwjbkhkY
4BBB/3Y//Q9JnsB6Vr+PGNA1FiOvoAvgcm/0hTHvVW+0NgpNVDajqatPozw3IRaPuqLahDkDip61
2UjbU+1uCuN8kqoV8DnCsmiwJOOi76hE3vd/UoHBLfa8SSwsZFY1sVHcjxipUhlRww9voSB5+yYS
A8WkSs8uyboD4OSuhVabiwIZPH0fsY5M94a3BwiNeYJNXRMHURB3g2KKGesHmb6yLANVfh0E5jkg
UtpNOWXXvnGlXZlv7ecWPoA3iajqhpPVeQBQ6ADC3A77QkBsf1MDAj9X4SQ4w8sp9eZ66QzCAVUY
Y7Po7S5riPnBpqg4cH4sjF7CkFy4HG1i9S9lYFvwU3UjNsdpOuk5e8aaZ7/GnYJL3niAd8w1SxJN
4H0QStFQXI5mIJgZlctB90hb5e+UPcfVd27LrBZvrhwQaOqb4AIQPv9M3MOYLYb1zDYivs7yij5D
eAieMKkGKnV8ZCpez3S4Y11jyKbO8g0XEvafqxD0CiAvn3l8gMVqx7VyYFDytUPkxOb1+1f0rF6C
20s+ALOjgSbNusA8enJRpoBXh3D5N3/VImzGgpW7GNsW+LfYkrStwfkjtwn6AgdaFMmuIhGmAmcq
1/NfafoJAeHBkOcktV1iAy7xX7/X9k9wOV9D/g5jXVFoVRtrq/zWMsnlyHnfRF94SEElNbqTtHN3
xQAgrk9sdTbD1NOq2Me+bp+YXO2yqTuajKRj+7FsgM1Ufn0JG2txaOYP0o3SszCvD9ADOfEVN1Xr
ifpcD8ZcnYD88OvavMIbn+ed45DQUZKpDrTs3/fBBbAHPo0LZned3SGwqqY6oa/LofNfHMk44TNi
JByq+t5/c3r32z+id5QoLWCxGt3QYSi1sdMny7kdrWbJg4q9nGqry/DXWdGPRAjdv94oqja0Hp7F
4M0lN/Q2KAyBxJPBmhWVzqaEdaxCTQa5tGmODCXXSjfnI1hYrHQY6eHydhSlAAMnX6G/vXB6sn04
mA5bUrw3e+/QR6L/GA2IcJXXOaMyqkgIsyL+TTXMsPXl5BlYT4z69WRggepu5EpbSWjwLIrCG3xw
vwIL9bTzvQyNj2d4JwgKwUzeCH2kSkJIxa948xoa5COdH9Z8Ot7cLtGoe4hWT+OI+sN8ZzxC8HdF
iv45cZqqQE5hG81UQhzoarEJcjg3FTQquOUSSFIwojATFrKVrF9JzbCoqhsjkrkne56xWXl/GC++
oG0b56SKDveWcZjB8Qlxrq9OXSjgMRKKg7y8o3fN9zI5Dv1DK9JGnPzh/wW8nlms2JApda1XLr23
sybr973UU199+DuKgIi9aM/bmAkPcZL/hZ/V13eVfLQYlZlZtDE2DQOm9Wo1ZBAm5WZ/EaCEmbSd
XS5mBsC2jYP1SgtHI8AWFN7rbnuT7AqnmdPyeSLPWvIDtYnZ/JbRfDYqqphpQDscakDpyemKeEk3
fvrN4Ah4T2lKr6x7lTZ8g0ZXoJfNHqJSsZTyshEPoivRmamSe/3fJovAqQnYGC/o2ghOHsrHk5oF
Cc4glGgicaoYfypNXkyli5Ywsiu921YX10F6KOAKtrYjFQJvNpj2YrxNKSmfC3lm2Q9566OHkTqX
OgLGLrAv6zrGLObKokXMDqSr8ycTEH5Cf39+AX2bjXCOUxKC0HdrJ1AOiT4VWagdA0Ex1tDm2S23
FxdRAlFpe6f+4okG50WWWCVcCLmtql/XXYuOq1DhLJ+sAFxOim3LAHOWRr58yKVmsPm8Rm/26/Hn
moOc+8jgBoikzJvpxn8dY0ZywTFzPpQvk9+ftsA/ujfz2tvFYXarYeRHb6N74No5r+awyxO//qA9
c8n+stdrOTNLAQy43OFR3horUcyKd2MNyoYDiYPRI6WUjnvo81fcIteBOzH3WDvtuCdZVHEs+Zpy
xm8ehja3thiRioHXtpLt3t0QoEYMJOFN13mKqR4ByIjnFsVolEAmXD1PLy5EFHuntSQapDcOeNUF
xlE/iVbYE3cB80On40JSa1lGPM8ga5Y5su36/b3uqutI/a8dG/hf7MUmRsrdlfWb91dCDQJlgqR4
BG+qvBZOkl7VKL53gRCRu3rp58z17Mbg/8F98xH68WBrYQ/suJA7Cdg2Vjy3LarX1M2cVM+OSK9v
PfmufU2LIbEkjuaiy0CRlPWXMtJwbZtgiuKzvDHTi6oJ+zafDTih5LXKQ02uoHRjh8PfCy79qI26
BbQ/ipe4OaDEososJluP62tQ4t0lovacaPvTWw+yyquKheKfFnr4+eIvn8V9Cnb6e+ua/uip0xps
N92PWhIX3YnrCkApxjUZmtCOaYCFv/+pH3BwKfq2DMYdS8ZqdboQPmkTnPOHXuFkZnt1cohl7NrP
9BJMWJ4aObExczwkINlr8YuDGcLxU132+fK7XEAqOc6FOYtNtrW4SClXYf/7v63UI7NgbjxgCCra
ppEkAewSpmEEWDyK6ADbA8X9uw/ZDyeXLAt7NqUqxsGLI2rAqOJGnknrBENgmoqFaPJ2n3TFSzFu
lK9ZIDYVBVu9u+XEHPtZugBh8nQG0w4MopnDfdfFER49BHQaBljKyrjjBiz2Cu8Eo6yEg9B8QzmV
al2fLYvW64VxmIF504oewzunRzQNsPGYMcn7V3jxDYfKjDxPeWDe9c0UuqnYk/3m+7e+ykc0XpN7
aNmserXkcNgnEoyS2uD9EQJUDcgTCRKSaXWSBvMXKkvQ1ZCDZsCT83b4McO00RXwPkgv+4wn0RhB
jKFzOYUwAL/X45uH/Lf9qewmzZx4fX+Nrgri3IUJJjlZaps3CeiTazEQUx/N2E7Cs2OlA8A2Hus+
XHBXSUOtX61aMBnJwfb6cDxR8bV90kQ9d/ZnhvGS5zvV6BDM1ZtQj3XQAS+/Pu8m2oxOmCgfVFNl
bCbg8eZdGMielOwTLzYM7KRVIcPLGkQQR4GRJrZLQSZOEOH0f9XhOZIsKHyxaa+6XE5l9PeXU20G
lzBxlCVXy0DnE2MFcXoJ0wgLz4394mHT9PhDXPghaYhgQ1uBajKgaVqs+9zEcOFUN14THiy1Lvok
rTnTpSgyOSMKEPMAOeaL06YLgiyEwHN5kKwVjAp47Owl6IYNDbWyD51T6gbp2svwHb1hhStiiPFQ
mtmEYMnHMnuRyc5ZJaMqtFeKLPpIj0mGI5ezEkOkIpSB/nozG88ChK1FyzFPDIFcMyID/CXGFt1s
r+E6u53sebLbCL7t0aNxCMdpbTGpxGNTJbVIFs5cTas3hKR/9f3ZJEoSxMAWyi+BL4Q8D8MJVh3U
wc8+PtIVw0s9wlfXZGKHlk2YiJncdlrhzToAhmdX6b2nCefru+/WtVLyWWHsosLXlr22Sa0shZOh
jjBGp4Ya278KQAmRmv9aDqsSzbcF8RccOiasQ4oRLRGuuUeZLxvOOgVf3xfRGJhcxOBKwiQ0iYVs
Hi6+vAYaERf6sLcofP8XfBbL/L59AWoCl9ZYXZM/9tZ0p6F0pfIk8fq5gH3KKlVOArKI6Y8ZhCAm
8/aJASTGIpwHC5QExvKyE36dsCcuvbKnlopD6Ywo0nZzIgD+X3Kjmd8m+0S2yhepAXAVeT6xuf20
OGwCwCefcBPEulxd6zCG31hK/UiS6x7ASMM9n1SjIU8XprU8TWeaomERfw4Cuw4VqtEV266GFfww
Xf1YSAG1+Ty2sO+erSrzI9kHjklbTVCoEbycmKoAG5zkTYbI8sdSG0PYTMTkA7q+1ObKqWnVf6AZ
ekfUdcQu1YWpONVur7xK5H9McTzjrN/tvvxShXrbFlfaoyGH7bT2J/OEcVAUw/NiLAOUgeIwkFF/
6hhboiNfCu7eYytQJ51X7xfZZAIj6ZwLSm/2unUbYBMjtIc9YeO9RDvo92XMW1vUzlS7BRL7V64i
juXYf3A5JY4Fin58Lle2KDRL29qOz+nJ4pkVmPviUk4w60J4pJ5qEcKd3UQ2c+tVbxDd+6Tlc1Yw
AkFSwqCAfkDjahNNxFxWpLToyINs+mB83Ns1TnVvuOOEssBzjcOX3vDN+IqGppJ8fubyfCCwPerV
qU6jXt2ji2w1fFYmwn19roAqes4QMWyIahcasKr29CFp7CjHDeixDZ4Y53iUK0YGKrb+AJp4VCTb
Te23dkNl5ZJSSVO/RIFdtVEA2YDnKl0F4T9bvqVhZf1v1D299/zAuBSzOMyoP0AnL6eQOZBHxfYl
KvMflzrcdai6cLK1nwK7SxwQJQUWJsH2kh8/ImthPFr0LNn1xXY+gtUKAGwt797D60BPhkv6TP4b
+/sce25jOLSsIKgQSorIAVljxTXl1eeW3ha+fePmQpIQpiiykEtF4uK9XaoXtVSki72SdZb1tffb
qRKnYNLw8MFeh9FjJy9w5/RXBpmkG0Sq/Vkxmt1Yw3HeJ6J/38znyNF3rPtH5rTOdfHb36sOWQxV
tQLGRjDB2QXSstwOY5frl8YQPx1lR4pGR4FkHQeq4RLKuRBiqhx0+9lTCRFU6PojD7s6SGCdrext
f68WkaB/l50ZEAd+E+gGYK1z5/s+hamnbsVlqz8Z9Ksl1gn2gLkvo78vAMfZO4ZEM6M40JLKjY/M
EkAKn0c/8LG+ACfAVnwCeoDr8nTe+XtXbiUpL700+3/5XdskaLHzRbhDIZKTTX7BHONNaUNJr5qr
VvJhxUiAR4JTAnrf6T67T0d0F2xvrt5WUu4Zs2XQ75d40I4OIvVnXMeZmCD2NppCYuoZhP0i8P73
iTMnJ9ovuVqL6KITVyqNPHtGGqXRKUqHQeRwy03jWWuogATpuYvOL5u23bNOvCW5rU9B4s0yZume
H2sQtiyjv1Da3QTAMtc3MJ+qjtFJdm92gqTMIuL4Jn0fsu3rr/BxEy8IdXtUnPVaBtkpNhbnh6Rz
TAX0FPnlK1FG6X7DsGqaan4u02n6YUl/xEcjlA/yhKXNzHMktNXdk6ULFQ8vNPiyl6hD4Rv4eose
lvCtEAWKS1vtDVpsDNndFO2QUcknx/BzEvJMtk91FRyOMskZ3OG6J9TGjJR86q1d/FoEcMTHWxmu
LNSTG+aY6FlTxzFTNQwlhhFBhZMD5yQbohna4X7SQShVgSPnNpsBTKDmo2kERIcPkKo94lYVluok
ieJvKFXm3BALcOBhcIPh+Y0pn2Ggu6Iy/BwqXKvWCiIxmofx7pNCuDfL2YlyaILrmKPAAOIB0SgN
WOQMvqp6evW0qlins8Ue0mUVPs4VzbbQcFqny7jnL52TCXpbrbh5ZW6CPTbfhj6yWo242JHfI5fT
mjaoJ/wsOJEORd3S/F3wCebAwIIz9jnFJQ8hj6VrJ0hgu9pwDfwhNL1FMA5NHtOVCGHnn+FixWJq
5R+Q+RpSWrBI4DUhIvNDWaqFHJl8e3hCSNaGF+svWzK0+ofoqrt51y8sjcoWrEsz8a06at4KN2nt
PfT/KOqovywQRDt7W4+5F8QrlMswynaiTmljTDbu21JINwiJsoRfid5UVJonk58lAKpynii7dUL6
pWxZWTMbDFPR+//WKO7DVLNCUs2tWepHYg6DR2I3vuhSQyHSBoETczd5RJN+gjyVTQHyw/MvbS8+
jpcVrgt7Z4jf+QthgYlBYZMJJWEASZCLJf6K//AOzhJ+SbaTbiTwY+3UMKdjTue7Pr9YhBljiXif
LqKuPt+3fY1S5nMAJnXqW+j3CyC364Bbk1aLJZsCUn0UuT4wicEz+BkSXO0EOdEgHo3pSYlQxEdh
Zl3Isyrvr2MttPZc3tdlRZYBoaZDNsz5zCzveTVpC0FyaY/q8hlqwyzrQhPzh8JAhQelCIW9eBNG
6uN+Q69O+1V6Z8f/vtN2xhyxWOtAS3c5RNXT+S8rZasSu+udWrc63EhTtyz7HQPOP1cjmNMRJh7Z
fdoKa37m+GyH709THUCuGiqBVV76IHFPzO9scQ/PPaaI2HZY50GyXLfIAr4g9jVA9DvMI7RSu80Q
T/s8KZOqLdIasKnmc80t/G+Tt1EvtSYRDgbVrJUpEyIcZ0F2gvtN10HjJL2LZj88NWTnqYmMHseC
KRaxvsimhh9ZMWSEjK8Momp7XCzY0gkhPe9PaXD6HUWP3urWWrJS8qYJIEpIVgRss0fYVc1b/45Q
oi9qWnSWfPGGhXAOY9L/9Vv0LjTsgFDcyCrwi9I4SRxz7j8tg9NE9eRNcynPv6NgfoxU4iCjTE0+
9qOCFSp6iYjJcz7yqpF29S2jSnDVMGDq+4J2e+ytS/A0GAhQZGF5UC0XMgxEFN+TVxyRKKwgTtAa
YWcEc1aSc5ZF0tBUqAyJkQepMOQObLBiMbHYt+VVvEzPelPRQiGDEKDIfTCmnRPbbjYN8mtleJ9Z
erMn2x7FvZS7Mgx27ELzKdNcLzg/7IQ/+38DOMY/GYwIJMY12B1RmYm7DY/AJmvqG74hSciliTv8
Ze7qnulocN9VFiDLDvLq8KZ68CKarUhiXbYxBsQVzcGwiG8k9Uqb6swTf73T6hKqzeEyIphYnSad
BMjYY8XDFu54gWVuFIu6EH0PEXoyxk8ioxv3MRyGg6IRaxToaiWalKxsx2DYsWrji+UIVt2c32vg
AWDVdvV3DkSFQhc/1edi6SuM3VEGTB+Nuf8AAXZc8+HuENYIkdkmuXhjSKhWeC1QF2kIlFoMZP/q
Jbk/XFlbMHc/nO1ym/4I+CxR3iZXrB31RaFVmJegn4JvT3E0tPhm/0nRtYI4q0lP4xwgAIUBooD1
+jAYZ/huqAmWRFvCHSfpzqewqX+t0d9uwGpgy3XmprPLIDNUswrZk7tqvvXoVK69j6WYmyVm5amq
5j7Hu4kfdIVgdumCqdjiePFc1mV0m1GPke1OFzgkpXU56aTxjCFv79VUSNy+ggF2Guxz/sxNFsnq
3YLIP+Y30nS08SdmYS6FUG0Vvrthh52tHlhwlVlBnA2bpGDpyolrf0ifB7lejGxosyDd3dGByEsn
6I1Fa6ZX/OyFAb+ISNB/hk75yUQgYnd6KrbOgim1tlx8vbnljXy+0zv7UGI1KWFqZPkfR8i4loh2
UnAW3mWCxXo1h+4cXDHlfXQ7NlGlBZVT78fnJ8DOwTNoT+AYzyBRVJDMm2DJEjNZMkcWI2uXikXk
7NPrZSx8SJO91i9+mgCW+pi+MvgK2GHmz57uHf7Yv2SVCqmti8NkQUl59hvUy/JG1n40YIKg699T
LvzrFPDgQPE49PhSArg8DccqWlemA/KfvKVwz36q/bWkLiW+Ua+cAO6eI8hl9ht6xTXglhhe8M3k
SdzcQsee2btTsezRbnHAo73lybEiBht2VGxGpPDxnGBthDqPa7sekBz7JMurEuaHJHc/n4PlIzC0
93kxaaJUwCQioQxEh27531Ma+dHtnCBFS09V1alWO76X/RMWmGKlKxCYHml82Q02mj831+/zVCr3
ze5u7t7wJBH2bWQgIEyHZCTMZoWkElu/pV99DGrnqCxl+2LvThE89sUGs+mK88mR86vyhREiP0tC
2Aty19rrMPNhMuMC/JO5GBkpAL6UgeTWShHnz3OGVC15CN2ZOoTTHXFrGs5SKOdPtivkhxDvj1Ct
7kCAtd/BogjSt4O3NW9emzNM0IW3ydQPqlDyGZyvHD/Of3eM+oWTugVLB64qDJcHJyZ4udtv0pmc
drEznQggvfm0Y6/SzJud7zTLuf4Gozo4CWrcyunpfh2/lkDg6YyL6BX3sxg/tuyrRSUNurL90t44
YpB9a6LFnqnz4n24toX2pNoEs1NqaEw0yJvIjf7B1I9rJ8AMojAf2q8Rh36aRYt1FSuarjIcxHgO
HEWNhlpSzMKiBzHRJXEk2z+AhggUuBf2m1GXPgCr4eLvWs/UJnokuE8+bLjzWUXX+IlCv4DtEWpt
iRToc/Kn8rqFz8mVu4fVIPvsqOq3AE/wCFwpCTvU1Y7r8a7Mq+AekoQ/EGLSUlZvMnZbi+1Ch57G
ks4zW0QGe4TMiKYlwxtz20sfLZM1p2654r52vmNaTItdk5uUuuf2XFl7xAJM2Nd5tQg57F/41W/+
ZmlvBjU2WxQTxD5Il6UaWKAGEDucjOtV7+AOnoDJger4U92phB0H2ORsyo6SCo92BJAS34NjNTas
6CCWRdXa6KgYTYKbWm7b9ZPvci1YIT2cdS6wcho0hq7RdS0sBMCANyv6CvOtoNdLHLz0Wg7PoiYf
+mYIbTxpaZon/8vD1g+8p7IGEGoRXU9fdsedSaSWuWZuOQtkxlHk5oK3WxMY7y1N2vJWxgra9zWp
sifeufBXinZyTbB3vaEqBsdiPsA0gxUD3qqgR34mIA2C2nZdE5HOMpaK+vVI+qDNKQ8MqkuTf6hq
RW9TeJ4w3TAn5mQ9tvf22oYjYtOLAy5wJxO/4ExWbh7xvYfWIFjeJKpjUvlIsrP2gQGo5nHjXVJC
SQ7yFxEspJWKOH1k1qfUAMUvIDg4VAUxld3AgQnOQUo2ubwkmoTpSLgM/aakvw1jxP/ziJiwVaCM
rKCvtVgPpD5F26SnWSDTvYLYB9iqiI1ORNhXfPhOKh2ur3BvVvWPeVjCSPUqTYrtLXnoN1bB+myL
RaRzCbOrGKEByBqgEUWlsBzHvTmB1ctwoACnUMN9DnbLVO00mI4MFSshl9VdvlH0JidFTzdK51Ar
Y6Ng47G3QByv2MrTlxipcR97P6qrmKmvVRl9UhZV+32bP6w7iKPwCLBp9KLnsc7FstFIZXfOy1ky
ldMFdU7LaRcxmkImUXjO3NEzgp7SNP4+DrZRTiVG0SowCzszcsFEdTuf0/XYNhDRoZAOG0ue2L3H
HwANOMBIg/PT7D+MVbGTApYPp1lzi/u7TBwRInq0jdBVvJEv8UcU8P5lbiw2id0SytD+R4CRqgA8
H2MLNmZ+iJxQVSPFNUUcCt1gVuIxesbdii9Ys7dfKVjKjAAtHk9yfGqNNrP2c60ESvCvp8dSFxxU
PNFjvcZ7epiOgp1jqN1d7HI9yK5cQqwfcZFTtxDpdIUNd6QMn1E5jZWYaXou2q5LzPU67j1Di2s4
/mqdrDK1Tvd7zyNK4ORoT1YjB2xmCKDEq/Oz/l45OOqzCx4UfNNiyrDH7zlR1TjmSFOZtb+yzbSG
3DN9/i3PgoOUn+QYQcBa8oMS6phLaMEliiVTfNWCCyZOwNt875yWwS3AII5O5q/i2LwIMRq2DTCb
DzNSBLBFwQwTiTPtYR0sLh4JNCQNjOPnlSZCBlUhm0qIAwrlBXuhR7G5UUWdWNOHvHMx8a2FHqyh
o2af0ad24FX4IFCA/FLxvdSVgv1PCUD3YjxPePSatciLKUQOgYxodiuzSivZrDk5LCoUvnYqeean
JzmobJ1+HfNDvuHqY8GGNfRG+cxI3OmBYoy25WTWSgK1olMOWNMJW4/YLBP3HDFwC1ruob2lj7kB
PSTz19EFQXfR2311uMy5bUaj51SMPfch7HAmHi1FbtWnxlht65+kZCbjN1HqjTZSXDWTPvYRi70m
7tCwwuF3ggz0VQNzM4/k0jdITvAIaLrkTdk6Ab+y9wds14FH7VQ2oIEM6ZWw8lAkkXs8EBIHIuk+
MbIwSCCofNICusdoAPdLj1RQ25jX4Ss9e15da7Eh5FjR5X2rica++j2XFnXNgM163p1C8t+YjPb7
t85i/uDQwicDpUQVEk3RmK5MUj8EvwsjbGWbL23TPruSK+8wer0ecPBRDQpcdntdi881ji+M4eq0
Sf6sTeL2tzCMJdVIJEdnozxyFS3vB2T/rGIUXokHN+kwkTwYbYmJizxS3rMbyZsCZmQ6Oc6deluA
V0etjtE6amRMZ2Q9SOSPpUKNvPK3faUxKCSFOEajPYdxj9Dz8J1x5ptwGsJzfuoAl+8gtyNyrd02
8EqeTvGYFoD/ciqGu03R2YBkTwrikGdfjCrlwjjWoq4wT9uAkDr6p71o6js/pT2uX77wjCwVcKol
29eaSWHspjJufM2Sig7364bkXNnReV87mjJKbi/iqqZYejHpZ+96hBYUbCVuBBsibQl8mwsHs0Et
VG7L188VSUG9Tocgxt88bKDd8Ga7e8xIx0H7HQWy+vNh/w1AgLMMm4onx/oZMI2EspsPKZAQBUVs
Ei+Qmk7m1Yz2+t4jQpXHXAlryGxC9r8EzB1uuon31ZwolCl1WloDDqqOxBq/PMn2rBAsIJdemNtn
i9WzD0JGo8Tg6WPXnrHssHmDYmrch06g0gsmKzcaJQ6MQgXZrEjjPXN7tHgzGR9oi3Vlc226SlIy
TUClI+5dV3NVlGVP77YW8ZF4jgpaSC+mjj9KABXU4k3p72wVn0fvgZC2HJVOOeqc4zgLxHgOrXyt
PrtCXmDICRgZBeHzS9hlIuCR4xU0MIcoizC4hwRoiX4xK/xschynq8oqozk7fruAhpClKvt6EUMt
cIm8eCoBVwi3vaL20ALeslKrQtH60elohMX2Wdpjf4XEaxukianl0iKB05vrMd369s20aImNqS/6
jhl9zEXlUgTe+bI7FcwOtzB5XyXxXy+/URrOsZpb2HmSmatIQjQ4SMmPSqDI8lhDcitgg+Vppnnb
ipoXutjxMUVRyJKTT0+JXQTVCWVQnuftEZMkd1/dqk5Omcg1TAqr5F5WUfvNyLTE81bsRP9bvd8b
mKJdG+bHvO0rYkeCj7a0ApeM+Vrl3ZgUJ+xhr3Qo9nkd3zhx7NVJccmcNuVwEIk8KYYz8/jgf6oo
x8xwBB2WQyjJ+paiv0VNxmrbPtFPW0VNFuOL+SwJZbbj0sZVZ3Lu/LVb7ip/C8ril/tiTP4FgbTF
ko4E5KLy35NEH3TXVaVE1eHfaRVuE63mmoYbngmGSl0TNXxKp7sQfLfHqDEdfJml/sjvfVVvyogf
GKWgvavVScxAULTDKp0hWYzY4l7M5fp2PYdY3zy9sCW0k7Yoaldul9kdCu7LW3uap0I4rkOxklN8
12CfTg2bpVGEwIs+LHG02DQbFGOjlrwNsN3pBCTddWv0ExtCS5J4U8iXIJ/Uaf/D0q8UPfBkyXkF
ueGee4ePR5zizrnyyNDMAX8LWd6Q6NBSI4u78PNngRRS1TSdkA7AnEb3TPvID4OlGw4IAH5qI4hc
+dmA0+benBR+P0yWGiys6+JigYFvgkujjNhA+8Awm89TGG/Nbg3XUf2VSuY6L4q0KLDdyuBDK8K3
ixj8yQDwUVyPJMLDyFDOs/8ParQZ012K+ER3QLZJmjH96L0LK1PRJ3UixZ3IgZBV0+B2tz6Qp1HF
eO34wsrQ68V3GCQPuae/mgRFwL0H6uBYkgc9ttaOitHWFQHpJRNQtIWax2e2mP3KVyRJNFSiVgki
o6gNfDcLrv5/RJLLjVkZghBMHlE1iHlyw6+EtBPwe1TwFyPtgFKsJmiK/p0wXw49O5NHm1FJ3s5o
zSAlk2c5kEyLvgaxeWqdrKw8KEC9Ezd26lj5cWdXMi3KS7EAidvTakt++TP/gSwhTMe7MG9OaE19
wBBxVF4Ck6fmnZuMJ++k5g3lYljK6HWK92Fv+K2aJKTtayW01FSvcQFDxiN2TfOCsVU4aWT3vmIF
0q0OK9HmC133Ab5Gbjopl17v0nklXja43b3mLJiHC8GDwt1/BIdP+fzkr2ADnbxHegSH/Nr7gNhh
yruFfC3xH47WOMOgSJKWDCfn6ZYYtR69Wsvs4VrshzK70Owe2rUUaVwzLdsjfPg1JDGNy6xCmVPW
b71i84yGroJuX+4OzJuSfiTn7K+3EYYJ6MSYcX4UBPajKXfl5BIht1V2BjA1DiaIZaoaLX409A+n
JRt9ztQzbkpX2C6lD017Gk31nuHv6t6AgX8P3yMRVmb0Nvi35oZES4pzyOxTWCAT0KjW2anXnbhK
p0ja8l/XBoYudUC2vVxUQTyMhw1qJIxavPPnD7+tPK7WevcQ6tZrm57qtZzHDu0dx5lpp232G4fC
iW77K/n4uOJ7rj5PqHQX2tWcFGCNeWYB/L8OQm/DQwsShhuzoeA09GN//J+BeQgNQyMG4Hs8wZCu
E2w2TwidwjEXxRY9QL9mWwTxIw8nX0m8Th+IHIRb/opdyU60sRAHYX4nEGgxcRo0S5tE0dTzQLfb
fmvPi4kxcsh7cuylH023bQFEOr/9jJPAgwuGmgIU9flw3V/yfLapNa/o1FEchm2ri69pUdOXyMAi
4anH/lwKX76FJqs6pRQdqCQSi8lw96yjO/HNu6yqmct4WFIjSvBqA0FZM+8oXryATRn4+R51iabf
CggeOXOKNc9wgRkMXiQ60IrRcN5DE6+5efxJ8dtDh3hYONjOD3sq03Umla/QC1xJfrfAO5jMkG20
lSBrd4Oz/rbt+KNUDTW3CVn6GsGa0xwPPPNgOt3FBxEhG2fkv8N3pvmnfxax3cbVuSqxU+M1XY2h
aErmP5Jn9wdsCUGhmeikF2RFcb+KSEvNakmB6N1BHarcooAF6eb9J86FYkjPBAROnWh0T2PbBuLX
A0TceuJVD+40DwYW43FG3f5lqfRgAeqQ65mxrie5hn8fX7YdHZSYyGgWo4Jix2bgs7x5kJibF2Tx
8GqmnsW5qICOK0ZAwOgC35pOSyr77cdEtcIcm5GLV+4bBWbvThKPfWfcEcY0DYoVez69+saA+KED
4EHvkg7Gj+Sph66UIvKtXOpPkzDmSCkHztPWeNiI+7xjmfcM+HVVHj/FQSK/fnUe5HoEDzQIUGls
VsZqtfA4Qzi7F2kMqYYyiFrotGUVOxpbG8Hrh86wI7am+wpn3xRJIDUJELGaO6310k4MEumGkdp0
ay0IPOxHDljAwzezw+s9KuJleEhdAcotzlOGZTsFw6a3CaXVwn4+jW68BymtKqSfAUjJA9Cr/cgG
C43PdR11QzmxGiCiUOCN+53j4UlD4U2KDjIQ5NGo8gF523sWmjG5ocqVtD9nmP8f4zecIRUM3rA6
MXEdzbEGTo56Ez9Rpb423xtqsWnaGp6vh2nzM/lRoxcXAQzFG2EENm2PU+HvI6bXpcxJYu3P6N1e
thhmVlEii890QAbQUR0PM41ElJDKa/k5ctEJnNmO8AqxBBNh04/2xhinck+m4oOFDf8pKmwh6Urm
Xhtu5aNH5GJy2XHtbHu7l5vJjGgVvaPhfU4pGNaTtV51+O8ESkc0IpzHlGpsMaBLsDQKOiRTtNSN
CUWRkh2vdqcOPVU9HZdU5bWUzhFy9I2ylc7ceW/dyLsN/8OEYmOs5Vvdfh8/D5yY3+fJj7R7opu8
976bnOZUF3XwBWAi66wyDHMl0tjWdTVu7spamqegrKK5mtqMMpFeofILLCOXmYEfPG040d15XWFd
XGzbvpWxabSfK785D81mgST+MUvtS/Mu6KcG1EN3uIJFs9zSok52Vs9Wnzmgv9MvGfj4yH5qzpCA
7s4ibQPWPoqxz0GvmzoIy4APvLhtIDRmJG8aOiZwAeG2swnEGvO+Q3gg1qqVMMi6hFOm2CEx60QX
h9wFFrO6yewXyiSx1o4OTzAwK2cSoLGq9/7gaB6Ip6i/3erL0CCtE5xmAk0eAGy3O/eUULPjQ9Vi
ZlbE6vT16D2cyGWXylgsrYvqU2Gt8W7NoK9a09WyETeUq22CjmOdnE1aUF4EMhC7iPFp0HcFCA2J
mr74oHvcxPedikfgZpnqX3zLBBj4jH4K7hscWvLPaDznm6rEFNgauYjo5o4S1I99V26QoXHn0M3G
pNrfRZHV645TkrcArbXf0U5g4S2B+YNJLUaXGIUuDtIboEyE6/2ah09eZcvQjKwmPF2NfOXrSC1G
mm2XOT83r6RKsCiKoQYJML5cDrsdFaUClkC6tzTOjpmYMsgwvvOvc2Sld2dsTIIk4eCkf2sS7KnV
C39MN9yyTQcRbRKFncS6KIGh4VFjSYNu3x1Q+23NnatVoNQmVnZTnkqekqAlJ1r1u4wO/8Q14fvX
pe8HmATnkLifpN4gcgEmB4tt4YuvK4buxXanmXBPM4C2FJ95w/K7JWWfs7BDwcVJC3iDbXDCB+Lz
qOlgzH7NEQ/1sBcNSuEIzCnfZ/SvI19pCXBx3htITGt5UTDDsol9CneWULKr1+cKliNUCLncba2d
H0hZZdiujh7V8LH3qv0IFhmAiD4bbiUIf9gFgLBEzYAQlQhvbii1NuIrRcpi4KzLwISbzmLHPi+T
LnT7yVgIh+OkE90zs9FQSMy4Rr1J5bAlTlHQHnlqStJZ2L1/SKZRVJlkx2DinJOcnXdjqhhmSK0H
vlnflmzSJiblyAwll5BZXO3Bhndg9zHngyqUpowbo6MGzqIFbXzVVekuQObCsr3udbLu9XyWEiqW
Zr4UaMz6Gwf/xReAvN9zyQ6wnW9zVfypr2dwIYC0ohpIxzm+SgBDvBTvxR9oEStIVIl87DHvZ73G
3pUaEVtPSjNg5zmMyt8XHLfoXE5H45/vXmCgBQTuPXYzFnX/FOzGHMVtrKc0sie6WeQ39iD5s1Jh
jhJH6bNxdp3zMRybCMYyuDMIKudelKEdBGlMMtQ5IQr/Z62lSGDKTpWrBEikprC3R/29Ch8f1xzd
rH+sgv5zjmQTm5Zy4GpS+xnMidOBqcloGq8xNiUNz4+WmlpFzCZHTwfkUJZtJ0b98gQFKoZU0aO0
L3n+X+5z3jIu6R5t44Zt6zKg2AuY2g3y4Maxd6fgdKAxF2E5dpcBxIdk7HsRvclqjkh0N7cfknj9
1/7nrQLptD9eN9KxD9pvURR0SVmFTCbYRlZKlF5itndQkmJRYp/lOlOEAdfxMt0UhAepV7kipO1n
bZh56zP6rASSMpbG8hodkI78HQISaduFzQQKTpCGjzvxbDm2VhdpbF8gvp2AXCE/s8NTurrXQ6Ja
B+oUJtTWd4UmaafGOILydNip8j4rV5wtkRxyKt9Pyxu5gH6+fRcbdctpwelypOscf6Wgd14xSatQ
bDUm/p4jP8vPtZmqTBxiRfxLiecDMjfIjroM4udqvB/VcBkO1nlcCbpBz/yHv1nlDgUI3NRhzQzY
q4zMy6ECEi3nLxkynJfeii/+N9G8zLPzqOt9j04ceb82yAHQvTVmGtjBVdjUH+H8h9LQUZ1WrKS9
JhFI5vFtc8YaOVR2biW9b4be5iN+NjErcTvG5MmK7FXeYuwmCWG1kdI7bYxSiHH4bEtBVCr44leF
ehD5t+y13rC/Z04iPmgBpgYLsk6N179poZkHzAVSlxwmnTU/0v/GbrCKVB8Hr3blmLatz+VskaRU
oTcEKqSI9f6hQgsXvxnkegJLeLaQukS8jLLHvB21YGY6Au+3yO/nz77xftvkq0ua5Vf5GgJXEsmR
+z2v2iJGS2/CqU3elETXljuVWi16dA4k1AWCQ9HjLDKrtHh9hI3jL9RhU9mLQRmbvKJLagGd+yAc
vzoow7aRCv9bQ4SPut2/HH4C88z84i7U/6Uh5vv/SqBzn6MtvQ8wO4VOnsD4VLts8FKtdvtf8OHi
H5ZRKIj5+eHPx1ZWDr24dyKGg4sKlMCq3YNV1YyXa+rNH1B/ZQTexbH1wIdsugTB267Fha+NKWe7
lkO8cmwz/zLXHkNuRb24S1L0cjV3Ib72LM468R0zOEnP4f/rn+udxc5bqYjff4HJ62FUOPTA67MT
JIc9QaDSTVE38LVFGsUYA115Ke08Xm/q8/81OCwuDrPkg2GXdm/j1w++XJPtbdQwAkliOCidIfqM
TSqZmZR61tVgVnPi5eSNvIshkX4NFdeiuD8xAUlhM9O0ZlcbmcWskW/bZmkRh9sEzphYpO033Vy8
xjFbf2vHT/c/Drw2MyBjZWLbgMwRuMyyZ6HeUAlS8z8YkPCKmxXARFLuOeWH45tk7/qKli2u+fS3
3TL+q4ZZQ7gZECRCyTQpQn/GUd3sPDi6DHS91UpCHSWCDdrrqIX7gOBVyu8EWtZAp5uaEVD1nF/j
BYos+rPRff5arzIakyrnW29GdCNNFfpwU4RPCQVlprNN2Fk21LxPsy2RdXBQ1Pg/a12ytDKHAivx
cHOdkzRB0IA5ek9mMw9NErpFkpprvIHGmtE9qmg6j8VEGEDDZz8eE8pBhdqhXFVCXl0dMAw9IhGt
r4ynfTMsWDAiNCUIx8OYfFd4Tv52wl6jxRBJ9D4P4FMROQ2x9LNnfG4DhvAoZPBWFJya4Z6faqW4
5iLOmc6nPymPCy/ZNElG98TReeRYLj3GeElmpjV0DiokmBHxMnl9mzryQ7P2k78t5shIduFyA3NV
EPHAIhXo/TTdc44WVfIoChTIy1wbuFQO/cARHLod1aIlbcr+FlBfShR08iBf248uMl9nxVgiAncK
/q4/qkhZ7LrCwsOGLU2G5qOC1ziws9kNsru5MseI8YSIE02OfdDISZdsd+2v7mUR4T6/dWk8Acqk
fFPmbHxzQptY7lcJm8OUkCQZvpJOtLG/qkESE0fCivdrcQN+XLrWG92J1HmLXpBJcmZayH7Mr4as
cHPe+QZUbGUiZfdKuQjFhfn03VyqQuSg02O7etG393bB25hkV4Tls0xIB81/+sX1pcJ2E6BqPLTU
UpW2MCjMxOJdxZDZBelGrAbBv4hej67ZI3HAdX+NxmPcPvzhhIDrazXgIX5Nm6z9FAvJl/MYfVTp
BANHlCpGR/rdId9wFq/ZOXYHzsEdFYKiZeVPEboeqO3VOXjMeYp/jOGsP+EcNG7xiOCMOgI4d4kB
idbi1YaJ1UAm4PCbevhSox8tvc8a1k87HKt6ecTBb0L5nQyCKjVQFrd9bh3JEZem1uo17AuT6TD/
qzD4WYkSUwWKcc1s0wkGKvdBRTblnTs6GKZS8Ectm+1IsNO9PHyHUrcjWZWjn1mSluPyZxAJlzgr
buKttSSw+2Mns7GNoIBcL/aRyEFq8yFStaYjdupvslCQ+P1c4nQsxGgES++yN6HnP3ueONTLQfaS
scri1Tdo98d0E8XclCSN1azNOjcGVGDzoSzDR21nMHYbTtlep5ToofSYUBRqRVTVwS8Og/mJ5c0M
h9b8Ansuu3IuPJ6pYUZ2uAkPuzCsagn1AHLncadtJeRZg3m5KhAYDL070F3bhRVCz2OHN/5K7vyX
7cxLTihIMPDQI4HvpwpaXQ1xGN2VKYNNnAATe7ZIlyD2Vgp37TlUUf4BoPN3pkzkkeMrpzJDyIZu
gVYroVZMp2d3ZS9buZpOrcUqZOsnjCkM0eHcsIsh9Ew94c/LPdhYZngOGY2nR3ZV9ba9O2zFSdtP
IByc9B49mW8APwT9pKr6I49paMvW/f2WllPVeUfZEtByU1SsrcpDgGnFtezs7kmWBuwpyQygWb0w
vmUNJVLyFhQlLo0QMh0QbfXCdyMYZOeMPm4GHWf9Z/LNXcNGRgzehEqSugx3xTGlLVsjEK3ngdc/
CgO91tzYT2rhDDtpVESvb8aHg5rxHXeqazZnXgB7/gdCDARt5bdGwCBGa09dMqIDwjmFo3dq0meB
rt6Wkr6Bvpp7ojURP8XQ4C+ZE5EfFXkusQjI0wOWEnYeO8mBw1wIaHdPQKRYJQynGe4NFIUWBgVn
zSVRp6J3z2vsPf2JJiYuNc1MG76XKXzH/ltrSMOZ2bZ35jC4nw8HB+51TZWyXWVx142J2BzZaOLd
tFP+MnhgvExLLvGLDZh4PBIeTJN6J4fvOyMUlI0R4YLJ/OzRnUtYE6+m2tOdhk/W/8Gpc8gQAYHp
Imi+r52DVvo2RRbTci1aVUFxePDDk2pD/3JsFIx7X+66jfRCULpMVQ6923gshX6FI15pbEuRIL8c
t/R21HdoCgCHY0Tp7HPzpVzV4n05qkpUHcg8fJID1Qjw6vMugvAlWtjmMWMPKe7GWoASAZz2IG2m
8pXWDMhG6ZdPLPEOu38yQTKvkX5L2cdcNAUz6sxP94cC6rmWhsuGtYs3HNnAyA0YUdmqyW+V1svr
hYDf2TeOkFVuv3lJjxPmr/whI63VfCcNE9bTpDQJ1wYiUvLD8J6sw6oNY/GvBUUI3RN2bPV/XW+w
mNzvJLl5rLIf/yJj8iS4B8ER2chsgCzPkDNziP0tZkHI3vi3wGOd9JdtYVt2sX/8Zm3ZiLtWDANS
2fQY2v+yGQzXJOg905KHMy29WESHP0mL4Y8Bj6D6etqaPKB5nlEjZDgjCKZ6ye/miS2YxCaku+yr
Bxjp+27WKYn44hfDMdSNTZfK7K89ere+kODjrxiLpo+uBopCxweMoru8x/1Z5COP+fKMe88X2j7s
csJRccwmzrlCMfO/AvHrfNQfc78vgDJmm0fG4YPRG70msF+/xkixLsIZ6hC6At37gp2Qr/St237F
e1SWkQks3JzO61cNbeBvlSkcaNwcyDhMCrzY1Nginl5OvtGsEqCabk7Qmd44So0LHVAZ8T6u80sT
hCvb4uYUQUbbHG9kymhph3H5hgzsQTe/MEzcypZkOIMaAgBRhVszcxTooXX01iIHDTTAxW+f838Q
CYa3qFaBsdqQ17EynNb+U4XdGH5kbFnOU9kDnf/RwKLDM6oMaH5x+YWPhNPGuwYiWja5UOFRErkP
8dzu7ILht7wBOHc1SHY3+ecatOlV+StvzglQtsaYyoHdMGQcSsUzfS69uHviQbkdNnuGtwwI6pxy
VAfPZPVZ9FMCJuGCvNsyS9oPrRTxv7wQujd4pHL/WDCpuhG7qV2YNdhD+eWPpHon3Yv3Fu82dyyX
orxFoMBhcd2AKkgwx3ZfRRBXPHuExCE1oOZwu4yzO13vC+YU6vSom8s8USvBHRXerRnxpI2bxsGo
81MD4d74keVJzlBa+YWHftDyjFiKr/C4SCniFINGH8eIRLmTYXZ+EJxOGXKKfGFHTVr/hRc1vXNC
2MwMythnaJkRkF4hNopZZfhBLut3JtyfqMwWYWe19muqNII1yEYL+rEmoMZlUAFkEHtGqXTHw07s
JItWmAY2YUqQXAp7zODV4AqwDXcWA7gXUzxq9BvAOg9f+YkCBHexNT8DzoFNcRmbzsDyXPwDvPZk
2dEE8sDTPMAdQOtkHSu1iQVJtNkhFBtv//SuJw6TYI5of7ZBjzHEYSaHsC11X1FhbhITphmKbzd9
UdHHBUyyltpwWLx5FwP5rTY9JJhUK5aZMJNTzQbcCNmue2FucegSHgT0j08Y33OtrQ1lyCwJS+/M
aa+2l5N7Ig7WDqO+NqUSlPea2wBQk38cAaM9rEBflMJf3T18Vu4T8ocBRMi6tu42kB/PCDfai5jw
/NiqE8iaPU6UbmsldoRS3YFrHrO+KkU/CoUpLfowxPVa8SUUiZ9TGD5TuCbXXAUH3dZNWToh8VOb
zUVlZxJ2DZVfHxSSb7JoB/oCEut+PHPinA2uId6yfrA3bkQ4A+2YDJ2yF9h+g/34p53CRLGEMkd+
E3b3UROGLEfY/00XlcZLbvf38OeZ+pudv9sl+5zMaulb9eqHSVSKgF2WvDLxobQGoc3+DdYLV3wQ
4sJIu57zqxS67tvpUy2NM1usxdRsPhRGbz6c2DHZstgAE5aMwNKbYZVFvSW6+EkXmjGLo36BNddS
Ug7P9sSiIuKWm9GAxFbFqL1VeUtPoXaHgxHFjQs9iogN7M6tuNWC7JAVY013jjMBh4hLJ6iuFOnM
yZi7harM4RhWMwywmxiw17NJVB+cu/S1zkkBj8NKl74cf9PrmY1VnDfZGk3MFzzpxH9JBGvmz0Nb
1h9QaOBH7oyD5ouY6z7nvtfA8rOttVF9oUb+sFKUC2yqlsyTb8wwsx2uIsZ74RQ49d7cvmJTptMh
w3txjQgwgDkaXF31Chv2lZGG0FX07l2oVGbPZ6KUDbLsukd+PPrzl7F4VufKXD23Hj3kD+2VSdqa
EsalDft1yUK+yhF4/ZeXHhu1KO/XKaEJP8e4n7JFhx1lTTCXVdYizej3NnU+AI0eNJhaQVaTntec
DbvHt3bjCWNBNuEgOGSQXNSCag62BJt7WXLTBlcj1MpI44HCCQa/6b9Btpr7lEcqRhFA1cI6auE3
JRVlQMnZbMfe6oklS4YtiY4bDfNzq0DcBrb3Q5+TDRCYD/xYLfbLFfFT7JDnlhkc2VNodHttCETB
QZkhxD1173gWquO3XM3iuOPIZ9+UC5WafJGWc5Jr9UzVGONJEoSZUL2WVlqq1eNme9Zw64ot+7Vh
PL9/an8okD5dHIb0zTGOQljJZD+LvgPWxBsnLAT78NYgihh6/RKNwpfLGi5Q+rRzSV9iwkM0ZJ/z
es6pd96IL+9BU0cLtD+QuM7O6FVOcxgL3dU0g2if/VxRsNvtj2jpvnvXdBpPjwmnIRUwBN4WT50z
haz3TT2VqKnvGXjC4NgEZou1mi66hTFEsd1Ur+77zKCJOCYYTFF6fUXVkXdvdK45ruzz3QVYbeea
kr1QBIPYZUXyhiIQsOOMrLWbk3/DDTjxqMS2aykisnbOYXp93khofWk8estqpCwSFzZygfjf/dlf
TJTTx4EvXLMPK3Mlcq1IwTjjwjsi8Fx8agBVdwWPp/v3yZ09tiqgzqAuW6PMeT9D4pg19S3cVrhV
a4qP4XYWydGt4knulWVwcOe9UJhdUGxpqQELpxDcofqHywte7X1cF2aPpHRnxuqNQiQoUF+oFnY/
yvdJTzbxfl7h119YIbW7HlfnX+62IYvzG+SXfhU1MksSyJS9nCMeDChUEfTIxwMBw3jyj69ffZiN
voEDvBDo4PfdDEC0XWgQwEo6UwOV7aeRGeN3+fXWdrft2DwgeQul2fDhopYTKYcC2vln6+KxGWkB
2wu3EkVWXFpFu2lK5mve5Ilq7KidO4Yn4yLC/PaO2r9ZJoB1vAexpt7sLGDOfYpLsdY7qqLzCoIe
17lL2MtucUZB5sQLxUgIi1aBWNVfTzDhblG2mVVm5O6o3ThFMl5myY9pHWrU8F+m69SSoGQ3J3Qs
tX69EcDcbTJYzdGPaP6CwYqwtbim1MRxeqFiOa8j0kBSExCfey4VPtK2+ZNJMVRkWe+22QNPn7a4
ly8+fL9ORLzM7sYAS714Yw3sb5yz0hpE7ZkROXwVtTelM9aJUvH5SYoyk79i+s1NrdOMfmbPZGt5
Ec5uij5RjKZ5qV8XGuOOlELtAuEttHCnSGElc6KQ0uR9CXmsxZOvdpapQLagBlKTMnpwE/xEnprQ
L6V3/AVc6E5l+0RZiHGeqckuJHiH7M0nhwc5OD8EeVuStRy8687A/UTzmMGFrcJjEMOtccR37MHQ
r3fPKNhgFMScQmW0By2Ki1ljxlvHelgqz5YaJGQXK5baRD7RtwWaI99bbuNt0II+2YnBYtEFLLYz
yij+qADSa7wRgEucQwV31Zh+IhL1GiNACr6G99YSIocSVrxG3bK1IB0MIcLIRF+6Hi5SxFUGDrzC
5HtwRSv7LNNbf/JJCFAae0z3h/9KiF5c/rspvt0zxXq+GtYKazLe+ZslqRExFr2JLK3wFYsCxPMm
n3jW7sFqXBL2Gm8zvxyIvClLdLOW2EQjJbUz1goX4Znwyo2eUGBcxHWrU1yElVdCqFpohiWYuwZ7
UX/pWqPOaZ+zcsVcqrq1kZ4/KjzpoglnH2a/wvO/2sWmLAnfWIOSXNtn+MjxmQSMdeH1NY7yrxnC
CVRnFZLcDiJJdRc9Ou1orVcmO1kee6uwYdVUAoRoeLnDkwaH31JutaAazR6CahVhu5f7+p2TEztW
3gv0ld09Iewvp/IfrT9WrcqEVslEyJkoi867L9w77h4y7ccGavJL6Wn+4NOOBc8x+oIvBNKcgc7N
XWjgy09JoHLJ90Xwj04d/dIfbbZbb0GLDU1DhMJ+KMBW447dRYV0KZUZ02gMWkc9nLce2sXvTgEs
Fhu6Qr0QHTqQtPx24IprZe01wSUkFDrd4fsjT7cHb3CPFHPAUGHWAE6xdv7l9lHYC4bcmziXuER4
YZiPgPPzYsA9l3jFL88RhZYr6M6RUZnZlw23dIwPGvx0v+5VcRAajNZ2zA9MLige5jeiC1x5aUCc
KQlwByeT0hQvau3aykcJfYmvCH/GcBt+Fo9a7oEOnD7LNq6H/FCcnme8rDjgJbr/+khAHd6JOXE1
ePrHDb3L3+R5pjOYsZPVptYG4sv3KlAfauF5f+43HnSk62hjAzLYqmKW0zK9xYqJeu4f7mfQcPCZ
yGpaSKVD75E1jw8EAMxJN+/eOeutCPvSE4yXfRaiKEqqoJ3kVoROFuzc+Seflimh23vidlFGSUP5
mw95DbUtzYRcCk1UU8RseRmf9oee/kUwdMTOPLCU9+a875CtB3nDkvkAageqVt7nnKGHmFU3oiWv
aPJlOAF4Va0c4Imp6wenc00z9M5fIyrJIwDulvDiALjn2jWrjDAIICuI+rVBIVH6umE8owK6aRkn
fSrHOYvtOP0YaYdMFeySWc2tCeGkXH27dCEx2I7XpeKzEbplSlJuyIkfMd6bmey3voiYSR5U9aNk
q+BoNnAnTO+oBHijvhzx1truRVOt/d8TNGVg3jmBaVQJMV2/9FxX64AJFIOmwzTuilqeSnla7twC
iXlJdTVhhVz9z4dHckwBjvqTwcxu4XLlZahOUe/7fDa7ytdqT1K6kFWU4QU3ELX1bxTxMzcf2yQb
iGRBObZdabj79AsY37oujTNoiG3roV4Q7EV/OnogWy3BDcPgC+f67HQYrMOuTBmkXPbTzlNpBzig
cfG9j7gy6WK6E++DzV74MQHlUFs72gt89yrGL6AynO0HToIgfc3pE+aiYeHbp4Q7luOot7aQJMVs
AxuzyaIe9SYLe8utJVgOwMX81Bt7w7AqLVJ4/Hd8HzfhTHemKfzkLnyvwiHTvd7v/MI161ipFrji
JaZZQtjMa8Hf4tPg0UDcmWB+SpoYP2DsU+giCzh1O/Z/UQBnCeoEwShdyQUHHZ6YN8iYmLVJEJ27
sfmB1lGoRJeThTp4WxsPrQJ5+mxljY6vizul68gsjef6150+1WfGDQNAdILKjDJcDNq5Fv6pMg2q
XL7Fejnp29MH8BVQ+q3vtekI70a3XmxKNaE42Ykg0QO7bzhyDQzd7giW1QVhe/O0DUhlFzmKbK68
JSUPIeLFU3rZe0HKKbgOAS9pyFErg3zQIACHpWUwX+ifCEcCf7yoVheMAUW9EHrZDEir4c/Ik23Z
oj02ZTKyEUCRIsfV7hRATaXcCFCVKkRaZpTPNo1EAMnIcOehVxBKrqt4SawiBQwP7nsRpDp8yjVU
Ge/Vfb8eeosB8/HWPrSNXb36cSbZ3z/rN5ozi9VTUkTU8DZ2W2vRHOuYwIbFVNOWLy+El7h9HgvJ
sG7SvwzpoC2qsOJ+U8vl239kTvzJlep4XWL5izATkWNdxkKB1+52L4vUbQC0aa7AFHct9nWvNfV+
rQAWAPn+XODUiOMW8iSPq8qUiABZj7GAavRCp26+xRANV6lwsCwq/xilSf8Tsp/s7qqXn+03DyRD
y83sicIPWneFsasXyR3XfofDryWcO9JkhTHLH9Mlq6cZiqriGcQT+63bh2+Hz93R0kDB0RyLRRbY
V4a+wOZAkEvg838jS2DFiOOLzAsbkCzg9NacpR1hHP22lmbjHbl8Z9+I7uC7G9sELU7SUl29hzM3
Po890peG3GSg8FGfhmQ1tneb9AjTDFDPIFaATdd75MVJ/i8B4JahK8ToYa8MqRNW6MK4TrLYXpVZ
xvfdnoHCkKPaWfPDLGkrsK8IF2jbOHWgBGzuaALdc3YKNCM5YD5LOMyNeMuj0cobUmhGStb44SUS
B0tmJFOT8mxKKA9tBDBUnlj0qiXrMaHF+Y6/QfeX8mGekd/cL0UjLCjmI1tuOy3TDWsCmq1ic0pZ
jH5P8+HVdSbCByldisdIRpZXmKacgIHHYZzuYZDTsM4v96gLVFMF8Z/NQ+Syp4oD3KamcbHCJVWx
c4DUekruuy/CFyrSoV1IFw8CAwsJ4xSKScM+dFAlnUBsbxTwY0Pi+/dPcMPYWHwDY9Y7G4vWaPM/
eNgSQflJp38fgIU1NayCD7kEOPRqTznnDn9ixoaxolek7WlqDmA8J8r9LwZSvboEk1v9F3TUHiCy
ZT9mphGyQpnOlmrmJDSlzfxNNTgOYcT9miPl1SP2ULP+8PzcZTtOdRQIIZCiVtOJeKsI0JGP2CqN
z3jm06SB5N+56FaU84JJNvi/iG/wDGiLiBvzVXH907VyGo6Nf3RSBxdgqqnHgg924a1psBynIr6C
C2qZjF0MMRwdC7d1QfYdhD+8+8sXHGLXsDPFr0yMfwwCZrLNb14U4KMM2Nupn97pb0yhVh8pzPk0
vrcoHmESJbDp9FoZNYOTh25SmmXqDctVcUI0piWXhdaxx0BabB5eC/l2oFXtaBhVoYG0+hLgY1lj
+CdPlFryALKHizFJENNxUdLkuaG7gDJjsCU+p8JiUaqPoqokl20QDVCm5mtQ33CZ0jat3bDqBokO
z9WZJL2g7reCXOgxr4fRhsRILnNTF66xwoKMvv9Zl2SJEOKJur3qHc3niyoC53qiF695CzNtZEHE
4etdgXm4DZDmec67gvsyBc/KttlAMWElXuO1zZiRRAHVVlPPl/7H0a87qOa3Hn0bn2NwI3p6uGDY
/l3gnCG1AnaiwDG/9bfB7eRBM90qokPkZHGLf4nC8v2ktk2OqeNi9A5RIRkEcQhK9vgGmQ4USnTa
+zN8sr+D7qUNKteSH4MKcNhsy02ybFX/kVVkhPD9LsCES4AYPyo5RDQ1JVHISsUeTRESGctW1Zaz
aXALo2SCq7jteP2n4IVCO8I9aiNH6V5QnVpFT01aeUuRn1PvVAGHIkrDuERDAKLzC9fUNV7kBKO4
Lo3AoEO5ZMceNtCq3eD44W/Zee1RhG1gurT5kJtlq8g2y1ZqHkBIKV2eQi424EWlAdHbBWkqheta
c7748R45Ak3Wm9Z7JEJZZvAzcG4U4WOvzKgW/4ZdqKbsTDEBAXQmUI7W6t2xUeTSVkHhCjie28wg
JbTB6y7loU3S62CR0SQa02+137WaLG+sYZlDRb37urre95aeIvYr/gaXZS3Z+Wj2pFN4XKQsziC9
V4EgOtL6ByaxHbKqjGsYPBD+GFkq09hp6U/BOLgJimpHmTqpqiAkYgb7gWzPsA9vrqjX4Lw6sAZA
7nOsdhFH3YlEInaYPoY4pDLWedAF+frN46H8kndN/nFxAsqJ59F7Z+f0v5x7FWMuex4a0DL/CUWn
sag0LWqfhvwblax+/j5n8Fit9n6qwiQmMPjxlwelY2bTTtgIOToIkwlbnsxC8hx05FHYP6Fx3RWK
Y/9ptZONGySPzXI4HKB7DxL4CqPpEgT4VElGEeY1Iea8eJCz8/Q5FEsLG66Q3xqNwMSfBLrG4wDD
wfvsiMzhHT+Te3mbhA7IlH+hZq4eicu4FBPUvnaVi7ZsMuM2xSF/qtYUfNS55YCtpJmSQZTYpCBf
oQjcA6z2w6OE4QV6BHelU4MW8AMv+uaUhywonotW6ZKKkZexR27gVePnZYe3ZZtBFvYNCURpn+7t
UygRMdVuR5GNd0iYB34hoAfcCQkrklEvWVCk/dCLZT5n1a2seOOvMUir9CDVisc8EjVwx3pMrqmW
IpSezCiWY35SaTQccsph5JzzETsIjb/8kh7d4bEcPMkiIJttiYLwwuwUNaj+WZkXaB70U1R+5LZp
nixPSHfj5Lt2B+ZM96kV+a3s+4hMzTPftn9UdMhh5ZKvXMOoIvOI6UD0HT41dg1uLk167fPyDM0z
D+b7yNQOmN54p30sa+o0g7b/Dr4YrKxL/wTnCLEkjhiy3CfY/AToM1BZYiJgKPj43wDXSL+/ILQ+
bpv8Tc+k+EZ2HMpc7cGCi5gdx8NvHlYbHZE+dYuO7PJbDdf7hoj15M/CdUPS2yH/I35O0PCTHOGY
qSiGD4bDjfRYBYdeTnbw2hQUHNKRotnp7Y/dQxSOWWJgqDfBEpO4P7A2EQdNEP2XNV9STuyjPPTe
yHZkZX9FAMHb2y6MsdveQU+IIwvQodw1R/7VJJ22DSwa/Q1W/CBlk7jt8OFmle+mWMez3Ub/B771
9eIZp95ikL2DbFzEpoRbjJujdDhSeRML1XFGfH9kzG9hWT+2ofa3iyiBg3q22Pa7IepGhQ/M/gau
xTc1kcZ62g0Hd8yHR9LM1kiqknB3TxlfYr9nZ/BFmrXYkuEKbDv+keFYup6KFJ575r22oTRiLWju
G2Ak9qvjdpklKMZzemO8R372D6kCYIhmtAV+iF1cHystT/Ue91Mw93jLopgc4LxqZ9Llr8S4aE50
7P/E1nAcjVF10AU/6EJcfiqvty5UdDoD6dCISeHdk+IyfsN/5koE3cqV6mIfdKfT30FtVjMJVHCX
nX0AzBqCnSUkiyprlM4NNuFcyOSAt/m97ES2mL82Ol8KcoCMfhfmmPAWZIa7PPjdfEGMm3hdIOmI
aERvB13Ekj/9wDZhqFtJpqitA2/ySdt1dXf/DXAQN0y0szopYS6NssqUHNOuWDeALKxWnImSnloG
eDNjO7uz+O4z14zHB4T7K+xePl1RjQgfEp603T+nxkiUivLnQhkGTwgWQywimjoR7+Eqr64cIRHc
E150hzzfFu/9jjeM53ZLIsC/Yyuv7Pi7H4APtGfzxstYUKqVpv/LTUXiAfAnuD6e1ktscX6endcD
XHZJhvTgiwXdRE8X2x7V7xQ06xGcm/XiQ+2duFMni7cYbXJLGGGqV/Z+czOWQvvRfcH97O2A2Wru
WCfVz9xWhZcoloje13/9YrTuJ0GNDRiD44QKYQpfjopmj+KRsYiPeri1brjYJN92wHJnPqZ3WCel
GfAhKWqbE1ihZMgI2+Ze4Q1QgiV0fj0JC+gGStIKN+unCr7Urb/S248z66ChBDB/z3xWEeFRVmgr
iPnpF0NXGn21lg4DxZyO7rKOrsgCm8rFDZzpHGjH9zJMNtX5+0vI/UZUAKiv8YCrDj5hUVXDGyJC
KY0zB3NOlXPU0S7qBLc8iqPyf56knwoDnvWWVhD6D6o+Q+pv/pYyZC6dUGu+Z21JbwR1ipcOTuHf
lP8+euAyOgr+VzRCrSUg0E5GHNjztZsvVp6d3B9KSY3hFj41Sza/V6+MpDNDKMUWTfPudKeHHcy+
/ct38slMFaAa/BE9sxIxN8AQO28wmMbGa1V42pXU4sUIQdCapXWnSBuno2Da0xnnocT8kKHNfAat
npochiot5aHxXLXO74YA+ra6BELqsu8nn8KTFO5FAGdpolhWdMf5AgHoHsrTMSjQ63wLM83Nmd+n
aYLug5xzlGjBWIm0oLpm93c61qi9j/+qhugSESmfMMUeafGYDGOBS8j9BCOiBelghDoiqC1fEaoc
pTF6lfkKBGW8sNvntEPEjP8/KMtZKbWZekmgzuOji+kkQA7Wvh7PIV6rYw5j74i6NKB6fZ1w4MaU
sptHaOdS1ryn1l2N3mdFpPCOR3Fa7gfo6EfFb9/yS7Es8ykP2kiWEg3UXGumMVdPQEOseJ7z4Afq
WYEzv8xi0Q+V2cUmkOeiyA6b+9iB6re7uVsGj38wFD4IdGQEAfep0k3x8QMbHC+VaVv9qbI5vAIy
8X1TBaivKiurovahXLNsgMel2o6lR7VyLQLghvyxiVbwIashhv2jnvZ2F3Ns7uSRsAIezFSrlX1K
38QdwOPk9VXhxr+fQVKQDU6ts4ImgNmcD9AVhft/OOnIan7wGm/cQAvVpyRNmskimpvi4lA7KLDp
IdqAs9Blx9rpiU3Fi4XUq+MkQleUZ5BoZ7O1Ona96nhj1qJsTGfCmikib3z1BxPO6ElGfWNWQf49
VvRtO+lcu/MQEj84aqLLQGGv9VV1TBOm0sgduxiu2VU0Q3uwjpBIVlJvVoLu2WE3GyUwroZrdnbM
u/1ynUy8zu88oU5IbvdjUVuTtyZ1YcAWQiYouuKmuSOFD8I9mpAhMAIAIXsKH6XM4KfYy6d3OhXq
eaPdQvgfhi2OAFypQHYqrna7Sc1KUFaCltMoKlnSbR1HsafB5mO+xYV1k5ZG/XY5J4JeDAuFuDba
wD01II5Epm1U3BIPEF57W9DlQwYLgrW8/YBjQQmNCvzEtXwb2il4MfCnzqWf0I0df63g11r7Bkqo
UM6hW9lUX+r8ZKcYIJ4GshJtCh4v34/QXeRvQw24CS8SaQQYyQOFAXNvTz3XpvR34s0r1oKBPAFu
Y2qdsyM9xtw6ZkxCO4fo9G1GvOwPjF5WESqy5V4gxrqRArmlroV4L3R56Utac0i2+sEwfBNZOlpO
0TdNefzxNQF9yaM+OH9Kzt+vYoBcs8y/ezRKqPAgPdq57jyn66SFWfrNh6aSUx9/8SF8GP9Er7J0
V2z3I77LzR8C9oXuRz6vGh/gx4Hi1U749x1pnjFBO1k+xas8p9aFc90EoU1JTncFaqMWcjGv7QB3
PvofDxwNZCV47PGy7Bo+Ma31u1/J2wmklc7vSaiAR8eWog3WWNBO45WGNh8w7iTHMRAxUELOM6rw
qx3DPvUMF1T/KOzybTaPeIb+vObqNuHN7g9fomX4pItNdPuslkJ7A7pC01r0pO1egIcdyc4WM0VG
KrGUwQFfvr+Gog6OImaPN237h3GV932gQ9mak73D6AB3R+M+9t1FrosFrfn1f6JE9lLKFi017SrG
tNiTyCWa4xuD3PheYFtcZdg4rkkwo6MKIf9nGAfVn9Jp3zHDbS7GqqHAMRdmKJr21dlmgvQPeUCb
e6phZl0iXga6aEU8jiQer0aDL7K7QnDN3mV3hZ5glE80xSuw0UvP1fkeDdBQ+aWGzgqaP/U9L+B2
XEufHWDysMjJBeqeDkq4wKEz/LlYP/yfSwgsut85zVH6fsINvW1jTgWuj3B414TjFW6jAG9vJcaA
k/MwU6+6TP+lqhL68VPEws6B/F0dHPHwzg8RrZZu6dsvWFafWDpAXxSB8tgNjBwr/XURYntuZ6e1
JinVGCEnphJTcP+9WIJixaZZ0OOjIynDzTUjXA5p60EPYSnv9xIOTMIoKAnRI86cr9PsYHl1rYBd
bl4ijes0ehZdO58AkofcPwMyC7bDSe+l5IEH4x54GAoOCJylmxmUGjFin2RJfdf1P+BlY3BEBR3m
5fZrWwc3gn1mY3RyTtiktmRSrUDNeWvnIZcLgF8jOtTOr54rzmXo0LZy0/YDwfNGXXaZOJd5TIyc
GLVPjbrXSv9VLFZ7erOHUyZFk0tXDqxVpMIG4TvrvPZzZ+JkzKdeKsPIUb1A1DyJhEW7VhQf2CjR
u7tTtTpQOOC2a41rX9thAu2yITOWuCOLiLM5IOOGLkfZMHHUsHWQIYoXxy4gNLz+vM7b7SeRrqgd
n8C1oeooHh9CepNrur6/A6UZNfl5Y9HflrEFL6Tx91lrHIt7kbyy+CHyKK0A6+nx9quM2vmMx1Pw
eHV6ybdbk29YYZyjkn2VHPwE1yH4yIxGk8WBm9od2HP/deokObCXAfcjxv9VgNSUTKolTJTTBMsj
9OMOV5AGsiCZnR2rTV6ysvPb7F9rHw9bwwQh1XdSPbuxbYzHhIoicvDDARrBhxCSP1ePdncmrk2h
9ENs+nnYPeIuTV/U9cMtg2JhSi26yFu6HLUmq8vYfESa2ZXISmeou/Eu2/P5E2qwl/YrU10C2Dzd
EKkTivSWgXjdruUhkUSosReJoii5ZEaz40+NZ8zxxoH+EDdzI0MS607yKLFhKmM3gNieDqAmkat3
1QHt+PglVy3/Zn+NQSptXuTfdiUeM2B2kFRQ73vGkMU9uf7EJLrAfSeOIUByhDUvU/26aEbtbJkU
q6RFd21GuQq1UinciHpohhxT2U7t2/7/EFBp9seqZU2YRiY2GG4UcSqRQuWA4eYtRahas8gGPmJ9
9ktWntPlKPfiw85zAravqBhBkH1gnMYUo20/HJe0RRqLVaJV0mRYyt01NvrFQjDXpfme5fwvWd3u
Zz9nNvj35d72CjAHpwAIjA++2LJHKjM6SMelqOJwnEZPMV+fTitkqHN6lK4AeIGZ22aeCCqx0Ts/
bEiXmPFFBTHKHkQSQ8dgM5vll06vjCG7eLcgX0E+BudScNGm6vQ7ezEUHA3YhFXov5AR9VqUwDLB
BmMgb9no9CfMNZrkK1LV2wx+xxpK8m+rME1WTKsxE424Mw31B0JP7tq+yJqhVBSAr59o1maX6kXh
ujg+1X8/BnQmigHqn5P47ymYgfk673w42Su0BkogFjLaA1HbILzJCjMH+mHV/iGhjMaxigyYSalD
dzfl49SXuHyVayrgKKowJ/cIsLyrvecO23Bphukk2bL6cvuhqb/gpZHlIZvW6pYPsFKnUwUiw8RM
M/ji3z2SNedECq9oMOsYUxI0kGsKifSl0uihrMZ1104NY95GAh+Y9MnqEzgeDyX6A5xq0DRrUQ0m
5aPczLgI2SVweNOppSks10zPZRUq+2BRllxO56FNhSun3U45j8ikiFiBfEQZ4M9RjyD4mpTumzn8
aHuimQeUiNOkwZj/GC+oVkWeBiPPU9aGU21yPe79kAUvi3jBOouKGE3JhbVkG6P34Yk/GpmKDphw
Sd5XfUv8hr6hYzNsD6JLRtIrU/1w+tGiS9k8Rt++bduMOLW/NEPWWEGLhmuWyM/sqLKBamvO3bDj
szw8TmufzrerjgkonGgP4be3zs64qhKEiLyj3TJpLdXmafp73ve2eDFQVji2bx/88Ip99McwygJ1
/7o3AYMTtVP19mcVG4oJZcB3/B08diO9nxiNC7KCnHANAfkYb1wWsUBkkslXIJRIK1ypxzrDvrfu
0qKSyLE82wpiMPcYz5Hm0siO7+kSSjGPyzr6EfzhQqXpDEPF+dGizddxOiLKaUPHxn/VMnV3iThF
RVEOcYr/CnLaEOzGBUlYmCgluQLdE6pdYQKMki8xKAMPjKko4aqypfdShGsn1PdFKAzfH/Yzo0ji
qHAbawVUaSOTBcKGRsXujf65TUayFWuJVJKNwLuBeUaci67ZZtN3plSh+4bwKeNqql40lk47k6bD
pNBaQJVmzFV4Qlq5t8zyaUfgZJfnvGFBH43RllDN8WbXhTrDEViptY1h0ZtcuI7RuGfMiVr6lSdo
AtVTx90Z7PKfqe8rEv83AoyBOgj1J+llZLMxjvsxwhXMLysEH0cz2P5ESvCzYu3Zn7v93bLIlYpZ
FXWGgclkfULWv7FlVPwv4DX8QMnOnjxbdYMf4sgnHwXV0mPzXWY8wx6c5H3QzfbJk3+FugsLKFIB
rwynIN4NOP6fAfyzXXJZj1UHu+jiJF8iaHpGfmM6FmP2S/+Wzvnpmu7b2LYnajljeceFZHSKLbTB
wrgRnNHwjS062v3wkP32RhcsNMQ4Io3m8MvYwVlC9AowxeQZtBF9SOXVu/9clr48fAI12VwK5cw2
aU2sZU0unidy3Zhrl6B5uvvoARBKevsgFKeKFWI+PFlvqAo7RYXgPaeyBUs0iQcZF9NepES30Yp8
bZXmaDqiVhLntIfN1aKdHPwAQLzrPG1KpKtQTxerOiXojMK2RSsgbp7sFkGCE/Yf0LbJIEKRb0iU
yAGK+QXfY/ogDznE+/VnepcqB0ksGgbvMuCi3ls34SyfM2LMUMLlgvpVo+XBvY//WKZ4WPELY/18
Jr7zd+SkrImJ/gN9M1VEzCpRTil6IxGiDh0rNZUdfTlsgiNQQ3tASVGcbARu8xmWXbMei8CMDkXt
gRTcjdUqI1xZArM06FwxT1O4SdELMQ7V6PGE9CAwT6QkxJH4U5qkvTiStXIGHC8O5CZsbUIYYm2O
vBl+GYGtprf18/1v1+ZON0wYypcbhPnqccn2O/q7VbWhl19IoXp9ACjuMSYokMnGMmaPe5v3/BIY
hwcbq0y7NQXzOU1k7Wx1LqGGh4uUlIDOTHvmtFjR3Xooh9MkqnnsTzWH2ka1aR8GXmCKVl5+LeGk
YnkvPuQMhlDnYHRNU1xuowFqxwWqaFbwjoapTrq2thlHioaR5C/2BTevIQEc7FR/ok89COZJX+sB
xfG8YiYiyM0BnhJtfWe85fLHoPDbKd6/NhAauiKHd3zkg4FCy8IfoxMPKh/MqQOhR4RVCvbyngWt
Dd0QpYqHPrFV97xmMrgMV6fFkpyTaS1A5ln0q5V6fKUJr/JPpIT3+V9pmWL5dzWjtvwxl8c9UFd5
RMQ3P25SsfgGrtKBGbtvUM3vYbWrU82xTYScokvpz/sLdn5Sy7caYhaZXDihuJGgDW50pjuY0Apv
moAQmlzlZ8s0gzlYAzaCKwYSbVYgaMi7RIU+Lx3DE/T0TsEb6GKAuOUoKas6CBILcYBSJ55sn1JB
c/jRzW18JYZvNnE4KNh6FlY9A4iBHZI8V+erOySFWI4B36FEK97/GOybgZr02d0QUM21BoUoIY/F
YppyXUn4taSbXz96P6Y+RWQCOa1P4N4A7/m4iszkgrxhj5ivhfnFYK4W2WfKG6Cm65aN76dg2+SS
Yn2uJMVJrdBjs+zUvhm4Mdn9k00/DkHcMTUaDMxF84k6YgDhVLWzQwfc7zL5KLqJX0NDZ2niwKNx
9M/hSsTFwdVOoBOO4iKNIbeMdHb2TdlmqqtkGx1cZVazJzzYhnfYe06jQGhugyfXbd3E4hA+yyQv
tk3i0tE8cyKOtv1LZXHidLFF1JquTD8TjBZPLqm0JfqyHmhKeEKRfc3CB4ypYYD3++NfcE9qy8x4
ICdg3typuuPxu1x1xIE+6eMp4ejgtZaoU4qcTIrmpITrM7kkbubten7heMS25Pgr+uWRPmxel+l4
bewZ/XCxh492Vkx7sDCGJUjJoqBmzTT0O9CmMdgukc0HH3I3BoELd1fflaBVaMKCAC9NP/OFgdw5
Ph1Ao3uPnLV/mFY9CJna56WrJexT5j2kM1ZWa7rBIoXSu26LfWaer7NIam5SzGyeMtQ2hdaR+akU
MFXHxQrIZ015U+z0LdyIm6YaSlHwiLWPTBG8dl2tGpe9KbYDKUlMd5bUGew0OV//ts03zpPbI5Ep
+tcVyz1usHRiYBSg4Ab3C6yK6zxwuTL5sBfaMXruJvEI71MzUJmBO9ubUW23qDQOnOkVfb+P5VVc
Ahdbuatv5hADRxaKCzogl7D/KqO0Sw1ul8gyUu5I5cakXmc7sNBjtEvaOUiJurOOXRfE58MBhPKl
eJxXp7Stg63Fkm33scYKhqSdLhBEx1NaJrzGX8x/obv8vc31SrQDOG1A6AjjNE7n/NadGEi5ELQ6
wxoQxxJL/zXPL4QLRDOVR8WybbvWtZj5/QD4h29jLVeXX4otNaDNLgfQshpEVmprgl6yiwNK80P+
7Klj1IP1F0ebVuGSNZiANeKCOCcJYUkJ4m762TvNvcKEfLljRUsK+aLPQQBqN8GX7L77z+QBEll2
VJwJjksVuJspHTLXkJ1XbzDcmkmO+ghjS7Uto0egrlNmEI1ZlTwtrTinPBsRYXSma7zBLAJgVdAT
e1bl/s3rhvw/6mJCvIFLgpiHqqOv3bmjfT0dGcFQtsFqnJalJUr231/6R/SoNkVUQJ600wcXriEh
e6DTkmJ4ZqWM1QU9P3g6EG9b+mvIcBCV9y65bOqlBvTh4RIEUJa4BVN8A1BAnJQYGYZCeYeIENK6
jwn31eTgS3AjAz6HlmRWwRdqYPiRZkJK22wAgu24e8K/346NWSVxltqU5EqauvMZMD5zMMUCSETv
eP5cJLKT0EfmW+ML0j+qmlA2gZ19Cl0DR5Y3NssPwK0oObKZiVQlrJZVlCCZpCtyGdFkHSU5DbG2
Tjyh0KTgiXXlv5devlKYgxC/p3DD0+0I8n2ZYqkRs1o58zJdBzO1opo/eo0e/oyLKekKviC+Ib5a
aJEFx7UqATH6bG2bUZZ9Ijwemz7q0lCgQ+ceytOjqvlp/atgcdR4NpCT/RC/63+u3cvXnG7gn0tZ
QjEYdYIL3o1HUiiwsn4mf583HrJx0mGguWjrrbSemtIafiUUM15bwMfGQtK0FyMMDlfYQXKfcQh5
NNQNM3v4fJTKmDTVoJ8YvOZO6a4iLjsy7iSTvSxlC5RLYg1GHFWfn/pyjJbk47CXvLXdfKWu8zax
2xfDud8OJeN4StB+lGU58XbgxMfCnU5aJEGuGZyGd160mNSFTs4kD+gr56wWYgSQ8Es8+n27wtWZ
z9RQZgXrgieqgGDTNKJHWmA7e6NVFVv/L8gPOLwV/7kZ7e4g1weqHsYy2n+XQPYCBZHrljyCPC4N
1Kb0pBqfoVZsHgBwwWQIPzoJmoAEkL2+T2JyjN/QAAsElwy53Qid/MRvhWCaK62o3sCWNuDflJQC
0g7xj89hpqncbBQ+dfdV6DSwz+Mjr0KsQgYqAyDvBaWaKHW2MGS0rY6JStONPL1Dc6HC7fh6ap9A
Row6dSoReSL2KzfRLQ7ULteyKKmoTDdnr9XRnhpnolIqTqwCh4Y310Winia5Ce5cdETJTBMrADSV
Sr4TO4qF1kEbi85qTB9OW2gPg1rzsq2SIlqUk6scsLPDkJDktGx2wyh5ZzPGU9vq2ehyMo4FDw5M
HF/iG6Jw3XPo4TS10EiUk0tnfWbS9I3wzyuw5RY9rBCDP4ZYBoNVPkyruRT7GG1KVZOsre3gGIkn
ykzSda6nLJG9S8BhlxvCVATJ1tS2IoHAMt6o332RPbYaCRyEnItyNSH2twSioP5Nv79p/PeZ+xqf
8J1bkdMBo5Q5ai9a60m7Bi1/DcFWDCVH2UGVA7d+YEyZLRGg1UOIdvwp9v4XEa4eQ9JTe2+c+GLI
qnevEOyC5LQGZBzwQEe/Z4vKau4ERBTH6uA3A2HAaE+MRXhjI97q9hVIdJDwwZpw3/lZPGp5eD7O
aKCArO1h/OZu0DiYGSAFnln3AB1FACJUgc249q8TSBR37hIaeLPQrg/ISOBjqq4bontlvv4qCpMo
YFzgUjWzihFCM6suNMnlzCCwGkZpiAGGNT0wMjbi/gfOOV3krFRB5Ht23k8b8DkkFbDtDZunDrfy
5zQDlDjJyYVGdb4OmHtwTMUqtLjLl54OxdBB8y/o4F1VxzGMa5IQEpqa8CJrDebfoe5uxLNjaW/+
CwlAgaYsGWXV2b9GsanXFlOk5IoNcRtiVm4vraBk0zOThWdeiATt2dNYgLzNk98RHFYjubJKAOt1
IQUJYtQiaa+4w4ZDnC4275df+PD1GcY6A4hPF1hdOuGsxBDEE9ksEGYDbfC/YphiW3AcSL5VRO/0
AWpyGmwxOvhu5tPcOPjs0nUffusa2VfD/eqhXOQRgVzUgolX+yeSJ9ll0Hf6phdusCSMIhvCoZ2D
okFxS6ccX2IH170c9/1PGd/DM4trFsYg7lyN+XXefTLRgsgbnN1VMomG9YgSs0zWhk6xpO/uv+/y
ms9yQwuGePF+sCv/GTFBpaKqVxJSpjbuqI71oCB2dyfofjUU4zNsD5rLxVbT6+dITF9+PpnDy/Vi
hKtfz9D+FkZRP9qP+Em230ySikHlpjJl0tGH3W6QIl5aRznLpslNbOQUjHG4fGYShqnspVGEkaTX
nU3iawkmbxsvVmraxVxsfSfkIvs5j5RY25IMcbM+SNOvjI4BFdlWLhyZkVr6/ZBoS55XUIftHaT5
/re+X1IMJxJ6dGaFlvCO+j4RyGjBjDcvKix9aapPbs4sfJIylK6rv4G8wlscCDDbCpie8C2TzIO4
is3Nffhb4RANZhE08C9tcWKxMlh2tL5YVhTNs5gzth1vncK5pu4ygE+i7LZ1NeP2YTCxSPkSv53s
awo1v/haQMdt/9Ia1sZ2HJORSYyd+2b3ds3rA14QsQIVot0ySsJqGAiY22QTqubXGtirBEr0IVlp
JwsFrKyb1pGP6fOgip/hal6oAu5FwhUzkeSsycOmBHYgHxFKeFczsS+duXsRZyXU8KXhvnH0QJB1
KHiXh8ausb5FfpscB8/gizTjJXlX6aDBR3DS980OxD6WK/tLeTT5NWxLdlyrY4dZRIP2wou29sOS
V6OUuI6PHU4UqcrGaiCFjFVgmvtPywHutzLSmJoL4oO2gFvNeZJAt58ch47Rj70i7dLyif6U1NS5
n1MdZHnMP31ugilyDY9vJoyDfgEFou8KscFfllOGUzgKOdz29UQZuyqNi1nU40z4ptlQjfSx5v5R
IIJz/QW1Va0d7071xKR50+2eJyBQuokUIPSrxK3LTLz82tq0P5JIRyJawuv4O35ThCJI2w6jDWUH
6fjiBTHdfJqathS2TaCh15czZfZVWD/devx+cN/89zftd4JjYgkk8yweT01NnUPYYjx54NjH8JFW
l1H/Xtd22rRcDSgexgyaNSlsm0xVkHdOT0sezl6l64Yr39zKuNo6mYxu0xFt7HhJTHfexJZWMQ2G
z4+o6TtWAwwuXx1c2pgWVEdJxtPbtEaghNT2X7ZmgLd9y6FOoM3FUjh6MDJpgTM4dLATAAkhv25h
2yp9v09t0R//QDPdUUTB7rEhQT6UfAkOXCn2bkuiSVu09hjWft3psPhW7kVT9vU1ZnOGmkI9X2GU
y7TQMo2y2TlO9GQH78viwwyo4Hsh91csY5iehlIWZKdclG5AYtJYCzFquQ+30YP+xdPwaopq4458
vtM/T4H0eqyfORlWe4FqUo0CeTRFbUtVvpqt5OCvE4/XahuY/pMFiLKU++ozeB0jNEAxuXV2fKEj
o1fm3oNFxAUQpxVMNcfPop+lllcSdExf7oomgqJFB/PeOat+V0TICaivd9vXGotnUlOgYH8tSsGj
i5fcwaALhZi+cta9l2hfCg4V3dk4dV0YZEhxON3vA7DdOlQ+4QAw/sh4dRidH65ZV8iSd6VbQDDT
2d2nzIuCD481QlwPC6sDQcOHkUrQlRaZcGjzbP/EG23hdUEft/u4G4p8Z/xbuyuSi0quHfdVIKnG
vX6nSWSlcxQqVB4zec8LLx3Q9y+iwAZVZBi+mE48UykbNL4LQVlvF5OxHOS5xafRobICvcPbANCT
FZAOn2d8N2vQgNZVXXT686HaNOGKpfdU4btS0ry3/vQ7CHRsTz5g1ZRKBRuc/jZtht7o3H+PLkKb
hiKsRwon7iBD8EkrMcTxFiRWD9so20hSU545gLrUXEh/JSxNK7v6K0/yA3bCMiNIRxDKc2jchjx/
l/muhFsxLSeBbBmOrdNn9SnuNE0mIuTwOIUowFEsjch1FoWcm2esj+65TfFdPc3H/Kc6Au6CXCRz
JkFyP6leZuUxSqsn1uwXH2Ux5YRIB9Syze+xOrJ0NiI0F8eTT2yYS5kLMZfWwYYjdsMqwHnoBh+s
qEuys5sV6RgLko2KeHcKsLrFkv8+XF9nP+hh1Ay0d5eTp72Ol72IiODsTj8ce/TPHdY5x0MbkoWK
qjxMA9MBfwjt0JoEIjXkp8ilVSw/8rv8MWfcOpjBz7mLxOYWhqLgIZb8JeaP0FCA+xtcL7nXLdwu
x842er2zcTU6bEsusz7P2Vvafvi9aCEnRsElQ7Mqcdn+oDN7pSh7rlbiLVJr0WPsqXIfiBVByFZI
WEOO6EZQk9Bg3I0kBal9uCz43bVhOxSaYQtpvGZ2qKgR4L3BqQiULJDbOzl8xQofgZil9fNZQmmx
ju0icA1ze85RnDTWv3kIHnlgYL5+xu5mtX9ipDzU1pxkMB6fjgH5TmEJ+ruXvDxJtkO4zLDVREGq
NAoou/8BN0HbVBg2qj+a3qsm5BHGPPhEHdtT3UvVxFT/DqcT98AQiIjoUHhEBb8+MZjin6/ZgwhR
jJvadYuC08D5L3IzisqmitOo1eF4NEXkKrQQASRTPlRdeSr1qH0pUmOAe6cwBao25OxE0XEUTkTy
xkNn/cdAEH48gE/0QTllAZqUklzeJwgQ3TzIzG6+cumjODkYwXN2g8cWd82PNDUWc7brhRWCIQB+
sRWKluAmiouIGwVIVdAr4Eo9UIW0dj0lfoVR9PiQEJV3Kh6hzrQJqn8eXuJjFJVlgLKjTRekjN7b
C4SPUUGxcrXnmstUY3IKHX6guVG23VJUxxKg36LE2x9UIUPoPSqXv3hMRSyk49Hg7Suaa33NDGRZ
TbQYIkfcfBILR3xBmzZQawvOshPj95VoMX+QNfQmS3iHtpKK4sGtVGhd3F3S1YOlGDy8pjFkAy/4
J8lavdxITtxp8e0EnZuc/ow4cXkbZgnuDV84BaKXMj1H1jP40LFsYElhjzawKLmp8x4fwjQT2dp6
bhXcj+zlAxngr0XJod4ZIIhagp4pQtIfTz99uAdceV1EgyEOSUS3+5hGIN20JHk6+okuRyoo49RK
JmG0tbZqDHCWZWSmOyTFPEwA4Jg4HxeBytwhN/QH+L//URdCIu1NPUxnyW6OKqO2WI99Ny+cPLet
k5SU5ZVD7bpmctAjTd5uzPl9ZHSyrk95x3mpCBi6v9x1TkgueT+GldAINq9CLOHTREuokE43hcsa
MQ5zStkEwuRZX11aoUjtrSVr3Bfo/3tKVHHp2MeIsqhXgku6rUW/uJY7XDVBVoBY3JVBdPa6HNgG
JtIonnRSRbZYe3iNjj9yW5aCIY7DD5BwTUdr1XzWna2ojIS+R762aA57pvLMzOYjuBxJEGTis0yt
PFDxSFD/LqQe4Om3UeB6TP/0gZ3IICFcNCJsJclPEvy7etvM8VkpqvoDbWfXyQBDZBTg/T7S3w9z
GYwd2raO9hF6XdwPJeFdPpqI3pcYuMEBeO/FpPQvWPYpWAtbhVkiu2n7UGWCr8NGybEB0j0520JE
eB0MH9F8rx3cYcakErqjaSoQduk2Am332urGE8KQBN8a1AUWjAEeo+AFZsdPY8S1/jA0dian7Sdp
JrZQUTO9U2/Rc8o12Owc83/6LwWyjbbTXVgahyQgFp+tEzUzyfIjkmcNL92gilwX6vYF3vTWU8rp
rhcSSp6KBfPVEHboTn9saCvtO31hCRiP2pxdO1D8dz/zCDy1cFEpJEaPU5j98+YRCjeHKKYhnP0y
zmVmuuQTUDwVV7keBeAePRbc8RZLEJO1Q3Y4tzVxYbg/IYqzPzg04klxBxZNkMF3kjHd7rM9jLCx
9c5p6i6sPZTWsIgSB3vmqJuPq8LQ31QBf1UC4zgY09EE9ONJjWe5MeOVvcARV0GsLNxk+oeYsRsS
tndstE1ZHYgm/OMOU52oW9Int8QjuPYZtxESFzBrEb7ubj1/NFk2kutoVjjppB563H+6rU2x2fdw
XaLY0c/IB7fhHMwQguc5uKsbC/J2fEKdyZbCh1IwH82vT9O4zrvJM5Xc3vrBZgWSMv3ToKifewg1
x2NvEFfUbubAD34HvsLlyH60s1tfSkUztAaNKinwNMPdcZWGIzKIVMUhkbfegAb4hiPF19FZlQYF
2g3+JGsjveSjiyHCxcpyzFilep4GUM/Rsq5WyMqZ+GFutWXe4OwZZabyqUMrT33i3Ym89P5r8Qkd
OdU3cqlGM3DYy1F7yjnqvXIrggxp3gKRior5mhUTONYpZVoRv6ZCdNCnKX/uBOJQoI8gEhdkVRRG
J4hZwn+doObW6BMJ/Mtz+H53AU7YkS9VJYO2VPJkz+QVP8RXkMxHEeLriaCOz/16T/mXO4uGN23C
4nN3uo2N+PJ7wz20rP+KucB5c2keL0JQDTMzbO1a4WL9Yxzj7zzEN0CBLn3Ye7vwULyQVItH7V/w
8M6Jp/uOazevolgYo5mTITq3+0xGrO/ETOmViibcrGuMrK17zlys6F6imDxe+U83gdh2Hp0SfB1N
waR6brbM2lralJpymTX25VVerAH9mQzDqH/bHISLw+kU2s262QqcsvQ5iGG3GbHP4dFqlZywShBN
4aXiUaSc71WU7a86RMo4I1ESCVGvypyHvKlHp2FY3gyS16nOVISoiimifeKBuNDZgzbL3onGoupc
oEbIA6yvEsl0rI5LB+HVmawWViBPDj5Y2EoQW8Q2HGf0eDTaMnKo0fO9ZfpzgbDM55CWLUYfBuee
hQCzA055hr8+GyDeaeZT82MzcbSQsnBiKVXvGIKENdM5zUk6B7hlk1HW5SfTzXp7J0PuzHWYQDwO
vC1y3DE8PQHwn8BobkTcKxBlQF8MWxX7JQvSN/kpsTRsx0822o8mUOuPnrR1l63tgwEbjwfabhOp
sYgK5QBBeU42bf+DQaBdfnHjktSJvXktJumGQIOINes5OiYbpcfS/ugKGE6DTlyL+4vzQ8SNnXPh
oPlKUGse/+Ac9qpiedi5JMJW7wps2b1RryfRK+fH/lG5GIaEtpdt1uqf8/zWDhPVSdMvx+VzaOKL
/HmfTU3A2AN2H2EQU0sY3Z3C+9wRUyVkbwIDNW7sytKr0Ze5YQ3k0fcIU2vryCkxpJxrDtbALVCH
sBQfPmxbI6M7ZI29sJYc1sSzFhJBgEsz0gyPatRT64lG5XieJlDZe+dYLOu+MbYSkjGrNfCmXb2U
m8Q5e/S7wuqVa9RaWvDN/56sleWLYQpLFuTkiTHEvpF3Ccj0Oc2lPODN1yXi7ecVKfMknYCdQzh3
zv9OTsF5r2LzAFd6zDXs+kfWqyhQ/YARogmrBu0p8r3xsWqipoZQXaJcGruKhydtat62ndxBGOVh
IAjyyptU3Q8FBwk9QN9kDsxl+0vmIFU28EIO6/ga0XEq3o6pYQkQHhkVRuua3OA1UDb7BX4ClUFt
qPhmtnQNqR4Fs5iOqwe5c8AVKYs9O0mFgEw618B+w73WUn3dGAWYhsPD4i50cHT8aGngWAGP0NIN
6WPbiJjhDnir/UxSLBTarYWI+HniXyd73imA/rxGgCaUTddxqajdXBiduKS52m8LWjM0+euOARAE
MZ7O5AZmqMV7Ui2i5VTDpQ15j8uNRYceLkp3KXwt7j9YcbZdc+TP4hs/RxtR7E6AbrR4BPR4btrf
x1gsVYFcn7zcLVkKRfOntsuhcR/NYTxvL8JCE49EYuirW85UXB1bf/cxCtdVNFvjSFNQiBetajjj
tQ/sAoIFmitmop5m7SlypgcUQ2tdJxJ0x6BHsN+VliV8dI86RAHzvFFDOPT2sYlLPp/WXH4sBaCB
B1Ik/yYkt+PhcHzvJMTZndrGa4LpQaGrc1jZU8eCZp0XLfBgzBbwv6kzSc7/iTUcibexyN27fwJz
HiuzqJ/9K7R5vfy000B8dsx8WlziDIdpmisqX4ro0eZtyLMh4Ht/HRfElYMLibntxM/CkdH4pWX0
D18gcoM9cggfyo5bLTNO+RFVxvFAdPbufqmumgdX9j+GdTCpkaL+/Hod8fnGklSAoxtrzJrlEhsU
za8hlT13dkmtsf27ucDEdVbJHVAmbJopGNNgzZuxjGaHGjOBer8n/NQEOnP0pgdGkuhGdVskPNiR
cx87Zqc3aCde8MSCPOoEv3Zoy3RvT5huV8BiCyNptCNva1RPVP58/3UxXzY2m6+WlPYcFOVaTRUh
wzQRDUVutPzKDfCTuOyBxp81pBZyUT1zG+zSqqzmagrbZuSWdztbjNpaE3ox5I288ODDZZC5ckIR
t+uNC0b+kCYOoPBT8YcZekfJ887Qq2sMofiUNiP1cTsvJIZVWblkpvbwPY+ALHXLrBt8OhR9ROsX
2rfEtXkSvV+1nzntpEM934pW/3+4UsJv83D8KbMHOStvrgXKVZGfg/tcIodrOBh7/MO54/XWCayQ
uhYfCX25kMAVS5HQU3pE7OIs0lBpymxw4OB41QGMpCJhNPMpCVj1R7IFK1FmiG5Z+LjGxBOOm79A
b9ryccYw8xbF43ZdpjJO7aTHeWpaKEghr1J80uRfDcgthE35Q6nnjfA7r9ZTUyqDsyexgDpH5Ghz
uycpj7G3kVWi1KZ63eh76QZbRErV67BPjbduF10BGPbzONHI2gmv0jfBtPgiLUzTkA36xEzgYLiT
TA0d3T86aIBxJ7kp8+Ic4XK8HX5/alQh7y8sF/5IB4dVL+BMEaZ80kGGFv6uXmG9a5w/u/I4818S
+0B7bawy7hYLBG/sf9asGN8N74KjHf+UsPEPBjwKtyuRhjiZlhERk/vfQWzyryVXdsObQ+tku0Wr
gAfqbK2Fop8rssLofe9s8Tad3kRpD82fc014W2euXgw1kcVa34jQI/0bM6gN5fOzFVU/dLgLWa8n
VYTx6FqaXBSCTwnxJOlQjobHENRAXf0vZcZMOVikB+6pxuncP1V0VzprmFlxhJKeltINgfFiZB0T
QbFx0a5g0c6p3qaaoz6oo30pWWmC+QZgfQzo58FpPzNS/Izvn4BjC7Ju9+1yjRtDdSP/kOdXb3KK
XTR4NUNdkYAIunHGY7Vznv8UMdVwx9R8Lq+UlbJuAYdg7CBCBDlCoOOLkDOA/Y9+JwerXczW0yob
vYZCjsLAMstnCMmyJqC9nf7vDwtwRYkDnWxurc9ZIw9I/7QRB4bEH7ykKrL9vExcCEjMQgMVITBy
tg0kfuxQNrUR5ZX1bMS7X4OrPGS8NTOJcnxxrpu5CSijYE+6zVRUHnoeOLcri+YncU6GTOikT/Di
3Bj8szRcscx33mYAludsU1D40CZtF7F6ej9tEYsifByjJZ4z2RyavDFkTplMgQreYzkrtsbwj8tF
ELtJ6AZ0y7FMzybWPP9ldnad2itkT2Bqpz/rhi6LqKqaavgicomRGJzC8ishHD0aUEsgDfs2Z+RM
LIsJo6rsvF+STuAVXSWIOjPF86QwB7YdF7wgVC8eFj1lmcT7vOwwBMpZ808z17Q3sgBsN6V7JH92
r26stfXdHqazYl4+HtGzAxQuU5bkyTgnplwv3b5FtcpHViEh7NtjkmqAJcXVXRdxS4eGKz4ONlPu
9IDj4Y4g09X1GndPJ/A/iwDynppUnI1wmrNGZVZRNwKdb4wZgkyBO1MwfXfcu+/ArggZNN75LdpE
OvhlryWY3IWPqJ/Wwzdch6JDMJv1/3w33Qzv6vPimXsANQzIjnB+VJSN02VI4K2QkZ989LWo36tA
J52zMjKeeYcl/XbRaWGt2dWkaCj4aH+XpKLJtWv7ZseSgyzbSBCuyi0ZyjPqlFN13BJso3bA0+J1
6qT1eQJDhYlzAxDSJGOMBwFLZfWIyTrBSzk2S5PuWDCwQaqWtZHswRICEhZqRkZtLc4pfnmOzEOJ
3Rc/Qzw75ms0hWg7/7Cw+RN7pCMjTYPzbKnxUrBxA0mu8D5PljOr1kX7hjysi36P57kGXEyqSijF
GUFeDB83H4zuU5JLBJX1IxzGG9XLogIEC3QwfUDM8nRejyMHJZ8UYJPyTesCjARNHHaZb7J+rJPn
70H/ts3Uedywo0/zcqBLd0yOVc+jPq14OvefE8z9ItDB6WuyHk2Ddbl8abBgrLDgCMLCz+4XzEdd
mxOizC0pGXnOoqynpszwHMS1LBGk5sEjoUbY/S28kxtI6jObEM2aJ6l31WGsnVYj8/xfdzoxoywQ
8bcPZVbfIS2qv90Cy8Roy/gFC4sJZo2LLG2mmzSq2vXA4P7sKB9ZYHVtFIaL/YXIUVGhgEBg+SaH
iEduH4M1oY92AlFnSG2SbHH+4BWJrpL5XbJKbyxTZ/ItZFzIwC6OnVjqfnqOw4ulxPopwIwrv0zM
vAK2ZZOO9NRmCCFACiasZ8TNpZQk/kB9pTP0xohrBalHXYYIc4lZybk5izKt0nQGsNr26XZXHY5V
bnDb8VDvXVz09+TsN5z8gx2Vizif8r7sGQRrekiIrztQvfP42dqliDve0hycbsMYNHHMWRR3lbpL
SW6g1TYbJchR4pXGENW5iP495/2siq4I6y9f5QCLj3DUEa3DMnrUUFIaVL9/d5arxf5MheYQxBA0
UsO0pC8gEQ1ikbnznkXKTgCmxZUCl6fY5uTm3KsPzOpiAQIoKy7cssUD1OXRWzNVKmPAej9kny76
7Zz1dyq4maoqcvjNnpzyP6eaxfnFjLJMWgcrkVRdW3p+bWn6wcXYnhl/8Q2Sot+bJnx/0LBKTE+8
Cs/hBQf5ON9YMEbWUTiVnwR2teHNDZo4CVwSyiGG7wL29eQYuhS4JKhIvtomtmZHfTQ2U9LCMV36
z5nzzS40uUGfSqBfKy+BxvXGuckCm2TiUPfAilcjSDwxzFQ5IGDA83FpGkib5kp9SLq5d2FtQKha
kHLDJ/VmVPPjJ98wI2JAemDlw70/iIdQUNXDxWEZdcsOrSxJaPdhsOrLZSU5PGfJoJDXt6eafu9d
tvr0dlgVYMrxrnsfvra9jKI7US8kHhe7975zpYI0JNyC5G3vIRNHqQQ+RbpPUTT57y/TBTFPNgCh
EBqxMI1Ws/EnQsYxW6TDxL3M/lMcpbOozce1lE6YjxA7hpdtfG2jqOQv0kNw1BsRxbUydmz9TPa/
5KX48wwrA/zARVBpzPH00ZySvyRS5zW5/C8H2wokQmcSVUz7K9gWYqPGMaiuG7Wnffc1oxbrsL02
qDLLQA5fqVz4pS6XejFKxOhTmb7FaEDJzZDaMhC8Khu02Xz6iKePo/Ude8N2Fzk+N3IA0VSsXGoV
0l0o6VPMmUvq4NNNKHUkmEEGlRSXBH/tLQvoDmQWDxzZuOL/1OsMBjlalbZQU4Ja87jqCIhNSFhh
KKW3yNM4iQcYl19NZIduK6cbopGYYjWM2LlPMDAIQFkNYP5dnYDHuiZwNw5UhCIu+QKqtmDE+C/q
Z+vupEm8SsCWiP5zawphns3zSH+BFm0gFwoomTnDMgdw/9iOmQYvgkQLFeGxJO3FK8EjLrNSXOAn
HEE/oe0NBg793E6zI5HXNf+BODUC0zasC4p7PFx6Z+WsssBV1ZNYY6Ra4mMrFG85ePL4gdK8gflk
CYKzuU/e9Ssmrnn/JC282S0D0Qu8LhIAXrBFeqY+ScaNTp2nH5V2A/JhA8ubaYtW4enrxX+EvJQq
PogeFriYvuwCWnC23wF3NTssw2xB/mhPgt025E3G3PTx6mCSbXcPgNQuXOE2dBxq4Q0IgWvTQtoF
TtQGuGnawgIyNFCJsdQqlrAqzeNAaSTWVgx21Tnvc4AthFn+BBaO0U95Qv4Q/XumEl2dvzPm6RJk
T8ldh4zMAduRwWgg8zL1PVGuDGcNs+KhhwY/5kvpBbi5zBHAcwuk8Ys91Q4uEQ9UyShzAENAuthH
8pPXQ98XcjN5dMCtrrLO92RtRLea1dILtakjCVGS//tvhsFy3yp6mNV5TVhM/uHQ4AY4yjIr+Bf2
0T5jMW2UEUwCiqiltZe8ChcQ/I2Hd5zNu1GuVOdgiB2nmF057O/oKPZI6UqEzWyremPmtvHzf72H
MK+hIYB2IwJ4NhVK0zseTQksj5CkvR2KXVtO3J1vHq3h8H8m+h78QeyGnMwHttwpJqJ5dp1TSYqs
Nx4FptcqE0CXk74gGj5xORUlm95lcy15JIw19TvwlBfaB9gM3QObi3JuUgdjNTDZpIzNF7KBO+kU
UgjIqR8mnq0BSiaCBwNGyjTYFKE5ZW2iJEK+Lr5VGjEBsh17vHnrddOAFQgeSfV4JogwYzRtrNxG
eLzlPMPJbFFuEA0TFjfTBCyXnQfuSzBhJlTcqP8GferdFvW2axJqCLEwViUwit5yyxbSpAeNiVuw
XcjG74LgZG5O9fL31wcUKs86KfXPFO1uhpdM3NbRhpbLfwLtetDnOD1mM+ubRj+eGCRBQ+tjrNFP
jdmI365ETJaO11yyqsqaoMYK6RPwrEnpEOhQqlq4YHMC6ukG9M6cY5SI/gHwsq5awygOctYqqqA7
R5NT0Df+vPAu3T8zETOIzd4gOjvFql/AB2/2swLc2tzln3IRjz7J2Y+GbFlhQZinWXAxU7gzaSe0
4iT0OMvsf4EOfeuvO3cuNC/Ghxja/1JThZrAHrVa6N2OH6xh/0aByxAwvaQVpHq1ip7FGXfyXS0B
jH0tCJiIn2QmG+YifUhNkbg26ndbMGyzDBQnaxhKX9kF2RNctGfnYvMKjZGjpapYwfLWPH9KLNDO
66rS4vQA+fZ4Ar+hDascVYr1l1YG7wGSXP8rVsbwU+4aPHDcqqYyjFVcClAfjDgntCB9/0FKsvHy
qX1NLCXjscol/LwEBH+MY9Dix5ZSBsDYsQjO5w0HtJCw2rpxl9v9kBgiU+f2/5nhsnrq80KhIT/b
0B/MDw63dJJZYj2/3ciR4w5btM7NyGoVZTdN2tGy7jypK3CaRjWzQ1Zy+CNJMYcspxGfI2qdBxq/
ii7Bamz8Ud01+Oe8VQe4hR8zJ2/n1Gqehu4AezKmasBvqfKoAY9hEGnq3DIlbxLVb5AOWMx2HiYr
q7TO9iLtZ1MUHBxkoBplL8CznBlNNeJmhj4W5vA7TobnHgzWevLapLeZ2SvJWY9tiGP9sg2Dgtp2
vLT8xYakwX2E/OkR9zNRJsLWZlKX4jF2HD69PWv9gY/MmI7mJFQ+9lLs5swfSct5edtyoBNCsS9q
K1+HkVmSj2wLUWYNUbKocln7C4yYZTtsMu1/SpD2IIB4lpc0OIofXW1MxWEKwkgITS/5WNLqyFey
HfmjMI7IJQqS4HkIQBsOgxfgbLJ8coImdIg3etke/ZBPI4t/pwzU7jvYlXsVyQjn1vgWn/Ra8rqS
9uOEDSJDzjBhtO8S3//dhW/bQUO++tgALQ7Hnl7TFpYWtsr5x640ZMcCafCfpxTwOqfLIeJ34pS8
e5aM3sgeepYDLFmtYOwoiAKEIyfcwp1ANVVHJmxOF4urPR3BBIOS9w/kNADRQOfynBtjDzMibBBQ
mwvodV7RLRwhC3x7CWdkxu9H4F1f0Cj0BLb3KXjrTNeEvT4+FQ+hqxo+XTvUjKU/dzy+CIg9bsBE
DMOLFYiafSacIjeJLo70ircNSqVXpIwbmzu4fpMiCDKN9ggs/e6cvtcsQcT/fDgbAPQ4Gpna+94h
r5h0Yvmo8yIUl13sozKEnFQW4VIPQBU4aBHGjOGVeT/4uQQ5ABru4PcehH93/AqhUYy5gvvjV4ou
SSYHtfySwac6d0RUr9tud6htUs7AetwDf4BAagcw9lY7BhZxm7VT0ph6Fp2PUinmLrVuSZaZKtJL
pDl/3TdKrNcYxJetxCofPP/NWXzCLGhWQGq7sxPROvqqqjLudJUj3CKjTXiA3E0YErqY+t177rdE
akgk129Z91G5iYFdBQLwQZGAn2R1K3yDposIkSRE0qjjpWSFz6nC80xxoYEqgLvNoU2kCW2rH4ik
Mgb4nWLFs52iazK+icpOfKCljCSrYTDbkgAbki7yeRyoSSoDjwNA0o8uQIUjMp2R7LzKfOCwHe65
cKQg5ttamvrgUa2YdAdBCgxl0uVopnTYHnXcUu3n/7fD8K1jpsA2r8WYcpbC+855uP3k4k8XqUuk
RSiwUHh4tlVY8pu1E+xNlxtpC51Dh9Jp6FZY+6PkQNDRfivPjdkl5C/154wLyhVWCmww+qT0Bjt8
lSuUQAqjBjhWCLfcm4cqQof0EOh2kL/D8bEy3GcKPe5FQL1ADnmgBYM8GeXYI9bG6gKkpv51G2ag
6dh8qvPijIBK4nMymaN04c2OzhMb6ot8Dmc7iKJjOnzG3WXivyTDME/1/sommF2X0RxptDCEq9F0
e9yQ/vxkR4eITRIV2jyyS9QJTpBbgM+WpwWTnQA9MzEBUdn2tsfi2ztcmGZdlcEHXORIWoSKiW5R
bSSnf8mFXw7UR1/E0qd9f4ZeYanbl8dMcHp8vi114wokop0CjIJhrENEPFOZg9Iex2pm2q//G6E+
GQs6t2b+iVQoaG17XmuuBG4X5tcC8XlLdGKfFu7F7mTr61jqqautjIRJnuxppL/MEvggCqNECH5i
0tg+em+gfkTiSHImkadRNWkkLbQIJ14RlVJTKQeLMeQZZ8N+XHJqjJiWyArq/yQ0rEIu5wSBJL6G
MFm5Sn6hmy4qJ/QS6eRnV6EBp1/BMT/tIvezgzcGfyDQK22+nHbr5HJLRB22xG8eECsgZ4Lu4ZYD
dgpplK9qYlulpFPFkMPsVRRZ/fIx7hbItg6U1Aa5D6u2+uxleLeVHOgHXBAWJbmZBWAHhqh7TnYD
guiNaZlP/fvG1NU8FiHJMcRmpPa6HvjD/g4hpT7Cc/hHBmRnlHf8n+PVcowqAhum9HiC2Es/Tq3+
7IBkvUpaaQS7oEb1jWdLdbJPfO7vH2h61Tcg3L83z+LWhxAc8sdPsyFjE7GWztv2s2ZyPqTifIaP
haa6rLaFT9wGf+f7CRxf1ALyGXQFc7ogQM2qeUIKYBPtEzwQCCkkEcEXwGJ73KBiKTsRz0ZQTGVY
vdien1jPxL4/Xiqicm+XQZv7YoF5j5lwub4eGPiOX2NQvLdDnxWTGoekePKXUEFc4jzs45lXnuS1
nfd+zZ9Hsk/qF01wVL39dQlh/JSXVtO+PBqZ7TeShXQMfAN5qY7lZ8QalgMyA2uKpjnAid1MokpW
00GKVEfGf6ZCQ1zhWz9jwizI3CKVLxj/2x9VyP29eyjxHTutFr2mogniTM+0BkkNNdZUSxeMREM0
nGn1N+exNfNj1A6pJ8FkCz8u5J++DFl10uI1H7KAdyG9umbD9kbBqhlsE8s/u/uFpnMXkY/XKf9k
xkz2mX2iEluk4ZAKQ3qFr34gYzScYhRphKiugg2FhDxRvu3PfZKcYsrqw3wDVWPP/UQwSDQ3J0RX
XbeL0xpok5mxazwEVj1YqkKnSfGj6T7aZ5glwObwBQMbdRFTly9n5CqxmTqPJfWuZM4Pq+rauuy0
bfK8Qcvh74LRJMtB7x0CmHA+xg4Eg9/3BdQeBZqcSDUdxbTU7XlXiFfySwABntcAUfgCFNZNDSXi
f4JFLzmQJawdFZOuqyzhfg/4bZVeUDRdbaXNxxbT32/6/88MabZklKDwW2DH1K3gmPkFPMV3uQi/
h5hkzGl+bpxnxQknRjlaf6pIPD/bKSaTnUj/gL9ExowuJLFQgy0lAN5oyMsyGVdtbzgL9v0KkCCj
1ZwrVyovpykkMzwS2+sp8Pd19ytXYV77g3NCGd52gwRjxEU8b2Na/45zXmIp1iCULw6vQQ7ZYbUn
gW35vXPqypmZ5mcPFApUklBZc9EvcArhgFhgsE3Xn9ehLjcjUlfqbCXWBBzBcFX5OMqVxeTFD9Ja
V64rvIvwtWDghBhpCTseKTs3mWZCfQlP8pt45GhacYqT2wvrylQ18N0VxsUwSHZAuY4e9B41lZp9
Tb02bWB5GR1zP2N3FVgz5bkMxLW7hEdTN3JAMCMdJ63mti+lgT9+pMv+lphEewnhOLsnE3JdzpcM
/V79KenHKHTxePtZ5oDDsWhNoSruL+WF4lfVARDKcHltbfZorVlbpNQnsL5B8tVHRCc3z9s1qY3T
mn3+avgSkuvTjcQnqBhJaVB9Z037b594B8VJiBqythMDd0nYcXtBOEYuf2sKgNbUitw1Dy6vlzN1
ZX0oOc22W6TLxtA2N3WTVfpq30FJiuEcyel6Qe3J+grCWK3wYvanWoHwU59+GoIDdNxorgq+r9p9
bLHjeviYl7Kf6oom478u23YfZNCTpI5A4qmLVtU8TLBnS/7GrY9uiZu3TO92sbKY9vh/GFYSXlLV
wQbz5rDKT67gLmInIaACZFzO3cLusn/crvJEgt7CGI+BtjwLiMKJWustkNCI5z14ktbndz3DeXk+
cSx54XyGuvKIUlsjTt8tpnSjqfo9LZ6Sv+MepgQI9EL9iO0tmSG88dnorQhJ5GrsY61hxxLd9XP5
mIx/u4ME3xppmYrCNN82YHGVx0nLyjSQN9AbgEIkFDQyhUv5cNC65LdpdGS/nrtDi5fPK4NMuMs5
PsEEjQmvrgao4+zPGt8OseYVacjdYtGrcb8l4BZZ8a0h0Jef0uwaYps2h8yT56uSE1nIM/T+eNXi
O4eJyFg2UOYyYeKoBteJtgagJr6iXpWZmCh1iwC+K34vp5gLNQapNOkm6u8xObRVJJxaogbUi9ys
CUd8ucLVyRk44umWuGTHYseHtaQTVZDlJr8jJR3g4HPNyfIPye4G0oMTUkmF1K241T8Zvwe/JtQc
GO0w6WqByWqA7sE3YLCagJhF1BmYrS2pBaxVzTIYcDkHO1vXPSTcWISmoIcMVpd+urhWOaPDQiP3
ZCkSV1LM11ZtCCebKPza7HQISUlJmciVpZaYZy0AhyqboIU+EPBf69ov0RNfRi0XA+7MG6Xw7ING
4JDcPSvujjpMEqpIhncKWxeYWCnfbuhP+Apvi1nR5LvwbzB6VYWv25Q9LGczRvKFrEMM9ZPqLxYL
Dz7Bpcyzyvzvt/ztFl1qf9iYiFiO0koBXSDR1cIclFzlThd9a6JsBisSmjut1fc75UYbdIABVap9
q9J2ZJ7WIa3R29KkYKbxKmE2fJ63dsDb0dJbrhwowMe2ebgsVSedjOpJDfcuVHPiWhZznCvZpvrB
LmUxVY5atRp+mTBFLVztYSIKXYGyFPl3YdaTWEvUYKd/9j4tL6+hhCk2idumeazVb7VXiaZk/GDw
TtrCRD/1UoIWar67R+KML+Kv3uBDw630/ux9unxO20146I3cC7igLkN5TOZVua+FoEys4VPo6qBi
uS8Zo3QkZwOMS1BmEaMRuF+LMm/ddmEpGEFxbfV4kJgayPWC30LFn2vgt5O4BML+icX3Al7uGRYs
xFdkXvdK2IWWrH/SAisBIh9KTIsI0/vdw0VA+HqfXjwcL0K6s/HSNYhWWq6qTCI+eMgnqULPXUyP
6vcbDNJACZy17K3trYcaAB+nECk0PYC6UomALaLCT9exlTDubOXcwzLUQ42dmojZry7dCJfMsAtV
jGiCxhNSFGfkj+xrAosSEt49qPfVPPayyXpy5rdg8++BqCaWlNqSpA4dydXH8piyJk9tGnN7va8I
KqRg+AKurZDOe6cYEjrbQ+EcP++Jgugpse5vgl/qcL9WSkcGqcqouHV6sqNaO2v6dapQPJlulOl6
t4Tt1Befl5IH66JLvv59gSIyRTnH0L4IKS0oGNb9RKOo19c8nfE3KyBac+4nRizGeETKJZkkgUkw
w1cPKr5oN6axRz7ZFnG9/4cpL9jVrEjzeaFuWtWQHKNIBJPb4WnM9MqYbYY8vE9Q77w7GGn6tOir
vSMFN2XJoivhMTf31wS4qdbBDiTUOqaRenhheySJr3emeeHMKi0ASKa52zFmgdMaJ0CNcCdtMRUw
/IFpIvCdOJOoVrTj2rU+PwmxZjYVh2FMODo71Rz1diLp4kZa+I8JZvI8w6LbB7+YjBe938jPPa6q
u8LIaTH3/RrFLgTBAG4sCJJPOxme9FF7Xhkd1OrPH6uAN7frJ9DnS8q7INBaA4wmsZUjkgeUa1k0
4mZd3hsVlbficsItg9TNcpSEwY0Lpz0IF4hAj5+teKs1mDllZE3VPge3l9cnk7Skju6A/g9Fvlgh
2em+5NoTHtrNI17rlEfrMh0KASLN1Wrpo0X2lMK/HxD3LpF3sC9tieTnZKNycjl0E2n/F3Co8TKa
5/Aaob6a51hQ5Zi/o49DuIYQIC9XG6VHU2LQzB2imYlcGlOwUs8wMaYJMdnEUzZv+xGCt7om6pyG
GhwQrgvjKDZbWcXIx5r7sisVY1MryOz02R4mr2iFwP8iHH882Ls7KrsageRIgsTWsovbCY7712j8
uaqZB+lJ6D0fSduVZdgXMPQrglW3IbniVy0mTDfFu1dq9DEu3jPe1OaWAkZTILqbvzDheDeoHgNV
zUNBbE3fSn9wN9SfbKTQMmS5kcAblkxK7pT+pw95ZZMi+MNk5h19n7rxv8nOsEDCUiQ7OQq01Xdp
pZlM8K9iGwVsUji6uya9jJIHn2PphNrqi8L7bS9kt2LJhfDI3FTLwZDGspYgHpDGeyUzG/BKmDNL
QnI8qCqhJMZ5YaNS70KrEqaDnYmr7O6bbucfTQERwpqusPzQfF4MajQQke+f6XyjKbHMo59HW9IW
dne3xHnp9O3nTJoxMoTBpgJczNZpd44dg5ELrfH3HWkVRT5zk8QifF6vwmFpAJf/4V+kKPXcFO5M
c1F1ibbyS4NKMtlN47q9foughH2ZPktjUmFS4rmkxDUzbDEX5LKo8bY8uJhW5wQHQ6r8fNmF5T8B
MxHm13oGK2LUhZA/Mv33TDgb8VlIG7jDrhioQEgdY1Ti0XQkuir4aKEq4WHpKFOTzreVotK/i1l8
hoFfmsiTkZYaVfVV5Wox0KYjiuU1qGg/qhv4Nj0udiKqQ6tsMSj1QQ/tG30GGfopbK/niHZNlW33
qJhyEcFYU51ndPVRkgSaQvwlLLTpUMZqOYPUgRPJqBeafNMq54mHGRQzufLn4OzPAS6aGCoXC56O
kWHVS55pV6Y6tV4jXCoVfBZEol+KVjpjS3TwaxCKeu9x6MkwsEyMcoh1pmBdUu1GaHlbXfUJD4gq
+PMZW1YK1miYC2YtR3w2bjyHf5Pfxi+JoiH4m/Oik2aTbkunukmmMfDYq7q/Sk/sWtheNmeFeLq9
RHwDpMtGmtRgn90ZvJEe2zAJe4L1bGX+KisScjhlFUMiVGyWyVjWOVuVGj5uzS5iSfOYITWLD4MG
S2K2C/Ceq4lDW7m4ztSdWx6Htle+NRQe1op30lWYMaPWs1cICUD+mRSAZ/saV5dmg5HUnNaAzbw/
cyTAhsRIhjEC1XsbVoUAEZSTEUBqxPVzReZV4LwJMbXQL2HrEV9DjOGnMaRi54v2jvrUxz6Z7cNa
V7YWWIruDJLjsMJ3cSozZ7/2oUz1Fdts92QU+KAzPeSrs/ZqYocLU+tymfYAe4keB9ZNsEtauaXX
G19VL3cWqb3er9Pmu3FWXWtndl3IMQo2k0pBoXScY9pAyUM7dzwQILsFZBkV4RhYTDHZvyC2CMyZ
AOScR2ct/lfq/SJg+4kA/4zLiWe/dmkYpRuDc18EL872pQqdLse76ryejLtKaM9MeZLKX3dJs951
sxt71XF1cPuERZdB62ckpG9b5RE3hfLdcBUQO7cuWG2txxJCozmFz4oG2GKW1WEPRUK7hQnOXAlj
S1V3aEb/4zixQj7akt6Y3yx2luzYEQ3Bxd9en3HEN9kD+nbJdKcti6+L91gibhPnVi43Ch4ruBRJ
7qOstlXXOFJOoUwOadN038sRppOGczV7JHtnlo++b+q6zHtrI3i9ieizUwgvPfgsTj5f2XIbsVh2
VIx+WvLU1sAKzESx3JM8brQFEI1FDGNqwQPRExDXGzufHsIcUMdOjLBvDEblot/xG5VXw/BnAcQl
k69rxLEueFJYsyeVbrO+Sy2bib91v1SfgBOGpvexJuNjoPrVRym7vlumJPfqh1HYNQZicTn/hqpH
UgEcGvsc1jhvANkA0anikZH6PeNL9GnVvltduqJFZlXjXbsqg6VjOWACTAoPzUooG+zffLPw9Xxc
3w9oHXRF54hWD2LZ+UN+PNCa7Tzxqq3iXgLuyONcfw7L3xMfahmS1lsErZ6g7QxuFZC6NFaBFARW
qLNinKsvCHtSl28slHsYJ/GiuLn4r3ho4wS6cYolcOjkgSqmOK0VGGNP03PVYJ8OTb+UVLCqm7Dl
/+DmMuX6Z7rclJagK1xK8yF1EIcjyiGTEAlPdloRnYWSzi+u7uB9Bq4756PRYNd5kaKUeawMI2Pj
EV8wxO9WAo8iY7F9WwXeK4AbWSizMfTiik4mp3p0ePumMJfGq0FicaR2xNhbqBCtvgIrkLLrehPO
AAPDtrFAZwydJqrcDPp/oY8wdG5W2+Vbnmu8O64bJS0O//6EFUt9kd6ois3BBVW9tUdeTwb8cFGp
0QbwmpSVCa9JNtEQm1xXb+wvk9L//V9p/kbf5Y7mymRnfOcIfqd7F/Z9E3AKY1LCg+LgWrxJnIAm
Z6wwNXsTt/UwRKMx8VoEALml6VVhUIv6p6KhKa1GB/9fWvwt2WOO6kP3AmX6Zwp64IX4LILAL9JT
g3aWPl8Ylhz21npW0cl1aw4LDLfcz+tLYS8lsiDxpfY3Gr6TFHzOfW839Tc7iMtK5vkERs5obwFY
amn+t0n310+QLX4ASqWn98F5c5f+S7KJZtZinn/CCUQ7ozukqLjfMqJ5Psam4iST1SMF5MIrwox9
b7bbFSrCJX9n+VkxoO0Ru5C/d2G+87vbZx3FXoDbzY3RUwNXrYIUBVT3kemD+6//I7EJWFtz+cx6
v4pdowzebV9xyclHlnGFalUBu5ZHcXEsLkqB9ewekYqWNTixsLYAh/6gToLn+oq37r1kaw6xSLAd
vlPTUvhF8/uilEluzh86yIr+0P+bcIIvc6sOMc9WgMPl/VEqQDt0k+2+M22ozstCM5buD6iv2ghI
PzM42lszCXtizxhCNzrSJXFYsbJ2HON95qGBwzaNVRea/yLv+QXTyv6mK0PSA4xofhRDoJgcwzpr
4gEYAsttbR6QAKqH3jFESFWVP7wegw0Iymp8nJNC0aDDP8MKRwx78bUHeAj2MWojPeB5uUlE+rhP
4zfAYm8VHk3GN6XzfN8EjAQqNmEU9t5MeiVasrRoT369ZiAQTPhmeqJOemLBo33L10jxm2OWP5ak
rxtNDom2Wba550EoXlWge2C06gyYly03jN8mbFf3N5JQunAUsRykvJWJac7yKBgnRHbRIg7/8j93
P2VdGt0yRi2EzdgCM+moSR5//K2xEGzHC4YotRtJYlzCwjnrRrcQ9q1ToNJ50BqavhYGw7TddTJM
pYalvBBXiQgmKCncXWEthVt0xWNaAIYSZjyM8OpG0zoS8OM38Ng6ZCQDacCBVV5VmKH4l8ejvInH
wtpg+CFcd3oXNvPw+iJxNNyxFS+Z15bgINMEsj3dBnyYpyyj24HZb9t/A97z50r+/7vKh5yHNMcU
6HUCap7hKAtVdpRzxSSI4M/f1b/gfV4PFDRhHhkEC1ZrdTAlTxHlfcSbp38zZwe5C2bHyjgCzsaG
EPdumuw9lmcsWUe2e7UFbk3X7TUq7SwI/+hYgmRQD2hgOQsVupeHsFv5O91izE+D6ZwFZEKbMhoF
Gti9tLu/Da6NxANRaZYVBeXHEA6CXg3bgitJVpW3+B1C/vv4CZmVBh/LYF3vrMjAc7ydDMXqNr4Q
/wBErLOjnIN3JsrztuvEbE7Ebp2R7/xOE+dN+2VzvT29VVA0v02HATPWykMejeOsdehh7yK4v4jb
96AU1v+qojYKek0qk8CohGHaD2tikcU3ykyJsf6kids2STfl0WkISnTBQ7EB+dABez7Fzi7nIut6
MnksN3WMlZ8EeC/RQOPQzuhV5hzt7RLzL4Zi5kmxq61N9CpbzZpH1Ylhxy9a5zoTgOMhttBnHq+f
s3Yi1P2W8g0HAIwYkGnR9UzxoBTPqmVLQp6gLT1yTs0COQ3jfvscbegBYv2VNXqTwV5Mhz2OWo/q
EJ5Hg4uZZYTsCxiVykpJJRfA3l0Jt00IBkdSWGUiw3sS8pkwET6QOqWxv4+Mr0HvwvAzHCYdRLJd
WbevhH6Z6LGjCLZvJE+ZwBFMeKskQFr2itPmeMAUNgSnoi1RlPwBLRIKlN96Zfa3eMIJiXie/4L8
qQn5lkWmiF7BMW67L6oQrBwiLR9LH6OLJK/+x1Yq1iU7awHvSxfzQ3lj06Ga2MUGMov068nlj0Rx
Gc+urIcP/HOTPlCDaOOIKvYG2UPzsxwwQ+ILJZXjmiM3dhr8F7kRaXt+8mDJk8oeit2Ynpxh7fKs
EbKuBUc+yHapfBmczqlhOrfiMEZUbsEN+T/XDUZHZjSpiPrJ4MXRKZNxoCSASLU5zJTtK+hDG6Vy
JpCgn/RGKMfPa6VZAY2l/rLB9H61uuu+nE9Hzob0mCXSbZAYjyyPUl7kDur8/ZjkE8hKT4ewA0Zw
+kH0gO7pRxT04ilkGwl3Fl0qiFvrqvqj8BasTJB1WOLnw7785MR/WZguaIHtTwXxnQByI1gEG8qu
u4b+MyWTQIPw4fux6E5FbQRK3Zz6G6Xg+Ke3nHX0ba/VICNR38PDbKGqqpvtth7Br1h/oFjcKg45
SG1cWHxbZuSelNUHXGQu1Mpa82b1iWzwwSv7i8zOsmFpE+OK8lcnzWCeGWJtdAYcVkQDj6MfQUjl
+PwKqRRESvXWS7v4BR6eVh5FNudRJH9lgWDdAv9c9lxFGvdHadHj0Oy3YxvxjoVXwDSkRFGI/0ZZ
ITZM0sy6oTHUd2/Gzn0yWtKR/LVKjm8CscrADcAW62eUcpAfBIRZsHteJ5/LHqnEwpSLn0HxqFrM
aHGlo/GoXvlQ+QoGSuUarZPkE0c0U0Fmtvo/hF6Uv+4Ipidpk9avAC5LUWTjMahylFTqttbspQ0M
pEdYC5uKL4MtzoYP/TMbmZxcnHBaIMDSvihzcqUcxEH03k4pQEEm+d5AK7ec0cyGFvnAv9BEC8Vy
t//M1myu6Q4jhGk/UVXmRs/GSegXx+EOI29AHRWR7tyvaTZLF481kvdQ9tk40rxNJ9hJS/iZzP/M
aw5Ahv1Qa/65uw2K5vHPTOMllqhvZQiZInWOSsL6md1VWRhEwPYOjpKIL/aD1/LqqZqVP/fo2Iws
IQNrZSsiF7nVoa3HIMmIFTFd0Y9fh0Aw8F4U+AAzpG5zFeIvJ6HzDH3IeYye2lKaBP2Qh/YOfSFJ
49PFA9/M8ZEtLE+ejcWekeVBkpGwgIoPB2O2hB+uHKSpN2/M7RgvcnraGJCYRqjckQFuGTs478C2
cARWOMrDCSHrxohhRNPpLQEhB6nn7MN7WLz9mZZBqV4wMthXvXBQIGEKQXozHAOTIwh1K622aWMY
+WAG6wvWuho0WD5mZ78C0wGU5t1zDRMn8CHL6FVr1zObdHi/WnjVKt6Ojbs7bfDDATYUWPVYVGhW
d9uVrsFifW9eipjKxcTlAxlnzArRKm9ngyPsllBHaYyxa1NAwEFKDGLdv/O/b2Xi4ozJWEVOn95S
gD9YPd7NYomYmV/13UvncKkTgnP7satCCrZ2mtCu4z8fHG/0aIN3DLR1C1uBJW65RAch3zjh9jxD
S4zAoxaxaHoUTCS/LrhlmLIXzsLJp8AFSY0tJpjUQ9iKEsPEI44usLG5FXJJI6PX+G8HgBZ+0WdB
077ivTqfUbk+DQoyfo9cJrlgCvGpDMb+oxfUzvr+49h/vhpt4OlxW6OUkjv59UN6Jsn1i41iVLMj
6i/F23D+mSCaSJLxWtyuj5dVEMRPc6eQ00nfVugJc/VJjfx1332l+rsKgphhaJMRzgDrgNnYZJZD
RWUMpNjp66Sbc+qzOUZ+OLlXwY0QrL2FELtFjTIP+A0Np7kftd9gQmVGKDaTn0N6K7qpV2sNxTko
GO0QaR/00U3O4k+73JBp9sUrgWLTC6V4mzQicD7dfGLuVF2qYk6FpdTSmjYbfpYNTqGCR+EfOOKk
IEu4S9nK0pcFGnrzKdS8Ycav80ZtjUzBQRrYtT9M84N9+JenN5XLaGIxYJjKEXsEszWKMFUuq1fR
6p5HNV2I2b8KkqLFCj0HR64jyyve4YFfCfQhMfE6/UUkSXsKi+U2z41dMn9jxerxQf53ksggJGmi
Vh2Zyusks5y+9B2Bm4LopA4KZax08ANOODC/TzwgF3vW+vASjnXzuOnuSVqA/p7OPmKDjGVSab1x
pP/ZRoSUgXwXbiibJSiPSOr+wAW48ARcHxbnnT5VyvuwO0duvJyHiVWUxbej3UD082iknIRiZcx6
tSN7vrnGKjjHPHJo4EGUJarDtWRsViZUUZ/T4ND2/KV0qLPkGJ77nhiAWPmjn/TReiR4bxsOLaA3
Wt4FbnQJxmdGxp4FUm6JRpxDuWA8A2CPpdbGJwWQhHkKHqiHwDj8dnwLZBCcTFy+ypduiUauLWoj
eVV9A1aOi7Z4euhPKza/U6XgD/mGWjcjzz7CB3+6JPXH2RTMwhE4FWB2HxJKVmy8PwPP/zEddA+N
497Jts8X6UfwEbHnAxW02Swg7TwEw8yJ4Oog8+fd4i9bw6luUwx40AwtJxefgWfhlK0j7ttjQ297
9vNstkdlHPbeGoMrJsH46unK6O/hFp8KPIr8WiLjGU+s+JCaaXJ7T4CTPXXWu3ylPYHKINXwIP39
PPV0+NmNCqVS8oPC5n8p6UtN1sLXaob+Ft1l4oyjnGNs8hCs9DXmQ3SL2OKguVzZxwQv/67Y4Pyp
Aby2t1xDfSuP7sDNA6UMetObzzXjSs9czxcLFOhm5RPOaMxEVsK410p47L84jqyRzLXgd2LherL9
mrojN8tfB83YnOcSCiGUHoYmVZKYVccassQfE5oDCkcfVs4RRy0iykKXERDVf30+yc8jsuUgAjsx
24URGp67cWqtRRXbMicg4mQs2tVUDg1CsMiYhov4sKIr0DIy/tWohrsKcc2rfFIccGXshn+GCpfL
4nCf9XOZHyu6YjuEqudRfDyHDo/ChRXzCLaVOKvxBGd4GhQKMpUkwVK+LY3CJwxzME+62/boruIw
fwODFhUX+Cog5SfuQIt6X1SN4KIUh34o1xZboxjsMciwolh86mJRuyakpVwqgj1UeLAWFsk1enRn
d4ekKhWdBGDhquY5TruVHRIZQcGH7PC18qB0FqYZ2Q1p4FUXWEvpXxiFE75ACk1nb20wOJbo4xH9
lAj4vvA1C/Co4amGkm83Hj9oBzLeyIBf27+AD8eoEuzBafIDNzQ0N1hoiNrvseXjRWRtTLAMjZgi
MW8CwroGPnpFZRpFWZGhYEKD0bG2P4lUWjfySODHfZ3vvMsvbfMRODHAMVYlRm5D06wuZ3Zw7YXn
4XE1zmkK/rbm/plCrtKILcn4MPc+lOePgxjcHLh64/4CcVEk8j/DZWu9dy+SI3GeeWtxAIOXIy9J
Eicn82he1vTeERUH0nFTcvVxVBQGJ7Pl5DBDX/+hZzSBeQU+HxzFgA7Ate1/fxqZhsZ2bPx+giwv
cwQxZaKnIfp5rsdRgbuDWG7vqhIHvS+4wsa/EIV1xdBEiBn/Kn9HW6g+bn05l9PCkbthNTOO2r8o
D6On7nDRZU3nx9Txw0EZOKs7iqLPMVG7eVll7X4TdBcoOX8P8/iUI3trhIQfDvu+kuxjG5OcdqP1
K2wb+YXDWT0wBNikLe1kK7DzzLTJcV/ny57Ul4v0SbOHwFzBuHe/yZC0MA4Ga9yFKf5jfpU1yNym
YJb8jdbD40D+LV+/fsK9MqEip/FKvp6Ss1fCf+7jYbkwScQ7j6OdRbGtiS+5KRaSN+kPY9dEdLK3
C7ce9FJVzn0ls2Mw3kKWwl02EzSaMqWFFNeu0ajx0JM76cle3IBQu2vLc/9xdJbhvkg/gu5VX64T
yr4YGz+ZAJvPas9Hfx+K1abPpn/GVPruKtnJSF05fYWpB476hS8J9yK4oen0KBbScsbK7BWjSbX1
w/PLUV0pNbPrhnMeXXPpwCwXVkaj8zSKBHs8UIkZIVV0r2fknSoIiHiRda1RYCDFDbnKAt9v3Wtx
4D42SnsOEf0r1p1uKqIGueor2jmTAxhNYTDJonMSVUodujFRbGUJtXOTUZlFE7a1Rhb6hguqsRe8
STI5cllgXdc/fUdVMr626X2HaA3zh46RQCosZkQROCS0/Z4JDGows45BENkLoJUyHTFHxGUpdqxx
BHV4WPqEkke7oaG1goORXIr25aM7jiQdb+UkOaks8JKYhFioOpQXv6czIgbBmCuPFkV6Nb5kN/gB
9xNju2NF8RcYB8eYk6rUD7hpX/3nNPVeygtevIoAxKFim+z+15xXeb0h3QGHHJz6FkJDgffBk2CV
08IP6mo9ylXASWrQXi/GK0OJYLvjd10OyGSD3EYnCHxXDp5jOQUHRQc4vOf43tPw35LGUrZVfAoD
xJQHf+/XJulT4eMbRYxcpW5NlREDArooEPdJWYsf7H7b1j6vV9TbUBVgny4srLCCvLNmfSUX5a6y
0FXy6auuA17cTnFSolQw1eZ1XNBKcK2E1a02GA1Aok6PiJAZbk/1KcNB+lZdJx8XHFwLmrtS2CUR
Ws+NfopZh3oDKiot5scQuoG53UVz7J3OfiJfOqSBcix29yq+33bbvxPrJHFkmG4Xc7y9xM5pqXvI
+dN8Y3bmmlX7D8ET49JltGOwGHIkhvVSMvAihtEhOR0rPOUZY898i0OBkKyN5UvALipJ/z+vLcC4
LL/xA6gXKtKm9FYQWWjE3nJM8cGzVjUsCcDYivBadSGawO/yk/kJKXWjKfRZHgfrTgXrHiUKgVsY
N9PiFVfDj0fwWPI1guOyOmr6hw4jyJcFaUQxLWx1cspGZfLO3gc1nv8m27wUDpycPVdwGmwefPy/
mnHEOwd6BZWZenaeURryLLKssqTFteT2DigFlhWguAHD69V+gjWuh+UzDAvHtVHgfOtUy9hw4YIy
f23ZCY9gWJGGgRMgPJ7sn8n1zv3wRXl2vfPSe8Fa3bZAJl9Xsji5q2dplXc7E3T+JB3naujX0e0e
YcPcLSx/l2JdTtnS8NaBX/2q1J6RkxQzgLhnnXgjidp/meNIh10miAWhE4TMOgq4h2AQ5Tg9K2mi
/w0c33pI3AS01OPsqgUbaXkHx76aC7k/f5C8u9+fc9XqEaqhmw3V8N1YB606ONe+0qqTkam62g0y
CsuGH1t8CvHKcvch4XN2KzIAOZWwmpLraUYVFWnOqQQW8P9OkLJ8PLheXVRVFzoZuvoSfg6icWHQ
gkF7jOt7tHvNopKM8gLvTX72dt3+wIU8soYQvJLvmXQWu/HKIesEDq7NyghbiuaTCXJsQlsvt+bZ
QU23iY+BPP0BQysqs9LvY7+1SBi+h3ydxDXKwFd5ppeK1bO8HhCkK4ICey8gpgM1LfHaRgy06uJX
Z6MYIJ8pNv0YwCbOUVb6EpphnG4r38jQlB1Lit5yGhUnk4FUyFb6l0iL7jhm4BT+45P4Ec4RFCSd
44OfYJT6dIBPQ08nTNlckyMEkc5rkacqpTvlsLZHy3NsG9HVndUxItQjWhzXPs0c5GJqiYHlAi9G
tkzyBY5JWD5yweHyuqq3wMTMhRlr88ucRE+eAXRlVkp4nrqLdiuIdyw5qp24y011P/enUGPIlHWx
uRMh2ygCD4olzbgUSUmWX+kSvdwtWM3RaW5RVaNZoKwLF5lL3Ql0Y5wUVHD7CiZIP0FrjrOgNG1Y
2TeFSGXWK5Ld6RS32dHcGyRhUSYtKbY3ZuVAdfUEEorT4aRlvbNiosTwdPhqr+GwaR5ycowAVlJ7
eWOex75gINZmy8pkkM87oq5lfaLqFo43gnjXiDYYnEul1E+rZc/i4Mzy2ZeEec242ZqZyRPXYYh3
/zOdMChMEl4Xy2ex4EteHyuaQBkNNi4mJ2h6AUoREtSBljdxAwVg9mVAsJwO81uBlKmyS83vi7RT
XQAvvoNw5d6Ex+716pYr/vcuBt917+f6/TZ0w6hLGr9XgzaRcTBQ3F8XDPIGc8pb4MJrTCkCyeo3
P0BW6C0NPpIVXHdLj2Q4Tbn59EU31BS19UnRkSIIsAp08U1844FjvsQAbzgZVooHP7r8kyekpqxr
5td1LV2keeqnmnYy+QewlfgnjGKKtZIk87wjv9XU1pqZ1EFPJSOLuMQ2l6WYigxzSDWjs4y/yVfj
CD0J8MxsrgPerR7SMlcP5BJJr7rQm4EmArIixL4IjawsGawirw+naOPA18n+t6y+jaeRzaE3Rg63
dTFopsWcixmh/tcSOxV6POV/CO7KV57f2ApeDTssfanzZoAmb4xPupe0olwfmVpv7V1q7OajYdhp
JO9RB1KveCGlqTxtYTD17U6RNujVskVTl+ssqoOUIrD2B66Uv3QDvuZ/otTmcROmzbLE6PBfsBtA
G6xFtQL13oVqDq7SBmtIrDgAfmP9uD13J8I2Aysder1mepRB/INs8UUV+1AY8Xf4+ZT19O4RBYUv
HQWVQVBSFnyfcXGkt6pth03iQv04oPAZKqUenLc4+gHkJ8B0xJfSaCbzPPFvQ0+sl1RGmIHr8cQu
TwPCl6ssyBlNCZsLLGkXjKFCGk5fGHf4CqKWUcjg928gwiUeFUPQG+2+o8OFTzTNKEHg4IRIpXcs
LIcEd1IXEW/IzR+GP7xJ0iAMtCpSe9sfDBzX5o7mlWa/14EM7LzxV1hCukJtsmZOOzQZaJj1Jnug
hECq05K4fTeJHQDA7gXWsThJv9+y9FBEy4q3arCqjrTu4tTsfRmN1MCHUe9GeODFilRab0vgGQBS
OL/r0lZwlpH6YqXyHgt6KDiccpc4Y5oPEa6LZMMNP2222+gkWLXcgXJaatDzcwbntErO37VfASaa
zNpnWcQ9dMvXNrzJrQNx5jk8otcaO/DN0Tuf1K9oe7xmDbQlUjZI77A/+8FJXG8b3dzNpd9n66dy
Va+kr2UXThRdTsZMGl0w3Fov2gqo1IpS/hJkklyns/N96HhWzoyzZNmRU9ChKfkov5ovpsPmuyzh
aNb5dSC5olQPwbpgIMy4KSWct5xv6Sz2aVvmU3b9ouA0gSTbapNNjIeKlNPDkav0vZDRCq1Aejfm
XaZaPspmbELOsTbfSBgqIKciNQ3NzAHK1MEmYAl37hfQY5XjXR8LqCI8ZkSJzse1qezYvR/3mVbx
djzEO7+1wlhAuXTQTTeJz+TSJPFGyCW7OWuKjqexU6XUrxLcstbvCv1eoGNyXMF4LsR6MXcKwTVS
wx08blp96zfqR0c6xbqtbjiDverpl7IZNbsoa3XRLms9QbxmebOR/Jw/VV3TBQrY3DHYi2KCduaa
ImLcn9A8OrRPGm1h1rIakru0Raks/m1EXM1IfjkU5Mr0NQLmKLZ/rWvXClF4QKPDQX1J0V+BJTk5
iVP/IrcYvsdN66FQyuIX2BOjLiOfSfct1bPQuVLq7JB02wKlSaTI6/mIMuo2z58vhCblx6RtoN+q
umrppf6jXoR+wreSpz76SZloxGI94lmooswxqzyuW84Wvpt0oB7CmOHDszQkCRp1ADaFbaXUeByt
feDmau/bMrONyjbexS01U6OBJnhARHuC809ZN9YpY3Ozc9n/B4DVyxNNwdM4oeGPe0U7y41vzN9W
5dpm1wN7oH0Qo27YbZAluoHOFJO0TQ9iYTMpHAU30IY2CRLdjdzpJeRqnGeJFuwxJe7xFlcjgnF6
ymWLM8zbdpGkO/wCUHUdN+zEZomLO9VEiRsd+4gde9oL8puRFesK6XXHkLAzQWrztIS6yXqQQxtR
m7kb7+BspE9ujQARLpLs8ikYM7LAr7evp8bYEO96SpWM5HcqUh42CRGnnwL7r/1DXYrWHsZDQ7ZU
uFbJ6weh9QRTbPCiLw+CAqRJsV/oiHDVs+TQXM4FZLOzdUqlbi6RSJAlTsb1G5qiLoAOVkfqp71S
WTn/S1ggvyhk10/S6vXuTJeqUNQ5sRp2Wphnxpn9EAMtmzGsRP1gqC31FVT57HAj0361qbIlfa94
HzM/9FDxqxx+QxxZdOc7UH1f5aGH2DfI/LaqbBquyIQjmg/jZ2qnKvngZefOEa4tuXlAabz3FjPO
UiTcZW1EcDO4+Psc94KNLlp2+3om7tjz/fUlhA15CELoinOesCWBIsEWOjm69wOEjMpT5FrHuWmi
jFFo4WjL1Tromp1dxQS4PCsYrWZstqmDN2zntc6+iHH2jl/wAAjK+4xLJJXWiiCjjSTAHmRhG9Uw
SQly6BIKi5SDwf05TZI5xHbAZ9qNO7o96wEc/EPu8K2f0QDkg/HucdmKZjg6crX45HfrJzxyo5Yz
q0XisakmcLboXpe0Re0/3JYCsetxPH2oQMpzLUgsFJn6GWBSEq2Iv3hOeTQBRQoTgMmUaR3irF+M
7wNUdQmKJB1whBNWzVHewL4Bokm5byCPjhCn3YhT0BdI888S5dQ2vaetrV6T6L29VNb5SKyv2m6B
y5N8E99KEtNj7+4vDSrVfZekQYvkQK0Dfb3D8xPDZa6jd7KNqqm+EJsx2wPADXF++uqvHy+jZ/iP
B3DsiyfD6ysWysQChQU8kFoT7YFH1KI+3pnMBq1wlkTzVztDE27P9KqkbpvdjC+BTmehFHMQpJpi
7I6r7i8L9BLgJKEwN2u+B+9nq+pkO4xcewYhJ0ld+d1DuTNIULg95/qoZkQLvd9vwC8yXUQqIFW5
Mc4ueVe17/IMnQSGkVcpSuwHa8Y/a2xX94sQLCyMvVtHJga8pJfbiDtBkJhEOhXdOYOdN5Bs8EXB
IU+225ueVoqpiBAgX+SGmPayzisW8+qTyJjBAG3IndjSyKYZrx8qEItU3izeZUWgYtvoG4/SMInM
dlqqU7u5pRwr5w38cd2Xnr894oL6js1Ol0S8zi14FPUGUR0kVYMGCjthttOxnUi0DxshCRRNKfHh
IPenULa8zuv0I9yLIU4YGA75SCNqUK2/SwMfM663PAk9BxWiyvZI/taIChTTO7u41DQ5MVcHXQXF
HJAEXW+Aj43MeFR4ZhQpRKJt1iENi31F+2VU+NxRvCeKmH+dGpOfsw5P4bSD4RaWWOaIn8OvAw6S
gFqDW9iU4RxfswTZMgF7j5Y4q2eIemZTuaN4TJrEQvELloT2qCDlFVdjT/e43Nk9g2s/24NkNg7u
7ArRdeq6IpvFKl5655qHEg76FdQYoTBKUaT9754CBcLEVnczra7+VCbRwYt00/3zDSzsSVJ5PN2B
HV7TuTGCmFKEA3ZxMrqC5V1lESnWyquvCyimY0i7SMA10qEe4wtnzppBLxdhbd3xYXRgOX5DtbSU
SrkJdeJ2X1o6vrXZGrgjkH0ptyCCRCe6GWQ05q2QM8+gvdNc/KLFfCJuo94jG0CIrC2jtT8suNoB
B54MdFa8JtqBj2Zqt0JdyP8Kw9vaHF5cSGhBLcnLkJIyXnD1R+DstroPMn3P7ps+m0Esidk6Q4DW
NgmIngZ6QxV7oVwB5buV+8w7k7kFnOuJh6HstKr46iE/SoulqOT5hKAEw8Hjv//KkpFgiZoirZqj
IDbcCpdI8EGPA99uesRX9kWjyC0zL8opYUfcbVwJonOli3sUt+vwfFqWk1k2+6osOHp1b/n/fjAl
Da8pgIJYqcsxEYh8bDKRPatowXr3c+PXfdonlIxNuGQei9DnDkDKtQJCfwWPnejb1j9ZV4u7ow5E
j6MwAsELsYCB8C5Co5RjjgJcZ3tbo5dtuHa2kLT4t2xzEs+l7+IF+uLH+hEkTIO5EqKlug2byQzq
5bgQDm65lDM9xZn3hIIp7/iQJE+UyDzfmT5B/NLvxw9ytJCcvvzdV9nlN12ZUvGid2lgHTXzyklj
NduQKKRJfB+RcgqZaNSBiIIPJ7XrQCalxjqOYoX1tslwGvEcEFYylhfce2VM6ee4FJ4a16BVAkom
Q3nfRqmjDwUPB/tY1mBmW/8hzgpR4kEvyh8nn7GGP7baZtIgr2ABTloF3OZLoaHsNSeO8qJTO/tr
RyfYe2PqtZOvfy6eTumg7v64j2ikzgSmHUyLzmxV2uYZeAjWBXpx9R4fzE0Bq9Ug84h3CTYk9phP
OPYq9rtxYIY+c/MQ2gk7KS0Q7Tw8aBEIaOQ3H+qL7aF1Xy3P6TtQS03RwyzBLfyKP3iWXvUIWN9l
fE1BEbJJjz2yTiz8Pg9b1L5TbjZ3eAfDOKf6elce8Bs3TgE7yIFIev9zPZEQRNgalPyBUs4LPMbg
/8WkkSCa0/wTCJAc7AlJeAfFgDWLaAsFpy20Wp62Uv9E7p5Inz6AQ8g9jnQnqSV8YJeGjuLfLbMh
h/PrlvdKA4XBp0OlfU16CwVE+MvIPBQiriwUUlvOs8pjjdYb+Xa4WOx7aComsl77wrA2VkTfHRTH
0NxoyzrgODbSm8xUWMQh6q8qF7TdKuKMxu9zJN4Dq81kPWmxpHbpye3BZQNlQNL6Gjs0H2BFC/mx
auJ7FRbks+9dEhgOdzg6Rb4TwY1snSJwQ8P3Mlo7lqWGgeXSp1wRdEwtomcKYMoXMPVw0eukvML5
vEJgCg+CMNfdb0ZcACAxDBIKj9/V+MszWHwIFYwese7xLqM6zOVAcEceXkfv1pNw9V82wxErLF1q
DKpmHS4x03SiGa1QSttm39WdZ/bl4WdNdQJRkfUDaxzxxv/yGNuu+JbdTVuR2gY8W/kt6L39Ge6i
G/dVn4RFqHZu7BBZAwFfqZyq764jZbi2Bh1Nd6nVDOjP7TzuL09r0MDLl86xb0zC8lGfspPh8ze3
E/aDuZI5PYdvqWsxgp2cEagfukFK9xFd0ESlrepF3JaryzEpA49xB/UdOoR5r+bc/G2bnbOpnijT
ZiKMByQQYA9maKzdQ6GGwCMhHjn9vsH5PMqPjTvyhZvrr+3wqiLdYRYsVOSd/tZI402K9yTQ4JUN
FVKC/qja5Dh1fpBu/AocGzUe8Da/nmat4Z11+frz1ql8gsUU5Lcga4UEeyHyw3U7A2E0hecuhpcL
bCJVk2nkKc01EwxvKsVjbyh5E9spzozTk1cAvlq4yB6Q/p+YQDSLDxCv3jl1a+xBz6uZ/2jp4XMm
AZVQS2OI72/IOjuGEOT4gOwT7/Fsi3sQSbMuEoNAXKfT37DZRdXMlqeW44+9w+ZfdQryKhSEh7SA
fjQyPGxkNp44n2vBKzGISh4bmInRp0SQsJFuFk8zvoxjgH/mL26SxvFAxizz4NlbeFf2rj1Ey+BZ
iTuOFdnpA9gLDrQEoFDMba8EBuwGzKup9P/IepMASurjj4C/nI62fG5Dxe9JETws1fBiTd2jUNPl
tp4hWf3Wl8jFkAwfrY3FHv4Ak9xHkqUh8MDQaxc6t1wGbYPrRuljmbY3jGlNeSMW7DOBslo587KF
NiL0ByZXNypISUbZml7k/rAbLHEHt35fQt1DCKZA/Tf889HVeDqH4hglr8wdGXrYNqD0P125Lyik
piKFCMSOqIOqkJ5PMoa7Vxpo15Ay7x3P5Dp8R57LmrVKur7f5Oir5+vFS6i7QBlF1rgm14MU9me7
hOmG9s5UdrI5iGuF1Xd5CF1xdNCtRYuk80QQbpB1jE3kT8ANo2WCAePShP9l7TJuNrfBgqa69bLk
wQGNGha4MBuIZ6fSPigzK12VoY9rhSVtfrsfWlswgiNzWNGyoIesqgzAhyLtFT2/V++I7czbyrjN
c+MTEA3UwyZ8+YeE85sO5Eup15FGwIDySYdZDvVnIERtsIOxGgAJ+oYCJvAsaMiPqYd4YuSa2G3B
vgW+GYbamZwv5YIJR+20qENYa9q7D2gLcjrU6WQuWJUvtTJnZXuJwVy6cmaKOnN98MbwVI+wDuAf
qx9um9zsbi1armkS5ogVNfYQCyjaw6ob9H29ckgmLJ5KKiblbHrA6I7SDG8koiM/16AeQPtrnb6I
FZ/p56/fLgijUSKNRpolaE3vpjyweznFMJncPVN2qe32XiEcKc/egb9uTg/hRlhzGn0h5bEqWRpU
7QgvkQ/pSDGZVZjDAIbLHNe4ecYPeG/sm5C08KbMFOZQzqX+Zl1ayEZOUMEMKTSD711G8xh7u6hj
MyURVM7eZ+XgzMz8E9TEa5/T3CZ+IMgbnj/xinRaHtFd4SbvX1qSkeryEjvHUdZn+Cam1KEP4mig
NU0elfBt7iHNbptkW3M6pIVaN+guoD3OD6X2JD7capjNxy4JgOsCPEkHgQHlbYclsvsBtvPiEjvh
DxQWWfpddgX72UZ1UiXu3ECaVrN9P+fgnbFW7zApvnPLgyvazOV2yVLxSnjpYgrZOSX8AOuL04yz
nxRk6ZMT75kAjEVkBBYSlqygw6JSOCGIvIj4y9jySMjZGmJV/qK9llRNgQgd9vo61YeNmHfxv7hQ
UBz3p1WGVgJDYsG2r7dvb3CCFeVRS+sNpcu/QwzA3irdnUcHGG898fQdg4pxq6cUAgl/x+0bVt6n
H+at/AyLBxdbFrYX631d3QBsiTP8UlfIlNYvn6MEW77bz0GloGknY214/TYcpx/74ueiw8j+Qc8N
cSkbJATFqDBYuD49q0nKILFc6E3s1EQzogt/jTQkaevPXpC7y6owTst9tB3UEPjbXT1iw4o6WmhG
ZvBZOmkCYrgvkv6SrdGJMmuicfQNEJ9uoDH1uFZaA5yXJvZuQq4W3bU5wOxCiTjZ1SvHK0Yz8gQ4
9WvY4GPKB0gktzuvGyaHrXiyQsEQ8YYQQBKkol/A8AOF0SYNNGeaEDM6nilNYQZymU5pu6+i/ZxR
a5fnjYVPqB52laBc+KYaW0Ax704583bxc7YYtnoZlGh+cR1wa3g5gVTwi6zrqNLTSIWauVGCJZzo
ch361D7Vv6yaSERUyKIg4eG4/pGZ+oaSpeTVeL2jjPgHiZ6fcm8sf7UvzP4rKiVHm/APINjIZeM+
nqg88dUgFDmd2vz/nGeOnaLwdqJ0CKy3C1zp2RROde0IoJJuA1AI1wBBbWrFDHNpqZbx3Lf0Gsvy
pX2BW1h2xX5hxrVoC8QHnzecGhWvwvPdUKZSL0r9A4DSa1yM8jBXNCXhSBujFiuQK53VOEGH3pkX
BAnDI5pjgaXbuB+4zmWY8a3pjs4+L3z1pU5bCUyyoUcglEgHjDRtiOVsrBSJIC/9hFIPgNC/XhKx
B4xfhU+1kTuS01hvg7lmorbAnHB6/IcIG8hh9FjeQaWxl/6yZ3AEXWpSuwA5cpwbs1oRO5mtUz8L
TW2fTlLGIywlPEE1wxzRuwwxe3s1edZQ3uIeSZ5VOLq/VxL+G0k/oEO/fEgsZpPkA8WOZoxSEGlg
z+wRhat/PIt124OjakJJvhOBGfBQGOG5R04lCkH067NHll9hRBmO/cLE0ENL7tSHXt6aINHb+RmJ
4zFq4IKjJIk30G73waq42se/Z1AxpuJ1AJa70f3KvEIc4tygaqVACLD2vImlsQV7uUii8kmy/+zp
XzDNJMW7S2MwCYG0jsI9a2hfsBQxh5FIBA++quK6E+H9Zd3MOlUWp/owoPQPRE3Iuutadr4pEqTq
86MXMFfcKg2XCV3/+Th3JYGSyymx526Y6WM9Kz/7oUSefQS2K7vaIBhoVCsZIEVKZ6GfukruL9ij
fq2XOv6kICwgri9z2Dl4jm1vH+a4OMmg/eq58RrlXH91GwUO1CL5imaLF65Gq6yVXBvpWvsvs+Xa
zbKCZ2twNBio2ycAle9PrPqj8SPqPtQmV+sKEaoF3116+Q+4KjDrc8Z0tMURCUN0egcH6m+oRe5L
8oulLKdCEt4I/0D7e/nLKKTrCjQEN5nQQJAKYaslDDwjYaVoXYg2vonnXfBywLDQ8M7x8rZbvlJ3
CZlleqpcxF8wJu8pYt5dfcloZtNarzlpX37pi7iLJeNKFvMS62lYqN7SMGhkxiWeFDRj7MfOSmXa
7U3RpkkWOGtTIpLzz2/Uv+jIFZu0bpVYOK5KQgwFalRb24apbSmeNaUfaKh8/iNM+THKPliovNgZ
WCIdiFszX/ZunycOXae6Jd4DNjw5QnXknxiJQUPo0EDAwoowdHGNrnGzq5s57MwtcuAsrrSJuOWn
5E0KdoPihrmkng5xE+4j6gXjZkY7KDHIAWhuK5wtpcUUfrgEn0wo3hnmygNCqyHqe7n1Jg/O2lsx
zBmG24mZN+VoGjcFBwHDQ9ltt4AqUTlkSDPkomdUqtZo78XRSdlbJCGhrDhXPyYqeiGgsyonR+gS
aFIpz5c7O513iypHgU8FnxYuuEEvPeNFNBym4mfxklVJsTvb6e7iC7U++EUGG+fMmxpPApxlaEX0
+jv2wmjj4YsMhsb2LzdypeElxL8EDZ+mjtBRp2aaYd5/VUe/lu+82dT/UwLav82cTE9UXRAC7whK
3ofQbW7dNFfIrbcjXYx2x/GWyMtNlOBIKG+UB8gZ2NzHJR1ZhWqpHVDH8MEq5IONWSDbROTqW7zC
v5EqHtlEaeZzaUt8XsMSJUIplGJ7VNr70L1RNOcV1uXZQ+/AYJ2Rrbo7sTiZWwrn2hk/0YqAnJw+
Gt5nhfpTMWf4edlIeFad3NwRFMUPP/V8we3MFKWcmqg5ud0h8+Qxylff13RexzeXgm44YYLiI1LM
Hr/BvOtsgKmyVPMmF44OpilzLUhT6aWHwY9u2QmaHMADu+rKGuXGMBjskmV0nAlhe1eeOpFQzyCU
odnRKiPPxq5DtnNiVaDyK1lND5EasZquCreHUwoX1kQsQm35bIWJ9y0Xfl1MPtY1HPEOD4NDQObv
yDtAFf8bnBkYdsN/C5r7JWw6bXXvTaYegNCp6zWx9R4Z6sakmQ9RutbelgFXyZudUDpkOGlJ4VSv
27OfVojxNkdn1eMPPFJrKcBH0Q0nE+5Rb4LwhIkWbbpHYLcg63vT7ItiupbhZYSpkD+miI6RPUAm
LBgzyg+b837tvK6GB3vBYbIa1no/y9+3E9NZE4ReWv3g1NQ5HEhHLJpZYhmXP7GBoHK8KOg3gMvQ
sgdEpOAQ/CPGAaIbdMms5v9XKiZR4YbCjPk4tYYbYKuzUrb7J6zJdaMNkfRUjG2FTAX3wyrD950H
6rBDiZOeR0e9N/chB/72QVzD7VlYIDbllbePafl5Rn9EJbL9UmWDX7ugYBBhUrhBP6RM39OHjcDJ
qwJL6izZg1Mz0QQckF1gMdCxCF7Jm+WJZZCfpht0jIVfEdJeVeKtuK2SSAgrgv16tQy6aPwUtgrS
eJjSJEfMbafV4VUiVRHkipNC/Sdl/NBHVISMHxH5kxf4uj2s/nBa83bGtvI54GBZVVragigWJ9JB
EY0XiReuYQxKVvCL+ac0RsC+AcbnxQKokv0BX3+HqkzV30eysNF9UZ8W2m9dKQQyKt9Kxw1puJCf
ZMExLd70Z9wM3GmX9BhsVWLJz6QcWWQRpXmSl1Z+gOAKwqEC4IMewgEMhsKbT9rcx3Tzb8KYYNjs
FfAE3XqxWsmNLbCGLg7EurwgWSLVd4Ye9nhthWZNkPr6/ln20tfCZHwFZqcj0dzKlL+kLPoFYFYr
VzXJM+UYtXf+R4cCjr512hJHYbNSjX75vAX2uXlz2KxM1ZRJ99Etnm7BKcbxYU6KNiivE3/0PAvu
EaqTVx9bfHMJcL3a5k4f/8oL9rwzIB5kJuK7RhmpO35rTO4/r9Vvf3UZiZfP1alnvruqNJrwuMG4
n1MbnHdV6SNlBb9eGIOEqIMKPtM0YhFCVwKUi4HVF/5afAhdowM5f0BA8b6fi490x8oEb76r4kKV
luBqlJgvb9bpabP7+DUEWpEQjj7ZyBe3+ipoWRm3USjjMx+jnzRK0gN4qDDrfxz0nkOxsOdS1R15
GzrYknTeZR9wx5Hfvvp0D0fxoyMuw70wgEAgCmU7Yh0wceKMQLF4x18GfsN6PU7YQbQAsCiQjXNy
f9e7dDbSSpt/8ZKntRQy4gOLBYseSD0LPGf4QDLUzMuGSJHJz1Q1Nl85RB/wQp1g+PVm6SzO6PYO
ehtajy5t4ug95J6nneB45oNGmOj1eA+gB/bgnKbHlysyLSzgit1Kr2XNz0WsCJjqfp+JRR3xCZ+s
5jV8ZevniLeTrL0d84xyXX5NAjzH9wHDO5Y/7vlW0XfDcS9RXZ9DgF7TlDvaaUxjYqwGEuZBmmYg
70jbMctXnt0A5kGbzfTIS1ZJlL9/FcSH/rWvHB5lFHJyv71my9oPZ3h17P0j1Ivs6bYRUbTZdgh7
77LVTA2QAaZwQZ6IBwEpzUZ94O/R3ELZ6HhVRf3YsgKemOYKoBNk2dTCibkNAoYOvXj7xTQfgR+G
VcMxA9/T64Pch5FNG1ybJ4buunTLONyMn6/7fklbEL5pKxrehcIVWedxaG0ZSG1Wg9nXV9LbUi/q
gNrkrxuPNaS6YAidqOs7rjVjQiwGte6fjxheNyL6jLUWTRcddWmBSttsV5fFtsPmOVD0M2GQlAVT
BPlRb1SADOm5yRRStTtg1SFmGVCed3vvC/NMy3C3JSUK6tiDMeOi/VG95YSlYeHVt5wOfyQdwxUS
yrxgI58lTvB2EEBkhyC5H+8dnCTm0GdAZLf4+YnYiVBJCxkO1McS4k0USDh7EP9pzuRW2Xp+V5vv
2LuvJG7oDpXmI1khCC6KZsSSfrIPXi2Ud92ukAvxFGREixnzGXC+Iuwrhni3Th2q7bETFxnYkiUE
D+Lw6hfRAGKo76wy2GG6HfTU8PSsyULGC2J8qY9UZyQYPQu5OCy+d/IfQZvWShjuWI+znKNAfEFa
WQfEHeeFBdWX46aEb+jT/NxEhJXdUTXam2g5A1rUZZoUlASvFVUkiLLQc61nqs7VzCzxqKgLCK0c
PTtJW5VXFltD3J9ZSOCw6INycEp4q97pBYJgJdrsG/VG4QIu5VU41AkMqjvGHqBZYiXufJpAZ6BD
9KRrUHY0hf1ZY/krLxJC48fxf849uoRefw9nFi1xEyLUbwCmKe+vCQb0inH0OyIkooRKkjb7JXlo
rMaN2QtB/SDZac6GkmcxGxfmnhWe4SUocGTKOnDEq+vyr8sxRieCW6GwKWZCK2cJ6QJNNXvhQhuJ
HQgUL6d+S/+0OSR29JdT0PHEofC/FuQL0LZvZ9Tg3GTHf8fxc/oOB4AFcHDQv0B6kdxhHxOYMwmF
fOBV/d0stRFW6C/uA7J7depbd5HoppGJ7NkReXVk+vy+Xh2B5+Q+22HW/CGPAGC9lK1Zk+lrRg7Y
dagd6dECPnw/qvYyibttVDyT6ASor5pzYUiz4ztDQ4MVrs1W5bXyATDPWuBfIufe/x9ThJuIGhm6
rdngCwpkLYg/FCXpRJifX1Iy4HGWEiwM5hS0CgPw0fqxuUosNfOeDwAx3/us/47XIFIasQLmMpCG
ZF8K9RutsTDGorwT6MBRQtnS67z8s3ZK+geMdNVm2fEWKoKNkat0KCFwAtafHxZVxho0HPNeA7ah
/WHBp8IisT5Vjfk0jm2G/WmVtM3mcFvkDaIklII6e46xwZLGST3V+iHfJKH0xQFb7UsORdWssa8b
XTlx6MGjnJTbgpsP1nAd4LMAnhU+YsERmdOvijMqsZ/HkDxR/9xjRPIYmjdRBMxdiSXFyjj0gzxa
ihcEuldzehG4nIUHOtd0d1f4rPFswX2EwiJk88XzTMvma3wHX8j57okzlvKZjZsgXHBzyItn7bfP
nIcPPf44MTHCG+9KdhN+qk7xvBS+kzUoBCJIxESDz9DkDzYHh0iE8BMv05D/1V20JghzbLpMJW1P
yZxpm6rKrzypYYPwvCujRYzrqYXvLS35aVzBCc+JPD1zwZy8VVanFLGxKiDK2ycKct3vpZ6N4NvG
gK00O6y24erNrNKSJX+EI7rf0KGt7kVr4ikp58/YFroMzosXDhvm2Eanfy/wEf4qZLelqbLx0QGq
mGIffWBUuAxDsDXjQELUJO8Vz50p64V+lM+hgmCnO23B5eTJ+szupfbdg/1l1BtZdJrfLBLmGpR3
ox5RuDJbn915LrOj8fMTwAh+WsI5vhqYxpkG4L/6JDSNr6b1807yq2/LZ9dWqNfrkmB2W0twQTj+
sB9cBRWZz7zbcDZp/x6nYgiOtcDLVpKe4zbs5D2o/2o8pYARMuxAYg5Sl0N65k9FOdm/ES5VHAwy
MZVdRVnsZZkXIu+C6ljLPF2b4ca1aXx4/uMcu2baZftXHqaeeE/KHz9hq99OtUKBEgUGItbjvyux
QkjRPLA4hbjQweHsQjnIqfL1OfQ58jtwXOmGE9NgrUBONkAxgXE2pTozF1s5NLqGKJVQRuqz6H1p
qrq81jMMDkJrXDtdy95hkbmqQqBjR8H0RrMNY6AACDydedF3w2vALQq+EwwSA0/ZFL3ryq+KYco8
2JALOSjbTT/Ynr84eBrtI30pKK4itpyDHIBVtv7vcHfpi4c/xqLxEbRzTfFkjgdXRfgNyJVoD7qe
3cputXhpTq5bgVkicO9limbPGB7kJNzvBMOLaezXvA8ADnpCa/Su/CUFC9biWkdSEd8EotnV6AAL
Llwi3+jvSR9ih9aifpE+nN8dqckg4QrcXbmGl+LeqcMS8R48yRI5AxHvpYTlor180f9RClPA4iG4
RqaRl0LT2qCC4JEcW/LE+gaWNZq8wbs4LdR2bpUV0rrwYP7E6+QB79te39OcAAE9/NBocF3qO5fd
NtHYETzvbwX64CcMs9I9qh3EE44mhNOmkPvKY0Hys1YEXIlTcUoNuYz6xAJbxJXNAKCLRIozXxk3
NT+OmzMtJCx7qImPF+QpD3TI2m6fAvWoYU1Mlr/HhW3TTi9rfZscpyoJwSmRP4y+jZFVD+3e7d4z
NBGSBfilpDcBd7bLwHS/arQ3ZuJUwkGeKlT4v3F+G4E5ucCj6iZLIHWqyuflAfRz3TIDOuNmzGf6
Bb86IfkqMw7OM+vDP/LMLn4+N7uYxZOyltqnz2TxHiy3ZGqTqJhvoF5gTSsmzkhZXZMi1SIyseQi
bbjdGSoaHjvm3anO4OPZjQaZlf9in2DL+aTSFlDFoywB9rRBKvCRLgF0eKBIOZ2/ilt1bKnqaCDM
+mCqYPdOvGjk7Bita+yss04aCqqrryVzhvv18WUEwvRrrqF5N4OUPtcXTi+wnh44pL6DB7Ph7RSb
eVdMMjOmO3bGbdAvOPB5ZNl5KO4QpoWh3U/BNWwlHDwMCZmPSvae67+tmQ3ZDyVygD83ax7Ui73B
x358bzPM383OXzehUqSI9fRDC1z9mCwWVVXeRumrRKO+6K3n92akVGW8EikZeKJoPrE7H/lML5xS
7tWDHap9uNCNUT+ypdkjCYntl4oxK3liQzBGR+531VktMZWROdAPySeT8/cGvDH2F/b/idM1YrUl
acSp5R5KdHUTQCZx5kIZoOuL7+0L3sqzzj6VmGgIvdBR9aIatA5fLT63Y8lQobS8Ao3FrxeiuNS6
kMZbGSzPq00+JA9URFZt4gXtU3W4uzLciWs1Hr36uakPvaKX2Ll1Y4xnN1dX1XPJYfRPN5ghpaZz
8odLKRybQKmBxUTgBMnfy87dbZXHV/X1DMtqJKN3AJ6USS+Abz1QRCWKioGZU1lhOfxTmB0dnLg0
km6ErGt6RPGkKlppoYHsTftbKi/Q3KnZ3jw5xrVJ0APq7Vp/CMG3FA+E4Mm2K1bcfpdifJylciuH
ou7fI/LDylgBk9mqAThTxxcKDgkuwEPQSa7wTjfpkmXl/rHfAAW+EIP5oJuZyVur0TzsaJRX66DO
y0+O1BqrnfNhSPTRhWkL4a7vvjbgOBGTBSv7cZ4/+ulIMoU+az2+m+463ovV5B5uo0G9CwtVtE81
DyCWjegrgUpsCmyUluwITgAg8kgsPwtqgpKVd0KzbmRMP/+XNdTmKcvmMZPv8E8muOOo5aP/HR4e
B1FBQ2uD2n3EyQuBuLuxrvIdH2fTswG25BxDWFZK/dqzCr5vXfEidEX7FNjXaXJ+vpgQuZcKD0gN
T53kLyeiM9/vfr7H2pQTS8Agw8wu/R+Dy/4okGJ4CJB4Gt0bdcPtejXNRPRySJFBFoIt1AaBCUvq
oM2WZ4NkZIku1AmVwqHZo66xMT3XfIajV/iAcNO110wXXbqlYecXPeEusJODzcLsTQLOFmA1+7wd
PM3jEgQETP0LIMWlsr+hgYsQ5qetZrGyIwxhrfB1biFF487qWxgCh0gBrGTW2kDLt2XOJlNXIIG/
svUPpHwrC1o40+LodmFmkkuLusFNHsYDoKYYWiu3XpZGpzXqz2DWrXxaIXQtloIY8Q/EnXaWySLa
SL+i0zoT6dTZp2bHMyh9hZX2Gut6oCuh08XfgkHiHeNHif1KU/5DGLEY0kVTYD+TToW5OdYKVodC
yd8CNE4s9GVj5sgNJdc47dnAR25v51a041HnjPY2XuqaV42+n3Q7ff9QnKGqF0VD5k4dIPNWlzNo
vxDDpJvcVhSNEZNuZywoPr7AEYbir4Jcf45XQXOt0pC58qh1Q57AwPUcc2MRdpHYrkkZXnPX1EHn
iZ3UTtC7ImZk2t1zQsIv8zgizfG8q/MApdCtUS19XjEupDD6zA6B1W15KCxBf7+KgRK8O3xfnljS
HJIBAJB4DK7UNosw5A6rU9WCqdPvzuLvDDnVK8EulbfZPoGt9zbWA7DW8to9KqaTgVJOFGY1EX0l
e275zcd1l8ZVdYWCX0ywOfZa7mpypz29oZs4gLgXWSV2+yEVzy236JYacND+7cSMsB/ChlvQZtOD
mNf2OnfNcqnLIma8p5R6YlSiYu2XD9ht4bhCCXaJVehEV4YO6nk8+U4ZBhRQmaLqyBr953BaLvMD
Rk7pn+qlKbQmIxKBqk2/FR17MNNRZBvwmlvgBtk1YOCpwpNNQD0HEACXeJ0Od5il3uYI8hAbwfPm
PeCTpohptgL/f3JCuN/0dE8Ao2ebBLiIs2YCpfmURoU+FT45OvCHG+YX0hluaDeXTl6clKYssTFw
tuPavUv23b2xksYLPR6AO6Q48evwbsEkqpiDERkaaRAZB8ubdZYFJevEjqdKSP9QygXbK90jiiZR
QTZy2v4s2akuv1YVWLA4t/PeFL4qDJ2qxTVEiE3xdfNl7hEJ1EWGzSvc4Iy/1UXkMA5olxJvVf4q
3rBUTV4pPjtIJAMChrHO/l0RVa0sr0x5CWi1jqCcP9PL2CbQvML375EAjNyUFGR402oecTEaSyj2
iL03WTwlmNpXabmzer4FHo/RH5OWrdWRT3Avz5xO3mYATDAwR6NWOPtIQnFfjuWe7BWUu3i6gTfT
xxX5HiKdMSko8nP1p0GRAxW3d7nbyJt4mFcsK6B4xQTgspVX0vFXCzOWtl1esGOGXSu8tsCh+klo
xf9e/PLHih5AWrUROw5zhb/A4doasMJfGxKvLXSN0Bcz+dN6Yh52MX8JVXS6rrIgFO1ye3gnUI3K
+V1luPUBywEMbZ5ddirJ0cljCUuB/pcJO5ywXSakUIAhnh4ktDb5Blwz/mvfPCwPU7ABPCkBDYlH
WYiq0G55f392l3jGA2bFKAQCAcz9jo4QUiWCTB85mAgAJGPSZ4H49+uJSKRQtpiPTjbJVFBZ8Yvi
V7KRjoIflucxKlvHT6DiZhSidZFIVMlxsQVceXpvAfEtWdwH2CWXuTukOr/joG4VzF1Dt00Wck4q
CDfREEQt1Qa0YkcEcK43AHJuccgeBmVgpyfBuCrlUlViXt2GELfwoQjSPT2lVhWljp2G795T4rBa
UPKqYpWM5pDZRFWDbXC+5dqj4ApQtd6Et5lNanignJpRTHcLEMNlHWmvXrNr3PseYDbNFj5mR76G
qDp14D1hFtywoXn54ie76h+Q+AacyoLlgtSnspKl5hA38MjVke86sQekCrZMWfAzN3kIACb86hsg
L1pOjJCRpxMiYVvjnv8ItekExQDC4lTHhp1TN9rMDhNs3whcm7b17P9mmsHfQv4lFNEwBAfkaf9/
XUI4Z1Cc0Mb4IONu91JxAeyTelvbsqELrWzUrZC9VuAll6VeG73Ei9XVhK2cEP4jgfT2DGS3UtWZ
kwOjwcdYqnmGhqedy+FScKG/1I4vY5tGGbUZ4RfOz4Ne3bIQxlWSCF3tV1VMDoVifBTStITiDW6b
/i/xYCQM6QWhPWEZLt72eqQSdVB1HdS8mGIsJMAHlOHcYO2r7YB+C1hCXJ6uSjd5O5yl9jVoHM5b
4qUlD5L21FxiOoskTL7iDR0/d8lNG/W/wpraJZULmAstsUb4RSY2rZZvmdczzCTSbV/jBNo3h5cy
rsGfZRKpiwxrUBHIQR9AvnNkZkt0BmzJX43fbf5n4mR6cLo8lFW4GX14UY6MJNhMg0pGUP6Pd/wt
GxXjSwetf1Dn1aMxkJHa0BgqtH6NinKblzTsj0jWxrp4uKYndqwzRP8d7sjfq9sJS0JRpuwQSjra
LXyRCUYotBHLQfNf5I3Qy6JpLUv8EcvXqFAVecqbvd/C/QlFnIdt+I+SLE7LlCgR3ojWNB76/v5S
aj4WZ6t0nYEKIJwBveFTv7AmuHp7Onc7lkOt7Dwh8Vz+QqeLvLNdqVx2UVld83Jw9FQwyYydebnq
GT7i53C5U5ZuvWPaYHbLUnWMXUybiopAueCbdiXCNrcV3jDp7+u/LzxJ4Njt0l9G1Mdft4jcfgyy
wZhf2dEcUmAbi/gw5rmbjfZJaG5Ae8DDO6Uc18vZuGPMO0dHAdr9sViMdKL4JVV84Psg6y1h2tcw
r0S0z9PUGjqm8CAIumAE10TeSIAnzauqNO4K4IE50phdHDRxWO/w8VAlLdXiZYLdAS1NihcYsbtY
lzccuMHq+V4gYmTPSp639tSxULXOsVgWArT4h+EJnzR92IMtmoEbqarSiNr4pU/1C3s7cIdUiqiG
KQyQ+7EVqaNmskTdZw3kofnG7QoV/3uNXGuoLhSORHN2QwSLUA2v5whRHv7AhapKeLX9dTkNKCCB
2TU8ts/wf+U1LGgfVNZXZkMsDJKtyO32K8LFzLHYJdHZZZZXFsO60ayTo28lTrfANLHrwwNkY4DR
FH3u7UYaXnhGZpaiLH377RuLmjI+jEtVgU5ODwQslQ2zpUCAf5ExXeENynkLlJJf3/oUUbvAAM4f
vwE/7La/9S9BFG5HypOOO/Z66WfNKDsn3te2nCE9TGow2QkYqYT03fG2JK7J+wa46Vr2ZsbgL4oy
dztE5AYcEjuutsTbsBZ/Vi5OZVZGc2Sq0Rtosk8hSuDee86ewCJ5PzhggkqEYVvgC5tUaAV2Krzf
YJ4LbrJATkjL5HmKjIhWXGh8YHjxQY3/2v9O3k/WvvfFfYYltH0SMcyGpSN8ZLrQ2a1lHPy4oo/s
ZD0BUZl5zqrXPIzmCcb0nUPXNkSw63AEIHe/uYrx35mN6PUBOqq6M6hkaPvMVzyfbryGLUwpPKIP
0s3zcG9SfIEmp7M17kBtksaAhCOC10RrxkTnzfODRcHZN+Dt3bEpKSLiCtW4JkgLem4qwYhyzIjF
jOvOXN20tc/s/hsntFfnomlHNR111+PEtd/FMvMTDG1AYtfoWWhJNlWDH2WRqdXg9ClE1SePv9w6
EGUm264R2Lfl/7WRHF1qe+dYpR+7D5PGmvgsQJyuMlSDlmj5z5egexT9aCZIv4faXxSas+5PLRRh
2omMZZvhD+4WLsRugeiXvCEENR6l3Gzgt/xnJ4WV9haLutaaRAYd8tmGGsdrDyBhcCmuXNmY6egR
jmkaScPm368gAJma39boPzlULnUnRXVOJ8xMzDzkw/Y7hhuVjTnJhDjgWuuLJ+xfxT45p4m9gBG1
k94x5BrnJeSGI4lWTIBqy/RpHiDKb7F68DgLm8lg28bedEbBXUS/JDfpTlWJe3KTfA2sMmhczanl
bxpaIS8ywkuu2m+4t6ACG0hcsyZLN7QM4mdV1zOhqGX8zfuKWgvaUiKt4dzMBK4ZC8TJSILrSl/+
uh83VSqODFONHPGqiDMlp1T280vL2Th5mHL5UofLy15oERMNW9IpoZkYGS1WpHavNjQ39omdBZ3K
ldT+vaH47CAKsk/AVBaL7fjbb7+MSoZdxrxdLX+7kqt3xNkdAk70MkTFud5CCGsf+p9N6z1HGvpw
AU+5CWPPoN9quNWRyoqltnubxfrLD6sUzkF17OAEqmJ8tcRlpk2D1/BqqqVPYR5QKFCnysyTfZtm
u52Kb2x2k3jWTgXjQfUB3/CnfLe+lFgLglDWRacLdmiJQrCQuzKUInjCKIV1SsVnOb220CTWgfcQ
C/wZQTZu10qBaqYQ44Y1OUfepn2jsfhpVSNakOuzf4tkm9ZQnnu5aVtxTsQnBRILhHZRIyvgaYLh
CneSfqBCulW7f2i02FX6d78uW5yA3Re+38ZI0VQO+qmWv0Ctp5bDwd367XHHsYDf1Wyqpvw9YTzr
Y52s8rudhUSGiL3l1RXy9peN+yzHmQ3GNzyxaaIvnreL8kvPMLXrrTLO97AvCY1y2WJQA19zknk2
mRqGWgxpHkmw7P/7CkjZkD37JS5eVlAkKGK20EU5/bFSZ1DhFGFK8rM5N/wC/v3ZpBCwZ4WF5mBX
ffQadIJdKSIP/Rm6QqWnccmZm1mqnLdHE+Rs0nmvj5/6Jkf3qWPg8lVdFZy/+DpjIiFT54XDhwku
ovBQyD7dWi13QPggfmkmV15lItyeLs6BMvcjbX5a9FSDHGaMN4y2AXVzo8/WjnRFzwdpQfJGdILd
W2H4s5v5wWSfZvp+hr58rdTxXns434aQuMMp5Udw2AeLJ0mmWAvuL8iiaBYxF3OnLSqBLUikmRca
MMVr6RJ5GWS9uyfBgMk2njX5lYvvMUbjqw0o1xZzTBc1YcKfl6peHC+ri4v6ogzlxpNgJCqTRSN/
0BQ5HU46VxZuqrpskanmeMe5BpQb+LfesAxunrkZL0GgGpkmNQ2zRd/tFc76jGEFoEs8nQQg9dng
uPOdPdjRx0pzM8GBlRvyZU4F7m2YvZFVzTpIdRfTbc6SBhxQtBqIdnQcFZMAWH+GHpErEOffz0vF
j46fbNsl/Anydif/suXs728ZxlyQ5aGddaBAC1LDAhzGRWQ/ZaWVRAE4VaUeEFamWcdn8zuxNtBh
/0HBpt2IZntlDvxeehEeAHMadbnYrc7qZyWPy+bGyqNoG5vEBVbDx78pNx7U78CIkHrCtExxECu1
jpEvT/GclhPY08kDwj/quOxsDmepfI92ZdtjyyR+FbgzEUDDgT9NyhQnDeJWiB/INT/qZKqQRc7r
/GqvnTNRTS4V9YZGNlen/kQ9ed2mqb3eM8Ihyqt06sjBuT6K46hEZJWuoSf0V+jTtUqZj68ZxETA
/r8SI3WdB8IR/cv3s8fPQ9D4UWQQt8q5c+94szCnbfbbbQkFdTv1KsRaZwjlRPdAIOBoApQf0IP8
rnN+FB9FxyBfhiPanibgDbyqrfiCDDeLcLoEyue0hMIXo2bqsuGvOGB/g+hf9lFPMfKlxweCx83g
MF6WEeqEgSo108ggONLmhB0TzyZafSMIIoTreUDpVO/bBfpmNBJT/FXdFz3x/Oj/dY1aKRyloKjD
7Gw7LDEV8muQYYO4RHtII9DKXaDeNeisu/ROF9mHC5qOG8JP7APeqz/WIY6Xc1SfQ/q5/WYqU/bg
dLe2kJtbQoEMn/DjDQ1BnNyDhz7EJ4tcRI2vPvUsZNDT5FWG82Le9F4Q1KAD12Kj+1NWjzpDZfe6
gEcF7j1vHhGF2vZ5wZY/3lMAnxqQXhpOyYOK6vRBtFh+so3sTlM9mNHMV2HHiS+WvgWvgoYc7UFY
tI1OfxkUBk23CCJgPVwzE1UmwP8XgpfRrXyUSgsRphV7c3LY+gpnveThnyxgWn+FWyRu9kiXOBo5
ycT28SKvxfxDbHEzEQ7P1tMafZI+ZJZKF/Q/ZeeHYlfouaAOLg3H++vLqFAMhaCPr4VFzwINq1O9
CYlBQ9GSB/Kr8uChb+OoeIZCznf7fMg7/Uj3yV3oFb82AgH0eJgHEn1+n8+4kkCbICtarUbw6X5l
rxlXTCVoL4zvuAXpuV5yEJPR5qbY+8b2pJ01FBgg+AjN2N3MAvsKFas+AiuaAQykOb+GuoOdPMRf
hUmwKhWSaqvErPfhK9OeDyaPfe7dSxgT6Ow1aXTMujGXOuGbylCeGEqZrcuPZhuJiZJmTxINVM/n
+zJjLpNzUuI3IxJps0Fe/Rr1mC+dMU19xb36VoUkwVu3QwCNW4e2MW8hHH7WAA1NqRz5OflxEUdA
SYAGaimmax5X6hI9xRDxHFAhOqXoCz8DoNtEGgZ3g0epI80kejKoEabBoqrIchuHTaJHuu/CDnzm
+LKQoYDHJ1W5UivdOXHqttgXb5rtn+GgJvwxIpAl8Sr0+vcR6n6IrBTQ39kCjUtkc7hq22fI7VpN
g1tzD+7cQ5yFqLAi7Xvh1xuqW7vXoObAgTvdVw1eBxbT06jkTa4uak7Q1EnCf1LT69RfpNE+CDKy
+XJNr+JUBG3NRrVLQ+1tAgZKeTD53DlhvS3u7KIIG/abINzgzIj71AFGD1HfCnvrngH6jeFUAD/v
hULq0ou/UjMrh+B0G2C1eXvLttDzkZczMdeMue2b9YL/B6ys4hmVlDmxq/wBW+aAfOhl9BQhl+gn
hYhceDseQnXx/IuZOe9hLRSlWCRhvI4rWHjZ0rYDhrulYz5YLbT/cB12oQ09jkKaBm+ehoCZs8wI
RouC1vW9/cRk2KR7Un1jQ2nsLGtYTkx8C4svdQGTZ3ojT62F9vS06YF+h9M/YvZQqAjIn1RO/938
Y5HuxoYL/Hk0u0Cdw9u4dKGOfWlyvFQmzFYAO3z4Y9WxXygMxFeZCY3bb/WlT3zd+LWuSL1JyQUl
MjmmnpW2u0U6V19B6mY2ggzdcYAELfktaZE/YjugYGxLMSF6No/feF6IagCbBnJAxVeMnLtbUyco
vsO9W4U9ZEfRbMYYbemGWBUjLOHtJ1KBl1+xO2rDP6AOPBKw2U5owDtchbNYcAYLRr2+AKBBF7GV
Akek+Qb8rv8RSJ2/wOoLNehE0j1I5UUoxPVdkM2BCiJX9k7KMrkyzY6dp7pt90cdsoqHpWHhk1de
fEyQ/HHkEXEI5i8Q2R2KWAoP1Ry69H9uKYBBQUOxYHkc4JRxby//YLEYOsVv2kpPd8f1Lnj6pO0N
EchhnURqO1n8jnhRuI19Hx5/pG3/YNprdBPmceqDFDegrN+/Eu8cUofYQZVFfOWeIZNAXUTfXtVJ
So8pUeH4bf218FH4K2hSdAuNCOmXYzzSPwksh/+5n4OZMQuMxlcJNEysl0ECs2tOpTHj5E8RRyVA
9u3SiC+ce7YT47JW6/qeytS2fMKl1iU1v8W+chusyfpXwUgv2TWX+DNyrurmP3IBEzPi8n6WRAPa
FyrENl/65ix8VaBwREHvzRU2/X6hOrmk3M3CLMWX0UmofgzRNlOrH6Gu1Z8BOtYYWS36caa0SKiX
rpw/J4z2z+vlrVX0TfPlVLqZc/a4OQYcIT2VoUsx3ztJCcuZ/vMGFVypH1U/IUJNdE8jqZlxSeka
9Ap1H02R9LolLL+x9JBTKVv9ZOa1GRxB95SYJfBymow7L/4LkaBYFRRJ0mqJ+HgontwjmOWPXL9y
2OP/ukIg1RhqfRgPSmXK/6FqqeWykyv2NM0Awzc8FEdYmdTV4KBKHEvAF/tO4kvDsVrhsUSbPAvn
iq96g1UZ51ZyGia5Rot3f+BcllRK28tu4uuhmP89ZeaaBf+3ts4ju8hmYivN/gzPxSosiVlcpyAq
nDixr8nzv6Bmooiz+jcBIXr+9oaaKfQDtwTRlstnycgpzsDNwlaxQGpB5ElBLi4hseCnBGdTE2da
R+SWUdOjSJraO4nl9SCFFNrPjqKKVLBmnsiE54Kx7IkEzKPwnQ4irnWohQoE2kI3wbTmRmaerada
rWp8AccA6l7ejoSgVe04CtU7WUsG300j6NLgWaMHpnmNZl1WChPnN26aNkR5WUgfHZLuIqIIsjYz
N+eJ4JOlkD0ogRIoVg/51fvWbhnfwV9ErqtW+6be1Tqn/11Oi5cO8jjBjv/ihD/J73qWcKZYY6S3
K2VkWrsfF0hXvUajBTuI0U7tRvVfbTO0fenI9BZylSb5kaglrW11+vFRYc8MMxy1D42tb9wQyNJC
R40SqbPDxw+QhPBeNX83hdvJuZjwLTjAEuSDvsYzajjyPhFRMOqn14CBxAS82YVC4ZGoYY98Jm43
8jAcilR2L/LH+8mV9SiNqXktCnkDdBabHar6QCe/ODZQ0cC3hORP5FD7GY9m97srPdkOpGAfUQpz
1T8RcqKqI0TvhmEBvOSpeB7d3bWS7yXDL76AnUev9kHEBolmTp265rfl9E3Lxk2lKtHdMWELwNUE
iIKWCKmIRU+ChEmYuJbnM/H07+AtReKAHh75RzNKUFZmlZhc0+6vaScdDU1Trvg09ykqlhnmwqlD
sK126fThmbpY7csCo7i8q5E9G7y/qGnntFNObtasFkTZqpqP32gsLf79QVXlx22ex5kDjbgOA/8T
8swD2qzGEM383UAhKDtW1snLwOyqIMASizwH8YIZ/lmeKMpGN4HhtcxFNFY04iolxBuMfNhJ1P1h
Nj85OzOjxYBjw4jMfBuUntPwEof+AwVZ8vwZoiWvD0O1oM6D7V2OyhgdbR6oNnptm4CWXlsA0F2i
CXz6tAmAl8OGtfaq28nRILeBg78scP5kgg0cYeqFL1C+VI48m2WpmeU2cd2QtDom8uafut8nClXY
YG/eirvNw/3iy7kU8ardJACziivr0T+tLTS1enF6WoiLOB7ed0tglfgXI17m02WaVS0gQxbOzfCt
4areWgX8gfxaTXkLmVjbCpKEJmffS547Q1xckvDXU3zQFEQM4pEHkmkAHq5uipGPvhN3ktLeuyXr
GWHWZBdEQJ2yRxjIOWhxr2/GyhWlXjw7IZ0doQwLR9UkJRkx+4iQp2sJNl/QO11wsAum9Pu+szoo
C29+kBlCYvS1hBMEe3IVV61tnY0wudWIPahHVTwDTA/GAlYOWeSQz8JSuFTaHpBipfSp7FPaMBQP
MzaTBCjfjdKX3cdObV2Y7bVZ5suEy2DWs2UOgNXWAPaTXdMTYqvc7d7Hf1AnPfHI5F5Y1bWqngr8
1fVcgbuDNLLId1WNpsV/6LI2LLGbRaruefzjqjLM8/YTHdbR8Hq0GSftHX/0p5rAkxATlm4h7Wnd
EyeqUFycjlXIAbNYODOy659GI8szyEDJKXiX8m+kbbIScQAiME//c4jYcArm0yHki0ZULcJzK+Vd
o1D136bFes/jXBAAuuIxH42EuRhbygYYwqPuZI22Bp3fXqnqYWUkWFxdlZCx36I6QY6MPiHlkr/F
3cZMgLbMNhM63874Ab4VsCK59Zc9JQrjeyj0RVxbbsDJOrUfR0Y1Fqdd+Ie9RTpnk5dcCrmJlIol
Dd2b1stN4u/ISP1IoT+2Z4eejeRb5/NTLr1Y2ZFC7agFLkp8kZ/AI+x7zuh0HAlfd/fHk3P9OlX0
QiKQOGsCHG5v4Gg8syOYSpsQhR5KQxsOa6wWxmbGoiP8EOc6brxL5UMePSawruVL4tkT1DmQASO/
WnhPz7MbQtdm3wHzfYLpWCNPJWqBDEva6nlNNn6OSwO8wh05C3/G8afLqIo2BqvTgE1P+qWYUa4W
IYdpLP2y4IlN25Aybt4SZ8EFq6gbgoSGhdXJpfEqldjEVK2hs39oo3yY/JPLnh5HvEhZRavttdTh
47wFT4EmHEJGbagGpUFbDKlmca1PQ2dOICXCl1wzj01715e1O1JgO5VvfFnNXWOZMCoOWwPi2N1I
0rdQIOgDteF5ywcnLgOow3YW8Rdtaj2HvuDUVsO94h/VCClZ3A24kol28/aeLvRZQuw50BGqx/GL
aaSDbYEMzqE8PNR0QoWQmvIVMirhNloVP1ZzKFMrYewU3lxGzNf5l8R4hYtzP5j5cHZcDCf87cOW
jFM3boh35I1Y4iO/xWAJ5L23qxvBNNGrpmPM6zT4aUJMNJLOqyi84ZXvovfEc99VWxlYSkcySe3L
GjfwypYkZ4N5dvX8GmKGaczUNjUnzjcK3KpsuUeDB+MiWU+Q+ZlPZjdZnwwpiKX+buQS9ToPmL1G
gqF1zq2IcoxxBIEqGLkgZnWJz15lsjH29yKgRUMWvDYzCADyXmqTsJdlUgzzPxs1avcUwJivv4n7
pGBJnvgp41u9p51If9jOg+gWwV4cmDoo27rVSklRyDIEOCeFpVpai+AVKNkGVdIMG0Amrj56v0gv
7VtVKrxDpOiIG11wTHRoAiXQwpkOh9QbfFepwgfCHc6z1HZjoCzkeATmLQ5DoQ89TmZCaz64tgtM
ULiOX2awdJd+r4pjXCMtO/zRofO/DfOJeb6cSoo0bPre6EihUkHsb9ELoH6QAxW1yYmPKXKxLMei
wZSFzGV1zvwOONxB9I3b9uvZL9zGEguVXizCbx2N0cpH9WvjPRqWlRnObXwiPxX9iG4ceBmX4EoY
FfihkidpBWCfRYjqKuZ7CVtzfSrgIGMRseBP16h15/BGtMFLUhVm1SiQC31tbEXBS6nTghm7fuDm
VwkgSs5f+evukCrk2moE/h5KExhqAaMXKxXIK/QVSd2McXNf5q1CKwXPrmS4+3IfyhTQBxYK63Ej
4/YM2R50qPCwtavxQRSGMAEvRlE3iiuGcZPoHn1BAhyYb0CN0QAxMrOEF/NiWkiMUN+VJTklCfnT
nOkwEh22q+sg4dmd9UH5Q+MUZ7qkMzKNLWVbH26gEtZL5H4xJ5WcKhniDNmFrwbweqRkFe/77C11
BTBtELzDKfDEGQHOHSnEqBo3uptHlJDAeC/C7hQM7wnQzPoMgNOqExPqNDV+ivRZefS92t3EzgoM
VlvtlDL5bbxVxlw3dBXaie3Gt/auqLlLyuPVSdiJyBwTBbIw5nzCIcExZv3prdh335W535t/ic3Q
h0N9oytOtYCo+TlJlX4QCy1JKlgd01A8+HEEhQQl4QKl4Y5hr/STRrlo2uPDA/Zuni6rqrzJl/0+
zlobGlROMKGYcl0kWFtMdb7gVzrz7IJ/xG+xiPWXjXWKWZQ9aFatfSHtvhChicFOGyOSTbLbH7td
ACDvwBIPYX7TdyNWf+SjFW1FRH2hTQLAGYORF9AS2fp9et5VS2ByONkmQG8u3MfveTesU5kfx68k
1GPKVO/rbdrFrERckjdfLaDpqBd3CkkPl2WU0EEu4Md+PBQaA7n6+6wg9qskKcK4ws97Z6tSqyh1
a/IfGnsSO+217pKGS50F5URfBox8CeeoeXqJtJavl94cveQt+gXMCsCXa0DX81hymoWARmfDBUN1
qR9mqduWRPzKLYjj2gjQcZWjj2KF7rNlRRFTx8d8RYEHgM7bg+CyYjFRLPw0bz+yGp8rjn5KHiKy
TbRKOJPPiTB+RsfbN8YS+5TtGa/uvRXB/bFgr469GOV6L/V1Rmvj9weAuHYbYwFKPBc2W4LZwoKt
e0kWCmPq8pjlSae8ggT2WbQHEPqBXwfryeWQU6IcWb1qhVk9CYcNXP2pBbOTzXUiePN+52usf+6a
Gr3gONLehkkefvOPyaEZyNGFZArmDBvsKh+YrBBXIkiDXqDKJj9mMCptvoCHHE3cAPiql8qtA1el
2qznuNRe8KvlFM/EGQki1mR2wX01FAs6sDA5Mn492xWc/kCciwTGLGNM1Yx2brtyZrO8H5GBBwt0
q4VJiwXHwrDX6Mt8AOmgIupAi+T+okkbehyxPObhdCZADnnqNKmCubYjUX3kIGE10P5YJMgWX4pq
FiiC0/MxHm1k4tZEBzHYvjE6AlwkJdj+hyusw2JcIGtVyjgecepgDHrTL2UkqZySRj9xovcvYPPM
xHTDFKrkV8dshqbhODIwn3eBEMD2JomO4jeGdtKEDk2etmlIGvjO49ZJ7d1fUiW9Dp+2vD0H0/yt
V/Sfwz6rb6fyYnrPGgoWGlwhLw2R6vy43MR5XzKtiNEZ6yK13kn+oAtZpikOhFm3ygOsgZkD9MmK
zOv/ZmS8wKWf+uuBoQqWOYUQsIP4JqSvGHRUdAXEBmziSJk6vgQhup57g6XvVxQc5FDov+h0KXFj
S1WSkKK0J20Qh4Mn/6QkBhcTfqtTKXeJ3XI0y4trbPI1/vD0t3WmieTNUlxerjYmeKoiKqpAUMBV
yiv60QFSO1/scnjZWGBQf4qLELM1vP04ZLQLK4C16TAZuIhcjn49XKpyNtT0O6yQj1z/WcR8ZEI5
JpH9zeSyHFuofciC9mQ22z1ZVKt+wwqALoj5Gn3oQ5xRPfvqzO6TBi7kjZ+Dm7uo2rkspNpSfENA
eXJ7GwWwVaudDdQK/vuyRyz46LAjh6QoeV8JQJy8d7ehEAxJHR/zFar7R9F65Qk9AJva3O2jTkXM
A+sZfdKwft7qaAJepukg+DMw6J0QNGHQkPFPnAIdH0DSHcrKVRGeB1En9YZ8dJ+D0GBiJz2Sndfo
tRC1TSJM50czDWSlvStBsHEgNUeqZYge68n4FBm84WIR1u1kZhyCs7Wpdm+9dR+bFH+iOmt55/Rv
OcLQBnCFjL2AxaMtgkrPvzSc6lhik8nIQJ+tJwXgeE+il2yw8AMRBifztmdNHgNZUltW3wqqkEhr
TZRSG+Mn1c/yLimisVnwfQ0aVttOB6xtUUu9MLxcmakSPKEF7YHMIc1UpIyBFdD7yBlZ5tjvYRFc
w+VPeeMPQ3SHz2K2LX2qQv8czMMvqeARis2RsdkYS29q8AB5QXMPFN75u4R/cqn9Ur/such3RLc1
Ft5nK/5NZn89sqst1Xqhs6QjG5Cfc4N7Tn1uF0Ji/uywKoIGlHSAN2R9ib6dd1s1Bk7pW5yHTzGO
zh1lOEIIqAvCJ9Ua/7pAPp1oYfN8LNCuxwSew83e9TtwhMTYW16Exc7IpuhxQFMDOVE+E6WvMA2l
bWGMOm8QdtoPIPtdiWoXvwbEulBfpr6meVAbd2Znw8puu/imFMiaEb4dWRaKfTQhnIMIQuWYzbH9
SurMZPrEJBk2JVIfjf+5ZVii1aIubyRqfXyYvXGGmpmCcswNQLM4XerKXmjbQo/hyX/oUyAmMOiS
hiFPbXqxnkmeZiqv2JYJG7nvnLtxcoY89E24svojjx/WM9GgDIMxLEalWYPFOE4RXBvvOIWepB6s
FghSrg91yCgmWfVvR7ZkMsnftGRtYuSSEnkXyc8dC2ffTa8VG5urVsAc8s6YNk4uMi5qz7KFX1AS
DvxOZnmjas0sDeUQPdkVTE0izJKRzxagTEGYIFMHy7SJcvjz6k788yYqOHWW1cbXwtRCBa3u+nKK
gs/vGmwYcIKDBKr78C9U6SO0wmFdwwz2E3SYug58sN7WGI+3zMsKx5arFRYSS5RFD1XvLLrtWVsf
/h/WUTH+2ryY81qt9Jm96/ZgMOoeLCZ8ky5J9ubB5a5d2yANeAZWW9JifkNzLV826Ho3eD6j3NPf
DOlHm42DrDCHHB7H8gMQX6R+KZO2veqWLZZbO3jZBQq1FPJ/49svEFmhJ2egC5jRUMBisuNpBNws
muzp6meX2eHhJdrAV3lzbxHVjKxKnm0YagBkZ7+nJbENVpr8uGIYPlR4GN8vT6h/G0zoOrPMNxjn
tsJfxH+ut5tXU0fZmSy90UCMOuOUcR8hTjQBI/x/Q2CpPvTsJ115IsugigCUia31STOUazsQtAMl
zPr/okqTANLZTdcZfkSXQRsnHT+XmSPTX5ydbSAKF2VECojbQHZ4Sr5hBw6oUaWFabZwYnm9ysup
mS2prjIhW9ha9Lan7IGenrFM1f/tsBmx7yOI7zGd9qB4Fx0Mek3CrTX7+nKU478V33Ca6dgxdCvT
27BJX6LflvLZvzfXiDQwwVtg8iwc0M7hvg1QfSg/Vdv52gUs8SYveMVBatC4I6kB1duAzogeoRKS
G8vf0/Wkx+qw4BGjdN3WrITQREF8n5A58Acs44JFc+Bf974Vp4SFQPnsoYm+OCwZB9WiypgDyAZh
A4OrWgFlLaSSmYSbzYOESL3aeDt8eG/zT8ITl4mM26FnfWYJhh+2x/tUqknoQxqOFMpqDB2o3qUK
50cWzTNOmEOCA+nK0SNukhAm3AqWvRkmwxdYQEd9Vu73Hly2hQV5MkVvnAqa2t2lAptoSMUO32t8
SaSibpt72HsGBNw3WzJOhChpZ8ByzyQrSUNTsQrNgiIaqLSnfi0NCnPhvsN7yCrA9Wl+X9lp1hoT
4BSMhZMxdmjx0MM2vNxZxAg1OvNTklOyrwcJEf10jHWr9gW1XgEMeijAA7sHgArx5rUk7OwmH+35
Me3sLS3TXqqW6LT+rvFLaJD6rerYL1vGY8c2/s/DR/zH7kYxYb6T3RzisxdYLc2l+EkpM5Ynm4yT
SdvY6D/9fJiJKqveAhPKqHSQ+byT28FJV8eP2ucgEkcjy5+jZbze0nRPbiKRQB2ZL/pqfLznOEFI
VxekrWhFYYkD/WW9vNr4KMcTPYsD4c9Wxzk4EjTZxkpsNz2ZdVSTu4NAhq6kXL2HfsBNfdpIdeWr
lLwPBz6tE6qgR5vjBnizXtwrWhtAdGVE2+tBZ4UNNUA5BeC+GXhPx5cJVWxm3kFgw/PIKn0RrrsR
984V85wB/r7fsA64kVEaEKp3owNZYcMRVEPWwuvXQrid+oV9c0DeEcWWDJr6/fwsNHOM/BE8/SQY
iUi9HtGbF0Nrw8TcLnQ16Ih+asong3+dIsq8VsMHK52lneNzvhaa5qgGLm6IFIfPWlHZk6KH8zPC
RJa/A65wZqeoM1F2+C/hPBi6duNMYmNvLUCFMWID3sp4BaAtM/tqduo9H4L/kjpWnrH7+SWiOYC9
h1DLH2cFn5vXj6uvWKsMc03Qvjtqjo1kWH1SoPDltDJUupdWji9o4hokcSStgHFhtM0qfZ0xRNZC
h61AXqhWTB/Q5on6ev1fX6ZvxhsCUoOZHWJnIAzOBAHc4LwKdhtCjqvu5k2/4BkQE68KAjmbIbrV
3T6bgXkDT3UrLBcD8g5SShA22gyTpCrs3XUqqtJga2IG5jIN3tfgAqlISSXvWXzKq3gSV0RrW+rq
iodDkgQJu0v7y9Af7LO7ffs9eCDWITv5KbFaCfydexH8dPYhndHrDTAeZwevfvm0IHDdcOlbCO0e
xq4Wmx/Y2EgsBGpERmbjs/zJwhEiUf4mUOa/8pNrQOqNEIoIgrQVbfDcukH/rp4sXBlAQTlM68RL
EiJY54UH7zdqPtuzWbBp/pqnTTSNIfRxbu3KA3+fJuAhWz5e8RsYTMpZd1tDhPM8rZa9FTiaA7zj
dgH+R/EkS2ubq5xkoJPEY+A7QUnx6K3Vllcfmy6B+pA08l/TwtotiXezUUGG8jHHLjW3r0ELW5Rt
Yr1eTaJJtJiBVhu6AWjsO5/RPEydqk0zWmXvg2ogLTYu5WyKCn5c02sJVnwVc8abaHjxHvmgFPvj
PhDYbSPkalLo0MBplSTqUB9Nk3tDtUZaMK4iZ1eEndtoRr90QJ+Dn05W69CbkLalzX0gZ2lAKl+M
MbHxB/WT4VVAmc2AhL1E6NtpFGbujTgKTzC2R9WQdupknIEx4hxMe2QjLexCDD7rwP1uhwvnZlLz
bCqB/hCtVB3YMnyrjTzHaMHnEBMXUM5Dz62WE7eqFDOG2Ikswzd69YoPQZLFLpMB6UCcmLxuwSZn
TUfxeAJaVlHvEKFIjJ0H25Gbc2tmMw/04vmOYvPxj/+GEE2O2ew4EkrlerWTQkMuABbOyXQAHKhd
XnIF5AbBdJPKp04VOWH+7oDCY198KqUQj/be5fQkxMBeAEJL7acO5wB316NwSL3ZuxR2AhM/Vy8l
Xp4eTs8j46i0gdmVgk/99+huru6T8++t0QEZkSsPaW9JyM9GCvoRZNkiHY9Y8yAhqUucQpO4Y3Zt
jZe5OJybtFxdWb7IKK1kLMo0+lg8blBV7V/bYU/XpA9swtPOKIG8b97v2MK5GMpK0KPqujCUTYiu
NtzMxf4wEIFngJMtOkpxddHVp7kN4Rk3er9X4E2ZcBernZNRXFuEMOURTWn0nnt2TfK/zA7cgQG0
LKeTOAJ4NumfgUHr70CYUvh4vL6h53XiscWAP0JtQqbQfj0QA3TXXKmCx3MJgfWaHFZNCaPY47xb
yqEBSeVsw6Xe0N1gG/5CiUYBnUvG/zGgKTEArQdV0vaONXB4drmbE1qCjzbgdw3uJVL+V390bevu
SjlORlRkggU4IlgL/2whft0LdBQR7DnmmmnNs4LnUZcEUET6o8DwzTyEGX3k31luunUa3leK5IBy
YHCVqWIRlGH79Mgw1gphxLYl1nDR2MtkIuYT16IYGshyUWx7eJdVw6i1mRtScGR72NbNPYDkAGvk
qqvEB9/bz+B6qQe7OKsL4gHeCYZGZsI18m+9JeFgCtdP15D7wwKfjotbr1qePK9heKEf+Tt0kGOP
YvxE2nLGoeESEp5QbPxTq67dLja0UunLB/pDbTwRDMMStaG7f861a1v0uscUuNpsbiktqRRjirY/
ROS8yMy/5jWj7oRZtplQcGIrG+pB5q++0sNlpIB+ykYBRX7u5ztXaI0OWzzGjj2PRGPzuIPPhJWS
9liKGFJGiX4o9LjzLZwtqdzwQUQFKxhV4xh8WOH2wrnVpL2uRG3Am7wxnOxgQoROSM0CL0MxgUV7
BUeRPf5gGqKFPkAKQI/xh6jdsexofckQtQhkwTPS5THQaMgpfJlaEHRTQCUoXhWyjshtUQZbN0Rr
2sa7jnMJD87xzZQFiBbpSb6zRHzGSTqv1bzTx9lwu48JVyEke95DfJCojGwmnKzc54AzGhCSXBa1
MSKsf6B5wuPVN2XM5BaSOu5WbIoJ6gjfDct6/6gtQKaXd/HdOTURyKcZ6OsZtoQ5tTywfsTXuIkW
lckmWKN0XAgWII8OwXko1L02QNXxp7Z+mk4Ttb+tyMlUKOgvgEAYN3tXbrmIUGNJEArPwoAlAv12
Uz7X6KMLuurjUhGFqCHqd2K30hX4fn6PMx4Y4UnXG2eNTTLFGAa0tjmimC/QbqvC1yURxLTrn4k0
pECki8fqaW9WwE+iMKcCpkyjXeWfmQt/k8bj66piiF0pZsDqqwNcHoTDbON0ijPxLrIPughWbM9p
1SOpULUW8pnq+cPeSghowFxCX1HyD6BHnB9f9l0bCL259JEBRU8aUsv0C0jG+fJ8xI1TarsHIFNZ
VHyVe85d2jPpOyvPXCT7d6Ix2MXuWl2Xdx8fP6nQx96sbnmFXenShL/gSgBdAPnZ63FvHFalz3Rv
fd0/UPpK/cY02zrfQlo0/XPVIY+3Bv0/Q+7pMzlF9zW12q5MEJuM6iZ61+htM+MfN02Y60ngc+Qg
9vsPErIO8xkfIezdIo0kKG7PZm4OwNkp9bSfYyE4jiE7JsX5ahx3pEcDITTmj7bxvHSiA6Bs2Ri6
4Win0/3ReiaG2lVFNHi0azhd/+E6fJNlaazlhzITAVzj1WVAsJzCBtdhI9zmSxzy4w3X1BKA8uLc
zlHMjp6P5zO3Rz2QLa1MLARqnoja90iew/KpazVdOTsV+5yUWZDe9IIRga1rWqJQCH05MevSGiNM
sM8X+GX9ASJK7/QyH/9URBWRZotN8uep375ezl7anekjTHgQXyHWGtct8ISBNPZ5Z25JtetbXBOe
Ga5ucw2xSAErjqGQAS6xadw+/ZgHHOHz1sNP9jNEku2AGNDaFBs+Zn6yVCXH3c0GSgrlnb5Spf7Y
stMLRhWWpSRCTR2oTmbChDI3KMOfDaQCsWKcPML4Fmho0q0ilTEwuNJdAp7BNEGM5y1ktir4ezF7
h5mnWbpYmcSao0XQK6iLybf3nhr2DHMKLz8PFBU7GEzW7zsEcpr1YylvM1U5KZBJrWFG2mXUHEWc
H3F5n/koj2jQtIVLBeu9ddbcLq3w3+LrekKEU4vl7CHGWnaCKKrmX39Ozx4shEfTRWa3w8w/RSFy
7a1c1jX90QOjQ0P0GnsXj2PttSdE3hw0BkLBhT6sRSE2TxCYbt4+CRPT52lYWwP2/iGurut6K1wL
8Ds4IHxPz8PtaPd26LiT3AoaUBnmXyAM3gRIwnFiZfEzZseVGVba6cspZ8QSqOCdgWoPm2L0XY/G
+aq5h1159H6D8I6CYUzZtFmgZqnkpNCS3dgotZ4pUgdSEFgx1a0JrdaKEbIfREGnHGCtWweBMbXy
/xO6nz0Fqcchc8KK+Fi5621hLP8OLYGDsCLMq4h/XGcJu2iUeJTbUa82O7MjlvneTow6giGqMKU8
OgIxaccQ4STdDuo6u0g3DIIrIuvrpssAKNLFqqMphKl0EdyI3wCelGqMShwYo1XHHK9C8QhL97rC
fjS6m1OUhDKyDYcgg7bmphAmt0WbtLTdLRFoDT8sFhrHW7SIkJPyPYo/3utBkYzV7rdLyBc8uKdx
3ptic9Kce9a1QuIYwjQ4q03hr258my2kdsd76jKNcpFglFC11LjitKNabu1mpG6K/9lgW/ovchnm
Ytiuo7aZryAmYFd5arpiW1MpYZf/g3K/d9nOyGZbg6355fwV3Bg2SmoXxSt6ZwEPlc9DVyIo1/SA
8EYsyCLmbbeDeEG1vdu4R/x6gGj2Z2mjsP/STQqyu12fVYtJAKaCCRQGoAeb3PyloYwZfNyzU5uT
vFLo/piQLJdGJPCsfgvwrKH58m5A8xIWi/0lbGrX3q/OVS1W4tZjuCR7JJYe2Yl6uEI2tnbTyO3A
Mh+bk5xAN+BE5t8voTzDpzSxqCVISIJL3mwpuMmT1ZAprHJ2wAHPuE+CqhHjSNU+VMX0KUVKwPAU
6zrK9HXzBzbU2S7VKpX2msvnEvr0tEwbLu8wIAojbDcbCcTV55vbzZETffV692JiSErk1n9ME3Pm
m1pyK1H2yIHqNetsQXEY9heGSeuEY6jq8xWVdt8+DSsfeGN67gCQKw0IodZy2uwJEcE2Fc/0mNsI
dI3GbRNmOjMLdMxEbVoeDxj6TQ8JwUdIfew7sW/IX5CKrAfmkTnB42oQ+LdcYmmkAYzHNWuioSGM
xdBjyXicwRmVfHgu3C8B8eihomxqaMxk2QL9iZfHoJgo9+LlQj4Pn0l5dXu21B7KgOvBPFuIR1Fd
Gv5vFrRrpFy0B0mqkyEgIZ1LnjJ9+k9wMh909mP87Cie7JFGPBss8K8438xTezZb+lf6VH9Bn41M
YXApN7+em6cZvwBQ7cv2+ABr52/9bzfyQie4B+5eYFcwAuFF0TDshrWRYO26q64sqyD/MRx7AoDw
6aa3UpssZ0hI8IyqQxTn9X8IF7smIfEJWZ8hGjQueVpAx6RdjztxusyK2wyIhVcdoDKwxWrFpsev
FZoj44G7rQrDvlQeXc71b5mCq7sLMVNPuolpTWkHxwYnkvS/M0Ky/8oRZV/OBZAu0zylwxIMokhV
ZYDMhHMwzz29zuQ6LyKijqQkCVC2ykC/md2eHYtGLOtQOCt4WceExA1CnpqRzchtDqpNo0vd8NWy
x6+4wE1qFTLRfSYDfUOYC/RLcMlTk1KnE/FnJq6Ez12fneC9BTsQQxFoB6OK79q/DQj/GuQhNbAM
ofhExjx0jnNloAcwBD4AnjqbGR1nQytBv/IBFXxWZvzaQvTRZpsR0t9Dc6EylVA+Q31IlbDx3qJd
3u+GdBwczV7QH2jDZHHzQUN5iCiBYvyCdLrJpEWUKBlWuH9ccP+JIsjC6AkUF81c4hKF/mwCTtq7
7orp3dhV8YlrwvIoztJA94SPs1AASHMPwtdPyNppyFf+PW0w4GSD37ELNc1lZhEZvjxl1mD0JqbU
zA+bcAjCK5Ld6xg+FQ2QbEjmidw9ODSP9ItkBlN+WJQFJFqhkwIwUthpdFJugY028nxlYXZqggXx
w0676T2rMX9Ve7XBytZn4PLFHCK/I9ki71NXTkKIm3Y+vf/eNiUY3hRT5s3XucxBM0z59US8FY4l
/w74tDiZfs85fyu05Cua6TagdCDg+pmq/x9KdEOhbHpAgklQNr0HN7bhHN2uAlwErHQanP/Wz7H1
8xJYGOLhOoeXdYNk0LjW6kC2p26svJ9lq9vXt2JcK3t1rxnEVGDRbj8ZtJ+B1NyWo8qADy+I0Qq9
nQs/yh900ZrZrV0vtQ+3NohdCZW/gwb0xA8Wx41QmNaF9eLxBtJ3wtWRSRXcRVuHhDG7vL7JyWPa
X3TeLbmyDQgI8pCBU/YzT5xZvdhObvXTNRxIM57aHDduToXMAHCg5ULL3YljCoSHgOmrBoTU+jHq
qFfP4IovtKqQ7OOyMZwWi1muPO4WpgzKyrl8NtLfymfC3IKuG5jnk+Pmbin72g1+idfV88KVRVEa
FAsfBnr1prS/HybKYXytGxOs9zx2BLnIvC3LCDEO6p9MkrPeUf5mGF8Ogy1joY0w80+WtA08IlKM
wsG3rH7ylc61NsV/gEhTYL0XxJUublNXR0sopMYit/v48Ox5phvp7V5Sda93ezBxlyLGiEczaaxL
5dOgVsDekYg3UNhqQY+tIxsM2Lfqhs8aJ135A9RXBicv1UuitfZeEyEvCJu9DgsKYKvi5iQcQmnW
dQqOVyrET3fh2gAL7VHCpGosYNl4PTUtC8X/gWdBXhx+I7e347xeNluGYTwiQSpkiUo8Pg1u47zV
SUV3p4jOVW4sKQzqiX7dYvA+sNgXTVMMJXd8DI8Fgo6czvm3sBAoyUOqvzMZhjMKzArZIVnlWW/e
4DLjY0fUL8v/gNIlCLmN3BMzsn2bUQsQxR3a3/h0AumTqxrlxppR6R82O9ozHvijc5I0rogumSPs
4TaY7cofRc5HueSn/JcyPPRuLaiL7Pf+EyPNuYqIGHca+JgaC38vMatR+u173g304XfHLgMOeylg
LSV0pFGTRZkRSG3HGunK0soDRmaFoId/DzsHPnXzPeWHycI3JgEp1Uy8BHwv+es9/KKH/98is8hK
RPPO+XVepdZGJyBD8UU/bxrHEInxtyV+D9YtMuq2hMilhkCZsjVIrR5yzrlnZqOXDPySkQXFLxas
pzPlp23j2SGlDoV1VtPpNjVSxOy6N5mDlcK+lB0PZiFWWtSktG/xFXHImXdEMCIt116MQsKELBqM
G09y9fUgRojNpkdr1lasmquEaRq0nrPa+/4e1MGWv7uageA6ssxd8EzHRetT65mvBL9N1efwcRXA
upQUglNd+J0DiJYAaaUmyAmqxGAue3BUUZ756uOI9kTb7huEaOkDwKzoItNR6yW7nIwVkvOlCJX4
8YQb0dJlXquvnCZxtHwKtLtymrN2oLqTIyo4oHsGulrhYupSN5I4lupivfBLmG5OFeYQvXsKVIMT
yINy/bAtdcrs/2qo7d96zPsoX8zfIrbceADVFahK/cEFzxvnmeMbizlxa6p0i3PMqpn+XIcBiNc+
ictPLKpdPTEf5cmpd+1wFJA7umqw+Z4eI+lZ1F3EwlcWOo9Sb353K/XQvpV3GlKgbrh+yMIbjcCY
dAFjLzxwGu+mH61gXx6O0vqb1Bto016DszwWS7TUQjSB2aU8ZvWkNgvf3VO6OiR5hdrRCKEPLFcL
+mGUkJ5n2c3Y6TccXPzblbHYNn/gzxBvRoTIvF1AV1Wghwe0VgzYiQOc65/U3LsX6mrjR+pRD128
E6zIc0zv2gw16gkNsTUnZOuYUCraa5vGuO29V37InvGTjx20iu+8lxP/snYr58DBkjGYycPBWrGE
swzOAi58uqKTnHDZ8pETc7NM1mL+tWYdu4TULk5vv/s0KIugD4xowRkIWI9ZIEMlEXeMZBUEhqpF
XHDhNJNNBnTdOXgG+ti0oFOklmsjLESUx91o/3an7AqTqhPxctPUv6ql788n2G1ZbLruexQI28Fh
RP4BlUbypsf3z886NAttO/CuonsqCQCNF3kGwJZDKC7RZlTedE1eCsohiXdBAYXAC4o50dxh0STt
SIydvppWG0aySTxKo4fDgAR6Tojf9umKzSAxvo4B7Kd1eEIdPQV/3xjav/IEl7gxLYI3T6brLSfj
mfya0r4+Z6LvKCPBCszfLoS86rlpWfbiIFXFPcKy/uMUmRtt9vSMkAhgitzkSkjGUpjRWNJeYAt+
G9tNgURKKrMWsSYSvAr1BgqKCQQyT1zJPdM4nCmofmoFTrYHADmlExjmN/6YQRP0XA0HV0o6js9Q
/vTxCoUJgtppITacDT6QjvI1nXzmEn33Td0vaBg1VICQQ3FMO6s3jfnrxx07wnKM7AXATB3izMb7
X8XnE2b/kjXby9XgBvbd/Ge1eCgkd2iih+m+pcZHRtzjSI0Ys8CozESmG6Ok6j7X43CzFP3A8yZx
BMqmj2pxVWmCZgnqcjUrIOZ09NdRYmc+pwWkAyVOo4JQaWUCX6Wox1i2JNFN7Qm0Rf+XApoE+A8M
IxHGKbzYkcMgXQLvxV14wVD3R9ipwks6vZrKdU2Z9Vx0z7wznIbnMQbWza9Tv0F2ajned5ZPh3xm
EcQk2HyMmlZL0TVthkkH4/v8aoNlwz8HMAM+L4dDlRx27ygmpNqoSEvT2R9xXkT/P7AdBfUKYVDi
x2vdw/U4tiOtLCoRg+ZJXFt33lbOENO/To1inF6C9F1GqktjsvErFq0TDH7k9wmMIS9xlhOaYB35
jVNHRXgdy4bO1KhwkNKwEcm4CtF+jPSWUN8onbn5nSNDbYLVWRFtjyPTln0fn8M/F5O4djx9lEG9
VVwdUdGkQmePLtDq7lKptl75OxBYgCEGPphLHjNFpNkfnFZ7ZtuUYJtgqbbdhrbEO/B8BVzFC8Qy
p/rINmu6y6WNtir2aZ/2vN6KmtYEasZmLL1S5PU6o6ndKLpSaswLytPCJrQTs3oxQI7vs7Z2WEeQ
WkqoSfqaPOduWqyiIP6fVN0xK0++qhxtO+lqeu0pcysvHvx7S+NgLo5ZHV2z2xiNFeeVkg2l2/md
R/mRqQJYE/+mciUURhpUHZxjSWms9pcH8o5Z1PTki8qjEJMdyTUHHt5H0J8uwdFWkdWG7uUwiemi
gpP5v6+gDkZL72cSON8uuWJyOntdTIkd5BxrXlp7vjJOJ+Ug9jguQsBxxdDx97F9PfoRSJT5bjue
X4VQNFCtbqWvSdgcPv+HT1lOI5zxzHw1w6dEA+qiNVGohgLjf/LGD+ldLzqdDX9PiGDgNguIcFb7
L9/7STqU3M025nELcKnv9AitR8GAyXQavZyv4Jvfn8PvKukvuZPrEIWhTQL5lEMwPIOIA5W4WzY4
TzYZfcOyiOYauu6cvYDrHuGMTJbGH+8unxtH5GAa6WMNUHx2f6luO1NZk5YHXHpP7CVpLsNvUcfg
BG9xKSM/9+pMWFI+0uqEsi/57+A2ZZqfNUxEnaFX6GhXTQ/cjnPRL0XCUwbbCDAYRpmtKX2A/Yqr
9OOfUM+Bm+ZaLOFXeqto9Lqe7LUoEmcT24IZe2fQ/HAxZ3SnzgFjQMvqVdOMSmnFtmVOou/e0ZEd
0spv6rN/H/vf1j+rGtuGx6ZXEoQ+/aGyIdqpcDuEBxphE6IWy+0j6czaDttBwgaLfGt6AB2T7WTu
lN9X7yGmRVLFBHqicjX2mG/KKqKV2G4+1mL1GVxdQawTN6xdCM62x+jwzxQUBouHS0F80UuVPRFH
Vw8xHiS52DyQxFWK5ZX0x0oMnYE9grhlsSD/qEiTeQ0FvtLUQPUYiCV42Lntvasypm2J0TQBw4lS
gdUWcW3+8q+SCcvf3rQW2LinTaQA2yPZTk3sOICiPF1W5y9hYgl2xkOPbN2M15D3DRQ2OoovUl5S
EAVYwAF3MjTnTL2YKbvHvzOksoYENtEWXzBDWYYgK5AllsZgWH5JoaTfHRBcE1sXkEeqthGLfCQW
51agrOk0IhhCbFcTdx+aRO1pduFK/6W0aT+UjhaZTP/6LbqWmG2stXcO1Yylovv349ctCcvMS1nA
yMKlHnnVBwhTnakhxsZEag7Ur2HDNYaIM+qFA9AQAAob7JaiRaMUisNV/04E39kG4/WUp/VRDXYq
vxEJu4s+qm3jicmsbz4ip5pm5m3fSBwxTffvcPwx1lMcxtAqde4v8NY/oJxJqB3HFqX7nt/DWdf3
aolISZO5IbqQC94azTpkxqqNuSOHFE6zVaFSCEDhivSAYdJLtEizFJMyPr8HUReACGBCxx9RJA4t
5m11bnDBxxUuZqZ98l67NV/nndGayUN861QA1xjg0wvhOOSqRgn61td3OGXTUzJcHrjOrHHCJgGp
CtUcR5T7c2e2oj+igc6tXS87KUucKxEWtwioy1/1iGP0SSztScO5D2LY2GuX42k97WJIMXGMcrTy
UFPqhwb8rqiSL66zJNTzf4HlrL6nYwygy6hyFzgvEM9JvAQqfTAYOHj8e1Exu9yLNqaR/ZzAA3PR
tr84jrHM7WRvWLVbLHmOSkn2V72tGz9Aja4o3MDuwmJf8LdQ3uhcF0tusQAdnNMr56Mpz0CM5bLj
9mXn5GD6it+S/d8GivQpMAniSisR83ntYGAXolZxdv+E/XVFDJDs3zi9NgoshXquuMqk9HPE8Dw7
bJmV2CFAo35toiJ1ULid4bRESeUN12HqAOKCsZGUvTfsz8KWCu1uHwJ52DrC5QvIEnYl21y+ZZ2S
5kxjRVoeYWdJs25GFopvGheSA/7K5P1AYCO0NIYX4i+hfbNEzskDEOrX5+kOFAiVItkY8uvu6rWk
gG51EyPgBq2tfQ30zhPZt+gFDuwo/bnQ81z36J/KNN+8lXRo0nOZtodKuxkE9ZWBIfeKr+Smm2hL
hzYIHf0heHz+BpXvUWzEHV+GTfstTJIzcuPFUQpiwmrlh334zN+LHyUupOdoRiJjuAGwmLAfSKCT
9eref3DA3f+pRzQeseR3K99kbs+I82DUvZ0WIGjED4GaTP0iS6SraSUH6f9h7kRVjmZF/FvccbT5
ueqwzbh9SUrWPGgQ8aHN/8Q5oOWw2wY8Q39AYOoo++xhUP0dD97GFiHIF6oBtm/KJtLaN0+JGC0Z
zsD0DZtneq1QJqryAJNRlhTAu+V4d2Zv69v3PKalsMt4BriQTS+bCLI812XKsVK0zsWIUoUoCI2H
g/iA76TUIQnkSUpC25FJyo5oRhsy/vDz1iijtcNBT0JDg5SfV2PP2TuIYfBOXuS/8P0vOsQ9sTaI
RsZ5c01SOk5pT/hnXNgOUhe8lrPh8hYj5lxgUdy0il9u/SamZU/yojQ1gmp3JqAUa6gSASk0OGzl
+rHJKVeSTH+kfDB3l9xWairw6uyzrU2nQV2Eq6Mrj/CBK4B/7VFjarEUHuAmgiunWxDlKzrhxsQN
lMUqKGG7HSixU5CcRs8fi+mXfucC9Zb0KvHbWhZp5SrjLa73pF7Z/SAp3ehkl6JEBxPzw8VHXNdx
l+HS/jwXL0ZOTAflTEQ8zRcV9GjHXfHuk2vHgnDs+tYSwhiU+X2/4XTSDjHqkzoI/E8IGiABKhrD
GB5H6BCZ915Nwz5baqhrhRcMRbrExzd+rJLMUSmducdioUrzBahcI6VTV7rQ6mXncxwf2uOY8fhe
2xhzEAGWdOYQvAePaEyrMyAOmtZ9GJPb1xk/HW3U60F0sEAMEWEaKgwKkDDYah4olJ8H1XHZQdWf
cvn+gPtk8MvUJKUn842HE44m2kuEJvqqxbIBO4x4ZQ+kDIEOtY9bsiTCOBIJx8Kjn6n4/ktieQ1I
sYDpgn0kfkTZN/jFgijbHIEzrQoX3IkQbz6YNAn32yldIdOuQOJeuRfkswAMJ2YtcIye1Fv/NXUB
u+69ninYLSSNsy45xd4uYyQQbn9esaoi0WzJPlB8vp+EaH3uExcEzhhziQqScbDzcuVxgIhonbyY
e6FOKwGd9GrkjggsEx1gzndpv6+FVaRLBP4GSUOnIMHkC4o3G2G5AjQRqlNZ7pdD6tx7Am161W0z
yEIr0vtYq23ORizyiILFH5ArgCYk9XakgdRQz1XUFiwqzbeie8KO+nIM3BjI354/IUjk579uRCk8
gHgNvJyGlgTdQkqHca3pFuajexOYesvzOf/+Jgidf6WfzbVpySoqj6v2El8kpqE9WNf5X590dCEJ
wnz03idb/SxPSDl4xp85Kh9+FTPWU3EjrooiP24yUO18+ZAq5dI1SWxSMxlIiSmFE5LOWwDM5Vqf
4J6YnX+iGRufKVlOFUqI3touHZ6JQ/g+3UvvBxqRNS0xlfphv+G/TFXlW0RWsT+1xgoQrGKkX63/
95DbSRNIWwIJAjJ7tVNyA9ZKkUVplLsJm0ZmW72IAu0ml3DqOFWBJL9brmPj4wFOD8HMeIlfUWqG
Xs29aQZcSlG50jnolsBV6AJUIGlgCnYy/btyBrTRLtHYDlDY9OSDzcuky0kGFiwR2Dv1/qj5ZqOs
QDik9RiCvXUryZQQU09qp6MR9p3brzhBkzzXI7Wfhkusro0DuM0G/uhvg476lf+WRu5hf9J6JVuJ
OQ9t9/PibN1rrAgJJgV5nAWcLSFX19iImUt/EgcC7TFCdoNCeoJo+Aq1Y5jVmUeF7dzuuszAon+B
4AmnIZoIxNvGfRPHMb/zj9PuJdRExpmShh1BF83678h0h6o3AXFOZv7oxdpDYVQ2y5K0HpkIRt9K
jA9nDDI42460UaI+WzFctH64xQxp0WWkVdRZmedqePxZYON6qYDEr/FOmD7Yu1Q2Zxf2+BmZt2Si
nE4loUbRJpjQBSfgzc1p2eKI7e4L0F5seW3iAhELur8gazaaPxkGqvW82J1i9FNG37ZGOUxemyHO
UqOZbWwvP0C6J+qSC6gl+brJ1fud5kbqW1VR1Uhn1B4SYAHuWNkd8h5t3kdIOITVetYSV5UXXmlN
VhKN3qgONMDEpgGP69jQjuWMW6f4XUQt7r81gEpstOHgoXAg9PUUJYvaMCKAwFeGT/IWgoDebU/I
EQRY8gpO/WIY5SnRG1/y9Q9EeAv4RAyzM7CtMP6jM1QtnYErPbI1MmY9g+p6hbwCDI+NJ/X6xt0c
0r3Xsdt+m2hCeq5lEQVdc+txorR8MnJ7NJ0TqEyyX5rXp0keKgwWmNl38tiXlD/OBOrFlJI48ZcU
w8GMj8vkoNoPDDl4wpBB+7MqdbAn9gz5IIejfZXhrVVu3ar8Tbu7ekHcD/jKcZgeGg7546b359OG
mfwng+rvMLpv5aDSkohckdBFhwOmTwjQaSa/xhMEvpMLHigVTKPafprHG9Cv18z07qW0vxM97hoo
ZWYZVB+5p6BHnHeh95v7zTTTyi1zBQQsurk8j8M7MqDC4SdD4vs20SNti91i7M9VwsvgSCM24/N3
NWmOnOWArD48n44DEMKgBLB0TyxLY05GqhcmpwkJB5HwBcXGn00slJnflhItl/ZkjckOt/KPFoUI
4kzi6HS4oLIynzdF9Y/af0JbkwaXMRxvt/gxdEwiOJS39oLxBZlsu0zLG3IfRqu7ftmjsxyGRrtC
zJ6qXDgbrusIzVAFofgFK9XGzI6Iz2xKyqbKygjmjlz9Nv8tgmRmV5q2jgD0HvPYN3CgBTFt5fAJ
jawqzOWRBa+yAVNYai6/KdPscYT1KhZFwrrMoLF8ewI51ZD5FO6hjcYzyWvRSIPkTZ+A/mWnmHGi
V8TnhMDOK0skrsTBmYEzxfdqHLlTNk+DbA17QQmlxUr6UuauvwnQCXtqiIOTtPYyYc2fYpQOXd5o
OcUGpHZqT7PFr9VOU5jk/NfrHxpuhN8lxio89Io3ib1zjilr9YeAZyscWdIC4Luggf14gd6jPwyI
+U7n9Y3cxF/OViyTjFQiPGSmSjr8+Wl7nbepnIEqbiL66LZfk10nGbyvbfMxgAN62tAaIAngGgdv
ownDvl/olP+50BqaM6NA3OH1g8rUcOo+C/x7h5Of9r0f80sLMKv7SBoBVlTDFE5+a/WtmVAgouNe
JgmPpgqchyf2xixSjwxj6OE/a+/AGeEZ+qsGPYebJHgMB7l8TRTtinTab/0ZT7U02C6GtDTmk3Bj
sbclgoUTw3m7egCHvt+dfkVFg2EOEI4a0n2+bZMYnVkUwfVdRGB367T0S+QqlMzixgEji8wxB+sd
DflYBDk2Zv5QB4vUZ29BhvOlPoEVk8Li8eYIrW/cCLsH5oKEX3RmuZcRgKPSA95AdGcGQRsEk5tD
Q8CNllw2v+Z4aDz4gSGBkrcxDuLXRIju1abAgy55LFbH15nv1kKOKav7lKvEU+W78bkIyoVE26J0
Gb//y2SJgSO1tZLWcxKORTH4a57v+DkOSk0PDt05LGCd8t5cnAFD13xr5xEtYlpkOkoOj7XmbIuk
p7qYmmEl9pgRwEFwuFhlDW/3GW/f5tMw2NfOPa9PKGl9nt8IzYTutH2V+vIhvSc/zzMVyB8Z3p1G
60LQY2tn6jJ4V7sKtaRMJgTj+K8YAux+H09auES0wNOkagErakL8FxHnRqJi4dhOmLtocWQOO4+b
ISH+xzAISYCuXmrkCe7gelVjiYsASZS+wqraPc4oDFkIjVqJ530zLJGQ2pjWIkj/6TgCg3BDi6NU
OgFJsL+h+o/ehSSKeBNMrUpWw3cOq4mlGn4DltJCQoGoI9j5Fl3mzkLQ+ogMxVNrOD7eBmci51cS
5GazDKcLvlvF0Rfs04zDOA6/8RssbMNugSkXQg7TaoQ6IgMFi3Xv5h/AnLurlaTjtqA4zjSiO22C
GOfvMhBYa+4Kl1WJUZfQTR8BlI/pIHtPzsLVDjEKbLH4KkjzreBwtQqie0umMQ6yb/lG698GiIJr
WSFGgfyKBCwpsxgO0RrJYRYNIig9t+unBtLcXW5X8zCE5G2dXNoyWA4SdEi/tD4R6jPD9/JdYhjO
t2w2VhDx07tuw6DTM+TfYWRPxmwJpdARS8wQio3rk+5cTK7Sd6n64kDFLrl2ANF5DBhDC3RzKhzL
II1wFjIYHaOIQhyqJrPKut1c+SCfCHXANFbRvxpgjLfFD9t3UtM3mrYg5zB+YUfu2FEju6L60/zD
urY3rx4BozVibMvVyQ6GRznDfEpZPfVN9xWbkNu+Uzv5ckPsKttXVsTaZ/BT11hgco+v9c9LHqq3
2Ek5h69642VavZQFa+T2rYVU4hSQ25wpkdeXCBkrdQghu+MsmlUo/pguB6H9oUeYxYJH/U1cdHIK
0xiflC5v9Rfb2kmkLmN2Vg+TkiSYEIJK3t5f1VWcI3a3TJPJIkeBYfj1KjjeFqmdRl0qElFVvdVY
tsq65ElvqeDpwL9h9PUPmYUcikPK3HCCe9fmd0UWMzE5Nw/Owrql/sqmNv4ypDDuV9A407kP37Qo
btS/uBFKPn4iHN5HdjwRXcW1OD/elnKxcYND9NoY7wDVkDdAZ+IAeiNSJGGfjoUirVF+UvbgjDKG
Wu6bQNAK6GhR59tg1Bs+spzbAxsmqRUTxzURVa2QJocDJTfgNIud4gxSJYraPRfuiblqVhZBxXhN
dotMyWzv7wALGPlkdV24Smvc8cXnDcCvumP7u8MCHrdct9np+9kRP5bmxZKN56RqGa/AlfJzjtw/
tGsm1MlfxwxSEqj9JXHJpdJK4yLAcoKmaW4QYGbu3wvdlLLZrgWQhZQDv10N9tlotgmsSq4GFhi+
6EzcQzoSDCMCiuYOyFIPooMmfL/AiArmistTNzMDFlv1Y1zf0DnCuUgXmzpNxhYdvcNh8Lx/A4No
iBsXVKelmEMuxnYc1zv0xEumDNyDc7IggymOGqB0vLailQLPYcyMEkynml0zTpcAAsqNQ0tLqmzA
OB2TSt/lM7dZ7Zc7PmrPVIqxFtKykFzeszkq94p/sqVyHy8ngWRQeJf4OLMfIdtPTHdWdPq8pFpW
6pZcixkpQjIuecGm8IXqqYs9x98CBObEREh/xODxZbX93vDu8QjIwku8cfIXvWYITI1vk4RQ5OEM
9LmYp8YnOCj4m0MVeaf/DsmhghidkxluiWCaf2CH3v6HnYpDleXg4pdFbto1QKMnICDmYMHi+yTY
sdPBN+iLXKAV4R631MMU+WeIVauGAl7QpN2f8fUIkr9ntsjMDdS99mx8vAS37/K+/QVht0SG+WRT
e01BSzuyfiJvhQ8xQrfsP737Znm3sqRwfc6puKa8VM4fYrfEFwB3uga81HKzq81pFVwWc0bysyrZ
TaiVbQiAaW48M0lH7Xw+9eYYSN65jhe0ZYHL0PHHopx38NtJB+TPfwit8DC0PQY79UYEb1ZoNMpj
AQHOy8uMrzBZVqraP+8DNd9Jdwik8b+IdEWxT7MIIhz+Ptvyrlsd1k0qLvUKaVfmojavMBXkLgdB
nmtBI5z6lvRWCHpGLHTDxAR3TtU/9yPcahYNGFRdnCdOakoiPttYVnvROI7rQsXm4knlpmqSoFDd
m+YUjHc745ucN4rMCOo300vkoV0BBUE1NJe20Bp2b+gWTswdwXgGSxJodLBW23mfL6cJ13hHrMTL
/e/7r7G8NRGAQFJ0NnqlLlzxcZJdNscBrwwJIsnxYmbj3Fiy9UWQQew41sMSCV9cmmRWpr/H7Ngo
RGm5if+R2gnhnR+NC2SQBycFdc9H7fHJZcR385TOcXMdz2I6DQhJx7ptF+QW56oFXCNi/gpomkpk
C7O8CxFGLh+K/PNYyEgAZk2bQwFfuacnbDDTNH63zMd/ah/tsZw0vzv3Ne6nhhcNLG77OYcrUCym
RVRR78yg61arPml3L9wfFo5GS14kngCSEkUaC79epiRMKDYHBzQzCssublStZJl5RGG+2YzzXds+
mRt15wO8ij4qv8wv5l9Ffz299VB26X2QrVMFna/kAS2wT1O4h1rycwcZWihEHtu0lZBsyYc3dTBX
aBAJcDlv1yCxRlONUtG0PatEmc+bciHgFLLAIrJEcRUh1CUdiNtmxNBEeVgoIpJ2k7TP/1w6g6qg
j9wVzRs4llmHaYRJuLQCEOeE5q1pnYvsRZjCYuhmP79xiED2PRnFCQyW+S0witcCZ8WCWRLeyRI5
+r19O0KXvms9ac9Is6E8uWsyyu3SWpPK0Z9UUDPSRuOAgHN6Kllq1urYrv/UaYsG8Q064VfyLz4r
YnZ/zC9z98NXqHBvcL0JCPFP5vZsD/fNARsC5FwCVWUw3L7pvQvAdtL793buYLVoVNKbBjNt+pV7
m6yF0Glo7zRckS+bxker0v85qpZYeCkwNQ6Gax0dbATJQTvuSt/jqPTfkBhyawjhoLb5LgcXCIOW
IUKFw5HMWhxSF0iWuneJxMOmZdvTEmhbkIsXQX25a/+2yZVRiaQetu0m3a7RfRHWbpm/JGYqq2Ob
i0Y8wHbLsk79/xtZ75U+z+F+gCwKcIJce3+dvnm1CZc3RYhOpYe81kpaKEEwvksCzat2B7OjnL/i
wQ6J+AhFhCOyxvFTQRQSHHPKqe/6sHfWcWoeKtxh/msZnJELpz87/GQyyzOwz5sIRC/RZUyc6qbN
sZ+PTmyzrvrCPqmvbThEhxmZNqjAPOJmsoxnDaaIOiXhRF03aHW411v0AB2UyG1gR9izGgULO21V
e+52AcW+zaqTOS8rtACjOsjSlGNo8qWMWqIey4WakRukYp7+D6mP7CyOXCHCeUYx819C7wWTo7pv
hiGSUEfrD0CBiGJDfAuuaHmaOhl0bEUX83IigF+mhAAvdQPN4qawqIq2TejH5b7FyJjjAMtadQHz
2o7oJeDj0/izdiYVyOdDRLXzB4Ca71y56/GGAdgJFhWM3VZgxMRzGBZP1TBYlfK8yfH+MYH5ztEy
a8/nPnDYMVWFZH1Y0Y5NEhujCLWA66bn2woJowmMkZG2rgRu5XDixaozuBeoi5ohHE+Lyb4I4d2b
QPlk6Y4zkdJmbAwb2HSeEkB4o1OAhM3oDTe0Te8D5kATRCncnuJaD8WPZdQYJrhBuyPvkQAAAv6n
7EGxnEOMNLkYmHhVOg8DEEiS0jZWmWhmEz9MNYinbt4+g7Wypq1Wecquu3bacChhEzb4uB9bUQP7
VIoNVOPTAY8cg17WcfPx68Im0M0LCDPhInNQh/7frS+4m4/KOiGp/4cxTbJ7V+wJu1pOYyHgenBQ
bYfPIlwa6GFN2Gnw+2U7dF5WqBJuYYBcLOyhPA05HZzaLP0SX+9vtKII0JedA0uwwWkkhKTwSLxV
fWsGxefUhvVsMsrACSGszUny79fW5Hy8ND/OUEFRuoPdQkiftTWxPyxa1p83sxXNX91Ut4GWqy/x
ovZsZn0gYGnh2yG6NEnDHvGRDWLnr4LBk+41Z6kgzwaVEFP3J0eZE1FIYWy9LblYbwXLHanhDk9s
dCEIe8A5d8ukLSVOIyxaTaJnSMwOmjRFeEjzdVqHHnWeG26zCC6B2KFhdGgoDTM5AYS0Y0jsM0VD
xMlNhD4zFjCdedRP3e4sy3VeuaQmFFE8pZ/aYz7VsllPK1RfT2x/sceR/NTpf+FH0VedIaYkT1PJ
oitMb/nUXSfZDyckq/Je7bNymOsof6R39ru92+NixJCPJflcHiPHoXPokJNM0wp3WN7e/8OmiBL7
gHPG4944Dk3ttNDtTVTajqNcfdyRNjWrEbdS/MQoOPbBcMY7DSIKMk9YBU94viE9jbxM62lLGAcq
P5p64+gsasS4aeN01fDvJ4Ee8mh9mBVafswtD7+f8Y6uqZdM52nwBts6PIHWbObBRI8FlrEBOjf6
4uEk51L/Z9JRSVhsrF7VEJf3X6bpidOJWhlcfsWDMlY21rLlKPdM85a/g7rNII6aWaWW6n62z0ol
ZMI9OzeuhFdEdYzvbdqjEIgYuggw6mjlwhXFWhOgF2ojRf1/QJhnTxoz35kNt7+rfWXOaKyQmud0
yIG2qpSXtrGxi5LuQcpOuYOY62JqRKHr8QdlQ2kzHdUtf0TGtxbdExT6MDnMAOhIZhjvUe4piiA2
7eg6Vt5G6b6r66+cLqH8IGVdlf2xuDQPRkTFxB1fHuA+hx+E5yqvK0ctH7cxnBFFIux/emBUziRt
i34k3NMvDYQXUPJ7TZzBV99VxjTwcP9lBa5vZ4Mg6SvaBq7G0mDSE6dqqsl66gv/h3JLpXrQbbwc
3SPEIX7/Cgy5EKLnUIOpAfBMIuKYgV4BEen17ABKrFDiDAbOM/DySynGB6w0qQz/t9A2DGzKJ7fB
JLDQ90EUaRvGc3rbSJ0H9M4XH1gdqZB34Wm+FgbWj0Yk/p1VzbxaCElaC9IvT6f5lQYDQgDV50Ik
wplrozN8q59sESZFrwR5Gkto/Zciho0JzGY4XEnfyFR6N5L3S8i8N65yv6Lq2HHt0lVD08QxjKC4
VYkW7VkhT3IhMI2W7ys3iXdGp2rIxc750bqaignLe7p6bqcouZ3XMA+G5gjr12yYMSZl3FRwZ7AY
D7XqmT9tzSCiox/O52MKH3IyY1ZJX8JkUT+jpfqLdjrUArmYJ6djrkqHJmmr8vat1CDiMbs9ceLQ
cVe6a3iqh5e4rz5lxbkWwjMDOchU85Va/+7T/2ymffnrqB6BeyDyOxAbqL/K4c7mdaPVBWN+NFDC
vHapNH/3+1+FW0sZKPzvRQESQcu64nZBgHzI3TS6lKMd/19TPOF17IRG4Som+NGVXhXq9XQcHQUl
ghQhz0OH9Q9oawurRwE1jQbHl66fA35HbgohmNpGUeQ+kxXarnZbg60tQV3s3DYHWPcCrM5W7ALP
swQzwWy/DEQ7UZjDQ1Cy46ywjH4N8IIhvJ9zhz+RqDjxeAwaoMpcZK34eN1FvAryUr+Nyy4YJ+/X
smlrtSNQxGUJKuuKCSQT7mKFKtDY6NPOeNtkklLSkp9fq6XyftmV0JcAXp9V/4YCAyanwd47itPL
H3oSdKbyglMfJOZ8WKMmlqrtoKGGFCBguz3p5HCyGjMrL9fAvOAReJs+mJZ5jaZvdriHp3bXRPSF
EBGZBsfrlRDAKEB6i9c3m2gPnWJ7nXXFTQWZyr4I4W/RWPdj01J3bUXvixqbsM3UkbTAAhsRLkzJ
AWJR2Plo2JpT9N9ibAo6vWW7aJVrAAiC/9yB8IsrQaZMmLoPfVx7RkhvWgACPlStHxKWlX95AyQn
0DEE1qHpwHOAs1VP45nXTb+bNlPjRw7D9NTsRuae1uZ+uxE3ZxmErw7RPQ1HQe0sEu8v/3eGqFuQ
TOZiAXOho8E4zMncTwxsDW8w0Vv7QKwS1OP6l6Ty5rWz7grW11RqGNvLIm1nVyd0K87+B2x4KPnJ
NhHf7Fa3xdQghnXANs2JFhO86WZ1YhrZvlputOUm413S0VdcjpzcW4n87lCaxWOUXtc25tCdanrv
BSvPcGvZ/BBUZ5EvqoXryWaRoD3vL51nKn4z7OfxeWY2P9D9Kw2/ys3g3FRP+oomkwrqrMwiz6UX
A5YctVjW5PbfOvpYgpYcCVpiJQFB0yFW7vYrP6MIgiFytiR20irBI70WsUcYRajE1VPg1hDQlzUt
Ib4FiYqbqrR6gjWcRXXDYbjv2S+gL3hGbR9uqpSTpWBVbPtCwpstUBaaVoIvU0oHpitfU+/713za
aFXqjOKpPGZ3GUGDn3JXYBhZ8Z60qSLeQPaL3JVtZQGY9G/lrWZ5cuFro5FP0Ed4diwmL06aaQhF
cP2lD3Ns0tX+vRyUHp+QISL4N7Xj0f3CGKBLsppJTounhawNsekX2ErRX+uqSVBLWZ/xZUR2iBv5
WfXBaWvql+5/2DXFCPcaEIyT+4CrKI8qXhuceFW1abXOvGQsv3MVwAQyzr4FSIwCBkk8dHpFNhIV
ZgeGdMs1hq76QLAoOV1+Ik8YVg5ymBYB4s9AeIT2kkY7ZMtg3IYioA5b7dPiMpPdtfjy+OZA8ULp
I/DQsifKhRE1SQCzHqX7wR+it7tzE77KRfB7Nxyw6a5Q6f4FsL4//GcIq0brH/i2U79oTzzvgXaL
SUN6gXlctGGIBahlKBF6bp49vZdn7Fqv45rygFDhfVQyg0gcHLI36YYQSyNSnBa2QiqqmnnSrLkf
liTpP0NEtDZ5ylOyY4s/sPasaC0dKSCfOcOyDc2y45ewJxJUIUwqV0mAApytZCAfIreLl4EVZLzD
ynH8uDeESzBxecVa+vfuTBT6lLHfFU1MPL5RelS7AeSzXl6Mec0adNoztWuLYFAk3gUtiemU5zBe
ea0Id0BhUZGuj8bEs03exRQ8YfMYWu4EsuRFYpn6smqP4zt7Cpn9YD+Vse6gia5Ar6K+5NNKUQCn
krOMBkcxjI11yA76lwz1O4FvZiyZpkDzzhaB4NsraNCay8n3IhZPnNkXZx2LXnrx6+NL6VWEypTo
b/UF7amL0fG//XYTc0tXdqZ0WquX8+EWYPOPAT8hWq7x3XxFYccmKdS4eXX8Cez8J+2LLjWMpXvf
IeW6pTWXo8oQCEP3Nr6v8FE1FmaksIxhO5JnxfyDolTfYoyrD+2WYyqe0OOl6kl16wazEprYN11m
epClMyGTz3DAbh201j+6NyNXbrcu824qRV1gqQoJbNUrMD/HFLo5BNdYoEuD1fConiUFX6UAF1FK
3k1k55sLQ0/YkUaekdtocoKrDb344Tlc6oZ9G+/IOIRlUMmzBXQ56LlYyTsvMjUnxCE2lIMgrjhA
uIKzmR6h4mhhkwTU9PRXwZz8LZ2ygzK5yvECuOaVoNSIoSMo75i+hYGoOztehQ/6N1kh552PHeTu
emLEvC9TpcRGxQd0sTPO606UhIuMLjiW6qv+y6x5ZyStFyEkzGJ+vIbuoM+ixWrm5Vgh/ipMMZ/j
AwzbcN6y+FEatoLGw9yOcrhRq6O7ngPtC4LID2j3XTzE6uPIY8vSCU3rQmJEeLvL3oB0Ae0LIiPB
qiMQdJucPFTWfJ+EBcpbNpz7Y2hnpvtwETnse3z5mWY6u1x2+KAw4bAuLC4xkRAu94wCNvHDBPS/
fHGLhnC5gQT9RUjaKEVbKwhlbi/sZvgS/zzg7uBlrzvYmZC2ux9Dj5fY9YCMTCcGZhm/vGAMKYc8
xYFAMSSZ+1xMToKz6T/XHjZPbC26xLszvw/LVKB6QI6L8SxJPG09A2TFM9tC5TSMIKQk2eKA8JwE
CfZFyknOqTwDzoipppfTDPxD232AcS6GHzYVHlD9WM0X/mNOhwG8utpmfMITNsKggo23gb5nf4m4
AjznYfFv9ZkUchqC4mal+GfHC2o4OgCBF4833+l9Klx2Nkc3P9IEvRNeTuPwSLXtCn+b1N3aYSWi
cKuGBI0xtJxxBkyu+G5o+WpIvBLa9pSPCv6zi6mTjbv2QLHB5vs8gdmyGn6fxXoIRxdWqiPVvXG0
1bxFsQbb7RnDsrsijEhOOZ36mWjOcSpbzl02ytRKuEOREz+KiUU1mz9fMCy7Bfj+gmSLCjersFG/
MtvdxkxC41goVy1QUlnbWjog7ZMCH8YFJ+nn6fu51FJutn7qbZ0DbzdFtW/nFBWhWP1Acef7gvPe
XD0mku43rw/CYg7KoJe21VeLg41CubyOYPJkT9YQOqjS8jYT23eFXulg5M4YgnUuNuuprwTco4P3
zJCkVTu1KMIakWUoluBl4tyosXkjbg+eqO9/7voRmgpJviop+HwpuG6mqBEHDoscffjEBf4vsFKn
p46AX2grGo8oe9d1SFRjcUHdrLsmIPVs2fQYziuoeJoiB1rlEtenAwmMEVKnYB9MBdPg1XkuM53h
0tnn0zTlUFxFCBJFnsRVIlzf+O1eNRdJwJA05nHbyyijfjCCtsUteVoAWa+ivuAyr8pllD/U92W3
Im5AajyNj1TgGHXlsCjdGzti3s2qfWrlnq4/ZsmycuvIZLXqxql0rWJuXFuVFgTwzo56CM95OM1/
CxhZBAnfnUKQYnjbnRJfVwRYNlSdGcHjLaWoYMtbGBud/2Cu5OBcmw4GzZf8Xtiel2s9Qffpscx4
LT7V0opzWn/bNAJTWOjn6HFb7Vy7oLNO89gd/UC3VAVhl40WmrEqXYX+omQAKXS7D3sW9Dno3C06
iN0Rl4pfxPAyWfJmexqygMC/v9jQeWwYBlkTl6qZOZ8q2ANiUTiYhqi3/cttJugQTN0M0625cubc
Ip7tZVihTX1xhP/kl2SYoMYgL+G+tjzfXtuOF7eiAeBo3PKKdQdgDn5KMs4Fdz2ZOjabhOKLH+01
Yore+BqO0axdtMiTrBG45U1jgCthEmLQ/S7BTkhDxNswPIjIavbNrhHA9JGAGpFlwKXxF/iKpVVc
ajmupbXZLE9EtB0m5+X/UMlV1XiVNQSgDQYWX5CztAIJtqx6Wzj4dUJZpPOqYG3Qmk2263tu8uAT
v8IfBj+yBJWLXhRy+H2hMH0onOBQeafU1KhPe59yzvEC5bS8/s98eGjxNRTF/XoBPVSpD1nF/pfL
ICcfoNw1EdqOcsgRfrp2Y9rFtcqT/PJnDhpNMUFW0iPaZQYJ2dfPzBXe1MCFzjTnCnauDDKilfZE
JbcI/oaCe7aaXkhDzAXHHnOgq7sc0pSllguvLbRVm1UvWGtcitVP06Sv+IdfYfg0qNijy65z79gu
VSSwGTbmjCnrIhYBA1+4TJ/NDcgy5ssntFLu6ZpUOXQU7QihvnSRTl2qDs7AGpOKiAe50SZJnAiu
ilSJpPGvOu/8pUGRruIyKQHj5s1ST/I2tEy7PU8i9o+JHTUDyzOryu0CtC5draJoFjz0i+OywgH+
JcmBUGAK+9PXD1H26UpZhrpJ2li2ggTZvqkyTEYISayi0QHwoexQBZ27MnLaftoXGjA3DSLrYtcx
TYxE2Tc3EiabNG6k8ingBbhssdwsyn1SedoaVuoF/IaTA9v1DdenE1kBRR6uCZqZMqhHGTphAWC+
W0sngbFn7leJXAxysOgJ7iOIYFGGUUsN8dR2uqUezUT7px9G6q+YPKwhGt59iZcWrBOVFKYWR67O
PV/KZVW7T+8cQxULdXO6n0Rj0SPiEVhj47NBRysvnnVcx3fhFNJVg8RjR2HL1oznJ+mKkKiQaiS+
aTAWJeA4A26FYueU93jNHE2ex8Q3xJtFnKs0/n3/XXr/Kv9VDOp4+000Hcx6G2cq9zlW/JqtKyYW
i9JOI+tlsXBobXmtv72w0DE217jzPOnM0RR55oTUdFQ8NESzSY4sOkisO8Qm1Jjat+kf0niig0sT
ON9QeNTK5WrZxPkAfQ+qai9WOQR1JT35G91dvbIyfF/kDyqncEgRBG2rjBQrVPSCIC/ylM2/Pemu
m5ANOx3mab/50aMSNyWudla9tpvm/g4y6hzxTJnhXxxHQXY8M3j8OjecArH4ZLhcEv3EXDybnNCM
pGFotTKULPOv1ctyz1K41b5NQrMhp4Vg0vvQ/gNKHSbe4VEBBNEmQIdiS/Ksd1DPja+sj4Voq2lT
zPW3zjS8e2iiK/Vu56xnTv45QUnO8VJqcTIM0hiW/pTqV6NaUnt42wkZEln+/wJZXCAoXM/s8fL/
6xZk7eHBRvzwsL2tah4Zyj4M60hMwAH0pO7iqzPjfrzpIFqCtWWFO3cImfV+Nc+HMKVNUOPrfKqc
A3/Ic7wufYLNgBNnNnRSIBoS/6W1OomXfQXPCkpBvLalylHcOa1clBmuARRNPh2Pb/3yQJiGc8Fc
hlmk8qu924EnnigQROzJ53C36Won28+kfYcm0Mc09/T5Ai2AGBUmn+tb0F7DyXOG9WJRyOUPncmV
K5bcal+4U9U3nRlRYFHXZwFdK/aH06G6Mg6JHJrv6I1plYVfCloswRbqaTEK42JK95R+rP0zAhA4
vTVDft1kzBLXPW8cdBG2krgm1WQcFVZcgy/xezPFOCQ/V2LRFc2voznEgcz8Fdc0kQIlyg8lJ6Hv
vdQZkmsv6J9jUk0sHYBlxNVzHuDLzM6jAN+daCNouPOVXjKzx0INnrW4ZYr5PRBaEOTS0Z9wtJga
C6EOlpWoUpq8kemzbZg33UHwx2yXKYnvwx7tyF/qUU1PnYO8XQNnkbxGcxML6clPaqs29SZrk+vV
ogQcNt+UjeTXSP5/JxS0OYDZ2TMOSyDfzn3WyVwwGy5WXZ6FBy2qveAR6M/k8pfIKV/8QOGQS7pU
jYdzmH2E9RjR5XzilJBOHz+lBTx/W3h3U91F10n6Ki66A8PYNuHOWqm0kuZraWDjuTw0zXQhr3W3
IZYoOPTSXZbu3cndxOkaUe5jET/InT/0h+MkmNINHBq/ttoRtxsFMXUSVRR/yMGQ02mpncdovd/p
+Jgs77DBmwG2PPfSRBqxh70rIgevgsZtLNcMAwDrcNPdUC1NMIya7TVUHJtlEFi1m+YQ1kHr9j0P
Wnt8OlnFSr3sGMp4xvQuwztKqRpymaBhB3uL+k+7bpmez6IP4bC7oqIjFj6C6L3wu2/0HSd2hhQ5
Dok3PO7cPDlsoygnQsOH52q31ZJQpjLe+JzWVwUH95j5ZDm/3LYPKVsOV0GFjVJaQQNQyNm1fmsQ
nCWkDI3+XfppCuSDe8Zn7Ybfdf8yfBc0zp0MjkcPYL/yvN4pQT6n+Bo2QWFZ0xqcYh33GSNRR8eg
BTgT++etZ4t8+La4prHSNlwdZwIFq2DhxkESJg7H3k6MEBWirrtDN3yP4gfFoqoXGUPrB5dVB4yM
7DPBltCOkJ6tEz73/jaSl1I4EjHzZSoNERCmb96LUoWVuzFrRYI5756HRoSYIWSHU65UIX8R9Pvp
M4wf++Od45/eyfPNpi4ofJd9q6VXnqeerTq/Wp+U3T4igB6Hfr4FDg2Y3m1nOcjAjBgFOjlT5iXs
7sQ4SxGFXl39V2vpSMy7XTuQmvIkQXRqex4RdAIQVe16tQ3pxiQ4Bp9nazcK/en/fcKH9oG1ecgh
rYaKLYIB8e5Yt67/NheguWIf+mFmH4/hreDrYTMke2mj8RNXd2g+A6IPA18C29t8ASe951e84tTQ
HUqyxB4Y6LW9/zMgj2k5RjHkVxyIUzzS3SettKvBSY+1760qsoy86g5j6Xx5Qt3b7sWzIdAZ7ch+
lZJ9NjCH+wK1A1mkGGxq+LJ7MByjN2UyKwaldqA+ppJEfDnSWhNVmi2wmnbQPGkWa4C2oqLQs7ac
RlHEzbaBPc4b8AnIMFalRpwxgd8k+zQ6EdLZxTdRyPpTmxXc8H/TrtKBhRoP49qs2VlJBrCLOzRn
l+1ab1xs71PNZkVJFL6k3+0SStEHmsjCIJssij7t6Cs1TVEn2iU0CSSan5zX4IGTj1Ot1G2fMtU6
H/ebMgQPvdiOTo8k9Lrdl9ONFKP5GzusIiwe7ukb1EyB8uMd+bvo8U44g9Ic7eB2v5msimULET9i
SDHR8YeXY3X3uHdlM4qr88J9Mi2MNVwp4Y9M8tn0iZE9fJP3hSQ78nsj7NWlCmOk1/F1IaGWRjG+
aPIE0/Kw5KvvXDWfJtJLjPvN3gcU90L9559e+M97v2FWCoiAi6SuZUteITIljIgzflnG1Qjcc24+
zJb2MnvCXbAj7csa/EL8jxFXngccmOW3JJc2CCwo7+BJKSoXIej+o1/eNOxSLq9LkTWbSrxLnG29
DLCQyhB11gShC95zEo1asDO9CNQTCfCssCJ4hx/CUf20vH2sSaAt0anjIJrVhL+iuO2fsjv8fnWG
A39yo2jDT/IfSX0s3HN1irSzZoBOllegvzcIVYGoP9rycKrpZThneMOqb80HzEKzoDSs9MRJ5M5R
7U6IJTSBWC8/Vw74Py4NE5Uk9rlsxatUAyqj3RJZ4JwyADnUWXU0kk6Y8LcHiW/ZpFhNiRsoaKu/
f9hh9JIW19W5uulmW6xHYrP3v8XwyAcQBtQilN8YVpEk42N0KWBgYRv3zF4kKlhEB9t9eE9R018Z
XaPZD3t0o/HOCLuns+Eg7GX0y1LCIELmAT1oH7Ru2oCAfBAFWqHB3EpcOE8h+oqVOZ25tt8ym1po
pijqwcE6i6RBJhUYsz3I25NXgyho+/6lYFNti/dEvcemQ1mEqmUlC4EP9PqZ4v/Cv68Zg8Qt77dQ
X+BaTR54sOO/W5st4oPk+qTWw3K/V1DFuKjk3momJ6KEEuLceUeSDo/4NQX1LBPKOnXlnsAqBzEE
lyCMfOFUTijA9o7YEPzUmZT2dvb9yhqkey1H0vWziGgmDFNK/mEsFtne9hpDkPDRfMTwDqnV9S7B
dIxrSjLB8ObtcLifRZYOG++xxNrDCwCghfoDFw/WdwJxDzb9DGeRDpqMQS5ytzxSE2Y4TRDrZpBL
kr+9r14efPFF0t6S+0LYYA34XARGQ0yT4A23PyFhMpmJ6IiBRXdA9YVOnGPHxu6NI7/BjOOEvfH+
dJ0g1NszUZmzWdL3DNnXOWTD7+xght7CDBDDL5mJCk18cjYVf7zR7grNgcvDXP5kGzLB4QtUcCAj
wPQkc6busMGp3W9izja35UY66u25eNk+Y09PgqIqIFVT4v9ILkgcUT/46WGBbPl0HE+tbxY3SRaH
hbsX9PcqykTP28ErCAWZ6I5EfL5sNNfsqiSRVYmEyRMtxpWPFytZGv46gR/4R0PL8Pr2if1ioOs5
A6Es+x6LrLDahfTiy8fujRS7TTJ9ubwTRW91c5qNLxZCyPf8/Z3nWqMXsXkQcPkvhdTEU1Pjwvkf
XIZWPm92UjDXSp3R8c/SvPQ6VNde+rBwS8tWexxnXPe1P6oij5c6IDohlZsmBhQ9m2v0dtGQSEBP
ZYn/fLqH0SqnFiXn14ev579jC/JV6f7NDEX/zp2OLAPCmOdDrrwM1U1nO4wxJ1/atbQQA9KnK9EM
vSMtcbDuHOwBzkXrStDh1mIfZjHr845ir+mNcTI7DxeOfVNqoiatDWhQr6xgU8hjCTOYjWtAyCt7
lRpyIg65zZt3TSLWjJ6EfzGlBWsP6J/k+6jvYE36gYyVKGMxUnLwy3ny8UbnFZ6cEuDR8Faraf+I
vxkSY2Ho8snKMqB5+g93EN8TUGdA/ZntyjBLrTvYYPXQzIVPdNAPQdgdd+mquIeOEAxRYeNt4DpK
7NM/8eFGaS2LiH6HXByI/g3Euu+3wiLo3f+SjpUSBNRYZ5ymj20Pjz559AEWxbLHvUMlA17JEkUc
PPCObf7leU9KJ6b82n9I2Aa4IliNrA2KcAVe9zSKM3k7kjw56XI4M8n4RjgDs6NzpkXG+QOBNNqm
8muH9s4z7rMDiIWL4saFqsLkjzwZZmDCCpZRIcTiUIHbdSiHfMhkY5SOVINInLUEup1m+qIvjX9S
FQW2UEn5180prgBeasRGC829MTTdp8dtARvFcTZRSqGENJWQHWO6GMXJ1TSk2912SoSAkhtF3DIm
T3gLZD/eUxEJx1RTY5raGRuRSmQXvwLOXYXdDV/hHJUCZdljHJbNRETbaUN36QYv2A10tSoYwX+9
cyU3Iz+b2SwZY2mMncDah9/q1wDHlO8thbnOIlVdNJoNZlJ+oCyJyJz5cAUsddCi81n3bjVntyRN
nfBG4x+N9UE7dP1gbhboww+C9VL+8dxVUh2hsVD0cxvp3upKtZuPiVIoHWZ7Ze0IZ8UChWbNqACG
GK7o9tCWgtDwh2kh75fYg5bgyapT4MSYXnxhuQ39tLcW7+Fcrpl8jrULYNgNEtyVZV9lXPBWSXcn
o26al/qmuQvhuPJxyG3LfZV0VmMovbDDb9o+9vMmwMWlD+AeZz9BM3IbmkLn1aRE9g6kG7PWka0K
yRGz3Qoy8yiW+vgL0D2PmWSttkV+Zyzoa2mtEPtygrkkMtgrIbNzT9HcVcI100VKClxqpKp8r892
yT8gTIQFLkrVD4cccWPRCZse42/yeht1Q109lco/Y/DB7lEfdx27Sym6AJpwgO6xv9z2149uaMeN
zy3T9I6nKrZnZ4kelARTekF9j+SAZ+W+IaACmg8yD66RL9ZNurEbVH9VweaqHo8w7w+UgANbhbRR
Z1BNQFtWUh30Kx1xfZXnGHucWq/UVVAmyYsf+0spMLTHK7yY6imWPsn5AXQQrLcttuKAzekSmUQ5
CGXRm4dojx9lGZKvjC8lfBPBYZTEARm3Mu6W5yh2Qu/CcNQm+HsOyNU3jqtCZ69KgJ5k1hdRdtzQ
Nw2+vvfx2Bl4iWS1tyvxGTm/VJu1VkXNdx1vW9MJ/dMDzCvkkNz4n4K2bCCPC++2klzY/yvFKcDC
XI9qaaVgGVgGcFCJ9/Q7UH/h8TA770satUfZiR5A6JONT94z29xHKWsB82GWLT+MtEd1zp4Qgi/L
8gicLaAOLLPM+jDohWNUiUl8Xhn54LDi0h9O0jtcXhIeQubZ3USvsWOLccKAsk3rE8FQD+D5FUqM
+ibUsMqzjH/xyQ07vxIRsYp3HMryDs9PwBQgzxY+oYIxaLA3Q6CLNuOJg+1dC/MRA++Z6bxQObtx
v7HfNpfXRRMokkdkRB8Ux/yxfYssaFz/lAugdynE4WSt3p8rywhD7/ZYkX35zTTVNL8fec3TBEaa
uyBISUd++RkBUFIfWiJYixuH28stgE7bV5TUaGU1TJ0yEs37rPev44DGJ+ZxpEZo7GYZgdx0DCZE
7ccGKj7VKMhCd2ii1lrgELa/4GCpfjHcJ5TV47plGsajHc76vFqDnXGIUiddf4/ubQwBsYDMUE73
/cxglVL83NoFdfPnjb0O7Sg/X5lK8ecB1NZJLcSNlB9d8uwrvsyyq0qaJhqEW9RFc8Hxs4iB+eGK
ZqVY+mMAifB6mi0G/U+oXz0/CTsSowNXWLAuf8Mmzy3YAhiLFGlDsbRnsvxkOECAkqhXxl6Wt+8v
YxnOWMJTBwBOBulwu/dHrBgAfWDqTkP5nz7bjM2z8Hsehetqh6CYxtjKAzeJ6xYRvGmcKePgqhl+
no263QQLVJviNDZshDq/G66CCov52tUVWuCdnqZ+nTRH2nfQQiJ1E589KZ1huaHLM1PfvumDPnn3
gNM28BdWlUg/q/ML+DtcbbPu5rZvqugh9uPn0U5as3+Y5RhOH97nq/i1sYDVD86zs55Q/aTQINR9
W1VB3LvGqxbtb32BMHX0UW7tgLSSj2P0WmPmGrB+wfFS2AZTXorzdwkK3tVaIltjBFj+GsyxJHeH
1jy/ZClgNvBEAGN5FeK4cvXDH1LZyeV3egCh671EJFUFciTQnCJ93q1vaNV3KwiTJ0H6whXmG56Q
5nEA3F+l1ugThylzO2bLENDSehtI7QEg8SYHDkHcUcaMUBuyOnHq2ZOFWWKpcjQzrNoZHViqVrDm
+hIpLr9egjTG/vmM8+9KUa09KfYtVYqnEtCYmx4XGbOn40Fu7iijX0DNfKVek1uic3JCRDtxIiD4
rLfh/PK3X38jTMI78KvHyZ1qJdbjrtg/a1gUMSUYAelkxrx/CW1v7SUKUtLFAui9SNDEHUgiOWUE
O/7C83ifQNcxNe968GvUVybrjQQB3qM0D8hG/ugXl153ThNls3k9FBq6lHdkHspZZ9XS1MrE0LmP
IgbMYyY6C/IRwCUpkqPv7pO+F/x1yb8RczgLbzZiMEHdTA3SLOlb5zcTbzm00rv5Z1QV1kcx2DEd
z5tENMD07qBUuaT8WxVDP80AywGg1vo3H0X7LGcXBIZP+zfatzeaP4uhloiDZBkL8iTfVGDA6MC3
JY3WFez5FLmh67AE9pXNvw1bWjMVHndpuXQlSRMAe2zqsI87kWAZMGAwJCq2gLodMBrQAaJeU+QK
WGbiTgAYpUg2n6NWgSgL0qQFWwxO/bQwjBQDIznlNdiYoK1k+bDd0M4EeVqICRf5Ut9x5izrQjYh
CN2rrP0FSbktpeZj+M44YCOcqAwvf0C3SQ0NvivZ/SJigVA/O3bNWwymGKILS2VF+s9jMCl7Qbi/
TvxCwgJB1mBSvZ+W7y++Gqd85++UFvzJCDFyrRcRChTEsFkTmJ2Irv++cHkDD5ersWEnHABwy4EK
bQM4VjGOoIrF4GNJlKs1exhH8JYOgCFwjevro30aoNHbuhGGPqIEFH5JSK5Pd1o9LYhxY1B7HXBO
o+qdg1XzKxze0U0ny6PtoGuO357sYYQDu+rbA9UqSxYFhnMW4+kd9GZ7B+x1wnz2Yq4S9cpdmVuc
Lr9VmfU3MBxoses0hUzWKTqhkfIHFdN/+uOG85GIXyviPJelXd9URutT/6G1RvUgjMKRbSj/ESFS
uMqruGgOWA79/zDn+dNS2vUwLw6UWuduksUdFOo2beBBXr9dyMSIopH9m8g56oEwxvzSjcmMZr16
eDzbIaYedmmMt5ETu+LAdenqyFkCWOp6QpD1vr/gJ41t2NEZSoRmU+NGNXGf8oRIgxx6d7iyrLMl
bzWjWxNSaRI/FBTfS4d0WPammqUDbGWXamlNU3hSPdQx+rgH00CcduWghq2OGZj8dMVYBjM0T0/Q
ZjoOet7ykU4fHNTpQ2PI3czEgysYIgaFtJNy8TpoxURqBpjn5FObmP39DkxR9aLjtJOC2u4L51iR
9pbmkFt1bYQX2vVTW/mHpC1N9KhhW28O0G1lRNZ/pkH0DVUN3NLTdFVr+tiqwa4SXO4UhfD1lT/T
9EYyN5LR/EPFyHqq9QKVdKNBUCnXxquxHhy3UFWVbT79ketm/UXr/8AT/Z4f1x6QUIqf8bXIKhR7
1JExZB6sQBZ9tPCu1JiciLybUskKocwju2Y1oKjCCDIuQnKep8A5aoxbPKpgtSvxvv29PQgn0pKc
SaqrFJM1+oaiXL9M61w7cbEOxs9P7J0kamSL4EViT9EDN44QZhcsBLl+UHHsV1iT43RKwiZ15v4z
KGHbwX8NPG+pEjkAcmNhFr7SOidKVSDHxIaBUVghLjy0xR9ezNMQQ2bxsD3bgF/1Un9UDh4z5PgK
vNvMPn9hz8AtYsLl1IJJBbMvWzrroyOrOorBEqKbx5tm26KCZY1mJOuX3KPOXx4vOTghW75z5cUT
Uk/Ede/zV7x6wXQVkOOx6ixZz/3X4hFejqFHbFNoupWwXhGP/UOzEzNERztu6DD18ELFLavKviu7
EH8B1wxI1ALe8KS2zkxR7BTIMLifLdkLeyH0kBFtgCnUh6W5B5wegFGyAJSgFF+yUqkLDzBw92kg
G++lg9g3qw71dNC7WhLKFRMU8Ff2D0MK41pbm+SCNIQ2RxVjk+cUPyUiiVnhPfoHh0ch85mffMXO
UErqYqhQZjqTjQd+cr471nu8zyfppu0c5kF3/MTDHvihI3faTVkAB3oWCR+tI7ukhe5XaD5ruXAh
97Z/99EjzZv1EMiQgUr9oSjJgFgYwFjO+LR8G8XPBGvTEckiU4QJ58CAmIC+yZyjUQfRvjDjR0MC
lN/U3+tsDP/4zWEQDVZFtlhk0+2dd5Z4rBIHDIr/PDzvGu367QxpFGZ2ibnSjvuRFGR+Z7Mzekc/
nWcda6CUrAfj00eyqoesBQznCcd4m09gGOtrt78/50rids9P5LWDgO5A4tgbcxMSd0myi7GewG0G
X7aXw+utZHVQ4jJz9Ey5X6NdZ/IJ69+M6SlHSFB8nw8K77fHkdWh9eajoK9OJo8C+BiEMo4nzLqh
aVLKcYOLd0zimALyQ9MiedFqoodcTo6CDNzaNwCbLUfVjSFySrZFyU6BecJl8rgUVTVpJn+Dcux7
HKdDfb7czXx57x3Y2tJfYzF26bae1iK0gHeqVNcoxFWNqDPwJXQz8YDDVU+ekKWi1VdqKIz7mSQC
r4lt9BiBlO8UofodelJzTmN6JKvj/uoekFx2BMddbx7NCpZxQVCr8ZGBYbppsgvkkdQVN74NRP16
cxyNfZZIj729v3ISfTPAof6dJVYRAbummP6Ug3LGDlJO+XGuKC4T47aztuQaJ7gPuoPmAFhPYVn3
jjBwtYyy4uLlrmcIeVomjQv3oqG2K1CT+fOjV+72sPrZROofvfK4KU+usWEZhwHCZ1XDXEYwlUyl
fG1JHJEXhV3f3tq+YtggnUj1UOpVQG7UluJAT5JYsDBDVGub/z7DYYbrQx2yZ3UUhzdXyuG1jF8K
9Wtb6vQeIHt9Eqq+4lZNsWSCfToa6bEKhblcfeHlyxZfImNF0iNjeldkyBPMP3Ww50+zKd/OQ+yG
h4idWHuItbPeVU7XPk+omaWHBDX5Fmb3X5EuXnX8ue2ZNou4nHHo7P+pvdGllqo8yD4zCFfM6G/X
3cDknSAE1hn213j6FNUMa44FztuWErWshQLz6lkUGakneU3bWHTaIMLSibqhX6smoMr5Yv9kK2n6
AAR5sfwWlytCsA6DtUxW3N+UmgNx09dBqaC40xhtNzFyWdPWTfemoAg+1LJQ1D8YNSgPHzAHhOBS
Ncx+SVOGFqTJP3DmIm1tS4Z8uAkXxrrN/Kz5n7pnTxhpWcj6C+MdsqYVc+kw3bD1585+qpGoXoum
gkkIzJY0j5L1MRkwOWmJZqsCs/Uq/l0FQV7knh5GIML74rlKfxSp/xtowKudENMms5cG7sTbuyab
JVAJpA2lZi0Xcj/S04yCtt49HzCHqw7SyBkMIU+4z34wpg8OzU/UZGmak+HLykBlrZClZBia29yi
3eXsG/twfDdZ0ObAiKBaASjCgYUhG9BfRFES8/ugrvJ0nlKqGc+sFNu67P72Gj8icy2cGuGXPQKP
lWr9m+ijjiUtmV05p/zr6zVsNfFYRfqwwIw3FiXs7Z5RudmvVTmzGVK22cx3c3KkCkMAhxIwhq02
nT0PqgwbHnjLKF+x26ibQAzs/zR6ADPIGSapAcAox3MOKkkxXYZRYJART+ODNFpmq0XKLnTzgePj
U0gbzFHE+ZqVJf7hZYtsh/2hpuiMEPgbor+oAwSsRtf7ENLdpz0zdY9dIpX5z8YhkSTp9Dann5ZI
prjBrxg7TV5jzUticdBP1HAlKGWsaJn25/i/qI/oaVX5EieAh7OBOsZDtGX8KWQNiM/lIusOvkvM
F0zBqRnr4osfiSADQKWjI2WmEyBjw/pTwTueswNg4plhdmPPEfFeg5rKEM2kos3UOagdFuY5/RWa
JTMDIVKc6gLqn/E9F39RLboI9nk/piQ6k5exkxrBz7xvW70y97Wd41DopIer5xszITOslEeFga9+
cD6Kr7F4So83S10x+aiQWSHfpx41Q558rRaguHjZ5Xg2u94g5dyP0/pJRoddKx50VJ06AkHIJ1Fr
JOmypef4BTZyjWSOHlDz+9TtGN2wwCSMPeaZmZ/tlqQnihxHL9ZgWakDJxCtlHX5cf8NiMb8aQNI
IAAuxLlZfCTrlTaEhupCudsmeV5vZiDtC3BDqQgNW/YB8mzy2B2oPE6oDxoPFHShSoNYnChzL0wO
1jWWjBjplGKsKI7mMj2z/HTmdTMyWMinUePU17D5hfcZMudcPhdBsPwpyHeYrBTBuVdkvsuD/Is/
mKORrVjlf26ykVnK2PCSeKGpEXPC5l1eKI/VPUavQ0YMW11jdAUkZNPG+JEqagzxQv+XFqCRaz0Y
1WivYPZ75TXGK2GeZetAdDhkiOjOz0nPF11YLfWMTCjaLGlOsAXmbRPiyvxMddqtF8qiT9HfC1wW
4uSMMAJ1XlGJbzdAedU+mqmX/I0IWrePNUyPxLEdCizI6GUG55+8THVlLQ1A0HkHvgF5idcTlo1d
38iC74IVSmE/hF1mgwIHdKsPhpZhpTVyvvUvCFxJEbHjDZ7JxLXMi8Bg22kc0QQ0Tv27EgEZAW2E
79aGdD0ZTMIQ3nbmScn14k7Uwzk1G/CdWR4W4jf6F3m0rxiF/jAFbhx1AI04cm7g/lwFXEHtW8AD
R0oH1hEp+AGdlbnCFpFxcMWW70XfoG0weaJAYjsBgasxC7fM1/QDH0HrxFk4F7lbNZkd8uDhPgZj
VQcqQ34FeW7lCX1mSng02W0vn6fIhNk5f8dL2s7mV2hCEHe3QuKyAN/+TupXjlWrCGbJ600Amdr/
iNyFgrbf4rIaZGHKFwTZdCVR5DRqvMntxnRQA9bWhSwgXtVBG84SfV2F/1MkIvgZu3CsiDDUTKKg
O5YsqC5t0g5blKKPL9ZCvmMaCpEINOR71KSS+AykZtwXV4s2nrnZtcugq/e8/EuJ7U96OIAoA0HC
4e8SONeNUSYz/0gc+MiyVLbaeCiuDt4fv68O8BGw4+OPytDfbA+eBkptqoDAFnj7x6vcAzXj399q
6ujD2YE5JNjbLKxF1kDf/GWJXp3JgQeoPCUvG0MDrVMtVyQhrA7WtMMxnHR9t5ojJAk9XnQdls/j
QN+OHfVF/ET3BCnJUKeM4NWOBxMDv2CXwsYiQs2k09jRoulnyPFZ8X37iPOLDgY91R+8YNwxN2/U
BEIIyb5TP42gXK7Bw2qDIOX+CTNBG1dyTWnDpLKtQBOtoTaMHg+OVh1Zj0IwJ43+PyO371Nl8HGV
WQ7dnF1E+ekJUjL7vKd4lonq3ivb2HyiuYgPzXoEDnCnhAYyW0m2ELdJWhXZZrNSO7O2HD/eKUiM
BPeLbrt1Jj+g1S/6KFtnJZ918/VkeMmliDl84syPpL7zM3CM+VKl2Y1O3SbJJgSM+/AMRWejbtuW
yhHqF4jVGfthFcEoBuFRRCeJY5T3U8r+uI8zgCyIPhKDRzfVcxYn6PIJhY+R9b8wolEPVBDR1SeS
UzCKWA7/X7vphTgxMf9dD8JO/arYcaogoIhKgbI0HLydNAQdnEmzwPKCr4ytUInbjyt4VzvSAVmr
g2qwMoPXT3202ZTbBJsRBar0OGhCA3HLBqvrq037rDETMFEqDsVYtb4vas332ugB9opvK9W0qqKq
OPxWZiv3I7C55APhDCPjtOr4MBmxB8pdCGoUiEla70IUq0aCgYE/PSHDDxFPsZJR5YxgmynAqs6R
IUbD9/0lRfZNcV4sJjYV227M2qp8UpFOAOWi3cQ2blZsSOc7lvVTAJZ4/E/dxYdcwghKlKuWy9kJ
9ycw0Ekb+v9iomqcA+8qPgqQ3Mq+186qDT6J/ejIbPUaT5lr3vWobmUXZWrLgDCFdCpJKcShR99K
lFssWJa+r/xNoS5iXYQYHkAJs46uBOyW/w7Ktw9tfOGHukB3DjarE7+j775WEYBoFdYBLcgiQ6i0
0AwUX2F9TguoHszULvYpPChYkrV5eeQFHUa5iBgzbqyyzgkcmrcn5LvnxMMdNJETBeLkt4aN3T7f
hp7q4x6YymDY9ifkUL3sFJ6KXNYFUemWxMpL4ra1Zoqr+hFlXavWTueOH57k6upQD3lFPZZfi82u
c0PvVZPmr9lyjl8V4StxjJSWDtf2CcvIEJS57qqVmi4lAmSuEOkKDQmxBbk8KD+AEiqSjXFQU5TX
EcmbHEmMqbCBiGlc1T5TiFMsLFnYc0QDLEMw6PNut7s2VEW67yFL90K2igrcuYEYzFtuP3gitMIC
MT2nck4oknB94qIGLfe5yPqbh47n9w1l0us/lWhX2Q5bBCMo4p0FB8fapBnZJPByztYla6zWVWsB
iX7UjVaXBiCC4N1DfmNScBIlK2zFEHACVHqn5ylNYue+8W9kF7mCu9qDO/kN6Gw4ISGltIXb4Rf/
B6UxvZnoo6SphCMOqsV8HE2cEMpsuwaQGcfya3cJ7VJKX9dl4s7GzKkV+oZpO6ut9Ur1ElnVzRH7
RCnqGuPlOPN8Cm2ryLJ5N7cfirrhcdW2CJCsbUcN6n8Gr3U6xOGOEMiMpCOO7yXaa5H1/+pr/+qf
s0WRCl/e3nCBahlhH27G0yOFjFSRHupyGp+elpZgy4ouewzoNagrEUKJhb3AzSl5eNT+1yxuLeY6
tfsIPjOm4X469AzzZTR6aQN5h8IE1uc/vDQJq0HbSl0ljxBMFYE7MAi0Z+71n0LCG91mc1qRE2og
GxWb62f5tPFypJcfUMP9HZLpn5EE0YzL+g4BSFFuPKT1xqrQS4QfAPBtG0sI0t1W/LRKiqkxj1MR
POCvpylduG7WKnevczPTK7aneNJjJG7+SILYY3KOxl2DhNrK2P0TXlD4t+289EwYysz8FMPfAiLQ
ufKrllrKYP/lHH9sZn/ImdACul+eA4W4hHeOOJmPa2UYFeBc7Sf8pKGTh4CvJBrDERBfudaBSX13
BZhEWmDwifcJJuf8FwGPL8vIZGwWjfqEMUliggTy3E4W3NNCHVLfUT42CaGU6tP/nqOYjIZzErYM
HtysPR5SmEU+kFpHVlLpfH0cBJToRA1LssqvyD9i23SGtZOrYngwKV8taVhB0oOT/iIbgEKZnhs4
RZvDwIA8pJUT21VyjhSGh8RhGR2Z8NewYdaVPv1bGI/HKmFF6rweOK0yujoR3+RKvnzYfAhW63OF
QaZdnotzERzUCrQj37+RuVr2u8ab87SnZIILvW+hXKChPkSoop7BfcKejbxz4P5ekvAa+toXoe84
PVqGYPc10CNpY9ZdtzGCsj094prfc0APwrIPMMRjJFbELU4b8VfWc5q0eHw2turJFBvDHb9s4Vqe
aEcC8/iawhVHWBXe6Dny8LgzdrOAGBWV3vX07bayHt5n5aVykxPq6l2Q1mgIfFfbLmmPzOtCu6y6
031crQ/HZr9/2PWuJd1VLhuE4KUDC6Sv6FzWfSLBLXtxbCFqXXl7EIptUQ0nu9w4woSXGhYmWK+V
uFQH1FPVat3C5cCkk8PEG2/q7Vk6puQfFzI4sZA2ITuYR28B6a+MjTbK9+DudxxEBzlDBeButaGk
8gL+iDdOZCdyQWI/p1KnhsbNBMWVJr+5NdlFJrD0KnrN8hNxfJuGLoqY56kpQ439+U/neodb+JEq
x0idpowJKNeQ2asos9EFwLLY3wTYoD6AJG+NOWzlS7moUn5M6gLpdIr/ESBXuLDOmHFGUDEkPuF/
NRC5jeg7Z5g5S6tNYlc967bPWdMi4JI95+iC++gjETDOC3pwq9+uGDBGh941TNg+6idFBouWfyF9
PVvR9LYygFEiw47ExK28QClboR6qgb1pFlAM9Sj9wiIly5/5yVKu29T92oJbOdT9L7F56m1zLx9j
k0LAbptHcHrAlg7nrWh6dqPZljc/0pYC+84m354b8LJZWN2siwMEDDilVKiXmNZEloVnDNkgDn+7
UZVfVP4+/7YFDEfXuTtF3x2KSre2PvFSFMpoUFVS1XsL3YTZQILXL2Py6xUE8jkRiKGItvLD1t0x
mPAezHQOthOoetXPWBhxMv8e3Ha+w2ncxi2Wd9fhHPHKmHp4tyHmDPovG/EE7yivjvgIucEHu74c
0KxWqy96sxGK8kbLgDjggIFBmTU/eHc6fg44lu2G09QYTgx66R62tJy+KYPa2Kf+402T9qD944xw
Qaov6id5RqOnm7WkG5HGGfDxZg+6bhMo6ech25P9eEPINTPoHe8n9ZBeYlqCXhdwBiI/3nwUlM5S
VJ6wS57JOKpR/WBmYE+fJbd327tZXaCEp0aab1NFehhtuRld22oIsCc8FK/M1oXfbEHOIf+cjk7X
nC+w+TcLb9bDKsvJqLXt3QUaDm4WcOuSTfc9VbhPCqgQg647FfU8ivL0yTr7BYD1ZSPB2karJQyB
OrEfwxxj4za0hFnnVN0W4OWf7TepD9T3L4xi+i6go+O68mA2ZkD/ToxkauMjaufs/vmmmaIQrt0v
CGbGEBrSJselyeSY0SleIbQMgc9/amYDEfe0UdqgwS8Y9xgTIxqWTj/0UA6XcN4Au+SrL+NdT6xW
6TMbqrsq7E66W9GcSihrc4uLo5dnCKb0vJLb1ZV103z1Q/97Mc1aQB8WyFdlyznMKh8ermJF4iPS
2B8rfY9M7zBA2k/3ojYjWijLgChYxDRhUM6GcrTVhob2/FR0q6nULQZCc1GPoxA8GbNjdbzzWHN+
NePd4hPLzCiu1BCHl0tjKMFaWv5DEWI9QX6q6Z+M4lGrLGYAuu3mCNAO9Wuyn12AvTHlROxHHQl4
Zf/eAtVok54DQlB9sFN0NlrwVfkQZXO0/TfgwkrvN4vIFkEEwE/9gBG1DLyHi0OXelpdKrjFJq6y
QNRZkkoaXn4uZ1xs/m/dGtO93d500clgWiCYHFyExC/nUwuiyD2o+MEvAGSkxKyrv08Dke0/ptuk
FBMG4e9kQ49aC7Bud5aXPzN8mTfmDeUjx4LQyplCmSNQFQm7WXXMMOUPVjoOu4fJtdvAcbEYlKNi
L5Dmq2yAKkx/QTjCtfYcJTWwKNz05WnBCQ1lqKas4AsZtnoxQ1rjbj99Mvj5AlFwMK7i/xdGkwIs
RAKiUNMPspwWwPa08kXOahpUOXzMihkH4vhW+Bl02bQ6xYJkvzbiFJx+JOC7hd07CLUEscMe+v4B
WFMVz7Z5oX81fTPM2YayA2t0fiwE9/bfuZmNLry5/HnnICknpqM8wYVyrQBUsyCK6Oqy3B8SzXu7
Ge2wjtWcjYuTvs0fs/6kydlmiR4LPrTsnxNzxisPuuatLar9RZFmBW9964BgM2PqgIU07iKAckvP
uQURsXkIDgGDbnO/Hv80qZ6sUkWbwu9cDP2jYeVeOPViSKut7Cj0FIEQiJdwY7GVpNOwwmO7oe8F
oQw0jrZsKEutWbomHYiMiadeVEHkp/fpG2Hm0SFnJfICHaXZUWbehsfr4JDj64ejZRxnvQsHNx8d
8NEpiqyH2hGFKMWhhrqM82ouIrq8lttYc7dCF0EuUKExncPGcdQLsn3Thj4/5kYulT/lDJUqhaVh
XfI8ZXArvE+qA3srr0e/SLhkoWVW4//Bsz01HttrNuHJUAq7gc5QUdCa8QcQC5B+F5szhsG9C0tf
J6x3bC7aUQxtxCvNll+i0RNTAPmk5b7bJXiNDEkar0uq+nFHe6prv2XgHe5sQ3bkFB2cF20MNRfZ
ksy4UqY9ApJc4jSiBTZdG1gBH4RDMR6rawxH5X7FROh7XGucR1DrYMGAZIOWZ7uWqTMKSkfsvvry
0/5MvYLNnzQFA04ikqm87BdKHVYi0UezIz8fOvNozD1QI3IdpXH4TNWfe142+P8Ui+rX+pXygaFB
fUbwZm2V5nvgfqJYnnKP7jrHCPLO3sRGZzd7iZsyMIhDIqk45fiCEdStXrPXqiev7GISVgFdaQeB
qs6t4PU+bHflkCMO/XqP0vbCEvutzgQ1Ecd4HauLW3bZJKTGn0OMb1942LF7zr/gbC4Hg0g1rMlx
sveVR5s+0/l1P1EyGFwzvb2ppmnawkM3kaiJucocdIPDWG9GNeexnCOvQnbWO4WRFwuvHgcEnJ5X
YALl2vWh8L93aBC0hAfK0mJx6o/tQGdEzy3tbZIQ7QyQX2t5fVgtlN+tDIIbCm4+51CcnBZSTthZ
z6Tl8635uwTa4puimX2dnaUhlTW2X5KErObjFsfvl8fluiqNT4GH2qF4xnJvua16RyBeLfRlb9XS
sURqcGIVuXCUWqFZfBecUyPW8qPu5qdVLbMdyzixqnvGeQxev0URdlcgKTWqkg5kPaQw5q+UMmAH
x/H/TbcX8XQHD1lLroE6z5bHYbkUQc87uAplfI4HDQQIt1uEBtFt3ZMOPjWexOdLxMev3T/7XmXt
TkiGUV3zGmmUQaq1DQF5Z8yJA3I7JiZeA9aZIXLfd+KLgXK7A+te/m8KZ4dhdDQQ/GUZflp0JoGV
NnfMl7JGQlCFwvGTPaArL0hGNHJ4IpybncPIlsfb/bjKgNz43KnqIsNgdUQ+VB3BtT8dTTGzZRjA
raNA5GZ2uCv+lvxJk15Nd3IY3o/WY6HAGP4PNF+NII1LC0csu9PhTspfIKgszSY6SNuHotq7/WlA
+lvewIMZcm7QVpgpYjhvrcZJZ8LjJsRf6io6ZIC3Z4Lf+DyL5itsbz1SFtinDF2JAH9bLFZf7CgJ
1nH44lLrGbAa0XM8dra0y3LHOK98nATCfSSnr0s9wBt6BQ/SesZzChPG08YkcN8Czp1Deb416pAe
CRPf1RE3pzFINV7NzReus8XcbaXv8Yk+/gPEfMJ6of1kWYpctRopNRV1krpnGqTt4+H0lOIlrwEd
i5NzWsR/vd75Iv3m3UAd/kStQZdXTbSQ7d/jfGKOHJVb/Cz3qZA6XOLhW17Msp6QLZfhdxAw396L
KqQ0bCizgsjRPzXXqXppRBDhfzm//Cs9cA5jrpZBbJTtFSsU2bust3ZrwrUISQSgSGdji9xfKSV6
FN9xHZSNYH+UJVNNMZS+KW97lI3CYvtv4NG0VUTH7AKost6W8hJsRixznqQ0A6OIkXAAR73+hWrF
Yyt7lrVq9uBPjKal+4kYB9nHLNjkacorsZTDrIwcQMtHDQ2adfd6GVUq1A3ltcBxFiWMvM7KkUXJ
Ur1V5d1N5ltM+RXrU23fRDuC3k1rg2tNK5pSQT3SS/xKow4OvbBfaTwiM6oe0SSrCKifOFgHwbHE
U0gn58JVVLwaOdK4+sZGj27T/Nxbj405DAiN9U6+RHYbifSKps52pakDeS0CsN3XJFx9jpUAwqZ4
FXcai8hUp9jFi63scK2fau+o7eOvzqs1udzWfv11fxe2l3ixXBv/UmMEpNT5rv5Os722N83T8DFI
4zKeSNogsyj4iw73QI/sJjys90h8mDl7IJrOXG7zqIi1MovFKt1VWxeqqmEtPpmuRTE/fJG9Ok1F
Mu8k2MP3NgsdaELgF/DuuQrALdJ9+lXR2q9Ehyx2H0I2tRUmk9IEFXLYyXmQ4KOOrOyXog1b8Okr
Sba0QqNToDv69TAfEinAiT7YmCnWseWDBdiS0zR23dsj2eFjNrXoe91zZxJlHfAmszWKWMSNe3ig
4k/x1/wTEL0y6MAy6JSYJU3cKh/0BwS8nbz45iEr0QAFJIHMmeBse9kduUebmTTrBRBJJk3msncC
uiX7KnrrVQ7Ty2/yT1f6y11xwqMVn2345CsP7plMTLcgYgiyWCeUw5DSVIvZMskU1n10fu3KLX19
PfiWIAPN1Y2POr4FB0tCN4uYjYBUlvD5g8HeJQoERdZZX40y1PGvUORTQiYR3dUi0TCb3SAEaF64
q9Z4Bp0cd1zmh824bBR7ZXegx8ho3IrOlAon4x7Nsp2NGemCxIic4hSOHJOg3qVz6OJFP48/KtUh
kv3Xa6tl9uUa76qa04RlTIMug0EAbbh6XtAR+4WTIMys80BF2OfxAlp54mAknqovivOu2BDOBe34
61Hawt2u7+lBFM0J4I3hPqJNfGHge3vaN51wz8ybYoPHcwfbhkBzgsDu8BwoOk/Hy17HE4MHj/3A
Dtgoxt0g1FUngvOZC/DotOdtL829+4ldSV7D78J+Au2LcQczr7prgyzgExpSQtv0H+muEYmcootI
dmLCFeHQnMz88oTLfua8EzLcHw/6N7t+0nqPYI8uB3Sy5GY+5OmBTB6IpJIPlqzmRkJkc5B/zA63
yWtKa9GJEtVBbSb2ZY99O+/lRu4u4dblTx4cFz9NuaSnBdXdOkGexmDUFbQVME3ezu3Nh2Dy9ayr
x1OCM89vUQOapo4DXhzLUEFX7s7YGA2M5rch3UNkXwUql8VRl8eydPaOZFj9w9Z16lm1Fn5ugnfh
e5C45y1hiNPXDFY+QzQeeFRO20ab6+ytxRtThQWZiQ9C+SciGD9JIWhMXVWOlbSzjIEjx+a5l+Xn
jPxSU+08sMjzTIzzwu+5pKrstPhP+VqSCEb0TpFeQUAsg5bO4UTX64o47058FZazhwpEp5SFgh+k
X8Bea2duuhBXrNuVz9ztWFbgX95mK9Jao9kJJ06l0pXTvdd6DVJYvih/EslbT8uUaqE+ILc6Lr4j
ISEbnCDzpAis22J7hNGbB29/DoB7BBVev8DNPOEIdUuiv0vzfa8bGf6Im2yPhXoellTNUzNqD7ps
vLexdVNU9QakwOklmmMIBv7AitesnvzJboSbbsd3GVlEFzrvJ8WwhIOgR0zytGRUNBHqMb2TlaG6
iuVC62MK+mGdzIod2DA0ym7gRjxVtWq1nLlOKR1WoeBOKxi1aTQqyKFNAqa93KpQ+Svatlw+i08X
zMpSLglNegYSk4IYr9NekRgwwa2wp30toQPPGZdoDkyXYTbvG7zfklUlQro4uxy8R8PTjbYfv2GC
1y30DcGC8olxKa1+SCTOBQyf2172Zhmb/6anAXyvd0zxEGKbKYjfvMbbsN+5LKtcWEQZYnka2TqW
GLGG0ERB3eSLyrGhD215/R2RhvjgAiFrTzrMgAyXPvcFgKohXsK/iCeMWYx9oF8gdB2Nf47euLsh
19lY7GMyIBqEAXRkpe9TeMYPhhwUy0AKuka8a2pL0nYmUV+4VIxoKEkbXrOvECkE0xKpccIyUn2A
lVjMnJgtr0PJgC1st2eQmuxqQz4MvR01SZM8qf3Q62AINuXKTvj7r6smXkCaPUmxUchM6Fst68qF
4AYDT8bKbZgVKmnCVmb8YbmbYVeFD8Y0MKQToimHlm1OBzNh7iuYE2wr6yOKNEalGqbrXcnGaUfe
w8ChPXJZpRrN1ulm6XQPyFPET/qSd9/X1ofFPAi8+YpdttuD+Q8WMaze0ID0njSwXvilpPe4TNwD
OaUp9RKlhA0rzUUoFTNHiwi2X75+yP3hwmuYRuXoS10z1pxb1sImU+jVTH0LR+L3vqs8XuAdj6jh
+LmPMdiQaWFhO9u///n/OVPB6ZZWz8oN60P4BUMDJ40aFAnTFs1djkCEM8r2vsfcdbrOLlk2wp6x
3kIcCvlWShYCmm6dIeQCoCBO2k/Kqq2QhHdN+57oIQE9ObcaQTbKPAp8CX7RBJlqrf8TlWTY3bSH
D1zq9OJl3mdc6PLMX68NJUn6NqICPH1+dx/kXFneV2rUTydgBKOdpf7CeOGQAw0tVLAbhdU+7j+Q
qDr5Rik698Ky9RHAwPHuqhPzHckTJB1McDc2fVoF5zEIoXFxNw3ABvOGCP7Ks97AjO4MwTTfwr15
qC2AfnB/GMONqQ5b6yh9FcKsckOVY/sCTysPIklFJxuHU0rVmXElAiEBEztGFMpkMjt3HJGDllYW
fVCqP69Iyd8SKRbP2wzglQGnbhDQPTlDX1XYlfRdUvK7dGmrweN8KFj/zPuNp5dE5zPcTzVlJTMA
PblhfKcL21JU10ner8ElVuD553JrNHbcVh+xy8LrS8WDTCm7JgmY+Oiiwj937GpHIFBMnsADeHgI
waW6LlimkjWgA05qxjim9VAVC+bmNpOYSJWgkYXacH6nPcWOVvn+s3s/p7VyMfKaFLt7EHg8c27B
lb7grhD7Wxw9GoH56UxYrhQNVo3neAQPk9db5MKrO6KKXQDWUlmW39Pg2RXl88e+Y3in/V1G3xz+
8kQ51CKGaBftPgDGi0f/282bSxGOp1OyYhBx3mWkBDvSTrZCB2S2yjlqtxG5VVmVO9BOjZR8HVLw
jY98EW0NRhamrm8ItevLgWtR66Dk3qDjVvqkrmw5cEYXWO7tId00JPMWwjhWPQDV5Ec/60IffkLw
zUN1ZBwzLRt8SVzsDvBs2zY+4fxf+F6PxoCL5mwSxWSnCCWDQdy0/itId52MJKNKUYnyKgRnXuxU
yjtqw/muxwwYhTVQYZ9c+NJnFVDrJptV8JLut/AqPu4gqa5zHJPSccA6G8Mau1d5R6L6s1GAv7wu
f8NikWFuScN1RWc5wIiqozzP4aBnSlPjAYRnP93J+a37CHQMHT9V1WXVQ/3jkqzrMQ2VMOVIRiOy
0EmWg187gcSV+q5vRx5PWfZzEbzLiND3umbZVhUwxQIyY8B5BsZBeL9rpOdojUMF6FbH5Jz4uDPJ
anLoLpSu8cFFHn7XbZkTOCjOqQy0GL5xMScr6aSAg6zPS30uSn9DTKSu1AbZiM8vCCGcyDlJVaxs
skmpjuQKzIEe4+k4jsXIPpMmnDXzizG9yhlDPejt0a61m2T/3vYqdJZuFYdm3BknffzbzACTHIAJ
Qh/iPmYUqyv/AEEHZR0g+4xLH75bF6Djz5ED7BMjVY/04Hp6z1iS97D4vUEawKToznxaxDgiC02l
ZCRoY+ZVI5uiox9w3nlEnDtfTDsoXwrz//okDnFmLU2ctKDgzqkqT6aizJYsfSObdWb5HpIsP1Px
5LvLl2lfJmiCi/V3TgxfY2cbGqS1NDM4Zsx0mRbm9sifX1nLJEBp/0z7y/eX0qXfZaLOsSxaXii8
yGrX890GCiNKpFW6zYnwqVPXflY8jEX03SwAj4yxDnCgCozYqbPuolsukbpwEe2J+V5haY9unCor
SUJ1L7y4aOpHyOAAca9I8gg9f8F4EWFT24HirAOcX52yrWDKHIoMD/ZGMPoblOAfHsfpSH9U2j5z
b5/AqYIjDREB6I610ZxqBYlXUL0CgCq5R7jTw+hAMJWjPrhqZmF0VvsrYTu2W56XxsxZijusnue8
tqtMBfWOynySP+tLBayUshoupiIArya4K928pU1GBc4YaqyqTRn9++3kJ+ZR6lxegf/7qrdehxvs
G2GZcCkSEgasLEm/NKwzu3+pZ/X83P6mNfY1SNS77rUc+Ih8LbDHkbspHyamV4zdGt/yLZ4tJGhI
7Czw4hEo3oxKjxbM/rWNV8z5K6ifYCONyKoJHfqDnfvUJ37Z0PeNYuEfYF68hwKF2NN1X40LI8VT
mv3SJcCt+0g/t0HkPsAy+crO0x6x7KUO+H3mDfdQ6pxdzMXPMf+Ctqh1v4NLURpaz2dsCg6390Cp
VuBsTMSo6qfKq7lDO2U6N/eLaGuk7j+0A2SD2baGcL+j+B5k1id9IUabTWNRMMnRaxYdAHil3n2c
R4dGJqiVoS2ZmGpOK3DtkSVI42GjKrSjv83VS6NG2+AN7+PpORDDIxI5/UHsvV/3z86IrvpCfDih
k+qZMpaevakuhxD8PO3qdh7jAdxjK83VQs9lW0/MEwuwo+/iJyVZ55TU3yc7fwY3BJC4d8mUllCo
912cJN5cHE3YXIEgN3SFj83RZyW4BzNEwaw+Efw65yfA4Rh4DfmRTncDj7JqzBrYi5iu3DJRAO0E
dSscH71fmHJuO4Ol0PGh3Vh6nfb4kbPUqk3tyWxGHV3ZxVxreey3HAoAIt1NKwvLBV2+SEwCbLmd
cj5t5/bJ7AJhktpsNv1Pkd6FuB2mnn8A/QJSYeNJWtrKOP1xNy/psoWkixV1O7edGStLAs31zTCO
+RdwBDGGDZyxnU7HjGe/pFARN2fTJG0fGOoXJc+FFBDF6VyaGRoq3+OK+zsBRzbEzBKREs2RfXRh
m+SoHh2sDGW1MpyT6y0QUCBjxYzN6m21K25T42ZcSwrl2gqRYtdeSljke37k5I7Q7uTxGAZC+8WO
GgXQX6h3+U4tQj6nOM4m8L7v+coRpA0dXYfYPBqrqeXnduOHRhqQ7Cmd4slvvHme2LmjamJxk2mE
5699MYSlZeCbNwNT7fKsVR0/RnT6nD47IJPUJIEfD1HlH6yWer4+pXbszl/25N1RdCKskwEmJ2Cw
iWV4/48wzRMmqIVoFRXiKcHH9wXw+KXE2Je3nrxdVFyDalERjbNHNkk3+R+Cw43Nfh/CAm3P1KQV
IXF6q+SHuxdjR3mBZZejb5SFEKLUyc8tZogdJeSfGkeoZsVMo8mP0e7q7Nu5dCemyMWtbDwUDj9a
xjbn1aVg4BhjA7IMdUjSaiY0lrP6W4eEukh3iQhzYirGN6U9doNkgybqhuWEsLo9XVR9K6vpxKM/
J9GJcUFPw9iJj4IcwxqZgLLMW7/swtBwqy40MphWfVWDkvGgM/+4UGJi12lYAb+/vitBYOhPgo2d
04KCo7D55J2k/nuYhEpti/Roig7nnkgoPG/7S3Ejzxp09cOQEqz231xtQOH8Af8DWP2wyt6ygAVC
ktTZVCGrWDiHfyeMtH1EPGebaPC8ubn04r26bA984si8Wjl2JG9wYfIeJ49CC91DZjk5wZ+Nt/0A
akStwzJbwyWEpTNLwQDVUyWFbzbjojn9ksDasG1tjlCjMa171I4zXw2GMuyz4cki333AwA9O9rGp
f/8lGQkPp6ZC5m2UhbLDf7RpJyMu0KDLYEspAgVGpmSgt3WgRGbckx4zAzcx5waokUAaj3+5ZZas
gu3C5q8/ct94rMovw8QBBjmSb+aQqDwgDpACC60AVRtrMg8FTCJ3u3rVekNGAZkK2EDP9DUIxzg5
MfQRSpoBgh5tYgYumX5DqNPwQ3KRt1oLV/tszEO+qEEkncvgzfBuhYnbNaJwyT0zhaODqTKzo4Hm
K2aTkemjZS+Qs4B/LRa1j+BZqZAg5abCStQmTrz9hhcgYOY809+90QPaRYKWDTaR653Gx3VHCf+1
PX7lQ8/tD9ykrpf/Th+BLno/fNCWpMc3tApF6lclsAeARGq0LIeaiL/uIjuoHtv0BH0pzPc7unQ2
RjXqctiRlnh5slRp27sLFpXytOy8Qe3FyzjM8g5R171o58Fk4EENfAx2pbvdDG+aKao8ogbzc2Ax
UG5xEsUtNbOIXyaDECr2qpI0Y3eGVeDEyFHKo6Fr4e56cPDTL3ow+jyUfJiEebYK/PQ5j0tx8haH
SqmEDkDtMr2lveKzDSFQ/B2iwZrLC37i3qvcuMQTbJ/yjNmVK/W7ZQTJ9MKZToJS958QxjSB7Yf1
dSjLmBb7ksrG82HxyRVDAx8ecd4Dz4NT4i+5DcdyrM/lbL7l73axiL5uAMRXlXp39EubIKhSuKSt
yGS9zVVwPVHPa3FzvWn8AmwuDtp2CzuTxzT7aGZWjds1d2vFF09xriTeRIuM8YE+nQp6SREA+2vI
dFigFIkPxAoUk9IbPrIayBQ/PfrqXCiNR6dPAVJnxUhoGTumngcwby34Ic2bV5HdgxHXQVf7Y7/x
lwrFc1KczYvt2lHEvJd5SBCr5OYjhPWleXaViX27Kxqut9c9KfxbjO2Mg7qEsh7LAkCvkPItgeeH
bEFSmnyxTJJ30saEfnh6P9dedS5eUQYE97wSU1nSuT2XXDFTZQ4CnrckiCoi56t8+sude07M02cm
NpXjPhrfuuN7hoQ/IwQ1ppImTJ5c83ilHcPOMcJUVCmdcG3UoAEJN3M8UTl0eRbTIqqPfsrsyMMV
HoSp/S7ihc9F7P1nr+YhR2p6NWh8L6SEJNsM0sKha0qI+zQFFfS7HbtnkYlJ4Msn52RrKnondnHI
QrwAGqqD9Fw6sILPlAWXT8kKoBfo5PNwTOpevnHgW8eoq3G2gFb66E7ig8LXpRT7CoRQJBzGChvY
khBJin4E+M0WvGjVo7egpwifvCOo1VZayirbyCQBOIkYbaFNfIDFEt83nfPGwPCLdKkfdpyXmspT
Hd3egl6Sj4WAif26OcR1jb0+1gvFpJmXuiD6oCqvmx3ftY6SyFTT+K2LP46IK0e+jmcUpfcufGwX
jr5BJrR0qfXwGGcdzzVgtP8aHrBDHrghU9ZpMcJ6vVkqJIAXiKeM4cLD1B9wG+3EaLRCcb1P31pf
Dqnk0DTy6pEdHU1b09TIbfjNPnzEtdDclUFAyH7hUEKutaq8kL7RXDQ96DaNbTPFpcIF2NSs1cbS
LzLc98JOTWqhiNjNp23ZAZWXfNsGfAQ/zZspIoVFNtXB23ICyg5T/TTOc0bE/y7iBDE9utIgUV5+
JCJ62bMUc2EjxBoIEv408o2HLIbof1lAeMuKk1/owU66jOSIz81zPoSpgGP06wykAnmUzw5lJFwn
qW2FsDtTdRLfVg4fmksUEFHsYQlBEbCsM5s5bKjswPKXFnxWMwI/7s0jEEwpWXAd79MAL18bBAWi
yNLLdBMe/1UhznTfYF+v7Ta4gCvRTPUJVHin9+uy5GrtePKxfRPM+8M5c85aYNX1DsOftSBtwgWF
Pw+tboD2DjEJcpKJ3xEic6HjP8mjIVTD4H4MN8/MfB2/QIUp5eJCP5ZnaykkpYq5WT2ewVLs8LF+
iBPSTDuuclZRIfw0Wi9I1bEfLnjHETj+/bHq3t8mxvg4iMuqztHLQ2l3JE64CtJog2k6WRag5+Hy
QqZEaV5CuIrJHcN6jg92+eXYOaCFj5QKSkzQvSSI+TFLl67fnkrBQs2ocw9Jzj0gmEg7qOMDmcaj
NmXqJE8+VTgdG+pQ6clryDK6TaivDTERVEXOBJ8U8+fIoF2/qf1XPCaFq1rbJ/ISqX/7+LdEYlLh
cum6uAOMErJiYPqKz2h7H7oWSXbutKaqCs8OmTZtJ/BcpYUjdQjPKrrSYT79ay4jnr6rJ0M36aRR
ZScPFylayeFuv3kI+Q+OXybRA9C/gn3KlzuPXyzs4b8tZTADmbPwFCRCACmGL70NzMezYsfYgyx2
S333LEXWaHYmmclbeNgyVTkKZUKmK8YAMAVJQLbe3u4Ll+manHWGNV8SNws8MfV1zVnmxg6G+OHA
A7XxC5OpYETkCDFW8ehRjmMEyqc1BRInhJx3vflXmXuDadcoZsp4HdcU71FTOHQik45XWBmh6LoU
4nrPAC4cvBlEfAqdzKUV+0VmEavjTAN5sU4QK62vCUvJlrBo6A2bcRYvcA/enIIeJoqi7ldYI3OH
jMOf2n2OQ8j/1zOssRRhv7ru2GlB/wQ13kyILfZ0MbatllKz2B3MMWpeRPtpInY54/YchjdbuTkl
bt8IMOVKpGfWuTmNrvcO+JXi28QpKAMLNg1b+/L1EDd2090NrDOyXbAI2FJfExG+59GmiCMhuLrd
uE6DQfR5QL74NigsaYCWF8+dFNyYXzhfe4BV6GkjFbAdvjzjh72VQJI8JfSdz+jjhdOs/Mq447dl
91puHiGTYyslGG2cNoznZ1yNUtLaw02G6vjiN9s9sH0lNtJNb+2CkhAiSek4PyRsewF/hyO4zIAN
bqLxDY2ZQ8hADgSqh9GWsrpPTS0AS+54ET4RIX9RkNEYcN3APml3mUl/7KRFeQ41uC5ur8p2Gc40
SefzRi0a+0e+X3uBio2fXxB05XAYhM9O76r7Fp1fv9BsBI3VQgk4Y2VA4XTNdHw1Y3Sx/dsTCdQ/
VeWQdL1CBU8xSVEqCDWKT0D9To1LyzPM/OChp3ud3SlQvIjh6TGrtG4xHPs7qw6tBElVIRHKqV/G
t24hw4MJBPDtgD/La1kYqQmPcYgWT0oriWsmC1UWNcHUbECN2RMR8KbBdU/JmSfeTQo+7A2jMLkk
E0m9c0A4amUurbaZ9qM8iaCYjpwdDMHV+4a0HoRwo4Ipg8oUoNVaxA5EZ/fQNYakla6dqH4a1wo9
xAox4dticypPJRiCHxyqW/GDlvE8KZyNWWAEvpjSTt4JCH9K6fodB94zQ0kEfmkfggSNdMHYNFYF
Klt8NPBrUslix0lWV6S0gBHasgBKzSQueNX7j9U3HmELw99am8MHM814yIdX2uIZUJLvRcP69Upr
fow+5agYyYDaRR7ZXYqkaNcJVEuBXrIJpLswSm2tKhftTgbZVhB+K/Bd8WKn1hen5HZATAut0p8m
sS6fWkks5xKMDKoWcotxe/bCCEDigm3mzVbhjGF6qXq9FBas+HYRszZU5bSncGqyzWRP/bFmmq7c
quPr8bTLq/W01VvCFfIOn1A2aXmlMl3D17BbjCCOfM2k4D2/KLNelVFy0kCHSs2lpabg2qLjFFaw
f2/UB3Lta8Pd93VTHQdGRPaAsf2F2L8x7mxPcUAqTdYS4wjzEE0OJlcW0D6YlPBsIVM8qLgPRotR
Ym+pKthlfgFaH0GiJl5meLaznxKx+tngTHpA/cPAhkyQBfSBx/p95KDJ6f9MPZ9GzKY4CU2H2vJg
T1E4VGEx7x+Oqs0mWJPlg+py21pjWK8ygyYIgDVqpO0EnDjt+9dz6874Zt2iTSPlKTyx8/YqXwki
99taGm7hAJa+SYqbtuQf9GFN0EKEJrCBZA7jMT/pyhLHIK+0hplT7t+u90nP9J7Dlqdy7l29tQ94
pAWuuKqoYi/WCabaKChzVmfSEACUp2r4SXzhEsewdnsjxvC5b2uOn165JI+rPn0FKo2iJ/ohTFmW
QDoxaBYck52ZPrsvjIKWFi6WuLEvO/ny7uuLkxiU98bFBWKPLH5F4zvBcJmz5XvXuIyMP+Olobgn
TtoM8YLmWybIZ5sVKD9Lhw1x6PZVEhpHxy7ndxPts8Ei0vQDczGiBXPHLX66Tq5M60FAur9PIcN1
xhBzHvMQKWVzB69qIvGjxxDnkh8wNGay9x0uCfREwcbqgapMvBdphPeGQrw1C2/CLPze3v3EMv08
B0fvJS5Iefq2HxlEw54OP9d+h4qW/BidCEJ03Z1lpaVMmCFPbo2Kno5RdRG3+z3lID00pUMfwdhJ
Rz9RoT8drEm3VPlEJiWd+ej/Yu9Ad9/MfGx5R3488SxBZ1S1RUdpRU6LACPqPH3/9tOYJLEBK5b/
kLKM9AyyqJ8qgsAjWk2nwCeQpd7sLfdlIZwQ3prxX4DhQfnqdX9+Afw0I4rcQqUTasWIaQ36JI3N
H8CQgOY6BlUZp9EfWLj/oh/Mtg0TbAsMZbhRgCcspMxROtpoXTAX2iXirArPbQB6CHg9OKxBIRO4
QTft+miPAnO09z38ROcAg83viut3B3pUuXI+7/qSeqUlYr/7a9Vu0+vKsJfLxnictwAvkDAn1HbZ
CjxZqqzussquNmCcy3TD2SQPxvJ+MehVcNtt+3/ystuIBIwTR8ndN1GshLTkKRBC5kxC6xpZAqUi
qE+Ub4eUmdxocF2TA2iICdX0ivgXK2QZm3Tnt7SrKNH/PrP2KtWo40hWNabNuL8779GamWAoOicU
D1KEE7ciCDFcOq2i4xUVEB+fvma0o0ANhN186u7W+qhaCtwxFnBYiciP+QcG5VVrZZGzM7iZhi97
NKdxgLs5J79lgNhcw5EjCLlg09oKuPfVMyd+tZzC8+S+I4beTOswV71iRDDN1EK2JmsvcQWx60Xj
uPyPFIYk+nN64lhrP2i2zjc9xCQ44ppvlEdilnchXcdl1L2CgdRIXmdlE71EYj1u9UJ+7PHKY7Kd
qwcxmy8Twmj5kU5HBd/ZSrHRMNL1qG4xje9hjxRZA8GwkJjeo4S6pP0z/z1hKctsZ1v4kprOnWKs
fCmXH77jpHfIxziTcGH746093sufbOVwCMnELdmGAj7pORXqMXLGU2Tc9FKJGHFqoKSd2oEGlq0X
c7DTzS8rBKc73wdQ/bRcrtMPJ9TyvMBp+NzGpg1pfYVObdc0C1g0FqgjvH7R6KEBW/kJy6w+Y0a9
C7KH1T+TK+cjyRFxKD1gcChZp/iRWwuPmHT/D+fKin5o4NjZVwsc9pevfNiq+CUAG/rdJp3rT/j+
BUyZojFrTtxe/Ccr0j9aS7+SSY45MRhcxyA0nIy8zyuaf7sVHMytPYaHTNq9Hytv08iAV14NBXPR
5k3fu3+9X06b9iWIG4u/8NnxzHxZW01J4Tl0XNi6UyFBOMd7uqtZb94d6euxpUhv4RRHorQOODHN
Y2bxhuyVmW5htwd87GhTFKf2WUsq4znpuDVm8YTfCtFmHpbFxYK8oL+6OrM1MSlF6mtz2DWtXuBA
lg0qRDP5RSUn1dPx+eplMWAKXA9E5SSaPw3TvyhdnN11FlbYxhFhpKVHlVBTH3G9j0VwvnelhocY
qxLaD37TWYS97JoE4Qy3jHxgh5h8/RaPfu/APmaHczENpgqBOIHbPjtgOtO9lm2otbieSvBk7rgQ
htEvSZl69HRFMKErtBFb9nCmcX+mGHkUW8iPfciN4EgnxPqbII4pJYez2ZAmOLSGmpOw5L0LsUZU
ZGWuYI3C0Vu6tpG+enkRjaU5MtB9RwBH0tqa8IGpNExkunyyC3Jt+2gHTphCv4VNcbpTJeE7yvk7
JKcK4mjaMLiBLAE5CkWDXqVZO4T3bqH9Q755MUEFZCprEuyr2+WjFG2vpDEv2IsfyFeHk9gv20+3
UStGyH/2h6REXME29Vo5qEmG7NE09l1S5B+sYM3lR9i5bK+8RU29LCMJv3ohhROQB6YHdlFzkAcV
lOZTR6xXHsRGqC405IHhq0nVlBnJ2xwlA9wwSUsRmGX0893k3/k8AjDhNfU5SX+wDRgArG6lnzrn
6LhQJiBkszYBaqbmzepKygXqN5fI5u+aK9rtm9i5AajaaElYhCYl+HX71mG3UAkaOP7JmEOY9nys
SOd0lYYleqUpl4qzbJXYZcDwkzu3QwW5LECzl4Ke+vA3kixgljzPLQldtLsu4TymaZubRJ/PiAko
MpJtdaqjBySQBMB7cdb/9nXDy4cv6/TvvprLHphtmsfaOF34JbWPpdHREiBzE2peTsMNH4AQ7oJe
BZTimn8UDxd+ob0wPnoy3b73CFADjGbDK6/qjPWf+GaxtMOKRSfnJf2a8/3WpHYnuBS09BBYCZ8f
5uzffFImKixaknFGGNEek9XO1bmCkFnVqLJF6Ergh+d/rd1QsNTL5tM95u9NJYuCV6GemM7CfF9w
DgsXC5XvmqPdN3Q7sq94IpAQpNSkuRmL12Zqls6XiD4H7mdPvkYlaacRlRye01l+xatSqjjVBJgr
rTF/tkAbueV0jZFmgtyzreKygPDVt6+CUSQnkZ7fHoHVNpAHaPMq5n0cVyV0AdhyO2KeGah3Lc7v
503W7ZQOqQtvEOU81KkeoeA+h3kuhOkSLSzdG1TD4Mi9XtrnO/nnTU31XZS8WZumQ2wFrYyHSz/9
wUMmjcYPEGaxZiEIR4qYvvxNGifBB/WxWUJ0murqXzuNgnb3vg9G8jfIllMm7BF/J4sNhuIeen3C
PFsRlXm431hSLAv9kTfL4s3OG8tfu4jwJdfoJaqUxNecK9wKvuJPCEyl+99OP7MUHG5hkwAVNcZm
bXyhs96/lkBQZ/rREcD3EIF3WKuUQOvvU+cRPZ7paKezbLt0oG9FVar1yqCHrPo3M6iZbKOPx9zH
H+0bui2N2amiw2OPw4lSnldUdr5UDZ3A4RfUIwM6p/szfiXhH7ZDLpVRyvgaRAXHv7LJ5g5Iemfy
jARYi3bHxzE1A+ukXES8zrjjSofopNORTwj+RzeA8WnbYQhYYVc5Ex1y/ED/vPszrlgdkfTTeGR2
Oe3ek8C0OuUImjpD4QThkNUt8a84R/2zTur4iaxxqv2QwiSINrbQxIBZljBCgnMFQIQIEZMeDthh
P+Q6uq0w4pn79h8SMe/+ShggiJNkQHIpmHD3ClJHw3YR3QnX8DxZqep8d3e926Ip/rwd+ynOUyOi
TKl4ktJEfX+V+HZOOxrgOiSER1eKLjXCSYNldAGsSOW39A02o4uvHbMb4Yjdbg1mqIQ67mVpQv83
d6QHSV8b6839TElx/iAqwGhfvhFA71FjJUtfEYGE49Rv9OL6/xHM3dw00B1TYeTpQCzVB83Lvqco
3+EEGZwRYzH3pm0t3Z+Ph/pJX/z9jXp7o8oSqnWHLbsBGXV5rATCyUJpSQsqI5gLO/VLslyHGfOF
8kVSX+Ef07oXF5aTwS++6gNBWCU6FDRSPOQG3PfTqpTkzFMjR506eca+zFRlmZ7ANQHK8mmkwgLV
bAYyK1FIgpVlvv5m1zlbUHuDWrqOnOjWdQr7T2UrDrp5WcT9yRCqU7RTGW4njI0GZ6Dwp4/ZWPJv
BWDpRfdsdK3q0mCh9KxZHo1uYtAhQbLvc1g4f2mOkAuGGT2Kq++Do2vb363IPLJpGa5nW71i7k08
P/QdBbAgeAjouUDw7eMSHov2DRkVmh/moXSa3U8KVW23vuXZXVDUFaO5oJVR7383ekb00ehkZEth
VLdQLfZDD0eQTnLE6OhK0OH7CogU/zHEq/ACb2JdE8Kv8fhPOml3YsfkhUnm9axMPmpxMMd5fygT
OFeU41ueryvM9K4BmX3oEXv3UbFqwudGJRuuPt6KThytpbZydGMRWHAIwFZ8Nn2sYbyqxqjgIUy3
JgFkiOOQHcyCh/TIwNmk0bWdsWaz+XNrqRRZvdzifUPxLc0IxA0wvkmXYRSmuFLW8SiI7LovsLrv
YFd2spnBDa982ZDBdVcl4GYdebn+yRUWghLQNG0QpyX0VgbPcSjsO+fYyfb3oUQ3xALAbXygdgkh
mYGXhZ/EXLGlf5wMk8OG8VxR2oHHVqeS1lFnGcduXjDiY0VjlYYdvmCAOX61fG+rgMvTNHxtK1DM
n9uz6PbB69f0WkLCF249Ag9VYxkwyh60eqLUZLUc4J6mgtSJNJ0w+zZ11qeACqvnMnEm4DkTPwIZ
CjiWM025SQWbw+RBpQIe3geo8GBFdhf9icxBnPiS3R5fi4BBt1vEP0u/HJPftj20FXY0mo8Zv3td
VP+fZgsa+dB8ER+/plGK05OkzsRlfmFmgRvzBHJVfJjPKDxyLvm7nZ54UbQpKDIpncYj7W1NBBD0
s0Hj29d5qMJdBxPHJ+VJ+0ZZGbdg5SB1sIL/CT1DUhNsz3sMTNfhP/qF1AmYPy5z6RNG7ziDt7ZJ
HAh4zneDIac2ABQv4CdkrAdqXqMKFTsrq8VcdxmVb0a9cBGQDIJieIuLW18abNKqhzyRXwPo0pPX
jdgiAXrGG7b0bEpAnWZz/bVsoixncTGf2Yl6PJEtqTVRG7Qtzw2zg9xbZDZV+HSVzzCbWfcnMyJ+
cX4N8IkV8W79UqaIUo7JXmPiCXAFLCsdUd56OaxxtzcHSV6aqGtMUe8Ije1xNJj0wWnngwU0Uq/3
zcnUs9uBAXFr0Rjtx9sXIJGxCKPctjSwnPiTp8wsO9Us+pbhH8RbOq+wcvfQZRWFevsx6heNY/QW
rJuaVA9tKMQFV3lDnvLH7f66AVJy/BMhcPyqazq32YCnh41FSMoYgNO0/u14+yA+QnRFSqLprJD4
gJsUauciiOVbkM3OkP26zZxAxG6TOfVxrLyaLGfX+Tsp5/Du1K+BAjmpsLIm7Iv0yJGm9sWg7IBs
KwuAuk0N45X77P6fQ+1/AJXvZDnQnp33BSIxu31DJh26HwwtE3Nu5JC5MGfHzVgiE7OIjhES+p4J
0vvm4maXJzZ2PTOPLSC1ZUjsY3OvfcmCauUhnZ4lAbXWYWITNYZperhy23sEFKM+upM9lBRjNQEZ
TNge6X6qStiTn5oHbCMzpGiEnYXxugqSj5bgaeLdo3ksLbBU0f42XyLoXgIX/mFzAWGsd4Zhxnal
WXEZV7cO6kj8TLMoJLtW/ZSsiyJA6NV49qT8nmL410fO7jt4AfhmLfkcE1A3rFmF5z5KAxydSCWE
gs+8U+6EjEZDIv3lgyNqAVcvmco0ADnRD7sSSGgJgvSosDIfHVsdFcINQXOsrpO0bnhtnGLveMhL
1NMHfnrrAVDdbp0Ckby6+y9hPV9YefPRP+FD2jZqWHsoZE2okUu/FS5onWRWmoGLoSQ7Bmh5XauJ
xhhCjKYn/6WtH1guA8FCcNBYsYMPcK6BRz8cmm5P5cFB/RM/2v4kOYK3orAgymRJp2d6J5wS4zFE
qnkxeuo5MNGNywoSWCxBowwuNtJoMzSkAV0c1VyE+S1gc/WQ6fDYva4r4groVbjSS2l6gTF86xgU
OvTsclo15M+TU/rPWZ+5+joqClarQAYDs16Im5Rypy/m44xTa5CQwpBCL30zy9h9TBqZiUJ5ilkR
g4vnRCgfDzFhNq+qeq1eC5M5ZvG9KRyaf+0lbGZjmi31cmFS/8OOHlICBMVIHmNqxybcRxGuUrxJ
a7KfbamntYp/KaQYC6qioLo6oUdh5JpiaF3zxaxAWwN1xYeJBbhvVODlNkp5iZsU/MKw8zL2eOAq
tGBDNxv593h1TYBTo4oYh49KMrCvV+6ItmQYMCEf7Lq0jjJN/5ZOeFCYe2OB1oP5K56wL99wACMq
cKvBp04gVV8nm8yAdX2TI6c5TPTH5yjXK/MwC+VU/m9SOrK7oRayHBukBVh5UNA2cqKNFhsz5Im8
LgcGZvC9WnGN0S9hKEErMtzuIBl6LstJGvAKmI+3kMTcOrG1/I6Kswj+YSOqLJzcjteh/N9UmHhq
mLh3gMhwSYoMkr5VAQwHBKI0cZFeNyoDK/NxcEjalnby76PM9mJB6pHts5CZdV39Hi5wHlF7YS3m
mFyy8PJ6xkirVImTYP5ZK9misFKVdKI1iGnb46nCj3k/Su9PF6AVgIYBG/8D8hEed/Fe2L943Xon
EQvKZsbtI3aw7xgdS7gbqKuAiG+V5p9ydOgV2eHgntgzoB+jI7ctm3yBcY8v+rPccAYxQD30rdkF
1uc+yzH3LfMcrK49o6uOR45ylkoLNGOGEmmFHvanncdyGdeEzopNDV8hxtUvbYkmUN8l6XppX5Ls
5YoMj0bMd6NJ3je9MFpYMg8UpfAzyr0lv937p/32iIQzfaAw4YaAOo1RboajsutAg1DcKz4Ngpkj
RGxp1CxLzIQbH+mFB9piPAhIjMB37Lax9amHawz9InVYpVI6CiiaDpX/3ag7d4iJOcXU2Gtro8aE
qIckHAUlOGXsqw3bOsAH+wS88RyvnduZScRmZjPOSp4Xjs7StZKcVMWWc5QpiFy/bIOsFqtjIIdl
b/aI6QCArM6QLD5SOVKjn0k9akWtKoecK7u5yB64M1eojdJafqxPNQSLU9p/bdBXhjAIlqZLcF18
ovT+fN2g5QngyCntAkGM7DABUAX89A5Avtq2oAj83b+9dz1PZb/4k45Knm0wcOdC1pdQWYTvUmPA
ngBy7OJYCNg+TL1xp8I0t6kRssE5qzRPpYjU7yx+n4etKxVjS0Kmr0VGNrujSVn2Z1FDl7tLTyO4
ahy1FRoWVGJRtBALKI18o3pTXAWL5Q8UOSvSccyM6/KwIoXNWg3vtowgr6qCdLQ2zNpsrTICUxA7
XfX36r7u4zDpJ/yeLZTDbVRrE1Dvm4QYBkp94XbBsgLeihvW+Ed9TJBqa10VZdDKkq03KaurxwcB
bi1gmvI8uTDLPgI19CntOo975kT6zkQ7y53T0KXK8RAOTBO0TxdRAaRMxlZUlyT9V6HwNJ7roPH5
//wKWYT/7eLcVxr+JwR5fYXlwz2Wz9bH7HcmHwp2PVvNkhvvJEUaTaX/yLzsUp+yVvaXiRYNZXiF
W7ZbekG6Ijmgdk02esofLZeT9G3ODaC9D/MObahhwcKyCUZFxON5LfNNVHrzr3EeULAs9KeZiGw7
2H9HMRz4aXUXw8AGNKpXAKHP7nRNqElpGLej4WwjvRMkkgwxReqePpU8vTqp8LpNcJziqTmubFUr
x2+KT0ysJMbcpCm+2IXhF7JsRS+RwLlh8wN2Ag+xyIzayA2vY/dQxUlfGXPcqyb43x3Z+xpBRMLI
eVl9wSf3SnaRAJAnGhpCA7Q7XpZKzLIgwof85q57EJyq1eJe8hy9ozCz2YKIf8ALuoszhdm5EaW0
aNKFsG5574cngUjrloE6kQ8LOxS3aD4niYYqoKJT5hN5Ryb+MOepQd23CdAskznnM0N1/o0jCLk2
HYDYU9/mTp5T6W2IBMe0sMkSNdGfjL9WQCLMYO38HVs8QZ0EihZtayG9nEMXyjl+G209ksPVPGC5
Xl67kqV/R7BBE4cLy4F2yrKFtpwAPUBTABko00UDL+eDZ8cCSCQeIv8jUb7Uf/43cY82lHsx+AfA
dtsXZSA9OkgLPckyDchnQO3S7BIhW77pAqzmUAEjqQoFzTqTuHQWTNn8d6eplZTODNr/X4QBv1Hr
2LLtiPkHsa9KOtwENsKeDmHlVwKULzOmBCF4Z2qLy3jTkFPtpoCdf1z1y3VWWhZaDIFgpvEci8lN
mVYUx+eN5zeWMjfcVe5DbEXkG9+M0YrAkLwJMa4Uefxq5p0keBxxTiU1fEfeu+KEJntxB1ac0VTT
XhXEkYDCkKojkXsEsRw15OR7jxjsY5aTuO03k5TgJimMilH8rKve5rciE6UlQDESJsNrvGu/aR9I
/neLRO1aoTlJkHaLRNjcpwm46UHBkiJyvPxzDq3GpaECzxGkHbUHHkPBnw+oI7v6jrBIlUOdApaN
EzhAw9lhIDceP//ViFP+eEtm/HGgm32zISb61a5+k6UPAklECP1YtkJF1jyd9srm/8dFt4kno4ur
KK2ZCHOJqe/2LvOrDlxzaOh9q9xYlvgg4SEK8VTohOi2qnzAuqScPboIkdJD8NS1H1jc8J5Z6Y4R
+mnBovRX5UKqswt9pkdG0BwunHe2CtYfmj1xM8O7TCxIDJGcXqtZixszBz4z4VJf/7iCUi3SghaI
BOs0TzvAAJ5l3EgCreUZWhG7lsd+E2AXlpS+mzdjlN8utJkHhHgLmNUkbcED/2VLf8CJ7sd4GYv7
NNsKjLQ7yUJBSEWjmJfFveo35zIZLif2zo5OG2mg8fnpRdEAsZ1/ZTzZBqVcKwd2IN0uht+oHYwz
oIgsSQas0qQiUsR48+xVApdzEk/gpqtcA1M2XgKGGk2Kwy7UJe6izwcg9URxi6aUnS/dWq703Wzt
d9nJGL/s+FNTXij9pDpNOazn6dkBo9ZpN7hDh4VCEonaxcJ1xi+pJC3FacvGHA3dEUzChemmku/A
sfEgnwmNHmkqZ+2OyFegblCLtnBJOMoS4yiqSGnmvXW1E6nJ/uNHXiEthhF8UgT8QcbR90j7VO/z
w0h42PPUIXr4ZlK6I0bkQXB+Id9m5aZ6mF2rR6mWZQi5UuziRzsMYdkzSCQwSAtb95w7PEBm16OB
RwqgBwfyYw++O+r1HuJBH0uK50E/cMielh4iGU3GELHBwF3TFAJTdyl3ccRymsdaiRWZ/VzQszAt
bNvY9YJwRuAuUNOEaT3CXyEambIlqeg8AScSTpIdAQfCCZc7vXTn4tMTQpdo3CScRTfdf3eSXtHD
xqdYIHXxBHAGj2D2lx1mk00POq39AKnj6jYWZNBQTTTCmi9mzrHUxD6I50I9kASXLG8INnNY/d0o
oG1CwkUyy8o5ddV2TYb+6Ua/LZzYE73eBl4Os33Y/3eW5wImP9zbey1W7SPl4s+0Y44xFoq3nUt6
9aK7tW5bOo7xol+HCluZl3siijUm1sbHgnW5DV1Psn79HcEPNsC4sJj4j7Xhw3pKSDj/ZyrYH1lk
AiRUvNlsB3M6iEW75Z8iuEa9b/RTeMueP+9Yzq7SixL2ILYALgtexqJCEnctjNjzBXfdjgg1nlKU
rWtoqzH4vrCbjfvwNGLfKYccHHHPJC4Us8JTjGXuHKDgYzfgUZ5HSJyaSLRdmII38LilM+/xSCLr
4G+Zp5XsJxfpMAPiPKAxTRg2i/SxMPwkQ1BYq8mwzY3XDhXFjXgndJ7HJsL8XLANPfpCAjJhahAj
MlBsFB5jtIJ8hZSYRbP+pcnLBoyIgEAOa0AuizgGkH/c5x7VWb/xKEeJuAJxGSjzmsIfh8/pWKBd
AooaGyJm2BRqDEkcoEtdVj8IAuboYuwjKhSgO2JNf1Q9gpqAZWe12J+glmxzakuzmE01uOVJoz8o
J2UDBKOzLFoIVstUCBRNkGQQRv0RR8wFOB5QOTPpGVF8NCxt09yXOm4CkH0AkdqdEQD9rMv0QGLD
KLiZX6Zcn9Ltf/T1N0qiWXAJzTTNvb8n9V7mNaUgpf42kGm5SUwOs54XX84yddofVwXs4I2wPOGU
YA8YnqzCRmF+U/rYE52meMf9ylkH19su2y8H7PTjw4W/1Uo88FMq15zmg9trl5BwDR7oiXfbvenP
bTl/rYAPsvJ6Q1IwM06IhabstSleDSDZ5nsSyA8TTKCk9s79DUqJnVD3s4gCDEhpPQoETURydTBw
U4pHb87AGJrDuwXQ57dN6rbPsyohKNdBZkEYpcDrLARckUlgZ9xpW/XPQ8krvQMLFF9QGQiS/vwV
nHS3XQR3BjlNAQ/7jCFtAqVYQngvRn6QFtuwKIm2Lk7MJ7wOhNoMIT+K+dOo3ajtQwzLvjHxEd4v
ayIasQGoVsrlnyeMDybWNxKloAhqRjZxHsQskWM9F48/Vz+gSe+6u5WVo/7pYTV7PZd2KwQy0Hpm
LhXX+9WIzpYK/IA2AHtcKtK4R/YcO8qgntlg2owjIJ0KqSjNNE9cs6WfjyheMZ/UFu7sAuIF8VD9
Xyt9H9gQcOc8+l7iiNAaI3YOqgIAzqcU/VOF+DOrPTqHh0QLkBHRouo3+glaWhbAunh8xDKz2mu6
O3OJQQqey9zrfo9wYthFHX5S4spzSK5J/wXshvPwO71toKmNylPFxcctBYJ6/8tJ+QV/DYTpXrDS
RCSr4dwF2v20pCvE5SwKIru72IJHSu7445wljPne2EAz1hP0zR7lw8zhkxwcaqE2t/EdnJmbEhcW
eACmknA7pS7tVGvlknhUWdmVITK1YYspM1TnEgReBEsSsPnP50RpV81C6gEYnOEFMBEs/ST8zuIq
eoaGYJh7um7c5VFAJcMwrpWq+Xwwulah+vxoNRf5zgvg+rjQQaeacWP8fn431U6nXdqY7wMQf9du
OsU6NhyciVlgMrcLZe6u7dUnG93cef8fL3JFCkQ23W5OdfYtLXzuP7P78sFItZ8oFUxssoNv0dVZ
KnyjedxXHbdDibMddRz4UKKOkC+axVt7f1S8aI613BJ7vf39J7vV/FJFO54bhrJgklhfKFffV+x6
SWp2aE6aPPAYix6k6BIeEBiWwFRjecVR0dy9zlfHjsMyUmcE+xxPa5fTnJwuLbefF4CBg3bUc4KG
fnNMkojkzko6H4SYTbLeiDukAx17dgqrasp7qZm4Y359m6FAtgh7h/XTjH7NdgprjkWqJbMeeTs4
0m0NntL3R8Rsh4H1jb0Nd1c/bz/r80iCyJMp7LiD3Kl+zjc2k4N6IZACaf0ts2FOnJ+85zgoe1o5
kKgnq4QsTMwZP1bDmcqJTE+o1MZ2SFGGGu8KKvE6UsUzyownSS6luuh1uP6CyNBUCFZNdUqkM+jg
1NPjMTG+vVU/QJDfkgEak74FQFAyGx3ZJITjvomHey4cVgyeLAGHUlvT54xgyMExPMMx24wt3lwZ
1UkHL1DCGnfFyOoWpNsuG2eEliZrZIN32OfpQCVkaa7SMMXa3tjuQ42HzMZVnzXDduE143iWx4BP
CWATOS9L2GQp8T1JjRB1+M7X/QuSGU/ruvI//3f46ob1DH0q2LjO8BMftaR47KMrAU58CyuJLtcm
j9WUXBj+qLswuja49tMJfZZCzL+VTXvgMdq+KwSyEEj3Jm74EKQvsNCVSiniLPCJavK+Uq5KsEqV
Sd1oCugca0sDNeVytmCBA5siW3Y9NQlWYUWLpRgwWh/2FwjjEdO8g/v0l1eSpmDhajaE7ZxdKLRr
I7y0uBron5c8I2mlNyy3Ar3HXpH9b/U3iHAtYCnyRpAGeG7rvOgpz37qvV4UQImOXce3YJRSvunz
uYBDrPf5vZHdhXlMWVPBfcdBeRn5dFaND7+xnQDWnFbLBi5284JQLAwCOO/Pc6kelYjCHDLg45FR
FswMy0wW1oVBvsZkcDhNzY11o2qsKRoSNNLtwVdgizvDHZcatkvKI7JmT9PUNmgUjIT9Un1CZ3Ml
lXIgtlsy/E/vzooJNq7mffuqUnFjXPcpy0VQ/PWC+7xIhunhJFQZ/PeApFp5pHGiTXWojSQsGHGg
u2kmUJSyHFJgdRq/Lhsl8F5BW1XNj2tbjXkKl16E5YJHZwFSD7Q2h8iZnQyu3rf4qo4yBNFCEESo
76IOKwCSFvt+CAYTmFoPotiMiUudZxv+2oveT/CeYokR2I+uQlbaN7Z/KujUwkG3ZbwQCLsSisZD
FQhzAh0qYWafR8RNS9DCq7Jwm5D+G9akfn+hBihpftugJShNTiNg2uiwo6FH0YSUoqpHqtKOSudY
Dx0zvhtcHaDNRtzU42RvjAcFeON4wFY2bfAYxhUrBFvR02GBoTO6NFmxmz/U53GMgx48Yr/3wrMR
ZZwOUJUimxFd5tt/HDPGRYqqeGA6RKgJhKIaHW5M4lvl+9ggYCa8lCNiSVGeZaEZCTL5dJfHFySH
NcR9UbFCYt+ze/ItZT2YikPe8YJtXVqFsKRbBxtk99RCeYeX8C1hEB3TRlbGWpqmVYxfqYIforoh
JeuGjIRPmQ9rQw5iw+8Xilw0CS6X5TQhtYg9em/CnReilUmO+J97SGyEdHEy2P82I1TceWZ6c+Ep
tUdhbYmpWuDRXJ4/bUIsFLV6KKXvK2kubyNl3mRiFs0AOAfIDVfZ5g0Vft44wVeDI63cctP7Yga9
WmqpuHDKULKk83pY6m8E/cFFWg/8JLfjMBtUXRpIXbksJ9FhAGiF94eUL3yTYDpC8MvIbAH7AQKf
YuXf10/mCtphILGGYE8jrbF8ql1Fmu5G/TnJ0LBozPNPupdhJNyflbFk0Nh+fYYm//P9Vb1GSNVm
kTZvT0QPJdXBg8uU3KHq1uZqYzkNQzm7nE3rOItvO71Wm4LKpJyU+Suo+iB6tgqid8iEfyoMTfGc
IP/jSn9sddAovxV4ZLu33hMRy0npk1319gLba8nabr1TtL1AqbeEc9ZiXprB/aDLcJ2DqvFQdYlD
kHtnIKAjugzByPLjEliOF4kFed8Sb24ygNCbS2urdmuYk6LzsYDyhQzzxTQlYP7HfJ64UweDknJM
rTMNGcMgdYm2jJbK2R3t86ur4gxD7hwdG+tm/U9Of+FQ34XLfTimuMxohu/Cq/gxl1ze1KtJo/F5
Kv/rS2qMVUdYif9McKkP7bOzc+hcDYfQScdHnAFyLS7KMwB+QJl3Hf66FKlFfdcuUvk5JMwddUyL
sQ6Prz27Ja6wQu4WUv19t+R2sfJc3Jqd3KScBmD4ApUu3SS+kZjtKESJ5JTO8Sb0GECEGlhp54QC
lbyo+HgjAauH+j1MzjCWHtqiawil1M+udIEL2h08FH9e/Lbgo0YS1eGLc7os8Q+uRYLB3IO/VBJh
VPVBfDaKc+ejtDg/stlJDs44tTrCdOH+BtP1M108Is9gFaHc50ZeZ+bv008loxtvUjfEpAgwXfEz
E0klGeBgzXC66v658FmhZkc+shZcYo/PWH1qetNDkp4jWMperLXLaO/b6T4GTXRxiLludcR1kFl1
26F1+qEpEKrp2zsjRtJCTen4+VR6OV0UYomw+NBt34v4qsdDX6sW7MkdfbyKyrlUGTbt+N8NuSMi
Riqo3cDwhXPSqdeFLzBdgeOScu6/5VjNZVlRgRftKdHp3aRV5O4S0wdLTltywN/sNiQV1ypfWoEc
Em3q3x2UtSIcpY08EsJ9iDqI5zyB5EdC2KNMTXz22MJ0kkZqjeq14c5vowV8/07pggxMqUrYHIZ7
rjq6V8di2PUdOXATkjaIbz/aNTeR4F/UarkQyVOCz/JcoNLrOSnQbT+jVGSs/x3qbBpRQ18jC8dd
tIUp4kIamQRFgaKb3x6oBDIR/j0JBFYZ9PYguF7ueIO2O4gjJte/zn1Ir+Ga+f1VBbUtDZ0G3icC
pU13vDnPiZReGDan6WOgupY3yrSSXA+8JLHZBxOsXjU6LphXUPhrOMV5+1G1+NQy0wMdGpI0XAFf
8PtZ4lgvIcunSn3PD+skHBo4YEOw/bnU6IQcn4wkoZ6/1oGGrQ7Jre+nWilzKgN6oiklRmx3Zqt8
0xWw7xgsFh7A+5bKVCIhfNIbR6fRkrKHGLixjxsVpd12FDU0CKh+nRg0ykvkJRHJRKLw3eLyCFBL
LPIJISWhGTQI1X/WPY8w/Aa8dDnZzC7mXPYP9zvMXZ1AHBapNwsDzyou0haRwo88tcooc03jDqDy
Vp2FVBcgROJW1JsjrMKgOjRGm9Ef0/lbTFW/I44ALQltj4gmkuEaXKEBehAL6Hea4eVgfF7X0DpL
lVUAjb/UdtiWQBEXxg6gEWknB6u0CplnXXu1CCN2BemjYzuWjUMfyWZsZJCqplrardBlmNZFUwh1
T7lbsLMb3N1CzJWWD3wEKCY3GllEEBjJcxHaWRH9iEGM/2jHygtFYZQJO9FAwvUqSlqPe9MOnDm7
YCYo0+x7tNuYVmYeuwReU6hnSeQH4+iAQxh1A11vUZlR5njsHjIgU8dK0XplHmidjmfMH5hnyBxq
UfEkVRH7Q3ZOxBAzLICZ05ks3Ibgznz1xIbaC57BVpbPLHoKHRQjGI56c6Z1YCb0S3coCirPJcK+
2bJ40mJV9V0xk2dQnADnbuQX5T/aw3z3VAU/nQ5hsrn+moE24v/p58uNxxBKp4QpwQtQve2o1Dvq
37lzzl3EztVXWMxu0c5nVAVp1TOglUKmgaCX0j7Vq87PZBTvb2fBAODTq0inkYHYf2J1VmmeWnxx
z+b6NnQIktiaTWUikQDeZi2YngLbk+P+QP0QyF26vhTeqjAQdBzQy9LoXxF0Q65Wu01gGbxg0y92
gs2OeMmM8B04bmrz8KG95wFgeZf+7LEN2ggNrFCtlAZRuCS/f5PkDLfosz8ABTyF72/jb3qUQL75
XlQzBdcK6RNH9mjcM6hDtlsmySiAdS+R1k4E8hS7PO3jsjban7DShDm4+s+xveuhLxt/fIcGteG4
eLlU7Wy74GFKeMqJ6AN0vEnMHpQgOkU3cquSfvJUwMi07Wo19CiX83ccKtyY9KpT0a8oz73R9mFM
h4yPAqhfXqKpxmoa3G6ITVmvhG8cFGFDiIuYV8ZzT3e3WMSbmjU8kOosY7MGOW5IP9p2poZlJD2O
UbeCJ5wLbNjQP/xNG8L74baBtlhQnJ0Fo6b6oj9cwVO7xDjslMgVccjlFBv3gvmAe+muQG0VmoTI
X4jq9yZtdurOqpH4XPVBgipW8wzURNaLebZuhNYJjgfmzCBabAr1fWHCFY2/Xull2XV7KY5Qe9Cu
AtfhRHFa1AmVe5tMoYI0vjtMf+KL21utmnC+DLRvNh3PpkjQTEYd9fygKKfu988ELYvq/SHIVpTp
fpfT+RP5bHcjNki7wtzGMoi/tsvepbRJ876cRa5klk8yuqQ7NoiuIg9ujvh70K7NOmb9HaBGcuiA
FoYHDENp/eLAQNrymCzjQeQRbuX2dxtX9UJXf//3fWf39JfiLK55o5Tf85/zlZxMwaYCi8PMC0Yg
k6zIbLHJBklvBB+b2YImrJoiG5o/Zqdw4lfFst4hm9wo5MTRVIhlvbFdDqtS+2MVfNT3ZvS8nkJf
9uLYWt+CxNg9A77rbs0OiEcldbL9wHrVuAfGgEEPfn4OKHSiVJT2eTt3Fu2yiIXDx7q23Gt8/bhR
ZPGaGcG1CH+Zz1OmYKUafjlj361JbuEolvtDsMr5YdoE3/VFpllAEsK0saEmCOm61ZaojseqWl1s
HUArqvJ9ZGJ+HYR0MyYpwgajolofSoUG2n8KqNQx7ObQITsx0WYN62xEw0kzAMMgaugT56iU3pZf
VcQXdKWbpg4mJw8Qx7bwwve5cCbEVCOP/QAyxcdSpqvqVjyrT35fK7TWElQm0bjMQwIYzV/ZdfgB
36LHDAg6OQkBrEw5GFt2r4pakQMu17AYdqmG8ZiG9xDCOWmbbkq1H8bknP49oLGGfm2uXZmzCTdR
NfL1KzFAHDZTo0yGEPCJA4v3R/iNx6cdQDftijM45zGmRURQ+6E9BfTCgmx0RaH+Cy0MFASoEZ+u
E2b03ETvHQ7s8p+4dINT4h5N4pHK5+5OdIMUPz/EHjXt8zmNIeCYeOcbYF1U+Ii5oVUReNLEkN0Z
KH23+YkTb7rfGOPsfxMq7Ft1gCkLdJRvzD3pXcKAONl4fcZ3mpzO2tIe7JfgZ6/uamAxXpgL3Scx
Y/v3Fjxj/nNfCnM0VpL09Gh3j2K1TYLRWmhOET9lbOuYk2EpWSyw1Lt6eFGEjirdCv/po2dyyrV0
saI4Rs8QA3R79TTOKU43YKFcJVY7JfOdTn+v3YmmEEXpNLWsx+QapxRFHbPCbKddo6gZOdGvlNu2
WOq0wYectWKClPkDZY8oTL1GY3QfHzZ0Yjr+VyekjT7nJXtSiVNDWoHNhIdCeFifl61aSm6uZGC2
EN3OtTZRy9C9uin6hsniWvtbPiFA3kgGCowX0mL9kfbZH59RkitbYf4Zr05CU4Ps1toB3cnRnBuQ
O92eWcm9+7RJbu2+dx9fxGMNHY4sgjbSEnCLsnMiCOqqFkkl9SOWVn4GNZlVmvsnxNKsqhOI++pL
6/OgPeKk9IP4FVkq7VYH2T5eeVpcO1aHX4QSes3TOxpRJrOhQSGRL6F/Z5Q84b5yQha6KzgP/d4w
XVjIIaWj/S7In20Hf4X8WCBPy3JYhOMkr8AL9Hj2rwOxeFh20I+Bqea2dxemmjCaKQrFVZX44OPy
/UkSbMnGMfDXLPfjWbEHoqT3CpQG0O/3BxDdThoQOPdPMWqIBaZqyL8xWNB+7XwQob4OqhXrLiY4
iMQIL0BxHj1Mioai7W0QtDq62wkEiNzWmGodYXdYS/w7g0ItaGeE2e0PCSeHAc045qKIgsrgQMfK
2KBjcbEeM6A+jBFR6n6N2MPeQcorpsufz3WschpucCSyP/bEAep+PCFfmPM3Dk03niqYUEZdyvdw
Sl8JyfSAlZNm2fCsP9Q940BoBEm2HLJkXJva+xIUuphlsUPs/WMeFNhtIUbJSbaTCU5SISOqegxq
eYtEbiq2uyRzy9Hjn/iSY3MjdFjN4a8OXPRgWpDYM+E3hZD0vDiAbr51Jlo8GVeutw3WBu0H7BUB
BVOkV5rhLxkXhACT9DC0Inl78VJMUlpm0pBTGlqgn/EyXjCCIeZKPEWLAEz/nSWGCihRItacWeHk
VPxuIak3WOHoshWKj75e5fY9PEb1VeaSQ5GcNTf7LWooPd7Ruw9sc90soAik9uGdw8JbLOW+JwPj
I9ejXiZ2Avky3gexEYCqEW8PpI+P5i4JxyqZ7zHtEsSHtec2sx9BygeOULMqpIamqbM90tyPTJKR
8KkIaHAXVjTY2Qk8fPdVjmAsr5icmTXAACZ81dTbVCorNRijGR9yMYXbUXOBGsgPI01muKhWLS+s
y4Q3+2J+yC9PtNQM1nYVbSVOR1XVkBkmbd6Jx1EWRbjt3RkYYBUc6J9BMfSNbjzKIQLu2XsZ/clV
6123cbG7n8icrR8jzfN8fBzeeE8yMseCqqZPv+yrJ7OpmUHP8NrOPIqhHxgTHbmS/c+NJ6+iEimH
W1iq6cmlpGSs2aYzWDFKCGQ7vdK88l3/qWYbdvJZ51IrneiIvbOUpi/A/A0OojtYgtNyTglB/9zG
8UUAcD0NH0j8+MG3bYeVkc1jBOAUL+Xd2xK7+0bQ6fYeomP6QngJ4JNg5FBm3SkL6oqmuQyXIcyN
hdYsOTFVxxBXEEnwgYls5ltX2Y9BioRrp0BjdRbtZ+xkFmI2oNGPiNpGFX4liJUS5Hu4BtI04USV
ahWXSmLDhx9NwTnJRC9oOKWFUBmzc7tYcYpsrxOUZkpF0ZjDW44fkI+ssA9FDnb5LK9CYo38Cbkj
uRVxRlkRDMXXciwhn3JQOJYoOJS3i91aeF6RxPWXvYyRx9WN5WIdSnQ4tWR/DdQBKXDSlEbnaQvS
mPgiCYQmqp/iNPlJTUN5yMgXbopSS5Fd32I8TnQMTP8ozjHn264+Dj4K4rJfMCtA3PlbEbrrvaNo
ozIy9nhHgwN64jkGzPJUnj4vK0yYOcdEJapzYRJlgsMoOzAGk00DlWoLicw4QyaqP9T1QhiBZYR6
V5bvBrTRgk6x9YuP55JwXe5dzseBhqKtr8VQ9VYsQ9gJIakbWhhJnOMYFavoXIIcew001Jv/1ho0
qLtUBNl567NpakM9tqSDwZtHup7G3eFsK08AHmk8rLa/JNDftaaOSCRLF001gY/OPtwcinAwhyVc
h7CkxoeSF6cZapVYRG8wp0O6A5RbR/4wMvXoIhFzL39gX6ByU6/n2itOu847d6Zlw6+2AiWpMGfS
3uJLUyy9SjC4UPkmzfgOd0T5aEgImz2rUFa+EJKzCV8WSAqg7qbHIYgjPg/qDhHP1FeZ3MDaV/ay
C1mk2uylTpRQ9eK3+6hGEffIeHVo2lURkheG8sPow6NNf5sarDaFk8eYolpLFv4A6gFYDHKkrtw3
3hFdGMbQgt6t9yfnmZFdX9c1Ej4/Q1mNrLq7rWwbQqxDMtynP4qUE5JsZwMrZNpyjM/HXWePsNHK
KBgIh/0ytZGwA56Eu2KNPPnEkf3T9+fekohKrVgVVD83rT9FhnDJWxCOmYA0Qg9G0JeFZH6loWh/
huOQeNcUTkj8HvqIIL8SSyAZg55MW13K6QcOotqcDPR+xlMpilZmD2hp5zWatXNoEo1vh3pI4dgr
Qi74jqLaLFi+yl1vHpyO904VOmPAwtOne7TvEbg/ip7V+f4K49Xy4tUfK7YKWcjLPC5ImHwMjV3f
Z8/dxXReWxQjEgTneSPzV0X8L4N9WC5uzqlH9dowr9FhfwASJ/5txIdjXqLuENAyoGZfCYhTPK4p
YTjfuDGKxl8FzJ/rYCqYFIkqEXdxaaYJYvFM7QFej7Q8ZUQ/kVacKa3pAOpOllQHQA4KJFnvveR/
LyipzqmzDTmqk9Y0V7Xjzs6UpG+3/9QKIp6W3o0rbyRgDI9rCSuZ4TzJdljLSl24UB9WXxuE0/JN
bB7faLSuAVE5hcWOMLRvMZ3Uo/DzTlq4/KKXZIgc6LcqakNNtf/gq9YI52mjulP3uxORYLQKB1zL
kNfbe8PFV1/Zt+k6l8hIAnIHDOeH4PSVc4/OvfbjQowzyv/RAVP3izsxPqNzPlQ15fuZNWsHwqYm
BLWfYcehga7t8X31REw6HmsshEft5gmALlbHKChcoVf5rkZLAZw8dl0dydKty0a88yEaIyNgjgd+
HSyjq3lVWMl5+tw8G/CWLF9AgHpQMeZ422topOOSI4cunbdG9G9Uw5+hM4TApylMiCAEMdmXsElb
TjQVWWIXhX0cf5ks+7HPlY09NUL0CK0d5UhJ5VVL0OD3xaxiL00YDNnw5T1y4hJajQn2CAw8/cn5
BIXHWNmoW2uMPv5KAJRYEuU7jbNMVo8zLD/YT/CIBi9wWPkVk10Uwq0hK9gg2SKxaNlADZJ993kd
/5e6z1XOkbDKNbNc+ZWe5bvPjQUNsu9vvPqrYX1592hhPef2ja4hhZF/CYvu6R3NI4rdhqF1X9KR
Ii3ULCJ+ehWYK1dV6VCy6jKr7/NgmM6YyVXSnSu6nqEcnssDLzPapW7xXy3Sk9k2aMAUzZbK6M/w
8ibhK6xh9WK9P6ixesgWo76Bv3hWD6IjV9LcYaFCHUJ1ByE4bZ5oiplNeZrUsZ3d2cRx9RqpwtV5
Ca6uFqK/nT4PRs8fyCqWfM36L9bBhBPyJeI9qH13rSZHjxrVmBEIo1diYfJ0Mpq7DmCyL2q+QW7B
qKriNZgYhIlFC4jUFHRk3wR/Y/wFmzQ1cVhItJZtisQy119im3EYPM3hHRk9Fg2HPscoq8l0wI2J
J9bpJzfPD3P5SO1OgLPA5/BFAQM/SzV40AZw9fIk3wXlbYH4jHYFEcpM43ZT6glbidojGxNOUUdI
EJQZg65wvnnO5O03qpn4dTcXRX62Uz0dTul6N6IkQHoDeKwOS2wa+PaE6r8vytf/g4+YEt+VCVPK
07QExLblm3lTu4AWC+wyVfjOirtDrcQcrgGXfVH8x7XQK9RyjagEMp41+7CpfRpUkPyEC1cIc7g5
tNW48vukfvX/ZEPGajDFULEzXBxtHECFvRioF9U97dx9quF2APUCMkPrAa2/Aun90V5yyTDeaBli
OHlgom54Qwns7iXet3iB2h+zAEJOTdUxEENZnp+0HzP7svpzjMinZa5wvmM8Ao0pm+2gkrpfVIY/
8FiPXTP4w3N+BteMSohDyOCw4K3tMLLUnp2n0uDDrotZmI6D/Gl67d1AEMJQuxzJHNuASXhNDZ+Y
DJgTpiMsusFvgwvdd1klhRfzOBbauLnfl2/JQhfqAU5gePDhxijP9MzikmCILm5BIJw/GVBqrZni
mrbjzC3w6DFKQQCkztG85Z2K+xdT4wHL8UNiktuVx7RkFQ8GIyPHWDubiW68Z3rFC/BKwyqzH4G8
/B9oNs5MSaUUegsKx5UP0S0lxf/QqiPnjJIJHtNNcELTEkxloE6DQxrxr8u8YKCQci5qDgmjnDWG
B1GkMUPHVCVmvgqUeod9BidfDP7twGMkp2sO8pbP4rgMnBUDhLnfuCeUDoZL2IQKNZczgtk9WXUl
URJGM7NP4iMXRgfy9ovQ914YBPWv5oTXSNX1gikfHxK7VtEGa++gFAdrQMq5VGvRtOsLNe3hpTub
SQNoOGcV77N33dzj7XF8SJ3HwL4qE59HbNJkYi3JEsugqVvZFANS220TcEYsog9cC+qDaBC5beE4
FjE5iltKxV1Dfo/Kkz4uUOOINKVYcIkkbOJVAEgU3jZNy9NAd1aoWxvjA4miXRrYLQeNl6zCQBOx
5JiISTWTab6nogZR7OhtJYl2yQ//KlLZOsP3e6fG1HROsdtQFBZIiMwQZZBbKcrhIypoTGHgrGXn
WsiRuaRVBdBMmDMVfEn7rya440msygahvzKcqvdc1GGoZA+C3fz4G+K/YtF3gOOxuRzWtY7FGqVN
7yz+mEcSgR+0x3+tp1qkuQviZZHDg6bP2o8zyMMdUNye9fqZ59wTqjwRvJZTRPHdSPBpV/yRt8e1
gFhZrjwvcDW9sxfgMluSCwBGaauOp+QXHRG9OYOdb7iLjC+z66VfJgt6UHbs5Q0UFLonrWeq/ZQn
/h4OPqs6Y8giPTcbg6BvBAuKXHgGPHBP0LGiiljqEBlD71Xs5GoJLpP6Zy16NNntHXmogVwiYxhY
9oLUBHXl62+6hHix2+DKySHezofVultTsCdlN9Eg++RJnz3nBWmfg8H9pZWFsQ4ClZ8sx35yn73w
1CCFuYF8d3jGf1//q4zNDqQXPd7Wwuim7tePtOmuCkWTZr30Z7LHP8jl0O6vrBCT4jLaIRwwZOeq
3GHlt4VyAg0+RKsPgUbbtR/Yj0smw5O0SzexZ+/T17oh2vLGWBVOPqdcfZ3ZzmUo2Q4+bth5GLTE
So2TAHrTHl9hy1fpm0tLkPCZ+Ce3APKNUFLCzHhct0YFe1I/v2HLDbRhnzRlbfjiKhdCjlQh1/+u
qDJ4wlrNwctEbVPz/g4GroJb5CyJ+2UgWLolu8RApMe+HwRRK1i2cvi6EMyFMcK3Cwtnm8uoKd57
jBF6VGY735jSJwTAC+BEjY1dzK5Em46IrJM1L/K5p+NJQYrnF4ieWOsB4Po3/uKgr2D1BINtvNtv
SwiEABy2C474iJbiUPa4cnLmXzHawx90yBdFciELdaxUwcVe4BHpNkPj4uR9uT2JBkJTM94pUknt
9RZ9hGYF96hYsfcklJn/eokrZ4CgJ/Y1hnE00Qe2UVkr5+iWA/9uneTtlc5lbMAN3rEJ5S+HKNpj
fi+/W7RkS7Gul01/r+1McTcElSS/lQEzhUI+ajSpYxl6ayxdkBVuocb9dZXyx3UFVlqKSFsm5Sdx
h+ahy8fcbu8ZRjX2mDw8Jdce90Qlxq157U8LjGPKM7vp2g4D+64RTQvUSF1+1wz8cgi9tFzpR+J4
/0pgyMfRLjh3mlE3gdNFe3jFmeAXjkzifDq577Y4ibNqRFPWOXl2tTwC60+UN/jAg07+aF6gOXmE
3oqJ2iPj2Nt9ntMzxRefUsH277oiY9afUMAuO7YVZzlFcSuJ5Asa8uPIPnw0zdwiEb9xiI6BGEUI
Xf+sBU9phssgMlDqKzjoK7KgW0fjctZTSzS77eSS1m4jhGhsvYjHyOzPEi+pH4EQrNhOHUJNtCjW
uh0V2pil1fKC0+wDAFDbKPW1To6xsgSub2k/Q4lQr5/j1LgnDKa0kAG/C3mB/t10HeHvDQdW/eu9
5tMS8vpELt5yplc42zHOJCbAq6bWwc6qXHZYH1uvPiPsrdjZKqtdXisLtArDSsWDHYeKhV+TQOGY
SO2otHshP7N/DOKvKqsBNWGsl3DtpU+0m4GrFUkuaPPgjajMg9yFVFqx1ce5QTHvy6DXBtwsKA2d
lp2iVkh1JesRO6g/PH3sWV2xqbtoXkurtZSkRS4xc5yOkkWYrsqq6mQZVeZZONxJPGF4Us9ZS1WZ
b6VS//y/TRvceURfvbPSomp50CGsq2XiSHCho17R6KhI5HMsIA6iJcf4S1WPqR4jcRW28o+ljr9o
eFlCn+NnMHMkHUyXTY8eTJ2IZ79XjtwyEAAbHnyRfiEeEyBXrNFvOvzK2g1Jpz3swxTvfQe84AsU
vgb65yiX1aEjN6t0JnPixYJjjKSnl9LIuzt+vQ4J0u2dxdnY/ro2HmI3H8PjbphkDnThFbnBIOln
Sz/1GNVE4gXo7DRBwoxjOwsWKriZdHxm2IL10NbE5kNC30gEpCPQqeNTWXogFClcHiHwTWnfr10Z
/cmx/oZlKqnLZgLqkN3fMOa9p6AVzzualuiqESNsAdCPjWWFAsBDGM9RzxgM7FcsFLI/MlrFPXDQ
Ridw0GgA6rs86OHFiuDcmUJRWDuPmvzJTSo0zjaA2vqviYObqYsytE23s51nzLOPEp0PHlQspYr8
eZyFqZlp0awEWxz1DXLZcistXXLM4/glH2/m2fyD0FOj5dtNXO0B7iQ4Fe2ilx9EFnJ6bNMWo4hc
vPxSWELYRhhsDWbwSym41tm2W82AmiynnSQ4tYsQ7lykkoGwPOTU+AiDZY8nhhOR4095Slt9Iu+k
2cI1xwnXDmrgp1Dxx7wWhIfQem+HRJZOwlaK/4fGk2s0bala7peYN2QDBzfuhd2g6Gx9su/Hw+jq
i8gOQWV5GCBjBuootlIe4eyCGjs3kR5yBNWD/K/EJhdfXLlDz6iiOgZyQ77T2nfYMa70IwE3Lxxn
ENPb2SObGEhDg2LXd7Ky6VxHVohvyn+XQNiY0LvB3rAdmDSvHl4Zw8Sw0iRFIaGAoBL9rg0SsDTg
dt5Dff2UuL9AI7rZm0NXOBB1tY+VvfJXbQgM+P6F0HEOm0uIQ7Bel2D/lvHpUwtzQDnaGeICyC3m
ng1N5ym25PfF9StUqUAIhVv68ab7errKo+LD9ARS3ur/XTiFo+eHbc63c1aLM4zbdE+dHUnitGPX
qEXM0RuKq/dO/pE1NM1FVkRCemTLCZeICdYNGqNVsv4PEsZKqoz0FIWeO2hErfNbYsT9FlH2X2ls
Kv/twv/VWsw77oUW63BZlag1pJ/qF4dwtI2t6IQJeQM0bpZdBC/ZkIxG+sGvwNL4YeXZsFbps3mC
HT8WJSVOkEAK7/crGLt0fomR8ReyMUQROzOyyjoaPMY3wrWvyHucjmdvDUpm+2r5ayVOkSpGN+aA
ThcE8MvtRRK0R2RyxWvJg2jU5dzNB1/x0QIcX+1vbv3bogE6arY9RHQhZkuyTTp96GGRWVdzmUoQ
bpc0LpbC+/3NrcWdQjrM2y47aINbnVRJWpzwt3QJPl7yFuBTlNN2kOW8VKkbDsouaAnULPxMwERn
qKHAARzHVBnfiQuMsJsEJ3puxi02XJU2/hU84mE29pUru95tc2Gn/z2F0uOlKuZzeTlcpkolyyDj
mdh3tKQPARllj3czRh5CydAiLBCK8BX8NQBskaNZrZwtXnrxOZuT9595TGpfYND9W1OLdDLoWCAU
OJb1r65E0cQtVOI52bKyJmKZJukiDUvH+R+ZNYigyPi7FLWbcaLNkuiZpgffGWXkXO8/oS3/fGag
/b9/XI/6qKbxsmNek16EmdDWSgDrur1qLfH0ATtbFxgGAcuM2F1GI0dWbrZjO5ImpWFMu1lKqoMB
GHc32kQwMZY0jpgfEyT/UU9gbH78XrSlsOghFUMskJivl4HtF4AKxdZiviztcLroDRu8BHU29CeO
ynrQzVGK2FoX8vJIdU7qwFPjw40/8iO4LBzD84v5zEIj3GoToX5WIXz6GYQFu3gAOqOYyQG0Ps0u
fvgUudkpMCAlTrrAxbNHqw+pSact9d+0Zt6uCa+F3RzlGdPGdYMkFQdnyG0TU+nAubBQwGDM2lrJ
EljmcpALeKPC94r5HY0kVdJXTMr66vWSF3OEU29h7IEHUKz97CIrobMErN3ZSvwOTB/3bThMrdOb
mu0M82Nu/J/PcI0aK8N67KN8l2darDcbrEDwjOHeNkFF1HcLwHHtJpgLdyC7FE7jBSSWZknkpTZg
GnF7N9+YMcSekGP+TxFOS32lCiUlxc1uNyamCAolRs60f1nHUsbGVVgOEOufH4nlbt5vH0ERmOhk
BvaBItIiVhK/f50R0qKSHExrCXFzQp6tXNNXWHa8dPkhHI49SMgIuD78O+JoJChXdyBWWpVZO9F5
l/LMUCYOCMw5aAYCkunbHEDSRmsOFQVRqRBfBOrpE/NZjBLYDEWAxVupj7Qj8i1n/mWtutgf/qcv
A36uqZdGTeIu1B0xRpPsvu+lj9IY3RBO6FQzAhQgtdkRELGrJpRE8RM8bSBSMQEqzcbtVi1yHRnK
+2rej9JSD+Ut1E9fjgwVk2Ms5Fw+RjDPrkPFa+Nf5qLbtsNyeujqg/HLrZlFxi3tSCnLJY8D4ZaI
SjfPU3p2QBT5VQvzQnJT9J3bXEA8DxXu2MklORsVSU12U+mwI+awXyUjbukEYEDdPAC5xpDpb8j9
m6KiF/+7B1nsIjrxg1piUMaNsYXIhl8WGli4FV2jWkhx9Vf0EkJTNmDlGuo5JmuNXeCxgQBIvrR5
T5b8FMrm9Kgkjqgq+iXoKgMByzlxeTiv/97x1Nwfpaz40P2Hll5iE2AfIDZyAvZzifSSpKvyLREd
Zec7NBsPtT/Mvlq01zS+0AOMwaZn1jk5bCHk5AeI+BfrqWn/ZZ+tdDJQxvNhgEz4w39rfekIOeHh
xUWpNtIHoP/nIWm74zWYyW/zMyNK1W7HYoE9ADHNu7HlBOazUmsLhQ35cpYu3ssnVEk0E5cw9uI1
y386vYadsVKrmi+hgXyMXQFfZWYTBSa2Eaq+JDPCfZp3noHvAtbqPXFH8mkjvTPrpSMr4bZawXqc
rfBc0fmbCtoGyZ4MXM1wQKr322hVApl6MubiTJpB2SMzl9idRIrIgbm3bnfWHdgEBoJ2b4F/Gx4t
6LsGS0W/AP87RqkxtoBHdhfrcqL4J6WFSGGyIutm7BoD7P3Rtys8LIgj+NnP8Ozyez5mIU5tfmkM
PFQxpB1lt+86J9TTVtcWOI/R1fasKKhfdVdqcS4Xgd6dYWciPxnd5ruY3I4X4ZIgl0/LvfcXGZhm
X26RyysUJld3oYywVU4ZYawEKK1iMnAG4hpFvz8+lvY8b83b9YkKDXuhZq1Ikga9/AYpdfpQENXG
4YhrSFlCKrjPU4vuX/KCiOBVZS1GdbrYJHkOtPzHGRx8J3ydq78/u8gPuKGEl02I0xNIgcuTAsoZ
NKkTtgijXlGCMtWJhpLtcpBku+o6c9niQ0M/P2wUcBmT542NeYvYLoVSLyPv8zo99Bq/8uK21COm
/Lxb84UzFq+C8jGaoRoYw3MqLiPDALpQWsgRFC9h/McCmqxtcNOVqHhvQ1RKp8ec7m9JBA20EAXL
QXXpgLdGycYJYP2YEM4R0wwCBfKBu6E8RJo7Ntt3DMRxkCi9Pe49YztxHPJ5gSk8haQY94LjfNXg
iA+ajoGWoEqQBZrq5Lj6ApqtlG/PyjU8rfAeO8vT6/2ZYF+wo4pUIgvOdQvOIJ2ZfOMRYiHWp9a2
JVlBFALSg8EdJCiOLo6WVy/tDs22wtGK5yqj/VOefMt5Ia/lsJmlIDKThQlD/gVxO28i/A10fPYP
fLhAq5LFX1qyyNWXsvHOfQfQR/eK6hsHf8Xj12wxkpqGn7PfdJNy0nucz+nRRd/4kkj3li5ubYBj
Am4m94txrtmTCPDtEWVALVFrlspcB4NZpbzha9yBotuaJpQlNDylRVdCiH1+QF52zHfra2xlpwmr
uwkEc6iVAjvUAZL83IUxOPkNEuIrQxlGk4HYdJ8VJxR+jg/PHHPATm/O0cayiit6vqOxuLPjZZzP
6eHw7WZCfCne0XyFrVl0JWw7RDD8sPcH5Vo57h+msUoP1dYekIK5fEEg16OoMtVKhkBo6QGxP3uz
vTwg0K2ahdBAyno42Gx/JUPV/tjb53qangXZcsUGbaMdCYL0wGQM0le5XpKTat519uNIPpx4Tp7N
PXkj6mqwI+OvZii8cwhDyCksGuYKmIRSusrhyWs5vmAjO2kNet6qcbWolDxbm8OzGtuMjBDtKwf5
jRbaKyUP72sFaFJiV0c7ez8tO8riA54yl2p/74oNmF4s86lsh+QMr9T0JKhJ13wh8YH5/OcoNp1a
qzc1B8XZAtbRGmHnhS3WV1pgpb15B18XFeAzK6Ss4tivLFJ5+k4re9DQHwm1pl9bDv1NWqULpbTl
jC2NZAqlZREBnRG747c5ILfkHK57XV5SNhm0Iz992BIe86bNvesVoh2etrQQ5kCCzFIGM2zVqBZ1
B3AQuFenhe49nTI/gMESggvdw9XTBMOMwu/ALnwvqeLYRS3XS6g2/neH+4Muh5sce4GjQSqKe8hZ
70Vc/mUVG0iZ9PvbdBc0oos9NyT6XxTEsmcgiPhArW2yWRfPsWb4J7crdWrVh5oJI1XCcudDlLVA
HAP8VTDeM+GmKV6bGCVYNM5JRcmiQfrSHnZdKPodO+uCMa16QCuaFPPalo0BE+Vz2KKTXAgPSWNL
8KjQHWvG1PLdmZ/0J/zTy94dOcDUAav/wT9Y7xmtk2txBUF5Y2wObtSqGRPNCPqfXBkdK9b8pNHw
uiuE1Q8Omq2TRQb/Us/gUprijnLsAHHgGOMOxXaJcLtoEY+wIewaRRGyGIx9FQwCtLxwdl6BMC1b
F7bLHOQBES/lJwAG/Xd6hp4N/oZZf1bDzoBJLepWityWErpdFPIY5/j5BU/44JoExqUl42AtFmmj
E8/1+erNnFf9XWHiuPWekDd4kyobPFOHh50V9Raf7XoasCPlcesWCFNlV6WS1csusYllh4Zb+mSh
H5+LhoscgQX5D06URgxLev6IaWHHJblDnPs1VC2eUv+XX5MyCH4KtD3RpaHjK8F/OHlcD96ZDLiR
YhdL0hdfk37QrTYvwkBy3ok8ThgqCtYRn+73dR7anPXe+c6mtm+DW3MA90ry1yp6nKmLEteudGYu
XPpaaE7Y417tGTAR9YRG+n5m9E2h6CQmSrJGdXNFnZz/nSGrAuisqpibm5wZIxFbIc/UU8gmAZmm
FLYK3obQRF0FI431mE7MUXFMNnekp9xFT2Ex/blczvjXz+rm7UZ0Grs7mAdfEKUyL3GT/QYwrOpw
snZOex/9fZYPxg5dmpMHwXDzkR76BlvjEQoP5bbA/unrA5LMKzO+AqKBtPnM+YznRR+JgT6G7GiB
aG7ouy+TckISJK0+HGvk6ZE9nBvVDSEBgS4/gYA1u2ZGbj0gO2ty5Tt191Uklwjg8gWYPGI3wyJC
p33NtJa7HOBV6PdPBQBaHwhj9ORdIvyzU283BSOpkYe8IiTP0LWU3FgAn/xHth9iFj1rat9j1bUw
xCnzE2vQ/9QbCDcLVOWFUJ9I8gdPSwaQuv8eNQ//RE/ju/TFYXfb4AKg8O+E+90XtDbw2PBdHcJt
hae2UIUrabhwH96w5NWeSi6/VRYpyRRqLzMWoHMswj+3a7eYQ8xDpe5r/zHGFFE21AuY44xlCw/C
rR+HRWX6jRoFKh4sgvTBXxNPZEefIGovSpaqtMyimSYh1ByCujkRgbon59QZOjge5wTNpc8tuy1I
ojwjdb/F/R7yDQtGMfV7SMkxLecCps518ADunzWwBDFMkkiaXVSU7Ae1MeH5HlpMBPVlW91YuymQ
xtVbaGDYyPrV+ATPGG/JHyFtqoZ0Kh2HHZ5VEQqXbj4q8Gm6EnWe3bI/hbGSMsoadSGXG51aP+jS
PU2wof1oPeZbw5p8roxjaGgJN/ETfqzZ8NG700AmZvM5datgGWDnZznnYSWwwyYxjs7/zSlAQzzC
KwXXre/SWWQSmWorTPgoWHk+sZYJCLhlBSTMMru2Plglx/qrxqU0Jrx8/raZ72w3nEaAmk18bNwb
48LlEIbXSsTxzEXwoAVCmgS9fasVm5w8n4+g+S6Ze6oJEdu2lTqhIQeOzDTYyN8gpU3qOpXlOekt
TxXxJuO6aaYBZhQKLMg/kcJ7qQNa9TofZebwTHn3Gx8z9TmsJrQWdu1rk1Qq7L2qOQTlq8csNxTQ
jh45GUU8oLc84qo67gioxQ3P6zRB8jRW2mTJeFn0FHOiX8urkeqJqtiygkCwC458iobhRRgz1WBN
UPC1EMnv8lAbS0ZG+UxdnsOXMD/fOZ4VqPr3deUxYrh5uh/QK4oej64ntG9LI7p+ICgiE3VlNJY4
4k8+QeJIBu5spY+G9YpJrdEbYuKEpw6hJs61YRgAwIOqKjQNXKatXyCwPE7poK/qyUrD/je0D/FF
V0I2bXTnjFOxPjClqfqXFcScVNWVJ0staqo67ZUHxrCR+RGBtv6lkU9D87u4PTwSj2bZ6OATANo4
pt5TogVN6Frey6H01ta0ju5fZqasS/v+A5j5AxzjxdBy7zNObRk1NiKTnUnQZPttxaP8wgSzN8R1
FC2O7Eg+m5QV7DF8On29g4RixzpfYpiqf6rpJVL0bMbyv2NIa13R6hMoLPc7jvcJuFk1+UFQsKW1
V+NJLWYBWZFlo1oaIDLo0KMceGDhFgd4LWniXhp78U0SDm17yhqd109BIBZ3h56Iu2OzgChUnrTn
Q1K/h3TJxoVy472g4KPTqo2R370ZY4Yr6oZuntz8lAlRIfCsH1oNdVEvmVaTw6UYVUCVwFC0Rnb1
k8hgHNkEZ7+hnfeGZqaHibIrTxDs7Zv1n73zcyJgdEN7dLn2vtqc8QKCGcvx9Hh4/FU9qwU+skAo
tCTyl0rjp6KybMIKWjwl8C1cAjHR8GmaxBG/Sv9wcAio0IIBtVR5Oz0OHotTWTMxwqEcMzZQh2e6
XfvRmTJdPErPO0cIJwseWiUeIPX2K/6LCIqXpwSHhEGgRng4diq42Lum8/IFNtytMuCyaD+c8Flu
mj7qqvxKNDg5zaBmTW8NZ/mHI0epcsW4rfv4yDvbsd3JqfZcNXB6XUEmAxOF0gmOA7u3ewentuUK
IoYlU/SYwQeAG5/8+583AL3piV1e7DT8o+NHUujy7AmyCWNqyGD8iu2Gev/WbKQnjBd9N8l0Ria9
VeNqpNc0m0OhvAKt8+HPrrHgQPXCRushvAgFfq5uOukRgXe/YfJUlAGdgr4BYbGHgNdtmFgqmKuj
gnYjdQxCZuHRqI4J+iFaC7e9HMw7hNzPyZ6fw2hONnsi3XLp7c/aSENa84PUtN9ui0Uicnf7e+gz
KDaXXOZZr6gWXtzFIcDR5fxzvS/m73x6BHU99mgweF1M4MVETp8KzOhpEWzA5qcmkL37HvpAXyMc
m7qQ1gQPdPgQiv6kNEI/UmuFs79zuY/33M/YSR+03oJm4ht08M1qTgL12B5pRBcBfeBxMNHMcdQs
twsb12AD+FZpvVAH21R7jiWzkANkoQA/6dJRyFyCWGy8w304HWfoTcL5NuVaGbcWHu7MDjWPj9zg
nV9wchgCPcDwZSgPjzlZwc+PcDXGG37Z1on8vH9Ige/7t4yDyShlFLxcDSRR6KoLbKmBbV8HI5WI
XzMVUZckRC20x71PVvMPf3BilsJiQhE/2jkk+T7LW1Oow+Mp6yz5/cdS2f3pEhJeJeF6Jjy1KJg4
m5zewYf09IwAhR2X0LwDVxy2b1dWtSLNYu1WfyJ9p8TNRblrcOtcZWcT4fUcU0SNVkYFhVewQcyb
0rFcQL5ygG2A/N9nhzZ6K7UPDPB7pxsY39JjhXLYDDcNHOKgMjZioiUx6TxeIO5sjHlZi7056j36
sOcG+dLHhJccFaW+nheLScucV9vAX6ur7AflAue05qXFZCnER6MqIlPooPg/MhoonO97m/Qj6oOm
OuQgCJ5VUOMynxqjLfRoaCxaVvWm0IhWrx9jXTflZxvffuBJh2PAhJDZfDNr3S//LrLv0ZF3g1D2
mUzNZW5yo/hVKvpZtZo9L3yWN96BW86OkVcbdByPOWi0tMyRpVOK8QZ9Vv735OjCxsJWsHJZkkFL
LaiGNS9QFr/ko3Vk//08FPNPtROz9PpWo/RGPojS2nKCU5YTqtVQBcPbo9tEwlMvZPTl12Bjerr5
wylKAv+CxoxPAw3d+cwL/gDUV0oSU4r2vN5A7iHZPSOc1D76Hx9hf4l1QyoPlVp7aTUUVW0ExbyZ
LMC6Y0WGGF7+AWXTmIZnBEpLk367RVefuE4GcgyHXwSZanyNXMtNERNdaJ10Uz/IJDzr4U7GFYvk
llt8ly7ICiE715cUCeqyZYjG0lDeIP7yVNbRzUpT6m9twGKu1YuBpPoUKpZL+j/+fwgjKjsb4Bpj
4RUVir08hZMaZlhhBi4sK7uWvXOuUUTqBdpRqczTLhE/87ebLOha71EyekGk5HjNlBXJjniXbNIm
ME3ExKIPW8Jg4VqSs8gTQ0T1iWy7BrFZyDhFQab/Bhs2aZm00rFQ7/Ip8BcFHhbmmqysYkl3d7U8
14EKJI38pPO9jt3cq+gYNd7DOU3HYK3U/ER36VmlwoKJCxOy8AiadkCECgQhXTdZZaBbUdnz9eal
bR0uTeFR3XPbtjhWCzHFjvsdEARaMNB2Y2FbzzjER5l0oAPbs3vGcEwxQQz0nOhFmWKSNaGdbRBx
yOu2WlewIyKTjjPcICVpWhQc3Msv95bURbgA89iH28vb91pZO/c1TGAD7Kmt0gKfleCzwnPRmFJg
X/TITX2R7s7ytfynrzPgfcZtZ5kBdteRaN/VFB0vyoLOZcIOkypRd5ma3k9qhGPUs6Zk/fiEtR0B
XbY7dNKWYECmYMuM1SLLPZthWy0jtH3LJnPuhYS3Air2YsDcUzoKornTRCCzL4QD2wIr6OO2GuHs
lI/waWoRnVdZASeumeWq5A6qkWT2QXDS8seaQNQLOwvmTddyk3dqm0sndeFpSZAurAEZ1Eh6ZHk1
K6DRf4l0lqUn85F7Ihyq2G9Lv5lbyDaInuc3tVR53Yi965b/Kvhq6P7xeY1Nt3J/bYp/10BPTSIb
/iJcleCcK6cOF0ikqvp1Zarr8ultnR3nlux3PKUxRarUw6RMT+13Ul2jQPdINYF0KzZ3R9cs24CC
c3gKxmhuS7TMNL7KPl6qHD7Rvxp06/W4S4Blex4iCrYJNK95RXo92GvOm5rvs0lKZqqA3cvHTM+P
fw9fxH+GC4OmXUD19vobwIRaH1k/BU2NggKQ0qQYlxZiLjrwsaMQfQhr4aGNup2DrM7GjukEIxnT
KXQcqPZGUzCOvVzOOmFI4vmPmxu9ltfZTcpbSZGpK6X4yRmtfJ0JFMpW56CYCcnWC+tHrmwa0c0z
LA3f5Sx/WC2r4AsWticon+u1IS7zchl1keDg6BNQREjfFFcm4u0OoPdE64ygl4ckAb+wSekW7KJ2
rzOENi/X5X9ehmyCSllD5gkZy+BZpCPOYBTRrORYv/APHwJgkSudYEE4q7wmH/8uDmoU0A2qOEI+
Dg0cG2D7tX44akVHqPD81O8li56Bt8JR5WuGrv4PVdON5JYD+yjxRWJ991WVWDsNEa+xtXIbiecS
Ac/kqMFvWJE43ny7BPhf+mC9JAtnr/ixSK8DDcDRntznbVw6qaR2NezkPf9+hY99jKxpbIcbKJAt
rXcI8WG4bRijvP5p33pSkBpMg/zR69lYgojRWsX6SAqouanPUKx3I2dP5EOOzQT9Jedsdc8+KpOL
k5Ma4e28nDmhEXllnvAKEzgl4zpnL+SZlBiuJs9GIZVHTHSUB1uhQbR1vYkVH6jZeD5z850SSr77
/jas0Dg1q0Mqw7DkHGhgb3dJW8HH2w+tnrtAD/2w2UqummDWRNHxyGKRkXdf6TLImJfD7tNXdBIb
kEo3oiaYM882LyODDXzsPYBqh0Q4lnyYOq2YLoTxUuToM0rKnChbWAY2dOLTWBIyW5T6Qxudnc4q
gH6nxxNvwBxE0vNJtcSY4DrrIdlyQ1ExQ66Ipb0TKVOPqVAG2sS88Y3zE0GWS442Q8Imgh+nHZiV
9RmhePNmRt1u7W2BhP0z4zUPUzBTGOGtr6BoM2hYcts6jTAuJlUmLkhd9z8OKs2R+MHwUEcRdUbe
5N0LYABtH2w9kxesYzJxJtEqevRP0ETTP1mxe7acNpnmeeZuXA8s8nC4amq6GtS4xuQ1Ga+KOb8S
Rh3QsHSHQ3v9Fiifkzb0EtIEgxIsD59XX/a8uqsrLRQeUpsJe0EB7nvmyTDUG5EjEFRVNxGGb+8R
ye3QbbNiApOT0I9RjQte3PgAuNixBYgK95haUhQ5F1USUXZpqZTJaYqH4rOspVcqpeLBD2QsZ3LT
Te9HV5P0A4NkFKmE6eoe8uLGwm/9NCBMy9tll11nKx8tOLjldgIKgNoPlB5wkoKEshsNYI4bANPw
XavdSVx9qEyo/EKvwtyHb7HmBRX9jElmxnfdfd2lFVx9zjjyFlA+O/61R/+OOR+HxnnaP6DDIQcD
kpAFSBsNaIUBAYif0CoX+ZvtJuDYMlh3OPlnKxPVWi2YOAersSpNlXjrvunkrTwuCkZ2cJ0hJlZD
UvIjq+itrHr8a7a7dnquf9gD4lgJfCkltxYzvn5oJqIE62f4TG30tEF5KGy1ifmHrq9llZlqcPAZ
oLNNLRQDCaS4RCMl845c/GQOGYF6F6v4IRYEUAahcDd0IvjJEoUQEr1pDALTqarljjhRynm1l1ku
9ZREC6QIQ3tN8nNb5d6lwNzymAMXRtbHfqlVC+dzNjlL6hHkDertFJ+Yw95pJclKcbrykd/rvcm7
7+9ACvBwTWSidQwLkB0kzOzK5l/wXkK4cMc5DK3ptWAXZZJRARjKONwSej7qa8n02abtRzekC7kw
q14ASFd/d84YVWl4R2/fpZ0YJzrHAuwMEXerfdTVeqQqhEl8wzBnNWZTr6cItzvzAj/rkLqZTyA4
89Zu29Kq6bkgqUYwV7phy/C/ILoK/wZOAFgj5a5xclodV3Oa0WN5Hrkr3RhKCb5GtIhD2WnGh2zS
SeDKMbesjcBoK8KlP0ELh3JpE4SKYmfBGIa0WeBllKl+tE/EIfWjh5pq42vffDnkgoRqIRBr+WK6
EX15R/DYfv2f5VgDsFsiC4mSl/3JUpVZspIuiRjAV/J5+IBZEChpUCRIr1tHQHtS8s5ykcIfK3q9
VZ+vT4MaPiOodXl2YIioG7OVh1JfAGdVJAofgc0Gz/pJwTO2oc2mrWIQz0ODkgHSi91ooBEDuCzk
BiZ78Bw+65oU6D5sKXnILogi2SuJn4Py4z7S1Dl4p/ledlbuWox84fe8Duadd4d85x1BOnPWmSxc
3ryVYds2tx7hb6+vGVKqDVsDheHTCRLd1pnCIbgj+acsIu5O/5Dg93pf3T3pyknSfDwNZ0jwprxf
lKpg1dTiNHnKdAI1IPcu7h0eBKdOS7Wu9qJcriCw205aXM+QiGSikTAajnUw1cJiZNNEZCKsaJQq
tIGmFtCTRyWIKbWc9EPdRyEx9/WQPsdI9RjjF0RsrjBGJ7IagAdX/w+2HoMpRltUrH4Aw94OIfHZ
RUXArVWmsXE9y+0JxbyPAb9qo1FavnUqVDpang8pUyMI75KdKsAFrsAipop4CyAWYSbfw4Nxnhxb
OyJGUT6TqzUvSNLJzCUpBGSYpIkxcRG+FwMkLig6pjELLiTbmt1TtSXoTLcfo5EMOJvRU0QZb7am
yniyt59dO5SvjhrG/sQcKYHNR8cQ9lxD59QoURapXzriEWDVEk8uvSuu0+UpdBxv464YKFofB4cZ
G4ojeE30O9rkjrP9SnzjjL4Fg6Z+YEKIAfXlEMsUAYF5jkZP7Kg0oXYGWDq8B1Bx3N9bG2p+XS5O
1cNcvq6iqYkOxuFUuKiHACEjVjauKkTIt2TumZpiDSF8tYV0ytf2wIlt3bTQFCDbGY/TN/5WTrI0
/bf4cMqS6h+sGQimSMhnoHWOAAylg1Cw9dPOlMj1jsJXzlcrG+FkpMwy0/zPtggq9PqD5yFM3bE9
5tupavEwrw5WmCPzFhv+woDS3DL5mTiUgm5ueuMpNBrOEEPkuE54YBzUGfuub0AlTKCknrueGzUJ
WOJ3cagCeYWOErOcSYRPaCIvcQ3ARL8RkxJvuxAUGgc3cjgwp9V1jqIdy+kQIeZT7A+nE3MifDDM
gseBmlLpoKwzPvlj9epH3mAQi/9dhN+tc1i4eOvAQxaDuXez60cQZ+AF2Dtc8E5UIfDiuvb52C9w
zIf2DLNkD/auW5kcFuhE27s690GwsSwPalwWT94v/aDAQzIbY1G6cfGOJTtJ66dMrpk3OapoB/D8
6fIQ25T/uSlean65ZyapNs2Wunr61UwPLwj2MT1uqkJ3+4zwYL2MvNRNhh1l+geqPIGu7cRObFHr
HuVd/wzi68AH4XnMUnU8bP7ITsFXZQycxExqL2ECFx4VVfKFIs6ix5bj09txm49XBIw9nup1Ro4e
y7Q4zGPl1cU9OCfme7tIY8Kf1J6uUOqU7mayX7mLBVqM0EiEZ6OqyruZiui4Wdvpi9d/4iL1yya6
FOtQ5WGsIYynj7XSs8sWIrca3s2x9O3Npeeb3SmydGhAPceU95bTuc0bN1akm3eFrtE3/xcWqVv2
TpWweFBHgLQoWpizi2XiD7vHP4QaLsw5qAULtd3gRkiV8r73/E/fzNl7vVHheQ08hDMFqp6JJeZ/
SwqJfx+QuD+HBJ0gt8ckbGv7LA9DZFZe9FAek+fnetOjwogLfuvOKmLtPM2AEEfeKzD1WyF3pl86
VijtDwRpiL1fGR3Z27eVju5qkNgFYEGbUUar8cvkKloj6y0POv063V31qnw7mAigcmhKso9wPxy1
XlaFvzI/4ZXhtiIQxfqosZsJlHs0OfdOZPQz61xJ/QnFjA6Ak7T1nLXEtX9nx1y6U53EqGVuSD4h
YPEqgXYr5LxGR71ttIjFnVieX+Naz7O4gSTzj6qc7e/2Cf68ug4DvIyyZDAokl6nMv7L76XEtzJy
FtmhVSAnel09hfePA3+U6a+41OXAkmHg7hNiWwNtIhBCb0qDGat+j3ssOxKydjrPuOE/1GJXkHIw
AhGBw1bOXrS9UkiJEVYgTzpUEKN1mUERD0XZra+5RmQOh7pPpJxHrnVMKH4SYwuIEC8vKXQEtxIJ
kuySZEexTK4ZhZPGJ7vs2WajlyQHmFiAiGoeOsW+/a2017J/5gsKSMYqZau2PflMzC1SdxZj9aUW
pYXo7unBxKD8w1Vo9qE+HcMSmElNS4JCiU1+ClxhFuKDbAjeeSNir8ryjbBhw9dhXx9mCiPE3fub
Mq/kDVXwRux+7RGsHeEbfrY7tJ3rkqvLy7o+Tf5bfYikiH9gsjDbj4/DAtEqt/3D2ibCqX1tx/nT
i7d55x6/3/P3Pp0WssCpIANy9pbxCfiGtOiZzU2DXcn/vOkb+f3tkIMXbsHqbl28sQZikT/3fQsg
1D85DcK/7qK/pP+1EKIdXGsCxhYT6y4Nwh0BobGt0DSri8S7vFuvukGKuQ8WZ4foQMivHR6vzax1
SuSQyIKuFGE+uevxHhNO2cB1Z7cwMdCKcQDpu/k04QYvTWxxISsroDeSTTp3D15BHcAjcEVO3sFt
0qKGvd/jZ2iOR7jELaPfmBT49BAZ0yJPq8WHTx5s7BlbJ25q0QgZhD2BHWt4dI1DPjX0wTyg6Iyl
XjdHLOz9MG8oYc6OylY7/tMb0vItLyeLVXRSpiYDK3P7+nOlqL51d7aOrQjffQw6wRifX6uMjSoF
2tlmUej1MDfxeh0/uxP2Q1Td7A5hHgIIwuw38yu72uwBqokE56YjqUE7rZUUXoDVN2IMTZDHACWe
U/ZS8SdggvFXT56ScFm/KEo4tUJ2HPXAeFzcHVGWHE9vbiyb5elKGxHgIRYrnvyP1uQZvYP6hcoD
C8xED2dwjR+CzreBsKp5kI5Aqitgru2FkOg5MknrvydmgRSdh4kax4K1lWm3KEXMA7fd2WIccYPH
1f6EHNvjSCZFxPTWFo0oH1NqTXR3OvLAwMthaYM3/cFAKzXfEp5YVmeeedIE3UPlYBpLIW88JbIt
tj1DSnx1YfWEHxIA47A2NYfunHX8KWyhyTnhTwUJdsnRcI+u4JLZTNufY9o3JxEA/bBBL/LnUK6Z
i+oorIIkbxR8gM1NW1oV9O9bDt60GaSDjNEXkYMUISZvbymFLU0f1777nZJsbx4q1B8TY21ppmLY
+dWA+Y7ZlrB2yA0vWGBXxE4b+gBr6tuPTMDkEcjbcmDtYlxR5EWM95vpnNue9B6Mw0O/S59lhuJP
ncQq75pIlzEEbOJdMqhoBOhbYC4/ceeVs3R4VcdT4Qn/+8ya3xS9eXnsmE2rJ24uGdku0hfy0YiO
zQgco+mF0kcnVMukbe/UtEJJ8AgfTqUlbKYvjJOmUiRm5vXksHmmpBXqOwtIAnFQBs9jeSgfexhp
SAgKdhy1oE70cIu6E/sy4xxySHtNGQmhoBUqytoqnjA3DnvtaMq0oQ4MVF5uNe+TRPAJ3HKE/voI
jdSY+Ql2zKNEUaaj9+cL5vkF0h21t/n4MGBw9k6XuXedycDx3roD0J7YUmu/nEyPo6cLfkZf4KQz
AUeMoYUlVTSETzTcWilHgw9wJGYwbkKgdIueOE9XJ/vrERLjKz/2vD7Lg4BEE2Nh2X80LmR2zPL8
Y21UIsY9H8kSuDyuUngLwdXAIe7zpl2ejNUU8tcoMLaI2JYJ19pKMbnNRJyDyEmsNC7Ual1AXpWV
Ua9VB6aEbR4NpCZ1cNGU0toSfsvvrPo96g51bvF5pn9c1g0+lUYFuFIygKg+WuB7UVutB5jcjZ2X
S0mMVDnqii/KhAaz8FMBSaY4BNo+a8FlWOv8L9KcaLiUgmCh6EurWklvDDovBbyn3sCGhm4rtXGp
CQoUuuCwIZrNJchTafVjL2gt2GeqkG+HzdEP56mxKqjDcaeXXr7SlqNu/0E8lz0WsBVAMPgGHiIF
ID0XkXg+VymI7Qc6qBpQV8JC+Qpligo3G3gJMo6UXYyIhIv/Lo7LaXq8mIr1ttSt3uectQJK1Gbr
cviC0qbllBaggknrPBomHp+GqI04eGYh2h65SyYRqGp3+TMJ8VbCRNIAd2wgATY5+Ltefa6RG+Cz
4uoFhSfdbhUEVcX/wvU9dbIvYSV7X7EgRim6G5+7DDapC9s0FrTlvh9BIezAx9/xVCvOsALPtHtL
KkQVQKHT9GzyMe+pLxuAfENBd7bbjNIkHXs2ff4EQSqHrXtY9rsrCnZfxALNX1qeCY5/Nm3jHdzD
MOmZwCDGqVbH95iLr2WE4TZiontZ2KL9bnMk9dh169KyzCLQNnAdCvFknatY8XnbBLilDOTV5NwO
kjJpeWALcfIdpc/NK2IRRwVt44ejL0HmXar0XB7ddtF+EITCtRXFytiI/Dq8FuXVKahwrtW8zz2p
o3OBdE4D/FnyG12FKPYpulyqjBM8mVEQnbGI06YGNyND/Kn30uccgbI6/x1f61FA6ugwlZ+NW8u8
HAUEhmkLkeYIYYj/d/Nd80oXa3tVEb83a/ycx02lI4yYf2QSw/K20l7srwRhWg1Eao/QUJQpsLqN
kOHnThKhu5yt3oTVWGt+fuqLOD41TNjdSd7yH8tZxMXnOrv44i+JoctqDk1yRI7+2aPjhjVj0LPn
v3LzXDi1gC9IrBMcxkp3iq7O7HhTKSrCvrkohxY3mNPyEDoDQcodCtazv4ZtcRWOHv8k18xtXKlB
sc/uamI0/mgPJK5jB+DH3FyF2x2WKLZrpwa6B93oBlosLI4s42Z1VxwpvQ4uvc+QSPEdUvz/RBXD
mnn7RYn9uBRaqumGUNxoJZ4ivbZeH0BM16DiyENzki0ba8OB639/4zRz2ygw5DYhaD6lGkbEzuj5
GcaKw26IJTmQi0mbgHjl63WeL35QTl4/BhV7e7mMVXC4N4R5AMnsxViRT7MK1rW+DoBU+8Z8kXCO
i0qQoUtayVKr+kCthxpEMBQNniXRSKzP5YCmL0bec0IZ2madZ+dnHoFQkQYqsCbhXfAXgoeOL3m1
ZpVxr2qjj/26Bu+mqi7JNNk5HGA36b9PDJem0no3IZuLXlyb2BLBVVnXgbvEIPAy12aNGjOq/6IO
k8NDV2SWAR+aKUYNiuMmAofd6E1t7KSTbzWQe6ZDJQ0m8BdYJMDptnzvxH4YZ4OxUYg3M3FHhxja
6HcfvHL/9AbqVmZAtgmyiRITc8X2R4ISsJmCbCNugnvfY+lbTdFFfagFUxmIwLIgcRLKLRkDrPig
+1FAgKbubCMXDkfrlLGORTukyJmSr3swD+sg/SopiZJ8BxGsZNs8NfJkiGOnuDgOeCLKcrhh3CdO
3cmfKIBsNR0HalmvfeH1rS5y+iRNiiEZWIaJjbQ2i1NmGX9cQ7XEuMC3MXXyk+rJPBaCLVu7BHLB
Xg7+4IxGi5Fs3rJITijkKfjhFOhIWv/EpmSxYSehjU9Mlbxpe1yjGIwLQTYk7+9Nut9sR0Bmmw6Y
z3KGjzNnEpfowgzmEeNjI0dqalbfhDlYHjP4Q9Ph6m5DSA+YT98waE3+/9Rnx/pofMwhg/BPQcLf
0W2YRDYVtJP8RPjk1uR62yjz3jz0j8/2qKGhNMpiXJiZnblYwKKFTPEruXqo2gAMcPpxmpY3Klvv
oal5gX0SbzLOQJdwaydRPcQFcRKwyNwetpnjXBhFutpJZdhEN8jNUSjY7cooMMQPF9KlS6ZJbl1J
Zy5OwXYJyztTrnMfQ+JpRhAN3mSI35ieA2WF6flDivOP/RyezTQLuwWgwTlpCRUxkIgmXlYSz5zF
sq4RE+NJIxz7VmgXEfVEdQ41lwMmDF6Eo2+GhEKGIpj7acYcme2aMsfTsV3+miRjDwBecFvrUaIB
kfKlTg/uUU9wCEbuMQG+CmRFYlDM5UXs3jqPoQ/xvWkSMLqMQO98mTyoOSCtd3uTdWhLay148iG8
vq7q50aTh8lkdv5S9aGQBgcsYHdHJh2mIIktg0xljrxGcAXUqxlYG+0q013yysfgz1FXT53TvIi5
icr3RljmRhKEmfvnIE0jIeQY9d+tONxZxyxhNQ957dZSnDpz4FIdLVX3Advj8bdMkOpR1AVTl2VY
6HuD4ptHxGK5iv6avS4wKaKHa98ngDxm0XrLqx+8//YUgC2He2ptlpQ++9kufDAxKuci9ow1RDlP
j8Z+FUUCZIVSm9ssXuJfo0HSl6Dnr257Ruo6J/FN2MlW3Mdm9QiZr0gOAJTP3zuVRrZpjdJdPBy2
quq/pEUvBxZex1izJogFUvCFS5HCPRTCcd+AXxHWLcxe5mWR5KGxm73aqbnjRrvytYzuoHTWfp7Q
ECE2fW4hFm5M6hdA9LiZ60+RwhuMjJLMn8Gh1nSRrxT4y5FSWNcR31nO14X3c5dN14HjB0pjfID1
P8mZFTt/tPYGGVR3/vqfKhti1t7mIZCNHmYI8JtmKFW66lIeugAeo2LrZumh+W0Rw1Rd/Y7Erq8Z
82l1N6zCEIDLYT8LnC+MYUFkYIx+knaNgIGHgCufBt5V7W4zUZu8YR1SdGLMjJACEt8Htmc+3kxY
yAY/Z4RUV8PrNMwtSLcKRtGTgXt9LNGYSzxyndaDvJn24M04gE0v2Ey0P3seSKQ4KLxaj0KrePCP
yB8vQyngOLHx3fL0WDNzrK8UnPG5nl1qZOGxKPi1j4QCv215TiYzpX2/8Ib05XdWXwELG1/58IWf
y1yqExtjhj8wTbTI/fGYXD11O4kpShDTpr8i86Euf831k6IqyzKuICIwkLh1/C3paIHkXQvQrn4a
WvkF4SZgzOiDBOpYwvIv2ErcQBQqlHzmtoMe+zBYOie198MTsZpc8fa61t08O0inAg8jQA7wGQZr
Hgf3r8QS2BdN2plKS2HDtSznBGJNTy+3b2ej5IDa52RryQrSeeWErtYoYyCQ9JvPAFmSref/zyJB
xTtZhiNBO30nZGVKvw1fuWYuxD4NdNMJ/7GTLFfW4SD6zsVnjlL48r51BP02C6WO5VFuMTssSOKz
OzwsXz9qIWj9D0b9/euxCmtGJrXl4gGvMQre8njJA4PPzzEo+e1hT3wCopjlyld55lAT0iwFavkq
lZ8FOFpDk/CbA6ozJ9i/7wNshgNQegQe36/NWKALokZ9d0WqDZXfCn4spvAuguGvT+YhxswYLysV
fWPOshUS42baRylK4OOcwiBr5UguA7wbTxyuikN0OitRQfMdmql2tOmgz7Btt5mYHXxiLc4tfWcN
5eTNrWEB3ZalndQ3c2iU68D2EcZaktAUJ4RPj2us5SCnUccSglROhBaGDzGBo4BERhK7L6xGune8
okJsWZJtVgCubyT+M0Tvo0YtgfLvZyf64hpnwiNn+cygQG5FcWYXObIp33ibFb3/Mqib5x7OJUct
Kmj1QL7Q6FSbNi6gBHg1t4gurleV9F10hyQfS+qD71HmLGRDv5SiOEorsfa0fHGOkdJH6POkEDcM
mxrfjzKchMVeR3BzON0Wcsn7tJt2Vk2nsouWoj8xxsoPGe04f6JihXpAvt3ZyF76XU7uaI5V/lwx
otU5RMs0L1NCp+oNqlNNo3/fHZc0sPTMwcdHudu+C28Gzx1Cf1zQNA6mV9xhTPpNYyOh98S/5Fht
ByV5cfBFyOkFuWciOJWcV0wY4Fd0wMWbGdFN8HLUT+KS6qP3aNo0kjMuU3RZ5TMI7FAGib23A7+0
udDDeNwVnvD8RidfzMwPg28yg37HqfBhrUrODzwxtcyfU0g07uIQpjHo1bkIytyrcBRNIUouVhBT
g/PVMJBFtiuexoGIgXvNCY351x6J9rBPRl1coXtmSfTazytX/he9S/AuqOU0YCUCbEi54+d7MpZw
7VCeRighY/iv+IDK9hqo/rpFSInouOYDVVIEawoW/LIJoIhDuhtvBzuRbAjw9YS73nbnU8mw0O5x
oIU6rg7O7+UPqkBNEJneZDA/QJeXdpPraATyHyAfNC3H1LSv9QwcEd+BoQvPFi2vL007v92+fPfv
e1cybkgnUseB4g3rM/RuCW2YWNDvGXGvS72mYuVfqjNsLka9qcRLqYQ9yTH6tBwkejoWfE4bKusT
W49cnC9iNKpqhXjdZMWPzX1oIiBgubx1CmLjNdmJicUbgyk9+gu9sxk7PBTl+n6AJwZjIc8S5hCP
kF7RDsBd+LAT8dgl/GSscy2B82qJGfks8T6zn8djTP66JAiuDLY1sNu3DW7vub9xTCW+fWKK3v7S
BVbuJzm4TFjqIjqquO43CdJuccVPWUmmbKECfFwkQe/P9ZNQhdFrdMEWg8DT7fBITLLyPMqndoMr
LBToQhjXf+jtH/VNAnPo76XQUT/+NNNYjB278z/KMyE5+9A3WsbfxE1B+8M7YxnOfCB843+lNHjp
I0kTOpDfx93pyt/ps3dHElnvNjwm9rgwErp/tXS7qoPbL8m4+q61Kb+tNV8KlqNB91Xh303iqJ+W
puVVIwK8Nwt4/iG2pSuKp9ZSSOX9Wx2F7d+o4CWE+gXR5gX6jGHbXlfESM5E1VifANJcxsg/18oB
H4vwvT+k7AkRfd67K630qUo9icLxPrmOMGOf4fx/hRBFf9d6X6u1Dgmgrf0jGC2KsAEjvSBlT8sm
bBcknhs1xci3Toc0E9ELlnuPVSptBsseVVTJgyN2/8oPlFhJtThwubQseaqe02bvsKAWg288FGKq
l81u278q+PC+TNCAYbQN7HAdEIKSUKs+GnfkZZo1Yh2oJ28cs/MVtFolwYeQjj8FamIVfp+r04lk
9UTNkBNVBCIATwGcTQrL7IvrPMlOXhYoIO8T7BtBa78gJeFHQXGLlVxmXaKZukOtVjEha4GkQ1Xr
bnSHUk0L7+osjqY+ddyaPYwd+RCqNXT7U4Bp1irjpzJru92b6zNniwzpTqVtWamLWo/eVQnusy03
fXTZTh4xrXMev2WyxFdfe+1NZgSvY5w+u/nLI6WGy9IboT8yJeb+n1JUjH2onxxzmY4Ph87FxnZp
1bTn/tQGz189kloe2ZqZr+GSX5uMJUMpkcqbPijaKoSRnQTY9QrE2TkXyz111JQqTilRwv4qnRlZ
cqlODbcaMlNJehXIFKi8P3Vx1VEvFec5cvtGImnn2I+pEGQCImR17D0rghR9n42cVhR50YxFIeWx
V9ExIg25UtCZgwFDMqXK81rbexZEvsGkT1om/inhdP8eh7YlJrOLnTVajcMid83G3E5Ga4we8kbW
JqW4YjeHI3Pr7h65tiFFz/+1NziT4W/tAA0I56q0kQPRpxg6Otn5jagKRtOeUrt1+e0xe3T6ZlMh
BB8djdLgJftTi/jWnKMbgNJQ9qXpMuqWA0cCSkCd8q70rnbiQhYNAT72/KDi8W36cWUEY5aL43mf
FvX9AZ64iFBkyuaP68PD+AN7IEs4YfMItGk5AJIbB4EBP+k4F51ZdxkFPcy8wGup6GV0dj+oVj3E
V+yByZnkcwRmAd2749uvHW5mQeNZqDAzUk1aPmZfk/HS5WJsC7W227uLTCfr0G8MgL9yYB33RKfI
VmU6h5TgadvKW+jpCefgrYggUmOvYqAB2Zp76YM8JsmF+DQD+KB+0aZrRzOpwyZBGCUnvYlj+bGy
v01wEtRFmxhvuM3QlqNC+JW7W2gDQKEu8Awya2fV9GC2iOJpG9K8wjah5r5bZt3uXFrQx5FfhFnV
gwVftJZ8BQGK55kgy3PEREg5naeTreMUY1RCbR+TwRgOx0k0Tz4tPSCHKZYxiI55hkwTXj/9vde/
yRklrQY4a/zCeSgHXuqbhyoaA5y520p/SvzLK7rsO9HfR4oTAdgu1PLpAoENTSbL4lVt2Uf4h+Pa
qRKaVNGnEHxLePuXq+gRp1mM/lU7q8Fr7s+X8DKcI3on7yh/UnvYN4CxjUOF1fVQLdD7uOsNw0ru
uKDFoPRm6cshfHxT8/EgiOlCXATnOJTkw6rqSLcgW+AYiOdo1QqsEueuo53J3mDqerkm5n4/akKY
DylWswZsUUj92KLdrZuYpEEC9IcQnXV8PBEOWJmzASfzsMBwTB/Pq1O92CxhdpQfLwV2tcCNxcn5
zYYruAuEwl/SqXfxy63rLmTMEjGWaDTbbhwxia/AJ5/pH0PTu2w48kK6EjTD9LU5s25Khz6/6G0E
06/HeiORok6yjlW7FPLm8FM29sUWmkw2TbXdUZffAsC8QjWz0wGHIA6x4f+x0DAGNXbgonpDRA75
TixmZamfV+SPJd9sV/0/M/3VdHIibNqZFilOOWBbfyTQ8rJ89Xyhf8XaXlY3cRHgTAq7rAKv/f3G
yC0p50hVsCLdSL8r27Pqh9JtrzYSjNhuMECQuEXqAi7eJCEpsW/chCouM8Og8ctsEkNZCaIKFS/X
iaagtUqB2kzBHoUHsInuB6+b9Tk95FbFz0mFiK0eEwBXHayr9yCWliK4QIDNhbie5OdW4EdYP2Wu
imGakMFrGshjxSkPs3yhKHZfscztFd/95ggt23iexWj56ucUYNZjjleG2wTJBz6jRrDsOOHrkr6K
Cud/KbgwyfUEcX2v/BS3eZc9mp2VLYREIpTPR6oU4YJeyuGwbJKGNXZRHNJazYu7cwjI8lr5JJrl
X5pQeWDMv4CqvyCDk0ZE/33/U3yjEnnkjTIp2r/PbGWAUXYp2D1WnC4a/Xm0rHaeZ3wUqPtynj2K
mjsJsvy2/Bc5zHpBi7hDHTXHTR8uoeQyicRlvBDliGQ71KQXhoPZzPwc9Ren9YZfRJgIopcEJUtM
2Pk7LE+UJax+BftlPQfkQx5SnhNZqEtSevCyJjBbTXXSyP39CMJAFE9qkVaVDV54DwnSrJgM8CDV
CHMiOcGywKfwIOpvs4HLR9n3DImYF6sxNZYVWIzPQzC+qCF3p8uPV0adZQRFsrmrpVuDk0b/m4d7
ds3+8OJ9YaCOEkulSxJwowQ28Pc+d2/KknCKlQdh29PEnSJuJt6H1zG7hn0j8nRSIQzHmjw7J16Y
Ryz5h0YSt7BJI3cEV63pHsq1niMSgrVGZBGQJPAqzGDEtlarg8nfiETk0Xi4teKQDVRM0ouYIxJ9
HfzfMoNNfA8MHgymcRizxoVNbxd8JpufQmuDJZurbQoduufe4RfIRYYcmwZHHDckmS5oQKBRq6F3
RxFbp4QgyKdN3qc41VissktIIui1LK6EjE4pupMrJqwfG5+XMb2ID2GmfaCvPRBEAfVBbEgJj9Pd
OSRanxCRTU0JVEpzGM851fy3PFu/KZq4Esp7r/sBuJv/JyQvymMS9cUOclgzdBcK6bYLKjLnse9x
TF1OCR5Tqb0enTGQdKEc/emvp+dxxTnjqI3kBoMx7a0faI0LBhUBSkonwTmyDgRdgcn/Q2cN+Om5
Xmz/jRgRk65NQMDm64Mssb0GBkQP7it8DmHzBnRdPN8BoREcCbMqs16LQJmlIyrOtIAkpykB1GTj
MmBWuctEaXnpV/uTr+CwI25QNKVLsP9YkYXfkKikW9s4Iz3XXzxOrHd5ypsQFs1+WoZ8u9Vz5YmI
07Hmqi7OfHxYOTsFsO9CstNUByb16hxbAACiPVxADUskrEtKA0mBtC5IT/Eu8bjvmfB0Mc4FDY9U
YJm/u+C9GvkQtnfw5E9NK3BRIr8X/ilJQ7CUQPvVNYQGQThkogaGmyrKVtWrE3SVzCgzn4N0yylY
pFMPeh2rgS1Gk83PGV5cCbUThJ8CE7n68v3EAh+p5id89Wbl8wcF/zjz4SXtdROMOgP8vshj990K
xNW2gG1UdNe3qIyuny83LeeVt8OUiM24RS0ISZt/a/jUEA2IhArRgv/zal2Ki5XKO5qhV+eLzx1M
5GlWRH112XK93LPMqt5DQFCcOaH82cQGKBqJUSPwCPbdr0WL9rcrTMhfdcm4tvpn6Kseb8eASqkl
GdYPp9+B5/1xj8V1091J1GOXd2gnTZum4ko0Gx4DJTuVoElLirS5j6TLoCpUPugxwsfRJJ/vkT7I
RfxAMHy0c2pRCj1RtHRRuW6EHEt4brGR+eIuzDUL+xc5+G9bMTyTodYG0dnbjIf0PEn4BM9+T4WO
y7DsWgJ5UnpcOKvsCJtC20qHky+MeLundvABxctCVSxqGjVqyAxA8vVEgZDBGQbIjmHFQN/Ehyhr
uW31biNdSv9yUYZYaVfFqvSpYJGLqBaGGm2azhnuES+aft/7/VrRIkaLcM+aNCfsUSFkcgYyIkjl
TaXK27dac9DxNQxP4FIWeI/HV1qj1jdUzd1uE7j5LUMMzqu5AslQQf1JQdlA8kqAzW4aHe9DtX7+
a3Mxq9MwQ9VQMos5f7K/WgjPQiOFQLNsbctFDnBOYmyeiuyCGSyJqgbj7AAVCuC+h06j/Er2WzwN
GJiccGhEOD/4N1qkeB/KGUq+hBaQn0HzEXSpnahBXw5U9j4WcTxga0kDSyotVzd1VOiHPY6l9XZy
WMvMJNmR7oQ1+vovYaR/tK4tC+zRTsK0yjSQ8+PKRCjbmSG/WYa46ZsfQTfhfX6gcbXqmtGYnzyQ
pMm/dCIr3tw4bQBZouXRUYqmS+1HAiC2fBw/MVdiq0KCX+pnbpa8fNkaH7dgN381WXnR3S1hLj6R
edSkKl4UeqQd5d4g8/sfCokdw8FtLKiNFDfhT/NMWnOfz+O/OfGufZTpWUeR+I1/rKANbQsgZkJC
lSMj+kBsRmy4cj75WSrSw8Z7aH17jpYWIyRCNkS9ZKkXI6k8r+bwitdgEao6NfyBXJJOdffXLDIr
BMRXgJVY0zoQk8vd3atwfmnVnlHXJKQqLS7m6MaqmI8PtEJWeQRud2UWE/OuD9z/rU474UE29xc+
0sK54kMt0pIx1fIhMdZbuyGjGYKuR0Aef9mEUTiIBswuiVPWeF0j25zRXdgGVCqhk7ic/SsKSphl
GQh+HI5VelsJEs4o+ahymhDdUsRUV+dCjvKp+86Sx3vl3WsLm+ANH70qDVcC5+SjCUgeu9DwdtbQ
NlergNkXyb3WqjGMSVVFsjSu7eajePJ2nRNLnC9kUXYvxoAPKsjJUCnwOgH2lWS9M0uETW3h4w6N
LjITA4TCguXR8OpjZkZ3EMTVNdl4zdjTCJ2rHQ/TTeS88fYCoVZGxaAeR9eYK1QVlI1Od3hwCt1k
vkaY6Gi5zz7/z5sBoGEfoO1W/Myq8O3gLgXcyO1Vv0/+bQyUaG9d10ikV+vPXjrI0JVVbW8/+Ptv
YvcZa+MJorVBXmcBr8kkbDv51OA8TRmeJyMmlr6zTBNC3777/vvECtLbbtLlXYCzQ2MM7TXvqdoZ
T6ZQKUwD3qEwd6GhBwGFtChbkJYNM3D36iM2z8/KaW6oBB+b5bQQxs6nsLHM//dkg3hqsD53yVyL
TBUiJBqwxS/IVKAuKQKLEtYIXgNjzmPTv57mRg9Q9amxebOBqPN5jFF3ftM9fwNuxjWTHqiW/kY0
KXvowlo+kx7aHsoj2VAFHHi6weM/jinBFrGJnOgGm6+HFjCp3XnjHbZtZVkeeturl/47cm/qLy/h
/CaZD7xMpe/Irl5Ov5oz7gQLAf44/RUZEpmauHvIBvf1e2tgMSx7oty7dt7Syad9uFcNmme/2vvW
PdD7Z7ltSqIp4KjxE2o1/wfcoFUzklkWlv0/ZeEZr3A1fCoHDJiYdRRSBLT2PDf2kSaWzFTz3/TI
JAsdG7sPnhjQXdSmszLM9gquMQDtQDhH7auBPFIPSrPK5nYvmhw2qc3YEGECWMXJnxptG9BBeawz
QD3n4SGnhdG7Vf4mTUpmjZQfV5gxBQMM9zJ3oQ1SMd9Tu9K5O66rRIxqTGZlYjPh5BwoA/DAxeYR
a5gyA0xZTUHqlGTnOyM0ykGWYd+5O2sXLEH6QuhJEhNDz7c2o9AxDlvq8muRhFHG6JEXGa5Oe3je
8qpD3zSrNURKoq/LskYEnETlegqWSe077AYbgIKmVbhXjl4MuCd89F1SR50xDQvxcg6YGkzAyhXa
ABnNeAw/Eonbn/s/CB2hHUuwYSPgcwqa9Hd4GbfVpW9o95mn/HnRDBC7Ys4OmMAKQ3LVlQWksQG4
PtJkbaMETxEh2gHx5Sig4quGS1k6Yn6Y94snfGe1neDkq47IIrtOzII54NoB3OKgIcDMAMzTtbse
jtEeybSaf9epCsi4OL8MpafAi+uXYoyrbCZBIzGUbFnGQkv7HvBmmOWf+S2JI2VILNPg3ALFw4ir
6lbey1IHZ+pXksjj2/Z7WGTbTtpIg3/21iWVWFG0oS8Qo1TLkCOO1GoKdqD71QizBwib9tKm9CDb
erXb5viHY9u5wKe8Lji2uZ85OVFAjxaxc/QTVWUs+Sw0xjQY4lrLeOUUBy/mxQhZGzxyK9tymoZf
jN98yTO9WcUcrnTk2p96V/3TCCudYfFTi3z7SLIG/1AT5mOKQyw7cT32mLaH+5jpP3hoY3MXGB/F
10O9TK8Ayeal9EtyQ4z4tS5JeZVh1dCfZJ/qQ/awSFExagohpQQjFB7P7oOH5V8ItGaecEprzBMl
gxC9ZW7TNt80e4vHLHc1PZnBwimeOwEUxlsSPs6XIVqUQTTK3eeWExxB8Y/yScg6hAlk+iLLupdn
JLjC7pmN1A55IIZqvFlZQpLbyHYVIR4OlAwLI/u5glAxTaNKDhTc0s5Lh6CZVC1VJN0Ip8x2SD7c
Q++kAlD+sAGSYopZlZ+v+Qfr/iGkf59dLNJ8gAeaWZf4IlODrXlrmMU56aRNXPY5QE2LDm0vPYRT
8+LJdzp2U2YEGn62h1l3diJfgqhT6E/pYT2xAOKn4hIN42I1cHNgvJumslRCRB2clecIePNHqqnV
5ScoTr2lkajj0DMYxVPBheZYZo1mzGIBCbme2s5nGTLfzuzVz5bXz/oDyn7EWLE8gLgqFKLQOGIl
LUYl3ENFwtYco/uJtuky2jKwn1VsHnGr7guH4utS+iUA4Z9eHLtjcd4016HsH3vGs4l74BRWQOV6
IuuTeqMimZs9itvXmObySjEgc69UK2F1fVh9X7OtAckOA+lubNEV8N/P2rl2Gyuo4i2Tltdxi6uS
ewX6KO/FZFj1oCt+bMrgjGyqTYGmExW2ztL1VSWMeFxT69hG1xqL2qyF+ozooUF+8QqQZoe6R70O
/JJjGmAj5kM0G2S73zXL7/9zzVvbh7KMBHD4gMziFuIytWNoWQkQqbBH0+3jXA9p1EEFfjiHdRn4
SolyqRiP8NKUUvHDX0DNRHAENNgODucqZbScapY3SmPUfc7B/xMfUkxP+u5+Q5FJNkptGbq3aOvT
v3r5LYujtpSjx6Uvn8WeFM/5zaowSMmRVpuQ4KIyuxxZkWjHuRFy9lm/BCMv7ezqNNDePKbGatGh
PIlshFUX7zkpLIjtkd7YInbK/d5Hb9foQUo5y3JGB+hEP2n6JuB6Drie3WsQUI0aI21vsfMkhQvl
ofGvEpf3zxtYsT1I/UYjZkocKrb+zGyJuUECsSGkQiJUGYh6BRZreLs1LRZMXOnJOdiN5oM/pS6x
N4f23v986VIniTTT7cRjYggGgU5CedktRfKxpKaUzplCOhjAK3KenxBmpgA94EE1T/xawrAQBkKD
94MQNJClshvuEPHqcunktnGPqYLGy0pYre4Kqu3KbvPmesUWFmDO3Lyvt8s/UqHyfgW9UKHpRlCq
T91K9NGH33PRRkm36Y3PYQ/MDxJmTZsvlQ6vB/FQCd56XRtRiGyWkyrl4laogw0A1PTMW6Tzsjx+
ZVvDisswU7qDKWRXAyoG0im+5B/HfV7ziPOEQH0WZ1bPOd39gBdBsky0n4FBrvWw4OB8ueRM1AFI
imBIvhftzcOBEGyoZsl6hymVtLtfKVi4EsBVzSMQBYgAbYvgeva9mFdPjGsdcYGpY+Liwai1Gavb
MdyM//5RS1FPFAmAork24zW3efxVSwaokU3jIsO2o9E+Z2NjW9r5p5BJujybWLB7DNEg2R3BaoWu
RFRNqPdHr/V8F3Fq0cgU2w59NiGxrGaxHLqigpryv3EybYhCLV+3o45tHZlAWVfxXjZbntdwNFAO
bQe1emOWjPRv70Lp8iwJK7sYsF3xJfb4V9caew+K3uRTERY6R1z6hpI71Ffk+qT11Eae0SN7isow
yx0vn8m9KyaApoZZ6hKc/lkRdoKtKoEyaC4wdrLO9nendWHQK0N9x4wrTtI+3YeNh57e+D4bFqfp
0ttxq7r10QXV5mC1CrYS0F0y7vqHlXV8QswJFeTyb4WgsrpyTfl/kyYis4evEaYzEfvJlbxejdvk
N5kQBSna+7u4TpuzTv1XQ44It42kclO6e1KgACVNdGfrYQq5auDn4RfkeR12MradSwP01gwWAch4
dxHJVuOeQ2gneaXM0xjDMCUw+rSVCzTna7IEfqv9SSmtoRVvhlE/p32QxaGvRL79a2nM1dDPnr/g
mJeq2+/pJTzg9T66BJq17vQrKoHLigyAZ0yPDyVq0tgFFhygEWBawyuUADWIuTk2OFKV8QVHdWah
O53IFQ+heFDJ/+StqsYoHxFRogm2tbnRDmhjmfvUg9+Tf6jEsUK6gWQwNp/bL65MSOx6hUH2Uzw6
+S6+LeK1DnOA8CK99+N7AbRxQOy9EjMuoVL41pJQvbpTHVsZFUjDWWAhBWTfaa5zNzQOVbXrls4z
O9BsKXLUmSxWF+M4/5xuBvew+7MgR6aVIdzpvsHSmSliLy/CIsFCtXMysqWqSAOX7ktL6rRc+NvT
FJnqsQeMHTKt1fbSsvrs/S5sfu+rw2wCum6zCuKVVYHoaeZRLuG9JX5apae5Xxee/FVmtZBErVSm
7ZB+ZcizVp2liSQ05HOu/iC3MYn9LznKNzgCHLntK9xJRmUXi3NipkxpCQurHpEhkWVTGkxP+bwb
+3afnrGTjIq6T7Mn+vkwPALm5pVWaVCsJp3ZH+EEW5zs4P1Kurcr36qhrnehzCGaBTGSBwZgv3Xi
F3PhE8A0LezKyjCR8v0jQEv4gyqNy/QUid98puaxazbZIem8W/7DC3g66vCHrj9MQxPOqiEGbigN
RO6PDZPES21lEMRxrFR0IJuSbYL8/ZHtD36sMO612cnicfikTOkWkHmB4Wz3EBjDUSFbKgllxpTe
Tc+uunOAEGJdyoaWxTLH0/9lYyrwo3OQGN2WKF80ycW2bqmxWa15JW3dhsVoivAYK+Ic3P/6ep7v
k58PVkUAEf7NfC81diXi7s14SPm0Lq5jgISgT8eC3Q12bfFJwF92S3AbtYadYrRxqTR1hB4egK1Q
dZvI+qDD7JTdfSuoADLbp42iJMbay2vKmEI1UaYkE8QDDVI5OFT8mjLLgeP3470ZluUgpKgyx7nE
UVbjIUGKewWPHQYnN6KcrX1HeeKtSFAkwR/X0GhbVy+hgAHaQFyA/r7UC1+heZ98sV4lDxnnRUGz
VSJiQ2EfYTS80ZOF9HJOYWyI/wtItpjrDNYn9Nxxd1Dp+viYyUc0rPNl8+Bi6bkq7h7lgkRHYqem
PufGwsdVjdOENBgJKAygb1z3EoK23Ibhf/KZgDwueXAZoeA4OFxd06RsUcymyM7sQlV3/KBussam
K0FuAW1EOj4Vrng+7e4+NxR1IRkVb+wV8rHawrEQ6PymnYpW6X3bSF9R4tznPohyvzuqQrxpd6u0
OHkrf/k7SStpAuz24bzUfZn9AQApFG+Cr048Pcea26uPclWE87fwfoL/pP7UbgvhQQt8u6TxVx8J
/62yAxFkQDHBhIsExmCpYr8XqM9rpNNWP6OhRMjB1WuvK2wNtX84xWh9/MZ7kx5Bk4HRkHX8nEM5
rUq4Ub+vawFW5WqdwDd92LtU656JRbIeswXmHpPAOVP/+WFYwWT/eKa+aK88WWnn2FGUtqOB4JU4
n8JGjDeUhGhVB00Ir/UfWKTfzY75OUDeoJWm9dplB2KaX4TwRoTJ5u2b5bxMf+1C6MzOvw5tTrvn
yxBgEaYb27gO2M/vGqgS/IooboauvpWkF6IKVWcQig//1bMauArx2B+IqarBCRfAjauRAZXkU910
JRDk/IACN1t5jgAOsJe7IbNog6grOvsBA97sv2JUNARxs4BIOmUrs1XGSY6P/8DCYlRqboWje+j6
nz/tAEz58NsK+6i3LwYNqw4FDLyMpeK4p8y+daWnvrU6Gu/hsAhzsZQ0yyWeL8upWsmd1Tnh0xvT
3b7KalqjM0GX1CbUdP2t1rGolwha6KYzamx1hO8UMyaVEtQ+ld/2R23s+0qvFgwuRaIL5vSrYXyl
dywCN3z/0hozK4DNH7pEhGiD9MFZkN7Uy6SNXuT2Ir4UeYlCg18RedO+L+EgfEBh/T4QmFsgJ9rq
YzAW/VpnWEnL5eM1Tmk6m7fkg+iu7lJIDtr8jVpq8UrrKry/Pb98m3MTiWwQ3dRyNMtcH7G4Q3L4
JRTXYG6XiQ9swYjOmtasenhzBgrsQeU5w2eyTNC2+BuYMWj6k+bpmNKlQI2SsAZSRmUe26ohr5y9
We5wN7opVUQK92DOsftc7t7JSrdVrYx2MxoZQT8G+ldDOVAmxZpOSfFyxndkELbCWBVXNRQRxJg4
fUdemUa3M2uKNKAtgi8vYnwPwQnGOmB5W5Q+xhJR1Y7LfwF7B6N+z8HKkhdGa1Er3c3ai8Uwfnhn
jPDOMdKUvhRIzu4pKkHo9OW7mg4WnB9AeG5FqWGjdE4rR7VPdDJuQ8UGbKy2dPDYzYo3blKPPPFi
oHTihkSAaTHmgryYgZQnLodTezICHAfBDZ6h3eOEppcChD2fucS0lVeZLUOlH2MMJACwLB0YRcci
SCS816b7II1qEDNZfhli/TKwdItJQHaigvJlZ6j7cL2jxFJNIfxGRwJnk5L11PxGY+RnAYw5nrbD
aEfJY4xKKOFb1TLZAVzjXbX1wElBe8ZTCkwh1U/KHnPRScncbvE5oUrIQtDgbZkIC/VlxwH//+EH
AtS7orwtAnRJGWvGXWzo2Uuo9DgLsxo6Ct+kQFQ81DemX8zzRSyBADvRga0QollquLrnIVBODirW
NXVe3H4q7CzjMCWVjfnOD7Im/Qnt/goDKEDTnQ479ZCCn4OF2Vi2ktx1b0lM1mFOkSIz/EDbwjMX
DJrw057cDWBlPdUzObQUcs+mt1toJXC5mNh64mSoABJLJYOVIPkPDaOBUVGwHmaYUv9MuhTPt+Ch
4B6Ne1q8illQ61mGGWp6h3FS9P2vXL9FP7OQ6rmYB5WnvIAYQS62/i6VP13odqYtCEl7Gr8mx1Xi
5a7SX0UdbzuWmn1ls56KiER/TJ1xHlYZMPvaDKPJKC0H3/vsK0B8CD+FZYf1FFBlh8qK4/4GEdD0
nGvcnTX3LNYlq9tiwjuCV2AoshpXcLG0Q1aSqY+MYrH1PFNEVSIa2k4QmIWEgFsbnRxHl+4l78Mq
NoMNMoq3cL/3A0GeY6wLIM6ESrRWdy2yGxsL9Rsholfhj2NFrR0P+Vvy16p1mYYmNrGpvLy4QUnF
yWbXaCbf1WTBT6jckmsE0csE0zNJjs14gdZ8fq5q+aKrIIR044N75CXOp2MmOlvRzoaYVKYDFlMT
fmWNzcAafQl5lbsRe24Wi50k+UuJfQr9hU05aLsDZJnKqFAhu7NwMYs8VDGButxYOVaFr92Rv6UQ
BDg5qaZxVYSKC9781ZdJtWXxm4y/t/F7K2dlcR7mZbUvsKh3K1RjqWZ0gAXZLkrQzE2L8ALQsu5L
FWeUTwoK1gpu0IyXwqF5oKcMiuhIX2wcbmx0p38JbnzN/IzEJt4ws4ldOv+XU4SBlrf+yovUWozR
3bUPHOLtMa98c4Dguch2STs9bPaRGl9txIfCplaJhb8FAtyCyq1AvNkuzu92/LFmiQft3xygBcfF
j7RqpA0lpS5NrXJGbE7YC8nJnlPlbL40eWWG8mGbB2o2uEypvoTV4rtMJXO48lvl4RqLIw/axzAX
X/izMzN3aAWp3fe+AkyQTun1oSgM4pNxRuENDkudqKGVuWdaa2uao8mIMD0N1SeqaTF999mryfcG
DOuAAiy9tl4NY2rVS7pm6P92mjM8rb67P7IcNGW0SAypUQ+nJS6sLltJ82j5tR5czwYYmKKKw1/7
jOFBhSHRJj4GlIRrYYPcBSyyT/RMDTUDIkIpDHPfYDpgP2yarzZwnjbTpFDuk94VE18xdEl0a0j1
i2DPvXk7GWgZW9kIpLn5mOnqffCH4AmAF1v0Da/deRqfny+Ng4Wnk07QSl+bfz15CCV+udp6OmbE
M9qjcArcXMrdk58XO1ntbW4PdRoO+yY92LDDRlOyUVmtBmuPvrpTxNPOP81FyHGqrJBbt3vxPFg8
bbFdT5yQmIHILeXe7EpKO2l/ZZ1STxRXK2P4p4mOkFnz+s7ykVZxPEjLt6qzdrZcMRuwAv1cEeAD
gxgt1y91tJtNnVIEX/16gyPXHMxKhGofPKGgB4P0KdGJ550EJbBhAn56ae250nn+TK8OLJ44C2pH
6h3wU0a9C7mVp2iWVj1779WixBBHtNfFXPOvvh0KMGphgGQCSd8gYOhLQLAZE9lCsjoiNyY5tKr0
j5fKaCtVB/8fhQNJ77oxgaNAHPbYR0QXnizMsSVGkkeqJrf6VjC24MdyLi+W294Kab7Vz8d8S5Nm
DHckTYQfG3vuMKYXiVekYoc6xct+ml9Tua+/BXHv25advpwhbHvWXH4Ot2eiQWY6UAi+4GJdBYdQ
Giojt9Yj9XEUPPiePJnfX8w1/iTZdxi5WE8/ST3/b78DkdfoONi+4d8eh8tMRBeou9ZfppBncm8q
qjPouMGkvmVCz3+x6b4tPRoeetSaZ+QRfV2VPOR6GfT87YyCXiqnFo9QYt+f50PNrj8e3Nde7yAY
I/KOcjhNGn0A90sqWm/9UjOJXcNWW//p6cjdardoOVhJczTakxLaUd9Jt17chYl0pjGiSf7VjfVW
pg6x0oi21C5cbAk92NzVCz4Juj7hhaH2B+URKX7B3X6kQtbs4AZjr5WGEAMThZQz4Q5/F5CcDc1E
nDKt6Bd6ocJktl4+5r49ih7B7ZU4yfny5PjsZlrqy+LJwCUuiVOfDtXl0r3DYNf1f+p1LMfPuopy
9qYkFxiGTVu3VDPQbTwkjxnKeiCB6y/sEMaunCcZJhCIy+vq1WoToKknUU8tXGEvtQaJpG9ciPdu
Quux5lysTXSjnCtTYljnN/ewEvko2FiB3ZHgtJqb2WGvjMBcy/iOPmW7absNAbPB/hCFFzkGIUyC
8oQN6KHHFTnYwJgOs+5GvENxscLa9TncAQW61eBOm5SDqHqSv15giOC/zkKtK0ul7fLzxg5luntP
GMePvPwrqTVO5zW5Db1/LV9ObhzleHI6CaVdxNqWk0MgLHxJusti+F+O6M87qucGKBPXyW13jH0U
4Xbe0UFqtP9srMr+EVCD6RMCgM8mXDJszWIyFksu3DEgRXXLiQ/ab10pSxEjRXwwwWmxBC11qtP2
Wj5n6b9jadW3OYsVtqnwPUpQi2Wea2Rj2X55TCvGjeXNsT3VcYq9ilR+83IgRViKgWN/MSSXEC4L
eozlwaac2dhZKBf2Jr+e81eh/Lybb54hNSKTj0Mz412HTb28xBA1s55v+FRaRjYoG8ZKvhiUhMQA
YND96XKgIPHdwXTjfxzVCHt6j9N2l2z2vpeAQsgaUWAfPidd2owTatNAWr1/BJd4/1gjcDb/upkP
PEJ+zptolgWnFpdSQ/1JGcqf60+n4zKkoidfEzJv4SOCaQpmBbmv1GkKf1jBrGNd0mJ4gVrI5vR4
PPl9kGn5e9RIb8k9tUMK0OldlxYKYpW4eHB5+Xohetsb44u1RaOVG4fjlfxYcaVsjhVev8RAmW8C
RAjEwSLR030wIFkIAR1nZs1W2rPaJXTdPV3eWtWtGEQAX8EtjFxzhU/JrF1pB3qh9txT2SW0GnGU
BIHnpq3VDNUfeoULxRDYjIzMMk9uAT3ZGX9U9QI8M1dkaRd2Uvzd3tB6B5rjUD8xyOWKVsZRKUAA
SPxznyPX63y+e8k+tyM9tlF7PdJkLb2xlNbMfjkxFGCjWwC8Re41/rV9sIaFBUPi5V2aNec/njWE
Oo/18TEm8Qn2YUZDWp4rQauz37QfvoTIU1Iy0/KD0Lcud1WmMst32drb1G128/2RYUWCeRJbcFLi
bsyou39OIrUNIYhl9ajPMvUE+pBEJD26NqUGq4Ffi1hzSkED7KgVWiGL8KiJbzKY0WH8V8sdUd2I
9PstmkApowA/1CogucrqjZsAs4Xgnml6aU8vYZCIYVL3PS1TFM3j1OJzRED4XADj30ZEGyYwKWB0
0XDIZcmUuQcilO2ZOYqKzvu1/zWMhwlXQl37ODdyPv5o1L9h5P6BbBDfaWR6L6eg2ivUd/yjkC4B
PFUuYsVViO7rzIdk+r/Pf3Pfrln1ayMC8+9HXwrPBBTtHBVZOg3Bd9skkjHNIyNRxcRUnPWP+NMG
RUHNoUalxvuUqHvytNNXNJATKSLxXPm+c8iQn7N6Ea1Az8FWCqCM6pzsdw2ObgHMAYtpRDQP6lUR
MXm7A3XsSH8a2IixLGKTAyAf1t9JGXTowIegU406Y7+hQ4fVG2hP3dQHvIfCE2Szm6b8GfaJDSZM
WBqWYtuIjzxzvvlKFmXxHjrMMgvFgqKktUC7mmFaLqobfyL+eRnI+58ldOXp1KPbtiE7qYizKSjF
a+xNbNl9+5wtPayiU7NsiwGOACUGus33R+Tm3ACawviWT3oaBNiyZAYpqoBffldE+Xii4kwNSoMW
wUZOEMqrD7aMj7KttW2KJvgJcrXDgdt2K6l5bAIEQdClMfb+3SYJ5lRHqn4UZ3a8y68ZMxJFyiQD
KsFOwwtGen3SdgkcO5h9NsOfiSs3oln+Fu65LmwHSJGDpCbAzxxET9Qm+kPzBTocn/dHSgfotHAz
0PXP8oyUOIJAHNufDOS5mqqxxgGqJBueBNw9iuX5hrHvXPVGdoxA9Vm9c28FaA5yYMPXD/KXydn+
GBwllWFM8JOxRybzw3gAL/w+qnSC9nZlZEnZoTlEbXHzv3gpAWgIdiA5AbxGpWq7zvNY9j5njFwE
wCs7doyeVHq93S9deuHDAEMeiw63eQlKIt9PXMlbljaokRmc44sozOI2thybHeidM7vLZNkRBppj
QD2HZYJSUXyjSlx0p2xtvPqCKN/7Pn4dksPJ6jzVyFffMF/+tGfbde5QEFsBtTzopolr3wm96g/p
QsuqtlfXupjFIZWw0oQ7C54pEHQPt1blop6FHcPgzQfMw2lonR+slHhIIs9kVlA2tnNF5jRhuj4p
AN565F2DDiV04JPAKy81dUdY0SR/0dJRgVBpPP2uAS+0C3z6ozVYJOZFI1ORS+X24IA5YflJbHff
Ktgklsitfop3+uNS5kE0GoWwLiAdahfXW8G8Xc57+jv4sx/Plqo3AgFPpLx5i7oTJWzbY38ptn6S
3fjoI4cPfSI81bT35iZoKIcuvvv/2i8SDfdPnwSS3xhw826nxF0O9+7UNY+eDefT3EtyM/NE/amw
3EBvB2vaOGxa7D9RFHgmHI3eKsD4F09Dc61qI15zdduW+YcGLS5uHqrQVS1mfU2QN4k/bmVHLjEH
2HCUPJ3kFox6r3p2oyWYqoY4qI/Pf/4rMy8eYxu4s2ODAFBB27v1DSCYNxB4SFeGGB4GbkTvoVxX
Dm1/5/GPMKI9sWYZ/y2v6hTxr2C5F+b1Qvg0OPkVASZHMakLHQnta3D76lDKMYl/bGCYZgBqqB4C
P2txX/qn9m4PRfWzc9hM3LJSPC8eURaGNJlIRzhL3Qc0DSSVV/J1+Jssjd+6yEhHVtLupPCkknBC
OuktruneS5HlXg00amlJ+OgyB3vkw+dzXDTuTiRdzxGC7dVDTpHFeqzvhJL3+zpMSeCdwxTQz+yi
LhUHziuDiZZ3lzB2UHZlaLO7tbNUdSVpfYwsN3rrfXQap/gCf6UGS8naYYLyU+NAbHFUOLvJyhp7
XQMfx72s1uOFt6izRLSufH8HH8ImJ/LGrPpxGT6jWSMyP9G/QSUXo9Vqehlb1GBH7NhvVmk6THJp
xwyQTeB75rNMLh4n87QtT7DYediP5jBPXu1jBO3Xq90dQOtPtQtX1qbhPxObf7LXH7UvVyEklPbE
bcjxuOlim6ODyx8f7ft2XtWrOYumsi+2gWbEyMtWnP/gDoRVVtU0dptim3QDEhGmDVnIUFG450qq
Ev0HAYaiIHk5EBsPFecF4r2yRi8lc7LVzrhVj0qJD5JWwDW4EPw12sfUMU3XY227hdwzKxBO96aw
4/cqJMrXsS1xXGQe+ooWdEm3sbIfjeV+a+GuaxqD81U4cejxaWiRy6LCSd6yqGSf+iR9an8Lbsby
2bVkFRXVfW+V0k1b8S8H5pN1oFquX23c3q9VWfjAVLFHEpQLb17K3ztx9nVPc1Drjofsavcanbec
lXrEFaQ4fXy0nK0C5yadJVH9ontfXI8y6EFQu3dNJWLf0s6EdwdxMwFoQ+gsjtwkh3o5xtXfSAAJ
LkRhOgUew14DRag8tU/ubB80t5aQhJVWH1L3McbTFdgKhzaElVsm29dcHXoOi7mUlC4VWTdXHvsk
4xlPtPIKAWFAWsFp+dfZddPxfNAfMH+xmnonLwv0X6ZSOnUpxR27ugbx8aPmdIjWHZtrBAxhGRww
m2omWvsSpbjT/A0IvbrTz6v0ES0ZmykWUka9NkMAr1APvyKU5N1a8GY+pK12Hu+/dMFB1Pxy8Gzo
qWxEkI8inRvCQxdlU53/eh1pb/NpKOZt4/4LRihPo8nMI+3ziurhtMIYvaoTAjV9dODeH4IGrC03
kNOLNTu1eYBe3M69fTw1FbA9PdUYTVZSYtCk4d19SmIYC8xmELeWjWXokBxgPGEg/055Nz/R98Ah
Ho+pqr9d2Aypws623BTOaOq4uv59cdfQnw3VZOZhXWtcdOWTl8lYC19VCYgMGonbrciYN4yOtoY4
1anbXfvX8x9RJnErfKr+1usjHyRVknCovUrPn878rT361uBWKI7KN4M4vg0bPTGg4svhuquagVi7
j53nlMxiTTW9F3pwG1zePcWUeCAG5nKE6qYmG09/m1vmXC11nV2bVDLS03VakjvIjJVNOzZOhWis
b5As8ncCBIg/aCPwprmn2d08tQ1ZLss5OwrCSloz1KWk+PfdKr6HyTrQtdZGorNh4ZhN2WMyrs0f
4j1CKGHxJVpdH1J7LJ6RXVzupdiCFdCfs+986mCfv8W8Dn1qookVfrYpk54k7VPjh/rlbezD52+I
vOoZxViYu9b+dqGa/MzmJDMBX/oNyzn3XlLel45HVFLUOIOw6g9bsdayRwtVGvk/OeBiqwJA7j0e
hHUTw8YE/0P4pWAjsU5XOxM2g4tBHZRLgueOxeXaPu4S5Qr78Ocg9Y5swNnnDawvR/mCQEpWjQNY
Egylq+Fr8PC5CDz/05ZpGWF2FStG/sjTlNi+K3beQfjZEW3ep1FLJNzat51vkF4klO/fMQyl1rBs
viR4iHvB3cfrYTn4/M/3SrBsGSEqlMDXLWf4MN7OjfOTFi/JJExrOPNsS97d+iTkiRqVjjULT5BQ
AmEq6IrCQ6nWke43qsPmyk3SWOpXnrPsigfIXXeCgcOX1gA2vCT3vTcXKny76obDcSpepOsdcwrB
cgw4qo1BnG9pqumhoOSw7FIsOEI5LGqJNKf+1qB6tBPTlNieLcgFqpAsNr4tD7J4SXBwfy5h+V0D
yReAl+/n4EcvBPgpnMQgyouw0cCfcE1clfAUkPyvp15iOcpee67o3mhkl5aNX2snR0jNRd5okoOG
FafnbAkuTTtJRhJZFFBBTTMjpWnevs1GdA5oFsI+a0bm7lLOanNDDwOwrXZJUbhfJRTP1fvEqxZU
nFpAXAjL54tbwkzBRtMxT3cqRrZ3c4+fUTZNbYZT4wM0dnN9Q5v8f/JjRX0aQm0Ez9WR20o+R8y5
2zgTsLcx7/1FTjcfKJMKR3dfQ1MrfyPZ1mRtgP3+fb+7zj+MKkUDe+MMomGwwRhUYHuUllGd5CdF
KJPHQ705WIJapbgEzkNurxAUDpiOTmkV685K+kosPo7LbamLTeqRAoyxDTqcU2UnCEywB2F1R8Zd
q0qzophl/jDSJk24GYjmilfU8YhDXFO/5tgPaidtEl1pkGBiI7uscSLHlpxbBObOesR7YOW8u09a
7Ti0Xd1/1RnuD4LT4cgdKgNhcDDgkIpkyPj4fpjbTEyJ+DEnw1sxraIKhdG2yX7a/u5meaj5egj0
gAXdO9LdAhKD+7nzcE3mt1ZMCoCJ+YjnwXTnCJCai7EPiAiKSSZ/vKczFB0DDgrV4dm4CFYs0waS
tjA7edYWaNUi+WOygk4fxIsCaHsXQnoM4IM+Y6ByoysgeHN9SzPxxFVmh/Z9u74aXXldM6MAGyWR
Kci5PBb8oDtcf2cvEZD3W/uVI+alDDgAFqaVK2JYQf/LX6URusxw0Z1bp/9Uj2+D21xs4BkNUy/6
2ElghDuvChR6dGJfQjYRMtii4EJggFVnsujFSPo+ZxNtoHFx+g0rHPv3edlTGfvhBfapMHzOdbOG
Ay4fjnrMNQ1M33+u1K/fZh1REJDp53mYCu7t0OXReD9DW3sDD9QwWzTO6+sLqgPJsCrS3W/pWPAx
+qqnJaKVVL1ItJx9jiRvVH1aLUsKMLXKHTINLMhXfm/Klyuz3CMACxRTiMrU6y9BCiMKlXHPiJ3S
4z6MqZ0Hg7TTDCdJjtyMuIyn6ykJVdrlWxN1wugtvtIpdUoh7g6u1dI4G2AAWoa3cgt+wvkU8G3O
/EfX77j/qegsq95586r1NLbu8S+0IIuuaLTVyD20tlg4ZwFwYch8L1TbnUdVHL5mWeo2Qk9rVwSr
TGrt16Y42MzxUN1w8HLm69M5BdiDXEPgaOqMGjrB84V8VvA7MFqrVxoOJNLuuSBZwVI82SV9lxUg
lbnp5WQZLuIUCwU5Yo22MM1ieW+JqpUDMYJdYEHe+EHapZUmTrxSwgqK/tsjdF9ZLqfUBiw/xY+n
wHuVWmh0xoY/BoIlA9AjRUHFbhCkTC2FkoLil10An5VfLhWDaUuGYoXLW6aKYqU0Rcr1Kam2p9tg
HBdQAuAGiknQqYdC8MNmAvCLMraUPypzfCUdaHEc//IwcyPhmC8f6EzAbVrKC/ZiXY8JvMoQyBks
KBovzzoOTIuyunqPq1Hz2QK3sr/uEdI2WkoHHsD0C6XUDqvq8AbswfQ8rUP+Eta4goJtKhN2VKht
kpHAENI6SLurkEfbxhXt6GsVXTqrn0xnMI1qj1YTH/6iMJIrEET3Vhh4VR+KUfiisWsY7DEC12Ku
RNSVdIxpHW4xintRefEUAFE9X8NI9xyx40O6uivo85Z2JdwVMnzZjDXCzv6SmJpBPD+c9+7hIs/7
ezxcDx7DhRWqwrxAurFT6MDV4XEDBKpjDwsFhLWVhJaxcJSMNUtY+zAppxro38PZqT3z31Wptbla
dDSivZ0YOdFo/IJPp2F7fv/3gjbV7VuShCUHFgmAsv7BaZZ5sm5jfujWGTzgDKVjFwQAiBi/WPk2
utjFbxWZ2qKXMVqJfr2vVBszVVZTPQE/tkuvVIUv+v2KaofN3H0IwI9B136nejfYVhcKRq4kZ2Sh
sAW753jV6KwecO/HMV1KacBlW0hnWaBl2WWEwkQqoLmGockOyZ32O4QG3GQy3PpdBZMvyD7t6G5X
XXz/D+Ws9KNoI6WFx8yBd37Q+lScXxYgeEKKczXU9ArQ5KMDdTDvrOCm2PvwoPmOF3D5654eqW99
dx4jo4RTIej0PgmCj6roJffwP31s/VNo2zfwgnk41hp7HCR6Q+gzn+EbrhCXTxC0WvgqCTHE1pIO
YuJxGkDcjypvR54KwKsPCtWUdHOagCJCEkhncRAEGTc1c7nrzZWZ5rKT1YnlmXyENAsZLfzi/ReV
nWjx/5wfS0JPH1XwZUcLR187G8xjZC/GCv+H+/ieQZ50StfhfgOA7rWR31UutgnBsXusFZ5CHjfL
C6Yy0jbBqA5UWMc3W+qhM3u+stvkS2z/ImY6U9EZXdwy/SG8Z0oRRf07CtKucivdxaSsO7bl41ma
ryR6NJxoR9wdYkj46nYvudIqkar+sR6xDlMoYbvx7m7YuKERXapWLGNACIseWlmHVCJlWD03qFgB
lfKUXohu/BGDF5zrlZecnUoCB0bJlotl0ObBWXv9rMyroIRgcdJLfJ7I+DbAiRBBAR9YsrgcBfJq
B5of4hqqU1p8OeHShfGx1hdu5l7l9AvMic97nEG3RAVWvnVRVxPK6pfbhbZHY2Gk9/8aNRJi7HBU
bFDSJKRv5BHsNNkQbschFmajbamHKj7UgqjnJNGyGi1eJvlKGO1JAf+uKNEm6fFbxZyakZroiMuE
XawzLJEeUmY8uktXDoBsYrksj0///P7HMLDoAFDfL3D8GrunI8Lbb5ysg6W4kB7j2mn2hD/O0WwC
9laxFpK51vIDhKZqHYJw/qVrY0A8Sq2Itd07sZ7mzKv045T0zwwS8mWyZwZibV+K5OPlAsnCh3zP
w87Afnh2XY8P0q6zKuz7EQsg5HIFP2yfSz8E5Li4tDavwoYuDfP0BrvAl0Mc/5XFm4aVub/NxcWs
sUxZ4FYO5jszy6+KFFU4P4TAWX9XCEvtK+rHl47Prj2wPvzy7L+KqcJAM+ap2rmTWqT6mWl1l+mc
kUIAK0XQ0RjlKYZB2B7yjrZpVmfbnHJX6jXBlsHibBmw6DpTKFZCqGcn2uraqepYHUDbaS6Db8fW
5tTkWVvHdr+HzUXOZV2rye9titVBNvkCjFBXq1z+ly1KAR3ACI8RtpvK5qQToYMVLUvBZC6+6DbM
OQgs+bnjaNISbOhG3euN0V4zpJw+Hx8FdwACrq3DBSvy4zgID7kZvkLeoKf2R0sYQy0LGNIWK/Ab
YsXIvHi1ScNRBJuitwwrJR4MruF7rKj+StB4Kh3RAL4J6qVLcpaV7KwfwmcuHVCGIT0bxBvhpLK0
fR+f2mRghmndPiRmZORrz+t6qJUgz+/Dwav1RzB9XRq2x9NrdvRDBCfBE7lhsksoScij6FPMoI0v
hYUQNlo06i67CKBheNf3JEn47DHwvuz9cXafpkmPSW6pEuKKpo1da/paWtF4V4GZyM6UyXLJWXC6
VKHTQQnge4CU62RLY3mboFhAzOnR+VdY+tloJUE8pwOT5ylHV/TVJxWpBkDDBeK7AFrZT+J3LA0R
b6Y9J9xEVmxao9j3wWBKdZkd3JinbRKoC8SL5zTlwXHdqpue+FZCozEsKkUxJ3Sb0is0+51FvcN/
d124MudpZ4QnUivGWVCr1cuIauOf1xdN+dEBYSSpRHzZY68JL3mmebzZ0o/TnYdSQ5QkJm3JxyiH
Cv/CV6uLUZn+om8z/9ZmLXocZAkTlSiK51jtN//l1sBUTkeVMNxquUL7VTWjG+AUXDZ92IUxP550
IoNNc9l7l5A1ESFsatzEDehE8CH9shAWn2NeeAJD6VcM4frlnPISgydd4wUuWF8z641H4aG02CM2
nHLG8E1thiLX07WkqAQj5XrwxtGhevUT0DK1K1w+/1fBjnooJzD8Iv98+ng/AhK3ppK1gYZjgXbp
PAGtajHU2Sl3+TCDeyzT64Xi89kM2lR42FcJZsd18NAXAj0zWP7m7064zXmiO9Vmkj4jHEhVp1Zz
8e75Ywb3OEyOP1PZpUK+7saRq5/B0rDveIrcMIaehpevQqFByj6sYOhZccFRIDxZtCjAUUTZ3UHl
/jkxz/iglQFQNxD3pWjrtdQcrVnS62w6ITk/qENbtrhHy4ry669zKUwkReBDBK2cuGXoxWmhrAY9
Z2foVLnHleqPwJS9Peucq6NKeMwdMK4J3o9zKD2OtGpOf1oI/SlsWAALBBy27qwsOY0BE6UIxgbG
uoGUZLcLXMMVBJcDHnVOYXY6jiwMt7dHaU46A+/lQBuHqenrGv/BkkXckrvNGT5n4tXGY0fzZv+7
6ktdH/eJgENgsKdweYBGyDjHqF3s8nsOMolHlXBkBqcPZAH/leWLZ45jzuGMugdbQtbxWWl6nmS+
7SRqW2fylATEEW9UasWEIvw3BnuDhsWs8/WXe+gRdn/ocAj8LTJse7XdIlqZJMg801LnyyrKXbq9
+VOPdmnz5Q/ZwKLMOu7/wXdwu3d73Vw123nIxQopRt0++bVM4GcmwuvLY1bhxbbezJk9xExcDwA+
I5ugCdP9AaAqXeHfGzKGSlBzo8gQgMdyho5rzNf0InrrXI16BGtXuQU5ghlOe7WmIIYfiVREN2jr
PAW6A7m1Lb5Co1b0rf3WXgLZyly9p2qwjOHdnm0GaGL2wQUteEkC9B6JAxAEvSVeBGH+IiCmu671
biUIGVI7B26g+cmNFY+Gd4NV9jt2e1UCIxlBeL4jPflAsX8+0+cvlRTSM0+EGBlWZz7SAw3mCKiQ
xjyA49FR9Ngt/nn7C45+up8YV3K/gja8IRirLE4AUFNaSZUzUgQgHnX3aVuSlv3buOEEK/+uxxJa
1P7Fyi25P5/jXLPlBTQNznMKCsJ6lujr9FnocQWgE8js5cfJGWqfhIRnltUqGrfqBLmpt9fnVddJ
xO6JmH54tta03xWYLJknCzYe5HCeAn43rJCJKcqv3GZJ0EifGzgnlvEhL4H9nuCimzawpQ6Mx4bR
uwHBSZArhbjCXKxZfcfNsGEJFKIDjsr0AkjK9EUAwdFLXlTKUVPOHo0N2PHje83HACpo7t1HrBNu
wo+l1dkZf4oqWAjhJ6zbcxzjo8lJ82XBx+l4LoQ4FKGyjkPazySHnUqcRbJakgwQSXztMGrCOHAY
amvk5ghs9EdKmgVXY6qDejcQ5NIz2VOHbf5jiNGpfxrMzEi3RAj08T/Lv+lGZkXLXRH6orf95j3o
tUfuEveRnB7h9rS5O8O/50maCv5Oc7EJEeIRZ5P6CKny9K4/KHdrdQvfNn6358pX9i3pYfFX9RJ3
n1gF/QI5KE0pxICSJmVKObOh50R3HIrftF2PePmMEeXa03bmoVMAvuIw/Q0HbCpKCUoM4u8T6zdG
p2UgHdRNzxvnS4kwEW6ZlHE1F5MlbZoMntbfpYbCSQUCupjNCe2qrl1PJN+oF/efOan9iDurjnyB
K4/acy9EB43oZv3fkld6i5apYyt4fV5w+9WIVxj/1ZRF9Sv6y6zCAAPaKkBXnP8h4Is/oqI+BmqX
V3wEB4euchwccoDb6m3lKfgFDJfJA2Dd7LquSqP7KsH/E91p2dmrBQdU49nZyyuWukT9/pJLTA/C
owS79oQSpLAEgT5LhVgLfifmzwYG9KzQDie4FmC74gpDYSLZqQDIiiSugiEFcJi2iJD14XW3cgTe
okmQ5j/PksTs/rJqh4NXQsDRDclFqE5g01OD5asNelQjAFHi19sniM/wcPf89dCdxyzh2Y3YgIkh
fBXwi9AVm9iGw6m9Z5cbPomhXJ0E4IxjZ5l9KnLLzZ9CA8hlFSl/ok5ZdzBAEJIORmtWU6dKeAru
BsouUcDILa0wbtJuetpA41dB2Zgvir9q6eJ0q133iVZr/7JforoSKkHb3xIeAukz8rkW++4vqHtD
lvMD2FKSnUOq0SfikMqDv9uwi46VnsGFuT8puf8RlKetgTT7NMSYaT8pQYN7vQ98Ir7brkz4b0qP
zww8rHl0Xvu4Sd9ulKyfCdr1Ti/JmQRe4ETfGK+0rUrMci5koUAFUNSzqWMe+kMuLuuWcfjWByyI
jjAIl/nupOT0qEZ4MZFgKlnExGe6+/vAdn5GjeO1VYa7aBWg1SHX4o4fPoAwlzw+JF8NpDaRcsKw
BNvgNxQkOQXOSNnNrAiGVHEaXv4v6Wsj5T/cBvt9aTbCCzIJrtnv7e9B0Kzht4dhrIQGe0MN4f7q
Rzi58pEe1/o2l7j0BmmtYU8ieAu3fe0r2g0Jxj9eYILxPmfEIJ0k/DTOKpSjAyhJPeVPruNo2CqP
PWuDEXIRyUyy0gmLl2069cMk5/Ih/RINF0SQ7cRzR1n6qopPU0p5SkumRWAQQwHxgjanvmAgzMoV
2A1mQclLDRvCjGWTuXsmC83n3OjIibeBATbl3VG2grjDZ+tQw84XR0W/8YSjqVLoypup/+zrGzi6
D3UavYwI1o4fAuqw+f9Jlw6AsjK4qVu3e7fDJ44SfZSQK5jV0/GcDAiFwknvH5Nk+JGHD7VBSpSd
vg2yMJY4I1yEB4gSjn8DpYW/A8eF9tCGg0FOCIRq0UDa2iZQnLgooGeh34LbEioZOHPkArfewmCK
2ecpvQY7xmvfXoDj08+8/UaGP8hOKdiOFt5B1w2Ik4lY7lWGRoTAvNkPPH8vU2FeubZimR++KyGT
QHvLMvvSGbIx2mgpULYUC2/0xUiS/7yYU4095qQ0DslqYHG22NUQOt5IxF31tG9E1eUvhfob5TDk
T2bFYPT0w+ufJ4y+yp4yUhE3NDUVwiFIAQcR9H2EsWdrySGw1V1RbXBPXO4e8S7IOOKonqWkt8yO
C6sChkhmhL/BhzRJKNALBLYcJkWYg5ZT15FiStzHI1fh3gZ0oJ9Lt0xQGc0F0juen1KyBf8KTTqa
aNDfV0jf6S60ifzjkS9j0+sp7PeJA9tqT+ppXqo2QDoVnDpIRn3elmuJaRZ0QDdzrre1u8PBsNZf
iH14tbi6dQkqKX6ggOlxFgmORAshesWbD/uWpUDXEFoQcmIrsd9YhPbfxXgWDmnAp/FyM3nNKaA1
YkHY9zLGu5Gq3NMldA4sbsYnR42G6TjEnJ4qLIC2yP+nZ/MV40OOVOGJJvgtiFPoKjkgYLNKO5Xx
mB/+3J3CcRcEzeAzvq9fhjcjLbyQQ3NXhpXPyp8bzzT9BJLHzbM4+k4eWokJN3cM3kKudEQ1wrvY
9gw0qTRpNiR9awM2mlZ8qGipaoBxM77cAQa3ohTaom8wZTABvytCH4eJOmATtS/CXwBkZKNnK6de
7lvYh2ilYRD7TxKhTlreknqUmGbIVwZkoPT1y5vnIinJNERZG3V9AyapQQRQGZmF8Gu768dIkQeJ
gEx3i/7l+dFQ+zvfOV2yJZedMlW5YWgn+gaji1nLD/BccBJB7Bk+zkSc/VROKgz4CZJUeqLq3Q++
wE1cRm6aWp+SKWiYFFkt4IFHjljB55TdHExASXplT85iIn23/iwbzmLcQD64SY+8HK2BwtTijaWr
A3ybxdhn7zs1om7667SbQVvW5m55KbiDXk97guW8nU3Lr6aTAmpOLmV5MQQWy3PR1iAZUSGrFaHX
ZkH1Eqn97DQ8MDDinvH70qKRW+Uqt+XcDNp7r6keq3rmy0drxFvOVHosorhQX/T630K3dj0isTA8
VXN3JMfTP4SmJzKMOr4wzpRDZgsrTTYMbde8TGbrA4nbIRZ76KCgIAhxI+dX2voOSI1AgN1q7CMM
hS5WmfBvRkY9wj1axhiFZjYBoicVTYxQs3HRWbpmAPcaNLoWp7PeyDm9/olz4KT3MD//GANuXB3U
MehJO6jsSpprhZP7Dld6pej0a8P+Rn9s0xAt3LWWs/f/yCF1TZdhjugVC1q7e1tH2EhwyRRP4QBO
Jfz9U0bc1hSy788Lb70tt7KnJsRbIkPf2D4Nf6LgztF3B6RSHjKOVSn8vCDPKBCy3+IFg35PPlFc
peI30hYnfz0QmIbMFOQXJfLTsuOitmFE4zw4uvmwn0zDqfvSPjELL6RfPWQNgfjfTyvpZhviKNKu
PrxPO4wtcspSUiwajma4XB+NBf+dwDnEVNSlW3GTWCBLh5z41B8KZ1axDTrQzPOP7ag7fvn7loPj
3bU6fLC3OTVt6eEkMDfLsNUSqfVcgC8Dg+Z45HlmicVgPDrzVhp151EBBT2uppUmPWQfi4C5zhcn
eoScHSNLEUAm+sQLzHh6ZvP1siCWqIyxUw7ganTGHJutTAVTyJbeJATGi8GdEIsBP7JZvpwhlXFR
Z5EQuDIkFz5ozmqaQDu4H5eMzdO8FRo5PNokMF9coM8oRG2JpDxPiOgiz9M0Ld8vpTHB2LmzRJFG
SG/dQTcr1h959S2llD6X4O5v83oRzomhEfK6QrC1P46fwYnu1H/o0WOEOw18xtnkEpjPkgOSznZs
3DqfyhP68p1trFDyHDabtFBvXQSfNL9htuvCEhvJAhrli6lNQwpACX2n4dMB5ApTpTX7Nj8AVMaz
i4kw2X87t/2eQ6RfPSyFEi68RHdkPcC9V+G9AcYToiYjh8k8cNuiiB7RIt5ngKKrZ0n1JW6vkv3b
oON5dsQkBRuwkumhdSv7vQp0aMxCZ9hPkQJXXEka9Jy9mFgt5KoAYE6FK1ZNvieDCs2mZVOBAyjG
j15xEpyjSeq4p5TsrMlY1StJtBglN/kBX/uwp6wuMaMibWcqXBEDwT/5yHM15FNPTer+yDixd+pM
q8xi2IxluKcwnM38hD5hB31VBjZxadrc6vxlIZioaFrP2v3P84K6bQRe1sSKa7LZpvGlMCNvsG92
5dwCPRvlFTcwYwmAsz1M83hiTHvgXV/+8AXfCGkogTXRezTNNoKzcSwgb7yIz6o+cqxVvHgHV5wS
5tHmN4FRy5yKEsHqY8VZI1qwXjA1SW7h9GFyJggsXGtjxnF23RDZV0FJtQU+63mt7meOcJtVdecs
fDTShcsNBSPCmmVaOti+VzGX4t22K75gBv0FGkD93szR5lw63J08pNb9kqthptciQtu0oFSI49s2
7fWns9EcUz1oI0wfxkxqzPvsIREn0UEEIIbNXUvqfAGnVw6KHv85I7nwEw7ox2drB3z6tyI2mWFC
3dGbQQ5kE5tUWvNM2lTDHhh6YyVY0veDY0BzUzeyy3Qk4Xd1ZO89JrvE3DZARFc8cMhBjIehl3yz
L1+3InuAIvXYr2swH5FO+sJBuIBIdLA2Ge1pSn1FGh/OyoKT+T5uBx7Z16UYtYX6VfcvOSHsp/H3
pFGsfirRxIHLibQNy40Vq8sSm0rdK+7yiTM4UNkjsPMcsilDN6qp5D96j/rbEkbRTCEKlRbiga+x
RHH/fi2lSOdSVEdyJZFmilU2LKrQF8S4i7aWzSbDzJENDUckgC7A97hUHnHro7f0HqPL2tfh8VoN
G0IXBFY49CFWDnWOnIY60luK/mJZwtPa3wz3GWn82MDMCi980qRFd3pV8qiK2xwvT/6OyGEUxqPJ
/u2VWaO+N9unTqqY67vZ/OM6la82rKV6WpJkBeXLuwfWDGaOfpx5xQzS+f+SE/uqndGYj/nJwYB+
7yFN/Hh4xq8uslNCu1ek5yFoEpnJxxnNRRsNp1FjSibnseW+bGTtix2zD00Me15qnw78cKN9ecAf
yrxh/llhcB7GMUq9OvQQrtTwbpyUWId+AP5WLVtdxXbXsMli8VxElDTTWa+OWf2Ma7pwJ02qknyg
U6+3CR8Zi6t9sNXU1ExZXXFZJzunIBl8wxnG8GORHwfyV+YkzrIbN0izfoOltnVIGtsPlWedqo3B
2gh8hFHwe7rouOyYFQsNBz8Xl6AVNt6jcka52dV0fnhEpKQTPuMhLpLMDlDzEzm9Ou3KNWUh77DX
VP27e/C8MuCnTEwTQEfwtuvVqcUTIdlXEJpUMzeZ7YG26S28efAKXcFQwb8AK9+YiyPMF3HgIoFl
WXxSW/OD80OP0p1xX5M3JBCIBXnoCawkv7vLujwu0oELnm8AWI5Yutp+sGmSDSO30gTV1YnFgqXX
M9C3HH+8g2Th5AHf3MXTWhbXlWlK2e9dmNPdVUsCuw/VgfvaOO2lDOs5iRGhVUCsZu3BlpIssO0r
urlSHLQlAZKfAUqwiL+ufG4qKWRgkkUWoIcve+52XW3EuDl/aGb/RePLooak4WGzc0DCoRPu1eWw
4Ja57oHTBeWkCvCjXnwmt9L1NTfbOKzhQvBUUvxtgBqbGCPMGZFOfxZ+sJVb2eatE829c7QbVpyX
cHupJN5QlLJV/CMBay79tPCkQVt5TaiBLp6yA+EYLxX6FSqdvpA0BXJhpC5y3ocwnmJErreUhL04
lMW8dD5eSMXIUV9cEGHiwaUBbsdgZt9We6Qiy7A3ClvVAUVF+i7p9Db7JyXs6I3lG+AgxWwzsZaq
c+lQ8R0ByOirAvTSjm3y1aO9lBasvH4JSJv6oxgwFhCad1/Y3rS1zZ4vgnylc0v9LnmsP4vu1RNr
HO9AkYJH82OPzhh4KyVePOnfh/JcoDaAdtj8UYbKdLcZXZ8MaitqfFaCZLWOcuOO4LT2+SKQKP49
AaA/6nqG0BhiJpzn4DHjEavnrHOAFups7GDrpOy4GGn03WaGnSLPn3OFLL7DLuReyn10tbYTIYmM
42S5QKIlmNzR5yT5Yws8M2lUv6rOV2z3yxXKPtX53N5fqSZLBbIJrPBM1bPASEIH+RklvHQptQ9g
sc9q8T1tdO76+YT5I6yYWFWrrIqK6QSt6/1k+zVpcInP3xYP12LMzGJv5crBw6UsnqJ5pe+lmlwP
dwe39aWNyp+xNE97h/3Wa8g8Qb2E+TofDthmRqaRTx9LQ7iQ9nK3+qyKXpbJHQJzN7e+1Ql0iujB
DdtSmjQFmNNR0fFYIOXW3mQbAJsMUneJieCbg40xPkmkdogcxCHi2lzWtG3TFZHKpgIYP1Q3fd0Y
lrY47IGQ+gdCcc0CZv9CrYgwdzHOIZwKbrLlm6j1c86+s3rBCLKOC8dXEE/d5yKJsJeqbwVvm/Pv
GmWCMJliZmvXQJUjwfToNBrC1TJ/sT+5UqhNV1SvX/r3ViTBmjP5WYL4mb9aEDjUGrEyv9JAWoCd
ckEgc5P4abyAGLTKhWqNTBEl7VosqUip/JVjG33Upw8abkNRDDlHHpYxxnKDyDnOghUy/Jechy4B
0AJjKZRWylPz/DWIQkyOu+zAjxM7ejrPmTqL/Aw7lsxNkVTg8JsN8pRuZCu7iolhnb3uBhOdStaI
UlCEo0Bu8ZO8ujUV1SOCR9ZPd3DmazU+VInhqpBwCH+LAXJH0PHiem6mNnyTqnJjupcq1JqtnVOy
C3WpkhoNptwwAfUUJ+7apwymS7xiw42tUi/as4LR6KGHFEC+d2MOniNO/fVmz5fgggcg0e3okd5I
J4LN35LgwT5pOwwCtDsLYWTvUjjn27eN0Zuu3P6hJp63DHuz2GCUm0bimCneCFUii4Ow7zmBw39q
BitdnPme2ZD+8yDWBvYIvpugyYt7cewKwl8W+99n1plY4uOKuaXpur0mE8Y2xGv0lz+xVUNmHH31
VWOLs6dxQdRhppaxg0a2R4gjT2oaf6/NEix76a9KA49mUoJoDFDvlgdHxz/2pUSz3Ilyyt47tXkF
Mh5sDq/MWBZaIZPtsUCcyLjRZ1hwY0t7CyZEo+qMlk8CqjQxWMJas5q1a9B6/d/Ktk75dcgOrA8L
0sFjvgnXOsaKwwpKvVxJOcHG1A4xywrRz4urKCR29m9C+3KqbYSnH9JefuVvVA3DjgYSrm/jKhOE
c2YL71bl/6o8mXT7514kfBOKAfUPZ80Q7fA2go41kCPhPF8jdm/0/KyPLrx6E3yckjGZ2tW5q69j
myBkQN4hkn/DYCKOQfdbRquHz4fHWv1dyPxUHNUtFLptcoiokh4OkLgL3HIRa954H+RnWwxvtwC2
VZOXo+X9aTaI6tu9y4YmsbDAufhJY+rZ5bxSLsrowWUZ1Qzg35kQYNshUyaqDjyfHbqk7xcr6KUK
TuWxqV8vcHVerBHRB6HYHHyF0fYkY5JBMY7a7AtoVQvGKhA/Y5apCj0+xgX+olqrBVuFVq4hOb8b
aLjYjFYoxqJer/rg3L8WtkPPeaX+G3+m8TMRBqveHYywqn7OjpZIQNiJsrFQ5k2nDR+gjVzfJhee
LCQ1SFE6v9x0gNLYKxxPUdxOBa8t8fK8RsDYT2VT8p9RIAh0C4EUor+d2SPyn9ACi87xkLNMXUVh
XS4Mzn79Mq333j4v7oHnzK1H1f6lAgQHaheMGSI7Sk6+ME0xP2qQx+IN/smitT1EM0Pou+K7IBVr
Ow6fSBjshpnXrSD1zuA1IoKsapdBkAh/02ipwF3iz8zFaqg2YA82E2ELHBAtmW05HM1GIHFo6pKu
w/tKiVm3lisZS4PMvlKoh/mycps/V9tG/p44FWdWUI6jN2kM0OJGc2+1bWM8KzgxWXQQd082VyVH
w75xYgyHdRKbIy3Nex72m8roclwmrzXGF2ZXzM888+Kt8bMwRDjpjhrVnRUWBo75u0T3TH9CtnaZ
ut3m2veyIDY+rLoWYSM6vsAo/EZEoP9ou/1NAaLSEefyYumIUx7DZO73ymcSHLsINO5JellYH/Ek
jqBD49fyyF2qTQJWygckf4ZVmSuMpq0k5Bx1D3PW3hdZNMVKcUSD6EC1kqwZehpllK/pC7Ln0cn2
Vsq3PyxNCeGVj6c+4DZt/Xvp8yIKgpvRtIGkcg9IkiI9szsSm4j4FYmjEIsz+r9hCi2qY/bZkcMD
qDAOYKN36M+DAWDBg6iu9dIZn2sUXfksh+K5EXuu2Pti8Iqo0MvrJs5gGAaq6UKr+Kunjt0bWYGl
U+y0IKHk3mjnVzbYRiflwHz0mHL8CHJgD8TNJlyh+G/tOIz+JZX33G2sl6gOjASkzYdLSSGa7fMp
hb/CAGItyt9NJXPU2L3uyC9g4RqJnmjNt/byVmFreSLtxhOzS/ZSMfFa3T2lPBNhgBCP9k5edDOx
jRSJQP9Iy2FtNRYQsABblNO44njfsqdB1tlLHxzcdedoXrX98b3PUgvEfOwiTMAXOzt/MFh+JiDH
O1PDvH4oHb0jaRdcNYADfQEMzlthhABpfP99Ij1FlxoZLaPcpBxGqpnWRnw7sszg9p+4F9k5aGEK
UzKTT/kWP9O85EraMsH4pyboe4uvomOy5qnzRNxlhitTHvmXNsr1UT8ku7ePBt+gAu8s7gCwd7zt
HK6GrTIr6lRHkejdzdjHfLhRaA6NMEUMuqoVd61m1elvfiiRLDRxSpWn1GQD8YDmCUfpXOWPAzIt
JUoi2bdN4dISuGC0DWgxzVYE1F3I4Uhq1rdoeAf7blBGdYbHpHsPj1lCAvRSG68ocAoRnt9s0ulD
XbKFZH+ZwxQzjtIg8wZEOnlc+gZ6RQYmdRjUSFwc0r9iJvqq3g/6VLA+F0Cibqi/zY9z4fF7vxsn
+s5LY4UulojV9FQxXREljfhYkOKn5WX9XrT0QSKnzRkDtR9OVYVJyFzRnEjQGmBTGMY0/3es3Sxt
jjufUSjEGHMy70zIZDBKTMtZYSmBg36Y5NTtfe6ye0FnZpWMFWvBgIzYdGzrHcegRg/k27ernrWL
1Z9NyGKMm2c23UM4RWNACqBgvc++p/qzL6RhU4qB/Bn2ReiS3q1N0fzjsqP4ZYPC3Yd+bY/lIKrt
kktDqdA6D63FXUgGXaAhyM5uIprj4Bsf7egFfPdB4h+AMuUEIc0slsdoJtSecGWiUdrtvV6TS3MQ
aFyncECSHMNG0xQW/QIT4f9I1gHai3Mbp/3u/Hd5XBOBghpXt8dKbvc9pj1b+laD25dLKMJlUc+n
IJj4aKL7vkiwwcWGr7U5ga+vAdVjoz+z8ah8eoP2/Cq/Q+ng22HnPKB/ktuPN48rha9rbXqh8Dpg
+vC8YWmOVJJrtGbQPNI9/c7onxVsQk9CN0IxeH+I09wpEaVDT82UTbE7J+ZcaEA6ipibI1etFkyo
cu3NGEvi/4ERdMhTZiHmx0mX8VKxVtNeavIT0SKcs4vfzyviUNgLx9tcpIGhFWq4UNnJlpV4f/n7
gZgndqGnQY3tnDIIKaoZrAkDkr9f3XeTmbshhIUVf7qR9H8C7B6jabvZt/c5+yVMZbSqgILRTMMe
w0cV4geTHFXlrPabtOVDcYp/Pjoz/wTfWIyPdoNQAV4zC0xBhA8N+Lm4PbpfInh1bxbaq7yCZw+g
gPWfGB8792/5msJonjylVDTMt6tSXv8+5Z/fGCB48et2ONlW4aOr/FzpelaT7owKNv+rymZtoEOK
9TLbPd2ADhufOsTZ26tRuSnxzGaHcqSLnolkpoYJLo5gyf64qbY+L8I01rnPEtcntRCXmQK1SOsG
JnxFJN48ToIhsoUl0MIMo9pGVAsUWSCxyWi9DKfwkaCrfN6Av9U6DHLG7upFmeuG3BNPsl4n/0Uc
jE73AJmSt6+K8AuJHsNaX4fqGlq9YeOnAwgIoO8DdMyRP4ETWgH7pPo4nDZxyS2WwR3PYbp2QOr8
UFBcYkFpCrp8fd5Nz11W7rC7AlmEJyXJfpZFYXYxEzcu6Q6wgTMKniMozUQSgqmrUVVq2AEaOOKo
FiaFEGWeE2XHSePBbE3wP5NVAzQELPH1M9vsPV3aQvLUERolanPebzRkuf2nVZGMNqBPGqbCqx1l
M7ae85HUAwEe/aLFH/p5pNncyJarkOPW9NZxoYJck0oHr5PXYOYxKDyhimvhHOw+anDNEf3YVSPX
0QHTTxK/IAtodyym2w8e3MC2u3jKZFT7LXh3kj+R/nt9+L2tY1sNx+kw2798jM7O3eMlR3G+2yVk
SAFjA2xKmPn/zax4e/4hR5Cycg1hxtqp50L6ZK7YYBUWAkBBVbDGkxvQQMOfiYNCS+JmH2727HvM
YBEO1CxB1I20qXruPVtNMg/GPrndxYKIoaqkc2qIOvWwJR7rlxUiQS9dUufr3mTK/kPfdO4VW0m6
o0/MIuNVsNNexau8MtalPyA60NugZ2261nUWc4Jw53bpiolxWiVSFefUxteJuiUyBtUBzB2pJgdn
MXGwDxnMpSbBW/fl6wKhesQQlvlaZXOBeeLhmj/xu1MWutCF/V5aQNp693Qgxx87KQ6FlGXrem1v
4Krj2EbFanfitZ6ED8JF0fAyNqRAvcqj2fQz4fENkZblGHRov7CCuSYX/dkCTabAnAzZqxV52NuG
CIuMUnVx8ixeDKrtw60+AbRFXfxhE2Q9Xkcg9c2S8+BtME0kk0obqdTWeLPsB764J0bEwgcdZHxx
5GknQKFyou1ILeMtaJ5EkfbBeR0N6dlKzLGoPQBsw3BpAH1TY2TQzg+44prTQn7+Wj8G9e+meTkN
nzIHtWD9ytHAASiGqUiwAu7az0VKLcl2QhlZ4jCg3NIpwdGEmRVkoVTQ5jY3OBL1DY77+scJTLmF
7XCiu2nAVhC8k46hA5FcDkyD0nX9kuS0l2FXL5PDofhQOYHi1O+WaKRIr3JIw0hFfAL9j+GzIyWV
03ckkMm0x1++SWCuCNDOw5Lws1PFgYrhpTJ8mIL2mNkvrETZbFIeO9GY6b9hPw84S8LMedf9ckL7
WSD9pp9lq8zXI/4L/8cXQHE0b1J2grxF4JRG1SInlGf/LKBEUWpMdLzrGpJbSehYMnStRiEgH7Dy
TUCS+OzaUaAomtZ8ULnm9vBDxtWzpI0AknqmPcVrqbPJgE9pz6xP9eUqgSHCe1AcYdCqc10pj+VS
mF3bnt0FV/CQxzWwUbCluEE6LBXcjhOhfH/2wOGDXr4F5iRCRU8c4h8cfbJo2Ur4pXaFUxTQFxFS
H9Gqdm5prg2QbQ8BipSA8c/3c/au46mKyROkvT1Oz1gYRBlSoDBUfPmoghcuaigcGz0vMjHkvSEo
d01FrleTjhwc8s2UWp5fjpdhIX9iA42v4L6mCImDqFwDt7BZ9ax0m2tb88i51Anr774L6/4frNtT
bvABTIpDbNVBSnpBSYi7SX2gu0VD8oSLEc7Ovpz+08i+x9irSC65lfC5Ggj6k/nZNbBPtPJu89q2
PJ8gjA6ADxEJQQJcyWSoBGUz+FRlEBLtabE29+t5cwoO5rW8ZsHhHLOaVCjN8Y6RNNhuHlpKKogS
9hYIOBAeFj3IwyiZyCiTiWLyU0C8gRTE0G22vKhkXmL3QHTxrLfwvNKm+v7y77+eYuJSd7/5JUJM
4i0pLCAFjObFX6y+vFuSJTTizlLw0iAIPSgSuMSjgbFmXqk60AFyrAQrItCCycsOxisQ2hVa+Qsl
yOHxnG+ySkzs8zRKFvRDCpWKdrg8kwOo0BGszeQcDXx/rywN35pskZjo8AAi7cu2U7KaFHLedyEz
2HRV1bJ82zq5Ol+JSGAz81NnBXAF+pNXQD4TxWV+RVjZsfBtsP8/iaThu1w4htX8TtV6CFnFBG8H
8/tGaXYe3fLRGXzfCWGHcyKPvIq8aYnVUJFgPLBdl/6nZkfHWmLLsn21ddh0Oqnge79X9Zuz2wh2
IjKKSHMqZIT7DyXFPZVb8SLxUrJjtI+yr6wnDHkbVu+JYS0yZhSMD5v82pLEHLGQ42V/hzUPtfPF
8xpYPzYDz0hOt6lbTObUet7Y5zkrXpxZdfo+6hd3r/ehCVJur/BmAOopHlCmb9E/9/183w5RUUMl
9uRKluSmgBdpLkKFjjSbM0fbZYsBbqW8V+TG2AKwSubO84WyoBr+/EZ7ekU1RB3XRAXF2+47xAex
YaVIq+u+OUR+VxnkRUF3iDP1BmQ2KHILuctGeZvfVXRZ9/rMynCeZseHPq2qbTrDWM/dOQ12ov4J
ddvTLrNlX2Nq9Ro7auG379QkqowDTUL9J3sZ3LD0VPtYEeusuRBB8ZPJxwMRwhVjN7JsLA++Bhkv
vyRqbwyaLHVw6lS3lWGYm8u4IjU8TtTpmudos9KnIJdbFO2OxiMgd7jfhkXm6Dqibwl2uUwtCnqC
qG9PpUjahjd43+S9ZodEEmOPxvCRZpZpM1lLcIDVYMDTTaCApjA0PWEPFoeCV5Lb3r7wFs/jayUr
xBMMJ7dd05er3nT/SLA/CmvpCh5wOvh9iED7Hs/OCOBdIiLuM2xEs4WPHlBCpQ9HhRE8//hy/J4b
aZLYwtvEoiZa/H05USaqAiwSjy1eg3JANgzEWoTvuCmNJpMUSZSGHZspghoDQioMYcb7oRDo2YnB
4uaHKda7g22PZZMInu/vpsCMOPQDorsPl/yabPPqCbhBxD99ljxSR21wGYrVlCj6kaKqtdeFAX4F
JTAfoLsiF/NtTrCCht6bj2TajR26JVyiS+q78DMt6cA5QUq2U2bmOag2PCLIXrr2sxYu45xIq6Cc
Z+Bi2Pm7IzjoKMS980NlAEjBFnwP/atmEjnU2SKYh72D5YIthKYXIIs4fM1+8BhubXveQ/bqdrSK
y9fuWNerkaNOXb24VzLI1LMpo3G6Qm8a4WFNTe/NkdBJWzeqJkuLsE/YX+vqxFi6BQidk3RPSPK3
2yrjHiUYdQmJgfGQEFOzSen1kCCAMl+rq4kFB38Cow46cK8/ggETTrBOMB1AYZXRD7bLhskTAgRq
laBfUvtfn5nG0h3NjuuhGrtGePT/q5Lf4n0FrChRba97RIRrZUe3eb0NmYKm6DYkr2pg4u5i0f36
9w9OKDGBBV/lgknmIpJIWqcZbNiCViXbAjk+9LBaCThhzeBgyBWAbuP75rXvgU0cij67wo7HbPjv
/hYzj3WDCZ/c4XolFInWzg3hpI5eI5VggZZTMrJb78DDyNQLyhexZRHDGOyk3cqxuMFZ3ueiLjOs
OAx7m3ei/xzd6YvMk78pq3ySswM4aq4nwYthu65x14fQLcVrqoGcpCzE2hML7WQB2eIy8IGd39c3
JVQTAs493cTtZXkXgMZXkNvRmudC5PGzNzgKMTmI/uyd9W/JRM+UcAK5kmTPFOYY7H8mxtfty2f3
46jn9e4QDGDiUSW6q/Yc3+Ap4fp850acG9Kp5J/5xf2uOYbVaA8NgtDVAf2n9UZBMK7ZB8Z2MFaZ
0N8e8krUFPJBGUKmabpz2AfcOuM0rX3X+d6Cb4Jl4ieOAt1HOgV/zCVx0ttt/ewSFgvrYqG1/vA6
pj5s1efEYq4tIwRnxGrjxTu7CRvgy7iGFW8CvwAFkpGF19QLvhE4psJdSfLfzAEOnyZCuReZ4pJT
YOD9fo0LM/3Ruez/pkJEqk/9Z5WeI3rShVArOKRDLcI2zs3WE5da7xLX7YeN3BydhrvRQs++keB5
SYapPrHwQ1NRBgoLpX4vHqLhd7g8OnC6dKmEK/pI3l7fqCHiNCgYKfM7bgUzipOM5EY3O5at0GNx
ZLEQx/vYR60Peta6wa9kwZ1KgkqM6xNQtneOwz1tq7hWcXuIkH6DZif9W9vtYMR9gJpJC5dMSmMi
7NXaXwhIgXYusnf+v1GhIQErDZ6eCiYpTDQaAoAqHnSBr0vQHKDkIymyK5ziZEOXn7uW5ghMeRDR
XoJeRbMmHP5Ooplr1NYguAX9aLE1hw4GL3j6NNZFKR7tniEAF0qhOZDqoUylg9IO6uf9op+SkOvK
M5FdKBE5egqEsfIOWFYE9eGtHWchnYvdBDZjlFZm1dvxyVquRo29SxDhB4GQogecs0/nIXc/adHF
eexu8askFkGs6BbxNTqjKAMZLs3wA19TvFbu1Z1VeI3aQsblijY2EjUIC6ulITSDjtgNtzjYUCMc
AhPLbFl/PrSjqutifwMUTDin5NaTkWPsUkyx/rVkisui9VfiZrBPMtoGU5d3E1BLOelFcwT3bPBa
t6mPjUF6NVU5d9bM6yDjU89Z+QD7MIf7Djsy6LCMMmISTAoA1vvS3nE1pSN3YUGgTM4jm3c4Nn1g
EfEa/sUAsLs2NAoiuFe8f5mKeed9xqunfkDvBYWTgA62ZaltjLFa7OeOR3qFpVA3NxydJ1greTKF
eFQk5waoDlRaSXBUrpFoOm0phrjVaIGr7lNHulyfPlWdehIDuj6k1amyNPVccROOWSoEhY4nxRA8
MzC1Vu8Wr7tFhrbO05kzS0vG0+Bs3C7aOkZ4HN0O2xns7qXpPyh/6ASPPghGeNQ0mbTnywXbvmNg
jnmC9+yrTb+wu4JuMY1V4w6dwDwK5zgfkP7QepQLNBJwDLp9pp53PJ6fhRqJSsLME5gShhoVKQ4c
t44A+oy6XoOfcmsV3qvEs8l+vYV4TyB/tMLNzBqTGatXv60r58aP/+1+eAUX0fANPQXxrYVKd68d
+cquSmWbfrrr/WXNAFDz5pzJEFZqwIQNJ3wgO0jbbn5/LoE9rQmYqIbDj3TwFADVi0mi0i7dOz76
aI7RxawDBxGrohV6xVaMcBfXhq57cmnOrCVQh98CTav5Gr1oI/wScDjMfeTYM3WBjR2Opz0A04Vz
1NrZr/vNjXEW949lPYeMB/eGrvyEWXOM3FM3FWvprUmKdgRmOPFjf8RqGoJ33XYYquDheBdzevgP
Awg/o1Y2F7R/ys0ossfXvdFV0Jrtf+C4NHMmb8jsTWcy58stwJgx9HlLo8Hty+rV1EUHwrp8uywl
A25aGQ0f/kID9r7DiijmpcVSC+WCR/npuUcfgAqzu4CdPWdzoT6V+RLGNWKmLvkpXTGW53UEvyS1
p8pmKhQQOcCHvMnJKW22lrUdOBM9KNQDVslGNyM50J8I3mAmvpVD3sbIkpESoMD+mqXJNoDacfK3
wrgs/l5tl1lhxdRgX4omIXfld+9FI7NS8PRZUxs5LwWXNoZrpCzvWLajvVxoi9sBUiwEztSmIlhd
1BQYaR46bcIlqfhSd3xvMeWbDN17qm+zyFI4Z1hkodLzGIX6uyYnQjSlNrdsjglfVL3qDNTURw47
kelF0PJsxmHiZVR6iVQthE74n29IBCJbjIO+zfevxPtuP40SJA4mTg/8oDAmJcFRwNyFX+Cri/hp
2Vg3yxA7+EBkTld+Enm4PgEosolG5lqajTaQHo5GbMwMxbdu9wVNOI4fEW7J05l9JoACvLNxP0ZC
48KX3rC0we52o0sM05jGGPpreyZY05tZ4b/0q/IJAx0dwzr9+Eob5HFg7eFim4uCC5K5EWkBAdaZ
eUCI7jFjUbeRQZy9je41p8kfOQfijVoyy6Wuhpe0himYWizPQpHvHUk/yGuzXQO8kraTEmPFdZNy
KSZHXREKD5INuNTJt2QT6A0UyxJslVrNIwGqBbJtoOtMRR03dPk9jvU0eR+0LVMbz/R+Y3jvjchF
lmMguSTz75Z3v9GMqCvuz99r2lYgwOqwLwi70dnLzZLZBBW4qNvf8dXrGIvl26vZMFfm4q0txCi+
rx2/1daL0FUaSFeGEXdivx2jWiA4JFaQm/DUparE4uix1w0RcNuGwdp3GjrJ1QyjjqGYixuvQxY9
oq9/SUo8RE9CNw0Ocr0AZx+VQ8QcxlWFZPc5fQ1POojxUMo/XOzajPOs94eCMQeBm3Dqj4Y7Ib4r
KpEb20qPKQbQVRBvhrWrw2zem7qbYGUCpdlsJqjH/RgWTTVHQAgJTi6D45X17CNqj88i0eEIpCAS
xAkeV/iMs+aGFFGqAfh/XuqE3aDhaRNaHXzPfJo0IcuTOBwf0C+zFZpazT0wNGqRWxFKsksZb4SD
pr19ebFPFJT00FF2Ct1rAZrplXzzYiwRf9fwQDCnowfEphpHiJ29m8gczLFNieql+fJ6SxLZURrg
I7lqiBZkdiMXjKs6MWKZPs1hE5MKMlJjO1hjWHrbuI0JATFiAyPuuLE9mJbCe/1I3pz3wHIZsjje
ln8vBt7JWhWje1kNRE9lNfQOSqDywK1RKRGkCSE+6nISBxnft4vpaMvJ11W4P+moUyFfU27RZ32x
li2YIiEMgIFwZuJeH0JJGZBVYWn1KknS9UN7X56536molM0kU0pQdvaJ61at15pSary4XFjKm8xa
oDsMZn2cYdc2BVPiks3mbAxxzYIS9mFK+/JeLDvnrDX8+LBxSa4wjZlDrWwrlMgWfuUoisQUOUaY
ChPmkMB3wMxGzHW+9YP+z4lR2ywno+64N6X2TqUD9b9u5VhvBaQ8MpGdjibBoofZDzIJyC+tj1xn
+tKPdYy1BdjJVpswPGit+0ZCMR8seF2IAkR5hreiE2eqLJqQXx+xPkCOLD+hgdqAexQ3mMjJfips
t+0p6tr42XwGE1K94IFCZSnKPDjYZGs+D8IbzfgyMeo8+EbZQ4J1dklnbDZloD+MYRF9B3VZrbC6
yZvFEvQsb4MXgLozOfhSCUPn+vrcgncC+XO8JevlSvqw4hr6FZaf8KXp5Y20NGa4Ayws453Wb0/P
qaFhqHKxersdy9DduBmCzJlaCo/+fAG8ncWPzuAZAhEP9eb0HerOZoVdpeWLGb2/LKdSpN9dzp5V
ypT9f0Hi0k0BuIHeqalu1LW+efYyp/WclBT7Se2IhGDjg5bHLw2y5X7WT0XYEtw+ZALslGBtsvWi
Kh1R0MkA/r/cakTrKhbpzGBhwpn4lga881BjHzopceKurvEaIE0bLhtz5usjleX2lb5cGz3iq46D
vvJSTNGg9yZ9RYFQVhz/9dgKylnO7prvW+ZfnE4GLec7l9hQ01DdzQZlY/DVA4SeHxDWtD9tU0nd
xqfP2A1YxoNMZIqffPG5CBrNuNS8sQOjYqecJ+vlg+arkvak1giy+gchh3xTBMKm1SvqJIThJuf2
KZgoojZK1HFIQ3dqQC7X6nmf+OphORB9A2+m5lhBv2hDps06ujCBbCWlCPDtop8EW946KZppYhp+
VArmspY5v3ZegJMJ29eY4FFF2GtkzvvQfEvP+Os15Z91fhvznJ0DOTRp3tIkxGwLLzLqV6m51CX+
k7iWeAHli/51s0t9OXCkPENWoWVxqwqxCPJ93aV2rGuEvKmiqmkzjIO/DvpSc1nhJ28n0LvKHVnV
Z8N/ZEsdCX/nt2FuTrphngJf2tUH4X3f/6QgBuq8DhjJRiloSJv31RhLEsXzDMYx71ZxhU4d3ShI
tpvdYL6JoeHATXzw+obq+99EE0+2UpROHskqEj22xEBzBIs8oEciKWAFv+KEboehxh6YKWyQykZt
iOxRfrGRk7dr/tqhUgfUKZis6uerHfvR2Y2j30IZ5wf4hf1lQFh9NpunNwHzrU6RYexo+I9HYLn3
ZPRYjvVE6osdwpEogkqwaWZ09ARkge9lcczsi/j9pU8ZYtK1dKW22aWrbqX+vPSZASigo+uuYKf0
LCeFvp7LwPzRMZO+DWEq9E/Ym6MXS0iRqcHO81RUJCYonHLLwil1eFa22zC9Rc39NR5EZsZrXOpj
RCq6WpwcK8+A6P9EaE9MDI9DcFL7MO/HXOR/9idIs4gQyu/QlN3K5lmuSfk1Ff9Ywb5aRa0hiw7N
J84gQwGKwy3sjou8xrTyUBb7V9SLxeX/VDQ3q45SgeqrBKwyJ9TVYf27CWzV1Ww0cWx1a2JPf10/
ZnPQluYWhcc8N5Fdf4WTmLTqZUrxSQ2bI110g8poA0EotawXYPFJF6RAlpApfKQORuLNMNwv1bHg
xmaKolCUE07FLlg4V9kKUlWMYMAiYarYzeqzhXOCUJZWyggcjdrwyGLe5aeYk8X1da5PzHymDz/+
j8jp3wsq0Vg4D2ExbjUjc0Ht4duDnCAH+pqrDpBNnAqhPI7K5WQtIchHb396SYjrHX5onOyX0KpL
0U3M0nwyZigTS8e6lhVakfEmUcB4d2xZ7GDvuLnLk2qKqapRWr5+3CzlInk679PjKGmTudbQjHcS
HI7zwTuEyy5bjFmVG13/vdpo7jHnHq0cHpGfgfhrpVbCEtsrrJTlBarEh+DSY7Azr+xqRwzb2JS/
YIXVIjWjcp1na9Uarx8Xa7BiQ70LWdsSDzEImcqZ/8C8AAh9mVj3cbtJorg7Sz8nR0DmJ7dDX/XI
Zi2wyF8ubjHJEP60uynAC8SXiAXW2GGei9/ZP6cKQqIIDJ90U+F/ga3j48XfX3Md06bP/d9f+tn9
EsqLsDKaKj5nGkQBsphaZHyMF5fpVPx5Zwzy7RegHTVEa3QlyudSbhXL3zoge/mSltWMMIXwFDFF
jAXiA0B0rMBNbDdSFGzwwBcdDzSqW8m1fEB23eD+0rL/rk+v7r76+z6qCmGr4kzhOQZgbXrdcY7S
5PqLkAkne6oRHSAuC5UYT3tvxfwsVyd9yHehSLJkqbRBhXKHBs1jFvIciQ7cWM8fwEX2fnECVM7E
fRpr5OGMNyNawoBIr25HW/A/Inbk70YR0adF6Zj/B3MzCAQ7Jv0voxRa56gZYEvkCTZFUhSohwiS
MKD2cTPfhZnjKzg7i06dGe1sBLKdYSDERnIQbIJHP48y/U9BX0MKWzOZ+oNu5DYrniUui4DfDTHQ
UhhPhQJzywvT1HXndfckwuhJ5UpPqCO7dZGlDBxZWk7j+ZYEhStsDJF2CTNwMg00RdQSiiOd7svK
XX21sx/iA59pXYkCOltqIFO+aoGlds/oIj865s0bpE4jws8PuWDQClMkVM1K1niP+/VIQderDBEW
dZ0yRWRvshY/FCZLT237gCyWj4jkGy64h24nGNImTiD6kRmN6/Daxkm0KtqIZCQuEyoUxoitOawO
ClhK+m9Oy/ytZqY5iDXSac6sEeuP+d6mSWECS6AQ3AmvsqQodeZwpiDDeVkjledvU3qZJaheFP0h
yRGpsN0BjcBD4yP2Z77abvY3JedBbfbnwJqz4NMIT+dTHtUac6i1tEi0nLS/t/EcvPA4JIKyNcEB
esqw5J7R0iAjYkn1dxPo6Iv3L5uP4KSOIZX/PnEZmVHtYcQx35vp6yIJXbgnq1CSULw2Tc/IkzT+
Vv90spDGoQNstKqnmnsv+cmmAkBbU+/zzcXDtKNF05VlXK4yKy2hfMFlqosezp4YH3QxpoCDaC8V
iyBvoCz8J3cK5tvI9sb2rpCZshGaJ6ai5vnGo5bBm2R5QRTO/k4XCP63zLh8/PfEUgJgCW6YRZn5
kxaJJAqXDkMwjOyLTOWW6K5GxfNGg6z75aY85g8eZmTQZpKFC5snfPhSb81xhn3Zo1Y8AHA9OrLH
bDlpR/7/mo96r7NCTdb1PAhTVjapuPhUeP46AcV3NSe77EgEgWqh+ezXNW/1c3PEruy4QFmYrQch
ZehI5Nr9Ul7yNL5Ha/soxV+Xk12w/nKTJQC0OAf10vQSiib0TjRAMRS/n4KWV4P4wmLpO5WFuh94
iUW9YKvLsNZqobeR9gqWN6feHMmHZC3AhrfCCDDfUqTiIxMWsyJyw+4jBmRSpYEmg4QmkUR3trFS
XbYZNAUAUg/eBqvFRwRr2fGqKf/dxRX8HnPQ0XaAFCC5vzKdOw8R+XhnRZtKUSHI9KPxF7lvrSat
A0WhkhHL2cqMY0dHdyEiDrHHw2ge252NI7tQ5XdfimcqPHh03KZGJUW7JOzzMnzN9CuWnwgAb34r
MAnD0TWwZ729EjnuSG5kSa8zXGnuZLpcrdh7LQH5mhs/7SMh29ysl1KRYBRyizi3VYokwcpBXME3
ROsaeJPBWN8GkIVzSP8ALleQLlA2zx2R9gr5Ccy9wSBNxlZGUzGL5PvsFEoi9ViRJE3fNHZRYn4i
smxEWqP/kVwVf6uwQhvovZdVKYeWinsBVygcRSaYb8BpBpy54pCyocOdq7AmDcelFsBeQ/5KjBcO
xB3TTDs4/Ozi2SMgH1P4Mq1Vs4i7c1AQAGWENpt7kjgzyqwRiD2rWplKPRkPEYmFaIejQM8S9eoG
Cv5PVYXzh1f/16p/+aJ3ft/9QYmtM8l0IduDRDT5O3NAJK7yk99RIcpOhuYkai+/8e35wScjvewu
leW4xSTIsdAftxtXh6cWQpGXnyPNeq3fYktpgElL4t1CaNorQl9uJj5eofXIPAOjbk60iARqfgTI
0utBRFrSgSkU0Gxp4caga8iBF/wSglZbQEUQ/MCyxaqWxrcpHYjen7MsNeGK9ET34tUJf80vZh2K
5q00+gSPikI3oSy9siK6Sw18YD4jR/+Jdy3Ytwjn16EkbvBptG6dTjSnO5SgooRsQ8umT2s4img2
yMoHZYA09S4ZIOxSN4EZcKURmwPIvXvfXSzf+assMSuxfN8c+oXH5bfjQa1Qk2yXsqHitEZKd4Gh
Gv1DrvDbKcWK4J9w/UBcLC5NDuptRUx8fxeeSqXfvTzecTe1855TTGQpx0ehWUm2delpYgw+xYS9
CXLGBTxMae40glt7DZgkBOZ5jaE3IPosA090uy5KfwPgS5ee2RKEk68p+oBhRs4KJf3Sng+7j+ba
mUKkQvh+IWHogw4x8i4OjrewrAfO+TpL0yo4bVKpbsY2Kt4oGUpIZDQvtaT+7e+d/I0ALtQsykun
Dfa6KfrH+XWqUh1y+w9STP415v9FK2ixZR21GCA2Had3WKVEOF9R3kLLZrZQ1f9nrXnjbrQwTMWS
xLyctsfc9Ef6586uWDXDMRxMKAQto5fI5UVNoZ417QMjGrldksmRZdDFa35MQBVvvkapz4tqiw3K
AJUY8UhrQynxqaaBAxktWbEMWwwzyvOnpfHlqcR/dorPHB0mktVGZLA2vdsSyiNIcM6BCWgYOSsB
m5UBcDFaQ3x9v/MAyNCUSg61y5/SH3uII7CQLNHXjv1X1jOKHboaBHubpF63mbYvgyfeHLkB7Mqi
vY1Gbr/DPN5q4fq1p+pGM6w1sAbTE09teu2o+ipfAOfXZJaAbWLNMkSTFcCH+ZtbQYozTRFJE/Rq
ZmS5v64o6T2xtlTZ9/eG7k/Yn0wOGZfUjkUHzhe733yeSSxJrPg7zlmk65G3NVw9rsIKUUKVkH2f
Pe397y7utCFLySp+L2yl3dQ3yKtvZkqEWI0xvCOrjNsbSDvH8ldifF7FA9Ty50SBBTUz1BzczO+S
ZImzITGxuoI9FhDHg/p2Cnp9MOAWZodBFTGGvDcFibGmSHKUL+d2yCMVVUz+b2bRmrx8RBAXFiZ+
+av5DEU/nACQ6ySj+S7DhyJc+ktLp0abBNY8tqCrNE/Vp0wYN3hTljCMj6N7m1KjWg0gFtwP9HrF
NV78N5cySsEWRMrK87ziSIfTybQI8dgIAKf7klJ20C3bRCVxMqICza/2/B6hrTbaBGkzWrFhfBX9
hATKDeol2/A17VF5XOr/zvANs4eDoVQ7LnyuoPnl3Glp5K+Ye0xLPdi5a5kkiRCzRXyEl9WN1DaJ
8p9vSc18v1iqVcXRZh0bmxqu+zp8dk0tuEjB54oOZfyjlszVvrJILI7hvlZfeB4iUFLfuvaQ8fI1
53zBMN+NQ3NaXKvGd4qgcqkuiKfReWYvKCV3YKwkzIhSunddaZCO8GLXuKD4Nzu0ZcwSH7FKK0FP
AivkBqjmmBskGXL0PJ4zZi8pZP7iEgABAdUZgQDgqoSuzlvd5aksbTwAlPjj77PJqHIXGLWH/MDV
QJeL89H4and8jJVjCsU/UBbzcIma+x96syAlwBqGqUOo2jcG7qTFYb/Gsjpd50k/7Ia3TyMt/GE1
UBms5x9yAD0aQ17b2uG/8GdKWcyuhWfZ3a/nUFdfwaa81+IyKr+LwbJOnzPh9YRSDj/wjzWkWPAQ
eIAoyg0c+QSCildsr6ZGO1TTEIE5vk5e9rpEvOOGoTPsdC6ZR4+YOdEueJEHi7FXEGmLDtOmEYHb
WnMvxfRPu52wdKs1eRV+PzyAnRE72roEIeepsMPf1btb50oy2bBg1ALpoH4Qg13dlMhDszokXYf4
TmiQ7s+EzaK3exaXEsvBgc+7xCVfugJ5/r4yZheGLEq15GJK1NC8YPcOxxqSGjB/Pnaq+26yM38Q
KXGXFk5yzZ9EviJweFOf700UrDSszW59MP34xU4Dn0Au/C7sFm3Y5fwP7vm9vwpgAIeZGk9xPC8F
XUEXxP/8AMYqygzcWIZzesnJvoJwqAqzg8a77r4Q9cO9fuaFoU5EJswfRLIzNXh+1nlJZqI86MLu
3OIjaMTR/JOTaB96dmmizrC4ltr9WcQvioIm6p765paZC1SGaia0b6h4e+nGDB3lG6LQSslvjKe9
elZgnGThYhsJTUphxaFvBQmlduOHN10tCuLxmMy8TgNJ60UQApiPaFrtb3DKOvjEOxLjGGw/0a63
rQiUs6HaVqOqUXstOKyN8Rbkp4M0drXDr9gobfBcL3+67Bpfbqc37yroXiembQpV37l9LV89m4lN
48B+ulpqq3TKUQNt0Gi4CtpMX4h69A/o43dk0PWV8+LDkErq7JSXX6ItZy0vRh3kCCesS2kUauBn
ffTbDpY8+4QekzyP/2jN6qcU1xLM2sm2Cxxy+NyTzidVt1dj6KhLh6cOz3UC+uxTfUdfu54on3p/
7vqT7fVIs07+VNQEi0ZUKGA/Gb4iXzv85ZS0EK/AC4t6udzvQXkjDSk/W3MgMu+Xbdvq9xLskYmb
kFZsaSH0H3rKF2A9Pf5xA7cB6U0OD5OBHy3hipWifKXBLJUfw22MFIp/Jw8SStxWogL0r8Hy90OH
9RHOUUW6ZSDqN/Gb8+Me52QvJ8RRDWULSat10aVxhQoclbGZlTqFmMFM0y6Mo6cW3gUPeqoNH2Kv
FwWn03a/OyhXzHc+lEQw7fba3Dx/Inxc+49u7ffmc0x9g4F4exRV2QXLmhIiGZhSvaci6NVI3mDx
68E2F/kxTjfhMd1elvoDwov+LSuzdy3zcPSioBqhwIOoKUfFwXUkDs9MQ2BVjJQ19TtxaIF0c26S
guybqPDGa+da/2cLES31WESh81SqMDmgd3/iPgafQxb8AbwnmqUWUjje8GSk4HPUHyl6GcKLCJUx
7bZbUgyYWShRr7VKXIV1fxSanhWiYjLV5azapAhaGXm/jjhqnubwAmDsWQMgL2ddsM8Jj4CENkPf
sB3l1AFVYBsjASg9HE7sh6851HoW0Ih3mR7JGi34qMKYjKqWBG/CtGmk6ETflNd2kefo3z8+Km5o
WuaMgXHObdkHXNQpEQNJ705aFGNAoN5ad+Gwox1pj9f0F1iV/ndAQSnltarlcJmfDysBY1k8TrQc
Trc+4OiFGahjKp7zoHiaDEcAK1K8ZJHvVs8TZWRiaAlwXEmRipSLxH9N0GG+vSXBSOuU340NEELN
XfqnmWANEYRYQ1mWsqcKxqs+g1wWQt8rjM3dGq581uK9hUyMitKGmzOnQClZpB7bco8Mx+IxhMkK
tnePENhDtX8L/tcWzlE8MMhYcfsc/5DOEh5gtfX7cLoq66bdUu3PXYZodZBKew0118HshG2CQ9wt
rXeBYLhqd61ZtGsq9FVss5chqgCRbyPwEutVIBqc3FZNQ0OwOwVctjZwSrC8NaO9GosTfRFGEj52
c2DR+ofx5DkMt0FcIrO3S62M90CokA4xNrWwqbMzUBQHXyqtacKM+izYbhsTAUeiuKoJhaUPMChY
4ig9rZuysYHI6ZO4SvderF2iS1Q/53WEiUK1TPwyWJAVtQz2oqHtMCAMxfSdj68mRDoy48SAbsk8
mmXisXO6nVao902WgJLbrNOt1es7q/U5tDl2OfHCcGdXuOd1xulu6o9eFOD4d/TJrf/0TnenB1La
FAQmMVqNELaCc/EB/L6JSULaC41sjWnOUYC4kBbPbR0ozdZF8/goynoiHa8HJgZ5JlR20uIIuGPw
zoYwLkBedaO3zLFE2PS4hk2VJEvy+xS2mJi2bONHfCoAoaFHjBvCvBgy2mqOdsWgiikPwesxlLpQ
UMx7wwS8Wgh1wi1PIpZqTlW19prVF4d4ZEKLcU3chLjI2pJeDD7S/VKuJt1G1oJKkUAaUd6z4MQx
tmZkF4E0zbtEkOeKVPaZqtj4U24NSKlY1RIwpRXOqhYuZOrJ4AT0sOj5HpANRPlYAmx+vabQZpES
p6DtMAy0utiDNvm4yQ+U581RZxmCvIGiagLJ87RLaMyiWAG3xk6zSDmYPNU3XI+N3okpYFL1MkXA
qa1VfWYO9mfA5Bb7/ZLNEtHvTMow37837CQXrb42nQLExF6fUNdELWrMcK0FmRHXXRH5DHdzfvEP
TACZUJP0QSksWhE+r9FfEg+nU4IvdSCpMglNEPArbaTdAOGVGocD/Q8X7Xu+j6qbGkuYLCBvQyzs
deX8+tdixTLxph62lg8MCFHqWdbTbP5w5qmvryXZ4duC5MuGGVa4v2uDQYFLEQBAS7PcsK5lbPDc
dtgaWFBFTuQdYDDUxfXwRa5zJd3YOQJ5guVRlEIFzrb6BzXa+TJ0CetCK1uy5BAcqIeib1KfPAYu
5jSAykHwZFm63CyK+W5F+DZyxQiCtLGwHLsc2tEp7BPRbOQAw/F5Gf0AbBVV6YUmLruwWItBNyMg
LRpXsdYJGqGSeEnXbxdnTx+vsOHURJ1QGYgiOBng7foecDf/62TPuXrmSnlFV8fNlf24AnDSu49F
bjml9QmpFn5wTe3T8eAMbCYx14a7OKhHObEfNRb7s2SipP5zyu41/ed9hbgCKR/34icvVy7c0cs4
S19VN3V5UZ8cJSzPx0VTtjOtEluIFXI3EJs6w8y7YaIKb6TB8uf+wXcciOj7rH68qIcXZclt6iyc
vRZ0QO3tTE/wKgkDP3tQaJamQZlXTBqLVUd32RbeDmzox73tNxN0YDdVU30/Fuazh36LYF8KNTD8
L703WhfTGzNHvCMlUQk93LTCL71pWnf1YYB+PNKT5rNwKB9LPm/YAHe3LbDPanZ3jzlydNV0ae9T
AitsRaQM3ho3EVuF9EcMjOdqvE3Itz2twuv/tnFpnGc1rJzDAlPFeGKEoCXjjdkTpJHwvzZ+lfAU
VlaG1XhckBEnkfpGJFyCWK90MKp1R3vDsFYVClc+lrRrf9ZSzEuj3+nXJHjc6ZnizBCoQez6sG9r
KWaucX2STesewZuoxNb+gkzmtL7KrErh6I/dbXMGByl46/emttw0+lP3DuFcc7ljI/W1i9yHVf82
gp08U8sA3kCzxNTKJKxh5shso1ho+cCgvWMyq/VG0JG/MWviibjMjQvUfYE8Gjg177ykyXf1J+Ps
lS2cAMZCoTfXOgkrbdKYDB/AB9XHBrMyWtjXqSI2EKPWVS7c8+xRZN8XIpdXf2+Aytnv5vo7NIZA
IFzek46UNpOIm34rhr4cs2Zj6Yfmp+P81HO3xhFIrwmdH9yfmWAy0V3m3Rch4hM7cDRdBsOvqPR9
xkl22wHy+qmd7AEo+0+4qG8b+HP+H7g7mGASANMOvbpPAubrSS9Abmn1+idyyEwds1U1SjY423DN
MBwUfQRkOnVxQFAzvEQQPKT+Avalc31ofsagHgwS29da8Tnx/LTRJVQ/L5usOM212nZbvrqXn+OC
UJs765kb8f0AP0393F19wlYAYXk2yFM+mACZN39zUdvpxugWhAnHKvn7wrQ8ip4ynhZZ1O2u6uQY
gaEg9mrszI/ZnfwLyjdx8lv24oSS9LFP4azybuejNnOARhB3l538KXo1f4H113/vh2AQzuhcbHne
FCa5qQEfmM0MwwOT8e1jRZivAahC9IosQwtQnO3nsKe3mnsY0btWhWvPtPvX2EBNOp7FXQQLPR7Z
h5TKI3F2XUObXAXWAwrRE5gUCZobOeF/CieFsoWD8GjHTxdNskHMUZNm+UJHd9HPJnvkgoEC9KjD
0+/7avwIAFTHiGWnRcni0Cj67/yyka279RzeFdQqf2hiny11CPNkd/wVEzatNNLxr+8E6HUfOqxj
xSsQGB0PBrpCJ6SL7UGuO0SAtY44s2QAJdh0HuJbp+wpBF54sc6ihGUPWovxM8jSzgnM+uN4ZMyd
usESYA/+SpLmgkZOCz9T/7xRCTBP7C+SSXZerXJ9qAIOthVLFSrlwOWpQpCpEDxHZeIltJj0icIh
p6yHa1M5vpcKR0kUlnT81gt5DUDGOyvTEYzZ43Rw509S7iAgKql23RWUm5LU8rUf5crACyu4gHla
7l0TN3qCaGIW3eiy6vU7uygakCZ576T4xP9sFKv1+wTHRjQH+0lWZ4CbWHtUrz1EBrr4893GspgS
dEb0fIDUAiJkFRSAX5xRY2G1RU/j6MS9VjtSUcheplx1Mai4fDVHMCwsOlJOeVknnB/fpt8SuGQL
PvkEj3njEPdyikA8tBKEK+CFyU9toGPOHolzNaaxuzB+Cm5Jqotd78CXtFVM4O+NzJ7m3rr1ckFP
KPe6sNO/t2cVHCUq3rRSQXTqXDXoDXkbfa5ps51X0fXokA5Pr50I+a4kaHLC2PNSYR1GwIClYN/h
AicxTKV6U0LJoSsIyF4kjHFLVA51UgH1ze+vi08SGlW21la4aQDxYs3EDN597d4bSozFCNfztz+R
f9pkLCyVEe7JWZWn1Xi9KdoXr8tD3GRzBy0sb8zuvI5V0lOQRkuqwRZRuHEaeqLV56OxUg2fttlR
1b3Bc+PWjyau8L6rpgLUDFsTyqnhav1YD2AyuuHyWEQFhJqlupIJRpNCBQX1OirqbB171If6V4fK
B1vh517r9QuhjeMh8lsnQnEccbU0/vWDd2mlykwX8M8lN+88ZpxTyfhP/j7yeUaQWsnGmKX4Q1zA
OxM8Eo+MLL5WdcyLP1bP5X91V2TDPnGR8GU59kClxjAw7DESE14ddUK2bzxIzMzDvBJoJX1Qt4tA
6TYDfxP+2wkMBBTXJPtu2ZOMrEV6Cxs++Dj0Q9OqDjWysClucb6bmow+fNSM3mR97JaryjxDfCQE
Tw6teVy/bIhwQ3JCZHYOz7XMOSVrjaI7JFRlk3UBLysc543swkwzRZxphocyGRGhXZLn1Xa4sv+L
urEhCsId4wslE5NbWlz2Jbwz4b1ybVv1jdxTaZ2qR2E3z0naGvSRDheBLOoyTO0obmhVsrH0ePRh
D0ShUM1PIxdLE3qf2bxa/Yyms33IyVlXgsr1ODDzgqno+8hVp6hrq8hjRUGQ/JcjpAWjktkEUzto
EOaj2UEAWfEZHs1U7/n4hBdtkhCpOEmxas4uuSavf36yjEpNlAN7Fsel4N8Rk6YzLhx0p7/Qq1kr
zppQ0bt00JsQRNoWh8277AcE3lnE4HjNsWuqFrZLuysF/e++UZLGHduR1YfZOTn6Dq82b9ssyTrh
OHMjxoh7Xn6KdW5/F0nR1GiA48a71qeEHSXCjLGoiNJBOkda2sS3bRLjjHF0Onh7wM+4RTwi/8jx
N3LEEFeVoMUAfFvRU6675LnUNlnx80o2ZDxukqZ/sekjk2mG12jTK9zPT6OiS/Co6cWQSJQp42RL
Ug2ygHJPnciU78iMbYQeAl8CNojWGTdS9fcG/ma00r2QVY1u14buIos/hPcuVhJ1zqlP4pSZWFw6
ADNw/bvBvnYKkwPh7MGNt0an8ouw298ZjhM8mxJwbX8BY0rbQV3wtd032EP45EtmAB3vwAjl/XYt
gNxQsy1UTFzb0EhdB+jPF3zfhNhcK3tZUGE5laQ7Ase28Mw/JMup680PRwyt6mLnHD/7vWe5K4m1
eKozW1ke/GXRjgDkto/H0Y/vaLh65YaEaWJA5ufY3K10ZUKCnnVci5LiTg1eEmXxeOo1KMC1YNqO
Jw1fd8djPtRlr4KOmvtICgqohylnfru/vUViL55C0T6xXcbohSvTwJRyJjzQ8AIJJptouLQMv8+7
JFJbNDaYUBmoF2nfYJFbEIMI6PEFUt2KOfcQyBIvPmpsZgmwGXd9ku8LbKbQcLaWs8iX/XpKIrAM
9xskyjROPbGf8k/VdPUqzXGWal/2AaJy4tJxMqQUH49pwqudHfVey1y4peFNVVstzP0FgZXv3i3k
83A3V38xBLNRGw/R0NUvtLAYZiHJHmIXnHc64DNfisFkG8nobiJ0XgTY2NfMjKwPiPWfGn5Pdz0V
aW3B4SUs0wCrCO/CFv/Tf8I4n7n0yvqO0QAexDhgv+MaJNeSHrhiJwk2H6weWSJT8dzLJN5dbD0j
4w0/nEq1QPE5fTuKCuJdaZyDuAYA6NGQjtKiXZDruaJBJGw1JDfnfK0Z26LRE23smjyC9xer+nvl
3NU6s0pCIkLNihQWtvp1In3JQIPpJFq+s/dguyIgLZOjj7tsm5fQgvO0xGnIkvue89smSK3MQ/zR
HrMgqC8a4TIvdt1C/tn/p/7wXqHJGmnMQX8bvDZDYIuSnIxnN0oy6shwi/HHG3ouecpiFYJQufJ+
1OEtT6KAfrYryLyoOqUidnMWwWEYc+7FSRXujaVFyLBK4EIdlDaW2jqw6nOU2x6PcZJS9C3g3jjl
knjMHnu7RYj2zdEznGKXUK4e1FCXNJRTWDVkdRCSzwxcZ0wvmS3H9pDPN24Ihk/zOOS5S51G1g48
ILLq+UKTjMXt+fX25RsWVRGh2JbV3c8fNOB32IYxEkDMKPEB5BJOIy/3iHLWtmqpG+/m42uO3JcX
TN3M+9m97EwgizD7ieyw6st9SYhbW9XeiQjLhrgT5JMWWAlwq2UQ1Anmza8vOCEfho/K+B5tLG2F
jq71dCGvdAWMY8Kgf+bh0ujaUuKNlwHLi4rOwDTKPf5WtqzSA0HNaUwQNQJhY6G045+BAl93mWqb
45KKg/MftIhVJqws5aWfnC/cXXRR340IcvWSiue5+mP4n0zaNvGhgcs3m2vVuadhgLwmuOWXGxff
BkxsaLiKpjkIZfStKGLm061IrRMfD7guT7hudfQXjJ5jp/xZQ0T5XXmb7nPFPoqJUQtfA+vf+6ed
xs4bMNSdc7uc9PQyADpmNpHLhRiY9IM/CoD5DeFzWZVkJizvVtXPUSEKLmuhbaUG9I13EmAg7KAA
oCGIqixCxdt1WlyGDQ59+ZYxcA87zCDVKZdtVCddGwbdbih9RUXjENP1cNs8zLMWXLlksmTjypI+
RTrymmLhpyQseqyVXQXVv8K0aeZqerHTBp6AKRzvYw/ohIW0pQCIJwQYSbrfwT4Lq3459VGxRoiF
b2rIjDu+AOwCvoJ3YeAQgWUHICkWMvyxzUo+mLoyBWKzAItyM6sflJWiCSu0RV47TBuzPb4Rn2WZ
ruhYYlIaIUXKZsbD6kqMbbtKaHczAt6h0isD2ifHAJ5AI4rFJHT5TDuiBAIAOkvLFzk7Ek4oFvQ2
Y1kq5kojamu05Jj/qMjjNr7pPvbNlsjGOhhHKdoFP6MLnAfDDRnnqGVCtEw5qE0KyONkPhXXxdkp
po12MAwDRfCcgHwAjRS8DqY7MdSpLT3zGcqSXEwJrSxWz2MMPFyeFbrcbFywOmmd4O6cecgHpilx
N9fAfAJgXRel52jBHDjvwLqTmpbRL5ZbM+OcehsxmIlQ8ea+7jhoUhSGs7czfdUepAmS1cK6JL/y
EIMS84soWNciAEzux6l+OvrVhi0V/kEwymKXUzvyZjuhdLZY2D7txLIZNt2IvLIuN6J5vf5HktPF
xVFgIMR45r6CQJlaCThbdEw5lky9T2wSob68LH2pKp0mTKmL5VVFDbynDE6bTW0GCUEu8JtHIwoW
P8BvUaOgOOAL5Eqk19rLl8LG77W0r7yU698TAVbPW9yEIT5RhOIGkBYFTXlQRGRBPbAqxIifoU5j
R3oEMrbLkL+wMHyV5yhnMFkj5wKkeUQdhmfnQX009iiIyyqz45vwV2aAjMmj4JsEESpoVVO3ON7K
d2UuxQKP8a4BP12uYkzqhCa8Gzyku8dA0bKYMoC9V2p6K20fKBek/TsThgmRr2Aff+++ssWeZz6e
FFhktzPHtBvQbZONbFb+cSgnjeANUs2J3GexHXhlg55puw35T86iAm301B/6ErO7EZbrd1uRZVVn
NX44e2K4Af3mfPgbhAizsbPKKpYXCt+ug/kTY8bchGmGqsQ6ESFpnJvSXgfY3dlvl8YIwCfB3jCF
EI07b/PVD+5QgaByGZZkV1Bv+oncXQCza9J0MzDp14shJLzMAbrSmefjj3EvK6PgiVKqtJL9n9jV
vlg3W7XuR68A1TBuReDbpULuMz35LB6jOthylBqsIOJKK1okZBsKAlWP0kjOhgsQd7HlLljLhwdF
/ySnmPEMm1OQuNK4ZnKOPc5LvGJCJnoHK34sshjiC9qgAn6Gwic9wRuH1rWUf14P5GA9hJTVr4CS
3QwgXYqd1r5CB3JIL/CjpvYKlkiKbsx2LLinL2MQQZDQ27r2eV1wbyV9bXFv+xGvJKI8PuQmBlQ/
0cBGglV8N/V1KZitsvN/ZO3g8jp7gFYIRcSJu6dlxXEYu9Co5sGYTLoSZtBA5iKnJ65Rop/gmhCR
BcAJXjXClBDUtUdERfqnKzQgsngMu7VrmbCR5UsRVGjSCnnHr00tEMXo93Utr4XbKnjB7FuKH3ND
comdspMbV/1Ppk2pOb1n3AgAjhgN24RjmuCoaqp6Rp9ewWzDgmmolQvz4g6UQ3aG8XLRfH8GeP+Y
yzDXCJSxe/9rNlRu0xRD2rtXDFYlEBlbyjhBqA/qMyTADGBbso0wxw/5wHsLcOw/9f7Glir46a23
odbBe6369kR8k5xmSw+nI2qT56/kzvToEuezUAnYtZiTJjl5OJ/ooafkEK4Sj/2HyAtTXCciCGUJ
Ax+7p/XP5xbhOTZig8A+F36puHKQnmyxbTIYp1CYuNeKLdRn20pDbq1UHZpLDcKQ7m0LFwGIje/V
qK9CzFmsx4B332FGU75KwygWIQU0zlneVs/kTyS67oAbJ4Z0IFmQFdI61M9NC7D31OuA1Km9P74/
Ws2iSwUSRR4AS8f/6GiuBAOL1wYtMyxsWmRIIZEAWWS4B+g6+jGzVfPZDwkYqbeJ+zkEV4agmqkZ
cgTlC8KAyQOPuzOlRHPDPgYJ8wUxyIH03qLE03i0mbqZLreSOOu2t+ydcGJOsyG4iYhlnzJXeJj9
2afHyWYJSn74oTjVsXGF/IBG/0gk+MPBG6JcXrujOxoTx8IbtCFKVxx6huWZEQxB9zh8++W/+gkz
BjoVvpcxmd0Qg0yptqwZAWTyjrotyI/iZ/mzqrnykMN1RV7BKRQHGUkLerVnD1q9qCTHRb3WBnWN
OBBzJmTKOBoIoWKbL8SkjnpMlP4RbmMRW8PCvxeZ2NNkfhqAqbcP5+4PQEcI5TzSEKf6j7+Jx+Gn
CLJ+XEo0khymUl9hoRPYTXq/2Rw909ZhxCEpx3d4ivHUE0Lk0QaQLnHhIwuTcpEP2x+BqsrJ9YzC
JrZpVlXvru8Jg5HQhlUg/7jGHeCtUOMG33NOMo7Ip7Vi2NhFXfkOPZWGNzpuSGkUngvDK9mKd+/S
g/YyLsv/4pn/gD1YrcUsgunc374t3IDx+LJ6/clAZxs8uacZpTTCwr1kGNdAhbJKG+42RWZbzQz7
bt2eafOt2TiDCI0vVFnoW8DTqAVytRLsB6jMkQojNHtFr/qVUEMk2bg3ElFzrh+1McbpGQu2tXag
QqN+1tbbVxJnP6HHSdTEvlyGQvx2IFmvAMekZP/GupbAg5ju7IZ/EwYKwzr3sJrs192F7XzlJCJj
tl/jg66bzEIuPRvJw2x5qOwBQMQ3Grf1yuD4qzQbBewHS0Xi5yrvxvHhA27M5lA9ACPTkQ8ZF26M
gGecbCHQxkzq9CKYGwVMSSn99dQVZl3iywLQARgWVlSXSNsbgcQiQ3rbz7k3kLGKbqszCylx7eCv
YvNPIMVr45L6WNUsuc19L4NWE2uyafxpo8Qac4b5NVLkbEeSX6tXTtdDEvNwsF/I+KksadmMOEku
YjnWRLKBfKOJQ6ORMk04CkVnvrriyY0jzZhWskG0C3CLlf8UKorEO44UWXEYGCKBvDNChuK8dHo3
8bT0Wl4lM02FC1jaKRx4QRLJaGshGAC0jVLZR1n+mZ6y6GcMmr6UtjALGwe0Tpcv+LXQDOy9NElh
yRE3UNv2i3c4ta5jXM7C7vy5QrMbGCkTza0HbKdRTADyQHYvqMJa8T7IWru+uarGvfHFE02WPimw
lJxdDgw+v9y8Jekxyjrs+KpB2lpThPLf2Ifj7CcGbZj9LaB1ZysBStQPtWQthNY8Dzpf5BOP/rg5
LOPewPlju7YOIKQLAMUY9V6AqKIrNS5/7jxgfWWWWIZM8Br1Bz3DZNalKQB9Sc2TBl4fpkLqDMuj
OtAcw+3DTqNHo78ukIqdqbMPS04tBH+yhPedRUnOfKyDO+kexlBa73Np2Xc9mDZS0051PMl38pON
9CSqpdARvx4j43LJCeEX8LQpC0iRTiFRuSUh+F90HTTdbKqaDEVS3Fgx1LNaFTN48psmykJjFEn7
nQ+dxQ07zFSPN0yOap23MX31idr0KSWYrpZ1xdK8qJwl69x3E9UTTswQzdchzb8i0yFiwmGf0iNi
5jeAh9hzXIx0K6Djceeu3jfzMLfpaOdr9lkn1M7nFtGnGw0YcfvyAiJ1zH8NDnikGT5KeuGjBgPV
z6A94s6NCJsHwMhD7eGJ3Rthcqsv0SyTr6BzBVKiBdOGv2sP3YISz6q/uAOd4rZXKXvLobKmltMJ
FmdQHV1OhLAeJuoO2KrVt8VN0HBsf/TNx63qoZKlrt8uPB3NRVC6nBqWpk1mN65PIey1msAQuXp/
mXr3n0js3Y/7ch3rwMuZm1AFK+2/m/aP9CAPW7nOv8Fha3/Pt/S41E+vGp2eV4sNOsMd3ZJpAP/0
UnV5lf89FEpQZLFohyXUWLuYQXBRpiRi8eJl8KOdW9AA0mBWsUsXhrX/VF7G3yboJ9W9BqLqcmVF
4lRtJYVv1+/GvUAUxjzANr2dxD6D0TmPwxqR6Gnw4uCIi+iv+Wx8UU9oqOV08R4Tt2l9VvlgloPQ
8U/jGi12jUGOibEQ+YF/rwwKG3wN01KPl/Ksta2c1aU2g/OE72VNAZRQ2XpYK/SBb+O5OE4iUrm9
YwiRZplUo75W0BEHOfOT7HNPepyzff+MArL+AvEupDvQYs+E37rInwfQZqbCb4DaD73HZDlA9JvF
24w0PXGdtF+9ZCELAgQ+HST2iyKdwJViuwcquc0t77yvsDOHVtPwHT20vsq9WUtLem+VQsKcLK+c
iiVVxcrhqdaMHx0zTWlLYFfY5jH7RdwJ6Ab/1dMNygXTVz+ZT0Phjt8R+ZfqmT3xq3ZC0UfKas6t
mrz05wHfA9PiQzF0xCkhC5m3ofgdIjlJlWY3F/Z9HbwkNzNmOd32IfRVI2mB97Eq8WUBXawpSoIu
LYU4XA/2KxaXELj8MPX+pGWQO0u5tYcchR1zjggQtRlVyXBCb9wJmD/mJaoRvcS9p5OG+vI+Ouuu
yjMKVi462kIdgIPFPKCynpEPyGVc9J8RqrF5ouInbZfiDieEVB1qu1CQYwAKWcd8uGsW6PTJh/VH
R/acV0kBVw2xVlz3qn8GDIGp+CHpFAHxB8ie76X9zzgyoCZMW5qsCgVZq/0FsN6JPEpRTTQ1o0uI
/pzEP/qOrOPHrbvWNwZm1rqkgpoc0QDM7rDsZLU0eB851fMZGVsVQUg/cwT0M5GLHl+FoWAihVtT
jxRCfRVRCnh9bTeNQt0hhJUzn8UQlw1W4yIlVYvZOc87qVwencopafR4BLZum5mqzQHJoZ7Kq0M2
ycAsm/3roRMMJtRPZjQ3EBqXCMYpqN2qOT6yWUUmSxbONaNqn5L7IqhfSsLkIf/LBw+L8cKCsL1x
M5X4BNxqK5RmtlJ9y2RTY+/7nR4HNYbRBfE+LtWqLhjYGMPc7iRfF7IQW8NpbbM4P4oH/AcY471k
Ocxi9pSraJ5E/1wp7xUh5BaNbaDkfdy7UYwCjHt66csG2vb2D9MxXItXv6eMwP6ko8IaDf7lUppf
rDORbYAq0v2c2s+wrEKrb+x5G8DppMa+h+KPoOTD1AA8v6orymcGqKRnP6U/RkLcFILe30UHF/oX
NheBqiU2WkP6UoiBaWfLIiRydQY0mGOqKW4Z5MdbG6+L4PuRiAT6xOdcrFgmi04ulvkc4YfCdTY0
nKjRrkAr+GCXzyq1sRLPhRUrEOjwYxruRc40iir+4LSL+sRq80AIJtEo2t9/fCaqFiONnZY1IyOf
QoijT5nC6UUvbVvDcLEn0NA11yYLZ5g3keh0G7rYWoTnBGzIqy25DVj1UCxqjmAb4isFt44rxcdS
s+vbypIEpsU7pXF/YVYOQ8rRa+S9NDfqWyGtqAPA6jfYDPsiO9OuelLrkBmEo3SnTZB89zODkhqy
FYIRG61MEaBJl9yMmAH3oIIk7wXPhA4FZls+bZbd7QspkJ9U6kfpkd0NU+WWAy+PXhCeYUEcmaZZ
IRBTaI8NWEodNqWA2vZNW2cAvFFKdWftuOpxZpPAWThHcGoyZgIDbAcKCM2o+6Vd7UHubR5iGU7w
2QH5Ocm4gNH1dbXM+BtfLcWaxwdUGHvBq7uslQQ/2/vyZs0OLhFtIdEhdc4Qj9ge18dBHvSNSfyB
+f8VnAGqE63kFCSep/qRIoBKU6YMxL7PX3fQs4xWkmeJXzdZt0LEDbDo2W0C4cZfQaegfMdDCHH6
uqkB1/LJ+0qT/XSq82UYCpz4TWW6Cw8Naeo2vsFwWp/sYcDGqY+iUnU6Brcr5YnSsmrWXv+8YW3v
fl7GLKWzrKCHQtZPrSaQNej/HzDpo2VNFo/sK3PNXfWJ0CAdkv1rNM7G/Km0w2F+A37bq7ccDBBb
TaN+7Eouuqb1r2ov+HpG1bJijR8uwyPSEDBez+1eMqSrzxYsIQmAC4hkys7vc6p2vyq/X9eo+w5k
xcmnQntp4Y/+XNYMETDbXNgDQ2VS0qCiCJUED3PuY8HVDImv/E66u7+/UxI5OZBtEDGgzJJoyR9J
PbETiUnIaue72WemPXu0ZqWdxKzh/QpKxAC7T+U3Cv60g6gI27IR1XehKvIDXF9+nKxejIHzxLOv
Q5Dx3Zv7oMj75fTuye+y9gAMEQ4uJVS7mSqVFXreF13MZMrQ8/+EQUbFpmewuoe1b/c17u7MoAsR
I43MuUJzKIMBMAmEIdADakauAG7fEP66Rk+XHvHXvByZ5UyZ+Q6RYEQzfDhpyjubYXglomlKOy4a
U7/foiegAFI6vMng5TDiYaR0UM6BqAP7cO2HRF4Vk0nim9VsQqg3ILjJUCQO6ZC6wDtUtWl2DonQ
SbXLyLCAUJx+iZWjq9tKDk6QbCsZEJBu86kE5dyaiiDUcxGzAPtsAR10vxWJwHpy/yE4Yy3GJr9Z
x7vZRzBlvKS9Pc1JC9ES6Bul4QhhqFb90/5K6SUWylNKEApYstAgBgvQc0dZuixAD8vv59jPKm83
rreCnAbfnoffi0B4VSi2DaS6B5aS2l+a/papA9TEeH9vyb31GOeZum0Y8sy1+Jv4s5nbgVz+C1OS
VJy32Q7xi7sLuLGxoSOP/UiX0ayYEd9GkwxIjHzy8iujI2JxNsxUfNYdKHNxrxDXYzwBdjt/Dxkj
v9YPxtXUsL/dPKpF7buRWC5r3LqOp2JSyrLzA80C6OnK273yBA9JKT884ouAijoBVeqJsHEzyw0k
38hC9H0gq3OLe3rI4T83txy90WCZoU2xuOJE7+5Ld14YBhuXkTm+rSv1Q3PjQ+TjPEZ9/9sosuL/
Mwey2+pu+D+NoDi5XMwzv2jHLxqI6Qf2AX967SpewY1Mz3R5iofNHkCefFh5NaHvU9wXG31PE+yI
WznlpMfQdkEqnJmFRliFN1PkjUylmdu2Vnv+WsePqLbPKJbnVbI4RoG8/6r4ux6msg3FmQA4yYLC
0fn1/91jJcb5xagp//ezTLxLNU0pCH2Pafy+88L9R2uEx/OaiEi4DTNa430VavQPvFv4S+Iz+9T+
Q+JHlF4BV5SIp+4JydqyEFzRjCe90u5r4no9Jp/S7ZxpHrS19wDxDkOsiEn7JgEw9qtjkw9VI4C/
7aMSvCz/ZM5PYhhZ3TPzvJ3xTnfTBFoJ1xjxrLRNDMaLCNScaF8WcnGW0tjqxVyalq2hSePZQy42
XSm9bb964VicKKpnCQhUlaEHzhXV4gpVDw5utZcjtzQnwaKeZw3LN/xHW5sX8uu+hGMDkrLxO3f+
yAcqRK9b3ze6jGLpZpHrLgFkVunHOf3DunnGXjbtYAfkjlgRQAOfeE6xE9TRxud8pR0r22VZoFmJ
VukEY479WMbNczrykJYqx6KuwAZj9+oVEmTe7cEIVzzgHo1gN3uLXIc0YKbADq5fUtIr8x6vZIBV
n9eaYF0v6QvPR8KasVasVStbS7VyjnrQDGgaOvKNummSzKAU34s8Izk/B8MKM3OjlC4/Mx3Fu4WI
pe+f+xFcfvOeVHRMd379f6kPduAuQEMZo1BqEtYEJ6JZ4nmgyKYDpWU4H3nSbxibAI0NTdM8ghIs
beSw+n5U2jL5LrT0MDpbhmwEGbfBsiv0RIflUFMFusSrUUEu8nzF8MRrZuhzCVuV5tvq2+ZbIwdk
WV8HGd3PD1bASCGcEzWSus+3D1mwxiTefZnGh3cyK6K6zy3iXTA8n0yWOeGl19mXAwixxfRpszMQ
Q2OYIjOOHxhFSmTqfPY1Kuqnwl7Jqu8ju+sLpRxrdhKVE7lqruS1stpk5vrqmo550fRQyTbX0cK7
lUa8fGUNWapef5IKQMZK//dpBqXOXpzXGvwnghmn8uxaHj8HtUB92HsG/i9G8fURwn7maABzQ53m
RoDI2dBkrYYjGBQpjg+bCm1r8T2XE1/QpVHV5/pydWKyOXxIVZRTtH51Cj/aYStaitE3fcnYquPx
9ijK8+Lxzemo+5vjnnCKhk517HjiJNXKFdY2swRdYMwXBrB4oHNh/ZHzU7Tm4vPQDhaFbHHjss/2
ywJcIYcqOa0GkwCTMSX0HmBlCvnm99zxncsFgFBg5okM0riXhoq9ITW7vCtUURPpK+TVDkkILQjr
h1DBNhprBgQJlwFPRURyvG63i0WZ1F/MQ4+4oyfGzq04zq4676KIDThOEdDmPgK4XUQUaWxFatkQ
tsSCbaGnui3XugtIBUyhOV+D0oEOdZ0MKPV2u0LJGbdBZiLdnGmpfOWl8RhM5MGaWsV+ZNl0rCbV
9KUX3IOCenYzZFVvQPugIKvWGGLBUMYmGpgUGlT9RIdI1Uyy45NfBjUgpOhnYHaFsb5gYQsnY/ma
0aRy401ZUgwXrf3bS0I6wnnARFOf/RhId/piIOdw2vYqO6ycCTztXWIzcw/C7SHJp3w1fskLBR2L
kmU1PbQaU5snm/w/Q6eFtTbAUAV9maAiTKfeJPkbtOqvqS5mp4q7GMWSqU8JT3oWE/FukO7PzvHH
vt6kXUhcj7njCqBuBzgyOYAT7br8QVg+HtJqE1XPJ11iVB/hcL4PcOdddGal8x7KFPPXwTamxKbB
a39PNf9mhcLx5pAmWnX6C4MiGZ+E/OHsk0+MmoYgHju+s7pb0UJqMJJoGP2sYK6FZf/PpcPztfeM
YPZw8SrzWtd5reyb+anVFhszSoh8kRfSphcVzD9RlAfgBxxRg2a1ffibJ70DZNMWKOqGR1T4JU7+
q4PjfMyqv5lTCiVu8LQZ6MdHDgjRoU+k91yrz46Bg2nJeM706t4A+fsfq5qkppFMuDUvp3RjQGLQ
bt9MSWVjz+1fqnlaY7OwsX02EqBmrAOpaxPZhyIlD86Ix0hPLixJ+1VlGeh0WmM1oS0VLRDWNeig
Glz3UvHOnORz+2GmWH8P1uy0gtiPLHt1Q8LDNG+04oDfDGFoG6xdL/I5dIfER/OAlCjvRsV+AT13
mskeL4cFlYL3Br7L+01ZBftk5Ya/biZ7YEXkgiZirO/HTzEAdJh3scU9bEBVt5JuCDuJxSQxRZFF
/IQM7/opSCBPeJP3V93BXPIh7/MgiUzB7wK4kmyHQ4sXJiodYsBB36LybFNHZCLxeprfukDUQcyb
70vzfbqeedpCL3ls0Cq2OwxEd4xch0TLranlNXtFO5M6KlEgL4U2nUUtCnUklZ6OMl0fg/5wXJ0W
qBJUVriEJ5N1HJXU4lb3cWUMUVAltwv8MpE/ZbhISIXsB3Vd43NzC8TO/9JbEq8Zt9uRskhOWwuV
to0IhdSEuiCKy/PrH3aBgbza0r2QP7yIJIaHJsjzA7PmySQRrRIlMuV/0PTTZXEZ21uz3nhqNKnv
JwXTwxEzaoPfN2MA/zcc6mVxWob5pzUr7wVNBmgitbvHyY7P5b18uQutJEYHmAWeaZBB8pivV2iU
V9j2jPSL5KlwXZNkZ0Oi63NyEH9xaKhdILJ+FrtBwrweKWtVccBeQJnV5Foq71lfARMzGyMFQ2RE
OX91h/FLOSQuNB5zRdy6A7W/ucISVBNhchWaK7zA14LdW5MfcD7KvRntnA+1cac8Zr46cr9kznwd
ShdV792vfyqE+7Y9SHDaJ7YwrEeK1r/CdP0NAX/8UswIs1r75oI04Dz1xTAEc3OCwqb47xvdaDYw
RkUdOddD+7ggU5QdYaoK27lDtYtUt14k3iQmVvIyBQdSxk04jX9pjISW/iI+LKi47ZLeQ+WNRg2D
ImaylcbG6i+3t4W9jLljXKrRQmjJSk7HK+JsjcadmtR/KskZ+Yjoitw5Ue7ES8RJI/k2LOAsSmfa
NyJva5oNdC7Fo/PhPADS7D4mBKDnSM5EZvvDm9mPDKy2OINiVm7SgawaEq4WjZ+sC7+7rP3mhr+9
mUqFfdrGrBsDrKtG2K6YxQDFxieqVZgdPVUi36g/j9f/45ZdnAyW1noWeBYEXicV+NKtYFiKbF1v
w0L8IxTK9FKGyX7+4aJpFBIeSqM3A2MyI0CjSJLZo9j39DtWGS/8srk6lX6joZ4xdHKnYYUuBNsC
G6yqLo3UzxJJ4uLzPOEcg/muYm4GgKS+JpmMrWVdX5Bs1B9U4ArUEaOYlJz99KJOIWGmP9ieuGFr
H3fiww2iB8OA+gMEHZSFwBQjTtax61dKVplBfQuvf+mjxDepupeNPWMLSzcIvDBpiHP1yqXlNYN1
GJDM3a6U5/jHco7v5uqk+EQftkDPd4s9tS6E9XAw0EB2/vCbCH/1VzCD0MzLxaoMuAr3A5npk6A0
5veVExLJcxoq6KxZqMfTyT0+4xukcGlG9AS6Ot4S+ikiIRuCU2lY547KlrAdexkssCtp0l7RAVLl
FBXeePHuEq6tZ7iC9ErpjeJCjvdwQRWzZOw/3RCMIsjOZCMT/oYeDcPXa/8PK66Yk5b2mpzUZti3
cYU+49cwMrl/g/4KtusJ3sqbkwZEKJnPf/jenZr7HtpLOYJmrcXjnKfNU2hz/1CkHvMYrzrLe14u
P8v6I8CEojzqKvPZtTnIoIIuHEsDxTNt9FtbxTyneUMWqE2S6TcCZQGCUjC6xfYBn7bsgR4/coMJ
1dojDQNn7HCbfyHEGJmAuYY7aSe8boUluYGd4QTPj6b5Nl1/PYdgcVCbXfkhWfSWnlWum7fqyT9q
sms2v/H5Y1vSviQ/jVIcwGWZY17ea1L2J9gyrMHf/eptlXLJ7E1jpU50WQx6bj9jLoL6QgLZhs6Q
BVJ/LNsPmqqtXDia/dUofEA6sEkjqHHBdMeMdw53OK3rNNpApvJV4qHUnG36tIEv2RAS9PXqZPX5
MPX6iWvbmzrvc7LM1V+mPWuFMaCT1p7pBeg54UpGxR273lhFs7TplC1QNJPki2pthMRgezBmfiIv
WUa+Z2ExpZtVwXkb1vsRK+VwdIwryLeTjKRd8WZdofTKtB92715tOGl2eSRBoxWv4twlp3A7EA9c
FVSldPabrTBLu9DslYB3vNsImG0DCbum+ww+DsvkNT8Mz2tF6YOZm67T+S/f/pqeY7JAX92E3NU3
XTT5hLYbfqRDErkoJT0ae616oB7Tz+tfGHkZ2WSCOEcKViCE5EXE+YLdsxCSgRAaSlMKJaMFgWwP
9chP/YU65hstgrWT+Vg1TfBMuGjtZNl5AlFujiaA/+yLz/zxyZMPsPYMglA/shF8cvLZKJhePhAG
26bRv3IzhHOBv92x3xQ6baQXk4QC8HE7l3Dmh0Vxq1wOZnr2rzabpK+rWPfFLY9UziAAoZD/Sfe4
GPnetg2bGRiucTWS9uGNtCeQeRR3rA+zq8vrbAMDpRTxEP7WhkJduSTzFhjNekiMHdJZbR2Qt3bo
pCDeNtPpx+Q0yEgAvaXBi/2enUmKCgDqTTWLVsb8a1bzMkzM4V5pldc5hJPhgG9XtrFcNfbzS0Zs
eWJCcilFui2FaDDAOMQLkXri7U+CGlUPri5lJXfViGcAudzEySI6aQhNp7ijXJr7ti6sgggjCkYJ
cfBGgX+klUH3Q79NHEMUX0hLxT4z4ZFs2tRICQmBatK5iET9+TAnBvSPDLE448ltKWTTG9tkDi6W
r7ogPZErzGWFJ8s+Ks/+oRcaPJjFfZ+FMXGToniPC9VOwxDP1ObfHyODgucr7VVHPF23aBE+wpxs
xuCPGapirVIEG/c2SyCw85gEiElPBX0TMTpjMa9qVyK30gMsrjXLL35PaM7FbQ732xUdZwFrhvOF
jLahKda4VbJgbiZS0TZtvwBNU6gt+d6kvkww3aL0gtYTT+SMjageRV6Ko2fiEA9K1cOBIXnim7qe
u98u3+iDKzQDkY9c+wfDHJ0g16QLZ/WjT0QtX/1YfAdq6OqJ1UUQ63vyT/1rlWuE64vzuHkZXa8t
UR+c1KP8Dvsng0+ISicNYZi+RLAhHXhHgOWFsbYKjNhoAEAvQ1NCsGgh3+wVpVSVgqCO+tdP29Sj
58znQox2xY9MthAz9ayXqGWTcu03spYrIyLwKnHSdSJ8luC0spcwiHtp1VfCERqHyJ+5ZnBwLzic
RdFLoDEPAJvAz4AyFXrg4aROjopRkCjtK/5Gb2myth8Bonm/M/Ob0FJiBu8Yx8lPXSxp0417CpWl
GrLbNmfXWX+iGm11GGZ8e8/h3jnmPagkufN4QCO1NNdPFJnG8+VVFQCkeDxkrgp+pxsdj+bRO0GF
/6VDC+ki5uBZmVGgEh5xDuOHTn3alilGlEe2DLYCANNNPbJUUI5tiivXsiI9VG2cqfZUt91tOMFh
3TiH4uhB1Z4hl1TEurbQMJUJHsvSij6WjKJIUGt37fZoAi6L9mgSaQ6OfYbTqHNYhE2x9zaY3sH1
JBvDuUi9U+kCOeHyWrc/6OjXLtCinuZBz/aUjajSlJSk2pf5iI1WGg532tvHo5elIzQoLE+jVOYz
l+EbUGwp4PBG1PYbUtVSP2TtiEaF/4VENw92gJPgECtows0qi41SuOzAg51HwkX3+sOC6+yEvehD
Lg5DNrTGBUq9uwNiORSp8FDXFX3sOcyb1VhrSndOLPx+1B4HPxpAHjrRqTPV68RoEpSG/g8HWuLI
Vt6DcUTrsLLiVAhFiilwvmYcGKxhwmCEDg7EUcIZENEZi/hoGo4XMJMXY7n0OTyO6U3Q63xJbP4G
WifLbAfSr9uOIXT4hXnviYfyn0HKFRw3U+he2jzAVM9mi4JQSt6fjIgls9z3sYo71uHExgEe4cJv
TbpfGKP9vUNYkq3958UxoQ0QTxvT472Vz1p16BE6F8hLRgqKxo9EaGL7/kKhVYcQseAs6S9lAhuB
W4u/1gzaAke4if/fQLg2edmu27Y+pAOIsw2rjX5wPYClGFBN1FKed+0bZnUBgc5oXrBx8PeLj+u5
7gnOrMEvpVb3KS3WLmEbQzEbFbC7MwbEZKadBfo40cJjP/f1rCk41de9K/z3HG+LLHry609ZJPcx
vEJdZ1yIZxWo4EHe0mzbiA354jJ0BvRyehsPhUwJjJrnlCCYRTcRIBT/kj1UTVgak/+VGCkqa4r9
n1ZdJjBfL4ESUFa4lB20d3NN47Jo21E+s9sMJFtIofeRR1s8FJDKG8mERu5ST0ii3+S/CLhsTsFe
Ci9a2pFul9Jy3SWwEWmP6wr4PDGXMR5diiw/sSWNthkU8BZXfXR9wmOTCqihYKeGLk8+FKsoL2SJ
/V5HuNE38dGzDSU/BI8hnGE7kuP/JpLgx8KlFg6RYZkzasK3jYFjwkuPLUhhCBJpInUsAmhrVkkV
6jCgju5chHphpBftAC022uBxpcA4MMrNEpOL9l3bGftKkrsRzyq/aE6bL8fVdR0+as3zPaERcoCg
U6CpCDhce8t9x4ywsoakTEGuEJ6mCEr+Noyl1bh22oPVf6pXDf8pWiVIy+NVmtWK2tzq/RVUndPj
elcD+Yt+R26mCkgygaR2VcHd29YR8p7y5zzbc8gXAxEDsWlQRjFiXHsPtoqEtf6OQXKayW512Yoy
1AdWYlk2zh2O0X8SMhv8czAoRD+aPnhAmiMgCCpfgwrsFItro9lxix9nBx4RBVCMMZ3Yb4ExYsW3
myXyJnReLVC59oZwYvUUdFesOLgj4dtZNfkPcU4yvPkcOfCD/Cd/ifvbpJes9TDt6keY2n3XaegG
o82N+LpfL6SHLQtPuwpu7I/txKLptNQBgii6FD00OJfdvPU5PogAWXFEC/P3lD70s3PKFiNwzUTg
6cfI+Cm1RO4cuzfWLN79pGFoiyZ+wFuNkCK2OLvQ+WuE01vjn/MmFfvvD/T8yC5TuJ5HBjpsoaPR
spHAx4BdA15xaQ4prGq0nDUjEBEvakkZwHqKopXVd2mop2sdOGA3oEUZrSV9N8DQPPtHLR3BaMpg
+w7U8FVws3F/EQGaoFUQekVbgnvKkGyuPR2EVFQJzR+yaL7kaG/97lPUckJxUqlH6S8QxG3m3wi/
BHLrPb5ZYPuZBFDIt+Rpq+AmNcbegmxySXGRsn9HeTofAlhuFLSEBRUsdfi/GSZAZN21R4xrjcaO
I85rzyIKR67UWlVBXvYPO0J9UhocjMAnPcRxF62Vf0o1bv7ye0d9ea/aekBYADJMuBeq4dZzwI7C
+7YuubzC+CmNV+E13bNK5+wzm3vEO6b1dUogBBdtX4b5uOilXR2i/+1pRTWioiU1mYs8aXdsSeod
6frDCPeqaCZOZ3RIn2Z1Ax+xVrnjXUdmeRH2OpSUtaGuFEjtvym0nMBZqhPLJAvyDndurOXmpzBZ
1cUtWeCn3OVbB7CP0wmolbM5lLEsqofeGoPVNgLrviSBeViBQFIgn/61sC+LMLqEqABWJmKCUyIl
SjCqkBQg+xPmKTv7DFnptcRXstsi2oe905opGZn3i3dNNavPP+8kkaiH7WzK9u8WLN1Sew1xVPpD
QlJV/AT7ub57egkgh1bcQUtiLjhcTkQ0PL6+IAVR5fHdwKiiyldfhdO9r+/PX1NR2hpZmHbKHcf8
qC3EjzdOXxXSAYLoqZx7u2IwBuX07kTK5jA0CYK2lczqd30dQrT3mbvgQfc91ls7YI2f9odsFrkY
sixgMITv8HxjpMixQNcJ7/bDUJMCIwlHixBF/eg9h6D4gG+w32HPU3ll80/1wWBao6/VbZiO/rrc
6bHRzAE5QbHiY/Gd4s6UVfyTsDL6XRwxX8sbZK8SOdEr8PsiaDXP7g6tEL4/LDyIeG6sNRtj9XVb
ow90SsS7zdxuVVivrHQ1mVzmCFlJdgibZg20IUmsNA/Nx/bUiRwG+7KY91IiNZp8T4snLWEfwEHS
+R081Pe3YUf0X6lV7FIpMA1hlBc8/mfDJXFe7wavztsNnT80eSJVr6jl/rnrVupbi9sqarkdh0UA
IWEqj8/z7/yt2CZGqlBlYLYJH3a8dK6RSpr5tkiyEI44fWTp/HNSGbQDxTu6d8dn0YPh/r4DE2Fv
TnWKsNfeZOFKOa33UQaTqolde8Zy52kBM+VGKwbOfWtP7PR/fPRzfPRrNzxB5FvUQcN3hNuHFZ7g
j8L0cO3rBDhYv9GfLG6lc1caCk+CBDfk7dptnkFXNC/jr7b+DySLixWl0zIVklCitBmX/aeh3CnB
OURcQamiScnTYFqmFtIjDEmO9/Eh2Wcp9UBSvNCTFTP6R1ZK6vTMrTOgnEoxgiIRXcBtC2gHXhtD
4dFPpRww1NosQ4lV/zNvyyYFZ30Xm1+pqqQVrBLDr+ql0JABvxh//KwlxsbGNBk/+DkcGEPlXjrp
63NEpeLRuIQFbNTfJxLojJKpWiMxPkkQpO3viQ9+yhDIcojYeWy0mloNrvsxiKREO+oVr+O1ucye
/y/nycia400n/2aGR50mA+TictSLqqQ2auaPuVbZKiI0JN1TjN5ipC5kIh+AN1SCfKCHyQa0m9R7
VZcKHQxFQoag27OFEAj7WuJI8qXWemHDWdyycxOE3MMyZrsNc5rJI3fr7FMcU3+wUfdbsJAI/iNC
zvB8eXVtWeN5VQkWcw4qck/byPROOcN7aRCVfzqL9V1fpuxfQVJgWcM25ayNkjonO0PunIV1qC/U
MMH6VxjyG2gdaq6rXQ2bw4c8TcxPiPplhS+mdSAgTJKdvr6zClqfNCjDmpkLwNz2eZw8ue7peihV
z3BoEKg23UHZWwDkHu4Yq/E4/TR4GbXXsX9I5Omk2NARICeWKca1QqRMBj9gDy4Szs4GSWr57ZdR
johX/WThuZd/tFztmrOGhZx4A6dO9/t4vEihkBZPt59xFAuGd5i4ua5JwADkQNg4TPl0k3VMesWg
dlseZweoR2bwrHdMcG2xyvJBYGcCquq+ZXaP+RZZ7JdYaPylXJO9Q9OcY+qLpHilDcdnZOXf5TuX
11J/6qbLwhrvGieAxKNHaKjcHa2rzm5pJAq9sOUitFUFF+a9TxfkdESich+swgI+Qh3fa7/zVoMh
+p/bLY0LbnaVpvq4z1r/vS6tdxEGRqtzmsp1CNRBDBNEC2UdaOYz7YRqvEmJwq1B+t5zjvsqn5vj
em7qua/IL92/COG+oOK9Z9xnhPfomcnEtlIn5UoPl6N5Nde3uD/TJ2A+URaPL4JfjMoQFRh1rey4
fd9NrK1LeLAhU8Oc0UUkKPDqpBuY/vfXyaojTKt8LUe9j2rRYUNyyTtbSPrdh1cjr4wOIbPNFUvQ
RiwM5LxZetXoG34MfbZYmfv1k8NfWvfeQ95LGdW1aG3FfqR3+KVr+xX/obeII6fEbcbeht2xWBcu
Up34/Cnjp0SAzGEQUtSs03p9lNhM/F0bLxpGTjQb1neWyuKsu9qIQVAO+eG7QvUvcHs/LF4PUZyX
fd6l0ThBxUrxa05nRBYC3vWcvuA7rcPt9CB94yK6Ao0+jW9QtMq7PwywMBpfCbDC7tWNQ9GI4hdM
YlJCwcYj3eIK0+EkpsU/ygThEXVMi/tlh9iWW+ullN/o7e2CCxz3ZtFG9Abgu6rS5siDnRxudIa9
yyFYv3Rmwu7m5IZ7G85dZC4wYjP8mOg8h2LG2gM4UZ4LSKJTj6ULzFqekdXpB0Zov8DI5ycwcY+p
KmjLeiBeGIyEni50MjAyUuN/6mH+UASYR7P8KtOp0K74cTsxzNizP6ZBUPqcbLaxQrrVl6wQ7dw1
9B4XqNPpifcNrssA4tuVCyalc8wjiitxzZdA6iFVHW+9AisfT9RbuiblxCW3L1d3U8hzeiHgwR3i
X8JhF5TQ/dEgTT8E2DrXDVFdbglGXGE2DdAE8AXC5YGhf0wcz9aA/jH0y5LCpV9l12aLpCsbl1iX
aP78uWpP0nBSQt7t4AFaM433ezVgbSLPxk/10edi2xz4+H0K1CJPsD2ciydwZC+4T11T9VI1QpOK
pdoAW/+ULD8YuCicrgBqFLYCg7+SCbxw9NaL4a1OhJtpL3vux0p0fbtJvtJTAZ25aM4fmPStb+I8
S/LlgUZAwKsE/6FRRLIepVN+uCp3LGxCaeyjFcG00QHwhfy+tGVC82bgKLcY456PZXHxmjTWSmqb
5OMVOptOdTIJRY5Al0gLpyF97tKaGV3E7LAyAPdNf7vlrC/9f21Z+ywU2BfXrqTi4gIEqXJJ19M7
yQ8BRPmxdHpOfuMKw4zxcKmjKfuykOUCcCFqBf7a9DkYhfLgelmti+n/z+B/AxI2bTC8rLDrIMQP
w9wmYjUjTXUNhR98t4+c4SOF2oM9obW11cVwMFmg0TE74VsBv+3WfJ+U4Ih5W5c2oW4AQpF94vmj
7Q2P93UmqK3NToy7lLyemrqNIFDfKYer9oo0r39bNdOEHJmU5KBrgg82bASFSJk1NtvsrIfEYVFM
vnA1+s0vUZ74D5ngL9fR3i5PwUAKyI3HM+26QYiVKOi3s3NwHIxmhA985bZY70KhYRnuIRQHs5LQ
csirBEUJHcXI3avyOSkNcLIcDbR60usuwrGbIV3/hxXqBHbBp0Md+75bfw1eaSo7XEjJuWhrJ1Ug
SVIk5v5d6cyn7uWq+HE3+s5THDq7lKgvQn9UPOAnWQBzOo3AX9fSsFDrfDPEezaxScqYrrYJABes
zuXkI6eSh53Xjdvb5dDvBvaD/V5LW45eJDqLMuziV0kGIN1mJcFnrb6e1Lmtlf6sASnLUUpKs78f
IhXfjVFEodJH4gF+FfLQgQxHUjpgNg66gLsmMIjX09EfscUYZC90KxdOtQ1SGwG1tglJcBBTIrSl
3o13v/3LSdaibFY/vcPGD8A9XLCUvAvWMvZDDuzkrtE60/ZhRrz80mxW0gdlEiaNJjWcHtpcirHe
J2WcWab8oUaufdh88RyK1Qon+shwNHOoGzpCVX3jeAovr7R1Q//nQB9XEi9jJHTUvBRVFQthOQw9
gVgqyREs4IvxPraa6ngM6zNDxEGSDkxtgTwLWKKINw+mjgPAkIE5F3dslYDCMuHYHUYUYlff0r41
/5ETtEvsCqSUmsB69NiyN7tAqwg0py6V5bHyPVd5mijLoGIZ4FH6JmHSbSEKyp1kGW6GfykgK/T7
rSYqDHQalr6yME6QHAsl9ymb+ab1RTSXe/Bn3k+zZ1mkYabDarNlr8/wOiCMPhcDEBeOJOYf/9L5
8IqA5tjfdu3OvNt7aWT7aGgEYh41JC5Yo/ucUvyn5OR45wAlHyzp5wfCKRUHSyq5dTDR+J9yGbNd
CjAA7AlFdBre+PVrO3H4kWUASfrk2s8b3O+TI3ZvAhndQ/2aGDY0ZCgcZcUFjUZ9nynBW12A/G6/
hFGqFWVqMhUtyT1PY56QTDWfDNUK5zL0iWzeJFLbf8tfBclIC5auMh5/rmXCvhAmA4UBv32BpOMR
MHRH+2PiqCaUbVpuLANidQNKABwLakgxuEfBQXDOxA1x07BdoWjNv7wa6ZY+w28XziBDIZ5ZxSEg
lF5PayqinpZAHIk2hxFcmx0Rh6DunMWvBd/J7eoGeVJjAtuaqnEsku//wINP1p9721fO10hyyRSu
ARonWCI399JS9b51rwlFMwF2JSVF8tTFsa4jg++bPvBQDWzJw2Lcw9dHqkfYeGz82CwPNXoidgZ9
Dodz9wilGUDgy6PePmrrWjt+uQx2NGQnT5ZqEbvubcclZ27Gf229rpnqa4DnNkOkXfuOdYw+vHwi
z/fhc35bOexEcaIvtBsfvW5EmfHevwxQIo/rmNjYvEMexs/6DXkcIbOqEnC5Eh1Z5oPWqBLKR5KW
306Yr3by3NKIhPFxENMJVqaFsM+BSe8+xstsH32mdfdhuKl/o2cuGkzRRNC9ne7OidPFdko3mRW1
Ih7fBmMstZWtku+WXkKUAI3HQnk3ykJfnPOPK28Pr1dEFfWjc2DHYoXCZO4ctQ/1Ls3zy6FnWh9m
iA8epb/Nh4X0BEQ1zjDg99ZRvu/sdc3HuySOGQDF2Dg+BYjgXQAnIGNzcIfwx+aFP+8jREx89dUU
I+kJ3XUte/Qttl5NYcYrkxQk3JY+8698AnSji3Nk5fZzCTeWk1pBXQl2+4Fz3WQZvjC7nd+o8c1Q
FaBzV1xX7qwBfw74I9NG4VGWspN7+sV45I/21ODwxUd9lBHpA0ag9byUZsu4j9nsScEHf9EIDuT3
znkBDBOFNi3/sR6Cu4jqKFsuY2LcK0dq7ucLop3hbOrCNFDGRB4E7jgaG2d1tWj3ej3eH3t78ta8
qggnSBDUhKF9GWPS7sgOa2wLARmGi8syYcTU7uvJhBm7xvJJ9haRredtqkp6QCj6OXBU6u5XWvCV
/Ele7bbHYFDmwjLQPADtEMD19+c8UQS80iLuHTLGaxcYK2TZZZgVAdbomXdPjq31c637jXEBQBk4
67olnojiYlsfGkFO7oGZYWfU1AUaO1UNKNF2GqzTiI8tFL7CGkvOHKD5xbhsVu7Jc6HLaQPC0sic
froxeNu3xvWS4ufpSLex0v3rNUwQ1e1laFMFmOI3eBJHII73M1SnHh0AgdkugQf0crsjE0MHOexS
M1p/c+yKw6O18WuuSzrVmjg2CklAfxHP8UBhZ44fPWIOODv4HjRJYaaZOFJ0umc3M+qv7V+sE3ll
/fRkkTPj847fRl2d8XHllKsJD4NdZuM+yVBZxJUSCUFv8dKCQaITHsRJjkS5o39ZnAC0ZXdZRl7l
V5V2ICwiqVB+axxaTOYt7fYsX9yL9YaFLq7hLv1l8ecU0O8hGhd/JhfvguF++IN7trFlJAFCsI81
mxZcKvIe4AFoJYyFZZ3MCLcc3HMQVfQZmqlzHS8oV7cTrO/xaDxBMpVTgFdYmB8RUEfn7/UffPf8
7dfrYIWQYaCfeOQQs2hB5b9W6QOTk7vTKIsCG/LaRM8NPOOhasTdTzZmo1E5c2Zn9EkbhpQ88laJ
GesWQh70fuS7S6g6u4R8rpLykn5P05zIg/QFutymCIvp1fUxZFg8FFghbfUHRQmyovAT7F/McCTm
c9Ra9OyJP1wjoowH79Jx92xHqNhNmxGj0xYBCrmGM0v2rCOvSrL707WLMC8/AwX+9GVU93IBm375
1SlvaFWzT/x8pavFGUeAeyP6H1ns68Cu5dRvWd+of9gxZUQPpTO7TL14soclvl+oknZEc0yebvSQ
8dvkOC6LC9iDvNr4/GJQzzIXLd1+yiVGxAFDkpjYfOvuRU7fXheJoM+qANdaWgxSlveDiCHHEry7
HTvtLZ/lT/bgbSnS9pd35DWaHddNTfwomIuTMaiHKK4cay/uhIZXufN2KwohDvhvaxA954go8Bro
iBEs43aLCKSN5QcpBvZetyT5ZcoY+rXah2tNwIH9m+RF0ZEdnXqvzZd3mo0Fp6DCrQbxe1bnjH8u
WyopgvLHvaRiY0ZeltGXtZkJeuJ5+G3Iv5UBB8+EmQ854cotao2DzdRWms5bK6VesSQ8Fsfj4Nzu
Ha23cvSF+YaP8cpyjwybWSmplf5z5qhHLZ9xP3qPRfdlxqdNBaWGqm8LMff/me9ZwaSSuWkG3mGd
cq2gqdfSoqQhj/CvtR4qOtbWQYyNscHCLqsPTQdFrlavvyH57Rmzp0V5DKoPekbncgdwHjn3ORSV
mwDsmNibsoXUnSsj5KFzxAvxPzcirk3kBTRs++2SKfEOmj3DF9vpBGL/T0TYT3N53/0WLtNc/KBl
0CZSytzkVq5lJp1f0TFl9XHwVmo+u0EC59sA4tZPe0P7woyXKLbwiacTDOGX/skVLiGPljxZ35if
5ZzhlL9gMKr7U92W2JkbEyXWW2hcCbhjIIYrWQy8Go9fqkvN7f79ZidjamclaG1y4ukGkzUpkxlo
PrhuwC40Utk5+iVLYlfO9duzi8+X5GMOHq1d5vTEPZmq/N8ZoBN3uJhVRjyUPDQ+4wnSX/jpyHJj
bAD2IjcIzQZsoGBWnxRPYkM1jeb+GyWyBnGeTtINZSPRMGpojW3MvBm+fSSoAEEZgohnn2syRyW9
G2HNJVyUYkQs7WLKCOu7DTNN6kjdv5DT3yCv/1pWK9rhYlcPHOkPD1KfjfGcuPo1/QmE0PLNH84+
BI5zRPW7WKExW//uP4B+05CPc17vxQ5T+1aG+JxR9Zqng0cEJEv9dG0xZBYa89RMa1FWrtHjBM5g
doI2QPrRNgylvU736Cn0mUUcb864qVZvJWsgvmQYYsxyjpFBOfO8OejGuXWhWd0C/w17jCFsjuy3
4o3CunQp6nNaclsC9E0rDHDQh2dxSwWnkARo3T6JQqnokEMYhfZrbz1KDnCoDxZrl84Bu1E5Lhr5
6TthMnfdmHAZCbumHv5kqrO+NsXFG0iLdVEqM+9qa5oH7UplqIL8DjVnCG5u9+5z4xvwNA1jGNoO
FKoywP4xYr7HBLQkTcOtAex9vqe5gor+l5pg3c4XF/ByzqMdKH5KrCfSyD0dG8TM8BpCIWLMyPcQ
VVhKBv9c9IIKrf2bP3ENuX85gNeVpTqkuSplYP4SFDN+FdCVZJGuBHBkdKOQSLi1scv/B/gEEDKe
qVkpxzopRaKsRsKO3RObK7zsSxhSc8riZNmkr7wGXI62qVdIlRueH6XvCSE0vp6+aCV7xzDvIzd7
SDu5P9XJaB26j0h0CvWMUoxH/9sLUQysSRcS2Za6CzeqkVY6wJLd/aGi+ON/eI/9BY1i3u00MDxp
5HjZCDNeuBQFmHmpcnPxrJ7HAebk5PV6ZkjPCL/A2+otvP4aX88d7GQIvaks03/MNkYEpSbVUeXz
Ck/AQfdeqUTrRot5X8vpGwFP86a8Q6E3PHFzPAaJPzLR51LyXSYduEJpAAcx00Kkeokr2YxmU8Kl
EWMO3/1UXqxQ2eS2DUgxd00P+miN9vIucK06mXizl8qCGZQ4rbHCBhBx0AGphy9nfX773+gTXZwD
E0gqqhUamFvyY+KR3iUBptBcESCchMJE47/7AWz+SSLtMr4sxi0Z729W8ihNoEwOsGAliT9zzkJ7
ik4V3oOSZhg1ZSTUKn0gDhS5GY+B5uPcWifRWXGv+OG+Qw4MMQ/A7v6Jjspn+a2PSP4F65KxfJrU
ZEpG5fMih/4IWyzdWGgA5erxGRvJlXyXc3N0TLh87pdmd8P6RqFLYBIR48I1sCXDYyUebKiObrJ7
pOeNWZwo9qpMf0/J5/weps+CwYEDxGl0byDl+EmmDJSJ7owkBkX2holC7sIFDlWWvMMysl6cEKnR
LcCiLoc8lhATr3ZTWiZbp89vF1ZiHaEwSd5XQ6z1F59TrL34GrujcdRrGPGeId4rn19NjZkjsKRi
hzKRVOfHO1c40Zu1qd1e7xWzJPabJZAx6D4+DgLaL6pbnKGcRXcsg40de+CzY+4IrWVm3EpNiVVY
RlYnQH08mGbt9Nk3/mNX6CRVzb0s0P8AeL+D+hvZl/jXxE6fOJrHGg/SN4YPNaDzJ11ywKyh/sQc
fVwzSeFTpdQZLnWokvjG9VhAyI9A/PCqhhGYdygqmPANOhjAfvicoepWazRDtU0gFFrGSZprUvZZ
28KeCSBsIpdscsr2aGdq12gaWsjeRUNywCDFjAWMTlq7R5ruiT8rGxvjr43MxcYxqs6NcPcw9OTg
FuViafwnCOwGLIRWMv25jFtiD0gmEBnGnbiW45zTGM8q9GaKjZGSkrBswDC2xv58/YURsZupQSLw
TNK55XGivtiPMQuiQyjcJ/mL1oy3YcKQ0tIGhLJWJcquGI0YZO3HJ7SknUPRd00mg0emJLARJOr5
97R/tli63OK3yj0DDW4Tx4OC6M1nhXbWVRlQMc50Jgvuad6dbJSslUQ29QSoTi/3BwxhGrCfp7xC
mpbB7b80f7FKUZBRgTHU9N0fAvNdcOic6mcYmZuYRXo3zYnSfAdhvn8B795gNmSEm31IuRfoAkka
vFa1WXRuMAR/5zxkakKYhgvcNG8Ga9OJfdcFnJDJvO0TWm0KzRRES8dqthSYpDkhz9Io9t0/NXCz
yM3sh8AaAUElBs2mE2KloUh1rtH4shpmT2JUFOKPeGlI2agzYSzp/0lNpY42+rc6Ptzv+jmHm3s6
sKjHFKBjRv/u/M9mCTQSn6mxTzeV1iyuhIWxAqhCFNeOTFr9nbZuRVoVXem7UsH8HxXdbXNrRL4m
j0bNHUngmYIqilf7QYvPQzySwIzilp/e8s3VpaZQcHibaktz/kYyhmdpH1XMTiYTBT3lfjfhflo4
Q9fRMwvQ1jcIZr0OVLjCKXOjdiTQYvXjELRlhlxcwBemyIgYIncLLFqFinrWP98S3g5a3w3awqlV
RAXgJHvxAAfLMO29aBwmT7p+fPijIA44agayt+UJcXE2DMVp1wvoNlcxQUZ7Ao/R1KHBabGc7omw
uHtzYcwGCdDumqMr6njS88Ts9rMOI3c7wxK6lTplXLfE89afgKDRV2YF+JlstAhZt4PzcS3j0o9o
uSy/1MzS7KxB9N8WzLmQO3oqXdx+Y+5pVuCDUEBZvWKbcTFtwFKQIqG1gFNx4FsCc/tzSElPmGOE
wvKuqrb5D6J+q5EyF/f31NT5HGFqGN9N0zR00TO331itUBpLCOuUAauJoAbf5y0Utc+fzQF3nXzR
+ufKRcTMI8NHeA7fvQLJ3XOYPDwMmG5cFEZ/9r9GpdW2E5qQaREF5l8TchJPJ74MPRyA8/Fq/jsr
UAyVC03SUi62MHtoPacjMknBibLSbI0ozxQ59+y3Inctb3U5yiILt5/s31qy7m/T+X8Psl8Dbfzn
ioGgjj1wyOzLU2L7m6ERtzb+bL7NTGBx9S9wHasoajONaQa32j6veH8XOC87sZCoGYq0YjoYvzes
2XnWaWo2F+TyEGiUfSdAdLe/JEK1Kv5FnLrKSMm+9nMY0qtyYW7A/WpaXy7zI6MFhtrMK5AMp9MF
4k+7aURFPqYYK3CD4L6aCwu75uPw+Io7/5FTFOdL42mtBlURGzRpJGS+PV2L8nKEoqS/ai2XFFRw
e0y/s/oaybjlFFTP2mqtRX8sDYBPI24c8O5TZgy1TBEu4fjhJZwrSNNIAdA8iUUZsRUtD0wL5DMQ
VufFW6fWQo6guo5ue3kXSKQQDrK2/XrkbTI+uzZqcYCjOfjYL1lz8pNZYQxZIieV4MZzFn/kCSkT
3tOosdI0erhRIOY3wxUci3ckmM9Vvu3sPt9ZZMbM63kFhh9LdGofRHi9wj6his6VI7ZtTXojLzJ1
B78y3kVzaz3QUdefb9nI1A2/xXEvWTK7K+Y+TJmRRFmISsRcvsbTD74/t9/6/ATAvU/BYIKYwK1r
7FdzI06Oe1QSh/xYc/ojvLTVs4C+5sHsEeXFL6EF7G7zpB8jnngT7Z4DPC+BVmfmhAylOKqJMd+0
6Wc4tuLHNjA1APT54ahQLD875LkrYGJC/Xsjs8SZfZbAfJg6eUg4AVd5eJsy8XS3AqqZoFdxSB/i
oRwCq7Z3YGVvBy1QOFL3LFVMrob86IaLce7igqNQ3loKKsic6i3muTmd3sub54ayjVq5WKz2UrnU
k36zyHIeZZKnM/P1HXgLNOIlxWThHtZzU+IJRlOKvyPpomu4oIbGua5LlCr6gi+O1/36f9gKelwU
VgTA1Sq9sU5lId+Ab+aKAzzx3htGck4kDiTn69NghoCf7HXLMBIE+/Hf0gjekatUn//stmX5Ogaz
7W5uRtbF6mG11U0iGjvCR8J5f2ivvhQKPo4E+BV9JrWGNMGgRj7gcoLDwZ2mdIY+W8arSnerETeG
M9a7M5rgCyrAd6fpka0KvY5Yxo+khCDv7Jbis2HQHydDVl0G8l/xZjYV+a52k65ikbbxttV0t69T
KCKF4MRmvKfcN24nD2fTez+msjS8uxV6oCuoEltbNFDWfJrHaaduxk0xtQmwEfTVmUvO7SO+0YtF
iAUJTWiX16e8zJfsJVj6L6aQHsm7yvGQ99Kyuc6JmHSCUbuTwgxqidt9DwEEuF3FbEQmVUk0vcUP
RDkONcBJCIH+Ahm9muRkBAOzjP0kXC7SqlFK3Akuzy3DYfA8HAlyeT8x9Tw5ZRxCOnD6Yt7X9fQD
HbIKPa0xTxfLvAaejil1SiSBS1oBkRDFPEBEVD/HLnNd7UU+2HwOQwLpbSOsjO14i6x6BVJZR6PC
rd2WEMsaACBVBExb4w/13O4rNeOpPqBkHdTpsDS35URiJeKtTqsUj7+7rjoPXdAHX5H+2f+bC7b0
bu7p2afoPJH31Ii5nwLTY4dY8XPmD3NQf2bBM3tvJ1mEQAjB4ErqyAtqsraDI037EQyHxc4JQAZ7
M1l2qCwE/t0ybwabvOmnDeodP/nKMETGeYmmwKjJm9sNUz3tYhck6TviVp3fMlJbkRHcGqQ/7/kM
xkrd2XsN/leC88wTCOqMjYOQiEMHPN5g0hBsDINVwKhEDSBUcTYWkm9syv/oJlVnZJA6xFR2hFY9
o6zYPs+HhTb1nY0dJy5Z8YDB4t+KiJsHo+jtmiviZojZj54NUGLvjF6HG68VqPtVX7Y81HmyvaQi
E0vONrGwKEmjh2JwqKKThufGMder5zO6dwcvuGjlWiQ9PfH416p34JHp5XfvKu/odzdLd/1XJ0Xj
BzC0AT3u6NruDkV+o5t7xBGll46DsSXqA/IdQPNAor5KbaBdfeyCNQIINbaUc3PegDZftABffol+
AXP43Bc4rdYdwKMb7u3HxGhVggeVGLDiXxbGxSA43UJgleBnPTFN9dwUeghMBrG8LQO1gta+w/uo
hZWglOcT+sLnEBv2jv6k8oeiCDt00cL8pZdbsEPxoIeFib4YjMHrxGPWKM7OVTxz5rrb6Qt0c+QZ
edua9ArUK9q3uS5RGyWtAkPBo6RxFYc1fiHdAOa3gnE+G0Dnzg3vSpKnmB2YPze83Qy55vLFdQDF
OqLVRqADjYKfBBm+iZXrI1Wel0auHVxDiO7v2q8mm46b4Z8SBGi8sRSJtQGhrEC3XnUQOkgO/diR
WE4tWrJfSgMqmoyKLPITA+pm3QhvQoVHLp+wltbbwsXHAr2x0isdpAmws0EdWa2QuNrO+RHa74Lb
D6tD08vWfDKMr89v91vgLjI9tXn7tcp5+57kTWQPIIfZEj5Y0uOKzvev2Hcp+kPn+7lvHsmGgyyp
F+tlHb5BT/JUtuYhcMkk2ODzR8yowpV1KkRUvNKuK90afKvfuyTh9lD2LL/omxB0BiOzZLVH4wPj
ABIVnMluG+c815b/EaC+PnTOlBSQU30jGSh8XT8sXnR2OxPLkIn/ZWx1OzcmPKi154tAsvPUEi8N
2DiFUaZLT8XF5Kb1ZwIGfRkGw2uD6y6Oj+yRvY5w7QUBLKNl/1j99eC/y8uET8uj7gFKFgCqWYGz
7KbkSV0DW07GHf2Y8Se921S3To6i0NBFhTTC2oa0GfgfGLMMAG6wqrh4DlgHK9MK3/A7tqsdbGhv
V98rUD1unXuE3Y20xNvtrrpCcfksA99vG3/gVi6YbK8kVDSJf93myqjYGwPf1l6U6XB/tYnPq0si
TTTiLnb3Nc0rsdKL9sfg+xKyUb+iRl2tKAYWjSdunf4aakTWt/SJop9pN+1KmRdPnYVfCIXG8RYv
/4hnm8WodMK4O+J/WRTEW4AVPyQdlIbNH8V6QJ4Y3tM6jOzi/px0Vr+n2zWY2sgELHhPY5hDBLAH
zXEJzeE9UkQKh6kKCXiOySvbNY2usEJAc4rdHUYYG8R6HY4UgBSlSLPtwzxI4gO3BHlveVqAeVZh
B6IC4U+NUa2e2bM6keUuzw/H+4BxX5SIoia/MBkYfSjX1UBbwwtzSqq9onNunhZeu7xI0FJymPx6
lvuueGH+2MGi4pPL7/cLG4Rh1lrWDiSGDHdjJe97nIl3nyHQ/8tlm+KlYRf5X/mC4l4Q5ucVN2dW
xLPGSQKCGof/UUoU5+jmdL1vzk49JDpHMVtrzGkUiGi5waIjK+q4U4J0oFUFVJKvxaz7dB6L0P03
g2ipZUnrFxFWlxTC4q2PUKgB59UpE3wBN0ACNpshyCpFwnraoFovFEdyaxIP51P5sPpnfDiv8wD7
5gfVaDEkhrATuIUSGoLQESCI8dzPSkjIPXuFDoqiQbJH7ykrS9CXWYqfgsMzyJ3S4PK2y3ItVJn6
2e4oLXirjwMUDCEUF9amFnNeC0aChgkHUWfiLWMEl6xeNUkgo8doPMAg6g0w/XFpEgSs8xgP2OcD
p3MjBCTp36pprIrQng2KianQFZAj8AIcIe5uXMwRVKP2VxkhFKd133BepXcGDeQGgb3DDJlxU6/d
8f/zN0rS3nXFVc2VRNHAekPp2u8QmP+GEtad87wQR50GB2+MqxlRAo63YvLwQiM370y5Me9YetTA
MNvrL7UuAyfV4z/nPydCp1hdCNujOdytjzVyh5ncKADjC5EtRTbbymk4kZPjessUKMyrH+tCzsAH
LDW2ac0F4GTdaJRNIpfXj2mwpX9mzCKvRxQpJ5VmwajYzSv6aQG7PNvmGiu/4oMNrpjMmi2hFXCL
u18mLMa11aqYnlJ7s/UwK/uiejd/I0hjmNpfspKQagmJvVZxrHN03A6PbY0f1BzjLBcr3B7FFc0k
aqn2SQ+1lKHzB2NSMnOVDP4rQXqw/W6Eh1vj9t/SFmmINw6lLrBcC4CUD6n0k2ztMXpxBy50NpOg
Jg/216fI/z/jt0F+IEiV6ZyFX8A+55VrJy1DtHN7LX0EDsm7i2blyx146XNlqiQkBH4YoprQvhcZ
KEHS/jmthdf0KiZcBrSGp4psjpM0x53yvVLItxbgoqxg2YC8dNcwc5yVEyhkG5K2CRzQz8n2ucNS
VqaU0DfCMuf0lEN3Ol4/WLssP4NREf3YT9/ndhaEL75b+OO0X+sSEljGeoBWEvIDMwPYlKiGNP5o
a5SUvDVX/Bo8TMoQaWpbtL9l+PIBhfD/34rmPNKZMAfKutElOzRRV1n8HR/nrU8p5fmBNghJNcMy
tj3J2TR7rxxCl4dI5s7J06TH+VtoiVfjfx5MYXx/spRD2IdW/fe1BcFzXUheF84SkdHAwCV8PrWt
BRcNZtcAns5GRJjoUfWl2dtLFzqZ+C+Hl+FQafA8+vgrPrW9MujhnQQOwqjenJ71jIbbZ1VGgwkI
OJP4zgXOINY/l2xTlzPNHUqxBnHMollx7OE7GQ8CjG7IJjxcJeCLgeoufpSCa67WA5TPlEHw7OzY
YRSiHMG2duoan/EGC3qqgUYlquDiT9dg0JNCEWxtHrc7FTuPxe3D8SQIchWbgBKoAqAG8QC/cxoG
aXruXYel4eBATfG722QCqf/Dw2IMKUkrDIun7Bi/SiD7XM/i6OIJmny87ZF/CeTeFY/uM/zl9KBP
Fk3aRKiwOwRlCPy+WCBClsQoXaoxHb9BJOY3sEitHUH10KzfziWwh7jWN3QwMg5Ae2+NyhCKyOhP
PAVt8dxHidiyv8YCEHapG1OpDvY+m85qBbpKx/h30u5TuT+NcnhDcF3T5X1IlfOpmPgKHOHASpX+
+axBiA9teDyaNrVLdwsJYcUFBRw6cMfJICjOQGpU3WaCCoYFI8c9tyQgtp4GMLy0X6MxLXr8+/R4
Uq/RAG7KmGVFga/xwRawtFJvOQQIP+3Z+NzaaUGg84ZF6xofEFIuJy2Aq2fgOMmnx1FNUz3989hQ
dETRnfcHT8tYqIDwGv/VNmh5XlexIFfw5vT7ZJC7xbxwsu1/JDekkdzOHLECcAPqRgXB3GJVoO0+
DmEiPBejYDGBTBYPxqBV7WoP5RZIvhRW5e8isnyXEvwvcz44zun7t7G4RvlCglQotib0Tkzl6x2m
KGmAM2A6kpRZHks1H+AouxxKM+ffOEF6ml/Odfm+lDP7jhxebe4xBpvNa7nyX3ac9iWDuDJ9oTUU
G2HunY0dRamz+910T+DIdQnRU0a33fo6QPTGb0K83iVqIPyxHeg6qTFfo6D3+4f/tiWoj9gO189Y
sJkDZ83ROL+m/qHV5wpeXvlv7zr/Or+dwpyfeMnBLX+k0UqBr4CZ+2JhLzVpCM4CoqhmWfDNBIDc
foTejIAGLEV+dhw34u90f8KmXxfvz1xfBAWlcm7KFD44PLTscqM/TnerbcCMD2Q7oaOuLXGKq//W
rlXxtj1wFehMxl269f1NKEzTuVbT5p/9kKWVlTUiARiho8lFI5hcGqhYWP9kGhYduqO03gv3PCOW
EKR+DGxqNq9N4Q0s+5FFgGg604trrap3SLZr7DIJ3YHz0eLqE4pSskvYP+vt+xQ6B21RerFBhxeW
Ar/DjSCST2AQSVpQidiIS+4UJDGBuQNwwpnjOlfEcazTl295EhZNXvB4r7SOlrQZOxiJvN06cf3h
4NjdDFjViV/elo4+2+xey5VGBOaNS5324bW1ebzEyETdfFIoPQd7nyPc8GLAE+e5IJnb6SNGwlJC
QWG1kPdqNmyc9lRkXW3udAMIj2sMdfz/p3XfCFnhagklwsQRKXXH3v1Hp5dkK/ummY79tx4CzkmP
HeH9UtkJ9+UYKspEiCAVNrd+A/0PuuAudhR82/9JI96kCpGfWAxEbeUzApQYcB5JdlErtPaD2CCn
izsM34Q06Jfopnu8f6Rf/WtiLrEqxKHiqg/juivn/FFdxQvjmejUCJiTm/jw1SkgF65jA2pERc4S
VZB6zAc+U55XxqePUS8B25TQwbXHwRCeadQE9K2UpY9REW4EXQxv8ocoqObPrJwahkpi/UyYJsJ0
5m3BO1E69AufLbnwNNm0nKr/pQN4abAKfPjJ1Q5YAgbDbhfz7WW7LzkIx3OjATKdMjYYRIQ6TD3P
hNv7v0b/6Bdm75GLyX9vMxu7G8xaRlB/RgxdJejvn3TkE6htx5wVlbnXn1f8hKOyu9lVViQflOc9
mPzmOUMYq+RYOB/VKNGtQjZLFZXzmqra2ddAgB/sMbCg3xEKUV0dvAMPqMMhjdYZ/xXK+FAfBRu/
3GmMSX5cnf8/XJOi6kAs0ty6/vlvgYfmqiiLZqVtFDJpaWMK2DIXf5TeVeL6FadCB6+AkUw0syic
svsf97oZ4lc+Pl2pJKB83TSmas20F/zLMMhaKsiq/Z1HIQujE6rbeco5dRe2DvqOVy7jaVgZiGcb
KgjS03NqouuDGbr/Xfim1uWAu02kPUQM8EZQu63g9Eo7SoX4aCLEMVb3QVeLXL8u+vuKtrHz2ain
q0vtIf6q1pDUF6m+nDk9DSJPlegdbsDMEUT7gQaXC8nurMXyIzH5btvUgHHreQA9r2/jUnQ+GndG
hOeg53EoqpC0H+SaapH0AAlZaq4A4bgN3AoMr3nhZHWyf6UvrJU191ZM13VbILs6G6Tv4Hd474Ll
XAPHI/09U3e7R2UAezKBCWuDACt+njZ15ntjuIMfFzJ6zUH0EuH1+BWMmRElVdHtnAv/ysWZjzQA
wYjfPkShGpEVgzPpG4jN81ankIn3tuaVuz9h5veuWqniNQjedjb7xg/l8xaCRBF5IZHRg446lJao
8VzJYgqwClOpiO+S9crIwbsVyIP7X2T/ANrMUAbJTEamLX+dXuRtPOPKmbge7uaVP8X6nozkenbf
gmHc54TzWbeMrNrG5MQPW04FhLloM0V7mRIRva1EVjapdhkuyolBdjcamdt5PiU//GdByUH5ZWkV
25IHHF2G+uyHqKTlOtEdPcnzP3G+Vf2FORgP699R5In8K078JMcNXdstnI+M+nM4oQUiezZYlBm+
/lqRdsBgnlaZW8C6DdhsjaEhW8VqJLulHIwaOySUFNI+e8Z2eNj+RPHZIimHdL6OVvFSUf/TVVnK
F8Kt5C9f7BVBju8Cs5h9Un76wOrRpSXPmO/uVkZJPBpmcksMPFVE6YANlZZm09ygfSZYb4JRo4DS
DFBG0tgrYurjdFSulyKEFWuQrpB1O+nz6ySIffkQkG7YcElYv9ful7V+LVYOmBEXTYEei0djxNzP
QZDGKGZZ/Og1dq/5kvclFPlDkY6A1bFOsDplhbV8lwCgYZ7WVYGQY3k8F4rNf1doKutM8iR4U2JE
okTUciV/CwUuuTe5D8aQXoevQ5AtSlztpdSG87QurVrg7c5b3x7VyGXqsI3mNBvwASZt43o3Ra6M
EMCm/3bdogsfc8Qu0udMWpg8a1AS/NK1Sk53FKWlD4EMl1l22ChpOQ8jxbyJ3a1nD7LBHZPQw/MS
YXgShBGZWaAWwDPrmlkcLteSN3C9Ybs9gMAsbceij6JPUmWxovqOSXvmILxl/TMUhohfuu6jaaVr
J/SXEs2y+0PlY9364bnnRb+nzkMhOS47mjFgM+dHdVVtaiuK+YDE5929jVJOcfuAE0Mhf5sg6mGm
1ANr1MaAvqqVwQUSyUApDlbAJ40wojFVxF2X53pYMuCu8Ceu3K4eE3vZm0QuDDFQpzGyqLewUd1E
o76l6vbRGDP7U470N+nbbvjFtPqJDroOnWbyXmhwnk8HRXqRruuBjZahSh+62u4JdgYdVfcTTCM8
FLbHjFyoyUscR4ucJgQNqKQvNUasogGAHDpqyx5PmC25LP1hBWZnjbWsuqTOZEfcOEvY2tZdgF9z
EtVisBlVGW2qwykFzEqLSUYFlhmgNwfK4gd6jDmf4QJOfYsd4W+EWIXw8lbsCwBWFKevfGLFcQ2K
LhH7M/bxiKTQhnntJB/nHaIXMyHRlz1mhvapJZBBNmhUjkPbz87oCuowwPkQHilOvgmBliTnQ5aY
B4ap6EtECjCtxvyKxe7CFo2FYTzKhkeoEeklxnMqggRV0Q+G2c7ZPQULAJGDq58P9ooF1dC9qqJp
u5ZglnVGhgoqn9j6dyJ1e5X6sGX8AHsKn/ROV6Eyyla3/+r7mvkI7LO+y27g8gPobQNnCQ7q3pev
e5BkaM0f1qamiaM7YxmE46p24qGSu/fA4hRaBSBHjLyfiuCcQt6bsBX9vIAp1qHZAvVMBcGEphPS
+oYGUUkrIRoAc/BD3YfQqkvgv0YoBd31h0Unp6B1PH9KO8XP0kK8rggnQ8vXErJ7xfE1HM5x2y5f
MGvKX22x/0d72V+UKx3yQT7+LZpG9IChRweAH9pJmG5C2/r82zcgprh8rS35/+4ZYJPdKq13zA1y
sUYq5jzlJh53iHEwz9sXTnobhjZWfp3ZNvmpRVQLuXIH3zmvZPuEO7ljcAwrP7jd8ROfrW+YfsvL
dW6qwVjqfvrHNzwN+5cpRnUN1NA2kBTvzPPE5fQoTmnmgD2w+zIthgwb1fZ7fJdubV/QzDZZfqF5
ciiHiHkUyf9PoC9hQzHpMJ3WpnwTtLxBOCIL9taj32Jh4l0q5Lb+IAW+DaWPGy/I8yqgreUB4BxI
AfPCkUI2KYlH67KJ0b0i5sszQMSI4necTSmx2R+gCMGoJih/sHqZd0BC8FbJ/jIKMGneYDdOejST
hsLvAF8uBpwht/6qce1e47WIs/J6Xquk9/bFDasimYPT/chwZSjyKw2whQ4GySSOZ+nJ3Xlp+c2o
6plHerXdde6vdUL6rzNRf879wS7lzN2vVfTlZypoklhrqQo++3sdTyv99E3BBtrwU8C1ls5Khd8h
JtJsyw9mFiup+svP7T371x8LiKQVIQUEs2wcQSl6PyK8wekjsr8Q4Hj6pWqsInnPech9IzPxn214
iU6YY0XwNCVCAt1e5UWXkmxQ8ubtKr1q3E38UjNmS/gzHu/zu8RsSH/4Nm12VSTypaoLamVbVBih
KNSu/mJeG4SR5Y8mWXW1f6Q307KziHTAqAvqEBRhFgwg8CUcfdXz0bHO8SVnCAUaWZN8CItree16
SaWvb0oNMlHcVLu2CgViDBXPcwykeJ8v33Tv41fgn7IdQ+lst+b6Gc0SipztyXxDzEoi5Q/Nbl/E
PPfSj0+pRjmA7yWSIhKaScxRFTXALr4xrqtSfBNqjbxDq5fuQYVLySePsOfL2m5TPoMGlSQhQ6RN
cFAp+fqo/HOyBOy31Tn6fabt3dexTHrgy2ZHYwFUY3c3TLJXPr1kCJuucgq1MJ6OGICto8HMycG+
VDVCPSLQucVU3xpvzYWxAN3r+UtYL/VoAwe3iQfw0heg3/XM3YGmefuY2nqdUn385ExMc5GmoY7R
2yxPjGX3KKpivUVdwhKG3Aot3xIgz9FKVPSY6C85Io1yDwelDcfTIg6gm5R2M/IA+0j2AYpXjVR0
DUamyjnrm8JjAwSepQnkSYkxOKMAO87BdLPmSXQiF/3xWy+kCWKkvSCA55rhFehVOalnAlMh/uFs
qmnHeNn0lr12cpKbiVdDgsmtoobYfCd9/869zl/mwR5PuAylvHSY4IbLntjiib7U+HdgWDqY6cOf
pxHTr+pmIOEEH3r2antKTXDL7hshQZh1M1GDamTO4t5k4bvX+2tEDbWmqfnUspaZGqN1a5WCQ/eX
kTwEqz9pnxdqNTdLopZwxE0lma2JfYpYggnNDUOj1s3VvxoM182vBPteDadj7YNsU5s3gYF1sYGh
6MccX6IqOWq9edA82fCjeQi3Bmkha9ZHvwGeSOsODdT8h0fv39EDJiFOI3IAUz58WSH1agxnvP9Z
XVrOcIaD5e7pOnUILiR5NkSbt8QUA02lRgaM6XF4csoY7jrC2QURvuTnF/+klKRe0yHkj73WqKsw
esooiNw3BB0MGrM21RqqH4Rz92x7c7fHQGNYWhm3aQF8tnHKjnN1ugTZLm+8ap+u4e91mRVV8m5U
zxX4N1gidJMnPi1bUQDbi4HrcP1G/ZdSIzLRI6fcz5FqRi+dEoswBMoI+nMruBnXnoLgtSoknuer
czS7W1bIEtTv0sNcY0YafIbUIEhvPoWJ4D+UKgG1zvMC0al+ToBECOP+UzWIVeyK3J4ckCK5LNWz
WbOzn90wvV9vptsho5B7odQ/Ud1Ba2fbwTKrXVz9U1+8Tr6jb/DY6mKVnhAfnpnO9icbG6SiRsJv
lOckRHXFrKLCI2F2cQwhRInMIHoJRVdZbxmtn83zfISQVeU7GiZH5E+lOTkzqo1vYyfVUCm9I4Y2
9ZpOQFVyQcYxVbILY6Dzs5TqYlcQMyCpU3jLmjhGxlq7jMgI2wbbvaiyoVPdC2btCtFJjGy+Kxqy
gA+835hE6lMzNgIM3TxRjIPFrG7TPN1K/T0+5PNKKYI6vOKsgyTpygKehsONbuHH1nJ8sgS0UiqW
vtuAxDwJjjGWZ02RA1tNA0y2RFQWyJZAkNzi4vf9d5B+3653ZlaGbhRgVDTD2v6J7XscpbGocN+0
Dh7Rbv3UbJh+4C4h2Vs0D69jYIowLWZYfCzUewNjrAwF6aenNZbKXR2Yv2/srsrmhGnftBoc64wH
yJcRv42+6XY35IURb3XvaL5YOcVB8gpk0rMBWV8WB6j5zWm7zBRqaIEEhdYf4WTQ9iZyOJ59Z6by
heO/5z+rdCu4VxAqMlbbKnvBRaoSB7/FfXHE137fVt76AuHU9sTz4/okII1PVnZ1RtOMiUoZWsGk
dP+bZlvApkFi2tkyAZRWGydcJmTQ2qAqWszqEtctv7EexQkofguu6vh6CDlmR9FfROHMCo3917wT
EFlRwOckEkjmaJu4IID4Xju78eq2EKp0q0NbvjvEfiLisFnbYxAMV554xVzDQ++dVrhs0uCl8Mle
FffDZoq+rhw+7liaruB6S70+XUzWb+hd8jxEJPddwxuKWffEX1pVLeD9tzPxJfKzxLgIkf2bkeWq
xnWyF39p0NMcvjnJ2xeU3xs61PMX4+tN2VTjXXO1ubCjruE9YMJY8AOD7cil17I1E+j1nvDa/Jg6
7nWjuyjIPwR2ghMqwtyAvdsgYy1WHI078DDyrlCrN2FLWLMnr9xkHBuXi8XdPU8aiRKWAFXCD0fa
+ixR5qYM00g11yctViB7m5klwQ3KVWyAe+lkgtFtgMHmx7mv6qlNJVlzXUtJstuNdSbi6r6yY3bl
Hj8EeT71jJUjLJHPqoWXTnGXWkuXb7xXXTpdvgjf0hB48Ni8JwKuxvEB53g2lecQ87LauTvbWcwl
NDC09xZ5jzjofbS/s4ggX0CxpHsnDXYT35o28wfEP5MiS3XpZr/vmqM4yPXr/+K345zU5sp4EWPm
qSe9kNyzAZ8qzfPuUisgtNyVgRBarBR/en+l/KokTxzzop/PpC/NweLcR0j3WW611bzY/INqPsl4
TwjSwyh4q+zvekHJv+EczT9iqM3zKnJw5RO6QJMMiS3FZqU2qYoYTMfPfnZbvW3EmsoRO1TmxB2v
YkOYoSWklFGBPz8WfSxprddkgsxloHVTuvKaqinuNtDrbDq+bYjSZvfxyCTOmGNWCz5TVmBSMwY4
fcpITly6MM81+BET98p2VT6gtI/I38EPa/StO61f2Rzs4NhiIhkZLwNHFL9i16xYH0nWMxr4T0Yv
M0qhHZTbRe0xzPRz3ZV321IS9i+aIEpm6ofQtA0po40hJKwBg17BlRFfVcipNdYvEBJz3EIO4tP+
tSQqXCBhhTubpnG44WENFTOoJB+ojaJAKYLnn5yO57Gyilyva4+gsJW57PzfBO9s386Un37Shsct
S/SVA7KIHMBagXX0k3GpBs8vz3dtfTtlY3fhfYbD803QweirROCzQ8czXvtudbdXnwqD2aVLfeWe
mReVbYhToeoLQ99EpC1BrGKS3JcuNygmacCX6jycmgL68dd1G8KURRu5MWhGdZi5fmTS4cHLHx94
qbk5s3r1PCgaOgTkCKAGRJgg2nh7QIRFOPk+y9a48meu/fKWWhfMD6cS1kY5+7+7fyCgAnKKC2Ec
l6A2AMIqTgNcGzXeB4Fhyall05nvL06S8tIjALJAlKn8kY5M4ufY1TJAzMM7VkXqXmwUsQaasQtd
vVYqOX4Xy8Xj5e70C8lMMqhp2EDKBYSlQKjXzylHYfxgArDjY7MaNOpI4xZ33ywdye0l+Xkk9vI9
jiTfI6U02RJd6TwHnrqYxoKkNTk4Y0zG6fLyPMJma1fAY8IpvAQYf0oWGbMaxyhjJNpHXLFa6sXH
MOhu5eegwDtSBWFSXO9x+YjxB7JAsppVgcXKu9GT+Yr8Y48LnjUkS17zt/LOOZtC3e4LPe4oC5aV
aKuytY3Bb1FBd3gE//M+j67qzj8t6bhTGHFRRG1iTBhUOKBPVRy2EsgSN9/uKBTapWhV+/A2pCee
rw2ez/h7egUOb6OA5CqDf8z0V9Hi+R7h66JrnLIg/e6EUHLqsKoh49YrQ8zX7tSVQ5H0WW2YAcuZ
1PM5cyEPJ1SOWGbNB1G1rCtRDIhIpuX+U5n/LSZF09IFJOoDG/QulpxlFj3ll3Gzc84Yovlc4+FH
w5i5O1CtxI0BQN1Kn0AIaN9wXemY4Obx5udHotVimj+NqsIrX2LEkYq79wSp5v14GuFnFvvC+LUb
WeNmPZHtHICnYeiBnNEEohabCoaSmMonpSd4kWyLtvhd5DKQB4rv6iOiYrztsbDKYZkvKE0gaiJX
1oKiEYRGG7AAA/JdWY/gxiW9Wd0uV4Fn5MPxc0T8ltNUYEU5lf4FlPQgq9Hho7H8ze+l7xizzFSW
vAmcDLCPJ/ZNEZpcT6MMsb4R5gIWLvkGaGfMWJbON6xRFr3HXBsNgzkSHcX11oczRlbJndMKQGYc
hVPY4S3MiWZttysBv3SrAfIU0OTnzUqtsW9svgEBuhixjQHFrhW2V5Sela5O7RU/Uz2By8oy2B4H
ZqBZjiGNld3VVr2ocwgmpujZohXZV7sjzetBbAJSO2YCnVnbrvkzU2zRp/iO7W21/nLlxiZXCI2a
839+GM2fJjXMsxkfPFl/JNeWUcxhCQ5vD+JlJWf+PGmKucaLyR1T4WRmYsK45xiFt81lg5ofl6ur
W2VLi+1Cfdbahq1O+FlMARRZE9PxEZ6MvLZ/qkRp5Ee8Vfrr9CxRQbVFutAdgPIB1n0a5zmVJqTm
9XQf8G/QyWcHhm5joU8Er8RkYW/9NiInm8dwE7jffuWffgQFgchsoZFL0pG/JlMJ/Zl0GSdrel0j
V3jFptLs7I2deXH9GQOH09S+BYE8bv01RB2Ki+HndiGi2fCJJUchP7pskWgjTzFuOkCnKdBzVrTc
EduYqplY9ZH5udCuNjR9Uvs9o0ccEazjs4d/kAUZiCqJwHMCp6QgIM/BPHg5N+7k9kYpaWjdSmY6
VWLLyiqNIs1LKxG+v0ju3+uok9kyZAxkEbOlx/pBCgC+u3nvthqkkUj0vjx7wgnPANDH8OoC6hAX
1eU+7lYjhHOBYX82fjT6+b6NO49ACAzzIZVr0gtoXbg+WaEM9U/NhA1HiVtzW1ud0+PC7/n+7gjo
XHuvZAuxWrmCW5yTy4cHTV8xhp1EXvnpdAWkvPf+VE4GkUitUmJXsVE1Q2wqt4fMPlJO1eBNXi/6
aEsTMLk2bDfbdqEfg37zmUSEA9kqV5UapN+b9J89xQpcS4Gi7TDklzE1R38gBvboRHo+g+G4AvcG
/ZqllMbO2Jpkb4jN4IHKDXx1ifrS+cDyG7Y2qu96BnpeyxbrE+WEN+RQEpp7KKEHkLdzPjnXyoaE
PAiKexiJAbKp8slZMDm8MyT78x15XuA1emikACb4+wLOzl90eQuCkKLxmnKCG9Rg58iQHENsJZ+F
lkrJO5LthSDSYnAQx52aCtNOw153OGTphWWDNChy+BmzCpO5sHAFY3hEr6B7I/i+gjB/jbJZSJR3
mxF9EhSiSHUEsdcV1BP2/O9vGozAlA+hi67n7yqxSPIvPymmEOtqxocvpqw1W+sKvmCXMCHLZVPc
cKxcdj2hXuyskcitnztT35CCvIoxzrsIzBXm6jhwD/TNjiYnZpd+Vflwk05JjTdSn6dOvS6KUOUs
DTwXKeYVobd4xR+H6iKFUYLUlr/QkBVbzLi+wBoQrbY0EPhuwx0xCyXlZ/SvpklOR9cV/8iBm9H7
A5yZEluUKrpP8UI/KJ9CIIYlc0s1dm7oq6X5Si2g5tF3WLF/y5BsB0hBqAtP+MHWPz1z6iCTB3Mm
3VIAzoaEp9nn+FAXyaflxljDDpotB/TihI+Jk+GDFo2diBpFTGhJwk2s8CULPf0/yQuZpNF/+twD
n/dYRqBpte3v8wkU3WRSK2hXSS9KPo+OHV/apaXUEeZLZ83ba0h6ZawPBtuxItiyZGyqdtDNlI9A
GJr0R4NW4lzFqJZbYoEkblpr8JpfW9Y8tKkNuAt5biOiBRidlFhHy/qN8JtttYcOvAQugtnXofdb
XpkOSqEZnGXqtLFUFNtL2iG7m9rLVX2jq52yEKURRGU2C8eRpUhF4rXAA5sxgyVXHGnnXpq18uEj
e2ee0IgyYFxZzYwlTTMD2Pj2gl7cu0k7kBaaYxebAnxByguCFUClwjGE0eZ+ESK1lGQP1bbz14tI
ku2AaKGXNq5p0zr46LmQxLwhQkt6BVfjp2zk0vVe1wYaHNc08KXUSv9bv7xAvqmj5sBXAC24xG+y
L8CX2qtpD8In15BLbW4scxZKsGKNtWCjsgmCvPz8poXUz5rzKVe3HEFt4sZncZ4PmNwoGdpoCErw
YDz0+YjwGmiqcipRBx7ZheFVsjyQxg2Jc5IDZbLVCx0RteYKHXXMPYaJNMwJKljACEZkV75CzpKn
Zd13WBcNeVtoGoLnDZPBwnNLAzs5x4HIMPorqCNg2zz869XPTLq5gUuCUIl9q1eoDP9n1hngNU+z
3anHYOuwqWQzoHJY1N5Y6sDMDBXqCcE72YYqrjAau4BkzFHX6WrNix6hv9nQaPZdbG8zihXkW0+Q
GiyLqwAaIVhBQ9kAge3ftMwL88oR6cq3knp3pZ91d14l5fZ2f5Q2fLpuWijBU/p6v9OYA39d/6Wi
ZlB36i3O2/90Z/lCQ6zsbu1RtX5B1hbxyji+aju6LZFgIk8WEH3Qpc1kX9pVEX7JzhKEYiNSZ9Zm
XJndq8+WNgN51R7QnBVoWSWNiZ7eYvrz5srUuZr1uyNw5SMWVfJxxjq4SBrLrshge/BaUVxx5QEf
122h43HtWWte5+fVflgWynkipqhwvvYKu0FWBLzUKbZDdwniHMCEebxP9qauVxLDng+7TOgAE+9W
WxL2t0x9I9ssPDV4KlbUemGd5LG7CvgorynvRT74Li7tHVxjZOt+0+0ErJDzaC3xqX9EbJpNP6YM
UJVMoCYjFab6c7iNspY0sHOdcgQbBoZ3s0YZ3/64JRGJdzlqT8WUq304F+Gf1pFDcYIUljdiLp2d
xUEtG67aeIHGnVm5AzYGyWWC3CkTmXQzqvNmq/bdtnvb/Bjuum4s9EeMQPNTPjL/j2ZKYOFleT6k
yoOzwlq5vlRQ34aB9pKwkUbpz0dA2MrXDZzQ3SgzujNTdbnlHTIRHmaGIs58NXYTdl3OGh08t3xe
TIMbjbPTDCLpMrVIaX3rj7knU+R738Ow1gG8LAfS7I3LYWRuVDLaqd70JdEpSkz2KqXxVhav0Mka
a1aqTzCFev9e27ci8kq2huyHnABlv1gV7ZqwMwORvsElXDu1TzYI1JcSCjs17kUjyfmVjlYnj34N
myB2clWTtBg6xjVggWHNl7BF5Fa8IGbreQvrnBSC1gDDW6XxOH5fIwPl9f6KfYnqBgFzd3G2ys41
2gfi89MHEcCZfMW4G1M4ZTBnV9Laojhv5y1BY1vniA9zrUMLq+Ml31aJbwYxYMD9bshVOjMK7uqw
EbAhu+Oey8JU7Jj8vatrFQKcOTBFcRrNwn12FSYWDCHnemt66ceq9m5+XunSQ4vSWAJzYVaqyQ/X
1QajBt+krSkKbKnymsz2d5zkLfo1i5soJGdCYSLVgr/NWzbUxcmSOaHl4Iz8ZmSPnLeIfneiGuty
7fdyo0jp1ZioUlQ+e9LVEI2EQOfH6+jRTaz0xS1XxhhHD1gHkEPaaKZdrvGIDNyqYA6J18gHnHo/
kIPhSHmpecSLcfTKtrMBu1Bd5Suvmgp7M7qTwaRPxHOp2RoqZiwqxWjU9BfWaBheMlINMQKaQNz+
IrB3MzsPXaSp2QumV3ZFL1P0LzaoM8FWg3lJqPdEjovxJ+gpiwnF0zUSjtlRq5cKusIEUyBqe1r4
qaIeMETBDLZ5vby7G1aU2+2iZGNgWIV0jeTAsWJe0Gct0aMz4XX8eSC7w+jNTtqkePpzk4eAiESC
vaw5nP5wTbyTOZ0rsgMLi2ApP/M/AA+jYnGvb/TJCfQb4ge37fXFBxv3aTbDdnDt+mQIc8DDg3P1
LMRR4Yu6fJeJ05mRI8C5fVnDSk7m/RFQ53LqfrxGwuArauuLGoxbAsPr+RN14iC8dLzDxm9UuHZA
wCQ+cFROCm3EgzpwzFAXxAVNJx1AC2jGoOMSPXc2iRt0P/zkSfKw6cCA9YBCEAj0powZI0/Fy5Cu
pm6WM7bbqqlu1XD1N0MaufTbDgvKrh/ORwOylYNABCNRqOGtK93F/UhlxbFExdvDKEaEssQAz+Xr
l+KGCLRiiMzHMLqH/ttkRm2nyGvBXXmR8uWVJ2gCWcGYvoRTooDAn9dycCR1nr6H7Hm2M6cA7dn6
90FDg6ysChnR5GvErVgh0xP1M8R7h8VJfRicq81gYrYdOUF5Acx00Hro9KyUoQy4wAvaKLgIionu
qestKEqo28c5aijRckCL7QPUHZR7sct97EBUNKOAKqmny68whPVLoiMURpMVpjWy0Kh0OgQpmqGz
gdKFyo+CAFtzbPmm2j2bf0ja0BN/BPNqiscjk5sg/FYJGJGZjdHT39p/Cf1w2RV9yrqH/QESgXF7
wCszjv447plLc+TsrdQ6kdABBYpH7QMOhUm7sFW7WzaUhNqZUnhDEn+McYfcK4HZKvSTI2+S4aPw
ZThjbRGVHGL6VCSPKCgtYJDcfjnhzj+3v+B87TYZsyfkMesjfckA+pWu3iJPMilWVmAqKGopYK7d
XaoVmuuxMg3oa3NJpxAhPE/kI/b/Y6/baMQtyLPSy067q+2HZoTcstT2RntWJQpbxFmfEd322kg4
1bR3F6Br6PKSihOyP+Icl8WS2aoyXHpfaKVP9DflUMsNqRr7uuBVYv966j1APhfuxbg6IEBvpFsD
loL46AcN9LF79fhbSMEGXD+XJp8GMNllFqzgaK7sWYMoUGkNriU5ieISxIkkb4pKugh7rsmHMahw
wknpgCQwvsvNc3r8+KNu7QKTlTCMvNWy+eUCTHdBR3qbR6ANvuhfNGrTTjs93h8t6Z6eKbMsZmsu
qnZXDtqFEFOIKXp7VOmvSA/2EFJP4Pc8us27fAc2gDt3zHrZc77lT2spl64ar8+yX5s5umzG27Bq
6+Y6GA6cxPcYy3uW+YEaWH05m5QdvDg/0Imre6JZKKFQwDjZe55w0LFY0V+Rvq2X6gNl+PExmnnR
+gDeyhvx/M8lTMnnt9aA41tJMS0H7NDlMuoFc4aTHOLiuYX/Y8a9Q3/I/7Bu5dTAn41MDlemWMVs
J48TXzQRWunqC+X1/KCIGoQprQFemDARh2m0vhoJAq/tCTk+LY9D2z965w4siIB14f8BOjDDYR3Q
0Yq4DGC3sjLUYDabgY+1wau8TnDoThB9rH9P6rn7z6GxuvKLNRStCCczLI6e5R8EUmH5WXKCvyXV
bi2dPW0EaoRlp897ExcxnWf11TX1JMGw4Ec83TpJczWMW2ojr3DxnXRyvN1m7/Z+71X1HzWAwzhR
TE7tb7xtjPcHqFVqJWXBPYlY/BotBoMzajTuo7u15UCrnCnLwLP0QYrIQCJphQgoBv+gsy9H6gD3
5InZGpIrYelcEw/LMZlBCtl9+qb7me9pAC09Gm675BiwfGtpNy4d5oy/kKRV8IM44sJgmzRsHPs1
UUAsdKzLMrHM+LB+EGaIsOr0E0dDPymp84wX6ww05QOfxaXjjtCZAljYcAxeVSYHQ/C3y1GeFhvU
3gzBiGNCoHToLbX0N4EkRSoUGRtUOSbS2Lcw462WZUimu1FS5XXLQWPvhETI9WZ9juZyP2YfGW3Y
+JBiFCfmNF86NVhahNm+rJ3edLTLFtY7J7eTGs2vhpqcJf7RGzc879TuKHcPBquNGjDQspg6UwnY
TE945eMO9RQ5j4mqLKrqWn1q6hUhkE9enHENdez4mGOLp0EYZcZQckYvUHhaPfOq0QPaLmjcDaLi
rCqjlkmmQDNgG6xhOV5toIBuWMT/6pUKNpqCrdneUW+kGrp6Hv4gQR8mi5+Y+kAa4iCXX0sQ3qEm
DoqP9/tLKJfv8EAwRooTnW6kuLkWsyv0xUDJTLe5Q9WChP4iMksiOacfK1xbB4JCZxlmuNFagr/g
KI0QJJkuP3GGKWHpIW/MJNohb/zFA2KwSqLqZGDpH1m0OuhQWsu2r9rF7F5LNfx7lUTna1VfzDjY
gmvSltrXazWRoEPsqVnf7rvx/Xm6EYOFCRVKfZcNwrSeyY34hX7Y6A3PuYFhBtdvH0mY6gbzypZh
0OaRmJg7wEPtWwjhbiLHFh+4+lbQj8537MSM4WIEfBFBhuq4APqdLYv+G24IOUcghFwPR5+oSegA
iQWt3d1EFuX939EmO8l2jS+tMWE+DO3IkWPzsDwudIBAsNKuNdjfkFzF1A+MiE2luOc8euEOpp+L
JEf0H1u1FV4kZOXViMvf6J7AW5kB0AEERTS3RV1I4VS+bdKvFK6bIgVtQshE4bfkdvn7DHoKvQC6
D4lnYIm3mpfihRIQRhKboum22HAhN/MIMyHnaUMN3Uo6Rwfb07gDr9QjLRyzQEwGx/Vi3jfkstXr
1qTOz9txJQFNoP/YpeAqPl1qZYeIje/ZcMWGUwTD0+XuQuX816rU48U9P0Jg8rdt5StVq2cDYpyh
+/6XGt0USEsDcTZj4u5xNgoF0E28EIqWfxeT9lDPUE45Nej2UKBL9eSo9MB1t+p6DG1gRPuj3m0J
emCXDmmnGSEMy5MX1Mcp0oVVtSQaTKcqiTq7KN19AjD3ajWRXOzVb++8S94tYDWzHdtszpZ9uvNS
TJ3ZGrcypie5+86aJlbfM92zTcs3s1kSfyaNIHrciTJDDXEtZC0GoGS7cqvbj1KPfTBJWNnj4ryC
6WFcPktCMpXYMqSONqaMWCQbCU1xqSFHoByGQXkORntJgKL0OJXtM7yorXnPQ8n9YNWZBBTXHLCe
avBNyinccTtmQbVnTTVEUscsTKrHzXoTSamuxYD71UyQXdCee52nMt9Njix4K2CGNRqbMqKNTMzA
6/2RPZmK9m1meLKla/A+Cd66LY7Qt6I6Dd16amh7yfEGcJ8zbdi07WIPtaDsbO3VbwrAvEJIkf2j
SoooDi82RDCYB1pruS+JM5C/XJb2ZyJ3IE9dxUfBJTVWq/zmAaruT9JqSIMfyfaxXFO3ONiMq3jL
lLdjhWXbQEVTMLaDpfQgyjYgcmV9GUoD+9QDSGF9nvcMZlmWvpT624hCh5OSiEnoBPCKnv38HIWo
oSbS7hqxyA1A9g06GQTTObD7whSE2e3zVi1jUuoX+O+07G6wg5ViKOX2gEnbbblXVbJWZ/MmLrHE
Fb8rLKPuEN9/P/ZKtRiD30AGLxkO3uA5m5nI1LyGkD2iHdoTlJuoVDZoBwk2Y5/h7BZWuGLdpAl5
VJZ7OYUCxk/z9zWn7uLnkFkAzzKSNCk0u6Xpw/ThJDmPhInymIgnbeORNkIsALNfBZbVoHDMpqA6
NoYKGS/VCxqQVGSxp8ZbLAaHDyUpB5ONdV1wQ90qEWDnfbIQy01zA8nLGwG3o7UedFj2kSfzsqKI
GWW4YPKaiLWtEZjInIpGUwzyprJY3f201DBY3RSV1hbT/8mg3lJn0odB0sdLP8StjzrjCpTk84gb
eAJQwoCnvRzButM15a8o/OlucMHJtjn75DguRm/UV4ALSYYZ8Eg+NCy/bFffTK1KkucywkMWmZ/n
f1MeNx+MVX/SgdDFY0DtXYIK8+07cpTYYQDl7dTXA8kcwdr52N/Vt7zpkpqUwUOCAYFIQ5XxMXVr
2yKC3yp9L0fKeFWe/+xeMWqa23OH1v4Xd0wl1md1aijZ0koUbKXeyHYyclSzFUbIR3BZm1NtU+Jl
KoCPXk//Pb6kyk/wgCXDWXWeUQCiE+1UY5V+JO6pdcLuRlwJxTGD8ZGGvH0H0xjI6OeDC7JjRR02
6PaSykD5hQ9SGXbqQzRudLOCkXe0lLNYzhzw1SkFR1wsY07v3CloPBPjMGG0OQFsBppEpD/x0oVN
iw4WodC5q9j7C1JT9b6RkXlwfUbjmhc0BQdRDXrCzwJzUvWMW4hdB7eoNP34qq0Ih0lxStnMJbJW
fAGsIaNGCRt/VBBX0KXfQD6dH9kM3iKKXebzyBt85dJ+fdCdeuFEwTgY4hHaT8pfuZY9fuRnyzDa
Oq2OVuixSif7zjzYvIQ/CPAOBpWsOFFS5HQgfZUCAHRJue1k24WYKV1KwyhqCLn0/JXcdv3EC1Cw
5bFrLgX6NSocrP+9l1EYxcVZahglPclOpQQHs4GaASol8g57dQGzeNfbYYyYl8UG6sb64SOaa7xY
xOCrLrcojs7+90H4TP8xHTnPfSqoxnhDDz7bW22zmQ5Q8TkotGTQWuWG4eDFuGLzg3mxaj7qxnB3
vYVKyz+S999vsUOOz0Ts53ewbLq9rdnlIrOzK/DocLltLUNA1/SNYMOJGzOzw/u4QsiKiZ0mT1ti
3DJFTN8zxB0w8yJXmLfj0KFUJmXaPxWwectRQBx1bR7SgMC8nDt0Ww7G4ETQMwYLMwSfIWyaQ+gi
BMf9IH3pEXGjfKOOEqgqXy01LSJ8+fZdlPo6JEeIaYqEUoTItJDbBPNGVv3c0L2VfD9UWEFINBhK
otOhZ6W3WZ7HN6DOOtdrRdzPdPhASlX8BgSkMZfxlzPUr8zkZ9TEifNREejYBrfL8xBUuQ83xDTu
7Tddeait25QaEQwCZpuqfP8OtT9zRT7+ScUAgN1Uy3iBAprTdk4xkhs3ptNJ1AmElSxgZptryVVA
gAkRrt4wq2pfUe/pKpdolIDB+5XJKMUq67jLz8HylA69DVIMhc3UbR6BXjaKhrFnMxW7US+HpUO/
S1CelRqAJLu+czyhYwVdxNP/XkjnbbjWfw+5avOCZldcebHaVx7PpEQcQxXHOmJZ8kVgeafS1Hop
yDZ+BFcwbDSr8JwDGLxaFLhqZt5A5wFKrPVzqS/efMzPAWk+YXlRAVe4QdyuNbIB4fjUW9RlJijC
mp+ObNymM8B6cKHBv2bvhgbN/+reH7AKKwv2/GjkEdVyQkUzlrxAc8bF+cJn5i1QsNPxMmlF+C+7
myzFzywRqeklZr71wJ4i7Qx2lIxI+W+gybBEZMgf485zV/IyKLdCe17qt1K99663fmaR9tj1boFe
7Kb647Jxb8mIne5Gh45gP/0tCVxyP6NU9PamCv8ay5hfTjRVzwjl0MIK0chpVtb2q2/L1D8uhNd5
XtX2r7oRFw2xCgTIXqOlwoPsxZ/Lc3xi3U6T1L3kCkcibIi0IL5mkCFg9k0Z5jhNmfXbQ4p28/MK
sKxJeQ2HaomU5Sfel5efpwO6PkQicbuhA09d2+qU28Fx/Yr+ea1Tzx4Z3w6qI7wXXXzJKG2/za1w
Ldx/71L3piUf1k+5fDw/VeCEP4+f+BAwoEWO7AYkupr7Jy95RUyTjLjN3z6VZB4rXn5Tv5SKbD/u
4yDR9++5VKPL54tenmGD30iiYZUUFgI73UiQo8Q5U41VcAzTr+BBPB7ZsdyCpfXJjkLC5k8otEGz
gIR5GRmnWHu5ntjMs4L+KK7M/DkfKG0WjTRhCnBCgufvlmAUT6L5BokJFVJ46+kAF1p0J4NQ7Cr3
8xqsqiqnDWqMsLS2zu1K4MjlCZGcl/3bDRuA+mEiWlsnJ57T12Gvq2eMtz723WioMSypRIi5jOdc
a6y4qv6THP3rMNgOBB3rrP09V0jojR4O8N2pZB7r3UoQPyHHT1pA5jX9FUHalp+PXOJcMCiZiNYS
TAESQ3MEJSo7Rtjfd0OQO5LLeWqQaNrHVJvZfpWuvPJEIHSr7g4yPj6tU3uAdQ52Cx0cUso3zrpT
WqdBPV+nK4x6IAnnj15BzTPctjncuZjtEdv+7lauQnopEwlS4Hw9O/VtKQk307N+nUSu2/a8o/aM
56c5k2aLbpPautzSpwnExgqYRf2vZuftbgGaPoNWDivX3cLrfp+uaFno0WnYzbUmaZyRfLJv9+0p
pvcN+5ybpaXFEPNknEuQhpr5JHmbVNU5zLa+5AflVd5Ue3gLQCe/E7ExOZBmC6Z9BuUO7D8dm0dB
Y142ItQDsWGqcA2d9OjN7j8KWKp66DFdkdTBsavlDdfoJNOyIMqim7aLtvxwXNZDmV9t7PTrBPuF
iUsmW5xN5PiTumtYBenihxsmX3gAlDKSGffA9EGlrHEtnQBCZzw8BtldwWKKOI8urPc/iCZ+zf0r
vvFHUTPAqR6c65h5QJ073uO5y6dlmoLkBxrWnCy4JAEDGw81IxqMIX37i5BH16NUhYRH4mBUit0H
VfS3vsY8d7iVMvVxCs/ZQxAVmhmGBWGU/CXuj2RwbcWYzG5a+lJ+69vkin4WckV9YJY96kONGoLX
zy/09gMFWtZnw18DGrKncS3eg654GAyth6z/VCtDsw0gb6qrzzDM0OJdSxmjY46yhbUhhtKTwzkJ
nNtJzh96VQHwbmppeZVYUHm1PB9EZMtHmtTPv3n6BpzvoGrZ2fbHX9el8aR4L3O2qthQNx6PWENN
l3uek2QA3uadX+PtEIVQGfcz01P7r8duLzoLAMcnyN5Yxm+nIelBKzMhDygpB2nredHisd+OxKkh
uW+rE0uFq+29dybVE1jiVSZaV985COlSlMmxNgzQpH7+EDdSI0YCBpZSEdAyAOYg8PtPP8NPOEhx
vsgEm83bTj7fZ8NW7SXzG5+EsLPDLHLPBTITROPaiqdAVsThnBuJt7O/Knhn+097U4DfzELNUSWC
YpD1717mY42Nk/DIqZGwBV4NC+/39h3msijcJJal1l7JNExbhNNPC4ehNBQURb6gjrOkSfREnjdm
RSULZYUXJVM1YQk9HX7uLnoKuN8ESQ191cQckknjmwqX2TOvaYuUSWYzgsQi+sdXMZlH9mMkBgN3
lgEtpvzHdRSig0fE/DjFVcPytNodAibnvFxCmx5prLH+FcD3ryhpmDqRFz2MqmK0J+fU76RPjG/P
kOglVmZufcjoh9jKG41ffO9L3PmLB+Ur0zYynRO27eCjDUkuVZDxBY6TbsTlqMDJ3oM4WnOCFQwc
PzgG71ZGdRFK0t7F+fBjZCewUwX/I6H5xzbwq38gJAMciZwykLRMzSL/YY7STGEq/GFkeCCQ3If2
JMv37c7wUtbSdFeMGQU8cL+5Fy0cUEAPN7m0Chd68wbRyOp9/f4fdp+fPDsFlo/MjxoTAen2S6Jf
dcizubZdrM6uheUIyhQoeAWIBhC96tmIeQyoJDWqVT7Ia3LuhvI+MBXm/w6XiTMhghVWF78GrzVD
Gk47w9UPilztDqeTgJecI97mmd4FgN9NKlmMaTRF+WAHyroncj7fIg6JfPI5qO3v4NjlxmF59arf
TYUQ6NNXZiD1847kkeMY8CHD2nrQnGFxy6ozouwiLntopjo/6KGH+Qq3zCZ+9uM/Glvue9/bKLc6
1iLmND1EZ5M4oR5o4SEhUN7PS5gX+LxL/Z3IxpOCsNvZfAg4xijcrEQDWz+y1HMcGKQrjLcRBpvu
x/7RaZTr8MY1YYbI3JYNKyVzZlYa1KtlyQsUmuUl5LGcM521J/5r17XIfDNnAXil++BZNFZqubGP
iW4jlyUm1+5ja4rUy6px7YU74cWmN+InmKQqT1KSWM49Kn9zcBP4cfvpVG0c/CN3bDNjcHTfTXTO
tiizXRHi5St6Z0fhC7/ow7bPmQ2dMNaT+w5LU/RfXu7fzT18+JteZsgylgEAxddLuCIsWnComi+0
MwgxNPD5+NgZNjgNlfskBZYXRgADq9ApHmZpzcMOIUFgJRfNdqTsoJWetqu4QK675/YNB3zcokFl
Z4LBfCKyKFctorlaOgk8LndS2YFTmtKRiPXJa6A3BPbBEAsdoovpAZAy3T2FF3c3pwmz+5UWf7Jg
BVE0J5v8VITOHApM8+Ie0NEMRnnL6I5TqlaDJe6IBbLRDyXrXxfL7+x6YmtWy6JE39alLdIUa/ae
fs80QIRsLdGmxq8OIXWFKewzE8LBGgy79/VAZrjOt5S7hY82hYxxXF+USVv/iwhYsCdBywWmcc4B
XIgstyvYel3/qhQ5OTRQZLUZywOjiJL5a8xIoRtUOyYgo1NkBkifk8tTawXeV+rVOvy2/9u1uik4
kmwovaMtUTxUNKGDGZrKvpyZemF7pexbbE3/V9KEJ1NyuQpyOgsuDyCzsA6b0HYHLEmTK3ubEuJZ
W35CKcR2NIuMg8w6R2fsvdaB1g6JSAZdkjxwcuSSAY9q2BBfNrLtWVslibi6x6zIqzmgG+v+aF5S
OkhhrnRJGOoegBfjDvmtGAlV3BegKbWdRC61pBWiOaOqw9yXIa1kf9kctsJqLs+81vTobjw22CDm
a40ubF2AIozWyR8J2bwrhd67f5omouz7NVNeD0oW86beVmbW1Nz0yp+g4dmi6dW+ltcY2SUf7q5g
phbhf9mw/aWlPQ8zhypBOhvF8yrV60wofuI1+DOBDvseE/emnLM2AKDtOxgaFBOnklnxnmB1DtzI
1U9FL1/AQK+ROgDXVBlJ5F9/OI+GmJZdy9My1oYa2uAWAoPA1Onh+t2VMVr1DgOr9VBZd8LFuYZ7
d5Mv5eleFmMmTxWIZlnL8h2WsMJxldZa/+yq7peYSc82Z2EvBroj/uFhkWNoXW0J6GbDl+mVtyIF
fZTMSM4o0XQAOyn+Tlqhb4458PhPBNRnlgzUpJVUEReuNL5DwsQp/ib+QxSvwDI+3By39F2lIwK9
KIDys9twGX45RLZY3ZloAH1vwbuKXvzf8FOTuEmYR2tlY0uHafKP+RdBFTL+cC/Xcunv0CcjXX6U
LJH2Pb0HR9okOksEzH5h5/ppRkwcE8eR0RHdWedQy9qayjTsotE9cGlY04sJwAaGa5YNnyZK2Um8
+mAvC02EYfPjlLopoXgT0o5EKPV0eS654vznQjkcLsReFJkHBqrImbiKfQutBmjfqIHGc66UxN5V
963V/VXQKipgFTnKd585bc6ANWg5Jf5vBigh39qv9/bp7XfjcpZ+YHcDTBbIdnWzqHtJMBUnR8lv
BpURzefyxErykoG0g32QzSKay0ekFPtclRXBa6464+mH1+AvErcqyk/q/j2nxWqEl+S6YE5FAkcl
N9L3oEKvUobbmp8rGdOG/Gl/DhRrvbW7koYh2S6XT++1/pq+oRm3wd/VwXJG7SOsswF26JEh8Hyx
vwCVvutN8HK3ifN++y/JVHAE4ix2QbhHEDYRvDlzDsCE1ZverMhIUFLYrwa4P8Pe4GX+o4iEZHrz
wBuKiiJ7rOvEVdyjgPertps+vzeISYh20tKt96h8HzunClRCLU/urHBI+MHoMqkIb3f1b28K93EH
MLAggovM3yV7uZMn37Cq9dVh3j+xUjKfHayiy7zcs033PBl76LMOpKQS/hnVmz/1XuBsCHtjasoU
RxYD8rRWr9WQ3kW6Vnv1v9iCcLV/8iJ8Dy82DW9uc5fdfgq79ChJD6w+4KH6z1q6NHXp6rSoGxI4
v6xzeuJ/EFONrc/xxy9HfeK15VbnIjGMBJHMRuQzKpi90CZC60Na8ZmpWeAOkx79d0Z/iF8oJIdL
Hg2TRLM60e+kSjC4oFrUp5xXRC8XG81uyV/L2W4uOcb7IuAQN1+NwZJ1UqWOcHwRPV13Cb8F4Pmy
35bB5U+U7eUgUwspOxdQHlTCp7HMkzeYfWM0A2gxRo1hjCZ4f74X+hG29bUbaR+iG/afpi6mmULd
vL1LHmAF+YJbATzRlYFxQkmA/QMkoe8mldAJSttCWE8BRN+hXD62w7nY7MPyFTfsmLU/4MCWlzQV
7/GIBt6uAImuvRZ2FwmWCR3+uMEmk7kzLpWOiAo5WdSHLjhGzJqceLlKFRFyFHCBahZUNls44IqB
kbHylCNxcw4xqDYonxtjl+k4xqetFaQhlmyAnYIao9SPa78qImzPlFa5Mx5YLtPaTn/W3jJDK8ey
mFRfUiJE01773r/1Bzk9lYAXJrc3gasj6pffqNYcNt4tbSJsg5z17+2bO0VJCJ+cFQ6hQ64F7XN+
o7sdVJvbgQgRDMILqSMSkbParI/61QIibhqEgVb5Y1mKwMBV+KhOhXMqaIi/ely0Ls0wjVzZoM3C
ksTmn1T02TEwQrQikHwPssOpfz97Ctz8Ba/QR6zsj82FlejlTyQY7zFXFbD1E1n3UJeNA58wpzR0
mSZU3wjk72mPe4OBY9DRGo0YFtW9CRVJ1N5V+Mb5b0Er/Hs7ZxxHGGrUAOnQgGuha064iJw4zWuk
OT5s2dp+dFKrQmMGqdGw6e6K3Loe52Bhcz1MsXw90/JXvYmaA3Fs77d6t7ZYuVfM9FCrj9D2UpE+
rMNblkbIjXi+huT3e2PdOkBC+iMQPF+LpWyDKd0NFCuiqxdYehOOWpZxoZ+lot/rrJOsuR14+UI7
VjpDN77OQByBQGhomY0n2kxbhaKVXrmKuNtPUITPxIXyBh9incYmOxHutRTtJblgNw7KPJU8XC1k
EznbTE2IadmgEfckfZNKcbd2r/dYP9FdSXvrM47sNGHbgkKnQqzr1q2w2K8WXK2qbMGjN/cCyh1z
m3GS+6BMcNZn6Zza073M/cINILyrHMBDrXNpdaTOxggyqF+kZKV+pfQiQuo+FtvaWFA1TyUrTh4B
fpSbI6M0s411avZBvd8+sBvH9KYgjPf6c276dHv5qgQJ9oGRkuHx3OYmj1GdVeFHteVp5mHb/iTl
vhAq6nWsfbPMQu98nYIMVSP/U0S1j4DGKNcfKxDLCQuljICpasQkOghQp+MTUTUOCsTWl17urM8G
A7EATFumKEl2NmkVeuuqlwpAQ0BwpW8ITE9v5n5Ckxq/zCzJshL7wDuGBj6fT3ENVNIBmfmHcLWf
VlFnsU/f61JPVTFhADT5MT3xmc3/ZCcQGU9nTxU3qyNIGwkyByoM75jKSI7QQR9RymA/BQpYwdDx
9p5C0yva2pFtvbmxM8eXec/HzrV0Z7HEqO4Bg18KdRwwxkQmRgEz60vDtHPaxcHPH+PGe2nz8sCy
wa9Z/ecI0ppVopJPapOt3xDxO5qenEoYimsFnN+S4CrTxUis4sY0xCqSq6kyKEcUmjcU5f1fA0TX
ddlckb0ZqPplDUldhZ/QAD06tc1GwurtczryGTrPLUCb2elTLT0VqEWUixUQFGdbyuoU5tliFMGI
SVwS+1RL5MEy6SFMF6CCQsOdh1+RNlT/PbLD/5gI6ff26T91mT7imm66d07CtKuWIOLA/z7FihFG
d/C0qPYYsW7+D6KTVBO/cHhFY94vhiZsAsHe29YaIjJaHjmC+qVDz9Jbqsg/ccNUn/Utt6vGXts/
lcp81eJeoDr7qaXwxUAFIiPb9L3a+9bd6xgRfPy++sJXPJ03+1nW6oIf17FWOHR63LzUuuPTLgCy
X8cykQxbMYcD/+HGAwhXteoEcASyciD1BoFkNhdRcRcTKcssdPbITVwiUkKCHkmuaTfeTqUMNT2v
Z9rSj5dfLY3+zl55ZBjQD86rfsXi4EB3BCMyYv6bDjUu29OnJY9I/NOHXUQqNJEO/Td9mFj7ApLC
cOWtg2dWIHKpURaRL2y6QwR4fP9xBR6AYDOEWd6T1mfgKbefU7H/USbfXY8CunFO5F8AuVYjk5aj
xoctE/x2Aclon3hRnK6O1+2K2dS0G/81YUs4PuOTvTuQQCtYdLGYs2j21W7yq5jA5JEcl2V3NSfn
um0tNRiXmLmmr3T3i+L+tvQtzVpAruMLGiAjK/ClSfHhnZPEuJvlgxsVaH2J4PsxykPIpI9Hu9SJ
ctmdohjH8dVAcEMKbd8Fq4/hBt1nLqquQfggGdvios3BZPRmz0Mej7UsvFy8ZP3vAuRtjvfsPUbq
LPt0loc+1sBDOMr4C3CjA6iwGrnVUaP57pZTReJCAlHwx042aD1KasNu8mGjEH1gv3Yit0MEf0Md
ngw6kh/GagdKqhlr4vjoSuO1wmnvUf05dcwzDJVh6wBZl4BOhxXKERkyNcO0loZOhyh+bRCKTk0g
H7/TLRtYYGGlVc9fSVkYI3SXezm5s4sxa4Ps8w2MAkHBuF39mK1rAJBySHyFkqjJ8fQSz06/ptA7
3v6iXDLsY6ucRRg8oYlBas8lmEx9K46183FFef80bGMnqRfBnW+F1wKK+vhqc1PUF0lG+8crA/Ih
RUKR7Z8PmAoWvZgFebUOaFSsXVejqEbv1AFWHcJ0kHhuOaQDi0HNiTgHunoC1wnUzd+TmJhJcH5L
E2J3yDhhSXT5obvPvDqDaYmQs5gjW8hOJ0FEZ8JbOZcGhq7mIDGVJCLu7TdEBm7rQtEarwx5+8gO
yEEjP5qFJAPLEHNQzvl8aerhBhn3G1rXel3D3SIttCtBCICDh6EYzhgxFAW5XNq0LMF16Izxt5mF
L+HuJ1q89gS5yZKIAzdb0z1DGHH8FoGypqXAgy/SA7a+ZsD2Kgh4tibf5TEZ6wzmQkdeigrkCBxD
BiF0l5qSve7d4brAex9wGB5lU+SdnSq1yWOiX0JO4IuLCtXTwb+q9qzGqP3EYx2i0z3uuFg0o4oz
fCHNP3nHoy4KcDJj4ORV4wNtxatnktnupFeS7Hra8VocsImHGComu9UFI3rjqx+xLOQnT2ItfvCX
63mfw/fMg2Vg5zkmbcA8KJ+Q+b3UrAp7Zb+FqFayAFA3LRR8ynyascCuXKm5S/d/QktBHzFkJOBb
u+tCPn93/qkd6eXg858N8Rh1NhI+1Yy/6l6WvLfSzArjzbc4kAXYGlGmDMcSbuV186XcYiLurvI2
nl1JuKor0+Gr9i1ilVTKt/68p+YCaCSv+acnkwO5lkuWIbK4ReBiO/afGim4Vm44r1yY8cfk8BqS
SqgrqiS8cAIAjhzc7pjYvT8o9+YX6wMmRFbfqGUwCFadL7pZIqb6QY+qHMyfXWGZq/QvLmhB7Hae
Vrj5fDqPSbEineOc4fWQezWcVWEIPHCY92ez948FTDzAKmJXDeMnAJXzaWreGsIreN1vfV4YGyP3
xRcwJ23pXDTlqwhYaVEtT3Wfz2C+oTFwroOt/PtUi4l5kG7Xk9bx/gSP5FiEL+MbQTdR+xWziqmh
SWKyWS+qZu7SRsf91BqnVXGHFOvviBKeFJ+qVLrFhfCmkiUq1pGiRJQOHe+EMhKxKeG5At/TObA8
XwjnK6DhTATu+5l2V8MLE0XOq/OlqnYC1LrustL022asYW8AbpuMVFeX8zIA4bvVvarVELM/KU7l
gvqS+vC44SrVgpi3ns8BGxVuvDXghnAoMkgAchn7+hrlcs8jt3yGt5N7HOT2/6fW3UxkAgPY6Wiy
Nw/Bu8n4FAMcBtCdbAUQkSYkpJwiMpxCa8ctX1HiywYr5PmgE0JEeXd9zt0o6XLb+6OOgf/ulXh7
ekIWuK/t4JhYgIzfKHxVgtaK0WJrHekJl7LYJBeX3NfUcwcNB4HKOCi94vlM7PMUv/Tb+J7LcDWw
f9RGARvG6ISer8rGwVZ5yK3NoM2Z2iBgXjKAG9dD/PplN32L9b/m3tLqF6m/yg23Y7qC9f/R6S6l
JTktGbO281p9QlQzFtp77HsafhKwTCw/cPb0xVOuHEFcQLQgNLnAQPfO5lR8zR/l7oZw0cogOY9r
VMnJ0LHW/fpytHwP+IzOx8N9+B7P6/gVAgOPhNnjPitca//5DwZtYA/ZxJ9nIzXNG/G6GUE5Feqm
l3wp5b/B3Qv8sMTCD9zTqGbQKl/csjDlSX4dc77Cl5+GXAS1Td/Cwkdbh2OG1sSoz9CnpsZKxQCG
hOD8tTnblw1uCRdE7cZsgnqsqsDRCrg2GMOkLWw7jHHP9L9W5Ud1PnhKN+lIfrrZfR9cdOTnMten
y0ji+3A8l8n8fEvYuj9SwSjJTRFkWLM6yzdLLPuEP22k5geghoxPK+enit7o2yQHguwRLgCQUdSm
twRWF3AAos1BxgxsSALD2MAJpjD4Gwes9H/yOtRKSwZxpvCkcPkab/3Bi+GETV3Ys303JyOSEmfU
awK0EMSbZYV4oxx/wg2AoaVhiLaPHY+gflHtnm/IantbxbZVTNy+fQer1WwbI4d4e+z5aAubzInD
L+suiqJ2bdhVBQ8CR+aGNDwIYD4NtswENMhw6sZCN4iFUqw9nLXFM/6CCbY4819vmfygdKpqfGBB
PJaD2BeaGqs7FS5iB7oubPX0QtWpH+JXnryXNDF/ykHN2lhS522fYJxgQATFD04sqRPCWbjo3eOe
3l+1m2qR2orDKXeOnzrhm7EvpHboARaQRCMhJzrrGmslShYvoRv/NS1VLDeNJwr6Zd/cttFOZNJT
DWNnd6V2BVf5WQ0f2AG6/l8fWhQ3sSHypKPw1ChbYxHF9wpZtggV6Xhxn1YblkhfPxkmWb3IvL3y
4j7TYLnT4BrSOpKqvpmKQMQVSujwc6F4GNRVtZSzg4ndYSyep5GFuY1E285/jCyO6u5oX6Vu+gON
Do0lxwnG17Q46UGyD2OIwyANfxR0RnRrOgChWGrz0uinr/24pWVb0/HsHhaM/J0rhuNnRQp5NQS4
oXabxcco5u25tHW7DioRYjeLmzr+f6mQ8yargZXlRUp6CSSqCi26V7q0eYwRVY4dWLmQGW/E0joh
B1AQqrtcqB9VIcR47JmQsazgc9jVvHMbGSVr6+4ebkGjL66FCITutzSPPx44kNfF7jxCNfYaEbkU
SzXYVDjiSFx08DBMxDhJo5U5OKs/tHY/zhtNxg7gqnIzeNTZsA1Br0KsrKsWzY1vi987UEs/CiL2
5msh4NbrzD4KBngvCgn+g/VOy0TvXSFjnpbM+gOASkMluMoabe+hz/LCf2WBs75n6eKS85m2rJ0f
Ki+QfQWxdHr2Wd5Q28FALBtFCL0qrjjm7fNdCeWUT2GiR3O6+XaY6aXha0Y4UN8nsV6XTB9t3G4b
i4m4q1tvDfktcPWYHj1ybDPL8dGAnnopIIZ7u2pmIXuddKW4idIJNEcGbzQu9HFyAgDOUO+pI7UM
2vFzaLUMvt9QqweBzTk+We4NVjuThjszGk5aHPLNxZrloKk0POeNwEdEJWxuv7qpp8gu4ta0verj
Wv26pMIiRRPiwuf0e5uPEKPsRIeK6yGijLNoZtpJ+6THzkqAcX6jvfjlpxNHfjsRILwHFcCoFM+r
YAKCpcSLi2F4syf/pgGFDkDDkwEXtjPvT++leaWcBWOJ8knWJeaXgZLGAqRIV7/gyR2Dqp7iUmwt
/xiNY46ZTMoFUfkN2eH+2t7718lMUC4e7HCC1b+DezjgSThiBVtSQIPdkm7VDPkVysBSs+Ek8ZYf
q4uf5LmznULBEdwZwprGzI5siRLki274E4QGE+thIa+x1+lsqd79jk1pvm3awdIjuTKzGXz5R7wa
QnmYFGGtKVsdlnhArj865xgnIblXo1ad6uXhmNI34cefriJnbZ32Jivd61Z/Yp0iJhkmxwRKfaPw
+F16lI8ejZUwgLYgsPy0vDpsLa051cQGG+Lth0Z+yDIq2BfI5wH1NcMbC6dhatQ0ZyCl+P794No+
xrbFQEOTJkTRGsqc7anqdpeqId+lUeGOCBBqq9QvQd25THTGGaXWRyM/9Nm/YYaU4B76oVvJ1ZwL
c+x3qH0rHAKDu+TGsgAHOxXQgpKYTFV1+r0fON9wft9D7SgwxPQshQtCc9U8EmjJwBW4xwGuCjIj
n9TC1Cd/YTBewLJYLUerkIT8UO66q6XIoyZb6PHh6ZX/k4ILeE3N9snayA25rpANHOAfRZ8Cx3Gd
X1JO/tUcwhyebAUKJbpbybOMPKJFcQ3nU2gcsin/Cy67mguPhCMgsLk8+tzpl/oYTx5YDKqpUJQl
5UohIoKMepZA1QXZMlmOmZD2h399bxMJ6oyfBl7gtnEg7XcA9Ab9xuvNhoDdSS3Y/yzmMWiezMOB
zyuMAwuahDub0w9mnlA+aSZ88Vdfbajb7xebLwVeLscbs7Oqm2LgnxcHNvIwpZM8bi8PE6HISjvo
PoOLT5XtMREUC8YBK2VGVhICtWYwTCdCJSrwE3EmJ1N4zjyXeKrO0ofq2+omOAdFbF6Zs7/ntaNW
0WfibmTvLwkaHKYS1vq7/JpZhQZO2SAvriHbFY5GrRkXc7PFooOhdEXAOHal6iPbCsLt/ll76Ksw
iNUwK+ggB3KR+mJVATOIoJsne+WDPoti8r/UomC//lUuf04gHAKx6u72zsxX2qxFbw8pVO0gFz7f
dWTsrNkhLffRcj+YxeeUYL2DJPpXDjr6yeu3wvTwNrTMAIi43g/3FuiLUJOkcXt+2etC85ydXr5k
tD4WCRVmcwmRy4PI+hot9eQhl0cDQSimhm1RjGL3OVTTELNMtH+Pz6phJgZp3YR5fuULN5Fvj6OP
mapx1yJplmc/QZreM4h28ObD3y49BlUgOpGtgcXSt2OIWT0KEj6Ldqahyj/DqTNg0/8aL8jEmjWT
GZItxwW1pzBaIqMYMY8ThuVZBMdlqXOigNPJD6b37TNIyDSu45vjD5SeVEhH9HSp9SjrxtxurTLJ
YrPU6bYdvZrdGqRFLkCMYPgTPTGnvsFhiDG4W2KreoN+YesZd8n3OWf5kEx9oFGV6X/cOZbFympl
A0lGlBuYnDp8gWL5ClidwkWQXEnyQvYzb+SOOvIOqEsiiIksat9oN1ooHdldAr2hENkJkXB/P5LR
Owrxyi/yzZGfsO6WeaotLbW6ALlT3DHMo8VqVPW+gS7LO72kVzNFGxQDQl9+3mJBmTwnCUNs6813
FZF8Fcy5BYJooM2SKeoZK+4/WnK8Py0ylq7jrfzhP/4TdXfSO9rjsqSewNMhyqQNm9lhWkUnWh/P
5AevMpAPrpVeXvxOcXt3mcVBMtfW4ICgaV0qOVKqqeX5oskKgjf2D+LMezutFysazBuzkV6ax/PD
ip3gID1p9Kfg2HjTFNm6Oh8yJZYXAMCFFQQ4+QUQ50zE4Oi05johIpqcwDlkjoxiKXXq7ApUKeuz
hFZiESBnVqQFIbafuH/ldiBzpz/u5g0opR+5tYjAfEyq54e9pZ3tmRHV1Y17iMgWhoMjgul3xppJ
M3Kr+fskipZIGf93BgL5UiQk2s4412JBtCc6blULkcILDIV/3T00FuVH9hY8WB31JrQfOOXheJWm
abyJ/v13ImODO6vL5AwEtmyeB7d2ScMd4AWN8rGw9WMh1/7hdSVMOtn6ZcobD2TXyd/6dDDBYTZJ
r13YI3cwcBVvnYFU8Z19kiMm6y+OxZ83/Hv56AyQ0LsWeyugIn4EL6bbkxOqxjQT480KyyR0+yJQ
xKRezEpvZ4Hr0N/TZBD8YADb6ZQuikLJ+3gPqRwJEAl1DJ2QzMg8UVLqZJXQlTprOag7jZ0hQII6
0ACpy/knAO58JVkLHfcx+ikmt8B0zRyZAhSfDx7cVGowVHswNW9YQnypsjyPo/ws/2vztOLwChcg
igahMiwv7Ri4mMFdPnGr+G8JBjM9ngNBnFhs1tsMMDblhmfLLfJYBmWWtnAIAiUNV/wUMpjzkL9h
M1yaMTLFXxLllCd8Blb0WGpI5uzyAcavS4NIVSpbmwsW3wqAASn8aa4PNm56z1MbJ9gKpNgBVUdg
chaZUSkK616PbGHQBOAoWl5WFOC5D4kBpAQTdyBAAUb2enbSV86geVDbWaucwg6uAIaZ5s0KB6yw
hR/GPpOEqAb/9NhcsnWTH/t8eQPccjsB/9/e/084EtRPsGaU19Jw96sxjmkPzk+IxIHafq04ZSgk
SgtVZs/TVTBXEhi5X9+zUYZkTxrmE5JW/hnR0GU3rZGYMCDNi3iTWc3TbaOcPA1lEfs5ZZOgfl+6
WT8xVjrcYtmvQBMbPlTO0/n+XNyg8Uxdv0uJoux7bzGSNBKipi7iD5/kU5UUhY2hM2PgZXQJgcnd
q50n+3dnhGjR7SG0vrBymWvlVAr3wgpqimtS6d73gxca7fUsKUUfwhuCOWZH1aRqX5pt/rdPT397
jduU0ftuTH/pllckhctFVuNND0mW0JVMl+nNnyDgta3X2iy5uAbxrTredSZqixxrRxd9otGbNCd8
cEkoAXAs22mn8qWAqNKZOgfIdFso/1gP8gtS1XsD7fItO0eRPQgiQtib5Faxfz1snraoKLCW3EfM
NuuQOKKx8RIUv6wIR8KTln/uZrK0FLADfol4AVBKF54KJC/SWKgz8UEMSHWQqDLK6RE8LGTQ3B8j
+esU6cgUaPEG+X4/jK6/+Q+e6LiPnD6tmvDKcoPYm6VC8XtlBa6CUTdnQB9NQ3g8RwxzbGkrUUsP
P1+S8JD5MUpSkrHJTGWxLujaIB3nReB/QKTDkpK4TtdzhsZ1qrXtMnPJZrvDVDYwjkupYk53YgY6
20GuDlEEfYOnA0YfXBG6pYOwjmXDam4p+hDH53BNuwcB3W/Dwe03t4F+F8zNYQTWsD4fXS5MhInm
teosCmRYR5L4+XhgnXCBDloQmMRz9ChSgLUa7cpMoQgD04U3CX9EQ9xZCLVTnnqpVixB+3tOdd1F
5qaOjH88A0Pe0ggYJqPE5xrsR/DRg5X4i+HFaddIWHbWtU7x/zmV3uV5cy1NT2MtIBNw2txGx7I8
DcQAsO9qrT6D4ZBHWwK0L1orNJtW5BjzTZMrZ604gZaFMxNhKxBebbrnunvrH1IyDTAXto9yG/os
Iqdsq+vIh9mnT4MdwvHV8l2NfSk90RnXAshBJUBxaZxLPH98kIOnylQ5DtTcoAgoa5c4DUAFMaDK
ekP+HMVblGWEuiacGlOkJSeoNnzAFMdPfgYPSuTnR3gYoh8LWaBk3qQHFF/eQ1NRi5UmfEmgYeX5
Lq1f+B8uWdfXWzAbe7k+pqFmQ68VuxsB1FP7UbbTO/UAdWk54tzvZelRooZIdE2avBc7j3RTr/7N
fkDFM2Zw8Rtz/ugEsZ9eKkZMVWLjVZwAnjoUQUzdpKHn7oRf3Vj8Z2V0jBv7c4sidIHSnBqBB2lv
fTH9QYEBrGCZxasB2xgRWQYHzqrQeYb7+zDmhpRAQqDl7NG9SFMKpP9qiL34DKwMD3YV3e5jiTML
golnsvdgQWdhEuH9dE4xTm/DcsUL3fxfPF58Bax/AlpP0Lj/r4wgkCpNnkcjwWfUtO8btbOLmagh
4ehz2s8/ORFIlbn/dypX1zQWv1dzcSasTDuN3huIQ0v4w8bTX12BjGft9xsN/y9dRjbn9O4fUHUE
Uiwdy+5lEaK4zeSr/4M3Y5O/9Q1uy3y2xfykk22TksMAwQw8OvFI3bwRheb1Tt193UneuJ2hPaqf
wHkp08lBMdXzEAInBZyT3yhpKFTu0baW+s4cz7j8riiTkTWoUwaWrQufecTyloS7QYbeR9aNIW29
II0KqE3p/dNjaBKDw/ZZbQzigt1MLBQPkeNQEqJIPqQJBJa2RTFN0HgHhV/mtfr6WCd/JClTax/M
XKDIoh2gbp/FjRkoxtPlFUBC8Zc9zvi13JjdaL9Ig3ZRMjYk2ktnSp3/etaN7mbrXRvTchCtEBUi
ytEqLe4v/FQmzOjALC+C0Uz0AzzBSYl2gICR6L32VSSTx8X4fiFtW3Hx5oIiHUqkTBkGQcAt+ra8
YbuvIVs+7faBB+CKIdv8qZDWr6XT4xPhzvVPT4/2Z+kwQgo/AA7vg74SNCpc191QvKxFImiCg//+
RIjNLHo0zMBFBa3Z8bKtoQ9wL0BYBe+/uySkGieG/icikDU1PLUZ67yP7b6s4u5ugW04qTDghVy7
w3zo+cO4ZGGmtb4oxvIylR0IKebSK+ZrotenUDYMYnYrQjyX4C9sAal7Ufh7e6+rF8PISX9lyfJL
KbXrr4H2BBTcAYOSOkXhGwI987JuOLP8GDGAAFYco8RTUJ6VtDov9IFvnIF08yKiHUc8+vBqGJf1
NJqy9YM8AZbM6iLJQGuMlDAtMYr6F1Fac7CLifpFhDXsUer5i5xFKZQXcE5y5zngad6QN4Etf44Z
QumYkvRgOTDJg8Gslm08mWa105EmPK5Gka/HlI9SWzzd9/pYQMi3QefhFZeMQPQcPXx93TjEQ4R2
XCpyUkmBbqaAswJSTIdsjNMbja0nuJoVkjOq3AVFwAk/R9y6NQuzpfSGGhXec+YPyoWnbl8YSfu1
q5bfkUqc6oR0spabvzUBuUQMtt+gFeJQScYis4RVSHtdFK5k3br6nVFv2A0bar3+O+t/Yk7oNiqE
hdC8Ha2BsDOtoQwZR7Rys1mFmpsghhXd/Xyd1iLdqud1LDJfF/sChkUWlaumcS4jwVanZPPfbwhc
kSWPlKDT73n30IXLEke7ej5TMc+909YFPVAQw2B+KdsLH2vlotkFr+Td7ZVB8bN741hB+exzDujU
GpptPOcUn1vuZCHmPEjSjVm5dVuDNqdoN5edNC8qEvhHCh9rviCR12RHgCfNKOvM7l5fltkM7KZ9
am9QBlr9Z04POISHX8Z5Ce+ry5U8EUlCMFRpj/3fb+L9liKX1LMuiy6v48Xo9hlGWG9yftn4KY1C
WSmAFkv+nvixFmxhA5dZ+HbZ/IaPiEn4J2oCXtOeBi4EGWTRtCeMN9Ib/FO7ReP6Ib7aawChHNgU
f6xgDl1PQcuRwosU3QZsEDwl02/sUpBG/oX5lWf70Q8V0Ebki1aCmwgIjzoC2G440xLNpHTDRdyz
yAX9BzB7wwUj4ItHTM3aX/8pY+dEDBEgBl9yH9vTqM/KKRwR0eMn+FszNRodn8soQPFWDLk8X4sz
0/I9B3Q0kGqAt2VYnGALEJ+IpOsU6QGmblVrHI5dz20yW99sur7E1tWxQGgu8SnFp/JDq0q80LEI
CbN+5P8HFqBFiBrZz+ZOWBD+8y2JQMgyGKwnefFmlVGQbjqU6l2aGXSu1fzXhVq3Wa/XsK5pbo/F
T8RvDeReWxMeguiXtr4P2fpTgCbdl1HKCdXiVOGEnO5AWKcU3eF8528H75yJcVepK+SxYKqZdBS+
rcF9QT5H2Illz/i4MbTfN2S6inrVwe8NlrTji0RI/jkDsLtuuS2rFosPoHpVqBSRPO3Z1/VJoYMb
4YtABs0VblHCsyxsxrzdnjfJGegUs5mocfbHTdYkstlRglV0q/F/5UnH/LICaDmK4H4/knT5VGFA
20oHmj5w5Lkh9Fa1gNFN6WO4/wHrzHMJuL6ZxjMvKqrjf7fzW3rWijvU8gGENJ0GT0ddf6JjXclN
E+M3kiCJPQ1F2Z4b/2NFC1Ls5QKadra7k7GLhMf181KKmtWkEuhlE2Bd1uIYUrM1CHnzI29oaYra
+JNAsbjq6ramy9d2JXSzUDaSSDfkiVjnlWg46ljI0PJsy4b0eupLLLjEP5vkzlInyepEjiN+Kl0Y
oAhQQOHcWlG/Q+ezSN3mlrU/bOpEChIdHWv5PQrEsBUq6S0ahgQAeUUUmI1uYSAf+12ZN0HZ/6St
VPRafLP2YxakyLuLj8dzIVWEDQPEQKjmutVdYFDzfTFB8lU3cNDln+NDXla9hpLv5MizRJSgKBz1
xUOqd8vDnOf7hWfRPaE2Ie5rYVI1nPuGLErwjq6WNHL/M+Jxvo5qku7O/JEzP9Z1JwyGLrxNF2aQ
Jp1rDAe6jYooZ9acAcL3NJq/C0rfIXkRFONdRNe8lftLkUfLrMbUd5XKwjRqC++cPTPgDXTpdAkp
SQZuqL+FTAQIKHvHXiL42JeB9QNBUCIvb0etRwlH6WuLJyDRIO1/C6ydU5nTKXA9vka+6zMVwZHr
ru925FlZWOgzp6IXG43fP4tCgROs8Wo+gfPah2hGHPCpcbbiPEtXtt7SuAl5DvEuqed0CbZ8ytJC
66RWDdOOrDBxEiTmE+etUPpgKa8+1qMlH/+nJMisXcoCuzlJb5iTjRFCLzU0VsiMrxOW5GJOhLd1
Kbba8Et5kyjA5TG2cmCemDjKK72VTFtbyFTAam95jNm4Zdn89zHxbK98yS/x9IBvh1n2gSWpuvJC
p3pPM1JtcR82e1u7X6SpZAbhJX3gTavdqqsGsO7tJ980A0kXqvdMA171DInWPMOmvXm8fbFdtdHM
B8nJkdOFy7bOkvLgeH24/RyODMjJ+vr/rOvaT8ou2xwaoGc1/i/3putfDCDQT4w1v/YyoMmnTedP
49sN0FeRbFwXSIkMLGqvsKcUASo0iPkvuRiYxzwNJkDaSx8vjQBMo3BHR3EwpWBUBa/2coCpqZtz
xqM7q2r1fEB2zVWAnNyLgAWgQp8KNqiNwZ4Wt4zZ/U2tJXqOWLh9AmiV9oNU/PyRpD4XclBm2K/K
8VoIgiuOk8yK09En8jMvlJRiNDsLASDteZuB1NZpbZA2gS0DRz3frv0UeaG5ZVXy8xLKmu5r1iRC
cOtlVfIYRDwUQr6/grO9Hi+Ocn6xy8Ni0nLitTSbrLnVZHJdSxGhZ7tDS/pNOHYBgTcnJTmF7Ybx
qHgKkkyNc/cK8O9kKSYt6EPCflIVktKESVY0f462FCwgZAz9hjVY54AFNoOgZz0JmnMxCDQNFzYF
3GuLDbiOh/PDZhTQT6oMvkBk/ZMz05z+QG0Wz2rM/a8/e8P7bo5TzegrTxYTUKQ2PDjwkvpfWT9z
anUjMPf2s0Jg8bzCyPf2uzBqbQB1WiSIouMGfdA2GSYIE/C1F97NaWF5zv9AE5nITgVxMid9F7U2
7IDqXc3PeDG0I0Sq1WPQCbnVlRibwFgZK+6xRezhVKvdNUByvDVwtLWU/axYGaeWsjtagRSz+OTZ
JCIYlCykxrFOIGMJmsro6EkTJk5SLxyWnQwVGZPoJKQfU6GCWlXASB8HfUPXWqstO9985Oshj6CI
5KE3tw7FPPx8v33VQ1252JGymjvgO4at6u5paMZwGyXRuCh5jx7oqyl65Al4+iTd2KGsmJ3Qjd9L
q9T7OghG+pk2cAFvNK/Uqund75TyWU0UxFGar8Aa/mcK7D6rokT4VRDz9nscKIYfDF05Nd7Nlyt8
IQ8djorxeSB+Jb5qLEpaMGgnf7mfTqQzkaz2cCfV58dSMipIeOGdNdLKyjyLWaC0QUEgh9OFWDOu
Mhzv96GlcnlwM/nQEPyFpdDzNd6cKTfuDTG+AFTv1qJfj2+RPsXfI9mNFdtweIIP8YdO6+ONmVvt
Owm5n+ZddXaHwv0BIkXD84Gt2/lbAP+ArUnOQ2xZHSnNTar7Zze1gZ4cPblQ35mTOUMO2RlEWzZO
v5E8iHggA0U9CdlU+F7mojuVQ48AjaVNvFtnBDKXMZYwGDn5lybx13535oHLlC9BYHsv/Of3WG5H
Y+hqjri0puHNAPJbyDsc8fK3bdZVyd/ZAmUb3d9wIKRix6MmFCiajZJ2pxjO/XXWAR+1Pn51eEwU
8X5H0ksNGv2FaCsitWGCMQfBb1/b3m6/FcB59PqnmjYlrAt6Mfbz7aYJM9pyHBBIKSi6CtuC08K+
HOoOV7OhPfcZSL9YQwQgohfRkRXnebg9rzhQg+ppVcdXJUomF7W6IItt6vhvyg9XuY32LSEwh4PL
ngYVMJDAzQ0AYPLQ+iUjilzbKF9ug4ZYY9ypFja2IuS98sgTA8YpaTxwISZso2pK9jzUQDQDqQGI
b8ZxEd6KB1OXPbVs3kFmFhNfIQmU8ODzCxEunRH+J03BQIeZVHt/FhA5WnwxT2eEJC3uQYt/uXFF
fXNYyOdk/OvKR7fJQEO/a7ggM3ug61+ctzkFOCjffXfg5keQKrdeOjyGfHZzMTGcp2rkNICVPztT
0if5h44V3f6TygQ/44NCPurfHgvNE/ZBtdMlvrvd+gS1MJWF1tq2tSjq5DZbBprvfr1xWuN3Y5pe
pU+GJ8AIyi+JkLtrpUlxEK776fGE/4U+lBF2UhU/e5cKSJ15DFDV7pFt01/yLhOdl2L9/Q++J6wU
/1kGA76A1S9dAzzR0UnGEwYvfn0h4Txiiu3eg6XQ2TSaoEX88rygJxa49Y6SdoIikH6ZDzs16m6B
GBQhn0re3nkbLGzGc35VQpVdGIpc+LecluRwDLaLg5n2Dy4+7RjMf5gur6+q1SosMP/b0hhoQFrW
Mw7CQN/1z7prufGFLS8UnxbTFh2XqmQvi10CmSOCVp2gZyYiZWc2v3XBKw5s6bVA3rLcs6EhTdcu
riY4ie1fVzXUcEX7YxHbmiyUr7VJKuGnxe3yp6bj4ur7vGDGqChybfMsBMWlLexE9XE8hgxFoXuN
jmCvI3ErEt1nKShFzV5gedqRhywoixzWm7mBgq+QoXJldEAqi23S1mPQOekpDNgeQUs7pks7Cp5f
Csltt9tLs6OG/av8AAWTkS3yvGLlmOAbANrJj7aklUTIoAKupr/iychp8WrteCEEFBiJRo3xKjpC
XJi0wOxT5l8qs4lK/ke0XZKp7STYcrzcMBrFTshX3LWmeMNj11Qv19iOWnSMk6jkWNURpVg1tTKJ
02hYCqRW8jH3ZLuOsGuOeyyP2GTEPYKPFBDqdfgSl2J3EOxb0y9AwKSS69WRlUzqlURt/yFgL7n9
UOSFK08/9LJQl4kX2i5Wj5TvhGHSTXS0l7WhnJ2Dm+HAn989k/pdXfyHKbGpHmgwBtzHdYrph4l+
Hz4r1pzjCgps/mFgcxPJ/JGfGvY6F4lZRV22lSjHe0Kjs7nJiH7NeCaziEoy7dbnjoOoT669Gms+
L+LgNPPJDKhAvZrHkHJsFGmM4ojqIRCWM+kxeD57YWR8iIRZTkjjHl5Ss7FMKZBnZWRY16lLq2Dx
26GbMgXX+r24D21pRXjr7RUiiEbxyc+B5cD8FJDaIQkX3M5lnIDmN0r+a5ykzCZseAuN/Ef2WYn6
lrZPkfpKuTrE75N9QcmqaZG+w/K7lvAwoWGAHvIKDjFbMByMzhZd86jYewaKn4xVX/zfv7SR1IVl
4ow3zms9zsMdWU0fN/hRP9mrc58S8sNnq//OVfidyw42kMcjS/Xv/xmH/cJnGSE1kfd30fERQ3fd
cB70ih0ZMs7Pbgad1E1SoGuDmPKDkGzV3p1TMcbgwxAt8QTW3kZkHNc6HbKlPCIWdDigBV9AnBoe
Swxd4jCqZTIfBwoBe3SAaBi/SNE3qcsnofTPO2xyYjrqxqYllDblM69LY2mMlQhC/vDrywewlOlc
Eqak7kPBPNgLbyQ1PRXRJI1hPq26ZsEjq6NDFiza8UV23CTFzKirD5FiCK2VYduQHUu7tZqhWEo7
Lm3EoTbIeYUXyOnSX9aKTgaoTQeEx4ixD8cLhZ9odUF21YTY4EsDJ4bvCIdtdP/4Stvr0MUQ6QNc
cc8akXExI+Uo2O4J+5BhanIEORouB1uWxLDQyaFQ1T6zw8+JxnSiBI3op8Df4jvmjsd/AVwBKHhT
yH/jF1f4hAyPYfseGGBQhASx1YeODmMELYFadcFMUyWgCORWrpwv7fn77hPLF5pSW41Tz+BTw7RU
wCVNcFuc9p9v6ydOZ9gYcUgqB8uC+xbHqlYE7I79F041HTJ7gZpajui13hFbuq4I4gkIjDlzbiwi
lAjme60Dfm0KMpYlBhOTLVDI06JUXmHMLxgyiCyxXfUEob6HKZU7bXX5BcSyTekxh2PaaDHjP5Ng
v0zxUQsEzFuMUnqm3YJTiKvhuy3/hhUn5dgmXAd81Odl6x8HVjLx2zCThEUwcH+m8Q9qTpMv2Y94
yG6kQogepFvTRz/QNu56l4BWraHn0VXAOg7T055ZXytJlCo3HERUIQCyeoNbdUqnhBjaoCycgtfB
vdbsKonDRsgWZWzT1Wtldmioc5hx0SdlIZe7DRH2DqveDQU38NQeoFs1fyotMWB88pqZ7+3Yv0pA
cL/xhksbBUkJqjPWw67TkxXUr86/ZgQnQ+NC0FoEKgCo2HqwBMIFix7lu9rTBuM4MC7mr02GrzdF
Zm8v9T6OyZzHOH4arbPdBtAvZeq203FleRnKvNE5zcdjnlwlpI/uvD3GyhAatm+9mvev0mTFz2Ep
YkXgXOZy5po2WZjcTkjiFlh6c859J7CTGgXequXyEs5VPZzaNMZfuXXpq+s+EtijFcrBAA3sZ/Zb
Qj8NaDb/HObMDfePEP14UdoE/oJQuZ129WEqPNOEPi+xepj7K09tfsQsnl1rzq3oC9b3EgjofkJN
wHrMDd4gOOE0TsawyV6gKz6EB4c/nVA8qfKg04hN478vBRGJ9+YCIDKr1R4oTDeaAmlivmVMbDlP
05L/Hw90qzKtNPGYkpIsKhQKwVwdfVp8wTWuNjDNe1DFd85Dw7m/8oM+18Rc1oCRZXENsOueaBeL
MOeVtBHte2C8HfuWblLGNeKE3ZFmqdPRlUCeFGUOaZg3Utq51pMw87nmrUhIQi3ARQJOMd5tRM98
7LFVABgS6fYdyIsBi1txrKt6Yqk2/9VvHhuqsIFcbkdUAEWK6SxricVNmwTPCPCnUym7miEHCn6u
a+QA4Ko8Mtpbff8mO/pB6dpSn8VZLB+mBF+4gY2ozbBnclF6c4mzVfhJ30dQAwZVlPAMZBMbDvWX
5n0NQKQw2Pf8n5pKjnSE/1UOb9/jhkRY3EJ6EQ/e8SgvpIpwDaLZn/jDkMeXGAm9BHQHqFDbY0Za
lLD5tiMBRNLSDEaOo1dyG5Fhwhl0ncEiLqEUk3lNsOBHbkX3IdCRyiogySh89iJciTR4VhAang8m
0v2puUJPpWeFdF7d7LrFv1vd5qjpr5pl6tFpDp3JTYQWYPmRDLjofDy6maSiNwhDBrAal3pzW8Ni
R+vGfqB/Q09hgJbCXB3xlUE/Ak1mIskYCOBs+ED+HSyh9cldiT6W+2UId8my3gJ41CDtlYTSnIwI
S9RcTrrVt65TXCi9dl4zXkL/YbVKjV8fi0kvZfXxxnnSQuSCTjWOhAImnUdsQbmcQufSS1OlV178
+c8WQWx5aNXoJGVzpTLdQztnAxp5iPCKrYDQAVTI8d8uNVexKxxNL/I6fJKxio9DXpPgyWM7vFc8
FUPfxlHXS9RKWoQwwjl2YNOg11AwFLgKLmbPheMdwCdhQR141oO5/MBhMQz6X2adnOvYRWGipsMM
63J5zzVK2PTs2khVv7uc20nSmhXfcLNYXaNQ1XXPawJO5pDL1E1KNWgr9tj/HytuvGYiw0FHxx+L
ykdij7dKvwwOU2/Gm8Z3D0heXs/cYtMu9kvJg/6fybnDgg2fYseCHKCyiK5duvgoZ9kFp1HkSqL8
A5LodgpPkN10K5whUnev86AlzhkSidXWRZkTZfxCJjawUhowlLxOzqEkoquhlMQGPo30cvzDe0JT
c2DyBfbzIN0tdOJt50KiJK9d7HBs55g8bvcpu5inKMPjaJLJfRP8fhJ7vS4vCnoU0/BQJMjFFcfn
mrS178NSek1ZsmXVI7vEV5LO7uAdz3V+/YdAZQWY0tITMIgEba8q/vuIcUXAUYR6wp9mGV6trq8R
ttUVkGu6Azy9YQbRYaJJwkDZHYKIlQT7UyzQtUevBCar6kXMSy+AodUZb5RIRXK+V0f14IHfDmD4
Vsn39eqRpKS9wFPPO+qVsE5n6dVNNgWszs1iyBxDo+S7TN8L1omKtPw0I294rKAO3wtttESN0Nbv
P2dDlkfrs+2Zb6kBnKPuSH/EvvvTuXzAuOzFHHBhnFD3Hw/Nz7aTejLPrLI63yVWVQZeAG/wTWJP
6FSuDFm+dC1vCV1K/3qOEBWEigNiNTw9wtlBE5nqq1mYe+rczEYJHTChVnsj28Kcfj4he4peeeOH
QJAz29kJ2tSQlrblQwOJCtBKGrrKbOh0kc9guTNZi95SB9C2Yidts0cnmaLl/NFzDQlmpNAIlRjD
i8YCQe8Hdrw+muJ2yzUsjP2HESTA+QfWm58wNIzLpQenFL+YIO9tVRkze5oOo9NMTex/XvAePh9s
OTYq2Tk35nO6t1sfrChHJLO5ZOak+WNCLAB8SpEPmxRcj2S5SuLrNF5IT6uNVmWwy4M5ptpYndFi
3kcFl54yr8RUyN6jDa80MCTsTdXhUjWduyl7T0alzxmrd9P7GC5jv7mqNzScAtNpPRRUaESHR1d/
NYuWgp0tPXWU591stf0anKPhkuWXbJXOlK7mkcqNL1tphBR0sRn5S54/Z3YRddSl2De6QRRzfOmt
otQW5iZFCmDfBV/uVXtcRzUzqieTnTUYl83Osg05boG2d8KQ6e5CYn7wTb52zmsju5b08agIBXSR
0DCaw6JQ5bVPie0i/fn+ZRSlzlAAB4MKrURTFjlSq88klS3QzomC7bZ+UOCk9KMIMzF8mXS5rbRX
athYeoZ/dkfPe3AB5RNx0R6xdrChIUmN54YN98fouX+iZMrsd8KZrXa5h9RMSmCTnJ6Sbr3PCCWr
Yj+8WWT1mQMgbedv9NlhEDTThQUtQPHb0xZ6Gkil15jmFl2Yk2LtjSIfXwRxVqFmsCyOkiC4td43
zYLMmZJ2cbDVk37qdKngMyqVc+6R1g7uHzKP1rOVbEjpU3mIGmcNizDE7mtNjKdPKlTGwEABdyIF
iayVfQpcdBXqRqc/9QGjmCox2kEOCQzCU+yApzXbopquQA8E0HNQtxzIQXwta0Ojjb/0nRgQhyL7
bppZapjLpIctXJRTa5c3M/i2rObxYhqSe0pnmG1hMpAPOaSsNEI5yWOML6ZsShlVq4sCYK+Rt92k
AYZi7bIb4I0MNo8JUCTRAwI2q52bT4g15jyStISc5lKnmAm/osHnVukr7PcJAno5CH1u5E+1W2D/
1KNlMDvOycSiwA9Ddlqev63fIi6q3LrOwAg11smGIYxncMMfAGL7jkGsdBgF/GtP1p29txrhegnU
0HvFkb3216H88biRSNqOD8FPvxs0HYQoxmu0qL6ONI0UgPgkK/9fvTkbkiDM7O50jOZOzL9KbAzq
nhDEYUJUEx4llV89UwSSlIhnAnp2LKCQ/Yi44MM+P/fmnQ0BQLMhYGRHZTM+O1n5Nw8pDvJR/GDT
sxXgyU4C5F78CX9ZouB41KSmishOdL2OsVlg2XvhhY4kPltGYQoaOugU+XXUB9rurJqQdYPT7MyG
Em/X4kuxGDUq5q8xw1aWdz3b5rYJZQ0nKImIA0TU9QVTXeaFXl3/Hs3VhdIpdZmc/hXD/ejbvAC/
QpNHGKqvq0eQOx6REeAtgUB4EkmPyE/twc4CWcBngPtf+SdO/Bj0xQm7/P9gRpLjI8/Li6IGxRvd
RQ59uBSAfiKONMm/HDlyhArRIVAKNzs9yHu9jl4exJOgIlCkKf3XpKS7YVk4HhLl3Ju8JJOCuIwb
mkHnx8InAwOqbTvyPiwLrQNt5OXT8EA8vMCu3l0OYjDVy/iNhwvm/3WRLVxt5Zy0LMgFGgKL5Gqw
h7+TUGW/2cEqiQd6K5lrauBucCYAlQrKvlPqDJA6UfM67vNVmYhsNmTmthwRoguBWhO5x7C4d4Gm
pSUOaGZHD+5Jd5BTpWaa14C+tGvwcwVgeqvsT5RnsXtlkgnVQyimwS+riue231CtxYqUS3EdaeaD
64XWoD/o3Sf2EAwzcZb8EIr+vJSiEppS4eolvkIpWZOTn/+yBkv4CsBFoURqZvX5xilZMPt34RWK
8GYDr49krdtLF+8xZ1pqzWxTw6OgtB6TIXben0SCz0u/4q4u8J5iOsA09bJmHHQ5vXbpMhp/we1F
tBTCacElcuRktsk2IvA4vXgBn50mxtjjOiP9AX+FRZ+7C0VsCGoH9igA17wFugWXm8lQTggpXGis
cb+/46C9hxh6RU1nvRxTzaMWa9J9dIlfaTpSmCGI1hmOdmE5ZF0LhkEtWXJs7Xt9L60QT8Hcosbx
SCqD2CwYC7Jpjb4opTlvBMbiB7ZkHL/Zfq7rctSn4SZNNCKYWchXnqws8BWxZaeDsnlL7RXZJq4M
nwpQJmLCN05aL6Ks/rMOIcSL6UMCq+fcoEOw9YtiAp2mCKB52UKRs8+3A3m4c43NSlc3lCZy3916
oMU1pSGd1pfVli0O07F33KtfdAe9uXv3aSIyjRnmrfSLjQ2fnIZM4eBm7xZp7Fo++f9ueiazXqMB
Sg7VXXHn8VNKCQnvJ4jMnhO40lP0iInsRHxjN0samfVm+3r4x80KsXNsWRh2f5GPM+/FeAHF8GH9
9zfGjdIH5Xw6oSEDwZOG+WhexXNpkF2ULRPd6Eln+dobhL2gESv5AHRaBkmqp6Y4ezWSMwJJviGO
UuciwhFTtug6Zsq5yF5X/rlUOprVOIQ69OCKavhW8MsI0W6ILyJImplG5DNn7xQUyur4L6Oh7jQp
9sclMgxID7y7+2ZqfegZcqn4cDegRwui27/LXDp6aX1XEFC710TMuJXvPPAeP0wSvNov+oBLzB96
lLnbJQck2y0qXR5kdtj1sVIKb4WfDTloxbGIw2EoSw4gUlKXWAh3CRx808+/ozoccrEbI8AG4kod
jXjeD7OJpXPRndZP347mQHL65a8bZftPkaqc5zXLTbbZQekBaXF/zB4195H82bFem8x8P3lteqYr
R/hqV3mfs3d08FNnTyU9eRHYWnLTvnRG+Sr3N7uhjQ9bmofswa2IqVaPpvZ7MZNIIucztRnbcLIJ
GfxWjltWuS+7yxkz6DEElr9zd2JPKzExLKt6xusXeVynDNZscQk/Qneq+wsPoSBW91jUbz6HbY6n
yYO1chPZH/f2SDgw6UmzshmTWB83Kk/zMOIjq0pSUdck3+RrG2ghoJVK/1V7NAhK8Yu8kenzCF7T
8WOl52OcUhZxsqpwcjF1YX8hdPwyaPrgFpZXF13S7SE/ApOHgNHaaymAhtgbQlK8nVeG2cPgIjpT
WVlSdtTZKs0BpDViSL7oOy27472kA2XvdTX2XVp4Hj9PTm9SPvngCuCVbm0Fj46ss7diW3zlfQ1Q
xMMGw9rOLFSId7WbXiX+FVSreDUx9VaBR5WkFSY+IxaWo3ZEntxx8NnUQCV3OPfbkB5gPIgfzw3D
o0rBeekrPzm1P2YUlRiEz/EJE+YliZ2kV17rQsbP0nreCB5bX+CBeoRPHBeSHt804mWS6QQ+nRd2
tn+tZ2ESsjlpIyqVCzhZyWPVDDNFqrDqOOtNmwydC59eFYZzuuWveC1MgWaTn3boOV3uXdJcjgPJ
a6QUawHWuHc2CuMjazQaLhepZrBsN6oNAfVXfnIfXydwk8hhteJ2w+YIZnp0zKmQ7ButCi4KaJ9K
LqxHuIwiD+h1AScepWKtevgShud63ry3MVAso+dqw2VJMRRrYBxj7zTtn0qf3EoUWYa4eVhJ4IjI
7yPI5WfZvUUZn2ZILPP+bwN5dU0Mw9eO0OMczH3zcrnYzUIl/bbmlaaDqtRy1tUWejiHS5riiCaL
Lpwogfrx8ZWM1VHdLGH0aHvwcHg1V4JWeXLo87ApwbrlWLdo89xMw2UTaOy8mq0aROrV5VmxEpSg
9eK+MM4HEeK1TvcuvDJNiVMinc2kqOTV2HEBcdr6+EAk8QvXCwlaDdErNEYWnF5hYeKGaPGHOMK9
s4ObjHsSAX5el6rMGgkkWxSjij5kaOVaed03v7aZj86Y57CVy+TCfo7ZIs7L/Od28slwop3f13c/
AaWMvJegZHu0V0WHEbQ3QXb3H6AAydZiZVSH2++nUsAeZonRw+/Wvt2EtGAuJs/mFdcy1DtAON4l
scXdv2uKq4lhL5IPMKQu6S2w20Y7nBioHSoaweO6BDCl0DHfe4JeUre0+UB0xLHHW4Y9RNFg5aXf
GiF12gg7Er9caMh8UJAG/vfudKtUXTwciQbKK2SSbWNLPJ4Yc+jgMgbmCMKYtF3W+an0hBrfg2ts
iuu3lWJP5EJ+gnYpdcSDw/ttcXRzmOQGp3WoaYuESdPZL8dK4UKWtH6u//QfYMNb59ARolifWryC
N5/s9/WT9SMG5ky7T9QkiDWyI7eKaq8E3A3UgzeXrSBplc4FoLryx9htJXpuQRUfRq2qKVT0crTz
9KXtEKfBsJWhM402fJ7LxWUx7lM1shdNPMr+7AshPmeVNb96hNG1Pz0HXB2+XbZfyU/PoHWa6ekN
3cGl7bR4ulyCW0Ra/VIFqJ92IMAgdWjylXyP/QnrAiMxEUolQAmHk06Otwz7cW3s7zTu9nW5sNl0
iFmekLZ/KCrzrUdRCid85bqJTWuddalap7AWUioFjlGFjBHhfcTZP5iqVw7J/BN2FVXHmYoBPBKD
yS9KQ5LNU4KN0shMrWVr2iJbmYLqpuYXIsL58bS78AyYvmzsY7vyhog/reTYOL87TGHR9iRVH0YE
I5huR8xrVVJBL+2KnkTRAD/AQ892rV/q4xLH7B3EOtk/ow+Gm7HZAHZmzramirlnqreArICH40mt
2uU0a9Bv6zclCyMJjCzgtYshxgB6WfKtYeGyE33kpL/d4eqIV3z8/JWpbqk5gNZ3mTySi/LuDOCp
ur/ZP1AVpB/VZeRAxE4jkMXgFjrixA+ACX7n/2T5DB/u6UfNLM855RlW1PczHIwfnmhT9seKXaZj
Zd7oRgE+P/Q36+cOwFT5wYAHUKhwhN5RBr8cxt/nbscKmXhyaCep/jGR6yZ5Ve4jKSq6+UIT3M4S
trgYy1HvptYjH3nQm/DrPlSENhtCr1ZNX63klybvKgeRcDiLziHNn5C1dbyDceT0/vwJaTGK+GS0
aNuMBDIghasieJ5awPgN8IZq/CgqYUZ0+j7ZU3c7ccw4SJiIV7wE3BtCrR7/1sGY+Aus88DRoDkz
INEo22PQA7VypEd4huoB04MF6ZiHKDpD5kAUMnKbvOrdoR6fT4fpoMhpX+XTCvaM6aQoMlogVuRL
vY3YaCocBNo+wfRjgdbgQTxbTVlKp+2u+ByqHtmGu5RN5HvWPozHiQUuEyQTClJVM1xcfahOCzwW
g5tDA1MYcJuJ3fs9kduYHg560u0AxnhJB/KOmPNm5wvLpt77Ht6MqIlWRbgv4NgdpX8RB/ArcHL3
9cqNH4FUPiOBaElA2t/oqYdpV3401IaA30Nhx1+t6v9C+Nk0KfCJme2iuicfgMTq3Ewx/H9O9WiK
1+twrAGxqiWAuY9PNl1PVO+1Ro0lsrRAmlPmV0DON4oVYTiZV6kzW1dYrEuV5ArRvciTWYKS65Tw
FBCL7Gji9+zS5AjJ/qHwvOIWP5ZOt5AK/Yg5ZfWaD08zA4ecuHhq8s9xSARrGSIV71MnlgDVupul
4KJRrbwzAybWuED5i3VkwAxkIyBco9RTFCsVD5JxdSh+2XWtviTtin30zoWDsdJhIAfte8jLzI6o
5kuXuzJRhfe+okqtBbCY9fnODyykpI1W+omiCDqa0Jojw+hxvvmnifGhFZeSb3HAd5Ol22Dq7PhO
jK2n5Am43SzyphqMac7sBOxjcPTPmjzlwMXPbUdJy/q20j0BHQFlB+7TbDDn9KoDJ1vXVlHqFTpc
it3Wv/rudE21Z1ec7/onxm8A3ThRU5HdskpuYi5cDrwJd65QvRw96pHTeOfVVj8I8hUsoXYXfqcD
Qxm4nCaDEb/gZyFkmYH4eYHDsA9qLOjS05vGvJXWuXIdsUpkoT4Ey1rN/7tN7/S/hhn3yaE/Hb8y
EeVSTImdoHBeY5dM8ZrF8cUUxKC3W3b58Xhac2kFX9XNt2j7wCpxuJXBz0jGZqkhAvjTIPjFgj8u
fy5t5k38tLhuwAbpcuw5jrnWV2PDRi5Q8rFMWgJWLXCzHqNcXtREoxj+/MmPaJ7VjCMz8VqvXEmv
qBVNAdYn+Tld5m4C7B07ptA9pWldj9uaGNtbc84KP2KJCjg9YK1IrEsxmo+kICMmyVD9snhrWHfE
x+wllnAhtJJNbZm1vqPzDjs6h5+L/wWIgK5ntOX0+oXg1bncRhXxjvuFoiXcIG1Yvn4Fqavm8okg
AA6EBMMQGkdr4qa0ccFK4x/t1duIqw8U8bsTKAoMfufgBisICqiMSRkClnepmaMQBCOyQDAISNTf
IhszAF+ACAcWDDXMW7W2xFleaCGQraHM232tzjLvUDT/kE9us9Pkfma5aqcLbr5C4xlguwBUhd6C
3wBEq1W8MVGZrVK6u/46Chs7N1UB7zLN7lDQgLrPwXoYFbaQ/ivWzFs5L8xK65rNvXVsgOazgmnx
O4Opr5i5o2AE2317TDQrVbRlcOSIZCAVL3smEghCZP6wFgKRchLjfx2ybwDtGvcz6j7Bny22JUKW
v3Rrwz6P1Nf3WmSFnUIojts0RNEwfoDzoTEur/qRdamxERZHSACmR+9+1dV+wn8cj/oS9/iGzXz1
ys8F1VGZkWArURk73iKGzl+3rWg155lXZB9a53gGYyKTn3ZouTOGrNFexZrqqw/J/uiCJQWx038y
qRRucxbJPRkF9LcbvlVqcoDQBRxTYXJOgz41BHOu0BffY50CWKxyyaNXdhqfQAGndbjBDZo6Q2A5
1TWKFiL4gSZbEqRs3b7e1+3mLM+r3PcAJOsMJGOcYpDD9dY3Dtjm97PhMz4jvgjgf6GYjlxIUWpO
d2/Kh7JYsG5WQKH90FC6I9HFmqJrNS5dZbO2ogV+wlVYvfrn4iUvY5MDQv25h1moQH11EqxzlKbd
iqGBIuGBsNA2UXuHNQNFOppVCsnKi/Y5oZrIo4Di9CEcpMPTOyggCNidrgRO1nsLcfmLz0Ewlodf
HxlAgVK31YjHypoNVXl42S3JWz8dINinLqzTmqK58qF+9A8StokxvEaGOF8gduY5M0R2S2tDxa/v
5Hz/i680QQe2FcG9rtXWBjLJQ22sZFHsgTgA/s0QxC1hFOWdFt8oCcsIb2tpzJJ9guJ4VTP2CyEL
8YfK1jWWiHIVZPqkdB6dhVBJJ1ABYmQtWlcmWyW0bakYHwefbY0OrGWbM2lRPjvXjVkckli70pMc
erSpIw2FffIsSfHkzLDCU5d5urgZ2aTlja/1/C/nAsepbfhU2cohjCZCaMmY9+H0+K0WOF7nQSae
vkEkmmvwHNz2SJ36YS6U1x6kYtBnzsf+ahluJ9RiQDWbmIXNzeW0LPBPIUSexCrXB8Fu9nQEFBxd
vnBw0UyxTAJ0GMvjnqnA4Zs73dDbbmPJnVnF9Xmxw7LYS+k2GEHaLAa4o+KYodfdWaxFKW/mDQuL
srZZggzbYP1VKB78o0nnbIN2aD2ZBPulEe4exKcezonX3xqoE4abpzn3uNnk12pEXJ3M9/0Rz9Hd
xtaBSKsZW2AWfRntzmytdVcvbOtCE1fcRUWX0JFdL1gNd6ASzEyUdTkTWSmGAi3AkYsrclyXQfMe
Lj7K32pn6G0Ov1+EcptJij/rw/MndgVWeQPOZEGjChLoYIIlxe6hZ6Mfke3FTu/lgz/Eumf8VeEu
cYwgVV/KBgtChqXGiXm8ji/wqLV6Dn0zBj9lUi3PByF38RmBXXfS+SUxKFWJkGARLiSJItXVPSdU
na9uYKi519MvZSFRaN84kRIAodghl31qJwXW+QD2F612lAfhi+dcD33FDuIWmlnMiqV7dwhCT6C2
Cf5vRW7DQgS8K/hPsr9yPKwMMoww9gERPlcrD5KHbF4igxvmyIPTRiTSM1SQgn2fgYjMRVagGtGs
NCf/d8NXwO1fWIkCOSgu3Ks73SrbwfnLFJFbvtOsf1z8YW+eU6L87keefAAuXPhLQptI1ZTZKmDp
M+jQJHa6p+Ieu5oi/Qc+UvGHU3whteObp7NiKK0FG1Eog3E/L0XTqK+j80jrcmaO/Z2tdubM+8rE
7G+qZOiQyEQohtA7P474InKY0htkztHid1M9mTHrbBLo+wTkvkbMQ+ykQXKqQy7vD2ZnvvFp/FFW
BPecmy9eSj5GbcW1HBDNWlI9yVffFmoL2wvwbUY/0RPBeqnI0Ey2a/f+6gFYBP3rHfptLQoiCc49
e6uOE40gu3wRQ7VEr1Rmsi53DYv19p/mJc+I5Eub2g9h+t0EYY/zDu+skKeA7J0GMYsYXjRVv5jz
jH7Cxa0YS+GKBA9rtpGTBuDmEjpYaVW45PgDAeWRrwHKrLD0ypGQrILGvXlT2EYY0yRspSJdUeFi
IINWTJsTv2NlxSlnO7oJjNMCG9kuEntJxHTwXiuO2vfJ/pZfpqC0MSVYdZG3edZv2dCa8DfhsXCE
/TGXiiAZ1C/kp02sr0yMexMkO0OpWYIZmJW9s5L+G7ewBCcEkIu53Ahksk24eHrA0zL3UVGgkSPA
kZlozu1yZkHqew5Cs17xr+Z2FdVzKuO00ZscMFqZw7IyTbkkuTR5VyPRiFbVH6ZLKm2huW5nZp9F
YxnMJ9idNY8dUd0M1gb69OQewcHAfoH7NVyps12MfZZJppCYW7Dys372BtbNN6U/VKl/8/6oqUuk
nBofk+c1NAHeE9ZAVASZjiwopbYI8/hv1IvvAvgN8gNvvM9XswMZMWyleifhoMU1pxys4EvgvWRt
5U61ocsJX4JOOuXr1TnT839l1c74FhtXKLKzbwGRXph9xl4qHtJaOYAKvN9Zct3QJi1UcrnxYhyG
aUMVcy4478AKMTCqy6FgU9EHXUQs2kMF+G9HcmJSJZKMbdO7q8s2sMSif3h+q98UuB+IQepbeetj
bW6nvEqEt5Pa61PF8frQapeCtu/MYSlJsGye3VJNCR5ZcIabi7CF/Z/6N3vK7y/3Xe8diqv9wJbp
XB9HLnpI6j3HronMHLRqBiR/Po1aCLhlh6nVq39Pqg34kMpTIM0H64R6tb4pSMU3wG7n2zn25IW+
WuqjVpSGlwkQKiW/NBH5BFWNDC0DZnoiu7GXcAq8fCg+HnhVYgW06xyMtP1yXoh1cNYdrQBi3fAG
Id+xFrGTu3l4RAggQ1oNjD5fm0Txnkj8aTtnH+jxmCQcBF7W1XQgUObq7xJsocjN5x7Hk00eT1+B
zV36VQKJeYoFE7vNnehZgMAf3Fj7H4fR2qFIdpmUH0x3RZw2/Ls8VTXFrQdUH+lOwd6YIQlfvlkp
XUUBL7Kk1ijz1kCwFoc6InP6Aa6kwilMvp84lw5yDKzABFW4w2inTzebcV7hWYENIEhxHyt8+MkR
vsPWkif1HT0lkksHk7Eui/LDsl6o3kyxtXVmY6KL75g4WeYSPlKfLp0PWQ9Rvfcyh7uBsRPjkfM1
tyCqeEMbeKpFB8fjsU781v1sFq3APNQuEGYiOH8vQ42HythmmTU44Pinl6+RFjvDubFqvBnYKZO8
QpX7bsX5NiFWAkRU7550J1lcKDADIWm6OxM7ChWONbv9aTSZCS9o0skLwTjbku3YpxueMQu1V0Bb
ETUWsLnhzbeuuYNZaJB0Bz9iIQBRAZkecpMkh0g+KPVh7BEMW4JglL1ozPJNPBAE10dV6KN2O+lK
RhI/0go9lACTSUfOy0teK1jJMa+FmwIGCXaB8L1J5AcP8ScokDQTDvWZeR3SxILToeBrMFEvNOFY
m7ANCt8wgwCpxMRN+MJjRw1/S1v4kqha3XPSjShN4bcXrO+/vlREAQL9pu2amnbZCgtpZt8dgWhs
cwGrRZzvHSg23jFkHjhgj4n3R+huFgyH4WsHYhA0unGOcHZc2a/HC8kvRkfdL7UFgLkxtzT/CjlP
EmeUCwqQA5AkzFa6N8cm7ZVeZVVHYnOXiDn1B8uK5rUYFDm2NjMNpIzZdSJH8PT3avQbIcXEODLu
652HyOjepiY69BPeVBSFMFl2xpXFDFcg60cJiZU2adO/gxIvzzQXoVvU5GeAAEA4gr8j8hM/N1tW
ehn1bwrt/p+MDwoLxfw+511jg/lqs0fbgEsQfKqKiVPK1XnJTy/mWmiXO5jOjgfonzzPR6jcyh6G
SRzGALy9aum0mnalsdwILPYd5IpQj3QuClBzo6MxsrNIY74eFJVlxw8NpOBE/ppD35oPHKdpldmb
4I/PUSZ34gTnfbjgGt4xsksFdvGYbeHFBfAs/L0dmPhG9IxmRqMIF71prIpv1+GRGCkRGmXG8Ysy
DCSPzjXNL5VX1ybmYabLX2bms7qZATgymT9RQQzPNPSL5GCp9ZK0JnusUlwLJ8ha0UpxZsqy87a8
egoMw82ae1CrIzwX1Ou427J7a3TaZSOQpAhwdUQg6d2/z4qh6ZwLyg0j/rNabkD6F2CFsaCmwIOF
yGpvFJ3jof6908YOI45uvdeRwQnwRtJTGMfhtSFdvk2AYthc5aur1VqrzeNd9C2sV/jar3TC/4it
oVa1Q7N3SWhgLukFKVLFQ9Uxm+bFYYyDahngYHEk32vrSLzemGTwtvRGWZdMCcFLFJ/YVzukGbzR
063cTAG2Rpyho7LNLhkQmtW2YuHFIsyRv4rbduVPoh8WC7MI3IQdE9bpgUyiYiGxQNk5SHurd2n1
AM/KvLpLaardkM04gqBKkQnmuwLQTjAXPG4E/RmBZtodiS1AswW1cDIKOoFN1ZPzl8z5fwYfj5Mx
pG5hzvgFwatXpks9HHOFxb0Pw9n1bWmfMJ9IaY6hdI3UGTmkpSv35KRipHny9Sg2HcszbE0uyN0j
czeBqZF9Z9gu1EnoCjvi8afqA9CxWFOrnQyODGTQuQ0dmdDMTDd/Z5uFzcgK/yoNgZtPsekYYwib
zn4BNLLfvzUJ6GWdmB3l+XTfqDrXMccCNbI1O5VYl770/3wLQeabSpQ4S8g6CASmXLCLfNOQUgk1
TCbe2Lld65WXgY4NL1fGXVJ9eN0AuFiFVGZZdginUPddZq9RyYx53avRJhry0XrHhxb/8TGtl8RW
+UfBdZ1pSV8Sn8iFsvvEqO2KPFRRj6Tj2fXKiUpfggM2+WSQe6h8XzMpAWEXtKOjBDPL6tHXb437
5B6hN4SX79Gs1iSFRlWDcMkbFovBfYHQu4ReOCFaS6XzYVVvRqDhtZERZpSW3jbrsBoh4I4AAptl
FRxmMwwS2XKuzpEZvCbduk1OzJjo1wwvXz6yFe43J5IF7FbUPrEgvrgJscKM1KinmdTDm78HXJoU
oC0m31fUist0Lyt/BiSZ5cCR85+ymOoOz1kxU5kRaRwkER9e2guSczWeoOaCnugmaTnU/b/2x2ya
o3BIFyFs67CyVn/MdJJe9V0ujS9IB3YmODLihYZzxW7IIkuQicUTVwdqRmMBizuqGLTf6/is4OP7
xTVH4xTnYSKYWP0bDQ5nGhqxuQ+jyE5ysgSJsgEQ7icvoaNYUby61Jctz28DRPkz0mouD9vQkzgE
8w4JczkkM52Ed3wO9WHNm0uIT/7kLAL4w5QEdalwsSM5nZ01bTBTJqPAWEPoLu32twR2yheuOeHi
VZdmBSr9cxZVsXNxLugCmykv0e2YNKY9Q/PWhIAq38miSDT8kIm+o395SNWUjB79MjE/r0iUvodk
mmWb0HS3F5NzBYf2r4Mi2gIWOpqpYNh5QbwFPvLZC+gAabTnDCcitbBlo7EVW2wIghWKRcZLhr+U
eTGE2ng6/MzCcCQRnJrmsjkQ4Wi7xeyxtBw7ArorsOKkF0zvH7ygXQ9pYXq7pxvbHUWP9ePSDXbc
4l6hWE3S6D43yESbDvKKxAr3ML2HwdoXM16zo3SmvpgyRDbvyaU9urz9TvHG3EON8EQdqjOUc6xk
BWzyxbsHnCMNxtVs1wBjhs7vuBHcRjlzGxl05Ye7V2VnjI8XAX3YXV6oVE4k8Y6bDW0nCWC617pb
JDiaSMve3Md98wiHsNjLIz88XMPlwSEashs7ZcgpVHbNixRQDn7tH6LBv/IxclOO+CsGgOhIq572
Cs+j7b7Pp+glzO5BmzqhTMJhhqHj7CxMin6mPmnqHzLjdMJa3Wh3GRFfTUifsRspm5DHk7/drOrW
PzySw82bqU+cDVuJtCrg6ro04vPElgS2FA7+JXpmvknZqUjH1hPZ7nJsCZVVBhknbfa+E/WbrFs+
yHULMIr7rydJCEdctjAEyO1YnhOdwxBT/+gRqdKiLupWQ/9DeMX9B+twmTM5sdnl9uSxrLWieSu5
IE6IeTjL1kp0lkJdTnK8M2TkAqUzdfi0yNHpmmqXSCvRz5orBmf/MT3gNgRvZWeBvcIKj+DgOeS6
nzRLcM0CugBKcIRWZiuAgBq+neXFZ3sfG2pwpLfGqaj9q6mcOzhlRaWUk3A7Mx4wMCwtfoMMdJlk
S8Vfokyf3WygcGuOZRUiEid6fqfq1hAZfAhXMgcqApMAYuzIyTocbHilQbQ+OUm6AQK8BKEcFDCC
NXtHNaUF5MJrIlaJle/hLvJtWg5H2KlNRDflh0bb6qadIxyyrNqlv8O7Y2pl34S8c0HdPp2q59dN
6oRRcsTA3bmBawgA4ASq5rmvwD1MH1f8+MAf9Rf9netd7HTK8HX+bjF4/pT9lP5rsu53DHw/57bK
jQmrZj4FDNpCZdOQyUVgGk8j+nBZpxGtFV8VTSwtNOF3iMhjZYKH1b20+yMt2mGCo/2N2gJGwLYD
emVM6lCt78qvReDKqgyJ/cjYWXeFBY2blBRgWnDLQrx7lKeyG/cTRFIqKEzzzCbus7UvqfFYp+RO
HhV/XMHGP7ykj54Tge7HwIY+4ZPjUyTEN4oE9EiUVp4eqA9LgTAuRHD/o5eNdUHywQtTOGSxdEBo
DeoDfySHYyUScxaNhLkyCTtzDhcAsJRjUFsh9rv8DAu+kQCoHGVIdxk0mLyB7g13XssnYUT0glEd
h59y7SpSSJQD3x6UgucXN4gJ81DzS2vjs2THjcGR5pqcUvTHoylkEbv0pEdR88Z++xB6DL9SM4S+
PPbjRsOPUiJXovJpvryUZnJIJtcPOo8Hu6nLkEIPs0UY4/XnJ6t5Heps9SI397v9N5W4AwkfIEpe
VoSzx8usz8Ky55aWYp6o90Iwj2+3XeDlCa2TJWCLibx29XWPF4INnk4wrL97f+vZRAffg3M3WB8q
yRQxs+LEkE/R3yCW+ZNRd00zdxmAI7A5WeP2+XdtRTRGjxqb5bSbujeQ1dfHnVjoLFHmiTODLDdT
0cHzdRrxEghP5ZREMABrwLbUdLMzxB2wPvba7nvE+Va5WjKn34e5xFue4Iku0a7IShiKdwfvVFuu
oBJTc2LXEPvQeo/0XvLiOBdBzUkfwWhN+fzNJc88nvUOADCr/o7Cja5QuEag1eB7gF5t+v7YJmy8
fxm05f7WAuMGQdZhkR2hnNDqlIDadHqjNMu8ZhoOd+3vnf2VqWWQJ9ZUoDew72smh1VnFTsaoQYR
Kkl0sbm905o3v9iDKzThIJfQEOMsySYzvd9xaXhODGzVs55TYdAItpgvesKMEddXUSbCwDQO23B6
yD+QJcrr3GhpLwWCgU6WN7g+oT9SNNCFkWdEC8nNSwFSd3J2YBitkMDyOTbbZvjo3piGW2Po6mrd
p+Gw9kGwbU9QsxOfM84Pbxm0FRVKR7XMp20GmCc8pP9xY+keTUa9MKcqMwtDr588o7acKlku1Yu7
nD/PdgUE2HlrkEz8Lv/KMuKtmSKNUFITm6WMze9dozrVspmyaoeLOO8VwoRVtsuNGhude9W3hvBt
HFgtTrI2uIXYUxZMXH4IEXKBpdsI12yWKw2PhAXKRnI3PS3ooYISReMghkdOQsL9QrAFExm5liDo
37cdIfC6QEMTrSqvY+JSr9G0koa8rqXY7bcFIUg2AdR3JqEhh4f4ojxySgzgwBVjc6qCYwDQiZt1
xXkAhgQtDz+n7olFEwOMFJkSAHG9vhmPJdEMxq56uNbStH3HNKlw1/o3tqbPFfVEququH5bFEEwI
AzFRKZbZRyi5cZsRqMgnkz/4n1jQ8f9U0KQbQbkM7cXe2nAMjDnGtzWIiu9txAeL33KFcoGdV4+s
tS81AT076gUfLtNvXX9CYhYoOWQcXm8MolOR+lewkz5OPSHSLzT36gaDJtv2cCA5H3dXw+Y0h3CO
pyXwsf9TuINg6ySF6+z6AofG1KlnQlpRu/R3VQ+oYUIFw4D1b+vU3Dv0oFQhfmxZ/Qc5zTPZpQyE
68CLc6ntCkfGEDIL+r6N0IhDcnNAPLh+EIiwldmmgn+J8GLpNRsJwQb+K/X0MzuTJ8IaE/z/6Ytu
EUflA6pJjNr3FoZsEYGxpGLUshkcEbL2R39fES7wdW2Uvv3H9430CMUDmx/CBLiMtNq2i4vdUyEZ
1rsWifQJi/KYLyBPI3MNRvReklAq+Orm3OnABYXHe56WMnEnR1ZN/kA4Ah15a1Qmf4fVA9b7JGwS
1eTYOol3pKphFDT/krJmT8PTBt+nCH3HRxVJ2KQA0XBiCzaS1PgHc9Pzcc39YKpIiP5hP74F4I6h
LUm1WM3Z04tKxDb7ffXAwu60C6TGPrDvKye32UZA4W88ikcDjdaNWuhGngepc6fbUwNXV7klMDuV
sX3koDTKsi60WnF1crGOocutbapThdgG9tphwIMUCuq7asqSYWt6R8RlNMsv5gBT/+OFwxrdw0r+
TvQXinPMUJ1V/V+dqg10jgKsjJGjMdVfY7fdhWMds/xL7VIysZqQL/ZhE27J38tx2lf2coY9cHlu
Rkb7VfsdTiQ7YNOBUlvXNR8ycGRrupXxztieovOawNYyjb+5FYMrMxlBQtrsui75TL0cpNKuXZlJ
zuXOUKPMvDtM4FxW3wUXDktJ1gGUw8gWIxmJ842RXvNfqCKhIWRcvnH8XkQlmCtwRwCTi8plJu1Y
y/LcCHPyp/iKbWYq5kjKG22RZdPjsyHvdbtIrxQCQjUQpN+603xpg/8901C/Cr8nibuyGIVw1nwr
hvi8cCmdTVAs9W4mpTroy7l1nNkHXmY5Uo3o0zqKvI1Bq/uPATii8+bazizCKHy4PkoE7Uc+ww8v
kgNn87WX3u1/IJrYhxVVbKTHStBH4w0tmHcmIUFXymdnqqpBfgJNO/0uQIF2AMKedgVseWTqa7uS
3k6AcgdcDA2M4BFWc/N1snEHzvRi9T3mi/VOgaCUgVl58zsJ54EgXlvDLlfUhQ1GYKTUAUv27SFQ
zzlM8uXeS4uuUdO+ywAQ3AD5hcEk0XsCFShdRM8UB4+OyZxOZeRr3wtLc2vdLzUKR9T/cj3tD12+
0HHooNJNcwvgdjkWpro6+ikCpBWvjpMvl1GNVW8DT930Ot+H6fkGu+Z+1nla9Gz/A6j8fa+9wzny
DRcAbWDQnJwdUlfNt1yHxxK71QtKT2UKYvpcVeRKMHAK9OzhgT7rI8xVE5eo8darD5Aph26x2p30
iDKdW/HxxaUmUjfbc1O0WjXn6BsSBbo52s9TTmNcrasYkR2Eq7QfCzQZx7OI1B6Y9Bne4geIDZU2
Fkh6EP9hQnYwNAq6SrUOFgovDvEeMOR0UeuEyuSuLN+UNQPhVdb2X+6YSa7l9qbclSyKnpmdLl1u
IzZzeumQiqQzNL1V/HpaCGmzrVWKcIyTu6KOtpBtxn6zfhaDGjtbeIpY19xOUwM+sMRj54RSJSLi
NphSn5i8safkO3Mm0258o2VKrY/geP47uDI6Xe9jVvzUajggVx5Vgcv6TVHO8wVyHB8iOwPV386y
/eEZXgQthwPtg9JSX3zqQA6x//SJ4ULckx6r+Kb9pb2mGjJrzL2SncJ2gE1GePpBAMu7fy9/LrR8
SfmpZwTW68A7r28n3DLQaCoEu+89rMCsuSvo7lXGT2FKOfAjsyqNH+tMUGhaJkrl21UNohCsCzs3
wXGPERN/zansX8hN8RruK5uBKBcopjJpOp1rcUJWLNVEoNN6OreB87aoZhmu6xMPyvg3r31/dQGm
fFNHg/RBuo1vJnPOUJOuZlWfzXBtLTBIkOjelnB7lPkzZiWW8hV+pdB2/72TdY/B/uFpwXDEOXy1
YvZWfRoekSzz65Vy/cD2y8Uf/fYdGZf30CQ3POwecgeh4WOS32OyNrQ0ciChKWHnpsv8SARdqiC+
sOJjVuLP3e6wXzYBtJ1pEEiGASXZmjm9HdYVJR67LrJLiSfl3TKVJeFVwhN6y/R3d7AbWTQ0U9gZ
qAc0i3Y3/k+Wn1pKAdvKu/19QyRcKuo9ZcXWuPq8inY/TH7MG3AbG4hHU7bcRzkEbUJxYPvzGBET
CRj1tqTOr4r7kMOVMxrbjOE56Pd3VrtPGKYR0S/c08XsYGrgN0bgNHTj4gmL4zlc0Esx6Kq1f4lL
j31LIsEfNXG3AVQ3E/I+3opJGiJdkBHnaPtYLk6wOv1eeh7NuNRewvZbNzjlpLcu+rAJOumBzm+I
sRzf+O4wGpEM+gTB81Encfh0eDhg4qoZr4/PiHnHP077VaA4tirv1LlyCKlu02N7jhBC7T/lkQiu
2J5RUgAM/uxF37OH3YX0PnkHy6ZNmUcSfSqq50VTTE5Uctjsgn9409+P1d5xigte1yPMzqjLWJ1E
99eB8EkeJhK/dNWyblm3noZ+pwk40g2REjQnQ3YvG1ZfDOUjgZn6LbwGAnX/mElMlZaJcpUILOKi
1RxhW1TcKnlrwq6Uae5ePmahB+bRFQc8/m5TExMbBE4AdO40Vq3tw+tI9AZCGsqWNTJgCWX8Paxt
oPHsVq9y/oSLjB83u/jslwkBHe7q2rSk1gHZTawUAzQsb31rvgjwEnbjWSeDWsDHp5/18Sa7PE1d
ve50lm9aVk9/iAyur2DVI+Kwwd0Bjd1GSWFKB7nUrhS9MVycD15B9BRZxkMPAIaPnDQmtP42szHL
QRPVUDJ7au/GfOaZdejO+NfjSe1NSCEWaHNtPOFbViMNBuoGfjAnSVEn+joo0dLOYjqOceFk8mQ4
znIpU+gkukNfgdhVN+e+vrqMd3+t/Gw2E+nmezl81hdNgVWAOIyISn3CexUlwuGDsChzftVZFU/I
uJLUEIsHhuq6KNpFBAmH2PahGvHptpczoFEQnSSAqh4j39geM774ztqr5tYQubMbI9TMQX0AQ6UU
RXLWBEdWheIkzvNJdtBlIVPdSKqAyrNSFDMxqm1pFkqXbaoW604CmBrQmbtzwQxWwovmYsybyfcM
JpI8N92egyVBdgl4CHKHd5N0XkAxopRisPXfWLAHY9oppk4pkHeho0E0RmwSVDpwy9Uz6IG/phWq
hIqQn7O96vtTO6G0vAvX53Dm9kY9ToAyySA7ZuDrWmI3XJyy6oOLpQoaf+TC41ZH6kWMXuxRlxnl
7eHJo/kGQiPeobZyIyzHVUTkIMmcyy4lAtRcA25UC1D11/qvNYLQO1DKff+pcTc8Zn/zA+ais5Uw
6wHaeF1RsyvVr6PYYlwGE/ZakeSzJRneTuoWEXq2BCFHutQPIg1KqS8n1CVuHvpT9padeiWU/6vY
z2SlIZjU3PBatpG1NF95PUOpVwvD0mVQ00+3WgpTqe1qnBNYsqfycdVaDhMPp478UUCFEPpFUzdP
ysrNYTI3gW3VJINbCmi2NPWlKD6wkrsdodjlICWCfsbdl546iUsVQnGVkMr9TCszOCwLRDv+7UFh
SPoAn31LJZuAB7Tg80btM8aEouvVQlIpdwZMEiQ0CGQF+RLIhwN7Hg0N7wE2x+N5UT6q9u4UdzNp
UO0Q6cDTFSyY8fmu0bUu/LyhWqzHdoicxuhcvhtijuLFSGMb2gvZsKyFrxPy6ZuwXGUDg8NYrFvZ
78G0mxUzhXC1tujWBfyVVGqscn8EfWs2XItlSkXjTttAYyhA4k3JD4FhQrzIsl1GZixde95aOnNr
wPEkICiP3Xz0uAiNsZXpxUIsY5ob64oE7fGW8FwDn5t7W+ji1+vJK5DGMmMWY2ZrTAGv8cSCwmX3
1lUTQuBftPYDynBURCJIQ91Tsj8KWiwIYraIC2nRjhgivv/0uHBOGpv6u9a3jXfbuRoSQ4OMKq5k
8NjGpL2ByBcfC+oYHtzYPEdRJCl4EFx3cECr5mVoquQV9X/xDZvN8k/l+G6d/UI2gGwjx4jFPWsA
MAae2nWilDT1eBS+kwI2t0RkNDk0X64N1Mhw0D1+LC73adRYGlkwVA38b9tdAditV0H7ibMCAuJ0
CN+r/sEIyTZouhDwgung1Y0PilnGNtPv/JTwOYSXCBhTo2uUyQ34ZmGBDDkU8sYd6EWPgWDun3zV
CG1CSiphCnPLSfejs9zagF/WsXm05HRUn71/duhySfJRLzzauxfo0v+oVwNrvF5SL0snAIdfax9G
B+aBKnZB8QP8szv3vlP9xNSoEuzVhKsMXTR5rU1agOQ9Y+iiPVBY5J/U5/zuPxrnIjKxmp0lI6qe
VSlz1WLY3UL/TuwZ2lLYtg5+tk2Md/GGM+mjkxvL5tAJfG7i+ElZWGP+uiKfE84oq76kWuh23+rW
l0ioEXhqxOqADYO9pKzNqV+9aANAuYc5BfoRWx2zav6BU35VPPN2cGimChH97v5cQ4VUu0fPtSPj
aoOziBcdCrmZomRfSNuxpbYk2PJ0DJq/gY3HsuTDVJp2gOhnL0XOJVr6Ah25DxitQ9QjLBYXp2hO
/uEeZZz6Mr2C02yKYcqLCLEhAVCd12DBrF4aIwctk5/RK9LPIoxAG+5+rmbMGhGkiw8clliNPOjt
A02f4ihImWf5A0dFsVAsWkVcuXJcveb0lqjVfEMBiN8ojrghjdjpYrEraWbdSrcCvNNHzT9So+Tl
klivAFtFJKQCKqb3DlPOuyx6G3CeDyBgkGRQFENGaI99ypmODK0xlOaaMujMjmepPZ0vRG4Vtm58
OIY+k7lV3JiHBvYMaSuswZWqWzPQQvap/gu52egVOJIk3ZjpVBZ9JamjOKvVZPQSUMn+tLlfD/Xu
ksBXssOqmWyKZ83ba2OiGGRbaMRA0xPpJ24vY40VFlhaeEINGugV8iYCwGEQZU7xPvSQXvJ7XfNB
slc29Z591bqqtPcWNN/po9cCIKGeiOlx1qqFEuFcCBYdZws9pg6cHZRo1/87xMHNhGu8s1WtVlkD
E20SC8I1c1JrTpu79uPV0j3aIG0/P/Qf8Y7unZuycRkY/k0PNCOPDUQagrK4cKsy/6DvuxqZl9Ii
CgvSCdAcYAOuuubgcLxUBMmH1AnPqyvvOuFvki0yV9PqDjb0da7ZTFe2VwbxPn/F42BbjfkAjoHC
aRmA/aY1LKghALNsHo3RW08ipJFVpJ9XBuC8XfWGryWV/hAI7LuqJ0RnZjpthjs0H1Vmw5yIMMx0
ifZf7HJk4LbRXgyVSuZGgd3k6M4uVeecOAGubhM93oukT3OUyq+WxFWU2bI69qALJ3Ejul10vnsB
Ek7NR9pUvwPbZcls1vJptQRxtAomps07ZsVER7gr7wK13uDJiVtwCEJW0MOO6hXuMykQCfysF0Sb
oZfwWRhdJy5riiEXiv1LVyS6gJ+9MD35Eh7thfMgkOiOG7RMKVvjrngKKnh10J1aWzPZ1TAUDfo+
MtDrzM6zc15R8uEF1vJfbbNrIhS2BRqg5Gs+ZOIhDRNY4DiaUCoMaf8D954rbcZgB3R1wwMyM22S
UE6rSYYj0t0BL1rnN2dlvAZ33C47AcBhg+WCOtg5bLtm0FNt3FK9FSJc0TXJ5KGGR8HoDDKOj/bG
S5wXZc2qcEu+nhaNEe8PkQJYWeLItxW4/ziVLuX8maYs1sTQp3XH2ezew+0uumC2Ocwlhj9/IJYB
vLV6arTh5ImF4jQjcsDdWV3SXnVWJ8DyDEFRdlgakDk7tNhBkL6+lRY0yF5U1+DFy+GPUAuh+O0C
iyGfIGWhc4zxv2pH3abLRrkn8kTyrQK5VFJK2UkmNELnU7oA8vUL3/aMKSg2tTT3aUgk63UqOLfd
iiPyE2MdI/GFtQMozWg1RZd5sbhxC+AaTUqq7NS4civaaNJgxuMziH3ncaCVOMI9y/uw8jQlD8W6
DaU7JnKdm/ohL2u/TLR+9Xh5zEkiZ7leQuWHmUeySr0TDWuyeSZehZ+vjKAmY8BuPUrevMBfINh/
fa/XpFi1Xj1C2xLGEAzm9Ax5e2RzI0A0Kav8xZquOJaqtaUiB5fKNpZAm3hFSmiJEmDWKSrampYr
bZ1uxWp3fm7Dkn492e/oaGvfQFd+c6AajltNO0PXJTQ07zPO6Pg3BgNtqUYoyXmlwjJryuEydNhp
RP78gGo2gMiB4r6WCHAt2hYbUQZMe/kjm1zfUOfF9Xa5naWDs/4c9C6n6rgjzvUfCyF6y1tCI4c2
w/j//EZN9NCeN32tFT9fYI2VZk3Y9sqrdQOIC69JUjhupaD37c6UymYH4LsN4lfsEpt9CTzz3cWR
NRYAC30yO1+70x+XhyBqP3bjwuV68giXmy16D5qfzSxVCypawWhoOl8PO9Te7/95iDOroWMXSrfI
vG3n6lb5Prvqd6NEMzokXGZEsShCmhfab/NkkN898ulpYrTmy7Nml7wmWaao72aGc9DaN4/he1tx
QfpMjhXBUyrIbqbbreskrDUZdhS5tu7PkQ2vSpNzNy3xhJs0WEijduaTirfcmgqkOHOE4MAYqo4+
DTUkEAdI1Pp0wweuSl5LFuV4VDvNiFqYUVYgMRYL4BVchRmq856JDtlajTtyvAn9jQifvkiT65fS
4HAbiG5nPA9hX2LKgaMi/E3pzayo3hF3yG/k++9xMDrpXUrZr3UoNhGsK1kFLi9uBt/nEbdHyr4q
ty3CmlRovXaZDIxqt+fXJ10ZjQGGp+mvtVE+xzcqDYtu+Z840v0NJeoqtu0naj315RWRKUOPLH7a
m37IMB5bbfGeZbbD766DMtJh/RcOqo+tvP5Qi76F/V2a1KKDx+t6o6SiY/ZSxrfzuBL9W98kBGxI
rYzHEZd6Dse3jqJrIA+AHidOKuWikAiY9k2g/cePoh57t04HA4dX8/eJp2NMxj1E2+Jg1R2Yn/4A
1/xUeF47758tG9vrdZKslcNykCNs4oqgWF/s1R9tpxTChEJwiqulLnBmXv+8AAP6Eim83SVuQ7Pl
KeOJ2alOjPkqYIa+E52whSLNo8L//cQm41YnlPvPWJoCiFrO7lsZuIz8y/gQnl+/1kwKtyEYx+xr
2F/LzzrasZtzPcrydMJbOOvDlW0Z6Hd4j9Q4Di++iG+J4QYs5VlNOno9hUFII4Ws9YuPXC0qwKdY
v3Z8qBPYMD2R9Hr5h022/7LUTyVtP19zXIDH1VBYt/5nNPc7uHpqQbiH8w1hTpCEPX6hLSygAlNG
mEv35+lPt7NmGBYhtf8STLua4svCzcHf0ZsrDa6u3A5uotWdefkhzkG4ZjdBjvkCYoi4a/I37ooR
OiGA8RBVpkK9KOtbdYToJk0RS1OgYdWK3W6WKR0SD0viFsp8NzpUxD689oq9m6HxRP9RsEcUS4Y9
+FFQBFZwHaGHlOAXFp8vUXE45KX4K8sI0O+dyR21r91oUvUGz2BMQkYjxaAvoTPmrTPvtAH5Yb9Q
aLW9ayAWG9yxbGTX+Yh/LobtxmVzxQ6zmh1hISP8x6Mzo5xrb2W2AtLeVJILgS4zOSUyroQUDpiG
08SB4c/Z0aNkh/PNnhv0vsCIixRyDbxXn99asuKtGK6OilFT9R5JLxJVKPLv7e4HSpGlFM1yO3uc
43YTrw1ZFjf4ZCwIqvcByvdO5yHjlfRlWV5rLkPJLv+E4eSv6IgTfzRNBjLtuzUGGsdIgRbxJUMt
LwgcVhODg2h/xh71jmDJdS6wo+UGJfi3x7OXFwlik8owChIDTvHAgqlAWEttCay78gq3yCuB6dzR
MZUh27AxutEKfQceCG60ud1SQWQv4TX/5SiyDnH4quaHobvWBcLNvfIJ1qAjXI7IpoynxGNCA9YJ
D2tTFADfhdQSb1NdwgV9aBYBSlHfS9LgcoB0lXRBHqEOeBJR9uF3VmEPhk0N+3ixvv+uQSgpH691
yvbInGfxUvKytmoKqATf45EVQyleVLjgKIrDXGGRdvCct0ADJ544GxcBgLEVTjokvRYEWZr9W9Hp
jeLh0dMRdaO7LUR8aXc9XPtGMsE/bslP7TY2Xl95Bq8FxdAhwzkIl4+Iyrc1BAgw2jVZWMibDOrb
nl8EgIZ3GoukbOFE0rRE5VV7ckozm2WE3wTA7pPY2ZV6iCwOqCBjQA2IygVD4MPAvxu9XXvH54Tu
2clh1o79GkTe3qfpriQhxO1vBivnhcedBFw+HOuwuMZYx0FSY4KmcWCSxFjvVZup9M1Z3gVp+AHd
5171sujY/lW4xSDmYMuYK2mSg3Txi9Xlc/xRjKfh0XJvlFbCBw+En9FeXV7Oiz4YcjF3LNO7SKcI
hQPiii8sAHU9gBTba5vwxsj5f25OA2CJGC6dmL9QtbykLRiQUCnV/F3veIlJ9U4KLjDcX85+uQec
ma77pZTUsP/covY7qCfAs27y/xyHC2yQxqcGEocLQNOJwJmTt8jTOQXGWqWIXJayN85P86X0uufq
KX3eyFLxMzdYesYPmQVSDa/uUwRNBJdskc+DYrGy2rS3xwjnaz7Op+IsZpFujSA5AcH/tqngY/lt
DmADJD8W79gYGM6XfslJRt6Z/kZsk6zhBzsP+b8IL6JzceCyj0ALknLcubpIOAwlF3b2pHPBrDSb
iOY/iF4Du6g8h+WE89uBfvGpZE69Q1U5fhpz1h+vDxWymEAUBLD8jzNM7zRAVE9MpWuLgXe5Uc1s
+N53fuYj3t4N2b3ZixuC29vPIVipck6V16zxpOnGRrFrJEUT9K8tJIOHFAJeth3alGo6RkNSis9J
VoIvoq7qvm1K9XPmLLQSgKohBQrZIghDUZltq+Ie/PtLFQ5KxkWuAm8WoLROnNx5wzCPGiW4Gsdk
HOWTo+AYm5rrXWNiTeX5sed1TZ8cqCSvgpHpXitCFKubhrunMFaoIltPPMYp6X7SehutprjoaFYO
AbdgtXy2jdx/naDhNPHBw2EDEcEutu3V0U64mU0KCJr3r/zaOTjc5akw3hHhQYrMmzwIUBgWs+Hz
X7Dr6Ehdx+JQLjC9wvaz12E3E3B899b0Vmu3exVaRobajfLX+4TPMk+Fee1aPdtTfCo8xL+Gg2nv
oy3xDymeS6FXKDN+MWyn5b0tYZKot7ctr4GKCWsXOgiScJA3HOJOG+gfes55ruFit9hqcvJe36ac
wrfHzx1hIXk9ODGxwWsr70KjV+iqwhQ6KLlHbmUPAhkvIsOYeJnumBGhIiEDLnwVs9GKraBtWOnA
FHOS4ofu5Sg8q9K+VQ8SxSHOD/wRB9sHYMbQUmRK4HadVVp2vF5SzSmSrxYtzU3LhHRPPnj+jzJZ
mnmEvuVDXf0fsSRRaJBKRevtlmkNOQinmljzEoPZfnrjy2mYbl11Ov9BG0eXpDSYBIgk6A0DhrWl
uKhDX81/veJIGJ+nW1n9TVlUdS6zO4PDC1RUIo7M+52QHsF0pf2cdZFvKtYuc83aLDK6OIdPqb6V
fhNk2Q60Pn4trLCBPrQ7psgrLf3dfI7MNv3GQtQlgEPU8HKRrgoD3YPY4NW2PWpmoJxpbJPga6UH
OEv52nRVWaKxLrSA8ZsIKErxxAO5d75LOterYvR8U8xLQST1SBoRkzoea4LqoBnHKWKdJBWAIn8J
vnJaa/d8+OvgnrFHDyXPCYGkeYJpIIHInqhePcBbbDAuwMZcMmFRTT8EnTrpjCnSoB5nZKgdqPes
j+jNqERg/Ek7v1IZlKgMmv+uPD9Miq9fFF5dDyEf6Q/3hw4L+6MaBZnotHfgdts0ed2xA4tD1NY3
Na0DbR4b+khpygziA5dM60kHfvBm1GIhyNq8adqOWEpwm3FDnl3Db0mM8qh7i3f+FWLadlaGOaI0
+M8Es97wNTytZUG45IKGJ6B/CH2jcFK1HX8pXdlHiNceg5SBWFXpRjsTcaqLrO2cZMVUnS0EeD+a
zeL2PDEN6e3dutylusCyNVf8W6vTONrAIZAl8Xl2r2+vsx/LHVDHmxi1OeBvdE8dbRG0QPh4H4yL
fnUQa0qP+2tQFTYqNxzdfo0qlHssl6k7z7qPnatQEqb4U7SK5Rtkw5Y0asbsVLbvoJe2xHx7rgFp
3Bp2bwLeY1fYKMbpQdVGJissqcCUIzLAJW2f++E8LQ1LCbaDdqPw58Zaf6Vav7F8ZoOzeGruIV+U
RO0FRCaGXUtexm5aUyfl5i4bZEV7F/JMTHZJm3jRTuXGsD6bwi4JjgFCYJ6aJfwP54+B/ii5VxoH
Xzanoh6pX3MVKVcUsOMAOnFm2da6S1TLQEQkKTW75sAKM32VUn0t9t7FlmS/1Lz0/3daLjTWhGLv
dGc+co6Zx1IEQG43Nuw7cx6Jo57d0W2aJY9WTiAQAhl18tf57kLl9AZP32Fke+8CiZLPTIZ1WNpV
lvboVQHSZ+9pdDIPejy17sZY+y5q7oFegpSnvx56Z6qE+NG2ZheCrckykaPfYUc54z694vqNE1eH
HvmCBwQ5MrGB7cwbpmiwKfKg5VPZY4IhOS3Tof7Fhd5+eBJwAfKCcZhTTcEpIA6YUv8Iyy4rZeOQ
IQog4GRvbU7tIi/+A/A+pl3PafbH1nG2j/fwVONglGKlNLh0+9EVdiyoYpLTET9R+zsAK5g0MLbL
8lTkW6eWAY/+1XbuCVX93y9gG5w1g8u+WwHBcr2gX1Ce/huvFjQWHOQgXVnWLpNdzkIkgLZk+exG
omRDySVP72Q/Peklruxdhu0P3OKamfq7fOu9ovpGnXTeZAGVZjwuHCf5gy6PO0Zb0nI4JnugBuwo
CLTI5uoMMoWW/F0IrQbJCj1lGrkXCdTlPcWHSUQ5uTCVX32Y1+buv3wmRR91RBonivXR+EqQDslU
DqHA9nCcWPwu+pEbm4GkDGKn2gJlFDlSSqO2/Ck2lSgHfjAYVuEWBeSqBiXFXyD3tifl/2vT4YOH
CaBiank5V3wZrDbDuWBsK2E+B0flbQTMcCJCeSAhr7F8sgrE9FerAA9byp7/3Dv18ZgyzYOXtyXC
kjzbOV09fAU4sAyclQRXnXfbDzCr8D+U3V1KFCqMN/O9PwGOmZO9IVEA6Z2RZQazHWwFVqWV27be
eplM5PY8ncHvgQyzi6Bl4nPu7tcY5HsnnTQVQkv+O9/DgYc0sKftXBS9doONx/2hzdT6THxRr6Uw
9fcsbchHbH+c6f/+FghmhpUD5LbgG2rF0GGWVDf2fhc1yHSV8M4fSCXZw5ku81/cNVXG/VeeqLjx
mtbXZ1FI4iNN5uK3SsO6MGL+9dNgGhHP9AzQf3NwMCLoroYDbIUX4b9nzjnSMvYuV+JAaZm+8SXL
l7ddu+ppEDBA/Ds/EZ9N0WEOC6qmJGpfVkZRRFWnJjTdgtU4t5m22GCe5u2CjKgdBcL6fTRr8ZUD
CYkmARZK4p446RbIbOCAB5CRqvdIWoBwJHt7YNe1KLkmgpA4dP0qnPM9+zNf2YLOwhiq6ZIdvug4
yiUAAZjEor8Y1dFv3oQUzxsPhyBzB7zLLO0BiFF9/vwC9XWivjjb4iy/j0SeO1hZWf6VsWouq0+4
f9JWfMFOflSILQ8ToLn6NPzgzgr15SDi4N76RhVfOfWJ6gIxlG1mczHF5fKX6rAdajpOz7ZNnqzY
3tCv738e/h1zKrt7fJPv+ZUPSiJ8AGzLimCT+pG5jRs2of1K8FoYjD+FjDqSXqp/uEdTPlaRdfx/
T92H6ZPG5QhvRgkMlwEmuV/4TMWnU1hfsdfJu78eQXgj7FFkBZOm1KY7zCDtnbIXYY00kY4HHBdR
7eaGGYhyVuQfxOfDYCI5kgJUYf0uSF846IHLFdnfc+jxLcndJ/iMA0JIHh7Qg06OJ2As3mOTa5s2
JwfVP8vZ5jNjqCqiaIYvfGalUdMWiqrMSAuw7ckKrKqvLjV0WydEssf+7vz3R50STpi7L/nwf3bI
O/oACBDXdGJUsOMlqAmlrBf3ImvMNDE41m70toksA4GjAuqnsvJl9E0plcxLkcu2SQ+fXL0bXoSs
Mdg4n/jnbo7+BWWvWDE1kWIwu11Hp97e/1fdj/Z3tGpW9DL5FWHnJtvI9i4tjdw+nbPr2fp7rnYf
ENuGvfibxYX6BeUNEbhhIk1ZMe6gi5XIyJwgilE4xMl9/myEBI4R1XUZN86lkiNiOP9LwN+Bb2yV
96GYnAP1SsedcrEzneq3jnMYprqS4mgpfNn+gxHmyhzFahAksRJYR7u2zFLyar1CCPZxvxNhGCAF
/JQZZCbTruk33XDjgI7RwfWLm9X9o7HfoOTFIClE588u5I+DjXXbtFVURiqrlyLCkutZ89N65ejQ
FS4P+krtJK7DoOJD/FKtWD1XyZwwVjLI52TeqJQQhb6eMfFfe3eDv58q5jfhipcBp79uEWQQW2RP
wp/vI+wDXJgfyL3UcaJFq8lOnfEKGXBLPnHoKtAaIJf+LT2PaBm4ffNT4WGEmZsi96Nx9UXARGUL
nEFPyPgJUDsyEK8FFG1LuuqR8pGoFGz0GZhD1iYahCR/uNHaGe9KsgHpSS2/vLRmqHHoVgVXN08N
J5y21A2X3ZvFghYsS22tFWEs5NhHrUzKddOxKnwyYO1LNp9ON9WQNK/JvSCqurgigIPN22FNMqw2
Ohopuh9cHHsWg87lrb474dNdcPOMmEfXAEETBQB00lzsJCB0dblD7RKijk/7C434037Hj+0grNiH
HsVkf+FAH1Q6kYY6eDM8fmroNMHNB24i6fKuAppDMiCjsdCkd8OPLUSeRXKPX3ZX8DhguA32O6w4
RfD0SzfdAffZGJCu1WqUmX+hA1NLlQdhithAQ8PorJ1WgSkkF/vrGcM5hkGnQP2FhvRf/tTVFIor
TZ7yJ/QJ46W0ZcI8rZrfAZADGZXaqgjXTufASY6b5k01G9UgojQ0cMB8dclSANtawoPF7vILuEYp
e/Gm6osb9/zf+JzK4/Puhha/2Q1/UdupIKVPwtN+JQ4qWty/NBBYkVbrzYm5/7iyZBYiL/UurPjj
J1O/dMbZ8EP4HbjJ/GRc3v5qFSu09WiexguzEOtwDq/JN6NDMTphHbzVv7IpUKoS4ckCPTtJxOxS
QP3dOmMdxQ8ZZaM6liPZRSU2deUbfBlUmYNwzy12T8ArEMzS8zD7RAYJRvFPRcraLr7qKAz2OYOq
e6L8deNgyVZjEmlFkJGGRl25IVkZ/2c0AVXQkzEOIAHFRFi+UF7UTD/rFIOyAXpVUY4EH8XF4v4T
67n6BBis9q7EI2PmI2VSDQU5UR/HBpAtdq9+mSblS5kq227HI3w+G9Uk7YfRkjeC9Kpn65N1b8lg
GkfGVapSuy8H/uVdBy8R0W1gmVzGw9rnyk8JPVzu8uk76e+L6wrhvnnKj9gBFkx/wtPn2yLgXzP4
dAn+2KJ1NCVBjTnXfoZseYOvkmqZiGjkATPoeVIzKZTV4cMjugcUvBAU6IXEgB9VPdlTHL40+Aoi
QgDGVn0ctSvcTovsZ4K7dbk8OFnhxNNnSS84URvf3mwEK9Nl4OFVSlGi4RJ3p3ZjzIjvvfHVSRxc
k4tUy5aJQ/F4lm35dEmVY8X5VtTqSmoUSe1qn7wvZ5ZEPaovJKYrRFvN/1ySWIGN4HpIfWyG3idJ
Uq4uHZIHL8D5mvZ0B73x9JIzIZFWB1w7Nt68SMzKKk8IfQkQhX8/4RT/kZEZ/Bj4Rvm40sh5wDKz
b4Fe8WCFtieuwPAfXQ+UllMBS07u7jkDkZ9N+7zhjyq8jKkvW+CIY3NUH7TbQ3FD9/z1nlLibnUH
65E+tIQa45c2PAlyGBfSUgievHhiP5AUA2yQIv+BBxi+30Cic+dh870ximM+mXWteRyg2e41D6xI
MiSOm96Nx9vgkbyt0JXQLt7mryM0DjzhMuUM1C94Mx8U9XOuRvLv1yc89JUE/OKkT8TRfkCFlqgL
2vmrMpb5v1lDEgONDfd5IjZMaedMS5gFBv5jq28BspizA5uxgFkIm18pq2V79PKuEsrO9x7uCgd1
ptbshZgEnPjH05oqC1xL/qC5NoJb2Ub+KwBPYZFUL0lMQYWLsj2vROr3/dzzTlnSXMW6VMafnVQT
rQWMhvfPII05ixewTGAgo8mXdL/hKnyHBGJypoouswsgCsgsYhxMvjdG1oF70uBBB6jo6midfJNd
pXF5BCz37P5HPdkA0M7hThLsWzuf7uz6a5XFPdZwvizFB8YmwbvyMP51b8Ci5PeKxP0tZX0iObbB
8U+oJfyX+3lCOIq07BU0kGKVOcKxYFz0Di2/6Bq9MzDYOgdX6D4jTBythhVQD18iO5281Lk9n8Oq
xbpNIj4M5AzCw/XnGZFbrwdgnn22Hokv5c0DQRzH3sNS84i1nd5kvrfxc1erFWIBt7vHd1kEz/lM
wuo/rC/vFRxqFZ5QVKMedTbaXK2JD73FjEU6L0HNZItXpbc2+fIJUV49pRY71ioWfT5KaA6nkwvM
uEZP3Xxc62ukRk8QFoZKjme4odLwHlPA0IG63eb/2lat5W1j2JDsh0lqdqF0WoTZO/xtDMCXZW/2
3XOFUJmDIU17OluODe7UC1EDmbnCG0cFfjj7+QAzk4NBK09KkEW8uPScn3u1iAnWxQgYjzJr+IK1
ZNYFChxWUu6qlHGrTduadILi8Y/IFY1tFMK7SgYaMf53DnJXRkBZhDwzZKZm4+gaBKpMUZ2Zz89V
FaJ8U/K/kHk5vpFRiwmdDdJdoUDem3+n319T0sSl7dwylejP0VSisn73niJc/PikAvEXpKlIcxEx
CrsvRWvYW+tWw6W0U9A5qYA+zLhGcrzyT5LWCqDLu+ILDefsNHYWwfa0gZf0BZoDEXH6n9LkRngd
RxdDSlP69avR3ycfoxFwf37qZlLoxpU4k0pkWVEp5L67gVhyWFa1JmnThFnbhos9Sr071PEEiEwZ
ib1iqwFW6xUI93Dns5Z4BlBqz3Nuy+8+ikhEuFvS0RAQ3Y92KHKz4UTsMVID/yG5m+qfd5tgiwV9
jl/NCgBFttWBXpMIcVEbSDnwff8jnntvSzK3Iqtw+en5lyoD1DOSrvC2TzvGCmFfaZP3DoKjY740
X5xr8plMHSJYvG8PXmOZEk5DMHxqOPXlg2kCacX8RPJduEwvbRSOMIqkc8DlDqGrdW+4aKykUrt7
gYQ+uqDEhrdk/kozPUw+J3pt4j5d1snPzTubvSyKXGFjV7pj1zr+psFiyepWDU4+ladXAdPtbySI
s8Pgz+kUUlHIMQB7nxN7meLOyR0Q8fobNeeypgBS67MRCn1Zp/XZfRyyuN3G3cfQfzAm5tPZWojA
3sE+baRQQWv4fxrHNxshbiQAJ2jNFZanekYgS3LH+JmAUOYmSw6TEATM8DiI7nAOBalCVtIWWkGD
x+jQuKAHays2rOguRIZlysajdlj8YJBYQfaeKudhMOvuJii6hOqZ9eBqEl9xSB1luktKuQcKmF2M
60L2utnrJctKtoWYf0iu0VoXDC+dVNc+OS1pJc+x1ueSzeNru+0TnT6plIh+cSM8Z8UpLS2xjuHR
soH96pDzTAVOfoheBZkAM88x31Eq6Bec7vXyK0ut9DYa+vm6qbfACuCl26bbsw6i+AvDeUVO6A0q
EmQtIuUDJLR3egjSblU05ULUxAG4bKoK3VP9TtAHckqyc1M1l4VQRIWQeGeVuafI4KXGWmvFRQkZ
3a3kr1wGoM6PCv2+AJoo8DSd+7si49VduZByXfr0ZgbryzrQu31mwHNtBT70+GXoMYiUCV1hQTRr
E9xtEeMkYDefBC2MOnxt7Sx2btCjDjcjYJoMoyQzunwAm0LrRnt/eB45QI0fLcZ9x3ZBTNbfgy1z
s6blQ2mgFCJKMRUgTqEPzlyiVk4qyoxHKj0xAU27XTVx5iXJVYFE/vw81/Q/K99Ekx+6tNlKI6RU
h/tNXvguF6wDrQY6Lqlms/KvkwIk+3dk4sFqYrWyDxaCD/vYfoJVkc3d8xBhcDM6zHI7ZhQSBKY5
xlDzPAyL0sAnYWvAonIxhtJ4mHQdcgVCVHYerLtJ2wn8gMXaINvSMF+aMt93kbvUtmV6QZGArsua
q05bqK3+HaQlL+MmONAWyTLeG+I6hthJyiehUfuRf5c3z430+pxkdkDYsxCHsrYwIhOMhzEZn3LA
V6JBL6ZZ5nU+nktyx/4hiKn4NbqQmInG/5gQqwcKEossxEwG63zLz1bCSMRgvfpTmwdUCthI/UGC
LunVP14M6NmxgLJRB36Cdjlz54m0yn61iNHqY8jtPk+NM/MOBVsi42lpNg9pieCB4iyWTBJixKKY
KaCegBHW2dDB+JxuWBTE99A/iK0wnX+8Zht12HhDF2hQeVCZ9r8xJ0C2VBPT+SDGMkDLwMAxDyiA
nzi+eaVq7QzrnL2qX9rYadAarIPCTMbiH2/V/vY06IrBSq/TrbhgRBHm7b/XREl50CbylOsbP8KQ
VNx0KAbzLXz+v31kTqVNBHyGQGxdnjBXjPP13A0RmVH2A0B0pS/+8HovFkDqZrK9Qyzp0BTWf3BD
xPA8f/E9MGThJkXcuF66jOHEafVyVnDEMpjutpGcF2Eh1g+SFhFi1LDVn4zErr4W6cjF8WGdxwiv
Tt8TDTupwx7YsBL00JR0iOnM/mCF1fkSt6NicM+I17z7vRVxlu33E1WGBQgh3/k3KeIGd3NeOb2I
W3YWaBGEWLiocYC85MnKp/QNQA/OJuhbVjOVwvwBszrpKrcsPKIDKHEIP00rOjdnTDCBJxqh/mbR
tkdlLCBn5yWYFcKt1LXJTYa6BVxK4fAlUh4Mq1RWPWqray82Wbx3q0/oCktDEsR1/DTwFE3At8gm
wY25hLIa57nB1nUxyN5dSQGcyc6l2PYTX9wdAb9mxUseeX3SeLTtxItrLoWXydCAgv2Z3vvn7SBa
uaCXJYzOoI3rwuA9CeSw50gO3qpQ4Buz5vhgpQgKAtwhNdEVCDTZcUiVWowrHJqLeZy6ZyDiDP0D
+ruf4io67Neu2hQbcJO7I6if3i77SBOR+L7C2209atsFxEb/2l14p3y69fUydXj8Uzs7Jq6HWwtk
SwFOSZvRic2BRx5vceGMl/cYopdNwwq5zZcG8oggh1zD4ApaUQfIS7R+Idw+2i25tChgbBKR/kPI
Jckf4oC/iCe9ERuI+jV9NFFmPRI1zbrFKp9ZGSlGsOHtgnhOcA1Pr0ld/2FrdVmKDnHpR05qn/BI
hpvG5k/3lYtBkI8qdpONDy09zbrfCwXCMhSP3MpCO7MRYYykf04xv53GdZDhpQdLPW1pH2BQ73Ql
p34eqATicpf+JoQTzKQlWWrICUjfHuvVGYojCvccKtiAdkYOn/MR5kNbu95uAJQ9TboqaZomiDFd
9FTu968S4sKnndwY+OIcDC78Ghadgorb3fONZCVJXb1dbsqLKS245YYwQYNRTKYS1I4mJ+FQ8OHy
NN2JhnVqxtqlLhW3kXlTni1SIYt1jK7ki3MvSmV1pOAHFmu/bMtUZ0cLZnx/lcf/xvjHr8/6YU3+
7YrXCPGNjK71KVU07XxOAU475jO/mD0NqMUr3NK+db+CXNkaaGwJo47jKnWse4gaCu3SU9B+oqFA
6yLN6TpjNklAVTGk1jc7Q+sWWi978QweJ0zBYSJBmFHJJNA+4vz1IEsoBnmUXo7fvV00jEAqYOER
43Htbr/hq3jgMwWX+rcdMlzikPwsVWqy+qRRwBvADhGgU8xgXuy0mlfd2Bea8c2UT9JGAkKQbEgR
2I+0jmV7Lptq25yUt9V4pPxfncfEoxU2ZYUH/DLpHouWbeMJvVze7NZbhq1V4fGFcrQElwSM8kZM
nKYCQrHgcZ+GpLW/44yzzP5IIjdQyZMBVLMDpkQGuSImolaWG7WnQ0SkzlYgNpJkEqJ0Q/HuGZfR
oEIYhLcQ1yjx0U2IkYbcDkKtEhIIcf1Y6b8cmOVQN4+Cusgi418Jx0dFu8Gv1Qswo1x+4RgwX7NJ
yqiG7uCRXmgFUOPfF3hMGH6OF0E/bXLjks+qC68lOuxEL7d96YxEZ0KXWJKyY8vUoUlE1wMf+yPJ
BsBp7YSlHqoVsOxbEGhwvo74KD7CH/O1csTB6kgfIxszjrKwZNOKdg6G0x4YsZIlqxSH8oW89XU4
3/Im9j/s2pY8xnhSZ0qzQM73qhkzU13HuQDKXUNp1H4Ok0FiAJNbhFZWDlimGoSns0/Dzy143YwG
dec2ZTZf17siQF3LUrtDvORT5BYxfUia8QqxyzAjkc9XZF3y4E8Llu5pqybEBTubw8Z+q2NpXApX
ScY0mWzn1+f1/ZeMd4HX+j9bkVBLwws/QttnCMB9DZMTaYPwee5Sx1yJilZoPIm16nomqL7L2BSC
exQIp4AQbL26IyV5J6rxOrrKAAPNe423ygLtID8GUJtBJyPWyuEkGNedpMW/uNlIK7IzNsOjZq/C
WRFK8dp9Rtw7RVtLdtaQcu6u8mtMpuZLus0spVB8HnjpX+I90loHp/DYjHyVDXAs2FtyqBG2QGKV
/jpO3I5LBXb0pua+vriEfaKHWqf5r+bGshIaF0HEByWqNFIY7NkHP8ryU2xKXdb8Nc+ul3Dn3nRO
t+9G63qzKCcULMwE4xLGNSvTrq0uOtB3xLqYLlixBHTKtdofg64Qq6cAyw0s1gDXL2qe1Edq90yX
RARKBwP6mc2b+0lsVuPy6eJwaHXLc3v/R3tpjl2L7zAyIYQchoT/aN3qwTjjqYVvueVyAvyOkWYN
3cX8YFnYZyC/75tkhqayA6g3sSfUythyl+rUrUjXNgErZ23KLAnKIAR3hAQ+Xk9W+npfuG1B3+mG
K5hsZMp0UlzgbFPy5OZVJ5D8r0EhLk//esyMGx+9xq0B82+wbGDZrmCEDSR5Mhn/TiucN82I/puZ
0KPrF4eB/h5cUT9OiobsZbyJOsIgueJO045FdFmy6gBNFt/1jOaeoxyHRMnVU3xcYWjJpmvLDue2
eD3cZ/YovotvdHMy9JnO2PEFOZupjvpBm5OpdJ4LMVCgULjhohni5bd2d317o4uHF+jo9rPAz+vC
joNhZcr2DOvduAhOu0RMwMLpciSnUYUavHrvyTZaLms0/417ahPZI/izibPXoGNrGpHVjQ+fAiXK
099P2KN/SpEFG8zTSZzAX6YbSiJCeWtFnlHuFybkDNNU8GjdbDTyCAAO7gg3tcfxo9k5q4ICZFS6
eRF6hwVkJkkzlp/vA+aBgOa/a/GW76W3z8c9fOiiUJTn70efLRy6SmYJc8gQBzFAkHpKgJkPwQUP
ohVCOaItER0QNhOgglN2xq0aRZ/JiEIaBegh9Q5v9HJCpa2XvCyNjIg+subQixod9yBb6P6K1Q6E
NWji8hcYgAMo0EdqPzwwVqZLywu+SePOujwJHLU4r9o9iQptkKz6hZevHbl/y5FF3nedqIKtetvg
uJdv+aTFv6KCPcVmJVaynVaNZnUn4odMOJGhM+bSka0EKSzArLyLc7GjySL1WYA+Bqoh0ggwBfCS
TWLxumJhlXwP3KH2Rwmj0dSlE8iTZatpCR/vepMMfoVu6SK7lvVrogHbzlxYGnCFARJZgRYlkRnn
qskq75MSsFFxvn/E1UFFVrVQKCB9k3MXiVvSqmVDyUk5n/90x8DZimccltrlH/qdVaKvWEvd89ST
cDmIJ0wAEw5tTi7jtykmmRhZPdNjdxKFDcAOZ+r2K5N9rXb8pRmkQ2SmXyV9QZWGuSX+/kZODyuP
QZJrQODZhpFuw+eJ2CVBkqp4gGjmR+8hiryzY4BblQmpPZ06MVYsOyAs5uuE2RtRIXblc4mGjS2N
G4ZrstPuZiSa4UZCjrPePMcOBhpELNe8EQf7grv91nr/oFTUWhBjjZjRrPataC9GiN8CpY0+H5BN
s3FULqEEAwEF88QWf1fyjxY3BfsP0nUFYuSxq7DleKqbf+8LsPNXdC1HIc5prLv/aWwpAsQFKzu7
NrCUYwol1eXsBUf7m0Q+PlIONy36js8za7LvVUcQ3UIt6VMSkrvjIijnG8wDH66+ct4+DzBkLWIg
ssBw7KotGFKeQPnPxMnsNVAtEYwjbJATTGwm1cet0AVk51Q8/hdPkZIXWO4//YDORTexL2G4z1Iu
fHSx2wsit2tS4S/FQ4lAg0pgENXmH8rK9WhNNKK2jn9eiD1GkSPI77OVPLWl32+rT/8glgsx8aaS
5zk8HwgktHNiGYHuXyXQ7pXW117+imzexXrhdIhF6WkydnpRBxzYeVU8ybOUpfT7JkRixQpFh2FS
7JdzUjaHc8oqnbc4rFRKWlCLA2waJJ0D/NzRJKtAXzELYuOqcExlpQkSwzlHPsiPUBh/Dy3A64jm
tG5MCeCv25yL82XZGutZPq9f/jUs4JPUg77WGWZjTnHSTrnirT+FV47qNKHdpZR6eS7W+p033d3V
fvDyfMJYUmp1BZXepP0JUGwwEnx+B8gZQDPyZ697n1ue9Sht750bI0IytK3Lh9mSpgZPphA42eMd
CdvKV78PiWQfY9qMw/rFD0XthWqjO/PoTOpslqpyAJm/u1MHlIn1/0odEA1M5aalxwCQ/KGij176
+96RG5r9r+xQR2f7VXiD71tJvi4QfsFpkQCXR1JElPGWdnvVZq0H0LGpYhgGNDeJelv6BxLXb71a
hR13pyUbKkeDdW+LIUb0mN9xyQSTefRwdIV9+SHH5K/eX4uFFqzCYUof/XaIYzs7vVhIy3iLo1ui
xIiN/pK5lCqrAnmeLr6EFTA5Ir53CXzabNxfzUmyLIpCqMyMu+SvierIkm0O3+6pO6SYDAREmYEb
J2m5BODqAvZGt0y3Q9O52eDDlObTEUo19up44EKMNi+Br3ukuh52BDH3VwxpabuJxnlbk/Uw37wA
9uhYYAn+T9H6oW9ihYw3hPOV4nOypC+84f2gBDk4c6MKQoU4MlnXmTRMSji7W9E4XTapLc3DKmwR
1cvwogQ+ag49FxqPNmob9AJDKVkNVbYnN/GCYXo4IQIRDo8CEGH2i2DPs555RnV4v9a7IHr2Jzv2
qxa7vRl1pySDMpjgyA3wNoA360setegMT6n9Igv5y8X6LrZ+CEGu0xjrb3CAl3/9UIGRJnSv+xjE
DSWkyN7omVrmIMSmyGESYpinHHSksAQUmJ6T9Ecg+DnOrBlQ2WlQmHpFvCCauUpJj1tS7qlrvK9H
3iEopHF4tRxyHXbBMSBuz2hOeaakfDhSnidmxHU1xbu51dw2iF1fIPfIZ005oWZpYJShSkbRkY4v
DAZjTxiXWQBvWBY+taNGxMn7oWE/XzyLvRb8TCSO1We6TYkD3eCnovZWfvjAuD0b9JuLRzu4OMzx
IyeADhjAn+3dHOirAOaYVZG4ZGDKuPJlCe4vs8suoPCpkx23VtAJDmFsHG4ca4jsKF3bKf4eGgW1
Mjc1G+5rVGXI1tVhuQvoxcl4XFUAGsJBidHHg6e/QFk4CSXEYoytP97RTuhqP7MlfR9i9Nhyq0o8
6U1Bwfw3jgl6svp8eEt/fucNUkuhjxwTS07KMWyi/0IDDBJ2tSOxIeSoGqY8DhkuFfv8KginV+hg
WN1sgHwdElzAHePSybzvRcnrT3aNDz+hRKjYxsZOwK/9UBDkRuHRNcuR6IKa2kvwBB8cy9Ct383m
QoDxHQxgWMMaBLMpyTdoAMK0L7Snjt+DrWVFDfeN0A0zdiEHPvkiUx+PdI+EQ/petB7A189cf2KO
UxtQT+fXepsUTVMYsap7E5tJjMboepFkeZ/hAEmNOJS1RU9GBkTFZ5j3R34bgo70SnH0db+go3Dj
TaGfXqBhsoku7XI3IFYdMLteguQgQeTm7F9VPaeJxvYqzacFb17Qzf+iAJyAZjC81sM/UAyBWPih
8C+Dnt31sg+4IpiASjoiQ/TM3FjAuejpsXLxr3Msv/zOu0c0pjlo9aQMfgKaQm91qu2YllMv2Pyt
Wn9OE0ZY6EtnVbL4MRmrPuPsyfLPDh8/2azn208zmwqn80/L4yvceX1EI7sgzAJ6kMaRtOtVwMF4
W4n6Wbc11CXlHHt5qWAQiqrhfTPgWtR0I/sy06rpiOw2Jjw3g69TpcSHhEr7xUdxCLa+5tvd7ddr
iMl4icgMf9VVnvMWhalXoe4lHNceC+Lh5VAJCBZpTjjEJVpS1HX3fZxrgQdY3cNIfbl6gbRK8Q/G
f8/P0RWsiDaKvMrNXjQSLTMJkwEiF32E4Qh6fnvU7r88oJKMStt5oi1gWQ/NGxm+EzWmjKFw4nJI
7Qm/hlXstnxKoy3VUbzDpEK2ySpLeYgXYTBPCgPlr3TFxViY2jy5YVxKmYY3OCGIorvKE4jLIbhP
Y+TOvn7iNz+roSE5SZm6WnWhz80Ne72QU5MKxzEj7S4U8psW75xLXG96DTJEoQZ8Rkmfqda3P3zf
QHv3RiaPuIwjL2oipfhDIGnWn4V8k9rMcM92H6r2+KAfcVEYFGzuyJW7jIJXLJnSzjWR+1o8hsTn
qCDMfL9l1f3TvpxT+xljaYR3m7V63N/6IKRkEfWDi/ROxk380rcEFa2TnrnBuXVLiqX1Mx3K95lY
OnO6VBkiZe6Zlx+9jInnGNFBBNVTSOLV3K1nc5God6WccMKnzqeA4a22QQi3bFPl7QM7eEerEdXz
LMW9Rzvf9YGCbBJ9oFpkT0OSdEb0PK3U0KnGgTaC+h38aLrI3d3Zx2tBNr6mf08LVHMIlERZCf/f
6OTE5bO4vtWtYE8ensGVRw2BzOGtUzJcRp0muYKoetHqCFg/CmwbOk4roZXXgSK6PNP/HbFoe8XF
EhEAXxNWZJeg9hEUs7f2Uvt5HdNrH+hQGtxlBUuDbZPbpUZoht8np6dDWh5XdnjVV8OyPPDbrSCU
6PqbXxTWPfaicqzZ+TBOUPsAYiiBvO76v5046ylxjAVL0qkB/TichX62fXSj2Q1umbHF6ElpFvSQ
soffMbTeknqIFLIb/7NJOgTI/eGyh27dHT/qF5ku+B5K64eP3CvBbA/Zo8ChhER9O49V73bx5geG
wbdF1bFWhr0FYfgp3TYBDrRyREI/iKpuHXMflSk+A3VpsA7//S+H2cM+yOrJSEtu1c+gclaMW8VB
kuBoWrgHASGoSut1z8fBdohoQJxnDQEofrcRZnNNOJtj1aqAKlZWVyj2pGBcsxGt/qwwijxjIgQv
HSaZLgtdSk9/I0pcGSK/chAuezl5ofLniB/WSobAGiMftrrh4YkIkXSZkhP2E4gmEEebDPCqpwc0
/1Qz7ogAmfi8bgXBPl6g6LSC2djUDPouSd+J+SQ9v19pz3V89KeQxEDwjkMIfGNSb1d75u2gNtSB
e45GgXNzkF9Ic5oCj65zpek0lW8ROc7Yzjnmens+rvxGnK5BwXE5X1hAyfa6/kFiSvqbdKNxaMIS
FV4FF3y6VAlBeo41/GV0Z5tsDH62/fqzSEmJrhnHNRGV32BdhLI0WxVpR9iJHBlXdWSnTSqB6Nxx
AjS0oU36m3oCa/PtYcssG/b9F+weDw5BzxVdMFyLi34nJ1Vy1P5kmn0ySJDl5vrAVHK4fK0cX5+O
cs9p5dosiYqMyeNixTIZTVVEO6zLrTuIsm4+Qkx5r2nS9BTRMKmQG+CWbzRehf3ivyWY7TqOA+N6
rseqxd3C+EQobNcCllH2PhA7cKsZIAwX277BRY9ya+n04WE754E3BsI7hCUS37uif8mcsFsgKQ8L
UCQieRH75tFUI+RHAUejkty9s6XnZmIUgx4Ljrk19RsDHLyoA51LwAmX4Q+QSmAYgrroJzC0buaS
Ys63OnHGYYsRK0ltQ1laR7Pt5Jr8BQOwESjwCEKQQ82yH4Ul9XnixuBdRC4MX7QBiM8c4qURYVTZ
kY5m54VWOxbiZRtoxkTGC5FCfWmcP0cKZ/Zm4ybqqc8nkoN6W3WtqkCnw80uEzo6eRFpQq6JN2du
FGPvvgnxVurQQBprTfJ+I1LX9FfCT1oBw+9OdSn0fgvsdyD27HyjNDG0Sd2uR9kLRKOvpnZeFBek
t+A2NdrpsIylMWvIW1LuCJDFulJZS5Jc3iou/ADZSvnl6IDZYgVh9Nq4N4K2TPWtndtCoRhJWvhL
r0hSx54BkvlCR0P9MZmK7aLEJ3On5oFDlWr7O9AzRZmr/lF0EalSIcSmDT+0YgauwDHVulIlkctG
uJ9ku54Kvn01ecSJ6Z60z9zwphm0GADqvEcmp3uVZOebFafP3xkPYT7GCr1eGj4507WIIF4OUOvJ
7OwXCUwWx2T0VSgjCqwgUkRCAhMXwCeKp5xODomqtceE8BoKPOBwxd2UB8UpO6KA+i20ZV25YTw3
cf85vU5ym/Ux4SE7Oej12NRE/Z0u5TsQ6nFnY7smkC0cwDWXnA2aT+14fl1TVO7KqpwrwZ7j+qn1
Pa5Bl3IUGrh3jPBH/s9ABC1ZSnvhq+aZG18arNltPGzwXhHtwjLS4rsW5DUJxeL4qyS0oLYVMCag
189d0AseDiK+0tqFjYuJP8JKTbgUr06WbujCdwvW7d9JeBjzsremFmq62xPdr/uH6WwkQr/PLlMB
UYh9z0+2D7KyGH8Fb1LhmM4J+GZqtn0Z70bWO98OWGIW0/gKyqcqV4mZtClvp02Q88MQ7UmkfiB8
1O0tzLq4OohjI3kn2tksb13Rk6TEoOtmsok3Ty7YnzVXDV4gtit6ceLXG4I+Abzq0se3eJxBSgkD
H7cqSFdYRnghjHG9nU5E7cqESJjM/dgFMl2Yo4O8eX0f53TE2CMHXciEsgdfndxuJrKC2WJfjZ9s
AA9267C+/AKpGOIvUqoWHqCiM9AJhni+VJY2hYJWLUFIAO6xCRIfbs6DwL5gntFnacZ5b23VmbCj
7df/Myo94L4OaTBqtgkutvBobaIf8XcnHuA+nwp6LF26ZR19enakuo57oaS5bOdBePApIbKouCKk
wYrf9IaBPXUWesnDe2m38EOZAdxnZBtrwCKB23OC/lVbAZ5FncnzTmt8bKfBNzXYhcgT+FBQ9DHP
u60GYHiP+7MDywIakFD4QYODCCP2bCMTyaV//+JTGBLeqONXSl58PAmeDpg8etfa84BlZjsUhYvM
ZRO+wEJ3khcJHuQmiRL7NGOUoHTcYz3z0IwGBd9Urdr4NOrkMYia8PEOCeLfmLEQUHjpW1OQLiXg
yiR8gtzabr9xFmkyQQn97+/JabeWpiv+DVeNhkIegaUAPek6lfVQeHT4zP3gsfaWBVb14AHJc11U
C1i6rqAzQ7I72SthkewkrgNi2iWNWzY6uSnbHJCGQnTdxiNgXR9YokNmaBg3zk45mD+AMS8cB7PK
TRoWdDhL8jeev9DixNGc4eJnRAy8xxWWIhpVBY6NzXU1R2pQ1SkPX5ltcg3SP3qzTDrY4P8a2Le/
/yI53h2Ht9Uhl7kqmA/i3QL1440Aw7kq+WKJWk4nH2CnHdJvz2A+khGH0mHjKHZTKbfOCC9DLTbY
qMS9PSEjAl/7rTpEU/6U49Yy84at8BQCpzQEQoaoVd7wXLPmMrU1Aql63/2xuoGmdAuDlFta19BQ
RLqk6VmyMkwW+ea2+cGCjL1qVY9EIdpLfeD8A6E4SVq1NdI4gksa1YmCnH48t5C6+v1GzrJipwGg
LUHxX2yBzFCiA3UlXq1nFUhVbT8LbMX2iH9J/k1YKPgDV8Yw5z+U/OzM3DdQczkxwrdGa8ufWGk/
LF0cDULqxG0+aoMHGMQYnh6oeF9alHXZ3PL4mpl0de4rRaC0BF6t+WrVxtKzoLe0ZxU8RzA/eSds
hpJ53aPxB1M49d2kNOrit5kE0xkCJ1zQdkJc5zd5A5rDTVe/++IXFFPE3VFGl77eMvtmkLkRaT/R
dRN465gMGd/2z4wFXb5r1Yc9kW6GIXGeiSUB7QJn9ZPokQ3O+wtCsfuH7Z0OfswB5EIdvDHjFl2/
y/ANZardpzkYtjPy6JcJl9z3HUUQBIiUK4awUyjynocDougyc4dOEog1Zn8TqUJrlR8a7KUrMTp2
YGfwZddaov8Gmsnl2Pjy4piIuldln6p2jpZinpidGFsI+PQOrWGr6EIh55rRhS1tNVo/7RFYYRd2
vqCDVJ0FLUxW1yLP5fozRmSsis1UMd/PwH2c6iAsg8X54NxJROeagQIKPVXmCkcZ3e4remHvEJ0E
zYbbyQOOGJt86Z0tiJ/4Q4RcJJ731yeDwuPLqwTf1M3wbIuVJfN1g5CV/06Jy9g8T0kqHM4P9OUP
ZOgdc5ZUd6Y+hMUwG2b+hEbgfbbxeQJDK/EODjzP/Qc4SiyBiNIs1tHIXhzakYm9Hh2WmnV2j/rm
hjewRK87Z+0nQDTo/QXdIsvTQwlb7DAtdzXFEQDCCJAnm0WX4O0DuEfpMou2KEmLFhyOlZq82j90
CczKQBJMtFARZjNZJO/yU3w2IEM3R8AN/8ZJ/FNpXjvETyTqpFHxloJHxnd5XfhnqqRsXCpxNFMh
Nr5/DBaqeb/Bffs4YcXsgO1yDJnSHodYCBxijyDNsRLjIZ0IyYlu2WC0pdKI0eNIuGra01ot+TAO
h4yaqeWyKXFqW3gSKNUWJSqorZa2Gtr5+7MjdWx2c601hwsCMdQNMON6sJNrlgPxHJqLOY4XBJBN
f+H7FB4gk7iz/IJEu3hiBZT+Qo+nekAsZWwl19QE/CHDBpCA0vCCgX/ZyDKJmDxHR6IfSbnFArhF
SKX/ME+0RxmkCKB8xVzREKjAdKei+kxYI8kdrj5sOMzpDJo1x/Xwha2xcDjmYl1unW5GxE5WRWLI
YnWmSfT8uIASpMRdZ9R/3mfMEdYyJYBVYpxOn0m/IwCO+lJvnH8oxg4ZtxJSDr6faj8vX33PGrlM
MnbjPattAnRQzzzFp8ZpWdpHVDsyoX9RSXAQObCtSACVXHgL4am9gQuOn+D+Vl5+4OMdIgg/PsF9
sXBH7MNEdSxdJVYLbfQ/Cm1PBGiFUnbIXHilHEP1jwS9qm4zLh12V6S3GeyHZ9tyR2z9oaELSmAp
g8UcaiJum298sWlsKZhJTy4NH+iU/FKiQbcIsasysOFqbn/Pn8mexhSuh7Pqbq3VLlW1ngLz60a0
nnoqU0V8vCS6Yz102N+Ce8lsktWN6gYo2i2iIotrBa3XL13ub3owoHqnGMmVlsMh++skgiIm/6aB
tCA0j8vxqGXnJgZGv+2maIIbEv5oB6j4jb4G95mkmbDrSFEHWKJyV4428yXDRlgI3a0WS0/gEk9R
Bp+DnrNAWpnvByUJHu/km/stBHEo8LmTrMQA6eLOBoJfINSUahYIt0lgGGhaSjYbgGdIxjltjLRf
8rWlp8DCer+cHO7sJXFRyACznFr8IB405Su0pwOfJbJEo/smHW9hmq1JUqLMuXh2bPHsQQ39p0p4
eAtmuSEtGCX8YgtqCtnxAYe9mhX992KVGHFddfSw5XS96YBa0+HvqYlOfxmVFE1IeQ602xar7xdO
Xs8dOkNWO86t+6kBLshIlXOl9zaUY5y0EKxEpNLE+4HL/UB0+Y5m+eWlqP42gCOteie5MvWg/uI9
DZiDAz4Iis3GOekNoStjR9ULNPqNGqEZjRsdmbMqESjNFg/V6VnqRHoahHLHiGh9/GJ8lcqFIqq2
THEHZl5GwsWNWsdg7llIKrgfmgstJGhtDBRxiHCqvgcINUvDVVADoYORcl/w4XoQtD78w/Ar0SIf
KqdaxvzZCye4xnuZP/wWXvwnozuIsfx1rNIziL1dNt8ca2hfB6obRLv/T8+U/6OmH9kB4WxfnpOg
n0npmii3mHAgHdAa6WzhRAtLq3r3Idp7MoB4gDYsHCObwH4QmWNKOCnOhCXGOmfIjL6XUunzwaLs
r0/LW8WQZvcZouUzaI+tzvEoTbC2yBluX4VoVtg7tmuUz7MJ5AI5Kma7JMkn4xbhSqFRNWO76XeL
2T7OKAHVyJnb8K0Q3bzUd0Uzma65ax04gXOO7vvNagL4AVH3KZ6B0ULEhp21xiZXMiCfkcZF6c51
MIOtGDSc6Y0shXy+p9bGuYYZUzbTfuZ/ZNoUIFFTQG9y/J2nhKZhL9E/75N1Kn+JOEXsFew0bPo3
hXVpoKUeG1V98sGdxAFuK72xRKIY+63ceYs1A4c6YrCnVh5kUgenJQQymSezTScW4EoLcruBg3GV
txDMafzXvQD2fchkr566m8sANvzo7YICn3p3fdcR8AJ1z6NJz4eCg+3UOYqQPMrGmjt5Z1hXq74J
PcETNK1kiIvuyKOsMxbhHWI+Wfomn3r9HkKNqJb3jGBxOIghTzIv14s2mC7n9azpINE8AYMBHIPL
XQ06ge7OTgyJQW6Cf0zYpszO5Ke7o4uAtqrnqfd5MsknqVBe53Dknty2Kv6lbWeYgKFE8mn5U2rl
nSbEPg8qoD/8n4YLMz9aV3PTZG/ppeHMxjKkA97QTPa2qiOhCXA7dHuGoMJ5LM64IW9x6H4BEeAE
POtmEIcrqDOw/PrN3RKv/PsCJHsycHbjADJpE5o8EdmM0zU4mHDs2skUm39yOMbqZCKUCrb1zEtC
piYs56R8GGOMh6U5jJRLaT3xjmoHIP8n7i36AXrS9YC1B2b3rLigZdGR1T6RwmI7JxVW6Z4445Tp
ftnVHcMZ0pGfFvWV8qr7G7qXglcF4CWrGTlND9KOIGXlY/DFaQDKCN4oMCdNtNe8DIuQkyq5wj4S
8hPppq53853zAfdWINW+r3ODziUZw9Uas8TMr1SndmwZyFPh4fOYnlgT0mUdkv5oE+4TIG1rTdqp
l6V+P3jPVz2HD5HWb+MyxrZ2yezv0k3nTO5EKMYqf3MsL96kioiVg2pYrO6N4y4AEC6LdkfArjEn
/c5HleP/mZjwmooHW+Lxoskvu9hiNnTz7MjuOdo/Mbn6f/R83P+cEhyT0gnCklmBRWO/FI9+dWhN
pmB46e/B5W+eOL2FxAH96t/Y89ZMEBio56n0oxVP6yU0IuyimgjKAXDSYGyikbO5hwagxI641oiX
rd8nV1hqG4w5k95E+fI5mbhax7TK8QWxnI4u5EV6iTlJT1TpL5T0jkLfIujQmKF+X9rqiIlD727D
lfT5+kuMKNhLd/LSMp6fHL3yhi/BlDN/cj9yf0klizJ2omHPaixo4FhMVYO+dgCDWvKjVYU4GZh0
A1WcLNAww1opQMNsmtoCfS0vfG8oOI11GL21xB2R4CheIs2P+LQGPs3/vuZcHvwl3g2tMg3U5TIq
+MFfmVrV89nLYwkuu3lBe4KJipqkayoz33klEZ3qyrGHN/1WXtVWo0zSIjNyEzesv+zTNUJiBabn
pPbXXsqtS9p2RDROUgo3+TLSR4rGLOXjWO2qhF8v9qEezrRAaid6XAnFenuHc4/ncfA0SQj4IUL8
PGZfiYqwEzmklNwg56GzQXOBIjO5E/tbmr8RNfx3It5QSlVISQ58KN9wI7TgkvbyWU40darNzSDv
5v+O1+C8tLiMF1d+v7wqUgg6N4dMKXDOIOz0uKkQvqNYFBjhzIeHBA/Vb2hYzB6U4IN6V2PD80qT
RQUjV6ctq8emsR8kvEaIa+cbZwSwKw4e1LNKC5d9M0/AWdWRZjHUHId6LRI9ROv/dWalL6nOHVGU
8sxY043mfc1I4/o2b+wM5KlMdOzcMAqUcYDyka4yY62VK5tz/Y3OeNXeNW/oD0mJGnNnGGHp7vRd
tnHx38Og4SVRXwf+hR00080/7P4AQOFatP9cfkVfaxgphSRMMUEs12IGEa3hbvSJF77aRONmu7TW
IjXR8uOtpaaVn1vyi37bEwIFZyBTix25HJzzy48vXwweB48GH4yoOQM/P0cFAgaAej49agaiuq6S
IR0YTVsWzek1ePOZ4UER9NxXk4oEhi37nFJmkAyRRrn8TDaMhCzv2eOGMp6DM99yEexlv30uKTab
0F3wGxYwFYBRC585wh0V7kUVUEk4GxK325MxT6MCG/702lqW4YIZtFpOXGj1E8RQwE/QVkFqq55h
cDHB8JiHNx3IoLVt1T5PvdAkM3Bar6878tLSPsVqbxTvR0NdBC6FjyAZ1cyZmqg5dJPWEyIzjbq3
+b+ryvAgPQzbxTmzrAohTWHGxp4jdmhBBFKZUyF/0N2NIpJKA9L0tg3OPPVpklCqwcmm5BMtC77D
LdQuxfkfPB3z0xpkakhxrWPL5jsz58DFEDGal4gItuebweLcUTgX5ChAojywtIeUVeKIORdt/HJs
4y3srRbZZpiAY8qaqX+hEL1OCar+dNTCf3fOIWkUN8ZBYzJ8TYtN1u5wN6Tl/XhpeuQiknU36NGI
3dkfA6+tcSDg9XNJWXF7u78ikwkN3o7YOo++B+NEODITsNNHfwuowxnfpWcpqKjOrrClPfkLsrai
r8MSmMJnPOU4iIOoqEn3b+l/diqIUAuAHixubAaYHo6CL2KAxLONuxPFw/xrByVQLVyLjugXwses
1Tgq2zS12rRwCU8OmTt1tM9BaayTDtY/a5rrCJfxDxtcFY2ltvYk4qDU5lwZKyYT0VhdbDY8oMuv
yiAX4i0uFbeZlYS7TFpLcGWHLlO2MIVRujpkEzntLJCUsaEdS9OS+rS3+INXB83+i20cG0H35L6x
/iRL13Ea4CBmaL72ZuVGvJ7eMFmo9VD7TlUBQmfRhnScPklFoQScv4xMwVlXeFSWHZO6ikxjHh8a
K5W4v9NUPlIA7SsR7f84Qz3F6yeV/k/9IRIrb9EPkWPi0o41uz9fmLLCEyGWhkw0xCLhp/Jc8vUv
p4I9nG02Ptl6hlwbPhFIiS+eBxNBPa2BHhqOtE6MrvTXB1h9lIfYUA8X3XIaUUIwf7nN6QugHB6Q
XUO9tw9fxF2XeKInH85EISkkXmkiCqzE+vY6O2hxugrDlaMc7WnM4pQmvEUt47P0kLMsBYUoChXN
6Zs05roa2MNPGYzObvX3h22lV/0zaKHnUyqQPD2ilwE/gVSZnBaNhlPiZFeUSkVxPbI9LkjxPY8t
1thkDUCJCsLSTOcRkT5HbBfxrZ54dojiZjn0IIjw267fm2ce74ffMsx0UY69HnONTgYlJ/1Z0CRJ
nLeq5QnKsfPc9naG3dHBqq3+cf0ISZQCui07RkkUeBcCVO+/MdYAX1b5G1LRpifEHzTVrK/r4rcq
QoOCs2zNXMsdDVcSfn5fecvdPWoSrGD1gNNIu/N40QiZ0l/ojvQdW9gl1RAXnHOIbwhhyv3xdtgF
Od45Mfy2cA6YckrmFshPdGwVOreqV0BT6uYPEi8iDt2h4DhsOfpOzvlBcvFsjGMTAsB/XgToA6zU
LHjg1s2rni/CwP2OJ6pbML6enc0MhKwhX1dym4gvPgAWbBWuIFlI+Et3ZZGTVUuluK8w1et0XCep
f+6B1kc+teZCRZ069RfpW17yc8Bh/soeajPegIETIJ6gI2C/Q1n7pUfqJ9P2OV0MStY94bTh+Cti
djl40ArXlhURYuYc7Zl0diDxG/iReZDpIicErGEPGRVR0Ev3+m+D5nToepB19cqrV36HVIblDQ5N
vp3JeKsuDai7xoADeeSxbhGHT2GSNSyzAjgBNBSOvsgLTT5cdyZH7MLl8AWpxslLEeHWefDDBXE6
/LEeiLRpLsmNn1oV3+0GdTTJvQAeaVfSOY6ZUo5zU/KpKa8tbIrSRN7ATOdAo8Ta+Gb/BFbsvt84
vO77P2djPg2/eo3cHRwuK+89eAA+E620Joa5DST/ee9kOiv/HtnpnyRLnIGbr0NhYpSzYSzvpxsk
HmNoqVpwjlAsrK5SdDhBSy4zlyL/jJSB+eLxw39i0MopLLi5TG9asN1ttjCXU25xpxstreL3pLZn
LruX5sSNkcpFr198aNupkEblwmMHL2rRF4UWf5gzxdsuyRe9yIXaWN9PSHU9rIknNLaIdMLAnTG6
iAXV5nAQHE5A+iqCc+ITW6e4sSa8PdaY0VJ4HZ/3nD88n4JnDUs8lDDdRgA3RYdO/e7T8oZr5s3l
OZ1tMifqKKWNmad2MZMYP6Me4xIf+36WMzuNOfZVp+rPq5lY4AQ0ivgzAOEOrFRzJfKSVepx+igh
m56+VG/zYfGYJ6t2bdnbCroyKC0B7P03i3frHNIfazeRj/lLUOiMbCjmlF4Zc4Xow8kQzedi8XSp
GYi6DI9ng72ojjr3o+HyDSXAj3tIuc2JhnhkDcahm2IO3vv43U1P2Sz7RGSDswykoKcx5hu9fmDH
N0J6UWQQDQnnz75V+uP3H8O/5aPlSVfb1/rAmNdPSDM9z4RChFPegh3imOUocpIFMBwvQJEPBKYh
ed0QOKdim4GZXdn3Ymm3TUouArQHxnCI4OuHpCcaz1vI6AT1s+1PwG2dk/8PMaRieKryQWAm1PPM
5ONu2IhxyTw6OU1v37H1JZ9ko3WL7+w+PQuWb6QpYx4AyUAh0PsxkPXVaKghWvx2FSW1VHRnwukR
k1CTBGLQEulpRC3dQFg8Y9lu41gVigBxGeNCefMudcDipcamgHtlBvZ4t0v582FZXlWpnRQ0hs72
HKBj6fK4V3xVYTGreSNvzPZLFueljmRypyNtoAyLBqV3rfeeHKQG0cJ/knjU+PUmaDWVqja/XGH6
DFM3i/3YoL0p/w5rug+VVJhwbsRtLQM0JpL1DDYnc3yckaNtScs4LoWQ4HL3D1FZ3X+Hlzw4dSjg
SNBC5T6hx77DbIWK0RtHWomq9yiz/IVC6jeoIbe8iFL6s2aOHWT+7POAPCyYzp3wihcP95sbeW3p
pOAfOpGslvX6ereqsifoWwAQPylWx8llVALwEABp9OW4z54Y79LfK5SR8RixxvodMEnxvy4ZoAyL
7l3o0FWnsep1QCbyobnvhkUJb/AbkIadgK8V/EqG3cxLTg88WvURUh/x2TYvUKmlyvNayhKJ8Ip/
R1F1DEKkWNS7jlvyvNwqDS/MZpc2R9g7uV0Zc1g2R8dGWb0Faw2jGFy9as+XsZuADNL37RGhQJvA
/UueJ0qLQfIOmuY6rdZtQZrtyVr6SZEMDJajfE1lsM8pZvOLooE+bjRFk40BnERRO6ufiO+mjWcY
JYJEpuIkse4xHns0c6OJiXV/Jq7/JpeT6OPwgnFZl2DCsHgUHkjiHTFLV01Fk/Np/8J502W+ShYc
MbV/B42IZQc6s4qMJTouZ5KR5a35MfHp1zAC1Yjp/e3bORE2f4h7q7hkTWXVlap8rP64MW5bHk0D
eKx4B5PiZPbufa+F1mtPU2um6zUFj5lIM0PcAYxhEw4BhGTLumlIKMCHaApQR4dn0iptibfKoDhW
bSkvPWVnuuh0b09yaHesJoSLlNlkwpnUQNKuQT5TJDlQl33bXSB0BMyi2Gfgllxh7Xoc5gx+7UXT
EGubcXAJs3+HICU2a6C1lqJfMZxlJV/WZGM1uMRa2MDBExbZztrTZMpN1JWzV/j/FPC/fMQqA0yP
ZwZ8rTcKQWfksn1dXYSndInXOEkIWN9iOfYzTJZne+705EuPELWPwwsynEFc5TFo0A0ezNDhdBWY
MQ/hRzf1r8m48UQCkKyC9s+HDsb6IBxjAwUITmJNQYN8Bzhv9t+EwvrfCzViLpdKRJf811TX3JjI
sYYOtwkjK7VTENvMVw13s7XCxW0OAj2UMvPsAnvWvPLa8UQtaC2mMMWkauQKUoO16mns3RZ+LCmP
muyo2UrvOrThfAI/9bY+zRjbJPgu4zulcMNOKTvf2RsBx4qmk+kJuK0RC0W6fM9avi8WWdUFmjSU
pSCZrXKcWrihNVkivJdC8yWjieatjNZg70HGMSpHOKpPbUu8xHtZmj9qtZLDlpyLaa4hpqzlp9X0
BkHPb+gukvEOLYNQHB8h+N/Sj2bnTkvy/MXAPtIJFu19/XVBqsEqbRyYfEc9gNN7kyf7nJijeTnt
dSGsE1HgR06rCZ81kupN0qtbwPkipfQjyPH+/eZwGnkoHU9MkT+RPw0SR7PYbk+X7iAHlnlKKkMv
HMk5a/nk1X3zaQGv6Ag4DGgKVFHEmAHYHhRvNwSDdWwXI74oHlhJ8nMkiH6LTsW0ep32X5M64vjR
I65+ABc7WRU798dNUDKcssltXbsCBqZKSfsGuI8bYzvZiqpmREYDmmwNYvG829y8IPdHEzK75Qvn
T2Re6ZDUSz6GDTfBgjdWzBelCI3VvAc8eSTqEvu5oZU08uYG755XmtGkEDP7p72XdNZxx6PY9xCz
vHL/p8Trf31+7l+lMtbXhNcGUy1JppptCs0ly1h5AnlaAkvt8xJ2Sp+XcOrSx4Wsi0IFzkFFDyJq
MfvI5JctfLZ19fPnpuDBxX+cbWLheL9+N+rt/h9NG/v0N/95zJneg8+7zc94zSqXOZu1V4HKhkNZ
cLCpx8X4dMQ0BwHWpFvITKjtXpX64DDObJktd+HAYIwjsuXVSFwfYLnktGSQQQPLaEIO+YjLu5+D
EqI7uIGMk71kdVi/CvMO9nErbDW4+JBsv9t53LyOG8ubBmJhM+tmgcysVjf5Vynqz6MSVytu329F
2p73nrJ/F2SfmI8xs75eI+RnJZoEUvSrqpTuMy0vTXs7GfOo+dci6GIDcy/mvmkYEIBhFvWHA8Y1
A0cGc2oXHdvgHEOQGC39yX9zISnvZhD6dfXLOcUB85AKrqplefvQBjlmYAt1BjRjX/v/pM9iEcIQ
JYdmVP4PiEEyS4AH5SM3Ua1YXgBECpZ3JI0XPAD9vi9m8JHMwDnrmaHMlRBSKU4y104/emIr1MiW
lQtGKnCQRB7+AQAnnFFXFIkW3tgcsxEVGonJhg/7GvfgOwYh57hrMOIY8OZ5ypUN3vlJfdC+lyVK
npx2+p0Hh3Mqxw0VjOi7RSO4Xuzzs32Ze2SZVoiSvMNTN/DM17Mrr6MvrsuPkPqeEA5MOT5JoULY
mETYH0E/j1k199xjKZD0FqY/j99b+72k/x5LYlQnjvw662UfEIpToyvCJdrGkOciS+E2qPMA8/Is
Ns43Uk60dD7rHxqK9UeHeuhm8bXtMf75esjh1eKrZCHfecn3j5KtnHxP/Qj89QaJ6hzVOutlfhYB
yDRji1cKrYk7IKHKkYV0FOKEXiJK5kmvKpQcZgEj2fwkMYZ9mjVvour7MEIcMwYC57VQYw8Lojk6
Cq8711vntNkHhjwST/AOlQFikZIdAIiQWHFldOXHU2RAxXAGrUz9jg2h/YFBinQYkoZvdCRieQ6l
s+O1YsQ7ww0g3Vj5Jv3kkCp+V3t+d+k9a1Kn1vB2SIbH5kBi/w9lQ8Y4jC43Skkx3lxINgrb35yg
wQuYhrJNrY4lgZ8754gp13T2I1cCiHOUjSugK5dqdCjrshlUNeTafB18vE1I9YHFy5sXjr7T7rUx
rj9ZQO81VyfTIa2Lrj8K7Ca0ZdluDNWR3iyUfr1m68/sl32pNZmNGobukHTgzqMWYK/XuyWw8wrO
FJkQKui7lcJVW5C3VorDWKiG1UNSgbuygrxFZNTwjLqaresE1hQxsJK8KXL+r990FM/FtjKqHhPn
RsJSj/TRh5Cus2oAYFiE2n5X45LTqMhdHEmqaAyhJsANPpbZmtu4FN36XTD88qoFOOP5YHzsqlNB
xuB643O+NCWIe6lzXy3m3W6wvbuohW/w/9bo400gV++YU/mMB0xsoLlg4Q7mGNhqoIaVnu5ztbOW
WuqGTBIN4xbxhcGcBCGQCsbvo/8ORY1ENpLd4oQzUECSnzGrnYz4Ph3Yi5UAnVrUaRlTeXuVwdlb
Lvt8uARBEymF5pM4WLuF0p2RcSatvUx1xSar4n/O2Z2sEE7LxLzSqMywZb4Ah1PEcfxVo3bmIu5j
CgenUM2pxMW8tU2XZHqaC9KxJgPC7/TO2hqHetaUs/ZrOv6A75+ijC+AA/rrAB3M4Y0fQVNUp+Ja
aj+UiVRhm51sIUyQAUm+j+jvUF2sqxMG5uO+CmPTZMh3fsU2NsrTWeJiTjFSgigpAmYJ0yqsT6Pu
vgbn/VCKD/pMQ5HacT6m9KE+r9qvuQTrPVyjY2nH9r/Yah9EWXlQ+yZfLGYM+RXxiYgQB0dlui9c
n1KuWuGpRm4Mt6FUuwqWpRB5RmBVT6Ye1OakFQeNF0XD2klbdDFxFiA2A99Cm6NrRA/s9AKQMlmn
Nx2fg0UUUU6ur5tw/XvkmsLJdETqZ43e1UB6UdXMH0+Iai8P4D/kH8r5xkcrMUEzDGm41fsyJZp3
2U2dl/7efOnaLT2EwuIvV7d2QXld10CQp2X48DyYgrMwBWC+BUdX3gWRhvnrXLFT06jBJRSe28Zp
KEFYDjQwH6UQgAGUMGgeAN8x1XU4IyVsdVY7xw8acRGJ0sHrgGECPbql/yxIITfVEFWN8KtgrkY1
V3mOJ5T6bChJHJfW+rlmsuzihP73T4psw7bhnl7cGxI2u3zp9wzEIBNt4/jxOr5JHGxKcZLovLG+
P/R5E63G9hcumcdLvVshR1mcOCgumK6RMk2TvFudLw6ws6DpmCDrYMrjCQIPswDjXL3MYB1HNaFS
pcvDfSwQop0YZhG/s2wUlWcNHM/FcsZZdhlFTw/Mbuhqt4Fjy0OiZbk0ckZAJTXBZue/ycu3BRk2
qP/vXzgDk2J7Ab5vwrLjVu1pfgOmXNvnkeJYJOMCSiliK8ixJIXaR6ixvrv2ediUd9OFQqlI5z6n
BOLEM2scr2astUbWo0PkvEsPSkblomphWPETBeX6Bk7hjzC1j9USLhG3x2obZOt1xzc6bg9qowcv
q0wKwyBA3TXfP7NH8LqfYnk3dj340BYyRYjnKiFpQxNuRf8Kbs0KcIrmZdNzbiPy+V/BNfsoF3Lw
RizWXRjyXlAiLHQPcQgfRfyF5lLrq1ehWDQV3Mr1tEdTlG80vd2IWNsgltUCm/S8RySfMzVLhJxh
7g57vF8Wk8ByPEp4pJihXSagoWrLCxx86OKmcRiJte4ckv9Ent8IbnTA/WW8eixLxqfrqZhOvg1o
zb3wvYQ6kIVbnRUa1kHHx5m5s3Nv+joX+6U93rOXZ5JjL1pjDzPnIfanGDuCGcGGMHWUXZI3pZ0l
pv1BiIpd6vTmH9vXQVE1SpcPPalI+EYnGCxibumvH1dHGGh2/156aDQIen5Ve41BeJjZ+qgDEqd3
RpF0SOvMn4IsAsozH69/ed9QufTUZsTdPrGJqFY5xCGyB1fFrJ7BfTfhgi+dRNPy/Vq3hjDU9SrV
FKm4FY/WXniOxoyXusiwHzC1xADKROev3wx0yFg1CtTtZPjdspPuwV525qHrxC3WsUqH+hZw6vFA
eCSsX+Seizavg8i29MNRc4xGN526TKSSCz6cHqyv+icbFrwsUoSiW2bNV+LxOUDigpJqzMh3GGQn
S6x4+j/9Gjzdjrsrj/kYy6ldpOkSVz7SOwspUnSz06JR+h/NZlAeLE2bWQaTRK30BGG/71RinxmO
MOatP0d+vOx6tJ1FY++Jh31Cy0ak047dBW/0UeKA2w8Qwri5ZkGqP5qEPruRVhBH0r9MjnktfESN
uOlwOd2bghaXKLvRmMER0/S8PP8+gEuK8IEtWBX802a1lrNl3rzcHGCsCEzP/hkjj8o+7uFEuWZs
qdBIzchWFQkJwWn/BmSjD1/36J/wmVqoAKAm7RQ7NoUCG6mTrKaYKCH9boQj8joNe9oJxg3WB0pi
ia4NrcF3on639Tvsxy+cC19tmJYDh67NHn9hZHHG9gxogGPtah7wQOGb15tXuD454OvcUEP5NUOj
vz7y1l6xM7OZnojc3cCSjgOn9VE7ubQJ8mqS5Ojr2MrT7Yolji6IQcNHBrxl1myVJeB/6pGjYljb
EW1BYdeWnnI4qzioEZwULM3g6bTllLTF0DHKkzhWFZKOreV9CdIPLhx0vexPZXk64+Nadtfmj9mr
tnxs9pfZ0l90vkfMSI/6+r4LCqPDG2tBYSrdaHi76tiFoYjh9PLUejeJN6MnFQioi7Tz1F87RFRG
uGLH0lmS6sg5+N3UQjHv51L373cvSXgYmGNw55EJE3FP8S9A1akzfRmccgqr3SUomZDFr/yilH5x
N/VRRCQpv8Dr3wkTnAWwa4EN0yUrgNCcqh2JYDBrtnsjkZKo6xPGHeQZmmSMdNdHRkw50suOiwEz
A2aBdQJSGJMp2dn+oXVWPOxAbAnuOA1fZuy8vMetHzsvRshrcV9jkAsbSOcABp0D2pELqQfQQlED
2MWdPnFCibRnRUklrJxmhLqNafLwqny69BAoUGISjKoUaTC/vguARN28kHjqaGPp9r7hzbBEJNZv
WKWhVXtDDxaHdUZkWTotlkqvY9OwYW2VNO3I5g336hz9RmCcGCL+vrXpj9ohJXPzAySE2x+1rR/i
7KzKa+geyJ8+jF82pg2jJzFXqvtwrqPbhOpa3VOvQ4akZ5z9UVFSuS1I+OtOOOLjSJNq+f3eFf31
udS1kccX0TXAjKFTOyY+Kp70M92LiKBC6OP5ndGhYzSiNWY5g05yEYWvaaWg1G+F+v2GRx1tLlpX
cduiKhseZHPuYRZU5Tf4DFVg1I6jF2+/NDBTaYvsK4HrNWF05/Mv8Z1Ca8YE3HNHMST1bSfAjsln
UduuERbAFNHtqQ/jhLCl21OxNT+lMXtRK38L/SS6ujPDMi+2qwt6BULnAVRqzv0AExBzIKfsoVBk
jCmNfuVQzXjYu9+qHZChc0n1XY8j0Ur0z0xpiqIlj3gRzk2/lqIIoNqBTA8yFuUNn4juuIXjN4XU
KzhT+ZDEUmJW0m2COxKTE9aCXVPvzjyyzWDpinoAo4E/TLGzPATlzyFfRB5iorxmJeEf1FN/sK3p
WEXMBpEBepdjCW9pyYqET7XddQ7+E672GOIBfaZ6+8+PRlBwLyaL58HEm/5w+T929LPIVpZV2ndp
LlFA6sGpAMD3S8OreirPySen6iOMA1IEDiAtvIyuUdC8NXfCsAhFf0zHmcrSxjUJluo4w2xmQryo
0trl2doUPwa2fZvW//zRxnKzXx3d6xd+qHWTPgOrbRuQnQC+90CojjyjNYkTz4ira4GGcUxylsD5
EWkTqeHdiFIR6Uvi4V+eyjbagOh+/YvM2XK49D3Z7fSx9Y96FpGE11EMJAgW//CRGr4XxF54n4uJ
TqAoHwanP54pRsXY1juSL6jFOzyVIjAHPPBdskAtZ8mb7jG9K1OcxXt1ZokWRDsVxNPOeO1DaXm2
CGAyYPpA8tFwi5XR8aKQFzIVjeRW6gbkq28rILxCcl/+bu+oz3MFRaS6meLtpRDrjcW/QRm8AJYW
XjLxSLkZduvrpWdp4Hjb7bnFPgBu5/aKf9keu9dCWDe30XspZ92nU1b695drNuF9j/rQ0lun+hV9
x+GDeAWw7d/VV+7lGxWzBp4+VpvQF6wliThcce/f0sLXiXt0fomdEejeeiccyxiPqutVg+KV0oVV
NoI+v8Qcwp4PCUa2LwgkJJg6YkfcgJjEnMHzj3tnl7TBjsLCL5/mBSxjqqM2k0z2UIPYy4xph/me
53NhT4VKrl+VfLLKFLBeRmmJ4ZOeMUXPsDXWuP9u633LI4tIceScLIVPjM5ps4Qve4x9EkldZv/U
H0rr/2PUoVB1g681O/vhRcpLs/DdG0ZPUvNn54t9U82HieWHclfCRBe7ty4FXxgnD7KlpO6PHkKT
9IYnXjqhKj8+TWz+m9Qwx1KKTNSMP0O7zgbFu0QT+WGUEN/WNjFbQRzXWJmEoad3dpWUJV2rnV8W
Gkz24dp+0rutpePo4655JXzuP47vsdFdLHUiiYqdiPElkuWx7tUvcAeCsBhawi/cjibeYSizTPI7
56yPJd4kZIiGrWiFnK7KVYp7q1lskTSHO7VqDwX+/lDe3Dseklo2MRxTgnQZ1+JJl/Ngy9PYWJGI
YzSIqlQ/mNjbQkOY3Gx+FliZuKOvbNN3g9LL63viPqX2/8nyuJMywx4z1ZhBr9M+lWGzlhHWfm3K
t8hLb32CBgtEK4efnR1UcPZohJXf9jBKnRH6WwlArHcmMZvQ7vz4tJYbNls6mXIU2KZUNv/Pm4ia
Q7+R+B9ZUwGiVDZL0c62YncxMSwwdQ8v6/FmATuf00YQ7d3wIWkfmhTsI2iQBeyxISr0OseFnJwm
cex+srg50wh/H2bUd+nts/if0X0oxmPh5L2ubfvJw37o+tQVF7psL9Wq/2AiidiIT5rw0docLSjw
gxNWL8mOOO/qO0QK41S7CHjNyrwQ1u68e4JJLEIoXc+spfOsx58RPvuA4GJwTK5EpL6cvt+cKwFU
7BUnjk9mFhS9Wkei+R97nqdp0SmjBoI78CxZKRONObymfTH8CqTF9CT9haOP25zBRS+5wgXXB9Ws
TYdJb+Ad9QbvfQOKNLyjtrqyK19qd10bg9pViX5BARVWuw2DDShNMsZ46YGbsysBosDKmc50smx3
3x00JqJ1JZkqenGYtXLPz+UPyQCVNkSL4fECbV0usQGySQ7YN3uBW2r+ZLClEnycDrKMrBj2ltk0
eminEF1/k2pMX7+SPNYZruCnJIWICbt7/nnUJh0yk6cVzO2qV6len4fDVAwU72WlPKjv+T+bDmSC
88Mamk/59pW8cfXaiJ11uluv7iJ42bAuTi/Y+hGUvWB6SQ9isG3jDpVryQXl453TX6xx8oPXnXGS
4u9KMRSzVYZjhkxv9zkFHpUpiPCyh9oyCW5UprXY/sA8/HrczeB20qO/6WpwHCEZ6oswB7kmQNTb
BI672V1wcTfx7xwJt3lMfQcdv5/EadpCpukRI37bpeSUzst1S+xIL36i1sXKmz0quJwZcMWIvnjM
ThaFOfV+rAUB2rJ/pep8Oafo9FHiSHDjBy+hvxGjuOGwT2UOAZlitB9ArylkjCqn8eTt/LEqiA1v
ctIihrePWK37gP28n6PE7UKU9vFUU0A9XRVAsYiWh0CAhliX5y3VAvTJwG3iRInVdoau7I8CMCx/
HMo9YfmcA5U1Qt1xvgxLnV7ZvyWuzXeH8r8mloUDOfwJlfNMFigPXtyDmax/SzfxVLIumGvZ33Vc
OY8cJqB4FMHhXBHFY9pWmaY79nGAP+t4xVjvrcCuCZeBIoyUW75qD2o3Tb4ae+n04EVc7jiIVsa8
IK2P45aTYBeKuEwB6Q4Jyk83/f1vM/NkoIsihTFief6psxkNfLsZMte72sMOnij/KYk6fpqCPEdQ
mSItjeXWriAQsQZPylJO+3OeEJ+oPXBy3Kg7iYvVoiFb0kxRXIKuyBzNaZBbfeJo76QaqTsGowh1
9S15HfR0326fZ0Z/VlAkyOL6RwUzdkOfI1RBBTLN3VrbFuwrcEkFrfBB1Ff4QARUhUi2dN/EJjCo
JReNkGZ6OPpRN4GCuDZRPHx22PS1My5j0jol9IYAgXahihpvjALoHPMx4DbHAlyhp5WHhjZn2P2F
uzV+Hp0313/oLPOnIoiuRaQkdaAo7bnHH9urqlrWFWQkYToAHHVUfNbT6vnQCvyNuSe6/LzNsZmh
oGfeD6eYc9I5FHwtT60hLE1xbpuoSBo/hwfjkeO/yTgk8fiBGCT1wylpygFQd6b4EAaVpQthHCNQ
yY9SIMXTZc2eqEzNxtmefD5saHNaVOIv0/hojfVrX7PFFNhh22L96oGamKTZRE/Fhl3H86x8j0eK
ZE5t+H/AYcxZIVkoKFIeuhuzQJtzX0UaYzOt44zlS24MleVbs6IPky7mO5v5CysKx4Qyst7vT7eg
4MnZ05E/TKvC5dxYHJ3XVTI5CXdPzX0KNwF8s3ZUJhtZyPyH3RlN3LvJARBl4va5zZcJ3e64K1kI
2eyjNaueOuKJCK0Mu4aO9jQoStSkVm7fcHcc7Xiur+Jxr0QkyPT1qhM7cTmExCcc7ipjBXNOpU3w
Vz7E/n2FNQj6Rfl3PdivAKZsu322WhPl65Wdc9nKFD4kT2r+7OgCqnUiLhd9k5tDyDTI/f+Sb68H
bX/JB3xzFc/BjCZcOARHZa6EzWdMXK7DUgPa1+KDYQUcStZs7hLbDztle9kpw8oDpRyKM7wYd9fk
lgWt7juJPDS3xZMoXmXpdg4znEICzkr/UxE7atuNp2FeM6XT4kcrC6vmxxSuOr23aqXon6Lqo9Kq
OOBDsNJrYWhsTpXXqkLSPBaisXE062E3jEwvfh9/7fpZ3Vd00H7vQtmW7kiVvntcVx2qJacV0Tq+
5q6IMvCSQ8N2t8LRdR9vvWmVrMBPAiY2aLv3Vas4ADq/r8sYH1h+3/3B9Yymyb9MRj8LPw+NPSkQ
k6gkQnklJaBdF1mp7MsodvJNnEsyGrHzy9gXW/PtlnUUIJe2ashbdtF4ZD53deStaOrFs9p6byBA
zpyRC0E6bILkkkAQ5/CA3ploIQG0KjQMEIVzwWGm3A3Y5q7k9/xR3NgtIMq90c7B5/6Bu64JE9LT
gh7pYXUFMJK5zSLD7UfEr8rClydQAoUqZGeNU/ie8/uNqJRjyOChOmmJha5eYv6ATA6JSIc3ZC3h
/ubK1B2Abm9YER7Ek/BfdTrm7ptavAaWLDwXfIayrlOBGYXeVNC2nlTWkZJIw3FtyqXYZYhsnnXU
Z9TGgq3puXxDg4kN43YMrRK/9UAXjV5CXNuZO6cvEPife/pYCiw+yKVH/ezM6rWkRvX2KYSZNe9e
UGldd2PxjindAqLWXU6LXDgklO93nuKThX3v6ubM6E3hgjVkVPHfAo07Tj4juQYBH29UC3iZikCQ
GsqZ2iatusrvqn+20OReS71FvJhgteqKwnpSq+uUwlsmBU/4gRU8mW16qp3zi920mgv7VeXn3Mbz
tic/FLAoU+BUVQVt9D25mZcDCPFOCNV7CgYmGJDRD2wDrO+FDa3mMDA6ispR3r2Pf2nw6i66sUQN
u/S6+R2Fs+FFLeu+LR3jayIWZbsNs1OFJNmEkHeNvZ/7q6MYNk3gO8hEa7LTOrjYn2/SeijWnR/w
Hu7zq/3IAaku5NSRbVhq3boBRTcHrlkPMNHr7915lc3kpqy8ju3KrQyASC8Y2fNogRiGsuqfHbM2
Wmex6zSWC6NWW4TfXH9gCH8pwp9yJOAl0fccVHsZuUT6Zv5vHof2YXRXuCY6uxNWCWaFTu4wOgdV
2iLltlFq2p/5W3diW0WYLdlO9lbN2FmnVZxe4Ky0eAPpTBym/o/Um6fiH3zJDATMGVLGbx+JndrE
IkA9YKU/QYriQ/caBKd6IrlzJW5dOgLgfA+1Mz5b/wwzAZMTP0jydlBCG2xrdwfbvoQhcvNO1U0W
xIzL7Z/zjK4kbWfhhI++yQICyzneLZ4F5RZtqzY4doF49fl700snFMR/zK6/b7HHWviUbPeWuLXF
kN/83K5ROlMZxQpC7OGeNc7uH66qTb1YsBqc381B5cTgtsNMBGubIR8gt0AAdo9t/wKfMcswbWR/
E/7k/tEhtHGvMvW8ul4CTEBnJxrZz2/q/xil857I/mCDoKalEsCm0dSeywEvyVyMGPrEsvvqN/fT
aMMPJZXsjp1j2zPDASM7JL/UFCVQxt+luwcbJRRarjo+vtpJgTNBaqC+bG7RCYntIyA3bkSEM1cn
LhLuFwM1UWmo996Ot5pSUp5jClEz/5AymC+jmSHZb8Vb7U5gb4VRGrbe/BYwE/ak/1JFZ8pWhBiF
01KpKeH4VjU5/bK7Idv9sdDEZKmS3jIddozseI5kXqvOlWwcbbVX14QexlDskBWZP+8K+1YTOEoc
nTTY0UlzqvlJ5jKwCuQsASnI9LfrRDiqhkKmsuDHIxcPwL2R3KQ9GAhq0pQ2hlkniEfyLzdKIEix
9CGOt8/hE+y+XKuXu0IYhMyNmUXJ68pj5D+4a0DP9zQZT/zAFT55w912SVI0a8RlE6P3qEOGLOsr
SXhzI2fl7DyC6cu8DEJztEKalb5614QzbxpilNiRgNACgarka3bWRn8vK0AjLgX4XhVs8tKYEXRh
00s7Hw0uxM0N6F828QGQ1k4AOgvZQ54vLJoBzaXi6wz9bVpgxiGo45PdpSDYpePI6DY8tH75ggRh
eMHPMhfpwymDNt+aoiC716nL61P0VnpfheqJK4sfuQ3mhW2AXBZWn2zf9TzUlUSRgXkHlaZ3+mi4
zhUv0Do9Z2QHTP1RSgf+WLmCWkPsT27po0otRwVvAONuf8KILPCJfD78/t14XOscIzF4Trg8OBAp
4oF/HQZOhC3sauNdgXmxqf07rL5ikgz/7I/K6zshYLEaTlmLTT7eRn279Hki+04AooD3H+pH/GcU
oXcllR1JoUO69AgnsMA/BjjGC4n5dwe81oeP2+k17ZUZLNK3UYr3YSrUo8uwNiEjSX44Pemfb0re
ubEMuwodRO9sPU6/oo7iQ39NB2Zub2lO8bLHzLmHnNnpKGHSgWlwociS8OIteIxwLsHM/O2y3wUD
C9QaTE+GYaC2pafjmCVbCzpvtq/6yy6q8b174DBELc9/vo61/gUEF1OQWJIOOqHp1H+RLx3QIi9G
UbukAkJtwLcL8CnGvZN36prfxQqZNy1LSgBJF+MH9cVi3PpzV/YKJ40l1CAAnp6xnVA1RQYnjAf8
bqkljcMzrQpuHUtGBypagJoLcZF6ogYJBpFgXjnRxliRKDjYooXgfOpV8xqR2zY9d8kguzysp/b+
0C/s4CyNfo6X9KI//1TLnOZeo1PvjykrukFEOThbjFqdRe1jvKBV0MQiZ/Wd0t1pL90O8BK9yWXx
XMhtCKvVwcgrtIGnBuAqW6JbwCpSBi+Y95SqARuai5x2I2b/Ne8PcA6cTth3DBHY+2WaZ60LifQK
oI0UznLlJYZouJ/vjM/kqVvpSlNi8Iz0ZFedTEVu5a0WY85hxrz67XAapUMqHQjraOreaoaAVeX6
iNV0G89bhIZAyw77Bnzthbra6q5c5RCsthIPRs5+QZEFFS91TdTjcbgHlRo11IuLFE34ABmRK+wH
Avoc4Mp4b0ixXmY76x5hNOpW6fdVHFzzdvH4Gu345HBHf/Op6X33YASyprQPWmwL7jD42/JB5G6a
+0hbg4XExwikamxo3a/ro8Y6ocZSIo/SAE9NZ2F0N5KWFanJS2CwdKoOdPDgXKLNR4gch4SMJdfO
oy+TD78xaL4Z0Dbn0G/gwOA2rW4FBR4Vocil8flFNqve4Jp3QJsiNSniv66muoajHZEL/GJbyvbS
+2R2gRotiAJ+XHPJHX0SVDOvoo4i+3IGPfw1yTC+qQglosh6UzIJ6CeTgJhMp90NkhROY/hz/n95
Tst3bKVXgcq4pZ95dbIjXQABu7BB1FP4IEjrP+jFkMaVXfiAfgILM7oYVuu/IzN3Zdg4UTpIN2RL
pQJD95Xh3omrgHNtDMOPnH1uAoGXo3JQKjcX4uInY05BVWeaglMU+UFFHFXfLaIBqkQF7CaMJLPM
p3pY9NYUg30rluwgzz8GRAGlvFf20+Vs0WPtzpzOIATlm+dEOnrWkZ5NZSaACaljZzIKT1qz2G2n
O9q1ljVDlrBvmJEx2tDXTrY51HAqSpfcrBYlkmUTID+6AYAYy7arfvBcXZFTDvX7jhyovryl7+Fi
ss1mbom50cP7SA5wZMDrkEYKDnbgSvxmgHFEZiVtOJz0tsijsRF+lE2JRXh3TcSH7ywcBaNQtYcA
aibaUOQGFgDG+qTs/KHz8OZG7/QZGs1Ml9TQN+vTKbezIt2FuuyTboY+cc/2bIC7gCNKfW+aavxN
wYLbaPVsFyW14jHmfYNOOClvv3sojpjj1B/Lbd39IvyK1jpT7TNR4/lB6uZyxWqXKGcY5g0zxrdl
43x8ZtN3tT9ldrP88tPkaRMoweqFzlE3ac6+82bR6GsR399cj7+6oSgqq9ZXXPcLeGU+B8lQr6wM
JvPXGox/GmSAyScFgvP9zn1dOlDP0jqG0a89z8TkjjbT44VrKcUdCcPmUFyj58cBvYqAD6eu5fsT
lqExs59vr3ZicmTnnWFSoj2hi9fvpb0Z6rTKQP/NrWeqhpWM/utrQ1q9bF7M915FtP4aYqX+ikhq
AEuMuhcOQTIcZd/VFcb5uamBAWqypKt3ZoZkluFMXU8w4Pk7falWL+zWZbVe4vPqc0iHU4yOiuuk
TWaFAemkztGnvNZaYO8kMAHv9Vyw0ebtJ7juIc4hrcbB+v3hnnBJDE8WICc+hFfqrzbGhsQaSsX/
VDsDzarB6+R3DzsQw7rghqYkwrXAF8enOwIZlk6ZfjfQBfPq7osCmpomon+icFZ7sWdfYTp67eH0
dBQxcJsY5HXmr1x0r/G6K/6AVxsnqiqEP1TbhJugpUV1uISNbMPfjVit91yFsbSPILuGKjWzJtnY
3KPAT58eEnaltV3Wzp1cy3Knr0kcYgS1+c7a6zw1AxcpicSzJU7ikIXXb8IVVGBb9LBpm7i1W71x
oq0PUh2QRZz4PG0r+rE5fIJHJMMSCGFo+ugYLJq+AX/Q+GzvC2zWygrke80pi0V9QeDYUDkgzmxd
6HYxgdvLbjTcMn8EkasQSq7gTKCJ8I6U+uowK7UYNrx/xrL/T/RHlcC9T4J0Mwm+ZxFlFOykLdjr
ugiVtdIF1WV60EioDzMOPj/ds8SxC9dPrs2RzAktP1EZjxfuleijVKXZnwJhs2Wd3LzH1PG5M+E6
oGXMfNXjKAusfxXQBdAMY0zHrvWq6cIK+MKC35XJoieB/QkB1Z008VnNH69FijTVtrDqe0nfxW+9
vmzQQ+tYFMCfUdlDUgRyLGNdaGUFY5NQ8+YKVej1nIPHsYU0NfBuRWl2ZuU8tPNfO+SXIvA1bTwb
r5UcxYtF7sHOmC4SKeGbNWDVbdF4fXubeo+eQ2R1eIihaSgP/mfZMFpFBuuOYGadkJtje7wZPNH2
jybBuZEU5NbYvyoZdslxNbUYzaHe7PEo2rPk/kphaRTyqDIQ2gySiWGjpIMKpvILzB64ltZWK1gY
0TDJpRC8u0ShSwzf41LLwwvxTMa9JfIDlC2m+8HoQJHzK2XScBsNcoH8wt05UXlhmxWGPAC/Ic3u
6PiUMIFJYX/k8x2jia4oAWHIy3gbdgp/S8H7+VUvsq0Ak/bv6ckQcRjbQeSr1xTo426HgtcOOurc
IdxWS/gX1/Gti7ReLVkoo3+7A/aNeYRqJ9DnZgAQA9RQnGhEPgJnoB2FsLCle7VptABsYOnbD5AB
VeA+9DalaeAYQTuNZ0qXOXhkBlQp4NuaC2M5k6Ug50GkhoLPOkiNlLvI/BZ0WTdlXgvgCL2r/zFi
W32jY3qUIyoMf9ZneQZhxs8RS8HbmsowuOn92SxBlYOib6td9i/NAO+wQ8uyF6X8FyWZ9NeDc3Of
lg4lRfdEcaWGU4c0xvuCRnKB/miIr6JiMMbtTBBhlvpUM7UlEN925DwBVKzSLLlaY51viJWepD1/
cwcXbKBI7GDeoqBA+b+6JldMhkOPgfj34vcY6MkmsDBFXSTa7HHN2Z/6ztVfb9JVAroKdohbDW5V
M/Mh6GFT2myvodUJky0SHesJFFSDo7+16pQXM6P5Ar2jxVz5y6AkQ9X/O4BFn6eX1SR/Vw4Ucpi1
oyCsEYFDlcl5tk+1po9gMdQSTraPR/lp+k8WfIWz9qumRa7nzLbr0g7BYBxyoEz3pIgilHfU9gDq
HgBOuOCUML7hXCZVKXvVr8n3Rb1GTWKKM0iBaRD4pUfeZ71ebOPnDqEsFUInuArqWmfQPo3BKP9p
BhA0hmXroO+Yuglt+mdBWGyTEmwfHJMCBl2yW2bl1hB3TryJj3rDv/FCXtL8NOA2eKmShuw4ZphQ
4OShDDACAGbN1tbn9XGICsMtb18Kma58Aocos9Vi2TIwHSEWPzrjkDXmgZZo4Avhu30KpQ/vxp3F
KOh0ZAXEqASW1UBBfNl312Dp4p/LZUkUp6D39LFXTc6gerMMnmc/z8cqfwhfWC/fmVW4OWrgvKZZ
qxgDj0+7+LhgW3v5BgvCQPfDyUmvZibp1G+qzn14DH2fEo3oScD5q7m+tJd9Zu3rrWh+5WQ6CC8l
yoZm1RQ5b6CM3oivA6cTJ+Y2h/hWTjcp8grxmKgyv+oy0cwHFpvrRrDotHYnjyvsXkfTf4BpBuZt
eT5TUk8/MI456bTGWmjigyHIuCwglLBebwFe+5wDzk6tPo6mpVpKEWIhH+d54rqfsGvrN7/VaWvI
zELeFBK7fbkGeJ347ZPv0z1ZU4iOkO6S0dLh3tPX8JIP9Ffh4OxOPJTKFLS1hbQ3uCJXzHbzUMUq
0MmpQi0PT4S1wQSNY3M/srkBtFRgiO8HFx70nHuTHbemMYpcWaNRtt/fya7wNotbb35o3RCpDEEI
GnoMNTbfba9Mv5sOCObNbjd5vNQwM5qVVJZpIt+y8U/iKq66JYAN4V6X67yVfAM+lB581QWZ9S/c
sUHgrPlRRio0Lu7EsP27AcqR1CRyJEr6HB20Gn2D1ql/aliHesEN8jzWNA3sgSbb+nV+dZRtE9Fi
2YwI8H3rah8aIzqbXtErvcJf/cxDZpyNz9pp2oKswJUe+f1f7cgNLIgS8GkjfYvK2vprDOTXWyxb
Penlh7RpL43huQwd4JYBAna2na4mB4WFdRAGZ11k4j8WpYiIVz5PNR8PxxHXwBA/fZBpE2W0tOGI
FE+uF0aVyVIWrmthdkv2gvUKCPpRqjYpp4blH0UTYWW6y9C/XgHF7ZFa1f4Rt6y0O2aaPYnCmVNF
0iE3DBAN8tEmJtxllcccKcMWZqIHEcmruyMC6wJMKm7Lvjr/PYbeufcOxjCHzzpp+sm5GiUNEODJ
cvla14cSqm4B5tIilwCoBVZfk8+FwkGyzrC5U4EWONGpEmKBsl0zuMfRK5kzFbpahlBwfod4NFRt
2fJiFTl69ZUeCi+DNJ5jidiWunOTH+9evwPQULzHWuq/MOs12C6mgWzMEetG5DQV4suV+szJflJL
2jC/lVHHY9+WbhjbX+ikFL72FaZfRizQPQ6vviDuaRVwmvbyV7Z1wmCxoZZzh+UmIwTL2q4KuEo8
80YLs5+GwRIK/+bqG04MTvxBj0tRbT3CPiX0cYLLMHn1YA5IeXjNjzxslzyoD7PmLg92xaOX4qMl
QiA/POY79odGiCcpvHv4NkHXoQ977VgF0ji3TZgMiO0W5SiLccFFG//cZSRf/hi5QbLfUgmy8Vz8
3TlYT3JcqMIWBmrfWaxd6HLa871jNF89upmxzACMcTA54DZyrc5V5OD6jUhEYln6RMdCci9VN1Fg
KtKTYvZDZU/dzinnQbjcntZTuwEWYtocjU0yYxfQkhoGE0Iw3+maTW12VtDfX6o3sgbuKKD23gZJ
kWRNtQOFXeJJbwcPQinjWugLHRFhnpE1KRkKuAqoN9e6D1tXbNZm4DFj0Seg1L+SclnjlFyFHpuN
zlIS4xWoq/D0yCOxhik7RyQPvaoT8MX9C0cDxjgLhB75w9CPShFXKAKfe2fayzagRNSSHGbjP2tO
kJkR24psx7jYBgkPHyHNq2b7HNrhlbTGQCeQO30Mliu9kVcd3xWG0cahMvDXF68u0qGa6NeUNXzU
Ktman0qUKwhs+z7Bbgb3UZv7EHZP4z6lF54H57OxE6LcXzvS0N9HODeE9FlugPIOfTwWYEcG02bC
ACsZKiorwCtFwx7+/yyuabbK0edHKVctE4FUtafHw1wi9ErxCPBhIrZAiYImn1mByyPF4Ct1p7Xg
tz84c9g0TDAP/4RVd7SFYuoG9cTvrHo+lNVioRMn05sPs7HWpHDoqHXo0fE2HFgcALVMeFM3Is6j
U0ddiT0o3LAQOoVpH5gUuJQuFOCernK10VjSg1qFQybJhJiaXfrxEFzU65L9l+WfelKPybqB9Xm4
NtA0DtRWoVxr6uWpZ9NoUyplUlDXUnRIIbzL94I8bD0xDPM4Hz9B1l9YPA6sbMBifzNEKVmowZPp
6Wj6AysiSBj+FK7QfnIgW+GuORl/DZRTQ7gJ2wjihOOhcCZxaZQ76uXaqTshcheNRuTv19avUVZi
2Bw2nQf7l/g4yasrwEbNQ4cLDXPLi0mieYkdpLU4lvyRwWq5UDWwLZOza3zlTcoEy2wQknY0I2Vd
WmLYtHJkjIYv2IBHOg5Z4lqtCjzr7vIpc8K2qyzAFeOXIe5A+RpnKKSiO78ENJEb1pjMLuS21HSk
2wGOIVOotsCLa4aoaUXoNS8nC/yjmpIwfxYd1ktw7yYnGCRWut9scoFacejodov2etl/uq9qcNAz
Kc0KBgzwA31SvAkjKUyccJcPz0FK1e3s6nEQhjTdypMH32kPGqowttAwgqjngv9Mk0klsnFMCSzc
haIvJTJF6vOQUtIoq7w5Rx3h+dE+Lkqw49phnvcnY6nnVsU3PNKMDIc9hcE15GJm1zBCd+qw2V7V
yL+uZQICXoaIFcCUnfZWleuhe9eKULtWFSn4uMLVmyGOCBZnAhQL1HyUVY8LYNkT47PUl4vlLGWS
L98i+sOzOpwmZJ4g8GXm4OZ+qBKqWezOB6WELBXSeRFJBJc+11qbnCvSDICAKVr1eqnHOvQAzpLh
CRliRUkq9DaOgPsjA2yJzf7bqTs1hKcEsX9dOEVbpCvnMRxg41xJndew0driqdjDFL0JKoBciDkY
GEMG7HgWmcmU2bKy1y+rzbdQbZi9A45MTpVkEu1XExZ1IP6a98OySCufb2QSxousZUilL/rz4WeM
IRoA/GAfIBBF/O2wnjQnn7agzpLmOTT3uDgpVLyqLZlZNty0qptOF0Tp1HEeIP5UhlO2FYuuIjGg
XmoNg2uwQToZ8QQt3JoYHXXStXTk5q52OHXoiOvxPsZCVEdLUZ3pA1vzLQLPURiApB8uNkRm0Cse
SZUpm3mNpiPnZ8rZvanLVwcEzUt+L76NLyhunRpdI2s//Jjj7d6eRBo0uGGeZSFXFxTQ07/tLtVO
whCrG/BIhcBiKI5p5Js+YrTfeiNYHU2ch8Te6WHwiIh6krXyoKEeDsCV8FbhgA9onnpRHAQgDnsk
rDzVnN5L6BXArZJIr4iG+NN7MJG/PpWKqiM9xy9SMZgeXM2nwOlW34ND3HrAaFvohGsbY2lkCqKH
7LCX7iXvZY943C5xLjMNM74KSCyxf2e+IyBipNpRheakdlbnaSRoDxxwvt1bJ4SuTdjQbU/0PH71
chmLeuQUYZPBIRBOFi97g9Zymds7iJiZFJ335XiCZ/d4NfUbJVYW0dsOEsAQfL7b7V+h1QpmuCeD
uR27hreAgPQs9C3nOQi4jcoW/kWlneifyWwDbyBpsHHOhiwI3yPNNsGb5C2Y8uN8aE/4UJ01kX2y
NifBJg5AtQoH+KdhuJHvDSVrJQK5I10WVjz3Tt+sZGEkPn9fCiycvVfTVfMK+9uAior5pHUDL2oy
nS1X08S+M+DxTTXmOFWVHwmcBD8PXFTY3BMgYGlz9ZyXCY5y8tqb87etd/4se3jHNxTHesFXZjyr
49UgTm9C7Z8q2ojn/QrZ4RytvHK7OdVGdwAibB691R5sttjOTPbQdU+8xwAOgAM3md/p8SGkKr6F
wfSzKuMTmTe+lDB72cxUZYJ+otFRYV3IPZ50Tx6n+cx9X5hv4vkxIpw67bTXVA+sGfI7zRohiR12
4EixcKaFa7DOhsEYjEIxOh6tPhl+zS/n1i7NEMbhPhfNQaHkSREmE1qI0hZwyeOrNCC6KKmxTlnV
6JU0+LCkzzas3dVwHt+86MUJBbZkuCB1vwHZTLy5YfuULiyUuEFCa2fDa5paKyuVRjLMc/dj7wd9
UfSDS8hc+ZFAW76fSg39ywY95yajixzXQ06JD8UFf8kuqfBM1b51Acl70iGqanbXuHrm+0kuyhzm
euoxmbbuml8FJgqYSZtZPdzVnG8/nETDrJfu270tuCeZBsAd0qV4zC1C5z8zwsdRLPCPn5VyNOjH
Ulg7N9TZ/jaKOZQV/QxkST9Wg/dcwTCv8gveDMZxy8puPoZbA4QZCnUryoSVIYRmJRFPbH5CIWqg
UwFSHAse8cVQUWWXXonWOfZZ1gvVjNOuZUyRg9d6Aq3R19bwuhPZmPVfa5KbrQjRa3I6wq2a4CGm
A3tSVxhy3SHh5TnhUIdS6Q3xsDbIK4JOrDGLLj/n7GcXAOP1cvrFF5SpJXv2yPQ2EiuldNnU9pr2
DCsdETVqXxy8DGX4B/5yjhfPGXSD28Zl3EOVFKCIDKX4dP/U5kHBGpnnIDhWQ8hX8SPi51nZyktA
BkmzpGHzEI4aVN20kVjxzAmP/RVicAf+Y3Ao7Xx6ya6hJiJ4P8f5mmplJgyfYgmdKXacIYhEouN2
aJJxPIbZ93NFoMD8pd2tm/2bvylUpzguagThu5oGeCuaOSqP8xCNJNajoRbM1TetsfTE5WR82Wn9
X1ea2lWvX5wPKlBt0khAdiPWUHKGs1pF6WZrww3G52H3ZOQbn6Z11L/K0/UYChEKJPnJ9IftMBwB
7pqoe3fJqLctCOKXgwh8LDcJrfb5gyd+C2kqEM/RQLvQtEXv6iLYq+aFbyXT/0aiI/NAoXsXtktl
o7SZ6/ZvZDrs/7HGSA4Ib/l9jw5BVbIwvOaXhRsJ6W6zXN0WauqwSSZ9hvYzGykfEIc9pI/0Y+eF
l9vOxGzkj88/dsNOITsr8qe9jcmvVqE855tJwqL3Jpmx0RjPGR/9POY6Ug2MPlCiBIXs/nE5VLZO
//4PYQFv1qAf4cM4ZlCoFHtYXLYm82/Qemx/CuL6W1cHA28wIOAKgwoBF7gBEzg+sp0fV6QpUXEc
DK7KCy3qL3RnL5HixyVUqGBhGBPIJa7+W03dqfiu9AYqdxH5Mpu7zn0K/nXkbSC+SbYc/NoXHhJk
yh8CNKVvxNsKtA2bemes72oxeBN+lQci1nMRxPRTBwwIKm0IXfGLu8VUtJhdwHAJYu26W0/KdZNM
mqXNXokkxySWDnGcM6AwaUNy05WrlwJ1oNBBrgFqUkg1N+rF0W10FroDdnEOsyins3YodJxiEDvI
Z9iMR4GmCzKL2DL33KgIaJm8FI4AtHTM7O3FjOqISlsC760s53HycAlIu4aVaZmS1KW9eA8vAX2g
OnwiKpX17QNUq6HQRgeBFr3GZWirKNZc2e0HxNc+4uhTEChyD83Lo4z8FZ8q7M9ooAd1zX2v6FQu
giq2IjNjW5fO/1/SfpqZtrGD03tMexpERUtLPF0O0zY+KhMpJqIe/nfwd862+LGJPrAv9ArNCoYD
GbA4w7tmDctjCvZa1NXobn1eF2tzX5lp6cMgykMLmJOJkN2/ueViozgKzsCGICkSnH3ujc/q4EiQ
Duu7dWyftgogn9h7RIoo4z3S1ysgg5jvQ6uoiZ04IC3NhZTmN32KuC6TRxWL7AxxDnrGPQ3M2XhW
rhPCx0cI1/eKqfVUOEYzDEGgSR/h9jxVNs1RpFJ55aJtxn6ws6lDQpf7fl8mQ6uc54UX21043J8j
X7Lwv5mo4Mv8hPudMH43665gfTsgD6NfeTHNrSr/yjv884gfPf9JpbdnZw9LEhgDuD9jkmBe91LC
vRn9kkVYVji4gk6voKOm0S39MUudbyCly23IAZ4TexgU37gL/a0GwAHVIvQlbAQ0YdDvk8PdaJJR
MfOyByY9Fyin3aiNzV+qvrkP7pKXPk8HdRbmjmuJel4wh4n4vKWCE4DZCov+yXGzdTOf0+zHt/8x
H55Lvgb/F2yo1kA0/rngtvWW4zhMzP7/1+Ibe+wjVJsqIC8c562r3FI6Se888/exVEMAkmOleH/A
dpdTfx4GWupDS7D1IY3f2AJkpUmdYwut7XPL1Y/LemugeoNlkmCCo1xavDgWb7B0f1daoQVolPKf
3pXhfHg6175AJYZ7EiAucwoFR+U3FvqT9pRN/aYQ//q+a/Hii3C5Uiyx84ffnufHK4jPkuYEZIhm
DvXlcz40oxA9l2ppHyzKGKIh0/b9wGitsMSDtZ1oyc69feHWsHfDc3kl0ox+C9Lc2k+5I6Gi3h6u
FYals+o3lQ9CFyND1V8142OgTtFsf374TpJ4D0UT9fL38nN6nnBaNNxqtBRC+vqRaN4y8xKbA8U5
s5xJhz5MuM6N5v0kNrZHnkPXCdb6eh+6sDOZ+eJrAXKCTAbQrzqkCm1xHhNbRjoLGMBZe9kQASWP
ZtBYSY1/BARWWu5s952DameTvQ4rtL/DCIaN59bcMOVHH/6HQy6u9tTCtaaCv5o0H5P9DyCbluml
+ev4qw1K3wdcgusmYxUD4f0G8QuxZkkWhI/KS8hjB593I0wy23+Joe3NanGQysFonCdJ8rJf8N0F
pjzAUTVKt/cGg72jpPbETsGDXe0TC/ZF5pP0LoamI8VB8r4DS6EnlHFQuIZvfFawKLcamo+n6eZm
2Xs8ejXAQf757NhgrLlbQ9CB8N0iaYhk+x7EDq/QhMldkDbY2vS33+dVeJyMM9qd29eeEXcoG9rM
tValM0/QD2Py8ho+C1YyGYL9WIjdy9ooQ5nLyZoUQ8LStaLsXjeVioVTRp5xyUvpdBaSPuHTdoGF
OHJLycdVlbArgVGoo11gRjpq+7bM23VFQ01rPMIPdXoj2ttVwJWE+kl3qRlIlfEyVsePtDIclRIq
hX8wQtQrnb8gZobafPQOp8AqOKV+lC2bDogwbQDHwUHljUlwF80fkovyGLazc8tFIhBeV4dH4qsE
iz0clURH7p+RQeqjXUHdX+aW8E83+iabAwImLrAsiHac7kWgM2O/VIAtoyXyw7SLGxXuptus1AU3
tRiKuBXGZGs+j/ajtXgYE9B2SIkzRG6Lsg/oUMVkCgOIUi7CaBxEfzTyhxlRwJXWPaBthhaeQ9B0
k6CPZgTbKgtNyqWny4WZEhl79+tftibwCvA4P1ZFdLllXzWRJgLjsUjv8aRDks0FRBkW7c0PCIF9
rTYD6YJsqPMHxfwXemDPIsy+lEwViPRRasDQJwWflSd+8LqScfIAFUu03LrqlhdrHB1nDvrph8Tt
S0asiKkV5oD/VXqEDz6OMUU68QE19ppYgS+nBKvqafQ3T9BWpz+VgHHq/jTACeUvjZH+PbsyFlCI
nhS9vq83B4MjDDc6YFWmgVQadb8pseJeZkZPxnRYBhu6JCNiWVuISgPouvNI4hHSYaXJG7uCvz2C
c4+BrhDrFm2fvsAWCR7ZaZ1SxVGn+J61+uR8O3Yi/A43DSH+0O1EymzCVX3ipBiSXIF7bD+SctdA
xrQk6zLx0WQKVFAn88pho4wugTXDPZfEp48z5o7JHJ+xFFNIfHXnR2TXFqSgCp/EbpmJ5vwbz48q
8KkXoARUSvKvjjDCVNP5JRL9Rax3rJ1+ApoXInZ7nOqu43OcHmZYob2ahN1r9xQPnOrWQ5BqXpx0
sdPxRiJB+60vLoDJ3zju9hvOWtNzheT/f46SieXsfKD/+prXfHI/1OnTqLM8isZ/2FcbCGsAXmxb
QUPU3tjS/6vCvucEDBo6GdVRg4s5PiDGJddoEjEF1OBGtKD0Nr78yP2swloxtScW7fHCgknoN2Q+
tjWVeS8MsLBTJJEG8GgRXm0MCWkF9tEgeCULGki3GLenNPH0nvN2BHfuJ4za2/LWqEHos7ZhPpw8
DWtlsEb2xCvPVnPE78wYTpbwOF4z5CGsI70fDS4KhHSUrleoygXv7S578Agc60wsvminMKZOmsGF
dCwdzemV735y92amshOg54CDGXuEhxTJttRP6+CuFKyCCnNFQFmc8q+nfhhTcWUZ6AyBmhAL25/H
/WugC9aDbkcIYA6WlVOahNk43TQaV1PX2BtQ2f6MyHyk5E5SdXFf8FeCUpzW6U4CHGZVW8kadBpD
XAlXo510YgqKOYwjp6+pvShn0aWANjCaD/eZ560dc9HiZYYA4ObiKLj6hjXx+IuowOxWd8GlfLuj
3RINetL5WdSGj0nqTOPkEFCbjRpPKQIeX3JJXOS1tEh5nTdesDrfqXn8L4EXWYlAR//SXifJI2vU
1SLQgo9fatUPEW4bG2YGVkWtopaYEB8N0CT2SJDHrxQKfXtM84wDr9JzKBrfji0V6xn2LVA/HxZG
NAPjIQP34ER5UCN2fYLMf8hcXFxxMwmP6EgvAdU0nDlKdKknaykAWDq0U1/0TYw//A/d8w13v7nQ
iA4tvOk38pqsl8Fo91CBx3Fi35LoNEBdE4LhAVMBjfQ1uZ7ApP3QNLopU6H//hFsiIv/sc+4MzWE
IJUygmwFfF/C7TuznHNPlv496keG8xssT2k799Jhl8SGxPATCH11rhtWOW4NSc2KWwd5vIo2NIC3
HV6dLzRvwS/4ogG23yAEQz2z7wDlHEzfQ0dtihXupR0j2eU2rR27sUkHqRXZkgDl2lmDs/1YeyvS
q0ZoJzLcAf7Atus40i3ttkilTyfv0IiB8ZiwzxZLF7+LxQj4F4/3MOumhYbw9RLfbfJXw4DImTdP
Am/ykgCTA++3G2qMPUhtQGWxh/FFDNy+DUiR5TSNpm3gF944ZYgQPmbWouadrMFU+MWSZx/NziBO
jcu0Je1DSgzn+oL6TKFQ7TB9MYNHqm4S0+3f5OXHpAw/dZbBOiqk95SiLBqIO8F3OzerOQNWNL7m
ObCcvZKpLNgtoTVuxIo76R4u8XYmXy3t/OCCf2udPdhBVy8JZw2J54avzbo9oNVevfTW4ZQljkIv
5aDGbKSqobmXcEGb64G9dPlwXyAHQ1FIHkWWeElgSQRWnXfyXziKxMPdR1mH9RbFzwnzsAImlL6U
4G2Lae0ZEzhjCxffmLMvvWkutfgJHpBGmlHB/anm+im+LrMKG2m363IOKPV3Cx4m15U4fFYN3d1f
7ur5Z60y9y6N6kq5jJFbeGK7GXFG8brZiqHZCdylOGEJdyZ8QTSlfbAc8COxSexW23v+0wVunMLm
UaykWrg1EIbFFPqpnxjv+4xEHFNeThu2ujpTS72/QFr9vCqrEgsUfxP0XaM3jukVH5fly+WcMHCM
AIM6CD5jPqWo3te840KZQqqj6Wwz+P1yxv1nNz9tgV3Rvppf/BAUZUGPfOpE3AJMxh1YQQwQ8q7/
h9HHG8rYNJs3SC6LONg9p10TD2SrN3gbCzRZgfnJbWVHM14e92p8Hei6EqkiE21T51J/7NURG81T
5snqlRo3BgIa2xBJHHQM1G0yQuFYsUzgeXlHPnQ7vldI6eBGtGmnF9xYwBmLh/z6og9vYkZF0twl
C5yc4Tqx9UimNzOqk5yqMUgffidTK5tFkRUMR9qKhi0ynxXZVTeGExJDo8K/pDgTX44bTD15mCph
620qNI4wR0rypXnkSqfDlrneefJ8+09BqxkAsP5AK/YvNRLauhYqazUTRly0kXxq5kjzv2eFZFWQ
FstyE5rLq+uIDxN2HhQqzXtkr2kdjXgNQqiobSgx1RI5WN6wFTPLSBgVX6387sJbzT5LiimeoKsx
M7h9vnWNhaoSEEP+iKZGPYchR/trNHoUk53hK2uXhx//03ZAHM7zovmSW4caF0Ulb0CwfwIgjK0G
oRIsaA8dNC6LTpKIXu6E3kBsBMPmz6offdI+sWGffrRUtzQp1f92rz8mysgVI7a0twdrsXKpXMGC
VyQmDqObWFLgTwrOMFIdK/kwp62HiTnvTzbzGZhZ+fTNel8ucF4f2q7FXy2E6e4saknT7MOEVIrB
ubpXTU7JVywh2/o9ia7Xue9rnq4P9GFby1MP5tyGLieATz3YTmIo0z+hlPOzzV6irEp+s/NEL0j/
eMsLZRaVFMFOvKn869rgWKQeOk5o5iUU7fsYc3mtv1KWcpoeSmvkCn5X8Wh90viH9I97TUhFUJ4y
ro8Ud5YkyfWlfcOmOwfja4z1blTN5dBWefPNmS93lpm7NN2eALnVpVqOi1qzXX/d1ZRJrO36QcY6
U8L9Vhh4zAZqbU7LBhGiHvI+Gi6/cThQOAcjseyNsBCp12KrLlzzJu2OhwdEEsWUoCXT7l83ZksN
h52mFA8IFilBsG0+U6Li6t8S6ryzVb0rc4e4471XVl8V3BjjNNCfjzEIc0Fp0Rz3wlwRDD01pC/k
P+mlfQBS55B1qexkc7IiKMtpHOhO+7ARZ218wa2+YQJKl7qQlAaXoddJ5NpzVfBLKjUz+8YX+iZs
sLpHluZ0TliQ+o4EOiTQunb+O2dvbVcPPvVFfShQBygPeoL+bACPAjH+AWTSZ07uOBoriVKDWmqM
AroJuc+D7GejCvGa5Ccx5WJO4pakEmhRs8/zTxBKcRBt1MD+7m3iMPDdSKoGf83by5+H2P1/adj3
RntTSO5ZKcZmWHXtCAbSAX4iDjZhdknxpKO526tYu/ZwSbrVPk6CCyqxqoFihirDM4bRPx/edG+P
VWOFON1xzs7xbvSPe21fTW6uy+YCsu2hsNkBAa1EJPLkOpIevXlCxK/d5R9+ABqkgOa6y3QvbVrD
iRGZtfC5HZiMnJcegyNzPaNUExB+opBoAesHfgaObdYxHRh9aLrRKwCO9tNOgoAucGSmITpjZTBh
QIaF80Du4JYtxXLxYOD0ucYft0Q+OdKF6tWvZxDIntlzuLLjS/s7RnnqnmT75jkrbpA+AmU2b+Wa
HMn+LDW2bqenj9Se+EhkbQNoYT5zjH3Nz/pkDFGf8gN+1/nA7v0huRBxU7LkuXTfeNZkWzqUF/vh
qHUlUNy/uoxR4ugz/CaNt3YUzXpZyucKwzzB1X5w43s6AsENfPX4NZwynCc75iLaFNWyWAuIReEY
6YZjOQc11phw41YZYUPL7Lsm/fDEovcj6lWL3jRI0vfwJd/AP5QDJP1gQ3pkEGhKm5j5F/4F1VbF
QThLRxYjqrwpBHBGv2hu4veZGfEGn7AscvPwIODa4XJ6PhmLXhdeGBeZ9QCJZQfYTdXMiMEOAIuJ
d05Cp5JS20ZfH+EGZ/rQHX8hBPtp5xcfY9dBPXmeRX1wDB7sPqifYRDKQXNRNnSMkrw3tzgxXn46
DevsKn9o600ZwCfXhRus6eyjFt4xo62ZJguRa/JD/qi3c5bi7BvmqHJlE2bq/b1/IeitbT9yB1g0
84KFLiGOkJQiNxPxDUv6pNIOI5+VKU0WCsI4gN9pXd1CdRpRjc5BRzefqbYiIrN1lH3O3A/9ruNS
cHOOfKm/xJ0XGMCo66fYwoKPgSJVC3Xjm2cFSJn2LQiQw11o9gV2rQD0Iv8kVVTovQbLOdE7OYPV
+/OZ4ZP53M2rU5Snrnn3fQy5qEeKyigmzgC2yFmICznlEcw6R4Fr+3LDWm01uRxMJJOnB80hYanb
1K+g9U/vNc1lb5pxRkd6r2O41c4dUCfLh6eYyLGxJDEUlsYOTR39CNbE6TwmCNGb5UZ1FL3hvcWu
IZ/Kaxl5KGnvAyCi7EMwRRPKnuG3ZOOclqmkzxqgtHA7bCrOgCxhm7QZ/SDUzR0Ubmlzw+zK4DKR
2xXcvSATsyWapF76C7yhPZTJLZrmjc4pfUowvv3GZh5vltrB2+ea/rsuvz2a3jQYFF8WnRc4kfNv
yMPpykLABO6qnYNfp2o11WCdcD7VVrRFodNSv53jyhpbzU7twyd9bGM9YV/WCp8j4KOu92XDPYDe
NHdZyudGU8wabVxUaRmm+rWIdI5OGSoZxFKkNRk/ZnN4O08dFBp0V749huNU5yP0mnR1aBqLFYyB
KvmkVkHfeEc3rEcvzzNwSf3kMhvUFPsce2KzyfNUdcD5FfD0p/epYojP9tm1rN+KHMxooKX/dT8V
5ThSjV/KlZKh+4bhCURN25DJwHJGXXmMAj3MlWkxq8VqDLCq81U8e6J3v/ikXfzcY/6KLDMjONXz
FOumCAITo07RmaTHXcUqIihBmmUem+0KLQWTfutJ+mme401QGUDaOZIn+4dXa69u+c1tB/GvP5z6
LN82Bp4gd5cPD5w+os7pW2ulznlz8gDeVC3SekLgtJcGKUyaOeIKVWxJUbsq2R5OkT6goifILFvi
YpFc2XJaiRk9KrycosRWLKCUxxonvxlEp118IEQ8AFeYNyHowWst3zpCXIBS9ff7wsV2xABMiSNf
a/AogI1Z5jaE+n+J3zV6ku/cIJyHN4FvPg8Ck4hd8gbZVGESejuJ2KlGzSyaRS+TrxB7Qy72WCNA
aihQs/1qGtePXCD2Cgcmlaiiuj/zmrOKlt5c0wDag+ytev71hzEqhoPfoRmL43yPSTAv/nuv6jlD
VVMKa7qpMy/2knBLyhVmd9/x1RFdSGXmzDzxvBlwZ/J8sJcL0Puk5YSbAqxASmHmCZUV2SshOLog
yvHJMH/UeeIYFHkh5Kxj5/QT4QCXyfoLv9JAjyxKIgnBAXTLLOqrd1pRYg0VWY+sQIR1aM/EWeKG
WeV50FwBrep1YISizeatUF7D3qnJuyag74gzFjxB1cfXmfjQUHmbfp3TMjwfPQkBkH1VqsscS1Zh
88PKNz2a8Le6aZepDrVE9lU2SWCKxC5Xsg0dkC48eG6vE9Osf0WxDFQWuvVqAGFX1u0PvZrXdOuY
hzQSVwHlAezZRMcYWsSD773CQLjHfGNa6YfAJRjx50H81GYE3gGBXSzwTu0oDUPn6tMQ0qPyExYs
ffOTJE7A2bKybLscn0o8wy5ce89N1KBxPJjqeNz9ceRPTLCH2jpEHkoxlfpSxcFEQQvmoDtsIMjA
fJeYIDHCHIzV/v4foAJGKSwt69R9WWiAuHQ2CGfq7reKalF7WZB8bhTxkNuZ27I8cNBrsAEPKwwI
Z1jUtC1WKbXnZL2xaR+VnXQUFReWyRwFhYSI15BZuzr6vJR/jjBRVKA9eOuOSDAvyKD7bhxwnsxe
CL46a5vI/TTU3lvcfXLyW4TQaQqghr5AWR+xXRWsmszcln+7GVZzmnZ7fUJP2GJoQQZxMva43G8U
I6lwqxUvFqslawUYtjrH8pxjyiqYO4dvCOndtUV5eRvUQioxvgEaFbFCfhPqM/4vKQ+RVPRZsTfV
1TNEaiTdLrXDfNnqlcjI2wmlqFF5/qRZCI1yAH9u7/ouzqLwy6j4RZZea3CdsbBFT+A1D8o/DAob
GNQ2lawQNaeQmYweT/guBEDCpOSFWwgE1H0COMHnJ6+5hxpr/thGYFuYqVzmq0YtjB0Vj+BvlbzE
X9afHV6VF7XZahurIdZZXb3anUZWTeBRb8GZpX9jGyVQzvwU8XhLjGmYbNFZtvoObrYbZDMS+oBf
+BUG6YTc9zA06nNCqDhY3GgPbi4QRoT0wDfQ57fBMnj0QITHJvPZOcerATQ46BVTQfKEUrviOE7Y
IRt652VXsI7kOyrwMCf96G2ekk+PZTqCWDFmrAvVt76w4TQ2yQ2t/QQ6f/B7LcPG0I2YeiQmjGyz
niG/pPby5w6PfFuPvhGwQHpEvyenPs1bU6AevlpupCoO3aWaN4tqiBoItHPDWcqGnuGsjM6ITA36
Skzca3MwapxMB3FgsRwhrSVnM8mV+YMRmbZ+Ck5FXyOm4U0q5bHmfXI5XhqkgVReONk+ia01pewl
UWjVMo7zaemQYLbhwmhbB3ZDvLvprbppwdor+2mOfqZl8ihLDuafVrLU3UeY95TZ9cd0kwMln1sD
PetkA9B7JBOzylZT8ywshex3KHsS8JVyuRfQ/vOoi949DLQb0loDZhuP8hYwNlnXqLaf1MRBlJ9d
zHnKuczwAxBCEXoDaYlZOlm7pJaRvNXLK/jl4biiNCA/IFViTYHSu43/XMAaiwZ4bpdqNfQQFaAg
DCA/xF8skPSAR6YqQ/fP5+Hpt2OeuASHwgCohJ17PnHXsbxTn1usPsCEPQ5DRSAqMlkTVhYeuTC5
ftOZT+12DmMyI45Qegs+Wqk+EH+x7z22JIi4n7N1xSpW3UGX95UtdKZ8XyUteYbZyt52L7ouXMeW
q+kcQc3T7f9kgaFcunu6wnnYRXw4pg3QKS6nxxK6N3ND0G++TyiywcvPwuiLX8bZptxkzC2pn4H9
Go9QXX0zHuTmIGkaTyMpvr0kRqeGLJDzOp+fr3p51sXO7grcI+LOth0jelJtSmwrhUJleyZcZrNw
q51x9gAJzoYVKQsduKfI5sxgXql74BK5Na3Yb3FDGoGfvgCdRHkZEufqmHj+fUpyu4HAUf4xJe1w
QixHOt7HLfi4qOLXj+GdcpNsXS2xSlUGPwiAuKkCAq0oPQOZ6f460afpUJJaWorp0Lx5A/EOcEi1
lV7U+xbnl3d2CCK6FwEbxpoDUBu0NHAqpjv04UaxgO2NBaROCPG+aOXYiqr9+FoMU3r4MWYSayUV
SCAG9sFwJFRiR/ojYRA9q1zbQfzdEpBlzjnneZsIszdIR+nX3dQLeZPi5H6vCPK1CB4QD85XxW1E
vKbR+P3oy9sZruIVKx7bEIw7ePj2yb68WEyGvpx2TOZScl/Z7tLc10Uyn3whQd7CBFpi63+wyszV
NzbhAnAWWN3lnvrQELrGeaRA9Z4DNOhhoVIUl10QGWBA+homA37TunY1m0GwW8DbhYimiZvjz6/h
pkx1zgqP28KBhULqcXauoJvq7wQTgJYnNTMa1s148exKI1IfB2x5jSgAUFVhFK8XrL+d8cofaWf4
mpTOvLI5ssKkJI+5DXocTI0dPTslzJM36xZABLwSPEYSDYY1sQFbUWoIxZgDa2cfXU5ARVv6hVuE
VoHOgsxtW79f4Fz+aWVM3Jypgh7JEt/Y3SEROuTehSIHpgPfgg9E/FGpGG3P5v3DIxYWejH27N94
ConJ6Ohee1oh2KHrXDayBl7nC3F+RnURFfbjE7N/bXEzAqWnc4nEWV8GZyT4VQZDrcQRMREM8QL/
uuSWY+B8pf+JwBG/MEBWsxZQ+2Ro8Mwl3Sz+oWnRBHRDAdAnk9DL1cx1u5RLI0NuOjIchAUJmp7l
wIGj+QeGSNfNt5xAKiRIU5CtDTQoBsrKsBwWuj0WNZIU+h9rFyTdTyu2D/Zon3H/rGwHZva+4bTn
79H3v0egcozEegw3vfKeE6IfNFJFwaV9Eu8Zzkobk3mhp2rpHkFURM+uQiu0BXXaDfK0jErXPQ4E
IDbJxIjV3XMrl3Yxo0HuVub4j7795D+xjTbSQpEpbvRA4EGul3DlK1c9mKX9EPfAeKt7EH9m95ak
CbH5WHtAmMT5Hi5PqWeim6PR0Sf6Q2hdE5q61jhYBBCb/VkaWcrHDL1J75XQ9AIPuXBqjEb5WE0x
v5FtDUqffrn1oZbcqrxzgSqe+8kqkTwdCyCQ6d1KU5eh3IgORmIiCZ+QRZsx2VrRC/sx6IpkspRV
B5ZMMy5EID4plJn8bZEnnXAm/gnNiDB3YUtvbw/pt3LRSvabmlbB2IkXLGTRSV1suox+KQ73JlUr
qYQI8o8JcdfP9R5rP/195YqcEYQMg2HsliYGAVQNf1qlird9aaFWiFP4Ahg/BcPyoJiSXqHF4tEi
3wu2vNGav+8uJZZueDI3F5PjtcsMC3yq0rqeTNe8LgyhgUBOenKLvpfDysbEL6VXoEv+js5HghQl
2K5YTWFa4h+a654lxlFei4srkniJyjVFJFOetamnExtqC4luWZgkmIvvkduaKmxcXkvsh6IhmTVC
ZSDf56Dv+Bb2VzsqhFtaiUDsdRaBhcsZp0BF7IZviKrqFlbnBOId5R0HH7yTSwCeEhW0fksQzGht
OPB1zKxLrCVrKj8M31JBULApoYeZyBGZ2dvX5PHI06c+4uXgRXO1vuRWJsflPULfPAbl4JJbf40o
KWpdk+nTc5xP29RHjzWF3uzb+1wBx2X+oBb/AoHBdcmMIQX2h2DBCk1sFHHWV8LDuEIKfYvQNWZA
fhjbRWYx3ZJ0mWCrJAW/MpflSKc9g3N0UMwRa4qb/zNFXQYYDe7Aq7ComU8qnVPzuH6vEs9NPvu1
fyw4OVAGNKhYduVPCgjd3EheokFrLdg5vRjSF2tnCRoPriQaKIfQQyEVMayQK3ziSlpxDQp+/TeR
bTVe0KPPvUNcer3xWDv2lHxsRW/hbhKHzOyhct1Qgr4U3C2rJl2EGJtWEHyaOk4NJVMzcukpwhhW
sReQsBQ5ELUED4NVsvdGipIO8zvrVNse38aTqf9t8tFcN5doMYLdcox9f2zRUQV0JjyFF5G8GJTU
Bsysux5moR5iPKDrPY25JGc1z/5X4tL7S4KJcc6tb4Cioj1Hmv7/UVO0Psr8jjE77D1ag3q7stM+
03659b6pUfEcREQJvrAh9r5bar9VrrJm6fmLAIznTfb9kUefnq6klajqxoOsqOLi03NTN0SccQcK
V0GHL8vou8iLu8WfMkuyQLly1UV8qAbfskMuDKszOO6pveAMJKyHHl52DHfHMVlmNeuUof28c7tR
drvb2rBTYG2R2Y3s5p5Ep5XinCwW7eygigZLkORKg+Xq3+Cco7J29FHYKpjfUN+jFa3/rgPbuJap
Aub7W6kJG5dS4jcPL0skwNhkRc40Cz6VAT7NN2lhqdq/XEiEKajV8m3bjjTyAF/lyP38DpJ1kD2D
D7xMrMx47ghWPcHiyUnTWgbuTZcAGvd0ZKyiC6Hwjhf7PNn+OupR4aO8BWCGnaC9YIglvWQ332/i
oscduhG2GYJ3408292mKVbdWBRjKuMdnnUGn4r8UO7qhbqEjH0r54Cy7qbjoYIErjqAA0OlhY4ry
+fsG/rc3H0/RYZ6Cm8wG/CbuN9B2bhG1kY1L3JANP4rMZTcIwmdq0mzQLMSQU5bX9snqZE/tgCjE
T6MQG5acE+E7L8M6c7yrGU+/nPSGUyfo04K7AeUtVgmw4fYKacocc0Qzquri/gCJKgu2tq1GfJ/L
P+6FeJzmGWWlT45N/Nehi5b0rA0Ujoo3m+aAeXyqCtiFu+NUvZl6WXbOlsXUEWOKgaF7dz4a9hv8
W3xNDDtrwFiZucDbaTDqeRSZXXlJhgiVIZni1xhL3zoN8tec+Hrkr3Ai8t3FGhHmyIYzj6Fl5js8
E7QqgA5D3XNTXaMirEDDAlwo6jeCwv9Ov9p2+3xtuQNSf3VW4PCqizl/xusL7a2l0fy3PmA915PN
HT09GaTyBbYGq1nO9RVyBTVQPsC1vTTX8YExHmIYfhIyTlRrP9ZD03/VTs8epZ7BytzBIpXD75zG
j4VfeYqIjAOore08+Nu4tEcb3kjly/PXTdfx9LZQaclGfoiPN3ieBliyWJSnq1LKGHZRYEz6/gj6
vzA1Pv1tEoPDpHPjH8uU7QwXpqttIRjI0AgTpTA7rP2Gr6ICRJDuF5PL3syzJGh4tJ0ELP2SFdg/
52AmAGV1CDO9mZYf0GGcpAIlglbKbJjFBADm55B45negV8g0KojXerzGY+OuUsh0+iHyIVVy03ht
iFHPfdKQ3IdtGE/W6bcxcYY4i5FbzswOwpaSLTsUAcaLQ1afhcOG0Gx1WmuFoxsXKekySjmflh6L
Vd/Jm2vrDjXiQBmu0ArS5O/CC4VuN1DShTyJUbdkiaRwxP0n58MuyT6NtmcZ4+KiDsASGBh6MsqQ
WwxTNNVvlw2UB6QG/GSRVmQWehMb/Z9OaVIlmcXil25vTMyeq95y+9eWePF7+u2B+RKP4kDqAvHL
LDG0lYpqW6QqM1H3jqis3Bh7jeTGr2hr4p2ukdxIeo3OWuEvYUlfUAe13ruoFtLDn1nvLhVZ2S8c
3IaTH8Bj0EFhEK4cX4RZ8dkGQhtl9wOKPwApb87kzxOONsVqA1+kHLWAI5VaRnRYYCUIO3ZAKa7m
G9tLcFXF6RESZ6x549Z8x98WE7ZaDvNUE+3Q/PQGUZzKNVGXS8ppkHnAUmlFZhj+AJ0v0GoBPGKK
xIqi3+jx31nq3UpSp/pnHj1M89keWXGwaE3xfiilNnAfVyOmtmqTud7qjTRupwGitQ6EZC0F6gEi
/KEv9rGDgr5eAH/DJInoWhhFnauIFsvRQPesr9cS/KjqmoJBcmJt3MIIAK/Aqavk9SQUtlVlpHbz
FmirIJy3PoT4qFGctnjNxW21avF15tc/RoYvmwjH6k9jlw1pFiIs8jcE4qVLui1K0TUw9CLF6Xbb
lfuYUZ4pTGljTkodnDDw6PuYLr0K/kYlSZuONQsF5EbIvxOKqZUI7SHvb4vmgB7CiKCQ09oeVE3L
54aPuIzroLqr2J1J2jzyGocyZtncsJXp67LBe9JER6f0Z0pZm0h7R2ZxfRR4dae0iv0UaohUDK6G
ur7Io9gfkG/Im00Sto6udjFUei+2qc07bGSq8cVJmpVguad29dGeZ6K79ea8GNLRJlVR+DL6GX6N
HbwFWZx6GQtl5yGw10S8n8iV8NIQf5HLb5SZQxwkzcyjHO/WzR8kaL3iKXxQJsKAjIIRtVZI/viR
cNSOENKRRjuJrIDk/NZSGN9IRfiPTWsZi1MAakzWKUWi7zx7OUQJ2r8u/i+HSo2XfdliQXpYs+k7
FJ2n+W5eNs9FwV62IgRgxQsMEzO8YycjO4Fq0zMk/QXfaUf1tIjubc9pr8kHe0aE9R72jDor7c7v
QIpwD5V2wE2VTcJf1c/iEJ0LmnngfNfPYN44xtCGnmPyfHpPzD3g1cEYP/rR7M5R7JwapWaLkC6z
ib6hE0rDE8JCIseWJaXGSBh7s085efTyjJbUJ9+o0mBs+Ce7MPt99bpp5Brw7M9DFxqsSuHc05E/
0/RGwpxnDSnpYVBUJZEpkGwxx4OMrtEl7M+r00n0M7/GjfiL7qTX4S/LUTgmRS0kR0NmAcJlf4Ox
EDTWzZCS6GVHC5QU2qxx09Up2dDhkhVqIwoFsJWvSOP9BmhKzkgwKDTG08fYSnzNytUjbZBmWDuC
j6u8MRcyQZl4WC6eLv01OSeEfH9tS9wv55YhFkLO0Jz0A53wCXhR4dY4WYT5Qdjf0gWts74/4fuI
dD0CGrQ45Ucn5fsQF6uJT0Q5f2cQ1P3tQVPIZnKc8Q02IDq6z4yjjt+qZnOGDBd9obClkUcM0s6j
raU9BCrVBc3/s1mH5gcHNul/mcVxRbETdxAkTQWQX7kkakwMU5TpbaF33X/FojuA1wYlwmoyO5mz
UywxxmZPzzv9dMaOPzyT97gFqE25U/uduBplpoQ6qZBfGYdVQ4EMfhPChb1SeTtjexR36mqgDLb3
BrdKpFkgsMTkvjCc6fgJLpBuVxqpepPuL4bpmzyMXWkW0YlnopDg/C2nHj1mYqpNyzNRM3r6lSsr
wZVse0kDc8X8702TNwIVGPCIfSCaNY+Zy+iXeAQNYgRD0tNbiyu7rP6VOTyTmA2N571mMtYJgXcf
HbElpM8YMCQK6lMUc0r602blk+nYC024tG/oWwAlbZAv2CJiE69sFcwe9E+s2TqqHXqiFmt5a/bR
ia8qj2xP0gDrRSOCjsE3OQ1AH6eXhkGOMDNL7Uwfp6WGo9JpArGDK81ihV+q+6+t2fCgNtsNd6xX
MmCqgRbljPPJuuiIKJFPzyxFWCJZDO0kFwhFQ/6dvGtziyIIoIOgvSEWCy8FlS4a2tssk2fs0d1K
pVExBwi5VTB4OfkGDSujZTNq+NVzBou1C6RDbTWDCEg3I25B+0xKFZYQ5QG5/f0U8rU5m3SItNor
3JMvEI0uYTkiqxBj4g7u5xlh5LcCYVPC138hsuAwE5sfK0//s32DRfHOmmUccCxt+esnBKcA/vvP
XDwyFQUoYznA/h427XnnpPRz/cnDHfiia5yizBRSd9cT3GcMXalPPwUPUm8f2GpVCiTKFVJPlWDv
KXZx6eGYfHQs8rTXkMCqIlHSdqjHoXySV/xQ7U93p9CJygRSdomQ47Uq3qu/ZGVqddqRpipCV0uH
cRfvUcH8H0lGCFYa0E5NZBZ7MtQkcNXBZb+moYm57mLKcMoZKnbQRKO0GH0V2CBTDDWKo710v4WV
yk3zTGocWi8ySPtRgkejOM853uPH3m/QryGibB46Yzn9OEaY/tWFvDKR7pWsHe4sY4rkCTu78riW
trPpfoitYuVper5tBWORF2UxJwoSu4rE2ka/gxeFDhGWDNnUtS6sOoVoCDjY+nrVQeFxnMAFaOS6
Q+WpWkdHbDtx0mKH5gvf0Ixy38gRkvPD50CR+iYpvR/jPj3EpLexpVWYYMx3CJIbUziQdr8RcK2c
6unz+lniqIqAlWijeF74fF+cI9bzmDH70wBiksp67tuJ22tNmIfBakax+ZzMG5Yla7s/PqVCDb9i
p/QvICcRe+vovalO1ueWnV9tk4EBEEXKxfoGMR23KTQsV6+cwe2c3QIEd9bPwdEOsTCUHqwse1lr
mYQxBjUE/Qgi2HgUI3lk+5gJ9F0U3RW1LfFIge74YeOhHzZHE/Dv0EoBf/KEQvbCp/Dzu/WT00Gv
1SzO01cyK5bMdoA7wkE7roM1ZdqNdPkTBgBxKktlD4RAQysOUJMyIj6kWXlmT0E7Qk7gECYUsv2R
IFFN+LdUIUk6j3m//kRi0jeIyiGLvSLx3G/UrZwaBiTO1Gmd3AJTcnxLfRDpjs3e6ri1bM2HSXtl
oCGSoeVYY/ac9r8olx2e98qHnWLrlANn4ZelsLxjIWdLK9Bm7MsZ4z2C0O/4RJgBJnULmZX6xfWA
RZ8L+zrtQza4hLOb1I0ySCTWKAFH6Ytsr5oVIhM2P1ml6w/czbTsB4S5CUK0fAjNlrf+/fuqOiPz
423cHD8rU6fsrrUlSbXYhIg/HTQbzKg5RMb524n5Xa2GvWNek3WmmrqT6aScyFPWEvFdDP/raRAv
65uCMppdh8BwcVQJGCizU7VnfyCpsl9qpSgXE5Jwy7ZnckM0MztJdUBFxtWxStV74FWSZM+AHApo
G1QdVD+8nsSF6TMUFmrrrXsWRTakzFKd79zNyewAXp0lxit+7LcuJZd77iZoSHRYMuysAya1+jdp
LHY+q+f+ojeCzDtfps2U2TzKE+YTuF5iRZ9HhJ50LYN0XIofmYGrsvqKXp0W5XaDkwoIOIBTsnHz
J6YPS2+/lbUkW2swRdRTcaktfCsvpXU54VGAHjjU/BzUdZgJybkg0s8d/F8HqliEWuz0g3XIsWcb
eKb6gvrnaNASyq9S9X1q7UOS18OhjiTaGlCj7t43ZWJwQBiZuGiWy5RY3pDp3Rm0n7Oy+YkODSwg
YARgnt2x5yg2jllP3t02fUo8AttNILGwKSiUdev1OLxT8SwJ86owroDeNW3RroCrmedjeDGJKros
klA0NT29wiKUAsiD/eyRQdbQ+zpaZXPGwr/EdZaFquYi8Sl7n3IpEQG2op4l3yGehNEdNFDt31aE
GyZGT04/u8a9VAPo53CgomHbn+JUpv3eOc945KiKF1XOll2OYKxhnWZrahKgUAB+7Y5tddR+yZoW
0+Wz1SDiKRbqa6I78GjDl1H6AJFfTJCy0iMxGfbmoRRs50HBPHJVg4f+C3quke02Is4jhiMkg41u
U+HYMAhNeI52C5cCWnjvD5Bu//cA0zkMLCkT32S02yXe79ZUfAIyikcSbOoAjWjFG+ouMgAFVxGH
EjSXXQxVCcPoM+iPjcgSawDuo4Hxnv3Yc55PlkkSA7gnCVUwL6NWwV52qbfYE3bjtpDSMODYg1M7
iX23B73F6WWJdtpDJqbQvqqgP0jaW6ObE8wo2+mzumYVkhq1IjNPh9GHHSq2Rk1qnrI5usqTFuv4
xGZ6OxfkNeuObJN0s2TJiKuqrqTqm6eHslBnghv3t4jf8CTBadRWsSWKzuwIFWk80NUYncS94E0o
3Yz1ZTbFWpVDDX0FH9UmL19VKXxwtV8sDndZCOf6nPUXVY5Dl1kI3Yxzg8hP36wtdiemIZf/qO3L
/jriFzX6azbwzB+IQY/lbnfayWeS8pYlsc1lZvn0+YbKlo0fHO5D4Up5ErMJvvERvS+tLh1RMrmG
/80HzzyPzhVt4CsrFis6slYT5SZgIJftkAPTadkyA94ovKynFJNhWOc/Z3BbqKXSmji9sn5+KK8d
EjI8kFH7/Pp6B2K3rfFrpRlYqYQrFJTMjemvfloK3zY6YeVE2xsgo7mnvzTD9ZuOuuwZ/UatKR8y
OuQCgAuALdadPvtViE+I9w8wcXzXhPF2a01GxyWc4pEgWu3EbSmhySG5WsOpJqWCjQ6OiSaU9dYV
R7ibS9hrtkryxkhC29C2zxIg5QLA9TNvIthIdJy4AdHvTOHqb5gVxdEQaPaRgPrzFldSVB6vyCWB
CraIVPcPpsa5+sS3meSM287hrTxtxWiS8/50N8J6Hp/AF0O7cUYuSxO682cZxjmdRc9/gbn6IsPk
vrLur8Dmov3cSbzCvyZdG3KAAJ1YPyKeN6E3PidQwDMAKx8j/2YqNoVq9BMwdshwO6VMtPAB2XOW
3tHgA35ghGzPuJSw/kKi7xG6P64LcHW8n1Ud4/8qHG7HdthSWGEEsAVytxVG8jJVoy6ahpPFvJDU
XAMyeN8hMqDS+PQDFrao2jTyD3LOVKoZ+W58V6Gw1XfzEwYHpdvXBHCRcivqQnUrtJU21FGdGkKv
fcSgYmU9ZbunYK3ygzz1bNoTNTj2GKsfBYdGUFG2qQa9l3gy5WKeb7l7RDidCEWOrpCxt8zsPc8p
Cs2ozUnRuJUQsPyooYz04olf0pXluSnsp5NvUYQ/fSrsg0C/qBTvLv9zXZyhDQmCvuR/xJRpBmg/
5hvpzyQUPM7ZKCM96eDShTutpLjaMTK9wZcRR0ylApb7fIx+497XCwrdev/EhOJ9LCUD5P8m4XaN
CT6n0CHrge+di1K0m89AGnaLlcvO8MJAsDDTC/Vc1cvRqkg1i/XCq7nvnyeBkSsMPJAC8I+LRPyk
sjG3PEglGNNM5PuMYifcJMhjUNbs3aHwoMF8ebv26bj9qTI+3wlDiictxh/Z8bfdz1GqJzRXvwD2
df/BlhSPwrUU8+CvFGrfnM0lH5Cs07BUEpsqy/32wbn2/5a25hycXBnkwx/3HFVZ3O61Go2qKVbK
OIi19SJ1YjfTuInisZfPkgyDBJXI3D1l3iM2bDW9scX4pDyjnhprmHaRRQZEM6VXwo3vuLwyraQ4
y702phOi35jDlSg/tV6XFpozUoYjblA9LNgm+o6cHJ1t5qYkgXBw6WI9fsn6D5ncR3SlX9NZwh1t
ennPsV00u9u4El6NwU7YR0H0YeP0J/FlDoLLprX/uYvF8f+NatVjtnH6a4bbfBjBC3CcDMy+Pea1
i4kd1AcZckeGs43u1+oTgKo538gF3g+odlCorB+ewQidGNs6SZE1zrKzAiWs1JXGsEyUQBRblhiG
DkjzJyYNCAnPUPJT+Oeo6LVJkK1krRhGPsIyMUriim7Ah67ULZVRkU7NQ5qJeuB48sr0zhcWmjxb
gHEnX0nn1sAjssL7NpMlCsZJDU2qLwCQdCSaWvuCCP4lQ3XcUUFQC6KEHtmiGcc8JEVRE7tmrug+
IPxvQFaqTHX8bDUkL7mO+QUU4fTEqPTNQkT3mkSmy+caBcqj+tWUMSQircwVt5QOIox0wXL4t4X7
gS0E/jxbREMz9gQirmvq72qZ6prUVTIN0C1dF8UgE9TP9L3J7n9Fl95wb6rGk6CMOgxnmfDRnR/z
IuF8HqGixdPCTAKP0XBhz0KO1kdqPe4wexe0fWhKjqkwwSLX5HrIGrWkZigdnebtN8hLcUGhgKKE
Dp4qZcy/Lo2JSyZCyuB10V2z2Shqh7jC0WeZr9Tvzao4qhIh1N9qhhXOvseVRWiB+08miq71vmle
y8MCoanzao0eI5RaCFlaixvG54nqMInB8w0hJLEikHoOqHDI63EFSppN5tk0ORZ6ooMK8llTnTop
DuUTjok2yjqhv3bMGgoJ3wHq1ypvkOd+wIVbUQwBSky0kwhfvvfJotfrPeSp0VofCGJf5hBH9Ttv
l7Ziy3qGGXUWeyBwJAAYtSEXm0p9C+MuEYJ1DE8fJwA30Ss1zGddlKdbXkn//aezj+jZBP44ywXh
MStykKYJWVFgqCvb4WW9kVrfrJ4IRAKsZH1RHdU3eS5QZMguxOPNYf2PQN/kinl8LAekUDlfnrOA
PePyJkOX6MA9yQ1JqRc78cBi7Khjp2tWQGZx9ynYnu6ZQyFG+Y8fx7xI3esOSIBBV5OblgFQLErf
xxINADYB999V8xk6YYx7fj4bmlLvImptywBsT2X06GZcX+oHx2GGiFceAMNd2X0xbJUx3PewB9/C
CfKfwJw/WaSf0v/Tjpw9WzJEsznecvMyS89HzqFfwpM4G1lk6q3alROGXcGicbkMIWn+24L8PVOS
J9r4IROWdBdQHWPHSrfMeaks0d5o6kBxirA0pZ5iZjgY34okNpIB0+ngpG9L6YLqfzXInN5umZKT
DdtuLi0Ep3VUVGTNI1/t0HjfrUxCS6SW+YXN4+fFTT9oCRaRRFGGKDqwpXHD5+Ms+7e1nf7KPBpA
LVPOr0VfnQ6gUYa/Rfuq14si1+KWjXV9umA8Wryxmhjz1CodEVqg6Ax0D/v0ZDDU6Q3QMYXpJlaR
R5t5eDx0m13ohkUTsJQ42QcxzuRyKlbiKzgNO9Tbl13OHxRx+Hj2VJsBnaH/MUsrkGSjAYXIL+Vh
GIc49KUC6E4GGIw+rrxdRwFVzBg7yk186UimIDExVwSsfOHdhHCh/6uG/r7ly9HdTSA/o2jY3DQe
Q0vvXeNndy0D1Be70YJEjFKCllBx8lLOEd7OeX1+GboL+lfw5C5LhHwpqSRAiTuOVYqWjclykQrT
u5sE59CwlL+qwymYyJ0yhEAwdz/R7rAJMv0f3qz2oSMTJK5BZ/7QFGhUCGc8FfxFnda20kw6u1Y4
9gU8CYVbERBXIarMT7TNwSknoC4WXT6ZrsjA47vpjcGIOn88wdoZLwJQajsWJDMfvPp8z6NpskFq
ZuHY3ua8Ryc9/7lXxFwig2Pnyc/sJ2OoE3fZk7iwAEGpCzOZS1I5c1EFlRUYWgCEmovpMYralK77
ATB/a6QoYLTL/iYy08/wZzcp5ltL0MH9ZizzGojPJDk9frEECgkic3WkTkCgQSm+Iix5aea87Im9
a1RrmRBTw7Qiu6aAi+zSLfe5bkWhVNCyOBgkkrwTdEHYSRoO5vuxtV+2hVZjPAXWpHqLtiioG5Qq
Shz0f8ysnBNzkiMC7u0fx3Ui29r4F/G/CKcL9grbTICff0eqcEVLIMLmK5io3rwk83acCp8OVe1p
y9kbfqBrkEByEKX7gj/S2UnBYdxqMpRtXhTXa+sDXo4tvMOLv7lpXjEMfmbBWlXqM9a+Mepc7RsG
2C5mSxXO8e+0Fpsqw40vBIC+fR68SyT0PwLtYAInGnhg1b1UWeO6Sf+D4lUNkV1rlOc2ZIAiqvAP
rUmGGjWX4hVSNmgNFuosIqAUYQwgZ/d9ZzYydTn7r4AoXvVYoPdUb6qZDcOgSjtee+jLWSlI7DS0
gEKUH4d6brfRDJZlL2WRXpV4nNSORqp4FKmqMZHaojCPWH9PrnIIo0UyKqyHrZy4y4zxCAukveOR
ORXeYIisinVwz8GwXTxGVFzvCnFzKKf+0We4K/KnpVGnOfFC3SIg0NzMQw1f6Uzq0X0y4vp69CMK
x4O3O1kvnZH1TYqehPl8+YIwfD+zuTN+Z6tjmTza/ahEhhn68Wu/AOa8hwLk9iylL2LFUzVmMCPH
o0Ue1lOCOsLjGcihJ7i+l5J7Xi0PD0dGnk5MVVUh33hy+3MnuENTsUTbtA/LeqTZf2xerzIzOBLe
f+X8NvepV3ryHcYS5TuzkXmZsO0IUjVWpR0Z8qme8B743NXW3y456UrBS2URTHjb8lv9wqPk47TQ
VanjbZBMwUEgHC3RNTP6gZJktpmT3ZH4iKbvHzwwkZU0Atq59u0THGhbz1uVkbCGybg6pdMuVQXF
20V9lp7c4n9ei8lYsQQBv+Th4Xh29xMJ6b09ta+e8bbDe09qx65VbNQqlzC2DcT6Jqm2ZsaCuvbY
EaMSFLNZxrUnSiYkSiY54ENLaGv4dfJGLW6Cc8ISA/UH99dFFz34tpIIKkPHMD2RJX9utXNAlCX5
OgFPxcP9xjJ7rJNLO1izM509caoilDxIbxfUJwbwKxtSU16xHBp/Q8IGIGdICiX/cC5+wHMbMBUr
ibLhGxzyoRmlyW+AgEWXynFw7LSLZkEqzMUSIt7z0gYL2SJ7iqvLWjul0dLfs1v++oMnblSO9pfY
wdgs9lvo5hX1S6teOUdhXQdK1NM6A7zyMSWemMNp0sW9zFlOarSmYNX0eCv9pnWNk0kEzXf6iNBF
kIqCPxYv6RhUIUXT2LigsShXRSeXvOQC3Dc6BbE/wUNnZgVHVGsTUYX+ZkVDgqcV4bs2qz7ikZLz
i7uMHICt/Rx7DNtFdQxDP+wFhdy1vX1O31V3WUcJl70IcEKAza2tSWwXuhPNNaYVVWj8PAoXiWMp
KDpPNdYA9vM3PmtSgbmgUk3lw5g6mp2G2ZIeeWln/zFQx3DxmNbCWm956GiNQ6DbQF0jfhvDsVr+
0rHTqNQLWabTPYvskivnr16w/K5oilQ7GndRz3q58q7zK3Vy0+73b+ZBxkuEeX0BN3VaeeXidp/S
bmMyWw/qSkiK3E3KT0EpOVJ75Cn5wnXSMOEibMp4fw+cCzLFauoa1GpGDeK0+2AlSddaU2d5V7AZ
GKBHa6aoBuGwGdlRrY3/ONFBTGxMl2yzRXu5/bFnTxXWIqwy8K7URP2pnHA+8XQMG8rBNsqfzkkP
RbTXBi+jbTqjNWy2PZDYXRt+QKy7kRF/R+Ra4Qpfx0KpBaeFu6APnWVOvwZygLMoF1gCEHyaUwFQ
mjHkA7Y3kAQbfZw2c3KQR9yUtdokJRCm3CCsvw4v1q2j1BUeSdRyk+jQAzEgzsqRkWhcIoMQvPDE
BjfpsdihLPXzSbmyNd+3OalYqmBT8mXC0m5FXb4E9I9w2sudfjuhutbQLG7HdSR12i9IgJMQtzZd
2K4IA9XRK1kY+marGuyC07YZWQs692UF/iigAjI98dWfTqDWJvam0jVgkEeeMaVEJGQ1z+wLKfW2
PBdQEgDG9sls3vej4rr+h4MYxlFQnNyVSRTkOWiMDzM7iEC9s86rwxi4atICws+fOG1JnGpSsNy+
y6NSbniOauq1YuWchDWJTM1HeuZoNo1zKvcLmXVfriztnJ/Btt/19BL2SFFtE3YcunFmX8F+x1GB
v8xgitFzUg/Rc9wfpwpbrtYpWE0f6KjVRRKPSgzC3KZtOqQLz3dyaKlFVq7Jpdh1Zv8ijvngc3eV
p8StXUXCKFRwA/QVAnx0oFN/hFRhdW2b0ZpnqmB5ZPZkLagt56e/WrfhSR+bPUzp3cZLz+lcBxRU
q2gI/BS3h7ojWttJER5+Uvon130jf2Xy8kfg5cYEfji5Wi6KXFoSmZXRvQG/cOajf3psKf4I1fm0
z0E0f9AwPmE7SBiFriGGQLJoEcV7IHJ7z6Hrer9XC/eUqZdyT8T2krSO/kxS5TpNvVuSb/5T2KWP
WPx4Uf2cIukEnK9p5QitQjucrdrHEot9c6Xm+3CL8dk527Rb6yCs/yMP9l/FtZjgzFSyXkChXinb
FuJ12xBHJyiFD9/YIRztkqIaEYkmbzGYRn0EUPAI/78tcyViP4fnaApIMimiS3Nc/8hfoTx5RiFn
3ZL0FXU5hYWl/fy6NvWBm8G7fbOgP/Nu7SteGTJAhoB1fpYdyD7ogGD9ietDarZjDCwuAkxWvZBH
FEyOdqNr5YEVhC8k5kSrTiMRgY/JeVDRjVKDDeGADvPMUqJP2BbrmZ1LqBf/fDk2JJdB4ggMCRkc
SDQihCLC9cjuZXcZWRFwjoILZ4H/bPAG73AQciPCJ3wdL2qOT2kEHuDd4brTx1uGBCzK4k50fD7y
XqEKkStpQDX002D0TDNK6QfI16/N3in6CoIuCzXGwpQms2xR7cJ+srQMWwJN2aZQWEqPxd2lTwLf
A41jLDMeeKwFbHJBitiRB3OESjOnDdj+8pdfC5wSt0YgZFF7vOeqUePhZujAvVuIU1KQTVju7dCz
am/STIRD7wTpgnMX0ZSewUnGvyoH3FyeDZVfGwsoO6GYI+d8kPc8SssQtfy+kySs13C7BlgKrbra
mNKga+LbxWg/VA0VxrJkBkvhy4YGMHCLhwj2b7l4OkmOWV2hpblqWm1sPoziRaT32Bxny/qPnNO0
77dg8C3/M9rfcSDJ0xY5F+G04tDNBjQPqCWjt6JGE1sIoUAt+uo92+qaNvsRAKXbmxgSWD5epN3c
5YASY2aQrxrtbBcNGSuVsOKhg7PKRqImOxA1wbHiXAs5eV845XzEW7xiBx1dXv0G2ot1/MVwtlwV
pIdEfccp4RvCPwuWIwMHXiqhfPJIu1rncOPzxRyWRwfQgXFqZj9EioHMaJYBmRrRDCr5JWH2x8jp
o6DXS6WCkVhXn6PNi6dV9peNS7jC4nInARLBw51Ah0jcJnVpAfJ6ksGHgOTn4DuW7Ca9qOiVmV7c
yQiC50FUiPYZOER6IMN6oRkUQhCdg3e93BQy2/w8Y4w8Y7932e0X0EJB3dtOiPwZWKj5qGBarQB2
8TVxvLym2ZinLtmiGyW7Ouhb0Ad3o0HMzzkXFQJYawLy0s0SgSS17M9aKNQfugNLk76I112TOm6m
EMGsSNkw75w/8FJnT7nVd4R8SnSvsVBatHJIJ/Ia4H4r4KcAofhmW8NOkCjYIgahG5lNUBWXfB3y
bt/6f/lOYRJesD6r4RDaXao88dQqPA4hhRPbIhagnVKA6siK0iva3mOs4uvVCXeDLWSZPy6xAw35
JRt4Q915wwJprZl2RRtm4iObmcEOsHVnzhQt/SCctM4oIdrWUCmX7aFhTG2t8flBIrkpobi3BCCm
EA/pQysY2fYW6ElIUeLXKyxFvESPBr4oJv5qtuHt1GcF5aLcJEj6Rb6K3iuFWoirCubhmfZOZJdx
jmrX7otkX2cj2yTt7bl6eaCom8sOLZLxjj/X8RijJF+c/czcKJF4HQOSNyGFFFJUfxqrvwd2nIZD
DYLRmZ/ZhsEct0o7l52uq+vMXdye8N64T9+pw0y6CcKeApInfTBEqhvqz8Zb3Pi+5vSZHLsqugZK
t+fUpz8eUfmkCijTjmDedunh6PWkfcGN2Od7ek9NBUyU7f+zVvNSUmFY0bGFaXc5jrQTqCS1mhsD
PNODBd1IfbunyP/f+WGWe3oPHU4hULHzHUOfgXBChyJfGqF1YwJLf8rz+PyYLS+0OFIK5zNnGIRY
yu33XreFUoFnVL/kyRtADOXOUR4/vkVKTMTdJ+gtOUaST/nKfd1lRHHASmOyxlo8V+y94dmdtpzJ
ta9kDnyJErjnBpfoM07yX9HyXaOAn/YWKEx5+5J6DU0c/kaetdlpckjLT3vkCjy+4UiSZPU+93OY
yfXbJiceuAwtX/R3rulBumxjsfReJUspAUARN0sjVj8tHt2VrGUu5MMy5xBW8g3BskM1IN3Je+0T
jUktDmIgEWX+7T3akjbhizutJekRynOwNNNHb9Pa1mAqWeXq3v3nSx/kSPAbqVcE+of4877NxHvi
BY+QY7m95qzga57BFnLs6EU6XLCkVK/W74X+PT60jeXzlHEs739p/DZAH1M+9NnFfFF7+B/zNzTQ
sDpWUOX309SRYxHstXLBZ/UnI4SQxSU6wOJu3JQh0xeo8TY+A3fkrRRHJeoZG7Glw0ku/sMmgDgU
pru0o/SdKxTx3H2+CXDExQZqJPHvdd9AKAWZUAs0UiAhn/iaVjB+ty8h7Ji9ZtOq4NNQ55CRV6cg
x3GEwrg6FibmlyaG6g29UBILLiA/fPhO6Q63HS+4IwfJao+qMlC+CVCyoV6a7kB1ULpM+pHpvfs8
Jb7Piac//TyBnxvvbhuXhqPBX4ZVPLvpK4DxqJ0BLBuqCfzmtJAB68BSfmhm4ld2cTagI0ZUte3X
EWzxeB52dTbM8IW62Qg2GhI/BTkrRw5o/ToVM39kTrfcUY9AGQW3fsIR4L448/bHMoHZ48FE37qJ
LqaYHI8BW1CGMTV0fbate8PaBMg/xQvBFg5TtNg7el/FY+Aggx1ZS7yJoexPXo/hi8qONqpICkgu
B2qAZVnScwfZHOD/gDpigIXohRVGq9tdLnyZvz2+tFJTQ+LeyycABWGAUtBqO/RlHC1Wpp0y34/8
23WEp7LAYBwJHEEE+I7BhSH31XSTi+Pcaj2rs1ncO56KpLMfJnrpYyy8xxVMAGxYD2mjMHtEwALA
lerdVBpCBTwKjsGsRoUa0ezsrOr8wvRCKZ4yihe7jGHD7MIztJxsjePRm1Kql+EGEjWMtFrLtLkH
8hNuBOdPIO7aJXaeJoeex5D+bDR4YIjjkF+RaXcK07Fokkil60UEMDg/xuiuiM7G3u7pEilvhjZI
I0PZTFOdwv2SsSoCH1pX/cFIP222apPMtGwsp4KIKRt2CldOLdFMW+2PYI1Q41pJmll6dmbf95CP
r7RM70Me7hXCOHYZGOUIs9Vn2TlFVDc6xypqTk6jO2BlVrOnDXJ64vclPgD7T9KIuWZrhjBR/SFC
RMQsEn3JVfTG1jdlq9RB2ec/L9qYgKziVWvs6RnLcSqDCuEkAMQyz53r3tg2eVpyvkJMRRQNbcku
8sWy3ESEwnc9qxp+jVYOEB/cXYkjBIRru17yWPFdlV43B8x2GitmSiIMnqbMZoBH17ykwTS0LA2P
FK92CWB9RMik9oklLhgEOs7FqQiCcuOTHoSsJ4u+we4QlvQzc7To1ZrzhaUMdfbJHQj2VhLNvj+F
TntT7Lct8vDchPOs5AqCPHx7pb/gCPeMlL3j+1TxZVuYtPtvojOnXtCs8lTROmNGGpJeYbbYbkDT
W2/7oTMiBMA9xvfNFycZ9AYcqxj5I6esI16x4zo7YDzDp7A5/etw3xzf7D2Cs/IJx4w9UMQCVFt1
o9uv7YNrN5rruBBHpObuOYJXoV5hR7ynz2ezv7InU+5PapiOlq2C+oMSJn13rkmA3MYXA9jHJ1mY
8ZvHDRYaUjjFHOpszB8Lv9lYw73xThZCGPj6ju4Qc8VxzGNEPDSOnsxyHZWNP4FX2d/QMMXgSLYG
EwS1vtgTpnXSS3TMSn3n3bdRtDx/7XDpI9AFRJzUGR99SDU1rt3hgtn6GhaKaIufv/WEY693On3R
dJMMd+dv/ofjiHuJapZJFFneciyp0Ygn9d/xRIkU/vSCkYbBVOHUPxZa297Q8YE3PUo47/nTOSM2
kcSabVu8LnH29Q0Mjv7UGtlFXOBkQsmNQyV2UBhQhvc4P+rlM5f1M2Zg+SEG6v2fNbteitF5vvwr
K1AxCisptXsNVTkGlAaawdI2lQyffdf0I3T2XlcMRH4PD1MOLutOmAOeedE9FS5qevjrAEwR6UYX
hV+yP5uaxIFWLFgMPEzHQbnzhww7EsgRE9kXN6RGQcAM5FMTCBq09c1CnuSlCaayzVqiroO8n8tk
f13+IKor3HB1ZsVJK3ZLDHbDhbQrOMHIwzcyvbZy4EEeFQtRrAaaF7v1fGFj1TqTovsaJJWONv5v
BJ3J597+3PKJrdeUrfvs8NcH60ecaWlHIRu6P8RfhLdIFkzYsyWGwhVpKXIwQS3a5NCz8R3rYhHO
xZRixCCo6tqrH6vyI295yyAcG/FoZ/+2eJBGvh4Bmu6fpbTKdJs3Xgb0NNBafzZYlpdX+LJBgBXT
WTwY6opNsdCzEJoK1fdC8kbnX9qyjm7WFkV90F1bPLpH4fiXPaHFIbJeJHClDBesboYvlFRBsKZw
rbJNlQc2ExZLB9KYBOeWJ6HwvJsQ6Lrnqz9iFbfBwC0Ut1JWWwlbieSxYAFsL/w50Lhz307SpyN3
R3ZuINBWKMhShd2yKeKW1dAQJGvfsVAUqF5rXf13EU6ojfvxmlaElFf5uIqqBExFN5cwOabEDVPL
8+BLtKksmeM0QhOZlYuO/EuEIxG4iyO36W7Oc01ugXsFMXKFpLaxkUa+ZwEM10HFQUIoobZgbHpr
6BHxU0FwP7qhvPF9Wb8R8Qwa8yPhT/MRZmGF0DdqaYWpwCzh6DHEqAV28wlWUSmsigHnVsQvo62M
A8xFyXmky6lq0IiLL+vBe5TB1x/YgDw5PsfJ1598P+fpkT/scfA3jXqqT4sKHf8gLMqFzP0ih3yP
i2XfBEBDZAg9RPqhJO4WP/d/G7wcSX4xUY+9iA/FNhwZeiPd4bL295f6w9CVmXjAcnQ4mhYWyqy/
NaQBv9jX8W1+GQtccTLNgtKoZXUxKCrsBUk1OQrAvRo9SaIEGVBqPTwuLSGTU17FuuHXfV1Y5RfV
Z7F1GlqFBYOMbpEZ4Hp4xzIWsV5gA/BePHGARS7Fgc8YUWPrQJQUZd4HZWGdS2BO9BOGpE2ctCNo
IRI7cCYd7R8K7ZeAcfGGyTwwUxDrEse09g85EW1UpLQdDQRPzKZFuAj/S2d9TfM80znzm54OQgZ+
08BW0Ako9ip7O32PGAkdOnQDoflqWMYknLCcmCK/CYf+QaKv3/6NSEO3kR/UFmQLJP8/22QCFtWA
Wqzthox3W7rJMrg46gvk/KpPn7mdY6ei7YhDMBBDo672tn5bdSUCSUInEpME7TTfMNuBfMBI6BqS
iEqoZW9zXSR6R7BhhMW9h9xhuFJBIITyMgAAwLvdaRGzuMEQRgUkSSUvdC5reeI9L9YAQ9Hfr06s
+VimyQ3AHiHJjrxQxHQiu0vLZ0GJp3oqZW0QcqbPxZwu6mA/4+UhFhoBtadBVteI/pyg0quhKg92
cBNtViyK3wR01FI4/vxbc6eH+bbpMS7dlWEWln7ruXIMU9zBKSZJUXSuCX+e2AOTfvt9W9fbKYN/
09b8+2RCigMeCA5n+0MSvpS67sCZll+ZPQBuNAXJ8+6fcf/95wsoAahlOAyAR9GIVBEKrubz4fix
U/6MGvQqUibbR+XgZcGR1Fs2j6CQ/eNRQuYGNwKoFzfBGNkyaUQgZZ5CGHYUAflDjLTRWxqR8CP0
zSuweq21NygI/esGldrHjQpEkm6EIKPgj9+84WahAN8e7oOzjs7IveTMr1m/yPZDg+9Hbc212Y9T
MOtgmyCmUlSgex8hkgp7akW/W0OqFCBLmZcnKkEO1ksaFvRoyKwVGglYoZlx55uw0SFtlmXEY/ht
dy2QDxlI02Bs4VoutBfJyp02p51yaGuYZEFPXoFVpYqPpdP62pKuOJ5M//syHg+qMeZXsNBW0/q7
yHIPTxhCZWsZQqH0lFCojn30qlsUhf/+qPjMyY1L1xtcKgpOn7+fqNeJkghO5zHmI8zVC58NKd3l
QV0xDG56+QoggwP/fGfLi5W9gWDMY8o3Z6gs2Q0T9NvjOX0kYyHyQLMt3z2CIG7Ck+Yc7Tri8Awq
vonE/hirgIQ1yVXgv3nyNn0tUCetuG693LdRF4eMJnxImbLVUYeuGLBg20B3n0I2HzcA0pBPycJL
Msq2KlcVVHhPY5DtnOp3Q6pYBvL88sCCOr4XVLKa7LIec4xH2RPz11HW9QctHorPCEaqRzUy31Ed
I1cPpYkr/DUoMyVAKcvxetFwFzR/Cqcsz5s801BqrxoACU/kXDYju4rOjSUBk0oSlPeXaHubN4x8
WCoR9kdaAvOYYr6umTjzU8UclQJk5iz7g7Si4ovbi6Bm1Kg0/esWOjznDoIpZTH2yHTRjZzwPb4J
HrRvWxUIQUwOl/kOr09oUcKQqm77LUxedU1T8F9jaaocKWd7CjLxcZ5cn4d+ZZgaIcYQ8+/zfBW+
EGXjQrRZnngeKY8o8zeRfS/IBvM6lBvVNcMK9PhYGy41c0MTc6kTVAQj4IIcUK/Tb3mPJJkn8shv
au8homSjUyPiQ4PrwHTdM7Ta1+VDergPH7uKkRPteeUIG83tvvKNkZdDk02aK2NNr9wjWnsfv/q5
mUThuNngnZ7GRR3hiovuYM1Pk8+/0dcV+ASA0C3kL5ZWX10rB/2HIoEYTfwVbyKSEWTAl1jjLvrM
SP6HwlQIjICCASERan5wG9D1Sl0Ca08Fq18uppXovRdz1WBVf0ZZY3YLUyjVk4WpSlgPar03KRlS
FWqmwcdauPD5koIEC2FWEPTPJLzVvqnHuPbcDdxwTLclNrOEgquE+w7L3szYcq0JPmKefQJs3Awl
WZFASVN+YxyYuCbt1VxLnz4DD4F8Y2cH55NsTwQqevhKY5Yi1Keu3JsgoCZSnRw/RweR9hw2f9ga
YvkNAsN4wSgQ0Wc3V3TcJQWco0i49DpsfxwPVeM8Iv/QR8qiXFkpPGcb4G8so3/7oxQeSuqBx/6M
yXeEX8tTWVrrTI2qLPBl63P5cuuIBQz5eLyXXAMVWPLqVYlZAfvBnY95fougcgFT3B010RkrIbxK
rucBeKf04CVLFd7dQHqSBZtoSvBfEckaiLLc2VI3NLs5N5ENdMiMnQhEKwLkatq2qPQbfrmOtVC4
tvKslOm0KQhMlCkEtiRaueY9yVpSmB+B8PR0jNbXQUDg10ER3RJHdg/u43DCCAxtfa2uBXDAZTfY
/O7Y8y9eAH2YyvPlNWUQr1IA0x5E1T6frq3Z5ar/7BgMq3r/kH1PWEIl1pLkggfVA8gTV9OdgPi9
G50bWj99ufRvIAe1cKLAeYhaI47pZ0uGGsXMRMC0/r1urQGOhE+ebzlenvnAoP1ydJHB/2UoDWwC
E86qnt+rgueaLSKNG904GZbgMVZ148UZZ3fQ1ni5C+91D2CEFna+Ed6GWS0HsDVYV7YVFqcfm5EJ
pvoUBAW2L+GvGoQbyWcpT1XU5RsBTQ1ebTdBO8QQXHJP7TIzoY11km5P9O85SRDvHvYL+kDVgvw5
d3Xfe+IFMa1LHxdUCjr+k9PkjomLQp8b9uMikN0hlAJtsi6Jh9sMZap50gGxq/nV1yMpPGC85IuV
wS4PX9w4sbJfoi+CWHw+/3qDtncecpwq1NMT4v9vkkPcQOKf30projg3rUxxbf24isP9K0+PK7hm
LLFsaIlhqcpRawVLRkGE+Mf3Jn9rJJESceE5WuH7YOnfz5A5sPLKIH5P9Twg1rnzlsyB/1nQl8w7
k0fDqVsgBZ/hiSj72nL/Th51L7+oNPxsFsb5+lTw6jj4ATWSIYLfeQeW0B1xmTz3FpNKWo3dC+iB
DV/ddFd0jZ1/yFJ3A6e6l7stKo2x9Kri3j5seE5r/pH2T6ZPrpO0fdSK30VJHFEEZxfH5dtKsQ0x
CN74fJf/QSU+V1KAxR6aTjPrvYWSrG8VHJGJxIAsbTEf91wa8KXErYin80AuKS2N/unZHunxhPYV
fX3/BIDy8UQjRzsjFECkSC+8WbIWI4FKgKxdT/ReouibZ72VUHFT4GTR2V6fH79vfERPx5x9SwLN
curb7lqTR8QCXPlB4okOEDq1uhODwFj/6hw530b0b13MmjAgh6hQ7IM/n4/ZqaIuI0MLVQLPIClG
6ZURgWhGPKDWK1zFC7T+TD0Uk3Sd38Be/IPKWEf7WPD8NbNGxjXlKMPMlmvaMMm5rU2kQs41KKST
P4jPRL0AK2j00ICN4YzBRBZweYArO5dIRReCZuZXALsxrUkSUBDD8POMmDVKIMTude2gWkGr0JqA
oiXPv5ljmE1MztTyo5Jxsx4/2dy7ghxkGFSd2+oiC0lVUv4Z+ZBIczVbwSkun6oy8FZ9KTFzQnAY
D5dFxcrBmJJCDTGSM9JMfzy7kFKtaPgxoDsnabEWDTEFieUZYGT8XeUsesXvAS8q0B7sqqmFZyNH
NxSa+xTY2nGTU/4p95ZsO4Z2B+JXCEHAeLZbSUzcPBwOOHz966K55IADxGidyLDW0bJ6eqK6HL45
zh8PFHq3o5FDiHaPghc1gO7X3fSG7PGrWEJS3FASZM3gs5CJOhwzNoKm8/AgAf2wfjR63YO6E5BK
xCH70MUx2fYKUIFZwJmM+Vk7GnYJ2ecQJZ4BzvB5RWRFf4O0LvtJWW8Z2XN9GDmfqw4hIiBWQ5Qk
utXWXCgNpDUZEus6i0zPPsC7QcWfW1nkeBnG1mv98Jiizd7bPY2jnoPXBex0GUpsYhQfmEnb1xxa
mk/AZ1oApzceNylO07q29qFohUOo9cO0eaJxhIxFjvrPNTsJUMOVtpBHfnrgD6cXd0bLBc+3BWKQ
lTF9ja1YXyTUctb8mkjyHMFFW8vvmjnfaNgtG2V4VKk9DSLD5iShZ69g1TT3fu3F1/zIQ96U4DRp
T/CIKKMbiwUAENQSYrLSBAkVTWJK1q6iJnyIj1IbaBcv3Z3qjM6Zsw+XTmeX8kCBGzhbUnAjFVpF
2vFNm8+sdTTRbP/8rFZLElFSq67fdOOr86YB817yOqFCPfFTGJaC2hR/9mKXSrYEOcZloKQonnDB
GSleyJSKQW7Ai6ZSdJkmZ9J+xb4Qw66OVwQddns+7FRM4G2ZyE4lrGYF7UaWWBvM3nGz1MGnIIdW
uDMzUh7aoM8FA9seNVBjDskWaM7DzUMPsR8nUW7FfKOjto+qNO3yDqhR7UJHK3HHxvElY+EW7ALz
tVIT14Dn5LNHbzj0CL6skmTvha2e/jfC92D3nfGfPP5LfTaV51Js5NckMQEwN1ckM8f0WNIJMwaT
bqK7ZFe89aZYXCgXY363Q5B/YUSi1OaRB/gcyKVCAkBRTkeSmX3Nu6NKzhHfi3+YXLgn1mSMhW0U
JZSGCV3PccsePzjnqBfrnSDFNHEWlKKpGUr1FwtVO/nGF7Klv5SpPe42gXJjexKNFptcLqvA6DUU
cjOgfRAvhzoyGy4ydCFaZ5SHhasR6zGjKiAodlkCLAxg93YGcCAxOck2aNNXl6f6pqchCCEAgGHI
vsdUhOsvNRMgf3RffXyS09WTmY/DA/xc0YN2WGUCe40xmTghyAj6pNBhLQhVTMKFG0u4bIDs1Y4s
zT4j43PDKTNkG8tdNgQrzDroz2CpnUAZLh5+ugB7J8HctS/9BQgFg60J9a8GjClh/U+2RsJTENi1
AiNf1icKPDHH9qT7aqt/FL6OqJd2YgxF0KIOgdabsgjIAqSXx54K+0lCzSE1Tw7b1v7YS/pOheMH
SU3GU91/+73/VEJkm6+92fxfPl2/MNfyDAhZ0w7Y0Qa3rv/24unRWphhxaxsq75sEXBj5dEQHvkg
zK5rL5+x7MbjOGah8ZM99Uxge+Xhif6+TwUff1Y6OpT6AXg6KvO8kqGbistI1gdP9y1Weec6ETZq
C1MW5MXSUL3X2RDrV1k8AJyqLG8MvvSGwDw7DXlSRsSutp2G9apryPat5k5swX+fl3GP0e65m8X9
8lIdICWYu5/taqE6jyvj3GrGG+NK4qs+g/2W/I6HqyKAVv5HqgIBb80Fje7794RkbuoN9G1aZfHH
ggcnVIt5dRVcgzI6dR0VKq7uS2fyJqdHKnwMq5aE3ZOUkC71kBi4/46eUntaUSbRVLJbLIGOf8gk
vnUgoZjg3FAB6LyrHqTWGkBNA/U8HPcOTf9Oi0g4LoxmpxezcAMySUiRR7SlcXCMF7UnE1Th9xX+
WuZAknLeP6fvDi0MJBPblRzhwQ5diLr+7Ku27ZFg1wYMk2Z+k7M/XRo+m3zmvAJb4c2RZm+oqG+a
8jQyQrbw/yaxFcEIZnomrT5WjTZ1U4i2pyRN1tFaAolq2IGkf17pgpMr7HdHtoiUTbfseRpbBWP1
2DX1SAXmuJ1QZ13BJF/occ9vIR06mmWgKp9PIuMwTyFp3qA07glIsFSk8qd7yvytPCwdeHjrDrnV
aDbAUAWwgsuLRoflCMwfd1mY3jKrsMIKxhpGFgJz9mhzCBr9FaK//gIL6fP/IAMOW4XUScUoBDV0
uJY0kBjKba9B3oWeVqe8MRDzMm2fMiZf0oNF1Df8Lj0U99CQ4Dw26YZH637Mscf10oUQVE0jZsSJ
6qMa5BRsOVjczF5wHOsWIGSQg93PH8OD0NadRVLDxTT5+MetkgqxDYRFmjt68K44nezYItnYZovL
VSFBAsjZuthlsbgdSHIt94k9ftT0nAJTjNoiYVN7yxcgsf74Nj212wUxgkDU5uCMStkhmFAuj2g7
aK/xlU+zX3Rcf/nD19BoD77r5X+G87wiiKJX8B3JaECv1CUHFjP4Xl5H/uLrD8+iImmt7jMLNepl
kjNFFsmgRMgn8yKEWnV6ghPe10eXI1CDFIBWmAYuYcvqhGobmbnoxMCbAixsm4QWvxH9x5qD8+Po
JXeA3CIXp6Arnn9oNT+ReegL8VFVpKXPzKkpR6q0GrsZNTajrqn5ubnEn8l++na0SEvHmJdH+mlF
jnTXSAhFa6LCQaDh8E6yap3z5xpeTQGNm+5bImpcAIIovwUYW8d8JTPb0mWpZLAMvhw+1xbtVeGP
p19jbXTE/R2xtK6my44qB7nj1eUteS2v7ig3cg5kppvJ39uep2vbPffcXvWWDlI9YD+FxLhtOeOg
1l/l82dkb4dUBHcqYD4xeuBMhcWlWCEcrLeYsPkjq0dwibRCJ/gmjkrERsjah+wWj2QuCY3T0ME8
l5OM7OQpo/5MzT4Re1loeFj9Sg8459ZPORV7GdAojggxE/VFNmlQ7coLZwUCCSSffzLEPV8xeilb
fivr6qtarNF0tYJXz9HKC4dYGvxmG+3asj6X/36BQ6CosPSh7tp0D0i7/A1eRyYn/daN7NgeuXRu
Y8cL1YXWultFANceHO/aIVBIuU7bC88Mdv1Yj2PA2NHOFVcjmTPPaYASF4hByrbwpxJy1lgPsq7l
wB3jM4EzfKryQKjrQ1mD+JA28GRpOqYheSZxs0K2Rz8frGzmDgELTQb6DJy8MhdpiHZcHFQ3v6wY
nh1mJaW/SlNzvvzWvolWrfpwSirjM7skv+gZUDfq1RHYqoee6K8vZIt98eWefShywmlVikcmupr0
BgRHskzZE0jJBESFdLyv52XGz/DT+Z/zrOUEQJrF7ch7xnj5Ja4I7rTQUjxvQHt/G7B6Bom3vGkN
wH78y66C2QJNIbxLDEaNbgHgyPuKRXL3vWlGmurludJ77pdwS2e1GRhjp1wT4ULYIAPJODlmFJSb
LHAKNUBS/eo6vb8ql3eCDGk26cWF+cla05SU3LFkSmBNC84Ozl8rf9nvAdr9GQRSVQjPCmgWa0Ms
GjHhA0D6t2kYlUa/t3mQ0McEPoVuMHmyoaKPGrOqO5LKXIEQbiouA/EBPfrPSqjNLKdWac/tbWQX
/wnxDvExmcZItdsyFJGLNZD3SW5xGg2VDd/wIdiLhLqTbDwG5Q214462Y6yOPfzAFZ3u32YF/GOF
0Sq1K9SUjB5N6mGcJMYJF2KrlRabEAIouQHzqRFQ+DfY4RuEgqFVr/Y2F+BQDaaJfRsz4gtzUtn8
WN6R6bJMLspKHM5qaxBqmx48RDKUS6hK9tXDWexFlWq4gooA0f6cRAx3PZEkBFMbzLLFYzIulPCC
L1sZnq+PXMb49DaSuF29MHZSGncj13Tc5QXS3OaeoPDzb2R+RmxW8xpV3061no4P9suC66ltOuhB
o1daIMaPjO0f8D8qLiWjX/OXu2L3n5FUv5OQakMd75jq2doFxzsN9nEV6rscfY+EJJa0l51TtB6O
Gvfvh9bDBA51eyhZpMPh9HVedPYYf7/Jrnmt2OrT+R/mMNg456pzYl+j97r1fDChn2u7N4xSdQDU
QIlpm8lmuk6YZGUk3YQY6bZhyxzoG+Fs1yZWwG7VDODZ8FhKqneKsgNz0tSLIcTLoxOQMA0dgj0D
HIfTQ28QL42i4BuMRtCaWZcfYiGt3JLW4n2j5sZEGSxnBdvMMfWHDm7nNtjGWf0D1FcrfmQ0u1yB
BMTJw7JiWJ+D1X0fX8oH8NWiO2C0XqvHYh1em2RSAbKyP7U+VOV7VHMzhsuJx6gkqQpSBz3wd6zP
hudfSnsveLH7LdDjxaGwCo1PGb1pEV+6LaAJcE9Tvh4mL94keyncIVrExxANWRzQcGMv091j3eCH
P6rWg/a3bGmQzFOrxqe4qQsKaK+vWNZZs/2Ehlfe29Bpzgnouwv4S7Po3OpFbFPwMfhlmjab0Msq
Iemlc92JMuit1rqKRQg+DoxOJmh9WaIr3ASu/dHxHwJRV02I8cVUzWe4JsotwikWilMqwibAB+pO
ze13HRhp99moL7ONs2/bTETXBlKaOrHBwv1LliqyP/IFsCpWfctaGut33UXWqn9/14WcxtwPhevh
egh0ok6yj1x4JYBLl9Dw9+90SwAorSAoffGaFuBvvKOmZAVLQvxh+xOHPOlbEoqYC+Rwr7+X705c
9rOB2y9Tqdymj6++AEdyA6drVGwSAXDNR+hMmqvRPvk4JyUKUXZtl7RCr/HTFoORNeNuoRQ8gXRE
EK4Vx2BR/nG4ADyQl74tlADyFZl5uj19WMSAhQHD/oESMOG0AXzZAZOvzvFzgsWNGCWNiMiUF7da
XaWqVq9JRz+40taUCNGf1Ezt/AL2FBfDrO076Bsbh8byYKMJhvpDpqkhJOwTtjRa0ZagYj8hlSLI
U4YI9ZWKLUToMkWW1AO51cQhTH9NqbyoKBn4VQ36WrPci0URFKszLtTDXHs4eyq6J7YXMrLykBGP
QnzU4MU+Eo9h5bjOc3az5yET+FAKUDQjYIVTvgmcbwRWBqGUTd+4xJhJOHoJXmPFKc2zVMwJ2+HI
9My5XbyJQH4e7HkeyxLvVmGp0kmOYawp7v69/+jE8z5etNzBKbeL3lQMy3wnXdODMoOijK7ZrhiU
jCPijASnbSk20WBjHPIQCkXkkYxWch15Pqr5Jy6E5t+j2F9ryJTVWMxNQnMLjzTdv4qMqQwlyyZn
slk9SJAfeBqDKLGkVnFgci1w0vKQ4cHBg3P6FNJUY72cUEwuJLA/DcpJRoixIrVzt3SsyBUUfJHX
J4FKAUXP8r2mBvX7bH6r9RVSKPcYhGnulDoJDzI3uyo/Y+DefzDtXCSe21Cw8G1fi0dqdnpydNDb
4Pl9vtWwlJR9GUXI/21P/cvXQ7qkaW2dOHHo5d9FuzFzuu2sPubUcOABeGWe4m8d2fNFeDKTcMSd
td0hAIvSsehKS3oOGOtAeAJJKFmGVl92xmWh71UaYtxUl4imkfuSMBg5BdS05xVMG5NOLQkO2UaJ
TiQKrRKVtk+/ZP8N9GvfDC+dfsSB2G9BCo1u5ntlsCD3yWS3bmebkK32lPouWRAB2zq1y4e72EH0
kw7i0Y2qOXtqSJQSn7VZglXahNEHE7sxTOJPkjnupp6MqqhkVQtdiJ5XAtowxOHyZTRbNhhkYrmY
qnOP4gO0I9hcmpp9EQ400fO7IB1fowmf44PgruHR13o9Hcv1+aCSR324Fmv0OcM10Dgaz8DtUDqt
PciFCSIiW5btY3BcsfsS9sOBQMmMbjnBU6iXWB98KFq8Du6nLXMLiCXrzxLiaA4WK1mZVzqtK/ow
GZ17bDq8GD7QGbA6rO3tPXQEXQh/7Y6+vztUa0S+79WsbokAlc7zQMuz7PWQx9EnRIuBDm8FOXPF
3RsA4KCoRFyZ2jaOTpr06fYDV3l2YlOB9o3wPy+aHf7sWv+/ufrlySaGYOPyrlO7zC96gzOaZJLP
rJ5nrQt5x3AribFdQQjyISMJ59R/cRstrVt8YZi61fbaeZLAmhoee4U0ZI2KGOlkZcf9zj47sTzu
zQWPIq19jmr/ggaIA6/GyKy8ixosxQfejQTSHaYtDmfBf+CeSX149kt067Wc1HlQR+5mFgAKdBmj
EVboDZZUa4t3y+3RD6phusunygJKlhcvyUu8P7jq550gn6eFmapeo/ZLMqDw3k+Dwvjc59lyB3uG
yhFaHaLoG6lKUM7CFTlY14XeUHseTEMktZT7KHk6pqYNBEnEJz25znxMMi/T1UxCHIIFHBpBwyTM
1BOff6DrRcHv82zZuYK3/guJ8pZ7iXq/sw11knBf6niT6C7P6HIuUbI3M5KDKDsgLyc8HxsZmQdQ
GMRHTvO6XtNEHiLp/Gh/tz0xXWRIp21u/vJFiHfNOeQyiMDlINtHzaLYTw8UHyRuLTpvI8mPiBVJ
gR6uJZq2ekJiog3mvVvwrB9GnnTRlnXTLDjTbkKViGFsy96IdAgVoAlI/5H/iwT4/SWWrNgGt+GU
2Cr5VG6FGOlLQakALWFDUMsKyAzeMH6Zx/33cLtCiJVpR2as+xwS+K2WjqJV1zt387MOzgAd9RUn
SODj6UQJ8zZtpA/fkKeRrTTKk374ws/dLnyY/j5tsQHvRJeY72CdcpNWa3gyh6F4n/Z+SRzrki4e
gKVBlNMmAYpABiZwXPkf5JjtkeJmVv/XRiu+P8COPRhkAbpGjYpqnkWaF2Dwtkz66dCSpYlJuHVo
Vmj+8/Bdg6wi82wwpl22FttOSPvn3tJctvEyyd7TAFm1vaUcW1bTxf0qJp5w7tixX6CmxGEOZSV5
SYTB3X1Iyw9NLS716RJjwH1lJbN6X7hS+4QGLRy7xbHLCpK8oXiuh6p4GypqArdGV9gnG5W2xbbi
cdqJ9KhgPvuU/Okk2HoKhJ2ugHAbiQSPV6Cssr7sSeO3R4OUJjVM19WlHZ/8iayxi142d6ibdeiL
3x7WgCBn7zHDVebslivMTiWG2qKkzYhUUHrhDjggVGGETj9Lp35GlwAu+6J/yyu71LfFSnamfHEJ
mdYP0P8R+L88gnu2Q76tMCdoSV0e+SJElPXURTNQCGzlazXPWA5016PH27DUfnIWo8bbCEEYhdZb
4+CUjJN/1XMpT1mpztGcHsRBP+qiPVjKNk7vhfKGe+CM0WMkcbVDQ7ggs1/cqoDrcq5E5chkl82G
N3S30RDf1YK4ceYelQV5YInF69qlQxglTX9G37TfPG+efbInzqOwr0qRV7yxVdB8oXijrGWeuv/e
8I1X3zjGtPhlA3na7VDjZFqkPOdCtEK9d4H/fLk58JhMxxUsQd/4/2ORN9zOPv9yaKJYXnSYWOOc
RPSOgv3+epyReS12Uh0lLms3rzm1Wa+e4RPq0joT3iUXR/3Sjvln8vd6C4RVd16Ik0Gxljlxuh/3
y/Cq1hnF9UKgsnWqv+Ni+gg/OB/emeHpCoJH+NANHkYMGbE8qfwR6E4CbyNRpNWNQg4gheVCatde
ssVSwAqolv5lZol5gRkJ0GBNFtKeQIwm4Cwsz4ICa8qii0maoteKj4UQtU0BjevGTMA1jNgCds8F
LvqrIYrUL0BRdlnpFtGrMQ/ydMZhNG09Flwt4xLtZfLHOSNTMyh+sPh2+UUhLgzCw1/NEn9OQ7KS
ORWcW6y4IOWeMhgHOAoOjRnGFFLB/fTIlw9AUSqMtLA+mbyne7gGS9LJrD9mJBY5GN1OBFv29DE4
Ne9nNBJfUdfjfB/zzJjR9J3ZxKqlsTXf7QP32RC80m8lZ1GwR2JGnAp4ulGKdAV7XgglcXetUZb7
pe8166+6qLCX9ig5ajneFZ4EPkNSxGxSxBFVN5NdgsQh3EyX7/lbT2uzQt88xuYHPQnAr54HgD+l
6VccQO3I9Hnifvxz3Yu+BTBj3CwYQs0z+297CxJVxzOzTm2kh69YaWl93+yO1D/ZlxJk9q50Ij2r
VfnZyQIiSSNf0hSo4XilP4n80UDfslZrUbb6SAXafdTXSaJ/z4sV9B+NZHACBi6177K4H6zuAM0C
Lb//+yt0Dj/lbv7hd4hbpNqSM0t35J3fXqS6+r23L9zqW3sZJ91+KMcHrS6tKwRvqADDa6pAi1TX
YfsafCk9pVK7KFrNzKR2ZBXWEZItNzOem+MCXbFGlcGhVCp//syzMYdR1uunPfImDWEwvC7VEJok
lxOfe5u+K5lSIFbphu+KGJmEAlCh9xjjHlsQBxMIGbiskWP6YdJ5bETOytE8cJddIXCAVJUQvb7h
gHy6joz4KGpKSTHOTxazsnDFqwRznjxJ6A9HhBQk1hYudSiFPfndJukE0gnm0jpa0hI3ZyHDPXXi
m/ZHPqEB8bVHnsdNJWhG3dduhhTdIhsO50LuN/kH/FguMQa5kdotwyzQb6xB4QQ62vR0gOCH3J2f
Mk5u1LDNGFPc4aCNcnBuQwYhrehcaLepF6a0djsOCTck7OnnnNiXITkpJxQ7AB+0XZCmqNmwKLGX
cp1w5ebvf3MjRY/YeVT+dD7/s6e3PTEWCjIlflrn4/IlKGRKY/pBV5oX5q3V+EjdkOAdS16FyqYX
NE75r4BBdktql6fvs4rejk9tXP2i1VC21ylynhkY8QWuhuGn8ckY2Qd+SjbCavbYVbwIhPU3Drd4
W11J4aVE7juOJsBJhJA60q38HZg5YGsyLxqSlQaEFXW0IuIzAwXo88elZqCmmXoG7/Sq/bNhS093
vsrX2Imjcix5tFngjVV2m3wU8k0fKztL0NcK4GAJMoxKzyWvmor3YCwriC8OhufXoa+2Xph3fsVS
z/IWwxp7634iA4aT4Uv1VhpAtMLIoxdDTs7Rs+eeFFwbEX7xBeY3gG/vs6zPLYeHvvrVDfeQNxZH
qiCV68HyH9BwSFr0f/mrmS/zqkRlcZLhVV3r/+TXHw/xk7lgr3H/abduTd2M1zLVugbFFaNmgUFY
KtYkvDPAtfpVeFnxgiqZwdQRvtcxzC4VsfSswRzuSEiXOjLqJxZHu3Lz05IAj9Xz1/tv5eWsvLzY
zcvKkLD9opnzGUzQsD8r7NZso9MDHHylDryEdI8GaUb+j+GWDWiiUQidfqPbmWtUneUdtQfxNkPY
xVT2xV4/JFrY542cseNnpp4yBRZNGWGWOAIpOwgXmggEQk0OJJAi9OYSWzXV5+jJy6hk/ow+Syx2
MIU8IiS7bQq2LkbHXVoLRw6go0GS+BXtS7vQfZtKJI7Qcok3qCdyRmv+rMBpNUG2fq5AOaz6aJBI
/juHEari/JtMlrdauDSdOg/8sUS5tLN0VLFkKDbEYTVVNuKbSPykcyqUkyReYyDiuoJIRVOkhQIP
ORZuazkRnjv0l43QBksWnX0LpTYy1ziZBFIHhHpWmKgDyJdDk2tZflFKy+K5VJjDf3ORz+HtGRQb
WZslta+dB0HK/Sd7tZget9mSQP7Jin0cQxLPr1xhCqMbdg/wpPFsQxTd6PiY4sqxqQjGwtWcGgY7
IpRdqxsr48cr6WGI0MKfq/ac8jMIDPuTaLrh7s6vPkk2IMkjtnvqSqqCkD/h7U90DT4TWslg8uO1
Rgmc4gO1CRPU6zf/1vg6OmS9nXE/3IQKbENZucNdLZRPHWmYnMb+wPX+TX+JBlkhyMPYWWyZC+Nl
LbrAovGTk6VRWxbkCxMOi1iJT6GC4QwRddB2GjZj+iiw0I8UddQN+MsIu4aMOQBYML7Tdw5ij4Mg
mG0ZVTgLrScnX7eMkx88yTy2FGMATvEZ39hSEcnITw6VyIK7+njYOw4unKVk/psFgnu7elx/HAsw
xFYoRv17Agrz8+vLfwp3B/W2RMc0qthrusO7EXGWBQF/oVe4SKgFRvlnEFK10Jugi1QlbMzo17FR
ed81D52tT1dM6RECNk1gIMsz2akBeJs8c85CWUNoJO8mvSOesUfFdnk1XqhxUSzrzmXdC6Bg1vU6
XKGVDGqcFWNcSYq6K2nFIVt84P1dApTy35CYRQ5gRX81Lk2AnV7fbY9B0qkggzEHHNcivlRV854F
sqUN5lAxCUmrxpW3o5Vn9mzB6WbTMJPEGj59hHJPG99u6GOxcCn8EOEIqtdoWb/ug+ore1GhC5hA
A8Oa29ito0WAlYJjlXogOUKNG3kIULYvDJCDyvhxfc2IlMmGipAfvykTKZY46nQFt0t/50TnRn7r
NhsvUqbL4+lpl92GVz7klg+lr0GVYBCw/wXw3JNVfQeYTGjjy/+DhK9AJIFCVpOOaNVgc100Cjt3
dVq7qajQECG0YrbIX9BQyGHjoBqeMqVsAvEUEMK8kd+QVO9z0rCBW1fW85nobqZnRGM6GgyTOXVD
JMwO/LCvBCjzVeaFuwDjL3PDwBq6HYZ9XgXJyEYBfvUffcC+0obmeR64p47K7ki/vFv39WjkC1vN
L+kka3zEqglU+f2PbeG5hcFNN5AMa2jGnruWZSt1E5AJY90820MNenBKfM6d0v5JA+KygP6AlFMu
h71sQtOia0Q1jh7EZVXXTfLj49ZDA5DHj3v2n3uOPD4v+Phz3sossQxJ77H54K1CK9LunF8Nbbke
uNFZJCzGDkTJFvbjRz1UJJFccYtU5MeM+qYTq4fvtXNMtwmEUwnuFVv08mbIBtJJkeixWu+qGOux
cubHQqszpUE7Ne/jOiGDzJl/cyTuRm0eypp3ZfsbF7OGdbCfRollNSb/kySJLbbdy1zcR3On5yNR
OPMUOJVfzR6iYQv80MdzFhbBUGQgh2oYrRyHshH3FUMDa1/Y3FTc2uY2EWgcMDl0HT/RRTiBUR8d
HBwTyWevi/32qTK0wwKflVyg7eG/s9iEKDg9y1S0ugLKjNe/lW1pGjMPo96IxdnXc/mEUgvZziMY
hH38SJmCBydfLawAZR7IxelUOHzOQoCURymM7IuZ4knZ8a3vv8HJ2LbDDxpsDHIVlClfLHU4/RnS
oi9yBVLuYtplWdWMl20H57Eu1pWtUn+fpOQHBLpF9H1U4shHU6PwYmL1QmWZQdA4ilicADsVjdhL
ku9vM8cxHyQDXErXm3xHXTWjRuqSfXOWCEzzbRdTkI8/gBI9s+qTnDdsatHIgHkSHn7b861nsjfg
iwi/LgTBav5yy8WJVmNhKrIeCA1F8SX3mSTyGD4+3u/Q6SlVQZKuYsrGKkYL4u7bh8M+z8BNmQAL
IqHwmoVrGFmsICFj+Rdmxq/qv12NvGio2o2XYWmWlEqp0oajjLcMMCu3b6wP1a1/48q2a4Blsww/
+jhmetEuYf/+vdvlEqJhvrNvBcFnW0zBtrjWFs2ETGHLAjRBgtQ+CWPekPpT/YWNV44tiSyvt/yH
r8azy2wJn9DOVUTnLrrpyEaOeFp5ac7fYz2IMJpi0QUir4BHDlGLXYBfXPFO6ltw3qSQFJl8Fxys
vkOB20mb3uJDuRZ8Run9JVjqxtNV5bTyDLzJI1B/GFUo3WTnD8+EPXdhKOKHw8ZNCFciJ0P9z+oZ
JF/Uv3fngESsg/UmSYDEyVBKH8gQePHK7IwXSzDT9+CgzdaZrZx6TZGjrn0Blau4Zd5si0NYDlxF
LwtoHBLS4iDBc4CQPMRs9f2lHXFaP9zUgh0/v5Ap93DsmCFV3mbQen3640AHjsopldPaAsitqlZ3
zXF9jwxoOaDmtX9HSfPKhwTqIn55+DwkIhvtvs19u0LuDxJMRQdF7ne97oHVZ5coKttgj7Lmkorm
GYypwwIaZRiVt3e+U8swI5RHGCuwe+/F2Sv36c/KY5hGaaDnFA0VFYBnmTB6GtVfSHF9IQQdGV5s
2N/6Czu3QUifndSZr/2blOm3WPIV4d+JWGyWqRjDwYvxbDbrQ6wTc3aul9VcJOYDy06Duq7n8PfT
NRaI+K/43yG0N7ocxK5dZ5kWxoJEiySSHgxLEuPAZ2QeD2YVH6Ivffcp4YYdX/VjwlSDwufMxzla
mFHEyyswkQILzKzCuO1ljcQHnOwDrUp31Udd0bTCwSHLtabcMJ77h91eQUUVSsZnuPNiRszF3G73
6QfarR05VhVhEgAfzg611nsduLA4Ue1lx8yX0HnzuO3DCiRCZa5gy72n94knVI3yzMumBzqMdaWM
AdqPUyj1Z8veIwC+coUc7AzP2+WkJWFsM9NbkqG7gcD9YS49CNtRTMNbyWdG9KEJRrZfBk2hcN7V
kb5/BsQ5IJcxLrlWBous8kpwuhWkEU0ddWw12K/nSoH4ux+qHB+xDdK7yYPpSHProHUz/LAaJ47R
NP7rk4kUpol00jtvbXPv4hIekTunsmjqaFqQ8uwh7LDQVYKtvwoZy/4U10Oazvyh0cj5pILxBrNC
lfj8Poea8jqaAvacL82AQ6NU/P6cJNxGpfor9IuDd1etlR4UbB3xYw50vZ1R9KQLqy9LFJ7D+wM0
6jkXWCVgy0I0AYq1axWPUHv4cWP6i7RJZ1jtwyqYRkhfVhK9igg9uCtMHXc4Bmf9hTTUfomEr5CY
OA7qXhS7gk92QjS1+aAjDdWR1HVi8K3y8ndcgrH2B0F9eERgp45xklEnOw8u3SBY2tcchuYG4BJm
N4+s9NASxcFGZjzWCBRR2hlbYR3LsBCEXXeZSFRQMyLlt0uFVDo8EWTg+ZdD8WUMNJhKKvgXqmjw
jxR1KoJs1FGMrRkUcc1j7lkY7ftRTWv26McFggQqxG1pIwBQYvooGQAGh4H0dlUv/aQizWXqciK5
fSwCYxlS6F8pwHC82ax019WhXbzkIn5Pdv68J+KRNOWtGfsnehbiwIu8B4V0tEG9Efkjauc/qESi
GClxGwaVbQbrMB/ZXRTSjy7utgZnq0KWMimIFHoF33/Ezvc2+VZKK9jFtsjXSAgIHSCsI9nBa6A4
jvIriQ3/K8LvGwXIqOLJeGxezjM1NAUj7Fe0AXwbb29IvGEkZ23iuy7olPbyjud095AW5c3lURyT
cWmvDkLFtHVKzTnig99NtBJKTzUHyNRC8y0TSUODkGy56NSxg/x4n5ZgVmw8ympTZErfzwpgfROc
PoRDZY1P/zS6JeHOLBzgAbN8/LjtVivxZlMJOkUYkUROFfi77XX/kfYQFbTiWUQxWl4yc5DH8No9
ajyq5Jd4FbE1YBHywp3qDdiNVTBuFPs24U20sh2R31SNtQHKEs9zM6rD6xI2YhLI5BNDwF5a7Jfm
+nIlviERIOngd8eRoX5WGGVjipEA+UM8awBR1+RXhu/Kfbso30NbzDjGM7Vb8rTRGysiIse+gVmh
UEptLfuqpEKE5xT8morFUFDKHgW1tSoeJ1bzvbgxAxq+EmA2T98Akq/4n8QBjfLa3gxuBG8XHLxs
NziEodaEWzolQvbTGJ/VBwf+IANHlK1vHOGowUaJY1MvCHuiQOc8e2kjPWevdyn2I6P410mz7QaO
vCg/roTJV6k4Rkno0MVVI6xgQJSuAQ7QO19xRIPaK94pJ4pSC2BM+dEEOvMg8NxQ9y76VZpmAs43
LJl1GbQmAgiG4Ij+Tcy18uIyJbuJDTzidkb5ZhviK+uNmUsGFbbXy1VpbhQyyfJ3JkQFDiYzSrWw
H7RtN0hJkGPJFab7oKvdXQroSnHCYj4hmV72wd5cwWakPMiFl9TYXWqu2o3YSZkKHf2LulJxTGaT
qicGSln+5twxuivESufl7jsPA10BfBaHbgPTY0GTUI+hcWsKKnBpEpadZaQcK8fJ68FKTBrXmR1E
cdHOR95jnyfiV2GdF3X8RzCnwuYQdF6S+UK1AbcB+HAm3PV4Z+ejIQE5ErNarLiVtasnSmqGes42
gZaXyWTl6NW5NwJ50vXo2hvCNHJxK4uh2fWUoqV3Ql2u3k2QvU6bYa/h9fZeOxU1CQ3jxPrNog9G
mr3aN07mr6FGhI50OfvU3SomtwbqwQrUFcRfbpknZEEBt7pOdgiCnXyDUX3MXs7N++T/oq6XXaxm
EJXt7uuQCwGkVKrTjSnaOj/1gaWlgywF43J9P8y14uD73eUbtKnJNHyl6Qq+ARPZ/13f20bazKJR
HslqsgA42joJcdbE4keAjEj9mudg+vbaB18oQDGcOZfuJPCXDYgOci/4e3AAlKVCEWrY96XEg1AW
2KQef0V7tR8ZW0dJWOjaHvcfB9pAGbIfJdY0daCqv4st4kFGlsQei6M6US1wuf4OSAX6yERrgrsq
jtiDbKdNW6fjHqHgFEuDyQnlmyR5HFucGKkNlK7bXD+AT7gYVzupMVLbeIMDwrKDcswY7quR774L
ct9C8AURSfS/N80ITEO2HRjc3PhAdlxktFnq/V/uSoXf/iAw3ReRay6+auDsqTcyIUeCjO+e2UsM
eXdHSq+sIwhawiRE4msFcquLWdO0ydfAk6l8FbHXlFw/gmgrFHWti6bbWUW70WjQ7FQh8PvF5jPl
fzkyVPYkHCeuySLTsXARmNC4hPr76gHL2IkVO7GeN29LyruD0uRuov1G9Kx7MCxa8uBpUk3lm4IN
2dJb2ACVum/GomAmfBUGdBdTCSsHh7gaptb7Ys750IaZfuvnkTgrPCQ7/UZzuMF0lSTN+/fp4j9n
u0PJWZq7gBAnicD8JhDkCsZQLP4zq2U6lbp4d/+GEJm7mVi8scIAzaTygxm7xJuweMgIfQlTyU1a
NRpBaq01a7E3PfGugh2R/JcfKId7rhLc0KZH5Ni8wG/Ec7THj5+GbnyMDH93eXPpetsakd75QvIn
AdivnbKm7ri2gP1LILFcVNUfz93//ujQdsrtkgXnGiGDkI+FPVkkPT8cu/f8Glo1qtMNkGGK7jFE
YU2PoOzOqOlbKc8i0TyaSiMPV8qNZIExC0FcNi3qz+gKsbEP6V9+ckrUeK9Pi7Q5L8P9UbI+N7fT
/SS5+nh7cW1fHfO4PomkaYV0wo6+wf+NvaSefflQhJT2TYyFYRwDdgC3K2Gky54vHd3HE78HvKrw
8Vgqk3xrt9h7qa0a4vkTMOI+UNyI7J8QR1B7pgn8SOHdnrwFPOcgOGGf1yI06HbgwyVV8nLN3/k1
ckR592SObXrUB3xkxOt6x3dw+FtHLoabw2AsDsi6jVKs/Jn/WeOqT5Yb9ceqnnjI/X5UFiAodTWT
BhFWH0emr2UA44tRm53lpTgf66+zqnxAVIq/Msjyt6XVbbWS5IinoTtg+IAimzi3zTvYhaMVei5t
B4qDwF9HtN06h2Gktfn95J0YkA/TAHk3KAo6olEaCIHjV+IsKHiDmFf4P3uRlFtuZj5Vhi4TIMYA
BGgcJvlLsZBkqPBte5iAyL2OEj+2F2AiQ7lH2b/SHnSHtM/e8RHBTjCUKfApoZtSC20Fm/9Exh/b
+8KpbTAoHncOTL/uFAx0f826V3iyQmkjis83Iza2L/sk+PpmfT2MtIUtW1iZn+zK1bKR3n1eWlmb
+8tkv65n94FeGi85M5w5fzYs465isfdpoj6N2w9bYZBMLx5TkHV/CjAXrcl1On7Z+VnseC3YrPXA
zym/ta6KlI1/TQSRpyLjnp+kQQ4hXaaDgKaJ3TpehK3y622Qm/ld57Js54wPHj/vJWLC3Rq4y1ow
PFntvWbhM/W1Ickw+dVjxisvtC+5jqIT5OAAzMrVgPFlP6pfqSpGlbTloo3lsNJ1XPvthtEMF4ak
0bY5pjaaekYjYaaMFPYi9cud5ip/mj9j/ja50Jv4AbhpX0Cm1YpXGBLfoEmdGEX0RCRry1oYgXqd
iLOXB9egxTX4CjHBoXr7q3FThD1cF2YdyBNVeY74zemTYGiqY3G/zeI0EX/XL8iqTcWyowu2UGBw
7FbulXPo2bT6a4+UqU3pKwl2By3kxnKXMscA9ujZ4ZZeQ0NlZgHtQ60EvUnMIPj9G19YGCQvrzGI
gY8o6SRQmR4xMIgOx0ujLfKi0eGAmNYuaavo/frByJ/+CmuhuIvLC4+qbszFLDhRDkdt6XJjZM5f
PIjhOR7gifrv9kKZofOwoAtwTes8/mgafATJnLuwMT4T8/bFpqpFQNhMaiD5hCR0mtKw2QL5JQor
MG1E5dzb3kSlPyJYHOOo6GkCGCjXG/sWq1Uu0vRx26ZK/638DGNhk7dyRInP0kE1ijsCndCpvt87
xmSCMyts7dsD8xdnLfzTTyBwjew3EVngvzsCKmVkuPra7/RuDtIRnZBqFIrZKQPo+MFdVNMJ5fFb
eUST7m/TaxhHPeQ5M6I5DsjW1VlpbkXRclYuughYI7TdWlQtJkG5pLwG+J+mvqbAs1aCr4M/c4O4
PUDbECyT8VLH1ufWgBVTS35yZlj+DWowU/3POm0iH8z8YGD5Wp95JvD6PGb6J3xPOk3j3B6BgOX9
XQYILfn6QSwa6repC1UMlFomuubRXNvucCqbLviMLa4nkuF779SAn6MdQ/eE1nYDMeNBjJPtVRZg
FZuj1AQvQTDnhiJX9iBiyI5eD+trQu2GedBGQzCwnCDYYtK+ZLYVlIUOltwTbUyVnv0ri96UUssz
snV0bLkuAO7y6fb+XLR9Q7wwJFdbx5e0EsQZ/G4+i5EyIO549VTOPY2lYKeO9YDvjxDy7vPdDpPZ
+NntxAnsCCxv/gJaAelEwk8LdgOuxeLX2rhN9R/X9VfoSuLQ47aw4fKnVss9iY317ouKMjltQsD0
EKZka2UVrTcm60/pZDDFDhZlbksOWfCho6jI/dr0b8ruH/snsgdAWBzEHu7bucs6+5bCoqEag09Q
6I9415OaSYg9hHaP7ssP/3AcK8HKxBvX5XL43s7/51UJOEbGXBm45qtRjZevPHfw1rqda5J48wsg
RU5vs6vpV+2piSA5CaSaRm54cQk4tVf7pBJaofEPDAnstFEIMjro7UNF5Ja9NfLeFvUpND8EYelz
H0oBtBP76LD1XpNea2SGQnZ8Hbr4fUsoBMUlwZCAJfrPilTq7NcSTSTVYiMacBht/SRa4n6sHM3o
6kX3HTB2JqYNi2M8UYjS4yYCv6zP0aalFEnB32xe+O0en3CMgurqHVPruCu8hfPKgTZD+38Rjo6A
jm3WScXKwI18yK0IZnYF455RZUd4nyeVWmTyqYWmU2lVAfLyWP5e85qNAsAxHLO9JcYIfy4FqofH
fXoUE64bwszE4bcJYng4+9ScrWuK0AUDc286h6KAwG6aupuIt+QXkcl+npxGvkmG9vlThQvbwM+C
P0UReuRLBnHyya+brl+ZJE6HTcSmkOI1N3WiF5ENAVgPPfAB4PTjnKRgAjtg17aiOJn2c2NesMMf
G7kpJ6kpZbM1uZmTh9j6zqersq5bJ/2NcSub8EwHsw4lRyP7LC2k6zk8C+U7PXcgnXUqz5pWN031
a4e1EuPyWXYmllUO3t1sf1Bd54mTKYfFg1es6EhdsMyJVOnclaCFIFRG9ivRTmSFFlCwQDrwoAZ1
3LHQ+hLIMkyT3lqO2ZyS+DLLNlqZlOTXaTjkVGZCXzmnBMlDDY2Q03ML5T4RSQ6k7Ojag1bNCANM
hbUAvjitooblVr7pb23wCZ48W+yZBYAD65DuUMeEKCE08fAp0YUq2tqJtN8u8soXGbK8351cw5ie
6kg9vGV5odJI6/nqCmeksurZ4MrF3J4rv5cvpY924XvW/aF46UmNnX2mIM3YaOYKApm83ADn4cjU
kjZh1N8NVcYVS2E7UW7PI869YEzWfp1pY5cUPUsI6d0Hq8d7X+4C0kRjTY4cGHFhRh32AujR6GJ9
MCiyJ7dx5obP81WDriopLxLtYZhw/96du2giEE55npJXC9kbOxlxosI0n3e1K5wQHp3UBJZIcRpa
LX3u84/Kj24cyeypeJa8HizX7bhBCbM1hqUDSjGDoUcySls8wMfIfsc2PqLnNBNOr47vHVDJDOEb
Pe7wouN7dB5kay9Gbc+t36PUqRbgtI0duVinYTWxgSKmrh375d78WGdT6SahC/ps0tZE091XVK4W
XKZjd1lxj1D2hKi64kJuLctP+dI0Do5arBgbF4E+jMx+SkKA7ob3xMa6yOled1j+QhOUcTPNUUVD
aKSLDHIrQZ/wng2GUFzYD/ilTQcv+vzGpQVaydmqV/PrXeb8r6XxrBQPrGFYlGZzFM3MKbr9Q9KJ
1YYKA0IcE9T1b8YLS1si8A/yp196dDC2Dsgu9LDj3x5X4l2kZNNSxNidIE85amYKRPQt7SQ14t1S
Wi8Zj3FPERWgWLnO1uuzQR4LSLEq+7JbiZdUekJrPUvSwcr0QGEImqb3j4wyXCoB87bt+WMoGL9C
8wncZy196Jd+tNd8UY0qnXZ69VL/GPJMWeBfoeKw3LOnrXUK03PF5f0SVz3mdVr82Mx5lfyvSdHF
WEESolO9LIP4PANpBZg5jZ4Rykjggm3avdkt4Iae5eQX2h+lHHK8Dva3URu1uAV+acn9tTmuRKHr
VRhzQl6Fp+DfjkIu0wQwb4nVkltPUZRdwY/PmGrkgC3o6cWCSwtdG2ejsjgiIrA7pdSLgXY2+hrD
ObwUo+FMmQoiosvNqGypOdt2Aa1ZcZLddHBynhtFmLWBrzjMfjtSsGyVxDz9SV8Y+v+is5IYWPdl
+rnkspMApNRwLnxUGFHHjcnhDnRJ99BZRfdoTcqhirIwEufrORICD1EcmnGelqgAF8+EJNLmpl1X
bQUbC6WKfZty4yKnCS8pBkjClRwAt09Jtf8uvLWqYsJ+7gi4iXXIYYN4ibtGGBO5Sm54XwN5Ob9v
awdwSoGwh8IV18vYRNLh9YvzgcEkpO5jkUdlJoZg0MiexSfW11tVdyFT3mZziKNYY3yl4nfQJEKa
twRdsUroUIylnEI/YonygGLYvAn0P1YzqJUkgEtRVjAB4+4fM/HRp+Mc9wFjigiREhM5LjK8xXGG
v6GB/HcGkYWxHlLWgscEL/YxtXh/IYV92DUKbvN55QXtlq/axPocbuVTQMlfY87V9lO9g5/k749P
9vUg57M0+ZO5u4xD0f0Rz90hPW45OX1VzV1xCxlUkoH4AWJXg2dIEFiYHBNKi1KLtw5dHqxFc05I
aRTv7iiFE8xnoExhGcv1s3TYnF5yMl0gpMPTwAVzFjakG95H5L8pMecvFTirrmXrrE8DKjPtGutk
/xkZ0MCMf+AOgmCeNet73UNWa7EWTUguPYLrvv4k+OB+G88+O1m3mjzWsN0DQrYwXnC4BWov75bG
/SwjAksCwCv+83ib+rCTCOSIYKEqaaEXeVfuVlO2x4u0O6ZUA/tNSEjFllmkCWDgbwmJ5hRtQkrh
eq0J6/cmxR2k98svnWr+PrOH1ByGgPq2aZmiFXIuIcVXE1ipcR0oM79wgaXeYixZoEK1jfRXhhTL
3voSdohlnK5zGEbI/S6Gv27IL6hDYC9PtIvpelJl/h3IJKk7vhDCzFMZvHjvj+tGN4NAQczVUJA6
MtWdDIRPx0S2kJ3za5a0lt8dPa6rIwfh6nHtadYOH0e56y3dqGPQyMwYgq6DVegOkFjGo3AzkSlb
5t+K4aK46jwgI332KVYMHd/hiHHEm3ItkKke81EWuIDMpL/A70BzyEq8WhHIQ+dlSav3PZjTGxV1
OY8ESEr/kivQ/QeM2Z667QtsBuOvnB6NYWRIwZ36jBb1YqXtMc+fmiYpx1y4MoDW3npPUBfsVg1k
/lg3lhK/zm7WXJ9unM9BMi0mRxQ/AaheDvM+6spdaMGhfjtUxhunh+kO8jxid79erVsDCwZEVF0X
+Z6ZcGRaPq2UoG675/yFIlpGQ/ersR5J1fZOyHywyO1zCQkkIbXyP6iYPNrUmxUUIi/lRoO2tFc0
vfx8i5D+Zdl19RBxxWODA+EAVjHIKSyJr0ft8O/KzPkgWMtitSFUm7nFiOhm1qPXD3wjpiTLuULs
V+D714sFN2u0BxVT8Vty17dbZzQCDXYrlBSVpbmsJW+Zum1qoUBvPPen5YYfLmbkokiqYvzhGhqR
rvbGi+YUp6fvH2s+GsDWPLqvgEuNBUAHYJjXBwKlO6cp/zd+4db1S9+052tkPJk5Dv/QUEpOq4QK
lh30zaUl/3C2f9w+65X8Qi3MleBZQ/+EAaT9vVkWEB0rAgYTe4z8L5bb1u4Nt4UHGQWNRpHidGL4
cJwTR4B3gFkZ2yi89Y5jqu+SrPGkiYfiX3Qti6EUCu9dlGVSJvAZi/CoFAm4a5s0MMrw4X2Yff3t
yrrKBLi0H2Hz2M/mtXpjjXycbnkYRQO9YSqrD1c1Y/7rpkKT3pMxnsFLXCETWhBRvBt5Hqkxuyzi
lOWZGKmPKWOYYCfWnsFsiuh+U/S+xgGI2xV8Arh7rHU62ZpISAbZeBWD9ByiQSHFlCDlESQOiwWx
0/4KlVx70rTFomNFI8aXDdOEz0GwRMAKdp3U9z8ccyu7s2hy3krswxmkXs67rToUJvdssfel/KcL
x9o5aDXlJNBLxCbv8+T3RYIzfgy2NC5FnvF2Zq7NQLAcCNoTZoq2/od6BNG3VH1Eg4ULbzXKjdKj
1qW4Ih2Yp8wp2mwgKr7k7NtKfD88dBk7qpYbUPpSFuEznkbmHBK51JoAvxuw614fUiTjuAygvuXa
hO6XLQvRD0ZBwf6xPh+YiZKH//S7xHsyNs6Q+JCuGUnclmojFRZ61eoapp+HSinuk5M2erJOG+Db
Yx9PbGwTA0vLOJbsSc++ZJiWDS0QRz0huTqnLYFimvqfoRmvSZrRdszFRiblK7ytWDpi6KuX3sVb
FbP6ks6b6oMb2DNqV/HekQ93afAF4uo19hB/IpcUnpjjImpzTVg5jW4xxuI4F2twC9B7XSCmjQMG
esEqiJqthfE/krL5qGR6r+y8hlDfsercyfb+qR08XvtAux8HI7KEYPmnPeDBBZJLe9bvdgUeK2J5
zCHv03x1oFnPznK+n0Nl1sZ0LyU8Ek+sPK+hmLIuYcJ1zSkGBBTboXB33lCXc68O7CJMfCnf8kZk
UIrUebIQa3XmBz1qi8aRP5O77QDwcx0YanjF+Jf4BwJEnTendA4B0mDDbypurl3hMsLulr2NJYI2
xdsi7AudTS4nAbrGQJXzStUVvQnmFYgIcL0ILZNnoR5CSySj/5X3A4ohV1xpVrXPnioEz0uev7lM
KPIELK2Ad4281IpgbMg/7IWA7JXb29BIbiph2Uhrz3yjlPXtdVz6E7KtCpwTwR+HJgDL0jVpIHGq
GmjO8qncjmRdH5vTmzMIskCJLPEUmST/SXoU1JIWDy36TBvUs2MGaRa9QS3sqVar6qEh4efh/mJd
GGk13BhmEX3GahNkA1qdwCENmdwLeAfVSGjt8BmGd0RcmBLhVaFn05om2IKRTqQFmhEfen39r2DF
PIExQ5CcrhREW/2iHqMUrZoDlBt/bHqmTTu5TN6Y6icNklKW4qaUNWkspcOF/N7tEeo6Bdk3OTgN
JkJEkeKbz8170h1duz6zCFRPdC+gSE/bBv61CxELLkfPH3L9Q3AqXUxQCCtV4OYubMpVqWIEKDHA
Z+cFvSCza+jeqSK5nO6VTBO0ATvu645yiuYeeUg1eTD86WuhsqbSXF+3V5l6sajjr2qRWYCdDTzs
nzFDJdVBJpUtoFVGb6E5Z9PZpDhARoprbq8FaE7UCY3jiXDk2d6AfsHUGN/4JTyAl+ZeHghn9q7P
8MUR3N9vrBPw8pMl4z8M1MpbRGIrgkp4enDU7en76CRW2wK1Gc0Pme3XbyVFpVbSZNKn79k7M+H+
ZQZydvlY9gQ+sgZrchfIL9f9f/Z5/92a2onmVpKyw0UmR7qp5AK67bRrR6CFxYqBho3CGo0NWmD1
KTmikvdKTSxNNEd54QLSv8jFvhQmD2QuYJQlrYiQ57mq+Ti3zuo9dfeRwnxqw851J1d++qh1JL4R
TNTyuOvMD9ZWLRmQfJSPcesTyjF/LBDgj5M+t9RWwwwSwOMcOlozlXT3cVEjF3kAd6qKRxTQ5CBK
P0sD9TN/HmfccW06neT2DP0zzp7Jmbtl+dbfDCO015wPUhrrluaFaB+vIzGt2LDwshy/VCJWhNLs
5xIaAvAGrWV+CeqhBLm+yP7SQ9mChnl4Oiut6pKf1xDJGV7LRwbhaJmqWBP+zYFY3zZo/6JugHB+
HIaq+VxBrbt0wbCX46QIE5XILFCHhjOH0YvJeaZ1R9FYNwcqwE31NLpm/Vstwa4XOVZZJBntxYGu
TkQdS6vpAgTu3sG6V+ansN9KyzghmcjzHeXvZ2bPJRZcfr+OCdnCpw73iCddw/F4OcuGeGnSzmys
wGHQW5Oh5oov8yX5OMzG+GOO3XtLr0N77d2vucr2Z5kDShiKDrY3bw3aRLt+hal5fhSHkTp3fWLL
EtfRNt/rxpKGDEcRxJGFXFG9qflWYdg4rjn6zxCIwBWIX34LDWBlqId26ZSi1JhD8qji6Qxo4Ftu
KV0KkqLrggGsyonwTavjrJZUtB7TUqqD1nNwNP23yoIl8sFc6JU/mm4KgnNdB4MgxWACsHSYwObY
Bn5p2tVJzl5k0HdKKIEj0TmmBqKijzxD7JkrqYJbvdsHqZVOuVT5R0JDi3zSBtmoYCJfr1GH7bD9
D5s/6HM4pKorRraDBiEm+PcZ7txs8cU8N62sMb7UiAIdSV/9JxBcd9atDHp8c+8eJymH/E3Gnfc4
20Uo+p6gURRWjiDg10QlDEe2Pte+XFipd+zdwEX5RvIZHDBUm6xRF9iqEpU9axuWaEhxv/qBoXYO
5veC4mDchhWNLAnAZCPgqy6cxvAUASKm2qvCg4a5HCb5R7tR05Jns2yEwksIAz4KuKLzcuYcKOni
5g/WByqdMQPM7WkHAAbthQei6pmKiBctFPR//VJPe9na9QwVSaOFs/xlHnJ6kX1xcy2WirZutEng
aHW9btwlXe446W8FTRH2NN9s7J9tEqV22Z/ZJl1oWzYyDZDv17FGAj2zjchGM6NImYIFWNrV/b3N
T5OnvLOeUXBSO11vc3fN51YA6Bv/0K7s+4xjD8Hv6GrZO8YbQ3jnQ2AHda/G+J3btsK4c5+o5m2p
SNjE2EhhuyZ8WZCbB8YPNb701SzrfmRQre8BWv6eeB8F4RxgNoYZktLrIr1KRzn3PM+mooq5JZCr
sL6zWATjSMC8xMS8Y2rcYx0HZfMEeQX2OayaMx1KJr3M90ooCPktXFX3IpgqO1TnSuXPOSTiUC8g
xoTi6hx9mMfJsSIBAw+89rj9skQRXabhoAXtI1m9gF+2eEtlaMSwLXvXM06iDdUp2kbX+ILrMAyK
PIUg6/OjXw3c2sHg/oOYopGBT5/f2G1GW/KVBUeYOmG+3bSBz6ekLdMPjGxUerwjStUGg7BmpI2p
wOhlh/IzjSswFOfYNYaQO1NgSDH998cjoZOW+klUnfWofGF4Y7la+jXz9sp8L4I5jfDJ3i1MmTel
s23Ls6VLbQFohueTiLDrIFJg+cjvxYZw20v+bGD3aL42t61+o5lGiDI+5qqKi3T+BhMJsc3Ta+D6
RvyvAlJ8PC+6/Al12MK06NLA3Ey4GkGapM1hYUfY8wBrDn4MnLXq3we0MGwAQm+UjAq/98Uo5SeY
HqevebqQK1PNf9TiwN7C091lWkxFrmVS5syn72cjOPryrvwdN1LbBaVQ+RQhzml0WUqXvw/W9LOo
XG0tGYTxM7ZIqQx8R1kLkjkeHCgiDU42vp6QHJrKq/U/qbibsj0FiS/DRBN+n0GnZayNnRQDIB5l
DNmhOx23xFAGEOTmOEYsnCiybcKMkYZ6jqkdvYHn+6ZuGCBGDqHH9LqsZcYWOIiqwLSmXn921YUx
Oged7XjMEjBdwGnqbIfxSgrko5YpYRr1ilPcLWH1oLHlF5BA0iGiIdcjCZ5ynH2v4db5fYuY11V1
TcLtPWjpJJHUXMlnQzs70xtTTJp2K2X/VUMuiYCKl2I/zlzF5ruilKWmoqbZjM59uI5sjd/pvAlz
DsjX1lEj+UBS6e9ePosH536na9sqg67WyH97NMQ1q3i4fSbF5AcRUizbtygcNgLQAsErMxCcNIWX
U2YYfRAxZLxYpszr6OCShqD2ERqUL2obI2ktBsv/C6zbYOwIrokBG/pp+5Dfaa4bRorIj012nUts
sToSIHsxk2ofm0MPSOWYLW5JFnj+W6k7S4FxiTXTFxRbC3e80CRZmYmVUIZ3m6a9WSzraJajWSWS
5ooAyVGzuYBDcsWslUDFwXehtqrS5BMM0D1HaW1VN+NtNK7abN5w6OxgTLa3sqi5XDqOA4g2pNJs
NDBCIdZnrjs3/UY/4xUeCjQGyMN+yaYafzmy7MjBGCE0F1qqZG3/6rp+ukTuT/dMF/UeqcM7Zkze
f+3ufEfDL3lciNz+E5XrushkPrrLLPDvflx661yX8/94uFQ2OrOYJth00DkxUZkM2Fes8AgeycCO
aT/oPzrfMI6InydiSQZwCfvAum7BCF9doEMXRNw66kgmhT46lYgO1CBBFvuZtD+ax3vsd3GqS8Do
ReP0DNyyzwQRw0k3Zfrw+cy2k0TjUdKKlFfBJnMTWObiG7OreXhUxDcFUbrr8LN+pZB7PnYcjduI
ItQUUap+qcUyn/PwqfDcxToj68Y1jV7K+Me1/hfBSQ/ZMk8QRQAToKVgiTb2eTCiISX+c4YdXdpO
SsQnorFyC0MixGR+l0pwnnO6N2l1qd6q4lnwlQVZKmdY3mFUotqfT95gS78m31AFP15ACoIUNVHW
ILL3Qk9its76IumuW3fnU2VO7hZY1/ui5qIZksaFy6/pzV+tgQ2yM09dOZGSWYY0P0lhDtXn6WTR
nUq7gl+HTupZP5TxZpKxiMK9SNNjm5xp5r4yw9FzohIUWLOxEsjaDlEkuaX5eUVHgo9f/4XYF22H
Nw/w0fXPKj6vaVx7NIWhvRcBynZKBW7W1PGIRiOxwBLyRqQ5eyyXeyFCzoIXXGWXZqp5AKDZlGG0
bi8bQ961xk99ACNIu9xyU1HOI3K0gsn2eUXBtUY1WBJI64Zvyh7dxXApo9GnguCTFOHM/FhAEBUC
6kbD04d4Klj2q+fHPPl08qsCJyBF1aSNKcgHkzE5t6v6WdW6XWN3RDjtiHKKOxetBV9DOPoxWeqA
cW2QFPu8pKNUs2oixjAuIi+FaeD3GA4XCu7GtE/JeMtNntj/N/YcxRC3zx593V68kjoHtIY1S+7P
IlbuAvKxtpF+k9O+5ztjRvOa5vXdFuaU48O2HfHePh0wIaoAZIa5oFJemExdd8CmAzp2BtTcb8I4
gESNapFyS7XlXQCcA9H8uFmaGQZebxiJ5Y/0FFNZSP5RkYCd8nb4U0GydwpQComjx+wsoSlj1TRY
arMsDbkwhcl/BS4w6XM/b8pTizx/oFRRvesbuiNsd8rYEZ8dDhrWOykUNJJcpgZOxXXbaub4mtLv
5aC2vRpq2CYuMWD+3qNhNUzfV1TWtHWbtI1G/Ed3tFyF6alzn+pcPNAK0p4pddXZ/hufbRdvflSd
yPe+WI16tAcOTMg5U8qp2PVV1SwzPEySM8nlOMQ4QdVj1feoZjQmviidVhmtbho6R+/7277+OFhI
B/a1FSrWpwlED9pUeHibJ3zFbsE+HuOHVz0MZRhB+TrKR+1RQafWJMYn3xuyPRAfg9e1MsknoAN0
mApZw9+soWdjREdullnN4yXfnVH+DcnBO2Hynv2MDJTT5qOjQ4AcTFFv/FczMjGa/g6ScULfG0J4
yYQx8JLdg0+E1lU0+QDX/dYzdSjYPcJ4VHTuGdPp8u4+YbLFEWwflpgLdE5+sXGjtf5XBpxtUnd4
+Q2RpCy+K1ecMBjv8xslLk+CtDdnUV5CN04h2cSbAU0ZkmCHaAat3z6q5tcJABk/YdEe5Iic65Ej
GE5eHsUa+7/0m86clpTh0SiwlEOB//TOSez9+K9C/lFvQSopVYvMK9601Llm2CWgVTZs3g2rUMtl
vHWtLGeuj7DiZoKpK5iCKa0x1XPP3w4EXqef8h0jGT0JwNR4bCgtN54eINcECI+ZO6kjv0FVkNhT
20jbiW3WUjTZMnS2HZh12TXHq6Dj36t+MpLPUT3tDAIS1tjtLw9zVD05FZXwvuc9v1+xaYA91U9t
4s7kfVEhuTH3tHkxpaPXy34x1N4JvLej3rt9V9rLuZMtFIqKTrOU5Ekt6dQtz8VcahL3/33RouPR
gtd02nmmBElcvQWD8J/dp7IEbU3lneWoX2IUfsVBKIB2RzWSVr51whybpuLRx6KCN6nM+Vqr1yva
kTyy3XLr5zR6wtG59/FwmjsvqFuLO/EFvFCAhfT6U3D4OuLpx7cFkCPzVVWj6tcn5POe4XbuqZ84
1ixZTcGEldWqPRgJBtd2QmxqFDRz2o0aAQVb5Ed16YhtfVYknekZw95CL2DTH2R5XY2pvvv4pNTB
vmlkHJ0+BiqXEMAxf34rZICDsFjzB65YrwJLtcvC/S+ppIT9OxMvZd2fv1J84Et969SK1SH2fCu9
4b757nNWjLneOMgVzC/Ds66dUt665lXXmRNoThuDQQTPEM5289pwEEfKzBWxpGv7AwUh4YV9UPik
jd7udJ+lK8MFO0mx2tAfQPJvDnqPQVBTonesN98UszsS4BKhcdqXULk9nbrnH3kow2vCY/ovWsbL
A4xgMq7jwAQDQLRYdoZ8Tha5ycwizKIC2170wKOtpWW0pY7RcJE/58pkzkw7tyAhNYCKPsiYIxoq
SnZt6fwu8qcBGGc8vXx0tWpe/FvZOm0LCFIAAaobYWwlTu0celVqXq1KHpo97g5C7WzUCUNOPHw4
ADwQHPD8JxdlRBNI6MD1eWzaZpNgwVdahvVmnW0clMHHRReoRwDfUVe9sxqqKcTd2veZ/S7xl3uo
Ph85pwYCfunrhcV0OAhWX5wtm6kLFiySlqBk+JG94XXx5xH+GJHShvm6zsMbrKwNAPbbYye7/rbT
pjte0U6WtOqpRUNERh0z5J+PniZNFrVIjqyzbROQFe5aO5uM+e/bcvQqFR+O/cFUWefiePhMtpT/
C3KaW354pMQOyANGUsVc+jC6KOaN6S+q+F8PpSIMhxWV47Y5wu0Ow0uRfmGSeXAMGnVN+JKM6aPk
UNNWDIES/M0dP3eSKvLdCsFKSPYsRypzsgtLF9E9gtJiBtRYeUoRJG8bvpkfqDvIqJWIVIK1p6J3
UdfCn2kpwvFD/7AzZcxyEKPOL6JL8MeEN2t+JyHCOX6KhPvb90/RAnvbMXZ6E+jlYxohyhR86bmS
+6rfaEPMT1v53v8dv/OqtOSBLoj2tZM0eUZqrdUiANz/tM/ZaRSxpmBHsIQPetlP+1lpyfXvTEgM
AtKjAZanAzuuTPMkxmeIYQ21fJHWHEiiScdbeboj2nijfluqqY65RilIZqij//W88KohBgm5IJ8S
4UB/i2dlxH7sPVhg+Huh2iIxqmBZjINgUfRdep0i9NOfFGI78bWW4BnmB8xzckAYB7gHxYhdxZVD
IGFFrYYUqORz+YwwXAUNm+O0RUh4vV/To3z0Ou+JIvVEZB5Sibu97sZmES9EtZSA5B+vNRLrw4C+
5t/KJPxNgKO4N0YsZa1btbchEXxr0d+7ItXLeV/qLP8XgyTjOI8kOx3OhOnUho8P+0XR+1JnnFlR
Es9+By4tfUxWrwdYgBUteg+f+n9QvPL/CTNHtkKc8AbZufMcXiHla6O3KfqgU2qZ+1xbEdoYesNQ
aggMlzZDJUQr+ZCESxye/IhgFBL2VBioPgWnMt6Ranj61rgfBkU2IseMmTos8wiQpB6G52WWYADT
MJNdprG6boCFCVzFAcaRcIB05CxNBu6liJOJCI6WthPm4n/JJE07uqrnttSAuVTklChAxvJNQicO
S35jg+ru/LG5RyMwsTHrO1e/wHblkRrGZ34kErMMNnK/mqKLeNV4UzmKaBTfTWd0I3di5nvs6wd8
QfqGh6RZG9cSIZ2gERFQ816/bk5XeMvYikofaHvWlLZHahRssIoH7n3YeZd5P6XIxhY8CWqKPeNf
9fBJJcAZ3yut+XK/32H08MRVIoHJ7UozgukN2xxiAdU7BnyXlfEfvdCCdAfFiYMZOel/C18jeC0P
YeQs2XoNmnxmBQ+dZ4SxiyfQ/1nAULezXOcMo5FKX9PFHE26S7Xr7kETvNrfH3oCkUZwTxtYTFg0
uw7gdu6zx6SGU7M14es38OIFrJD49MAi8AHAZnyZijSx2e8iab88nhlp6v0GCUn0bEYmsD+XNhML
Jc996c94bnlxCQSUwPTm3yh84rXR4cIy693bAEkV4G/UycfU3AxcwgyFKQdymKFKlT612B9aeJwl
Wh9/kx38PIUssiiHMRC4unyDwS8f47vLtyK3s8xc7S++3n+RmTMs+BZgYKYrKl194Q5VHu46nhfN
L93pefg+z0dR8A6vqgih4VFr2fkHikUUtCK8dnsbfMFEDnQm67mNyKp9pWILGBQ6103HgeUI6Kyv
VJgDvjAnkrl7YrIe9qElOyfCGT9qmOs9MP6YrA9Lcu2TZRQcdhACFji20R4HhdjIGLJeNJMbZs4j
cvzBj150mnLbRMyZscTcJBXUgywC+gXzZjWwlcumHR0t+W89wNlGizIt7CEWnSdxZ2O0Kc+PCb6+
+SMtTBdleOdFleceH25+FzqlvuQ3MzyzbrdZERVH3vZytsyGso0M50ckBY29tGKl74luf0wR/VoM
TgZ/X5lJXhkMuUmgftwm4kS1RiamyePrfFFRy6eXUKegN4XFKtQa+jdzvJvm6/RhJ2xKnvyjUWBq
ATWGYSO5M2Far31hB5XyGfpRsrcUhM3j8Avns5hcRbN78iCQ/tdI7eGYp/ITUyo4hT5xp3m/vveS
8G5UV34WTGVa5w11Nr4mNP/w4zjxgGXW7AdBvhB/acOLnmreb6+DK0zsFtug8RDAtG0BNvOuUVv/
jrXlA66kjhsVGyREuHxIiTbq+U8wb+ETMS9/ZFw4Dyo3GpsBlJB+w3C5nekGo8nxTNAwNBVjzeKl
xW5SDN3Fb3kVJQ4bYO17d01nWP91nQXvw2dB8ZCi/XrUa+WuhvPGeTsOWD7qvxmivvumHkJv1Jde
Tx3ZakHellRjdOBAmETZGVe+7zIxcZo5/p7jQuJgAEEnPGCZ2sqHdJjI+32W0RCRmgh/eN0IQd85
RZSA0pQbFlo5a1M83P5JjJoUhEb12mWl9h3PYlQ99EqbNknGHGqlQE9o/gP6cqWiqYL8xQwJ6yAK
0HVZQdtO3V/ovfMmT/EGcTTGcASs5AFpB/ePwHIv6tGWKhuBpSCqjEHpmD6ctsC3Y5rcRLltOb5b
vz6ipJs11sSKWYNvtx8dO9A+vSCiPQ5O/XhPoU08Xce4tRF8IBinHz2gpCLwzPsWeOBj3Len9hRR
Wy5YeqVMsRecEhzAPVnB2Pc80M8YBMI5hf/QXqLO9UogVgf/N8xUCQmNNOJiv2d/KdA6sNSPSdCc
s+/Z6z02lp4YFOUE6YZxtPTUMba1uoMtATZxdEleYZO2LWViIFjjOo2KcQnXHmi3mZJnWOdKxgQr
Op8V1UCgmjZ2JDzHyGUhvrLfNQoLWo/fAqvwqQrtuCF2y0Jkv7ZMDBpPjG7KDel10WsAjkyZtjK/
cWdWa0gddMTgtmAdxOWhdoY/ZoHG3eoNQqoRWi/dMWv36F91P9YEb7mH11HpOXSOs9iJS60PLycD
Cp9q0r0yfjet9hKsPF2sv2DJpSO1op4A5FAO3sF6LNyL8vjfyRazqMICSUzpQsaY/7HbQmLGGBXo
Az9eUTt9RiV/+OiG488allDHuHFvtzANYYViivgSph3RQ7T0m3GF+vGQvzwuEssjNDMll8GNa2k8
DTc5C4KYqohUnY4jgDNAV34Ca3CVdfOMbgZBweFKymTZRxMbHCtTqfK1IyIqQbfbKJXt9XEmX9rW
HlNsbB/8sBI1DYnYHqpC4NfjzvUPqAJOND1B8l1vFPiQjq3Gmn0u6t879STjabR3mK1utffuTl1K
Mk05LUMx9VXqZm5uin65bC7iYlU7IY4U/ME0PvmUtdJ6h5XS+bPeomGB8TtiHOJtnTWVbjIX7Nk2
HuvpwNi9/ps+TKlKmR7iZ/QS1XE5uZjyBbGmXSn6BsQmjJJHIwSevkmD+f0qkeej4/QcAno8xPOb
T86BKpaLSmXvauSHXs5K/kqfH9foPug0yi+thZFTdlvJAkkEayy8gsEShOthAEQ7begoR/2cITyg
UVEUmZGo80fuOOuQvD8UFxPU7cFY8VZR3NAH+8MbS/6VZjLcGhZhrKk1lbgBxjCAhUYviJP8nppU
KQlNjIZJzNswILYPX2aC4/M0T8P+EpChf90VYb4ZO8FL9tlyhyE0CE66qcQqF5r4/MRt5aDnWJCO
yNACqr8YFnBhdgkNtqK3iCrqLo1VZ/WPDzgVUKwAS9sruyF/DFy73KSlQDzKIftF34AW/S5iqLFz
TNRxcNMyTIBWCAoFOqxXxLYZYTangL45EJoRUAugXSj6hrexKYg7LP5YCiikpjOGhLb0kiwGxGqG
aOgNaQpDbxkkOEchCKdOon6C0Byqu837adtjNbHW0ScIk3rff8/CWfh0I20YMqy1LZ903DXmZI94
cPsY228375wwkQU0rkQzG1Ybsz0GB8i2vq0/2MldugXLkH7oVt4gYuUthNzTHD+6+vSxjLtz0QBS
rL8YMlH8KHevfRsQHpWSMXnOW3uD85JgX1EnMp6o9pCHvZrb9zhxEP1BwHyupPqPncOO+qnfasCX
ZUaJpe8wi1uWI2RxYMnitqQ7cgt8QEzUcrGXAhyn0PoURmUGLNvseg7AFi9gTxnkPHCYGauyjT/8
+KbeJYoKvJcn2XFE5+7CYMA2I6TykD9AFgQltD7bmoyzfI9c17wJ/1KSNAS/6LOypIa2s4vGKG14
QA9TcT4VG9CbrQCyEX3kBbuVVdDKfmP5dUQuLWhEpO2phgHbvd+kcXyn9H266ZaXn6nbFPi41rfi
6TJaSB40z1IiMj42EQi2gmykcyjEjOzVfChcNv0guCPLptFyH32kOGL5do6MtdEVr1okxlGlBXFK
jhZeUXR1Bd60s4hi4nXexM817q/l6781vtUetRse5y9h8L8ynsSuLNwcg+iwvk6CriV2AIl7oOJp
Ugfh0sV/pznxqV+lzLKamDTXqiipbcb2nKPy9pNIGCGzKFNhfJbCM744RO7iId4J1B2yd8jO45qX
LaXyh1QB00T8TrLpk97SMaSTBySD/weHZEXokIfLSPId2EYR8tcDuKCV5814wRlSDb5KFvZ/ON3n
8BID8ojrXGi1sNcIVgK2+87HpP/7q89lqeEDTuBQ2BNm/dloxaukjj0A4RxSPZNklMhJgWvopd1n
XjxzuOTAsxmH+zbZeMeNpqJlSMqmVnq4uOiYPMUZUDU9t5H1zf0/mKRkVGWR4HDrKrk6bTgRf/Mc
rlRbm7jH0tHPZuOD6WjsK36GMDhGBYq3sdSSF983rNhvijU/n5kG9uR2UdCwlPA0oFxkSUvEAc/3
80oFxMoIwebsd8SONd7WxAMO0D2TWApuhPIrrASSwp/gXePkcBiuxlrgTBp3fUVDNiBddECYqKiM
wbZT9kCCFpWd83yDsO/uXpck1pK4hXqm32Fyoyh0EIxwBBShKgq11PPiYk6cJNoFCnnZMghdCmSN
40E72VvhuXizRGkT4v1YsZPI0Lz8sOXw+tWnvKjMuIinuu6UOcygdN96paqBlNqNlXKSWfoK/KjY
7dfL2RujjN0i9G0HvHpW0EgtBFmPD0J2rx62wp4i1Ks2fFxHs+f9JUob+upgPjcrU5Z81vrb9R8l
AnxSv0GiuHqqSZvU/KsIwl4lymWREBiaEUdukhQbWH+may6rdvMNyDzjapD9cftMZgIsVk3MkLBG
Ye6piyYuvW8tYUFGk7KpgqcmL2wiFqeNxqJROgMj49P4rKQlHFzHhzs37KFnCbbk+sNU5G5H+TkA
pfyH+rAFOccznaBwRtQKY0sxXDLsE57tUP+pGSw+DZWfC6hVofxBGtSgIRZmlsB08HoK2z5AE4SC
JfpN60IIUTNlYxz1+2mGV+HqZyIX6ZLnJZwm/q3rjegJKvKagOfFdJqoGHjuPZKbODb1507Udkkc
43UHAFoiJcC+xZGSVAAb9p00fyHqbNnH2CP764ENq4A/iY51l80LdtL6jp9ZI4sHQwU1UaUJzLS5
L3THbWd/Zmt++X7C8HinP9kCPjaErfn4RBG0FA/x8pdzZmMEWyGuWsYl+BClC0PYM+nEGSq/1Hyc
CmNQvHOwmBMTNlSkSMPengw2JWTVQIeupNxix5l03iY1nnC38ts/Y7znj3idcuAtWEOucdHBkyU1
vI8va3OHjenU3sDKKhRw0Z1aiot2k87Fdo0qmNn3Ypi48xlkAVSkLt6jBtQYbH9GAcQPZ9Benj+E
+ZtqPl5tymf8HdNK1CSzpghmi5QcXPD5EWmD4I971ruNYFvk1TeChnT8GgMMAl5nuY1jCtUO2s9Q
dYjHcTinht6ZP132jpPU7GXybUdmM3HkegVQOJBR4eh3OhQqgCPKaGk6SU8JVbm29j5NgfpSxnRH
Xky9KRuDKzj+eQiWn1NVN4p3Q39IzhQ1sLyAhCX849fsBwMtyKiKP3+zdClG0MSU7P5fnT9qwkzj
9wbec5fTvkkbe7WFYYJINCis7wTf4sLFZ+POJcf/Jq//UgvgOXVqqueVN+i7nxlj/L4qpf00DHJx
iblzwM3z5Sp4RZkRGTz5R+EY8BvP+rKbrrClPeyDT/Pa87g3sKA1WAL3MjBx/AgDXQSMEsbSGN6m
SR7Rt+TtE/cfAzNluDkwVF4O//jA/LzYChOMg86jxfc1Y9SbC9nAs7a/2t93Fpv8I3NXBUz8A+qe
BeLjHPWGJYZz5EtBvwxjFQWuCMcAYk1Vsf2krqSpBPENOye5D8B+6/b3LJHvuZVAJDEy66NvFbei
JW0e7T/NPS5he4B5sHve2rWnMhKdTKtlGQliGeroRXf2esV1ZyTJU+COecwU/xsN7/Me22Xl9iL9
hAbBYGRFMBAx5iWlrrs3m4c1Kj/yg1aY5mCJ/vTLAtVeMe1qt7y+QdvT4NNkTp9JWHWTBmY6eI5q
T1gUxH//4+kZpgKUdl6PAULJSjcuyl1WDgTKmgzvVg6beJ5fPjLkWwrCi8NawKE+AFJbd1WsBiAo
OkfQSjTpNZsC4wd/bCkXvJUaSfucVU5hMkW0j+X+ChKsLRmNMd7+eoZUXNWdRqRYSLyCoDyTN6QP
v6EDBhJx0pr+eQoQkosmUejdujbgiMRJQmgwgmN9ys2fDScK/qT/MkFvAd7V6V5SqqDUae6/yjKG
PKX0HBNObe4xBhdtb2LsC8Dy4QNlLxQejnseYhe6K3bS+cvI7dYm4tsTJfi55Fg0Yk3MvMmIhjFH
4IrBSy79T9F+p5WK2ZL9N0aVeXfgwCxW7clMfACV/KtSqxVqbB6Z+ewyqAPtEaIlFf3gPtGxQR1f
X0YuifLPXNXePJp225MztNtFk8P5vwuTNRyfxpij1z7FDgCu5Ud5Hbz75lJMLp3lfFOKHfmmLOEq
F4/osf+kY2sBK0pz6UtgUFkkCIqF1Vk9EhztUzfLERjnHFC7AKpS9vANwtf6uieNFKdY49zCHfoO
4eS7T10lo1ndonF5z84OgpptuhhM4LcnbbSOT6oMm50z6ZNKs2VPheRpj8fYcfII/kRu+wbX+Gxi
o1V6r+RhteuERmxFGio+36otKFT+Es+2L1gPEJLsC2Nxp28VqUyBNY3/PTYiD3Z10PbvTeIYRczc
p+Bum/V9mGlpkJHQ1WX2XGENVuwqS+e3ajvlU3oQiskgMJac6y90wfBn2h5hALuTd0V52SPFHM5D
+pc949R7vZqcuHlbr8lCRVRbbQw3/ojNYtUmHqAE8KpHkkhFwqWs5CFqvq3Ms6Pu+sXt1TumWToq
o+cI8d2zu8w2a57ATrADnH4WKOeao3lUhj5R2RWgpVVIaH8uBjzpTKQ9AwU370ClTkPnQAQjYcXV
xOdAwJG5VHdBHN42860S+ZKEPjFdeAhiILUTgllNdWWIMgPvNx6I7xfMewD3Gfyj1skkZXctg7Hm
8B8EEfeEdddY32G7kG3b6ZCQteZt7GNThgYXYQBZnuC6myvJ9KQhRNSbWi4omKl/olJxb3wsyqD9
bmNcVWb3LDvFi121TjtW/SGNefpYaEdXTIEN4Cb6fVSZck1tlfFrSQ4tzr7gteTqlyVELBlj3COT
g5p74HmU4InyreHT3+sCeabDiQbGYpTEntuwh0j7+ncxAsneiH/Zs/NwKig5VaKQzD73mn99o5UK
mPV3+ZA9/Bj3UFXDf1ZtGMcCDbxfVKpH9FlcG1f8A1i3LYF14G4sW4pztMXhObeGhqSdes+jQ8OZ
OHh0DgXltrhwZpWhHEGmOe6dxS7eDyvDSKlpZ+DLqpH7ZDN7CmvOyckXA3ZIpehjGa2Mgus7M/ic
aWt11LP2pkZ6Z/tdu4NLbUO6yU/Yd7Ox7zcxzaYWg63a0WO3/RTZ2vCiFg1YcXBad0Lme0MwqgVl
uBHJl8ZfQF7YGl/OtwsqPmeFCLHM9GMqs+JAnzMQRn/LCBwGH+XhmxpVzaTM9RkSb6Rbuza7rwHB
W6Cs93mcTWOcXtyhFlxG+BlI29c4POx922e6U9/ZR7Dxl+prHI4lMTL3FD2Gt4IRMmyetd5/9g4o
mpEbA73p6HcvYNPiBFmzWCSuy/HIq+30SikfwGmhMbgz/6HLHFJ+OO8ItrM5WTfS1lmRvB1q8enc
9SbPne2OU/Iq1TPnCF07/i5qEslBBTk68OWrvb+f3FAzl0uKFZI81j6/Dge+Dl9XC5McPD+zHIXB
AG7LFdMuwPIpcdB5uCBO1MnQIYNnLhe/+CA5Yv/1whiNw8JaiSmf5qxfi/Ejd1w71oOmfV5CV+6J
uTjVXfpcb5KzJxCA09XmBj9jF7deq/uOUlyQRA8iOGeD7WoSjdz7hLoXtTSDlcTU2KIUxQs2Gm5U
d4FDYBtGxTJiK7x/HUlm2arHnw4anDuHEvSA9dAwpLfcV+6jJcAN15n08zoZYZE3AOUob6Tucys2
TxBunj/wW95NvwNkG3Zi0Ny26mj3IHKGt3uc8Lm60H8UIjAuA/pdjhvt8aZ2zkEBVozDfNP3dFEi
aSkerTnUI7WAHfmDIM05fvgV26N6rW7Z5xrmw//71s63KXJz8XcbS7iSUs16HCakHi7pcYiQUahT
ZmBJLypEpEklI9dexr9L5bMh6csRmYVhH7IC9SEH1eKSzXfUApzm5LNdGzgyS1tMvRDcuG9NerBl
s9zHyGOcQiCFYDZn7NbfZdXLqD3jlhyZpdN/BJxwhq8XIMb9czMG0XW+N3M/7S7xT1NjB4t8sff8
Roi1uG9JGEUjVOfqCmMVID6ZorycliSNrIwVZEYM0OFpO4ixktatbpeFYzZtC8rta8aO1rdGRhEM
up0FQuuhUnLj7gGVY5jQIiUbqEMu49HZ4Jygk67gc4tzgOzoiC2+bNp30Lx8mveAVws0tR5j1sOQ
Y+jJaQXDKg5tOhEqlUfJOIcxcM1333KjBYLCdqSJq1Y5tCoWqO5kFLUPt1LSb3LaUkJ1hICBs6A3
dWsoxMHD6uRPMNX88WgFK+7+BhzyDTLKoypmAuyq+DrZpnjO01SUNKvl34qik+YSk1ZqQSkjcIUq
Q28084cPESMKJUHHk5xOD2jiV40gDxE++dEn8QNnhc5piAScYxbsqrwScVhqpnSMjaC3l+HxLvLp
4Khv0niRIfENdu5nQRIWBR0D+yGig4bb6vhMWStU9Jl+KBIC3eWC8WyfQ6K6I7u2EIGs1fm04/Yu
HzJNFCPrnL2nD3JY+3y3DWh+YzDRbbI6lJOyMfOadLrXnboB+rXmymEVnsqW649qm3+g1l8fQ788
s39IO6tD1WX2BNKJOT1xTdKSEQU9SSlCXnfnuFuOlJXCBsxlaillJWA46kZu6M6DnT8QzOR8+2e9
DQeJsoJpvM7FSmCltbnB5yf1ipxo1EwNVuBEsKUIcacRCrOsWNYxRThbbQ5JpqclGIph9Huq3SD2
Y08h522bSYIxvpmcN3brSU+OMIXf0horwo6lagigrucln0BZ2b+/1E0jRT3aq7CmaghBBbB06ZeU
PCETEMCJb47q5+/9O9rmcows4/LRtaMLmvVfaIHF2e4w9YJVgP+hpK8llVhbgbW33nIq+2M3jJCz
3j/LzQofYUYSn0cw8jfd+KVcBoJWUudZJlvmVDb6leakMHVrjj7m7BKvPUJYHIWVxTudECI5JlaW
yLphzmWeAL7bm+G8cUKGdarwehVs+5ISVswEF+xCp2ZXgXaYmWaJsbelmnLh/DFNFLkYCZXwSwwj
4QTQGRe2pnidxTqvWSqpYo4R9xt0P+xzoM24Z3WtnzyAXLMY84+7p1MUPW23Y+44zywux+ep+cql
oj9GjTC+WMY9NhjX3DP3kYpdoby+dNL47fpKsQFhmbZVvHx3y63ufLqCJ7OgzUAEX3h1ElkhIj+v
ORae+pBOUh9gU7OuE7ivjSx1KDW5mLFLUZyI0u3ZKZqnXkz4+sPoT0SAJQjIpAEQdKuX87zp9UzD
JufroxeHpJwcWJCvKAi7DZXGgzzl0O0UzGxbxltNRfU6jmziy9qGrTMWh1DeEIFQaZdCkWhylri+
N+gwX16chK4ARIMBIiaPIar/ltyFMOBnpjXaiVDvL8Yj5EBkn3BIzUTrt/0F3vaB0rZFvbYhfm5e
vAHcV1B+ulniVV7pfZsF57JOgnk4+YS8Sj5kcl5iSrzw8H0Z+K5sheaXpenpd7P39W+m9BOrAoqg
qig7V0lyL76zES7AIokywWXHCvg43FKSWWwNmUqN13+7kPEAzewjUruPZ+AT1w9sXjE5huQ03jyy
Z5QGJAISIAdV5D81xPIoteKs8TXW+LQtnanZMESivfjhkOtJ9Q1B5+z8ATzdlX0IjBRscIslQzAQ
m7+8cO45gQ/DPKEMwvzt7M/kyw5A21kIrHIoFtyCUOa9u/YyasavM34wQ27bFeFQlUi5+TqbXq3P
cK1/cla5puRRn+uJpTpZr8YQG6C0Hdix7V+tyFiWthmqyeipry7es/fnrN3YisHKkihYyrEUOPCo
OXhXT4cDPkIyUtcaQ3o/zpvbe91gxljDh0wZSjtipv9j8zcuU7rGiuP1XcIihS6Bx3DQ2gK7rAFI
CwnS9IkpyvieW6xkQBum+q4v8gXiHpR27lF0/s9QPXtCrHrVlIbyQt5jGj+56pGeN/vuMPBCFSUC
h0BiO4ltupfaJySDGI3nJ0xA7xC9lN1fYZKSuCEf20kLVsu//psrIp+tdGrmazqrYa1vCtJAeDOU
eerTRNLfCBf8kJ1lfOnhKRF+XRAUPEUGKR4lO3ZC0kBO/WHxD1cVZa+iq6Ch9eJokTvV6LMRblD6
HG4wZWfqW6LW1rzBsZ3hzeADMdUYB4A191RSGNN6T89h6srSP3NZpq5ZorsqbMR0jcOBYbkW62PX
YrDvoqcLCoxuRDQOeATsUEm9FcZylEMW2wP6Kf1e1DC/+zf6JZ2ffY1adqvsLE98gEO/iCzizU1R
hJWxnUm2xryLVUNtqJvrmhZjo4jzRCLIBIH0qFrK9BP6BaH9bL3Srm58fKS+KQ6MuKwyJYlEat1N
2buo2htI6Hgv9t0W8OG8cY38jG/9aUpnFYVolf1q4YCCXh3r+ATe6INutmTrhvY7kZG2fbNL8wbP
6HyMPFx+3rWEQLOiZiSbgH8CH1fkImX4gqI/YNra0VOOXF4gIbxslcD/NYGAOTRUSepm9RdIXLC0
WkLeQebnmxORlfmz/94OJfHlylOmbN6LIsRLG9EXQwbDNbbZQA2rTJGLdGzRLiqcIXMWm2dNWtS9
oRcMR641ZECyVQS8Dq6bQJaMpFJIu0PN78rVCCV5bg52nHSIcxoh6MyThWk8eFRt3lXpCyZhp8Ls
6nMCs60fPS4y4US+nljSsd4MvbEH5EOE1Zzg9tEka1iNoTDvpuZ7xNk5e5UMvtDwZf1jY1r45nO3
eRGykvbCQ84sDLl0eqOzPL1nV6d9BXPIextCC4BFT+LALe5kkt3j6cQRVx7p1GE9IRZ0rkfEJE0e
4WUqtQuS2pU8Dz2So+z4Q9DCyDwlw6zHtX+2TqNIOwszlIrtyXDft3oPaIaoU9DUckVlmLfZCJsf
7oG5HvcLbM66AyjHt4Uu0JGR7Dnns90ZY+e3RKFUiSB49hGlqUKQYMB3wjV9AeLcwEIVsm3QBo04
fkiJMZy2qLJEsiXs1xPnPe5mUTH5IW5cPXPzC4vj4zzPNeo1N1OsxbaJMT7i67Ng3kHR0F2t5BA7
At/Y4zXBhfUNagzo+57TlTBQNpxp6/iWxXpGnOGfTKntS+oMOgnR51d1520/1P0tel1bGndK7jcJ
d3SdgbXOswDtB0LbTToKSaoNqqMZrcgnvZ1e8ihCX4f1WjKLpuEjGZh8w4h/4ryoFBb6pUnClnt8
JRBehr8lsd0gOYdZqxbmJ74/BQri4O34BaibBXBb1iYkbRQ1E5yLmAYfZOj1ugz6TOfyPTO5VTri
XfUSfcSthcQCU9QJacbbZX4STspjRMVMioLZt0WjSRce5u5of2PyIHF4BffPngb7ca/77k3/1cHB
oxVnfVkI9KnZDU93npc/8C0US8yvGo+rQmXfKMBDtCL2EAKqAvByzKYxiLulhhmQqmc5r8ulu61A
2C+To+M6WiEdlTtGfpLOE796CI4Mqf1sHYy2jIFAn2OkPKveTphwNxmKRKW7QPbfYxPVJyqB9wib
++Eac1NZC9zvkMQJVRhW+eLkG0eHY2TOK21dss1UZkm9l5HIaYfebfKPDtc1aUMa3H9MblYXDgmn
qyVwYrSdtYmg4HN2QQm9hKX1tmmLgZmLLdxQjRjdBZkFIF5BoIN+WTwAykQe7oBbkoJeZpvPJ1GN
nWePiKJMHiBCiY3zwr3S1lWLtJ4zR06CIyNBeAjKEyevD5VHeUX9I/yjDbIFv0fm7KAYc+vPSudh
qfQgt9AshhF59t1H2HJ/1jggbHkXXlVdot3URmIlFOJR1K0PmfbqRr8er5uN9D4wyDaqCh9regcE
aBSmJEFed1cjyd60EsbQ0uZa/mDyU7iE2VoxcQwPZWlWUJ6tKhwUrFPsSRUapYMvF9CPhGUJBKxO
K8j/ilu3dWC6j7cZNkEoifm4bAC1k0GH8oxCmPo6OcW4GT3idKf/c0FlVzECqDZYi6IvFx8DKUsM
BSgUNozn1O+Cv2fzpD2zpU96rfw+8kek7sNtrkE68gPTgz4jF+7FOTBYHnxA1WCJuG5YZxf06RMu
RcIRPjcpoT9LPXO7CVSS4n4ajrzbgrbH6OhzomYU4ady0Fu/dtBnMzAnBIhCWp0rFQ9gFt8hA3AD
0sm5HCt74KshbXJ1nSxzIyVL3q+UlzsP74QSH0DloD8pPX6QD5RD4gVJh0esdgrP3qhMB2hkfTgi
/cLNuSfxieEEKGwGemVWA9tM7O/iAxeI/TN20cQosUZcXx87qWHnWJwSYtLOP96IIfUNxPrHjejd
DNska8Q1AbnoIViKoeJWXoDgb1o8C5IhcaqhiCUP19wSqYsPQsmw/S9u08E/FiDNtA6fY9FGm6tb
DzsbzIqZnSbVqhLLyb0srb2wUmfQ0aOp8AwFsobIpxpCOnmE8hDrEuS9l1lskKz9K7A7UZn2YI7p
dWsqAIw4E25F1P5jq6LdYa7hyjMnyfjsnQclDkDI6/EEc+PW6y6FRL2AaXHk54gjJtvMwAWVY/Fv
VOHfMZJ11deYwllw440JlfB38jEJgejU8MKet/bKaQ8m0KsBKCrigfSDafSviG4Wa/dTLZ3cjmhB
rKEGNKtal1CJwALa2iDY+4LmeooJFbYMbVBMkOhzVs5dWBqAptCH+cdKl9TAE4oXIKIGspg7E+2/
oA9dV1+jWGFidoGyHBr/Hhqb3v6e2qPLdiVa169F+uRx1/otRORXKtBf7Lb6mbvp7Rwd/BBItdsw
VKBoe9SRMGZUUHM4ayq6usbzHVwrNAZ0hp07aGBb9ihixC3WepiofE97rBcpzSanOHCwfo4L6EBZ
eJEXbeg0oWh0bELmNTpzaSe29eEsuxf9XIi8NuyYIHDNQ72vm0kjzso10g/P1jaUP0PizmaG9O7t
9sQ3udXgxdzC3xt6MJr6sIr2zGMaL2gGFCgifnkC5RDD0gVCTSsslpj1O4n8AbHG43S8uJ68q6K+
VTzXkqmsdLYxkuOL5CBOau8IhQc3df6BX3ABcSCsQmKxoOzck+eORZFr+nXpgkaCiAyhjoEWOZhI
utv/P75CRfi3ziXuL74e3wfZ0mcoo9GOJBCgSGG1uFq+934t/nyNUty9FTrQjLydsGtfYovvlRA0
qMLJRnZvXKljMPkkCGYfjEVcbMDf10Pt82T6g+Fq+Ag16FAJszaEab+PUfmZYOYciDz1fUzEVnDF
ZcP+sXI7zf9/nSgTyAl/SmLFLYb5XH0KrYd4H6dUFU7fKkrVZkeIgXBK4IlDI5zoxKCQ3ZDnBKPj
Gb5ZA1HvEFJmvGZw8IfcLjG8ARg/nmKc46Qf5iV8ITDWpS7wQi+p1BcUrn1A8wM9r1eiC5ReRjrL
/7KopQF4lIuxzF4YYUbD/vv5Q8PRmlcRoO+j1Kkn9KJwa+s7t1Ofp76khmBbODNR0HNkkwBUtzvB
ZSW0xeM/5fFGGmsiILpF2gF0FR1PkawRsMArDO+JQrfCj8Wa0BvaWYcd8VkNCqZoiiARLZCwANAq
iYbObmte9SjTiW1Z53rx9m1pwlch+vLEZ07jGe8j/4xyPCBhQu4KtwtKPqfhyCzFv6I22a0FB3E5
f81Fr7sgBqBXLOMfmLfddGM6x4qHe6eyaH1fc6k27iQoj7qNfLu5FTi3yWSTjcdPINmLQNe6LSqj
3wg7bDCWW4SCHL9DWkngx07pysy72Llvr2yuZJlR/9XvNA16DbnN+n5tTfUE6NjG/CZFnn17AlH7
T95DXvTL0+Y/LYHsLMM01O1AqJ55sRkMotIItvbDt/iAnJy4eo+7vkqcqFMNhdA/STC370dPwH+t
abyJS8FLVnjUgrSxYQBd8Zq9ZnarjCWsVpiyFZiC9Io/SREyWCMIjSNOktp+pEZTYV/9Mf3gjFR2
6NjGoOZ55ZnEH4C+4nDT+J1yWv7Cj7CAUR4iZPzMg8VLaSZrkThtmkiBRYKDyPFZRu0z7sQVVnuu
YtK4wDPHrHclEGU+gV/9uV9hoRoPGk6WSiJRAT+yyCoYNH+9jiklCUKxxQgNbQG9zjxLtbbFy0xc
3rA88pVH/cZEOF+rQ/WqRddksZ8Yg52RrORRbNrkyLAlBBwpqExh/wznmG2Z3Q0x5P4qqAMANyI0
SNQ0PLuzGHg+Ge9lBnX5NtGNAX9GzBBPtHOXfOdSF5q8xcpejDPBnDt0e+JCFE1+/k49aQpe2SzW
5vgqeyBd4n7O0n/TGBlmqoz88MawElSLDqyvFMTBSJCHXtyD8U/88Tc3tP+fC3oSTYT9omyFNBbh
QcwueRhE/VS9rN0lwzsAaY3iQP2LCsMeddEwToSTpTFp3joUlErOVDefXgmw06ZI9YHj6VNkBeb+
p4/wi4Dy8T0tIHk8OOZWZQYrBWVCOHrZzHYkLyYK3Mn1vII0Lvvhw/B4EMyDGTmk27I5UzXS24ad
4+tL8706EDq0eqDH7yQey2+v5UbAomOBRNCsv0LXTXAwaQqEHe/RUL7qFJak8XeXl1srhh1nkF3A
nGTV+mBdNu2StpMBR1g3K1ZUNKUgWz1JhfXyJkj1awCmxsDc0uKamleqL5pRH6ikjdJnGlkmqi2p
bHCwuDf5KSG1M3N9JoscYs1cjxed8Ec3CH8WMpiJseCebHPFuKvSrRjxMVRRkuq0Sx51RSLMhwxM
gR13nTCe8H2zpBPu2SqsJenytNcfp128rkq+vvJsGR6z9U3bEhRujKacA3SE04p4LNqTbqvwbIl1
e+DnhLl6OvK1dEvt1r8Y8Gk/Qm0+hVLb0sMBDbJ9+nuil/RYnkno4Mduxwhu+3EdO76uQy+zjyyX
1+YNXun3PPTujbVZ/4NMkzizYPTlWT24XQoBi5HAqywyh+o9LWV53kmSCkTzSQptiRB+2RE4HACH
P8AJ3LUGB9dxYi4EroQp1jhVf5YCFdple5HcZgiqRWxf+mSwGEto/6ctAwIoi8D1APBSz+jLaFqy
di1o3TB67uEGEz0e16Ge032g8/8INZ+luZB2pDQhdm2nu+6mxAAUlH1g87j3u90kWN2E8OK/5rRC
enGtadavynIoJTtujMZebsmNYrUaKMO0fVu4pRrFaSh0veKCq6tRYUIfhZuIfRdr72PLeKILyBT6
HZOtaQTxIXyIHmZEnM4JwJYVZyJFpW9lYQ/zXrrAOrKixxTOU9KQHyTYzucVLSfgFmFBVtXzHI10
9TVXJ3bc2UeXFe0OQY2JxX4ymdiX7ZWRkdsJb0SJQ3s4mkeVIDhMkDWf2egWj+LyBSmcEd0HENJj
0MLV0juy9jodA0uvYbcO1sEW2wotQZlBa/MjUg5CHAG9D968P0ZwGvDmB1GxEfn+c9JomHO7nM2A
CElwkHAcRugGLhKLgK2Ets4AtiBbQ1F9aNFGGReQk5+v1sAwVa4ScaijQFTqbX1UIqiHeWSOW3Qv
kDoauxWHB32gr7MpMruj7WwpsTPpfEUa62GOoT4YqG6vxkupb/tTxjeX0WAIgwXSHf9UyXHAwDOI
UW3uDREVjirkAyYcepq5+HmLQozg8/x53tmHEi7qvzXHqm2DJqHbazIYWzVDyPx0CYGLHbAf57Dq
01Ob9gpAPwptLkj/wevaIM2Rb+682fjrZa0K2TdrXt+48qRSO4oBbBT+hbXcyZN+eGIoVh60rT5r
Vvh93NqfJoa3zva2srZP80JXSlrDSyn/VgtJHcKhJhJCGYdtt7e5rUDWGFG3UqD+2QBHDfZRzQ7V
Uual0c2D71Uyj1N+c+L4dXk5eFZ4bi7Q3gEtmyr0EkfKlAJ6ErqFOnt5G1cpAhyckoCYZpCDyYvH
g9dX3UeIHhyuHxqSk0GQkXUOVE1BKIS31blP776wXjHwYm/DghHUTeWanXhrqH+RWOXbIl1zrPaO
My0aAuWhlppoI0jfvoQtu36dq8fqwuxGTpwO+VMFQdclXky8b27Y1bjF8Ma+P2d2eGrc2hXT2/LH
qBg+CBQz/T6PZ/p0TVMKiQmpsh7j2oE4HN5Qz8uxNMrt1i/4lZCTpMBnUn/Pzj55cPVfmxW2OVqM
1MPeNFXg1h0cnnhQpawgS+efmKmyK0Fly93V9vPtFvywdWOK/f+9cjPulW+sQrvaCr5JDP/YTmjP
010jxGyE2iHAxqFfTB9dtIMQ5h6VkUxtBL5RWP+PkpJtxUoMgPz1gVrynbgblKyIl02zKEovPF9M
qPYGkg5YoRmDLxgMflsQhVHXXdO8rvusLw8U1ZviKMxF2U+pWKVs6795sK1LxqSlkxNnZXqewVTq
q7PwERtSVmirDCDfv4Pq272s79FsUXJCKm5pYu5+iCBPCgQ7JjUQXS+kvY99XAiojE5XKlWxezKA
7gVukrnCKIxKfPlKHbVoCUD0dbMl/duzh3XNLEI6YeA9Dpf5wyuWtILNHhrkfJmoOt8Z0glFlEUY
W2I168oDjeY1de0oE4uUxnZP4xPf5ShomAVzfbOY7AcWA9qcFPTAd5ZZ509767qM3CqXRdarVwZK
xSdbHZuojo6ZUWjKs21Iom0K70t451U2P9KqG1pNPhNsFwdMIUHASYcjL6xKRpx7sMlRRgADKaT8
O6qpsmVoLwl2eJ+0VzLIwZa0pvP2nFDauoVZqrZAk5Dwje0U7wstQHQzW3jDWfSn9l8jE3ZtIJbZ
ZB/LrP0HLCsUbocPb0g9scotiBcc8L2sukw46uR/0gISxEnN/m5Oxj4WaJmfUrhFQuWvnS9hPt0e
yzgSm2E39gX0IaCT+rcwjVkkHc1PjFFQ+CcNkRcDS48WfGIpp7BoHfOrTN+RikaXZEuNOfuIpPkw
o2UZrYV26u/XlziIpZfHiPlZ+syzzq9RY8WrvFa1iLA6uBCEHRYwL2F/8idg2AokAltAhYJ5qKQj
iOOvFCdlcKeslI5FrmgDTrlnQBXRuc+96m9MIbWb3N9/cLRolXhlYwVe+67ocgvffsmWnynJxuhl
FZGon2EEqpkK0FNkpCXTUhuPt1GHYQWRkWcp4j5o6Htyl43sno0SPlC91uk5T1V7vEsJweavqUiR
P3z1Khn4c8Mpxu8rldapV+z6PpSLcjlyzLntoxN/A/OL62Q6STcMYD7KVzi1UU7Pcr57twysqgwZ
2ZZSnEYmlPdi3jL2aI1Fb5E/QpkaJRe3HTFqbSPleEfHSfjbcowqhDbFPow5LNcpJMhsNu0aZnNf
+ufPmkkVVYWdxBXhOivtEsGinZ8Ru8DXu4tLu4CcnIyD6y5IVVrU/bO1XTiWxm2VYPzrK2pup0Nb
djHeYQOqjwUXXqT+8Rul4RI79HhiHpH+ChDjPyx52dzZCSCz5CDeyMFoXJb98EVBbMgPwl0KvG+z
UMTkElvMpWupTxvZi9sSWYIISxU02wLquSwPQc5WFtEaywHZWwKzmwa+iXMv9vrVLrhHD1ynWr5R
zD4HppIry4V/sJTxDK9vJcLJf7AL/C9xu29Ftu/xy6iYikl2EJ2YVtYe+BXRLfWw+8u2O0NQakRE
cOoeqAnzaji1Osg2cKYPRiCvrJl0WEIw0r1kdgcjojj5xLBH5/PnvmUFG85/kR356dEUMyevxPk+
rjpQMGMF7s4xQT8zxvmDO1fdQk2AJBrthCbWik2Sm4meZuYIffm/gyL9EqWQYcuoknn9BaJVHrsP
U/ntLVaiujTD1o3Jr15DygemM9HCQ7vUsy2lweDfL4Gm5eJPf7bGkO21GN1A47JDOotliV5aa/uU
r0NYX743iqxxl/Bj3gLY/Bq2LPCEEtrrO87vTldKXqLQdZc/kWyhllopPT/+IkvzRJyS0OKvc/y7
A45IQoHpLIv9tLqdnro7bZhgp1AfZJ8DWlhRXH6S1xRMLOU/Tb63NrvjFvfoUKhKRyNC5l4wJw4o
i2ia2XFwRIIfBt8Tc5ocIO58ftRjqFCe/U0qXkejS5PvMtCmZ6dojt5QiJvBgj1vpO+NdzLhLJK6
HCanyJjOseiXmxPC5S5K8VkxIsjZALz9TJEIdbpKEe8FI6WkgR4Dj0znt+JjgJgFy423TOfGGUyA
KZtTqPt5KqLZjtFUJjhLpP7bCABGhsfaDcFRHfplAqCxkDqG23ri0OVkZWbWQoB+Q4auaO59qyn8
BPeeGxfA4qMPX0+dNISfPIFKIAtuEV0ij36UBqa6zI/yP/AKnimeNT9EezgNEdfEcSvZl8VrC3u+
oejBsM7xm9g5jdUd44ePYDD6qo3TG+gXWOH/IWZhSbWmqJW4j6DpZUQCFII4XxqJBhKwAwoSp8Cj
iG3ieLeoPLJSeKEbnBwVYbmgBhXKsSubBlC+mhq9VvmxneoZ+jnh6ZYD0AKsVw1J2sIcVzs4qQyq
uh9qR8haBAVXxBIeUc9+QXPTYwjbhpMMeC3KkuQiY4eJ1+uL0H/DUqpotGMeCIGxzm4Ceyk7jAzE
7ajf51IX14mk0cLvYzo2ilUZRM1kz3UbqzRbqMydEk85T4+hns4bw8CDVHZwKBbVKoImYW+dV9Vh
detgwLENfUmoDTRTLPMNkME9OFPnRfth+exezAEuJldu8Vomnabo3c4gOYB0MdWJwYuBS6cJbf9K
JWm+ZM2XYXH5oXn60J0SWlAnC28IUwx6Ns2LYcw5WSEGIfD6Kl6V6yrKdmWQxkVWnBV/Q3bPinEa
YzBZuY+kQrbT26VoVEgIUzuoYB0XhlrLOJ+bSyAQ1ykJtOsqGpPyUWk9TB8Iu3zMs0VkJtPN6VK2
BIrFF0YM6gYUD8UNnleG7zAyw9o4TRl9op2YJe9635XdL0pTL5kIP3+FLKFUTwL1WV/mIp9rooSH
QUXVghtfCKXr4Wd66CbBAgRCzf28oaysnZ2p/tKN5lV88W6MRWzWo7Viegka+3JHzIB12rgWkz3O
VcHym0zhF5Eb6g5ji/mbWaMWozm6qgZjKt7hRW1f7DWu6NYK31AdGnE9Rrs5WijRd/x2j3EXvCRS
T26re4s6BeNzY/qMo41ZGY4WMMxjLT9+iVkoJD8pGp0PFiKnGOx2EJS/T81LgHucOMv51JMjcQXS
MxlsUxUZ3m7yjYgPPchDjHtmsVjAjsYsWBjVVfKNvtrQ/hwl6uQ2Zg5JdhIzjeHm8GAgb0v0mNkt
Z5UeMioCFsLuZaxpjXJaUMqxIN3ysc8hWmiBK/7/MITM/tvGlnQ3NFq7ueK20HBayHaxz1EB2MEu
mdvJobBQHqJz2BW7gX8C8v13RTz5FUakY5/ADQjHYywJbGodF7vT65IBDjHUT3ukeHaqA3m6V1wV
jhU+sRbJjQWOFxctpUjbd4a38wtOpwIoEMadY3nZGXO8wtf3XL4raer3VdebbX2v8Rt+vRmLSyaP
ucO7O6NPkaXeqd9BYpJPnlUX8NYzJYeZezlJWdNCAJSyYNXa7LacFlPfEdrEFSbcECILn8vaRXq/
ImwnI3FfUj2Xv/u4RJ6jw/b+YwWDXZNjBPq7UAoVz1zwrrw+3ljcP8MrpWwx5r1QvfMlm8SlMCV5
QcQY4jUaLVdek83nM3wkFYJR3wor4Vcev1jtFvYA7dcbL00lmSyUZ9WFxR5cSXTKUlYGS/E+Mfzj
SEgCWLEhDDd6joUSd3XQyLHDmSrspBGTi8tW9S4+qMVYEcVhWhZyzq3lq1NOmCVw7Pzj4Jv73a/I
6F9UfmWoQVXQpSxiOED2EMHB6xy0Y7l8tb85TytHsOP4FFuvrMHgu5NVguKChMxaspKQI/VM5X7F
RWIT7ZR7AI+H4BqkXyWhw+dgjO5IxZ2jWsReSTcfTHvCZHBBMHqmaCYmWQiZC0UXXToAPZEU6QHB
d1GAF3IGKpuRAJmnsOEIqIutWB7pNNPQWiTuEix/BZZM7YZvrDNDPJ8N6ZKHh7zw0H4vVDoi92ox
w/dMOZ5j88BenVIjUR140S7Xatw7Aud2lBIXt1JTR0gW3buC6AdhZGFwPNfOec9wyEPTrjWr9EO9
EKyBQDa7BdvYzbRJD5fZZEk9nSyDvWopYLdkMm3+78yBcOlpXCKqAbkha54sPh0lJcx5wHpCTdWt
snmQ6qgAUSPtYEgxXU8HDhoyAASwBoX5p2j+bwypScSwAOO5t7K/dZJiCUxp5l8wjnQWu84ZrTFP
qUrkRnAP6EsdNI0gwpP/PJgNl4o0ojOPYfZyz3mYJsmerVOmn8lppia3Al8uvEt/kiPwi4+xsED0
LWZDWPSFbYH5TLtranxx1Q1P8StziwJg8gqMGXyrKItwtpj4k15Pzsh8PgsGWlKWDPc0/kojen0r
JcSPIInmXaVVhK0TeYWUUNgHXPQJbDCGPBpxM6j4ISO7eIYWV+fuh3keIVFYoz6MPaiQsLCj8Ynn
jykW/gOigfg6AVVeMg1JJwg16E3LYwJAo000+GrpCABt9y/Ih+dHpmxN3pmNUgjr/S2gTdKgrwj+
ZCOKZFnB4R9pibFYztVCe0yp/HjhNVLCb21CgtbjMTmfEheNqy6x9Oxjn5dZ/VubAaGYi2QTJJHb
QyCer/4gbUDxztsGzD0VubYcwIXQJRqXo7TQrZrTXq5JMmFkB2tV6QTn/DLwmU6SYmZD1104A1XK
t4B3ypAqyqm3jaeCzaTibSFFveLvb0hqCbMzMyKd0KKcQw6H2/9glt0sxhLTkzOgnulZCSMtppcN
9LaWne8ih98EEKeUavffdH7zWB+H+2lTmkZmN6PiwHF4TMw52q0QHS4VCQ6iGdoABK4Bey8jBv+E
usWM0sDC7b6GeXTM//Iw4W5+cRCeeNrTd9heW6IMbMUK/RQv5D6P/QsSUYD1hZ/k4XMISwofLE6E
hgTmeKUo/9zLrxls3QsxYjFMnbzV43kjy0uca0ZpTtUYUMm6d3Blh6S/7ITjGct7EkMH7hjeHD9Q
8s5nkNNdrQBPwNKqT/aiY0/UWQ6exxzllYrzxSrmgtCD0bx9pBO+g6uk7iKURKpHF44mLAd3h4kP
HKokRPrx3jDQAaIKh33u7S4XDw6lC9uRC0j6MMXWmxPCmQgYfnKbX3OJ7UY0fF8gk2bNTp81u0G0
3kbEa5hCCFGcIiSUSlc8ssOBdVzHpHAPNn6dSWTzZfYXPl3q8ipL9Bb8i6lp4aN8lcn/TApmemJS
nymlSrhhn4YWLDxQGJl432QMX+EW/iY8PkY+hFsa/MDHkVhnqMSn1po8AwUbdM4xoMdyTNRp0D5+
7Bjt80rZYxULEBceHfWYWFsJElaAnky3H1fSaXf7Va1D+Gp2a1Z5ZKpP7FyQseTsI8nGJT/anlOr
uBO24EPZBWs0Ydvrda+fFB4ydUImVljpGvMTr1RPxKowPPCwgd8O48WeQlZy2ZdVGajzfGXecBo4
7SRoPuCD5Jl9qx7n3vx6q+wEcD40MIw5tDIBpS01F9Oqn5bN9pSvmfuf+1dv4gif5sfciJWaE2wK
i17sSkj1D/QKmec8gBasv4aL8jffxHKFBpXa1qehD81/53mDM6wGkgP6y+H7WMe9v+Dh0hDntBr5
rpMaswHTkwiFu/kUEP0cVeNVvs/Y286xiFSKdwd/Rx0l3HJyWv2oTRuCjy1mXIqiWM4pZYhA5qz9
VjmTbSA3G8kBkkuSENcoXq50rLr7R52TfyNhCIG8rVKdeXWlWVRF1tQ17Q8xQzgks1v44BMhTr7d
tyv4We77kOJWtc3IAoQu103N+kAolxhrg+ejJJVzwcNlF5IeTfVFrjWQjybmhckTDw8ryMtsqz/c
hNMX1zDC2waeLhwstnDh2oXh062lR9Z9s0hYnU5ZGS+qo0gIQVs+ANL0s4H6VwCy18FNjCGDMb01
r4DIedFutSTaz1O0V8r3OSKZ68YSyvnjAtMepIo+jLqLPAR6TMRUzBTcClT45V7O1OAWbq2CeUaq
C5nB8jOPVkxYjjLa/0j+WP1ACyyffYnM8G8wWaqJuJdv200ORau8EYOYESc9R1BXmxPfm45uiz2P
zRXKe9xLN3nRNLubbsOAs/jjIGVJeDHd25lYpM+4+Ig2dNoM9/Hp/H3PTFBWP/fWS8CsOXXiLuXZ
SX0LW/EEny6p3qZf9EXNaeuT6dRVaYbrOy0XSojnfzm8owkD15YwTDjPL0oc70fE6pHRxasS1FKP
idwvVPNOgBDcSr9EUzXDZE3IbkvZiPwrH2H4k8paxdF9GFdaAH3zRQ7VsvbIDTF0Cs/AZs0iQxUE
drqWIQFnzUycXSKAX71bgJGXBSaH460m263zhHkAcRvhw5qUQONAVoxT/4rMI6zrbAEVD/AACiHE
1qoPFVDY2KHaNF+VKhP69+owOhucT3ARGxpmtpe98IVuhxmUUHrAI6yj1CHw0HSVNPCYyz3a9wUG
5QZfDQfb42CxTK/g6PiCTjxX4/tWL5bv/4RG78Wmu+SqLQBYITPcCt5oQKSdKM9JE35sGUrUEB3/
YJjc2CkPKZXAzu9jAs+CbMZpSNpLvIfwOiIWG4MK9Spw27R+uE4J9Cke87c8M4+PwZe8XZruRJt2
6Wkqr4eUYlyk4/PFqD0d2/oFkkKSml23jQxIrxwJWlZAskc+Jz8SwixV+cKcT49TDn6lM4Frn7em
yF32oICQmIhGSKbWCTvOhDiBx97LJkdDlh7nyMkTTP/h7NAICho86apVA4Znkv9vhvhNFf3OzRI+
jijSdRDVBloHYVW+TvZRFxQsPIJwtcX5MBjd7Zt2zUpyBgn9uDVdVmNmMAidKi6/o+BX+vtE1PrR
BglvtYXRU7PsCRdM6TyfQGghEJ8A11irfbP/XpeXfP62qLeW8k1gpchefSnPXNCVhlkDjM+i3LiO
+W1Zo0bZVsM5ta0Wvfq/zA6l9lD18WSa3gcW5rzsA2Fl9k280q6DBFeFepA1gWdHQQ6fYHdnEIHR
QqLlynVKTwnLj/4wO0Bp2cVbEZHYqtbz/j2dfw1HrWEo278aBY8WDkDNcDU3pOO21yq2X6/iP6OC
BxzApK8w1cKGn/dkZSQOmxcTGGgeJxFauYbxD7HSrphTmow+qP5KKs1O6apduXHV2sAuNBtc2wAq
BqNWjoxxcC82UxDceDNHG44U6C58ydEGyYz1k632XE9YA6BFdO0oW7uKQsGDOt9gyXBWA8agpM3U
DpeqNhi7SCwkFu51BczKfB/HqhOKT2DmV4zWrxzG4IsviSs43/wEUk91yq7g8Vtsu+QFVesj52GD
L8zx80Gla+j2oai6xQ6lrsQr1AnVjImd/ey3/UAPWyxtBNL7NIVLMvHXZwRiVbKt4DXw/roBAsj/
c0RWmMWICNTznpJvsuDV0V3lfsgps6EcAiw5pN721vkjaZH7B6ws/Ghdh+ge1EeqYDGyexACHtO2
TEdXGMcI77X2V2n3u6MqrnKo0IwZKOmvatfAnGW8ifjplgY0hfM73Jcgv76IOOZyFUhS9xo7JtA8
SsnIzvMzUWetTDqS964t8TWignZByuaVPcE8/c2L+CwGalWv9lR4oDOikAwex94Nm7hmv2JKBbq5
gRf02dkRotx9FVgi/gOL50gO4by1bhuCM4q5ClnJXONdNrMYVS6v+qywCSJExlckINA0inh77Jxh
MHXQh0wKriXzQg5ZaN4xnocpWLRfc4jEH/JiMeH70+01IQWuE29TCU+H6H8B/zZd9LUfgPzeUivk
wbXnGqw+Yps9iLiHSodV1sRO54AFkRDSr1wYF3f0bXh9u400dBmwFJ2DjbK2O/72Uyyik4KCh7oy
e2ymmyygO7nEPIKx4dgICK/YtLnIetd1cM1P6+4QcfYm155Xp/nzbRjHUzX9mSzq9hYQPcfGtg+q
hOa9N2jNfKAGy6HfQjfMDIL6pF+cyjcODUf3kb32Q5aj9ZdBw2tqOWcVGtMi5zN78vajmwVXEnxG
NmE+fm60QI1Xpb9AKE5yUtAQjKMEb+hEkCYNY3mNM4VWnuzo37EoQKXMMlU5IyuP6akwPAUN4adV
EoNEaijj+OshyfCjMVB/H/7zXHz97iTVAH6FUYfiUOEMd6k9lISGfj9SP/p5XunEZ66wE3W6d3Fg
ltOyQ3qG25CdgixNrI7E45pvJBEKqoqiEG23k94zspSVi5k2Q041ui7Mvw3CkTp9YzLeq6wbQKS3
x1y1Mi8JFToLx/DufM9wu6EKiJrdjY8CSoGdzUDabiOCJQ6d8ugwM4ux2uDanT9tOa4BqI+AM55e
Nyt3DwekzXxn9mDz99++BqOI4Q/Lksx4dcZ5w2msDjEzJ6tV5dQXLjz5thX066tYmnKMtbUjG4FL
aZeBUEX11DGy767QAlPj8xX/4UjBXcZwgn2K8SPinYOo+1mgxpdBta8RcKFbvMl0lHzbTGmDjTzr
lc654jesPix5FgFjpWAkSJ5Hq2we5YA+54WYvuXCqGTfVOKy7OQKrYqNfkIkbZVhvNRdFxQsmov1
aMo4sQWhk/6VtZZ8giq4MAMmBvYSng/BviirU5tFKCZx0iOMdPIxLGdt+SRPK1nJmoc5tqfhQAeV
p/wZ8C7m1P45t6FL3AXHK9hf8Yqj7K86f2MQNZNtsKfCS9jIozJZxwDn6xF46pC8KxnP+tgU+S9M
q5y/XjHFqHBkLD9J6CHvrP7U8LEVG6mf8h1ngVNCAXkNENF8cghut+Kq3aGxSH7ZEz0O/br8V7JH
10jvDEu956zivLawuTUjnzZX6575QyZNuJv+3R+V/60Xx1qyUiXzpmULVw0YyLiG1okg8xQ9bcPw
CS2F63o2egCUbjtVO8MlYytrZVEhbFqYWIqfe0X1FO5t89TwmySmcohE/GAtA+LVPq55WDZCOOYU
4ggfuTjGRG8MvBAkm9CEFr86DlfOCIkDaGwWzSyGt1idDMNrTveRoLjXtUHcrBirfy937aRPZNQY
6gba1Y56uIjOcsQQAl4Xru2Nr2xZJvRNPoKLVqOsaj3RdHMxv8WaFNh2r7986bXzybZQRuQnxGT3
lpITD2q+N97ZGwhaxVXC4TQ+bz01dVWVqk3USzhcN+yKjW5EaAi4NT2vjJwB+TVg12I1fDguSs0K
W8dxoZAb2KHt/Dm8ffUXT6iCjopjbtW63+NPcu9QT8VwYEKUkeHqIUCcIBdOuEvVjPl6JiziVbgj
nVpwtyaGzKEQlYuW90O2a2RV+07lUKt8f+279GZP+CiX/+sfftQAukoVpqYKMgRLGeN3uYSwda2N
tX9uVTJJ4urnjO9ET2IG6Uhy3PRYF6pOS8LzrCuQQQUrkJfm00NsWTdx1torX6JEzmO9A4+0R2Ww
AC6NXY1KW/UOO45J50ZUEl3MG3f2hEy19dFOkPCD6iAX5mL55Fagkr2/wP1VQLhE+8U+j4RViBjk
7ChQLFqeCbEKBn+STE3N4rCLhuzL7OrAlYb7z28L7Bi0/IKbPg3YwGkU6RuV0TmlEfPURpwmbAia
8SkdYTB8TB+fiHjufqOYPUU9uYuxJ35y58KP6xey7eS5xoLMAdxCoUaTUajKP7Meb0Ih20YLlL+2
mRpNK2MrB2syO/GDAahDHmlzMTzspASCTrhrXTo2DlG959+kJoxi9J1coYtbrpnvyCItbLVFbTnf
9B8cF0COF+yJ5i3WxZZo54ivS5W4j9kO2JkJoGXld9nHZoSKCz5DY3oQ0WFlU2UZ9xwT2qKOaa6E
91x1GPlXHQCryNST0grjXipquPaNiSrQQSgz8dw0d3+Q7DF0Hg4rvfry4ouvl8aG06AgcctrAbeZ
9v9K0gFutvrTrJCszXOxexLQ3m3YzPUFUEhl1RMLk8hZZi+Um2Hnty+TFEJXIAr6ouvBliDPoOWS
VCNA7B3NfbL0K0nXhuWqO+3KVePOWHUhm1WouD8D00q/3aQLWa27oEvw49VehKwoM13CVX/KGVmM
qUqUFZmk3FN9KguXJ+VrRThcuV9pAor/WA8+yQRhHKMbuZNWoeFQDn0x8PhiHsCcNJZkPOpe36Xr
EJQj7/8IujzScM96OLOW3FaN9HbXXiRJfhrsLbah7uzgFILxkUW/oKjyECvh2WlQSWcY/E2iAPdA
c7sQCRUsuO1e0k1XtlDA1WmxT4vmqbj4DDw+00pEhE/STgNfdozayawGqpTJ5XjeRiCXVihhw1y1
zSidbhpN02NeRl2dXiwDOngrmrNgGKx+Q6/KoBmVRW9+YQT4ac2cf/1LVcBaryNPd0Im9htjEsZG
0CJqHl6WSuZyNRZnKEqSEnEKUioKCBIFzKmoM10wd/dl0NgepaYnYbkNbcc5A45H3zpODdePdEVh
h6w27YPNh6tFav9FWVGFPQ6N/rfFmUpjljZXNg2mxgzNXXZa0ncusbSwvl4M4G1CgxkogwCINVx2
wF3CA0i4U+2cjoaJqZX1Ju5xCIwPqgupKJD00nUW6zJCpoJEqONRVTmM+E3MHnqU7rsU7/LUqj4U
XQ8+WtoNScVtw+xoNiiH2YCIuvpHwsLg4ij2Veav4OttENBvZzXATJpfbMuDJxhhko+7BjFWBWyI
liHiBzfHi7OOmxQPDgQWoXlW/PMibv88U+IjCirfsX25ZfW7gd4bP3VIk0axKZa22L8lIUZZeCp9
r1nVIq1vAUkWpmenH0FQrAxjTjxz4Ucwmvt6uKrllXr+U4DIkMGvqnRA8kNhH7d21xvmnAoLcK/T
xAfptZHSSKWx9KJm3vlKQwo4fvk2hZfTNgs2xDtWS3pB9a51tulA6n3jQDaucqGfLG9+2yxRWNZ5
Wx5EhqLuryo3RsANTzv5whtIXmUsLTIkgzt+k7Y0pkkhbN7dpBmjayXERWsLOCxta3j8NlEr4lGR
9V66uh8B/BIu8JVMcCzaXLLNAYUMsom/BFJBU0gM6RS+/1J1YWhGLgHrhS8vj0L7s+CJ/YULheoC
V3xY86zfQxo2hCQeLxDV4RxW41+i4kPIb4t8UQPQM1znCjrDxQO+PosWEYywyK4dmMHdWNnHYhpp
3o3E4FgS6THVHtVV96kmV1iHWTaB+N1PbmmD5vpjHxNhFN8O97/Bq1u5vjRJle25xyEs1Ihwh3VK
Wb8Q+hV0r28TYgTmrfvTg5ktCI2hv0EToOyPVc/wFdkPQgzZS+zyDopBeSaZb9ICM6s3sNirkncF
wtNaGOWFcdpg9IHHnHyF+0Hj6AF0Q1xwucb3J33zh/8S8kEL7piCgx0ka2XkJO0hh3AN+oi1XT/F
MzIiUFnQdJQH9KGm6KW01Vg01Y+6TBI81p9KEGDEEFziH5p68w4XiZP66Ziw+fd5UwXJ4Tg7BVFI
XE81fqYtPal3q55LEICj6OZmTRrhbYecvaDxjUw6iVONdR6z3FYFWz2mANGXn4umKX9tdK/I7qhN
tTFs5aRTXaRikJznU76y4+gZtycsiafQvUT7wj3WKNODcziG4gE64h5okoit6Jm/XF1sUsI1VRkW
OLlBDlA7+Xo9yiZD2rjJ6hDFmfOuWDMSo/E81z4e1QzdrRJSt78sOVJ8kOFI27kREYdSdFNSr16Q
Ovqmi9VCs6Mfj7xfNvs+v5PNbU7id5sXna1gY0/q85hSeRKjcsVdWKZjNA8GZxM0jOsAPzt1Mn9M
hadXrpwKmNR4edDyie70Ku8Bt7ChhHyD84XI9h2Sh07eegneBIleBqL6zvmDq5V9OHGpq169eV7N
BWcKQkeigWj/DsZ87KEKtmgfcli8+gqCSoU1eHUEC8k4UMIBqCpTkx45iwqujWNClmrJXpso7If6
JvKePTmo57RBzekoh9bZnGizEHsWoUZftegbmK6Z6OqIvKMzQY099m497tvkdBDqA/PsR52Lxc+X
2dc0Hk0YDi/M/cR1cbIz0ZG72/BSAYRSSpl8Z/kuEPuzGDBEMvEWcOORk4w4mpYgdGIdKFmF6/1M
KXfWa50qWsjbNyTr8EcRvhSqw4/qd10auhGbUsy5mLFDw+P3edDPAPaNfsSowaFGGg/lU2TzM8PG
5COyuaYLpzuRcPzw3y5y294F8qgIi4At7Jz7Tl51vvIEgjRJTdH6PZtFb1nc9hQmsDMcbpmR2kVj
1NqYpY8PyOJgu0o3pW0vomLXoRXBJ33kdSn+zXKaW1i6agmQ58M7LAjHPOX5IObej3tJwbSRldhR
7/yWUBE1nurr+BeEno1i9V6wdef8qG7yOKdzZc3lfsZnQraz2HtNluRhORE8QkSQ99meBvWCEGMm
ogCmulNhTVDY9mMSnUWgTMKIRv4FxGVNaPbOg9gKI6HYYt94+8p89eMoyAnq2OERDCJCB2I8vN2T
7tz3Lq9iQeLAuNRohw+FjhVwISoaWeyRNf7Pl7H9r/xGmLOowWIjteGNIt0prybok3HPPa/dfQQV
7FpnBFNNlz+M/KLNXL+fXOO2DcqazJycKS1Af1y/ttLor1+mKpxyITxHUwm7EVsNO1bnJx0vQsLt
84wHZH/ugGXhTN/32tqR58OwoLnjxSReXsKyHyjm1xEyJEkB4i9tmylZEc+HRygzz4kVrlaEoAN8
9DTdWdZQYz6AzXkrhjYzBm0H5ovY82EToskkZuOfgcD2IiJU3O8HBEBROWT/Qlq1K3nE8Vctr20e
ePR03MXGz2/Ko1HKwE4cFyryVM81D39yvV5aVfY8wuKmNrGICRZ1SvRhw2AP7nGJ2xpDWwviTynB
d9l5b2aVEQmPVqDjS1eV2PvjPWvqJ2WlMoLjAus2eoMyHA7LyFNnu7/iy/a/S6CH4Tp6s4YbxjUg
YJQtwZQd9lxFnBMoOPn3VQ9bcPPjF0lmmTzye5EvXjj2ZURukEsydhM1BpNg0YVbfuqiSjK9Rrfd
RSPhIvB0eK/mwOS28HQkeLxeiUxoeVZAU9Iz4IqJ/2gfDJKks8t/LBhcmrSn9U0xrthBhimDIUlX
oCxxBXKOo3Rmwq5IleyAruA6LZbsJlCUPl9qtlcyig3XBnjdb4fzafcqaDYa7MIJeIJf2qDgEOoB
AgYCXIszLa88NKtiz6Av3uNoy1jZSRe0q59uAHrImFb+/MyEH/5G09JUw9WGLEU7tpTH5EAgNU5v
4FurS4nPmnf8m2GtThtZIsHji64Go+kItmkYfy7sm6SNEE9U9J5X+Bfmdl7qYNwMPJiNibF7ookQ
2FK2h0yceAj7ST+abqefpWoe4Dd+YYc7Kaj0dAATyiTOyqK4k/MONg4/qaetgpxfV85pqx1xgtSm
AHHVok3Z7m5cdPEUgrTFioiRk9NW9OArmiFlZ8MXT1ZAy9ChibChtDd1SVkwp/l4WxuGvI+tfIvA
MHKeFmxbBYHu0RnJESTbTKgWTxg68s7zgwjMMhAutL6MoY2nRYx5TJNspRJrugzQ3GtDwyELFYPo
yer1GKUDzEhScgk/8HkXjqyG7HaRwH5FnnOM5wCBk3Bb3c+XDXM5y1zY04MDYyO/ZdPMu66CWZv5
2ndJli+RKx+Su4c8J5LuxMH62U+G2lqqiGGxBGCa/QTWEsY3X4aikST51PKBBF3YFuerPkch5N+6
nyX33qLLjyLgyEDkOimrLwO47V+Lwta1TXupDeO7Fz0+XsucSNAMz+HW/JXLjeMYu0mL4K0Af8xa
ix3v4ARiyqitl+JD6JSzdy4yeTfXgb+NZpSYJrVsPAGaT9B0svfbWdkK2ZstrkqrFeMZQvbLj54o
OjmBK50nedVid+CShvEuqeCZ5oaRty6Su6ZTN7ykvwRN2QOSoY1Pqfx8s1g71ci2RvF2zkB89DgX
VkFA831CjL1EnwsyP5LEvHAYIDXb8Gi0RAyOu/9wWl0lr2RxyWblL+QT3fQSuQpj1WmhK8QNBUut
/Pe1ebOmq0yA5LHpjeYOdW0r3LO5kTFLMbJmqnLAS6Oth5+VJRrVJzydD9ZbE0+HldSI9mJZfvA8
vYcOuqr4CCDrjNaJ3YrZLcC/fCyKnVkunjJJocw2jjqOY9F2WNgLDOfs5eljT8fKmiIey22/45+I
KLeYPGjHZbYw6/FTt8ntIHEXJudw6whXGQfBj29O0Wib1fcom+Rv8AVjbKEdQSedwPnMoc6gBDVH
zemxfDS3foNxnOqx6zyG3KGxIaFYGO2VIGdyTSWYSwf4VB9JQMJAwQrIO3n1xAwwfNqngUPZKrem
MVlOzFw5PjWAaggVPKd4LV0OHFTRaTPpIgLvE8cmVFnQxNtTOh5nbqSVRvQdkw6Hnf0z6uZyhl6J
Qaz73di8LGOM5ZfUvqeChJkk9QNsyfXMl56Bd/Do3FAka11sM335+CLxjjcwFufqoglXw+UA+5lL
yr++idT/XKJY0dNkLgVGtk8dN7IddqnW7nm710UvGxRyb9MR9ubhOelXljpcvY5+z3Jjahy6OrIj
BdUM+rPlJkA5LGtNmTH11woMEP8SnWBGYvkxT9wlHry4JmbhnGbY6iUB8O3ZNBGB8vqfZZjygDbU
MgrTQD29vkdAFUhyJkM16U9AUDa9Bedy+Qfb8XRFYXvXsq6eCZnNXBw5wDClK5e0gP82gW+PJXEa
Alu0VcIDm0RAG1YP/Q5GTwmcGPAH8MKnBUn4mj98vDmaKNR+jZ2NgIqsGkIpbSUQbBIvTkRg9bys
fvDGdpE9pWuh7mMP99TPmKA+c/WeULTGQjvJGH0d9OAz258vswUQ7NDXEnNTRbfdtuzf/w3HXp6Z
TvgQaxoaLoA2xJtj55+fsiiw0O5vE8sg3Qkk3ZxUZDcHf3X6Tzyuu3S33oIfdyZpknIUcuDzmZEi
tDYTDNDmOGXeHrFJNtyAHU2uyifXJopjlm5u6BZSLFUpAK44goTRYqpc6SNnfzSKdKLEfwENa8Qq
CE4Mj9CGyj7iI4c0wu9CvDqQ/uPkwJPSaiAYNMLUXWkwEPHdGr4PDjPMHWkRNuvLX42JiKgYQMED
zKYtavfdndaNYaOA0K4YCnhUDaDgJcdeV/nvmoNl8diyRSx/1Iqnfyy8dnqK/6LE148oJYFNlaOC
3yPihhN2rI9K9EypITn/QT4MOiYOc9tQF64youINZan50rYaIpgrhMi0bp/PFWrD//w387By2uWS
kQTiJf8IQ5DOBU1CmLZqUgPLrHXNXZevwa5EWmflfv426OxASipOJQa/eqiwqoZf1KUdwGqTeeSY
p+DINRWqMSqfxMSqHOy9F/nIvlMKbHH+ucpDISf1QsmU8AlIjSypiv6bwWt5n39O05qNqWfin4iw
HY9D6sE77MyEhV3o6d+B/4cI+0V/ShexkyO9okeGf7ujTTeunCM4yuzTknrDVcSdw7/gEcENCUfd
UrELFlcNOhSQ4gu2Inteo1e8aMwgZSOtl9wK2pAiujcGwuQ2jI5R0gfpHKjoBK5+EavJpIUJrHLB
tsTvhpKgP55bxT3BfAQcwkRGPQ3443qbmloBnc/0ZLDsCoMzPeywdpqVJPPPnONNFv7/m0pgfHbT
Zu/eFAg55Y9v9A63HEL4kXz+NnreAi4NbrcmJ1UaS3Ic5Es6klUb/ZpM/dgWsChRPZTkZe3QQFGM
zOta/9aSmScD1UJ/p+pm/X7efVjPAZWQJqubVWyngYjDovXihK2NI2u3mL3UXR/0kirhuzq+6n9G
UGJ3ox7zbdt9n65Wi4TymWkHkts8jUWLzq6LKatA1vRSAlPTmHNnuYrqVveO0uJ5pda9JMCIOKdX
hYgQd5pqkdKeIraoDuuNUNRQdY7W4ZQwVRs9ijvLBQgPPouc42LGy9yHKffyZN7EiWMKuh+gKpCX
bJuHpNGwZul9AJgSeOVM3xX7xo5JzY8IKAhkGkptd5vp4tp56CFRkwlU0ocr+mbign9gFymdHI9Q
cG60lwnOG4HTxok9B+KO8B5EMcL2Ai/rJ31R7uxAXjJ7uiW4lwOreHnwW0MiR7E3IAsMIbpvYWiN
NPYwS00kv6rT10jPEIDTDrCvBud0NvCvvMJJkke/j8yZBqzU24mECrxENwqMDVT/aVVJ8+eryJv7
shWOzSP3g4EbnI9PWtmDBkOgyqlBkvMB2jyTJI7GROLLT1JSjuZwKFn+cQQ8Hb313baX9cOeQIRd
8P2IanwViXPJSbveI2OJXA3i6DW31W40XOPHpevKfy+8XwbY5esJtv9vP/XS1efH/xSDYV1bAVia
RCU0VF9OdPaucmkN8fzR/iWTRPRz1xsZkz2YVIbm1pDXV1DviGH5hpRov/ZongAEqolzXApzK4a1
ZcAUJAVFLFVoii7x4DgC6iI2i3KVwJV0Sm5izpnCv21Sjkv/RX1BVGaY4+ygZlORpGpmZCarpCnF
gExaWwkknUFgASK8DLWm6jZeexZ4ZIm8k0P03il3n/int3GP10uOYb9HlggxK5sgb7CyQ+8KQTeF
fKXRssmDtk0FACQO6RwUs/PYtqs4d7kdJKrNwEzGBVjtI0I0/huuu82pYKE32lHG3CWrC/R3FWPS
Dd8bmiibQheyEzhcEb7F/XZmIXB4mHBFRkNDvVm6jB6TajS2tisAhDe/8uh4JHdWmowpjxNQ3Nq7
e9Ow++rIzWhDnUMsBZEBkHzf9LQFEhUSumL13ClrjqF7b+FiKYaC/fpC5cQBDnts52lM1T8GfdV0
AZfU1TpndFhAhs663uTdHBkBStGz6Uh4fC8UTQ27XRX2/GeTAQhvUGFPeNkmvCeYAgtYgDisuClX
wzzD1NszXOXK8ODNknjaQITWVbwQozvfSrjTpCjizT7AXXSFUL4ok0URPBIYCZsbN5mOM/cWSiM5
cm5iLl3s1NAXv1mVWfBLl3DfcceNBRUcc1N334gfD2aOjbxZ+KwJi+tLC8H3V07cwxntVSpI/383
KDLDj/uJmfprxyqCa++luKGAaH/UumP0Uno/El8Y1m8pWHmorUkdsmApxYviF2VvkOdvcNls4myR
2jCcWMfqxq/LFDxSkxppef0bqh39JH9wjobey1IqRLoUcGc2K2yvGYDDQQLz5Foj9KgoCIKBuaq7
O9Rq/PBgNKcYCgeg1O20ugcCVFSyhZBDBUkbEtz8YTgnhkbpgEScbl0TOOtRptGhBC39IRDwc/im
vZp9+5Tu8T7Kmry2BsYkbouAvz/KOF17O+hypmQv+rsmo9LYnH/LgQogTNhd+R734TJz30Brabc7
HvHXezpGCDp3S6akGXVNFvZfhmVJQRgLT+radjCUxDnx+G2scoAsUllW9UzLp1QsWgIyllJe+aaP
G1xRWsms9VpDsI+eqwznIdnQz9P2BRO32jxuXVswz7CaG6EQpS/NBbhRtvP2BdZKm97QpUZTIOhZ
GFiTE4omqhMb9mPluMSPjzjJD8Fq0eQYpQS+F3hBOruOVOx+SPXv6IzrHiKM3pjVOfo7fS/PRCB2
RH/J41tzOcIfW41qfkCrkLagCGGWuazz63rk9K/humRQ11/5tYxu819+QTaf4li5jRqJzzde3K0p
Ax339LoW+eJT03j4sWTVsu+Aq4FEnM1HqoK6wEuVJui1OzEpSGtwrXB9i/63yYoJceGFyJ6AXMRG
PQRm+RE7NS6U6MBnH/7PZsU2g0FIGtkVcfElnQJatvKNQc5lUq5lQtPjZ322SkDQ5x5sR0V1OwFL
rYnLwTsWCGzF3XN0twgggXFaBvflcEVVeHtea6z2zjElh34frEfHdC4frxw7Yce7gFTtMxHh3RIk
RY1tc8ueExA+fTCh3hC7SjD+Z+1JiwK9JEjhtkCycVc8/tszpWX94fTwPzmDriFB7Nsq9hBcyRB1
p0XyJPH8fS5cvwbTGRj7S6UNeruoADdaIVzZSlbqPRw29B2P7+H9mVKascWVzwukaI5CNUfTOPxq
Egn7Ktm0fbenLStr06RyXjEXe8XorGBoJjCW1IGTj+Yzc5HhK60tXn33XY2hSDeXIB3aqVxg2KAm
ghtML8q/LETSnUVNhKEswNMaWFasSLEnpKeWBzSliMZNi+WNfQpJHaK8MjITXKbc7lLYM3pxDykl
3DeO0SAY82qQQDRN9rL5+3Kkchbnm9od2Q+64dUuftZsGH+m42Ck75GhlpChSRpTZBAT/DKZSGrk
baanJveqVq+sct+XDkQIoS1mWE1z2XFQShXOlDYiYEjTzpEcqZEEi0Yn6kE5IXvzSZD8O27amOo+
sTB+GzGtD82JynKXQnGButdfZbOnhY2O2O8MzELbXd4nV9KCUdBJWFxfACt+/IqRqT3HcrBAKPBw
FT/8/iJGlJ36hPIxx2AwRKMhWYT7E7ZMrXFzUH3GfqyTGC0aOZ+Wfv1LTrOW0f2hE+plyUFPWYvi
pDOuEvYf53W0k1R9l8e50pB/RzwZmEKviKAJO1UnJz40XiuwGzTTW8Gk3CpiJMtbzR2eHKqnZ3D9
qf13P/FvV56kd8KfsvhRqDNaV845+kw06xJK/D9wgmq6F0/EQ0R/Bl88G8Ptc4wozaIX9EBYUnyE
PHRICU5WawCoKp7IYGE8PM5kUbLHLKiYEqx5wnKCi02ZQnODqZwnU4ZlSC0oUFTNZDYtzm0laRm2
CmcqWbVFy9mp8/ByKKGLxiOJPa2I2eyn3e09Ac73+e4nP+YcMbjgVctfgc6v1zpu597jMot9Vdio
JXj+Sq72Ai46kxHYgGNkvVok+2pkZREqeDebGQrPb3LRt7KG+tGwq/NGsAic5bk1HUfKhW/8/70S
Kvio52yWAIZe6NtIi/xZrwfQPEvWmtfg8vtvwjopW4PjEvYqyUgOrbIhSCZmhsIipNvEHi6D1Wh3
lbttR4F58d8MGnO5jvEHFcopmu3KS0rrcBpyU3tddYeKZbWgrGAVQQwNkUzLZrjq2Lir9D11JFPO
r7Y8LuqsVi2K1gVYfI052AuD9A2u9vwCvHZDW3GKiqcJ0Xa+j5UzK1RJwRI2a7OHFF9Bq5a+33ve
21vERHSiP1HmlUBNB963TbWzyrY+scj6+jz96+4MVXgu6EyXDFhhQv9MaUoMDoQCAzARCQ9T/1GH
yIXemoUZvLjwtpbXg70aHglKVtuM8PKyEqQWi6XMl71DCHpDMGLl8KOTOOkFJentOtTx+vikrUd/
D/XUiiUkApFrjikDBLrith/vZkxkd15/2/UMUsVGrxMOr5GgLerRW52jxrqcl0u4QJXjC1c3wN2n
uhDeUXdV41geja35PcfrVJV3m4qyfFCmDv1YCBkcPqPPhrXCJ+RKRB0PR1AMlJmV9xo4766sAqj8
wrKiyMs/v5vnY2AEa1gzeMF8tVReU8ZaFBpYQwpLQfRooiJsRnskyT6Tlg9lkDMn3Gix8yLhXTqo
k4ing5ONVW5B78VEEVJ/4QB5RwskUOpj1aV5ZUc6ifzuNnhgepT69PRcFiOEYikYeDiUj9mCaK1E
LGqZRZaH78xh3TmlfNvXNKITXcoRLIgJerf09qwm0EL9kbVRYV+2fxn/wJWBRajN2yptWSObevzX
WP40BA8jQ6fS+Vy1P41ER364IwuBCwzfRaj04cQ4joek2R994rfLyPBQnLVIMqQ9Ke1O44KSpaRD
TlU99Nz0FU/uQDnl5ycdmaLd1q+rUK3jD6CXZQhJdYF4YYran4pYxx0B6RHhbbk6xi/CXP+irtp5
rrSMfh33wHmMlF28MQYfzqRRlWsdUO5tizEjQiz31FUQsSN6t0labxLNus5t8dm71G5HxQd4QHHH
traayq/+nzGxACWoEE2qcI7nPFJaAhdcg8KH3pmm1ixPGiuD4Q0DKoxPxc38wxEg9F8Nfi4cD1lG
gF27OGrcUXf6RvyLGD/sEljWtFrHnsx/HO8Oc+IktsG+KHH+CqJ1vLHj6BE0en2399cuh8nN6r2f
7GRvR7YcXGNHCiyul21RCUqny3MfPnJ1J+iPYZqHThj9tjI5WZ5gKPaghuxWyoiTYrsP5XGe3qMN
1jWbdwdMFn1TvKHIZqmdGt3yo8BAEJvYAvxN7ALPeVYpkUAMCGNTJCyFuJUgv8oB9+3i3ZA+znu2
GzN6+7frvSQAxHQEPw4SREAkX/+1DacO9Y/cJTRLl5Vath93hOXPTiWtT/DrrH3Y/JGSRysmJXDM
qd2QkIB3ca7bo9mxZu9xm63tMYft0pw60NdahVDuvtSk+0HnyYbow8ZfFA6WqYG7obz+hgYw+u+x
gr4R0v2tedfEWKFl2InLmfRuL+BROiJPAN/+phWmrIDKyV1BVBYJBBbmlnLPgDAWb/W3PDLZxheI
TYr8Nu0mwbI/HUD0g9RPE+xXV/MGKWzNjaQgD+I8o0ZZ246+4/0DpnFqBPtyZ0yKEnxtagSpKBmT
2eEqYSz7EXGxn0bnkkKjDsOAIC+r+yAkQ26qbwwUYuoSrahlcNg/jK65TR0CmsEPUC9CmnO8nkbC
8Oq4AQVngkg9SA8zjkr0jvE5tlhUMaZDT67ocdW93hIkhFr2Oldb9apPdnreGG7JqAOrxqTAwk89
LdH5ocGhhOGqVEPH1wyyd/BuCj/EeNHBuDNDeQ8hcKy1pbWxokhz2+IttZMb4Wv1enSpQyzKzdvw
LXhbYFitIspxewwRb9FouNDDcunXiyXjIschnydMQoqhb11IK3VbqfJV2OYl65BC7YylGrEVePkw
57Xc5OLw7hj/JSFrcXvvsmpyZMiQWY28LS+YnNBBn0BoYqwS0w+Ibf6hUonJCxcmuQDMSYcFhDjA
xzN1STJv4J8gW/O8rN1mULp1co/M8UmQWy1ZxXp+aTFNMtdgRTiRpmFE59qVIV8mKuOmDjqM9BDE
T2EOodLiX5ry4/N8JhgTH7Yz5ltcRdiV67O+Y78ge4h1Z7oVfldqKYeNtr9SdVQgpI3wcAQafYcw
DbXE1BUvrWXhTvaaeugcx43mqCVCGDX1ZPHrn/9fcYDPZF6SKs6urchgeHuXfy3BvMNY/rZ9QX0t
JfmU0Zpo3xWuk8gr56mJ2jjaz2cp6PwPTFG+Z7OZxMwbnKwFt5GyG1tik3QP8/OPa6uCMKGT1AJ5
TCPyFGjf87JzxyfE6adS9FDoE7aHVcv4VBZRAF1yqJCwz7F71nIP/M9fexOVY2d7upokuWkFDpBD
pBbEGZLN8GdLCJh9mksNPvEDp3+D9ysQP5zAlorV3MraBgqmkQLr5DZzJqSHSS12akVGu18DgNin
rItAzqFSzorZqLkEt2Z3Bz0M1m8PYNjlgG6+4EhIKoI10UCp1fhO7hIU1dzPjvlpSD0JDUtRleAy
Soi+fOvFp1F5n/KcAA8amdlgrMibfsEUmdjvVxmPKnk/gxsEekeU0BVg1t/aVHjRK0jPp5Vr12Qh
e03X4+3Hw2vXl1IvRQzszBkPLcTE8esPhGJhfwu2rQ7KzcmHyLC/GIonv/aYsLu9WX34GgMtfDEh
7wzD4HDip/PIeXTbSxCT1B6Y90f08+6L0Y5SuVOXzSFqtynqJpVWLcKmzf09i5WVhIUs7jauW5qE
0+c7O0ikM3TJywA3Ame1yHL13LS12kWJ53pAMf3MiWXxuCGJ1RdNX5gmvXQGaviIajWdQmZKIRzj
YUfBxOtE99D3dsgA2ncUw7kUkVoX2E//hhqxa0jfsKn8kgC4PXVw9203KzzRfypAByEblYxB7Lvx
xb885FmOK5J2cSe/QaI0yna1KWiC+ouZyPCnae+q6b9W3D7/5iIcSXAVztML0pAyYIK2XuDfGhGC
QdBI2n11FkJhsyqWJP+vOnVzvrYI2W6nB1fJ5ms1QtOYV5ViTMy7iaTyCGoIlxFa7cu4EeBkDJZQ
DS205s4skQoi41pM//jn/TiZpid7hjhiIlhE8EIs/jdONTLaRZqvwCEMUZtPi59Ag2YXiWaPEwkX
Snd+/zwhv8mvPUKdx8gVow4nLKOza0pZuP6YbydYJvrtI6HT9x7hXmV7VDsWEqHzaQvxaGKXLwI/
8AJUHf7qH5nwXcPTzf8omqsLUpIAA7ZopsPhWoo5pcS1KvlYI4BkbMz87coe42iRFX+L83/GHQ6/
hrOVdp7pkcHnlVPt8C3b0iiLSzj8e6NIPf2AM5StStX19jyRaqfhnNisODNeUtGp//icJUuokNAl
s3LqX9j00QPrfMRg3qRcjtjyCwRRJoNeU0mbZysrCk0ZDegJXaDo54V88VfN/6Ogf58O4cXLrAUm
HpZbvTrqT3v/KMXm0mneqJRSHIte1MxvCyMNX4/vEGTU7C+id4LarMEq05zMknQ23zMBqzHhYFhw
u9WVg66a+z+KdDPYtvipNDR+l8N4lbQzcTw4vD56gZsTb3tiof+8osnPTOEuPX8Sm72sjBw0Pzd+
sPex86Oe22AaC59jM+2tGzM7lFFfDr58zrNwqA4mnnv8e8fYKTjrj9E4ivIm2hTBKCSwNAdDykig
CykCQMBgAJwmiBI5jsOPKTFBF0z/xqyIgG0bTHyNsWnVyOO8EUKIDsNmGkCpFjjRHKHVHh4bd8UQ
p7IvL8kdDXdhe54dggSTHK5lIJdCdswOeKFzVJ9fUC+bogEhiLtVOb6SpEij2i/EP4rStNVvsv9s
cVq6TaOJIDfLTxYRHemJo6pEIrTFEPH8QSeaoa1RJYcvcF6P1NJRbONANhUPKwI2ARdDnruqVOXf
c6fVXRaBY7/jRG4Shjp/IIO6YZUnCSUWe4R7OxcyOUG36Qlgn3rzjqmDL6LFnJAe19rTATrhllmV
PnQs66PE54353ODy2dGagZGMTULpqKxoIwTrX6Ax7Ma6eU8I37jMCoavAof6jIU2Y2grDBb+GNr9
QB4nD5MqpbIx2kf32I2kdkOosG6LfGoUvbQOtijwhLlXh3hRTHjFNMw3UBt+pqrd7RSYIOqy36f9
ZGThMBEJNLIu4tzBFr9n9iyg7lgs5KVzcQk8MVtoKXI7LH77V9eSitmnjx+EojjpP780qu/Noo7T
s3iKVh73nGOlpk8mKoYECcQBVvZe62pZ5Tg0QAxIVhpR8J4Lwb1j1jIzLBIzJ+aN0ZqTm2fvToIb
QBzJaFT9nivWXUq4PHHvx1kI8EmlCZwhnhghN193Zwh6xjCklzoP8D7WacsKKIOSaZG3+Vzowxe6
xQS8w/6qzpLjhcZAWfQDx913Z+Y82A5+M5crWmMHxQ1zxE6Gao5NMtn+wcs3diF/eBee5gfDMGoC
+4QPDt9+Na2MUA0dyINrJ15dkrATtp7279Phkj0T/6y1pNB4Z4ud8XLGRPnkXe1mMfmH8N4Mivhz
yBF19mrW14gkNvxQRqXEKZLnGEKL1MGb7V5eowtulb2RZ/icK9fvpcvp0qIZlZ10+pv2l+zSgrJQ
wembXFB8d30An0I0WlZveuahLV7i1KZY/LkVv7FH84Jq+DUMPp1NykDZoX7yVEMDCra3EBE1FF/A
UAD4JmoQdpbJttwjhG+Dbegp52OJ7RWNunSOr4X59S+L7goXrZ7+pboIIimEtHp2Ufcl5srICNBp
LaczYU9YTJOU5oSvA7phuaeBO0HA/kmCJe6jj+srn1W/R1bwV9boSxeunqlsE28nun7/IFWzKnlh
Dxfv1VqP/3l1VOzdU5Q0qcN2YZPYbuZ5tMKx/CoBDltNDkOf/i8ZfXg8nmdeZAscdTmQVg0RSjqS
H5P8AhukL+lJRFWzS3r/bDJ5JyBTrVuca5/gFUM7vQXVUcBaqgPD/otXZ+2P8pSXfGa9PL9i8Dp6
fz9j6v4xpA9C6wfvWdJAG82klMsor01hMsn8tr3xZodygjx6J6MnNeD7IBgcYuFpUo1SStpmY9Lz
SVeHil/bVR/9Ziwhp5TdMjTVGDtIzVqYoORYXWCu1C8aVpWAUIOuLl3m5SIm+NccgO/mfoDijq+x
RLSKoTgJJkvkLmGb61uevf9OU7MgMXIAe9ExxXm2aiXbFLxDtJn689cWGiILhf5M0ZvcvbG/d4yM
kpSL1iCweSr9kb4ApMleYY4Rckzdmnye+L5L8B+IDq3zJGAyFADIdq/vJtqSUuNUzV29xoIbGPH+
IxwGFjHgf1bXVRZpPUpW9VyWvJ/u9/WGPCGhx99neWWtQkusbgnJ6S9lCDhvmfOWUfSIdxLB3xic
V0ntQgpN+RqThADELoRhQhsBNB2cXnW783KfDexCxo1v7zw538OBMbuKpxc0yMb8Wr9iXn8b4XLP
7prgzakMwkUJjSQLoUv1+CrbU69HWgqLVrItMck7nblGF8AtimRU/WQSqdPqFxBdLamvjUL79MvT
wFF7bNwrVfTOZtKpcx1xUa5Dl5aTNOqL4i9xzw/YBsJETs7sxzjZ7og3WDo+CSdEdM9ptw6UX0qg
7E20kDHLZ7ue1DTVWmTa1p+50k7HwOLWG4k916r8GPFQH5Sm5l7ExpGi98fEXJkoJHAbmqxiIvHm
bir/cavmiSrSK+qIXRT+PQ+/QJ/N193kI6shMqJfQ458EIROsg4pCg6CJjE54auotm7avZ4CHpvN
ohMNA/xJajV9KyfVjeQmyb8DhBu3zwMvmgyhTQ/tjKoawjQ/j+PCRYk48h8V/+INDcX/7wAojO4A
82VhgwawlvVuHIxIZayP/tO1wkfG7ycFeZYXhwJMBCY1VXNrmnx3T4+iIYpMlHOHTAavZVGXZJBI
+BwHy+MSI8gdumM/Q+PFNhJ4fN8lAQwOdNjPwLn4DuuPsPfJEFhzvXVyQ58npEq57rX9N4d29Op7
r67qrclSFCJjBttoOW8HaCQrcvEhfw6bEQhexGJu8SqYJjRrPGAJSd/eI/NRfhC0sI1ixAcatIE7
vOJD4tHrhSZ7EWjFdAE6OYXa2vLeG76SpRmQYOyFc+eYf7ciW6ZtRQCxwhh83MMliVLaTkoqQdB7
pNr1NbbRUSQ7yPf7U7cNb67sesq+mF9kmGgyvwWN4BTGug6fVqkbAtZ2Qi8RNNY6tJoC8DzbkYE4
qYXeZ7m009MXNiNP1a2wwBYZPTs7MsllaDONmBSqQ7Msl/ooN0Ixlpa8a1apQUCoSRJP8VyXADon
GxHb8LdHbuBeQhJBoX0mAns3DqQnItCX9K8Dz3t4tM3PfYhggk3oGRXyVcHUsU2/gSXuobYKuZjM
0YDN3ui8qRhg/+E3ZUMZoJ445b1I9tre4RHV7qQCmtJnndcw7aO0mI0XVXyZqYuDFIc63ObEuKGS
f788ykn9Lnglzm3+bisjLNdWsRVJr0bgrP4e7LupJ+76yJVMZRCixohwmceff9mkf3mZiW3Hk0vk
UaVHgDzdY16LdZTjf6n9GNxXFzL7xC4TtFvDaoDe6ko4QyJfH91ox9vNTyFI2fmFk39IrnzystWl
vkBKrKdHy5DuAb5CKqu/OcYJe3cEcWnW/cpDOZYAoxtdsYQpZ1d8wW01RIyuLClf6h/UsSBfMx3R
kaNE+yRs31L0myUX/ZgmwYVk8DGGwso7+8o158sxqAh+wGWJQ6flebTz4bSerX73kMit23mNcYn+
6vyRCwNZIoypxJxCjgwaBTBcJ09XZA9h6kCP1YOmJ/qaX0Emot/kWNQ02X8qlMrSS5IJD0FH2qWa
mVe+tIvxgQ+w8VYoB1EqNyvCDiYhaYHRGulr9IE/E6132mV22fd3YOq5ROTHpbrXzxpkKvQqcMxJ
RoscCuKLq7PC+EjDa7oh+YPDdvk6eSSEdEhjPPQjkNH+clJakEZK0DGaEh0tnHwaMLy08KHMc00U
5xLHIE1Se1Us+GkTDj53KhoER19eeyogTkWT6tnCfGZNqSeGsV4axFvn7fr+crTYoUjAPpqzI/79
JcKb2lvnMPZT2TiCjGye470l5hO3dq7ZgGQ7cQJ0oCCeQOhfkKdpL1Xu4UUaggqvPea/ujRWapcu
LlFp+DKiO/Aod6PqXsITC3l75WoMDRmmqPcM8Z4pdQrJI57vwlTXkeV+415fJgpxliuSqvJp0owk
NrCMYyWcrKvFSEsOKh3PafVflAOr4mt6RX2vaJNg5YqyRVfYoqIDrobJyhOvt798hIan6cFgW5Ea
dW9EXVPPc8O3MarCi8x9Duk8mWmiDoU87x9jOtiA1Au39sJUM+YiPb/1WLRKSKbb+dn+zXG5joIw
M39n7XhkrkTUIGa62ZkZy5aeo2u/KVycb+390hIm2Ub8U5168Xpt4GkMbaoUHihTNrw74mXyZGxE
drIdrTDJU8+IW8NTqEwq74xUK9JH1biBLsSJo5gOPILoRYTV/bK7zncENNdqpe2gAr5ic4ORSiv/
tl5OFYNiJOnLTcgqvBg82ZP1hGj7dMjWid+f/S4zA9tTF1NQhcw/KcinEf7TuP7SaJVvrHvgn1Wi
OJRV8rcdbmWK2mbfxTSXR7ewKomlJ0SZm8L6t+TkNCxG19xj+P/0nuDoNbWCC4MZPxCoLucP0TZT
G3cyjF+E/g3T9D0F4PMi446BEXt3QqaTGc+gCzM930nT/irge2WtYukJdftRllEeenxOIDS9s8xz
0rCznZhtncimnOZcvRa6etA10BdDpe7wVBrBGapk1GDS3bzdPhBjlKyK/+PQTkuOTRCYyZ/j4TyB
vHeduC/mBVIVed7JMjOm0F11NQGvq0ROwftA+2Y5zdmW+8v6wNxIJsDqVp2KgJZ06XhRIZ8awWzJ
QJ1PqE38HzLln026KlPOa+nMz/klR/T8DZhgbwxjMXmfZf7R9yRUGgIQr2PKOfyyoTy289GO3ioh
JMYNy8fH4Pbvv4wTObHYr26lg7Z5gZFq3W1d/H9f5ZfHjFLSIYDOGUzzp6tpvRRqP2aOnwG31h5X
h7EzBfpH+FWFYFZru+0sKE3xicDjsO52k96j9i8ovJw6t8XJYN2AWgpR0VgRQ7rtHumh5G3qDF2Y
6bgsO/jGUvx9e6f5VDS22qCLAqDrCx4GuVm2jMqw7FrTeEuP8+SlPordP89EzOzSpI20Ixz93zVv
9hcu/NEm1pEkSiGLK3XQCpBZejqUTZYrZV86OZ/JHICy5vM/aLVoqxbPQv/+Sej2t9+AGA+T26Ho
QozovNin8XgsbHXWx3APxEPBxcnNpA1KSpn1bxqWLAGAGVZgvwiXX7VmUa7dDE+EQv00g1D7MDIJ
p4ahV0HhWwIpc2c9tQDhZdf4lvOY9GSPCyshURMWE+pI34/mLWo1aZM4c3eFGzEQnLFHf1SQi1pJ
ui9+S1omkZbw8gpPQRf/OAf6mheYQpeSw45fGPzReytuO5aXwb6KQq+kThKBIRS702NoPLGl6MDD
2T1iCGOR5MYOvGBgXDDqDAJTa59oYwgw9XLi4Y5MFh75s1NgIKBghovxuRV2Tk7EhMiCpvevHoJe
0T759tLwV50JTn9Jp/JFHlPbO6x8HRsH32RIp+RfYGn9AA+Ie1Z9HGjPnxPIsImPwLq9fBQdPhus
y31Jk9bIdKEE2SpeD4C5Q8E/8r3r/LSiUyUoaQK18QsTZbNA6saUjx/40IGQWc6lUqCbddqtpecI
cXjkHO4Odcfn+Ui5QeUuwT8PYm+pd+TAQ3tPhmlAxGRLR3VEvi/6cLF5vyT18lvMEnIUCi1cUrEJ
JdzlBvIXpFO6GBAbHIsfzdWfH6Cpe3Vj3yUjMssnaRMZvRcY0yEIc9joS+gt8PDj91SNGuBYPH4Q
2nSF71SqMMwND40jn9k3edyoJNU2ioNA1P/dGyyTDseNrh76SeJNtwnAANHi9vM/F3YDSykwr7tM
MIxRE5PCGCF3Hv0UQqKCPcweLh8/WLk/Emah0X1IfeyjsfoWHwDWXKp+GLWdqzaUAcMT5E/0bVq5
SUj7Rg4Id91heXPyu4SsKyBCCk41vf8dsabnmteCM1XY8rX3ubu+GKVsVGOlICo5HGr8iu3j7ueD
vdbj/nzkD8aaO+X/41O9Q/J/3sLe78BcSQ7PuwcegFXwPOch85vMCag9odRfOydYUSGBnIf0xcNW
HR7OTZ1+TLN6Oy1p3jcVcDPTFYiTEuMYg82s+obOjx49PJXZt5Od10Vcx9PXIS8am8HkCIpGWMQS
CTPpwTL8QOTS8kVy6+bRPPwpCYfhTpfhFOiBAUHd5QsQB5Q2fbceGdYYTgwkZvEPBZJ5XphKP7Ir
f1WLKrXzMZf4uPEHRNVmvtLpH+poTX5gTvcHiOAWMVjV8E3oMloudYyYreGTdUNq4lfOBneK7YS3
rmfktcImA9ap5zzzI/CEV/d8OeKO1/paEtk87C0Af3xuXayq+mik1+yWCYq9PBqYtZSGfPnfuSyW
+RFQo7ihygqSTPjP0gfHgcTttKtgNMBcUs08PB07TmHa0u+QSR/8Gn/zJ0LLvH9g/1cxxEgdBNk5
5f0UKSRMDUvmj0Q6NN3e7fQMomnpIDKlh6vKiwG0wSztPDp6y2uA6beKrk5aLbXNOq/3EBnfouFQ
NznJNwpG6jdnXaMAK9Qww5MRCc/+63RkytPn3EFieZdlhh4WcGqGYqOClOZ3iMY5rjE+hPTnuS4X
pPfMHxmLdq+d7nseVEQru+32h4bEOxUm+Bfn84VuAl+Io6QFX66IWQRC+K7CtZ2d5Uph+O69alx6
52N1gY2jJf3DoHGXfegMxKosjyKcLV/sLuB56IdpAV8tE5Hxz7B6obOFKIGFx/7J/HDRsLZTCMyO
b97QSTG585Fhf+l+gJyBPUwqkJ9ZWyY0kplENXbWEs3UpA6A6m/xWsX7h8JT60XCJur3C5obn5Kz
29u814CqmzxDdL9mtqnhQtXgL8PKrrLpjdJgFTIq8KABBuXsdpRPjnHbajURYPGBnz1rQuWUfVbB
2FYUmEw4gw+/C/I3OTe7d3DOA2PGO5ecdv+jCHRSK+fEBhry0Bu/9wLpWf6l2bRZF/URDBdy/Uxf
SPLYwnMiOGkZ44oRorb7tksp6ajONU4KjChyO31yPcqbmbWcQNQs/nydP1FFIl8AOyBY7F6O8MDT
zlGRbQ9wHiGs6UjsbEUnYeOZScXpeJBkBdPPYkI77O7PMgm3+1/iOlARtntfJUildtq1wI+3hRKP
gjjsYqBO3rCA/9emcqZdn4oCZdNOZz+imhZttvawEQU29AfPMfYNJtfMLRwJDXAqkCKsr/7Evv72
0QTIQYk5zDTx7cRzmZH1xtO6TnFd6rBfDqqrtyx1yEx7g4yC3umxrj3jlVOtHMKG85joOJH5ZDHj
DqW6guRcImuYg6MFCf0SKyXptmt1istu9b0HTtbNOek64TsrKqeCSFGZi8IvVfaJW2SRBMBP8hrZ
UwzwHF6B/CxpkvGoy+KxJgcUXE2WiqecyGJSxfTrMlY8tUTlyjQ87XdnmSv+NDRPQ+imYbAUEsZu
DH0Igsdue7ipvjbsHuf13pBda/+CgaGRnC48gMcjUHSvTyYNwZa2kOmzhKW6IwtOTaCT6LnNKH68
uCfSZ+av+9Ns2nA/N0M9ulyyiNfA/iMqe9nFqOi/g71oRLXFwIbQwFl2Rjy5VDaLJ7+d/I8zzzxv
SLH9lD7AJp827PjEmufZuZ984EnMMwdecC82Sb28QjagbpbjTgD7JeKKSkBbM2V1nWjQtZihIEzv
aZ44rxwqM09m3l+AP+EwR0lQ2II5v6bzwxnKWjJauB3QvYcStzNLrIp2LKvne2yisjMIsoQKj8gg
JcBS0C3ekjskmBujKDnXs5iZ4DTGQYBYaOwWQ+oy0tA7PUaZqwcONbNpD0Z04viv1T41D+jpI3R2
3nUD9dAPLK6KskLe+l5g1n0mOTkVCLxEtnJVjaLat2C37cbYmV2kr5rCu4bROwlCH8n8svdNCh/2
IfH6zxrtvzYyg7SScwLO/no12TWkiRlv3hvLdIi9wlq1Kf1nka20uXfmJMGr7s0P1BH8Kw19977W
CbaMUHrGd0TuufLxXXtOUfsibfkxlPmxXgaPjd5XE9BR477Xji5yROna/fPwG7T22iEBdczBd9qP
mVWn8zb99OyAmxobGQQzrSkLw/jkFpYMKI4OXIS/sDmBnpyuqewzKnnccEFLsfUuHzeOgHe7bOq/
hrt0ibJ0ltLobd0PQUO4BIKYJUNrmj9If7Rq9LTYvZY99jfs074jHfKNiAHqnuMTFy0u95Fyiquu
S5ETdiwPd5mEqZMACcg2Nxuq9nK+xYrkTHEa1SNoAg3tL8tpS3Vsg0Pw7z0yolTGAFIPWcgA4TCa
Uh9NXVzBce2zb3q+eTaZpT2mAWUo1SGYBdGrh0h4Xzl6ml4oSgBcMoTtnzLM1w+M7ssxhR651hiU
BLWP4S3yQBcJi0xfassnOr+qTQzuGXbDiT7lzmxy4RKjZ5WHE1DjC020t6KKODpCmzJFCagTSgeq
9LkM7KDYTLhY45wopKOefYh0+jPq/xZxRWoQxTw37Bl0lIGKm+v9AAqD67ZCEBkb1fs1DRaYo7Zk
Yibylo7z6lNw9huEHU9901UWAwqDvDkhuWGKjIe+8qwWFMc4KVKWySpNKzYo2IGVZ7LwkeMeq1Cj
bqYjFQab6y9UV9nHx4BFvMbJb/kHKQHkwM8SyTwb0F4qgctDhEZa8VzCdsZKJPJpZztu0a6b0xsr
l1Dig106WstxVX0Mz/Ginj/8/eGt2S3Rn+JYjUP5WROCPhu8NJ7n1n+a5T3b9RW5VBb43Y+2O7vk
d02EfRJV4dqRUXGdcLQN8nGW5UIL+Fdb+W54p7stTy9XVvNMzJnQTKsYewawpA0zbL8PPwJzCOak
+65hdxIsysrgVW62jX/oSMRnJgof4YJAGrqV1JkxCRqLPU4a1Ek0OEj31o0OEFZpPoV+o7jV98yY
SalE9eD7ZgGlK6AWt6NV2bbqhREUSldUkakbN4XEKCwn59ea8nW6FrlrQrZsxKdl22K4ufDY2XxI
450n9wqcCpcvov2mVVqE3/mfrQ+jeA9jX1ioRZEjdz8n+UqlY5D9+Dur1JQEQUP7FapXctIbsm89
X3H6HEQqiYeSyZx4E/UgzubvbEjKHJd7PhO+PaY+kg7YDKuEfNm+ljJF3cOr5I47MAk/k7xxuJPf
44jrOPD+e8E8bihcs1gcLeT41Xpn2t1DxNGRGqq9CH8+ktEt4bohJGVcSABFdOCr7PldOPuLLliN
lXHvK0ZiKYvuUXubDSK+LNPKRjAv60V5dZ3FI1ON5u5Sbtt+Uh6HuJc/3k4YtoUYtsEEsnKc5DpL
t60AibCkwJiqXaWtoUa25340esxju+0syxk/H1s4iNVreD03RUY7TkkdGDmAroOstipi9ejBXH/D
9cY8C8/QoB8BJ6jo3wxsodZh2Krp3MTw5XKNWhjYc8bzJWZCqu0Gj9oYRM3RU1XOObFpK88QLaa+
zAkLSKt6xuSg+m9TSajccFUQDFoBOFIks3jIl/vv1p70QHMxFkPEfo1iW76AdEATxRV87xbYw5ZP
LYM1aLc0d8/f4czX8hIJv43U4IB5f9Uux43NY3nF3ECifjuxVNxCJtzjLI6xJKl5DMVOIdkSZzZC
X1YX2r8qUreIe4/e+rtLlIswmVuHK1Z8AYfBQarXGtbbLd5w26tNuNG73GKy76Me9HBQhLwNDZ56
9/NBqjQLTZR5mTTVJcbHDYcCMIIjjFxc+G3LPB8KNkTVeAC783nu2zwVy4raCMFAE+1ZOa08fFKJ
NeDoKDoWxtRsw9zfMjyl2FWI9oIsydDMDNqUoOMGMHRiPBsrb6IKQpUQLR07IiluhFl+kX83Mq0W
NK9kW4Nh0FblJkvVqsgBtYHtyhzE7HRrPCBlNTpMLQgLOtL956oQOknAWi18g/5aPQsIpJZ304FJ
bSsu+lB/bUIr6rRKZPM5HzMhXG/Ts+9sy1TiVAd+tqiKeIzTVFetbqIRAxfsKI0hu6Wqfxeq0JuE
S32MDmi4ZEPOID65NiDtFLqNF0/QaKl9IbprAmbR73UOwxKAZoTFCX3r5krkO5jh5xgsJ8Gnrnir
8yjro8FT1UucwUSc5aKyW8tPYaT89uLptlJc7+bhA84n/h4Vlvzd/WaT9rml3VBl5I9aJiB2SQLF
p5Hq13I3JtBv+HD9RDY6jcG4XEi3fSUjVQXyn7SVjJhl6d4xLJXh5tImbyxZhaqttP4IWGSe05Br
mklAzSkYd1WXZ+BmH7FMC+sml4LyJtlDZYly2vEFWWqExR0GB38//uvB9ZoLSBUjfjXZHb1Dzdl4
LqTLUcWs6rqkKF8RETWnsBO9C+uVsC3CW4ezLQCgBgB5MkS30Nj9d/sJkT2NZhQKTIwqp7nHGl19
JqmiEM0BHCAxAfHiCTGhAXlt9Y5qhbmxS0ZtR05uq7kBTqflV+uHq3+aZLWAfv5+ZtcK8pNIN6MB
/tLDJw5OmyFsnX9hpg9uTvRsnvgYksNAnrikCp4/V6dZdfeq0tD3KsCM9IRDKATcgnbSMT/NTNbz
2gXtcsBidO/0DDLXm0+oVUxouVNPdJnDOJC5gpPB9/BDs7qLy+dV2z7RlJNI4uHLM3mh/uPDz2Fm
esY9OcuWo7OxGHw07qS1MX7T1ehSi4iGEUM/NO4mNui0wlDn/T/imgzZbygesyQbpLxk244G7I2T
ZIOfrlXgiB7KWY217aDCFnoS3OVBWIfV1jp1B5O4F9igzBDKEK2pJRDz1Uz6L2Cihqi3PU6u3W/B
FInlnicOk9XAJRM/DUwmgP4u4z8fssvRO70ElVhZaypUBVCM+HMLqvX4JHh1EPZWEUynTgFPdMZl
OQfI178E5OEVrHseNGRUaCAPusF9GzLDPlPM387ipwqHzOJ5tECK4ZHQyeC77BDS2Zmlx3Q9NGQ6
oURYmi5NHHUI8ZmzjgAqw6xQivlHft0sgQ/GVyisJBmFZrLwxGADoj21ju6unAwvIgbxF+BVpQ8a
hDY+62uA3jUtdbLu6M1JvHroS8jwS0QnkylNxAFBHtknIrgA4sqAzbyh6OZpoSjbrGotozMwPilp
Vex4v8KeyVmfklQDjq2O5exi3Yu5zMYsSDr6MZB0oyQ2SlNmUrIKs3YXMAgmNLawcIcLlLgN2t0r
1PFXQC0VZ2gW79hN6VjGv5H2oTbGfOEj4rNhZUwB4Cbr5Gdk9CuRfQaG0gD+BEkTDxp5RJjm1k3S
7+dA563VWNzPddANQ4TJ17Tz3LxFcaOO1pZxgiwrwI/7FoC8HkoQIIKOZIxXbmOia7vMWWjSJV9d
+ojxFnWHJB4rqvWtFR+X6dew9Ep0Fqc+2djz6rB3xZbyh826OqXsduVHkQPeI+5e5Oc60cDNWzZS
chRl2FX5+LASIDdt08m8820zBTyfLoPDzIyEeTTMZjt5FdMqYDTJCdT/yB21gqTwYGCzPf98n6Jo
9khTA9zXXoCi4OS5p6NOoinyaZTrh06yhqZ/9Dff1ox63wfwC/bKzwCGe7fBKbVsU7hzTpwBP/5j
3rjveY3KCEdx0x6Bneu5Fqr4oGH7dRuRT/gSR2VSibF9Tqw+so6kXHc3QD/eMH/QyqgYtmZLkW/l
aHedhvEX0oZ8BkXQii0AiKSgtzatpIAfeNhwSZRUCtpe2hUhxUgckBQNeVwN+yXx5xBq7PVVZqGm
9kdy/sem4YVSw5VqJ+8cb273YmnnYR07OQ0MKSZSro+u+kIgNx899/E8vpldUISPddTUTXpvidhO
W3Zl6RfMOMPy4P35r57EhFRJ8B2xSud5hPbsQNum9JtXdLSQmGxIEe9fqyly3LChUWh11bmA1uoP
qLHh4hO7Dle4YNAe87RN7GEJ42MnurhrDfOEYSNH/B3EbvgiD+SLFMQJgGN+6opDMsI2giIs3GyE
LFZC1dvU0OcUUP0lMla6/QLjjL/mOwNxjt0v7n69CkTBktd8BBTUQkJOQIIsi4/7ZJeqp3spbLmG
b/o9+CLlMwURgRZrZ/Ux1h8fvhLwB3CWqoQ3Ewt0cYC64S5Lnu1TSWkbce40zM6DmpXZGAn+pyGA
eJslxy56IB0laAvQ5D0dP/rs30D7YObbUyqYvdvo7y3tTS+XIJeeGifcd2AWG5DG2OwUeIA3KQXg
xNV1SrdpQggQWxGc6nOmb19K2qNlA0n5ScFfe4buERGXB1SkpGz/qK43zRmhasOOEm2tgsIAxAN0
JhqPgCSFL3UnyNYQkYibT9e0s34VtM5TXhdb7PVBrM1R3L0iusnkwzu69t4/jP3UTFm0zUb4/Rjm
h9JdIrK123bQg95QmpNZXlTmKDSHODXVL/bztQxCrsHNl+7/BjAFAepP2GBT8BhOgHhbOJKiIlc2
NRCRgzZPsB6SnvgGOyfQrpAabTQf/X0dtjYbj5eGywrOVmTPVNrchHc16ejbuJ7MTY3U8dLUVS9K
jZg9xgYTsLEJmbi0/H9a6JkvZNim/Aa+M1jtaP2eJeLtS4eu1E3umNfdBj1HE1g16sbpZ6OCcS0I
ZuhWvmVpolagIQpQGeaGk7bjWIK+H6Zyd8u1DFp10ekzUtAI5JBjx4J4r6k82OyVLIitEgAXL3Dl
j6nz0w1+2LesGS9NiAIaXmDnV/BWg8riw9j7A7yl/tOMALVy4P/Y3Uk9QyI5JAFuIu4ZgBO8uMIU
dshoz7l9lNRjoUok1m3ohO85/AyTDPRY6osmzmng/xmizEMpK1ctWVwzP8SnIWd0hPXbqMOlTzYu
BK3V+5jBTPJOxcnEsmUdq+2yHqSq1TBBxYh055CiXEgGLe9mk11YJHrooK5UxTJa4itiHqRuLcJe
2+RweTUhMFCcd4Hsnd3ANq1dGktog10jMw+LBMxDrFQ7GvsTL9rvFsjh0mFWoeKOWsLCRABbMsrR
S5IGoC9j4UNYEPwGRbxdIyGiLT0YV9CfpfjxC+2xlc2LwacJbyw06hQadyJSu1hPEvn+Fz//eQOW
09N/JVpaRkSPJztxjRB0i1vp+veQsFDlohO1iPyVK4fozAy53hKZoUv+l1d2051iBIJ16vlcnZsZ
Wcuaa1nWCJeISZZc6qlbTFZhQZfp7Jlaa1Ke2qKfnIVt5mWCPxecSPUCwuwcNUJQHp0HnFMPySN7
4TaglsKgsURJBa0XkqpmgOoOTdmYS0a/8kYPdxJairBEwFHG1pVgkqK81/9XJLZ7nw7x6eLBc+NY
jIpFqOurX7l8sbe++4QecUdjIhNAh4B1Z45fT3iWtllyHRCv16cQ2dek5LHLCPfj+YDS9q4exqOv
vF+toE5+5OgbRDOeqekDNBFF32dJQrLfowiQIstGzj44YXO0eLtTTkshVKUu2JrE4NXpsDBUggNs
0jQFsMk8PvEs1vsyk7O86dlFrh4MOlOjF9aKQBx4J606Q5lXL6bHJaFLZIwq5EuNZADNvRym+q55
Egn9nzfVr0JAIWlbS9Aj7Nc2CYmWINgB3anc38bBDXPUDi8zxRQYQz7agbWlEtiaba5q4eImpvw3
B0Qp3xQOnwcFevaOu3+Q+nRMTrBBeAgOCGiBkKLhKeNEyKfEsJFF6m4smVdpXGo+m0V5JvMh7nXV
v+EFQgvhYrLcqBwrYLjQjPwWyuuGnlW8DKrBzb3r2FjbPPphs6QAKgsVbVNfVgFej6qSWa/hg4cn
NX7sGRn4NRv4+Hi68tMcLvwlOHwfbpQBwLqZLX2HImh3EF2Gr2PTQYnG7+fMh1eHV0qoW5Eny95/
TPf2IacG5gsSz4DLU9/QJva0j9co2aEu/2TbEkOWeNEStvV6XMnAF5V0XdO18+7h2IRYuuulHyqZ
GNtXuzXt+MSRwhV7M5Aw154xSK1jrh/8jPMSUNA9ILDjf2MYaKjr3R2v+kOCgaehH+J5jVQmv/3D
FXDkl/Npm1t+5CysXLqdC/6jQ6tiB8BRve495nrWGPJWaM+iW4XRyVg3Ny5eS4gAuhnVFP615JEc
Xzx0brWrNqPY/df8iquc+4Zjl80jF0zXarBXG/yJC7D/hjAXuRN8hRQuWmCce1VD+w7+MvGYBxkX
WBCFaemrM63TnZxgo625TU8gfhtuQJC1b3jsLXqZlusC1XYVmZABNKrcWFpivAbSOl1bkyJBhpcH
cPrDX4rcrjsz4YlP3xE4325XNnmD4/7uh92/zqWccsLg9DDNqGDSlgpGPDPJ6E7Od+uMqangPUy4
x3ZgIOy8b9tTNg3Ah6DocbDgZdjImuTas+th2VGXTgcRWuzR96zTV+BSkdTSYOaBpyveqAFcochY
YM7+c0k9PR5Vng0bM4bhsJ3OsaDseV8dUxRMNCPstqcuosmWZaAaU8LJug+07T0oOQbSiW4Ys2t/
/5qhBT2aidW7kG/99csnluZEvBkb0VqoXhYLoj3Jn0SlLRO3KvsdF+5jWvutxOBenWD/nvawQM9l
s6aAWinjGpFVX7OjnVqikoVox0mr9wAHaQ7p5T9rZESQ6oQAoNi7HsLwjM5SclmVyXTy9jhBdr3k
j9Xz/PyDoTYW6lwM9QnppnEuwClw/YjKkYH0/QZo0S5ZSUmj7L5maFaeDa/Dgald5sIs0j5edsEo
I6WtSZgaJzZjym+LHbbfCi21bLvDsd5ni9szl9NB6cuKhhv9Ew6TYSYz40n78ZKKfxQkvWNcBOew
PAaKle0H9heap/t5duXTSwDR8La/ZhA/jTakSkX7Ka+Pt8Q5LofSILilsygstSCZlrCwvCYK5sYA
Kt9DWEeY9xihF87M2AAUpRUR08lBGgtYCZpefUx2qIfgUBzGYWAXEXgAnlKRh5WKdBok0i8kREjx
hGHQlARYumSGV6f4cQn6/k4/eETCk8AFFRJqaymbcPSLL2T4BLpjdXiyzt+6PUS8KavKhOml7Rgf
VXo8QhixI7Xmu88bZMDfCH7nVgruqfGh/QQTh0j2vmrkMyTu0xX86U6eHVneoT63onAYu8NOvq+f
XgcjDl9407tyyfG77b/5D8oIcJG1XW2oqNrRFlEtW/iJYIBUyMPiuJFcjLiqY5LGyPyqeKCu4nBJ
6AjrlfJ+wek9H6ZBKX5p79Hp4/xr6KNFHcLmEAdHmvBTwPSRcRgyz4zp9w4d9mydXkfA7fw41hUM
tBVurzoE/ss/Niui+pr9W5yke8ZkewENXFENAgFgEKs1jiiw9mtK8Wqkelck6XtP6fvu6BziQF7d
J+zwDqfrZzuQMPYQMgQdErVgbnN6Q2xXpAyR3CiPxQ/po+5VH+qQ+iOqFUquGF7b361j+8ttVXb8
WZtP7UCU5ix8VDdR39L8cwL3x03+8D7c+f5YOn0MG0SO7Whrx9Q2cARijfBGOjOPkZQA8TJ+iJ7c
rdJVMsVmVt8U037QJQdRgpkDFeX1hk07wQpjrlPt3BsjEHK4R6VOZjsaM5qCsoDl4xC0NyjhK/5O
mZ6BhHLz5WPOS3LeP5B2Q5c17GV3R6YyxR1CpsRCeR25mxUV3X58lbipBs+wA38E/lPSNJkWckTA
budkBHFPCistQAtJuAaTMLGRddwH7Xr55G/YHjDZfylnALYLnl/QDVqFBKlkT0wCZC81lB9L2JnI
MCy+EcOGf+6FCLEByuFKTAI97Zz6Xdj9ZZ/TKlx/f9SOrntn+a8Sp8Y71hejCsWZ96mhgfD9WR9z
zTJxg/5QRNLVbOAGsk3SuKWu4wpYme1LAPuNMm9qqVohAfCZAktlXogg4y4MLiwRR91OGcjSti+P
4M3DfGN24/+OvGZOmdz/Gihe9hfrQamESMMk3AV9zHqU0mgWPleuX4+RG7hpc3B2UWPK5m+aj6TB
2+fPv6bkshGxF8l/NrnW+F8Vjdt/mSGZgHILuvG5dSUBJZ+Ra/OHbvV7K5blKNKNyXZfaTXgqneW
Qa1ySvDujm7OJzkmWD7art88opmePN62T43g6HLttyLBv8s3lFXlYv2ei+dBVEmO7tjBT9IJPANw
FMlw/61+v+YMY1pwjY/6m2+W3rlqFQGYzmrQjXcpE4NVF4w7LZnkZ8i8/KYJcJC0z7IvtiNliOW/
yWCtYn8bMQMTeWIpyTwinzTagcJbJWXtJNl0Y2o8de+bKMmgCyX+avaqTBVhrabkYUJcX0POvliX
pzKihB0KPnrNC7/tBFYq9ek4EaKRTWQi+kcSapZSOB89hWbAOfGbq60e1Lx44KscnDPc5hZndwKw
RXQcibvJZU4BTOJYz0mc7i/e7ZoX+6z1y/82T02sM6PBZ/+IUcMz0x/s/zwJUrvteUsRYYpP4KZb
9/l4i/NjgJDGzd4DvImwG6w2+pICNmXiXy9+n65gQ49dATahhzPPdgzJYF81tJnF0E1cGz5YxL7j
1nKVOotkvwF5tpUwYyDNwUWn6SYtKMoW0o+YqG16KsTob08I8/9xRC1Mx8JtaFRSuhPsBpUBTDg3
glV90XkBclsQksIskoG2b7DDldKoj50trRK7gntzdSXxKWGbNYB9MIAciz+VhFUp3aqSNOm1qJic
PUKhTTYFVMrTPcOfzIoEz+iwT3lxQN5H5GgBi2Don/+tjyKuzpeIhSHTqG/+FlVcvex1BDoaXPja
r+YtKVavCbk3oVTJjb0TC6xzjMLAXUO8c7C2LL4SepbhSJ+yrIuncOjeVznY1ABTKz1mGlf21oAp
L45aR31lbnkgZEDWiXbFT/y2CfAY1UcGLpzDJIeD7FUFJxR3ms3DSX1EzsVA/KmU+FJx8kYcQB6Y
x46BPbKDqG1kR+hBheKvB5rpIiGBF4YDL7hnyEFDHgYxGKqZJ5iKbKg+pQ3vyoJyss6l9x6sWtqQ
AO40GQuS5Ev97szucl2YX+Gp1Iw2ZqVwSg5fvsrHheJoAlScnZo/5r6e8XoG4eDtqgeI+xC/rOB1
4AUW2n7b9n32mgJsaDyZn3kbuzWqj6Vn/adWEApAOoXjI1Cuo6XR7xDGnoLp1iMkm2Nv3Z85empX
UCmXAnfyv1wcokZJfzqVpmKyqNUhrwmNYGHBr9zFw5rRhDWdBTQvMzBFO39N5cUKPHROgobpdzgD
/fbTH6n5agjpHI66X7O2FSINpl106oMcdnJJE+qgNeAnS3t0pr44ygLgyuemcjS0dLbTDIaf1LOH
Bi1aGJnqYq1EeYh7u78zY+6JPHKgixm0XtPd7WtNFIndypjcEa4jcL0sTCUo5ROaSKLPZPesTlWZ
CNfyXL4gTW7HLLiMpNurrUBy8Yzq3acQDaALsmdwSNOph3mbTdkxjfb2zwUjCvuu8gU5ytNk53Pi
ICniYIYw+/0In8/bProj75ieYsnJ4rDHtTHUp5SeiwJx67sPZaRb2uvwSy7E5ZkP3sEBOqPmrw09
ep8/iRUoxQJWV9bY5hIWun5OWgVU5wKBlCBuIIjG1/Kcn8tffRiXTyuWzmRaCvK8FvxkDI/tKhfU
+HyXNzf5qPsRTQAwzYKyWEconNOD2BxF4aQ8EyWK7oLoDs42ax2csJ8muMVaInyRV5kXSjTEM0kG
GLWxHjpcEXMRgNwmjC5rA/dzaV7nZ2GBiCzCATG7M6UENf/FzDafIo1ms0G3SxNzNJAwpghRSXEs
K2Qf5EsfCS6akLQu608gdfMVpdOKqfERMyqkEuHfRpPHtcS1FP7ZFihRvKAl6YxNsirAn6G59kZ0
WgVMolIioEE/l0K93RasgnxOGavlF5bI3/KKPRwZHVNvxde8E9B5HvEb9GiGAy3JwH4a33zu2hdn
EACaT9lP7T0CvrE8sctQjr710XAr568DtZATY9sKrmDjKynqJ7zmwqdQfp38e9JJQwQos8T7u/e+
XticcqJ6z7IKRUC9UiESnLZ9PfPPkCtCqmo8afZlFX/NuVvAyGI6PlzeZOyJK6g4sN+denqaOHDa
i4InXIBuont9UbhYRy2AEMLGJJU2xmo3dLZLP6rMZDtwAtmb8eCf8XjbFe+s8eqmYRrZtzqusEgS
ooUi5w1XDB+FHgs4UBPGwUs2NcKtZvSdXMEoRRmua+bHmVU+KT3P6sU7uKqVXCG97RIwlofHxROR
bshtnPUjLiATiO/khH4Fhi9bHOdjNzP3vCann+l7f4NsCSJ8ma1khFKC2gfjE7AO01gLrAL/acjD
FG+yr3/WZzPTMPc/6PS9+xnTZi1vG+ZF1/2M3zLcDCalHlEiCt3BmT3MVPItNtuIrKo90i5Cq4p3
d1+aO5dAuJtuiJ53HRrpU9rWDZNdp+tfCzkujkE1t4RyLYt5s+pHsLaGQv3PUE3P49BY+l4mRR20
qi5pSLxy91q4Ej3AdhwDYTBSY8ov6tPRUK3SC7YG1eHtu4y5TXLAHoAqxP6lmt7XeL9L64DiNFja
My03FeQkJ4LQxcX3GObyiEQZr7RZP0O/RUrLS0PvIwSP/iwjownS4q2E5nMhh5uQneN0o4FBUf4S
2tdZRoR+qxVH5vvcOZ4wf4uGPOJzdXVp+Fu928WUdDUezYo5HYn0E8HDAZS2Quxp9mJTTBx8ecO8
5q2el62jHFeRnBreFAyULW/4JWk1Oz41tLYNZzc5evcP4Y4whKBiMHPcF92PYNyTF2FC4p5vj1+Q
BEmfM4QOPU0GpUxS6TwNL1u47LRoBTAisXF8+GcV+OgkYna9eBe76cfdP4g4ORd723xkaY6VhtOX
8hdtjDjtRK8hXWa+GTDVImnLwtBkduXGKVIoZSa4PcHRvr8noP8kJhl8zMM0JrhKheHQY2RVYFGa
eaFT49BW+todAiiUakbj+eTUKMDw+UjEjvLLBa2dlDMCOcqMtfnqHZ6hFYSkFH2cG1TNyIneeGBy
aW73wNQQFWivJRBwSX/nO/XyjIl6ZL9D0JNP7WbjzpbAqHjyMph+N0/rUPJvkB7g7z6jk2nsh5I/
SqWASBaIe/k9ZGNrLMwjDErBEB6F+i7E8qNw/760HtIuMUEhJ4G24X91JxVbhgQyWn4PhJ/Hzjku
j/blQTxUFYL5wwok0G1iW3zmOaUeO3rsfAFCA3plPSRkA0PEVjdARGpbRJmWg9eLTuHePknpAN2o
F9JDnHs2nggs7+2FqamrcUvyNDITTVb1hc7Jg4seinl0FLUuu+5+/XzuZuLKrj2A5EfpylD2aQZw
uW/rlul8Y7OLkE5m1VoFtMwq13L8+EH8AgEZHznNItwD2WGgHj+S8xeglh+Hk/e5xoa52lBvCMV8
6IVc3lnMN/mQ7NbhgEeMkRT7ULCQ5vOaRZeQ+jbmDk0a2CHyK04WhsmP2ZSoHO2l+cYKDh4hjVHU
5ri9W4BHTUJPfwbrp9ikArLG/aXykHbjgZpiPVuJQpHGVBj8s7zDoUVlkC3ebpVBMBcHzdjlVmYY
L0rvQCiaYHC9+ajTsYy7GbWvBmNqa1SnxVwUp8jC38uhORDjk3buztJivSAlzF23mz3HjZJqkQf7
J7lqTW/H2DFLzm+kqGnIvVkhvzysiwcVB4ZwavYRlEZDh2GFCBGV1AxbWtXiKtTH8K9rH0jpHpXN
P+qyu7fGtryg4s2k1ow/9S8T7LYC8cE5vx2HsE4a+3vjvLNS3a4YPjetDMRsrvOxe916tPb0IE0J
UDhDRv/9fA0EkUxOXc7GizfhQMK+5QN3msD43IVHDoUwtcx2xDnPLNIXVIUBl3tkNcbmQxbkPDdJ
8hIijQIfGBOJ5Ks6JXoLSM4K88G6hL4h1eKEq4In0VJLAK8hhrnXUrYR3jOCkaPsJF5q4gNwtB6d
oiGybvXlvp4BfZMtyROgT3nbuzZnEAwwbI7efXoGiQm4Ed2oPV7qR8Cxpxj/1jrISc8vJKN7a956
PoyOWLfJxcmT44FMxNpLlL+GvQOiFX2bNBtz3sMbgmmPA+fuaOlOnLI8VP22P/z3dtgOZ6AhWucD
LGd+m7sYEz6upzRblrlmuRIjjIcLIwT5ON0OpnDVLVm8Afj4RC3fe1lwZhPw2kv51XOmDGPpOfod
ATBt2UzNSWFWyhEaa4qc4WBv1EJ6epw3jhsW2oFpuWXZjNjwmPvuPEdAcXiDTQ+LkmeqitFSfgND
D28Qd8XP7IVyZ9t/3WtGG6xkfFvNN3Vl3KierbBeclk3defgLM2bbWX8OaKcSpVmE6HB8Kwo9Wln
W6jOVQwG2jKhNFSRtKa/gyaUa7tn4R0bwSsljbz1ECpQlPWBW9FchgQ3nC0DvVy0/drbbtVOX/h8
bHyvzhmFhWIr/QpLHAMJrbFhuIVueaCnHjhsNwIqvuNO19GeOF5wYFXgwj4XoTeqCYV0ueVgr0/G
4dahoh0Drm1/UH4K8QbHSzY9Z4aU4p5f8VJvSQSZ55dAhK2M5M79ZblOBAobhrXcXkSnsof5uyOq
IaL6cB/0IGQJUGhp3ak5JXnfkuecEQ1DVbabwaIq5P9aJ8NppcJc7bZDhPXpXr2zZAJ6e3SixKbl
QZsSMWLQ7HE5edhKLJqaWjuFt2+UYjIIasAstI5+6v+8bukBBJFKSo4crvzlQbtCfyiMsc3cUE+9
CVvl8GiIHBHvDcslVHKeIemmKlBbCwqcUVaow59LNpEmGG3QwgUxI0K6x87QRH8DPS7v8O/qns7p
6DbxOj3CFLkOiXl1/kffTJNhbUVGCDaoo0PH6F8NqzrJRPsFA5wV+IDAhN3HD1yemqDrMC8k2C28
sNBHLcEe+XBEkD/VRAODEogVHasFhdwjHZJnGK36rMAf1hAAedgCO8hYOFHE+mn1toLSjQ1zijgV
ch6+fRs6dLxLWML+tHEO09Uubljce4MyJAojJlv9RkvP6cgxwOSTQlP9902MyoH4KjUYfS3Ke5MV
50CvmrWST0WHlgybIuOOycOyCGY0JJhFHoSkh21N0rsk1fShdKNkNGq9FRCXcnAtRnQi5z86kgJi
izyr+Ww4WTMDydSZeE5TcX2YW6jWIcu4M5MR+SwmtAtT2Btpwaxjc/NiFhWhhGtHoikhOgqK2bCy
ag4e1682ZX+hVgKDv936ooeLv325N3n36WZ6u2vH9be7WBlHBHGIsboR52dly41pBF4CpK79GVdn
yEmm11Mv1GtHVZ+QRoJhCDcHfJH/JIvA57N3dfewxs7xmxpEsyWcQGT+ICuMuB8M3GtZ0rm7Hp4S
LHseOF7qb03yL8MBuNhUvP02GLDD3hRhFAL/nGHPC1ikTg19P/WtmDkgDSz80XSV4IjCis+YH0oT
r+K/cPmQvorQH+oUmbQCxck3wXn8HxYt2zarTtwZRWo87L2uekoT4A4E+F8dH6nRsq0iFwxd7PTo
3Zwv1IBdSEhQH+wIBcol9Mg4ZUtYC3b6+Jdz+ODeEP6odK2JkHhkPcj5p6t+l6WLE6v8eL+/7g3a
CX+1K3n1hiuRBnqB/6pEkeS1FZ/w3oSmKoR25s2lK/PSZJnBScndafvqqOiVwJYTsQBthjUcMzFZ
jDLvTvsaWPJM9bCKym5fkfCmn3pDRA5F8mea7wqmenXDstLcwhv6HyIobyW+cLt7a2gOee4QBrB/
UbbfUAh6mK+hw9nqu9xkWaeX1OiRt7cgqN0VIwifDpCXRWjrwmWFA2FSPzpM6tYE++mXHTwR4Hw4
25modWGQughivl9OiCddJcNtUqM64IQRQzyjEBZN8ZogFDkfmtM7WmuF2BDEkbF8HtBoxkfCacUo
DAv+TCCtxC9+LajexRUehssuTF5gGTV6LcHF+WX1oMHJ0poxQ3/sRwMAaheYuY0xUTVR1kumxfO/
hvH+NL7GRtfDf23xzova4rKKLcwVaaxMrk3pxNDiLRw9H/u9m7fWntvRohq5DPZFGwlN5lnHtxhH
AL1T5pXSbraMRZZogoV7Fx/jK3rH3UcLlArUc2Bu/vHzPa5mOlyGqk2/Sh9ieWWAbQA2CfMcNs/k
BIQhZmvUy8+ma2w9Q4/WLdJf3awAa1K51iRUZheetAEWebMZkKN6ZE1tWIcKJ8s4A0dWmul6Ggx0
LcpXQJqzx4AVVDo5hkPArOvWzfFU3vJ7BAh8SH6u8NEmeSkEWOZSfypsHFs2e8nfOJpZqxi4C1rK
HN4VU79T0eUxmbikblQ+PgjvZgO2k6Jl9c62iLx80ybqKEoUZDG+4M8u8aUXtW9liFQr5R7pHToZ
VE2zjHC5PbQcNPX55pGaaumCa8Q441lnivDAvjFAegKamtaEVW1F+G0uZVBB6XX6w02RgJMb9aa2
+zBF1vVIAzHNQOic8770tk9wfjdscqD5m/pG9/ynSGq3bgJ/2hkvA6h1qWBjN6lPLqN09Iztnp2r
FOIBYdW5jxAaCLy2jfgwqqX2ElOl+AtuIhKaAKCpb+n1KPtuDXzNZbUugp5IlxGleqk8p1UX2vDH
70PWY4MQWrcLBPYlZDkFKGykYiCl443tGzHnr+LxSPWv4n524BU5/gUW0B5nCxM650maIKMtN5Qh
jQ0zgw9yOkAxenj+duMi1M6ZA/oiwCDHCtcR8e+bbXZqtSAmEoOs0yUzoJ0vE7Z9L1i3on684sHa
R8qUplrrsnqAJz0L7t9eLDUDsVP4Rc/3yOb2DSycxmeDZ8VrLIbBfhkhViX/mTuDdKRyvfpnFleN
o3jkN8jfuz1AU4NnjJXuywFuOv9q0EYNcwoJOSMLBO1FmrfoeCF23UJqjjGnzi++9Y7jc4FOA2Ar
kfge9qlLbHdcF0CibKHpm2so+qP/g+OmfYKDDfbUqk4OVAtgChaY2U0diBydBjgzqIK9+DnuiXvL
rBJLg7nrayYeocQvr3utm/Pjm+hCTJH0gvO4DPDambYIX6azlgtl8IaSTPjGFlSDcw1zlzkHpZc6
LWtreSiTndST1LmTdyzmyK/+YvdMvsZWMGkp5DOS8nAbz+N1a9aosZQhlvmBgF8XfX1ure0G+OMs
s2aWfQQ/sZjuSXD5/smD3I4BLouNmtr/kebU9epTgxDiLZVnHgJ16wZXWSPZN6W2oOJMuKJ2Ztzv
ZlFTHu7k1qURc3+Ua5J6cNDnOSdlUfjGceF1s/uxrILaDyKeTox0uSTvhcHqK8bcRppN1Rf3KEjA
K6VPq1plRGh33RtfBGBQz+ibDLNkyRBtQx9e+sxz2LO4mUqRQ/3atPlu7seTCJ9y4wJm//G8V3Py
yK3CVREtCXiL5nBJVv3G40yoML5+Wt6LpHc2pP62wsHgvTEYrGUz7IdfbvPLqVBsjfJforDSWYB/
qRfsGj8yxLiacpd6tTM/+/lUu/Sn00nwSXN2lFHsLR3usjfO4MhykK3ACUGiRhfxWVCkMjjcSa9Z
pRO9wxF6jHcO2EQ3VM1iSqmvJv4q3yXqsPbaAwwGYPUGvH01DY8WR+uHJWRNvLTqaJ6jAYM2+sjF
XSmRD4MOse5us8P7dXm1NOTqfK2xDEfVR+ielI9mVKU1IqfgGxxAdTzTM0oS5AfL7uKE8eRxoW4P
poAfNyRTs/oZVkJN4Bt6YIYFuQxolyZ2AZeoO+eNp5pfkCwZmB0RV4GX3NfFCrG6/d6/9YkYGFto
WFTyW2D3GJNk864ESEf+ISIXyx++H3fs2GpMt4gZN7r+2sYpumhPgO89ulE1Zc4bHNnohcp/HTgT
qzTfdMKQRkznqAnBt0rloSYvb/jtB4jJHth0f3gR0HYBilW6xaetBAU6oWTj7XO32alg1XlzPq7H
XdRJQPgFeU7K0JTFrS3gKvBHX5Af+AHRGZEwKnwE/1L5N9NU8tHBx8AiqR//6p01NtML6VxV4YE3
XBMFIE/0I1PbxOcxWBjccogScPJ/Iuj+gZh/I3e6dVemcXf9ufWHxbWp6CrdLKFbb32NAPF1IuYo
KVIyx+XsX9se9QFqXaRADKI5Ky5ujPMzciUkXsp57HWKcTBmUsHJnmdszw/akeu12f+WVMVF4klS
LzEVRbr7XoBaAddaXi2vdRW4WPLV9VRbG93gJsXliQL9VyD4WTGMhzJgzky8qtBgRB/IomYYQIo1
1Enu4ztWj3LYyaz1PdwgBLis4tejpILMod7K2RQGl16jcaqjh/8CPZ86QMv+5tTpWxe7XpyomToX
BQaKk6yF1sLTYvpfDVgrPjrlfl2N/Mm8ZZkrCSAF/7E8p+FGpR+IoRhYy2oz34sK0kDidRFz+71Z
hgKfYVeGYbm+hG6wQ6aXVx+4WAJ58T177nVsIx66HFwNUhegRJcOJ+2jPz9h5Kw0meUHwTyUJ3OK
PHjxHNJIheWMK0QGAbQrFCG7hG/L2jMy3N/Na0KSGB4e4XSnjM3uxWAvsMXZrhVYPXcOw3gmxz0W
RPUeHgFpBaG6SJty4+WVE2Gh29fyhhJomfYYnGsweKVU+z4uoD9oHwU06aB+DJS6CNhSDYmmI2Uv
5jN1thYFgYnDZ5zqxKb6ryGfceuoZRyBA52SwoHqhSCkVmil0r4msPoXLBIUs2ABKKEUkClq23vJ
x72pOUqNlyUBrCXCMJB80Y5L0yKDSvpB1P349o1ai80cObs3wjB/5mcg0PXfpy1M8/zgDVlKcpGD
f74eiEO8FOYOyXY3ie6vRXUstGNvDyCqN8imQaLxDzRvgbZZf6Or0Jcw/U6kgCgv0szEREbZjJOn
TBQ4XGpvF7qNI/Cd+rGOJRskGg9zW5uV9YDInBtMLZwsfdHAtqlHGjaKPLa2hKMVaoemxHXu9Ha8
CYLDH2mZjYUftIArDGGW468+i34llqG4nXnCF1zKeKPo4+LkTHuD+785Qk8xXx4Pdal+cIDY2xJ+
2A+tYMmxRFyGNHilUx3QjR2za+gkZ3+RCyfDdkrjlf/wpJgRvrJc03NChi7jPARnC4ZEcHVWZtOu
5Q4OFoudsLSor0n/5KDe9OnM1fBCGbBx2ixofRyGe6/U1Ficcknwghg24w/imVL89EPAhL2OBaDK
9aeNTBv8v5IVcRsddenrqteOPLRhqz8umKwExOcs2KEX2IcaYAAOIHOYX8T95209HUvSt8niMQDY
3D1OpEx+jLuBdx8LC+MRj6bKsI1BRqrZ3gedOGFY3zwNZho10S9HuQ6r4gycxzoe74gYI8mJShBX
T2oM1IJVuGV5lFlteISckA563LiSPaMJqu6ecd25S+S/3BhJa7JDbgYpDLi6KqM0Kw5AMSDChtmL
HfFPs7DPIkRkHyh7NKfEVKXB2mF/htNMvhD9wj1z6Pl94NXmqbjC62HKCz2oWBSF2hR4iFZl/fZH
4IeY90wvNoeNCQWhIaDmCoR2YcpJ/LOSzaRLwLRH4xrkoMoypyK8jO7YrQiOlUXv0oATRkGK3ww6
/lHDiRm+jkTQ6vCa5xgoLjXhQkkeSDhuzfJuVqCJVZrQERqgnNgs9o194tvGepKj7NsWjB4nSW9k
3LhuwFflSZNzbCSVt6/BuDoZVJ9UDLULCn/3hJ8dp/EWIGp93gkGb+udHa1rHYTnLtt2QSRILJb2
L5EjW94QnOvLK16odoIxPiNOnKar8CEJwI39bWMwg8D/MVvfzMcizwOSx+w6vQuNglZuRigoB11t
YUnAOHHnqiZ7LHuQwU7LdBxeWavmAize4IvU6IH2+/ZzYD1e3xGOt66F/RG8xjgPgRZcdLqIwIOP
eDh614G5Kacaqs57ViUxVoBbdq/uURvcisrk11MRyUrpvhgIrQU5cMAjCRmAawOt27K+Hpi/OG4m
J/SYsANswo3Ma82wmkZGKAEULzS86oFITn1Tiaat9N+6x+fnZ5IYla/0tFrCbWPqvVt4NK6Jp0hA
ybOoGgE7jOFkVHSQpNj+0K6pzYkReVck3L2bYl/vS1jqCHbfnPe67KqLLZJ/6rDFxyJOvDcr1W3u
ncBwDQgc1jty7wVCBm+fu1VTaumUtd3oZpA5uKvMh3k2FVlQc2CLHe0ZtozABOM0xw0PdxFBj+B6
jtqUNP8LnUIQFNtwpMZq768iuBy+MQ9uonvbyKTCgNTbwubK9z1z7VuA5G1nrLxQlSE3p6Y1q+6q
/s+4OmoFR1yFvScFb/Yen/x+JLUARIDL4sxvnMIlzBmspUJ5e4aTny8RrqU/h3GUrxu/cM/WUQcz
dYezc9+yUOBtrhwm0jqc4gwRaoLJ2b1wGchGxLZJT1wqQzF7YcQ6jvMhYr499aixgWYQDDEgGKn/
d5YBrDZWHryiUrjxLjm9TobYT/dvXhSLvS8RXWS84eb17PSC4FalnKVr+QG3JNR40CRueekS4xmJ
DYQMxmJ3eBlCm9tZvzGp9vfBObIDT/ptPpCn/iO0i/lO9jJdgKrFwZJ/h1+4xkwE44LT9vMsFD3s
Toa1FbH9DdAKjN2Ocy90TnBgUiBouAa+L1/I06R3TA/HyFkdRTOOanvce5mZsSXPb11y6UaSD2s2
HiCAlkejBPut8gUDXrUEjMb5UymyKzzAsAlAdu11/QxzWc1UwCmAah+K9kGeQVpO786g8Z3zlys9
SRMaCSfrh4YJSXrWnXkUHiTlvIbHkNuKLpdOuKvZ6Ah/eD4xeoHjujea0oSBLs4M3ZqrKMCn9mCg
F3FaPKlqH9PwZPpWt8hFfG9Mtn7jStEYETEBdWxsVjrmJrSEbp74shhoGXjI9mxHweDZtmmC7cMP
UhLHnvs14ypLP/unRXY7oiuI7sOGunNzTzfn2WSE6Vaq6GgqD7Mc3rS9QbdriFiyYOa6C2SlATHF
CLqq7A69FkYE29dz3OQUcP1KDrk9BG/kynUV5K8vhYL8atvCXbXr8134ebCSSDO3OhEHX4lz/zJJ
hhokVdbeN0ABh3qumDLZzamhy6GSUvWL7PSPqjT9GYwu/Glj8hGXoPsRclgjJs4HMtmWuRYvbFUw
HeZVKfI/CoKAOpDjJr1F4QEnalhrnQqLpvkLitrUyVoEINTqMATK+kZcNTKKsurhBVf2O1LZ0OVc
v3yDVohgir3mzK9p+Za7yoU/7fhSnUDDaZzLmaxOCAoOT09F+ttknU2GbXdnMun3SyPGSGk98YD+
kPcCa7TO14rdD2QS8L8l4jWfi6tzmQRo7/WFZE9uYWKd9vNsF4CwOeRohvdQh0DAd9U9NNryDtnF
/+XreFDhYdEa73F2q9YyvLZLaxXC46ACBMkDlqy3AonDzERs4+cO8lurs2Zb06uzc71iBDp5FDey
BkCWAP1v4EVn2YbgkERqLnEQEG4ilK6KVMUqZp/fjvvzscvFiYYbb8ezW2o20ahpJ5MExVlG0+Xu
RqG+LW0oNnffQjTtJv3LqefCXTlnFPmJWi/IEmtGEXVLnxe5DPe8WhHoYNr8StuQg9rO1RUoipDs
6azgNSSQY3hRUW2+4scUGBjJeAeT4vxQDv/IwSLR92KfLjn7aMofIwvpgKhpe9lWeF7yZQmJC4vE
Onhf+YuZY2aXoa/a6aT+N3pbOMYqi6RUowoltdnfxXujcmfKZRmTs8ObCZjiIA1KftX8NfUrgPVT
K2B3mMwYBBcfjxs9kJcxwES5zasDiy5FW1AGueAAogCyk34Js8VP0iL5Cvx8VmlIb5wSa2m4Y4Dh
zbY4ovVZ9YXLulgZsMKnS0rXvLwHIPG0rfg00hfirIOSuTwTpmREmOQX4hJGDhNZLGx4gs9qASAk
2Ii8idVg0e0Stu1CurCNwkBezenVKLnR1S42WH2iwGddilIg6eSlyC5NLYkBHIfMfInIiNLLpTWu
EolflPtDrEUG7O38sAA+AJe4COeP5I4rYqNyPbaJpDwI00P9hzE0X4gxHg7lrgQNT7/Xgf90BQgA
JSPlBGW51j4ygi4w4ga+eWwn60yY1iEt6GSMYEPmvrOmvJE9nhKGiYBtbDwcJ+yQxK8uvGzLQG8y
vpVszv5POqzi5rnMku42AxjQ0r+mHxo3n1O9SRduIxxjvTXDWf8VfKHQWNjJWWlq2679qBhSoB2d
xJs6MU5xBl11y1Gr9ypwpnugyAnuZq7pwRd9z7ozf4O0Km1YOyEV2RCfCtPvSkfsgLhCFiy6l4oT
OEH/CrQ8J9P1Q2G99qbJDYLrdrI0Y4P2H6ht98qBqXnVc7qKmZEcGaUeBe2Q7nGQND5q2rut2fho
15fWY42XBdaVJvHc00d74akvhJnrsEwuhVDYoGqWh75qXXHgqI8FlmoRqclogi9oTSb/jr60xdqs
Q7VEsNlrLDPEBrvECFZJUOnPS93XcOv994UMcXI1ZJ1KfCZOk/8+Y/+P7A3aJU+MS+cFpLvxCYBt
lBb4lIOse9UiTjxymAcpvfp+T53A8HG9g4VyM5iU5xrbSfFvNNrPl7wDo5s5O+5+UHXtijjFsm3n
55Fm9g1oq6563PvTVC2vUfRt/4+7hzD2g/xQhif1LBYI+7CmGrx+zQdgMeVGlmyVxUSc4ZS5bPlu
gW/jREwRqVThJlyTO5FIQI1XaavHNwdRB0RLPPTmMnXoFz0DFtoD8S5LgJduHi5+JpDJJRIf16ax
JjpZ6fCP91djVDCh5oUUzrODJvfhC2QIW0LSs/oEZ2DF6hYMNIVPCZe/xqezZ39YuGwD5JCZr0n/
rn4orrUomru20/cdCwzPwZyKLVf805UB7BEPh0MyC8VigKteg6V8uQ4t5SZKXIPege7LxwDk5zRD
chXMffJX1CBvDuMS1MAbikou6cQmWQjQb4ot6P8JA5S2BdaLjCbuebRnjxgiTabmtmUvbsigrx/J
YKjWgysrbvKgCX6RSvYnXC/6w8Rm7Oo0SQH56cA/rSvrfhh0ItWOHyyqB2iKPeiGkJcraxm/S05B
XnGY7iApdIlm6lppdJUHn9rnWpaAhFwCE1qA/vY8Ul7uGJ/OQ7SnVaW1glSl6FZmedw8IlZilgT+
q21YMc0/qkDgTNRYNyBbFNfydmecXExtq1uHLxNkHcNVvDt92Uv116T7S7GbEzxVmL/9Gw4nyirj
5sTJzwlKFVAgl7Zb6m8hp12mVMqAyBPNLMN1Rgz6jkEIETpOi6+tyEGoGpzQAhBje9nPT3ayHXrA
QXhelYu2iKIGksLDKiResGHQRHumh7zSndFrXSkaRwcvASELQZR8UlVMi+qFxQh43Db1E9Hi+4fE
j+m5Vyx78XILUhNfcA7QfxpK7R7eonODKnVoW2wAD4Xxw8kWyhbSLSgshtcHr8mWjnZEz3zU14gs
D4A5Uq5mAcXYH15i3b2kj2B1sn1yedKyeDML1ntwBn1YGMZpZo0mMKLoiKyZXTmHXnSXKkiB1oKQ
5jOk4lGFI2x9sjUvR1r1UUFJh9EwgSW8CM377s0POcdz3OZ77gOtjOYAlI3e/rcKSB0GdDQHceuP
SJdzhlYSb/9cAL7iFDQMxMYAvC4BP5omuAaxSJeLrXbgjrD8fiOuYzgOW92l+gv/OmziM679DaL7
oCt3osO6KHQ2SHCKYo2hsXSB2LWbTWkt//J8ySUo5qWAYka+UAMxe4GZKKOsJFYHjs8EXaMUH4oV
AjLaZD3y+PZZCgUHnPxMRKDRRDAw5eD6dCjB1tCsKwVbbz0EU0hb2so+UCRaTQbGY78t6qTOyZVi
sysjo2slnWfEP1U0EsJLJfix5vo1UQrixsd6SykvfQPzkU2IXVbobHK1S3X6vh2/4RgwZrDwz4BV
ZdjpRDM11hPUVLNv7CBeLZ/u+Z3fbwakD8autky2SIGVkyRa1UpsQ85A1ImZazEckCZl/nv7fISE
EuhTTOs6s+beqAUffswiskHYdHENsVVJdNkdOmCY8RJRw5YokshzjvwscteQqc/WBT2JP3fGYgY/
QlhoyEj67eDAz0Qb6ofN8lDKWgiN9GjqrqLbWq9oD8qaoA2QAXsqtF7/rDjtpmFQuW7s6FNb4JKs
I5G77Iyu+temTGKEDzrD5irU0CLBGzwEF4rzVllT5pZFppnoVzOyimZ3Ipqh886dsGgj+2Lt8mq0
2rz+hhetMtNW82p/yNpwCj1VPGz2CiFUIKe8p8u/0sJIINOVU+hC53DgPf+wvLfhnJWWzopvxlTp
C49IbXoftQXXfe9617PqZOetC6bULyt3dGkjgx/D4n1u0GaCvG90pcPbhRC0SrJz2R6oNV1ifL41
22ErfQg1wcf1DSc+1bQzflyhPywxQSfFUyVSuXTh4zn9RcKB480WP7jw+p3kxp1h1UXJgbVrwVKe
xl9S0n5MqcH0MthDM+H+9LR93DVf3+x0eYBZR81nG5JWKQmwu0kpGQU2+Mya9UKD1cvh/EOmV1V/
2+Lsa/7udqgNscBDNNAEV5qL8zxQuXMWaOhXm7iRoxwPa9ODZHW2C+2xOR9A/qpQ/c9ZO7WzVx4U
FosluR9R3M0CuFi/LQn5rrzQDHfefzROmzgLjE9su9VTSo7WTM1oHNdTgh5Na6QmzQQj5WDIxCHH
BhX4yleYHbN6Gd7TXYFgfjl0uGPYeX98oteI9uqAGsaUptxEVlpA4yn7rk6/iZxRaZ0BrF1dwnPQ
hJjspCvRDeE9QcE9R4v5jZragF0j64hl43FzoAB8Iy98lcwmOvVuIjR3klzhTF/uzKBW2O1AfVwL
78p885/Sg+v3rnFhIPdp7rlLc8NzIDoJY//9VRs1T31UKsbdCh1KAUU1axj9m6fJ8zov6IeHN9Lg
stkv+1sdODb2A+C+suhO1+ixgLu2YSTsrSzaHexvdmj/dU+sgf0H0E7WVpBkIMqovupgNlsxzmwk
x7RyoXjNa2YGiyfrBFwsGCtZDLyVbFJvUoY44/tWjcYVUOy7ZGrzutPwwSEcCM/ncHvgvbFksk+X
zzaiPpYX/8/JncvWMlzn9t/SJMdJh9kKohezmY8wyepiKHb6Ng/D+QBoo1cytC8PUCZHyae6Ywoi
GjADG+zDz5dznyTbhwfxVf0NGygcvsijPKW1A8FkjtaMKGrEU11Y86geSH/QsqYfxffLgor4c6zk
Iid7fKLajKG3m2cORP+T/nlAv4y1HWupYykvwuhh6pcfxvTTE0970f15ZTI8ZkGQ8BMPdvUUMbD3
6cSA0eIetdS0HChRXDvDLRwZwhblqkccWehDz/DvtK4QhWQc24X8P0OdR5Tu/0NqV0hjn9fWxhaz
CzHVOpMesFdaKdBnvC/rzuQjxb5uPc0j7lD5iLwviL4fF53EEX7k0Ynle/da1ulDNXTZeiAjn4Io
UPwxRMbLhIJm3sf0l/cDvJNDII/D8sskpbeyk30o5h8168uutvEKuLPfKdUrGPWTzOfu9DBtNHQ2
1nZXdTlsQqTM4Jw2g9ds7exfxvkiJ/unx7FIsPEFpKCQ2EQMgNyJHxogjb1pGTcQdkaQPj5RaJ8Y
EspA5dO1fv4SYVBhck+eMkio+tUiO9v8dnwxN9nCawNnEMOMXw+I/lOeGBP0MmcLgoI2ZZD7A5aI
+hsXGJgQMNO9hv/88AOXk+VzRiHnlOBOUvs3IkBzEmm86AUz7JvGAbqV9HuWxwgLTTgm3wanzB3Z
0rGCi6pYqHjSYF64ovSCQJg44eKYvg94/gr+KlsFoyQRbl7HaAIjHnIsbrXDMQ3eRWqr4QKeHi3g
iS13S0ZwkrPBXSyCPEpc521c/DYrHSHPMnLO5mqWeabhsAJclP+FHouzEL3j0pN5n7ZSnz/uIWAD
W4jfwmDH1vJX6FStoRRWQBPhG1UaLQAlHhPfgbv7TpS0Pejf99mXkGSNURWmUcEJKxsSh+6zmgTG
OKQJltP78zsWQU93GXYZ41m2LVt2gPUm0gC5DC6fcz4ipqkuiISKNzim9rnhDwikUAbXMwlJ0dd6
gn93/sMBqd3n92Lt00qJcluwFZycK/pUCFvuQJTwc83Cg0t4rbbE5uxxPNSjr+nxDKEk55uw+swL
VGGMGJZu/VULnQntseT5cceZknlIAZGF498O9rJR86MX6dwxOw9aaPXlbNBE0qQtL/SJmgu5UPpk
gRRL0In5SmJnfhoCF61yN5jPUr5LNylTtdDM5KMm0FyQq8AVAaWm9b1RtrL0hcF0dODWjKCkDK8T
qZ3QqyZRk+puhuFgEsCnu6tuG266oH3ZKQO/5gixeueTOIB65KPaqbNu70+PErFjehWKO0Eav2k9
ronzbrVSvHcfMzLO3HPexdB3cXWfEcw5s2BQIcdj2Rqkomx+8SyoZZB98IsjkDPtgXb4UbFHvx9F
ZTOKQTOsPAPaZXqU3t9zoYcaHftK48/cJ/MxhEqhaeCVoTUCeXbJ6kX+V8eg+Ny08OmNKrW2N7qi
/v9T19BqNDD4qJkh4dk24OsBH3qXKqdVKatxzV5CrD3lzqtFycqIlioMPBjD34jhqpoDx3MTPCWO
yjOgsDeyIHDzBC3LJyPRez5QqTW6XyfUU4CF1ZmoasQwz0G3w+MuJx/TUg9H1NFyZTsLQv1ieDA7
7D+eAT3zGS4iAlINAx6PYioJ85M+Tc15Zw0hE+5YIV/J7cp0emWLECxbYZQ1dxgJr7x2ntyeZ07D
Xwh315M/I479/aMLV+VqoJucRm81McnV+8Cak7rk2eFtLB3jrk9trKwGZ3GOhMk0dk88SpVys+Zu
JEC9v8MLFLl+ye4L5o7HEVcSQpD8dIxBbQw3rgQJ0FhSUQk2ObbqKMH6YtdTgRLABbwuEVUdp2Qv
RE/qPxijfpf4oDKh2viYlzqZrctBUNsVx2dJcrJQqNXiUtVW03l2GqxKU3rcV89R47GivFD4D5G1
qm9RSNYzSKVVi9snM0uEVSNxUKZewLUVk2OTmWXtyq7CnQSgcrgmxgSGgfdaI/Zx19Vaxg15klLM
NDN+kd04gOAHgEWHBk6VfPBRtkoK2+oZXbbu5PyHHPhE8Fj/52dQOykeXEmOJJFaWUY/0oGUCL7i
NlxcW/L4YVuDGnu8aBUMvJc/tkzQVJbI1xBovm+EZ5QqS5rSjqEtFUOB5fKZmybUKb4wWbEt4gAp
nJ0Kdso/dXknh++P+LlgrJvTsi1OHpP+bjkiL69F1z5jnryCWaauF3kLR3OV4xZe7WjEBhL25lYi
8d/+AGcT/SlRN7n0eJp1K5AoIdR8B4JUuFuNMkIpDdVaQPHF0DecV8nvA3mxTFVsmerCtKcduzCS
hP+XRgwnhNGRYiozJlb27kPkhmRSgEeepcq7qXghNZJ99cvw2BXjxnAfpCMxG1K7rvF5OqjHEQGW
i2t3WSkJC/bgPAKuREYopyxQ0Lszv+pZyEz7yVLyCjH9cU2EOL2Pv+LzM7hN/6ivWk9xiiZsSbSE
kM5XZtZBQZGEh5XHQG75ug8O4mO5+M73JvNpqR0uANGwo2eoBPYaOtk3JQTFIYch3AaSqMEYim3V
S31WW8C+094aQohxp1Q5zm4m9yvHNQOBMMbuksPT5oEr6psaEp9BUYqKgdq9b5+f6gTB3DeceN+4
wUDyTI2wOq+azcCq3+LTvZGEtTuxGpC0O0hhAW9RLZdZucR4uyDR7WxH+Xd6hPcfHDG10vRTcnU4
DbeC1CVBfOEwJ1h9vC69q6hyMVQd3cPH+y3drp2NdX+CI40IrZnw7AjlxAopfg9QCvD5OYlc5cGa
F1XKgwuN4tEbj7W6HuUH5NqY2xddy+LwOFY14ZRXgiBgWUw0YP5laA1TH2c4fwa+WqO26PYOn0nA
7shjZScMTQ3CDCvfCQIaOvXKeitqWdkdSbvYC3AvZwgW+RzJVm8UQotc7iPhlmla6G2xRjrwEjmb
XxyKS3etwq6RLb3KNBrTxDRwy/PV6ZtL/lxRko2dbEN08D/vnNK7CCWbkSiZKAX+tnVkyJoRts/Y
ShHHHgnxBAHbCoI5G0r7JkNWziLNSkdFfa+sSXeiyaCLM9zD26+GtQZywzJMib22fIgv4huFSnFM
KOMTlSZVzMu8NWUdPkbRtYmgPoPmMZRDdP+jBAxBFLBt9Rr5eNHvtEJSqlURzkgAej+7aY35O0tY
YbqyByMNRjN75V1HaLAQ0DQLsL31t+1to6Y9YytqyGaD4/ZTaWaoXRLM7XLZf19UdNQkOffxsBGb
qmJ4PNgrCLYt2L6r6q/3iUMBXVF+iplGlEQoIj/G7hj+O/8FXJdLT5wYjgBTDkNZnThxmaJ1KIF9
JYmDgCqo4RYEEh31tZRxknOdfoHaAsazyimZAmvrt524/UQLnva53PgWsSaojpZhm7ocuN5+7aHu
i06T5rmlsO2aAG3PEV4caMO97pM0VrVO9CHacxbSKhKxzuUNQ+Z65xLznnNO8mz1QltAdFIDKsBV
BXx3fgXj+PFBnAfov42tVyK+8DU0PM6jNn7RyHS3kER3KVlI/meU0XFPVRNQy2Mn2P6k3JPLoa53
+3pnc9YD25gMgmArAvNBuv24rGVW8valsgYFxRe5YDqmUnY211Ja8UGGjh24b/B7yzYPrBcZxonA
S5dW+mYzn7rxj/j4JwFegWiNDT5eU7CYgTm67sm3+K8ZO41UqGWOqmOHLubHQywLVBxRswkAVk7D
v1+N/pzcBTZ0zYM7BP3IoM3JNtTmeadfscmh361sCOVH7QcQX66vCepctlIAyEPU7/xVb+V9O8Ai
nizCumgB9X0KvXa/gNCrzxchUEEGyiZwV237h1SOc0lvFr5HPB2Q4npgaeegZD6PsHy1p5SW76zH
z+BEOL0KSh9oszyVnfXMq+MR0xEqkK1j8u1V4QZiNfPQy5chPmKlTNx6iokg0k05HObYMDgmkr0U
CP7ArDbyRQdg6djvIBjQ+Fqg07XcQktABivQegtpuZp/nQGd+g7pwctqYiHu0KS3IdypYjECBUIe
qNoALvtxFF0mq/lW2NOCgrFfe5e7pGQu1a1lNwC2/77uDOerBV/fJvAlpozwqPM7mIUtwoEz+sXM
9dsO9gdzqdTr2JhaF+fsS1i+6leH1+x0NVNo0kzGpfhGfrEcasmhb5xOIXXEIZljer9eHJJeAfJh
zKEP5mdahGEJe4JewOEkSmCzV6Q+PLW9FWE67d02GCJ51kuKGsaQqw8ukMgrGVR2sI4NQrUf5+CL
jfXKFzOHYOGQcp08D3lDJ3yKRWwnZZTuw4QM1vUVugjfSc/kbPEqYTO8UOnIDlABsH5rn70bzbcW
4qSP9CzBur5PsQRkkvMJAOAGLrwwHkmbuON+7wLp8wjQv9G+c11gqreOl0GQ3tnoLzbdaYO1SCvU
ENnb1ZheG81sVaFb+hgFZZ/tN6I14ymqM3kl0ZLZEx2JB45mIlgveij+BBMh7u6gTnLPsWv36LiM
5Z6/X5kACV7IbYLEnV7l83F5cViPdOlLZGCJmn9NNJdShEAe5r1iVY7kq4UG7Uxo09BEK2gP8XlR
Xxt6df/xugy2YpS+UWBhVLU2aPQkDkkjXZBqEP9BCfXub8ESPmVEJaB5b1KRBt6rslIryakSCWOi
YQh9ttYeom7Zo4dQuzYHMk5ItzopuidBqnj7n46NSct5Jp8yiLfkws6J+zt/K3WE7+jszjXWgIBx
shiEwBy2/t9lfBxzwfBbYWqPHOwAUjBmDhw7GaL6OIMW39fP3UXTyDuYnbLb0cuoDaH1gOpxLJZz
Hy/akbOYSeiAIrLtcpTXV6HZ9XgKpzOBR9X2+zyczGsk5KSWOjrKNGqnimoxD5M9jCn/sMVFk6mf
stghyWVeIaqA9iaShbSgkV2rLXQ+UVWFPiwQ+UPmBARzbz1GkQ8EY82Lrgp42IkRiZU0Paz+MnV3
VQf0bcJSm8OusvEG2nO/NbWVW0A3CpdAroUpsQZ7CVtF8UYVYV7AdSLYr+y1M9cuSFCb/w8SYVnR
QLLdojripWastV5r7Q9nOhTMWHOMix8NudBMoe6RmoZq9mc0Zvsp1HG0vNP6JdOrvNIPQ2+8jTn4
/OFgprn4vhUFETm0yiexsGBlpjQ+V1IUNmc9M7RiNZZ0nxRYl0ADUU3oP5dl3ZGxvFKM9s4gJRzW
vO4HJwB/wnaZ6wLEToYGsm2N3ygryWPypn4EbtSmuyeEv9FbIjTLzdWgXFeze5c/mABI09OWXUfy
DoiwqnzqeV+7s8Ki60Ai2TGppJeR5wR83L6iqOvaxf5/eUdGBLuxHxSGF9m0Rfk8U2jjXL+75zWG
ud+oap7bTExmoPdLS+nqd3X09pORZm/3sJUKAFFiizedYr3BWNokOe1a4V1okdTvPkJxPgTa3pmi
PSdTyDfxypzHFYkOIIJ+mDbKKM0/twxaa3sT3TkWgLpy5+iJRqmBJvJGxu2FXenUQAiGGwcdJETF
kVuGf+574E2hzLKMdeFhavpxHCPxqFMjsbhvu2NYIUGNn1jVUg/3olcBLKz08LMHZvGDXMlLt6zf
FkZauhv0ZjvYYg7r78KCFRuUSsMHE5uT1B+tSZiE9td4tIzHSVnqfd6I7OqP7K+IfIvTekNYLeEn
g4EXl8uPHiYPMe5148zsNQtUrkb2qsvbo+3MwHaPbvibP421oupCA9tMhuajMpZt8g3MXr0WDPID
RFkaW2B6qATdhY9DA/YPw0cgOKRhiJuCU3SbfiwU9JYD3Vp0UOmn0Vll6VELCMfJtkXjfn/oMKOA
qL63lBR4J9JFJZWWDMiVyK6HHF587iX9eLr5MB7vGkSvg9eJwpVb5s0yOmRHP/tLdcsQrHR79BP7
EfdvZRnfSGN8Mh8uO9jtE1Wxx+anJWYNHqpp2bG3fgZjL+CRuVXwvt5WL2U5fydep3EgcdW5WwB6
ES63mhhCgwVxTiVCAeQip8JDXw+D8tE0iN1aWQ2PTHNnK/NjorkkAc9oZr1pNTj/ozKy2AWhPypW
atfnOFx0AmtF+9wEhh+jbEuYlYt6xkqp1rjej2a0beDRB6mR0bq0Nw8FgtYqsQcHGH+rNUoQYA3c
fx6sQxABg2sHd73w5z9dT3zD78kEyxUh1ROqsJXi/lRoX3vHgBhWqHhvmgfckGVTMyzY/qonjtXP
5Tek0ICUjuI1ADGrTqsGERRwqjgP3k6AJkTYP7X1ivO6gtHtnx8CM3fgkxII06T17nOwcfLJnWMR
k7MhG91Bx64jTV5f4ZPcUX+HrMUQ/de1ewSOPLgQKcldC+ErCXE1mLCv5gF6sFj1aZcRuacB4ObT
W8U69460FjtSb9/HFeOqbZti/MlZtO6l4zhygZWF03OYAq/+/yXYU2aC4k3mE6At+Di9Tf4Loy+Z
pb1TVEgP6ipXIqBofX6Oh/m4KxwIFVueCeYj0eX1KGIMcrD7gb8TGHqDf4HqIBVDOHzVkcyC+N0H
9eeuAxbIvpVbBNzmwtp4cUo3s2F5Mm181AZIGqo72dgq1Kh10pg3dI8dhYgFSrlO7Yv5KmVcPf2s
oilclfR5eD/GEP4DNAD6zgkSnyGoplnMqhbmTeQzP2UL/+hBBJFnUXPvpx/sbGI2aHSUf4FwE1AF
362P3nVYIw/zKoegJIntCRNutaf340bdnJKezA5GM7SIUpvqfAzDun4fqaezckaII9hUJGZsINB6
TGUxNT0IuVO2fHxIbIeghpf1Yldx7KzOjjIL83zlx+TYTQ4kSTQgFQmloQVvko3/vZHBL+U+ga9q
nD+Uv/bcOblza+xH1mTC8U65Y3GZIGBT4+xpIcoX1eHGLdAjbYKqBO5YMV3GGxJSaHKecJrMtPay
h7Z3auuvcJtcADHlpZ4iyLdEUbodl1ezEmx5ZEDtEKnxfYc3WvSDyB/+uvP3u8pZqkgN0gX2L4v6
Lndpa3F01NgAFhVUAj0y6jzB3bF4DW4OCFe11RQZlNdff4l+B5VSRIOdfG+/zI6R/GPbzN6EwJQi
xENjVxTVocarPKG0jrgLTmJ2piqxPhvX0pBUUyqVV1bQ8gTikJJ+Bo0eBoz0aekOQw/sT82TD8Q8
IXq6KOn3lP8bjx4PS0jsnKV5dOQgLFBB8pEC00ERzgRdhHqAFHEM/orat1Cfdul/p5bERG9DnC25
0yV+dd1ujlO9ZR+jPSyYi1IWgbwroCoknTwCkJolv7O+XNYOqVeuCFqs1QqYP/zON4WSN5YmhVFL
DCUdWgzXcCcYO95fJY3LkAasvad4d33tCDy4HQVx3lKKOM/7RUfYiUQbknPRE1fth7MyimyWy8FF
JcpLVmPTFRL5clme8VIRYGx4hgIQeb7m+1sReplLxw+qCXlbGHogVgBhKy/PMNQ6rRb8IFmgzMLN
6lmoh/H+Sf0jvpeAm2QCKmAm6Ce6LADFjrbD4ZkvfgKo8gI/tCzfP9Oe3MAv2l+PrsRT7Cmbtt5m
L9htKsIbQFgyDAukc4+I3sXRgBI8qDJeUAaUYnI88DyC5KPRxljP9oeh8BdoSuIjj3bojTBNxu1g
//poMJ83gcooK9KFrq3I5oBa7c4aiNveDkHzDwm1W9tWJfq9ihhmFKosX+ZJdypQ6DYQ1U//vpe/
AicZL9rDO7z0q8LfrDEJ0Btj5R4LScmW0Lbg9vSCUu0eVeWwi5CKJQbfOokKyzsOVNqsKZ8G4rgM
OX0vjwKD0JB6u4gUdESEYEEOB4XazNHYyehSKFgRg9JOKtS/Btf8938XUeFycvOO2mXwmqQn2fAf
lqHCFZ2fVBJFswzTfW01coNp665R7OYCD2apD5zKk389qeqS9gmg23ULkW5d+a3PnvGItKK/9X60
ozLIllqkHJP74SR7F/FiAb2sSxS/9gdPmAP5921nCdo0SsWUPeugjfkkFL73PvyU88dt7HAGwtAM
8S8KU1T+fOiGmLhGd3QEJn6VeAYka7F6I30IeA4T2QFXBPn7iGoJXrVmuHWS88ee1HwX+VXo7ney
qdbKaeLRpvGbwYO3qtGDgzzGQBbKl+1OVq3nC6/uXrc2E8ptBqzihPupZOG8cNY7Vi8TwDofKcQC
k+4qpRRrqnWXBDrBUMXOQzIWG45S8j1a20vQZFSFchRFzyXGLSwr/yeDDMBQRfoinU/9DHHPAwbZ
7LlE3G+8IEr8CBPCXKUB6zoow1p5lozJweKfpoDp3Eb8jfzztlejbttyPi8B4ciZyqRSMjBKVGea
AamvdKONHee7nqFrAGQUSNx/YqZcTxPRAtGsUy+U/iBXl698thQd+d9nmqnME6wvp/YoqyZY4SbV
kGhl1WUAy2v/3qYLddWIGMi+zvLIpNlGAVQ5J3CTyaEA3LwKLw2wcuaKknjQaOxuRmYL0WK3TUFQ
7Hyf0NRiL3mIBD9nh/YnCUQks6ah8jjwp2twTP1uNgyJhjTrPxYveiJRVKPCl5yNBrEVme027t5A
Go4ow3mlExtuO/VYQ0vDsd/qy/UNl2+8SF8plCovgkTHSMBfovucgLikAHrhCcWJ2oyocPhPycsG
a53WFOGoeOe+xe4BdFqpVKp86I6ulS+IFh1Bopa5WJQa3o2fgFYWYdkZI4aUGzvLtsuXWARBhzAV
H+BCjpjMWLG1pil4+igxJpOihxCACQWgj9zvCHAJrltAHdIMxK0VyI/Hlb26XDETSw8HluK1/SPK
NVA3fr2rRgzmUy9kydGiWKTU7rdgt1it4wTFjig7vnXOOpOS+ayAVOxiITWjRRyC2jLPJTWpQaH6
TBHn7J2joEvPkS3pzI+5/4wZ6bzTG9MoZgbLwIdzHOn2v8nFKm8vyVAaaGR1NTo+RW+qi2PjoWCj
wG4/uhFXFtZ31DWfZINFIl4bSA1SXRwq91Y17f3g97evUN8OJK+hIbTwt/dIDgN0deqM8zadjdz1
VEZCAW31q5F+vKKopC8k6oASygYyToB47NXdqIgW/KR0eMoK7eyUQlhpo03TJnPBkodLQmVOQQtp
iuh4vyvi4s8dbvZiVs+N9jWsBuVxGQ2dMrshV9/ht3Qr5KOJMPsWXqkgdmjtgoevn5d1jB5txFz9
Btvt30ahnAQoBp0v3MSNCmIDFahjCRXrLD3R36yNOPt82lVxK5LLFPyOWLE5qmYuNQg+Fa50phTa
nvHKL+huk6D8bartF6KwGgoEsPwg+tZyMwc4qNRE22uBmEckpXJH9vk25fhrN1oS75osZ/bBBx+m
Jimkfk0OSi3MhOxxicV/EEjY1ZVypqGi/D//C3uccGcYPuDgeQY5LikoTtPY+RJlTLaifT6V6CTM
7vHAQRGQvL9rzvG8eHfU39cYJmhxb3a4uI53fyLW7LDV7U8GEvSbk8SztlPVtj3crGZZGSCBEFM0
h4konEQlkTptRDLaSJeBBKjpMAdLzEIfd5EZOf0GXqt546Yj11qn1g6wXCkg1p50/mXUEIHYgVNT
82eb0UMPZDxwRMgPbd3UjgMxVuavMC5Xgj6VoRYyqBfa6YdWjj/cE/VMjvYv4QA0IcNiMfRuOZLT
glsWrAlOJ7Ozzk0kLNu8cjrtW23TuubCUSliniqhMm/P+oj6PK3meHbT44uw4He0mhjJI4gBvkuo
R1zsEXIXH5r9ZMACRxY0WSRbGxWLFu5wm7T/HH+ahU1Gf0co4EtF+oKx7X3atOLCehXto0zwQEre
dNDQnfclcurSSfdISQJxyPj//+QEnMTRrsuWtQgXXwdQHdze4nhqkpftZ1Ybb33+p4UoWWNmWJca
Jq/ONnMfjoXlBM772oZxTHl87nc6sq9yD4IxQMh0yzszl0bGNybkxAYCSmMMmBQafRQiVq2+xi5z
j5JCqNFP3ytbj6GCRTjeKNyvrK3xkSlPMHImmqsLGwpaBzLpVcO+STRz2AH1mJzntvMhwtD+Z5tQ
nrSgov+fld3DTBywrw2ZZ3ppzjSfD93sku433CrF1JLlMzpmQw6K6DOKAb9w9SLixI/RCL2SCVqU
C14c62OKIpIYP7b5qa/0MRwahtaPD/6+NwCxU14gujCED6pU+Ayxb7Lq5buWjTJ+g3MiYE2SAT8t
HvEmXX00eojzrbMF1FKcMoeCM4tf0dJoasNC0jEos/7XEq3UF2A3bg+bE+RaB5u6XXuvfh5Eqzi+
YXSuBr5MZ7iuo8hp8hCEo2LQBizjFJF8IAC+M5VgYY2GRLjw2PhKTclskHGH9jCfQLpBCDQ7Jagb
B29yZTX3UFYIgqWfqpzWze/KhTAmixg8ewCr5QBwFBOjEhVnEZ5ZQc/2C/RED1LXUZ2S0KUXHt3X
XADLEq7VloilphJGOslPeTv6/q4eWTxE2cnhjLyr5Z3rZaADh1DXkzGLwy4uwipCC0bY6gH2+wp8
dN/ufg20sVqhi4Zxt6MPwX52ziiFxs5ep8O8u2l3LFN7BSdimt8cQ9CKs+B70sNBhq2WWnQo/2eN
QWc4m1m29rqaPw9Q+s7zAXfaHj61KJhWKp8xE/i5Q91MP7G5ISlzJjnWgpZGxdvsG6Lwlh0hlsji
taNEgsOxrg0LoDypF+fDQM2gwvoqfvGAm+G5Co3mHz/SV+8uoKU8+vG2CDzlwZTnLnAX2CHLSvj5
B/SiqRd+AAEimF+8OvZ2wkmgyj5t35p+EL4A2tNSBpLYCm29zsoWtiPPWPbgGnCJeflhvPHVhD3X
gCXhcMRVnNa3X8kutZ7G8caH29ee9zMUh49dSQ3W6hSge2DQYVzhusP7ew9y47vjMojuLER2ftxW
kJ1LWMPtCgv8Ff3YgEy+fB5bVItXuA/vJVjzk2v4+3bvVbImNO/p+/eejXCcQQAFjndtoJ75sNzd
wgZP6u2GpWuPfLjo6bZ+8QJ57y8PfUanq53isqoHL5jhXSrrSItqHS81FKPHMe9PnviGBbtaGKjW
q/CREqDQgWqFCCtcKOebo0xSQDL27/Kqmr0ryQSOHBwXACpyL7UDu+v6ui+Ph9tZIwDlWnGzDarA
6AVHpF2fDaeqrv62K/US/aPY70sjby6mbqEvrnco6YOAzGCbsnXx9uWxtCsA/M5gDFX5Ir5ZhwFG
VypRuG0birlzo8czp2gJimtIg2wLmNgVBOn4N7ZSLGXmEH9IEYPBPWrSRAgmyCcOf0i515Ydivx3
F3t91JFgOq5tf0G10rEUbmwFIhLYa9BDC17xWOcdSjVsuTzZYWisFZ6KSA82fbffpAuhEidwgzmj
8RQW6SvVj7kGMSiRGHFXLUDeME4zqbc38qJTt2JvAIGU+dMPWasGARGlzvwRBu6O7cGDZHiL7OOz
fD0TSbdaqagRBLqP7uNdC6R+ACUtJlHf72+6y5Z9jeAu2QnQE0c0BTa71RzcmnNQ0f+uaHDySNWr
tnpu2/jt1ayTjcGdowIZrjBxWdtNi8njxU1ZkdJf6K9hV2JcsSJ6LPSIjzoT7vHV3Llqfs3azacL
mUD/eSkionq/xIFDzG8DudUCPzA7oqmvEMgEKJtZX4MXNKD0bSdOSIZiYIdx/6O+bxthIrKi4fK9
+28631twRCq0Ij/mS/+Zca55QZ1VXhA1MPK6sUlNws0CL5XNAO3Vtafo3VHTd4k4QP1P4xPsGS5a
Z+yyJPY6XSQlvKopzwG3tErbzoVYtnExTQJPbk0Ou+wbDTkXBZm9NEk8uQgHJECbL2ExRzz3YhZi
rdyKK0tCd91DcYWqiR6cjOz3ig38frLpKqc0QS5bFUGheNuQWQzIhwojebtIAD8hp2VDhNcoVc6+
/Tubds43rT1tjbFQAGv/HA2T1zBa6IFuyDCiX6WrDrx3zzYODTo9FWGkS9rqx+o8IRYqpzvso454
60UH4kA7VZAKBF0HT4vkvROnC7SWVZJlad0bcaCBaKN6DZLTIiAslvKDqISdEZFUmCQD2mm++ZGU
kVOojvmaers4Z8DzgkyRscYMPRb/Nb24vZlgetRW6wlbaFJwbLeF8O3fyftsp86gCfaKD+kP5Szc
OfIlDKy8GJs6BlqB6kIqN485IgXGnUo7zp3AlhQY02M/lD/kkCU1D7qauphnffYF8iBfJHY+EDDH
H85qphaHGq1uP/o34a8jjhVejyrF3NqF0HD3Qin9/j7G3zNTGjHaLMLxM4XbmjFjfa47xwks1XaQ
QddypULQoCqWAV8VXkQj8A+cMQc1+Zq8M9/haEHl3YOrAcTy/5dwTxTITr+e/dLVRcXiUEv3XiBg
PpmZ5XECzkxBuxeL/y2OBRWGZI0vSamHdDGeqo1/AzKbENPBLsxd81fdEbN6nq753vh+vHe/KGAR
wYSZoBi9I6c//ulNOdT/ronC+axrZK5oh+CtZtmbQ64WjskBA2XT7Bzkua1Lkj8Qif+eka5wLynk
Myq9+YfKyqv7YI6QxKaq3Gq8wCudnbWjK//LLlFbDeZIBIJ+VyuqEAoKUdPJa6+c4MWWhJkpJpPa
d8rMgg97n63kG82sdQv6zTIa43YcmlU0iC37iijFfv5lUdjWsgEd5NIMk/R/voivXT25/i01leAK
M3ZGoNc7dmY7b5CA1t7Y4cGRZPXry1Cy035B58BGWwh4w9dRPtYMG2iuDzIGvqpWNqhG1dvXbtRR
+kNGQRRBGNpPvO4Dt9f2PFuNT4DGV79UFUYseWVNg89gm6D5JGN7ll8DHrv00SrR2A+vJGha5uRi
kSwbnDpUwlC5qt9lIciZStnNAvgu1kXTGVKBZTEePvffDbPd/z0Gm6q5nvwqp9Ari4ds+GfIT97l
Txf100USW1AU5FO0mfZn6TG3/5PF6EsuhgkgfVmUzFIdb+P5aKMTJXqxcQ4xsMioJ5uALxMWErEf
VcSYE1etFq7tZNmVyCHhS2s2PLgHcE2EdVKAFoXK3rk6t/WpqlDmT7+6xnWnHsySgT+ccFfY5QA6
Gv41gFCL1ovmUyCbBb7YhkJ/ZgzslAfR67vHthcWPZ5KhVlifWpoSqzsARxUYxCLo3HFe7Ar85ty
cd4lFbi9xM9xqQViziC9DvQE1wnItA4uRCLXxS2D8LXqyynnBE3QH9gh7idhQNTYNaC0Aj/W5zEr
hkkeSR049sXWo/kZDCcNznVgEbBDu+Kcmaqv1RGItaVoXsUDztCuR0QllE68HQrS7Y1QNp2xodUm
xPwraiRjaoXS60P0BvoU9DvS/pIo9BgIEipHywJ/Xda8oYDuBCJi1wyGSvPHluCgK+o4LeWkxQCO
rLZpXInk+8PkRisrTV669iMa1CXNg40i3QTUTY9flEmxHcrnp1teh2Kwkp7hr1Uhin/EC0lCTxFN
Ep0lVdZmMDX/2UBhqIzHct76LEaZpNn+ezzj1L8UpWH+mlzGnNLwnVaUJ9+jxDfyBaQmQS8ggIiZ
WSRzoh9GSN5IdrvVL0M9p9Ywf/yVCG7pYkxfFYe4nUapByxZstuGuCF4P6VecxEzA01n2pFhlctg
mQlWjRKfwVdm2Eq0oUQ0H1OAe26QS1cMeshNtsU8vMMJxe7hW3H7T3qsCS5U7+Jr1AIMoGsTlAg3
Gnzoex7Zz9tURgZqnVb95Hft0x05XOniaQLAZceck4+Af7j/qKON8GkkEwZsbdZu/QT0RglhGkJi
HMCH6+U00RdxrCmYG8rwKI/UCY38/6IdDkra2OnNALEr81jh6QZZHLN7RIeGpUj+zC+XpPcoFCFD
LZSsEXnKtSczv/O8nKEcGv6W3gRFqrmdl7oxkJjXHaYHYMb1DoGrgfpJy66g2vF72yIWbc7Il+Uo
XsrFvsTzt9L6uNxKDnmXjHfM16b1VS9aVzrcvSTM78bQnntaCJiO8QB6b8WoYCCyazLObkxR+pf9
zW1TFZxPjiNLVSlW7mcAUsyhMTvv7KvwlG/bjRBsESJXREZ8a6297/NJU+PBoaoIY1howQD0WBng
83yc0AU0pQviMZbQ7lldu73dKHtr5/zcptJUkkDZ5wvyifJ+Jd4vhEJS0kyuJr5PqFlgQXDLqlxW
C0JybskIJcZ9OA/C6Mykqp4ohDP2UxUAVb1wVXrZRVvBff3cvJMX/iqVXacq0WOiB/1OGHqoI68s
64wNHgz+UfK6QOBRTE3coL++8vAPINaA1vW3dtIcZy+8EXEckVSd2JjxxeY4MdpXfVgDzOHyWsgp
jCzqgRtXf1Zzt86ej6KwYtCGHnWH8U/Kqq+nYv+ecbHW2UJ6rs7wOtd4NwkAXlCbW1tOASA+NtmN
NWoQuwfgUjQIR0/hNV0s0uz+KNrD6GzIX1TmtI5UHrlzsbqiXzX+TAsskkVASZ9eKFxSfhnQq3FD
KCXxqAP8vPGr3maqjtNX/6CiL55JJBzF4UQPzDqyO6d47hzrdon2dgDoNZU88ow/jtAwU0vvoimS
pMuwBieMnvegu9OTkS83JhPmrTlPI0kH71sg5f+0pxB8v0xDDqWEZujufoRlo3UZJG80ihFDaOJH
99PY8Hz0AXilJK2aiVqF2OdleeplUmWeOiJhoqyTAbqlAj81ERhFvE75k5AalZSHpoEpSfz6D4yz
OgyfpZdSkySVFa/XEhHTx1WNLChTf69O4Mbu4GJUCXl7+9hxW9CmwzAELVAiayW7HOy3d5tsMtvi
9vL6YqYA+bHlqzvyhEW7uzAyJHS5jzYCUhkPoJO72TGrhkt6fY3bFWtbKP7ltc+hExvey9CPGL1Z
xFQRaXAa20FiB7eq1xsD0q0RqtJHcwFWzI6SDaEWjGQjIPMerllqPXk9mj4TYR/G6lXOlXTQ8Cos
zsoo8JmtVPcwnnSwbOifYT025weVvxeXmLPHIlJnziiBQgmMG0gD6vGadVyDcrSb7Fm6GNRmrA1Y
p0aaTRgzWTPc82JfC9BXgHO5bKA3CrDfQt2I+rhi60RD/PnzWGClfsvdrJLmwLYZHmGLG8LfRCKl
5U2BdaURfePJvPxQWTy+HpuYXGPLig8uVRvrBx+FFowTfxjG/NlWpzE0uj7ipErcykhNJbW9tXAf
RN9wQgqqAL+BIQWrNRMpmSwX6k6GcrF017DgOatO26B+24yZudg5LRxCgWQVI9y7c8R7Gf1mDZLI
xrgPB7sCVsuqjCRh949MdIKTQl6sYZu083tboYjOcfRgPNZwcBE7mmy346Yvd6Zljzaf7b38FCYS
noBuaUP66wAze06OjMPkCa7oIIHK6OC/aOsOaH+u7uMVQUBnqTv7vBhr81/SdyNEtJi/YJxqRy2L
LBQkGPEVOmDCuIAzuuH+AtUbEiTbQEWd+cntL6O7KVcF5JlxMr3F97rNHYbBiMg11tZGgQG/de71
ahe/Adr5mg7pQVbw2VngPin43OgOZiUG8dVFiANI1YNwi6sMQV4qIgQ8wP43NzhriMP8r3BpU+QX
YuVTm9mYfsL+/jkFUu3Q0FR+BfR2nIdlNXl7bwBrKoHqsdXj7DoCqnEk6XTMDDvbSoDBoN1pguHc
oBr2Fps5qJ9Jav0AnBswFKBjVXqKvQpuQAq/KCxuXt8Mqvu2ixqfaKzsyASUqnCp5sDTowZwUMkY
KQXdkLUuk6c3cw7yhsOuDHsA/C4U7zKTF7aRyWkgbc2lrMhxK8OH28uVa+JmRk2gTNsIAZTziBcM
IwncWxtwlajUJZ1C6c5RILb/tvdRxrZMtVym9+rsD8P36pg4jW15uNVgxFmfdbypQLiZUCGZweq0
WyMI3MdbeRpSu+AEbEwUx76FslsFxl/5t4Cr35kxd1gLoEdvgReyaVaSJuBRprKbSgep9QtxnDB8
OS5NrQ5If+EWxaTimnJo578+0moLG/1stPsio3dax00qO54Dcp4/7ebdv3PAi7Q5EkAlkTaC0Jxf
iVuG9uNuxRlsVSBe3L77Iyt4uDNO76xCllnQSRr2X6kzrk0SKRM2mZiiiBHwfFcTvN49f5dbV5q8
23Qfm9olqySJK1TdJ0i/28FfgYCknaXP54LtxbnbS3rEyRS7yUJKLl9T3SlxU75ss9BGxAdwbDeh
XFXLeKYU1IKgGvftXAK49IBX1+E5RKiuGsnofdW7oJdKaR/wayRyjRimBSEproFLyVeIO06z+3ZF
oWEt1pt9QrEzXB19la2oSeOf3Q+O4vpKLF+7qKSrUPDuYOfbAJ6wpDpI/Glu3XQXsAx6J0fzgYe6
KtfwJ54FlDVL6vJRyMQo00WSEqC91/NOnynMCFhwZ+i4oK1J4Jg85IIiwYMRhTuJU1jWOEQSX17V
pNadnackzadFDP5XBvg+Mb3sI1KajWTiW3qVHJoyYSKk3IRL0gphejwepZVEeNKbDSXATNifrFta
EL99yGY6Hv7vLAM/8juw/WFeoCrPBzWVXaxLTq60ZUA9/6ieqnGGQMsE7eraXQ/C+ZK29GXups88
sbJjVUj2z+RydFnT+4YsD9TvBPgWbtHNdwSIQXt7Jt1FNzOQ02JPDdHJ+P4/Otofvh0lCBEL0HKL
6U28NussXzxJKRephS5vZK9URpWgnOvR3RrGBai1sd5JswxsEgc5yIxYJLoCwKZ2X3zfAColI0V6
56LfM8WDwaTHDxXOnsu5I9mD+W2AkMDUqIXaZffPmceawEbhu3TVF+P7uIrcTuibbmFJnKEmlu5j
InUJ/4FjVE/fXxHuL0mliSIu77FIhNzhtk7aDKEAFlJh2t9ewxdtUeHCLxfVocAkckNnYrCcYTHD
RbSy4yHFnyJySc1k/NWqce5RACkeVBZnjn2JKbq2CNlZYvYqbSAx/JtlK4SUhjKeuZYvNS2XqtCi
Ub41QKKKhWRVUy3qEX7vOF1gp8VgB1EGvRKIdQ4A76Rz9E1gYvOwt9WZFcnlks/99PplwhZZSdAB
DV+jPz8Wj2dyTQFZ/lIexqgSsmWi80icDFFPgIqXQqVAIFueUYY+YGgdEP72GBYcabuboLZYtYNi
1ZGTpGxkkIplYICSa4i6P7pRw0Q76YGwXMWyI1AUd1ElT5TDFjpTI0UHnDOwE/cCjxyZ91V/PK58
uRNNw5aeh75UNaze8bNcpH4wrHBYx1RdLrLaafa1nUpUD5l500QHt/lAWCvZzg0uJABBMr4cizL0
vPavVUSJIbM4iLhhk/wYPDonUKtKJqXeRyy6WkEPd3Vley7jOvUXkdiith61hPCOCon4c4e8rpnc
+1v5W+0VuuIzQUaHtIL4KlnsWrzpzzQFgYbjXTVM80IQiFR+sjzHdEKIQCSVOI8P+aL8lDpKZWDQ
5fm6qF0ihz8EB5Afq6EaactAmMwBY+G0L9lPby1BPAawW5FClScrAClzi0vgpTXggptApANp1MrY
KirjhzRsTbp7Z8bpF2Kl5tOzCLhRanVsdtrV37oZejKnaIq/4WLZ2kUggR4RWNM65GiSAigRvbtD
fhKehZ36bjS5F/7UCTYRbYcQzuedu2xVGuKwlBOqNEvrlS52fPgxurShFXaiOvI9E1Lv9NdX4+ZX
WaysY1fzcM28t4DMsAaw/P1PqE9zqGLGoAPtkcSqGiBsPPpf5UVcg9e/6Pvr2Xhne+gCJddPiBLe
ZYxI1L7EJllK4s83lYPoWv5UO4Y7JLbw1ZI7jIdqT28555F3kDPT2UvUns2TSK6wxK0z6ryWpUPB
6NSN1KotWS/FW8MOMSLa+yKVTgwGtEG6ZgwbT1h6wW0Hm3FSyNSaD15ExdzwDKCjMNT2/ZJZbo6e
2PScDjhNXpEgpcQAW5I6UIztIf5xN0iCAUxSFqn6Q8GNuPz82WEkvdZc+sdXg+LEFflODB0eMYwI
vpWmisfDKBPTAk2YqkQGhiNRT/q26Dnj132AuLY56KVxjEvmAhNUe0GbEtst1pq61BVorZjKN1cl
iaaZhDVAKCv+835REf66bxi8O5oHhbXENCGdE3jemsdoZD7Ij/JVlgQ4bsMyXWw24IEuTzLHEriv
0CMhazXMlrJcI/G4ZoTrX2ysMezVyPhUR4dWOT5m2wPRZbbMJk1Z49S87txjGlpQw18m+IJHToRb
bKs1Lo2N0eazkkmCHS2p/HBxYIPgtih+ulHjKnvsUPORXUwcSS8hDHDCy4NvY2GqMzDxDw1wAWP0
jnvL21vw0Bl35HCon2yzIeS6FPd/4WG9Nibj9Ei6nkTYr7/DNFwak7moA2FjxXUa6+TVC0yIfnPN
+h00awQibkiLcRUwVndUzpvTSmTX+advy/ykZvTX7wrcATGB9DBeHNA6AUGKjxSzn6g2GF3cHIFu
ThoHqJby1OHLyXdepvXy4OcQouxrLQcfA+XC5hSzpoO/xfVXQ9lBdAXHu0j/mUP6kldMOc59cZ+q
x/rEtnRG84q0d5s16TJ/qHFzK1jdxpxFS2+UW2Ok8z9vWOr7PaOkL8dGmOGMT34Qtjmq/lmQ0pnH
1SrxPROt06xVw5Y6bCwevTjEJaNdwA02P07noQPjCZfv62MdGvSINSP+xM/fZNorNC+PIrwte9lL
IknwpVkdBSjiPWUXhderu3bPNIyH7cIMvu1jUXT6xLIzk/h1voZvnyiH3CfOeNFTMcEJ0hguk63I
RP5+0EBQ2QiavX9OjmIhbtySpfMsx0RxaEN5+BoX8UPbL9ZrdukzdeWfr3XHMzVwd2a+dl3xk0Au
ezPDHTR7guHq3KbNjRItX+FZuW/NMRvNFflPXijaxmzRfxapZYgAhEMBdJ6hgHTNKQtiYmvvzNLY
0IKZy+glx+tjT4ULIU4WkSnhoowSiA4Xmfjiq+pHamZAQ9XCHyoIs6uKxTO9DIqvEyOKnhbZpK0Z
XXHs46lW2x4PhNzVgQ/n2EqtxNqk83q2ymyWMWo1vMFLY6tcMXMLm9RJP9LML8ghrHUiKuWm/FrP
EstKG0d28rk5ye+EHUtIIKQX2uV0YJ/Ok8VdnMtbhOUqp+QUMMbhtWI+Vs7ATZ+BftHix9tcU9GX
EjepOV/ZfKV3x+HHjhVo+h1J976r6dHP90zsAdbyP3QIHlZSEOPRj/sSJ6qEigm+5a9W5Qp+18wp
wM1tRdic4YwFPJXr14E93SpwFl3MNMpPgA06v3Vf/O7bPyJkEjZrRlnx727jOaSKLno0SwsFeJUE
ugUDClbb59TAAkEZfSeiS4ERs39Dx8ZiM73oLWZY6aEYaC9Iomp0PID+J7Cv2QggTsDOBqCxSpZ+
5J9UPg/C03xf5/GcMaAYpP1ZzGAMEEWiOdo/i9o6rfE6x4wVh7VugabRFHqVdnY2lcWDfz9QE1Rq
ZO/htzPPBdZQQ50+elF8tY+940Hhyp1pmAcoyNWKVb+lOiberNXbDCLEnL5BzzJDaoabpDjD4PlU
Q/J/jibiF7hRB7YYPhb6Me3VpV/3X63gs0D4k5FmHptP8SYhdnAle7lIUzpI+OCZoMs/xaTnVIUv
AAEOOxQWGzYOic3zwz/FM8MC8g8WEBirWmmtBrPJqsN1uslbxcPgTSJ0Y2PdrbxUYOt5bko/XjHU
IqoQH95XVRNqrulKhtbbZpBde4sFwnSSyneK0DwUX/gXMGx25Z9dhH+mhvZUyzMvxMmPG6+H7Zyq
RgjXE+7ECzvR8lW+GCgM/uBgKzAxCx1df55X+9K9cNik0Eu+0MtWFmjsSMJPmJpW5vc4WyjhwmVp
8wXuVd4za10jaPfNyiB384smUIV3m+o4DB9TIoey3KmuSblzPqkxxf3KO7QmxrM6u7ZfDbhWAmUp
KTTIk78vrfTfV0Omn2UemJBZWa88qr7bl10GffWDguMee+pCkP30DK0x2uULj6xloQ8ABoaTo4z+
C6PzwZ1CIKtj2XI6/JCNycDej6JpGvyhIp7QbtfEPgxMbcyoqlH0Q6Te/bXu7GRocFOzZTgFLOAA
s+X/tzEmiWLTKZEvbLmJdsK9FnhzfABYJnC71Q3AYbr6Uj7YvFMVdX0lZ5oMfSqUmEtXUovwtMn9
0q6Oy127lBSwNpTUJGwitKIbUl1jY6aP3o7NtIwJy3md6yuCMKZyIWxUxcNLXF+EoyUxOTFU0A+B
IefIeQXRKBVahMBjKhcxbRjJK/E7G3cq0kv9vhN4lB67c4PBjVtTwMp7Cf7CO0XC1ciHiME60Upe
cNLK6w+Y7lNAsP05cX+NaWqjZV3AgqfNH5ny8lLH/9PqNV8A4xR75KRdvbyymskkehVhkpXzG79+
PdxAoH+UQC+eR/fxRJarNRC+JCwYk9lPHiRDmMASbCW8TzhZDsHXKuBPlnGWH09dvPKIts7+1Jnm
/gOWFkBe09WMfn4fEQMWrtaVst0ZMZBbfJG4ns/YZrr+LR2cQCGrXk66daDJLqEONHR6rd7GBeuy
xI4A9UwZ4lPDDX6Z/7DUpDDu2UmvnIqZ2ecUG6l95Dmk90xqNNe04VUP3D+RZMZJpgXBkcyg0Yg2
EGkTHdRhq67ihO86P/sYaRll9G6J8IQdEzoQTfUoHxsEyeg0dJBhxIZyArpCmEwQQ6S8z7+0ov1N
7dQ4uWaThrC8BU8T/2ybpWG/QKbtyjJv36NSlQBUDVhGyeI7RcOoe4OU322hPFoe+9apzcplbvcw
0NV5IDthNLFHrnCvH0aiho1vUZK6I0+42kWMdUnb8RKQ5RTwpQSxInDIVzd+z9HZErepvxl4zEo+
H0QWltoM1Z8RSYbUlt4NhURPCmnacda7nOXWfX6vwS47toe0pjMNqpRFcEoTu1x3MR6gjFQ2M2Ey
skfk+4mLvrOSnmwDB4fB23VQ6cMxPDHLtkfOWCDVHeyEwr/MsujrzDrL92HFU774JNzkKQrmVJ/u
9DmGaVjzTjUHWL5U728pXf5qHGc23eU33OL+qvQvc8VaaMuO6Jan+gJqLgPgtPWeOYeJqwe5JS0I
O9bZjpK4iMtpL0+xQ5MSXa49N3DaPjhsbxJEAx6p6BEHzshykRIUuGXfm6qfbRj+aeEHKfO4S0b7
RO2sRaFf2xJ7p0bING9dEKNlkKZSFjynOxjfAow1BE6S9wLGzZPn9kJXtW3AX3K8EyDLmxccWnSU
CsR4v/0U07lx/qUUz4Q7yHYhInXz1v4AI0wPzyZfiUaHKl99vzaWPqSMJO6FZ8oq7hr5CTGvGf0d
gr94BzPkWv3am4TqLW/8LITSQJcUMlKAe4NN1NGov3jb2m0ufw8hHgQ8xcW4nW6ewX00M9I0AS0s
AHXKm5gQssvQ5n2dUun1pmilkdyi6MfM8PmrlxLI9d78NvJ+wz8JeEXdyKic023dk+L0+ncXTNPf
h7Oxc1qe7qakD0feK/UUbeQD0n6XS7vA+6a7f7A/5hQL0QAYx7LrhDfEBbMO4ALfkMUB/ReKCgl+
OlAuC6upOFUsu4eKht3fUsp88dmQrNC2SqAFz28qJa4SfWUb8HSZ6psVDAo9wA+MZdhNwdE4bXq1
zNxOSFWEWQFlNbB1SrzXK8F+sImHUv/Qv9DqYEctqa3o+csfG8Qe1wWl5pVgDCCZrIqitFmmLkOf
CKxxOwp/83l8fvqR3DRMvrG2ZZzGkorI/ha547vb4ecn3yMB4SHvIuOgRm42aY4pAZKzDMN6rI1K
DvbQKKhIMGABSlcLLRplAN/5IeVWAGovGgL08SQB6DvsJUj2E+qotj5IEeF/2ol2OoJrPAKxOjiz
wdese6SWCVEswZ7ZkqdgVG1qsvX3z8abGq7vu9f/ECmIANFQdrWyv6j2Ic6tCXOIz9S9FlXHkhYO
9Qqj8IObc52HaAcIExTSZQVQDWcu+iEuXHu4IzQ9R3ARONpm3LBTmLWrqexPpNzzoXjUiQCBt/Pu
RhFz4nyXp6S4IzUJ7Vs3Y0dUB/k9odNEtKaVozvW1YVg63YkgFoz5X20vL9TDuroSjAQtPSot4Vy
NC7pkTheB22hqv7B8DWN3IdE1DlyNoQ/hXvR4t5syjVr2yjHj6fmJdTh4aASMOPwSE1h1e4Qzj1/
aPX3SwR+VCykZKBn1LgQmLC6kLjv7jKXuTmV9XUsjXbw/bLlDHLYLUrlMIaIHhX2dno2KlYIIXTZ
r/sFJBhrP7gUubBHj14B1zknp8luaW/2/CEty8c4Q081PO0qqLjq2c1vWjRTcT6GSej4tcYZCV8q
R8kLdEZykYAhOLtTLAmr9EHcpi9mnysxs7rUWLiCqIPrDnHi5jjobMSIGur4LfLLdXNeX5R08Zlp
prjY1QhUoVNLIn5waVthfqtsUkZKkeYJGHTspcOMVPkqBcJFdLCeOvB8+VczUGNQY7TeJGWPxSzA
EhaHanvoRoSuwn4c2EKImKCAAyKI0vqt7GasTyPT4CFYehwPwO2Tc1BixSPb6BfbD80+ie1WQd8S
zy8G1S4gSctWatSpMGV1W2fmbOzTugCXFPp1IWT4bfYSPu0YvTpZ59V+kZVGHpkX6OIr1E17pM3a
GPaN6SGnRGsA3lCNxggtc6tRVo4vat1jmOiScJ1Lid1AgRfZTxwuj0s0EbDLgX6DG/1QCwThCcvw
4dNWGzZ+CM6/QRX7fUFfsW7okS2F+hp9r5oCRNTUGrUfBDD9O5JKTEDiWudnnof6Sta9UhTEnF8X
1Y/U+iVgIpiJLHs9gCLGrdPfAmFEhsIbDxxKbf+PiI7PFQo8F2mClYrDxND8ZPH0Qi8M0C/435hN
7zEaBrwlYBoKH9Hc2Hih9tnBpa0NeJviQit+IXijoGGvgLscqlWstyqHY7dx2wZkR/hz25yUHhhC
6pHe74HYgRLgYLqPNnUtwfh01yeW99D5BeNcNQLLcGhW6s7MnVQXHl2wdZ3miAEsD/7gbrSll/Md
upKs4S5TBMoGVgTNjRbHO0IiQkkRfGCfNcD7/7wtYJJAOjfeFOLlndZLE3INHw27XF+7m4b4Xqez
PIu4jGLReZ9t4LpUgpattDH3ncjLigtMVqPRFWhxej10l5WQ5V2tcSN7KbXw3HL+0RODGiodqYAi
kdlYyGYIwY5FVcGivsUb6ib5QunrkP5L6tw0CWGB6eluTgTDkUcnpvZ6JTNG3E1KjgieK6cKz0/5
YHjkuqRMCLRhmvcL2tY8W3Zc6sXjhF54+++B/UXlkHUQs6cKk2MQv2XYlo9xR9pQl648VGRGLLck
BebzHRFAVzTXKQ2mBUtQ/LMktNukMw+X0k/uVZkZHd0H0Yz5qkIEsg7kh0RzyhPm/OkALUh4Pp99
FemBSL7xuZgSVqNP/aAFN9ygC6zJmmXIZWGA2ydnqtXdsh60h4eaNHigQgzW7IrKb/xdLprcXJ0l
QTVGuXW4+xG+Ma2UYDUrFWAUDS5+/02MQJXM5kguAx5vfiIj2esuTEm+HhrRr/hVoeCl6WjasLx8
Lqvh5YRfKm3Yp9uH/a9HWL/atlHXsA0vn5mfw8aVJPCwoBIk+80Geg7vZRyJO30yU8kojH+MM29L
OR8o3BZcOXmMHoh99wYruo429+m7Dqoi+SI8meMoySznknLBMJtDWeIk5YJQbPVwUoE9kgkirf30
2Jh7lT2xM6LMq0rKJ6mM9KsHiIxgUbvI7ufQsj0NeYBz5VXnqO7hsBciXh1d+JRk8Yd1brAicTGV
88kYrHOQpeirCIvn2pHql1HElMgCn60uRV4VWxu8P1yLVOdaEoFMjtsgnA9rKjnQ1lBTCT57HwXH
lq8DT0Ybop17+j3qMUnnJ94uyxXZ7FCj5zIwDW2Ih3zkib/4H5NU68fa9jHxKztktu27NuXUCqGk
NoukPh7GxuoCkJkRKbh2W/bb7VKRqbVO7+6OxnYg0peqneOFQcLFFoAhEfYQUD1IAPB7+1pA/weT
G++OygE+Ljk5mshYuX2egvgW2aCjphncf/a1mRO7Jc9gadZZ8D7wOWYZ8XoDLVFQIMn7wN+oEK1h
7ueI96NdcKOwZ39tx9A1sdduNqhPVqcFIjfDQC+iE4cb105my3LYmZeJ468JS7eckngB0gGDxTlG
G3Ua593sRCvO5AlQ7oiUlk3N5JHAA6xH+ppSnIjh9IyDIACjHGM5BbQDPNm4IAK+AECynl+UDwX4
8FZq0iDfZcA2dHBVoS/WxTcmDgdRGiCPfmMlfe4Vcl8jvVpRvC9olkNiW56wXFy4c7SQ9q8tKWCb
mfLRX7n9qg+IOTICN04DPYGASP5awBSSHRism0MxrhpO1f7bQkvDd838v38nPn87RRHqvHUSc6Sa
1ZE9v8W1B2LoTzcUnfnOCmPVP/9Bmrd27iAAyHZxkiqmCWNmLtFr1GeULMl+jdHJWLlJ1Ewen2gC
UmwJ3KRW8gBMw6eusIzSQ5a+Qd83NpZt9LoRnNNQS1CAT6fd3SSCDEL/CHvOzmhJQ+CNzJZWIy1o
sDuC7jd1bchVWALd6eU4PVBW76Ld3fWpsxqi9iwno08zD9d6O8cTdT/TaD+SAOOFRlYv/PH3PlHG
fFBHDGndgZsijSX9FKZPxrvfgHMrKVfHGEFFQ9w2snOecMWvyRlIg9CHAVjVP9zhaJjYTBNh+0zQ
OtEcHQq9p6QtuZey0Il6319a3oimyxj+Q6bQY1mBJMu9zgDx5PHbyIgPUEw01DYYFRR3jhCnOjWP
4pIxDvN/AirPK5mJy7LJvKCsUC0IWqfc2GodwEksaZ/TtG885aUqF+mjCksRgw5/XMYl2JVZXhoa
dVDwNmbcQ7B/XIcga5mg17ABHg876Czttw5/rrrE2JF/hwZMlSIoNfx9YXkiD+5Z+joBLTJQ6Dy9
yJ1pXgtSSIenRfcoK3SYJ3PRJnCkTkb/cD/yyTu8oQjm9mf32owONy4YQHHs4kmP/F0RywpCjXTb
I5A/SRETR6flxwjflNhh9M9M0oQATNab51yq+0ng12e+BH48ct8ViPCJkVBOKHsYmGccGjOmMX1a
oFfTACAESy8XgPSIUEy6UYXZiqx5P0MS7PXTXlzp0bMoaIW/nQGVDHwRGV8tefAzEA7enS0SOLLq
jKj0AVgLiiNLhFZahnptDsWQ4y3S9MH5ka6Wbjjq0MkKa8OBnCwXoGQCA5aAriSVI9IGQzHXNFKU
nq0M7EP7IacPrWHhEgzjSbYMOtMpMZZH5s0BCCtNukFSGEgWXQBmV1iqb+ZVsctEk+bYBNzZO9mK
LrkowoU8mMbuszGfX9M8r56YZpzPplfjQMqgwYLyGYFY4HXoWK5pwSDyAjAWFrhIlvw7r0MJoklQ
RUAVjz2zoEL3MsDZ7KCtrNney6+u9GQs4MwHXgZ3mEdwC2xUEmyH5PxIbMyUGf6qg7VaIC3wsdvc
xbyo3tv9gWNiZhtDYDUk8NeQ20bknS2oXP/H+/3ujAv+IB7yvNLktVNJCWV/8u+JQtClgiKRk6Ey
aJ0t0BdQuOOl0TNqYzGg0iTsB74a4KHcTzxF01630XFp++5LxXTFecQarI8ymnF810ksqWrMwKrD
S87uPQatgTRnAlr4zJ2NOfv4hzro/h4idRT1pB2xhUnb5NvkrJLOvCA20qKAzAUyCprWZ6TOj4kj
nu4T5QmlCxTltLyoLc9XZa68isIYj8Bhw2La2csRpFGHLOyu9fahgXH7rja5HA4rsthwbFitwsPt
OlLcupBoWIQmSQr9V5Jp2YvjmPUwDNY2qiCF0hsbqG77Br1gGz3ipx94lSx5xxoenW7Uhiy2L89J
LCDWAer/hiBJawksmJaDQMOfJGgnSmrJr5xzYPc+3GRzeIL1iDpfxEyBBCU3UdJcXj6ZKiLbM2Yl
5IPlTHMYCtMKqZ8XT3H3xz5LENeBRyd6j1KVnDHmPcpz0dgx6PoGv+nYRvZ5yUciFkfDFA8UBxvN
WTtNOoRjoVI5x6kUaMs7HZcU+yqu3t5/w0UhIjbhU9e7ouCN8mxNnZ7NEw6a6gibVGI8YcAY6nIP
BBFsq58UbPBw2MEXVXpJkPHvjfo4EjI9rMqlPI+KpGfjS/aEWlTHUhgRfy6p7NwgyPovcfhmgtsI
iPRVoSrQQX+qnaXiKMipJiu6f/t+SJJ3JV4O254DFDnIukEZdv0m7DdvTN1KQeOGQKc50RHozcG3
xYFrXB9ydJv+9e1N/yO70pz3LXxHN7mIQvR5UgVE1cyBG2uxhPc49udjxjXCaAi4HzF4fnoPNIao
4TePyDpElFOvFTV0aEcXw4O8eq4F5RpWplBONHN7X3Gfce9vqMQUiZNTsWOCb8HhFL4yNSRx8mq4
7K18S+BE1NhSxOCj2AFpGANVD5TZh5GO69kRtOVfa1j+hs/kKZWnDtV77ZNCXw6rzM0K22yQ3HLP
OF+eLCD2L+vSlndXAKgg6SJhWVwk4E849LX3HxYTQpdFlRIJp1SsEFN4FAwT005ZsQlo4zqyii/5
uhAoEpKsgZ2Wp9zSyor9kjVDqCNupWy/o/E6X3vofmAuZMcodxqtEYPjC+GeltSTpn/edjYY+LLF
so3aIMDwkf1PD0DXSGsoNmMgdiMhS4uiRy2MqcFLcrYSiwcJLzqg1poGPgBUsi6RSIWYHqJtRp8X
QJ/hUaLa0c0lsTfyvbTDX5BJP4XGG6/YjpA3PYPBvqgOprgNMUkCUt+VTKqG/ys4ktO8N/WLRCBC
l1et+rI6LKsYzivO+wiyHVpzW59tYb1fcP5XvbIDrtXXl2CWgYCe4/V8k8bUhmaegyhFooKI/E6h
fAvmaWvcKZtyQMXbPy+T5zRtFPqa8wV7P+O2Dm2+iOQ33sAvlt3SjJGQLEnP2bTQFpQIZeE+JNlp
mshxbIgDFGec5xc+gpQRAf1BMfeD9/hTKnnGUDJ00B2zzfoSE1tUUzcju1KbKiER2E4N/iqzFZlL
zuCtKLBjjg8Q8jhhgqq/dc7dE3uJjdWkkKI+t6Kda57czbzJL3XqDK93Mnk/cSNZeyVo2umc7esF
h+jyuM+Lbk1F0JUTo6DBjchSz8sOm1serts0pifNAea6WC/zDXsQpLtE0V7ESm/swj7Bn09SpIK4
Pm8/FBge+cs3liDxFDVSu3wu/UdeGF9dW3U+RbIX9iMoSudkBiXObpF1FrSZbZn3zZPvWtWUbzKv
bX/NmVBq0l8me9y5zBZs7XAanq/gpTM9cUPhHHKdJoZjWT/0NPaCgc10lW5C2VtDr0ONrtbpQnoF
enrqx7lMj9B17vbX8dgUASJvK8TrdWc3vPu8sEVrRvLorws59ByyQuhWAz3NxMDbKRT1ua9kVYR5
l4W1noZD42D//lJINFc7vtBNhXVPxfTgE2c06mSkMlxPibuIGKSor276N7fhOviMfrpf6Mxr7Y6G
8aFrA7U26G244nO9cKt/Nme3jBaKBIfOop2RGJTWEHNj/WI8266J+EjtKk2+aVeGL4ZJTZqNKZ0q
IgoMtgj6oYvx8VyHP6yFfZzN2MrYUlN5urT7FIvgkdjdkrE3jdqaRhkyWyrnHXW+Z3nbvW+dmRu9
N6Ke02i27N6nWv0lwQUMFWc+KjgYchFJ2Mne3MFR7GmZuz7K7gBVhhISZpURfgZRgBthHDiLPt/b
wtuD5rkG3TfEDrr3yAEjCViZg+l22J4MYaeEkd09nqmsC8K4dSxq3W45Ho5pp0UgTfRorByNZ89k
p8RcDLX4/BqB/qvBNC7yJcIeuGhCX6g+soSpyDrdOUNvoQYUlJpEt+0SBFqxqp5FnAM2KByRxP2A
xU1hP5wxqApzt+iyf/bdEuPh9oYHSi6+uUMiuuYt+ohOKTHyjpE39guiFqQmLffJ8W8snQ1RFurv
EUkLPTqsw8HI7VLzjbvPxIDSIpSpys5nfxb5RN1RIW8qNn4WK9aghCS+tS8HiLCu5K/krVnUrKFM
KOFvNG6JKKO9A40TYKqQrpOD34RrkJIXfZP9+5N98xKEph35QAguQGPV2tFTW+iRgLPEn1W4WPdu
Xid7jfTHmoVSA9+AgyEOfvrUC0dr8gDLEo+Gi/+749BD5DCAc33vP78gl8T33Kt1cOdrXlhcHL9p
YFPyH/qmjbeCmlOCZ+p3IS3OsNgua+qD3+ccTMCLwP08T5V9oQMhoPajl8gSNyHujBGNaYVQZMbp
AhjdvYWsh/dVJJk+xLEU99vvL0s1hEWYvBL0WdMtDxYarDGlARi46V5e8rgbhe0zmVblBfWHTQ+i
tlOYdxwCtSdnsJlouitOTd7OnfYnqSJxYZMrFhJ2n2XH6bHhqlPw+XdwuNtvhY8GPdSCoRxETol0
ODr01PKHIPWKhesnGInbUi//PnEmfFmqhuD1cF/uBxxoxBVPiuVuHTXfKciQSuTF9aWgpTqkF392
9EsvSOqDXID45P0DynPMGZgPMGRhIWSJTT5Xp5BfV3cY8XtAu8sjmVJkHXsX1rcB5KOmodLnlTSM
Pr4vA8ZDnxAX/hE53ucVSp7OSwSxkANxRFqTn5XPSE/XzTtwJfIObFZge15aQOdcPgzM3hgBfpck
BKxmVgwKP0cpo4s3t0klNH4yOsHEgC8sHVMzniK/ZpMlVgSIwJb2sMFUpHroDNaX3lF2TspYA7j7
/Oaud6hoIwRKVG9clAJypDHbPIysfKGO7C8COetUWPU/gKUsDJNVeUX3sY0m7U/Tdu2ALKoug+3c
gFrReFn9WOsVtC5CuG6d+FegohXhizEllI9j+HxlDUbG48zu/DzkZdYxgasiEs2TCtJHOw2uQdvH
JoKMipFN9ViiBdECR2n7bBY0QV51ZLo//TdKBPMX9FTCojz2RZwLPQHGSEIgkqu93TA3a423PtAo
pPKIN41NFEJkeJUgNqshj2vkDaeLV88iIRLjy1YZ5IeqEVU7fpDsBX8FU+UcjNOe5NFoYpNshRJP
69XniAWvoZZREnk85K6G4Cu+2LldisH8joFeBDLk9RW8fBHSgksjrrkIC1YU9aYNgX3kzJlAGAzC
Njw8UWS5cECPzVrhMM0NdkMADv6nd/7AmbjWpplOxRHLvgBnAumuOrND46N+fJfDYT03FZePwmM1
3sbVxkmp3TtcFr5/CpWXuwqkicxdNtbEZQC3el4UhKqHJOIAWb2/HYY9WUkEfWmMSHrf+JES7lJa
eEAq633byh4kmbaA5KG/NoQ+fQ/Wq2KuUlgOkl4e1AEcJq1HSgVOqiBdo/KfJvkDiIHP06XPih0j
NObjAiZFMdorXI/Uw45QK8pUoiGdcNcyvNjdfZYMY8npCXObk7BiRrYlIHXQcTd+0ZBmuyOBcGXT
sVVJlXydvb5wk+nFrbejHTJRD1Pq3YuG9mCSWuFuNyEvXRYUYdK8j4c5G/SVLmzLxpxdDNfb9dJU
Z4WzRU1ZlaZdHXQJ9MWjCYRq/+AlYTbq6hjG3dJ6WJM8Ur6yXJv6NYJz657IAPdbBJUgDsZDOIsw
dMaw0zGv/cn343D+KIwtMnjiO9hnY6/sd6AZGUBY/lbH88tm9A9KeVtO912mMHUJHVSMKQqp51Cg
vAeuz3U9bpiLyBdnL51JjBg8zf2vTROKmYGUTSHf7K4NFVBVI9zLvkqlE6XDOn4TecR3GJAiCZOw
pgt6XnRWfsc533+ACejVqsByzttXKeWBGggb/8d4Zn8KnfQlWV9ziA2b7bGYvmkSGByF38lKWJ3N
ulRwYbnp9igLUD43LJHHVGdWjVYSi0g2ajDCSNILE+pBx2znhJb2AxhKb0AcLvYWIo0ZyXXa9lCa
8yO9in+PwAA9xxST+75+Uda1qf7pV+9FwvS9Ud+aUUFikNDPkDGIO90wQuNckVSs+Y4S5/2L4igo
cU65ZtsTvTGy6HM65X7D/MUJjOsspczMCkZcY62G6c6a66nIoJPxn5HAaof+2TEsZuVV7uU3xWBt
A7m2EuCx2CUSyfSPVPMyPM2JyoppP7af23mOxL27jC8YmePsssuzD6eqbVOG4tEVck27BIrwgpCm
kAummsyr1nM1MtQcfioFIPweQEee87G9PYzLGulrvCjHQR1X+mGjbxLiBu2MqiRI2Xs/F0a/U4AJ
wihq1mx0Lt/FH6sjDqVi4Hwfg1u2qCJsMaVzvEPnxoba8tgGIj/DNsX6XTdNZxh0mKVnPpfRj0r/
jrLKzqD7VNb/+SX1HG5dEbeSuzzwBx65ldKl9lPaFtKoMIn+2dftGJqJ2WQhGHcTqwMbuyVyOzED
QgmXn0gCtUBw4QCLaHm8RiD7Ra9uy2Ow996ELAscpdu72fCt9yGL29xU67XOzs8gbshYL1Kw+un3
8/Hy4Sb4gLyKz9IKeha10e15p0ez163XP2XHg5jcGHWNtmBjx7ofH/z5szofEFI7+Ciowl3KLLW6
m8M2nKD7ykKKkAKb6PuQpgSYhl05xmBBIFfTqYU5fERv32gDuZwxV+pzPLaNin/2LTX6INgx/VQ8
7IKShQ1qb9d3fQ6ZmeNty5IJDVMVR1YJ2MrCzH1etnkBgtN9KVmHgxYOUAPdq3GReNmhpXRSDlcB
kLX1Ya1R5aGdmCoO1go2laef8+PQhjBj1prZQr17Y18JBqZ9tf/dIOG9CNDQU0TmXXBC5nVJZ9bG
DHOHgUQ7yagxB563ssgB2SQINKh57S5haD3n0n01sLB8ak07YytnxMdxdQpUivy/3ffAF64MqgWi
yKLneS4CwYbfwmoKkV8WBRt9olLwU3VZMqW0lq9/fKP5eYkef8iPeBVdDWIFP+v93L1ZCoy/PEws
nfxz091f5ze1ZXwyp+i9+oa7f394K43Jcl0yFmAxRPSesRZQmvU0474td5q3eCHKlxd9CJjPMC/I
GoL3ZKQj9iZ8EqcJkqei9hzBBYmjRQlJ2hPTBteMOUhJywvajh6lYRe6kbgN1UBVuC/MhDvh/F7e
H9Ud8bHWdeO73bqmy9zLJ0F3AwvHa9lSsaEsS7nPx6JMJLyHsqutXQHsfCOQ88qe5sXntctKKLxk
BXZzvMwOVJeGy11FknRxaEUY3m3lzQk/SpH1wvC7e1OpwK6EP+UDFvsaxajtoCCWIgBcmnqFQx2o
2wCS02h1O8z+SkJr+OLhzcBW6mOzOUaqJTXTpHahBJiRTuEAy5DQ399murWeKtgHD6vMITcxTj+l
cPP+w/KGgFtbEXXWmb7i5GdSDr6uG349LCuOpvJCvQigjaHDvQ/1IWxfg6epIDDx0JhtsNyLH8r/
ssBsVzu0nWESN/X6caH/9pmOES+n5XvGl7eGTO85eg+38quvPKnXT7mYbZJNSwX1ttHZ8iYM26LQ
hQm8NvCFOq9DEEo5exbmftWZiXjQ5R7aMQQpsmMp9EwAHCUMWKOynDINNUB7xc1yzbXT3Tu7SDqJ
lcOmeR8JU54pHgXtFKqhmvXcWLdd/k4IJQ0A0VJTAO4ArT5snqfKBy/QEA3txj0zyQRPRX4xzOxq
WaUyoyrZVZeVQpHezGg3mbl++inXlj+TQ8o59zhTWr5RBjx9vG8o3zX5yMEwjIwUjBKbwtfHsxxI
DMemFuPbA/V4IlxGtHJvecvIhMge+lb0oqiDRRYGik81JUqPW1zZbKhCYq6L6w1hEcXnmSWsRBxg
/GGd8S2qftlN3i1yiNiPKKM9CMks4pO32KbA5YTKKr/n+ZjaKOPpEI296S0ZYgjf6zQQLDJq/loz
VnUsJkJAnVBAyp8sSQHzYbxaDwrgvJp9zYFoTFPJdwu6B1cgMNfcA9P24vHjrgHBTAsAiVbybrZ3
P60evSZOv1RJe7A6qOCS2MZD7251N0ZN0xOf/zmqQvgDbMEi7OpaOJ0uofj5Db0ZEFkNhrIv0ZJ9
uur0fiUD3jW1/U2PhzAGYnOM+r/6OZXNlpq7HHdc+V2DrCX3HjDxBPiI1ndJgrnRdgYI3YCwMwmx
FrZulVU6L6pKIQqllFGGPST5rZ/BdPD51MeIac/SjN9b6qKtNYLhgJkXQhJ+FkIoXZeKUtNP4JMa
XWcDuYFwbS8Mh3klN4HVAkBKu6t1aq0qSFsb3foyf/FiUVKeFiju7XudUt6rvnOTZIcrxEzX94Th
c9cQ67euLhpZLRe6ohvjs8lqvIi3rG90ojx/6k21ywet6t27hpZENk6opkDV1AU4FqcCvGg02U7M
zVwzUB3JEeXvw055Hb5b0/Y8X86dwcR+dxIYtuA6KDNpeVf8auIYy8Fm5k015nR2CXl961JYTPIJ
Rg9tS12CuQuTw2cY520YbIDkLf7LClfm6R/7rUX0KG6sWgQZXpE3OUUdmAxpQ5NhaM7zNMfQktD2
alcFHGOKWQmKR/OIHOmM4S6nB6BvA9ayLO8VMXAvWV081SDqr64O0dq4HJ9f/K9vGAyPdmSPifuR
nZbXbOwyf6K4KO3rm59AoeE52yuLHaCDneViC6YffN8T9wxPNPjP7uga+IQPdTqLaSeO2+ETfJEt
9KLgAx3ILjTO9vXK6vcYGEwPw53TyXQNSZMRDxSqHci02gmwtGLh73/34am0+vbRzbCmAL2JXDTx
XyBcYN5pzTQF6vwQSykKKHjESxYZ1BWaA43J7Yp6HrdiDmS4gDGZQtkk9x/6rp+EJGlQPj+wk1O4
0JdZ0OJPpsErxmwYd2dkEnlP9HEmsTIWwV51uSy3fh+eJyhaFdskhJP8+h4VstbEHQyf+MgfceKq
9vJzBcW4AB0qV4OKVt+EWaMjck2jEH/iUxWfhA9iVXKQGNI7nzqONhS31TfULQLr0Z1MCD0i4jfr
m2oEza4zb6iFpLaU9RsKLT5hUGUqmQS5msc5CXaxknbz2eOVz7He/SEOGI6rGzhUDJn+DpPwRYOd
5D5MunZq4SFB9H7K/GicK/CcMkAvwMMYUvqj87DmWz2dqMIm1zXIARM2NK/+Q35bGdK5KiIJ7/c9
/eXNB/+ZJW7H+Jh9m/ekwx8J0WSPGwqZGSStQoVqOIxyZu/ZtVVQrV9uhDm+2F6ECXqPKyA14lhW
1r2saDdG0srBnmdZza4gxnkE7PvpGFPCjXkIXLiIex4H9KO/SeoS//8bTZiCnXSq7+LUdYLhHjvq
/ub3mzDACy+teKIdJE7c8rkQ7gpoOpZ9As250ZRfbH3TEGsGMK2j2FdBAg/8WX/PXIuo3wZgzFD1
C/WuvmWbmMmmlwaaVElGt0VORRq/EqRQJWd8mkGePs8vqVtMQDikZBYXoMbqPgOnL1VMZNDujsEu
VWUbxsHhtwfqBDLGk+y/N36v10H2wzcrmAPOrRdHJfpUeQWMlK5lhgWHEk9IEORrgTSrgkiLamUl
YLkXEMv4t+0r6bJHHTPJgRFk3cJ0g04CLGAYQYfuhhrFEnG9eCnDTyA7Ui8pEi3moH4zECPb4de4
4HPyUXHEobe3J3JoTANMDQXAF82SeA1yuNnnAN5tI7golt4VWcFm4Whl18bs72IxgGva+4Gi38fu
INYeOLLSoBMpRinNL7Dw+1C9U5nQIfFXysHiGCMHJkmHWD3Fn5oYwWQk2z1a4xPrHWKOqY2/H6ql
af+zvtI6nJUIaEE7DpClP999gqR6NzsuYDH3Q3jxLpxMwNgjaqflAE3felV9t8FFhgF5PSwWslob
nlfRM5kJQzc7GAAbgMU8vfGmf89SFwvPnf98OX4CsZiEPgDZDbUOsL4UXkR4RmnfzfymiwgLU/9T
3WCBf9Y9S2quMW6yJzX87pnEOIIZidNRDU9sIFhj+iNobEcTrMtuM5iavdeCcZVXqGscRBMSquY6
LgtuirOwa04WFTJkP2KPn5QkIX64e3snYTlCeDHSzG6SOLQ1ZS+IWLwkk5kR4hT+wOBEPJ24SS68
O/5/gfPcVGiNsZpjqa9EP8CV0MYNq1zWl5YZLDw3Ep9e8n6TNThndCEBH82nvhwy4CggQX9PzwPn
KjqJ5kMobxz5VcWwOQF/9eSK83NNjKb6af1+Nuh2qIkq9Isgj2zopnXFWoIABXtKAM9o612ttdTE
u/O6PqUSv+zEPbxX5O/pFA7FqdxQ2cCWwJ8yyeH4YrTKvDWkR3DacErF0gD1GgqVwaiJPSq3Y+9n
wxA8AqW7ALQfz7q+a93pwhbGmcjPS2bipMWPt42q27F0+tuWsxKKYo6fN0/WfCTtHEUSbNHqe16C
I2E1xhkh7wGQaGDOjo8ivGbLWbxkuvIwig/jkgt7I2W7gRl6ULzoH7meXxvlkRE86Ht4Ev0NOLHt
sVAcrcdrGOKPsHmy0UZp3W58ujD9BsaIKa4s6Hm1rygH4FAun4yyiFuXm5/4nQ2E5F+6w8W58Fmz
xgPES853RslbEMe/KsAOmKKnVZC/8LTaPOmao+moTzCNnfdyYdMh9QwEoftB05ljQwRW4edB5SlO
/hMP9wA9YREOZ2G+eEbgRSUVzS3njhSLs1lvX40eF26GlQCNoPXjPXm2+oyyIzPLtLqVK9FhCsj0
oVpVmhuk42s4YNryqUqJ94yHkZbXAUxxM0mDVCYjqrKCGq4GbuGjP07D1uj6+YYAk1pj0ZnB02nt
2F+RMD8kvRpzeIqWXYJa1rB6oM5d0kpX2v6J0V6aChL9juZ79gImZLA3QIVgwn2zV83CxvysZCoV
e1yDTX24rqkcApsuwmTN8w87J7t3sUbK6RJLJIA2SvCEXDLFb04asXa/WpGaVxtInBlcBIvBhjxB
xt2b53GzEz4s5ERZcMhQrzrzfQiCNxAG7jUpmc2O+OckPtySCwVSdcREl0CtLRK0y7idmVWk52Hu
mjkaYCElC81abqi35rHPMcvHKFlyor4SZlWeLmwoYcPsBvw2PrVlwQL+wDVRvNCK/G7Y2lLp0UP1
NyRcz/WesO3u4F42NeTLMV5llDTaXs3qMQuIxKqsyLcIsodSpo3CYL7/Ki2lnCHUW4+VxMCSWLzN
HynkoaFUiI70YjeETYwagbG16xcc4fm8uoxHUbOutTaED1tOfS6n6Vq+N0UQfRw2bLuO4Du0WFCe
TiOAlHIFA5U2xrz/KV7bA4sztzUCBcm5uvjSMVcmxFO4LEcbZ4oozM3PGXtq2CKA/Oj4kdLTLedT
+NxHpI5V1BUIAErcRoGOExyvIgbPjbiamLtecL++aOpVOKjm4ZmzcN3gYKJ68YJhi9w9yDu1188/
2JduvkZ+DQE80y43dqFDCYrOBtiN6atuL/wxgbUG3a0HBOEQMlV8B0lDyTnVC29DEX2vPTi+iY0O
s12qSgBgCRp4BtFmH984kaE60aszwPUpclYPINa62kqOZ3zLdEFNlseSumbyrjibuk5ooVSjJ5Bs
xH31spPoC8zocdYyY8QnDlSr5G8ddZjN5jlGuQDxLVo0VrXj4djemN4OOoN6PtZVNC58M1HGACTR
A/OIB71MHMyZ2R11BULjqD0XdG5TAqcn0QvIWbRwxh+qVt9evMY6k4SS9Vd/Dr1OEdXEG/7Wq/MC
/Wu6Vs+eQ/X31YslxwHc94Ck2eSfYml2xqF8oS9KuNAL4rP8gfRiqSynrTnSSBzBAY/P4IOU8jon
M0qo+BjhWEVRpYjqGEvS7hcc3eC+Z+yTgE+zt17347xfB1Oj0rofaT7kn78CmXWiwR9k6FJLXFBt
1fb6ROXXBFdoxlNHQdkdBBHEpYTqKesL5Fry/DYnlmIvMGEKFmN6Ww3CiraOg+mFtUHqXfIlXhlL
HXfGSKV6VjBI1brAdFxtsJh2qxVKC3VlYt6xmvzAudhWJxD+ZPOZvZFv7b6ABG/1mCA9HQTLprLi
LwDicejgmULYOUwrDjf3XXSFjT+zvW9kDrzYSF5DqKY8eV0bMAGZyR7KNnWe6Y/6mKFin1o0mEIR
emIjbNfbyRDoLRmnYTsVfDwU8s3rorVQu++WRegznhmJNLVoJhN8SPeoOKJFEOGR/HVy8Fo56h7g
6+XZ67EncbDZNL3YRffBvEWGXQ1Mr1gH8eLOfuRWHXs1sANuytvU3/hWkFqV2iM/oMSzCj0lmWDx
67Yye4CGtfvIeFXE5YIEqkCiK1M4jGAczBZ0v/+YESTJVLTf56Xls52wEEIHBoDM0RCo+zlpNJfa
b5xnrcTb4FBv2RqwhlccYf3zgZqR/echnOt7t60HdoX/qAzU/hdMszj3rXD9yaPm+T0l1x/SAaly
HGv49Z/5UfuhNndzCBivVKawCe0HfM/ivMAPQqB0ICREBRJPoJcoNawg2I1CO+zKk1yQkr6/SIIm
aXXiGD/dOc1YFDmtL+6KIB6IfpVG9M6ZLK4D7dpdQTfgzo02A0EJDhvKvcMKLg6obh++iQYPEA2G
EQ/Mu9yqaeMXkAkGIaZ5EPWtqdMqCBam6HMlBgvDrt5a2D/4gXdKRPi1L/oFTGr126hxgTrkgwUr
9JIiX7kBOyAeKCPmUaFzRPJG63mQ37QM5Ryg52LyOXV5fPWEloorPQdsKe6VODma9O1I+dugCndP
ePfL7x902sXb5QJko2M9PeonhTTCHGKaMreKYydgq5rmphv2BcIDbbdRG5alF4Y8AU/3X4VqlMO9
T9Kkbb4otRHmUb6nJhG1M6AJR+/jAMitdDTnAy6PkO8/K32JHiXjYnVERjCmGhyh/wp0oD6XubI/
FygOn0oaAEbCwNyrjEvoXE5oKuC5EYMoLcqmzXfZeWHdAMNY9zK4DPtU4nrVkS2pAD3MBDO1Eegm
jX3e8QAEu28ALTwYoK63WWDz0VZ88Da/csshrsqwleWnpnCqBVqLjYKDdkLa4avp4Rq5uVFD9Edx
DPy1r0zfmD7i6/aJl/HnfYMDQ2VBadMIOADzF5ZhIXawSokB2oMwLKBCcybRSGanGKfjz2BRF+cz
KdVDhtMskqH8HnUeTYjIZirydwYTr3x6LvQVbTZoU9gcVniaIwkw90SpTYb8HnOEQqSxGJ5hg4cQ
X7ws8yn0WX1o312NRKNi0awkO27AFTp28/fegA/cJjI8Yn41ygkz/iCJk2wL2TV4daaC8YUCj25u
x6L3A381ktDS5iOUAYZtEJ4swQ6a7E/0leDFgDBaQpO2HHXMeHK/AatAv3VH7fQGwqtfwIxgKiHi
wJbPIcqTnWfmp9VzdE2r+lYy1xQC0EcI1EQTipN1ITDrEDMGMhsmjbfz839Rj1YCplISn5/M6utr
69huhzvuVQzS/4mbJbwgOiENCXz1VuRlmUA6L5idkdHFwwkZXIFfGUZO/HeP0W+9GUy1ENisYLBt
L2+R4j8/EFISCdfHgsqqL6vRuT2MEwBxGKFfxU7vEVNVvXkFcXa7eVptO9psdsG60Ouk4zu3nSeG
jpFFW3lF+TIGzTCR989qKmhHjCMpTm1WjnBLvHPBSF7GXetfbmmjtJMDKxRdsh6gC7wQnJrCERiB
iru5H9++wph38qJaZYIwrmcyNjLCOrFtkL9pUXqkyBP5YWc4GYC+jOfa3X9jTGO6b4dhPt7lgz0+
NldAUtTdabPnNnpv1rN0brEBmO6S3Wi0lw/M0MliNbkENYBQqbnTR/TzcmKDxXOzd5vOS+Vd2X87
+JSZcMKVKcE4cWpDTCYU4rQWZeL8Zp5xiazfGpnWR3l3eHSBycrA1t00jVGwpT0IscRt2kIoLIiM
KoAfIZ7Aiqx5igXsNr2PJevJdQ7WO9y3VB1y94BQ0zhIxTjQ5CooW9YwfPwdg4rXlyXKhgNpJ/2b
N/HNvovlSPmnSfZIPAQQKsfmmsWQQTK7Cjch/UARt8Na8eMCmxj8XKNCSou8Efq2GtLvykGzwzds
HdaYfErvvdwL0OCABmAck3USaY52t38EEfk5bFweh3XuTu9wNHG4qG0NCGSuZ0gvo9AxrqHLUc8e
gIGW61msJ2NmIkZD/tLBu47lmeYjjOeaGcSDudN48EjSWKdW2bgR/XVfuz4ItOI78wkm1i0TurhH
ft4s8f2V32xTEg4DXg+VHHL8CMAhIlN5f5a/DhBjrCyQ1kFuUjfVYow+GfwOtzzMZRiOelh5S5FD
ketuXeKcbMSR8eEPTHNBZY9xwojiChMo41AkiHa5jNV/AG7dWf4b4MoLTlHAStCBHhCtk4xZ3bmS
VtSJJ0tV04SNB4Ulleei+/5Sfv/4Jn7WwPpvxk2MK5VsJT+6HLo0nXma5qRQrlWY8Z+sjpzkCSA6
yAGcJ3Q7u8a/p4mdxy/brbiBVK34vZCq5pitVOZaIbkCoBtrLxMkxkMRauzv+iaUKlbxvb9QaABq
zKYc/id5w5ZDw+V1B9BVNWj18StGbDTVDEPDlPi6o2kisHnRJw1YNWjUCHC/qlh5+eWhjak3CcRy
nX8fvpKWhcPVs/tVSGVpvdL3qJmwslUP0lkFvaqXFfocenUuGcco+Om66ppn9J70Ma65+HiCZHRU
4pDmH+WAUfDK9HIMD+Tn1T7DRHD4DCtYbKtrl1E0BhXx398dvf4sXOQDgjHdIQtLILlmfXCGo5kT
Tj8IQagGo67dN7Dj2PNR0HInuEjSfb6zIGVZggrNhmAVI1TaFMTAzlAZi6Xof6/HfVpQV65Hz8A+
X/FpdgdAbVv2eIi79XuVfO8NwDYxpGI8UmZdsq2UBx1e8gPj4gN6AlJoICJj+3H4F0tdWhZlkdxO
EiYS0TgWLwTC6rXTGirm3YkG8cHCQy6cEE5vqPmja5jZDFyT5Eeqz4PJJmXAoT7jGvAIQV7qfpN0
4p4t08zBIpzCuy5aODq5dPQ17I5g/KFkbTjCfuhLoecYQIHebhgzBg94/wBv/vVPu7Lm3SDWEWRP
BLDBiVjZ5yrOieanEPMSpYoUwcdG/b4SJ+o3cxxmKicTub50lXaa82r/bqw9VcVIEPuyxSZXTaSO
5RFkQVGWeXtgFpOzfd6tENye0SAFX0qUutUVuIJKTHHYRlrFpLqlem6WH7HwBC8zB/+YawWQv+Es
KEccbtrzGBibww2aPc4isCYGGClg3UF77w/A+1uZXjLo8xC4fjpk6hvUnqRChaiKFJ/wU808Luzu
mwyddQIEhFVVq27c/7TbEpDFf0TmG+PtrSX4/Sv3PIUk37wyLMuwCXxtEIJ/+ssgRGdf1Ntlp1r6
3m1pGefSF+86kq9onAqBbcv42ikz2+eOEkJMmHq+1Nv8YIvzI7pNfV9yELgXKTDWPVBLua6DgcTL
nxPcdI/JXoybQzredGv2MmcX4BWArfNnG8WBOGBVOTnVrtG/bbnV0DM8EMkKc9xeF51BuTQ6K1tQ
dR49QJ7eLkimw5VcZYSWfYuiMaCBNGGYX+gW3rBx5VkMDQdWuZ3Jaq7dYGGT9x7bR5Vw+BLu5os5
ORIx9YUytQwF8IKlxwrZLBJ7DPVwvO4hZR+2VKs0kVy35vDTrxAI2Un8AZKwsY8juOG6dtaEXVyP
AYTFP+aubmxfcVILpQSLlCBvhxQmu7z+djhm8v+OhN9U88lH8HE/PcPMU+drn0sN0r1sdd9y36xs
egjvwvgKA4fAzoTyP/uWB0x7N+uNj535kp+u5aoAtAp9So+m6sCNeuH+339H5QzdeBSC4hrKFrGl
7JxpFf2hgePcP6HBC7nIB4XKYZX0b3/0lDEvoK9uTvMnLAFcjTZWKKymcoOYeauDtcqgxNuV1x3i
2PNFnCe/7LwYkSHOv5ah0P9voR41xRcSTKETz/4f0ZvYZf1MWXJitSVqiIVcqOiozGRYoMm9wDj8
V92rKPfNMfe8TpYvXSY94JE8f+a1n2R7nUdNa/EBP3/sNmaJjMj5Gfl04/+B6ndj0fG22R02XpUr
5/7gAZZJ3cFKJj0vECLR4Kq4WaiPtEW74GsYPFQKsxU6KTa2iOOL1HK93ZSZKrCkIqEIqCLLgVKv
j3hGuBt6PoJBu97WFFWvDclcEl+fas+EcCMSUP5UqMDynD1Q1Pd/wWyhfGWvLYiw/T2AcnXi0yJs
QqrNfagFdgoonUqFwCIgpoh/Tb5CGYjNqz5yNuG9adlQLW+SN/y7N5ZV6dISS/WpdLBY/OtSXu3a
Zfm4AkVXBF+yrXhWl8Ip4mHUEtHaurWAMrRpVbKTkWc8rkjNho+oSavmjdNHZqgYJb94hGgcZvpI
uXaM+WRZV58SO4dB6sl8TMzqEjHzpbQBdFFaf3SNs8DNqX+gaxylHDOYD9H7c5PW8CZXjrq2AnBY
uXelJIcO7tBEPkJ9l73nWhNRcCYxTBnrG9CvdZBjjiA0d8jlXV04Lg4H/q1fyII9W3h0jmrIfgn8
zRTzo132FNYZ3dYGz24eFJ28mh1nS2JAWSf3T2bxWbCiRdgB+xdJARCwrqjoJtSiDTEg0I57pnpA
T+bqOzTFMP3XN7dIrHlUV1VbnAPsPlGGIU1ielJMoatXYm2cVqD5gmD37i/NdjMwLjfMdolV+8ao
kpT2siWh4e74bT/Oo2NC5FgoOrhFWToR2PzVe7usuD46q349Q4x9oA+9mGuEusStP09jojBM5Em/
RVm96TCYlU9WHIByGJ+Kd5eI2ztCfieIMPs0jloH0h2Z1dvu82qf3KuSfB28f8BokzIqt4DA2QrF
0akFFV645yDVFjsQoeEDzCwudFl52VK+YruFYmy8/Hp53kwdlW6pTN8nLwAtXcuBW68QQN63vcLC
BJqEsImYdJ/TO1aryWvh739hJl6ja5xLbbxN7roSfTzUX31WUY2Tz5/eOUlfARYhobIU1VoRTPVS
0HDdwCGg6DuAfO8A3yOFrmlWhSc/hPY6UxAs/8ymEsyR0HN50tP2ebnc6j/vxL4Yl+sfL0XYSLNw
nlzzeyLQ1ZYlo87c8WDz/vD3bV6ZVWcYV4AVjFbdZM/UbT4pQkr9JfDSyE5X3S+hFhP6tCFwCWVz
sPXeTIlsu7/KOafzJcG7UJknRfORwaJNyfy/tuT2G/mkCUl73PxizMya+aK9pCic+jXNk9Udc+BB
+5ShCnoSTbYRD2oAtGQlg4lF5SGmsh/31ht0DH9MMNvTEjhjEBmQoGIGz7JCYTp6nwZcOfnzYEW1
h53EsgRd0QAgx8ROEsUNm30M8mWahCaeJb6A36QHFac+Jl9nJ/H8vvtyVxjcB68pZcfvoTwP3GvE
RlKTuBWp/SqesnBAv1WlmfJxcDLEsAPFfgFr/8QsvRNOyz3ZXyCVnWlZrcJ4rJK/i9Xf3i2O23OL
0ouHx7kYu1IGJjoSxG2a6d6KgMuM3QN2osaAcH/w16MB4V8F8ifq18ZNCwKGeLq7n6Rp80fmznx5
QlW8XRkzk6srpDO8TYMUqyS9awN+FwzlynXypfnextp4h44r94TmUxOoQRCbo1j17tX9XULE3usH
9gFa2RuUkuHeEXtv06UgNYDp+1MnO9qW35rl+NHP6v+eyMXcCoHfzXxhbNwslHy6D6XLP+of9mlm
gv5Xom5PBIUtc2uRNO0J55esDrsClpRxKMRkVeAyw5B6yZZvIIOFJ0Ug/fpI84v1hJAD30lw22ov
vd2XciYD0EcbPZnPrCyyQI3x+1t3fGQ7Tb7hNmGVz+cmXCpdkAQoCQMdM6QwCjULMOILBwsDs268
EXisFfpP088lwXs+SkCKR0SP06V/3vAImAkGlAX9YLGrCAOuwg/bx4zTpP/VreP8FDjXUyKuHlqR
yz80yRnjAI/P9B/JlGOUz/7LnVtE4uY6uaw+JDD3nBHFolOOeWi2KarLRjY9ohDHHsLYNvFrfe5c
hNwoUvR9zR9QvItseLz3HQXiOqZiiycHlZp+SSvuZFFqOBZasAQ8CInfxxnt1+PyF//of7nYgfw+
8VKrMc0mYmWYx4Ep8kh8+DhVrD7F9wnOsuPvHcWMMND0vjhdnfk78SIvTkRotuGT4II0dX4YPzSY
RLPQDT9B2WYdK7KMQXOBE+WpkmTK116nVRq2Hl6VrWvzwSh4uZqkwJB//+DHeclc5ukUVBuBrpyh
F19OoS6HIt3/fMqh9KG7ADhSzx1ub138fqK7LtrsUQ8kNrzaVHS2zgK5eixM4MwAVkXBoVYlLCZ/
gL9yUPED2vMwH9oz25PnGK24C9MeEzbBJFlR6hVNCe/uemAvZgx1m8UU5BBIa8rc9cTegoqwjmk2
WKWPDFVMiqcQHwGF6zwRXSboQl4pDM7Y6iWGnH2/ASp7gYGKkYUuhN5nrQxAQLMhKVwtgIwd1pf4
g+3M2/wkAIzqyqP8anPeeEsPn6/jOT4WAVepc+Fuv2v+D5Vj5cz/md3xnzURV0R8LKQk5xamtfPq
yPXXRrxFlHc1Gwou3gt60CBzdGT3Sc4qhgPbFWs7SbXPa/V4S9hgrppcAk1Cx0BtZPp5rDelpi64
WH9bN8Pfaj5MdZPONjoMwGfC+6Okr8mNPIqK2r7VKpgT4/v2qdRiKii5cIebdbtkuqPjqwGwtlcp
37E/OUcc4dccNWJfwcecfxCIJgKQqrPiKv3lBGeAyodRSRWpOvpZSFEOYrAXx7KxCiDbAmCf2/Vd
Vh98AyjCieCYOlFyYmXVLwZfRCFV6nqq1uvl+ZIKRx/WTFJYE1jPqLvmBxfD85tmqAJUj9BePHOm
uDeQrcvu2k9ZBqcToya2hJVPEzj/FoSxBy3Q5W1Zgiht2BzUoeCgb19M9iq0G+eSWGrcejGkW/Vc
iQVAk63h84oJTKc2q3Nxno4m3TsHWbO/UcDJ7bgMJhlawVh46Fn0CbaeficuksG98ej+5FdFwK9H
uyfGq9QU6xH76V95XiVK00+xzkYq/rQPgW3NNThkEgYBNEnK3caVJgH0JQz5plWWYI6ltyNQiZrH
FqQjMOWrplp8wKdz30kKQMFHWN9u/vq0NsflqncFq4JC3x6hEhMoz94sKlsXKhptEbP/BDTytXKQ
0BTHiRL8RT7SbjNN/FDTXlG5nTRUTAnCxiiH2Kyg+xGSQqsG5YcVzprEHrWDbwCpSEF4dYb4SST9
Ij98j9cLDvBuS6qVLwNkWzH5Z+MqHc1dvk9qm32Qac7TvoB59IzPKEBswVUPR5dfcEl+SIn3uLky
QQOHH+IxvMwliToi4E6JNBfhdFFaMDh8Lvh7XeVBAhJVkCyOamZ5nd+Jp9kwRWykyoCgWczx5AzM
7jzvGKdGFHCWZ7b/ThyDtXCAzcbU16GJwbcESk5/NayvThYLg4pDrWoXX0ovh4ShquTguJGE4Fxp
guAxTnI7Wu+5k/+81kYBg/J42e3EOOJwAxksgyZWDSvAlZJbJ2bztmUIFLDxbIh5a3NhdHHmNIv4
0ud7wOmTk8nWS4UL0tofyZuNaJGYbvQDcwDLlVIhdiIa/Rsbe+/anqCokFmDgFuP9D1f6ciJbre2
Or7Dy/UV/jC7fqVv0Gd+WBDy5masrrZFAFtHqFYwWRq01EsPeW7CdeBt4CqyXve1UTic50m5qvqI
Z8+Nt/NKvWvRxsQl/UXzPDDvulu9bVVzkAkg66xZHagWfj6X6v4hAVvrLaQr2lsOnk88xpJMA9Sx
TxT3+zKDymqT/cTkrQCJohpXipbmswvSNPfKdFARm3xApfkkFdX/PsbEs3df9by4PXqcnF1OyO/U
nk/1tntffePXYi5WEOOuFJsJ64x+wODNmgaITRFduXI7j/sSTvWw86/ZKrqNfOJknMn6+kjLxUE3
uvZCzuZaknBlCATvHDEN2WEpFxCAQ0WWNn8GGY0yBYVr+bcSDtrrH0gPgAcSf6X56wUl0MCGOKuM
MWP2U5tZKXwm9ITE4UVEK4Atn5lIxlNN7U1xAz9IfQEZA50XY4gnMKpThmu0BnTmFS2cn3L52rFQ
USennOCbObr9aX/WYbgyAbdf1RH4LsRFGjb2STm9ph2KnqluK4he/wwz0c5O68IsxXw0nTLwnzDq
gTWOswQlVdozVSr/sGvsuxMy9mh4kCpqDCxdwUdPfcC62PGiTzjv596JaosEYgu6VOd/j/M/Vx07
ZFiYOKlGZGJL7nQnZTEquP19KHAxScS3fVyVCPrajYIXGYAoUDRzpIaswrmrTOgw3np/s2CV7BcP
aeMUb/Fa7pX8hbVyVzijeMrWbEFdZwMi+TpP3VJlfr2iV2UPGfFuqcYxTdhEVnB85WEJW0IzCK+X
pU4CnOuwgiZk9CPNmzd51flKBXxXKNq1qVNrb5w2Y3KHdVx44fIrlia+K6jCEJMmnELWnMEO396o
YnvbxxbbA32IX3cQoEh/xa3dtvoasD0EO9s4DvSIdBjiAMsEVQh6TZEjG1yu8aJWbrFxuMwOIUEJ
dYxe4ZTbfLNFB0li+6ao5uXdtFRBbqkYAuMyCnlfpWPXwFmXPQ75DEM/LUVLYfOss/UfgVlZZUin
oG9OG0uftiSi6xroT++lBtsb2iwLxrDi+qi3LmSlu0a1klhRmkNuDnWRCWBKDLnIuFlCy0upRb8O
df8Y+SRdgork10txnyRbtN3MEwRhr7EdqDRkDTy0szoSalgZydQ+Ydt2Mem+fZMzvTq6QXRwDgux
4uYUHBOIP+flnfKxaaQ9Ui2dXe2/BA0POZ5uwMIkmPX/UivHnNewrcQ9ECywcbf2NjBbWIc/nEcl
OxXcPEIppyZmBRg4PLOPc/gNgHbW1jQjNJFssqEUY0OjsAcpCCWWJ3EroZNkXh3b4TNokcE0vKlJ
iZylAR+2dLcusYnotMZ40jtdds7kNk8HQ1B2e6k0/2VKWcAk6yO6f8l4wpVmuVn/vw4eoCST+BdE
VY97Axkc4RwZ7YAg+jgc/OTHPKOFC+iDlYGbCAu9APPMalG7QrCjfryQTPwpD1pmNqkR0CbL/lq7
ADiqUXloftSycRqnuQZIc5Hwps3i2m0W3vMdDpz1xB8YZEa2vmy/ndFJSI/kaqmoWNluFvtdvLvD
Jpq+j0YLAXlEVqQ7H+tVT1/hD1Ou8z2H8ap1kE2mbXX1ff/v5js90bbCNtWvbYtXSTZmqL8oB22Y
A3pdntw5W93rHqVomtR4I/fJFP2GdyKSWwZi1ThZnEH8iIkS/dwg2YPQfqkGXZaYf8xPT9u0NnNB
ndS2FIct/2/dYSwDLd7bsTf3Nktw56jut9IZ+LgwBn946KJTJWB3S4A7L1sXEORjD6LAZlPPAhJD
Z/KW+jxXrINRZpk9UwmLWTpb3+xsgsK4EnCN+NOmS/FfMZpnhFiyL3VKE2nYHpxvDLd8z054eKxG
qL0+XvCH7VEvIHHfn/2MsTsy0JjS0VTbXmrVglk0Zf3GM9rL3E1nXnZvHTfsQMUn9kVlINF8kuhP
QaVcDZnTHs9nxBAV6tOMz8B9m1kwURy3/hgMHx+irjobhbfTBeK4tJ3IVYTHOTHahm48VjdcUWPh
RxZyhy1xrdcumg8V0QtYoiTyS7tfQhi76R8QFbcQJwtMinI3wgctNGrYhqFmiQfAW6p90yvmUW6V
rTi0VAAzWbTdje82A6SrqWtaF4n0p44+99QM0gnYzGIpDJiWjOlaGQjrdOzy38AUOWv16ST4gcT/
ZMm70P9FJ1OSxHbvVMBedhliW4Hcc2Wui3+OTAFCohcIJxmhTixuRtgaFUCtNYh2uCF8D1tBxlVu
u3Nk/tCxICl+e1Qnqyn/NktjwSxgc5pZ66JIvFyEfKr12TuO640M8xbiV600hWrUIKw19SsVsYub
f0nYl6wODXJRBTJUUT3Fb64jOYiHRDTSZHSzkpFqCr5bm+TFRQAoVd+Dq4XRqTWZlwaoyTrG19Ak
8jMcQqQzwtwllAV33y2Q0cHy8zRtuKmF3k4cbHSLfMF0OTKbefS3Y7TmElE4Smw/xVRfRiouktzd
ROEW2JvdplhEhyeJDS23oeP37gftjZsw0vXkfPU8ChfHngxGmRyfiPAFX2mYEDhym3l+6wSq/YEm
DLLQhJdDVgwTKkLczGxI1bXoxG9QP4Fs2nOhO3iIvJgFycbdUH2NjkZeiq87k2gCjbnbpNclTjc5
VKNu29tSIRaGRf51uugNfyXRsGwEYJNhgnjuwLH9HrNTmVk+v+ieNAS7wdnWMHgzXiomMDFi7mNJ
5HId03kzIRzkMU+2+ozR5PgxnNd6QIYVxmsFdCeK7eJTc6mWOLAR1G1tpfG9oa6/8pweG0xJ7kAZ
DF+gj2SBdKg5ZtGtE5MHbL69BjJuTVCvA11sOFxbCc0ZarTsAfMYoHwrR3ARCd13jvXjdp7sKQzB
VUjqKBGu8D9QVD/X3/A3XI1T8QBFwkcmA7UnpwDaKRN+sizXOJoNHPWsbHZ/evSamXeG/pd2OJxr
kHQ7DXLgrUX3oJkRTpL0vpj+4VPfDtRz+LgMF8T+CD1+Uvc4BShMfxFeg+BJ6kOUtrUHnBM00pry
jwdkzkVpp4jh5QyKz9Jw32KEuc3Y0MNm4PCWCb9djVL97x7q2Fk9ZdbpY6d5yccwTtuP/qSMgw7g
qNUwobwc/5LCRZgkj4CQj1hwuG4r/YPYGSkJaUFwpwbgwREa4FckpSyn+RQHf3TmgRjFyCFZeYNX
P7ndwHOkmTjVpG6Hb/zQXmO9Vm4DAfV+aO00R2+mJHT0i429zm30urbAlQxN0L/yCotNDW8zVIC5
Dg/MDe1XI7ylcMmD/0dljKLVTE0BDBRafcA5UTNqos4eL0CGngpAJ625VjEvYjT4L5kYt4dR5M+d
r0cQRvLr7Yj2Slu8rPbVT8xmjH2AatoOWASirkHhkD766Xnd+WQLVf4G9L6DuuFEQxIw/ZUNoz+2
ctTEyo8gtp4LgSdpe5zsWRy53Sh0odBTnjVP2RhWNYHODCs5n3f2LwKzeYWSsNlQS2sRTJ1qchhM
TEiECpqP1XKRposqNom8Q7IMxnSM7tJ10ooldu8EnJKe6dlwNOHZTmIlSI9JLlEVc/fl578tmcDJ
zCjM4obcO++j7Yo552M5jciNKmXhuQlLx4pDVXQNNxIcgeDo79fwMwrtfNlGadqlVlSu9ZijO6DC
Lj+7Ild+29I6MYSvLSWIxzkH9UhyeAIx5yCba6fWxa3EbTFxiwaV87eWuBv6fozrFJQ1MEhrr+/0
g4HrmfWENNvbVfgN27HlcI53tS8RYYpsY+cFQQIDynipIJMATb7Me2C2AHkDyOX+EnCAhUhDV/Z+
TbpiqXYS/+cNsE9TfWwZnBxrglbEd5N6WlbO75q3kBTUt/zoPv2hvEB6MAZoIMLDLWuEu4aqFAZ8
qXA9bHdu0bKqLzzY8HueTstvB23jgthoJYWI5MLvTBP5xyWJOO/vNZunasp0pvgH5cXKAqTq9sVT
MECVkQ/PKVJGArzfrshkjGXAKdn6QDI4I72a8E0kn7o5PNpvnXZkiF6Adgh0ptENLqEkUQoDwPHl
M88RsKfc3h461zUlDehHjur/q2gbdBpOHCUxOjqNLqtLym+RHgEKin0nQCV/oD9SW+4FJRYcYUGb
GYY6ywCC1Srz0oed5VRN3WyJ6sMOQpqEWZEVcq2Hgnr9R9lnajn11Brpx7168PC1HlOyxZbIHyEd
q+8bPWwke0OJPWxVBpPvobbIWyGzjFPbK7hcUNxf/hISPfbOO7kzagoParqmGvo5AMh2qCeLGmDm
5EjPcztGBMJN5q12lnaPUMMalUE1IPTgazYeg2tsMxEkL0Zgq2cXKOG1WpvIUGeTdXUZHwYyCzC9
KnlZPEgLFuj2FO4Rl7rj0hs8vaRNUNQR0vxzveqOEiNDUPCmRH8ZnvGoonf/zBkuAXQ5q4dkJL6L
r4Rbba8u0/xDkAg2S/PceUs05kOR/UlIF4+yNcKtUi/6C2LYt0MopvPiJSuWBB+tguE9ShvfSbci
SYeSCMcBSvDWED2aKApqdLMpvCotfVl48FAJOuZEu2LywL3R3KWyfsWiiF0GZIes1WO5PlaRsVU5
6D5mxszhblckWgAb55LL0Em3zK4sYk0f2gwkVkIT4M9k0ncTvmf4CeGSmeHMvJXSixrK1E0Skuxq
bP+/ujPqwMEEXKJYD/rn5T4a1qyNt95VP93mml0wARczzqEyIp5uqAqJ3S/NEKedFoZ1WVhIaXRo
3jc6OR7vbG8f6aFHV80ZAGck6sailoiR2Td3rx4qERltXhLD76DhPr73SpRkQ64eDYC5dRKDGacq
a7Ps6012FfsNeweqp3jMQ6WEvi8ANgY7ce6VIulPxPPI+Ec/Dcj8FyCOp24iMLeuCeKV+eCiF/a1
xvMRKLXfcpZ7Xcq6OM9S+dc4j8uvYe3RTxc5zuKdSxwNS4+A4TzJILwy6N8QsdoAj7C8Ud+jNf9U
GfRDnAswdnB82UC6YRdmJywirWX0L6yuOWFSaqLvxJlXBAhFW1Mr9/WUL/aL0w8M2uIF4vsnl/Oo
N55/FmY0aSeTVNpGu3/sLEE3ETxIjjmxrM31a3dRwBLv9SxCGADy2zLjri4etJMgVBlmAg6r6f+K
2l5szuyDNSIsSh3+HtD7dRtX+RWF7hiwgvqW7ZRtdHV6ScQ3HC69iccAQVaiNNpEjqptgPWIBKsX
DaJ1WKD0um+6RhYOAaznh/Q3lq0DtQbAfKkHN84yT/JXZhuUo1RKWjf2ABXQaJ69W3rLrx+iJQMG
/6hdPVai5Nnht0B2XglZx5xu+neySTM0BnxVmJQeIl/ieBuX5nrZWBxJThUo2CC4Bcxl8eAKnYyK
Y1NrnbUs7MxKrHIkZ/mMMVv1CA2d3bHZkCgXkyrf08Vbk+ZrRK0c7UEgu156w7Rf7bf671ZEaL2c
SaX1OQIIhTB5CefrYGFnpaRorXkqsZ3NpwQXKA/iFdv68eMZRUeSs7V70AvHGiqo3Px/pik8WfHA
ZkHfAaBI70ZEGgO3ONLGUJ/pmtSovDl/S72lPEyuJyyP+WOkwdf1SQXzCpTLpQurgOrttythaPuU
jwONkFcIVfMPy1ZTZtnmLZz0kkblFzFkiKNExbVbt5X20aY0zl03adFC/nX/mYsOlHbwfdMoqPJW
36ZcR2038JjuDNGvg0VGR4YejHOhRmOJ9m0zP7zURgNKVFYAmNcznp6S3L67PMIdnrSlSm6lk199
HPO+5uyfD+15eCistgJmSl9+OvoYNhDYTSl1ylow2H/2VgQxz/0TaKQ08bjD5SPRg52gRqA+5tcj
zkNp3/NuMzYFs8Gowunv+hRzAUL1mzxlbzIxwkKHazFLDPmdPeUIJHvoDQEZJEtlDYObALHMp++g
IsByvadJj71o1G2NlY+DrzWgBwu0UlNUqk4GhaWhDijrT9bgNW0EwIo0irV4RNgssgaKXZU5/Pnd
zTbT3btav/O1MZDyFchY1jRWZHcg/pANWKCG3K6ZBMh+r6ssVHe0GFFsR76KBC59NcJoqteDwx1N
EwBkkyykgFND32E0HmpmJ04P9TmZmh29J2zqhX7cNzDwzxMn/C52OGFl5sLg8lJqWZlh9DebNXcu
/Bln7a+yr9Vc1IjC/Hs5T8VPta+wB2Wu0LKUYWcryYbo+XDcgRCldjN3tBMlIi2oNIOxA9XSDiiU
7xoa9T+YjCXGw4CtdKsDYda0K1uEzp3t16bJUO7DXqIUODk6xwBG5G7v/ChPeARxTlJxMYhW7JDQ
5LQk5YsN9Utm0uwgA9JyOQQJohB5nm1duQS8NPoRTLNq15dbKjYJH8SkYOZ2RyvhS0yIPEwAEVbJ
QwBO2v8gOCEySnuCFoIZObKqGTeEIeb+lMvj9pAj85KUQV3DAAVv51f7eQhqE9JJp/gvEXisTAQ6
mR8aNfU1ESM84fcfXPEgKkEMPX+L4vTEd8ew6U6hT/WcdzGmlmRb2ToUDiqUSSLnrI5E3k0AB1jR
PB9DJLkKyMCMeC4ZF3LrynA2gQHFLqiS96vymfrsw7fRqrKLNeQaKXJTCuA0Li9Ne3sh8EqBMTcq
lRMaTr1QMcjBF019AUSdLaLt7Pdx6EAYE5hjv4+qP+4lReOfr107We8b5K4zbdZh2GJyWxDjfV4D
cZ83Cdcsz6K6qf5zpUw8vP3H816krtKyYzf2sXM53V7k5SIDxiPDFG5Csq+UQRVPxNkv4fW+5RG2
bjLkD7gpXigLVCi89AUpo2Zoxi+Wf29ObtaxbSgQ51itHNv6GiFOCTwV67JCzZKNm2n6Fmdo2YEC
TGdZgVl3nIdC/FHzdK/T1KroLtHLW9GU3/SVgvfWLps/z0J1JBC1xB8YysZi1GM01P+g/hX7hkLP
vnkK8IUzIsojZ9Bp+ctQilMuLW9cFD9XS30Q8a1er2mYxzuIJRr/CksQHOXsohztHPZchbUtF4D7
Rzc8qlDPMiwanjU4Df/3bsRfl7VyHy4rT2RaAqb+fbI/1rmQoOM6Ij8RASM3pL2cSaAbuGjwpxWR
J2u9uB56DNSZVolqEYndfaM04vRKItFUE01CCU8+JDgM5nRvXBV/YGlWT2RSs2wgIv7uzJFTwyj5
Ff5mQVFKjUcere6A71ta01hn2IzCOysWk5vxyfXjI5MrdmABQyVhzJiGdKckpaKnd3xrPENvkPJX
2qQxKAANEOFkV775G7tIXCiJxp1qbs0biRq6JUGzksQ38WEE8Ps2Hi5RKBrgMmbVsuR/1k6/FJe0
mQ+NnKXga4Idwk7ggwkhN4HKJs2C6mul0gChmPqJMLlh/02bysENcMmT5SyVD69RFH1fuk7ga/VJ
mbPWVFaWuq5dpOmXuordmsnOA+RbXl2YzXgAZj72eJA3QAEvNHYFA2VGSj1fumRgx+Y3gXfqlXQf
68btNcx1gNVS5RpgMDz31yio9O8xWHhKZq86yv0VxYshAnJ9psnmjlmyrO2gbXHnqFSyL3+8+EXk
w8AMhHrswx6t4CUVlPAkzht3SoF4TUVtly2r4UEt2pDjppr+zPGh44F5OQShViQUglZ9NOBrEb56
2zpwB0tHgb7rguybU8fY7cm+OnDZPYNJjiF2Em7oTOrC1nT/1ct0+0yQvIRvOy8bTmY8NOsrM18e
qF86hN6SgI75wvGTlNlOLIU7VFHISfKKxD1DFhnr+V+iIniIq+9S6u5tNM1XItvf/u1yb8XvL6Zs
jHXQzVtQA3cx9CkwAy7U8pFzMkxkoa6j4CBhkUcSs/lszcdPqSKFrjr2NBNaS2valYhl98lBrjDO
oQuF06gL9rY/ORTOI7UULZ2BTk5Aiwt0IpyOr5NhK2tBeusXS0cy9clkCOyRygLWjbm3w62HT1A4
WvcxtwZk9+384QNJrcMtLIHfOeWjmaz7k2KBXjCSqGD0ZDHgpRW104QKHYxYP6xwDCS7JyUvIQe6
w73/W/IM8Sy7nLaaD3TOEWBqPN3OoerZ3lI4h30nAM8epBVOrpz2DWZWtNv4WcvCYaR+fzCyrMyX
tQ9b6MpVtalEVUniLqeE7fGpAb0Xiioe9jSU/OszTe8XmsKaHci4oL1hL+q8sN3m01tgf4AQTxuz
e7nwEu72EjZ7bckF4ahqY+VNUE+EMf9vJ2WMFzyVwBjUanN6HcGcVWvBx5R6+v4scCeYsdDvuGTk
vnhGlr45dJt9o+QSrysQp5YtF5U1mT+9vAZSPbI/hqIbYw5xeL0iNvbZzSgvXdavOY85o6i5xrls
R9ujBqISwZ1UqcKG7L2WEJ7+ym4MXD3uyI+ZzZdxVhlaQs58KrNbfi1eNxZHME5c8zXXJgkSC2NY
IFK7fs+tQzLeZEaSp+YSCy4s68g9yUxYxEPIKhxsejZzA9hkk3MCCjAMq96bp4CXywgoYk/K6t7G
I+N6/+3cjE3ujAsIKXON6Q1PztQ821ohoo/h1XMObAOvKBkanUvLTrAaUJJXxAhDE/tSVugH/8nL
ku7Y3UTvtzt27h4qAnu9YbJXLvEDP/Blnf6DQbQzeYm6KAIZU8Gn1xpSj+n394idPktGpom7Ne5T
vymRZ8+WkkdxLHJbUQbG6u1rktnZzdin5cfXmzBJh2Az93Dcn2b3x3r2/d+xHXctCgfzvzfVn3DW
mPL+ISK76bvwQfHvgkKwNTq43q5SHuN/JvPSNAjNH+cLKUCugW+qQBy20ObKPjfai/GpckVhapAW
utF5ymhWeppLoRuYFS2z1uP81XamBVsJBHXX2WX3Pj9qJN8NnhAfRYMgcMunL1Y9dwoFui3txL/y
vXjY9XNgCu9xLqi5PhT29uiOtPIdRmgQdyCcJiL6e/vYzH9h6gQdCHNIy2QWy43PhOybL/I1OWI3
KPTLxYYb5vX9RDmSYQtMxAT9biBsRm/ohUBmDND8maXpm0Eg17zpkQG/4msMUdN9lmu7rLWRNY5e
kabz8V8f135i8mkf+6CLbINp1PTM4IdYMHHfEyL6G0w92kcspzJp6ZB5PrWQgsd7d/a3fO/+bbHt
JHQUPNtMkYuUFNtNcGNUX6/z6mnLPw5uAQSIMroqlXK7NErucIPzhi3eGywQB6ww2mf6twLIZKzl
6bKm4h0hsdmLaqUOJL/HuA/65JHkPwhTmjNlM99B1wIWg+oEMFI24+upPufUspZEDGOpSzRiZ9Ts
tnU8HdM+3R2FYX0k/b8m/Zgptzxp5jco8V/8np2xmsTc3WJcTt2H1LD+UO60kvi8oLw95bE2eLkQ
7cb/KNGt5Cv5dcT/9cqhSnzMmWiOB/qrDVtBF+fjZOszrWHy2kKU1BfYFp5GugBDvJT4ltX8wj+x
BqEfGdqKnnB9s3FYHhVMEf9HIXcpEJJw13mH8ToyRCZMRdp5J2DOz1hIWkwNJNg2tZA232GcHWiF
LNRANNZ6thf9p+au2LEQTpH066lFdgN3izTu1RD4LBxzfbvOY5xpcaCHVxck02+hfEBwyRLT2VNF
RK9TMKNnleUNQQorfaeNF5MbCpXT0bSse3KcVMk6oIpL57UdV7HehW2cN9Noda4Bj8Av3vfO5als
2mAAHj6sjb3kjfzjWdKdviyitTkyvxxYWml+oUqmVge1Tmyr5Hm3MFXGhuMxHDDIdDfsJOjNBZcL
2y9Q8L1AGWd95gdBZR2v0fPPt0nAYAC0pIKkQ+YBg7uxcrWaPZBt65SUOMH2ZjPbfUvAzVP9hlmD
E75V6Re5DhkSBFDrQXdYgC7gYQS6qhO9VdVUzoI44BPExJ2GdmN57T+ZqlUgW1x/fSbGrb/rUs5X
/+unVCY3NsIN9SNBlFuJyNN9rwzWK39u9TZJuMFhZzabMrVKu6uscOkbAbtjaMs8NOnNMC/Wsp2q
qzmmLX8qBns472FDaijMpra2Zul8VGCYW6eGXYxcJIJbqLkG39h0LhEjdGKOyGqGHmPdoxuoonbU
vu+gFGoZ7r6peeWhs7PVZq+sY4S94WW4y2I5ddeUIAygCjFsocyBzoOItJuTucd/C5pVoLRygr2Y
BJwdf1FMkwAE2RFP9Cfu4mqslDrSitYdj1ZH4nGWl5JyOrAeFxJffRIAjSYaIdX8ZTCiSBDsZ0b5
yhqaYal8hIbltYXFdamM6wmSnOC2vjWUvhcXhaOaHBG///fkezXTyMwjLFzIqpxMQm51H0m0VGyF
dazQSl7I4qyME8K7IXdJXDMX1nFOF/F6gP/+uYXtc/vcBQNu29NNdNmMaCkSCec0RxjPDgoZ3Gcr
NdmHaXfIZRrMquo3LsbJlXBE/hO+rQgKNB4g37pEz9GWftxmOJrAWteHZdZ+6FXZqw/GuEqrtjAA
MiFAD+51tqbEtyLvNodGHrFfcqDYqRicHLdTTctzBXthY1u+GplBvi7/qAAp9ab3Gl/mRTzIYwCp
Ce/zEzbmTaIdNs+WIXzLngvH5NYQ33njeHcPIwS7ny4XKflpoXAH7bTTN4Oun8TY8aYA3ODKzRGr
f+vLhWj5AKWBR9HatoKrj65cvGbe0c/t+SHkv5yUySC6h27S9dTQbywn7v/4TGKRm3zG7diHM0Sf
w7ZLIEmJGLvQEGn55uRJSR4/Xh5u9bPnyqGcXNGHJdb57f0Kouz5QP3fmmPkPSy5dngacNaSKgew
KSICiOvFc7h2KqaDSxgCah+ZsDavJdfI+qlcUR18npSAWftoNBGFH1dw/o73ICF6ftPlVgETVhwQ
fg07QnPhgJK3xI0WaE7hXvDPRxqiJFah0ijIAE3+VKgUqDduGb1qmoAgvYiElk+sZVO7IiNXA3Tf
+eyBn7BqXIJLE4FBVJfwSOCDhcCJ8nxPiNXT0eYc5/OnjEHg7xqMb2Y3kDmc8GmuhYUSxno87I1N
CIx1b05CnOXmcMuWU/A0Q3AJdt4X0yS0jZsI/IqaN3OnFzp2YJm1Q1jaoeK0kGmSFSibiC8ad/9I
WDP/eunGknqymLIrjjLetwogONEtnxNO24lrJ4+JvrqDJFYCLA8BlXZrjlVMlqAg1Qf5LQYSd4Fj
/4Hmf9S1kDTY1ksN18AtihxM0lEIaGAAIwhjURKEcLroTIBLETQOTRkXV2TWR+05/7JNTgRWjyiS
FL2WlGzd7uHLt9u89VUZT4g/0l+SxlZRv202TcqM3pubZLmu+e75tOTBz05hVlxxhOxYg+/C1fzW
hNu16QPZDYI+mSmOjrhOfv49l8ZioZuVZEuwWe20BZJXtdtKePvnXUDMA27ksRFtoi3vcCWbkCSP
cxTc5Me37l15Am5yeBIHPBETJ+fAkQW+feseg6o8+9i3f11fd4e1HmjnHBoKDh/Zv0M87zg5bzBG
umua/iqUt3AX+2ratal7tP3d0DDPYlZJSONrAfDQIMwyT73q9GmmRwJrg7oJB54K4H5CPincmoCy
xSFqLXY8Ebstw//B8LeA8oFUjfVbUoBG85WCWqCHShEb1tpZtRNINZwKmkEdSaw2e2parWOCKHOg
SkKosF+YtNWy2JVx/ALercyQ74inbQhP18UXTq5T8+da1Ud0egdIJc9/19XgJ9GQ26oVi+JDDV7t
LvFDuQRcp6afoI3A3vbxDRoDM1YrtDPk7n11YgGXYyP4/0Ozwl4Q2eIU6ot9o/9RHYJl4VnGeb4V
BS4oueyHtfzu/H3Rs16WikbqwhQKxlhZiXz6wZdh7M/fC7S+poYjUs/3X/aTTxlDlTQgpd38clgr
D403sms/6c9KNyK7jT4gPJCbsuPhgwHV058hNEMwHhtpY8Tk6e2db9DPrpPzw9SqV1gOSvvqDRTM
WzYxspWytex4QRgxDnv7KB9zDzxlc5KPh5zPEhMZZCy0t9lL00QATyaMR9HuOEsbA0soRGmvbXpq
lqETurMrPQgkJRL01HizNlWA9Ru8BdMkBDYeZ8o2hFgND1iKyuBY2YrU8gDjJahY5tT/77ODySYX
9d4U5r6F9lQbHWPnjd8qRBL5cA0dubU7ge/rORxAuO5IkO9gBwMAhwT/Y6yWHLkxO4XsQmujM0AW
xrQFDaR2TF5lbTkdgxjZLprqGolzd9WXRbUUtSFoIw6PqVAyLp/gtri7DXuqnOa2F5pZ9GUCsp+O
5WAB9uOgsQ7yn1UqyCxXw5NIPrKJJJhxX2YLaN6sX4lnkHDJLxDwMUfNv49ytFlu6mIMgYPqZMmr
ximQFK91Eqz3czCXabmcldii8B5sYYhIsHQBlLFgggC3MHqqBe2x61d1dO3QKeW6OkBn6UP9TI2u
Ff45KATq+qERbllf+OoP5Kzxp3eW10Fq6RHNhJuPdPdEDvtjdXWOPQhkN8arvG8eajTmYUtx6/Xa
cpD+88G5sb8bmO6i4zAxwNnHtHuIUaVlMyWU0wfwTPOXdc1B6adjRswy0vdE2O5Nc+OTj6VRy3Xq
8P3WyAvSSmOAscl7GvjmGm6hjajT6EylZzUowDwDQS46IbljOXhkgaIEYKxuiLT2eT3vEaZMMb5L
0QGUS/8cCOwKLDPANswlV/+kd4xN8ZIxuFV8hcsws6L9NtQUwHs0mLHo/OzOWW0xGaMrzkgHYEd5
xt/DZxjP4Q9P6ZCSi6CQz7cMlbnwTFVgfLF5INeXvBXgiHPjY45Ll2oq5+a9avq2iJgq7gaTc5m+
xI4OR++jY8hPj9UmvlyjPp9+RMfXt7a6pnxKrpjp1gyzGOwlovM9eQtYCndpscVQWRkk+iEcTGCR
AfwG2CAoQlqu4uw2fNMuuCdJTDfSnFrovO3tVTUfo1SKoIdw/QSjiE0PCj+cSVuaHkuWvfxFV4WB
PFQ2mpx/evuHww4gLbyUTlZD5EGQ6tuA19CBsQnABCddAQcj49p2HBK21LMsbqRGDmzkHkXs01CI
glClijFN+CGXbucAG+BOEYxVhuTWwZytH02KtFOXooqq8OWr8Ud6ngYofY9PZTO/kvgP/5Fitx1c
cSFiRbqd3jF9iWofppN7TmWQZyJnvplcpvPacbB146D3JyeLukJf9C1E/W2+ZvT8zOI+RI3UnMpX
GrRvkHfYwZ0EKReOiKXdyTvPk27sNYZA20CVOohLd9Bg0CaM5w9ZmyGn9a40N0wT9Ml3mfD/+YQt
Ena7Bsy68puPjJ445qRFIpauMsv59vZ9t8GynYZgnhXjjyPwb/9gqi+yTrpMGK0OmjK/q1EKpjaD
RsQyrpk7e2IX0/NWqq0Fqw/BF9KHXWQPwTtNU1psxvHeyKpKjd0HZV9ZalYEJ95zO4ya4W4PqKyF
VPdbqL6xpS2GMX4fGWTC4mF1/xDEa1OsufT8YbmEJqLmqnMSqN5ggMWMI5qnERh0h0eLaJGkYHp/
/Bbb+zGJKVcUOe5MV3J+h4mV3mfJ0gUs426KPUrFfBXWP0yNXyZoQtvNh2Ulp59i8+Pa71NYsnuE
UhR6ePe7QnFEBa5AAjRuhh1G5Qnu/+3Zcac/8O3MwEW0WtOok9QUe+oUalqFN+NOoOnT3iZ8YbDo
apHVKdX23lM8+RV7drgTz+MM40v85U+7BsxzvFr7To+hAhYZnYfh/tb2NHUvOsYQ1MhtyDyi6cmj
YBDoCyK1+apsR1cFdkNvqJ2W54EEUsIalEjSUjvuFFk4M6WE6QhhvdySrrd17lUsY+w4FOFQTY9j
oADdygR0BCsdJP4RRduNx82zr3wF6VFkzjzzBwyD67z/cmtzMu/mgFsd7E1Ou0qd371x5ULJ+dze
HxTppGvn8IMK5RuOJN965n2oSYiW2y76SNUt9RAM6ITvX40N/CCsyCFOmf4ELSq3/P9ffwtWDqit
oHCNcbhFdiTP9lcBIrmaP9h8BErmGxZbaUpjdDvc1DtrAPA8ltSQwYuXY+3Oth/EatXya5h0XTcA
5gO+aSP7qqXaDiQoejPYDj2QwJ3Ybst4SnFPrO32svzHWNKuTgKjei1iEktpR8NVDFzQ54Ncy0U2
UhC4hFIX1b5gRMOaO/kDVZtIs8ps1fIpyDZkV05Q0bzCLPSpk75sllKEyk55BzzTgzVRB5e1WEwC
uyaFqhd6VHzVb+VWMYP/S//8fkQt+N+JkZd4nPWecbwPCyuAORA8mwGuezfkE1QZHFqaeyqAALYg
W/2zEca8GVj2PKDZOCL2pFIZJg817luxnigjmuueUYvhliEjU3szFCKFlMp4wnxhtW6nsGcwkOOM
3OWl5Ri8cy9guIonoKb5Kn3D9yhcBN13695/Ne5wLMJBxgjFUwue8qDjg8rBfX3bbRaCTjkjsH6G
a/Z5dU/iJp5wCt1eoa+7nKxgHIIwjgy6Rj1buKA25V0t/mYJudAs+SHLRihoLACkgW7VqB75ouhZ
A1uQLLzyoKGd7N8nSpQeApCV78gBuD2Yw6zXi2KNoER1Kf5Dd1tuplA2PkMd8MEV1PxIRzPVrZ2T
y5mNGWmGJCyzKAJntbIIk+J/6mCLv9cjraaUBmFR/B82yRLAmxh8mXG/8Y1oQZYBt3gJr0RdhHa+
Z1jSBjIpjzs2vMfrv+TeGeAgkUDM7EGFr5+nhf0sPZ5Jg6m28PPGfwikECYQAXxD5OIatNOPe560
hPY10c3XJ6pE9eqxS8HPcLo6NkgYd1TEvzb26za8c3ANJ7KfoRJXxffLazsB5Jb35IDpETqBWMcS
/VeIOM1RmIsJYc2Pgap3UBWIeVElyswFoDwSnd69xsRdvaEZyNsulECrtV4CK1HE5DdwioaDE384
xWCGeOSeo75B2PNxUlQ600ed///YHv/QpJdAl+IXqqzjmHJE7poHWWCyZZOKDAhzGZv5QRF0rfv4
oZhtW4OfPrzMOMotBoyx6e53ejWFFT4rQ/FUZ11qOzbv/nFxBWx8UTLG/f5bkXgAJcV3ET346ocw
nc0bSJu/pc3Uyph+Wu58rI67/J54LmcQX0Dyf0YapJH97BMJIg9wu/WXxg7YqOlphBj1hCoq3IjV
SajTIR127aEzfa0DrnU5M/JnzXzjaZvZ74VYf007GOvtoSzMaKFpOCHe4bN7VSSS7exq0Fk2hESe
4shrLmkyZOrnhrU2bF61j1A70HoUTR0BUawqldXYB3EE5W3hF2TlIpg5XxBq3Z3ldpXcXJe5JG2W
vfNWbMR9QDncgn/0aH4aaXkjv6toghiHZdqwFKIWaXAnI1PiI6vJ3zuUZSNLr+Bx+o4QBi8r5GEB
I4sgLdRjdkyK93aoqwlXQBQmXUL8JFezbyjOw3RbkbwO1mR4Be+BCbCaYaqZcWQLV9Itl5AfGQcl
NosSPWLG4MX3u1eIIOXwi9vuMFXlZ9GcLXK9FxnXtCJQBS6WG8JRHUxCISd9ZsgIOXSgfG3DKCHW
FcnFUnWT3BPP6Y5bAHczO7Po7xDoJw/MwFJCEjPYYAVEIcO+5oZUqChnVcLCbBoXugcS4sS4bOio
p0MNtpVhRIrFnA/AHCxalhKVUfRQ2NGaQYOonoFmireUPQzkoIzKvVn7+vjTpFCIvtSH1fUo4nqB
/CMwUhTtuyUkloONA/unw8ofLe73TRJnue6z5t7AdmYB6BiN0tdeg/EHSPButyJ7X7IBZvFCM0Se
jejxYjQJg7lIOBYKcqcA0RhxoXw/e0dRZB/rfaW0eJiA220TAIniIQtN8H+yfP+GllkzvTepIIsI
nSrCVDN+qpo/NUKKjcKdXqgLMwbu0MAo3GmHPTGhdrlfpWJL9oYLVI9K8WirfV1NJainnnd76iu3
iC/86/7reNiGa09GjEc9Ln6sEG8Sd68beAeECBUgVrw6XPJNWuOxQdp3f3Srbw6zgIdfhfv3g1qa
a2eJREeFoaOaddyppw415F1YtO0HbEJDXH43S4YsfOkzurhnR0VIpdUDIP2JwEo03lLvyVpFFS9+
eDSbhfv4sINpsrYDtkpIR1DHPu5e2LHbqGjFfP3WpgYi1b8c+U3kEhaYCkvTeBYqtGMsz7B5Kb/l
ODtV6BDfrulmVUXnDBqQZo7YgokgFJ+EvPA4NqrqJ6TDxg9fEZrV1P8Z7Ow6PFCEvGKA0ysWApMo
DnJ08Kb8rUii7F2i9dbVtcgB/i9O4s03bNCFw2IGJcCWjaAnAZKrS7q2srRiRJoGUgFqanoFSu2v
z4eWPkeHBYCpnagHjj3FnC+lMukRiyaY9Ns0oTka4kCWDlr+I/8KC+/gO/MZ7OAg44zGX0/+jhcT
WDUI1+ypAYf17bF4EXMR7kjwKTbi12KJdTqR58Of6/kyw4vdAFbyRnkhtH4TtjaYe9PfiBfOF+jT
aknA52tfqRuQ+sVfdEvRItVhhlmIGUfNtMEE8N9VGyQk86j8HqV+95CT9CHKyUpT/LK5VLeDEn2/
sTDYbAT8+yN/0K57zegkworO8RG8EBGgWH/Vc+lHAums62bvJxI91ZtEuxTEEBnOM2tQAMO4FECP
pXnfZ+pCJ8QvL8D1Sw+ToOccgoEp3Cnfkrjmifm/R0ewxhNgiG/08xtBGHACP8Fh/xgcWAG56CIh
ST+b+NaCLBTb8tosIdqBOVkcjqUD18V9lgk5JNd5nD5DBxPevtqsB7bnpmL/p01eBb4ybGh2OscU
7pqxGr+UZVMB7YKf9XZD4s3Mn+Ar9XRbcC6E3qeigTfjwhLHiUEOuP2UsY87C7j4wjkul1ZV/aiX
fP7Al+J6Cd3NVLT9vmwvEdYPmyV+yGXDCWhc1iBWk1o9kgu/N/VboALzqggoLbvUZ/mMm/a1fv43
fwBijHhukZEeB+IGiRQAzrQvFYDimyqV7Vz/NiVu95rhi6BIEgqwX1qf0heJOu0zmN8MNWXylBBU
bN+OTBv3xzzXIcCFMFuN7afBI6K4cVLRhtOfFi7albjuT9IOrB547NmkFhG+yxLn/lQNwtePT3Yf
1+UZS3+6ec8a+mP2vMrp1g5HelX+5186h3PWCpfPceXZaKhNbOr6xsxdhEYdWY8nRK4VriyWHheS
GkiC1R8WV2X8xwtVcQfLH4+eOiC/QZF0QwAHxOtNr1O06yfATkCR0EHKzRnZXxj3E1n6lfoXazGq
Jw5mxc48WGfIAKlnfIjYqyz9lexy568CdRJwchNcMTEoHQG7YtYHvgcqocmzZslvgUj8yI1E45Ei
sTg2ZdUaYuFQsITD5I2BrP9pUvWLG8jUnb+/SzQpCsKfGWgRhuTIrhkqRMfbMdEe87rel9J+wZxG
mzeT9hezTX+K+5IG07FpsUZNCGBTbVOWTQRRqXIaPwkny9lbwJsk2Z637UoDqtFzl6aVHK0/imfg
wWSnGEOZzWYfoI0ZvXdoiYR8k0JMC/XSx4Vycjh0Xx+N7TCCHU3I6vRFCy0Ru6t0s2cUdGyi1i4q
FCuY8FWJBnlEQSHYNVPUswOCSgMH64N4WE8Ra+vvUpw0ZuGeBMeSOQSeULFcpAnb9QE6do4pTNFV
1cmM/qeyemTchpq//JTxsn6aQXpArsx04yKkK+p8SdKoQ+6kAmfrHrrgxLUh+u8CbYmrKykCP2yH
MTbWkjsmcRfpOG1RBD2R7QsgK6b9wPvW9jWHxz8I6WCOERINwOFAxKntEvu0LTETimweMJxnR9hR
0wL2iiaIzV8bzC4TT27QibELc0hCP6xMC274sT+460eIFqQIjGqV18hDjIwAkeJx4Z2+MHsNGesC
S9f2WRBIvOoAJUeBL+dCHv7ZyX6bNsINg+rR3k0efq02IHKHInqXGZhSdgQVueWrhRnw7tS/Y1V0
aW74CzmqiLPuf0Wc39ZwIaocw6xF3AUqYTTY81gD3ViUh05csxMlHOQwtLlU4UHBbzG7ruEeFryk
DhnOquoqJFacTnH17BEAlXNhQZeQGs/mqyQiZ2NFCuzebg3oIkRat02c9JYtIyn7zQuLubWvGVgH
9jO59fIY3q9T/WJGYpN71unqybjeB4eVFi44dGLlnkcwk8vPJv4ijIL1WPoXqxPAQ/3qUhmjmNUa
/dLioXCiKcWXHdBqW5SA5IoQkzCyDHilTcC1ky4245P1Fo/gcxrouXp6lCg2Jp8pUWLDAI+ExlYa
Y9OxlxXs0Vz+zCRmYksNRVh0M8iMm/VD0yT4XDz4ylNhGDXfSaG4z3A4tsP7zTMQGzE6otxM47tq
C0n+rkXJ6dHZH88UVQ8gm9YmVryoHfTX0Zdz1GCpFQJvKTPeC3pbEmPDKQPyWBuook+4+OOoYr10
3OblVPshOTbg3dDI3dVUQ4MpcIV8NvF9gpDH0MQFaxtPWkAAPOoABadeDCyMbOMQ23Sv6/dk76i2
tpLJ4tLU/R+2tvrqBVZUKhpvcoY7uO6dkkQHLYbPqV05zrsJEect9um3YRF13iIfZiEojfpPb6Ot
WNEIeQMkrB0jCOIWcD2YyJWj6EAZrR1Xziq3XX8SEVtPN23HVhbySBXXxDWM1bLdtysPTDwVW6JL
1Eky/fGTsqy8+ntuSeRDJTIsIC/wJQV2GRR2ZgVMq4yiBtrpTJNlnw/gZjvLxl4ji6fnQ+GUlLU7
WQ+N0Z+g7alNLdt0RmoPk3ivEQEWSk+HJVcGCF4xFkx8kNr8PPHC2lHg8J2HghbEBdjONXAKBhNX
2N1g1RjpQ3efTsSgsDf0nMoBSYk+LPon7BEIo+PrsggqIGi9hj5DzZd59u3hHQWRvDp/hu/zniQW
DCGme568vZbOi7z4GqJmq14b/+nr6UnsQlAXybLA3Vr/14OfDAoBhlmcd9nl02cZOJErBpTlou4n
HA1UdL5vRXjADic+ojMBhfSCuEOtK15FaMjLOjIUJ84Eas2/j5842X/0EjyEevE9fbzs133cwxRO
GvS/bkwHzYb/cyIZRPylxOiY9VBx2avkPfMEdrPoTPl99dGoObT0C97yeV16+eKSC3obitLi8Ki9
loToVw4O/g+eWW3gXzSI2RoYbaRit7AFg90jy5OgZmXDbw4QqRCvoIWWQ54P2WhP7OraNiMNhrfa
3jtEUL+MmKJb0M9WbfJahIy9a2Ha7+6wNCC96uyDpwO0p38DMces6JZMWRmmIx5dsHwWEJ0NGgkT
cIuJ76xT4avNyT16qtri8kX7arxEwEq8OL7TQtl+ymP1N3o9hnkRV6hyIsPLTNnjuuLxo0AWD6uT
BZ2bMWLTKNOOuGESrQYIyjHARgXom3HG4WFOjS9AKeeCGzpec6YGA9DlGUq0m+5nLrt1CYD2+mfB
BjT85uR4WuHdBC1KfkKyhWTJb3sgUtvltevWwm99sGFB5Au/QraE6iJ+4dPrrI8BL5hyKIiwfSR9
yHZwFwvKz+JGePd8tVrGIB7Kq7kHnpyARdfDIVqk5L4T4e2AEmlZ/xeqLlHdQQE9x9FosVSJ71MW
ctP08wMdAR7JU7u76xoTGQRXAmTlAbzax7nn0QLjiN/9SSR7hgvmgNLwU5AAI81YpFvb+kvSZ1bB
BCatBTAlNVzbS6qvkMwq74/UKjTSqrr2keOr5oXS63DD6J9Qa05hbPQxSH5T6E7INcly5Fv69cls
w2JMTL4CRy0K+ijYes+dIRH0XOUhWrh8M5fBLbhQuxkcEV/rZCyQgyVttV8585vN88dxCpWFcecb
fiE4MIVhZYX+Jb4jYIHkxz1BlMS1JC1Z4xrkkBNgwGsGj43BxTGAD9bMShQdETdubKm26kstxkEo
G7Jw3VLfPz3/Rs/y437+nWZF44sKxpETnEtHo4bHNTqn4kb4+z0w4qlsFdqXm3PiCiGXiZsgYS1/
6MjavNy9oZXyFQpjvOnyICszIp4r0D3mVKN6RM5yr8flYs4QN33MuqyE+HrEcSw1tSNzREItF5qC
VkqJA+1QSLAt651nBWWFajCf+5xSItOtBDnhGRT0PUrOm0bPVO6tJiCmArjjPHHugAM7bcyHdl/i
4ompHBx/NUI1jMrrrDeoO80hxRhwTGqntSRQqWZ67JufPFO4/IXvfgL/DNTlU2Lkqc8BYx0sjLwt
+MIYHkJFxdB854x03qHXBxwI50L+HFKOi6sRfQeAw9i4Q9HxTEKZl7E5jRjmf4BmIhvdWZSRYqr8
y70Tb2uj3iMssoOUcIFQlEkGt5NSXiaMrYilSaBlonYGmUpeOT+SU+GMe7zNri7yS1W6Ak6H1PG0
Cz5UTPmiPwAAnRu6XItjz2+lf8dmhKuyuuMODjsgqUcbToQWe+waIA/9Y0b6w81uRNggUaw6ujjO
2zVEHbQE4ZtW3WTXJdR9/xWbU5ClYYVWDy9+A0ob9ic5FxwboVOPZj8s8NoYPQDJAksteVpxNIpD
+obbC9NJ47jjstn8tb6c236XlzF2/ViawEUiU55XHBl3hR9gsnZ/kE2Y3ZJ1Absf4c/VcOvw6VKw
zr1O9/RcWMD//1x7gzqbBg06KwzClxl54BEAQrmFQwXkpsxcr70Gb0QLQwANNvVQcBji8pcwQyKH
dv+u3RIiO4r0RsxvSjSaa5DNbGeN7WZ+WkVjxNFd+MQpgoxGDz2FEpm0WR8gZGDtQkQCMbwGBJUO
iRAYjWszaRArwHtnj2lop1QzPvWuvtdG84hJdYx4DmPf2ZPJd7SslIupSNyEmnwsxIZhh5frcLWg
2iraxYH1dlugM2suDLrKc5TiHWOGpn/OWsZNknBM2QxzxBiSCImhcwCh1u2m1RrVsRYx03ZI0vkc
eqgBDM+YbVVKhrjT9ubcESpBhzr3nDgjgf9I++iPXJplTgsN9IIKOPtTQUpIVsBUOuTAnw2JpNLR
7DIQtl8UPc3eXh+nQZWnJdkexUkrSWgfi74rli70Zv+uDXuskplxNDrrF6SPcxS23XptPk+KLXly
/1kjCilKTtil5Nd0mfEeW85VGqCMA1xqecdN/7U02zQ4gVXf3bUm6F9/gzVu1Gr+z5d9yxTNQ9nD
du2BfHEdKgYj4SH3coWBoMTMj58ZEQZsjGl/b+lgrU80SkTL/qH7bAcLPnUV2xrQWFtlBiqPsk48
GstFba2kGdcU8v98SHBz3zJ9ufn4/vPzV17QVRfHIRqSrZIpF4pZVTiHG2/sEtRVHHkoVWAjMVB4
E7q5W3wX3Q28iJknDR/4RDfPz2WK/OVjdgfwB/bMpjjdDUun0I5WnZ3siuWBLr7oSPcdgKks6XpM
d+92AICSd5ZGGXzJzRap2n6GP5MCzMoHLRfeBn4QNW6Exjn9scyerjs5goksD6RRFDPbFWIT49T4
cpvpsVk7OPBOOHKxLbA/8n1Lyt6V5Jo/sgCpLH31llI2+RByOXikdks1t1oTx5V85v4DrwC0NpX/
VHVA9MOO2Gr9y0Rh+mA6qr3nvvbhhmf9RJqpoJ34JB9Fqkl6tkDCJrUaB0KwZ/kPP6g7l5JsP7Up
UoG3tTqCt0BE1KPiYIIe9V0t958F672lArUhNPlrP9/VWwEJJ37YR7rilreCB614u6F7KFVs+LfM
d7+kMXMt7JddLiTzi91aS0BeVMkLfrnpykgDwiPyZyFjawECCYk5AZ5K3/mwdEGiQxiAvmb1WnlC
Kaw2ar84wyYI3jDdaVCILFcBWr/RP0CrRWaMsnfX4UgigNH8H3TRTf1NgLZCrYIRFZF7UCZt/+CU
0BtJIAFewQIkJeEUuty5JatuH1Jr4oeDh+v7c6fG2ENHymp6EQPgaXOlKUOp1qtJXBTw/Rb7wRcY
MhmiqOVIH82BRK+h/9eyg586vgkbRzsNt8kMGZLZH7pHWuX083GffVhIEosqyLUcDjbrm67rbW42
tXOLzsoSGhp3Glms+5+HuRsbhln5hKxkt+1jeCmunn101n3FJx73CiROW4XVAXNbtkNIhlhyYL56
TfZhuJJaxcpOt6AubFafRlv76VXTAuiaZ9IDJO0XknQo7DY5r4dUSzFhbW3orjEpeePQP0KC8QdH
+UR0WGa0Pg/NBY26e9F4YM8qqd2y7/BpvWF5O4VC2N+rPGTo3KDwd61qGKzykemMc7uzuIOFLAP4
Enb7dBiElhR9R8C8jRuCxWcPK+F0Wmpx0lrkckhOd1iSYyIJlkVCR4yokX5R98yQ8ZmFQZF26KcK
lrpoUFaB/2gOEdJVVwk8zB5/WZgsluVhYT+SqKe19Xl4vtpvsiWGa5ktUVgiZlbm15ioQwWMINlf
HSBhfgesj91TYD6iImsUeNk07yFPcTQg6HXxKikVZSYnFTZ3WvhPy1EEO7b+ryFBPEy6S9zbXccN
TAP8Sevhmdg/1TslMYjbK/V7d/rVlgXCE4uJjcZzDqUdFQrV1BuDbBOlqjl1G9A8IB4AhSHVYEgF
OhJiQq0mnfj6sHGSDh3037OsU/P5XPZcHyyQG4jPkqGUqn53cudu577tgZAe3p4t5DJIEZiY9LW0
dmF++glN2RlOA99+jUe6GY9OlXROnr/xh2pLpUngshOoABrfP3kaZ7NsMaE0kuKSO5OqmJI+jMDe
QcaBc9kzlts6kxesGLRYZcTzQY58iEfmS++LxVNKM34WtPVlQpBlUkvdlR4D18kMpammSDNuH8ky
4ufPKXEYsOYAvVXB5KnrX/S3Ngn2es3FZNgUUUNpIZE4vzhfNrMitP5eDkkEorVdAqrhS2IUjpYX
Ow4Wo3kvel9eHUUHWU7ZoX9Zf3BGIPob5atFShWu1TGynab1LU9xYEqwnZvC0IinOx1Z8XA7IiWu
tgnWd+Yz9GyeR5aZbkEVuQ5dgLO+Fz9kC/U7pWbcGlggyV8csoT3b+lnHKHXP8AhGCRPuc43Gchx
G0YLR882lV0IP4jxR6x+qgb0pweE9jI3SBZMeY7D8B0bw99USBBOzmVfF9DAdZvTJnsOuHRe0NxS
49SbNjyibK/+hsYHrrKYutQ+fsYQHDdf7608ZBIcDGdHNuDyYJ3nd6vAEA5Sqer/ve+RMnKgJvJJ
pbp8QvC/YfzuFv3GQM7TqBbhnoFLH0a2ir88mJw8fpoQnLGRFwL6VLS1Ip2zpMEYnAzthVWMm3xk
Csvl52ub9mbfRo+09pFyP5Vzm8WcMDnDU08HCnGAJXzvdSsMy5//qiWpVDbA6Zgx9IUzEiiuE0TR
CsbZLnKqQ0wD/B4IgoaasvjN8Lg/bSoMT1UZ2ExIHL5Ck6PLHz/UrGZpk0gtNuTg+3tN9dce3k5b
tBWuCZbjywgSlouN3keJ6A1pK9C9mHmApeyimbIQgtEbcK72botTrlgRCfUh7pjDqucFS8hPAWdU
/F7blKbogSVi+26kz4ipdwyVWnr1JAsqUt67B1ekeHt7XrpOLc6jn9gdeF0WsKl7bGf3m+W4M+hW
hwgSPWh87KRykqQlCa18q+AVr8aBbLNDRc/MAN/hznXaEHlrfyGAngYjCiI/ujd0NiTJMQADiGg0
do5RAOFCA8YvTKj/c0zV4ol3ZVlkJDLuaTXUSsjP7mrusEgo47euMl68oa4ULfM1Eg5bTc4OniQp
RO+SQV3Z50Exi8ENULU0RtO/mZgCNeDr5fhxWe6cfVcQ+snQBQxX3AuBwkkPInFOI4A3hNSJp2QV
LnAS/vof8IDtZH42Tc22z6DoGWNQhjU/dK80xXYlSmSWbtsBYTpumX2puDFjlcL7b1NG78ummrki
lVFPfPuEPPHCh9TaTXkJ67EsPkOSlUCkihxB+OWqD+gbc9YEQSSwp2a2xzl8Ru0GgMB63hkfCXNT
hd3DRD1P+FPoVmU7mLwnLvf/4WX4sXeLD2nLl03HddTFTLcoLANmLF8mWdWUzcKPX55jA+KACc2s
ye9+W4RVY2rc50OY6NMCmcC+p3bOHqa9TC+LowlywB5RN6mIftC9YSlH0oQpxmTYdh8uLIKx5o7Q
geRoGkxibCyQli1piOkw06AgX6DPVJgtDiT+2Mgd0cpyXZRj6RF5uJqtBt4kZF3kU4p6Ugjn+Gkp
z9KF4+wdPNuiBJ7z3VHGSENb2Z8+cr37NjYsyP87eNX7zztfXf9PyW2oUyszTpCX27y8RQDUuWUF
LmCr11oRpFpZ+lh0OsbTO5AlEM9a+sTTDZgRwFHZrN8Hs9O6Ba7NwzId2iiM63eQGCi/xLh7wqA6
lUID+X9TG4u00/Kig1h3uL6u0nI8i3pBs9bCy95Rx3criU4sSOgndxeKJnYLTjim2NmZRp9Z/0t+
yLGz7oesCH/LJEdrkYPR0M6BVAFtRm0PcrmDWQtpueRcTt4UO57mDfOer8q8kK8vUNeeQvV1sGh5
8SVQddnR4MVd/mO2HOtAaNmbxz/YX1lfkMMGrDuZGaoUkM+dNdEBjduIeBCIJaBl8p8VAOwZlcEe
9pf3MTQw0nqcSxXx3EwI2FbFAwskZvi2u/05cj3vsmx9rYsgoR/qYttTZGeST5rA+NgxTIFzJERg
TRdynnbIlTlEqPQDFQr38XIu2EWUUw99xgLEScGd0eJaSWGS+F0Fbly4t6irx+uHlp8v63R2mWJj
6g3+iddEBcXi5IfUbMSghEmmclbq4o0TGfluibi2lvouSgNI6fF/Sq4sRY++3VQlzPwInR+gUcss
lYL99/ORtk37eWrSyEv+SR6cO1yCLNMrewsHH9cavKomPL4VMsLnRv0M6/WEogt/nakaDJGL9PyN
LXA5/cAJDegFt7cncceLdrh3/7g/SnsmjhwmslCKYhrPyVT/lJX7+5pyXcHNfOUCkZwWwHXwVOlD
bvQ/ygCN6dNZcscPpW6vtwjtpitfGqf3+4p7e1AVOZDB76YuFFObMCFTrgIIS8FLqhfQAl1FzBqk
AXJ7IWWAP/dISG/9p+CFgT5uw4gvdeN/0r3rPY/0+3aNR6043BczYieuM9aWG2SKvHwdWfnfoOGy
I8ZvW3DcNK10210lWJlb3zo3ZGwhfPRHDLau5m2sR0qH/6t8RU81zxXvUEvgbl5jK8KQKooWRDUV
dKezAaQwDl+rYk0+ftSDST8Nsxf8OHoTfCgwR+W4HMPiX3uPLomX/6GYNwQRh0KwZqA1pba9mwdi
Oy3gOGAmsW0364xKxjDUhmXLwLOtrV94wWOq+b+19+njT8yjUJg8t5AvKbxtX8JrixSnN5Hkj5aH
oN/qbjYKGX9R2/ztcEONiwJd08iP2u3l+GYan6YTBE3s9TVce0naeWYStuqLj+22IrIKryf4UKKI
jsoksP252dqFsUxtz94BkdF+e1/xFtf+0zkdVHc2FdudeuIF/xecW1EcwJdHSSB0Dlyq20PfaclB
toLoVGIFhoOSrLdzKJAH3SHsPWj7udmGnRZjIrj0MPV+nzZu2tK3bZDpNa51L6dEIOp1ermf0WN4
NUF4YJW4YrTeXAEIueuV8IOF2zKjZmVmban8bmTHeDUAJFsL3Prn1jex1RiBZ5Ev2HKEcQqrTqC6
apLrXg/oF0LqpjAsBSb26DFVj4wb169FIISFNprxNxjPToXam3/HgFOltVciyA1HIO2oz79h/Wau
3p7iT85uhe8RqxdwL4JDj+4ONrQee/1LTBzkwglGurAJAggy/TlVfruvrSwElqonVKN+2zpZbUEw
d7U+yfwqxQtNTL6Qwc2qW6HKL+ZxSGcDyyJ9HMvvEOrFy/vnQ7S2mYZVZdbOs67UUPAx58z/AYVH
tAyNVSHLE2N9Wg3RWW4K1T9ITOZyyRoc02F3Vwe2/nDS2gEFaTQdrXNshU+06EF6DhratMQocQBx
MYlk5XmJMYA7ANZRUVUl859Gm8aSPkColTpQqJq5cdfv4po7UT5dU4xvgk2U0yyKRYIhPI7hgJdP
sPKLpT3idRZqUw3PIzt/aAYkkuYiEXAF6ZrHlVG4M3FLQ/jHtsziQi23Az5dKHq6x9ZnUPlt5TVh
PVmuibWklyXJetPFEJzhMeFLDdNjgpmu8whY5DbS5sriCAoc1PzH95dJ3DwmX4T1MPf+H+pJTeHc
5nDHrY+diFe5w7uZ/q0cYEJ5WnPb+ZigycocgrrUYqgtsZU+WlXun+f3dbDMgNJE5k+AZ+ArjIv1
oScrusB6iXCsFIHqs1wdO14THL/UXssYr6ZjJaqY7/GEkjHRwZxTGTO/MJ9jCJ9hxGRE3ZIue7WG
F9Ky87F7gbhqjKQp8ku3FgB1IerZ5aObD579EIbgOdi9h/FCp4KIpH5DgGdEFbYm7wPe/pkcYsYg
umH420GuUT5u7xaH+gaIaQT9q7s3x4CtiSa7+T44FeurUc26mGuDsA0rYtL73a0lmMHWHN+NGflq
QVrYNMc8O4ulQpeSTiCtI5hWl1lkSLYvdgPLwgDJf9VIqbETDjZJowSRBh4bIDCwJRC8Fiv78I3c
c6ETHcAN07dp1Cgwo/UzOiB8wzaBXi1PP33PqYfxnIYq5ycua23FFKkC0BZ6sqyA+k8ASlhL5itt
AahHAi8O6Cv+4GmS996onOp4bYq/ZFQJNI1cboo+iPyeof/2tlXKrkN1EZ3str5VqalnqnnXkntu
DPhCkhwjWFVJ04/K0SF1pNCsEAkTzm5u7c6YxAvCChRdOJiqKdP2/Lpm+fWaS1JPdWow67i28tvS
/9yMtVbgpL+WwNK8nGadn5ClTfQJnagOQX6gewaowGuzwBakoGCyI0hYcgWW9LOM974KpXl6ikab
tasKgw+XXnEQpMVCnpgogdmVioV7Jv1m5xevd2McgBD+hMphQZ7YUK1pop87bnCAbNROQW25a9cv
QSGB5UZ5SmKQwV1lz5Oaw7r+frwomxjBVHc/4bOch8bbQj/PxvvRpi/7QXvOxRSVvXP2I8g/Lh3X
2pVXLjImLXuSKxK0GA79PWesBtPe7jt5NEdSIbYX0wdIw9ubbciNarTKlxmygLkeRTORqGE7fKGr
ET4ki3haBmhocXk0UjOBbEsDV7uDw1zs0RDymQBJ74YPWobcx7FSpp7OxL68a8v3fmT2/W6qul61
jNe1B+nXpsJDigAf1xKZvZaWr5SKrGB5PrjmBVZYbtPmidtqS0oY7dPywr8A93slmmP7s3OxKlq/
qlCgrHMJBNWvyo/WObKu6nSuYGQoUwyFW4qhZou4+1wc+OBKTN4i4hptsGD2L0s8ygzyG2qGCxbo
VT+36Nb/Q+2S+YBDKCVpxxPYMh0HWWrFkvKrSRGBzGRxrqUIHvN0crkQhg1s3wkfxwn/BAxKAlzL
q9Zm0GRrYmmKn/cbDCRrgV8+906TA7iTgHPSBrP5ROPKvZAjxpAS4vjOi3v+4aCkZFHACfTjfv7Z
O8Tkow5RvQWfr8w2miYMAGdRaUojTlFoSm5FpaTmOAal38u2TjHlMowqL/tNrR2M9zY0P1+DvPjH
k0NJLInzU7nYvjDBvjkbKHKX3SI+FUUr2ZR9PT4TWg6ehih6WZ3e5rVoxGkNx72FI1ny3t3BeSCZ
Z2ACAw3+O9wMoajDR5Wrz2YbTxMTpHB7oj1Xm4r2qt01jxQqse4hBp5GLQciC7o0pC3nP14ts/XV
VLR5tcctq1ay0D1xPa9ZQH6qVXAPIfKjdvszrN2DkjkXWaYD+6Sx3Exmg1CZ+5k6lg4tiEA3Y9Ug
/eBQ+9I8vxrIPrKlCVwPtSsfId5atseU7o/02vssV9m2b/CIgHQuI1YzvOQ221IDLIbKxQlwR5Wx
okVGPXo0s/zMeoy1WgvQkLYUelSDcjiVDfqth7cpW7eycQvT6deQVpO5BjhJWhdgarPkIKEFa7i2
BiKdAImpqBlbSqBIYbko2xpd996k2HWuh/TWBeBfFGwKd4lKxf8hnqLZrBcVMpN7KaDEeoH+c7aP
6B5xr/8lQ9QR3TN9nzULnufNn2O6t6phRxYBWHpfBcrHBXO8+qA3E0gyDsfZPg/XQL6FBq9J2bbG
caAJRgjm944LdpW5uIU2RNCsWD6UEvphx4RPhgB4R8C1URUpq1Gcb4lGuDmjNhKpqTKxsaDfyCzv
Pvn0Y2iZwV6cQCNILtIxwyJejJqJCA4RjFVIGh5ExZU4UHLlz/Xz+ZPYXHD/QS04mLW/T+eTBP1q
h1VxNKJNJ+eAUvipe24Rs3MGr8UOJkqnV8c/9XetTK4PGnOuWrxN6n+F7xpFm1vShowlW4BHNmXL
TYphzzIwi4oRgQXcfHV89D+W8upW5NMqE+WiiJsRnmxr8tIpDVNcKDNm5cRqdDb/9wiicG85OuwH
/B2oyB+FBzlxLC4FphPKMZFwb4SfYglPmY1y/KGS3vgC5tldgILzh6yAjB0+gHm3a2S6CwnRehOP
tcTr8RtGTzvwhdB7RlQ/vgF5uhAzUPobI6nudrGvbL5IgGCn0ac3waD0DyoVxBwUfT8cHZzqu77e
t8/RvXGxgGzsyWMZll23Xuk1PQcBI7BaZ9GBPUVlOaMwGO2C/JBfxSZTP/7Zi8q1KNz0BqF7dD0g
Mwfv7U6J4FbyjLJAoJnnzVcCHu4iY+l1kEcczHX0Kbl/28dHeAib3E5w7lLXHVG8peA7KEDbzuQD
LaFS0orRqF6d2UGKZyj4HW2Uq4HApTPKOjozPStnjUX+xyz4wxV3UOfT35llAgp51e4d4w2F2Iov
z+++bYQknpMzjOR2/jJF2MUEtWtmiw1NTVdRwwSiRjxepFsCaNLo2NIJH0aGEb+Qvl/k2eq/DTVM
2wa+Q2RuQBsxtkhIQ+A2URooe8+96tUQHi98lrNCaa8hFhZDX27lEbeZGTRQBH0R1WjTyxV9IJt4
RR21O+ELCzZ3glqTf4IMaTF9GzKmBhIqUkKFaKLxfCA5z8eW8ZzIGdpR88tOrLOCWRUJXtr/Hius
RSGjHtHo0bTOr4lQNtPoRIrEWZCsAd8sPCcP8B1Hd1cCQCar+r/NTJiowQjQQFckAeY3VFgW7NPU
FZOLFIfRUgob9gydGgYNLJPRCNGprQUgJm+1Nzb1mnuhN6X9NoLBjiyv/O+1h/pUoG7m8SAyADfN
2Exfz8k83Ruo7NElO/XFcvYFYZo7Ds1c945B8VD3YawdTfOlXkSlTxI2weK6n/XtK0fvOoHBXT5n
UyC2BSk1hrTg3Ydx6SAbuk2j473MHDMgKNMHlpIDYjix6AR9H/7fwsZf0TWEqIvVc1IuzRa0WFsJ
7ZSBTsQdBNfF0xWidAEzjBwS5O2loSxFH5LFdhCBWlzcT/W1hugHYzIrvaAB55KdklHY1dLQhlaa
oDwMx4p9l6f/wmKf4v0MXNkkZTXE6ZEi0WKS8p0J7WXxe50wpMTF2S+4OiQ/p5SSyfiF+HoMKOK4
eStCQ+zxYjXx5jLa26ReTK9nBKNJTJ1l2XMGtmZ1uklqUCj8QsZDc0NHHwrfjcq7yBTsCnuDayrl
LseCNkG1L9p8Jg+i73dQEMkq9fnEh/uk4MNLooD+emmfFQNQX4ybqc30PR5DOGaPUo1ywcKW9HNS
zIgfEu3zcGm0a8+EuaUqx1PPVwO+Y5YtgL5IFhcMEekLVzSM1MLFTuq7Hsr2Ev7m3pbLldwsDlHs
hO3fJXEHIbh1v+mIL0Mr86xjtF9s3RJUu9xhI0q+GDtY9r1Pesfezk+xrDbqvIEzqpYw6ICkKUAF
n13iqgu0/fehaG2WC7zXp4nj54VPYk4QY9mMt8E1J7b1OrSExFm2BZS0Kq9QzCiO38yl2qLA3/vU
RBhHsBDQ4ROBOradxR4PMstpfsstC7ZunN2ZkT2TV7cUgZDSSnxZk1v6ppA7oDwxDeTsoofQqbq0
Jn2EEA4LxmnKHbwpnVnlVHg0uexmQpHEzQJUJVghca/j+iD8L+5Oa4gKpvPKbQjVgcfNFZur0MAR
yp41vRsx8mkXDr3ZbwF+IrgipdfrPzTu7syHgIYw5p7OsmsGnhg9UDMCKwvbHpB/TKAmw1etTykb
FZruaR9Ge0BtVWQnTeXT8P4NTnQ1btxa9q8AZyI+LIgMLacltqrjPnf9PXqb0mvnWVBB9l/BZUst
yf2Ic7Ja8rd80drpLzbdiPWuvjek6pfUbLMeQ8wVNO1bT1xS/MRgx0KJHu3UswRa0+EOsTAo0wWM
/qihvDlugePEE9viCdoQ05DgsVrvmBb9nV/82iJfHxZkRkrbrqiG9T37Wtt9nUf6Osm6EfXnRJK2
HH+nRAtlryGKlHq1uHeixWylxj2CAuWkommSSvLaqjEFpcZgDDTmzYDnWQIvknQSHPVSobyNYpYV
3jqN09Em77WjJbRvrUfCpLK+tBqlX9B0U8CaJPrYW1udB1qtwalIi3OXTTwZ/nd/FSHP7G2L0dH4
m08iCBBtCtQl1ODTfaxJsoQTY4ZUUIczpoegUIqQnJ0qjObJTn4USFpc+FLDgw5kRn3zIuhsPrmT
dZJsPjMSakLEpy1xFwphw0XGBvi6JRsI3v/RZ1wMRr4DLYooDEC8i7JMQirQ/MaMIN7R77jv0coC
5jYgaCUtX2p7qRQnzOqZC0d7O/AULplsM2My3+wpJKhuNYfSa2CIpjeTs9y9I96237F3sQuJrjqW
SpSiflYA6uqHY0eOjESwIrvA875oGbHnmfA8rEO5VIK7k9fFC8Tlm3+EkXAgGhAq0/JJ16DE1HY9
ifAnAt1Owkp1MEK3kxap1K8iOjW0mjit+U56tJrkUddDRmdMOKbwMLBFPvvqc2y8D3pE6NHf9H4t
GLoVxcAAd+UunK5WwvKICeTdAe34cg5lYPuK1NBcVtivBcWXAu0tpvndhVLoKRSN+aQvKfnHzHx4
biCuTrlXNgYu0MqAatN0R0ISCsqBw1pd6uKr8usXYu9Kj7LYLqAYM8ztNsYPSVRP99v8eqjS27rH
QsKTtewKXO5/9og/8dmvH7PidzPLLTikPN/Gum2jHG9i6+XAIC7pBUkvjeQrZcGf5Cruy25gCZl3
6FmGBlebyAzRGDkpyLX+ZKxgZ9zsR0bUKaweZhKMmHUUGijrQRMkyv7BeH67CEN2Bs7Pb/pj+IjK
eZrZNF7tGZoCRXpwRL2yFbiLzqxUkgqV4WUuHgQ7YEtWTvQVQLjDZCnnrds8wzn5NCJrmbS4IO1X
SDBH+3kJXBaGlx25860eN9Nvz8S4+t8hyQMC26ZMiBYV7W70X4YtFzV3Yls1CfcytXBpwH2faFL2
Gvv9kD/pKKG6DLcjUL72bXNMvSg4Bp/YaJ1qJH/aJAHK7UrzdG8IhoE/C49UXZDtfJGwg2uJtfJx
vZIJgc0CVQn6/4TWN98KOW5cOLDXjwWdxKr5mKsZYq42UHcy32aFhoO6TtkuW1lKssNtSdgLIYCf
ws8d90m+lkWA2VFp6gfMLLeoxa1iHqQZjiC2BglU4wk9DnxQK7iF7IxkqLPjbN8/lMYJcMWqMJS7
98uVXWqTRCqaeg5rL37LMtBccAi2W93bjX10wg1YuovXbMFtFQ3UHZU9hjVIDeoPJrPps34nZYz+
GjMldQ1EGdKy3UAlyEjpYuFKtRyjweZW62jCacoP4mD1rP06ij7iJQ1pWSNlPiVj1iFlWqR01Zsf
ZdXru3ZfinDWZ6qKypwep/u3HzRsnZ9Q5NYXWPMcxdD+q2o5sFwO+7UrisgAUaKzkfzbnEigWjky
a7MiDeH9TYu+IPFgNqtSamP35GKhM/bs5eQ0FlfzHn1K6VvkKUJbAMBJWlGHWwl67Xt5QrwV77iu
4yvIgwjvcFQR7mEIdcTqFjpCnlbyhJgrshUAcV5tgEQryefQcUIrWE4xE8cp0uMYizKEezj3MkDI
tz5bNlHvnKYzwSbCLlGbT4UVDySNLzHjKNPvvTDyVp+3jGr8z6wYl98L6T1xBRlwghZ6Anrgn9XS
tBzrLMHQ3miCrtSGSs7uW5uknJIKHawvoSgkUoXfAW1vQG1LfiCYauAZLGPKcX6RU7/h/y653LAL
fAUA8dYgFo21WXYT9u4CO3YJWIuVgrL1584dc1HEdFs2i2BYXFkK8GQGcZAbz/CSJJCIn2a6pne8
0LXZWIEOrSZX1YESWOJB/ID1RhAO65RyxwZwSEkSnTPcbxF5B+7lzA3DkwyWD1hdrBN9bnASymqP
LP3O0RF8cvGJeu1n9Qm8Qj1tz5gkfXGbgwuCzDIx6qKV+cz2wrFEvuJdbnAeGsUTd26Jwb3JZzOm
GUd/uzrXbX+dMXj5hcCmAcrKxhVYfRq5jh3T85mUHfPz50wGok1CsnX1gMJBRpHFAuIPz0mFJmm7
dtGzGRaWjQ1JXPrjFt5wytrbjKVKJvCWOaJaw3TQYv7OwlTWXYpDS4j3mtiWBCaWmHWPKqE+exFy
YVGnxzSd07YY3bKY4Xxc+bhkTXCreq4/nlpvG7ouzQncBp9bUioabt4Pu8GCVfQazcnMLWKUxbkG
23M5a+02MA0u1fKV4Qgl2SEYxw1Ccr4zDx1+Fu/90aAg0jMJuzH+frabA5PweiVNdXQF7wyjvhn7
4W90R1lYUN0DOgAxKVnXawYs9Y9etPuZ4apxOmei2GrmY24ekDShomPIKQLr3kFF4q66Ht2rs/55
3uUuAskZ43JgHaFhHobKW6N7T9c5dIP7yIKMSZouecQbfwjpAyMdKejyNgUp0Kxzkcv4U2RYvLHb
EKP+/RFcmp66JXyoPYOJc7bpJ/gyS2jof8xwVQxA3GVR9EGhEy4WbvN7WCV/e77ZcIslbmn5NRX6
A10ghz9/OLkeDtmOKfQ17cEVhnMenvm+bWpnsamKSFYeg9Tj6drUM49Nda6QzErpnH3/zHeOlKs0
oiwlF6FrtN8s8Vh+V3dYdIVA0ebMf6EbQmYMfFA8a8DigoR8dQfJh7SUiHXARyRwqi7Jcy3TaMuy
wkJ+pZdGQHpWImMZ9Y187ShO+QpZHwD08JzPBIYsiGjloT6ZMv1PF4ZynbGlSNLQVpzl0pFE6XKf
cqyA33jZjSDV7KWZgzX0G68ztZ57esz26I1AIMVQFnSlPEFjzqCOXLoKOhM9JaNeQUG21eGdJnA7
Sm3l98DhPwdCnne1XGQOx+y1ekq14xjulAToyD4azKV0EP5k8vWDga+fDcVzDkl3iX191jqHlt+j
JZXL+OS95jZqBj2PZLcZP0uQXzb9KWmLKw8R37PQtaDyWxNxt4UB2U3g50WWg/1Fqn6HEKxGQcRr
bFzU28/3oNhvauh93I+tqjEpAOyvaSGgMA4im/5P9Ne44o1gfRFcar9Po7yFYMMLgeFq1XqjKJRr
/9OJZIZcat648i66EDT9BhUcZmTvIA7UaDMc2bIN/pnixUKCa3jvy8BEnuOUDr/46GhYjZoZaCI2
4PjJXOdGHNS2l3jqp6IVez1L/f8+0y3x3foIZ+iDgPQjSSs+3J8f4IMOix8tkugsH/bh3GwPoS28
Fryu2RpsOmCxP8bpDT2AXrQ5p2ptJdWCfgg9ADOcdRB67Wp6Jwauz4SLIGKOFyB/M4tMZ1ja3gtT
o1VJamxUWjtjYpQrnZEAREAkqEC33vT+rehfv2aVCeVjx7CvxkJmks5vzwfeRDUhEqfyWgGtthAm
znszv/2L0pZORjkv1kgp8Tik+IOI35GHHZ0P3k2iRZSnmz788u5S2B/OYE1PyFa9LSwuxCTklpwq
DzqRSQm/kWih5k3QAaxZb5rWAsoVrlAFBJD5UaoGOaNEJVK8BzONip3I9//zXDHe2fxHiW1SNI+x
m1VsnlT/fFlQQ0xYqDGPkPXGyda/rNioW5ot3PtODOydfldu/c4LcLYbln2i1GLlQKC0/cSM5BG1
UN/rv8+uDNIXwQsUBiXTUMnFDRh1jatiTKfZCTsEpPqSvsDQZaZt/vaHn8Zi4vSL/aJ+UAL/RQJT
ZNsDYF49eAjn/tapGipM7+C8WB+NoZZLSrvaGwCTaudTEJWPe/mZAD1SR/V6rmfXoEx9Y6qiK4+U
oGhXJLibGnIeN8OSWP4l89v8dabt2RFhsHer2n8C9XwNxfElOGXVoJ2TFURx/7Y0J0Vajj/IWseX
i2ZPplTAcMgI5qh49qVx5G+fJeVCldew4Cd+120o1YMDa/VyqHkPzKwZ9n3vctPY00bzOwFUCP0F
3o4ear/BpMuzVKagHK1owDC6jGVY/rY+I3PcFLK+hZSZqQpUfI4Gj+H++rZKj/cKnPuTqz+5RYYt
c4KJT0KVWxaVcVEWGPirh7V5NHOqJ41fFWSJarBzJrmh5IAxL5mN2LkfJT8g2mB0/Xw49zIx2K+D
ll9JpuvJgAwnnnIbIxN0pvHtPsysY0kO9GGWb611P64woFWEJtj14cF4YlSCCrKeFHo8yNiVIp4J
Wjir0tOK2PeNEHs1PHlz2yfXSkI2MjZllENyQ3Dc1VTWBmCSF8sd6u985f+8xZPQt3GdHUWgWN3Y
LB37yUwtNdCrf4Zltwf5D4PhfE9CMVhJndMgmFRXQ3wzLt1j0R06krKXY510kMMD2ESCwPcRFQnq
HfZJtXAKnOoH56AnQsUldMLPoizIP4UMdFJUUVwerqwJ9lUQIwvLorc5l0LrlGYZ/oMLbtG4+wKG
QKj/t3TRM3klCE9zNUiKLniXBhZnwFhlY/Fqzg/isPohd/bwt5aZrbtPgkm2EDaMbppEDCMeN2EZ
tcMEHIl4ei/kBjmtkHunTZGMS4PFc/r9akfaARP2BQ8v4J3OZuiwhbn9hFjjDgcRddhjmKMQ1thR
RX1PZ/BFPmoenPKCdoDU1KhlkMbd402+Pr2Du9AsKrrkquwQOkEXJ43LSDYPriu306yZM3DoZBLg
kn2uxKcW6LyHvXSPnMmrMoMAqwS11ufG2+Mm4coWFIw7W53KhibKhbjkGQLnQl09ugCXJkNsUk7K
0/TQYuYviJtB+Vc+fjTyqDIW7wnuE+qCUymM921L3zydo/lAilLY9HhOZylJsN1lqZzcH1/q3x1e
4AAww3Fx/ibuHVBIN6shBBnu6GCnSJdvHIYdI/q7EfbzCL+sqJmj4A05tqEaHpkbvpG4HpWnKo4r
AgFzGN2orVFqTL5RyCsKB3K2eSzsdY0d+pI5Qi3UtNaEcWYHm+i2bjJKmfKYFbEkYPg5PipIKMUV
UTJ4FkPUOQ3dYdxZapwREJ7PHNpKgWM7QVRuFvkmlWCIMcLPSXuwD8rHM2hLWLilea+sfynHd90C
/uQmSendIWu4vW/lcClGux0YnHaINleCfCYeKZC/GblC2IayY/sMzJvMt2oGwgmanKBZzstIrO9e
riKQzqK6VGxqKH+tMev1rhdwIZS4aSO5UragyWuVicq29GziOmFHw8A3UdP5TjmWj2dz+fJIKY7+
VSMQWjfP5UBIheQqa4aX9ke7b9vp95mC25jMYhszdAlD1fhm/UJE0Xs9JZasPmftGdYFF0QF9qIe
yXCuxErBx9CfTLyPO/dX7VJ0pKCpitAfzCMAwiaDwQcUHMXMHH6DjPa+O+3/OQ6fHYNSsRNoZbnI
ZWM3p/hWOIvQWK2Qj/crYcrBe+MYHR8iqraEZphId1a4LTr6ErPuBI1Qj3q7FBqk2gjl63SsFOy2
qywxtv3Wkoza6UbDoELfNTCunuAmjEMEkMA/xdahniksYOGFbHwHCHHjdJFE3m1wXfzV8DqehBqT
vvicoirKjpogpquTMqaOUtUZEemibvS5UghT6oJq8ikSLnd+1ebZb41ITgIVrm874jckcpwDD1xk
DRUNHuKPtJsj2sguCLri0Gt3k/6FkfUtQTSjbZt9lvsecMZypXb/tQgvZncrQI+jooCt6rVYhyxW
7T4kiOTRbhdDjS3m/z/yD2n78n/KCLZFP5foRiuUPcFsYAuHAbhXMp6stis707hUdF13U4qXRto4
OfPHSMKEa1nYyjtcn/7CHmF1p/OMHbv56mOUyUM2+NVjIZTn/MYaLOmdECA4EiYo8mqrCvcJ8NCZ
dsaH15vlIuG3btE54p4T03n5Ib3KTwrZBDN7Skb0zzEoIL4jxOAQsgcz4SF8MDu/JOFyeLj71pIS
/w202XPzjH/lFQ2J1Up7zQxgn37wgb2a6yIlLO1ksZuljNCR10cWppV+yTbzM/LejkdMLNmMcev/
4YEVuiUuOjsuDEAW7CZThUG6D2/DzreW4ra8NxiBqOciXbqhYmthhnJuPAos4YSiAwzSwMDxssSo
kczqcZazFoYhKM20jpDH19IA2/LPhx4FWT+xM+nTONhCGVD/gZ+5HPyv8KZXYWyxDm/12A2KXANI
ei3QxuCGZlxptbPuqillmDwTBJlOF0Z5r3D5fwgmnoGYJnB3PXHdAhpxtewHJvSGFv/G9mAY0XCr
tZ13pGDowi1ORMnrjNbHhMOld3z81+fyuftUyMusx+vfe3w28lO8y5Yd71KaQIbfkdvd6V3Xw2gA
Al6fEclef8LGfCk68Vs5qMADw7kj8dBgUwiA3Q9cpC68iD7PHX30syizaH4vNwJDlS0/I2Hh87FM
Y25P8O+8w/8Wdeu+JaRamwut4x3n7F23/Ibu4KU/XNDzq0klNg4WEt9AZ18eXfxiExNEoXXqJuFd
j2HEZgF9RVBcb2YA6sK3pOjN3ic6kDKkdQwarsPJ4xvrXV759FPn1kdw4kJjOLudvVE5plhn5k97
t/PQp6rrXaY8KSR7/8evQJoBZ3nemkv2VUapGefjsIoAmcULC3xxM8HsKQSvKKnz73ECuSEMT4er
jgmWLtLNiOzRW7ivsQ938RyoT4py6KVSKS2anwj+SNpB/XVWfvNnhok9AQq8S8jQ36WgN6ptH8DD
R87y9grTQAD91TxZDPetw9BD8q/ZU85tNGVhTT/9tLrkXcWo2pNIojjiqG4xRTLBaM4eNRi1Z2Mq
W+xkWMzQCbpUuqxf3YY39+AgNWhzdH3TMeojKmEGCZdZR4fsZ/wXISLLDKEyFQfbL9njkoSC0zA7
znrbU/DiDk4WY7zaIRu3gfncUZldwQ9gXrHUXsqzi79RXA+Vm/tCjN48VkLIjVqz0cHzRkjRxZmY
4Tl7oDE5XhmQgpWP8MshPoAMha+SGRaDzbaQlCabWuUL1OtIwadyuQb9XrlNdv0k6T3sLj1TblyM
HEsX61lHumpzqa1qZkEiyvtJkGjWIJ6xjQD1svwXQ1NfxDPX3/1WL7tRwpcFSxjkN4haT2By1yWZ
7KEhtuS1+kB/yW0rFBB2ci+5PNphq7d7fzro8ekssqwnpB0M8VvBWfZu1alEiwWSQPhl4cskkG6B
oXK+xDHf02whiOcHT23zYPjI50icNbvhLdACuvinI1u5d3f9wiCTZ8SRY2E/yBcL8umCFbG2PeQt
g372cf0DgEB5/nAZHwipJAaNHSzFA+pgzFycTiDABUZZnglqhayJxCDpzw6Y61GxZsmdMNdKqVAq
+AKR1uS7pEmjoiDxSl5dMS2uGUiiLdJHAi8fnFa5T20ceHUHXZHTGpbkwo+BH8LZNErn4mUUdD9w
HYxS4TGZ1w9sqkLxcNdUm83LuGoxKfg2DUp2SlAKIA1k8U6Mev3zv/j/NTpqwTzbG23OlH2w/EPJ
LeYbVA/B9LHVvQaMTdTULwmjAolVchYo4PG4PUMp2rDRwv6n1jFkRSV8trHFPJ61PFxHnX0rlkXm
AFN8pmy6SidMm23t2rWhLsFmGEFc+LSm4vixBxbfLn4MQv8CXOK1c8mPS3iX/ufeeYIDq+YSLDNV
s1KYV0wcA5qnkP7AwgEX2RzVu1imPAu4k9SBLMTVpYqQURRJn7wmAc8y7SaOAkzk2WK+s315X2S2
ej7VTdE3xa4S2VQDuGVutYEZIUgviNFBjUICzb8eDFN9gcyBhaHzpu5WZ2pQ5+QXj63Ct8ayEl2Q
pLcV2xEI4GWX5K+mTaLZ9a0ATlLu3z/5vtgKMi0X4WtRMpHn4H6ZQz/pMS8balbEIQiYj8hVlwsb
OK1Hm+SCcFHt+GxoEsBqqyQblLsz7Hmdh7oR6wZ9XtGuP2PbUJFtoZ9+LBZMLuwfMY+tsonlIC4V
sAKi7AhOexg/VDaodiLJCVcFX+cVmu2cfJ7yD2J0Z7MuP2BS9pLo5kQfhk0GjuzDjYKIVqb6tFkw
tluWXg2ozMZDOaQeMTM0hBM0sa3NrCrNlRZ6s9jWx+QzDgWl/68DiDxTN4uMiERRgLwwXE6osyIO
zqWGtrFl5qRZWab9xFE//3s9Fbr/f/bZs32x59G6UY2unOMCBC2tLn2iEZiLuxqriV6sOx2SEZ3N
kxIisz8tceoHm54daghTFPAUtCQfLr9xQxYxTft1vJRKKbpID+qkYrX5jn6YbZ+0Lbe2PlO+up1b
6fEtMNG6NrJr0RFGp5Yblj9R63T8YZGxhEctADluuj4snn9J5G851N3f2+bsHJK4cafL6wAKlj3p
35M5C8+yx4h8Zf2M6mwskQZV+gMsB0B5EDcliHBxgC0VaST4k/n1rjTtHThZW9bLGgd0/Hz57ecf
9zTMkrqPB1qsZmJtk5g6yAon5iHHzjb8ijtl99HK2hGiO1V4GTnjbinLS1zBLlfhzj8bVUnzRaGg
lRdBG6OLZltzIbrdZFu/AfelM5kk3CVYHl60jNlqoC5x4IWTfO96cyHxJXPgxT//TEOY/KA6jOHh
kI4Zt8sl/KoxLmQ/BZo0D+t9+A0ptyrWItebPQ4r9MrX5Dl7MhxZ/VmpaI+KZT6S2Xc24wsX8XDF
Mghl7uUOV7bG/1+AAxXPk14Lb6V0Bxief5a13tzl6YeDaxC2L2NkO3U31S5pyM6VVj7W5V+640q1
USYBZSNAnB8MHfl/JzfgpwMaGrLwPUJzW68gmcc1tsesbEOsMuv6Dwjfz7YBzwE7iN7eSKsQheYG
BNwVRmif7rQWDS8jesLlVXvce8SKQqNVZXYjyqy7/TtJmd3LKMpFqLvKg0VuT4PcKQE7XiJVxkL/
wXbHl9UD4kQ3n4//pfygreHz5Xdr+zTs+LkUsWbYs1SwY7ZBIh5sujP8JMSYTmWX9IEdsp4AQbDv
es7ffzPGuK2iN8YegxCOkhESn+Iyg9FGzT0WynJDNyfjUdp5yo4DBuHsJE4dlVCG3c25cFEGiP+T
sPrc8yp6JxlQfmzDaLcoCdB+HpXmWIsravCpe4kNTtFSs+TdpEL4bj0dstgRFjjF3rVdb47nSQu2
q0xFfCifgCx36zUv7rJc4W5Q38Nx35KAHv7HwqgjWUV+IgoNT3YnzBvtzVqw/NMqUHGVZH5HF7Rv
vVF0mKpS3yV5REnY05C2E1lXNMbRfKf/7gLP1BIh/NK92Zgd8GopYnYG5sBEj/gpIjI/0PvDR/1G
MmAXY+cy7Jy8kyM7xuY/vdVQ7gbIzjDfAOYQ9DldoIoGCnhFysan5cGkLrwraGYrC0cJYH77tVp9
4OuZ/FvLUW7cWm8GjvGysXsOTKOOTSS/sbN6SxEy6NboOURMLvbVYtgtT6JKW5VwC8JHMCehiGS7
eX9ry0YlJKxcz+hiwTt971ybIDwAThqQLGCJXNDZ1zb8mRV1I/vywghexAi2+DMRWrEX+5idsZ/b
kEkR5N2HNFvTwDY2s0C2PCPc/z6ao1iwBITU/lTJ8dxt+0kKrG8rbXo69wwT3sSNRZGRDN6t9HF5
2b3crW5P+CewJdxFvtIG8UPTm6IQWlhPNIyxA1RvrHoEAlEhsFB659akfpsuJKMWr5iRmE1jiZhg
V7aThg8CjJvnbh7GPi5CVLBUQupvsDHbMReApk8lb66oKJWWtkqR+AzXAFOM2Y24nYbYS/Ymc2cf
gQII/v9cyuxKJlqPjQk2AVQN+Ck0iuj1AqUkVtTIEuNvZTyfv29KfvFnAb4VjcWeWPxJLKcne+op
a3pDd8lCnx7k9N1LaTVcFVA8v1R+Na5Tqvux7MCi9WWr2k+IIi5uw6JfkNJNKaZy5tpIZMIs94v3
qDqu6ucNkuESAGjRqdNNs44OSzUN8j3fT2p2RRYEzxeBp/1Ew6PzvKF7qd8MWhD+0el8Z+28ds4f
iwcNt2F9Qxj9WQFoRfrni2CiysRFvqqf19pgsLCcUlVMgjT0V48aLHuuR5lyey+xI5YvPfKlOEo0
HddZ4otw7NHei6ayDHvXKnU8FfUEeIkhuoPX9PXrTAn5QsRgIO9WS2FZHa0ryYOxfPJgfd/xS0w3
EiiUI5bNctqLow7EgR+mJANZNvBJlyfXPbZDKXvACokS/q7EAoOPXppRcxg0rL0nX8mvOqmiFJAT
okEeXulTQTMUgIkOSqOMAJ8Q9maPPvSxFCxdic1LwplKV+wYGZ9YkrJC0mGqR0PGb+gvNMc56nXy
fenoTffSTty08Ige7MqvKyD8AaIn7VfrDoOJKSuaXrrFvQUg1J1NtkD/JP/GVglSznR3FJZ5P6Dq
RnZa0PUUijt5ee5b3YF2EywUbcBFpHbFnZkHxzB2wA/K1xEMaKm9IQBhQ277R0nRLCkjGsiE0EMM
Sg2u3hRNnNECnQ1XhVxSW2WHox5aTbBt4kHVaFk6TBk7t/sswdu6HyNSWfq/GzCy4t7FdHg03FiB
EGE+y3uiCf5XvwQHGniD0+8FD4RWXhSBhpYkdR2sWU6cV7Z0RcEgslv7SfaWT02QKVOdLafbv6VO
/m27A0fkOP8oZyDHLT5yQ/4bnh2i1viRjqPLRTcY6Gbvl4fMxbxkR1OulvVpLAAjn11VVY7qsvfD
ljlTViNqOtFQQsZLQycD5Grn6pOU+JQ3C0hqaIEGWaahwq7wLJWmFtfYcVoOeG7Ooer9kS8bBfjm
tofbNj7LmokuD2/dXTHR0HscGrxA+/crwtJqIxJBfX/HrHot5VskBq8TXeM0gBaqenslq/FpP2Jh
fIGG+W7pQO+UhFufPVKe47BV2l1nezKc4k7Jwdd0z530B6fdD3wLtfaKBJy8Urb5do/cKJ9ZcIFU
Erb1k8JjGBVM6S7P4fCRYp7IcYslob6KcoyOXRqFnXsL1xfsvzd19P7T9+aOyCu0SIcGUGWNFY6M
tb30BA3e5HnjQRmU7lDX6k+0Xdv3pipIX797erRgPlRYm/ktd8kNDzb0TCW0w6XVlXnuDOkZPFLw
KeXxSNxwn6fxh9PgLstdn16f+gq1mMueEtW8g/tSGgEZgMI7NlG5HqUtD8T88we4XY2SKcUTOcfQ
btSQk6YSXlE7oC6cyTPbqIbXVB2IfaXDpVd9dEmOQ1yN6zXZUDAEVepexlKnTJBhnoYMoo4A5KFd
jw6OvjZ9rL5GAIfxVMpEe0iAN/1ea8M9U1yPX+y58qqbCSiRsoljVR1HCQcgpI1jW5WsXf1AS0ul
AZknl/KMmt05UI8GM9bV7DWy7nxWUK8tmCzQO5BsVE6XA4ej7gCqFM4OdQUvQHR3i5oLmGFvrPJD
VhDfZu9xUSdUY9w8KmQu1FA7GKAJUM2Ye6TnRUpkwAoCGg9nMEUezHIvuElRWE6eM9HP0ZrB2tYq
tKGkFQwzENNDAvu1B9MHIPeg06UigUFAZamO+Sq4g2l6uYsPW3EH03uf566IBQkTDztbYh3RqBx7
SBoiUIv9WKkZN7prR9zwInojZjlwFy7DCdyh+ol1a3+h2rHNt0ZkrXXkr/1k+0+ha7jt79AUZNcq
o1pwYIDBvvnfGtFYGpxIbp6qFud4VSn5ePQz4NvtdwXMRSabcuoYJyPiP8FWP3aYG87GV1hTx683
ajuIyIENfdumQnwG/28rWx0DfSrorhiDja2Ske5Xp4VPWK89JaGnAVvK9hpUTucBPVtbPtgV/Qvt
BU8qfdMOjZcJ4U3KTUvNX0DjCLexgJOr/5UIWX6WA1Ir+Egt++AqZaoZedpVSww7yZXwkbFGut/w
xihoDqCKajxOUADmdjkakSS3lyZ2NP+K8Zix3j3TsJ9bLtuV1d1xnTHHgAFShsuaoElBI8hdlbw3
osVmb91seiVbp7fO5SYJTLerdxiLksS10rkUFm0bFM9mkRGCsJIir4MOELLUfdx5ASHQmoP75+fD
cuT4EVR3upNYfLqW3HkEkXoL43vi6YbYsv04pAs5HPGIbCqqRurpojICJcIuBYFV5DqJEnnyI8EP
zfybeDFf79TJuJCWh8gq79m557PFJA4qPm632RZuPwTTqLCJp9CRCLBfRH/uEsLeVcUB4IvZqN5m
vhE+JrWWaIFWdi17WVURz0YJz1wg2Cgt1jK7iYVtAacBLcRwvEXfw19rn58z5rWOQWovb3yfS7gw
kVWuQ5/Rzep4C339hKIWZj2xzFXtNEkXQ9EybC8t+seNH4UVcSN5Fc5Dfv/CSd7MeczemV7vsPzh
vIa6HhTzqEoE0iUih4803MVQoL2XyUKGsmxsPVsBNYYWTpfRzTFU974bpUiN4wNgV+MBI9nQGydM
lfNiwp91H4fs00xccqJ8BLGCW1krWGiNDvhcZ1RPkh6b95i2sjfHylncQ5ndD0wfrkCGlj5pD5cx
MyvG52lWCBvaoiGZq5kDI5rhab7G6EDR/OhsBM04YbxrNonN+zH3+5JA5ik5jQbeCky8OlMzYUCd
TMyy5lxU6uMSC6n7tn7FhNQBTrXX9wNjk8EEv8iy9QzhUwd31TLFQZOUSUSWQ+CTKpGPOdMhsLqt
mXH4j1caj07z6nvAwSPh2IkbZS+QZ2LSlxjoEn/lY4/q0SLuDDvtcVrlu04vg2sKHRd9xLmdbwp5
8C5s8tCXfwjC71gb+IvsiXFlXonS/n5zhrk638t0b8QPY+Um0zjZ+bT+EcYQHyzcp78nE+F7Mlst
mVrJM08omyGIe4FRZo5jQ2w0bstEhadvLT6mGc6uKLyRL3Ldu5uXgE+oEwjsIs4cXt2kPJdq8jry
i/xf+6mEWpY3pKtaBUl4jgwLJbxn++asd4Q4OuOcgt6xsDrKQjwuptmlJ/kpi4GS7C0XxcN8g0/2
Xd5RErp7UqchfBdV9r5hZzdhwGxXV4v6GdSOImXGHqeF2t1C+vxhSEGIN6m0t6x5gwVSzQlPxhmd
KaIWE1TPUggd94PIY+YmA2f8Vx0qLVNULI/YQxfls73eMx9jBYhQIuS9X0TB3F17om6gE619HEM6
kwztkllZDhjQaii3g7KdEbG353fmtbkS/CwBnkQL+AXbpRhe3QQDEZII86SmE39yUxCTbMmq3f85
PBOSx1CQ4LdS+eYvdTwIZ6zaps/WVgyHrbLhU7TWdI0DZ3WgqB9nhpzUoGNCeuEfldv9H5VJ5F/x
tFgwp8he7jN+l7f4wTE9UDlndW/vk6EK39D5rBKgxWzxHjmw2Gc3tteiRxzKGYLwjWfLYs3N1zDg
lm/t3cR6Hva4EkPQk59VjxYkYoqLRAwaxBFnMJoX6ieF5MRrBoe1VyXmWkHbh/VzBtTD3hdMfgbS
PZChT9x/6+R3hYwdVzEXKbUeCb787QK1t75x7mq0CPeHjVZpPSsD4Mn7/JLxmDDQ922+7yYYwxaC
VGQstXVXau3vAE1o3xAcL9BIPdb/XIzaGCX7rjPw0ui2MLmhv6cGWJ76zF6/ZFO5dmK1rf9cgTKf
pFNkJrBKBykg7eXd9xXv7wG+XDqKy3SRRIi50Cd8uKSb3Tb8lGLKWntWDlsEuz9fv8f1M/APhvCf
mI634f/Fxw1ArKNCs2IejHlYn++GNZhBPoNgCdagBFmR4C2Kbuo+g9hEFGYw68G7KGE/xewYQcjy
EYms+YSLEGbLBgk39f85/mosx/SDq0TY4etknt7k4cLem9mA15tgvu8+IKS8X7pRzhcX6XsSLfLk
KCVOtsaSD1iTn1j27u+vFWYsZAq7rkrm93HUIU3ZwSKN+YniviToxxOH9FpCDozWchQ3gk7eu8EW
9WdHlznHFbertya2JsN9rA62je2PUejdNFvezAVdXy872mnEN3sRkiORfs6ixKq5jQyJ2+OuaSa7
frdc23f0cK2dXtPAwP6vHM0jkm1CC/HGaVpK45P9wGPFgnmH1dKl+q/COWM9e5vaVP4G6HR43Zda
RwRA12q7wNIX0yBajwtemmzNPYB7TyfeXMhmY86iI3aaa2+4ZmsJfNxND53mQ7bvwE8SW3nxslOg
ZmM74PvDmep4ot4TcDuMAJEIVAfWY0RBTkAQbfx/A3n9sYafTwcHKcrRtwdJFQfT57UKTHHLdgGE
9vNZhbbNBNPY0DRCezw3NmQquX30vEcDVZwlow5bkI2aHP/6EZIzuM/QQpmArIy3+ljIvfBRNRua
hwmSpSA0w02F1rq6Fy9LY5aBH6JtZ/4yBrjolakiksm4Kx/qu3GOhWdRTMWOC22uSnk4QDH0gZtx
vl/joFPE4Uh1W4FMsdQ9c/kpMa1sV4mA7QkD44xSfoTTPx49KtRRAl2piC8CNiLBrVUit075J5j8
jTnhBEEh/sAU4ZCh1TO6cFX9l1X3gkKctKrJtzaRM5lqLFlCYBXJuyeSpkDdKdnmIkqDywQXoXtd
VbUo/Ud6Rih3LLmpfQpxiC88o2sBPRRTUAXjlUqAVRCchH3YWW5bfYCZTZFq4MNmGq0ZOQhTQtjS
EmLeMw0rjPC8zCbTzfMgkLpF3TbVAa0XWTHK+2+OetzWhFZPmoSFYX+ypF7mR2w1HscHQuoZ0wIv
saFKDL1tV1WXMlDb+B17+5bLoPcmVbVWwdf1ADaPuUPp0QybNAmgFqTbaBZ2NtdXTRKwdnFPLs5r
eNdNG5AWa4vOkaYcw1dUu27f0HOMgUV/nTzJ+wdZRXkIj9SwB3wJHY9nDG862EIryZWsI03eZNT4
StcEAi36MEgZOVxZ4Atxf10NpRBpv4eIzvJ1EDDfa6n7WG0/NsqAtYI9iG8+PRgpRx9VK6hS6uau
pPpRKDkpEF1/eiEkeHabplRcn3zu3d+k9s2V/c+OLRg5xjUEkTzx3kijKN8KyB8U1GY5qb38GaxM
oIboKzts1VpNHU8sEhzqhpp1r89SfXcwKwDTWN2d+5/6c7oPuTh4SKSEwnGn4CRwRT68H9BsvMiS
mqahKgek9jle1UoVQXHQqPWhE13tkd+dFfv6x483Y2Sf1C1kudXgCWGQfhOtgbexb9PoDUPs05mN
GC9kkLFm34J4eOISKgcL460tj1N0ouEyUXvismHSUlSEzC7hBSW0/TRW2wYolAtb1Ep5ESkecjvX
PksslW9bB8ZbzLwvyhVe6G4yEIh4iu8E7eP+l+/bJ50G62d6pECzUzRU+AarDLLMOlLPAXuWwapn
UtS1j5YXYvA8I0gHIHqEJhJa+DuasSnFjlr5w5nivlS7kfHB0ImnIIsnPy0qJVMnhgCDqd6OnM0Y
UwYQEvDcMRpJSQH9cVCFr3GWZjTD6z8YEwtVWDodH39LDc+Oj5gpsyjsvaGmKRny+nD+gaIOkfXs
eyHOWCScEilHQXtpLizhCIdgRqWG5+vHkPzCDWiE6/ox2pBIzZ29an3mbJ6ZPuszCvldlz4YnWed
kCZuZHXKvT9T3L/MhPVwGbEo5mnMtLeTjA4CnRuNfgPQh7yvuN9OIYWIjRBg1m44642etCGt7N9c
3WArhjb31brv2AH+sScADliNtJjA2d6Vin7Cr1uiyZfVxsQSVTzDE0C1LMparhSMxuexJeNlYZ6H
zhax/XKebPlLp5zJXTXC0yfZRGVIykyb5QRKfZ5TlWEvlIYFvt/iUOA07M+/mTJ/jMyACGtjQVjG
bTR7CaxZTB5GGs5ecl44XmDzooCHI8O7jf+uN61j39SluhPhcJGIOKHw2CFaIOwarUtokZTlHKPi
czX8Aez9declWyM2NBFwbsDsYYBnkr4jv8uNB7iSWLbybb3TUPJVN/QlfX3bC2WggsUM/MUvcMIL
B9UfRFdMarugpq5PnNfmNQ8QVL4TPtQWevY1/Iyax23b3QO2vvUeZQdKxbU+UZkfpXHmXY9fRWUG
V7WEIoF1ezdkkqBEiGcZnhySKnSW49oFq3Og2IkNwZ1tj6cyTPU4X6Yt0dwRTxdeszghejn6wExZ
k/7nFw1Q0HgKNhZ9aGACzmpEP+AT2Q6fimv68arV33Wpf8G314EzNbv//waS6CV00sNUPmEp/svw
H6ecWR7ivry/Tl3O48MoQdDi0AnEPcJT+QQjm5RzJgd4/LFGg35vKg+6xjlFYTx4p0gV9MKvxjyt
fGCDSAgWwyBcUbMkBMUXN750cTsyosVovJ8Exjt38uAKWS3PLOSZdmIoKcf91NenBNcHsLh2ZO6v
UFsvfolTys925gNR1oYDSVtzatvSzIozNGr3MF6lorh/1z7KOV2O+mNuR/n9TfA13zGXjZEakgEf
jzj58BhzdsslnFvKYMhnhDrc5sq5sya+1x+7GbQL4nf1WHQjcy9f1TTsjiLef/tG4eCgmXZZTeY/
eDDZEC5+WfyXAAf3zE9eozcc02rcESdvDpMblpW4j1jERLPRvq4i3i7Zw7LE93VJrzCEOE36/3Hp
ydce4XbRdJspDfEXm108ukTdiBr8x1F1oKtU4g+xnrSWCVGRLFvDjW1ZSGHrvzA+R0llSTnA1gl4
eyZwK7KRCnQw1slqHPQZq8d8Imp9u+b3hig3/x7WkuGK7cz7IiInDNzrVZyQ6WZOGmlRT5GQvsJ6
cAbOu+D38RW1RgUJwbxNwJaIHr3fjCBd0HF7M5bLz+ZadLzVWuqmDXNBksuLMrMtgRW0OQOBPXuQ
W2n3xox18n4Mzu2NdWS0qpBV4f2xJaB3sS5wfm/4zUIKfPwXf46yqv4n172SXDmGCRi8OJpZ+fgr
AQLl+/I9tb1xodky9DhyB2beZW7I6qaHeh0fry1B/zKiIbo36J4J+zZOB8tGY7PmvoNskanYri1+
3vqGWZ8jWkUpkYKU5naOnfDJu5KUNec3xpC8klSIX50yEIOCEOWva73JsjwI0/3D18/TGtbVQbhg
00zfrosuISGfHDFwOAWvjIINeHLu5wxbeCRYJailPZmPFZe8LSwIj9LM9n5RRmkp/RT2mlFZkt7V
DsTHa+wAfsF8TVRrOxahGEVSWBe8tmHLsybL6WbZ2axRP05eDDYaUjgIUpECllzxEgNRKkDPWza0
u0+wdDEzymNri/BcJa0HUeaAvBZQtuedXq84Mf+g/lqARwlpGrhQfMnKqFbI8ekQanm7SOqt8ZxJ
EhjKyw7nldBlu5I2eGt76y6Z146SrOtMo1W5mCriHf9DtOgm8Cl2YzSlCTsM+be9LiIKbqwRIoO1
uy2hoO2Rcabz8WAP5YqNwW1aXiSXFhBcKe/5D6my93H8NZWb4Phi/XPhOmzhnxR9RxdmKSnht+sV
Xczs6ksYZwF0YyG3XJ8pYLlw/KW0hG22lIE6whebwft5PiN7TaVS6Op0Jk8YTCBw3BUIHz3G87Zo
tvDMV/aZN3IWxHREID9Bf0PP/07qb1AE4jgjnei3ayNyEDuO0IRcdZroFmDcAuPrLr7XTk/s9O0f
tnjgqaQwX+IgeEWYLVPp9txVobdLw3g7Ek5HW2YmXyFKlj6rEBNkV3A1bGJu0qmwyKue+6WmX/4a
5mqUaChcUG4JfI8LTHJvIhJP7joF46y9ABzSvzTCkI5pOJNFy84a2NG03by++DSotKfcnfVI8TT1
zKDzAze8uU9Lrr41TxVmQC78NshSI02cPhdVhgmtWR1k4sW72v+208TQF5Pgib6k+lzrRtnAPDLq
Acnk+2mlWyYPPXfjxks0aBwGzsr2ZkOAPdmLK6+pVnHKQ12VnEr+FulqdppMAkU/tlSNZoHdFOxf
NQXsr4/KU4iV3RYKmQpDMpQxLcybaOLw7tv/n9P/LrbeyyHs4wPnEcRSNsWXBRLIFVpxiojjzQGq
cYOVI7BEM6AXA031/D1QgNEHG8/LJGkdgJ/W6KiUY/SAcay5ZjFTzkEF1XdXMSBWpYAiogdAU1Ra
gSb47UvwdPQt/derdtFvVmDBS+BQC8GF1KHLiGzBMAXk5+mmd33OB3R+Gt4L4WoVFL0Xjr/FYIKp
QArAfSX/1qXLH/R7YxFYcCDBHYBMzYFkNrkEg+ebimZNhYTQvBHbJKTBp75qqpHCSViM6dpayatt
opdHIW/6aaSzqeO7w2LWfswGzNt4eXYOzsyo4rphTAmuUg7hTWQZsTDBrzTGrywmgM2EkgPFKC13
2Nm1UELkq7k+6TP/fnIcP/Q5zkw/Hxl/wMUqpNu/zgamtVieqmc6jwfK+y0JywYB6do69sOmO8ov
e9tXKDUHBU/UAE8qi8smKiTHaxUO/P+vA7HkbzJtXDgKIMEXUgD8k2DypdzbeX3S4QZd/6P/nyRz
w0/xMDlpg3w2d1gM3kcQaQbKEt6WPsKTFeOh+vsY2nR6tAnOF+0QPeRZe9Od9oKlQj/lNFoKej2t
GLy+nPj4VegNB5g5Rdj7tjwEJ+XBA3vPcygzLgz2+KRiazTjD+HpeWAikrYPpe4RWQN5A3VZAUhP
4gvY9PJvowXNYGL43Ogfb5zb1vQGsH34M5lqscwr0C+DjJ2L8HycTyqcFwOg72vz0TmAUo81v2lb
8gR6XiidKbTcuWBvesAaPSf7JOmuBR7K/7Re7O2eZtZdtB+MAjL+zpbt1AqOJ9HiWpB5h6+B8Ex4
HicBZsJWumXdqs6iOFdMHoP7PoAL5dkhz9OyEs6m7dk39TpGg8v2XHGkn59vBj/XDzlTHN8iPP3a
hj9Ey2WiBPijG4RcQUmMIlo0gEMByvZWdFoktYe9MCnv0hSuIDP0jLb+ajYd4CcHTU/9nlu8qs/v
NsXmRZw+g49/WaGA5jkptSLvCVbMwiew5i9eWgLSNTa5ipI8VNg202U0yRWMkrY1H5MSi0GYc8bN
fKM2j9CXjaTqDsH8XRy7bpBE7mgx4WRdeH54HZ7T0rAPLDEDWRJGHsOwzCGXZyokzImCI/ArcWfT
6+ztS+dzXrZPhjlosYg9+G/5kbkl6hUaI7K8utMM5p/fILiFPL51ZQRKT1QvXoyr/2Z1ZQhTzKUJ
8iZ5XcXN6xhaG1HdRSDukGvTJyuIMceren3j1vtfEiGJrZgwdZSx3Y12gBCBCHXWxFIeVETAv456
l7sl29L0ZSa/O0rszqgbb7Lk1u8DlDnJlXZrN12Op/+g/9aS37F3IDS8blEx4Ve1YqGrFzP/2Jn3
UbqwmI5GNMpI8Ubakyf9KRUdNMQdTxpfglEPEAEWhfW359hlO+fns7O5YzdWw74Yw6j7nFLPUNcv
LB07WsheM7vqqT70Q99IfEOkGuyNTOW6XbONowHAzeMfHv104YMkPInYXN4gl0NBCDb28e7WprkV
XA9JFO3Tukj0Ivyn3O4ZCyY+UMlfXHw7SyhrDm5PilZlldM6x/KIBZWLwYImbmsyn43R9HOLEgD1
9CCYbpb6LPC6JupKsYfU9DMA9pC3vL2OECwmhcK04xptpkhS/x1OJf4GFNaKM57bVoCxkzL6nGP5
sp8WWO1S+qRB4vLfJ4K31UfKxXDws31jnXVopy2lzfiudtiFQ3McrevLMfn3c5km0SUTLifBsxba
cj5/4ihGAVSW/hX1y+om8aQznFdWgLWFv+Xgq2ee2elELE/Vdg1+42VE6TLTDrLVqknNjzt0q4mt
ICdv8XT7MExWajgH2OchbIEt7YGsV7W9iG9CTgObLs6d0rBQqKkZoniUsJDKE2wXf7hPvN8ZZHxJ
EAQxrzSvEJaBqtLsqy0oDe3fQj8fHmk0ylWVFAfpznzJidSfN3TpOgCtgQlLuatVwfs941ETKXuB
nrglIGzHabJ4E2Jm4U1/mt5XTKtpnmKRC40H/lPZsrRScj4mcltcFnU6sc8VmwG0lb2EnpmRgbSD
pE/qZLWliYt90u2V9v18eMti1o6jtbwd/8J3pmvRdweDEKa3QxJvZIVBly7T+so4UuATG36rsqg6
veritXrO+CuVGH3rSFe3404YVR4vjBjHg5eUr5b/j70IYBJi8PmlN1P4x0nKuAolgde6X2pUcIaY
pWKNTh12wn/InPNEn4kTh38i8Q+WYo04EBDsvKz3rCvAi2NS6GYYeH2PjDXe6QC9sirk8UhH9CQw
K8JTmhOxmfbDhHwJNY1wjRBn4fnWnjpFq6mBq4DxPlVzzvE926luRvi30On19PluzPe5SLA9tqGz
JUcY7jiF6sUtU3PTRUQKjj7kU3IJgUYKDLttLiTt7DAXKwwGeaor9ZNX7+aTueknmZj+gTkJuc4l
j6aYM+GW1bkgw+SKCF9DafOkCH7Zs1ums0JuBetV83VrzHH7CeUWhR0WvFuFrskqGWf4ajWObuIK
9LpwC91jz4+3f54SBbQ/+Cuo3tQXQJF09uR2w6eGl9ovY9W6pJLy1c7fK3utPIg959TGEYnWd+BJ
GO1D2M4pabC1DYbvJwf7yWm8c+eVBZ9qiMBab7kgJBRucmk08L++3KjQxOBVMtaJ4tL3NsbxXnB4
5U1Xs1tQMAhZznqm2LR6sN8Bm+2fkf1wTbz4I2Cxnhs0v0JJ6kHKrYbcQdOGB2ildikpL4KP04Y3
zIYDqnpI+HHEDaR5NgNN/X9oQCMnpzPwnDK44rcciHS/3tLDS7oj+JMbFi3JeNGQVi91ivs6yoKi
Scm/id30Q5pIHTJE9IBK4/qIVFcPwVGDs65t6I5M2k3f+VZXjkviYcgwa/C4y0LuFxxKfhSVVBMG
ZUDNh2InXIqZnrrQpA3OPEP8M67RVV/nkGVNsvc+rv77mphXnb/T/C8oEf0rEr9ziPH5TFf2f/e9
Q9cUG0nH4+yWLVrv9b9A7zrUX/AX+cPQaJeZJM1QWo39V+JxSX5lEWrMHftKJWXoNeMDyPjQAwuA
nqBUySXYQoIxPVZuNVa/fc0Kk/BDJs8mWnWIlxJRTSZw+CTVQG0wmaqpzC6buy0NWLBmEyKJ5z/9
Op0BbmMXy8ddGnuXGmdetD/Rr5bxGqUWJYzaK7Ub9Jgf4ZzpI8agx6Gs1JJllDu8ykqqg6aOlzD+
EeK1644RftwjoiCHABSTfSAUsMgOW2x7MGDMF3hWQwMvXhtD2TNjNMm3Ne9vp3eeZXApzHFkCaOr
OveJFNK6McEotaOsaI0Iix3hhdRUmTWB8NgkRy65vpLhjUAgBw+Kg9Gr80XKF+4ImockZcnDVHSl
qVDDBDMXdNuUbWo4p8qgYxePET210C5LYwkqTbdp5rQkmeAWK/svxltJgBwY5e+7q0x41KR9hc76
aYFsmNbI1/CUQ+xkGJwumyCw4HvRgmft7XedDoL/Zq4nXQXrODjI6oHB9aJ7eJMUZtTzCDP3XqqO
voPIIim1tpWYOGRVZNzi61SPoRZnEwUVlHOfOe1sxSLbYxgUHy82Po2dDfMqBkFXqZNbSt0XRtnr
Vup9laJicpBFlzG4K12hytv7IdmNlwtd0DpMXl2aDB/ZwocPjhIqRyDsBThf9HCLA+WxcEb8FSkm
sm+KCePQgqGjaAtlXkvQbkEQYJcpjLMYWEjSsBv8N2wbuEQOrcZJj6tUsJ88l24jEh/6Pb1yDVU4
A/8zrISqWdE8McdQOsnILjUg5rqNSXZcpYN9Jll/X87Df7FtWhDMi46vpABTZ7julzFLJLekt5iB
gM8GXfcpaF4ezxUYrYZh/QjzSVUCfzo97Zqpov2JhyaniR2G+MVGLkTY2SNYYRtpMaQR5wbuIf4e
GJFtMyWQsf+Az6fctFGR6//r3+1BJMfurTjHgQlUap7vYP6BJIUmtNiZwYCVaNIP2CSUIV9nvIKj
Vnhc7r6BAtx0Y1KgWwQF8iajzDSEqkUSqJ8r+BhqY4ztisjHfgaYRdsVnz1pitAgwMutvue1zwvy
+iZF3dDtYbQ9fQfxUgYwyIPFLAlgqH//3Sp6OrwYkbwEIMO9FfSF1uHppl9PJLozX6UahDasA0zj
e1WEdUEb9xZxN31WUde/w8uwuFdEEhcdCHM92VoHhBNwttcM9+oWnAKQ93x5R6QSq8RrSOnSldHZ
f97jzIPASwGlsJaNhF0RVy+AgKqhmynwl5KnAfXnvqomt3kHQBmzO2g8e023QjI2vG3Cz+6hdEMe
aa+bf8yUXN0uhG9aQQ3c8Z1VKBZl6Pia1/s8ebn4aNzzdT2gs9stV9Rd/V1SKdgPYf4x+2JicWZG
LYtBRrNgKcg1jgk3WJHv1SbETrxTpu77SYiH9NT4mkCtHTFQl2ilegQgydhHAZjd16odID9Zbpfj
qtNRe4St+01RF8F4cPymaxljiqSqVyQAoofgaO7zapxMKCBY4Xj4oTX3frxcEzJCfPulrO8YiD4R
asUIeqxB5H6cz8QF53z5OWh2/FlYyL+q9QeCgX408/4nHvzSmN/YcDzg4y//93mqauKI4Eb+ZNie
uarqXLqNyp5UXYQdHpwHBxzAC8MU+kNPTVylYEAbOWmWWW4Vn6lRDnvirJfYlrIiFNPQb8OwDArJ
fOqFWKD50UlYwh/ARkiPdoWlQFKfNNmffUKSm5s6Y7pAF0lF7x7sykHLM0Zy6udGiteKU2ARbCfK
gBAUzHBhVa+4Csxwn4NMCq76iP8Slr6GZwjfiFC0ReRwub19di1rWkEpLhBenQMAbavMBH/GFMCk
xkUJthV9hXh8mn2mRwZxWN/Fq0Xy5mwJJY1gRRLyO70aKq2LvGzVoC21McuBOBUDwtFtGXDL+sCk
PsckOIGIfdf+eQ7vKZ+XRW0+pph0Tj/W/m9GdSSD3PZsihbiqFvTIgmTo4jFTxAlYB0CQ4c7ui7w
FMcL/N2zCZl8JwHT2PML2wEwBLldlitvq3G5SkyYCE7fIB42rQ9nO9AATTU49GxG+xfYUInkKvDo
eJN7RxLw7a4UBqxSJDzTfDH+1j2L4dyiEJxC/BQSontXQ6VZUI8Y6XKsdP1NJ0poipNIeD7+VC9E
MjG0QG/CAqFUmNTh8eU6vGLc/+nqwxB5E0j621hS42Z6FQTs004IdIAvZo1PzoEEZv0i2boraSGY
CqQJOflAx02vmx4LGAa0XtKrX2IDuICqZAzSI+QKHLxb6kjObB33qgoKTONYz8fa7rNr6QlETZC6
CtpuRWc8wm4/Zs4hIQU/+N/SGhojwpy4zE/1sZEKphxx7XP6fKFmSXLK+cMiVcnzf8pd8A9qS4rQ
2ht6AhksiTN0U0KXG+pYHjLWv9rIileLCnCf1MpITnoD6ORMymm0cVqB33+WVqJXKjoI18GRIUsH
j4axd9Vpblc3OWSkjqHf0m45jQrEdy8rDMeNDYMi+D6/wsDlhQKyVdPmj00OCVcOGEoflXlplxfO
CJd1zrt7VLDKWjlcA4INIMEOXs9PPgwLQqTP0Zebk6J+rD6nywz1LMkKbOwRae24YogS+oft8Nhs
AXnKnKPgvBcro3JvkGuQglyaLxK4L5jDO0VPOlgUIM86snNg6gybZ9tH0Z3WEEtqu1p3ZosuvuI+
1BZusphJCi0c9LVWy9PyiqISBnphu/g3h4w/RtISnJ+tA1eexvi0BW+9YxJlT165NrNpsf2onRoB
zG1FL+tqYYjcntVX9aOugkGUx3SKL/PbRGOM5KlieffkfKkwPb6OxXKuhR2O8yMcHhitrg5yk2Og
FJQRdGmTkDos7oRfn0Uy86zJFNjjiYlBGYpZj2gJDndphHpOpwjkLLIfUkKGcZIve5Axts7cMANO
igsOpPoYYhxytAbEiqFq3ZbdS0Lj4qoOFTdE8mj1TztVDA/RlE8NSD4dE2uCLUO6zg9qzv/qnJn6
Te3m8R+TFCOEsIdEpk/7HaOR7BBetykmVldDeOi2q9hsfSHzybW9L6dvfJU0uvdQBZ5q++M+Z1MN
L+9PTGsE3pcg/uHouSkHvFQPnqk+FaXQUfcyOwQNvGggw1pd0pDzslRu9a+dWB47noDtAy0oOwMa
UWqgP3SJVEagaiJgrJ80EdkdWnN11BHEy84IwoYlxN9lic+CjQqvrFwYSWRKvspvAvAjemxY1iqU
DEGELegaWIGtj0xRoMC5vRquax3meidHrbCdL7xMzusk5rThmKyfLJnhoKlOQKiLG3YRt7y65XaP
6MiajUjbRwqGBSNt0THaW1MHgjSaH70tndOjZaovy79Q1+4yQ561Jt5XEPLQhiDFP8HMh+qwCs1T
hkiAWO6q4W3EesRjq7pcfhuZRofvARljWXgE5DscfJmXlE9Jw6PVo58GGOvu6QG21FcyUoCJV2c6
wN7pcyCSeKqmeIFVTqUB9Nu9L+b0qD/EiSvIEn/CnCZOBhWcomH4VdL1Wdf9Kt+Wihjl/Us5F31z
CZWVShcyWf01XtBKV+aqV7uJ03wQ2q3d46OImwWpkYdFhngAUw5gXbvUNhgh/Uz4AhY3MoJoxZXQ
s7U8F3S8AhKbg31gchwaar9BcEqOXZGRhrRirHudiTMY/sK3UBLO1duFLF3hNVFK8gn3SRaqNHuN
mZ+7zTMnjo/Lqwq3CLXCo9v1YVzy98g9ztUGtMY6Lv74ZsjsEbsAYr+lq5eQIhmTk7zMWMZKvZzL
LENZxWDYXNMlK8uOkBgKyR+Cpk+SOjAuotGbn2Wm2mPiGo6XEEAtAefpIg7X6cFlGYbVE2LbQdYH
CyqQDAW7+f9egrmQXh5A0WlJmBA/rQBKlhq/5MjXuBAG8AzVbp8fCwaWghSN4JMqF9vKcNFsW3fG
8IJdPeQnBoG63U60QUP+34ultwkhdPdSP9JHgkkOtHhJZDKJn9kWSha8TBg4XQn8h4vW1LeSd/A7
cz/lMMnEJR3B1B9Wq72WMBRDu6lGOGnkXZTU3NWAfx08k68OzmOLT4WWcK383ta6Ze5XQAu8oX1u
wBUdw1yOLVpIvWer059Q7HHSIgGugjcjR+5r9OydbE1k1bQ4W6OuXhGo5hhmBY2bdI7N7VehnATV
UVle95SMs8YSOi3iEsi9PRx8yAKBJfGtRLt/7w0p0lLHt3cKMNrFtz1qKfW+Gj9R2bMKKi6nlQUB
abmDVxD0nch8tNktI21jjUts/L8aMAoxoGBZyfxqx4Dcqkz0A3rBZ4pKxYgDG3vh+HGSL1laP4Og
HzI3Ce2QUa4KGG7KivskHcrAMVQzmGUU5gHGz6CwzPriTBfEkJ/Jk8tX+PU7hgNHE2xfoOu0BTrN
THcZ1UYBtjl59ZwDZOU4Mh6IyD7NnKCnIQycIBJJHmml8YIRsBBE9MQoA+d4a1fHUEIK0TrIqdcp
GRsCyNeYaCHyp8c5Jn0PUvistY9ooT2+obKU0bBoPBfJzHPn9KUH541Ay0JZjFI1/5t6H+qYKy9k
+SdRqba9ojP3PeAmxP40UCtDP7YChzyrBixsVMtbt2TpVb2ysb8josZPNEAsXgtzdumD7Z9DX5qk
AjpFWhsinaWB4heW7pg/eBV6AgwfR8J/aiTfoxB+0TpjFZnOFhba2Osp98BhcFIY0XJ5UquUYQq2
/Vg6f2aYXC/qX7dR4JlDvV9f2/jJel/CHqQAkhLUiD4YBo99HBUFLQ5LXSbHRvinrqAE2cNeu0vg
WDSSiZKRGhlL9+0pGbrGbY9iovaj/ktH3+71Yn3/wo2G3OFIPU93jG+uPGh/Vgg7CvHe1ycEtdZT
A9FPFhxFhi433DgF56Pn2nyVqdWEfNW3OIuRdlqitelmEaFwVYqbHFDRPKts3nbxqM2J25pyH8r6
B3D04MlR85c8FFbDPwH4ANPA/78as82ixUUfWd44wj5kqLSciwpG+idRIUkmF130OV+pokalc7M+
nDO3CsJqRcUxxwzehBwKpnutw+ZAKcUXepMQVcg4H1MtMQLcF784BkSmIP0v285KoT+b3ZwYkHEu
7hZxjHF/YupZOwJxCF6LmkAUU1RPtTR8AxVUlAxvLJDnlh4zImuH5Q8rw+5Cir11HK8KZugBBJHe
PZlzbtn1t2iGSDSzUyg9QWJFMBjgy0Q8fxWVDSn9J/ntbfCySi29GrAhXpAJ3ei+gWsMYTRaPDPa
Z/rOMYl4/KapuaaAt802PjNF1Fn52pRrDUTlbXudWMXrD9E7tQbEow/dQ9q9tXogjRV80+dYLZY4
kgd4XemEjLLjNUWJhuAur3wxU2G91oQkBeut2Vxj9mz4mMTJdERMr2ScRu1TBi27gweKTztpGVgC
Toy70oAbmlw0Ucay5TG/yyYghLJ66vI3VEVbpIYHUBHetKUyWlnsIYpjMBGWuKjnXuqyaMKW8q6F
vNp7PBn+T9sn29892NDqmyc5Q9U5GeK65HIW4hYLt+mZGyBsviF325Crp+EaaaN2smyF+Dz0o+Zz
sY+ARg7hfvb0ZvBVkt6+upokRFyH7Y58B8XNXsZFu7li0pSDOtT+WsdvB58Qtm71TBoR540x75hX
59w2W98o681YurW73xIls239ash777i2WnvWTFGB0dhpCgMYJ111V2no1BXHwJwqhPwgw3QhyO2h
1B+JffFwLKKh3HM0PgzQ9aJ3qsWF75AMuB/xEq1qwbCasy5UTwHt/htobwQSuP44F3Llftw+JT6H
XkATt+dRQPZ0Nz41ZrzaCX9ybVoQMS6mlL+CbFZZtY3le92jKUi/d7lH44AcAMXihkcq7C920wbG
igo+N9d2nr6RcrztGGfptSITC/iNfcP++m4LxFVpQZrR+/AgR+j7ZH4M2Lk/bZJYAcNbm2YHx1VP
y/wpE/9A8ieMfi7pjvo/27BzgdLmuJ09y/IuShyCoT/0zKihrikx8StAEKXBlcYPTYl1zVVFdwe5
hUv8xwjwY5cO++fPC5qLAfD3gYRmbrvB9JF3jnDcT1qUPTuvMJzMm8c0UFP7a+mAKHVhaa628E2q
Fdi75cnUIymq0RrEJedoPZIZzRE+GXOiN971Am6aFjL3Un7ag6kQ0EfjR5yqIbH9HlMSr4wtth6J
u0wOtf30s6etw1bn1AfKa6wMOzap8n0558uX+ExPX0RSSSNQn+TB3FvFujhSqleOjCJ0UyUbJxyt
8WHAqJVCV1ulL5jASupqW3G15Y3YBW/Tc9nTNpHJ5Wvd2LdMIIxgx11VKLO+7OI19eGSVzjnvZND
gxXYDdRSt/AKLi3TI+ZT4a9S2LkxfKq+NyTqUjj3Lwg+/RrPA5U9eTk3vFW07A8hX+Ttx7QTBSbf
UWCeRrCfOjsfx56LyNHhY3FQ9Yten8A4VwNu8RsEoikHZOQz2mNoxkXBzgQbexbOIjIjaRN727Lw
/YCa+F4H/QbiXIN3M4aWAFHLHYbgGKsN82BT0cXT6DzqlusxlwjFk2TVaYTfygpx/ZPlTqdkSu5o
oCSfMTaztdcDDb91vw+Kh08mwFG7Hk7kgU8f8cnQQU86ZSlb0q5qNhJb7hqEBch28xvgjcf2Zbim
D+iZujD4P/4aShXxpR8qaL3zQ76WWffipB4Oh/Zm/iF76/rw4DElhMcuquZODrFt8QEHNUdSdHV8
HWMM49hqRo9rCjDbHGGUWQVwybe4+UEZUzYPYeT1Uw94DMA3EtWQwEutagDptcxJVnGHf2vdKP/j
Ck7+NTr3fH4LcVJLydfvavNTU0yfDFa8jk0XhnqL+VHS6PbjXwIXkEzQ0vdeXvqw9jCt2lsXqh4N
yvHqMK30Pe7OVZt1jTjunf3LynO+KfmEmHFI4MlgPRA4/XUllzsWzSNr6IXDWRGxBQWtX5nA/Nuq
P53pP9MNG2rWr8RpRTMIXCkJXo6nMcI4zUaoLFextHuDLCYLRz+T9Tos4AfTbnHdIlCjmHtCo2cA
14OvIw1pm7SBea37grE79lGBmNgacxxa0QN2Mg35GqsXJYCR0Q+w6vMzan8ikCeZm5LZoI4ydtHS
yfqpmt8JPNgRMhNtPn+11kh4NCYgkxp74cAzcQxZDpGsTdNfsmQ03PP+Jn5Rtwa5QGD2jwNX9D2K
qnj1RjCcwgikvd1ipNZU7+ifCsI2DKXwckjR9wt/L0dLihJEfwTsyh6Hex81UEmoAPPLXVjofgj3
p0OF3ZTZcdilV5GAJ2MdHYng+12X+BHtS9K9Dw/cSN4J52mJ+bo90ddQw7uxN9Pb15Y9jUJ9Ma6i
v/3Eq++N7BxrBgyrKZCWsMVryJNd1t2iO55o6armwW7yfNbXCJKv9Ob1ygTwjever4aQXFkISUci
UuD928kwu+0ERF8ktyaphHpjyXBp4MIo2pvUttaz1vMrw+teQawQDTbwaZkr6HKyT3XX1EfSXiQ2
BkD+4QbPOpQVZ9ELBkQGkXNqN/1YzLCL8/svzIcJYiiHOL+LJhQdOm6VkXRbQ7rKA4ccZXEJ+Vx5
++8UjEWWhi1/kBgXdy8EFwheScOkKniApjFwwXhnAHQf9HGmHurlE2CHS4AbOZmjn5eciCkxX8sH
9ObTPmJKUSikEgkSXQEONw3WwG1Aw13++IEFn/LdMUEj44RW7PImYiOuBGYpSwFdL2ziIq9zgFMR
dqVZW/hErIkwh8SnwDjWysRJYy6xBKBzmomfCT95xKs8Ia+XA2CdakQ0GxAt5JzW9eXJciObtd3I
x+rFLcyv5jcgcPCnWS24Kay1yBnlz3Ja8Ia2Icb0pwlRT35c+SpXERwgEy8a0nmBwGkVFW1bYGgh
Qrh08IAvXG+xLqQL80Yb3+xdyto0P3pX8tTySRweTvhlWpPKbNEpHihSVNQsZwiBuw0ht5vh/+Ge
g41HywUs2TcQTwwfac3As7Np2+m7XGlQ0RL/fJZDBhl8OahWARjIFGlIfbsYijOHai+hJQVZJTpc
YI3QNx77XQxAo3dmVfFdur5g07f3SLFBoSvOX+9B2eRTYXvjHVUr6dFylXYUe+7AmNbwTxme/xes
yBn35I+UrjhSEJQLJd2nHmvvd/NRJlWUZ3mnhCuRN0wADb1aZlfRQBeqXiQQCMt/zoilUEzWGGTD
Aw0mDQt+IQ6CR2mtMTmgD24feZ01u2+PBmgxqU/rt6dVIC0BziUuTePZSxsCzuvkLXZMe5b3djYx
pdKacQpuWLTaOlBCM3EdGm4ZFx0CdVLG/P8k3L5yV82W6xUzVMF0Blb23j+Z6VexEsphbA2MZ++5
i66bZ7npYqBg7YvmgDxNz+Q5YEUPTHBVxyIJSdnHdW4HbosZl9JS2d1R07QfsdhxxnGco/7gSsmE
qe4H8wQg5Y75wNNQl/KpK+8A6FRp4qXMZd+PFyzwiA0tG+UBtCBUW+GcDpxsPegxM8UCK1jEuvDS
383/Ip0kgAD2wrYoQNILCyPCtebdI+qqzSz4RRDldgkazEi4K+18Nf61ZFdUj57mGekEJH9Ur7LU
yvLhV0k9BRbTBtx0vJ4/GO5RqSZnHFvxcZpNLnfO8sbxCjHfL9Zv2TFNqNYWhDlFs4Ubziv5x0pO
+qDHUAcpI6f1taevRrtsEmomjx3Z0FuRbPP84ziOujfGXR2cxjADoFyQCG1CHeFfbpP4L6m/KkHQ
i5AKQO9KqNh0aWcm2fOrzSferyw2dd1U+LGfveU/+vp38huxqt0RR3zSWaFTgMtaLqIc5y80NQo/
YNSCRasDnUIxo0GVDBvXiAKHoHiqZLXvaRnAjhC0S7e6tzncyFVDbF91+lPPKnCEAZVhOQmk+bI0
88uMLw34wUEAPIu8L2hR+BFYBuQlNvuRn3X7LH9+m9+26K1hdtZV4mYxcuVDpBtljHFeapB9b9G2
aA63tgu5yB+Nl5g4hgtaGyvVFVwSM81YazRSpIghG0KfOYMIQfQvtnoEZnndMSrXeB0FkVsPZI1F
mpxwTOugMvrR+oiay44PPR7u/IVD26eN7YC8cTHBC41eUb5nJ8zbOMYDahjKYjOl7TuUsP8HeDDW
pVFAawtJ7e332oG/w6axkPJZy39oB6XWZ2OdEPLoeVDo+SLXhsulMnq5hqMOdy+VYtiUmL7dGZaf
CmuXgNYGYUgUOrxDl3eTXjzMPfzHk567rvO92jX32XDeVDpd1G66amE9mQXdge4v1w85ruDgHbIM
mxiHgc7sHT+AVKJiXMQDXTG13Zb0a13QMLKJ0jceGHK6p25XbZ+5Kg8udhHQ67TcXhAlNACurH5C
RLMe9T8bK+cshVQ/fFc4o8iNg5R6mHnqOyTSz6S9Ue45bH1pnBPFEySDybYQS2Wr+NdZVw/QfUDB
9G9ENEpjDM46S9pCEcnoihzE6CsL4ZMdIrah0q2ABZnVHHrUlj2fs6PHoaq0oCgwCqcvoV9yv7FU
WH+4paybHECvuWqIqPllcvvO7okTwYs+I9+FM0GSG1yqpNShkCy/6K3bMeQhEEC9488wjQ3ngcjG
bkXLV0MacNzgOimUH9vZEiArnsgPV3ORwb5qAjqkw85rVOsmE8OSllc7j3oJE8NQLFL4dsWKOuzX
QqFTv3nJUdOJOPA8Hb3ZfLOEzSoqrDU2VjvXiN2tDMJLxgpPYVLAEXwfc87Z/unXjm3MTOvQ8cv2
cNA0NlClpUrlmF0YWZ+2bSRJEm58v8+tFTN4McWykznBVjclb1YnfsqW4LEiTqe4cm4Vw0ftYdVV
y2Ou0ZOKIWjqfGgfEXo66nq4SpbzedFugcCXFINjfcWkznrQOLJ9uC8iSHT868MN1yNMViXdnHon
Lo3BEjHRmq/kELLwTgqBdnWUl9HNmv6+kT+MIKHQYF1CuXqMAJ4dzslV504iql4hvZc+1n+IzSYM
4Qh/Em2WXvRfGzEh4AbEsIuimSuWBoSH86UEO40cdG8z3lpGXG6LvDQopTylpMIciPybFlnj/1pU
OpPRP+9YRgXhl03SBgik6BJ19NtqFFQczlHoWJ0BbCNmZ2885GHr2I7uxgqQ/6CdTVQeL3ThRSgz
wGCSl8g9lvNsDUoVnxv4HvRvVYrl91IaF23mAJHi1QzAZQOLt7HKypMSQ+vXdTSQHn1vuXVMJnKE
ZRafwzb51O0rnXYRHb1DHP4IZb3djN3XpdXtMYPdt+AykzAcsy31wwmghqLjpOPXRWMrlkhBs0pU
OQcFLzASLJTasUPrt7wjPE2wLDfnFrxrrY1+AU7NCMezsoYbpd+hl1UUXxXSZP3TNgR8t3VN9T+8
aKLXL0Go6zr5/ZF4+iJMhFHrUKQC1P2J7+Vy5ItV8knqD9mBTLoIFzuh+u/io1ODvSxv6SwJEkc1
h6R93TOaI1tdsWnvKN2lXaMCsw8Juce3vqTReTcCNMwcwb0uLp/+h8P5rIB8+d3zboMntIk0H1si
eqUSQ/9U+sygky5T78SFdLeSANnpwDYKGEUcznZ3TfZJz/WEzVKutIoUa7R/OKWn1po34uc6EPhm
5dsMxpxdYeFW4vGrpaR1JV5FqlAA/0o2ORGLK/CJs4lxeJnbT0qQLlruErsQnUcg/8+Tb/KmPEuM
3swtpy8c9DVzdP8JUcuMImY1t71IQwc9w8rVVQTfThUiH4inM1BJMu78vCn14yi+Gm7ojFcv5ZNA
nblb85qvby+6RkIHeMKbLsgpuX+8EowscmOoExX9/f/wsUJhfF5T2BHRiTmcJcz+2AuHYC+paC6T
ranLqQPr8REJS57DEV7+Dl18D+qJM9ldU3lMV8Mt2Kv4mt5HcqodN5E5OtQNT5xqIVnF32YRHetm
kLFprJ9pevDyk7oM+ihSd4J491OcoLKrfNMj9ue1Yz0lnp6KXE6A4pqi4rRLhHTyxqTp1VI5mGkx
RhiHAovZmp0qb9c76CwBLUfTIsEZKZE2rtVcr+bgt3PhrraBBeqVPWLmxPtupdUSJj1/KQSIRRID
GXs/u8PArV0L1PyNlhb7oKR9O3YRuArSDNGJNjzCOMOlkxafYa7fhKkbijcwOKku4cbTNF9ErxaB
SW5GuR2ousGyhTJkQxsNEUdXHsTWAuX9t1c204tg3+VJRXKjtzocRMI+uKysfxE/7zcrLCvznbBj
/opAtHJej1V9kGQNIfZ1mG/kkIH0Hf8I0OQ1tKmNW3LKscFSPYS7PlyhhJ77eWMwey/wrYL0VMCF
TCW7KQUKTV4Gnmka2EajmF8gj9eaInDagiQ+guzmWtOqeLKjIFhkCx1DOz/YPG5AOtvkyfgssec5
cIuwB7jO4/+EWbb6TdhAwi81NRdzJIwmFAG6WMYrfWJ8AQ/po/uz1fqEgLQQ3wcHY3K8/ZGnV1u5
mtMpOLj5GXPFlSIjbesoH/MtBI5sBABbDQJeJIr8CZ63vSQfNyc04UZC1CJ0eYTvtuMvTXpZfe48
jFX+c/Y1y8JdcxF720DyKEUgM4bi6txrlBmW1dv2gl+9erOxGUy/T3z5cImaWAVXVgt+x61238AE
bVKSfFRoei9xtlMf3gyZeHbhyDYAVMkZ9nuZth/RgHO8Lkd/GnGF/LUKacYQOkhkiEyogF5Ak0DU
BeaRvDcFyTg8XzsIe+tuAHV5Un/BfwWJq3wMyGVtMu7Ad7JPtDBwJtkehurKssQVdFlSG5QEYWuV
bNNTmvlG8qGvX+bLqu9qu8+5PlWA9RQCYBZI3e+nJ04eQ3IV29bKlrNAP0eLve3JpabMpbBelsAU
Y+LhiFjfAxVjr46atPK5jeLw1QkY8MBWCjnoOtR0Fj9c3BuGuLRqDCQ9mmKE7RWsltuWuXzptppO
AnWowAPqyV3whW+kvwx/n5agpiCr2Vl3xwCYcwrqXjunwLS6zpX8XJqvBiCviJsi9FwMYIypcLlZ
7AlwjGDj/Xnp4yabcUpZVHns3+/HIoIiyUdxNAyGa4mPArGe80Ay3C3t11oM1+wzO7mkFZku1e8t
oRvKD4kvWzEOhE6h7eHNLbrC3xag3vtY6WhRNBtjcqirn8mcObKrzwrEiManTDT3CE3phC4uVRhS
0FITzo49+XiejG+QcoWzC05VAsn5UEpf4Jv1rnSPD0Yn9gdtGD9IU5sVtXGu+pdio3OXEEdWLLpb
ER62612YfrhWEb+DcmIYdu+LmISOrY+T3FU2v/uNWysYowt9LTRI06uRajYBfBwjBNwD4vSOUuE/
m2XJuVfIRzqZDdY3/WxNlkJl9pXEoklLFKQ7HgLWX73aiuV7cs/idpfiHy76VfPF4Mfh7PGhCJbI
G+BmsqHvW9BWH4H813uQddGPFLXNaAe+WDgoAXAXXatQnO0pbCalzjlRL+YWyo6Baojfzq5iXJ8p
41qkIdLKJbD7sJ2ynrozCnJViqE9PFWyZ8iK8nA4XD/RAVpCJGiM3bijM7U875bc0yNr6YV0gHhU
cnh4zpYVzm0akVPVwNnxXshYvBOWY+5gJpyPU2I6GltnD8unp1csNVSufotQJEMMfwUlFwleyVTT
ERWjDUAElngXXlKoXgKD4h3znw0zjzfjlIfxL60jZpk4KWIXvhJeb+8MFdi1/LAMinthNCdYIp1s
P3mXbm4iWcf1eIry+h2OmlF/oK11Skosu1xYRILRFbnh9OF981gnQuB65y3qz9C2GJjUxjCW4Pfq
RJXKO2cuc9UNA5rMmW1T8F7vdvN575Y2xQN/wV+ghePn+cvxpnxNrRzHhBkfUFnLInWPMlrpDsxJ
QmPc4yUaIKSA8sOe7OAU16oURsdH2rUKa17BpbnGZOFKSfrQQHmUpVGbuspZzyjIHQLfxm9kd+7s
GIrkHXgiWZTacEpHNyoHFl9oRZFdcf9hJXOwtIHziNtuQr6vhVoYsUiLwMFrEPfjPmcgF6WrHxhB
tVRuyRpop+01DV8YPunF8yYdZHE9/bErytXaQTVdpQAC9JLsV+1luyim5v/YIouBTdhxWc+6JULv
c+HVfhsHWvrFnL9XCE7ExDY+E1Y3d9WPlj4MJ4ln/RFdR3JnQShmUNRAvbwO9Ii/J/M/m9WDcjMU
9youhSlU0n3G2Xc+cEweqDJ2EfnvK3PXp+SwOzF9dsEDuhqxuTjErN25tKd/499MPgOYaHGr47Xj
lQehX/qtxIkPMeES5M2JZzcs2UU/vzZzeWam/1V8yn/CdqkjM/N6RAlKiSO31rezyDcvavMXKEGs
cMY3FDJK7aG2peTC6EJfQZ1E/6/1RihYRIiuSz2kK1NjzNcU6ekoRg6wwZ4Rv8zSMCfRXS9jMaxT
xxeZxqYMO4doqIrPh9wVyGRDtY7guthreAa7Xtt2og7as9OgrXz8luQJuBegOpSmIgCAL2QXfVTi
XXR+g6rjdBrTEI7doQ7bA7kdGa3SdUaZdm+ZyJ069LcPw2XTDR4PGwf7i2PmpZp0Y6p63kVLUQO4
bu/1CTGDCOJOZ+PZzRCEXXVA26YmiIA2FvcxeKyGprsyLLqy8qQlwaoQeMEFysh/z/Q1tbvaXKnD
NSg9VEQnXr9ZBag6I3uINiFkLs5kXW3Sq/1zYSHlRsvzl4K1gdVmJMSr8A9wXulFU5yqCxtAOBAd
Ljr5thxzUtNX7UEKvEL2TaTaZgeMQHr+AAWcjyz2oyOLwY7y2vLQIhxLoMn2Q8VzybNaqzRdbEAu
ch0gR7G4Dm8St2BjuupB2+hJOEIo/yQRekOFwCFVnGI9SlP7aamQ3DG2Ut8lfynNRju/7ZF1a5Nw
UlIcdcAJB5CrndUDCdvqDMY3Pxc21c3iXkLQ7whHFcqdGLKKr4vVG1mpeTVDmSDVETaKMfXsQc46
WffXQ6z13fIayckh4lOTifZmHnRUr5/rdANfvCXGmAW7DD5Fsy51piSnKWZmIKCU9+y2BhANfU8S
gmsCcI3gR92WI3ygRkWvT05IJGrQ94vh33aWo3ezC4VdfW6vq5S/ndAgejHtVTEFkz1ID0JdKdpa
uhnlV28Pihbysf1xBAznYIwn0hTq0V++Uj5sz4MlLXzqDmX1gJqo+o7u8/5o3B0SvG3gX7N5pLwd
qDU3NK4Z0/7tML1dCdhdHUC2e2tKmPbeO+Jxn+Wed8o21hmZOAiUBMxhAioKDkDWV4hOsvcJ4QPt
MFW5FqU9XgMBFGbC8Brd76xwbF04cM+UePjxjw/J7QNphEQLDbylweUn0HNk50cb1pxGdrfKQxnW
5UyRmYONnnjjG7K7lmgHMUfIH69OovIaEVuJA8y9RAZ2yMA1YXedlqlmEc1Fl0HAXf8FZbTHCQpf
IvB1sGX3o1U00o9iATs4BORNgVLlZS2Oy0FhNn6sFNnaZ8m/EZJ0mpHAxK5bx6KJg3WgROnbK37J
AdS3JIW3Dot3s8D3UxLB33F6n7gBT/QXtC3dsfpjxPIOM0V5+zLLO9Q4OyaIoSzpE3eC3LMEcq+O
tOjIbEWZZLtbJBfoLupVUp8Deai4HemrtMaZ5vxFOfg1xEX/sHfneCn+ERWtJmG8NR1BIafAL3Aa
/8kNpxgPhbZINP/JZhxPoDBlUzn8FXPfLS/FF2nTWsHCX/W0muLic776EsGvgtQY8XMmVYupw0vM
qv+KtBhDybJ1kU0R6xMuk4JsoXNJe+fD4LZoMR2b6bU/5Ps7OLpppQ7kGeSmVouiz1fEkzdLENtm
IZX0my6tR/3lJ8mW9CeTkw60mLXEh35W70md5eLZ8K3hyppoIi/KjA5aGefXHEwJGf0YkP51ssWR
kT6zhPcSoriYhToGYKmxCjyByIMPsKLalCJnkShyqZVN8AKGUc95UtuJIY3m+LkHW29wMAdW+4gl
+yHKdhpjFoL1S+EdtBoSqCYQuFTif6UrOXYCMm18gRUfmdgo6w52RwqKMVGU9KeMRjYDXyuDiFBh
HHl/2o0NQ2+2yY+XpcNsMB3KrvKEv2QFle0maoFfLypUK0wdYEbFtnimBDEai8SRAhL2MtN2R9RZ
KDw3s5idb+BPQE3YG7eRdmrpbfZpIeax7l1IfGYuZ77SnO5dE3K80aG7wTSXLohzxijxc0JE/2FN
n+SISKyU8MECgzbIzyYfnm83OoP8MY1QO/k75MQEPhC5BJsjI4+bCpoGq1q8ba030B6pW2XQpuYq
B+E5x8Y28hRV012bcxr7iDOlvOm/QaFUN+639/lTG638WFRPyYh7bTc4aGszJG0oHMPtG3tGoSd0
2hLjCIqOq9vR6R1ByHqMZNb0aUSL2OoSt6CYNINmdKF6mP4xyg6XbhQaHveJKKSBQAPAw33PVPS9
56EfUqQdFRj2TvYq3mXYOmoZEDzeUbAiMYyeqDvqi7MUh8KYn7cV4oUl8xrY0w9EhHn1otQnbwkh
63rHDP7JHBIRXnCN1B3r8UVa1qw7sl6ZfOY8N5a9DjZ3hqa7dbanJhbLV3GrRrEBlfZXEN2EQg48
MuvFhkElv3JGxByRfy/2wMOeaf7wbfRW3SCxJBFMsLjUeozVsX+8gcO+Hrw8UvsgCmq5b1uBoZm7
rzc7IV8Q1aDwqTjdraH636/wphF39EO1JTAwFmXaa+rK5uuhsdYiTS/9xjWLwrejDu20hC8+Tud5
cqQ6SUkDlRPLStfVhAU/rD8HXmiJCkCcvhfTOB5GK7MqNb8KdsY+QcuxOQU1b7sOsM7U1hkUZCB5
nvHhm9EwtlHvp0AT3qblD8Vc9XSX94Cxec4pHWXVH4qhKSrHjmhAjw9FOg1WfFMy3UIZTfMPOCkF
KHPEvCHkZLwQxlPeY0tTw/AeCuv5zMdgD71HBibCzT+a8l6Gq7URwCUCcRyGVwTr6UI234zTqRsl
WUFBTQnH8eEvyzY4y7j7bvATXzgQirK3rI8hJD5I7A9LFoQf7iha2rJdP2/fCeuaCA5yuKFwNhKR
A/NiWofgPsVSdJpJqF/obI0vMbaDEEU6nQudODk7z4SyHL3GCDYo6bTHiSVd6qaQDha33sAjoIaW
9BsFfNtfTP2MPnVJ4xlj4Y/LT0txZKScWNAkxuO43e0ob/4QNeJDfnHhmyyeuwrSiVP3HiCr/iXC
NID3nwrT0X32sP2EgPif5yQ3m307AjgE7VpnDlx5TCBa03hvkwIKzlzcYt98CcPztLNI8bEJyiKK
dtN0U1icl77Nr+hS/tz4hTmclpadZ/W/Dp3QDI5hnf10egMBzCmeEQ9z6rwtI9HqmA4RTcu8IWTG
UjJFVo4OUAj2kUc8TGSvPxsqAI+VL5nA0cUJEj1XUAjHjnlNAhaOndnDSUqbzR4BmVgsdFxC72uo
2eTjBrx8wxiviW+hcjONP2tD0mHckuxeP1DJ6+TFbny9/dcN5nDsPOFctVBGowwOAGnlpQfEuaw+
c+tvb1f4fnuLwPO8prm3MP/po2XBo6FnCHzSHegUMFyxwGOoVAl7C5qZ8M8v/hTolz55p9xk678+
JG/No0h8NhjnklFGwguJ5etcmRjpMUOgS1ci0X1O3KcAzwvFgaJjkCoGi+qAA8ZmyjUK0jvA5ux0
r/Oaufw1VOVpmLiydrpGFSX3AH0kcjkujgA8vqZobi+Mlby8BQUdxFteqq5ja0XUHndyUyTHMqyA
z1oIfUQahYoO1uiJ5N8KtZzf5isWTARuE3/w8DQSZgTq35G1t13LF861RdMzhP/evXLoBl/9b5sf
Omp51Q0EcQfCy01xZojiMISaTxUlBvXcIx58Y2lSqB7Bax9WznrP5yW9SuRoFPLDqWXKjNsX3lvD
woPpnoG5CeMRMElIoRJ2xS5PVM6ownFO96PtPcb6p6WmjiKhIenMIJny/RwOuw/Sr6FHiVRymgOg
Xui55u2XmMvqymcMoizUTUR+9JXIN09k0eU4vj5dvzMx8yDSEb9omGH4IQvD/PmntXdb+suqbBFU
uz9lQSG1w+T46ktP59cUT1v+PldPmCK2W8Hewr6h/5sYXbOnsClMziEF6Gzn0wf8k/O7oem8UGmf
orot9aLl5pBHxUzBxmVputuW5uHqF9dY3t/lUj6iZeDtEHY3Gk6p9EaAjAquAuOBgtC3nbwBjyHM
1Z/UmDs44Yrr71Ri1XoMFdIsgFIOXug9Ycwe1nZm5gFhwVFrymTzhfCmDQYwYWzjfaFxkkJe/7k2
Lmlp49pRXGmCuPrKLs3PTsI9cA6OVFIMVvvK52iiOXp4APn1fN+ZwxNtPXZCrUuo1gT+qZVgrrPv
ZDErL9OB510x5pr45SEfXH2Nr2KGt2pPiaVciF8/N5faclRvrMB38dD1VnZiR7gPPlIlBNG2FKZe
PlIulFsUrL1VL5L+DPk5/QLgpY8zheQTMSO8gTNbEcXx828gTBBCkavoJaRqwmEfQH4+LaMPeCkn
19gZdI09qrBHiRnIDCiRm+PFbXmiLNkr4WoRVl8tsH20WcAylyhtjk80EbGtNikqYt067uY7PeFO
3kZTlFUem6F35W8Rl0iDcfjT7bPJMXQ/oYkf/jjXvOkd4EVdf9F5nqEX6ftJ3rXv/AlWKkORkKnn
UgCy65brtJsKRKYTKR1fIm+lpAWlu3PXDnnLa8L5/twKNVERDAZ4RcXBwR9cYlOKklhTbZt7ZQ6a
qcpgQsaRq55DXt6evE4UzmL6St+8nIcfKwP472r57kXxCQjYcxjBdbxG3jN6eiKoeqSOE5V7qfpb
M0PDsaTRWUfqv5eFIL1uhxokQmKLlwp5HqWXQlU4paAomD7+1dPgx7S9ARWgqNYHnKw9aiuQ4vn+
Jkxoxoh00lS3YYoiLpNruXbZnkX7uAz68zwcN1bVe6QaLNAgAjT6/qnbbllkGUNML5k3/3x1ceEv
ZYJ3YAyuNLG5FQkvPmk76CRUKxX7VPUVM2hNfaGfEw6sTf96OsTcthtHU7jPlYryXhkeZTC4a0ot
J3SDoEzqc18sZbjSYwqLXqS7rYuve5yy5b8R8SBUmi5RN3WtdDm/NBQs7CFo3a7TTRPL5L6Ze99a
z+XiZmetMjOcxAd40JzuWM+RQKu8/AhG91Maqeb7qUlq/elmfp6zKt1DzRRdAmW0F2Aon4kb+hoz
O78WJsN8OHc3q7eRjlUkblvpdLRjO6QCB2m+Nv2x0emflCPBsS5+AxBaAmh+2RgeHkL7HzMJs0oq
5ys8mVMUtRQLIHO2s4dGOO7e+JhoLsLsc8zhJn7erB+5oNOnbjGYvnraAX2zMMEP7eZf1xw9gLHP
hHe8bJ2kfGPB+nefVNBa+rpOCD1HcEruOaQ7MTe8PSBg9nqoJzyPfIR2vSm04oFKdQ8cpwI3W0wl
UKI9EjImsrbQpEILIg+rG2fZq2dU0nFuXtJ29aN1i85iKakyuBT5nF1QvoECwINmM1XR93RA+m8F
Sk14NiOWRoP1WTlMpl1tRJcCzvg1yCilA6NroB8CkQaDbnJhK/sCbQQVABugUxlL0BsHmeqw498z
sN/hQWNSwxfROz1I3SqWjC97Qc2+3IwdTnagnlBdv1Tzpv5CB5EmA3yXRzWN8qOIsH1u8dtOGQo7
jGOpOywcKGVc20FKIwWFt+mwYTvFzcyIrabAPpePBqG9js9vZ9sYMWxFMvIYoTbZX9ohs2T69SE/
qMB1kJPt/TpsqNOOoIqhTD/GPgBiOQ5dE6HoK6fUEl+wp/2IFUMmr4Wg2Sf3DGShegm2SARlwJd1
jkx4Bd7tCWwcORcrTVbVw4rJse64burTEZn0YA6Px/A92lHfa5enY6nQGzaA7YhR8rhQeQLZyE+o
y+3dz5Wp99WogyJ91pynzUup8IszfNft0+gIBKsKWkgeZusrVHoY1Dqy7fwEe7NREi9Nm1ZM5Gxm
+hk7JVP0PRic9ltau8tHUIC2shc5VaMB0LLmK4f7Q/Ca5txb8b6JQRumuzCbKY5yjBiAtsHqKFh+
zhBi0cSxtxrLudGCAgPC/9GwgpRwo85qyJdBZa6E996Si7Q5aG64ZNYbldb158CoGq+q7N9h09rS
krw94IeQFbjqGpV7XDcW/oPswX2BgJL6FUfBnCGPQO8IDbOaiQAxHp5OL/scCpfqZDh0Qioqilqf
0hTtuSFKmZIDfSD8D0Uu5zjc9YVRhvVK1COW12fZDiXL3ut682n3HDxYGD4bZy0FkScIkwSNKWvE
W9UpyDnt7GXY1wXZD/SJRvSimJHoQe0HY1HjIxQutPTODtNPRyQV3lnIaO0UYzkgUhhwzp19bM3r
IRyaaew7UzYfhV6ZLMkXNrFKSFtqkRsLdRifkX/E9LWBnGf+dfVT9KSNXAeLxLIwJCWVDAfQPCgI
X7cbvMrfBENc00jJWOtO+BhAFlKIpPKBk202Mu5AC7wcNU0I1W+mG6+7lOtankV+VedY8SbF/hrL
S8VSD8scypVnaG2wMizwJAn9CoK2Sv0ADwXypfR98L5yjhK9Tb/v+CL3h7xFPUaZRxwZQ52RAiiI
CYwHADcfyDcohn5EWKSSZ2WO/jTrwdhg0grhG58a9kv3CtlJKj76cJhKkLpFVdSc36zMJ2UWpSUw
ksRvNFUNieR4DCy/eOUwS/INq9OJ/Gxh4W96jiP4jbRwt31CxGHXjeYQ1JJnfUQDTD0C4qEyvZ/C
FADiqF8w44msrmyp8er1IAzWl8TAFR10/us7zrzJwD4HAI/5Ngv9TGGaQtVPAAXcb54tQ6fMJZmX
rgkjlo8z5EQS5wkTZSxZ+w7lji6FOeO3lQMeMoiSYi01dzUkH+8yD5TNvbRkDtQmLmznWUDH5a0Z
r3wlURLj68+XRKahYgZ1ZiZWzf6oT/lQN/Ylir9bAIz52FIZBtaBguNZJ9p2R8k827f/CxxqwLkH
T4owGgdSCENx7PCS+jfLrwebTqwPVNFoTuxMbNj6plBdehIvE8ADwuCB+9LVqRxj01aYxQc1vr7P
UOwlHjJaXneYUTLo+3ddMzk1lcTsX9nWGuSxgC/wikLO6x9oELwzPt1qeL1GSBYn4GzjPZN6pesK
5BWgpA0ZuKKLNXhchrsCP59n4bSfoznoIvpLLv0LuiIRPPQSYGksJdyk4MONW+vBDOBsWl1fLYci
QI7EZV3xqCiWSqf9IPGa1mL03PGS3SDTu1P6dbIzQWP692OyVb/XT4v5YMxkOjTSNgUAUxfVrk6X
ty2uou1YY+C6in4yo5Bkmy3VkgAD/dPNOezlhcowgNI/Sby7iLE9a7mIj3XbzqlydWZ7bt8SBTdq
UgsWPdq4+tabTNiTZOfMIUF3CcUDMphEExVJUScZ6BBvvoo29JdVPaeKBZXGh8cIUgBSc3y92AS0
sZ7Scmah1epmBVN+nD5EbspopOIeSbHQhtag1wKI7P1ocrqe+9dHkvfe/zj4ohpUbpgbt0sWGVXv
yReMbzzkM7MLm/PQGwoeYMVbGXE5FmiT8/OaOs2NovYD8Gy9XMnjXEURrN5SRsJOqEWVYeAgYzJ9
vMScrAEreb1jx0SyIn4fI0BFBpw8Ilo2x9GAZbb2pgrx+jYO3XmNrlWMBagPgqtome3gY6br2wlx
Nj0VwmXYa2z1Xml2oT5x0FRp+z57bLxmtMJcwJ2sVy39H9sJvpWLV/J2s4FWQhnG5wYZJ+WvinI7
+vqS8t3+XxwJCpAhLCOUwQ2Z8ovTJb8cRsm2VxpXzKVRGAW5uy6OPC98VO00R9v+jWY8wbJ2frqZ
rgvrmRoEhPkMQ8cWsdp9GNGe4GJ4yL6tYeUIiXMQyiUaOSuFdop2SYnwIhSxTu2tmHGwf3Ttkoa/
7FLcUV9Faz3xW9efw1XhaZCYpKbU/OHhVEnMwFtlc53WnsXHlt2LbHyaC5SRkBsQtpK962LotbcG
aSDjbw1S339xdHBwcjw0zgyxOe3hwxkGAx+XmnoYNWOIMRP2KrXIVNjmb7fKjrw7+zzC1UYY77J5
McMYxiYGKy/toMooVhRKN7QT6ASao7BpCylf/1sqvazcMG3Ct8039TWKHtVqrd68T1gQq/W2IcjG
gV1W9ZBDCEtgNXAsxb1e3ORWhpEbOEoen5K15TFOipERJTHMa60S6mFPL6tZ9pFmYWnLfnHf7DKf
fI93hFm5CB3MxWv/+XzxgkxBATyUIf8Qej3fwcmS/SfjZlCyWwTWtS4uA+5G8czcBLMYDfw/jlBE
Kno0izodECzPUyrxfe1of3ADKXKpVZmaARAJWGZy0AyJiNWb4RP7VsZ3/IwSiA4DuK3fuaKky2WQ
DInbC8Va2Z59yUj0o+qQY/ecmznCwhDiTw2M6vqiKMIEPPpzDfK/tgw6IjI6Zv3UXfqGFdV92o1h
9RI0Lk7n1UGNiIQEDncGg5f+o6su3UtKKM+quLk4NOSNec+1Yxz8YY8/hDTBh80tkH77BI5SGJE9
s3W09UuwnHPkdcBjiml+jAQwMaBx09yVXX+RifaiROdsKa/umuGmAGXFfjZ1iMu8+NzkRBLdzxaM
pAJLrqfboKsfrn4MrhhecXqrj4yDIv3egkCaUiJspT5cCfSopvC9i8ghkclWMNXyNyQGpAfDUu+S
1Lq/IMAWjivi+wuQQrycRv8chloK/bKk76PQIVQkiGVVsVPU2dyAB+LF0W1SRoseE0nSgUjWgj2R
+MOngwcIa4VCW45SPwsCqZcyptA//qtIEkqUfNlEsvbApQ2LX2Zbv7+dFU1zCunXluSoUhl8DF6s
FLAjE40ds0YGa7mr0vTVBQZi/GOmSj7+18fndoEr/lUbyblK/GMpVC2tT4bmYoWbMcb7EjoFape6
op3Ye1Ecpigy9rj+EC5xBeLTS81kuQdQYczgH1uUIpS9ojkwKfYcbB5c4igDhacLBE//jr39B3hf
MQmTXBDvowTqfGskP6Q4JCzMHC/IWLVSw4Re7r8BBxHUAdLDvVX6C5RCM8eENV9TZOSUXQLBE0Ou
9dIvoND06ft6ffxlwiSA3dEw4LLB97AIsq0TDe2m322LfYh9ahl3Bg7BHTMC2aooo8gLzIKL7V6K
bPNRm+bZLrdGRMhfgDf8Lb4h7Ad+iCc3+wIEgDdnbpOJUeYmaCvY25Nb/3MnVbezILpKSzv/nY4D
ajDjtAKgUFeR+S33RBs0D4yU4mdR3208il5OQY9ZvGWiYblfXiSS/35LAfhXaKUgNY2KamJnSgNS
WUhxPR9MvF8d3eYMxDPjYi4ZDenZThD4RGRE7/AaaKiIkfGHH89nvwnDdgvv20zqDXSI3RZgQsFE
NTy9EKAr2F8W3NJmY8/J/3TGjx3S+OgJBZIS5EExbqJJ18ZIAWBahen3FMrao4q7nBUy+GUMICMR
ZW1I43Pt5PWk+GoZnaGNmceiR5oTeXDMy8M/QwY7cFB3GoxY8Xsj/sr5uuwwtO0vjBhUjUjp6Yp9
cUy5/MLVJ/WeqHPBSRmRIaphNe086ZeYvP13gNkvYj9iLqXwwucS76SWmYVlqBSBDLjVHjQxBhfy
fZCokAp0upFYdOwbjpinYPI7HFdmoM3JLuaQBO8YC3Th6Qs7Xn+15v2yARtHKPMeYPt2w9WfZgCp
7OA+IuWvT+IqW+QNd3reXLZUNaeMfFTvyOksVEcBRxCiDTcUi9ZJksSZ8pVRD827CTj+eib0nT6v
VYJMkM71heqpVzjL8VsnvfeN7/LFtRwmGSEUXuwyHf63NDLnAY1748v4RNC1FTOO98cbcJAtTxW1
PxwsOrvMsPrLU6YrGmatsVukInnZsyJOp9pwoh4/Gdq9Mn81G9V6/DtMNx0lqYmuAiGffueOwiFT
4ishcveshVwSNhJCZIt+S14mGpA9QVjBmEVBNtOgxq3GUroF/agj5L9v6yGTH2Ri/UwJ2a4pk20I
NK6zuLuRlNEssFAz5lWrsCbGItm6h9jSdZcb4zucwOwKYKr7Etp5zY0RQYfSCXRzR+Bq6sqOhLLu
pIiEZ0SzSTo6hEG+v2UounnRg2atdd7F/QGOhe45ghlL7KgMCeOVjeWWuasaacjTkhMotWueOD73
kn3CLRdY4vjDKwo/1Exr4N88uC69+Vw8vM/oPVl9Ls0iQk6sG3Ye1ycXC6hpDr/rixJdG9omstfa
5HVT6JsqLi9bCddrEbWrqoJD3FsuyGVndf65u4LJJ/5/PtATFq5IJab5F8p9Y2GDUEMQwUvm3TtL
6/CrSS90RSeiyi3L4x/CUhP68ZTzFs4924VuHImlRX6m894dHbCNo3aHrotfeKiaX4yF7fajuliy
JqS20yG3pKACEw8XiWXhkLcDhZKGhwKZrUsAASZRTylNgf9tKq6tRTP2shYrYeorsOcIsejaEz3A
cvmZ1ovRxG0X7fPTEs8FffotrZUpUaDD2RbZkNd2Xk0s5vFwNFeAS0p7XOar2caeaphBQ/xqDXxh
1fkFhF/q6sVnp9xAx7cdV7o1L+shbPB3YfAjKlKwNYfeKg8KnMEDzRjfvZ7Uf2SGtjEGUomgJK2h
ktsfnA5bbMbxYEKt1O9QcgbpgL8he0LdFrjpWzwk60I0kiq5MLmR5bj33WoKW7Cwt7ez7FqWmET+
+K0ZIAsZxXxWQWoyLQLjzdK+Rv97uqobJCbWjO77E7kMBqHwWkh2d8lmMp55TGkB7mnX5f6EXdRB
q0ZztUwxzhl/D2gfhauWrcDWa8kqzBTuTy6Bkvh8TADXWodvKlvNAafdWnst7JnXxh8WRVRkaAev
DMOn5oDsPDlUB13O2eO1wrGkmTgVQbTM+pX709md1FXIdHOKK39kl0kp+wfX+61bFf4Z/r3g00iI
QriM5wXx4/eCWtHEcBTsPF8ayu6suwg47dTR1iBdkH6pZfxid1fLgHq0cM7auMCHBptpj6GhJu4X
irAID0WQa2YCCbgCIM64+2GzDmpJMqIPC+uj/f5/kVyQMn2/R8fjRy+EVTVHSNXBtFlK/+S7OP2C
ALGdFheklbg4rdRp1NLjx24rX8rXzd5Ckleb5UoOvC3ZamG2N8Vwz27PprUJA0eDacuaj0zY/H9Y
d32AApl1PUhJoZKdSpBvgHuOvwcPphIocuwrMH0yhPXtkUq2naFCrjjyJmtjq2wrWHXFzc4Layu2
IYCP3zvbWj2pXdY4ErUfttCQ2x42n/7DbVAwAP/a6I/BEj53fjP10LXytZhcj9xUaSwC7CMY3QFx
kb4uYVg78BB7txtBtTpcII8Qg4KMRDlCyfqDwyLWmuXPqPPIwusCRcLTg4T3DkYvg4IB598IHBv8
JkJim2JCxlToNUhAk3N5dTN0YFoOLUT8awX5N0k41uXdjiYRhZ+jWGPJGR6+ZZA4khnU8na+mb0a
FSluJbf8HRbXLCon1LphiniKJrsK23doThZ93oUKj8WpRpWe5eK/ZvlmKBEHudy17y5QpntPh0wI
7IVJPYL7KH8L1C4U7mu8jEkEhkPcNAo3dXlpA6QBq4xLqXE9i1Y4imgZsourv9wnnu/A8CcVXTnr
I8EgOnlhOxeAFjVHk/u7JlqN3uvjCePCG1RVZF7lgdk7e9ttyOSWd8MnUARAoMAgtoOOu6MibUBT
7GW0Og0Ju3h/Bqqo3qgio2KWGrQ3nzK76K3aU7pRsnqzaS+6bGjpPDGmsabdVeHKq88xLkOB/Tyg
dyRvsUhYlrAQLSiiBSa7nU/wu/Wd9AWP8uJVgy5NvXEaJNsRp5+hFU4zp4/DW25dQwhbZVuSiJbr
Biqn1WIAYrG44HCogiUsDbWOR0059qpHJkuTGEnvXGo+FPuTfzedWzqxRTSjZMTuoClb/uf5789Z
BmRzTz2mXnP9sYpFHjlDuok/siwcz3YTFF9dFxId8pwiRQRYOObD9xJf+r8BN8bJ/I1HjgtccG0Y
/epI+ogXZuSlLd2yFg3Z/YlRF+jR4UmVQclwQPR1ntJXdYhJFj2wPvNKGzu95CW8BxTZXTk+nKOs
V/Gdr71Kjp1o30zngltVFVRwqGdEJl5+KgvY5LrX0bC2PXOJS0irUHVUzqOou/WruxG4VispHKLR
17BJnCUBr0QZg9hAgYoPj3P5RCTr1N8nSaNv1XfXq/CEh66+zduppSl9ckWT6Ror3I3ndmCcG/mJ
8vbQK9FFP6R0gzL+xe9p0PgoI+JuMzNA9BxcLEeoCvfP7AHJpVH++eozxXuu3zwyj9lgg+nPgeqQ
iAk1yIwNFFA+qbB/3Mtv1u2fHghRRtI+zw6TttaA9flJEXiy88pUKrsznaf4n6R6KEb/kaz+3hoM
zHHfDU5f2DOp5L7BaqNxYCYb2boqoXWcsmt6R7wcbSpPBo9kNyucUpcQeNR1SasdeJ7RTAz81vpy
ypcZoAcmxV1bfMTtF37Q4l2u8q6NRaWOrZAkhSWgzjBZRq5IWG+9sQTYoShGZlpoIA/JAIWPpku5
sM8UVfi7mdyl7mkGtxfrzGQOb6gdG/A2oiaKHMcuwV+hQsxndDrbo/jCFowiGCyX0xMZNBR3a5cw
YC2xx9YMaiCsfpfzTwSD7rU9z7RIObrynV3hwiTmeYF1r3sJ/7KQONeCKtn21di5aAsCL7liv07y
LtdTYS7A9AMwZamIsjRD62aNUQn7woMHWgE8v2W7eNZqLL4UPPoUkCsTChlXjPg+BVeJECL8fS7U
rafn8P6XByZlcauwuyUEFryql0wOR+Gaq7l3Jo7H+Etw5ELF9X5R1oqv13YyU5DpgBKm//AiCaLa
bBmI8Lls+npwnUGxoUx7LXx2WmY4yJ5qO9HHOo+acS2voBGTnE+48TfFRn9JS4wtEiFro4UJ+xSy
lG8sa9mdqtAPgLmXXE6mLB+u9IATMAupjEmstAZj6Gy3fArm+M5ulpd0GbyT3be/c66wlimKSQS4
jhgPX/NBN+woR1XkeBW0k/6JH1EYwyvgXx/Sc1Tgyhxm3kuKXTJZGcfjQ6pfMoO87kjXtTl6HneE
hUrmAW8WbB30GeUGHLU14nZSdvnQAltvxZ1mf/A1vlZuuQf11l82UqeZARQ0BUGNM8M0JJCNc1Rg
DXcSwbW6sjk3VfpETICVzadqJrAIl9nzRLXNVSM/Zpy8x0EyaW9XjlNbiNMWPlI/S3gB8vXM3eLq
bjRj6/W9WQFcn0P1MoCigoTZi+pfDrxoJ9l14iorUm36WBCDU5F/pC6YE3f6IlD/Z54rw30rR4wB
eL6akJxcwRJ23OZ1tAyymLn95Pd24PPB+FmE8ULiaQ9V3gSha90/489Skg5Gw31SjMUstkEPMc7m
ltwa5fHcQFqHvAVLl8d0kC2wgUqvfSw4WSxlHWGVlUP5uMD2fxVicCRtGcHBzL28CjzxDeX3wknJ
Yc+TfgSdzEXfXKGZQWaMivSJGmWi9LuRcfjy+pQVN7DQdAq3Wb6d3BtiPyx69QoptSmzJqHuWtlr
RaZ1Fb9wOhlnwj03jtdyGokugqG9tL3w2fF5PBoD8xTWNwIf5QKDwvznwwTxf5sfO73lwjJVyOuz
SIX5cYmIVh8orrUvubV2/OE/sGwh5z68rPOU6u3Sx+FFzYVhRo5drhnnWD/pzkOxcrfqZQiU0sWl
frOnNQcjCV3X3W24i5F7l2NFKXj7ePYdny69PjymVpKpTcMTKt8Fx1+C6Mhren1RzJ3hmshYa96X
0YQ8F/oo2vboCqVr6/rm4MVWQmAwQYUXo9npjFzA95kbS+ACUCVlFyz0i1nF0a5WR6NMrbwVBliw
OQFT1k+Saz4MdqeFkhtF1KCzqxoeUAzdmV7QbKZmXOq9T1x6YfedxXFMjcETY3spQScSX9DZKiq/
yL1tlXkLL1DPNM6TH8J6mOQqKuR9lkXf/7afYgPhqQx7EvLMsnyY5oHStyPtjpf0O1TRTIvZpvCU
GllBSduUyBhEAKzCf+22vja7/a6ZHpbOOfp7v7u0l32nYXHwROJKO5u81jndKkInSWsa7aGxRr7Y
l/z9/dYRxCyc4/5HlN9RjfY+kgaxgTqBxMGTnovAChG7t1s0cgvQiRcVQo87C2Lq/izBxVUFPheD
uDKuvvVA0kZ7llGaj95bsrP62aPXZRn4OsXXN6a8Eqr3UErNk0wuVqzElxNJ2Xr0p+yigWlX/NNE
rmhXNAXOyCTlIXc1o9IzzqxsyMrSrrV9Dr9Dm6mxT4afT97Q6gGwgl2f2ZfRKt5NwzGc/8lXu+J6
bxdavAYsx4YtKFtHKQ8U19XZtqjLX9ITA73YWJLvpl8warxN4BH7bVRySQQYH7cwFPLmsCK48l8u
SAU6iE03qX6MT3Kt6JNpBuxFX59fngP6wgSY4q8ED2HI470cB2P1pMWGUjWFNCYxO6gkSNBq5oer
deU3Yoi24sHt5PLhqJgIEbvznraj6T/eHefseEQxLF+f89e2cqdyW8eJjH0VyEeq4crsYWjwIOxH
jc28E292XTZiX16jnj0X1jfP4JaLbMgEru4yxFZ5WZSDiJjLgSqGAqHgr5Zf5dnzk6eKO07rwcBR
nhSm5PxWA5pYFEo6wFym1bmAc/qqTQN8ywMs1bSkNZTuLvzVuOJnqXQdwxta0Sq8YxQ3doyB0Jz8
do5xzU4TOiVrrg6lNGK1YF4B/xnVanNYCjp0xaLWrfl2zE/6l/gmm45/7nLMIb8tGI9zz5RSLz63
7v/h3XZatl8OQQV6gBNJOIAi7Y4k7ECfpxau9s53G8cyjFFmjSUOfDdp2lOnSz3CPU5uDibenIA4
IT/99J48X+nRGqMz+2QSGWLxrsA1dt16ClyDutN6Ae2MeMRnu1LSzlgGQAbaaAglUXfOYOFwHhI+
2Zn7doLDpMUOz0dth5hAEnLYm9F340OFWI4dLTIy/AwQSHA7OAu5Bs04cgg3j1DTR/BSpJ5Z/hjo
Cufs2vw1/+lRuvx2/OV/epj6Jaiw9iIN++1ArtYvRha0y69eK0F6Yj6rAWDobetrMFBb/c+HyNQu
mhbI8HMfSFnasSAJiaeEJNLJvTyhvZvBj3+qyx4XTEb8GDdZP6tf2RI9oZI4JyQMUgdvmN8AxhPi
G33XP7PbzzQxvIAJ5/2dZAjbhzOaXJKkNZelbMjM/uyfS5HHXh4moydkUHkaemdOm4cdgKQ9voRP
0zRYkRvdWonIr9LA8nwogBNiMNdZHAVU1vnkF0FyYbOOV8t6n7/Q9DkoBlPHtMf9q3FFoeSS15cm
RuQxGG1sufbmLy6cC+6vQWx2iigCF/MEn+n6Yz9JQICQlqa6367jerHvQMnWXGCS8e2SFyDGIZKp
uW39YD7kQU4gn1YG0ZfgGtuuOqbzcNf94sylss4PZXxCpcIwJ18aolLMdx4dG0ff6RU9PsWw5qOR
4mJ5YJMexunYAg8GEnJgkuoESg905Q1TNht3gwlEdZTjkys1ZCtxl/gHTYfywanKhyvHDAmlI1R6
37mfZdHOOk+mleYazZ+9IHWxLZyMTKzgj4W43JirDbsnJ4qFH4RlFOgfRUGu6PBq3W3e5ZTNHPx+
p+NwrxRVpAmKOA1AWv1jBgfoFe0RcFQgfA4HDzNG7F72RDPtHAvWZJHJgMGKAIhf7Ir3zb0aIZ+f
l20nBvoTmVQYBAZliEsxbDAdVClPWKJhfhs3hsham0PPILTp9jBRwAGwVGFvOCuDOncMkNIAI7Nq
qefvZTkXixHjqX2QtyDRBR3OM0122+4Z9iLraStleKPLu0YytcO7NA1YnjMDc2w49ox/kSYR7HOv
ODtuUeO7jm+Pff7X6Ezb0SaExFMQThW6BVugTAXPHzNg0DBR21ugFZyv8Bk06kjAVcwseDSwHIfg
xdk79vvjXiFxtY9ZAaw/KXPkKms9JsbJsq3OzEWuLPsW0/dpzs3whl0oQSd8mS8ZCSZC1szYhN4M
Qgf5TiB/Za5lRaeF859ZW6pixgrI2jcJ8lp6NjceyajXiFBp6d5oGsfrJ4W/+kDT3XZdRsohbRGO
22Yjukj9Q8NtpvBDh+kOjEQWZtrxzWrdyTQoncMZHpk6ZNEP+WV1MS8dlFZJDcxeZSipX4hkrP0s
xv3wgLv9E3yz+DZV3fuigBZ91hjF0DGAwDDO7G/IZ4n/Ua9OSwkUzSsKCxT9LsPP7TxRasu4gulX
XKy1Bi54filt9ND9STRGSgrt8QUEGVtLm6kmHt/ClEeKwiqetFes4rgHtbjfMWEA3O9iVlMVKnh1
QWQr14JwmzWgOu4tcz052YuPpXJ3HIMb2NLFzjO5VjdO8Q5cwvYrL5aN8dk/B/ZMt6d9l/NlJCXX
1WwIt8blhbjdGXyJ3Z0Q6LE051RhlEyA6i362dSVTMeRkLlgOxBWGR3sVD2RmZs1JOGXg1E7q3PE
0M7WiSWOTJEsr78RHZ4T0eQu38/DFsMNWOEvfSNNE4cYK13iiPyXOGkJPsA3ZukfzfaucdK0cimz
hiasHjhR4HfRy1/OxD5RWlBTdhAp92+/kezuzskZ2+1xl5GEN1FoqljBn9YlMFHQEWa2qHCZALYh
NtgYVJrPqZP6LdlrdjMv+IwhdOIRfcBUYXdFT24U/qDpu0zLo/u5wc79jo6I0NUr/3VAVGgjix+z
EpAeVi8dpHcV7jvh/FyGQ9tbEToNG92/iCu3/kjrpYrV9pqKWOUDOtbZS23Wvyd7rwegQM430lw2
H5EvYGMRYDI9pK61S2gz6ZGqSPQP70YQhmmtd7gAiGuPDqG612Rnp1PkAV98pA6QzCln+oKE9Un2
UYpHkNpUygFlAwGDryzpOafuKq6dRY2pnpCL+/ZF37ArB1KIkiBTXdwTf2qr00GWuSAd1knqNo2s
+nvxOmuhmqKN87Hg3SaNxHuXa2iy8dXQdf1ygezMktAb5WoNNCeV2IG5O6+SYPJEvxddaGeEq2rM
/bY5WDiacbULxzmqj02UDcsSjW7zGJZdvFDlcP/+Gd/9q3njyj8/xsB5SfIu88Mop0ySsRak0c7d
OXBMjsC0wpWsFASa4eofBZN76SZ0QD63whcoXvpz7mMCuuC2QzGWpZafUrICXFd7i6Bsa/TjtVZ5
/CCcJBxcfCil5KTrVU7nyej6ybUsv7KDOp5yBm3yU63I4owmOhH7c28F4L63l+h57scO+hVDlbr2
m8sVcQMpN7gUta5vka+RlmwPuGAhPJRZIfOYsTA0aFuUCb2zNyVGuUY+nf47ptSSdKlAp0MMXoLW
SVQ5xWOVz7g89sneB9YTJLgQnCk+q3LfTMdSl00q9VxD2frmKs3gUWFMgL+ISlxRcVOFG4wd8kd0
sKuVWRpsz5lQKydW3FIEIGh1TMmutzU9xv6TaTMH7NSxEuM1JoKC2O3n0XQPCL0ELleR21zhWjjQ
aGcOng3jY9Vx/1Eb3Sl5fqOWoVqisIu1nHJgWPCvjQt86AXHqMt95b+d7xyC1hSGNRFZayu4helA
7+TbggpH6C0/sOk9E/2vmGpJoa+fYqWe3Dw4cqatM3L5kdMVMryPn3XBXW1ghx4tOEH7WsuIzDlX
3u5L1ewQfE1MHxwlkSTrrDOIyZPI+lwedy7E02p6caEXs5ySqekaRjXGsI0YvIGI5qcdKVCDavCS
5lRq+EYsLSGpo8VacBaFLDiTy9LkISoG5K1Wm8gFbWa4oC2/bQcLwHUndlw5diBvCYIhJ2B809Lj
iRZc57nDVwaMhODk9V3jEUapLIQ1DaJjiewiDZPgb2x8oN0DNw8xRwAPCU64DjQPOsfUYEFNFqjW
NUzWjW9JeSdR0U4T/jM5VVbD03KfyXyYvLELLBQInWrhswdbTOHrDxX+8LM4ZOif+O36RO02v67n
U+4qZDllXP8s6BWdqr4hwqrEYLquknigvOfz0emb1xBG9m5Kwi6nDPqr4GLhXtaL12jHrBnPJZV3
7nWD0WflbAa0Rtqcbh5Nwz+PPl29YEG0SqEreZKUUfgxofXzleLPgYjZhdNjXKEHuEx6CtlWyrUa
DkILNC5VNDMkn0vn5wGLyS0Dq/tSTmPsdnkvJKNidTAuwl8oWUENW88KX7xwNcd1/o3sesrOXam5
oZq4+WwT6lXfrfw5HLUN+Czyci7m6Edux9xi/el3jHOc4GgAKHnOgtRN7FLjUJJXE70XRLdUd/Xq
qRt//YGX7RCk6yDPhBVfhuCvwKltx+ajGQd4Lhnflaf+ZcVVrZ/Eo6526XLscMSIp12cqo2za1LN
dCcwbANpUaD/FHKnJc//PMSMF2lzOnQlnCtVlSsq9E88Z2b5lMNiiLetJ7F3kmSN8P4zsgftBtfd
2aKGufUIm5T1kdT+NiMwLB2fcwIGDXj5yxuSfRnUv5F3g/xDPE5lp15h/JLztCTtbHL6zjqkLBaw
v0nbKKdCxZJmR5NoX5jQ3xvsaPFa4KW00zh5FGVeVbA3NuE1mGRTAa9xiab6sObbuwhSLvW1Zymw
fDZoCCSNhcsJsD2ghlO7LLWvjiMnu2YEV9JN77IBiv9bMgC2PJngm8UVCpEk0QuHMYESkIpvgMEa
HM1cYNPjlnOS2Bq6Ly+DtpWQXLjw6yNvfQfuhPdffhuk3s6Ou0tQUF7WngGcd+THof87S9RrwY8q
S7yrB5JcnsT8JS3GOvdhabL8bvKiVxR6VcSkqEc8JZcHhC3QU+U/eHJKFxQqTWSDDqu5V/nbKxRV
L3ZyOAlrkVWVdBz4FaR9pEUnnX8hwUqE0gGvS5mhx0crzxmreuPsg3SwacykJLQBb35dU7o3t0Nq
CdRTVZxcdUf6r/EMf3/V6ZU12PXUlDKj6LgorQFxspjoc73v/kQGMQkkMxW4Vm1oDzAdWXDtZSaX
2DX0nF99nl+UNRns4i0J/LXy7ZHwQEWODgaPF4edQWeDXZE+9wTO5TsADWKmacQKqOJM14CD3+S+
Uv9JsiWXq5+JImz5FnVkZrpjlewHOJzzkKqfDbhzrN5Z58A4ppz5p3FK9oLTPvMEVufdzihvXrex
f2204VA+o0iDcS52kzMiF6zusYkvFe3T2Uy6jC+WFuVvjVKLJRwzvws13L56xe0TUOCpN7/fsXrx
JL3WpULZSO2dVH4lrBUgwF+YaCsTfx2k9FDzihkijuuoabTpDKiJibuOa0CyDUKe+Tlt79PAItz/
u3t1tlxzjXlYVu2d57a7mLwYmotXn5Kjd9SRJLLyFrmker5tvW7ZRokcbV8aFXnGeJXtna/eCTq0
9AV7CxjuL3+h63SsfKwNbjqmYHDEWiPNDmqyJCr75nhsMYUu4ZaYQ74jvq4u0hHHh7+kqQ6OS2mf
us/ESn84U/i2jLRvb0q7EUzSvlv5m23UMHRE2GD/J0NQL03hPQp/h+5vogmqLEAOs0Y1o7pyNV9B
hyoWZ+ACPYXu35PQfPSbLu18zobZmemcm0VltjALGvpt6Pry2ZBc9g23xKwRl0X6Z4FhWINVD0p7
WSeVo82RmzE59TnOFz2vxnT0uvJvyi2BfLf/BOeJ0+8JMNJOUhgMe2K0+/Q2+RuQwoIvoQOGT8W/
Pr+4J7mI93PQ9YpjOkjOnZUQKOlyOn/ptV/AD0uqedvMGkAwbaE7jFioi/Ke8rkbSYn+0oqPSHlQ
4jqCMVyhGcK5Mdkec7q6ySORQSwrs5KAh0KlcMaoug449mHDgtNcjzzwCWh2kczv9t2w3bDKAuNH
im32IFZcdDbX49kEVf24oR20hoTPquh3mxum9XfvkTN14N95r8Xofs5qPzWoPSk1tfCpEoU1u+Dj
V5hiN2+L2TG5cJWUVPH5YXEL0koPu8odEEUkH+a3rJ+YZAFjWkOBZJhsDcEGfyY6oSHFHjFQV12f
X07m6I68AY3s5ReaicVZkvBOwzQpMiEtBfW4fFmJzPJcNlB7XbcnmApRHh+3VA/aJ4gLYUi6FPjm
SHxKCf32ZW6VTiB0cCVCNdUFHTRY+5Yp24XRllHx06E53IA4uPibd5r8VJ41Ivx7arBvftmSYZLS
bFLfE7v8Er9W+7d5xXmaoiNBdNUonPfB3Xx5LUuSl2c5m3QhIgNkD3EJG/bC2e2ZGVy4xAKaLDAK
MmDlDkO1S3dcoJQgnG1DBk+CPyESu1/2EdzF1zl/n0sCq+U6Ttzz6dg27XPU6jVW1QNsFPod+eTo
TMRoosiKBPZMPbtaaGU1bwrohK4UcBBir5kZzZQY7YOOjl0yIIPmX/8Rog3g3L64a+7EzNEg20KV
AgLjqY+sk4aRkdRnLLxdeGtv+guH/mRTZV4YT3xGboOosNRQ82ortrbQo02nMtP9Dg3Zj2J5ptbO
iSqn5alW7MCpMuJBaYlch+tFi9ba4aRA9d9N9TK0JHphN1PZ5yXH19p+6WSjDUfrd8z6+5VC94Er
YtDit94uRkSv5+7m3xRJRKbklz8Zy61af9H+5fkrI8mekUHgQTV7qXyXwLXyBBmC6paxOkmLiCd7
YLBkcZVWbrVoYBqjPEsKw55KP7tw5yNbMkbot2KplIQlfW0Q1hYwT7kv1pL2gIta3Z8uaXVS6JqN
MXpHbszFKBk+/e1bJO6HplTRg5YpK+2qUYP1hf/u0BhIXMdTIL9ObXtJb3VZbhxiumVmpPoJRRIF
bEGbE0SHi9BXmgvjUvtQLCcnS0c7cznFjIhc0F9tn9V/BZ0+Ny2rQnNhICoP+qgWo8HTLCJtwPKT
51hCYrBO4BqI3H/xlpTnB5guKrS4v0+YkjzpeER9C8GwjmMMz4yVNBLcaHn5yOkhG3xX5o9HjNIZ
LsGerGtUcXmM45tbj+v39czfwY/iaxZZBbHvzVnUYHGmgdX6aUuobE+/sP50D+dJF1yleSF0diOb
TjqACSyWVY/5V1dohe9hz7i1M7voevW9E3lENhGOTzmQWv0qjKy6blCrLcTlzlDMm9Q435ybKOzO
QTB6glzipvehM01afrWw6Qaq78pkRLDgJ+rvMsHDh83l91eRI/+qJm7KjWV6oA1RVjghlRlr/lm7
GewzVYmmJj58MzKVF0R6KEle8vsjdFitLsjcQXFVni+MkBNiLrjovaoJELIhk9Ec2VRj3Feo8BXA
q7wooHT4RkEbUekzs2PLxnfYaKfxgKNk0Loh1DqnmbsLgddankcFBUovJpU7LNj9lUJL8ih8taT4
abXfrMMUqkCD3jA1LR39CX+6Ie93cS2dyEUNxbLTgh3AoNrTa5fL9PPIAxeucIiGd4fDirKgcswv
oy63MOk81GFoN90x54i4PwnQAceJbf9UWGv4b6CvWJ3EQeILXci5MRD1KB32anW8pUoKT7/aWpNA
Nu8rjwR/7r0XqKJkvSuZxAIfWQUTk9XSTgQE0QtBU/5K0euXhalKsos1P5AatD2BCKhjjywgRQPv
6ExRTUyo/ojz/SHSHVQje2Q+kYfcL8x4JRNvtXfXNUi6rPQ0eLkWGGYoUiXht8KaKWkxRSCvles1
KJUV+Qhw9v68x1Izf31gdtwfTY/oP1y/eZHSMchxTfkbyx3drL2WZWWuJP4mjaHnSPo6n/xVddvp
sxV9h2VV316Fv7EETJdv+GHm95xE8iRKLgmvo6d+O8qQ0zFAsIrNqiOu0d67gaqK3T4WZTOag745
EHbvwEVEAbn/Ny6SzCCEG1/TL+xtbSnG3bUZWwd4hUg4QoooYg4NN5IIzAEm4oxCaWDa/FCuI5KK
feyQ5wHbgRSZD5fZ0bseTfuRzHSrYT5WBnI5oCY5vldjjS0VIJf+NAyefXDWE0cjyyE3lIw8VJfW
mDIiUD81AY0HDYxji4Yhp4JcY6KMMHkIKP8rwIYJt/febBNA0LTWyHhn5hTzHjIkCenLdMXmqRQ4
JwlwrqjDi4yyYEykEekjE/pe0KhAFNzdDtXLwUJvgnM3jncYOIKoezf/WzOX1ms7z3OJsc4TSvd2
Q+8vr9BXMGUeM71aCIxyjVaS3ruwg0AC6G9aQVLFwfiuchfQhW0ySWCn8GI+omiRw7Km9WQY3JcP
KaHN3NrbX9mB1fnQ5XwGh0+RTu3vQ54UWLdWp4rOxGxW7cpufwpF8ksuy8QtgQhLDiyLFAVEnpS1
IZUo7PibEgj86TDFcxseupi2Wg95QpYxd+8277C3XLooCKvdZo/4Lrg7a69qwpKvEKkmtJA2SUSn
uZ6VrQx8cpuGCCFHNtSE8yQMhgVlkcP8gomteJmudf632M3gSwrz6oLXpYf93DwgEWw2CyUhSsHX
zM321pyP2HzL1nSOF+2oCwCELoF6uy4/KYCmlIGId1dnye0kcP3lUCtZX/g5W2tCuuxGIFBt30zO
Jb3TuUEA+m5c7h1YK+5H/cr7EraO2DZ3bpubWd7U3+ZIQ5q5BkCdhsGai7CWC3iWCwN22eCJSo2p
IBgVu9OHqKUPgfuVfP6XjM7Vqbr2INJ7ENjTc8UDuZPudorm9oGhFcKzCXpYtnpZp1B0/uEEY9sL
LYEphuGdA7pWg1+Fbam2v7k5E808HRBNLPk6nrI1Pvlu2dtQLzRBz3adC0irU20fcnqUIIMx633D
RCxU4uMlGjST/WAUJZ5Fb3NXmHZBdIyXrj7xRXnJozJDMql2KND6kDJQcrHsAG8ZNOWquYkpp0ew
OJKPS6XDEz1rlTMIfkrA0MtqzPkXgMdQZpXKBS8tbkIHti84EjYzWIrlZ6FQnmcp2JahB0foO/dv
QOc+vyvFHMeN+sNWCsjQ0mJAjG9BQOhDQKO8c08+yIcKjOzCyOvj/uMIIj8fY7r+uqM0F2CARlRt
Ey6CU1sGM/We8gcSZI33ZEOReGYIWtPN+F2udaV6Xm2Hy3IvO8jzK/M6tlODif4GxQmWQAUgrCOK
NXLGvd70U/xVOMW7uE05zAD26/PRRq+eWgak/0UODJxZceGnBY1JbDTJx0SL0t7FRScvdmGcY2wc
yNEZUJM+OY6xHATW1F6/YGsCkrWA45Zezb5DOtxrAujJl9pPnWZ8c3P48wg3hKCJo8kdPMPH12oB
PdnwTq3HzDQoLK+gcQxcCt2pk+MpVoF2uwIDLjJmr4sWHVtK4VO5sV/2e1whbsUHcHGRixAQMR+I
+TuQa0tGHDyRXRfFZ3fu9Sn6aO7xnXQ1PhaQcKW39vKNsVXkq33tdl+kOIqkqApePhXt6mxCJcFT
txECwIIzn5Nxt7opZdvCaDN86vgvj6sary0XlWvcds+nSNkaIU6PtSFS9lpA2wvCmWsG9n3TKHzo
uUj3areYUVyPlqIsmdXtL1oMQ/jv7+itMn/UfJw3BHb0STVumcm96vZcqXMDz9fXg9pqUDic+11C
xFDQoyAvGcAvAeR5Ep9IWrtjetuF8RXSxeDkYgIxk5xmFwyqxmuejCaacZZ2TImDDrcuyn37ruNU
m6eph21sP0Z0g8PT7tPtSh2mqGM3ygnQXagxowCckGQfWTm2yBEPiJokfUkek4BRYAIgz4M4VjB+
Gz5lL1MOBNJoDqlpUhHq90R7rzXlS6VSpy8+d08DJH37oA+ImDIV5Rvyb/d99Y032p+PiH4BXsTt
xyUYapfJu/wHARTAa52OCB4MSaGrIEmm5314nSM3JVbjWhRMWG2XQnjOPcPGwXYJjeq9OzPy5WQQ
MFLKj7MDg8tCU9+I5FUk/rQK+uebfjNS1ANzyLQvFI9dHkIeGQNF6StXrKlPWpPPr7q5nb5CuJg1
7VmJiIqKjaY1hpT0SX4id6/wSKuQ8ygenDAhSQ3SMurN04EA8UKbNRE6PjblwSr1fkeYV2cbGIRQ
0abmsjfgjkB1DCzz3ZDhlQw69i6fuWtecGzrqI0dDmeh2TrbuWVJcXXMHmj9GblhKjWEHZfalwEw
spIwVcFdQtXN20BqpvcnUfwhaR1qkXztpsEPumbIMWvsb1k8/K4POX1TnJ8stvZ8By3iP7Vs4Jf9
0KxbEb8ZUO1U27yuP3Q5GU7cuQscLMY7VPgOV8q0bn7cnuhuTp6YDx9H2WEIqOnnuBqvmSOQr76S
J3UrdjGyOvbw8VHnGXOfYDeaTrcn+/ACIpMGx+J++vxclIB4flfAw5rDf/RvEmPSIc094vNwklXE
OHaJPw4mTqUnlE1X5JlRllqEr/bc8gkvxLQdPblsN0bQ7psYLWqGr2DY6HN3WtVPb71F0hDT7kfi
mU579iOh4s2+/Ou29VlFUV5zrKbEoPw/QK/lQGyuKERIsneSJev6+ENLYLt4mKEZFrxo/Ikezbdm
6/Wh/nZz8jDfralaLxrxlVCq/rYk7/WULVfmFRixlumuE7gNKMwYwZtyXUVPilVos4UhhKxffRAs
pC5rPQryaZOqY9N0AVwGKx58tZBYcQBcJp2pGik66bPDQTBLSxU1TBpJftruLWpBQzq+mI7nJYZn
e2WAHxbN1zz3B0zk0sKNpX5dDadM2m/xTNDPu7bKo3ml3C1EzUP9uKnHY/5j37IKfeN2xKoUxxht
3bWZ6N34/BSYVOgjFuUg77SZgh9CdeWADyEfakA9o+8FzNTYgEsiK4Zh4D5dKFLLeRWHsz3xXLZY
XP8s1Bx+eV+Q1o8CLpCEMTUgq9pBaITJsBGhFYk408bkeqDx999/N6RMXM/YK3IdzqGgCuZCCVLI
UCsvRfDHU1VB1VkaUMdRjpLXLJoEUk9bpCFuPJg06b5k6sv/CwGiJCp/I3z4fwtq6Qv3M0c2Mvw5
0Iq0nQfJHddpBW6+YZ5tiljr/nD5vgF4N8jwmFDyWx8K7ZQgtZKLlEBt8d7xnhMbn7+f2WFzuRTW
hCV4QIbALhM1jNEy92u4FIM14hcVdyyQbHDYQH2YGXpCD0GhhmjboZxSciV2077/fG7kiu/o6eqX
3fwVaPPQWnYLhZ5JIyZqc4VQOwIm+4NcwDhSrpQXGVOLTMPPGz+xa+ZWIqi+HxzIfYLz4pD4otfI
O6/UL94/fOFjuABiaYNFXGSc/BEEX04kO+KkuUJ+2BUoKkwhGl0IhKlfDA57X4JgnomfIMK+Tv/s
ZjQNIXp9OKP67WUOEETgR4MHxCIf9zyIbc1t+LOYrrW3znA8HS6XLgayDHDFbfBz3Ph+kGViMHsO
hoLClFmFBj31dGJenMLHUg3yd9e/mUs79Dp/6JV2M831o5rq30DR5J/igB9QvmbZkkeQ1R4upmQx
2vFgIFqtv8XQO6WsjsHtcjZCnDsgOsmWYrxOLeP0JdJ74SbVzDeNg7hlzyfOANZVyo4emGqbiD5Q
GPrfA6z2N5MxClob6tNRMKP1Hhg7XnfeAZAemu3agqNtaQ9+FM7qhG/kXfOApDBQ78bP4I1P9jIm
yEEtq1H9tjGoTGXEXuGfzSxHN8eg9xfTD5qWzDPPLTgM/Fn9zfh65wuimoFGIRHoxmssDtcWM5Ov
f+pRz9aOXtwHWqb8b9ftC6tvS+OiIbP2reRsFjzm5wiGqx2sHb3vNqzui1V/l/qapAMhB8T7uXG7
lLqEdFx55vojfnnVSQcANYj5xksJvArFLLQgFSx+TbdxvH0V2Q9nxltWufOY67m8CzAJGjJsKGhZ
P2Hth97K+eLs3uBh4iXGgybNYpyUKwUnS1VUkI1hZRnvG0Nr+P7PCc8eSUbSxRretKWztgYXVgs6
IPyZZg0YXUA6v8TM9wn8TnGXd6nOjCOnS/54xixsk55Bri4uFTlMhzjFbR2RRSToaITyVbpgFl/p
Errz8bqtaBAh8iJB6TK1QxWZpvUbV2HmRbGcFbmlnnTlGupzCkzoKQ7gwY4o5fevk4gu02AC4QD+
eyz0YRJABc4Ff8QU+KDEHwrjIkelsPoSbqmup+rIUbH7YSJ0HfpEGVgbpYIYei6Iyfr6NvOwG48g
JHm/sR3f9+CkBaq1Wi8lQLlXV862RnYJkRTVe4YE7IGsNGev2cj3OrHgAhAGztthNtbjB5H/g1+P
GzbYvRLW2CadLuLsQGY39hN3+abrhBr1FjBU/6FxEk4JTcoYVtQmnhh/YnmXs3rkNhWnKjUsBszO
LBEaAqRdfJCx7QnOgTIZbzWQOTglrA+pN4wCW8+qB4BD7besuo6mmGMsDiUnTCDhmCxyHCaw/YX1
t/YO7/3+rtLFAAdSLLK3o8Nhw3gPNzkN4hsGg0FxiDYh/1RcTutZYs+slyQFjkguWcF+3v1f4USC
wC9sMhPSjnp/sm4/U/ayL/sNbJlelB795BeCwN2fRyBOrCSaN9/3B3YEvxyQTXqdP1E6oRSf6721
jeuddtYIvN3RnEItA7n2D1RvT1bDaqtQqHUwUpcAnXgQQqwx8kyQl2hE1FBWeKebc7Ilr5FIN+nP
BW3lznuNCITZd8XRJQw0qjL56NufktHlPyWq7AhkYJPmCFeOGZyU/CpwACkzRHZSzT3kViylyjH+
d1hmUQt9O58Qm7qBpTbS1i2ll1pYPytmv+CScFl1sQ5tYK4TqfcSpzTZduPCDA9lmdJESZre9oQc
yiRJq05CSZ8OBX2DVXKTjFTUX3Rk7mA8UAxmDwypo+eKSMw6mckWIeMaGBuYavToxnIibGyZZMW1
3xssv2GHQ+oZsNSaqp7OX72xDS/21oJKv4/mBEurbqdaim2lXmJGBhNunb/O7FeEGDbF8X/orrI3
w2IClkY9hDOMgmFDz2TT3zTQixvhVu3Rm5vaGUBOoPmkv3jznDtJvA/LlFbgE0iPaz/+A0RFVXG+
+5eY5GvpObgYetVQr2d/RmPdJ4BL4yi4LIf4iJmDxWIvOr7oppDW1ZOsk+b2FBQYYtT1Qad98JlC
gxVKWEa7yPDkB/Kuw5E422sqzMDfMXskW5cbFL23gJoQ58V3yuef00o1f1gA7FcOpsrSVME2opMI
Sl08AJO5EhqEtrxIFUBbAZ2fG4edob0zR3ZHpeEewK5t9HOrHJTTm4vAYKoquQkKpSy1YPmwKHfk
NnzkM6M9eogZ3kDJGYrSiN2vFr88pjz0reoIzs+hkWZb8wbIxAGyuF86ePcso6qV5oM8XE+21un1
stZ1I7+k9vEh20Hoaxqxc2ASomVZqx7L8xZO0SMQDQausD9Q8bNfh5Vg0+iYg02nTLrEd8ZPNF0A
CApoowa+qqARbMovpIU0E9D/6KRZhjUzbmUJrFbUGIIoqvS6tItpGnnskOWZkoPn+5C0jlmRH65j
F+bx53e6uslkUibVSMpDJ33IiHovnH+AB91C7KPxEi3H/O5/cneIGtmRjtsq0DXAitIhc6Eomhe0
Y7mEF+TNshR26kyr3W429Qpn73zJyynXAtnZWZD6ffksMigP0BFdL5cCkn9i1YXYDMRWspu2RWQ6
k1y4zIRrljH/BjQ/22HOLApKLW3s2yNuPOT5gvhYtQZUDrk21evlZpuM5O1Vuzy0CYacR0PJzORG
YryvOFHpVNGhlyzauyqoryyZvisKKycc2GAcdG1mw0n0R/7KoWmD+TU1ZcjTAGr46rxa1pd3lhDc
wMoCaxacMpy8nPzV5jrYai1d9aUIxT/MV45LxK+jXby/o1Suc7QgT/G7+8gW7iw0MeS8JDqheT0W
qSVfXkzHSRdAfGcbEtKji03zFxYWuayeRsFMiCs4ft66CS2UuQRMiM+EHAgRhmyY1TaKxFC+in3C
UUirpDTdrK8rE1tQSLqfSnvIEM6CBdIl/9MqlTpc8A+jK+qYkIAxUINLGltcm7SWZIVRTvqm55Ny
z6/O7KvOXgBuH1vLDEQU3Lrt9ZAdGVaHkK3TmgGmmfOpvqLngJ/NjFFbX4m9VVP0VUfVjN1qOP3R
ky78H9iPBrnGGeB5mcpZJiN6M//+xtnmMMUMOYV9mR+8baukmCuJCtKSWnFeGBHF+nsrqmPIzdbw
vTWjnD3CETb23NuTaoYkblXMmfDzj2YmsCgv5bBQ1ZlAyUFlTa17BGgyizHYAAstWFrHj4+755EG
oMkXVf64n/8+AidiI2X2tHvLMmMtTHn2kjbTeXeUzSSFr5c4orbRmXRR9//tWaKIHoRq7BeUKLV1
wWjFkXAB8WKGyuZIgtIacFuqflsrKkmlXUELpohyslyhm73LD153lq3bWUN9CAxiIsBlnxydedMs
5MSrJ6WcocF2WENkVQ1zBb8S67a/iM4NxzIljh0n/lTAjKCBnoCmfAAGX06unrfwxSIZ1YaIu12w
8iz0TuTCyqjddUR33oAwLNFv3uEnnvqFrWQAGYstYyAbwVYPU9KNtnRvSI6k0Ifc4sPZaWXhMLOS
Y6EdUzkxFV4dDT4qOlkpJlGWoovpLoew7zdO9WCwW7r/EyJvOUZo69QZE7QaWRRxAkNQwE64TLFp
0FnewkTPHKugwpguwflaQ2rd/oeVq9dX0vHAQhOTCsye+eoqLZs+nhX2C1/nfo1Ti+P3K/GsFtfL
TY8b3vnHSFH+92Dr22HoKQwNiOWdd8e0cfPu8uHQfQggUbOj9wuDewWJgSmOOBPEaAdHqwNvkp/i
SUmSzeWsgmINmRTkEM616KaJMRjvLd81oR95Cc1jSdQpWmCW3Qli5ATnXQcZqHnctHv9JvwTVqAn
1UW9uQhzeB4ke7nMlKkY3j4BALvleLMTt3lCeemyZHvqjKUIT5dthTx3H03zfva4qBvWOhhekFOT
lGMxVRnjl/sAkb9SRurOFgePhGZEkDSEvX1Tan3WFbm72sHrsj8pAcPw0ztJRDwlD/N+zJD+Jx46
jlU/6pzBxfVHu0it5Il1HiRywO8oIDF68caxcd1V5LcSXvt0SEOvd8gj53L/sQXfWESIGm9+sOE6
4Gnmln26DTBRftudZFLkoLTPdOdA1umCEOoXTS64zXplUA1V01xJdPe92zX3nY72PcSuUTnToeC0
bf8vw8A831PCg71ENE8mt94fwcQGKZT7AqrUHLNvGc4tptCA2w2RnwoWCgmO5bKQDBl/fnnhAy5m
7CKvzRPn8+6dCPfM7wEsf4WYYbXmpPEe8SJbC6R+Fuy4QYnNRKMaMkJu8Q3rGbp3/LDN6t1fx3ho
pyoyXq1HlcKe9vFJlfTmmJa+AVEv3TOwPUhyzhdFDKPauT64/KMMmcloxIl7iPN3dlivYFAWzXDv
/OAk+H84Y6NK1AdkrQ323jVD3wreJ34fs7CX42RKvRgL7xG9tfD1NhbKDtPOyxokTGuETR6ziP6F
eVdrDwUlJG1WCNei4v8lUejxxJuOirm/yL11B4vHmSXjvnsBhnTe13hG7/SkarjgCAdyq2XTjMXF
Z1OgSVnL8HIZscIboThK2NJ6qadyb/x8WwOK5wZvruR/LukaZl6Q8sspwrm6NUnbXNxbTWO8tXgZ
BkdP6lDh/pW5KnW0/yaKV8dzRN0MulSY2qEPhiXlS7+gCxTivBk0mYRSgBCrPudAMpPJMfft5ThP
PZTQdZ6FylFlUrwV/L3jcr0+HG/FUrWkfnFFYuBI4mj+gkuR1x0FHGethMhf1VjIrSHAXDkflFsQ
WXiNd78v/r8ZEy7I7MSRiS6LvnJw1D/uE+HuclE/Cu5i0+OtpQT/li3u6aaG5pKBo0h6Pdm8Cyed
Xva7hJ1h/o2DM6c6pu8p6KmBF9fkHG0hUy/nF1Pa+pX0gbvKB9eQpw0n2vdJ+gQiI5BBIUcNs/lq
4YB/tu6b1RLvOSXSsReEp716IPo1HbNudNgo+3liZeG/90RG8v1aRmbE/w2T8Xg918/JuJGzOG2v
HjxIrNMV0O+zl6ce7gd9bWr3O9bb3k0rMWbqoG/O4KyG4Ea6GXyL6wZbRoqnlf+j4r+C9Oym3oQq
b10ctfEQOD0Lo3AsSRu1EK6rjbpEH/ll5DwDwMKFto8MQy+d68U77ChV8ePRvwockWu8thYL1wPP
fQwzR3u/ApEuL0UZyINo/jKbxp9MRmUQRVYZdsiDaS+8XZjP92go5xr9tTXsw3r4snQa6pxVGv+J
O6rifxLxVQS4YfyMSEQvAOboaXRpVYhHDayFFaLQd7DkPWYqbzGHmGzzHBr62d4BlzbNsTmndvIP
t+NcQwK8Uj0fszfMQoU85orhoPCmk7aLsr+m7Gp9FcCkBZ0KSkra152nRShazOA9X10iL1UHetVE
sKgD06TeisSTeKHV7XAm3GTYwyhQBs0UrgXkoBIwM/qb2tN3EA0I8Fajec1a03MrSmVhoYaXQ/ea
eswLgJap48Qs+7kaOeK7GKWYRriMDzun8y8txf+Ds934iaXMDUdeoIf3fdQOZRA/VF8LeGTD3Wih
O39koGzT8C3ajytwVMj9qQYLEDcgGivXboZhVobRTaIyd9GjsiM/BB54z/TGckP6vDaxCy4vHp43
DcSMYSvji/C6tPQSKFnc+Y1FH353Nc9VWDESXWf9oEfiwsENSMkO2JQrwwPJWiD7bqzWTKSGk5Sp
QqoMF1inzAAUUJ4F2vvCNKeuwNHIzCZQn1FZsAmyTBIAs6GzxmfLM6THNLWRBZ2Ih7nvp4Kf3WW9
FhNOGlT4yfTpyoBPU8ay+TEObQRHSK5TqDpUGqUadv1h2W2j6lw6lvm+nvDHdHSjpPrdR4OYTwx5
TBhK1ggkrgx6BAk36Jj+xStVbdXor6JuFoO8xmjIkCndgOfRSNWHsre1q2Dns2V2iJZ4A4iwJz1v
fVdy8AI3omJ8sWUi+fZn0mE/zkgL6tQw0vIMxV6o53/5Zj0XO2xidXkkTfi7pC7BCBM+9dWehy9V
NQ8qbTS3msWgPWPUY2i/p0tPckJj28ZS5d53Oae2DXD1+6j5aK3vaeeVcTjjmR07NB6xWtn+xsTV
joOK8j7NtVp/udfKgQkgkByuR0GabX1G3/n1VsBuJuvi34uJlfuz1M588m62f8eU5uXk/lnZ9yUj
6w2OOfEyTFC2Y3gMB86J1JhDHqx0Adcw/yfxCXutpDp6KTTTX03dNCeRk6Jn0y2mv2/DaBlDmtAj
Qs9aUfFyHNaTHFMdGSUeMrNlOUGZNgYlUAIlnOPDYTWeF2AScDGb8pQW057VhYgy+k2hd+vlh70c
rPS0smoiys8aETQ1fE7Anbm1Rud4Jg482gbqU3b8hQgksv+GlBfw62XbZU+GjfTVgpmn86NaT9sl
j2gbDo8Tl7pr/11cEPAUr9ImwmYv8M87iFXo6Lb7VRCUvJR0jpS9ZON3rbhhsuXabnGqDEVQ/fvO
uCBBnIwBSWktSPl/Ah3+HzotAt+vaBawbGxDURf+cecPTSTHwD575tRCjT0bbfgbBiebOI2/4p1f
HT4naOBjW7ituvaakYPV1SCN+gOHjjt1dO5YMKuShCh3q12ff9Yvh9pAG1TipUFB3m+UGvBwTm43
JGxTaGZe2LhV9+6e6M6oZcY5+sMoBZl+kwwxYKjIfaNrCtpV2IsrOdOJv716imurByAuOwq8ykL2
E4WljluLDQJrPKlpz/wfUUEoS/pGfUIaMnHDQ4EtN4IEVAqnVdWfBrCoLodyHMZjuQ6t0aZ4lMpx
ZcTYfy3x7P8X8DVV+rtdMaeikNdkmY3/vFmLvEH69ExHjXYkNJuY4WSwBIO0hPW0GaIlwA1AA0g4
U9znVGACpO77ALykTnN3WOpvwPnq5cpSUP4gVhfdCq0LoYY8mCraX3YdJ4UaJHCugdYhpQfBmnaQ
IRLGeRh1YS1Cgl/pPTu78YHA41b77Fxwysjx/PnElR4u8Ja/s/TnPack4pASPvgBUUzTCWWYVIWs
oIEJ1vnyR514jJgfoGGdDa9MKSv4qKP8agACJS3plrmZTm4ifU34SZMyw9J+3+UIAkYmoI0ioVaG
dtwmtWRXLqQCkATC/PevWoImszxx4M5uVRgcrnlCXsSpnGYgk42erHwdPolxwcxBBU3ZbrGVMOUF
JfyJYegr3VASJqubYcQu2MZkyENfwALDSdIxw92kouH68HTZFouwOA8tpH37RshkGkvoRR2i0c4V
gSGRNity4/H+G6L0I5HUlyOg2/wtDD9hzAQKY4lNhnbqvyh8erjD0fmx64HOsCafV5/MFkpXPk4M
SBaIv0MOwcBeVmp6UBgob/d1GE+70KGfwil8tAuN1ZvckKtKq6W7pVv+5Vw+9uCMfl2DqfrFBP4Y
eXsJTer1IPEZweP8dKf2okMIZCQ3mmwcrPjuPJKxT2hGp2BX6j7gZyNwnE+rkdQIjesBaYwbDAAb
pGXDMu26dAKyD3Svlm+ini1Ge//drMIOJly6KELu4eCKm3s41osasvp69Qr9RfUD3lMHwZIkxmZ/
03tOTRgiROA7hlYnkFjYXb1ayP75Ig4HNyXoIvULMHZfZ+zwJuvaZZ6d3KH1TMFwrKugeg/ITkhM
+QCi7Sv6AjT5DMFgt6RUNGhYl7y4vUinESkpUswfH1E7VXeYKkAnp6GwdbK5GQdTivBhzArf8XiU
nz7ZE03UncKvz/xpP8FokKeSIIgKXrH2ta5HkNxu/+qwZ5XbaLKeRgKhWv0ogmXUOYFiMKvkGFlK
oqwCYPNeR5NZg6TTqB6lcPOANm1tkiFYfhl7hLPnsYY4aD3E4b3KRBF+BaOqeYlE+PPwI3JwibSf
0u+8pUY3StX1Qsmyg8V7TNK5D/PTJC0xv0sw5YX/m1yfHcYTP25ZgaMHmvSRTSLzqoAai8SvvZS8
miaTiotr4MrIIxdedDyVJ3HiX04+gvaz3CZYaIuF71mqNRAPatJ3rubYpcpHNOvCGQZLktiwiM98
LnumqX0nQrCyQRUh8HvYKg73jZECtAQ2QuqyoH31/vhSxfx2Eme2n0u/Gnnbf1qMiiHdpBf27bBw
vteAL3vRiMoPnU/NQ0L9uk3sIAx37zeeP6GECX3CDN4Ln6yG1EL8lY6Vh1twqx2GadOSeHxXM9Kj
RSKMXA02ygOHL/S064y11OKAUDNJU8GJmtSgvM3X0bmuZyHsTbGdW/MadsBAroaZj99GvlCenD5Z
sFzcU96Z59B1OjR9oKHXafLybH9zkm0ku7TPEVED/B2MRGeOwApNP8fPLPDQAsUI/+7/YYsSJWVn
6CYlDmNT37YEo9bC/p3N5QnOABa7ciOTTCnTcixDIH5GNK0KYjqSIvgCrzX6t5u9b7xiwK8hJN+Y
xMQ6kx/saWBE1d1kgD/NqI+p7Dqe2OWjwCTfXkDIVxxIm/OoCL5L5nuqC8n3CdbBu9rzalKyKCL5
tnSAwc3gtKUP1tPoibKzH+teHeRDwaSYW5S3vCyvnTM6EnLNmSufwsM3+hl8yDhNeSiOyTe30cyP
o66Pa65yd0iWLASlnzk6tGi3/CCuDjHzLXu9rEXf2iCbAg5dC/gGZGvz4f2gs98QQ9Sdcyny1YZf
YyZ+zZDdsSXmV3/UZlddoAgJQ0EOXljblLVZFpJLwmiD+fGsLzJQwSL46s1H+jACQQw1N2W9h39A
W66hZtLrvFLFCWjqes6Nmb+lAi6pN6xneofQOFM8SrA+6xbM+xSzhDhMBLAIL7Cw7NaHOkBmOK58
5fIrYMPh9Hu0MH3d2aO8XTacMFZFk52g7h9HVi5o8QOblkR6VVHzE81fF89lpNHeKqzYjU1YG+js
fnUK3dNItQbOHFhXKmJaPqpk7nCOpfa45CEfNklfLabeA8CfGtCz5P9iQQ6+T4YduH2VcPjXcvre
WOb9/Ys3vjIf13qDXbrHETfYvMwspiyQnQOgXnYAQFCk2QyJLvAEokGekF4xYn23roGPZpzfaAMu
zjpmIurc8bhRkxEdlOqB4RTWlY2ZbGOWXCyhG5pWV0BUsnPjEG6Acr8M5lIA/32qraguDfmoqCRC
of6ZoPzpu29UEeO0slOm6rjUNijEtw6Udq5f7OSq1RzlhfQ7HR1DZ4St6oj0hTk/xboLnUmI188g
3R+iXMXM5lOHGZb8L3n06TTHZHz4mjU2p3ftHabEEd2HVrGrV9UYXxRDJuPd5h3qd643Vn3Bej9g
5hsUNUZ0ZSwyOJcXr62hnyIUzTC8pWw11qzRuoaqCXe6IA0RIrpdll7pn4p3fvZXPmEc1gFKnKdt
vGTDLnDwRe3zQpK7sGRhwsYtB/6wx7d+8F7Jg+upnZnK4o7N3IgRZhXGWP+CBjiGCEvCcWdWP2XU
jj+yOMdVMfH6QFMwEKzMAdbYqPY3tdg5V+4sDcu7P8gKEtk23mlfAopVAGcFVytUE21cO2zhueD2
OsVCo92VtvNvi8ARLahFmz2b5TWvG4v1fitJD+NdSE9oJp/L4zwpoZnOkfzr8hQvnfZgoBwIK3ZZ
C1IDsG9fsKdeF92a9vBWI/dsOJm9HhsLYyRVWjWsasA6DaPo95dNAAVvEPGxeAcmr9s2/9NiJKw8
t6fEt8x5zUcSHahbtTcrsO7u8L65mhI2bHTOLnAQNAjoiplRB7eMxs7m7X8qDjkioZ+sqNy3Nqry
sBNJs1R29nVzwH60PXUKM8yoWlgt4w/cEcsKSWLiW8f+wN8gmihjTgomAAiS8WhVm9YzexJfLHNp
Aee/yNNFuVpz/uS5oQZp+2wplhqTwPCfeAAEmLX5uWboHROWRAVR96OJQ4fPLzwAadIKJ9J5SmfP
oK9XeODTDk6ABHdtYDM+TjMn/vGjio3x2wT9GtuPom87+lvFSNioxYuZ4kt2Ml8hNaKAfG3wl6Dn
l5jtVS3Tl8plsC4uK8ekSiP7Leh5jK1O3Hkj3Zx7P3+tw/QQY/5ZNy2PivIQ0fY3OlcP30T0yt3l
s+cj2jvyUtuD6G8VmVjfbRF1fEkc/gcTr9joZc64JQYku0MbE8gFQSUInYYXMVwku4p9NiWP+H1+
xOt7nHQRLffumAMx3KF4snU1xb6XVqllmR0FxJ7ESRYgdEe5iH6VJg11bGVNZHe+o3c+FevgD5EI
m8sNQj0noV5V1HTQOQ9J2hZ92pJ6BVknZbydrRASy7HES2mbgkCRkR8+aheDJqjgTEMS+sMOG5Bj
jlIt+L8teSFj5rUspzBFSDqt9ko2RLRqvKvVhmNnZ9ZTh0o+kcYQKQkaiOKrIfjYx5vYN3h7hcpe
6BAQeF9iniUdHQ+FFTpKVI3XO1/VF5Mmicc7LGHtiweK7c5ygLTVp0HdzQqhLLkKNFrpwg+ao4vY
ZYzeCcnWp2pYE1rVufd2HhgLpVIyZ8c/zQ5O1kKvb+o9IoAZvn92gkeII8Pfjt69R1Ea3fnNECny
muQTZeBGXjuBruM4tJ9gf0Fsn+Y4b4GBsaDXVcVWz56asjfgso85i9FmyQjS/2CcQmHuhB0dAUwe
p4ZjACnrIsoBygGPgKQTKcWvJFVzr3bzbNUOiJnlwGuzihODRscID+VKLP8tTFdE1zmSeI28Vxml
d7PmDcmHe2/dSJOIh0xHfEr8jw/ZiMDa5ieNwfVvkBZs3xTBSW4U7BO9pCcyi0o43cm9DCigW4VG
Q6679qaO2Hxwyx+c86dBQX8UEo2IpTx81yEoLg1K1em6+seoqBEv/k2yKx3kc48WPgNbt1FBiOYy
FQ6f8kIoJXtWni59x1TSHcgwJ83H9sTssm9zvVVXYaYO99bl2XjMwHmw4+WwANpDWtHcyrFkjWe3
tr5MAx5QfxybKh+4ACLYC4tdvGSKacZvHjE5W/N8JbsCGfjkhbRlV8Gt97rks2RDipNvRAlXoaI8
DpSgfp3Zx3meokvCL30LhOvBCZzefdRL8B+snNCI16knETOUbSb8QiNGGawhEhtOQRL6stPBPwIZ
VnPDHMToIGO0wvRJomgP3lWZhHR+C5xiDfiFQChLukI2oAuE0D+GDZ97bZ1E7e/ta6LeQS6E4QYB
KFf7lAT3gfi/bmL8dhkvSrZs4WvqS8WyFGLPgnNt9bWexaPjsh5A4Hoju8qiKIsZIaImxJU/M4q8
KReIAfPjdQyhQzT3k/HQQ9N0/931X6p0NJcBpGT2oikM5vgjTxArNLXJV65RaU1KWblsO6QB5c9f
W93CkMN+Sf5mz/EaPxSFn9RdvbVaewODFz/aVY1HRphoBSy4hsaXbOgUYezRPQdS6jgkYmqu7rzu
/p9kyhqpvgv0VhGkw45mBGZkZbUT85vnQ4AW0HCJghj5rWcGxJB6sjZpuXnY0YNJwUY7gaE6/SB6
4uBAioU2VcbjoNy8A4Qs288BCaowx9lzExJw0A6UHMgoe3ykr5xn19UpkMVFZzj8dhswp6yEACey
hOzMT4JaTqRH2tX6LuEH8Zt3IDvIPm0VFZ7cd5X9HHXoWAIXbHL0sHb6AaNkAiiD48p9yfkZcE82
Y3KFfbdQXTj6MWnjUBANGid+SlBXEf67iRPUfWfCbbv88o5ULsInEiVtXTam0X8/VnF6U9+LaPJk
Md5XKQHK2K812JYFYuOQz3Blqcen4KMb416EXT5o5YCD5+dIkhxgcSlLVShP6VJqu8Pi4XxNd3us
OlUsKZbZkZ7KT3Fvqgqca+cEvMHmt7RiYFEHqPBuP3xmocBiwwWo5ctGdSphgNSLrftzGg8fvyj2
9ecWkExAEiZFXbXi9KddalZoAcFc3+CDJ8ZvaC4coqNvEQpHTy6FO7Ktt3KYRbkQsOPmzZORplVd
/DbuZvlNtU+NdJYPAwaH2VU/E4JAbun6KueCszwLh3REHHxnZvs1bWZj9u2s2X7ei4oOTKp7hy0u
P0cltdxg2b9yBHQXwyttNF8wKfjcuzJVMzQgTeRAvZ+SPitn5kpNLBCWmvrzaZfmIMcvxPq3msqn
I6YX0u2bI6sHP6dAYpCfq18p9t2hmPuE2VwSKDkt6fd4JiT1EBrPTM8ZU9Y6yVLO2gLWAZpTpMlo
0qhalf8WkAhcQsKXUxZflW4oOwqjPpDK55uJaYscOe+HD0xjhiLPzjEyX4tRRY14EqZWHEJLaj4G
xnrp6Q+QgE28X/s72GsGmrDnfonkPw99qnceXhXfGORkBJQcSLBmHBTaZO8bNq/rjugeNbMwMfuc
ZAYjoG+wsrHSECS7TOVFfL6YTN9N2yMiIzQAmbgtmpBkFQS+gGSJ2LvOn2YNnvRPv/n7GR0SrswT
ZIilHUJi2uj/wZY511E33h8YUwPsGkB9ONlbHRj9L+xUz2M0jgTb44MqEo7/qiEQnSincFYPJOzi
lqCD4hNUR/1O9PDmxEBRWBASWVQ27pAefLlCuoHkzTJIdtcWage9gvmtaDblKcYmwOu5IK4WQOjq
KmXwYnsYgi1LZSp++q6gU3Fxn6xULNsAHaZikZ91aE8W7XD0nZZOGYeg5i1dnTwKn2Su6feic6MW
NBYUqZGTtOaAPdT4AQAgQAuJUQYJnl9dglPcg2sCDtPsnPLbMHqJqQJu1MX/I3PErqRzBCU/skEJ
Gj5nDLXCvKw6eAniT06kTBzgv/9Hce7v9bRpIVUPdtRTHrbeGXC4GLp3B6VCuP1upW/1gJrVdwh1
tz6+ONuJ2uVtGVAxjgM8dMAaPu8ac1Fc1+6m/zphxm9NED3T84Y4twMCgvZUiGtVzG1RbKLhjFfE
BWbKo11tl5TOH+JRcY1mf3tf+zQB3C42Aszo1FlEm0pKcEXWPqat37DAGnf1kzWCz7hZXzLzY0n7
PiUr4MhzHYf32VwUnWidgJ+AQu/IuFQG10cDIpuBEMkIaUCqWLR4bhaDryJPmPBpTG/w31GorGoQ
lVizIFrOK3C7TYwnP1ZYxfsyTM7Z/DqJU030/H3vVgADrmCrmYyEDeTFtpecDvEI8Us0LDUKQNzm
Gc5o3WIPJHGW8d+GGKEM/qsoRprZXZZkwV6SZcLYiBZc9tkkbuF4fwaopCVguDymB6iJ/hgSkjnS
Ijt/+RE2awN8KVbv33Ef1EFvTW+AQLypd5jNRrUUIWDtzdYTn/QmrsFhnMrGSWqeENxiKCcBcsTY
WAuD4wqEmFZY8fqueCU+3EBUexwyJ1juzcSowWrzQM1y3jLY3Ih52pGBrsEj62BAJo2A9QfWxoqE
uv1hl5dbdeN/sPV0XEDgrylJnwauvyBrg2x2q12TF+CshvEbGUjwfFO/5j44vv49mcTnmvJX7D6w
aAZhJtie4/rVUdACG+IPxN2Yknw3s8rFF6YzUUoNA+e6vBfvh/R7UhFBPp9O12tTSRdO3MrfisyH
oAvayKSccD67FKq0ERRz14VYBgMUjRiuORFum8N8xf8r853/3vTC+iwtcUX6QiTgnK0BCP6dU970
rJgdJgtm1TD1Ox9bwVfDhMQ+0jAeC9u+Xj5d1u7uWjDwF8IjQnr4Xw2Qx0q16EJ9AWCyzDQ93sML
xfPGCsEWzF6qe8ydvW0gkIGTHbMfd2tyKAfEypMd04IBHJEDNnjEnad0QyOFn4SM2PhnI4VSEiYO
tTPEKlYU/mX7MHWYudTgU8UgRqwVAS+UvfXv1dTMRkbVbTxeaJtRAfr+YxHzqiBi/Hp38GFyqLpQ
gqb0eu7WXXsRwiZW9r8XyvlswT9pi0FXZLNqt+9BdK0m+ahulnfM8HbxTUV6nGHWQcygOL8IdsJO
q8swcRNr8nphblaVlTkTfdSdD0ZTxKz7l12tgoLb5sYNOZki+tcL/LrQEeBXc5fb/+YXl8MkYyNS
oKHqx0lYiU7WPajiBDSmei8biC68fK9QKoLXdLj5/SPaCM56Jb5GsegYW1c0qNMCUowmGF5sJ4AO
mXAiWIegVN8t2ftyQd9pE/r7HC5VsxWvu4Tun6BEF+rBzHsNUIvS+jFlssu3AxhUyfnB2BOgRIEM
ySSoJ6Sj2DKv0tS0oLpKI+OTPIcdJJCv6XFbsUtEe9ZGUWe8HjNiqEENaiY8k7YYtfKcRNTN1dbw
WLt/zUgnsTfxgFFsAXG67zlpcXK5nL+B8GYGu14mzwsFy4eWk4xzNBnBtvvUQZHLRYXFxqLAWEed
EflZzNcBjC4UAwTzaIKVKlua57nxd44Qd4bYLFyghJeI6Rc0tqbF0U50vjxCOvfZiQU2oh1HOxoG
Ign5X/ZTb8GBE7JsKRkgYiFBBLnDCMNVNmQDQU+BA6Gv/HoAAmoWPKa8taU0+CSlW7jPB0hThmjr
RmBQNxPHeJ32Dp0Z+A+/UknQiQRRrCBcHz0eJKi3QHYpqBZivZNKX4ggICAf6dUkB/VygE43t2/1
Wxf87wxp38HTJQods7SLMgBNrt5cQy868Xb2PK3p+a2+vHEyVk8V7kMb2fFU8ioQ63HzY3ly33qD
mu9n9x3kUlKvXUeMSckzyMkwf3IIWS39nIYyyWuDsqABHyOZayFK/tGvEIFdZ3f7JMOfFAX/em1f
z9hY2zhAvesE86JgRN1QGsd+vibnNV0m/0Mng4XZS14RKEUEN4qiq/k9DNTelV86nmWqk/iluVRR
ag0lEANLl4lqMCkY2vcc3eb/ZYAqItp2gg+Iq+xCttoFv3usnhEGQJmyE49n5kXKVwrsrvoa3oe2
EMTrdXlKIBZa1Pku40cH4g1c5OwuwQ++Zl0ZZYnhiZLPWOqyUlx58OzyD0W14F2RR7Bx8S8mtkvh
ys5uPCbn63Gdt03tMJh3pkvI5hQ+7OiPvGj/AMnuoA17qiIDl87dLWG2zrGcoKPv+qOrT2utJN4B
70PNmHWyeZmixccULhnMAj+9t1CThAIJLd3KMuenqafmje5DEryIhsQ3apMAEwRQxYEzM85vyfB5
rUyZQixM5DdIhLNOdiLb1RfarZcM/fR4YBpyFnJ4FlQ0LXzfXfkmETKFEEUVbn03KyOv3v13yEwL
5cHft6Nk2i/yh5uJkDknh9r8gYt/gpM9Gp3lIHAusWmlgfPpI5CmMe/hmEgW9rOjn/dKA+8Pj8RD
is6wMS5VRLfUJfJEmRTU0tyh1GmI38S/0Tk8HCB2H7vw12fu1o91CabiaET9RgADlE7l+6dyvuos
tIhzn3G4wP/6fxWS1B9ONNoCv6AyTWvJyZ099i9/XfiXr7yLC92++FfymMK4bGtW9nMbyyFT2iM9
yg19eRH7OdidaTZUiHo07RCMzWYjFoyZCAIqhJAB8leVbX+FtKsWVaWrBItnO+Wn1wxRlCNvYZCT
DB0fERS+nJhoAvjNjO49uY7nq+lnGwdBKdNBuAZ7L3x4wpNplqNAGcEMycG/ZNbtljF5/3KsaKRr
Vbp66VZV1sPV9fgDwMjZyPXd4GpO763ry/mbR+8x5yUOFiipttGAyq90o06wNoDbnHmkzykc4Y/e
0MT/H6npeK1fLqB3mG3KuiiktFobBgY2YCLnd7LHOcGz+nVDEl0IfAM58Tt7sY/JZ4rj1eSk8QAu
1YJ38YXQtGwMIqyr/fEssZAzcEzw4MuXCEkHpN/zYByxttdJDYFmcPx1HXQvO25TUnYVoRS9sz2c
FMQwJElDE5LKcViiCaFBl9163eDwZfV/yXCDgsQR+0RiAcAMIwmQCLUiRjf/z4INjM6YHeeD6il8
2tsppHVZ/3rzcHaq/WXLAHKbVQetINjO9HyW5vrxA7W0EhfMtzVaXwrx4NwbXVB+0BnvEfrlCWIo
aKIjTgOc6x3aHhPTDb/gx8pR5W5/T0L4IAJua1+e5VFEhwetRQhPkuhr8rShqOj4HOdQXKwpvlUI
ickzNEu1t0Y6OCbNRuCp7z9kimPg1tiH774i0HhOjwhOuZNkBu7pdY5Pzdb3N/ARtD9Eqxe6iaOv
LwvGVYGN2mZiD5PzNgP8bSf90ASFYlZ/fqqWT57QxLtYa4WOPkudzzxaMZzdfMZAup4afvtZq/ke
CBWgHdp73hlXXBJengtDVcU+JomGQ4uMJ6UJG8tk5Py6LE+fz0r+1YGzvKqPR5eSzdcYL4ETkZEP
XNFsaFYWjtxnmkwWxCYHz7f+GZsv75+nahfKlaSXe5fKrakDa2xpJkaw+eDqHMDuVSuoiwSSTS0g
Ukj7AhhhxC6rfNGFJPZHMDcu+VPwC2bTUrncTRKlV02n86CI13GcDxFgUeqCCcutodWjfarM9ZQ7
gYnIX2JC1w38r8A/yJQIgbEGHlSMnkmIu3iC9FzD3m4UVuLrVqYz8J0q1+lZTOlIC3/SMn3QB0NI
ArPifoVBIOjabXIZ/xrxbmVdRxoPotwdMyLPvdqm9sW5/DWff5zMfrgg37rbfMg35kV7htCIB4bq
D0A6lgo2+xFmUHew6stwRUmGe/XW+GL2iWnz/HI7/1I/kG6cAv4wN8wLc5PBUWqNzRmqKEK515kb
kqF66w7rk1ZOPgbQq7JzPQzCiEk3lGp8FHYpTejAoVJbMShvTg1L7Zou8wZ5Nuu/XsHlUVxPURPd
tA4YCDEi4UMGge4BIuiAmTGnnguL2vGyZE9iMTQUjnbKeakowcz74EDsVHxy4GTlIt3ueoCLqtkZ
/8+aAAf4mjc9NFO2OwOEjYpSRe9fbJF2JQgJUMHyFyonojSxztSUm65J3bBPfBugcueob2lhpkul
5JI3u2QCoG+V4BPUyqcjn7aHa7Lcfx2YNvfxhXU+ICAEAeQ+x6XWTlxab+D0Fs0yFB46ZKWplvIz
U8M/ZU6ARzsgZ/ADWsA0tlmWHYM3Pghcnd6vV5x0slR0pJvWhH3FQMdRhjZPdtog+BaW4hZWMkdI
bVzlXQGKEl8qCZUwYHgduQZOz1Yre1aZugVYYrdfkQij/nBtiXLblxWDUB5/dWzuvN+nN+wBXZ7S
Sc6HfAQ5iSMSaauEz/HY7yIEGy6qRnU+hnvjDu20mVfTdQAgfbFhI3eRmXX5PmlnNbaVRLStj4xH
wu4WK42CaPu38hJY0WNQEhtAtVvu+jCbE4DZaGhNHjrYSSQt1kqXs5dwiKqg5cF8MJCdwdUm4mPh
4jovBpY513p0Sat1B5VkNR1DoIrNu+jF6ZidUFzWBw31axy4A4hZQZaIlaYlVxvwllop6KdeVCZA
gxGd0V6BtYmh8Yfj6MBvfqR6t+sH4wtBuQPKCtO753FXvZfv/NZoYaVji4Bcq7eOQtTTMtBvBmR5
NvkzHAuh54azr25FH7BwpMA5LdWTFX0V7s+ZnOSWsLomvjf7THU3qUqyC5L5bbDGQ2C4etMD6Wf4
Od4zgYg0sz+u9PKMTKq5XiCV1/HTVFzavgGMWBGyKi9t+XbDGQlqP1ls5xMye7LBXAsie5y/VPLz
8G/HvBlCZbZ8w0eQxAPUFSwivl4wZYm9aMeLF9OyzS5ZzYl3STVi4deStq+A083VKnDNZ2TSTui1
/n9rQ6wr/zLeipEFQlpsVSm6CXX8qUTwVaGNNJXfUY/wq6H8p71Bn7GgmQqtguapFds30qDaI7Hp
PNs3WvRiKM/s+9GAS8bcIijcg0B6fY/BBFyZGyRkqt74FC7wGMAGpj+kjev3+3zmN6xLOdfYSMVH
AnXE3t2K5t5sBPht8qoQUgS0RxQiJuZEORPF4YqdoL/+IgTBcote6TlW5DoiorQpxcQlFij1Wuor
6C/6uIUqi2P/VIgAPuFAxwlFW4SzmIQbfClDzqMSG61MPi85nmVTWzNwHuNqWOBC8iuX6B/4lW6l
LMtLGnWskMBzIwr/BlyNVzeBPY9/fAZySBzVJnntuEAZKnsMzJ+oEo2WjssHq5kmZ8Fd9i41YYF5
OtFrsAoPz6F5EDvLQDGhUqbcD2WETSRpl+iXkXl1itTpDzTrH/r16vy8/nQ9S/IZ69jDcpMoNRc4
gWHPz501/Ec/gCWhyIXuWyyaO6/gFSQ1zy3nRA5TUjNDvp07DQ9lAO2xWDVNqnkNRw3qmq4RmYjC
hrt8GOmscvmAidBbGStMuux81X2TWmQEg4tMAMAM4BNVvDrzG79QB/7lI+ax8c1q7ZYdaEG1yJOy
xitwQCovaZ9I7Yovc3YVBrf1NmFmCP6skyh0S2X8BlXVf5umRyVa2fNwfnZerHIwpBlLY1segLOd
lUdHvAytkP2OxXa9MvRXI9Okzs7NqOLsvLqM44ci4ZGr0T6Hn0klQABtf4lUvseXZrCEUt4WXGF3
25E5NXh14cn13UXvBYS6X9bJDakW1C/hCdngEch9F9ezGNttme+8oBbgas47Hi02rSVQMT0x7O79
nv7NBrbstDZcPlwUBSFMfFh7WRfcqHwdV8uwsjM4UdusLcIBDZhNYpaD7ekmy59ojupudEQ3mTGe
nUb0KC+vyKAaejpTIQoeLmocMj3uczJMIGR5AnxbK/spWlEc17UfLYWZCzhn7bXLr2+fDXfKm7cz
o5phH0mesBMeSGuyMdtyLR2tFzvOXZhJdVoVbYRLvK8FjIactJVg34Bs2IIeuEsquO++inrJMcDU
bXAI98lUlbyRpCII4Tmy2LkigrPsXsTIdsLqg1lxqOs6wK+YfhF8YEbpxGsj4pilV1LgHo1WMIZC
eI1PkqkBnOS7q8CPAJaDJ/hAxv7RKv7lRBaq/AYex2q90am7kwcxCd5PNgU8/TFBHGu+icG7/9/J
sNdweTbrdHwBZ5w5VkuUSFbVe2WH2U+1xsYrCq0iIPoXYirlQPOaF/92cfvokw0KWX87K68ey8Hy
syGpG1u8+DFp851quDCAPU9RGrDqTKt9bWb/HrPesbggt6DOA3H0dtppema22WXGEF84SMCWoGqo
WTgs3YDaNY2O/1bPMNCq2/I7Wnt1wex94Cu659v0ZxqYRv12IjrBUc6XDvKNyCiybUDfx/zGlthZ
pU4+bnccVJOjnojLeNUn6VGZc3NUKFhCgUSfZacNm8hEpepnR+tt42nzGRKP3QoBEms4nL1WGATF
uVF6Dha3lWk6mzAdgxT4i2Pv+jGBG51HVhWUzpUkPJk/i18TlDbYpvz02Psxgv5PfA3WLEqGX1Zg
5DCx2vIwZ0zWjRi/xpVC42QcNdOhh5zT5GCNSQ1QaVtDdZEEQYerQGVk+6SFNzjO/2Gd5PadoCbE
etEZLWww95jcWe6riNirGsnB6XEcMUFmA43x9PdAOIpozRCmAvyHzdXy1Gme5A7CRf4QZ3ELWWuA
TWs1JrftSYJroqfk8VvC5mFvGtMq6e6QuZwsAtf4VywOPlrahmK8IVD2ZPkKkKrtih23ZiUsje/f
H/EFWDRYFv8FV9GjDcWTSn+/DdJ2OIYA/KtTZ70PLhLHtpCgdbDPiDuImPuOQwNYG13wPVH8vvzf
+wXmXFCTfDb/F/nK0ERGurKDmf2ClntHxvKcPHvpNVRVQ9ZWo7z/fSQfpzDn4b4GBtwqwl8fMwb9
vbmnas1x/DQaygv/gUU0GW1HlXPNOIUn4ZHJkeJCU6vcHWd70hTT1xqq+AHtBFQk8I2wvSkMDq+0
kVfKKwqz3+lQMbmX7i4fhXTjNn3H3b29cB2ZumzkmvmIHBSEmwu8TU3Oxu+QI8/fTYT9zMMnFZjg
68Q8yjOmaC8OGrXWszdD0oeJKuL9yAVt6Tr5n9oNeLdKzVgRCz/D1m9yM96F9XhjRPgw3ifUm8uY
wvl/erf2+U3GBaSVpW4JqmEUYYnuWapnDtc61MREHbdSn0V0+OChliHFzUhwgmKTuNW8SAZLJZHZ
s1hBa0Z2fYXebS+rSPQ3zYHonQfh+toCbkIIKkAOD1CHJGlEnlbwkGZ3G7bHTYb5bwV0UBJxUrbW
b3pqcnbGVjwJV7Qfz6odrPAzHYbkQggcdaFxzvtGcIpX8nnsUJHlIZsLldvuID3Oraz+SFI6k5k7
ByGnYbGFMumiLdCSUIwsM4ySAba6brRF+HrPfDTFb8PnElCGMBwOIwUKtvpXw6EIdBdelRSTk3jQ
ccxGCBo5/xn9W18ks93WjUUlE45WzjBSNR0ihRbsefPuIyspR6TIuQNIk1ZbzkpViXdSFC5zHu5k
0QzuMGbkHW900JJZfs+zKopvpYA1XDGdFq+CVkfILUuMbMkYTMkytY3eGg2dFnUq7vxy1Jmh50MW
hoQT+Jd3y271CQZdhedzWY8WuUzFYex7rWvwKsHt9b96ZezUo0bQiJnAzUAyiGvI8uvTmY5fqA15
P5oQWidazolqZvy9pHVXyXj4ptRNl7Fe4Mebx2R/NMpBwHQxe+GTzGy4RDGn7ywd3DcePVhiDqfO
MAVpVg1tL2F7j7EKOiIwg6Y90yOkDCKFtV0YaWpK5VYiaRGrXYKJXUZhwpp/hP00JyIrOpGJHTUX
U6n6WZUr5krXbrHCUNIGl80jI4Xs9caniMgoCAkI8ptcMlgS6j6G6kvJDkY8wuh5sXmISS9ec4wD
/Kl24wGOTaJtCjdrDSHbpbCXzcyoeymiRRPXjklz6zTNgV2zzP7xPq/wfzG5zRPL2nxJUMvzJ1C4
OgnxipThc7e86vX5WjP/LiD7Hub1Fo+vDGG+Jsh9DoLGqNLPMs1hxcuVvMA/4GSljjsEVbjBPbw/
Srqug2mLQqMCso25b+LX7Q+2k+hWqNHgTVusZ3xf1SqlGYfML8MdHxoOlzBjoi4fEV2IfW0nCUUI
I9Z40O8HRAV6c8DNXI1m9Q7NIc23lGLITlcaI9oN5TtmpdnNLv1sFSWiuyoXgMwwMenrB9D/aJBa
zepBEiWltVrMVXL5ZIotLXJoWryxG41vT9J6r99r5Of+ZIHPZYMJqOMb/TY5b6qUvXQRyRQfcJBQ
8SiK1LZTI0glzXg3f9gBmmcl2V0ylWFCwPs88I7Rppeg4WtoqgmT8jCk6UXDcEhOte6kSin61h29
fHL3nKBmVF3pCMUnMbaH7lVi9+ZEthwWWzhRiQnhE+d0zXAclG3LfFRNgPbO4pPUKUAk1t9mkAAs
ysRaHlWiru9Xi9p6Pgqg8kziopGwYrA0MRtGJQMXkMi9EFu8Dcrh9a0532WXR9QveHApMwL762Yg
zaeJjNcs9jDjAQ9OhaWG9uiCXUzCRkBgf0fnFFzkmewGR3F367hiu18AQOmrbfq5EM8zsLlDzSkI
z/uI1CCe3wrH2UnNT3xPKsHghQzQWf5vIpTN35fel3Mm/9rGJWJs1enpUsTBqtE9joFDg8uMo4Gi
RvOPnJEJmO/YkhHxCEVhDXZiPuPgGaaiJx5PROVYGi5pDy/HEzC6neUKdHRbNpUwysyBTuQXip2/
L8V61kCLcS7J/NYOJgUue4dxQqgmkBMFdvog8ogfHCAm5XXIm+D9Cw10vGefX9SypVWbByqbw25e
d+BxJeLU58mXHg9t29WZOmxugrAzW4wLH0FaOQXyGy+ZaasAqe3RGesJUKjtCsveoQxoZkJshka0
SUZ8ljy9G32gDsLzXMwYqCXsByinEE3zfQc2hXEkwzxmink11frZvwnv8vDEBFeGjpbxUzMT53Cu
c2OtC2kI5TRW4Wh50osekDOZ6YUFFE2HkO3tGdyBAwzpz2nn06HyxQ7+27RZRmSvxTZu/PwMJa8Y
+pjW054uKIekbjJyc2NWdsFpGo+rPCQBkKlJ+rT0eva0x7op5zrKHwkD/KCV4EaOpi6PUJEhgnjc
VSKCKfLdH8XGF553zAI27hKTw+BvKlZwFcljuNCi/DcL6eL1fwv6qr4Ib9OQLSV9Uk3Gt1Edb7FW
8EzhzPG0dPLf0TUzuu8cygWOB3wiea7934/6SzaxHY0ijEU1zNcJfGXZ6Sg12el5mgVIZX0df2XA
IK5OX65PU7LUhgx7ybyTi7m5bzFNa1QUCVPU9FEHkaY/6uj5WvGAWRljJD8WcQy1cZTcacAeLJXh
qAAZIkwPS0YmVDgzcNnIldRtm2wgwmuuTD/oZXoRzSRjPNloQfGz5heLbcMBiQK+EZ001/izRni5
N3cbk7SS++9Dw8e3wS+/Gh9vRcDkNxo5FOOCzK8zDC/svN6MvJoyvIOGPWvreszVySRsW9+j785Z
ojOIunVApqUasVAxbwykqRf0B5eyggxxriDHi2+/HVwfXWA5upNpMYv2mT6Cpt0Epzr4y7A7Na1+
Ex1scngc953P8dNFlEEF6H8yuc0C52t6bwxxkYRza8HVyXnCQ70frD9etr2xhnWNn+X9G/fYZ6XG
QTsXhgEDZ0fezfYsIsjihrM/OwBd6Hbq/VwfopzQoushUVA+Zo+OzFwcm3uywWgW9ss9Y1tVRzje
V8+u//69Fdb1s4uqXw+c95l0XO2GpyQDV655kXXM8DlIIdJj0VKZs4+r+lLDB4hOULb96tRbNPjp
1Qtg/UjhwqhW9hOeQ/ePKhj0l325KO26vCIgo/2skgvPTQ9FvjXsrksnR1gsJeewHWji9vIkqXN+
F4aIJl0dr3dRpQQWV71AefBl6b49Vx23Nw68Q4igJvt+XTV5Wnzcand0aT0/Mx2BPi4iRNF7t5cr
gS3XQ+kk9tZxMJjyaogfJ8qSAC2tEm3ObKpYkFgW/6vIEVC3QWRxfg0SzoiuNKZqAQVhF8qgn6LI
MCv+HucPmQ6Mfyy5QGM5Ncua+3QAcgCi+furxyKF9fsmdRiNlXJb+gAOgGXO8LVY194FENYON4d5
PgJ/qTYs8/I+PprV6H8Pjp9nn0gxxJ4dfEyHPy+Ekkmw86LJuIn5Bb8150aQVp06ZWxjImjnp1n/
rEL2UYbHT/MzoO2bwwRs+TSWTtVyGFb7hqsKWIsFbH0xXnXGMp0MqVFK9YWMhb9N/6tab7fgnZaN
R8t6T49U3C/VmPKGUpdyBPKNGkAhStU34tDzqHcAOcd+63Y1oV2Wgu79u6HlLaZH2RcJQNtMG65H
2LwFgpY2oXJcUn3qNurfbJBI6f21I4s13t42wMe97pmLRxekl6SHSPTKelMo7wwpiGK39jC9CNxw
cWWBNTBGx9yrWMDMEJlib1K/07kc9n8b0jTCMpg6nnsNUmwKjSAb4fnoxpVyISeLR+cChC26mCNT
t+P0R4P3K8rLsEJI9fM5hTTTkBIVxB3W5KFzmvI4rZtDmtNPZypZSHCX7v0ZsOFJZZNlmANojx+3
WCusb65GaBLDTpvhDJ8TxDsLCGG5juNdROwqhEVrZGz7VQE+Y0w7lM8EdOiEGqUnUBnvscmCAWBt
Nq5ZJLViWd/fieqByZoe8IjlysHimO7xiUtl+u5+mvavq7CoK/RPtNYSUDCdbv5AQlkkRwG0klpM
8Ui3SQHkYCcbrd9biIJkvFilTrZ5CjfzOCKeOCrMRKMTK/rSSuejt1Vwcw8OWB/j6xGDqYdRvfqV
E19MwiulbJUEScsGcDC0H8GNhQOmFeudl7/uQNRBVDKHwvqz/VvQEfhcKBna5wsSEZHBSNqqgffj
TtRY78bQtiu73suUQtL6d2UXHlLJhiuOHw7VwOkAEK+vhQcsWdXx2zXLO9GDINUSpA9lOndOMppO
KSxzWqSWmQGtwPi09daUnjWEalpNCHpp+Hl4VIGHVNY5TuBCus76u1iLFXgPVKGFF8Zz8ogJ7rko
Qr2kImlUPVh+t0N/Sq0n1ppCvpHxXdRW2r3QljNW6ou7VIOLilAX7W/KlwPD95Fi+GpmaFmvkdDy
AlIPEq6qeSI7bGCNGisz6eTyoHAjBJH3dQGU/0tc5kiajeFHEDV73ZycdXRgZ//nQ+OdgFJuL9wj
QV22o3NyOWl9Zvm0/7s9IvtrxRTCBi1+bZHfv7MQAboTaLaxl21t7Pjh9pyCnq7HY4RDwPWOWaUJ
riAug8pBPT92No3aJsMKzDhiS2zT231zkYrt/XrvZcUKaoxjbt0j2NAtYi7VtTccjIA9kVovEsoG
KIibeDRjX4wuU9+TWRimd/vwztEV4q/zkbb0FOATdvcHkFyRt90wbNw5Au0SOeGglu6KLpSJaGXz
g08wPAypoIFdgzdxlCeM8/Tm4Rp2J3oPYrJc1wCzGkOtfCyo6XmkwuBBn0hCXbNcnCsXFaPQFRHd
ZORGyviePuyVcyTzOnl2+qF2QBT3zLXg0bCSxwphRIB/NUtilzPGjs1fAlRcqRvSLBzARUHPfuzh
7uDNOnQoWNDDJFIZtg3S3Rkh291bhXtzPA7WvzrvFnn/PeCvPeVxwubBzw7V7DoaHV6DI4wzCaM3
kRPT8H36Spj5xByZAIQ4R1HB9wmEq65uWZ1HOLDj+dGsw/Y1ngmCmwnHje9P1SOSEYMyzuXhiGIp
WBEVYkaMbyM6S2pT1FQia2Ga2cG7Utb3ATEePJ1GW8tF19dlMCRGW/vBgAfrJpoTe98SBweP32Bj
qDkdzApwWtQ96feN7dTvvw9O4VHyRPuoZSiL5n+Qz+Ympc4CSltLgRgVdLmiurHLZ7v3K73DkTGR
POL8vcvYiB+mj++Dz/W27kxhiiN283XeGG6SKKfYlDDzHsYR39MkBPRDIotikL44E2A2s1Rio/hE
pF7+88eOxA5Gon5W1GzD76FvLHbY3BhpXpmpFFdDYAO2N20oKKoKWO1WxG8+5z/tropaeUwzjNke
n78A6aX1O3oOJojhV4x92zWWOtbQg8EPvE/sTfKQrFVINg9ipe/HSdbjgz/KB5oCAf0Lg1DClVSz
CEhMNzjvaBaBISEtrOsDT8iEIwU7spnjnxLltGRSWuFHr1KZRrfHuBN9K0hiF72gWVA9Gm1hZiFp
toEq8qnEMTJmuXojkPCtRvJBA9kmp0Pextw2tuE5UpsWOZLEWzQcRFAlunciMoo97wKZF5oYsEvH
GEvtFo9ZPO1Y0BZlL7JRLEvOmvv7TuLLOSUdeEO1ZHr2EkcKp1mYQ8nHnTYD4ArtQt1VyDIDA+7X
AKXHsT0hXC5EZHhBYWtQD2LqVasKgfFBLoiyAiNwD0jU+1CalhN831ojvGq6Cyu2JU0Fy+OWMHR8
2x9Le97Oziql3b3v0/oXMoUZ7viWS0S1nSv4VaBeLaubIg8QwRCMT0C3aqYiQ/aXs/0WQ1nsBkZJ
hsQY9Ft8tyT2ViP0gXYLYP3EokkoUbD7vz2PdYRTzy3ZYqz1viv/tCp/LB3Tigh719jAE+WnCz57
vqwS/xSrMHa/5JVejtRN9icZy+6sToJQw6WopwP4n6W838tiORuvJ6oRbNoLPe5NwVhwUR/beFyf
USRb3WaL1nmUZ8kJumsCuvXc99WMBqDZODku3EYCoz5r+vHg3tYx2zYc4BELXaa8boVq/hah4gyb
C5cQjjkaNHAAu3GCo8pKVj0nQGfB3Ndp2Dn49uPGKDCvqMFRXeDd2d9uvO7NhpGJxto1OeJREBNf
wlIRBjw3Yuv1Uz6yGykdzwRnAT99sPmYQgkX9D7JXkOzcjy0+1JummGoRMA48mOjJOXO1HbyP9+E
9/ivjbgYt0A9l5q6rNlSQWpU9xfB4Is6FZXpB8fwO7oRq4zZUxw1AJ8BkDS2hrMEVYplYa9l/CXq
XoP/u7qTSXQYILjf5CBkNTkG/cAxL0cYHG8yFMxLCPBw2IPqYfLBIL6GTignNK6G/WSNznVs3x/D
Q6AOdkybgCj6aPm7rfO2MgDzqzZSsnZBnacsOWKGG5yrAbxhQRFnhS9RejjVCV5wqWLft0GXSDhz
vzyYYrzPTKntYIYhw2cuWdhgZ8G7jFpCCe9z93plf7GjB2y21lfUOcU19QFW7fcMGWcBiA1H77R4
HsNhymwhkOwoR84Ujez3o9k8k8hzugSTvGjnVkCW5n4SwB4R7cf6s/LQWnusItFEaFDct7wZ5k3G
EZLgAbPWy3PRlALYPPedNh2GIiOP/IWvMgwjiJz9gdajL4zVtgBBUFdK/ME8l58xW4Y27h4QXaeP
KXCtXTC8Pd3WCmx/+SyoB7PdTw8z7RDIZv/Fq5+iGHsnq7sU1+eVwehfaxzTRl4pMoIG544HUorX
Cepd5siahHQz+L4b1rQjRvkB9NDHTxtCYZb/qNu/m+Y0CE8oUcmyIQvZ3KnIhhB+RiMu4b7W/A1u
T8Tcdpgrt1jU5hVGzrgo8EWM789iBwfLH0BpYAz3dA7HjPiyxv7vJEBHri18gD2esg/tfz4Dnu4l
IgjemrXqWrBefCye7JZ0b52BsGPdZP50Q8q2JBd3pZQ57F/KfS1xe4kBt1anDAJvEa79xdPEaSyj
r9gLEm7oQNGEqokmzeHRXNodyKpjt+2h4/LJFqZgXkFySNrf5/aO80Zl+LHy+9jU5RgX4C1D2bk0
pau0CBAoiZoPQS0zMD+FKXrcJfGKvWjw+I7PI+YY0Vn8rseOON8934h55ePl2YQjhL5B+yWqbGQI
DYWQ/Xu6dQAiPOi+ZYUkUXxqp3IQfTHayoflYZLDa7m3x+HQ7pl39cqsFzZArNnuBVNscC9054W4
TiSHLvTlt1En/cDt8s2aGazC8vhlOee45YQU5ct987KNc/JwL249ZgAMeuk49T3fnJGFXSDXflx2
21kdzNgf2MvfT/HNgXjY0arqyWce0AIh5zRYqjLcW+86CBRPGVIx3V6Y5qJhurmDVhD0ezY2BKG0
8e0q3LFBnd/hIdb8UH2LwRD+fOIpdP2OYfujJOSIBOSNg5SlJEEE0roNebIHpNxpHV26bV9Ld5sF
oHiwCD0aFBKrK8VgswHVVb7lIngBrKsDkxrn3cMkY6qZJiJo9NhBzOHa2ssV4Ht9pBSOY41+sGjY
Z+o8fcOfvPMnWRsbiFSub92JVuC1yE4CtKtQNcdCBwPF2JFHBveLjhAsk1sInkFFumwRq1eF1qiG
AT4gEmhZhggdu3IKP9Pt6diIF3Hi139b6CKX3kiSa2BbG4t7PKidyQlVwRe4Kkepu9c8v6h/Ee+l
S2PJt+/5b5xoHMdfAgrYCEJ8KMgQOvj8yX3Ygilw1LzHXk1wf9e+t/HR0Zheq2+xvaWejXvCY0CR
h74pQh1GI9pVXcfRydb//LXTOgY+2DCnfuCQ5Kp6ua+WvqKf7xFs5meuXpWojC0sHW3eBrsnfmCh
sFb/c3O+U3vdOUJtzxA5Q/SnoEFavUCcIPEGXgGPTQInnDben4gQmu98Fhw+8fjBEL7y/ktxjpAu
s0KqpxsYj60ilrEL/F0qWrhShsbk6hMeZZSJyvAUdmZGMPn0q7W6oFee8fuQR3f1OodKct5MYcav
TvXRSwhunHY6sn5iNsix2Fldc/TN7fQEGjR+nLdSHQR7DhywRyHiliy7KytiTzucKZVscJHjcNTU
CNBiPocXiFrukqHOUwi6VTw7gYQJC/7SlDI/Sveg3rD/J5HglDmSCMjEe9ApHReTpm0GDzC2h+y1
U9XZb+VE6V0MK5sCSOtSBPp+Nc30u4y5ilADdJ8dHNyyPkMB9lX2J8iKWghVNKXhFdu/kH8aXiaA
PNc+o3wLZqvGzlatHi2ejRM91ENoCm5ob9xfTysEJxCC6bJILtWTHmrHoKHNFpC6T+ZB5XRZbfuj
Ubze17s7OG/rqNXjrEGOmBH35AitSqPePdI7+8oossY43ygysKfKPIAPR0lDpQEUfGSErN6NzlWE
dePAe/Vlh005b1Zixm/GBqwxVCT9wJaFR0j1Y+brRW0CEIxBEVM/moYievLXvSb5YzQKgRGdfi2H
V1m1lc4ATLV3RYdv/X0J656HdMxBWsaF5fq7s7Q70+FdPagF8Bz/8mc7hb1L0Q/J8a7qR5Cet9B2
1Yrea7/7giMZwddcxOLVQug86GAOrHkGKQAQfFWZr5Rh84SlYSIrMyAfAEUAjc3KihwskgaEWf9t
S11e+fCuMw66t/DqABVpJ6af3RXKQAF4CZx9N6kOC+AyIV8qaiW+hjNc8zbp2nvxJpdpzm+B50OX
dvS0NOyT344tQGBm7dPQoXrbIQl2nZbhs4/LDDePnBbqKARSBpo802llslg94mzYH6SfWlNbaTY/
OyYxE8cB6XDCY1eQtmGy3WqSf6QMtuJIKEmS0GFNzbcgDGGwtm60MDMFWdS+1LxD3+H/ZRx5vBhu
j5ixKEbnERAPOz/RoJcg3jrdOOOZhIWRGHkwbyS/I6g1dIEViNrBmslIyTEcb0hwCbEtGO2Ld0ge
Zf35nXEOv1E/xlxw729b40TlWDH++NGFko3jYB/oGhNZqtLOmxjwJQiiDBVVV/wv0wbMd5TncXLO
oF/cCnKoRoQ//osNA6/cAAqJ5nL5VS1weMoOTveDylqlQ1e+ViRKy4aMkRKaoXv8Xo0e6I3bBXnm
MWGUJL82QLuB3aL1lYLcbvp47hO+tIgeeCHcpQXadXpLYGQfrkjzx+u7e/dcF8BbWPv54ZCK99fG
d1D8UXLbUtoEBWb3N1mqNbRwcox8+MgsJ+w4PdTkrQ+xn5xIFvrQp6bRPqkA3R54VkWcsao7OqA6
tA+FNf4L3uK82FO3Y2yDyhTgF1Wcqnc/rKyEOQ+sRq4cR9rMAVhSLp+9Ag5jNh91JHLHDmyMEW2/
e+noWveuqwSQlcsYLic6GXg+WfpmetoEDANi0amefuCJcC4GqeCw0TmH/TQ0IOhfWPCfoBYRK/aJ
dCgFY9rH+QOwJHLmEr+Vb5zTRhIAEq0JY3+F4qE/zF0+IVStTbY0LX0eZfq0qIVmP4RMesNyydRS
cbvb/cVkDcXhckfidYBaaE0iLChyuz7FDQDKBJrUQ+aDXi1OQ9AO2wRMURRzsa1IARMnkkUdS6Ac
PBGTjjYp1HZwsDJMVrFNkyluKEowa5sMHmK9z1wrM5RiEYM7sw9TDaoIkO3I/rf/zRxYwe1KvjOr
n+gD10rmXzuFFYS3lslOz/mGgjSXa7hu3MHXuHT1ZUgvVji5VqGyi/jWHQs2k+pxOh5m0m1PlEEu
TPUZPb2KkVfDP2DVUmro5LKFEgJA6gFEgSGyM+QCC287QRJ8gxoB+Sp3udyMFtcF3J5fXK8B4tGs
sPpR87RhoBDvNZkVHULFw+oSPSQiiC4N5D56qLXu89FZL05dHtyxfNKGbkfMyYkb8C+MaZm7Erkt
2gZ07F//G1nO0fjsP2O/Mbv7ujwETQV0QhV5gxyocctN+VDIRE7n/21a2zXV80rUuPqg/zZ8VjzX
DOhHJUwv30gpMDpsNvHzzlwOLxIai9AY0r2FURsovN8L21vElFaPtSrgLGlJ9FuxX0MnZQSIvDWR
gkSDm+fuPnbVnm6PF9T38767gt8e5ZUzXBSebWkK5YBD1yWg25YUJT5borVA+rA4nGPUGiuj4//d
dk3hXrst2TqxPJrfjvxTrXTUV3lMGhK22AtxA1fOyZt7nOAj9iNv/j8JzwTvYisxrzicQeCN1qsj
07W+9WhWQSPozD30dk5+pLxze+24mTeyNT+hlKbpcAPEkyeGgjXhwnS24kXjpt/qTakztBncHO6O
MB1nuFicBeWaNB2UEGVGsR0aZQ7wVU2CZ9TElBTd8Dl6/5LPkB6dPrgGZoSF1j0UHQpXXIvef8ZV
ixZVGP41RdTC9D559XUfqtjTF0EbU4u8oSR7VzYfdZa+SPZWpW16q6fEd3rB3pyEJqvCbT22P5Mf
ZkJ4LiHGJ4eAFJryy9DiJxTRjytJoowIx1oZKTI0w+11OjTAYZ5oq8GolQC0T/mTXFQzQ5yDgQ60
OwestQvXQAzxUpNdR4+eaHgDWxmnG6c8td+WkwPlOfQ1S/DB4OT26oJxXVNw5OeZSnzbSrndb6yZ
vsFyCz1SPfLDQASlSTzSI0VXdKXVlb5qKzSQbMwE90oyHyB3ZP0lZYPYcJ0A/o5Pd9xdDgBpsSlG
uskkldnVqe4IZ2YgVxa1ENcVPA25gYr9dm/77VkdIG3ZBolnv9eCaEUjyhVKbQZ1hBd0bXzTDhYn
o3EpHDdLwC8RdTaLQW5P9peVycM6p3sEtPTNzvu2P8Z8QFQp7RjKK6ajlX5hl8z5j/QEu9verAFm
tfWVMwDQyrxtukXH9Icc3L6FH86GlFl0TjGzKm6+hLgitrwow6YHpuglcFjCegJ9WjpQpYzchep0
l4drRLixpClYmecvc4kkTi3PRGjLyyxCdVYnsh71e3abk1S3y3V1p9Nh0iulf163a5B58bvYIT5t
JpGi4P2U3l1RzN1xbAwszVMcUKVr7J9DrFBk1FNsfEsKzeXKgjopAP/zaE5LIKxYUkdas7t3+D3a
/hwKez2AzAPBi8Kx8hmiJzKWlf2v5x+Pr/95gJswg8oVcF9XDbLMAJoBjp9ttLEZvQhgxec9OSx0
FwS2hxcPgfzi6bwEjU9X4N9/Vcf8DwiE3EJ6AxnTtrD8sJqNsxYDJbt7nAnWRmNNyW9EPgGSMj42
ZeP3F1AhVynzO8t8MBAUfHyPpbImYkE1XIAJBOfvTQkooWTvDOeTZA/gI51XacV5buGfht6L1028
XLkDAZ3zOihfEAVnF9wTfzWmALYag8B6fFUn8GXLPZm7+M85E5PRwFXHuHIBCoZ9gIFy6nqS4x8k
nYpuHEnKhswF0GD8uGYxkdsnkaf9EE1NCmSToiVndZ5L5HmofKji6319ZDooNAegsv3gYGVsWqJA
VbfK+s/XGtA6ni0eAF11NnXrBIypudA1cz9XOD0QyaA8Lz0+XeQerk82xSeZ9FELjDeKyz6OwTLG
EOu/RK35ol1RxyZrZLKqFSEuF1qJW0UebJWOrEj3Ld2J0Uxx4mhBWkYsAPi1SfxFdtbicerTFhIJ
qvIFYWw2/UGlR2F/ba8Gurwg2dpQ+ZT0D5XeZV54GN8EvT42dWmeWJFJiB7Cl62ry8A5LPDO9FVZ
OnaE2TdPi4LhdYPzWggrocpi6Me2zgTNgvEQqlLS1/e5FPq5Bom0r8OjK5A8zWv57C6wE638gAdX
hMTACoIzmBBrYAVrH/6t9Agj4kBZfd+0hJ8z70NWeu5n89DGiYbuK13s2GcfVA36vzTZrIXTN3xs
PYulmVZBVQfx057uYTq+Pz8VInYCTJkx7eqfHBEanrmIoR7WNtmgnKcLdIlyC598T/PchVgZiCnI
f5GY9AaJ7nYNzaUbmHCHaVlF66f18x38WrYtlwTTMNpYOwnkynh9NC2Oy8WjZ1DAJq3Sn1EkLSn7
cwKU5Rek6w5aORHZtDlEGvha5k9DJUNMWHy7lk3yG5ZGJGaGBAw3z1vVipC8NcssIoG5C5TBrALw
BSkJbNiM9aggHxTwl3qWlpQ8iE7d21wpibDBwfhfBitCKzrOQDDiGEyH3ELM4D7L5vTslTZBQB4a
1i2vSAzgEYVsTMuF+tFJk2H/ln/w2Bkw1yZtpEmqVJPDbC6LpvE7qGXAa64FgAnr6zA4bnJRRzeV
StPg97ZD5vfs8F22uOgVNI0vTnWzr89r/Y5FzVAXax+c4DxXCCL1WDXtG7enV/kbyQlUtYTLMRmZ
kCszl3SQPthkF52D4EdprwkvO7ntJZGww3TYJmx6ZKAilIz6cerUfnHcbkxI2Xs9ipap+zZ3F3jW
2s+KXYPQ05E3CMBV2cA1d/rx3fPT6MvvWqzRNUIU5N6I9fH1mAwyP0D19/QZqBLpwNm66zbAL1+r
KidBlT4gyoLG9oFqK32LlK6kpclna0ysm0kN8rHZQp6MlkeXTyPEbJOUwfSLhL2voZd5H9V4FahR
ckZWVjH64CTAansw/onyIHpHIXTEchaawQytfYRO0nb02dVw1cLB9Q0kgq12T1Rqs/nDTGkGfd+b
JPbUozR7bwwMbhSSxVao13WgKiMzzKnMKQg096Ydi4k3+RMthY8EZNsijKdgwWsrV4dej7FRbOCT
lh3Yx454ghlmmb5ySpg9bu6IXHVAlsa6i1t+zvq/fyDWLQh93xyqKNKxQk/rqNPC173frqUpIbBD
0ZfWljGUs2eoxaMTToWG+HZdKd87+UjwkiBfWaAgElpFTor56FjwNDl5nZ+n17n7erZIYv455tJ5
JxKptU6EzwJ7qcoCWewRkMzsfPCMXVCx8onDKwYD0SPNspXtnoa25ljEQLpXVyBw+XzM+j0mMNix
HC8Cu0z5ZBCL8lMCsbrWVgWEJAcGOxyFauwmr16Fft6XYXeB0fTKpoOZPgQsFx3an7t+vUUpgZgJ
C5IGNMfe99g7D1MIm/FJbOJL+m5/2Oknkk/BWQbMQ/fF9ium0fF5kOujNRSDJ6nnmIPMqAiEMgW2
QTlii8wuKDoPfGzjhs5iH5u3IMAlpRkh0VdYoSF8BiZo9BEU5Y8dGTqDM+nTrTx0g4xHa77ZGomr
ZeM+Xr3KzH507J0akxclmKjXrvMFEtmEvy9T5PrQGXxte7gS7ZT9kHvoCjXuJyBt2PN9yRlW72nr
iRNNmYQemo3L3gPxxl8mF0vEgGni3KdsLL4hwF6254aGC6HrM51tvFpWXro0XECTpZuyaf/LEgpt
NjUKyMXXXBLdS3Zoh68Rx/Cnwoiv+Jw60Mw/FJqxllrPVLsVtPqWgeCWsy75sqrN2/fjoLa4TkaP
DKsNNWimYcY4p+3BGhLvGoUibv9UN51umtt1V+jl+dYHVPcXjfgZwhTsJkGiMhP4Q818nCSUcRhH
kKotGyG+RmGX3C3r2r6SMilE9Px3yiSxpMK729zMfdKA04RYnaciiZhj68PWSKgUud7c10JqmKY0
siURHeCXcbHByZzxzqVDt9IyfHlpJmoULgoxAHLFOGpToEvuSl6n0KBfVdv1pvHanmF1CgqJyUVU
/XZjREttRpTvKZUIcbePsFTdJT5YRXmIRkYXfYkYonWhtgqomCupSIyJx1LNcE3PMd74oRuy+Y6S
WYhs//Vw8Z6svdH6/iGeZU76bBlVTEUhnmYpdX+jPkpupU40efsvXSmOG0ftEvoAeNSaAa9epPKH
XbXKtZWuTqG1Wc0wjI1lbdyH16EFm/AhWO2FIitSpzchHGbSDZMIlpYpaY1ylXA8MT9qtdbm3m17
FAx6dNNQw+LAB5Af/xz/Gg17hXb/GlUWBELi3AdSifWXl7sF4v8vdIex11Ean+8tzbrvRWXTmgGH
VgiiElZWOH7OiyifGi0OONSae2hWUHpOwqdXINs5A0uGqln+XY1n85Vh3HFx8nm0nH3En3fyF2qz
shRyYgf9uiwDbBVrIFzuP2qoW/4va7dfkSTbyqF6/tk0rkD1H1ICXBgDW9VjdiWRxnDxfKRGZWMD
I0P79F4DnR7rWsfb50+VuXWjAHvlCRHRSZepCoLy7VmqMC3hEKYwizeUhHknNMsVHlScJ2vSs0Mf
rlIOlUqatzXZP236LpOg/2lWgzatrUQZFb9BecoemuZ09tJ6ELs9M/qKu6TPc5wNwR4rvEk8thNz
DNrQr4tThLFFdDlZrG7jYYjPxmg//uqgYcTMIYfaNas46D4nVZFB5nX8w4uI6acTRYoKK0dmuCKj
AZBTBbmUd7/yc+RINYNzRrRMuVJtRMJxfgKC+PFjt1QTfkYQfVlaWRVJMcs71cHKXyDj3mjMPedx
WEzCghYnFRkzUYQ5cSexo+1uqVtGXSwXdvn/dEcXxwpnofxGqFqtxI8pCjq7gY5SG69cL7ONieN+
pHLrKzAlo1d+jHNcRUL1VTxsCtrs3dmlUTQy73/twWl/k3EktJ3Jh2BCQT4mx8bobMEw6vjlj/ia
IbxS4ygrBxj8XfriAi4lgruhrfC6JT9rZKbDc2hMADjpQ53WbdBs/yJQrEhqzA1q+4I7y8yrm3Re
/YxFBzjta6cfD2WRdHwYLX7+6+X/G4aF7sCjXs7/NFub+saHRyfsom4H/u8AER9tK0is/GwQsqT5
rg06wvwe+/GF2w3KPMjbllMk1WBUex9t4Us1J5aanfidd+IL96oB5ft/3s4QOtvhTehhoGQ/SgvN
g8ADYgMq7+px9DaaVPI/4kslHBdvYAVdLe7BEt2dvgb2+W7R7HfdaacBdTHVCHUPWBM30dZBc4lL
OFOQy8HQ8vXqPhlkZuKmawMI6zX2EsuFxXV+cvIlwsDCXJ36wPkhkk3f15rsjbtbIKlHLfv321va
WBZ/UzEgCSdWb3dRxPTLSLzMPAKYn0a6Hex5/Kk42ziHR4RUzVbYhvTkOtECxJoFTSRuIYHK7MUn
7dZ8jocX2mZFrxQbRbzmaSgjwUHvqAwybnijuV4yueyd1wf7zT7+J5dequ1DE08VgkoWYqvB00nZ
4pYzZExu92Aakz37KpoKgbzqpL+CnpqvhS7eCjhwaqaHD795Fjs51VfHP2S5hdo2lLGlyM3PRos2
gjyq0hFKr1NRitbrWMF6ajZkIdyYFFYBZwR1PU5FBfmRpVt1YG7cDLpd+mzZbGTUBZY8qRlpwbor
Orpow3F8uxeaRLku4vrkw279c7PkH/I45ZnUe/kNRaWZ1nV8/k78iEw17uGWG68RecWm9T4PUatN
plemhAQ6vCsy1yyutlcINNQ1hc5YuxoGt2jUe5mCd3n4rUZMaDgL7y3T+H8ll4K8AHAoadIqwndM
xMLqKDuyHfV6UjwsrPyeSFfPWJzLeOoEC16MnSjNVHmqWBzMv2ZIJP6qXE9sd3HUyhjtScem3VF9
/129DeT7vKYXdTUbGee1jszxXVT5CafqBof0GEwNNm0FsGW5V6NQRotnEJaqVGnwAm/PwmJS+O9H
RTOF7QJQ4d1NneSxWcohhpOkl4yFOqHU5I/Ap2EK4xKkqRvTqG+egJN2p5yxhnV8HR3f06DF/kw6
43qjrp49b832crOYffMJw/t3XK2TCX6cIlVbX0TpFSjbEO0x+ZqK5y7ZYk6TH5DqVXfDslSHFWg4
KQnB42CYDYKr3f7B6jfX0YQr65ugDJe4JHE3wtjz1LYKD7QkHB0c0lA+/nyEZiaqEof/6KwHg1Ai
2zDqk3qpsieDUPtCl8/eLW8ovEGomCFQhuCFVU2zZBvlCcA6A8X9QHkef57NV/eB0wUB0XzoBEeW
dbyVpOdwH7b3/HUwdJKzItS/SgYXi5rAeLWvrhs1mMB9prR0gbNFEM7/Q0M/X1Nw67yewDqjVYTK
Yxl6WkUuXQqzduB4qvLkJWdbsKJMqCa9FLuaOPAlKJMIb8E5gNvvc55rYMsrMbynUtZpqE83rXy9
+nhk7cwk7gm4Heq95DGQPzGph/q8qlEg53AiYKMdEd42jRKjARwuyEBih9VaBdtZWzr3aHAORvbQ
FHEdZPv/IlrpBsBnDz9HSX/06UemBlabP/qdxSkwskttvscziZSjOqvYtVRu8tq5LOS5f9GJLZ0y
xESR4q67Q6b3GiryhXo3xX/RbQTan6nLwqPLt76F1lq1dRnCdke1jumP+wV3zimXRHLOr9gUcGx/
Fbckvj8xYLMHNI3Q1XqsQdGyQUuHEo4iUSA/zlkkUTAYPl1P6BWMtHK1If/9XQRJDZTLGHi5Rd7J
W+OSKIJtKZEY+LUuKDF10jfi1vpSAdjMKl0kbxoRITl/KlOHwURs8I1WIpEd/dWScCQVgxIh+woa
Xom4qq+Zu/2fsBZFa4YiAlXIMeCthvos+XSshhNZTSQOGoNVM/w3eKhCNvKSRH5B06Zk00/2NltA
jTn2mswc0gVmDD4CAJNxA4dVpc90eUHBFgUiMqgXH01QXxBZFWnWjpca4auW+E9IlmRMoQf8cxvj
oX83e348nJAcXkxQbEI/6AMb0UZhfP2T5QMBlqPUtq2xPMa3KCamScwYcSTb0lGKUqa8hCauhSoj
3QV34rilaBt7dRVU1HLBxsIJFXeflZNiNDTKF50DMsNqGfuhitr2CgNZ/GfOHwi/PZcnckhDUJi8
RASeZYFHYzsjhbpUd09lrl7DxtJjIZEE07CCnjM+IQfaHmjXXt364MMCZ9d1xAezOIUwEb0cjMmG
1HBMcAeXihnRVpeX3FRrpGIRCknZRqajkwIQDiD3xHhZ22kpZt74zD1d9meCNWpxfmfCxedk6nIN
bSv+dMFW52vG+sBb3ks8IO4eZ5XNUCSEnEF0H3RJF8E16ohlr/+UoGV5nm0EPqDlDnDcFoLe1qsr
r/Jc/tzJrqdW9sn0mLYDwha48lJox9dYETVrt3GHmSxbmkNgGF7/tfEHa/Na6qi1aHmC10uU16wz
3JBNcXQ1qz3/OiSc4n4cqs3CrtULzYwGVcAEqFwXkzKGoppgUpZHucVSxULQdLAL6DGnpNmT6+8V
2MsqFW9NFi/Zn0YDVh3x8Y1x8APKXHNF3w+U/uSiSIqA8MgmM4z20qHIpB/w7DcOdwYiMbNwpaPG
5MCv4a3AcKWWG4u17igHbhdT3UEWQ1V53WEvCYlEyGlSrM2SMyM7jr7lABvmCwONEFnKz78i/9VN
IMWrrk0Xebs/RiEzt4XDMW/9EStiYbBevEPowlJiS3L/OGVkHXWmzwv967shEkwQ4gV7e48miw61
sp63k0wosUKacYfVRJMwi3fKGdqpeHtQsMTwuzEiFzpwIliaajyAoyHkiAsIDtEwqBQWaXa/UVkc
eka6agb9MZfKv7tXa85clLFdix4BEffgwQpWPsfmLiDEI9RhnvZtoHBpaJf0gTbfTJOTjrQ89vc3
sHrZiNib7CADGYcgZb2WBwZyC+UMtfy2DggaZVj4FPd1Sq7dtcbqGusf4Hrpn8STFl3Fs/hDznHD
CEP4S/okjcLncVc6d8YHDKv3nxCr4D1bsUXdPtP1bjZHIP/KgYRfy6UvsqW1z0ozZDX9SvqhMZ2p
qZpWrVDboy2MBvoRmrVP44gPCb8zcAA3KhlqLoCsAArjB9nZKty8JylKkxZuuZzLzjsYYYvrAMCg
/KOSztVMtrzNa6HHnSRXVkckh+C67NXbsEYcRvJ/p4m8q7junbdVMuYzA7vWU6ktGMKFZsytjFXo
lXakfmPWDii4mqh5KFF5f5n/rEiOdYH+7kdcRx//+581pmB7Ku7C6vmzDEkrHsboBgI66Sw4rz32
i2cOKFPVQ/DEi1fMZ+dqmWze/vs64Th5eVSzb6NRCz3opvU5Yljw5XH3+ASYtZXEb/yyHImH6eex
Yp5MCdy84US5wDr6pI9oF0dQKOF9PTG987tOVEI3c4CFFEFsB6z2QEAFduAbp+LiwaiqMgFoyD+z
rwqaifqWmxJ+WukoLUbQ2hP1RbjwnNQgXTVCfp72pwFcu9vv8Dz5eFbZiA2EpF1XGgP0JPkq+jIT
s6Tjt3kTn0PxES3nkns+vhZnH7Hm6nI6qG6SnLI+jDgisvVKyUkjX3m//YVOT4gsoSAnh8Qq6Pnl
nymnQuVrTRmyAQ7vMcDo0PWELo7HHKJiEOoQPUs+Hjl20OlsKIRL406Gc/hKhTrhx63h+F9vTT/K
jXQHS07L/KEamHbsmt9sGhZ+cEUbo/IlxJj7bxTbtxXsUsW8aWh1xGYniQhJXiJUhJcpN8TmJd4+
EuFmCfzShKqHrLXy11CifjfF4/Y8GrFlVy5iY0Qm9k55ZHS7N9CUctJAoKDyEZHvXCLd+ho3olSs
RBOQ7j81sR2ffBWkiil1RpJvFqhW6WcFWxdm4HSgFWEIKh2EFQjD9jNSpK8w7X6g49n6IarDykJr
eEyuUbMROe2/5NkAGaEljN9o09HjiHmCikikMm7jtl61CXBmNrWFsUxpH3wVnMajEHEEec0f9WTP
G0bPOWoCeKv9x41IpYaWNtwlXqHVv6VyuADojMFFAOpbxKMUO4OSo89F8JdB+4B0g26gfTMvB8Yz
W5vwdyzzfCfio3Bt/ySTaOHj1sMxZ+84aCHqMO2zHC7QysUyCTZlxjCaBGIs+iG2jPFMaBEv74Qq
RXlocZwPDg0vmmUUt4TCTrE+Tol7qzQCfIN5J4Hi3c2zUIHE22rccXCH5pd1vQs1nkVKLketChfC
QZT8o3XJza1h0rNQgPyCDNDWfxmju8hvqPpj/Hl8xdZ8EEkMblmSuOMBYxjI1hYeGCCr6vMCNjt0
TCxTA/+4RmGWT8JhAqMAPok1+YEGFoDfqAzJNksqH63gbR8dNg2780Q24hI8ihu0tUtICmKjshac
c6Un2dUPMOjRU1/Cwjbpw/jRhuXE2UhkT91I2FnHum0tl607ax5iLkVVKSUA/JITc5xkNH4r6kv+
UWdo7rOox+D7LNzljz+CItjZ+z0afnxKn1Y0mckG3lZuvGuNxxRHSSUUcfMaAMuTU288zwq1N59K
b7skoYupWMeEsU2tm5107BeSODmZRwhfXVTq7GobIBLDDXalaYCcjPq9n9fj1w/0lq6aq9IrIqFg
1LPLW0AoWhWQTI75nQo083VehJGxNfaKCskoqPiZDK/YGiS8JVZyaZncopVfqmHTQNB0CNz3CHmI
0ZgNl5soGgv9ldyAa7trCOxHa/TuzySun/tQUky/Abzp0kqca/nvq92Vx4bQxvH+DW++PL1B+uSG
fjq2elbhTw3BLm7RiO/wal97KutS9gaoGCKeW6ZR0augthBmVVXWEIMRog4UtEKo0a7mpYIDr0s5
UPpmIVnkFARt9lU5iYIyi8p3GLFOhxllEiJN+kXP9yqS+9gTWC5+SSa/K37vJvlCLtM7Lk+dzamN
aUJr4uwnrH0w2M/GUDiKLMyugj2OtihrTPOpvEcuiwk3KfPTxk4Jj3tl7mfsLQAcpuE47gTgC2Ow
aw4YXS881yPB10Fe4Hu7lYTHU6g9YFIUNl5xk/whSjDw7p7Bp1q9Bfi7mBslOMdhSygs4HoR191E
XqM0X+6ltaCnr8iQ/tl1aQRqEdYwrXS+85sCNOKVeqPoAsryxWkEfjRA2ZWtDIJXSBHu7GwvfzW0
mM8q1SC6SPQyQjOO/l5fbtHql5c4m9hGrX+li5QPLW8cFdER9DZ7GWJAo5spsgu5bb0WsAs4jfwK
8sQoDOQamNV4nY0ZplvVYMPWgZlbH4P6wfuDQ6cc9BRkI+wStaKb1qQiJAz2r4VdWJYxT/e09GmN
H32gNcONe/K5zPAD6Z0wbJ0IpvJ60uc7wpH+XaTKF6C71fkOLTvjhxRyqfiH8SVswTMk0qyZY1Tw
QfRcANww8R1KOP8W3eTsi9EC1lzsOR2CfXaFrN2gsTS9sqIaG47Q87VzyOezL9bj3wkFyPYJ9gQj
F3O3b1MAu8ZkR+h1LpGJmXnF8LiBElg+P3AGqRon/pOB5X+YZOAj17g9mac8+r/XNewSFO0o0urh
pII7JxrC8zzVl/sb+iUywqjlssli4PESSs2k0t3rMxKeFvyFa+CYJbF/QYaFqusKjZM1FQelO7iV
6xdb4lYq5l0XnK4WJ/iaLM5lB/injYHA5ULlt9kF7fxGZgkCyc9/lkFIxSMj01dUIRbsgm4u8h1Y
ZdC7Yl925REKSVpABdOvXnXQqdfMiWvQYxc6ic0ZNB8v0519elN2zP4pLzzoJsUkb2OLT0tbAAGE
EYaad5yXNkAFCRZk1wtMsMS9WOe9y5AI7d2F5YOayTs/8kRerneA4H4gCEOLetwahKmzdtgZ2o/N
p8icmBMxT3ZDds/c/2Lkbr8X33F5v9ODcHmGhzR1qW9CDzSeIcSThvJ2dJPJK4qpm32Ge9T5yFQH
9isc0HT4+i1XE23W9aZB2a8xgR8w8QBWtuHaT6X6Odcrdicr1y2MU405JXI2Lkwpgc/LCdQaYIHi
VHO8IweT7Kpfzgw0CVb18NqgiekPc7HEfDilTyBE0jwcBFltL3KtdvJPAaTHsGM6TkvDlNPK8rYK
7t2JfXRUwSy8s2SIfovfNNJEcqWPNJKAOJlhtiDa/EB+dEOfF7aD4JGK2j+wcKA96LZdAU+RFVuK
6Z18yus7uDrPGYeC88nScuxq8xNdmCRZHE3fcik1GzSHXmcFzkZBa0tLq01zOSzKXH60F1N3Kdu3
dRra6L3nSdolAedaNMUZw2EOofFlGuIcDbDQZuRA2Ld75Q35KuZ2gAFiTV1htfv1i/vDPI96PlYo
P3y5YYXcHZY7oYDdKN+Y+9G47TB23LrJSqaPczgFCSN4cv4cdoK4jf9oflblSCZK4pAuvsmgnB8X
ysVilnVLFCHTpsvCgWJhKW8LEvMrdkoleRJeLP6wXz+O0cbhMLci+5X6m4BbZGtBUxDqUApnkTSI
b5Btj01/d0WMlZNeTLhOrra/AP8jfHUlPHlWPxyQcrrz+YRYBNQfjzIkyL/w6GTJnKDB5vNwiY7A
WrVVYhohZYZ5MbhpSnqw5VlzriZMspJn006Pm/P83y7oIQQkZLkQye6rfTwlxnJ4jBdH/WQGN6y/
k6Hh0sRSFuaeCCr7fNtW2ZizqdS4uVlfIPR5FZYgNhC8nbEHPviGm1etEWvvvA87xqqI61obqvFu
7iU4tlvvfZz35WvjYbBqSfKBLPBI/3bcGS6keq6pKypc5/TWc9ZkBrpRr+QSrQh7G8MFCmqILUbS
XlED+wMwlHfq0/23+e1Wb842w1/0lfTQSB5cSjtFMEraxirTJNY47ParWpO9v2L1HhBbB/3d3d1e
NNhYah5crNs3ErueMAkyDjjokbPYLx/m/ptt1B08bW3xFQPriiO4CAs4IfBppixnR6k/l+Rk3AiJ
a2ARRT/ZAxuKrqRDfYp8FRtmgZ96mjPr8DSRIfWT1fF9w4Px+byPMea8UFYgvBw2olxHs+K11t2a
3PbZPtiGDEYknh9HqeHOYyJCgMILcDnnMmvtlWMRZjDvqqRhKL4VeT56mW5XEWVhO+eR3Fqk9wLa
c+msQ5v9h5gT0/iZhBuDLJZZrKajWxeATnZrHF2GEhopflnLk1K/kONY8xPrJDuoPm3tTd2jgbnf
y2XKYTn3ueRenqaVxxEE2arzXQkrP/PRAssYk83oFxQmme9R3JrayUhGzvhwukpkpM9Ok1zDFjom
J39t4Ao8mm756+fxd/471IOPYIPD05BahMBlJzDzvwE19CVSulU4XFoUkojHXgnvVnGXnNu76m6e
hhLTWXa0XZb0M8Aa5CRofUspuP+WxDBeUXPY5wMsaMvpFSjLGr8Uvf4xTVjKIts9zJ51YRl5Kfra
4pr4z2K/nk0GEdnq75QOXxKsmSBEdVB0IEQoXWvUPBOluo1QSwXFFbb1e4fDQYw1LMmmtT6xkD1S
rkO1f52wPDen6T5uY+CEpuCbKmvSJs+MabqyS0wWqCB+ePq2fm3Gnm2s6MmRpMwS6RrRDDc2qw/X
QGgktWrn9Wd9jIHZiqseEjcFX3lXOAh3JeMCIwTenOIh4djn6bULDXIlxYgdrsdvSxMVCabZVl8X
U0WdfEbLssxNVZmvYpIyklqA2cHf3iApOxjAIi7AwCJPBwGAhWbYSsKTXq6UrqFYneV24R/lGdms
fyurnkGAjtRyzTeu677/5XxsyaOqrRtJKECYxsyNAuPITcddXdY1HCXojQv6iuGa9EscsdPxROlE
KHiinz+cfiOuq4r0oLuP3hgEHFbDcFBRRVEweju9FmvaG0HZUXFfMTchDGBCF8KqFuZ45Xi6RpP2
bvlD3CLxd/VD5hrP2Y/blx5d46ntbLoj5DYz6FaQbxZUueLRu3iJN8jzn59shjpw0s/IXtbdfuoZ
Cs8GM+pKTci/6knQ27mAwQL1py51U94N9H01GBXIO2RIH6+k5U1a23NzI13G1Jq0UplfZMIHmh3V
LsK+80/zR0P0Lqi7e0+OmY/6py1e2FRJ0qzQqeq1/QlpM7IGLSaqf5uAtlm9br0OCSt7jPXztuIR
ykwLL1G2RYlSklRZBNmHe/8FFFO61Z78wR0ZomacvtJ2QyN1JmE01f6HpfMOR21ynP4gIXj6MuxF
T9eiL/p3UDTh51ktHSreQA12RW0CwPruJpWHZhSNWPjLwtFKmgRdz6I6Cy56ByP5kBlv7ENcukmE
Nr0Z8FmRuahFUQIQRHIYdlA5sfk5tLVSyAkNS8ijMn4Phrj4xWtp1yYhdCrGOsh/rgOnz7O80H/n
KWkxuxacaM67ZEFf0YMqu5bArPvS6SzZMtdx4FAdsgTablx589KuNOfp1i8Hp5Zf2edXONBoCcVz
7hicR3K7EeIMeoY0FUICgkK6M1sMN0mybVGPlYY7R3+s8S8mJTmM0YoWy8fy05sLCKCCwvb/qOGR
4LEXPeI8Dz3GOSPv87qFfSQRTlGETWu50231o/99eJbcc/2joGAk8iKepBWMUpgHVVF0nazFsceF
ffKB51qdPCjGMm0rM4NRqXyurUYWryKvt6qKbRj5zWEUx9wAE321fh6b8Eo6cSSnLwJJDB+I7SmY
KA18RmV7Yi+j73UanbAEcf4l2sWMyEu/nT05hvbVUnFo25fvMPHyI4m66CxKwX4PSXD4cUfXZgV1
vhs3tH5D4J4bbTbksS0mIAjg7+E5c9FyZZYfI/Q5ndxXnsuyZB202VEUw63zj9vWBfEj+4bQIUYY
LNTjqPO3dh1Y+U151c0Xr0z13Cxfg+M+rww2cH6OaoMPMhA5Vh+eCoI0IzbCPRmhG+RQR4Z1c7dS
A0TIXPKB78TkK7htH/geMwFsy1e5GoT88vRIG+VfYXGBgNVTwueJoVJb9tRvwvN+/q/PCebunOc8
OvYlZWNspmUplfk65XKakhJgrjUUtvPQaTpoBsdzr3uQEC5BM5oPAceW/OMfbLkaDaCccdoNlsSL
Y2wVYM8R3bB4ModN7WOa6d+Cn+bIxhl8HWhbDe8REnzNSNtXzZX/V19xLf55Dkr7fGH8KhHEhKgU
7PWii06Ua9NthIp5Xx1ZOPf3C3eJFob9v5MIp5FZBnBfBf+2f4yB4tGlJlrQM/9KVEBgJIwbpBec
Vmiu0XAZ5gkCQGeGHNUqHfPWgyhDRlZ78cw5z+QghizJIlM3z8Cy70WjNGa/UAx6ilaB7Rl873BX
/kvKh/vMVlp/8I6Cjz3a855UfM8zeDluxNIK9DGchOa7WHZ8VjZBWXXMFDRnYxDXUI9jF+FXwPAP
GF/j33JWdCU0yajuqBpu0i0y9mbsNscr6IQjLLmyqjr8/H95QCcUcnvQQl25lVaPnkEkCsv0P4eh
yHimLXcrHy+noeNJfeLY5aUPWf4zrOAJHbJmcmEFIxBJceudyx2nCH88MEdauouJOxXw5oXOtja/
DOPRaFUBmRzlYSvfJkTef7EXsYloJCY/Ilao3bBhoHaWLo1aAIMhSDXlwfcpvGLGpqGTCDGo1x00
NIXfeFt70vWL+AWbXa9yy7C8xTKf8d/CHow63nclJRPXcm5Ahk7ozod9LQID84gRDJoPWFbLw12h
cbxPSzgWmMmslRv0ZpDFSHDW5d63tFysODX404vPw1SueP2YLzxQDaeIa0WpaiTGfGzE1CByFOZi
rBKxWnQZPDZh15OuX+EaboeA/mdYXfpP5bseIlITkzL1dQ5lyyvXAV87nFGkQJZdYQbufEcMzXE8
CxhbqdXHnOemrtYXSybZ46V8N0HnMOzciD6UP/z5noXJTyGT+hDJAwsJfo1tL2a9RUsMx3fFDEA/
/hlE+gT2EHUwHpkkYqILjwF21ZYoF/d43CZE3pcUwnJRYwFvZF36/3wfULQv4PFYQSD4dXGbWMyB
BSkRPQjWeSy1AquFGOh4QMKZQFBU0f5CLI/r1Thz2bAxzzGNnffkAXhxjCTSBcH8jf/NatkVDSWh
OBXD05IcObToo04m8SG2lRNw5BXhPCOHyX6OBvAAgSEDZHClgp2BkHmgtKHZyrq2yM6j8lut5Dvq
OWNR8ZVTl1EtUVCwh6HDFS+MTuImuhhv+8Yq1LJnUvm/WNI2GwkQkpM3CXrg2cQC2fneEMRbuZ10
hbdi2U+iq4OEsfitb/LYo8TG/HNwucbO15TCttiMR778T0t8Ipfqh9HaajKbywWYzQu+3j7Lzusp
AbJuB/xWAppXa3iMtc6HWqWDrbruIixds4cPfjSRy9ReZJ0s0bMoEjJE7THk/3Gpydvi/HmvvXOm
3cZGHqx9I89jUNsCB53yWKiBAKiWPTcD2r3cXYZaIrMrzzv2OTyHwHIpOWMS0PkDzUpdMdzMpwHS
liMH2pAWm01epGz4VppwrnYZN0DdC32jd2IAsjHVMWm44VwaINrZm6tBpVZWUiZ5df9Z65ecU+tw
foEOO294gs9TFrBG7w7kaD3VX+OP/qA/dtMFa/e9qhksPmm8ngKdU2h0sL1vn40SSofjoB8LmRth
ji6Q1THo8GlWe0kTGVYuAhS6DBZj9xEgTo3JlXnh4YZAwqV7qNTuKaXvWMB9WqQ58pG/wjRYSU4b
uyMhLEo9QwIYXpPp6iDUdYhR8PkXRWJ/Odp3KK1uCU89BGnsLyHLTQMtlPoyUZgDxyXzEiW9BpD6
UoNF4LcHh3bF9DQzJ0NXZ0cpR1LeGx8gvuTImJC4fOPNlOT9ouclpYaCtzNN31q/6gtarYbh3R9F
rn++HAvYAOer/GYODGYFJ81BxdAVs+zGheMOkpTN74aH9EN6Yoj0rQoxQTbsZmS8DAQf911aK9qf
Ffv18wAb6Ye5IbdDBlKbcw+NuPvclX67u831iiXeRj8L77AwcQQIP0pKSngjUAzxt7NZqQuvcn6C
pdl+cyTobw+gdsy9Izx6sdjqM8ZbCufpYRcH3lNn7PmfR3TDwItrNnGCButO0sA6XhQ6pq0AsBJj
AW9e199RDvyz52haQnbCCqNUjTQ1tg7xBKGcAo1+oMueeIumlfp3fSQrQQK2qQ8E5dwNwxbMXrFM
GZ1BXJ/Lidb/TnGL09ktD29+NLfxfurff8zif4SL0x8oBbvOcfTAFtckyG6HnPvXKMG60nI3rxUs
Sx3JUxIxVh/qnqu/CXWn+oLnbMOm8JfUmpSPBDkctBC39PRvW9P9kHmc4RoJZMYkonODFVLyp02a
hHcMqhPUGHZX3gLZOcNPzM5FEe3D4dWv4m/Tg/zvVi2V7SO9XPJZhOWU6zQoUCI7QhHC5GlpyafD
BvkGm368AknnyT8UOJmkW1K6PKuYL6PlceVtagC6Efb4wCxt+0Too0PoeisLSlsufMhQDN+DyN90
YyGfLwHh1fuA2AaRUbjB4+tKyXeNLbk9HmhZLvskuZSO8PfcQadUvLRkKwV/ueUPQklNshzz+mOM
xXYjA4tmg4kmhPg2y43z++0uzDAnrWJ+eOSslSydFCXCo5qnYoc5dJqZaXHfuNqRF8IR5TIa2QnR
Alspa3EGbb73rRFe6NUtE3/LG3GLmfy63LPPFO/HFyYCCB66aB8k0eFfZ5MLKbhjREBLvzTTbd4u
vGjOab1VAZbrHjtCP4HwrhUxM2TafBUWBed1A5YnCQLkEsWMIlYZ1Vrf4NUmdrj/YsSIMedCb7Oz
EtVWimOk2QQMq8R+Yp/gEkOb89kWaRPbViLKT4yCEpdNFnf5zAlAZNsRv6aFNBGOAmlHnNhvUbGa
JvPGHOLhmrHI9oX3Hq0LYTdq2fFDnyPN7KrvKLY1cXW8JuzxTlhQW0+7RMFtIrIZ/yjlbBziy1pt
al8Zl1NpUbqUb3XWzM20vkvsH3HQXM9egc/svtCi5FPtL0aLiVZX/JBrlztkgVq8jjRDsKoa/0lx
9lSPP9qPbqjmj5+yaFJVHpcivgmu5yL5r+Jk9dHPKsxGW+Ac2TjJjDMF5Jy2uz5yqiC9c3dyQ4VL
eZ7zNXlJmlNpVmcbHClYokKrHRMwUSLN8Vo/H/2r9XTf3AWKrxlUeCc9bM8XZrpgzcMcyZ6sQt4a
svQ2f9jH+5rua6ySqqIiacYPaCKSX4qPhSFxUUGQ7fhLcZUAU18C0skeFHMt2ysvf95DYEsC8gfq
14ukPCTpOf4JKkE017lQj9kdyiA8devOxCcKn624aWp5lfZgOyA10wPQY5lYIIukE9z38sUBlZ0M
JnCs7wZ9havjiqaNDuX7vlRCHQDsrk1Rebs297UbNbjknr09i0H5FReL3aV36F6+wAznMvaOk6ds
zxgHMNo5s4pcAuOMv/6y471rpzW+2yAmTjdov5PuzTSHMmWrhTsrZRxP5mzSS3SHWLyItnvV95/X
PxoANCuK7a1QZ07IqVO21FAQGmroy4QXm2Gt0MYpBAvf0ksmX5Eu7KP7wEx/GbAsSXG4VuwP8UnK
5B7oAjB6ikwXXqZAOZKHROmds9H8HxR5QxykBfqwmvtdELlboAE4T1HbBdZCL65gIJbnVA9lIf69
Mk3k8bv0SvSiamRIVxUd3tGHWh9dl2DAHSrU7HT32jbCkOj11M6Lv+kCVmgPKhsmdnSjdhfD6KHk
RhZc4jqEJwFk/2reUltrknsremIDVU/L5EYf6ONAnMxxQ4UE9mZJ2I26GLvDFlcThzSIpVv+fBzL
JZszvIgU80vCcydRTggj5isqHFbPf+Q70IR4a/yXX/Wb8csPqXlKvM4uHm5qBUZgaOCtwT92w8bs
NqbIYIv4os0CO/PWtJ91ZJvTd07lTYRbUqgt838N8z2yzeeHY3PUQ6yZCg9sBDzSl0h0wMmwmIqv
ON1EqwYnnJw8JKY8Mk7VyngN4eTmGghEU0VcllxVLUaHUaG57qXVkilPf47F1f8Q7P6NZg0oc9Y9
InNAlDp5SkXXP5mI3HJbv19zknpO/3m4MtXzEW26GLCSGGoVNlxPjOlMxKtcIfvYyahNQ1ZTte92
ZWl/+Rwy6LMJMNRSTbqSZdMX3xGRBdV8aGb/JV8aT1nYf+6loH1bk9jW6yl7ib9uCoV7QlP44B7v
rSXJR4OjuKB0zKdwWEZuVX3js7o/1A5/p2080XAzEQqLqgVp+enUvRh+0tzPZWXNWJvCEem4Gqu1
iLI6qEWZnWeZot1GyHb15fYdmhYQ/fmsSiDQuCBXvVfyYdwyppKH+uQBaPVTF4AVC1qgOaewQU/l
Jpard80+TyIhwZUam7Nf4NFdBTVy+Q1rMJKX5anKhFlOcaDTMQ7sHNDtiXU+/4DqdvEH8f3gtMLC
BSmrxcGhBMFrG6p4aG+pG9iTmb0I6PNrqpL8kw2ZSqj32uEblJ3rIAsU7qCzMa0K2dxPpg/KbVZw
IAulFWdmBhgaBOgPq1wver0ZX/hIew6N3ZGIP66fYB5621aNkPc+DrgZJmBGRKgPfjNO8CiYyQHx
MFRehLJyMKxw1vLKRLjOlI4UOqcpNFoYcgYnglp1NvAo4ITcMVPY2T47y6JcJ4TiQOJQLwWnoR+i
DfxHzfq/wVWiK/Nk0gmvrA9QlZfJXuvtiLtM2dvQFHZkAYPYuvBVGOmkRQC8RTu2H9RxzW+u/U/P
mVImlj1G0o1YeX0IrSEjy1thIg7bpS5Uk67WlKVkVHWKRZu1UnT4KpqrLmnsme+7G/oirJQ6wgCM
Wml1uUSdRZN1S2YiodP875cw5CVTMhXanAQz1NbCKNcEmcyzJzk9H37/nXm00cldFiY4hVCToE5M
QaTgFAX+FunqqZsVBJFtsKtS6Z/bAvCX8DF/ENyxiEK3t8mRolStmrR1rTd7KmFzLc33fcxoIBkv
Hk08a8WrntEQgjsyVhGR9i6s5Lqqv8QIo1CVncsWHvKp/oFt66pKdmF5ZZJvp0GQ1X+hO+AE/CH3
fW0f2vn16ySoZknMEF04J6GjYtD0G83oBBrP4HPwDeA4B2HsX/wE3Rs3gZ3zVIfQXX2YFteIz7nh
kiz2dSqMMgz1ceI75oPtRohgR5k8WtO2cCuGDiT0eOXtyvuLEfL2F1EDPQGeTUR6+rMeQArth/NA
NKWUMbeEFwKB8LKIelGtmNaPIoXShhq1uwK1W0oD3qyERAN5RO4v6f3rlTg6GTun95/Q2ivfb51H
QYg816dX3u12cDSyWqMmUkhpCha7i/3+Bas09/Z7qHU/+Fm7okwpWuRGh9NpIa9g1c/cjqCTkvRE
V36UL6R8Dl8D1J2X1mmcwKFCiovE+Lj/8k/I3Wop3NmZ7k/JwPglu8NbkuzVqNVaRWz4Nb33apI7
7cOTN1ul6OCOoVcBl6TTLOl0E5BDq6pNg4iofnSOMfJlr557PejbiKXLZDPiMjPEA3Xpbm6BVMeJ
YuWRkH0wyMGfY7Yxfh7p/Zl62oW6Mh/B7gVJNc6Z4pXogPQHsJuAcJnpCrk1vDczJUbKaYOtq2lA
p/kQ5k7aOa7b7Bing5DCMmmTZh2ezj6DQhpNo1hqCzazKpaoNoZwOtd+NDBULMWuukow5+3aNthP
rDhp4gRPqF3milONGTfwcoWPRjl70rNxCSzzOcJvc4oPD+iX/Pgm9NjscRFsJe0Ut3IQsV3phXsp
c5vjftwZkGI4PXqCjKePk17PVH9d5dQJiLNYjVYqFcHg7ugRzBI0AUAm6hURmzyoKIS7k14RXDDw
pdb6pP5Ajib5WD+KaKN7TAHXx2sB5TJllNcPUHkZZw48od+TQVECI/WBEMox0aJQCsvkawRYFb0c
lIosOqNRscdKzqrRFHXapQ/Kw9j3nRgrIkcy9//pvWCyBq87mNtQFAFBNm1hwOz/zWdhvlBTh9ss
q1flU4EJAnUSReYKFqG9j825wMRhILLzLe7KMY0sCack00LT6WAwT+TjgbBU8oghfOlCRnBW2jh/
2vPF8/82KAxVOL6ucGufeYoVRuAwxWW9RlDyZIW0BrVdPOh5Mg9HWjzd/K//GaJskm3v85MzsQha
BCFMyIqfJ/DYYkM9Mtp6krt19ysn+Y6NSN/Ofgk4YOkcne5BJZJuM6YKjeup2DGT+4L7fgDWe1sH
cjzWuORjTRfj5Qu6j1F73iWrmhCHtFUycTkWl0V8urbSCVm0+zL+YVzPif1hKIrJFDixnbB9rjO4
mtVZyQKkZVpqop33EQr7o6jHSKmkzUYsAdTAB09N6hnEDNNGbk41XVSxCfgd0IKrIdZfDF05AuhA
ho18udf4AOjplpceBVl6i3Tyzo0S1tf8dK5RLypllUqUYEnmYf/6bDQoGFGPUJv/KEJ2vuXLRvUj
bFByeqMUzKiuoDzTmgFPpZKpZQpgXyAWdH2jco/u+dbkWXDUBDy970epP+iyZonBpORu77VcpEiB
qYmcK6lrlEY1sBF1+6kfXUi9vb/ZLQLTnOwUwvvRm70xXEJw06vK+qLLRa1Xc/Fjjmydz2tEHnvR
tg/yblae4TybBaMLn1GTJeY5pmj+sFEI6JUwVE/UM1klBF/pZKBn6lsertp2utCGk6m98tBZIyZh
vZrtM1iuciJXVhcC13jUYnbPKl/SY/SqBPNDrbvrLiZLfTubw0s0fetuY2ceHfSu+YcHVuDNTbYi
NyZwljQuHim9xaXp4HhdWo0AWGxAIsWYPGE+3WIcSsr1+ZdqV9mHNNSy/ZDOap/MovFGh13JFjOe
4G3B+1oBad1AoVjtUbZiLFGZlf0t63EBMSh0wXK7Dr5ZXOJbjwbw3yQYpaK3wAYDiQwsFqg6S0Vp
N96YayP20DmJRS03gDH1Vfdhgp3acuIsz0AxCniyutiaF1jBfdsQ78Qlqsu2NfIBnbwh3QiUEtfw
ll+cn0onXFDtqqKyCHGvX/AWlR4K/qgzl+CnJX3SsBBgiP86yUI4+rs41lETqSL4FmpAYioi3JCr
rvJIh3LOwKQ0PL6p6uLwfkorO0olt6qkyuO8ylxd8LBPDmzdcPgHEJMDn0ipdwlHTdEk2kz2QI1U
LLME6rVnWX/VDllMqzEdjATcimWyzvR0A517yiQFl4X8IXWBWsVAMFvWfXUplZC7o2gdfDUeg/5e
8/KLg1ZKOqXskt5o8EErXsBP037cnWBtu8KOBXE8/XukmltTdC6m+jIe3/dZQgrPzmWOFh+OBDHm
3sEnjuuz7XNmRYhMXsXPvWzH5vfPHjLH9PNPllymCugaNg+qT5QytTTvX+3wjjtupa0juF75NOUh
e6SOOxJB/NYoIkPG+YSl031rbCq6bsw5M5RtT4ngcMBk2TtgWAVpTIUU5WcYijiYAYXkKS3VxD2M
1yu0FR1OFH9+31UNcVx8UTm7SwBJEOW4cq2mCIqBkzgLC3y3YqxaxGww88bASTElcFxEMHf/Dz/1
0dyyvV0b9rr6V5AL8bhVF8sYdUFuHv+pf0eSSNNEfIjfmHEhhmjAR4OdYKqa6Qxw7SJDrY/qYS6/
H/K0ewnu5pJKaCk4sUvB2MFqLiMaNpjJcMOAt5QTbimDJn9RxIf/tBHgu5mVDucLN7vy8gL1R3i8
4PhNYZHR2jigkYj/ZZpr2OPiBjLHxdPqScaq3jX5qgQ1pifp98NKRFmPw8P1igOMibceF4OhCPEf
TXOKT6f75F3kyHT7xm/GzJgIHzPY1te4EuEJUNv5gJNmktd1gg3h2HzuVWVxj7i4Kvb0zJJv0r9k
J/76y9oiMcRkWphL/PwMaSXSyGdFonu0PR9iGRvCsIncYTQpN8EeW7XnAjmb/0MFc6rHNIp9OUdL
9cEDBqUd+cgpBuATMUk1EuZQB38oBtz4fduVMR8RbeSiJvnJqilAdw2Ls6vVB+E15upg+9BbWrWV
fTKLfrZidX0yRqBbLdhcRRv1g4pQLOlfQdEvN6DasU+idbPUgYSa+QLBa7GnZixMCHgeW0iTNq/H
80RNcFM5Nkb8r66wZyD4+ozfJ/PiDVMS02JbBcfB86OAUTWMFhDXvw7l9YAM4/FbhMRLb6y/dU0R
GV/xV7EAgW0yiagQfiGLAU+nggZfGuHpQYEN7tLL7ehgXHSnJYcHjQvkphCuPQK8X581JUN04py9
wBVWoK0s9T4BjeC0lBafPZar+fCQkwtQCWzz0nK+iU7ljycjt8kASZBjR42dGA0NSXH1mCGD+oNN
epggAdG9bsQl25uJKZzWTgET23jl7njdFfQxPcm+Go8FoAxprUdF01L1jvi1fd0cGTLA45aO9vxo
4BG9KJxNb9+Ve/GL5FTQ6UQbLBT1CD8ah1gOfaJhoT/a9NMkNbckPfatM26q+xXzfBccbE63z7v/
QK4rEG7MveUhy2hQ+hV4dUqH902cnBr+WbSF+8c5qCa91WQ+/VJSxZjLEnqlX5/dESsZiMHazYz7
28KfiGEoYeUN6hxRwkw9P9+z4e/PoDb0zalYV1e/1IPcRTmGCHYEd+j4JPNLw0O1XdUNe7SUulAl
mWciUsA1PxbgdhDaWXrRRHK1sujo1kcZDa5XVACu0vC/TAGzSOFrlXfpTRwKURFl4KqsHtJoc1lA
Pun20qDjqMZqwfMFcwjosRlooud6wyuDuGyaiUsXRipoFQWaD/lGuOHkgY+Xs2BSsHsiX63Mu7N4
ntD8r6symsVbdt/Epmb2xtKy/5/IfvB5wW4T0YPuSskq+wC9Q7WhdkWfELd2vOgfG47bGmas/Y0m
u+CJJTFi0kFWDLn1JlGY6dGHIRWTFmpxyHjrWqLJOoYcWrE/uRSSCTvMI0PGPsgi6RzTzhpskZfm
xOjZp85wb8jX3AjaJfuga4bKRFFuQ8T02jzAlW8E4Qy4l1DihWaJX4TQPqr8knxwAo/bVvElQn3V
1Ykv+ffpB+412QpivyeQPdFKnWnjmSbsgFg/BGbs54C5T2B2UMFtioXucpZMCygFWzAGjJBuQbAj
C+mwi9x1ofXmlxcGp1YCpLGeLijFbkKZ/R/vaxPJdsqXz6VUvp7xJ8ZV94rCO4fg/l7jPkj8QPmC
nisXAPjjaamfqTZ/1xf6wGuCXh7W0d9PHMo3xYP1w0ayCV5A1KXpZ3OmFdXROmtorTffWvp+cTx5
6zPT4zKz/rH5QotmsIvsQudksDcnbvHRfT1Qy3cXZfw60aav9bAUb2W4qf7Eb5LGmDGOGLnVw5ES
5/yq1QloQ2yR91CFjmZ4OjAC/wdhRMLRVzY5RjqdWSNGkSO8ePi18jyyQy25y7jGnp8g8zjv6jSj
7k+35te8Kej5n3ld3zy290wYa8p3uzzFc1qruNKC91nWrahyGAnb5k0YLBscp7Q8CD9qJqIo+f2T
GTBUD06l3W7w/XP6mMvhJYv15J5X0WllTIjNfSaHLeMLqCDPbT3NkYAWHgffKj7UFd2fYQR80MGJ
1XfQUYdimR8Q1fgNrAVEtkzc9twJ1EEwA/qhRRCnXjDOBX5a6lDjmNTht22b3kaOhe18/wGoJVeY
wgZWYv/uCK1YVotAWwW0qgA8S6OlqnEP34HZfyDQgn4ZRY8LFhJJ79aoMziLUI0QUtNNKNTpmtD4
fxWADrgidia3OT2cvgoTBHzEiOeAQqZOdyi0KrFeY+wlGhGFoyLY2ATak+8TpKk7lXuHFdRy5J3q
6MO/TVeGUxI8jydK54b2tBHvZbBpjnK6zWNGdcn1OKqlqBCdBOTT1zWwEv+pvCYk4pC6dkkmtCIg
3qjoMRm50SvhdTzewpS8Xb8DZA/3BiYVaLIgtCgMP7LThkudTDQtOEj/cLqXIEn7+PdrXH07H539
e8mPv2FA1WiSWAfJ3s65gjYu+czIXGfhuujpEfrBNZRP2H/D1+t2N0jogJNFHLRmE+d0ZK89J6U+
/mXKQyE6QZbGaaHOB2w9mV0ebcUiuWwhD2ro6n7FybaJnqj5ve43vXS+nMhYi0J9Lc7zP05WZ4Hj
dtWkyZRLXnHPmzapzDs+RQ8CUyvBcBWCsDp13ZBqlYrkaZY/3Eu7aqFUotGYw/d8bi/Rh8UNpGvX
ul/Z0Cpcq/TapsKBliwtjhCc8RgRIrxYA6dSceBYro1uxVvzKUHXGwUaU9Z4VFsSopFoo6ajqLF0
VPKVFJ7LbES6EVgeW+M53vmLrfgcrpZz42Jc9g7wMDwMWGrAVPuN9pabOPNs4eoGuRQj5FEAz4+8
lUWhRM1N3OBpRaOK6XyE7l4vkCURG8lanumYD8gvssIQZD7s6ttlHp2stecG5L33IGZodlO2P6El
Z9nRq2+jZAe9Palad85pv9+/dQfnxWYwwU/w89i6XB/eYkDaXDpedtEwRs9SuK5qX0HXaUKBAr8W
e7DWrU6R8jG+5ovgvHQGMkA069tF1FVv4zjldoC0c7hcHteg8p+EAP1eJQStfjZUZdYdK0CUMbX1
i1l2D5MCf/rJPktHRgZFwAmThPGSEtfVrr1onqNXYfvpZ+o78q/qVxJ2lX61uvQfmHbFVCfhtBb+
rDaHhPsp+82ZeiIQdM6NMLnRcGZfLEmlYa1LxgJ5NHnOm/UQth7BqiqxjkMLJUw8I12xbze/GCE8
Sukn9J6s4J51QClOEgDgIqo0BhsB/AbsCZ9CDodB5hqJYm5i6Ojv+SvJC3zKAoae9gl5MO68qwJZ
PbqIFdxLKe/4m/yyPOUOdJo88FAN42PEN/DZNzV6jdfEA7M9IwGZN2zQzwKCnTfHBKqxG62TzPtG
+1EjCvwWhjDUzme+maExwOx43OS5Oa9GlGD4X/W8Aa2j8p55vxJbSUxHJEFTqfzFSL2nc3jZ7PK3
oRk5BAq23p1jnjtXkIMFVAwE5IyoSSUXtaB/mAjg8BwtTD7msPyKFHBAkIszUktD6S6+t739nKwR
GzhP1TAnJ2TbbhPmpXrzta8/zCP/7SScqcJ0q6U2Af3K9/Zsf1HntILlSEnZRMi3N5cJPWbuZ2TE
/lnvMC9BwtPEtLn0L/pitTWOqgV6XtIGU+DCI0cU0FjgT1b//dopU0AqjiYpwSL4rcjS60cSZQnC
DWJatUGvtXc9RBxotY3fNYM5LMzIsUDa5lERtHTrl04ZUhOmPy7bMgqxTmnWhwU4BCdku9p3o/oB
QVH3MGeUkcP44Fae4s63+LUNWGPogpp7FOV4EmWvERKqvPk+eT8nPoKW6nzPuCfVIqT3T/uT4pBH
k8j3lDoabsRN6Vi4Xovkp10NJVcgeeStU3TsV7J7UkmjsDxt5wC4JCpgPTbr8k/EoRhog9BuXXFu
/yoI+nEyKLVsaeSnev0oqIyAw+h+mcQueOgXAipiHZWV96qI4RebnYj08IzBG4/xVHyXUenjGoua
+eDcioCdkBNnyHPChj+wlZhPdcVm75HWPiVYwA1MncYUlNJCMZhIslOzjNOHMJlJEYA6+a+Ao72b
2+EsNFegXNdRoNIcAjA84lInpIooQhRg+Hmx0e0wNJMrAtXpPYey2o+w+AkYAERqpn6iJ+bxi3F5
2nYPVI1zyzYUfY8EWjBD/b2BMEDinFt92LnXnm4zd7JTNuGLNis3cTGTVyOAbqXGcAf92pVnb/2g
mLmbdlDqdGMM0V0DaqtctXwuswX5w47/yju/LZmmD1gq65mi/WO93n9DBnqM0MJTF88rbK+J9MLS
W0ZwG0hpjFF0dG/E0hRLHCMdDLHV0mLCBpwx1cpANqcXu7vABeB0Ern26qmobgvo2H2am6P/CRoi
HrgY9qJmyoHejwZ6O0xm/xc99HJ/Y9eu2p0ZTvKbbpnTFtjFaKzb1rg+88wcpQoTWhIOVJbe8F+3
DobDxy+6HzsV/Jt9tTtbZrfz3ZaUt/fr/hYaVN0HX0iJJiSjE9i9/84EDf3Mkfw88BKCQ3sXjMeb
mrflaiQlBxaRm+FiwpvkVAHtZzwM5FA9P0UYDXHAnte611XrIYOeJSPmXEPxgi9CbrRdKs/niChk
kySZ7bxUAqJpsdiAIZS+Rbn99cJepHNxAK+HgKthV9jwrBYBj1TevQGVqlRvVGZV5GoHfqgmGnjW
BTxDWD/fdLHKUq4FF/8m/qdXYvU8y/dm3LoQ/ORjoKzl0buMQs7RgTQ7MCwjWGMroO/3LNO+/K+G
HH5YvwdsJ7/BTMJVhhxCBu5c0ZENNEALpwv88GgA7+TLgSjUf1sW+1qO9hAM+PV6+sJHrVCKVydU
gsELYwkELs3Ye1E/cAx6NCftQNv5LaVtf9lZeHJeXYJY0JWXJ+yHFWf9e6sr3U+gJpzT6kp0GBdI
pbqM35mGaT8t2Tsiu5JSnzMfYQOlNzanSobuT2cp+YRAY9nuscDWDUouxA6C/31Pv+2Ia7vDEC5W
xx9u/2HIPYBYcAQEFZyW0bgdZH26o1kTebqeoyblfEpGNK0imKNva1Cpxv832nCOTM/ukdmAqP+W
Et/n098pTkwuTCkmrazop7JYU6ULpjb9lpeip4F7NRgAt1VDzYOtGgSRYjTiiWXAWpGTrk/XDEBQ
cQ3CCh5d2fgPE5V/tHmQRPkPECmVAsD3h4uH2pGMWDTzlQWTOY7tMhmgRh98vIHwUO27aZUGZI7S
ig0vrD5FsFVsH+PTsZNOssGdPaegWI67Vr0cANIvHbVjX8ukiKMGDSecO8nRauPbSodkteL+oFXt
LcAvKw64CtibWe7750XaikP6L0zA2g4IndZIpQ2dsfxbmcx4giGyR8W1QnncR1Ymb/rhI3iDjFIY
X1vGcGNn1zOgRUQDfo87wMxqTapTjmS4kG4hMvCA5hHr3mPvNETshBRaoHc9XrWYfBB/mcO6NBrB
6hW/BEg+3/CnePiYo1EdLo22/wpR2NdlG55I8irIvQZspPkdGUJR9xE8pJxi6yfZ20U7nC+ouH5O
z4B+eR6FdYAABZj6QyT39seA/7Co8N0gOQ5m8uxw2jnxG6qzpGsulmA83A8vD3p3u9mF5jMORzzf
Hn+jNlk+qVPjmIyi/fzF0o5G+S9nBIzzpmaMGmrFFK+sgK5/mlQmAat6IA7D4wicgsdrLDrDGChD
PmcCx7/toVjh/toV3nGfDsud1jko8dItW+r6q8kMIF4g0rwrL/7/yBtl9WyjcggSPuoGhkTw4Fuh
gMqA/Ca9sGH8LM5NyywflUXM6twbif2i6INtQuWVkzinuEM/kwIagSywxc+FE4IhQC2v9h94pabK
nJ8SbKmNv+T+ivmTtSImwqBI6x5pPnhanrxC5vyyWEma+U6o9apSCG8Sd8NAOt520L/+uJhnwKOM
wikPW6sE3T48LPFaRlS0auVNyZp7m0am1m/zXrfohWcH6tMI+18v8Ux+6dPa2GFcgG4VRlIB+BJE
UpedeMReEuPAQU9sJU9CDNHdNp1dl+HhNbrESXn7/W9mhY0QZwNARuQ9MngnIa6ygwcznuRoIdX7
+QDy62PaUw9/40/eG/7hHv4M6zkqPvecsi4kV4iBKw1eSfH0IvKGJMXEtUoseP0TiF508CKmQQRW
8lbQi8PEN9wWWJndkOWvR5GKu/Ho2p3TwRRQSPUsYWhyfWgqZmaUgXoGDamIDUtvhLtvL4jLr4qM
vmvflibFH8ftpSjmcbcuOmpPVCPO+CFPHqgmOCuMM4W40J9SfjAA7mNSWyg7PW6u8z5l+ceOM3Z/
+2FiPmb1A/O5pWPi8yeqy6Wb5hbfb+Nw+XM2fSLnYbcQK+bLi/b0k14yPJwZEQbNKlXA3ZC/zxDb
w0HvZbZggJj3xktcnMelau5xKVtob55dG1Xt/Awlf5c2FGfGXxSZXc3oP38VwFqUP0JhZ6S5lDAa
UBKnck3QlB4JN+Io+Dy58pn+XSh9rMCSwLgXBAvS4VrEHjn0ubLwrjPwA9vBX61LzQP/+Y4huJS6
h5+DOGkCDN9TPzFcvm734iOnpuFsMWtgv5f554aWV8cb9iN8TuAUSm5vojGwqScoDo0YT2C3l5cN
sl2okCujg+pqHR0nGh4GJAgaYz1HuVPgog7dUbpw+Q8m5axZdpNccosybnUM8K1orrB2zPblQVrE
uQt+5PNx+hEZkjb7GLk0XcSu/s/yHU57xJqUxb/HZbrcQbYZ5BT6A7P41gS89aA/d1PzKUXmcJo+
Wpe5fFI5kX7cfttqe1az6JaMvppheknb14aDFomR4l7ygjSFUcOAYQ4z9dekNcYWofwS9hjO+SIM
ZgJr/OxYmdoODwHWt4+h9eUmHzJ43A2C3Io6SU3ujaiOZt0qYeLU/zpjeJdoyCQ9cTmvyeWhVajn
cdIN5rV/qfJrx2Cf9uWw+sSHoGoj96eln+cqhAj9X/FvYyVbeYUpGs3Y1mAV3JWf/oX2jJrwzgwM
VWZCAJbmzRClxgGaYLUw1M1DfzT6NphznG2aDv4N0AyXpf1G2PcoLlL12MpMg3XyBBV96MjThdU1
icVXjTbFWwMK6e49Nhxr43EDFlTSZeUWk+TvJbD9qfLRjaZKYXS1vNPh59jdBDU3VCCG0aqyDHVu
N/D5HL3BMHwlxu0cddQwDXrCNQPXevwEnOkgsIlnbXWebz9pi9c88RuY2HyDw6wao2gxBxjKrDXx
2671yqn0oVWWE0ezZPP8nlD645ilrjNS6TC1yhtoehwtS02/jPnkER1igvWpp/3TMCbsCBZIaj2m
1Z6+S/u8DUG72FTfD+yipXLhkMuZmmr8orIRJ6fDdWIGUZEs7f/jXIDYYSjrZASXFHx8w6umQToX
/x9RhXpKajVKZJmSFMJeJ8qlIrTYh1TOiAk9AmnhmSAP4sAZ6mwemOfuDj+MDs4obEF9peshwTSq
qxCJENCbpcc0IhBPWYpPcNwetPMPDaxLOj3MXhhFPMdBSc55WsxA3ETiCwkrQHjvNniBgTHtk0mw
27LrfMCgBpZc6tlQJdCQy8zV3Yg1RXAoplLf00Nh0U9j1IdPXLd6gUWi9kdLsBerf7ieZiXYnOim
nI6xwvYqVStTkPwkzshSLiyMNZqdD+mF7EPLwCI/aVCtjKBvSvFiaB6VsfU92ARxufpWIMPxoM7X
7aWQ2iAukZAyQrPAafdlK3c90/aSshohvSGzYSFNJiOQLomCjxRzPACH0zWdbAdYu+Gs874txeJk
/1cwZBe24G2ANP9bvsz9NF+TLlIsbKZ4Hg8tdMfHHt19xCIW9RuPHua1B7tVCEZTBMUV8eCAMc6j
uCfdTfh35tAF4RqiYBX+gQKiSLN27Bfn+PKPo2e15fpR2coOTtYZOnM/g4AMJAVFqIoMcvuV1JaF
OURV44hjb8ZIeGRKiGkXKPdoPY8FpVBeuk+MtkrDr6tpbct+soyDQ2vm02hE2FyOYo/L4DWFukvA
nSfAEIhxVbRkAgJJz9sLidWkA1YwUHAqccUqEaHu8e97dIaCq2WH2lTLnEj+bV1HmCnLoypdtWdF
PsOIn11SnrsMNSDDtRX7npTxRuxHk1YkzfPXY6ublBcf64+LbFpPnTmPBd+AZUwStf6OcVUf/twG
qVhw4+u7N9+mK/Lx/XPdKsXOsZS8jB2rDF1d0JRL5lPxUQiiovTL9j3LGwRxstZKm91Bauk21AfU
f869l4haMN+Hq11etmoBqpykx0BE2jezSJYcquzRKqhvGGoqaV4r0pN5aJz2uIJPZ9ywrD4Ablf1
VrQo82sVlbabtUDPnzPK9S76Yv4Aiyb1F2y4T5pMjk7iCXPJ8x2api4w71aQB84SXyQpvbOIqxV0
w/UuMFp/zwMfhpZQCkug09wP5wCcyNNn+c0CkzmoVfhUvHObSJ4/j4KHvHsrE7BM7XGr/WiGCMrO
+Exh7HkKarGjXSengmrAM/0xq6WWULOcJ1SpSomTLaz9QmMbFucz7ne8ysXuDHWSQKBLvg1B3zoq
W44DNoJmIuMfEvTqaTMza4amX0uSRlJDhBI5LStXsRLTSjkuO0/KWHT7G9UcvDW9VVqwUB+nQkLg
qTJsNtYxnmnqRHeGq+pxB7CYjzy0uSLtpupUYhXC6hFVmuYyDKQdqD3WmWwbBbP0qh70aLTn1VpP
EQsnUsf+LA3TPRTtO79c51HVA81cjQVyYOYnctQ5QA9UvLtzyVNbWcBqE7jVW+GirH3I7MgfW3js
DAXxc4a+5gNP7ZMI5pjo8f1cH+HIJzYcrV7vfhktkAcB/HvnsMq67MLAaxwc3eh7Er302zH357A0
FiZUyA81AkQ1WhDVH5FmW11CWTPVXApDWSHCAWdNnHU8ywDvi3/iTtEC9sOoXQOM0Q+yhFQ0z/rG
RQt6MALYvYFrPwfcT8CinCTTMzb5Hdpsyy7HpYCeOPKcDUBXjPgiFcgF5HabVNiqhi5AN4A7RjgE
ovKE+pgTFq6TGKaRs7Z/bXPCECkfUtFgwAM5gvP2f7wH0w7ghqB/5qSmQ4wZw5o9ZV9OukDQuK5k
3/BtIx/BOlJpdu5fvONz7ZH/hgn0X9s4QhvTOIa8DT3AJ22cs5O9aQADjHtFlXpSF24poW//rwbV
cAQ5onvczDuY6semxzBaIL9P/6ybu3+ThHrCwwVstJMBtF2kqs81AHNyP3KLNItT1zjZXu8oJwqR
GbacSmGWjXQ3SOQU2v2/k1DeG7DdMHbnTT7vnfly0tBJpjNbnLk13AKrccVL98E94PcLpyktHUoB
khGruxGu44PUQDHIhgEhJIP9S5/0f+hXdbgodcMNMKqplLSqSqWRqL9ycEvnA+3OID13L+y1hzgB
sIrpX6+kiPkAyEzI83jQMS5xdFfFi1Imkxdrl4ij2H90ZzKg4WSWVrdqN+qMZZYl7mUpemUPOq7h
gMuZ+3xSg5WcEbArRpHGLKNnRBYmzC4l5qqwEnxK0kmd5vCpbIKnPRdPJ9upobU9ibcZ/Ud9X5eb
JL+eXj8gVEOgf1cnUp8sppzxKH5Thk2h977vyQAQpKGv3zHPvA4aGC+5jEVD1UFwYXaO5f728c8/
ZPGTcU6GDWna5WiDUW0PtUv/z9eTbL8G6d5xJD+DMbR2UyMYCgIWT+Oif/NJ76ZP7je23k9qKOiD
5iseYW5xzWBnwoBjur5vD3MXFi+dny2eBsKFdqmz929v3JKwZ3YxTtWIDlEECOURmoLfZc2thbO6
sHT3vGMzr18xghwd+QEpn706pYB19anmAOZ/1r7hSzpH1Vz7oqRsTR2mQp/jcZcwUwpWnuPbmd8W
H2tNN+EAGD23khF0oBDkesX9dXtb4FdzUm3prpsOEs2jF9tp6jH0rzNLvIQNTvYh0Dv43YpLHD7d
5BRUJTrB2ezbIyND+zjUyeP/f76PpCIt7ftqH/Awhf6g26567hQXvalu6bIvcYt4HrBILsDHv/Pc
YPMn+ateqq6M4OKuWo98bfBoGp7brJ3ezKS1nLZ0EiWLxepJWDbHWy6Vbus73S9m5oeZZx8GZuI1
0z1ECaak5POb+FzCATNefk7kNujmBK1HxjEswZwzxwDZCpQ5yb7OXAEx37vciE4QLu+V5N4034Bn
2l3tO/Fx2Z42G4Bg2LD5Q+KOY0KGr5qQwYny7vbmS9Z+tv6OZA8qDY4GR4eFBXYWqoUsB2wztuXz
g5VXsziuwOzPDjl7INOQ7BJgrUFNhCOytT6Q6r2pafZvYhu5kSR1F/NZG+9PBYms4gBsegpjxpXo
DhvHjBJNKhWR5wqBPChwqt385WBgomms0xXXoUxkv1Fn5c4re9plp2UYM0+OCYtDCRa1TvqBJsiZ
GFPYkdjqk6Tdbb4Acaj+vgyh7Fdpfk3anSt0tGcW6TziED95nSIFX85/hS9/X4V/7PDcF28E1N29
5afPfDtUAR5Sc0YaN13NxYphRn/24s4iMxncIA88VMVuibQKnV21WU8/2ApyX1ATRa3UgzfYFaA9
SQmGMG32h+t1JgBi1V26EfnQOWMgQIHGUp9qkU1+uj4A4zLhAW3kt6fgjMgsyiI/xIV6Plsp343w
cmV5CeMfE5ADFXfzN8D826gc32sr8yUsAWn9Z2gBtqRNojmz3La8zXmxqNfvGKbnfcab7KHYE0y+
P7tN6B4OeDqgEREZ2/k7fR/oyebHuN2a92lo9cExM0HXT9KPNSHP0c0W0FdgT6LP0reqzJl0MV8E
PmoShBATH/tYUmEPsZgh6KOKJO+zFfXsZGCEAfWnrAYWn17fjrI9MshYKrvLTnxS2OJmScdpkmLQ
RIKGQDMvtsYCbhd5AqmrxnJ7y0YG/rfZbK47yUOKwG+L2O3T+EmfQcAm9mcoum5nvUsXR57Tx20M
T0ZmgJNyYkalfqUDWjB2Wpn6Vlg1UFvHNIzJoYZwDfdVDy+RSrTMLkz3mXodARUa+3dYEtOESiDq
CFBopEkKrEpYftDrqV8ZO5mGRdkt+m2BNT95RjnSAMgcUblZ4HmeZ8V4/To+SIBMVZfKejdrMjBm
4pKX6pEAWmcPYnX+/SB0gUct3Pz7Y03E8WvNusJbiEUtA7t72lzaHOdfWLlhlXPGF7WiGqQ+7EtC
cwAbVVgVy29Mpbi6Zw6xtXQMeL063nosd1cPHGr3ctr121PG5+uPBkZXNsGDkxx2nzpJBZ2qnIZj
uy5fAPTmO9cU3iHTd7k0izEU2lvFZGYd4ZBPTHRMWtY+ceT8JoNKcbP1tsRZqUFXh8jqqWZAT2Bl
kc7MO2sd7VBtiObvPm4UNDBD5WliD1uhTMQJAX7fbbBHSoKo8rcuM13dzGS87wSZo6OmZsMBy4vt
079D70VzHDYkMB7iX+rbRRHR9vAX3ZN9AQtWYmtMv/brE4cRibNMoYZXWH9jCQCk4u1x2xts6abg
QWH8rtZMF8qetn/dLSgpDh5EdnNd5QGrX/dPnVRwFFalfyev2vpnWq0x5xqZo3YxqnBiigOVa5nC
rYasLAZSrxKalK/0AuDvj2t/8hWrMrnZu6JBQDXJWpWzXCT+Ygr4WBTG/O1dYxf7SUhAgoEZWziR
5iXt34YCl5KNW+ljgNJFjLXTh9/LReGPKkxsXMqfaJMSdlk58ytw9EwngjKeaGPnTDWD9FZdCbTM
QNjs93Syzvj8paKZLaqtULYIsbIZBj974Uy2P52aqi6hgmIDD9ag20xA8QNfzqVm1JeY1qtFtjdd
/warg+J4JDwHN4lql05fTwHnz8H2a/2fYA1PUQ/dINmMh2FPB+vMjFTJ47FzTpI2FiEkdS1m3hC3
PCapPMYn+32L/vdJEihqpYOgsKGocKAWzW8O2amBWGVAnqiCK7UVEccjQ5wCYmwcJx24ayFD5eVC
esf7Vw5L1G49XZQQztQdvEDel+QeCinF66rBZaW/gYlTeHEcuP80mfiSQC6amfmGynXVBMTaFYzR
7BOMKr1V4MookByqNkH+27OvVCJCZW0cXAvTvclLPbr7q/jl6x4o6GxXyEzp42iel2zlzUcmXVwM
ysrbHwlNh2QB5YOUoP8Ia0RolOmql0Z//kV57gemlN+th3+U2zSdM4g3zIhvGc+Z/5ZbauK9YBZn
UMfWxkdmgtksgKOwkakEf3Xk2h/qWMUUWyVRn0iXI/zuVV+b+CnQ6XC4lV2upZWhUM9xhryiPhtr
3wtPJHcvwYHo68U/LxN/x3Erm8owPK7F+9RtbkpVkNIBiRygaRee54F6jC5p+GNGJzdRgCNkv4+4
gGdcq+yih6MdJ24bwT+fRIJ6Kszjz06hubW+qSbSQA1qZcBGO1tEI47Szv+bSKoWbI2ONYp0AtSX
0u3riwx6qVtR2sAQpE5MqGPMP+NtlBp94jt6Ub/MPbD6ymxldTrAiRmYjvFZkE2RIqRkbJVnKlHv
96gNnsVhf3ops7fp1HsnDLolGvLYcom4Wmzjra2ZxggeDgaPkPQo+r7QU7V5ZIcFJVGxqhe6wVMM
qp+4Z13u/S148kqhCTbDCw+33R2KiO+aogyl6NOgGVfVD5T84l1FTobRJDGzWYcAKjiyMyA4XpIS
5StK5Wau+BnN/+vgicW4Msl/I2VbGCTjLJ0PoF/KAmwzJxCA8U5yz4NT9/Bjz8NdguS/w96B/3Gn
/c9NC4kt2LFFZFkF7wzkd8nUTnDx4nTw8EZrRdzEUnX3HgRq5ZaoKPQaAXltnoabdG7ZNi5rBfH5
oOW7X8JlmYRcmYjvsIncT0kFF1wVeDVHdHUuSQVDYoRIz7OZYnhptA16txfnt9ZBsSNgO4lqBwpH
aHK/UIGULvF6l+HIdUP62RuEvOfooXHbt6LUipvnRT2PgGiTeBFx01hfecd0bY3HKtE3RsGaZFjM
1G0JLp7LkYpquQ6UU0p00b5hHdRW+V+ItCP2Vy0jpxGEsuDTAv3KckoMnNx2IMnjDRILpNspB+yr
4SBoSuyhCsQI3pDmaFyRpwNONk3EDuUbv8LXAEW/3EU/2D/1b/4pmadQHsVmofzOLRJlDeA+M0n+
U08oanJu8TU/EAbaB3emCefbrGwC+7dbQ3DhPWJUyah+NPZVdFF+/nontq24EySebrpJ+0dh6Wbj
FomVf+l+o1x8hPjbMxoLEup7f/HkSAd65JNsFX3zhzTLGe0YDgKolnNYD/NYY35fxOvegBXYyyoR
6uSRkdcUlaOKpvMSv9mhMefqeP8UqdlE1uzvdZbgvfYGXl4MkzinaPLilFzzowSPiTUnj5CZ8xZT
DsEY1y1D4DiDL8HpZ7dG5cPIhuPJWIaBVrgMuHMGyJXvJUiFWftbwKphlEYnxGqRjvXHXvF2uvCH
YVsJ4d+nX7ropcKSR2WJMwmEkjUIELAcJM/LQBytqNn7RVIq3ZWZnK4NtItdI4RiqkMztru7uNUO
Td0hxV1WjAgZm1uW1IyLZs7EhWayOy3URkdRgSJoatW/iKE66TWhRzoDdfFOmX0MzcKOpOP1cLRr
BHf/htYRkFf6+AqboU1TVdDLLYN8q25zpV8F72ojxWE3OamskfSZgPfzexFZ7vwWpHvITZbPysSu
6GKY/6UBBtcSVODZLMzgyns+a466OyD0KBxi1CarB0m3ZT82OtliCt40bwW7SWKxlPeOVh2YOoSL
1X7/sienn97CwkxAgHH5RaBf5aCIf7WOiYyiIn2HrRF5Dwov4dhZfm9CKr/JUk0s1Upn1WgkusFb
FymlUNUuKBlDqARPcEqHq22ij5Ekg9RxWMyiMDJD6pkWDR9a4Kav38OPMeI51M/wfm1LcwFQa3K/
fD16Bje8RtA9EHfXCg5GRGOirrRLlq4k4IpZqJuNSojkWYTtXhiYD3jAT0AFlTbIf8p3SphaAjBI
Kp7P/9M+J5F3PnjhIKt4lMLx+CuDZiCcqKNGsAnSVnYCA6OQnWDiqHdVDe+JY2S7EBv3sjHIkzSg
E/OLAzUHyti6u1OefjO9leVHLxmtcq5QiPNbitzi3Q8X7Pp36HWoMm0ie+jXTon0hLCR5ym5qr1m
wgGdS2unaLBr0P4wBJzmyWezCUSkUW0ZPvAfI0GtCEXkEKhfIF5LMrhk/kxXF76855mo9KkPYKEB
M5ihD5GBKwuZF6pD+28lIZnwlI4dli4043bRzKE39eV340m0wOR5dZ5+AfT/Eopn8huAtUHLCrTx
K24ok5hqhYQe+FwBBNvjFAnDBcQE2R6g7+Aww2O14sHz8yDvZPS8IsNzUM8VkL6fRO5vINS2LCIZ
qu1BzVcj1Eu+fr5WeSFtO2pGB3Vs1Dv5TdDEwOz60EZAxVz3OI9oCvRcL7uDxCoxH96LWeL+Vihi
XMwGoKX/t3ZVz64CHdRbNH5Hbjn/ddjMnR7NMXaA5HvuUCVv9BW2k8hv35Q8XNVDc0pDtydS79vM
iTDyKidp8Ggb2zISg22PrkjeXdol7iCpnU8aUBkDDyj+v4g1dQFvon4CXu079xXlfBMg+A2r54yb
+Ji2YpZSqAImJ+vct3wXFL+7eKRoLTbhZysebz/Z+jIedgsux5j+W5jdtH2j271Ds8WldshyNGSr
UoX13crq/MM554v2CQYJH4m4f1PVX7miKGLWs7psh+my59TXFzcEX9ZAgQoB/hJl05Bf77A5Sw1h
1UwZV0JzrRvjx4mOGseDdDttb7cUuUjYeZsuEcYu0ngj2NtfXagsSdZKcwzTZrUrpbBAaOmjkqyD
c5DRfzsZ0DT//rWpdHFpZPwnowFJaVrnYyKN1s4cIyZ8fITKN0N4D2XIPNa4K5nh06qdaL3XLpCJ
FRgUqfjkhuAeXt7o/JvQdNY1lnFJanV8xTswIenNBtrnzx3uu7ntswA/0PFF/24Iak5IpkBkZq6h
OKfs2zdti9PO8TNUsnynMpuIP5xpcTpSE+PbIv8EQQ1xgUuSIsZISkSNPry1Cz4vW7e36xzoO7+/
hZGVfQvArDjr/Us7IBNbtt/T0IVl2Pad2ERAy+eIurgp2RTearF92Nl3jisL9vWXQWwJEpBx/Uzq
R4AZLjQ4QTLELLYypGZEAZY09JUz1cGA4Um2eFSmn385Czaq0no24yT/fxaaXt2+T81wweNjKI8q
QDq/OE35EL6NWWR4vtV1jwaU/6mhGjc3NlBA6qwqXsDh253DZcNSEwkp2yOYaUwvgjhFy7Ci09yd
A6QDK0Vvapm/9SyDoYvC2T8CElOU7YZWmWcezyjYaSzENWdeZ5WkOlTNa91TMH/5Nj5oaYVDLHgG
A9ITvjiRl0BN7mhJR2mVmchZpRgIyfz4Qshj/rGN5knlXdAC8nyh0aB453bFgd600n8mErnsnpG4
+qk/R+UqrfUZmSPbYCygqINdOU322Gc4cSYqIQkdqYXDGfag5fE+2KjL+ThJJ7veHmHN4GZcqV2A
oegqoZ72zmT1qyFHkRKWGX3NDi0ZFPvfLxj/D4IO8xDnkxq7gwWHkTWZIH5oqdo5xxz1Deh00Csc
DXqem2ph15KQF1YRRFo0yke2rllINTyPRFqzS05QpDiFoRaGmIKLnvvWRJdVV3Qd6nHnwhX56IEu
Y0gdNn1snDzIHR/1p4kw9hNHoX87r/T2/TTizmz2DfIPuct3tulSgOsKNfnEo3cmBqiCyU77kHBu
lOUiCGL5Q9Hd6w9NGJ33XHmBMl0wFMeE2dPMxXyHcBzyETyLlUxNpOdfWGv/GOHlKpRvmZ6AOYWn
hdeTGABb0rUW2DVhtHA85Ci247vH+BMUgKEhsAHUn/s0L7YJE2YbO4dt3oRx2bi7PHnbFAo5ScWz
EPBSTjlZ3fZY6bMtC8ZyVAAJgG4XDcnLqHyaXSR85+IFPd15i43GTI2guwBwvBPZ5Uj+jEvcd5Bi
h01vYjMXfIe6U4dfgAYbeyc65GDCOjsCnCnbEQU21k29foKaPlOiYYpqV8i7axqQI32e7k4tAJIG
926/SXtKZ9NqOyyLtw7X4D2D/9vt9BgxIZEhVYtkmaPmeiDm/ioK5xZYSVbZLkzHSjBN72Skwi3I
noGKr9XDgHcSxq/o+uRfBRTHdk1rTBqWJdSau6YbX7XJxI6O2jhaYbi99UOzwHq2zsbWrFLKDEA0
ZLcKybjFwc8hid2aVDtJZjk6unUWgi1hQadiCKRUJJUZqf/qqtW6764JOuLtjxnjqDTcFaKpPQBH
+3yZkjxAHdQq6+m93DZd0yqA++ExT9VCCmdyrhgWtVoQ3y++6USNmXpVgwNXSHSCG4LURDd13OB2
tLI4+e6Oyrg8XmTaswUXXQRMpPDkZfptyu0IjeufMUoPBGWTctNw748oemMDwpPnS6/ECGkRWnnU
rz+9wIaNToWD23kFiRsc3xdg4sRNRJFh6D0uA6f3BiuN5v+OdCh5orN13y+ibqoaBjMbtbvuYZf4
ZEx/Nw88AH4Nw7BRq8RIErWO+KikADL+ioUs6VjKJJ1frw7NoPRN9az1xragEFLlVpDYPkNICl6R
B2PFbocMhNcXTwDZ/WO9p5bU1+frp7Yun2fKY8KvNqnqpGtSd7ZDy3WRrZ3KLnKlFReWvjOWwxui
SfXNpk/epmKZigD79Q8h+MbZbXgOdjcm387/Edm3JjehShnjAE+kCL1AxJydoYFc9qu6Lb5PNTmG
vsl/SdbNWviHVZB4xW2WDv8wSf5VIWFdD0xI8bfEYjS2tgjscMskEseHELH9xRGEwrDbUSnk0uav
HRVYV+uSW3hhCrNZnhpfywBlo/q/vP4OTDbrxJ2Qh4DSd3wlelVHQ+yaj/qYObwDOMTmTfROJFd4
PdyJpGGleu3qjcUgSPQzdIpvpacszmCWqW5CqSF66o8FMjfh8gAiQqlJ8BCe39a3F0g4tG5accYF
noP7857rXaVfhHEVexzDaoQ50hHUNdmJ7mZ3/Asp5u/N+OrOj5MQFMWmBTO4pYULee7Niq+uL93C
gmKrig1sBlRU0lmNU8Z5N0H0piOjfYbgAJQ1uDtJKOEl8e+p8+vvrSzxrEJUON7xhORs8LXF+Luk
Um8aIbKDgbzEDmVAcQQTUegm/BPANQ51qeEnGey+EbPFKyx3dhS1iEDwhnHiQj/NaQt5Tb+a1QX+
Lu10icYTID+kA1Ds87YSPLYgy3ifTm6DXxxdeS2RdcXNuXNapcg3dRabsQS5O2Mi2no6FCWKWYMY
MnVubcUntyGVKsF9VXfDIrK3I+OeZGZDV1ExBOakyyeUVLEpBeXEuXulR7Ttiu5NNzT5R0R9NqbE
k4AwB6OLYY+Bio5ZIeg9bqkDb2tYDqm3s+czc1SXezB6QV+QSh4sE/aDA/vZAwzx112CBNVovbV/
eF8PKEiP24UnshZW/OFv1uMLc3vQuwsMljCRxDtKURKxHdFmppWd6oIBYZ1RBsSmcPEEqf61Wc8E
me4q3JaguDchrXn+oWYDuLjfdkyn7/l9MiMJV9EQL7QunCr8Zu/Zw+cbdlmKPTC1iID0gvKhFVc0
ejcBVmP0QST0F+L6GvvNBXESqteSrdcX2GyKWTtZnb3IlvR7vv7s3feLiPIAMZF6v3ClgB1jpJlf
lJWCJOHNVUmtoITBszXdWdw9LP6M0WupZ8UImevM2Gpnzx9BVfyndy0hBWJu/rrBYHtpW+/THjPh
5MZxy47uI4L/dci/lwv5mIQhBuIx9jtdLKElg5xGXc5McWYNASmsrkBwdgn2LPah5WOJcwmypNUE
HGiawY9niLRWhNb2+o6Vrg7g+qmrieH8LFRanMPJVhT6XdnTisBvuaguzKuOIZ+zjU94DG6q2UbP
m+/HTaV4AboCjqB8itQ6Knag73LbUbUnpdHV0Dl+31hdSI520pRmOjKRZW0+kbS/eBm43Dt2DSoB
ygXMTloR0M5CzIDLehs8j8exNCViZ4cv34XSreuaJ1gWWjSQ4pIy/CZhEuQ6ibdglz2IzdUpRTWt
8xduX4wpWGgVvR9luLMFk9Ssv7O+BT/1WvaAMqq5VI/o7qHlDb678ifU9SmiTGTkexSBrjlu7pH1
mgvPfXHEO5z6CVOBHNxu9bNL9RL/r+EyXH0xAXvRQfYDGR2CKrkz/BvdYZ9bHCQIA35Tmsgz/zxo
QiLnBtXTy6Y7I+FziHS/t2AL60rWyNOaCMz3vtI7FO9kWBkUpsl3r5PTq/AIPI41WSJGosLnQcFb
x+tP/k9E8lQ+fLsNityfk3zReDAydjnJBAOwmG6wQ0nC9YTgcnl/iPhaIG5eKaglsf1ieSNr1Ou/
f7EB5mSW4cXNvV9q42ZPZlt0duoGPsVb7dO5bPxnhkf9Rbnb2SlMHlH3FJup5tIleDAEEVHAmQYS
IpRNI14fwHRCbRHkiIfqIzkzaIcCtaZFg/3mAgI9gq0qT8MtqPXSWdq0QG0dNTZsvjUwuY1LpIaf
xh78Ql/BuXmQKaqlV0zuInXA1CWyI86i86M7011MG0HiDcmVGgx8fzdkQ+jGZoFeuw/EEu1WFKAO
7DpF8kruOmnast0ljr4Ei0L/wlZLXukfH3ZSIKJ+Vy6z7rna8tIM+HOxpd2+TRySfz2NIgQssz8G
JQ8O3z9sH7YIauPW6j+EZuuusnA9B0XDRfSBT2ei8E6yOrb+CHiwF9ckrApwZEFk1IEbYEVbv+Y1
J6kcpfdDS6K7aVsBhErDGZJ/p/Emum67Gf2PvnJ1dIRT/pE8UjXoxF9GSZ2kFANgyHLQ0mfir/R+
2k4Vicn5Tt/0YLvUGcoYUPPuzKDC2Vw3IaqLHiHC2gzdXgvMVRCJ8CuitueBjgHfiY4Xod9xJ37h
v1CwLgZTVoHsAlrVOrxJ88rs5xwIM7xomKAPM6uxbatMPnDdg5QjEH2zegt2w+GplasZp2Z4gvoI
rrvlo3qiytElabCPGoCiMCt/5QljOoeehcUP1SRvMGf6eiN8ELMNc2U7gsDSdpN63CXQn1uMmZnL
BKnrn0U7YnbB0RvX7T2V92NqFj/KoaQuQtQxxfLfaE5ZzWTs5qhgdepu+/yI48Kxoz4ll/MB23vV
1T3gf6DagpwljMrdbeJ3QbJVwTDTk7HcKDXWotzpJi68FxdAkuOTawrD7KLlfh9AUCR0ymyogLdy
H6yzPgCSdfh2nG8RtuXDm/1qZENa3Hybf421lcpnEszn6UWFdxsmNYtMhT1Tr+h5KFuCstRkEKLJ
mY6dzr5M/SFLKDuh1aLrrAS/KuC6FFpbDyd6K8YXnKPOyEBqQYdAQggMKGVA3NDc1pg3qUqyD0PE
sCTFaCgfvsYMmZrfa/QYDqy2nl4FX8KCe8MSDgAEOxowVBnId3+9HILAW2ykBkUlA6NCCROMeNzt
bRPE86qyQjN9wc6NU1S4O03evYBGYAbQo4SqnPPIyJqDOKN1AQygmh1cXVRyd5OTNTxoDkZU8/co
gN5LmZ6uh4RkuPJnli+48x5I7gw9oXrcOEVhvNHGYnZzmBlo0+bbEWVeVURyMFv/vEvkgIxs1vRB
Z9duLvA//oDk31jZOmW2GFJKtvwI+aEHYlLhAODCc7NLKaDfr+VMOuVkgOcanSvhVdR9nwLBqx+b
p3QpMMGl2I4y0PzR/6WpdsXLyiXTkx+Cq5nc0rQ1Yey53nVDaS9IqMOB5PI3P1nbvL6gnK8PRnAu
5YBR9q3HFvf1WvxYAOXbMHbOz3pwInXzkVIPI612rHDkdgFOKXorYltuoL31Lmugg2oxHdVkPrAV
N1YWFEmcQKiZiWsBpKsbgG//Bxr3M6KN0gVV6IiO5GRXo2LR3ReQutQTfgteHqCqo771+jBut09e
m5Zxu6Xw9k5LYjjPLqfRUp/Mq5640eDl6CVDHfj5BDBJ7iJ7Ga6RLPn2+V9VS8WxYAJT2y1lJ2B7
qfkfDBxA4TtxLZlZpJ3y691KFfq/VjoDlruThpXRd2hf7e0fyFq2C9rYS/XTTZzr4DmqvbmcPRVf
n4iCVe/Yf+TQKTnY68msjVP8PVeavaPUivmNL3dYnRMuHGG9wyOfnVwbuQ+KVcAhqDVhvqE+6DT8
+9QV1ziNv7K+ViYn7WIniHI0gxVkNvb251tGPcbiumn3yq3E2fRgVCYLdqUOxV2WzD6GRRVTuNcA
AL8X9lKD2+yoqn2BArAN6sNvee9dWVbUBPC9MIH+1ps57FywLcijXQj99BvjyCCO7phJ9/qVyScw
2k8ZpBJI7wlJkuVsu/bXdARwC59V6Hv6Lrrh1r/iF4jIdKmHvSw0OSY7481DFrQlEmgW9gCWvAnj
alk+dC4zxlA1/apH2ty8MZhP0IOqNeD0LCdWkaCjqb+dwpwTmDXqrIfotTMXmNhggSU8CZV3VZ3R
iOWRgksDNgrmGrl5mkDXuUSruKLl6sFeuKJI8/+0tkag7JPE1CLSygACJvNrDkUqQlE8DLpxTKz6
nhE+No5iWjarlGUfartbcWM2Cl/cItTWJhFxgIcA6OzMatp9Y69oS61aL9QntBLGDI+ith7CXVMA
ah/UgWYjHlx6aKy9apLCclEZkQUBYupe5ovZwCH+8IEMJEBp44TnxWCq77CTDqyfmSCCokJ8owbL
gXhTvrxoQeDsV4HwEh/AUwNKk6NlsNqdSP8wBgJtR24pTLVqRxzo0ErH5tkFNv2AXxPNpvuSoFpo
kqZNWCaxLr4vWwgb0H21JTMnawLnrGqsnmCjNnnBpgJuCwlshT7uDl4fDkFofOqqTAAYdFg2HYd+
CoF7ZRVugNlB/UBv/X4kmFpE8MBxvU5di5+5ZjAsw7glPa8BNUFafgDQ0MaBPjSMGQjggdQfEmmQ
Hyrn5yTp6OMELEW82P1MTsS8PhpSISvgHvJXo/l7xA6gJRplt7ue8V9UZXOvzxgDuiZ3UnhzSjZ7
iLSL76142XNcZjyM3zmgNh9xMc7UNIAD+tH3yfcEmDl85xkS9VnILZHzSpzft/Yiay4vaMOUmVMr
RckY2aimR5EcyWqeFhqSRBsFTJYnpwvzbOH8TJJdN9QLgPF0GFZpbQMSlcSEGA28EjBsbgMH0wwP
SRPfWWZJfwqnoH+7ZQU0ITglCDRI1i8xRP3o0CmMJEKCc8m0ijyqDRg26GFFiCZBh3VlLaz5UgWm
G96mkDZQbEM0G5RAYvWECdPqGCRH0IKsK6WNaa5IcsRtKmxsdbaeKQ+gksChczkxzfC6RGdhkoHN
UmrdyckiNg7uoU7D+IiSaEE3fx2S7YAAFdkk1jOq+GB14+nkG4RcjjDhO01htztveqhnV3ypWnwn
e/bbnCbxchi/KfioYUqdTVOJTpxjYWq2lREVE0o2yndrZh0olms4sHPnW/g4StdsNve8SPEGlkSN
zX5VJ+cbKevx+nD6tpeLRvuriQUyN5cbOlTKV0UIhuMpH6X6BYpuU3pZhJa/dSQQlu9PMm2GqjYU
Kq5+R/PTxMwf00NlFklAPEUeC1STYNII7/V2wS56r9b5qXTDZG8uPwG4UMt/qp77CvgRKJ+rLaJ5
EDKhc6AxolNyWbSTNbHYMXqFzmJ5qdZ5ZZ5xxjkFgyQnhGFYFYJCicmzRLiFmvNw9QMrkkKZC7St
l4gtwSOQSc9fgokRfcCUTxk2h4fb+g5DSv8RzqDB6RhmCJEMDvl3QnV2AMpWQyYD/9EId82wrE4K
1OUHPy/6A8sPjgONjTvuVs+C3SYRIBN9x2o0iiX9PR0lXIaF7Ehb1ALzeBNus5enKrXs8g7lkjbF
vPqpJpbK3MDC5OC1avKU8qMvF7tMDEAtPGuYZIV1hrQcYUgeOl0S9YAjp/QSxhnvF94uNidfbMmI
zhtal3EoGay/qkb26Y6Z9uGieXNcPqD/wVaUtmwZo87RvxNoCE7CeSN8ltJ9NSzI6rupREqthj3K
st1FOmIUMHuLsDB06T0v+MKPb4OZz3MDzGhpjymhJfYcBvqQw93GoTkXxfYMi9cRbx8lJ+a683mh
TolNSR9YkzFKvMyp21CujX91QL0KBWNhFGss5qEV2fGc76ak9ytz7xwEuh0yY7IScw90kwi3QQiv
vbJbMU6wCYxJiJ+BEk5e/cK4yVGAYAzdTWiCevuuqsgBHVw5gYxeasMhMwD2Ln97YyOKeAKko6c0
74uiIV+QpNvcbcpcL0M58wBKpOjOz2LbCJgSzT2aI8erPfG9qbRPKJmzvgRl9w51GJGVgvKXQVz+
bWmdxZiO0ssF/477JF7BiSvOwzAug17VSUZgHZE8dP9D7df5lecYnsjBz+Aw8OsG8z9xAB7IOjWa
EsV+nAvKGvJWX15kTU1LHQ9qrC/CVLMwI2+N/VtV2fhmxjR3w33/G9UrSzuN/92NQtk1qKkrV2va
+VtOlpjygWhvVcV32xdNbcSfRRmZXr5Bacr0fDzWn6l06wz51bMAnfPDdARpmgnF8sslqcH9jb9p
PIMrrRRM41vtjsyWVPuhjb46+1dC1ED7tzrK+qpA1q/xDB5k347YHllwKLlBW3VT7p4g99ntUWGB
XlL/xS9oG5tamENF09ZZwsv1r4wtcoNuScuFw04QSCBS9iWhJQJzlmxRA2APIq6p1Ldb0BB/OGyD
5V/8KgGwPb6drP1T5fXTtYDc7AaqkMsxMDYxIv1aRWzHqESjPLxsCGPcCHt2EWIIpMa0FkpKPOJm
y/3sg7oxebZzDjPq9X0rs64eLHmhvFfv3YDvw+z6c31wFPFdKOVADoP8GXetxK0f5RaZ1fySX9nL
/3ArikB7x6peRhVcZNK64SkoWfJ1/VcCsq/YqW6fOPf0eueGeY7tcoqn1TUKo2GokfkWPk+cVoS/
5KfqJSHVckdf7UJOx5/MUc4Aatprwzj+f4eSTDrma6ZSxmCfBi1BGkXzkecPCfFXiYftKYvF9vmN
+zvlU8ml/xkX807gmEpHBWaxVE/MaDjw5yUiRT1koDlX0azkGEsjqVOsWa/hR6IiIVHDNiPywfjq
G7mGNsC9oi5VvQUBiLhyajX/jvrdCmnNLrxFmoxAEsj1IrNgx1n5kUfHuEZu8iR6E4sUnFFPhl4F
gsiJ14I53pE2aunbtCgHUtKTPMuzKfUqSRN7Om2gE/XXnKpr7XURlVeZZud05rgLbK/z1Ggg4Qa1
xd6GC7yDTL2bKbKkGwrxVFZQ/N8qQfMCxp79J6a6SnwAIO+NLK1af0QqwpZHFr4E5Lp0GX0/pXSS
jcv3+bqsNTTPnNMmRt8T/y72mxnVeZVOeGlPvSRT5QkCTjm4Kl6YK+1yTpM1LuhFonpMD16qtKeU
0GNFw0hzHmucf+thHEDHsWRbn11Vnw0LNnx4zZYICIT+hZ0P+WkWUo8I3tzC3Fln/pZutwUUPD1P
olrWP6CW0sJt3O/cFVcSZWHT5JPShb9IgHTaiorGau3t1QUV19m93p4cF5y3GiwfDqJFQdCm5bij
VyacE76CkzJAwyKwVln899dfeMHLoVsF7WVkLFKpWKkPmZZ4xQMCaUtvxoBS/BEsjPGa6KEDL6cU
Oi33UHWcYEYMXBTvL/J5E+Y0YTBwtQoZsLEhyUpJJWAsdDbrI4p8LxN2q19mhgs3zFrFFXw2svC+
nQcpRT3CtDXpBOUhjKvlfYc4pZpUq7LlxHG7LnSClLC86QXgm8HaN2CAvsxK4vngmJ7uT1fCnVqp
Z1PDm6WTjwMgN8P1RxltLkz2wZpQ4OpL0FGLRZMHQALTaKEGbIMrB4FiXBcKXe/VMOQDO6S8VQkL
zC3oxv8rjx3PuKGvj8ABYgWbULcazsnqmVCaZC9+fxkPxFzO7cliW6neRRnwG3B/nSGIkERInOJZ
1vKd0VZZF9B9kA+abA5TQ9ZU/lbJuVCSg0pdNYqVb04UJNOhWQirmKvBTRPQhdCMx2YdZMSrxmmx
OWN7nfBnQf4+eeNWWd8d0CXXKoCpwMFXkfPgJZFW/uAxK7shO9M3Z6QzXCePbX66BBSITWJ3o6wL
yX1wWEBhqpYRFj556nuFyFInMcn8HZ1kQYN+NRNocMzgsfMQ8sSd1yd/Q6lc+mRONgvNagYhWZjJ
4qt+tLiDfUxfaJrOPPfE1zg6ttOCQ79BttmsGTRnlXWryGaW7w/chfLRGqGmT1WaBgEsyfDKCY/d
ji72kq+KayCua7ooZ8Rb8Pvt26YgTldZCjB5CxGPt3QVplSQ/t5xarKtnCr67QnMzhBocvdUAUhQ
gMblP3VABQpUzOP+2O3qw6nPI7YBDjGeuEfZEczI0eeki/GhytCg3bHpaiqbx29hsA2iBScjg/sO
rB4nxJJ17egR8Bjrj+0V/z9XNSSRlnF+CxD7GNxprbwDNQiWw79pTeugNaCpfTy3Y9tAW1hGDV7l
AlmW1pcTk9jvwFiAzpdu6SpiStpBG4KYeEtXf3cAhNeUIeMJoKzLV/vsHuFUUB0Y8vBWnhhltpl4
wz+glaVE3tiP1AsDh168cnUS9pJWok+gbssDFhH+m+wUPJKU4DJfECVNS3qqiGQetNMFruJyC5Sd
0gBGDhbE1Iqx+kqMDL8Wa+pIsVU9UK9iQyLaaNJkOD9kW2Xod1dC4Zen0duuaPZRU3flmlwhtkEU
mRHQIl7EbbrEyQsN/evhjdIsR6h76DdmmkAZd1M7oqNFDm7Yog6Vp0uSZFiaf833VBYbAruLEPDb
Ypo2GCAfEdSrpvdugdG4CkvYO/MBC1IMkd4ocUgQTp+Z05sClBHLAUstkWTJrQtxjMhxME5zZx6v
NjC8DnMjOmWObZ23qiEjQnnLpvhGLfFg+9sqqR/W42uwZqcM3gl3eJG2QEfdMzZHXasYYCZEnAhj
L8fToz53sQB4SM8lrW2sZxf+5Uvs/895SuD4oz0I6Ky9yfQIkJ5Y03bA9t+3S8U33ImyWkxN8alR
x0ukp17oAGPoCnSasVvTBMeza20DUAYotypaCiqF3ffooyZQg/gFoiwv9b+ApQyWAkIdSDD6iUfL
RPsxlD5Rgyg/Y4lu/+O29TaCZ1RKTgTb7PYhFlSsDj8eHb4StzR08rBrMx6+wmAF/C9FM+kobWsu
pP6DV6gSyu6RpZvt6glEii42pavI8kGtZ60INia1ohCGvNfzReMb77VbEci4ZW1fDevuaMy3jt9O
3m6NiC8o5HqLA5HBa54fOiqsnZXsFb64dsPIeMrR+B5dqvlQ24Y0Ta8hOkiq9oPAuiZqHdiJJS+0
NXJT3BIuH+YQ4l6QE7PjMKX028/jQohbfSVqQV4tnxPq3IRKnbuv8tmGr+62hb6giEy/kvzKQCgX
+APUjksMvNPWOBks5gFNlcmSdHbvxyFOHlcsA0v+mtzsEg0xijp/vZbxodgZ6ab6vr5nvahT/FGt
1uWPqL+AFXK4HAiy7NfI1HJEvmsbSbFjEq7gMAEGOG7B08R1KNkeREqoAIDO2D8FEmC0cnuoevwM
L4Zx2/EIbyDFyfHK5PXbGdKRhTiVk8dN3hMI5T35xjbJQDcy1zfd9TjhtfiIeSGwqsr58IIoNPTD
8IKIQX4tBQ05I44N9W1jZI1SC5kv0A9HsWEzXrSl1v8gnZOfbvn9xkZMcLutMHIIfsvpqMNDmc4+
OP1/tZksAFGLvoRKNKW7toBY7IE6C14xNjP6guw65IL0QhrKwnnpYPTNumlW6CoVJRmelxJeQuxY
2fZ5/GnsenX783TCnkPhnM9Q6veVRyEX+J+nH2Hluaewx9HAG89UWermi6KpDMrqkz9IWTe5EjWU
HbgoaMkE76+DlrBoPxPxWunvuRN+1xyriGA3cm9qEUrwxR0rzF1SyQ1gmqdbiCDN6rrV0UFaDC1/
5DJXf6YgJetLMfklMLecMvIOvWFeiNZss1Z2adZztjtSn4baVleWDIwYHlBBAK+l9FF2HozY7pQ9
PC7B01HRInMkcNqEe9PsjLxTOpnadQybNCR9EnR1AbZKl8NU+hU6c/hEj0zSD3gLAGb6kt/hKiKC
/ccXj+dKveui7h6U0MGKC350WycEibJqJrpuAY1ysNwzHav0oAvPMJF4zII5gBj3S52magpzZGRu
Rlom/kb0NGzDTpdWLeuD6gKJ9DiwYn+LBrqb4q8ZzMxhCH7vhK5zPZuf+o8I6E7xxsKwUNllWM4R
Qm9BmMExYk0fsaDsp6JUJu9vjrnqaNORnY8wEEVBhBWqbq+aUHeNehDP7uZSxumUmyI+QT9mHtPV
UL57MHN90sFWNV36A5yKUL1BrGct04RS9DBcjjo+nMdrEhE+25WhABQ1JdUNphzr32OItCzk3El5
ty3QBq6VZRU7oQ/LqR0bgTUZCdPA2x626HRiLfh+BQpo5fzLUJNAMdOgJA2uwo0gA2gz7+PKlIxv
lIEX7n9JrA3XjtnzsYoaw1HbHNRYT914C6INfwWYoJo2110W/sRCsKurz3kyH/eEs85PzwZyvJNA
3ixt2O93Q+ga09yo/ZZMgwlZJz22U3qX7SCVrYLOtFGZMHdpGv+wxbRvvtzLGkrl0G8NKc4IyFph
uXcIvAl1x5Gi9PYFoafa/oX/SAP8PxZ1lfsg0SYq133AaQh4KQ+u+HvFeKE8o3v8iW/X+LGuglID
AciDEszlKIhy8/EBzH+tiC68+TRBXtxIdsSR136picdhwBjyRvqn2CkXbpHQklYcYUxie3fviUZR
Xj6ko6hPKg55DyM8BvagKa3OewTjZJj8+ML4iWD7EQO8o2UGkyIwL/axdbkggbdxNIBuPqF3TNhe
hgof8wg/niw/ZNxboj2WlawpUgdNA/KWmexFaM/SrOJSQN9ypjREIEtJisNvubz/DDfdfGSwk7uE
uzPx0/qZlOtcxqHijVyyOBQVcYKFrTN6OEjNbiWLp5ukP5qDI7EA8qSzJWrHqTxXq44jrAntMcp0
TXS5mZyWgitxlqHgzAgYsJs9UqRv1QqyzpHtaxa+KB4qv4FXMI9dyFYlk5ygXXsq2B1ZXYqxc9Uc
aeoP32aiQEOLo13gnuwJ7DenDpqRAVNzlMr0UVt0NKLujNGdBvGsXIpDW9utQioS6m7NUWA/LMZr
I8g2kEv0u83IRSaVM8hQHWNwB3F0Evd2egQhnRS82dwHzRi/+jeNo1c5abHSKFTFEsARgv8833F7
CMG80ohXey2GlF3ax9/pRtD7wxX/R0xHQSxqaGUf6XzY4krL7GQRg2uS9+KTF0lzuGN1WDMN5h6e
S3vb0quXf4nyH0gJVuXyHg56fnrSd1oV7ltgqkQkE1G2gx/5PJHvdfpw/MKoomEfssJU6bftSFy8
CwERrFhGRKwKcuM+nkCMCexdfhL/0HoJ1+fYWiHbYgVWJRyaAv6R3JZimdvgLNSEgIZtWfI8up3t
AyXINm9tHuSoQG/qEPl7acgTqpeobdUK27UNuXyygvkIkjkkXACYtZdKObEoAKbxn7T7Gmr7947X
m8/q7LNiZaA6iSnpHnOzTaMIu3/rwhc1EkhgWiEBNwUjDpBc/84gnZpb/FSPtFCh9l1DlFbnwACg
SZb24EUxw6Ro1vlc1XryDl0b1KpZ8x6q0fXG3VLs82w2SNunq0qquGg+bwBg1yzugUdSxxVlB9c5
rQHsqXxF3oBfsP57eKXumDduj0JcsRRFVgHqzqfKyhoiw4X74eEsd0ie3yemx02bANyPyu+ypJLj
C67FttUo3j1lm85RNzc5BHQ4esvcRLS/66icLtz5JBc2osrK8kRZmQnDXkXO+dk6MMesZ5/6b5CE
6RKjg7WbtpPp4MdJeGJELHoDjwAqMIRfuM4W/HKnWF17ec4A6rzOL5RDjJxtFk0zQlvs4mklyd3Q
zRIVnW3atFawhx5SX3yDzXcv82OEiWp9On2KlQMpAdlGa/iBDzaYW4V3pa1Xpa4N/5reiHcsUead
J3IQ4ntOD4c4U+Ds6RkdGiijGLc7lNonk1tV8SRtQna/61qRHx/3h32nZ0uctM7Y94VuQx3qVVd5
8PnwZNgO7YmwxQCY8tScYryLLumObN4HvVq+BW5yRf+3E/D64Z199XL5KIQTbcoRKhj2xmHzqxhE
AcEulrpZVu3//GWXYfbL3TD30VD9xj8oUCo1P+unwMTvCTPv4nJz5IEtDsWmmUC5oIWcqd3ahTsk
KDYSY7zxgbhr4JKiO5gSqsnjKNdnOo4v2K/D4b5Z5yeeLsrtmY5rKTTBQkAt2vscuNR8AicHNiQ1
WONqUHGb6m2aAS/9zRxXHcTfDZ6hAU1nSI434fbZfcBnH7YR4ONPFwfCZrE9lA0xmWMyach5YMgm
jr6z58JX5NYsVeo+ySArSVINsD8VL9rjcpx4KvTTSqR3ZoX8YEqQpfhbmbrVBIpO+6Uu2SWbQk/t
U5uZDMC4V+qQGHaq1uOIkH1TJ1NkhHF6f39vFaUbVncO126nzLf7kD8YUFEJkwKuUH8lrhZKQu18
XhRPMkXRPaygrLXAVg2dhRnO36RqL1Jc+KwPNSZcqm/SXPWmc4csoJhKI/dKhX04MJKccZptJAec
Amx8gB2E52JlZjGBZg1vdx1SKoq95jHiqu1Qv4XnmYz2cHQV+oOfaOtEZyS6E5WP8o9HsRxTfhLh
S23VaIsTudEAVai53vrHPasqBIIO/JSpGdJ4IzEX+GY4vfyBi/7BAjRuPoQDCCkH+7Sb9A/GovsC
bF6DiIk7AX8gRlrjr+xTQcYyIpQkhJkznZYqqoLMuWDF6DZ0DhUaqh4ga8BhR6wz5dInptJxEQhf
Qa3OJxuFhap3kw4DMyBqy28AXANQSt5n1dcAjpZIHStWCZJ0Gl9z6JMW+HvjTYC9iAlUADBupdcl
dfHU+c5/44kWQMdXeqaJ86HHBfBly2mJn2jjFfB76m59dIkbCRS+iJZazvchkmaLIn00m46B4n7B
pWM9ABO4E8InvltYoBa38rpS4CopRLk7vC5kCnGFv0uaZLfv1ajKJM8xoeSgDn5TOb1h0EvFCz5h
62PfzRBRsV77ocXdqjCKqOck+6L+29WXXFUnzEJz3Yk24fpMWtiKo8RVS9I7Ys/hEHQyB4BAUoIQ
BQ0QhutXbyr6/MhbbjyUqXfazyOKdrrlanIzMkQ0kfEcqEa8F4ULfsDdX9yRmeIKG4Qhzp1F+G/r
toah03PVzYyly5aV3Y+/KfZDWUOipXkL7sX5ThmcRpy7j2xUVLWFXmTBCw/Gj74r48fo1eFXv+qm
iBw4REaj8RTgHlVszjfZ0hlu2jOmQJJJ3wFqmZ+EYumcvB1F2x5Mkq1QTMos2C3mfSsViWJkAxfd
wT/jrC/WomPsroGvqCzfaL2wAni8LCM9HYJFLzHo5RrSQvKnVBoX37KXsXSi6W6yQyYlx5se26BQ
QdcAekyJ/gbbHUUzGt2Kfe5CmH2H420PHNA7iYxGHPbs5axPXbj2GtBJs+9Z8xo9TRfitVyNxMb6
hOKctEDXZqFPnRH/D1JFAdIRfjh0u3Z7lEhDNrmgl+FGOpMtr5TtqUMTgO1XJ9Up+RyjDm7x1l7X
5oW+Oaeyu+R3y/uRqX8WG16J0rlaxcZWTYsbvIdOC+WpzOR8Rbrj6qFy3e6AetxCxNF6SN2zFHoV
0m7cLj2KbFMfiSzT0iEYMY3/mN9ZzSGAQ/Xqvoj/eJclV9IvTukZJ4yDDKdOn506JuMDA288M458
JxeRpMNY/PhMhFbzwk1p918izLh4VtgNTgahosiTyZFMjyIK19JhLSH8t/MVtUF1R1M93Ki/KnTx
6W83q7zDgPqqOqtaBALpjbGWFawwPU6bZfpNCyZ7xFM4JZ7bhEefrLhoewzW4biH/ExK4Abk7cn6
+qqlIfDaOPFMS8a6bCP/Inl2EOqvx2WpyXEXEyrFHlR4GRoBYig3ZOfSE32udsYjPDKb0AdDbPkR
e62YHNJ1ocyoCzP4sDSt+fGSSqH4kFqQXFYUZIfcCboI2u+n398wHV+zmIFwPqtO4W/Q3ThhY4pw
XevAC0rTjUu3B5ii+CCZoizVZZ0IwuS1UQ+0RM+5u4Fq5DJ8iOvOdMxJ9Akz1q4oyY/foX5V2dDq
L5h7xGNf6w5SxhLa6y51SwdhXkCazBghXchfFa9D1rZynfTd4ncSMQKWUi3WMVvmBaXxO9kWoVt7
2PBL621zY3RCYQwuPY7OPsfJHP9nVngrjX2WtABDBYQl5skBUZCjF1rgovyGvUahFpYCaPpLXh8J
glNed5HF6JAZPNuG67LwAZAgf2U8Kj+kFZ31TjaYQFV92EgxMyajfTgCitLXZCNMjqvlWBluxVmC
apA7fBmTNw97Cv91RS95XeSOWUC15dEt+/YHiOMZWejGyutJdzvd++mahrky1Kg3ydMbs4ItXvKk
TxgCzlpjgpZ3zrVY+vr6hzicFsGymuLamf7+LIzS4QE7yWJ83A29193zw2UrqaE9dGOLoMNtnETN
j+5vZzBruyzKuEwzLAPjgjKUre09/El9VDZKRdy5SMmQJcTR7Q/aYZzbTA894DTDo0mkM0V6LaP8
XtBbgJdpDugH5wOJRwcOBXfdgr9ec4X9LgOTU5XFZX1q5DQlPitWigIfHvpx55IFiU/22cakX/vf
iXG7S6POyEWpfHS74lBpeZhP42HFk89/r+6p75SycwGwkIZDGErr3rSQN80AZtDsfhMD+iibrWLa
vLapLGZxJ0larfX10ZhF9ADqg16oeynsS6ZE+JltXLD4Kx+ImIge48Hz0pQyw+IfNf5j7mMUBjAX
EjENVg5Byc+XTl92kMmeu4Z9mjRS0+3yKbYDUIMA687ACZbmiH1f4QgfIS8lqfg0go3kNEuXxoJn
vQGTx3TLN3md2qqKTAMKlbuCFUQC4oswVf1HXZZ11+axGi0klPmGOvCt1Fxz1yDBrLvcRwWQQ0xW
Qq3/yQpaiBhSwAZXu+oRgz84LtFrA4BAk1phRT431wSHPFs2PFayihQ+cnNvRJGhv7gkMakMcXIO
MTzeRWyXo51g/VF048guVDw4Jkalxcls0s0B2t2Vklfkizf+EXaoSxhAyOOM2UF+S1GMl7SRTqeM
2nGGyFy9xJUi/KKnR2SxDv1MX5FxUuDXml46tXox6Sljm74Ut4hC7spD9SC5hs2rUp7VPaCJQW1O
Vit9pML2pQYKeHx7HxZbXSqnFh03Yiz54ht75h7Fl+bbcnIT/mBu38PT18hwZbL+x+Sw+ihQIyhH
lkGIrkpS7OuCAW1ruyjPr52Rutv299yPmKFhHa7d4jzawNdoZ8D+yxb4v4Sn+YJ/MlrHWzkjBjaq
mH4Z9XRPcwX1hPexVg+vheL9mcrsw6QHvoUzbPPtXNASuBfKfDeLyYXz1/bzj/rMAT8FrpHMBVIe
ICfEIfK26e+5Wg11x6IBDjAeOkrKHTnCEjzrPsJyzyE/EdxcIbERAgeRepRWe4OqjXSvG3QXMml8
EfTqF+pq2SDK73EPXbe2aUqaRmjHir1jQLkCIF85Ru22aHAHIl5bsMunqAhpt8MroGo6YzMgZDSy
HOuIZnAUp7eXoBXBMaLXe432jpuilvZa300vXK1jB1dwxz5Js7Q7o5gM7QFRHutYWSfWYFWMlJmb
Mp9LXPlo8aHnLMv+YRm9GYCIc/CzXQM8QMaoWFI1kUw9rZnlzivNAZWTe8A9UsuQ/eYGmhpXzIZa
K556YuTvxHY7oKpALCV/A8wFM3cGH9o6Jcynw76n9bAt3DxawIX78H18sfHneKvKTCBde8OMEZPm
sd80TQFQ8CUNVpYEHvMWOfIR0EviEmFrh8Sm46IN2XJBkbsLY5V/ji+wiNoq6kpmz5t/G27rK3Jg
eJocmPZtNMfv6ZJld2WrUAgsfjyDg/AaujmK+Gu2LKlfHw655MxC34nLHHswTJr7Qnvg4OW0tOtw
xDsZnq6UIc66YNXk30lC0t3uqD6WzgGtJ6E+NQNf1eAhuernbW6rcj8NhTysETiFTZP8yOO6iV/x
KzNNQCgh6fzqO0Stxd84flfV97Y13nUWS1JdRkPPcfZrrxEzcE0x21XGV4aRdgO2g/SRKtrFEIEq
0CijOxX0TL2RLqcG6VLCByoGtM3QYvguf9uzeQKebsfQXeAwdlIVlvzZQYZnOrSktHhZLntJCmKa
FjWCZyxQCJBmbbgxKEMtyWBc6j4sN1j4m/nokijsGk3nad6uJiqztJyUinjd1V2ZHi7vbm5x7DEN
UI/jvZZCBX1r3DwPawp65yrFp0PijupwmizKP4hStW5gEgA801R3O904sUW7zE6TVx24fdZGaCVd
T0TxFwVVU9Y0KS/igjTSJZc8j6kobO51IWcnjhKQ3KhJSroXoCc41wt0eRpQh8EuzIYGfVDqeAjW
ngr9/xWUVEhX7udwlZAwhi+MAGAr7nkQbAECawRizGGDsFmnmbLGox0+sC7yHt5n7Aawy/npD8p+
XygcJaEAI1eYAdlsY8S+HuckKx0KP13narW6HqNiBiL2X9Da0ZXIB9Ik5LtrYb7X+9JstlZ/q8wL
clh8zpMlqWU6hVQnNkuR7mVpWRs6LDofy9uUmkjsUPoMZt8gcPxjolNTOF/oPOiCIVz1pfJ5YAWW
jVCM8j82AcUjCCaPBg4For86/U0sWxw9IrKXKLS5dbZrqbcTwPND961QCvotWFmAqnA4cc/dXjYu
t5HuqOpQOXDxfxApGIBtILeHKUzEzZAoRPlegb8ZXzu9+BhbaqbYWimERI1NtGMmXMDvfC80Kti5
9Ty2mqg28EvSOcYbf+4SARfzMyDiiR2W0r361UG/yFJWrZr7z61O4kVt2RyTQ3nkLvrxlNrIpnHd
gZIVltq9WaomFk9IK3ul8PRl2nwIFhZdzTjn1+6OeKqR4LUF/TD3Rl8uuWpnJ595PNzfM+v1W5QG
kvLC4FaVzhs8xtjppUXcxUrrsCHI0IzshUXrmSzUV2iLnwaJAF61WHJMVj0KGzuSRHwsRoecEt+d
/49uJDJ6GDn62pqCBtf4TioLDvuI9MvUg24tkIIvxIIjgJe/96ds1GryD9FzjksfbMBZios+NsJJ
n3SPWjjgfDcdZiEZ9LAqelF7WyXPOJOXPYHJm2SJ70sTRoefwSDfngrShAu0HLjsDrAw5J6gkYVL
nUfQfFWGJwWr/4naoF4gHDoTxW7UVWmxzlGHpIZTnjPRZDSJCr0LD/JcJSS7Fe2vKhhe6dhu4UFH
uxhjxMGEw25A4teyu3qg6x0yJTiIOHUSKAMaiZH8qMvIp4S4GPvmehTGqmwX3fqxprfnISHUwgL8
eZl2kew8MJJrfcdAbRK7zvdWWslF5kKWF8+5639UxwRnCiTmvbT5WU5gZx0BINN5xO5d8AKRGPC4
3JqWHkdOhM5REGFAWDsN9w9VJQDpZPSVYxNbpP8B+nZfvHjHfodTfZgS7E+/A0wHvs+jZzFVCggm
dRFjjzzrfIrxNwCHR5rwou82iZJvoSkNYYKezopXp5Eu/lrJJhdZrKwmLVowiZIXp0yaZsNwqzT9
3qc8csixEYShElJVQpT8k2SIcMFnyo+7QQoZEGHNJhzDUL5ofdRaJc/RV91L5+qw+eNTWVIb+2PG
3TY0Xix0Qr1z1wPEFKtrU6ZGEbNM0bfFYUmqLo9Gkh9Re2o9siJ4D67zCzzKNobFfUinOJ3HozYD
EXtpXODjhrumdEEWda1HiC82Ulw4THcctV1AMXot9kyVr4lkpcI2Dj7wS7qNw7yAR0HYWsaji7Cb
kYykSELBLsMSnwuD0BcwXR0YzgVJLlmbrdIk2QfQz3ykmMyi0RAnVyrOG1NaYJNTllnd+OAa6rYg
d/0OqyH5k9rILdhs7XSFxQ7uT42XgJ5a/Nps+7H2v1sdFPGZ8oqaRdaCrca1BfNe+LXU/tA1OOmd
jxG3k3RYVwa3iObyxx2mcmEGV9r6rKnW3ZTTVTmB38K8AsFEGU1gfTy9QEoAqLaFxXFQV4+x0r+H
oRV8YgQhX+32MMgODpeNLu+uqiQhcIx3qdJ1/zF8FPdC70c95zCXdZkHlSPe7Aia569u1HmYBf19
tUGIUp7e9RNL/9HJLW2L7uLfMV9qT3Y2a06BnrXfQA2FhtEx6GNApMl29J67FnzRPwJegRyWleqT
ulCMfRqsXQesQnIyYu2PdLhoB8gxLazIhWpX0cknbzAaGMXKS1A+Jb5KGe7UhMRh86qmtiN9brlH
t+7qLtDMOtFiqYTgu5pdUyOUzGeNjZUdPM6z2VO8NpjhAqlYygZXU2TX3UwUOQyJNaDoVOCgJiKe
Ceo0btZ7b5JfMym7uXQ3A3m/YzqGCzJhOHHjPM4g7pJ/Q/jTfTR/5gvCYtNUDTDCZsMYZipsn7rD
qjzwFziy3tN4E9aPJe7cz/B7QA8Qm+3N+6SQpiV8kPZ3HvT7Fq7G66nogKX5O2EzCXGdtBeJ+Hkl
CvxfMAXkZ4WmxnQY0tSl0QTYQlV+fT25/Fc37pxYUDRilVWI/+Det8TXEih3E7DYRL8oN8EKtwra
h2DTViTDiYw3g4cUFf1WYVk7TGY8rxmFkLKjtqHt3wq0Yt+RdrrrXIapKIytN4bnqzm87Gbw27QN
Rmr71l82u/+lIbpfS4rqnrDwswV+Av383HZTgmkw+RE3U0XIFUlbXYFOHe7JMifPqNvcFOsPGrAs
4KgsWWTsbVR+y7rBI8SYNLc6ofoVVGNNcvm76UyHLKzZsSJCEEnnehCqW/JrnXiJf7F20SScERVJ
Pvy2PBcWoZU2viwym8fYyJwtuqo7i0uhd47EFclUcchRBfozMc45KtwB342rLu3SYIqLabiBcu5R
Z4R5Qs+5a9WRlU+6lsDj/9YVB3A2697GLPs+7JMp0rNtCjiH+hEsigYy4xTP9ZS5nTSgSpa2amJS
I7M+mu+3i97fgM3M6kGB8HOQNl4sIl+3Szuv4JQV5WVgFBovTHSycLtivHYE8Ua2t8w23KTtU+s8
z7Cvrz919GzSFus+Nh8O8mmHenXLuQJUgflOPKoFeu6rvxJns8RPYtyTIBM4m3IImVolBYTg6Ebv
NIXaxE1s/2yeyHIaFSb4zSU3aOHAoCiHZWRl/7VjYXLmdvcqLV+7Xo6L8hwTEzxeftcb7z582KJZ
hCJyEbhP4NIGR78WTKWJJJR0s2k/y3B65vCTUiDFX2RDi7nOAEKXgktnL4Z2rYfp6FQcyhT4irJi
L35e5xCXTnuGItG1DOwzBtD6DwFQBBiMHHb5/eGWOxLvmT3euIegme7oDg7APowPANtHLYsAGAWz
MVDNwvI9PE1YCdseNyx39LC0EWWFbW58VajNQ9uYtF7MIF35OSiY5WQLUYwZEquWBvIWoFFv7bsx
jJSUjnDxR5MkeS1hPD8OYW5VZOE1/0aletGIwliOBEybwgHXjiBCWDwDnQO4ZDaO2ZUpD56lbO4b
1gjPRirPoAxtCy9AEg9TctGNobax39DM/Fl6naGNMQ/a+mHYwsHgwq7xFezA5FFDML+TQh6OapZ9
gZW6kuqREdgk7M2khATFGFxwg4oBiSvDSTpuUW8txzmK/vXLL1PhawoHOyv8rZphL5fQR4IDIbaR
0sbyB/vME4w9y7agfEGrXJoFxLYWV9CHUhTQUuxfJYbt6R5RKdUNgJ+mXJQLYG3jjNBjHcgAMafe
GitMLnVJJmeIWDbkxErYUlT4qYy4pYdXqg77GfBPHDU0kfcbEN9SRnz1fBTzaNSW4gp5nVeINiNY
0vYXGpsTL+axwIuO1OMGyqeHW3T9AgT2PynMH0Vl256UZyrbzZy7OVYrNUkaA3pofRTq2lP76KpS
wRx+cAZK2LmeZgbWcQvP0BIV9eggEySgYRGfxRcKoRP7l779URUzcZXADm+U0vHmEpQJkaNBqSat
w2VVT1cyCgLalV8wkOTCArq+mhjFMoVWLTS7Dz67kQYfMpc01Tm0+NHnvfhvz/b416Ud1BjNeBgo
XggoDJmttbRnly6GN1GjM8ovSDDt6iujogeN27fBL5K44SaVYHhghVsQZw8GkObJGn09EQA8UFkG
0JbiKoINTjXpGtzVFCkaUSBMEU0cJinUVSyETvWzI90I3JaGfQsZ5bjokRn+P2Ew2IfKSlZaRACJ
jLDQdGvrKPNCCWD6IUE9wFuLDU3110ZEBBAMurU9V5tLHTuNdCSwXgGjlpL05mAsek3yWe6aLhDE
EzSEECmvqTfLg1d0X97kvXBfd9UZeZ221jz27gDKKAzEbB4pc/ZfrTeUB3ohGv81MOaejQVZun4E
w5Q5D2l7iiNoYjXcFD4IEvAK49ffS5gYedszrX7kTXkgIwEfV+dAlzz7ehKtvkF7CkMTlK5tlDVG
57dxz0l2LLfHAMXeIOXS9A4ePV6DBBLmoa3sPUIyslV5O1DGHWyM7Fvqlojo2BpA6Y3MmFfKgSU1
lJ8bzolm37jxNSPxAGpkWsTijEekbY0ZMrNEP7o0YsyzZMg3R76vAzBAxcyO3oGSAkFRDGhnKuOV
0j1UuNLVCIT+q2hkkopLoIg9R8j5UNxgdC+aL2t9/vaFC9mVz1ahXs2jtW4BPVxcP8MDyMaN5was
p5TCLOKB6D84rFOseFWB41KqMx5e7mWHFHKzsQlH15076+iM7xMDcDf2YOQ57/XpXhLo28+x4V+Z
awgi0k0UxaS5E9iEBmjMkctnyq+eq3ecNXic9vXkRNwBUS7jby5sEAQBdB6q00HsZB8AOEG1G+0S
P5e5DFQiRpHdWLJUinjtViayk8IHANHecWSiN7F98p2rJuRaUbHMePJ4jtWENK9XmNQTIFD5DHLT
5Gj41RBwyNWdruEMRsg4T//jNTO7t8M8VrKhShtoB4BT50pfiPnnPXc1AzloSsfYYkY6cWrcYS7i
MwHi0xBS3q9gXCTW1yvlLjcYej9PFwZQqTg9e7mEJBsNACLsMK1YyA2adymMVbkTcdGUd4PY4N2/
waqhtgbRSzo4YUvfNh+JIu15Y/WnZmMPdEPCbiqQtGq+OLp45v8Bk/lBTOPGOgtuhrIsIDUNMlfG
vz3RS4LT4yQHP+bnw/5CAEup5LY0noHfOQEia+iarYoH+YFuzbHYyh9oNnWryLBViUMOVgNSpXiG
++MK/JaQjBmI0TxNC17/f8Xsen2Hchp6Mqwd42P0LggY2QLuTH+2BAOWE4aAt9bQ8iLTVHzfaTYa
KbAfI7tA+KeCK75VfoPZqYQOT3b4v1M7+/3C3aPH3Iu8ZsyRTa33Rf4SO/JH3jyO5kNR34IfKL/d
aBVTjTmjXpBlV0f/FrMWk8OxVR5g8uwMRvbZ+wEpQCZq8yQYLFL8p1YgDsIoy5svy3JzTyxNbSxu
8fs+M4IrUuNr2m5nLw/WjkoT+H8kqwEQjy7KYYUWBKQdSlJMJTgmWsYYhp5S3Au48wUPkQDeG11M
nQSqCUnmSZgSh+HL3D+oA3AGKf/NI29H7043HqgHbtxsJsCZIj9SzOepB+8a4SsvQTWkbUVct1y4
Dt8zUQJCbddZgezNwleOT87niCENfSdGO8MTUnQ/CdV9y5QlV5++rxvpNT0xPi9bi/ZTkVKNQ7mO
8aKDzBCpK+BR3ZmUBu8LY/xj3x9gYTyR9DPOy3zZw6CLfmTU/SgdW7SICsMrF7sN+n6K2yAZrFe5
Es1ZApbhr9JiTGkfu8Etd3OG1CzjqsqaoDk90HQITF826d4nGjNbzy9M9buEJwOSoU9/LLpZy9I8
FZvTTkTW706UHGD4qXQp8DDsIMKRGbAtnelt24E/TCpF3vBSL5teBCYEl6YYP5R3cEHXfN/O7aI7
IIR8LfOkxyF4uP2chB4zH9J4I4fYt+OjuOPDeahKCbB/HgNtMdx/af9vzkaSnmmVdMu6Chk7HaP/
cJnB/dUQv5uj+EF2wilELrdBGCXNzjBfIi04fECxTJoUxwFhOZ2Nlh1v4wlBDwmwizqtP+RouDn2
wrMwRWApFgzEypucqjg9jkRknmdgqz0hwMxWd0hEuwrVB8cm+YzRsGdeZDJXlTIzMxFQKImMLCr6
nPCFrD3AZmrTmrsXL55ZmuX+yPwMtTnsASPXuBJmDs0u4aFUfO0+rsiNpwFbqOEB1IDGbK5aigXA
AxIqsFEv5zMdpWN5PufStkA8X0fqZ6xQwd3BcvzAqZOOfHcOoHAJ+7/3nzCb77Uzc/9lruKHgCt9
HHKIARoi/kN/Dc/rQ7KZ15L3/KmMHNjluFMgv17sgk4nYXVGQGz2UVCHcUaNGsZq2ZWSdEC+13pB
3YxB9FJ3kC6FX+l55TyIRLFjFTIAfPtS3gHnipe4iJBsZB6nobhY8GYU8J/KgyS4jdFNX9an2ftu
dluvuwmAStfO9PrGhgz8L7xxDMdsv+aMTEPHrjNmhSd4ZRPmrfAxar1cFWzcMlAdmPtu3Kho1hrs
Z4W9ji0TIH3F9kdKtvQUh4b2jn9SfMZDinDFpZghR0kgRU83vIGEh6Zc2b//NOgAeq8pf7Hd/fBi
VgHHODGnVUpCxIU5S7zPgALd9Oj4VxjkpuOrZuaNR1fjyO/oYHmNJcSvZ1UL7H1zyYY6nmsHPw+3
aXfHZt6oM26R5E9QQyj9YiIZTwg7pVrniGoNYvfscLpYhQWqJTxgbKT2EnlXNBBl3VQdv2+xgLDW
7EFQkdGCDBeRP8eZRsFhZZs3bwYnBmjex+fWScvbnQMeO64POwds+XWFZg/D/iE07nK9xaaF7yWV
UyEIKyFf2ylh2uFtFGPikJ+LW/wa0w51XrSXbifI/KFre0Zz+tsronON5BGm754btJpZXfnvYI48
Tokd4LFgJ5ELtVR25d4EPHa15A5NGVAm4St91+nziwIV834zpv098QUJ9l/DnvhEIfBuy/tdzQc0
51dZzGxF5cSwALMTRq5nEJsRSaL2fymZnFW86dum7LcumkwyKzABmBqPo+Jajd2Qcaj7MfoOsN0b
2ezYrbu4wkQFRY6I7my9Sn4uf/c1DiDyBmd4qonkVW59mAIv8XVcKEsePCuNnebsWTnY/HHFEwcL
3gCOmB+i03ivuPRiq6t5rYXH/KrEzPmegu83vAGEg6DWSZRtnwfLAJ6DDKkabIuWeRAHZTvsk0ex
px3Rlrun4kwKXr8wFZTiTyJJF7A8C4JFCCJetT7mDkN69IA9VaCKeKucOY0SPwHhhl6SGFgd7nlv
FlmdYDv9f8FBbyuChl78cJEuf80f8F+7ndQu7EXgDHWIGndSCwDK9vcsyAoIpB3RncLA7ALboprm
f2aBzyvP4/jzF4zbG8CqolowL0Ck85EnHZaY+ztIb9vsw5dUqnTteXOyWuO8WX8UgOAkwBfCTIyb
qJHPfr4k1dABJRPd5w0VoE6FZLwigenaXA+MZ+uEMinFMh9DhXbBY0/G6FkaDJzsOeK9G4ZZo5yX
XPq492QCwA2nyKr7k3QX/mY3ubuBTxLmub+0OfIPatK0bn3am00CvRBSOPT9b6l0Tc7Oo7LnZrnZ
VGR/keNBcmSqYaMrH/2w9yM/zI+apwSRM9d5AfXNB3UbcjQyVWsfrGdS5SGEe4TuAhJQs6USXmQb
71r7t4Cu+pjeQQGeUmRiHFjPtLAWTBVrRuV3etZWt2CRb+wJDfSzSbaKFnfKQRXiWjvk6hoFpGcl
PqQnpNN+BOHODZ9KbTK7c1kVZVbrs02opE42aGGhhsbAS9IjUlfQTF2uSFewFm8WD0msAWvUu+Qp
1Y42+2eOzEBgH6Bkxk60jbjSaY9fWRSnPh17Vbnc0qmvtDMkMfg48YL0vj1Cdcyi7feBd+UFyjel
VVF0EaYLVg1lY8aHoEVUeYDQvSFT7+1vH87vtBU/R7RpDXY0w7MY4wJlnPEfL+QPMUax/RcPStfk
OyOwwrZhK6+HceTC/7f3FpnlnL7CMJfLaTf9vv09dLfhQXfNpQfDitYpkrOjwqGVrb7mAwJzwLH1
TFGCDR/jE4RahwJf0ou4xnPWjzGsXuUjbyRhFOutiJ/SEk6Em1s0d28Xj9mKn6ldJaXrau1z54Lo
0AZKvMZ1GUQuSiFHWk9kqWdDvp3iffUBlDPxd2fxIC8ri/cEQ72LNw8F2T8/Run0lmLU9KA5x65f
t3eTJICAaI1O9bIPOc/Tt5oSMVXQmJ+lNtrMp1OPhnJXuzKFCII4aYe8+ko8kh0pDnec4zayxjGZ
waB4TqgfLzdcBw5Tn7ZJ2cvmuV4k48SY2W07dhuvxh5xhvKWPN3MNVkV3jny7hAiwqQoKwUEfwBw
pZGLGb9rX3zsViNL4h0DMKzZhbrBUXuFXaQuH1raJhyGPi/e0XiKjwXpRysp6MGnXO5huOaPwirj
Me7DcpCYOwt/65oZTUS/h3WJFSIbWiO5w351Y/AkHgdh8hy/CgABwX/U09dwBoIFHSjHQypyCQzZ
rRP7KpwfAuvCO4YsrRrfps0UacY9iuJLyStEVDHzgyi67B6TzzOd/ePkvDQh7hO5PWPN9LnL0EJz
XKYAaRIg9cai/N98ie7ROkRO4I8DGyHYr9qmjbSRhOmC7pBoTpJieHjRLtA5rqWjD0w3FSQW3RGn
21mdJKW4cgIwZIsCq4wTdsZIwF4gQChScUvqWa/MWR96bdXCPUhlQ6FfXwS/cdpK4pi6MJXvWGsz
EmX56gsz/4phW1+yWufOZK/giTU+Tp5Ul+4x7OffsP67eLNyF1LQe0FmO2+NCPQ/SWlUfLQIVWZI
30BVFLinUnxqEVidQLOqCulFTwZ9oLeXqj9PETpRgIUAuFrShyawGvsp01qfeMeCN2sa89pHp6+5
+pxQ8ALJoGo08q+MecJCjMgkN1v9U+klCblJHstz8ZHo3bmrk9qyRhR0N5WytnDVaLQ+19HfS21I
t+YDj/jVwByYqpCTWEnZNukS8X2tvuZVzbHyR4v1w3wbj3TVtNxp75idcdVr0LScmNgDAedq2FwL
XtiMjOH1PpU5LhnTPR4OAGj7kTxrxJaUqILTbbiEDGjzLywmzzIW2JQ5EVpSYMxkrfd1R47f/M9z
ozLhcug5CeG+qcy4l2nynO4r+RD5LgAvN5deOgfDYbraLMA4B2KcNaVJBa8xaIG18QrZeXQzT5l3
fpFCFKmH/3f/v3AqWUt0zYD4dDRN2xPiqaB4GQJ4fiefPrMCs2hqXMw7mzUt5FfsL5ooCv50dxOP
dtzLcl3V24W39LElk60G3stGV8yEt5lKT8w9Sd+hohH+17rBZ730gcWubF9FYoNQGh60Aa3HLUP0
oYIUNJ+F4WUpT7gSEfZORvB+3Fesbtnf4KFzTUKoHe/rdqfiGIto/wHAKV/G+b3E+4KVChTfgh6R
LGhiPE+/iG/siSEV/ufpn/O9v/Y+av999OqtEUjARvklwhJeBBTK1+TF+jFuTCaIOPFetDXDKiox
FOFmP2uVoch73HyHyPugeHvfmFpViabElr3FBh1ewRhgnVXKI71rhy7bblDpq6K46dtldFaZYXIr
TaVC22Tf6Kb+flqIkGknZePIrcI88PBNvEKDUFkPpw+09WJby73lgbjZ6NC1pBK0NDS77H0ccun0
5cf6zwcUefy5dC51hENrVJRKxRLZx0+W/ldT+gJIqyL7GeZD6j2lNYhXNAxQ/WyotSd1/fPQSKOU
zmMVjOjvAoCR6yC36OC9LR7tzydurjZawHiRNiTX621lBEpCp5sBM70EVg9yJ4joypRogCRRO0Os
b0BcfUzPbs7ckrJ1MEKfxF686KGaNWbNQ0khaZeak2oHyKFiLRasUYUf3s2CP/frUime55S7nBZI
Zvz8NvusdiJWdhoWOG2c7s/9SWbq7X7dU2K7PItZZFn4e4iKoC2c3W7DqEY00WvVK2xNyMCd51Zz
8SWga/u1tDGC9DipNHRBiQF9TZQujDqFvH4c9JlZO/AMMpD42QnZPL3GI/duCRdoi/vrn7Ziregn
VYQzFV7ezQBlzsnkJIOa5JJFw3Jcvq6a68Px9G+A7FHTY8G+phEzXjQP07mmjkxL2bh+RCUskRVv
bZcwdJ6Rkmwv2bK8dHvh6WjtMXtk146zFGpgVGtF78LXFYrr8aU7wECIK/9/5R5xP+oOk02MHBs1
z0I5s7y2xaVbZWPiCJNOAW0dkcdVIEGjEkiP7i/3pcrb00TmPF72sg5xt9SMDU9YlmsRzD04tjWN
j95zWC4PdPotNBDCJFQ6bNKOIsYEiyLO4Ykirhk5FydkDI5B7BnBcPMqFjeWIS7Z0WSeM8zoAmj6
2pbeTifIWgjI7/LMjuxXqSWKXNQQV6kt+2/eVNrNdNVrkfUkgyFlLz5zL9r+1fqyzAQhqanqAze8
T9qP66czSzJnkng3AQfUR9znl0dSFkIfZtD/StSUhb9aKQ38pdIu1tTh/zJSsQdr0TWk8pdV6Npi
iWvYhF+X+PZOM4MI2hQBs03iFOqeQfzrDq+QTZovEwExmXJJNRmzjR0pzTzQT6YR0EJNsiz77v6m
8J3bP1g07bSeyPTd/dXvjSbiWdVmoNa1DdSfUhpUOtnBL+00I4V8IgmD4BrBYHiBh8Ik/cO7tqBK
xMy2VfXEeADfEnLbzjAh5o14qjj1ZYCEgwLmXfmzNW+ZZ7TBNQxbTHQpDmw9LH/v5Rl4LsbrzSrB
EOgNEqBqpjsQehpFaOIdHhDd8KZOcBJWCZdpLkDt6DI3UNWtxjPejgEHddvWCNWTucMXaGu5S0uW
r8SMF9YFxcSGNg1PjXk6y5c4IIu8+ETYek3wUBBB4GZm4MWr36UTiKSc1XD/RA+Kzg7YDt126YFN
tRvwR8dp3fKMPqgRQU/ZGBeVvSTU7y9juVNcTf6Kivl5wYfE2pwu0jiyMH+mPYEBgMCrGgrFhUVR
qiB/Va99QJk6QReagjyie7w70Q6P0zmAGDFG3EkqDPyV5z1aKGhHX5BUjX52awaPSdB7GPZoDCpo
l+zri+iYJzKJfhPO2fXfoy/4oU9k9PiIysggOIGALslIv/xItp3vRc/3q7jiiILolWf/Ji1VharW
V6dbknlro0qL0/J41jBC2JBgNrLruDv+hpGbiCKOA8Ow8Ax3w4kpiBr7b9vlRWq3icKC9olgv4w2
K7KA1Qxy71WOFNDx6cXaCCnxX6yA98vgQVMoJH+PhP0htH/4X+wVMLBwE7u/fk/MBibjAfH7SOUL
9bhUSguQ0FEeUoSM2sGrrVu01M7EZ+TGPaPdF4e8uo3kDUVcPqMNj3V/QoUc63EOPwlFOiE8yCaJ
YTS2kdj5k6+dzJQPsX/FSINg7+WoCrU40JOtsgBv+bA1ILOHIIZEbfopqXUmHyhATXsdZ4k+dCNY
9PXTs7qMiJrCaBccK+3Pu8bPucRpQQvgUgbUaCM6jYSx/VNUUWRJ7Rrsb85kxsKqRoMkJK9tLuRg
fjGzig8r4d2TYaqqcipRjmafIqcATKYroQYSybtXxIUvVkzqdQP+hpnrGNvHPjhevMkoxTtpmr0U
hB96kzkPhP5JQvVi+FFDxDh82IBO7cdTnYP9IpaPH78YN/oPCzCUmGiEXHqgXj5Wb27TTLBBfqH3
VCqrK5giQvvEpN9WjLM3DMhKqLNS3j4AAF7C4sGNFs6DNFGSe7WW5Bt8rEYyVTSmp0plZoAvlWBa
DXTHq0LsqPnAMPD97WG0Ikyc5xH0qgS7848UTYofIszfiiv/zw2VSiVOoJ5tQ54wq9XieqPYongj
rpipDqSDMT50ts8+Ws6+ItDElUdr2SVHZWFKmzynbaFB58t0rMxeFRn7ndE9FJN5hlZfzQ3Hq5mj
Ypgq/zWL9GnYnNvD8qpQ/ioeTTTisvUHodCTRxe3k5wYc+SriIJEC4UXE8vQlCVvvMKKuNiG+dZe
WlWXvLRhIL5YGslQEq/yK0F1/P63PCvT0M03n4Y9LnxYgBD4jmXe7RS2QLyVTfKKCLWg6q58fluc
0RRq7gxBL3S37T5u1+N3UZYKfQe8SbJF1cDEXBDOgOZnBCYqTb99ED1vLUiaHts0h1hceJKwza6j
6McrtEdHuhTZ66JOe4cGLiCvAHED3cacYFPG4xZw+aqh6w+jBiKkmiVSwwfK0bMPYgIlxdKg2WzM
4XyGqd3L4vyJsPphJlwRnc4NoDR95XmG/+F7n2+4KwuNigaPPK70wpjeEXx4TkrTAjNHjCNZwKCT
roH7u1Jf3+2Ff+58Jv4WU4YJjA4rFErfH32DKgl0eIItTIwk1lFK8OiSZ43sxbe4ar4knH3kxw55
ieE9src+UEuwyJBIumef31f178tfMxbNQnziBklCJSYWNhpefnrkXw5g1kltmANeQPmctAxVGatu
gtkFyRemEqoJPce2dTVPfHkhL21+qkeL50UOvSLQo1ABpDSHEYLTD/4zkAPJyLWkuYOqAwYnw02J
IJzE4/HWiaiNVuoU+ICThTTOqcF6NhNVLV5yKizI9xDiOYLaWWFcI19ccc9jHnwHiKVITAFkc2Pp
jIAXDmTdunSZOCnHd+8b5r8OXANGlSIxJZZnDPszfQLMpeb9mfAbMhZWjEeiDzBUYKth8SUr8OY1
2enSbR6DuvmVVhKjifQCFJ3jNS4Bf7EghJQENN1FikU2FwwidH2EeXl6lKonDJ5Dym8BjQrWfHNR
GTclf3/YGirHZmOQMznxdsqQdcNpPPZJErm4x/u6CtxlazptI6txttzI/llHg2Ogien0mYqAFGhG
6BQmMpyb7J+qY+xoFIRQnjeIW90ADzs2xSpke9JfGi4kpyEp2bzDnVk6vdUVoPOq1kbgv+TEdQ4T
mDv1jhwozyF060hHdnqsEdYnAIgPAlaW9b93Q7MpL1dCL8gprCDOJbWUCCm2bO0PF2hCPzLsye8B
0DrvbP/1FyRzLvL/k0ddy+mesr+mFr/NNXDLKJS2a1KaEuLJKhnQ9AYEr1fGx6iweiuafY6m8Rg3
mpeRp41k0qCuslmyMrYJESskjUr4H22vnDTDSYRMSWQ9WbZWg+hFaaNMxE2PcKU22h3QHA3cZMgN
YIMV6QVXqsBSSPmXKVQiLGGunjeV6vogQ+7qTCT2v/0fr6wMskqMEY0gCo1OO4en20u7YxHmLFnr
s0T1RB7gUSUTNPmBGH/PO1KiPI6C3LYzFCK0hwTX9Xm1E4sv4ebyVtee97D3iyA8ektPd7xEYh4Q
ojQgLhW27tsUwV+Y61iAHjaPrqwFZRsM4z4TunG+zZ6Hi5r0UYE7cmdmd8U7JASwpmFUe6Q3MECB
AFtRkAC1ZhhTVnYpWdlSv+K6VubCyoah8al0iAGVlJX3qp4oqVuQ4/jFJNEyMLsir886fiz5xwOA
jA3+5wqa2BUnphImPlVPDY9RDWH5oaBJXnsxgEfELrkL60iqoLdq79w6Fi/rq6mSKBRGEWsz/awz
Kz0TnnXnlqv3lk1dB73AU1VB7XJoqPRO/CeYr3IkS5xOuNk6xOQp7nyTVRxRJKDWlTIXzRaYSiag
4lopyvGDQNFhoHniOkJaQXEWYB4CVSKh/rQzkzailYoajzT5+wZDCaEBAbYob2eBa+v+QAjueoVZ
qddBAO/8/klTZCtQriFXx8luaCF6Ykj0cR0ZArf5OcGhecTODcJFRAN2sed/uSh34Y3wuR3e6LRv
AkzOLhBV2mE22sPFwu+cwb/vR/Ob8I8ixKfnzw/IGD62+JjtixLij9g5+Y/WNtxIqorddny69kLv
7xpRHfXfm9VGxX3Tn7onhIl9B9SIVAW/h9OKd4k2X89wG/ZtJRqMhMC9fMKtfbyh6+r3P8AsLXTP
QzQWETMDX5XhYoEYAKGGxjlS8VpxNHGLaifDpT4snbHtjG/JrhZPVHghgZkHEcxnmfZ8ZioFWWkh
EtW0erpGp0c5Wka4QWdzy5yPUAU0MT5c4lS/RbcYBgZl76LHkNgxrz0x3bZZScKsKWJUbwHAgcRX
wk/AitA5JnAHLPI1yImZfHBXiaBY/sOYxIM2tnDsmFzCKpUxvm6gW8EI65oAzHD0K21NY7tDbWhI
kjS976f2uOOVbNyo0ZUNETA6xjPBy9YzAvh7PEY1wkHfA39VAztnR3x8xM0ZtuKKN692K7ZWH8Zj
Au60qeiisCJ+9EVKPrUTQ/+vvshBWQEin3YHb/cqWd0ko83GFDpyyKwers2OiG5/vI0tGSF7o1ie
WvCfP4ovzaqaYeONml/Y2Gl8FevkRcSkO316dl1sbDNAuN2M0DN6LgZ5TIhgKeFV6UYj/pp4x0UA
lAnFD7D693rDzuGgaoEKrVeiXJvd4pAFlBKD/CKC2BdvtW2B7V+47LxZRsiTWWrEetHdLYEsDyOK
JH6NS8bd6wKO9HSAUyMgG8Tbgc2imuqjVgmRRm+mlb9h3QD9MnoKcpD084YbrG0+rkL5iWHfJ4Ag
yMlHoG5x3NpKjPvOBu9dzjsJztRn8x1ol84X5PQksRi1uluzd+p1+ptmPzEXZfNvfxzKfPgJn/Yh
1fh2oB/DSHyyTpLUnRcTtPZfLEE6huZ8FbvKHZGfDX2EUPiSxXSN7RqLwIHKx1ivFxQ1xjucxIdY
p/4oYbpVGFOvawHIndxwARotOkN0PbOcvQMcpVuwpkEdyvVmNMwTyvfCTbJxd2gZuEqgZnZawuwf
mCcRvBmO4C9QDF6wDXZVFaoa4/yiX9rb5BpFH+YU5WqpqxQ7TGgq+KhMamgyN8fxBfLHBJmZKCoD
7gHp0skmdSwrnRJY7BD4EfSOQ3QHMcm1ny6dLhZOUU5hmZzfJdnVM7UpIrcLO5R2p07rPJiuZxqX
Va6ypv32OzWmAQICxBv3z6daS6yY+xe6S7Na9Gm84l8vw3yeKzXlfdN1+whjKNSO0RA33iSu+T8c
qhIS5x2/bWy5TRKgtSxh2dpWRkkKR1DpDe+PRX/EoAVWL7i9J6QAehS2cozSlhWylDnoupSF3hU6
mjJLgACNK9JgOdeVo8GNhfvoxfrUl1xefnSIjo2rdHXBLRrQomZsfQR5Cl1qFgwskC+5h6tUbsgp
/rI5W3C0jKRJ9qzIFgPovX+HXzdHSs/PNViH4aJowJW9BVbv5WIbG5HBi4fKSuJdBo3n4YTWC2Lt
jrIw45PJOGlXGqhtbCYwF+cvscpDQeiCZ8xaf+GUQ1dQErHZQGHvm/7gfCjYJuG4r18t9dVhFjWP
5PdHoQ+/fC8Af3xm5y2HeA3GSc8z98hlBohUXDbv6umkTtuA5kj1GCAQISi1N21pNPT/Fy4r2BBX
3k50BKGDprVsIyqt5j5lazqJgcGVyLXIKgkVpV8chP1Olb9vqPjIQ6zSyjGZ6AouHeChzeuXEist
cP8OnGrjmAZ+jRAjUpuD/8HuOR2hMnmMwHZbx5qRoLYpfBLnqnVyqd6lLuimOACU1WAU8ICgO+2G
shie6dyVuQ3WCH7dQgjXjKnrTJwlL5WxvkGdmXZpuxCHiSl1uT6FIHNSpst9WGJ5iUYxilBVNhTr
LyIqyzvzISmvoD/LGag5L460/+9Rs5BW2Ba/H/DBGL4imyjjirt7dRDe2R03azSxh5xFJX9oojAK
Q9z9VAujlwRiK/hyjQHqzAF8PPaPpfn9XepQGr1xardPDmIu4j7rkdi2jAF+ACHB5pz5FXOhQfF8
7zE2OAHO5b6FWk1gbGKy4KLvG1PSyDkvSMbLHBsKHkztY7qrE+Htvxh6Qck7a07Df6NyUMPe5wvl
F/l6TbRJ2bHQI+2Pv72hAt/cd3+7xqaggvLzXKUHPyRQ56ssO7Ano9M/sMwFdA2xIJtf1IB6WfjQ
3bW1MkrreYfO1+se/G9gX2QOfRowgOwVkgzlLwXYDvVynSPcYsxP+54ThgI+fPOXrAO2ioywfs78
tJcWjTcxVu0BqdjNZQsxGMaguqs/3v9uXMZ0agWQFdQMkK9xj1AYZ5Xr+guFi7Bue6sg1jM3P6HL
4qkyglRM7kLrWHu6FmKfxDizA/MdjFmAysgroBmopbN/7w395IG32iSKDmA9Yxjz/E4GQFtU8kgO
sitSA6y7COLpVEyONoDsMe2fJX8OyPLv5BMYUbG/M+bCAjSiarwUjKq1XC9sMle/3ciaVHoHr6YT
yLeQaCh6vdl3TFiBWH6ibct/2/qvpfeM2sI+NzSPmIXAGGy/Bq9KqmB2mV1yn1bOFjn3Htmf9bwr
bzyeYYGIV//o9RKRyiVtDi/6UoiifwrXuc8KXyCX9Il2gFYBQ434S3cAmgi6aZ7qMSWzR3hTGo1c
7O0IE0e2mNPuDYB35fviGTlmIKV0pp8EC551qGHzpjEnXzU1C7NH9SkXBmdnMmwclKWXBvjLc33E
EnO6z84E27qHb4LSTq8ZK5hStPzn7lipp7iEVnULEEnohZldGpQDeTgo6EHEo6E5HGimEAaAvqvg
tWLye67JoDuQtaxgzo5e8k4VoCwuovtf+XaSszJ6U+YCA0F4kab8C/N2TwZaJAR2yzsxfoE1j/jT
+L4OvAfftRVxQPsRTYHG4B/JSpZj18FQAVfq6BdE5hnolCM8CcO+fiPFL3f++n9qhkBPAVo/ym3N
R7Nx9g+8YZcv0W/la3rcNRxNSzbaQsmszqunufmiuXMEO/TU9TddfrtNXXzHG11XUGy0W/mJqNw+
ZTgAkbbJnaGIHTUKtm4jKLavLKKuJreWLrp6uHv1Hnx7hEjSykrZw9dOe4o2bVIMPYQRKQXvUouy
FF6k13r5VwYl9RODQ++zxD4AE+CGmLzIR0Ke7Zqcr/g4TStHdUXWJDBMSaFPn1uhypUdMfCovegP
kwVG8whgtbwvn2eXvjuLJvkv7E/Ja7CmXBEfl0ZLeId8yS0QFbgJ2DEAldVJjJX9MpmnXIp2RkBl
QXprwFjZ9SWaHR7ufYMn3Wx37lf83tgDbtFufJkYSf/GYBgbZtGLb6V/U+DUb/bf0aOqRZ81JY9V
/V5EjkzA8B+bxK38fxsZluMjYsdaoPtJFA7IQW9su76dln7w6sBZhUN7i/1MJXjSyXcKC+xAKX2y
JQY3QDEG/cFW1tDAv83+F2/hFt4W2GXJzZS6kC6ChfZrd9FD0Jtfruwqbyltl5zFjFz6tcK4W+sR
Xil3kkOk9ZQWU6+/cbn1SJWQ7uREF6C3IxDrddSpvR7ymPwfoxLBPyIY9wbTQq0cd3JmGioyC8Hg
rdLUVWRlac+0kyzgANZwiZkd/UVdQDCRs8XLk5exEM3+mxtaNY4SaaDSOxsA4Lmc7sqRDX3zXlfY
kSNci4nJgKBEyTwTTAizxaI18RJPnUVG4xag8lkmLlrPQP2EeWKebRbYqv0+hzcU9batnh+d0QfH
FzSoJlLiNsawm/L5uxQNx3dl2sWNAzXKrhLK4dm6ITn+heCUjci0sKqBXBqP2UDqvjhlfWJ3FZkh
s/8vD0bqVlS+f7UVfax9GlHZWZm94T3CTtBUghmcV2CShWHsGD5+Y06xOoZd0XvOAtYAtldMT8gw
20BjDo1iXiSaLhJIHLQIFPSILHt9wzxgOaJHLUwNiXMFhAQjBAtgiYBm7gvcyv8IP1O3M6tIYvXa
AYJpEGIkWbnsU12lfzBSgyx58+DfKyodoYbKjPwAyECwcfcNmeMDMZ0p19/JWAoGs9HhlVB15sMG
LLfjfTx8CT1KumUOeVavMzT+PEvGCihE3byJdZeZrefFXYvlQ6w4CmkyPEopTk8zsB6ClN+I/qnH
CG1zAr4+i6IcE2X8G2uWUOAFFyf/Gi34Z+yPuyCqqNYWcuQ+QRPJNBnMHRiW4lFFKHmLs0tOR0Zl
Xm9c4XgRck5L40OXTFiJbaw7XQao2WzWpTVbDoYHY4os16czo5M4D/8ccSw3TD3tIBlrLdJpif67
GYLfguJNkbcfw2XzyHE1qD2oKRmX24SDBKrxbT7ZOm9XKrTjnGJYBSH8E4qSqQQt/3+QNzjbH3HN
NPD+bruQ/FGPbh8qTfiHpvRhXiAE17cNFmubmnNJhrYg2QdicGa6c2oEb3hIHCtmubP4/6BPTech
BNc5eptDqfmh0bNp/jT9dYE+GaIJGFhkf5Cu/z6v33jpZXNYnrTpXkXpV8PPeOUDQZuTxJTzpC+A
NxNzLuhJaX48W8UgH5Lcxq2KML/CsI2PxouE2UGGYvMwtSHwr8SQscfELLwVSexgczbKLjxvR1cr
p062te1fk9xPSGBufT9s+t+IdRbwIl3+9Ik4JvgpGVH/CRgCca2O8n6QX6kRvaAUadGAd+/Nmrfp
sHx/k2wp/MqIZYT9vWPTWs0KsQmut9ByvMYETzYpfQAMILcO5PRCrLFgKfUVLkBxLjYmGT5gA35c
F91ECA0Y8omfibQeweaY+sjeflVf4GvY3gd0UTeIy2ecJCRJyv48FZlhhEL0i6n0l18uOb9yaBQi
DDk3p2HjjWYCvJ/Usp7Bg6XZ9tsGTMJnN85PbLuggK6h2NG2faQd2LI/aPfJ+nNjsOTWAyI5mqP0
MBte2EH/9w9NFMedrmRX7wal1wEsXp1e7W6bLl5t83b/gdrXyaXB8FTnVoO2hn/bkIYDzgUPn3UV
VoPfZmWZZvdpXMvzl1nlTbw5+5XD5jqc3kt54tsOfqNPvxv7NbSBKt39DF02H7jA7SQpAJPNhGCG
IVJSEyZsZsoylzk7mfwgFWi/oryriXL4iuKzQm3nGuLdE8DXzjccdrHjGOeOBm73RP8AMxt3sN9c
T0R5wcVOzc2XP1qT326mOQPjfjhYdEnjnaJ15psggunmH7K7zFfFC3e64d/+nG7sDe8ugGH7ucy6
5kz56I5Okc/AVnAUfCyUUaRRoV5CJelRcMDE1kpCjnJ0RkziJRsVEV13pIYoQ1mpu93ZQk4ARVSE
6IkHdCCo08dcpma4ois0D5xaubpm7a9/I/aLTX/ZYBpDSdgVLjYE0zAYQkEMOYorYdkuDyorbTP5
GwGOLA+uSIX2wn7vfZYbBXBx1ujU79E1Y/I5MTgD9gG+EQPhMEybsZuvEQ3VZv1dm6M+bQSvj016
M1tROSxqDTfqSYhN0UlbA+LpyY5UOlY9e1hWiRy7jrlPYIjam67zuK1k8weXbg4KDEWhTtaYbtmM
+AyOUf2lQUP8C6Cv8dMzQspvlA8EVBsv75tjqRZhTIuVndXOptTULRSAgezE1E2g7xYGQMzPzzP8
4JgFFga/2GqJEb59sCk3erH+k8WTL+RnMDTLYatgw4cfta9jwOHOvVqTBAjK3mGFIZd9FoH4pfRB
4KbdJM4DsI+HPSPny40zMRcx8NiHB/FYSoLuTwsQxEQOYp2romAcaGyjKzw2neSUEoBa/g52PDoB
k2k8PrTqTtogBSdFsXD13ixdyGxLDTE13Z5aoQ9vSW/51cntb80lDzxa4kTk4vAfmYshzDWMA41P
hvfHW+XaRA0ZdTtwTagbjkROd/kuo0ERjpChzrpT+kgupPMA17GuCjaj6XjZvBZeELAwWCr1wUgo
pmWYn/dF9E8HiCVbKoJU7J4vrLYeDwHy8nOIt5Xbo5TDfyD1rPBwj6kaaoQYPdoCVfaKKVQl6Hr1
rbfec4d2kHy5REXT0vdQVw8cnif7zxQ9/Mi1mISOiaFV8SqRwZzbpx72gEJAWRS/VV7vDb/QznsU
Ru7TI1ebaPnNmBc8x/yfImhBZa80oF0x7DFajtj8Wg50fQlnZYm+LmqDk2Hkq9arZCHm6EdoXHBz
ynB5emqqUJ8fdm+KLjCw6+tMpP9AaGw3yqsyMLBcmUqghXxOAEefM83k0+i9A4+e4JDuVkIOOglS
VM1G4Qu3WRDUqIbmHQURhF9UjCPaEkZgmfhXQSXNyUBlkYVhhMH3nS/WJMYrKMYkHii1YYXs6NOk
tLQxNmbpbz6ExCN275lnoQjEP/iPQWaDFIPaN40WfW1liwn69NJDbp8XYuIH1T2zxm7fNYLUZNSK
DTeIh3ElwBoTonh/dnxeD2NEnRxcvKnLC9jr2O5OGgzY7GOjScAKzqR6LV295GDOGo612jy/7BDm
RHCaEnk2eesKw8ySOHuohS9SWYBTMRlly7p3XPKepgOJplCUQMjBUP2D5wAG7j0myb6LbmGSe1nm
KXcyaKBTbKkZvyXmBXjry4zysj+BI34wkdPq2uv3nwHLn4Tblpt9OoHSwu1DoctdeGLw4cKnsom0
lhNE/nA4GuiO8PQgCda40HjaR8JI2rLjiy5/ADaQay8FBrUQKl+6F6jfFD18Y4vUYr6NJeDIgamh
xzmsPWJu+u+2rgvbZrhS84cXvy2b+Zq4gYP2VtZWC2wdB2rE7U1DgIJ6Ojp7TW7vKIxGSw4JQW4w
RNL8uSNWXr+Z8GKOmlNUC0hmaRdTtzhgqXOqtq00bTH11acQRGZQpr7JS2fBaFYWoJsTvkpdQp85
Sbg0CwDnEI0p7GFWNsUVS0ypYUQ6rlVCpVbIWGWGcjQr5pvKHYur3A0o2ZeTA1NZm+E0XoPxRlgb
0hkSPqIY+BdHsbaKOr+cSPWsQYMzRLiKVdsF0LVI20NR4126Ougk8NSD39jlKi1RbqlVTqSmDvd4
GrpfnM1ekF1Vg+Xla8fUooaZ/FHZ3qbkN1gR2FPdQTAoMj551DCTuSDfjc3x0IMjaW1kC+cFVTY9
kxpy7Wq9bqGgmWpUkVQrNttGGp3e+mIHzuigvnV198kRO0nGmytN1Ig0y61ru8PyXmT/LyhP7o/I
xjDvVnroUAWXmWI2Ms/KlTDcCB9GcgTdcwS1Nq+mW7AD43ssWSxLRAsOxBITj/k3l3OohIDz180E
4B3GwobFS9s7Fi3CGCfVUIohMYaVPB+BZ0ORt6PPaI0DYMMOw988Uc5yJDpaSowd1lz48rq38Krd
oOLNdjz7SRuiwuDHxLbixje4o4NumTTnOKaSmUneK6OGebom5GcD0lhd6bxielqF3iYGxrIUr2J5
CXqRoSjnldz7EVA22yLINvmGpR/H2TdzO3rtyYWXSZPBKHjEFJdQ7UW5crxSZX5nJnneHTXj5sCG
MxvsTQ8jjEbKub9+aEXAG7cZbfN7IVPROqZYCsV3ttJIoH25ddDrwA0lqRN4cxl1ND9qB/mwytBg
68cql+B/ROW5ATUlfLuBW8D/lp3uHZ/rEKtlmhEhRJnrcdC9gSUNNkF6fx5JNKqxAD1RKaAy3OxA
SM/ajYJ7mF6Q2R5XhwaQDNNVQFQKydX2UtGKk8TpS7se+L9okWicSUulTobBJXEeN5xeIpba0Yxu
oxbaoce2buIuver3yF854oEdSFIqrn4s6ipP8ic1PxBR/r+NyBRAL96EuJTwu4ho5uiutvuJR29K
y8PcKjboOzXdVXMNsvHD/AXNVQUFf40l3VnFwbmUzSAdD/hoauqhcltQ6AILNxWjs71PV2v5W2A2
jyoE92XMEeVBiMAq1xhA5/iRM4tPRx4C43xv5cL9+Q2rfKN6PaE1giaiZq71LNVirEA6MJPXJs4t
j1nc39VEAD6rDij1q3M6ZDdXhCI2U/lNIPhl6OO+k4aKJefqq1mvsncARSkjhAwtxv+6X8RKE193
ybCIJSuyIEZT55nVb9ll4WLFDdcYCFKBQsmMAlK0ObW9heACDeBwRt8b6VC9u4rQBML4KWJajn+s
QwvZSW2lzr43wVyfJ8SnOdBXH5on7GXGEDXycJ5qzecVBpWmrWpPIZ/QPlcVfSvrBJFUf8rgi79F
j69WOB2Fw8yVA9zQAVq1sf5WAvOA3whIvRnmr8LwN4k45LikpQ3HyYliO2sqgusWlmJ75vhg6pm1
+aqnNDSdpKdWypgiflWIkwMJ8UcS1JzuuCyzfpOoDJr1V/NYaAT3QoieJSvkE3HucW67gtR/gsjv
m5cr8+DpUXQd8KbjtiDnrMyPdksh3KNW3ZIGTJ0h4xN8KqzrvLNpSXmuBs5kl2n8xHHIQS+VXnqu
VUmRSwwoVu2Oqc/sEGBEaUyJy8kGTPaIsst/u48RcpsRmzteanVKJlw/tkNEEgVl+ZjX34y5MOYn
yEyKWy1twbkM/XdKwzTVsmh9w8+h/CeC549/rp35VDptBKaa0HmRKKpSDNI7jRczPc+HAn+H3BLJ
gmYhL+quU5L/SfBiB+6V/BlblYVPBr884DYCki9ZNufXCCjXdaiBu473mDto43RGXRwk8rjwfXQM
IBfjbynS4fVDxW2QDiB6KWG/91uiN5pMC4swP+jaxeOxCdpvoGDEXMMKNvbMboVam5utPw2+KFwz
OmohVPModK6+fi1XcWL8fbqyR1WyNoxscW0M5Ya/Tf5wdfX9zDTmjozQJKhcEiQFhRxZP1DtP+Gt
HQxxVGYKUvYzS0B3l3gH5t5dECdEQ4sQiz3lxcHrzFvTbHhtCBSj6H278rYRaFEfkOyRFXQLz7V/
DQPSSQBg2JfQiwMQRTakS94rBCnAaq6sUetrgDAfhA0nhV5NriqoQbOBav+dIdqUpTmWTuRi6veH
epaoM2deGmqypycUOx+2EF2oPiTAO6uhI1a87WaQCsEUdeGky3goweAMElonenlo/p9+toRDtJQF
RPHQLSj+Kwv9ZKA2N0OkIlUZVGUasII84e/IyUcmVimGZQHF3cIBOYjz88JYxOrYccJgMT4j0LoC
nsVnZf/qniCZ157EgF+lFIM5ngh2FeZXT14KYqA/4M190SetjN/unq1t+BO2BFlnECa/xSzsQdtI
3zJDQ2aCQRpJG1/cqobKVmZ4EuFRkPbwx7WDqHaHM15PhyYxkogvTCndPXRBhsRPmdPEVc+Hx4Wc
z4Sp+/6AD0LIK/EuNSxs9bIJfnAm5u0aVsPt2lOoUlgw/HRQmpzPFcM2NvsHbB9WJ6+axodF5tRD
oz0fYaptlmxW6F90zBE19qEMFwPk8N1z7T92GVRcxVvIw94DilpRHvHfKYh+xNbqjrpuVvZ96MIT
H5G7LmWL8m2Qiw1C25Mw/ST6l7kpA4JmWxj//6t9Yrc2Z50vaYD4uRZwHWV7ueS2A570O/vBoGdu
uin/ToaVI27fl9dAgaZmFTRLUWZUyC7LE5699U4WN84AwlTXFIjJOnR+NuSYTWT9zFrvXbvYdFAt
wn28A4Dfe97LQeDDb8xzZBAeqAyt12ipMJ8s5ycJDr/ezH10APyJNd8VpiradNkCmrcgbfk+ceRL
+pExmmgXRrpiEFR0F3z3E+FwzbEUgr1jj3Sn3ninYH4v+yXjT8ovVro00T9NmRqU/0n/7ITJA27d
oY+ssdwjJDWTGkB3TlNj5CtVzfVYzKgK8BUKMzY8ViXuPPsmrTa+pchHZdGixkUMgh06T0EnO2LB
XySzbnyouscegwrHcPdqHQxp8k+yxPMfWnvFOa6ptDFZfaEmObmbfv5Ym99Oz/qhOdL2I9/f7aWi
oVBEOe+BzO88iiGGhv30zLh2N7duq+2CzxGxzUHSNno4wfHRWiMVHDQq2HKg9F0JvuE3TBt2jo7+
xaMxTosgs1+95xLNUXTbm46ng8t4nLo4OjA/w+/IymQ8vzk0B6t38frjoTTi3smJhxVXL4JPymL1
fbqWhqk7eWZuSGQfQ6nCxTPPhhOzZ5awNIwBWNP740bFV+4pQh+K9Y8YqXB9THThtvMbBJQ4uwLg
qPX6RhXUST/i6EXRs0EQHoEii0yE7wicJtBTWDpRinbo0PZo0ywUpJ+vuYKXZDpxCgqNrr4bRal2
z7q/PmxVvVg85O53gjYQkSUJuIPtPMDpuFkenKHhE3CmJJuy7DuRG6aNTLYIZ2tozASB6uM4+xKS
TCtGAejxUsWOHN9V69NLvz7As2C/dPLofZvXC6W/FuAImhk8CDHcKKLeLawnCp9qMyLg0UOw32qB
LCBMl2N2yh0TzCAw7DYLmhC/IH0iDRmGoN2+j4Zk9OuLZrMt/s63hGCxx4BaKYBR6IoxhHkHih9a
OWtydX1mnjtvwbVCyfqTzhzKiZX5B9C50qPKM5sQzV3mkoOjy5ZCyNtJ7zQTVSzeXn1XiOBhkWqu
E1/A7UUAPtmkWxlqTamQvogT3NxIejlL+5wjSVIqlORFtFQvfSKn86Phgzv0uF77WzO4x9YzRLF6
f4J1+ruPHIiTPOCBDY8Ytf9Y4mQovv2DXbFXVmuPYt7cMa1Dvcfc3GqKz3OmLeGPOSBTK7hZe1XF
DVmmUtNSvcWVS+fcUxKUfq/6+TgxmQkB3lIhE94oHenqqd+4R4Cu7tgMSa/hBDZdCdwSZ5nUDUzE
c5qtACIzt79IWpqOg4nL5EfIGH1LOO8a4jVZyeHl8G5jpeT+E+f8MrcT8++SZ6bA6+vfb7dmI6mt
O6aq/OXghwzgMtw5T9jST7XdX8R7KOA34hLsZ27kk0UQu3XkH9LorakUOotYj6NFJME7skvwkhCj
bTXNDH3CTQ1402jQTwLjzpOJCjhLmmQZnqvNz4too2tE4sNDli1yyFofr3sxpEcyhYJjvdVpaWYC
FKe7CSoEgUbsTV//26tCi+OcWo//COtVMi3Shu1Ih+kHt3AK/zw4S+UVyK2jjP3cKxFvoPG0po36
PRPfvFcY9vWHZf0NN3NEobcblphNRRzLwbvjnNSLn4lffVXxXp1xLiap0p8za+OrjURXAi9gk3+C
avn2xGzJ4VbzPQjtzZyLZw4WloqdshW0FaYQ/pBxUrk4Lv7n9WTT25GrbSVW53paqAZ0y2MnWsSk
GlziASUvr/KDEuLXW0NE4swqw+eiTmFzXs0GN+4vP9aJirQAx0Ry/d8QZkqQb0jMhgMqble8ZIdt
uO97qu5A2SPijXa57QdpONlB9dbVMXydr1e1J5L7gCJ3HqWF2+FoU2DJPOkIyA0AoYhEILRnIW+B
lm7E9zv9Mr7YiddWDtdXV02QZGU5R1HOnVBkgN5XG6Vs6rYerctNYZSM8q9queqewF7Kdw+/IF5M
KbrHT+hnKZcDU8QLJRTwK9j+wcrJGftpJHKxW6YQrmwelHjSIxyf/kfSRWu0/XSCRBsLpTs75MeY
5qj6qxLLLp6S/L9ulQaXVBNp9DtO7jqWR2QWK4WAbJmh0KnmZHQkBRd++OC5Zc+YAqw2xqJ3hOpv
wJMm0+ITogtQPOb2kUCmFr4o08Fv2Tulh44gM6UA5prauRUxf/IOdN7btfqb2CgkmE+LBjbftuEn
2A6/agRKo2wwdcXO4mjGKVf4SLFPCSgC0A1q0zHN3KUg8XcxD3QxDCzfcCJ7/GINDF+99EC4cWRB
gvDs0PVFlKg1SQSknjriPCq740XIH5LF140ASNioyw2EOcsr6Hi9JP3ANs8CcML5xgoWyyHmbnHd
BnNVd5QGdb4+Eu5sHrv30zlVXFIPoRARA1f0UbwMqy/TjOfbN/xK+gH7a3lC3BFyJYyAFko5p4M5
x/9PsaR+oCSg1hvodmLkBgDHDwxrr8zXmjOdJ5u8q2KXQs/U30lnv61iIm60YTwFkXZICA0xjISQ
kOs/qfqfQplGlikitHR53pHw0J/8jOdOusQ+ooKkVpKfeoeQtzj6oDN0cs/7VqG+GO3PeZtYi4J2
QxFVP2JW104+RQW0961waSBHZpaHkPr7aDG3U3OOpqEcLB4MSqzy1oNCgr/oZYQA8SXdOGWfCMEQ
MQK1idD136USCLBCqjpFpARmnqz4wHuIS6oPtH6QDhuBe3RGEKvZcnxCWMulRvK+GDa0H7mf76J1
9Vj8ZLVvvkw+3bqyDqHyzv+0jNlWKo/upN2LEwnVS6IJeC+hY9/w/dSFfmzJgIjLk3L2zOH6jpnb
fIKICfETGArzBSuxxZba6kc6QuFiZIVzFM8hLHCY6Fc4bNDnEKl/9SEasOhihUFARqlxcrJ4+GPu
zfALL16mS5p1bnl0U3RUfjcbbbs6KCquad19V1TnhJwHc00FQ8Gp6g6vVZsQqwhpN2HZ/KFSJuC3
cyHxkSfmbPYZv9PjA1v9Ewh1SJnIzxqG5++frTxZpdQMqJY9WKZg/Blrm49iUdeOzjlZLas6GR9B
ns6XL/R4BulRJeL6oGS0EaSRUwEW5Ndk2koAB2v2XA8urvka4YUoTwjmMuhfGyD6uaDMUV5chRRJ
PiSpOZ7SjAy03HmcDwdKf8TuBnbAoXibPbD24xSnASt4lPxc8FtV++tPn65i+tzs1TcmF9DpKOCK
pB7AZ7k/1HyQR8RM0kfo6n13ip92jyrJ2kikU1oxF+9pRwLhH/ZjxQv7EyJXjvuXlHI85y8MKwpf
+WyBqpSxl/V3EZUFpQWN2M2okAoROl8pCiMVimfG0t+l+R25NxBn4aA8bYrN2HExiNXs8T2RQsUW
MId7dHqv5qLeev6G25z+NvE5E8PGLOGOlihMQcVVnUiWqDBqYtm3KcUMPcIVbg9aVEbVdLPBwUIE
6Q1AT/mRrKOmPq0Dcs0jTpG9n+93BTt8s6rYzTUM2zhWxFBytrjiyRrlQpiIJIdbJsq+x1cWVdvG
ahoiPRrQAzg46SnEM7WQ8eXTI7+coC6DZiDs8ChPhU/p2P0Gzr/LnJzNsuS5IYExQzBorVC+OoUJ
/GSEZKea4VUovg2o14kNZGZYEthBwmeoWS7t/3rOunEvC2g7ZEqKqCtsbi75iH7KdB/cOV40gjPc
0MTOQQIUJ33L6/SkPD7GwxwauLtgtyAXW8mAhG7nQhsEdCRfmgVPQacGIJmpN3bGpd4fNHAj5/+W
eXnFjj0J39xSGha6o6DHkHCfI4CaPl+Hb9aiYYYMAqw6Jd/apj/VvmIaAxtQqJZIPFYs/HcyGtGA
voydsbNW/qywz5WV8MsMMRXiE/eDQ0Rj/8S2Kmyzl5S3MeEmwoxpXvgUOMpR3UoE9lSx8il8YD+L
3swDTRV00tvMxUURhYf9EOV0gtKtyRM19CwPbolGFUHPYMn8shmDxQtvdSS/iKrXuf/HNgA+/TpK
I203XAmFhIcgq7K/klghPjUhgSSR9jINOXFXTcALC985uCoOQVcOmGInJVb1jHaGApHtPvKWZeGM
vXVkgWyVXH/rgFbyqkjHl7r1FSr3X3GDBBp9Tu6ixP1fN6OjCCamDrrwwnYqQSUp6PY+U1ZjYptR
J1K5po4/H3R7q+UjTh+ri0fvyLg+2W4Cz2PM2hFroK5kC8LEkb44mU73Yy50sJt//oDe5SseELwF
aeNPdCNMI2xugS8EQ7uUXBXVK6ofbCcCUmrwKgDMo/9pUfdIyMlaT2H9gW85JzXkhtj42iVQHeGN
+0EzHSBqzLrEApW4GGphTmcFg//cy3miKGHfmlmkVlapO6yBWkJEza5qVr4JyYzIL4/2s0o0iDuY
j1RiS9GLgbMRt3ktq9ODvV45fx+CWxSclBBXq9Ao3COdXhv8qxAgb3rqC7V3APcDKiF+0PfxC1Ku
QaMkBWF9GtlKax2OUvppEhIMz7W4UGrqRFQ7Mk8SIz00AFEMPNSL65DRn1M7ipui+1hb1k72M7RJ
S7gnGKeYT+OAaAGpwfE2rFoGkezYOFVpgyAG8D5Va1YAfU3RQb7UAPfHnTG97uLtGrt71e6B4ewD
bImNEZdju5ozILGMYvma00ubK2QIzXMAXh1skIhmnbX5p6jnk9DxtULvFVkznI/Uo0LdGH38vKJN
Ojvziim90SgQWdbkAgK8SC9bZeMJ2SbkN3vf3nMA2/HL+VB05TJaeJLA8Q9v6aHvzXYVmVdDsdr4
1HNYHeb8LrKvHP77zFJW+6bKZcmpdPZ/DT216tkOv4Q7jY7cYT/DXVxRMBY7ZO13Q5qOCWwG/r0I
tLtBgjdSTg87LmgOxxWrcYRYy/1fI2SyQ9oD7g+YGt0zUQWWtsaVWGg2j789qOR3ldx1tM7TaA6S
j8B0plaGt+F5pDtht9zROS1eRZY4mZhzXs5aFna4k8iH1FlBR7+dxKflyHdNjSdBECkPjNyvDe/F
oVoEyIit2fVaHQszGaVu+4n0uF9ahATtWBlW3EzfbUgK+IqZSKei0o6uf7NlHYiBQ0ZCEuJ8sXzp
nBRg+Kv1vDI4nk+E7zjYWal8SF31If4/nWz2pigJXVKVLbxx1rVEKtoKm+Ej60vUIqvvuIZU0oRT
vZw+4njnSpq8jWw/V0Uo71ZzCMR4ccTWhA4hwWUjAzBP/JVNYL2tpm1n3PJF7e+LKHR0MxR0Tz/B
E4kaA9by3ya0s3QRhVQboTX8nEcsiWw5i1rLYGnpkwDMcTh7oIcQbPFrplDEegGGN0v3A8nELdke
u80P+YHjNiRs+gFUr8FnkUO/AiD3Wpml/4sSOcY+IkP1PiVlFmLKQaqyZHI1/BM/pFz8oh0NNx1t
jH4fSx0vPnBDiMnLz0Aou27tY6mclQkyUQIYlgrjzw0omqOe4O9ZOZmD/Q9rMdlAj9wNxNmqqKZW
9F7eAWM5pja/ohmVorTY9EKnlG8hRdScyEWtwZeflz5wl+ycmThEc6HphvkXhq0s5NodkqR8WgCK
kuotn3nWzC0Aw6MFeaB0brrHLIneK2bgu4/gmJ++rGmICacC6UQGWGgazB/QQzdCgSywhbqq11FO
vXdfAPl8BOmoBtXosak6zpu/RJck4FKvjMECVZ3D6PWzmz2QpQ08M/FqQ7qu/vjpPzmBCvuKcNyf
1gVmjckNc/2erbQAX3KVbzXfPdcFrwkTCXNR/gm+Sn0JkIAuDN3W3FE9PahaJdvbZ0adgl3cGDhs
5xLZplZlxj64STpHY+NbqGnbMr+3/7ETfoqnepmOpvQ2K9He+Lf1/AvAESCOoanClokcY89qJ7L+
BrQEIeNL6reRlVUDLqEwgZ5Pl0IR7wq+EApmJqs5IAU5Uro58WN+sBGGF5qHfhP+GWhEMkQXCOac
ATPu67rxWtqRo1zd/1U/5tkl5caG4+OGgfnhT8szcAutbWE8MX/Tw5SVEj32qGGE8zVVBfXyGPY8
ZoulGyf5yflPDa7bUmGDF9i/otlQisLI8V4Tyt6KkjHHH6QuhwJBPZKlGk/fOq0IbWBXC0zUrxE8
/Ni9xDqSE4IC3rfWOdqEYsrNaeLXz2fpRoclBsXLrNbAfgidFpp5zCGGRSgZ9UutQaPb0zw668Yz
2wbqxX05q6nWbTCigesQQJm1ePmAWtOEJZMxDR7F+oVI9eYMSghttXTiIpFva/KBhTNLwED+mbAh
TYzjAMDQffH1GuFcF3uNwIDz6BbZKRppBwD0eL2Fvai/csW/AVdIYo07AKKaeXnhcSm70rpuSCdC
H5ByGjOKTr5XOlWfpmrYCqDmjeJOjyppCzDMbzJL06FtOzX3qoyi+Xr2fMfiv7nOB6wCtnxW8euq
Y0N6Sy9dnXlSHmZ3xGR5SrZpzPuYpKqHoiGdo3eDLg0NBI7o5iny57n4stNcyOXZMdl3kJAy4rqr
+ds29+YwGmKogPnZo3ooicbo2MrVB+limn29iaeR8t31DPzRFtcYPg23+nZPm96XkcVI0Buyk4/L
+nE77ai9flbZENKExOr5VZA1vqMXys7eP4NCWhg0xwp686maa4XjVq4XCjowyvIU66/9DzgNOprP
J68B2sdGkRUWmJebyEz8HfbD8G6251iLSzyny5tMzIi+/nUcgw0QUmX59SiQ22D38a2sCBbRmsnc
H1Qhu/L86srSdyjiMOL6fCbHcJPsh4plJMaWdvWcyHrU8Afjm7EMu6QTRFMjocBYAKy8SO20sfh4
eAsPngefw4ifco3EiZsVDU7+B9aMtOvwJQI41p49oX+qiOr2UGhmEckcK8JK0Q4KVfcSVSAjA5Pa
uURULEJnlu91bCYq5R/fy6D17XCsIUFKZgjnHGha31XAwYIwnqzWtrGQzxybSDRmER4xgpdHsYRZ
36npjFZxV6I57WwWvwxHQioczfMxcgEKHxubMr2VzOufe31pw0tUNBpL+5UyE0S1vrj0j7VVVJwX
0Iq/hhJNBAGIvuM0ICq2JLUXu6m9IRY6qeVvVdUmM4nYJ45IZBKb61FIVUYTPSKX0TWE/q4VmicH
KJB5gKa26BaWCBq+xF51wUmuagmxfq5J8tDIHPrY+kmHccFGPBw1z0XQZ/GERKfImzeKfeRh9Anf
gacl/bgdc2RMBpUsThLKW4Emqst05RtCwjx7Dav4FNweLct0y5zXPIK8091ig7WSPkWctS27NMBS
sDx/xZxcjCUlfofLb63JUOCQ7EGyszGCMpMuq4PEls8v5WvusB6jOg1yoRGhHOpEDEoZ19Go9J3N
evU4WHvkEIw7GLvzPt5mHCTQIpupVqSyZa7JvUIRM6fZAuXwLH30WRVHKesgXeG4JU90KuKfIlUj
dO76rQF4Z3NdDD+kJJCUyvoOgprBoiQKLEjS0LCci2+53sr71wS9SXBWXNkLJyW4tTIUdaVNZ3pb
+vtHWNUJDkbkc6f+rh29cmA/m8YjuaSxNRBVvYEmRvVB7kkDV4GmhUf23jSSFrO4PaDG1/c0funZ
LXLkx9vtGqmF5u8ZRfqzxR0R1mk+Xx2KooUii6htV5hyLorfAg6GUjsH/JfUAh1zY4YXby1pE+2I
7ulMUFdb7+TEs6vU5blXDLbU/lKfnypn7eb/wuHMVkEgVSqGfTE8o83iDLy+zcbsFEnO4IrH8j+2
Eypv+cRcg+bTMZ26StTHZElMORzYDsrJBQrYFEKc+p8T/Mxw6pArReaDAGQzpdyiuPCWgp0umADY
nlT+TyOXClpVzpdoRxRlht/2m1G/AjyRO1qkYInU7KJLmC5UaYU3qhgUUJ136CT6H87HC5qSt2vH
WQ9PXEubZsvuXCYHDfoFWn9dPsPlEkBI22Sad1uPdkSa85yGz1WIggc1tub76lukdJiMKr8steuH
hTg3+HerF1LyiUz1oQOPtj6uSKovzNw1jWphXC7n7WGQW8M55g0SKKWw8SK9bpCPM2X0iKBfRZGl
MmHAptNS+KaMkDiSz6W8MFMq2W3IvG33vV0OOnJSojSPszzEvMvzmk+JQ3bmWSV5XYg9dSt0QYy3
vR0V8TjSPLVVpvc1+Z4KgWrkdv4eMfaT01c4T867SGlT5cxDv4SPmx8x2aBT3e67Dg39Eq1h67Bz
V0WhA1LDIBnXFxHRbzN5iy6AQabtJDr3KnoRT3JIRIfon2Bpf5FPy26ojaZhhmigg99XiDmTsWFw
U1Km5AhZEUg7bc9AAngq2N7D2nue6z0Ipzmu5MAMDahqqhur07BZHTy1WhCleL9tjCyoa/yXbecb
FMVkM1dznEKcmBQ2CXSnQ6Re6XG7H9HSzZVxl8BMZNJnZ3tfhQQOy7YJ4L1Dx+m/hBbGQhtVUglE
ZcjCwO9H5c/O3hnafXmAZoZ7Q6yQ+gwJYSecYPFh4aU0FmK08YDUv8+q5/aKVdYtmZSHNoHdpAav
Q5WC1LC2ulYgSwQ9vPPydl14RXvLwXUOeD4XNDSdHtyDGRZuifWB6lpbbun0ka2Se+pr9G9k6lWb
AZeaELjx49uGl5SfeZAo1sq+fvR23RxfH3baPF7TCXzvCJac/pPn5L0n+HNybzlF/hnk7La6p85N
KeNSOTde05E2nfrbA5KTJz9mFevSXqNmRSWzWAIg0FB+5Jp/K9zAPnNJvOSYbjZhBO7xBd3G8paI
Bs6EoCtoUw6B48Yua9oR5GciG3YbNt0cYqWCkSiZUY4xxj+3sWlkWs9D4Q5BhyLyiWzraYWeAEVV
87jPCa6m/zC3euEliiFiPn6kAMNB8Wlvh3qJNzru/0YwAaDrEz29xwzaFuPgG4QrP9Knr8Ratrjh
OnU5RyDnUs5ztz6WRzcG6SXIE9DearR3f1b9w0PqSZaBZNBnGaGRjORLwp6Vpb9aV6Nei6xc7Lw0
/XyzCg3EowquM9/IcAnhVX29BnTRo6mgN11i4zEo0xSM8dAimuXk0G+MM+wfoiTqPrL6m6SimWmE
n3gM4VMnsjqI/L2MAGnh+bDV0vQnNN96aB0xy9YsbggTjNuPKZe0m4icBdM/6lcjeHWN6rMbL+SH
fWtW1H6g5GXi9Sy/h489EUlOpiExPs2+zEhh++JDxryhiSR1FG4fncrXiz89o958Mw+dO1PTisyr
C7/ZO/HVWAma/NiFo4Z+LIBls2MymmRIUdcRU3WNg51OYaluVEneq7zcJrUgn3fZRjbEr//tz+jQ
uuxEYoYkYaYXWzWE1Pnl1CUUF2R2mcv6u51ix4W3kfROtgiLNfIs6BcCJ65Aa201elu9t8HZhKMo
YPmAWUDCm2K9Wi57DwZLu8GHqjvUDNVIgzdg60BXicYvsL1BCLYee3/8pdPuaeWRAbc654HNy4Y3
4JkxjlLSGftYgrOTX89qmr5uDUHVlR7zlWIA6lzWTvgp1OSsDIv1i4mpyVG9JkNGXqBiwFZy1Y5f
VxCKhfuzy4fa9Ak9PR6onVUMv5c+6FB11o5dyL5huNKlnbY8Eeify4gzyX4JLCCFsELwePWguBvO
x2ctxNm+oHAueenr2Y6LI+6ZpSkAczr97LcwdTRRXm/nU29JIh2/JpjtCYuAze8mK8KwFiJHC+4y
h5whGU1MUJHtBaqTuWMpmo59nhnOFhjoc5hJXSyIUo7XPr30d360ZPBBy92FUsMpT63AUhzqUXh9
CaVt7HzWixy/b2GMhpXEvttIGTMSFBieycJbRtv7vfPvT12cQnE+bWlIY5ICoV/e6GT1tt/yaEyB
73cITlwOtXriykUqLoFGcawEPVHMP2zZ/x8hAVAVqFOrGrGkVHSnT4sWsS8O328Hsuxi/myCJAQB
ud4zqUWbxT70sJnyns1AxE8A9ubbtJiGVi586r9S5l9H4yhefzG647++9zLf+Vx0tfGyRVPyD8BS
wzuXSvG6X7kHfytERniMJlR8m8caL7N2LxGrMvzaZ7wPiG6i30KbuKu9jb4Bv4Qik+ZekmLN1IXe
aWBHCWzm4W1geWOWGB0+IqgTyPcuM5KJCiNcQRb8+PklSIu3m6f6Wd0cEIp+WNeM+Par3YLEE5UM
qAdb7OCKxZJamfWOwIWgk876rPRuPT/ia9XGEngTJ0TLmiLoTXjU92xvqQw7ua3Vqiqv+liE48GI
myyDaX61bhqFUSnemCTSRvIOzJrUrCOmFYG6suDzBBiA/2Vkwf+PuvMpCyViSCFuRC3i8/84+sCu
ablFpPHHjPLYafyQAZ3fiN3KY19DNDExGhPHjht6QlAIkP9kyvuUwAkk9j7ulVbXtGfETZsF4mR+
uVeQQ3xomW/LZlPdj+kRvcLC9pZjfvMs2IMx19X9e0hPwygXtX9iFpthY8XNkt5nQvH5LfEeSRTp
d6p7lxWIjbUzWXmp1RqH/2cFb1Br0954fdU/XquBD8i8qk3rWTQ2b28gkmtfrTUXgxvLCYoQiXX+
4enfXt5BZAuPRYVGb5fWimIpYgpZ2GU7bJO8l+ax6gJq4A4Lv7CAWEENKiOMrFinsFc26VKl6OL+
gbPKMcwfD0zKQJuj0omHIV7BySxr98ZK7syjx2vJ51Yv6OwfZYfX9AbW8lA8FpFviV7WitJsOv7c
QR4VuovhrZgLFGE5DtQTlg1Q7Bs56C9fKPbCaQNF5qe14NiN7OkaLyivJu1DGVF+cENIrMGDx4ce
+WHRwyMY1bd8kTi58gCgrJIl7PJp6phxn8LEbm151tQutJVKuI09pxaIxXQo0EeTuCY2LuMT/2G4
2D/yc4gjuG/ZFLr8F+Tpm1nV7OuQyj3RLTE+5S2zjYrLgl72d7pgygp2wFu7/oN5NWZDRiKC3DOu
MHqqmS+1AeHhOEXzoA6c+XR/oENpICbIoZutWQeYNBOrB5SgVGv4zK5HlIFCwDZAsiYdrGy45+U0
aCI1eKQCquF6C+LRuUSshA8bGXcyArSIP/zpHWyQUKyBg6s13jvWkONNyeHUaZQJovtpbfMvlVMb
+DcGEtaDzW6eElsbzZXfoHneOgmieRcupdMs/uhkNX0nsunp/rycgTxu/XQdOyKk0BYWWfWF8D/K
IChIAix0hN2UM3boLFH5Cv+QGz5Xq/VmmUKhHQf05Q+JLPTpUhxmdFu4FN2QzJO7aRuMhGqdYwkW
WrcGU2eNuvGs3LVQzCNnxOOkAFBNuioWqNOkgksCwxsOPU1yu1LBKy5l3iR+1m2/o9Uj7PvHwped
n4mS3Wl+Pk0reXYKzA1IRhdXY4xBrLJbZzHko81i2lr2Gm8yPqORL8zyyI7Uq4wiv2FYSK9Bi8nN
BLhnV+on7JXPGKNtBjMTWxtTaJ26U5QelY8M27RxxlZr6YTL4dpwEKula7xUtPZwPBd/LQJ6OdCz
uPjvSbL7PhWftqP9Tl/S7TGAMQ7tZS4Up2fzSIB+nCS7s1J9wWwnrmPhOmopA/8KoH3wD9ybyH81
fBTvKZOjQtFVL6CNyeaYdZvLJyOFhodn/JD8cG6zhvDdi/bhIKn3NWV7cN1bWXn6P3CKc7S4MIDW
5mJ8kO25ZIIeowO0PfJp3k/uW3Avst5tI/ggJnpyvsIiqGDTBD6HGmCWNHoH6whaQy/H8NI43dK3
BPF/WJ7TVeLhScm4ShAIoLzhoS9DtsCG8BZPDLK+UhnJuBxnwvaAw41WtaPm5Gi2jEUHINL8KozQ
DtolmIBSjzDrYDW4zbdW8q7f5S4ctn0KU5PiJYZQZTHnirKa8KMUelY1fzJcMl/pEKep3ripeF62
3rbnHD1Xo344qukGYUF7FvSgVhknKgueIGHrfqahVWYraNjQdslp+VIOtXst5wiQ5eaiVMgrq7w/
eeVjfTSAA0QfMNa2ozIR8oRPnznbCLlgBmwaOYmhWjwVa3OcKfSCtkBG+xpj9izYL9YEPyo+2OcG
iRIAiheQ/7KL2rMK7dH5ZZhSgklhOSGOdgoI18nqlEvnq9onrTOVDI4CEY2zLcXhjPYbh1GaMJF+
WRAEjhZ0fzI3c35fo8H0Md2U4uVqwasUtluBLzmfU0bPjZy5YgMviW27jHWWqnizdjG+oPMlNGOn
6GO+VCyZ4Cn0NGJSZ+7p82tzDgLnbnk+qPo5ztRSet1PJgmld9sRNwgm/mzeTZqQY5Dpu1QqhW15
omgzLOrChfKXbUNdlKZrjPQYhDkylm8q4AYWkV0c1Ed6ezzhBLY0hwy9V8pGLA2i6udxB0UPmmbr
0VS7T/7kf+LBz0JPW7icrUxQxCJvaZTbTmDK8kGYDpyFr8XRMl1eL7SnZu8kmaj7Nz/VJ5UIAnr1
gDLBpBYkZu8b1B7j0okOYfzHREnPATitHcblSMXrlqcPV/neRhQpSMS2jxfdqnXc+Y1mi+pQpcxI
VfjSpZjyreS4GghR7W/eHoU8Hg5UxglXsLWBj2UOcxMFfb6JEFCNS5Dv4v7SsrrgGBfDtOGApTMy
GzO6kkfhPiFeXXtUf++TKvDzJ9RPyc/KmOj32blwE8uCPGp8FV0MviI3A7ThX/hbjLHdZYNlvIyd
m7CJxg9pHiPaVqa8FhLwIS+VAnbnLFb7TFmg0KF+m0Khg2Ky3VfheEIE76sLTc9ykFwzrnZyeN7p
GjqAGhkQ/zSre3InfYRTZY2ZscFrohUc+PZqdIiYXS1HBHqcrg47+GC/klOLO81tJeSVW2R08Lp8
l4FNL5wFDKshD1xxvmFQ8eaS/Lt0GYugIZpCYw3fAZJI0e1YL4F82lXLQZ4nzYDJe2yv51eBfWp9
rPremBgQKFKJ3Ui0Hlr9oFP7oMi+rN156KepWpXf1Cjk+uUhKFuO2L5Xft9uS2lBpUct36K+M7eG
cqrPxThWQazvjnO+oy5zosXOtMr1MJr8/a9JrFcIoPdCDJT1jHzOYJmbOpmq3SoUVPKOeFOiFfVe
kkW+7pvcoEutWq2eKQdIXApSN4CGdlDU6NRgSBm+7BbvNV7cL/0AxdhiYfJ9A7MAWjmSsRRR+NV3
Ix0hdA8PDFdWfBbAeMXiYs6NB58xXJpk13G6+/zcqP1W8aFSjXBD+H9HfJKzrgTMPSFYKq4dQGxK
90BoUomTBRBsv8rz8LAizQvkVBikfzlbJ3EPGHQPxVz45s4hxr8SnSUFCJ3GtmzddzUT8TS8blCo
bmC/QjcGHQOVcV2inIfIJHpXy94tjAH3CSvRAS4T4GQaPx4BBNHJqlUWtaJb1SX2nRau7bOH7tdP
ki8YjwcxD6MucvraLjW5AMBOY4NLztKSLIBMHIs//EDaMTyXf2dXUHIcRkEvbzyNPMGeKQQ/LeIh
mbOv+m7GLB+ZfXQij37tqXgfFZGFYle/NR1lJ3raT8U2R3WdaQV+DEI1DasxaBL87pUfh3HJ3cvz
zfRoDvoSfX7+XyOKsGNMM26tdr+Dq+UdbLRoSqQeUYlNJ9sjD61dIoTp9QEx4T3nPCRz/9uM6sLX
Jg6dPSwi0LVHhmg49tD1nKhkm24LfnuWoxTWZtkCOLLXlR9LsXG+hOaoy/PXez9qz4Tibk7xdl4s
XcC60ogLMJZeUz+b7Gwj+9J8I5bHTmTBDxncipDmUclKRiLmw8gYCHj1Fbluw7ZLZPTpX8K4U2Js
NkMSSxdAsgbvwj29GbojuiHvakWILhtJvuPliMJc36g0yMfGZiBEohTwReiUUoRFKOqjShO6TA2b
C7FVGw7IFUwvha/BDvqxYRSfD37J2w83MHkV6cGKueypS6C1Bq5yW6Is2hggB4kX5HWYWsSeoMFo
M1sMuFXloMBCH/pDK1Bj42d+vNsi6wstT9mbjrutAbAEbwvH619o46GnDfaaCZYccPsLlPWeMvTH
r39qcMI/nI0CQypFBm1di7SfUxpzFCTTBPijiq+xa/FaRcAalQE7C5+yDQ3I9QBTrGxBm/d5zdp2
ZIFUizIVsiBWvByvAeNrJ4w/hsMbsMCOOe3R2GTiKb33m0rhTmT+OVDUKiK3FK32VOd4A5IBic32
bnt/+xxf4FHleruNJeYsJOr94/WIXvdrb5tW0OE79hQ8Sfaop/Rl9f6sEwJaiE36xx6qrrrwRs6y
JBwo7ru4qYgsJ+bhK1SZjdT3UP2cUjp9xtDw5Cn2cHQC4jXFSjOC0wy7nS/gd64AWpPUW2OIFm8p
LrwRcq78upq0OutIRecQD7f7f3NpnPRD1uN4XZ20q+6+I1Y6DY3l8swM3w/6DROdvr37mAz2IHuk
YBMFlBtNge7xT+fiaCEoN0+YL33VmMCOJGxprikVb1lTg5OniSscwNq/GL7lIDOvVtrr/iGC+ugV
3kl63spAz0TO4o2C8E2/QXQntmNXT1595gM2iHKzAi9KIYsiJCOeePCT/aJ8Bz5UjRUvIaUJDh9/
zvowDXiRb1OP5UgAfuD9XWN7HoFEcpF18Iflr2PRJ/bGvuwsp7DZq7Cf3imwKHl1V7ZdHvO5adDg
xenIKYGUhibkYvEm5ofoWf9mYI6FEoYrVCvMqd1oELy0bVQ0ka4BFaND9C/R1K4WdisFSGgJdpaJ
qrykTB8NJXjzIpEtVIFFRB3Vy4YeRBvat2XZPdN6xsuwylxkLgv8BbgvvUJrh2VZ/rUaL/yYYL0p
KaKtNZdbJf/Mn0Nde/X9PSDvbDixznVqyvd91/ekq8kyOFedURRZCFDlg9FD3UqVaywvT07txP1M
ROm7dZZsURb9J1B6CinPF3tA9g+5i7fq31bHgEL9CmokY7g5hQX/F5ZH/UYsGNxUNkEYRlrEzgDR
GcQy4495a5NhF7m7Yn2bYIuYBa9iJ3uOqOP8Jlo0d9Lx8saFwYP734HIJ/xbva7fIEViMw/xepcS
178wRentzjzUj8yoqGaITfkG0F+qNFXEH9MFA1feeIx4NQkgf/fZu/vYrylUxbM4S1qOFVCyZbjs
B5IOWIOqEuzi//19Hdko3qsN89kd76J4R2kj+HfqlA5XQLucXVEScsVImK+YdP0hEu73C1JPCbk5
Q7jPgg2Es5cTdfP5ArbeA60oEvTkDhjXYInpAQIA1BBetSYo3sI+kcyD0tSuAu5AE3bgIsMBreLI
FHWqAZg2zI6rjBIcTTn+2/F2PdwOS8tpSxYiVGhDSq3PFaQnnQjWcd/mwG8UtSCndQQoeJ7kSuul
nVVfbVPZzBTca++QsQdQBbOOHev/obiXvntiv25NgK2ODzMJsfIftrCaA807yqeX9MLq84PAL2Fg
hcqjB18g20oDpyJXOP/urhvZz6J4E3TBfCHevzjRjdaQ+QG0At58h56EIgJfTWwcDEcW/VHMi6KG
Sg31eHYCMlVG5j3Ysr22WhavKcQyT1i9fAWXEoxoF2vB9i7cxbKil/GuPuCtxSeFAYXdQoRq9teF
HJgw4byRSgxjKqhHbBT5qDbvkEYX5VzKCXd3X+5p12tES0ukIY8WQ45WnP+ppvQVJ+lv8+rFKFwJ
xs26JNskwOFIynQwYjaJxyATq6MHXQQKSDetQtHOWQqgxXn6KFuSgpPNDoVizbK6GY+tFjxkONsm
MV2ASuSJdeDyRF0axiZcVLbuF0NghmTGiliyA9JAm4E54nfuhCdnPc5G39K5vRU6/0ruBBHUmHv1
+Y4zK7MYl/5ggTIVvWe+1DiVaMbjWITXMuVrg/NBzi0QiNu/r7HyIqjsEKW4o3npnZIPs4IYNHE1
PbjPhXUidj0ZaPqiqgMwwrvqEWSP+yponDEarT7bTLG5162slgB2DAw9qXkrQAWUFsk/UZa+lBEH
WEi4YX4Rh44WdJrt/0yys5JqH0R2DT4fMpXmxbjora8XBW0D2nh2SBE3+Pd6vgZEVY2WCBRRC6d+
h6CGoBBsMApblFvFMBJ/6HpBhLYbMYGC+BDOry/xdRVSwkcQbSUhQX/WTZj8tn/WYlkAhm3QOwAe
M/8j1WDqICoj1L613rYySdEumLLLrGxZiqGcV7xcdlASK9Cr3a35FCUDDvTywT3xzhPkVK3mKl/w
+QFdXQITYtLXa+w6obkrS5rY+OtCKnP27EtKmWjynPQhFSG9o6pV01k9sbMA+5PrfoWVs0pAZZ3K
ljKbiS8vctZrzLV9D2pt5n7b5VI5T8DuS+U4VB59K7GlM9mtrkc1LSKfblxxsOeOJq/nfzjQWsit
wQNLKlFWKv9bSZPl1696WuzsnIoKCvd5wv2KZqoxUvf32lLrtVfbXjAbIPrhQpakOughR2Cpkbfo
d5vFa4ogpqZVmHWXdUUuieh2lu07vP82yCuP7q54TGZvbfAgkVy0sgmPxdr+r6DMAAyHAkl84mka
mhznrkQvtThdsI8G0iT0VN0lROGNRt0BnLLLwFxf9TkAe8lOjEDfbAI1AQhrNOlAPDGaR589UZpF
VKJKp32Y7QeO/Yly7x4mQec0YLQ0iYeJwnkAnWGX4OCBp1qV97HSnctAaCRiOg0Ngb8hKPVa81C3
caNoP9sxA3RC6PSH8QOSMze+hIblEc5ToO4EWUwJUm8jlfaHGh8EN+Yjz6MEnC/gYjUmAI8iBXlV
a5s2YIqi4ZY7ew/WSm5AjLX+kNrXuQy42lmBCs+Y8WrCaxV6FsNI9nKv45aVal3b11siPl2qPTKb
aExmHnBq+1QRrRVkJw9g/3xK/eUP1Xva8TOfr0KIDC2k0GWM9Dp75wQ9BvLgfRAfx4y6Yo9f/Ypf
C6ImzOFHual8iYku9gQqjwUFK9S5Gz4lvU7+SrF3fGPYgVZe3Q6ct41K/lHnT0haKWxrO6+8KuWE
gPoIIc8SlWPSKcv0bxhn67PnEmONbLY2WLxhXuzSm7sekWdZgzZ/X2MlO/w2dDkbkTgOZPTrymWJ
xXaFLey4E74DJd3SECSfFJvBSj65cQkRmB7WP3zMPYBF+pRkQGLAMKbzzgnLSoiaA8JdSQBFvy5x
ZQ1mQ08Oq2qvYzFSP7TOyxUhorGPbw/iNQ8q4o1luvtmJRwpZ1W78nwv4Ccwwfjy/3R8enZ/OxY+
8WkkWI/ERr3dte+kt9G5v7vRpQF02BO4oXwfw5/Yz0+NzB9Wlxqykmt3E1DxBvDgMYybzj4icsXq
iuhahjIl9d4tfXLebRB1Z4/qp+syEvmmq0HAw8HomF8vB99D6Cv0xjV4w1bV/FsaIJ7/UJcSMFEd
/0rr87vsRmWggVqPue9X7lPkKrnqq4p33a1wwo/20dJ4D5r1mmDH65GPJOzKYlEnqGAEcOaZHRJC
gUbYCaDz0YyrJE03QrBCMSbP5H1plbl4lWRfRRn3eeGwZBxGfOgFJeObkbwRDW0s5pBAmWfu0qmK
BQyJvAXygTNeTEvao37lr3SfG19ph28WEtOoDAPVxvVmJoG9Hp68v+ZsVhiXNQ5LII3ZRRJe0MQb
zcOwunv3f4jnMkoM93BHbpIMdr82KjluCZDlyfUgDdzOm0jdcgKDrWTOO09jeCxGzEShd2vHXl/o
XHixtzxhV/EaqDCABDMy2lnVC5yszCFBGVrThX/O440wPVblHvF1W/lhvWDrm3hrLKYi6XYS71wZ
EHWDxrdOZfDmqC0o21QXKzu6pJ7TtVZCk2X64BTFW6nqMpSYvXNmExaOtPIBpF8z/CEZZihA8HcY
pnggKtSeDEnQNvh4fmdYUX16nmnApS91ATaJQze/sWUCX9G+rGsUtwb3OAJP9w9TAvGW3Uyzmzww
hhiiNS4EUa2zY0PkEocjbwFdJqHDUOiREL/A5RZ6xlFCoGtdKvLISoVweuTRTTbEOFzJFcD9UeSZ
hMJYCCUsnZRUNjVyyL6PwrpUt1j4Gv8xh0bT2zEP4TrSLT7uG0ormWpvqq610cDNMdG3k8pRu/ON
7YQqvAKO+1o9tuzuLkHNdR+PXaic5WqdH3wkA89v3RnThaPDcxo3UMO1KA53tFvBTalRRCnu+kfx
ZwQK+n+gQF3btEERZxDonX6orwOiAZlRxYvceMEMS0b5PnATVKaVZaWkMd6FYUjNESwO2qC5w79K
smuSetzQrZD/2LDuwv4AyhwCgEIe8oA7NK5TFh69FX2C8IeCJeHXlS6CYoh9d4TQSBGc8vxpVKqJ
y3zyMYKsjABmgrKQMiRzQOihnltP4CBHM1zKMN90IvCJVmQEQlZnnkCPAO8nfhe4eJwXnQY/jBaN
8O6VbeOaR6P3SpRDvCgC13oFlnO3oUlyJstqkc3XARJn9ZvOyBGooe7tdmB59766LHyMKCNDhLPN
Lg7PSSMfvMA0DJ6A7u0IadzWEAu1AywiE8RTugRiYhh0ERwDKyzZ58piYLlQifjagG5AgcPXeNB+
JpCLiBy4y/Lg7aq276zo34VtHG762eKG3/o7mZXt9k0j3p0Jsm9T0ygWz7TV+JDnsFj17GPMEW76
Yl2eS6bpN+9ntWnBwc4TwhCMVLtVEY1GS+mT4IONkTfwFHvsmPrGnOjm79yl/DR7JGC2GwVOtQf5
HaV8nhNRkhkVMMZ7jYbenOEHVuOF7LVUugHd0POTu9P3zCbVywjVL7Yy/+wgCqWpVW7/1eGtW8xC
1uFn8G1foV98cdEg+0aRfhWJdc3Ty1ciZcfWzEel62f4+uGObklQkbm2Vgl0OzJ4WTrIIFKSM7pW
8NvV77qyovPwaK1ITuHh1I4jLLwrYN0xHREEOm1vaBlm3VlVdD/9B0wPcvZJ2dmYJEGhph4jafqj
2rwe/m105xxxl+dPfheP+Uts1CYCFW6hJGlpxu0IgdCp3vTBmZ5rUBC2FyubqdWlwlfMCrXbhK0f
EAJvGoEIPz0mAY7LB5P5DgdHlGMHqsfQgkbzqb5Tlu8zvXNZacEqQT+1LIie0RuTYFAzWIcxMZj0
MckM4cGwNjFtBtxBCvpAe9Gm3kpeC2WjPusSExXeb08vCYKmq/El8WmWi1BINAsBSBPDO5e+vmM2
IS9C1mlmBQNIMQFEM/zxWKI9NjLJKTzeF/ONzBYq02WNMimsW3t7Ku/Kou2o1B8Zh+6EvY2xfRNc
eY4fvWgWa+wKiSectMfLBPDKdX89uFVUi1AwZx4Hii2D/XYL6pnweqo7zxh5rJBHWWJXrlRR52Sa
d+WRbd2AAPnwhYpeHycpqF3Pm4c4GshtMjkhHxwlLdnP0Fij58WhnnOACyxIhj6JfDaJAUVHmNTx
urVjBx7LkqswVvG9drEv4xUdMfv615OyLaffpxS7si5y9a6l7gGijWDqqxw9XhpDaER/BjoubUTz
IUkVf3/Ek1hU32MHEttYJt1cbfwF2Eli0Aeq9joTMPokG6a7rzAGJgsAfcnUdScj6lj3mAjtKHyx
F8vuiI7cVTaqvqxFQ1aYMEoT4YgGbcuN9Qp3a+XOYqscFK8clIYnoI4JH8KfEyOEZLLw5utEQO6x
K0qHCRsstUM5lNbXfduWx3ZrQ12NGQW67QhME+bO6GDa+P8FkbxbcTzRtm4tuO/Mu3jGSehy6T6z
3ixrUjmogvYrgY3Yt6k7JZAZFV6JLP8xpErpsV2lMkkv0ah3TEMM/fXAx0rxHOltUJr8g1e+VwKW
7TVQRos26+pR/RZmii+78tgLUZGHcJHs67H3UWjGOdXiE7dvCK4zGpC15DM5N8kr8T8ZJH9d4kcn
Xz/fUn/ALJRVbGhAlauOzZaJJwjVxrpyhcKBXgJsEZb6z36JY/nh0LNl9xULHUVzQdfmJej6B8x+
Qilu4xzfBpMxweCKckkLR1w+CgOOLcfoRr2RBIzOB0h/0N6bnHlAQFi6xS6JuLSUakCbvQ4sumI1
ArWVxFCX6/ad+o/oRBfL5BVMDji6e9s2wIpgkMi+tOUQ/Z5jLdAlXIrC56fui1xfaV/rWjRmElm6
ZJpHYwgYx/xK+yftnNMhJ6pd7wdhazJ9oYtzaW0urhmcpOQ/PWtKNMTXPE2mzk6c3u0vwBxRDbhM
Ux9g9qK+u9SWfGMHm7cRjQ4rlCVhi8nZeyzYONspczZlGQA4iykOWKTOBZkAfhV326b1SRRFTL3p
wmMi4yguFu1eatOnI2zW1c48RqMkaQcl+miQjvTChuA0qdRUJTk+gPliA7ruMQx9v6GFoU828DcW
aHFW5jeVUJKE8ERTJI47MdurHr6okmwuxpVLIM03add0R6L0OMe3nzlpoIYBKqbbZRZVdcflzsyy
WrmPrM2zyCBgQ3Z8FIPegQxhVlluvKPGh7PdZBbmuIq809hti4JtOgCScADXIqUXddD0sZKzafF0
AWF+ilpE5TnchdAbuTlBLfxb6co+E1vkpR9GZKDW4WBWUvO7gD6Ql2Kh9o2XsePF9v3WBSZS+QIg
KY/lEtrPWtE1Zxn21iK3Ecc0MCkYAXLvoX0pXOxbQu18Rjv/lY7ETz05dxr5bSCqyJITyVmMu1BL
CSjr8we5rK6Xu8MGQb6MJN5RBAeqOjvZgRWaG/qK0GM/qzfn9dGbSnsDY9gt1ZrWARCtuosUWvSJ
PoEtdXfjHZBchjXTV703/HEuYcGAJxUvJWd3JpPLBwhZN4FOl3fAlOX1jhOLV43W3Eo3ElPYorLq
Q2C+iQCEiiFUY8zM7jNThsHKpMmTgCJ4lzXanISZVcdOqrs0czYVwi151gFID3Xd9nowMh2Ww41Q
A4fo3Se5njGJPyzfSj5l2poX0D11NkNVyF8JHzEtFN0KPgBFWph5J3ScQx8MlNkRvDcRoRvyITPI
b82KzQGEKvPEZRIGTL/Uzc6C9Jwtu4jMD8FdbAO0RIKMOcjPM+rHjjqHESTN0mdSA5V9AbVTRjqr
vBkj9gipbQQB9tozJXAUeMvTv6IIEK8bHryP1XfedeFmNJhayGWxy5bQp55IEmtTvSojFMDlAwA/
zL8GZWhJtmfJqwHWvChRZ1h9LdEFzDBr6iLKN5koZ6omXS/ofqZj0nTfo7DFx7whvc52x2hb60Jg
n11vpQBApfQx2O2Mmrv0OwX5D6Miqw0TC8nTy/3fULbAckthKB1wGUAohTDm70PJejVftngEwgHm
C+W6OoUnTUZzZV9XNxK19Sb+lYwnR0bRCi1XHx4tcsILDWg1ktZ3EdiBlXNm+3Rc1D91BiM9rKAL
p4bYwQMIQVSJdrmWijqdfLNOCBi0SqmhGWP5Zdf5h3M0wZqijWE3sNHhuctT37t7H99HAfAFtKMl
e97higZVLUPy7q9gLPNqVXndhx5iueWPSgDfgucm5lucdIdZQzIHBZ+1z1Lfph2MID0uzlu/4Yx3
FsDMLr4SHg1N4UlhXzF55jGATjP2uZj1G9JEMOiw1OPZDCCiJguacyPTeU53mAZ9WN9q8cdpco1o
IqysCkePICNFi+mcmB1527JQ9z9qwpF4Jm8+Lmqdo/d0jCJ+KNTTuVX5tFrZVzoGAIi3zFlceU2I
TOejjUUKjSJemGPrPZy3sOl1DIgbUfeHBzy2avAgY0GDNppwRnPLJdNbanqlVctw05pGBsi45Di4
Plxg/tBZb0owHSxwIun/jm9XHCB/RTy6eU5hk2feDdYVnn47aT9yj2MrIUQiB/mjx+BTDMg8UGAJ
3wMZE3j7L7smgBsrthO5LLguFesbRPmixizUIQ2G2ROUJsYVzuVvACt2lETZc4D2eTN7DEorYGBI
q3KYgxHo3bdqyH841GF80W3c0ZmitO8A+D7z2CpRN4Y8U99Y+ssUP3wcteVeE9U0BmxTFOXb6wu0
iBdCjZtOQXDqe4w+ovIZJKc+nfMLIdrTQ8Wr2c8uxlDafgBz0qx8T+poS/2SJwaWE4Nyw0YzEv9n
hVbmvgNSFK3X0msRssxtorAu7ugRLqCRS6g5tv1p2QFD2c2xsDoKGWEifo86Kt/Xdi3qqbEpky2y
Wb5cFMAyVvuNlRIRoLsEUo2q1NHrTb5MBBU1ueAp88+25Yvh3MLdBpysJgqswYRVowYHy9d/k1Ef
q9gA6CrHvrUxI4sn2s0kxlBF2LU1KL8AN74v3Dqfci/vgr0mk9rUC+JWzBqKbIrqhooDp0e/I7SV
KbL8I7OtPS/eYYBt+lM6lCrZe4j5bddEpqqNj1oRBvgnuJKPM/GUt3iGSbb+krMz7Xy9wAK5vV07
M2/LvKHoQIad//h1tpxa0xnAh9/oCiVeN2qRfEw54p2hK4ahtOvYgykjNAhGAGTmTyx5SBmY/SBg
v4MQgulGn/jXDaErfKgbtFuQwYdi0wp0BoFO5udZNvGx8SIBJwgYsgcY/KPsYCifFSFV+a4lf8fp
XdTG2CxkDrbB//XwtsxPIyZ3oWLs0eCNTkIJp57zWnps3wDcNKGrArCrqldJP2ArEqPkQkzV91tl
x8gXRhxq7gENkvCqH4L+wKcQK/oA8q32FSQMpzX20cX/8Dl6wh09wvec05CgAPyRjVZcG6WN+p7+
3jnAlhi9ShFQ25zjkr2d2YX1x/o0NxEG+Jdm6WNp7gXpbUtlDh4sHE3MUWrgzRiRUqwcCRGWzJd3
7CWr1I+sgST38xRamNQCfW9uvKXYBC3MN+6gNrE0k5joFP2D6h37FdfMNrvhYzAMBKvLc6BqJwYG
f5PMWmkLhMBknsyrMkPMRB/F1MOwAzsSUMklHUiyRW5pPoQkNxggEeNbFWv1P0+D+Vv7GZBkDGwQ
JDb9ZVG5a546MokW+KyoYTp4BvJsu9C92et6j7oTYPoeCDhgW9pkjcNHAMSlK/nypsBdQLCbSuxq
MaK0A2lXE+/4f79gevICDeLasteX8R3vRAB1g3tdzbEIaB1Dc6cfTZ+v5yEf1r04qBQPN3h+tIq/
MxRJ6+H1Ma/TjHgiq8+SF9d+ZfnVVs6pAE4wN0cLzgHr1B9VvP9hEWEVGJnpBRKze/0d9x6td3UM
7FRJIlgNs3px/PLxHVQEtOiodgChSWbk2ckl+JN6yPYHPdR2ozl+iVtd/a7IbpsxLiy1ygD/b3ov
Kc+sR64wsRhCahIwCUjyH6oTKe/Wvt+dOhnEGCphnI2THiWCm/Cu+LrsAOfZN5nJsjaNV/K9L0/S
7iZXkV8HTJOF8dvnmMmmcit8b4ApPQaYFpO1a/+lkioBBfxx1DDtkfdczxLjy8sfW88Z4W43iOvO
HojLo0NFcgbxAJFCLT0h/Ej0P24Jh7cV0kUcFDU6folY9gii7fw+gShqGRRJP/wqJ+a6R90GARSk
DvNM3eIi85mzLMCqXBnJKErQcb6n0FH/I2cVnY8GlufnfINvTwPEFsNbs3d4jo96KNqy1tFi3/ZU
0ZkJD1zejDW5xFml8hI3aVYohBTpyL9FI8k6KysU350rdtHhAUgKlGwV4GD1+e/TUr3T+D2To3Hy
+dHsuT+qNVsYLDrFNXyuudXPxQe4ITDxe2iAeskhKXOlYnR2gPBm4+wOEiL6/hkVF8JKl7w0LdWg
1+kN7fm/DdCE/+6EFW04Q5I9orCeJwS0R8Ni545YQsCGWdBAPupbCkqeZEJYRes915X9V3P8xunw
Gu6H14oW+tXFVwAvRfzET2FGDlERuC+Fg6n3x/Vld1lay5zIo4MAhm8Gh6znTNbo38Ul86QV6KJC
2HmtvndlG3DtIJDkjiBi/mTfimki5ean8jke1QDQZARxtAt5YjFmXiyNXoWjj3xmxx1Lh/KmxSDU
2oo5IicjHwdF3PYfxZzcOXJ3WC+cRo3RsC9V+WsT/T98KTs3Ma/6xFvWW3Nx0SiLohY5yzb8NKQr
ZGC2AuNyH1GW+CF2wvLajKgDejhlaP2THWIl+P6IEDV5413ygmw7tOEbspk9TjG3wFpHq758prqu
RgktjzgGJB2l2P91SQYGthxd+bVJuCYqtZAgl+3dPR3CPNa8V3DjkMF7RL3PVq2k4VGRR+epgDOV
mlkConZ1xVgamrK12daWb+Uq2X0ShEFDEghsq3L4SRet8roalC/OZKlz00TWU+rAh8+QgGTmCVT/
/dKSzoDLOWd3ZMKT6zzwGn0EpFRSh3ArTCDG9FPD9nkAwPG77RUjwpVE1b6+K0wfpy/FhOw9YZMT
lIk09mCiFrZ/YnppjfeEq5LRp3jj1GX2VfIPItpd8kJ7FXfPWzLmsKd8FFBW+qcu8Zp2BC4P6Xq1
FlqiATJGkUAfxpmzXTg45Nh3ipRqdi5oizAVSwXiL+rAlhzRo6FLvJmKIjeHKy3i+VmLxm1Nbstn
yW7u7dmtYkLjViW6BfZliGzJteFevmVY8UlP2FolUlEEGlKP7fWcDv6oiveN3MkCZPxZdRaceC/f
iOSnF07Lr494836fBKw+T5DHl1VxC/T88T9N/FVYZ9N2ZFXibX8FQtuMdEaYxSflpaGrfLRX9MWd
C+KYa1DZtQ0Gsch0Zs9Kv2KjoQyWeJH0TvJnGSkunxUV8OmUit265aLuSit3RL4ec7giZKqUx7RT
bBlnTRJ/ujkHislomv3CIoLbG6zfFEdKra4b6XR4Nlv4Tcdr/6llrHBFo7BdPgjKOabmkgNqSRVO
ZsieTe/CZR0mIu8czgu4vXatlP3DOF2gIR89DHQu2WNm227bkk7eumuzrZA0n/l/6oUDFRxDP2a6
rfTvcaUg5f6G9BBzcCoX0Uhel+Bf+8+f4X+Pojnzw229EFapRkOKNSqfO1CXMa/aPxT7SlyjggsH
ONjHxPyG3CX4QrdL0KOmM1MfbQMR1TulMQDs2N7GY4gFagQPlp6ZvjNoAV+Q7dx9VRvBTVco1MVk
VWa3VYFuDn4QyATbK5QLYVlN/TOn5tvSf+WnMuLRdOkQDKWq44k5HxMFwwbhbh/QgDSr7uPOCm0P
ir8tB1VP+jsuEYOeUQ1NH5+L0MjYd1iV41aLmbldxS1riNRU0Np7DSpCoxn7tJSYFfTjhZ6+piYY
nbUhm5VP+UI2d6mu6yZmhEZ1pZUGPGNmkBrFlCQdGdFg3PsxVzq9RpTpIV7Ym3mRKt6ki1H8qIuh
oFMpcxgL+9Y6vGdizPMOSH/9mCsIPDiJ2afYzlfvOM4HiJJgmv9fIARoquZ7+UefpbwePk6YY2Dq
9EXbmJYesGpdh/eSEAFTPuYnScrC16AARXVWuZJcxBdrnUI8PeD+JeMmuTCIWdNeLzXrwkhpjrE8
PxOd2CxlBvmV2sAq/2FHp52zSJjM4IyeYPtIEKkWauHTs9NjvRv9M/JiQGcj2z9EsXeRTEqTyEoO
rZQR4h5JBKGsXWVQ/1QsPbiBuzs0R85CUyeGLwdt7m6h/mpUIQ9DsaL7X6FKBU7mHt4E4OKSCnB6
dRnaSWLXyzwNlqpK8aWUJlJUgIk4mixOdjftmCU/HPpRP5M83uVQgWqGIEToepR6RXE0hQN6nWva
TdyWFo8t0v1v+I1SE2vbTWZjJqY7ffmrufA8As3A/ne9cjwzAwDkubHxNLHbQNAqLKApDVZa+iy8
5wsUgZG8XH6Jl4KJYTcEHjAcOXACUhHTxw+JI/pneKFxOETtuKoSNmDNFc7DiSAVNCoVAQAovLhr
fdaAP8g4UdoYHqlBlQjqnMGEOTIjad1E1BQ/Pmm/tYr6o/Cfz4fqPxJ+9NDW4qF85NmPJiOWi59o
oI0BdE2Sa0e1NAeMvVR5LLB3QoR43rn+7yDDBL2G01Ibh8V4AJYYnDH9w13lJeyzsB8IdjfRWQ3j
37qST5p64ViRRcFH+DG1pdZT7Teo6C0cgpaA5fht8FCQ1n39nwvl3J3Pig9N63BMFz3RrBqNlgxi
x3i6rhhZDbWhspMCc3E0R9LmFyOIPPbEQ/rV2Za+4gksW4H58XyXbYQGrUl4KIEydLKai9IFd2ya
cw59iqDFv03T4aSfYvhv8H1Uk+vOhlx6L8Rz2d8o6o0nXn2v0aWTvmL23fcnJakEuwsa2Klkv8EK
t3HxLqSLNebYF5RqM6udXIxMHUTHe7T5OyfpjFQ4XB61+AAm/t3yGAf2AKSuxDTUeKEPS8zONTY8
8E0KqsSvHFb8ErGfFxkSKB18V1ZsW0fx8KGrF0TNQm93Zn+iRJ1ZfwCIpnTRm3tq6yZl5XkOer7g
HlCNg37ZA1LH5cFuSnsL1ygTHAJS0NuadKJ0FGg8I0DftH032+oufaj5pAhTKDG7wDDsMKE/M7d/
WqR/BlmC+/st4Ls1c6iBJcLCykfm4jNUbUB89Elj140j3JUj113fOr0h6Pc4NJUMeJFHunV6imZU
RzXZesJ/D9ZcbRSgTIuavLEbuJfykHEAajd19uZfai5PiSvC1jd2SVusc9RpQ2A2PVVI4EK2BD0p
ylIpPJoC4aL+teiBRtytpWAT5Fo0nb+XUQUG5q0mksOazKzVN39CblR10Alh8EwIUQLoO0J6Mw/o
AgxCnDBWI0h8B7EkYNjDIe/NFsLRNB82H3fV0EZaOVdVDJtNSIL2cimfDLGcFNf74YZV65S3wr10
u//vwnOGuT2vqT6cehXp3fGKw8vByBLZITOSk/chMGs77mquMZ5eDkKuAuTVrZKRwp8NpmIXmjZR
H028HkkBhIC6nHPgS9CB6vqwImyFkJwOSe5tuYZUAK8B7U9OkywSWEB5nE4T2zVgXKs1extEawlD
4iODeagDSc34WigfkzUYsTKPuKa5o5/gHluT0Sm0PVZZIt5ZDRQj3/x40dhgRaUsPr3rnBUa6Vei
4nWQvvVrLd8URM5gdTrMma4+AEbMxJeSLuE9xFRLk6hqD75pHjWQlZU3WwPB/vdit6humxlwRbly
MvbX6SKoMrbKdRbiXygRFVBuIqpAOxzUvJ3Trc7334fXmhaN94Ebd2NStbS3wk5Lz0lLTjhtjLHD
/dyV1taOoSmkvysCCbbdhkfrorUKbxg2Ov/h0U2K/XzQH0Ybc2zJOx7hSIusEWxfO568sr8jxZJs
Kd7E3uODZz+dNonPiSbIVthnz3RR6L7aGxzyAyxPu3RvoEfBEgcBedcJL30EtUAquF6cHzQ5cbEr
LVrVIiFngHhplfOPNLsR13B10P/Y5F12CEWCExA8ECCrP4s6jIAw/nb1uDA6KfTkDy+M8CC377uJ
FMEmTz0O6S1YZ4syOJMfv/wVXMp7V5ZlKgXhNwNsGOtZXgn85c5W3HH6e2bXbWxJfC/w+9uAUoq/
MqkAwH5sjvIvMHPjXmfJ1OHPi9rFTV+AwBIe5X0/9njh//cYtdyMj5Seu7jc5nbUAjR9c6yXE5P1
t37Mdwfqbn+SF9WkLC5QzwsOqSfPBK/LkD5/C9Fe6Ce6UH8+bYoUpQ1GrLSJKQAUpjNVyoo4TtfD
bKGS4kqkzJLYtvqpXjf4eLcSqrkvRw2kYNA7rs/q2pYbU1/FRebeDmH/WIX4hK+3vDo40aDVNXS9
Lcvp1jd2ad0UPyu2jlypjFXd7+VvJp6K5eJAhuwb5a8Xaw0a98BOOdwXMbrzAjw0DDAk1MO1pcdS
zHXHATrvDK8zCVfyXy0iCj+alm2vCCyq3+FPwsY1dnaEwj62/tmh7qAJoLoAOkXP96Ze/s43DDlu
T9EgZN3MNXanhXj79NzUxgNP0QW2NfUV/jqaQMFmsnoRolrIrsKMEdr1TqJtVW0jKJ+QZVK7bb6t
StYLqYGUpJEvNBFTF8aVwWt24H+DWum1ZO2z/qvq4EZV+DE3iSITBJRk6hqxX26d4NhLJDcyGPWI
q4rF9NHxKBEwJcRMrO8Zdn+Yy1orGA9y9OPNh3dS8G+B1Fip0VDlMrXye/bj7dnvtuxIkM5UVSzo
VERnartbK9XOLYSnSyTIrQ/3OBTf55Q+g2JhFb2S2lY7t0QR28w3XxwaWXPfrD1Qc0T9Y++ycCyT
DcUjQrZ9EOu01+9YK2N4eFHnt62fyVVDIyLsAGI7t212o93aoh4BL62g0uPA2JyPwhuHXswUIccQ
snmcpStKbYgcRuT58hs2Sq79pswT9P+kDy2LagWqattQ61ewLyq4x5E60UIJIW4JM0173tg+/AEU
IfMbizehbggsIUI6yLWuxd3fKyo/zPg9Hyagx1r87G+ZxvBmsASHvwNJ3hY4gJd/0NDLRVJl3BUZ
M7xtQmXOzvgOXvK17uOR4fEahhs5X0TqGJTxcvzzwRVGIqOIpvaxSRU0IWA/uXhYRvcTJvnNXdPI
BbU/38DvBOZwtBDEMNI3cMiIi2dq83WmE5fejWq2f55BVJKvMsux4ja+tW8Jj6A0h01iCd5CD5Tt
Ra2Yg+3iwbYatm7yn8TQmErbI/vjoMIaUEaoXAmoOiB0+2YKbcf3RcQ1iLwcXPRh5I6TzH9RZsad
THN8HKUqlUOHGSLuLoyoO9ncGO8+3eXwo+mZPC26az8X4Zbay+03MMeu8JtPyymYKX+pGdR5AhB9
AhQhy74g6Na2yu+voxmqDHvNjjDBLEE3C0GZkr3lCAyYcD/mU1azWY1x3FSUnDMmr7Yew2jJ5gI/
F7mAzK8cI1AL2knpemMWLKhS/tb5p6uois2pUl2l5fKV3bXJKGjlT+zBMS+FBw4zqzhKePGOBg9Y
gmRCvbBoLmnA0Rto/UiYo0l8C1X/OIxrBLGqh+MkyrmWByFSV3HGUxdY/NoZ91wDyZoFeWE/S/V+
R3cvCCxh/XvGyxSLF7Xq/tKioS7X7Qpo7OBzW8yAJKmoQAwnzo0fS2kVufM7DAXOqIE/a6Jhq49b
MOBGR0pTP1UetPsoYMNbAyoAwdFHdcpzdl+TP27T6AlsDxcp7NoQawAJ2ynJr5xHMf6eKv3Zu8Fw
0AQq+8vFAbQA3goEc3ENnXFDUY97wgFasmKtgJ8FO96Z7C36Mn9fbNduHQtHeRFeIvDdpSFIAeDL
L0UUm2EEjPhTAfnDeHdE17N5y4e+gIDtZYScy2yJfdm0CWxO5wppkFua8v3EoI/vFpe3SgOOH/W5
bLpy5n3nkpRw1T+1PzyEs0YYze6y3k31tOF3MemKwv36tzEAajUS15WrhIz/aFFoMvdKZ+snjHKF
JnSBPOlV9ZiQ+WaCcUcv4YsOaYeh6vAHCPkbRI/3my6NZSwcqfxFNMdydh2zrtR7z0gOoy0Uy3eT
b5oBSdHfPbHRtlxZ+MAGPAUmjsaSX0GvU6OBAMmvH49SMmAgkY6ubpjyimg8907DZVvAANSQMgJN
3hK6nZVtHmYqMk++uYxYiUB4BzZ0Mmeo8J40KFoXNtXTlcyaQmlxjsqGH7gOjakbZBZ33q3gR23l
QK9xg1o9EE97eFFQrHRyp3HeW0l84cUAruZXgdl0Ds5NacDSnpqbqDhPZ3RvyzMCfBoUfgBoeSfR
8TOXs7ewr5oeR5HfiFItcq3C53vualCWfAKypY44/c0waZSkXwsBjfL+7oF1ASXuo3OpQO5M3BfT
o9/t5tPKD4pHmNjbC+Ci9Lh/ZZ5OhLFBjdVHRRIvAXIDRq+fFxUwDyV379aQO2H0lorjojOKbuzu
ojRo9aHF3rVriRpsVi+iiPZwFv6djuESRgsAoQkGsHX9jS+PCExWYDWkWBAfYwxgwlXnBnacbVTt
yjIoUCXl0mRFa6Rt3tWWR4h8k7rNZ0tQNqFlPN2E2ARaeI5gixuzepwYX1Hnhqi/jQHkyj1mH6kO
kf469VBIVip2kv65SHs1m83cxbZKVh5M+eQSCtd6Qh8oDVTFTud4rhapwARKqpFlWeHoDYvUG1YL
T1zVfBQWccRg1MihsaCorK44R1THZW4ZWDgvUWNFHPNrKg2CKj0NxAlOigKJNdNcougxh7ZAhUC6
b212oHSAZN1qrDgT5YBl1/mkqxSoCS8P6wMFMWnAk74qtFfrFmtSU+6TDIMJZ+/34A4qAYQ56ANC
8JBokyTFp0/STbYTjiBNZVwkgl2JQLh8qmJ0xYxTBPt1yk8Xoa9VghuyFqQWE3W0ORdWctr2HBm6
5pn7lymejN1KJsN5/3FhMQsqW1Ncot+P4V30K/82ZdUvYjUzZacLBpTFNcWzbrBLk8OnOHEubKrk
moob8YSg2tlgeYTXPKg8mJeD6tKqHfA9dcacStJ/x8i+xcbOYwEEcN/mhZ3k61XKEED8LTTDfImv
+2djlGJzZT5MnmPXol+9nMPHApYX4bRGM7/dFqhcTmHDUCHAYQqw9feQyzlzaLTKJLDJPwN7SKCx
A4WohkOdH+CZWrg96gX/iJ+AwoHBSCGtgq+BjgbNM5IZ4cWqdKldf3/2jUDHLpdoxseO3Q8urPDg
AIyNybxmrMo+ve6T23bkanAkfiFo95CC+1i37vQ84eVrIqWplP7dQAdiyCnfLiIkq+nLKTzEzZaO
iIt+ph3dG4CSET5wZgVe4q5CRkbGd2QyO1anNAVeKGpuLWPYCBEJI56uO9fxcNXyy9hAoOxVi6X9
d1wzI1utTivP1TUFNc/PaC/t4NUzJR4pFAwuZ/prqV258DDOamwqOM6SqdmMjv3s1mTYngJ7D7jo
hN/8tlm6qFtuHmyvF5XkiMhnmWPbBzpiQTx/yqX2CX+EL5k+9xdUxpqmUkbgRfviXlFL4U4nMwT4
ZIzlFtpfFyfy04C14Y4EPGuZ2lijVIMANvOt9hFp4RohyfIydEp8rwXw/z61qPFp8qwpg72XEWnN
qNePbLamQo6aH2voOVBY2wLTS0JZ1quuAtX2kJclMbDMTPc1sqj+UiNujuD9ESuyfdj+mhHAnhdD
NP71qKVTKWTdzcrwsifLPfsWGR7VUXraaIOYVnnWe6DOY5l28rczOfeDmyqhYzuk2y50bFKKOCk3
MHqg8hMDwHbAoCs3v+gkkYtMK8Ol7ZNUqj8RBusqMMvRKkYEadpts6ruweTEgCmYEgxdEio30Z+k
yqEMUeEDtP+BHExziSOU/H/EHoxzlFgYJ7lcLNV0bkZFjo9xRRE0lVLw0x/iOJYjRX4WsbvFwSy3
OcAjp+Iw6Y5T7uCZVzKFgjGfa1mZKwxTcQFzuhnrKDima9Lq6Xob5A66C9AsM8k92C9m6yN4K6yy
W6NP83p0RWyTRRUaWqEnUeczi+eW9zAZ/pL7Q0r41laT3x1QgjZuiTPzIqeAsKzvdWgOSe82x/SN
GtyQ3kGMwX/qmQ7BZbSOHfFZgLWgNJ43DR1J4gczG9d7CiaYnaXqzoaJmezO/fDSfBiE5ch36mYQ
+IC+LXRbUWihMiPTfj6ze8ZVDOnXQYMbVbWfq/ekc0b32+eY9k00eL1e6/l71wxu5+ah1YnfU+Tj
zQPt1rhO0sxqM8d7g9mIev2r8lLsGnF0xHgy5NMbRwoQziH3CqSnSDk3kcn0HcCCgifx16cgb+78
Tiu/1fDUeaHncztZD3RV6FZtXDwtcOhtjWkse+E2BH8BkNpiYtwuN3FqYrhtiMgkIoWBaq19KtkK
IEfvGOnj2fJvLtJS9nsNLa/TsbUiTmpYeTID7ktRoV9v2Zc5J5xEY6SdFvGmP3q1gYy/RIJclbLm
/AE+I7MihFMJrhzNG59v1lkzJt1FD4VzPYfZVwFln93hdPtZMfwEwqmUbIxj0gys11Zy3O6ahDBc
Zi8EPjcowOnhqr/e8fs3+ejpVY33n0B7+Ju3WV2hlSL5fR8aWeVamqQN8dwvHaWuDrNQgh4e6y0+
HlwutwRLyaedlGPrUvKaCki+92rHQj+bqYLOUyOE+rWuYo1+/aGJpNL698Fu90G29cwuFRKJkX9k
MYgHh1kTgJ/7gtgmY/lmO7PU/6iXOtYd5Y97PgR9TMTu5ytIKe9C4dDvRStxrBNo0VXfaevuHC3D
W9AvrWfKm6oq27FfqFioPA3jpoHvWBe59Mgik90I/Xn5W/6du/BAtd+Rpc2KRlYKARF14Vy0JlvC
64Bz+hMEUYpQZPyJ1O27HSLJC4nT+/VgIOTvRHTP75JO7XBMy7X04HwaeUvqkqJNuVGQh7+BUl//
fbSdYQ+R/W06z93VmmlkMKtQnbZOOgt+EOjrxesrfi75OoBcZXvMINtfj9WzZ3onYPcmLRz4hhLJ
8RL3pL9puui5VRu1AxI9Cy44+noiN8bqZqsUabpANj1GqjRbo/Nk9pjey2DRjJm8wDvXvzr/shYl
KYQxteLVxipc6tuaRKeNvfbgui+q4QTHkonGuAelQxllwkxacAmlKrR9MewJQq3wGd9+Qq4lthd3
saqbXURdXmAklSrGkuTK4oBOxGBKE4zGqns9uABMO9C+w10oaB0ifKX+y4+cZmZE5JE9dpQho1XF
oKqfHj3SmQH3ectW+YXHIhF+A1dj13bFS7uOnPLrVIELoAAwD3ZYilFhS1RHFs2De5hcRGsJN2vi
CMuLmzibfq7WlVVxPNWvupq/LjqsagqU+7R/5jRkroOXGkeHEffhc+4MnLuHz01nxPCkm8WwNvYG
Z3lDuyDNq+o4XFVmghCftB5Jgj9wE8pZPRL800WaDtxmVOk+vc8i2ZbHoY4ovGEOmeDKhtM+7IRt
q0Yo7Y3QOXOkzPRut2R+4iO27yAMUZTIeGmIGH2gQcdGkpikwq/knEbshLIR5g57jQKwl1IgXYA/
2QdimQgRUqpsYg980hR1Lvzc1rdRXNv0GqUO03dFJFXQMziVqEKprttN233H7R5WWbD8o+nLMZY+
vam5x38Bq2WkY0pO6GT/8FEWCE+u+7kLAn9TPgd0NhX03kvcY/vi/aim8Bkqou6/QVPwMrnIYnpP
EBchgSf04c6SW02E3XSXeTL+a2XNpghiw86O6svOQ60d5xTnZ+FNgRkff+lKUOSlu+7ic6Lior+f
cnvIS8G1vQ3a77QKixrP/MXCsS+2te7hpKuvGcMHYiMDX1a72ANYs/wH9R7d5miSmCsX77ceFWEn
+2SOrxUWV4YkRuFaHASP+9NIVoLXeLwZZVu6JRYphcGqaODVA03Qbu4F5miA2fU7jxndUo/3KFkW
HXSPApEHLThuIfLTENjv5Pl9ehL6G8n5ERMJlG1gIxPUmv7gDmkKDzkiuVYPKtR41iO7r+y7RAJV
ydd2KVOivIAH/NJJ+JCV7SlpHg6j0DF86OoCbeOffqxHkFTvAPSgbPUjoboIYN4ZK1WHS649nIFS
pafeZPjcYndccDeRbmaRA6oKC+uw4sDhs5iImKP27PFAIuvxDAcoKrKrosN5Ssfr/9MGQjRaUw+Y
eNXqr7QrhUJZ4VVKEck48ZfF4xQrcdWF1gHPug+WmOuxZRlFEv0qX6qov7TALRBK76lWtkHtWntP
6TypLqejS8hNg6AzF5iBw1T6ySjczKHrwyLqvVR3KEMQi+Ion/Hs0BGJL31MPGhwJFQLnHnRNtRE
GjaywXs8uQLK9oHf5WeF3w2WXYoAKZLEjZJdTLDl8NYcxFAB+4mEnklJjQNWhsoOCrYkRjRHAgDu
zT5E9ACbLVJ6N0Zpq/3Vlzg1QSkQDYcL9Aqazo0uLyfXSKP6925f/Ai7K9gHG/vUsvruOYt14izY
9LAUGYm4U7lDdqn9hGbTF6K+lyFAH/ytfiGPU0Q7PH6X7oyyywxiYw+3tUaLjJB8aaJhUmx4M+4Z
TZLxU7+um7yxkVoVclRg4cONwB4wxv0fTm27sJ7Ph35zXI62+ooVvHos7mVi61zMDCj8qVK5qu1T
d/4IeQvUPKxrSXBA1lgjraNSDRuhNfICvOpeMi/SBlv8vt7j3IAwt2AcuwobaNc695BJEnf/QeQC
cFoxY07J6GiYPrnwUh3M40U130a8dwU1PqGcBlCFq8Ftx/nwblZe/pPfwvSPbhXp95RObPZ8pWIb
1sGtXeyJsu8P1R0S/AIFZ6Jr597yKr/kZTH20pJSUUpFDUqbYZgl9o0EEwOFADuEn//yKTbMrBOg
w72cjhq7bWuGy1m5VjCVyUw4asi1MzgpttsatLkSBwheLyCXv/SylNMISpmxrA1RiZ4kKEELiRpP
zznJLRjfsHx6M+VOC80W6u7iocqwT1RHhEhgh1NhXawQR3skEYgs9kCXJoc=
`protect end_protected
