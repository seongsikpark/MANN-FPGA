`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Nr3OBgGGKnxUK1X7rOkaBJKORz9hWxlVg67yU84JjPi+qqIY2BbPnqxg9btBjHSbZTu46aT9YbEF
/t4oFGAb8g==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
K1CSK3p3xsaXQsNgKc2i8PRS39tU1RH++HdpwsYWaN+qNGIVQnVt+JVoAzlzBpj6Z647QJmWBFno
UGBUjkMbDwf8bO6B9myMTDnd3IZBWKuiBnOc4OVBTqrv88TtHVGIzqlWb4ecD237g+fkiJn5YG1p
rffVTwfu8WS2Qs/2QcI=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
e1PvTVFVRfdh1BD8STKPLjONDFsN3HeoexQQfdlCSmg/DEWm+hRetX5NmzBkg88dnafteg1P/aii
wRNn0c2v0ZKmCBkmHOC8POUoDVMv8dEmEj6sU+EUGG6BfaiaLS1D/nVamoEHCCcMJyhqe3GJJ5vX
6UK0Ycy6bqzUJLiMHDBESM1Y9Hhi3YaRAgRsVAxAqLM3DAMOjtKpgh1MkoQcNQh0/+r+7qYDl81n
PV/R8RqRvodx8MLPyA83UYDFOA9PWbXF3qfLSyVcilwcXgHr9dFLx4KEhnECHNwDSMg4ua3TfcUD
prs+Z7bn8oJ05hvJXHPBY+idRArS1XZvCxeJ2w==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
X4SZefV6hdTXXcGMz9CxJ2xcEYY1/phrYlztUOMP5QOjmpn1yAEd4H/QG6ngBe0N5epfPSq6b94l
ZN+pCWaqCEQ91OGK77HFbZbz3u33UjGzMmyN7pdilvV9zGMVWbRtxS9TqXMwioMfsu2H+Tmw3mtR
3+LfpRnArcVOUo2d8UQ=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
fXWIkerFrKwodOugJDC76vUXNIszcxCX+/rNseTQVldCZKHKiTV/1A0+nCn2TFEkSkiSd3AbA9GT
dK2EUPMoJqBX0q7VEgPgaA2hSWqTEm9VBDCbLTgf1jld4Pir31JxiP1JQRSvqHaD+xfup2dMSLUY
QQ6pi1205XTteR9+lCnOE5SaEAmypd0cGp/cceJCYNQA0Q6VgI9tU5wzg4fPc0Ou8ZmIBrrjLM9y
rih2RaSOUNGWP+Jcakpkye/rHnqEICyFUdskLlNXIqPZqaBQaF3F7EaQJHe0YQKiyami8C3VFsaC
s+scVitA0rdcvRPUDDG2X+c2HdGVVN/RiJU7Sw==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JS5yxYkrBQG93S7nkh+CVDNZqZGNl+Y1h6T/6Q6ESQhZQY0lJBggpF1mdae7aV4oMa7U6LW70h/V
Wo4XBaO0UTGuTgHhcxN7MT/UM5fry7cOKS69iQAQaXum9BdVsRqoSBkXSH6NT3kMKW9nPuHNVVIy
GKhOjb8Ez4UGl2iFLHnQnhJ4QEIGILiAaeme+sELhZoIV1VtSlWndReDw3sUtEttCTB1RAKuQzwa
GH+BjvtsR0CO2wz1CV3zGbEUYzxrypq65WvQlLDx0rHRq+CS1Tjkg3FXN0S7lyFicIWVC5qbreK8
2nvuBv8Ys0qewZS3TP7p9Gr7SaoWzxQNSyVgLQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 114672)
`protect data_block
C+47WbjY8HdoG1QKCzY39BFqcJb4mot4LYiLugItx59JV+INFbbMh4wefAZJWORQwwq5QpovdA3V
xWLiwI1gl+GPvpl8wZiAwiYcBZxNt5+iVw8FOKliAj09Bc8/H1zI2i+jB6wJF805NJuqpQr3/PwQ
zcgpXs8mxbhXyUFpMksCGgHV/XIc53NXr2PCGcii18kl3FYqpee+zRZNckcJkNeZCTLyE7LjxL4r
hKeIMXBLfQm4w46iEs/V3+7Ls3V1AvnERhdHLsjS2eYNiCDMcSqm5hF7hcQZuRl8605+Pxi3o8ep
2fA5HkkTfYiBhsDsKdwu/IuGnrALqCCXwkFPn9J/GB37voxPnIsrZrWQr+VGVxkHIpYnVdJ/6YPl
etGzd1IBra/Ih6QPpDitBnFObt7kK4q90Yqt2P/2oqYoMib1at4dEvJmzzEkJUMJculoyDnhJBZ+
zv5BXQPXRTNCXNCNZURZghy9jcSfp/FJQ9DJw3uu6+KCaG3hYY8OIkF+nb5mrgDFFUMoUq70SUr5
dvcbsW5BJZaE/oIfNa7iSP1ZEKHB46F9amnRlSL7aTp335Kqn4pCHwffYzs7q1WgzslaoL8Xk6mh
cqJ5KoypHoDKKSNJDvMsZlzcHkwv0rGd2slaSaybjgsYu0aU7g+efJihpt8zqr30Awv2hrkn9g+L
oPcmxlgt9tVi47OhR3NkEnxgFbTO82lPeAIXHdYFp//P+92sdIUGVI2Z3nq4Wp3ain49/J+eyHQy
mldGDZ18KuzsTgs27k0PZ/8TAwK1m6r3TvrealIOiowTsXQDEZhUb4XKCuzT4TwEoLxKRCSNTP/O
GB55SLN1i7hXmnxNLoko6HuJKYHV7JoaBKfQ8j7HtbOKxz0eDo7WakpA18LjDZJDaBmXhLhKd8cK
tEyMxw+z7g1F/Bos+Cw3mN5GTmvXF2gkhpDYz4nJNMJ/UxgoI570qmMD8YPR9q/1KwirPbYUBY3E
o/QtILrcx3LKDibVn5yCWQf32IvYVqWepxINyJMcJV7KuJgrZzIMOmrl0WjfZc0hCYnd/Ycgutxl
P63M6POJo+HO/DvCcfjGGkJ6OeRcSGog75Fa8i+ylsNDWnHezlzpFOlnDrMrTyVCp5kW7YSjBBoa
jZH5VTjR3p7mWAs8mEWz2XBH49yxzO2+Ye3eRZu6216QU9FEg+QSHsVlc+4Oxd3lrV6JRpqqyBme
9sfK0iVsIVhsaFgYNf00tFBLdU04ljn/uZ11KnO6cG7zU8IRAz8xL9bwm9yJNRrkObNWLaH66tmX
x0l09NcKDFu+KeSB1d9LbW2fTjGnx1IAi5j1Sz7jU1WEnajMIBlN5Qm1WILcGPAJtPlj+YdD3Ing
HRBUlFss2L22pz+Okm6tvwwoEu0XEkAdW2JFipnnhTbCFnIukX1W+dJyrEu4CYiBAnlwGr4PAX0C
1wMzObsWMh3NVV2JzCyliUKAryVwfDIDi/FxPt+fulIEJSSx1LggJRQOX6Onq/A2oeM13U4Y90an
R4CJNwPMKVcI45PzYWsiLM94VepyMMStOkAUmn5A3MQjFZHciiyMYkXSGlyQFhdpDHKyQnCFOZp8
jVulCSMPwNfxl8JOOxlAVk51cgsELr29vXoHEXPQQoxnzslwIXXCT+ybWpbT6Xj5KLSiIjGNP+AH
IWnyAvWUAN8pAaEi80w9azc4Bhm0w1cFTgUmelHqST7FjnfiRO9sGmeH7/zOj5OtybKljQPz9I7K
y+Fkj8FUDBb+/aTBglETeeMCXj6+hIoVDhR7lYNO+1qKZpOmtN0htyaTA3fzLkhkrN9L96SgU5GP
ytEAyW8f8oiQRsWx7UjwCFl4b6pS0DDU34MrF8eHtBclFKoWnMjDrHuqMVWpBGcOYyBdgn9731g4
ATwX1ibPWsXjRNqfuph9UXQ58EH1ict8symbK6JL79KYLIbi5Ycec5C982lFfnrJdH2cTNfN9Mjd
Lo6idmH8a/Va5cbvo9GiBl6D/tjz1stvnFXFBsmqGoRdG99BX+mw2uLXDuhxSeMTxZ8xvph5LvY/
tCNE5T097CFWTK3O5VImx+og8Rqtbz2RXWsO0bC0s8wFFyH6HueS8uqVwfkb3GE5PSrgWQ1TTbWz
Cel1xBvml6Kt6S/zdyhDmmeAV13++MlwdeQe4e0T7xo2RyPehHs+3nVT+WZg1gRWoB77Hc9js9Wy
8WYfBWZR5de/d+ZwTx2E3gvI3njlDMT8rj/inSaHuILNhOxxvWoBaWKpjA17FbNc8fqFAYayaKzf
kgwG+bp4vmyFN7r4LfdkglvdzZC3JqNhygUUES7FB1vshhTjo9ZR2b0mEyUeSTmQP0xg3n0rV216
zIznRxj5xbZVsDQOia02cGSK4HYqzNfvClfaiOhDbXGcL4W/OalaJbk6pG5Z1IkE0OzBP/niuqG0
BziWr9AEXvZei4ELaU7UTt/78opi06/AXyQGhtlTFXVbba0DtxWuIsJsg5f/cFuAKMw3aUaWm/rQ
ZI3TjpN8sd+p9rLf5u6Qlly5vmxqhnzFzeXKdwZWTnQoFCj51JbKKu2J51kyozQA+jmLgfr3wy1C
tMC9DXltmnFLuwBSGDMISaC0LIXYZvTKwoRVmnqhZmW9TR2UblRSElqaHoB1RjZrFBQu+xzUyy8a
3pi2PGDbFa99cfBSiWSZcqWaJR0o0tO3NhLQVURHjX87sh/8l7d8N8cTW+sHRrxxzdSva4mG2JFH
mVvffRmogn2pVmj9iuJkd9TGd/DFdZQhtusBvDr9WkoRcTL2ktJWUsrSgsDFn3q+yTWJ6NGc+DsJ
4FCGjBQ9NQ/eJK46fspQbFACpxWT2IOeFGwPTMbm7tGSqKaQEwIRz/nQfgDxXVxf6bpLdx4jVAd/
3TyiJYkDSSAcV1coEed/ONewcJ59GyFzi3PaTXxddrG+ntHOcyUncLQYTf9uxPZ5k0lNcgHCi6S9
eGMCO6It1HKjrlaWHvrfucYuTgsBTosuXSpoTwGwirDWsGS4GEEFYolohlWMf41EfC0P1/GmHxZq
DVNBDGAqFXQdikw3kvBGOviWZUHk3wFEJUH20ZVmhM31tRQpBAQVl65Rd48cXWua1FS4eJ06Bj+g
7jO3GL00OPM7+9vuOtVw/uegY2VwyA51o5RwX332J8BvsKyPx7dic7X3epuk9vMJ2Sv4Co+xquTb
jsXf3SeqJ5bw/ozaE8klj2y7O4h+VcVuAVgV8RMwpUV4mPGreNP2ZJq9lEBiWroKXiCr56iI8XUw
ZmXFxQcNFMf0dDuNq1QbeUGr17DxbZzCAmb6Khw8RSByzBgxBh2+fmfYxk4+oaXZKTiwC2sfmH4a
nNEo1Ro1F8+f5JtaFXcIcRRCYhNZeC9/WEsBKUcvRwqDNsF2dg8smEQmnZrKlfO+BbBYSfacoTer
LkGLhyRxVT5xNM4X5y9QP0iTk9DG+n2yjvfqowZaUAUmn45FSSPNBAjpcCe/II/bN4RUkE3uoPAg
RwLh2sDDRv9RUCR7ts6ujUX3L9KArD6K9OwIjCWwUg8Kd3K/cdxXA4+tGja7jQA+HVKWNiF440wR
3/BptwzV0KzjpZwC8+dmhgdwrzxTTz+jkvmoIiBvPy6Y0kBdiHWIZ0C9qgjlThzrpoKrqg+mPivc
TAfOS7UdB8u9/B97KiUDYJWWOH0k0lUMVQLwWT7RWrG3b4HbncGH9/z9gy/4NIAhLKJuj/yup+kM
oiJC7+gcQZo2wI4EJo05QmlktTXcS9QmNnsbL/V56sYDBaw+OpLPXNPobxbcDHA8X/CezSzQQBYZ
rsqGyXDRcPLsZ1IDMuT7M+8w9xSV5Ew0mKH41mleXnyV+f/qDO/YLQm+3W7uY/aPNB8zoS+Qhcur
h58l8plAgoU8goJPAPitHh570DAKVT37xYtZd+Cj9pbkh4D2H/BAsuKfdxV5QcQzw66lvcg1y0TE
A/Qa0x8pebypziLZx+SqWiFCQQAL6I87L2fRO6G9YtjiFrxOFmEbxlAPmac+dk+VGzDkf67JiUUK
NOcBj4W2s3lYA7YlNJ7lGWsifexNLas6iDNSNRrwP9IxrVqzsaXwlrv2UTvZ3QmuMIu8eEjPiebJ
YjLn0zMG+TjjKdLpWokWz/3oqrf4A1p8+8QQBVc7F376zg9hoG9SkC0YNqL9jFBvwN0JyG1fOkE6
yv0TyvuxOSb0nU/BVxR420KFSZUQG8ZNC6GADaHtmoyw0indlY8DfjozgvIsBB/+Yb6YupdRokpu
wHQd1vJ9z+gN3gif3GHRkHWkGrodqAx/vyD8Uvsv9LudDVXnj468zqHKCXxv+Myhf7VMwiqs9HKc
gE4AFiihE0UVPIYv3yKwva2fbhDCl1oSnzarS5sQhYjUHcoFSget1Gwydxo16zXujggjoGLdydWI
A/hN/vvxSHXTSgCO+sOkeDdgECuP6EuEXFbikdb/WXlKBg6JJ1+To5B7NK2vLxJ2pB8WO4OM141K
x2dsu8tBOG5QCJv0vvinipKbEgR3BXUtLm0ADl8i0jyxORgfhkF5KIG0Mf2WsLa+B/lfriLiJ7yu
ZFMU6fHv3TUqZzTa+nNn6Dpg3mKGSU2Psa6DlNWmoMjvsh4KM7q+2SbtWizfLSCsKLgv4i/AS+3m
+B+AepIwnRAZCzn/rB6SWcnrkvKofdLOqAm8S3GfGDiedGSUuiNFM3/RtYgvHrrjwO3r+dQK+B3Y
Sj6fRaEiW8pDaZRVCLmpRWwIJVL+RSOxKqiHrtOZk0YZQi6buk1wvvVflx+QnpRiX6O3+fs71UcN
mmMKZjPQpTSXOHwBNZZcVMrWKjLzSpEnHVszCfVzHuAyjyBbW6B/0ji06eajbVTBq6VlgcPIHJeN
1yAs3NZmdc02bLcop2t98ctpVvSnc2TNquawVSwsqOiXX3RvtNZD5o/mEHGCBvIJwUkzB7+qq0fQ
AoqTnYek9OfRxPZLrsgMa5PKWRBfDtDwpNc7VAzuUrVGHkfk9XgVPQOhampVEhmsMXIwLsBs47gw
0LQW1pagC1rpVkSGJ9MMeNgerVbBF1vdq0xg++mNG0EdBtkEI3cCjEJqmKcYjwwNMH+p5HeEJNTo
CCIvYPI5Uh/+0Cvv4Z6TY9knEowicHsr8zf7XQ6YazR+zNspbRaBK0+hugajuGBfgpA2z7OTghVE
OFfW8/3VglzWnLazmGsjwB4k4xPA3KqP9+rjQYhjrz0sU2bJ+zfAF1ieDeZo7wNIWEFFl0hDs3Zx
GYWX8Hdr+ycF4xE1fh3GclnYY5b4bOrvB0qupBboOWra1+M+G5YvCJeRBxBf6pf8ccGIdb0XanvQ
uP5jof2ZthX5as613x3jWSrM0aCgEQ0mTq2cjFY08ESAyLzpdfcpCNltt+JBvL52CobwbNPuJaMO
kdnZcyuzcjkWyFsvxidcSoBHanit+MqQzgCedWFhjddxxVJF92sAh1i1z4JRdVKgtLIvsQ7fOCTA
JapVr3tu4TsaP29Pf7W2O1K8stt+m4Z9NZ1RNEROlESDVQ80fWKZRj3O09Me4f8OZKFv/uqSICfP
QZsx4MTPfKshrir96H0pP0FKciUyLgv+ou6vV2wK722AvLVp4Vxi5eUOrXQurnLcu/F340HTqmjU
OEI2NxLFapMlbj9HkO4ZY/j/qbwC3qaoanYJWg6WB28DcfvoEjeCS6lfrcUBTniWsohQXZKqMg7t
ZOl/cgDzC3CyqOfxhlhnBqX6UkiXMTymAgbZhyrZoSreHN/ZqxHrSaS5Xz2izGTnRgv1PsKqJi2r
sjT/4mly7km1tJoovzTAY/18hzgurI+XW63Yqirc0LRIg5ewuXMZcSxWbbKItSEe1e/LyYg2hGC1
/y6K8rUIx8l4yY7n4iLMCPHBPE2cwcmaEA8rKslDJyT+48/POiTDOLxgl9HjLKn/ITQoAkLB0deQ
UlG0Wg46vcQ7y87IhbofvN6R1fg+rO5Ph38FaqBOCSUrAwGanHbdfZAxaCaggNQJhDLoB3mvBf1A
ztG+rmG9ePiHL7Y++6Z8XEzclOqK57kVjuVmlbKmi4lg4E3PVlTd11lQtv+gydwkT6dutNQ9BcR4
dBOJNxZj83eEKARpdQMzlRSUYCtl+hRl5XpmkwsGh8ZFEX8IkMzz8dYn9bpmUP31PNpVPegzlLGy
AziVZ5XAUkOFLm4XmAYgLb+i0Hz/HAnPkmXuQBMm/xoxiltIJt7e9myEpkjuxEXLFRHhZwtaJsfr
GZ8jxzf5eRqP6WFyrBUpJU9ZJVllh5gvaJrcMReUVCe+yDl9ZLGsY0P1LGNmKOSOy51rT2jGhaQJ
BRgkhHG7JkvM/CvDHUqX0gGFoVEZf/gYY/QQMQ9Nyxu4NH+43Nyymf/hqQC0pDtG9crDSeSHQ9gh
nP2QgM/h2fNKKwkiC0jIRMG72j2LzivaOMK6n0opbIBwLw8Ta/qHxWb39RxQE24zZ88lLqXIZ8XJ
WdKpH6514JugmkN62zZaOJHZ+NlnNYpSDh6B1KCTLAZ4S1bLe6URuW0J30yAscVoRKRrSCwjdUfV
SbqmxQ0UE4OyB6meZhzubvvGiicEAMrws0P4s1eEcjL6ea8G5xOQ0sqyPC+7aGe3BpFDUqnmwupQ
G56jVdW2odGAJD7hxrOjs+qtH2313EFHI4DPEWz7VXQTx2TJQv0cBEorQBxsj24jg/mUIcKwTTtF
ezqC0t3GqI43WQbPl6OZPFdXnLhiqlMRF8eM/8XT3OmkIJ2d0PPx3INldekJFw1zQhMzw1ZtYo1N
AuQMkuiiU11bwnds/kYnpRcFHsvk12UhPe69XVtgLMxgyThEtWg7+QHM9Ufo9ryiLF1xB5XoBOrM
F26cgZjJgdHVhfPandSGHhRgPhP5Jw1GAxDXNCrzl7wmla0KXcoDDhEHiJVCTI6XlK4Qxf1uvJeJ
Z25NRfd+528Wby5hW2RXbgOsfLjY8XnFQ45moURs0dpguxS8QqVtaZbH/byHudiaHDDCz8TTwit6
GtGPsS3Ecj9w/ON5eCahDMfmgXxs+ECBJ1+NHBwQwAB25q27zbtSfe5C/KLnd3LWdjaZjlHNRpq4
tafnZ0k5qW9tth3L1LGONYUJvsg1gSIDCXQdnlfJVSxbL4w4mZ5KFbmB1qNrQ3I+KXBktmx/yYNV
Q1cLRbMp7SOwX0Zp6TYmcQwxM5rCirq6H2zgjkyQA29a+gFfq/nbu0oltg13N/r1EDd3asWJkd28
pn4NcPRKIK3OllErWM94ttM+YmTnUERMgrtapKFGedzjSLx7tCkxCupKZULjD7uFl3KBmrxAk4OZ
sVSXYQiTuKlUFPD8Sq71aTtmxpzHWCoaTc8mOu8fCaVfkX5PwPpOGG1rIg6UsMmSlU0rgwC/Dlef
rOW6ysYEihOiOJmxBjU/tSWc1C2CgH43akiYgErKRao0wyZWWGAq9pCpvLbKN8sbfXNAC6YhsMUN
1w56IQ7+JVrZYA7nV+4WYMHFdQlL9jPcyxx7nwUwEel40QGJpkgcnBbGk9kwh3AOtBZchJCbDh88
IJ+ig+2dojLpiK9IIt6X8z/GZ6sbr5ieMcVCeVll7lRXGtu7fc4c3FGb2BS5Jj0UNVhP8ne9C7MQ
JrHZ7rg0a+0qqNchhCv0l/kFIsOqUwOwHcI5VhMEkk1skHCT18LG/tXl4sF7NaIshmkUtCe+3cfh
pkV0kIurv3/KBgqewQONGhiG7PZEZkz863l3u3D+7hkbmWd/04VkzacjBKcZe/iZBPRlcZpDXxDZ
3uLEAreG29bLJUBjutMecSqCVEbNw/JUgcBM6BQGBwqK4MrBpogEH815/MNRnppKj4+I+gGlJUjc
K9ngBGACOuy1vQ/fRs92tAN28XErcxveu1QaZDX85/m3y489qCmvWrlzmiS5zN5NXb8i2LPHDsWS
GS0FH9DbIVdro7iNnZSqbRzDRS497AIyXrqKPFO+auXAV2XHal5/eQUpTCZs3xvOcfUOF60FEoqw
wK7ogINnpq+xP8rq0MCpWxhqWVrNhVF9W5j0j2lMs/e2LAckl9Y5pUK8vwlguFWYOI3ttQxQkTT9
YS/kL/Jzx/xTHEVyVgTjLFZDwpkY1YQy7b9fXpiSvqezeLud0GXvYf6SdFQKLaZb+9RdBwTr2Ne/
OsRdtvw6zCSBNeQ3xNyVdszxGZUw8z9ynhNti9v0cnqA7QEWHhYb9i4Il4XTEjcYS5SVUbGie292
hDutxBkX5wIhV0sP7Rhupp2y8f/32fgikI7RowI2GEHS6LNaTVZAWkTd7Et+n94GltINfOitKmaK
0IHIQm8guSVkAKhoQfPXkuv1ex6HHwGi61OrfcM7eFgak/kMGv0ydVFS6SfKkP+Cnq1fz5ugSKM7
MpJVEvVvwCFx19ZbbV2DdBbX1n6FwoYwYdWsM4yK7qoKETZyFUXovIR71FbxmeTzd/ZzToxsGTSz
w7MNjLrv6cOv2+V17KY31aEqPxG1nuf7WEmiZiA+eWOq31BsHpB856gMpMaq043qOgbHJprHLlWy
MLnMpLeZXb/sYfbUjVINi3AEhZJl3TYSALqGqr8q6zBzDVNAc4pYXq2z3cEXDkHelxUiVbT4k47+
rI1DVNALT0bTZHoUdEFYRNS1KDcC9GPfw6imH0ADanF2QeIPUCc67G39+UrjQAiTX9ckVh84KDwf
rYBD1bITex+G6QJ2Jq/qfyZoDcSwZFaTyZGTxEkSRBKpFzxMTUhB4zpvZriHB3s/Y2dd2+iqyxbV
yhWY8YGzBl14F1gj5TS7ickt5qTlsxTKL44q0fnZoWoyONISnIA8dDAkSN1umk1XWXsU0uqAZt2I
HqlMV7r1FS6AuPaylCnFOg8zh4FRwW+3aTd1LgB0/XgdqU/hKY23HTqm4Syawz/EvwR0QP6wVnl+
IpT4BzfxJFMMiL3U75n6sZDj3tHW6TYXHXpePChFOPl08jir648J2Gc3ddCUrFTz5RLbUIPxea8a
JOkpQp0ZUCDdeRXRpZk2S2+gU2R3lPKTQjEVgvgnMRa4HUq9QKRYXRycCq2dV7XRg/BIETzNu2do
EvryOO2VPLTid49Rbl0IwLmmEwklHPhIpdGlU4vZzonbcizyygKLont6lcALsrKZmfR5tMU4A39J
NoEirDHEljxe/EOeN2rxAr7WzCRK8bg0j+qrj7kuU/C2nTjb/gpAeBzGRIY8DvJ7pxsA0YSpm4Mj
JZ0P9BWnc9IDeU0tbmGO0K9mqYOTiBHQ7FPCeQhnT4s9o/yZZh9e8n73xOMewsfBfPU7WvLexeff
j0nGonakLRRynN7RezLWTzrogRGe2/lHsNYjSBKVenz5rdFHuTLk5SApraRWTJHS3aB3iz3bP1OU
MRt/NvEHznUWjl5UAf0bav+rhqwC7ZAIwh7RAnRrbmqsXr+jDq6yVXx8vR0vIaDpST15iSWJZe3M
P7Wmv2BBqF7WVYSeliOZdeuf06M3lXBYUc3vFBpComl1mxVqcbfv4ftZVLusZMHb+KBimdwZgZu3
F1OtmkXXz+F82i1YcUTLWHeli7QiKjrZhAQH90DVW4fVja9tiFhDRdJW/I5AyLeBWIsue6ZFtHLm
VM2OKW/C77hJRQMLVluCgE6o3TQGUKBNMq6rZ3tMUYSjC/thmGmzWoL49f8BZJusMONzGS7JUHvY
rdQOGcp5DMNRmj2979dLGZnXATr1vwrzSMZaHGdAsapnpmjHPC6Y4Qg6YaXEjKI06IYoF9h/MCS0
M4RF1gZHhOeOyW9onF4Kz18/cQMpePpRbFhKEqZ0EEvU50HImur1MDhpZbXRay9YJAFZOp80z3kY
w3eTySsbCWNTV5YBkpqKJuixlSnnYceHajMTke2CX9HBtV1l7LbzAvmiXxvG8Eti9xzxGMJIuoqX
4Fsm8ZMpdGCjfqNpfA6W9Dz4ObM2JUUUCXj4eeh27BBuvVnGhgiOKbW5avPBDc+upMUNJmvVTn8E
OIDZU1hDHquNQU4Cf2l2mHL1pzVPC7uxw8bS5LmL8+xeGZm87PBG3m2qU/hKGuqycBEOyPC9q0EX
IvPecB7D3gOiwFPz2N6K4/E48fXJ9Z7FUzRE4/ngVnGbE2wRAeRzudP9dpwB7N8OGRe+84SmYNMo
uTUjHYHQ0AB95HNDMN4PIqtWuh2Qjmq/a5tPJc6zHRHL5ns/n41QVwxHXG2gf3tLAq8zoFlGIVYs
n/NqSSPxUQ/6rADyUq/5xDpcNBWlM2lhHQQPsQ9e6R5kpndZcf0GeojPxWKbKI9FmBd+JJejBD/T
xfNebS/V9Vizs28EUaZQWJDg3uBmNGWAT9+QeIsfkmZhZmIHG28T1zsbSYrzZ0qbfPCgVc95QbZc
HtJjqbYn9exE4B7njyA3vkCyOpwf8EirLh4vwPigWQs12Ub1+MAmn+FUdgVsKbKjstFf6t8A6BVJ
t8q5Gxep1VBhAG2xtTxLQgNYGIgVIJwLGDCEfdM/lgpvLpV49f1KZJWGHRZu+Z6otPQQWeUgNJDw
RjOZpmxMECeo5gr9SUVmhYp77wjz8wzdD0QwAQ3pNWObDFbfIZBFBPoTIA088PBVYYW9yWSXZcoj
QbJBe40cgVc000T0X3rBru7YSk9e7WdlUbFb2TfVjtiEqNqDFINte7192m5jAxrS9Gntfe6QhT21
t/SlUuBcWeRSGv0c7DbtAmGYZgkqKN81IpeEtCYAtRH1wt78bjjfSkIVilDdjFdg7Hqk0l+GWm+2
CyjqrjX62jsjdxl5aZgMuzfmV1xxaZOrB7Pfhnt6/+8SeJPJJ8tbsiEuI5zMKvMbCvdzzprylimw
EpXk7ROwT0G2DBtD/xBmh6CUkH/DHaeM8ibBOynd0O/8Hq+wwkwQvRVdcV+KHK319cGPFbj4Rkdu
+Oiz356JopkiJhtDO9WdfBBb3/gYl1xo4ycAmyP4fX5iHRhuDlweVh5y51E4rO9p7j0NqWfTwLWG
6OleF46/F/JTjFeJx9sgNQgi5Gvtglz/B14vsv4qswwaNDIm8St7iT/9HPcH3llGZULWtTprkxW3
YFPBqKNg+wvN9PScPhsKNlBQu3KoMX59qUGeyru9NCwv8jX5zv/Dj0RNEhHuVSz1HM/xhW340PLa
KABQ9Nnyv9g+W7U+sIa+TMj9hV9U2P0sJz+9lUFp4suiRZ8Gz+tJaRoI9Gj2BIWUZhfakvGrETON
ic//rug37FATNF1cli3gat8ATKvjvE+kHQsVVRx+WeQ2i8T808oX6QnBzTYvySEP5f3B1HM2d8an
rtRu32IJZKywPEfp/MGNq7Rd/VrHruasOsclEwdW4FnIqhimXtTz/sPLF/vf7jX1+U115GfnWmM3
IV5+vL6EK3x47Cl83JExcIkgJDuNLrM0GrVrs2tppHssEby1D7Xlz5VIh+Msb3VPHdMLdCmLjUVB
x08Wv3DnPvPQjyJzICuLbmpC5lQedIKXg91QDrChsh7m2mRbB1eir8ogwpFaLaOJcT+TmnnOXO/v
6W7QCXPAa9ieA8o5yOBGIJRHLTCL7C1rLXT2wrFqONzcZrBThroLU+m4nltK+hzZmiKM1sz/QHdv
/E4vkewXECatyn98QXMZO5I/gazx7KulcEH3PSgwSkpQbgTpQdlu/iqn3iBIvVUZVxkXbyUlbgGu
ISMh7vQIW0W+t/c6L6QuyKVBfUYGolFMKRQ9TIjVYaV+UQAIyZXA3Dr70+i+8e01dIYddsNQ85Xk
hW42HuutI9tfFbp3A0SBme1O+diPq0NZ6cvL53WWRDwGTRuCvKyQp7R8FbxoDhjeykEM5ZCuoq3a
IlthWqptm3k4TibPCwoCUryclUi/7xF4XpHBw5V2FKukvRvkekUMBICI4m7MGo4kYk5FdWdfrQD9
CFYE0o4Eh8qdn5Kt/6bx5LfFmnY5NB3LaAFbeW6JokYnQXoVxpMNM3puTr90zYp6MjJmq/sZyeF5
4U1swfg5JG7/L+XsGWeBozAnNFi5nqMNs25+/4bglZcME48ZEnkyZlxfVIDbq1RNmG5dR8Tp628e
XkPT5iDQm/F7OxjOb7EJJJgirKO2LiHgJf5Eu04A7xDM1niquwEPlo6W0e8posTjO0wU6m2q+T7G
gi+evXIUa3tUkPH4iPv11m3paf4EVzlXIG1zHajvjkZ+SEUM1NRYmdV6FfjXAVRNUUKohWyqg6XX
r/6lqquAe/v3+XO28C+J22Yw3+mugvS4iaFADb/e6Nj2fGHGim1dMKrhZB16KVqO0eHH4u5i8ZIz
UTPD9kCDMAPcS0XGyelf46DyVLpmWEy4WYUjNOC9MtwueBvh+3GjAa/4A2v1CuL6eYXWxhEbtBGk
FnHoShut661ZmRXhD8+9uNm/zPWRF2Dtp4CdOVcWXdhiihl94Jl8kWKG9ppf82205sjcRYYNkMXL
8Hr+0I1+nSv1gn4qBaiY0PGs/YBle0B0rJ9IC+WKw+t1sl10TLM/nsOEmQoYV6w7kIaB2sjTPosx
S19iNAdd+9gvQNCX4r4lcVrMk+cyVrNb2IEbrz7THs38fLODRBM62pYQQil/FI/7L+5mQ/Fxt17t
D34Mv6lq4kWwk9NvwBdiiW9XWfC0HWUqvLJnM5vWWirZceMZzGO4u02XHrLp+Rz0n/yzS+5mpW3c
tiJ8CUynz20T/6vtp54vKRuOO/lYAYwrLZXyrbu5kfBP0jBwrcHvaNc3ubNzs5CLDFOmsIkFMpN3
yI/z5ae8yHFKycVhdqo5SHxPGTdqiwF1B7QwFKomIJ4QlWoNYWeJdkgByQyaVC0n9mzQ8GQ6sOar
59TZqdeBOvfXE9TH3DLQqRsT1XQtP8lQEvg6ypDVsQTer1laLlzJDkXhHQ35ZYWIq9mEmJmwTr1u
G9rYe9SmeLrRrZ/4v7yqlqBrKJjpmjKISZxCKEPoCdJoqICU5zZPbkv29L8d9qWDy543wA5jMm+3
UrXkehSSSj1YxU4vEjY/eEjDtCeqKFor+U3rvIRS8zwyoXhvuyNAQjy1e3TlYYE+r0+6nz7zFWgt
PjjHUe7zzbTwnanKzUpVwiSyRN2mumVaztmJK/7U6GSvIHkWPUEv8r5w4Y1jhdCo1lTYonXJcka5
sspbyeJkt+KjQjP92TKWTPuvnAjO9vMj+DIcIv06lXTfs63FnAtHQ9Sh7pQ0IGi0I8TGxIxx5aS0
tobPKRnCY01Orz4dGCzu2YNoFvcLYgoylktwxuc49hf1q92XzSSc82degVz7hvqdgvrRpXawtk4O
nD4m2IE1kbMFqgtkRhw/FR+HTP/SJxoivufjx479XZKisdT7wW2yAAopiW+xxE41Afl9YG7xXyRE
IO/E1zPodCJl/u1UgOK+U3JcTrkCkZ1vd0w6/bpEX8rLHaFwl1fA+cY69EvU/9EnKNOHAATt6xW3
PU+Qm9DrLVQoaeyCa82b5HW/JsnoLfGpiLSneYjj4jBERpgrLBYIcWp/VdxVEibHIX1gtBDPrCYY
Nj0rFJiDdMj5UBMp4+eE3NxX8EhzY0vkWQLFpphsKU27ig/c98m45y/tw/HrH3AluNAn1dPBG3Cu
rNqRSuX1p2zzV6I0TK26dIYOwOa/m5rBnnV70URHFPgVqbdbBV0zF+fLRePF993fdfdsxalBMPhk
omxvrvKcynBKiNQFT9c0qf6or3OR/smESlACx4C3eH8Q/Fn+dA6cOIzoQTdqp0AqoepBAjBSOVAd
1UQYszx3IyvnkrTXzDcT5YgKx5Hy+XBLR56Qop0wlsT/8WfSLg+VAbCObIHH+FhVG4XXLdW0lCON
0j4JiHL7sqyakshg88sxt2IFBDRlwYv9zXYTJ6j8AMz1+xKCZu+VUFzfl0oJzWrt/IC+98rO4/fJ
Rg8T3ikgd6DXL1ava/gYVqQZjLMc/mpktUWKq0pQ6z9OvRPcydl6CnfBhHYrLlDI4lizBc0A/7Um
fmhPAdVysZwXXC2fMrN4Z9IqFpBvcmMRof3vv9u5USK1lZ8eyf79WOPehAPbXsHv30hWZJFCgVz+
B+ikGPsoZnrGGtTNEv6V1ZjRBa9wf2zQhxUJLuM+isypc01yqSnUFQAQK22nQJtxTZn/fc125+ro
5oNF9wdlTcU1+N46NDyJnVcDpcjODvWO9Lk55nez0ZmR3r/NCAwqiThSoMdBTvkm0/QZvVFkVWRF
36aI8qosI2xxbwIko/eA4aW7f77TpMhit2Doe+O5qklXrEOLvvGdMMLwV85jmyjYTbzviIkk5z8R
nMQdrGji/kDmAlyOa1CYV/2stSp7kX3jCxCtegBk1am8gEvC72RMKQTElCqZez/bkhY+fglmUgVK
/lLg47xNNhKLY3LS8gwmJVxq6HgFmMjKgpwC9jU38AlL/Dl/NlJ5Hmmm3SgXVDi/acxn/LIrddza
/rZq+bCNMZXJFxOsj4HDKJwVUFflHWn5fvD3tzlVeVV8NeGkPJRLRUxVjIb0C/XbfVF4mn95NaMx
4u7i/DEMNLDXaPtyhStmkhy/jkZ4Qa9YDsZ/N7RK28N/+Atr9Hc7zJ9mkqRCANvwx77qhzXjiU6d
eaTCre+pK9Tomb9Gu3WMF0nSML/ct9RX6dwk1eL1f6jhMMEBED8lkSJo5l//sSlBjYzdhOk9Z4gT
clQBEA7hSmdy6u4hpnkGb6TL1/yjRUWMgmI7Nwy1QpU9TN1pbBfZWSidU3LY3Cg7cVtO3sVz+T0J
UdpKyyp/918n6DNqMZGmrB9GreGGlWb4Efz1dnICeO52PLMRoXfEKoxVqn7OwAJKliDK8j3ZMWmv
Bd91hYiUeJNvSo5voJzvqAogiXqbDCR/fOkqChpwEPhVLkE4yLVXzsh3erga0BgrPmWOnmvms4ln
7GcUz5AfIojyN8WFYslN9hPtLjBl9nmlzYbZDL8T1mUg1hJJstzaYvifR2u37jkaBqs2wojNNLId
zyV2ccCJiZ79Qc2U61MPhcEcas/uLXCgZeY20MSG5Nf/Srb7h++RHZ4WRybmTdsQy6BJMDL+cicI
aMJUQJcKdUsHlD6Py6o7HEYfBpG5bnYuzqwZfaEGCWtkwDCQnh3ZefQA7REtXfvyd8xj6RqbH0yF
CrT+r/Cy5PJTD8QvITgvDKK+5oPm3Bls4+RPVLqpSkI/GgsWxuhB2GDNr58XvUXnXftOPq/htuB8
LOUNFdYOB1gomOxVLKMbimsmuAcwJ2x2VS7V+z2m/lH565ZtzkLDSYVvoK/1C1sNGECy8PTwuhHE
7GwsUkbRSApgEhXV2CYB2PiLG1TkYmuFduKiHwkiWMVF0fmlsqOMzqra2EK7tKBB1sDPyk3bxMaD
Im8iQtw4iqZlEX1Ofi/NJn5FjO0nkiiyAP0QpgRxWpu7HZ0mPDC2e5gMScG25vOa5nFCt7vamrx2
FJ5OByN9fNR/fIFCQc8GcVqJtwGTSQgjOP1KWASEwP3kLPmkuoEAaltRe2ZYkhpPo+OCnYNwbuVY
/g+oh+RoboM7uOV+91ZFBz5BP4+JWBZf8K9X+DO6MYuyXOAxAcD6093uHGmz9h8R6ZPhJ1qoN1XG
f0zphoW7qEL9rB85UN+l2MvxEflcSOnqMUSczgwi9hls3D2I21qmd8WsLUhB0843Cjtny4g1ocZP
u+8zXCiqKVagVcfZrHnczmZ3WVqy2WoFROhx044fnnUUMxJp8hZpL+wBtgvJO2mOxZRKrfh3I6tC
D1imyBQvUjQBtMYfkr8/6fa3UdVkHTqCSpcFHQ7k+XCpW1bEZu1hVVKZQHKT0KvKtORjjhvzgtgm
BBKKpZst7TFzzJ14X+3ebC51aeooGY4GemG6/S8GZ1ojo4nKsrTlSVZOpNUfk/v7J+sxgpOf3N9N
Tr8PBKsQMFYTn88fRzAnNAFVq9n/N07cEk0dWOUVrZFyo3aYo8iw5AYIMMlMjjpWwqBDc77vbUKm
fKNwvr8VMZqY0fIskJLu5R4U3Ks2zx3nCptUcljLGzCTkBf3jaoDyikZTIdxpC4sAjikMVycPWPj
8lz2cASQWopx0AttNSPMK6FMtlq5BFe3/WojkEHfTOSE1FaesUjeYGGmX+ADm0tmLGJQ5LkMf/2u
ueIUYQp8qjEo2jVV44r3Ku8aTs4ZGKxKJG4vfbqbZQnW/IEEiN+WaXdORWlU9usiYUNa4914BkY4
2giScY5u3xlKc+FDcevHw6EGGZr+eSdSRi04H6SE4bS6SyCmiBYTiYGV6e8KFkEPDmG8OyHuh+0S
B22hMuvRKc2glHkxZXafuuJGs67B7f0reoCRqDhcMUjLqNVv3PPmb4lqiN61Gr2F7kOrer7F25ja
uYxyMUMQtSWJgmJ/mYrtRFk44Gvksc4Ztju2D3hL5d0g6J/+TrYU77WamlX56qrd9QqHgrULBFgg
koONwp5D6z0w86gPv0WLj7YcWoPlMrDHP1iQ4tdjMpnh9wCrTmDcdnthAvEHIlO8igkI25nHytqr
Him9BGrw4jdzAjTFZw8fr5rbGSICiXUx68U9hgMuYm1XPHZqGRmVslbhxAG2+CYIT0mQd3QEHei+
FaqhkdAIpjN8k6SUKz7bvGE3ppWkeuajWCxLlmBj3z8OPx57A1hRVcl2bRFDwyzjJBygSWZGrwu/
3W1eYyvzIIcKtGrZCIaoXICTcbP1kNeWpOldgvm8DgcOqw90IUqog6GNKHKbeMDdwGIUtAMQsgk/
CHspxA+v5dOkY4JdtnKPzl9I2LAPHvx7j5NTdu8w1hNECMkMa6g0AD9yyCgvhMQGSLlO9JOMsRNo
DnQNtG++8KOX6h1TLyRQjKIkdj5XfWg5OljMf0AEi+wfhOnE8UCCNyenbanl6S7AEo5oM5FaCP5Y
BzZWxUeskl9ETEqGfMrKD6fNPv0LCcJob55uT0o+SzRIfbZm4SWhPV0oetsv+Jg+RdUO3ESag9fO
mes/DAZDEtjkAmCdiZRXvagHtGoILQYgc/6CTaek3mYKO64OwDsgnbJ9SIJm8p83bhY4b+sPVjGV
S2F2m8FRztxCE2aaRgJPaMeqtULmQrnNoFegIjRzWT7Lr8slSzWv66PBy34wUkO5pTEPo9UbMmjy
n4JSch55IOqLVfZ/xDDBSZjbk/0fDCf6UzXkUkLXmTwdSgDQaCiD2KajsYRbEtQyT02O25kLBrtI
jux/0U+Sv/5bwhEO9uK3SFlwMyqwM76tR599DF4tj8C5N8O1b1PhvTi1uD0YnpPvXwB04UK5FMqY
3UcT8PmXgfdIBOwEDQ2UKXM1kvnAWG1SiuESpekR568iJxkkxi8ZHO9S9oIohUyHCpr9HxERAfiI
5ofB9JgUxI5QBI1MN0PDL3vBPhyQuZ+robtuRVTFgxgwAiktp3usClrBRgXWEQgv3ejdCP5cOkJz
0wmofoqjenM2z2r2mzeCiOyUB1M83EyGmtJBL6m9GL6qKEwosZ26CgsFz40koqS7eY3aQL7vigc1
s4NvEUHJ73pcg/sEQZMoEze6M8cK7esRi2eXVICVTx8UQ7MCaBvTwrZ3wCH329z1UTCpeCh2xwlJ
dUfOY5fAWoMLTkfxd/GlTDvmzpTaxxKlVglLqW+cwezSALPF97IcApoLtxgVnfS4F89yGlzMxSzk
FC5gN9tuisN0xsg/kP2y+DBqy8BFLi+OAkze3hC1Tt1DcRjyx6XGFM58BdoMPV6whtBBSJodT7uq
YbRfrJBpgnxFJXbAeeAnkQr94qNwBXx2TN5erVyrkir8MMrdXTkZ4h0Zw4KcH43OunCDTvrkI8kF
UR4THbIjKP6D5yLLG9e36iXd5f+ek2KPvmEBGAwKgnor/NQjiht575rVB45H0N1CiRWyyBuW6Bco
7HJjBTPVSTWa2c1ioBn7dB0C5ItLL+fuPHS2LsAY5uABVy0fyePlY2IIcuXMAJckcJ6xjSa1RCg2
6npJBqOg+AGeeWvfo9agY0pgIKxifUR+C5VQI7NO2Bj7e65xcKnl/BTYwaVH0GWa+S/mBAQKu+3C
rXi5hdN3IBYZB3EWDAXullTmB7WOfN9IwQJRYRgEDpoq32quoQEAg7/Pti6+/7Og7eMJVxuE3RrE
oZ8cUCyZBo9EYu002ZwV86CUtbTwZmU7kG3++VHmXwslKzLm+ebBOGGWez1w/Vl3+eOK9rAxLcpl
DF4RlZBFuvLLo+aMpsIsBdQ9CPZwn1obhdh5PAEOOk64v3v6pNxtQ9QZsnv4wuRiL0EouIswnIUQ
b2ZL5kDtTkTr5qCWDWAILbymupRJVPObCx2h71f91VVTOaharmqUWS6WYe4HzXpE8wq7tk5CSdqZ
FR1TGLj72kIr2rWWpXPo5hpo12qUJE8EaPtTiLvnbbbpVyyTwJLJfrxjHrtkK3kQKOFPVpNpBOu7
HRcantAmsor8HtQE9D6WJi6uZEgiWRaxQhUwb1o1rdkKpKXYFcuAZK6Oz4ddXyrKYQiWPC7YGvYE
AkBXYDdvzjqUQJ9eBOZj+6IE+c1B0ifSwdeMepvTHgsNjMwMjG0419PL0qumo4F3kD+3zpOrG37+
ePqIvoAmvW7a5eRt4U+NBH5IxVuXYqPxhyBLvFsAQRc9xZUA/+WdWgF4OE/xr6GYMYw66L8NvRDx
XMU/S8OjPNXaHlpZA3r9w9kxyIUZgLNlrp6ICKa8GQZdVhCF5g8e2KOqoYGICLHihzIpdSmaOuVw
naxXOafdQ7+B+bmyvQd7Bd0iumEhSnjZbNXRClFTEFh9Ap+MLuwS+6COR6KnTNxi2ojpQMUKXfdX
xialCirlqB5/6rR9IiURD5yVOt6faJZ319TlxsMqw9xhfzBT/EzYIrLn88ZEjzbssNPwYqc+Sgvb
Vy/jSdXm17S6sLbU/ceFAgRJZdNm2hgLAQpvWdmC6gnKQvSIyrNTDB32PzJ3OQt/ddn1IweRsNTB
wnmfMulDFsXVQJHNheHGDKhnOmx6fpV/g3x7gRWs+SbKuUULqiiDQfrpxJOKsOkIEf89kENvTn0W
ebx7r+VgBbjhAliX4UJdwYH5Uqh9xQvY4iXLSJFvbHdrcmGY648epdwe9qJtJFKe0IyKxC5vUKfI
5Lzp4tpXfj0eVHH57Ilxekd3rMswYo0EvFOzgsR/GipteyzfxPCsnCySVxJELMOGwlQchK8obOfk
LpqKm9Q2EaQK2NQUG8RLytaB4jdsmxsT1zxnWUaMFxnvI4sfZSLHtIrwXoOZaiEONLH4LwGVapaP
juVH42ibtc1qt4Lt2xkon/Dsym++pUQMlG/GChCzLipzSs4O4PIwJDe3hWJ4zLenADeJ1403bBMk
p1dYT9Pu5NPCVzRoZlqMa2OEesC5TnxKnCr2mLkQ/z7fFQ/U6ltw4mjRlX8ypaHwJDHr01r9IbZB
yBeLQasg8INBlsc5HMndbq6y1bhL59r4heaNRlL8t0CgZYYmdsZl5b/4bq7/YhBV4moiRjX7KvfD
23Bc9zZihP/ucuccJ7I3bHeRstcDmNA0xcaZrwHMkZVSNt66gXtIIrA63UMy+NDkvJelvfPYCTtW
MZtya9sbJK9Aqoo112e6Iu9s/zb45d5KEtDhrylRQq6po/bxArCPWiCSF/bUhH3y9Yss1rMKGtgH
1dJmOLu1t80QgYWFJDuVfyE/PGZiUuY4Y24mB7F5zFUzTblYtREsz5qGahIf/l/X1WzS5mg98u+s
wPzscZcMJPuzhvnSd86/MFduDKD0hvluIV3q/HJ84iOPeOkwEHTzLwW08HIf2YKnLWCBnUWqSfQb
46EZkZbYZN1SA4/HXJd0Y2UeGZ0Dj6T6lwbPC5X+E5JwQLuzQv7861zNAZh4xrOHJZ5qX7iT1zgz
flW7y59a5qF1EfQLF0O4rpbOJeLToA+56dWjrz+rBGTEppNtN0pQtdMONQkRRCLfp4Fw1Vjyd2I4
lKoXMEji8ilLIm6D7yopgGz3ARmWBn6TNzfrfeP6O2tA+hqLZ/zXCEaS9LZdYqOjZI0vuNF+HXz1
fWpT+r6epujY8L3qCREOUmnGUWZeJThUvTFYhHM9krWZ80+Ai0j2ILIANX6xtHBxLAgsE0GT/N8W
DBpr1K9QALPBMJBSdrgl1EUV2g9nx6wQFNNZuOxQrA4G8S/5UY2w1BJXmnTBJ5LETQAl0puM/lD4
XMfl8DVzvLWl5NhpmNnSebS3qXpRYyz+Z56IZEOnc6ovnc1yN5D5XklcaDexpp6iNjH0KOKtp7NC
TMvf93PBdkHCY2VZv/flDCLTLbiK+fhF+5v32oZiLWmC0jpQ7kesIt4LdgI59Gg11/AuybBQByY2
H4RglqSE1kLSgou0Ps8iphcB0dX/kt5eq0Q4NheqhAdFMTbMwekxIrZcY1TGk1FoIZX4OoSvMSJ0
E3rmRCtSCgHxjhENxe6NO380VjgoGaIN2xpLgbOolg0OMwmJQDJDdESAMU1Tr6DbJpcoSU/av507
+kT8hx8xgNCe/QwXrIUSwRDIyF9fQoRjAPl3o/kJGd/wRrRNJHucWPKzEgsUM/wqSmMkT7Bg/ljw
3psrZ22oKfKtrs1diuiIQDzJDy8P0OGgIDGOayufmAJGwoi/Tel2NqRFFdKMC0asQQcxTJqASIK+
OiEx3upnl9dG7HmRdOreZ208NI5k+Nr4XnjuZeexy+4AK8AhYGnfAGIb3TUSCQodVRqSlkxy2YlH
XZqK147nDzRX1g0sic+WwgzH9EneMxZtJkDJzrhYYBS3A/Wa5PBTjrLFxYZauDiUxOr97FPzqSLP
w6RxxBX0yz0vM3SHtl06vKkUBYyAK6iQnGXPpLf94SJQ4RhfrCYWYNdFwyVV44DDrd7tnf5nqak7
8kAloj0adhpkCdCfhnjdAsOZ1OKQv3Q/iIdD2QUt2ASNRKgsufcw5qcYbmCICPbvdvqin9fkERbQ
EWYM9nVER3vtjf3BT/1wB7EMXkAciEwRUKulwIXaPkmyn8shYX6mdlUglv1LVm6ZJRlPOvDn8VOu
Wt7RG7fATBUwMX/9z0vnXLN9ZXT9Uji1OmcOvxOMaXrQMI71cUxdMsoUXVGHK3csOBmH7O6J0Cua
H/LtD8BDg5Ij9R1JjAJFkJmnaTHWEY+QGGw6WOn5tfjCMRFoxEOm0sfOal8GJqL0JChBjElwnqmo
lLLaVl3o3WrG4QeAoqIXQQ4mbQo7uyw2PplN4wjY1QxejTUACJIExNXfcLh9NDJ+md6nZCgEC5Fq
VqRDktMl8IOpajgoTzL/QEw31QBQbqzcj6drVA1twF3wJYtgve3Ghhos5Cm0IlsVGsc09f04Bxba
WfruCq4lS3fwf4Dw6SJuCIXGMuXzdDO+KxrjlH+WEU+TW2bcFG10EnBFldjFtAbS6vlPrHuoYN0q
KRPuVHxC6umx2iRCLmyuI59JkZZdjVlOAOpdT19IUcxtNqgqO6Gov3I7yXHyApU1E1kKlzPNV8Ag
+tloK1VZYto0IFRmjp65vc5hvPDwV7riRDrnj3Dw7TJOjOtIUoKjAW6f8bkrbe8iFD3xFhx589Lf
oNHwDH0lrhIIz3Q0gNW+Z9lcZaJBumkVmlna3dCB07nmtE8ypnrbF1vG0lLUbNjwJmzlaYwOsm1Q
qEb9zkGfb6oAAqitoS+EXJR+D/hDt98A4zU3/sS00BbM4Mctxmt0cP6zpXSr0kgZHMd5aZ4d6Rul
O0O6u9CCBuZj1C6CjEaIepawV5JUD4HI1MGKLcCnZeNy7VgLSh7Od57kmL89EUTo9jSP+N5tqJS+
ZEkGUonDASwdbfM6+Du78PKRZ0fbhdGSALizZude0ywj3YRp5xUzErinxvz0ArLMPT/ROG7v+2WC
RmUR16O8J3rx01MRrXtZbPGzEOn2LacsQA/5MDP8K8/QbOuyAK37VpM35I0aJWGomK3hEKLgTgyo
+q0CYlTv6DqDY3ygMV+LmKK+c8+EnI+N7U6058UFIGMHuHGdS7ZBg2fVMsHxY67K9+alMhxfXN7P
o5dxno/ljFezeRGMjJV6/vj6q/+NJx/vfIqxpD5C6Ha6ABap5xwOBr4WbPEfLnfIV6/eJZGMA9Df
Nvyx8GNyBqGTNfgRbGyyXZuDGQY3j8fYZbt6frL6U6AlqDlPD3TByHxOZ1IplXgP1a1plpMRj7XI
G+IX2/TuXL95pvHAnnLtti2hiw/C62D1a7HEcJ82vdpMPvfk83JH72rnnesNrOEv8E99n+FXOfUw
qiysd/RBdPWjCon4vgpszngMFhYOOsrjISQYsbzgvp0XII0ByZ4pQv9Lr1FDG+lb7ep/2u1U2eMl
+50Y2uSnepvaBl9yGnEcEEtkNTUiafHLELzKgCfi8hvzJt++O0hF+YYXAhziI0KlN6J6bdrRaULh
wfDCmj19psGCnHQ/XMXlwLG+LmzP2M7coSKwGgoZJthYvsHF5dHni3Tt2YysKDjXP/t7YMsPhE8w
uM2KGMlgRgK/CYC6L6CvJcgxub+HlzGbqMYfRzL/9GKX2vNpAmnxAVaKG6MBhicLf7OE2X8lU+vW
P15KnuB7wLI5t3GsbU/6NksQzotsFl/dX0gD4a7wLGmnAVAhaxK5SEVN7eQ+csWmV0Qj2e3WU2ZK
IyuPcmwWwKEMfhyAq/0IxL2pNknbBZXmjdBBb9ceYIFm4s8RbX43zG+eUQJcfpQ2l9K0y6WWE7YA
STz1ZTTUf5/2v10CaC9mEZHtKej8Kq/ra6rKV/kpHgiok2Ztk67z5phwUPK0Yj/5MUeTnkTaHkrK
gTiaGU9VV0K4CqDwoJnObAJBo+5xvuOAijd/Q6Hl1ntdAkR28XUWW6doreoT4uVPDoO2YF7vMjKy
hd56JDOEy1WQuTQUehIYeWGXqh/OqGJNLDE3crxTK8SugekxFeXLWt5m3ncd1o49o+8dQfT92ORH
3iKyoPkEYFqnDip+dvW2dqOogcophNbyjFwjzAtkNr4WSKmkqlT0HkLinQmRCX9NuVQ6b8VR4jVz
444aJdWQPDiNxNhI4+P/FNuzj71c3ebPPqhDzkpKryR2zsfWjGqtF7bPaHVAVMTm1mxB4sOv1LLG
N3mI2mV2OO1EWDlcEGtrYrkwvM5vZAlGxT3Q1sLm1F714Cc8hrI9mkaTLz+z/p/oXa92QYAp7acr
uNcBt9kIUhqm4OwS08Rhdl5e5f+8rwRXxkHK/75sFNpLIO5kWcIdiRWEnzUf0HK4p1AOp6GcVgtC
xIw0yiEh9X3NWamVUlBQiiUpZA+BcerSMKWVYp1DMnscq0Kt36N1m6Q5J9TWzw6KsmWB1uM228+Q
MYMxnA6dFnCRsVOS06usfrzEO0KnuNuRquYV08+UhL6RLq3LHnDZDEdGRYq7QQEVgursT4u0JiOa
YXv9Ft89rgpccxHzHKvqmTKh0wVHD5kbV38vsJNXiv0TTbIXr73uu4FlwgniEqf0X1HGZQM556/S
+e+fGr8Rp13nthD7l3j6IfDuUQlhfOjuZNKk74DxpV6fzqnxxdqsABScG1O305MnnhzBXXk/pSfY
3rPnYOQTJq0GyAwtwuMbTQMeC1kbja1PS0qXaGGGcmiiNCE5+3GFDCSzg8Kr9UdglVxbhhPBVVD7
Xrxsh/IHzzCJ18kwRshTuvwFkeHfwyqw9sdTniqg3k3sJoo81Xxykd+ueKqTbNxRuofzPJDNaLxf
2mOntC483bCguwk6LCqh/XaqpsJmc+aX9YaOxIAgI0SPTj9meOYY5QQbPe/KpfP320HjgE4JyQ1u
8FwUz4qUFwyJfbq5JUT8h8+q5532I0TAvKHp4o+uj2tR5Ee9L+1pOd+w60eb6tlv9oA9bUfnVha0
RrJLdf2vxLo/YPqMpWI4xCG25BYwtsgjI40u2WfNcLWzu9RHEreijOVV10MlKMVLDdtpoHPAxOlJ
YGOxg4gZLziJ7DjF+fnfQwDfb+keiqVrNKG5IRBgpOuuwkdiLZakwbqk0AGAmVBtxId1yQurepd0
ODaelu/HiKujN2s0KftKP6uZ+3w55ZlS9o6maXWhuNHQHohwMX9f5YcRs9yxITHqjwcamKRORfpw
biO0sQLFSFxwKXzPnTMoDxXFQxq2+nOJtRXo862P5IRA2L1f6Lpjv/WkLNu4yh0cWRMbg+QZu4hd
wIzgIdiz3VZ1LJ9WfFu92bql2jOrenS/6+8EGkUGbFNWd+Nlw+3RgnKAB/J1UfMMJOWRFQLQWVqf
QZpGOs3TMgt9z84DVZJV+iGdw3F7PMp8LeD98BbcRmplUFYPs//dy/c6pgoDvLgfDitypGXxCkSg
4VdRQf+ONG5gKSEZaxd92yCo0Re+GoNMYfEQa8iF5V3HK7+HX11HE8Ni7Gi7/2JnG14v3bAvIQEJ
RpOCkHuTbfPKBdlSzHaNx4jc1K5FsvLGFkJTuiuM8tNCmgfxDgmJqqUSLeXFJJTRisLRcZpiQrJI
ZDzGJziJh+xuVlCW9V5ceisCGKn6nCUk+xeSz4tU/YKmT1akztagcJkFsx3flQWv9t+OlwqrPAly
oEaGc8U/hsMLbZwzlzZSU7UHtsUJZqchNebIx7ChQ6sp53oTJ9bP82m4EUC15vCi3JNd8bkgyoOp
BEXA8g58XN5X980IM+6x/1zEVqL7glBNp+eyqCrLkc5OFA0uuKbkq6bXK7uGCQTqmDL3iYpbJibw
8dv1NLedykVTnoVdQ7V/mfvbvmsAdB8EiXTEZ0bm/a94UH+U4jB1PRqHYdX6Ps69J0KA+9Y4XyTI
DcBrnluKRDCDEGU1gozoJ0fHrWzQpXWrFnzSfXal1Fc46rHX4j8/60CBq4XW0xgMAdgIYksoT8WZ
0kHqpPs7A5UlNjAPOtK4qaVi6ZnKPeBoNKO1P5xm6Adq5IVbMjm9RsxpE3P0IaRjXnyuCVG0VNVX
HUCFBRO84XlK9TFbhPe6Vi2MiH4HhGB3OC5Nlc8WOBOSTE090BcohZ/6i9+RQ8leFhYltdkTu8Ic
0YlaCT8rhhrVbevJp2WvrXKm7yqofGW7vnRYftx68+8a/wosVI47+UN5GrUcJDfi4kTsK3c1AAbf
eOyxjvlyU5c6+up/3cd/d0T6/J+2nsVAQ7WgLN97FyODioEPYrXTrXwAYs/RqVVlCYjFlP2OD8I2
fX1HNVXxO10Fx6ILiNsGdSsvPPs4KYuTOVr/dgNkNivLRKST4bsVz/Zprt6SXKcYKMrOzufzByJO
0Q1TWDLjEUq6OfEKzsy9FGNGcT+g6vdFzYbKNRS5Ar4kHT/kyyN9TeVPqnO9w33T81/0pscsrYbZ
/K+MiBaLf0pYv5ofX0tvers4hRje/LRlS8SYPmu8I7JxCuR/ZmiLgzBOFFW3Kj6jYi+G5neegWrG
sfYtuaiNCkJjeG6cMqCwrE7UT/Y8d4bFYsAbK0sU6JksRwt6BTcaqylwJBJlRetg6hKNEnOK14Qh
m3Wni40++4HBiFlLnX8mytY8z4LDL6+dNPEskRr6hjRwEgVLQZrey/T9WR6lTZETYcfym4CPSBtF
CHexWWstlooJ7hpeMyi2mrNhM2Z2HY4nzQicCsnFX+eR+ClyMOJqY14aqdM49zE3Ll4VX3d2864x
k0WOTUXOuNJPKRpRPTwRF3h7RUlNtpMXE8npS7CP6+F3Oakky1Jyr8grt9pqjVzjAt8WtC4a/eL/
BRrQmUDjvuPQpybN+9900w+1EvP3xTy3xpqFNRrB6HMVy/8PDSI4lk3WwXcjTSRG4tczbfcD2Wph
vk0oRR9OMHDGsSiZ84uD9VbQ+DvDe2344YYlmjzu/U7wjvgz7XXpHzVS1AehKC+lYKp6izNv+yAu
UjEGBF3pbUVCuSrxytrBtWhNr/EgaCSz+5lK95qpqJ8dcRfLL5Vw52YyDs5ntML0SukyT4mCh2At
DREja2IgVXC1vUKcAVQmzbOKFJkd7OCWPliq7nbMAQUWaBqAbuvPOJnCf+afSdl+Bhom7RcWnVWf
kk5jEmFrx7lXDf1m0//xqdWc4wa6UVfdVoNMWg5J9saOfSPBPMnUcoHo3I9AWql6SMI+GjtGkDm9
JJbOP5N7LaxidLtL0/4AsLP4LiM1HNyoyw0Jk+yH71/hggNvQSQzEgPg8YI4Nh3CCc+4qOZCvpHC
WfqiBXfMO9fhVjDXHkjRgvHMN+1SJXTt7brdwvztor1M4TQj34B/4RI8xdO3zehGysWFuSy9Rq6E
tOGtLUbcTk/p6cr5JcMtyhPrdMloOHfsXjb8y4Eo6In+hjKTf2Py/GFop6nUrDNwwH4RZ426MJ56
ddRm7TRfhpZlZ596G9nGrHD8ytoKZpFXuG77FsIt3muTN8zySyq2w8+YQza1kDRI23qCfazGpljo
o1H5+6YXwIojuGNIhFYkQEdQf3uj5kuXelSJUVNkaJF8ChD3W2e+fcrMaaoLWg6gPwktLCiLrJat
9jFDy2iXn5m1PuCcB1JfaFo+EUE4MWYz1uGRM5J9jHdkMH9SUeUApA4b1uwcW1xbVkTqMDhTvaYW
UUIf4rsWD5BeCWQ3r0h7zdm6C8skBfSC6xDyepWYMZ00q60OB4LmDwnYLuDvFALNK8qU5kmTiugO
wyWdws8WxY9Bx5xfsaLqnfW3fiW6clvV24ILUGcjAqJAVCUGxbkPOwke6pTCJCiKM0GMDm8/fw/j
9+9dQCLH2wmY2OZLsY0ZHO9gm9zTn+iWB34/JTB37JtfpGsFyzjDs5JCMZMymobhfsrZqDGypjBT
daFUVg2nD/bGY5yd2KyWd1EaFTYKV3A6kKHkoECm6po83LshA2zy1Tvnmd3AuPXn3nflZoCVtAJJ
09G0Q9z/hDh9dSwmyPCU2JDuA+slDT+X1AL0Vxhhdod80QXCjdewidfGZfPn91/FmhmT/QtfPEJi
lrP39l3NGsX5v35VLdsn8scgj4kIoArTX7Vj68z35x2EN19+bVLwrTCmdF4BEawuyz6Uv2IontA4
wvfj/u5f6SQDIXrOvjosP8ApettnMr0SQVoIsWAjDRLpvUQStdx8yMlWh3dhpuG3GHj3tBH62Y3z
Gbc1YzJcbNk3HEoUAAo6BP5dlAe9SJ014UBfLN9M+jOODudQm/+KrT8KSHSkMaH692XJ0RKbLNsN
Kqsn45Z10uzupYR3yJOWggCknQ8Xv0NnKgxItvSQLoLIWGneUyUHYfbmUaYvFqRGzZ6wXsr+rwhi
FvUorP9kvdcTV5H6AL2MiyOUYT2+e1ptNZRXgiTr6j8Q4Emt1pVOeG3aEcmg7YduYKGHFg0o455u
IVCRbf3FZ5n77T5wHgyoHPNnqsbt1AL04swPzqZxihZa3/WNsBlloqf409JyP3np6icB85kXdH7E
XmPZ/AEMnvmsYcRHnJLKlSglQoZOqvzBU7FFVBJTc1DRDDs5NJmlsQp0hzXEp4cpaOSeU1gfUBFK
bjSiyq4/hD+8GzVG3JJQD4Z1evnTBZS85T3+2BJHpheIv0BuVkGeeCSBei+mMjT+o/1vKYiC2eQB
3aSAAxHwSnN1EGrlGR0pEmksXntGXBlqnJGRpjTyCU1fA1CqSRUKmK0kkVclBOfwJZrWRBCm1BSq
Wwf5ggtFt7g6TDJRE+h5D1z8ncK2DbxPpMxmtViqBERZFof6N/YEDfdMHuPKqzdRuG5SYECllBR0
+8du39E5HLopr/5LrxNzrK88H8Ra2N4MddNNasTvGBOr/ShP3O1YJqf8wd7bZKl4w8SbFqusbJxZ
ThGIY9SLG1mjgbHhyh6WUN2orXIaXjSd0O2/jbvhflvcjBgh7iQcKk6Q2VlNUXA5BI2jQSljhn8j
6n2jLqZ/gXMYNI7BYqItFC/4eWGdff2aQfyHBCKUod4H62fjAOYY5b4wWkiM9SbeQVI8MMlC8F97
DSWbZ1GnfeBRxo6gr6N87faJlg1kvWWUPxWHGxyZYKnD5UG8uoUuGYjwv1sbV0bybNrVNVKXtKGJ
5PVdivBa9tBhU3gS6X6KBRGJhcpH5wpgul2/beCbXLV4IJd6jWDsk1+4F6oquIXnY3K5dVUx8V0j
Cw3ckbXd4+gFgpskBQYHOpJclda3iq7d8/PPN5fivnpZUaqnGux9eLp35QBjlr5Er8J3Sv6Xtdnn
Ki7H8XirkITU0ROetqL9Qhh1gcOxK4CjKjHObVx2jt9ZeWpxmsfqRJqVAY+9prKwBLnbxVBswfXc
IhSeOXVF1RkE9zK1P4MotCc7opBSjQcb7ez+8u9JhJlrCclaoB4ZX5FKgz5BjGdYyy0T58JPAj+v
A9oFKQMy7ERE6cwKyJ9ojDKmoTppxxBbeBibTC+xEzJgSI2TOewlkKuXXo/WP63RYVBWM/4NORJt
Nm/FpTlfNJaqEetUOSYOdWoxY4OVhe9Y08w9auaeuCEVzaxoiSyVU210Yu6mbKKl1mzl8fXWS5Cb
jTObDR5xU6QAA6zsEkBNomAO8BWD2L46rrZp1qRxg3CZC5SxmXrWDy628YonhjNxs4KxiUs0GnmB
iCQf7Q0TA1lamC3gGq33CmTwAglmx7zG3sw9EPEccEqdee0bMEdSNB+FjumVgkCtZcmHtcvLoQPm
X1wnRO8r0qXNgoxb6kLw/G4fWeH/TckyGCwhuhTOU/IGXWoIwDh+b1AH85MIjbhCjOp3f19NmQqT
TjYhXJ2HjnIdpGT6lGU7pl9w7jUX2S3fYN4sk/Bso8Qd9z53Uh41j/S/3CoANRWPDLMG7MGokXSw
UUDknWEDIRQ5/ScpfhFCX8UdIDEPPiL5DKlJKWKsjsr6vsiXXNR8D0ybqnvd4M28+IoT2Qc94wJJ
UPhQYuuWmNFMvAgt53BzMBdBMKNrIs+oG8bIzQTwBLrtuJD0p5jw/VJ/jIbbR+SbZfhNv/zLoNDi
6YI8bd7pFvGXFGsu5EcOQwjWzoFUhIRjEwZhwQJgBDqrFaJv8bfj8xIpp0+/Y0AdG4oP1lZPmbJp
pnTglhz3Mc44nNO8v9LSPCAOBpj0+XNubKVJ5/sUS3tFulYJjSq7D8ARTiN1FmCMeo+QINCRp7Iu
LSwMzpHkCqAG97zsQUJ+WKSyAHA3D692hzsO7xRpetE5sd05T4itXkTVOEIYVHeo6NrqOlHLNUKA
PXCQR/6PGO2jKhFAunopnd0XHMBcmBmU/OkHMP4Mcfk8xpsu3vFg4yAf8I2kdgBMTpHDB1BWwuJh
knT4EWS/5nwcGgIn2ZqoQGDJX4PjtYpsye6+p4vqp0qlNkHrPrwdONYaumTI4ViT9cqM7Aae+hKa
M6OrYK4UEaeJA2b3JKgOZB2tk4hAU4wXys7/jljUQI3ZXBzJE/oypEtciNY7L5RUBo3VhCtQ+7tG
zai6o5vn1UoR7WPorq3dfqCFRf7Ww1Vg34zZdZNvlHYz0xOd9JoWsSunawZQfnbSFHMGo6E8XNEv
c/68C86LccBAJ+gMNdMM9IDSw4PExWSNRIbXz+WwagUMcfU6QRT60DiiAgUjkXlRg86cFR6X8ZEu
h7Ki4jyufzdUs6ixll9ZquthD4YbNemfjilF0OTwKgBXT7j+8Lv8Co1B/1Q5X5Hs5uMKLbFhSqPP
6HhZwsYZru7yoQoruEmO5k/+5udmPnxoc6Duu1yevfOCcasMps+c01I5iumqP0S/H0HtCTXjeQm/
yNPWdqSDq8DrUFBcQ5rRK/i1s8s472pEtxzxPWorQADmCBORnG8YfsALm9uwPFDTKtIpnnSFRh1R
gPwvHP8y6KwiaD2mhYxwOfYmU6sQrevGxPLE5/KBjECVsFRAFOr48grhtDj3Fkn4IXSbZyKL1kKh
dlurQfcx61kEqy9pgVfF+ujxWOtA9caI+8GuBDJ4IRNMOf5G4ff3PNZBH8Biu1v27GIwRiOvGcaU
mqwop7xRlLunMQ/4BA8BGYf+P4yTAOaC3lOiUnOORW3b3aCJu8Lsm2+3MBxp/45Ud0vhoATso7Nz
SUqoS3/HA8KKtGWdytZgSKtnvE4q9guOzu/ZP4BU+5ZqsOpK8w8WErJBM4PkLwucCFBgnpaw7rsR
0Qx8H7kEqKJOQl5aiDW1Ye8w/OPxQK1QdLdAi3C2KP7Ocwfcsq6jcbKkg5gL5iGjx+uon0JS05Q/
Gt/tUxlNOkbvtFfBWM9GIQ2AQlKmMOAF8rdv4E5wX5tcbmM9fQDyUV0AfDlfjGgpH3tVPG9mcM7M
7zCEYwMq6jHNXNPlbm7P/WFDSMiexjv/VnYk7awmjD6L/HcPhQlJRdaEXgNMf9I9ddApXgLjWGCW
enM3riecGUq9fPXnQW7nk3zeG+eS7vxSI1VVdj8/c9WPEARPibhnqn2guzx+udUsb3zl5sPzK1LZ
+YJkCQISTk6epheRgD+yfb8OnsS/WPvLSXMTrvv59FzbJI5jQVHU/1YTs38PI2T8am4ZcbalZ17d
Oo4yC+z5in6HWWWMVq2vrBZmVCUuaiN6PSLwAFghI5+AA0hNejlUUaQ8BuwMVO8YAL6TCpo5bGRN
JCx4Mo/ynzhweVn0wHPPs5UNAdL3wU8qzR4L1DAEBHiCI7/FWLXfP1o9z4whkiYeeyGHS4BvSA3q
YkihGn5SodME/YnZmVMA68T73Bdx60Ya1uwOLP9Onot9IasUXjbOlyuqGt94KRZ2LELNUQPF2he0
K9seTpY+1ADZNsHWHNMyySdijUJDVks2Ww76bru8CbpjB+1nFm7RBWwF6eyMCCe+DRwl5n/J7daR
UPN3W5qx3sEU4vtuQewpzwE1WNCrrfBSrf/ehlS6Xh4VL0BW/DZ8FY0PWbJ1qeyI+V+JYcUjlYbP
ralH7SE1YfcNZikbrB985KWB6k56IUdbuf6nV0mRVUzpJsoCXIhPXFpums/pDlOmuZsaxhNR0M5A
vuiLrQRu20Ks/f4Z4W2tuPLwEYHu+8frQW0PmXccdRj7AxSlfeaZjv5l0SQSH/0ibadYfvXDlM7a
JHyE4dauWLt2Xgnba5oop4VTgHfNo7vtmF1MEO8pQ/NxG3JsRQGUdNksIpUuwwV4NDUrcHEUMmlb
Txbstc2FzeTXmlRAE4pv13ObxOsW6lCdWJ7viswvuFeY8C0ZLmiEBawhXASqOLQV1W4wr2kkkiPd
lZqdT56x8RJYtA6R3Iv9fQb0IdYsrxPXz3L4wcYrdxKvYrr3Uxr9eskH7wnptSvZRuIRtAwevVyi
c5znVFi3EXfCDrDXrgeAHT2aXN5LX3Vzso7UvL8YkapaawzIwHLJuS1RjgtUu6EQsht1L8cPQbwp
FMyXKV5u4vow+4TY+Ke6ftMJozjIWkvbJC312HomOLtvL4XCdW40Is07GnRiwKZhS4RVOHH10Zwt
YF+sc84Bvg7tAe3nQChmzgP2A4wWLniYK7qhEQzlCvvI8IoTp+C5Y4Er5roOvHOt1n14/OoekN0g
XbFsYcZT5FButhvnAdfBzStIIiK5Zxxd4tmLmxwi9gEkKfyFx/ERmh87j3xWIUaNdfb+n12L9VHA
ScWWiKX7Su9eJMLJg+ZlMPlwOwI5D3icI7XONTSh7O040W3z6RhlVFExsIXVEcd+6XXBkf0NwMj8
L87Ry2Cl+kwvD9D1TosdMJSpnnwbojr64Yy/xhLMGQmkC8l3inzRpOdQXo0i+BryGImjP4Br6LIj
W6DGAkxCTMqiXZiXC6MmuBD2uqOqTkhtqRaXIIVPzUw3PsUyyQG97suSjUWUWpzorYBSCKbNZciV
r+FpA1CeRdjeU8DI6CA5o8FIjg3ou/fKLXZLLNGGheJDyItosV33jG+SB2zeQGnjVBFFGq3Eq1TM
9JeM8Ae7awV9qu9jCh1VdWwgMkWc5OXwMlcLz5kDBFSBnJn71RoxanjSYw3diY1AtqMUQjMOdErH
yuCYEHinDtIOYNGNdFcB0KG3SSIPNXFpDkN4sF+M1MI0Q2zg5iYDG92WdqATN7M7ymeFabNqIx3l
M/GO0FSNnh9lwzdFzzG4kfZTvkBf3E//ZqmZjU6N/atGMC+4uAmuVdytD/alz2rvKjc1BrEvI4hF
sKvBfNwXAE/nu95zqUQGDtC0OAnpFtsPQLxVe3C15oDuwgkkhJPkjMkUknU8J5VF7kID4lv/ShGv
us0viOelSP7GWZG6aovHh8pAgpypRIdPc6zsMmuSThnQL9cIRuRLQj1pN1fUmGw7sh/y5FVKOu46
nxLEWzmEUBEMBSJU+S5iS35Y/dGxsfttrJkofxeQGtRjEwj603b/6j2EPwntFi197QbmbRr6KeBT
+k1kS/CeK1UwhqCzWf25U9Etx8/P/MRFkxn/FhMCUUTjVj7vnAMX4gneyEV6fu+Vd9TmvAsWSBVd
rROso4GRUruQ+edj+FPmBA9b+iOKqg0AqzAReZBdBrzRRCCO+ksZd0J49DCacmidjhRXQB7f7bct
cQECYxKat/ZqmBWYUMZk3lA9a0L2AYCKyWWIhDgcxFrYiTlBKl5E+s+SZazLjaBYgPWVq9DR8Wyb
L91EGpAyIvNxVqu9iu+iB9v4cqID+CGz/wryaU28tDJOes2dSiXMBqKqCVoI+9OV2tqNpY6YuzPt
01nRe0w57/BBXMDHodWtPzqmbt+Sv5mcLtdwM2vvyI7o39WZyJFEHsEtfMH4kx5GaM+YL+qb27NB
YLozpUzeUomy0plRoOhALhk6ri/h/qp6ZU8KL7NtTRm2uqDt5kweyZDNdF2PsmTT47hcHevtya/9
zEMNDYfjgct3SMhuC762jtK+BobSnQae6CnS+KK2+47QR9c+F7DDhEtZxqTZpAKSLjO8FtTlGcC0
qlZ54fQ5h3IjOkCwC8iZDJulN5W8IL69D/NL7LBdWRT85XR4XQsnUEP1Qaswuxk20iu7m4v5+ZHc
0cESTP0ON1piYdMTbroEz4p1dQLUdVdwoDAgT+eOuEGVENWYfUZYi5fLZN51+dqQyRI6GA9FNLRy
eBPYSTo0OchlJgvbt+05wtq+vRQpAqNrsQIg8wFU7zKwQ6CsZTqA3niX2zjA3kHyADZ498ocJ51T
02BlToYDwSZiXYW1nJ8sQVFQAM3J5yrLDwuX/yd4HgWKvDqFzYXIzjkBYuhFL1vdBizl1900fFEz
PcvpgvXa+b1s9Cksi6JMBKbFmdQ/qa1bJgF8sxACw80zQ1x24NCZvL9lgD6IMbVMoXElO5YO3Xoh
p83+0bq1kwKZFwo1grumGhcr7S/3aNrkqteBdBe3SyvVjGfihO7aNL1IvL/rVvZ+jA6B0tBeA+3a
kgmGVq4tIabjxMAMcuaoHFTZgP/KabrUcRD7bKWd8nrWh8TvfXkc0ppfyqR//yE5p6fu9Z7fL+NN
YIEvpQ1Uwtoy0RlLfTe7R/pKTQcfmFwnbtDkFRfIs9IK8apctOMMRqGIDSsWje9s2qP9fEOFM85q
5p5LdtxjoE4v/J1U02DZyrZfaL7kc0cO95WCzi26F74j9GrZKl+16uSSrYrV7kmrmgHgaJTRJxBZ
cEHHUgDcC2qkD1WOIrUY3+HU+SPajoKxxFpa4avoGAtIkAh5wgBp7YXp6ZssxYApmB/JOnxQ2wxY
ONdIVb/+Yz9GYf3qhgKSi44AQ7G1/ltFWSCZwhy5Tt4YzuF7G0GeO+ld3dWQkGU4zYaqVl9wj9vE
EcFIZpNjVLs641/qp+kDUb84bLVIJwWxYqI1ANV1QgoY5oxFi/QviOuTciPAeSjDAcLQvcg5Pp84
FaPoHTpLlszsnGlxv+OkM4eHsow0Loe8hjVS2g8/4vReTHBQH2IJ+QqtHu2TL9NRapnzO9N4Iy3o
bXkmcPM7FzD/ei6k4MuwxbK66D0MpMfnK3vbIjUpQcN1YFTDevV129/SmNFl40pgi28CTj6nkIdY
G08qxWSOwaUIHQaVZ8sYaPW+Sc0Nb7YURshgD90bm65h0jxVmTFHpKkXTAIR3WeG8T2/wGd4rW8v
Gm3xJEyaSnqPJdw1oXPNUESKAWRYyC+EiaYFx2g+LPp6pNPTPaiIHVA8URldfSdviC8b10X4D8cw
ntwc26NST507wfsrCe1Wujh1W3aB7OsWjDli2HkLbT/B88aO8H1sHT72TykFtWR4UdP4a0LFM/TY
EeFPMRT0ZbXw8AO91NjbMDi+52M8j18A8ImnbZDK7/LoN7V95togeKew1AM+7S2EoBlJf6JxjDZo
pgM4ornMFDX5q/odI3jKLxu6s+bDM/DYjxqumjaGHRkqZ7g7cr7wZ/j1+5yQ1xBcHFI+Zt+Ben12
7+cLCCK3k7OqnLcr4gsGl8taqqESd3bm6Vj7Wn8+ehEt0rjq0YSiiEItvaqR/pCmDdhjxxENyUmU
sTmxWdUD1BJcAlCKw9XV2j/u876JgPqCLn/M9hZbhviEBlRNmEnufJYUeUqX6kARfTuRNt8Z6gSU
jgkHwF03iRg4pz1jHxYdhHbK8owO4rPH+95LNDBnP3ZNPhQGndMd8zxxbw/RHb6dUf0XGENjgvFN
/NADv/DaHBwAcgLiefZT52aK1QfNWswUCbWZSGF7CbYNGBuWjwA0D/nrvLtQOuBnZcYa5jD7R6hv
0FvgztSKG1TJkUBQiZZcKqJuQkeqpUidjulF3oMyITk2Dg6V4VDzTW25xdEB2EXvBghawUw4CK3o
Ckq+YAYhRWxFgU5/HGY1Bc+OQlWNlKsT2A2T87evfF6xva8PTjsScIzSq1bulgjXYwrrJ98QY6rd
qpDhjbMZjS8nMeKFdXNfPr6P6OcqscKr+ZoRoWNWh1VWKQrz8EldX0m6yXsPjUOqvxclQCC8C5NP
ijEXLWSNkXDCSRVQs3a2Kr1hXPRFsZC8IkpdPDkyaGT9gTJIok0t7skKxH+vOt5f5IVpdwNxbTrr
foJaoiFMVCKXoW7uq0pmhAsbvKJ2ET2W3/jdNLjvsEjUOqXsjegdjCqWv67Uwz69SCCTVMk5GoyT
o20WvKKatdO5BPE81LJ32A/uGBn2KjVedy3tHeT78CnNRl7SHDaW7LcBV68mjz8gEMELSzVaWAnM
wWl97HvDF5m8Uo6MWD0VKMWDZ4M7YeY5DkQp3nvltC+Bqp9VBclj+APRIwE8rRVpDw/EacmZFX+t
T4yZ784/adc0hCgGj1wruMYdhg+TYDXI7U4g5bVd3BQjh25He2ePrS+2us8NEh+y45vEPGuGJzpx
jdhvDwbsm8aY9ZCzYCDQdAHFkXayBC3m4lgD1dtVMfILVP/Ut1i//x3Kw5pC7GgqVlgt7F9p83ux
ZYpfS2ZSD7bWSv0+wyuf5jdEAm4k+Mx43rcjeC0od5ZzzjPa/s8dPrjvtEy3CJ0LpU796pz1THIR
/S/+MjOrMeCMbR83C1PvvHAyOyF/69B2FdExg61PDThWOFmodju46jyIC5ozo6PeTAZUXidu6m5B
8hHF2aSo/5uKql10NMC0zFt/DMtieKBNql3Yd2jsf74eEJ1SPQs7DXcKbhfWQvW12TYTHr4lNR/+
hVyyjp+VGS7I7X+7UtNW1V61CPBCfVIv1HPRCRTKedFcXnn5SaPvo5WSnS0dflRlSWplPop0qZGC
EyTe2wYp2UAa6MHWRGxMT4Tk2T7BanTPHs3mJFVvMdMqQs0nKOmqD5cqQ/FDTBA3QUfsSEF42PYI
ovygtIB3ANBJjrtO0Vf4x2FZMKcsAM3q2GkV9z5Et4WJtxPl/O1AVhuBzZieXwtpMfH1djNl5GAg
8FXTONclb85MDthqpvsbV5Rcef1BHPyELbQhCisyjfBJQ30WX13xLTu7gGuK2AOyzF02Be5MiqDC
owhrq7TeL3abJHnSpTpYtjsLqpSx8mitaCf9wbf2lS90/LXSCc4ERHbbd74llSXaDYtPRls8AeBS
1FloSh0fuI0u/G53zv3ijxBgD+AZB+NqNAFQQGw5pXYcEHRfNTmeQQkgw30RIugFYI8bs7WBK1n5
9SPCfZlYpgDRtOAgWSAgZjxt9pDqqhZL42Swj41urPqEqlbAnOwL1D4+lgV9LQydwy9TNrqw7sRr
GZxcHO025O2VVot04dABLd8FE23RUmyPt4//cxF8rqDLI26Rfqy7fP+BlqGT+Vum8pXZ+h0H0aUv
cw1VE3Qr8eBg++ltxMHpXo7uRGgMmA0mPi7MGACSlcJWw/gZrioEojWErGRrQRMafRXbLimc7uXx
6on6pasuQLQph5ULEJxYAfExFeNnaABXy2jc7tkxPPgL8fgTXYkBHK1+Cz1ELQ2wV7bYXKAprGZk
8kCL3R6krg1ui8+orsuCVjo4ZtXBUcWEdVR3Dik4UEBEdabaxWTMzagq7YXjtUhW848OU1MXrsPa
RY6NO9qk5XZ3IKLZWWYrWLnQxCnpk9tdehC5AYjVfLoCRT+Y4jpkTvG3tP+Gpi3Ej6vNm79/JQXx
kEYk1AnmNFuJpJLG5/rLCOueFyepp3sN47IKHhjGVczOxQsraxdy0JIoccy24Aq5xESep6PdxImq
3J49KrTTVbkQdUmwnJfyN6TXbNeZ9OOfMbuqAN+ZThgjD3pvJgrOOFhl4m3y61F8bvubSiW7a6fR
9C9JbDpSV6y+vRcFDaFv2J9Qto2UZW7fFROyUr8GBLDAt7JmxxyfDfFBgL4ez76t9PtBIk+BkDYF
/f2WHzXJ5QoM6dIsNpHj5OWF60S7OEILZsseYmkpI+0BGUkes9thrmsuvPwdW5y5wOKPxXmyc3Hy
FQrABA7XPku2VbqoOdzfMt2NtqDu3U5dCA9vsK8/6VfttrkdYAOkMih+0a8ZAKkHt9pYLiZogBMC
jETSxOW5Eh0/uIJ6Wx5ZlOsAptpB8U+6ux0FRuTuX3ubjERLEnaboAlvW1MCtQYPrUGgzOU9aVEK
i7pBj+4Oelv8iKNfYfLcFnB/0yaKKtr3d7MMCSiRqpKDjRD0QUZuEwAJer5gQah8bziwALKVrMYo
H5AwgN4lWsHRLZaubOerjFlPonE4JdxtywEUPVAnRyVkLioQUBvGmgsZvl9qeD1zeaAPYUdKSJx0
57Qu30XF3sWWNv/wULyoI6NCNigozV9Pz3aXfe20wH2GqBbVf5xtIB3TgyMUyesJLcQ4QR78UpHc
rgKQXd5ALhZ/s6APOFxuHHiONLta8wj6/lQgDmYKPSjbtWqHBPYzM9z/8Cy4Nw/pPFKCN6UdNQEl
tb7eOHHu104ZUWVXmZrX+wO4n8Ox2AYysL6F/1mhy2a3h34sy0AjMs+ABGkLJIePV582TeOdW8fp
CarBNdEUMEkgaG5J70VewLAbJM/WEICTF6CbYC0Nt9a4nUhQogmU1w/0GmRlAs+FL1s8kTXSzUHb
ohBoEBf58uGMEBJZk8ZHapAEt5eGoYJx7dVOIADdUHfBK3hJ0U9vrBrs5o4dQ3IfiUuvVDy2rHyP
1JOf6STG/W6XFXM2m5wVsopjOEFI8ZH4wy/JantGgWZm6q5JJlslMTX/Fs8q0Ue1lZSFCxCgQEBs
nAW8UmfmY44f95VzlpA+auCJnsFAGSYhOk5sFnA3k+nwpFjNj4KznEn3yB0fuK+kgzjLQhkqZhsz
wiClrAxhrrv5+K2UNOWpaZu04vzzbmwWnLRKjl0f6q+inSoFR++FWKkppSAxvZaMoQD97gk6dFAg
z6IIF2Ok+OfKvbr2zi/pi21bf7tMMhUQgcXPuF2LjrR8E+venHFIyQ5hfTnpwd6UErSIAyW+W6QM
1ga3hkDRGc1KWF2LUG3tKPDlTpeOD52UtvTJF04zl0PjcQ07H8j4gwMEY0mgC1cQh22t9ioOV/Jb
ifrLB7iMh1ib4UcWxyGnfLVVmScxBTjF6ybaUJHqA7d7ybXz90FLaeHK8Be4GHw3iR8oJkeMg50C
QBjzJEKUsouKS3UszucFEgmUJbxpZUihyqlQj8VxlytSIbNFDa9kjn1cpc9TeebZOfSv3DFboaPd
dH6OH7IsrWPwMeHDCazmEzixC5A8CTlv/jYFHdft+lltkumWrrQISbNyRCSJMkI38oZccr8FU4IF
tYB8HxePKzXRTPS2EPFU9uggM43udl3pQblRqZhiCZCcF2klg/s77xGBg8iQ36E6Et7pWpQBcoL2
tFCkdEJZtY4CEvape0ImYjIvcHX/9NQulZjvwBFIZ3pp7eUcCAgpx90KHlHd4CnIWvPjQTUauKvi
7BDX9DXqYThJqjwHLHAW2fuUurWOXDT7kP5JfVtfFHYIwHiDc1hQsoQXHnXjmELQe/D6g7BsYM2G
YMFSn/N0VaPslaSgrCx4WfIIbK/NcC1fzfdMVyAEpR/v93cNypeeKSrmVfDPoZiL/wtSouENx/Q1
nNfo182lJUC3BiHTuQFc/SRRb1OeFiQHRgXDkCawqVQt/ZI/l6bvU2pBwVxWOAz/Cp5ki4W9bk/A
tLhdEFQKMgb4MpZixtLRqL8Um+cEGchP9oTJm6qmP8U7svk95Ld5NVW9Vi0LOFBmbUmlynva8pXh
/8waLAR83XosYwZBUFDyWYNU4F1Gl8XUnj5rwIhH4UcpFhTV5iLPuJLKi+pKdShPlGsd5pLkTQLw
y12GaCsEdbrv/C15rD775/h3OvunBP5x9LdAIiSqYzm6/gDoaxzYDUZXf2lkAwRob0WEOg4qta+q
GzW+/OlvjO/iHA4RanmxINVOrp2LkyTsOTU7JTh/h52iXnhfjXg6Bt4sV0tDdUh+Cci7EjgTp8Vj
0PBVzrzC53Bd5pR4AlwaOwSCvIC+WXtaFF2Fv9zd66MT7elGWLs6fnx51dwfuZcBl/kjndRr33LP
FUFlO+UNdrN3wuU9mGzhkv0W7nyZxGN5DE5Xuih3zgX9JNnJWjdx9iuawg0CPTgEL3h5zE9Ko1uD
4AY4AjO0aC7Q7qqtmqzrloqAZb65YSg0yFl964eRyaC/ATJW6fe88B99nRoFqzsPvvOgUy5ISDTv
0KQ76nLuxJ3T/cotIeO5Tbs7pf9f1hI/kedpkcFZkjnDTBjXd6QBQP18qzwvCTahiG85ZbhKIdo6
LsaTyVokf+q25vV4d09X8DuHi2FtSWx0zRpQj7kVWpK1UTUNkJ/LuiBrf0P7MZYYiwHWemjKO0Oy
mSKC/gw9FDTTe2cQuRRpB3uz7kXPlxuBfJZL7i2MdiT1FlreGn1wI/e8CA1OHoZL6yJVOHjtLSXz
0DIwCJ4qCd4q0TQq6lm2sIokR4VmUmaUmEz3VuwMWoi/uwHLQTecPfwVSGkO1Wxs/nz1hpkJKxqo
8XIoQ7whQdiOfx/XSLzYkYsqUXGFMupHCQeyuEWe/HwCFyJOdOi9qcy6WNY/hybl5rdECUz7Yl+M
TQtIDat1GLyCUsW+gbCOCV3ZAtXlU5ijug3eCRUdvyXNa+fDCl8v/EyecQ402j8jfw+ozpvQHuVD
Ew455ur+a5hk0boBIUv2RZ4ZzSdT1AVwQzWIu9LwsiAYCSU8eEPdUCDZAJq+XzbMzyg+UCMKyfeS
jtG9Rd1i90XuHYpQulcLZxBdyjHQy4WyK3+lFWHAF7LrdIYzj3Ug2GdwcrrzXfEW9VCd2sGW2h2J
dgs+GXzXljPvjyFViwybyLsbxbRwCTC4rmmcoIqcwhThQYlw07RkKFnUiqCQ7FTLWjKDV8kbGD/r
DixpUrvWKAv7JWELSoCmck4k99la2ey0OLF4Qg9amVLmRkVtOjWFWQXoyRUX6Es3DzFk/O5iUUSs
wvh+wtyQk94iQph2XaAQIgxU8WzPcKnQ4rgdZiZy1SKe+LN4BcgTnZV4EE42KtHGHH5IXaem35oq
nsifZRjp+ZOfcKZIuFAaaqM+ysScC4h7Iljs+T1tKqW7TscV6WbbLEtxGMucpOfsIpM1MyjLwpRA
S8AR7vBoObzrmdbo+Bh9Xb6N7dvyz3Klu6jz8X6ZafHYDDH7QlQxTK/6CK/RFFfPELykbiWJiHnk
rz0lpd6I81ZHgThM3JK02j0OxLDKMc3RH9fkQ28VaJ0cVng++hKzsrefrXz0r0cFZ2X3p0REhCGM
qgTTGTbKGnLQ/0s90GJQlBmQRVeUAF1fBqNsMrLcPzwG6RS3Up//psqj0neDHK2XKmAJY9PbZrCc
rn4ZLHVUCDqvEgP51cqyFVYCTlqIX+OTfJKLPoePTc40ggzDDjLpceTDTVrQ6XV8K+sTepAGmpvJ
xsoUZn04HNKKbgy1VfKmQrfw+1yRYQjiUy5ctUrTtT+pB14sMz4EKY1V6gT8/SoU+q0QXXbFmM8F
DyCamOoEsqp7t0PXpar0XeJHufnPHemKI6OLz9jzlhk8PY8TJSdXJebkJtlxzgbVFtu37gnKcMx2
RQp1kMsBXjSTv0mafKv6E61cbb5NLpFyfpE31/URNZIjD/LIMdiAr3aByQJHCtbrxvDmDkOCKZku
NOnNORRM6T72a0lDqBsTSePX713daBQJynSbsF1ljilg3EXvSsiHA5lzXKMbmUCY9JXyj6te1xL2
WMaUKB8TJcJoIcSFtbKolq3ebpzg7Vt0jcSrh0Dl5OzD0qGq7XqGtrbVmJ512kxF8ZS8HTG0q1pi
cCtJJBdlS3DKLMR5OyiDBFuFDUk+GRha43l43vAgQUpzDVSr5nzOaMZ1EdjmkhjEFHrC+K1QKv0T
XooKLkrBr4ZjO4T4vI9rBIv4Hao9E9COvEzuNvVrzTlAcSS1SQQU55WJyQRDiZJMy4we05Ona+0+
ON2LJH5kEttRNEEUBoMAjux8rBP7cxo5fQXUCoiGdiXVPHjNj4+rhiJXrbfTooEX8kh7nbodAPHN
s0vYPyjESjMTCMOaTSqRQW6ONOvSuMemUSuCjvYvWAVLj+5QiQVqFOpq31y+VmFteLYM4PYHAb82
RvhKOKdtLpV2zixq+RrPoQCarM3bnQqkMqLNHG64qXD5fn6+PDwTsbCsExPBn1+ZHj6lVZ2Y7NEg
V7IBXty6a2LTmxX1ig6GyYleO62pQ2dlcRp2MQaE3TFZX5+IJLBTw+QlDhyOFO3VSvt0kgRirOcz
ZxCBr8k00bNdnmWP0jGtt5+Gf5+xcegoIlFo6Hte+5THP+PTSykkXHYGFuTHAh8KN/oSjyJpivkH
Xrss64oQmDNvbcev7lNz/uT17wPo58LdINTR6QxxBWwhfAsITyJeZ9eD+0XoUK0Yg2Zkc9h81gGQ
5ysDCNXVWATeIzZOQ4J+wd0T6KV40CUzjYQZP+30dC0B3NdjKvIsAy2UGY6VQYM8QPI8fPXgIf7e
+uH4CCq7Ulz27pAj441h2oCGG0O0RQVN4s15CfyxRABEmffBkqZFs0GAIg1N2QTx4KkLihAhM4sT
2wFq7J5BUal4sPz1ldOagAydLPMT8dttpnZu79j+qTDWDOtj7KaH619//BLl2hzypjPWGFoyM0KO
/dyE2gCAXI5XVjub+jBMiEzWpCfGsePMSnzAbpacRZbLRe6S0+eAv+Wu29STSq4IaGmaUuPPaZvg
iWw1V9dhcEHgoKRq8FMQKfn37yMuxuqb4UZYntXB4ObBAgN1qCOfzpdnV+kwaxkbmduE+W50ThTo
ultnkdo1jqB8TejMS6/YRQ/UbreGLO5ZpvywJDgMk6lUNio+hRKg9NAdpfjlFtoORG3cpn7jEA0L
cH3NwfLj464WBPG52VYTEyPjhDUV5nqu+GGiEbfk/L/row5bkQ3b6TtbjIMHNdM4JNzNQIaoezSs
oPIJM/DGtaM6iM/tt3mtfFYC/IMFiYdaXl1waL+8jS0b+AaGMiU9K0UmXMb/dg5eeBD0RPw/DJZU
x3fp5RRjxjzRzVHZy9968P4C7njaL7ZINE0jNGv7K3VzomgG5VWW6YE8lbNlkYrP88140jtD0JsR
zI9T83xCoTfDInJXnELh0rC/Xmm6KnVtiPsnWW/PZ0W4PePyFUQ57RVNn3G++XBPVDZlOIQUwVY7
B2lmTsxyROWHkBQdVkZnDte8XOfDNoAZjjXzuqMcHQKZkkHUOIbiIjEeEnhmoPSnP8OrWqjhWHeZ
YUZCJ4vZmQRPz2R2tnz/GMZVjX/V3ygsr3ZsE885Vyzg4I5tbC4hEPJ0bWIZolUWUZ0vWIalGv2e
oznFOh+Nr87UHoMrhaqyvDr4QRt8udvyS6EUXN0IYxJC72l+BPm6pdaR58v6mMMkPiTay8pozMRC
3io8M9925VPbcPhhC3TLdqFzjguS5urBNtJc17MnQJjDEw/gr375fsSxHIaa/3FT+GU9EwuCL17R
uQB+bhV37GTQSabaD5JKIJz6Wh5qSqhbTgR0JAF+pgjJza0kcz6+VQ+ySmUIQKvV6rXCdYaD5nRR
39ks14LIJdu2MtuJV+j/6iB97dFcfxQeiJ5d63VtMUhaeiPgbGKsD2/V6K9cmBPottVwZsnQrwyy
CeniA6kiDDycABLwpsDJIJz6rIYJZ8M95u5FnlM2nPgSVbiCpX28qCOc5PJiDWG5xal0Y3iopy4F
yQa5NXvosnURO6mg9Kq6drboBsrTWKZ9+M/kHO4e11E/w6vZMBLoziqZDWVdSdpgXd92NLvXiiUx
ilqmdc8i30qDgeQ6c95o1mZcFU5L70us7AIsBXtLmtxr/Pt6bwxvytMHdLZUyUzmL1+r1ItkdoJ6
bp1yLJh5NsQhvuV5QAMPl90uiol3Rn/H53PBCVPpYIw2iNUPSHQwS3YbX/6ZXgGidvKRRKfXsxvU
3OCr9k3HlS8jyRl8hNhatb5e3MMHONjufJ1prwWGLUykHD9W8cxb1kjEEIdX60LvnJPgjuxB6dtV
mMSHI//c9RcpiS1t4jcf07Cvl3Y+S3S+M8zX3USirIHFEmQj43gc46OqqaUtIdhbgm4K0YgAqrgz
y9Yxd6UfzCt597Lcm5F6IT/1bWE+JXV8t8kULa3pVHA28v1fkEbIhIoOQcrDbYZ0nFSHLso9LSfW
KfHL+b/78av3Xo/12dbsAclv07qreuRs7zAEjylJ+V8kIXsG/BjTuearmpkjvecBIiqHS5e2tKQj
fx97+99v3uyIJP6szVwDTCrDWoaLUWMvBX3PmDhNQOnCPjui1sSwz7FTJVzPBYgy7wucH1C7Zdhc
c6uEei1F/FfTz29eHg/WRx6KgrFAuZb8+7LU2rr4uzide0/3SaVHh9RluiscLQi5DVrf63JaHjoe
eYiU3rxeS5sckfkiyoyczD4a+UAk74LM404okZz3DEIOJaTa9HFHBC8qH+Uiw+0gOKHjs8jdKDzo
lK+8RPZQ7w+gMonhOHyLdjUsaH/9e9nDjXJIMMW1tpioKpfo1SDGdOq3zRvCv+ye18cuf5SQgOac
xqrXI2wX0c8CHC1Lpwwc13LQ/COxslXCJUvuZGMJCRkIhIVFnO+FWZ5Ga2hDIH+OhP5UYs3TPx9v
cjmLHVd8mJbEQZPpjpbpjhkfUDMoH77xhAq+jS/mV9ZJHYukTiYLiHzyW8e1Iil+X3t53NAD2shI
BobPEb05K+jSE1HgzdTVT7K3lLa6eCxmIl0HAjVn6Mdf9C/s8H4s6/IDBXJQCXtfIXsRi6U6n5Gb
Kp9UHhpgOPyerAZJqEFAMGM85S1zrdbwRJ6LHaY2ILrsU4KWR4Fgo4Hlj572uzlTwzSTkpEkIG20
vxQOvyGOdYXX8HOw5pOKrvL/O/CoAFyQKLbxYUoR8i+EWUDlsQ6zJUVVwSE09DV4JSMN95MwAPvF
15VEbqs7XNh9ec/m0tHTV+AMw5g8pX+tOpAwSPirK4GrV+7B1kIFpJ4dDnYzWW0zrbvxmj3pHe3G
Mb0HuAlK6JFdirL6ZZpDelIuCz3lqNzU5Hz0GQmOR7R8QsGERAokjioe7p9SRElDLnDgRE2/7kfW
nL2oJLD0TkxcRThW4BCGtky8SjCoMp1VF/MTxqshrhmQvG236r35xEMXxsItwKcqd+wSFUmw/apH
apareH1A0zJtnvUS50Q3y5IbSUJuiOVLeYPxz7EZX1/FzUmUdXqNak9SSJW5fXBii3duPjclE/fw
vIHdENRk2xpK8HegJuJ/z4lVAIssT+La6D9/OEzA0T0cD1tkGFNSnSj6ypyb84spQGSRYBdVi6Yh
BHiV0dBVdLmmHedtaYMZn7tHO41A8YfTV3elC8G5IW9ZWv9jQrEmOtTsCmKx8tZh9/FDRIPp0Nn5
HTZGTHgQRLBduBCUCWJVy8EK+cSlzsjcnLeWui4zHJuQ53kPdvm1cDwNk8qguPnO9IARnPbfw6e9
4ttLzBSjFBsnJ4jKT5xfmLlO/TxYNM5qR23z4PEE/aqQOHfGjd73ErS5NvA5jZtc2pEs8NW6xw39
pB6t2TSJGo5A8ozGT1yAjDKeIutpPanHkKE0IDwnYiXiJ/0zqyznyV6DNiTy8qKleAhpfA/2999d
DQiCIfzixv1V6w4d0S3rmTSRDuMXl2A/bT0giWwh2XsR7QpVNFebisIakoDYxVej6JmyGaodbmO0
FGjR9BJMVKmAdbbxfrlUptbsrzQmjMZOraH77qFvT91ASv5glC5KIVo092J9TSulGKByUsuyJpns
PGHjENQzZTK9rqgAxwhFquD9Vypj+b9E/5CrrwIRuJUOPOYfawDJuwNARQRlFa5C3GFga4bIdxSE
9d/+HubtcNcDfBnhSnjUX7uBtlTyFOmzbR+uPsYYx8Er0LQFcbqHYkylqQXlWUA1TnI8UDg1D2bM
+6Lo5g2bT/VjzvvQDVJXa1kvQ6/5YvNbOVgOXP3ppxLuSUdN3ZZu2hwN8i0c6SfVuiMsu75IZTFB
hl1XlltE+LNIKLLLba5iF1GPDxZP8AJpXVZmsLZR0RkKv1vUIALttl0GUsj17q1e6mIIJEranxpz
sKVTKIDlyMKrrEnZ2luQCtkiVjQ5Piii/gxkVOjzf8WsaVm9aD9hGnbuXQQITm+k9+zXixu3frDR
B8+o7KYznZJEqQpt8s7JabezwipcoHPYvQ/+vja0naBeK/Tf2+Ps9r6dBTyz3hwxybeK29Zk0D0q
nXVbE0pMN5kctg7eC+XLvbMQ9ochVD4fBufQnz3TUBmZRpKOoW9tzbGNPquwTbihV2gZyonQUHxl
J/fQOmiLCvCURQNAmqm6XfRAWsDCAFBU1dKIYJEbUwp1OjR8XlBE+dARIsjCDaK56FN/yaLZXVQq
5BcWkylr1oym3asg9TQBZ6KQn17RVdgvV8IpK/CxgGRzD8kB7322Uc7ehS0c3Njdwgx+bTQk3Llq
zkPloJJMXEv2GTE86+uLOgOYHzJvW4KwZ0B9t2tE+28T9DCcgxft2Q4h6Dr7i6bDFIYg0OvaLi5c
r05zpQhHahTYX2U3QlcDcBWN5mUiebZNgnipsrI9pTw5Pvp/fcTIx1YkbxhOKPbMudKhRASEgDGH
Ba7Q2iikm3Z/BE+o+WBHKHJRLh7UZ6s3HmYqDNzlwDWgAB+Jvu4B6XPECchyDdzu8GsZf4I7Uf8z
qtHQukhny1a0EOjVTswgCvCCMEdjYKf0vsi1JTPci1e5wFfjbgJVkfmRH+zQj8t2qEqcIHYGWaU0
4uJONpzNDJO0LCXAbO6/RDpPGWC4ye6cl77/TX7vcCBUlJ63ViqDx2u049bj56/ZYeW/xCaeJ4GN
y4hCSoSm+1zhx0TuckaZLnFmsNE0hmGhILb7QIysNu7Jx1e/ZNfX313F5wZJ3afVlE7q/2duULWR
3xi56yqpEilbhGJNr/J+3l0TWuBaiWPVD7U1LxBkEX3B7t48wIICGZJJlPDPl+jJkBl6UeKBx02q
0INsCT0dI3I1Kw6fyDv+t2vj3WJ4Bi3JcsVkDfIQTlsiPs5FYv4OPerlniix4r5d6bouQUlfs8xH
pmae3tlD/vVXv1X/mD1nQx45kpevhdhxGUsxxAvzrOrpxStSjbVY7aUP1VY2yDu1vs4nZYfjtXdT
dYYDG8bQQkDQGMyYjNMFH0cnq6ELt+R2M3/im8WX0OlI0lFPXPfsjuDZfukY8tQ+iOFEUgCkk+fY
8reQ28/FyS90vr8l6VqtlVxz4Au41bQ7qlqpY2wNP6lamRpWAfhzv9nv8q1wLxfRkXgz4MntWIfB
/E+oFqfbeaTyXLbs0MZfJbSo5L3XFitWCxtvgVaMcgMVenX58i1Fg/Z+rk9pu4BG6fVkZvCpZ72N
fwYjBpLTLSF9POweW1AGXy+XZnGUBCkwVm3XB9T+fFF42ipnwohgeK9QH0mVDB06oEGdanU+021Y
sZg7/i1W604CssmBicfDWxN0/AhP9D3pu3ZEgDU8TCF27qlo+HQdSli7qP3uipS5jksbdGTT9PS9
48b0GHUmAgbTqNmKDf0OtCV93Ftm08n2FQrvTa3bJKLe99p6ldmrQHoTWsc9wHV9yS0xgSYb2eQS
Ij0oW9lfteb3XGWesN83K5vsdqU79TurGjr5JXFTRudOQF6Q+Hjg/W2NwPXOd6OpdBlrHYrXGZuO
3NNeWjKVKWNPf7u8Eg5nbN//IYyV/P+U7Oih9aXA+uU0qzxGyI/aZH5SDaia+Yscb5ViEjFumywd
p/l//RDfHjIKVdcbl5jUpA4FzJQSwjxK+HFwXeIUma1oOKGcPJ9L+SRNw+NFtjRue6RouGRACUrD
4/Tg2y2mAziOG9YpbBmdpR1tSw5MfKB3XfR3NPzRXQAVmENnAUEf7zSphNkh4GNCBJR/O9e88E8z
/8r4HnDfbqvFmj1NZN7BmfczqgAWyxRhrHwsBclMfudARDlppO9z4qteEvhFPIC1pDtLRzhb7ZEt
8f1eGXMcDjGpe5LliDb1uM/ia0Kb54UM0QPRLdfDV/F5wPIikF0YX2vVVGBglGW99nm8mQEYqqqy
x/dxz65EJczN9oVevlZsaqvjA4DbKZMb8Nngb1QFsHQZxsSlGAVp6keBgX7X3zkE4RjpnIHD0F0X
tYqGIgVkERkJp7aa3i0gWGezNl+Z4mfwS1Cp0NtbnbTDtUZ4hPhqwXhuyaTqZS4joLOdzZ11ngAC
37CysByfYjLZ3w7aNKJRSCFUrFt+N5Sdjt7ovyWAr+zzGst42JPyxcIyJQtfETNyVBeNrB++yx4R
3xpjsLSBcoWHKbdZEoTLkOHGL9LyDjH8LFkizFBypdN3ecln0VrhX1igZKhyyljTg/HRueSK6SDl
V0b6OQY34SvgICo4cq8kGt3PfrQj7FA6KYQk/TxFl+xgNCmd5h2/eOVvJXdgGfjEj40Ul0Qrof4G
qJF2QwjzvMHIKqDDm8Jv7Ad7eSPDOhwx18e/PR3Ji+w6Va79AANyZ1aY1KRGvZbuvoTvbgziNId5
MXOSzVfevNWP4+EMFJ7ByApWruyIzJqn47ii7PWtzF+D9fCn7w5DWkHIE9PZ4DP5c+VLu1qSfUDT
zqd/uWj+fl99XllyNGdgU0GbF3mG1oV9uttJ0pLU4elGVRnzTG+GdPIZJzvKjvhgu9m+V8Sq9USK
QqaZCIDdSHLVtqeSRkVKuuPRgJ1yDhjW9MrWb8Yz8FlZxja8J4kr+vP8ive0tDaIumN8sV+ur6ip
XaIYI4O4ul1WrQf3B3HWlbw3ijVuI72Zo8NI4umD+wvo8WOC8sZzegJH+ZMI9RCPRKwdgTUt72YB
Bbg1csS5ld48MYk9Pmxz1/2RyKHBgkHgzLK4tOhzE6dFNQHvBZQ+fmhxQ15QZ42XnI0GPDIlR84U
aE+4MPXA/LtQYWyUEYP0eH4CPjfX3wqDzkfiGZpDRfArdkXj1tPpd2k15TJOfOm/fk75t0gOu7Eo
CxXovBoJeQKL2K7C2Bcy6UV3lGzNGVT1qMgd+G54tNsW0dOqV2kKrskdYI9rYfEMJZsU3vOjRMQt
tLUokwrLRizCOtJQljbNAwDOzYDOkuv8aoPkcKe7khYGr+v42rvNaGMJwnw2xIDEpZL6MI/JmQvq
ZUurtKS0e9zDcspribQE+lF0bSxiP5wiTqWF9WT1iR5PCR3np3SfNa53jQ3No4BhhKWw1yVBRvX2
j/MC7xPSAy0brRbJHHHTVoDyDdVwIQvrq239RFvP7FMtPd9Dv82IHzjYUNo6MuUmyLiDwFVxhBPu
7EtfdCufLx/GVq2hWiYxB/2bpUOndyyEdWNEuW3ZJ+N7EMYfwcEjnG54I/ZNli5lYzlO2YLWE7K1
O8CbwKTDOFxlymEW+gxuqbVKann7X7C78Vnth3Th1VPDrtd0x6rZey5QNMa42i3C0JKCGgBPjLAd
QgRgJcor8+n6p3n5td094C8HfjLP/eWKXHxmMJiaSnfSSQgJ0Xa7jP7nUZQH1ASgr22l8M1Qi3eC
+alOYnzd9rtwvTWGzjew1y6jOjTUEwlPUcCSQTb1yTqbCfG4s73Ia9sS4JKkUSsgMiVhFP4+G3ej
y0/DYv5vIS+qiUPO+ITFOmT7y3TaOyH1+oQSmgFCPdSTuCwLLCWLQ/tPK0HA952vvm5ITEIvZQfY
IUNr3N02uxx8cfNRCNrd1D+UGnNa37oJ8dfIkkU2xMR8SSx8X3m1GC9i0fHccGP99JX9SumnfMur
Wf9YO/XorU60Z0F4lT/Wthi1mIgD6x8mqrgELLAMzE83nWXaAYwlrEAcNMEba5V+OfSRfZf8fjDf
idvj7QNwigyYkifQ6BBVhDG24gKOqHYI69C0tvoEqKL+AawD+CiF/w0DEjfeQDKOhTcW1aUGnfmM
+PL9N8g6EEoCo1R063IwnU96ETa4xjFhJb9vCyNaxFejPT4GEbaUx61roM4Wb7Ue2pCAHzHdq59C
3/hAPvlC0kcLEXZiriiMDbU3ZR+or2v2uo0kjx7vU4MykO5QpCTi13sLD9+ZFiMg+sZ/6ljEfzvH
FY9FW9ZGV9rQCd05NOT9rHbjL6+EDWVPPEaNl/0RVY1oRbaP/akb/bgIYz9NbUWUJII/Px2FPPXT
Hu5+aETgJrOVDQQrzpw1PJ2Qr2dcXkNacm7iBgY6N2yNoGA+JWugxlD2UmKguX00Ue3+cLPCj8Nl
0BVbYH+RageNEWtUzpzBoNA0IWHIFMski5i3b1fBxJha8hR3QGHeTKRkTaMTJwg/C6OWxd+dHPTU
CZg5Un7QG4LsudENPhgPZSqFDv/Ol/z/PAqBWWcLyeIp6aEDZq+Ulac68RCloUG1rTv6Z2A727Vf
o4MqSwg46TyqWuOzHPwITddhXLw2Jiqb9GwR0oOEhD2STIHKulZf2m7bc13kcaahlsgXW2VhbJvQ
Bdeu7MqrPOgH3ywjKJ575X0HgELIH0fkg7IZc2jNTUW9mOXgGNqykVnTHWAyAZJ9P3/B80Z4OQhn
eTayQjuiYhfpeoaHAlSpbpTzCu3a90+lyKEVgzhsJa6q0nn33acmcDsk9/8hsOZ1wXNrZckPc+/r
qe6YPFuH2mUvtsc6xV79eWq0UkLgNsC5dO1JHLbrRIxhq3mr5/FfM5uh3y1Oo2/XvY1Z1ZY9BJlT
glPNKBGeNQ+wouKosWL2AFj8kp+NimJmx53wptqKoN2RA7JCBLxoexEWs7n0JxFZszGVkMLR0rIw
Ms4cudx5ALGjINg+PQHvhzwFwvrubzTmYnyYxvUWEmUJkFMcecq/AhpUUD9l4NogLSl0Ewtt0cYA
pfWgitk9VB7I2i8/lRHeE1A5RxR5ERpezK9UIWXoGnwrHHAmfIrVxFdSuIAwH5K2EB7hgIN8zZPp
zb1CYuinrr9CtFVxAFGwzKeJImf6YEogdhIic1U/PMFvYyRuypBoCkAFl7SiKKrlvofcmjXfBY/T
fNovLag1zd5B1411j8A+ZhFA94Ny79ANEyOebs+I/H+0XCTA4CltproIpRjIgTTQzsB3DI+uNsNK
cEJc4gHIr2BlSnvAj3AQh0FcTxo2fUetkeMPwBP/t9iCaBvF8oSZvPI2B55KwbNvDo+BAPP36EcU
tQ9TnYCGG84JS6+rnRu4OHRsMHqLgZrrKWeCG8FWcbh70emYm8+BarvWH4qBcv6n0tra7Oet1WR8
yNFqruKLZ6aqG3glec0XkqcsmeWmRBtsrFsQfHytD+0KjyNaCZbSptApjYSvu/JAYDumvY9hpk4t
5Ltea1vshEhm8HYJ9D2muLCqBulsL5cPuMcF/EmT8R8Oojpe8/skvTuhTzwREU6jbjsBasIaV009
vdAGr+bjuprFc/yhak5D2SGBX/jE5tKFE8ftDIWmD888ni4whh/nICNrmdTYIMKCPBIgW9wMXR4P
m1sV7za14AcOz/Ws4mrbN0nzlNJtFQyN1s4MFWs7JKg1XixWMBKWOcohK1QOM5veSXni7P27hXGR
mJFPQN9AqkvVMJCLeU+RwjO3bxEuybE8ntWigYI7fTHbZN/L/HFA7Msw9o8fJMNkuZGg1BqjkCMQ
HV64FrWtki41gou53rzFdw0C3ojUyXVoeduZWuFP7ooNSHu84ATi9QEgwQcx9qsR7sexDXkfia1t
Hb7o9nDqyhHYx7oyCLR41deIFkjsR9Qvrv1g3jg8h2OzNm4Gr3Uh4b4y2lbHF+gEUsdxOnjULcag
BuYzzSy6dNkjeBxwyNkfU/YChBB8JUMJZ0PtZExxiZVjhbu+S7V4l8GaC1vV91SsWCHF7c7EGnJS
zOHsecURv2XVWuCRxuKXbTRgO9pwz5wXN4H0ZldBUrjVIZXtDTb6eqfGeLfuF/2KTs9Bk2U7lY9b
lb5JBXNTEgYID3pMKJ0ECOZCU7Sd86C/7/f7PRcQgxm6zCidDnkQkcBHLLgNkoUqwYs2cDSmke8x
E/BJA68BoNOLrLt0H/zXSzqR3HOjPGDfQ5d54FYdQ9U4tVZiaiuE75MsXftZPPhmynE2FvU0pN0c
+ppLAmuhOqfahJS88bF+SmmfsMovpXXH++XxrhHC/lpxW7D/qKOZa6A+aPjw5rSDDHeX/fGtXTcN
GfloJ53Y/tA1C9HM0vYUL2Cs8nZ87iM83WFXX12zPIOzxqunrsojCs+YNpdRbFWfBgb2Fr9wN8hV
/PLaCSt9IgzgWLp/UFfR4qweZigYgGYYL5/j5oniXjSkojj6fYxNglC/iR7Exk6xD/OAlcEarh05
Z9qTL9t9lrot5ppA59J7wP8pkqwDL3rhXbeYDrt+ADAdHrmziJbUn0R59sMEmBVbjfRAkAtfCy79
vxr1q65BD5P+0CYpNnDfXWyfp69SnMao6v30+ilH/V1C4ogHx3E339vysZa4veTR3TcRhUtMJa0j
NTFnIGfJoaMj/xeqOg+1PdiatSiqA3zl6137eOzv35G240icH07NgHtCM2PRfo2lITVmwsWuE0qv
2krmfKItkabwxpGugwNEQzxzdtQ9q9kVLZ9f2Xr47yTQPtQ+bSbAmX1aR94c/t/gq/DLskrtezvj
h1/unqdJ3oIlXHorWcMX6zTnkLT/NP1WFm/RSAD3PXc70yAJi5J7VV8eSE2X1+fIFYOXOCtFaKG5
4CRoLR6C4knXCUD+VAz+cDIwLb53hxwncP3nolmT9l2NTEMzWlCyHi0FbUxMVYiTa2oZfQvubYwy
NyFpbwNlb9r7othkJTgBm6t7X79ViWkYriVr4xkoApMJ+/fnkrgBvJhgZYPiQ51H16qNDkGypMDr
diOXGBgyZYVk+vSto+MzJVoa2jtLfjIs6WYeoQ8KlylHqTKuAY4P7fzd5AmOMFjmrjAui4b3opL8
R1a0PxTQhOZo0r0UcLgFvo6db40o7Wi3E47tZwQWW5g9+wCDqvL3eTJ6niar94eKkqeC06c7Ekiz
Bo8Ioc+DNq1WYUX0QqmI0wC2HYmH4iqbtLPVAxVm0LndtcBDdPgUemj4m7PQwuDeSciUnI2q0+1q
bY4rrBrcrYL7LHOt89o50qMI8wtemct409oi7ze2+sjNV/xCIzhHmPB1fXasRiVP6rSb4IMxXskd
rVyfu9EGzihASf62pZkbQUWPKsccCYRCPqcggfD1Tzr/YqClr2OA2v2a/FvlxGp4y3/My5d2q7wW
DJgyaxbIWEVPG92xdhCZzdHtddthFK1lkwkLL1P7Pzm6Jc4yAezSbAsra61UmnqsRF66CEal0RHA
5UzKqAxWCF/JibNN0QHLPPcjJGmjBnRMakx9r9AKqs8KQpMqKonRjXsyFfujKuz8R+rmi9n4Vj0G
j+xC1+uqxIza7nLT2v+moUS9ERyzWbInuDgbFF2dKBXy3etJhhI34leSQ4BF01yXQURQCMrbgW+u
z1YKOyn9MiHh5oPW9hhJJJfBHSDma/lFr27CnFFlDt7d3WSvsBU7nG6Ue5hhmjKdTDP/4lOIrbtF
U1T4X7p+n4lbfihDWvLlLfPM4YN0K43mDPWtJQNX0p1bTpqiDol4HiVU6XA9TgI9dmO+pJwu3tXw
c6zCtgJHF+Paw7OnFN5ztMMNMPElMmZUQU8aM4L3eQzq6zqaGnv2FVvNzAQMBVw08SR7v/DpQ4hA
xjOAIyKQkha6V7xI35BJ0hynCThCJiFQQStv+N57cJzZxbmPMLvl20+iOCklKCHqgCSxJKseQVIA
iXnyr6+hx4fdPRTw/2GqqH8mgJ/gskKRFDgluIH3ri1dt4vVVCxdsz8ks/jYgcZa+Le6TR/jZdlf
NZfwx/g9UXYt+tLhMID9lY0/jiP2bWbLQCL6EsEUrpxFWblgli/zDQWG9EMroLSZ5s6Ykw8b2opl
oEPP9gb3oAU652y5W76URQIW+SRIH4kOIXgBqTPoH4Ts1mPuk3gKREj+BcwF6PmnT3qYEhwm6O0A
2exxh/8Bb2gRrF0uVTQeM4QZeb9qxF3AMMQMHO2X4ast5CdMc8FBHO2RqPzTgYHG8D5SUTtqAOTN
mpDcGA54mlfOmfmudbgWetxblGjP7/xzmF771GIy53HFYH2RPn24fGV4K5J3FU4LqumfzyWr2miX
KIkuVniMytV+kA6rtUpEchYY415TwSPSBu+5mNAJFzf5kcM1bqF0+F2WlD4TlgporRdeRUoI2bII
Ak2M60RhU/7kcKuO07mCrOvXTrJ4cs7OkQLpGhxUKyniBJV/oLJLPbaXNN1cH2YWn4JpmuZjXKd4
o+7CHcXg1ylcJhNzkPEZmyrhvJLvjhHHusntrcZowx9EvVDxSYC3k7d0Ri+sPJ2LgwR3qHMUtHyt
gJbbCXVTpx9pReXYEQxLLMUDg+NT81emthWaJIkO8f1+6OeKGeA5U7wCSi56dKLLCref5iLU9QAP
iSvb0jqeZ66WNKcEmLE3OlJJoqTSUuAzypqkyERjOGxCa+F0ttIDiDvzyK16l/RIKH8yqU9L1HXg
AxmNzNRrX8wzdpkfnsn14ZcvUIhuhREWk9nEuP28/mEGutUu9/aWj5QXEB5sq4NxtthM/qKSncm2
yTnjrllXsmb7s+Qry8p57tPKYzn8lTKI0adueUKa5lZ9Gjq/e3K39Pnv37qBnTHlGHE+/MOryIfE
cFEbiq/T+z1xCtxWqqrpBPdAbQr/fAu5NpjKG77hawkFWUWW7mcJBVhwrzOl81efnutpfRkC24MD
7i3LH3SZwk7fIY921y80ULyB7S8bmXI+X2Tm7kNjYnbCcY0ZJfJBRV4hnVGHQiFG3W6NdBm0xg3J
M3Nrpg/c2m8WCu66jTLYamHpR6HhTRCituVyvcyAcR0jpW6xD/b1t+VxgZiFOg3yTWBvJgNVzbC5
4C4vWl/84+3Khsgs1HkrBFKccb/E+hLZZbiwJG9FZInvlpIVHL5+Ku+6bE7aJsoPjsFxtwSFPz+g
lxNjhnebfPnAbRJK2wHHYNsfT5DZFKuXRBki+wj2AD9ixRnDyXC+f2+V40tjbNHxA7smSvBS3YdY
zqYLJBq7q0wn627QrBruNHLFpVfWC/Vl8HM+8FkwCvT3nCQjyUy7cZCwwcqELmVwuUmQCaIiTB9/
8nFfqQ1GUHeqsUXSs8VEWYHTy1KPouzPwjWThRn3oef89OUCzhCpuOZC4G1D6oobXAsqAs27szfS
jeOfiQap2h40GGDm9DKdaoCb6pNuVnMd2+svLNgfycwBqcAEqOzdg4yz//wOqvRn5Mcp5b4kBmRI
pb9tN4XuU8yNQ0b0Qg+hEjDI3OQINiewzk1V9kP9fgIJCDlA9rvdArWrMxJpjdOjr5GF5va//Z1A
U8bngmz1xFaGyydqzWr2b62X4TgkM9uXFfPNYbEuh7mvcoJjlVZ8kTyoYXiCT3yzJaW8y4mEZ5FF
FdDE5Ts2nPf+R7N9bGyBwmAxgPZKNBkJbfLkp5tjyOP5yKs1lbEjT4Hp1+1YFandIR+Dl4xUArTg
9tSpIxeCxKyh4izO/sK4cFjU9vM/7PPjSNiKCCjkuNt/SWV+2Emc3pgyza8uYpD37XJYsrVLBuaP
DjHn/OUKR6u2/OqAP61acfg7VcraXrTy6d0Ejf4PGVnurUcOJrwiHYiR755jXjU/WN4KjmdYo7mn
ZAFnm1lvxCMWiul68pmIH9aaozlLZMu70iNyLdVJuMre+/yvZFPQ/3ytTHVmo3/x2sszbdy1M3WF
aTWone2sELWSVxenzJa3n/wZdlzA+o/ZIqxkeGnqpyRSJlYXqwvaycrQEqXfS9ItoEigagckXtSi
JbjW+Pj4lY92dgulzuR3HhVK+BskfJpjE4qofRA4k1LnZJE2I7J1JcvvVtLuIX5iudS1OFovZ/vl
2GqoNjgwtygg+L0sOFVuNtXDL7ae6zN5ZyZaL85p2Hm3YH2tGKBmeelmvvpj0OjJ+3jXvL0/kab1
0A7oO1UOADULM2BnfVXe6IYrVNhww1lU371z6BEi11rXYhyTR4+hslXa1Kx7gb+nS0e+y7SAQqBr
UVWFbTilx6fFjXtLXlbTslLVng8GzBeQkTu1CmBvK/t4qtDPMmWoJC/+f7LFjVgmiSB3F4NsCPpu
rPec4n7giRq9L1MLul65ROp8Ba1eMWKMpnGb1G3abHbVWhIwMGu22SfrfxaPVaycN+8SHqwSWc5m
8SrwQvthg1JIUgAjifY2EoGgmQGpKbhiEKUrJ0K4zLrMo1zDFnBwJnpRDPAJheXzNOHoQL/A1Jjt
P0Beg7BdLZATACWtFgDGyGC9Fi+feVrXfWwt8NbuyoRb+Lqxx8rfE+wCu/fnci5TxrWt1scE8i0h
esZXoTRxikDGgWZFzEm78NOEhO2dTbIvhy/XkBhyIHuYeYlHjlca8CNLdPHO2oeEMQ1OHmz4g/nB
WpiqFETjzixYUkCyqitMSrdLoAjnFkZJbkkZzIRb9pncmTkS2+ts47bm/eHi9e0YS1l+RbJZqmqg
/fPtig62hZOqh+kUCgkaK8xBLnt2F4LRD9kNmq44hABzqY+lcX/QgAgh0G+Il98QYHcBttMHyYCQ
vmz73xC9V/EeLBWlAxYRNnNIpdUpELL1hvkUOqJDm22oflStQOVb257F4KCyUMSuDvs2dIO0A8FH
ZZz4SG4mYuJdl6wTbgeWTySpGq2H+BqcN0eKkaPN1dlKO5IUq10PhY1WsPh/ZBYc7fcPqSfItmtO
FHDBm4M9EKMogZTlP/2TPgL4hejt98wq8myZZ1eBVY+F0oH+ZwJczHD4F2wMNUd+CosgCHM4AV4q
ZgMSrF+iXj3Xplc0Msn4sg8eAOG18WEs6i65dt2Mct/VKSrQ9q5Ux9gfl6sgviZEsYClRT0pOkXU
BNcMSmcYenZKbRFPSVpXYuwjuWneitjfybaTfSBLY29ueLJdB1CYDGl2rkA1AHeoCE7zlF9Zyozu
XwefynkIGPB8VaW4aQfhvl75DtJp1NKDsAOP9srgtd880b9TP4YwxZgpZlO1Adsm80xi0SJz/mfB
BKyIdoSJVIVU5jkcq2gtHllwBUryfK1zGxxlW4hJUdP4v+Nx6fwNcBTBRwEWYwdBFq17GobRFIqz
wEMNxGuWrXYU7V8dZzPsiofH/XFvB7lwQTeAbq/i7GGzYGx4K0Bhlcy6MwkqSP+snHwOxXraDtFV
KPP6r4yCih3nbhz70EksUfQqtBeAK02hRw/oZjKEeuvh5NWREN2gUjEWq42YqJkvkOCR98IQvl6n
cd7MxCN3UUXTJedUPznAjpsmJGg8iBJckOI+vEE3mAr2+9XggczwKU3RwpIYZi+eQe+tSrBx1wfI
Xq5MxPLbG4GpH+y6i7TDXhoK91j/Fqjt2jRs4TU04TN1eOCbXS1gjnfKCVIdtW+uhJllPRA3fXN2
VeGb5xAXNN3UCOSXjC7TN5jyHypSbnCwpQOyY7sgmfWh9iEc9twQZkSzK/W/eBOQwHbEpknNmfig
426uY+fBFz1CU4uE/bo+YSsZZ79izmPxQooo0RjbI1WCUVTBhEZKmTpFQhZ/TH+uDrcCXwrH8WOi
ILueUXFGvd3WSMd2Jh6upEuJcLgP/kZQrc3EESVXGmYz0rNngD/1qVNonoQbLgz35PXB0RetcqT1
P8C29SIACpCgejrs192d1IDVbH8f3h0c6ijEfyrP9wKC2St3jD7hY7GYVrO7RxSGDFkjzKrNC5XO
zGhIORo0zT9l0qBsV7xXip0uiDHXiN8YUd2JBLJCIHW5USRQ6ZYHj3jfdVkCyRQDcmVZrsKs66yb
qA+qhV+6oK4/Nlv6jmn2IH5mqDzDLZ9suDdDsueK3trKwzMJTUpBGMSUVV3sp/f7gelHBMoOwnPC
uKJfP78VcMn0PlRdEuKAFDs97rW89Yw16MVrq9XujdFdNJTTyiKiG4tyFSTDphxKkQ7ijD0K3T8O
QSmxswNDcrcLY46m7JWa7TtHqqB+FYVB8rVY9OK+OSABgkA32T3nTmCOEb22M4UuPSudYUD6q3dp
JmDCQN+6HdfAOb/TgWoRyr73RkHLcg5F+bzgkaE+ZcO+4v1cxs16y8inMoDofdyVBES3lZDJnDlQ
zjl/+VF0UaOsAcwDZKPqJA13qGYbkH9dGdlNq+gLgnL6bKWLN51uRDJwaLdwQsVY2/7cVYpe1ejz
qQvXAzHovJi7Nkpu0dO41s2BcWMXXKe8vdstdtANkvjang4VYehwPCVQ2LzbxALqozVsSzfO5BRR
+9NsgHcyV+Kx9UNb4Bn3HABj4ykt9paWFub+8goFs4nRHuW7dems6zFoEbFa1CRXMXmhxMS6oQyG
4p5TJQO5FFfujKfD9hVS94k/Y6lo9OGouOO3JRGBras0K7+JPWXrlzTIeIyVlmKm1t3Vb/4J5jpq
QyD/ZjB/T7UKRhdTmnkDj2830AwqmosQWZJ79t9BHpF6toPlxpXzvbVF4JeTydQSEiKDARipRaxv
Rt4TCEkdePep1XQ1chOu5B7U6nKpoKpj+VbeY7aOxyx4z5DptRjaobiDgK773ru8b8DR3S8BfSKm
tPh/U6RDTwT2+AndOeJT3uIw/pIkdvzS+cMuZGeolMd2LsxNCQuU/ixXaUwrej5/JYbuuDJQnfT0
CnufMPljkLuiTeyR5x4gDLuGVPgl08IMCollt+EgFChx16U7yKOPFhNWS+wEe8WZyYd70zGfqhrL
3xybFqALVH0xigeyncyLbn1QRBfqhth6bnhw9ijlsHn6ALD/U5z2Oe+r5pzfcJYt29xe3Eud66fa
ini3yjcDFlPs1G8lC2VkcVp0m3l3iiEUXF3iUfdSnZKI55Cbgiy5LY5PMnhE4H0ddNC7svjnhP+a
xDPHdaezyYI1lMmdpRZpTbOt30NybQgZZyt0unIexAOdlfUp3hXNT5cI0XBRAS3LexWou1QuwNQp
RG3zjIFehRQ0umU4xNvvLwF2iN1oufYaITcxhLr9WfA0IqrKjCGnQY5Z7spfrkcA0l6WhKybQ43C
xbvWUjdcioRCi9pg0YmxlC2tbtGbeq1Lwz+28JSGVdqhj7QsKON5RPgwNXC/q2DjrzUm5U9ANlnH
yVt/22RTwC1vUUDOrO65ybOooPFSDqUxxdr3AQrzSue3bD9wKHEiFiqobXGtiXBD8MgdowKPewaT
FKlLRZ5YRGjroYhdFIPqSH3kkz0mcXwhdLA9MIbQtEo9PWh9rAdS5yHICZ2uwWYEFfNVPiWx8+jf
NgynD/gazAIdB0y+oqdC02z9kkSnMm0+2T0eLt91XYtBqouIrJUomVrQ1WTGc2IU2hiJqvwr3rOu
xTq7R6D0Vp0qrVpEQxVUS+rjVrnO8xV9hFJWRb3cIS0BUoQHsP58sQ20frVZDR6+q2shxiDuS2F+
OIV1fjUXYnhKbs0yX2AQwDgW1JZn9eYAFRcCoomAN1afvfOzS/z5XaL5xi6d/k2OwE3JVsCbuHY9
+vcSByWlqRSpPaNVC6beNSvo0QGyvbC6qVPkFLzyhBugKVzX0LYIW3bt+MP66hqCCrmhZycHVMKb
nrVPjnlfuYhF/8Zrl1bPccXrMHXynoEQGk/FdE3tjlHhHvX4YqacMPD2V7uK6S7nX2bSz8sSxAGd
NgQuXcIZzuZedHKaSTGQ+hjfCZ8Hvdh2cF6QyAwmPMZrEp7h8Ucan++CMHyGLR+6FiFiK1T/ox1W
Orc5QlonkdKiHELJltNcWKa72YUFLZ3lkF6BuSc/hw0GjeFSO3FZrtI3M8iBZZZIoc5xcT+n/wmj
zY8RbGSimGKoW8na1mAk1WfXopkWZKr5aYKMoF8UnGKon0kU05gRoOirw4k7ENYTlrEFjOmgv9jB
MfpquPUyPF10Ee4K771/eyuTRnNpcKO0wvIvxWYkN0VpmIbUhdcvGuuZPdS4SDo1X0PlXtMHt8DJ
Otbv8+1wLWYj2m8wFhvUupwItMOqV3MWi/gFWYJVBZWx1AVB1XDZHi5cnNzvuz0iwiL1uShx2lyE
uVvSIaKwQOqg24sr27h3Wq6iPJjdt3HaPSbW2aRug3QXTV9/kS2Wt+sPK+f5JUcq+5N/myEoiCko
5C2/KKm6l6VddNN4aYG4lUr3WLeCRD4pUb9KpDhWWsK0aM5b2ipfPxhWUZMC0Liy9vvORZAIa0Dt
K3dR6P1+OVe9QchFm+M4jFWgulEZCjLbY8FPM8hK1qTfdkGtBnaBN9isNta9qQpanzv68WY4IONh
1/otlQIhh0nBJ9JaKhahzOF/7JRLIIijeaJUky/gUQtRlwf5KT7p00c73NzI2F0Bw3UhxMA9TAKL
4NySD0QvChTxRKoKunhXyRiLBBq5fZltfndCzSkKkaYog3I6nPuK2Q2SNrcCfUOYRtzAEgHhyMIk
HaECp9Msxxkn0z4KpaMs3nP1uKyObkXy1ap7fyiFCC/ajM6XZbre/BZSU6hX00IWB9VF5Ufryvh4
5973PCAoOi9b5ddxz+J90dshDcENkeN1srfLiCK9K0Jw4lntpAeAFdaZ+gDGKT2nz+7LukPThYTE
2wTG3zj5kjLH2gLOjlcN+s6AonTM1eSyS+/g8ZaRgh6k0tllLXjdsNcp3vVnMIqILj0Fr288S2qa
3Iw9bZOiWmWIXmpT2KboM5emg0OgS7XNMhcpwLN13Zr9BA/2544QsN/1J6s8YV+iVwj4oYVqW2kw
A1RKkCDqhoQZlSeLScVpb4F8hPQJ51xKWSaAx2obLo5AIz7hi1IRBqdvqz4bQ+tzY1zBomwSx9Zu
2KCoJES72NxnZFvM+zSpAiM7xg1r4xjVSpntzEOodZgdC6y8skTk4d3KKlPnuC0+K2VlkcdWL8mo
hJ7+gp3Z3vqqlOBvVWVydD8spHxn7fiDNrfqRAt6BALrPGWfBy1QY8i6zR8SFSoIvbba9zWNIHVW
2bc8xz8YBhbXmtbB06Xy+FmhlZjwxYBJjE2YmKkCoRdd+oGAkYqAC5InOORsdIdEYpVXTc4KODjm
EBkDx4O2epB4FmBDItqn9O6TF1QoasVSXhwGpukL9M6Z3n35JRufPNgRtQGDIWfvvqK/2gH9ehWI
EZJhXkm7fErzQHAQAotQNOtgj7S2/YWiwmyDCgrOkOSDRoepCfRal/2cfKDvKZxpo2A1pIIwjvpx
Cjg8qghbK4HQD0ExDeX4Z4KE93gQxBsOvLx2zjwn57TGX+314WZjNVOuN63x3GPjVhk8SWX5HdE5
FUaPqvmECtUIRLPcEuqY5CzFdklhv83dbfll+MffrhnmW75glXE1ScRiu0vAwLIbgEnPVGd74+jN
vmkv8xhnscNB6JgdSs0wersaFInEmR083WziCZPdCBOOYqrew4IMhYt9NiU1FjQTZq9iGAUVZjtt
Ac6YTHAo1uu0SikZv0nc/kRNObMsTg5fGj1XQmQyNbbaLwCK69fdDh2PVC2Vf9wgG5sIehaxM8DA
MGcz2keFR22Ck8Ljjja7TBEXRnSuMiPPLIxVSzLj0c1kXC7qZoBs0zkMT73O8RwJeSU4szv2WStw
CW4ZXnEMOL77h0QCHJHr9/50Zzo5A0nzvS4pqaMW136sVnJRJv3FgniuPbprsBEOAYy8HF5tZyDF
+K6AwGrMGNXU37WaAz8K8zO8WI4x1bIhzOTKafbVCdtdN5wMS2e17X1KRRBh77A3C86E2Na0idiF
0tPou/sW57qWTHk3XdEGtRAGCm5W4XkySLkdAAaDplV+k+iwvdp3aqOO8JBKgRUfRC+tV14vtn8I
69Pt225BljYkOUJfPRFBRdCwb4a9KCodk//jQnCPsp03jLnplnAzqjKiCALg8imxjtBWRwhiUug+
V00FTS3srtJg08HIThf9A6WkJQ/pIqUI5THB3vXwnnpJpadMFp1N7pJrcPJhPF9Gua0xrYZ02DCw
GwM9XWzaQ6gbwkvHIcokcLMmQhoZFQirZmFLjSHKY3xfhMMtiMvldaCMeMsIH8LoW+eBWUguVL/B
J2HMbONMsFdi4jDILL2gEtOBnqbgcEDlXz9IajLG9oDY0v3j8Kv2cU086IqUcPvSKl0xmCMmNeJ0
+mcEo5sUl8DbXiVwu2DihTjMc7AD1cSV4ZHlLBNk3ILAPpnh8wNfuL6fb1FPwu6OqV9JphPDLGXr
waBZyoNAKsAAPelwRVGly6BcN+mRU+5hi+SDWyv6n0JBPhWTgXhGP7RBPlCpgfBUTvbWCOIditqA
zmzlWoRyyR1UOuH5gzYNF7vORTQgp+pUtys0gIesaE3vl5W2X6Iki3ug61oEgiSIGlZmAl1fXwGa
o1ciUyS3cmBOtH4hKJEUvqTJUgkOfCguh+RHSNPaKFmuaRW54Sfbq1mrL08Igk6F4w5pzWuiG85P
McAjydwxGxlOID60RjwancS2yso2VxP6Xqeith/8VNhz48BFQPOtlpPdb3lyjjDw7L52sFZOwojs
fja0ajH7xDSOJ/g0YEsedM1pQOvTJ3Q31u//lbr+CY587ieYvOk3Moz7wvg29lpkWtFtIc4uEEIa
2XRJlh5XPw9xWuKGQVfz0hHWI4kulbt9Eu4wHEUNC5kbNrsmNARTcGFYZUqC5hJf+teQP+WyJsJw
jK0pjinmyeQ3rhJtiKxUcssUvUMqB3om8zmarVGNqybV5hgkgHoXY3j0wN4mND/YGjbkRhMEikgr
HcVQZEM0L30wu3u5o83E3+4Yey5lvXQazKEU/NtGezhJF9bRDZoH+2DLZpdLhHIoIkxOq5u2qsDM
FCr0zNEfsDoPQf+hkoc32Ccp56dyeyIywWDV79HVAP5TE1AIdceU/ZEBLjR9mVtl8OGv8hgEZ6YC
RVcbKCYGqgiKAUyF+JW1lpYjnMk3TDARigbvDYRrfODxg2qYn2gSQ3A3byD36df3rpI5nZSbJjVS
5vSJ4KWQuN+Z2xDR/lkOJxsFisiQ+QTk7cZbgxRMX3Hz85pR6O8824GyPafCepv+rjPVi+3NqFHW
E0i/awpKA4MjjgLt4C2V/daByAT4QJbuwmsfISvShHaXnSqd+Ighe7UOh1SAj8xk4KmD0u2PK91v
HgQz0DH14UPfHl3al7mzRrgjWdlbkl7VySPLhbJ/0a6MnsvmX4WVPx7+aP5PBdq2aBydNxbMZIUo
VzVbCme5rXGLwmtDm/F7orlWDDOXUntv12hE6GO0/Miu40UH1ud5/ri+5IO6OLPVCtl+ZNwrScpu
SMaSpzEyUr0LbbwwBRxrVd9RjhC5PoEGACaAbr22sSXTjHbaYPHj2SphKClyCP4ZRLQwqlxfkldS
lR8zENMGWk/DydM5eOqYky4TCjmYeK9qc54uCAM3izJyyJV4jU+4EPaVz79XXsIrh0KQ6KMPHdwG
UmBej6r0C3DbGnHLNWnpc9/72TCGze/kKqpsOGM4zwjOFHWWqdRtz3/ZTxfIZmicf3qWAe1QzJDh
xnys2WEPuS/ODnF3g+W81EYrslzR5269cbVVff5HmFWiGAwkgptGsIIljSlRgDncLrUksCwkYxZQ
tKMHRE5FZRUZXyxVogXxNjOCsBupdCQw3KUWepBt3rzXKShP4LO7ztHDsGF2PeCQU5JTovPIrZaq
n4zFFDcALA7sSVO0raVY1ekA3763le5CiVZMYdt6GwKwMGlC5q5If+VbRKxjF1RRNBB9Wz4yDRfG
mWHAly8H/xwLGeirHxSAXLZ31WUN/X9FA1HcoFLvtjJ06SNGb1FMNMHxjbz1th/citsBeky6JoKG
ZInpgUW9D2LCYW5Dtdj6WvK/z7XOz4u6b3Nbiq62I+NSPD4jszWM0WMInUTs9LKUcocWmu58XLEV
CgD3uUb6rQKxiWxmuXZZV+X8z6D/Q4Gp0qK9JKNm34QhuY9Bj4EwfwcZsmarBD12+xjaCVBHPOUb
+6wWJcuSVYE9uwy6+Ph29/VErJBE5r7EvmqHynhhKbAFaQEtRVLToo8XMqZJgQh5kNfqzIFiqQJu
/eNoHqCPnCto01J5zEJno83pKpx0qUAVmRZJ5hLXvXTfcKd6HlrS/awgZsi1Gp0mYvfiupViXBcS
gKU8veMdQgvtgAP8sHk2MdyQx9bXcRS+EfUCV4zaojoQNqgmYGPKwWMhj8SK5xxnuE81vLRPJbuj
daMt3syrF0l1nYKMJEaC7XGlHjWltUqOnw8qJC8Gp0vw1QSfwb9wnlFfP+JlWpIXYg07zPrsp9Jt
ORin3HC/D9IAon79IlzFHftU6M0HNjHmvjaqr/ldh+1k677bF7268oWKXxmwoD297iQbgmMlyYZh
RUM6QRhHTskt/7TC/7IX4wbgnVYXH2JWUaPuxSuYLDJr/eZqvzMmOWdlEp/1I+3xR1oz6SQ63sfZ
6j8vkbiqdauZrZTw6tgRlDf0JPeqbaUDPWYj0jcBetfOQ/W82G/MqGnvvS7QrstfaA5ni+B7Eb3U
sJLY5gks2F9sHWsPhQYwwEhAdPwSNpIQsFuw4G8PkUN9pS5igh7IqjW8L7glg8ZBVssYpd8Kw7DJ
hPnIHx1HMGqp2YUM91BMcVIe2EbtWwrCAHICAgpRb0583s8puT1L+J+IGTWRZ9lKfL10uSAg19zv
x4xb1BdTwED0vRNLSGQcPpZ+OQZQl/BzF85JerXhNvR2Tw4MzeaosJCiwouvuY6qWfDHtv8mcvFL
8hq+ByVN2sPbEzXgbXxk14+rKJuavlL8tn6LDCC0H+nuxwHZgst+eGBiIdUT/5brJe/w8QbhSCNN
SGzCmQUs+1/+t9Xw9Nkjo4O+sgxG46n/wKbl4QyWkLQwLOZXgqP+ZQAikjdaxsej/tRlN3KChO/c
lUrv+gUbFuTcNtzTBiQM8vK89ofNIxP8ejLzDEjIKjB81+fwP9HYFdk6bM7SQ7aC8mw5b+UnNZF3
xS4DlqdtCa/hPY1XZYxzONZCLMKH1wfFBYcV9S1dBjcfz0C46QqZ69BrEep+WqkzHD8QvM7BRFqq
Q2T4DIpjGGosvR15zA3tZkpC9YofeyWreKFQwVEYzgfUIY+qK4jSMBJi+OyMOSFZ7saqx4pxQlci
fMWug7myweuS95gg+AyWEpEevGKI5TVBVActDbEst5JJA6fBYqaPr2vnlpPHWd/Vpjr0NBE0WvPK
eYmX2ER/DcEnAXmtxhTMMb7PnowSiVQ4mG9uqdSMrEGC6SY8VtNgYR7PJgDLLhNn5WfY/sx+psC9
eEHbDoJ1699+vNDoAoD6+wQJA/6hs6Ae8IcC2weAtfRe/N/qUqn8yv+KBtorAyWtjoLxbNMKwbc1
k6SDp+cWNSrrKDQ8kanKfIMvaqt/c6VJxtJE03yHqWt/G1oCSLGUe15kKb0qk999ZfQ+EJ5U4/DR
EGlpzASzmkd+qtUJkYaNzHzA+SnrHgc5oL3s9Z6ue2yN97FfgtiHI0jZSKPcRwD939k+22aMkiyi
g3gXQgNSEQRJHKVUG9KHxeVWE6xkIIlBS8vy7Lu57rEXAPu5fvXXchgFEa32dHSenWeULMhtaGwM
D2uHh8BXVFNzDwxDUjxSQOkU9PTvuR2NCBmM+jbk5IY8K1O07CHxwNMy7ahgPokAgR5x0TNL30cY
qE63IdXDZbnSzbXp9dvPC3WV29Nqj5+ClFj+IfXlaKw40hqkQQW/rhiqxcLZuqxrnkQdnMr3n06o
C773DaxPejsOUECLAD3jziprf091E+WqY/3KZPPi3ZFnYPTI7ugRG36V1YYmaNHboB6salsc/8vV
ijeVsUCBUncHSaJEujr5o4uUBnoxndNIkiGh0gyobpcbOPdiYu8zSOacX4eII5tp+6viK58CtBwK
BgSiHMKBZmzulJ8Mz6MV14lV4eEH7C/TrjmmcAM2KX7KbnPPf8L5H3P+itpP+U91YB8DFxrMZMmh
BYG3Af6bFjyMgqHHyLEsToRc0oSxbXi9W5G6dWZkS7YVUWTXp5WnIkjfAn2oRQs2nB6uigJiOv3y
4eGL6MaTaPY+E1cUB8/3fQOesNqOoJkPG1ckCjl2PojOwovaquIgv9wBafuIe1WN2XBgYuV1yYI7
puzbpTUU8M7iwKzMohEns7EQBW3zvo9HfYH5krbofyOdvTuOvRcUrqD8hvA5KiRodAhHXUJlJHZB
7XbawHENc6drQOxdbsP54AxU6VQoH+9ieJvM7CqsB9VgJR8j/ZNhp+SL+aEgOCm68PJzrvLWqmEL
Wl/wjp2wUDwvxH+q2X/GmL6Dw0/4OGJ5yramryszxsySDy4DDctlcOX3XKcy1B/Vsboc57uXwmsC
I1DwyGLW0H6+RB30bKwWBFyEyhfedC2cx76XOmHEvxu70Zlujk8cYUxCDJdv2NizeBT0KUzjAVSB
QXPoiLK4uDMpTJ9IcevUnAPLPMRdn2b2Hlbwf0kmxkuz8xEe3ggbakKx7V1cSJXzjpB3LjO2OufV
/Wp2ebgFxSk4NJB/kcWGTiFjb9t+Z1dntk0d6h7R8xYDlHZ/JfakAp71XOfhQZ17L3N1jsKQp2jZ
UDt0Pz4mtxsyKQSg73BpjrRcVs2Lq1XTgVPUDbNadMiPzlWrbzOiiYQfLEKCrc1ABzoKzeRIeqxz
UboKmZuSwVDVRRwKEs0vBslJkhbd7zttfa2LP3ZCnFkzZ6jOwcjilQu5IjhlMO1qT0JHXUTO3XmY
9pMv8hwnM2TwgUKoGooTZ3U/ee6rBHvv3TSOquJOgyugDoFlvRL3u/TGCnXDdCcVzWX+DXOJpZ67
nXCIMflVARR1IBreSY63bpgSkQ7wBkJl0fpX+oJ/5W9vouJUKnPub5fa8V42eu+ZxPNFL9/lT/BZ
UjRlZngpLo2UfhH+T554aVE5DTFJ9zdxvssAy16jNatmI92b+8cc8xFS7HqIwzAECg9H839yQG66
As0vAWCj/XUgHpLFyQPCqMIYnhHTAYbWg6LNUFRU0XSXlh6zAncx8VnsahxzUVxy2DbVOPPNrQzm
nxZL000eFtPvK2mdn2rTawzWzkRcvDNjEWIiY/wsTbjkRkge9TpyMglxAEEu0W79V6qyON8YdW4V
EsVmpX0HSi3g9l/FQi9lu1xvP0qJYxS4k8d3eqp8125YQCjni5AvTKoarc6QKQJ3rqyeD5EumuDM
yabKl8/4zUdKuP78Qwgr8mFz7Goeb64CJlvxnZDruaejo1+X8ENCoAwM++q9jP7ntCzW9qomwbuo
V2zdIIu4SqP22N7iui+isD03GlmRp3e6FBCyIa/9wCRf7mrANvK8sel6E2IfGR7jxPOuZJwAQfSK
z49rBZxyFjm+jV9aSVa1nq1oYthDUtOKZRZdjgFUtL5XG/YYKCapww+ug9fm9Ip3h453XfdvVKn9
Q3x1WO2HvSirMyunvk0x9MSzaNbEjQhTLXArm7pkurgoji0aol+9pV/QEV+7scLXEYaVuE25BZVx
YfZREMzDXuTcmD3UQdrYp1eUQhcooOY8o4LrK54bD1iL17DUoLTb0tJxDepyO9irF2+caI1w55BD
BfgSdvEAJPDx2dJR+O9yiKG5LpGnAB9QZBPZMesg+sDyl0JtiaNu9MoHtBz8nu6wYHSZTpAEN40w
PcLjOKG4cr+fERdcvGy2QhsqHsKA28UN0nHfSkOL/2WENnEa8abHOJBqsnTQmEwT0VR/M9lkBlsv
vJeBmbqJtANYa7cMg6bp3U3tSE7+4XPJhQneo2//lfWern9j6ry99N8r88OUyPdd2/iygOYfWcHG
9VlM4aV2/21rSgy6xg2iwspWAZyBjEKa19iWfYE3YDTmOMJmN4Xo28pKVicoUmKzOEDd/rcqLiIT
Wath/OrUgNttigH100gOmxVG4o9Wg6BxRTqyQ7TsqXcx5IiixJ8+zL+qSjv6M7VztsEg/OArIeDH
gtKkOrdWGWRy/WCpkr1yMJolxxnV6dzQEHZkk3/tA11IDP2FTN8kNF1qM9kAaeRVG6kZqyfCGs4C
HASGzxBio6boxI7K5jT/tK7mHrbyW14Mnnv1/3lcX1yjVLEyrRWSbk6dhtV1iU9dX3jOqHP+0Oqd
501/FnZVng0da52SQbHtbP6bVOVdcRmj1kPv9AZgdaHVjYq6dh25rsDpydOobKHJClZz7/UtzNb+
Gwl2zT0ZOOa50spXsgSAkOI1StSzqzmebf6JuaoBXX9nhHaTk15ScrdenyVEzeF6lEcPA96qo2ZY
iYrwL38Nvkvtv6rLy7MyQIqzfpd7gThdEk0bVPn5E36rpYh4lzrk0IcanwfRjyboUj0amvqPZe9d
eDqf6VZNwBBMX6TQ2Aa8MopKKJwtuTKRxkV5f5+6wU+wjyYuamP3mcV/inPqqrzOvwK6eTUW/HJB
hG211JPMBmHdwxJvORj5/VYJvY65QKRM6DRY4GE/BtgBkieLOBtnCZvvEYGkIZXT60JTRXwokocA
lwYM9atTP8+gJF2CQxKhw2sdZNpCfgfS6U14d+tywJRovOmi8RJd5smOXv8ld4hR+Yl711vWyRQf
oOKQ9x8BipJYDMutB8KYluOeCee4lGLAUD9lTxxWVzEGsDYV7x4LInpTssbjLSSetoisaVIoRx2k
1Q2X7NHy8F0YjrhX6Bpx8a+fOil+AR0Sg9UDxF9PISr3Ism2c9uoy8UpStykb76RTMdtMtNx5Wkw
KWqlgP4LVka03vG2OpUQNfjTaz4ozJO8huVvK4TtjFjxR1Vjteo3JcJ7vz9gLb1e2uLYzO6MzA4t
17KGpjWw62zMDCEqWoj3A2axnGEc8nk3kE8blBUfQPrUy8VsRCvN4CopbEZqv8AN7Ks2ZlCwUgit
39ywn9QHRUtgYNPPZJoDHuSeiFHqDcnrgLAD0CpORnlQ3pK7ykZzezfCKnuO3j39g9McvlUt5kmB
lid7xIBibRH4Et4+ljELVh5I9wG8zB8QOwqdot+jEhUCRrtTcdh9jATW7ZUK3nrraRu/nQdEzWjV
qOPEcryim0dNMnJzcZrtmGOa0aV/ImCKi7372pVszuSOz3sYq9sMzOU3keFY3TEi6Yrk8ysbsAd1
EBdAQmmQf1HXCtq8bg1C5WpBpRf9YOdRPKvVmg993fcp9+znYXH840nqaFswPPlEWsjYaghEU/rj
15B7ZGNsf20lfvYZjnBSCuupSltViBCOThE3CDI8KGatk2Ix4m/WvKC+4GxXaK8K2cDgOfe6hTCZ
KswU9Q6wnmbqmjSLKON0Tyi1yHrmQmW8Ds0fN/gOkVTztFbTIOzDmOvpZeVw7eBjFwyZwnjDeYW8
KK5ia/tgnR1eU1OJslEryUFu/30scyRbHCy6gDcvzxqi0D1xR3S+7ejghgs+8AHRwXo9eVENNAtV
S9JmiaqqexNa3dxqV6bvDnpalZScSBNLiaAKP6kEkXDbjlkqy6nID5Je5NQeNc6OzKO5ZLiz1Ga+
tj0QlYp6OiAww8RuAcHv7fRGqAIkIrEpm4gt3gJZU9dQRvF6h08jd0chJYjoYE5QzrYvdtupQuXG
riL+RB9q5VELlF3y8zMRYmzkxnmAHRbYwFTx0+Z7OrPiBEcqezZK9V3AGJAx41JW1nE27L2yuM3N
FYSYx3oc2nYyF8u77zSez10DgId618d+dM8e8+cQ03gxZtwWFkDj+Wot6846FqTDW0nWN0RrNJWi
SWgBvGFePxtVzg7Wce0ONpr4U+pgKehOujuLGia5ciMoH3MhP4Bq3RJ7LEf29A373bxlC+TKlbJK
/xo6Is+Yio6oOvixeLHAGBGx6nXT3RIEBb6iW+Bhw+6T9BAcSfBq0yeqd6XGQ2FDoJ32TBxXCX0N
9+XHUdRMb68HFBKw10517TiIaynDRJMQSR1RkIrHeiM3O0Pj6rgGFS5R+nnXy9gseAeuRjvtACrT
ynW54KcN/c3MoiwL8DMN6L5TN7k7wcar4pRzpsNjn2myBUwxh5KIUV+9MmGQSiFFrQfMvZDAloCl
Q38EwNc1tN9k/MU8vj42Ezk8rDlRtdm1xu4S6OI+6NSVWaKOxTNvgss+aJAfxsWeqJH/OtluwKLx
YbQc2hoz8whSPE88qGk19LUjrDMtA4Lp4t34LW1V0DQa3GrY/tbzTYziPNGhJEqCGPyjRSMTR1kG
MBWMl5Soz7cqFlU++/NPBZojnn+xBmaxELhUV/Yi5NQrY8XdFMfr9RHM8fjkfpNdFIdlg1CVOipD
yWPaeofMVoiJHMAvjB8iWQ0fsRBJsSguhD3sGevrkwofA36HOW8lU24l+E8irKL8XxqAU8Ff97oZ
a4snvJimNOWG+AqlhSHyzjcGkk4P+yz4dWtxYCJQ2N0LYRUEeZlCCezSA1QoXcQ15iAwSD1B4TLr
pOBpau4BeprspW3yolmqUN4TazbYybFemWz4ViHscyJvxwv8p664ieveI23LVQw+qsaQ6UkUO2vI
EhdicK5VuBTuInx9VnXNGi8JS2ntDBIK47t1ey6rumDW0hnwbStnt3JPp++SrS56+HMEUqaz1ysX
Hg2sXnu2IdDJNo60The55MCxPWj+BBfY7u1T9/u4orap0ur/TaP31atZ3hK+7UpUzfXblyN/hvC7
vf1KMFPSpJmKTOudm9NG6E/uEm23EYzmYn//FNRaW2fuzALGuxQ4/s/fZ9fAz5KmORBgsR8QYtNr
GsBcxfJBSoVSebvatxAVxfVBg/L94SIZXCtYlFJSTy2rLDy9NwFOBjk7tKCpcNpqzB+ME6lrFJrZ
0cvKKsWzw/9zcJ8ACdWa0H3EkyAttPlPd5PalrBZeiblkmNbZHwTbjNDBjMa8vdh0CWAevktqbRs
38L2uDMBszVIEuzC3S7qCEVsj5ZBrBLnWhlZfvpCF5z0n3jbPSCqDp7vErtVV+sxHsjnofEbwPKP
qYbRI8KTzL6eIIGyqR8YwAQOcY4I5ke5o9e0k584k+qf6/4VN3mGLwOc5pyn9aIEgSulTmXp3SjU
8v8dD/4fUwiE+z2gC76GljVbOCW8A985ioLM1IuLMxGAn9sSSBcR9z+yVjCzczC0BQi/S194XRcI
uplLQ5LrCGblV0wnXr2N36KSaqcNVc9M6zbax+df/tAs0Y/OonaHze28BdZS7qmDZNmtuuYFv4ku
ZtDqJsz25zWmju6XutUZtFpl/slPs3/CeWAM7H132xMxOEa4sgStEg9l0/dr2wBNo7iUqHKHfZb9
BEmaltPY+5o8BmlPGRsUTplF1xsAqbC4BxalVe1mOZfidm/TqtczXeDWQ19/jDl3pW3XvkoBF23U
eC2OM6rjyVXUtFecA2RPfu9s3ddd7ELIxGy+RlCb86MTEEZXWw07EnalP0/brxB3QGffH9vqlkWS
OF1p1ivkMgy7nPBnAPQ+uegCpSBHzAGOoGEw8Kj5SZ2iodHbYkGAulebnY8KZHNhqsxPOpRRECij
P7avyUSorzTqvQiz83zj5t34sKmxe8ObAKZlxKWk5p77hSbRl9A29OZ/vdS3kf2fafmTnTXvNsij
25Zi3HEcdEO7ZOrkA0RbGt1WxYqZmuBfHwXl7MBvd23huhI8kMmMK/m9VTOYtHSugLfWMwYMLIKU
qVA+gWSxrE4JRQ5op2hbBnAxldVuQpHpynNGEBCSEmng1/4aV7dL9nPiUdDeMCC8IPbgV8lGgeel
XNqbpGkSuWf/ET/VE2fpdE977xSMh1/gt2Y+9qHmFhCvMw98bDNG9l1Si7K/HmkNmomEgzPgaTkD
+sbgAUiGgy0xo+kto5bqcuEb9wA+I2Z93NqmPpNbWEJJkguf3PwleONJQhOcH6OVOMzddw8Z9WTH
e+6kZu+DHG0FK1bkXBOi20Y0kGdmcPx11yWRPS9Z7t470tACX0KrXbkoPF03uvkdK8YDEKNro0d5
T7raA0DPTHiKuA3KdNolamdUA8FN3XjtqERmjkPBKt5GVTBVksDjXdc9ojBBMycvLN7/psLVY/PJ
EoC/N/KwCjUW65SxYxKXVDlp5XCoGM0UPVgr2PBQfthPIHXfq7plm63ifZ36PjVVa52VKm5VkJws
3oXzaUt/iVOZpGFvxKpIpYgyc0z7EBnmQV0mYTCI1lSFQWu3qapHtpQ4Fjtr9nNXIIg3PPF0ha66
hvCxuYARXpOVq8GH3mwkrIttkQ4dukAGZzTI6YeyIQbisgzywwTmiISnhQ2ZDmU8lpPfqkabf5rF
LDrCM+SJaYjZFARUdH/Nf/p4h2EHG76eTLyIrpNWRDPDM2Df8PXsBsFUbIAsAqBkiv5S+xP4XKYy
/p59kf/A9TpT9JBkwgk87bVVYEdmORfG68p1+PZEfY3A7FHbzZhv86LQzxas5JESNaRiJtI6cQ3C
hqKLgJo3OGvSCYQ/4DaJSnWc84ph5jbeThvJHGuNLYWYWMNzkwm+nqJcWv3eVvzyFgFMuo5lMROE
MCUD5GsF0CJOE0258u/jj/vF3fk3vP1zCoDm6X0d18oLp00ndTSl0wSmVXPOG/LjhCoWaj3QvYD+
gXUXEEAROwoNsByopgh0EgCW2E4kKSF7ucxDsfJ2iruwDWIJlFk1ncakNvIKXSSV74SyQ9rxQbR2
g4NzmYZTSIkaNdw17rxjSY1WzNB/ymhqwj8N9711ybM5mibK38vC1tU3RDOU3kAXhtW5WkS/CehF
aq6W1cqwKVccYFECBs+vX4EJfRL/FNT7kS1UIIG+4/IBlSBeK80kteuHGTpVnjqUfwcMrqUuyrSU
LmJO9NfxTY/vep6xIWrX9vhib+aJUt5ZSuuKdk6oUBK+I6wTJst5awvKfgET0XWJC8LNOGN8VvC2
BF0x0d9g96yPb9nu89Y4dhkExwIuR59TIR0KMA8Hcob2kOD4FZSx1O2LrcoVKgAs7BFHd0M+n1Ea
G3YWgGKJdPggfVuf15KAoOv4lQjpHqzYlc/7dqSx4wN4dC3m6ydwpadOwRQkKGu295lhm/wle7oX
rn46T+yuLrzy/qMcjFDHzBmpV2rqh9trZeUsKVaagfVrzyApwdwYJIRQGL3rE3X8/ArT2c9aZYpz
YXr6DqP33epv2U8HQC0iOVSdiZ4V0dYv/QbUjTrIPTHz7s4HomG5M6r8/IE6i/a46RPBx8kRkD10
NcNa5DEmy2EQTmIkhLYtHJxEs2q7GJGCp/L0n68MbqmDI2e8MpRVbnUKEnJk5qJmhamcJSkkSo64
A4NW26wfjg3wJ0ulJYGq1TlKPJM+8Ujp+/eH02P7yQ8T2KeGec6IBHCeO5Xoj1Qd6OKUhHnKlAk1
HxQSVq9tWGOvuuwcVwqX5frBPdykGljN7gUHk8KbBK5/hoWY+WZGBzx2A0l70mFs+6SFCE2sUIlo
hXt6vthXLh81ZeJc2JIHqIZZT6UcpDy6froJVpEKWYYgELhzUbOX8/WIJhg7cCPZrLPURp2F6e5J
BGmZStQUKDBQTQ8HqFMgnUhOl6PYiPJSR++554UWUbMU5zPl7BKxJ+kEo2oToyI/3+pKht3gSAey
PgJIenmxv3q9sF3agIYxP1h5+++Gw3qTaPPz/uRKB2lWbpE6hqOxqBhG4PqtPg9pIi0NDax3xiZM
MwtNXAGfEDfXMW6dzmjv6xO+UtPBUKFdwLnD33BmiqSL06C27UPuVrSzFTmZQDnnVRkFESp0cwOf
2un9M1yw/y7MUKcuQ0lY61SehYzE2e0/qRRUprAyE6bHphutpTBy75DWvOgK7LULnL/KCVLnczm8
fANaFgD1p5r9xpldGJ42B2lLJ/FOPA9jauM01PHkkxF6mpcFL43eAFULpRN+vsiXl4HRVqNxMK7o
LB5bEj+/8jygHeZ765IIGX/eO7JwkDnm8FqYlDBKpCNC53IXM2eXfjZlqBG7KuGVJV7c/imgLJrh
E1fzm+lfdWa2mkWp3UA9r/KAOa1VdOueIXtpGr8jLhFHo6CBxhC03KQ8DbcEjymAYiz9wEmtI30l
p3iQPOrDUni5Zxq8B2We5eTikihjp6FV6XLewb0H/tvsY/wze4NN9c38EG0DRg0N7nU2A8b272xo
y+DZXNpn2lNGtY+oeg/N6mkFwAfboaX8wzjeHNoYKROuHVMKzlVCTiMDGehn1ccbGoQbYB6djjLm
be0VX2WD8muweToc7/FFy2VoLLSmXpXl3y798iMNSL6aHd5aclG7d0/Z2cHanPKaP3xgcVqWKvvy
wWaL/sjAJWpQm3ZXU45ycaOGCFn82zy5UyWwpcDnIBNSSrfQ6euljHH5gRDWO8fVW181gvZgdncC
rnrEQu9th0B9dC0jL7ktS+nf12VIr3KL4KmUoq4E4CAIYk4gQbUXvnekqnDiezKvrFcPsz+Q5l/j
b4mdByulqEsXMdpI5zPbWHuBvJDynx/0zHFv2Cgu9NuVK0bPOhNOgxBADaASwip4qKQSqa+oNtsa
dKW9ucHHDoDFcl8QIsOo/0J1xN7RmQcqUYkkOvVzu+6LBuaV5W1h2X9PBpzPj94QmlDq+t/YbeEU
r9oyVZTYCj5NMWKYN0PlTC+66PNKV52O0FTAHBWmAr6QdDQ/1hUbAJsGkvYwtusRrQ7Lcjm82v2W
zKAssTd13oljA1IN7XXow2mAqZ5KGC7nSpimOtV7TwyYlKD2a2MCFj06uhq64Z8QHOg/fUIFvama
9GzPL2n/56FA9/6vi9U0wAGes2MbqE6mLwSJJ+HZCkSgNjJzmVP4GbgZvhlXHwZjeAAaCEZkGu+a
HY2Jmz+Ty8bi+eWjqZnlECOgalCSOr/8iNYHg8qL7VtpqHV/Ox2rR/ZCulXKQ/20tFvbAF12zomh
uDPaXDhM1QSstyiAlL++QMCfwp7eiGpNq/uLM63HPOBIMRS5DWSkvRD15B2K2YFthEZVhon6NzTl
0rwR7Ocsw10L8iFa0TCxRCN9wim3yGcgRMFAVmxXywcp/UDkW3jhsDoEoCwST1HdNKA8OS3NaxRg
o+3cA6GO/hq+n5VsTtfe1JjPVfe7AW65YVZAFVyDuMtAXeXLVIQNqy4lrADDMPktBKwRjMXYNStx
drqBuci9rw4AE+C5VK/rmecel2jNuPVJwC2DbWiRVgLKMr6ju7pIHjbJ3CDG7D+oTgUwrP8/NmeD
26md4sh2tmoPUpcFDa3MMu6chEBOxSJIImFIgaojSiWguou90pBwyPyecgefq9d3vhkj7orizGTJ
X5GDhZtV+XZwM7t1fcwf3LNHtHHSR7XUzqga7bF2yjNmbLlJr6QW2nd67R34xbF7hAj4JLUiyXem
MxMjgqYdTIKYwozJ3C2GvqZieEmk4KQnlwdho/czb/pgKCuXo/fe/p30VY0msPjpY7TE4P+hbtXN
KWu5QEOQ6sPcQKHBgm+ntL2esGk+Q61Cc+CKRuoBnmnwU9GKjfcHq3siEhBM52f3zCCJcz28Rz5i
OdabG8cYYedRPGktWEvxnV7cDNzGl1j2Whr7caCfOgAt91nsU9FuTFiGN/oYPMO0HYvA05WgKpXO
rFoMo0iuctCYePuVyxdQXlYbkNh9SWB329MaAW49h60oFpaDOtbD5N9L49DeF34oP+avlaxJGOzo
2lEAbUlBgiSJAcCggUGwASDANKtJaYuMRsuN+NTciU8J/55wYA1V1X1OUiGAUe8PQiJr7aKD3j/x
uqld3FCFKVbRbRfA3EPOktZeMOG9fbfYKDc9FDbAtw8i/2fjstJGqKui6MpTZJ68esbJNoIvNM0T
BV4iRURgwnNSaVbUqU+f79NisLZTC2XK3yZ8InY76rEknusk4VwIYJuoBcyKFC5mjFV7EdQ91wCR
CkPWQmPnsumkELu1pXKF7RSUGn+T6ImPTrRWTvR3DSV0HrWYDMJhKN73iE8EehYgxN2UTqpJ6EF7
o9SlrJG/mb5Yw0eNtEQ5964xNIs6iarYSOBq9o3oLV0nlLphrvaqNRNjT5o1UbKJzUAfHfl3BPls
+p6vglrXVg8xOi1MaDpJTlXxuhRK0X44RwXG0dUiBqHU6VfyYzwcO+0xazABT5IrbRR4dIBdUPyz
0acbnRoodJKY0XRtbDc+d3ZAk69LrfS0gJuJoygw50HIACQ1wsWbin15+K1G+toZALXSQBO90CWV
nO2Miv+qYgyqMdlaQo4ObrApv5Ku/Vy17g4YZsFXPCE6boJU8keZaTH4LHRym7O07506A2A+ghQr
lfyEPWDkueyWacNIKWXSYPyp3GgkqREOctb2zM4pKptJ/Gc0drkTbJ1XcDEpBPlOdyx6SFRAl16Y
ZCzQbTLsollLRcfMmX0UXLTKHDmdcOzzg9oZoiHws92/kWmHBQPXlsWJiOqHLxtoOrEVtvrUljKX
CkXLAimwkR6Dl4rn4Q4/3wWY+Km48WG4HcdY698Pht8bT0XBc7qB0K6JyQcIj5CtbGlztySxiofL
hJLLEV97J+6DbNSrWN3CQuutHIwvfPjpSoTmzlox+rurnVZjMiW8Sf/VIOCJ7LGC1BqbOb+hmSzK
jx7UWUC9m/i3iElOYr2Yjii1/jcqv18occPJVxgP+OWLSEU8tJilEEETlwXp9wzw2gsuSK7dynft
PY2Nd5zc45onBCSPO1YzLhmqXMx75/oJKr1li8KxTG6J6gJHha3xpOQA9IeFWus1Y+IgAQJnCBgH
STr8+4g9gBsU97eS/6gx/ZNg4EmZXFhgWXC6o2Ma3CV3wajoyC3z5cp8BQL3Fr8JiiB5UlV/1bpw
52z7eh669DIgTu9Q5UPKVa6s1LlZSiU9ExkKdAWSJjl06zpNc9gem37bDbxZvi6k/OXWEpYDD2Ml
MNhXQvlWq2btGjQscSesMOLuuLd25bjf9qXAJQqDpWq7BGduUrrog8y+0L98uXNSK5c/sjD1pLEn
rKNv5G65Z2SNik1IBhbOKhSSKIp7o9qlEBO2DQeXO2ECs5xuZq3GXjwg5xlMtpaPvU6cJUj/egue
TkkO8c89XmEO5wWkxZxx3n0TXyIGM11ko6dbQrxpenrfCEmHQUI0hCP+Np0XHneITl6Ay1GrYHvK
cLPfobiscE9zgE9Yn2Jd70g7d/3dys7l7DFJfFPb0o8ok29mDs+C8oKfnW8ybxdEL4kGmpoRItil
Oet5uYaXMy8dDKiRsQoSt2IDsPBS0obc/CV0e+Us1ZxeQvg/IPm/h1MCXt2dYoImNedyM7fAR25P
qWyZKSGR58Vg0DLlJg7gE/J38/2SgrZn0QrsNeeCXFj6XIdApyfrXXovlIGnuHCJDsEUrqt6DXhb
m3f9hkutp7qSwtbepegFJzcPfPZ23UDJ77ftHRjscq1pBi7hdkoI+luurz/pDLSDtb3FusCcs5ty
++aBcRL6UURFYiWHW2VH0HthUiVoELQhJp1reJIdV+Qdl24emKr/Ug9JdsNfkuflCfhnaBAU2tF1
qO5Atw7MPxGC0gwoYidP4Rns4s2uuA2EpnYIeQoq6vLiwaiqlwtML3Hs/V91dhxcGjpqKDm/7F02
urteOhabYSbEGXBhgNQyOYMQusEsb+uTK4r3qygjkGYBLrnhI1HyKMgN6CcDpKrKL85YU4tn9IBL
naIacEXYcJ6dF/TBWd4sFxbfTT0MEMMTDD9dOL14cy4EB5zpmWCKAhaBwo+Afj+iuqNn/z+XN5IP
OKMfiWg8BxeH+7R7SQ1OOf2dU1EXHBub0YaQ0eQMwoQv+ZQwKP2w2HcV4GkaHWZjhr6v9tiQ5I/p
/drKUqq/PwYEPizBcRv5wpdiVuXdmh4e0NOkG6k5U3u2cf94ame9vEHxK9eITOJvCBnlHstaJVxu
xLR12MxSQja7lw7NVSR5cc6rweRCYZYG7L3LfYS6MSSSBQ0c1YmmujQl8De7jyqvfliJqFVhaisz
Vet35dIjUItbg1Sd65AxE4FU+2JS2KCOt8Uri5sNYQt2RiXjcsBQYkE0zR/mB8XPv7v2VbbwZdgA
vFC6E7/lVAguCZH3u6ZLQeAvMCqMkrbRIGv2+ln2DFolbZ8ZGGGpg730ptsZluyn4x2lO818AiBu
X8YdFtVz2U7axyRV7Qolm/051IRoNTePbAEUw2jH0tqieaKH6SoYwqxJFjkwtwO1QJa4IakYvBIu
wUxxrst3olUoKYnH6AN9GAPpA7Um81AGOLfYn0eV18E2w5v1SQM1aZ7yxf1Jch/mFoe4Ygm1/6mq
MfeSreRBUMGkNkAixnUQmocT079s6XBCsuKoDnfmzFTX12EnqaMtkgx5HHJHh/ENgZIzD5MW5ecE
dkGm2LGdnE/pcLK2ReU/PorzoVVO6QVeWZFXhkOjXt2lFUKYe2DOYN+/l+IJvy2FK6rbutS37n2C
9ZJlx9kcyDk4g1tpwy6zD7ie/v/cntDLMf8CHHoBHdfepDlseuPQvqZ3SRTSGtv+JdUOyZqFbl8f
sEia9VkoDXOq8rogtYloQTObUniqIiu3d3iA42U0OLh46xUUrRoEeWxyDxsIO9dNZuZsgKCoOID9
xks6Pxi+tHiUXZHHfzM2LCrF3kU185wP6NQsr76KafVOKPST2NTq+m6eDN+1qc5NCC/hqzjIGNkj
cs9Q5Bq5GfeUArRRJWxfK50xH/R17O+hJAew6EejCTw0atv+KziuJ9LwvecFVzPXPyUJ7JauG5XJ
8i1xOijyz0D2EDsVUNjya7agf7sdR+2i6fJnJccJVIJvd/qmJ73kA+F+R4h5OwzFGdLVfZcR58wO
UAW5DQfgwh2IllCZRb6ATjmc8owP0tsN/+V6aII/auq7en2vKCwDJXOaZiTgBNPWLfNzetfVcCg/
BYb5TrZTytQcv0net1A3u2/jO3vHktwkfCOvhn0gE4n1PnKdj1zIutzfr3adg0FMZN0L8Goxq5gw
RlhZYL4rT/j1kYr1T5/+kPkDwOtb0K3EG2yl2nvGwE/jSDNfTDgC6a3HdeW9A84ucnqSO2GS3Ifg
PwtzsA/zxxdz2RKa8fKNqdWbpJh5AZkLxlQECgYELfYCSxiCpgsaT/3iKZyoTOHTt9yDUebWnVer
9jOab60wpZYLOiDbTgHSzyOpmEWnA+qXxi7lvRBIoiAiDQTeFkBBsPvlvPk86Eau2AXmrotKQh7B
5qOGwzm8hJUs0QUKMyfMsWKP5HBWY1uHkb48hkEpF/ge2jVv6KFnzaxRtvZuS7TxqAyJUlU84InA
8qotqLPTQBf3+ZaV+w8RhGznDBRRa4RGhu69sgQBSqjOMwasqh79A91FfJ3SjKWr5bm56dWNcvcI
dEnDttuuYrSoZ4/E7J9EDS/9Y22wbDVPeqMWoHfo11TGPR5H/e1/q8a/44hg7aDtZRGdPjSc/UKr
YVmlK53alBNWA+qHI1dxAwrFZa6LX2g5wc92BCWIkjIDKIc+KUX6WOKfSCszaWTL+6uVihB6uxzZ
Z3vCS6xvbj1EVK0EANum5+kujxBY3bs+5sBgOf8h3chJrK3WJkyUpKgd1eoKBBo6H2n2E+yszaHb
4GRBktUMEQgfxlwzXKW8tU3sg2RhCzdL0zdo1JnJRkvOPdZoqyrIFAMeIB8tyTM+RWRMexKHS0py
9PoTrkXlL1WaiWJd2nwe5XZnFVAKGwxF1bt9t3q3xZz0l05wx+oBV+1D2UVpD6yobVM80UE5wwjW
u7ojAKkh41Gc9qsfhdravRjvb6DHrAorIKALRx34HYo/dHEVUkDjmbLva/L3/+VrRgvCqletlQTA
WUKzQKi2kJ1EiJ2Klmf5qeyy/8zCbYTXRJL88MTmAydEDeC7ekRjr60qTDDaWjMjBWBE4aeksQXN
0TIFccuLihHNccufzN9qXExv7+eDu7JkAmmoCw5kwnsk8pmd6C3Sl6U28yUMIX5GDtDrfQN8obMf
wEiEiDNUlQzhOr2p+2sODQvD3V8U++lBZogXtI4GAxUS/s6hCtitn9NNtqzldJ5dqekC+ZKVa6Wm
xeNXziOlsGPESxG6rQoTRPzbDKKEVuI1aZaHZNC2Vw4q+cCAzUB4pDB+U0u84Qun/UvGvw/rlaus
H8DY2bivpsPm4MT0M/evbswtL8hf89xa3figyK0KPqcJmaosXIgV6uc3ot7/ftdPCzv3NbpUe/kD
x1OjoWuX4XY4BUdPHGDOF/m0Tv3VKFldl+dWKFs9krEJv2zR1FPsIHalCJZ2lkeEP1+2KdjaemoT
Hn4WU9qwSeJhWc8xEEJpSc+AFLcmk35p7trZhNvx9UvhmUQN6hzEUi4c/3oDqwoBhC/25EiJpW1P
O2MjVmTyRHPvpYOqxiQ2kw0mQ8yqqf8XDBWHtsErp0dREuSaWrCrfeJgfKwoV55HzQBMSklSkCG2
6rAMzWEqnELEZTHXiLLheszTHxXg83rL0pdebbIpYAgWWaq0LBHJtRpmiSyuGGm/aGeFf1qBUWNA
aeRI9L8WOhUxRxsLIsQ0MzFfvxwdEk1UR7ZeNOIBkYobYQrdbBcF+dwDG67uyXVLqkCwR/GZXEC1
UJi2n5xKm4veoOTJt/GxhTAV4kdzjWuZsndHUE7zssZRbvh+/18xITw0tORVWfUuByIFa5ZvGCDr
9FEiXtz+obdBJXYU3hECKK5gkhjlZuolh/R8WSldlZTO2ivCLi+zU+F1y7YYXRBmMGBAp+UorfMJ
yIXTZuYOso6lIgY819qxKtj3P0CNBPqWJN8pqYmtHYJywgaKeKAweauENQZhTXlbe+eITFMtNPww
/zQorBYci+IuQZJoawfKwof5iJwy/WOOJOE7shVZYsLp6ArhoBG9suztzzOLfrmVXF1NJ8qlK0g7
htP7pg0/q73CBDb81XVGawGNJ4USUaQ2u/LyQ7mryCWW73ts6ijCh/5dxSsw9Sn4/Iu424jsjy8X
ordHqiQjcapUZiv95ODIJRwoBWl8qVnzBWUjFevkXELlQ6lxnNHeCzAVr2fXxv/NWJf+ChHYrOGQ
Zt7FGJ9PvMKk6/XqoNXwOR+pftlgLS9KHXdSXxiZZOcCfmxycva92Y/SjO87zps2bw60qeunLI1P
HCSibcwPWccxrJ3EGOAGe1LHljl91OK2yKHebrFf+ZSk3ovka0DFO+FMzqLskvEjDqs5HsvSWoi7
SOON+5R+yRBsn/Ip2Ow5mRWAENzDR2/hcQZ82WL9jt2UX+0JOZTpy5j89/C/aLVUMfWSAiVACL01
6Lq+r9PYxM7L8te5zgXnFtv9UWr5q+DinftPu9Qmt3kctV+jIbORBn7P1d8tlYvySbeFSKkSDWMU
BnzL5rbfYIzF8eF93n2k7aQd5fQuzIutGHsU+DlcgGimnoSfUiV6zvjguZ+fTBvBPSzgimloR+Ew
PyBwVrFh2kbGeOWSAbw5Hp2jQfcTvuvBVV4gDT8klvyTcALEw/J/RE00GQbDh19NMNU8L4Xi5h2E
U/6PNkhUkpMXalaFl6PgJOLBAeUV9RF/eLCOlDrw+FEeIl1nt4d7GSL1dsDYtkPcoCb5FbVoTjgJ
0Q0/vH38Q+P/VwFUP/e6Yv7jh0KVlAme6EZ8e33I9Fvrgmlw9jKp9WZlOOBuroekKV/y+yu03o3Y
rx/59DErJVjOrkBZb8vtDmKdXhkzGskTgH6IuD1cjrwSJ7hiXWxvUlDorYNv0ujpGTHfqZ02NtuP
ywiDXpPSEj6vw2DjWQongNo1ylqYJ2EUsyZ15vnKYJAR9GH4GPhJ0C6XT33OVjbETLni2vIogeET
1G6UawmWiQpE3ffL+bQfSTzam3y7rl8H2XvIvaCgCDM8DV3y50UeZ1y8mXzm+E0x9EsfY2PO81HM
Y27eQp9oTcNn+ERtu0E4nWn4FxkAhaDf1uphD5atbPBYvqNebqYsuTI42M65O4EiyKpOfHLZ9qfF
+DfiAtD/KIj6V07nj2e1IZ/FP063yJ4Vr+ehSePj7qt2Sp50dNtoirnzk2S6V2ji4566Dw1A/QcY
VTI3l4C5bgmNcJzFeIH2LDyvjBYzXdfHDTr3jJApSK7vNNu5bJI+yhgv4/QAlp4JGjtFFtITRsy8
1xKTyEDfj1aY0ErBTPq7kRrjmPR9jWuUnY7K4IK6choQuFUjjfnG9yxbzVcL/vo+i0rlO478nGtP
xPRpHpuWfKNFmJnyxtCTPxT0icnE1nsvzSAlQ4BBD+Ew4FyXct9q0+UhlYJ/MN2/H76FuVg8bNfV
N+LooHTbNvTnftIdEc9pQ6RFazBlZ7W0b60qJZCLGBXHCYQwOxDxmgNn6uTrVFw8r07zoNrcDVE6
JKV7GQeTOP4Mb9ELuhIukBsfpV9q8ckPXoVdUYv1Bym1CGuCDEcB7Upa79MFC0pxecutKrtyqbWR
2TL90Iq0Id9U0gVNkMyj2LtKYu2MSV54Ymxsq8Ycex9KC68MEGtqX16gjkG5FpE9Kkb8RZADuElS
hipmNEIguuv2tkvkGNLJv65pO+IbFruFDRGTjEpi0fgSQTi7IkkGEoHyWY60LcFyDKOAmfHcz7uh
wvCZVXRWQZACqTRNB/lNNV42FwOAlZ0Sr2kS01vYW5MA9fMF3IupPt/SrsAz9UCEe54Uk411L+cG
NhYk8nTkrPtjS7Bb6waa1LGt2YXa+U0qyVfnvHYThUAuT4KCxnEqkJZyim6WsIuX3GtfwnKTHeKq
8CdnlTvJnEbFFF63JqjBjbVQEZBePJUDzcHbXB2BycePiqywbQHGJ3UxrtX5Aw4mMXTbONbdIQi+
mJ5h59/78cTJHOiy/zw7VniJNNxP12J8jIXM20+D3kVq2PYkXJuYWwPOcjN+4bt/SicExe420v2u
5ImndGU5TnJSG0uxTceYItOwtCKnQC9nhNIyv1SWtxoT8wmBRTDrR3WgXmWxtIbcYGEuLDZ2mioN
cfBjY5a6H4ifSJWBjDRhtpbg8D3LnKz8UY1CcjJjvYf6qYAi8ySqZvAtbIgUGf1kxddGx7773h3V
8KEmFmb50Rr+xQsh2JyEUOFD4et7JbaypxqLQJUhYj1LMh7NAbvTzy7FXGP4z6i2wIkMsy6HtD0U
W4bOm9AXOTedexjjM/iXwXVFccy5+6Zu0YzdKp1kalmh1Xdv4u3CVF6Slwgk8UzYIVeuZCAIBv9k
wLqaY4vFJK7yKYpAXHV7kcB9D6sKR65gKI/tx7GB7nIS2FCvIyrJxyORnicWAcRM7julfKRp/f91
I2EzRNpIyNpSFye+ML0KAmuYifNg1oy4vMneAgmHAMxc73AVtE7zTSAUs32O9vEKiOD1OCEJiCtE
eYaIC9jgW4aCCsrBVCS5Kcp98rSiwp1yoBnz1WU+irlsWub/2tL9gbBWco8MkcMDagDehOsNm+eu
AhX8DGFzQHopeiptql75Ir+Qfd43Dn3gtzEdtsS44qpxgP8nhNJweKkYkRHAbCLhDw7+/+OVvsPq
DuwRCubD6M2GdJPxRQdNF3bkYrMXlqw3lFKR6k4fAf1HzkMtXhiwsTpOalSdzji7bGT+GVhwF6g6
FIbv0DLt36VIYckUzcb+C66jcg3kBhgm31qiMtmtDHcIm+SYzAajlrwlEDogqUFL0z0EzAF498p3
DtPYtsk5k7Gv5+ajfGbKA67KGYiOwHg8/L9rgkhL7M1tVOVJ1VIr9KzbEU1zAGMtN9Z/QiDmzG14
2bYl9fNWFqy5MsZUPdRL3SNP9Z2QQVskIYRzNf3qyQ2KDN1UYxrlIXfodyzxrohGn1Q3VKpzHmcn
Px7MBZKTLQiMuwvRYr3v0KeJMJgB4HcSWgQmkhnFrSTufFbCEZAzyVZSiln8jtIKIugNSn/3J1kP
LBGNw+zcb6WX2j6nYN3caZMkyBiRNU2a0x6t2ChQp6H75eCngIL61sNOCRJ7tKaiJxPd7Gmn4m7w
o3ZSkzPfut4HiFHUcOspjA7C5qFgyORSLh8eGkey3UTaAGpD/olgHvIYuSkXMBa2W5/X8iMoyZrm
Y5EtceJjX8P8TZESk8NrqaP7wwtuehuIl8TZ8BXeWBTfzJFK7QX+JI8ZTuWGW/BYkAGRWcgzculn
46dI9H2yOosphyTf0byXxaaboGSODBWw62SO18aPKo/dvSPDBBQuBtTVqklhI84VTGljaSTeWNky
EOK31VmueB9jtYqrlA1z9ucge8NHBmbMIX1+dn6jrzjUHG8eQzz7ZZ2jfTeTnDhHB8Ib8EsWffyM
K8DOExVtyRi+aSKd33gBGgIbrC926GObH2pIgxIW2k5AY2+X6YvKqg3RgDAgpBydGPjlK+/0SqzP
6eNdS0yqMBHD5aqPKeiBRujWaPcHBtNbtPehJte+4fsr+t4Bb1Qr2obA26k0Pki3kJIB8RQGWmO1
R9mIjlclR6l+etXgLj37zKhP3skoLiJTrWzGsiP2Mj3qCLJKZ76FSfMW6CIStckE6PktGi41HT5v
sreCMGSwLDhv6NPvO5qavgLtO517NMe/NSibqHMFglvsQvJny/2pyebDIggFvqwhQkUE0UfbYpAb
L3DFKeRXTAavxJOTgLVaJcVkxzQZOp65ykaiUqhKyftscyuvBT2ckesPO7LT/iGLzSlkNKuYnq3q
QuhyvOy542wDOImC749Wb16vlluaTRWnDjN+Lyk9s9T0+4p4Ou2Gv+2yTjdRzygjz9Mp0t/Kat2Q
TMHuzLTpYlDv6+BIokdTySceXEJ9WEsZ16BZuYgHx/dUJZeQO4bqeGnyD5MMTQfqNBnLfVjl0tLK
01m1mCpykrH52lGjSuktqTTi/OJjm9hr6ldELeGhq3Yyr1tC+HzBygvo87/d6aTc+IUGgfTv+by/
U38qOaUi68KUqDUhCbSf05i065ygREB6K3sONlNonV0s4wiYD4P93l1L9k/OI3rcZK2Eujclhwh6
No/5+oZTxDK/Kwh/QqclyKwfX32j5LpGi+3zYhrU7QmqAEJ6vRz5FGsQYEpNhujhY5WP6p0pqyY0
8SFepqWunlSyqBMes/a1sFSxcsA+vS1aComGUXCoyYj4mEds8vLvBS3WDndxVytHMOMRgFeuFVs0
IyhYJCX0VoK1VyJMxJ4bG3hVo3YkVIebApBDKoyqaiKDa5GVqFicdT5CH1De7VfFVvf2/jI+Ttb/
yGFhZcypw3DNx5ZO2jzFoOLNjaC1caXcup2/qK5dbaToZXjVXTMn6Raed/VW2xy8rmRzV4HxIynH
nOgoQS6/mUOdH6sbDoG2sjFZHaskypVGk8bN59YCtm9CxSZvEJRyFogQQbzl/k6O/Yx74R8FXupy
aCO9YrTz5xuz4JiUykOi1OppJiBkVi3jTu67twpf5tqut2byNtP28LvV+MyPAiYgfkLZetpDCiX6
GaEqsrWtd9k0seOMpLRmgses9E/Ys6YiDkpdGdMsV3274Cwgqgj9v+zsFfmtOj0K3DXrr/xFTLvm
9bHHanu0LVOhjSRXG5wl2pZRzSVn8WnhPOHHrVHDYGst5GsT/kgJtGrGhwl7SwbPIhPfiDibHL33
tJ4QQWAj38VOCx7uHOAczMNFMGwbeb+nFT8/IkEEAKj9qnIBFVrEO0kxtByDjOhKLaHDovwD/QPC
6XkF0USbQM9cBDnprykkH788F4Dp346AlZt7t0kUzxL3ryQw3bAniW8FV0yEmkND+rpWMFAQM20d
0RX86dotHCGNQ3RJvMJnHIVLEABQGoWEEKyn/TsVANXbgz9UohunhQCGIlpW5son4bx/l0F5qjL7
OEXHgGumQfEINRLxCttoF6CcJEZO+pWj2VWyyHnjekOeIecmjvbKojZX4dvmYVovlSPnQCc5DpgB
NRqCePOLC6rKwYQ17pIhitOphWBjp52YQTKXiwGE3WxndADJR82SIe3xCjCffVhsCDXggQiOxLS/
rbvVNhspjU6WPp1KA323kb90GVGHfa76I6tOa+5YBeuTIJH5AsgJi+XnCbpbtIRTkMBHz4PZqapE
Nd9AA+gNIkC6yPxCr/77fJHnFCopYY8KW7ZqQhIAnv+fXnIoyQmlKpC81xUa736ZDTfAyi3zklu+
ycEFw0NMwUqbKRgguAY75qCq37jBMwtY+VxkGqGssJ39Esabs88qVEbchXyzciQEcNaJ0GZqL/a7
qWjXEP5hYX1FS60+FHE+CnLhoVNBg5xA5q/FET4MsM20mgJO6M7/jbxwAKkEk/EcjSX8APeMfu5N
47C3/B4Tx5NuSHBAkFi+d4XoQe30aPVr8dNZgW+lrkV6kbfXXKMDTbatjlK9c/sVEXXIYxu7BqUC
/HBfpZp3qSaYimdc2nx2hnw/37g+hcw8CNkOEUexBaBCt4D+4tOm/QreGsaLcqPjrVH+MFAroJO9
xcddyfKBWFmT74R6IUEcn1Itkw6Vnp90vfhkcdxL+ewyG6wt7/KPTwokd+hvKj3MBJgCVUtnYLxO
sG4bYMbJ/ZSzk/hr2iyh1CJsMLMeIgL4cLaqWWSGxn9nZsVppdT4NW+C6NJbj8NzGxsp1kR99opj
bSLeJwmUccUzr0gOv4wru6/EKXSvlC3cR+sHJ/4A2O5rplF+Eml15GOJAxjEmgWvDrmrM/nWfEuP
COM8arkL4MbE1eo8X2wtKYWC9aq17pz+T35KsZYRZ6bqF/CucxEeR4cTr6ekrUqNf7INf6q0hPdE
Rb5YUX0NQM95YefkywFM6JueJzTTJ8W3lC4Btc0vby97JRkhqSr+oIxEVJFpR3Pjuo/0RMSn9Fzw
SByuZ6MRdCW2jnRlAS9KtQ9Eg+bEEHpuEq9mP5fOOYX3BwyEamD3oTFQ8e5epz0lnVYjFAsd2+Jh
oclTGP4Bg6sCuSaq5njk/TtoFt7e46lS81UAo9iyPE/cEOI2vxFh9c/EpwFyDGEjFuoDy45U99Jy
x8UhXtlJ4KomAr3h2TW8FsLOcpncTUaX4Y33IMBopDHDqHxrkWynOztwSXbc6NCvaV34LU4i6cwD
UazyZuC4EijRFrBGjRaA4nzchHol7ijYYZuM8S0e+8Zmu0toQ9tVfTdFx2N9n16lgyidEzR+6h6O
EEyUhIeY+j5oJ40uHBITAgbO8g69c/DvU5Dmd0L3WZNOHpeSfJu627ZoLM0WwXB9geeLKw1FUr4G
bbC/VzFRGNV5pFfaoxSWZShGhH/GitD4EEkg66buVlQcQZLy9tKWNC1rj6EsLAePqmKLR/cc/PWR
aVGnwIwf8DQIMbiwrH5bWjECC0BE6sZbusSf4LR9bUQdAcD7oFR0xIrboHuZQIdvB3t4/xTWIkG1
IG83N/rNYkoRNgGxnhPFZy5WA+8qR85RAWK8OKaatvuc8KsUVqTI5I+B5mH20McWpehLJD/mgmsA
K04ssUZLS7eqCh681oQt+s4yKtRbArUiGWybEsqFijkDXYEBs2rWE5WOcTbez2NYu1PVJJOwzB7k
UTiL37abi77h5o6rNJc6MUC9rK34pzpw7RvVDOsWAXrA/S8DPO1yrlwRxdgV+E+ofwmOApmTyjV9
FmuaOfItdDRS/hhxLOPPZFz106MSjREz57Ueqp17arCnRBY1tldMPd0tbWx3I68yVcXjUw4y8b4E
jviKQv8uZZ5fK5N+n0tPanh0Y08Ik/Co58Tanu9ansLCVPc6CNucnGPiit5t9l8XBhoN89pzS8WN
+fJwEhtvIH506zxE7RNaYuATiLj1gmJbI6c02Y1LrWh6VX3eUY1RwkOkCcc4uJtZbf91Tg7SB5lI
8tEDDu4KTtbm6uXAx4ThJJDrUEHS6SMdYnxZbx1pYES+0x/S0a9F6jEemH9J6qgrH5DqTaaw77gX
nNSrH2PNfvY2WHGFCYLSGPOI6T2oO4EjFNEOH5AfEt1WSSsaGZ407aTZNooV3KFSuRDaeG+FACgA
ek57GokeJ4scAEGeXOgidzEe4oRk41LELdftwIQ7bUdAx58KinBW0z6FmRozs+5WmN8CfgKcnLC7
+jB/cVgiVn1X2pIgMbnjdHBu39a3bz+5Ny0XJDVlm23u/WINpglpYRIxEEFSJ5c9pJ1HCFNl+NqS
MpNPu0d4pkOf9FejKWTNXekhrbGKftFuYXX9ZeBAcCD38fer4YhW7p/wel87NAbqrVbn698Sy7ma
mlpfDakagihdg5fwXey7BKV2JCg0Jn8STcz3znZHViO7TxH6Aj1f1HzUWTRjxhQl8IlKvqS1ejjm
HMLgaCS9F16TfXgJR38qRumUCZ1uBjgUtIpA80ecF9TQnUzZewNzoUnhfeqeQDk87agZBajnGh9J
3Dc0GEwhTUJ/7F0ZvhUcHlEVKn0exlVHsFFE1B/G7NDp5ZHOUMDnFEBCCOcjC54t1Xzwu5jf/VRM
YeUgFO0H4LoMNnjm7YijPnRTCiaaCqcyFdp0oQyd7222uQI5FQEikeU7jrDKy+eFJUVU7XHhLPLk
oeQD7mJc2EiZrRgKd2ux3HF5HywOhXs02JIV9xBktADP/iRGmVBmpCtRRkQSJgZ5nFk9j5eAPa/h
EiaC7zFGmnY2eJ84rs6nuw5F3DJmGpofuf3QqSpCVlEgEt5LM7V24armlWaeiOPIEXD2voyl0xKW
9ajyhGlBfdVW4mkhWOqjVW1r5m/8h4jrQy0t8aP4TVj/+ESmnrH6dZDRh0Znb3BaYkVIydNia9Yb
0f49p1v4E3grpel8qiff6ix5u+B8RQrXfsdYngHKLZM1kVp1IV8d/DkyaRhqz7pejQTPZXKMoVKO
jHsG2bqv2D53sJZaOhlS6jmZLWabIovcqvDEROCwTAn7y8h6kmIc/CWwHbd1fh6m6ZhDSfUHv0I9
oyzGJIKTaAqu4kRcAyxRRAbKar7YdSHjEYgRARAoTQ/44TGMFX5JSprTKrpWnW+WJwRMS9RnamTO
Vo6UiO2NslLxXseQddx+J3sU+PmWgBUp1g3eaEVJTa3sAMDdiHbwW60CC2dZEfeCzrJziu2sV4FO
UrtSW3qHIL3gLp8EgC2hdcWetU2n+JfbPFsHRQ5Ga78tr/RZInPyKNDRNTIGVYJ05/R7AWWeg9yH
4zyRaNcywGcVlgBMuBWHIeFkAhO1lUSoV50i/HoNlmJ1TFsVqYSAN0GtissCj6YIezb9v4McCah7
I2VpCjPWHx1ixXZLe+oxZbZCVAxN1u23J10HRakkUQg8UWCA0faxjBc+c/vyk3ICUs2tvEHMvLRn
mJOVQ6fPT7xZPU0yTUnPvu0+ZRb0vx80sZlc9yW3HxtJKgF12iIXniCQAPkb2aodUAQkirqU9/iu
5mQJrvWkErnHeEQBJpdRDILJ+tmfHR2TydFxQfKlCoLAxL63yhzayPMQT/g9hJjKvtzyeZiuE6Go
NTd0nuFRnMXll6gAm7e58N0Cab3xKhYGfpJX4MoQA3MEOHkhnl/ZYXR65ocj9iL0VVsNqZYDS19p
y4AKG1ZSw0qyAMmJy8GQMoSS9A+3NLa9qDqbS/1v3OsClWGI1S5mhJ+ffiRobf5KwO5ojQj0c9LG
LWFUlIstlb1XTB/zrsst8Wj8ZOh6F4eCC9XwD21bxGYElHzDiZytZeYUbHAo9ZFusxFFKnOM4HQm
mRZWQDPvss5pnKd4kYuHuEbhF8Znx6+lnNe196KQ/Dezc9okFwYGzaKwH43nBY/3XkPvwpmbMiNI
rDxMqh8FoABfG8H9QkIqVBUfzde9PBEKPUScpOXmya7Z0wAvi4cLaShXP6eEV3ZQnLGiacT34Oc4
nCV8yHi59MyL1f/6Kx0M0q4o1TSctWW1y4zh+uJMDx4apCwzQQgoC4YBxjA5f02NBt0bd2VVV7wk
ZUqZFmFC1eXgzf1joGJhQ2TwPrxU/8EdF8s38/KWqnxUTBHkFW+1Tb9MD8UllEyS6bC9vSjkJJJc
X/B3mpqld1mFLQahyDhXCovrVw582HwcATLiJk0FiQ7/SUGDcd2BAjo8ccZUueL/siMR0k7jqTJr
VHwG1bU2v4XEaYtrgCUF+27NZBtPuUp8228LHscUYjOTev6cg/pVLWf5JyML64t1TCBoC2PF1w0X
cFXbIsF6w55Ay1u3buccfoHVUmKod6FLFZPQKi8sXdd5hZqcxDxrB6/E94yxyN7amR+ZVKm/q6kw
PQ7Rgil8Y7kEaiik6e54DJkIxWiv4cJHR2yETfMBSHF3/VE8uc3V6OTZ+4Yc6jTA44BvUXBLwUPu
8ghiZzhdaWhLEQPttTHziEig7n2gsVrvnuddIHIGWpfp8YENB/JKKuuIjD6nRIA2LYDXTudhnTN3
xG0+mJ+/nJS2eYczpR2aD3AnDm+a0tOf8do+Uw1T6wiNIVy66HlTitAOvV9zQHVijJpx75Sb3NW/
geXW9FH0n6ET9LCVkD5OqP3HYbjXM/8Gyr8c4/IRj1ObXWvnFuU61CoxdSabaXmgSHjWRhs4Qb6l
y1Q1X0L/PJnoGV+Lqvpl4ewnHP2lt21QWjkZImneKjPwt2CsNBG2NAA+KKMvsPq/jOSAZknj1KJ4
A/fDMHpUmwu6gxvILNru0yl56povmP7O//6Q4qPLdjtV4fHTqAB6j0e1NTRIc34UM3YBgTrLOUKL
qNGl6DGBlB8k0STeUR92NsHmEhyy64vDmT6lG4EoBf/dxM092h23CG+BsEmbujcClXmsmbJX0JMI
rSDRGcXMlZJpaGRpRoj174JP24Cw0/9e61/aCEv4THTAWkh37no33pO/h5zY1O8d/tKu1kpZGyP8
+S4PZLOs+nPfWGayr6bWxzp9FP+xpdOcAVOSZTLh3yCDgv/GhVgJ8scAtmfLvvG/qSy3K1Z1fuuO
nh0SADKxVq+Mrc1inRZsNFuE/VoGGopsHkZ9sS80Mv4R9X60yN0ZsDZaP8xH4B6kuNCf0Vq5TsXg
dFXNlviLIEx5TYl7LYFx/Y1URRu+4Ou8obzVY44fWQ9zo63QzRlvr/gg0yjkKs/tNG76hKCJvGb+
3qAnbcqvU0uoDMfZC76uNRZ8haH/VN+X7gBpTot3TLAG6J1+ikWeej1EWERLX1nST3QyxOHAGrPP
A5V/zXsgfvV4Gwj3EoU7upW7Uiv2Jli3+19FEdP4R/Jan2rJFp4zgrAL4JA8lfJ+lUIexwJkML97
CqZjdUX7CO1NO8MToQVFFqADKHdPXvAHsrjnNhL9rFjI2XZuYL2Wj7zFoJKQcIBVLM+n3o1xSU59
60m8N3hEpjCaHjF3VywJm/Ir/uydpcX/9cxkripj8ecsWno5dqpBYN2McNfdnnZj9ciN4+e31TfH
GOVwTeD1Rr42+1O1GaWaO2nCa7CisV6riERiGanbH54uty8NR0TNkE2ZO5OyL50MFfKfO38w6D3F
2+lb5a2avGE6OF8G/sGpPlchgY3Pu111YG0b8iGPrniagPPseCktO/CVN3I9207AwUp2Y2Du+Oev
O6lxlCaAiSk3Ol1o6jdVZnybj98/6DACmOz7MWC82yX5p2ERo1dBpl0JEjaAvAKZISle6ESUvQGE
ZqnMXI6WOdN4Kp7+/t4ADJnc91WxkA+s52Qmp1LOyphH0gn8Qg7Zb6z8ilh2YJnEvVkLd7Uq1A7Z
5XVj88Wlx649EXDcr3MB8l6DDf5lPbBF4gbAzqxqrh2SWRmT0byWOyGRWr1/3z9zx2y78IG+uv7o
b0DYPi12h+QuQFOXz3NLBOYCjhEcnmoDywT6Tcf1yDYBPy6sC75n7zW+1jQsExkAAglcUtiuBqLg
C79I2N7z6OpssFkPgFuXgragTxp/EPRjTBhv+xqM9yVfdVrdk379y2wKo91LkQyoEuOHCk1gF87A
uJkb3KJ8HM6AXSVh3fE/y5k0iurScombbHeK0m0SuHXuNFUuOrUwLReiU2m3O2osgPJGQeNI2QtS
my/+DlocLmDzdZsgDtjrFuK+LDo85jco74tgR1YygVhvsHXxO4vuDzWYaKu9WTOOGXF4EtBM03rP
bsBb/GY/+ukCncmV8noVW3j8QfOGXFnLn1SKhvP2a2CJ6T8w6yUgKBRinVXNhFBkZ5Qt5bfA+R6a
zCanYyWQoGGrHXGAGgdb5YPsD7vyd/e+F6VTB/E1M7BLulLH4uBVvnNPSM4aIWVF8yKY+0TLg4te
PDX8qB7/LfjbHqxuaAYWwIA/Qi38nJADLg8CewBgy9LN/yr4d+7/jb7ks8OtHfo8bbIuLJj5H34y
Ad+DGNjuvDqdJLjfOCQ+XdmL+m09xn/RDyurYIeDwBURaWaYo11Z3J7smIoYufyuqpZXx/3mO7re
y1AN9zpynt6hpTSTq2Jmsb53KNBCrF+G/u5JvnzmwIhlOU1ug++S5GOZ4JL7prVXMZccnQ9tl+uz
r2P4Oxl4B+rr6HpCNB4sDTQd6f82fdZ5NfjRN++/7XzqQZiX5FrV5FxqzGyzeunKkw+6l243a8YU
0caAJ33d9whfsA2RhgnFvmWkMQGc1QZyMnxmjivZE236GR6mYFAT/cHHCi17q1rPjHjRv/w6DNiH
y5GH3L3tcvWf5cXLXJqBYbKB+hdC6tBWGtdffpZ0sccqEiVXfsw0eHRcKuogVN/3i2Ky32PRnsYo
UHNhrQ6DyADyLWCmwwtZn5Dy5/MohfEIEgifA4+oGvAaZKeKvpWd8cpkdG/KNl30XQrjJRFPJnI/
8+sITVp1YNdGBFml3vrKfsI/X8JJb+WN1VIf8BpT0giXpPy5yDG7+pB0nh4bwWh9Aoe5AuALIHVR
MvJOEeGPKgnuJSUD6bBHXxybg7nBZgNHXl5NdmdwKY1qW2PClOTrozUyTtaT5Qvc32hAwEzd9fIT
WNWGFHNhUDbsBP/Wk39J33166wsrpkndRPNcUVz01NRwdhR5iW+k/JZuuMtXfbjNU5dJFpcoupAB
HNRN/2ybT+e6thxZvegySUcQ6aGoNw8yVBk/juxxKCvEjrWXWXWEbITKwVsLvcQ//aWPs0VYGTkw
UiN0Gn6r0O/qjTtIRBnTCslMTX7PbP/fh+N+4nuk0Bv6N3S4R+R1s2+uGJYPYjtep4wXLVeFYkgN
nnZG4qBVXRC5KEngVk6dm6MwZdVZ+iI7h1Ya13klzRwyXEtVffDToMte/L0RJzL8MZ2xVLgxB7Wa
OrWSqfESaB7cNpLyF0z+/VA6H3g7r9L5Fk1l1RFEumDOyNNFpiH0nI0t7qGpHFPEYhsZwS0g4QWQ
emTukQpVE/sd8uR7AUpM38pDSlkO/qZkIJl4Kn4MvRjX2mNgWEqFiZ8YVZnCpFEMrzYd+EHidQr3
GF3LS9O5Eiwge/U0T3TgyEoiSTD4h/XXu7iUKu0HTK4NsXxdjQQArng7Y7e0EAmQJz91Ly754vuI
TnzLIh+TJRgJTu/7DfHXXXq146n/HlxpY9Wn9zmY4/zgXYiLsH6jvbwYDWOEJ+9MSo7x9T6NLO01
kT9vg+x/Y89oGNZ+DyDBWH6anpeDyWqCXyLgVV/hIpoWudO6KVP1eEZFfXzmMXGi/FzgSSVLntQo
CsvfzolPZByCoPKXbF00guTEzNiHU/l/2YqU/zGXMyDTOvbgeEHlW/4czFY61fzau9XshK0ifzvc
8vbWz0qxwk4e6zarBJI6RYWoSJh0Ny06wVCweM49tOp+lQEuZIKM89SurtmWCi4lEXyIWUqCeIdq
WJCcr0YBdxX2jUu6Cg0eqCaYUDslDN3XP+zJC0Zr5XH+cT06XpD4Il6g/ikPyL0RmmqbM5HZEJ+T
7eAuDDgxZ3ynkXkIlWUBmuuEW/NPRvtnQIaWI/9kKtkzJG9CjL3Rzc818Vzkm1cnSA8Lz7SX6ufD
/J/o+iTHbJRE3j5ZMk/gmktP9zVlA+++6XtauXn3Q6sre+aDercEVMGrXHz0bVxZpeyXjmsPsZ8j
lLzN+YxvBAv5Qw2AAumNjJJPmYCxkmlpANxbuv00y4YdalbtdI17xUnhef1oNrn7IvWA2cz9Pozz
gPJrLPHv9ovVgVs1AQBZ23gPEOz+H95TLVHEFU32Jytg8//uGuFGMiGtpl0U1spiNqmSpPnymyMV
6G/zVTXJyoIKAzx38ckpttK0PbGMtWtPy42+/77nADOAlWCqsO+h8yNmibQmWBMzEoNkx8Z6qQqH
OBWLmrOdopdQ1KaS2XxwU7M4Y6+k4QoFZSpqU+O6P2aACX/HHjHoCzWcnl1NySTJpsJXWgJxYyT4
vcZnGB5BqjUerGPAlve/G2AXbbLgHWezNSGqp4FSTNwRBhE5GCYKLP9vgWdwq+RyJEf7xOuH6ATo
PY/jmeJ3vjPnDRudFeFoBis1W89JHuGjeLSSCAw39OngMeC05NV1t65r8/1d16m6Ed+CmJsp6ZS7
FqVlr2p4PFVBl46HWFXBCDB+LTTN6CyLBn5JWR4vfz+auUpr69/0coyTJOLjQQ0oiEmbQDmFAk0g
kH1Ot/KCMjKMS33hRyWl3gR7ajDYF/RXz9dqP3CQD4ACxRChcSMXa0fTN0asWk1RQL3XvneiiqC1
FXcDdmGmL7ZB9QpZh99bJG9LrD137IaduCKZ5bmVNybxRvjJCddZ6C4Dy8S+sUvsm838e6kRq4lL
Z8AbWWX18gSbO5MZnUiVK6lLC3C2abfdUvEk2jAuMnLnVd1Ns2C2JuYXQ2cpN2pmKrR/JAhZzlmw
0qWew6KaAqs/nnpOKZlJoX738tq0a7CIIeQfUBCc+pxZLzWM2FSn7pzMblSnZpwSZ1AfSZyypuQF
fN/rL8bLNA7YBrDqrMFPnPHDrYo12mcZOW+inBKTpUoL9XSLZI6fEi1j5ZTZCUpibb60NKWRrCOg
3cDWEJM0NNIPMAwo/ODfkE43QorpnIMBTa7xgFKfdKV96cZWDKBW7rbk3p9lYKGYXKbIgzHf2vyR
wdntNZ7Vdu5TjTKGxM3ENa85yT5xYr5Gjwig54NPytp+MY+iMV1vGJ4jjy5Eh9ZCrZ+zHR1Gburl
jlnv07Nju2sKS3zIWXx0PD7cIOnx5AwMCTqQFW18r65/715HwOcTO7G0AfSPE841WxFySi3VqXp3
2MMExGzRN226OLF9xvjT10A257wK1wUcB+WbvVAANaugcqlXOFtoEyq1LjKT/NL7BzibfrqYAnss
Vus5B9LfL4w/jLUEbMd8yRDWv39ltQbmZAh3mFh6pg1pzYnyHxKOClbrKyAZgwNm57QBGHoUo5RB
M9Pvlwcii9aJdhj8hq5qUoH7OR3vDRLISJ79kXXZDtTaI9sJZdWvV+KSrUXDewXQveeqGR8fToGy
UR9w4H2A/5ngg18a9Y4JejXOwL3etzAhy2gB2iQaH26OAkP4uagz+NIyroFjY95EDBbtlXFoQp4N
hWll6XEEFjD82qUpFeaYHSxOOyWh8dl5OyjHTvwtb1Unq0DCauMJetI0d2fIgz5KACTXd6RPbQql
C9DOxm38d0su4OimhSCZAwwmM1TuY45U0pb+/PxlgJU4Q+z5VnqVokD0x6wscq/FZQE02HLwh6eS
SjS+01YtHQxBAC6xWg4aBWeeQmP3q7PKRR/PzYNt+Jjz/Lux/yiaL9yTJGqezp/u4ueLNgSZw081
Q37YXdMIat0vZUdT/avV1m2zts5C+JmZFUcJvnkTcLRNS8I4TY4jZmtmjijBj5pZzH7Gi00qbkLP
pdpLEeA5WfEZN+6wn2dJzFJzSSHyEW13TyqkRvVzAJFDJ6rwfnHHK+3sKYpZHQMz4+TrqjIfte+R
akfqD/z2G+ZEt/GYGXSKEtD7jBiDAuSUOywO43ptJOi4Cw2JusyBPozuxzdHDcyRRStS6C/ddLxk
VqalnlTphBRTiNMFA0WoBdXYfuadRJd3S2oc8ksf9p/XkrroiM7BBiD2S7XLv6ctmEPLH9vrx1jZ
iDw3pxxKY8NMDCvbl0TfHM8Owk6PRFkaFtfzQbCodx5bg6LupwPXnl9yOkMz7Z03UdYY8LjPeDl4
vG6iSCEdyVjM1VC6z4u4rQYAun6iLQJcLetcvQHly2d2ZQcogwHjhangDVHz5Q4+h3G/wnWF0+UN
wklSsfGMpC+6r7YYFyMseXQQZgGY3psnl6/xcwScv3qs3oZpjRku2u56FJGx1bd0GJctW9NfxQtl
mmgny5lB/qMJW/Ivksuz+sVgIFtMM8KKv8bWr1xCkJTMtXSKyFuExPUxYdSwFYleAeiR9Xu5VqjU
r2MYTomR4KjbtIOI6j42BXhHIP2j+1pvTLkz2xK2mJ6r9D59M4S8UFzSPs0hjYkdRZagzRZAZtHo
m2I4R9PNqFpGvofODW2W1iU1Yrl9AJXOUa0tKgLA+e72YtTQx0VfYFfNuyFHNNl5k2wzNgKHLOUX
9idrRli5uPeABy9osiAUuXiyRO6U8/jNh/DLWFBlthtDKfkbh4nKAQmFFHAVZmarKsRFzstdf4Og
B+jUnrlJOPoXiDPYj5L2l3K4NHPYbLjRV2kxJlns/So/MmhLlcWIHG6WO0QMr2CzJGjFq+WcJQg3
hozedzThPKxi9EQfQUNnTNxlBHVXGrmb16HGTgl2cXfSlRPzQLkRvn87ikRKrAIdHq8W13QHhRnA
L/smEQzt6fBhodL0l4/T/c2VBQaUlvOe9JL60FRNvPCBVpkDUvp6u3qsgu3raS17klYGYR11ZNUp
Sz4VMHdeoOw64DORMLUhgrMvJVSYnFs5lOBwiGkmF4QeyN5ZWkaTMLckcyCYuWngXGgecT27LLi1
zW+4ruwhRUCNjDdeoDUX2+OTUHT7DqOSlXkyvK3109f3VqYsK1gSx4SNdRXIbmnjD3TUHtEwPiHj
9W9+pv1UcmQoXgK4UYteTnGCLsL9G0k9FWAyxGaWDMmx5vMUCQ1bwccT1m6GI9VvNjjK2bHFIr+K
J6Ey2lWLvsr9sczRafxa6ykWJyOgyUnRsd1+xYm28s4ksdW50KdDHjUDzqMmMG5K9/7E5h/I4zw7
Cd6A29Z1NJgHsUyYWL5DfFenkaRO5jgpTeBKuWbGXFEirPd9bcQYh4w8lm08dNhr2/HpHaRsKlf4
5TkaOgadveLRcJXteuhMVzfypnLXhRFhifN3iplkNnY89vET5hWbjrTPBYSRJOh5FeDcPdYFW1+j
OsrzXfqX74j6bAUB43VWBx9f0eo+euarfriZ9B4xDo4Xx+EX+m0eTYuZ9TrT4Njog6uDnv74dz2v
I4jmSQeMNU5xiJ6xW58aZ0hG2B1IgW5jSeft7YWQdVew3dJ5oFDxRJDja6XTl0ANRWq9PZ2qEVAY
Ir4uJsC6iyeeGfDEO/edh7eRRlsJqLnyQo8P7JH/8sSyh8bPFAaji1dKlmO91RrG6d1+iraL7APx
jlnCUFe+dqprqSUGdWLfqFMYZMKasnPY3jcOwT1khP4yDsT1OxBt59runif74v+JGMY2Rm9R3N8p
6NS8cePvkgFDTA+NLnjqKCgUlgpsTHTWWxg38ab6FEDPf2NLg5mNnhGFR4lDbtRMKImBZ4hIgxX8
+H7ExKssC0EiONs79JHDuZ0jnoQCW5fFgalFBFJiAgdBnoL8NC7WfNhezl62imf8QkYW1xI4iujq
aG83AT82PQz5oxH+5+xrDjNKdpvPS1mUKtO5PKRWmBvQRgXZjNhXgIUPlI96apDfy1u/gtWfqOGS
xNRLCTb/Sl4HgwxE2/xgTvaDHjBjKolXdaSHJRrqAkuTZRk1xXHc9UU/zTs4DheBkElQ2j3/PjG6
dZfrUpRpJFyj639HlTTFqBjPdKA6iPVxqCu9qxBbIbC2EU4KyJE5lz3wGnvqpKnyumehGk1WgE88
nFdNsHEF6hXb10tCSlgLpcyYCYBXlPyYAiQax2XIWE+2POYVie/2UASvY+n3qmhZQh8eBdUb0oYg
CUVMWZEZWT3vqu/vzQFP+nlQeY1VOiu5lTi9gZeGKJZ0oFnpwOXGVNFrwmyhNX+4B82rcd5Pyoew
zBUfYpU2WzYQWT9aISj3K6Etsc7VcRCzIqiKsAKj0TDVUnLVfgdHWTlA1Gb5xN87Y6/LZ9btinQl
Ou16az6jk0izrm9mHaCoksH2YlN7AjShpLrVV0FmQT+OIAUXIziBBVtjktDjfijK9x4SlyiZpPUP
7MrAEgK9ktQ3f5byQ3IwJSglWHTFgvwZxYMwRy3sGJfWTPdVX3Nj4cTh7wbc7D6zYOb1rlyashTZ
btoXTZCUog4kSrLIZG+7AkIm5f3s+e6O+vIQ/qYQyu3UAqESjyn7w/vGv7AZRgmzuo1FryrMaj3O
OgEr+/F0O8DS0gEvumBDyIMRwbiyMHKJALDKjduR/BYB67qxyuFVJ6ZpheIITqz30dOwBgr3vShb
LG2d8CSSqQwCJnM2mjXVL1u48fTD0nvj3Lw7DebNkncZmL+pVtDl8lOu4gN0co8YGe5qsBaDhccL
hglOAxUF/ePgEGYn1dsfqRtAv65A/QL6mDCxvfpLA5WHTOlcaoq547TkL7FBnXIZeJUzUF/yOu1R
IuGGoa02HOe71uRFkwadrm8/tB7h3/rVhEKhxNTtWAlPd6cXp2w8ZZtbblza4xIhd+13sTUlBBFH
zURXo1SAzpLb23nq1RIBxDjM+MZ1Hx3Qr9MiU4A14O1XON91GLm5AUhjhJ51qorU+Ed/hGOr1Bh+
rs/OPzl27PSuXBdph15cMuG7ZYo6j91tK6ShTaEC1YemuAA7WFWExg7ws4GUlQX2QiWF6pdtuUQy
k/Olax74jeQSysoUkyeaTPgkO15e2idg3BuG8jl0sC2Cx1pn7BpEdymjJqktZbuLw2tlHnF/1er+
BQuaU19VV46RVyEpVJA+QFpUzczUJhphJjWGqNjoe8eH0CwnjeEzZHD/h83xZqWjVLCIK7teoCfO
LuvMJYaRiCv0gX44GNFpfgVNEpiqiPafkGnApAkMQJOUBfR1V0a7bSfbDmCC8rZ1TuxU/cr46wD3
zDnOVob+dXtR52IABfM5pI4FQ48cWiddkmUb/qgBOUsobwmEIaa9EcQ7PmRI4CPGbgrWIn9TjElc
BO1cwngj8pmVpiS0i/XT0Ql4/ALqiDy71zg3ePDkF5Ekp0gE4qvbE1ngjj3qWQxXjZFKRowLS9rM
V+p3evx5n1rMtAd12D8baj4rHTN9Q1Yf6uCTtyTmW+sDznDR57C5HhNw8cN4BAJZxAh0M33QU9Vo
XS9+94ZEbwWeo4RWRvREylEdABqgTt0cn0AvosXWDG4qdpl3HILmcT9mRlSUA//EcjDl6mcg59qQ
WMQSoeHfMIXBA5DTpTHDG6Hn7XJQ4csfppZRZZYACUJnxl3kv5x3vDA3JA+FKIFER10lfQwJq80p
ZmUrXQ27quIkcea9SOW0sk6Lg+TPGJwk0ugNmJg6W21E/nfXrdxApI5OeVnMyUdwOVIHMWH549rk
MWPsA3ewMu9v3WODsatd75Z5bng+l5ZJYucdwCwtnd2AmpjrRjvy6T4t2hktyHB2lAHCA+LGISxO
/zAswgVtNrrlFP2EutmfnCMFu0L6DYXNTa1t+noN97pelsADBkVDhDKlJjUxBevDdPG1I/CN1KCg
cZ1Kf3AzO33lx+RN9dzwmGz/TbGGBuKIioNVztUYAQ+jQz8Kt2Hc1rK6cGrE8OFwibIgeuSY1pR2
qQ7TByxbeuDyLK69C/F5KABSSoODwTVf1eQsb6eRp5lIfltAm4YgcNxy0HsnOVnE+HFF+7BfHZFs
QTGRs7nRD6hP7h1CZyOtsjfLuYXAXNqzJChxiuzbnfcuJ4rT30bgy9orqfeBDd6FSPi9PA796ul1
hyFYxsCIQ4mL9BJ+I7m3jasOX+7ezI2pexhTbU/KBcyb6MKqg5qzO3VjC3m7eIqrO2dYcCRGgGcs
NcvBJgVVha+k3NBTT22y24manFZ6vCL9qjBpgPhVpFPPRh4776wTY8lofercjrcCpiDpVYKawFLd
FFia9LyNFy6o+aC/kdF3R8LiCaMYcYc4pRQRTYpmzK5zMTET5XCZ+d+EgOui8ogovUDsa4OZAZzP
Z2yJp3GZ2VHy8P3t7p0K3mvOOkzyuLTUzVGDD+hHtVNjhv8M3OM9mjQ5VBfWVD8gPttkUx9RzTqK
yi3NRcnj8ZPggH8omQM5EwNvHxYiRypNahGlhdaFrLptGXcjiK12cG4YRN/+uXWA310ssNdsU8ye
7k0i1yZ0e3yXOaRy58qlIaxn46CgG5TzGA4CNMpkfjOsoJwewMtVr0ULfPay+o7vWvSNGNmaIA6s
cfAiho6wpbdDZ08eHOBoeiI8Frv1/8X5xLFZHmEnhN5Hnhv5fKRQFIaq8lBkG6MMLREhkZbAM3x7
nrsNlYhhstiCmkVQW6JkQJlmWj4uviQqlyWGj+DLIqeVs+DII2qrEJ7dWctVFnMs/K2C/naAe8+y
2FfL87tSLUEMpE8Qe0CKiEgesPzA9NOBtMr5y/Ht7woCAec37qg/B/YR9ZPfX4vO9T5C2rIxySpY
cOfJ3W9NSrUc2BGUtpOr5/6jaWmZNcZm+IPl7h0nzmzjYUynEDCZr5ORCuBzgWX+YjC7iF+0w7Vz
FvycZzNDauA5h0vg1JehdeKCqvM+2qh5KndcLWrfe0b/fNHtw+jPHxf0LkapsgjGYmcIiFyB7SLL
2NlqxElvORsbdYCY9qr7Zvco+EPc59AdA925DFXRE1Pl+/AmjUd0z8HR0SuKzIKOqLZoJt7biz+z
w1VqlWMJQCSeMyqpUrZAL/MDNaqV3xG0LOxlWK73zTU3G3uz/RyquT+aoRG5kHpSifHOCwd/OXV6
OC953Xct50RSjqy1sA+YWj7P5VHMVWvEmvA0bYgWob3NzGKMMH3enounvv7jlrYSPacrD85wnj6I
fKl9q8cEKLkADm+ufLpOTJ0lIbTZjZloJaRpJJHLJE1nWh1nh63hKjUCnPwNBpMLGrrZWrdyYllE
9DT4gl0sc1PoXrYHL7hOjRkyqEtUm5MU2xN/xuCLN+nHw0l+HGeluXI3I9WVhRmW2qTEu9DMgcYn
zT3ZtngEDT63zDT0Hx9F+5NBKtse+FUXUxSGas4yoKoI2SxUuozZ6O8w8CckmOI4Ft1gKFStb0eo
z5TWFhoKO13hOV++8iHWKlNW7i+SaVtEL5WTrptpqCk6wx5NmWrHXZr912/W76WjutrFjMB51/28
zvp1mLWuif4tadQjPXKFweIgOahh9qFeBccDnleIuz3zxhhAcY2T3jibJ0tI6TvJ3zlbYcNQipo8
kUxsqNByGA4QFnpvuAbh8PBs+b2PN/pT1ZG1KPmm+5E/J0pcoWh5KzIog+XA2wBsOgMDKfBAKJty
Yw/AYQ5DHuTSpFurKi3KXfNez4spl4UcOngC2rtBtW4A+qKMQ/JgBBVgKG4nViM7XQIHx+D8/Jv/
QY1LwL0kdnrILv4h3YoyoZA9/ch+y+WJhGOBTIFkjGWGrD1E2o6FoaO0PZqEXUtZQPcHIuj3ujKT
74DTikoCpEFZfNrWYbympEZwcsgGUbBdl58EB7GchhbrVf41Y0mmKRcCjC+c4RYyOllTulhUgGLa
W0z/XXmdOq5DzKZ3KeU5mljY6KVyourP8MJ4EdjZudNkm4bBvcYMSQYkD0krVjCZXvBbxv8ao9qK
6I9QI3zwV+wA2ykn96gsFjpY+10UdlTysNNtLccKxmJoWF+BqYYg8Fv0yDcmMSL8xtnG13/nzhsN
sKhOWkXPIPr6bBk29oZU5SqrECqRzfC0JB/X0ACoPVcofPUnsIHv7JhBekBMy1qGNRjk3ebrgL0F
shhAP1VNNpKsmTPQ72yuveya91Lp3s2NKve5avFsnB+cqf7cNbcOhKztbWaaDdau5vM0YThUdJBf
fexFn3S/F0mdIEMYaJqVaiLUemcP9zC3giguHD/vSovN8ZOm7SDZDwAzrjmzaYeX/sSL4HQDcLU4
8pSoSYp1H4GNn3G+YA/ZeOL8QkmzqttQu2ufLIQ2BmJhNCX6OEc/ZgCd0gxPTsFEzaeckADh3RGo
kxzfePEpP7YpY27+PaG8oRgxSBB2z5McZI0P2PfYp5yNHSKGJqIhWIHOrHgUiJVQwaJw9oFgWd6u
VjTOpO5FcUmTf5P0QL0xzw580J65hM4TyWbobZwLihe+Y7bks108y3QFdawL0W2srGbZtzWdpv/R
98DECvdajRJE0fhEYZenS97Wt4I+kk03FNmYOWx2BsSnKGMFC8+mpxLitHnHneyADvGMDcksVVue
IdhjqmG9vytJUZfWB4BBS6H19ZjRXxA+rNbGNFuxwFut3V5S0t7Ckqr1nA+5f4FpGZbX5caJ583e
nUj8VQooyGnu6oCqEnCEyYbYbuFXx18O2RoQBDzTSGzhMQhPfyaxMeUJQ/dKcxCEzmamdbXoJXss
tckUloWRTeHnjD9HjCiAWEeIXs3drh4XCS6JRqoMfs2dsbeTgmViE6Ifv1GwO2MC8gGuL6VqshBr
xHw1nCvYRjs3D+22ItL801vYObUaUrwz2Aag6ErFFh5a5DGtOYKM32KqGJWxkmpTtNnbEl1yC+BM
8XFY6rVUXDvPnl1WR0euUREKpNZIq+wOy9iM45GPEHcvk35a3n5Xmrlw4/vvM7S3p09xFhU16+r4
dv/CDIuBDl4zV+s5U9XyTGm4n2HZsaYdWSsMYDek+YVjHIcDaxHAsNoXonHCOxmmKE3IJdXS48oM
OHUh1p1IP8xblf/gCEbiLA66XgeXvVT3pkVNB3sD3KHOngl2XVOB1Xfp5MPbFbtnd0FC1SMQr0gm
lrTq77nc1KmgC4pbeZWwYfjJ3wdtAbKSzftktWyxOe3jMj/dD3NpGpbzZLRXvnYuy5HkooK7WRLk
L80X8kBrk6ICFjd6fzRzXj4rMEIgW6c1Ie3N4AaqL3q25TjXJHaYPBFhOZQ5sGO5fpGstfQtzgG2
JPEaRJMgVhGS8e+dLxlSOJWMbr+OYM0l3uMrz26E8YRyNmjCtJX3pZZntPt1tKlyq4qSW3akBfl7
neJWaEU6ScC+5PEyoKcGhA0Bnd1METm5vc/aoJbBvHAVISNcXa0PXGpj+//woQg6a463/nAozFgK
2Nx2O0u0sWbJCC+l5xikdLWVDcLe+GIWO37wKVQhtFMm050yYoloBwODipvDZOIbwDploH43JanH
L6BbwivLRnKtqoTHZsRCxEakuQq2vjwrOIUU1UdTiAaRzIZC+BTQvqZ5OjcbY1h3VIlynqL8nxzC
XhnIQYS4RgkHL0zv3+7kK2F4jJQKLv4pTtxaT1WzIx/k7s6OrdMUw5ko+LKS7YIQxuhrNJ2bzp0U
Rvptg6xk0F3FGyvI3lLflZzh5hBXcuWbJaGnYT5DzFEwDFKLYFVNJl5hw9sXpcMa/pS0oo2JwdK8
2XlkMFqVDm40mcLiS2W92sm17t9wf89oklvSsKwMMvnAn02thWH3IxRqAdAOg3QM9+WG8xwebW/r
PibN+ivX0ljF8kmrvaWzNiP7V9dayznlDqAxypNSep2VkUE+oZ28CGWmAT7PMGdcRK1kr/HrYDPh
ys/I8/fQHwa0RsPLYZt5e93DeCl8AhKYVrMNqSOYQBBygy8oqxl3bVwl5n9cjKRGhRlznapewLVR
ftAB6j0VDZAzw+hS7V8a+cGL4nRscolTkUFxRwJYCdITbc8YTyblPyGDdWOx14uAEbsUFp2ToMN+
ZXgrG21Kx5HvDzQf2OohKgohgDKSRJMrk1j8kG7cAi1rkG/RfFL9Emd1Pr7tw1ReuCeBrfb68975
RgqkPHl4DHPqB5BYhlFYU50OWO+ic/cgi16VB1qW3S2SZdxsx+vTY501CFElvTyNcWi3DJN/7QcC
RkS5BAgVlloYWQfQ+m2G0DiYPJ3QQCVMMciSKbS5IGxhmkb7JTLSM51UcC/0T7mYSdtyAaS1BWfH
tARj9UmFt8+++/9vjDHABwI/Oou9n6nxvI7cDk2R1fo9sLpg4uqO1LfwXrX4C0UuddVxjXgo8ZxW
To91KXosgo+H0+Kuf6nbyLsZeqHiaCxUMtZxmuPkzNwav2dnPTxtLhJnmkpwBOKY9jiEwC8yii0j
nmh3NZ0w/eEt//ziPiGFF8/YrtRSb1gMjCCWGGXi4xbOuSxwFNiwkLgj6+42PGGokNNuWnWtm1tm
dBPjnBhrnNPqaSgR25UkkC1PXdxvQhTQaLtVg6K65jRWqcssNNouYZk7MpJXK/g2VnwVxOKELalI
EbePTLupMmiKFgAVhzU1HA6+sPyhBxIWmtoNTH6/SqgBbr3q1dcLpWOa7/0SQU77PceT5QyWp9zU
tmiVcK/kW5ToIDme5O68VPOZTLeVI01prOIJi4yb8Ymxwkf2d0TZdVLW+wHH55kKCo5jgqcT0TFU
QLotlRhKBU7uSsVhDdUhnR+Z8Vne4XpD6w6vr6uENiEjfxc9jq/psufc1f+gdghP5IYOHUOP/ZOX
2M3lkwpAiK6ElavdMRTHH8tn/vTYDuv8bV5gk2K5bli58KHWlW+T3AZVnNlya7f09QocVx0w2nCj
7JbZC6fdi5gNQkahspgrSoWDZxlUi+bfPqZSkMEZiubdBuFlKcZAniBwCb90CmT4HtbTMWiqEsMF
g1Q20w7MWcga4cWraSSJI5rjRvhOJrUA7l+Bo5qJHTAle0Sspkut/EPZA4mkqIWKha9UTBKwLz7c
Q5zgq535An53Lcp03OTdNzs0VVq1MGdiDdrmkk388jAt6biN/OuyuISxOyBKe25njIAe4FqBKvUi
TzrBGS0Z6MMxamCSOEE54g7XEPvRVAYXhYCKSSl3EJB3RyfhRpXZNT2qMz32IaL2KJqdEx92AWUx
NxY6WAz2rRdoyJzEEhdYHPP3g6GH78XIwv1cjhFXYKU7d5ajpSw3rE5RLEarJ4Zc6sLJrWWbUuEr
HwDbWuAKEufe6UZ/JnUgSA4TaWShwX8eNvlWMqa1hO/C5KU4oY/1T+tLLgM7tDepa/Hd83FjRVqY
tOhd+5Leh09L6sRsLCenc7HcfxjHA8aRwCwU6C5UPOK35KdS4C98vQ5c/STW2rT+9skI+5ukPFet
TLcArhwfh9YhQIa+HfguC0gpn1+n5R3z9qaY//pwc1yNzzFwz4pXFUiCMbfBkWgcLN3LsLHoX1q7
1lNev4SBE1TEF4Hd6gS7nmrcQhfvcKOCglDV+88iW2vaQop0FF/gfFVhBYrIHwLcy69cW3xrhHN3
r3+xlTzt0XfyScZqTMy/Yqv2o1R1x9t2WtL9e4644H2ICpPgqjsXZvB0qM+CtiqcCBm7GRFtvHpR
wo2LwkvSlISm9jTUX3wXccgLLxfSZdf4pX9EFOqcP2yW5k3A2+8J2YVBLhfSVogqmU6qpn+tQ68X
HTOK/1FAupmS5hWrfdjk8/RiVsTWzZR3rDk/mM9L4BuROu8uYIxP1bU2XlxshrIA2UjagnKl8Dh1
L4aiCb3xoCXeWXLtO1Al2djaakfvaGFYbCmoVlDHx8hxG/F/JGUDZIRZ8KOW1XlWjrgp0fvJTigd
4N6FCiHP4nDqUhIm4jMxkvwqvp3zj/rAjWfqpgqUWq1ociUQVrQXfbidk3flT5wzRmr0E7J0b+gg
7LDffAeLQI8UdJXVxXgo7/cOYlnTfuEhaueY4/je5Rm1pzU23WjmY+/wf2TU0+7X80ODfiCcwacN
LPkFrCZ4Z7JuDdyAwkZpD/cJstFN7ikKofHMUhfKEoawqnPCUZnZ8+uHzka3JWzbMf5py/Hwb5GB
KiuQtlf0tnSLT+Yc7gqqBg/LxN1kM1rg2q7UQIV4sh1gBeBb+lU4A/pzvvWCPJVJf3boF9p9KeDU
d2Tmrp6xoGXWC5vFadISu2YfKoH5g9V/G0+yaTJwTughLOCTQ5+P1zopNTDRffLzYaafcpdUXkt1
s0Z1VkvfwnKO/IMj+1Tsc0QHEVXa+Kk/3vfjOpxCaVORHqiQme4DthsGCP41H0S5a5msM4e4cUMx
h8p957zUsZ14C2jh8Pk7naPhSbYT3bOgdT9peDuUHYQI5mLnKAXFTmoYikF1HIhi/HxgqLtm2nIf
Zb53xzo4+YV+OEaQXFnewqn+OSztGojfhCkZr63ldXYd9kT5AmN1GpCjqDeFhpjnXObt+xkunWGV
usyXyH7SfdOtVUxHls1OBT372hPVM4zPhlPQuUNCm6NAMeGIVrvSZh5Eh67+P/RD1WA/8S+sLTYf
F009T9VMxM9H9zZFJEeL84vFaCRivYvje9ayv/r6BQFek7xr0Mj5yD1oKWqitxN9OyNqktqsJMID
dPpHskQLAXfCPEKngwj66fAV91oPyvEHXQj3dZOx2xxtHUVNI2amz7vU/6ja1ZV5d5V/+PZqhp5s
uLWf5F2uyNtw+8z5boEMsc7Ikc80LRvI7nfedzLI746Ox/tQSu4PEl+Z2NVa/8ZWsvGScUZYC9E+
8MFLbbShA0d4qB3B4GGE7LfgtG2I5BlbBRHmUH/tKgyqaJAraZ46N6CIofL8ljAWQ8sP3dLObq65
eRw2y+uPx2AVQcXCQYmquzJuh4bVnTXl3hHmx1+5ESxjd+dQ84B2dH87fJVibyebhw9N7jOEBAsI
q81FYI+PQ2/RILlevEyVhPg8lhglhUFS1+tJ/uzC+HM9ON/xd/IGzoquFRFvmVmmdA24EBj2Ao1k
V+hdQQYyQ2CfttUcn8ywXdH7AD8+KicnRbjZgiJX5hwxE795+0/vTMTGVHbO1OMo3B9rauJ0aiH7
unZGOkv9EY11BPmxj9WSu2S1Al1KFJhuYBBGvKpBmYytzRx8Dfm9C1VIbNGZE+faFnF/0iszfnY5
pkXK2tdA0I3biG3mrp5fusai8q2o+mTloCJqoyhck1Z2KBhFluDG1sgX0OQ2DENSmi4GEjHVkY2S
PLTo/1OjrzRBfthUkAS4nhTgvuPIWDhj7PI2IvRIP2Bnw2viY6UGxt6erzdCl5MNR/ADwXN2edOb
wefJMJoQYiEVO0KUyAcChL/CDk+DwuNj84JuP9ABix+wuiC0IRPpEu0D/Tfk/0L96wEt5rMIgdNi
CCHYZVVoj/UdE21paxlTaEkQCM/UeZYQRxTgZJGx85f9Uhl7eE6USh1wX5ujVNhBC9hrenv++HG3
nSzTn7jSvTy4KUUyYxaFLaDhnLEOtohHEScawKQg/LJwSl2+MYTp1Zh7IYJ1cJ64DtsurDlpBp00
MMwk0VM2HH6oy+pw7bZn9nozc4onqHdGrgBOpwipLsV/WzRXusb8sNelnjyViSHYna9pl0w71Esh
VEdYTdkl4DnPFdHtGawxfeIhu4mjVz5kInoNr5waZqtD77LvUSSZGHhPKLcvh+4dabU5Tc9xQMM1
cXZfV07Gn2D4x5F3O+vW65cuPmFq1vMv9Uiqp6DLO5imMNtQoSvdsKxkx3FM7ERMInXj4I1+CG2K
6HCKyi1Cj1lvqaVZN8pEVoDitkSDCgLWSEfz8d2jV06lSIFmzZjsiulcnzRd5oCgwzXJrb2+DIAO
hFZ/QNi+35H2ydTghZF7lu+3tluzsvBbda8BnulYLq3czADOx+rxITtaGN6td4Rp/yOW4apo6IBm
RaDCbRw/J3Cnr9YiWDB1nMli/etTV8WMBShCVTc1lu4IKXJnPLVLCD58v5d2USchc1X/rsjKSeVf
Gq4kBYLttPgyXhxjqJcuNgoAn9Yxe/S/lMhwYSClb9QYk9k7dk85KDzZUG3omffNZGzG3HT70qkM
euxv9QfcXB3s9HtLE85s1oj81OgKdzEcn7udt++F1oVBATb/tBz3bVXyf6RIpiwxbTYNPuPlBKil
m3DHYQqlVunEOpal2aN1ikkQUtxh2Cc9Ex0tUjrax3N2ZkKpRMK2lFB34MQV2jM2KQlGRTNKCGyA
bwF4sWHM2w07u3K6NsbPD79UQ/5AXmvCm9FwGCkuWWB5oTMhxIKvGsBDshfDRCX/rRtZRbgzoysX
q/6OCWahoqBqr8lBXMFiF0TwWrd8KESklIPw4KBPV9cvL27kCXPgtULhWwEnXUo3svCaCNrgjEIS
2JZwpbuvR2g1Y4jQTP8TeFklZza+9Cu7CZhqz2pFAjx+/enbT9j4A+7aV4zkK8dUZeQ1VBKYxK2c
WKlfYu83pLRIRkQKTYMc1Jcvd4Xf+imq4RPfnlfYchl2yVP5TzTICn5ROnQrWfgyV/dYIYiEFk0Y
XUnzSa4AeG5d7RPSeidfCt4jH5oEqZgfQZm3Cm+O2Zr0J35+XMgtT5zNNyMJ54kl8BUovCb+U6NY
N+Ch+/XaSxgnOYX7mtZ7NNfmtfvTLPjna1XXVWiwmhsPSG3MoeRH57wtratXWKmnZ6tFDrEMMlgU
DdjlGyIJ1pCDFiBbxfTwdXVfw66QGpzZD3MSLuHM0ut1iNhsehz9BSgbxMzxTbHXp6O4M62JYBbO
cTprbU35aD/11aLPzzxWQ+7b1I/vuEJAbbjCWLgapWhaT2Ixoe4GiD8u1tZekw6+mGzx96PksGak
x8nx9q5nwAPc0Q4TRFq0Y5K+1alPHilraqPnq6LxOyQ4srlDC8+L/cWxajfmb7g1ICIHDE+rEmnL
ImuICQ8TE6fjAdleesrG2sInUcz9mVZTMTJSToa1jH4g8UBSDhLQv/ndsvzKIPUGuoEMyAuAf9A6
QRrnfR1rLniMDVZ+ZskcDMJ3Nm/YDE6Aad8wSIMcIXgafQ2P2cMcj36UVJQ8iSe4XgTK83mgcSpR
JAG2gSZZHGyKuoNPQEUlrkkF2o77dYvNBDUKm8Rtq56VCbgcdOJ0/CfwJBeHygxGV3GFiQVSwDBq
N+TtrwX/7zKyfKQOp5T6EOZLsEti2dYc1cIorSzYrMiB0ZyTZoup8XyI8+D6PSvil5AYPRQhcVj6
htuPpAUB/9JzlWtPq1VZiBRYI/r0AusYubCF62Tg8Sb2nQEvkEpCBBftxxw745xzDq7l69XvsvVc
VztT5cc9BgpPp7V13BUrbKOj2mmXzU53O5p8EUEbUWGl5crEzfWUizTSQvVnRcN9+fzDYRREB5gp
Ejl0bRvDx1QH4VnQ7fHMxEOs7vP5Ms35zvORAR1vSLrz1KE3sVHArc82TFhp5DgK50rOA5NP556F
5u/M9WReUdIdCUQ7cis3uzkIsGJcPEY/ktRmJYdYRplZrAJaTH3NjHZqEnzBs4JhlBFk3cFuRUiZ
AzGIQm+RrUJe9EFt0Ti4qlBC01vQJRG4SSMxadIZlypbaXD7QFEen+l7ML8drtcpSNOgzfStg4nw
zVNSa3mbNNnw6Wr+FkWToFZJYUxY+q9xNRgnfCh393G/WUZVJeYdUtKst8KNx0omHoC5Wc0Xus1J
vNYeUE2XFSLnP4gGD6ucrW2Q3wbVc4m8n1sFlctkbKeKXccX0lcr8UbLgZKuIlqwkVRNz8HFB/6Z
bSXw9HQflgworJlzaVNZ3jWUchKcDPmKjYxq9fteDjpIzj9PQxjzTSblsuahKszaQdlW1dG7Me0X
EfHRlkN/FFaf/bzAUEuKMC5F1H3Fy+2COpEzZRBJbkKs6A3U0Ta74moOVz/8MqjkHkWt9R/j98mM
EjzM2EwkiTgr2yRTQY9xIkJizZfpP0FWI/cKUOodcUVH3Pm2dZb/BHG7+AKI69NWba09E6LrKEzI
RVrfSOt/nWrMNtSNLYSICY9CakfQAonxTi9vbSINZZ913qbQwdB4eG4cAIZ68PrzYPO3kpJ65kc3
rSu4l5rd6Mwur5FyKUVsRvtaRcQYXr7Et7Zj9+TFaVuTX4ZtUmSB7O6lURgirCDPZNkOTiMfzbRg
lJg0t+8r+OrUt0WWoXwWsMS95pF8SuM7M2XvHNWxJoAfTttixXhsWYSmd0sa0ErRKGYo1ySswJ7p
6gJUa2EQ57ozjPHxAL9RYKvEOfVJelmqjCrGQpWEhJ+uOlRe5QQJ+8EW2qoLjTlR9i89ozB4EQ1c
n71/xqBprFrxLMW0XFOLTMO+FT7Dco7JhQI0L2l8bwje+6e/sXH1Ebqa32kx2bHgdCPYLKYBZuPv
4d0exEquGco+u6ZNI0JsM9VcYATpaXG9HbKKBHvJUI/PoVJHYZ+tk4/2YRkcrfjBxLlgSD37zoQk
6HfCqKWTbirHKhvx4IWREcn8hfIkUCG9uKuWlZ7Qdaq+TsNYRo0lzKl1ONpgRB95FOcdsHRkQToG
YJgLx7BmJj9+udVy48PbXQLFREU1/OhiHmezPRH2BAg2i8wKRPuIDZndW7BD2zRQgd+btj0aIvll
1Jtm0ihfeKWnF4un7nEdJ4IaVQENAo5rRMRJPnPgoBo+lg85/xl/7jEV8ad6/PzK8Yuad7LdgyDz
8/zBlIlDTwlLW84mLZnkpmVqJdtRT30OkvQOYnP1u5f1xFqS7LnQ2JjY1g96cW3HRnJm3uCLzE0y
EM1iOqfTC4KiOvKQW1eUEx2DChjrU1tDh/wRhnjDNIAACxYbunLhu58nSxKSSMPuqZBwFchv20NM
5DJ4eCoZdwLXWfyQ0+tn36Vr6LW++nkz41h9vIGHmC5NarzdJ21O4qD0DUDE6EN+hMhrzIIV/NPb
P0vgNQML4RcEBigFL6o0eV0B4qOiEMQQ5PXbRUwbh5tSVymthmimpvsaSd9bkj74iq62OTq9ckbd
LV5l4e/ZCktihLXmyMo9WkNpb207LKghts2IBySbmvPLP0WwoxqXKa6iwxXkhtwWrX98bdyCToz3
GRs+Q89sHAbx++W7pm8sGDuUXK2yO4tj5i6qRU+FR14vwXuhZgWy0SrJvx/zrUqfCMpCZyAnul2S
oTmRTO4gwfVWE1a5tR/eA+imldXfywE4PUdswPN6R5C/Uth2lrLApp+82RtnWVDT9VJUPxKLZieV
qQlViiDGKBgT7ccblu2Ckp9pVKrCD0btea2chNSU8USHcqBJAXBrbPkdIYebu81pXG8I7nfe1yXj
s1IdNRPWxnKG6Nlec4le+MDPeEVGv0Q9gyIxJJUYFV6QosQXZxqfLaZviYTPkfFlKr7UfUPV2xtL
qIWk6GGrlLZStLRujyVmGfpaV/+FGO/G4pgjA6TemX7z5hYfq1ViPdEtRYQYQ4wl4Vl7rbwZWbZs
48HsmmzM+VH4j5edYvPSO3WUk8UHGTQzy8iijxDvuj6Sp9mk11GdqcZZegM8bxCDDVIL01WVc8bz
1tHDioRXy0yUHO7vBHec28qA9BjY5O0H7TOrwbQ3EKdz6XK4OtnXxF574OwDIzRcydnfeqMDYPwp
4C3y47s8myn70C/GJfXTJ0eBRqwAralbz5ga4CiqoLl1dqiObs4BXaCqGeikzQj/FqEFGpCQhzNF
fOk3Q55bRycnq1OWEHKRwSg4Yc7bpsJ8m9WeJpcfe7BXzEKDd5fig8R2Yhnh4R6be1FJ96KUrq5D
qAdwRdr9CTVLJAvkuZmJ2Bi2RD+D62BSmv3YkxEZUyVXpZn7KMIlONEPEnW1XAEI2kFZjWID7B6v
VtJ7TuY5gfle7eglro74XreKh9WmxpH1kGpt8njO/2v2ojv+HHMZ6QHhvsTR3topAFDbvp57u0PK
YN/K9yhibwl/Hxp0/qMYQ7gq/27fQCntzWsWwLYQTJ6cW/O8mdqUCCogZqajL67ARGfvjdg++jsD
o/UK/l+N6LtJC42UTbi2+YpzEikF7TT5bMxqBRjOfL5EtGbKamz3Wr7OzhSKWjk+mqgL230lMdf0
2p/7MwSV/WqoJaB2Ji1zQdkTsuOPMct0veC5Bdt51Kr0DiAoNgSch9upkZr/rD78mBUTxZzCFlKF
owvDtBVNoifrFFXApWKcqPaiWwm7WuPUJ496lIePTgVUS6VQvVLLEh0O5Sy9AJKKjj3EQ/utdQ+f
LFeM7Ux5Z0td73VRoyRd3pEmFynR/V4nsRqtHVyA2fVRdCInzvh6nKqI8MzQ4nAB78LjA60GHKHa
fFThEEhOXSXYssedVpClYG4T5dFrhO4U/YBDOojJEhqRZvacdO71Ph7vXsQiS41yIrnjKtXXv0WD
KwfGL6Cxnv6IYgXk/pWhNy7lbOY0QfE7NsOckca4xwNzqVNjRbd57gTwhFYfk/Ia+TQ1/tKzNrjh
UewG+hNoPbqz/nznUl7btna2zLKDeQCt74QfdtKOJzlmoTusiNRR6fWOPAqPXA5U7hxKGmbSyWfs
GXXKZoQccMk0TbPiNkaDkbUYbcNZ/t0/i7D9taJBVNLmSl/oxs+LmtV5W7QfsQQIbs1Us5XtPMUq
jY2Yv24kxDF0LgCIFo+nuzHwgPAv6nSvldtcqz2G6rRuSCWIz9wjQHtUMNwdU94LFxMCWTATCd1x
nJiDo6I9opANh46PFSDvCngX96HuPTouoWR/U+J9hG3fG2PRr/b/RnrmQIuASjdIChQ2D6e+MpFG
oqFkSePnkjGhuYpt+JWZCwRHOT4gfnQNJTJrvZ+r5aGNSP1k3Z2Gqp35L51/2wVxo612MY1wgmdn
+6EbEo66zfcKhk1gcNznHINLttV3SIStV1h4oCy+yn9Lai3GmZTEayN4y2CUsmBW5atEsp5eaQOt
xbVisdJZdmnpO652sJ9K7ZeEXqOD8ZY7j0R5+clC9rqKMsG1LfEMCj4MrMbJkp6IHg0YsKCPToP9
Orq2F+HW5Tz29XvbXkh5QakqugpPk7cmExZ72MwFT7etkOauluvShDiQa9mN+khaRScXL/b/QNV9
Iu62wDCaApKqa03vaub1YgNllxOGL2EEMg6cS3C4M4DUUicUPN66zR8fnh+flhw0ZyDKVjbO6Bam
E9JZbpmHAC8+b+MAopT251bfr8gFTfkQgGH03f1inUWGcOmIPNi3phgH2xDC1pHCSNITlii26UQj
GerJj/xgsgbm4x1lNzDVxuIAIeePirnotNtFiaOWo1IYVzSG5ZQGQPOzQ/0H4vSeGqt9BU4bLL9l
IPq9mXI3Q4+eZDVEzmnfPfLaQdN82jpczDUrVp4zQpTB7RdmLFYIIfcg4heWUQEz/P0w7QSWwJnQ
tUw7nAExpU6kAigeshxBqgd/ij+HmqX84UmA8zZKe1ujmfnx+0pnpVNJmno+/QwKkREISOUblmB+
WTEuAfd/YNcqX3xXk3tPT0Hndn80C6ImQrJ45fKJ43iyG3U5DjKw0v6yh4H9AOJB+Nh83ltaZY7c
ho5192n+XvvxlJ+dv4RCh2bp6+hvC2VxLPpTICh7XKTfdnvkI2e4ChKlFhv55uOy7NWtPfhGIOER
ijhYPIo/hJOnRpg57VpK/ShEvTb1M6j4fjudWfCMugRa5VzpFIfC+jx7aTFgvODPb+ldz3KL2oEM
oX7gVA8enlOilVdNtl2ZREYf49LPvjHQmZlx9+I53jmv3uDYIUZd24e/35AWNe0b7Ko/tRYgAx9p
Brukr7qAjbOeTTZ6s5GxeVRT7xs8kSrD7xelG9YiHeXFJ7UtRZRuZ4V9Ahr1LAKZYcoShRb+ESj5
8yMeo990w7Ib+NEkRTHrGA9tB0W9XyjuTVop6NN66nQbO6+exB0G42k2+/7RN0WISnAQZiLbc4g9
+hERz5HACtc7aEynwchyN5Lw4Y2iMTRPR24xf7p1NuChxdHFZwfomvr7Npud6D6O2Qjfr0uGTp63
lVjnwhgzewrzMgtLNTeZe8lMSTILQSFrlhiaTuJ7+Kgnr0cnGWeFQa51wN+CIfE4Bc5A+RJatRps
BNnIpY8pPBUWs1X5sfD2qIysbjdvL1OrL4Ii2UvfO0Q9BwvERshNt+KOcZ4dAPU0T/v/AZhy6JRB
7D4drfy7b3+KQ7ISF0uDs6SFSyhtBph+cx3eyqiXtZPMFZ+Eluw3abrdGyStRfw+0Ygkmu5ACjud
18HaEEd9k2rP7RAJg0FpmmkPKb+knvuc5LYY6vX1xQi7juOvjOt8Qb47F6YfkoZeLwJfs+FjZfNE
AahUN93wEOSjZLXH45UFcygBDj+JEZzDPIykE9irkNi08TK2+jQIZ6pUJOLZPAyILmCTy+AAKeb6
mUz0bGV5CjZ5bNx3/Ft50xaReh9BnudcX4pRxAJ37ehArEcBj4Ms+CQD3kjjioC2QjjICs7tgeWG
XTqOP+gbuJSkhXV+N8RFwmZDUmcd8iNUGVyUbBbhmYgc4Vz7dkrT3lNK9HyuGhNrKx/snnZI0Wgw
k/7U0JstI/9QX1XtnXT6exSfdKWYgqlR+mGINUWCTrNNaXa6e+MTLMbAbCyOiOq4ajNhod0SSlbT
kJ65HsxuEKHLbhjkLGprCPHX9PBdhiLuTznGBAqkvVadCIvs0+lZV60c9xqSZHSm1Uy7gFNqvTFv
gZARXqWLHqkWzXfdIqnqyKnH1AS/a4XT6TCUNJK4V6yej1LJ/jiLiFDTD6MccDbGvN5nj/QpRY5P
x/kFHc8n6qfKtp7bkRqGpjMggWzBoVmq8Vf/2yeyeX9CKg3YEzFtrvCCLxSkCyILivMmxH5MCO9M
vS1uixGEoHubK63o590p6ufcXY107Y7Tdlgevcqkgq2zh/mx522BjYdwN8b8sOcPXq8EDeT6f17B
kBUITb6e5Lo/neUMRWtgOs+uafLLK9JeqcnGHnP0qyDNfZ8wNE4gC/etAqTcqaIYaRWSL+5yjPck
6sv89Bfkt62Dt6WAH3+1MJjV0iKKj7mnK/M3zjCogugarHPgKzLH0vJs+nIse5mBQV3gJi2A3RVg
ZkA0C5MGuXmCQ4VY6iUEj24RDd5nEqP8st613nhdUWMKXQvqle/yGx7zX3KD0DTlOdRuF4PEnFQ/
8WN79ooGN8X+CjNmQK0Be8uy1cOyKsLXsLLsK81ecWxZvxUntcdFrd0fnsjP0k3/M3q99DbgOBcA
gaPjU0II9KK9xfvqFVERO1RdJ5WN3oyvXCXqoeCY51QjFd8eLNIoNEWztT7ikp0uEfV3Wp2Xgs/b
LOw6ROvbeJsb23b8xzspi+eirdaqF0iL/gDMHpWWZO8Tpit6TZ4p7wfq8nWywZw6sI10puEa0EWF
cWVa17IbfQivPj4qiHDHWyDNgvc5jXNvplWK/dyFrPpI7INOcWECm1OTp+SRb0YZC7yJ8CIj7FsA
kk9P6XiFIL0Sg+NO3REPahd+I4puPIUQaBAw7FTyIiu4yUnPyY5lC++cpdaEbWbfZI4AK/CorR8+
xuXdawdPTcVauPGuxoBohkmvRWwJCEfyXElHNBLcoupNa24FM5HE+Gf4MYJq9zmH40FK6uewKtLP
WdqtOmtPmYeQkwM82NmDC8ArzRf6gwkIK12qlTmEyKEKXBUHxr1pRX2tWUU0kLuuyGs2k/gWkX1X
rIO9acAwuWCS02TCMMxL+HgL5chuF9TnRwhXXAkgTKxB0Flgj69l/QAvyVNp1dnpNoNsDBMZVP9j
A/jyUuqZOdJAC/E9ZA7aSm+VvaWM6bVcbx9w6hUgPbgnB96tBIJbXWaGHELFOvJfPaOntlA1m3pZ
HpdccBCHJg7AWwMjOjO6HQtPrDHEM1QotqKE7AMgnLnrkenqTXjHEZ5GYpadfh6gJxUJ8Bu+dL6+
mS/ajaHx7ucM3l0+7VHvRxvk59ALn1wjbOsw+hUbpEx86TnBxrH3mDdn5Fpf6NAW8oZTUJQJ6dIU
hgsCd64DyYSySP8KHzU37epfwwykeQb2JD+PD9sGQksQk9ef5Ta/RJhPQoJeeJZdMG4O0jy1+lyf
LJrHukw0IQ0IXLgg5wAQOTrxSZJQglkZlqAdw5Lc16QqEnitFVEPdqcpwmHpUeUVYPs1pHGaBANa
wVrTrBiHUulXAXXo7PmVQBnAxymAB1wD+jF+Hd3+I8AN3TO6NBHAsyJoQFsk2r80qLhD7PpyHbki
N5qD8Hq/xo1p5/QrLKlmBHfmNe44m0AxgPfESUdFJzYNDUqZvLWU0rxucnUTfviUuV93vJCXCYKT
JEmkTg8DswCRfDniN2sCuvGtGVCYCy6Q3hcDfShh0KoKaZXGxMpxtm83GRIKDfRA7l6M6doiJ0wU
4+iMVjNclu7mMLCGD0VzzJL9xvHsiI2tTUQQOopZzW4Aoun8okUcS3iaOBgLrqRaYJfAAT4OVpKV
AtO8d3+EhntgvvWBMDIOBCCmHTosE61A+9V983upbMCixKwGH9zn5MLUHVubLIg7y8TW4BUBrCmk
D/oe4m0aNA7sU6yzOyeUXLLlPsHjpnhufGZaNrkBE/e9G3+Stq5U36iN1qMwYbas1anw3IC6dRT/
zPPyBdQLNDmq3LFH5z15SUGANVE9/kElEbxiJt+4IXbiILN7MRJ56EU3nKX5RgdzkXZ4uLfgRRdV
/xNN1/M7oakDclGpKlAPHpMYjuQvTI7nXHh/Z16PGA0LUOweLrX+3MFUndlLgTHydLxcf+M3kHfu
HBk7MoZiYC3yZYG6r91kuTD9EEE3wYB5MWG++s4c0PxwgKQGMrX+esAMGOJYoU5DiFk2fWHsun3J
4eRSuyFyihRK7aUQLtMWIGukW/xbhw8nCAYlM9BUB1YGcimHov+xdnAOjeKi+10rcvHfC09Hnprb
Ep91x/ec4WHj+8UAIeauiu/6DkKmZRCNhTdZiQwcWEkJapX4C5iW7MXipPI2QN4mloO9114ggqFI
R6ByQ79rkbdJPWAEiNJk9ez1fPhe4t1f4T066xLd+aI1U4KIDmNgEs/lG3unZWmTxeulUTG+ftVa
xFHndteWTlE8yRKgbwpRVgIKvLmFJnkAwzMmqt231AU8ageoIhrPPfzQFIK2GI1CqQ2RDF25ppZJ
12ym6RZOO1Nno6KE2p5snxMA9MIcnsAuHWnB5nN635roXxR4f5x0i9N2MtpHis3El97KJtzuQswm
WFWBboJATUvIHS8d6etBkMwAseX6jjEfcx5Sc3mWprnDLbDSXCOn0ETzAjEZ70mw3aKJXQ3Oko5E
VoqXTuEx96wEIRDXY/ku8p57mvkaFWPIedZylt4ExmTlqAcpNJuMVZK4eF7HhZyU2iXf2/YNF2dR
51Mxcjy4XLKUWG2EdozNYDjehy1bgIwHsMC2OCg5ThXqogfWonEp5gbOFaHS54JgJGQDzbyqMw8U
nOr1FaWGy4sXSQlsSvtRD1drgJFa0RJjktJytXsY/Gfd/LlYrEcYyVAKZbmB6sdGvggTueNwj+qZ
BbyhnuUduZQ5MY6GgjLVrwFglpAmch5Ra3TrxTz1110pZIL3WjHvB6YZkqnmRSZ/5QfeWkuC1ygm
4IFRIC6pm9YVbpJ4JFNvAj1M+R2qwNAp/oF56rqL/xzRBxeyfNbxZw/IhfbJKiCXdRaOwglS8uVD
sN1P7/40K8yyRmS1XaPm/Ku/ygDq4BDbojdB5E+84jWQyt8/FqqsRVIik9RqWKDGwDSMpZmRM/mr
KBxlhEm0+NhiGKFuKfssBSKOxBCPX6PK3bRys/XlCMUL0Kb7aETA0qfBRQyhNrB0I3tnr8rop5IT
ddign/qpB61jjs7c/OmauCCn7g8lVJBNkBFKZkwIG0oDFsNjoAI7pYujMNnR1tR/epi5CcW7ivep
14HHPXMPRBDZwR761XvpwJSvbo992Z5EPJG2nrNwJxJszw8CZ0SMABHRrNH82blsgc2NOshQsrrh
NbclCnncvPnzVi//YnEEg4aoqkxXOslhwdvBtFFES9S0Ia2IBJM5R8xuly4icbPDKf1g6j2bhYjz
PDAIK4VzswD+UPFUWPua2rXhMlgVQlKbmkglzS9kjX4wuEoXz4/0RMSMdjgFnXskMRFPa2Pe3e3x
uxo104cwbCoaS8lJ4Rc63l9fKZJFgugh9VPPPjeaG4FtPNFj226UgA0bF1Q4w5zOqTEada5gkCbv
ugJg3YYrrVq/eOrJuRY3q/6IAo+vEmf2KkZc5sKOY655g0GyX8QsKlAn49o+Codrpa7FDPb1Lm79
CmQZqYnfIzgCEhUL+csCrcAtj+1As0Cwn9aEy7hoCHDGzRxXURJcqkGtrehmJBGFeHwFEFN9/WPm
2BQ4AANiyfSHHYaeJcggIdAosQoHbrf5V4gJHJ5xd+z5qgjSV+xE64ZJlaGt3w1Wrmxd8cfixZ3x
qg9fHLvz/bSR22NgdYUhdBEOxCiKmwbqs9avJivZhYKrRABcd5t6Sg5+xc2NzTKziR7Msyd6WDpQ
qRjrSTT+O6iT8QoGGUPVrNlhsp4s/WGmeQSYPrbNOyEiJPFy26DH9/Ssw/lxzRCpGRHobsFxvQMJ
NbokqtwUoxdABTGwzQhf+O1VD0tp9wz7NM5nz/5NKJwbUyBJxll7zVujQz4cbAcUeXxyRHSCeGCv
kG7Tq8u2hL9hbgMAOR9LTrPhtMb1G0xdzAv4FM0nvflTsyhflxwdxmXmevueZ/fwX2+YIMGalDds
mZ4D2wgycwh8+JHUGV/KCAUMWfp+cjbfjyjdFksgNN464buTdIIkEMVNMXwL5aJZY+RC/CMQ5Tov
XB4IO5RP1VNQeErN2J/bQhr6CCNTz3NJRjvaI7qLs+88zRbLQ9N7zS09utXP+b9sirtYF8DKU8WC
vEnakRbeqZG20zGw10UnsixNiyahQOvg5ZY8Mt9RtvwH88S6UoZ7KXyT5qnVrCzwTMqweRZly0XQ
8mstFySclREXUnl8oHLenY8en+9C8VDgtMU3aHMWMhq/In8ccKHmHFoKH74VKWx9B1Drd8m7quuV
POafbVOsaESdAcuJ38nkiA7p6stOC158Iuhv+VxL/ynqydBrHea404dnWqPDv8pHQCvVtZzo/YO6
3jlUWIO94u7i21d36pdHcprcfFm2plP5M1qGrhqD4+o8pC5oV803UhJUe4n0t+98grqW3g4QJY5F
WKhZuAy9rI5CVzBHdj+snVxQ4BMjySonUTejAPNTZnep8eScmsN0XP8sE8fah5qiMmjWseqZGYEa
rl7ea90RzfODT56RayymJQWBo91daPnpEabOHQzXIg62QvUC7lPyMRWtMlxus+nRgOE5udbWnI7+
0bJYeLPxytoeUdn9YnAm8Zlb4XQbj7V3oliO5KgyKwcVDAqdA4DwY5AOuyRxZJmc7oeu3ltaDNIk
Cnhh+gLDDnjLXv04HHon8EQl/JnQa3GYVxd71JrE8Ka56sQWmN8vi798YZ5NxIiKXBlyC0MoPHkR
4Ab96up2NzLNYBOAh0C3z+oSWqER++HoLhNcHioHic1idIaK3R2jr5pUJ6kzddyeEjgUKkn9/w4Q
oUZmLFEX9qxuqZ/FW2OBjLe9oCs2Hwdj+oyMtJUhaSO/8w7F54VA5AN8QvQ5HrnYfxVgxVsCUeIL
N3V1o0lkx0aYdaEQGtqo7DztL1X8C9jm6WfCH0NVj5jMwsTZUg3wRTx9irA+mlZNYgBFCucThSSL
icUx7/ZDgWfYscpIHx0JpgCjFvwkfYtmIcgxUhrZDVsVANpfufbMrPvYBrCCY8FAcJEkrmBLong8
SaASLwzUIUSZStNZIpy+Siw+us0AorNIKt4w97bzyNqQeP4RvSg8d5vfPBAD5oc0BVT8j/UUdXS6
y+8hnFA3Bs7o3oAj79UMq9BrePb8lpSFbuWZpiBGyB/s4N8eatAOxbYwjNh22qXSAJdXfrpcrKz3
aLyKLnot38vJaJjLe9xWcy7QoRgnRs8J0Fs2ZiV2z9/XnV+A2lSjwErUXhTNTBWsof9te8vWjewU
R5gvC6ZZaT6ACxyoDvmdXxxrgRuHV3EGTIOAjHTl34SgkKm7BYdf7y6vCUmyH5PbCPvj3mtx4Y5V
of3KoeWovW42mPXvjavs8y5P9kNU9qjminx21uUrET2AQf9oe4EvzGF5y8BxyRYEz/7o2BZccUaq
Mwnd6FDioOgIadxxP+FYNh1+9Y7XwTfYXsollzTWv8C7lEcBAhejI7xcuixqhgCl2zNf3+lUXUKW
IkiN9VQajElXgE8TF4p3LO86vTp09hWoc71dZ3YYKkc6yj2mvtcsz05faplbXqbqDJOfaoa11x/S
7Du5Tv7QS9BTcsoEwXkM20dtShDRAc5gZuhSEsMgdHuN6/PU+IRe1jlzcFm5GcKeP/jWs8OWqZsD
1WnYfsFc3ky4NyR+hTpwqBvuSkmVyn2oJisNQ5IWosgPouKJpoXZuDD51Mp6V2AMKIcRurJsddFW
H2EQ9Abec2QcUaj2l9pbivnsODp7i+hCikyjlGGZcI5I7xunmrEh+YW2Wzr6Y5EQfmsDCO8/eHpr
TRrfKp94DPtShLldDBygA0GxLo/erH6XJdEPZIWVUR/jx2c22sXYL6IhkUDmsq0fRdoQtKEOilse
W4wM56lWy4aVXgGrmnfc6nwImO45yTfhbDbFs/7403E+ritM3CJlEUXiE3j5s1wZItz+LQsJYMDd
M0woINSsqdFdgy7uq4OiW8Ia2DmRoo0EOe0P6dWW79vi1PaakdNflTmulNvUbjt3BUg+8ASUaH7R
BtqCqzddEqB5BaQ79+OVN+U4q5c7frY3XCk/QjQiD90olhDuIbUV9P3ZR1BXaAIUAXKsmkcAEBCk
iWsIUitiuV1hsIY6XRqXOAv1lKfnDwURU0RHmrk+k3Lo8p6oeRRS+5dRaRb33aQN3s+K0zCu/dS4
6k0O6Xv8wudd9zXkJ6PGSksxEdif9a1hJuFgCrYW4NUzjOKSLyYC8AUQtfqPinEpgG75GRtGGA1w
Mi2LkHYlMKh4kwkODuCzxqYGV6e5RWsQFjyAFvI5iJ0TuPQECe7Fde/DYYU9FDyA9x4ERfOCAsEF
M6duRndA9YfLLT+Q+QqcULN6Gty9TshVrZIU9HX7dsxatscX869Qhyn7vHZTzeCtFVYa4TnwFBPN
HwaiauIm0o0itublZw+o/VorLLI0C+1asYFdYfESjC0rSEf9mBFiZoOQqXWTY2jT3+XmsMFN7AIk
DAnp/dSYymsNn+8fKjU6wLD6W4RdJ3i051WkDRnTI46nHYpySyOOTru5mXbKpI/dO9TcSHiKsGf9
nCLrfor5sB8OOTETuAAlnC0BfEKIfD/LDj1thjNdf7MLz9ql2qS1UhzzyArUg1crORH2N424tP0A
2zMgtBkjPCd2ZqWJfSb3y6Uj6x7YH4mUatzCD1FS6QPG4mjBGiM2GuyPtCVFHqXF4YzYobXzrrO1
em1VKWF6n8VpNfjITgfEkMw7mN2TjFS2sMJgvLlrcsZDpKoRR6JhEGSC9h7n9QkFtRYQGhTYiHsG
KF4DPXZfELZwdy1uO/xjwfrgSxLq6rVjRBJt8bmqJYQU6vO9LvP5wnxw02TnFyVFZDDoTXPJA8uI
dYWmwjJsmJoqBwsmmkydPrXgKSDF1FhFRvzH3rtuMwbyUVj0n09DunOqZav4AVcvWVNJZLO7ba8f
/4XJpyoyCLqTOA+9GUZuIpZgGR268jSOOYEblzEUnoagRfc8oPpDa6mDbP5jn3vMtIOEKQIKDATz
8DEboo2xRUXC3rIUt0zDg2PQa7+TPPaT41pZffrYJxke2mF3fjyZiycDk35cCyswZ6v/tTnFQjbS
hDTn/o6riVstX6MHZUcWV9GuQgQv+tAzD5M+SBfkVqXd8pq4WmhGj2JxvZAIt6K1g86w14e4vZd3
1onjgxxYqkmhCFi7Avqw4cL6+yBqIu7cR/Mo+47kUqCDd2734xC81/bajbGpGZg0eAzCes+i6KL8
U9LOf5H/tU7uGmLEHpFGxZvDdBKrkjyfOLzeLHxgfmEGq71jQ488fTKonOH7LdATqAvUTZs9AYfV
o4TbxqyEb5Z8GWeeMyWoMpjmjWtwPy7bbWSydbEAUBoJcgRmH8UOGqWf/vaPmj8OyySlMaeG9z8m
epv7iLsl9wBUlh9CLGmFH5yevdskFa1IYCmxvvmcxzD5ynVb4GIEE5Lxdz9a1P/ZtzJr8QPv9HSe
LG58MbzdXUsFYPZO9myTdTrW8kwO/aSBvOEhmyuLP4Xe0k93etDEfEYdddi2DbnhvVjn5J4jP9U4
i06s9Fz8Dso2bdIeP06VrWUt9Vrq79MsP4/gvscZvLSseLaWLKoABKmcwjU3c7Fhz58y08rdE6p0
IgAy68iRr8xihLfgQhG4PCQQwPEiyklRE7HGmVmemCqEM2T5uFPbWGCW8FWTDgwnmjqBleFxQpIH
VWLp15dQFgIlp7S0WXSI0HBBasU9tCgTIOCmLM0RAK/zSH0bcXpZDsjgU6FAxNeI6jmDHV81orZ7
9gnT5tvuhTBxE5OTwTjbRYqV+ftwTeE0+AsuSkLBRklGbmsgMhT+l9hs4+MGaXmTrMeJ9pIoEcBU
uvoDJBf/5EttuvCcsBJtsME+r3XCUeYgozw2hiP278KtLfXW+SNAMHQOshb9686uFeHCDSO36QbY
Tfcf5ljojJ2Z8TvcOiCveK5aZajY/7ln64O/bVPB9iqajUY4yh6UKHiLqhVtVVntb+piirqp1+VF
iLvZyMD0+N13jCOED9e6wYcO8iGBNqk5MYBCsVAc510Q/unlJf18/76fPiL5f9kQU54uhgmdPIbU
beK+3T8mHtX6eOmtYAXAQhIIIUn3IJkaXG2ajGD1+wjtvyOalZJUg440IV2KwbzlXX0N98+DSums
fpXeyHwEY+58/tRA+ZwE03zYOzirtL0UDdatBqy7OgPtmB1qevPtNf15RrUPlBjH/qH6qn/D6x+8
olNkeyU2KjbmAEbi1W4V0Hy8W1ondUSk97CbXJ9K0Pt+1lLF7DvLcShM1AObaAGb/7/CmJvfNlxW
GmFYdjCI6ma93BuHsWv8a4BvoD08uD08oLm7xgMoPcItXVgvhSu8GiQXDWFoogrRUTNgwsSTbT9M
3OvPmHYDV/FM7Zx0IDX44/Ce5+Gh1oEmYiEsXzqWbrQOs8ELxhs0YsZ0MMK6cygTgOpwvtBzqG6Z
7b1K9L5a4MDdV2VfVlcwrO4oJdlMeVgp3cphg1qyzBL1XhYob0+77q0P0HKNMt8q6RqLDRbCOl5V
1y8Rtz+V/DPHiv9hba3QyhRjdfNOFJVGbW3JJovoilECW/fjialScoZwQyoLWWAIeQb11w65HB5g
V8Xcv4TMJzySo9RkP9GnY+mKJ0H0wVrrorQDC+DWyvWQ/wLcT54hdsopqDavKxZOjHSTV7RebMhs
KBpyKxu/N6z36iREfbAMHE9T9zzfPlRDbnpj2K5SEl7rgMiPAzm65Je1hmJPbqZ5emitsDlKlWLh
k7UvVcz0a2HiMNasH8Sg5VmtcLsO78iNvj1iNo7GRin/l6vghc8QIOiR1KIJturQHDeSUOAR0Y66
3tyV8ssElUuUnaikahRfoWUBwbZR4ztQXFJ2wzrgS3Pbrv5bJKtT/TqjfcNfeixoARjKQ19G0Rde
5+e8eBV4JejCjAUEgUrI4mFw2j6IYAohk/CWzqtT4eSDv/rlpcWqb3fHSjU78gHZkUGJ9gYx3bJR
BMIZAn9Rk8Cpa6BCl7yvq/aQAWaRb2FjoW1w8vvuzru8yQsXUrMXc6aTWgkowlt49NfeyN9yyzPz
D8d9ldeHgl77kKH8gbpu+eooXkkGEKbO2z590RJYjG1PvcY+gihTgrtJLZHj3xU+YNpHssMyt8c8
UShRyzo4wCpEXwmyw2rNu4xb2nZjlHiqy5Ufe1s5Q5Xx2eYaZqWlJ6hPLbBkXgptqwMKoBxb8/Lu
4ThutLfQZ9l1Ljyip9kMgX7ELZlyvB9ZvHG4rP7ZXcKKIj8KbxWtzAU354vzSabcZoey8EPqXaSK
ctvsSxqt8PVtnRs5sTeYDkHFq7ocYMT76BbC67ZkkNKq8xuy7tcX+l6e/dp+q3ZvANpbDEj3WrMd
TngSWebjWt2Vg7uj4FFiekcTRAMq1wAmc23rA/RMPcWxVEKaBeEsRSawy87FkDirNyU8S1Q3DkqI
UINRel7sdEUc4aw+Ykp6I+rEj7po4GOKNklj1Vw6uRV4bQDyE9ArrisUakR3/PUshYLgDQpnAYbN
biPAij+7rzkAkXDFmvTx7MNoxeA+cdmt3wE0oZilO7gCJ2B5zWgSKnrf368PGe6ZuRBnBxOepfpu
g2+Ptk2q+lfxn295FORQQbzpDF0BCD+VGzIR6Px9oVaISRCwzfhSTYFF6n8mjWgf2qTK9cYTtPH6
ccVBNQikMo6g44RaoGuo7q46PapNP0y2TjjoHHLO8b7UfRw2kzt10E45VcaBkB3b721+xDgZZDhb
YCaeXqBHJi7EtFnqw+lD0AKJnSWkOaAs24Q0TliKjGM13hYkJE+apevMFX10vIM5vK/3pSnZNtKC
9wnC5CyHspx43DyFDqLn66TfKsXn7WM96V8D08w4fJmOD/jzoY3saF+dwuJxVPd4pWMi7IapS38F
1Mcy0MVBzGk1iXcyhMDwxisn1onUKmzias94k+p5FaflNNCqhePP/H7VES1bkApovcO9aQBfTjJw
ewMx/qXbvrxg4i4BGQXbOT3qvB0bDBGM0mrXH5h6+WJ5MTcJt8STyM2b+1U3do6xkqMRGcl8kOt2
O4FZKUR7rm87+wzgDJS3l9h8TKf1ILRq8sd+MgKBsKtaK8BGNATqWUtzstyIinT6rUmteLcvWFUy
fehdampxJ3gB8NWAJfXX1oAFHeoSUybF+JpiypJdXyG3ASIYnYyw7iM93qwXJGuh+dcLd5FWVC/k
OI1I6X3gfVES0XTeXPj8jIdCpgdXcFX+3asHpJ03GGxxxsgpRmbY/R8vzBjyNc+Tk29CqhNWrYUr
tylu1S6OyNn3uqo3Wb3zhtlrLlNKb+TYQCKdFOho9KtE6llcCOzjHm2AdZ7zUlLRValpaoymkqtl
csowp/jFr1xoSfgoEwS8HM5bI83eXCEYArDYXRc/FAOd0WuypraC7TKzb56MkrkGsFhYHUF7jma0
FoX59fajmAqOxZYqVWPuzTJEdBCIH7g9wj00IvsGZXa5RlF+SInorXfxNZA804fHBNJUrDUx5JhP
d/tpRqnkkGhoXT7sQkMe7ru9R7wJhlnHj5nw7p0wB/UEdiuH7q4/cdX6kgaPFVEi5DQFjxfh+Ec0
b5PJnxY/lvTZbICbq7pnzCHi+cMuZlrepkqcJwhVDcsPL698h6AD9PfY53B5rII1bgKZs0Ibhs02
mBR7FzlHcpJDSpIUM/Th9fHE/K5ashs9EqRq9OR1Bhaprva4ti5ugNNDle/0YE/ELLk8kvi6CaHJ
pW5sBW59YG4htmF64R+w/beDFLjjkvGaLXmDDkPuBI5TDXqdM13ToAMJAC7VLCQJY9XlRkv90XZf
VKkYSQ/AHyZ4BzKz2o63vycaka1p2FDB/atJN79QiFFg/UGGnXXgO76PK+9I0Xa4pwhG5Rnq1bh2
np6H79IuExbHiLIh/29BTF4X+bQByptL6LEFTRgBTxrrp6czwoy0LDA745o1ngXI/4oZBsLl/EPm
5jElO3XjcoFmoUOR7XDQBag9UypKVTBhm6Y0lUp0tVlQZimqo+dSMWRwxxxmWoWk/CUxuRHocGfi
HJAKGjc0BLQXEmWRiszj0OnIHeOwVKFtXClh1qA9Qv7lpFFgMcT+gamnr2IrqT1H6+7+rFhKKsUt
m13Z9UxNJlS145yr3PcZRTcpSRopUGvvuKeq2hzOusC5DyReCBEu3fmOxLNKZPCmycr357vaEfZ2
RF5auvT5M7z1jCu9jWYAfZ6011ppRaPnUFwP46OUqHrL+a2L8nm31S9m7hhLlsLER4DZERLCxTgU
WEhBzUA7cHMBMK1W2jtQCtWYehTqoX4oN728ctFLHEvwWManTJBmuo8zVwRGL3eds9JtY+W9MoKv
Fdg5VhxNvYMX0xagdLOt1aI1wqUwGEFOA9CLMHmsPfldjyobq8DYWzF7NI7az1BW3MagivHKioDb
+lzYdf4fd7uy8iTkDh65O/PJpkX034DNZk4GQZLn/2IX6//zohG/RBYp4FelggrBtp1yzhpEPauU
2sAihSTiAnaEbsuzfRlLouZX25MfDXgLunp+LLzxdrNYWO69F0wIfP1seUmfC6WgwzKVHUHRsBDa
f62637PYseWQI6JHj89ZmBdZxTXpaje3njSsmVUtqlkEM/ao1jDaSHd8yg558ScKM8F9uXrwmW9e
VnZaxRiVwMzPijOvDzZ9l8PXk75NxU6q7J1aMaDTp8tAH7Yfs2aAJcFCUPZYsf6lS7W/1vqFI2rQ
UFuIKDulgEgJ0+dPDGts+gYVPFNRhazuea6C0/udS7KgSjQkL2g/Fj3BiRr2gXe+fWT1c1Hcxx9W
gbziHXWhKOPGQSGlLWI+wbv2KJpwe/76CZ//l75L5I5TdyRGL3XywmQKPZPAmZKHwausYJ6zVgT0
GM0YorBfEgU9JAi8g4Nanr/g414zbUcFYi3WnaxxEzqQ5uE1pYAVehKdDEGqLoyPbkgnmOmSHCqU
2jsrVy05J12NpC+GSvJGjpuQprjoTy5NcHM9Nn/2i+MwcNeTsuSbxgLe0pec7hpTY3HTZADtZ4BE
cvX73ApTfmnakSe0/xEGUJ6vvlfmoee8NxAuzbFCXwAS1c5VloXIAc2f6+XcdybuBZo7jkcusc3G
0T6aS84RHepcpsioaio2Py1DKtM19JHikWpKIrxL92D60dkMTnBzEHAXnut5xwHRtD6Cjm9+5uhI
+CvWyZNLAyvWtyApqdoVNdewnguGWdPwMMUiTTUYMeWaC1aA+tienCKIdglNaAvU7OM06TEVt0Sf
POs2QY0bec+DrMfFMnba2yFnamQvo3LiIrvSy6UdvlLMkxg6PLiyx89QpGF01YEzW9ZKadRL2KOF
7FzIvy7a+89TO4GMtnnE35mt2YIybuXjqMdGdApkPtVc76FfvUZanQoZSa7Yi8gaBUPc7Ac611F+
6bVuutubFY+CjU5V/lF52oaOAQxBlD0LEHRzrazq8wMLJhV7VW48hFdy2/mpEqBT/xKf+/JfkT0G
nbBXoZcbh0LEs5y3Cc0HRroHZ7r86hm+waLasAqWzA6oYXKg3sXRYolEcsmRuAdLcvOfYGecuPip
94wmpJiGw4hBAo6pjrLefkKCI9prViwp9WqqBF+jmACMLT8rwNDCiwhVh10xaKcejDWEM4wGhZ0X
+PmCNnhmI5NphCbTLzyejdSca6sLjt2Tdi0VyUMPjtBzwNcuiC81Eh4Dt8/h2h16tGkbxiu5R7uW
LhQD64NqFBkzpXfY9XlQGiETjEJufsFAqTHjMFX3KjMeWm328uoGQoYpMAq5D7Dekf/e0MYX78Ld
suNdF80hxLCDBXrXwyp8YgnHtpZnHMx9UtF/ZcfrJC9mgmTOm82J07MyAp2gsRCF38PmddOUBOFx
T34ZCpgZwpqOJBOEPF7/ASS63IilTqxbJM8eA5oXawKzmy3VPtBNK/D6ODbD5zMgs/6fOvIcVBYG
SOwl4/dKu/rbjHc3cuhqaVGXIbYEhwGuvvxr7YRhCPJ1JPMK4WkVbLSXvcz0TVmlpqk6JdvhKCHs
q+8PXX3HZSMKYANjgsmAfts5Q39HegKT00Vz4Si94zX/HQj5vKXuDBN5sDgCQVrc0ygbN4ed5MvM
cAlmSLIEQUWa8MNO2nYZYHYRFF2KN7NomDpQH1S6AzQJrmzAKQqzqB3hILfmdlwtRtmI2lxqIdlm
pF1cwRpzNfo5VwD+B+tqZ6VY7ZNVZPmHDSngxo+hNS0NZv9HdMYP/AyJwHak4TL9uIcB4GrizeL7
I1bkch+Lp3vNNKAXx+FJDPkHwuIt6XPRb5GzeqdNif0vyhgApvKim/ImUhn2faPHjbf2WfMMSV9D
2t0UzjBB0MtxdIdTG6rpNgl7gaF6aiLirswWGGnzpMbofUTi1MOPB9G6TkknkAYr7Zb8ytPkH4Sk
1Y1ufIf/hdfFzlKmKOIFyKiOF+Fqswii2M+wHux8CxJh2vHD459GI3Zdt2jrUemeKY5RMXpj2T8V
rV5pqmU7bmeFYQKnafvz6pKQHSSuCloXU2Tsvl31yRl38YDOKknTapuHwWGcW6/kQLKxScT3gDO8
jsCEB19umQCI5zukWvLkZXfQut5v0SndK9mLdNey87HqqeV5iv0uivu+VitMo0H/1Sr0g+tzgXuH
9GpknT/mzcTg+f+g8ZWqkqghEmYjELsowu08evJ3VdsvmsZH3MxA/zwnIq/+rLPBo8P1eaCBkLg3
no7ELDVR010T+WMre5Z1hRd7EBIv404yyT1DQnGn2wFdBvH5Dqe9haL8cvAAqsN2bpijrftasQ0r
oU+QpzkhvUbu0hxI++uKM7/qkMYkmfVdljnFSUnmIyv9LrYRWTkgFnbcKJJlrzi03h7o7p9MOpz9
GkRZBPJ5UuihHNKPheYsw9YP8UOj3RAMGK1Tbzmq2I04TGecd4rYg0QS46zAdgiV8Kj9+vs1Hhq6
pmcrNqdRE5xy+XdRpc/wAB4er05VYrWHFVQviPSAR4JktiDQYQa8zx+KEhp7Gs8wDLqmXq+pZMnn
nfibLZzSCQkKfJ/uUFzOu/iGsU8cTkUIMo0B5jV9LcM9O+MlO5lWM04eOSlL7ECyW/HVkHFOP0Xi
hPkLbujMk8uuuuycYRm3ygXOHPqCoTbKrw/66TtT8282GqSmDA8sR+4J0vqwxmxJ8FE16mAAHBHw
hdBsHw9wtFNvV79O9gP+4aZz0fTU6eqbH3pqvJGuxf/HnOWwbxoqXZQub97BFz+XwOtzYaoSifR1
7YDFZBmbiB/oyV+Kt0hJDJs2u8O54NoYBcP+oPqaWBOU5OetbvoPjCaWTO0s4t98G5Y0KszE+uxi
PhLIx0/KFlW5Ise6O+WnPnIUq/zSgQZN7TJB+eTbFH3cLCNd/6rq9ecjxF3HFL8e4u+aUJQdunuB
P0G2+bPDzo2JZn0D0F4DS8C64vi9++nbqqG9FBfJ/CxMqMmlVp4OBER4A/qpuspBSNUGYi+ZzUme
N7aQS6ibl2DkXdCVeoBCZF8CkG57KcwCq7KlDxTk2dttO7Qk8Tuc1ck+EQQAbvp8YxnvLXVd2ehk
ZW5mydC+Bs2RpyOKiJJS5HvHIMX+AHf03ijsBqB2qYvpDNQrpXeP6FEuNA9wrJdp4xV5fJD7Lk2D
mRCGnus2z8pMQ+W9+FQ0R6fBgBTq0VpfBaGyrveecSpIEu+r0p657QsXtVPmwE2LJzc9Qs4DAEDF
okjOO9wUjbP4otM7zVsXQzxh7ZJc1WuPzC20jQweHm+E59xxOeE/l4IekxyfdL2BcOJUi4M2/J+N
OPixC+cOEPllmh4FHZNizAEH3L2omTl5kiHukYuLb+BUnA9Uf6nT9/zWgMFHEWRHZ+MTuGYHwX5c
HIeYe2TKr0TYGMyV6q26hAWIyqjjg4l7mwFABQUdKfT/oeE4hjGzAlDUiosmouWFhuFbILd3eDl6
8mvlvpK3LhrZ0qYCTc1Kl02NgUjTnfS3ec1wHF/IhRhJtAc6weeWUiypKdu52Q1vJknaI3m5D9Iy
wBttLk/GFz0TSRneZJVf02YiL8OqOapdX5QnQMW5eC7N0KdxdB11/l1P/99AV3s1PUUaAUoS2JHE
fI2TCU5SipL1QypApVmLWZ0G3ioehz4WBAkTey/+8LSBCNjPXFEIWDC+7MiH9DE+U1rhnpxo5ukn
u9AqhXeI2juJJAk9cWjlWlaVCLsg6g9ZXP6k2gvNp/QgIZRJnfUeT8XNyooXuDGfME5e1FR2rMaz
WNG9Nw8kxPwzl50EPOVIELELJ+nduIuvtS5vYKg/K/z9KcGWc9gHiJC8BViywn0cQQ5ujHNr9+58
+rBrnRrRPpw2opyHEpLRCYFHS+jZOJhGTbjYniOzDm6JDmeLpmklLApw2CzdaS6pwM3S01PowCHG
Ju7oFPoSb3xKikwtVp5LKyEVmrJNM2nO89E/FdsU5gjaodi4pnSVtODo6wUNRjDYPqzYUu48cF0A
9icRr0TmLxcpEDAxVUjnhEsze4xVKsqOls8ew8VcLRHbjKt+kB83Y2RrWq8tZEDWeyx5TXFWBSwG
YcTHCMF2P8+GrL8vsrPqsil40ah1ZhK2STlOs7MW4SRUlN9NHOZme14m2XBbGe5InTwVppxhzWM8
ZKQA2yybO2PvH6oy7RtACyuElQqRtzVOjJxYlapEcKhxJ/AHbhWpeu0FSkqPn74MSrbt7Uw2a5aZ
INrlaKj9KhuKyClTSOoDpiuW5JYyxsUi+mbIVzsA9DzkBruP5OzoIEZvP7PyDuVHm/0bZxvD76YN
zK6aVOOVeov6AcbXbx35GKM/lO601icbKTL1TypqOOROr952Jd3Ty/y/Hsr7BNaw68zBe+Dua/el
sAS+DT8h0ynB59ouHUDT3cYydx24w2Cx9mj+7ltad7zazfKlXn45ldHapWG/3xupXjkxPNeCki2h
3//GgnpoU2/DALZMPaiBco3x916fd77rs20Jn82ydxZ9E9poeHyPYscXMxeOV3FPon9WE8BFdkSM
t9rli72w9in3uWVPX0LFpAr29GsfI9uS497tGm2fG2fAeSdLEBywt5NX1kCIcDswZ+qOWEVbrBZI
ht2nQ94sZyaoHOxTqBmk0d6IE0lh9pmXtnAvUq2ckKovERnQrVVP8QxGbGa5iJk6xEq7VPE0qE3r
Tp86R9NwUe1HOweB0UHQThZ1H9+D9/BvJkYxDWi9QxkdWvxAXDKul77Qh5iUi3dxVzYmCsz1ySVj
D9HlzsQ5xkhvgDXwjkCIvO1pT/JL1GTwEfiProxzPPtVP5oXtFXVIN4S1UDTPMvpekzSvIS/rAt/
wsGWhl/MwD7w8sty4yOPcbAx9RxBu6eGyc1wm70/W7ingtTRYZ4gkbil3S4gLYYqVvp10vBoXHDq
bcj0RuyS2kGYL7Lp6FqQyRw+Kbxbo2NnvljT9lQldpzew2EeAKCYCx+Mlwe+ZDGZXccbbzONmU3U
+P9qhdghX5zyOVQmevXIIrnZGZs3oyvCKp55ELab4A8IvbMrLLumz5cG8teGMj0eCrh1giT0Ry5E
LUzypt87STSE5i2kSIgMzG49y2SJ/JJhalao1caUZqih4WHO0TZc3mMQCuEuhm+c12nPr2pYfMDz
i0UWlWm3zMPhX26TyygpVimYcfY3KhKDKxYkllhE7vr67SSy20lpZoxXjCNB/0V9waXrOhceha/X
HzuiLz6IFyA9xOR+iYCy6SsfkCCd94uMdc/9CQjO8kSJlcUhsuNtVvaMKkFnapvOmHpkXtwSpOjF
qVpYCWrW6H6UklvYqCoxWmOP+S3tQdFyk7+aU44eXuymaWRg0zgxpMJ7e/fsC78UF+MOifKkHQhn
E3vdWT0U05d1r/zZpGDqld9chNhWt8sCtLSG3vtO7O048B1cHXVgLOBZUjV5uNphBqB9XWtPvaHN
h5df+l7qpTjnHAIFcT5Mq2khnhLX/cED1n5vHZnaEHBDcHclYAsqRCIeiYP7qA2j8eHUYgv2J15c
2NTrSOFVc8y7oECyFtemcw5I++yLipx6YqMle4rq1hzo0PX2tuck2GdB6QY/D5MAfpr8Ka2N87fI
WJb98tRnnaH2GEo0KhNeTz33Ryc+GDxxpRYXgl+p+nOKOFj02XCZv5vaqM6rMuV39YpTy7BCbXql
MJCaGKw8xLfPt4llzgOmpvuZNLgzuDoW7MzlY5vWuskvltpRBdixvZOvYp/GHywvjFfquv43y6AZ
LW7sRu0rOSSK09+QTsiP81ASGRT7caIBIpNwQRbG5fOZazs4ElqEXJkzMdjEMrisTEnn2SO8yFI0
ICODRTljvoOcS4HePTP5fm/LUHddRHwr/W74uj6WyM+iqm/MfGi9z7RdeQVZr7z3zVpGOaN7vf1D
Sm2blcPabqbW3+PvBNFxK17xau+qKOZUcIW342njPKcEKPQ8zJkWmf9Rk5MzD2tPE5/H7toQETtv
jidB2NxBGGvSYtpNKTPyGaXtThvB2UyBuYjdKnQaHMKWFsrQoBaxi3TZcLKMDHj89nUoSuu88Vfw
RpGhzoxR2rfYToFkGZZisE+zbt85XEfWcVIztFO9ezTa/KxldZ1xiKJeGR5kKiyh2HN0lgKejvxE
Y+fsH+lk7u6aXp7Kmjgchj+uYcPqScbGBW08MWAEyaK52n46nmjgYMh1jexXY42rdKJrekwR4pG7
266h90PKqQ9mby5JVUKDE5arxTt6Qzs8dG+c2fEK0w2tEBeZy4zpBi0MU7dGdUKpsov9Hi/WLgwf
b5UaCpksAriKgruSOGWno2HFENLXEomTC0gnD7pMXHsZFCOZqMpnccVirim6EpBpP2tzAw43rkZt
dec9ypT14W0pCCtYYtYQOFyHn/QvidHSZaS3UMBf/jJRVZFeUvMd2jPxlB5tnwZWhXqzMm37CdHY
MSLUm/m3o81cHYYLP8y/Dqat4w5qgANkRtJQK2vSOeEqZSatpuiv5fR4foafUL36wcV1Y7qBxBUX
7sZo88MY9cZ14zbDILbRglHDQ/TbYy8tGTyOYBs3GtX9fwep6gFis2qyxFFi5V2FM0KXPbbkwWzI
3s1phVdUx+3OrPhPW3u8H34+jq0PvWMch8CjOeydhUQ6HlQ/O3DHfbBj3nM6AP6mIvUInTSEOf1x
AE5qQqBY2Z8DG8FDkGHoSzYxPeMKrvFwKUr48pwYl6eDeDzTyll8+8tDpl2abHp07xmkh2vSemCF
3lZytGxGCxPU/zqwpSZ2L8gZiQWw24+aXa4YnNpAHxKnRY2BTMjjmApWBhARN05J8AtO0hAlX0NR
htKhn0hMX+dlZi+WFUGIev7At/ez9Z03xg4nJ7fSvtgUFtxIuhAJZ3lLQlK0EO2EJlwEJVMG9oPC
YW7qJ/K5E005htAwlUhzFYqp1Js/H0gLdQMRQgQA8EWE52lf6nHGpWg6eXqoVWdPuEDiQoSsA7+C
/kkH+QHhJ1uGkHX/Whk+C6BssxYe0JOuhipIghIAGC/bcZaBnsRvT1n4rps27sZ3KvEz7i9xCd9q
bPH9lubPoi0WxyCsnTjTtBSBvVYA+1Ax22ehGcl555RVqoD7H0V4dSs/djtUQJSa2E8cQYKNn62t
QKWtzs0CpcsQ2DgL0o68ke7bxz6TmVsm+JN7QAEvFLxMzdfSMKG1yc2awZG97zy3Ekxn9PSv3vG8
h1HoS7YkapgDvJu9T4NceL0Gxl2s1uvazGqNq+G5ET1ud+a9+lRB8Uk+QMGTlr4F7VTsb+dGm/RO
xSeeamM48I6xZTIQ8qL0Jcye/GkLVhqa7Ooa6muj8ML45oYfmsp4KJACz/0SiLB3gkEDBLoAoNyt
eqXgrOHcNb09C/JSUW2KEuu4rGG/zsxllCHiHfnvJ04Zu2ptStIhV8xvg0fmBxpI9MXE6AKulfqG
F+Pwz+6kDisBIgf4z422/stTYrFKfHUnb8EuAajyVTa5phxQSbe96tdyPryGw5tt3zLYwnosUZ4Z
Jq5+PRqLbB6MbEpcnJTcXNPDnIMjn1DyvwjwY5H2rik4v0K7Vgh6wZW2HZAeaLloL0sK1ChbTrKy
qaGDl2LAxsLNOO4/xkEUrDtwosEEnNcs0Berm8XyY7k/zQtca6atS/hZu3bLcugT/mO7nRlgFOYk
mvLWXFBqIQRDtUQ4XzsbZdCD6TN1k6kA0H2YRgFgrfYumNAmkK8Mc1e0j5PByQFFUuzm1VldXMks
jUYGdK5UcBNJmk0HetNJ1i/xf/psxLDcWcvltWzoEhK7JAMzsuyMR04Wa1FovDlk0UU6mNBcOkPR
VpAizdUfsTV1OPjgnarHphBTebmV7HmWAN+fMjZpTfT63REASEwLV1GRCKfZerSQA9weybfQsKfx
sEMbezB8tcKiBDo/icvVkmjLm+qBYb2h2J3OlBoNFXLR0wI1AmMoH1R5Vd/4RWllArbp/k3a4m/u
Xj1WcgQPqcDHTYad1lwe57in5/QL1tiEJhHuaYa5V+zL4iiNSSFuhWUHzN2sxaZZwgdBPfN2Y9DS
iZi3xG6Tuax0sJh0bbPKfohCrRw6jkPtbw+uTOhgzD6NF6Cpv/ZNO94r7nWYrol6ryPvrb7MTadq
s+YTkoT9+ak7xXxcmVqbJ6f7sB34mcdErbqYPe4kl8V4rlNbv8CRs9a+CmRyPKam5eVUiRWkF7B+
JhHZC2/KYKjWbCkAkkfkSF1+eDmrdZ0gty8PARaoqXT5em7PQ6qHKWviQzycbuBa/4fG/Nn15c1x
qmrDPRjD7DvT2c/1PkZ7gmTmvgTFDtNQcOghjSU554LJSYzd6VXO4khJlZBsAfcf2Wq3pdpfR7Wb
rmfYFKu06QxT+YqUHZUsoUG23eNr3AYH45Qh8S9bjAO7lniIxBjPrRjXNVSqow8t3rdmu1MsyvEl
Z0Y8PQeqrSGD8l4mM/pMZzSqbw5SPuMVroRagItVd4FcsakoSIsHsvje9hJc6DtxILHuWMdukBLC
MeXo+4mX2BstNAu1Laqz/gnMGv/Os2CXBSM9tNw5/MaI53zIZbQlS5Fd/8Nc3iu6R/aX3kyuhu8E
b0JfTFlEMqdt1/s2LdCsLxN2Uv94te4x9dX+7LzkAD+QsLTFUGCSCpuVo3Qn1aBNzycJjRwzOUsa
uuR9o67ZiypgYgvDdnAfb47jgZd61d0oiCdGwAWjUXNb+hykHMNcZzfTPaJCwpQG8lIYqFvCejRJ
WoEwFDX3SmGFLLdWJ5/JAdNi7lbPaQCJA3gIYUb46ekfnLUcTCJPQnPX2KILYHGTHwKP9pt4qZPb
ozTffU/QMWLRcbYnSOeKaWe0nP/anu9LUCEj6TvEjNkCUrFU/67YcYO7DfY8iUwk2Ye2LD8r/vKL
EHiwV1QQ8zf4bLdnD90eoD2wOW4crXHQhGIABC8QTp7jeTOjF69X/6ilyLAFgWG2LPGrrMi4SkIm
ii1T0RtCPZgDsecO3NMzhNvvGcZizC04bZOw/k35/5dWkI8tnfrwdY2pQ64A2XEL9q2kYht9uyAL
kxILXusH7VAkrB07X7Qf3PO87tEAzmHAyRwT5WHP+Oa17LjtMM1POMa14Obq0dR2KrBfNALiWJt8
2oJvVgBGS+hHljdovurmFjHd/BSNv7nYCaTy/PI3qPvOgAoijAavO6ClY3mXt+Kt0G1GM5nOp+90
M4rJLk0X8tSVE/SiEyMK/gpzc/8iQ/0wWAch7I93UGtDPAh5I/mVuv+EKuqkbpq6wjzY09wnnMLb
r4pWvIb9W4Oxzsy2xJOc73HOoVl223nubIvXYtqJ8K9qtAO8wHfwy20o68B5g1qrAn8IxFSmLEzj
h4lAoUaKZmn5CVEXJhPfoCyyFa0bKEISN5W+A6sshUlQnsXyy3nWUsQejvQvnp3OCi9YD7Yuh6za
6buy8G+kN8jd25bsp+q97ZRCkr433SzbbBVrTuBgw4maWBSU1IlsgsOqDoHqG+j/271ZpTPbY4do
PYTbQVg5e2J3Kr/aRh9lhzRAB7QVWnxGFk/LQ7yoIhKVv3XTiUQ0o1qI892omwTPCJ7vjM4BdNP7
e2xNy8ATTuqjG1sUi7gE8cAylTI4XpUd9MEKM/tatfKMWsA26nTv6jAWWgUgdB5j+eLweDv6rGH/
lRVFc77+82SnCFZrt/cvbtTWwwlzxBv+Hz/jh9bkCzr71RFR0m8vr+v93m4mT+O1r4m7pN6HoKgJ
qlD1H+5X3XtK3+KswT6Lrg3LYkKScJJALlNc1vKOOjCkqVPBucp9Wdun1dmW7g5eoA2qdd2HlSHE
7EIow1yffkyBwzKYHd45LuO/1qCG4oxHYfZyIlInRJc524+tL6jXTZT7oPDCZfMUk6JXxZIEi46Y
y5vX4U32bIi+VMRZPU0+LOmn9UEjrFRkuJl3xbzAV65TLK10oIR8pb8sUgqQkTuBtLuq8kaMm6jU
CTPi5/fs9pYt4OflgSo7j4h3sUZ4FO/2i01gTXZRvIiQATsu7dzdiCYEXO9CWHwqeq3MalYqFhf7
nNHW8rvHWbEv9N+rRJdfTYUz14VEFI3xDI4D0jdV2YRYGLjm7fjMy82V/7lEtrrN+EBJ8vYaCKY0
10J2ZMNt2DdmpjP2OPuprM/Cd8aYypoqXR+fZfjuCiVdqcphL9NzQLVfT2NKsK/GH7yUmQHJQwUR
r74ktVhCODJcdfoLbVOcDUCaaVLSppo2haSHyFx/37BJg+IXafjbw/GfCOwpE+0F10IQ9KGWtxF1
3R+L+8RAijw6hAGTfZqK7D1TFhYT9Oq3KG0BktpD5LIsU0A/bKpvLpl9bvZkyWUIcKrB3ypKj5/s
pvHGdOXKDYbnhD89Zh5poww07EgsWQlbRRH5TbJyypJ6Sx2NaD2LYal/gAFqBLW2brEAXdfeMqHp
0/LJKvDbN+87YUp5GSiVKh2IRHPXUhftnbZyq1WZGnLvOvIxDa+7xZiw4E38bIYklkwWIibDYady
ghaPCmXzneFZ9SBbPNpA7EmanphH7SWw8yxOUVBVaitMwq55IpWgDtD8fpniqIE8iC+E2BBQIIP5
2njEpBQt3ymi+2j2DjBurjCK+t/7xEWHjoRglOzIYTD/OgH/jOFIp9uqqSF38JoNiSyVUSNEdXCt
I0evMBDtqt3lSz/xkIKcjhuk7g6xM/ObrWAOodrwpn/26XV4F4jaX7JoGEg7jkxjHE+omenT0MIE
Q53xvaJDHyhfNIwDmvHYXwr8AhdFnbll5v3M9MF9rPfmailU9a/Vxq22AgLjZg3fxPb35fyyPUxb
YhiX1CdRnm+3dlDOW7LcDk6YfCdZxiVzMOVZUWbZpIdUW1hqZ283Qb6SSJueeEuVJDaYXT6EWccq
QtcF4JFSAzmRzXLr0+5o/yHHzdOKQh4RkQEnpWfql3tO/V/zHReCIPXQSvE/wcS8hP7oy+wwkNI7
3XkJrxrDQ1WqId4VXMaULhqoIMFhiraOBMDPJz24BX/EOkyjMmTzwvDIeglmcTaFnhv0VAsIttjQ
110zRjbALf3yN6b2e+RzRYIIkxqOtUB3kUAgz8iD2rOjXLRzH/bQYrEvFGB4FBOjlsz0imYNU/Ga
2R/cjM1OZkOzfTIc3V+XlyYj+clqoZmIkxW40o6WWUvsWgtipBRbxb7rF3aYPEYttMHA3auH2v+d
r8ID0Q/4u6Xe+QuY9TV1dRfmqpfKj4TpXDZWRBbnvM1d23kQGfugcyc9dVERmn1qDH+feT6SUCCx
2CZrwDZ1bcGAo9nvWuwTYBk/46xDyrVB9LMHs83v6xbKRbMjCvYfN/qLt18GrDkcZ7RaIRTBZY3d
8VFrdE3LMvBOEsHf1R1Q3CLq3RL0HlerLp/ZsfhZMD7JubYQlkwClMQNLxc/uFwpLt9BpM5OBVIb
0rw0MVmFgcZ2wa9VURGpjx54nrYClsCJ8yWJwetViKtoPapgqa2ETkaFuZX+dMHylX/wCMl76xrQ
+t54ENIJ1oz4ebwbHjtgD5my18tf/m8GJjRb3nq4SdxtO/UlF1jiu4AvXOPYZWQmd8ETJNOKBH+L
mXjVnRvNeAheBIUrEmqpv9b85O5jGbkdB/ADYGdooNA5YDz33XFy5ZL1QhTPYtLhKuwy8Re4Ya8d
OtRMnQvBojQSIFffG+HJ2AgntV7uyYiFD4b+t7ZIJ2FoSsP4jTNdadZmLnl87GlnmwJ1fqrpEcal
sp9cn3uPeSKJUcc8wYusk/v2cOCWftXjyy2naW2BgNQldAzJlGG2j3Ug0RyOc0dOkwsdQt/QQryb
QM3OLZP5famuaELc6k1uJ+9CoKGgsGZoMZo19s0Q4wKUoremnFQkccQHJPLtkqWu1a61F6RnRRT5
cSfRDaIr9lpMWEr3m0Qfbp/FYdtdNC3ILufTJyTubcbP4eIaLeNiW3zSQvDFK1rbcYpwhzGiMAec
h1dcLP115uMDptx6oODHph1Zybc/2pj/f3UrCohVQFOsJ0bSu3kRXZNekiVKYG/R3OBxFr868pND
Bjn0ZVUia461itG1rbiC+NSDo2To/H1h3qKXQEruF4AoIyhiYgoBrgV/cnF1HCK8z5w5OhHTwW6c
g95ZnXl02khPSkCAjUE0iY0NzpcJg1cCnCv30d7g+lVP11ljkeJ7bXoVFITM2I006yl03Or+/LcJ
zPx3YdJHEJXjPq8nloZMOp8X9bFN/aFeVAbgkFK0nEj5FhXwZd5NkLkr/C95NMADZdgfUhYXrBzD
mgLRtlbPyAKFcTQDvWGIH6V0j8hjAFxkfQNgAGG5VOW32OQelCNqxnI3g4qJPrxbVBf1CmGNsq+l
6PHRc/3P3UdbqUYFmwSqTyhGyrU1lOFD1LzM2PNVUJlkq9ohtMk44wXfUyQ4nQmbJKPvX45DCjj/
P3caclrcQdSdeHyQD5Dy4FVCzXYNlZQJ04rixxr3nX4hiH+0HqBfyi1IF5LawTA5mFnKOjg+NCtI
D0IxjeMBuWYEXJ7diKPh14GmI+CeFrXEy3IBmowVMpb9wZHm3wAj5yne/jlVgKmG+Apryugyf31M
DMYitN7ScGdGdKBu/mJhmbPs8MrR6Ly68moeaY7NqAM4KOgPF9ETWEZnGoEi1XBi0RUWJHrlK9H7
fOzsQPKNY9XlYjtA6DOtRUZB031whzCNFcZ8oYUwk9boqzP6jOsxqgd6jdjmEK5aniZqtjGxng84
gH3avST46xJw6FJaLZKuCP82BWi7YIGMlEx7JanxAU9liFe67EsDKzkM0MA/WsnAD/dhK/MxgSYd
1dmzo+IOI5ZwIVg5WudhZ+v8Nl4fyFqAmsTAecL+lSsba9hwKBtQpXuRi8hl3tBFxly+ZCFzC+vf
vvT2LUyF5W7O5eQFYli+0cYOZBPaYcyGo2FQqIKbKscsz8JD0x/vSpBpYO6XJQ8phYXH/7fNJyOh
bEjsgGW+UNt5QvUuAZSjrirevbqUPu/3R/0XfPSqfumkDLiTQjvGAxFzIgioXlxpBV3fXtaLmko1
0MqYgZ2ImWEOawueyDRYmoDJLYWlOfB15m3fHUf3OTyaanroHV9KNZvxZm7ogKwtMFBlnqzPEU5L
UoNqVzd2jvMNanOIAO/JbMHwnFCQAIUyh4pWzWvppWu/uOrvSwbv8+2s/LM3h/udW5T6jOS4luFE
iRlnp2K2NcnXbSCmEPIgWA6nUfW/OSl0HmyKQ0oE2cxznoX5bIbPofPWaC/xO1AmnKzNa6hgnpmC
IdawexjtOdtoPhGfHU/qzZpWZ6/Z9n55JJnCy50y1i/w9J7OhSamsGVsk2JOs0moCsKdbEEiHWmS
LL4YOxj/q/usVakquEtp20o8nUaAKj0/ucRf7ukcqG68nMOwvIrm+eRsFk5NKQK4bM0oOM6Mka5u
t55KRAeBhBHW/cAg+ElCOZo3nEfA4l3eCGVzfLww1vUavdEAQb4Pl3wkSFUxOeaXvuaKibAvmajW
BIjfW5zuRUOOF6w1wsm8r6Jrs7+GXb3bs5HGyq3VAWMaMxFjl/LHGlcPvpAGKLRDoLnsSWxAmTBQ
o222bFPeRMgUK0/M8za33L+nHpzJlAl/kcX2/6b2+a4KVA0nSxA4WrExf9rnDK7F0Hhjx+dFKed2
7rjPIkpJzeseu+fD0jPty1IZh/26ltsmx9GtKvYvu7viJYQLJeUTHPJ6KIXLvfJo52zB75X2q/1C
b3pSi3e+e0UIcrZaEK6Lef1q1vikAmiDJ7xsjwWbmMaPk32+038QjEYJqZyMZ0xKLUQkTb2CykzC
RIk7GbTwtkYq/XzGLHwZ56rKLa4Zh1RrNvcvJYoiGKAtGUOTp51BKy4exwnJsveSfWTKSlF+YlnV
C/LUsmPOzTZMzCP95otUAuWuPnPNgD8KvrIfdKtZLAbd2+2mgc0gkUN/XZOS5Ev3JWuI540hpQDc
DGqXVMLKcCUZH7AszYGmf0pUTB18edzsiamvt1HKtYp+MXU7pm945wagVsw9DuIFUe1Bz9tDT62d
EuTcq6Eij2xsaI0IPhLfjjJYX96zOSLiyhBB++w9ud9QCRT5t7juEWHnQeZhMeJ3Pijpp89nr5cK
vYIJkd9AsIddvxzURfFZagZVITl9csCIrRISM+2lOu+tm4TT6KlwtqpJf4eBKJalk60WtU6yHUg2
shHLZm+d1AX7FfYCPPcgI4NUqPbnznrk+vCiIeYWrIIMCyMcvcONp1c6TbFP7cXlVMCJHE4eaFII
Fr5E8opMG/ebYfiKnZtl1hKqEyIUmFfGZdht5O5uxDAmaJf/2OTpMtqFGX+QpCxG4Gayi/4QK3pI
+es+K7OwBhTcXYXuzYe2pHPau/TamiJG6TIICuBT31k20Nn9wQDdQSc7ZgEQ5cTd+9hes7uVkabH
J/7fMGF3x5puTCY0qYDJLawXVsA+e6SYtZop+EWsgpyMh7TDwPUOCNNmJdMD2jbvBhw9GplkAy8p
zldhaLpF1HE8uW6h8AuesCOTgCO69y0zZJddQKSrb5uSLVoTTM8l63ze5ljoIPKBGl/3ztdkG0RR
hVvLJJhvsXfpLmJ99uRKjQOS3WF/I5cwNAg997NZE7ncWG56PK59+m/DFcWmnvjyGQmjbP575VsL
qa3AdqN5CAzNZeffyQkE0lmFWtk3FF/CLFnFdSSVtjke9UHnZLfgW+Npp9LJA+ed0ypmlQKLHi57
yAwfF0bmmow6bGla0RaJAP/HXGpSV6QpXFcVBtoSlUrWK0Xrrr7Lmw+En5jaPQ6TCJj6M+jJj2w1
FtmRNdspa9YSVKnwReCrUtmo7aUxiQtUCQXgDb7cGdS/wFw8s2XLL6V9eaPa7AB9l6/DFCV+5oF0
OoLTdoep7FJNjh1HGPmJrfINLbXsjjad1QQ46+FkudHuhyzQZxgVzzjNI0D14IvQADkOr6HV1cBs
XdR86H8Kd0BbwXViP9ynAgn8JVJBC0d3xNXtPKx2gss04fauoZwaAHLIR13TlK3MJqMlbBCXyWCZ
KWHbFZ6ASUQLbfGWLleKr3uvj8Iemz1GqeqPcvaHe86gRbEA9V5oQIDbEJcYPJzSIYvbqu6kKdjA
w7Il4DtsvUsUNwnFqt6O0gFqq1MavB++JCu7g6CdHU4RpznnVjjBSqDpTlX1/WxN9dfc0OhgVnC4
tbKpwX7qshrLDUX4Ja+QXRRb7dElBswhAhuVn4nf0yuY/VSF+bGEr5xakNJW5y3oFg7xzFncmhgY
qO6rDbb3ZA+8u0Frdgo/HjxWC1bD2Zlfl6Zuqx4RapAy5fihNIU4O9dnmh2xq0a1Kp2LhFUhQWHK
AnsNdAjK/MG2q3FH6EL0/BQrQZ8ZjxY5lec4/MfXUo9KbNCu9UM3d0KH6le87tNMlIbBJgEvTpTW
eU5tCZI1LJaFLwkR7NaZiCA0wWY9db1alS32LPzxtFCUebemXZcRhtRFH6ZJD+bSVXFwqyuPFvTC
JVxntI78HZTCChqEkEeVVR/zqHKw63ginzMpyPxQXaXraEk6BZd+MIvHWltQcZ1xai6bVeOhIwUT
Wi3tG0nrv5gecY0myGyYCaax/taZ555TW/Kby1qRbWpmfjjOfFXaT+4nLfANdWwOt5GSCkc5CEO0
fp/4RUlaIT7kwJ18YYDUaqnSchkqFJz9X7B2v3hviPS3Jbs121QUf1Jh2n4CiwNr0FYU0iPqDaSk
b9eGtYpk5Thf1bq3f6+Gq0l4Ud/VLZnCfNkFun+CGMR4GISc5iti33lJCSZJcpFUI+UmKDUXzebJ
kkVILy36J8QYZ15J/nUbONb+UkQLyTSJRkFoEmMXVT0TpChO8V/35ZQXhL5OPKzazCKgPql0wN6n
G3UuyyfHFN6x/ZrtDGqNiuVgmK8nro3675xMtht7Sc5vyNx6A95ngBQPG5WwGGJZwzeJ3NxhxFsF
ymZx57Rq0RU7B2fkD3XhYh+2Zq7gVWvxxqpI3zcjLuhDTmx9VgXJ1fudnzqftpWqK9U+H/8qjhVW
mPnMH6h+KB6PIxUVZX5vfktyatTkncLizB1B2lNVq9VVZ3MKtym9N0Jdxr+/d5nopxcmb1Os6skL
jDFmL7r60oatVKtLra39EehuuOZZM3A50qdmacS8AipTOq2RXURFIP6HubWe6POSTnunI35c71k4
WdZ7GPzoU8kjE0+5alGpeZMwpjF2Prw/X7yp7L7GAwc886nttcdimoJHD8dRHU31SXAomFyaCGg7
Ph9fnkRWICAx4gVHqvEM/LkRUb15wHZG5JCLTc9FmFcOE5pIU80JHmLkR6WQg/38USp8UZr3aZTv
9YFUPeK7ry/2Q7ZAMp2GtuEKdP7wRQ3uEXxELlhzHy85+Y48/7VdgqPYA2IPWFY1uc6PT/TgdkKh
bitOjrFiI0zE0xo2lLbl0ABWxEDLxTK/D9y6tiSVsTpFl3BXYdSS/NVPFkbNZ7KX2xC9/vjhN1Bk
IHoe1piJDvm/asbFo5Ny+1An8i5lFURda9QwH07QtlIMiu7ssxE/W9Z/ag2nnA+cbwFv++RDetQh
QOWJvTvw910+BvBz8pCKvzjy5c405/0/dqTYf8CQUD2bIbkArexOqZTELnQPcIylhVWYdjlL3Gol
T4eDn0rU3M6r8tVteeHa3kMQ8cSHitO5vtTvUPED7BrUcHY1u2xqmJSnUYifV8AkxYSxEmym0gIJ
7WXdmLe1qTnfqRPP37lmFMRFG9JIqDp5kyGNubYqjmJ2ny/lKWVKUlTQw5tGK9q1RWZwGvryjkpX
ET3DXzB3gEXGQBKOjhv02jrVgqdITAPg5YKPQ+Pc+sh7GmHDAH3fKxhO0wR406TLlP5MhZKufZuD
oM7/vY4lxOYkbEnbUNUIInQUafxGjDsotQ79JX1BbSbW1Yqx/iMcaWBDaBdPE9dZmAbEZfVt4pwF
DMTAnVcMG8+Y7ba60c6KWIXF6fox6UB2W9f3aUaQ/wKP3QsykX8juoCoB60Uz00Nnl5UCrnyVmW+
zA/MgJ+Dui1NW+m1fo0HMM8VErusgNSv+NmvFc/aOG2rH8qvDDMoCTHXQlu25gAdlwze4AalJkkn
HfbPTCJm9trF2NbKWcIlKme7WkaKgXg0T7Fs0RhIY0hZTOtF7mYEfGinJ9TYOAdyJ71ndi/M0AQ1
DCy6gbuqoHdRh7ZBewGY+WJTTTuJRrHrMZibYnoGwh0b9+DPjzsWj8XqW7004AcNAOOe5slTo6Ra
b/fR0cwiB9CbL3PCtjryoiOHWv5foNES/TipWbSjH6Mh3/Gch3SQUgtVnQSZbyK3Ak6mabupEdB0
kHQxhV+uNcqUwQ6SHoCMxMjVsOruINTPFBoMT8DhkxRBdyLivOdPOk8j1d6OIw2jCgR3FBtWHgjx
KH6WTdCck0mLSMUsCHF161pXSRMwpP563KpvqD/J6IhLhb8NrFwufFroX3zFehqsrO0DvdlLDL/d
O3ek3u7xKR9NwfPfEeTwXSWmvphDb/5icFtZtHHOZrEezs7M43o2DwnMfdzkqd7R2YYbYRlOhsnj
HK/oaxyBNZRzwon7/PAhkgsHGZxhw5zbmrff8CFT2VNw4uDnw6WI+TOoIOThtcrsuo2f9H/Ar/YU
+H5a4K62fnk4D/Gaxf2qdbkXrKChTLpK3J52fIuO1ZKJS84fvMuYXlR66gLRgdL/2dG4pf1ojyJz
yCzrTiTo03Zm5jJymrdK7W5bYQ2Q+p9vDBRLZw+DkizRMzboQ7aBk1BMqGDjIMb81K4u7LGk7UIj
q7hbqlIVcEF7qxWmWkE51xf2sjR8gts1R2jmZjR/tkLfu5a41F/nNL/arc3HicLPoE3sr4sGHNAb
6xfrc1OpWYTMN0JFmwIxQNlaKNp4ZLOsJqs7EQcQBMJ6fDge1HZkEKMgRNU3GlLcGFoBC9V1cADA
CZYZFCkP27TV3maXlAHfEppzeSX0AuURALh2sMPngYnOVvKmcQNdsWs7P2Q6vVnAk+t33QV/WxfA
58P8SD1lXuovGMtO1c5iV66By54tz65H06rETESMMX7MqtkbwO6oiG7j0fX7p6D1psF/kXJO/YWG
oTghc/auwKvUGEelSwXLDhIdNfkIjdpwAaK+SP26mkZLPSqw3YJzZc1EZZhx6Jv/2RmneRC0GVyG
uqA/JmrxOV9t3uqiAaH8Y0+lQA3o/lmmU7thA5WawD3YbWcC2wbxD0ybczDPPDxi/sRHJLv+imTQ
ivlrqus5LNaIvxzaL7azCW3RrPG+CiwSJ6cBbQcx10fpEvTqw1PPA6AgNWSkipMNbxQ1J4JnCqr9
CLDivxY8OTmaWX8qEV6Mi+YrGqJ0DlIVgYc/2oM5vubV0CBqV0wWFpgOX+0iq70dqovj2u7Fq97t
YGmFtCU8HUNDxOAPCQ0HxI97igrJeooliHGNDnUPBkHH9o26LQSeV4XDl7cuSUaSzDnV5FZI/Vsi
8jYIRTS5w6MSaE6N8/hcS0v3BnUgwUikHe4GnBJjCTjVJT33l6Yr5G9o7f5ZSWt4issCXsmLit5t
t6MJ3VtIC13e4zLvL1te6lz7VMGtzr0M+bSE0dyBst4hUW9wrKClmqor7ZZLO1p87Dv03Fz42Gc1
cmICfGTGW0MKygKEh1LaU54CG81QkVA+xMJlkX84yq8rtUxbyTOc8e5GjIF9XkCbopadH2Wyx646
to40oyNXl4zEdZ66mplsyuKlYR+MPfwlYrDfD6vYwSXgB7JRaTGC6MrTkCIqnqoskmO1WN2tenxn
FFObuV/aeQY1488AK51gt7iqkKoSd5R0kjCd8Z2tCvSbpI1BVeygjBssS1LlSI8k7Y5GX/rzliLP
SIfjKC5nwAt+DiW/sUhrSnpX3SOJAOVX9RWNWA1ja3xxC4nmQVr7z5bzSPvpTNiioNRIjWvnIWxp
mKmzzH6qysPCGMH3NgtnMIwuxO119u9fZiIoYsVZrxY2dt03zHhecyNaXlIHIPMTTIWXwg9A7jb7
9zCT4PjhkqcJLtfJ10JsGChYh/r090B3hLaNZ0zur7XLRK4eLDJRtnFcQtThSejyjdrm0pWRX7Jt
Kgc8XjZZLyR4gDjMPtc/kHdAW3kT+tiLp5itG1BM63uNFiPSFV6Nd+Vbdk0Fhh7pe1Xwc0tM1FFb
GAhg0ygYpzK5GBwDtxgetmfcyXZqA/Gtf0tJO/5gfpiHzlMuRIf9fTZP0Mj/T1A0eJn+b+DBJ7BM
yURLI3K5taLfHWwNfK9jh+KLciomTVDoINB5BGcNKY4jZDsULuN1SLpHSqvhupv84ORDPrisji2L
FOKCzpfkF8XcXucqlGELz/UpoG+bQwpxh07YcYn6/i2Lod6MZGlpRHg36humzEX71uVqjpb7bBk3
c8acOsWVnhUIHm9MtRWiq0d1kyMRKVuOVxyqYL9y7Syt3wtseCh2xeYO2KVKR/g3nsvN+H+FynGy
1Jv+lBTFOSdP1bRFeI5KU6RksfOV2taiHOHe7d++P9Fzm2EUiQ5CXhqbmFWA8nVI4o49GtmLAMsx
lhSi1lYwIYqPDiYIrnh1jiIe9jK+Ll357dkqFHEc90GlKX0jSWBTlUMU7Yfj9XarE+L4kUfXjhki
3SiW0eXJAfPO83zdtQ/H9zboR7LHFOxxuoy/bBFjAl5feE4keoDzf+2FO0SCFizzz0HRaXuhznzx
5GDrrjQ/lqUtdFzclGhSFVf1FTKzYp/ZknjPzcVjYYJDFsrdL2sYuWpH1T/Xz22bjkpzKV3fHdIB
MRB9FtSvUU6GidcrkLAIEpw3LnrI/voYD603YT3MkmPYqMuuDGEE9NtSmmGBhc+zNRuVFPGtiT06
6+Nh0xigFAbbNxBPAaLp8JgC3hA4B9ID7JXC1/McNCJN7PNq7U/Fkrqb/JNLOSwRAcBFDLWdOfrU
RPK5H6x0D3UeEO9OSB9QgDXpyXHjbcxjV/M/IwLnxawtjSe47TIASwNonGB8Gc4dtekIhjiOkG0D
88baafAvEII9a1ATMCZD+Q6ckUZZ2cknoUMeSbal2aFjWKa6WN2g4v4HTCSvHPw0fRkZZBy6QB/I
iUnHo8Tp1Ks184qCFF7gNLY5GMweHGO1BPijmp2h7/vgVPPodspvnpYpk+pnVwOkBwj9kiS6zDoD
KxQAILzDBXjZ/v37GpGfW6D68S8DImGMedf5uLZ2z22j7DOV6XUxxxJ5aPjYSSJjIx/C/OwqkL5W
IIAu764uyRy9DrA5MkI27XXa/PSoD22WMzFtpDUkGlPBiJ/hj/anzIhjEMAbDCoWUh+IHoK0ArGR
/91jPcTWNFwjAmRNlLA1whLzA8Yka7GWN+nXXNKkESMD7FDF05fmTY1pMQ0tPghbbBc80KrP7GAk
blgyhKT65ugZN/sP3y94bPapkSX+qEQc4BRV2SYXwudJdlFvO1UIx0UGq88VjgdPHfhABvmb/ETo
h/v5AxfmCWEsk9S1zRx5FmtsaPFA3f+zTl/aKiENYqSJat04QrTeKtUm7qJBhcDUwIn7fN3i1AdO
Rhsx0suCAvyEICm16/0MiWzEKhI2H2a5xiKktbYaeaxE7NX09ImP1QfhQBlxr7J3iFn2Y4+q5tyx
/lyeWwVE8yfzT4tw7IDWm+iTAyHY5zVeIBqbo8bK/yyVmcht8PL0GQ4mGMGRtvb2n5qBfStLD/yV
FP2mwpAI9AO1HXGwYX6Mw0EVa/QakaELooZ5YUhLASCNFy/XZhMCAtLmq1MVL+yGLy5+m3XjqAcz
eXhOVOvnD3YqSXkQWqWf9/Hfh67mLZ5ry9hZeon2wXq8JEHKT962+UeoyS9ViYa4V+qKzBI2sue2
cjzAEW1KKg5101ebsrMDu5RIf964KVkDUlcAM+UaV+kO/Jdbf9MiMfWyl/9j21nC4cGxyRTxVM4s
Wkop9QobeLlf3CqBItsfFbr3wPJmai6Zf/oPbvh2S9PfAx+lFatgfjImbMJKlJtXZhVi0JgfLSwd
WDYqRuHHVeRJs7zOcBa2F8MBISX8b6TKJpJuyimPDdGdbbV9NgfXjIyQhKfLgYCPHpn1uHDTwsaG
MKoUvOpGduspRXgTBSfoSx4So0wko3lJHKmD5MeUD+JFZpdvw08xv9+sOtgQHqWLF4pCDZYgaPId
59AT/2FfeZ9PC9XHW0aL/qrEWlG3NiewUxftuMV/VyIskcZnqnZFEkvpfui2eC42oJxRSrQrKAm3
xaZe7D4EhuDQRO3YVsvT98p/nleOJJEhIwW9tKHoL+Jn5fTRqP5lK4Za9FFsvAPE7zbO7fabHhng
o0xLHv+qeY/4BuOe38hqe5vxws1VXxicwaKwdu7LD+KgAciqD+Q2TFk3uL7AyEelhJZ4hOzPoE2g
Z533/eU9KwmRWQXL3vji2zIcdbhu99/fK2cWFzLqRqIwOV2ZN8H62Xn3lJSkEjVZJCrVsX+E6EZJ
a+nHs8jqiQQ/Ow2P/zTsjvO/aNT+kbOaCRQdMDzi3c9lwjfKqUSNG8HTA3/TyuWOBjlGNoiLdLqX
2pQqqAASzAcCP4AdsRg+NOh29sXZuqDhwuSQ2Qc2b2XXh9/8Agq7t5KgZY2vzf0eXefcv+ijSTli
A4R7p3+70qBR3nd8KPZ/VYRTcbOH8Tqbwj13XQQV4DJDAn/Q8fUMm8Z0/I1Zoz1hZ2QSIxAInaEE
aejeLAOmkNctQpcBz3AAdLdhReotk1Iw0hSgPdW4ji4+lbim8q+FJmjWf1R2YbYznErFIb1/lvBc
wwgRSRQQS3tNb05XQiSUK0gIMbpF0BCzyb5uzgqO6a9RVwwbzVVjgbQrp1URDnkcjCSSipvSmhWd
2pQKRZDoHIk5P5G9foBf6GfCsG2XWmQ/vuc//oGp46hyYPRWP5Zq+6aSVHyAg5BNZWc+lNB7Hbam
VtmB7GDaD5kJ78nUHS7+LbEnSblTFRSJn8KghLCE9/4pXVSOnk/KYBQasbv56psYpFv3UFeRPjZT
cLGKPQ7hMt2VUtiu9u1xX78Lzgo5bMPr0UioM7MxBwFfsjRUZIpSt8IrSiXAGKfZSxrO4sNT7XAj
omWpwYzSRleaXIxkRvxj4TCVCTQkKtypinw8eEKvS6nX8ATuSmjV57SJoasYk/iLZM0gJ0wM6oNT
dNKZsgYSeGE5KmBpA+79UwWbDUlRM0zxbT3nEAwm/Qdpxy7BoNcyntvdDShJkySOPVoJd8NgjKXu
L4j9eWCasODiJslvHfH2TOvD5QGnDa4LrYGDOZeLMWlRclXgVlvQQHxeNrGJf7jgl0Ip387jaVvc
g9wTMahikmFXK9uQScn9ebw9jSh6pYT5Cdrt/oqQzux2W6s85Z8oXPRtbrmoLQc1mS8fCiwfTzRy
wJAyfRm653aqRAtD2TW2Oo7Ki/BzZix1mtIVhT0m2c+7zg0+PmW/Mwpj/m7l1l4t9SFnWJ6xaOyA
xuhkkEWkd98Z2uRFGt2xbwjK4teUvSvzlWVuDo/UwP2acQo2rIyR+7TxIlFmHl2GD46gN9zZxlxj
A8ii0HEP3HPJPrsygIGM3KEKNA81Z6K4l1RlEdbWYhoJ4+v3Dzd6VZi+SZCPRXb2jevwNDTWbmac
noTq5aMjG5/0L5EDX9V9YFUAQ8Ix+vGXUmjQrtOgUcbCaJidd3gu3yDyI1w7zYMhxPeV+AQ63JuF
d/lPgguYoEBGK5VYgFbFbSSdcSkmHHiit/bpmpFGa5IRQMo8sJszD7Eud/jkq/tFMQtgYX/yE9hg
dVShGo6F/QD0t0RXq7ULEH5cJ4Xg2WRAxTrmiP85wcLMeqJgzzSjLF+dcu0ROWsVU38Emk67ym8Q
jXcJ00IR2z0s7clGlbhSxBSDm1a4oNRCWUXZvmnmAdKaBWH4fet6p6da3YEJGbczgozySZERBcJN
p88rajg+Dd/b3sDl00hd0WX7WQWsQWkJPLxC/GWazFc77lk15J7DA2Ct4V8QcVnIhNdOvi+/47eV
F13Z1l3qCRCn78p4Vya2SLYIcYWN3G1Ma9mc8Kcv4nPvuG/OqFZktBQyMFE/deufgFUFseJFUyLM
cXrHEB0Rl2Bs7VCroFt0oMSiIqYjeixE+hvx7cX4jvHTP4veQ7Mx2Nj3IzDP0I/VVAdkqr6UJ1vR
To9Nq9NCYE+idulaLpqcQ1D8g74GZftWXFAaJDNTrhKrVaDRONl0r+AzueabtmNuEy2nTDHDQfwp
WN5lvPnyhI3EXpHYsW7QRT/U7IBEPTIA8baAHaaHJAmVbqnhAg3UeM9LKV0FFWdy29CZfzaOAkOg
GcEp9ChKI83wWenHCUcdq2ynLLUjdY3riSN8gdVNZBGlColPU7sIs8hqdPv04MOQsJRydUxDUrf0
eurkRDHC9DVVEvmLVWt5DZcXqieqeKirGK02mXraJNcY26M6F8xqBdxyI4vjEEePSBeRaz3U6/uS
byTQZy09KhK6tvBvNIzTUA18fUNYfAcBjVkB/4pnpkyKe5R1UbvzMZyEMZMeSWz8AlHMEkorn3s6
z1+y+phG4tiRSw2HFPjumkZbO7P1B8kriJ2/NrmoFCn/JlwX/wvxUxso7FYu5jgoGyGCf+I93SPt
OaFBF9xXrWaQiBDKVJLKbbz4cR81cFEyzqFdRwoeVe7UQ8UWof06WTHXrC5YVqmr2SVfkkNiSEXM
0j/xOvhNk+xwpEE0BSH+nqZYAtIPQxM9IRoTORUnSbSF7ybrzR8fmT83pefv07BuMkUEki5p6Dfq
F4eB5iBNoJFhYqu7sypmZZgpr4DWbzYnb9CF1g6DL8JpuN0Z14u+Aa/YmB7Ced9X9LN91s+XkjSE
XMhcLuYF8YO8W6tF+3lqnd+A/IOI/AvNtNDS5W6dRGJErAtrA2oZg2vxBIMgbJXXGRtnoEXFbKZq
Gj3OgBzeA6kKr7RcAsAVFWSMFjDg4djgxRTKArBjPKxg5viDX/rNQqV/XajEtcXb56uB+MWZ9/tp
OS5gYmQUBkkZuhRYFFgT9obwhjbQXwPJ+urOJHAunUHOs7eB21ZyrMJ3tKmWrIhfh1gjxUQlTEzy
TODhzJ03cCzopQ/CKQXuKDh+XHTqR1ethv3MQbqBi5GE0EF/80LHJU3w35oTnI3m5eP3R1lMnOhO
6tEG1MNlkFbfDc6RsYOyy0ECXwMLCCYHEsWTpJKauaJZVJC7TEFnvE8oL1zKQJluZmBHvs50TLpf
WN1QBwWzANhyxIIDI0+rh3kUe0F/dsWyQdRWxoA6hXDJbTO2zD+nFnDLuNbwcMIhpVEEeB1ILWEL
XKicH+Em1b2t4j8vGLF3fTV+NLSnEkgI3TtoProIu9ysl36+IuIMxkG/VWLTfmQNZ4UXQQhQipFL
T2YNvK5GIFdiYtI1Mm3lPS3hC7WmjXk90Wug1OYwsGNItpQPvYWkGh4DKMGnEdNYP9jdiqrr/3dP
K0JOJFkZoGX3CAUHBRVEqMgBsiRuhYu8PJ54xcwAFiQLY7yrdP8Y53W55zOlDVdWIxndijU/fvaP
li6dOfvf9fjx77XVVBXGpbJvHMkpVQ4W7xqgCJf9Hcq+V8Ul+F9PluPl6nfyBuY6XukfZGZ9osmz
pdljUVEjiDSsIqLM+N3gDjqLqUooEPkj2umZCIBw+AXweo8m13RqQT/RPj3Jv4bOdo43XcsIz8oa
nQurRdEtsLCUSUlIeA8jsevy716yz3DHhAWB0agxizs4o/Kv8YmEouE8BW/v/A1VwHwjzboQeu2e
d9GY7eb0M+xwk6J0DYzy+2IR/faJdHodOz4mIi/i0MRTI+QtHA8eJ1Q9ReLG6ib+J2Azo273AJCx
x27VuG+XsxrYkwo0EEgxWgoZucJm28YAUuClk498ldPFzGqDM8g/2M5TqNUQ5Jmh/UGAmhda5og2
f/Zb3dBVuIgNuYlU9HRP8in4h5//Cq5rDTj32fZmhhLO+n26c3weTY6NcOesiXXU8eBB9H6EB1+x
emYPa75wMe8+VnBRm9qTiGDmlHT5y9IaBG9kCuw3MarsJRbmKcMkHJQTRqMJWDCMXj8HvMJkXeza
MqoGECLPw/UawCheDOZ6FCXLsz3UHBV6e0EEqU961vEZhsOF86mf1Bbgj/kwq4jz3mWz021XVTPy
48zJabU1Qj7WOEZmMxKwsVDPfSbS5ecZsdina2Ry3YFS44uDYdYHsChS8wpvP1hmQSR2bM6WNJLp
UJEF8Kfu6QfhcBYXEk60WlTlUyyVGwt8ogbZdT+oQxMH1Udtca6wYzZCATZ6sgB5rf16j+6C7F7p
RdvoYPOdrCJVNz8AdBKFyOWNpV2lJw1ZKAFENzWBfcZA4WGI5QIKXV/erbBxBTwb1Se7wvhpuOxf
zwetDZikryk85vIrOmGTsKD0UZYa8zf+fu4YRwVhSTXmq6zM8CoU+w7v90DrOJLhpVId59ODY9+w
zFx6Yg9qY2GLWQfSJyBdtylOwzj6OfpCtBkP81nhrtTiweuPWtV4heHSpgR+lGOtdIsKpaH4oziZ
SMtRv3QMRCKfGbUu2G2ysMUqxFsm6EtLSeE8/EWqzdQjQM9r2tP1Ay7FONgD32hOdCcViEFLZ5MW
qC/vnXniwz+Dcuua+mYYWgWuXE5O3y1rFL6TEVC58rfcnSXRMW1niTmi5lG+X2U0vKNTpJqOw8IE
tVd/AT16Be9vZQeLwawmjWFdUH26CCKuRVjHms5xSeoUyCyhLKiaPTAODmnlWFyOr2FB4uPpM4sP
PO8BLWxv9L9IcItm2XxneXh1REBxNlQneKcJeObdwbblNe7PMJHVnd05ErO5M7iiztOLFDBVtJV4
7ZDWRsoVGr5VDC8g75cxjR1dmKd4QIKTkVpZ/EMj4h36BI1r6cjADbDHSq0greaGDRhvlLd9L4aY
AELE39Wp1LLJz2dsSVWpFOM1GeNegSe3vdPIhBT+B0SVV054yBtErdvr+j7ZY9H39wsCaFGhHeRk
g8Ipil4xNRhf2tW07Z4UjsrKGRXNP/TuSEd++pHm712mjGsLNW2iRM7ThFxlbFYnJQAV6bTd94lH
89okHn62++wEgsfZi9pFEKZkcX3s1MseGjxirIqZIX/hE141CUM55dPrti4yWrnlwVWAfqrU6ujy
Gq7L5UB0o2ft/DR4Y/YGbOnOWcTZXFytQEXhKLdyVF06eEe6vg/l/PiBIqDOoexYUw93BbM+HOTv
vISshpfCjusBrN3uVQ7+ZO4mvXEKA84TzCpAhUET5xhMI9bIsY2ftRHT53U4VhobU67TiBeahS9u
Ttxt+A6xcJzwuGqgYxMAJ4uBdtCPiHklJ0zTF34OAYFmO01knifF8xMCF4532fZysr4IsbFn6vZz
hx+VzOH2/bDQOwbQm5XGx1B8Tw5ylqy3lW1vRJRcRJmRy8b00OYV/SFncKRNmUyXi6NS6MDu5CJL
+h/2laknCDx6vtkG27U58DM2vd2kxl5PJwW30hOvVYTMU+kcKdXo8I5BI+OERWo6o12xxUTWjgon
M71yTLmP92PoNtrm72GQ1qrPylcYSJlZs03xS8FWYyaMBjXANrwwGRolka0ZJuebin67v9BtBMRk
G6uFVDhJ6oz18cycrroC6ie+h9LT3IS1HttI7m8HV4TMBoKJ/bqoiDEreKbTeWFq6qInueu04E1j
3bkEKGSNoR0yD1+YQ2wTed0qXB7n7tOHYWz0VSYyL5/m2PZBLgOTR5LgGNoZOBR6KztEfl9pz13w
q3yfvvuiqPGzO4MRhXYZkuXEhDhOvysr8JQPRE3hyI0LIZp5EcFTodOfgIC1uQxx1nK1vBVTfsuC
DYWpJTgTwwy3Kq05z4+n1Ht9IKyM9IHUgftbVhpHKyqADb0YY0TRKihn/UQUjnndx3uXVtQjCiI0
qL2yiOvWfkBWf9yjvLCDvL70MpqciRyB9HlJAur1z6suPYNioWYbqjJa2KNHDXbylz7vKzhJCzFJ
3YLZh/2ubzat4GOIw8zYOekO+2NK6p2vc655TeXNY5tMbWqoHJzq0AgFwhdEZJwQUkVDeAVqDSGS
o6BAFxcQS4WRnYiKhB64VcIDEM8z6JSqYsySzaEdMWTkjHt5d6NxlrPbqL0jIAoFK5Jwn2JhCXH0
+gQ6uQb6QdPUHzwHIhQs3m1JlwtMkYa+avhU87P2RQa/xcEAF3NEj4tLuA3Bem+QDDM2iJCleV2B
A6o6Pch+H7pEcaDI+LrZ0xjqdRWWWCU9zIHJdAU1Qz4ajQqolhENxVeSt+MB2iM1+V1s28JqwXXH
wh6c9YzUR7/kInVEem7BDaSyiu8kSk6eA6I//eonKKasrXw8FrWA3hiG/IgrxjxglcO9y/swKcEE
DmVE55lSnukfyR1Uem82Z8gXIspNJc6kawy/CfDGaa3PC0mdogldlauPKmWNbZ12VOu4H4DMvjFs
YbNpbknM39ZPcCO7OWonCLZio6yf2HjeYc4U3A/URYgXlJ0SFHm9KppiayfBPYBfaDiziz/niP38
RGfDqHOY0+F5Sgnd/IuFytKyHg+Bh7hCxCFZR7JNrxMlny1axQ7JtwNwaa4K4QY6bliWClTAWyoK
QFEMADzjjwtay/tUcXpKpqhzJvjEe7pEZ7m4oqOVa0Pc8Z9zbfolyUZhV4Yv8bE6b5UO9BM+/o1m
InmyLPPFPG4ueCS8MARkkEAzkJDhR/E6M3yRF8HZg7+wbv9PwYGOzAM/YJgTmcoJUhkgCDQVFLRY
uIW7Okj7fItbNnSMFH2VgiVgL72ga2XpLxekgrdUW770qTsvIwKTNBlWbsurgdywxJA9Igdyg77U
jyRiWAOQrI36RfwqOVvExQjLzZYeiQAJKs+uL2BInG2rk6wwMwp1zLLBLnyAtHn0yK+H4e2K3uMA
WUGIvyXPEavHqlPTUCS8VaIZ9S35ZlO4Asek8crQ5cGd96rpOM4uhb/KKwZLS9Az33UqO58yq1xN
90Yf1bWW8cS/MtNwkU8z5dsHA9DVbXoxaj7aKfkTuRhDr8TEm4OKfp4cK8adhv3eJB7t2jFuLUeu
Y4c+1G63SxyvcgXU3adIhychm+ZEQYt/o56yNBN1k7ZQXXoUu8dB1t6atjgKc0uJUIGlyV+QHRWJ
b2GI/mpull93LMrageSkAO+uYD6pbPewem9ZSGpbS2JnJYYKd961IVungNnDBltZ3DU1oo9VZ+QB
OH8+uNjcgUkbtcYn+FICb5p+jOZV+9LsiAzdujsCZFBhgZwFi1FozKZby+vCBlRDdWxmDcpSxgi4
BZ/l6Tj8BPZhLd5vdEjo52swlk1QHQQGBF1x1lBdk2ut1+3sgd5uBlr0MjqarjiYGeW6d367ot2v
NqwTVNsX+ZRl8ttMJKKTGJ1/78PaEjqhLb4spKmmfaXYGAoMTJGTzGAZHbrF3uxnVl8agB4EbPOP
mtmyoEIYmPSWdx8FEGWFe4Ke38Lt5JLbX0wo5v36v+0Q0JgSqcJdn9WG7hMsFmPS+XfmE3ivezXj
pxWLYBJdXrQha38/7TD5NVyVg7eM4mQsl/zHMlX0tAJaDZHiUQE7r4GaZL5MApjye1QAuZXnmBeX
0u3Spq3mD363snUozFzn0Ldk5+WDrmYYmWVgJwgnLCJ7mxg3QzYD7W0ymrCzjSegIuj1S5vqVJjs
s2U/ybHh6VgNIxerb8KBTWkfvDw6Z7mvrey/1hgxYRE2Bvsj/DeMLiJQ3OjWRLMS44UZ5HgkVKWL
nfHKQVfbQAEGyO9NmLP44x3kmRw4eBPGyEtIGtFZqMIp4pgNDtJ0Ay5JnzgIwkyn304ecnIIICN9
Dm5lZ40DAtAwHcF4BpVJFWIfN23+sXgtHdbS1CyfXJ356dQ+tTlfSl7+apcGoOVKUyqhvbBR5dnw
/QKklGKJEYXHFi/Lq6ldmI/M+7U44AqyYwOxTe4gQTVy97gOKVX5CaC4eLig8/HDIrpaJFAGL23F
N5VnliixgG816YQDTLid+tD9p9MQ0Co1yAg824q5lRbLWIc7mIZftxOiWVF1LK8CGqMAJXWk4hce
goq1sraR8Hr6f/9O7WDr+TT2WEpHhzNcquwRwBCFMoqRl6Oi5JMNBeOlEAITfu+ihUGpPZ17PcaV
P1rwCXQLLLPkA32N7IazHcwG3vcvQZolpNeTuDtP535ntiwVDHTojPxXB6RINNMA+JMjaMkNhQPu
uGfXiPq/f9eZ4RuhGEf4YFthtm/UTzzFclmeXJYqLv6OLs6mW4wsWm789Cq5qQfG3vSR+AYcMNLv
NyfCHIub5b8AX/UtOu16Mad1mq9xcHLk9ME6b+gEA3BxfPWTZVM17NMstUyfnXgatM2C4l61dR9J
OnWnzLwucS5ZYifZOuWIuckOZzkjwS0ZlCn2Ma54UPD6O59vM+mxnbd+6Tqf
`protect end_protected
