`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
BOb04KJRoJudBEfc67qBMx8FwmTzerWgH+0+uj4+2TC+LGlzLcQRUB0OXt7HbNZ2n4IUxox2e6jq
ucRLREBvNg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
lH0gRqNvaFU1Qe0mme5jG2jtlvHn6qO4YSynPKrvVlR9oq4NdF1HapDzWTPaC+4q5CIpkGDp9CM1
HHNxNi2QTxqO4QuK6GOtgbVHEiYkuqfnd+cTvrfZOQigvUD/qqL4+rzteP+3gjv6AlmUjPQCBpjt
F+ZXXtA44cq7Wff9sgE=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
B5e8yQ/VR5u3iQcjQZqSUpATM18U2VkWBwbq7LdjY4b3/OzvG3xZcbckB2JS1rW1vweOxNbEaCPY
/Jizoi4EmRy1UyiGAZm2AdRSIwYTGrqS+BdnHvhdDLVMW6P5zah/3vCtv6BvIvNMk10rOTAPe8zB
BsXnzSnqvM3+ibDibNW6wyeDDYu53k9/jWCT2J1P7zk5B7517VkxLySq2BK31ccfA6Ac1yZglQFx
RXWpcxHS3We+LkV3c1i9zOrWwXQj7xZr2KGIBYwu03dXG5iUPr8PioYW1f8hHL7wHIZgqtI/IHZn
qv9my9/bGlR80tl/wbqa/3huS/nR9s4EqisgZA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ao/M3SPLH1bCKHknOdawe9XRFnMpNLWuIi5eGNbohGBxefMLSC1YnCgv3r/UqBqbOUTHi6qlZ0oN
zm10tq5HBMwJQYY99BEL9DBde0ZDFQ9i8rSmvWKBioJnj274Cl6O5LMcnBxfdZrJ5sCA6TvE8jC1
KH5ch5ogHkyyXH0i1Fg=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Z4xJBBQDsflv3TritnbaHiNUw8gbGWc44bYVBY2l4Q602T/JkeZY6h9rBijq+CRkyKxBOfnF7TOx
Kz3fUVVh8vmFixf0mO/lsLDjY6yAndkdro7d1XdlsYR0nYk40gBpto/KRxYYoiP0Ns1oqPDG1Xfy
L7PMmN77S2D6PtixwKs5nbWJR1IY9/kj/P+NqJ29uAgMOofsgEwRmJne1g0dTTi6fYSlxfwXpWpF
SruF0Fy1f8mmNWyi6m32HosjVmW/gUbljtMQOIBzIjoEMR0Mm4MYgrbjhotdc8d+zbOoQAjuE+b7
EsgEcTuSJlOh+vBbfOvctIZwhq1IIRqlnXLp7A==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JfOmnB7OrPsYkjrR2D4DpqJsTszKORckIVUffs8tEkV5t+uIBh2gbrFyPGCo3dq9R3U65vQ71EDE
AxBRVk8H0eUOiu1iwM9AALMz8Eyvg3LPW8YUG0cHC8hcp0jq0N2bGiLSK5OIhNx3KCOoDCXNFRss
v+bbip4xlA1u1CqcbnX4DjX7nkRu4IbdW1wko74lHhvA96qox7nNT05xFD7Izk9VAbLixY655gBQ
dX3Cj5lrzn/YmrtITOxzS+aP/bgCi3wgdsm9YMHzewos5vWCyqGX9tkGocRxBaXMiNGsIxa+Ruy7
N3zc6Lutjhag81i1aI+q7z0qca0LucLZxHIrJA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 52272)
`protect data_block
SKPZOyLOb7zPzwQIaDX5TjA6CjFq3jsIs+L4CEokKVDpzftLdpdFUFayEvY1Sc5zbGzaKZNkjB37
IDYIGQaVpyujR/LEUNmefCfmM6EBBkD6+2YrZIQFy6h1l5oU54UGz4E8FTxIyh+1hkZuX1JbmEt/
C40M8TVxufb7ytsKShKWicavt+VZKBHxct5wrzDE65u5gGoro/WDjRNXER92Qid2lamb5nwG2A0W
HuKInGq6qNQn/vIiG2B+ifbKbEg/GS4Of9g9qrroA2bxqQ9iAYh5BuE4x45zHyk+TRJqPgXOQ2/h
bV2YTinJF+/CStgg3MJnXoy/xF+1Sx8+9iKfUaWLROf8XFax8mdNEs29JHAIqQ+R51ywgMPHW/eU
H/+YAEQ0f/GKhxgS7Yz+R315n9LKl8eZZp334jVHIjpW1dJYJwS+fPdbpHRRBIf8CDU3Xqo9OcmS
Tt7tznwdYwsp8hF91h1ou1Se4vRveOBfd1F4vQLSch/PdEusksyBvtmObh9QjDC1F4SBNTFpYS+l
FZB9U6yF3HhYzPrdQl5WF0jzVEZDEtTWHwbYCdRkoXp0X4PXpEtdrzUTeDisPQ0DgUtZb0Mh3lMS
U5P75ETMV5qZahROPCrcKKs1utg0tmVqlPwqm3BvZBlmgEyeGRhzUKCWAdkt/1N49W7QMZX28MBr
BmRjlak4NLgCeuOeVAyqVZWVE4vwwH7azvAGw2nFTEzgMgQYJXSD470dmMswMk/JwGkv/xeNalpm
w98kkhdDia783DErRIWVFDLANdrsteNztBngEeOAcLN2vS9v3KKXhrYkSyAn/cprqemPZicnzcKo
nbQ+qjif04+ccQPl4Tm3Zr3aWVDGWLpFOsPGrpnQ2X1FgVPWIorFQ5KNs1R/lIxMDUf4Pg2eXzia
2B8fyhldN2Lb0u+qkcx7p2dD4JhIZjx60RGLbLUxKLgvzXEbmor32Rjx3TioBaeHZ5SgHNk9QTNB
xtGY6FQ0mVpwl5RmPVfYJutdveFK8427/AIvCGgAPiMNdnv6uzJTH1AKxf2QgQ3RXO52Rj1aNNeI
Sy3rJtZdXD/vcKQ9q4hpD+2meQj3dB0i0+i6VdKy617USE7KhpGVWJYCmFmMck7Ds6F2kLSphFEo
NN1MNn0w4PlnOvUMSQveKbwCIHlePlm78KvbYwDgQYo2DuTa83BHjMrVAMcOSWP5kMN5u9j33s0g
nKYnHkhHgDNBxP/c4Ep8/KCna3xLd1TCCPP3eVfKJMW1TBlQH744fIKohFCWxz5/6YDJzocDVSB8
DiZ8JmpJ4d79Fa3TEJe+Cd/FPlA+W+fB0J+nvRS/V56MZFA1nuIhihhwSgjNRLJGAgGOT7Na1yIU
GxfKKEvjEsRqRPcr1J5UWz4mmA2MeUjp62cAR3kcu6VQ2K+w+CboIN0cRNeTYMYkXcfLeacqLGan
0LBdY/e/KTFWBPHeITnyjurMqHsGRec+s6KzFCbQ4ryYm41UJqiFToTcv149fbjkPARyL8XVhKBP
KJrXMGP3FzZiDIP418JygVLddk5A/hByBNuOiuuajMA9CUZ9qpY+hqjFo99woBiClJP6Xq0kPYiD
2puGf3Xo1xVdKSgzHEGw8lTSbkSdKlMqSKx2q6dTfqCjoEjz4Hsd/3LxXJ7H/Marqe3fMscF/bUz
fhB1Yl5PhVPcmjPwXx+nzJ6xIXxyZa4MOSnaO5ym8yK6iuS47mc7YRgTBw8rSU+ONKA6IEcbqz5F
1cDGk/s8mmycBl0pk6oAXzYuD2YPUS6KOSxnfeTzVLZNHMGqNi3n/ZLiZTJHD9qi9DOwEIt3RWnI
/XSuYp91gmEc8T5Ce0btmAS8I5BCtjtSvvxc8J5/5Zf6i+bQfAgTJOOusnR5B6lNPbcHW4Uttyyt
2COirWs7oe9Qz/5BJYOb9DMN9B5WUEVNDbAx/DUo/TMLVBzWgRVUIgCUrSf3gq533KVXAQK5aYmr
37eDuPqK7mQKn6E4YY95irF9D594u43SRyo+vcEpHKuahM7tYCz+MaJfjvnPTRrnfp8zOxPDmDvD
BewvqwODcXacFK3oMOIkAdWWxY1Y3BXRJZ5Mt5nYfbfjGAX0UUYWcjdhTA351NJ0SyqItGqly87B
TOAs+K8EBhnt1UpuiiQyKCAb/uQoNrBGK/PSL4EqW5tJP2tHhRPPu9KeHVZKk4gAdG8v3YqepU4N
zfnrydUAW8McrMy2h2TYOxg6B1/8V/SnChJ5NStk5w4ZkTnnlpf9KFP3Oh3YOzRO8Hn62QbCLK4e
iMBoOq1CADxjq1FdQ+c3fQj3yDOtwz1J66YpA5gzIs4u7VRJvvy4VhQYviEfDcWUhtqnahdt7xn/
YoawK46hAUOwobiYkGPa0SnUj6IJ2QFft9FiZo2JBSaPvXQumXJurimZUPkd2rcx5kbiF+eop1b8
6/rK+P2OrLgWx2FafXnJNcltGk99cXA72YogNQGgtQI/B9j67u98JFOY66+tSB3NLQgkpEhZZSgb
TWwdFM8b+JOuHQas+3BYQM/AckSooCM7wWyWaVbtOG+yWb4fsn4XFmOp87dh/+3kysWvaAQHLgrp
3XTKyaFvZBa5N7s+1U22d7SV4GHJmiwsBvhDVu9Gv7Xl5LCoJbpsSAKynNenB4ywlYFVbzpk9N+s
HBF9zJ/rC80j9NFX1ehZsQVFZSHjTDWgNkN4iKezQEiQqEtr4HhIjp/oamKyZmmhepfAd2OBl7Lk
RDl8GgEpi3GOm7E4dp9IdgkM+8IvAt1VoAvEy9nVs4Hhy3kNBRppFBUxttRuO8nFLsdbiZ9oNm8g
eItRl+8zY9pkJUvcaeQ3NAXdrU2rTf2ZmGIhfDa/EhrJ746oyop/64tTF/+HsmEFBBB6YG0ewn2L
/vex5ERkmwuLya0BzgEREnvf7celJWtxSQ+DcPNPN1vF8ANkHUmDP7iYCycxRWNOpGNfqXF+0yLt
6vg80mWf7/5KUUhWvE/pkZcY45e3KSh1kYxfdX84Cs31v0dkFaZQFnGEqz+gZoHTpgwHIwQR1zke
kDDGRqv+VGE1ztbrfbvlmYjUA6+3Bu6Z3re3bshbVvV8911GNalkBSuiNuq8LRJPePLEe/QDHDUi
dw4IJzhQTG+jlkdBl1P3EPP5GoCf811we59ywna/cxrBpKVRvBAn59MY3gZOeBvo/XyGqim23Ram
nXkK5ajQ7G8MDM5Pp67TcuYoe8j0NAFxWeDvyl1X6Y3zZQRufuW9ODEsa3l8mbHQUeurlAgXuL19
xZixy3FJpUB35RkKIxwG/TuQN0/FtzJokdz72xHvOb0zZxfIV6FzOpaPpL5+/L5Aa3pf6gV4K7T4
EXxC1MSe7/dlnVFSz+25uMzckCdS7PbDoKQyYxVPglRlRvECIGj74nFDwJB/gaDPmzH93YV0eNDp
4ggN7umxxKY6BxEYUZywmDUUnfrIvXywBPlhRP8BrXKjP9hJGUjWjAamMVDwPRFBxZRmXAILgFZl
DJXcSQRkBLfb/AeXT7dHIJngkmfUhIPWAaT7c/aUzYaYmv2pxIKQfnUs7ihz089adzqAy7nRd6bt
mae+q5r19r9C98+c10XekaMGCurwFUkEFA/5frd/BPBv8psWZLoRrx+OJw3RqnYQ/nylnxSbS2SY
l3q5dFwwQ+0Q7zTGjVE5CzHu5UrwNoELax0nUkAsayDaR2LRGbj18wELDPAoChPnkT1o87vkVEf6
LCjuWXVGRNEPVPAHHoNwPDT6gPvEhoyTVc13UdPrDs1t5wbywzNzQ6Wz403lobFf4YwJzRYPKjDZ
t6MNAZ0wiuT5fBe1YehdCuA+fHA4KZLbB9xbuxuE+rp3strLRGBYpmotnl4wyAKbO07BAs3JhHBK
/rvyukgCZJMISVQkLHJaLzOCDlU1+QZPUmmCSN9tgR60cbkSvRebjf+vjcfXFaPdAo/WE2fDAo/D
KrWYK4c8dL4FcM4RbYIt8xnVP9ZzBZLY4Ki8E0sYlmgVze0V1RG+25x/sPN6oIfoSe/TWeFU14H+
lr6XKciy4vsbGmJ4r89Ehx56K/V1d54fqKz6QWYAOLr4/8FJZ3mYxktcPUEDFwuiYB9PnRLbbpl4
UUtCN98jKxR6gmkLAM9Xkjj86tbvzuKgmQ+PahVKnKvNcROMDes3gXvG6lUPOahyi+12ctx8GS+8
ykgdl+o1OtYrFcD9f1IJL3OAb9pxKwr24iUnKUH7J0V6drGcuM9MX131CPctjHdJtpFGd2QWG58y
U/DlB9YMkZjVlamBaSv8Ie1H+jOSusQxaRekoe2s20+/fmL2QnIgvTn0qBMD7/3PHx4h1eBIEYO3
iGVZVKm8bdEloufrRtaMeYOcUcDw8Ewp08B014YHQwJ6LMFzN2uvzhf0bqnxO75dSdnK+GugByJd
dzFRjLsuGqYhHdgL8bhyWqkpNkmKoRoR1AEH7Xjm0LXonCiiAWn4LOjKqOtMP6YmNQPuGHfInHjS
+mFhIxT0t84GDww6kgr5bfIL0WUDT70oK86WPk8TNDndPy7i7LhiDFK9SK11Xk6eNtWxpwPSdQSv
C8X2+mDW+t9P0FCeF4WMYXtQJJ+DVDXyQdmKu6TiFkSkeaXk+79tTsNhS2h4j1On6k6u8LDaUOdE
C3NDcy2XRVfWEikeusd6PmqwP0yKRNVaqcirLpOHoVVxgYRcb7dVTQoSuf+M8SaXsC13GFyxYCFB
tWRHcTkH4R4KG9jnCNznDakB5dc9yJhq+00wbTVX0rU8p2HfGkzmpbPIMqwID9YFTBrw7cFyyTAf
2gZWOo2Rfog7aUmjn9F3QpOvnqm+3VhjdTVwrSnfDuJm93El74xNvRS6HkobkFgmk6f2015QmMCw
Bk4k7nnCcMw0HPSKxzJXwLk4+2SlWy7GuugeFPMsNi6qa2oW3G1JLWBkdyhxLuPnroG/QrYSJWWK
hKXym59ld1cWvo4QHZC/jzKL5yVm9Pj/5pT0FxCV89awa5JbIJY5zolJJn/IV+YEDXYiZsbUrHDq
JftRD0Na9x0OchMAw81jouTlmCSRux5v8JiHYkOHlTrT+cqgbyI8rWv7Lf82vMfV0K+lbddbWYe3
t0gbvWPR0Nx3JfrqKB+yAlnrxBvcEF4unZYQZRu1pwZRSE9Bxdlg5hSewZSvlkluSSGlQ3QLHNq1
iYAraoVCEhO0rYezbxLudM5gLUo5w/Vy+NYfVnVeuOWCzC9Fnfr0+lZjXcJaNGBGG8Y9PSkPDg55
Jry3At+/pdluoMBMz3lMUscMRJ4eZIovbw8jBQfcPCwIjX2RQ1JRYRTgSe2MklRjxa/jKP2oKl3g
gmYolnkGwen67Njv3nkXPBV06TqBzscMOMxkJufiKR1JXhCkRKg0qE2wT73cHI4ix/H0xAJ8pS3E
/FhgIM84tzBpG303j7qVg/WLUlVStaWFtnTw47x0waf+8qTiYpH8/N4XR/v7XI8G0DxQeh8yL7EP
VACl03NRRm6NCthKZ0IkmCxLc9uSlzE8OakJafRfBPQ039RoiFsEfMNRSw6Zt0VqNcztXkpV/PPk
QVRGv2UF0D94jwEzxm5Hm1wxTThvziUBqzYG9ujQ5Y5mUCAZxbPiTJRhljoy0KDJmEzS2FhjSgUA
gmE2dgbIFS+a80hjBJo0fIe/3olZ/aXRGI4aNyLFdUlydsHnSos4qF7o4V0Ug6OCqotsJP9G4jvE
hi9e/xwkJn9FoemNUl0c+YbUdzIATrWz4K5trDqJigqE0ZDjDjZg4lkXbmBgj2QLJiJs8Ptbol/z
KBJUpf1DdGcoq7raq0H0N5eFl3zA4p2rCukgWScQKqZyRTWncDMqitgkhv0SnUjCx5keXvM3jyWJ
sol6eD0ovlsp/G+BN8ccLai1QR8g6weKDe+VJT7QplopwNCSarRwxHPRjsF8dHizAYYZmoZH1Ph4
djLL4V6HBaBh/ZgyToSW993VDuo8ZYTQdRzggOPxGVo8gaZ9159bsNAgRkZlqTLDPMyHsQjY/Yya
aD1U2xqjLdvgen4XuSVjNRKJ+IP+CmjZsGjL/o117tKLF1DfGHePNXqiEVFvfd2ljUwu/XySQJGt
ozyFdHDJa4tXFYz7gDWdOvQBYFLAZWhBv3EZWKWcP5a6dlBkEeWzHkA4yV5NhA4lFnqgTtIFqBXC
SJ9RKaRCWAB+TYmgwKKJl7pbL3yYlncMT3KSCEZ+Re92UuUmwlQ9lRqRtf9+GNYCFfU/mr73WAe2
LSlbgvGjntkZ13HsngeRZDicgeZm/9fV5Jl/7FvXXXOozKU/IT98AFLTNwhvpd+uFgCxYNnl/Pka
cUWFPP2PS1F/wT1TFKRVE4hdU0w/Dej3j21X7KzQ31TPH31srV+Krx5dWuPi/4Lwr3ij2u/2nMPh
uainaSEJ46p5EqYByRlMkoh4wU9GWrYryPV4MRDd2fPMgZpCrwj1wBru486nKWn2CXORag98H0QM
zfsjwUYn9nSz0OhaXUNL0dpROQoRN+u9WqsXpsXk/vyo4s6LbjlHT0jpEtPRAj8GK8xXPT+2cWl4
V/QOYqFIlhuc7QqbAsEpIA481cL2NCYQrZ/l47kewDR7TigCu3Ph+KgH78agVzYUfmPO1BeSKHCH
1SXnyX9xolbcV9DQOKjh8MQ0BQmrEVDVtsseKcsO45q5bQYWJCrItcaPf/LHl5+JbConX9ql0bxr
BQDJsNtvN6NBR+ggzCXyl21KwEf9p/FKPVIfS1+AXlkP04PqqZh8YN5NIQFADXSHvEyavU1LEqu+
oxlOVpku4Oh3kFqORagPg2EwGtyIdRT6F6c2h3C7HCmazQtAg9IlJR8Tr0Zcy+Nf0DfAl3O1b7XO
jQ9LvEKFAkS8ggt4CDhcDkeMjmDFgt45E3000BHa0/v/HnUmuG2XDC676QXxgIVP5Q5aRPgT7NSh
raImwTlZGhbS6EDTt3lvvXiBJvBOlem7D8bCfB19sQBlKnkNclN5lbJoix1fCpCGwyJqRLBC34cd
cN4zSeGuYpBiaGcHkHIWsmh1DBEIr65567kD/qD8x3tkeDVF/DnfWg67LgVomqet8XM4D8zlaxHe
Ku4LIgO+u0XLqcVGezdOwBCtDNZWyX4hUcN/J2qOrJF8qW22Rt7UKT6GncUqTe7ZseVyvlZmq6r6
dsfq4+QO3Q3XPu5cTw8Sd8re3pM1/KlxZ0AlAcZPyqTA8JjPl4BahxywTcFuP63voMNryBkccTgd
7P5+o5I87y0a4OhuoG5yRxb9Rs3o33aQWar6GioK5qi5FhvNgBF1FaZTR6w2s8rg990XSVsmpobO
nmr9nzwNXM6upVg4C5ESzOyZ1aWqA+JEiYTVyBsVBPX1ermgTW/fDA4kBBOrKXrQxhr1WZLpdVXu
EHFNn0a+MahQlCEWhAt3BKckfwYv9xSL1bp7KGPEvx8KqDYWVkIKA41AHCynVmWgLpdI/DhfKkGs
u/7tu/+d8NIAiMam3zA4lSaPK8tK3npLnMo0SqI4pmP5Tiz9l23MV+CUd7LwOS9LFIm7OXEi/G+a
nEJiiSf6SmmZXE0ZvQIrLrvP94v96UZAc52TvF9uYxxIM3YRVmI4INmMZ/L4hKY6MFahpveDGsHX
iYvNa7h/bavnVsshXfJOlPBGJD9UxVNAmBTXRl3YlfwFWTx2hLuzdD6kML4VOZmAzVwYCzuZQvjT
VQGC8O6lkPyFUFo01iptwjDm55HwRzv0TQjk0P7fr38N5rKINQimF68ScxrieFjyj+9YeLL9VCZI
P/ym98hge7vhIN69e1dtQQIJUIPzpTV13GEu9V45LAqhS5G9HHVitUJOWDlisFfiPyTQL0x7twVg
3fPIWl+EZB9MVF9o+cTJEsr7Dw0/kdqYW3bv8CNqQ21E3OUnIx7TNJoo5HitaTDLLHUR+xumt1V/
n8VfBq1BgKANo/aSqxm1MI6VWkdIWTwcA6ZNvJMRTv2NXSzp6j9O3fwAG4XwuO30E21fybfy16MP
3c0ts49bH6dgzG0masZJii1zterWNG3+jkzljsVKYsNqQKhSEfcpy6oRVrUElxTIymlHeRJ6rlWZ
ppDgZatwa04M9Fv21C67kgzTy73MeLeX4kVbpYwj8GBtEdnmW9oE6GUfGh2NpJ/Hld0x24YivTy5
Aa2X1Fj4eBm77Sp255T3YjIat3cXVq2XsKbjgETiHjQM5cO29jXOd7L73t8mWE2S5NBtsaFJWWWv
Fcj2A3IBlecU/aGViIdBLucowIDyIUpVCgSaehd+TreeoTjNTdoVdNlOzhEh1DYzY8kSLcJkFub7
1L/LnjKz1sN8VehwQM26kGDm99lXpHKJZsQhZuDolpo7IEYIWeYh0lBLJnfjQXp4NO9xyA5upX/t
rlNilxEbAJZIGA1gszzZ/5a47mJzlbIm9JHjSWn4Hr/NG6e3N16j8LzEMB+IO1sTQqOM3eOwdTev
eK0DLVfE0I8wB/hrYH6QS/jN66YS4jSawtyhRIw8bI0mHvRViw2l+9f+XH9fM7SsGLy9xx241Diz
XNwvs38npmT8ed0oBhKRwcv3y/kOnPuWV0KIbopC+go4RfeVMiKt9AuIgSirUO5w6xYh5TU/Tuc2
pjcpsaKvsD4vH7UD/3pqlVTRe7KG5k1L3etRotiF74xP6pLzTaqJVSEws2Bu+8Asb32NXZF8rYSu
z8Beu428cqDG7SckedCeDIdIkZabFzymmojj0Fm7cbviJjLwUzp+cqFQxMPJ3hCRUAir0DmY314h
t0sQEIA1bQZb+94YyWOW/iryV3MJAiNfnsxI7XMmaPFGbWu2+q07e7JYj9qbpBLDNa2Uq5Kk6DwY
xBCIbCdWYWD5R++VPboe18qHqDqdWU5rcofPOIKjpYE989ZnzX9GreFb1yGyoeSKKQ8EfuOnfIr1
tk+Q63ZfgHzhV6crskB5l7xLfv3IMBJNvwTom/Xh/cjTqIKtqyISMxPC2dqpdJYpiZ5DvTegVsx9
KEEC7KHbko5AsYEbq0c35gzsFQCbOAHIecGxIz3IA7oW72C488Zg+tt5kXYdJrNuYoMBROo7S6co
Fgh/mHQ61B7kY+HFjpgjOpEqXK2RZqrb5ZPQAN9m3ZRnRDZCYl7PE28whLOpxaii6Ao7hTpcW2cr
nqhrUCDh44sjM8AorsX2Wnr1Wq8hbMqb7g2WvLML+Xj27mC7NQ6LXfc8b7iGWflqAcwpranHRxUE
bcdyemAUc7gPefEWvdNtpYN+BUWzQhq8Vi3jpspH1y4MxPNRv4rdW9sAByDQ/ojbxjRsa05D9Gox
+jrvUZDkHKkWkGnwRNPvVTuSnBOs8IWebMlrCkZV02aYwvR9t6t1b8tAflKmOFI3VzEmMT1r3mrt
DfwAb5IoXXulf9RUWAoxsEmhe8Ft5OnEuFQj50Q+Sn7ja1fRPqRvU5TisflOdU18DXKLpUGVjTe1
skYRqKtEfLoH9V2B8jN6XH3fM+uS8ED1PpXTEHHJztYAQHoK4gNcH6N3BRtCBDaDncUl77WM+bjP
AYDMtlM0RRusHFK5tF7E83SU4gwMKIfRdo0p6TpUU6NRb0wh2zyDoSvHV5JMUJfhPBtPbjeAQ70f
b2sERWuIRF83YohryXKkjFxuwnQcgoeJIbRd1Aum0Zwh0Bbnfsnb0UjJLSKVjHroxuzfbj8RQp77
mvybKJKSW9BIKKA9i7hvtLcOIBI9HeJYA9lqrXBeup+HXvuY57IEQX9QNGlu6fRerd6ZchuobTGq
p9i7AFTRc2vDEqbp3VKvdA2Zy94NCnr0jNoqTuA6ZNruDy96COQ6/+GZG6jKPJT2M9MYZlKdWZsE
TagXUg0vfqGIDKDeHWok51mVSt9UcynZmvpL7iNZ0TQH+bTl2L16jBXS0/7M+/757Ml/DL4dyGs9
f/gls6tcOEvgSafqXds/5ltfIzLFLp4mq12NCeI2AUBFIUmoH8yfuZhob5EcgpEOLnBzcOqyjTpq
IjBLSEXJ2G/aWT42XtLDu/CH6gje2DNHieUSMs/Jv9YUFawyh4AHt+3DAmpje216W9ul9KzJcKPl
8hk49J7P/LiElFB0nBBVzkHQhQwZ8ZXSU8ErhzwjRQ9HIokg+0pNsMtOW7XYB8lMakV97ko8k6er
H0UD3rHHsLq2MwIpDX8v/a1VMFsaWm+H003w71LMD+BuCexYRnOKtxKcbszTrOt9WJ0iltiNi6ap
tm0JD8UXsrpo0Stxqio4RHNn1fNrzG/JbYlBZq5kkDRFWD/7iEpKMWGYQGkdHzxpqjGsFgWdjR/9
Ac3nhTjREmLSFDP4d2LdaL/I9H0RIICIO5qUjTcp1UNo7zfquq7VxKjqS3/RavLIB0MNs3s4GCxp
RXALXzErWIDGeSIDkEq6Mee9C73Bat36qRMnFRBbsl9PEuVfulBm+R+NIvy8N/mJ5hcJ+ClIOTad
o6YjTFxIFySPdHgv6pXo2IV1LNVk3/sAzKU2slWHQZhZq5pAM1d+MTErqV2pWYPGzEhfxiZ7Km3P
J+WeCPpkDOfsem0HyXZl3qHlMO8EL+DFgAVI3ARQZR9iSee0w/WynhtaFIxs0jIxq1Mxb8qUWft7
XxeP0GC/XIHLO+LUSUPKhJ+hP02n2HkVdMLI539AvZxa06quyKmjN+krU6AFzDIKxA+6x/Qn4aOJ
7cb2RTGRtHFVEusmJvwlEtU6qn7bXKUVBAJHPUrJphGcF8M2mHMHyYtfySGCrQjZ5y4gZCY9zUCV
ZT+VYD3wWVBNtpyc5qRNCwQlsGCIbtxS1fWeEx+N5phBrspMq8Dh8/rheMxg7iF1B9RiydPesP6X
NMyPykbhAGWv6j2J1a9DnnOpDtSz+qfS8BYDMfw4HBc1jIrSgZOvKBiy6dbx0rHch3NjD0rA/DgW
R2x+AOc7ZP3vOvX9Vnbvc47pseOgbIhtw6VeZUxsEalIVyK64KpTfoi5LiWgbQbMNwuxYPo+fyzk
C+GU4U/rPGF9sHzg8kH+c9VYJGtd6a+fb7frfIXcyaKHiJQdurNhGgHpjdB8s7TmWX05VC7ALleC
YkGTfaXhXH59dC2Szi2LsKD3frMEkaCIbi1F9O+tc9cj6RjuAyUL/qVq9K8+ZbJWhQ3eWiR58uZP
s3wC7Ee88jP5ym7ggeDPFbcseOYRgf25YjC47PzaVUEIY5XgOE496FEiGPjmQCuic+Yr/cetHv1r
m5V2BOUOC2hi8q7nqwi8M21HpP6aG6iNRUGEWyPQ4HOkAD9LaJ1v+A2N50SlQFbWp9TprAs8KAFA
0eRvqL5wiIbuRNDCTY09NumYwqjIJ67u1Oy+1Wt2NSZTEqF99yQr01WokWFoDuz7bOZyyIxiz/mY
UfnaByWjPX/YTUMH8X2PaqH+bJpL0HtwxWrXY3RTiY7Cxc5nwPgRl/p+DiUbHywGFPTeql2zqJz/
TsAoxek4fJItdaJDycYVA7MM1oHX381lgiHXl1/xvYR6VR+wVHKAK+0O2Qqkkbgoy2oWjPam+CIP
K2G/mKS4Z54OFv7Lw26BVjl+of5Am2BprabAh/Jtj/UUNMwSHwcB4ikc1imrOi4lS6/nw+nTdOur
YpqpD8l+eg6L02gTHdO3kf7QP0trfDRqDPkBW1FEaGwc5sM/jUuNr161Yxy/HGvlxNpbAO3CGe6f
VYmUzrp/MK8TwHTZhecJkxCHh2ivUttgbO+112WUoOdQixalwaRJIe24itbqKxOkjTqNb3776YW6
gPbjNEmMsJWFeFwQ06OGjUlAp+4lKTmvEhJrHThi95N91LMOyvoPHoVXGmxxNqSkk5hKBJSzq3Di
O4tpd/TxJ34TY4SLp2Tz72d6BhBZVxAWuAy53ng2zn6pvbRR5gmMeDc0Vr9Hw/UsuM0D4otLpbAT
IJ/HYFUrNYBj8o12lz1YYOqIJFwyImHM8AU7Nllh39gQYDb0dRSsO6COffVAr5Yi9BEyRAUU5TDL
UkYdLr8miEWGiz8V2pIp1dUcTYj7jEStSwguTq+4IxrC5Cdn6jE15VECM4H2box3XO6PCjoG1TK7
mV2H9QOIaNwNidO875gXcMSeiBcuJxczMm6hTItDI8Qp+tGG/v8Vk+1Rpnxby1WjonyleTws/koH
pfTRrJ8QCwJ3y1/ulVmPnvMMU99LAVQtezYGgjj2G6lyKmQn/i67lMYFfkp01wi1/8m17JcJDnti
CJxEH+pvNZ3OayXC1suR4DdsfY62vUfXmGN92SQgDnx6UU1c2AHnw3GNM6Kdyx/Jcfw8AWfxSq5u
tyQ35S1Xs9QGNzv/I5tTF9k4SkCgvLUwyEPA66ddUcAuIyjiMNZa/6hs9jRhAhZCxYrAhcGjdzR7
bSUKHHpOdqk+rs76lSUlgzfTeMAMZmE8OAMStrb7ds6W2Lbe31sVK838WI0oFxmHp34pfKfNQ94r
Shjvl3UfI7JonxcIf9Q/6YNC4co6wTLLp2PTz4/5ZJmiWcYaSTBVx/wSpAxVne2jJfqsHgSf88Ap
wW1YuMCTmmD/lOTMiE4EjEOvrXcPHcHfbhr6f6AtTXPzITyEHvHoNfCV4qLOi68+2+X7pxVG2ddJ
GqK6OmIGa4uWrKDlp5EMqFeWVUGasbv3AdwifjPUaaJdoVKQkgQigBp9al1PW12ROamS8UZT5Qzc
3Fm3SYd+Zy/+e8epGrBTeITfqlnQxmBZmBSk+ew+cceEkJBIK0PLtQPpXl1nkc/Km52adg/xd/TP
x0oT4j9ByQ+GIWJugWBfHVbqTrWI95ua6rengGTfca9SUVxB3NA64nzsqcJ/CxG6wU+sZHcnGG0g
cWdatCqACQ7BrhP+VvCF/LY616hzzKbxqofAx56jQ0J8ZyHlxk9rMa26YLXJh1xPhM83986GzYFr
dkghe9JfLtNMJQbsBuf7+dy18QFOj2H5nxkg8dztifBDE9tWEbKgKaOK30p79tvblIpNnwiscO9n
fYBw5tFyEMF+XxzNuLFfulHcLypMwXyUhCyKCTtxuPhR0Hdy1N9G+FZDUlZcR/xBP4waeuTfixR4
wyy3jtLtD/vRLC0YuUjOsmv77UH0OCZ7sXyY1KXKcohaV2XwJoTytLipZere0AZm8JtpOvFUBlta
DBE5VxQeBOBYbZZBr51O9zNwnN3qRZ5D1nvMy0DHPAp3Rxfyaz5EBrINJjOKdoPat20nyhmWbeNO
MWGP5E/bu7WQacPA4rsqE7Pj79zGcfi61PIssBZZIQDKJfgI4hWLPDOgKJLYcoChd5fQ5e7ORfqj
cjNSPWUwXuXkCe0hXWrYmIMN/POGaKko7bRvXX0RyFfdlN89Tou7n92iv/K/8MfYGQR19WqRvvqk
pR7bBPsPNUW5yev1Ln9q/qFcJTxpOBjJL/OYD0whOKa4V/jEaR0bJhYhYjwpeNm5W3TFpHHhGWjr
R/Agim8xWy+3QyGc2hU0uqAjQsgpJr+ujinplABY7C2KJCezpCkIvWmWcU6lqD8zH1Ds+o0SSnJ3
PlRK2z47wsIYDgY2YB2xiV/iaQPShb+xVMGPIGOszorxz5nOMQEXomaiMGUaYqJJnZEeP2wuu64m
MVGc2SEZL0bicj/m0i5i63mXGUp6dQ9WbifIE7exzSHrvwkUc8XNMbuCgFt7Q+PfxuoasmjvYA9p
v8yyfLFvA5JYfJ+il6agkoJ6oT7C43hUUOO+kGqD/2jSoK8pM3WL5kQ4nO2skTUu2A+zOljHQXh2
kFjYKo2tcW4Z/THnYS/bx9xPiWErBXRWFn6hwL/PoSzvQR0uphyZjCiVfdIderIrDN/GCgFJOlyC
Dd/Pj4iWg6sJUwe0d8vbYIEYOXu9jKFD2VGMkJ7PmpiWarLeYft8JP3vIMqWK9YQ7mK4GgeqKh0f
DpI1qlcphfsUirSTH9iyTZvfuYP+wdDRDKnMqBZ6PoFKbrYaen0w1fXP/mAPzGiA5bTB4gF1YG8S
N5umP9IzU+05Ss7CRY3KJ4YJx3k9gLjw++Ebwtm4zDWMZUJJ9NCisw2hY7HR3sxn3eBAzkxczfHd
NMK95tX+u/3F840sdQAMWmHQfvkXfzx/xb/bR4e1GFEEnakz7833OM0aT3v2IRBJS4k76nwJkgaU
yKRofodIw5NdJPL0nZgbXbQvoLFUosWuXA0LV+CQe7F7jmPug9bhV/9L8+NYHzfAWSJP0ji9O5hj
wL/WoWP77UfK7bICc6KgmUnsW0KjIabQM34dXK7CgPG4vafu8sTsttjBjPTWzFlWxfdjzJm4kjon
EF4actpw7vvTzF1jhfOVLR4k/wAXWAVMP1ivYw/UB34bd/mg91zeZBG7pAQJ12M0SDw0eOyczuAG
QAMbZAQZQpsnbwbXkBUehSkLV60eSmIVv8EYo13GUYirApOk2bxfi2+LdVU3xPcsq0My7Jbafkgi
Ps85gmtrwFwhR57xBtdTUr6v/3GPOYENJrfOvdeVhxRmYK80KcopotON0zdjYMIJAw5FgL53sQAw
pFPGyokiGCwMD1JTQS1rOxweXlryAaOAZLyHsNmOLy38kxn86TkTWG6+FI6yVM+bCA/TSBI+l7Cs
NpLygQ84QQCTBT5ZEqg6MnNWLSR0YjKYvzz1adDRv01371+YTJO4/4NKHUmORFfNqqYY9wf0RZxC
xnGctMVAyztp5c867AsHklB/cSbISRvYZLlO1uZkh6MCAPqfHRemjaFSwhGr4B2lN3XkVRDH6GRX
8X3+GbMGQzL7ZlkF7NAVw3enG1ba1Ju5+KhQ0EAlGzMIHo0bDIskkihCEIToZL3Lqd3x8NZgcD4W
AJ5oeEuQIrBQfddY5kngPR8PhJo8zWVjGthQtQM9thUOjW1afUI9sjuni/dIBmhwFRWeKjbXb4im
SV04lhhJCla6LgD4bDA2b9PtycDJM1eW/vYjUr+SUP45F6wEf1KNVchvpz2pv+X5cWZbKdVC3jlC
Qe130o5BIjvGJE1UOV51lMPjfj0myaKxlierBsJxrM9u4gosCOJCGuk3LjI+Zra3acj/e7xgTGUs
AOqCnDfiXq/WiaXZaj4Psi2+jdg1dnk0o5VLhsIwwMvGRy45CVomxMu8X8aFny0X6a4wfWxaiixF
bmH7BBD6UpJxtLQ7pn2rmlmmXTJbLId+XpN0TqIi/Pup6v6cHb5EVvKMaSaOzz3WkHyXsIVKIllk
IK40BWGrTLSFy22wsMWLKVJheeWS+qPzWCN0GFKbDmy2r5wglDikUCFl76UZtxRoY0t10mC0c+ny
XxMshoKZ7+5Pno8iFRIR+Q5JWaRAeRRdXDEk+6IQWKUkNedz+HTRmDGnStMXmJbzYxnZq5Yhv91I
1+rsbZV65vOIJ9HKkhWqtd+CppTB+KeL0AYsl4ogt+d0bWZ7tKLFsyUunNH4xBe93LWo2Put5Nob
06CMR6PngPL+GWnAXIFQqYz0s0asBWQvqAfLJLdTjM/k7ZDTPOvvkUJBBU6PpULxe1ShCO1pIf/0
udfaU9lHmKJlhw5jBu/7wrwZtBp7SU4yppU+Pd/KXuq8Fy4+dtQrhaxK+3sI/sCU8YNbPvQnyjoM
HilERg6Zk176NTp/Cgjyf9+Ol86chC7XF05VeNz88MsgyaU2/hyyeQmmbaNC/IkeBVZELh6u0eTk
pv6ejNPjtDbCnlnk0DR07uHEOhiJjLcqttkWbzA/ZhBB8JvwY/ws4kAo2jG8PTkSTGl1oxLrzzO7
h5IT3deTQwxE8+EZsl5548Bj/Lf2XAR8JyOWGXqDJcHmc3f62+s0vbHAga+mTEkXit6C4VXXFVEA
mbuv8+ly3z1cFpryFqtE0kraCNwcjTsypPOjHJ31/k7KRJyaIWyKY/9jrcUmeXjr4Ief1ECqZcWy
dXPTKUEofa9bGV2Qbj4IcAM6aWyvtFML3uxq85k10wXujFDmFyqM61laB75/rB6IWxodMHt5/1R2
b2/fSzJqSTB5GoDZ6n63vWfh7Qjw/NSNgHO0csePAt6OdYrCY3trKFF7+r28qoGz4cubcvjtTTi7
hrb+8f4Q/fJggvjcqJdplN4ulHrg8nLh4dyJf8PvACm7q2T0bMol3xuEzKLnjWJthcsOjtBK43nS
bNdwDfPuLLbE6Kpp00BtHizllz2uPHNlXnpw0YUWc4NSPMn8K/fyZWhseOUnxhlZRs5FiYGASRmd
b/g04ObEEJEeL0a4L7sqKXHk9ICML44a0bTBVBWACnHpNpdgiTZojv/qZ7j8LjbL74UsxnHrlZ6R
4DfSpDmPBlfM1YuKldt9vae8f2RUKWy01uLowEQOlkszmj3GCqtDrtXeLROM82nI0fyIw58bsMzD
oQ/ERW+k4PX07PLdwUarRmOPkHXXlSthbQ54/ZS/+OSueZnjZRf8SjMiTD7QgG7PSPjN5rphTzfy
Tk6fe+UCTIggWrWBmKQJkoPds6AgE852n79Hxl8+nBkWSe1mlQFx20swf0pwtvPcwvr6JOQONFdY
7L8WyM2lBH0VCXmHyQkNHwPXkDsYBANk0m4M5AyWxh2O2h8MHFk0TBN1rSyRZe3WgSS5ziNjE5PF
ZO9wwxq825+t2TyaSOm/+LzGgDr9BghpHKpfSWMkFOY++WrKpduOX7qyN4wZsXmpyXEr3HuI2pLH
oFh0M69LOo2xu22rHO+nquwgrp+qJbZs/uU00h5v3jiak4B6v2VeYVicwbcwYfgUzpqAdJewu3g9
yUR8m0gbbHUp2V8FQW5wTLk9ERLEYWL3XTNzkcu33pAERBdbztT8jDIVFrbOsx0Ww4/Agf1c2Kv/
Wne6QTjoS2jdenjUYUuvbwYDYhMQE7ztuaeYeX0imcObEVQooio79Fy1EHz3Tzp7PsKz1yPbvMZl
LgWe6zYp1A4KD090cl4ECI9weQrGlNrYYoQkeKZ1dbU/vsYtpTKUhk5r+CwNpGKB8/jk5qs0z6Yp
uc5mwmhHHfTo7fas5VOneX4wWW3P2szbgrp0ePvcqLc8cZq9/ZQ5CUc9voNEFqtOI31gQZFYPoi0
TMHTL+CCr/4vMD3O7yynoROc63ZEqgPjQDvZ1il4LYtZughOWahgUtcplG5/JkFB7BDMajor3rzA
ONNMTFLDrtaZpharBNFndvuuFf+sH8HuH5EHEjYPijV9bkcvevMjbPnHuPUO+OxXHl52725u1s6L
80zpaSWvJ5LXg0jKiXo5H/pd9AisgnjbqdQyGeATHyM6gOc9aH9q0Guag6kLTFi+wE16DT0mucUF
4SUw+d3QJy/A6fnINAvIKccjp1ZtgiLpLXvyhv5fAvVLGOIMuLrZxN1srSqnvgFglIYtSMFi0uJj
RQ4Csbc9P+PRmgQtrSbxrxGV6zGNiHgSPg/3drC8SWY/Iejor/Pq2SsEMa3MtM7OBiNzpsR4nmf5
RMGEieIJ8b2zJ8VhyedNw/tjj9I385PGxLLluqJvEY9HLNGbhca9K/1jzyOPtiJrCTuPIg2Whb+f
VRkMh37v+OURZ+0vMmgWGwUpyBJzNQlCwW9qNlQqTSRTS+0rU9fcxJ62I01jKmiXANIdQWMkHavR
f7rAyERG43drWzPSwe3JeN2SOsgJKrRZQvNOSLPydF8hfgHZGCy4oke02BSOi74mE7Zh9b4S1DH+
InOYLiOv6NaTE3RYhIW86IzgCKaGpl1/5fKr+d9eBW7/qe0fJajNEFbxJ2JWVulJ/a8+3kj3Vaf0
rRn6dj7eU6PyX9s4jFAE224xjwHio3yHyjr6yCUJgHr6hllds9WbLbVO1/RyvrIWDDrES9WDqXUV
cGzwpyGnKbJeQJ6RdMd+nn4m6CUXZoHHKkWSkkvNheP2BmonAM7KWhsuvdt3FvoCRkltxqtSEfDV
nBEngsI03CM8zqWl+vzV40RrSsF/71Yqk5s9vXRxnVfh2aTszom9EqK+PvdiyDIa0EGQ1q0EslXE
xQ86I2D7yhQgLf6fa/7pdVYtFjXkOKGEuO3fAhCdMJnle9Dt+dhzdK3+P+TtExAf5xAE1Obe6In0
nQt2rLO5UK4GCRhUAUrZ7tjWUwyawr65k0QuC3yifGraEZrCvVhNv1SSdkehZbQ6eQNhhAU0iac6
/NLepBd0yMGMR7tj2d2k1aw5oVk/hS3ZAG7WErAyZYLler1E1WHcPx1v5ZEAGcT45Qy7Q8nv8msK
iUJI0IoJkyl4yRiNV6jnx6051m2fJ1idpNIZnd5k8PSCwQwFb9Hzp7VijffK7OQ9jaSdQKyhmVZA
UrJyguW7n5/Hj9eeCSGS9/R9fr5ZBgXIRe1x6cbTb1O6XF6mHM3wPsnsp5KHfaSt9Qom41QyLFyi
+W75/lwv3BKuBkKWBT7XPLGLLe+AmFWFKxEcTHaJ3lhiabrx9S/9u/F4sCUMlqu5KCROJvXOkHHc
ntCCbCxUFlDlsucwB4zLojJYcrCkuKQbXeg0p5b3D7vxkf5GHD/Du695RIvfYvgZ4ZtiJV/RP76G
XbHL4SXpCz1nX53tPUbfzxwrkazQPG6Zvv4KVrGG8+8lcTqrVksOQTgfXhIa+gf1BfnfLGiJHWhN
6Yols5WCVmAe9O8BauKC/dw4Z+DStKYWiNP5PwCglrqlIeb0hKIDaD+VetAugbQoR3vVLQFb6NUy
jwEeTyessms0FJQdggf8rmqPcaXkjqWEZfr4WCTTe11T52Z3GTqOhaxIHoJv8MsWXowBedu7FM/M
OQB0ZWQukrzio5KS5LTBrqG3QSRUPu/TBWpnLCYO4tJjfV3x6orKL4POrjz1LwttfBj74z/ccwiD
5qTqTwOVC0yo4nIQyQj2UChOyrN4PvN3VNUCxnq7Ap0k7WnzMgnTQFJqCwtCxNAmmcChQQpBVXu+
jqdyRNb6cjfbhd0g/jG2rW85eYnyojhQDyVdfEg7/MuRHE/V1wlrIWujEExN62HCyjEmQryUXvEr
QIA1B5glwwnsjKfVxUX8INRCe0L55C7TqCt7tYDN726fNQo09LkU/hy3DoBDxiQf/WrTQm5NjlZQ
Bn31RjQ/QllRthwU0vSjmvSZ0CpaDjLVhLtJd0f57jaEOBM4rgycZ71t69GSo1z6BKjG5/PRhTAd
OkS5gOT1hyqu7iRmqw52lMno1HJQQyPIstxatH5KuPOanwAVedObzQ3x6BOTK/a24sIZ8ftEXqsx
6aDhWGJXlCDnwT91L3t/1xBDSEYO5D25NSiQbSui/cLVicbjiOHFTzxRWisVr782eNkaMvt+M+De
++n5opsGKonZy0i1HSNaEgGhVhLADewBQQV2KsHMRBulRWiaP4q4CO4c5C+9eFnjM1krrMsu/znS
vbFxnJTbfcjwWlwD5dPuJLz0727jV4V9ayRaV7IHCHK8cvXOPp/y+IuqQxGG5bk/srKmrrM8h7qF
mP7ZWwfvcSCzODXtm7o40NlQ+oNXgBUKPBOMnvDFtSdQo0MftO6sQnVrmj80UlPx2fAb5jHu5+Cw
UsAZQvP4A1qa2gfzVPX2XGvfT2gSlCeUKDNM6A8bL86HdObDCgfA3DeKCHdV4V5yM86JzfDSBi6B
/MLOI9HATJ+MdX+o/CRLoRhu0/eFcr/iB20wXMhniMthKM0x/Uc5dv29roJqZlhv5a6r0UI9mMj5
gPBUx+W1/IfKAkFxU7KtvIRQ6wLrZtgmN0Cznxcm7aYgXxseKHvKAFJxJs7M8d6yj1SlVuITY4Le
WEyoUt36aHUkK0pCAw+QSLUD51RjnmC6dJz2vPrCZ706cZgdriJnyfu6QM980CGGuVX+7APcalr3
Mt6MhsvhkHrR/uK/HGS6Oih+Zx5I1REI32uIS+K95GbQTotYMj9J94SR9c9KfUr8VddYojv+WJde
U6f/2XIM2ItU6DlAC73D31tRStnE/vusANn41rudf02xqHf1kMSAJaDkTZV+JKnd0G4bayZkJ5Lw
0k+yV2J8tCxWozCOirIn0hmLWoZchLMXeTBQg3G9G9UFEu5u+nD9ue9mhzOAlMciqo/ed++Fp0nV
nTBz9Dx+xWDBynwwKZvU9Qd4Wq+mWEhrLbJxsCGOeTTQH/iiHSWWpmDj2gTySQbL5xHfYC0Yp9B9
pwvvrYIl0eMnmy/Eq4GzQDPz+ZiFd/OjtqgzRu4rHprY3iDwYUiXb5rLD7Vqnu+r/y7fw6H0OosZ
MWgGsrcpv1av/iIUMw499L3zIYPxDcPbF6qhwRIHIriowTZF+5IKBcIVjl333ziVb0hICJM58HrV
dj1ei+s3/I1ylPxVUv69jV4xAJ8l8GvHRZinjKMEMSS+PD4fKNXqza96B+YVlL8FHUtGG/0SK+Ht
CSZRwQqpMq2+LZqe/7IqTqOm7xEaXJFN+1X9TXKSAxHTWerjqRqGdzjOrOhvuEVCzaCb77IGu5ro
lI4t12llSNRzIxpwLguoHBySU102WVdlskggqZE2wurebrmH7a5nwyaTuCEEEFynvJJxIfj/SviT
h+qJ0yGra1zm3H75KfV5PjPN3QIcnqAT9LdOpBgBJAzFstiyQFKqJVNxgB6GRBUoKpcbhAJtd/9E
8DlejZHO7ioGbyTDL4hXh9fbs7h9Vg9bjXxghCBqJT1FoC/I554lAMxCxtKskik6EDaM6bkz9kYg
JYWZfAe8k+fxWTjiXNNwgn/6dQO2wA7rGNlgGTdNTJW7RMqi8c0iWAWxyeNt9qJ0k7SIMtyQydIP
i09UwdZW63KSazIBRj6oTo6akcPdn1QSvKMPrS1+t/R2XOVIr7URItp6X1Bzknr8NVtuzk7qIUbd
g9hNgkBAYEPhZSPY4ikoSiylOhonFYx5WwCnLex2vHbdzzpyZb4NYIJHgJ/Vb1tSbcvLPudIXRep
SwDIIEcKzzEDJYIcwbJ1btgMaemLtVXy/EHmbtTijF7oCGBth4XRpIOqEmWi0TW39nkMBxp5hyEp
mMDB7xSE48YHtXREVGrEx6v9bxoPFt5BOD1siZlKQ05oKCfNGMAShvrEMFcV08CAd0P5k4CxG2V6
8CTi3MlzzIqabddlIFiJFHnN3IEPCPfiJPTsi0N9CUbCHRzeSz7v7qRwRUgzzlB3I0ifRruUFE+E
kmenIRrrACa8V6nPc901KDVvt8dwBsNG9gdvbEBnh5KDz7fWH7OQcqkSmLrjkENcC4f6ZWOfrmu7
Th3rvvCF+UWFLETUdYbXws3RgTP+lxW150AVpoX9mf57QS6cDVA8Ce7FTKfgRUt4uy8KjRoZGBaK
ByBUMMRSBi2UkGhC30hkYkN43x/wxwsdF4SifQjwB8aUXCodpvrxhPlCzGTD7UvhkwZOCZ8Ndc3a
UZGJDhlW1tXlSMtNptoq4xflOCyNtVvBU1t+MmZy7j0l+9BMyuWFqxtkbrKd2CuRjcIPLthzXsxv
dzbD/ZVDSvyJjty8rif7cNG7Qo+a/hGacC0/zFmvqm1dv5cBUOIJoAMgsB60pcDuP8IuXBakTuv6
sbBk762WQhPj2PmejklCG14ffvAaiBOVeE0oh24YZz/slotfIL20F0D9lTnHddxJ6Z/6r18bxybq
tdwjXiOoCf0WesjCjNvMLcJrMQ5Cvsp9l0tl/GnBJXTHtnCGNhLfkarX8mhzwV6I4lBnPbX1AfZZ
8qnT6510BHSAFF1wJDCyH95EJ4XbJjxt+0qJGEkCYYSKaV7+cget1YySxx5WsJjZ6bna7qvgw+6q
rYhvlbjMklVGQmAuZDBQTN69cphBNd1ea0k3A3+uFlTPXDlO+hiMtWsWvzMSwF9Ox8tzof/joiy+
8vt88Hg5aWn2keU3VgyCaioxXiBUgxN6ECd3zq+PVMMLkJgMlcrmRL5mJzUslDHmSVxlGwav/DqZ
q0KlCEP+CJv/4n8Kb16gBo0vvt/xfX+lXFUJnHLYUObUqSlpgdamOjO8j/VENZVjTOnFGeTjzvQx
Rjv8etVJodwtOeEOyuhPqsIC4gr6uX1JmJSlE6zhp1A4MM19hgRL5qb//vPqNvVZ7myfW31f1VVh
Ma1wscHJGpapk2zPrBZhvwvTf558DIT6ECoQRLA0PvaxlqE3PdwLMysg10iqkrKzpPvviEPGtZMm
KwoZq4hsQgCeAfLzK1ztHx/4iJESYSgsNDUUs6DkG+lgxciBrcMDJMNP8Xblvu6+wSJCf2LOVUlv
rsfr8FgmnTTFZD9J9aA+onFezKi03L3dR+9uW/fxrl8GxY2vuIlHoqCvBpUJVRio8sPuHS2tpZFb
LsdT/whvwOAHbGXV6DTS0ey9q5L2nsMgGQSO7P9Gk6UbE0t9ONfBDH10qIyiNirn1BPgISX5pk3g
3JslJ1Gp7fXWAYtXGSMhVJ+9MFv9krmzTNfWqDws3AK9GqxkRQbyhLQxkYc1SIOr4ukCafJ6hRnM
7+SR6VsNlsPGhlfu21SAL0wE/Y32o3pzQhQxpei0gKko2C6FOMcr1/64DZsqaYLrbqLjND0JI7R8
whYZtW55rp3QIPDLuJTHtYSGq4/Wvm8b6JKHQ938XEYitvPpOtBzJyWGNq4muLFQ/6HaaCPh9cDj
6Mmbq8ULSiiN9cop/tmUj4pziR90ePDA46krZ+/0+tC82sHbOiRGhFfJC9GOeCJH58ld2G6JvZCG
fVzIgPxQfWtAiTKBJPmf73DbiOT1OEi/klVMH9yaOzO92ZwuZQiGsBLGCkxj0Th25Wb6RKMlx0wN
3JrPuhvNcMhxTJHGUlMxE/JiHunAppJZgTXjWycp27lAtTsQnZv+2LL7nw3flDUrsgD3C3ol8HWp
OS/IeMgFHy+XBBJsVXxA8Vjqf7pxz7IffJami6cEE8IPG4AC4BERycuOYjAdQeCPwYYUM1mzWUg5
KsEd3lNwJYnYe80enxnlQE60GWPUyfbkdbDv0TEzLalHFn3SoyV8VHkpn5GZ7hWmQ9/Dr7VIhoyI
68deicMLmXIU5/4fhRcxUEt/JFuB/bkI4blFvojQzmX/TxAvhWZhmP5ACxTgChuI+7KphA7pFct/
8a7WkbHeSEvY+i+lA22VKqEmez5vjyLJlRf75GYIZtACOSf9f8nO3lgP1CtspC7Vr6hROP5OaIrP
Kf+EAAZwQXAuwLd8bBDvz9wgf6UrTBhVEtRQRiiIZduoBzJ6k8nqIT3YeGgMLhjhe6kFuZCHQvU9
GjtT44jMkLlkpYdLAC5CAaaU64q+f8HIZ0YPkgyILhFjJzNoq8O4rwQH4AsSQePNY7m3VLU0206t
oa+QcpNFxfev70XVrSOwkYK66aEAFUmMnLh19uAis4PCwCeujqN1tU68TW/GstMs7RCDl0XqnR79
D1SNxFxxC1LOqC1+7mDnu7LZi0YArAanNw8I62YsRQHagacnPIKhmkC5CiKIefxZ4QOyX7gzxpwz
tiW2AfoboHGmzrrciZbZ4LEn09dDhTZSI6f/GgEBNs334bVhxxWIAK624eoUantH1eQ8AK06KxQa
KdvMuOZTHmbqdc416kDhWalZqMaJE+g7XGWLjdr6CwaIV1Z4dWbk/m9TJFrHJLXzok4zz5AGXAF2
0Ubpa+rlaQIiawSuxdBhIPZ+rIeNtprJM9JXTjZkOJ6EP9SYLi9eMWE+tgp7VQ917efdmGn7CiiI
C7qrnIkpZfDB4wvYhvL2R2cMoVr4z44uAZoZOGcgAJLHh37A54KqDeYwEZBuKlQ1iubbYqXSa5fq
fi6OnzhDOZH8uKncpyyayLETKVFttHiepI9M+9hzzIXdeIfjAhp2aioycw58xyGuVeqYYXmcuDkW
rUuYjPG2xCKd0ohjCNhmNysJSnwegNwK7OLjiI34LM/w+yzkQ7yKpHzo7Ca48d7U5C1x3UgkTeli
tcChZePCDoUYxGPKX7IrClSaONaKHdpMxVnkAV5HV+TnWnMyy63UTnCcSSxGATS8HvDamKxesiLp
L1SmK75oWJzp3scHdAjq4okBJ5gLVgR5tQ51dLlL3U/sXpbWYBJ6zjfXyG3Os3HQZo1CMyhqNv0D
+svh5bkcIY/q7kNIvk27JQHyEUvjHVzUpk2fxngvOvmZZGyV3H/HwsnIKc8gIbdYx5tByGM9yEL2
aeXRo8iuUlhsyFwqCxpve7EHU/Tm4Lw0ft7m/GSNxdHlphvgiAAxrNLcVaVxrwNr5O+teVbkcD4s
MyUCjIxJ4kJFq39pT9C7uHCP0g61k3MdPif7jNW8IV8ig2YOwBw1xfYDyhy2CNSw3uuZfynD3tbN
IjF4ILoRQUbLOCWxHCMo6fKk+DMOdmTPRCKCaos+1RzQngDIn2cpO0nh8Nf6AKw+3WfGypWU1KlR
/hXjjoNTHttgMESJWNydAPNDSf3qZI5mXdUTFVIWWijCS1+A/iZktrkyO+nVK+djh8RZ8Jo8O1DP
wPf9oWPEF/xxW3G61iSO604YBBEZcyZmbAYL/zVcIj3+mUj/9XQHIAS95COBvSB2tCRiVQwvLSZx
NYsCHEd4YjqT3bc8Y4CeWJgUrqw69PMkPsPHapvXfPmE6mdh5GE1xHIWEmBHMU6j0YGJwXpxY6cP
0YCSQ1DJc4KXnL9tVv6zfXmj+TLP0hHk6E5dcDHNnqV+G2YjfBj/KibP0K76RyZZXfKarofJ2srZ
dipJPqDk+X4/J1D7+9n+0BllTSGzxnM+N6ZcdfjEUxZKoz2ZhybdzssM2niFBCODB4cBDIZGmAon
2uwIgXOtcB95JdrVGID0hOeYAe7w7E85iP8VzMhJCHhHdmzm97O5roy78RrKNStKoietX+B0q2J4
APxNpglEOHb84HjGturJDfrV1xM/Y+caX1BWGY0q2eA55+z+tUykkF8thD8V1TGKtpzfq/6toLhV
/YJKYcbBqSEJDTLhBQCBoFJzthMCK0NQvI4AKl3zzZkGC1fViyITC5ph5eqHQdLLA6fWz6KuTa7z
uYwtg0sBY88uYRZInZaikfs6IarmMRbguwk9V4VfI3+pgF8EZAwcWE5QaVRWmNW7YvacglHWJsOJ
BvhvPSv0XkH3qvFbmPQIfL7jSdurWx3uivFYrFS4SMxXYWFesbp8SKvRgXQRqT6jRlYdc20DClxa
dGFIuRa6EP2PiN+p7hH3G9EF18ZpfVU0x3WqBr1Y86LFPOdzmuH7niEE2VMbQvvO0YJGWdqmCS/u
YSd8nuRSJe/YuPSqUg5xFyZu9BXQHRbpip+9BLwUTYp5LzePJGYqT6I5OUj3LlCh5GySHwApaaYE
qI+PnYCADOtm76XSpZCY9bPzW89WInfhKxhIff+m5vD1Z12vy5r/gDJ63j8hkKhV0QimZvIbeJn9
ziqA1IYjoruxc/Pc4e/hTJzxwA3MFtt61UPztCeAIfJin2QBbLSfBS86crL0EeaxJd3SS0MHtFo1
kGdxkRrkucxY3Ax1dPkLK1YY5fRoRmwMFDrhUdA8sWGqh4nJMbIHWoe7XLSVztumv1UUYCy3IOcp
Gchc8ieh/8vUjNYqy5n2vAbKAfC7DYBeGKAWP4TEuXrqUWTiTVUx4qMD7sumxmea5Ty87S+3/W6g
FtiIdTIaREyRS5e1CGZrbSb1fxzmJShJmjdAb1QlUBMMGQDXysdL877e+BjxdlvC/zlpqMBiCvzW
0maMzuQSwdkas25NBQPq0A7PCgRwBOw+HR8wN7xe5R9f+NO0AxvzoeLiczgVnRmcVfyKWLY+6OTh
Fc2cjPm6seTwAy3b5sJzlJjiis3HFJF9zItRxr7Ql3rKdBXW4L4EnaR4BY4B8awdyJAEOHHmoW6m
ggijbzB2lR9oK+JkooBzq7Q9VVPJPppPwuWW2GOKJLkOAeyufVB7zhtohsZYzW1EjpeaOeeZm+iI
j7pTYBVrj8uypRd4KNeMr7rFqwn9wsMopi6OsqXAqEN0F+OzYdai9xiajRzwGHFLUghSUWrDSxec
TqrV6iYH628vSJD0K6kW1+j91YGmYzPDSu9onaLn7Hcr6+TK/KvWPkhXtnwyiSePjDrGzHVoI9Rt
OgHetXeP3KaRPPVNwmdeE+7DiY49R5EGPeRBeBfmT+Euqdc64rvUmfQdmaGV1by1X4UnL3hjsrqs
FdfRWurUHchIv0iBq0dbWcxMs6widmCms7enCiNbNkMeBh4pjcPvJU29TM8TrHAbsfgxuiQ3mpBz
zGJCLOanQCg/KkGqYBVs8mxKx+GnruzTReVr/gKYW2pEM0/fPNqRchxbc8ddsW/ZM+CKbGLYXrOh
3tQJlexRsAInKIkb1KKMDE65aGHdsncjHQkU7vJn+SfQU3KbKVZG6oe+7q+4mdHY2yfhZkrCgOJw
ylNILKC/rVtyefU9Kfm+3FFr5wgPU8ZggYfqlrb5rYgrUrQxyK5R5QfyB1JKeakCxHQGGtMjvYGl
5k5tzXq4P4BdljGnrnpBBD090oxxWfu26sekKsEqjb83sO3goc6i6TGrIvpQIY2rQa/tBjTQBro6
P4RimTwagwSy6aAtRnGh1MbaWrr5gn8HKeMYwiV7DjR+8E87SxWIqznP4R0DHP3cyJ+i/5F8wI91
SSvm68q30er2Cv3jpp4ydGX0yT91+RxHGiq9yYrecOBdk2GiMZh7BTqT8SRJzzeE9IgzsfH2Mjx4
eqA3l8jv00+TJ3/NmhaLYAuDjurIKLeQp2nLvIEl9GTED5R0RLY9k6YENIjflQjbzHYle8nyPQm2
hm9SPcqbH1puYHkrpR+LEkqCq6A4tcnkWheLo7f655qkIGevR4FH9wVeWbs9ivnn2vOBpOiDAjEw
EP/PPDMP3xzuCI642xKUkDWxXsneY8pgiHQWyWPaB9Y3sxmRFVnnJbQH1mi5gqCt0NkWJbo1JFsZ
wLSgjUi8u3Nyj3jYJBlDj1YW0HE3MvOGImnO4pD90+gWPitt0lPHhCQKg5KKBLiU069Lak3lRStf
NDUjWketeYXyX5VGuTmM3szSUY0HWwrU4/+hp0aBu5jtiPc+OTGraGpwno7EibdkXM5hsrVwv7eP
94rPszn6UPdKOazDMm7ESAMHTruX5L6Y1AVf50BB2Jkk9PVNMYEuWOaT2hmVp3NJTaRLjF11d2Gt
Ohxv9vqhSHYOW3avt18TLiHbseJd636IiL1m5zDzGvfT8RFGEufWzVHt7gFQobgZ9xdTLkkDHRRW
Y7UXK6QOP+fdISGRi+03ZG1AWivR2noFYal07SvPqfmaWyujmEZLXarNIk1uOmZD9JxM/zX6E2Kt
GToDo0boIzE/oGHHJh+x5dFAyHLiMnyL+dGOJDKKPr64hG9lHrqsEHjAtjntx8xCGnl7wfvK+20p
Zu3NR5aDKQ5VcGdukyPnnojarj/YKf6hEu/Hjm4NLDNV/zpLwBiuyxik5eE/N68SJn913zWZc9dF
eumX/Mu8iyJ1PgtEtJV9RlNoMfFLZzoH2Py2tmLSrpfQTPqrZir+Yao2YIe8cMbZrOBiBJ78br3O
zbPItqta4FHiakb4FxOadwRABSL/gL7u4BsiDq+7MOxt32fAXCFammKeedX9/LQydCZvNDdkB76Z
K4k1ByGq8lbxp7TYqfvmTJmERiPVpyA+LL7zp/qi2qubGzw8MXU5++2z0XlJVc67jmHvVO+F/X1F
R/8bfPRtF/c5UONXQG7uBxP4n1vZV5D5J7qhdJumP/mfucDP1YXoDq1RzPjYK2mDgOI8svTxdmq9
XEsP8jUxnTuWfYNBxIGsnwKnMjtHNuIFcnRlGuM41atTBeuFbKmoLIZfzDk2bUEnm/gxioW0ffgY
R258eIvQ5Qg0sTPBHTDr7YwhNb0bBVsoY2zWklUqyn59qT3azXXLCTP0YdQwlKRf+0/6+ApyYJs3
/byzyCDHn3BVkeFUq9caiRKQTIc8dTWU8zBA/uT6nsYgpsgXKjWSgNZ3Fa1ARjmVwEfezw1K0H8t
Us+ccyvOvlaJ0ZqJiJ7vyochDQeeWvpRaQQ0s3YP/FUD+6RhJD3BY9WvQioALUzSdOeCq8Olat1d
RVN7ovlYtP0EM6E0/JXXv0S9NsxRnbeJ+STSsd/XIibXGlV5AbpbNnCktRrg1wdJEp9R765taWjh
bjq0E2VrApMsshfHba1hprvg0VKRfmXdVWFCZ1Jp0dhRs79axo4Zmi1OUt7SC5lzmKp6hD52bP5H
DGXL0PpXIuKUX+cSjjwtGKV0n/cXkvFhUzYBFBxFt/EudhDCdFQUM8cIPWlpk8G4GDdNgN1jJKbk
oAItz0ounAyfllLkXGkWDRF4QQtJw5nLBU/GA1/kxsuI8mfp5+MgWh7Jzpy1/C6Ea0pq9bHU1KUq
UhDSaw76grsvyR4YWgZJB4fjEX50nRk0aLdzTFVYFMBqA3ALD07Wfh3oPUoCtAfbQc+UO04k68k6
hdDR3Vel6EPIDU5aNxLvg7oUY6H8kZxUAgmpfAn/xrG0vIo79MAxiif69vbPDVVAyta/RiVC4ITN
tU320a8d+NeuUsoIXsIsCTTA7qblvwSI3z5F6RuKsSJttPZSZ7gqadGkE8H3og9+BVAzwV0nWBbX
w58F24c2P3h4CQaJ1NXLl2i/zIkuHHs9z6t/4BQQhy+V9Ds8DMr2T5U4CYdpildS8oJAD+n2steA
uAPrzFZXc3OhL16SMweC4wqYDPqTkZ/Ffc6VZ8yNQ6mjYkPTAeUk01jI/jJuG2mFxB7jHX0QSZ1N
U0C/CA1Ujullrgbl9EjpuKgorliOhILsti1p7PHLsoEHvoKOAqtBYyxkBox+XNd8qhvZJuHht/OT
2QFyb3x8BkcoVbBkPRASOVRYecJb4Y+luU93qY836JIZvcnJ13hPrwn+6B3B6Nw34LIu5TpLCDCt
50uE9Zt2HNUcCdQpkwFSD0zUHpG+wNfyK/vrDoq0voLI0yTJp13qEAQ2A2y0cl5TMfziIww0e0M3
DPbIYZFu81nkkxDU5ekLYSX8cva9cO6ycmGkdoVXxYpEcNpzZrHVKTCV+4oIfMCAWV9v0e2l5zf5
I1/8q3lXZUhqi1BqmhUfasKXksVwWbCzvHD6eid2GeaSQc2RPI6skhjukKlghSH2DzaTtF3Pm4Ic
vPEaq7uUSbqmHTaPfJ+U0rInZ6IL2pdMvVUdpuetxqc7vZ6J7RD8Q6wcNgkg4PjfHL5xiJuXV7pl
4APARt4UV2Gm0+E5sWBI8Nm0fkLw5TVSDBBO8p3b7gKNMUd3yR4ob83L6dlH3TY3eF1ukFSHFVzZ
TX/FnSo5pYZRBcCzsQYVlxzruEwkrUtW48FAWWFdvtFjO0P9P6uMN7RXUHG8Yj00xUf+aLR6vZ3x
HV5xMIbsFZrei8PDlLnRDs6Dc3eTWL5/gq6lKwUR2WVX76GJH2yhkI22vlAEzqVKPEuf2E/nUJCP
byidmdM28q/U98LVrLcOTMM35q4EVdSyoTC351c/OZJw2m+cUGQDtTiwGM2w4O/YkK6yToXp0ZkK
nprHu3IRqhguFAsMi6/T2Qc6E7tcltqceTfQOqS9TEki9ajKPrcvxXuCYsdyWySRuohIXzVpaev9
KCuZ/EECTBH1YRzWHZinNlRiyGcBpOk0q3N7RCtePmh00oA01yeUlEEDc2ZQXKFXAJXU80C2vHBY
a4+0DUXgyf2jr+QCinapk3GFicKLYh0PrudjYxB8FLzItOlnnxxff/iWiB/KFrBtnis64kaMHgHb
x3PILK0eYYCSVQwrY0sw1/GL1lgtt+qN40mWdb/MNgPDsyzlvKAze2r5YhShTBhflMukWe6f1oGa
GBuFuC7XAW4kO6dcQJ61FKf+xNyOhj3bVN8NBCc8CcXLbQFyJOwD1L35IqR73Oj/LjUhDLdvXdnC
Sj6zLxbdhN1gyaTGuQ+s/kxsJ8+YYWP02BX4YqoLtLWUAgy0GA8dYJk5nFk5iLMrzDw0M8Ryrc+V
xJOcBooCtjl8QvV/Pp9OwdfyEewwAI+aASwtpg1/y5d5exCvLKIDEPVusEps322GeePy9bv+H925
APfMB659Hjed/FLnL34sQfwxhG8rbbN7UZGwBjvDAE22+XkOdEt9yA6cCsY3VVnUL21Iy65uxk9f
6e/LLT5cM4QIcJqkOm2ibbpn8yEjBLh7emx2gL6eBL7R6qmft0zTQ5c+HPGs3SQz7jxKrVytxSwM
s739USZJHu+s4n32kBbE6V6E+x1JxVCYdVJtQk5B71+N36zm6/ZQKNEDmHUUQI+S04dMmh/pNHK7
6aQ9WCMabcbb6MzMAKCt+A3rQOX9mOm/CgH0d020eyUjqqziBD86PesV85gpcRRjv8Bz5hFXm8R+
SXS/2tjBE3R1Ek/iRx79nEY2DOnrve117m3mUY/s8iPF1iJQFBHtbHK+XRsqDVD7FvDYbiq3jUy/
N0M44/EmnjIn4zN3cZbh43ZNOQxr9Iev2kt+O0UCxDjxtq0EgNxmizZ+nDwU0nyrB5Nd8eW1HjMU
V93VQucVeqHLbLi3i4RJXWT4V3B6FSiLugyp+ysthzclKXIcwRepnMi/3/YHfng5hLp+Wen++De0
2/N1slHG8CZGPPK8YDpvrQu/PtUkRdr6eGo00FTN0sGJrAbBQIeaAS9ikqF6+NWdZn+DH0pTDf2I
R2t5gs8PR+7vBN12j3xCcwA8ew3t1glZBoV6CIYQEkh9ck4jq8x5m5paKHBljtNKGPJKFh8hMFy0
OzPC6vw29FMt+RANjpgm53p86GK0/FMrStEmwH2N6jqSeLBqKzTARRL9pe3hqzYBLztu26CHMjKX
cYboGCqvR9OtcXV6zEVghjCHVqYvZSr5+c++0valE/WUanoxQbaM0FeH5DoHiuWZWCVqUN+vV4jT
94Qp8cTzE2ly0yPL+sHu0Ntu56i7asp6LM9AOa6BnoV91YfsYYodU64ymzDPXoed2lnl2OlqFv3h
N7vUApNcMFfJ9J30kNnlnK6PkJhPXcGGlgbMXN0CZvhhGJ2cNSThqwNR2PzK7YOnq0iD/od11zvC
CpAsJ5N7PEfmNIPNGvIC93Tfb1DZc23qN7K2gX6NjxwKdogR0qSnXiTijYkDOjBlmowNkPg1D/dF
gw0VuRLOJdydQc+x1TKlQWoAlT8IL7pLhNWn4GsyG6TV78QWyQUt3jPN9Sv4ggdkB9LfVMeKClZ6
LvyefY6s/h8EVgaNkENC5fHlnrTnJl26TIunfPCmb3d76soDqaZ0kCUKvsLaxvuDK6JRASJhvNdn
Wye5DMBrdIcGOYCI/wXTP3oUcXcl/CrEWY0/PDLA9eE1yMeO7dYXQN5jHBJh/CMhyp9zgS3a+5ga
e9a+Ddd65EAkQibqGQFuyjauGy9N6DOtq6Q7aOKHYz26M+hsoOlE+w6NfP1+f1s0JQj2KHWzppvR
lQ3OUq+fvgtWomOmTjVws84UWFSXg5ORn1Wm2SEX/NLtB1QeWvug2WnDS7A5tDpGHHrcnIe8LXfj
xOYOVwVM37hDumqWobt0Qgcb/XrEPyotc4aOgDYeguIcQnbt5sd8NZ2FY1bjUEQHoAFgiaYIrsXG
LPKj/4Ww6ITtdgoXLQqG6BqpXzJ11w4gBaXzhM2P6gdLKuwtCpVfTztysLi+sQwDrSGiwj8mAKOA
j5LUOebczvP2FohX8MjFmsS5g5FZnq9lPyHA9o7Fm+2URe3yd3g+GeA493zZUSzHXWjooykaNOtf
Ny1oRJ1N4dxsPmk49EfnewWvGSHrRnhAj7EbZr6f0Kd+tzTX8SChQxlMmWwZDSpq1mGThEjy7M+v
wnlDZ4qKu62dC76rS9gt+vcbqN1oVnoUennF/Q2nsf7svM0FmpWVLYr24qQcmI49HceTQr3xb29c
FjGTE/IuUDi1BBMecBQry3l0kzJqVv3hPNxkoBgkc7L3r8PFyMc5B4WoFIlaBZzTwjrcpsxFnfD1
uCCahxtLMdGr6n32/CHTZEBgYpBlc8YeVvHFEyiDfRSr1nFIfRfQsij0FQU7nIOmlk2Z/CQYx3lA
sla6pcPYA2JuPBgyOvTA8kLWLjTNK5WUIxJkk5Em17uixJemtPod0jFhJD+kNZUKm23CmX9rFpml
FvtK7/uiNwYZMHkDpTGFtufZ3ff34KNKje8LeqXtXj0K/sj8AhLbwJpHw2/UpfPya+Js+q5CdSPe
BEEKncBwS6sxZnm/EawoxIvShIHbqu8m33YeNxRamDD/zWPQoHvJj7MpIaYkQlhXKvD1EkTKJ5Jf
PuH8R3qust1WkjCbXkd+5f00w/1aN5vsuGB/vM/7cF3dQ17AWB5Xvfoh5yoLStqCRnf9pkoNLC7I
yGCCXojsW7JGf0v6ShSaCmLQ4ryDr/GVaOXJcs7vW8chOtUSNdMk/YadOLgldvFebE5QcjUVLFPU
MgxZStSZjeAJsrNY5WXrxwMxh4VGPtSBVIp8gDFIYlQvImJcbve4yM7d2/KiABp/Od8WN9xLzJ1j
P4eU8qxg9bhuMzCLUjHRYUmkR88gPHRvnamET6zPc5gLM9+BSQNMsNEBZdAiaLIw0URJizhQOxJU
QTBwZb9mKbn+zbMqY0jq4fhrWKffmESMSsxgUl+HrV/S9yKIKIDlZoS0oR4UiuSiBBsD/SUxewqI
voa64ujE/STsZrIrzQ6Crj4ipnepd9EQ7VpzPFgNI0FQqNJ1sWDIlhPACoZ7DE+WSJtCTbWaEvDq
9pSEw80Xr4zWlH2Eque4ipAV2Qwey4/WXDlo4xQRhtc7ZomG9ovzoUGweIFAJaZfqShXvk3mQO96
JPocmkp9ZXgRMeR5SJ0vZgGCufGxPFtsxVf7xTJE7fXOAJl7r5oihaDFdAHhvIPAOhUEflQLrRPI
df7da7yEOtTZiqyezeF5xulGvpivO2WpQ+e9jVH32f52pKrF5L4N/DHhmV9QIZqFmQb6BkKMIqg7
MLhR1g9HAP9s4dHgbiH7Z6ARJO3mWAl714GmNrLK9c8hdI5wQFdu1yJyZoGIZfLH+nrp3wAECH00
Z4gRrsiVZv7/TMVsQrZrj7OzytJgRsqFR494rU/N5uvgeR/O+kQ3v/QOKzp0CSoYTYv8KgLzRoGt
O+u/k1E2dVPOEPCuZ2BqfUxPUf0g2JIJePq9LydX4/Qxf1t+WMgOPRF+e7b95GwsztUnmUYfdGfk
Jj1Vhpp1DqOMRkfaDApo1ZM3HDhzYFuzGyMf+qtMYXGfXCfvVBmr9pJmMzydo9S53k+avSr90EVd
U3QuA3HHxIMZwb3hJwwh7bAmduZp5otLKGqUJ7DgM+m47UtFtm9uUNGNh3XFyPYpOMhyHLoA9sxr
3NAA1XYvZ9IHMCN6EhNNJ4Y/yIEAZfWo/wSFyXWI0BdTT2DOfC/14Fw8t4b1u5/kWudj1uxQxJun
wq5Z1wdorisDTVhCwgx5l0ffmfj2XD4iMARtMTx33r/GU0UqK3kEBRJpl0zwiqcwiAR9y+bX71Is
h0gAj7ukjqVohT6DxDmOOWpghiCoC9jXIiuH3m5pfwuey+NdPgM4j35s8iql7KScGU3cP++PTqCm
1bO60RaQkLl/oQUSGexg6IwP3ek9Ok77ssqzoLkeaF69IjA/F5GUv1EPhFg9ryoBUwKgvy9cMWfb
L0G3GKXe9UCXZt/6BpZ9rIG+5Qfs7Y2OAbbVEJq6iuXospZ9GSD6lsGQzCSH+KprYWiweKoVN0Ig
zEOqHjCW6cj9XawElB52UdrISeJINuS9YnI7kg2uJWke8Mx4cJCzAsfIPKhHBt1tY+TgYymriZft
LZuEDrG0nYGCt1MHqoEJhNZjQjSOuFQIEoI1/gDXmlB5Qj19nY/ZoN5t1JiYdVSJPHWAKujrCMeT
r9qAXWfFT0aFx6lx5kA+V4NIKF1QFLtNEU9X0kFl9sQZwnfZxCKFqCPR+cEn7ekj4e70+GdoU7Qt
sFLHvx8vjIU4EklOmdCesAlwKTDIh1pJM6/T3WaG0w2Pf3t2FznOdrhJOS68Wsm7xovSAQnon9K2
jG1PB5raE3yvzI1ukDZjetayjv6daIYh04h6rsTPMZcHJ3/rCWCJjAw2ZPqNDkXemAP5OCh1x6iv
+vQmMbQs/dAb8ItQ6wB7Vy8PaqBayFNti3d9QQla2zEn27TuG9W59POHHtyP7EjwOPjNouUuZnCy
BgGb+1Aa1YSbBLRsM6vIPdyB6TrSsVW469AklKFdh3yKLb4hvIDb/7nbrEwCAIVslfC9Nii4UyRR
6pV5Yd/+L7CJ+adKKiRU92LmKYsy29nWeN7f3XiLBX80ysECkJWEF2IM2rN43NJ3IQtszYJqd64e
qPxG/JJbV74/6WsmpB5SLc1VXa3eLxFHSpAFNwXZ16OeEOkFN0OMAP4GhI2rq6nLoT/fwCHW5Q9W
pwBwTeXicoxozXdv9TkE12xWOob4NoFmlLBBS56qYgRPBYw65cuD6JkRk60RJ/Hu8G+uT1ldfWJM
tcxDn1sAQA5v7z00oX+Y3QGWFcJjNdj+dFs/Y+L1db1IW14gz2pDch+IoiOZ+otLFWb1WxSQUavq
yNmpknDil/vi6mpdY1YLolnMFpBJi6u55ETO7EaNas0BrvvOiPY6xbB7OGBKz3aQ20FBviz4331W
rWToxLvnwL6xMJZZX+FUrpAOoihIxOIqROJg4CV0/On6qPrZtMBIEeb4RRUJnKF7cWm0OXvQQRd1
fbLWz/MEoOsiRMFNEzEIDIS0X5Yiw5KbXMBR14tjjHtcW6Dvk3VTJSqH1A3ITt+7V9IEfMOBhN8m
AUpKOvERxElWGh0DhRKCMWuPfe0nUwBDn0Ky/U0BEvZoE19lOamOtt+CZ4JjQ/NpcmUY2s3CL4Bg
UNrEndWnNdTkLxWCtoFn6gFz+o0b2KRLR1Dgl0lq8MP6PXtxDjMHvqWSjAgN46fzaDlCPrC8JMOM
KDsaLr6WFOa4qz1oftGuVlajR8691Me6AdS33wE4yRIbA5DFX6pxK7rqE0ePe0hJpqFrvAHsvJdE
RPra/5VVHBLmdchp+MiCk/TqwZLX6rjmaWo8ne18bXYeGfNjJ3ctxDnN8KR5b2WP6YpFygirtZGE
mxRxQaJ6qLTb8w+SD4S87O3J8pJ7F7oe35sjNjO+DI50JEOBHPg2xz5rBXeB+NHZGgJl+2XAIZlP
YsYeaOMbEJCLDieM36XWopGFJiaX7BjbTySJ3cW+JXt2qOhwKq3nVYqqnRyR4r7DDw/FiCrr3PC7
NMfv1c0ffsvQYXgVDR4ka/5SLRShLbhM+cYLRnS7FeNhSd6HsOr98yRp2wB+wWepPsn8MGqRJrXi
+Cztrg5bJAdZDyRyQkMp7xxiG0TlkZ1/UbrpbvMzWrBsw9jLDKi3xs1ERWRUnA22aarpKh6tNpQm
rUj2E/flUwDAfp8KftINSpstGZrWyKBmS7KXNmitIaeYDEAE97ABz13RlxfZNycBI7kMfaNxA/rS
ehNPv7le2Zx10KJ2f5uJwbDEbYJ9f78ov3siwolTYI9+E6qSyLFIEWPHmBuuwkJ/SQmc6LzrCzOF
JLMy8a5yV+wi1VBTAjxE1aANzIbMDcxAruidtORBvV4eHKWj5yzIrCXEFuFbomY/ML7o61uEJqyK
vgW2ynamdsX46pNaOTXB7G9rdRruboL9skl+iAC9iEN1ZVfODSiCrHA4ukdFzeXWADHaJJjKmo6q
A3r5EUriAB47Wvnb1EfglkyW7JVHiFErRlkn/6FcYeQ7aUc0VnV1ltA2soUJhymARhBtWz1Qde7b
luGVk5A37PWUCwQAv+liCgkY1ZD/efuBsthKFVk2TPAwlJE6lDRO0BdZoSX+c+kYKhIAVint3IrW
HiTz0t6XbcU0ttZKnxWdk8ohzPYjeuM7U0Z4cYEeUwb91j2T7hZFKLe9lEHeqTBMpoSNenTVuPdw
BLzisLbhEBKQIV0/nGrxMkyvjGcEsDvSI+kgzt9SqUA0cAXH8typeNxbkvYICQOvdtaOmSG4Uu5a
cVo3TtMFQpd1cXTHK94IzBBafHRkXgzF/Q82N18x4xzHSz+4H/AWeC73VpceWE2QTP++jsfKURsl
anhzVCpM03joJu5i+mUuISCZlX3FMciKkdwFN75Kx7LDDH4bCqj6dYltDjYd4wwWUSJv8v5/5Tz6
wod8NsQsV2yoxwA38zwLMhp3MR5gzcuRZlqvdvayVyx4WPGFQpChhhK7IkKnjYr2gFOZtQXGLVrd
5K7D8AnhOl1UNLjp5lpocw/EVJ22pMvd3Lp47UJZog6CwOtMJpfQyc1Le5jSSVGtL2qgX+q488Kg
K5aVNH1dUOCWQLrefTXp1fPgvnm/Y/T7mmWL+ww5Xp963ONbJ8Zc8EtzQAOzPbCc4CNjlSNJJV9/
w0xj01cE8Wl/H9Nx8qXYQz9CNKhewdGA+Uv5MI7h7PooSR5iAt+f5JeuVZVx+VLRZYhuaTkevlRY
n0GAAYHbln6JgO+8zyy7aCD8m2PvOfGJ4XMxVAqcVMewBwysnKkBkWixHAuoyZWa5Bx8mpDrcYua
/9xirRtQQCsiPDwx/d18V3fR/9/BmKabhDEIQ5Fh+xB5P7wg8udm7mJexaiEK0ZT9xlC1XTVEfDi
gU502xP02VKBwh/jTSYtkQVz6SNmlTm+JGjn3yMqOzTp06FvkBkKbfnquV9xmGVEJsP5b8/EhD/Y
EY7K5SY7UZELiCOEIT5Z76WKDCeZvddxMXuDZsY7Hk1w7/xG07JlqkRNqDGGhg5fBxV4TCkdsSgt
Fn8We1u9mVNLpqVH0WUDCBC0kulLrXgqKPc2qUZcZbGZh8Z/vHLZprkJuye5pvHpFXkRX99YBUsT
Go4OSDOeAnu9HWa/651ejJf94d4kPnszuXqlgWnwHjPJZyUGIEuW4J2ZD9C5Ok5QciBTNoTbTcMJ
a3K2CbTJ3X0SVzSbz37VODQM/YZijMn83VrK+zHvbThfyAzvazpCJYJvJ3487lrZcY1UkD0VmcoE
+KlCnFdbrUPU9+xY8SxhlSNFME0aqdSKnPyP/m/d3Gq7dkER8GTFwjD4KwRMGDcnQSFskJ8Anq8k
LKhcIp1sTM9G43cNF5gqte5WSZuCNpJZRkK4KCc/dTe6rkmtbC8xlSGQzcJPwnLvC686uWGtp2C/
JnRxm/TQpYaxFaTSwdJxwtoQeYRhirAM9goht1MTEhkAbhpmflAX3uGhlEtRz5nLh5Pq49nIemmS
dx5glMDAyXt5FFKyF4gcrhT6tT0nQfnv/OBzb3zDa3yYAkYokM8kZhThzeCkdichwov1jIyMlMbn
beFg+eJlF8bVxKYLi1iB6kgZ0gmlUNkpdyenHByCRiT+yTicPicb8tUJiFMlCzwsvPmzyRYBfTRR
zr+cN2hIPgbsrr4/qKu3Yz1cbJ6/J+sdDJ2Is8HsFWLOidLH9NPR/N+B/lJWknD/Q5vBLNhqjPIr
LeGPlKDLJ3BTzl3eY8woL7dKc2nNZLV67Hujqvwu6ZSBBkOjd8MCKoNCWD9dblc5fF1yX1GC4qGn
SjnQC8cVTttcPMAHl4lBWuOsBleZTO0zvvm/JI4VjHIJxwM49D2H9SM9fpoO2zgpwLG4bbTglBpJ
5MpfndSm7V1quqvaZuBWAOttfNuRQTqPuIEg1f5Qu2VRiuKqALs6ZYCNTfpopsb22J39p4c8ewmu
XGF/Io5dkRc2einL7J1CRMQr8MV8e54LyTFIClDkp5tglSHRssDEWtaL4Jb38L3Ho0P65ksETJWx
TFXGVLLrH8K15lfd3ZSFmfUUDBYa/AfI42VN+KZHOyCK5rhSOOs98YjqeWhFOTB8z/jL5c4piOud
AVL06FsNI+V8X3Mpw8sIZjb8AcU+o1hWn7Ymfs6tX6ND8IGCYngnSoaA8bQ212fUXmNTk4tWfhfG
fHJa3f1xPkujCZRyInD5ftM6jCuvc0XoazlWAQAmS8+Z7YvNyKJuieG7vUwdlx8VbGGVeoQOpadJ
kIa786LQYc9SoEb+i/05HL3mrEtAu94hrQB0tA1Cc9ROHTZDy0l6Scew6ViNCWQXbUaRYMOZIQfA
4MQE09tzxRZfJTlnP3GSDxpLQabG6lmkpF+EOy5ork9TfMoD0Y8+wAYvFVD+gqDE8ZfqaPNw+5JV
dEy/jKg6igFGfWzD21W3mGGFZQjnDMV3LzSC6MIZKzBr3ZzrXuL4cNKo+sjoguG8idliJR/Ezsqw
ylbuRRiRPdKHNTBeWmRASi0l6qxXR5HehS8mxPchWRKvBpWrDkp/y+ha+MJfX3yO5d8QdV4rHSLx
Pk5yM8Pa8PpoPY1RWXHVfmCHMNbguzw01aeMnNGa6V+bXqqWP37dD9Po4adqxpikj93ZdecaMur9
YDUSFNhxd5rkD0UZPgMYyj1Dnt6WQRdd4zVYKEkDLQ7CwXpPR2Uw94JvPFVMY2/cObnoYHVwrS7q
QHu8nvp/ah1O+M2jtoTSk7/EJU4Z97c17hbyT2SLYJAodId2yQ8QyHJOcwIOX06G+kkdUNC0/jbU
vVKJ5SiY7t71epyTFOhjUnEU5IGEQEA/hYyCiyEQphdmSv97rTUScOHYypWErF4VgVYGZSY0NY1N
QViPx65wp4Rq+phiPNJTEn2kzKlJ8z6cCc7d++q0BkHBr3kC24f/He1fgQeiQvVUkDzKjsz9cub0
rEOCycBvQTyqXo0YxuitYdHO1V5cLC9b2z5Gb2M/Oo8nJ6KHjE/5bOg6i4oZ4JrVOhEVnwuYNes6
luo6kp2ymmrVA5RMZBO48bOy7kekjzaChpXEEgrhd9iqa6YjmHWLRSkM01GUPe6j5O7w9duZpS7E
NZQ229hEswJL5cVcc40Wrg4B5pUmAXvXI5WBw3ShLF/307YkDHkj3zVIIVKC4CRqAutUY+WgkvR6
IRq6vySWm3VwZ3i/w7oeZIUGN6macq2c0kkJe+uDbIbaXQUa28EYCZPUYBjGAi5Dad5rPthOQnfs
7jSnTgXzE4idNbC0clr7Ag+M0kOgYEDc4d+WKpjcp0RZYoADMXiKndoHMTYDnTX/PHD1u035GhWU
z1Jb5CzRRhTdb+11T6s3xcisKQ7NoLFbUd/dLkbz3u1gEpvwJLwm2kuY0A5lZvrwv0H91EpRtVZa
mJoUPlaOJzvaEsI1fYaLhKdRUyWRgV6YHIKVAETNNOezLxg1dhxmvjFTQDkZ8/tuzOJKPUaK/GHw
c2RDs2uXYVCccm7CoL1M+7p7EuovtoLz2Og9SawNK9lk5ePuxaAz8xVlrkI6NLA+VuED5gr5eNq5
tcu3L6+PGXsUcFb9fc/qBUV73Dk+6F/jtN6TK9pShiOKBPRVHfCYQ7yFECx4n6g428ajJd0Y9iGP
8J21bipuRozrvfy1MYMYlFV21gSPKIytVZkrCrJHgzIVT1q6iLF/jubfdOPPU/bl2oh0kjGMrXIS
Sn6DLD0SfN1rwl+HQcPIXSuslgAl1wkpGFnFDlp5HHZCQGBMbKqXk/kYAJvGLfbK3etzF0zYskTJ
F3V+dC1USkmVDPVCNpqAa6l4Wg5KJ22Y+tpY4sgAfzE34JNznDpBUknowkSP/G6s4r4/YaAVgRiJ
I0Z7lwd0/GwkZwSe9c1zISW5Wr0kvBJAk9GGBkavWTBdPBcyPcevkUFDfIwTJMpRIGkNsnTvqzYT
B3wI3soLuYod9LMD34QAq6QmWpZzNiOZebrcPx+1VjNSy98hNx4eYl4tQxpLVGG0VljsArKsHuPw
kSG1Hu7RJ31WvRLbF/c6Urrsnnzqkt4FI1uiHAuTia0tIvmdeyLVsH0DwdyvGmQNpaB3kQYHV1B0
mMcKCye4wkdkZc3c2kOms0KwhOmSR0u9AqzdqqAaJlhF1nUkVuDgXheeHLX4C+WtnkEoS/QpqR6i
Iz/Opwl4776MyLNozgpY6795UeWm/O6/woZ55pm780EDe6VR5cLkymYo+S+gAq0yiYUUBySKZFjO
PKl/kqEkEyXJ4Vxpm3d2+UXmNFtyOkrhbT11K7FR5SPQepV+sfOGfvm2rNvecxFNB4DQFiaJ8uQA
PXDTy7vuCoV5RcyNMfmdpp56J1uoAc7y4/VC/vohMk+cB8TTXJNxb5hHpkCukShCnNUBlQYJXquk
D6+OGMOCgHSYSpDclc1LY8TL+iwi88LZg9KVHVQXum+Da+OKBFCGxBIgIATZhBAE45TISlT/90i3
yTKyebu23Rzj5nkNIew2NUzvwcdU7ku0Ubg31uY17w+iS0Uqr34m367PKZyihqf5SS7IKIjYp+89
YGkGAMsVI5xZ2Fi9u87RFAOcxLuiuJcFrjRm1IyqZuJDF3NZnKqiJ2T+0y6imduIAJSzWgWR2sHV
ozzHweV/KkMFG+DDzftqrJ2KM0vL6YWmOOZoDg8fCFLIDFFM3Dh76hcxWSefSivqmQdj7LN1cZK0
ltKs8tZQdYyjrR5JUnvR7Oh3MSHLdtZMKMDaFqYyaDEP1VIaOdswf6CC6NTUEPJ9h2cPoznXchkM
agJnZpxOyJgwuoo3GqQMn8uB+PTc+fQT98gnwMl1IgYtoeOw3015uYrghMlU62xkN4bHy6Qsz0BL
74FCZ2/1aNl5UGJUABdYM09jjf/tcfRfxCHTpaUMrw2BWr+EZbWqKafPtL/cssFEfFJs5HRRuX20
//2sHenjTbCYRHm9tM0vGI/yMBQf4waX7IbX/x0PmEf81UcLBSOTqvREczQ1Z+GD9jpzJhc9Gm6K
n2q4G1Oy3KiTaFnumCi6k8pAm12JMMJLjtf8FN5PQwV86ZZkOJ3sRgz0prXH15Y6lB1YP12HNW21
NIsFNGyGBAGRw+inSY4u7qeiYNC7hRN5Sak5uih4jTJ2iRr2sHkW6TC1RghJ3uaWEy0P9EINDnxe
Clmcipk5fAS3xITF+6/I5ynKo46/FX6fQf9xIRiqqVZ75//3vA7UsneRHgsWPIvphsllnU7UmWk1
GJOQsZhcvFDZF8GFLrGZrBmCFdU0P/IUIO77oW8eOLbV9q2DZEF7qYhpLQ3AaqVvFyPtwkGv9k6U
P9sh54BpMYu6qC40KMOX/ICm5UJnT0HfcIrWPM3O3miMnioWu8EA9fkuVnaFMKmvyT3ooST7eNlk
EKkcovdtKBZH86HtRs5D+Rafdan/AH9xytjTCnBjPoQ+9zFLu3hFLZYZgMQH/7YIr0rYOpFXeHFt
LPNYLqu0KvltXTe64EOAMmjCpeVS20Yz9Rr8d6DDVPbD2vMDkIpuDEavWwi6cHmHb08H/dN+LdOR
qlQCurjeEq9/+gCR7WFfDr+yBBudBLgc/CIRN38K3dOxKlVBREOWSMzAJWH3Gwty1Vq2SnA5KL64
y2M9UF7DGyx80v7ULIxFJii5sl7IMFmtf9po0WHandKy9nhL88wDP1HEJv5oehGJ3qGcZLncSj4s
QErYhK9jqg2qVFxksNxGirWN9xmJ6Nn6/3PnL6lSCqZkaXok1KBhCweOfwUiI75pjf2EnRVNoRv8
c+JIA4tuyTjr0em/qv9YoMB0EljARG+fkZrkdcS9rPhOSK5VnediYSX1E0VOea4aMJ2k9sCm70b4
/YvGir2MB/WDuiUSZG9P3sD7XRnzYwNQ/rhlHRcv2Y19IC+DrrODxq+rtddWqkt7lhDxXMPJHbra
xbGD2ignHiTG4XHFALecdJk3VjtZaIiVKmiSM1m1RHr4+TO8Ateq33kyP0TXNj18O4BV7+CFiygh
rrrHxXmHdtQ6qnP5EtUVft3txMw54fcTlayt/FHN/bR+2TqSAyojm/Q2UhpgWO5n7g8hIo5228pb
N0so9u1RnFoXWr4Op7ge3qkxVAqI/G8S2v7LZ3jDMAngRBmodoHkicDpJ8hX0eB3XeCFai5Zr+uY
uTAeqOpJeP7MslaQ48V+hRnr30N/D9tRrZ6dQlEEj7P00VvXInbWCksE7h48A3fNzQpS9q+5P6Cx
Z77Cikvnp3nx6ND5ZjW5fDGHPr2ULC24KFx5b/X4Y4xxnvPtr4ZY0gUH9e7j36eTXVe/593cVoVK
R0aODkT564nRUCNTX+8+gYLJbYS5R4sYv39o2sTxjHgqtgg/cfFhmyFgmEVfzef69DGPhm07b8yR
SH4iUGBkdFj0Jjo6z1eFNeTPEwYycwrBPHsme9vcTI0e3okUNnO06FynAZMBHOPVz7oTrjl+q8dX
3lQY5li+VS1Tf1IKLypDjw9VB5gyE415V9FeDHze6GN8QsBa1VYAhpzD6cmHfzQjpZqVeT5ox9SO
10Y0ZSA9quDnxS7Ho0G60np7Wa02Ha0CqEqyzM3GJgnbPJEKIRi+JAvrkk0iPTjThz8jYr4T6Vuj
v3NmGu19BtD6jJ/Q6Hin8GyvwcAgECwPomdKtONkVHeQeDi6LlxJdyUj2S3rpklZ8sfR8/lm571V
RuAxp2OnQS6BhwkIGtXT7zYpenCZcvFLYApN66rq6+thpjbQ/8HGm6XX7HTrupuTIJ3QoLbZuVb4
xf/pfbnt78aYpB7AYmotzOvfqc84peyMAmHLg+2OXGXXGmuS9G668UUl28KHAZVotMznDeilQLtX
axpSgHB1tU3UMVd1AR2dQ1aVnVSzUqiCKbmDlyjkhYvYtU5XLnYC3hTS9EfY1MUDYrGPVViBCWIb
HWvuHEa/g6CkKcT668Ie1NBCyR50hFg+ZgAAYg9gxcWnsa0vc/3037YVYpFgAhaKeSmVIXZzmhvZ
tpSrtW/GCwK3oEgUChzMIPrFCi+WtJYserKxzLDt8khGxW+lfl6ld90KNbSdsNAbZkJLr6gBOloc
IxqVl1r7GTRt9MGrt4ir8D+aFX5zIr4cHiGIcL4tBxJ8Awk+ewlnQ6ab4oxgw9lA7Pr/5pLfQzQJ
0XHoF3llB58U07IJHlT+WeRKBYvU3GK3dhP1uSITek0sAJlXwC/L4QdR00KS3MjMTmvBmzKkLZPM
P9735ySE+8lEFggti1riIleHcx3B/cQwC3+mc8rMg6dabH0XGV3ZWpRJ/oQ6zOHLUrpsCINs9IZw
3wu9OomuGzvuEagQA2RuU88CjGAgITSFLBr83rGTCJYbJP7qUBWu4c5qywddgDQYGuwwMRDkBlZg
MyWv+wgBNuHaBsrIyLF5hc3qyYLMQt/4U81E3F73uytid78kL4GeboXY4pQLexEbs7b5NhBrkqWg
0/JZJPJLGh+0IEwS/sgeyl1UkI7PsccBCAi8WHPi2l1dvX1P0eNiJBp52GKMoJkaThJF4qGo9pxL
VnV8wKtA1m7Wc1IigHTbnmwlXTpIXyoBFnF7K/OyZpAYpNNS812aFwGadCjTbcZGzViEcaGQKvvO
pRhtE2xIs+wnZChVX/lAijJ9O+2QwY+hP2xX9JY3BtGNuevclyq6PCruJW6oaWWXmysRulsq1/vH
47eWAEBA69Z57/zXX66qLImrLBW9aDQq28e3v1ErTEtyRE7boVCv5ZYW/ScOquvtkfB/DbaPO7gs
uwHRoHcao2VX3Yvd34K3fNDoT5/klyiolMg0+4gfVbRK/ebB0HGoZZwGX+pBbwO7oUp5vMUn8TI5
So4uNjj5asrUa9bMxyjJ0lph7EARGAUD5i9Y3Gdg6OtUgjd4V6SO26dSNq83NozUNTmC0Vl+V2/V
B2lHZ3j8Z//09vOMztDL9GnZLtVICeJvoo5CRwtIS/dohjl63f1VN/pbIgy9/lUAbH+lD6cCvXrt
pqKt8Ci6ewX4q3rIsF6W280R5qWH4Gvf2e+9Cr8qhAMuKlbcKOMfHLlnpF0lghk1hRTj3UkslH87
CXBeusQKeStvCs/+WOLrQ9U+iAjTpvsQ0mOL3PXUsr/LQ8vNAkszCPv1cX/ePLluykMXr9sIi37I
4CPfIHc0g4G5LHGDglnMmyeT2GcLzpOEPz4qUz4AwELtqWs5wYdygf54xS4FGgkMNYtjVK8Xm6+N
rhlAVCKvXBLX6jEzNRvYqm3wgsVKzysnplALwffo0uIeTehXHrGTxhhBZcZ/TKRMi5FnvafhcP6p
8BrQ6xpgKvmiCSed9VIdLN4afe/9XyGcucctbrtm05UMQPhFbsi5fHDTVAUWSF6xxCGEQBMHv10O
6jmitqV52/BbFpu0ecVpLnOtLInDwX3ymRTymD1eR6nwQ3VmScQvHNCxNcfodcbAUjRWu1Cd0Hqd
B46ex4SQWYGa3+r7NPONnGDjJSxkbb5FUx8BR1vJd9Yz0YeN2vx1H3PRmB/0UwKzXA7D2Z6sxcUT
J7IfyDkz6TWaDgwiffwfo9ARA8njFTTm4wFhU5+AqG0IZ2i7t8zp32x4o7F9/yvb6f2yVzCTiE8K
tP4WiV/NrId2VVTYpj+IgfTwzoGOAXxVuBodDpiyRJzCZV2mX4dxGvGKobgmODcqyyoSRluZVoGv
fsNQrwORusH+J5bh5hJHT375A822Wug/y/2moCPHoEF8j/UbWyO81xACUMYGUF+fcFre3Z+0o82w
TokXWUhZQS8UOFcbZlapaVmvfaa2gk3G7K2WVF3ZFtxcV0LkDJUgAz2qi+9A1DjldQCijHJQ5/WD
0Y86bRYjg7X7fzGJy+SVZpTRTJSo4tlfEVNo0iKWX8fTo0SRNToD/qQY07h0Ia1D4DtYbFHq0PXQ
AoGGabJkPGQy9vwjpts2oBdXtnJyYOhWKAIMT/bli9GgDA1mJPgXgnOVmkPx4w6PpI6ax/AIbgw0
AZ9E/mDs0eq5mhfOMHwDQlmftfCSg7U4X0oy2l+7orldmbY8qBzmof2TRum28YVGRA5TI9Mb3jYe
tympXIG2mGH8aR+j+xP/dvf4sgnMjUQMrYKplQuyQL0U5xmA+p4/qVFxoTGOQHyW+Y0hakORewUC
QI46wZUwYKyM3CegGG7jGV4x3dxn3Rfk+dDFieiNmTHiwJRCyRddl3/CthyvE8D5TXyFqPbo1jNL
9ftuzzoFNJOVX5ojJ4ifYz1zDOBQzjNk+1b7ppSEjHAn3ARMk7Y82anSfN/GCBVLJHkak1JZIgjx
9K42YpfsHgYzIKmiuux3tU/3mWE50XX05UoRLvYBGYQ6pwM4A7h4a5YVhVJJddBpx7GMxl9nMOjk
A1Vo+Vic6vzpINgtyqqRaPJAwOmO2JGacb3aJLfPiHEWYXzUod9BFFaLTJ6nROSF+wvU/Fz9xR80
egxLNe+7W40Mjh2t59O85KlblYbwcek8gqwOT50S/uDV2M3InXB9yn3BkGK6QthdhE+P+xT+C+s4
GJsM+k7RvLogxUUY7x6MVvl4zXuJppPhbt7kSkBb0Av2xgybeLj3C100mex5VsqODaMVJbeNSQlN
SDmc3P1Ur2ACOsUfh3zt/rGqSv4QPtX0qCQNPvm+fZVq+60rMAevwLkyIKZAkuWv2lY1M5NKAS/D
IErPl1sFffpvdrMRrfXbfNm/eG3QYyFdZ7PA27SQeiKzp8xAKd9et2CSt/83OC1u17Zd2cnLNt/I
H6YtjMlfflHsqqeJeBS0iIR5yVUrogkfesdfT5QN8CiEIqUkh7sHaD53hNtSbSBU6/vX5mn13EFu
WoFd+GwC8g9nmQ+j7+0j8JIbqE1/ijq1BSS9TS5gCo3LHfMWhuxD8UOb3wdK7r2txTfjxTibagd/
2xcDx5MJ210Yivn9WYocWc3u4W0iOa3Jdln4mWMTpBmOqxrCJAM0eRO0ITxW0mIcDshImf6+kurB
HJ/eNeiywhPU5Aef0KD6YqsGY5U9c1KKCxgzPh8QUpmldl9MHY3ha6oGsv9OOq1eq+Ma9OHvnFa0
w7uqz/bRj624nBxp0C040esDF+PAAabe44CjqUaH7rcc/FzbjGYFk+6+uDmjoDUPkZ5VmwhcwoyE
GYH6wRigFV3qVHs8sBdkzp5IeHiGse0Wo1pxkASp7xqfsYKX/W2SYIbKk3iqLBzUdoTBXfL+egNU
wf+5VcAGDLCbUKne2k17WqWxEdY58CuX4VBguNEuRXT0cpi507pR4vJjAvVQP5odDsa2r8BZD055
UsHszU6KbE1a40UYDz4CsR1j5P1pzZrwd/86lnM4yPPfJdsVptc+1AJWs6tsDjMTIfo0muAsQURi
RK+Hjico7hxtSDhqr71Xlo7Ll/G9k/Ls8axwvawPJMCnntKkD84u28bfw5YrvWbsa8LnLgf8SFd8
blJ1SaAyfcnAFEdLYaPrDean9rFKl0cJkOuZ+TsHHuzRqGz8Holdo0QQYn6He9ienEeEH25ckyK3
g7keudvwTKwErmKqdKiGSCEmXMft+FvZXTShwy2NkSCwIb6m5mRBUs6aYjxTrnZhD6b5wUeuqyva
OpjXgebmHD38EBD9gXxuBPK4cR8JQNJ9VwxJtqZeSdLEWH3zZo3krlGy6l3T8cj8M1kzTNohJr/i
165lrK/iCH09L1csvHDFigoeeZx3Mah4m76X94uzdUdAeLhPLs4zXf1kQ2BmxTDtjevRF5X/nRl3
V3R8+WrXCbL+nK5CG9JmUff2XdDK1hbbVUpQRwhLVXSkQCtAqiqT/QlRifYecBTYd8zTf07Jhkjo
9hLer5SPKraakjGOpX+Q/TnHLNXhr+CQQoOzKXChnTDgl+8bsvN78r4Jb/bjrmLdVU4jQ0nNQoIj
y4kKKBuJqe6wxIQPNF5vEQpnv1aZ9RdzDR7EuPN8WuFKYG9phDoC8KZ8J/BxWlDslD8FjSJbcH4O
wvOOYnpjnp8niZcimXTRZIxPI1AubBZIy7+N1DIBlVAwY/FX/bjE9eOqxM2fflZ2KEpZib8/lZIh
pRe+x1MZmiAbeIt3Rxptkay3Dp8GR9HsbrAc36aUXMm68OcXjny/LyOS2Hm8VbOhlj8T7stRj1hx
cQxGvnjH3rwtK2xcACjG64I3yzeRpieKsqYqIYId9LsR6gQU2t4nuiVzx/ZxPJCw/17VFQkGaLOS
wB23GKaei17BM9fUCrkT5HctY3JpIk5crTfpM5GRK2K9xUcdOHFUOfZAFvrDVGWCPa5ObnxG1dWH
B1/oPjpID9kXVAjgoAm3IoFFLGQlve5/lVeBboL3JzUcDH6Do2zmNf+dTezMjeHcKMCKOr/ktWGp
qSq1qjuxXwbQ1ium6D4i0TFvIPHtQjz9PbEaPTF/3o+r1C5bTubc7IR2yZxlg+mt+pwoeRkvpb7u
eceI4u5jrJwSFNJE1deg7OL5Xc726T0eQ+depsuBYdl1lnBThN5AFgM4GfdYy0npThyxCYFErUAs
OmfeJo6flqzQJooePTiH5rbYKwiirQPIcEIS9Xv/nMEJOonxmdwRZinETc+luJn4hHApsVDwikCk
7rOkhjzCsUYt1fJ+AiBu5sUguHAmyQTzF0E8YSv6ROLc5J9m2OHqm0rbwim2aCERSLaerBCp5eDo
iL7kKMjJzlToZ2JEuijSOaNvViYdCkiSiltsVD+cCHcaQwvllmFqECr2PdUdeCcZXeycxbBsk0lE
+s4wvuJG/9Jt7QX3XjGKEfpBGFj455GDw+dWGoVI45REoSdxZojd3HX29IP+wvtR06T2isnovV7i
YyfKN6XJm+KflReMsPxmuIFzG4Rn6oAX2/H5fdH5RPrarJRisncsqhFgUwHM2jNk2VruKpOVIOtg
RN4QyMOtwijniNPF5cKDbuxb+7V+Hqv6q4kTP07wCVr76hzkQya7/NWnBEXwlTWzrTnrLYk5GJ1J
hGL9eH/nyE3aNWg8Kly+oVr5So8NYPOfn9puDTrhr/1WnJxcQ0INpgih4s7NnBB+xIJQYtgx2VFo
VnOu47aweNXdRLY8J52jkrZZqhQKUWCYsJ8I0/45RNr4avSckQpjPq//IWRngFQQdFrQKIGfWvXD
H53qCaNFk8v5tUyCcAdEGDfguUbpQWmjUFqPKTNk+OIdjub17OepF6QHf/nGPVZnfKpyHklcxi0y
yaXV2xYQgRIq7W5x8GmJlZRfwoNs8MiV6qKuvJKv9J83Mc3igtMqekaF2pv6TPHhWUYHhj/j8tm2
kpVtRcZdOPnXzcu0Beh+8FgiUqI45fhVt2uf5GIW+2Cz3aC9s4KPvTp/TkC1L1H914NztPm2LSYL
4phtcYtLNFmh37U4dvZ++yuX8vOyoSyp57HP2PtcYl0CZ6a+5f9rpeUh1h/KHvhx13PIrhOUsmI3
tEtaUdv7xPaxR+jQbwIyQbCM/63c+hgN8Ha8sJUNLhESajZ7lFYFzpoLBdCdhePs/eHrw+wsMReX
IoGrwEvWH6z9QHO7tjjTEGLnb25KoYJktSXMgJUx3KK9JcAdH+HFYgtt2M59JDV846dcwDlYVmZn
53LDsRzMCaafbDMbnAT9M1e7PsDYEGfwUapea2oejNRa5B3VnxpfbI/rSq2O4S5Eww4MYF8WujCj
qG1k4Obqr31443v13lfTGtB/mohd+83Jl/RSzS2c8tZ0vsinVMGVOp8pkrcnOCPn2t1zFbYDXtPr
er1wLsEkocuoKC6I3MpN8/kclCpckwcFKW6pzDoMOKXHxW0ItbtMOELImUPANvcHeJ8vlYyJs7As
G55biZShfh9of1Dajdlf28zFd1YnYkKAl/sQofl//JxWZoSH2pl4PGnfjxxxSmPvQ71CSHq3I4av
5U5kExihy/A/eB1Hkob/Soo87EXyxVjnAnPevof+QaaXF8fA5X27UuNzRYFHX9WHVV4lXbXmDE4U
uJ3QMxgf04wj4l1zwpJhhPVK9/Zedve8DkbgzWYvwPbGJFzyzqxXwmjnnF02CXL+XbjYn3+D9TWd
pjwSz2K6Lr59zeG6HVQMnLGgwqyhowJtcb4qATXWva/pMMx+ZB5gT2i2HkWTgT5eovpwxcl/EsH0
tGcibKL+M53+2TzKEg0aUTJeGPaB/7pBYjotaZuPAPC3SIpJklcRW+vzFC89Geb1VB49UQ7RN966
BKqZzGKNaDaIhtwC3GpIeWIhddwfFDwACvA2KVnjqxdyEDNy64rTyT52AE+g28LFmCVZHqk/VPB7
E0FOEhPAh7Hzh0hVduYqAIfi27CkpR10bIcC67Pquid/Mm2jA8I/lYkV7WczrfrL59cAlDoih2bE
ZxfXc8hag7ZCOS0Uk5QjeMEvspSWI/31bBWSUrfrutkHtggOs/eM1y+hi36rhkguyC52fg0ATIcH
2IpTOeaKlxO9WE2HN4dOsFnrxmr9GG5sV4EgxxQv1Of4YodbtI2H4xInyKDcSermKJnUwonWjWUb
s5Y12dGhcNBNh1RRprWQJuJe1VVdXnpg8iyd3M6s7fNR5U5dl8stD1Rpvs2P8mTHiovaMi6MlnK5
0NaiKyzihPhcwFKY1hOQyp3ChkPu/Wd0jBgc7eYo2qg802NTPALoV8Djw2MkGekgdYZqYfxGhuKR
HoDhcC8rbK2hqozW+lJKJ7LdgOeqfY+bMs6ceHHDGfG47BCa6J8F2dU9Jqe9L+a7yZDFgeiNxnA4
2+BTUnvaONa5mVbux4jpc+A+JYTe/qD5MnHc3T8KdI+1cGR75qBtKIALAVMO0hpVPEbAcF6CuFUQ
es31OpSU+rAqEHy5IBQBMInYRnetd/HntKQXDEKkKlrgXieUVTHR8WCBvQYYqyyeOT7MtQuCh2VN
YCBbYEPbevNSIUnbUfm+KMPWdZqHb8EVaMVr7FBnuNWhHvC2CdJPimpQCcN3uTdvWkTVEVNNn7Ik
IoROp0BnZGtfCL27nOLWvRJgDKckfYo+7HJPca4p5xfc7dar5gWHwBNk9by7fLVUabRow39ZuPks
LSWdcVpbLl5X1a/kxLhjFphD06/5GstznQj4P7GQDd1LmUVipw2yllRA04lyAgN+RdANI6rNw1BS
AqYDn7mmEksl3UgKbQETt1nbNi3ZIUE2QIAOYYiccBGwXbWgc2lk2y4yFCnM5XYadqX9AEhL1tYu
IkJdpBr3B7KQogi2gCYKEbHUyJm0wkG8f2hDsDCfJhRfrfLqP/J5+gjRj4//mSpWixOcHrELwGYM
Pv7fZ+FTMakLsCq5jZxmLPlULahqDw6t+GnzPRbisLgLu7yiIWotP9oWKZx7B1dc7q90poFGKz/a
L70pYtoVImg6ad4MhTlq68o+c6svghoUi3/pfAqq5rzAUCOpYm3b4GkXI2G92xmu3vh2Xn9YZ24+
5mYSS/5gFb2PatXl9UcfjP/R2gxYFSPdpWtKUd1wLnBhszPY3r1m8y9dizIpEnifX8DGvJRLZyk1
cnMsybw1/jIo7CKzGzzgTtvC8TI4DDKRCRz4rCcI28cqNC3KUaaMe+qDoQMuq8SfspIHReZyjmSY
C6eeNxI7UKJJ9YILVMVJa3jv8IzvxKV1HFjfT+291Qbb/8NCHLcEwGAi7n7nWJpoiBWLklpKtzxy
pbj9gMZRP8qshAnxTsAv7S5hcx34FI/ow5Y0zrs3x1/Lb52tYzEbbCGWVxmNosvjCabk7769/ayX
L8xxfY8zEdDU/6VcAeWXrDubaoYxyiUPXv3wsL225/gmzwUc6aOetMcQSEranWVFnmJrWTl3FQv4
Mq+YxAy25jYq+OeHpw+mAx3ueeaijK/YKwuTcSrOPgXGbRPSdQEEFI/kzrj0G12FepNEGSwHC97M
OzBfFVlDweA+Dj+Li9nF1o0qCfbMeboJOxq6dC52w+0JlUKxnuE/rgYEfeztn17OqZDj7ocUZ6hs
osufFVaRVJrzq/tWErGeCDrt8O47Ry68UXHGznQ4VypadTq2RFt9iIPx2prmOwDetkEiOd9uySJY
w4utouu0+OGamgVt1gJAMgY9ZZ/wJM8TvDnPAC4U9r7q6bX/ox9V0jOT5zuk6ggCiew771d8vlni
12Gi6QvZOYHH5+qp0nMrSEi4JkBVsvOnnwK7Zd9+3Lz9QvH0dlLI7SeMASxhtFKnTwJNINXAjoXz
7EtbSXAEIStJRL1dR4c3idTqWNVTr+ZJgolkte3rqBEC+MY4gfTqUAw5tsBbS5sWxPkrDKkVrWf/
kJi87ngiAaFBL3viEHp1MWk6E2jl84TISSpg4/3EDx+FIMOlJa8nkqFifF0M40TpOloKGKA7INPn
1Z43cnjz9iWz5//HsxNub8tT1dVcjyYBwAJ44v22Te/gc6iwbJm7+7U/HxQ6hjgw1KovElZTqde1
xtogwLsTxs6HRMOEwlNafr/luChUUZZkb6aSsmCFt8CXfP6MsVGdZL81mY+SKY9P6qzbboC/vo75
fFvcwE8JkBEkbkDvXFbzOBx81yQx0fQvgZxj/mCZbO0cIKyNMHxJS0L9rC12bhIT/JmlHEBba2Gu
SAggOhuwjPPM+kwjIMeciiKy53Xb+CbcwC+oUYOEBNicJfmebqGuikVhPSN0lK464YXbQB6fw7rz
I7i0OCdM4+uMrXyuvx7ILk4EKG77707eYZC33BBz4/OUE1IO+C2FNFvLDnstk5oVA2PwVLXoORqZ
7W1aMGJuNVSufRVY/gaAHiXKNhQKk3JuKat/3yiv6954lPi5piwr1KOwrXu19MVq9w+wArINqRBT
7QJvUbTCdhX1mXU3r7XEDGzVWynZDMM8eaLokq+xe8uziDOGDAEYVz9/t6Dxbf1Odk1o+rk9xWcT
/+Xgj6yV7806F8FgDEv1c3yuhtyHabyQ7BEVpHWFbAz6TfIuHhbHOYlDcdtwg82LqtxFgty9cnYJ
JKlw2vS8iQsy698DGt8wp81HuTtG2pWCnQG8M9PT3qXDSxX6TJ2T4Qw0xYpcMb8Zwy4UEMjka3Hw
DSuOV/n0jjUaG92A503WZ4FPHeCFUDyz13+YC7fCVL6q2ia5kvkxEdhhmWKyXUHjM+Uwf/psuBfK
RU74xayqeddw9QlsPFX+tT51HS85dqzB0Uck9IKWnh22hxBO769glbnNelBB/hLxP33ZiArIB+kg
875Lw5ft97brvD2WEKMqDDpMZ48Ja6e5nPcJJpbk16cb931k80B9wSdvn48m3+DwPLrfM6c8uQma
oUry/6FHyM5bVmmRxpqIBcXX6gQbfWQoWvQCE+LoJTzXCFlXDb7SBlaXPkHxyy/z6qdFTTPiIxM7
iaSPg1aLnhQ+TEXDT1QzDDHHshYHm7v/A5vqIQNrp2Zk7Zw3cOPaUaCDnXtUVkkW2Xx83oBBj4EZ
sCrE8akgJEKOZy3nEa3C2tbzpZ6BpQvdDTBnJWxWGx2e0YiWxPTAlgY1mJh7dpc0x38KXyClQOV4
6PEHb+IQBdej4hNByg5dY/gL2n2X1gY62l1VSG5wtCXrZGJnbcQxUOF15UIjOR99JFZySM0UAECw
yy/IyFhxV6MhvCJCtzn/IfuSyY5Z9Ukwr2xV5sW7tonCjh7PI818QX5VWWX8EOjZ9llu13/GmsLk
a0EuPrLQmo15uZh5FAgoY2sVtVn0PetNgP3pKDP2sN0OF9zLHh1jFKpJTSBvbr/xRkcJLs1wysTe
FlPphOxF0AmMfq6O2oSZKNT+7kPUECGZBl8GTAIv0Yc6Y9mtlvg+5uc9nPc68y31/5ZvjQt35Hd1
ZbgtZVAmHP5sut1OK5UDC4C+7SJyPonOsXad0oPyQGauh9Ohb1cnlIdq7nXyq9LioPctDSgVCgdT
Nm1zL1LNqhp1/4+g9sN6WQmfyucUG0MiWYJKhu5wdzHWD6pJ3WC0ADF8/F0pc//Rnw7Bku76f6m8
VVK4R5BT+uje2T8yKDBmSTyAdoJWSE84HsMZBOjpV+YeYFWCupduptv5k/9xQGQxVoZhHRAjgwhV
Ep0+pBa78V8r9NMpRzwtmMDC2o55pvUtNWGJVg4zG1LX5PIp6A5rz6yhGcvNXjmNUSPqzdT9MZp2
ZNQUa5GBfQEFelhm01OwufyWH1v3gcgPIabE6L785NFMiaBlDhjT5VlKq5GS5fS+IsYry0AEC34N
i4PTVoGR/HKN8dBeW/Y74WVXX1duoESAC5AUKm77ERJ6ovoCSudiiJv199DQo7Fjz33fUW1hDXOj
+D+V6lEn8htfY5I0bb21yfu9O4QQDHBQH8xhNee87qkhHGZGl3YrWU+euOL/AkF1/rodPFFMAo7W
ETR/Q0SWc0sjDjvbLvmT/cR/IoJoI+S8aqYKbNF/v2+vhnUaGNUPxTdedXeKs6eda9pHrNjHZ0oB
dNl65rlLc2vIDDYp12R6NsA2DVzDJhzRtxEuWrOebJnjBygCMLq/OC8uvS7EBMzGh4QEWqdrgxO6
pAm8RJQcwbVsfQ719mqPV0s1vp+Xn/9zPLanTmFsyhvi0vaezy/AEx1HM/jpa/FJNJKsVD/reaeH
YEZnio4mTJlte0w5K1mWol0dzvU3/0WQYwI+uFu1y7U/ksif43bYItUeA4jR2QvR8McRJtThT0dZ
HodbSUYvePTQPVhOny/Z4oelTMbmtiv4A1cuUJrvjPIjVWN+ghkfOOR4ne35MKjZ3uc9akuI94+o
hR//vHRQDG/OAObdn/ew9gIOOyYa+F1/aWP7L89HseUOQDv0vpIFTTvHlL6reK4ML8OEFtxyhN+R
SRjdulQMv+0JUGETzikT0Baz/mqTsvTCvIYR5WsHrn2CL9i3eC0IFsI9lLll3rwEIrCv6s60keZi
yIYFmMT4Vq9qf1289F9qh2Jf6elBby9yRs32C1PInpUnzQm1gLZIeIm3pjOc6Vg5CL1QYwxDdHJ0
y6dWZoGCGYNfX1yb/qKK4iuvsp8+rgAKtRlbQs/UGsHf6BorTv+9ojRkWKqoKK+tyxRAsmuqfM/i
M4t89q7qubHGqNyc4cAUKzJxSIw7WyIcIfsbkRTCx9elJrCA+xZzNLN6iZlM0TbjPahUzOazgY0b
tGhs886XkmhIS6CoidG4VOheMie+kwoKyNJkxAU7O2kvBpImIOF7OwgsDCqwrlrZFtG6iSdY+iLR
7BIyIuFC/uMg4IvfJRL0Lc9l4AWGjOt5nzHGpxKTbfgKaDSus3eqKcRMKUWFtZNg7+UG5edyCgzv
3SB0oNZBRCufdV2HYR1mQZKyr7BLtrQr0ckY/Jas9qC/UCWnmbyNpuyFs2vGoxInoSAdqOuNRdu5
XltOAJzM1gW54eEV23D6LnlZqOxitPKUGb7Utu8WdrpenFON6B+61AhHYD2HxUWi85zUUbLrOX3h
zFi1skOShSFtOLlgudk1GDWo7gpBr5KeRd8Pwssn6/ZvGRG3qeYPTJSGEpD0+KYp5jZQvSosBYeX
MGZKhcCEAlnJZtMlHfeI1jW0iNDGtQOSANG8UPuE+EyU2EhfrMP/3PSJGyOm7M+Ln+HvJJfq/Sp5
V5dW6u6/UTjNPA58eSomrcjO73JSytZZ4s42gOGaGfGj+aohaFW+gCSJ7ZVYmWu4j5niDTVDq7Jo
+732gMO8OFGtzRhSJnCUid/0nckMoTedUaV5r/qgnAVw0VvSzRnt47XGLhi/Dd26BgC4JZ/6SU3T
aC+Oa2e3gv2uACbxZHQ2LiE4CO2YGG5/cpvpiJ1vfTKy/Oc5370qgujpMY2TDJgEtyxaFcw1HTFv
3RBiBO0MGRR11JKaSvSZepKGGFZ+njEMwwZobcprbt4R1Ml9ylnTsJtszcwGCZ4MSY19fSwEWUFW
h09zODhpmIPs020a1uxayXyQJQKNVLqAoX+KnGs79E0z69kdX0miB/0DeYvB3HrfR0ag7AHbAIIu
9FsiLuYz+UZ4EhYi19U62nzTJbbmExG3WLgHnNmoiGGM5CbwvfG2+xm6sv1pvA5wyPSrm25XGLw7
vxb6MyZ+Sh+5Xfby+vTQAC8zWP2rW4OAJZdn6SyPPS2XsjglnFWHjrj3jOgwfvBCRqbXRHmiRuZT
cr8khpLDjVQgkqxr0kouuitLQuDJ1gvSA/SWf2b0eeZ+rKs81WzuexZ5weH7Er3jG8/mtA7FqR3e
OxvaIamaqpKrYkkP9sLZG501V8APpQQ67GWPxnaujPSqHlccwHSKpUtxHjImj30S3G5Wahdag1o8
oebNllW194Pw1Uqk4NdpSu0y+Xext7fTYPqbz2fvwIeGv0xv88uAV2sH83Z1qJxkVpFAIC0AoghJ
aHA2pP6N39lfQ6DnFaxNO2/46vxGfSVU8hSglqFl3V5/R4+d7/XiSDKE0L1i2Jxxn6TkAQYiWvE6
BSede+zdPUpBPTSOzm/8/NuujYOCaOYEXc1SFC1PsA29oVJUtNlIJsZRTDlcyaHM+lBuxhzdjptt
WZK/NT9kkqJyDltinJ0bZNJaEZevBUd31G1hXf5mHbxTS3or/a8j+9qSQXSg60SZttfGDuakNwJJ
H47CjpJ4TLCVCVI7EGURtjRuPLsUcuhq5SQA8yDsoU7FTZ8eLoGJO/3TbzCMzf49BrBNDZ0G7biK
mIjFA3ZH7VhNGyXbDr50bsyrujyRK3qmouerP10eutNP5pFrzDsz+uyajQMJd5OHwFJlVP1SA4fP
5r/PrZEt5X4ihxkqfr4zDNrH9qC3Z5w/AeGbtMCh+k/K1nC3m8Y769EB7GKVg/x5pdzCVZHo6I4S
LVLCADjuvATjBiAUz3R8uMhxDGRbCD6BhmUq++YLNAfwawwPlgPJ8YZqCC7xDGBhF598K0rg85LX
URLpCWZWMH29g7/i8FP6itXg6u87ecNRezRfUViDBs15Y+SNg3kuNcryL3eEhGBNY+TCk1O16Qdv
AO66wDzMXcOiHi9JMMpeKLPo8ikFgG/SSbzP27pXznbQyv2xUj5qEcHPaYPKg+5WUe+v2rE1BW1s
vywfFeXpJpVwaegaJhBHyK/1PhVx74jFsTqatLy515Mmz8XwdrxR+jbre8/FYj362oPCwnY2a0RS
T5jGkVTWnc3tXdEeS2pxxgCyeuRNY5op+99a+qv6VvIG/XzeAop6HxyL7GEj1Unzaq9bzQpdLOjy
ANYsrmMkisTFWM8o34CwMnElH8W9xQREKhK6LSUCBRVSCqvOjN+HT5VPLcYS7E4JEkDtINJ5P/Zh
uCtiGP7oray4W4Rz7eM70nyVe3jE8aZUvjZwjB0vF6a5nkz70UidYAJgfyqfwxYP3EYqKHu10qNt
JMyEBTmFOMoCMnhi/gxd9gdzjBjS0Gdcd/Kz74NhpACH3s0B1U0zSQ7Zq7gKwe7C9+q7NtI+Beku
1hGDIBM2lbCN96jj0Jo8UuQ+V+p1Kj5sNaV5KKvfviaV7rLqhHr8+O43VKMqGyGt4Q0RFrMlaiYm
qb73s0wOE3HF8Xv6UVsbRHDXb7L3ffrIIasRLIVqWC45LtfYF34pC93dyrQCCUeZx302uiBbtELV
etCDFgtJnIJnbwUo+WJ3asIzfyv/6C5QaVOgpeqq4JoVnbmiVCiWESTvrHF0OlMp5fv8U3dWP6BB
KbW3wPmQmTnimuntlVQ2vnVCsSVEt8znMOb9nhcyjGOFSQrELQRUvW/B4QSleQPgdNb2QLOyS8Og
SSlWBX0I827E2E5SlFbbhbTmDj68w/YkYH1JeMaXxZ6SSnP3MPuxEac1Wj8+Ks0MpeD+3HHyqRaE
oNFlwPuNBj1wE7iGm2rTeXTM6FXnNItx4WoiZF96K1+9twPnGDLp6/ILKWMQdjG6llqe1rtbWwFi
MCdF8ZRFKnr2FqBZ3srV1fwHzgbevWBZ5Co2WCZ2F5WJp2F6weyFJTn/qi9ZCtvIYpFY0I9Xw3eE
2A4XNbx4baxOpgEDgIwEQr8cELajnpETJOHTETUyVHNUaQY+kRqaaiu3DVjcbb+BxIZ1YXCQj+DO
x5Y3Aw4q1r3gNCCwJccmJUmklQRv7ov7Mf4pHdEQLFOl5g7cCuR6TCPM/B8r9yBvR1hX03qJgthI
6kqLkJJvQE7Q+bhfye8jeN+NfMv3cYOrFNsQOoRCKVwcCLCEjIxGtBWNH55+UOQra/uLi6JI3mbW
m2X1cOcTwyQ9TOWN1bWeF/H4eci65c0o/RDcDetWo0ZtQismt16L7f5fc+aRM+v05yUpa8ILwhaJ
XpJiFWJlh2Drymb7NuNbVgWJ3b98kayksZfOjP1BNBK8Y+TUjv7X32kkffb+QbWDbBPMOXNTo7Oa
dZJMi7Uop2ybQ2EwOA4ZRrUz8h89Vb/9msZpuH/3P8K4Ja0On8szpc1qWG4kYDWWQbHp2O78e9sl
RW5Lyi1eMNeNLjlruDjMaWFZzt/opPQjyL2taaiisxXCjarVr2Ble48kX8zYJUCFgUPeM1jYgx20
iwWOGFtjepuhy9t/jYv5tns+EHDScWwIrnQrn8FzLAW+cIeAFgJ5X3NhTezewmoMGAUquBEoSYke
tec9z7ILqU9zzGD4QotKQRjVGu/vQb1HOq9DJclOf/2YM/TmOJoUFGrHoKaP8jMCwE8sDcDvD1SY
Wy5bEBXeNncYHTOpnJNbPMcssNp+JaMxzUl3xMPNtYzqKBFDnuMTBz1hr303E1DfrkjQay7CzwHP
Lgn7+mRdnk6633yWn5vYoUETZiVau8G50ea20ncJXLCQGDJz6ozX6/r3UV9O3dVroPiqpQyS/F+1
o8C2mEJjmtUkaxzzwHehNyUp4Ob/3nCUFYgmR/XcnnX8YGFg6JPtVyfdjUMs/REiAKKOoEAB9LIL
rOQN+Xm0ueMIMAHR0VIh1IvqxHJfyGo2ySeg1z+yAh8NRPUHdXz/G+adTs4MWEbMBjob7dbrgc4N
GfzBZN/PFFeF7jKdvJkQctXnzNZhAN/0DavRD/A5WY0HVr/q1J6DNer513bcA7a0pNXeamtvY+RZ
ljyNNIa4yOZ9ilflQjO6y8krwK+DhEGJ6tyLnWtRaqJWGvFcHbJ/pYGqIq7+7pzr5hjODtAnkSBY
98LfphOWxv20UGd+Js1cksvekz+ORn4kyJzPDvzT6ep48vrllpBui/Ukbg5zrN5Ii9Y90oR41/RN
ngT/zgAyRy+GfLG4n/b0l556oGPUy/chZDsnFcQhEKqTHPOwnZ5nOfRkB+JuOsBGVELlG4pxE6j7
VI9xm+eeqmVaUYUKjSGA77y9piOoxpBxo9nNYdWsy0AGcUZUNeklKTjsIvwgHCMAVAYlJwJrzJu0
I88eJtEvxQy1l31xB2nC3U0Lsg4q/eD5dhrqBCF8KnQOil+91Y6qwtZHS4kt4ZnbZrLpSpiAccMK
SHOPfHavWRxxo6ZIWwdTMbB8Sdu8qSZUInriNs+aUu3payrF90msPfOKoiivaObajQ1f6IjwWS/7
9Ow0h8ZlLJ4p7zhKAMfIXzTtDmFUURNPZUvfWUi3/BhpraVPKIryYlRUgnL1liK+6BgaNCY+pH1I
TMrskfhmByc1poZzx5Y2jCNrO+ckUhS+BAvPypzwtQ+JGPmhe4/+f/6NbMqIgOeW59ZeQbYItQsy
Tvzx/C7TqvPlTL/kRMLsiJSr1T2r+f5yUUlzNYL6RdOVf6bLx6bN54QdrcxHao/83FOw/LvR6VMH
pXSNKV94zxQRMATPv2e+cMSprwza358Kn1iNLOPcE/IDVLaac/kEgiGZ80lHNjKdMM/XX5kxIEZJ
u2rtakFx2YCjtKMONIzo2J+ann96MzME7pkmBS7U+GMvpdNQHvq2kKXOozUZJ7x5mwWVnM106bkj
EtWkgMGao/sdHSL3rSoK3UvHoIBmrzzczFWX5B/Bv6+ttpPNl0IGomSbsXnHEs1cJeQ3Ikoy9Qhh
o3Jh+f+D5nJEIMuDEewaakWfv/RLeQPJxwIrMhWWTYqFq7mJzEQjKQzKNJ7R/IXzsxDmsGfgjESf
JL6CfFrLwt2K/a9QVdBkukz/y1LGaOxbXLfc7u2WeJuKMo5neHueNcGWkPuzTofuCQWL62XVeLcE
LwmxdQp7ogXEcXTzklp4cb3kgyWK0Fk6uXBnUTc1sLiKEBloMqt9w5jtC8LKqAPFxbkPi31S4lL3
VpYE718dArivnznpaRNEoTnckMfPC0pz82QvFSKFPKm9oq/6BTcpuYZhDrkya1A2DeuMfuJ6gD8l
CJfKXUxoDD7uSBkLFVoQuwMXV7UWsaMYY4HPD1jWBRwqvJDP3umPjKkW+hEO4h/tsPB5na1HyDMB
PGux9b+muqN3JoT7nRCBqP/gSPq3seIU5ISAo7lgNbS/VaYv4AneVG6b+f4qt5b97eJpIlxm/FCL
j9j1a0NLr8ud/UVgtWiR4GAqm1lxcMtPQo26yqj1/YelNXdP0qZiQYTlqZDhMvI41I2BWPFMH+h4
MSgCzNPFs5tR6Hdn/eIDDbLMnwwfEA7qaR+DhBJJHqxIfaZii+R8XaV6k6yv9sQVxXfocLHN55eK
X1yPrR37lvBsor4oGBhtnEfiQPun8DnqaZlsOOuF6SjHyPr7yr7I3A6KuUd4g4ezAuNj1L/XxSPR
aNtt0FZkPsMpCxSZoa6IvtuRPhm1hXm9sIWhAI+df5LHP+SC7DP1zd6Lmb8k0fcEL6qIG7asixeU
vs6A4WkePxoEN6UcWuZRtKJ/5ASFDxUsd7hQv7UDNoMFW1ey0A94BEoeYyMNohGfz+X+78QNTgRF
bG0MdSFcDi2oy8BDI/UoOwLTLb9dd8fnX2rPz1nami5JxR6aYYqS8Eb/1xfD+nntcLfeXC2v1HJp
gtszsP9Xa0812uj8jGfDr16Fji3B/1qY/vAh3CiDH98b4Z5+25IW0t1GGY1MDZ/hHSSeqlh/5nyO
4VQv9psAJD6bNztAZHPxjECJwBjXKkA+MLk7rJwZ1JYTVZj6N27mXh5Hc16NhuLB775S624Uh8GV
vtTnJR0gvCTHOz4KU549O7UM+lo5K3AuxVS72cDbMPcLnIPREz6Pe5Bscg+V34zlOmdGUiEKxbWB
qUA1iQZFQ/+qkJV7Mb00vPHifQF1jQwwHb6LGMxY3QvVyoCP26CDXTyTB0aYgZufZLPMQ+irLceq
MaIBZnjsWUXSQUxkxgnE8NAefeQqS4GOEGkJmg2itt6COx5c1j6J+lAZk5u/ab6By7uyQt56McC+
UEhXBPoMwLn+eCD3USrPtgegjb9UoWHTDj7r0XIBvhheHEpDGrGNhqwzXvSom8NHGa3T841gXtPN
nBEMT1sECp+6gQn6HSenzizHjjIJh8uCy3de/DfQDftzM+BCl6vmisyj7PZhndWVIvrN/nD2bA6F
sRCOe/ESsGIKxWDJZNtEht1LVYxFwhGJ6pyrPobpsaLchKstX2YVPfArn090YIGxnFdc+FfMUr/u
4fWfFJsN2PXSpFboZoF5icrck3s+hqm2pAu5vhfofA/cnjJqEGV4b3fAHvuz7ujTVjWomUQC/mAH
7XnCQLeRkVcQ6ZX9lAE2xFavAvW8qY1eOIqEL+4Ppju0KSW4GMJ/AdVCW/NDgPMZSzcqUgdSaX0G
2eyiO7k4i5H55alQJ+4FPkO4hryERT9Ab2UCM3kQPkgQthORVxmcBmTr/31LLE1DHGN+cULEqiHa
VsAgQWZAxxlvEc+pRGYuqBA4okolz31Ldplpsz6rowY9GT/ua+S96dY3SJlmp8E5ZLa0NjYslc16
ZPNLzVlLHYw4D9tqWpZowX5bPCH2qXZCfKp+oaDONgLkmRv9Ts7l5sAzgpa0+zcm9M4FaGzrtTk6
A/z4aDvp2aEchHKLnsALxwevyWLCONJDlM+8p5dpIJFR1BVx8XnTSnDzYiLZwhyMvX9iC1XqZUG8
6Bxly4vFyp8F5ujf0q2ah1xvl55SYoZ+bHrnB4yf5JePpC/17DKuq/5JA+II3weWJqroMXE6W+ku
iFpZKriRuwYa9QjJbkBagVbD4PeXlhK1obH/BkLyuyi28xx5XyKU0SYS/Z+yMdYHTcwNe3ObHxRk
EtE5OAVy3SbyVgUiIvaVAvRSgBNYGvd4TN4ZLmbjDgAhCmawUYXOvbm9qhty/tUfkpDuveZ9L/NZ
GXnLzdqqoE1nziZC2ZUuTQWP69qnGMLFW7itVSfWRMkXYXIgYMv5XGr8eDbDJuDNwKxomjd2W838
nXB+ejMwO/v/clyz5kLi912YCR9Y8A+dLuJu6DloG829UU8BIo1o9nSaq/2qpOYOuKTMBLNXEA2H
l6KUvgFUJaOQMs9xlcwsuTPK1UeHiekxFMXrGw93BCKJ3LsYnOWUOj1qlDwBiBcTkvEAfvd6OYTg
D22kqn4pQwtlpieLFw8SL5bGPVflbJQdUm0b3XIMrU1Had/+A7Cj9f+oeconiatCUnhiinTsfCDD
lTkfHONjYrqmJOs5f+SGm7fP38k9OCxhA0ElPSx2PLv262wgxqbXdRXgKLqWejCItgUCeBj0Uf2z
F7LEu8mEET/M87XkQx4Z/cpMSUQQbSELxr/ct5CEGQYqPatYR7RBeWLVlR6+Lull+YsgKtjyvL/s
sL4zAqoh26aIBq1UnamqU2iOOGrhF8tDD4CmUdvo/Mwh79h8Uk2Tn5KmZGx644wEeA9fufeN3rKN
6Q5bDoueNFX+lGhYrxsgVhIBKUA/onQqgIIpDGQlEPjj+sGO0aWaDD53Ev4F9DxF+kCwG1GaMZyG
HjRJXjOMdV/pWsxT7ZrdnysodYam9XB9V6KVSjtqdSFqrw6i9e4W66VkiwiwSaam2HkEFcOR2cVG
cbRyg76CkbcwBVVDqnPqn4lf91Z1sneH0a5hsaC78tjmGD4rePRxqq43AU01uI8KdLtsyy2N+qCE
t+dVFG6GXGjvdR2ZhomYAM0C/F819VvWQQFdcoRvv42x3jnNRYMEmeRP0nPFlqi4D1hHcuYEB+CR
FedHyaAIPMzih3Nr3rAve31KlGQcZ3yrvcx6PVmKI1Dm14eed2YV0veU6P8DZbZursqOEcK7WGjn
yy4eTvKT9zQHzoni6jXzwHnF+iBr1Ejcgqq0N4ME2P1/5oVacrmxXrNs0D2buI6Nd9gpaLCzpoqy
Tl2GHbYPkDaX1G9Jnb8ytLinkUiJcogTh3Vn42N58Occ44AkbSpNWxHzOCut+PT5AVq/DKcTOt1N
yia3WLNFeBL+MbVMQAr5vY2kYfaHMVyUcUKIWK8u9R1/6j7rHFmZIznbm+IgDM43gwDxjgf+1g/0
o3hOHbvwLCRfA+CEI8mW2Q9a8vRAMr2eCvHdq5ih5ZspQgF5OrfXZMvY/8arr883xgzEPyohuS19
ar/3dsTYgswj0FiGLbytF5SddQhmd9KctfCldHhx23sEmOL1Ywg5biywfqFxIcs+sRSsVtbC+QQ7
4U7hhFDks07Y61R6zzSHNdX2vmYzspySQCMJUz6MdUb2FMZkmjY6tUjlp9z2LHU8KaVDZ2LCOTxD
oPU+rZLFJj9/Amd2q9yxFY5PG5NtoGHtCP6GOlEXyyy1ggj/RIIySZ2YZlL1DmMALoxW2e7nvQNC
qE92PygJhld+D8F5MIcjH86wqVA1I6tXayo/fzt7RuvogUQ56q6AvgkNLPV/MCsw9lQtj2vH0HKp
YIdScB4Qs8O4CjcuRBw/EqOkin/TvIzm28GQsGeXOXTLTEYo3IhzQ2henXd/7erh+g+YJykElf0T
JAxGyMTldVtKaQEfL5dLNbC3+LDmyZwBBksVRBsl7KqTa3hlKD9dl2bqdEZgW7BwWby0QPf5Flg8
InIyw9n5mjblII5wcf/YokUVTOJuTgoTiiiOKCeQbu+Q4i5mebd5NzGyv1JXMH/7Ljcj+6sxL4H7
ARwiTWrnpI4Jk15EBq+Z6Hwy0HVX9Q/PIB33xGH5XdZjOFiPQa2dy95v8cMvg0hK0xd4wCSa6s8g
wxptiqOnX2qZyCtknMIQA7UtL/DIb+ot369MSNgbqucZZmK3b1Vgw9MVJW78+i77YF35gyPZgsUW
nEeWuwrVPSnbFjTD6yzQtW4k3kotaQ6u47B/ui3wyfmOWUA1NmnQ85BnSJfPslyL6PHtvMtzeLAv
cWFxLLNNKTa2PMqw9I0RV6nUT0fVzB3z61AoFpr0mMhpGQjIO0HLZeqP3MyDUGu+EICrjcZTHe5d
b1pVBrHwTqNBjdiSbtqkVCN+juQ7A6u+vrfqiKLxM7dOOtLFpI7ANSx8JnLFmQs5D7QuKX+9RuFF
2Bsmf0JBqE8KAeScS0hNasTWS8Kx0JJll0/fNzeFVvYhTEi5rxq8ph5bjGObZjeoBYc5yxX5sEyo
YN8M1aaEPODcOg/U1ZOYlg8q/lIChFzpFyxRUjMFsZwFdArQgamOe1KLPCCYr60cIEsdayWkG2t6
8RuACbu1DChxw/ifJDRzQm76lJa1kIqhJatAU+2Rgu6YLbwGm/wD44j1uzQ+u1tj+b/05h7mF6B0
KHBvVNRXK/+1VbVD6Hw4IT0hHRaDAJ8n4kuQhc/984nY/pCOENWrhYlqHboMLsFrrqewAVK8M0aK
V5UfeyP7iprTJ3n4Lv78XUGvwCEOEFxaW3YrhS3ui592iZ/hkm/gnZOiXYu7ZUP0BQ06qhYhpAod
+gZSjrBBGdC69zbrUfLURIuez7DI8CwFx8p/joQqs7CeTTz/zBSDByw0Rwjh+unwnKz4NZZaheq/
qG+zczfg7qRcP1PI4lYyGaqSZySBrgXr3tv5r+OnaxMEEyW6P7Mf6Ff6/cYLNVw5JQdc0pIPi9dh
8GDiTkoJfjKuzNJdxyyi7eanYTFjWTFeTiuScSLhIQ7gt8/tn3rdfxXBNMhzvYLRRvY2mcWLmGXh
UX5CB721TmC4kKDSXPYh932Sn84dWQa56iHKuGQ7V27lNrFDmJVX+tK1ERu+o10tZMzTZbPpjGmI
MYKvQnFpfGNS/qNN13ZKfeCUaw/R9pzqEhSz+zCM22GJJ7w04Fu/AEODpFbPvXvWtjzoj63cgtuC
Irgjf4U085HccWOmwL/rKHEn+PybcqwxOxDa1d1DToH1oPN/e4oS27yP3fadPsLD6NEuJ/2rWTsq
etvn7nedQF+xHQ2OPDK8zwk31HcVw0mrFckIdOiFIkI4RnluQshIh0P389h0JuU4t2Ju9lazdgtD
PT0vj94NtoyiytSEM9I0PfeyzTES6LiSf7xl9T7Bxy3sMEA+XgBF3tRbSYeU+80mmpHABJFsndFC
etbVwjr+ildqMZw0x64+bQdRr+I2dHzhLGdPgckMAAdf0m7fNsJ4RyzDCfCl8MxmSJtaA6gLkSY8
Z7IpLsKjQX9j0i/+djOAE1YeejR7K+CZEtjDzJjfRLDhUSxk1nTGcG4oHcZ2ATiaEeBW5GMrQgi/
69GVXwItGotiESYqlqa33sgRzmbaj70A0joPiiBOqTkvlltLYX33Z1xlvBfJe5NC3QfAEwnvsyfx
wo2oYGRGPwd8IqoLd+VaquFj0GovN9/lz/EEBwZfT+DYRvg/LN/ESwBT1WPwVAzn50Il2dlq+wR5
1vO6HAxUBhjT54LqYL8J70nprqG6f7Uwc7Qg3FUhK227lYMqdev7rBxjVyL8XCcMEe1fMA1RnpJI
FMIkpsMLlReBHKmQE52LhDrWMG5rWnlLaQbv5DW00RbUs5diWz4+3Z7lAVO7wewu461qbt+w0KI8
jWv4b/2sd2J+lSfxQVJ61Y7cVM2LmKgYSTD1aLs48gGyxKAM5xbNcJmV4pvo9l4NIEUpyvYuW9K6
mgnwP8HhmqtQ5b4CfBI2WuSASbPhk5f9KUcfy+lgp+vuG7SBwM+lmxBaYMnwxnAI4qFkTIR2cd9B
mJEROGoUrZB0C3VKp1DplpkafsjJJbu5414LUAaPCTA8mLM9n2aDuf1Bb5avAPU7OIjG3Cylrgdk
2oImwdaBGPhGXGssmBtGokiUPok4PM95QzlJDudfgu0dfuPbv0l8OHc1BqANHZdGV6IuewUqMJoe
cPFBxHSu8T62Ib5A6VZHkAv21tF7wERg5PztuMWcz+ugowjna/Cc6vLEr3GSTSLlI7yQq77bbm7b
N7U7NwAaujghyVeme+dDZNHykrOGpIQ4tqK2ZSmvS4Jw5Fbm5kAySDyOJpcQWBoH+1+eihuK0WgH
gZaFDwvtPzb+waQzAHl/kidE6dYcCCfRe6uMhYGtnyAsjG1AxssIMIvdAQB6y9w3THyvu9k1PaZG
IgqMhglNH2Z5zBoYncHJG1g6/oxG/Ztv6i1Pnnh3fsT30jdlcLQEAPQLWfZKAEshx/Z9McO1GEkJ
2kRRQkDJuMKECVy/du+hLsJpE3JVGQn4td23n8ip2j0dW83avSuTWDy4HxS1Zza4/ACv2Pt6V5zy
HrhBUDjUbfJF0lfU5K1XAX/QRNwlpU9jQ/oAcVBtHY752aJRqHiLuPsBCb3OTqU5VhoatdHNlaOm
5sI6gi8v+F3GZHNVSDeSMLYpD0SNV7Txewxb4HlUfW1FjOdMcL7yWF7F9Y73cy0NDVo0gtLPIGkM
MJEFYyoo1wPsjFZ1g8wJc28cGEQOIkm/NQbc9XIfE7wqmWJuWpxWWKUpV5dYMSVt0+0UnvxDJgez
FLojfn9n99ni/5tVx5Y+ZyynaGnbrxkL15YE44RQ5MdSn4cW+S3NgCyFs3bl5FLyFdfGhH0j0NiH
eW4Rnsx6Cp+g5R5cEOkXxwKaCNOr9LdHhxmcInrtlmEU4XYqFUpGDgd55ppoonZuQbTXEfMpaqSa
E7CWO+uZ0SQPsSG3D9LwlmgM5kjf66p3I6DwT1IHCytxdK07YmU98IGz0wBOGPskorZRI8Rd9jiX
3rYgEgkIytM3BYIXHepuYaKvLMP//Lea5kGvrxQxZSG4AA8nU/7NYl3W67PEvjdbuimPnccS4W4O
plv8coC4phyTqE/T9w9i9Xk6fIYl1R931aquSHWDlUmlhxpGVacKqT+/TfVOmjoNeV5fSNDK3c5Q
fYXNVFQJk115HyWXlAfnjj8ft14eHKLPOkLBpBU1Sc1dWoa1Gl7s6F+lrjiEtk8yvXJXanbLTQi+
yJipSNQJvZnH9BIYkKmPTQIIKjMA/YUrB/IcREayVmt0y0QtxPrTcdsB5XdMsa5l8klQ5DAP0gJv
LqRw2b0/YuyD1ThC1p/QsXyYOXimSA4cO85pBqHXsANAHCwj7OM/p5j8RrFs/5Heqs9Mw3SdvRv3
cI6dfr0RC1kFvgVpdGIi7/hRXA1d65AzO0haJJUH/uXFqZuvAOASNBg8zGmcSfpX4VA6aXtmbSqQ
Cgk00vFOMFUWNcAmDeKBgYrg8zLEo4BVDrDwrLRSbjw67L9FuRpaQMhk48K8LQm0Ln4Pg+CDRwQy
JJ9qXoVHJVC/F9x0kUtzCdy8sSNWWgzLy5QaSMS1rrP7xinCc7fV3+5B/hjbMdNaP6IwXViIt4Wh
fJiYVqXdRDC21M4SyBXoAd/8Aqoi3w2rQCSP5CbhR6QFAIkq441ppb/KXOk1dGr4bRdcXxAbVvS0
ZRoFKFaXuYh+IraWgIe9sTAcb/xI8sdgHFUpUGs014xR4VWaUUdcyWm2ru7en5Au6rYWJZNrAto1
1Y+0b/8RUrm8ZTMIzbRPBvLXW9sK8SdOVq+hsFkpYdamgl4aohW4XZ9HGASxYMWNSi64n2CcTh+G
b1PEvqc8UFwn23JyJCHwg7ujJH6vVztYU1HXHIKLBYd2BB3lxIeV8FPLN9YLK2KS5+HltsdxbneZ
jOzRjIyJOtXGua2lLZvDXK7BATiylLXMe8Mbp3e5G4hdYpHOmJxDla/zFtrwcrp061t4y9C9YMKt
+XkbPXB+OMRzDDwltX+iDXY0dYpFQ37o8r+oZ5wPBI+YVFJJNG5js5arhrZLsUOAN+3hkkzf/7f+
Vy2anYNVw0a2uY3XyJJkpXVt5fVsqTdJDrs23Ue+YOqH7leajPx1gLKWB+euf4VpkK9trXNbN3xn
ltBhLrOszmTUUto1Ozita1KXySpdOYuEhmfN4wHdtuDW6Vi7zVU1RzexeRU1izFX9voXohqzUyoG
JnMNWQDzCa4THXZNh/XzlG/5vCGftTXTndAVp6/8jskCIi73Rg4tgAdP9r4wcKPtZ2SykLio8jtQ
pxuBXnrCqwqj1Eni1tkg/7BTd06zymOEa2i3Hj0V2hQ3TiO2ptvMdsqUYpX+CTEkNlyGlD7mrrdE
ea537t7BfhTmfLwurMFnLWX3btYhDfV8j+ymm/zHdNwtew/AHzZFhrQ4s3gwukqtMWbVzJrzQ/08
Xq313bVxTqcOFXscdeLHZDVk6Kzo38zRAw7DoB5D8y8ttqHaitTvRY6/rA35p7XOBzrp41Syr3FH
85o8ZxXsecyI7yaSjoslYvfilveWOtO60N2elOQYa807zCM2A9yqd3lDM+IsxSPaW6WHnDcwYWt2
Xppl/9K1obJ2BonEgtDpmP8uegh7IB6w1END7xFXk+lzDEgMjFHxF+Nrw4WU+AItLZLaqSMnxkr+
RSjjWbonv6WR8/PUYnNaSaqN34N9Vll+geAJeBGBtr2mT+PihcYkh0Oum87Xu4yCpMcdEjhCDyvU
bPLps0OfKB33ooUYEf1LzXkMsu9dmAWulXlvGK9fH7aD6MIMx1bMNLmVgmetwDDxD5f6KTD+clyd
5kOqGjekn7i6iH87taOS5lut0Q2XmBkBeKxXtENPHUloKQhnFV54qdoSXYYWheIhYh3I4FzE/Kgq
TP/uPtptCJLqGdPxBO6fS6MLWfTIPSkmxOXgKLULbd0G2T3ApwQKe6gIoHR8125m9sEGOumR4eFw
B2xRqxKSTRXVQEAbSMq/6cBO6Wz7mArbArrOGBJj+1N17U4zIPm0LksZVja8dIPfp+FBODsRbcx9
O13+xpvndsbTISRJU9LJa9fsW1Ax57P2CIeG8x77mqWnRamdBScyU5OnN+jk3qJTUpP68pQsVWXu
iGlV/daesXW55Edg7mvKC7IwfWSdped2JyYDwQH4zfnKhvJW0+ri99QNlFAw7b1gZFQjhkwmF3zv
YZaiIpIX4iacC0mAwkdyFNmUa/XEZSzDH3HyykTFuaKEYFitOiS7vpM/I3bNY2r3/N2/NuncpeoO
kmVqmvPkhCF/kp6IXTodfPGT+tcaoVYGBCZAl6PWSnFdHuPR/TjFXvhllG3QRdMvTqfHexuwbNNj
0g/VbSRyI+QY2oa1cT8iO2HWRsW+t/cbmuM0rvOqLWbVOGDgXj5oqsyv9nT/WbhjXsd+v3OZDH/N
08lvzWuAtZXLklxS25kNzOJJanNaYkLrSbEnqBnyFakbn4y0uFSvKLJt4CzCokkeSIr4ccCackJo
fbEdKrn/6NwXsbXKDCRkQn/emCzTVlZkpVr9VQOGYbaQT7yKqulEUIWmU+N0eDu6Mj/oft3U4zd8
0OcBL+NbF9kase8cquiphBOa2SdYHAG77K1MG53B0wIKYRImhzf3LYgpSO4L79EdkqlQ2EBCN/z4
bymsgBArrhTuTXtjctU+HW19KoCy08IajdL6C94oIT7wBnL3DQ2bIvnLt1ONcGe9vdK4RYxqFHg8
BoVC5pwAJXGjU5oS9zCjVwSZ7lbot2gIzW3hVQE9FqU54j+EuHhdXFnr1gINjYkEPnt9j9dlzW8g
lk1X1yYs3EiFnHKyDBiJ8oVGW03IU8J5v+RAqwYmyYCQ9nv7+i3c1WsO9EfRWfFpqBjfBMk/fxhS
UWKDDSISh1SrgoM+0jb9Y3ZBj8SMvMMV0v4s2KWzHnGLZkDQsyrCWfTnADYsd+b52ShVRA5KhwJq
OzTjoYX3twMDW/ulP+Xq+kLCq2J9RCcYC7oqa8Vw8UuUGOiZFs3+blxI9hOiipVPLI7kZFKBI3wk
Ag+hsB/C17fvsg+YicmSIPXkWlgb0ZIAn6WGURAiPYFCLIZ7tVQvxXyamm0NYyGYsPMDB0/A1qL8
dvvJ4uqm0vA0DKUjKynS/PnEyNLc7mFESmSCW1NC7FKjZJh0pMhFBFcKt09n5Zaendp1Hj57ZmZS
BJqt29bOiSgzfrQJ7RvegaCSyHQ7VvXSP1RamIoZbqbv1TDPpOmrbviT2CBr/2wx+1iwWHf5vAd6
RiebKq3ovW65WvYMCUM7Qw89qbCzzSsvawr1yvDrudIMI3oqDqRwxclBMg/jXkBytL75HITKcOHs
CveA2wtxHkg5BdX/yWw/7S4l7fyB9kcWTa4domTUL1Ogg4MPv085K/JSOo0j7HueEBdHq0uUxoTX
sEBmohvMyIvAhPg9LEdPnC73sJI/VHMKAtoPGtBzIw8NIYAnG5hEjsINlL3EOxGXommF/O+c+x/R
l3wPhVFzHEvmiPAW9HE8hgRf44zSPUCdB41j8yQlxbK8PtK4SFv7br+ECJ8EpMWQSmcHgA0u9UTG
nWBEmN/+7gFdmyn24yviQuB6X435TbLnGurK9msUB/kyVL0FwumA91LuYsThUfbKnuKOZ0QgVJT2
Y4jbJu2sB477k5UI539MWL2eGBiMq9CsWvjR96yHpHfXxTYBNwzSvPlwJCUldxbI1vC0nsEQhrHg
syFZ7kDBJaearZBKpcQtuqlFXfxaQxMs8rduJaQs+r4OmhwzVlJu71cSrIp6MBpfkyRx7gJvtKoI
PQlYSoKMMj/2yW8EfPADWuT5EUNmPcJXN3du+yRow3dc+rxavGx9ofNY8dJkY9YGQAyHrD1VR/UX
KqHEm0o42meNmOSexOMfa2RS0qf0k7M/eN79w1brvd6YeSt7lLldQjcnHS8L55nsFHgvCl3vCEYz
sx/dZNO5BpOLb0/d3EZYGUWvBepVfbQCtjxysMQqcL5XXNjTs4OQx3+R4nnLwwPKWl/KC0JoVfiB
EX7vhQlWZGjPEuGYqmdXl8/j6kdy4I8b23mPwTr+0N2DT1JaV43yUWl2FvKDXV5l7SGMsBl1L1m6
WM1NwA3b3QoPiPuv/n35U4dtefUpjkp/5/cq/43XWbtQrPrNglZ2Pkbq1f+M/pBzn0aQiz5Wq8My
yB9G3vbtzJpvdqyRE5h7WaR9P5mnZuVeCzTpBke05cQqDQzTiQ6nj+5f7D49YnXbZm4n3RuREJ9R
rJGD47nNjApfGSKEHb1vi+/xTnA9cZPeDDhmqt+2SI9V9NVf2F+4zNrplQKay1K3pxpUaNLFiCFd
uSMLtyyPCb4vfgQ7H2E60DErTQWd3PLBlJY2PqzJa00SfT5MDEmoqLyge+hHxPrCtuO0qF38U12o
s+53/2e/f4EIhZ0kH1Fe5YvKJhzWtCy5IiFt99eYF5eejck+rTQtezpH4Ch7QbCTV9hnFA6tmkih
fAMvzp1voZZSNmYarkGFcy483sSto/Qu3IZ3fL9woR/83HHnnStLnBOopkMQi+eYEQrt066Kxe/E
Sgbk
`protect end_protected
