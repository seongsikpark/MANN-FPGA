`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
GRGBXwNpbkVxucRop7RV+SfHJkZCLfGw5NGt2WyDH1yrb8QNF6eSseMVXISjSCT397g8p+aLo3a9
3uTVbgjJSw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
jqXv65o/36Pie2pNq6w5S7D6a19gd8HKHeGL8B5Qc0AQilcxglr5/EhnHD57+hnX5FbNlQ8vGIt+
8bSKF/pWZj5Wt3zOmuPOQr5kxD/G+5jn7uryfr2SxE0GQc7mmbXjef7nWbcqMaUOuxIUWomz0t4H
jPg6HeICr2nLpsVXWY0=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
TfzJuan1yup9w7ghT6aLYcYQ6R3G7Uo5FJK9KHvMtBzE0bp412kN5unx6DbvfC3CBjrXy056qcr/
EHHUA/t4eenKDqSUpSn8f9CUZui3VDKReYoeVFWBgeweiwAararyvde9r8lq/EnSsXOXLodbLooJ
LNN/LaMjRu4eQW5hY9Clt5e0ZyxeoPHSWzDA8372ue0pSAnFOFss6WxgtAlK/Fr6u5oornUgRgn0
sFyhOLEKcGLqeTQbURRW4L0PKUNc1b3fjnOp4qZujQvpG5hRg+MmXls/8hJciyB99PRj6HDv2N/u
4geINFxUjci53hwGbZ/Wp+BNS/uZvhCtS9ZLyA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
c0hqogUpizbmrFNBiDuPRNhh4kIQARRfkJIyfR4udJhoaZFNH7ShRDpRSxccbrXy8LdZM+Biy9FC
FABpjTjAj+2apgNUpG/nPEQnKY0ftTYPCcdw31MdFZCZOBczse7Lt1WzV2SnVxh3+YQGB1s6uBQz
X4FeYliWH3dU3SfBPyw=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Y7nqguzdIGwc54lamT75XB0+JyuXLcIBIMtRhJRbXYBBD27qHStDUhpcBK+y9w7b2z4KtmepVvj7
dtd5uKTs0hJW3UXc+MRi86YTPYKP+Gixm4wz/Ef9WASeHN6yc1o3xZPXffXhnw0y5hpbv0QSJYKU
zhCZ1zZQ/vb6CrbXxvCFjf19uVmb1YF87ds304Mht6MZc2xEoXmxO2kHd1ZvxvgAq55pzIStSfQ0
C9jYN73Jq12FOe+skni1qbCkn6WKTt/0MshPX9rwnJD+NXwimHK06vWW4yaQDaUrXQBK5i1IPHkE
8h+RXPojH/iyDCwOjeboWkVnZbtB04ss+WGI7w==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ut6JnAr7Shq5pEci/hEuxWNFXPEzUAt2Bf3gOrXX5EiBeKCVAJd5Ao7hL2agWf8owf3a96xg9yJ6
ZAtgziTZfVvIflVoAwGBpvPdAU6yANoKPixWKitLd3MwC+jE+wshmiX0of5GC9QeBqeztVqEEqmj
D0hnAaPd1DtR1PsdPQxwPnkbA1p7bgGh1kZ+LI62pV9kdfrvKp/Nz4KDaz9oO1E73S7aI34jn/JM
jctgzx3BtLtwcfqTENpYznfDl3GEDkecY0m/D4qWwFIT+rZW50nDFFafvxM0hOdg/xyBETaYWqhY
LIFMqgk3MfDbGWnPiBSmDgoAVxuiyxFkaNJtDw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 103440)
`protect data_block
TXYt/J73KGeWvQ0egKiyaYnnc0FM5xpSVUFIlzIljyEsys/uthg4c3QCE/4Zc3F9grrswNRljEiz
K4S2ne+zZCV8/6UQxOZXwtWNxdOWvBJdQjzGcSwClDB3vjvKfeOOKtmDw2WzcQZ+j47mSe0rsv1M
wvYiEStxRgsCODmNegNypNS3V7ebGaiDTk+Dti6VTKlRb7F9JRoBt2TSwFQnnZ39EsDtUNEk6oAb
8I9oqPj3vL2X3xX8CfEBhs8NDG8t5Z/H4C3qi0wgs9j72kZnNuQJutQRgyZdyxgsu+2NjXS3jFGt
YFOaj16lQDSamL8w6nuTtz0pnJLu+IRsCOOyDZd7L60Vo9fXp5x7whtRLqr2ANGEkSfgZsw/n4uO
tbVFtHAR2G7X/QQzGbFt890eWTsljE/clJ2HGBH5vO9c97mESUNHRC5gFVizPUk7XMwSLBlgUIJC
kesVNYOZZ25eOHXrU9NW2BwRu0Wxetil1IuQPXgIFPzVT1tv055s4DVrxs6oRZeW9q1zW1nHsVEZ
M1nywuQCtivnpxPCkcsxX5CpPbO1utEKKGiZDTnFloqgcF494bGgFvPU03JXczxaHi+ZDpWYBlIr
EFHCuAMZYpoMwOfQRUjNzbJMp8ZN2kjAGC2RSuDmvxQIXYtDqFrErMfyPtw+68XvxOMDRvNlkTAT
rY18OKONzZ2Rn/ddMWqIZUPwEnlsOev3gi7jKq+aP9EKRwzVOwGkqPS8ZQ97dihbugZFU/ZVDMNR
92tHJrZ4oMFqvO726SFsRfvUxajF1pGVjEqHfXkJVuY7wW+j72vhxai1zvFK7XdDkAtBa6vleN54
w8vwm2zf2FxPntXI9uuAJ/TporQxPDiE/7aG0zADd8PQGwHzsqVacb40Hmeg+mLky9V36VGHa9iR
Kk+WIU0U3xOydjucEhu+8Ja/VmhH9gdnC9RkyaOT8JOWoZTsaU2NwEiE9mKYQFzJhTU78DbEw9tK
HEEBgSgSNDOzt+Pix1tjWrznsgFZ6Fs7guCpApdVLxZl3A3zAZkT6GN+yrmPNUioZwcg3Ml/4Ru7
IyjkRWYH6LsET86U7arZNW0QCY9VLf1is4gUeW7PMk3cwhOcekeGo6uruYQIwtxhY33Bm/6dhGeN
aV1pmnff6VzZ7nQLFK/DCbBIFlDlAF5PuZkV1e93uH5TVe686TpZhqxHQL5jkv4ycLqZrJ9AQ+B4
5RskG80e8JKOtjJk/jojOQ8lgqEbi6eYEIIMGgUNvSQmTrOwupwlRt2HgktZe/MNkzR7vheu7061
uf+12NbCji/CEWGVTvbSNYb4KiogYOfZyAHrc9EA9Cn/8JhwAdJm+ctwYnYrvReJq5+aWeA1Y9zO
iKewKggxrCbqexqiHuP2hdTrdEsA+HhxsLYVwhA3Nzh89qSxlJ111wtxfy3X17Jmsn8jSv+IPMJu
OelEMbbY/VWLOwfR+r0VFeKG/DUy0lkselSh+wRch/tpcKhbiHBXQXgqo6zWIzxH/KLWeubEgbzS
poK9Xvb0o3KnnS4uAxix8JNaUb+lzIBuIR/nNS6aLcNZyJRM3VhRHZRz4GyGNp5EWfWwgQTT8mZ7
bio4mJUnOtUyd3AKoxLEoB6ErkMiwa/3gcP2+RzTM+2kI9MHFnJ+Pk3LgbkLFFzQypEXULK4oBIr
IOvq8zRmRsxpPxWfr7PlrKWb95RxnxqH7oU2Op8BfbMBey6lZqICJ3vL0gqzdwPybzYqLKRp9TWG
7dDi9++GarrxKhPWQYrjKWxe4rrSAgDNLfJz0gaQqj0FvmOL7P142XLPZMwgfO/Xs2tzp2j3KmA/
woWiVVDMDsBpRF+q6FForKefMqkmkARPyI5fwaphkpi9bRCj4mL8ohu/LPhu4/nznB40/eA45i8F
/VyyXbFHi3/mTzbGPgHtmccZdTH8jlawEfIuqAqHX3D4BTgpIZwcRMQH6rEr0edeWDqpX/D75Una
8aCpIS5sdgZDWWyAh2E3PkEgNPM4pibPbmykVqNI9RVMic1Guq6dpNkC34z7WxaHNhNZjonTj2u1
b81/G5xia/o+po6mwNjo4HZZZXi3zDsBI0WRaQchiRQn2LUgycqDLr61gNSW4txrdoaowcvVz2Ze
syCzTUQRNGaGcTI/4M5K/LkxQ5iqVcL4EyJadqfa3D2hxnHs3nznFqQCq7/Y6n5eJbykoGViu+3T
31sOdHvKu6xAkFON5hk+RREq9FIN7H5v55Hh3Zfa6FveOLfMw6hZUD61Wh5eofV3S07Q3n20Ia2S
+/rSvSxWmtb5eqkYk9h4E0tGpJsXHz0qg2p7ojBVpwkBOyCWWkuyQDXSCylMUGaChrq145buU0mg
vsBJ3zQLmso2sJb32umNKpYhg4nfuD2d5iptI2g59DpvdvqJZJnPIUlMuT4XTGT2mdadL3RyR8Lr
3vo5JfMRlB55BVOzaNCg3yLDATK3Ylel2nnYEHQpDXu2LqtfdfPA/mavbffcOscY2knJTT4IcoC9
xPilD1Dvs9PKSeyhbBVvDub4gKY/GHJmQnQqZoKWNa8C7HB+cuC5WhCcuq5n6oR3ZAx51qizFzOX
+wpbqcrH+eZTJOzGE4mKoiKzVFYfe0f9+ktRBfu6B3MUWjadbmGCkts+2zZvwRftoBHul8wz9fB1
8g3XWgjB5oDoIRn37ZXhj9eO+omTJIkVcfsI6Xpe/4l2yXZkrE1OQw9NkR/Ti864OZNe1j7N3C/G
cW3vcDgZPTCcaCI9HbQO/5Q88CM5OQ1t7WRUievToTcGQLATpK8+uHV10beLHiEJrWk1E9JrPsaD
RP+o67xnA+qOSCm7KWvj5frjHSmfI1w/zjOJp1XE4XyDh7TA1R/uhYxF29RmLnaogqLf9kmVDW7F
+X8i3cR32HrBiBjvGmr2m96uo4FW71otUjyqz1XwhLF4wyO5p58ktzFHpIp8086dDHeijZreA4kY
Si6qoEOO3O55oq73KplT1CgHAeY3O/3f++TPRRGV2m750FMtImkJTlstFPudsQzRYBG4tSwZT5FH
PpA2N2x1bm+eyDM0Pq7yKQjmISKF2SUehL94PnE7og5D9AodTuKXs8pYdpXLkYJoRPAOPawkkKch
BCk6z0f86wLq2lCx05aS0Glzj20yASpZSRumq9uRfe+RHn0ENS8eHZH/caS0QSKpxfVyhKMiclgY
ycAuFFLQQnsj82VhkwoaRQlfxDk/Bxj3afvngIVcLDk43ZViibpAj1Cq4HYMBGMU8zg8D13qz5Yh
JY8VgiRId9EQ1LRibgy5VCgyNVW5v/PluMIQW4AUnJisY2c4OdtEu5A42e5YvMYs6m+1lMPPVgr7
zsGdy7uDLUJROOdLa4AxlzdEYhd9fg+/O3Ltd3up9URWv4Q3EGh5duuA45eeroc7+qHAUYcN1zWt
HaDI/miju1ebYxAv9nHHRttTUUOXPOwkAFGyMHM1ieacfP8gF75DCCVKt2xnsslhxQKnWmV5Gpvn
gk1h+gefn4UgJszwZlgzyCqz7X18NIluDOEg3gvf/TSHfurT6pyOTSh+FNY3w2tntCQ1HVIoYBBq
7R9wcavjoWncjJCi5FFJrSzXrmuGgYEyaUfPCsdUfjFQxOIT/YrSgoZRARAO4pNXXNkDNZRW0V57
aSjWx6q94TsWFprcAqRCYC/8AV3xPRKmX6CgKku4BYK7mQJkV9TSF4SYXJ98BFF2pNT4us2Uz22t
0m4Jz2teclQchI/wPIoHLWjFGq2saDqWnUZMtTefA69bOSZdkeC2AZIuaDVG7LXfpRdbRqpfL4u2
qLOmQTWzhEI3yAwBbIBqxcwmQIGvUEbDFx+mHVi0epO3xSXUNg6w0tCZbEK5N+H27incgmjHiCgD
ukpK81MICuf10jARdv/Ryi84uxtbYQNqvIWwv+aCG7u65g93Mj/J37qHxkcvAsF+FxpSM448RyDk
7m7RLsnyeLcHUEM/Ago9N0rCUFYpyuiwLyXpC4Il33p2QG/DWIactHbkBY4KwW4+wFvzgo/c2FKz
Y2jiA8kGRifNNGTE84oaX/5TEV1CM+R6RSGcckOH8dZEPsasEZLJq7T3O48Uz9yVqK1N1x6lCIpx
wEEo6sxJ7R2sC0HurAxKfTLyO5BJYVBvsLUV0enHFwv6g+JkYcp1fcUBl7hAZujvPdXscNZU2X94
PrpvXr+SiPKJeWAmc1rLoQnr2ZG/8SDlJ/PGpieuNf+zTBVZkbVwx5wMPTkTUw8OAGs06B5zfrja
r/frjUmbZqCXtvytOmMtmAz8twexw553Eq8/UZ+lxTZjpQmg6RvrHrWDvL3wfi5cxNu0OdR2BdIj
pfhw/kcphquhVl9v8Ie11nj4QR21ZM2N37AxZPnS3zQW1vNB417UqYEVvEsF/ZzOTcZV3vyiAb+N
T5v9iTfLArvSPmxxSP71IyvZgWekV1Z08SiAK1xRTGTkSDibqSUZKm1HSTTVxdHGH3oDrGRr+1mL
gOB1UzlPyIIfUKdaENOqMFOTlOZ7nuDBDanKZEn7Q+iuTWSDTLx3Eq1K8cGHKrIGaKAU8LCDe1l+
jJver4Oh8E5o0zrm+uly658PEncP4cmWQqZovuEHG4YNRe0swji6XAwEXpQlWKRPHLJo9rwVEm0/
N+2hueGXne59bQVozFqlS118LVYTcUrneYFcbxv5+6M7wL2NCmlhhpZbA1mob6xQYfVT7Ftc2EGt
ApIngDLxcyKq2THT+8L/x9ZemC43hNbPg5BKOIsik9EaxgUzd2LLJIP4AnEPjI5Y/xcnN8xzIv+0
LCXp/6A75TlWyxgYsOd4WJGbNCKlQkO8Ey2gQLJcM5bUMweAY1Q2OT5EY+FYYEGjv7kpOC91wasT
HHYtC99vW8z5jX6fVKkR5XNWB14ionznoXN+cESw7n6HQ9pS1M8OEavIAY+qI7xZKhOv1OK04xBA
xN9qqnZQI+bg2V0SxnnTELYkyZnFTJvxX4bWn8xmDWj/cilPMhFMAgUEf2R2JvW/4TTQiEiPdeNk
/XUdzpYDm2MfT3DB8DGhpyGnFdTJCEVBtqQa0KPPdyaU7jZPKR8QmFRjurnCV7K+JMGWdWmKkFFs
cWOOPAY5tZLm+ogumjBZ66VZHcy3loshPWL0QErTAn7CPIkWslKLMtdIUaM9p6rHpwZsPj1I5YZe
hCRiS1XNnBlNJ8MPtRSLO90mIbvRvWKuurRQnuVlQD4oOcrrifbL5K+PoJMcuoh/kYRm2PAEfDyA
QJJi8fKaHxfAxvepRfBqqJUtVi2A8xCy0jFwgxxTJAoZqfbhJyG+T8Ps4znc8fGp88mxJbDiRCVU
8RISCTt4MV5H58nLZrEGPLcqXrFgXLNvJ8K+ekrzc/MlFrfVBnmE2d90eS26s8erbWprfxgLHhFj
uQaKuuaR3y2ZxgIqFZCkdufHg9z+Jkj6z754pUqB/tyWS1XSG1lnkxkRti6/Q6dffWYrR0c9g67F
foL0vuq8DeD4wKLG+Ys+966wwvcDm+3DOe9l/B0hunVl3+gH1hlSYIR80N9bVfoT+Yd4c8KVvKt1
xN0wOYfq7tI9wSDabwsbjTFLdlzGZEt6KmVLSOuiGp1PTIlIa32/iYD+p87f6Kg6tidbxQfgcTka
8cUquyv+BOgntzyq1y/24XD6OxXr8HrmfgA15Aa4WGZeI8nUEod4TzM09agCAuJQZBEcuFCuMaQY
+mMzMOE/tiI7ahsGiQlxZ0tLJXnMGgxvxSnq6R7nJPcoTyGaf2J/Z8x9XDXxYbnK+0THixvLS16N
Z7TE/65wyewBrSX+VZ96TJ2ZCUFg4xkoYAl6u6gMPddlo7VcroBNUUSzo17ZV0uDXIWfvUkp5595
bOVqQB2/sdyWz6pEGkRv4tf0a7TIIiRlvvx0F7iRELZaFDycNJzGB9SEIcHks9WBKPtmP8XW9bZH
HiAkY+L3lp2FH8DR9jZSdZkBSvCMXcJey85sA0v0YjCWxxm1fsnt+KB3cTVkD9DFiSJS55WG2RAA
PgAOld3fk4xeN0TnrSKlNaM+RkHPNMT9Tfd+TTPfHMAPDgetqsrPejOthzhJBlEED6A+VXlEntYK
ff0YQIA8Cj1nP8nRR/UBpHg2corL117tVnWeI2FLWsOZjvkcKiX793PfK96zLJgKVC+CQV5TBWdH
EPHbOzYHPSXgZUDNMoLT4mbMTVVX5oZlu/YvOaRlGss8qkCa/WezzlG2sFEEUL+OniptOMxat823
fXPjhkJym0mZzDPMcjjjh/UtiYh7UHihplhNrA7j0ufGHghoclcTOnTXGKvwGDvfjhlt247Esuf7
6dHV9kBhbkQTEtkg2lOtdMJlgj27VFOMW0x8ninPUr95qA5s0nN27+XESR+d3eRSDy6s8geRBLPM
np1uXaUK3DUpLEM5wZAh3n+WwLaxxHODjpbKRsUzpBGn0C7s4p4/kiYSEdjffoC/TensbxD24/i5
S3RYq2/FaoVJQrYEtIpaMVZtk5TsjOu7Yi8UzEBEVmsUWm2bz+CT/l9nIH/fOceQ19XFs6/kO4Gv
KtaGI33i28cJK9uBzXxmctdDDbZeUWAcLMpkZOK6FvCi6WEhMe8aCzCziAhmLUIsIvkWG+ohujGy
JC384LwFys7T/tOqNMpt0IDNjawSC1mrvsTu5HINPrtkaljZScaDYAX30pcPJrVO7vCzh420D4eV
RcrRxrupHXOv0A7z8RZF8MpgRh/+5ZGF5UKchbR+Bw3LC4LqV2V+GDgkEor41u/hw2Rj1hS/5s5x
bKeQgqcdH/UObTmgMb+fAtuAepCNyo33uqdtsjMWZOuxNiFycTZ/wmmzsvy0KP6LDD3JfmN7ZFSr
GKYWCKxyR8cAoBXEox2KmaO5CQlGzFcer3DCdiZOPOOeQbzXKi1DN9REG3dbf6v7PPUK71dThxxo
uVDTHfp8LMfOGzEGzxhdZc1kLUGwTVDO8Ng15xzWTdZlAKqLh7lGtXxioYX6QN6Nl8Oox5H8xVg3
SGX9fX1qKvVU8bN78RFQZCzu4TLw/uTWiwR4bSS//OEXuU0AgC0f7DYU5CjGp6sfGbJS8mP41cpF
WX89WygHyKoHdWRw7KRJi5Br/Qrnfo0r5maqirkojdiMlnlAixHfYh5kAkk65rVR0qzgbgxRMU4v
A1O9LsERytGs0XSYPucB1JKPkPxBriXkLbXW7NCTF5nU6mWWaKYHbfeN7hU+N9DP2fOQ002r/CIP
3XNxRnaq+tmUR7Gw7BMw1m+ALzy5LXGVGe7axLVvrSFGzTufNDjvwpXAm/N5sydB+7b/WjqDGFvP
tYEvb2CgHFbIgqe9IZBn/kok8HXnqAqCvIHyb89ZZSOZxItycWGZGZDPZE7TFg8NHJGjdtlIz9tL
cymAsVQGYoH5o9I2uyHrnaNMDBLhoCJtS3f7PGuveA0XUIMxh1A48IethWq1JY2jGLRB0os8Hg+D
u/bDi+tsB4kzoRO8CqwiM00XcFvaTl0qhxktlTHlpg91VniyGu0IfCegY4ZKCUfje21ONl2abTwQ
AShVLsNdA9S/sY9EZ9kpqo8H9PycGfEdAEKrpH5Q/2uPU3wS8Ix3LdcaIZ22jYabnvls+eLncEBa
LZ6kD0rulz1KrpFZsnaVtBgt6CS3qgyiuARSXlAhhCsyUgEIljfeBYKSgVf/Gjgp4QCxxNGkwyLc
xoRPU0Ang+e16f+BwerY1rHOpEra8ZmYEHyUiGILuThY1dy6cRR/pcMg1xtuerAMZNpXCfMERegg
nGrFQQdiUF5KAGWKflKSLF7W9fo37+8PjVZRt5GTRAgGRQPJchonG5pXui0bPQ0oa4UKBe9K8wAX
QPYOPKAn/b7zFxfgo2pdvBxKx+qK2vQibDL9rvTxxQTo7y2ZbSLrRmEd5o3MHNS4Tyq307UMXGCC
jn9CgrzwRuyVyLhedj6ZuxKZC7hifU7zusy51CkVqmUj5rIjYA8bFjHxkgwiyzmqgxWu0hoqZkjz
K/hN1xirAnXSCNK8Xhg6P37h8mYbIos9ljsn/NAQ9ZjBJFF7oX5qQ1I2s3qLSIrlVyv972LyO4tf
tBR6X3qBVtpITRYw5iuoqV8Qc9I1aG77MW0BUx/U2RU8lBg4yADZryyKNpN0o3dBU4E/W6GCiVf/
lHIhsrhW6sjIsi2D+E6FlVyFfdUWMOGCrsD6ixlaZKe+f1Ho0jUmuSM3Q/f2boQMlZ3zlS9i+QPp
U3kd0ta84uoTzRCrrek1mqEfs7CQGBQFWFFPvYwajyClge9hDDh4tYfiQMd7e8/RnhxaCRZty0tq
TN8JDJohfLt3A5z4eDH9NuhhQEM3du10mD84dix4QeNHjfeJKcZsLsqnhbnVfrA1GWSE8JNPsZqI
FxHsb3P609/PuubfqTOYqs+4oQdW5bIMbT728qrZHkRbVKTUmQ8G7fR3vcxCUQdpLrC3Fv0uMAsP
ketckcL7rCi5Xsgm3AxaKRFiOzEtPCqQQ9042/uq1kUn1pLaq8tM3KTRTADGcQtpkDm1hsXcVZYH
eC0SDgXSA3HPJQYkyWYpwnaxbWfgnJPhSkxt3PlwVmhVoL3yLH2pwzj5P+ArFMqkaj8aleZf3p8A
vmAsg5KmuiDRZRI4rnMxnae3Mb4Mivzu6XUq4btTflC8btfEuDJvAxC8KBSnWwOHlH+Lewg1mEpx
IECHxuTpT18QOYY3qbVFHc/JYaK5WdcxoGbTzXzvqh5jXyvfg4quo4P7nnWysI5x79pCyNtdJgHz
El3NUzqOTUMLLfz2JhArqEOjM2w0SnJ/AfSKIEx82PCkS7hJztkQ9WRhl/Fl7YYpVYiPbMutLXeD
iuzggL6iYZ0SsGzhZbHqYQ3S2Kfa4aDQYeYWCJSqqirIS8fnDrSefclnO56tZ8llwWa1R5jKXn75
Gf1Kt/jFy2ZyVrXIcvnM48WxoPE1n23jeX0AqiUxC1i955skt+tLb6fnxwvefReLkCJN2CUU/BGh
xC97+rEOE/+tqcMsvjnhpRrziBpVyAwvW+DTX4GaiJw/+t2q0txuODOGdUeoK95/Jo/CtSKI1O+o
Noz0/4w7cOz1J+y4cj7jCSmnPLqQbtLjjUAaqXWT5HsIe9awf3GUFLdTNSjwn7W+pgLaN+RVmdrY
UY+X8FH21nOYuN9n4rdp9TPKsLWRCFRorLux2gdBVee51NXdIgTJHqvzC8r3nyWCPoBy+9JvL2NK
TQgksTKWPd23y8pWGO90QRE5AFYJZoNXU2p4CJsj85uHkh298cU7RXhhZxYAvZ/D+QEDaIVdTUP1
d12Fw4/lvjXBl1ytEfF57HS7DZtSoBsfpcKc6rDN/P+a+hMdLcjSRj3UqDRU4g3jvOlCZBiKh3K3
ntGh8/Hl8SMOdGrplwJ7WCKLmPzJq4mX4ZCo8efdhoHQqNi52Wm7bR49b0SEC5pme5BKQpJeK21Q
RpfwwCvLqHCkRje+UGD6DnNF3jF/hCLRL5bvunYbisysDSkEBaAWRFr/oK8Hfb+N0Vohi2Krvxdw
agmxPdmkq1AOtxJrHa2AqMZpjRIR6J6weJgMhIpDWNI2VjKJa+xvb6VJ4lJ0wp3BwFGko8W31jmj
WJbtGL8+IGpMZseDDXi3M0YbsfQvaPhp7H7xkd5w7Lx1DhTPF77ELV7dYfbdcJDsSC9sigkUMK/2
8o266C3yvvbWLznOE3VfTL6eJM9ubl2CewU5edv+gMDJesQ7JUiSA7Yv8OyWL9dvSzGtUY6rE7xm
NPTyoVKd9rpwVb1xGuGHUFJWpn2UgCyNTMgZ1g/h/O41ECgkZl+8yplOXa7P+ELCi3hJSXDBpXn+
JR+1t3ib1Q4/JiKIDb8ZQa6NAwhnBBk1aY6qqn2JbNi0CoSiIxpKu2x7STSPKrdt9xNd4AQ6yNg4
vJGzITg1zpR0sHPTMqSQfUI3Tow6Ic6dEyG1xJvUFzbVCyFuBCnt5O1vn3XqdSirJXY45JyR+k2r
eH2LCkTkG2QAf/z03iM1GYN3uc9cwk0yZlMmShEMEElkH9g+4lhuM3udOhnzd2fEDHKoeVShidiN
yHKPinBulNGNDpaU0VOSh3sztd2icJOFngde1aeHDaaED01yW5VWDsMPUOLHulCGlrIeLI3VRcqW
8SkFRypa/PdFkM/rXkRORx6lwyWAu//ODLps1HuegvzFjsjNnTuIkFZpnbLHC0rTctRgx2Lo24Di
4n/kYvDJrMSjDli3Tv8H75+9sQWIa109+2oGhuXKyFAE19ACMvVjCjBPOmZsXKZpUi7IFMxXPc0W
LJNlswf6as/WcxmfGOoogZQLNT0E3VCH0Cak7jeEXXGxXiLGFEw2jsCuk5KRG+ilx9ZMoZWPmSry
2YMZoe8iY7OYvRmcAi2emnOEMI3UtDXc11KYpczMT+M3e9+HtZ35rwfObIJKlQ4GpFi3rzKJwLtX
k2A6H8RB5JUkw2loqZYR73ogc9mnjfNXYZMJ8/NdszZVlN50PpM5iC5JNQqLNfWp3lvSB1gyIvFm
HEtNGdi8wwJ6btDfMn488QKYdNJRCR9HJsPxsNWz+S9/t38tlm6PDJP3yUM/OPUS+iKng5Ts5THx
yFgbzyQygTxaNVanZFDv/oP28ocRhN24xJTxeOLxKftp2IgBvTLhpkRy8qVHHT05zjL4h165dlO1
rjndHq6ATfTbM7COsBqr19CM0waEdNbBUXnMW9bcJBCTufd6r59Gj2mKuXFxiOtgNMPeu827J4df
BVJLOGatYZa4IgV3mmwfDPSZgZFXlvADYLesYGI9V9gym79XNjVTuyfNE7+yhCHpYoUVtve0GNCD
WeKMwALRciJgT4S88o8LrevHKFj5LF0+eanicPzvskjVcKGymPtVw4qxju+5RzXLg2X/t6ZU7iil
M9tir8TRBx2tN7XNP5T0Nyb7sDjbMgOu/VwBaATsGRTpy8qOBc8pNlClIu1E2ZNQFCdRQE+FP0xd
VK5ZC5XLxoxR0bhczWKydMbZbUZ5HbcJrRtoLMiQ4uzdaTKpOjUSQaeeIdEP9DwAv3/GqX2ewHP2
BPJ3+GE38h19uIbluQdiDliOrw3JtSnqg3/NbtX/BZ8cQe6kWZxOOdJAqLbawA5KpA3o+DpDwYMJ
Ltp8/LLl+hd69Y5pQxD7ho92soiSNyxiNXYCN2132wBbn5eB9k2PFoW0i1rc2X3+GPBPkjAEBrSX
xGanqxsKD2+4gy8AzUHLNb25EG/uAnufTWRfzjjPpyeXs5T6bLQePXKL3JuhrQV+GmxcUdWFezpl
48upHT3q1NNlcVhmwbHvEpyeW1WLd/TA9KQnmMnfcFYdbf0B8Cc+rH73J5vqpSrZ/RVuUwKskqdR
fGjvrVMXxZ1itkdHxt3geQ+d928lh9hk7sNiaYVE5kLBQcUszSFRauTm7HbwhQG9G9yhzHQd3c/3
EzUe/IRW6Rzt0dAJaYNFKAEWYMsgJZwmL207Jgv31gTVicN+7cLQrv76gWCUhzOKBETz4SBYrLtW
wQcm4Gh9wFQfuKBw00pXRy7c3Qg4iAjnIcZiY07TaCo1JaDBB5yKRl3kma7j+yQi7PxU/y1P2fL0
C+l+JdK+Bz5JIAZeU/1OobFsrCznKk6l0HCHTZfUQuNL1D7n8cRRaPyFTXcaG3OkY1bYuuljNBpX
OFWIFZK3WEeu5xFMsM2sNelJtFWvqnsKJW5iUFyksVxRXkw/3kx7lyhvqc9TKSow53F4HNOOJfYb
9r4l5bzPQg+MbnRjWZ7TKWLRZaAynx5J4QxWvSGlKfIMENnHl+S0YPlOV96bRnPzJjneH/zMLaHg
kqHFks7AU5Gn9hvLHti3UBWM2uOdsc/UkUGFVsSjxcwh1GUKmOUYhRPr9Y4agLzZ3EyPvFhSJ5NB
lt1o/QqEpaWZy7bvnmzwZ5nsykSBxjZTi951GKmHtE4XMHtKAJIbYCQHtt982saMPzzkZCi5LFiA
vVewcWlobWM89wb3pxTIcTCgp1Kg3dc1oy/F8qXcvkxwqpf6RV/Ru/JmURCW+qc56pjCBi+S3oRY
MJDFNCjwum0SWbSpJUuDjvNHxb31V7igEi0UyHk/LDWqhO/xPfJ6F/Y5Z6oYqnvrc1IvXHtdLk8Z
P36NS6ofiiYUfDd5Vxnj7lXDyPaKF5lFA/5ew6NF2SCcPTZDCbk/wOzEqxPUJMiDCKGk3/hlrZ2s
mlKDPm2IKUlVqDj0ACMmLIg1DnedsnSc92S/wJz6KziwndF1BA86Hj2fJIdYHDPXtA3PFaGiWNFo
NhBcP1vIGcFuQYmSsaPau+ND6iZLii539NpRAR73Nk4f7qhOwUkVG7NKi9QddVaG3CpeKd8+g7TP
Gspu9+9o72A9zsmdB0hCUY5Q5CP6pN8zVXPhVsnSvI6fnu1HUnkkkTvrQx7cWjftKKFv4ozU+tTX
OlRoc/Z9mTo0fX6zvXmp+PvINBcaIJnF9nvX6/BPQ6wkPelMmQ0tz60r7UZ7J4XXUSJ9TLMUh2hx
/j6gCmdx5lfHL2c2dUib5dHhtMUKftFtCbcD94mCmVztOWlLFziUyhL7VYPPjth2Z+5akOiuxGIK
S6UUBIzgsjIWJYIO3//AIUbBKS/LCPq3grJw+V5YS/GUS/r8atVwNNdVLBeenGfHz5JeLgt63FT4
O1ts/mRuC0FmTBFnLfLEkuouAEYob8vey4ATdLOLN0RuHReSM8xEGKBP1galu9LT/JlJ5wWtbeEW
HlBkZmyoBIghwKkqJqvjZh0CZoM8XeBK4u7t2Nzy4e4jNVoBHSyuR3Q1bpc4ULCu07zRQl5zhG2j
6CmG6DhieaDC2Vtrb8MEuZ4TLHSrDQnmqIgGWCTi9Xi9bW+I9HW5chrUpbU81MX08qg33TuUtnnL
taGRmGfxQH42TI2zqVza5a3SS5bImDb1/4u7930mQDOG8aKBhdcweuwrLLI7MgmGx1NkOa/l3ubC
zQka4KQOjnnnx2KMpQxxLNFioOlmVUcZr9wUnXsy1o9GidgF9gL0NMs4NVlP9ZJ2ZY1rSnFixg/F
VLWdn/wm3BdwEok15JYUSAN6hqlGM5ehHh4QIo79SuDISpH8DA9BpxWtMbGVJMzlr7AIjVMuB4Eq
ez58K26+jsCEal+aOSTRDjUmo+TJdpoVzOhRBuJ/aLraOGEVNdla20SybgKXHEpoRu/n2rR0lTRK
A0CK65DlVfnIGbpWskj2Zr5df1OLVYiw7TgbG3SaWNrBNz8dAZ+v7Q/d4+1q+78z8pQRma2nx6sL
BQgSUH8YN8GUXCYNSj4DS71O0XIp48qXc+MAt7COgQpkSb8+U8/ax2xws5X5ZRNfXFjESOP+gfIv
ex9itrGwG9YD8YnqmY56thVZtNdLXT1Upg9DAeZbZvMYtBOekIjmkQ/gI5zlxpxuh4Hx0HCkKrq1
pa/PhXHoC84I2EsNrSDt+iVrhnwam83i6WRp3sfZuDDVXK9jOVN740U+PfzWQWzdwylTd8gzwe4T
adtIgXqIMuyPvYfXisCA4jWSEfdx5uEDa0AWWnzurpcfgmDP5dAhXdMg1YPk7P3oHcCUocgOQ9pV
UHELbwmlOvTgB/DVJgP5mq2Iqxv3GJTVyJIrnUwZCrLI9n/LVVMVI8uaU4vA8M0LaY5SBUAldGcL
0avK0IuaO5aSxDtIhzWrUvvxO5IGU0DdLKp6A+fmfz6ufU6ZU6VguausJTmhrK+wKhsyihCr152p
cBGruboYJwhi9F2yWfHMr8uKZbYwvq3YBgP/fRvUCvCu4oZvqtOp5703n8V8LTD1rI9AgQrZe7iI
iGex7p/9rrWi4yqB6mwRQ1Jy/sJkSN1Z/sjYDzNqghDnkDf+hOpBePqFHOO9rAZtW4QEFKKCHP7K
AtZTe0/PLTQoRIfY4MzusZW4AwbpAmVG0nL+KV4AfXwbpGrIZQwaAE6M2KVfkyz3/QifxeNt6S4o
9QHOhPCH249FypjHnveYF6RWJgSsZOc5c5LxSR5XAwcwOh9Dgzh1Yh3LZ17CBRRHrRbrn2RrVXAE
WUFkHJtP8aJ8CkpTHbKkYk802Mz4JU5RlWvsYRjhd56Aj2xoZs78wGh9QqyFY9gwpmWgtwITmmIn
Z9jWlLLTtRdIKEyBYlo6HAxzuZDm82ySP7ComjivZTsa+2BO/m5CNJNiRy90acjXyCPPiowUVuMG
8twBZj87oeFTO5Q8rD1ckFVzyufrlPAgQH2Oc85DBhEJWhO468LWmALlTbjiv9XOsj/ll7VosCaN
TBmDxqE+q64C0+gQJfPNlmPRDT5imYB+dRasn6IU15iJ/c4DuNUDc2y1M2YPDam3kcl27pVP82Kz
XIBxfQFSFDJWtEGKAUns+cTqXAjFT+6WdcAS9HoxvcEZWeprX0pDKt1Z/WlkMGpsusL2CwSTMeW6
Lu/SHDSgYA0gnP/X9RUekw4bbIiAI23RRPYr8vwJkYHFeUaR4wKXevREk/e3aZmGTJZaihBBogJH
Llx5baItC/Cb+17MZoSkm4xFLjMvNWMHGSIOBnO9kl8+FO+9Jgpvw83eilYfbSenA1xGEQAfR151
df2ZMG41hfAKm6S3NHKTw7GLytIXqQxp8pXyazBIz8V4R8p7ep+OoqfWrscgwR2bZ9G7/hMOavuN
6KqsR2AYx64Q8KCCQm7E8WcDAealmP0XULPXPlfOvMHuaDRQn7TYJEy4wda/dUCmoEPm9/oXj2kf
NzsJT1G/cpvHiTjX6qhUh3GJBrSB421NvUs6K+I/KGIw+A1wxDyGvHDPFQv3hq44/8u3gQaGsgu4
tDi8s7r36Nct1SrVc8AZo+Dyn5LZPBpSWLMWC3PGMSn8rxRWE/X/y4yFlpLzbLvVB4mNXKIbzNdW
xOq+fArcpga/n6NkEVKbcjWRjXEWL2uR0fyExeoa8klVSLX+IWepqT2b1HAVPGMB0CIEiV5DOLZX
UwIscRrvpHY1EW1+WkzU/0jFKHrCDA99pACBkt66JJLqeXYzUpFQxwW9ZpqsROQ/V0xl8QHYP0UN
m05z2X8oCU2Uqm6gDI2BM6m/W5KXZGdw3KGk5U092jqU9dtCJUw8xUDc2qVJ1XXWKfucKrg66rR4
aIMhS6ukFm8IQ7eCYLUi68AlVnDAkdz7naz9pldIeial4bv/wPR8EO+Yt97mCn9yMIrGXTCsEboO
DNu2ssdUODyByT+i3R4y/yioB5xCqgrDDDFZpcGU7308ym22wrfA8Fmg2Bk++dz3NxL5tweYCq0y
Dy9sn++o/yu2tiJIip/O13dnihERW6rHU6KmTknmibbV/us+1+xMSxaXK73oN/PXlLo78vV/YAAq
DcqqY/omEl+OA5S2JAMSkcMMGzEQbM8TkMlTgabmG2+S0RYexsqk9IDNB79MrB5SsBbe79ni69li
qF/L4/6n/e4dl8vaiyuonv7bek2k1PtLwUfqtwkpvtdnCkIK5uaiEXq15EBGtprJeqfRVRoqZN/j
/3wI6F29p2a0k4HpmcgxV0xdEe2NIk/ZmbhKSJzNL3BbnXe1z+UHqz2szKw3xBHzAk37AQw2Hflq
7029kwahwmTSnBwEnlTr8EbVrMMhxkz4b5xHCmB2EmxdQe8k7XjhNr5ecMu1QCGsh+RBt42V+VcY
+f2FYF2+vs0XnzQVVyIFaKXN9eHODwxKiNms8CIrwrCvYeHWZyN5F9heM5V2GNAmLedcxkubo1eV
julvOTocHgTC8q1RDpj7AGgXITcHwi3epsLth6l7dAO42MnimgbBi9WHtTLKAUGdmlhGKvYsEqRT
Bfa0Rqyfr8rXhtcIg5SHR82tH5M0WFVdEdCbj5+DhOMANjEGDhlyt3MYPGY0lYOYTh9yS59kvUlC
/l5kBPNWOJLO3V5gg+4m3OeTI0qca53GSoE/tl/8DQ0KHn1SsWGw2bcKaY6r+He5IY1HAWadGeCE
UJO8wcpgxtC8QcUuGgeBO0KbOUfI8JcUMrRMyP+zOZWe2dFpq5U/J+gDILfJRI1p6RK0IUeW28E7
0tvsoxTVGxue93tTVzWcOQo1aZIhs8oRtnh+3gZIGCCWb2itj4uxSPe67gjDOwtPUOlB2JNHVrjD
Lu4yijYLKePUyIJiVmGFWf6WOCTOvMCtgNeINpZJwP6kyM7+TSCNMOtykoiT8PL3AApUaMs65uVx
4v9VW/HwWQK58P7izX5o0lSo+dQvDVwpjUsvazzqMK8ynhTTfqUH81CEzDpkH4nHBecfy2zkJbGS
/Py0rndJdyPM+9pMrMpPlGGaduRy6Gw9t0+/kjFYI9VfmejUSSC06yfs4mMXA8OaKdqBrOr5l9z8
95U3HoxM3cgol/yMZLy7FPWu1CNX1l2B6O6mxDmtQdKcFAXpLd+jdHc/ZxVGH9+oLJAxvK2NaGxX
JN8d3C+4OTt1/NSOPY60wUNJSE6iOdDJKMukQ+WoOGluvsaANpjb6UpJT9duc1UpbKzegL9y/3h9
ACuNuZKwRWkrF/V0l1CeSZa64RU2W/tyd0qLpgCJWrkfmYbM7RO4qW+EtBO22SEpW5yB176h4kSt
oG/ALWEUVm0PqyRqbmaLncMGsb+RzojR7hkcG2YqmHOqYufAWjXK5z5KxeaR3UkCXEqd7jhEMd7N
k0jPy02m8EG1EZY2Mv8UrHWxspbxHBQrGtd1VcUrezRq7lsieBTPePGvzWkxRurBDsy7QgtS1uxT
VrR6tFGSlqdPggzjaGPVQPBPdcL4xaL34KpPN0E/U6c1Dk2oo39HVSn/UhLqofr7xUpgQqvca5xx
ktqcmhK4sex6t8a//YH0jDCACNQHDGy9nSriBsWNUatYOwBQB0JuY9VppBpmx9S10QGN8s6j/zw/
Pcy2bLygjJIdG4CVfy4HEM+vwTEhZ+8chawdAGdvMQTrTiJNcBfBf2KBj/IiLjvcWDmmwKWB6VAB
vqY4trnwaTnwpHkLH99fmG01g2+9SHhqxulUNJKeE4mt9L8ldoJhApehTm8MdXXMsdsMdzuCeGZk
0ug/oQs+TQcCEF070NyOloLnZepfjd+ERL23gu4w4w6By5r8PHReeTrqopbPCvuiUAB2VtRJgiwG
rTswXTWErPqClb5v2BE1m0I+ql89mvl0W9wTTvZBT4AkWWXZumpoGZHvveWFCoap52TNMHKTc1th
dzItg8UESx4mNHX63U+3DebjlUEvaGaNtDfdTu8Cxai5wjw5i+Yj9S7E9Q0d+ATGicIgDwXcBx29
07/oSIgC2RKXgFje06AvD88mrpD+/1IJmFpRDa0DEja1/XebrWpkE5YhWS5Q11W4ompgtD5gP5eW
FSG9EuJx/IMHSjuOMrVPRzTqLsNVpGnxrzh7fsx4rq4ZrfOJNbRBpV1nNkSATszWEu1CeA209Iie
79LIYgDtdXM7xnyxxr5o4PiLYHEIGJoEKSSExQucMURPh+rtPYuy9GelzdxX8+hYvRhCFpn4wkDr
ZeuKLE8UPkzqIRudaWxPFCFr9c22RKS+PgX7FAMDyC/OAs1YnliXNrytSdo9Df8wyvAVwxQEnXzi
nMOnpSWkQeJDvvehJPLoRaf27r/iLYvmPaYHagpehbmZ05f5tN47fNpZSqr+5WoJEwuCvb+mqE5s
9q+Fy8aldsVpcMFGupw6neots3nL/OiPtVDeFMqokp91pdRfx27l4PxOLo3NbCZpz8NYgGRPlET4
k/GwUf73YimhYi4TRE43UNFqIDetLWuA+zMfGMKxRx7asCT87xseRhpm6or47YSLiT8Xwfs+T9gt
n80Ncdcd3IDPE7B4/TKovdkQh4b2SGDoKCF0PorkoFgzGgKaPONqlImjBLOMjeFK45j9UOfYq8b6
aeldXtwTNDGcmhYZcGQs7Eg2QxgXr1y61qonF3pxccUfyyzyOAMtupzDg0ND1KiDIyhwo5MH948d
R8FKr3OE113nwuASMdIu8Ch1TMYKaiToropn3WtUm7gwI3ujdIZl9zj7X0R3mPAftFCFUQfKjjh5
GNedoEefuC+mlHG8sL47peCzzlKQ92uUTS38sxPbapPersi3qQQBrzOEfX3eRfcZXawfttXbX4A9
JnP4zKR4ViH52n/tNOjnmKhAdzGT1YJ39E0cbCaShm8LdrVbrF8bp7XLH5EXxrrcomp3HAARlQGL
4EN29o0y3Ob2MjtF8dYFjmVbpDQu4NzSetLGHwZxIyI9Uo9dQFa8vGq7OuxlIa4fUuTsEDencuJH
+4PRtuOzsiqQ/j+/HZvDG59UonsDbl2IuPP8Zi9XsUzshVhUrAPbUZAz/Vx2Xvtjple4kA65igcf
CHOaCIsX27YFdd3dfhB0gsnipPaK+cmmrsCgYGAtvorqZN8hrIhuk8zJ/Cd3DJK7OSC/zhZJr8Fm
tqybJ5EvpvaOY0gPgpy90olMosvkx+NzgwJBijHIDto7NoQwWNL4FjvqfkLmwsybvSar8iqTu78R
lmRsV7H1dFGlXdLAh3P8Or7/61hO7S4Kl0WypkKMIhleQSjFHY3gszoylp/UjjL5T4O1n6x9vMLs
9nTA83NItVW16PdWCjz7xv0l+Y8YfrXa/L1o+YTixc8TJyB9VxZqHFl0hOirUN1yo7GL5sP1nSLf
nDGShkINpZ/YmXqpuA5BUB00SGNpbVerDXjxtJDI8Fs6r5EngPL+1If+/PT15RYjCjEnrev5gvYM
+1ppCx5JJUomkGHWMQSbsc7Uq+mARJyXs/yrXs9dTF9MGnR6lBLsQwgBCojxoMrc5Qu1vLCyQvLk
BqhprBYCXPe3QZt15ozkhkCJgc5QOI16pN5oVpSJhmVD7VWSega6A5uDNZmQYRuekxStH27gx7gJ
02whVAwRqDEuvR+/xWNuGK9R1Xwzlsx0oSDT66fBNFQPFuLd9GC5TcxLjD4/CNeaN+D8nDK+bFCU
4OKKXNT3JIO2wa4V1/nKZezW+TkxtGjiX4nzzlBUF3TCAybUhvzJao4kZXrab74E/5AE8acicLcA
bv/9It+1KtLoV8S/SghgJSjLcP++prtNdGFPpGBZrtwjy2PJFhscKpBIAvlNp9E8SpG/J6DClqk/
W1IHmtTaHFVnANwdGfqsgAgBaMANauDx1ojDOXSr/PftgG411s8zGPfR3ADcgYBHxNL+NiSZyzrv
x+jwrrpYn9HrbF9YvQu1OlwUh6ONGmzfwpy57NjLVZI9stBV0Kuy754MlSMMuCd0pjNx50fJuCKH
h6c04cujhvlDbSxfMQF5XL2yMmebJxTDH20HbMYVlSSpyH1qcJlZSzik39/S/Yv5YtmVcg/dMO5A
IwNEdPGkQ+wBRJ76g+m2nN7bbGkTgEn3IieOKvIce8nmysATAwlqF6etutiu63NFn8XkQG8j2vsO
d5tdurjqGzwiOx9XEZsWeWhdGoBfMaKApFL+aqZk8Miol0uJ0YF00v7fO7zXbeSSNlL5LVsVXPwl
S/JzGoYAYQ6MxOkmfG5ZznqQsqonPmIJGx1QoUYJk6C35S26XS3be/k5j7HJlioIjPbV/pmyS+EM
C6rRMzwzhPBNveiz1rkRmixsZ/vTaxMnVIOweLGc2SQ9KuLte/MaIQ3Ub2fQQ2oHvdCyb4a9DOQA
uUFOxalZjlTY6Hjk6erD9mJWW4KOfTFoQrg1My+LZnsDDAYI/vkTIqcy2Mnq8BlQO4Uw0W0iTsRk
UbQMep9EcUz+O5IrDTIUD9aYpMg9vnCZO9TxLT3QSBm8hOF7jdTxZtCZqd2A8OVgB3Q4OFmZbyE+
gnLa/+hPNkyma9iS24olwuSxtsqVPXxdd9un5zKZexuZHvNBySp/wzSA71VTThmhobU130X23fKJ
sKCsDD0B4UC8St/d4I2c85dxqJZsuiTZW3oZ3HeyJycXDbkV24M8lsiVz443hGO57mCmDV0GandC
VRuTnwwf4Thtt1e5Oa1zlbJMuMCz6QVEW+9E2oeJdWg/JiXDbGTZsOTjYJsSVVMyKp+j+Rbm+k6N
WXl8loKTKKlJ3lBdkcAVMheMAd3ybIJf79QZjMJDMH3/ODowxpb1xa5ZvTZIrGcM6MyBi86VkCA6
hJt5GePuqKPl5S9BfK5pChBpisAP5EAQGUOTaaHjtVEtZAAQMaC3v+GtLXmGLPrdAJCLaXsvIdHX
38YMT61VqGPAwSrx8OiLzXrG1wQ6pTHRs6wvP4RF23XDGkhRzJXUzkR+Fvk5N3MOuGlJmOjVMVwv
8hnNV0e53yU71YVKGLhU3kKSYXxIKkTaImxNz5ZhWEs5mKO+3QygGesYYG7HC70e7S+FMrWQCLTc
2Iv5ZZXIoZx3fI4WCjEBjxhK28KLHjCsOOheVNaShWPU3bvn0a60/q50PFc6LGo3YfisAE27U2nM
4aeG3VtJmHTFOZNn3tGH10/OmG8aJIJns0Mby2c4KaWKuhGm5Gwc7NcK+MxlYlHJtK0prktvjPhE
ImX6B2A5LMAQwjy8SQKlL8XhMhyCdyGPpbdcUUfGbOGsVT2qAW4WcOYHcEnKThBbHiITjHjhy/GD
GO1Pwunzy7LSKJMXqUyFwc/dklB1j86bQHoRyM49vnT9oaFtrmxE9JCWCk+yVOlaUd3LycRhTm1D
twHiQBH8vReqBqmBArNgqq6I0TkaGxzxnxwrM1fThr6qeKJ4JOqNHlbhemnzALDxZgxFFB5E78Bd
ayMqyNGRp2iiBMxhgmGrOUxMKQNiK9SnhX56JHEdruxtJ3Zg4r1fkmYJFYzMiCN/jb/t/BYshpG9
6uAolQvSIj9KupTaLVgFO5oQB9/LHSx2QwCfMK38IVe+xV58FfqEDgQ89vESpYHasx3r7ntbrZaR
F1e8oe9xIBgr34ivl6FnCMXFS8LovaD+FA8xpTpEaF/Or10AeHZTPTiUGmyKCH66ZzRpO0EOFypk
QKZHTog7JC3McMoshAR/Mg9oWsEwQ8LgVN7cNtt03sw7mm4EYW94biQvJNys1+XyXB56hlMDwZ8I
lkmGgkW/V5Xvb0yIIE4nfw0AWIxqWD1eR6pRUXeHhbIcqNhpkENvAItQLmFh1C8VGYel99Z2RKZQ
9cx4K2zLxl/Z1qS86xpYjPfLf3TwmiNzl0vFD2twTxtsH1GMtZL+l7p/x0L6QeFYH5oLFvDrdVSe
M5hoNjx+2nWgS7lXrC27VA3q2VOAhin1QAm46hDIfsCKkpT0DEhGti6K761svM12cnrTOgPp41/G
66tWqBHJ3bAeerng/3EmJ0Q93dPzSyONeRmBDJTWd1g3gJctEaFJU3Go/fLJ5zA1qrL2BnywUXRT
re2KecWCHt9dH9X61fQyf74p8t3tW4hBsfncmno8L/JQ//Jc+w1Ve0Oe+lI/IKl/W76e9PI0hWs2
3eYtwi4qVJciL4ICNdNeCo/iwiwGUHfzvfIJjrrSZyzyMLFJ/PerYRnj9lS9W+jcg/9yRMsG9TTO
fuHCoSJx26dExDzeoDwCmP0R+6Srr4lHCfEBsf9IF5ni6NgECBqq8OFl+GR/7EuitqUhZF71f7gT
VD22h1ji+TIUcaRJbrgCGDfl4Hd//6qKoEszhK/aTbie54JaTCZhUXY2UYFV4kOYXb2HWm47uQzj
2p+y+2fJcTef48CYdxolP4FMx3Yr01JhA99mVBR6pw7wYuF8f7yVFrthTbtuj2slXY3M2vFyhz6F
g7yrtv7GRxO+q6qnbatqYnQtFe0JJUcVbMP28xn+B2FyRz4IvPJwjcfDF0UBicInGCUn+/l7YBkU
BAZ8FyyNuHw2eAQllsPLI48JZONLl4AiU1p9L5uUtOjCoEmW/wj3ZHJZ5UYJZL6AEIqE1lDtRIT3
U9R+ZVWK9/Bs3yPoLVrWp6ZCdDeT5j1g/eHPEyxbjcdGkVY4x1g4B853wiQotAquJH7RPVcBoM4G
ZoHiuZVjWFSSnKO4g1crmJqBqKOrE6fmVaud83V/ZpPvJje6o8yjI8NfMdOsgO08F+hNfsaINsUe
wJcH5WucaXgFEBq34pbrvlcwpFu/ObIIu19mmSYTSnmr9qET9DiGLSKa87ZzYoBtoRT8rgZa7DDz
HltBtf+cZlKq1XUXq3ZBl9+QlBmQEZlfW/LAl09qfoG/4bAtDKBaBFwjX2d9eWi7pOnbgbVw0HqC
sxLl0IxyXUt+DU48A6CqCyYAWPJaDhRbf1CyQMKD79LLaSrQZum3vN03cYXuzoKSUE9DANsEHQBl
eduUI6kleNtjAS783kM/Lw8H6JwWhoD+gMX/3h8MGU638sb4Pm1bcJF25OiEisTY1pLlg9zwP3JL
wuBb9qxVz07iWNS4ZR0iqO8rcHY8k6f2aesdlxf+L9vsEFH/3v8iZ2kFvJrkh6c2HphiRDm4CRcv
dpNXa7tjvA5HMnylOkKVX9x/buU8vAwR9M1+fDZbvWPl4fse8whp9R+pdoSWO0T6MYqk8sC/nqIH
dObfWZehqopXjP9/50iDlnOhd+1Xg/MLk3DbZKrGDuipoYji2tz3P5KSJn+4Xla2U63cVq2dqvEA
1Swb2hWHo/oN5q2+HUy/q5Aumy1Gvd8FQ42pYTZGjO9GFGsJJYoaWTvhJM/+ZVRxsOukfbp8d34s
lvML4Hqj3UQQH0hEn1SqCSQgK9FtLW60L/czA8iLRbV0gf+n69mBW99FRQJ9OzZydKf7+yIDssGN
7Bsmpux+A+qM2ZHi9+/WJeal4bi5zza6Q6zBvI1X7Y3IDxNJCqzQdk+zoLusUFI+8v5TNgIqcD9G
L0d28kZmPab/QVxnXAmmdllNtR9kY1SPVNaNb+CPPmKBbec2y+8hptYpSXHJDnMrCJDf5BReB/nq
FxLcGrNEmfP4aFBD/C7AhDe5/tI8UqaKsGHr+wwzEgAxblaa+qR8EdBe66jh1Fx93F5FPDoklJPI
VgupvNzRBM57PCtDLWCN8FWcKic1H0zsKIl27PHt242ysQOqPOBBfo/khMOraYwLePBDA5WgFVX2
zFNLcoAhabg4m14h3rsRYDKf2DcEuVvMHCKr0teokLkdvYsmX9JFamgqjCEP+d4wriJel5aPvn9T
U8PxuWIy7p7wc+I1U5xpFcTpIFyy46y4FFi4SpiHUK/dEsjBayEouk1TshoIWpPLG3UA/I4auIof
Ah64s8C+Yl+ofGGeDvuW/nKU+QjPgbOKCI6i7cZaLrxkjI9b0C0SXiJ8TmDAiRf1r0e6eP15jyC1
LqbztfM0ZBEnPbDTEuIMdf10lU3RVURCCEBUlssAxf4U1nzTang1EW8M/611XuxyImFh3Gu78OU6
MPJzpmEHOsDkrufVpi2eiMzVt5T+rWrEG+qh7LlrMkP/rJKdCCuZ/vCwx2NUjFcbbfho1CPMNqfR
ApYJEweHvRrpgJ9RGA/c6eKiazSVryfJQX9acf2FkwFrkaSIs+w4H0kS+HhwsW1e1y4SThuknnMl
Bv045bKyumUsUSFOUWPlcVE+PV1iq8LBQawSozQRTqrRzStdC70k6BUmZ8TkFptHAJo+3CS9OMY8
Q/KkNXA1ed18zbd3UaZMTTsIzW+EhQdob+/CW8QkVzFNx3o+GE55F9VVNmzOr4DP3SEbHN+5tFCP
4Ra5MOtQFi9jLLedCm4iRJfzEnZXXwYT1SkcFzS1N7yg5ky9qlNhv/oQX8TmK5nBTQjrGa1ZwO9g
f4GBR7Q41OsVWuVSZVzsmYRKgERkWkFp2EirgGZpoFjmZigFge6VD6B+DtPLRkt0xoN9QjE/pB69
PKDVvklDq0SC5rEaS2WjAKn4hFzzlcYZkrK3XZdyequF1VaR3p8PhPbCBmiR5zc1sgYMovymiwXX
Wl964BpwmlXZLUhxy7YuQdpfMkSE2126eXxuHljtidODNt888v8fk1wrYkaIG81kz3czHa/fqH57
AqtDNamwPdoS3DQKwlFFfdUisHpKfj0jxY08N3nAni8VwpD1gool/JN56JPchpgoa5RvQOrMN1FQ
7KQe1xejcqxqkubmk3kJ9MucWC1OnefNRf7Tio1IN9Ht7HEn71UtkAaE0v97rBV7EvwOjUW1LHkU
LePSd9+3zfJJF6KqmKZRm9pjbUzMmv0I/LDYnvHy2PSbO4YX4eM/GUeT+oSY4aBW2k+oykoxUc4j
sciZyDNhY/tUty1kGXG2GTL15UKL3MTj+5X0F6D4hryWrHlGvTF4zXHbV+NSAfzxpoRiuEtdbBDa
vXy7b0lvvvaPflBVV+00rrmOvGPMOE1GL7i+8rJDJbUxq7gS6LHggLjj7U9rmgW6KhxkzxiRylWz
owpsEiE/PoQFnkO1VKBJYMuUuDY054XpHrDzOeqdsBqnL4xo/RP5Njzww1jPjk3uueqTk84vXeLK
XfACbyAeaJvQs/gD9FVMGvuHeLSP8XsDVForCWj/jB8Q1fOWi1vIFH0Ervt7bbRxXPjiZtDwHv27
4+SrCT6g8y5DIYuJBXrD2a+u1uwcrNFzw8dmGBQauNGc4THxBBfoM/7MM6z5Q3De7SXyEs/n9Ktw
dlUzztsEQ29u+Hyv6ykYoSSDkAzUTBOIjjsKDkIclwANYUj5iLz7j3sIkv9et0VpEJGLBapg8C5u
KVwVW+O6yOummGcuHWkyo6ITg7Ih67MERLmrWCzkeY1Yu1vRrKpL+AwqDQEQfndnwzm3dHGzmT6H
a07lDJR3az9aHAXlrYUSofdUj0rbcxg8m7IB2HnClpTJKWxN/Uwarj44b82j56wNn3cnduQKT1Yf
Ya9EDu2Ci/ad9qdRRGf+3Y/inyKJHJ8WF2XkBXlbzyDF6otJrdOHsTTrjItdKDYZv+Uvq4xWOnEz
S5L5G/L+g05FnREoozXh31DJr2U2QutLa4Uil1+r54RLNBP4IP8uou8JPMqJAqu7wLwJluxQ42zk
yMmo6LnXf74iMzrCKu2FBea42HLf5BOR5CvOvEDUr2TjAuc2G8Aluz3TMJlgvphP/GwnxqsjjSIO
e4S8UyzufkvH8her1kn2/btArw3eu9Xwf12hjFicIdQ8RD+ZDq3S+iGd0ogvVCUh3rj9gg9rDuAS
7Cl80nkJd6DpcxO7gjyNXDQGpndsDTIhmN+3ctHDzr/FQh7Fkm/3SLFnyt/svr7wI4C/dXOgVjmX
7ty1EGVmvx4JQ4arkG2jBUv5sJn/zvi/pntuw7m274Z/9w0wUnWuHzLplVMSN7x4ExL3eC+ag2Hm
nFqC+NpCYccgNmat6HYhLJ/qyp7298cU/NKlY3NcS+hRzfGDbq7Ek0nP5zNqZCXHd4lr5qJuiZnD
6yIivSVBJ8+ujiav7wBVgm8oXlWkLHTxz9yX+yRgV/Em/61qncHABC7H43VV1zVTp6T4ZlrA2JLx
a4TCPasgrk2uv3F9IDkHmggUsXdroSRS4YtIuqv4KIHk9V8FqTvjMWEM9OsoFmc1xPLHcWTI02O8
y6NyJXK1Ju5K8pCumcdbwob4kARF4l82NWd+GdX0uCuiOabjRSDec2ap4yEOzKaff8FdYSWM08TD
siAA1gDvs66ZN0l0Q6D1PfbnL1HjeQN9BFuQUYRsXrBa8PkYCivpuwCbLucIPHsQXz+KrFAMsa7p
O5zxP0pj/5AxPzpcjr8oZvl/OT5ec3dCp7T1J4gcJ41NqCfDUciSM7r2u8E6h53UHgcUOWEcqvWJ
htkacPqoHNSokO1XDPWH/UgHIrdcn0riHMQNoPztYaZc6ocS/45I3FZBiBglUgXiaBMtelOl0DLU
P29PjxHpZJm89dX8WWNlZq3i8usfsJ7lXvDoXSENS+RpalJaT673+TNi7JsLkPPQY/ftHxXYXmJs
JKo4mVJxv2oXSY9VMvSgLt4JYUSAUc1Cm2EARGAslC7TVtt2g8aKZXbiM2xZHMfSv3036EuORht9
I8ly249Q0bZ1VLtmdIrpugmqoIuK/JXlp0VRVN/X9qNaLg7D+lQ18W7hXd2pmHc7CHfRe8Pyip9E
Mdn/8KF/A3V5GTG6JICdLBBE2LXHwXLKF9Q/EUTLmMcZJhMpAMPIMSYxkHxmK834q2oTxq//RmyC
fU/1kB9CqZlSyLmQO/WoGYXG1/gVZdmrNpTgh7Fa4KuQbloyzKlraOzeDeMNQm4INUWvTqRPx5Id
oBfJWxbfQbqbVfTzqmAuIZp6HCX2Azerzlj+ejflqDEIgYTq1OdLqp3vkQ6pXVBhtQBlelt8zpJg
YUvV7zGVJlstSMI7hMfMWlXwUPeeNu4I0K49dNP1Jh2rFJ/LtYfM1AxKmRa8jJx+Qgv5PdzKAN3r
3aVO5HDlR5UbIgQLgBuhAgsUq7h2+6g1X2KSpEKmKuxdMwVwjSzRWp320Q9RCcE6QVD9Rhrqe20Z
wmNVzsK+L3i/ASQj7jDk7yaZ4FDbj0P5erlM9e/9MEr7Kg5OFBDPOjKomsnU9j5MZDO6Um1zK/SD
cg9FYNBbTnQiWmcHkKS0FhsO1xzi0mCtqBAivq+EhlFmFi8aTKQmHkzppDNdKgkaKkyTgA1/K726
ZvOkSC0II3dbPEmFsB5IPcCaX8pxWjYkPwAGTshfSWQCh5nC4AEcNtZqbeuhRNbldQ/rkvgBq2KZ
peZuJWucFaCBLUVm/W7+d7wK7bCYNfVWfiFURVT7KuFrdo5aXx/dtONBLG1v3ZmOpt2fvVfvuThy
B+AZ97oO78/hGHW71mLV9GpWQwpwn0X9afGmNi0MP7hY88atYD9O/YMLwUjBAjwod0od9x0rx2dS
2KjdRM6V+2NF6qBCd/DSBKwFKQ2spUCyJPCmaQ6WDMFjusa/0TVzwC8+GsaC7equUzYHzAK0Jco0
DFuiQLtg2tc354dgWndi1B1Tf6eIx8Clw4wglAlZIQXPCwH5ZHU15Kdd3ra/bJ1qjYkiCtSE5Y+U
ZKASR3pm360GIzDjt2Su9jsNVWTpIC2rhys5+h8magB0q5ZW57IyZ/Ygp11IuG+JFJCgpjTW9qlf
wrYym2esThWnvwPWTiTssEZJC87J/UWf0yn80vQHDvqdsvcWbtypeLP2YvqnnXOlTkHVjNL2IR0j
3kY8Vpw93w31Trf7Q38eUZ5TKrYsPCNDQn7iGLuGBRfKVtTfd/hKG9t+swZnMmk8qqs0Vbp862NW
jpOLyx5Op+2zgLgxeMp/lZRZGweSLJskwmXDoVGVCNfUKuc5aiX/Q4A8HMgS4NFt5DvW2XFf/h7m
Vb8Iw6D0LOxBm4GoZLOjBWaFIHvITx6RPvhedY4OlYndVoRm5YO/C5ODPNcUf7UgX6Q8gEwGDRAz
foNCEv3QB+W3AWjzKC+4ZmQmVswQg5JMKJ3rQ6AcbWnLqZreGCgafUhb95f3p+zVzOiPPiZUQ4k7
dUfQQ1VFv4zZSfp5+7TFTfObwKnDk5625YOowMKoEyIBArt+11Y1hNMFg6/XcdJECqVqK+bKM8cp
EqW6QiAxUAZY0W5VXTKs8ZWK33P9UYUzEATx5hxE9BPfcdxoK92ltmfQKKQ7n24qKDX/Hx2pQvNM
wZ9kCMFp/qq383a7xzphswoGJ5DyhyuV1XIJe9SowlCrCpjB+7RS1bQyVKWGqMf+qiyCD2lc4TQY
23xYUjkVMuAHB4I8CUiFsofJUMVJE1RCsFmRR5WFt/TFFY0J+XKlAtkf/nj1fYAWGQMKplNgYkOn
8B0skAYAxAj9Zae7orHeSyUMLfs2/aqWOPg6ee3EszQdRUvhYX5wztwGAjKaWmQmVrX9C6CgXR9o
KNlpoDLc5f1h3JOx+giut+oBrjO2eqq5Pts8rne/fFCIzkOzSNShqzyJYd07xtpdxstx+0u50gTK
lZEEh13KBanzDWh/HExwYo6ejW0k1JxVWWD9+g4gWSW1pvhWXC1fxwaauR8/w5SrxX9ISSlZXpi2
NDFppeqppgBLyeYTQa6XO/TvkY0UxZ/91U3L1bGbLBM/WmwAx8WyEZJ/GTmY1Z35BUvntR7+88ZP
cG7/ANVIBzEQ1i6evlSGC+6Apl4A30CUokjlgZFJnhm9BDoHhu4bJFEj0hrwEYgao7qHabkba65h
x/Y8cbRg4djzP8/RT59/EMHPoIrRgHmh3mNK6fIYXNiKmAbiVxQA7KoiPwpi6+LGuOD2vlZ0Uyc8
6+cvKTy6PfvVuaW5I8AvSlHXNA14wavXpv0nljtFaPYHptulJcz2+up83Tnc+qdckEG4bpjXOvUi
nW5cx6LWDHu6SP/dYVnsjLS2fs2Zymqfi5lhv4IXHmO4CEFKZLsZo0uNzPhISmMAEsXli+PmYclw
DNazp0YjPy5mKJOGtpbNJ1CYUs/WjuLmdQSydUfMtaO40hnZLFVvh0gjQxeFbg1z5ar90BU7Uoor
+jqoLqggp3X8kgiBkMb1+xdglcPfyd4vnCnLJYdPPCLuC6eu1c8KOuoxnxhdcg1S8I3cFsnF4whN
xzahVpA4VLf3CWhdplbdF+NdCPw47if2sRExeWwZ9Q9vvM72UPl5fll3r2ZDanRWJReT4wa76oA7
Xgja4ggq/41hd4LKn/GmNQSAUCxDMcSKtLGXzTW4e1fzYo3mnCHK3x6o46+cmMbE+ef1FikSnsTw
JmuKz7PeifH6huMlS/T6x7A6H+NepQMZqSLtILjluCJWUPHZxD5UXm8JR7kauBI3PvYcFVWXJJx9
Q8tXmru2OEJIjBBIRfuCmdZ9L20IMTl5APTDpkV0LuickUergY0P99zlqLSCcMSBJBgN6IAjegvx
kc4opyeNDRJFRkH9EUknQ/DDRA07FfktLK2IwQWAVCwpc7MORzdRnTuNxgM42Nl7tqjiDeiv9+B7
w4XFaczVgIudxiTA5v5IaGsOiSz99xA3JLJNEK1F20jhBWIRnfpyiNjZ2zrKIDPjtugbTl+BL1e3
hAu1keIAH/73ek754K8oNJecY4RMXOiuM8iUT86qNDLHARa0Yz1Tzuq1DBVsQN6AgG+9hMRl4YMw
McKBk+58dL4SNw30Py+DJFZ9Tmf1ZBxcfKiC3I02uzgqzN99Gx72Ymf1nOYQGGohtdnqj3/0DqAV
BHGwqrDT8BT0p1FDZGJvBdDZWihHt8HfGqnxkT3dAr5GloDSN6uEYL1uzrnmLviLpVq5gh5dxImX
D/nwytfmgnbL2DnuwQka4dkOS8eIs2Yok6gZwa6eI025oil2zBI9Vf1zMm74aipS6B6/Dk4pGOl1
ZcznikNHihQ/XeZlNuTN7VGvQmAus7dTJvXstk/teKhm4aFu1SpjLbllXYQ0mpV1iUZEqKBOWQMQ
jwg+syHhueRBuKMu/XS886NHjgumBJrIJVFsmMzM/YNoXKyYkVvNhfXWyJEuxbmAcab7nb8pmJWs
3M2jMJfBlNHVsNR3MOUy/nlxjC0olf5bV9LjVHeQnF1MifFVNhBAxhYQAf8zWpnFDMmSPqqT68Vq
cg7P9U9a/1doaufYcmbm5MRTfi+n294o9GoXrkDbh/bpUANoJsRTHSDo+SfcyGRcQPZAvs6ZpwDQ
yTrwmCZIt21Yio57rOPbqKqxC889g0VjbPFiJ8oKIYjzwHXFPrOC3o4dSCfxHJ/TfRejB6PzbkQ3
3PU9aGkzs7FIzDGgsSV4+ZjKZAaC2VmQLrdn2jP928WikfIcmLhmWDEmCZP3IbsHVF4tXSn0joaO
L9Ii5R3+6BrItlO1q5eG256Z1Ti0Emo9yH68GsLcasefWdaFsU/NyA9szwZrbmvrpTQ6bdwgyjR0
ellPdK7eNbto0Dvn5HeYBj+ptl9MvizCwsfQ8LyEYOIRMOit9noTb0pU562vamHfDPTeLYU/BK1Z
JlqvdMt+rzG8gm6X410qu9qs3vPO+nmdv7DKS+IRQ5ikFh8pKW/GVubKAqe+Kue+Ap/BarBU8H0Z
ded0QF3OZCaOyf1QfolfNWlylYcXH9HqqvEAVArc7ZZXn0upEHAIHLJLhaHjdVVrd8B5q5AXWm2Q
kjjpyFRILw7HgpSA5Sl4qd44knVO1tSBL05SkOBy7SBJ9kqJOTaEMztt2VzAAkSZmpK2VGJ9ULA0
meFmfeIwTlkaOTT0Xxr51V/jCbBy41cHqiuRr+3Qc0DuWjrG7Q0ep2uutq9DQxQIq7Qw3b+sxwbn
BjEd+mNeGIyrEiiMcB3vibsOTMr73i876t8dKjzLpKkgOfl60u4J1vWe4Ni+nnrroSKh++gKUeaM
LbN3rncyUuYZ+yn+oLwsLNumu9AKNWZ+7xdGAY/z8wA6+Rc5+VRbFsGuDKvIs8syXZsFqMC9sI5x
JfDkD4p+ln5PAv9C6+ELK5LMfRLfbqBq+ATmeI1nqhXJCDdo3RpeeDuyuW5+8T74h+z16r8P2ZQL
t+ezB8jlBZo3/8K8dd15ol+PO1R3+dwwOLIzbHBEPtoxGgnAcxaoWpNbreY3rkOC0k6GKunXOGfL
ABQTWWFZfw6GHf/kjN+p//RgqFrbBw2mivKO1hKdcx0Ph+6hfRiAvEnE1LKalHLSgoAvQewatUmK
WHx/jt+rlmc+4SZN/yjAtOeZSoNlrTBYfcdGBsRnIfW26TgF8yWCuV8ztADFT0krhZ9O6pqUSWNL
YmAzWbiKIjM+Mtkd7aZqmgYDnIchVvHi5M/bCqCodoWs6Z7MgbNoeJvLC9Uc6cYx7Wxj6WpAgjEZ
qqthsZvJaLok/xrMrg7hw58olhwo6i9o/LekiU46kUMyciQZV4l/MUrKEe9diJDkmcgneVWTaJhb
JmEF1w0yAwOa42G5x5aPJMTSz7bkKfgtc7CZDVASPHWOXVvjgViW739+vm8kftsmlTvpCRjg/MFH
Fj3Q/nz6tz2e7iqGSuZOqDh0sREzPB3DNSGIQ4Gtldzp4FqETpTBj8HZ5dj3Eefibn9vyW0Kkfk0
BO20q84l0NNBOxYPTYf9pHKFBxODuB/CgvGnU4+UyzBJGDr20I3CzBKfvEUovk6B8WroDPdYQbTF
lMhFDS+yoJbRBIlGUuDYC41UUAj458lSKz9fvwG4B1ZLyG7S793YqykI8CgSEa6NLtZJF+i2QEvh
rO9v3vOiryDVkD20EnAIReAjZ2eYC3qla7jIXUnRq17zVgbUNunrzdRObBTxxYdkMpXWqKZk/dwo
tI199L235IAsYOLxMBaIH27f2mFzwHNDqPSgMzFEI4InyENROzIOPZnrbjWRfu/194QgjhDGwX0X
jafG0P8Kfx0w19jj6/QcZae+vdmbo+Gcd5u08K3Sv4SnlK8YrrAW9Om9Yofei5IRJd0FunBiIj2x
a31PBJ0YxyaYH9DUL7ZN/J1GJJdi3S6S44j3lpSSjaTaQUuieqpW6tk84JxRXYy94Quz7IA7FpkZ
3Rad7GLeAMFBSENNSJwOt0XFKLeAmgwrwhG+dzs6NyW4/xdXb9PisPnIFG2xN76WqoJtodKDbYys
l/+uz3pJGMQyhKdLNKN3aRxtIQbRN0o7/y6wy4h4xSBRE6gfHKa98UrTiKYXcG12PR/r32sK6WwY
JIa5qUkWwqabaBSuWAP8CU/pCzBZQRudaNTQGndN4X6tG9GdZmFRNZW2PFzYltDWOKDufiL+S0nq
Oiup/jzZyI45//2Q3hgoriwvu0DPFx4L1VyMs7sADA+ou5n4REnaN2Hy3Nwh9P6DDGaDF4NkIGPV
Rm1YfaIrzb3B4nElI3PjyL/7IOmxVM5Yb1P5kVq5H/g8wbkDKP1PwqQPa4Ls35ajgWdrjXTofPxG
XvCzrY/E4epm/8B+QEcK8AYodA3xSRJufearpo4bc9Cvp/+dpjPR2FZMDrlrjZyRDWUlPaMkK3u8
KLiVjXTtJaJFU9VEvE7EUIMfZEFvw3UUF0sUIjOl++mh1bYJjqUZQJU+Bu5LYqfcKvA9uBm9VFHD
EaUm+wAb3WHPU8qe3pMu/Rt5S3l4BN1yovTeabA3lnrYDfzzxdzLDhNvY5uq1E/aM9lszTHCQ6Ru
AMaD7nNmDP/GFuzmJM+KhtcO4Qut9HATJaYnV+pUFz7T9xvwR3vs19mCWu5d7+upmdN6QdaFYsl9
UYQo9KMfbXaF+j63A7iwCrZ4IHGUryWKp/SU3OSKAsuTXwVhfgX5RA3abt9xQq8q+VvkZkuDAEnK
z4wcLS8KMSa0ApzHxMXFpb6t/WENmk5xBh7eqyyfp7g8Jnk8xGJhFsHeoOGihPw37NoGiB2Hn+dP
cszkLtkOdGDoqFCCQh8OpzSULOAi5X8zyEy3KWNSt1m33BjB1fkMo1CGQ1F/Z7rZ/imdfN77OZ4C
eO4xWg1uxdRFguuKcSxiMFwDYXmvul8rX8LI20CGbc/Efn2fuGNY9tmTfc0Wh3JfLFdVkeENV9PU
gpkMI/0oqAEmh+vmLkdvu0bygGm9ZMwptHuarsbl7PLEXWWdyLLi2rH7meSwtJdzWb2ReqspR1rK
xBqOZ1iOJOzwM++ji3Wky3eKODQl4bmjLdZdVCM+Iu9Ek2n1L52HcdHHwa2KK/5yP935MO2QfkfB
6QP68qHLuUI8+DwznRFlWAXtFZpZ2sBDd97aNT8sACxoUXNwLciWpC7Eb+BjeMPZZ/XI2VSSafym
m9jfrUPDkiTvuhRHVO3bDB66qYBLwLIPtzwM8t5Z08jgmAIfQDtpRQRpi/7olUOS/z71r8aHCcBr
EPCkh4LCrmWEM6sOkFI5rVBQYAI2zMEQ9/kQKc5DK8Q5ZCm03SpSvrJ8r9jII4T2NMwvG22vsFSV
ml2qw/ggpfXEl+fsG91/pOqFOLaeyTqcmibIM5j0+syI3tV78E2EuC6nQmcZ524bnj+5jGYGodTU
c9/tPmG2UdxH5C/F8ekGcgN4x4fAyjXT1fubYxhL4ZS+Y4HvCNCAg0ej6kTCt0wJWUhIi82PN3/8
5Z2rE80ORqMHUNlWoel7VCDyi4cnGxWROWsN4qRZ1mZOWG1XZ6CXgdM3LODXLCvg8JZvmWMbLGbj
o93mDn9SDan8tlevzrXq8PPArxqqhaRIM9YBWAc9yqdzsv92+6z+8YbnYD+RPifDGphLdyzDvLzC
sErPoNP3RRx2IsJz2N7GPJCT90GWURLvTlumh/DHtxB0t9KY9kyCgPCay5t8kDLlzzJ3QRha9AZr
c35EVNPUdbwFu8wvelwTqU4FK2JPSTMG5hbqntPNUe2Tj1WqXXJ7qygK8bijzOtNbQrz9H9Lx3vu
fj53a1nqz4RO2grl/TdTOw0o65fIw7vXxHmDvScZrdJsYcZvOV9bAT0j2Tc69e2GmhUtjfSCrObb
aZ6yZ24dxC7ZzRGK2nqxVRcfgrjw5DOchAPxndONSOCJhXFLGklco1i0nQEwzxnSvuH+XmFY1xgC
pORYiJEAqHSuymtOOAr8ws1CZpueiuU4kBePjWRkRe605ulbBAHR883UpAUtR+wlk27FVztJraOu
qts1+y42HLBzfxjU58947b7wSNQuAB42Yh3tqjetnCwmuBOmwtJNRiGlCX3ZpYUpexnPxiAl7ikP
DWKbgbtML6dcYeAn+LU4BscpP98OmJkTD4OrWwhScM3cLEKXsxffrRoDDNgmJyh3wPgq0PirTs7S
wsrFjWjdKPtbM3iTkoIwCvthrRlv6UDaZtZYmsphHlGAHti4pYTqE/htOfhQHMHtTAFh1qizLA/H
3k54ZcC5PhsqJ4LNv+eqI1/fj3579uQ6du+HPvlu5Yxy09slREVVyx2LnomTDu2bR9iL3XldIByl
9OMB8KFeMSl6Y20N+n8sJenWhgEJ6BMkT3hcN3y1ATkZ2p22VhhcEq+uzzpZiutBvlj8YSouw98s
D9FWbqx5xcSsh/nBEFCFxf/NVT2c2gSNRkRnRLyCIF1r0QfLrxEMHPCPKZ8Y4d6D4njbW5ukLO3r
+8a3ZY8nHk+kJ1rnuFkOX78hMF/vGjMQ7TYYIUQsjC8+ONNHGXWnOG56xrEHjFzPlOPQANKDR85E
z6OcJnAk+A5vZBQZr4L3koLA/Q1FO6Xir5BQQdKAIVdK3vbo1KmPU9mQQbAn7cXiHsG8wdk7LTHI
MCLRbDRgXsmQNmbYm0GXnxfUpcYiHU99KHU7qovvjgBXh/C0L5GamG5Nr71/6DpTwAIukFNsL7nY
pWV95+sZ+UlI4znWoJD1LzSp8JRw+bzLKuITht3wmEozxpaltRZLdFvAa8kKAS2Sje3AcsVpo/B0
AtNuEesqVL6wDbtC7i07yGcH/SqPS1bTTFvala6tJD9UxIV6tG0M+e+My9yMO044ImWdVzHjG29K
oZNDvGN9UNxNC4COph0zYdR9mXPHoWwErxX/wRNLDdWVYtydvyVS0wy705cZwVjJHMrzQkQJusl3
V6vcmsWuE5B5mKvg2K2KCUwyBgt3KyrhhWRMLNNHVnv3ulW3iNS1/zhnEs/nPgRdNU8RypckMsJX
qZAlSECyQ786R/uhgcsoXpJEPn8iDFkxJwyB+bmH4Cjtv9xh2nt6xXaFab8j+JOX6emt29z9UTT+
NF00+NLARYrQ14Gs2XwX51/2uZWx0xuRClj9oj6aU6SCcyvD/rxyrpqgY63uh4HKBJkK9Vuaib0V
UCfJNDq02vCZAvd1Imt9sVTX/MPO8P6R6waQnbaSgQWx+VqCWPmTGKNDZ/Xid6iAXSQphzePI8Zj
Xlc+hPh6HYMCYt6axFpecyCT59EPC7e0hepldzvWRJRETgPsqUs7V1/3BYIhimND32Co5xJfMGvL
qR63I4MU12KW92yQUVGeMkVafRqoJwHkAZ01Jkd6lRS3+6/aelS2Ifv9tS7mOzIQ98mmEzWj3jDj
ssVyqGZrFE94v3wI0FdYHubtw8Sn1jqV5+HA9evUiXmDyuXmLuJbwfbXVJVcA1okAGdMEddGfF5C
cdgwHALLpKgg8lztGoyjrZ+CvKv9+G48HiXDNm3vNcbuS4opLDGa7LP37f7ozcoVyok6IHbNp9QE
HaPAdHxP2YoPfysVCHaBF7XgQVqjBJxRjjXmJsKs7vHn3TCRZ7fF8Ysk3ABudBevdOt8u82jwmJd
1ARIxj21lLM4uaWiIFEnWfF9NtUMpdpLE2L+dn3D2gwq/5mxPurH8IAkVMKoybdgCRdzfjHGuUC9
hmgByl8a4M1/jMSymTQbT85UJc1ijT8KIsU5iERg8cOCsYwl4KV1TO9kr3b+FnNLuCO6SK9WefKo
mnv5ikYQYPruDDfpsIQceeLrcPfUVbGtcpkFqAfVWGjpTNMfQBBld0XqVE/02cf/96oAylWb7EJg
FoPBLT4FY3Yght6tsmjxnN5f2NGUMctimOYKqtJ/TdjQ9GAZzOJ0/3jVI8w7008TfN69NoknL4G2
KicxW5HtQb4/n5EWhHyFSc4U+Z+EZjoie333nd95AqRkVx8hxXHZ3HptuNf+By2NIMtN906IjHL9
txOnn6kZ+0OyFvVoSTdU6/2PBaHdrRzKG3okJ2nxSnJl/2S+fII1AokgO02nIMNNwn0sg/bbhwOy
PimYCBOjTqyVg2XiOOcug1rr8cn2XfjSJxMp/mMbiG7+21Ri4kFlyczyR+FDG+NVoByp/OFknmEz
Ns3qnNC1d9zzUN6nB/dJf/5sOHB+i+Esdu+udtMntOpsNhw9iNLWkpmLs6fKGKDGdAVo6Bzidv34
QMn6E+VTzl8oYM149XLnw8BkiwF6DevC0PKKLtWa1uM9ycFDGqcNKkZt7dB5EE5SGzuE6YLISpWh
c/KFXb58IiRZ16qjnZEAZSmmbq2m4TolEIdgtmHQ7DmZBJAqw3L83DJ7KCLewC6pPeVdSxG126N1
69lNREGp3YkoqOvZ+VxwPv7A2IMIcwmWUUAtTmWlNIsSp4TaFx0r2GikOm4GJXpsFjzNoCdykYC4
+TXWWDlfUVBZwgxF3GJK/Q8r20Dh38s6DyU4TwglqslsFu7Yq79/HPTOhnk8U+AgN5uVGrv1aYsq
KvSJl5/b8BvFBRNcyMkXQ8BNGz2ziwpcU8I7ReS1FyFRCxhTL4P14T0RUiAKGtY6ZQd64ckZhjMj
u7Bi7CM12blRTfgzahP6Wr9IWdjH7a6EHbQPR9KZoWUoPT+33TK4XONlcqbCPDpI9CHHOVSa/lvT
triBLJ3mKv+uelIAHprDlyH+PUF1utjK97mSgABzl5jrjvLNxlDtdKzSSRU6hX24oPjfeQukRf2F
gEY/MQ9j1ssl8/U7GmA4EgK/6II32AOuhhp2DF4p9NjfWtxAyXuTSG1jXwiHsVZ4czc/oCyHTDi8
M3flxMB89AvelL/5CAMRJiKLj0ejEqY6JofXBvMmi47KhSekl+Zifxzv21SUIstoY1S5Wh6dYFeE
tMz92//jshUTja4+rA9kJPh6g65eUczT1t6kPcqxBU3VRjzcoVbdottqhFVFZKXg6JuICUjpugvi
PgeBxlM6XRn7LmoOU9W4vrZhLs/jcV1UeE78JSitvcva0MQt2DPUtf4/MHzqTRAr7eV0UkW03NY/
pXl7JAR58OCFNMbH+JckKD1yMUAXBHvNqiIsnEJR/VGnLG/NoEdwQcsoIHYCFUvjhRZQnoHxxqlh
uyjte0sWbDWPwG5V3AmMbI00fkwTnH3sjnPaQSEfHmsKiA/+CxE5SdAINOdMDNLSnEG1cPXhvIHL
2/7PJn34zlTxFjuP3/OGLeFUIf5BfbBkX86oR41ld0CIGkfurqBHoUAqS2QN6uJfJAFTcrqJ+sT6
GgoEaisl9aw7OvuEh2QGU+PEaoujF/JIFrfjHMoP0aTY2OIFfrJ7quBk5m4RLMKu8K8s57mXYI3v
PKLE5pxV/JzlDWKFPz4tA4wzIwIWw5v9JN4obo9lOFcKe9+cFqly7ZdHKn5zvyk7fuf/ParxDwI4
NYdVwiV7ACYTWG1QCfO/iIwGgAnC30V7/EBzxAfXaUSr45x1Gi73v9BJk1qfPSD9mlW5VN+rhlAk
8w+Vq/vFQp4VawRoGPBq1hAlhyiN1mrvaM7eKwCOmJEvrntQCWv/whHBpOVhaFoJflzib/w/13iZ
rhA8xnoN5tHGpKic6a1HsmRjL/FZ3evbV6QjZMK1F4/X1ocjth0BvbHDVvENx6hMTOqxkj6ePWwp
Y/D6eEvdzL3TMjP16HLRaCqmqJcB/yGdcQIF11TM/MZuUsnp9bfoaa0wWQBIkZeluNDLnuMNWmQp
9nrsjXRrhWJN1j/NfQHCHqrJ7a7dkilEsnWPcTaNNMNbGn63uA8R4fUI3xri3pOB3vsku3yavxmd
1WLhBR7LZX/sA8zrHrlbL28ES+LN0JW4Daj9bmWLL85KmOnjROtTFGxSek3F5ATI55wi2yUD/9op
gm+hYsE7Cx+HGbi7fWtvhBBOIGwSWLTeITolTe4jRukYsqtl/ZJr2sC79+35PT5aET/gf1m09tks
pHn0NG1CYJcRCaqUomUx+Qkka0hFXni0WsfPs1O0GwPckZN5wykvxGEhdKW6+MOLFObLIg88HEZe
gCgysZRyW40FKinekrANW1BvcCNpRPq+U3J2CwDR9cQQzDoU+07D6eX07K1KKOg4YkgIkUPJzq/q
kWdjUVErBb1Z49yAzmBcohSYci7LuPFvzuKeYLUBMT3teSAkK8wpDVvAJseW6LSs3SHIiY/ltadK
4bWuUJgjCrKFyZWQqUjpPur/La3dymdW8tUt8BERd2hgclbozKVMYVZaVbJWZF5aOnJ1JFb0ujvo
Qc6KZKN+aLnho2V2Byy4XPAJYwkQo/cnwuXtaD5IkVO7K3P2FMPMoqIB3S3DaCN4Ht7bqvbfBjyV
ZIg94um/gEQwXTM2AfUoo+GbZFHqNdXrngA6N6I+sg6Ne/6/elh89t7DZMJgaTrl8gQ945Qjc0hU
MPGo3lSJWQLbadT+TycjemX6cJDz4MfwAhbb97KL/Zdnf/Y1tHfbEGA+mq60XloDmTbISPwP8MpX
DPJpOOJ7lgLtGacocFIMniT+9RYsc7ocIvA/jh3kwTHET+2JuTam/0uZI3ddkceoivZNPwSA9FOZ
7Yh66vzB1VP0RZYg6i2U03V8jYENDq/lcMvpRNQTiROsw2RwbPTT7HzBf6oOFALY2fh+uIhGzVlw
7HCuugfsQ/JrtnunvSN7SLB/HBEy3LDe4F8YtYe0a7hXYThS/JyL8CUbmAMVqo4dJjiPxDS0rXE5
XWP9e+uZcQ7b/MhXzjBuqhTiqVX1Vda4haNfN8qd0sh8sUoqLSzFTMCT93oSiQQlCqvUgLpdjbs+
DzLcJeF2cac12aJbH6TApkJBxEssdeky7eAn6T4fwiy30S8NCiKB8ld5SWISTMkXkX0mRyjkGUy+
u24/VeZ6RN5yMTRmInKH6r6PTeEG4nmmAwVv576iUkzmCjTAE4vr97DaIvvqhqHTfe+W6KwMLUM9
QUEhSMsO7lHABArxje+/wgRgcxzM5oPn8i5HmiQ3bo2KtOLQ+NFrwndWU5akp08GzbgeGE3GOKBd
rjxCgxNauoGIvTd8dwwfFGFCj+vpzxAaMRtnET30onmzY0UiagZ9XAX0Llhu9eOiWWlyiOl3/jUo
80gyDx/NmgvGAw/9u2n7jAlagPY+Lg726m3xO/cNUeAK7Qk1KcmMMs8Vp7iBjwpbnBzRdQaaVPeB
7vOO37nHM8Y7X92iG24bwpDVZ5GOt7bErz6myaU+/PzKaDh9atNiipQJl3hmTDxW7qCI6huDft32
xgR3nUWkgnuMrPhWWqomQ9WbO/g5qNrKbm76sttZNTyaUjXVVd2Klw8Sp6gcgIi8GOQFCHR5w+ni
b/fGf9FOm0WgdOz/wHomjB/dbPgJasRcoqjE2jNW3IzMpaXrM2EwjK78Uq7oZyLs5lb5YbkycXuK
mw8BPbHUCPifKAYaxRu3W+TPcRpksy994YaxDA+RyDRGwFi41vJsnMfsrZEr6J+t9DksReRDKlxr
RX2s20rjbaWm+dZN6s2yyOUYqnTZ7KeBNHYYeAZBk1V9sgawx//X764VJTN7Yrd+Djg9kmhcpxJj
Dla38idC8O0mnG/25wPLQbnWBChrVsEJ144aKHTpkzo4N+GRMVaCnoxDrVNdWUECiDdASihEYs0r
rO/td+ShbJltC7ZF7vXNccuP3AJbjp9HZDqZ45HRSAB/v6uonfBGswBB5PMSYxS0QXO1AaqLxQZJ
AYqIZPJ4W/73t/ETwKsk86dasTo/eycWwr1fxSLbz+q9bBicoRHY+R4tYzUpkyqr/PH9vNFnusVw
67X9DaQRKQR7fl61ThsGE9GZ6LGR8UeIkNB6Nfs/SNUHhj7AXTqWpTTFeYtBEJucNTBXkE5F1TIu
OFQCNEbUKhZmW02hgxgvpxA5kXYV/C1VUrminQSncK+e9LPjYyHklmWleoRWrc+vo6w6Jpcy0C8/
N1PCnOmTtOsr+IQuqsVFkw+28qh0wFdq8cRz/PLsLywXviRQUP3fy1/tiDUOOAY5J0bGA6nQ0dZH
PK0wbw4L/3G+srdTn5J5XgcnUA33Bd6x1lPqtGPYcuvsHxmln5g6evdzqYr6yZ+4iAu4E5g1OxfT
B0/EiBOoXVn7wI2mLl9DG1nY0R+ae3FHBz4Ib4txgIGOOXHEz8VFY+L8ScPOoWSkcTaGaWnrvfmu
A1T9Qw3bkZAgCQC1Zc6O6P4tschP4jJ20LLYFBz+p8+z9Wjsrdep8uU/RHHgV2hfwskESh7aMnm6
IR3Mk9TExu0Z6T4d06G4DbJfBbkYENENO0FQ9EZ6meS1noFPVvQMOIyV6vfEr6oZw+U2PV6z7mVr
uLEsE/oSt9zRuO9KHyY63+p7miyYmtqXZVD2cclA+gbJ7GZhYNNIBqRZ0GtDc6V0tqa2j+FDFBVA
Q18HM7ydv9M3zN6Wua94qn6qfZ8K7dVPCPXdeVnWl67wOJeWoT6V7Q1pXi/beTRB4J8kTILNC/u+
qo1uZGk6iGzF/mfDgmeaqvR41fD17gPmKSiKLMzXff1DjQFCl1WYJtAKI08wUSnE455Ihss7uOlj
C5zho/i6gwUxSvRLdOV/mn3gQ4Cq7GSBuzIaniEPfAXnnMRo3IdXA40w6HmGNtRYJGoRFkYi2IUr
eKBtfDknv1sfM9oYWZyxoON7wh36hQVisGPOiPyuD6OldDAC6ECFZtVlTr2pDyLn20nrGyuaiZBd
1tAzahsIEnT9ityzmW0m7oS+BarPVOxfnqndcUUcuo/oBiOR9/DeTfXrz+ANoR700+cH4wsWig2N
UIP96tbdqbhDtLnJAN7xx67E8BcTjUHRbFC0u8Y42EpIpgy+Jfd3GVKeK8A9189zLLWhFZLNUcVq
yDfH8zKDZrzuGw0+J9tJqHNyf0F+0SsdlRDhkyYz//S92OYGZgfEX0hRgPZuUsuF+7uIrfdx1YDP
xPQFXLNLmCnQz4LCZdX0lwrtkG0iRn/AoWfoCnih843V9kbjAguUczmAuK3OynrggYt4sYwCfSe9
pXy3ZigApddXiTVJsO9GLzXLF6jpuqHoFcPtZuI5iVN3CROeLYXYM96vv/VgzcpUVIFnz1QTj57X
G//Q2YqpLzVxiXNG/6JfyWA61m0AZSE4Z5THo3iduVB/koMDvKh6qM5Main8qkZWjD9BVx3QgOIG
/c9bvQMGE4bQkW9bUj9xyTHAMKxiJ2js9DN3QxwAS/FT7cgHA93dtGyT041M6FZAMhaK6SMHf3LQ
srAMouDqMM6HvQEYBPqZtmyj8ysJPKae6o8NRuJz8Vsv6g1NjRueOMl6OTwnLfrlmZeeF4vZY57l
yx6yVGxJ2RPbiZ2cvEzY622vNPmRjsGfxm3d/87Mzp5KKUiO6BwJz2QbAzeXiK/+jdTdoffMnhIp
4/Fyyn6bAJYF4qOHI9z2+vLuMvmqZNpGbzb/hk0m04lkDjsEN+HCe98lL4ocwFaCbEfUXR0ka1Gu
pyN8p6YIoo+YgBU+m320XxpdwIqv43Tx3cprCTzdrqqZLQJjIYMEJqS92tuGOsiJQc01gNeDXQTU
nwxOlnsuA1hqzylSaWwuk5xuYvE9z09ACmEq4KRPkE1MenoiAHMxBLM64mzugpk3EOKgUb/9O0k6
ww8y3mTzMJ7djwI/V9daEFfep62XkGLI1Xech5l9Krsa6GN38GPsxyL3x80Z5vdW4j5+gMx4XO/Y
WAOBEXNPGzhn56YRrRmosBBG7X5rV7cxz1qa1nfJ5ac1HrYwYHUZNc5dFAET9NbHNJibDUQSt3yl
EXx9Pgfkix/DqB1ud5bEDFEhtR3nJ0tRZrKST0GlfEFSPMD8p6xwvD105RRHG7eRDnaDvrYPAcl6
cZXsz0TfvQDocM71LrW4eujjBXL08YSlk+X9HLU3VgA1/ltuczMYpTRhU/XWeYvLNh9DtRSxmSKE
mj43S2gr4apq28nw6467+BwFMNrqrs+HjIaceSOYUpD6tsMyxOpHk86dxK5RqH6ak4KT4E4fnQ2g
22yWuo/tsxEwY3ze4BgDRi1iFYiPyq9ZCV9VlbjKJSfuJkZ/vDy3D4CdsOFNrWzTYMwBwD+gXBWl
t0EGAGyDSpcrVkSt+Vn31XRFRNcAwyPhN77TOpy1EA9AzhD4s3f8IZVaInFQotX99+awUDlsxIVI
VOyRFfvsjlOM5rCwfyMX5UHLRJGaz8T8J4sRqp7Qfnbv35W5oeJnWPgYrr/AEQl2WXN+LANVydUV
v5o3K85AiaJoAayZI8wbTXK5qsQ11r+F739M/dPx0zx6njT5MmH/bVL+iTmTouwsFE2GSdj9Kdts
S95L+IWisd4jkrG0zBjvqEXloOnDlYv5pCQTlhyfD+Xr8uKyyrrQnXGtUsD7oP0yD86nmd8ch1B0
5yoWDfX4O6CVOPYanqfgQ3UgJ0gXCjD9//IPnmNgr+bk4rMC++c6D9D4AcIn0QQIjp+56oVPrOG6
W+AF6cuYdmrl6J/OjAQ/Bg5AaHHpP37+8u1GMJuu1jlM4DTOXJ/fmfsHgHacEueV2FXnGQrZr1WC
3s6wa2RHg09Id1YrQu8PrHZVMlO4BGl2hbVnYfzeDUcBHHLazPY0IjX1ql6o71D2Ht60dVYgrqdo
OiliWEvA01PvcPWD5KC2RY/QCDnPOqrckC+x/OxJh6EreexOiplmEaSbJZ+c8fJtV+kLDlwmVIfL
tBRyJ6YPtdjSZdKVtibYoErfcKL/jrT/MVeWdDdS4hFaEgfO4DnW2+i7pPPSbZIRsN402xJXwrjS
TqOAZH5SQPzRpmutb7+6wCzhXtZUGQ8nOvFzFcNlvE1JfMgd4+KdRiniNXOB5SnXtw8LfM+hnzb8
glLBbkBuZbtX4gYA16L6WR1YHnAP5X07EW7B6RwEvbd7EuEe14+JEh/2mzu9tfvrfYBlMibwSEuO
p39y5pB5O0XZvj0zb1hz2Z5VSoSU0GxWSMmuQ11qKiJMoX28DMwmKPwyL3wZJ8YRIYMO8ffoUyvo
IJWZkNEuDBtWQ7P9uLpNnhl6xyn2v4SlQSlJvAy3NZlXacq3CSL0DWTv7a529GjLt+8VYjwR0IXY
WFxTf26KVxroDrV9hlrmWdPlA+bfzWO+AIFka8hYMF5TkY/vql9t3LFCV5nglIouQg2apdnzSZhd
OIgUTUiC3a72mHuzFAPo12bUGARUttgk8SA+oeSk1bJcMy5f6kZRwYqJKwyMe2ZgzxpRtIPs4Cvi
GJJTyxSgIa+dkpOHnHQLcK5+hXT0HaM6hrcIItMbjzZX711G2NZITvvfetfvwii/cVoCKVJ5eo4b
KBIfmXClAowxWtVy5JI8OXY9ixyCEiI0gvDpq4u4YJ5dDON6xSVtW9bI8Op5Ds60euRd5YEPsqXv
uh1Iyz9eNTRmwH7SrkdHfEYIW4kENhUAuxtGqxR8Hgg4ZoSWfKzbFIby6ejsqK7kKXJj3QFJn7yl
BTian2ylQQBtINDHXrzdF8EPLpxJddfPpOWbGeZhFf0XMe5N4booeUjej+eIxwPFbyqt7UO3LbCe
siRL95Plnfb14u8yeQVBPQl1gHXzL7ZB7/cJa+aNhSXF7NGBQiAsjD4dzOMgVJKejz86utrzR9v2
2vYR5gCVIIpgPdurYBI4LPmCQvCpj/Hb/+6pxmWPiZityJg2h6qtfnmPQHUYn1mHLYmfA3Y+YLTr
es/9ITOy95NDTs2BQWdrsdjSn6abTw0lQb4Smdnve/xopmk0upfwFSZx+LpFehOKs7esWszRe+Nx
YeacKAUVmoakvLnSD21//yICmF1u4HAkXRMFCg83fGYUGHQ4NMDrmuYN3Y+pEaD1nkuX7dtzWAJo
R+LS6tzcdtKIDBl+ae5dn91OuuMyvIaYuT7SIylbY0vmIqs+I+91wY+UYLj0kI+1qhrZsSpMPcUQ
4pbWEfZXTXVKPAjQjH84Hc3Vui0cjvqQlX7zVrMSsr0aa8zcWcTP/ZbKe+LOr4P7jhjWG7IBRFkX
Dt8uijgFDV3y10obuFgqI8oPFH6cV5gDyQB+opMQxwrIOsJ2DKwR+ed54MQ8UcOzN79DzbVxss6h
80RZUdbbT5ko7p54Vr3dQPIwxUGOXTmCVnyRGfP4Q2VZ9HEyBsmwpL0XCPZpdjid00DJzkr6NYjm
hFOVZVi0GwYRRZ4IAjou56O3pkProrFegLM4awujSDX4yJRDYCHtLlaqpIKbpWre5Dv9lqX79qDc
nqluCuoT9o4jLEWrCiIqryPhu2n8CPRCD28xTlHVXUl53mBf1G7j4vNGRYh7LoN1fvejcsYTis/R
ViX9vo75fttHW0nzcyjQxa/xdOBu2A9hnJTjJKN6j/qhhUcgIfIqRCZh+cNV8/ckvorIW8rocJNr
XkWqodBxMJjdJu+l88++Jgiz6YuQ1LVIAgEr5PWxP3+0IaQhl5l+hy4LqfZI+Azmxrkd55ddk3lD
ONsZhpi0T5Jwu2rQSYRLN/4aSRz+J0wA3PnuPfAVMA22ESIsUEAaaRQkp1+89BwrgsR2l4esE3Bb
8ItQn7sCQ55xdUTiah36vYXVz5e9Deh2Cz6eZwXH5TPShrEbaVcJtFptcu7VdSQykmsWZpuYAaGQ
3bVQ+krN9OFv5vvgm+qI+6Fx7JYdPcR6LqYFiJUANylOLN5pzeVzfQElOZU9uVzEs/6rGHnpeUCH
/GD4Ezo09zVA3kJ6GtOjQtmPz2SVPYVSza81Fi/c+Ys6K7qdh3lAbESkPOlXtk2z3U7O7W3ZgQ25
BLiUieiq/B4hQEh0QpKAO/haQ3z2WuuT3t5cfVBzOg1hsVjcBYVro0wJR3xD3XSbzzbFdXlKENIl
qLgSrLmLTPmI9ma7LQK7vdWtKdkqJs/CFTYH8N8SI+yG2aAhgNHLMAr2AVI+f3Tecl6KnfS3DjB0
YPLxO9+F42fuDjn7Wmga8J5Ej0LvsfH1P27+fUrzfHSTEZft5KFbUeW8j1fYxl14NS3bmt0QsIe6
pjrofdTM4JtNvxLkDwQ7cjau4byCzxKBYz+dgzQQVzfFESBYzgqAM4dnEYZdKo02IuKLWQ1dQ1KH
m94PPN3Sauz61Vm8hhUgQSS+1PD9RLfUv20xq7yqWTKcp1mxgeH1SS28tBV1TWj7qKyTvMz+2hnr
SKhuN72GJHfz4L1AeUGtI33f2iQiaAEM/q0bxqLWsVE9onim1pAZaBsRT/M98Ru2rcQEJ7iETVRE
+BO5WQsBCqexDpeR5Dr/zjIhz8G1iYrLb+a9U7XWAHJiOegxAgcg9YsGJqPalTatBj/4M1vDFAYk
5iNfDvawWLx3PsZB3XuZXjdtViHMLV7g0tP/JT60vmUVR9IVMa5dnUgAo4ExPQ1OkMin5I3LOff6
A26M29fCcmBYocTdIZIDo6hVbI5mS9ahp/kjXcjDmL6wcX1nKcyhA33RgM+vSNYmONBwZ6bcAvxs
6TSyiWKFzvapH6/sBss+yslQEsEOygE0WZxtsKZs8DYcVqK58IY4qCNm4gRtaprqbDirDxQtawcp
IgMIlCGNMpbxxp7kNjl1YbfwLB43lXfLnPx9ONUC6ci6IWUpcxfRk6jqCyQiGmk5iL4zX2TUSybM
wXUsVUWiny7JJaGdLhuLp9FUvEnpaIdyRfUT68VSpJtDfWJcDnJFwkWbPtueb37CBU63okPek0R2
q1E8T4A4snYMezcXIdXDJQGa6tf1uj+z1DFRUn95SY/wx1/BCuOsGxt4K4vYb4nnz97eYBOU9WKi
lxkbIpTJkG9h6Pv4epKGxKJ5mgyu7k5XJqhhUx921INy5VsCTDWlYAzFeM3CDmvxopE4UBtNz7St
QSV1JQ3OGOspOWBTDZzss88KYrqHxfGBGt7J2vhvfA5TxPvqZwawTb90ddTVJHrRukJNj6rJX/hI
iw1DBRhKB77xNh5UK1tjRN4GbbWwwnzkeGsV83mdpfwKT4fZ8bWkqUVenHcRETcUxWNsYRrOoyCc
ma1cP8w2zMlSjuuvr0RUVmMvgvjohaCIQ0WIkFXLIcjGSeyNVxNxivr1vL/t5cuSvHMAC7bU8nmM
DbVcbr1lB8EEANAz3o64hTekJM3+VEncbYs5qaAM+boKN8JE1EhQNNwybO8DtH3FUBdpkuTtibDA
XlCIC+cIhupQQwR24jMSbc/bpT+prDSqkfRChLiVAlMeqaGG7RA71BEb103Z3BIl44pXT4Yn3cGQ
//vTAht0laT41cYnXiKuDkq8PU8XbV6ayU7K0ReS4KXwlDWA1T7clEcq4msHb987ciey9gFb7PzH
gz6OsUeUjNPr/sV0/hXWRYYj2Mw6qn8Ns+/Qs4d+Mz7cbORR+SGUKRE2H+hwiaYHhtbgUU37/25w
BtI8tjB4ZyJmMvG+Xy71XLwxy8gsPdD1RVdqVaPfZ22LhdH1UKCZUg0bPvxgxeFhjXHO51w3ZqvR
5kftkE500d0CwOQr1WRbkseMOq5QM3z34pojiZShGh5Jtur5Y0exdeCpcbV+ZsKaFkbiOYqCwhF+
+wHsHcY0/Ojo0j/T6sQzQt2NQORizeIUTsCM6Ld+YCEe+ETBlR2RSPAaLCJ/qXBJ9d5p1Zr2BT50
3iGMX8Be1nlhb+i3h5rd9ZrTolRFCvCEWZQUiqAs0YapOxYzc9LWohJQyYqt8Mh/3dwtDvjwyeSV
V/i9GEwrjaYLZzKhs6CX/rdAvPkhuA6Obd5HyU26KMvGpn5Dah/kU7hZrOcg2u5Y6mJB2tw3qj8K
Ceb5rrJOLIipRqh2NVLqP1t6AaZ74+7UeiiJ7o3GSsmKEZJRxIlyuH5jF8PZrvxYJFwG6M4LAaeL
FSn9+HIFiVCYyXBOf73b1Xn9wk9Aegva5vPo+n2GpWiTXTxgV4rYSN6A48bErzRjCJDICstz9C/x
ECJiwFKG8lA6E3fk+YoRx/zVgaJirhq7uI8kjej25FHBVaZpOc7j7JmzlI/YCO1lLHKvU3AN/87i
BsN9/bjsGMu12jLZ11FSD/R8QZHBFnuz0ldZ8Qfekjd9n6kv7CjgzEtCbjzitqdAYQ4DnL0c2YcY
8IEeCzpulK0KLgFj5T8lLH5Jl8abRmEYHxxp5+MnY9V8CZgSCwjgm8fujGCbkWxwoYJ/aJ8sX4MH
8jBvjb0icW+b7WcsAus1uWXmrKUwoW01CWFTZMV+8Y832MCO0jwJrHUK9DYL5lXkZosK+oboJpxh
0uBdNZEfBBcF71JicbGoUj/XjerWjJ+DL/gc8zSyP4ClLuOfhsb/NKp40c2GLEIVcx5dHlPXjlQf
7BS9Jv2uNkUJ51RiaAQacgE3BOg1BdvKgv6w/2zo0wrQkAeqT4vj2YgKCgMQAh2v//q1LZ5DqxGC
TnzxBDA0DDHzkCk2+Wm+74D+l+HXUbn4NJmvrEXZkcxqrz1BVhQlucanuJ7RWEcaV2vZsSAmPQH0
YfUXuZrfN9QvGk5CsR6pRezvyYbVSsn6cJaXNuKxeZFm7UslZ/3LCzvJt/u5BqfcGo2wDneRW2d7
sEw+6bzNdmrgmBhNorNGgbz+34trQJMVDvs2Mo1jh8jpXOFvNmOLSPw5CR/KPNPYsJl9dUy2Ep+R
b+rEb6OHIfWzAM2wCQu6/GgCoVg16Eqm+OfDBkrIpVKD5yCEgUxUXYHlY4T/9W8o9lngWunojd+L
PcKPN+X6d2A9XrFqBQGh+Le7VIs8sguAFhtwGqD4lNcQthGKklr4wj/jrbypQfNYqOkyYDu+3skS
3fv7mNAEUMmxqGdtqFrq5ijqpVFo7sFu8qE6oy+9h4LiEkkVYni1z7+SNNkcPouyNO9czwQIKbQk
YYB/K3+DAs4iTNvcHiwm6vzHlS6nfjjToDAr2fFLXL5L9Zi+jHsEUpm1ibc6aBa1wYJY5L1OBGxd
5uyRCNpFb76UG83eJi59OmdVpnNWlV5emQ10oHBhkN+n9AwpHOws/Qre4TwoUkE+5WczgFoY1gaX
x5slLmrUPGGa68gxxkWzlJlAip4RZVW3CvCxkZRTIaMEQrg1+aSFABZDFJvYM/dAxOoKvAkzgu6N
KS5bthX/wdWLK+HUJkRvpQOeEcKfLoAkuvVUy7PZFe4niPXjU0WQu8Aoz38fUGTDhDKC8mPdc0tt
MWBCxHVH/mQy0BIj8uj36il6Wl5Ll/Oqp0/KkCLN3ED2suVNWscS3WWDr5Y6j8A/ZZnV4EhlP6c8
XJRSUmabyiVm3ipt1/h/Lw0mC5QNLxO+29y59Wc4wk6fIlUYm4VtfEjIlmB2GHVr7/9Rf4TsO0qe
NZIxbcpS5GFFKHXicGeo4zu1jBT71zKvlcJmD41k/3PTbKte20MHW1s6C5hM53LyK0tvu099GkS/
1eb5Ij+bg43KRk35cafKtf3M/A7YABn8Ibee5OacmZ3B4zHktkTE96ft16Z6VBCeJdLbmSEr3ga3
1J1KAOBeLumJSu0hQVp9y45BPH2Zo7fHgFc4mYPJcc/ug9ZxWw6hysl2EVpGJngQM3kzZ+W+VGKU
IiHBNqP4UNa++aoB9jzxVA/CPeplzPqq+CtGWP2saXLaG8TvXQ5iZsHH9hHX8OixrSqW8VvjjAaj
5jwZ27Sg/lS8UhI7QTNaT2JZsaVdJk71stWqmr5qK7ZBf/kTfNOJrY19t4K0wFx5CTCBescjuOou
89S7skU4gA5WYazjw0OFR3834k6rJmgnabC7uLNfVI4VfGQjD1hNv1jEGnpCWbt7rr3ewc1r1EUy
lszDhl5iz5wJ2bUwJGSFpUwV1rXdZf5SI71EgNIsdLxyULLlAgwiNLbAgoOL02LYTQb67aaAdup9
duuicVTZtHS2FpPouyFUes8Pf4OItDi4iAOQSRYXg+Ra/aAyoINiULbYIurQZzvzklfynkbTVI4D
y8pVK966LvzMtVSK5s8skHjaAgSSspkn6OmXdpkObByETCEAj1oCLJ46GFFSGpCyC1MM7SyrsGLD
hnNczUVfqx+6z1zhF+pnEoI4OjRL41IVc9QQKFtncXVWF0R4poImPsuQjDCKBxx0+GupMMhBDltq
93mnWIg4GjxwH9uACGuMLJD+JjbBDj7dAVd0kZpLpVvroTl8+ZqgFIPKTeuBJRTK2W7mhxxnSN5w
zV/FvDTr/f0H6pvWGmSjcaZzE2mUUoxdJlv5ZHBi7ZAHyq4BkobR1o4uEKbLxZPX7Z6ZELNmVYT1
dCRa14GniSAxBRV7B7giBhEsOiu6FASC1bux39scRuBOVsrYvwGAaaHU7Rl/NeHaasx3HnIsV3OO
uoivjDO6NizV/nnxAmjERQR6Rff97+06bj78+ACq87P7jU5Npe6L/teDLzlHOVmpF+/6OzeROEGN
JIb+3dmnjTnx4HEuB2pemewECsQn9F3Ih3svfXYN1CjR7lHQ1qSLtn0oRtL3fq5bHn8E6Auh5bG6
nXVa0tsBEKWNarO/G3JIiZ0eDpI6j8j0cu9Fvoux+4hzFvJtr08qs75yvkqf2gXkcmbMswVu7a0Y
AA5IyEuSLPkfCpXRkj5gcAZasHkML36NB+X9eJw2c9MPL8Ka6SbHmTYV6I1BQRecqPUZnIPRW2nm
wSk6jsRQfUScxur+CT4Xuoguh6Cwuuat96+muCdpjHxYZD+Jmg7qT0NcJLocTzY7iPz8zDNr0tVI
+HFic1ImfH28Ue0yWyG++ZCW9Vx6Hzt4nNh1rUml40Jp+wBdJWXecU6IYlD5slEN7ttsJjK13ONQ
+jKpJ5KIlumunEgDBMJxQ0+mR26HVAkIkmEDS4V282UH6We/YVoOHPDJiYyiTWjHClTDb21/VPBq
NmVu+GQcpFkF9RGLZHIPs1x0ZH0loTHK0l0kNdjdTkbaChY28g2Z44gDESa0gbCfwX1YSObFoVW9
cwoKOMmIypUFIDrjiUpGebZggcT1T5dYS5tfXysvUbXa3W/IkmL3NZ9KemU8uUgkezOJnn61GaqI
7R+b57tmHFJ9uNFWJHCcNjTCXjkNi5mWc+fgWtZe7t4UjjcqmGYk72QzPztTWEXgfpt9/PikYnug
dOxSCkjWVcosXlBd2IFvrROoXUoINYepEb7ICTGTPMUAUukWmLuXfaTfxSszbGwD22mCS6tBMuNz
x8Yyb1i2RtqAxK1aBcgVR/IBw4TY0qlsFvrilEUV7hKorohZjJlctb5lbKla3Bf0wYYe2lNDxJlZ
eVwWxZMv7Te9UFYVqgxB2aIwR/UM1mAj4ED19d1OxYDuRi2ApjKjCGOgFDiAy6x805lXRLA7AhW2
wHHsGIyKyuIloJvjWyXyka0RTbB/sXGZqH0uHfAGx1XpnEwrtrCr0qsm8GHeUrQb+FcjgHE6+FDQ
E51xRzY5f6CPWo9os/aSYA3Qo2tGdTEsqsZUgAaz95Md6tprz4T1Pg5YQHOoPrq2+x8BUPwbrCT/
YjkgczFmCpQqfSQiGljPDnTKBthrRXC9j3eyGklrEXvJ/ugk/DLhU1R2rFGLh7huMhrwvUlsth+w
kZOtl+nyg9EOnT22SeYHUmyPAtR90pEhzuQwCDuWXbI4cwviFwPc148XNTFAuYzNbewnArQd6iWj
gRkxa+dRtqzceemp49H9Z3VgUJc3h2ZZnG9QnzzunQk9z0+FJc61YuPr6t8USNuJFYvk+Tr2Q/D3
GSo1HuUko2vi464EFg7Rk4SfM2Oz67EcMb9lr7+tCkyFCmltQmBqp3gyjc9O24pxxTtFkeh4G/8J
R/Hb9M1cahpcJ8YaYMhWFWJFSuOWPQkCoC0M/D5Bh4vicn3X+wIuIbCZ9XuBJUxOli86rq+2Ax8C
NJqoTOYZsZAECUmMTE8VrXAU2n7oKbawnn+NwCPh/9lkFb5RN50JqLtRKotQILw1RowAOMvQqWhL
x24GIJJc9crp6pWi96i/RLASCF16mbhdrxr42Zk6PeFnFCEx7ktgbduxSAcLv2gIfMJM6+IJJCmj
nOXSiQO44KunEvdkkNs/6cbyHQvjBiXxQyaa6TylbTJXm6k8rpeLROx5TgLGqxf2RX0HYm25p9os
neCxdEAOOMICv9rQSgJ/ucl8uinByBrOGXGRwn7rL5zMminiTfi8UcgTGSv7vAoJtTSYuJ+Pwm2g
1wQWuFCiMX39va6/bjcsMXxTrxYZEaW6UsZp4ZJXB21wS3n3AY3FBTCHQIGyCR/6yRY2OH4uqAXe
4ntE9ekYm0FL7wmXwkbL8m/k3LBWXbVSsHu0UmlYQgOUU8TAmgg6axSWyRDfTjlnGWWyEV+vUOus
nIHhWMLwPVjoBj/foQTphVx6GZtrnzeakiAlfJIcpwX8LEnb209B9N3Twsj5SPOZvpu1ucrwh4KA
fYKlw0pdu5lnmcps3ru48tUUotX/Hlj8FjpZHCsnC7OyW4UPReHnYgUyW6xLA4PxscZ9o4kInUAg
cZA8Fqx7+AQ+Rx/d2SkB0/CW5NTsgVwnfy+8FLQiTpgStZB1u2WIUfY/QB6+KcF/MMXBjDRl6HBp
7gXmi5N/CjRyRhm1fE8laD785D8c/e2OWOfcx4qJ1oii+9Ok6wJlOuuT7pbv1KTW6LAPBHhgc97p
swQjhUmyC+0yh45CYZJjAgSC8BVtPhkGFy8ci3DTtmB+QMc1Ym+T26+0TNaf5+8hWbBTKZZoyEbj
sWWo3Um7TgZwnIjOG8qdXyozN8xDs/9QoehIlLQRUXMNev5ht1XvUUsgXkz76vJNtk9eLn30sGu9
8myNkJCA97KJ61yiknGnQ9/Q+lStCA0xLX6S8TuKFDZkafAiMnMC+I0n3UsDSWVuTeSip+woj1cb
NKsBqcVmVv5TU5qGLemveziKX9owylSqi+4QZMZsGucnYn/74Sj5bk534qpbfTT2eboJwKo0+Z2w
yXfcDOyqnr6klajai+cSy+w0Uc8GL6LCK5W/YHVQydaf96oBey00T4mxmuG+tVlDYv+vcUsha2B7
G8nZEGXqC9tf5fvwq6UdIxSzT/xMAfvM+GB5WIrFUysLtXA9LNW600/afe2Bm7Ku5RSz5hXWpekr
35fqVP6EihyyfT4rtSovfHlXakMA+I+e+TsX0fChqcSVyVFLMoekWHNqn//22XfRg9KSaMxHtwc+
/SBax1MURw8tmS1pDgUD0vW+nW+/towetyh1dTWEuE/HxdMdO5Yq4gHYhRrp2UqQ+eTXUfxOQGnf
okoqZU/fgymQirPL+glvy3R8dxm9PpF30f+FpyNQ+byd1+tzBEOT5VHzmQzWPRHPiAvetgQdT3OB
MozFt+vPRDRpJ+oeIVwNbWduWE6uQleHn6+jWd1maK85RTaE+mVePVlUvqvbdw79mzAtfVTO6gki
pXhGOcQJCfTQf0qlhq1Y7LavAcFt091lAgRTCkQckrfSPFyg+tEGDxQ9zDIiNdX0wTb9D+MyzAxU
2l9MwMSwULKadl4Trb/JJa1vLYQdSiiymPHvWSkdtwZ2hloT/vXFu11nIaSiccWfuX8Z9baK6OQq
6ZVaKdGheW0EgOtu7nB4VnHJ4J+d3fXpITa6z1xFKJYOe8eUIBhILQg9TsMsMGur94a2pXFBq+Sy
2G1ojiO6lamoUhtyeJfdXhqt8RaorS0ok63uG0dI06IY++xaXVW7bXzqpjsz3JZF2tO96Xk6zQwk
y0+OMAynvoXjrMvPiEHPmocYP9NeN28GyWgaewLtVlpOSRFyH+0zWztxaj3ZgS8kMokIJg5OQHhd
rtxhxyOyergykxy9gvyf/bJMGOft4mImbUAo6+SGytTRFUKXItW+kH+eRZHsMx7wfrZbDpDUiNwB
VoES960RFq4X2Pi5s0EyIEtCtwUUKC9j8770JYuYJnqAbAO7eCIXKNtzqekaw2tE1v8HJMH6yN29
vOMPtOjThqJd4HDjOxOqjBqEvQ7/h1nFCqfCy87CMJHEeGBCnp0wT9uvC3cZexK7U+X+2p0tgAER
8w0kZhIJ4K0QUjb07Cy8ESY6JzQQDvpI6bSuNBM7lxTGc17ZMQshxye32vVYXEEfc7W6NIh+tGIr
B6WOBSEnzV/Lt3COELH2+ouqnkAd1PqWZUXJmI5pgmZGjdUy9lV3Up2ASIIA3iwBoQz05IxKtFKe
sHPIhrGwrnxItU+yyqt+Vs5/gyjkpHxT0CCw4DnOzfRvHX70qhY2nEOtT02e6BAKc02H06F3/P+7
aMwal0eYMhlrgJy3i5HpSc1nAGOxsaBexRXxMzTas404qVmkvyNlMOsi2ygWcGWeF8Xaju/DC8Bs
nnSh8NYMdg+VzUwtL6oyw/sUJ5AUPXdOI6gSljH6nl4y6YKc1IqLNsF4atP4/piS7TshycCEX7cy
TVTq5Ub8pcR7puFFLm1tfsiW+SIA6xyxFn6VDS8TzqqUbD/SDVx6UKcUcdaGNytgTvMG2i6671Mx
nfNzD1EfCaIrH7dSWttA3heI+Ru4WuuxMfF70zVriDypLXSYFaWdSl837wlpJpRep8YmSq23lewT
HxcFCyyUhL3NYYJMpTLLxScl8LkxHONHQgdp9W2Yf4HGEzgEsMuPICklv/Ey9hAR5UKcGPyZWWLC
/MT1sqMgJpjLzDld3bpIlwj1sWOYyhCpWTdNcmgKREBjMGp8VSR2/veNogyTuy+4Smfm28VaGZ7+
92cZ9HKmBUP2u+LAoeWuhyOYehe7lcZSE66OB36m4bwLwEX8Ne1mB5Jm/w2fNFPfp0QFUXYK0rpA
aIDUdb3YoPLWemJvKt+/xlYchmoSmaK0Flik8UL1lgqRLyY3MU75SFlU2kX/wO0ofTtMNBoc4XGx
fX8ICEh6qz56vWFYKEZwMTOISio9y9E3QaNsRgURug+5cevh59QcPcK2a+ydmhStyclUcXPgGRoC
+T0VwyZlwd7Gi19+ID6etNNZ1romA419RzRwHzX12It/YMen7zPUMqQL3j9AnDvLTBg6DWzE5fGJ
GiAtn4fDpx7ZIokDSkF8nY+B2DZDY3ydlouBkjWtMJFmMjP+MzN8AcqifqOFg7L0H0s597T/2Cu9
3SR9aIvp6RkHP+5JuEFI1u9gVN0Bdh9zEmcUvHcQeqNA1bJ1WyAmh9QhdfkdxQeieEn5ZNPNA3Pa
u3oKQ+v+2Og18KTxaydrQDyFb0arN7Hr5o4GXtMdAHULGa63iRKXhnRprSBhVC1zvWh6n6EA9uMf
meVqq9exI+uuhZvxAao1qK45C90jd93wfJoFpVtSiU7/F/9WzhGmH+micD3Ta2n/ifiN/wl/tnFD
B7NmhSzouuW3mwDx0rjActpZgTtRzIjq+kcXJl3paKryjM3LZKGqjko8bCFvMMLoVpr8wMboT9/K
jpeZU9ojcJSsdKfkh/yhet5b7m6+miXe3Q100tEXzV4NnmYu6ihekfXl1usKz1DlSqSh7MCXMoXf
HgjgvDvQZZOPJnxcA88vN25nRcvNjqBH4lam3vN/F9t9zPV7xPDttMEFWKG2CZyUgqIUXmCosVgh
/502KIqN4KrH/HlFV2mNRBeLxrTvdB6GSP6eXFRdopaE8I6VK0BQ/fNs1/uNsLf5fJ4tBDq28VqS
c3XczYpr5gVEVvl/2D0uP3gRIwSbp8JnMUbf951fQJ6V/ephj+uKfaFXV+AWlvflv1SZjlq7lQ7F
a1aaXv9FRJOG25yOO2BeGPrP17IA3pHv3bGMMLBKau37Jp6KSJNkjXRDotWP7fG1b/JkOu9yS+4/
3eRkDf6ybyVJqzK/JzyER8Pt85k3NanIm9esj0VEJb+FBNFFG16xBiVtWsn9eM0zh1cBjPuLVftu
J1/LMKr3LwWL3NkkjHeVUgp5iqpE1ooEQ1vilkLfDECEOdt9WfHF2Kna168f7oIbEXsE9r6ET149
a3kaJJPLMiRsRQND8yj1KxKKpjW9vG8zkUgz/UrNXkPUDfU9xKaI/+mKYkUrQg0fV4l4LS0f16t4
yycL3hE2lASCIZOGECuKaJGgsCwFEAkobl9woYWY+OWRps1PGma74cHDRXbusWymFpu8i8GC9f+E
igcCX7+5asYybEZ15dlusWF7t9kdkOF9i/Is9MfNrqqfGMl3soGkOHjO+GZmv280K9eA3tVSoc/e
s+weVP4iVC9OQojfA4Ib1rsUyMAT5vHfGljWfCtQxmRJ3A+0G464iEnxEZzwOw8tL+S7n633yEPI
rsablyq8RDNLuHjVzcO4wzvIsAXZ4cnE+CZUxcfpAbeesHwrBhLQU9MvpZhFUB9rljw9CNwldU1D
2bberM1QrrHOgdlHo4AkzcOh7L70/GnjJD6zIAKP4UPbxXAHYqAfKWkf49rbkp7DmV4NW5QZ+ofO
F6yz7o1I5pWUqnRRpcf2dfxdRus4jriWthWj+U/LFOK38V4q5IHItQFJBOup18ojChoolgizenMu
N4/b8/K/4oIZ8R1KQbjDLEN3RWHWBJ4vO1gCB2IWEKYZOk/DARFeBdRaQFFFHCbZqQO1JbzUXVWP
yXzL2189kHCB4fgGcq4mB4MMNRfG8tO3OqMY1h+BZjKBtiJ21YzziUUItFhmhdZn7n7KUoJMhroQ
gpSIkZPdfShT2tHm3QhOH/KgsDW74+fQwjgeHeYbHJtpGGz0iLvM6dlbUFMr06cShEIviPlWin8R
Q22FCyKejtLEw1QR5f1SQcW7h8I//YCXkvL7UfaKBjTPDeA8Gfs/tFFQQV6ijNb6eKsqoShBWFs6
NekFy07rVjTxXZVVic+AsrNycl/U40/bn+rDR8Z7cmNAsJwQy7vhPZoX9xhjM0WhcORFyaRusbex
9l01mpciJCBY4hAwAqS4hN0MBCMORc2+0Vc3rL4BcyVieJ6qoS6DAuoWp8+v3ExhFKAovtLTcr2d
CCwy4Hy8RA5qkly8lEBk365Gn+BJJ5xG+Q4nxyxuyNWkGUdtEdjJvttGDVY9aupaOJC5zVXWC/j1
KPuo8wsgYAgaFDnsOMrBB/DrYaFVqvNbPBexUW1t1izuHZXZr4ICnuoE5YujNrlN+mBBpQBglI6J
kTlKw0bT9O6rIEsoqbnenXsrNLltiQupOdgNSYGxRlcjWJu8D7B5Rom95aAiK0DVGsdQAI8Xwvis
l9NKnrUJeWQ5wE89b2ZZcXpyvB7BhkKnCOv2+LYuLLms8RLUrtPoQA4D84wZSdNmd9PlgDrVw5k/
CyBOCtnUddKcGs8R8kmLa8BKCjsmqt/l3J77XMkvcJFUosoUPK7QwsGzht+wDZtkR6U3BkJqS2td
Hr06ALKzrzfeoH2cekdZoeERqrQLGbQDvyTsAdIaU1eWKFv8UcTrhJRn+8O3EangaCYWn0/ZHfqJ
JmY9o3UZ0xjH5Iz9+OKlkqambbCwtuEqiSERakmDRest1TcGlbMwO6SgtNKvA03Xqigov2bw7NQe
RDcMR9VIc/D/YcAt557nabOy1NroUatPH5oRe7ohhcY0TjQgOmK+ydIO3nFXzuuGtAksJILxDouU
eknULsKT/oodMKwl/wLDOVekFYHDK1mtWt4dj68WiN1BfUkyxWiwOYPVFPWIoRSkiUtlQwZKQNmi
CI/KW8fssWfTfpL/YSKyVAkslXMM5MW62ZBlh2RrFwJnDHB/ahVU3eEhNVpl4vcwpCoqLCOwQu/1
GM2JMBHSrX6PwTCU2m59ndOsOIRBxehUOszcJiKA8pIQIaXyRrT85TrqaPJcKOezfvQncDwXnFcL
REf/pu4sepZgyp19THD/jCf3xmu3ebEUN1saGon8T244RyHZ8NE0WQdSkteGW0PJkWprJoiE3nDF
uTiurld0cvRtVOpUOXQ0q264F4vWAx+zOB8rNYGBwU81dves1xHwp5kOBB88//+FRM0Wa87qnyB9
2JqFSDPCWgh/dZkK1QO9AKceJCFgYrH8/cN+xdVa9bQ0/mW0mq0za8Fmn3iGlT1mPnFTg0QiTM1b
D2qTC8tqHWYwkU0lpEhJFdie2IJz2yct0lFyGtKAgzIwI0eednwJAva2oMAxvXnLsbOZwA1bNJJV
53IU6cd+WJQsihy1lLKyLrRFZc25iQCc9Ke85r4VgxpYYYq/DpAXmCrugFZ33rZWoHTG4Bvq2Wo8
ru/ok5xJPZe1Wnyc3fU7/IXXIaaUcBDGryOLdAbf1nT8H0j6cbN+EuSaRRieRWIAiaPNSzu+4EHq
6jYsC2CvuV6Yku3dCHm7oMjIkag3iBtrA3OcnKWwt9pVJM7WSNkp3qhTk9LM/uDWz5s1MCqy/K7d
FQia936RxFhVSWRDXbfYEALG4APSAWrDFS1kQQC14U5EnjD+ODWjn6LPBt9mNi2VCeXNjzb0AqZd
CUY2iYUsKNnIcFnxEn+wBDWYacw5Xh82iox11PYFTVCjl0EBuKZYSXSiDfCeGiBA5L2haf6I5xpU
dkPw6vqFt7N0j53FYB/t55ZnIN3nHUPKn3Im8/9msuvplyRMbCt7OGsMJHI7nXZVe6EJRPw0wKFo
Yg4bL8mBmDCvzXdMRqLgBkCI6A0n0vjHEFI9dypfyYUEzAKaWQ0ZGxtvTaeFfFpsgb+Q+KPvrgpH
g/gqTdkOshUv7osOV+74xnVYHEpYgruqg0eHeK08DowwEFW5r22GnWjFYCecX+w+gKtalQjf8vPC
q9tJVoptGARg6ojraHeicyck+uyl+fvpyrDc60GKuj1/6N9iDq0+pqYbQ+W5fPYh7TtZVMQEiwQ5
THsAfbGyAwROJu85bjY4BqLUFOasCNPeZKJPosef8SrCBlTBf3v5h2YtiBC49fvdpQX8lmOfSdhi
h+VBQ4/6h/VACl5qXD0lAMNbE/wvB9Ag67raMba2wytNtbIyj7Du9lnSRmTLTYDNqL0AEkJjZ6QW
m+7/eqERyjbKuTV0LkU5SDzvPsHUR7cZ8wOMeZy7fHUoF+5JXcN9Rweq/Rx6fkqcnQ86UuEd7rwG
GFajc3CsJLn4jxJkAjHpd/qIlwiIwYxlm74ng0ArRnJkxX1txxKQlAIIW8O+QgKlVoZKjQhb3j6I
rmIYK5gsv2YnNUKWVbNKphD6+vgxjLJjsx/2c1wc4cb7NvaXWxBibG7PwDWr7c3/7fL8h9A9vFzu
nVPiH88F/XbfRhJVumEJnZj1tRFODNsg5dWUAIuQw4JVdUealvV/XsNGceMzz4LmYr5VkQxKwV93
UBThoQQb3/yxZefqWU5y+qG1V5tkUulU5CVIwGoDZY7+mlWJBCuHgW+0iEoPwPTsJDWFocrs3RhI
qG7eq09oBYADOdOYPjV/lGzUCu9HDP9f/KgdrMAKjTs9LnacaS+dZA1bS5JM48BRLVmpABeJY2Zu
+WOpokNI6wRxs/MH9xo6OP1g9ARkdABO06pwVEDc53fH1NkpsHbkeIClQzjRby3HLMknr8M2QlHy
gRf6LgqGeioUMUAvVSdqsXZcUWHNJgBJYYKqjA+U00uj7kYtv9Q4xD2eMN/Kr/O81LpCVcY9pj8J
Uzh2zUuAdXd9OupmzOjloURnTJ1ERJeYIzPDCIGIECRO+EqS+2f2/+GODLeY/CYc8zfdhbVIx6Pw
RpvKHFBlGDARYay+g2O9XO6njaD1dWqZS18uyWn4gu/64HVFzIHemWk+jKl7mBlwRMywHG4zugtV
3Cu4B0hkhQHEbM89Mcz7OUMwLpX4tNjUGWcdWYaNkRU7uGuWCPbo5MOygwcbsf3Who05PDKJzAI8
JTUpsGYW2mdEjxctzsZDHTb3ADK6B0LN4zybDUpIgHVgUQTWQHlzgjWHtTv24eIqmRn3/NOETrSH
p8BBd6jYP1wUtGu8Ed6oaClh9Vqr+DC7L2/62Iqa+hR80wbb9GpomuXzEsrE+wI9l1mCmfShdmfA
paYIQQcQpHF+dg06K04ARGMCJgB52p7fi0IvMWL/BDVEaIlp3jiNjjjp4AVrlmM/ILHCXLhzEBPe
d+P8bIUxFk4e3q4mkXZGd0aowm4+sDWATjcGslWUVgNtD3JLc3C37y9gXokgwHkIGlukHWX10Fe3
vvEEEOHKx9s8/5OyU4z9i8jYyp9fNsynobGUNRFWkm4YzkXieBuiT/uPlFVOk6VZUI94e2bP4Ezm
eWkuFGmeya8CUnE1vgftWRMGQbDpcau2hQAqqaq4Pkmvn1fliunfcubGhnwh8ILaGkHfDNV7ymIM
l5nDfQgFqF/lDgOcVBJonRYrzzqGJBnzMU2A+abkfVBo+5/lkm6Ug7BoK0e7QZK1R3wHdio+nLwb
GK7BGG9X8gZ3lRuRu/gkDG4aPq+FW1A4uyEFJ0o5UIKfU1jATzkvxH9c/7DxPaEJfYfY0TKLvd+K
+vG4R9iWzzb6L4P1Mvik1PPztxBfj5i2202B3MVwixoBDDB/hkGIXXR+alHoBbu41sC5uWYQf4gx
+KKCtXCtq4A8fGbiQ7ILoLDEaIt1owNO571Tv/hngvmQJklWgTKPO0mndmjgLbmEYDVJ1EwloVN1
UkZQs2/R9gaImpYOh2EFwLU00LA+1oiu9WYG4E3Esj6LNbGPC2xVsiCaOO+2RFv1//LqoHvrkpoV
WAdKHk49Zyff1ehMM4qPtoO/Fip/8K2PAKpLAbh9IRl6V9Coj7v7AVxrfn6JpYcdN9lYBETL2fEX
08l9teRFTIJwnTU3/8vVTjdcMoglZW7zacKUuSTbSH3GVTD/LuB14ngFxmJHYYuzxs5XzcqVXd19
UKjZiIStqrvAse4jtnRKo/GnGvsStMHIST/us/8p+LHYxoXNKJR6m9gX91vxpf4SKZmZblc9l1Rx
wix6EqC4wZdQawcPPpz5wc1SUkvbXGaW54amzYQuAF/HPQVqR5rhMJrvxD8XpVqFQjgQmA/ACQiZ
PKLf2EMllY7TyYcbDIaa6F/8vYsinhSIJ8UxfdOH0YKPrbqX1D8qyFQn2rbgJdRsAA00zZjChkRZ
RkTb81Me9N8K6QwBldM43omdaMrg5VM/NB/YUg4w8ciyJJAe/SFanU3G4Pm1bkM8SfpbqP3vKJYP
ORTP9UE7CVtoVjOvOHGXMl5M7ZOMU0I1/qjx68b6XtSEkbDwLQ68BKFjytGaa8wOlBolf+ihZggi
hDCUg9QElriucrEXRF+6Y58OPjxrk7K+fN/Z9hm0X4kOD6Dk1TlT27vTp6M/tdPfzQesLm8tX4NW
ee+IEAyicg+Q0jaTFO8B3zV8EDOfZqMpBiirgnM459hJ39IsCS+51gMeJGC+F9n/UCLvnS5KjRlL
sga7N8ZPxKQHMmNba/01zd1X+X9bDMg+gwWhZGo/7fPkNmGN30gzEo6pJK40c1wHhoQvpqPdiWxC
hf4DosxuQRitCvR7YnkMabKFwXsbsSBW/XdbcTYmHjfYwcHw7+45xLO9HQbpEqJ6DzE+VRihtZC0
qfRwZiwAV1LHGaLOZJz4bq0KLN/868cy7gooBooZJRVJjMW7Un5nEQmkWuxVLd9UyWT9W+K4QkOf
ZyNKBG7Lf45Yw1lOqit/DEPpWjjQ+d8PyEVVrw1FQGN3DTHz5fbINXrzz6NIGxIqp31Q/foPVqQP
lQxkYaw3KKtrWHXMBQ16zxO2WdatIUO672l0X2+hHj7eH/89bJyWHbUIKRM/YB+EhmJmeVSh+0VP
8dBzPbg978mr6FUqkKf0UuvpYsX0V17OhOFwGMFJzgoye91E3Rwc9rW88eR6Wqvf4uPvKkDk5OSs
WBMeWB2O2PjQDH8AIOXWV0nfsRabJZToLXuA7eBN5w4dR1BGp+u4MsdpCaLEk2xUq2lBtaEtcdS9
mwUGo1OGwL7YBxI2uA34fvn/Uz3+HypN+XgaV6YvC30D9qGrThKz+ZQmRrve9tZeaOXT0YsA53kX
uM9iNhyp1cWzSt5aAK4M8Q5T4bD77WDWcbZZ6JhfDlQOT4WddAzrZ20BaUMagkfLa8Bv9TksSkhG
p+D0Ngiewqfc5Af/QmhMD+oI8JAAyS0UTAD/hHZLiqEwWVm0zdGY2AtaVYjtkx0jibWs7YJiD0vV
C1GNqG3tLn/sWsiFJUAWIJ2gnEMcXgi3vTIGfZFCPGlMbCfj6y2+gUEXPjfvpbrUN/s4LCI/r93I
BpSRTmqKGvfwJZR7ynYqctiocMHDK5z+TndRuJbln8EJnX3Bq40Ik4XGaderoMBdK8D3+ujdAlAh
i83D4qZ4AYmQbikuYR9cZqUcFgy4p/c6ifmLzan2uGmItztVPnCicbsEzLtXv94j3PVDm6CXU8uC
Buq4qUrn6YO/lbIdFqCTKx5HLxTUbtK8fcvplj1+yRr6hpWa+LM7PVVcT8itAGtUiT8aObxoDE6L
zpiSuY95VZFivz35Ll5uUMLBggTqbkvC7Ttxm9QTdMCqMaocfadyg186WUPxWNPBMmebaaDm7QSu
XpeFIQT3Ho/gPhq28Wvn3P/1dMmWnK1Uir8GXXPL6gmpCzZgC4z9bpvXhDo3egvSr2galX29GQoY
yduQso8EptCZ3lK9NBdT7q7C3lqrj6rNQJCYqJkp2T0dvcp9e5NV7rxoEpfdEZVF/Z3yK/S2GXCX
1kiU0lWry292F3CTjxfAoQ26yA+VOgU+8iXacCshkXNlKojz8h99m7wBPRvIaWL2jMOKWMLLvEHH
9z9HXh3quYegqTksYietlAd5zbcclMAJEYy8b+Up7Xe2ZBKj/HSROH6XSfumIwOylSPkU7f/L0ut
R6LjnK89vUZ9q4YhO0FlHqPLt8/JsL6VOKjeeOSDmyQPKQpgxXBOKtg+1Qdk2v3eQJPhIUaFdrqX
qmN7jwTgvNTtEjSLXkvIYZtKqjHvKyFqS4+a3fw2mRxAz7tkiBxqTjexa9YZfikVyFtg1PdIOek0
5JW2UJVKH6VCrQwU9Ge6Z0Tx6QiLvGNlqWMR0yOKEhfGCPHza9TnCInDk1eVYzXTP4Z7OPwWlHiP
9BUrQcRXY/aVcqBeFWNZdUhWDesLW0ocUK/iO1J7tOJl1ZzVo0Tg0DM3tAdfiE0AW69wmpYixi2/
pA6wBvvZo3Q2R6iBHrAH0eZGoDnLvBlAH7z0oqg7/muxx3dw2oQDwZXleA97tlRTl+FtNYg6iMjz
FDrPZPIK/wMdA4hXTgMKbuqCmB7eZXIgxdCMbA828lZTPt9AiA6i3QEtJQc+1/Yz+zIjrwlRTKMv
lz5FYcvekMSqXonA331/pCQWIf9I+JaLBmFxjOilGBI/uzYhftaCH3EkB5JoMLbSXI6N8wG7Hamy
5i3ixp9zZLmShAUEenc8p5YXNwfVTjmmJeI2AcGYDDBPP1HQau0yh61FxxUf1IB9beBQ3665YuUv
+VHkh7uL3Fvp90UiK+NoOfRDAwMGEZesnUtP9h6KKexWXQvjhND5tLXObi41YgMtrr70/Yn75Llb
lGzcRycnoEOzEA9IeYRVdbO3MbpbAZKGcSvIH7QE9HwkMDrRr5Mcy/RpfrHA2udmGtwKE62t3rY5
LIk8kgTDqtOyYvB2/2OB4EGEaymS1UDdkjDV0KyvHd9RTq9eETOKRPWCA7JmOICJA+DYaDIuz02+
X/5Tl2bsNb5hbvSVJw4J3V6BtVDBK3MxX8GZuP9ZuvFp4huJX0wbpMQKQpDKZAqiq58Gpl3kxTwZ
SWY3o7thpfHwdLG2SqKUrKdXxoTDKfhmxHMYOlZe8xo5JWSgL4lgzN9lX5HNIQG8hDPazOgKRN2E
FeFNjbx4GNFEFsi29H0qwJO5c665CPCmDXtxZ60E69Qz4GlgPLjJWI/hXeGu4HGVQA1a0oByM1xJ
zEvN6MHOsuH0BTFd6/M2iZtrVaHqIX2Bhv6/728X1M4XlXWJdYLKNWRAaloRPZdcMJs6qeXPNSEk
t4XZ6RqY2N8H/cI7W4rLwh6CMepezsO0kvZ0DqjxYzLyIsjT9mPeve1sjEhHtAWe6/QXS/2SnTS1
7dTNAeXbEvedpzMfTnmiJfCdZT3S1f9Swcbfb7ROgLFKC1D6bFtqzahcFDpq7xglYF/5vV+gyNH2
7AZWZbIJbhNzrH0bkfCc4TFiwNWKW+qxSmWSwjh7rKZ4yP3LB2T7Jys2FTE76/jkd1FhnBDyvea2
sfrTbqYEW1qBM+HKXMVt7ZKNqY+TQ2NzAM0OTgm9spmeh7oFsdmhUJQyTe3TfS/T0A1LbQc0r+Vr
dlIbwbTPBkYPasuXGifGf8s3NPnezKb9xihtTVl+5TzpdbmOFK3XAvu1RYqSLadPF2gaifsskHke
JbD45+MX22FN9vdj4QsqAm4SWtPky8Qwb/GGCsBJZzcddpoMqIKI1gHfK4+XRZIFaGlfGVpjHI6Y
KEFmFsEoFzBF+YaCCiCvg4OkJM3CwNpGT0MWMJUxhE/CKx13L4n32JIZVSiitq2o4qyLkCz9lfr+
hTlHHtBiP+H/guU7GyDUC/OV0GQ7+mk3vHLUcDkx8TxH0y6JbqzpVvAMiok81XCYEBZRpprxG5Cd
fB5cx8898ibwgxEvAiSGV4uyJ2FtDxMBKXT0DcLaXl0ggmUq2C0wvymm7lnrlbfk41TjHbVAxL03
m9PBoVJCAUIFICy8F7xvLjod8kes/JRLpND7H05xLkd8mY5lXCC3o6rIYV+u8ePs0eJjpKOW+iu7
bAzzz+NwLCi8YEJQSj7kDjUxBSExccQcyJz9p8QegNWQQsvQxuA2PO11rkb0CDhbP7vSb0kuiFaX
++GOL9Zn1Iijx1kH+I9BKg47nHBQt0FkSqeUzqVAqTtgero1k2yqojfCqxjbdFZrcR5fH9oPfjpJ
HYInrosTPq4f/msal5sCF5qz+qiOMr5PO3qdhATKqipD6yb2zGpxom7GdGnk0D757m0+/UN+Nng8
E1nETn1c3Q/6piA2M3Lz09v87rEbtmcYHU4TxbAlL3SQCPk48UNHKOcB4hS05Wiq9jMtH8iMTo61
TRQSCyVuH/RoPAvM2vMXCsCmbvvf/e3e4ldQpQ09osdcr7ejUtftWHdjHLSvss8dcavWMMu/3SUE
t89cg9Tzgl/KHHFLoXIyzY20ZPZhqjOJaanHbWAkQgTPiHR5nEnSB1cUCc7RW7DQyAfSgcKvQjzH
SEqTMQR2Thv4w+vI6qs1HCOa7BWZwFcQUhqwlW0bLmmS57nvocOMGz22ch5pImLkVk4NmZEOw0Cn
FOKEg/ijYcrqa+luG3qbb47T0yay57giDL7JjIzVW1Nrbhv7Tzwl6txVlRnB/lqye4yn/fDlk+7l
72jhjuwNCUNtB46/MyWCRBfD7UvKiEdY2+YtPWCesRwBYaWkSMTWHbqUd/nr3v3GJ5IQpZ101Bkn
CIfLQGZtLqJ+ZmSqo8KSF0IO+gKmE/3vfeG3gLhgMkdc4I+HXnX5vhWT/JTgY8y8V/WYM3Dfcnac
1qrpiPpTas7QNOe3K++PU7beyXLwRB2eH+rRm24hKDOvRXovfju3VEbA8cuj0+j60/tQEUWYWhjp
hJg2Qd2eZZxasSbtMRMqnWV4Xj+SwWGD2+/SMdnQeFP1df4oG/i95AhQq4FEYrEEE6Nc8vmpzRCG
Tv4UrjfnM21gP1JzAq0HFB165OkFcUTo7vwDiBnEzn+AsqAPhragpfG394Qqlcle+YGlcYxgn62b
Kpz2wZ/cVc7NLGP8tuGkzmIREIfnwsxxupiTekUrTNxrVj3Gn6DzJUA6I0ZIuWspk4xLGWXUYtfg
NuTB5AUq9y8HaH5a0I/gjflgzTC3o/tfct+7OwAn7e6vizEOdu/oPvUo7ef5HZsv4xnUI3qhwHAY
6vLrJOpVd57CGGCxVQ44DAczehkw706naxZF1wD4kGibzn7+O3rnILev757g/2KW05Sl+y9uTkPP
2XDzblq40gox+xgQT5pGgXMhogDZc0AIK2zMVEE0NPRJNZvf+VlHYq4u1iWiF6XZjhYO+U1DDCU5
nO36X/Mnrqiw8/NpG17GMSXDwLm/f3u0KEwIc2vu6SW4OSd8B46UrVPWuk1q2AKiXEGjxToUfI3s
lYmx8TCL2n7gb4INCLXIvn7DoCHp5QX7Mf4sLHoby3x+5Ckdaylei1WGvuqaXDT++JxhfjxJzyf+
JfNhVqZ1KXH2+epKwiK78ZwNpTT7gECow+LEHh0/pj5nZOOiMJWLdc2cjky64ltwzh+2Bgn/6n8Y
v2NsDtIUPjCI0q7OmJFwYnIZwYTzLKzHlEj22qysmZ4KAIKizr61O5obBJ+2ENHpSbINB+4so11T
xNCPNsyjNIo83062xTtO86ta/QwcwFf2D3UxeIw7joIofyqTQ+RB2UJOF1A0ezSvvw6oKrLhIv/g
l9Yp8Fl1meZSW8XkMuxLig6SEM7MqvMl4u2f2aUl4cG59rtFLtK9BYgGsVtyCVWAGIdAhR5uwYqk
1W61QfbpGijeN7LpP7gKxumgAdvxRif+F7XIxpRZqr7+Tv5Ha6rxz3p1+3GVxF3OWNOKQ92ujZ95
Soy5Mo9l+NkPyXK0hRB46dPCjSXeLZZkq8HzwlJ/wJz9j/NT2o6DRMf8WyTUYmlKYuc/no6iUu3D
y3XXpHyVLSGBs5CLD2ABJ4nKt/7vz1G1Bkb2zpmD9KMueYHoqr/K0DVzIdfc5bEqtlfyPELx2I5G
gemwTzN9E0wTzP/IlOSPVdYNn1Q1e8vuKlA+vAN7eG0xB/u1dg5CEESlZNpTbES/9Mdu1t4UxV5s
tR424DN9JZwBFO690bM445ZqMozMaZWA2IRNWel0RUFZyBQJ98FA9bJH3MZyjvTabSPlHoIgoiHF
3iUym1H4CadO3HDgYc3rEYzYFYVmBMl6ZuO4reUzTViOCLbbjPjuIyLMpYmL1lfedXA8Ji2askyq
5nHGe6DzsiyufLzCHpEWNBwIBRiGiz0yw5Z3dXFi/GDAi4+kw/1U6KWCzxhL8P6wj4QX+/zf3Bqe
aIDpLf754K9c/vS6LgVruMTuBsTYCflXqB7BmQzNEwVPy/NFbLEKOCBZP/HpqhhbcSZ7wJM5McR1
EVF0TqpEQgMoK9PVRmqEMp3TtIcrDuC8xeRohk/k3LqkxrmdmBW7xvfcMQ3uu8JPOTOxDK2bqShc
dBeSKH60+VFghbq4aJThyrN4EsBzTisCkkxPv9KHoXafLR1vzFBN+hImdFlHfniGOoKVuIqKnP/z
ZzH925kSNw+wNi9OWol7TOetEHNjKUgo963kXulfqlTmDCX76Bg/Q5I+kWV9RXWUu57k4HIgrBPh
KMWSCQkVc12OwyssHcMIUrJ41iRzI/8H4thREyqevkI645gA4xdfj8pPdgBVkRsz1IbwbDMe0REB
YBajKJV+/cXcYpvK8sOpSkl8BTotZtK2RVI89T+hf4SskFtjyIVjKFff6FqNMHVg4MZ5mN/TB1it
Xg0/YAPcq3Cz8p8/yAptH8d/4qu7XH1K3ThWMfRFgYpcCz9UiNecSIoAY1FxScyREoC96Eqafwso
SX36AyncIeVugmLPiNV4tAWe9gtP3ToRG+mrwVIyJX6QlkCbta35nfKpJmHqXrD+zRN5vGQYCIzt
vUz2eDGjbpclDu9k7A7x5DQDpI7RmppRec0njk++Sc2C5ojCEJIVnQqsicBTBvTpocoVUwkMGChW
4ZJTjdJXYoKZrwV4gySb2LhQuLzpqdGzGuD/dNGBkaWqFJ+ng0kQhwJoqdrRRFo3vNEJJRmwknJX
qVgp6WJbpKuKAxYXHCAq87Pr1we8CdT5SNR6J2VhxFPu/oFbM1NrUUyb2xRah3gSNthmo+irIj3c
/WbxFXFFqiInynA1wg8bClntX/fbVBEDcZ2H3s75Cc3XLrBvP1vCsuBD/8NzpkjuxJL+qfam0W11
QQFHzUb78IkRNOB1RjcpOjjfexRUSYkctnprzau7vAZ88ZKp0cSFStAjBBXCZxMqBcba/bwAKjxE
0VBb6CgG8TLWI7ZfuvIASVZNTLp195eHUJ85EIbYFtJ6HtDp/mOFqhc1A0pWjW4If09kgYcCrP0s
LphMQUF44wvwjd88B54oEcyWgwfQemeZyvJBoig0TW2VGTEY6Jm2lGeLF+eHRJwkXBe1Xwoc3BOb
u7EXb1sOiTtgZJEHw1sIU01ObImlELOzDFfftASJMJoYQODtvxtwNCHdYmscWewOcKfoHJna8gwe
KJ6XByX39L6wRThaE+e4qxmBw4AZmc2Gc7PJAtSKT0QP22ga1CXurqGvjMxJ8HsJD8UDmx4YlKlG
iLg52095vnZit7CLCI2peNJgen+WVPId2j3KQY8Z+h3787yMgGUNlEEFHFH6do4AZFhjI8dRRVLY
YgltgXzGJ2pxZxaPbWdA1HT6ifWDNcoCqumPEuAwcgLslFRM8EHMmhig0s2CqdeGEWO5013aOOku
Ig3DC0irHx74CLUysSRxF9TnVbtZ256/lSbx4J8u4AwqoqCtmnsGsL9oO4kfn6YEwKPAQl6uqriA
TOD8oO2eubu65VuIxzVIjlwsUXg5ST7lu4pwOU2JbV12ImEorQTQnGR9XBpozJ1DeQ5A6p4PTQ+P
nk6qNWLYj5az1TieNuc6O7SsHdKlmWXLN2exZSJwiZgHZ/TKPe57i4Alsz0W/Qc8sVuuJ4ZhpWcA
gDpwzBekvOYGsNedLoYosqd18yLQ9Myv3kr0Vk18oLa+lmAwVUPzjCq+PLQTZTZVLZm6cSoHTgbR
F3IzbDRQLp5Ny9EzSYEoAat0Hutl+Hrjc/Ig/XdEWYh2pDP+M3Ie11HgWxx7zZo5xNvlmnezTXOi
FNMfGF3KEykYO3j1AhU31wLAPHr++5orCqqbQXbFgIBVhZJ7ns4RwcFZgK9MQUPsVN0TxKTbl93B
thlxKrqimQTRVGZ6pLFaEX6htBfA89y2LwZkRqESBUMMqVtdRgFu7QmgF3hbwqhOf1JDdBB0bZ3u
0rFIrCASU3oO0PjBp1AdQwnOR4JymcMnO86werm3uu5P0LmEg1AEZBwp+jqf1iEMwj22kYJpOIVM
+sftuHXhJShdNOi9Ay4VBX0swvNEjxjH9L8qcTkT4WbsHkdffCHAToYkLfnzYVejlM7GmiwcxS82
ZC1fBWZ9XPlSbvRazRU0QTKK7VrUGv/U4UJGAHXtIu8FLwkviWPCENZTQ78/uyjYR+FXlFqq4RqK
DqomnE/kARrYKX+dP1iHLioowU7VsKm2MU1TkgkeTTyBUBghfHWbmQBYC6TP/lt6rKGFExGLQ+31
nG04TviwtiszjULynetEjDamEfDJlke3PQR4Az4NN3/xQFBMOKjwCsg+aUvHlBgSBc6xCII0PrL5
N/GuOJZ2rAz4KwK/ATaSNtOf6HsbAb3FEXiHiKJ1jC2ffBtNEM5aubkv+7ZrfwsOMUsHRlMWlBgo
g+n8jsSsWQCCSJFdvJtZcvkXZo72PjhZTxUlhZpsokNe3rEJlu00fyIt4aLJrrP2xFyo3+189vvQ
UNGyXcLnWMu0FHxLSgwVbectrXdfuCUgZa39epYWB3XYKxJZfnmcBld584wl98XAT48zocv4h5SQ
S9LK8X/8X4HH5KEmNv5nI9QFaTMkUw59vptSRsjeA8V4xR1akuXvyTZGsBbhgxurNWKfgeCYPsQ/
bwo8mH9rF5Tcn0+NhKkRMs3ZRJLDHMCTFQbsfZ9oBCvgZCT1A45Gg3Pyy0w+4D7sUQtYkE1oxLv7
WjlgngL5/0rkfaztsyYeWL8fGcFcQEO5DnKYgTb6+W0YicJ0zBmnMoNUQKhMqAse5dSYOEV2k5c5
7D92dG4HoxqjzPEzZIeGz49+Al3uwScKbk5H5/t3e7J7JGDVxixuNoQyFE4G1BG6Y623/riiRdKw
E4ys9QWXjeKgd5dyrSlNQAzgAC6Fhw/0Q+ad8CbrVf7hVLGUBjwTkGCUY267T5R0GqjCLVjPpjj1
/Dh7nwAjGXd9eeC+/dhsbCFO0X4nVv62007Jl4z0H/dSNlaozEEYfeYaPiHjKAjb9J5itEvHPat1
+qdUy2GxAFQdwenXO8vr/y3dDCH5Wd0YV/OfNn3Dvuj7DTTmZyEWcwkObWGmaexnVx5B9ExrQzwl
t2kIIbEJPKz2iBmMFcuQXjZNT3pL1xraZYAYKTsXzo9DoBBKm/rkrweZ0VSLv4TLaODh4j/sbYfm
93fS/pbxzLTXDy6XquvjYy4urZpUqGvtap5QZtq4eRBLnJXzNJpxoTcogYJber1DFRg2R0jdP4Wr
xwxJqTXgw4I4tJcvQGIpeNtKcYz0GMpjnaf8usvy8kHsNRcFp9zzGKDVNCljpOyaSxxitxPm/BVU
nEXMD7khVOWyhKg7MtpJNGuJUFXBgwtpJKMKsRfF0b1B0HCNYagyNB/cch34opYk3CvfAysVEWob
w/2TQFmKEWEXIHTmjfcpYo4xfFcSjPCNRcwazQ3LZSDYezXqRYsSSwaqt3mk5gMJyG6HhZ5VLOrT
ZJJ8jEoZhox4u+q3bhX31Y1am9lpuhRX+9AbP/Hf5/EL3kMIY/hJhBCwQASxpcZNatosAnPSv6c2
iGRNbPcKjVyJ4haSdpiT0uBS4Wh+R9baho9w2MKG4Isg1W7fLCl6m79msSTniNv1HP7CpoeUshUB
zo1tOThNHQWG4dS4X5/kDSomzQkEjanbQJvZ3AcCTFNLvu2IGvw+7LKA3TrYaRj72Zajb/Flv7tG
gONwAqJsoqEwWQGCWWbvPjTAy8yYx7W/WTGANXJjaq/VH3lIdhvUzrMax+1AZ3wZjIwaZmvEWmBW
B6skCsarwKpsROEZcObWgZwCJvUp9A9p1LhKEMSfz9iDkvLCFFeRgNZrQKVVtO8a/6xvusU64+6U
fYfiFeZzZSzLkQrk6b47HyZqe56R/fNfRgLIfkVUP40crQeRpW9MAMRdO4oiolVoQVFFJH4mvoXR
zJx1p0a6HaNQ2rcb2qEWOmyF1qilIbPPY9uDzdADZLWeGxdS3FOd1dY+NnmQ+y8aY94orJfzN7Ow
O6vKNozdYO0A9wUx2S6x9ePAtH87Jm3DTiAdBwTJbMfLl2HTUe2K+Vzd3Hj88V0U8eKvQIr4Px2d
L8/O5Yagu9jjcmNaNjm5aI9YvX2YoxgQGNKhVhPmS8EZ76zxkRLlDkYgUtjnVlUvNwk1IhujsTM6
aQxxobmXmHgO+Ba8jxL2LjPckEslvtP+ibuUhlw/o9d3+nwEixz6n2jbo07LKgijfDBbHLeL72di
DMnexMT6Doh/M/CDgfG5lS8oxZ+Fmd5gu6l1etBlV8P1uEYP7OgcLxZSgWR9pITWGXKdpJ3mLzz1
M4wG3R//ocjcoScckY5UW8O1nAGCsnOjOJa7cjQURdtTACyHiXLTeTO1wi84NXb9Z8ZLwiQpnNg2
KB+ebLV9hnOt1mZ54Ej7mVwycMQlzrlrcyAnwKwyOd5QL0E6IY+kd4V1RdXcjybPmbCSsqIxiIUT
42oxfIZFlhOuJAGzUtY2RVbgaldCjEiCSjTkxesHQhacmC6LCG0RrUIUYIZK3Lp8jDqVXMpX1Dpk
iBxRuV2iffm3iHc0YFpoWwRaeZt9ww/8Zk4PGduUnMSkzUKrOLukchwISCFi2zpCC6HW5ZHxNL+1
CQgvwT4r1/YIUWWcujGDrBiNsdvqd80WzgtBJEynxnBs88qcHDWJVdRs/360ShZuJc4q73NtPyS0
qBFkauh18G9Qc+nqZW/Q4IX37kOfkp8VTjawP7BzP1AunTj/e82Dx1kNLaR+cCjoaPDQ6joaTxpl
/wwiYwNIKTh5dir+ZkzaODj+s5dbbZ7+xhAmqQsjFYOCzcQWyuhI/xrQ55IxT+6OXS3GNfmbukD9
tIMMZaudMLmHZeYh4jxIT9cFaPOmFdZOJyQ1PlL1OZUj5+1Lvo1I2sBYLgRsolhfqyR6LLIATZF/
0KtxT1SjTsgqIs9QQddgNGImLa6sppRa4U6sPAdDQRYqu5X+5ueBp8fYb15asAzMvYqeXi9b/R6Y
ZxtYx60td88qgKoYSMwZ0uFzBUPA7s/KgE7/jZ06TKXYlxuNDx55leHhwbsoeNQn9oiUw8OX8SUl
MAFlDTZJBmkarD0GiXJaXl5lOZlcTYz4d1QRpQDYk+cEu3jZMdOyHzT9N99ayX75Pm+wZlmPWPr6
XYJRD2GXtRNW8xSUi0mVVNlikpBQ8znll8Nuyo+mnfR3G67rLY6kwuQ5UnBn4e4VbXxaBitg7wnC
+TJRoLY33nth2FUft+ZZaPy4wEHmv1/0OLNHsqEYHnvwltVApEomBZgWiP23lt1shM8iFspi5PpM
Pz3ZPl5jkmBdx/1BgVwWjqlHTlHEgAR6OySU8rGe4a8AWEAkE/z7DEwep34Hyn+vUG9ByMNxk833
nMC0h/7ql86wW4xfVB3fCIw+HdZKRBXbaanAhaQSA/3zezZekjt6Z/Ya16IYjAHiCTac2/U4VzRf
ezI0yRmoso4M0SgDhzc2RzU1Y5Orr+jmSlAsN0oh+HTzqNkoBssnlcVdu7SL2MjlUeBwXgGlum/i
vf/XupY3ALKDBlGMcsWQ2kyi5eTOu7O48KcCLs8VhubHikN5CZSOWLrTBv/bV1PjHank+u2pMpCd
2sgqokbG2p3Zt279pc6n+XE6p8L6/zLrBBREAoqQ1it+gboCkgMYK3i9NKc0VkK7CREBHOE5XhuU
6B+QGX8k1r6JpjmNbtO+1mtMiTj1la0s7rBRq36orQYN38bUcouRGSeFcdsu2sS4e3gfnJKR6oQI
KdKXu7nzSZYKp4LtwOm98WRNYygnVbCwvNUJGAYI4YZSR52XI14vLF4N7C3tVEeLJ79lUJ1s6CUK
pyndLdpouJGf3qCD/GBYWS/l3bgN8erdcXM3l7lpqftKfxghM7WVdoK8UYsXSUOagXPIq8g+LAzl
Pugiot35hsVAzmffIFABsA85FxeeSqU3s78rHjdMn0UhwqwQDHh8bQ5twvlhZmS6TrsBzqu7Yx4G
4ZUPbBd9z3qqSpqCsXEcQHLY/l738/N4/jG6hDtkJnQMxEjmvRGt7WJbiK9vlJoGwAgaWeYBI7uk
EWcz0biwOol83g0lrG6f7mME7X/Gn04cfdtCul+CgwAWv2kEkKj76iNMTcGd5oE+6zOAFYAKvYXk
yjamrPwsenAsmwqgODq4O1fsn/M+SqVNEgDFqWadUmHHqgVrPUsvXaU4nFx0IYZrAo/qNj0fal6P
7R+gV6JEOpwraZtlK/uOm2iPJdkDy6Oir41mBjnrs+ZEgxZoIM48i1SBLasscdCjyw+6OjliUAne
ouHZqd0IsSHK6dkjTmJf5WjmOcbJGjYwfU89uPMgY2g+E8zi3/hRoOTcfgJMBRe5A+FARUVofoP+
Y86xIRBd5B911b16LfKhOMAninbp/UUuUa96nEc31elw0H4YveCymo0L1+1YBny8reQct5ADSxq/
/AYRNm1GrIoeGzi+1b4q9mEYn6fn73rbGl3EhtoL30248+G83+MJ0ivjnMbF039pzHi4LdctS5R7
gH5XoEhI5fCsRIzdB6Ogk1mQQdrSvuYclIcYCKqcqrPQ7RYX91cZUr9ykC4QEU/591gPk8mR7v6y
7lvW5wX/uWtQlGZmrjv7nHFTv38LsFOfMLKuaj6I6aKrF+QMjgNYlZOmSYzML2APCSptBw5+sjWb
PjdDrLfEzUaIzJqxgKyw4J4mzWVjtKTOFfvupVesf93zggHT7iadF/oIlmpy4cOJtlu1syizv8jv
Ik+pl8tF3ci81iuiR+Xes8Rapbtsm6ibK5VfEAIEtcYH+tCTkNs418K7sowtpHdk0ZGy/gVSrMC+
AxBPzqiThKEwIiLPcyPQKV8kzcCYJvtIsrrTr901IGJOLsfDvdvWJ0QiWsjC5SAD17fR3EPmTVlK
9mL6rH4BM9p7xMCMJD054+8Jo3PgFQQ9cg7j5Ya544F5D88/pgeYywBZavtjWXdhUkZsEVYIcr3U
8kontKCRBrbSKZ5y0rKHEt8ZZzEkUm/pSMgkgAG1gJ/8DVUCi1x0RUwTCsv8jXQucgSoy86pfHq9
FN34YspSibFWS2KY8OQsgHP2ESH1wG69+0nHBTdorCHePysqRWAepHS3erEa91eHQpPBSyQ8RbKF
1lYMeJDOaQ7pjRfREa5DRvukDacbNa/mFYEFpX25xZ30TmfOlg0xG6cnY9fYOkWo2rPurUIbcpdO
LWjBDTNG1huOWgtxwxeThB46Vm7QZfePYJOyQ7ywu8fv0bzJkkzIgnnrwq7iu9FH52cL2etyxVV7
Kb7lNpj0C+ZLKZoZdo2tcRq8T5TUjeFst0MPHTSMgF1IlnQc3oMH0yuvbIvtAi+m334CNeR6cros
XO76yOGcCuOlFci6JZ8gfDEaLYTFCgtKMhit2ZZD/gFuaBaHbxMhIZs8ku01sdUzF8QerXG92jvF
RoXnERKdJL9Vze6f103K9H1yc0XYVtT4ncemewzRsu1oWdsYbxE7K4IG+z8I1iJXAOmqKA03r4ZF
fiLrUDZ0RvDiBiKM0lEeTvmgnSIBJAykvI97YvkQEkswlNta/AbQvHdy26srOhZLJSmXqdgWGq5N
lHkUUG/Y02W2/woC7TXCnaFkcFZdlCsCW+UsQigsNGXiX5IYc/tNgMuAVhy8gY85Q/C95QH/H+iE
y8DokMlEfDti4Ht0o8J+8jzKQBGp29u+uCX21R+Nan9n6ZjcFQ2fjlEMVB1m830UWRrcrMw41Ond
rwrDijnbPPHTEfBpwzCi7/1J2KDMwYyI+FV6/K8qx4csQikV46IYQG3NpI2cXU2NhcXCWIbGAoF1
AXq2Wt8XVbpDXho1lurWWM7iPbb0c0CXI2tKDqWSTnuEcHyBWuDpcrGYjDp39EuBjsnm9aN1lelH
v+SzV+DlHcdTz7hhLCwVCRyA51QSDDxbrfZUjoFTBJKzqyRpvKqzYnDJKSjuR+08cbTSBp2sSlXS
la3oBDfvmtWNgBq7MON8i+HzY6poHphIWqBPT/3oKey5gmPbdBn0Jz9nK1tgnBrWcOz4xNZ6n0Ow
QZOMNx2Od7yDYaL+jHtIEkVnxvPnbPkW8zmhKuKyYiCr3xK0Cl3nm/kpqqOj9Hu8ICtRWytZMZzZ
ZY6IyRWWbxKe5Wb4WyqQhxP+0EFGj4UowO2HxBkOZAr9blPP5yr7nV0QZ8uDE+VDZrccA+WSO5Bg
KEbfwov5KDhjtN6405V7xotHJBU5cQGicvOWN0+dnwCNczTxe2rVmJYkSwx493XGWr0Wb4Mrz/Iw
mHX+U9Qo0E+aOQa4dxAr5xsrMk+5ynoDcU4C55t0dErVRAwfXAv3lfi1ONNS4PZTVcpN71IZLcsH
lQQlxqpTiXls7ueO44dF6L/m//ROYqj6zZ0LLz80B5GSjI+MS5RXf9z48rcQ0A6wBpFNZAwqqeQ4
wr8AjF4nLBPC5QoL6db074IRpcQnjaE7tmoWzVgyl6UjVPxGMDYL1eoZhEf4Amc8loIh1tKl8pYq
/QdXAFYW2aoZcoqzZ2n+7EIgwX+E+y+biKaY82N7ru45qtNY5napslDyHPLbKsczdI0q3Tyatirp
UieYdnwULDokXxd5KlUiyqzd1F7ilLRVFWxdVt24G0+xaZagdp0UEjICd2WJVIdn3RM2RkCdVGcj
lx6V0a5Tg/T5ccah8btTUJ5xDVwOCHNgsRw2kztDcgJa5ZgRRphE4Ejd2blINVDfaALbdM65nBor
mAzf55ns8iWeKAviZ2rVggj6wSk98fABxIw3rHndL/Ftq9hya93/45eFbSlcNExWqbg0AlHIS1lO
NrBgNhwljEJFmepTh7ttJPEBpp8QUTJbhHEJ7LJdxwM0qmtUgh3rM2F8L94zy/NwvFndYxhxKPIG
CszqedMqbZzc+OJhXvg2q6UpYV1AeuadAk5nip5zerstFCDXROY04OneOsmfOeLOY0Lv4KkG9n37
ZopVv+pUv5Y8ddmKmr5uUPJFPXija99ThxuCArm3yHolsEDmD6DQT5+2ThCPyBTULQKjjsy8AO5s
WAl6KzIg5a7R0DddK1qcktl5qyqAlXR1wZ33pGMHwViQlmzzV47axNRz40BMBsgDBcsmadPZcB6j
kn0ndIQREB3HDRl80TZJvNHdYYZwJoqsvofBqySv98LdM63+iKMzvVKNbKWVTV3w6thl6lfLXvYc
MiVU2ucttn7jsKvGNnff3+WQdevxtmxwtnpJmmjHaxhGpTYRVEGjh36RL8PW599pYo+3VepuUl3y
Y0g5LNbyi33a5+8hUMJQripIwIvifw4a9SdXNjKAIcz6bvX5B74y3/yjqW/oCin0jytNnDkz5mXz
4ffk+orFjvlwx0GAju6hlsjNlM+VE5iAUOnz9rh8jGxLpqEjHf/q2TNs6uLEuZLix69z+MnBXV/f
YNWPIOksLYZ9XBSxYdEP2k8lBX9YWkC2+5HFrnQAxWOiSzsBDCWt3J7b73nv5fRoL0e8SKZk5FNn
K7x+H9rP/k1gl59h1v1YQ4F4Pp5MIJ9vkP8TV1SiUESiRN+n0vVL2k3jhmRaTUIjJEgRHqIy3JNN
O8nVrSszXKI+cRPx2y5wzkSMsMM327PNwHBBN2FZ1mGYUQvxnQuYVyweZ8lb+rJaL9FRmn7vyUG8
8DtauaVG0pjc0FKCK5qfm+A1a8LrO0DzlTDDBgtatUIw18ijzb2FBUrNl+SiCBJslKgyZoA4j2Qo
tgK0o8FhONimrTsdKnXCtMYVraQvaP+auG1UQo15J1YV3KHYK5lc5oDVkGBgylV2zCnCjrUeCuKb
8A9DK6qJVqM0nN1UZX2K0gmAXsdca93FFs2TCToBbhh8a5eazDfM9AR7yn7KoCH7IwAMATFcgwV5
4+704PJ21kRgALFzJoBSA1FzFe391oOxFCW0fx2P3abmMUOwKkvs4j9ee+K/BjHIBwiPGP7Zqz6d
BeA1T9I8/arWpGEYFc8ZFFwIlnyfT9gkzLNf16D0dZq/72+fc0TySlArCeaoVym5gyo9cIerEEbs
QkMXuAV5bvGufVlHwq4fun6ha5ZHFSdJTVCTk2HYmicd6Sjl1oQKJ2ukT0RSYBn1DXHPqdp7YKqN
U8a9bHXkyOlAWC8vWT5cGtgygEUIZ8IcdPzh1SqeKNo+N+N01HaMHh9A93YyzRJZLFLCxhhFuDY4
EydRYXBx+4LJxfnFhFePQ301o07/2IX6fEqjnOzgbfQXBFqwrPHfLfsqXExBbK9yzNh+af0BIdfd
gp0SsxKdSd3qoyDJDUQb5SdlS9dm+Y7LjP1QU+hygwXPOGjSfZUu7gsWKrR/NDJiAbpBlw3T5Adm
lifpPiygYPKfKXvg2eDgZAPpvd516RJOEmmAjthJ80iWA8JCIKDxLFBH7erOFmhG+sdBWYoWXE3i
ynIrJcrf2sn7vYZdxqIEvPIGd2I9TgQYoqVrAiSiW//hbXwIvR15kH7B38ICI9gzhzTTTD6SMj9C
BmYph3swiybDqT3sBjYBAc5M+GLmJSNxw68aA0TPmurwjOE/bW+gJD0veKFH6PaLt3doKTxrL6em
QBy++Dvr3qhIV+Io1+M5OlVE21mMSCAO6ttdef13KkFh9CEYXp2DAd5btX4k62RyHYwcFK9TUdlg
rtWw6eFXBmakO7Fz5FWpwcFt+r93r7eBy4Pc0m6fQuqeiO7w420HDd6p4dtVjAKjdSEw3h+Jdund
FKrfmWDIdTqer4eTKYc3vJ5qjIQagRZZ7DvjfzowIn274GcWdqVsfcqn2bMivexD9ybUCStRVWvm
zSyx0yaBJjHt1/JRppmiunDIqwL5sZc1jqO1CKddIY8IDaH5SgM4nURjZ9RpMbASiUqV+Gg5WEOY
9S70WXSCq37DhDHxLIBELbGmuwyOUcxim1rRNcrWzg71qCdUMXQtIx/5hpkX/SoZ7MZ0Lb8Ss+tk
WL2niWCcK6kF3nqt8NLDxOJO8eUUBO02Pc7Fji7zyDlb9i76fV+ZCNrgTg27AA4sDFuqb2+TdShX
7t56revPeYPa6NZB2+vyAIYlXb53yTZgzb0Yvg+KhDjgFFESblofjDUcAgy7taYhOh1zadt4EnvQ
Gc7+ZNeKffnSmfnUHYMd+mdQCHiGnxzaTerZPxXWtKErdFnETcUpimU8v5yDJlN8vurjvQcAonuX
dNaXfJSohvcq8AABjwIN2smzi/pPnZGxDehaDcga07+KERaSxoHn1339e0Z5H0t2IS7TxzK71/tD
TenRb/PJ5Glog0TI3wDw7GzLn2JJbX29LEWCOiHo8jVkWgbOOJrHi1WIF/rnwfNs0U+5pvxVAbYR
EBfTcrHCwMdvFjOIwkerxV3tL4c2Ye8Y1ZVWkw8/JIV5xoDSUBZreJF4TEeIoJaiVCPnTEDp2c3w
ignaM2w7PXEJEXKZmp8qfHfF8EkO9cOW4BKXOTcJ9pTMdXT59vripD7v2BGeMdmuFuFsqnxAeyO1
7jN6Kb+TsoK6pR7K9uWY40TD28UcA0CyMVNlGAECj24X4qEREGbnQ/4cCr0/pD34OMPCbPpmIxg8
/FNcxaKeQoZYvwnOwhP3ttixpxUz3oGxwPsU3Qa/Ttjy+5QH6YKYADVu0oYyZ9gHjtT0jO0lkbib
PTwSoSZS4r3KA1FhajvgM/L4dFXDDDn2za6lrO07wu9NMlng05KKdgkPYIam7VpCHQsKSfjGZjP0
YX/8FzJ52XTxAukJdS6RmfeDu+K+pSQhs0kL3Tqw6Mz2znHC3vKavnhJwMJu9m+FwTUcKUBSlw1p
IWs2cLNklvb3XbULykilFYsBR+QkBChhIqd3J+yJabJ/zeqaXgH46SSjNFBbiJRMpOuXB95+lb56
Hzhb59oGWxt2s3gB1RjcjZMmQb0WTnQX1A2TCB0fOKnBuidWiPUfLFSgfB8gyrfa1nZkBA4LHro1
c+ywnDt2LMypTYsuS3l4te6H4EQMGk39VMABhFyRvF+suO4doanHYkhQRvl1ahQMuQ6ixxe5nrwi
qmt8lyDnU9gkP7JmAoeXDx+8PXM1gDS20XAwJqclgHk1RqZeNl47MaUW26HeSRBV2zo5iNPW0eWJ
O2Q1+uLWyeEqqnzLMwp263UOAkAFmdJaA04zt5PoQB0bBUNhiOBDEdLLafR1sEepmVAuJX43SeQl
kxXXs5ViOqp8P2wsPypYlgcMF1aXpkE1+7mqIyo0TWpmfAAfwkD8EqssqUr1IW2LCXnytVPAXjAr
5cN/5b7HPYWRI+SM/rg5DT+60QO+JQSqA7R3teQRDCMDsVz1NDNaq8BIc2yRwkvaNK0hyYc9kr9V
ZhRW6bxFBzZZDp7z7iav81eqgHEMQjxfCtPbYQ9BccHroCqyJaH/DVnOxJPYwIAJOoPBdNx+rw59
dxiEWUFKEYCdL8FdLLpURNhjWM+QXebR6QIM8mzSMeXiJb7L5xkMF+NBtZEl4dM2bDq4NoKbTZze
7TO0lRx0Ts05dVIePd5qK+KqI3n3MkGsi/qwB9G9TDpD49AEbHusvYgT2rwyFy3hdnKGzz5fXEZ1
QzMUW8reAZti0nyyQ+dDCezVcZvr6gOPyIN7CAdRflWxS8po6ecGmyZZ5Ez/C10v3486QLFrKHqr
jJeVOK+MmHYHZ/3bsrKwqJ3hPqUbZKuL2E5eGIikk4NOJ33yuc5LiY9JaFg4BiXQSiPDW7RCiGVy
5d4eiUDi1Cvbku/ZbfVFWiSO+3jMdKWoBTQ/TjhZ3aCoUSu3QvlAALiERDUH3YKqfxM59NST7ikX
1bYf3LHZTLXWhPysQ7WPwe9eLffXjAScvnyfsfMatUlDY5NsZTx9D4b+q53ukKTJzryrwX5hwFbQ
j54m1M3VS/SupVvfyBCYg/gVtYSe00flKaeehcGQueGx9dYuz1DntZ49pSnOovsMp6gftrxVnNA0
5T7x17BoUsAmxJjOUXhp6XIecXPdClO4/B9vhdmJqNue1fO4bNmgSarKID0P/KMZ/d+7l9O6jp94
l+957wkzpRBnwpnwi/c28shb2ICfV8SNsFgd91cX/+bWg9/Dr2iyaW+mEEbf6GzGcGXi1lEcklt3
auyuQ76Y3bWBc2g2LJKx4xCUoElNyRFn+pTP8j0qzjxcAazh/lte8Yd5xhZA+ZbiK9ryIQu/6Dgb
xx15k3GViVRGiQRBOsmMoIy++TzJ6auWckhth9MKt7iL8JraVOxvKypLuJ590HCMCGvGDxVuqsVl
8O+db6/dra4i7HbX42rsKydhHcGmSgryfr3zkAvyy2K2nyynsKO6R41/JU0cmDoNR67tBvWkJACK
PKG/UEvGtD7GlmecT8n/jQ2Up5cDs6/jP546vy3LkgS3O2qMV1QTnjmAM/wto/1j+5/o/XMYS2be
CBXRSjc2zzh+P2WFKoTV9BoHvzqInoPgnlScTN9g/7dKas7VmNlYk/zyRyFLdGVXO+2TJtE5mTvT
1QZ81ItDpf5gucT+ZdS5XVReFzFTrKfSF6yVQUpcGzOKGDOye85ZAB/bPzsR6k7hjLlHLW8fJKRM
l+wFKVE5xqmj1fpgtCAbK2QZTY4Ei0RhogxN6DSMmyheXWVqZkor64aZTt7k+LdK3iYwhwW7ig1O
AIk+Vfhh1S+q5vMqUFWaxP62hfO1CK+n7rb0jG668UXtJmJ34f4FycjN1H6RkSHJJMPzMVw6+2tq
b0kJ3tqHf77sRci1tvvywRa2RscD+91sXoo/XAiUckBA9DAtPiycoTatxSqy1dZCCrjeMyJJDx7W
o0GBm9eJqj1BllUI5X3KskM7f3x1cOYi20ht6n3+swIgaEkOlnj2ZWiPwGlqcL73UCrOr9zR0g7q
YfpOdGzwh3iq8+dNgpAbYXcCWR91VM5naKcuGCFIPyXZrfQ2cAPgkX+R/gBqtpuiYtrDA72VhFh7
JeiGhTzHmiSnrhQuFwou3FM61gSHPDTFXVoZ8UoHHuwRoFXllA+CEayuTMRkNRRntL6Be5jEF5eb
NWavkrVXinHaZGyddJljf7AqPYxApUD2TybNpDDFd328HKdpgu807yg0IKYa1qHXriRZi8fl/vna
rDDIbQ6UudM3am92zUzUDMWiATFQhiU1ccojHGFuq3GXPCYgpyInXl4jMPoWYJIlAY9KAKuPY0mh
dO3KBsuSKS/W9U+vjuDZMTa9YSGEehUJng65rny9uRcSprHqL4V7s2HQNo95JTEPpK67MiugU9zM
FWDK8RfQ2zT8TdDvvXMLSiFxJJr9s4xf19z9XVng9j0E959VnL+4jzYYaNi4R9vQIRKVkbqRxfcB
iqqK5sxyJfTxtF5GY+UmQQdVRvb1hFTYy73pKLnBsxS1cchzIStaKs5Xj6SnzGADTzAC4I86r+O/
fw/GNq93HN1K7K3GID6c2la9kXhpFELnIb9XVnmDeltS3Pt3PXOipm7oTPxP7IAj9MpEN7rKMZ5A
vov6pQLQq3Bl7yIm1JSLqyhORyrgW27wA0KvFcQd3vIdtndjx8mRWyzTRyqBevJgjE7T3Lfr8YsL
ka/7VghgntQHWGf+HR1RaBf5gC1TPsNaZW1AT6VJpsdMMTmop2fx3lvgn2NrWbw3sx7G+OekL+VM
omhR5zSP1OpAMbuqVMI/lPSIB36RlUWHxuPmFi4dxV5z/y+QHR13SzEspGK8iu90B/07EQjMXupN
KabBVwJeqyRzwhV9XVfQvCpPgYxVmAUDUPc+40HGtKK6p6pxv8vDrNOD/HsYnE4irxlSzeBJXwah
Gjdkc2VOenNX3yOKBqyyySz8vCI4INX20o8XPseFb34zafd1zk0mUcEpeD3YYWhVz+udc8vS0PRT
gNcq6ZZ2hkBiakNE5ISiS8XccA0JTCDdyqjjmEVpl0Fn9YV/nNgawAOBBJ50Ag+CRsHTz17U3pqX
MHbRK+55pc0Mcbyvi4XjMUTIhEbJFGhaPeNeO7cYfMWhm0PIhu1AhZNqa5x9pMqa4EHD7CG/XoHO
rJ3zTltr5mm7Ks5BLvJlyDIuzSWFxeBbEbksGdm+G46jpxdSjTZqtuvxFbtwVW2Hbzeqp60tylEd
GUb6j6rp4m6Cg81W90n8qht0ZJzG8OEh7DXHQZz4xWLvW4aK304Ssckc3lTzSOy9qASzQ8F9nKRJ
hVQDxcXO/5JIjLO0zjbD3rDb915fXM1Tt/2zSwZq2P1YKpQEtkjM97DxfsE0j29fneWBb0ENgQcp
wmRBjS9MfkSmIgieo6t+g93COQPXaCdZ5lshBnHhBoKvhj5ozLxoTx+uUVjZKIcG4ex2ItOcicvC
m+F5cCWT7cALc9bpwcd0QVvYpvExS4STMxwxvJQYMMIyEnJuVjXSZb0JKX97W9L1b4wP2LGM+rx2
WZ0mDaX158mBjP8NHkRIB24DQTYybXEN1295p7c+nOw7aDZxJB+J+TNsH++J6nf9mWQLVuDtKvEO
DCXhbIvyWyLhBwsACzpKLR2PcuLhS7ICagSN7uSer0CeoPgj7Gv2En9ywMHJHcnNR7zvhTsqIr3i
UUFwM4Wjh17/Af9JBF4i82eRkoSZcRhQTOKWJ5MRCTmE1kbMpVQ4wFjIGwj3T6WEbMz5WaPfy6kT
SvJ921iudVO0pR6MVEbEYSV10U66LTSvM5uxgYKXvfkU3y5kKYXISYknTJ1KYPNTojHHuApAwDut
TfnGA4fz/XEE2MicxEIWH030odQgal2s3K5Ya9CuNXnT8eh4WHP0XoyKcHJb/DtISIpjc871rP6i
74nStC/A/aE9F571Pztg8N172gYU7+uevcPgs+FkSMu5TrCIuujdepC84jgu4IjsIFCFiL9ro8nt
1AzfypEzOVbyqDOuj2VnRaY/3Jv1V4RFQ+Re4QM/djNA3yzrZwwOH+yuCjmCqTiy8Jx8Ms7nI0s2
NnTuYSES0Gev93glH31cQgSM4LWl/kgBq1xPcklWsHIP2G+RcV6y7l6Z1/6OBSchvYW6Ce7YudKw
kk5mHGcx1Jaamv0xrtCComN4x++nyU/se6gccWh+DFk7ZbdR46V+MFaRn3bwltccDpbcPs7jVjp9
k252mgWLN3Ca1dL6sji80VPP/iiLITvizdlxwd/S9uDfZaJ5QloGcjnf8OsjtgaQwqhsbHrxZRT3
djMR7DFWiyffhFAONS+iCAByuTPhjuJ9Oe91v1dJtq6YdftAHlgZZ9lATI/px0/3oVjal6TNBqIO
O4n0tvHxFO4bhLLSzbo2Vv2nejCJix5PFIVWEp04OFsV6UK2kCTW2M7bry1WX1NbHn5FW0szFlDY
0DIzSbXWb+GIGDNZFmO7weYWb45sygiu2XogL+0Jr2fsK9VrEYsru0/pYGgqOf5ocOtszTXacqN9
SfFyBPNau+MHYgNxVnqo7X9+tcRrQEhZcCNJt7YXXNlv0szsnRGEAJfeRbzMUid9jz/ybEwhG2jb
MXdpnFBLVmfJ9ndKtYMjPpmCsYSdCyxYzJY/lKrkpc3fdLFZVxrUpbE1KNMYHK+bTWplOSk/QE4c
jOnHFty8G4jZaQqLK1sObyI0vc04KWchtl02bOlkcW0WhtWFV7z5jplPidqJOJIuvbG8R2Cti96Y
ZKWrezfbUTFmCqL3O71+xPuxCjw9e8Krdk5kktT7vnv8AkPE3BLL7xJjc63dPiKVYSdkr0hDX406
0NTeGxV53FZpEwu9XIJ45vxeZ0w7+dNP+JIGbJWLtkXAwGeLL31FweHyjx5+ZAt4wAPgMOMN8pOL
xPPMwLFcNoL+USVLs71hVjQB02CK3pKCHJKhkx/lRKI2HSvLHQS+Rblwgi0RmUZ760OMchlpaV5D
dliao084CPO2A3FA3CeGBoWbklBkXk8vXNzjtWfmBXClUt0+oOP86ifdnYw++r/PLbw6BkgaIyvK
l+1JdysALWXZ8HuuvqlXYf/M73rkqv9Q4Nm3PsCBa/VUD7re590YtGp9XHO+9JMt8wcy7Z0sik7/
W77DFwT56lr/V4l6mT9zUk5gmc1L8WPlvDM/gVUAo7uP4nElNJ3Je4qwWDY/cLvcErTxh7x/qjLn
wFlv/az1xxngsVXrveIy1h8KARrzxTLe20MJUslHpYaefXK3jsQKmFfKpWgl9P6NRTa8o8bjloUX
hDqeqiBi4Kgi1Jf5qBG3Zn+75aamGVKqn/tZSYuUM99FiGB0bzQYNzEStt3/kdoPomDKyZOkPd8T
xP4as4nXwMNUDB4Xa99oqNtDtA3GDZ9+gxm1b7/doJacEz4Rg6FjahBodiQdUVBpCAU8d7spOSzD
WByiPpsziUOXteNdKlkJ2q9nmGaXitE7eWhrVIvS62zlixWeW/A0jaQ4QhXDFr4+31j21siXBanw
+PwwqwYyS94RR46181rVAF8WrA0YGgW05oAmB+sz6nRiFME+2Ifii2PqKP5WtuoVOgPeyU3+gtGA
47xSddrt3jOAcGfzdJtVvCJaW/ui7UmFqtYOaFfKTaCDqGWD8EAKI5DFGC8q9apJU/HzqyLMc4b9
5g8oKOM3gL5SBCV1WcBN3pAKGkqLdATOACGTVAEYtcJpT8rjYSMGW/WXz61sJZU+AFaSRc8559PY
e7Awef0W201VOSB+WYmtJNq6xmIxalCPf/tys3NyufTiF4UECJlBf0gh+tDc34ceJmZtGADIhgKB
Kx5+iFMGQ5vXHq12z8sz2b4Qm/VNw3/Nl05lfJnHuJBjbO+OCtTxRAF4jcOW60cIyG7PzFdwCm6O
uqiTY1bmDIINKM6KvT720dwh4gEEVqtFG4Z7MBuyQQo6oWtdXZL1lBWar85mrDiKHfaAEjuaDzNz
7Yz1lArmNHLdxldVgsAp0UL4FsJLIv4sbgvJUp27w0Q2gmSg8qMsdfqAX5nPhxTp0rol+ajy12IE
iw1Sa1BKjArJVE3+3DJImGYPr2NfwCghaukIINoYpjraXyh+Bo2B460EgmIQy/ZpELFEMl1X8eU8
FNiVjH5imbaSjH0+j5YteWGNEWMzVOzjEF4QdBRpsSt7AGxEOC9uI2e110RsYGYa6EKjPYHucr9j
l4PItlEOFqkmBh3Au1cdOssiD3O4i2UvAcCP2vp0JL0fT4RcIQe6v+3DQMeXEaVXzDpXsUk51cEz
PwrbdK9yCeLotda41H7U0AoH9GutBtXUxIh+39jk2KpGgyRsxktrjFw8HBCQVtR4G9dzO2ge4Azs
mI5Sq4HiVQrfGSCEYpmVSbvep0ReEC851UDIs4q1O3u4j96cali2knzDuvPyJZLhS3uowms3rRkx
RGY6JFX8SjA+zt6Qk5+zCIEk9IhfhG5K46tCWnkFS0o6aBWE2m8eiX7Nf80zMLV4insBVtjvZjYv
bF5X6TLVcgLi6HxhnzXYyDCvkR0Qsh23viwdtWFiNQcH/pN5Tamf/d4HyGN9nXc/d+ZzcYDtJhUA
3QxKIyCVQKow1y90tV2XqWaNk19cpshg+krwfq8hpQMD5ZT016Nd29ZDDyRbZ4byRkdXTPtVnqCy
1wFjonm5/EC5KuLvILz6LvARjdM1ZetUkaEnJs+T7B/5Md7HjBecLU85jGon7HD/9LVUsoMymMaN
VNsvt44xuzuoK+k1tQnaec5mN9RyMl70EA+bZSaid0h5tuzg88XDWzPvgia7vQcTKaz3UcmbP/ut
YmJcL4fwFJZ5PtfC27FlpGwJKWRbbkQePEJcYeJvXpTE/CWiS6Qc44USAatosMU4719kUirwaK/A
sGz3A4z8t/tx097wvNtATOp8lDSayL2ehyWfOFnGUXD3a/0GpY0OAb4quGXrCjmUF6qPa5vN/MxV
Z2J97a1pMoszf6M8HQXZTlDxsW1hYy/osujZbwjxu3UguzY+ix8GiDSL3M+rAirPv+ssHQdX5Dby
NxnwokDjPTHw7b2sgAcywMkFmalVujLJCOdH72qYmbGGv64vn9pJNvDTKzzPyxmETznbWQcTV/DF
LUNwWIkIWAmeWZk6St/miR3XtnbbP9fc/c28i9s7JmHFP9wam9bHIKRyTM2/qmKyRDpczMQL9V7j
lj2TtbS7QoIHABTWEKuhuJ7gqFL0Hx01gvGAbGuEyhBKVpujkF56rkTvgyinD+gtqoe7fGnrH6/v
57VO86B0qGD5Z3RHSnh7svpt0sbX14r4VAuMlwsQqASxlwFjpvaIgNmwAGf5fJrS8dF0PJoER8WS
GkAdvXiPivX7sOWAS19PlGfUed9Xh9mdkxiyn/Vp41wATYRJGXiOiZ4P6CdbvLkN+mMR0+FuBpK4
maqHywx/EmAwqW8qTn+WBHCenynNAycMci2A0bPpNDani0Rh84BfNBbM26TFo2lfdbmppjP9vE9a
DejCi04WIes3uCCRYBf/c5y8W9rm3TqCQjkvZPBoA7guubvf0ria3m1txlhPaAVhGmOq5yRYz9FM
UOBJSiqQCl+WsL4wyIOz7xmefW9rRW+gYbRK26vkavApTDg2ceS6G7TxaT5JpzM3+m21JMoH0ITz
s0PMCKYUUfOOVVpwUn6ruExxGl2Eivg+r3U3ln0Ohe/h33CmcMm2+MosqwjL+i2cC5zEVptFY2cP
Y7U6WVYOnb71cLwjqh6BXLK3tX8O9iRramSyXYxpQ0ol5eEHNIqdYrLZ+G6d0iQObFJ/ywC+jpWJ
rVhEU03HAvW5GkQVVg4j0VwiJ43OqxL6PGQCkReqRsRnzdfL1OUxcuhHsJV0+CYCdrpYBEcQNsns
5MqOxKcpJxdw5Mbfp1fe3bRfK0YBnXxF8NsspTN1eOhutPfFPK9p0C+H4kbnPqbKuMaPGj+3loOi
pePHKfYn8IX4Xekofcgllo0/tenkUeXEZeYk91NEzqUc8+z4CeOv7a7Ebmr+ZNIjXJCtSMRArqrM
ujj+xccL/gGQwYdy/BmbXRs3WPHUjLtp7PktvDak4Zn/4tBdiifpit1VOxetJTl4rJrGKIIpuJ+t
n83/A6GQql10CcvkbdEPFXo5sNp6LqTW1DDqzQl00mTos3WB+OnEeTWkcrZrjs+fsR1QMYjDzEP5
wpnJJ9O+j8zirT7GT4cNcN9P7m6G/kHBTl69qG2Kbkv1BR3zykpJO2l30ghgnO8qLnLAWUqmARzX
M/RTv9bdj8KRkQyaEqfwl/pZpcZlo6QhG8s91Kb9oNiDFJBZD+1ehHIFBcTSjkknFjTgyLAemYcY
BFnpNpOMvx8Y4864yMIjvsWpx8s3pRvaHWX4CjJiYkatkzhuAe/TjWz7aQQoXB8q9PlBYi3VkfJX
CAJZL9mVKmPtXoCG4P1bJCf0kx4ZVs8F6Q4eHdIJvm2mz35rq6ZQ65+Vc/VErPoYo3zen1xxPKzE
TsEIodkUVZSro0wUvN2XBcG2eTvso4Rx8fPS4qByKkrTF1M1N6183QAuLtpXvzAskeK04IoohHhE
qRWJxHpfYXJswZ93F1blxm+zSDlHlA2+tLYVYqdpDWhTyn9j413sjFVDG5Bs5psYUyJQFhHkU1IO
3JqaFAXpSKLgGjlhfKM18r+j2xBrIyTSTiK4y+mdODbGAiqqXeDvdbbLP4+1O3xSCWT7LkGCYlft
qRRJ/Lqukql6G8y+XhPMyGoTavRQYXm9TfH6UyYuyMntts5km3j/H0gXebCC6radB1uIIZXFNzqX
DRxEZkZqrwCMx3Ttz+krd7XCPnvthxk0XROIVCXbWF9SpwKlPekZSf1uNIcX/fmwtxoFp/cBM9q7
F8tco8nTSzMDGLDi3p8yX1zNixo8TZ3lI3VrKSuD2JvEvgPPIgoJRcNabImc/par6zDT9M9n0oE1
y5urONKiMXLOckOd7fzve3kVAsnnn/Rv+8GG8Pk0D1LcTMVmF1zCq66arD90tHnagh2Y9cHd62HP
LelMRCxhQox9pJzJWmb8174b/5jIZ3Pa2UaVrYpoYnengTytL+/cQDO76U5o34qOPJLEbpghOIeR
54kWr4NOrWqI9IW4nTskKYD9Ef4lkahNu9wV4abd20cE8x3kowgZB5HY5B121mKfYWQT62v9eZV5
EAa8OFojFSRJzwRQVfN5V3Uf0E8qSzYCrpu+AEaqa48ZevJlZjPAtU4f2a9DGxKKxppFQKL0U2Pz
aPKaE0k5YGWOlW/xwNGLlZdPNGIWPzyjZJNF590H082g12mymd9TgoSZiHg9WU5WOeWF4fNZGi9n
DZDtG64YOtQiwCeWVrfr7oayzh+wCJcr5pKAfqCJvnxTMF7p7SGuSM5FXbbvO4OMqO9Q2I3qR5WJ
MNikZRA16VHrOUa79JPQx+D1IZll6ZnFHgw4O4UissvFd5tAPaigxtTa2MW7RVXPGOmoXMkiEF9D
EN8mShBzGH5bm0FSapS6QfFTkpr6L7Z0KoDE596dj2g3lkIN0ZpiiH92PJsK5n4Uin9hXykS9RXk
TOpoSbOwg6zjF63kTedFK4F/I5Z7DKxMOa2oYIzSD77EYMRflLM8aBctW5uoHqjdBh0gGgLpdcT+
PgCfbsKFMf0Zvf2+kRkBuUObsV5YXIom6RZYhVORV3GHCRgbijkcCF52IN57TQeaW2vektc3Zwm2
XGrN6DGdSqwlOq7AgTuRur+WCgoKmfn2LKzs4rw/cW0SUM+GsB2bOC63vrLEN6JKOb6o3v9/SnmF
QXsVw6eWWCx3arZAI2GeYoM5UKd+OZtFlIURl5uJREafDDaCaZFW7LSc/TaL3XcPmi+JGLT5s01r
Y1LAoDSsLlxGCQvGE+CW3NCrO4b5vmdAp8sy99LH4lNdieG7cJQDRjGEI7k6AxaeDIxaMsM4G1SF
kRy9jw0zwaV1EAgeUjIL9oT7VhAGoqvL4N+nWrs/aXptqVtC92hfbTzaxgLgF3Ki+edvCgNpcnzQ
tZ+wN3UAEV1KJsLzYnk3kf9hL1uiTY+rRZFOsBPsBEvtdvVb0b9sSvPF5ZM9u2LLiNC/xUUgV2Sf
VKoWMSNJi3x3VPzPmXBsBZl30PC0CRmKnClNSmW5J/huRs8Q3345nSOCsqeobwBd4tL9Bj8IwQYg
54cGxa628dSgvVrFwXy3b69GM5F7qpsmLM0SJkbKlz0e59+DACW/KtPiRG67Wv6xRyJAAUdGyb94
90O2WyytRAf1bOqynvVNBs9ZyoE1V1sIpGLjpkivtGKilITJpHK1lsBeOLSmmnpEQMcgv4/OXacp
nIMYgsf/MOeOKxJQ1zdzqWAQ0l0C9g0SGRZuIalYKixcPcEbgSAyhq5trZJnzz2JQd9Fg3KLnRXo
SrGRHvxZybEjUCZSQI8Om4A7tsxO10a4a/UnqY1bLY4ABtPf/lgEw7z8tPSy7NlCTX77KTVWoxqS
RvphBCvKvQ6eea2x9Mkn4j0ZCtbM8ldCTMYErD6nxd/6HsSG+ORALnYstksj7S8tGRNrPyp0Ened
MV06WjfTVlxXMOnS3jp/0kdTxXpDtXALvwSB2qjOHE/2Tg+/wfTc0f4Z0PizZW4m4lssXn4CF8kY
iu3ThNc+Ld+MdjYBwTCB5rQ22/8vJ6TYBs1AEWV5tvJg2RxJPC3/CpxUBcuwit+N1Q+wRT/cSWVn
FzopB/Yg8BRce8k5ntPRdkX1PKe3Fkjge7Hy1sS+estAyBrL8D5PEpzAqq1b+T479MY+fOGn/qDY
As7GhrXf7JCxdVWT/14WoUsBKxAcGo4zY4hSChuGTDkV1nryZW8w/LEkKEv9DYrBwO1qHn7/YjMr
REyM3ibEmNwEL85SwQnEgMKXpCUUmLWOC/AuU7XViEgJG10LH/HHGpIcA/QmLZgKcOrjR4FIyYAn
ubGBFqf8gHk/pIN9kGWPrlOtZYQQRtHrSozPby3TLWPkDUBeMq2dWLcgMhIi/Omf7cuMQMnZzAPa
imrt00ukBMiduxKWCNCBqM23GEqsZhrqnfxzirich1QWCqtdRNKd04Za7MEm8wsxd0FsySbd2VR9
bh8dXRn6MVRcBYypr50/0e2BrDaDigiZHAZS+iP1D5ceEk/66SG6l3PZeD3QrawWI+wEnYQqjVF/
mmYOh5QAHNF3DcNj/Y6YMAhtMh4jQMFE8fr/YDXsgzAFTFjAXSXQ5sLgd1Mj5WU20VTWr0qfpnC8
huWFAZCtuijbfVBZrtnMPTetxyyQ2cU0rYkBSwIdEACJ6Ixk0Tzs2BhP5f1VBjZBiWqwL98zhruI
aA3D4fbgRQRtFOe49Kl+TzevodyRfyBra86C9J8/5svQcThi4PC4+Sc5kpLPs2Gzc/afQXp49Qhu
LBJK6htDuLGQ0U1MULVdg7EpIt31goDBD5IizFJ4930KEr7e5fwTvXKyto9OfTlUOPPaLqEvqnsE
V01ztZWpbBPgmE1Eco8jvclsMEYB8DBJ2fYZscDE5YdA4p1dTNy0zW5kurYXrUvn/LZPtt5FeE61
D7AjpwlslrT19QFR8miFy27qyWSPC+KDvxW9pa39RfNR32barvA/HMgD7VR6x7IRnJeOxPkXc3g2
emkBsOaTDgE7FJuNYnbQAfKXbZpIH++D+aznpKAjFNXtXX6yAg5trzg4S4nfjwpy3if5jCbr9Su7
mirt6F2LYRsIbQ9gZbRmCrumfZWcgYooMq4krgEQnvQa+RmHs+jX/XUXL14IBWAm9kM6P4PLVNmf
b9wYj4+v4kqD61VKQnNlWBZ81oepla2lsGklItiHabwe1US3njmEsHTlzIq1JfidwogIzWrZvD7C
aL3ZfROU3Zygl4Yc3Us/ACVIyzQZvDo2ZS6w6YbhOi6HwiZUwIg/eX3bYaFUsiO1KnC80IaN+ju5
WCPeo37cai90Am6IFnPlpPFonFB9GmowNjIzY4G0t6OpVsWXngYoiwcoyH9ol5N8P9p/VL6bM2mB
UhCGQ8OVHqi6bCDANloJ1PjM+nmgNhgCfoSyvUckvjeZdYy7pBfsS5/DlV/TmyQdO55qDwqgeK0l
DQvZE0p0xrGUBBhHxBJvxfUutijk2q4plgSKVe5pXpGi2cUeRTGT6Zzp2pkOKlRkqppADmrnbxQv
6U3fFPIXVdkOoQm4fLSNsU3R85LWrjyTuHa5oD5eiIc8S+ku3cUJCZAjMKqPo5ndp+n3xR9z4hqE
IH3GROF6RGp1a5caigCLfLg+/GjaHU6B03Ejz+3uBjfiv5ZzPwdcEAGu+6ACzH83HCw/E7l9T9jb
NbShWprigIN0ZVQMl0O0jYEZkvIC78ezR9RSbIJNXDIVBIaIJEMfvnUjQ0bGiYl9l6nw+T3KHa9K
EMmD5hRgjXGV68SEgOZvmmN1k/R7GmWCUu9vV7WjeDf+fVUJbJtTRq0kXPkblpBRNcpMi+ano4GF
5LtON50ZXnGcawcUZZVhM+blr81zdkvziml/vkJMGMvZ9qN28wzUXBcvm2EXpb1bBDgcdUGRw+d3
VafLPyY+8AEYOEPaggkZjtvJ26m24xjcf84df4+xRUxqQ748B9s2/3rXWO6bmV4OrMfgdeeYu/8U
oE/C/ssFeAPu6mQOKOu5qryfRWZjYSLltGUs6RcOYAxFXSQcqh59qmU7n7QT2O8N6Wbwry+UTMD1
JRuCA7AN0Sf8oXVrAIJGY0gf6mdTreWZBd8+YKf6LNLEF28h9moBe+/6SINgmf0iPFJP7dh8ljlj
XdV96MMoOTFfJ3uhO3ds8yCaAs2TabFPavShrouc/hNRNYfCKRCKpsPw4OsZR3UGxHrbJF2ezqHD
Iy/h16yp/PTNFF7dZsSm3PgrBTINgCTySrkNjvrauauSWsImOQleSVHwrSDjkYeN9vUKh3cdq/iO
28MVWlnsp719oWEBlwOSGMYXJRcXgxpvgisE0P4EaBIB1FTgyzz0EEBcmThVpnmuazigHVLcQm38
pBYZWbyLQRQdQLWxkXzSTqVHIPy2omwxjcLQgtqNVMiumKpqUmhTIQl7lMzhghdg34pPp6yU5UGb
5AofUw4sgszN/Ceo1PHRGi3PIU9gzMnNfcn8ZnbIfWFF8P2e+kzW58ya6BwtRpw+jUzaxP8aBzjI
oh1YH1fjQWtTvY1nnhQEeLPAEvKydM4VCGSwyUD5BctCCHPNFX0ohlEpMA4td7J4xdM9WULpau5l
vpuaXCnzmjrto51atg90vmFcNcYV0pQVQyLeT5Q6owLdhUF5gXAF0uOOIovMdulJysULpbp/X9eO
VaCiG4U+t3XwhxZ5l6b8LI4p/k3gGtG4fnwkVlZCCVIxZapk3/QerAdcoA5gz9Pscz2BBTbN/1GQ
aNlhzWZmwTySfBSqvZkxWO6a/UET8SslMY6PbnBNUBFSzRM+QtsEuY/bdDy1pF3A+LD7eZnhxnL/
VZkS33mG33oPBa2nAzE1xeTpSMq7mKjvnvgTV5BqHozUEYkdbpTFJX/OtMBjRgyObdB2KckdAZqN
V9u2y84ulGVAAdIdDVfQsmOi1zd1fVe+DPN7/mwKi2BEABXd0H9CYH1WDciihPSKzhUUyMl+D8hW
k93u/3VjmCZht9p6boJG2iRmDP/xuU7ONZOKx5wKgrPUS9v+8u6zGvNacI1CQSZskxAXyIwQAZMU
SMGMR1uoCk3uahTMuVlljMBjPk0GBLftJIxgIa6uxoXPRppj+cDkGPtrEG4NlMZauVI2E+E+IkBp
dnmXj2/1h6ThTR6KiZtd+GlhxNFOhl5yn//3bwiZcyABhmXbCbgTqpF8aO5FEZ7XFaUVD9y8hnDu
t4qEny6JxvoA61jgEXlC0VwqXqKVJ4C7grGSaFcUAPs3A4E9dgyfX4PsxsHFzUdXFqNq/OmF63+s
wHu8ouvs9hNXt7ERnKCIw4VDREWr10hzB2mdXcSDPYtcOiR8sHsxpnEzKjBc/EBHId6VoElVQ4J6
7J9+5ihrKBLG/PNOwAmC53+F0KZpyrxISCQzwokxIZgUjwLNJjcOQWHBHB2LVCBIgJO3PIIptrqY
dVyT26YghZTR/pXh4T0JHToY8+bqLEnrNSPKT4YnUF0SVV6sNqkKb16rHhtlWjMudZa2pJe9DI9B
WgqD38YNTtSJtVncTZ2BUD/2axTIRSp+Q1Yy9OOdYbXLyoJJbYb4hmgV1TNosLA7XuVqRgZKgig6
Oe/OCva1T5UsRstio2AeXisHZOJB4icV2a0KuJFE3lrOQwnsRvSTwMBQRp/15QYGhRCzHaujJeaT
NKw9o/SONOCjzAgOUgxk2D1Da+MUaMZwnsJKNbN4mVuKopOMco+ufp7mou8Y1FrX/VCG3S9KPK6D
zKtBOiZ5tIAr8FaMFLEG2grcpdZn3sxnDtqkdh28VsgyhF6u5Lz5RIuyoAbE4a1TiEa3I3YQzKjP
0Mdh/wzBSCMxPoHHFO77UYDK7enb1nOs4ncMzLCt1hf2SAx+UErOqwAtEFpxsSB3uoAAMdzMdHhi
5mZyk1M2y1wY+pWFkmNN/3x2J1ZcGKtIQImxxnp3jygj+WGihV5jU/llVyeRBKTZZPE87er4MPTu
IOIA4UftqXP41uuHRWt4CCD9qkauPbc61g02CZbpu/DTET7uCNklGxlqOT3UIDg1tlkWkqcci94D
O0QPhTNKb+4vqfKyuNYNCeHvJEaJzjwGmBgq1CvcXyjcunsyEeS07sa5qaIkWFjwPCB2rEB29X5w
imwvI86Sd8dx/Tv4hj8HPsRUWHJwS9j8U6vzkez4FevatgbgMoDjFHBOaEq+UHZaAGSRzP0aHpE8
0ARmb9sowpbD4HtZcqyT3WGLGEvT1TAahnBp5Kjkl0QASNi6yt0nfd+WD4gLI6QlIOcShSE1OlOE
aSIOZp7WBKP2IPVWB/7XcdwWwNV/DxvdtmtJclL/GsI0uG7w91/AFsk9gDSHw4V6Gxd9ZcdI5Si/
qPS259oygOHEg3K3k3Il8wYhZwqcYYb1F1NTrCbQscqfwdQy522UWnlrfC1t4p8adAtHbGc4cMdE
c6bvX2wZwsX4AQhdAzo4RPMdRGFAtYRASymKNAO1HJ02Jpfe4iOAWbqODIPi/NX6+7Oq5jx9eN3D
BTNoEtdbjAA+5xKWNQcFsQIlc1MixFh29IO5oWGagwN6CIAE/kdv77N/zAE2ib+fHhxbPSKgJUfE
E6fkcbWqZTKqAbdPvDSwir6sQrTuLwiOQ/XSSL7b0OdaG10XIT7dijTBpH6CuGPDWUn43Eg/w+ZU
+GwJbbYEf/NHYUC7VM1sgRnrbNGhvG2tNxoe/I1LKy7lRFWakzARp6vKcMwzJk85NSPaCqCM5bUL
2pRa8snU1K8Dg0rsadX6jvF1y86C9F4sPsOgQao0ci0N3lX1yIkzLH73nN+dlRd3F4SMJQO8p9BH
iLyFvFJzQq99C1cx7Lsrp4Msuk+AfAYp9uoTuRXcyVisneAKEgtxOmfr7/vSmNN5kyUQ16rfQi5o
8exFD18JCPmGUQ4LZQITjxn0JdxrSXJ5ksdoDuwWe2VGgzXpNMimtR8MOG8DXtElohK1OsAnkrXf
4RftYIWyAJezrhCR3sHVy9E8mCA8bglT3sYsAN1tKSXdM+5TDhd4SWfebpTk97S4YIUurVMU/4Ko
R5UbeKdMIIIe6047doKJLL5EVaQOjmImSd5+BgqUgBo0PqJnv3/3g/oWBulEOtD6mqbFm242fBMb
1xd4NRRlaH/cJbUjiPXXp/a3trdfHRyaPRZrGhUSNnmURrzgFVfiirOOV68+bZM/mIqc9694BZ2d
+p7BDNChcz9O1mGBTmOGLXnRvRzSZAIEjtiUNnPImRKYtwKrXRD/npd0duX6IeoS0VCJ3JU5yqU0
j/kzP+NaIG3P+Qoc6gX+FgBUnsnmAN53uYwU2c4lBlbz3EPMPKPZpsv3tl2BGo/+/W8tTzfY+FSf
DIBVf4+IkLCvmlswGlUbmQQywpSRgx9Q0NgJnYHDqfEP/SPrVAUs32QeYVaaw+vrCw3ZzAfCHHbo
NUc4BxIHTmN3en1T1pmaPcFqr/BpKiQbIMfJY3dnLG2NtemWyLd/uBhHJ+NpeZJuO4B7I7OL0iqM
w503xVsjK5s8Vd6dtmGrcYOEzeSSMqUocXszlPeuQlXgpFGHYQupx8udlEKFAGgVDw9O4ZKvVCop
2c2YpSxihaVte1sveSnW0LuhsOTnuzTzDvMulHpYn5xLgT2rP+29TiQhJIHDWDX/gucl6IdDSl6/
ijwqYJPkbiDxVJfwTki4f+69YrFnd0DJ19nUoSn7rJnqM6NvhQO/ku+9VOD60HWZNmZonrzyxlAT
Tou/6P29WbIgO+DAIrIMYZnUXbPoXuUJkdEK+AJupjpuKlC9wZtC4Q5dvNaVfNQ9H9h3PworPbyn
WAAcBWhvbPAG6OriLqCjj8JlJpOieDGGEuDQTX13rTRCVK3HFkN60jXEewKmqFdtkw+7q7/jGCd1
nqAjvxSBx1q4f1n/OAlDmYSHAPQphl5omBqwlEwkfSiEok5KZrMKvbw6hJ/SWX+3H+3ODciTB/Ba
wA7YIjFVBD1wc7y4M2ypz9Ec7tdWwAJ6Gc0WbJ8CO0w5R5o+gyzzp2W/KbliyjOqVR8p7e10RvDf
R6dstLUWKT+1pbuqy+dJI3BSUhbVkZ12y0KRSTW6elYrGEs83xzTgfiHuZKIG93M89tFQScfjvEH
nSbXYPh5Z8uiYWY+ZflkRosLIFjt5ZmcLAgkPGun0KcXQQEwAx4v3qMqmRsUZBjI2D8JmAeAZ6Pt
M2GjEnzqNB4JQjXKrhpfP68JZFhOPJPiKu1Vg/ajv9CIp0lec3FO3WnDaugwxWjP9ydjujYjW60/
axOmlyZphLUCnHg2z2B3CKs+/CnpLquObctodPE7Snr8N/oiGhExbaTJArnaUKZS78SIwVOJ/MG1
2T3fJaOEIbdDyHmLDVv/vUuXHY41Db96EQ0TBHGwQnR3xAnSeTEZ1Y/GEFZnrx4uKrpaUPYHQYAV
x/C05yjMEJOIF+dh5O9Uezy7twrGMr8y0UDmu1JpIJYzFNy/EYZ5IGRX0gnNMLZWvbYpG9euQCTv
1mMudXcBmXuXQdIC1cUuU+wNlrSjNOFry4izdQ8N/zSuzK9GKt5Ft32lVsiLyMpVAdNte2E/5lbk
Bap9wRjcwm+yU3m/txlNdcCUTU7I7jgwLH+UhVXjg032nLGd3d4lbSv2zp2gtDaRzWekoBjabGO9
QovUXJpwNC29jrvM9Jx7zp7ZbrTrX5uTc7VtDX0ZeC7ymWbx0ND6zEcZ0ni0FYHVVWb8WuZJC/ZS
kpLBxKwqjPMhvS16E1Hl/6u4Ru3uZ09adKhlAWp5cqe6hL5yqqdCkh9ITqeh5DxpyRJp8TD3dZV6
pW48mZzC9LLJmKQX6+SDsunIVIfwnCh+VECyxgaASkbkSuBE+ajLV5CBqiGetr8mOApMSSOYgoYH
2QaNEZq3Oxs/1uikci2nDbezHkjU1rLAdw/yTDi4gTamtel+Wqp4bGcq4+263GKuRxN6BF8pddXr
9xSMqO3oaDAwdRI7bj8kSppnf3XshPYXkKSAWBa8KY2sDrgRVggRQWkGXyxF3J7n4/iT8TubiP/4
vkYYG7rHBsDW46nLG7OOYL3nDGtbO+qg/onPgMxDwW8c4uuECwbr8ZMMPUS+f71btWjy/aZde96I
7oWMVGZcqF9SjHSjWP5enluxZ776YinLIBCEPu1EeXYOQKN6W31rD8GYhjAFG+4YAxUeD/igTgmG
RMNnoD6h9awQZelBilNJunaoFWW/zV8RfqAM9AtmDXOkrPZDk3J8/YsB1huGkpwW2SXc3OfOUqDi
niWZe6qdZCpGtxmDf/sz44Nsml2hSl/CR/QL6R1mKm53GwUL1kc+rogS4yUjjMg0/6wRyc178sRv
jOWHFW9PKaBwCAuwnPbT5BJIkhrkjr6f2ak3KzccMKUqle29esc+7TmX6QoaGGf5JQMLqaE/1Jeh
Wk86fffsOce834gMOOWcJn9eV5ddXwWTAy9PIqW0b+tz9NE0AaNw0xoKEUQbIu7HDHENMIZuaMIu
rBnhb1cWGgnobhjLw0BBZzmZ6BpUxkfpKdrNcgdt1sHnn8TNU8VmuEBXBPTziQi43xofGlj0vWeY
ggwDMWpxmMcJ6wj9vRUC0kY3iuFxiQ5AzM9lEOhqeA+/GW8BMCuXSwlRAHZAifFyGjOjxwhzIkK9
ZD8/2YSfq41VputAWpLsLoG5J52PqCowY3PKCYlHa1oBQGgYDAteH4TID3l9/WN/GpbWEnuROYP/
dHJqDhuOb8KPjPQ0TXU/vwh5f+v6HFxNtmSl12+UKGbgQhF/62XZTogxShxSk8ureixkxdumkwhy
pbxpquK2k9YYKQd+GGb56xT/ZyWOC9i335unxEOKglTMagTuMXJC3Y3dZ8ri1u6Jow5BEt3T2jjJ
rn/IbeCEJoQXXh2WUnFthQREsUhW5BZmh5DNKaHXEeJZ0dS/AHH197xHSYF8FSgigrTgC9cVUaAt
61BjadIBIUEY0GSHj7ugQeo9bGjT2pGbxWPOcs6xOzBVrVJSTxliqvUG28lYECi6F3go4tNN9g4f
Ibo6oPTpeSMcrrowPVuwnSvhMjReZDtqmwTojmSZIMTDSn+JcygjRIO4k0yJP6P36MhAfCaxri0T
HaRVG26rmosCynC1zo0DWRZLnW/IBDFFQuVM1R1ivDeR3gAvPrEQU6U4U0KECHwa7HB2/fO9QGU0
5T2wI66J3GokL3bwwb3fZ1Ex8bkOsiu2nqnbkDwZlZi0ZFwRcLQc20S2R8t+1ZzFFQk82Q2BncAt
r5KNcic3jBPCTWPCnWlMiMESQoTu34iSblAX1eyEtaNS/ZNQw4ild9S2KGZqnXWkhB4Z5hKTAidK
fMbFu+7fXgVp8I4XSArWLMIA0TxpL8tDeeKqt4QvXnJYsVCuv+oeXFDkkMSwzjXljllxc4hOkHQN
020Ns/E9Wiv7+o7b908/QYaB3vtm6UHRWcS1066batsPiLidZNYNniWmtQdL1FUiaIgr5GKKA8C0
uO502tpgRp+gvk+dj5ojNjdRcEdX2g/kIABfPCRMviq1Wz7wuN1mix3Ug14VC8hBBehMLhOUxWIE
v9zF9F+1NT/iVZx84vkbmoJZMqhA0Mb8wTZuSsGeGwdp7d933DAMQ3GeCfiTV6HwMTD/YGyAF53N
/vZw+9IGpEAEWK0eRALJmwzV7zvPWUqgMUXMzuUXOJ/nuu30VMX3KIeZsw9PvnhGHNoAxp3p/u7q
Hy8iQasDPHbGKhL6b2zJKYGCkKvUY54O8g0kdqSm/CMO1sK9fVqSrs2UroR372JCURUx1LhpCVAC
3UGiHg8f3vBsO4WnPseMjr7lugM/trixbeATUj4ht1Dqbgq0QEzXcK1XhdPs3VuoohV2tokmmTuP
TJbamsDeurVE2yGT8vj1AouM8MukqS/iDh8mhkoZLdb/dOXpQI3xD6wuFfPQiIx+s2kQKy4cg3lS
6f4We4FShiGgYjBP86XfsPX7KbnJ7XxlfjdAYeazgJWpYi0kAA+QEGihQs9xIbrPkXGhkOnZSg4A
M4J/kTlMYYCKGtiuiAkp2tXnepEH+SCD0ZoTgT56XR/QATnDbrp7QQtCRY7VGzUQijw9IYJAIrAb
3Hy1ZwKlJDbWs9oCHRAp2/I8L81JwUrgG8aOV0nm72Bv+5B2e8dx9hYZknR1bzwbJiQL61ciyQ21
Nr7jogp1n8av0DWAGuW4BoutZ5A36HqN/XOLj9saqZflxFGq5WgpNs40IuWhAd4wn16tuOi9UR/w
5kpiYaQuhregwyVnvN/LduMzqOuXWiojgRA6npvHPiK9/qvIGsp8ZjI65+KW38bvawZjdpe4pq35
whUp3m/2wDASYvMIoN0r1LSZ46KEWEiq3mR7HN7xbnaofPtHrcjUw5E/nwtVbSZvotnfoOL6timF
mrg+e90glF0kmRf7v8AdjoMbLE/E7/kKut8NPaJATKYFRRAPaJWOKqXZgES4z7UFoonoYzCdS50A
D/D1paSkHCWF1e+zym3nRwVbXYkv6fuodPgA/KlsvDBSqDY1JnS7pVjIyZnaB9yo3DVDOlPLP8Zb
lKIBULK5a7otmQ0DrU3fP3Q96x3kFHY/oaREDeFcPWePva1RYCS2ai1pUfkSY0oc7Jj2e3N+DftJ
9X9vEpMdCQ0lISHenpHor/mRFYAAoNtK9hyotEACeHh86c/+8R+fjyZmIKqNp+Enw2WLxOXoxpyP
Z6T9ITnTpJDbyXw36VkchO+O76YRW6HgGtxaGVFk7Yr/Pd52nqdzkJzHQPSppAVKXd9h+A6/Dzz3
XzrKqh0oQEKVLJC4QPRprr+S0Ao3g0FyXDvzi/sKoNoNI9n/292jkgoLC1kQ2sA7sZuRpJCiAMq0
mcq12lhPucl4NK5ievkiBde8qHTEDJy+R0bU+1a28e+HQ6zh6xQoIYjJEE+LfZrTzI6Oz1N0Qf53
SSCUs0mV6gE2abz0eOxkemJKICf1YJvfnZbMfDpfJa9XonwmnmiNr5ehvBud89ZC+hbxAA/OboiJ
hNd5CfgvFeyzLyX8R8fV2y9dGfYHEoMPk7eKPC3d1xNjkXE0jbRurWOvsHqc4wxlGm3tdl7J2O4A
yVPex73H/dHKIcb3zqwM+s93/PTy9xUMgVZnmV5cuAKkMJ59cBkXELvlq7WuHgSAUdQfe95nAqZF
j8EZR+hcF/3WBjoDtGiRYtptcxo8tgKCQlAJhiK4hXPs8GbWDj0UWfOPWgyakvV1nfV6nEBrzOPH
/648e+mX0dDo7xGdLUbIUhv1lUF835chVOl4F8413yUrFdd01xchxDa+xPFzrhrdDXTUKph3HSit
2+nvjVSF670WRtzgiEeR7ktMqxD6hTy1gQLzqW+T4fCKGwdPdcyIpvPer9JNkLvBfaQwxUOC2Qmc
thHE5gkAFojJ+2YMNRnU5QTx+ZFf7bQIBbLLbXe7c6z1J45rzNLlzevP6aR6J6oUYb1PrHp43tI9
4L3WPfX9zY9ux/BKFkJ1KqJFAK1qVvpT+hZfn6mbKz1TzUYDcEC3uNN+PjzgHKnYjh92XYFt+2mZ
OHAXKtc+ZqPqWsWElYtmwhnYDfG0b7GnnUm7dwovBYMe1nNqKrKLwSfKRvoWGqjuxQBNvuuRP91+
wJJg4I3hG5u7dvtGZbywwezf4hCjN6THwc+oXuHZbh3r0MUI1B7WrBOadeLXkYBUZNVGS+wyG+B4
CxbJ4uJ4BvhuyPWhr0+0s+HLpsQbLtW93luFlyziXAOYBe/57Hua/n3k9MSN6V/FEZlSZLAf9Q6p
H5Q8Eioa+Hqsn1WNblmO1fqvSxFYsE/oTiOwafM+z0U6EZyXB5xGHYvJg2yUxFmJPiFI28tGh5lb
NiXoUgmu93rloFmkGeU/+2ArHcbNuI/FTji3ZecRxTzM3AE04O5HnL9ruesBfh44B9hLFpCcXztr
D+7+H9yidNYLWl1o96KkiBmuEo5vsuh6X8nGKebxHm5liR60sQTQnqDpQj1niPlDabyruo2q3zGa
7MELbxmdB7u0dvP3dOV2a2wpg2rAFCL4HCrlPZ6Lgq9M0+OSHlsx94kxy5fJ0iQGmFjdZH/kma90
fJNLqgjOjgrOj/J8ZOyIPpeZbqw+WiSbr8JYHuc28DHUQ5iwKIOlYzEXEQhBi2jW+ZQCmWPCnq2g
MQJogND0XA3cLTApLzhM1dX/4j24kjP6vBhbzOqtBqxQAFpxN3pGfSEuM3qlc9+vf4Nk/x/S+1Of
H9vTB93vhjGA+jwnB3F/DI3oA+qVDvVo0U0xSpUFAFgKPTFZRlsaD/4TaYStAoEFKqUe2USqN1qR
+o6Q4TXb/AnwUj4EBDT6NTpKOCsN4cC2x6dSPnvicYBVi/wOIEb4TMNbOi/7zPfSvwZrnfOGBwhH
A9BnWLX5qM3tKv6lGtYRn3yH+K5/1FmCsS2VPnFalcoZbkw5eOSs4CsPnOS8dUKctwoCorG35vTA
OIhDPEXig2QYbr+kuHnxxi99S9efhQsoNkBO2gNuSSM7LUeeRZdQLyJ0/vVKAnwgW0cXGf7rbXhg
rf58mNhhJC0PLmvrD6h/QUGW7V/0uUR/hDXxcmlCEoT7W0nEFc058qqUTOue7IY58e1jtNid+GVy
Adjalb3fgFdIlDXjadnoYJh+zKT5zgWGUFuIKNsRP433Lugp8+bkWgM447fChyzsQTmYRHv+MMJv
Nbpl9WpSLcW2GrdTgfDgwSkwi4e6trFrfWa20Hc47HTtuYzAIlIFjP/jqXST7Cc69s1XR/E5eYfE
gVl508IKvfnT9oOSPfj2BbN99G37SlNEmHbtWToq+7u0VuCXd4O3ON2FsRA/zEBEsHxl0L9xj0uk
D1gi5oSqpAYrasr3MER8ASIx7JAu9rzZYZivnA9AJi7nNzqIBXw7TXItFj46COO1sTkxokRQmtO6
Y3c7/s0IDAGG3NgTXmp/JdLL4zoBUskzHDU9z5/vrKUVafNZEYStC/0KH7CvMhsz+//hQopvAyj+
F0USgP3Q97CGSXZiLl/Uo5OuY/OMoj/AxAHmxAL2T8jh3WZ15ctkgYKd0Llo3bu3SHKvcwxJmA+8
sqIXc1s7qSGImNXrmryDvqZtF1qcrMYQMSfPfxkj+13PEfzsrP09YntFLCHF4NKj4OTu125wft5L
OgItl5dOcIYVwHBFViPVhFwUoFAjxTfqkSiDvFAfz5M8yS2ounayhcj7Ba0zOMWTRzS6ExEsIi9c
rii+wTPyhCLiACDbVxPstd42q59qvGpZb4DJhDddFywqOTI0nQg3swLSBiIe42IJLqvPggTsxofw
Un0AH5rpUuASEuA8TvZY1K4MwKzQz3hQmgr/6gHMSWkjYzngjusKeR+AuwypNDq5gVQlg5HuOgtR
CLKbtoK6d+npMDwnNZKAyzd89jw/B7g7MWVF6nwEbIZgvtK0SeX3XrrJUkeJdZq9AUPx/dxSK/lv
SlaVkYeiduyWfWtZXU0YZazt+ZGrLPXLD209epdZCMwmK6fdwDwVuZwB+py0PQgAI9dq9t31lGW9
LrIhaPlp8SPhZR78+8y1SB597KzRU3LQ3l1Uif3a8qa2VjWNhZotFEVB3TZakgj3SWh2cIjKXaFG
0MjWGctot9FgQdH5oIHuNKV17ShN/TPSrNdi7DvjyiawojUxN89s+MnI6nuXgEqjcaRuN9ugm3do
p4ZmfTGxwQ6BPV+eH6VW0ftAKtS1dfm8EuPVajSJ9/EIdBK//vdMBop7cHEb7PsfoIox3A5faJpJ
hwQH/TS8iv4CsG/ddDW5keQc3DTyKPpPkJ8+dppFfIjM/8LESxBLY3/hnUgS4+fAo6Es/JvmNmEr
HCeF3ul86wa0oZGhWmsZacMjX2QvtiuavGOpcD4KzicJ6978EmLSLtzLqEkajNZElKbLRYiQXfAw
AT85vBQDlaRp8O1CKz691VyU5etU0af384nRPQGNEa5Ch8/z6DjwZhgOO9kilBfgw86TgIFOAGn6
TKOivF2hNdzTcddB6dn7oGPBE+fqVXOB5ZwHdY8ts2i6tRsomo0/1L1GbrxZ3WSxreCXBhf46USy
8uppfpM1Pc9vfpGmIljR6sNNlxLCWQAKJ3bkodF9UxKcp572+BVNC10RhJxDckTMp+KpJZ+y5pb+
Vsq7jt+Qpw8MmCjZOcCcBq/s9B3DoJ9LT288/TkS+g7adHYRv4akZevwlNprcFlGMiwMqj1o6Epz
RNRkpngWX/iJaBhk7e8tDOjFrYzkyiAZZUhUWoayIVZMrxY19gVHSFRnnfR5U4Su0Mlg+Yu87RC5
6MXCluTGSatIY0xcaDko7yg4kwtyZHxwPMNMLBh+ClOgw9a2hwB+bp0f9a+cHb0YYOvSKRUc158J
9eQaQJAcd64mmRRSgq9IvMshmgHu3MIH6ZO0c9VdPZBRrjdVys9cgAmvsuKkTkJb9mi2DSX+wZWk
pP26vzpKg8wM9dPVD5i+UTjn+OllndoiHRB9sWLn0rfsf2lrSbJX1hTP4AAoK1UiEFd/woErCDqR
ywTgrhN4AGPLGPU34yt88/Aq8IsGAQrxmO66pvWl18NJVmJPH+3wFjq3qqWWDoSqpYAbD6ciBOUT
HALQX3RhuBqJOXGhePMNB9Ro701XH3eziuCU8E1zbKI6tWaVwWXikAnwdchRoCgEGAZgRrErLiAe
y2ziOVnA/YogmIulSJjytwziyGh6iQGaV1oavq6tAecIT6fLzsPF75ZFA7GsoDT3hLJPXvk2mHdZ
FaGCA2bYUJPT8l/Lh0HoG8cvvP0zn3jH/oJhoZP7lTO1h/snTOj2oTq9cZRhNug+NUux8sP0ntxN
A12JqHfOnQ3jyBSwuWoBU1nMh9RJrLWLftJFvrWaeWpaLD3d3QRgWc4eSyAsYGTgBKOJJmrrxs3V
ETftbTQ7HTkuEhYxkXZOXmOALQdhw/43Vw5MkHiD/pVSSWW4nFzkDPFsRbZrr4pMUiiEaL6IR++J
tNvrSBKmDrWRcEc4dsta0VquvkX1HehQz9rdzw0YLA1aYB87YkdSiztPrL8G0OTaFaQKpJ32GDq/
1+0+5G3MeC0broYFHGOZ+cXXp4Ktk8LkzFQhDVPNRErTiKytX/u0h3tKzcgWQRSnm60zknhuO/QA
FGFOa75rN/fCLjpIRHDsKKR0knBIPl5H/ZSbL1erhHAC2Rvc7sTpgtA4F+qv9Ws2jqth2S0TTm+I
Fn4hB1BvtujFQIU1BS/k0aoRClWVsfKQGrnRHMB7CAVUWlM1idycTuLyuDMTBKrN6RQwN1gJ6nvc
jqHOgrpegsKYL19+mJqCE3icvPnloDDlHtNXcRkijDTQGGbbVI+Rgg/d2i56EojMy1FrWgOZWOXU
WSxlQcPrBqOVKPcLFi07tH+URk+wmv8/m0S8OS6W0NsxwT//P3JThpV7nPGxR9DcO9tXLASi0GxZ
jOx/j6fKQ2M97tu8RuY1awXvSWXkzS0HCShE2sNan+w2NvFLDk/K6Rgin54zVOOLVDV5dIKAlnQQ
GoesZISXOkxzGiKC8f120WW/7QTjQicpsV5f+i2BynV9rNzPTZMTPiVESyz09ZTQD9vuMafDhF9m
Qth6KWv1118zGO2Odj+1HAd2qduKYqqy2A7TVQCiPy9WinNTxHtInLdfatmvwW2UZENM0O/jxqD7
SNzmsB1SmUx5wO+mpMQpvmJIGIu6AxF92eFFSZ18RTiGOGgxABW9nxz1yncwzWGlC4M4x6ufxksX
EcZkU80r4nbdLY0MOuBJymaYW9Ba+OXU9h93SiZlHuhg+hqgs+vaQ9/NbmKPokXFmrNccZ3z3jnf
GaCbIhiZljyljTBJKKg76Pj8eAamfBSNOry0AawWqbgd1j55zb8plJFAmZyPQ05Xun07pS1hAWzE
HeUVPlRWmDbl64FhpCbQ/R1hfTM9UjxNJFgwJj/TCZfYwWYcJvVouumHQYgCtz/3oFrj6SHGW1Nh
FuzCvBcyT5YTeFjLvqSpfTULftQVlRAo2yvLycJzysI86BVubqZprOuyHcKYFhNQTZ2/VviJo2IL
GPPtVX1lWuia2CjNBk4Ze6PDZRaz+cl/BbPAeQSziVU2QjOlVnYrF/vCpTWXielbwp9UrHfEq8RW
23p896WMCwO5lbl05oj/fWjN6RRQMkyTxpyDqTWY1E4jqxUCa0Bp3+HXXOXvHDdPGNk/J8U8nHvp
5kbVLKOJ5Pcf0LkJ2mCc4prvmyY06Ec7qLmzI2btas9gfvhw3v3bKG8q+2wUFFnpgCMipynZa8Bg
CTjbtXHrg3lSzGg1SAO1dMvrpdx2au2CaMVqFcAFHm0yvm5wuGc79m6VSJWSlEsn1EbobYwQMcKM
cR2q4G/Z8O4e/JzCeDfYKzbTMuvvspzmuE9W3HdEadr9VJwWFvkeYfoqVu2Tw6X5unZP2XjV4Qxh
hSb2a77Wx2q3pZrxUEGO0lBQuBj5nba+w83/EoKUx97Lc3a2+zlM8F3NhETX3xfdm0jyv7kXuSK2
G2tu/PMXM293H57G3wYgCLIAIg3UR2KWGpGH9pheYI+1cljkUvofER+qX7+iZqTvKktCxkbjxfkn
a48xm4kAKSpxR+AU/a3Eyog1w3ed1VkudyICbj6+myIAXDpDW5jIoyVXmvSoJRE0uUnGssqFzYdX
I8iQ5Yy0ruKJEgvGKRCLFAHKTaw5yDEzchCGpIPt7PWEAVSHVh4syUj4fyKL5zoCJBBwPWm3xVve
g725uYNZ2slyFlz3usjr+GoLMbhc7fKHPfdothU54/KFmfT6RS4ocbuXOL4JUwwXItjiq8VLFIH1
XP0EdrYwkWO1p2vo9srTJbbZPqNdQUgQEv0P22B4kxm5FwdKVTIf0Z7qjmulZ/fHKc92KRCqhF9b
1dYVuV3WR8SKoQRcxNnQLMQPwRYkPZMD+Q6mqQFhAnB3J8PPELDhdjKCvriQEUoXXBHR4Jf7gOIv
592n4c6+UOT9Mlsw6BwYqLuudY0Q/r/D1MO+0WzTBRshvCUy3FO+WHQ0HNSMmijGX7AuqyDLb00e
+wb+Hj8Ve8IkCFF0bHYFtiCmUlYEQy+A0RBa1JIGEeovWYVUedTi0kYqHtkcVexM9N7j7I+IU9gB
SaAYGXYX7deP4/KqE+JmqWfyuiaeQz6C43uoEJ/9KW57hi4zRpyhmhJ/A8pBuxlFOUFpXA5gIrEB
UKPnWo550F7/ZZ7mXICOerVvEBrlyMW00DpFz0myvGveo4lm1DtqIuPPAGz4nCuutQKwbUFIkHZN
P3GHjZlmy8NZ2bcSpRpMJRgvcJnk77mErA+IDWPvhTx3ZpI8NalxpdhoxqsrcCRfFnbRH3Rafk42
ctRAQRPomPaAETjUz4iQMXqKyYsGIubzjyQ5FpVrrOBx1IlvHuThl9/JlgHQBq4FXH4A76Hj2/cp
06zLomRQxQB+DnzKITAvpFbHLyMnIhrZEza25Jd6Kh6F+NQJrsK5435TIiP5Inq91Utk6sD9QJTM
j3tYFSMwA3pwwMC4UZzdaBrTaBXnrkfNZ4JjqqBbiuM84FfsIsOubfx4O31hVlPlYxd6/2A+DcsI
ZdQopq/0Kc0GBSe+fT3WJatiXMLJSmHH7Gn9EXV+oy9d8CodBuVpZjCfHFluKiGjlBjWv+HfhqcF
mrj9QDyrRTp/n2l9QTG5FJDl8p03VD0RuU7+x8CJM5BdyWtqfPBkb9SQi6d/e8b9VSlwLYbNV5Ri
jsPlFSHM8YjPHxv3l6bkFPQiOvTuvdjmOMFyHyKee/xk2tSfmgGrPZrvhAl+ph0vef61aECd1Xzs
DFjXbe9fvmnxeHrIX7EOIwAO1o6QOJPK3sNd/MmVTdLJNvWInXPvJ8R0w8YtlT4m2XNFT14OnJOZ
UhLRitQWgGVtM15lVSmtbrZMAFErxZADtfZAhmtYihVHUe/E8bw4+Emc9tTLwpdEUfqeWTszBaqA
yV5i9mXa5oC2AE6g3zt69NvLOKJC24rMXF+cL5Dl/Fl4qzzKaNOwuEfXU4+tlMZL6me6SXcviEsF
TKk4oPLV/sWoM+MB1baFUeOF+Za2p6TgbzxLgaJ7Stsugvv3jAyvl+Vj5naArOKDfMOj2+JeWDB/
OJZRVO7kbeiJmBi0q7xsl00TDIYwf7TAhh9Qj+kDgQ7dpokoM0TH6LmsLmRAm8FAy3tKDTc8nR+K
xUALiMU31BIxJfYS/SAEOgAWHUYD9/d8H6fZjqRKi5nFhg/uUGd/gNMJXDzQdrlEYkcQDmFC94ob
8egNCrJ6bH4x6+3Zaq8KXsE06FKwDuWhUCgrQcjh/+NsGCzUat8YaIcXDbZcvDZ5+3FWd92aI9pr
jutXTxK/QL0uwn8lVI4l2NThCC0RZMpwe57kApKF6qm1HBbmKg2IB8XT4J9NrkejliPibZg12WDa
mR/Iydy27Urpt99INvAorfG2Vd2L+wxisf1M93IHnNww7G+SmAjpa7ZbZZSwiZdW94IcXvkMNGt8
XhoXU3IBHcKAgStzesv2rapKWYqlsXdBuVlRMMGsFaZOEHHvbS9cisAy3BlYDlnaRmxocP6gGdl1
vzA36a32k1SvBuh1dhk3UgNPNuiYgzMnQYsXg2S0jnsQWlLAyAox292LZ6C4020+eEpuTjV3NEkw
Rcl7/CDcgitnCjzCjYX6AYr9oWc2e5+x3zANiMrx5f1ScswsoqCXk2FiKwimoj/Dyx3VfHw39Gsd
XwribfLQJQcqf6DUDogZB514980kt8UGe/JXyerY7luyzO9hTw4JrlLdDKPJGxcp5a/N4wu26GIF
CfbxjUmzVR4WyR1v7RRRtXDF/awmhte/K4sKoNzI4utkWf6qKj59dk+dYHBfZSdtp++xWSmWC2u/
OUVtCioviaFef+r19owa26qjlg+4zOpJgOza+gZatnoWQDlfSdEwx6qpBYBx5tbhmEzz/XUEnHc3
2f0umHo4O6f6qV8t9alnWcnfpsAQEDZURATs5BZZvjOhveVCTudNqkaJX3oeOzTh1LPMKKSkOHwZ
2W+Gmgm5LLbkFjR3Io+Q8gBlF4maqrmTx/yEL8dF8oaWH2G7YS8dBrH4+SAVCBSLi9EPB1d3P+m7
itFrsixxUlZxPrLO376qt3tiEjOhWRdoXu0MPCM6JzlSntBdQJsbPQCI6ENwbaUAL1HheMD92GDe
d3GxBihNFoxwJgQJNBaXtDTuPyzVJ44qgbNaLo135TRrOgpBorPl51IK4GgeBFN7XwLVdGGRCanb
V/4RQjOw+w87+KgYrJX+/ooE/T6j4wEsCLyfTkI2WUk/jULFihaZBcpdadPSn1I1PRv6gVnzYeQT
hS4pC6VS7SQ/a56g0tWO2L0KXzCPI44y/qt18V+wyS7ohXoqNICwozOzJfZFCOFnbPVGm1ZJZm3t
aZkwdDgmy8mVa6+PaGzi2EIEAAQa6o+3MAaBVbMIGr469n4/x5dFKYZ1eWOCZmuGV2uyXj12Mzvg
i6oUHSAzTJNeIjpuuOANHkErwXLuIWvPps1VZZktzsNjcKRVErSE/7BNhb3Xv/SRwf/bs2hR4ncc
FOA05wmSInQaJ8zJZJPH4uO6jlWN0B9xK7n1m6l1n4aJVg4Fno5Wn3ezyp/OuHrs8rU7eIbWoeNC
ezSKRZG06AURQSEqVTqfrCfn24aDJMq9XDXOpm6BHUiFAKXBtKtqvI21BQt+GEk5PpnqMbPqPE8b
5Vk1s1CIJEbfR5QXav0RY7DxOxFVg4iSdGIzug0v6LWSimoBYypaKa+Gtjg1Wj6RrgE+P1GzfV86
MzwgYXqa4gMT9pLQoof2PHZTUGQiHIdI/XeUoFgF+PjsWevWW+ONzbj/Uihy284VBLhlzGXczoas
ExgVOw6U3xoqbMNGhLm8/wU7xxCPhCJHQeW5aGGIREIGN0wrI9+WECTMeTSPxkrysldy+o09l1l/
PWz7odqF4GhK0ZOl+p4r17ITxMN+8pX0eS0bJYJnASu3/oXkugTn7YMSd/htaee3prS8Zwt7KF/9
RzowFmh4gj6/FwG7m/if3P4F875aX7VIw1qiqZbWW0DLW31rRxhKRKzGJU8u0Qxtwz0KYCrZAWDw
KiUESelAJ/SmyIvDxVD/IeJKZOnKSJP5229yfKsSDEyjIOvjTaz/tUeLG7l288x2/SBGfJoedzCD
w+mNHDNpO+3nRDUdXdRjSJ579dRsMUSeL56PKeX7CYLgkdf8CKa3IANqJAQPmit+ldYOBwX3PWOJ
5vViii1lJiFE9z+g60ia9Hc4kwrvvccwwPj421as6x3obrupBXMUrz1QzHSsbp9RGWTrhKP5m0OV
aabKVPij+RZA4uE6+oIaUil/c8BqxztvO8hlhXysAvyvGnbz8Qkvh4GNp2upWLzRdL+4YtBOyWtm
GdB8Spv2aPPXEb1KU5j13zwVskvKlKO6G/3v/0kIrXwGkTHLOcqjVDzkszEncsdlGYZIoonbisZL
yMdeHKEahrws2+dCostP9AMJQ327cAyKFj41/B4ZksSHZTDI4SRAhpoZmLSIrnjYZsuNPDTXUg9o
NV6D90JwLI2VdHC5lV8ZBs88sdlfBsa/l4etjr2+wEVZIRkP+hYqcTCHTN9I1/B6fD53WMbtX1FW
E1FcMCZfJZgc7N8kynDK6NTGTTj2D6iN6HgqtLHedPX4sSlcZttHDDqp5teWlowDm53s9td4P4Ar
wd3c8xAQuSGMToPD/UtTSwZhEXE636oIhC6xEuVful3UK9jZtdBoAEtPTwoO/pKpiGd333MUwHHK
dlfGh8wOLqa6/4krj7G9J6LeKpRyLE9gBAj2CPQfgtWIr+mynxzzR4ZiIQ5PDRBdaStdEnaOGGGf
dQ/61XwCzTBo28OjkpoHp7GUa3sPr++EqZc6qmtR4KZLe16H3rv5JpgaBpDaIHH1CTtDMS0A8blB
P4AE+J1KUCijik3gQptZ+L/lHE1ZNY86Q942AmXaqm5T1jxd4SVDzhFvSsdzf7c0v97/o5MRVxkg
ro6m7iYiZ+T4sPhiJkGyieJRxDdTmVFw4fRCIOkNGabNlEJCJrrkMPypYe65jeiSI30h0WnETlZG
UhS3z1226jkFpRewrzegEb2FpgkTCm3XSM71PQdu2jU4J4ZwbImH0r0Jk7k8b9CWCblCG0o5llnr
fM0/v/TWpG7p4CSsxD0a2s+cNp1aDzMrPffJS3eBNakoSgVdl0Y/CKA1zJ65oKHUNj4IqA44CTGp
3anWcFSzd5fMMHkvJeexZyWBnm1qw17aE7+2PqHxZhPO/JWdVwaA1qwe6/d1phPcFNFgwYiuafW3
ep2cSaUz48RZ3rjQLEq82MlmTUQrj/ACJTm9h1y+SeXjoqYfvAX/pE2ecGG7NkvqNJUd8N9zDbc7
0qQ8Xy2ZV0mo7g2znIbrsIRGS/E7eEZdo2/iPaEEvKhfOlI8lvtYXywsNKd8FKX/gke1LEKCH4DC
Q/NbFvL2e/VGUfP8W8FGpBjO6wxaO5kOf3IoCiwyG65QWDOzOVmK8E3Zy6aTtS1gfgcJVVTZ7DRo
fMuwKj/7qJxTYeiU84UKtDjjwqQjOV9SABUO90cS/ejsN8FNRL+oJ6Sj2siHDDftG4VbttCxg2p+
iGknUjF6o/Kg7LQQSoJkrnNMa/qDxRMi02wUao81aUPxcppfU6y7ecvSNCXqw9XONbXOp8nBrL8U
rEEQTRjRpeMPoyBRTZoIR6T4/3rUNKYHHO7ES3FjmuzdJUPtfg9DjbLk7eoVZqINSLIJTwPMJEG1
WBapUz5eMTPSgGuUe7/5izJJ/aYT9EasfdNp4QXW6Y26yG5T3C6Wm24VyF1nQ1E4eXwIJWAfYoDA
Usj1bRGgUnKEJWBDoT+ulGMPJQmQfs9jadG5zueT1zAfULNo4/OvqKmbO3HDmQPo3OzNVxtQe7zZ
L4s21ky4ANWzwmlN/pYjbl49485NtYIsTPDcobkPURdBAabld/lZZW0IlNlCGy/TSxGOxZIYe2UZ
hkEHgDA+CqZWw3j87FD3mr5wvGoxCKD64FgRTH3lalj9C4pRolq9xQpQkNLx0aPtXNjqZv+gzGLu
TTZe+UjHxyY9BHDF8Zdvhr55e0bhzcpOd1jdLIl5hVjNlVI58DVK+XWjn2EKuQjBOC3oZP9rk8sb
ruvNpSfQX2kgag4Bj6OlVcN8y3pRUWkxYrXt/eQLNfkViDoQHST1h4iehQas6Q2s11ZoIYfS+rMJ
DNyQ6yYxhu+D9grpgT8zrg/Sj6pMbR67vUm6sjwW8g4/9ht+nXQA5D2iEsWt1Wb2jUFvnSTjp0Sn
acBw0QaBCa/kPPl58JD/9SfdKdAoDUQLxGE8W/gVenlErtQcpK/y/SkAqwpmBbRNf0/ubrL55km0
CZVgYohBj/ljMiGnY31M2UKPBXwqfdHp2Y7uZIgXy72hpzNcZ3j8Y4LElFa6uDOkNgzxwN9sTcPR
mklxjHkyPlBEaTy2JsfPbeXPQeEdiVTbH02n/jr7icRbC+mLGxjMcEKyomOpeTdTCybLFbhakUPu
HODdCDks5F0aD+lVu3G3MHlxVYjfzqnfRImzmRrYlPliwXX2JD37fCz+ogODAycFJUydVbct5wv3
twYhKspuiYpd12I2AlpE5pd0rVFgGuWbvFJ9UUYwJKAxpSsKaXLW1pAYXyV0Xq9/a4KlcS/edU9P
EnfECUOkMgrfO6XmOZqsMWFfPbHCm+LPTL8j3y40ELsF2grc+tgMRbSnjlNa5oIJlGVrARy2VrWq
zqcdS2vl0x5sKL24qC7qAEStmLiWBXlW22Z1kSeFh6Tgj7NgM/BbAXFg02wVfQNDYKYLSTP1s1QL
tWBR0mfGNJgDSDquPoCao/uy12AXI6n5vtpq//LcV34pUery43IzLvOZ6DysOzbFUaz3ZhNZQgbu
QAmzALIi5IBca9+zZoSr5lyTNrJlpy+xyCTKfAjUl99rxxbla/I5NJe1GZCqRqczEr4vWqkQMU3P
AuCzjKfFtFwrksSFnBhcm/GkwEIjsW7GwvHKKm2frXrBAmJV0w5gj4fmbjnNdlKSWHZeH9UjUkVE
1sppvdf7Vfefo7uoH2BWN8Nptfa+IqPfQg7iphQLTs+X9wllJ77P5pcBqoXzilTmY1xypAG3OAL4
5O076oYn25ifd/w3K/QdziTd50Qh1s2ksK/cxXp+b3GWZm8c00xefWwLOBSMDCGHMOmzCVQ+ox6/
FhdiiXD7w+W+7K8JRT/TR8uf+GspKfnN/0cgd6rj92F19OF1nXmT4yVs2u2PN4bM1LVsVNO1p5r4
p2YOeurmFuTmAAIlqsCn50yqiNYfmCOsNWgJt4VdtntsxQKy2dX7/OJVfcggIzHo0KOSxju2fmX6
1B0iMX2zAg7f3i+jExxaezlA466WadcTd9j/7Ikg0GF+kahbE+o0HLcAii9GdjzYj1xVDtC7dp/E
Tirg3xMSIbP94DBtfhKfHvVASWQb/+mWrHPEi+hQLoxXEQ2XM++3drlSDR/IXuU2sqB4KBXSw7W9
T2MLQaQdXfKoJeA84K/tYec9NOY0Lal2264sWyAELlh6QPvA7kdHCwG8wIx4gD+uFwGeN/r837cC
/Yz0UYlH7cEQLmAW7W4fPJYgYdH7ZRf12Mt2MSOYmx6dlbawT1EXXzIo1Ma3ToLW4TVimS/QOe3y
eJ79igf8A5gMOy0GFaeBPHfBoTJhMn79jGnhFF+318Q8evClKa/tob1kT3pTliTd1qgukz9qYYih
hOPBCjH6N2j1lOTUoOv+zLdQGY/mbWhFcGCFtlQoS6IMwxBUdnMgpy6gHPcBbmKULrBD9eSEq/vG
91LdfYAPC4O3ibsixEdp3QhdIj8i1o1k1uF/m61i61wj3ZocFMdPXSpIyqEEwC58RiHL8k4Z1ZsB
rowp/sEFYmpqIGrq2ZN8ATy7u3+WKUvmcvJ/DoOFihnYa8A5ftLTRnyWMwpDqmlWHdR0bocKbePb
EG0LYiPUSzlvjSEH4wGqzFXautZjRqwkzQx26YqQtSApnEJLxyMtLye+zFZ4/Qx2BLyhxtqv4ngu
aBwf5YM6tk5zTvfphBzKy2xhozAVLAsi6F3qWnjSDkWSiQsqMdihM5DzBFjoPzW6mwn1o0cIeLqK
pKkxP4gzDN/S+RuEO9MwXIHFNNe8J8mGRCRzDsJx8XpbGniOvIq+4D8HvXg7+GKfoU+k1GDGaWNN
D7h0Pccd5DYzbO+xsZ7RuUcTXmu4bn3IteqDHWPOhq5SUSXdCdF78+4aHeKyJ8+QIfyCA84ggiTb
a2eIVJYj2ZmLkJV2+2gGsPRhEdu4FmadN1g7uOcTJgWXLerbyuNtP8b498FWbdpKQGwXcIN4kW7h
GdBPxfcWkISQVvHAEy1fWQE3N3WciAiFab/GcOiipIrbLi3m8/mDaKqAn9jow/iGkgxyaSKsvMAp
aKAiuYz44TiIpMo0+ZfQZ3CEHPm1aQNLDAkKVkkOmJaqcB4bRCWj1iEv9NOSpFlBaFPQULaV7LjY
BNV09vzIZzBtlZgC0ZgJyScXlKJtVE3rL3dglFRW2UIK5/ntsZA+beUUtXjmDmKAviCEJ1aeRjKh
pUoTvHVQmIqYoOt/0oWZijDckKBj6ZmYS/RInVYHQwoYUCBIAdyWRj61RCKicBJWR+cQGlP8Iq3r
pqPcBsWpMeshAcNkgw3+A5JRTVE3u/Pm73DpWjZjMGtYVC0fxbpYOOeXbZvhOedr97a2dDePKh81
14mlxrD4dSh0ifAt22+ZYNiRmdheGJdhpmbko+iy/bOf0Te7Gzl83ltwLXwoXEWHo2XKVgHOWBiz
28sGGpjWM2EH726ytDx8PoRr++QoYaVTIZPcx9xEDJYL/PeUBz6P9xyBG+WgUK0Txa0TvC6QTNS8
y4QExUtLJf8sXA3EEURnrvlLFgwne0H30/+fWYHTjE9a3xgbispP4S+xHZJa6Q8sLrKyD7YDV/Vl
+veyH69vh4Se5pet9HWoGEyx5KrzVFjkDYJQHlVxAQLsuaRQlSfVTsNo6XvVkf9as17Cfa4/BWDX
6osHKvctyLTky4ny4Hfs+PGA+NM9H7cu8TlcO6f2dNCHIPgZWK6OnEfeICybOoBq3t7pIOoglhVa
njVfBR/QdVq7etKkEZVcUHAeIey6Nqe45A6ZADk9rMHLcnuDMfp7NigpYl7ZAOYixBnXalZPTI6F
zwKhK/azpm4RBJ/6UzUSMHimkJPW78I6s8hmGKftTaspKMQN0b+vjk5AafhKT8HomN0DXaWid0Gx
fgycumT3qGPmwte2coeKt8OovnuLlZlYdm4Mvgf6GSSEStP22c20TvHW8bgkaAhWlQvMsDFBOsbc
y1GZ+KgH9mZM9frBU6Osfur7dm9Sfqdfz7adsHA1cU424Ss7f+V47ou2C+XQpeAto1DsNH+ucjee
J5D9WsgGGXIRADIe2RNBJ1yx/ceIJDKAZSujk3VDZ9yMRgz1SP2MRHwsljtlG7Wefzo7p4bkhWDt
IY5jeszwl53lmoYMtwlcZP/AX4sb1jSlLuZ0aOyig9+E6FA+ypJAyy18nx/t+DjAs4butaeeIk6q
z8+W2V3t4Ih6NcafvaTOX2w0bkadF+CM0hYMUQzQki7HVCzUGgp3d0tmNCfC+MVsqdC8KT0tDw9m
RblSpUWrTrT0jc3Uu3bw49EbBTPMzKZCkCaYt4ZcKR6f/5iVOWKnqi07Mbi4wrTUiBUG0uR0sZBR
/8PKZEQioq8+7nFcijQ+MRn4ZC22WKGQ/dSfrIMhC66sQ1jbc67JbsGdVzPS+QPn5YOOPtKT3W1/
Idsji5/VsFDOLE9y3aohdI9a5ksX8grNcil6uns7TbrH7HW1Zk828qfHCMCpY9PxR6wPFCHInAb9
RsvO1xKNBZKsF/mrUjuNDqTRmlXigR+Wx/TBO8ddCUHPAm8j/axY64Gw6yMLSrUEnKUUTzt0sP9e
yt/5wh0WWjzvSoit/sJqZngxJzvSgJCeiJFmbdjhqn5BCMn4MD6J7XILc44SXdhER73Ff3O9UGLl
7/3MAGdaCR/LTx/5HfEeN9z5b45pa6dIrCfyO75gTL2TnD3OB9hFLXxxgDO6jyd8eIx0BBe04eCD
NvPgcA/BFTYbkGMJ2KPK41UzfntBPF9Q96pAq02oGXyremsQTSWgyTIaiKhM7Yt5jKmibNKNLdK6
t+jZkSs09YAa4sthfilJHrPOxqMTrvCqPEOYQFnFf48Pcw5VQtMTSyCeU8JTHJxwPkkY+ppVcdt1
cCx5ctuqI14Ah2Q+j4L/gnZ8KfC7V6mI8Jy+AgKIUdfXIJqjI0HmZRE628EsTzo/D84ihRASIHG3
lIpV8AdwDHMzJtSwHp9rzDLljdvP1xvvJfYkOUk6nqnoeZUgVcrxvmOMIaRNQ/Nktbx2mSs2xxZo
Ter8+sXDuMSWcqT5lqhUOOIlKqI2ap6fUEJEcAn3qYGT41KgjU1x1sZFy4wDGFfwz+rJtAEq9s2D
iijwao+zCFBXu/dFxcEQOsTnVAYqY6DaKReV5lPe6kUkhD6GKzulwafD4Rh5qm7A/aocqdXxf6+m
Ukd2eCNLOziJe0HRh7JAScROgill+haSQ53pYobYG7amU179XrPMbsO3uXinUALZqqSl31JquYrD
VN1sUnmVTuuJfZbeaWPddfflDweKmSmBt7lgkKi4ZzGVxbY5MVQuP+3ab7pNX7niGKjPrklaG/tH
MXqlFb4EcwChOt3BMXeU7rxovHhG9Yo8QoAM3iRJeHxGHcIPQnGnmMkV3gtstKVJM4HgA/skv7EW
tICwWZvLBhHm1G3x8sveciRblHse0IXNzdDjxXJa+ZsiWmfK6CU9Ctq+gMscdJ6HcB6byCwryN5e
97wHOL7Ux0/44OII8H3bWjzG5guXX/gztI1Qsa6SvTG9kTIhhsmU9F+bl0bWUN6V/tR0jRBCTgmI
6A0h+4OHmhEgTVtHk6i3zHnfFMIwWpD90t+th0wLMNeZCgGImSAgMrn++CE5cH6tjQbdUu+zh6B+
pUGCmTdzXe1FEzcgxJyvu+0EHPug7sICQ5g6KpdiiEyV30sctR9hrmyp37JNEin3ridCkKx0dZRV
IhWUNkqul4fv+7WupREwOZQGAqcr6xLQiaLoJjLQ1fh0KI/9FdOz5vf/mDLdr6kY2be60ANupSw4
RI0XiENTBzYFEOolA1uulkDbQnGBEAYS88lmp3TQuHInDEu4zubJGNhp17Ce36/BaDK9ft5q5aM1
UgX4srmN6mmI6UkdhfDAVlAtyh8IPzJLRHq4rbqRE2eOsDzYYJ3tb0OKRqfdpNMXUosYp8Tz/zfe
vGSU05HRuQ3yFhUhuD3qmydXHWk3FK1nHpIcI3lsb/yyLp+ZlWkDgx6ruH5LGHzRjD10EfVXXZzN
YsgOocTlnnlffA5k2Hj072nPcSRq7bcwVntD17O301+83SYUFw+7zrPlb4HFczgybqzJjAtYl+tO
m7+RduYhnciXT1qL7UVh5wdQRYcmkDN6tx6BZqRwWmhciKRc7Xtdh96/v4XQrCUSnGZEMxQnIYHg
RzDlKSRJg8ezNgw4rPaQSqyBabIa3HUkvu73fZsgBCaZ3B/+OJ7ozRLwbs0emNiAoE5fk6RAUlVf
UGFdhTUPLzym740qdvRFW71TrbsKLgP8bVIcb/kbANI5wn0AprnpY7Ng+lw3BxVjfioJPc3KUURX
KgdoMmKWysR+/LMo4UXVpUYRIV7kqo9x4QgsJoOGptgsRSmhW4akoteow8eL3lptEl818lkzjLEn
s2ZN0M0g2LM3KyrNvuDzI1DN2kCsScM+2vUtuKbgEP7RLPFbsm9ynWfTAwT6IqWsX6F0qFJjnNZa
26uq8NLAhZdQ96Jw8yMOK6I3pP3PoOykQywaCd2Y2p/osR6o4q3LouyOsjj5T70Zmy0+UDV8GDYb
VLIbmd4+SptiJxDUCZtN0CzkNypmeA0F6a6JoIrw6KpJWofm+l+nySTv9KzCd2MxdEptJxoincON
4VsCKhMieE2/9HsWFy1K0dcyqQc3aNUcrLkB9usHVMA8PVHHqyYyQymogjPpRWf4Rbcd/AGuyLkb
1JY1lMdK/OZ0WNxgvUnsclQ23hJzJUc5zMpOsp8sN19GmkxjNNCtf8NpzE+lNiAApGa0Bfa9p6+v
Fg+6oKRW7eEAoAayL60QFkEalF647uViOS1j7PT+sX+chU1ePBjUcX9uY0rcPyv+JrnJjd303FgC
XZOXqwdSYBvkqJJuNfhlelf5nh/JxwEll3GoGtRjAf/a2HBvdg8qRdlrgkjo+1LZ7GpgpmSBqBv4
wvVya3F7n9McMRE0g4+X5MUcj2jXVLrBud3G8nAA3cTGx5zxpbdiJbMI3nawgLtcxMxRxTmecLZF
j630jzbUMq7u8gap5/n15lYBx558Xrj6SjAjP7WAiqegsKxG8PIXlXvhPN4JC9ZmjNRMphZLTjGu
t1ZXc9bb3ZnS3iBbc0oMtY7rySNxDsQtRLRAXd+Xkuf0uivuIBL7YAhT5zlDeIvHgwGqVXun2qws
TS8ORa2H5x7sigXgGp7/FizUlR/q7EZgobS4n7lvwZz8dbqCjwtT5ohDTeAj/QjQ0/pw1enoxtkm
nZFD39QxxMdOAsposleS7RfNO2mhZKKMZCG6vCwdQDlyECPXH1Ets8m9fdG6rjy8dZMaKe1ZvLms
mRQkyV3apkRtpU4MvtWkViAD24QT5b9WwyDovpI7xJi8XQIlJ4HgBJow1emSxMvZXrlzD5VoyZH7
nBzSx3e9y+Ae60O6033RVxaPxpJdV6OtAzOlDOrL/is9aMAidin5I09d+cv+z1vkLBFVDAPDhAb3
K/wg1YAP7yKoNGcGzF5MDyo+xYqcuVZKC+vA950Yb5YOj6XBwHf4Xit5G6mbAhYxXl6xwjbWLIME
ktceAImoT+1KVFZvCJOR/HS+yZo7xpO5IraUNUFuBR42C2PwmG3rSQAvG79QQtn85wtl4CM6agIY
OnrqJmkvY5WA6G6hEGTONdkvHsHsYcz1CRO/QoIVQPOohrTqGlnRv+M3f6pr+MvmX4sMO8MWixxm
fRR4J1z1XslldVC0uaEaPOKXkKpGS29vk9BbOsC6jjnQfZMCP07n+JouS2NWFO2hGKx9Hvbo+nJ1
/4u5mGG/9xSQfFoDzAabeJn8IHaiz/qFQoYR8f81nehhSdsL3zvtTP3Pld7OP3oxg1BIRc5DOd2U
6S9NQz6vSBqpt0RVDBwHpRDGNdvi4Ovr241aJaMgDDoWWE347xoEOJUYMvSyxo7qOvGmthcVUJXF
DwZ3lMWFz7ge5JXLiT+uMwamy415A4gZb/Vml0BE3iH/qtekUOxiyjDqwhAItSO10FUSq+O896c7
V/47RpRka/VkEM9+g/4+q9ckii0ULaglK2Oxj16b1o3f6atGntKk5Q2YfdmaqrK6RjlJleFoIX0A
P/DGuAPv0NwQx1Z3AoePpXNONRmNu6rZM0WImojtXnN3+npA9IbvOm7hAEfbfxcWONZzzTogrMOi
s/7nsKAn5QymLViNDow1I7guywQI28JIp8Ndj8j9wSUK3NyOW0bbotuWtyGI/pmH2rgJl4Ug8Wl2
b+xdaxK1+HTrv9reqJwaFuSGOPQVIG+SkV+TAnUYC+nWDy9fl0unfRa05lhBTrByneIPaH3CO+FB
fNlKbEi8bvZDWc/rYrDsPxS4y0WnUuIDtl0PYhf24wYDuUNUhV2aXpxK5VkoP8ncB9l2LAwk3IV1
jicx4NMmYapi6WewBUUgSDtpkmTesb+UvWKf2wPvH5powlcAgQYNirV8EsmMVYZCqlAmodBft1//
8ryY+l+K76isLVQ3AmMiLNZDoSmqgQ8J6yBEwhimDQZ2RsWwNHte2BDDPefzI7JPVBwe5IgXm5IW
dTGBAdh2DTUTMAp5iGEBT0bHf1Lnu8QC59AjRFZ5DuTPT47hNkNLc0tbKV5bbpp63H5gU+mOjFeZ
juT35jZBe/iftr1sHNzerV3HZDN60WDWDHoDTEyAxOIelP8sGrqU6Pu2nrCptUrauL+UntGOwk7D
4ND/ZzsC3jExb7qOUCdFpHx73KnCWr8Nq7+QrufiSqE0IwnnocIxUoV2qLLePI7veaeqjrTggatv
PSzXQlMCckvkMV8zCXIUBaP9htoztFuXuvtOjvIDVkphSJeAbW7gCmEP7dJjnrWH5BrA3AVAS64u
GfKIAgzhE/NsL3Io8su/FmrKHdxNzhoYbBAhWcE7dArqc9cjcVparKzXoVL0gMOaCCd2odd1YZTx
SK+e5TH6vh55bQGXsfOLLNlk67Vs/BGl0Bnkn5QWaLhk1JCnAYe+Z0TsVpSdvGFhZSiRaFbSaDv+
3mCDdUB/fXRjrKKXZUQltl4WnndnnLpmvb+rP436HaA/AFN9LDQvC2qqRwOrMGAs05A8TzQ0kTPY
db3sM/aPfmKmiqC5BjaB9gsJDfAQEZcnvqWBj2C7+CUm3YaPor9xRaE7G8DKS+OfwDOD2PNz+B7s
N4QEd9fx3IqSz73nmkwj8wKbSvLOAMTi/BXsZDjbWYMGR6KOCAHDscITfI+WHOEKpdJm4sHNaYXI
ziar7MOyiedYhuwOKRHxxm/wYEKWl41qJ2xAN++HsW5b62C6GpGTKpw27CZQOMWiWuLnVF/9ePSC
UoOKOTByz+4qszOkNgW7gkmuG0CCpAx9ZhY+5fYqd8fu6I/zASw9+2HvMa6x5Qz+iVd8WIeSD5cG
1rjGhP58Mz2hblrVjfbfbOug91enEGOpKMqpG58pinaPqKMpHKXFUT7g8/5R/dXO0MT2dnC2GxCe
+ovKhD8KaQ/EOBKkR5Bk6PCsTvYukPHQXsvPj4U6o6x4/bT356KotKcaj7VeUKbSNOYIWijHVP+u
xVNx5PcaR4wJ5EMkXpyHAx0rBO5j+XW2tuDhvPbyw51ijD8hpetK98Dbcdi8jot2mqsRwXN+hOwU
atnIJvsoO9RsRKEsPuEsJPgunI2t4HTdo8viF9+kuS3Ruy3UGspn2qUsaSXGeOi2AJtw5wLtivnw
7B9Nu7XUzRz70qyL5ye+pGOYrEOMXKo5IfdAWpUDGt7TRbvJvg70qoi8BFLGV7pYeDrg275TM6j0
CkkleBKurSSzFAA6NxVyVUp22PNyqr2qQ7VOIDTGTwTDKCx3vZvSNRV1xFqOmOQZ9QsOCV8q6R/5
IJWX7WxOyfZlZX/8z8EyDEWCIPckbGQZHbaN5fZI9/VtiJfHkpFeH1rdqy1z0SV83EYCP4liRhmx
ZZlATlazlKphXXbY4hW2gDWzwBHl3//ZHbL6eNDI+FV9t6xDlQoDlMbwqHBx4qt0KtS3eYmMxIIV
wAwYBo2aMClG3ltzoiCj7dsf44apo9Jb4PwPhGhx7TAak57x9M+anVOBSBdhmu97wy3Vt9M4/cnO
nCvWoteIfonNEmKM42yzg+cDKngOGGm7CGM4rf14n0FNZRctiFvHYMF/lbki6EKS4ff6iijouEnU
6gOqGo27O+zsMpBIeMwF/QvuTVa1ApBqT4AOHQ65jkZp7ZzTPixeNYdLw55co1zXJGaJmo1+ZPTR
hLLysxre1kFXsEMQDuj/BPiHf8l4ZZXsdBN0S/MGRIgd1cgLUNYO4NmDeSy0RwcNLCF2DSCbmQ+F
FTYIlNpw86omv1zQ09bZFPQHZ1kyRMs98daYDpZ1bCGgZM+kGiFS1Gmq8gtuvyJwJ1WOlfvN003F
GApc7GkZpffO7XL4OrkrkFais8PwmoAG75hUoahST01puzXQx5ebGj/i6kQBvY6+LeE6v42oqxPY
CVYM4rbHy7RUomdPJaaRkHIhOQjiDJ0/kVrpEKoN8zBr0kN6Hdy9Kaszbl0iCc16GM5yR78q0aRy
wNKPMNbdi3URPj+0hEmQU6feNXArVJuW+mivk7PfbfN5996T0/BwGoicweUO5ptnTkV09WMFWrDh
Akp+lIfHw6oh7pEc8iA5feaxSPD7/Wp4HmFRmKTRA4Z0oMceJwIdc/hMFe/kiqlifkPYX/lEjM6o
PFtnk67IGIeH/2glasbnGfLMhiasjvDGW911G1l25ixlLpU8qfUK4Ermml+wjeB5WLvV7CAFsFF3
cLlmGKQt8FhN145IFhRuia8U4UK9xEJk0IAt1DpERFwMy0YX0W4XRr7pY6HF/v4YfpJ+lfKgm7ai
wDbChgDnSoppDm7nNcvIUT/MB0cVq7uaxIMP8UgilXu4EDMYOBXOwd/ELS9Ddvtu2EKdIPXqPOlf
Rip6z4l1pHl3FEOdGYqbjPHOvwWrJcPAE9i8wBgWNy72uQRaic/gSQgzAA4O97IyrIsMuqCVEGNe
1xN3LlELHk5ZlMCiiuk4Qan1jQHsBMzymm/tnrl0k/2i2wyE1eHcUHDeGYCKWXEBImRVHTExGliX
iDKaMR/YA7kxgYQbrEigr9PHWJH1KG4No5vdETk/Ov4K8m83fosERcExfG8/oPQVuDjcDGk7HHNx
jzN9WpCXCqu1AT5XQxDd7vfnDOeSwuRasgDqlk5ZgtsYtVVfFsn1z8SHKx1V5uKPXVvL0UzF9PH1
hTgdh1vGXIzIszSB3c6AEW0UFoq2w2yBJR1Cy27ibEfgepGZDpcxdEUMyCzOe9n/V/YSx6TT0hZ+
tqqiHDXnhXbVzAmM1Yp8NWwOHPs29Lg4s0CNWnyYFOKHTMBto4n2OMj+A/jZ9sEQBBVa0qQSyxMY
PmixJDrOMw3nmpFY/dfwkiBgNpVchfMvm/Cx/0YFa9PWBOyRLlBUrwEQgJUptBc0kbn7OjzzwA8i
5xjsgm8yikAX+gwZKVL0oJ/QuFJsx9ci8A2hrOf1o8gZAv2jwMRn2oQQ+QUplUsolot/hBGFsu5a
hqm4t+gv8wox/vEGSvcM0chcc1kGRpKcaG5dinFmsgi0cQL8gkGwueqhpDerb4TsR4zkRRIdNWOd
lawIq4AqIcU9OfkoSZC2n+B6QkrIefJBftn5YvR2DibVHPmBmEQeIWVpZQFhNFlimr0TMFfy0MGF
xFLFJ7h534FHEikdAoPHf58+1LtMnXn7aEX5WaOPPZO/xyU0it0YWNPeh85MhAjWDDGYLlU316HR
iW3ba5xfjkpdWP7GEBX5HkxCDdf34OdTH0OzHF4qiwGMVTdP4a+m6Q8pJTcbyD07ho6wLBo1S9Yd
ExRiJFs7ZTNbCm7TjEUF9GSBwUF7O1tGPOJP3gbCideF/Uqx7NOoNkqq5unEvYITGjzLwYKHrQE5
3NFRs4Cwys8ue2l/X4qGLnxS2qCrFTSp57LqTQCBp5kU0sDPMLygS5Rqt289QrhBdl/MU5kyuNe7
RuXRfMqLibJUdnWzW71O3j68AslN0vzNLK+Ybb+Ea4v41yQLy0U0yWoL3enO6Rq+wb5dgHQXCvcH
DWc99Gbs2tV81iY4xsCldXA/S4Bhszoy2P4NVAoplrmO35RUfTcB47gP++1gJu9rDOLtHQfvtHNU
iXPH3djOl9DCH1FNxLZEMsRPahmd/m1QbLyI3QkSjNJkjg1QPJMPTNZvecbBOXQxij2LU+BhAF08
WnwvaN89cG/XyozNeVvmnX/Eg+OFW4vFh/BBFIFWHk7pVlPFkAkMueDHGtPPa55tTLeAo+y2Ps5y
8/imJZTn4aIRrjUFE1ySEPqSHZNsB2tG39QgLB2nzhg0rTm1UC1JnmSkl/vEKN+D6UZRd5UxSeQy
LgwnUiXGLzurQkX5/gb4S9UeCBWN/wK6CIRgOZFxmXU6UQJ02bi0Lf4DbG286eHDFb6CbJaRrQqs
9HTdzaZWHklyrZ71F+Kdjpt7hyKkUD7/QQSnCIdC6WkdujB/9FMqIsx2VYgpimCwGmNJCxyiyvXa
sKMjN7xN/mWt+BO6446bQL/MBoN8TgJH7M+iSN9wbRYw/XO/GWsZULyVUtlcGFTV3g1TlnIAOhC8
JHo37TR4+mEVdcOOdDosx3FMihhCvLyk111X4x2PCS16ICcQsrO0hCIZiSRNcRxfzTeccTwCtu4C
yFnRkxgi3aI770U9H8L8hc/OItQ1vOmDjC11wqgjqtru9XVFWFUl2eFwUQ8lJX7Uhf8STZvuL+zq
/5RgogstXjXXJRfIJBDAzOFfJ0ewLHhiWJbWWCoYzl43apnIv8DrBjJLnOwMIaVSUGNTCdwR+dMo
1wqP9q8jX/kjskYTVkABPcQGyKBtow44us4lU3ZNJB8fo7y2ma0A/vCkE1uyHwXUgX4dzEtkEqYO
iDoKKVNBrlZdWAuZcoBY9flEeuTMZKlTcAHsPGzLALBAL5pfhFsM45UCjJUjuebRSxo8omA1jO9l
O2oCeIRwN07Qvl0DvI9mgKQlRx9rv7peIO3Yr+6sGT0as3srC/g99HmfdMOLj/sG9UQ5TQ77KPzv
uveybEiwWi8fddRbuzdDpd6r70tM9UR1Wm9ipFCK9468tQy4dHfOLbeWLF8kitvqHgo85g4hks+7
b9f8ONA6CM79pHpgSaofxeqRvjyIrqNTVm7rxbLkOAQ4HejLDUMpZQ5uu7LoIaaQ3IuJbzaaC8AB
4E7klLz+9X2CWpxLV70jgJSrlgepKHTWxuBLFpRA6cURuNhbQl74u5rgUrXc9u4YVWA41PIMGOt6
oAoC6kJIKGCdnxEODaWPUFmBEqM+ltNGB05qtxV48ggQNsAJyE0ofBJFt5KbDX+hQytWS8N7ztbY
6MF6wwETLjGIUkbuh2EitF0Lhp6BODIUdv7r6nh3oHXHqvYn7WLwWMaUrLFoYrwPZUeUmljoIwL1
mBUpV8g3Q/DQGi5sSXiBJxxnTdMPj35CBvRPDcO6WYTvv3YO4+UgRIuDxQS2+0k+p7Wtucye8Zqy
vltiRN5QOZFI+do9AxnIuXVJB+KMmOCuyvr53sYctbeIGkBJyLhsmZddrJ0WyZCw/hsQjSjdgXAS
RCjGK8vY7BeUveIEVRIGTbSo8NLeLf5cYNprUKRaS/hoIssyIdWU3EkrTGraqJ6SJI6gA6hj95fb
c2HU3k18S44op/doGHOcjFbdd3lE3x7CMC8XxI5j/bSIeLQR+TBwXWhWDSakqXdi+Z/XkFx2aGLh
uAzClKFwv5t99yMHZdJNWtGr4I7+5pkfoHfsyCysw3TtFeVz2/Ilt6UMTwIxivOCAL/dg4KInPg4
LKAZQHJ0/GnknmQVquHcqqKwjDWV93W8kwsbt8S6OsnUojD2ETGy3yXmdiAuTv3MQif7EThbBUUb
EKKNiyr+PQyc+4wtqYWOwDtWUjUgU/DJFi1MI/Bxt4QxG1NpyWQ9gUtsKo0Mk8msSFcVr8tI5eIA
F5JtrfJMhiRCpafyzna3IYIjRvSka9q0yPzOjFVaHkr0Kb06o8Ov/jBX8FjYsspVLaQyeOXPdZkR
w/dh2z4PcJMVnBwNoiNjwHLKXlF37s/42X0Dj9AvwUHWhH/HTiR048q5mw9M4OJzNXQ1V2qA3Ldt
ZXOBW8G2e3SmD6d/XLynzQt67BfWaSkK/o1fV9oDJFbAQ0R/t/0gyCM8eGyGD2L14uge+8U7yV6u
rEllAONefj3/RZrWqXn7mUkmf44OQBJBSp9HX5aO6Hm3Z2DCxEWHIbuALrvWD75BMSs/H5dtDD/V
nauf8ysfbQue3pX30Ki+YZ8p2kCJwGwpLdiYoF9WTU76/zmUfE7T88SCbAC9g2iJFNHVvD2dXcrD
RZK+ZF1wLLDRzNvhdi4YaomAF1HuDGHGHz/j6yLt3tJ8OnBEVa/FFIvt71pcme7hl68ViAzt+PU+
ajSqyCBvadziZlpFCDvIYroUx5iXlpzrm6+O+ZwK4R2O0liHumoh9ylqWgHxcVxHEXQhEbna/uJI
/MN02FeIF/2ZSrzkV6kNPqiqSlMIjGeeaHe8lwNDry71ftWqj7MBvEMxEsBaJEZMmsZqZDLvkP6H
J9YMWP080FG9qw8nwbiqLj2TbkKC6A5+2WSf2yFakP8XgrZJ6zC/GkA6bGC9MPjlqsUSfxnI5UNB
ZfhDHnzHdwTx8nzAa1BZmO/Y+NeS/trU1CtRmP6fOXkUbJ/84mzx4XsZjfeIXTR6Ud0HH9HpvHMb
AmRt7LDtEtU0u/gQeTd64sVC5R7rcYKw1Muyjh9VKLJYrWkgDP/ct9JcP49eL7oR7UeOlEGyFjPQ
IAwYrCWbr5xJL5aCq0CnEwfvmIvq/jx5wVvuosimDdK6PbyTmeqgkq5Gn/aym0S4LatArSRVm6lb
rGOsQSakcd2HxfxlTtS2avSxP6Qq9AFNdRJaLEcO5wRnom6zHapMLD43B5Ju/UWwVBwqJTJFVVyh
KU5PfWACeeYTVErooCAG20D5wYNKihGHK4kKQwiimWI35zpbkQdwuY6kiEKsw08C9ReahQLV1/C7
ygGuDw50lZL379XoSuhkqh/5xqDQLJWAiU46awfo7mXzErTtAdAczmuuMwPKj36EfkhVgdp6yBMY
/Xz/uJaAD5lXVMEKetBCpBmRGoBNk4yYENOzjXyfwHG/hKXb9Wvqk7qFV8zJp9eeFgmgLvf5UiYb
XBt9GAVWkeaMv5qMkiepnbasfR9UoIXBhcpPPjn7R8QQHaIKGLtOMIpsDPACTl5PPkTeEk+5nKw6
yntn/meQshxA0mA+YysEFUtqaZ3BVXj1YSsDx6coXp3Uc1fT4FQYu9hpBuHO8aSgrkDFwohMMrpn
kdNgG0Q6xL0cxyFtMArginHZvKCZiacC6O6i4ztfh5QFbowT533y7DQ9Mj02VOAintJxVzno/cVm
s6wz1dLRbN66GtKfl21jNl/TOR23rMT385EXULUF4sgXa3+TxMaTSAYivJVKgLX6njT74anlveim
fBLs4aNgxpWPt7GgLUY5/UEtYTfgBg2rav6yT2+LIxnnS+T2p+g6lenctv7xU6+M2tpz55KuwZWK
PkTGyo8zkVsB5jRQkBpN4XUQnveoGs4MSJiW4syr4LuUrRCuIwgNLMgY0BnpuCOlKDL4iumXKJeC
BMSw4tmMNWDb4uUXbcCNF+iYpeMIQoKznNm/F5gDLodF5IjOXnt8cEMtQIqSihFnCV/8xGhhKR50
ScNShnZAOERprke2pt2A2TsiQzwacbnKV2TSsJpjlAEyNuaawsztbPsju4qhMUP1r8VvT6QRpKlQ
3HkdvTgoqkVJSzETgeZ78RT6M1Hwv+kpamDtsG6EQpl1cXtlNpKB4KfUIMiCm5E8QwiLgTPWG9T6
P5BEPIq7Tufo8swdk8GpzUsW9cc9nzUreVjh8ByrL0I5/g5XLxKf7IH0J3zs9XWHPE6LeKqX9wnr
rKY4ON5miv54NYKR049gr5h9W5lUCdyMG9YGyE/cuYalTKIh2ESQ9fkKTlu93/MrHoDV4w6CPFUe
PAJmRxcIoiByw/LZLK4MBv4LQMej/89WplAVMKoZiH2TjhXulK4QQJx+vlUEMpgvO/D7sybK1kDU
g1rVNL1a824STWcyz6TKkD7Z6Fz6qZrbtN53IGz2P4fQdZXJQQBYb9az98ZCzwc5CxVAb+c5ZMPe
rfKL1KIu2JVSYNOypOtB003G2mWXEvTFdiU6VR5sTVQWWTYA1ZTAECkJd2VBDFU80cSHbhkOfAVx
mjWoTeTOB+r8DAq728rfyOtHAEIK3qxP/eGf9l+tq3JJj5tO8MpfZ5cP9wY4o37nRK40ayWzVu4I
URrz8yPepdLwzsSPPVjR3bfPjxfK6r+ymH+H5sXZvGJvjLZza2wwdt3Ri27h/8VX5v1M3mGYV4s9
STm+hHg5GqB6NX/07Fe8N+m2wYzb/I7Ix+AAD8eMeakRRWRiNL6mjrDcmSYx49uYAUTC52etcCXD
bGoxv0nBpo3e198ow2mjGYi/dGl7N9AzKgZqtLthCKzvvk3SjyrNHe4TzGCvXDnU8qFpJFZteUXa
aHB4iSffUCqL6yJBcx/RMhZ6IS5XgVRmgf/XL/Mlo+zfOrJ9eAu2KFQZblyTPJPAsFQKbormVxv/
Xb2Lcf3Pr1GSB3V3AOI4Z4EoEVewP7C7WstvgmaK71TdcememIIZzQZEDtpLjoeyms3iWuP+WhKB
vmdhSp1F9WHWScWd0wTF5JGmgDPCIZNK0FPpDjYCCPS9PSbnPBStUXMUuCOuDk7/FsBh6pLHy1cT
SFM0R4BuIP5aJGurf7jkFhm/8ejWfR9P6J5tdcSwbVVs4BRSsLFhD5FpsFJsb+OsRc8f7k7SPlit
CKJmAdFmsP75W+pf3CGciFNPF7/f8AGgMqt0avcOGsi47NzQIOlzSA9eUFdFddLIEKuPbkOCK8Tr
AbKigJ7OTph7AD9DVO5XV6ZiSSeiWvir3+A+XvGz15lhUpGdzgxayu717UJ0H62tb4+7clPG7lkm
+9a7szD9m7NRbyKdZkd0OE94Vr5n1nmz+wcbNCQNPnLvR2h1sUgrz8H87/4BtCnqhKeFHo614dMX
VaXBALkAn+Oskcpg+hdefS98qirN/bY/F2XpEGLb1w+K+AgiolUXAvv2Nn/zeQL+ckf3s9n8t1ic
RnIeY/iS5Q9p0ob6bzzWe+5t2gvq9cUIzeBCdSJGfxKBsx1WgrDG0oRj0/vKjzQxB1fcrpIIbm8e
TS6RC8pg4l4z7l1ufEz5odL+5asy3c8Kd3TAwqO48IgHgwfiMqN/hr8yCnUgWMkVUoVO6SQYV9ej
qwmOV+Zx2wWCEcyFO0BOX0N+0ZlpdAzsm5dWTz+TB5oBZZGGixMdfPjTPYuvjTQlXIJF+au0XpYy
eLpP4bCJc+hGS0m4UED2qsykACh1ETaoOsBbUdg5xFEQbb4RW+6QO/H2oG1safdz8G/6+1NQH9JH
1YIN/yE0T0y+yzQJp5hWNocwX72HW+viT74zcN+W+FX5pAuOZHcQMFhOC+AV7q8MZKosPito2khG
az/fTIHZMJBJebIqa9Catvgt1GRR2DCeCgrPHAfNgOcfV4yqMgDZK7fIxjHcfaBt+kK9qxJOf8AF
DEXThgRq2PHkDhTh5MUYLZvVEkX4nhlvoNWAvfRY2MvsBViQDjv/BHiNV3cmRWeeKdrdpcyI24e9
96B+trSsC90X+CbuHUBkV+Koek3DbOLIK0czWrgzTOlv2l0uZdkgTnMOAc89ZEG0jfdt9pjh3eiz
Rn0hFZy9pWDH1ya7oCvudvtWCAaC5Dm8jjJ7OkTmFbcSGFNQNQFih0mS9IQdNuzO+b8aPXI4HCG1
MuO2hUei8Ulg8tnK1bURxsd7R/Uzha+QEfj3Aff5CKdGt+tP88RKVLO1WHFf/6tmz7UdlyXC+ERT
3Wdrrt36kvAFneOd+9EGBsZO7PG4AaGE40di26YwQLVHXAQDHtELWOF/gG311cie//eCrX/Cr/Aj
j5w/dtERs1PdX+Xryv8k5zJLBpifbY7shlqd+pLVvx+qla9MmROmfTxFigfYSQCZBBXkAjwo8PwR
o6jJe8PAJk2wqn4RD3JL/HQacOn8DpyqUzLKD87eyPRNGUE1VjZ5q8nKK9cnP/mkg0Nvpd2QcoH0
+az9fT1++PfZo5PLI0n7dL4WsUhIKit5JC7gp7U0QDFWbMnXF2ESXZ8TvZireDijqz5xScr3s2TJ
mdt8r5YVodCRQK8aZOEIjh753p3euF3qEyQmHfv/Y2qbnQKkStxHXwjPdr+iRVOquDl0U0evu+UD
6szVWUYWE3MhP8qQb2nTnYTO6J2HG4tOfb8fpXMly188xYGLOABk7zGEhV5FViFl69w/ZikOVOmh
JRxi+cqu5ca+RSc5LSjctYrJqQe/2ISX2iPQtdqgFaTyhL+zepJqwS2RroKlhOKPeCtnexQS0qZh
RFwfpnXD9Md5OVxFMZLFcE8msN9x1lQ+DMILwNnDimFMN4XW/jlo1qMO9VHtdhFNLOh5vugX255d
TTvbP6mwOsQ5Y8M+Qk8FGDQLhMr3tDU7e+w8uRM+7Tdr2Z6MmedU/awEwLGjs9HAUOdDLFmUJHQU
NSJosYoG1zJfMPh73+7OpIDvW7/L+ZmchExTCB8K615eJKzlvUhszHxRHoKWoimKONEI4ZhDKoh9
r/Tw6raI5qRZh+JH/sxKMW8EskXgPgeFbvLUIB/Ge7hZ5D6gorFigw+vxEYCYzVThmqqNvfp9Kqv
bKgFzPf9dCWPc3wwJ24gosknbpPavJRultkhgqrXknnLPLNvri2ZExQixQopIm3/CaPnTGbPTaeR
0XOT4JVxxKIhgvQCsrJwOIMZexsd+taGEcjaCYEUWUQvX69JSPQIOJnytQe4aTZ6Pcg743vVvwZn
dF1ug9GSXKL9a6OS4YS9VA3E7qr735L0BSwvdOzWE870rjDR00IrS6LH2Zax4p4UKJYioGzNdYi4
Mdi4gVFZg6OEduAxHUy5pR59ucOy6KcIJ1JUDRs/TBgrPq/X+ZqpNNvup2nnYrabJlOH4fI6NVHc
JnVUuvZE8YbnnS+IUAhRI3wEPCpiLoxLK4vE1XmdNsdBQvQ1ZUaGcfJ2Di717sUkY+qBMu5xJdTm
e3qTKQGdsnNFDKFty0Zs0JrrM0IKdzbwhv67+9+l26PaIuXs0MQ+l4vpaFJuz6ZwXDeBCTAZwBUu
Ij+m5XQe/KhBVKRDcO4JTNT7vCeS8Pmm+dCk86+Ah8nXa6cxaj5UxklacxslJ6BhYPD8vSfSj+Qu
LQ2NY6CEIHTTjgRS+AXzFsuIy3Rf8CHTCSmxKa6ghzFbw2vHA3lz2nE+NEMKnu4ekPbIRkEjSrZH
a2+JBp7+zQLo+Clbz1D1x+bjnHHE3R1EV21axA4OdiJ1aKgXhsNjc62O9EUu8xE8oX0ZjaAM/YPy
lo1cs1BrA01DKAiqFKio+fnIxac953xXQRd7tf+3akRHhOYuG7xLQSvniNbNdQ2ynlaf3unNqG2i
wK0kOW5yfZA0MHRbtm3M+1ShM0cXbJvKKmfgSIqjg3KKA/88RFwqNNWrsXY5pbwuY8U3LnpgVD1t
aXm3BbPnda/6kFFho1mrqZTSI9tkQfxTF8mc/dU4+MnaRJgdCcEHkfZPyB6uDvH/PqE0PWbo6bNb
F/+jm7Kvh4URgwRVtmZshmA1xO1wNbuLEwvmhdgSlZLPZMaUPLSGVK6bzGERylKbhZ4A88cwAgct
u7j4aEWWlnn/Sbcwnk8Bmmnh6QEJ8c/ZfKj6L6dAgyce1ETQEBOXSOHsaeIYgHvNRq7i1ts+Bepe
tqM7qJUtMG31jYoyhykPvit2uZW4DVF7S7TBFb/RiRZ2jv0S4PaIXOD1BkmonY+8UcLSXkr7fgzf
Rl094+6y6T800Ypb1BrsVjZvcTW37jVy4cEDRDV9h/3Y+USb6XHtonI6I/9htmU8mBel2zPj50NW
SwKact2grJXDnjVOdhjIIqAixbvepj4ldt1EvkxHLFNMRtCSWnPSkZSsYQpOvmRFdBJRH3H+r0Sr
BzK8wWkXVu4QTZhmkijLWAlFsVMHdZJIUb19pcduc3Rb9Jwjv8oODhQf7ic2lPIkdDcaBZ9/JFEI
h5umCTv3dZOzTIEw3bb9KmsOk8guQgzbxLOWWd5ylB+OTZjZ92LurmsApZnvbWH5cQ8bIS5gv1Qz
VboiEJcIvA79FRTQ/e0ch8qQ7qFcbe5PNh/8wikbvRP7RWpneaaWGkSoVy2y4Osw4aiKMW6G27Gn
haYsz/PdBHqxQDRZMwtyvMq0MmqH+i6FF3aAI+cX3/AzHl+q6ebpcalBEydRdy3hRJGrXP1c2Yw2
r3RgQQeloBkAo1BeN6DBowj3lpmiguxzdn4D9QoXGQXULgT3tAl6xI/2jADEMqMheM51Cn+uzLuQ
EJYj0tOjTqy+odZpAKo76JRbbFvJ5yrrI2Et3uipVY9LWj1UCRcMfGX+Xye24fgMZmZ0N5wgrXLP
KRgeZdX6ccMm/bwVhf0uDWMUPpNZJ7YjuJBRKr0o8z2wmcmqRXLYkqNpccylpBs7Mjx1ud4ou3KJ
zakDenX/HUlwzf1+zx5Xd2JaPZZHZYlncB3b9HxDBpfPWR0zbU+2FQ/+JNvjnN+M3QyrBVNr3nsm
3INY+nBQn7yXwgSyNo/yeA3D+yrw+AGHGGAHPQgAjDpcoM0S4CJaKCbJuoLdWQEXrkTTV4vmVGdb
VXkP/Ifeh6+eub7IVXczioq56oO/HnfxLewLcBagyYROFaITVMIvX+g5nYBegnb26e2MGeMihCWA
1UKHU/IkATL7gRE1l967g8G4LCUZV219QL80cGjNHkk+WNQVPAE0ktPNFG5gD0Ppmb7dFPLYJfap
oDaZaVnTuWniRFbXx37Kbd2BGLMMv2mB1Ndh94a/cJ9xXtiKKcCREg07g31CjWhQJP/cvRrGITXN
7Fg67vJdXuvgAoc39G6MBWZ/bFzLREs9qLs4tB2UDjGXwCGVXaGRGz9CzETo+E+sSwvsD3GXirIH
Jo8tb1AbuPzpTC0Q0zWUWEPZnikkNox504hEhkXuTD+J5r9jSrjhygWnLbITy9AQFaMeCn3f+I5e
meNMFGHWBVj5kxa3IWPuHejjQbGuHS1CxvDebmDT9vVK/ukEtWSkYeiQU9dOacVLnMIZRKRmhQ4I
yx4pBvSN4+DKvpiaM/9HlebrnITzamvw2w9bkL+htEH8+5N9jgPvXxVsbOXlwr4Eeios6h1YbApU
Qmczm9gPBwFd6NaP7smdQhIQZXyMo18ozajfQBSKGYTeS/Ujc0JIN2iYIfgkhHFeo7X8pyg7hYwf
7WQWr3QeWBBwRPnnplXd1Rb+TqJ1uMtK7JuL7XL8a/ocF7A96r3p3Qd2L/mBPiUOY5S0HPRR/kUh
Obv46lgAbGyAPJ9vLojUB4okls0AC/xXROX4XCsilwlwe/YeRYOxbtaWVgv7hs2CNASQSeIPzpp+
gjLWPDe3j5nyLf5wl78y8MKvS9AxYIJx29lc/qlZGVbFGVOfHAkBF898YnHZU9f7s05mOJpJk6RG
qAvd/vgFtYo/S5zkCp7yHkZQYky9Zvmmd/hOsQqBWCm/gaPj54qD2gk08qlcXs98MAVaCZylJWeb
4QqfutwX1IWfIkE0/5zgV1VercZfSqlwTd4khi4j8AZIrjY5G5IVujTvszdb5HB7+hOW4C6wZ9Sh
AP49F+3OsAC1rpQS8jfwPx4Gb6ggRG5rA3lsOKxt9RXsD8fJ+n/MIhb05LA6cUSnshoMQ9k4DsK6
J1DLEX1n+uD5DJrfOPA/sb3eLsxyoG0puXEcH3xPmNpdAnEIotBQocBxL4Wh/xmwG0UeHw1n4Wjq
rxyRxfTk67wOjddQ19mGPQEjCFHHUAfQi7C7Ww5SODwdfwfoi/5v79Q4gWlVDqLJ1jSVkuURSm0P
zNdqk8KSnqEOWlM56bZUbiFNAXeGWfc9paZiae+vdyT6uzf4xPAePXPKzwblXg96GmzJbGdOu7LD
bGpc2WLojXAMrCiBVRkZbovjsd/b1TEfzQ2uNti5mHJzEEL2FUO41eDaj0s7NeElVX9Nj5H0weDI
qnr16iTqhk/AHasX20RnVKNdFRfFkIsbVgjOJDjw7vWVjDQD9em8HUbUl9qeHxHUdq2kouxl61Mh
8KYo9geAoaba+O6t0SKs/KcNS+9h/4aIdkf2kcijs3TzfALmIMcq6u5bBjDwDIgu2jES7Jserua5
Qt/huhVydtqSltau+fFeRCsSndmrQLmg1bj/HRPCkSB7jwrcfhIj3cdeRK+eHGQ4VA9NaBBPyI9h
YBVzLYshjDdy6g0R0w9I0PzoKC/RvHnwfo0zwLNUhBbCMxexcLvsrtHHglZQMVcW1It4p6cYBdZr
djPKeov80s5T3Ca1IUbAdV1U1mvIFnu/FPhzzJWiVWQoHxJ7shInv8Ii/+HHaHtZgqZePv1h477r
dN9aaQ1umzy3mg49wpkC+EUHv9byDS7+KH+XBGtsR9kP9Z+oKPEXkibQxlJatuTtbEdhRjQuvdgP
NjgnEPXHzp9YZqDV5EDF1ar6Qh0qqVRqda94nGYlxUvjkOHNoL7N/kLP+7GcI06TZTIN2chHfP8N
eswerSYUcGxVa/g62l5BaXr331HmqbxrLLj61QsLfInMtyDk/TQ8i2YcK1EaMtkDl1vSa5edo7TR
nodruPL7gWacZkPq+uMkOYULEfhjQ44Yb/p6VzJhJUiG5BUMxONd5Alcd7DlXdAs3ueLRBngHuap
WYkVIbf3HKtCTyKcV+F6TBaawY0ygc/7/W1GdURuJczLkKqM8ZhgFNQNH7EgDVIT4p5uuPe89u0j
05/MbIXNB5TCmncWTiy1uYp12KgHoAhX5ehqoFRioPgkoSdrfOSYEneXF5wK9TjyCseyyWgCC+hA
zjljAH8vQcjmISkW6idGRCQbafOsSASh9iXLvaO4sGYWvLLe9AS7Ry5GCIljPTRqVZKgeYoFDLg0
Y1z4Tegd+RfaqxKRgYamQ9jQX24WUvZXNKuPu3RhZoz1TYy06ZB3JNdrKSa0mmQ/TG527bb7kGO3
hvXYS3Y19Yt/oEChZY9npn96sA7jUNfiOSiRXxyHsbS+vgmshpXz3uVlYwv7kSX/haYfhKP6awmG
hvTRWispyyq+/2tr8kKKYGdzWU89N4eDOxpgfaONlUGA+iUtsVXivzku7kvFS1X9VSrvbttZgIzs
Bqe1lmi/eEdNb3roi89iyfcV+S+KPZe2a/id2znoMyNjKSMfxygsL1FbVB6Ygd1gYyIGS0AccicL
yoH2v8Z4ZJP77/OSogO2PyUPmcpw8M4EYhr7ZdFQFRW+87NDDVSuIF66oXZ6DXh/ogkD9p6Dn0Zb
yZmPs2rAprNy6jM+Z4zSWByjTiWa7xLjyPFWddsv/WaQJyEZtDbnDwFEw42p+DclYSrga28Qi6aO
2HuumYficPvXgqJV9KCD0BPvR7jetqrVxxCWrUHen9xtVYZ/89WSSIbIP9C2Sg6VSt+J9mxxzd3x
8CVNt/J83FCOaaU+giIpOkr/fZPBNFckuRqHWkIcE7KejUFLG45INarnXOBBkZz99spmUrkDTW4L
tS2DxIirR19GQg/oil4hkYTSEwzxDuO0A5Z6pA7wzxylZaHJ3lcB9sRywtnnuyJS+KtLPpjEQ7CH
iixg/2G/pCOfwi+uGaNmJtREOSQtUq9n98gxYA409eEj9WqLHNN+jtTGiAy20xsWhP35JBFOPh6n
gzMGOGVWMhEdVsyusBtsWIhxLRBIs7DgJr7MlHSyR0XBHlJdm7DVhvmT1pGFN2hhz8vgIwXocLIc
1wc+PR6hJgrg2mNqKcxIjTnnYjiG/c6l0fnjYLrjutdP/i3/eCGynZFnEkLfn9qEPt49lNeFy935
vmwa6neAVZSrK0/yNm0NTj/d3tWI7QkvNX0TAsEvD+0oXwNZrYbNPqrRKOvtzTG46VnIYzRHqPFc
ni2jLKkS3Xym+SZm8SXF/CKY2lFb/sceQFivagQj/d5Im2NL+OVChKfOU55MFUPxXwJvlSffPP9U
z49VcTkP2GV4k4WZ5rNJTYvjvhiX5atXAVfmlSDKMu/n17x/2yHG3QfF/ArVTw5+uB03RL8HA0M/
XydyrMgdkDp8WCSYFEwY7ktp5tZYgrtzNWxaP+hH15EUkfMWajY0UNzKl1Q+LJt35dSPNN1KIuCj
iftkFTicaE56HeVsEXQ0ODXtsRn6Kn60NdGuwq8sPmhpqvIhR9dL4hnQOFzgaWAB7ElFECEu1YWM
vgKnWgcT0zj80oRRNvJinB45PDHGBRzxtBFVj5l19OAZaS5LmmDxf6xlIBJkcs56EwjULwyx5CvD
G1oFlUIZjqevybI9EaBXeYUGB/UB6ni+yTWmR//bQ8pGwHwT9CjXNWZ1nszEh8GsqijFo/cwTPzL
juAQKU1Zgh12s/HYkrlLmzkcCckYMafsslvmneaY/fmRGuML/DD6RGvwJjO+BiCQFOLXKUoKDdSt
vL5LhUTRUHatL6AjnC7za3hCtYNpsmT6L6+YtPQh4TNDoFMPP/SyLVglWlMEj9GgzWEPxYi7Wuz5
azLQQ467wshJ4i1EpWyT+gHrr+NN6pUt2UDZfLJ86DVPWAutSOpwxTJkWbhC2FZiIgf+YUtJz2X/
6lswPPxNmkVLE3DEg7yXAvKmdigY6f3dowgC28pDVrZ0OxlwndYj097+HMcW3DO6Qprk+Z0aBcoJ
DOVESDMU2udz6Nop5JSf5aGZsGxRNX6K30/JD7RxtQ41LBCM5L2/peOaS1ssojlxwud5sCsp4+fs
mQPe5EyY+1HKoVktCAJNsDg7avu6gcJjp5XpHgSduvjMRtSOgqxLLUYb1hvYGCg6Ig0a1ptJw381
wGYbKrIchUUYFPjbKDens8lcUNsnB+C1CRMDBJHqBPFyKMArM533csAHAMJQK6u8OkvdJG0EOqrp
VHCEbYya4GZQek9AR1gPmARo+J4EyS5ia/i3nJBynmIB8MvOAXNUC2vMLplXerIHXHAvP6LF0/JB
ci/uSuPb4tXCr2aVE0HCkLXf/LSUWK9WtRuFRtWbr3PGqilenuKPP31MCeyR3xfElkrf3Vfr4ttp
FkNnfENL5j1FnULftYAaKAlZ+ksrXa2iMQpOqr0FZbcLTyNWJDgov/29yK4C3Lxnx1FxZK9IhXwc
ZCp9Q8Jx0fh0df3NUTN3eiGH4/VfJ6xQ0LlRDr4sDGtyDi05YKI8MFXtuHrRElvRr7dgqiSD+vik
w0OukpISHut5bUc2gQ/ynVug+RAjpVyCJ8BItHaqx8KSQ5lrPL0OsFlXbuoC3oOnGmoXtMKesJ0d
hlAwxNB+Z6gZGqX8Vlcgz/SPQXRtWxYEC4uVLZjBje0mPGR2syufCap0r1r1MA0sqLnSeBmKpjNc
ofbB70IRQqHQbTvpyYqtlHmrbilLW3t4s+ERo6blaLOX88N0bPHg8qz5x+C6lEbf8n+tzPx4452B
UPba/++HMBcNjfRcQDSrlmkCDssKx/hcvXwK5QrQ8lZY+8HbEF5La3Py2bUIiOmj3L3cQDNQ0v++
0vo3RA88OZUt4IFrDvP9lG2mS0SsUNclDSbwYCZqdaqrmZSOjYmNVAeHN4yueUdilECu3z98qliT
Y4G9xdnlYzAv2iMAnoHzONa/MWWfxyg3tKB3xKgt+/7FoDecoETsWntKv9TJCVcaCFOSahbYRiYH
FiVoRgwnve7FnoqFIqPov29eeVdhqVWj42n7HSpoexMloIJ8KBok0+gs5NBej7E7HD9NNRIM9oPB
/rd3KivDNV/YmhfMLdThUdsLAHsaipCmJ39MKmtrm63BNbZ4G4Da0ZC2W0AjrBdbpGuffPx+fcs/
cim21N7NV8b+QMO5On6DDfkmSVCuWzqBzPYOu5nmdvrstUvJYZ/+hkakJlJC1BLCuzS9N1rA73vh
N0kidbmuFh/3dyz6UAyF41UWlCfQvQVpU/rqWNL6fZbne2DL4CfyyYpgnUCdcKKe4cMWAUCJdtFr
SoqBcbgmjqYyJItOXZHi9xQT01Xw/hmA76+OSYSMcRLXkEZAPlBBAT58pXS0WoGK0djfCBfMRg2z
+pcJgmv+Xgt7m/udkhN3wRLpzlCCgYKOglvkpdJuZM5w0cE1sBnMtLsW/vrWerBhFcYICUD1QR0G
tc4MNnevI7gL/2C7KAawRV5H4c+q30xPil7nWE+EYy9CMf6G18kofw9+1XuoL48954uykD3uLWNn
I8izN3rnODr309pMe4h3r78duPnn7j4HpzyONytTUMX8S/akYxcwCOQ7iYYPyMPLZSSozsdYMrbJ
5zz/W8r4m1TbWhdKhUOI0koLbEcXILFMKWaeGVja2+RS4hZsl7FtVwXXX19kkttWzygeFgDclJiD
nSsLi9uwLkr65WfbWDyUaqLFdgIsF7F7diUf6jIYb7qEgu33uKbthJP+hIeDu7ECLaHY26diWiZu
KJaIAKshtzQgd4v8EEGceYlvz9WhAruB3gUjA6o37JNhLDrQ+7E8u/tVf2RYgEw2ZQq+U014M5aM
vJMnAUPAISsS/kKJpO/D/Qju3MQdTH1eJp2MY3ZXZ8tSd0GOTsOOweaf5aO26b/6I8DxJ7a4Xryc
NPGvhQ1IbI7Gjoxj5fWzQDFRB9RtG49rXQZR3ALVjXrYCMQZKmt6d4UMa+rgsxyLdeT8wQix78q+
hc8NhFttpFMj0ryQBSjgYYKfZc72Jp8sFoR116IsC8Ci7FFvReWGaJQXB8CUriB0wxd8qv524N94
m07EvtLKQfLbetQExLuqr5x1CNZ7UD4JCEVNjacfig9x5FXKXDtLeTDl6ogZmSGrdn5UPKUBCZTn
TNCrj3wzY/rXfFz5oRjpZlHB54bd7HDV/+YqExV3881OiEr0wIdl+eq4I5/8zqiMw/6hod1GDlim
gZ53Rc8Z+rZminwsTgw8PANMvEbaAePs7ivNBf4lyAt6UBi4uwAeX7klI+jdRVYgcsdJGKDeo1pt
Fe2gYjHp4S8PqgkuOvUTySJRMDpg4HtHkDVRGXLczEGh4VB7ny753LHpS2uiLKSMpvQHVF+12wv8
hMdZW33QwB6m98SLgIHs4kk90zcShgxqDHW43WKeKuHMwEYmiiQjN+hbG7R+crp6zt/m67/RUOqm
ZNiJsmTdapcQFWKiT+9JLzkKigwpDJoG+I+owUOsexD9Olf9rOIwsSc8vRI/NZZmUxDrjT10f06/
LYkjD4F8Wjm5Jb0Rh8PnKPz/U8LxEtYpzARDHbfaHYeOUcCO2wd1lUI7MOsl06pTd+V6jGLqgtal
hwxJQOEjg6qgqxB39aI8BxNCBvhbtcbG5GcoiUFyR9NjKG+nqHUkGGueoexKVKAmLE5qDoqrZ7M1
xVVYo/UONIkO2zCFtvwGYcPJKAAGdJ9I7azujBQfd9XIw83V37pro2Tcl/QGc1KbfFUdpNvKxTcX
v/0d+3eCiMzD+/PO+Ow+mWJY8cF6rCUe4/bIw4sQkZU83CrVSVxy4GhmfNWB1hIoZoFfamTtpQ9c
FQFIArP3lRn3yVS/17ybCxBV+rQgqfrlo8+1sV35N8fxLXyDLVyIm2vKfd9gGdiVqeFKREsnCe3d
xw+PDwtWH6Ccx7DyeSJeGq6Iw5nvjuz4MTuoDvANEaAZOD/ujeygiYqByvog7FPk2yHaS5Kf0OGZ
KK0XKGljAyh+vVGWyTKQdjac3KFVr+quk5AdAJYcxTezC0zMBpI9b7Iqjtt/fELaKAh8mSSUPac/
6CwMQD1ceGuUK9+Xp+Mby/s/EfkEJHJqXDbLn7/2eeFOI4E+1uuaV4gE15jTuoFk1TjS6KCwZL7o
EbC5AWslBnCePJOUJ8kQfMxb2Ma2YpfOwOUp1haEG2QNcU6s0Q/K/8O3tb86VNrZMmgY+ApqjzI5
vh4ITqsTN+dALpeY3nsN2siuK1vON8cXmdUBQ/Yt4aiVcqXneKXUIc1Qtk2xUyY7jEUEr2hUWiNy
d8+1jLv/AJ1s/Wyx2dvUifX3wQwnXhJJnLNm1/0LQgFcpDogHl6aEVQE72q8djkgKHdoi17dCdxQ
iloYTDbDjO0POZ0LhphCiuCmwhLXRBB/bAqaU/kBFFO1ZUVtOa2VMLyc9vSam5kCCYKx2MnC1RB9
9mkoRnXiF3Zf1wUH3HiaYGlGD3DXv9BS830I+WGpSmIFEBoArM3G9FXYrZ8/9osoTd/SAF4lGLUU
UrL6Nx4gzT9McEx/DvFoY+4gD4qycoZJVAhDH93T31kzxYSZ+PWWcNr+ErSqiM6/Ng83rlKsataa
G0uGHdFB3fRTRZGiyb3uKur607Tbh4FhBG3Md/4UPdDvg7dykkRJlUx4SmYTfkVYuwa06mQDDXyT
tuMs6W7MWDvAVkUeh7417hCde8LfD1ExuPm/xuThN3ED7SN5U7Xeck7cFHIrnj+H1yrfnTsXcSqe
tn/I/7ZgeAmm8KSE4+93zvA/V1W8MZAvf9lU1+OCpNiTk6rH6UT8NoHC4FwNFi6/904/8jwl4ycZ
ufFEtZg46I0OwDKjxv+ZV2hGU8v0FvPsAdFXw7wtmIMaKkEmmWKBIXo4Y2gSt9iejti80AhxZpAO
BJsYX3wzzLVnvM6cN2WWLou6eE8fzTdPtA8f/9ZKl1wBJZ3w8CEco2CO4fPCSZY9Xc5/y01QhfBz
4xy1QThwNjkVMETzvkPQLmFkM8MViw9x+pCvwhoCU78j/o8jcHuLsEfEAWunqtvh4yV0uMsPwwM+
nIiPxAqJPU2o4Z10n35UAJRTutyXyrekKO5IIgmMBZuH0xwqCY7YCWnPBLA2Qpsm8ZAEHrI5bltM
rCEl1MUOaG1cEwIQvaD6fldGNW5K/XOV040ZHonEMmhxdHEJJK34z0V1xO9zWdPtT3GUO+jzJ4eP
hJh5df+MU4TL8AaJmUuQVnOALqGT/L2eSrHOyzJQI2rblHNwCu66bOle/GvptVk28itdV/+JkUsk
28Kb1Fx7MKvFN5u9siYMmUzpxtYQIUMoInxRPHSjxFc2oTsVMTvr+nshifMBjCPDDkKuFUAZXcYS
vH8wUsojxUc+KfKcwIlDc5uXtFaAGP86RYGzfz26FDr0xCCecXaXeFLqwIb0GEL75n2zL4dM4r+n
Q23BMrPCwfOe273B2Q8Qz6iMJjV1qsWb/mUf7UWfOGSID5KrN4dlYJ1BUlk9aRBmrMNmlSO/ySDu
jcFa8G2lOIUh6FTssk9u+rHKVfkTsACPTJ+6Z++/b2lArSRPzTCjMtrr9O8CrkFmLiZ1EZhTtfdq
CIc+5hi5Yke6Xt9i9Z2Fcu55+nxWaf7wVPyGt/njbQNCVTBVsL6q4IRCVWm0jvB34cniwarJeHx/
iOxu+YQmbdCEKLffftm7zjvZL9L75df1K1yB0E7s30zRGIV0wsyZh4x/Kof8NFh+Q5wqscEo170n
EsAb6pSMCg3weAauCT1VDgOSJkvx/TU8zwZNrPcUA1dLETTqd4XSVpDKHEsYwRQNJw21sTF+YJpV
SsuL5d2jgvpecxMiP17Vbxc7TlzfTslZNuZK92ZYuUQi4nbXb6c1E7m4idFpjr7LsPrFuiDf/j//
uW46la71sDLVnpL3W/vgV4N2kWxPr0Ol3KAgyeayfd2gQKHvm4ro2QzyIC2YfWhB7MwpWHFMk3v5
8qlPYAzJEQs03yQLJxecax7drWeA0qzWv/HwNfXEgv1DHqUN6MPQ+Rf5gvPs+S6sVV9ifdzzBC66
4ASxND2tSWzJeqIcIXdnSSFXVu+C1NOGQK7fCAM9vIfaEIethFHt+uBmXOzTd8AsK+Oh1Xf/2gWm
hKVjxYmwSC+2n7ROJFd9aX5SDM6HiqmjFBPOjl59YAPMjS16uzwEGQGT1ZO7VjEMHYd4yWFbiSz+
nuPD5MA1JMAI27LONgm4ySXWkxL/m8D/6PVRg8J/zJfm+Pi45gDFx7o7p/MA8j/3IEUqkzCrsxha
aQN54+LEuyv0LcsXhcfCn9lrumZmKTu1Vkhvtfd1jUZLHvMJIdkO0lMRQ3zCXHTmfzXYrC0sYpDU
4zqb6hcqccoS6CnbskgL5eIn3aREWOcEjKytOEqcH57OetGDWYiBkDLoNyGIr4aWVIM3yQSstxEm
kKpeUfIJs8mmSJAiUfvCllMDRLkf5V5E3qbbqWx9CR3V0SHef6KQY+d6u9V+CCnV1KjHcxPTDShU
0SuxYyeAukwKNoY0C8UYKSbfqHm5KP8WV013JI6QuX91e59ogGiHlytYPe2MfNXUivtHFk7U+7WI
SpQR5StnYibswHh1x9e0r8dIH2Gimmff5A70o8DowjY9R1uOSyzzA3rd
`protect end_protected
