`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Vds3fYfVT3vmVmdeY8XKJ50w1p4S0LvPZsRzmB31BRMOdzNWQb3ocFuRH864m/QyDT/Tz/68hmeD
2wW8ef7mDg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
XV3c5pPgMoVk8UnK9dalQAhz4qy4xvQGSHc8VRfERmbCKAV7znQCmCs7Tsi/UozN5VqzL3AuVWSW
F5925WcXksrLLo5KSUbFxMA7z+t6e2XiVtdGrHtPEmzHbFlo+jwZUhnJRcXJIPLFBgoRC8JCtf2D
J0dCryGleyoYKWR11pw=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rSJmzkY1EW/eEBspr2ARhuXNq0qaJygX/yhD53vga8BFAAiPBrV00twDK5+C2uYpJCIUPIDGTiDX
cqH7mkMnjXJ5rnjba7szigev56e/4/EIMDeaer5IJgwAFTxIohtEdrBap/fgjtSlZTYeo6qH7LB9
CE5WBnDblYNkvWdxybAFIpvGnW4KzemcMK4jrs4n1JZNO7SgXawgPLapewUaQfDzcjsh+/RC+enZ
iAy/bDrOk1Gg6OfI5lApHgdj0KSgXswZk/hWIIuw5ITCV6xF4aTvpjNEopEGiTIgkyfMKv+E5+Bg
O31riS8u3g2rFv289LSJQIuiq6Wi9XEOoRafvw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
g6Awr3bIoKmNBpyopqupdpQjdZNVLkvau8WUEK5Hr0QHNtzwmXWei1Es0uZkMfRtE9JX9E0+HThB
4dYRSHcaodZO/nJGG0RIgI6JsM4W3P+mKCWOpkC8pEtJxMGZOBB+daNofO5BBjs12nVqiUCWXpN3
glBOq63JkrSsJ1tn9sI=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
IwoUPPRiKvF0uyTWb71LKSJT7cL5WzqDLUD1xz8tCXsVJVl0yqcTEIVryCusplS0aidUlp2Uem/7
+9ElnEViFm/KpuAMr+Nz7x+kDlOHPD8d7RB4tBqohkDMgzGCwLD4oFdxnUyBtGGXNmsPinFukPaO
zG3L5BAoDeV2QP7cm9CJo58o7q87vI6+vtRPYYOjcFzQHSr45tC57UiEMTyST9hL4GbanHOgt2eK
Jd1x15r5tZl9zRpGedBG7AQI6kJ/t0psvon8b3dy9v9KHPjh/nHMuR4TR8NkELD3hdnr7xjJOBhP
ieETCz+G2DLjAnvTfGgtIwZUJxM/crm15WMmNA==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
d6Egy6cv7pfi7JUnqoRdEky8pD21gigH7UkYJiv5Rp0Zfnd1ZSSzuQSsxsR8ZjwAFySetGwrLGwJ
1NqAvOHVMdJD8ZXDEvyjdUkmYkwJ4DMY/SOS9U8vyPZtGBIVtnbKAKv6YFRasliQ/hJoCkhkFg3x
oR92BoX8o+f8jfTrC4Iil0k6eWLDTya5YHs6DhqYOK2HxXtdAGe5OqaLmGJR4YG/E7n6pju2xu2K
+zWD2l7h68pDNHPzywwvGTraXm4t6abYjueeCjvwyDyHg/rc3gbCvso67/8a/OlTiSMuHjmrvdwC
WXb0uRD/mYxbG6/CwD0oB/bDbii7o831llt3Cw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5312)
`protect data_block
eGT2QLo62dMjhd1FHkcDUZ6BRjq7g4konhdhMPUkHT/DPxu4yvXngrYZ0KKKE1F33YRu9p59iZeD
3ZDdAIS6Y+jtov9HYEbvYZGl4ByI1W6p9BMOETZyyr1Meme44W4alSws9uPwKHcvG4MrEpi1cPv6
RDbJy+kCHN84yL6ZNuWVXcAE4Q/TZm2ea70Rt+rZiGmqzdLx9FeTfc1m3lKzqZ/ykaEzj9y729Gf
JRfilqkzLcU9W61az3LfvyJ0j7dBC3gPK2fQl4+xjWhBx8dAAlqN0kgSlFsaOhlqocdptq7q/2Sx
WBEA7Et8R4aU6aDKgUdeKSZcp9aVtcZXj3QMi/s2Gb/ch6Tb4+dt0aq//s1HXy5opNhv7PCXokzA
zF2ppp44k78xGVYcyd7H1WWZXck8HDu822VPNDT5/snrZSWBC621jwwDYCb2WcwqvbyeVefTg9VX
6t+aJVQ7KD1iD/BBM/UbBqFCRF+6qsc2h8NU8zbd1TvmBf319dvnCKR4nHPMhY3C7ss7VZzi8497
LOfNqxgBYN7l4qw7K2uRjZCkcHSiqst5UBPZFzc3mLKCPdJKrS2z08kh5ujGvHX9/hKLJUVFxWV6
Bf39f+3qxObLY053r5HO4FMWP2X/zoB2uvvTT5XiAWCV+w/WqXUV44ZyGmeN/mcwFh4vsywqMXrr
xP/S4Vp0+b3cF0sQvt+5oWdDcVvzQeDs/8lk8+5oraVJdMHLfU8AEvankJrOdyUQ0/d3ah5Lm2ED
veXW5t0TUFHJzMvc6BAIdDRrxh7bEqFN2ZfIP1Gu/+1x+Wv6DuxrbrU8bPDx2N6KkjVVBkiNHYr8
IFmtm03J4QvtjiDvduZ1SyoZ9RoE5deJ8+UXQLlSDKy3xJVKJsMI1HJwLsJN+2xDgM7O9qUYuUhE
qhH29oJqCPkzZT+GMPNxs00/viXXPc19V+laTy0eg44xhlXYQ0Xl/o5dAS/Fb5vFD0uGyuqpTpXa
TPFOijChgnYgut3vbXMWb3L3YxlUosUJ7hTonMW/FfzOeI/fRygUIsKZuuEp9jwgQUkAs4rh4kbS
oOj8nxxwjJSCsIuLd4OPKaseqKb8Fq3ZOQeZdoCUK/xTPMoQOeBouPNvtsV3LWS9n8f/sTCR1ETX
sq7qxAgizZQM0DRlhPt/gs9jitYqn/xtjedb+GveUNGmDTsrx/2iqkPLtFFszLbPoUuKh4En5TVp
NmGF5Dvf1HhDMxhuULmKcOJ6al5kiAraWBK7wRIYx+Wc/PLrIphEIyf+Pnh0KZKGRdmPkEDu6pyj
zL+SyVN/CNT7GwPvEaXqC14h5VX9LsluGNE2X9suc04vA0cDQFbbWN/5ykDsFm07nSMyPq+ZvjPS
HsO4DldBvrn5NcZ4t60Lq5zjfLyM2h1uF+BzGhtlhLN5dRrX/YcxJgXLl4yLB4KZB4ZfpH28RILz
FSRQH5FaeoUTrBzhDbWyuvukMsB5MDjMynrZ9oo1SEDTz2iUQukoD6vjMVgFhKVJZtBKNc/ketvi
/EW1xYRoEmAbHw+H43z3x0kdGv4n9B8R2D2SIfq5bf6b8B4LHCdg+fC14tEbUQO7bfqB/8cyGH0L
M22f0x0vNpIrB8xqtYP+rhSgQ2TNmGQIzgeWSaJemHFJ4sfwQLSFhkGxpehqiSnbYpd3hUmsvJ66
CCB/E3T4OeR8516wCtuHqXQhVwdzqAaiFucGmyFqIfYH4SH70hrxH4iPYGdciAjefeTriHnQiF9K
WACBBub6oKgcwrCXD/yw7oIvU2dWvUQMj7klhz32LyS5l1JnJkIViLoFTpvhMVuZ7rqunoG/ox47
0wNlddF0dEMjO+mvJQ2P2oWuuWOVzx+SI2YvA2d0cUEHvjiQRgn3964oAqd+x/hOv6OO8OdkQ2Qn
JE8AddARlCNCc+Fr3dPgwXxsVgTeOGzm2kv68pEhFryz6gOcLeX2gMxpoCcdcvJ50/zhOIvq6rsL
jsFkJLr53BW3+NO/Px3mtFVvUQofIMr90Au2Ctk5a4sN+szJw3fvaONdGnvIA6bNakhHFve81xvv
JgvFy6nS74AoxK1wSfkednUDvShnNMPrnUzz+drUTNFGnSck+hFrOePpCT97ObuAZXATRgQDrHRv
Z5GMVwpa2p3UKeJFM43/b+TUFpceI45LAcrq7jrxqxIaguqzEFYYTkSrcERF2YXY0uoGvCfw5Gof
yWOKOlJ80HvCXyMnZk+t7E/Ugh8Y6jAOFrKNT7tOz21bsomOc2gvI3NiXOn8sJ7D+MG4Sd37gLey
W57k1dfuaOn/9hcwZLTvM03QsicLiEaBosaoEFZX+28U6uzGO8CYE03DvdQ1nWuQZtu9TqTLBvmF
hwiuS9rZFkK+9pPjdoCwT2hdhQSIhKjk9CZXnWV+RdaHRj6rwWFuUzCEzVB8mYncBaIPZajC/a1/
ApylX/B6+cSSa8i4ZARjJEu9L2571K3KkngP02T4cStj202qZSWv3KwWM0nPG3ecIHc50CoAM8Xt
YiykOi7fP+GZMgvdGhow+Pg0h8H/khOkm9DdLqzJMDu5Rvug2dqWJsz/gdvvk6pRixn63ObjO63J
qiGSEhEx1z3ighz6Otpz6WKFfMioRoEmSUZAgmgIlEX7QCyX7hULpOFAUw2EiZFCLsovQ8NSVHNc
kJhywGZSQpv008qC0bJe+mhoxxv8DeUbja8pIAbZ2ugc17uKwxPN9NObipBFe429nQ8jIUAdUvkN
0Cz4K8i5BQ6Pyc1storNmhEFxpqUbnw+ztzQGR68DJpdt6yIfTrrQLv3zRdFHChpaVSkL66PRnyD
0UYYGKhfi6tsjTUIzkiYcOHALkpDBt+IHdT5MP3xTcAaA2ak/P8KCZLi+49anKTWEZmin/6ygw7l
O9ExlXYT6gRSjpEuhtlGDvyq5DRUCgFufP4CXFJ3irCg3nohhQYW7jCv+PKNDbaUL/2rIm3hOdUw
vglV3q061HPYuUL6bJY3KXfbuppGt1WMiZBo7ivijJoMaqUNzE4jrT1duBzYeqKl765voFJPCDu+
9GeAjWZwpiZ/U7rk9Jc/f/aZs3E/TAPvlGByfr0Xz6vYBG4VbtJcuad2edLpy4/UWdhCnfx6wSrX
I2CyUDa5zMjb87WNbM+bHilCiA3BJc86X+foa6hod0D8OGJS/WX/mXBECGo71UeQcMlpkEWpuBud
AI9YEZRrn9DAbpItPDFRkmdEfTtoTyjANCORZXJIXGShW8rXiW2yn7qge5O8aioKp2o6X8sj7oWx
N8KEm+cYlpHpR71be8BVFDcluQXYRoaGSVKdTVT9nXGK82Zq5dffK/J9Ja6EdgIhmLWFtJFVAYPV
nUAPPt1yBiIFptdbFZM0YcQNcO/O5bxdDSSi3FVG88XH0VjihDdb68HfG9GTMFet1gwUkv6Eu1K9
4ZUC0Q6JDrVUV+HxSmHzBN5CIhVZ0g02r8X815/0wzRcYSuDwVEioD9colN8VkZzkkFvlGKgRope
cH7lFAXp9aNXqXcjofVeBqkCcHadfTYfOaFAmPaop0rP6QynJsHr9YL/iDi6cpQTlvjjPkQilZsa
/uZvUpq/NIHpHfupmG9Fc8TaGvrC7SBbo+7NCb2uEFYGT/Ci163VHy/rJK/0DYEVzHSqjjyLvjDu
Ieho+g8O0Ieqlt7v1t20U1AqGh4wvMAwRNRLbP9SnjmqLugtXhtFPC7CB+rTbgHjtMCQ12qkkcFO
b2LVOLdLuFOndomU812BM4JKwWRFU4tJWOiamrP8G0Z5GAVynl5W5/YUYv63lAdSpTqZ4dQmMRG7
atGxRayWbqvq7R6mGnI6f0JNkz3UOZ/O8I+wPn4SN+sFbGJrxKjUB4HygykbjVxlIpYTJ5a8ehQf
MW+WwAj+KbzdwQULf17+5W/E3VZkA9RAyk6vGe270D5UVTfQ8F2qWzmQaCs2zDH3x+bgtg6l6IK+
VHpnHlBCm0nnJjc94j/BRXG90nSyNJBfJUtz+jKjGhDQYq9+Mm/BGOdjD3/8Vgm/CxkQOI3BkyXf
P4meRZJsf6toS29D6Kip60RST4aForoUxCn0KOvGs9M36B7H1HRc7uuzGy++RyW6u3rUYBzb9Gm/
s3XsopgKFWNDXj6NMAz0fVSNadui3B/lZkE+ZDiWrZWwf/S+w+VHUjxxdrc4x2vMvMGtgY211Qzk
UzK6hG8zvhF5BFY9L0XhKEkX4kbVxwrB5DsW34rrf6rTOQaF1mfDBoyZe6Ki+ei8hGPKsG4psBxi
QuZrGSqKybs4xxb/FzPHdKANXH7Jt38e85+Ify51fZaenPmt3QSmzJSw9bplDINXr5XvYA08FVk3
9PkgAqD2Ytcc8z5Jj0hPuTRKDPyBxR4KHpZi0xIaKzQRNQkK/5DezPdrfVpv+zJeSr4wl4mRTD19
UddWpnZVpdazO3ro6gAJDVK1jSCFBF60JiBHhqk1T1/ybfAF22gm1NoRWidv+OjjGopGsRRO0pbk
ewyZvY3sBR4OiJ/oZX3gP0pF65fqubC61HZU7hGFruE3S9ZczjrozZfXtiMzIyRa1zoQVVUqbeB/
bgzmUThuBG0uj8CNuY0kep8WjduGZE2oZTJRcLYAfQvb0jim1/1TMY8+qPQvJYpVF9IpRCVsVODE
j9/OXLzphC7WVRGVNnNeCSy9zHS8jUpze00lyHmrm0NkBo1zQ4oSA+zYhrBtGgICmdUvto56RqN+
jqyrgtseVPkk/xlsAWhxZg63zjxgTABrj9qSCD6xqle40eSNMxg4fpBM+XlWXNciImKbL23afCLS
6vsdi+qHc9FQGhWbj3d/2JO6JW2VgCi4dcCNYrrr6pveb2CvPHtpKFbNDdT6cZJ4xM2X+XvqB56n
amnSk0e8RqUtdaP0tOKb9xyjgYuQVdfUGbW/hbRWthrc+zvX0Zhm4Np8kqfkMQ++C1hNLQt4PLBO
2kaejttl+bKfOu9gr8CRkNxT8jnXFIUV+0/175atH6slIVm0Gkd5s9zEsFs7btlN5hg4GJZJyTV2
uRFmJ5AfxwrLL1QQKeZQkgGwacypq9Df74y0yEDtGVFGEIPDNoeQdIfYVFT78xDp4UiOU3RrGRHy
A6mhiRBXtprc6q92XYVyiiudLWpzzHxQxfPnkq52LwMaW6b+0ItwlpPOndd5fpAsz0kIvQBWxebM
AlMTZyoX+oWFsYGZF/tqHCG49fM9dPCnfQJu/Do+9/jML65OVXTm8nLD+ENrREaFA40NepfQGHn2
xkzRxm987qAviatw6kMYi0bNTtZTnMjjE4AxyQNr2qnxnVvESAYdmyIu1zjTc3v6HZ0tEN62lw6g
DLxfkmFJ5dzZDZwsJYUGZLEx+4qvB6y/aDkTMzXQN+0opyC2m6meKqOzL919cu9OMvl9BCk8Rjyu
Y4vY3SjZiLQBlo3iGG0GACNZ5owogzhiPgSkebAeUwo9ueFLzmG0raMkFs7kzt3Jh+LMta89z6gM
FjRQHOIXPmhh9OaIWwZIkyqorGvaxNgp/U4YHQH42fp5kJ7rO22r+5p/knh4gk4k+fVoEjdF0Icw
whOJ+WLecKuAnSXdqtoJwkaPxG9yfsN2Zk3N6Yr760vwxeesuM1eNoeh/97CoK/JzEICiqv2bmtj
roMB4QOXumcBkd0K7vb+/UmXT6oic6JHmkpzuiapBWvBE3vP5cUm6ta3Dk5l21kLl7EmduHJlhVN
Qt7mPJUgEOHRKufFcrM2kITvtNqUFhwDpMChJRZsqwoF0Pbq9eftClGTLHkWsgJMvX5lIzSwu0tG
RxNG+WBb4ItIFu0P//BNs75YciNzyC/B0+W7x//FC7m7aym3ykkSzb7IRXDUESJcRSFldB65OCwk
3GXomxDwrIp8yI0ZUGEqUgXVxCR46G6KWCCR4N5COwe2SLzVZydJiJZXcAJ0Q15T3HbQ5L2v6ZSs
idFFY/Afe/gd6Tv6cXsdlqZz8k+BSD/FCUGJWqa1W5VrUPkGtX62Kbd9X0LQFb5vfpjUTDB3envF
6q38zuOt4PPDlm8WrgAKD1phGkGDacJtA48vJs7FYyaY1nslBcdrTcWl06DD1Bq479Hw3Lmnz6Xn
oLmER63ePf4XF1FeOah3GbnU0jNHOTcVL5zwCkKUSRmhHT6eaEglKQiLxFo2up7L8V03m/0xOuci
fDPi+uxaooWHQMBSVFTXBcAPCwp8svad8IgMC1KUr3caQULLUV+ALfUI4MGabGD18ZjsSk9PopcP
mc6iDG5Di4f8i/DE4w+jQhqJWFjHJ4B9kzj3Z0R8Ng73/vIgs97rtmOcl873PoCn5CEm01mKZvM8
CFTXo3wGaev/HnYLId0fcvC06kVUmld01UWdhiDeBLiqVZdGfD2YxfER02ujxT2Uq2na0h3r4WxR
B6pRTGn1oH2wmV38gMvic6TQJl9xJrzYEEIUnnVAcRNC8iEMI/CwrFkt55NMpdJxqGcXKGCHBqUh
eSi1ToNl0liTQ7J+QAizBIdQwhqEqj9uqqK4hZSwYWlTxMJeg8wDetQKkEUgdGEQAvcW28vBSQna
DacfILRvcM9zmh3oUjRDo8KNphQuXVjcU0kgMabHu6o8KqaDtRfzZoppWa5j1+Hi8Pu2IXLXS2K3
ObfDUsNMqJX4uqOg0pkg1baOS9/sKpeQ1eToCUG0RcP/nC5yPrB6Ogd+gJY/icRKytbv1ugY1ZvU
bqyBrhmkhkx1A95AC/csCpFN4bXTp/hfAgsFmudTIZY+FIgNAFdmLTPULgt0suge+GmdQdWQv7FK
tJDhhxYvfL2CDA4dRew8JQN6oszc949VqpkNr4pKRWK4F9wytOJW1LqBxBfWfADkwW248jhmWp9v
KXzDpdTMQ6i3lH65FfCvSStKs5nWyUQrpDfnhhPqpglHkdpuolOOeoc81O1z9GXce279HLb0gHnu
iz9Zrkxl30KhvVp2hRrR5ZJT0Bb6Eizd5i6fQO4lbek28mscB+qYCyHpu+k5HNyBCYRl4D/8HTqi
XJmiHUflq+fhNqkjK0L7hLd9EtbHCDLU4YY6WVSmCa9b2sR1Sp+3ysNKTNCVu60HZTkmsVDdBjF3
b2LMxFwPI+1Viqs=
`protect end_protected
