`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Vds3fYfVT3vmVmdeY8XKJ50w1p4S0LvPZsRzmB31BRMOdzNWQb3ocFuRH864m/QyDT/Tz/68hmeD
2wW8ef7mDg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
XV3c5pPgMoVk8UnK9dalQAhz4qy4xvQGSHc8VRfERmbCKAV7znQCmCs7Tsi/UozN5VqzL3AuVWSW
F5925WcXksrLLo5KSUbFxMA7z+t6e2XiVtdGrHtPEmzHbFlo+jwZUhnJRcXJIPLFBgoRC8JCtf2D
J0dCryGleyoYKWR11pw=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rSJmzkY1EW/eEBspr2ARhuXNq0qaJygX/yhD53vga8BFAAiPBrV00twDK5+C2uYpJCIUPIDGTiDX
cqH7mkMnjXJ5rnjba7szigev56e/4/EIMDeaer5IJgwAFTxIohtEdrBap/fgjtSlZTYeo6qH7LB9
CE5WBnDblYNkvWdxybAFIpvGnW4KzemcMK4jrs4n1JZNO7SgXawgPLapewUaQfDzcjsh+/RC+enZ
iAy/bDrOk1Gg6OfI5lApHgdj0KSgXswZk/hWIIuw5ITCV6xF4aTvpjNEopEGiTIgkyfMKv+E5+Bg
O31riS8u3g2rFv289LSJQIuiq6Wi9XEOoRafvw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
g6Awr3bIoKmNBpyopqupdpQjdZNVLkvau8WUEK5Hr0QHNtzwmXWei1Es0uZkMfRtE9JX9E0+HThB
4dYRSHcaodZO/nJGG0RIgI6JsM4W3P+mKCWOpkC8pEtJxMGZOBB+daNofO5BBjs12nVqiUCWXpN3
glBOq63JkrSsJ1tn9sI=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
IwoUPPRiKvF0uyTWb71LKSJT7cL5WzqDLUD1xz8tCXsVJVl0yqcTEIVryCusplS0aidUlp2Uem/7
+9ElnEViFm/KpuAMr+Nz7x+kDlOHPD8d7RB4tBqohkDMgzGCwLD4oFdxnUyBtGGXNmsPinFukPaO
zG3L5BAoDeV2QP7cm9CJo58o7q87vI6+vtRPYYOjcFzQHSr45tC57UiEMTyST9hL4GbanHOgt2eK
Jd1x15r5tZl9zRpGedBG7AQI6kJ/t0psvon8b3dy9v9KHPjh/nHMuR4TR8NkELD3hdnr7xjJOBhP
ieETCz+G2DLjAnvTfGgtIwZUJxM/crm15WMmNA==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
d6Egy6cv7pfi7JUnqoRdEky8pD21gigH7UkYJiv5Rp0Zfnd1ZSSzuQSsxsR8ZjwAFySetGwrLGwJ
1NqAvOHVMdJD8ZXDEvyjdUkmYkwJ4DMY/SOS9U8vyPZtGBIVtnbKAKv6YFRasliQ/hJoCkhkFg3x
oR92BoX8o+f8jfTrC4Iil0k6eWLDTya5YHs6DhqYOK2HxXtdAGe5OqaLmGJR4YG/E7n6pju2xu2K
+zWD2l7h68pDNHPzywwvGTraXm4t6abYjueeCjvwyDyHg/rc3gbCvso67/8a/OlTiSMuHjmrvdwC
WXb0uRD/mYxbG6/CwD0oB/bDbii7o831llt3Cw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 961872)
`protect data_block
eGT2QLo62dMjhd1FHkcDUb/Rddzk1VBs10dc8tVL9CLGSchM4iifQyZg5lTZwaYPIcIKiBVD78G/
W1LE4GHMGp1tvw/C6GIqdWDRYl/w8O9LVFi1G1ogzsJ0c1E+7r+0zsUmf9JjRmDxoOowh8y4JtFS
BevKFe9MsZnTkAkESC1kZJzaUsIVTGvvsso59iYrtAfxLpzpe12SiHfWycfkFqpAq7gjKNC2tjCf
dZLD332MNtR2WEBrUXwns70LjnvepdLj8ZMPMN/lMbUg5fevBcBkTz5OzBH3+KDkw1hS4ZUBbhzM
KyVzZHSYZpFhzei6UUheXielPx8wh++Wf+sy1/CcMYwT6Uuj7EaBibb671gXKBlfx2UkFXarDCpm
GigJ4EPNSTA/g8gfe+1feKCCaErkRVQmNYQ15dCEdckqMHUBieGJwhDODZ3wlqIgF/jQL4GRbxF9
EPgkgYQnQoE1cMMk7M4aaq4klvNj/w+t3TeRceZvvaFa/mAg1p9Uo0xBqVOWIWxQqS3dhv2aBFQo
JrJi/WuyacSp4Rka7ZNTF46Q1Dx0JZu0MSuMwQaZFEfGxfxKJhgYCXBk1oV0pkhyFs2HJgP4mWbH
3D8VymJo8Q/QaY0l7O2MSuQc8W3uHMLkndpqoZ7317BxOnvOLYtlA2pDIqCwVjf4DYGFSVRFJDD0
joOJkHRyiAiUmnNalO2Bl0q4HlZeqsrZPgrGN7HOw1ppzmZNEA2UN5+FZCFur3ZRYcYz82/bRTBS
MDFo5CGUDmvRiOJUrNvJ9dFNphSXvfJMijXM41m5cXUAt2bBp6Pgl8VyouwtFWUy5NdzT6Ck75wn
dNO/3LLp4GEJgo6aTitCY9cKvWiYiiMIeHm99bxRMJsih1B9mvVeYBz4h7aylUY+p6OmOgJGueT8
XlnWZeA4LZvx39kCIg4RKlSALdtr8c38WeESt/8kisd4/nzOzWAIQo1vhLw8kiVkt63JuaS2EOv9
AIcY++9IQe8l9v37brCAf0v3jKI05twkpSXJN7VxQ+z4LmY51j2XXWyINcD9CvUTlomiBeo0ti8F
njcx9QnHzZx07DbgKw9Gl2ysEzn7jWDfxwNw5y6AF1vIAT8g98IF5GnYrYJZYKzsjDwu6pc8ThFc
oVGHSLrjtapr6plkRuZfTnY3SnV0XNTL25GCVzSaVPmVhctzP2geeblcMK82imfKELL5q67flGzA
TE/B7q3IBtbb/ci7hiheU+r4kTNqB4GOu14/o+r6vWReV43zpv7pnoUOfBwt94+/kj+33KrQYOm8
pF2MJsYzOpidDUZqfjgeN/5VvW8MmyoNzNNIBzEYkGdSzxRyWZrRhmSpAZYxvFI8feBPIgnK5VDc
w78+iLpBIlXMmz+ZkzC4eSKgA0f7F+XQzKPb4z6wr5OUPTcGJ/A0GriUt33bQF2lEqUAxkAuHbvN
8mLKEbbZWB971bjcx6Os9z1FTciMLjRcPvvO3/t8Qm7t1BbbfAJ+6ak821uTUXtNnSqlr/ikPuRo
nOR+qQDbfsObMpc6gT8xXO4CkH+l6e1wfBiQ/+r/XPZ6oRqxrHegj/UAzrQwQGYWG1Jtd9qFIsS6
o5uMLAw1yCuVE9XpFGBCLkBaQ9yBEl892StkDQLb/ylz9ttQ+eyywCtkL4ItlYTxm7412EGg5aOv
13gQFh3YF41RjWQZmXfJavReDuUbb9qxzLTK1afaR58+T6lO/qLGCEItC8Z6MLb9MmhrmhenOetB
iqHNNAmVfKi56ARZKMlyY0l+AtAAS7VhvA2y7agM1z02rPVxftVXWnFPzykRh3UrsGOpDSvnuKzc
Nvo5GhIj2ayPsYxdzJvsQfLn7vxFfs2TfJVXAgvMoQySHLWLD+v/kmUgS9cZEt/S25ZpNEmBjS2g
eVYCC0Vs9o2wAxHyFF+WjgrjxjqC5k5Bw11tJ6B3b182jd1XR/qcbK8iB9z3g9fC6G+4AOC5Gpmh
WzZkorldarHEZxXq2rUc0OKGZW4CdGc86lHZ/RrGvSAomzxz4Y1TuZOiC0BZFIbLGFefDxwVwPWW
7396V98nNbrapIUF21J3RD2dpwfHtrh2EaHp2ZVyu7O724VWL2Zt1YAK/Qr2CyA49xotNYcy4gfG
wOPXuxazv05OOJEMthyaYjmMGzPEVCMckiXsPe7uZ0zWJrOS96wGqExOPzJPY2lfLxwPDZdEib/s
qdWnazxKNqg0X4S9oShmxE8dGH9JH5JTZxfBXqR0sX13WupVwhZO9RVO09zJ7U2cAxioo3zMMEsU
/wP/VDoNPUmgDdE4JKQFsy4WzDkA9RvH+cAJVXsqwJ3GD01YRB2ScwQLSKiuAsA/yyQW7IHaLm6Q
okNGUOSP0vjX08HpGOUi9yaIiMtm+2EADJmP7OFHMO2tKwuaWk7fF4d57wheibeJVuNGjfWYo0bQ
TENh0Gjgja6u3QDwrcbuuvjF0ItTO1p1cZ+4wAMr2wDb7gp3gcEG39aiBxDI5WgYfacNmFu/L4fM
aL23RI8G2V+BswXEIMEberxKVgDGgWMM0Nwdi8lBn4Lwv8ViayXrMmnCdTR+QUTLlkPtvf0D7cWa
/JhfpDtyiIMypZ2W4diqdhm6L8FkRs47AOCTwSoKBzBZi7KXn650Uoqi2jSxa0tEUqSr7cLQ1LVR
vB1gYqUD/TVXgacQ8lSZ4cicKKZKx9JbQUYfO5Eksr1QOpbZID6WirAofsAFneIwz+R5fqnaO2SG
+PcACh2e0ejVWErcunLxq+68MPfhhBn3iF+qXYHcPGUhVPVBrDwCvqUbZxUjlZ9BedpWi48nghgK
4wp9+k3pe9F48OFCDts+rQnCtyM2Ckqn6Pv78rS8YhEXfVbzPLTkfWixiXkryqhIysHsGN1x7Cj7
GOQqve4fJnvZLqN1B3t7sJ28dUmc/6IqE5KafouA5rJoEJeiI9AjmsTJrPLODf4I+v4kCZLAkmlL
T43FlTylKdXdMd/R5YGyCWTVaI3InlwV5e/k5RbeBxr/41LI310I0rFQb7S1rIx04D4AZvhdc0bz
RNV5H12mZLnug3qU2uqWGzKijX1h41RCG0R6I7pvhNkIioHgTEDrrU4lcAiCtjkncQBFl1eVby6f
oj0VGRTSW8aJMOD/6m96RIEMiJZnSUsD9wA8TMpiZwWxDoS0i7Krg6j9LjZ2tixqn9E/hyatKoPI
xkpP7rHznE2e/VuF4t8VkNqQAGOqKnsOZM4QAcgAD/LbDeZq6w49b/J741GF3ZI1QSqhxH2HOAu3
BT5R2//sQtph4XK9bYkJqi3oHxApFz91lGmTfGhH/VN9OfPi+pqT6+TPC7iZ/xZt4wZGUQGEXDIP
Gb/+G5NmCnuK62RZ0g/jXj3lDdyvliv1WqPUJmQMm6mEypLe16fOVxep+ArP2/eyUGsXFSon1Bl0
Kz8Jc6+hpVis/36tIU2LdJr8tzvjPISZz9FkoT+zeGfjGE6qXVqhg07pDjJWUiLoo5ziQvAsI0DJ
zH6njyH99qtyvf4uwcrs4eg29mmKARQTO+UOri6E0rClHLdegAx9wmeM9XgeltV6oBx48Puu1OCo
CksVyIDztEzJOjBKEAFsLrbyI26ZV8LnpsOT7c1joSi/Oh717Ztr7d7P8RpdwYWUce8qPGcXFykt
fETFbhpF2KL8EYRq0V43sm4bR+/E4GoHpMv7JpmZzkrfVQn4l5NRkeeJa32eWwoEJLRIjzTniy4M
Z4KYrKhyGDGCfKA3ZnK0Dh9kt56+GNR11eunyb6ZGOSv3GJLflCmfKTPoI6HxuG7RIQjlW+bfm6k
3YAKnADpgEP7BJ+UtkmhgcMHoKK7M9V5ng6rC8oc51X3LRzcTYomAdax7iaWk/qeTw8K77L1U4t5
srGdLzcAsXcXdJE0UstLXbPrQ/xINE4xBAsoYO1+DJYaZsXqkEsZTrl3i9huZV9NCvhvYi5+M/uX
ZdO0JE6HkAPxsM+vsTUgCq6ViaQgRQVMpLRkml+ANQNqb8DFniCdvLIKAxb6haAFJxj6gjSJHoxG
j3KfgZb/ikDhAIvDM3FirbKxqTh6w6hhXLGJpbaeqUFu5zXVEEChdQ2GZeEQ5DWZCgssu/wkZlyy
1XM+4GOvgVZl7ZRHpsc6Ui9GD5w1SvUNQutC6q5krFz+hUWUyWh156/DacKQcAH7nq3c0Xb1fdog
jz/Rm2iMlfcOG+MmxdnDWJUqGXLYAp2x2QrRLl7m5P0nWhHtw4KJNMuvwgFVGtxHz6XymIIh4hqJ
vaw3wPkwPb2rY2oh6FeP1JZgqDbZtL9NhiGVcHI03/ti8WHY92fsE5UYj12tzNJjVEZKFA17J7lx
AlXMhFcxqvDgtMODqBBb/hRtaFVQ4mkj1hbqlIDFsdLHAub9o0ArEVAPQWp5Fas4vF49H+Cfsgaa
NjWPisDuAAxuXMTTuLwTJU0d69fFnZ2cTRtxWRxcm1mY43NPzyvhM2p4Ocdd8IuNNxpMpbhm+zRG
D674ITnxja7kIlVN3OG18UMouoxbDpis3noVfcXUPthLH6BkExXhnXrxdTfqXd516D8EPWM6P/RF
zS03C0/SAWzv4+RteJkWB0P/rzc8IYjMiNBFV/2L3J6FHYmotTMpI5Mw7CAxGlvG5HParktW3RdE
FRpQ+Cu2tgnnugbD2XztN2dqrTTVokuF0XzPsg3EEF8R9OqD3TFUdLmo1yORAkKX9+4VB1++4L1D
U3p4w9/Zck0/Jq21pbURHnsDxPzMoYHxED/RQtc0RHreDX2bc5HpOdOFXCkEtXS1LDennWLZjZEi
85wNcBVH+V3wLiCdyGLsmQFWzsFczEdjm63HZOuJqRVPSVF6r5iZu0su9WDeeVsXNDI/hxWy70Fn
MSJtvauRij/YSbqefeqc7pq1lMwc2PA6+fSzm8+qkeuRUr4PmB1n8mdqJmN0gOIQ/Gy+xUkm5Evn
lTb6R6jm/WqvS1hJftQB1SOvLM6VHlOzVl0n3KwDC4MwTxxVn9evaa/TFj9cZYEEVSAme7sH+HcU
eEmOXW6TanBheP83L9ylz2MM/jG+XDoCuoj88gDtNyK8n7PKT5dSLCNZk0HwQtjmnML6btxUT24n
X4Q/yGOeBjg6Dl/VH2JzyXfbgrSG30FpBprLyPcDxhyfyX8K1alfeoQmYUVhRRgua56cqBt5lGvf
SIiGhoAmHOPlHNvBWCu8lUKTAC+0BCc1Fb+tBDv5cKmqTmzM3bm+gh4wOy+dhGZDrVtw/thorKSv
Wa5ri3F5vBmvJWorECrRVSN0BPdpnLi8NcXo4VqeyxJQoHOVrJgL7Xlz1yo9lcMaDn8ejmIm/DiR
zsJ9UHMmZsnkztmlHoM+MpxSiLVcSNKkmlt/A5k2+LaGRQW4NXNvR7+4HfM05jWNh7pvnbDrRQFk
2R6vmXsU2l5kDXyhrxYbtIgPr7GZeSz6mHm5uGgtnhy8QlevqRpRBD9cCI1qTGWRdH73JJnRFlXE
dSWy4c9ashacvAwDX0Gr4J/BK+U1bI5N0psDetQmrxdMcQac+Wq4Z0PbJlkpmwsmEbIqNsaRbxAM
aRuWNazdyfxvXO4TybqThDm8Uk34SSB8n4yCDeh5YeVuPK7yOjwu2P4NMhZl70FbyzWvmQlKJfbP
bnplCXNeVeU2ENxmuo/VQQULQrgrQAAGP/OhhWsumXN5D+2KYaKmKqJdH6Pqe+B4g37nHq2xc6NW
+36O6FPeD32dSoRcLrw4LweNpqdfcrDZI5tPYDg104XL5L/COs7vvx3oKo8a5qhnf+6puF1sFB2H
nC17QJJ8Gj1twZ/eBqJFK0gbOPXHjC0ofqoqgdxr3+qFuUxGH2Rr52dw/qPi4niwOx9iKw7000uD
KdoaDQ/o6AyuuojS92ofzo6HCK8uWqnZaQ9bsk6poRSjsBVRjdsPXNT3ULoofpGfwcvCz9hUhI6n
h0vgaupALU5b9N2bHNQHovzVgoJU4EowBMZGgNMpNn8ad4057hntzzsiy5p4FxS9pvxFN7r6VC82
Jf5+3bqZ2q8UMSRWDBu3ZyHQ9quF7lQlXTVHhhX6iTuld19S+oMYlPEd14QodHEg76hfno3CnVCX
Y7Zaq2K991OpHl7v7CIdiB1+oobaDZYyW4FYR9tUeNktHV9jLNaCClh/+vzyfZWpCVoy1n3XI5aP
v/ksy6Hc5UzK2E2YwPJvc9ZMeMWI4ILNUWnRiIX8ReamzAAzcOdIdTqyd12LdV6wuY3CfBGecFES
QSKb9lqHBcDv911/luGHHSo+ltnydtHn1KvMsnGJGkJRw5W0Sw8s427lpuwOJgIGO+tPRBEwBs+t
bQeYEPAzi6sIzTRL1DT9xxk7rVfhDvRViBd45MAw6M5ULII9U1fCWrI8milJr38HpUajvot3qmNa
YI2R05JmjbyCts0Fl8Xg5Bzt3Rbg1fnfK1/HPG5+pnRFpbenn54wKwjrQUUIads8Y/Jid9Cd7Wzr
5M+mduvounBY0YcGqUC/Fo5QH7+JJzP3OWQsMzSF56aBLIDopzAXO3HfDIgNyw3gMcMMrVlNgy0J
KkuLU7/KnL3eAhwAiQPCuu5DexVc3AbQyY+VvveJKqtT0WOmho9WPHC+N5tjKAHaKTdMuu6KExbW
KST7y8xwnBQq+Lc3t0Huc8QzfxMzQkqncjKsvBvlqqTZJC9GcEdn1JBv0pmm1jp0EFJU0fvGpiFO
uG+I0mJ463tKHIZ0ojtqJ6k6V/yu4qVSeuIjAE+7Ts+z9COBauLvzN4Qu0HYBz2DAonFbvys9TjY
o49h7wHjOUR8YOmGjLH1OC5BIyEt4iywun3xoxUg9gAAcSwHsF1sqeq4hTv/KtIPpmlnQI/b6DSm
ycKtoHyFHIn7eeXlWg/Mj1Aann68Q3GWj+qfTLrBF68sxvvtvw+1otJCNt6upaQ/2wPpBHblG9pv
8yBP6wO8o37glWWfExYQz9e9LhBzsR3J7ciLFyKtNmSCWSmu9/O8kWuw3AE9WXIfFKswVOV2CBcz
mjcI7JaqPnig4Ey+TvMFWuzODRNHtbZlHIEma0S1jM2rlfLzUR2TczG2oT67hivdUjUrA9tiCjRv
vX2XHAEraMYSGC2f7FM86DHlTdC/2LSYtayfkupCzUuobPhIyW4kVxTbItcO0ENzh01CYHvEcInF
2TpBepOtSGuVNRsDVIwbDl0RY5CE4p2YDFywsmr0CBK0QHru+59Gp2H3pFiqUp4gQN+czYjZL/sW
2nAGM/uDo1duPM6PMUuo8AX19vpNuDBuk9BdUzXHojN0fNysPwL8JT6z8Qzfsn9rSSSRuXieZm5I
HnzyfC9jZvtuywDjvYWtEKeX55QR9MjN9KddhZughXt/jydyHHi14BwEsbj66+w5r2Z8XEnTMl0C
MyOfy9hHNcPyPcLqxmLf5e3Fp+NDcmwn1GTHxyAQCn9r3GaNGFIXiwEBSZ6Olc3V61m9i6ZvX3OX
WiD2CffbscnTCVk6xdKuT7F3uNhJ38qKNNtjiK/tDZ+6ekZYNuwxR6t7qMRkl8fjsQFAgFETmnkB
FlDlvxggl7yNWeOUz1RGxNklVb4c27buiuZOFmcI8mEB9okwBvrxgEnMrxrgtbzZpFVI3LwH5zXN
Oy3v060USYchQdyuCedIcJKlKQbTwIMyHOACs1lDMWidTHuvHs8W4t6j/xGutcxQUPzpJz2lLSMa
yuw3BruJQ92eS0Xb8eLswuragnnAhULFqTvd9Du8SqPN9rEL5HRA54zPo5m4Mf23slW5Yizrqgok
V/RCiLRKm+iaUCijnaabXIsYpwsv0H7Ilv5kcqj9LIARZb6He6UQ9TS2S3r4ysM2YolGksZKMEzR
kIPbtybA/hRFJ9r0MVjmMHDGfh+tGVeVJ/jsUUlCTlEjzV74DNV6q24NEGM7v4T+yjscX0Zg/Rgk
Cti5UnPkydJx4Sg250+/jmtlbnoHVTM0dvdEJQJl5M3sHWejH9Pabn+K9qhZdHAS80522tQgqjSU
ufqkMX0LbqL7JwNsogOZmQpQ74d7HYjr73cY7T+qv/b8tv+B5eBlgCff7I3FspD11sRSRT5mKyqm
/iyqmGMwnME3kqmwsgdgPEXTykVm7bDwX3fleJg31mFs15PdFBr6KvMTSHzxAnZrkneaO7oCceSu
hXj5yOQmpWawhWC0rEqUfamaxuRoPWCZAeuo6f1nowoJpkh5hBD0oDnptJx5I9y+fdtK5ShRJBhv
MV+fPVxyyJgxoA45MRYcnF1EMl8HEwbzjXpBRu/EjphJVzeWT/wqmkKITME4kLifWOFIRqXWyVfW
CONYfYtMXno2ZeuvN9dw3IqFAJN/0aTinSTsaVxH1Dusqr/ScmOs8JcUrYupgzUWb6PYoTJW/z3e
SldW5Ch4B6GgEf/Gje/lHdyvWdP8L+csHqUw0RMxvPUyiI0E+fozWtoKf+r03lKKoDJSnrf4mznP
vkX2LRQ/sNUbaCfk2cexzM0mF49Tc/mnDA2Dx42oYTD51MoGAF40iZHtEVMiov7x/mQ6kjLaCcpu
DyYhzWEaJaNLhyQLCpRM/Ma4kE9O3SJvbZ6nab/G5XtsslF+b19KaSW3bOfMglNHQ/zVccw3PgsR
ka3JMQwG8vqwZMKugVvBo57uBQTJ8/p1Jwaeib+yMbX3LwJPuxWKddner6VEK8yTP6GQOugE6lnQ
x1z4jJgHLpUM73+zvAP662tUJqAjjhubXoM1/uBVWI3Fxp9emm4+npPSqpAmIWXHBLmfxJDGSIyu
KG6kfruz3upZrF4SewdXCRshJorBlCYvwM+QjDvbcb1EEJ3733eO21UVNH26jtCbTrVrBXYJfriD
XrC4wrrGzpLJnRsbU/3fZYMC9rD6c2LWLLfL3exlfvKTx1L7kPoo6jZE4nZTxn+bmZYGzL4Qm7Rm
HxGhoIltSW7uybiowGqR5SBgYluDI8qwkgI63oU8+hVifijfxSqar0QhmtQKupEYJiH1JCLC6nVY
kgfqLyDF3xtLXrl9CMLkaDc3oJPfIje1Gx3O8uPj0Xot1w2dhd3+fkMUd6hBSlgBPZJHY7VjrAMJ
hm1O/kdoytqwdIZTMEss1kghZHH7owrEM0FxDViVSOFC1/8oRx4NRz21HF5VqNkO2cIbZRCOazer
w3oaJYIxnO+KlYCesI7KPWJvSH5L8k5JE6YJ7jyZqvQ5usMpc4v4V5bfPmwOFXn94fqdDD5ZUByB
SS0NXeGlNNKBoIH+wDVjWKvR79DotoNb8ipErww2VErl4xuv6XmvstQ1C3H6eOIIsCRLDqtCXeV0
boFpL7em7ybg78mH2+cmLyZ5zo5k+bDuqJ388Ui0WktBCw1a521UdOWyn/sv9AARYB5egXgCQ3cd
yEfliLRA/uFd/raUFI9v81LWzXrIfZ+92sRyH+HoQtohoryXe5sc6ofduTvlmjiJh/sVctH3lXqa
lZBvRNK8LjE4Rf8C7JgwmmuunHcnkLTOOoRBrf5I/QCtv6X74dSlTePNv1I4sl0cIMkoQnAG9aZF
QfRwmXzZlZg/Xfo39BjJKidDxotLOWJm3d/sYjvZmfcmxTSZR4kdwAF6XRXat2xwfbZg6OuW/Q18
MRNhwUVjt3KfSEaw4m2TnfZa4r4YjEbEAFQjo2SH3aPJQAQ22kzCJs0AzYYoJsPS9qouFLGhv4Ka
TO9D4OFgbnVcDQzCYUMtsq6dRcHG0M8OoXsp4yS0hI1yXOwoVjJGFFZZ4ZK0W/wiu5wjW2WHFCHn
coQ9xHRnSnBt1tqAOofJbZ/cpzDvB1FNGIFAkCyma6lhi7JuJ/Yco/HJGQFoh69vnuH6XkivvgrU
vQ29sE9dMlwAGQou0sHtOipz1fKkbmMzdD94nsy6lsnc9nUMShD4N5C8lB6YQvbQN9+faBrNxaE4
b2BzxqBY4m47BskeCTMsBW+1Y6nG2PFeUmXDKUhNyLIvPDoxKrt2jGkrkfJrZt958biz+es+Gbaq
7Z4c59RMt72j1L0Tg/jw7ddsbS08BW0vNJYHRVuVNnvANTWuUzrYIFG5KVsMp4C0RBTBnepEqZTu
K2z6P0dZe2o3RY4qTEmMve9YUwbjBgy4glOQAVipSzHcx8IqrHvrW94jkmZzIx3NOKqE6NOZYPjd
wqZJ04nXgBlv5yRHdZd+I61IZeNzddU4utdoUYYPqrzhdxq/E5Bkd93yqtSMAzJK2J4c5XiJcwwx
IqKVIf8sJv6rSczNrbtekYOqflnpLCSebSv3a0Gjv+GgZUtC5PI1Cvljgysj8D6Kn/tA7V3xksFK
/eRcTIxXSE5UizEtagou2cFsS/VNqA2aWFdLJOfGxNCA4y1KdE2eE+gYLDbAgvpsbQQGmt7SeY1a
cPpx0zTRZjIM7ON6LTkJ8XrFsSj/F5bfxI22ODJhwvqSxWi63ieaA3ueGTW0xa6+DQKsPyeVT53H
xA9bmTmzHjePFYfwH0O54mRQjRVcku6A2wd2IzBuJK7NejEdfy7Bko5oxVQZ4agxj8jSi7TdLgrc
1vgkvCj7AVg2tno5kieiK93imsCEN6d52keoDbCIroYcnVg064MkFz0J/gTa1Y8DfRcxOz/jigKP
57Mep2wy6EeKgg58oODxqHU41kFDJdNzKefTvzdJKYaCaoAplWkLabBsRIfTybW6uxVpZkVVkbQF
hZM/sLy7AZxfCH5faDZ9sxCN30ySzu05c/iqseyBS132IGE4LyKrI5KDS3X1quNsxinhrvEurnhX
LIvvhhmzd655kdSvDq5NBHWvN4sf8SK7wlrXiXjl+/fQct82WLHs/SR9hGJYS80JyhRtVHAaZYEP
aQEigJ3BS6TW7xwsmKzjG5uoJ/brnTuOUk+QS0ST7+UoWyqp64RTsUkpCZVXiqW7rzERR/2yGaj5
BVFsIpNQ50A4bO3cNK4zqueRgja0veH2rQ/Ku68Cc+xBE+lj0c+Ro790c6rujicFcOHriWIFXoVl
eomsHsMN8Mjsunn02DibmTEc400tuYO7mWA1DiM2A5BGL6JkDAQW1s0KAllHNmy5Tvh09teyQ1Fs
ISbQFOEatWDJVvKNAWZMkn4mm6AkkVOjtJRYxB0RdX2RiRtuqNSUM3OvI72gMpJ2yEytD82QSxHt
6JHEd7yy57xXsxDYGDN5+a0vXvL5y5c9xw3oJqwErJFDlpg1P5RjtWCa+khpORQrHbNG09yIp93I
p8hqHOoQGIVOOR4A+KDNPZYBcabY9NULyKQsxHOffkFZ0aeHVgMC3LpQaNFn/K0IvIPPpXNVByOO
Pco6S/Rp3+0q8ppsSolVHn/RAG46nzIGGfE3dbu7E9ir7E8TSzXDjqBrMJTIAulLbtAfTIjz0uoq
EYPaAq9W/rjuxljbtoY418SQcN45t3c4s334OMMcRIlz6jAbHWi+MBY9JspX4/j540XAu3b1oMo4
r0cPv4Lk8tBA5C8YXc6TYD7Bd1fMhVNNzL8getsDan6U115CzOUrYJiHmF8Q3oEOqr8WkKnGUHLx
yABH2B6L/hsEGoHEmjpAAMdptmtAxU7t23CzmvKoJmQeZRDUEUoVUdzWwl+1jOhLt+0eHSMqq3Cg
UfUr+3BJ6rjWJiS10LOwnkaI7nQNO332kNdr/pFewPPx9GJY4DfrRgZnIvvQhthrXQOyV4nq3x9w
TnigjfK1hpuyp/CFtI1sDEojztjRASiN2ckSzC+qjADdsd5s7rnzdTnnZ9CABC7SBIudOvYZxb1D
y3TVX+UfKWiVl7MOGduTgOnIZrkrM67mjeIMbXCuqnmbbHhur9RaHAE7jUIBoLhVfRNny+QyxhLx
PaUGF00GtgJwGO09sIRoS1q5yqHRhCDuR7vgKx0PCwGXGYs+6evFQZJaUD0K+NKW1UadMLsrkaG4
P5Rlu3rzc4s8/QZJGXEkR1dYjNby01KIjHMkEKOiLkGSZ6xqN6ua5xOMVlQPhgM2c53RFolYpQDv
Iw3u2A+uIoPokRUcqTAQuESAtLkapR7ttVRMMCTBLPaj7uhDtNEgPExAi0J5uOz6z42p5OjayZXw
+s4wR0yn7rjcWF4zLJBu2/H4EEZWK0KhJi+YBt+lVYc6Phgtmi6cRpCd853Nla2S86K5e6qUA21+
gMjCS0cyQWeNFnJ1rdG5MWmz71o8BIiN+Wrpn5rIPB4d0ZYcuz3EkpEVfH7FriItcFfj8aAZotyE
eNiRZn8Io2Oqu31df8IjvuIt1hmk+gHH1ghaivRgK+DmLvM8Xj3GjkbviCPAnoGX4PvPfDnBwi2K
+zwuThAuHMq6SpO0yVGPgdRv/El1I8oU8t0Ll5RiQqZ5HTi+RGWcZNB/lhsvy0eCH4YahbtV8Gpj
nAjRkdnCtVZe1GT5ZRsmM4xdPUKwOYlh82qmk2N/KNLlBu8e4/xek3yZ1vibnv3IJzetj3+HdYby
b9XtoeFm8tNLtwVQ16iT1Hdfm4ERA0sP3qoaaPRy2WDgg4s5QZySvgvjMlbdG/lWtHNLtE6mMB7V
PtLR8QaEZ72kcW3tCDtVneX2f1HY9dTyJ8KCvU9kcBJgUg9ycGzsfg2xAjgWzXj6Y7s+t/23QPGI
gQypRrwBNSYGXcceYV8AcjfdcRpNvV6zpRR3nOPYOjjg+m8xBpG6DwRkhpTanyqXXhEdw7COv892
9retnztS3yl7HE2aPJfnpUDHLTfIDcIrFxNv/kl/jTqL8g61htAeQ7AtXKMzVrIjhuBXBEMgdKV/
/F3tn6Td55rEXw0MfBOCI19gsE7KmaF2pz1fpkTewYjqIUKftTtzFT4qxgtTHtngH1OYkxa9AdZ1
tDJE7J6iRThsI54zpix2Ummdp9PxRnS+U6QTXq1GSDqL4v+ZVBb6rOKe5SQ0O0V3uVZMGlrOor7v
2zY58WT7u3JwWdkNi2PKYXoOur9o+mBD8/iWAUeofgS7HYj5sO93aOPgp+MryVayjVcGGDy2ExfA
6NM5EYGDq+t/ywmOTW7vfateyEn/e+V/7TmnGz8GzYOXr+k1NgzmXXDLeHfTce/nW7S4cXPe0h0s
NGz9TAao9QStVZeks2U1dcvbfTZS+Sd0l7h76Ir0SkilHPIWFZ1iP54MlBNx0lmcGS6BjWqKxkm6
o8maPXR8QADprZXJ9WrDCroFhxA4ZYSU5uc1XT0p8cA6WSd85WpENx+D0tCAIkOmuwg3sxAUnOOo
ggjSlP12zAWGQ6LTulvlAidKeV+pPgXBkuBTUNIBnvFNRin4v2QMRZKm9ofHmLgnt7ORkRbMQb9Y
VM1/xK8XaLafMf/yhB23Sywn7HJwOVsNBHrmUiyDsE/ohiHFaSCWfMNeRYFsoQAq8tA1EtDsnSmS
sf8LoqB9mb3uJJDtEKx86B2D/S2oTCn3rMR3lU8mhC4SVc9QgmsGKWg8CdDewAJQfKRVy59ZkIAY
jJ7Qqp9oRpFR5+eljRwcfDcOPeXoI52KJS57swFznfAURD/RhoXTP5UNuJTYr4Frkej+Peb5cnQh
VFGGbYrTWBTedqMFuJxJYimXxw6YYDNymqiompUrcJ0BAWAd72OGRHSRHlJaVl6uB1yJr4M98rJ+
s5NXbRxJNSvvBcPh4vviCWFsDtT6kSGuUDplzgshJASxmtJCpHd3WV8JpAyp40SjylffIk2dieMN
Su/sGVzK4+SnLYsJr1P/kJ/+KzSVBlvuNrNFwkXgYCUVprQFck5wThuaXd36C5BlDJAuweDhjhpG
1n/4jJhk4QFwTTMiMFQS2lEujwnOyJhGiPcQ+BcUTaPNSiOFbF0Uy2l0Asxexeh4ZOzhLKBXGIZi
WbRLFEkur23bpBYKLSYTqCjtfNyT0pz8RPYsAht+Z9Yp1FGEqEjqZLB/gKsqhrrNvTcgJy0lXUD5
RNGSgtn/kgmEox46NFeBUEUlxWRyqnqM2NQ+f7VEdfUkjPFReCxq8IviKJVMniFx/6cP+z4cReXg
PdPoaeWe1woIf/i5riyaps1MhVoGcTpQB/XzDR/bmNWlbzsri1uYJAPrw90J43HmFd7wCRj50x46
9utTt5yiW3088JHHf/PB7v1aKCoBwpGyPnrUuqhejx3Z73icJOc1wh+d1PSzs6JnzYQNED48dklu
Mi16vbcYzk5pNRJimXslKXkf8GJJ0JX+CKAf4KLYl56ioKrDBrW8oTBJ6HUDWQ6y/l08uFXeQJR6
gc7dhDSgJCVY2JYXzsS3K4+/WbUb02NMFCK6kzyH1TKJ5if356BGhLKp3Nm9UcbNS2cbj5KR+Jp+
6c9HIowtf5k3cblsvKBsmLzeMypIVcNapkmr0bx7piVODPHUnIjJ82ZfegHxVkl2sEwT7KCBB/pM
/zdlUBpziGU+BHJKkbchSh1dkHobwo02Qt/NE+RmjZvVHq3WdxqVbeAH7rW7e9Xo/j6Y4Hrry0l5
xWS7+rf7haVeKXHSCbdj8ftNhPmu1cGVekQx5F37qbfu03dXqUxjrEaESW06JQMyTqtO0oKf8aH4
TS+Vpg5gZUuYj8Qvcntv0IfT4yPiMOmwHrVUcMIOQaHK/rI7+DO9K2hfaFyNkha9PvUHuerLVnBZ
4wqym+LoXru/1ZuD2f41JZsENASglvWMRKzpD2L2ldLCVTICTvjuQr7ia/qTUoFjsFZfxMEb57Fh
eBXDgzVxwe6/uP3hSW+NdXrLcZsfGQwevruq6MIpvlm2nFrX7Sq7GFFd/Cg8c9doMmEXFbZrgQZS
qbxwfjoCQjhly1xR01VUfOdTl+fVsyQhZL+UQHJvY44Bl5aWBchAurJ68nujRvu6gz9mBlZvL9uA
hknmFvFvgI7PL/rF3nNM2fCkZRW1s8cIJgpwQPNPxuSLq+hU2w/z/dMa1QYfpooT9LIQg9Fb9kLx
ekjiV7J35kforo411/zOUVyRjqMBkBujamwYIK4cTTXZkC5Tpugl+ZsPGSfduPzjfYVWYdMQ2/Lk
iw360taR8CY5L1nP+Dw29WUNW/t22ppxmeIR2AG7lIPITALRq7VhMj3lEUoAIMayn+OCAtdLYJh/
4YyOKfbO7KybYFY3Tin4N+MzWT+NHy9/UtV/apUcJlH00ssCORmqmLzurZzYVUVIFnfHNgD6yXhF
iEvrtPQ99LCUOCyig46i+r1QJ6sEs2iOLyhcHxj9smZ/CIbILuKdi00ekQapMh6mnt7Vhfg0epFZ
VCBny+q81wABIF6qYb8pjg4GlmW9pkGNwRpmWsaZHNRN+d1K3I7M9xbVFDNuGJpPY9ahlKYoaqDz
6ogZruZ5XQpSp5dCFEfvsYrGxYlx+sg7aiSu/uNXTCKOEc4bx4L8X0pvgr/JBHyFomKLoXO49xVn
Aa+en3mX8aBdKs6FMUT6eNKfODCfPLmLpTL5mQJd4pNXL77TD0Kh+gW6gKwcUHMF5RwHeIqCr2R/
lkOoaBCdg8zIXyESyR9vQq+12dW9XRsVdnby+SMMELdAhRC3Mhuv1REpDhsy38eQQl9i4xZie3KF
HV6+e/f0vCk8B7G4lKxvodejwXmVQ87M6Tz93FDt/18nMl60MxzrCQ1yZmInAUVnOuGb82ZOeALh
/IjtO1zldPncBVNX9IlN/ZT0Ann3DmkkOdeJKitMbFCjvd0Q1M/9KDOEFe5c6b5kpcgrgLAFh/+q
ZOgnJ4SwFmMjoro/O6wdKXAMLaHeIPo2r9cOp5Pfrp8v1xFpgNzawURf8U3w0LV25tKS47PML0hF
ylnkvapiQz59xWmnGNzloaRE3E7FFdjTMlPoskULJOuL2UAwvqOBret/1ExZWeqHCs3BPkdPqhiv
S/qCiXMN1f4KTuRoVQuOwWZlv98Od85R7xMlk+QpLlWLe/k46CZGdgLLJ2J5s8hTzaK/v55HkdL3
wMhZXGMoR7skttbadWSai5OJo1CYUL8RrC0rot9iIvzbpg7oVyNEVkOc/ag8+hFjsrhNU2FCo2hJ
yMO2RiF7slzcn/5T/22NjM//wy1TcEoBiYLBWaaXKmo7Kt2sD38PSfrg03Xgij6LCNZMeW6yLaBz
/VW8SgJxxOACgUnbL0aMAtToJzU1OuImW9DybVrAxNb6bQB9gqOvxc2l7rp9U08xWiyGtj3Kqd7P
Jlyv6wa1a0f9MtDO34GxkNFIccJ6myh+5ZvWf2crayrTPclXpSTZIfcBZVlYws71E7v265QTuBwY
yNrAWDL5MV3HXp9HBDzDf7aI1fkxbau0n7hnhx7gxhwxxC0cAfrnHnavtEv1oOloheDAGJpljwt5
LQjJFFEExU5my45d6H4Bg2my+vtcvp8bMf3p/gBfVuD2z0emHQms6x4o8oduc9R61qqk5viMVTpd
fExBq9NU57rL69eVnVCuUjxwbpQrm8BSV46QFR+/3lZdT7CERRk+ynieYoVWmTJ0P1JyIY7Tsda3
Hc3PTpJTkKtYDPp7u1tJWEt9S0eV/Nh2chqb6wKnmSUa1Gg50OF+5GJOdpLsd5zTgAVYZt0oMasZ
OBXeKIU91QF4yElNShMnr9BhGvTo1ffbBCRcxwcuQVVskve3nTkFq+BSFEXk0Jrj2ilfb2f//Rbz
VC35a1IGIOhzh215n6ikr/TIHezGglvZme2Qj+0ALNDPZ5plg9IjARlnnrkxT9HUbe4QQ0uLzYu0
i/w+eMVBsSQsv9pbWWOHTcsoVmJw9LnhBV1AVpFDgCq+I+ttphbU/hcTyzBHUilrvF7OXM5OXTtk
VTHEihMap0U85sHrCdf8bJ/aij77uYlvv4ukwPa3H87MvMvYoLgpGtfsiZMwPpK9l+KQ2VxVYLIt
EfNw0hS0c9G24DzYdS8X7YeyZteM9JwOqEAVYZ/Q980ZrIqvo0Lh3diXt55dBIYWVsSLkc1QtQCL
07zfr1S3pRv/K2vuzRHaYkW283/ldU73T7EsFxMlRdLT1QhuO3Yb64uiCYrXtyUH2NuCORwQqdJ/
LDddeBAVLKFBQMhFzCPxo3Dexsd48lChlcf1i78KYlFZiPRVJwgjWfjOwQmRjM3eyWm0XLPpLuBl
o2Z0ynbN4uPyOduotA6VFP9Z4dG8hmRLJTbqgx/9hsGGh3an4KTEq/Ze+/feTkiyirn+gcRlBVST
89qOwxn0PfUpGeq+avIAPM3Q971PD82bljRr+dG1noDguyotOGN1h267YCQgHlolopgYMC3XhqSC
EZdTtKDLAqPVXk9NUdlzoiLLw6ONRaCsKcaHF3AfJnAKnTDYDgdmGS4CV8zJvaaNd0jyyyz6gNad
5KkrNykBb53GyPjq+0TU+Gy6W4VmI5CFWd7SB+ctsaingh3S/dHnZJN/+fTYaMmZcKoXPQX0iwjn
yctCur0Jf7HrAB0F4hB4nXJU53Vzi/rwRdWH465Km37IDB/HIiKbU0iNa1sm6Jus2Wd8xQQ+qD4t
d5IzzubXVDz7jrMN3JrZuWBdtKQt4uxqg2sxJOj4Vds9xTVr5KxBdT9HH1MCP/99Wru84xd62l/D
vWzSvbjy00RtC1jO9rdwR4s30xZPKXC3IfDLED6XluWiJUmGFZPjKeHJb2LBs7Es6K1qHfwQBGOs
pBRt+FHdufGEe9jy/JhlMiJkGFKaT7DtnTOnClr5zALgA4Hzr0ioVNzRtG/nMZEMNX2SkUghlHjo
9mvAB5bbXZlO+ayGQH81uVLhdYze3jGkoH9Td7BKYdIp8lvliCQp8mTHzj8madaMBx1ImWhz40qI
AsbuSGm41dervZ8EqaEdavvS7jriVGRWApti/ZAf0bwbULOIqzkl0+aLfUBpIqi02iNLCLgpS+SN
oS1UF12t7Nobmvq5n4GninaeB56rBwKFIZQG012L+D6jygnREGykjG0CwpV6P9+/AtFbhQR/RFYy
r57UsaYuPLq+pg6/iKaI3GxLTaanfu5N90aQErhRN2QBPts33PkoDSOl3Jbo01Flr0NgtueZGixF
QLBgnKzuAmA9O1YuOgKHNOY1v1xNES9TgOO/lRWflhXCWxbdHtJxqb71KzK93B74Mxus4wKwfnTE
s9kLSKb4VVef4a2Y2QtLEyoskWhDW/GRgpUsV72xOtvaDnSLXsJYePJY3hvV6f7Qp/H84MeZyW+b
5hG/lD2opbbUCubgy6JKTDu+Qee/3WHeX2QFfmm1Y7+xU7CSZc5EU1aGbe+OYdN/EIQceDGGYFUA
a7Ox64+FrCiZyOzixD04hCgnI5ZZOy3ls44AmKykkGP2fj75Ov278NxXPhpGHLn0KOpqvW+sGQr2
8z5x9IZc9XXKi0cCjrBCP//Ns5ROv4YAjmZoDHDPP9Zo6E2PW0JIAMK1YRn5GEGkQ0Idqz3kjixK
YH6ANiMXGAr6emifcvhWPdMct0fP3jaZQSy8bCkC3r+7j4ONtkJgsGRw7rmZG3lfMvcFKoMpVBEX
9KEgX1cy09fXYwoG3Tzo59444u07swVo6iX5aEtggW/9Gy1qX17+S90D6KJSs+vndY0PF3cvH8Jw
TYn22+1NfWwYn6HjyikDwS/DW6Um0fmMrUClVH9iGK5Am174E5C36pXSND9lJB2o/ZiIE7g8uxCB
/VPTvPml7IigJxeEVno7oDH3BTi0f9acDYNLTObvmcXrJICmoYl7jyJf68TDjoZpNlJx3I8nxkYv
EcTw6ZziLoI9Ga8QISkWFTEaDPwPm+Yc9af5WguVabBHCFM9rCyAoJtfIBfoM4/dSV01UNM+yNYV
q/I10gubeNXwHupXMMfRDrT8OxNTvPNOORzUQvHeAAlbR6ZqrXhXjXxBUJDqyVOdiF4eVxv/uKSA
g0uIzlvhCQrjSkgFr5lGQjkfhsb1EdnhdZ3ulTTEBeqeo+WxmJniGZcobrR920ZyCWh2OU5CTMNv
Pbb5i/3zcEmsOyVSjAqIJ2yZ/be4iZUAjlFQWGFd8DAbKdaa6j21fcHrlt5DWEWYJkZd4w6rLpZe
esCOJVcJ3I3Y0ug74uY161W5LwvDD0Y8XCWQh2c4wle1yWSl++tDWEPcxalpzwrrcELrpR2EwJdG
654QgipbCrg1JrVtPejlIcIqhiYEF5tDely9Kr7pgkigBYZo8QbrQ31HNqOQssPqBjYCZXqcrIM5
i23XmnNbaM8deyTv33L8A5qpn52fmdorc04pqntNtIZCzdtErLQMSphVrWlfUn6me+Ufu9OAPGk4
SimPRI4kpVxqaQJ8HxcmsBwy5NLdQMsJRDf6dyTQ8Vkknag/n+gyRziPIXcxh66JU9gEZ5LwxIi2
GoWecqYZ/a1s+XditoNiD260YjpT2HQq6Zjmcee2BvraN2Wkt1iWNzTwysSAsK05syyCnrBouzim
Wox2jafekGnCjxLuXgHhVqBImaEJhHutrYbcM9TZ8EW5hItPKFpPLQElIODUOrdpDeFsEEhYfpbO
MWN0HmAY2ZILaNpeB6lESo7JtBU4kaLX7IKXJJncW/IQVMCkSW7F0dULrEYXRsB2Wi3A1y/Qtt6c
PI0Fr/zC3CaihdglDysd7NU8GUFeV1o178HMi//LuDCZrAovSKK2jUxtUKnDOuoYUV0wFtsIHNhx
ECQOcV8sJEy2jK+SMve6pBP1kDNbZDwOIE62HmAzgZ9UDZN04Wa3vezIpd+YzgaaVu83pywp8ixG
TrW9FKBFl5asx6MERBWSv0YoBzvyGZbYrjU3y/sQlE9yU1XYNYHAD1y8Mbf9TqPSg0ncNAqyLESw
Q8mRD682Vcxdn6IWiwBE4A2v7BrZMX4UxLtoWEd3tsogKwOZsFUbhs8jaVnM2HOhWy9JyPRX0hzi
mjODLFF7MApWKoW2QukDjsEpywJL5la80znn6VWhc2Yn69RGZXiEnUxg0u57S+jRH9STdfyxZS4p
YlD79Yq+Tf0U3Wj5qMRyV1dDNATHiD9HY4+/ouCd10EyATnJjxGpUyOyO2qjndpO3VPqjpYOGK4T
QRLlCRegFH4rZlEW5auU07ObefdjYEsb6mjwCFILzk/rDvvkaUu9kNV5Mgg4E2qkWP7NPIzrajg3
IHenv8l4zNyjpwk/M5+F6z7M/dGG9xHLvhcWIYMIaBTxyCk3TWGxe333mKejWR8xznFRMma9OhO1
XbpqzEHA7JypjYZ6kZnpvTGeWvg/EJepqb7b4o/ckuFA1hJYodV3FqX0pYrvpVZUlglBIThAbtQi
I7kEB70PLCOu7B7IDR8y4DOu8uMaGe+XXZGpDo56+0DMZpZtZ8wzpjpRwdSbrcqrOJahLGHoppdz
4CiVrH+Abbi3vKAlaGc7dZj9w1fZn37kWam7LqSIsKXY3EEpu7gGmDKkM1xHHip5wltpAQCvdXc+
nBWpZ9phfGm0rnvFG61FgB+NY02CpblP59GTVwcMlp8/iXDN0aOjpzNd13WH3rfAmEL4jiHPsogP
4G36tNwOp1kbWoJ8+5nhFKvmn2soe9A8XfiK5anlxh7df1HxR6xfYwYz6KAHuTc3QX1CXPvIivOS
aGzMK8RtsOCQQuu7Ajya8FM5loX0RjPmtKu5CaANCDgpYt/WGgwm/gfeCHCWVzEjw8pWZvTkKvzm
bsGkFmm/2W7UVyUw4GlHIXGJuQ0z3KqymDBro7P0E4a2iC5oMWWo3sldAtjYwBGkEFWIDt6E/kTS
kYOxXj0gWkdFV+jsdnThl3nwAVUqT1f7wPyN1w8wBNIqtz8ZeaQRSBDYUU4PCvicCLpxBKCE4p7c
NRtKBFPwGR0D+zd2Vbi8gLSJyrEITjwSBCaOwR/OZuwWWByaeqlb+Ccr1/V7gmwjRcWcQF4uRVkP
fHnPPbhEBM7cjywv4XdBl3K0i9H+WSwRltAiRhi3fm037Iz+vrAGxM2I0oGfvHde0E6xvRnIaTC5
vRVqg1S6RTaeICcDQCEIouxYvEcdqpMd7/8ASljwuAXONN98usIcN4PexdR8lrYVgNK/OePKAduD
rDlE840Zm5dwxoSVEZzJkudH1Z47hk2RsM9EX+2fkqsCo+WdIiA0G0t7o2Viue8/eeQ6isXK1JHQ
UBSxcVODOpOqi2RH+2+5bjWTdaB+IAZGagzuUA3sbva1uGdfsc/6eKfXcoYlUm6E6n0sY3bIZFt+
wD7CwAD344r8ygispGLrjuDRtcRTjRLNncBlBuKSMUfhv0Pwa21c0VnZxyIp3rxbv0dbfwc4c63o
hD34Ovs8UharbXav95tTHi1CAW6OfSWREk1mDRFKLm/A7oA15Y95OVEZTd73OYsPtNhUZehT1+VO
adYGK0HaxUnlFd1+XnOFJF80sBtwTpf3tKVnqfKNwlZDYjFvIm8Oz6MPwhjAuif/mwU7umpnBP9V
OqWWtNJDiUP1JPCeUO5TOsF016CwfhmcjM7FZsGxdP72kSlAYwPMlucho2LEWniNTi48dWfY+K38
rXRXZLD33DqOX4she7IUs2Rch5BCraUweKMmkHAXvCOhezQBx4RTxcRfauFc4+jH+idKrFfoL4Dw
Tn3smeHC2+lyefymzUNd6cnvB5lZIOVrNWx3eGM5r1yHywX0ZynliEH7eBoi91GGP2i2RwI6a6+o
j3Aa0bg5HusALd5zukHHX4wI2A+BIetgy1oLf9s7bp7jHCVRcoA9iYI404/WKE7lUkcO6fHpeayO
ZXP5xZg/irzwuAP1Wpu0Z1y/aCf4QW70U7RysvkSgk4RfF9Ucc9G2D8fWvixoQh7tSvR79Q3zIkz
wQyYZtppqnpXaNfcocHrLqtr8LFkBw9a0yd/yttPUsPP7Rlkdx1ZeyPZ0rNFJAuUGNjWHq7Vi3XN
uqUQn0nOlFqxnR1XKwdMWrqHkxJd98W9Pzs3B+tTYFHi7XCVGUAwLei5iDa9nlSTuWO3NU37TgyJ
DGCIfxAp9eSa7B1+UDoq6jN7iESo+2E4q58Z4ytYY0uY6WeYLrGxefbwezYwQzdFyf4L32enDJcz
5I8dtC/79mjz3xG5/JEOwnfWNFU1VmvAFdKL7H4QWsFhNRrXTBLSAQPdWMZI1uW8l/q/h9dpQSSl
B7ld1xYfJGZZzEJv6vPlNrNrvP1cWyObGZ3/dWuiBM3n/BCLB6WcUkJ2wOCO+t6BfL7gTvY63Jxg
q4ZQDfvQrNsUPsJ1dAQ9QWC9fOeiRLJnOqmQ4QzvTQpUsfiCEpQvR9g6N35eoOwhEBmvXPk0fjaM
UGOYa7DCgEtZlRSgAvBJPBVaZI9ZXYZjH7ZX3BQK0/HKlXpwWdtbxGEZ9zsFDuaZaldRrqXYiBR/
pPFT7DoiJbfgReOVZ8GPkYl59lpopl4aYgIJTG1EhSnYIL3TDn7U6m0KvEszlNMVPr50j5IRKGbr
uoCav1MtKRryIFshD0BlSjORI+rzLsq4jk9S6J7T+N6a8YtdcvQsALsRL4j5V6NDAScm3MC12H8H
U03y7RwJHZW9vXYCbJGTtmB8JT9j5SP4TpiIutHfo1DQ+q3JD0Zsy2pyOQnveMZuhxn5LX2DmZ5G
QH8E2omh8BE/uxVkOEd5Bxh3mzmlvDiW8zH/q8NStdrsCKNJ1LHIfgRgPdY2DIpthkym2hthVCO8
ghOeUfNt6NeJt23zCDeckzI+tjnq1gUISuB6nG8ey2n/BSmSxUK1lFKS0mi7r8wlSBC1HuWZJnC4
piNMEdNM6cw1wa23YClYFlUca1+H3xg0YftDTlPddqk0q3yJPBhc+wWji28G/V8e6BtAg0Hqv3KV
W3KBXCc3pI/HpuPDC0UrxqRFRdhxVKCgICfjE8242eHA36cQ61D/jYHrhSFqXjnHBpUayXKd/CDL
mEUJv7peXKmH9Kd5rHNJs07jfpNDC1ohoqRehE2xlmt1NeX0BxJ/NLeXibYj14LFxWAQlx3kpkIn
EpOUqYoDzekSeTINESvjaEtyPoKhMRw6sVdeG2jzIoNflk8WNEjc2Y2q8af/3rUikV/+nSKmuo/y
AvghsDGI93zptXiMx8UrzXqp9wAC1XGyUiFR9z1wzaxZwKRsKnQDymYgWHcNuTZykkCa3vMFO61L
TwImcC7B0D5LZ7vyQ4Xw3X6npUAP2YRe+2Df3tQBI3lAfD7b9RPeQEzYavNFQ/lwtJeN6pcAWmXd
lf1i6jerEk6l9vg+Z9Wi7PMvj1clnT+d8ED7r/oWI3fuw2WLr8ybyUoJleajs0eF4/RqjTQ77t8j
Ss9oVl1JC3Hog7vUuabQVhF2Flu9uaKvoplocUZ0e2uxpBAJ2LDdoVBSnMLCw5RRXUuRP4H+Ir5c
ks5xGo9k/KTP6eSxhGhYXHiz/bXJbXpuYLHiin3HJJltrT8KfVpBWie5YhZDr6zz/mEArj5B7iQI
ZLxGCUSGA5iwpi5GHWd2z7fhW2pW8A+Wdk739VoKz5R7t2Exv3K5zbhInqYYQyyLeA6+bASNRjOr
oYKvx1TOJRuOWeidqDUozIxdY7xJ7d+dvK0VpA3c+ghqvRlzDzxldUFQR1Wc9MV9MbYRum+T1n7h
hfCYRjVPqovbTN7WVi5W7PuOvIe3DzdDt2N8sTuPu+F5EJc9AXASebgRU+0wpa9j6c8wA0VvSMLo
irBdSy+bRLIU9a9GkGbUyONNRLF9b3NdAPT+uidRl+v4717No4jfdH4Clzd4b7YdYmwQaPMGG3fr
QmhNRu/DXTnjfdu8ZCT8z7PxeaYKbPrJxFpzOAd27L5rFgzq5tINfCyNbu0ovwksSZCkEzUh4QYd
whQD/CkkkEsn+xaoIxQGhKtv/DOasaYo9RvRB6Ab5TCd5E6EA68SwcsrdSS3YfuAk0eTmvTIgZiH
Ed4QSibmKpHe11ylGHs5P8ShvPbu2iFOWEUuAA4yoIx9C7/+cXCsFNcnNhUMXfjq/XyR0B5z6ROD
tG7+Wz0rB59bCXmn29XgcDnQ6eArL17m5TtAIB1MN0bh9lFoMmyGAZNXbVFCbnV+BhkcT3q2+KIW
pg8fl0/aWAGpwcgXWIeWl6ZNixic4RWU5ec3ynM6+RUHWSNhEIRLtCx+XHSgEPrvBOx6Kg87r8dt
CEakEgdrSImSw6cbeqN/hF26NX2Q6/kqEDjzYHDaXBAG2xatMmqNCSAPHuovwhEso5JpPV+colg6
PChNJHWVs6289NQHLj9jyNmXy9SooTtcg+2CBvdtjBNOL3sp94TYN1pqAR+QtnBoPPkJGIlF54QM
XCIyVB+/VSMWXXaVjxtQA77/A9UBCKSDYmVmPf6WENsoJbC6GKJiBEKxKhHQxJ6dIELoaQTUryVX
lGgUjvP5vteZJ3GS23+LtbZgFjAw0U2F/bwQRVg4E+T6CdrB3nIR5pmXrTKJgRybNdbNjKhjC3aY
H/hpEe9iJUC1/9+B0QXZPRL5LckWe1B7s3aSBS1hX7CQPDuDuxAVgdhQK5sgbbLEQFfUi978er/D
nPrrNp4Wf2E0wRYhiYf2SwNlhQM3bjw7YInrBDy5h+Uwn2xZbeghBoDj6bctr6tUiHjCb5br2OBO
tW/SeB2+16pznLZEfAdJGor3mXBYG17Xf2mNoxYl50Dy7QeoC66Wkekte38Lx6rfefG0s4FuFolu
o8cQNRqA0vGEkMOz4Gk9YMYPjRII4ECx0Nllld9uzvEVgyMyd5nV0TmvgfFnX47tICcYOgJfHN7O
2reQoI4FVfjbAAoZctiYS1lTRx7SENfPvj75tSVIkMGxwCLjszzkTrE7W/HgQXE6yNoC76+a8n1V
HkJQlzwTWoNT/9lfUWQrepjh40rWwYIaAt6zommDXe6CpuqiDSxjR8meS10Qu1aIyvdZzhapCMg4
I1UuCLM27gZOoOCPcXfHXEN4M5C759HTjRt1DrABcbFX/wE5ePaWSdTcAumVygNeLfH6NT+VqJcb
zCUAggWeQG1Kqk6t3qXG6Lot73m/XmVB9Wpi2MlNPnUtt+dIOeRXhR6eYeVdEsWo6GNc8ZHwy8JT
zNN1rgeOFBI/CFlVR2X+mJEXTliXCP2Trmi6BZ9KZY2mvFSbIkLI0LIxLaFOXfq4e9xEgIzlbDg4
YthYx+G/lpC1bIVMB0SmbTA72KqLyRU9ZiLTlPALlCY07peXdoRWze2FvVeonNxvCdNEYUooR11e
8F/mKMH2xxgUWEBrCUspr3C8B8+G9raDkrWvo8bBezRFdxnA/+dcjCtYirvAsLhZIVUUHIzZr46Z
wkGuCFxElh0BUWg9bcCdw9hATQwx+QTQg5JUHqp63fpUQSMsjVpmbfsjUepU56dxndHMxCeCUNpL
OLtT3iUJCK437NNpFOBYTKMa7dtOcKhpbOTdOsUa5in3NYMLUqAPsOMV32XCZNOs16cDqzfZuq7G
usAqcR794csg16L4R7h3M9J+bYvZjavvNhWN0XZnMQbLW6fOTXiFPsoUz99h4aAco4mYLWJeJ4TY
zzUZhJp/ZyMWzMKXIg3wEh35SVPypvO6eusu2n+YM4zVgSYDI8P+hNsf8vY2ulnbOnX+0yDpmGP+
p+6QPU90hyvyUHpmTMNqzLxfEUK+XG7bXZQu1BoTSY+YSXf0QQblLUhlRxWB3XD/s1vqUG49TaU3
XYF46Y6fdRBnbwvB3aHl9yiNewF8JU+5E8DOP+dMWKnGdQcuO0Rg99mU15Zkzi14Md9e1T8Vj9QG
0+JyFlkjwXSRmYnpWtPn97kPeG5eC1NUeLtolg90ATF244jff/Zc1yEaVjpDaEo5sfIRf5KEg1M1
NOWDNH/d7QbXxVQxGr7pTtKA96CvJPun4KaudKKAPGnfkwTwmbVekNDsPRPhp3BsrH8Vb2vxARxZ
hevsjQcPV8ERLw+6QPOLMpmgT7ibIDk82c4dpWACCcvwUN/w7AlMjjj33ZMcL3EwGilwhPa0VhPq
NXIJCS4hHSZtgRbEcH8yngZ+BHo7fpP7MlrSYAHUu+pBLacTre6LumwxNjoaPOI5j9/gi9HSS6o/
/irknvf90b6TSBejCY0jM6NXVNEat1xzKNBzf/vCnuVoAG0VviGvJieZ5jwup+WQd6Px+1hTCclW
zH1WgjhDzXcZjmgVwFx6mFQRZDXV2LvgSlbv3BOMDtjXgci7MNcA/mnFmi5vMRC86SDBJxGmd1sx
uI6WexmaYnBVTNz8Z26krOMJeLTg+7zKWa94IYuL/TnM2ZPJDaG/OVl+d+zWsYhGYOrMpvv4SDps
lrfNY3bwt+C5TRpo+pQtf4otqkNZxI35FhhHPq8382+UJzKGsObEqLIoh/K4oez/1WRwC90/dBlt
dG5OmpyhQgQhxo5xGa2KiIA/1O5PgyPinrHywlN1pd2WQMqp0LwGtDfMay7OckMkQW68llCDtBYX
qZtXqHyGfy3/q6DtukvXYlRUYYzd8ZI8Tl4DgciBjFqhqrRQZ2kX3x3j3JRWp4TOGvSNezh5TNs1
CPYYj5GnKqW5ic9hGOUj6pJNVwBuezFTtYP3bD4WMFXbRhpP6gvrm47q6A5W40ZAUBJhaQHX8lno
btaBsATiJbOOt4l49eIyPFoEkiLoMyBjiGunOlgc6JGTgXGJP0Qi+v/t0NoISV61yac8+ID+NZ2t
Pw6HF1xGn5q0a4U+OCguRs3n81RdYuJzGUqApdUqrhk4gjT/M2OGOM6GUL8Dcwi6FQ+MaXq7z5BI
KvaF1mWNsHt9Yckq8orV1CeBbu+oxra4U5+NOPcU0FehHuMwbbRPZJref4m+AVe5ub8JpOTA2fEH
/kXzCecMBBc8I1qlnuVyb5qgSlAHvUghT9JTYDCteXGeHgLkRr2CV55vyGHry984N2OOU5+gPtMs
P8kW+wW944zhejJcjBvFyy6m4/GyjJ7+yOqzyNsKzU404zlMKF7Nna1TisAMDHRMTUDa3zbgFCxq
7swlsxvr08sdg6SzSfmzdx4nymCO/9uEMN4XhjsNxnpkhciRyACTtRY0yICB0K7eUflKjOMKapXW
FB9x4RDUKRbo9bSiXu9M329hKWn4NQAv9BlqgYyUJoUWwJ0d9rJqKBSRbYLsLsX3mXIYczr371SR
p76lLxJTmNEyGWy6ekVv2mb6QBcwRq09n6NHdsWAaxTlqsm89zEgAcxBf2gWRCh30oS3pXCn69EF
XD19OCiCzJKT13crLC67zYNB6/e/OLh9nJQoaIWqfrjxFzcnFW0YOZmH9UysqYZWEMdCZdwQC2F9
ryPD2lZM1OyfW4E7ICSeWbKONCVOYChhwAywWQrzSjIzFoEgNbNi5Y45U5RJ+nbvQMfpRadyGf/v
UxbPxaNrZJaBfWaUmemM6M+blLXgvLUMwPRti1TnO+9MbzT50DtpqQb5PaM8kHU5gkv/ui/TkeLF
GJ8+P5FDjps+X8EE3GVxnby7xiZonVoF2YhMS2WMLyDYxUP5E7HHCBa7BTQSBbUDnZTU4FdhG6jn
YIcps8KsmfeXccAiFXn/HbJb5aFXuKkN+IeDa5xw8eOQiWUM0OtKm1bUfKg5ZzgoritcaIpqvuuj
Q8QtU5/JItjYX2n+Hq1mUlqscqNzrA8MLOkMOFZj3Am3Dmk89zjYnJhpxe5IQPYXj3i+4B66+Nuw
R4T9FRpmsoNWCvVoPrmswxa7h3tqCGUA1ppzjy0aHAHLOu85yvzvM0CCsWTjQc2hlaIKArYNpLkf
hzfE0kvIgZKciyneimvJcKso3yQzsoYRpSnOVFyVW3i/SRmI1XYjKykfjUqjCX2wqCH7bt4H0HUj
ZpX2STMkL93rkRXj5SzE+8c1OFRLTJV9fHWdwrHhO+FogDLxrr9ruEdS3E9dwdNOAPEiq7gpc4zv
YpOYUKBKZ5d21wzey2tyQGDXgEHiGMElE7DX0sHOBVOq29+PC6l/8RXrAwAgWmxRKJzl4BHj8a6M
Dh0Y3S52N9HwgbNfxGXdStVlOIixhpyueDRcs4+rkd8yetWnihICMc0S1NUfIm5trzXOSrTSKBR5
6KUOOplojkKu1KJ1FEa4WeFY0qRLvc2z4PHG5SsULgPbY96Xn8qP1bjV63VC2xORS/BJruAa59/o
IqnOI13cetSgVbXR5Xe4LDJQCYybJH1HA+3My867bDK1uK19904ly/6H+UYKicHBXaw0Jf3MeY/e
iUttstQ7VR2bkG8D2PbxbSuJCXdstljWtZgHWWjKz2QUEB8XSVJmOTeWFITy2n8rw1MJCFKarpu2
PRKBCwGKnT5MeegFLdEKo/Df+jE0c8CLAQY0t/4uSnpIZPukAFwAyijx/KFGAUIylahoW/OZEzeN
mmR54ZX3FNzkuSpxHN8JnYzUQQhg+4O0lcRpEDyi6kwObcsJEI0DzoNVScjXDsMIjrE+UAkW1NVr
13PYYql0ynCPJ5RRqJiHiyRXVhU9vkwOJtyrFcBs1eUI0CxUSTrU8asEmUt/rHKln5MYFxeEHveg
xc1yfFl4sYhchU0hxaUWM8d6orU3jJF9PjIUleP0zaPTGq5TauDB6AMWZmMcCZsRg21oKzQgemJl
YpaaJm0H83VAWkyibZ2LjUvKPR6gX52UUwCVTeieGlx1vvmMCbm2zfbUcUDMauy/JHpkT4yOvUBt
a4Ze1ySzC65awV0wzUD/6yKy+ASdWRuNpJasYpgC3FCrV1T9nhTkrxpUvakP+D98zACqIvIPgTlJ
kIbEgb+Fliql/I0lJ3zZqP5f6Tlb+2a41257FufABF7WqQ12Lls17VEjn9wTjufSA1u1R+sGC5TP
lP3rUSo09a88B0Jiy69F2xoJqpJW3OkLsp8NyPXnsG9FY4nL9z6YCXuIHpFwi+H5LR6EZTDPXRlC
wzZF97dDlbBc3BusHAh84WSU6DeBJHdrwDBVkPg4DYC2pi5zKrHhLxK2HTelrfuckMz8XxfF8Bl+
6l41TZM4rDmn7QNsasOcKu2SGVzxk1pDVQ/sx3f3t9rsEOKBa8LB7i+3u3brTxkXZ+xcMFPUQsKk
HIVsNtfjOEwaU6Dz1Mu7z7PQO8Vr0LJX9yHJArtOhah17D37H4ZIsJyp3SmZgeRAnLcJBGNWGHHQ
4Ahp5mxln9wEXstAwb7Jna5YtRL7HqiBKK+VEQ/36JDp1PDViPcrl8OhObSHrzEVvzYo6qwvY3l/
fZCkF+ocSmgjX4uWHrQ39Ouu5vAGnfCEPbvO4q8/+3OzcM/SRRTtJnttSYFUi1cfS8ORhpIAIovF
TNQaMBiD4MRtryI/VX8E85xKKRwexpv58xXlMcGLID1zbOcn60vGf+ccsdsv9UteDszDZRujf2Zt
lB/YDRNSeaIM3II+tmxNPcF3w+fXL2JAYFZWIQY9uf/IHH2ZQdXCXq/pDpUt/5HCTN70B6hlPn9z
R119JCi4nKr4anDO9e5s4Ndzj9839D1qB+TJSPWx9DeZwX8y8p9wRfzebyhRVTu/hCo5SvImBFyz
wz2jkHXHSqxYWhu3DRzOJXs/wx/VKSuVcoXDZffXuglaegNk5s3hEWZOZpiUXcd/CtOe3NxV9JIA
hbi450kczcc/y0Yny589cnn71e5Kk2wqtxtptSARl91olX3fqpONWAcKjPYkc3AD8Bbgh2/3uD/+
yRObxErJ5a7bQjRWlEuJIdEchdePVMP+gLWmlpvxqhO8PjjmnHGkw8m5yRosD9++QP0WYpzFQ+Zd
0nQdoDufFpkqkwH7YepJflYEVjWF3D+/mWYnskzit+emZP6fBGICJEdpqIJgiomA/qry/TmeYn2H
pZK7DMoRcav0TtGsHh+ZmWCrikvWkzOEdIyyE5xk6EosAP03b6dMPqCkrqNPO8TmBDb56oZmGLAW
eb6788bPIGZE5hhBnoztaEhyVSZ7/Ss9ovGCBYdRm9YGcoZ6F03hD4dzjCyP4Q1++QOjgWLIRdxq
BeTb4Tv4toIUomBOM13KOMvTc+cpjtDyI91149048oEeUYmtq24qWNHqBikoL69jSRMg9eJ1jjlx
dp+sjlpNXAou2rYjb5elzwXlqto7L7V6kyDJBI+bAhuQqXflp59N8ABDyzZjThrTf5Z8/4VcDzaD
IO+qh6X6qpxbVuw1gzewwbg20cSSky0koxXpfbv2qcMCOvQFU4tfOMDDRGHQDPJemkQSZgwrHwSA
v7kvbHBRceXQ11TjrvyOeeZdwsJN0QZeZJXVz/ymvlQkZ24gvqWyPiMcLH5awbLHfAQyylzzalLp
fI2tFjp2/lAfynSfFk1BBstNDmgbeNOWu41/sCAdE5KMhhrpxnKSXxc18M5vZ69BHEeYbFSzA69y
bb1gqDn5Fd32/0UwEvQViEHNsGF+NfAivu38NA8GEIQlW+/feIKHrfH0zZ73LEf+p1LOrDQzLaWH
Mvl+Ro2WZ/Bq3YVYGkUbQie7MQuGIwgf06rCFDTWgMYFari0drA97LXLprnl2TASwEhMeLnANN4t
rNyjE3HJRAWgrsg3yA+zs/fLoPsCBzqLoiQGBZ8vBC63VPaU9R+VHMKroE6SAvcfuqK2A+iLTOan
xuAH0216IIDLrzs9bvGFN9JQfqKblKW56dBFeCVb8AMBe+og7x+A57hwt3PVCJ+ICAZyvbXUOfAI
NtlJmHytF2SOaNrQD5KvuVhL7JJizvT5h9F8EAaY/UkAm6rLlyJwes7qlDg3gM40LwxbgbKxKDd+
daFgpl+yDFqd4YPCGKm2Xul6vQAkXvZE2/LjuQ1MucTY5/A7thfv1YI1DQw6RGJw4m7Es3OC8000
3xXSHjnXcAyc3jQOQxYG0ZLYakxLDcesU2wVlV0FbInlEd7NB/7ImSH8r9YhFJNa1sHaFl5dG0PL
GkhbXwbgyMgjpzX4kTpWLlOPrJm7+PbMxWnNh2RXfiFbZBX2nzsh7wcVcXpk5p3kcPdiCDcdwfyZ
KXNJq05r2hnQ62OK+ODyCH3xlQ/gBGMzbUjtK9aw0TsZRCIGnRdUNOqQsAQZ4/LKfHnmwHJ6Fact
oc2vgx3qMeij5mY1gJKxrSEqJEdLdI+SFjGWnI+rQT9SVw3FSL0v/dW3Ml4oHuQXMtjiAEGP5BPv
jnoqwrnJdliUmFdIhpedfjxcRKlsE+AcKsX8JLAKn9FYutKfoiXukS/z7Hen/cZ4lFtP6Qz+xRgX
zc+IarCnDKdg+VIvVHr/xgsVa42yrSUcPT2ofKLI8xe4XlhoPfHbsX4DjXB0WhTz7DNeeJEeNgPw
r/5GXraOW78Yaz/ACDK+lQaXhMKxtU9tgpvbTZmtRZfE7OlJHn/CVa9vhnDYI3G/36wG8R8Pp4sA
A+l/1d4Peo8ho30OElq6CsSe0miQrgDU2IrlKm4nZBTM2SP4mx+fcalQHe2/7dVIPGL/sXyFw+AI
kf/5uWVx/TX5KQm+CS8Tiv9a/gg/rp478hRNz+kJ0nNYxT8E74LZuhSx4UEIHYdVDE/ysRENkmSf
juBV0CGJVUP1cHH7wz/JSzRLfVqbQSAr1Yo1H/wELwv7MfI0AtaDbtz/uEACtq9i2ZHEQnaAT76G
whDbj+DTDBKzc4jRqljUq+lXk3iFguzC6SlHtNHcPG89jg3wt4jbcynbhVknHerUc1h2zscoWsBD
CHhsmiIYJh41Cdn2Qk5jxdDSXVBrlVRx4jXfzJqwX5CA4IaxyTH87uT0kJ0G9+xRAx+LvZZVVfPN
zQfJpXOOPSTDnXlzLu6Fq2KndG5k36U2qhlpp4rPa7wKMh1lNwZxyQfM5kNTJ1TO27tUDRKH1Qh+
pBSMGgm5pNbf7PqlZ2tu0AQa4Y7Jal1FGYIswiH87MrKxXafEb1x+opckCFn93fOVGrHMh7fbcHQ
Py295qqgpXkrNd4sJTLCYiJXFzlIPdc6DiIm0k43v185T7Agklks9wG8oc7YxgBRSEwlQbkF90Xv
zyYR82C/4DckhvnIo9+o+daY1mC/8NOBVtAH85z3spZtjRsbq76OelW0cKRxOi0lcSH7UMEWiR1W
Zt0bTWNVOPngEnZxLe0uujMBCfacWI9bYpaeeSTJdu1xQZwiePDYq64DABk2qkGfD8dwv2lK1Q1y
efYVFg8vkKKaBwjtO+YTP9i7+Z9ohhOFiROq33LjIQadWCV83U4aYvT3829meQFYqI/V9wis5OAD
luBp5PDlNmKkVWQb71s8/L9kcplsNWNClZWbBlmDwWTCGA0pdB1c5NQG0SutUSxocINmnMQwWm4N
HQIjUDq2aFRff15oVhvJ740KZVXGC28Rt4tVYgeObsz6qTP3vjW6oipDqQCtVCbhtZ/3Y65Yw7sn
C7gzydKuK0e6yX3ARWMxta8sfO8TlU3iudOfOO2ueC6r4y3+CRPtKvzsBnRyGaogIGLUTS6BuId3
X8zyZDHlr6thkM8EIh2b0/puv2RG4vGhyFj7X/QHUpOtsdEUNScRlBAqz2tiXPytrXqiOyoMaYcQ
UCD5Y9WbG754gOkEf9ZJ+Qny1Te20ImF+ALOjW1AXxBKJQpfL0EZxXbMH/5RvJZCiWJTML2ZMTUC
wH79QcLu8zKU7jxUF3o1ktJ3KyhpURr0NduYja/i+5FA01MqtYAc8YF461rO1NzMbD5rzAG3Vkt1
YO4uo00Qsxdb9ipROcy5savDNLDsqVnLoRbmyRYBi5f/WpYLNDJxwzyc5mUH6ds7CcgTWPIFJn2b
vXAm4YV7EnsIxohVBEsOQLA5VWVHsjR/iZNnTmPP5S2p0I/3KiDzdsnpJwAFyzQIoRcxf7VXaidF
j1DTWrsDbYT2ltXMAbujjYOudBhunavTM/McDBFEiuvDkUIv85jj6v6y4+pn68R7V3ds4Ws5b957
+YD/YB3mbbnBOE5cFApHgq3YaNg4MSuGR7vXo6svKm6PJCHFq8HVUBBj+hCv9S3IdfWCegSoDoB6
254x0RTiI/01qzyibr11vOij5O2NzRRvGdLqGm5dGmVL4Kg632VJPQkg8rqas29YN83+m/NZu9Yz
G1G63/UTne94/Omb7czKEsPQwtSRjTfoIoj9iZEP8rSNHjm4ML+2qo50HbGJBYNhs4tOIXGNVukv
KPCxcOn8cIA3+YsLPD79HvNeUlqzi2PmFNpOs6FD59xPeeZXGxUpl5rwOuDinmXR2KEQBb/l+zH0
Hq8drODTgBxEf/nXG62KYAPmzOGkchthJtIiIPoFKCJcKffySILRVtGYa+VL+5iPU3LgQTNN4PKT
lo87qH2hrQ6X5sjGARsmDxJOY8DqcZO8MbsmbPfS5sGEOe8xRDz8tdMiLKifb9Y2QISe96C5F8os
h4ApMpD0lQA8nNp/3/PNaO65Fdz/I7rRNE9mYO44Vg3Xm3IO/KJ6NOXw7LRjlYXsAsn2zkDEfzuz
JFJty8KisuHWrt75FYQW7daDctXf6wGC12/nhXGC2NrOED2//baPb39tc7izyRRFFQrsjwohlnaQ
Xxn0g15apKEnorUX9lAB4uzyRxYrZZGWZbTyfGk3Dhl09EgZkQDIhzyJRiC9MRzK79QZE3YNz6QR
21edR+0u0KBdEbJ2oFhXZxWTdkexOsAmVdbNKZu+Rl5bGq2FmvGL6gHsnw2ibEhQUztKfOFz26Iy
VcK7iowE56R2Fqw6buQ62I3av6XBFK95gBMRzDjB5B71M/cJPbjKxW/hhFwcdp3fPwf452IkSBKb
q7JFIDMMDitawWTmzbn3XrcSYftx8hNGYReleKpj6Re0pcPXghRC2zzevDetqx1QzR1z5Rouarx3
PFj5y2hDxATMPa4XJ2GIVQFDbPnt2i5O0nrkB0b8p1ym6whpR9wfauzTC8j5lr7/KT776dCJtgR4
oYl5ELlYF1t950FbPRvwlUAFdGbohvm0VJJL5c5VfMEvGo8Ho3bqWHlHKNNU12F75+mgQQU1gIDH
+vEzxBDBmpQETC47KEYgHj4oDWj6i04nuxWxnnM8mVA1gLD+Pjv3xhNmdL4rrCiwZhJdfGd227bU
05whhkvT6cJuXOtmxAPQ1HDjhTl/9039Owo4L67cjo5y3gBsuZqm/70OQiDKVR8fZCRqY7nRel+X
hDLCn69ne2NPub7fGcEQgJnBm4PhIcD4/ZaIv1ykwWRTq7WON2eitopxlT/7ZtZTHII4iCmZGmZx
byyOkuwvIlc/I6FeVDDqVN5j7D5Fo0XHpDFRXOHdWUJS/BqWEUltXpCK8100wvONqrOVY2R3Vj/3
JE402oX7UrmHaf1WftHB8RudOTFUylC+2evmzsyVQBkv186yBQ3wvg500gBZSZfcIhMrpohH40IC
JQjPCVWiVHQHEKJZjssArnwfRjVfetyOfEjK/B6dU0PTBs7OnvqDANeOFRfCbx/xS0du7JUl9CXl
3IU541DvM+A9vfAH7qOuInSnwSPWeMjpCHCHxVB/lnkevcN6rR0ahUBZ264XPNKyYew+yt3daBkz
I1nhgyj+2IaBo9effuu6uDPpLfNk382SK73TSeC4+RqElB3MV4HQv90+36oEoqFg/itXkcmNQKF7
zh+QPu3iHH0jwSvyVZNcKoP1kKX3NDajcgdFihm7KlDVy6dt6EttaHD4ALuFPClKi9hWOdMRoIQB
t/5DZhTAJtz0LKez4FvwqHEZ09FqlDiHs/CK1o+anb6sWcWVe77ux35K2vix2PSHGH72o7OxefrX
9oYXgyWECD6LIdrzLyWp4ksSz9GnXWD+lh7gzBn8z2T6+WpRzqEgEkD2kDa4vgfsXuRN76V5EjU6
ogyD2vIcwUknFIM6uI1WmK49jKHC8TW3ltOU1UEXYcMyb137qc2NW8A83tfCoMvARXJxArxGrBm9
jGi0JVKPRCYIv4cetYN82YDVOapdNAHUMKT9gsgox0g+fpnyFCagMQAbGDP27oVB4YtkwToQ/KJ9
PtmbHAvbGiCfuaRs6k7leybw5ADASFDBIHnM3SBdSzgoUlOdOkvnrT5UURRfeFuFaXqxiKKvCn7T
FNI0Y5x8RcHNd/7Y2yWCZjbDi2xhqm49IkuzRrEionYDiN0brFg/gda05coMPGin5sYjmbs4OFnx
iTAsTvWv6E6499J/JboXYQhp34P3lszLbD3gBpQqHxb0hN3Zj8y/+mLUlk7moPTgI38A4FifVIgc
zeA28Ia6/FLmO8HINtglTqM0lUGy4LICx+bX2UwnTYXPPFAillmRKifRRrPE30K19KrVVuKgaBrg
We9TT84ny/8IXaX0bwvgDpu0rg3TS+HH/c3tNOEq6ewH8LKI5dtm6sKzUQCxrikKmWlSs+2B7baD
D6e4dZDTQwh+iVAeJs1vW+UWnzHEOOiIZcNikd/aPFVjXsKeEk21LAHnxwnplTQ2/GBdg3AGOSSr
TUNg19nwiDD8cBBK19dR9B+40+JxVlHNpOKzQvlOUx8b+A7NfArl4eJE4rRfH6s73QobDkjZxe3h
XT4qn+cc47+gqpp2Xv4jh+VVaEV0ij0SPwUKHU9DEPn7jCIcubeSSTgcGtfJdZx39IvvCgDR6ARQ
pGOF+ydjuSo+GFPkhnK5o+vj5qvg1qGi+wq4WlboYHDzThzw01rBC/KkJEVwpW48nu00vq0a6J/w
0Qx/QcvF2X0qT+kKaj85ZItQECWMXnIINKyaRY/14WX5UxM7FREJ5sOanMzgnbC5SHPGMRCt39Bp
eL5EqBQhqBbmXrm0ORNwmKuzZxUEItJZyuwVmz9ZyYuTDfaddQYwDpkDmncZ46UrrT7PASf/eNRH
p4EsEieflb3vR3SL7qlpD5b/ujj3aX+Dxn+P5vk3sTXumXYgAWmTCeCWzudP7qsQ7bESUBkuf9ts
4Guy57buK4rNxtxuHC9IRztVPFMxA6DxHKQHj7j3R+VaeytStFAVWW65NXM6ioJzLDH3En5YQBil
YswLKBHUZUtRFd9c8LQauWVZ5PlAQfsbULS8PqleOn2yMJ0VqAMkEO2znpTvVUe9C/4baey/Hcf/
BNtDeGKRHsdagUZvYxzF0xorlGaOababu8lvceqDg3J4s/mL8fdvn+6k6lxdlnsNLEnO6vHNeevI
4nb5nEV/gLjNslwX9sLul4r6BkHMeaSw7HjHeIS29sIsIWYPbmwx5UU17RoimoHjVsEZKvzumBTa
6IT8pf5A5rCxVYdglixdPDB+xcj56z7RKSW348v+R6ZLnbMVI2yxdU4aeHG1UGUbhM5n0LTlL73C
kYCGrII595QcgraQIWjBhWgU7p4uDWrZVCxx4mtB1Tf7fVaCVp5g9iuzXjFwKTFqX1VQrtTyFB42
2rLM+XFMrt8lL/hbmoQ80QIs4zcVfs6fXqr9TnzoXvj7w7I4afNI8jUPTbcxLwXMjvgpyHlqQZfC
/z2BOpxbIET9fRcdUe4TWWNjnlTImxaIheZdsfFcv6bzDvf897QjcwHVdBdoVVJSt3khmlcAufZG
FCQyhePhhEkSn3WSfQjAd4twnHhvOHsI0irMrqTkKr9E8cztaoUohYaspmbqn134f2z6TRHk/BR3
bIS0urMrylvpC0y1vsPbuQ4Wnu8sctZvjgq63cOLBdgVYke4VyQ1DazcITLUOHaAS6mWY9u8NsBq
HNK148LduQMnAA7+XLHqDVQcakQJxHeIpLu/jgu8ODmCHUYki9qywZPs1awyCaHR3UMI2aNzgXjR
44w4GcDCr42de9fgkAwIooGS/hNTXZf5o8zDJB+keSh2T4pRD2ey0xO0JAPzq7SCkTVEQbhrIV49
CE0l+9JsdUY/joVMYIE2NpikiE+aA+iF8HExyUiMXUdRTeGBttOxDLixvATACaR0yHx53dynxdHM
rSY71/q6xLGPnGdvXSLfEyunj1yXmt3CSJEjPopPiiUXbDkbjGUV13oV63DIUt+c5KsnL0Glwegs
4bm5lpahAxIqvZEij2grs9FOiFuT8fPLn+WkaxKTGxB9Bi6K/gvHRPZka15LzI45OWS+jaWVffY+
ymTZw/mOSF2ieCU6/87HJBE3P0iG54ZDuK9g8trb2EzxqmwjvZo0+oh3NnbY5TmxmY3CW/yG8xoY
X2wvw/PJ+qTagGakNzFY7g4MNPxu+/BEO9ly9xg6rPvNr1dfyarR6YMP6zCgdgzHCbPxyQYwJ0P1
EL5WwZEM5UIs77YcFBMnnZLlTmUMJ1oFTgUkG9GjEqal9SAkO//lRiQDnm8dRQI8dM4/Cld4w+b8
8yqsr5Z3TzVjebmqI7Fpr/841RN9TLUuVVHWkI44As2bITFqDlaMwHEKqCdCZNujrwgcFYZs36mh
qoZYkzF0sVe+TF8dXFZ1MOXPOZ7qnG1aF2Z9sMwUBobuoTmJqH2Q33DAjVD/cYcrf+hTOc3zEqkJ
vpow6+HqPeAuFKlphbpaQjB7DYyTfyee7wgzLTVEMhypY+JHQNv5IoJqmH5hxHBHVKJzgtuKkGog
JjfUkTvutFUjM9sCWkx85WPo9cb2kPjuXxRtfk4qKfds5sP/pzJpShmyS3C35p4Yx7CeCIEJfgal
PYQNOxCeHNgJpe/486pAVyDIcB5nGBrfxLKXuRZRxTB5PfWgqBpRAJzeCVQAhvre5vNPifltyqhM
W1cjVzfxFK0atm4X32dVUhu9N/OkBu4M2GkMy334kF/m9tLGJxiRcdcoI3Hyf6KnxDN2mNllC1cq
Pps3+QyjeBCFg+M/RVG6n/DWOHYQyqtaCRLHb4+u2d9RuWyZOZp2WSQ02Q0NGYJLtEDq3zPU5fCQ
X7fKhQ0ej3JRIRyRrI6I0MjsQ3DDqKPnqfK+1myUZGfNCLIngMwb4AMzedko4d6gwLa97h1lBrqo
L1DDW6CFdAhvp62RPZxIIncZVIcuIQpHh73nBOjxfjCEoGJFPa6UYeWIq5taL7KzdgfYseEjPd8e
IbBXm44wV1J5BQlck0jVZhQ0req3LWtR54E6UHDvbCvMV7MOn8A07k7xCLzeHZmb+Mvwt6rzo5v/
nVfOQC/CC7ga3rMz31cVVdFdd2nAud6Ithqv2vqDV+GxbkAPFQoJC4sQy/AA+5d/WrA9zYqU1mra
SijVDdEHKlASREebahW3n7FI1qmWmn4VbXM5h2+AjU6ClttlOTGBPHWaZf/am1DM8CG0y0SAGyDy
itSaFkyqluV9QnIuRz82nPVVekxdd4XIj0Yt2SQRk+ckhjnnP5dn9GcaII36uX8usG/Y1JOwXvwb
suR6phqio3Hqs5xp1Cr2l4Lw0hT2oGVR5TSJjZQi9ieBI7gic5KN7g1iITua0Zaow2pApnXIFekg
u4PIo6dWX7EiZ261xv2KA4QDWD1aCsX43zoVx1nCiELhzVa+Af/Q6A9yUPdzVlbCLU6jbtgzN34z
8PvcISdb5EVpeMcjJcH22qPvnPdHRiCLw48cKygABR+WXTPy/cpftOONWd0aeD0ZmXdFtoIsn7Xs
LAR6pdhRT5IarQFeJnBbKJyyeCq7pOI3qbhG68xtAInxkxcy2dTTjJGIfmbWAz3QY5e3AavwQaFj
cg3p5t9onWxD+m1PnfR0GMIguwydBUPk6wwhGfa/+iIRDdC6Pz51cxcm0W3PfPV8iJvVoqrMI7so
NbrIaoSRlC1EzcIoQL01jCJtWBlx42eq4HAHYYGlizlbz8iYeixHmPj75QrSfPbtXVrXtBf6CGdR
/vDLgpwtDx/sY0vGMUHPnEiDhgn/wdZ1UeUDYB2bEcQ2XHNL9Yq2v1gazvFEAJ4gJWSxzhssv4xv
6LAGsQNUU0uNSJ65yfKz6kS44CcVxGZClCu+warZ30ZpR+DAwU/JtmkkJXeSag2dadVDWKOgGBG+
Aw089dz1gq2IFnKNuy37pB/Rj2S0FiC8kUKccCu8SI+HLTXp0M1BslzLceM/iLzbL+DaFsTSdZsT
AfNr/sHYBwjeQNpkJJTgPnEvIcHN6a66WztQ10KU/Cr8u47YUUI2l+quMO5wXBDmmxNUa3Fyrm9T
OZ7ispWD9e7qRLtGpV9QmtxAFPkVdoR/BtJ/SXc8T3NDCwT2ikVTZ+ZKdl84uMZJcAzeht4msmd3
cME4voWgE7PtjIIuQY8DYC2eYi8qwyjc4cphXRhvkRLioEunOwqOxafW3mc0sTc1RsaKICJLBI1I
PiJm2s2Uhh191snzq+4M2w0A0A6qZb7lvo3Q0P/3G/WziyWTQFlhWZsORLAqjZ3Qq+UxRbj9EXfY
qksmM57g9Xxxf/4UikdbdD3wYIvaABtEtlebpO2dzXq1BLoanmbmCrN55+zOn4d5rYYljnNvuxDY
sdLOXxBVZuU5wxYBb/OKPAfbpV8xahh35d0/othuW/FrFm95z1bpJwD1TVPpWty8/u247mAx35Y+
bSIrrfg6Y+KzY8xyUiikACwvNufKiq+fzLF3+kU1puptXIUoYdz3PhPiufUcax7hsOaW5T0v4+6f
dMDN/hBOsln+IYjI0vRPmz8ZsfmimkclaXEVM/3n9zuu/OPFPh9In7k3lG54eFNd0wdTTGDD3R1a
qsFQtv5Is1EcmLr8sTDNu0SvcI2Ui7BjRLjGnGqxsKxEzmAhTEOPBIbB7eg5cRYQGK2JjkwAriwX
/j7hcNZO+Q7wu/xyEJ4o3ph3Hc2q8UHER9HVBcOqhyZnmO34IAQ26WIaWxfVg7poMt9cWMvxPr9r
uLQzkL8CG8e12Xhcc12qPO7xgAPesnmobcjFMy3bcZ7eTVaCgqUFKMvfXrBAq+q6Y4dFxeDlYNTW
B4v1twoFgZvE4BAPOOKcDK6xbmaoWbQjK+bLyILxiMsfeM6wbZ57DBBoFTrPmmcwMSGCNyEU+GfV
yzxu2E0pkCvpZv2nVkWfWXyXW2MA7cNpbLwK9mfin/iaqh1hEL84SCaEa9Uh5HN594kU8iuHPMX6
kqIcNXnDQKslk5+RieIpufrUwM5KQTUFm8OExB1SQhLpD44IkMGuWGvNZYfanYCAHnZrNg1Y8iYD
iA3oC22ujgYeP5XOzW7X1a9cIZLNcScIzWZSbplE8RL/3vA1zNaIrMyZ7A5UGybAIeDmmtUCjrUQ
WdkGli3HvOzsukmbC0OAwNHYcFmQw+Qi5m0LpWb+IW6208+ETlSgAeZdJ0L/KaGHwo8nOKBy/SWl
Tc+OFfHHDN5+9RjuKG7jNZVsPSktCq9zJ/wZsXu4hovP+wflwVHRlTzajAq7MGiyMAIZn4vpr1tZ
aFWxfvxw+0GStrsy8UM6ZKFuZRtb71edAzePQahFVt22As9d60OQuxDLnTUTeOvGZ2SrpR4GET2L
aWiusFhsZiaWZuBrbZPUGaS2UPxetwKH3iIo+7nUSSkHquoFsVkZD2ZoNPN00W2gT1AY6xlCFDaN
E5ghpC79BW4b8PUyF2pV+sbWlQ/L3r9vwEU2TPzQ6mFs7ApEoKhmJ1CQKD0qmELxgm2XrgMJsbjf
93ZD1qNEnVWAne9UqWL8UF1NLyV9mMZcUGrWg4biFpVlwe4YWi1xW48X4uEQ/rQ2hyR8NcRNPjMe
OhrSzvqEyXbeHwPQFf2qG/gNTPHkjTjD9vsot5lUFn6XDl3AyzX/soaO+r2Xe+7x/hmj1iH6UiMt
iaEVcSrwI/rawdXbhyvbSCspMLlev7fBsmJ7Yge1oEb77EE3tL2dONlu5Nq0/lF2DqpJkh3ODSik
UFiEcHEx6juHJL+E0Q0x9stloExUBoq2zgfyaST4AQBO4fBTbx8MdCeEjU+vlOYrk5HcYLi4GKGc
wnxFCA0RmKomdQu4+TzmD9evB1vY2zCLbKxC+BkOcZdUnEPn5OcjdJjaqyvBZh5KLF/9CrILbyxo
QYQMHb5n56hh7XFTHIuY2fEVIJd/tJntGU+/HzPdKDV2F/Uy943ApWNqNn/aKLRqeWXxJC8FszUg
ZPy/tqFuZ7+4ZW78eVSodv5gwNthUjWDmbzr+K7XSeoreomwYvkSHWFXlFU9xLt+38K+2zdUVHJQ
CvbELlPp0sWyu0NpfEzaVCoY/mYHbH8foRs13RqUCL9TkIbD7gBL1XkiJNOOXKT2H0qk1pSTwC+O
NI531HsqY+6/Lizymi+xNAaJl9cvoeGKq1FGYbDkojALBGznnszIMLrygFwoXi8zdtV+fx7Gt3oQ
E09MstDakzMwfmFiLw8Mgh95t3q/ju8cyegvkcVMOL3gp5gBJH5LAuy6+U7nM8hjoUKWjUz4BSl7
NUKb9PIeq/VifEpRzSqCDeE+WNOKaz5p8d1fU4Er7Lp8O/1r18CGLce6C97+XLct1ZRdYQ3s0N3Z
FHJx/+SxG50LR4TOsVDftIYFxWI7sclgyi4pXOSPnvljR4KvekFMmHfb4+gh3s0tm+4ndMEj4k/1
n4H+odbnO/1dbVLefpzmPgeG2gBWawxf/dWmMAnb6ICx1+oVyU7D24AjL/gb394iv6vWAeie/WgG
CtxNkYN2Og1niybKzpZpzUe2Ow53p8EPNQhhRTtHdtEd4VWvbMRznASNThZNrI4ZP1njXCiV3Luf
73BvjDRetXkmJlqeNx3GI8NYYNXtA/FXa0qpdP2qGQ/UFiDVpwB9J8uwPAF/SgWoZBSdr6MfvQ4J
f0byvSznqSYfA5PMEHKrI3gaKQEEc4+SE9vdeSzpSnbTOKAWyfOGFvPCEtzeOsFhmc0Y8rpDZ/2I
lTRlojK4BA7toig2d8S9XkpKWEH/AR/EzBw/YBE+RbflVdxGbaNoofB1ALTcVKSkbo7E8O3YuJuJ
htv0+lUC7MlWfM5QHlnO8lUam1EKvhxENxe9Abl09/xEeOThFa9txO2xp7qbmjgbdQJ3L/5xKIuA
VM38Trt+JPO8mDBkYABEl7KxjumEKQTpMasVFpCVZ2M7gUJESXd4wJ8A/uogulXo6D4xTtBqOL3/
kH5Chaj+C5JdflHfNmzFsUMK+LTnL/mbduGBqjp47J0rVx4mNnOPxs8elscogTCs99jGnMcLBu9R
I+F1rO+Es3Uo3Mg0dj2u5YbyCx22DbxbHmHxJaqFSY9NGCO00Gxb07F4VDhd61435/14AfdeHkyt
+WKfRw4sSYAKA4pi6nMwpKdkI5psQIneT5GWGa7Em6v0QR/pGrNTVFvLNicgwR/ID4n2Hr6mVj4y
aI7Hi2dJzfA4sVzGUrr3az9x/X16nv4cY9q7pvLT2PW1YsYHAdt4DmhopDkJCqqDVT48kr96dTwt
rlIBVOnGcR7aTzC0KDSxpBD9ENFv3pB6dR8fiSopDnrtszMTld5oj1UgwwN2+ZxoasmN+9CgmFbU
9RZ13MUhYUOjVAw0tvr8bykka6xPNJBWfTGosW9iMwXMFiloxpL7vcXr/QCG9UBe3TNanke60B+m
WSzS9pueQs5+N0B37Sh2LgQoyQm4tUVfcmvDTVRViP4az2YxLgHkZ0XvdtPr2VCzWRehnY5xr94V
1vw9iD/Q2SiDtxS0avnmI5qdHVDvriYggKRVh2DaKini3YgidwxEJ8BzipYPzTE8/svMmUvCjYiA
F6pf7SjpK9Iq+KRVgnYzcRWA8QvMN1h0jH6KuzbD9CiucHQkZjb7SRPqUFz00UHLOBPm2ahKuLqY
SjOdp+BhejAoJjqRbrCs9ZqkxW1/td0TTOGRx8DOjhHBnGQ+sDu3X600s6VStmBr6d4spUs9hZV0
phYPIpZuWz+l2qFxuSv8hlzf6cKn6ZwahU6V46N4rJZEReAhYe4hM8x4p8fOM2mE0njIl+4BI5bc
YNWaP9v1OKuDds3gsru+VIHGdI9nULpypiyyXBQGIOMBBs1xOZldYNmYVMJ7lz1fk+HcbugFhivn
qLDQ3umSFaHiT/C6TpTU/tsmGeQSGCMptSuauGLX4L+hYm20WWw42qXWOhEDmyyr7fhK7OIru2E7
m7DGT5+l9RDcBrxm+x2isDi1W+hB29lvObTdAHriB9NK3H2lt1x/eYdfL7L1jOqPJ9WobQqQ2igg
ak87Z0zX4KGrOwDpYok14yNH9oH59TBXgoxuxZg0J+8m+zwrA4U9oj4c4KRZxndG1S5i6lN6rrZe
aonyasLDe7VY4A9qKoLzukPgu/DY7e0HQRsPM2X2Xdha57HBj3T9QUy38c4WxjtsfVvdO7ZPUUSd
b8PuYTh8U/qtfzVrLOwfIBpiPzFdynLGWr2XZLdmSZNoIu2soDbZ5zXUSBawLAwjM793JxuSEWM+
A4RZTNUysQ4Mh6kqo1h8V7wrrawbpKOyVXbs0UBs+aFvcqfO9r8ge5Gl2aNir1+wZus/FOLtfrcs
bZ5FlwoMEKVnhY33A7OVRyWI8QSJCPKtoUTggQDXdk9BqNNdlHVuICukZhNaJyDeVmCH8cHOLvdJ
/q6floGIJYPt0nxniG767fwKbP6s0SSvf8KWyxGKjWy9ssPHDiJF1ygsMiYrgy9kfRWY3EWGPTW7
fc4ixlUPrcE9RuN8ycwsIoKZqGjJ+ZuJCDjs2KTklfQtZbpL5gwSp6tYOit2OzWTX8a1DglaivIN
canxky611kGYgN4AhS1bfE2oErjmiZhTF7Pp+psYerFYXcAL4XfEEB0F9/k5s2l6nJsYD/qAC29y
w1iUSSTqrPlSOwnuYqOlvRVccAp0SGHQ2qrsZVgsHqvsIZcy8d9GBosS5iS1kdMhND0d7UcyPOax
g+DA/zHHfvJoEYMATnw7cyGWaRa/6AE049Bbs9kIVi2Y7ZfrEUqXtedyEn2YWeMd1uwktdJvgrva
xu1Jjywr5vvit+BAN8yChue9wC+WNiHeF+oURHtvHEx1v5oJQCNVm+ee6RBk4kibX4To9vITbGl+
1Qj6HFLPz9kf93bArv4+5/0o1gxCjxHDdITgCKASGXJMJ9gouChIRX/lHg5fx0o+UIiiboqZhnBZ
tVHc4r/vN+lr6hepMqHjG2omsIMmZrYbst/3vPGNe1UXnh1vA8CgjfQOj1by19HZd+Jj0sIhD2DZ
nM9ZsGsWss/sfX+Q6PwkcTrW2gB676MvpxR1nH9jZ9GnecN7r6gYbywnatwdisaPgFhhDJ0VnwTs
gdeD5LwoD7r3iJgVOk0TRFQ7IH/ECJxGcgHzwR8HOR7ScZaEn/tYoKYo8KshaFdZ7BkMOXn0IVAn
VwDeKPWHWvxCNB3E5Qbm/L6Majj61NomK2be8XGQXIoifMqErgJaQBYUP6uWQGVx0Vs4g6gZ+9KS
BestvbF3QE5GRbPq2W6oS7ObkyHhb+1nYNAEXi8uSEytghsg3PIyd1f8f5/cB90+QBLh3NsJMyNE
FZjN+Niu7bi83m4HbJhX2wVpAU/SQ58GI3vteeP+ua73IyvrX3PglLzRRQ0s0Z0d5xQmA8J4fR64
rYXKKaCyqSq+dQvwKgNVrRFQNgAY1U5ORj51l1py5rWfvwRQXan59JjICEOwIY9QVTVkMu44DVVs
1UXl8tdph68IWw3ED/zPFrUcOHo9wJiqsRUacJs/v56hd+rTHMxF+O33EAKG7E+MK9v0ri9xZuzP
/8R5A4COTjpeLbk9GD7HOncJpsYQj9oHxKAeLYFbZWEeCV+wfdou2+Q75wdnt1mfZIDiOzj/majT
PPirvHfoURVzTpkkhsgNo2cJHCoMJpTBpLOnSC9jaUU4YKwnyr4/FLmP4CYyQX20tfTbr75EYbH5
czDD9ku9xDvWC6N4ZUdYNS0JLmlugBH8kn+BYsuTGnjzT08TwMa7WdaAv/OXbRY+apEcuJ+aDUmz
lFflfRNolV9wCJkTEx7s2bmT2NtjzilrPKOIOZkBfkdGMLTOMIDs759eeqb6URmCspa9LQmxDkEy
w0oRBwS1EcIrPRQN2L0/S/qliYvYJWOeZuDYwGhmvcqo1BBdM7KhAeaJfzGkB6GFv6NLM2ziot95
0k1iuVTHvD0LFLweVsL6dhl5JigWWNHIpUQ7/ZOlP7WyYDcUOW92py2hVY4eZnMdSllaCLU6yppG
w2txy0jPkmzMtoBvnUx2PFVs6d7z1ELoyw4i/j37C+ipmXWe62CpdWaaxDAKsP9FoYkkahUUe5O7
d90ASZODs7BdUoevLtabXbNInWg9h6dY0b4YXzGetb/ozB7VXCp8pM+uQMjkeuP0WbqM8I6LzIMa
Pb/BppnGHXQNk0Lj1WZBxinFal+QQGuenHx6ZhVv5nW9j9fhNDxxq+jJy0Pl7rDTBc/IHFEKBtER
4ghWJaJo6kjprrNoim+uS0aZ3mDY8mH1C9/c+Y9/R7bwcdc7blPNrxy8vG856MYbJ/JxB58VLY0E
zEfV5v38OQ+GcEfycPu4UblCtNubJPTOwHeUgGfZ+yLwZ98t+tiksG1+HAXEo7eGa4FIlwh15STo
Nr2Ffs3wjUGFD3ielVdZvv7I5Rn4uzdFCNeNOrtjG1EF8qcKZ7ba8UIFp8+/cQY3cUcggczilQ21
8KmHjepnuZb92ZrEFeST4DU/Rd1oL1Ibd9BrvZocnfpt79IG1aegzfbOpQrllmb/wEwLJQjFT/q4
Ou6APFjFWXx4zqtPmrMd70y+mmAn3gR6NLg7b3OszxU1N1i1/aTSJL2U8xNxiDY//JdAgHRI6Hgz
OoKqHS9PctkroZQQLWxLENsdgB5YPW8DMNYboiXT2354DoXIvuKBlp8banbCCL0UXMNTOCLJ2Pbw
+LtVtWnrmxpB3mhBdo+HMcYxehRkkRyJWkiNDnUhdDdZr1oIjmc4Ndy0tKBS9Gzsf1vBRR+R5Up6
AFpvx0AS49slrejSDe46cGRl/TX05TVreMazRtX/04pNxUPYiC/l+Vj0mNMZJUNqX0FiJnmRIx6t
6r/Se4gYqjtBGCVE/0lmgEPKL26f1uLrh1Mn7832kMVih6xVC5knmFPyGxBqS9ZcrUUVlsBEmHBG
j8rgmq9zOiPJkoBZk+NBfASiRWYudMEdtFFqfMmaneSbKpSruQ69fbMcWdODp+Bcbh0VetvO/ESg
ypl/RnXZQBtqB40RaWjXtFq6TxYJxSDTxpbF4rE16JjunweoEajvJbf8THCWNXX+wYoH5boWNp45
H0XLy/pyWYXJ5EtPZWJaOR/RZc3Pa7PmpLutirUPCDdy/xhvoJrLfWAyQynKd+oI94VAIAsdqITj
FPRhWMcETdmcXJXQupLcwSzOXIFR9+4snmy0Va+ROInrBqcqNbu5hsPQ8t2Jo+gnmZbTU1YLKAf5
tgLfGp2EW6g53goy1vkvZwzJl4CznhQqCXJc8CYtHedQirwK+uIBys8fyii/cn+yTHjHWhHbxQ9y
7Jtz+sxlNmDTi2kL15xLEnUXlapeeryBlBvpSpEQfEqlZ8czU7MeWvhAZyFjUgD/v0l/DsUmjm7D
qjUOtBAeC/eve3hs6RRPbHmu3qSm5F6wECEGKJIRmV2KqfSSFD9yq/497Yb6ClD3Ib9XCckK71rh
3xXUuBmts3sudChJTCWuHp0wJAWu0S/o2muRhm1Yoo8N+d36Obph+ePxsxVaVYMAA9kE+rQ6ac4x
ysHXAb2RMSElQ4gu9kkkngRUiN0Y7TliQRdAsqNf7qK3/vZKMdZGowEfZUJfTSw726Yr0wtG1ybL
6TGS9M3sOxIqiEdTZOUfzFnO9Mbfc6yxR390BRmQKofQTNHZL2l1i6Self/4kcJTEK3gZY4FLsMy
7idcP8Dt8sQocdxxU3yUQTP5CIO/aFG0CSVLyaZz0Rgo1/ysOSB7jw9pnmRfSLi2vZM4Dsjlqdhs
LRSCXwT6+TpBI27b8NDOutCDxkorr4CeQ0jbUeZZ+0bSx7anisc2nNPV0BUNrq7TrZgA2v+v7Gbt
PvUXY+v3IXoT2ULOW3drKevqkp7/jVc1VCr6RDK8Ny8UY4CjGmEq67cRCb6++62PaXzb6zjB35Bd
66d2bRDmni4wALqEabfrYBQN/HF7qr0RssgZIeJiqB+l61Jof0QodFY7GbhXiU86/RnSWgI8U0QP
d0aKnoqNbLYg53vGfKRenPAsAn04UKrKVmHZd1jlh7Qk/lIyZV8lx7jlULdE1wd8abO6Mk51CEGI
nqsYqoY2qcfC1yfkdcr2rGNJ4D8swVm9irkNDQC1tF/6lneAkGb073SVHKCQqcrL6hWNi8/n4qXH
y21mrk9OdHNKykvxA774XWhTidXpV6TQwggqerEK/DVIqA0hHVhawzUKXrAkwkUdP6DtXIi4V2WY
NFCDixlJRzb7MLPo3TBe9zhSw42PaxsVJDMkqacypDbEbmLUkUgJzyWeP+DuUNIZclkVYi6OkSdC
Myd60lspC7T2pCLCxvW0pz4Z14JQEvYzwlSRKL15IQlndT26GIrgxdSnD81gXFO1dlAIYqAkuFnf
AmkLUt6xyMJKnjXt+xR6sgn0iAKGRPj+wlsZoLNoW9fJADoOMV6KwSUKP95iD/3qPT/BFpaJTJq4
GOIMmHL+X7WrTWJal6f4mMaGHiWbZpVEW/Z9W9KmfRbORKBXEXqMXHFQu3DtPcOuSLMt+qxToOf1
jpzH9Uso9Qf18IHbTlEgGvwON2VMi8RVMxgZx3R1Q4J6pEwxr0E6NKIvouzIoSrKx5CLYUFUn9Bu
RTbDNWOJbi3llXjGN3M41T03l8D1wim/sifiWeeVwKGIFy2Oq29g5sbdX4+Ooyc772xfaangAGzb
eLyH0OGCk5LqutIqOFg+NfaXj/kbxz3GHBdneeEFtjKc5xLruhuCEvr2rAjl6ysdi6LIfEy+bzdt
MpWhnKb8sHr184dPBh093IkidU5Sk+4uVWAUm/h4bnlCmE0XZUb2JkRsiuNthefJ+v/0dCQ1UEmF
9rla4ericjzC1uarP5tV+XjrHJyATM5fNMsFowLE7CpfGUwOZ2AGz8rNl+9lt8OjQeWnSvHLuPsB
QeTUpiHyP7KtrNCO3IE02NI3Ij0DNsEiP71hZ2MVmDbtgD/0dlPLvX4RkoLG/dnUcESdBhWRYrpq
tVxOnVZxx+BniYvEJYq51YmXwOtcws/1Hv7Jmb+whf93suREgniX8NApeKy1aeKG7yQ25COwyw5S
xvtuq7f5GL03QlIN/cxZKbny+eibcEOd0+sGThhhBek4fOdX7GLZxTEwge+LFtcFkbfwLrY9lHMV
XAF97pZ8FBR9XZGtB0lFL1EJa6UHOPuKdrJSEv0SXbtWWX4KJh0SvIyIAgMjMd91mH8M+T1uSybD
q2+W4tnCoksTzVXWup1V2IwA3TNUFkpeJ52kCwV9z/269VZ7Gz4rmWxWoCnYhBBTRpcPFEdqwB58
Gt/vLrcdcNgRYdPiuZk6U/JA6NJ9bNgYPxwTckA+8CB7aZDrkE4xjzFuTSJuiEi8pjw4ZZXUnGjz
e61kchLytdh4nOt0Km4OgBxw9TgqXXO/c5t8NW1Zhqvdx7INEdLMFtWSQinfNmHhDDofDmxNecQq
gdqi9t3dA6TD/fYY93/Go7B1g20bl2dusjfWkA9072usIe7LXYWHxMjm6ZRiLxjoh9WBuidoETIU
KmAZqjefUcMqEIvVVtso3MJ0TKWYLUS9VulaiE4+AKu0uXFnj6opMCPo48f3zZYm1RXO05RImups
cnWCyAezvYNdFdqnuJ+6hbluhTJSnU76rJ7B/6JTgNucCqqh4DUxFJ8L/zJfKiYrdIwTiNAI/49K
H0HyED5K/WoVygoSC/xZNwZ7qLKjht5vMd+EEsL98aDasVUL7+YegwvCXHpd+Y1kDv7KGSH5HL/6
Zifj2DsbZJXTjxHcXcZnwgaLj9KuTw8LVR9opjyzG271WPmqCiyDR/GfQ00KEAfqQ0YtzR+Q2S4Z
BhW1R9BAnS148gjqhRaR4pYafBCfoFYwR8GSdVGeqo0Fg8YefMI59Tyv47WcycOkEeaREJUJ638r
X9S21EY2Fu0w32a4Q7q3Z5GwSD4OZhK40H3IFcr2RUZeG4MqwOy8r1smfTrEztDkb3F4nXIkKzvM
Y8MaZNZFxbT2bglvt8qoEYkmyV16eotyvajK3vL9WUsZiu8OMipXadWW0r1o5DnR/5O/lblqSGYA
1IN30/p4+Kt5UHsqluq8w/EV7uOO6Bkz5Y1jiOURrOJPP+d70icy53TyHoCrSfSBrSCncveyzsyp
inAjfrnjK3G0R0vjE3Mn8h+gYEEHsWTFfzAquRh6XZ4FvdMmQV7Vm5Ops/4jU8kuskpq751hEt7T
AxsyI22W3bnAPFe7/UfpB47ikgYY+2VIyh+B89wKgFNTF5yomyYLq7ke1ZXzfyXvP7UOp/ioa+/z
wjWz20gqxANtyt0MzC9i4O18/RyClUl4nsKmOeI+lsKK3dnxPA+D2WjkZHO9U1B9qQ3RdGCvtDcw
igbMKPzK6YTCRzdAsVVD4MUBe3amCW0IW+ivGevfvzSsRw0OA1eqsOKjkN3PPtZ4B09lLyPkINrd
epC/M4JYd1Fm8bNRMeCVr2gQ/CBQfhUbpit8RGRJeilFX4uQcUvbz1I2BRc8usreSEW/jNrzRVay
8ni8c4cVX854CH83ivR6uQX92EwrCdoB0wOTzwMDWN7RTjiBtF49r4LGKiBjlMErE3QXSW/Np/6M
NwH7xhNuCzQALB3vjt+nlLHl3QVXMLcl6p+2jxnxXag4MlmZGPQucndMdsq76y5G6qcJnu0BAY89
8X/BopwSteg/Va9K8T76dX3HPtNxP/N2yJcCFi64qmS/9yjOHEVrHgS7ezHK++ORaeky9YyT2l69
8E/c93MimpkrZ8YSVPgwzkuLq9n4aKrcXH5s4LXLBUqWkjFx0xT5yv09rp5u6wBz1I+9N+SaizdW
QanfIC4deVmYtAC1+lMGJId97StcXHOI7xw0fbd2uKyHnSRZgZrnZfzkT1zv6HP3qbAFTbrnMAgf
O9PP5xtTeTq624jTooT93J2Y1PkBfz2rwvfJhyXs54VW3BriupPLIFBw7jpqxxSPy8Q8qRvbqPyP
KlBNriWUiS2z6DBLc823ZOSFzhL+etuk88ZihYUJlLoFwMpCh/Nly7zlCRxR8VxS0rLxi0uHwaHe
jFwlBgqk0TBz3Vj1SG/zQ2nAQnkcbjrydJDJDerBkWbmzRTsIYIBykT3eeIHitfmUh+S0IkuxNE7
GSMbsYNhr3qSxXZuOcIhlxHhyztwNCiCCaOZVo2NEhGulZgv5DXGAXkusKNOwe8a9OB4eW4R1gku
X9fAJjMivS9LNl5QBpZLpouI01dmEohnsNOW8AOnCP/BZezCuqCzvIZwknuSRGPXH/tVJSn4nWK0
9+ZYwrHtALR0OVq5BZ8IvmBeenjcZkVmrMxd3HaSXZXzsYAY6+G0eJbb7Uk0/5sKnmDRWRj85YeM
jIK/j+FzoSo/yIViFpmNPrDm0/gVHk1vdPtgXulhw+9OpuSlz6hHe5N70ycvU59Tj8L3zJqu3iC8
I2oDqSKDN9Y2rA5n+xrFES9cki7TK/l5IW2W6hWWGwtYi4nGNG29R7N3+uEla9z53hxzOOlQu+CO
hgzt8zzcFYQX6bl5elfMLjqmOWKcmTb9+ZwoHfQ0x4yqbyvOPPtCpjk6D5krYTGd2gIGL66ghJgN
fNVoymf9629mEO5TwdHsSkLbx3JMqo/AJiCtm/P9QnnvA+g6eR0Wy0HqWkSW8z6xgCHXVpAyW3hI
XVd4nmXlha2TUG9CWjWp6T1qqt+Y1sVeRMOtNPyDdIzFzVv49o7yfc2/JfCZxS4TBKKwJXj68crR
WW2Jjj6KF8stIDGbaYMbJWwUI/h/sEFIFTqtlDSR/WZbDzomwrIm/86GtjDVs8lbhUb80v/aYr9/
qrRAdY0NmyoxnlS2RcvKnJRIAfFYQhvzSin9fdL/HoQXb/PLPmYLiZSvyX1H1BtLvDv2ZiqMUNGm
2gNkbpdCK0P2vX95N6WlG1br9MQB4EafsPVxbR1pUA/KBIt6TIarjiywf/8M2Ye7RN6/R6/Hw/8p
6JGFKu/KH5GjGDWyhryw9C1ZplSlj8FOV7htHRinK/n3yoxOsQjK+SpbUIPnWG0v+MblSTELPDRr
ZiT/lKvQZIwzyYigg8omkFC1wmeS+dUqV8TBbJ2qYFVmiI4S/lfEf7OtQ8cz9vdtOnzEhC9Gd70c
cfzVJHsylX+2mtRQRXtgRiDqluMEO+dqWAbYA6DGoVMEDWjqEJDvG8G7NYtmlW8YK6y7DOFN1buZ
Zf4wn+ET5FUBDOIUbGcO5bdk0oQraBnArKwV1rzc6WGdgMc6mJeHlywlzQoeBzHUjYbXm39110I0
3Td7I52WzQ+SCUgKUNxzoJbmtuX4K0dgZKIK+Dr2K9GIAqfl4XANxgNPqfEXhf9pQooj8NLpNrxG
ScZKaqsJUB4iNl84ZOjHBL2R714V6jDxU048snf8mR90bYm994IsWtcGdkFekVSYFS1x2OONP7F1
l+KgkturbKAIivOoeI3jODJH+wqjaWV19vMdYqXqS4xEPxejAVea6Vp+si6BSeFwvg0NCMvAQ/qL
9WWiAx3YVmHfmtz2qKq1aSEscVvlEmRv7vlfDCb5ySxQovtR5GysiJePm1iysS/+l8HL7tMj+0DY
DvSDsTGlj0av8NQOhta1e2/xsnC2NpKzwi5Bg0HMPEid5XiNGOCW8c8/SPM/ak8fbAOVouwsY5Tx
Mr3FYJqjabnlGKfjC74CeinigLLxdD0h0K3JTZH4v9UI5q2ksNCNWI4LShqyF5j9aOPBOGh2BkFe
K/b02ck7Ph0jr7+mBq6iJ/4bATGvLQJcL/Z5le1sTfOveh1EnxY1TLzjRaS7Zyw//o2mktFYomqf
kwDQSHDOSByfo1aP510qL9dXUGUe84+Iz94jNM2AV4g/DaBSB5hJR0TVnSIvNAL2T8LUrSfY+sMl
KFDGKxk+q1WNTczjX0OTglqHxfVM1BQs2KPD3rgeL+eul2xZaJOVhIbPVOvTVfNB5EZj04kCaeUq
siEl4NiHDAupvPVtDZua2WGObRap3MKFm398xp0Kh7reuF+LMGW3k05Gcbm2CsD9/kgqGLqj7zCI
uZmp8k+JYrEPahr5I65lqQxAz3MZKjSVfoaHaHKf2ssv/mdsqm9JslX2k3uAb3mQT3j6GTTLmLPK
aCm+OOwcipLRm3A8fDfxSxAuXuVViUOhlkIlXE/ikwuxNlb9VDx/YhKu5MeYQDeNO04jy0N4Wk3d
+lFC8irASu39wg1Hp0tbpu6wZnCjdgA2hbNTQ3aLvRmD/RNKsiuN02nizhIyD671EQjWWRuZnCTC
SZHCD/Mclm9/drNU3Q5XUP/0U6sFSl7AEZVyt6nrVS0lBZxAfp2YW4PKh4A4US8aZLR2QuHcncbD
1YkkwVWeuJt7J6zh+2jvZZOcSXEoZvWRyi+9W+d9rFFID8LlNft8cf0i+m8Mdy3Xvp8CClfZ3sSW
MK19GiuwPFW19IoU/GYs6wEw80sTjT9Qf+2+cLrzWtvgcENSbzO3ZwVsPu4zLiKS4T9P5zSPzO86
zfp0ufVzGax+48/LGJ/GguhCl9CPpD75i/B6MTZWjTnZyz1265btNQDsfoFbRSzOHfiiCi3u02ur
jRDYxZTVHZmPOukELaqcV1xKSMI+9rDCvdVq7GWm95/u23evSAPjqDZQrp708EfXXCJlq4Z3ddA+
5EAYGIn6hLLwACl8wShTAtefVVq1MBGo16zOWraxk8+XF/oGHd8jDQalm2sv/1+K/PgeBuDOJ3mL
xa+IYdoHDaamv+8vY2w8VtGIjr9NKL3/j16c30huaAAoE8Fv0a+MoRYhWKXc3VCGubbbS1VDKdUF
W+gMjFsiGj2GrYXg8S/pjV1Uj8uEUyFOWlz87T96pKnejaedKNTlN+nWsmURHfrCtSjo9OhrXg7z
C50Ugq/QE06Kyiz5WsD5BBCI3bA9jxjsSx/fvCL4vHmMT0PEsynq9ExcZR2R8KK/+ur2PYr1JJOk
IAU/TZ0ewxBGfSHVSE+R1iqRO/cFbMAb5A9i373YYprRjdTvilEdTbM2JDD6MdyhAtm7w4BoxVnr
ukhUwbOoZYRU5bZes1zBmIQNcmiag6hCm93tEW2w5LtXFNNkMEmLrzL+tbGMzkM/8q7XAZAS/HTU
PJZedDp/yVbtIhDrUmlIC8Tl+12oQiA8dI4YygTYrPV7qfUpGMj+uSN+M2wOYwFCsygcqYKQjDD6
WhfbkMwW4s1Dr/O2w6NaWSzUU0uI0RMrqUZNENj1b3tQTZP8ImI2OlOX0PFcT1KWk7Twzx9GWd3b
5eChX8Z83sj12YneCIa9msSsplKFLWWnoLRAg1jqHVzZfmt9FaFS/JGURKHH2GipQ6VV6xWUK7Lv
a7S5lzteQUAxY9LcaKzyDvaDfZu3hmFKLiCKuCrVBUSl7Xk6DLA8DAxgi4Q8H2/t7nsg/VhryrWf
hzOjcocwqUUdwYcesUg0yznU7Tq/phjklKJHzwLdEfn4SZjzhz+Wrb9basuMD1Ds8lMIIqdI1n7+
8S8dgBko5rT+nu6n4LQuBEeCJ+poHIUMrty3U6s8ovJnUlza025RqjosBDyCcaJiXOnlf8rFIZhj
vvN/YwvmJ6QFFGYgfwyUkGhFrj7w61MVEDN2IS/a2LBWQ7/p89AoRTKtdt61FKHoA0C2fLUO1NOQ
mbUqlsOLCcnTKNItTt8XrRvp7MK3+a6wA9J55g8C4+1e2YeeG9jm6gmhM0BqjGYXeyokzX5Mh/fM
WDgHqilI74h0+wkOyC/725x8YeTRCZUi7G+lPreKm2sroPDFyun1IHzQGhBjDS2ojGdc0Jx5cauZ
LZglqA0Wg5k5yUgKrGv/Xs0fHjzsjyTU/V75xMQhjzpcp7PyEB/gNI/ce63krDcKAFRcg65p8ixn
a1+gQKcngDjc2soe3aXtvGLw7HvkxYUte4vqmInI1xriWELmnN67xn0ArAOg/ik7NbOKbVmek0ZQ
sZyLdTwiK1F9A5wQAdXUQjDcSGqR/nVODOYY1/pdBiq9qWcLwwarGTAZtimyRs3AsTLt+V5WG24V
7IV+MuvKryst7RRkbYS/mVRbEveDT9q4YGgXCgikY37RLi59mFiKOX4xIBpM+7Ffb92lwRpaEONX
W/bSGc/+yi7+NjjdZ5vFGFiPst4rdnkXuvz5wGBFRjqoV6Xy71/g4nYkW0y/MYZ6uqrD5pNyju4A
fZ/LzsfnttpQ6CYOTN80LbvZL0CZaO3gmTmzajWLJaqu/d5/UgMALNbvNG4OugA71AgWdzTl2jjP
htOWd1FAqP37k8T1NdkiiDDZvSJ6d/901+yeBeqTTLgddE47e0dV4LBy+ZpSzBiB3vEKQq3xjprr
un8vxPLqZX+vZvvbWTd60v8id1UK+UfDnVAsc7VI0zbjgMgCsCWoLghI4lUyiK63IKUF8HIxeJU/
r5P5aGtyEqwbomRWoXd/L5CXQ3tILkxiWTVgWDgPK8WE6L1O34dHc9pBri3QmILmA7M5hWSbymBs
RB1l4U8VtgddDG1yaCTLcTM97TEtVLeY5DG264iHYqr7wj5gKp5+ZnTcSceiWc8eQpQmNytn5ucl
9Ol9wSy6F5FND3Rfq4t/mTE9NpE1O/1BKL+lNmcFXYHYEYHTNUX9tAUpnATMPExpp9WR+TA5cjdA
ToLWaN3xHm3PvjgNZrGD4ORhvnRJ3XPmAlOhEvy6mv01Pz7MlKNYKnDbglLKSMdMkGFOOw+A+0ov
rY9Qd/HrlmyGMJZmJTdYeBxHHlFFsj2f1M/IgFurRWBNK13GrBbAlz+ZtJx0IRvYY0ooymayFVBZ
emaIIlktYe5dWiNnDrQ4kJIhkq+ZjSSdL0BUZUKTZKwsDCVZhtWuJJLTTp+0guIX/3uhzivMERqT
hfELvkgs+KUkEAzS37wEgq+SZE9Inp7OKw2fn/Tzq4EMp5TqQBVZf8fqf0H8DWR/m3N2WRTLT75n
D/1rYrAgp73Mco8/WyIXk0LmxVMHsXpzHY8YLKjvZXmNyzfrXBsksFSSVES7YXHBOHMP4ho00mjv
1Ctk6TTbU1Wdk7P//76oJKXQCI6BfC8hCRbW3e72C8vF7BRgynPX3bkk7Bxdn+KvU5hwQR/8iuT8
6+ZjLBTkf0C0VzDIJYaB5xkxWSXR+bZmXjUX2UvJoSiJIn64mUTw1uZwI+DhkuGsvWyvnLUGRKip
Vl1hph0g1vKLJYgFPH3uktw4QNyz7ydnJ2vDo7+73nsD4bLGIPV4BJt+yvScCOz4+q+ZqS4c6i9u
Ap6kfU3mp/Ha1cpdLsx57Ex0DO/ioCZ61wLsxEkrvOZLqBESv7+gZRAVqS9cmJiG2g9nkHJpvvLS
l24mxSwaXDePs7OR9OiToLqLSwbQ4HFCYdB+4p1379/pWXJUsIfkNFuX/ueh1256TlLA3B1iMjTK
sJul+IzFIpffQVeluraLSdX4ZpMWQTDG4+D8KkEFujj7BTcRKOGJ7EragJfzepaGaU2QOqjBpJDc
9s0NeCMdo/VUryXT6kc/ZF69r9ilV+jzx2PPGbV41iKeF8ubt1vkumpKf5rtTuaL288EO7DgtGQl
ee7lNCTDFZUmcwVU6B9SjF2J8ITiG8WHFu4XzHFWFThxkOhxBpnTgeJzwGaGRKGiG5x+2iIshY54
m0nSXbEAdLRoY7jqRBxbznTONt3TGVeBSWZdLdWbQEcyvoO3tJuo9zksQGorhk9brTu+mbxLpyju
Yo8HNM0bRTIdNJcfsvjUT1lP071BjJa+fFujwmVEAnRC2oLlfBT61fprOjDEEvuRW9FDgBGSPjoc
s17nFPTs/0JId6yKTs7FORvnyQQRtmgU4ijEIcmXvzoJJnEiVbK49vePf7vnRopfk/VmBOQ+N7YM
+geARgEKfy5U69AOP1UYgUEAzAVUP0T+ufABmhAigdGcbATO0SLzbe+pc8/DypzYFcZr1Th2vNMx
NT9ToUGMl7N6dVaM0oc8EohbJH+h+HZgkl0c365Z8cUJAhnAgSuNFlnjofyQaywyislaolSfcyty
iwrwcGZGIJxZzA3t2bGF9p04WWR2J6QG5rzgFbLdEk57KqxmWIFIhRkZRcM7z8mhZvwJyEDtp1Jl
zf56bYVYMPar4V5P3Vzw0Ns01xXjDOL6vj/PlmKR9JeK+lyoVzEsCu8ozjZ9lMN9y/mEXMJa+wpe
iT32/nZC8NTFoUqbNDmxpc/utvp4Oo4u+ZVDuAmAtrNf2OA8V/IfVxWvi5MXs9LsuiskQFa6vSQc
2ddPoPdzOHruHCqjdIbyOYqmeRdLcZ0LHqikdq1TMiDbevfiR6/Oet/epgCPCxUfiLIS+gMgw+v9
jVBc4ul9jfobxIpQa0ImXU0Vq+Z1H5rCvEkAo4SQcLRRb/M6dd7kX8dDXRwCEoWcXkqWxysKItW9
TlaFctxV6w60GY/ZhDtPmfGz8CQyya9nUg744PDOHpmDqLjQqJJRSFrpgfXwv7bN5EEzF3U8Ml6v
qbZCX9svwdxCDIAYCIfF+GqbiqBBzJ9T1nS0xuFXEetUIUBbvDDrpLms1gTeIf+ewUl6QVNa5I12
7RkFMdNkQupUt6aotIbQPqG8sX4bf24VimaKjPkYHlrp9/w0BSufimTMqDNrvuqMi7r2QSPTEudw
J1pzL8+w/c9VgQysIdjoy8JPR63hEvY1f6SE0QmgVi1C31az7F4WzSu71FUH76C86ghtKk0QMgyD
fW8gbg55EIk7qQuDTc3iBVRWEnm0WK4r7q75bB67UWkTBJI41IOHvNm0uIEG1Fm1luSmoVrih4Eg
fESV9D+/Q/gn0+Xx5cvK7MoIGgGt0nYXQRVCajBebS895GCNbLds8VncgOOxQpOwD8MVZsqWVtD4
j5FC2l/XVZUtdOMHNwppmf/Ej56egUfyvyEjiQ3dajEG9HTaSgLeXErBiEn1zMFSMP3KrZCGAJYh
BNipeOEDReExWj8oMgOBl8dOMx0U2rWmI0yQlRA3QMwElg651NR0rCDbdHCAaJ2DZhdcJ3lCp9W6
8qWqtmJYIDgR78SxSnbnNbUFphMgnDhdHJC42MVEWNwdgXjv5GAPxNe3tRoltIWJeIL2xbT1i17s
k5utXbPO4WB6GRvjE5/Kadnhm+arws539b5E3RNAOqklJNPQjokhdIcG8SdQBM89H89qzau0lVDI
JYYAoqjNsqolcRk5ux7yxqdiJ8b5WpOBpbejGdZxLVk7IFCZAnB52r9XniK145N6PDrCDWWE0o0M
z32kOhBrjpoA2DBEUTnlwx+ojEI8+4j9rsW/bNP6+jH0EnJZJnBpsWffaplV91wk2+f/RBwXluDW
iPyyRKKeqkongtBVNqkBnaygcFslHxr0deatdzWVjSdJ0dw1sP7zKi5ZU6iwSQ2NxGyZTK0asCpw
FnjFM7+d80R83AUyND1ya2wWWPrYQ1s5fXJgHTjRRb+1aoZfU/RVDv/sziC0WElFQJtIvifYOGAK
FGqgAqT40OG6Tw+ZrmACZrgcBkyvxEOH/09kiPg9j3H7e78UGWI7/h0KJvw0MerpvZ/M5A0NWOtJ
EIesjAEHdwAg8b1c/Hr3hNRDmmeVl+sbBPKGnYRrxhDffd++HwA1nh6orIgBwnK+XWwUr14y3VYN
HxZ1IxTrvShfBgnhiDgw2NAUqH++8LxUuQ5nY8hFSpsXKKHYpn5t+qX8Lrrkfn6iqPlUxv6dCmxP
834cyPevBO0XzyrbYRKfzNDMSMa7tUx9wq8/NzcpeH7+cToJbcpVSi1gC0VeYTNWvg+B/QmM5X3D
8VLb0tWHtd92ryP4rTt2h66zJYbJm+lBDBBTrvY/GWaAV4nL1We2EdGto4RLnlpWMS761VQjtkK+
ezt+eFORlOlxCVuBoLGPB4RGC7fM/q3DLC/z5f6RkGQtaranK1Uw3/2ELkNHgkC9fX9DgiEfMvP7
st5zUA+BU0icwy10JkfQTpcATh7Af/7YrA1NFBGAfgVtMe1qo8yBU3x+l2tsn+zNcT2UiWIPL52h
aLLPEX5a2fA6IkpbCA+aR92EIYubXX3oSPuuVDBTR3M5mLL6wam9wm1S9Ksd5dCGCRWZzv5AWcUb
AkgY3wZnEMg7Wnf2rfze2GX1G+CuwhSAybFd5GkvEGe5BD/vd2ijryG1tc1/I4nt/97/pCEoLmzS
sxjM5ORj4Nn1so/npla7EXhX7pXMbbznbF3fi6idaW/38yjd6RvLuRy3d+cMcJ8Gcn4+CM2HhPNR
w4UXenihlQYa6Kf6N+GCAVUyCtK3gY9CTHoFteYhuS7W5Xn+haOm7LrjGSUK7uKcE/ZtazEf+hxM
LMkgxjXumRUhsfeN6d3fs4nQRNENkmolEjcwSGnNJA4vy039Ba3V6Wr1xCIul0UUhIui/SLNKZ2t
ylJgOWt5Dtol9N0Ji7Nu58Oe4Fbeu9BQNHlh0kqAKjlLBb4upJO5GHv9WAt/qTilXdefRJaRHOm/
bIWmM8hVPD0fSW7l2LD95wOPVrdXjqcQFg+WMAFfCaHMyiaorxbhKBFlRek1XRoceZDwy9LQhkqU
7BG5nu475TF63nQ6i1Venm/FDYRl+UWQzLaK+eyKLu+ywGgIPTtouecB5GW8T6aLwREu5AU9x9wM
A9+oOqU/Pol6NOuvt2GMqWkXimYElyfCWryiyJH8R0Uva/9cQcXMZM70XUlaF1shB+AHYtkSp6kn
72hR7Dhq7nDqUByzFdvOU8BsMtIOVV9XNNhZ9gU9shWd5gpDL+1CZWDvE/laOnDcJDJ6hbWzChUj
03b6Gix7W/YkuYMAHh6zCF8acjihVkah9FIDQthiNCsRKDl1n8q01Cl7gKylGgs9DCN4/7Y5/hVN
Vb/D5xUlnnI6ICucDl2IS+KisQ7dk2Wnf/IGiFdsfQF1iAHxQHvq4oKd1iGQvY8O2zgAMuiFrB9I
qBajVz7/rWxXPPn+/C0QKidtgi24up/XUBAAQbOXHS8LyjKL0I/So/c1omDPzXBwgA13ZF1bpzxZ
SrPVR1QjYOPECADo+ekekWsbk6MMfnhbezcERlkHWaHFrnssOZr6Oj+W1lXzfjC4TrGKOv1s81kB
snRV8nKOUuMJdm4wEHmCoDZNxYh+MeSBNHJOSG6LYIccxVLsaopLkkWGnfxPoYE2Rwg4H9Szx1bd
v5Dm5qLiejmXLzsaJc71Ruz4JqZxB2rxvEiglz++eafZA1/ri2rPzHQ6RAn2j+A628P5eeKC/EfX
HhMXc+dPcC6IiPDL9s7KSjp8IR2X9lQ1mdtj69CV+ZlIbjFF2/pOSQAF2v39OizZC5Zf5GCmFid/
Ij5Cw+ey9unyiWLVzlnJi8s7x+WLBJMRRQaZLeXjdzoJtAPKZ1FuPmGsUH4QtP1xSiOmuSant6nl
2fZzpNZNQHOIpLpdN5ZqpsfeLCVMru9uB3GmIoauscEwo5YETPkLHp9Whc+WDkiYPlrAJ/hH/EPp
BAnPhXjRMmfYoZe4GycT3VPWKUjfMDdOw4FmYUd4HW1xCmbmHix0RZ3WPfR9ujoZmm4p6r6hdGsd
hPFjRJBoSzl2QVU2c8annax78RK/cDrSb2VMWrDtFsKNTgdegXeJKBpM/breKoHqcYFFf5LonHws
8UMPXTfQ+39UE4qz3K7cKrnykXe8JWguNXPP2Wrb4FNi0MHs8k6cULK4RPfk6hnOMfvhGviIFwFC
exOIfvLD0a9VBErxtZ0C6tOGjt258bvZPfL0jMKH/n076yXTwwTOhLqVaU6bCrAt6YvcK5ipN2jV
yWgosjnri4SoJaeWQegH0KvYvMxH1agq1eUzE+nHjmNV+VOQOZgBXyaGQJwLhNKwlNb60Xm1gvh4
bVcaAZ4R2TRjKxzr8FT2fUHRT1bu7MCGbjND0nEF0LRcexlqePAjWqWcNKreLnd3hfnLRYTikEAZ
w9QWY8gNOniJGoZL2cqqt6eG+YTk5TeY26nQEAgMgYH4JLLuVWHH8PLbhi9jGYXAqV8dFlCWr2Uk
M9zjgohue6bwNpq0JJq9udLaoBEQd+ju5QeJNvAsKSGLRs2cQsEx02pkpN+pgDSeb5gixmpvwr+P
+FSoy0tDYvVQEoG2+BUAnq7imhFCANeSfFJi9XRNazoRQib1Oa3OTv1czy+LKtPJc0h1YZ0XEfc2
KsS5chp22J7dDC/hRbG0Wb4auEbTz+2osw7Tut29nX96OYA0KqNo+0HnniDQd6rjeiLt6JYr1xtz
yahgM0dCCKDMBvcXM1d8JNMwjCPcIGA8dZZa7Rx680jDWU1fvVJE2RdCraOV7t3dP2GS0NnTfgpO
gLC7ue1cdSed7MV8bDATynFnCrM1LkTe+CGm8Jg5woHfVCfpgpViXbXbymuSYQH9V4FVihE4SpMv
vI/VGf0+C/TdIbzxy/R8TtpSQcfVpiVNVO4S7y8W9/Xfxbs0g3j7tKNx7oopmclkkhPdkioooqF+
tclhWc6SiKWjeZFTlPCRBlV1eg5aYMT7xMB4GhjEGrWhux9uD75Dd3OFL3yxgz1eD1lBDnqpEHx5
A9p6j0BaDsJrVrDCexTyn2jNTZQDxiiV6S5mFSWa/BTpBsa4uAk4uam6IZWgA5TyXadsMeckPJfp
kt2CxTXm4jMJ5HLZe2Z9CNt9QLlpOikgPFnwhXuuTzxYsfOrHYsPVvtZV3CroOinpwG9KHt1XP22
zh0Np+cMhF0cf2owkt2yrQYidIN4WicqSSXSS66n4iqnl/KeO7KymvW2tdik6BkJkxOvLgxHM7Ul
CVn7RKdLfmtN8GuOO1CcsAaoswu1TBW32LEiU8L6P4ZZ77KJiczGgkTb1DkWz7YaYc9VQ2eqdBYF
pxH+df3DAHbAi3k9IoExv2f4j0hDibQAEs0vSVnzTdVjLRTCmV7koKSRAVniKohO3zp04Tw7ujN/
tmc3BiFEFcco1nGnoQqGOBDIi8jJ3D4zKiAmjbozjA6SC5NSOdALYsn6wEE0+1fI104lJ7D6idQ+
3kCNtcLtFu/g9kudrIG2ojjKju13M6Rr0MxvfH+MNNpfNn7O99lWL+7YQ73z9+IZjuNFMFQ/YiFH
CzwpGXidyRsX3WFiVocf990jJS8kxwZaF8jS3kWZdLZwEMDzhTADjk+6pZO6h2EPh+7vjca/4KnV
sY3St3PWlKgF30vXyud2Nap0W2X5fcSbgzt+hLuzRkYxgOZBM5m5RJcmuw3uaeD9QRngEmD9Y1uY
l+ZIezi7FWekY3/a/yjKPjH/hybHJX5BRbjEV3gS7WrO8CMI9TFkvsDcQ2muclCoBD3a84vdVYMc
iXx1lZncMyYwrP2Psbb84MruWMKD83a+xQVLFGAPytfkSlyj4ghuMH7WAOE1Dj66lNRgKdlv+tkp
XKmzNm0TVua8WmQSj+8LrDNN5yfDX2ylk/CgL+x8YSoaitmnHp0FDMflHkUsZz/nHYeJR9myvcpx
E2TtsgsrQyKuNKxhZtGDEf/YCKpTh/Zy0rK3dDkMzbKF51UfxkhJlkQuu1q2WL2owKlsVVDhfe/i
2EwmtZXwrCDKTg7jibiJQLlmbWX3lHmOu+MUUL84wGxMkzXd3AUO/HcEETLKH1DtWxRD0lx3Gr0e
iNLueFtQgmC9NlOA2wSKahy3uShwDAYXueAMRBpz35CGoNY5rBLsJJUVMr+x2SP9fsRqx/5yl1Pj
dOxe9Dp21BENm+ruhcCAFqIigPtz19B6Lt7ngjh4dRut7y2kiP1GIJlx0M66t3sFnD6iTeS7mB3t
NPGD2ulfBfxXbJC7qRerOfvRVPtxfYh5QQTnBu4KmLOJfFhOiioKhcWDNV8AReoSurluVuT7sanR
B53UxVEWbtiMS3CGOz3SqI7fyRF1yUIBLuhveb0wdHTOrKxcw/Lo21fBlyvPErGIIaARRptovp8L
ZVVbAT77gzbn/JTDz86SDmnw+7YMhe47uJN6IJkBLlcMTmOug7gymtpDWmNqB3+40o8lDWT0+nO2
2fFXZj2Ef3MsHMcQTlZ5sDLenupiVrFfVmBOoD6IY5kViXroF0H2zbb6ShMxnbd4RpgYZLggJKmc
cq/+b/9mF627Euq7P68oEpAw7ADRkMLHQih7yxORBiN0UJbnJtbleCgsYyza4PzKbU2SkYo60zqT
JdtjdkLN2qZ+kIHGHO2BCm2bRXBfwDE9iUXNd2+fDaQqNIUeO2ELj97GbgRRn1WuMvMMbY+PBM/f
2x/1hZ80e1XAzdHLF8FN6gLMb3sCHDUbX/qYX0ZKCyYodHejGPpmeP+UnYADmvIQ/1dziTpwpaAb
lcTLt0+S2i+rPlMhAcVuNKGtRGnbLmWRgZyKErkWH7ThEu9bK/g+3XxFpbRsNBMuwcjqm3tlLYa2
xLMSF5quwrcGn9ZPZBhK214tNVNXNBdqgz38YqBcxdV8hByYKAObpb91+APH8bWJwA5sbdozHARY
mPigbcWOLGyFIssLafiEJA9sm4zuUbYcwErRBla+zsentX9DopwVx7ukd8LtHHuP3UDQ19i0Fa7q
ysAFaz8Lryi4WXHIl4w46jqsMlW8BTenseLoJ4OFBDRjJ4VQb5yD2JGQ0ptuBdGKSMFTq4cvRTQL
Bsapglt9lWPbFssb1uAdkwQnfUfBK1CYLBBUqIFMpC6aim6HdjiGdwwXovly/sl4jaxfYc4uOh69
HWiikHbIC/twFY1s2wCNFf1qajmA4hrNPEyYhx2Cy7w97IVik/8/80+fj/ng++anMo0ai6e98R5P
ejIse6Jx3OBxI1FztlWc/0yQ1OYw0dw1FCO9bl4uPxuGUFXgdDtW0sKIUXHR+jytC/0IW4knO+Yh
r89ovWV6Kf9U3X5jnhrGh65K54KCKo8lzu6JsRBjCOJY+12bH0e/23WxuTZwlRaDtKCPwBB1ZcZU
JtJindu6Phj62b+FstgJepeGj6NHJZNWHfwI5WLCU+fyY6VHtLilp3L1og7RK+1dTHBUi+qsEp/h
e9WwtGfR63VsD1c0c7e+EoWKnMvgDHhoy/hFa5V8fKWQWGFK1tcgJ6HtcvMf467ZeLc4+ia6yjn/
rs0crlybIO9cjPk8QcN67cU2/6Jx8hUbKe27bEuPkjxUyKduSGH9Qjwznfk6Qy53GxMiMMy3Kd3Z
TCyda+3j6ybeRpLhm36riPcuayRMvUsOKN/BnCwiAqvRTirI3kgiPhZ79rvXL5v6NOC37moF/U4g
aHCMfjDZXYvl++mB/MvZZWdnVloz3N4A9XQJChuHj0Vs4rdMqOopUEZ6r3gK+oBJi9lXk4bMWsXB
TOLPybKLEhQNvypGaIdsH0lG8ImAouXlL4dDDj4K1JIFUf8YA9Iz5YJ7uD27c5CaJ0EpR8w9zuPe
X2R1h+qjpc00GraPyHVlX2GevpWLZ3tZ7EKWqu8T1uQVDfbmacX/I4NiD2p7Gxc9ehqs3Is4bacQ
DBEbN8qkycdlAqaooQ/o2sRslEteGTmjQ8qkB4P+jNrTpKSFCSiu1y5S4oHuoxCA9S5VYcv9tsIv
DA6soWxWEzVWvFDn56X5h6i2kU584bznswQPAPTDHcJsO4BfBKrdQZjfMzsgx+YsZTtifS3Y4ksW
fjGNhkP5fuDIRUt9mUJTpgrHeb2J3txquQggabJSA/3BoDCVZe592ABAD+jsZKE4XGL3oHKWwWGv
/vjLQaw9vjh9JB4/Da1hT8/X/JYaqNTuot9DDC+eHJBDGZBQrK4NnfS7x2Md5VcdtI49Fj3n+6kH
QIXULGVHDkPKnWz+kPtYTIWrequO/oF5mddvTV6HcUQgxiNZAjCvaGh72jHrkozTzGL7K/UVOgau
EMqFwGPXaBXWyidZz88V31gsgEVMRJGMQivSd8OsSi1kTVDtm1/fj5DBHzrILozhq7P47btis5I0
oUImRWIK3LZ/xqGVXMKUH/dTdeK60lhLyafFsh9/oQKO6xL0x9aNNCrMe7Kh7gVfJzOoUlHR/dbP
pSIXiuwUaUWXJ3aJiWDefMoH1oeIiqk4i4b/eF8G8yXJiNYmSbWx0Wdu+Gn1/1ruH19R5uDUGWwP
SLUgCm7UKHuxYmZMm8wMwXjD92cswN4ZQjY1AujRMLZxut5THvFevkBxx+fpMe438WaG3+vrbO+d
1TiGKtXcp7tCd7c+2YAnav2Oj+bavZYZnWV3/ktfY1yzDEIma43u11V0SpzvM3asIdDtPfS1FEIF
DXsxFuCjQbBZ2yufIQGwX5gTFthxs9LM5uzAYV+GHm+1WR2Os9QZ9nYMJD/NQWk6pEnTtVORI6CO
jpgHVhh5TdfA1i5jLUKIXw3I/dHzyrehUIFqX2kJnZqJelvYFSaibgwvh2ZEXkiM4XpVK1VDy4Xk
muxjLy7zk3kLWbJ5aertEgPfC69rmlPiUw7uIKjmnt5iPQAy043jYFYhShAOsR6Squ4R7Iw/tIoH
yPRQlUK9kjuwnvi8QRqYbuXfWiLYfoav7pV0+z7yHzEcYGsRKb2BNc/1g/39WSjNZqtWoEVwVOUV
Hp2pxXXjpRA/cme5gqaVH/7jEbRRlWNfetA5recjC6HZk0lTL5TIPkF8UR5F3XKSY9rbC11cE19q
xUvlqB0wufQT/sn+Um+Hc7sDRULyAvWcaR/3ICJLGde75eH0xY4xBLM0sX2D08yJdTpSsXWnbmvs
szGJgsim67rjRx4h7WeDdvWlPYQaw2RCknrSehzC6MLH0ItzcnMr5Y6HxAb0Kl090PYdW5AXwjMV
KFRLUUWCQcDOwJ9qIWOI0QSaqMbPsfrZVVO3eFY7jPkGDBC7Xw4WgWvlEHJKiG710o2xmkKySZLB
rMiF8KxVSjzMx1/F4RZyYcKw/SeWooFj5kMJCuedRTiV6AMH2PEDiFV8N73XvUDa9zfu91JdOu+c
P7LqGLWlamj1tSr0xSf6LVgYfyfB+t03wKxiYupgGxIVWuTEcU3ouUmczktGl9qzA0BRofMJFbMv
wIIGNlafZB3LheV27FWMiGwC9K10Ar9L445rYLXlF/KcvnW0Wy6G2orIxETt98ABkgU7vcDWM6bE
d0ihMBu+aw8/xgwPTH3S9hhpRLXCaBXQC464+g/NyQzKHxHwJWNPpTPtBHytfBnzrEFv9VIqC0uJ
F4l/mnaPZKa9us8JAmM0WaTsICvu2q5btgREY9/pPM3xNLVJUyFX54taTd1dXLtmWD09JcbfM0qQ
G/Y9g2HNtIeBu9bG4utqU309Mu7n5itYhzKADN8ccfKPym+SJjnTzUN6Qoal4M1kGW1FFmWs1sVs
F8tVNVuWl2DTx6sOp11Bc/cZes4+2qL94UIwtthW3r3LQyd3ZljyZyoaWcxvsM5CaJ9pRM3cNPc+
9a8BpbyFnsqxXWaPdp0AO3aOS/tAc44q4R5JShAs48ukudzSLQKG8AnErl52gTgw+g9m2HlFzWLf
jwf0X3rAE/9K18vb+G97PFcFmxgyOFbjoNPs/kUTV2Dux3C04SQCTV6XJjsL3vcGBUF0WtwNjDo+
RaI3JN8jswVtEtos+fTvG+vNBfGbUS5cpT90HyJp7+gRQVejx71iw93oW7m4JxezPOGHZQF9qgKv
E8iHfREZavw8EiXtzDuLf/sMhkho9B78PD0cPPVvJk1QSeWRvHwCbKoVet0hTwA/lbxx1DaQTJSh
+Bw3mo9H3W1+vFdiX0EmRJkZdmBP3Up+Nx/sAtAmhcGQLi8TL36EDVu0PlGAMWYNp+sLW3rBt6UC
EngbKTADGrl4oK/+vn4x4r/R4jkI45tSsGe3hGlhCNQDoWCTsrPWBx4bTNtJacgN/Src2P1jr98u
McHOrpMKJDlmg1LQ21vgvM3uKeMjo7s7HNprWMyT04Sm9q8/jsAIAR8Y13R0oOOxasZf5MA3EFKt
Q4JgULfiY2QQ4Sc/pmvXv+ZVh8XFz9yRpZUQyPvIdoPQqxXcbvOHfeZnY2vvM9CPGgxC6eUvcSeO
7rf/KazZMI+fSGL5aVkXpuVa+cbddW7FrW9kc+T/lnvH6kQxiVMyCuoLBIzl35toRu6XPLLp/v5Q
tGGPUMit1396BqFq7zYBgJzBZ8ri/hLdcXXmJ1Tr7Nf3zd9ce91Tqc2/a0Seph5EE+pV6GVNVMsR
OepwGghtj6i5HURfd9WaeWnCRZpoIZE7edNRDmmSYvZ/c9zw9SFVufVIvRCr26+jYyBHuID6UMmO
1tpVz4aBcW23BZ53vZUUFzgffAL4YguNZD2fI0khbHBpp9Qqo23wZBk0fmAxprbTNnFtCMh5UkF6
ziZEYBjQCg0bfQ7QQ1Us1iEqSppQCOus/b0xj0PVxkZdXmS4/uxNOKoe1hk5nFgSRyB/kUkljab0
0mlptUKdS5UUZr06PJ9xAFZ0WoO3hmscGEPTKD8cEUCtx7TiFgHOQV64NQqbE5Su/pJWK+dd3XWZ
RGJA9uiyaD7UGB8P1Rr+jiE82J/07XZlKo+iJyAH4ojlcIdgHVyBvB3FcondRrUp4tooWj3mxOoP
FKY6ab1MpH0QomJAKGUtFiNjIBc/SIbq60BksgIlbXvI1GJESpEBMgB/PAH+Ewqxujx5T3Uqa1ld
wexh/eapJQs/QtA8uOaBsrPLM8pC0Knvu2DqQugtTNfwgE6dXpj8LkdVJ9lhvdzGc+ElNR3TkF/+
m0zDmQ8SaUOuvECyZfvCHen7mw2tyjsnwsczSrKX4QrKWEoUc7vJ4JHhdfgrokLxQZkQ0gdzTolO
lNe+k9EZYuB/XYh1iCCzWjR8NRUvLwPha4fC+I/jvnba2Lp6uHNtD/wj8hS6/puvUWDKy0Fx5T/i
CfyqlDapjwk4GzyjpEYdIPzyXUq/dRq0auwDCg04wX88xwwSJtePjjvZVheAGTkxIpJue4v0Us6E
UugnAGg6zHRbvaycpSLBWf8VdQNLNnfrn+qYnXrrac3GJsVJZJSX52r4RNzKPNSesyEYXg+teljw
9N3Tlvc+OxL6wR8uXbXXmgfLyTbwqEfzCY8Ar7gczbKu5rsvEL2rqs07NJtYwOKg4sr/Hvksue3I
Gf2AP0keahWiNoSxRHcFto0aBwWN6DGNfR58hCDopoHdwk+Dp+yXcLhHsWFYWgAl4eEzO1jlFGZI
B1digfUS0ltQteKaZ7d6QhKEetB8O6o3d900wfNRVccxWui9TunhJP6p7s/jKnFpvNdbrnINpGTw
CMvvqp0opH5TlLQ6k43Lz/jtQj/je8lRBDDHy1guIyXG721yGK6f+JtkO/JYGo+TnnGKzqtFJV9o
/1HzuJ1+wP759XOsDZ5/wrsCFU2g9406E1BOyiIEeqmAeIPiZIuMDzzyLkGtEeEoKGZLnXitjPkz
ri/GhVNE2XjxkhfYCaX/K3iqs/Sh+/pIFNemm+BdKix+WXIxuNsIoLV5XARt9Kp6xu178WUCIZ3j
PFm4QtpFymLBz4QDmUPwxOehwG/tsyblCLnteD7VRcZl31OgQnmaXVYg2dOHYTdDRGWQ38rC1cm7
hLWNOjnqdSjg7HKChxy1Y14gJDDRU/A3O+LVV2CQHuZKq8EbqLFEEcZE1c3i/5Vw6ygQYp68mBLV
AxlxbrG3EsxWjZlKUjOAeykA/6b5m716QPj6mRs/coQEmNMkXI0dELLQvHYjTpWidhBX6Frq3q09
tal+9Ob/2Hj3DkHuElD5+rUw/x0EvE06BR8B8KgJWyC7bPvd9mcn6yPW4FKAP1D9Oyd+i7/O3rsm
MFYhX/D4yoCfaxkAxHSM1ONceD97qyIFH4onQkuyFJHPlCEeBz8IOHIi6JtgjLar90TvwjgOSRGk
NT9emepNH5QpaLeS6kh4s7bRRtzZ++bBWIlFE07ZTE16XMWbGyHkgOLj4mjjttFZV3a8aFnSyVcQ
SGmyVpIS3rqsQOJPrjvTO2vBnlYjwQfC2FWDMRH/BcERwffGofNy+2W9yDiQHwPx7RmZuZkd7AGd
JbXUoR/ER4l13VLXkKHtAI/3typE8QcobUNR7X+QbnNuJWxuumo/z41V8fwvUOLFrryznS66Te+b
pYWFK6J//ltKWO3NHr/Ol3PRuSBlA1hWycEjwfwIR3VU88rG+fyopCDuBRLs3GEf9NC+MgAwjgsD
9cle4ajliwHNo2vddVRDte7htXLp+kkWpeMAuIKz5rR59wk3VLr8xFwApUgPt98PijhzPyqLjkwr
U+wEOqOin5WBmt7tK2+Sc9WdGCNultEhwtnMY/xvP5KpaGbbdzlVDiIPDKTjbnOtK8VTLCIR0X7b
YgT/QB9zhkjseBIy8U3h7Hb02tYex9UYOGYzyW1oFGx/Yh6SoU36Mx3RlIx/tHiNpbqMSxetiB7G
FTh7ek8F26k2m2EnFqmVHrBab9Xc7rKolyIyZKuU6UhoFeWv0L29bAmBgmuB/SXLGSBU+K6ZzEzE
669+0kyLkQKrbCqoIQljO5gLX1oLeXseOICGfuAVuuVsPMHXb5bsGQYmrsNluwl7fcFQ1WMZFjmm
kIikySNfAtGXhqHieE/Orv0cEOCtNBlyjDePipivpHoHdMq2698xEy6ru/dZZ+jH7ti8JXR5cR+J
aU7ca6gUSiBR6C/usVSSuGu+IKZAMifvw9Fl6wsCbYgE9rPIgaaM55LHn6fJKP8Ae7CypL7HRkYX
JhE2loSwEq+Q4FkTywXBTAFUGmgC/nspqEWDs9ZhaoAOqqMuSltW7h/jJ/+lfdk49gavlPQsHD9U
FKsGev7lR0aHEFvw/HF3BL04md+6pfVi07P0icEa8NruurujrZfWxySLB88GphsnVEIoSq3Uy8oy
O0lqYT5GfB2owxTebueFvru+rU7sirLkunnoyoGS2sVgd0odlem1lujtzFXP1LklnisKOnTiZdB/
MABgg9GK5bKgscq75YkZAPKeQ5WTFY81nY4hcA2RRd+31HWz1rnBe8mVnCt44CHDFyWieJGBBXHo
BYYVfhKIEswnF5qE1ThRu9rGlu7+xY9/d8w7BUDSI4XNBVQ579KNenTz2CUe/2k8g2IZIZVbu1Yk
8muv6Z6e35KphxyKSA5E4xvcKz4wu9VZCx1SiyPu6VRD4fMt91LMGvOz7I25Tv7aUPEwhIQjhISo
rD1U01Jy76uVK7RBYc9GcFu/8wCArI2WCj/ihUm2umPJK3e5p48XxXUl0inyX69KrYyMzHkmVUPP
xrxTDMQl6+R345PtR8corG48pGbhZARn1chUTd4GbF88tizaPL5K3zBXa/ron0rlpJJnDgYJMTd+
YwheBLRovJcUGPaAUK/oANthUmRgWHIFcGge9hKaENIEXAEU3BVw2iL+48FOvHfd9o0D11wXbkiJ
X5n41LxGpG4DQjcAcERcsY6AKnTMy+MHbBbqYLL5m8KSStbwNTXvpruJAqcktiRUuPmBP1dPm+Cj
cHldEDxvwklA/XaTidy3vF0K6V+o8l4ln7KFrlqKu2KVZBEoXNgQdnMo8Q6j7P4FNjE7SyqqVBOL
Ot4FgmqLSXQ7LiYBEPn15NgEjA371a3mpJB6t787vjP5OOWGb1asaYzGhaYscJKMy9fSJegh9wU3
oBkbPXxGuTxnrPHSnuflN07tKBm8OQE6aGJTiLOUh34rHZ2ym18B+9rZF/Lwohov6vteRTjg1M4U
4LesKs9ouRdSnjpkL8ZafR2oH8/vc7ASeMPi8AZqmBxFLF+ymmtszwpJEi8WhbxcwvKHI49G+nVA
GLC+NcRBJiO28LrBYKGh1OHGIGd/biufYHZe4EhFY7FHkdIp8R8KyB7G6Hp/jZtbb4PWyZsRbKFr
BS5IIRMhFuQIYDHYTjy1eH46YaiDUahjvrPSpOg1irsapqEp9XaxSbEHKiIT/InsBOa9xCxj7SpT
jfHSqUF+R379XR1PMa1G641V3KokbOtNhnqDC3iPsExTf/yNsoyBYtu0qKTRwclrxVfAeR/zvb8A
Awq2a67RhfDw64t1V+KS+3xZlIEALdiezXkSd596CrhJJtzeNj5yD0GHCL6l5zFpbCyvzUwmjgY8
/wjlgwlzAG/4OLx7X2APwkuyP2PoY6emiEv83k/etEVoeoFA6bB+5OUEiaxpDBOTp92D3pdsA3B8
B4V6qqp95BbDEkUJXdKqnYYUPqVLebG0cK8wfoBnD80sWKVyKn9nrTZiFmGs8bz//cTlITd4+iLx
9FSXdJ/dh6tiSQQ6LQKVmkFdmW5vlqkFkS9J7DPXL2LqAoScod9QCyPZM0QKCGx8BfWR6U1SVuUv
6Cps5ovhvQjs/+Bxi55x05oBvP5vI7Nmbb89ZiwNaSoRTQVPdweQP62wM/RPaIaggrFioI9TIVZ8
t7ktI/MAuEMyOmXgWTKRE56oV5l5UWxsJNRmNcTX3R68nLrkINuLYUOoRX7rB2+jYd89IObflwvp
zzwk9FNxts4ypa0lKTDnfW6zPNx8HtXhC24uZkxpRb8Wwm1ENEfshLLhCvPoEW0spT5rvWRp0L8R
RVIRuGYkNcsBEeA17A5w+0TTQEgST28gIapJkwhuJRG6EPA9bs1Rr+vAp1cBOUYwclmbxfwS1KeE
4+97SAK6eGvJFLe0Gfedljco3TU7FFf0zFv/LxZD2HlgKJlvAn8j2j70CSUEWmGHxDn8vsI2oMay
FT8tCg4QaU1NcyjdpSmmc80XPbMTUeUYpHQIJArXoENCLYM6Pe3rtwuW6kt3otMBuH6T/CWgOtTN
+/ocd2zwKm2rtImNlC5Vi3+Ao7yRp344JnrHRnJjgPgKWtIOPoQLf7HzTAmpgD0NhqoE/tcRCuhD
k+QR0YpGIMmO2A7MvmIvwLnaxBMYZy2Cy++PeoiFSjkHSnyFjuwMqQAhsE2CccLDpt2KTxLzP25i
nL7ob3FxHS28uNQHM4ebaZ4HBxSTC19ERjabnTjctk03gwqMRjBNcWLUuZvMaHUctvb2bIbUNLyH
057xov/IMUKPDMjOn4hUiz6KSMK5usFbuM7dvKHEnqfqAcpV8hFmw2Nsc/KcKksyzL6ZpLvTLVuz
I5G24PdF7mjoNA4NKgKXrNyTFZlh0I1ezzUyC1e8rgpRRccomZtjo8cRc36VCnczVAfe0lkbSpEk
pXvOWkuysZz/y4KxjONq9DoLBY4qfGQz8fT1UpN3QTG+ITiv7NtrvqvA6fsxb4Zcf9W7jLKXcRav
jis44Yq97mDfysKD1aPTfiHunm4HvbhQT9OWj5jKFMPxb1r48yUHd37LUkSczDjhxTL8Y0udqAUX
qklYI9j1hXvm+KWmp6kUcQl0wHXdlyMaVDaTfuqEHVxSW7ItS/mlGEqBp+Fuet8r8JwbRfYucwHN
AgBDYhUvidcz1EzLG2fwlP3l4WLDQ6hDefn6Pz6c7Q3/ig1wRmbPwBOgttD3kdYiWpgUV3GtW6N5
v/sJ46IoK3D4uF5xekoyAGtjXRyhsoBc/ya6ze+0WzTigN4QHK3nTOnHLd/v0iuJwtp1STYAcwxa
CfIFksTsh6u3RzKhC3iqaq4/nhqhA00NmJ9DgrJKvWFYCHwx94/PljJWBAOEJu2be6cL2IfWDoAq
/s68HJwa1PEDBpePtjJuH9qTM1hA+TWsHcmgRZTH/SCDwpu5Ct4zuQo9OucAZFax9yVTDUt7wSQF
HyLcRPDyvV6CHhIYMLnGMqUqkjq9JBNILm2O4f/PyYm0n/tNwX4YkPK8gszJtmGTQQkDcgQFR1an
qmR5hUcpQwAxMpwAJ13zHTl22p/o1gu/neG04/16/Jmzh0gQHI+SrHSM4DzYA1mnSPdS/28VZ4pT
aJFrLHZEgIClhaqB173roVcWrFu2DEoyo2B46K+0nSZJ1q3k7grY2DhsB50ElN+61Ot3gmhhvBuQ
XMm9HOV6upSCL7ZGW4YLzvJnuLnq4JEJj9HcduQI0MZeXXlg7QQNFDVdDMvCyAh8N2WimiIJXyML
BkCNbojGFVG2IqYV1GKrAJe4PnfIO535SIKk8R4nc0C+Otrv//7DZNhWI84SajO6WLtvfZhPI9x0
CIsMq50A/HviUwmUmGV5dMPXUkGV3fP19/9uSLpyUZlAHLBT/Gh8i385W3E9mjVg48ZOkxMJzgRZ
PHc0F8Uy9BcZRfye/9PCDz4vklvG07yz/Vg7yOdKjc2pJ+XY7LjSmdMPR4Jj1RVZhuuzz2/HmpdA
/Vppl2V24Pr++GT+epmz1OApDrx03PksdHlWaNYWete6GU1G0VXHn1e/cgl0tq4EW3UySO8Md6/G
wcMfbntBQh3gnmQHbe6jOOibqg4d5AKv5mvNNPqzGvP+VvP1RzLV2XzIDVnsEBdo2U0k449pLenf
ISYVUYt99XwgTV0fBhCSO+iiE6Z54pNM1hD0y1UU7qhKK5Jvu2L5YgovPtbdEVyVRqtLxBSv0dXO
YncbaLZlFicL52DM3e3qIDvEdBXdaVJIBx5Jo+z/7lY0p4qgMPVpmsrk0acbCQURFwx3OMDBTt0d
sCABmenaTVXjWP82xzbWtDF2Q3TwoE6jsCF6TbSTMz3/nTw7dztVljc0KQuTkDOBz1X/cSVmz+U1
siOQxM8Y2BM5Lh8JglzYapt1E5KeIvOEnLIApHtC3vaPn3Oonm2vcSY2g2A+WwOIb8Z6GWnqqqNa
7gECVBqGhVPTE6WxyFfji77Auo29Kn3cwAcus6kaCoJhYuzpI53SjwkqU9OxFGHDgsKwdlDJOXRT
indwlVD1oz0naxcmpJCCrC/lC5sLQXLq/Im8JE9x/Vs16m8ZHsD2BRz4liPNqCMlFUYxgCiudBAN
0AOeUEWyYOp8Kje1gcZJ5MnhMDH5YHn0V1bND30SW0FONYezxgvHDZ7itj1V1rgkeGwU8f4bvscD
TV8FXwm2q8vQBXPyBgKulONMvTGO84eEeewFpwbvGO1UY2lcuwGxy1hZqRd9779SYC/PJdemvG1M
3Ep49qrg4ntN+q5s3nRc/gzXATUMRulKaADVt/eGMhzh4C6rtBSoJst4HQgx/+igmROZBuN/aM1V
0zwL0TzV6KbHJUs1B7eMPUyk+EjX7vLx40jxow//WNCa29DQt3XNPt0DvbiaI/8MtUzwJw3KfoIX
qjiZwCPFbxVvIeBo6PP+A6ut0MXv0yFPcnYPasYK2H24lAG3FKpRE3D+K8Wjk8EkBzxsSOLxbNZl
Fwwxt9FIsSWTTqnPg2NMyL/Yn15xeN+gOvoiR/EZNR/4A4jksbplVu5zZ5gzEoQZHscTJjCz8oqP
2hCJgUDzM0+21urmiCCaXUzG4aAbFY8h47yvxyUEKKc0Z/mgfe+plQgOr2+uq8cW5G8X1/dDaBFh
GM581vbKc4hBjZJY3uT7T1tQ90n1S24SFjbpwYfCmlQUYEDXYs/wlp54oFPfUjBAPhMlbaUdx/Ax
V86aixHzh9TtOwyodCSjl8CNE7E+FmAmyM2kEuKfQKULB2mfhaIdjPo6qMdHYA6OS/CvW/8dOmAa
M6Fa3Iwl9Nazsekm/NL0Lj+FevTPsy5EfWM5cfVVszMXtrm6edOTvoxZ+dA/JDVbwZon9dkCt7PP
NawFHFlml7OeFaLp2aLFMYb6RoCX+Q2yZfnYkF/mMLCs15GQ2LBEym7eBRtUbalTgBTJwyJbWBA1
OzGGO5Gc9juluvEKVFpibmwXCFgxn+e2uKLSt6RAYK3t6D4D+QtIYmU7pZijs7PfOWcXfiJC1fL3
GjZHyMhSU0jUN0l5IMaflldo6ODukm0r2VAvYqOHLGMZayPa/OTq778fY5Zr3ZbdHzkryB3v2moP
DGEDN6sjsc2ZWkpCg8CW9OW/pvVKPEkvyC++BYWuccarrnBiXOrRkOB7XGJhVDDdK8O0ZIrUCxbn
ptYzE6StwcVf2BuESu0KvSKvvw+NBkCbg1wAxKm+OQswoPEPqNh7c94zGFAQmocF4xYeXreRlVoz
hpAixfJOc7F6H3RXQI84IcUBjSbD0QM8zAYo2sBxik/X4KAzf0Pv8dbaLIsTFGX+8ljWR1Q09eJS
vb/+v3OVMQfwX9eN0bsrHoR6x+q4yKU6c/FCxGl7oKKd7SZ1k2muxNE0zOwxDNyEoR5stG5RWVcn
FRxM4JeQGGdpC8+PPt+swX73MkfHnatAr45CkQ2keEgfYuwLKnBgM9BGtE+Bi4Rt5UfC1EcoyumO
dfv+Xe5J5oecOs4b+oN03g48GcyzYzo18gGkFLEZIzbRKlapGHvfAt7kLwSed6t+VAuFy2ga4qiR
gd9S57csRchqMw7bbIDiWVY/ttPFXRQaB/YuqcN3w8XqxOlYcLaHfFCYnWnyR3MkPSift7ptIY/G
Iy4VwhXnHt9u8F8ri013d+1eqmS3BTDJwjuQzWtdwz7EswTgttfJWP8oCgc76f26Pl1PPFSamRIY
VGpwxdZC/mWoiG44ISZJLizKcF3D5UuK4e5ekryM25XiTmX9XebFAiSu78f/EB/RyE8IW1AGK6WJ
fdT3zSFFBoX32QlUavLmZUcq4br4zJ0Tom+bvplgxFrB7qrb+eYwAnnSR9HZkB06cdYGuxw5QZw2
vFwcljMxVLq5/PHrjkpYtSmVqmHCNvxj3pY0kCAKFWg3NMyfmZ7p3tbJ7q6oSbyD4VoA1wJAYm/G
+4T6e89OKiCcKp/U1lRcIaC4ohJtFPSNZmuhUmTRIDCDOYak96+M0JQP5aFXRkMLpvacmPOdgIqy
hFnUdNU7ckwj7IhIN9lSoFlU2avTMSLMfVyh5bHyRLlG1Xq9eBWLNvniemKHv+siVx9YDbDoHF84
Gi2ndDOixTVBokhjBuiYywDvpO6oOsA/sKlAlshfXEfa1/NqWHhqiUtlnR6vvXtnKRFir6/95QTg
I0bgrgqifaIYgSlPEIlXZv1XwTcqb3kXy3JQMUxZzEINnEWa12PyPchYmfrqbXKrZySC3XqKOisY
Z8kWY0vIgxTzyiEM9p13Lytl7ZcN2hlwYuAs4zKQt75XNHT4oBCnNtFyu/UnNhhBK2Va4kOiSBTj
LwJNx12irryb/FEwI8L3MrqlP+4H3dH+0CkSp7GKCv4M+Ja9ileyhLBsaUh+y9WZgD0WOInsxlZC
I/sWIafddKXhk/AVbIMzCCxIbB/aQviXy9HLl6MhRMVo7jVvK8WQY07jKaYQnyWO72cr97quAAL+
jNVB+31ZiKQNk8V4ZCpTJHpFy3E9spsgC6P1Lwr7zYlkOicbPsIKpInc1OhzSC6OtnEhbwduemoN
eBgk7nsEjG1DcUA7EFz05ei+BqM+oRPONQRK85oyTq1DTBwHC4AuYVktySQjKWbcKy7psQZ7tkxU
+cy5VOUaaYUbN+H+Hl66saWI/p89Uz1iFvG5F9eTxrxFQw2bEvRGBwZfwaKw2FvrVQLDPMeSpHE4
3XLo1zxayIxcSWylKkblXYj8dqBLlUKyHRc3YsXmj4i9NMSlP8uM8CSPAxH9exrpeqA6hQpMkKg4
ETLxhiaUiZuWvN7hG0qTBUcBPJVCmaqZnSF2EC3igDQCBjKIcqk6Ye+uKP6LLkkB+GImBwgLWd8Y
0eqR3f0kHhuUjK6B/KKdhXfCJUrL7ApFuVHzZa0zMw1YmmwqOVtX6LTYwHND7X9HRCl+cQMBakTX
Vs+tcGsRswnlDHAtD2MK8hRXqUnORF8Nt14pXdHcRgUq9/y+vhzsQJlE6D/idHV1PPycEeyzigL2
570/+P2gA0CBpZ22uh5o5ZLjVp/pdp3xXInX9d4zpuuAhEbIxPVZcrOk5qyMH2JXg5RJzOvCS5nw
538TfPObSxkg9AynsEMNmcYVpGenmnsjIISRNE0J/yet0Pt8fwoDBTyb/lJtMxg7hcR7t4zqJsB7
SAWrJ4tkZQ4kB1cgTL0OxGsL/JPtIBu18hubyJp7jccpCrCiupiaZd3MbaNYp/LfSHCbmUDd4OVD
p4CdZcIuAuo5a9DTRHROa3iyrV6OXdn18r4LLVy3frcMjVe3I0Df/8uljRwzTACNpHzNk8RMseSm
aiRYM8+tlIichQME1HMF2iNqrOz5OhKEwKvg6BEhz0bV0PC9Dy18igRU9k4jb1C49ZAV51IM53Pp
vnNFNE4hzVvqftatbr6goTHGJUEDm6lzZXf/N5JVgNn+pOuxQgy1N0rxLhFbD9HSypLSEB+VEFYT
K6dr9eLTT3ZoJ9CaZ7httHYzMf5gX3kiTJ+qC7GghSnDjZRgf0zIqL4iAdIYr0nTFsm2Vtc5QQYm
C126EQLnko0FD36d7XEgJsAl59g33lgSm8gaVCmu/lG0RFeeawy2VKxlU2ZKOWsjsLXcBGbEwCmL
yFXOgTFPulRg7859BsPKRpEE42x2QMg1uic+e7qyoHr85MZYi7co5S+1sggqsH+nmCdelXVXDNBF
m1uqb0nXjWHHcVXzQCTWFYwtoEMwNOXWUn3uT3jTM/Pzqqv4T/+1oScoqq/IY/FhALk7eaOZT1UP
cqykk2o7snHm41LTCXGWzKtTHWSr6wt/Y+5AnE6H+nZftPbqRN3ss7/Ip49dtsn1aZji+iNCRKPP
i92bSlgpUnMwE3lqgHAU61meF0Oh6Mt7HFOC5B04nNzwBvP8v+3O6oPWeLAop8/V8Rrdjof67+Uq
wkf/zPvDgnlD90LEqpBEOI8XnlFTXz7tPzAUxt6PVkUy02BMYLbKyeAa1jJB4dZrfXbKqRLvaVcn
Bo+/l/HVjKAhzn5zqvSpHUlp9IUW82JHAVpEdqMPrVpv3MmCxyaITxUThyaXRa/I/2QLV2Tg4CRf
RdW3xVqa9vtQjPuTKyxo5ToF4sG/+SKAbrBbZamqoJw7xXiBCfBoAeDcQuttPpCuqFGJGS7Vu3pK
y/eQsy5rLQ0GgAXlntjYFr34oj+vRhHr2uizHHRSaUuG9T2sZ2CN6vd7LT4eKn8BVyMkSf5eGzJw
ATl+z8vIITHEMuLdi7OPkP6LMC4hAxcdcgSdkQOXdFtiLlJPak6d2PDmsPNXE09IN3f7/3tuwtJV
rHph3sJmnYSY9rT08lNy+0FkHuuGDTKrNLy1tI1ktMpKdpoIwcE/DRG3W6lFbrDnIpZQI66hQxT9
lyTgabbm0xL2LN8XnEEofaicFMklbThCsaHcmsS4mJcrtVKAHAOyUAlD+6+fpdkkEmY0CRAO2jOa
ilQ+oMC8fWrjtPikJl3jrzrwvAcD76J5QsoxnLGlclXFPSmpv3PupVrNJQ/CETySMtP8jGa3FKyR
ZBF0v3SkDA38foxwGjIF4M8Ng5BXvcZJRZ/JXL2F0cH3tURmeJaWEzV7vARmOWU8G/clcZe8woWy
B1Ys/b8wX6SRUZBLoVJg6fdgaGg541LZnCzfsjst0YBgrCzFvJ6jHxYg/ER2v9fMKdBRllNzzl8h
lBwuufsdJquhzG1bGKvl2gMOSuM4Lx+b8ILAI0NQ5yutsQU8rt8I+FxuCb/thrJYk64qf8j5rT/9
4nMBStVACWSWGTaqJdrRSFl86S6Zogis7MWL7dtIzvxPuDNcL4ofgCX8L0Ut+K9QU6veR3eJBEbC
6O3qu3sceT5zXvM4CEl4YmXACfWXkkVnJcDfNBl4nlvGSxcdQ7i4xqaDovx5X2AyraZUqTWGIu9Y
oKTsG7dqGafEhNiRVyLDVFG094+iBQHg2Y9oaT55ifGy8qe0pxbZdAvAfqMRwVea6KrR0t3lp61C
xGC4cooXMP0KMclGW84OWcPKAo8LwDCRzvcQiThSFBobArY391WTDXBm0rlBy/o8qcvEBI5E1ply
rc657SBlO47DrXi2O97mcXycZz8dvQSFb9WKht7hXcnNlp1AhpP249HL53VOSl37LOXmYj6t0Rxk
jEaeqmX5tWBuOV8fEk6+YciVGPSNj8NBnav1v6/dqj1xUDjkPKcareuTrsdSy1vtneadteytRfgd
np+houvPIZXgofun9nodPc+hPyoRBSnCEIyIE56P7lInwcUS+LXvzpDPvoE09hEJVybnA9vL4lxR
g6VR5gO0eGwsTNtAK2buQ+fX9dlQdEDbk8MB+OXd+QvQNy34mbeXUyiDcgJI8Muw8hLcdi9GB2VN
OE+uyBiUiAjkMTlPbaGFD9QIIAagauhjmTKhAhLsaLt/Ef+tj9a3JEQmIdcw0i6hA5XxHyvBysaZ
MY+q06sl8Hu9ZJXNm/0KDb7hPq2rdy7aBrjFDXOcMnTq/Bcovgtq8B4IimNBfp0+OMIOeI5plei4
IfWUWrqoUjZ16kX0hGqMLI7ZjRDkzEh27T89NMM9w6TvQZ6jXuTd8rsGX9fftA0XGzXiXqtPZoyR
vwHZyXt4kQ5JHxLMkG7aJeXsoeqvMS0j3zSpCssGfLsHpxSgpCXPIGBq+bRe5hLef0GxpFepqMCD
fIn9xg1MZ1lonRRS1EhYA+o7ogfQj7H2srEkuZ3E0pvqLIibteUPapZSyvCQ2Vu/h41SPAF/Ztyt
tbghWjyB79AlUIrhJWj7YxUtlGxNKXxvMJwC7DhVz07DbzsXwhY6G1rk2EAC/d2xumoQn8jTvlz9
zj98gCh9LurmiNBMx+affW5w7YmSAASLFtpxj1pYytUpWvN2Dt+2hBjSbrYj5SDI4pjE801DGv2y
kFsxUh2DBDaT2r9YARqU+YPfUa4szoPJHLWeHmaLlCXrax7OqtZTXQj/XF96rqE3aAa6nuwr/Fm5
eny+k4DpNUl1jUnJCuy8Vh0BA1DhihZXcX0JKdUtdMKNw6+WpOx/jnHV7HjDU/kNn1OGQcSPwJd3
kJbI+u7CcTOlceO1Q1OIeXvBN/R8O9DyBajKCmW7xYJ5DbK6R7MF0iYQie6+udGXX+BLiccRytxl
f+61/o/Qg9ScfHqQv8o+6Xz+LFPQzge73PirNkBdEhe82d9bts7Ujc9Lg0IlIBQ3oHBjx/SzY87K
yfr5SX0VWvoMmslDlgJRxhKeGR2Y6MH26Via5TDE3SjmysNga5/K7jHj0NzL5QHOi1xKUD8M1oOp
LiDCyFHEtohxMMMPeuraNR3soC9vyDFbvH0h+8fFRwET7T6+kXA1qvZfdpcUMOMS5gAu5y2tcm62
MzSJxoWfWqR7B8o2Lwq/aUgf+A38WRf3R8w1FQZC3UIAXW7og7jk6cxOKx9IEgvQKB68LiH7gYg3
+NPcVlpPaxgQsFwR2KCMYB4G861IdUIkSflzi6etwLnrzP0vJYvrWaGPwgAl5dMRJ+IN/rOtiGU5
202tL98M32j49lGo2Go2kY/1tewadH3yL9te8X1dEFDNuXUwgk6HTYicaan/+KjZxJ8fIw94oTT2
awigk94yrHviXqd1RsGODEisTM2D0PijmhzVSpAckg7LsgbMcTfBYDGI7ewBMf27/oexRHP9KGxL
LAzpmCg3wzwmK76sr4tW1o4YbYBwcok0WBLsCTYasSVSwteK1FVEwUdMzGzbRsOPwI5sdA/mr9FY
woA9oJhE2qwM7xxNDpnTozULf83Lwr86TclaqkZSG/7z7e70zCpCqEUVDBcAc6CJH6jlQ/+MLZ1h
Cao5HEqbdcQFgLe7ZHoucP2GV4qetv6H8aCqYQ2v71uSW9K3WAF6DIWnR2Yu/S9nkbePP0JrwNnz
k4Cun/u9GsfmQFrhFkZrmhbfIqufKh4CowI7K0s0+7GPPgO/BxSnKzFl9Rd7eOMIPP5aG4kKR6/6
DFW40MJkplV0cktCTHm0mrdq0MvzAsUsF7TdgZj5rEim04TOa6p8gG4Q8K8LQWlmarUbaycU2WBJ
WcOLKfXCbkTFRBtAMXLknEYW0FVJSzWKvOqszFUUQQob6R/uFX6AWIVmdh1Gmz9dJn185YY6Tly/
6DY4qiQnGQhBU5m0sJOsxJBD2d1Zv8NztvodeNkqbibU0ryyq9b5neEths6L4MATqSt7SnaiePo7
2dHuLj/9gwX0qLHyAJCENUPgJMJH5hPvyFv9NHdrSQ3KA88aGu9NMPeYamK0J//uuOdY13aRbfEa
1nzZu98pzF5rjVqfhDoDE5FGnDaM9hUMYy22R+/TWzCihBqeR/TgZUVJhFrAXgd4OOQTAOBvJzki
xhniQV7oUuHowNezBQP1drLf+b+MbE7PeHUxFU6zO1inRLdkTJKC/mqRG1wJn4krN9T/Un52qUI0
bnH1Ik9sN+zuWRy9TcT/vamR8t/Jeya8AQg0fIl90rSdTrIV6yMGbtirlLA7jPg9eBtLuGLrf7vu
s6UDSgUF1nKW1xYTIbDWRnoJ/xliPw458a2JCVLnP1yXmGkrblAPDAEYwGgY+lGwi3ufOAI3d8Jw
omV2n8xHYoz2eUxXM7VCSyV0Zh3W1EBst6laYmTZK4h2LFfrusy2Y/GH3WJbyhpeuCt7fFr4gJzy
+YgRSsC5kaHHFp+aLwpe1cXSzl1Hg7Niw9v3X8j0xin2pzZpQnfylbq9ynvXMWysH4MBENpscdd8
SiDaVRS5XX2I8GbuKxomCcVh9fuXJZTYSMt2I4DkUNZEthndh8U0dari8SOdZEuMnuom5jjX2eKg
mIBro3YPnXKrjKkjn4ehJVvu+uVhNJuSAl5hoVXMNzraRQ2i0jIpyi5SKDG+jZxJSZ5msArXU0/z
4TaeTXkNY/Kt+e04KT2G/qCNRZgCF5L5UTDnrBdZg0UN8OLOP75++dIYJbDSVG5CO7tFx5CGjzpE
ZNzXZZ/Gdc+RnPsDC/dQcQZrtGpDRBaoeAYHjc/EuwoBWBnvuCk7Gexe5q69fnkDYRvYk+KGdurm
KrkBcz540RHG+ox/jNpUP3BwrSZ2baKzjDVU8G5UbUN3u5Ac8EHgnrSVgtnRS5ovtbVBJMIgmkzc
70YYVMPGVWRxrEKusBHWpyNsqia8bsZbpHVD8ISsr4JT3uKk1ODASetGsbH1osiymHHO1NE9MqfW
a9zMjtNAFnr0YqYgSsM9dmiftuPkkfSasSrOIHXnOWhcA/qHj3G/CIb0Jsb0h33Pjk+BrrfgXZ8P
a4/Z5SCyXHvoiMIClUFW88w4060y95HdL+rqbHKTRUF3ERKKCKnOzq7jg0N2gSSiet3OwBspVmlS
IFhrTjUtamjbN8VWampyQABtzamFzU0u7kPgn6GJrm+7ghgyOgp1xlcZurdmf+hTjuiVOEbOMnwc
lwxyKxeF6l7LAg+3nOPxbyqsxFVT9HCm89VdeqNd7J3buXcngJALSJNjSBbn8yt2qlmZnWvU7ZU7
8Q8aZmJRg5LMJ3mRNgAMLiu4x8XhHs7pkIhgsmSoNaHLpvuIrLNTFoelrnnYzOLipBUvFj+VMlcv
UaQdIgtN30quPzi4sWN6vYPpvMBzp4cyz+rAqPRUI67I91GsT5YDnrHz34eLslJ6bcj+1FS9J9er
tqtW4kwz6QrqqtbXeftUAAuEKnT3cw+5/EkNICcuVkHo/MgCTovg7UYwpDrwrVGTxJfeizGcaU22
Pt8CagO+HOY1kMN+cgW5xFtts6x4tvV8WTgdnApRzMOmfTUJLJBLX0sHW7n7AxNrXP8j4wMyP6Rc
orBKHraH+8sbBiSD+YgCm+5L6bgd4N2fYNAILF38ZPtvYF2a/NRSfsh20Ji61X6y5pzl6c95H+zB
RVwFBq2ZFvty+VOuZ9X0rbqw5LhZQAJhHL7xsItusWmxuMPITiUV9fhfvOTNwHLi3U1J9K60KvJS
Sgk6Dll34l8gb8YvJODrY791BLZcfYuaxGyDfes4IL02wcKgMJRT09KbFU1W/f10SM4y5aQPDaBr
Bga6oFgYugT7jZyGfRvyaqBVkvXIZayJAdgaH7Jhi8MPDBE5/VJoO9A/MVa7IdQ9ySFn3pBjEnXP
ti5s03am7wId5fgaa1vzHC7nhAV59V4ligZPMpu/n3Jt4gG2IBBFTNfJrFGPmMEHf6jMXtBRbENF
kRocVe+xGNHwtAtJiRo8HwvfEObgu1UKVR+4Nm+0HNBfTV6B8UIdi5HGFF02bgy6VM9jQUvM0ZjE
Q26OwJbmnHX/JSAnxWO79lbjB9Vd78Epl0jO0wkhsQb8H7oIAGhVLWDBHBBd9+neUidOdvy1y2p7
XS/ZX7ZsDtviAUr+xWOZgaPSNNsw817bZ1LRH7VY5OILRiwqInVzf9KLC5NEP7euFl5UgYU6UlXb
fvFOFUsEXLiVEXgZVYLksjN0d1No3L3nXAPYJwkbEbvTBk+zSKlF3KXJe/vLFzqMT0GqoBf4fy2N
4ljSbWgZe7crQOOk9S57J9cPk0QHM1EBOvcC0+NDYUtnm4MX5v9G96N16DHV7cgxx02AsYp2I18W
AcXfvtSvd1dUM+6BP/FfzrSzxWSz1YVZm4dprvwO1qcb478wWUJfzBn6CNqA6KghQOwgf9cvtoFZ
TcRp2jUdpUKVMJnrwPcoKrfYIHTH+LUNzMMxr++HvIVAVTOvz+hRhFuOIkH1wTLo626K+0H8pmO/
W3XZsKh6lPFCXvg+p0llDDW+rdK9AEqBdxEkcqZeip/xkaKAXxAvwL5vVRpecEAy0+xIvvUPksKU
OTlaizz89wnDUTQbpys3yCeZfGZL1OwMbqIdCGicGsZf2f7HAboOgTOBPWv7uz4mXzDSprekw0ka
6VFeQE+klNhwB+RAQPEed1hueWwZCyLeOvFoXZEpLlftNCbcUeoQmXupBOdsA/0wPaJcCSpj59c8
IUScPUSeeufY87cGwxJlmvbGaE0U0jOsnnWrna6T7D3tmCtwD8p/ssrKmZRrNa5IViaXZibXIB2t
5Aq6WvQhx/KcCTuMwHj9Z19cSMWhIbxClFmKiNd5GCs6NFsNfbZxezAxDQzg3+iZ9pQ/xZaA2XNe
YeDrRJ1OwE1c0H5Kx9bdi016aJ2ogXOm7DGIBGnIPm/hbaQpK3htaNL4OIl4ftmqEl+DtXiYR+En
m3lUNkUmpF90nC/cVefI0nMrgMG5Q9DYk6jNLiC0w6DnvoD8qjxEYH65RCo/F8XDFdXvpmSzOs7i
8ei3wt+PsW8/xPzzaLd5kHvwszYvOJK3dJYu2Uav+YhM4biL64JXw3GyJm9kkX0FFwYkfIVfK+Qs
BjmF2W4jXtXKpcyclqlGl6an1ErD6v5kBzyIxz1u+95YgFZEt8Y8HeOX+yYb4bLRv0VfpCdyIwyv
qOhoeUiPnZz4EPUCrEbfPiz2rTVXFHwwufCGBVMFkHgaplHLZuEYWtIr4OUlqWqGtZcN7Aowu07E
KHpFUatlO9gZx3UZw+sJoeGivYTrHEDqROfLdVR4c8k8LNikNlpaPkvdTYwf8v0mBzdDW7i7fnqX
on3tX9rofFjdcqdL88EpBXShv9bfozXRNm56RwNA8SikPfllk6uAyyM1u1ksTzwLnAnX9k/T752A
/g0XI2+Q27rZuKi4NxsxFRZ20vbJZSRSHh+AIufJ9sw0OmfpSsmRkccOQAl/8TQv+If+lkkZXYSd
xQ1iBq0LyTkgUMqSNALI8paZkO4YxZRWQQw8dQI+O5soQ2gm0bIgAIqaFDd5fC5nXGuRged8wdcn
4fy2GqFYPDuzrJsApoVCb7OxSyyLvH/01wL8Va3jASoy/dRoxNe+lvmmBpfltlZaGUAOa9gOIUYk
WAb+IzvdcQHgPExkxUQfVOl8/cMW/DiGvSAMlKjffoAx8rJ7CjpyFTrjNULvHFQxlVXEFbIcQhdg
p1uHK/AbBxIJneca6u5c1l6jBM1uKeV2yznPoOcu11kn0T7ha924FLNs7OZaQsBTbYRl5nMOhemI
m8hgMuCLHRH9IM04UEGfXx7gKFsjxL8MhXU2LNK+s7cCoCL1soWdDUD5AoryY7JE630K+ZiFi44p
ATICyvIw8k5Lq0tcWMDrEGZl+04YpUMDJXkgVWR7SI0+eKAGCERSxu7K/vmjwFywqHIFy+0zIf9n
3x9asIIdilmcXnYALPpyUA3uYujU6oosplkR222ejj5/ih6r+JZG9KoNCdbuR6nwFODHKySSq2L/
aGrRdWiGYeMfMGWhcoXfasOuc0LDp9/11SmKv90KByKebOpP7C7egzr3wPOAOnPPBuoPnpVvowhN
LRIIHI91oc5njk2rYC22wdEuarBgNnhaeomhujnu7z51Li4N+yKKNlzBZhvfz5mefh8uDuKA5YnQ
ePO/Bzk8G40LD+qt7yHXCjF+EkNspCBjjLdzLLooKipUIYeDkM7cBc4FmgtUDMqyUJI+XXkEdQv+
dGkDqWNWRs2Gu1UtOZuNGq6bHzbvpfieSHjCWNeGTA0sahktEp7h21xhjAp0TAgWKzsW+WK5H/CP
WRlRtEa1AxfrzcMzJEZBM7Vx/E0Ggz8KRVe6ClY9FLMNrztOlxQ2RMYoG1ubVZOesklw6a/UHDIn
YPIe+UawoqjlZi/rOLxsycBSnJ8TrKhBR9zt4Gm40tk+C0wBGUezE9BO/Aq0VqCA7P2SZzJoT2Sx
phqkyqRiTdbQf532LFjH8dL7iHeEhs8rIRNtqp45slKvdpblAr676Cr1rFPWhUVbqlmnIhNsLuEC
uHTOWv7bg+x4VN5ZGhbsDJBfc8jV7yyKMsVU0vxVA8UJi8JJ0hZv4s2xFNafgLmdRLG4tuif+XgE
fTTzNikYfkfmT/zBOLNE1W7+a9Alsz50y0MjaaTKtW7k7eLtYqAkGZxm47tpf4rZfxx8NrX6MKkl
UwBWtc61EXObL8Bx1wnRu9+GNSW2pCU+6gh0NPC3j6gBjErD7do3QRdt6wREPMk3KKncPQKKzH1h
wCZYTlBoo75oR8/+Sg5gzhJ1oxKUX2amzkYnNlmjdPkj6c/gHh1rx0L6eS2/3wSAKWecfTdZxO0y
kNeRNiasWXhW+5MkIW4iHf98NcT8MoqndKEzwjncCj3Tq3kn5ir0EWg3HeYJjJ79h5376GkjOfJO
2dP/pZGBi/olE3s/RkE3cABAUnoc7GfGiMK+xwo2bGnaqKDAV77jiYio14Fbrxpc7/TJhXHlCRs5
GIt5hwzYCIW7Q58Dql3aRVAdKt5HXy1OXSbbTqGkAgYxS1FPUNyh/M/0kduNRgjMFPhF5DBcbAXT
GVutChYiUkBU3L9Yit6kMDKOXQFoN52quDHLrF5gOATR9taGpEBIuOoXAtvA13TLXYsTfApeiTVM
RBjDiho4eGe64whTuQTBX/vPTAiX73774ysOhZBdtkeyNbS0fBfZm1tg3AUZhaw78Gt8CCiVE/Od
pVdaPTRyvmrAc87rfCjSgL4DUjbxFpSB3lbOjki1j03aXjQOHc+LglUEGH4gD24o0EpXY98E2log
3FpTrg94Sl2t/K2n5w6FjydWhaZvohTB+FzsxQbUThV58trkWUT3Q3ps0qexrWzXlbT59IJYHJwT
zyrKGgEUkVJSu161uvL38XOPVI0yvGabH0Eytjech3Cz1w+vZF7cG5GWV2oD7MoUyRraE2cpceO4
81JCcAGR+MtpoGj8OlhJh0kp8cSHdJcfHlS72NqbSBDctot24GGZI142WEQrcCBiPncILcTcGjHQ
2JriORacyYmURHQr+h1AmWfHcbPPCa6MGS7rxCwemhc0EynlP4tJ8FKY141ZKilw4lrc1TMdVxbP
OPv/CeasUVzGHi+Vbsoe2PXwEie8QSaYWXYpu8iWvwfQfbscb4xT2W7xl7nv33w2uCtWxjFmwIWC
uUpImkXbYjfups+L8BQN0Wu6BjXzbHzxWYcqTURuZMac4r+xbdAM+gFxtLXOCbCPDEVYrkoVLET0
a7u2mJQUSUlnjbhU1HN7SUHcS34Dn7N1LZTYXcOhinXkJ0bmt/GQrfMR6KrJ43IWEfZf0tc5v1sP
jlu6N4q99rxGWpdTRLoEeXM03NHMi69ZwAMMJgucxqaZIfxZHqTVH3sDfKi4EXf+k63rpVjgnB3z
ZND9pYRDmXbKeBolTNk/xcmKvmqt72ENseROx7feOpjC0hrRbHWm8MU0fOAKZ0mwzmy5NVrm1qU4
mmriYLfgxzSTeEvlz3Db0hryuARDkL9svh22Q76nXpJ4J63wk/1TxDrpaSTmFQcxBXuPEB5SGGZl
dWGF+T8WsYvQMS/dwpLX1i5oG8Zo/7G5xDfF/jAB8sGManOVxIGGSXseJ6pynNY4eCiZRm6sycoB
sVU+/+FzQIhbCOQ9/u9f77Lh69nDtQ5LNRfj65pp413T7EYuI7YtU/MaOlfoMRQI1ay17ochBxsX
eUGKfPDp+/pv7JyD/LKavlfQcsGEAgyO7+ebTJtntzQTtrNqdY+V6041PSUZoasZhSrlDB+MujxF
DkBkdHm8DoPcZFvOx8yCn9ZCaNTU0VSic+qcHo9vs+c7rInbXtte3m72eIolMSTUTok6pr1M+G/c
Lm6X0myViJmnN5BDXYeSBqSsYSPDe15Txjzrb3q66QDXIShrRZ4wW2lQfU/y6Tw6wXQf25VORbLI
rwmRHjeQorefDDNkksUaU7KOyMZ1h7CliBDC2jiPsY0FCYpTQKoXeNx6aau/hxA4yC2hNzb3tYC8
Q0axystlcooZOWcNQduuzYQUV1nRQk2pq4njg3e/GHfGQ5SSPE0DNFwJB/ayaNRczXTkfH6Y4NAl
s7yE6AvDQ+GnZtMPt9+6ptyxnoPOtoXSqsrkEme+Vc1g3ShecAHeE3gTfN++1nwYDzU9WagXoSmS
FzA+80/JMzfEQt6DFsc7AB8OGbINgN1+QtQg8XyqQ9SLRH9X4TmTnroMx+cGJVi7qMiQ4A6hnFHE
BrELHPGwHDT8Wun+YeiRq4w4SRBhfDOnV1OfVSCY/hTI+km/iwcYYBsDVD0RCCXCsvO7J/X+Dj50
iD0+jCoX5Bnd1Mzk0C5W8BZEKlBrasaikxFXCqOTRxyhSeAg9dil0AF4yasAGw9nxbHUG28lxBmf
bjR8DZVZgcX5L3nwQrlmg9WyTXvNJ5zevydShSmuvsf0IDX6j72CjUZKgvkBGDydIdlf4Vi+RnyN
w/HBiCL0xIxLENym7JjDjyzw9mJl/D0T+vm2+hYT9PgQr6TtJc1gOMkbSl1bGvFMyer134Bz44e4
1XIHGlbSrswYgz66Slt11IQo4+4y3KIrFwK8QQu7Xe215wmbHNUgZQUdwft3X+o1BYhy7dy9sfq1
V7FjKeI//qmr76J/wC5sQWxaiMuTeqIAmfloEVbRatZSVtZtOJIjeh2mhsJ225UfbBSn6j6131gv
fS+AeIirI/Eljnukhamve2FgoP99YMicyJGh+gYmkYby5Z5uDfavut1lK662vjN/pX38fJWXIdIK
WK6MZhD/9z7DNhysNgji+mEo9y/fCFUDMfmuG7NS45l90gmiuOPqshegZQTU2IEyjU+4xcYLu4v0
vzNArlGlftMBRc8PpuWBDLmO1u5SQoRLYDoEB+Lc9cFIt1vSocVg3kGJ8MGTNlUgx69EJjiJXwFj
/1RWo0OOJ56BvLFA82aGxshzXHdJf+oWGFO6imgErOJtzg9EoF0iys4csD76LMB6TP7MsbRHSmcp
fSLm7LJIcf76Qc6POwI6rsXFwREYxF+Z2GYgMw9bVWJj5veS+Kd2cw2cU46TFwmw/nBAmTZT0yMG
3Vuk7tdh7xYNdfnaDEIsmp1+xG5tWXtPDzKpswuoAsJwj0nwJ5IOGj9u1u43wXGQ6CVq4Xe/92q9
x288wos8CNbr028dsLCOZcHTefGBPVYkS1PGEWt2mU8yWvDUkZFtpKqubJBsYiMWy2kWmcL77Ok/
8oUMNfKJCKzlzFcYjEtVhYlKg7jjundvAvmViidjQP+BeS1O8zk28ybfJvJ8LHdOEW/BtDXMbZIr
tWqaM0GnaAv9iIRzRDad5skxzjQHnmKYJUGEm2rc+jq7+LnJ9HrIbZC8xdTCVAUIgCBi0tCQiCoy
hs8cG2G28av5kwhw8Wsy/hT7QaguJ/zW7OJDuLtfH59BPVCkWkoJAVlmiLAyFICF2/4iZLgKRccO
CUFKtmtfqq7hAJi1RuPHioN5ynsLZrc46/fLqojb/pdyoHwS7ENXkKbcerBxL/iL69w6zpc+QeV6
0u0hW6S0wjprqP1+AkBk9XUm/ghvvyIE/wpJ7m5gWoPT6XVhQ/IYYYwjSOgRD1LM/tz9GKAJ+1Kx
yMQPlM39ijNWZ8cEI59qaAsIUs/IsuDpps0Txe8pdRIIAsv0O2HHkfQNwPTON41i8S39rN2djJ8r
C2cBmtcTAFUHhjpma2HR9uP2ScfcOv3Dd3/V5zDQ0zYHY8it5l4ohVPMwIu+U1XD+qH1fs/wwVFW
yumczSCXuawmUetsv6eBFEYwELSdqxz9Bd4DiyF89OovpriWaDk7JB0Op1Jn9D5A1lco8v590twJ
m3MbMlHEVxmbjYXb8WvhokdfWtEiIZCfWeUMcPq5YxhtqgKydcqtC1BX0Y6HxFQpiwnUn1CvdKtc
plsMFMoW/2BRcwJoK//cGmDH3u6x3gYRpVJqrDMI9Bsb5zcpg2KKBEJ/9+Uasj+paLLis6x9lStU
wLHIVO+3p2gltXMS6D1rI2LyzvbjQ0enhtGATiYHLCJcnEJxz8pLWk8qd9fgTS82TWLZh++MvKxI
K7xgxxopteG5Fp1EdZkwnYjCv9o0PGnRiEFSBJ/hf7wZyrqMFJA2loezrWHaIyo70qq4sAQC/4fg
/KX77eID7YvK/fotxsdb2mB3F6EMQg3hjbEgx+2/RoxjG85VCpVj1i9rtQYEDTv1sc8Gpw/gyxaD
mpmzrPpmHcO/KsRpadX+AKsNS4D5UCSN6Shp9YQHkkujN2k4j974xLmQbT59XjlTR5JWRR1zfBQK
SQPdfMipBNCOAlwCUL1oJvqL19JfTrA8T45acKfuPIlHdJWoLrilzBu18w3eEyev9Ti+V/hKcqDm
RYDtPcCTIMx8tWgHHvLNfrUCdfRedxD0bt/s5cTJl+vBSckVCSya4XeUHj/OP15Z4AIntjvEe6o2
huBsU6bPMXtlflYfkiVGLIt0fZLXdhsBjCpZASI8SY2hws+YTkFnCJPh+BaW+1CTs71mor4nqKlM
sMMz8eegf68ymWk5SCx+emnXM8tIPqOjKwxBlmvm8omU1q4FbKNkac1fYK7BiIY3EHqq+ZQVSOWE
ev/+xy60EDCnuINJfXQMnK5ucUcZEkuj5yqpBNe/CMZuGb3BJ+Bom2iweust4OfFTGliupi9F2hG
yR81LWLdlKv/ImmOwG4fmjLOabFJHOi/RNAhcTXzjC/BEW0OPqGekBsZGcubwlo4aqX8lV1Dxmob
Kyirs5luMCEaKEVqf0q5r6tIT+ckacAy7I1ELXysdE8InlXHSsrjjr+L8K5kRQFK1hSw+ZFd2aF+
oK58U2CKXrF+ZDqxMPi4qRNL3lQLHEf25rjITWWwrBrm60KSv3GCZjYyWrfaxNqn/X1rG3S5sVUK
9xRuEuTH6wvma1f9L0rRkHT5OYsk+dr6B1nRtmhXy4Ksz8KtL7ItrdM/H78Pn00qPFjHJNom5CxN
VNkkHrHsHKsN+EyLFwdDiqcu5sW8xAB10+hXwefzO5jQAS9oy7KxYvO6wGFohZgGcat97tIAjbpZ
Y+krEes+CtFsZKCM1fCmQCoixLF1/1TQ9fiEwu2Un1z3hbpxOQATKojHJfT9kSBxPbKSE5umsOSn
vQd/Q7Mi1YCdUfjxLjjYuu9emU76Je0PhY5fzkXEXiTFZkDQ01bMo09/h7icgSvW0ALVzf0V+rjr
+omROI6lEZ/eERor1zQZ8juD0eww1uKrfxTE+P7Nb+jywdzK/OfMFRTF8Gv5QlEM5kukzRxHQiV/
b8O/qvOQ3USiQS/BzEQWZb1irj6WzFD8XaC0svNdE+NxEZkjKlybnISkDu5BE4WGb7t+mymVzSre
DVPkL/cHGADciy+HgaWG2/lQe3M/tQP+A1MwTGpljlKxeJx3hRz+NIS1pTOJ7dUCi169RCeEuvir
tmUrr99GLEKTmNFOdCT3QCk0qX1aMYXvuhnWRBCWMsN2GGLGZ/PapAdznzY90BABvyWgj6TzDprC
wca8BoMAT+sTMOMA+uLWDFxoNnpQWmKV3ktA9blQQUgduGutagKTMDDNgNqkBC3ONeA/JRvmqjfw
Q7I7fNQFCEBZHMRiZvIozSQd6+qXpM18qRC7TzvRpRfHiu8O3gmmyE66nTlG58oKz+pgKbEPhHlY
mL5R8hVynOq40GmLxfclgRG9iyny5rZ8i7s9p70yp0fbW7XekPLMlMDAEcKBdgFHR1ZodTSBuQfA
TvynpjVehQyHhCGKQ7rSghqG4KQYGdzQ7stRp2hmgjCwEBV22JwiByx//mOItanh7UACRROGCDps
VczAvBqVF4k0w8QiADVrx0dk4HpTXdHukc8XuF5Hqzn1l1I2u0U+VqdDHcBRr+6uFzQcRQeERWxL
rZg/A9yTaO2E1uC10N0sjdzNNxCCylvuev52zbBmpnpsmTH4dd0PjM2yPGQPs1tiYtt0iZkf2jVN
rMY2ywdOImgEOyYV7UEZ0f7yYyNooRV+DQccIs/ds9bPBzcYmgzjbBER/Ug7BJvYxrJo62te+fTO
F6PinRp7FhIAGCf5Oqta/h1fzIXLZL0Xfvmvz1/YpGDy8hrdj97RllGvvRqPaL7QPGsmOblAxtnH
FwJUrm+WTEP4o6OG1pSqyz0t8DmgwiSub55/WS8RaGoB7xWfHCD2iQC2AJeuz2t+Qzo+ShhB2n1q
nHD3Mnqr/BAZ0AKgFZr4QyWSngWE5UFxRh0Bx/xIQhfbDtVeZuHAn3WEEgzszIbOJ5ciSR2VthXZ
plExAfgi2l42kSrY1EnGgc9Zex5+9C2ybAuC2WhR3fKAo+ET6gb+zkUZaXrJwEIDaWWx34ftqiSG
Zp/vMvsD4GTAFighcEm3ENeVUh3lnRxiMW5DC5mFEZa//eH+g8/sXbKLbv26xofIO2IqPxTd54Jc
NlhkdWHEB4wQmJG73JBS8MawMSh4FJIaljdBNPQk87fsZKIT4DIc86GaHTHHSC/I6903VMlAhlZl
EY/yrGEsEGeHnuMNio3AwZeAHNALjIFIMm3ZmrdfvMZBeMV4U9e7NZFdhnieqzQ7zMO8pDo2BVFW
0xQhjA/XyJR7HNPoPZZ4HnIiRd49bcQETI96ZttsGoKJGuF2jRc4JXqHgIBZTFofcNGP1m0VD3ve
euOSP5BWTc5UcqqN8G1duVDGu8GIZtemuzyD5T6bjVZhfy29ea1pVZd8YENez6SgvYKp2TcOmIZK
iDTWdReKybXAGhOulDlkV7EJqdYbQIXuYxXMmK1bIs+Ur4SGSJReNc3UkBOVimdDXkZvoFLYEDCB
NnEc42evE0DlTmNnuHVZkzdjlTrj//Q/ItVMR4wwDklYw4701+rh8uFrrgl33CHEOvoeLJOnaPhB
grrG0tUgOOVS691DRpcW1x7dEyRqKUWQWqKuvvdwVBCjDJ9YSagPN2vIMkHSn/3Cv3+EwnCMliOH
a2QZrL6jrRPpj+Y51qEGD3P2vLGzOOTQwjFi1XBLsGqt7tOvRt7SbfpBZ5qHiRByu9cWmY7gykXl
9vb4aIlfkFyeu/vGeY5YEiHZL3KxvFluxE92P1RXiHviL2LzE8lFxnKS3YVM32Tw6BcxOdvJYx4j
gGDesRDNIcrbp5ALRF4wkoO7WX3OLDB55w47EfwWi9m0gtKpWvNmj30NWEq4KcG4ZQpQ//PiiAIv
iN60Y6nMtPNkoXUB2TNFb1FDuC7nbHvwXGdVGUbb68zggF/Mfw/rz0kc6pn7xuLpRfEehX9aJH20
uYqpk4Xp2OfqiKPM5gprZBrgF6OnvVbcc1Vz1zXHKmMUt3QwC3anznVgMLfriuk68z/iILp+xDIL
0+erG7z+aB4dt/AXaL1fqYg7wBbuLWyI20xoKPptgxCnDgBLQ98+TkFFeYiu31phUCvhlcybcY/W
vPoLn7PCRNVUBDghiDc/7mBPlK3rY+xTud+4etCTqNQL+2T+oWqPR4Q3eY1lTWquSEqVvFgLbwYp
NTwt2uW4LyrvAlwW0SbHzhc4QwsEhkG3Aj+P14QMIJpvCdJ6qAr+MkwK/ULpm0QnGmYED6WeSfQe
eTImicV6BMDpb45k4BgAGLt0jYw8pX6ezPbxjpYQoy/PNgXoybnvDOnw3lAC3YwqWL/9/EhqW/9J
jnFgNiv+J4lm6dmgw1b78rEiHJE6gYU2dwycmQP/gpktLEKljB6xh+cj2r9ZsWC4mzolxjHLWG9N
NntTjZ3iap0bTYQqULmFmiIqvdotifF6X8u5pshkNlYbjmub94WyCZnEJZSJXAHbHlHqtngzvc6l
tUoqSamganVWUFJSRcUcmqw02lLGrJHsCjcUJ/b23ItvggiymkivhzAoOzliCpgc1cRhR9eZJZUh
5ChX3nTkTX+oSHFK3yXjM56CMadXnmURHehcA9ovIYcVJcbzWNKpEoQglzrFDzBjkHzT1xS21RKp
M6pp0wBeJ1isggGrNATd2FhSlvBrUZq9pOPcak042Zu7qmVMhSFMqiR6ZV1lNi9kGDGUlWsQdKI6
SR67mlFrNRpTPHLbNF+JQ75hCX7KaJLgvdmTDbzyu6xR+zZgUA24eXRDaA54c8qqn5oEMCOtRhfl
HuBzw7z38IO4FBiIfw49eLic/UCv7uJCByuTMtJajN2slUPyvInvE8Pza8opEU03MqCRA1gkby01
mq9s/6ERes97h7xesCEENDFgOPt3R1g91cLZgUbqPiZ19a6lOx0SQAC6a21JSXN2C8qREIqD0v99
bRrj4vc9vQx0nE6Ka6qtUoYEGRcEr1wq3tLEwxCmZqE/kvjDN2yMfWJbnPIzDy0AhaFksQqguFZV
d0gzJh86OZMgD97G5V9HfWE42ao8PnfJF2p3WtiDKZYe59Nv4S1qSNRnd/VumN+ZKZwHFR4KxfwF
7Pw/7fWre5/mm+YrxhlB6cbgrAxJTipWoZn1hj8j2SiqL8BMIS0LDdCxer1joarq1VlpAkrn/v+E
CH8BQK6mPvFqOKUrt5FsPMkw0IFeAeP4mHhhn4uOFdvwsWAqbmjy5uf5vHNYAWTXe8T0VwzpqslX
X3cGrRLH1aJg8yLuc+yL2EpQ9Mg4s3GEnjJduBRrNWSGyP1vCdeHUoSBjZJd7sb6rw6pCDWQEGin
NzWJ/4UJ/wvrC85jM6S3T1WNKwu+HOkiE54yW6gkc9L2AiFg3zvps/9KUjLPxWqXUDo/aifoZlqF
SSZUFHU59NvQNS795Y+5mU8/bknonLNYUQmD1RKJR7PngfeRiBCwhxGtpYc0UAvFbS1aDyK5zVp+
Y+nE3GWC1SQRFVosB7vIVnFeJf5CZn6MuN5hBi8BSIaSgZiDMYwqkCnv7yEVcpVmIbgYZzVVMpw0
5pBTxQKgEg9CTd+hGZpxpIfVuHVzkjl7ADcT5r9X2kUZMeXRitftcm7y2RXWBYC3jbhbwCPfStpG
+E1dMlvbzpHb/+UwRiPtftQ0zONTqrzjoTGGFFe6ixVHPM8X4FkzedkUx27ez+kDFzs0QgBrb6pX
ZgfICvoUFnO1Sq30qJ7UWENpKiWNPC5cswtlRRkh5U/Yw7KYuZ+RmPt4EIoD2D4Rnkrj8Iyxq//8
34iXXzcbzWsA8nThyLedrtAkboZDepNIeE9WLb5XceZ/RCovSVEjaC4SZcYNhzFqAWG1a/s3G7UD
mcTJqllL5cY6GMUHXKcF8q98LNGNG0yzBFlqXftKZcW+TQaa2EsLEFxrM/qOshawwqX2Cr968Q1e
khmoKZnYsaY48BvghrtCouXYcjyaIbM64DeAccWYaU08N/am7HAsnwMBPKf3q8wntyuPlCcmup8n
/kGCbScSjKgGsXl060beRIpWLC3kzWf+PEEc1uGQj3aG5i/ftmBRZveSMA3+JKf/vegDcV2ZqySV
pBKvsC3t5lV4rOS7enKw36hDS2Cf8CFIXk6D9veJBV87kSNrm7m8iPZIf0diI5PWNWSYksPvowiA
ViyEFwdMDeOKd7GWwlJUxovz3J/rkgywAZl55S59MZz2IiIpHoNJcoo8HBoIwr/nllECWaeTrQRF
Wf1wOZCAqFMXgOcMMiktj6Nyvk9LVObOs7fJz31uIXPB/F4Bmu9ShdDYC8Uj3PmIXx5b14NlHuzE
p2KP/KPsmo70g1Ppo+4x7JfJWgGGzyK4lxNMmO2Y+x5LG0tL6XynoHNGJZbtSq38MHkKNNiyJBrp
l3GLtpbT6I7COi79hB/pcvsd1r8Fhk23XaHcxvD5hJLf0Bu6IAYH1jwaMQrXv8Rmc+inqIdicO1s
8xXImsul3Zr3Z9aM3TvTChUwgwhGPK/McLZ/NDi7ZilBsV1viwMyqi5jl9nLL945sQQGnSGMHmAz
fUtduenoLK9Uon1ju0VaicD5C/ItwnfSt8Coj5qwPD7vxgU0SKbNDC4heEFBnPqkhv5SyeengX+T
69AqhTCS9bHX+HfCw95ITTJene4R+JctvqcWGckoJrSn53QibQAdL0F774tCoec3Sno1E/31qaH6
nLPLhX7LTJG0KI/uA3fuIzeaoV+E8yjrzNQ4GQkgAvbPLNPAS1P5JxONbxGR2b1olPABkRH4rWru
xpiFJdFB2KM+Xvy7Nc4CWnoq5JA5QXJqIy831b1rll+lHXFtVU88e0W8lmOfQPvs13GNgnFOB0ax
ckyNS7Rekch9fK4I7k/2YSqIwFPqbjv/FIu/HaiiZX2XhEzUPbcAXDjdEvTyUIY5mfJQxpLxFN4F
QI3Av/+LnOQujg5+721gBy8zL220CYGoGbkR5we8iRW73kIFnEOaktR8NKoW7ReXIMaD3sP9i37Q
vjXbqikK5TXiSHjmwUMWxIwiJC362AdcsPxg7YjgYNZRjQAIDHQLbgDEoZDCY6uzsLMsb8L6LWMu
MoibDib/OOVDHrSQaGXPdt0uMzrAY/rv5WEVRYSYRPj1LYV8+0U+/qzYp9KT6qFnjpUlj+quG8Gr
+vKOLlY7v2opR5G9djKUhdSdv2YUtK4S6wC0afBhz8PnMR2LoFGGqXp6KO/jpKisMFwMS7YQCqQU
Uifb2MNv+cFbbfamE1qDEZ+GDHXovjspYj8d9w5AxhqQc1LPBccH0WxDQ1SLxDxo+0HtAVd6MQt8
on8v8o0dqhzJ9QnYevSo9YhfDCxEjFrMf+vlhUCeedoAJbTdOzGv/x1DaTbByKIRVFHukMLUEZBP
MAdMGziJt7Jt9HgiTRNQYcPoho4POMDkK/t0bdouMVVa7sulK9F+fHE6JFEvPtXkPD5RbCWfe60C
ZNridG72S3Dx1m4z4Z8atVSH6xmbC1O5ehcxCec0N8BRExH+EALs2nfnkRH563Wtxnm308Czu4MK
tilEnRQuCquIcMFyFkTBx9uFDXbv9JMn6iYAJ+cOCmpMR/sVHxJYIAWK3ng3PH8suCNZsp2ZM/dy
uTgZcqnnX3g/7aWGiqXoT44lQm7Bo6dQ6odkGlNpNWfr6rgPRQPNUEk5VWwAdq8uytmk6tPxMu/E
CDmoxkKPz1QyLoGGnii81sTnPy7f2O1+lK5/Leu/499YAJyW6UdkLxM3OZk/184Vg/FS9bfu61lo
ZUpPRgNsJQasiYU3nxeM1ZJB+HH65xXhpuFg505p7NPLznVH0/jBFlRAsjXNO+SjU+U/aCAJZdC7
FrhrwwSjlRsCpYsDu3jOZMhOgGEWS3EGGPP4OZOjOPfSiutmQeVcx+GLinAmfRCmvS4MPS1jdPV5
AqCL0Gh5H9+3H5SZDE5hPBk4X5BFIb0e8rQq2balqk0ji3v3yAEVzemivHjMTHZUgKOtIonbuvIW
eC0L0fl1NzExcvuzHTmCK5AK4trDisXxE0+AhWNOv0nuKpdo0nu7tjcJyOKGC5JajqLq5dhyY7Ns
UqZqg5Vez89/hR0uiGRjfng5dRAstDth+w03yyQ2IgM2nW4TTDtUp8DCCGu98V5yZmBH+7kmXEHY
+JK6LA/6jbWiZy/ZdfS4gxm8nbeRrAkMLNEHCdp1tS7iqSxitaUU2fgbK5cTbTERDnf1jZtjW2/t
mTk84XVuRs2CqEzKJ0jjDBEl1uCxH9kvBTBTxwQeASTYMxgspXaQke7IkXKtxJHwJimq69JKyD8g
fC9SyAjQeNXhjieD9e1CDfdlta/98MDz7Pa4DiQOxymagqV8+dOOpSFhN5RZt32TavrOv5SYEcIV
iwfRI3r8y82QSrYCASuzvTwScoJzV4pSbq06tw42QNNl6t+WvnUyIDMr/CWgkXUHXEmbRm+YBxSa
wjUdRNO+TY82At2eyvtbEJ5mmVD2pncnMF3SbjW1S2XAKO/2cXENUm9ctmmhnLA3VekghyAkib2h
vFLsTNYzUC2b0IgkMYQ7wh8Yfp2iDZxrVhCxykL6jPuY4M5sDBzUbcn2/8CAwixasqEVap2Zl5Id
UJHVTcziPTGjOCZ0tp/6FdSUl0GxYMnv8p7rxYMXoZKkqphCrFEpSeR9bGQCsrN+97JDlrPz7oj+
sxXisG+d7XKI35PYu1Ine2EtArxUPfezFCjiQ8R+qp9tAaTEzy6k/JwWj/gqLQaiOHYEZdkK+yZf
+gT8885Di3R4ACYN1hUnCl+qPRnQNUWqIKIlD+Ij8GPjGcCoi7JvHT10WoU1MAK+u/jHLQa0q76A
jiWPh1N1bKipkpu1W26McTyvR0t8xEEOICIhj5GvkVnp/+9cm15CWQNHmmwtoE4XW9GH0J5c6wex
mvnSQLTyTrZQKjJz2YvzmI/jr5EruEElsz7Qsk4vw5FeUALx/+HFJDAzeyr/JhY/t5j2YDLJRQTA
OdkyJnPbg+hApDgsOSQoNBm/jbGkLmuRc9k8rOthCeMJxLj5cJ+g0KVkPlNs1EsqUjfLBLxqmfCv
aRo4ABn1VMLzjT0h9ncQrmiHmtFBWehRMbxPgQdxLFRbXlNTsPWPvsaDIOgErqvEJqf2DoxBBY4m
CFI9fOUp55Q7MQesUaA1F7Ae8wGcEeN081iF4Eq5lM7KJmeBsweH6N50hWTV+L+fKFq+w6iU6/rV
nCZd+6kt956vlB10aTwMp+XvRNl7J5EiEX4+Dvqcl963cnA9HAwBP34tLp5fKILVx7yYRrk78ObF
CSghlDKf/FJaap/b3XF7gLV0qrvB0/aS+MeVYtA2S5xb69R4/q+UQ3bWKItr+X3HZy/2Nn33E4dN
A65mobEEvVtsXw5po2MBFzhgSBGpeAXcBedgyBseiNOAM8PTZuBwxdNJbqnfRn+8MK9+P9XdCtEj
0VBk2Ih6VQB+Aeo2dmdolAi52acvt6p3/gQPpKpFFNvcpF6IVmdepv1GSc2s9R3sEqreUqRvoGDl
K21UTfNX3bB01mFXN4/ELGeSsgEpMQxxdMElLxdBfckvDtpotCNFlc8v114gxcL26nQEk5GupQBo
tq/XGV21iL7FK3DBypjjH1PU6S+Yk5aZzXE9fQgJT9STmpTCPIIeDrsk7dQZaFPmzt0IiZfF/mFS
jApVr4F5lSbgvx5l5/te9EHe+C5/Rz8UxQad4fAYWzQME4ndsBVTJHfihA1OVgduSEhla1BrXG7E
k6KS2/UGE6uUqkUnRrYH/TmJ7YiyCKj1Z8MQkLg9jmA/V+jFHny1f8LkJGlGEzUxzFL1kgcoRFCE
4143hT5hGsmlG9qlGl4/RZt02Nyuaxa+/bduFOhWR/aAPwTykMAwiH0e0ETKT+jugQRi8K+03MeQ
BtmGcF6lp+ANl39HGLD4BeKs1Oi698D/MgWcxmKZrp0d0hJAtF7jA9OvRC+g6cin2xZ5S2TECOzV
UVMsUnLlJ3zuv23iiNDEWV2nxzLxkEMoejxhQkt3JaEcRtjyO8wCmvddGZbwbPNUa8O7Qh4mNzfS
ijMeApvArNsDr3B08DbroYH7xKSluO2u5nODk3OkqVy6EXx0g5SJ92WDmaUlZ6NIFIDa2PGKM60h
59SvRfTDPKjLDjDPQsoDszI610PIlem/5A7BAJ1CF88abmtG80l1ZbwTaxmpIl74iKfr6Oxb9MDG
HuytI6GUuvwil1D2p1y+nOk9k4T5yxI/0ZoQxmzsvF25c2jm+0z90cVxYHdFBiZAAgrk5wHoPa38
j2jLr+wlmsDvxatcPml639iRz9fTRyNPbbOXmm1IGfoGbirwPemmK5FFZjYEl6moXRLeCVGwiTUX
cBANCM5+7cEXWhAiOJsUXIIzKLZk0fCovEneRnNyu8oGLRobZMUTiWozd3KEQZQMl8swqIRTpatH
AUX4u9tj6y0Pqd6wE68FEocpbjxfAqSdUNw2dQRNSATeu7PE9Ud59vGC6rpbI4QMCbpJ15QoV6uo
3VgWeb7U4NB3TplRaRwgq3RFtowj6er2AY7FZtLhztTqn0wFWHE+OEa2FNFhtW8+A9OHvWfjuU+U
AJSn8pYgxsW+GGDKulV/J4jUQcmWnDZcoxKYbgBCX2okwmxF05GlDVTLb4tvGB/yuQA7z+7N4VTp
JmYOnMrLt7rgiSNEn/Rqp4f1egNbpfwYLgXCE4rqGOwAiOM0mqqodf/KzNneLxPqspg02xN77wDX
vbOjpFagqaZVzzETkumqyx0XfLy900skEmk3ayy41Fx9Onim3saFHdXD9M0YAGKWRNtN92pnr2Yh
HVxYjeY4IOeich1UN+KybyCm/uAF/l2YZWo9EYPRKmz91GO8+9rVorejTWaOev2cSw5ZAlf1tFXn
t7aX+7Gq3o4KFlIGtWkzy4G3NdxPmcy4mVLH5AjKatn/T8N8ywSFCnIyX4JL8Zoj3HM7su/D3sa7
LISqCJXEzIDBq2C7HjvLCPWjK4hue7n4FYi5XPf5v7BS+UbRFwOXoKgWFVXTN/nwGo22+P4wtqOp
MnOlXeVU7xePtko39ukr4jtdD1eUwegyJb2cQ2B/IjwZVrfNNXyW4GJVWxZXCHkaXMo6TJiSlY69
w1qD3vjWapvEOQeGDW7nhGZ6neUdE7xOpO50J3tdLPFUzu+I/vWN1xcm4vCT0c+AbIwy8KRPG+IP
ueVv5urcijVSS4eJFu4MG09xrhK/OFxgbkFlHNr0i1gEWrdJl/gQdRqQgblTQ67zv5ALkwt/B7NU
j1rlJ4LikBh6xrji2tj/dbHUBVZiev67+7+tzjIae8yFnketUbE9L98kh+u7XewiHjfpuOnwRM9n
PDZQEqgz9zkfXjCNcC0AI3WQig7KboCvZTgDlfK+qLDxKa/dlm9ywN7Gn6E3qJbl9+wBxOA1DySR
mqBATWZlqOzYGV9lb9rm5FGNc0cTOUpGUx/V8tWLITbJdLclSbS2PTI6XvjZRKihmLBumO7YJpgC
aIbwiYwqh13Wk6WXUsZrUOKRTOmluWS7a6BArI5bvjIxiB0geJKZBlBwyvmA+g7wNUa7DrK3MTg6
NSyWjUD3M9uwxwJq4p4QIVjkmvq6iWdttv3AYh+NSjMMM2Xm5F/y4MzDgH0vSjK55dK9sUApse/u
EklMU9Xw0LNz9p6kHX2vI8B6i1/zrbMOdd6PMQyuSgnFEOSopLg0cYG+MGKQCFfDq7MVYJ/yRl4I
u9X0SUR7DkMjYdnxfkBvlb3a2DHJpnbCj9eDq36ESXiTcL3laF7JdP0nm4zGfHpCVALZJzTKW9X6
KLEyo3eNVwo/+xqB26dTVd0p/k/MtPeOsLyN9QgAe7s/+vyWDCzSz4nmw/5JeprbdPQXd0LMu4CY
jbGXFFflNEmfaRyik/HaRGg2o9zy8jsa3AI4iNfP1Ki4dXKxUYJOt9GRhTta9kqWL+M5qS0cb/20
px+I+BAYbt7IK8B66l2qF7QKZWwO7F8IPuPnYARa+toon8UmiWS5R3UVu0exnL0JB7M0B1jhoMAY
S4Bx3eBggyt0Uep6tVwgTcbSGSzNqBtKsd7vcyVpgPtlK4+FOX6h8qN3IL5Ntf4pFzsxs+BTnzef
/50ddom1ILHOeSLJIji+y41vfTE+1dnpJMtXOLNNl8WeAv72lNTonEAdFpWGCX3qzHntCbkuZ86I
N4mM84BUUKlUxMJBEMCsjoK8Ktwp6ij4K+XoD5mqDfKuSV1EzbG8Cfiz2OmOryoAySMgxb25EdUh
e3VT1tsgbccrQET1iHVQ+kTPaIxU6CW1UglTZii8GX7uNYWk2+LxKBBPDhVZyuyu4YVCW8d+ZgYA
gh+xLkVSoWUkrMUgMI4RU87bAgzuqnyTKUf+o/vzdP8iMBgPNbQVH+aNUIBq8d9n4fqX03qspSuL
9MVBLpvUVXgjXZsG91UWfq2Ghp1IjxQE28i4xs9ldPetAUgxrlIoOFbjxHeDgXlVKIHDDpjKeGPf
isXrZBgyOelJeLUmtrzwITYQsnCWQU7YUOOrcy7Ri+4Dt425nDGtpUO8/95uSX5CUKxy74+qD/Ea
jgQOPpYUhbZodlaopDhX+C/2kF3yaCwCAPDAMV9B7165+2V1Ka4F8wXWvpgmkjqeD+JFbbQ0qwJK
N7JzpYNKFuT+3V6bKGYriAwNzBdRBh+C9PwOoT3jiXD+9p9p29N8Kgq8JMcxlr0H6CUx5oMI7PIl
rW0YkkTFgK3isMGDISDFcd4Sqyyv3O3yVX4G8hYD+ZTv7qcCv2PoGbY71c+v9kEUjF1wXWGUOUgv
bM+YFugC/5npb7+1MU5F7AdafqkrimTqRtG2/Dbz3hnc72LaCombQCf0x/x3Nwc3QRSHtH0RgmIC
vjafbNJw3I6xV4z12ib3QAAJnsOoM/crTMh6i3CGtF2da0YP9xQGoSmVMaz0U2XL2Da4OC6PJaoc
6Vcw5XrJfohbqtGPvkgYoAKbexxUzlPfQCBblAOQHoyJgNV2ondOxIJiH2evPO7MOystwEPtYRtC
cPTNO16jKJ+GqUXdviFcztb7rzgPzz9xvnjh/1UkmAi1NSxt+pdtll7coaEjdJrNSU1kaKH+5Cpf
Z2lKbrOXPqONbF3EWicNWk5GDXuBdFoRBqFqeST/DHkkDmwHrSnDfqgEfE4TYGkMDVPL9qJWlmQw
AJLB1+ogbagaTDUKW3tLsJt8Z9GYlTjFIVCSIrgcteU7ekdhjdmaqqer4AaQ8GZCZemt8PI7Qdms
vgw82u+EaXqfhaB0HCRdkZLuqv+5l5gM38rIrcJd/+Mc93b4AoKIL4EM41RSoB9PiNjX0JqmHTJw
KkbQ9CCcYqLbwjBnU8DW9cdSn09e0r72leh7u4NN9qpXCPmeDanYMuBuVOyUFaiTYXDUmrI+y0kX
hV/HGEYmCZX3wC4E6dP8l28yxg4hBo3HsY6HaGqglpWj4CntCYbMnptsqHeWHdAmIC9uNYnRvVEj
sx1OwcIgcEk2iKtjiPTMgnXSblYdYGJJJxzfW4MxGhGkBdpcJiRjfaPusvgaSSzhBFRTKQo0If63
EELTBVu7tIBT5MCBJqPRIJnqlxiWDvWgSgFMEvPEjQLgefOSzBLOSJsK00RGyG2MIpkVGfKZvBmt
ZZQa85kc5WejA6fismJjNkO3+Iq692A4+Q4htppJGz5UQAd03mZt1C6iq/hXwGoz2t96FdwF8BS0
Y6PtCXX2M3/B10oq+AmnXmKSCYKdce3RfDjkJHcs2qFhcxdnF1ldwbzpF9vWYFta0e31WlyYwYyf
iCOLp6IUcKR/RqZG+z6TP6Jq/p9GiDkcd3QOuaHouapuqWa6YvcQuiFIPIu4jwAoRoq+YNPv1adb
TvTmHsPIzSd9hG8d7P0Tk8UQLt7BDrWDrFpRxTkMkXMdGIFalnVrJQKeWdHWVGE1rySShMjA2Xrh
CKwy49MmSayDwiIoxI9qaAcNaJ+IbjW7EJqzgsyybQVHMvKpdeOAfyTKH2CPAm463XlAMFKGYwa1
7DNTNHrm/I+K3evAhvzq+5qqNF005c/FiPUrGA9AZbYp8R5BkH75hF8DVkLCKyfHwl9uiyjcETLw
Mr3CoKWbo0Im1ppaHAZYi2PnfTu/W9OTpW0Nqx04EtGVRNqChf54jZM6iVmMVNzTXtMlbAs1dE3R
HIIaypw4ssELWsuByC9N3EMVZaLHlL9lBi3tRSSCJfPMK8C25IOE3lmgqrJVrv725mOoYtfpKc1w
6SIU0zx3VgA6zlsbcF8/YzxNUQHwownLRpYzCv4/dHK3bCMhkeYyWS2T9hDu0PSSNzkO4+cHUvaW
AEmBP7+WKF2ETJu+8cFBX7CNwMnuRgzWNtcCToQdh09cbuXFtGh1WkLnmzMT5vFUQFtDtjJKxcEf
c86YLya5HgQ78wSPvfg9h1PTGcjM66rbVqbJeUjM4a2yAZen1v7QLW/KX8XvctPAOb0CpU7sGHl5
1zAXp7dSISwfkakUCEZHdHIkD6QQ6iMvOKCHIL1SED3xceAyD9MnBECM7BtCE8JQx2oNbMyZBz67
n47ZALQXOFRpFpA9cGyuLsX5sQbhnwvj4pUJFky1bN2Tl6OEmBtISsF+ECiPZ4/ch+e7h16ycV+Z
mt53x9MCHBrioII+4COU5YGqJDf//pVj4CunLuZWLPEnA4uDsRJC0EDAZPq8sEPPC9yXAizdVjbr
cUEGp1rKf30uEvzNxYzuZuhuEvygwUhubksiOkjjhCjXCB5jN4ip/U17Lo6PUMcoe46xZHmXRtrX
bPEuAbOCGmP3chH8SD0JeIf5q73iczgN7s3hO+nHOZtaZ0lrlx1SMSfy1BuiX0pa5EkFVPT9/1bC
LCC691OPDcNe+zP15zuOB7ZGGrFAqcPAXXQtLax0iUI70LYUW+3U5BiLzUzE1VBktnhx9bOu1XZA
vaZSH0kC7j5GHYneZbHNus1WD2ybS5wVGmT+gizNLI/wEqIZpqF7p5jVh90jTdDBi5C1n4c3tow9
HTOBw79rWkJHFmxGiQ61ErVDk+exVFG1g7kyjs7lmld2+RdspWQuQGUyGRjHKC8hMxEDIkTqaLvS
FafWF82YN6raSJTXsF7ql8rJDNX+CHU7N/Cion0jo7xzL0QWrN8YTc8EJXzGZaPqxQVQ9N1PzXIq
glCEA2Uk5ivqDqMZXDQKyh+g+7iLSbZxZSft5kQ3tfRQTXhsZWnzF+KR4LRt8qKUbg4l/LeKse77
AjFyoyB6Cl+SJvFKIB9LlHSb3OC5wIaOuCV0omKLkHZGtQkCTmo7f79yZ317dXYaM2Vy4pNjMGk4
MhFop1YLtaxWPO0Ip5Kp/nMxj+riwxEBpQtNY5qYgh7tsOs0wFaAoVk9He+di/0jdJ0lAZadbCRC
Gv9c3CDS7MEJuhl3gYj3rGfTU0nVqrSQ3sKgSW6lbEe7SrPcsJ6Gmyf8txRIHQaxVwjxlTWhu/aJ
NloqWeH8ros1v6UmMBX7Zwd8RzCJ70QPYeLdSQ71E60VRyf5hTqS+n0M0ymoEZq/SFUaih2E5Unb
OnqwjGEaFgzNdOz6EdKXrSfiH5dVQUJnuNTZLXslMd0xPGWF/VT7kK6eKr/CPc1GRR9XrayV+0WT
OlHYvYm3HSVgP/cloo8fsjzkV5W1xAaVT4tbQ/c8ww3XmKBZgRfV8JZWSRne9WIMJp1HHpeATgTy
le8HaxWYItqGWaIoZlyFtA7ocJiHux8v/+/R0evNQjuaoA8Kso2qv9ZoRcHwK1h96HoOtKqPCyha
lcOknvqG1QQvzcq6de8ObcaxFj1+UxKCriEZLaqOvTbxrfsVTHfOUgkARUVuVBqV/ywH4XAU5C70
CCGhsIjX7iryosv/EDBQEBraqf6O9iHjC2SFhtD2QrOsjyI6hnxQmy7UNotLOFNrD4P7DVbXllHv
YRh1CHYM8eVLcV5l6rUyMLS6hSyOXUe3jjuya+REbJ0bRuyOHlT/+tbdApBWw+qDi+yFvX39MLqU
le0kms4JSaf2yjb3H1hSWwkxlq3mGcClIBYbFYPI5c599V3gJdgtpCmvvqhbUHgJ1m8cjL46B4c7
7Rmgezg4CKsBeL+r88hySMR0bLVThSkorlRsAatIUd6AqNh+OQvx4qM9wGCd8IYaYvY0UcVT+Rl8
rpu6X4AkCFhipVQ9uA1jcJahWrbGs9M2oGZbTMISJud2GP9Z0aZ/Ua3FMwDkOX41H4ZgwSRKeFYt
RbCjI+c9VF/GfW6F0uraCOB48foWHXD680dQP0TRxszzuy2jPiyQsZ8456f37jBcrLb3MoEFXS/M
hKbi/JKUaMYhY4TthpAcVTUmshpCTJv5pAGbbeCO/CXlN4FrV+pNT9C7fZybojP3d7roTMQsFRGJ
U+rK3+Rg3yp759ZF9N4XxNqLIxndnRAKvniUDPYBGqK70vHcYTxNmTsBXyDVPcTHA62FkmTlbt1g
B3YlNWDE1jJltpU35L17iWX19XZaQS/ABA0PPs7GdjPd2HY0f4peZhMEB+TVxOaaiaFqy602kLKi
NbZfcSCr05sl874vSPFethNif6RELmbekNo+1fB5dCjRZbwbyY5yMXEkH7B6kYNXiUyAMQrjzpnl
rEKmPbUVLwjqiP1Hcw5r3e7yFt08ev63Y+GzbSixNSFaEig/WdHga95PyCMLqwDOjUVY/HexeINq
fZBhEquxUoZs3xqNIemwsTZtMdEiIbosQ7tVOeiY4iXTbMl4BgE5hrr0xLJAT5WNlnobq0QPeL60
dCfdg++aceI/00ye1xAjNvW6UxvMNRC40gLRNrT9sUBs+pCbpbIs5m/6n+qxwzrb0MMydyQgYnno
toqFH7/HmBCbHQ/dVBZb4G+dBDgqIJrNz60oCdcw51ixjRi2mhQaAq/XESl7QrP9GHDwYMo4V6Td
Gqy2I8yamOsjY9j9ZGSNdS9SpMzDELvpl8zLzRpRMBwhSyLymg7vccEMaY+BrfZ6DYbiKELmD1+c
0J7SYfD9Apil/q6xvemIv3aPFiD6bvNNKMOOfrMc9tPAv1DfAYnWCoATYKgSKf5FxGiUCIHvhvOl
LvjRJwIPm6tL5lgyQYSktRYT/JDBZFtw93Ykjegq9ShdMn4UF3cuhrS0t1pnkl69Qlm2WmNWO2K2
MPW7FZ1QCwUOaCGhew7Oqv/2xxpQhyHkIk/Ddhu6VOZow3Bc1cYhE9Rf7c6HekxgO/GqMgGMR8JM
AIDiE0UO8lsA29uzIPX8WGE1c94ic8uM5v0XdsP4o6O9kX5vGaVEtLnwbl0kP6TvLckl2CdFEOzh
yF0AgQ2a+cwRymPDY1xz4MVhVvMJnc9HTTMePmjSEOi78/RDbl8AL7NyYOEWUGJjcijz5rWkj8cs
fJpvgAvesMzCn3izODUkF+qs3KlbAAy1V9KDKqnbWOJuaXpq5s4TzfMGpVPkp5S9IioKZ09KsZIi
agwGQAJN89BYNHyGinzoTR4ueuEjZThPLennlO5yQOECLigdhEBcqCv3ukXr6IwSi990GlUsmCJL
xj5jsfOxAu6EcLuDl4w8hTT1bFqjoqKsngm0aYOHmwdIXtoES9BJIeGvei03MucxQrwmDuA5y6wi
jAbZ5crvThUI5ZaRwNzuL1L+5teHfgh/TSyicoX1JcKBQpvkr/iA3YulF90Y2UHHY9ZZf8AyZJPP
olui2p5eQYRJAmigNb8mP56J29v3U0U7V0eDotDZp7rkToFAa2N6ZCU/V29e+ccoFt9iSfNhvlpm
kAggJZ8r30Q+0Gcj+/CqLXe6vLAseo6gJ1m2I0gaj1HkVt3Ql7YNbRsOE3MgbfjNNQB7VMKEmivT
ZxyLRYLHdP9toOVC4qggiUdUDMONw6uIawXkmy1EzFumwQguhM8Lt96VZiMvog6tq9kYoQRNgNTq
Nw2gdd/VwXwEirZhqMRd0fZox4qtZx+rVGlq4lSYmHTwCZVuJM2i5G607/xg3veEprbUM9INoLoU
iDXBRaUMRb3LYpdIMGk9DG4XKhYP0LqYdgPMmonGJdQhmwde3XNdpEQvZZdiHFz7SXZf8yYFMOpT
aWe2WxoafOT4E/lAY8UyVUJApvZk0tZfCkkCp1mn33iDmFjHyJkWl9emqnObI4FM20i24VIKHIXo
aNmePaFStNExWI58RJ+zk3qeolZ4wXJoslcryxdw9cavMFgyG0S2gZ65YuQoltw6xNTlWneD4ZsD
eCsoVd9p9RBy7Ak249MUg1Z7BJ9TM0qnFkykqG+LPeaaJdhVNK+FBqgXX7UZ5SEG5eKPDzGWsIbc
EGaV68jVHlOYDFkssbs7gbKKxOCv1cUWmUTEsrgX1CSCZnH9lJLuqGq/TEbnzntOSeYX53ushvZM
8gzl0NYHyj9Fonr3E6ERsbXbbfgT7kz+A9u0Smw0I8jWi8KNd+dz69klVMrrWZL4L2821v4E0zEV
0O4B1VIVk9hjYAeAxRBxaFbgNvLgaZoBktnytwglB+HVBBQzj6EtTBLTBpcGpXPqDdIbuErFJEHm
wa242Ti6kTk5XcpXsb7IPUJ1GwaXU3d2vqAqu1NNXhibf3YAsv+BF8D1CJdQbk7u8yEy/7eIo6Cn
rSKIKxUYTOg9ZGzxzQhyE0Y+JTS6P1X+h82cwFvwYj4w6+zYcruRjQT2/U0j+56rGdknI/eD69We
lyqSSPD3BpJv+PNdBa+Tmm4xoPBjVdrfUq2lKXfBX6HTuftwZVt2k1fOtiQZ53IWVO1vHI8UJmgs
21EpL1QWXVs/GD31fShPCEfcwfG+EjQBV9flKqZsu70Is5olQfWEXljqNuyAtmySV5r2xwzfmvQ3
Dld3r1S+KUyrE1xUtFmNP/0hP0UU8F3Tdi1ye8a3ypfao6HwqA7vfxcnjspSvNoZDivNGrBcLaHh
UWQUQFNPQr0t1QexogX0pwfPPVprXnVYpAKUbz1Rv2vjyk37M1hrmc9NQobAl/kbDtKq9Eb2kHj1
MDURAvumx5/pznCkpE3g8IW8i/l2aYA38/iGTS/GnHops8XVCIfoC4E6+KdNPmtqqEfQxxpmcLkK
DG/q/1lg9ZYhkq/Fl9363gaRo3pFR4y+eSmVGjAAJqmqCF7TjV21bKpXfV/+L+E0xXTt5Hgh/sqx
eXieTExm9bAh+uZytcfTISyL9zUfnHUss4QkkbUJp7kZd2T9tQ4Tdq0vEdiDO1ELVsDURWwNGO6P
Yg4vxTyOdEO7OxHC09AHmuWN+52FjaY2zstqeK+GJjOs9tbSyKBsutUAhKq0gBKKRexImwFIfTze
No8jLrWz5+jdTpPW09EhbnxL9I61lhe5z+S23waoOK3H3YtkIszEyCLNCkYgOUOZNhwhL0w9cI5z
hEGfRXEXf5KT4KUF6gpX5dVMoyW7afdD2r7mGo/DZT5qTR0jGAGn54fdQqjLGZ9ITWYAJvRMU2c9
5os+4Ix1saHpUGpjtfOrhaDvP5A3WRr9R+RwbiDQknLuzHGa7D7GoZ1Ta8kBFrrvkAYY42faqthG
PqddvvNIE7sATfQ3KA09EXjm9ofOnwc1rL95Un7tvNztwyoUJQMV+iUm6wDAZ0pDfw8ki/pj9ba6
XF/zxZIT5aj9cXemy/uIsmkjTnYpcE1m6LviLjhyhDMXLNtt4v5Ti9byLce0X3v+Ply1a10btjnv
htJ4XFOhlyF6qv7ewpIqKEq9XXhSp5WT6Y1ZP/yCgb7QVPs52i1ZOFqZZhcaK6XdA3EG1BYcWDmD
uRj+uv5fmBRIJK1lJkTMF8IhVP0TnUOfQYmAPvLnA9R3UzZExVjqRijYrDgP25V+sY3P/NIj063K
WeaylvUAmnk/RbgfZAsB95IQSAwbjkpqH1ja/taO5YMlptAkkN4ftGVpmdxLIAWbN+wGO5AjVCic
dEEtiu65Z912QjmuYf2MXs3iAEh/c63nPHIBT7CAc8k22tSC34HFIplStoMQOGyJ/pEUwAvBtFJz
17vU7ZykvfWPBnMI48LLnZKimASxTjFEe74h5axHhqsyJI7uasZ9/x/8FvvHtZETHCryrZf3eYn7
i2KD5WvE3qJbi+c22AGR3exVVBJPCF3v2aqjPzPgWpaI/cSuyD1LZCxppp4C0L0OyAHtV06nJ6MU
eoi/vhKRcv/T453DkJAFikYdqlxyOBUJM4sl9YfbHGPeASPgiSIcVElL2azZR1B9zIrMm0XDtfct
yUdKIidjePkWNsdi6fwfr3EYY45cBGMOYDxQCjdPxq4CuDrI+I4mnGgvPoHOq2FdttomUGYcr6By
klzJ8VnJ08UyIZAr8xb0QEXRoXufu1SFzymGiAI25oDjUD3Xa1ouFvsnVjQ/5gGIeivZ9eE1vOKv
mo5dtxeUSZYrIBKLDqxpzEVnFG/ZN1P9Mu6iW1u90ghDwO7SAqS0thR7t/kSblW581Lr/X6wqSUn
ogspWZxE3y8aAw/WDW8L2VltDn3r+lo24GXVwvW5A9/gyRrm38Re4C8P7dxxySeg6Z1aeI9UqXa+
4FMWfJS/6yh0gOLL7TqI4ewnzMHWCIoaqE6t3RN4Ig6GYotU0EVsIElnSmp3VFSmwc5rEOvLuvCC
dondG/Fo4K7SK67x85d0z3CMtmQl1wug5ifKnLmmRadRhjYF3x/cUyI8/L7y8JubLto9ZhrAeCmF
r0kWEYfzxi5vG8P5qRXtHrhAoXe5PkP8pVx0MfO08jQD+qhqkLyR3PP4H/auW0sbzsUwr+crf+YJ
/xYPjRMDaV3aUh+76KJgs5yHZS8rl2T0nOeQWweT0ZgtEoWe8gaAztrqJvJIgcH7sdKg5QzatnEg
Fv/z3eLI7GeWTC3vTeKHzyhcPG9uy6/4quyWV+IoXZCQW5Fo9PCTkkVuU9X6YM0zY60d8L5LriTu
McXaMVxz6SvffMFjC0i73U93YaO1bHO+PUHkUTv0LcE6ER3/hQauJOO4og/GtAMvXGg1PHjDQjQ1
DbOiX0M+2JjTb4UbFlDpW/254ZeLN2ZeKT5VQPdWuqUKs8zNAOYUic3820qZ+tbLtMMGAkhdkgCI
6qqQVw1210rXWEZpe2MEaJIpaffwuvtqaQDz+wWg/bCU7qa2A/WPGVav0e+WE0ES9WYlhwsVB6Ju
Z88rQNGryV0uezcXrl5OxxrrMcVQVBRPv4e0aX9ji5w4lOFLdeDjrar2h1JC+7ZzWkeHaafWVu/b
pBXIjeLkHhlNhOgEgbOJ7ZmAVhwGAVWFszBYNtGwNzow9QeB36PLSmaYMFAciaRtAv5iMDaSU4Wv
YbkL0DpR6/mkRQ7VqZJeSKaRSIz4+EODy+rZWlQ4Sqm45SZhn9Yhs63ddRPki0kjOcB6uwr1OZxH
DPx3yelR2vQL7oEs4LepRtxm8BT+hCLhHIFhtQlvS3bRVu/kK2SbJXXbb4gA+x/o3h1J7gWvK7uE
dpDrywBReYil60hHdDeoLxekdR2My7FNu/e914md/J7FJyXSZhWo/pqtn5Y1Ucur+U5S0YTv3nrd
YMogV4M2C/SDjH4sWx6XsyuqnU0Uy2EEP4i58IlacfH/L/e4hyrbNOMlUETi9iItM/yUcrSPDE4l
aais0mfmBoMMRtemV3m3kJFVu2MER8Nl+SL9hJkPEDuto2oNtOhidiQZ2ohs5/u4AI7E6xuYzj0/
phOdVrgT5UViyx7WwNhu5SsfZSBZbbpzpmpWYZx7upmvpz3UxeEW3wDXwzaqwP/JQfil0iNVpR5i
CTLcEm3F+ADB+PIcl4xgz5dDzA0htkoYoCpRKgyxzPHIh/WKWMOjTdVJNCq1He0ioRekUf+Ga2yI
3x78VHp+l0N4xKijlfZcxXx1aSMm1lEUR7R2nrGCRvqLcR9Y06QApPfoJrt2jS4r3npSeg0TIBi6
4pFRpUNvgX42kRBKR87HPxaDC35CdQ2xa+EDnKzci4u6oLNhLYiEGlQSRVCXY+JSWsngzuOw/IUb
BX66iW2Uu0niR5pB7FpTrpm69CHczVVcPclYmGus3hOtqFjnJa260tZpl2p+nZXiAzHWPvhL1K+z
N3czwlvj0ZszIEr2p4xArwbJbHNIErsa8Fd4SvJUWBnLGlh6Z+49Ps0kpATgWUTZOu2/7qifteVE
SdQN1HWIQVABBOrlDQC1A9U8eHwml+DyNzI8FwNqs0ujkF+l0io3xzfuYnakADaaIQdBA7wxEb67
tsmsmCkuxq8MxCDH561ukmwGNtNYyss4H1O+jq6Gux9qMKNFoJIUsISKsRuJyZDV0TdmSurym6hF
NAMTgpas7HeSrX75yZB0CAUykB7yJVcFHE20IG4gWpBGjlq8S9RvtPum3D8dOpZG0Cs2Zel+X0M4
v3Q5wn0QHJxcdrgZYUUbRkrGqBycjsMU4yCeThD+nqhWcISurZEnm8Sxb64ob5MOoWLW3c/ol4Ty
SRNoFtjd17WWB/5AmVkQJ+EAcjB4vayQxvEDBiWykge2UOxzWkTRFz9ugBgWFQmvQl/s4nJHPPGv
GR2+VyZQKFAQktlkz97/tz5uGl1JNavVUclwirlAtmyQv79jhcrxxUEanR/kxhyh6X70JZ9A4Tj9
V6Zgfh6dLc/j5M3fvzmrQ8yqHhtBV222L06QB3cBykC4Ztp9pPR8RaWdvsPdl5N8oPBai9KLPBUU
eKZgw7NvCgwSCmLzbx9tUQB7UwtpSE0Nx2JJJ364HLhdwCN8TjabYpLt3PU6wnF1+rbOQL4OwIKM
ubTFCBrWSXDimTzX9kVZVKap2mBQHIPwEn0b1bFNLr19TtDZAh7x8qp3mZrE0fmAPPtYEn1AgOsV
RKixHwh8zA0BPjT93VYIurlySHhtdtyfdfAjffczDuXg74YIWt+PQ0wEo0Tjbvxy2OZdST2GmY3V
TeHQndjM4cLPzwgLvFPLT0SJ8kzbfIp4AaSMI3RRkOicjkubgyCVgbinyrftvSJRdPdfr8Y2mZgB
eqjrrwR4ptA1aK0zjJJSiczC28NbmyUQNikW1gjXt8E1DrDzf7IXGXFF12eq1B4kKL3H/TH40uy2
k6pjAFFirIyKMbRkeMORfVlsRQGHf8ixeb4mmKYu1rrS+MEAQs6oMH6x4ZrDaL4/kzCRRxZ6KV3w
VCQSHwlK+JxURQK9DqFXz4M+N8WSfqA/3N2XMGn0+Kkxt6lGMiAQ5RQI2+DiljyLWLhCd2nWwjnv
0UE5eLEQphcGaWUua2yfCqhLLcMplovb5yHYHEKIAfHpUVyv9AaunWSHMvkCVkf4aYfZuuQ2g1EY
S60jR71zLXOUSSU4jr4q3O0nIkXfokSxAvsK0jipaBr2tL35szVf8AFkDeP8kKG3rBptKapUeyCN
2pleUjFRsSV8AnZ8GcaGhOtkDtYoIAQr16LtoCy09UZw2AvDuTGSEILSruE19wCprFtUu0Edk0Lb
Q7xDClONbfFYJ2RIN7JiNdj7Ab6ycK+5LWPuNrl4Pka0LgkxyiGaA9blhucx1+w1109JDOVRMS7y
pmRxyBc6+LZXJjvrX/abzK4E90N5+9LL3+bi7EdPMA7Xd9uWLtghwO8YOP1KEysLS2Mz70KhRqpi
bf/JtTVdho+0FpsVdDlTAs+NkKScKFxvOc+dkz7TG057HaD13/WjaIT72Of/oWmoQdxf8a1BCmDv
fLRbN969B+L6d+QETzpUXqw2SYleT6V6XUN3TERPyqG950MUEMD4yawVv++IEfeuZKzkYVmHPFX0
+rygdlhBrdgwjdQQ9o6thp+YjQV7+E5A2NYzwg+BxFuc3nmRdAUGSyuxayT9JAPRVC5c0iaXLtP2
SE+XC/dEGMZIp7IR5Q8jQTilx6UnjlohgJrwBR+RkkBHKQayN/3+ja6fIS0ta3yb9y+w1cdd1VKP
xvKFd+Xo8JypDevNPwXIhueLiTJtdmz0jsHTKYZFbE/BojQJ8s73THvoGTOw/CQaOMYGIpSi29PF
R2ynZvOKzO0zJKyf6gCIthyPuuN87KG1wxfvxVI9Q+rDUvDqZ61Vh0Oy604tIx2b7HQnGMo6hIdv
e3gxmWfQAG6LQ0myQ0piFy3lRaExEQ3dRdhfS2TmsgKiXt/n9U4BDMGHderSHOKHqqrCdMl2FbCf
1IHMmW47kMtAMgRH7UZfCaTbMGFIvicRzDaopeeML7S7g/x9H6ms0jI8bIoqQHsmmNPT2JdYxgsO
MN1/C2wpIcjF4UmB3BH8BGIr7xauPGAkSOQkqFFC0jfevae3SWwWA8k2ZBDh0RlSseJ2aj3iBH/n
LXpRevvAjHM/6+qhlBsLW1BppgnLf7s00Gg7LElz7NJ/eU30eeNwTFuUdRh4ZQi3936aXupWtKQA
7UwO/348ktOSb2nCuKBaAm1UYu6zT1Sx4zqdDqLONgZ8T4jpVfkgOhorHWGX11nXoc1s4Sojkxv4
J127nTMyFhVTZS9Qvv/AQvx0oIlKPBZzVtDIFCM6ZjEizOUoVkAQR6G/BLFXEbYdYFvrgp+jPU+S
yeI4u3c0V815FEyf8XZqKEs2JfaieASdX3cIgXeyDoyj7CnPunne7iJwzU+M5aJ9MkbTXM/2uyVD
5RAA8SLtWP01YN2P8YevUhb4Xvfwmg+r68kvowPbEOuN55CF2RxgWrPHlw3RUcZiTZr/em+W6usv
ld+Zlxg2ebiBggEtA8rquLUwz7eT3MZo49Nm9Um4GKXooqQp0FNSv8pSl9dtjShTrFTjAdgT+ax2
AjDe0hphosuSPp0+L+WQeuLvLSIokRwFDv+IboZvHaZDwBwUk1NB63Aj3N2fXWiRoV0Kpfvtsoc9
lBrQqRhWfKCRzwwRkgMSa92Ws1dBQu9SHpfpHhxOq3wP62liyfEW3B5qvhLsLhJhe84GpW+ZHKJf
tIRBdie5MkBLqiIXKXprmCapd/9nu51M8JNjnavqRVZXb14BruhEvTqqw+y5lglnxKDcs9Twv/Uh
kPzTl5LANC7TCRtEZM/kxDmlnYz9e7UaCKsUdr35ekzWoYTAYAb7si9N/E2CoHmW2n6JyYMaNmLZ
3jeYBJtF9+sN4wPw9eNt+nTLQcfWaqio5gHbKDJgOXk/WT6qrH/GHBpUJlWxT/QxS6TRrH++gDZ8
GUl+siVgYJfUtNu/sySHy7qBms0n2cXzXL3j4wG4CRxrwrB0cPSIzO38651p0NboqGiGjs5UWNDV
5jyFom1tCld9I81CKZTxopaJWCmffkwhs+WGaFUhUxTmZWombXI84qsQERxgpp1nH2QQARl22WTb
2Saw0lFNFmnbNIEYg94nz5xzDBdmHq93SCGeI1lKWv9ZZa0ORKYOWu7hmOv2/EztoeLcE8c8TGgv
35BLTcPWZFfcnh+o0cIRaebhnNv3H8iD9myAMrOAY/LlCGuj2Es/Eirt4i++qRA3v3cOtnG97i62
IrNMrZqvDte0FccYNkx35ihgVZKAR8JcSOzRRLesJqrF/0So+gVtnE/nI0kHVD1qU7c6l0LKcF44
U+VvaeNJbJxJZ5NbRIxqRFpwVw636UFnSMkXOxpxYtr8pUAaQfTuwi9rNFovBoRZPPFeH2DUwPFq
gz0r2j3WMbniXqlvDtoyCv9crsslCrD1Tju3EZ2JswHZp/KYeUTTBx4yxvY+mjI3/sDi5QshiwaO
SjW+4ZGNzfVzI1pz42qFIHjONfEWXSqRCZlSAhn/Kw2yy/qGmqMsDkakNpWMiKquu2eOxv+iEFEJ
XDG2ReD3WRs2VV687xxeFJSGySspJgzjJcVPZUe5VtDlrJKn2YEbuyKUfs8w0s/29D7StubE6BVL
q5Kb+tUqqTPNc1byt6YJ5/+B01CXof3xJqGyPjjNYvr7gh7iIFz9LLqYSWEAmDZd+Nx0OQ5d+WU4
jSdt2Ac1aGR7EU+UhMhYG8u22b6HSD1GLQmHrPenQOfcgxRMQ1rnTYYdDAqT2B3c1zgCFONKdu9m
zMD4qXD8Ndx7G4mqcjsTDEIDs3ylhuykg1yYC3wBm7g4qRvTbhzAmd7XcRtGxP7XizshhPgrSTSF
7bcTQSd6lApuOCVc/9GqUuz9FjmWuhboYZSZhYX3a4pWQmBMIMmt14Tx/+uB4vooE3A+y9fJInNI
7L9Kn5RkuniVduLG047KMZKPEwgZizFxIke4c91CzCRad60XTy/N/EgSzxj/XhqTsyM4GXVZ1+n7
gvDLx0HzFPplfPyTHnJ7xmp62qexyF6EyEVSUMtAga2S2U7MnLCqWJHCNj8pkGsdyyNWDk+Ly/FJ
2wT5ByWgahpuVNuwhG1pepq3QObOECnMTkRYGtjgJwEjpfytL7rvadpUYsGjGRy3P2BUzFhIeJ6R
vsILbSKTtYAXOjWW1o4JniCF5iaVDM/aIsfnPXQZZPxyAQixbuybL9NEC1nLfIHx+gAW0Bx13qGY
uMZ5Y4pRjArUrkm7RKhXpyLJz/V+fOzvgRzulgcFlmUxT0auSbEXvG2s8iD4VoE8TAiFk14Jg+8g
wndJSblJdF4voNRfbdxVK+g0J6IxyO43YpSX9aOQeSUevIGyoxq2KLne46jDSt8AT5+i0p692aYx
+YdUiZXdtO/xeMl1V4WqZalVMvACElpuZMBJNR/bVFhq+W5aJzoWhCTqAiREfKE0XyBbFZg/scka
xdmFZaD5B7bkHhXjLpGghJ6GXwmQJVWTVUaEJp9tuuzWo/nIJuUgIdK7yfqmkQQz2jJ1kEauvzq7
t2f8LuvMiOpOR8helzkHDna4OQA/AOqhcfo6nl309Aw6SSRYeCddWtyiiRV2tBOaG11emXNvDXT+
KEBdjrEFvVPsFm0a/z7LzY73E+W9VRspAgAbSyrIAincgiklzT5O/Q081GRrRXy46jIq/UPL1B+N
dyc2rM7dyIGeMrVFZwiX513fLV4JDdZw7Vy3v0WmTzTFbApQ5/jbtAIsi/yUB9Zi6ANxyvSoWj/Z
loHLXKec1Gi1nm52K6/9gOlL90GYAnp6jl1vBHOBHdJnqz7jF0xn7JHJW9f0DGUJbV/zAGuu7rmJ
Dz0SqWPy1q5KMbBVZ2UiE3GFGVKC2LBExFR+O3tr2iyJWS3t6gMW7FA+fS47oSZ5CSIbc73t0idS
PsoEdsBYpPySyJxssv//2/Y/FdIf6bST/lf+dbOXZGlTsyX+YIKTa2d8WnBob8t6xg+op7zt4+5P
rDfNOLI53XSrJJdraMkjamcHBdB8Ega2tFn/L6sPMFAgiZbUcmKW2cM1e+rSHJWQ0p/KXOgwUKFb
Jj4+phbde17DiOQekvGFo34vnTrKx/GDZ/4OHH03/u8lvAj/x6nWtZ6jrl8aXAdbU+sWaFE+s7Pl
tMZNhayJDmWcwJMcOSubYwzhFUgrMJqrZIgDOfggP9fQiVttLSL2fL4FGm79gmZss5f0g01fHp5B
vxAAc5i7TCjv8STIduV3k7LosFG6gXlSDw12n08d9sOJzSbF6zPi5Qs1CM1S/QHx5bZM8gRC/gFT
jcV2WQzJK/TP9Z8/JpijwSoFioLyBZG8oKh47IhpJC2yCohCKA2YBtHC5Flf+VcFsGDkYtUSzvhn
l3k+H8HuIwFaOHHidjficf+kIIMmekU9W4mEpEKPKbV7HmPTM5Pm0SRX7y6oy9XZvAg2m/1lKNon
RTKBo++nWzPitEjbO2S/B6SQtQjPbbihVO82fFObeY8iQJ+4uM6RinKyeJwZElke/w+5oKunW6h4
7WLQAQJG0J7PjZ7pnCHsawKuh/k7dAJXOEJwJ9WI6vrqOCgDhdSTgGsMlElqZ3PDoVBKr1fPPDTX
nqr8ozmMcjTPtvK8wVhrKJ+XI5pSkTbfeDwveBZOto6eqTGYSWI4cllH+PwmD9LXSzdw8SbzouFF
Ybks6Gq8S/mR/q0i2fAQ39GcjA2Ocqyzk8OQjcw9NECYlwIeJTzFsTpgHJfs0iph5SEqjSb6Jn+t
898BRu4NZx1I8E0dpOvHwbdjF0nmOCaA5si6CgQ/RPrL+VqnAHTzoHqwQpFCgdNL2s4OuGluX8LK
5D/xSy/7uG1p44r57OkSDeyXr7btGMJOvy96IRsxdZWtjXLU5Hs9MjKXZgTE+sGTVCe4d+CTqGuD
mc2bdQWVarU4COVGGIV7gB1VwJyHKSKjci2LcjgAHo1RsIu1ZXCXbrPpzr/BokFFiZI19CcZwqCm
1oNqlIigKsbbCMeqvqyBV3q9COFUX/ZdHDmmQyO3+rXOa3iw0EWN2E2dU860ery6W4o93kCZgYFx
xRh4PXXhYTZLrmjxT/Y4GNkqQXy0KO1Ee7NEwrj4L2ovhUisCrHRTR/rAFPEABP+T76+6RMyv6WM
FLVKE5HgCgdbs9WDPbgaqWRJwZcvB4vmoqY0Arf6WGMS9Z6MKR34+D6hMuJSammZsGGL0y6bbnTj
hFnwZj73ZtqGfAyeRgDn888YYYYlb9jTBKy1U7/Dgs4GsNeGqSR9aKuIFh2B/AQc8mBcLSNqtEQX
G4tV3LzCtzqhHdk42m53VelH9x0nJpLr0M8ylqualJmjE+lmteziNrQCGGeEp7lrkoLQXCKn+DLl
hG4Cz0gJieJCx9I40Zn2dtgGE1FXzhPB0Da4kA51nGBR2l0eejJlM34j2TuIRhj6xvpJMBa5Bsg1
Sdjm7pcmEZgExkNkxQOWx7UfIY412Edn6RcE7/6Wf3vIC3ts25jstay7I5taLUEESTKB0oc0cS83
1QD18sQD851fD2V6uo0restCUxAYm2L0n1JL2OkM2iF6rxWcZtypycjDPr/zu92/8CobPmHk1wQB
t57xYLXzdsah9+y9lYbaBQt+lO0dBVZarpn1VYddr9G79fTJOMQktU796KipMbzjqZ8Zd1zwDskh
M3BLQWQTjP8ybA2ZACvX2N/Bze+n106RMgIt/mswHkZxbSzmga6c5tJcdC327esuDUmU0OLDLmcw
u4+1V8lerSB73eRhfYqK08Ljf3oe7ufhJBj8FLGaZ+ohcnhrcbqQsxp1UzsOcuY9k8eiVWrxLsGk
xsg1fkiTIlSxfZzsy/yu8cB2huCdnwp0FzgMOsWH+RnMlCCqN8e9rS08C98py1vcBsE7+GjpJSQE
BDewUVkeZ0mqDQM2JSRS2FiHRMNg42VMxooMQPyE/qomXgna2IzyHjrV8AEyi2AmNEkvH0DciUVz
4oKuZALLvpAzOm/GDSp3AYQoroRnaH82GeEe1qujyOmFTBAySiP/aZM7DEMJSc1uacO1bzTpJfcV
7cRrJoaSucKqGeHe1C2brh4/a4/fjM2zAgMbHGeOVJZW8CqlncUwae7JUTJVv5aihqQSjsH2tMGB
wVfQYySam6pIj9rZpr4H509giYMHUyvaTcd9qRjXPMINSflWKy61qMrvzMyYX7YBh90ZrKvzYgd5
XvlgvAENcw6DARQr+gwdR2F+qLaELsddEXLMEIqm+jCVKkPk1JJNuD50tFSMCg3ZYkFOrj3OU7Ru
s8p3++LHP34eYiURkIbIZA/xmNzE/R4Ijo2hRi8eBFr4UcipK2GHPFcSY9hSVM/cUn+EAho47Auw
RmfaOVr9FpDjsgLHJfUlnA5nm2laSUxWcC/ELKbhk9+JJWdgUB6f6dnijpb4Ok8otDjrHVXjZ7SC
9OPDpdbb+SaAljC9ETJs2EjJIXqfVcxgI0TTq4F3DzppeOaLtFbtBc3ZHDjdNHHWm2hyXCEW3t1P
TKRBHLTlZuHNIEGeiepZKBIylCXRNWhF9HWxrmbizlZLQl7dqDQamVwBg+SBO4cwI8s9I8TPLZyr
108g6oIAbj87JbPleIOTVcpG1nqP5Ol3OXepm6GzUgkPEl475lBUJlhwuiyRv6/SEM50nLLKiE7y
kh3OK4hAvbd7yq9TKLEw/c7OYdCEDK0FaaKS5OTbXGJ7WjdhN4r8EPmJ2xp+G7x5CzZAUm18T0Xq
c1fFN9KHmOgwgPuu4YnmzZ3k0KJZN7r4rWswOA8aln1F3QdtX0sGAuAjgnuIjOeWPMd4xpuBEcDC
NqWFlMozerTxVBDzcKbCDmEIwn8P5/SFIaf7FHVH6u945zTwowR2/hsFEerRseQ1RRVC4nbaKsvc
q3bnlkXdyFpGOrIxoih+PoYapezwk139+IUBiUuQDUmrv9YbpzZFt9a+IdJCjoekmrZyxiYP3tRZ
YroOBBzrBFXQyIZKxYNIReuR61JZ+RqtRTeg77pajjGklKq5LHHcmeRvZwtBxqShicViReJo8FNu
bWWh9lALar4HUi1IBnb/J7V83eJB8AMJYvpOi/Egx5e5zWG4KxN6jFKLLE3o4WKxcWzI6ywYs4nX
qKsxnpvP/wvuIUPBtq8RBSI1UrSmgIqUoTOYZFXfj8CNIBOcbnzjLz2Qia4Vh3GNfC9QERjSnACC
ysp2UW1PmIdR8lI6HNAJ92vQoFHR0YBwAsq/nqvzzsEgLDwr1gc6sNykJGXoLx/JO3QwutpvOzOD
dR4zAGRs0Se8euwbzUi5rPUtMXRd48zmU/FZxFrM4HkdFVTu+YNCOB5191m44KsWBFdqY45RXcSz
yL69bbwnnSblXYu43tEZFRPmUFk7e/2aEniOcaZ3Tz51W+GOk4/36tjwqY4wWN5TEDK0w+bLptGs
kUokdxWfX3romuZeDIViOLWFRbMWzVH4qZNgJfWKHswH7nm2KEcqQnUC0GF6Hc+L9ri+DAO3XPPa
4Hs7zeA6aR3R+3wplmNwefMy9OinSjKzBuSM+R4WnHFgiRBVZkUXEaEOhEGm0pYGR0gHyFmd5KcI
rqYCy6ih3Mrv2phb+fix4gwTC50M9EPfR6Sn0cxvywpro70v859ANjUgrHPavUEFmXN7HLMXNLTX
OmWx0prhtYWMlXthFuFws8MZNkzSgqtHrDQmwolggn8KOBWHtk7wTz7s4gaSdRtJOmrYV6poRNcg
Dxg0fZvuXWcALHUAmO8cbnPiyJlaJSPqqmPnAcm9V/orMtrkSXG+qf3uXQPlr6BZfUbDn+2ovpaJ
S0bX3kNZgmZWPx4K4w8R0oH4fvXmj/v5gAB0fXMr8h36cUe5hhy+PMgzEQKlZFDjshRbg525tUGW
yTOoHoNB/WUyQcD/Cc/bv0vcP+g9zDBWkcFlwgMK5wqOctL6CUuBIpqlyj6/5QYJS8NHfJ8ChRk7
vsdIX/kPEXdBoOSS4KOhiU7fvfPDjFaDuaJKUQgZ/ybgopVpRb0gRWNWWSJMF5wGbNE+/eN6R0Tw
olKYEYEbBQrV6rvBHnKCPqrAbLWSdw5p3FLPEGteJ/xuphHWqjMLS3zSFngClfU6MZWbY8dAvMhx
NljxZhh44mj7VkLWir+jsUqFFcSQMNeUpK/ZoG8wYYEFddNNvmhjxQqi0Mi7LeZjAJbkWEhUEEfH
m501WDKzppmeQB8wgzOvmlCwC7Ifn5HO9IKikHfZ/ZjZdr0oK6fY9K3M4iawnm0jIy0qqKFhJwgC
6QgHeQYpW0kiJKEqGt0oUGM0wHF60IUNs2W2tGi5EDBsn4WZC9SBwbz2cfkqm7Zc1IuDzQl5eQ/z
8i+OFmxwGvRsBR3JC+xE7/s7Zr2Nvm7wabCBI6a3wJdpPTaykgRUUmIkq9UaQSKjcETkgFtlOJxo
LB3XEqVU+l/6cD7K9itmzmWh25Iqi3ls2fMbYGtZEWY6SpiLp2pp3WtTv+bu5Mcnm9tz98Q0JQB9
vQFsEZWZr56ZNHkEDnHejHY9zRL+lhSRKcjx1lFKl1ToOsttupLiiN8LjwGOwdNgzVV8jmVZ0YAX
LjIipw4IdzhI3oEM8l2JtSlnnkz55j0nRcMUzHZbLtfQamMtR1U+3PFRQ3MCDmSRkZPiuHpbVns8
1hcim6UgMbJnFN105EQknCmdhQIO+AsSxc/w3GkAT0Pvku9pN50lJOLX9JAUaMdqbwvV4sWlVOMe
EZLSK9oXhzDzs3aVQX96OCj1k5k41WsXLXrE1uaRdJI9sEaNLsRj34sLk42IHq6kmhz0gmPrT63P
z2G4kRh9Pg6EPFC/m0sOU132cPvZVg/oP6k+ARp4Cc24eibBBawiOHhkWs65sGcfwq9OsvkwPcCC
XCWObshai7TGBKLdrVUfR+DN902LFCN7GLOuqyztHKN4238uc44FATGVxR6xZWP7yPnd1LbMfshi
sPnsKzYZdgHEWYv+TRAF1uH0YpsKb15ijtnpJfs4G/OjLjqB1SV3srigQTAf5NwsvaSXLOsuqgEF
vgPfEwB4SAuKqmhP/SvBvQWZ6CVMO/Hd7J14D8AX5f5YX/6QZVp0bi5UoOqPiYKOnBKhzKzX2xAK
WMbX8DRnFSe1jluBHG8Y/oVX/4VKunfkY7HFzPkiDQ/5/luXWWNEGV4VxHytjrRNIbFPNdU/MOOe
Ay2Szuvxve5DdBFKzky9SrTeGEVGeFa0Ns3pA1J2MO6tT58F4QQF+dwMDWpk46TgFcev9ENXpXTq
+CKgq/YGsgJrVJjP5skDtRS09lc9W3RWGXDAkDL3M1wHY/Rb7hsiQg1lFEIlYa5X7Y85XV/NXF+Z
f/prCbRO3Y818AC3R0S4NuxXxVHoaJvtWeEwSy7YVl1zn/nT9XwUdlMuSpmWH28+k+4fy/OfxF8j
9z4gKSkReqUiStbe5Ek5fUH4+rv+0KsFb2uPp8nui1MmAk9RCBJwAMcv6oeoqoCzG3Ft2rdemSxT
L06OToQyDrcmKwngemLfEMz1qLxUQBPnIq131p2oHdfTeu/8WlUQAjSMRW0HaQ+ft4L5DmI4rgJq
pELXgrUHPiubHOlcppTitPYNDwjAf6ZdrxM2cvkRHat3L5cCMesjlafjNGkS1f+wovMvzwxVou5Z
FzFZlRd2jtLH//qe+wwfHmQ1cf3r1gCINN3HSvpmCWn/zwJ6LZIULIWlBzdep1/0qQ/Pjt3fYGTy
mItGBhIXDTqZMaZeEAQd5Hnd3tkoWwM4BhtX38oB3+B5fMgOwl52SDX7pDBm80Ds/gF2jSkuXiaY
MNj83PXRQYFQVv14oWJgGlWrz4ehh0/0P7x6M5z/Rp9z/tSBB+0aVPgOq9aYCw70hPzhLtnWg9rO
GtpSBJl6uWnizi/rD9NqBvQGFiNlPqA2GbIkhkJgw0TZirAoieMAkssY08pUjyPp3o/YmorUd4KN
3FT2auVat+6fiSfmsRxLv9NQJ8aS8kxkjK3E3ZAS8EYs5xqNNp4rYtOOweLqTlCdCWfp2rHYslg/
tgpXzwMrpeT81wfIzGcFNnzpqO4+qiYNV2FtkmoP25o9CwerzahHILVnOwIGGey5mpmNtqKFJxPd
yrbmKE/NEEIEG3HkyR1s7ceWD/Zd8tgopTmuG42mevG42FnUaSHaOW8QI0Y2cneICUDOGxVkLJrg
PIRFjYao6Tm86WiY3+9rErxxUJnvdqS3o3U0/+uZUDjzcLeIy9dDriTi7QSsEHn7q/K1k0bJ0O0X
5RYzYK9179s2XhRFr5Gus21zd5ZrzgBxb02+hfiwXi7VtlkF7Fmw1N0jEEOEadfAQbhKsEaOoEEm
enRNQFBp6xIHLStazOzNFdMxFS8RIUOWn2TyLvyH5ke2m7iujQLakY36x5xsSdMfhEycj7miv3SH
eNpOxjMXRRrs0picrAplZR9ZOUKSOaqj9Typo3HaFMRjo9vLIAbxDSmLnTryiLOTjfh0WzWXVPKy
OZzDNz+4BHupUtTJ2jFPweGnZaFZ83160CZZqeI+TRRwUu4K/GIPDXF3FJSgNfiDZNQFc2ysGnH9
4gTq1eOe0QyLseCYChXxZZMM/Z9FpZ27jdTJFeAYVa708Ijb5UZIxS5tACfuJCI5OCfI+TKHby25
nTSQmW3ZEt5wsUhqQEMi8UuZWTgFewT4T8Ff+HJkgkdQWouRpWt1+a3WBD5W/aMUZjdbe7+tyI46
8akBkGaGZP+TgCYDUUYHYYqv16AoMfjLlxjvhDD8fTnCIRKRmNDpB58gy7DbjprqO9zqC0Iy4dWJ
hjnGI8uuR4mH3LIFNKlKXBZz723C+NtPc+jhGzCZHzcHC/2mYN76fyPvnfY947Rcmtxta+wxjBox
EWi8k1V1EpxJ3daKZQeFNWDJKYzM2NS4uNTlLtLjVQyL+IDqEWI23D5xkabhCUrWctVwUqh4U3tO
2qfGWyQgfhnENIp+7EJDUeljkEYAuKCZAov0xUOstk06hnAKFLLc9EVZiOlkxyNOdlWPsjuOvjdM
LBafS6eVhxpwooiUzCQOSeyV46peWyT6AFQWJi9eH92FY7fQj7j+Gf+CrM1cDWlmDyVOnn9e0gE3
CfLkH7tJyMxQ1uqg4q44F414Bxb5tElldLL1ujCGqw5oZ8vvZirX7DqmeFFjGaAn9zzrC/Ue2Iaj
ptXsX1zVbI1s9tF7L7/Z8oExDNBmEjIXbKBKTm35/1KOuHlyt7gmnKaqZ2xpcczJy4hwOZfYgqt+
eVA5xuR2yN5T4inXIDX5jeMRk5HcH0rI0U/30WGbpnfwLBmbxS1JMDz4ZQM61FpKTDq6pDhLBNC/
SEtdZXsQ6B0+4+AiW85csbgTZAVI2/YkZ+aYNlzUumHtsxWfumIpYLFGaR2a1voUDPzbtcW4lQQx
ALJ89/hJEOKprhLqqilTfR+Ie5PPFPnte2fkOVgu8ClWMP3Mcl9LPkhj/r8n/XNjZBVJgaJ10UIY
OxgJwv0Akx7322vgDGsfN8AaSAIHPCogWUOE3voYbb2pYl/dDp5HVv2PBvT+u2M3OZ+6z21cCuqL
ttFLMP80gNQuvCjoWC+EFOG9i4TYtR6a19QDPEpq+ScdpLwdXzwpDz7wEdsSXrKH3Tp4Sg8mGiSS
L4v3zH6UYh3Jxx2fyygX+Gw0fNJmaX+sutvEMROvR/k8siNeVB2ypQazHDAYeAX9ivsgWnd1/nvS
2oA43NrWyE6m75aBRdj5yVFfB0bFeF6uVr/exMyO6ZyGv58V3EA5zOUCOPHkQH9uup6ImEV/BYD+
k+ogDe7ieUzX491Jfjja0pW1bKxW63TtiAuUT0oEzloBtVsPa7IniRkq1xz7/wF03YCGKb2K9HXR
Mb0GdRIsKgkjtPCF4/4IFtWVmICHLiOpLZ43qUv31SapWVOUsHvANt09DtULd5z0kaGhY2mdvxLU
4jKhpvhtl01JBkseV5wWsru2Fu6NHz8x7eTm37T1oOcNaceBhDMoZH+Js1WpLbS9kMqaQAnnQzeV
l9MEJxylUQDPBh7mLJtYCIJdudq3OZBg6oq5NWcenvyFw1t1EGJKB/Tipujjd+Wqx9PivmJ5sDN/
pCS06NgdJxspbpsZTvnnFbKjRWZl0I3nvMKY3S/HJvcFYX0lNPvmA5ps8G490MSxAe53gzvnqYgE
PVKqqWA0/ZHfVqiLkT77CsT3DHsJXxLKWeZDY+oaIg72kQUDbKYTrrPtmFXDbHJFbMJ+F7D9KPe4
JbkIn0ud9BTqcJqZ/w6otB7aE9uK3YOQKZdM5xoPJVEJSos0ACTaWZ0M4bDtFOq8kgeyd0OsvWGr
ao40cQwOJttalok3q403YhJXXHe1SyVkWyO76lRQy0HildMmriNoVET3rjULaY7HCU1vbMDswWi3
8J8HY0TUbLDPrBreugUcCufiubwJYoWex8/CNsDfLsCLrcQC6DVLYOjOHbAl7P2sykgacAMfQHFT
3xBo90Czd7UQSEoR03eLmbd7IDE9YGkd7pwPX/uU9ErIEPe2simugTB5GaJJHjA1y9ETwP4RdqyY
Jp96s0bZrMkAx1rc2VwdFeM8Em5WEpW08YodoMc+t0BaTIhEtesjitP06t5HtRlPchtO3iLew9hn
S3TFtxLBEjDY0DT4/OhokBcpYlbqjiJ0QuoX8OKAyztvhRipJjefOhAYYDUT6Vw+uSK04KgV6sfK
4pgbi9hlXWiK70HMf5s1VcyEWiQzESSVaKmw8etl/+l/wnLAmOkfUjQhfVe7joQKRnVCNLvwm0wX
awu5hlgcFv1qgjlB8qd6gwfYAOjQ9AvfR0GhCzdwQENDSpaM9c7M2LOzSF1br/YW50C7lv23Cw2W
KQqS2W5QHt0R6HkR5ekVsX39WFySthzhYZu70Ap89fvDE3Cxza1FzBraz6IkIi9CgElMGjhXyfFg
r8x9abX5Ow1UJY1lPG5/JJ+0dDnBg6g0irwi2KXF2zIkFxVWVqZwmMSmDY6K/mKJjKh+jTVHmPGa
GG+nbFYFrPEX23Euyom4nm7GI2G/v4ekdzS6XUlYs91cTe0AtFCNT+AIxdUzWAKWomxv802reY7q
ZBGd55jc/N/vutO6NCosH07LXDwSSJIi52G0GRNzIf+l55/HwwUiC4RUeREI9aB4F+QebXOBB5Zr
vqqfRhmE3Jn79337L1FOBWGwNYO24YHmsqnIXcqidW3gdyQAKqQcnN93kfDXpSkPTLLftXdatnP5
K2p82j3j9n0RyyLB24PmsAlFI/5izjZYLsfYUBze/JM3sdnYak9e7ethNFkmcbe0Uup8e/w25qWC
yX/Wkm/zNIb9pbY3RGxvpZWkisjygoUFvsr/Fdjbjn8hYzBPNf4VQH6rG4Th4S5dERWRTkPAqouq
FseoFxkJv2rPPPpvbUJxDJ6z2aIHjlLHqch8vzPQkunp+dNjrj2KK1LJUdEVL7tjy0aJK7tU3cs5
TSQ0b0o8HFlpgxDW88VFfNj3GGSLlqvkzAhTh2HWGAOCoYLeZPRIz2+z3kJgortViehpNFmVF3NV
aPaJvnYTon+MfgUGROcOKPG8sRCWLcAmA4A8qjFYz0nmaiKHj0lQiDcQxo30r4/iJNnwbsW1F+/r
BU8IrZrdVS8lmon0TM4HUX02X4BdXEOTAOlayEbUR/IEUv2MZjEL2JeQS7N+lnSHWNPVjscNbhit
DdaumK7D7ab1bh/Xz7MNfi5c79Txl5QbSbmfgV7rKAvQnR07uIAlQcIUp6wu+ULwQ64mwrRZnqa8
1mNV2tgQ1pMfSrblKwgLVXwYbGoCZJJ0UHkjgXjqWr4yPuMqaFSMbUAU9tQhtu/pOBffJyRFq6UV
1+M1oTqd6/Za3HrOO/RYgiJwi+ohRw4biEsRAjYhcyVQeoVDJ4MhI6z5JEAf7dOBE67aIm4JRYbN
EMgt9vPkfdfUoEl369lXuvQS6JuQFEBtzS1svKHCk9fAvn1BfCqS7jekhL+k8hWZOFpsXYe3ZZr2
lecN3nqm2jH9XfiU333gYT1HrhUTWsOK4+tn50hbUqSV/rLtP07/hABX8ngI+6JTqNNSPl3cDZ6R
uNqsFlq5TsPy2pjiFcdcIRHnIyg/eQbQtwNZKm8HlYEpJcdMz+GlvPm3thpyjIcEE8UOFSQYe48v
4MBYEwqdsNQD/fC5ln36ytQnA+xJB3jZDMnI3B9Ymcr1QRVlqGI55LGCiBlIJPxrrw2tunn9iI7B
GPZ7x7+8UcnyRnvly+R+lqoPCHM6cFeL1uIF9ANLD4k5euJ9vo1dtPtYYbXP6uHLCubmIScgb5Iy
uCWFMU37IvVHmhhp3rC95ySjkDj9RUIj8AWuI0sA8/zaKAdaj5UV4qVqgrpmA7NmsS+tG9JscgvY
tbleY5cdlYtRPhVW0X13y2XzExkcNvDZyrCELcYvISP/Kz99CWvwCYsiVNhp9w5RJx8oRCp1dZ2U
SrUou0O2yi1+/bGNiXwO67PSL5S1GgnArj6xgelAheRce16MRW2eL+7ka2ZjfqeQgehTCkawl1nj
C0lHWanaqo3JNPlwBtr7daepZYm6Vh8niJJj/bmH0LR8glOEDdDWMKWxvgC25arGxJW3ieKqKugY
SQ5iQ7A1C4eKVxPFp0Wm5xUK5W2Cui8n4kUMrv4d9l///C9VnQYG33A+iDCQSp6RRJ1eydLo/Duo
v6UgBKrAv8GVCUjlrL3j/TaiKVODazJtmXmHdUO8UPosvQ6Fzl8A/K1zyE2zXg9SztuldUEOT9Uf
8Mwnd3U2gGHxNlYQRGOiaQu22hHxXlmlEswT8YVLGcwxcXgLa4lbyX9EjK2XqVf30XPhq4gVJUzm
hsdREGQplLWRA1Jat7zIiCtC49rkPUebP6dfob31VrNFilpht63RYPSKBnW64Udg7BLD6fSSVilH
6FapKDAW9AVUbQx+bGUjGYSOlf7OCsRKONAR0Ktu3svF1xfBo6rftE1MzQby7pnYQShULMnG0wBe
NHn5JuLXHiVCjvtw/snki0jha89Ga12qag/5BNC64uaf6+Bm3TXnQulMf/s6hFQnfp8sOAo2PmfA
jXh7roSS+wPa80tSsSBnuJwXs3PJxpOCzt07hWtGPDS8FiJawGn7UovJ+aUVIw0KDj+gUARNdk64
WON/sQ81yTZ97xETfPJ2aEmN086lnJFM3AkqGv9uX5kYBjkVvU0GSUDVvsqfGtxFtQBijWgw/GP7
CMf6kMjZjcKBP/WhcgiMJAp1WJsaoZDG6Kpnqa2e9o4v62ksce9iuY9x046+HG2nGsHnmRc0zzVz
tSdjjdA2fahUqvhCKKQchvALpMucbq/m/fpk8N9YiGL9syGEywNyPmKpqbE6oZCmjT2Ig4HpudRn
oxv9ZzakwEiVI0hhrPcms6daMbaMxch+xgbtBZ9xeeD/K5kupUgdW9AFMRabJp8bdzhY0dwFlPDz
Dqoe2/wKGFwnhsN2qS/HluTQxw6lNmPULV5XU+yXjA+xZ2SMOFOKAHWDoqHm/0UjUivruvOY5uUm
NLnc4+U51+JLVzQ+LTsXdpdOf0a/4GARFcWh4V3Y599K+vJdzm4ljVcA3gK9HNo9s7tuTx0UPhLZ
KQgwuv14RA3FvYbLSxvHWRMisb/mOGjk6r6iPDs2H5UQUx6J/buT+oVCxy9PCnHtGHhFAbHbHzHE
WfQNIH9rE5QH+aJiWuu3xzDD1TmJrbLQFuobhpZI5zCVv2bfSKWAp0vi03eML2E3ZUTcC4CPhFHV
aHQchhSg8cmVSHNQpZTXv0qCMjfoEhkrtztWYz2QqzdEcZZoH/fMQuu47igZ/9vU/FpNFBtPMsq9
UsR2MFIyfBUydoH6rTx/Xb9ZYWSccu8dvy846is1jYSAszeJQNlK5fvukwfg9m9bGgnR5Gcmale1
TIbrgVEGuHjg4dDGhBJhgto+usY6Bj+BiyIbBNIKmgwdbj6cze2uv4NKQW5BDwyPvzSPm85xLEvY
aewR7ElJttG4xiE4nXVGJTF6XYRY/GBxqB9NRFJNd3LQbOxFRxRel1h9FmRlFzEnoHkzdXPTDqVb
4doTT/iCuBlSGd1iSDPVlDuVyBXu1pAaNHOPnUE11qdtiMg5eRk0wRVmaqpl1Yz5VHa1bHCxmx/G
qfkV2S70qv0hUp+VYWdsBqoOE8aEEItJy+pe+FvxJ0GOrSMggqkVtUOxmXX9oCV+ingp1uEmV0xG
IwXgMAGFHc9Z4SZsCHqk2PY68eyblAQK/UfVx1yKn3Zq8x0ci6vBUFl83YJJqRG2QQDK4EIIz4gu
7Z4UiAPvcSo2anY3y/PlT8y3lGFAQaTj+pwLw0Mbb4E4odeFgr+ZgWAFFmS4N1vY8khA2DW4HkJE
Kfcw41+OnzSmh8MjfTfK49RVZd98zeRiykqH+RrqiX75BrnNtgYnjF1mIaTpGTlpMV7QQDFUtDiR
o7dY2FgveZPhwQEGnNrkEitN6SEHUhNm3CXroUqgXYlZqYUmTHEcTE5I2PuOGHlD/6iTd+q33YbD
8Uq+LqXwRlDL8tvsxspCUd45RXdMotH1/zv+nZqEDC04NMzzrQTieJEy6wcSzI8omgS3UMGKFWKU
I1fGYz6vaV/jQ9o5WI8y1pZ0sYkfIrCTKBXNaafEuCynOibApX4c23y04hfqOzfh6vwNn9qaxOeH
QOQvtQRVdn/lp4H2hD+uk16rq5eyA3gSn6cmmPk2d6uM3qeMmgrppNX9QVCI37My6dDQqwqc/2Kr
D6oki1faHRSrO/MT6NBO8ZPiUy0lDC2Vz9pHyqqRM9RJ0HVr5PjesGtzW2jv0z23x0SuPpLaI2oz
gkLlRRFxdSqOpqt45V5yvL962WiRGC8AEfDo9lpC4iSqSC3WYeeR3fawo07t/rrwjB0pREJvxGQq
Hkt3Dx+V5gpi3kC7sipc4W2Zi9uin/X7ntjuGEgJBIuYdUskycGXuOb3Gp5GkxzEQrFvGQSzu6J5
DG9zIQhojmwg8wuIAqbtK6yNsKvsDg2c97ZwyQR6seROUeejRKgQELw3WpjuvEvd6rg8fJpPqRSZ
MXe0DjFiJjNQiQT59GrG5K8b1s4yTuiZtgo8SeBzdeeLPLKQqZuCy+jTj4xtBcbFXeqYdOGjagjA
tLeQslQWlXx7k+0f6lhfavhJmz6u9ba3ONiDD4I3EeFcG4AWQ1bxV5BEn4uRAHazBxvbGe57ceFQ
VWqvuck+rPXU+eLwziGu4w5d7RKalirwi9dhIkwDwacvcBe+4QYxImPS+I62RsRwEYT2++4u4Oqf
7vWEy5kOHteLpAZO893J3LWZ93ya2tAVrz8hMGDDMgErpE+uhJYq8l66nmkSYttnho8NPGZaGWho
fnoFrwkd+OTCHZkva04BjDj8t0vgLbDKid8llLHEg7JHxosJYxt9iADE+h8tfv//U1eQxiVH/0q9
yoShDLm+yeaUByCYZqyuf0oQPu6CDhC959zUwwyrjyO9eTYcpinTabOB0E4wtBM3fS9Hi76TAqdn
QoZ6FsL7TyVGoEXP+fof737cFGjb9kV4AMIx1+12UXqCKkAamS35/gHZqo+ir9uty+pTdycn0Ig7
Sj0Vidf4NRaaNy9yPxWvs5maUk8jZ+lkqfzc+h8CVANb8cIhCWwxsYBDjU6Cx/T1Mi8I5SK38TTC
mcI3H/Jo9vWohEM5iE1zx48a6uPQcAJZuZeMlivqlEt0eOztZnwC8lnn2dGjis/bmow+6Vi9thSx
IWVc92kcM61Q0blhyjQQzap+Rb7AQawJexzeaJC3lf0Y0ubxk7iftiJOYCDknPr6TBUqHGzTLg/3
zXsWXEnDnW457dmcHD2WQVV1zF2grpEMy9jzjuPSJCSUSuzYSLFVDqewrSxBzuTJ5MnKlolCL+vP
kqSwXHOgJ2+bszWzefDkj26/j7mQOHv34+DG5EieBFv+MB0dAWBBa0evfJo7xLQcf2BOWCzfYPtz
5OmoWsWgtN84dkrjTJIBFnseMq49497CEqXgYGSpRVUAxjZ0c5I+6qY4jFt/0SoxopxoCKuc36nF
Vk8pkJlB8UtKRqpoKAg3TeGKfmtX/vGdXJnkeRUE7Uxyc1+YOCtjsX3udWNvqb3spyh6GOc3eEvh
j0AHaKsf34IUyi988Znacv4pbBg1YHVi5sOmMC8Du21gIm0eVdoDafu6/dfDo38E8gvhnDXOV3By
vKH91H0Ue2+sqStHKreISeLhJa/xihUgvVs6jYZ/xO6DpBPG5QsJUZpXY5RHWcbSqJYht7VDNCJb
TTIB0NEQEnJzMMHdzDNExFI36A1yhlRLljZMl2XA+fngv5IA3pNQp2Z+4ULvgsGKO/P7hXT5118V
+UpBqK8bu/8kmci+9oHeSxmS7RtSu4sP0DF4pwsPgNltxjQp8YXUIOE69mUOR1MMl90sqBAV08QW
HBT4cLnsw1D0ntL8Ixq8O9/1WWZNW6dv5dncJQ+cXJ59i+qcxTaFI5O5qbmKYhl08HvbokUn5Uih
df2GyHyYZAh7ihSGIhe9FwSr89Iq+KPL9lGRLEGAZ6sstuOOw2mAvQTZpWGbTuzgcAwmcdOrK0mW
Lz8OTLv/hCyKi50KdO+sZXaB3YzfZrJrAg+D67a1TtUdWrS1srDbetg1TaJu3xxnsIoDLQTfNm9/
yFPJu+B9EZhCo5wTy55Hnm/sM63HFSO1YI5om+cXR/tv5xkdQNBzE5dKv6JnPkw9YOyvebTlNzLu
D+tDbs1G/VEQY/L7evt3kWxn3GRSAV/uWJq6ZL2kDshedTjmmGF+u6yM1bHoPJiRYQEYUfjO0UE4
PaypMXmEuVx2DgVdX91QL2SoO/WWnuaKgK3spFCTspz0YSM/ny8s2DviqXezLv9y4K+0Rh66v+Xm
7w9jGhMX80IX0Yr/GWNN5YeXvl9usge2xw4VQK6egReYhtJASbOtm4rYGMqxCA/gU7iwt8J4luJj
cSL+JEMrYxtwumSL5kZ5/K6fuFkrhU8zuRbdsZCoSVDDp5Lj93CocImQKE3iaZChl+KlV4CBgd/9
XZnC90Wo5G2m1waR+nasI4rn2iFwUpjLVsernQ6hRm+9BT8uvflP6qy8Dp6Duc+GjUZJdIAqW2YL
UEOBx35eErcyeFlcdyJZBpbvFHjEVE9pUeZKhxLFAyrtxZnZZYRoqKNW6a2+8o3g2rKzIaC1x3GV
d/tp65z1Np15f14q6nNZH2wqN07tag+FzbyU0Xf1tQLQqUME/rwRaw2BT0ZiEC0dubOBl+TYtIOx
rZRygABGGgSWrmmEauoe6EHOPIl3MiNU0u+4sjos0lIv3smlvbLv7T+2Z6obaDvnkuqqM97rojG6
2afN275xUn7ih11vI2P/GLfiZY12s+e/GfL3OWpai1SyGx27j4fvO/NiPUtSnhssgLf9SAL9j0xA
i5gOicn9aSxN+08po40dMzMxv2MVm/roJlewX25vIPPPn1XWeM/wkteQ+FZzjpccrV7/koTNrhnW
osQvg4QEMRIGTmdQ8xrcMK3S0EjVq/iYcNTTo87+7GVGxKHJpAvboBwOGfYgRZ5F6aLfOrcgjlgx
m1PTlGcUUuDQ2YmstcV7fhBo5kouBalfzsfQOjbQQJ1kLDkfTW1iguJAu09bd5I87aQnRph6+IiB
JUXG5NhckK1IAveJorROpETfbej+BP9ALgib6ebqkpuqmQe6d+O3dS4nqCMxp/0PBbc2Gvl0QYgr
ek6tAjb5CtIFBRMkuSMQCKicwA24IcUWNq/EXu/QWUgsVfYj2PZHSAwuyZQ7nBXfyjhErE9S9/Bb
bIXJhSgFRZW0kOdAAJSdzk+XFD737Pj/8D3o2Bvxp83kZBtUmKudRSUucsM7Of/urhXJLo1EGCvN
5X+adVp3Z6OVKFpbTjUMa3q/qUMrok8SoiIbKHPsgb0vm9Qji0rBrhEUpKHio59mckuwFeQE9nqM
q/s1ODltnrq/9+xHipWvL2c6CbiO4wrKIltIUWKmuwPP/OtIg3i+JB6QZy1Rz+JmTklNjO3IzHh1
TKUfl+9pv/CmxHU8FiwVJgQc9onIsKzpnVoiOMjGGxzP1t/f/pVu8gmTmTyfgysajT7kTAXKohwo
glxWTakCJ2o2DRZeLm1whmAQDvbpetos7p0FyZzknw0NSyrlxvAyPTvXHHMruT4qN7RM5Q1pqyq8
iNlQJFqwTa/g53a+v7PBccsZGQ+9xdFqbtKFfQlmnvLVeTwoTcKW8JN167wVIUTAptX+b/xK6QyJ
r005Hi3yMBPhdyi5jr7z3uBwgEek+GUvxJDkboyBJiX5NAVxbIhsiQWo8BPyMjiNffN4zRFFQ/Rw
zg9Z8O59YyD/U8/IuCQDCNpeegaoDJDCFZNw6W04GyZK4sKfiSWN1jcs7s0aOSCbRAuJZC7UDVli
I48H8+MllF2a8TJFlzbVGEwKamIBAfs6Pl1IIEeqrUhnX+rTL2aqjXKC9FHnE0kisutjfVT5k/6a
H6Z1wjkRvfZ7NJfqQAwluDZgJtLSVYXguUdpYwSoMxTMyGcYrhBikt32GWUlxfDBtADJr7pq/DJ0
eKA8mdRnR8PircBKWEaX1RitB5hEDPEmoM8KCasX0KQGpR/D9vTTryhI3gah1DRT2+XM6YdtsrAp
rmQW5IaYSKLvoqFeHKnMJTh6WgRqtyGI4fNbqOVZNbNLh2SD/5WRZicGFZpnUfY90IVtxgGy1bAN
mJ7+UrVtimyuHEdsR8SIeuIqmbw4jAbm7FIJrww+oKmhwcmAxTVyWOYYDOucwxtbzwTUA+37eYfn
CnBavb+3UoOp1+r5/zkuAmerBh9NlY5C6AQ92CYcWPcu6eH65zTA5SC/ExcqFM20Eyj+JcBhFLBg
hCPUx1O/sp05yhzIbEF86VOQsNWdVWj+erSkrA5GbteUz/QBu6X9bReeGcBM6NpWgHbyP1f/su85
j5L2yu3rWru5PlLNUPI02oxmZP59zps4lee8U8+6r3tpRKgFcIM1DVbYs6N22LfNNqCqMTfQud0f
hRscl5yoImzx1qLz/xS1o3leeqFwIR+bTbhIcvZC67JfekHPSCp4Bed4UtFs0PMLVEZi3IkNzHGd
Wr9VmZPof6l99+5gwfgUvKIHr5Je5kihHNzpu2/lsDFfgl8YMorP2W0jp9YvuLT75Kbln10pPb2p
7uvncrCikuCGU9KyzEdriJwt4NvJ3RYo313ZC9cKYtMsdzZlsgunGxUDwBdV0qrQi92xKAquJRzU
LM4HGLySVml9OOj17i3MHt75rk1EIoUjrZh+wL9Vw2iP1sjpvUc30tsDJ10feU+RNWQ1QsrMFDDy
0oFnpq3d3Mbd9pt5CumRMTYJNHQe493jdkm3o4RkdXZRsIXwdUvV770sYtwy879qayQ04MRTHDrl
UnvrquW+X7Jtjb5I1QaZ5vEisGRJ2l42hmMwjW9HpzaHctLcFBLAT3RUuLTtDgUruuqlhigcDEI6
e736fjUXcbzvE2L1UQtBlFgUGxpAtsWtrYf5lM9RLmimWCVUDeshMOUTDe92i05TEdLODPZSun3K
jZE8qmxgzcBOcRtgKsf4Z0LjMk7DD+w3coTDHVJSjfctm99xR0atkxZnmkFwWgZ11ONj1zYsW0zu
Y9h9MCbUMSxogTMjUeYzhVIwvY1JsSI7uY/n4lpNJP1MrMrgO9egKb10PsPF9rGeZwFog/ou1g3J
MH5LY2uUPpc3CCMzlsKMhXPsNp3syHBJqfWBHXIftvnd2A0Y+PHGW+KprdVETj6vR65xszYMxbeA
Zms6m8pNPINePj60jiK7BgEtqhqivb7KjjQxFm0EwkMGIFrMGr4IZZu25zWKeMEqTFOl1ja5B6a9
1ekNWlzJyxiapWNs6KqmVaIuAqIRHMK/XcZa5zT9QrClXjOTioXGuWrP32D/GUlQoAtKQwnUtwoK
sV1C3+Eqrb5Nug4AjSY5xjO1XaPwSOr5v/lDuGt9beAXugPwETMoLxtD5FHbAuD5utPfsp91qilj
/tRPt4srSm5JWB6SwRZ+EFq5xbhWXakJda1mSOh1ItasNfngj3dA8YGhgSx352dzYjPaOtu109tV
5xwnLes3VGqL7QAsfrSVgYGho0Vp9pypfl7F/IhyJPHrK6zgV999LtG5fq6oiVFAQ5yaNgp7s4Ix
H0GEJUqJsFo70kwFSpRI4KT+9sB+TG8hrOryD9TXGaAydjXcud4RyJcICIQ1HEUWb9RmXB8qs00p
5sRy3a9wGY+kYdSqDI1PdZhI3kVf6+XEyPoyQNFMcEa2BBtr2vWDydwD4Wpp4MKWdcxg+ykKJTSd
Q7IDWlEioRtgf0L0Bd9NghDC3egs77hTzWLwyqxxCfkNU4HnqvBB3dnLfyne2yJCD+20mhZXw4lG
bGPI2AB65RfILUv6klxtc+wIzWQhJY0a/KVOg43+OznsLZwlIHGAAibtoTlQlfHHBgBDeFApz5jL
07PQ9ocLuWcmCIEe1S2bnwunovEWiF5zypu8iJ+EOJfYhQo0V834XDETZJkXczm0tdA8Bxq+su+n
1zIRiMwG14qZ0Iys13Qq3eZomTPf8W0FrrWigHj5mV5pCkJkTIYqpweQmFuUCYhi47pVtI7rFZFC
1weaT/GxCumuvrKK916DqeLshmuX0BMjNrp8Ym7wnt4/ysX84yvJCCfQFt5jdZ8iGt1vJcsgCOQn
sDVyRW/UV0Fu1J82GuuOJvPddXsJpArsLestWKSsZjjaufz140NBjJyGcUCFzco1wcRntNbceDCk
4rZFpjhwOaR+637fY67Z+A/n/gVZNsFxe+xARYFS4+qr+UmDduX7wAB62VjT//Q1aQk4PGB0bmMX
DKx2UlFY6JlJohHBW+TSpRkVoZZCRcGSxMNYfTw9QLIn++jvvfQVkwD+QuEj+T9QGZfjsd0UFojE
wzg9fIWq97xKJIzWsB5qxn+zuvD3fZfnUTCMuEfdD+U/9hv5RyjkXWCsrf4BmeIJYbn3WCCmldg+
nc5yOaHCSqRGXBv6HrNCy9wMWxyrYjRoh6aPTK/x8aQCgMOW1J3vubwuIniiaj4LPpgXFrL6SxqE
oywyQQK8U4PZw4VXciiR4GOxVCyZUZToEWS75lGCXh9U3Qmh1UuxX5DDk5Ek22BSSiPNL4EpGARd
R6+9nuyvRKpT0z7PsP+GAwmJYd1JtBK4bNme1Hmq2aOv+QkCKocMyP3TImt7zLnPCH0BdJFT+5An
jUrzc+fM1It3Rq+HZKFFZfOSZXml/BhDW2PmPZYJMBUH3dxknuh3KXIblZqlVnE5+orFEVN2oUri
g4TPr88sKZu0Wk+IeeGi+J0zu96wDWDZQrApxbsN/InM2Qnbh9ZHDNvAZ6rd3z6K/xeyzo22ocJ1
yKl4lgDslu1QBsNXz04RXbB2E1egSVrzRq2+D5XXA06fAdJm52TB4ZEHizlt6tu7MRmAcdGCtx1M
pu0ZNCHBrmAHajExymqT2fc6BadtL0F0xUaUi3QWPPx92z8Ho7wGUQ3Mm0qMZG9XtRsRoPtBBk4t
tZ+soQ+rprC+mrfh2ceffX3cAXl78lU7KJfWY/01WngchtCF2PO/Te17jcVwjKu+0NFfeTWk8duV
RBEkknIPJdF2saJnFLPt1W/StUsrKEsjR2+QlJudZ65Npqw9zrkKeLqRA4k+EVUISjxp0d/lKXlf
cgiXLspmhzopkfUGK2nbTJ4u5Q5s7eA+iv6MW9WMtJgBAUl8z09B7ASRC1imSE178cXLw44psL1P
tSIS9p+KXL90XHww9l+UpgRa9WyBT2Jes+12nmN9udnT0klsb59OdsqcebZnqrEuYRSyQNbiuIr1
fDX0yixmhqKg2ZjkP3hhfwBCfoXidshQTKy41ME+z1chc+bUWhNkT1o3xohAILkeDY/K0eQOF2Ae
RG2bfNxj1hoH30wqYRVvaHXogmh6b2VtyvrvnTU/c+rYoD52S4ZHHSGHAAYPps9nXDWqmOZl/YKD
nchwOrW5QXRXL5i10CiwU4BOv5ENMn4f49VSwERKIC55/3YokiPwTeBNWiBoaTL199jI1AdMlrTr
iInHsVQbqTDpchGo/z2wXvbgA4G2WWKQw7nU8x4a6mDNAqXHKfrqD2pHUp8ZShMLiEr6Zm678lhC
gsfLLrWwBErmAN47agpy4kczb2pQGGo6cX2Y3NTtgYh0b971vSDA80X0d/2dMkKPqJTuax3yomAp
eVPEAZbnLrIugIz63Uk7TLHPtRu4OF5WYhA3GEcBOx4rB/afKIWWyDg2IXnDMZM/dKTb5GChYTzJ
15h1+xOMem+LAGcCzTkVMTzwJgQk2T/Of2M4alIHE0xHDqvf3Ffb+RcRFpbh+edBV4x5zIKN8zVS
h4O9SGTeYlFoZ33O7XdLHckf0D2CJ0TdZ4FsZiO4FGD3kBXOAfzQ9qLL0cBvCdUL2vi7X6aujqs+
kWYiPMtUjVojhRS5kpZo1A64EDA1JAmMUc7q6EetsNYqhb9laXKU1IcYJZ2AUA+d6u/goDmG3cvD
xtyi4JN6QCtmtCrpb0Gv/s88juwN/YCd8+lykXcYrxDDq6quAQpJ9oEXT1URNCL6sgdN/iYweXDd
Eo/alLAQIYq+ZQXVOW6Yzjrvplav0iERRdsLxa8G+MJUAyEXI7fzGszpqAXLzZCTmOCN2g1UYtui
lv9rt098QyQUHr4ivfGS8BkVwrWIKKnwp8ZE1E4kUiFcKgE/RtsOifp9XqG3iQFQn2vNCSJsPG1i
KfX1HjEg6ZOgN7DJ3A6gWIodvsFHct0w4dEFLZzIL5Q6uFmxhslQwDJAGBsVSup9esd+g8v/lZb1
LAZoU1C594FaT6bQBCkwUZ52C8Lj7oF+bc/HW5GshaH88667NeKySlPsOva5IWdRkjFpxW+K05xt
HVKLk2WsadgEWpRbBRe7P7R58T1qcnSe04/qj9DQkTqnzV/nzU9CISxEhcrosGMrrdUxEYiiaheG
6aGuHD4nN2cTslKHqBORMeDOIilL1bDZis79QL4CzLCDLZUgH2Nbt1bQAA1Ds5/l0L2hWLF5WSEH
/BL2K2Gu3+TCZMX3IPW+7m+d2lWYH+7c62faSwALOG4KwBiAN0FfjA/z2V4aSlvceyOxeVJztlB1
eFQ+bKZgGKL/vrgkeBEtIxaF419rEvi3uLTvmAKetEJOb+UHFate2MQ4CQDtVbGdyQ73O1QvnA1P
GXV6w5YPggiHxbXYDocOCjda6qgAMUoGAkNqCc1MSK2RdcELM9VYxa6j6agUuzmj/qZ0MhIukbRS
Kvcx1u/l5ZhKW1NMjj2uhlnxdWeCkCKuInpCM+99hBceK5EiXYR3mdXaTdoGfLKesPvzij/XABSE
p90vH53fooIZrkTJnb0t6AZI0rLSiQxfu+qEPOHZk46d/n93QYlcuK413n7qBDpLkupuwe3yrm7B
AbPUY5DOoMbGPm5PBIYpymlQ042ipKfAXToeJ0ef/PBnA/kQBDrvSIio5FE0maRdfoUp0NlhDhsl
oySWdyqe6vg21jzveAf/Avcd/0GeBnauKmsHISgaSyhPOJm1M9XtDRLfhY0EsR8iawm7cO02FIOZ
OiZfKeDCHfrVVxCTtTcAa8t/5REeS5kBvP5mCLYzAHWtCJWWNulTGtWUmAySivAY7la6t6VOOIyR
YezF+UYsQVpTao0FWf1WE23EuohDaToCtJEfn0U8Vr4Jun4MZuxSvYycipDr/bFa6yjLNgUp0CyC
PgdRvdtbGG9H9C86xU0oqERmXMHBCKvM09jedeb19GlAolMJfKvpsNquMLQ64XkfzVuOxdPaHhFP
TL9a6T1QEgHGX1nJHzkrOh9ikhf4UDNR0Crkkay4CMjJJAfocbqvolRTTK/L70cL7HJ68e7rGLNm
AtRzWIQ2pD7ldsZT2IdeZW2D2pkh8MGE4qwztOZSTOxWTT4zMrvdtBi762jfFmS7YL3H1GUdblIp
t3OY03vJfptC5A6UDu3hR3TaQ4x7Jqsc2Nzwd/jYrr/Ifg8uH4q8b55dqjkpeDxDz9o9DjiNUE/n
7ig0LHzXxk8eDzzDwAXhqCrXccy6ZbQcXgr0GYCC8PhejbFIXLsRvgnHNBaJGaZ2uFkVR8GcVKDI
xiMY/jjQz7xXrOdAx4acOpE+UN2iD+e3J1sx9QebxFpGxBInRXY8M7TX37ig83AUduJqjOopzUBa
xA+kiO7C0NIZ3gIIaCeHQJjB/3SygQJRxrXscvGK5KSx/JxPqe2GYDnMhNGmGQG23najMtxxvVh5
6kGPpeKfp8LyoBuYTDz7rZxdSTalcr+XyaSA0LAmlGpNPPV0CojK6DKLi2uzPFe3hEeLg6/D5558
o+t7zg6vspqt8Vt7XbG0fhtr37zrlFI3cOwbniRCTjAGDrfomTgIstikgVKoZO4WCEJrMQVq2bkp
5m/DNebfJfqMnqFQvvaI1hCpu+kq7ggHDXKfD5vrVyQX5qrszec4GAwWHMbMJ990g9Q00m7T55F2
GFYHTXu0RmH/kJOUY924j7fs542GK+QI7lqpLaI7+f0ZvSSRt6Qauy0n3TXOkpNVEELlPZJBKuJ+
ONBL6Qdqxcx6FsgQR0v3ISQqPcWr3LgMpl0TK0HG8bKIn6DJ1/aDmHE4pvKdXo7hTtNjQrsFcd6G
6+RvB0Kl/Lyq1zLlMEFgjhCQw0K2Eil72R1fwtVaalPogUBikTXYvNHnx95v3g+9L/W9qFrQyCZo
Tr3dELSssHr1+njqqXhGSpt4E5ealQliY163Q+0TZQ50c59V3Xib+7ZRm9m7GX0Wdy7DcTET8vos
o0O6t0WUcHdfrA/hvysQylUAgiWImvRlW0bF6EH4Ya3eQlBHXrvz7SMexUB83CNgL3xl+npkjryD
7u7XA0D2gra3Bk44egsecL7Vv+M6/sKIWg0sC3Hu1zJzacqDsL2nKt6rth5XkN+/fd/ThF9mJIjf
/vvOsdff6c/jCqRS7PytDux4EpXVdoy14DYJ0R2cmvLBAuMHCMXRaqY/tTlEBQG+QliW04+F+4xK
1qdR16S8iVYfIIE1015LhBwZwC0huaRhi76n4pCwM+4RgRHeVP8XkKsZzhw0cH+QZHpJ2pTNlqK4
GxYdtnFVm84ycHQ2JHLws5NAsjG/PYxqOzDQQm3K9wyeZiQ4JwmXe0PbRmUDsJWW2qSYUl1IBYEH
vxzCeHN/XDn5zJ15Uvb4lrH+I6I3gQANTYeYxaYETKej6VGi8x1jPp/a1KJnRph2lFVYf9Om2aft
vsMiSC6hBmqL1t/GuRjO5WlSpn3eX0g1wVl7x9WZZ9UPQ7e2AI6Bz70kLacIyK+m024mZ4HSN7bf
srQcnA5OkbDqb3O0CmbJa+z5ECkpn6u+7S0B2OnTTzkjgawD8y7LoSWPk12qgJpU9lrtZHqipno4
s9rWeh6ngKqF8/3JBmI/TSTuIe11ZN4A6aWZKwXLLpHgFlXfdz6bPzGA05FbsEbB/NH9XOO+nxUh
1g2g96jhPUVvYA3trOCgN6RQ5rKw0N5GxhI5nmrHY/W0+fN9svbGlPr27gMCxN2WVXv3VeBASClC
TPGDwAjC8LSHVc2xSJs0C68aAUrq50S9dXIcNC/WeQfuW1Yljfw9U/8HR8vIDXC+L3fGYJqd4HKo
ajx7sQsbuqtYbSUYG6WfNha65INhcIGO6G3TWiC3WfGe55TnKdAj0TuUCJhZqCMo7zrK8NUFNboa
QDGR17CM8/kn17gk2DH6RyvdAw/INL/RqSkAPc78C0jEQOepcTk78WHzHlqFtPZwNZOUaubbV3Fo
UjjFDMIYOvqrYVk1W2t9V11gsZN3bhjAwCjbpZw6yLVTOYvf5v4DD3/zIE8BNn4yTc1kGjoatmMp
dV/7vZRm620XCVIFE/h1/2FDYJ7HMAPpIcttU4rs5ICjSDRWAa4cernUqgBWb+SXX/egJFV80yx5
2juYw5J246x/DMuNG2ipRocB8o5aI65pdxGYzqJB97qpJEw4/gwbA5lD9U1S+5jR7e5Gbe3yysn/
7YvO2VEHKvTw4x0ij4BcYRGFeEYdO0LFb1/4bUv0Ep2kmw9lkZJZ7hujJ0cYweUO60vkWrz5VRVu
2D1hFs51KHbSmSb95qB8z3/SAkkjrpdh4GiInunRvZuWXZ78C2TdHViYgce94DFIZ46SyVz3L4Lc
z86xLMeAy+Yz/SmY7ismVgVQxrmIggnlll0yVkH9X5HJMRjta3jlreLQ0S0lbCNdUBOhWrTPbXrU
2TLLn4ls5VNuXGAeqp0heejgTboIDAodDrmQrilkazk90Pc9bLyvPUYCpU6UWwsGlBKKUMr71T1a
jrweORpckNgdDhD2mnfxaJkdEG8UPu0xYG2yzkIZ0LFWQnMyBa1pOWw66xDB1efHneyTOTYZAHSd
XJB7pgOGzedlKoNeUPDKWghSZ03iNavuCx6a574Ktq1cEL6WSnhk2EC+B3DxbYykkMdS1hS8NYu9
p2qp0vpV2JwC+ilZ1s0JLnOCWMeJ7DmQ1d2UUuWdLsQq7WaMPLMzTmSC5HG+YiA5sRQ8WqOPo6AR
p9NlmJCt6ngS8SLOMdPo8nheT+X/u7Xz6fJRQzmOmKSJtgwkCbF+zpRFZfI4INv+I+SmOKRMdHgT
Bd7hLdFkODK5TL4rVv9rFiZjXB8p+Hp54LLMA3BtJdkK7SQnnWfp1oAwLyGBMAjqNzVS9iPC7LW1
1/MqPynBZ/TsFRVD3FF4LdAQsTvWxTQEPD6ElwoaDmF7D3a55HSA8CVUz1ulRMeQcPHsOuMqglKj
O9iCcS5H9UZ207AvTc222nFi+5EpO56OW/nkWHLZ2Zg2hsn5TKk0lUxzjwWplhQ04ekDWnF85ZbK
z4gfH4oYR1wMkda4OJT7xS+owL4u7L+x/zvFyPgKY1TNh5Sl3meQul6rilTSoQK9R6pyK1t4tiKr
eYz3/z2qz13KBYdx9KCpfNIU7Rr6j11oHqrlkOWUdQRSaLjXQu+5Fh3rvB3wLsKG00VoNd3aREog
EQP4VbZR41+h/du4nhDtIzgg+1UHo28dT0IOKqe11bhKk/N57C3fmdEyFJrI5U8N+HuOQArNt0sD
xqPbDEXV8kZGJdF8suYQBLSCyJ0urE3o9rkm9jFICzAi+XzdnfIP6Ywl+WGc0qi/YDEEYJCKLkds
oYURTLf4Mf4hTr3K3qFeLYw9k+09+Zh4M40/Dw+xiLaELonz6k6P5pNrugnKuYPDFvPpqSIaV141
KWnQCzqI32jlEV8GZgk2wq64VqBIG+PBlJi8hEt6peKSz/9dLOu7mA5pclkfLoa+Z+yqweTgBH98
n7sW6ke4BYo5hHCR6o2v09bU4md4uwrxEdhvGgXC95TN3fhI47O1buJ0yzsOMClj5nnocUjKnOay
LI3PeBIQcGHlZ8dZj+yfZ2m1ceXhguBZrp6Rdr0eIpSj7y/mlDi3hxt+eEQB5lPIo1llwNBXBnWI
ZOMEpZ5ZfuXFOTqdyIxqrv5v/dpymiLPmOK0e7oN/y7cOodfxh1GXYcrjc3iwIBa7gqj+bicKDjU
jPMA6yVjHzCG1zmTOWDHb5jIy6HeO9tSoUWIfWLQLitDKe5n3Ly3RGP1nUXbiy6zgTZuKhc67Muz
q0QqIzVfPd078ypyeFe9eKK+G+2ZZ6fUNYmb83UnIIkVVPWPNxedNVJ2pZ4cT0w9hA0r85yTq4i0
A7gjO1anpveo0/cmwpOPdLV4898BHknq+xaiWV+0Po3JIPQEUPeBwKIR1OcK2OsE3dUFl3FnHmTs
h6Euv0sBDmEgA1IVJvOznyTjZtdJYyKnDlr6sqdejGZXPvuAv8Bui9ssvjVpOH9iknARYNAJUOfa
EEXfyyfPhcak/lR8GkBpSI6rscjqFx2NAN9JA6+CWMpHt29VI4zpNKFm5mV6LIXvyaVFY0d/GRBt
IE/C3RiUAuwvqZL64Hm6fxCdAXJqgcIELgR5udDAqRKn5oybAWg8zTJFz32bPbAbGwiPP+OADgBe
fTxURQCu7LFSfDAbcv/9NXmTafVOr8k4m1NsI1bOf7ocFVO2CQSnu6UbHRD0p7lPMSySMYI5PJeF
yh/BXov3IFRECSCVb0oI6ULqo7EdRjczshNXgfaLoVBEAtirhXlmYxoCFYGc0Tj+ONryL50UB8St
u/cFSTyOeJ5+Tsf73hTgFj8rvVaDthNnVhuhDpOwwnXN6pERsrwZ27T01DTxrhlIK4aGhHR1xlw7
NC5N8CTipBImMUFY/F8XJFHikHqz8gC4uznrlP9SoG4KOzR8yGL0b7pjR2My5LYnhOXPVxpKXX3u
C1kQC9zqUD1n3B4dPFqLxVy6iY9ipDhybCcZTXGB/P/uso7vos9u8CY43vLNPtCqQgc4W5Z/xhEC
7+JUYVZX3JS6N0RTCwXH3+4ItPQfs63wC/T/GBXCJK7c8ow5BKaDN1LWdy5iix+eLTkcHFtaYrYs
F53CNHwjgHGJyNgsCCKD+Q2QrS6MIlLfOUK5+WvfLN/tte01sN5reXdp/iUs1A8MOmfrPhyRu6aW
UqsXgEYEBVwINTDE/UBfz2uYIGz77HEudULrsbGz/0XOinWadyHGRa5d3sspwUS9nicbOQMSnR+S
VKZd3vDQweDDSxqjD0ZcJRndR4THjezBSHUd8O04l7fYhssN4Rlhnohi5HVxSpQdSoI/F8Ldkygu
Kpw60qvdGyCPcgGTL4JPG4MFNtWWvEzsLYR5Pq+k2I3ckpKXZWW6k+ia/AExT0YCZxirL1X3Nyf/
JVGmD/BI0/VIKp1ZFAmU/SJvCCoTvWqbhBXKPtnSXIG73vLUWSh7FBRGfaxTLgIUrUSR8701/NWu
QoCyRAKhIUwMu4Wcp9iibFAB8K2uFqNAZUUiDQ3KH3VNImwfj4V4KLIRt7Gt1Rcpwlt+4KeSfye/
zFtEBk64R7FyQRID4V30mo4kXNY0fSUaENGLUZq100hrMytffkvk/m+PFoHPZUbNdy09nxdOAJzH
yQwlMEm/OR+9oh7Q8bTjcseAyB/4ErMpGURzfO7q9GyaTSpZbIEXmRY0TLhk674LUhG69/pjb3iy
cwhMLDcTYFDRi8U6dFgBCcKfQjXGTMlFKrJPvPpqh9GGOKBpZMKyLYn+a/BoMa410SoN9y87rf+s
eT3jQqVsG2gaJG9ybXJj7unfW/wWrGQjE3Iz1FO+g6iGN46rDlIcpRuvHNJegKDAr5N3MSxs7lsu
sfs5EiqyQi9ZILlNusAe/+ldchUli9Wa/vTn4af1LT6H4bvvowcqe8TGBOLhBdpBsJ+1W5Uvgtpp
r59OZW667/rkzHV/QuJfn8FJHkQ+5bFAQ7lU/sVyaJsIgugI/jJbTAiU8s0ls1VGbcH3KOCnm4/v
VYSrEvGKBKbNXUgQRA88X2DCRE2n6xOt+NQMhgkahl6xoZUrI017tOfJTy2zaWVL5+c+0WtRxNWb
Es19W5BGzc+MPJQs2n9ZVHfj5UoQUurXmkQfrfFE50qI6SLznft1xjon9VqmgsLf68LHWWZoyZYR
o2A27rjK6snJ8l/RzLaINrsj75DKD0vJJzWABi5MmxxBqBxgyeOIRkBSxyYgRUG9CMoUh76pMQCY
VxJr4AtEllgUwlvLogSUplVFjVq/AKu0+ccp/MIbRD90VwkU9dj1W1ATmS8IuoQfI/JMRq+rJLnR
oCIQT7MVxqUdJwbnbtJEhzlo8vVKg/y6+BsdvN9kWx9mcUS4GqZ7ztw4w7chttMNgdRLm3ptehXN
IVjt94RZnvAJq2DRY1yTJlHrT/Y2TJq/c31axAy7kVdBYb3aYTzitYgIyZNPR7P/6Dar6i/0ARUN
z57wCVEdX9XTEBR0met+C3nk80ox8qHQbhuBC+tagqe16N5E1V83NYK2vJAq7+sn+waHLL0ftKFt
7NvablA402JhYyqPOVyxwYVFVI1RaXFedUXNWikUao1TqXXHhDyRgqtvg6kvvVxU3t9uoWAwk70u
Q8z6zPxtGM2XpZ21iiLeVJf0iQ78pUpCvfVWJuGraM3Sz4eguMV4Tw9DVTb13gz6zfzOpH5QiTbn
l6pwPRO8ZJS6DVOlrT/2lLCyXKyGWAEpNS8OcztQVGSUALcMRj9JrUJjDWz70YhcyiS5IwAo05mH
c+v/ncpYGKCXTv/gwoXcSnNb8EedcpipIA/nwu39xHdc4ReDISKJ/VIR5lYAb6nypNex3w0gLXQE
/p5YWRpMe22yuyIFDmBl3ecVjUe0bNEeqFrWSt7aezsAkniZ5LYtlu1UunbS7LmoqMmqajEGdgRG
M54vTt8xOZe9F8dJ5C9+3qjuNOLaAP7l21f82eOuifibbqXkuuxCBuqVPOO2ZmYDzF45zPOUH18u
lxx1TB0Tc6VNGSElPl0ElyGh1N1G1ifERI4MyJhqppMk8+L8q/9UhVoQnbPUoFSW/gEJyv38eIYZ
Fjcyi3/gjblJ0TKzWleuBoYEiRCDiZ/s+pCfjZ/Nah+x5XMwNee0W1GOIBWHxDuJWhTIzq7761D9
yDdhF7ZwMpxnb+1y9aYRgmhBcK29gSdKz2gkYIUP2DtryunKPOotFXP2fIzxP+QqaZOjuwi14zjG
7PPML1LoQt0BA88WzEybAre1kJRQzXRD99lfr8K1m8gd5L0MkriPdsGpGilQRUXMbsk7fcFxdkHJ
TgaQokUXHZmMnK99nSZBUxOgxURp9OoJ4gE8PR2lOFbQPK5J/waQcF5uh+lmTrc0+zf+OaPzjNe8
9PzWjFgqcw5k2ouoKlqvbUnNB+/53rZvR1nNc6AvSdQtL+EgxSwHEVo0m2ms3e5a3dhil2+Zbh4y
5Z0WhvABAwtjw5TKGHbBruf2as7WslsfdjB/obmOISZj9VX6uLkUw4JRHfuL7xeZf1yznCQwNKXe
5ilt5RJOLbZquIXqOTyimlIogIAAD0ZA8/lv5RQR7ssun+yZ8lDAGigLTiAqt5x9XitUQylPIIDx
/uK34DlMJmZ+svsGAuiwuXj6MW4KfMFS9NArLjuPJ551R1XUpUZBwBEVFLy5KOCLnuFjfjNz5V/8
ER6hHer2Q7gUt2KgUiKW1zkSVjhg9FTyMwgaVhYbrgChZflPLpALQ7OoMtp1Z1LsQBVX+9pI4dQ+
oWv7Lxb100CA8UNsdSIsCVkD6sGlKxOWNatzbKBxb6jfBHXNeLszz6WBA2pK8jY1860/CMcIyqy1
pa4aWozFfDQsE2pmZvTFTH/ywiSb8XYMD0bVaNRNBzjG8CGWWzXKKl700TuSGDLPMwOC0tdQm2cG
kgn38S1JGdSLOAM6JwlPrO133lqeB87tUn1eTv2OqKV2oOfsCN0cwGkjpAlA9ZY/zul3DEtLSeRE
jE6CNCnreG6EHXvu1HtHattOCxqh6FDd41ygeXlqHEH7tBygfoy8N5niP2hczWJb7t18Yqk+oBxe
ER25P9kMUtacWBhqzH7MTU5XB31dPT31in/UF/739N98D1A/ZO9aT7JG0u5uZCB7YnCUcUsg7U19
KDOx0ZVcGvCXCT1T8rEbtYx0D8UrJ/rrmS4jbxUF3j/sHASOXroz4jXgMUdG/5ZpYneBYiupN42M
5ZoLZBm4sdWUudgK/Lf8gX0f4pm+EcBPGFcHmHVXLhaeB3tXHDSOByB2X/VxQe3qJepHIrT8KqlD
C930IPY9UG237xcKvhCXZSiwC3ZBxu3oj1kbkkBjPWE8re2cdoQSJAAmsxtMfX8qTLBkT2M/1EEz
21qVPKJh2rA/DiYuaOf0MY9P5Z6Ad6n+gzBIex3p1mzA8MNyUU/M6UjcfrcNnMQzYRNmTpKxxbAu
tJ3JmVMFObGnXWeEgwdSDCWDrFavLuddpe2n3lawycTMOZ24TGseJH5n80MafI7iR7Sj+uik1xEK
3We03g51TfEp21UDixtoa8UAqEo/QwMPwKkCWCB/milteV3f84gBVZjPbyNj++8tYivOTOn7dciI
9M5iei+fcg/xlgh0h6aJnbxyhqBOWrJUvmKRWARA4gjT3oJtobqtWb5eK8HCFzGR/am+c20mo+kL
PgU4ikwr+ahKzlOwaT9bGL+4IB+ReJdQdfpYyAmW2qSDfmFhRPR/m2Aw2VqNb0+pW6mcoCKgF70m
ancN2lhpeKfDZP42DtbcCsJ5keY60tIq5VxzZVGfYkgbJNBRbQeKeR7ViTbq79n4t8oLRsE7G//b
KJwhCj7tDOjjExe9vnO29Qy9vimB677adTegqA0wa6GqtRABD+owyP5QrM6GrjlwTHLWdSSrp0hi
BvLDVJQ+Sd6PkIj1xYeB7VZSUoRM2hpQllOD7W/q1LtmYlwoy5UwXCyjpTO4QE/divRkcQ1q8RuN
GyHUYKDQRPJDk2eW3PGFp28or+O5fegSXxf1LR/5QL8pv7VR4EOZGudq18DRseYcKeeYrY+ZToH2
BDj9MbcwGqh8dTqnDu/A/m6DFtkKFf8a+XDn1sMN/Rdw4Yhk4jK8auj7GQevzZGOwFN2ecUZKfaI
lG+sEbp/cVlbi2o9xEMh8/fJ/Gjn0UuJDYI+QStyF8no7hp/cMb0F7npTUgvig6+G+wNTEYCq4E1
vFA290FSAGREOLOguk2VetjVA2IVuE7Rm9aL8q6NVWXvRguaFLwyyjihn6eWv9x3E4TjJdlj+NjR
Tym5YgHnp1GqckDLTumL1hEWAHDRX3DxRGUL1eDj+Zzdn138f5nVRK5Mz5Q75mcYW/bfKaCfaZKz
BX/rv+YcipnvNAR/OyZkJd3qBHyaJFry5/vvi0IiKNdiodvbGbBDrnlZuFNi5rvL0cdPO50qHH5U
H8feJNvkAkP3NGZOrkM/5aTKxcmmGu5bnHisCE9lwrIdkRBOpauxT1FlvBj+5G1AAMCUiTTuOIj6
1J+iM/oLvVK4BYCIiqo4QJ/jhePEwhOuHi1xcRKnCPb3E8CVowP/40deZ4GQerUMIFd76Q7HSPQI
Xzy2rIeh/PDL+jwXVPA0peJIeE1gsoySu69NJVG1CgYlzZBddN4h2fnb5ZPyxwtnNpG0qoUp644D
Gmg5WGd6ph9NfWauGFAqdeC79jXJUleUCSWTsz/ne2kITchKh9T2LmTcJBkHImRavu1tkW65dPHq
lkOUWDIo5m85gdDwdZU7N4Pbee5IoSORSwaRdgw9EA67J3FjLAV5GMz5oc3xGjrhtGZuNycoSwoB
/83hHkNVK52M5KDohSr3eEnmD0P2VNillUy4ObvR8BMvisOcfLGujb6rUu1EUvMsTXRgjo4fxhL1
c+OfTTNb11jLG7RJdCHE91LDc2vGAQc404EULlk1cKDB4ype1U/iTV4mEg3YplLD3xOqeeeA21Sv
w+IKAMa8kNLEgT6W1PnjTshXfNa450KrNo6kceEqA9Vi7qIoUj5ldH6USk9oczB+b1++0T2hM4ix
rsy+MU4WdzUK9LSvv6z+U1H3Czo8tu75jdFOzBDdAf9PbfWNPyUz9yZGMedZGbQe/Vgx8lPL5mQP
rkx4Tx1XqZY9efPCR2p4LepTn6MArliD8Tp/+KzBQ7E9eEbyFaoiU+6ic1oIijj1R1HSAx/Jyacp
7FBpTy7oR8MuebQ53hYfz9rCbvLUEwONBsz5LdXn/TinmRKGJMFpkrXe0GQqnx33MfYTZyjZr0GG
WTxO0tG/aj6a63Ge/9tml9bX3ELNSs3WciHw4KoW+j3DtDhAyiUBGKpY3/4kJEvzFzGTolkBgq63
2KyXeL0oCvQlr8wZREV6IJtz5AUDlDOdfeVTdrNsqFB4bMhqhsHV7sDkuV33NVl0BCxwVTL1fAKj
zvc6udMEZD4d8jW5YXlejsytVjm3AORW8ukDAFBLuO5+thJJowqHhwW4ZJ3ZkVhZPpgBvdQuyVpK
UFGNZPmZh8gzPgVIuCbw0Bvzj9/yqbTqc3Zdh1pdhRGdIfTSgrAT43jhgH4u9j1jcav55P+9+yeP
Ss1vyUP7FyR09xXGqWSsIbUOV5FahcTllf2lqXevJMgs3xiXEU6QS7qJkvR182pzBaZWRyE8C08K
OjqFkZGsYopat4jgRE3zIs5iiDxjNSqzq2FmmK3O/Rh/X+vTIdvzqlJRQWBRpU/ZpnvtCAO7rjo+
WQETN/S6KO9lqEk2koixueGP6ap1aD7pJfSzTke/vKXcYE/S3W6R/3pEMM4OYz7+sz+Bqmr1ILa1
HgTX8ZCdRsSXFTTDZppRei8aEDMXJ5h+asIcaZFOUI691HNZaNk/JRe4udoCooo8gF2U8eQ4AOEZ
aWGyWm92Cqh1n+4YDaB02wAXKTjTqLsHDrjFY1Mgh2pI65NPnKzkRKa/9Y5RV8WiNzKz5uDtWMWs
zuWaNGqHa3syU4w1chjPEzwSjLSoF71O/Mpo2cRM3rCNhydEFMflqLOqoIoytVGkn5Y5ltALZQoe
cAt7qoMCpQHWJBT3yPve5JvTt1icDxC7+wYyszaq1lrCE7zUGXILvKd+eyvKyJFf4Vc8JRjeqbwz
raERTjaMF52J2uo62il1odEXIvvTNgHZbfQcFTyrlrESIh+YC1HfFlKT9rKohBQjmv2a5gVYhg/r
wFw9Gzp354D1BzP7nIJPFTfkfPQoOsPDgTnkQJiLbmfEXbyPVFMRL7eT0lxPgimdFasAT3fgyqWG
xGbhv64uq3fTlgdnuuGZTul572v/A10E9d+uF5F4bVseMAxBgIrftFaSYXpUx72zCFf6NNQEQpaB
v3twPjbJ9akcedNqn37dsU26G1h4PN411Qmf7p25q6Zts5q2Dvl9kr6Zb4GaHvxF9W3cVwYYPQzZ
atnugR1DB4PXHRPkUo89ELgCwM14nbzaee2uE92F9MKmDoOGu8+IHnUy0vXOoR0NLzb+hf2S2ebg
DkydBtZBg8oPyMLRMjALd7UI4vm7L1XB3go03F1UkPY5F0en9eDwaW9373AhalG9iod8cYjny9Bb
md97ajDICPUc0ypveJOuqaoT5XvgWpT58cxbSzdMIvHljETFPsfZxxx52GA4lvnBnJIEZwTPZl58
LpgADPasBF+w07k7YXsGhH+SHNgw9Z4mry98yblKwTHosXW2LWyAIAY2uOmxjEdALSfnDQl9cwAx
Vm70ItQf8sDUYuyGplq7rv5JGqRxWq+nL2eSsyHwyc9o2l0+5kdWnvRaQhYPeLv2m0owWwLNedlc
aoJcREtq2KKhrTZCeX5x7TjGaqtVIhhzMPOt1tgSDi//lb9djaqRIrOfqGgwRkPehVnThE4HcXxo
el9DBCm0+J2uZD6wQfglhQ3O7tZrPB/M30aDjhclqwXJRuBv1S8NqMCWu6LzdSGp+zW0sRmu+3sE
DTTQBGf3uNhAN9iK5LZIbbNuFjB/bWKKSLU71vnYC8YhpQoshQ8Scg5K+UUYQhzIb/pfKUE+9J4s
GJvdM6klQY+2JDat2YDh65Ta84gqQpK+qzrbvqliFlOBAd5OXzuA7nr1In5EzPJPTxyavwCzYaV4
XNfygC4heokr/jNFu0ncSZkALfHxzYNVFKbpNJpGEHDHK8mUiDmlDBTwD9LUNiIgYorUtJcQlL6C
iLv088JUTubdn/3CrA7HtTDWnN4hU1sNmSgRbiPuDdV28ktAq/2ezWzBrpcO06r5xm2zxsy2vpaQ
Wwx0RErYEXAoUggfKvMg/GPJuok5UphT508fsOmDfs4UecekLvcyqVfkC3wOy2KPKTKbMQUszwZF
/shsxrlVQ98lYPutXhbiwHywipS4hBLDnAJX8soqadizw6QUEYoPDJNv/eFvDKhfso1U+GCPoj3D
RA6t00di3hsPEuXzZP0GrbkfS7ahZehsjrMR14g101FG0IhCb/3hz281JSXCSHHxf+IGZnpCUfNf
04xGhbdHbtC/64ZuvXvo253R17d8rLR3cK/JlSaxRmws5wN0eDIUkUNCZDn417MpP8Gh7Z2dLRN/
RuoIvKiTo2xhqhhp0oEt+XpE9Uoo45YGjmWACYfmB4PnG5Y+0eMLzWJfEdW7fiVQi5mKDFhVD8u1
t1TgxtWehXhVa2SLSe7ehc/dLy1pZ8wOdw1vPmf97yLRiEcnlR22D0S2sLktyVAHVpEef4GWwdLc
626SU4R6W1nD/ohTHAt/Lyq2lonxqHyHV8hK05NQ+92XMv2PY3MFifoOha3tI58d16MoouqUxwAK
u5OsDyiO6W+Qv6jNJgcitwDMwTjJnxHvzfrpZLD+DdHl+aMOwu+h7SmqzC5Fmw6i7tjh00dkX0An
/tZyk7MKKvgP5bsUbZlyQ4STWDoN/V3nSBHpEs0rs6/kIBnf1c9WL90vAghW4koZteR/65NcygKO
f4oDLRUCp/yAxpXSK7zfHBM9adCE+uISVuzZiuaRJHkaNsXq7UIZo6bm93pPE2sUYM+XEiYcjgX2
NghoEiJPogM7C3icEFhtq9rUQdL4jOX+bKfFwKoIkVe35pD2AHrfhWRRn2VVV2oi0/yfGN7wKtZ2
xzmGrUM9DnCbQZL6aG8R1uJJo/w1goJxs0vjjKaD9P9LYlMcVt4fHjDwRNzuWLsQ5ZM/Q4NWhJbz
1jARPOfYRwmZC/MOD7pgB9xk8rGqw9P8ea5zrGx3oKYz5T3PmtJXo8PDzzt4gS9AmZTe8BY0col+
ElbAoF0tpCHViHWbAW5Gi3a8OiJieQoTIY5umnWfMXJ2+1BeSrhNSZ42WYneUxA2JNyk6RvEEeGq
7vV//+R3zahk5Jk9HP76yngu08Q5VSUCTNSMmOj9HoGsLkWDm1PA1KeX+4n6wuYnWmCX281cGY/9
i2H3UzbVWbUbn4SS3chPZCJ1tnZi2LxYwv1IRWgaRtr/at5CQCN2EjyxsvW3U3K18xzTI9geecfa
/ti05jUvoCoTvzFKGN5KIurjcxRzF+TXGcOsdAfENAb3bwC6IFrEEVzLAnmK1EPDXrDCVdDQK4i5
ipAma7R4aCbxMs1MePyLiGv3NAzYStLrzbsywnDYJQv0TRyqaOfYxFo+a77+zPlYjX5s0W+FULD5
4/a7ob0Iec0PRf/nT/d3r0zHf8fUzrBGPOuRmZxMYjP3Wj0N/zuTngtbBez0JuGi5zPgOwce8uNj
lwt29dlheP/1EcYSsPV5vMRYbk4c8gqnsrOXwNAxNL76PE8x2ZfHRo2w3G6ohetKqM/Xnpk8bP9y
1OTwEjyCNbmXmcs70D+72OyCPD9i8rgzFLmWj7oPrnZFT7P7P6gt5uNppfAiWz1WcH+cmUtTYbzI
1VD57lmJYPtuSjElsNoaJ5UcZp/OKGhjAZgTTmK0Sqx9ctBMXRcXYc7JR4KucsXCKz5t0D6xB+7i
yz9n35iJU/ydP71tCgarmBxl8ueBB990kprpylzxGXoC2Py7EJTbrZrz8KoBqF7iN2i6f3ge4Bct
rxPYDbtveLjsvEvWGFzx+ITlUkZpZZexKEPCJGH1sv9K/okzgWiJqqYRliMVyDaFwWFtXUKgl1Kp
HlrL5IQbX7CPLMxF+qX2PBZZYuIPbO9aG/8Be/G9G8AxLnxjatk8EDHYONhT3f+Jbhhtg47394dM
lNPV+iV1LckDzkNoPmZqD0ZiqJARVz3W2Qi84KSSs7mk/zyrdfE5s8RCJoI3ZeQho4Xb9CuPWo4O
dsZ895V0oDIHAtplr/WfCWLANSwKA+vTlxcbGuIiWkaMdwHB1GbPOjITkjE9NLDBk8B3qbTRnZlc
G/554G8AEfKZzm6h5dCbecg/OGoN7HvjLQN9z5zUSJOxYcnm6Y3nrrIs6CYDRvwnxxzCJ9Fs+0rO
Ip/uddZR1P2jpaLy1B5GCa6wLpqZGPdvJZpRdYSWhzeHbJgsOMrVqfnbLJPWU/hKKBsllZweVnzK
SSw6ZApcuJ7SOQBGRc4mWDcYAgTXW7ZEQ86qvRhglKvU/pgFsYNnfwnVqavJD+Ghy+GYNO3D1BuR
VWRNEXVMS6b8HeWOJt9JgvlpNQhwQyQh8ZS4Cs+jrRrgE4L9KbQ292jDJ0o+7pRzxRue3MT2hffN
Y2Q1RzpH9wAVguGCV3zDh5QNZs+qS9WLyYa2auSwwT8wkgmQU+1EkrgqHmbnPzSHfQDTpG6J0QVa
s75nI7LO10Af6Zjvh/JZkHF/RWiB350XBsaxegOXKNAaFLfLXey201/g3dFvAGW55iMbztTFwEDJ
5+maSb0z/qJyEWzVhty18jnbYovRsd73FPW7Alv8F+uW0FQirkLBkKhTjcmV20DuducpBG7zI4nU
trBn1tBLcNLyQZ8HIxd0zx+BS+AtSRGKsejTulKQpL+MUusQCyu757yrqpVmM9peOkrG2GReuCNF
UZIaLlXAZK1o+A0+O5NBqT/R/gedGeuwwES0q/tYR5NvJejCEhqIvoFAsWvAqS6gA+e4MVMmSx6i
G9izermUavPfG1pYWfrR8WIt98reQkMUNqoVW60jx0vzx7h9mintC2scNvm5OOjiFE3EPEpiR0bl
Z7SDhq/pk4yIAMwcLyidGmGjpYGPbTHREdCKMVkO66vxyaSkwr4bCStj+H/KT8kWzq5N6j8UrjbK
QxupzEsEOpduCNZiSD9ahOelnQcI6begYO02SF+uuF+NBMx+OQ1WyOn8mbcqpgt2lInKRxA2P9vo
pWU0atEOcpEsToBghXIlj1bJAfFuaShTc6Gq7nv4bOzJJmN3Qeos7pD0ClDObqS++89NIFEg2lNq
5R7baRtQco4uiN3asiMV76dFbCHO4jHv19qx7gf8b9JD3eTQ8uGJWxLfXNM2ahByn7xdQToT0mqF
ujS/lgAo/XMLkmLTATrveTr8DpFTUZ9MiBBMe1VWpZsCh2YvuIyrS/dSQ3vsawjOOV56lwwF10gw
a/OCHnSgsZliUf9mXPUXUGmadVaVbE9ByS1dUFxdthEFrjBYD25qzxgIett+wFBfiHc1+9r8JxfZ
YwGMxR6nlqocmr7OtkTBmDZCLQFoHSFNvmEXBatQCsDWv9AsSDO49UUiUuH8BnZ/ToqKiWiuoa5D
xCqnXUxKiighGwjTraQ8juOIRyzGxpYf8danPAVGnsGQ0cPaPJicHFFRwwFM09G0EMmU55Xl+RcI
fExE36Cgn/jkMiJmIVSIpWHEbJOmTZWnfEMBo7997cSRQr8wcMRSWL5D0dTU/PboX8Q3uurwgsUs
Noo8ycpM84kfp1SS64r7dfm84oVYTO1Gle53zKQSq7o2C/I5+JlpBn+fyWZOsZh2vuWog0OtLMED
2Xc/gyeaAfR0s92acS+eiv39FqneuBjZx38S3AhhOpMx0n475VWS1kKTTu/Pql8Ge41vZFG4EeX7
DUF9Dq9q3N9eK2NQeogdpG0/Tmir6fmKBOlBvdJVM7Gasx1XGCzxxYv5EtReSy2JiIDdnpg+lLTt
P47MC3qpztJCO2KLlOlpAYCjtoAERFLxsXhjqz1UbkI5cTHcE1RdyHTC4sX/rGlD++3RXARBvMZW
DPU4ONQCkVPz/qNmk3nvAfpeS2iHS5mNTLM8WVbOYYd745CKlqO6HrjNc1zwSg7STk5Dcz8IVNd9
UlgEu1xfT1NrwFEyiv7CKIx7AgHhke/QKWhCzapnaIE77lx9eVH3HrOLRahcOE7P4wHlM5WwYlKr
1XnBmJuSIFhr09SsPcKm8PgsJenOFauTenLS5xM+YJOEQkqJhaAj8OiG21EaJX52C+p7rTP01Iiy
bpzI25yk8daBWpB0fNhbHTTLvo5UVthB0leMBtIyeSc5sEhYGe/DrzVUpWmFBRBw+ouB/4DM5RyB
tQSnOyuLqaZw9ayFi+OT0Gi8GvZd/5bMQjunNBtj9rq99Rh01buotapahWD5FxG4QfkWRFlr12fW
rMVqFNcpi9pgKX+oIcq2wX2QVW0G225x6VSddUY3jFvUXDO5Wd0y9hP4ka42tfYwaNwZ4YDl1ION
cBsuVn2lgFQUDYmjmDLjno1aIefwhIEEtYTs6CCUeoptb41KDjSjRUcVTVFHtofaAeT+6+LBH32M
DVVY+bUxH0Qvx7ECug7hbju8muKXP/mHX5ceWi2ypjRDoRnwx7IxjKsggdK1P6nN0XAULmnIZMsW
7Bq3eFgL1o0IKIcpIiKLNTs2bFdkKCpUbwk7nUaGkyhBOqI/dzwgUnCfN+qTj2Je5qKH8vwS0pD+
/RSwt36neh4rMjSB36mM5MIArrvC8+nWZ07GRfqJdp+/3cm43Uy942ubS/FVyJkfAh1gCEOQvAYa
E5+L2BrREg5dfvgMmITF0Xsrup6HSb8fWez0L+zOe+R+Dxm33+r/UbxLouLQ5NbRDOeDNX9yZobu
KicnCP0c12yLMDRecDkRH6bhmxxH9A9yGN0iZVQshmY4AaLyj0KxsOzVoClIVx/EHIWDR+nsDxAN
/xugWmp586hL3eFQ8sEXXI9PCfgxNYAHNDvf0/qLBDI5vQa988IRrH2uvaIm7SYn/ubdS4bNBb1+
/rJrfQuIBTq4y4vIBT+QSuRO37hvufYkk4Wd5GyoeHEJUrXwoAdesJiJOEb+V8rro2oV/sCUViPq
hsrwb15Wo5GJJiWTxYqCebhkHV8ZJxYkThbwTLZV7c4C4W+RzcFvOOXqcqEUIYt4ADYjZMuFHfOU
Av65Of2pMNbqtyBZjYQSb/3x8lk/IjIJ1EC3CJblPrJN+FOMMLP4edE/Tl6gj35uQH6lnNbMiYBM
2W2yuqojy+gLotiLwDYCUvqAUCDf0O1n9fXrAPm68gcGMqF7t7NfPemj3axV50iDkRoTueQU+3Q1
UYmvNHdC8Qs/syVjkJlbOMyD7BQEiOBIV7xv/Y073OWww9EcST+OAOVWgTieaqpMGj1/ZsHNPxpB
AbaI6KTHnNTdCdKxYkuefJmF1eZFy4Evql2bnrtxdlb/IvMJ78eyPvBCXkKDDgLGPsQlSIvyQW+X
sMwQNmVAcrL1z/yN8n88XwD9MF5jh3RMFc1XyI1pJv+VLcawwnwY4EOXh3Jq/htSeNVex1KHarEO
hCB6JZHjAylA7xFLCF+UAvm29W0PMpQoZKLNKgTcnQ9ypeBwQs9amNmDBLtwvcaUcZGoALqOO0iG
dT9i2LueCEukuOe/qgGryjupMyW3e+3DxqCdn2BR3TUiDNXPTyvljdMKcqsU9OfZbwmDnZHzu/e0
6P1h6oVcYdp5bi0okejzG/rXyEpaPaRbYpsnhvasnuaKGRxVizPnEFHdoRRgWPff2R0lu97RMYGW
+KbKGFbY9pzSsBkFn2vIR1nzut0rMs3E+1SCwIKDpP6bzhSayAkxHmb4yQx6+10T5QFNGjlkmn9i
v+ZsjZ9FOnD1+QeUbfvMRlYuKJxm9PrGME6q/8RJp8YFlCMRuQJd5FzbMrNoMgHnCXJcK2/5Y0+p
BZj2Np8UHBTeRdqcskQJLWcHlKEYG9N7j2hF5dSkwGpeYug4t6dUQYLRanDrIV1Ip0zJXrmRzZNn
O67inXDxNgk6jzU6KsynHUpu4NHJFOe80ICkRQP7/D3uEAxWULilz/dQYBfLQrtKdmPw9uRb5KcJ
36h1owTjb8yaixQZgiky5uAqtFHw+CrNGUmBMBdfQ+HL6o+KIh6UmL0UUKtke8lH7caCBWZeS/wf
5xgsvOCWDzni3TZaXMvUrOo4KEzf9f5CghxJchC5V7Y5KVisKHJj+U8FHmHfLlfVx/4zeykTKMvh
VHhZii+t+9MU3QKljHbhsSQVGx/LA4VMT/z0ENlu6wSfzz+0zBgRTK/QW1cjRd4EEDW5E0lBDYeU
SSRseA8a/H9GJBq3Ku2llYMyr8kt6pxygJd2cU1HLxAVxIU6BkJY72OUAlq7fuqo0xJjFhquxMyF
TRvooYpRWbTHwai6IK5x21fus0WvVwI5SNiSF8Y9mgC2/y9K2JrFO5DRWAee0cR/Uz6Mv9nxt22e
IJfKJUl5h+YhRt4eqO421mBG7gI+SN7QQW5Wq5yzb1CKmHsFGdEagh7Sk7kzFpd94WpejYt+hkxI
Gfwsl+gTE4uTxKIJH3/CAbybEdQJLK08GHc4iJ3lShdPF48vTwHrMAY30qwetBuOu6h+1+ksRuPN
sDS/DX6yZ3pzQnlEL3aCXxRBP6udVGrQ24DO4aVIW4JiPbjcWDPQ957KEEVYrlj5+b9FaW1cBpdM
ojqFjKx/D8JV7mzcVse8BCg7UMbCCeuLPwhkdC5pk5JVInEBWfxajxBaO9sUPpK+4UCW6ETiwwiG
k+lAGQAqXVIwCVDKoGwnCld42rrTI1ZEpyUeVow5rB/C1exsF+eEHpzXxXUnoEOC7VjTvACL1GWg
BQxqeyvefy8r53UB8qt67nrywvzf1VdNhAVgxD5HU1L93f5Um0ddS/ogsL/nXEzpmQ1+U9gmHlZ8
k0pMGMVfDwQNg9Dhpd1bxZz+Ni3CKmmwjimUZ+mcpZoU0pLg06VIpLJXsPYu3JKX445frvVBC1WC
haNYS7RVWFPfyL+nKZmBOM4WcQ2oCTfL+aPBJh6ihhEl6oqrjCasOj2WXoQMmGs1HqwuKAAMLEHV
H/0s7ETbyDj4ww7vORoaVvwfJbedhjG1wPnD3ngOZbNbQjDYRpcUDhTf+5RalyOW0M2MVm4lC7Wv
vnwWkIl8wG5zqoI6na0ZBLPPG8o2A3N41LVF1cSXVNtXyS3j8F6C03v4BC98UlE6ZNHbgNy8VNy5
XoDt4BG87AE4HSGtCm+xVFeHGBXBEQGZWhmm/4HBhfS57ds7PyffZGYjm6AZrWaxhHfIA6Ee8nFq
eCE7YgCOrNmBH8mXb9ITmloRcSMsTOtOt1zXvLJdFDzr/WnsIDRwJ+YLZckYKWiIiH5+oS3rjk0p
iAnjUp5eGrNzEPnJJ/8YBhZx2lJV1CBSDBkEpO7dR20NaxhOzq3dr5QkMEq8jeCPw5+9WF99n6NZ
0DxdT9BYD4XVJ509j08wZl0aNh0R9cGCnE9B+HUUTZvCIouvoKnwtTbcqICexr7Qiz1/Gwlp3ynB
3IMrt3Dgan7ri9KEsN9dNy6ArY9E5HXvomjE1KxwVDcppotwoyB/KLjUS2oeT+BISvlUJPHRknb8
kMVhOtYAW/OQYGZWh+cpFfWX0P28rApEea0Qd1XrixfWAzBbq5cnzKWkHfWrPDEy1sC2XT9AI+la
WMsB2adz5QYEzowRjHe0l99mFHszJE/XbRG8J5wXAnSfyMi97ZZQ/Yl7kgSgHRMxp6NkSoDynsL+
LrcbOK+G8jXd6apfUZPyscKLsuj1/6E83zbjXPY+DU/QOwjnHOdyvGMnT73XOUco88v3S61/MWpo
i3QsBdIv4UFq9qjSO/q/1fjAXNqX7h0IbqvROCwFC2Q+uhywbg2thyh+7lF3uNQ0b2EvS+tc8wCy
F4g6yrbQm2h+xAK7Z5TQR4jlwbn+ok5nlzHgkQLa5DqV1ZS4sAaUJvk/SoxOC6f7+dk8eOZmLbj0
54pZ/L4lAnvYpusfqc+n4dygpXRmzSR0HLeTw+2PqjM8f6flAd7f9qiiH9gT/ZaCt7srmZPH/vMZ
mqjQrd3G9K0EJCz4rcvSJcFPMZTbGu2z0SOmLPOImZOSkmhnR5z35h88RUjQyR2cS0LUFQPYt2Wc
slxTrOIiNv9dlT56MlzbwnygZPm70SL1Ni2UBV2Be5kVQzzxjhdx1U2ZhsjU081p2yxD4LQukUiY
FTFVBFy1vc0HrwJseNHNx5++uhJ0eQDlruLv6pMozq/gDc56eD9haBifLZEDVusq1SyG4CnZvE0w
BZoKHMKVcvBaG4bsS+OmunJGdesCpdblcHb9U8Ug61bNb1/kXOg0Z9y0KpxRXt/mgmTTD3135vAp
Yg++ca1L+6L/QwfMwDy4FawvWOrwuLqXkWJ5joCaEkZ7LGSut0LhusTH1d1LV85zJ63KLY+OBwAZ
kA7okqrzr38lzecYMQ6VqamYrt0rBtND8cNk0NelWrvt+QY3wl6B84SN6+sGIqgGfQuZ9DAx/TCj
ztEwb57sLo8kk7+Fbvvz13yB+vDvmiZ8P/A5JN1BCX1h35Ww/1eKTKRKChqUYkSUzQBZ5sDoPgJR
unc6IkcHxqfAkPJ/JZ5oPj1z5+C2tnfS4YvSS7h4JfQGozUdxH0VCbvd2cO8Tl5vKj5dDXX+eFPg
w9db3FdNMXJhCnwN0euoHBP4ILUHhk0RAJA0lvvAx5lgNUs71MLDPMsqf3lSru10nDbjAtdsKBZQ
1XbR+QmRaeAbse8N28JoIxJYonuIdhENnXPQMx3Pgwki5eyTUb6cBz9AiYf0G+xIWOgnknZhHHiz
3C45/lsr/ksucY50SL71Vc0XuGSI2mM+NLunTXhuGCUFycsXAKcgtoeZMEyfr7Kw3/8vpOQ2/rpG
xfHZyzAMBqie9sqPxMljcOLjwqDv6U4e2x9+lbxwcMqs5XfZc8p21thIq1Cqdtc0kT8tmzSBPgwv
I4tFR4ZZLhz3Tmc5zo46+H3Sn0A83GXKeRu/p7CbzAy5p16q8OgJ6M3FMPFGhVEdpr9LnrOcB1VH
fdrp/mFGYjKndrygb442N691zzub5jUKFW8IaWATbumqkQ7wHZLGFj+6RDv3BO5e9emSvLlR+YpO
LYlN0rrCQmDePLNgnX5ZsL4bGp4gHVvHBpjpV67aJhSwybriq9jUb7D32OUwMCsUonhDtTJqI822
MziEFgtjkPCFbbXqsZ0NjTpMEbdJF0fGzsk4rOrtbbvWkFmRL6YpEed4W/z2wHUD8vSQdmyEDsb7
VDJ4Kn4zwRTaD9YtbmTU0+nqAmuA6VuriyMq8atMgNED9JIeyaqpX9DYzL4Xk1u51A9l0yNcNjQQ
cd38pJ/0Dvcm04y60Rx9nif57MaR7KRZ6z2MTvZKdebP6socxspIOheVPZedqhiSGEm4afMSVqYV
OMEQWaKVURAB4soZcCQD+ERR60aXOmKx5UQ5dObKG5Xjze8O8v6M1X59bYsRKcpQ3cVinQ/eKV+L
huz9000vOzp/dnPA7wbMVxv1rtKjnSUuAbdSFb/6vpjjYiWipolsOJ3bMd8y5PA4lHOu3fAeOkIB
mly944aRdRrXPw2GCycq0w/vZuKtRmZ5/Sv4WjFa8zKaZvzwhRwVSdyJu54LQ7D9TNjN2PJiAZt0
BvT7Wc5fwmN163LJwnxxVVm45ED4YQwFTCqvJZJFpNRQZv8xZVA9WSWocviDL7knVq5wV+AXAfOa
U5c7+GnZOj0Cn4ynium9PwWueEsCXRZnf5aPQoi87zK9l0uprf4v+Jmj71YIFq6D/DSFY2oR/Erw
AbatLkfHc6IDQ3eGoiAnNlCLevGNkbeM3VacQ0X/09/xUC8PPiyJKXUJdiHwMkxHYn3r24Af80Hg
tFOOqIsyv1citSAfhGmqvsgxFefSqqcqMhSiu2Vr23PRgVQa9QqhXe3aTBYriIP6E16jBxg5wN3a
EZqEwvNFLVmDl4E9BYHHZLDUNXSo/XODASbwGQ4MNNd1J5+yGEsFlySIrRBMDyszwHCivvSLBXc2
i/C9vIFGNu1nBcQ3BcssMn4XCRU86eP88at++orFGDyZul2/TEfkmHGGOzj2X5z1mRdKzxxOTIPy
z637k2sUDH0O68Q70v9fyHLbeyoFiLJRu3NnLs8SoECyaMeqMm2PDgkF2VD8gzLc/wswf8KtbR77
eqpWsy8Gsb4kRD7rqlLxWn8daNZoTeAPsdu6KgtPXBHh4P/VSbVPhdol5ipAybLgvB+MQod/v55+
yCShex7jOmQaw+o8O/Mb4t41CbVir5e1hUZq+5wxA/57X7SwTJMsQEXzSf/xnJOtF1rbikOIlQDU
TSUXx/nPfiQgULNJX8YFMe5NME7CKoKpVY5F0OlLRVpfvHi9CE/vfQP7OtJSFvnVqDkNNFPykxoD
tbn+zIUWFTr0/s6QS/+DeEDWIg0IhSfT8CU0WvCpz3//Tzdpz7e09g86o+gRl637ctLdo7vKUQrb
/rhbuC+o2KkRUa3o/Tvi2CZQrOCYZgsFGfdkJrNvTTI+hIqpnAKRTYWs1s2Awlknp3Zz1cQR+GPw
zHbOOGGUKWIGq+sdECthlsnKcq4hqyzX6qRc9h3Irz3hA0pEn7IobQKLLJB3bxzjlyX51VOhPkHr
DHLDZydAYWDcTzlbO+9ZD5IQPg+9IdlsmTC6u9Ihj0t76GAck0fk0aNJrWmFoFkc7yWQiBuHc7x8
pmcorA8ZkqrMbiCSM+gt5xnRyRsWjHehl4XKKwqPmaGhOvMYPovT9lBnqWwMX5JbAaNrGfcAuFxh
YV2fKpuNCxrGDJrYNk6Nf5t7MdOLmferwZPI/TeTEJtopwgcCLDBLVWIs4OUGWKpBFGQuLJ4k/kh
bMScUBlZOgSBWbs0JExuAQaEy3XMCwqlbrbBHkGMYL08RCUiCZv1MUtBUjec6+W0Znmsu3hOKcjg
veqH6Gsf4SZW0f7IJrt+QP8H/l0mDEZWf/+pRfhYwW9hfKnbqL15JmhhHB2QSEnjup+uyxqX87a1
4ITczsmNgTWODMh0Bkrv/9aYjLqdT9y0OW57ELwgNIOYNdUfDyQU10d28IMhOgl0un3as2tj7fD7
2pHxcwEyOw4M+c6bcklFCgOud/JmoOapkorZzzl9NjD+OuY6sWZl8CRj3yQ7CUKjA+QY/q1vP/8F
R9Fp+rFGprQeAYM+cWO9CNkF/USbtPHJ84vM1MUkDDNmpALsWhKnmODRUaZ3dKWq9VQi/NHfSXUc
+yuPyM1v2LuCNq012FLMOpsUAMncIBVAIuWExYxl7z4Mo93SeZgLxJscGpTdgHgcbf+Y0HDLAwVs
fWpL+Rej0kDx6emL5hEuzCjRrB95S5vxlPPSHtOwJ9MeHPC2dtxr5mp4N93F9K+RImu0KSF0pn7K
ooqevkN3mr7HmE+JWRthzY/Gt/QwI4/P+fq0GUpAVYuLEK1bO2UT+VKHgFfifT6Qyw4iuEYTMS6l
bwdG6n06cjRIbDdGTNkskt7+YRuWx8FDUyAuU9qlL4XQ5fqV2QHjHS8wos3PJTlpTSJ2hh47Kw+e
1lfucVVGtPz4qPIar9w1uGtYMOov+rFN7r1En6sPYaSlAJHNL5CbXpBX3X9SGYuWwWxllJICq/ZY
XwB9rSvPjeUnGHc68uiE3hBN/ua+9neo4R1F/3Phic9Ed/mF/WueTjKZijBOKSu8u/J4wHGe6Bjn
c7+7lWwSOp7xS501tdNWaltwDXjWpF71jCny+3L6ie6xnQnmVv8Iuz+zmmRbsQsgczUIvwuvGGRt
afHeJk7PbjNEKEnDzwk8iykDoUBZUmNuEA7f3ZOWZ6+yt+v3Ku5y8qj+T0eB4/0kto26b6VUXaq2
lgcakH5CfvIdoHuEd7LmdqgrkQKVdp4ocrF7Zf/Uqr19s3eGdz8h2Wz9jbJgv2n6HA0Am+WJy/uy
zwEncukH3HKFdp5xVSkGtKkhMxbnNfjEsmmIjd8Jdwxmym4Nij+V+eJ5TBIIwNMyC/Ow65cGfzz1
s6gg/Cqj8nrrTT5xeNWyYw5zJe7zjl6kJDXVr7f1LD18ifNlcvnnwb9kLLdMvHr9+dDSgXPpy7Uq
DGuJf7rMo/wKtCWQfK1R5RDqknAzJJ8RPCsrRAhwGBAt1XZgvp00xRTVw67lvfnOHcVcXui89cxV
90uvAH+sttNEq2iE1SB3S/CaJbrYCKVyoW2DWtrlXJNoYHDyI4QwOoMbSjuKHVoFoLbEal/OCHIJ
ufh0IkeP9NZOMcHE09b1XoXUPrXwgXkOHXCWhdIB+hRXI0FNipV22m65P4ERzOGKXS1MAvBGA8T1
TVaNJp/wOHuGJRRt2mP3jBQB+IgQYe3j66ENwnk3t25vf9a5h9sBwFOZ8h5gDpkCKvRNpNP5ppOZ
OlrQ/roo1Sy3Qax2jz08vEcXxvuRmp5CFt1oLnPVhhXYrjhpiVjdIUzzK6zCWs5CgHV03EgDrd7t
yP120XAbXicb7MxS+d4+ikPyPk0iPgdxfVrAHoaWnbk4IL82VUwwPdPCmWSQFVO0NGTXe963CXa5
5uPF74AZz/ed8uSOWHNe0Kjf6ltDngFMCXZ0uBg7pWOWfiKF0p1WqMklVF0pju7x+ckrsaNTscoY
4URGHBLauClp/6zQuaMcYaUCfpk4QXxzlNRs7MmXfafiBoASg32HHAvMH6aY+gOQQpfsrYNpzHs7
H3U3FLCKYfGEqYKHf6d+UmbHcQ5F+OQdgNhlFWD/Fc1wi9QQZQFK7KqzeooGgDBURG/dmvxI+yyM
YpIxzhlCT0LwO/rMV+JYqO/grN3XDyxSmvDBRcYjeO0pfpJPhCYnBH95vL51sLUZONgjOuTWqlH8
GcR9Kkm3U90duJaiecSWFCpq+5OcwuhIFWbC60nlLtR7Bf7/i4OqYQ8OzrJ0V6xhjlkGeRAON+iM
ZXHsbW0b4YSIYrVepCjDofaFvcO0i5LYHRHjd9NRZnaMuk8lS9p7cmHhtEF6ylSACkMPXS2m3mYI
lwaPmEU5QvfMyMc7MJK3kCvxdN5SgRnODDNK5JfYW0xq3F0OPEhA3lLV3SGy2z0qGDvuKnLZv1dh
ef1lCKWviw9seEsaksnHTIP2h45RCmIsq6fGDHuwFJ2HcyyQH+jIAuzDh9+r/CXZbL1vrguTa67C
E6EK55yk9wya6m7XS52kwC+IuZZfAgHbVhrtNodoYDn8sDLppmXFVD3ZaBou7aZG4PceTThfc3SI
BmnkVsAiSzFx+KFKR/VEpPFEJDI0+U2xK1hMy+SOoNStLZj3paMbQwSMPzz9En+9xMszZdk63xDU
yrb3Vevf90vfdTestLoo4hIpvkyyQnKSqYJaD7rp8TpHrkQbbq7K924hV9M2mZUeSdRzcwzRum8q
B1Zc8PfRSa4LJBdpVlv3w/lR/jvwours+aSE21BLJvRaRJ41pLu/ftFJ5ZcUGPzq0gOCDfOLrepO
+qrdYtasWUa4vimM5ADJVi5j45wzGs/qJlSa6fLLFnrXXP40LBR0XT7Z8XTqlKzPtmrTUxoY4XhG
9W7oeWROojRjItu0KS5+Ocq3pkCOA3WWDDGh0HfMtGnSQqEq0I7utBHKnrn2cOanzxzeZAClLDbQ
c6xmDVKz3Ci8d5zitRTujyJBqLpsP8lHs7gVLclOv+bhnny2VaudYmPh8cdu1k27pPAz3VCw946i
xwh42F9MO9287q2klZe2D+ILNADlyQYFMw134xo9P1Z+x4S4GL6OD2p4y4XhFfVkp29Gw66awcq8
t7P0Cpy3buTdalUDBsI+Q0AD9KrOqehoSfFFYh/0+JXSoGMLXHZcfOOOqR7qB3SG4w9mntO1Vbuz
Mibq+3lXDez1aSmKLT1/pyMFtVKO4YV6Z4uVXLC2Yoi6shZ3GOh5+h/GTBwAN4d/klnQn6KcHbGE
8OpwpkY/BCIBux6iwno88alhT3Ql5jgnoGCQOHrLY1QOcYQPymXVKRxDNTQTCa74idMtmPADp+oa
FzMW4Fr434LY+78ME2D6t3ki92oeCNXeD1qdW95a53S/BRMA1dFgE67p6tFLGJjHVjmG9MT+Bivr
FEfZX9eX8n+30TLFhTMyhBBNwHDIxTzD8G7Aeu0x6KLxwQjXVULXtN7FkbkRBkzk9oD5WibMxjpA
JgQAScjGbM+mJlpz3bPZGuN87pr15ZdkRpxKO3+kOiUrFdHhZ/zxgdWN8iVr8z/ZJTbhJfz5p+sP
L3Z4HsK6EqHqtE843+2xgSudEor1INya48AxJz0Hs3fbYaGt9KwCPgJ9hr/3WdMCef0XihqTED2Z
vfK/cNpaJ3nxbnc76c1BtY1Avx1ZvVz11M6sd4yfNwE9RM622p1TEZbVAnwQVnsnciO9IT4axUhS
zXA05a1g3m+mhRNlEb02HZArOvnU/ymTqhC6XI/gq2VqUr3ZPy/Z+9jXYJZWPzg7w4mdAZBc/guM
LCvUmHB7R8BeKP60nhB/MmPvAvSHXTXLrrrBa0dY6ZTIxugwJbBXM0SSp1UKCflHHP5m7IcEtUI1
/Di5essWkPM18Flw+iEFvRYnG0C3mm+7bI7Le4AH03yzAh4sOLIghS4eqwgWIovkbqeD1konY4IR
J3Db7zTF8T/m+W3qrptE+jJasGs+QzBn5NkMGpNAZ7YnKGJcADm1maGL9HPhHeRAaNy+jhZ4xxy0
29D0WKQJ7KuR04nrx4xG6HuNjePdg0VhL5PdY3u8s6cyOVSZ6aVk/Fmaif5fmFZOFL5HBsKv2Ast
8SbhSpLKvT1i0QNI7BfRU8/e1ZWWdm9qfAB8mF8YYITQBGtjIoD/0x+WMyOGBaSQEQBDjrCMP8ZD
Z7MyzHTrDy/c0bCOFDiNf5476DsQsbYBVbvlmVP2GgXBJxllHLQqI7RyMIa9kgh/GGYc4dqTmb1k
hBAho6GDGzYOJrQUAYG+vEOjJbdyvU4zzVNN3wRMfk4plmOucdmT/dx4Eniw1q6dACbiic0sXvYs
fd3PMO/EcTygtcFS+U4DcsHgB6sXL/a7fus064Qpv6D5Az0BYUDFjGmFqRMkPjN0ccGr34UPlywG
RTe/C1WegJynjdDgzXsaIGI7IfkB+7h7Hxnpm2ZcAtpquiBEoVnCBTrrdgX6liAGx9psgq3iW4MJ
a94XfJZDlWQGAJtDpzxjpEFaiIbIr3DmIpHFpXqJ7/OQ93/XXhGf6pt2Px/5Eqlt2s1vSbrK268I
xpbkGVdiVpY1lCexD8ASOFBgNxl5bjTm674Is+iM/0FADEpdFPaq3txkBPplKLd0aKOMgyBFjpie
ApIuoStyppppN7DCRSwEh8IZedHqbDnRW0Q8ptfjoF1Lt1i9igttCUZiU68RPV7PfrOBawT9QS4i
xzwVBdtkDGh+lqGeJ99Et4mUQQuTgC0qja/oTL3pm8ADMuU9e19wp9wNK8n2HWVPkmMYkgaOFhyE
l3cy9lNQKbUxycwjEghKM5qp/+aY5uUOACNJZHfLULlIa2JoIsukUudt1HC/Y3sK7z+gDPBwxW5M
tysNTR+jpSQpJsEnMcmM478DvKeTYSI+Gli8LNZVdTirsYqIvFWvclbn6azxr5xVAgkkGZfu9uYo
mpYd0R+evLOIIp/i/WEwz5DQnRbpMaxEOqKdgsrMAMx4Yldp4ZJ9a7rQJb5cnLD0ppeJdyvk5wyU
SIfEoF9uKxWAH91P9hHqN4+liIE981cnNj3xMIgHVyr3ujN1d8p6VGeOhyPtihV1D8F/d+D6flbE
TBKAwAJ4XGBwnXVxE1l5jSWBMwrWRogCqJEf8KClWW7QscVHZ+7wl3ZRMqwWkFqtX6ujcvvSXG1n
gZ+c7ngv+wm3GE73vnOTKOfVguVyQMxV0VnWnPpKJG9zXFpvUDuy/Z7bRHIgIHDH6tdozE/hmd4O
Wfhssa79Oyr3cEO3niquEcMTZ7lj4kTpkDBLhZdjQSupaS7++E9EyumwnD2N/lnqCAT6VBwloNAr
6qtA2bcuh86sXci1WlWcAnlJKGBWQJiiNFdKM9JgYUvlDd1NPRMN+5eG/DURY+zZxhJUGNudqrQd
HF2ZwqyVwWZWBuyu6HHEycwSMbK5subX8ZznV3IqypjVke4ouK5emriRpZUhcf9WbWLVRhnGCAGS
yABtCw9Xr4tYEys9aSVznLxumIAOeLruW/zVGhnuj6bEEt95O7VoUt8XKBD7pYLxvXF9vAsEiraP
IrjZtbAc6XrAHjOjJR2aQeHEWRXBFIHkLDK6C3mypitOmXK6KMuTMrHC2wyuM89nvoXkjUkw76I1
yCINbMAiBIUVrOI/9pcH6oacklL6plkb1aenumvDp940vs9v4kKa7e62DWYhwzTfM1Bdf+s5ZxbN
kZiKJKTdB6NpzXCci8axQ2y/12fZgVH6RA2yAJGq1jAu/4geiIi5mIORQPrp3dG0oR7LTJN2N8+N
iBQJYuc7z/njKjtznJOupiLoI8rxTjFcDE/U/7BGTxgcYu5Sz6hOc5T5GCgRdbkGlVWNcOJrRZyv
UpKf1sh5C2+c15eAFh7lSEZM4cOPg5zP2uEC/k0AJ9hG7eMbMZooe2akZolBTG82uIx65+yg9Pcv
+wTQxSTviPk/rb4bBgVV+efDHNnoDk+tvUIeW+MPNOeslHCIGse1vq11A1yRthSvzdZJFon18+R5
cUyghECFwjAuDbVTtWu3UuljZIBp3BwX4QOznk/2xR/wuNpaCnH3I+Y6ojA7tJOASkNfUgaTju2g
DEJAezQybwJrdpLG0lIjb30FgVBV6ApIlNTh1zbssLYcz1tPSLisnz4TRfIbq1ywYD5R3Yxe4HGR
Dmagjh0PwJjaP+Uf969Ryk/zg9VRf54STXSKA2rPT71pkzsBeGRPbkGYlFLW+rSv42KD/26MzB3h
hTNxVDKTzoAoUW02/3YlztPA2kRbRSJ58Gvh8B/s4LwNfOcqhNJ9MU4MrtoNSw04CbCbBXLvaQeX
L7Qpi3tLb8qIXPt4bYMTce291bKc5Q0kmQ0eDjZdO/C+wMSaZz/17qD8qRPTz5wdaidy/bIv8f4j
Wx2bxEvemSlX6qr3Z1W5mv+J0XLcDTZL3aHPyOcPleJKnh2uWaRNvy2MLcmIjX88r9GqpOD/9HRo
RzjvlSQZlSJj1HXjDyom5DZhQsgpBblzPzxRjF9D9pncfzFxPMHwqB8BFqLJyq8wINw1eAvr7qyS
zMl2GNfy/uof1ha2P9mQTEpf7eQJtF95HRUib1fXsHBsbfOhn3fCzLJdPa3anAGXZyOvp7qjtDUh
Sho5s80GgCnFKXRSRlFwujwFh8SQhLWWGZIHD/uWL6sGvoF2qhd6RtORgiSxf/toJFhpw53ZWgxi
SjLn2qXmhXyj16WZjhuKNO+/fskhvPjTpWn4aCf8sXQ0Iahlxub0rSnPTkICWvzM0Bzhls9nd93G
fxtMz78LVYoAPPP5/Y884ABRF4y2/AJATZpXHc2pchwjKQ6/F+WeNYAUFKef8YbZSbAv3PaMTFMg
bYDy330qn5sek8k9X0NVKPEnQsgZOSTQf9CdyivuaN0Q+YHP3hZUDnF20XZDhE09Heucd7o4Z1Sc
kbZtRkr31wvPJNBu8aSq5slpFpJ9lhWCG861IeBeOFVm44rAEA5XxLIayAcVAHP91a2b+BYOPIS5
GNoX9QD2x+2A6WLbS93kPojd/gib3IFPA1RA70+VLCnyFZcGmbMHSEuDXxaFDp+BZWdkpPY8IJ5Y
k60hFIurEGa/Y2mGyZcn2OxoaPGeJwG4s571qhjEZDPp5GhoU0+PwdnuzOfPMrkVhaqWm9TU3B8O
u7iIhMHkUnVDfEorMmvmxtfeKW22SLKyDaqp1JXXq8i1xUnGn17Zy+Lv8+CnLtv7qK1U08JcFSXg
mDh8GbE6j2fwv0i4a1mB6F4abfwjRkR3SBQBX5PyV/R05wyHjGoJUAonQdGwgsZQQL02y+c5QQtJ
lV5bYE0BT/NbxWnRlF9PuSK22IwHEVST5BY5xT38bBnpvz4fyKeaZSGr+3pTeLRgU5WYDZeFk9ei
64SdGpjo243CMmM3l9Hell0sneVY+IXYdavZCde/B/8M0vYbCCmdNUDQErjXDFImbQzD8y6qJhNg
+asQ3j+pwu4QljMjr5Rsc3dnev59iyCLtj/Hkp6IYeKoPXaq4GQTLnUbmlcEKkDarZ89o3ECvQZU
ILiu5WRekmuqhLdafgqC859dahgkV6LnKZsTwHZ4jmA2kw+rGjgx/FR/O0/FkipDTJ/jFcQ9jw3n
0E4D/wcEcgVtNDkHoC0RGrP9JSXcdLwMjEWlMwjZnrtOW5SrStLQON/CK5O5nXIcq5tIxpD+cz74
GTL+BRJ66Y0jjcfFLoo9K9JGBCVscMOcXv2puIC0uxHEhIfXld5HxFchM0Gk6KMMn7tLyMqHnaK+
sSKiCm5vJX0fgm8DIsBPx+54xf8DohnUdk61HEiwjNTPMRpVK1JagZByWAK3ERejkJpwgQI6g5cF
qlsZCbfdCj1LC7LWvjfZntLzeWkSr6458gECa2+oEexeYTGA5c9CvECydspF+TPxHyk1EDTZgqzK
KmDqiU1lizkq1vgsIRHtW0b9E+fSH+0zg6eG+0x5tAFpuYyeWer+ib1Z6fno9lr8yzwMP1tP/ecj
DXrFbz+E5eUgSAWExqhUH7ego3sMxC/kWw55S1WM2Px0cfiUX6hrFHYEF7i3iAWBH9QoZS7ZQoU7
mAy2QXjbbDlM8kJw5yizlxJbWQYXpWeJkgOLDbDQqfOwooHpywneWv/S1TetTVvGAusZJdkL++5U
aUxIn9wfFYkuxOH27f+BcdaOFnvcQz46YZDChu14Q/78r+Qkciz8TuAZDr20YESh7ygqbo5Ezxbt
Ote1LlMF9FsRzb8bSF2D0mFiM4jesk/tJdqDeBRVzIKgGRNHxbzeuPRPysCm70K4oS247esRl7JH
IkmOfIrbqsVFnFafltV7tu6qg8UKxyKVdC46PK/qcpNFsVixVY/rqLzO2/JEtSuZQE7Gm0rTYFSc
tvZ5Utf2i+NwXf2SIHSiMSW4jsiIQeBtcdZ9/J9JCO5klOOdEyDry0ewK+qkmu0Lnpp3ONyAMZro
Szn/Z1QCLWtC3N4w2k6ris0ELEBCA+yfMuaQ+qFyVwAYJMi/ealR09p1lS6dNKEv+JHcnkvlE9oM
yHJl/YG7xM8vJVjjbADasYCY9t5gxWMbrwdwiQHIoh/x5J2IpkjJ5xA6mbYcFgfKNmcF77mnX2X/
QBXpzFBrfUKWhMdW4nHAJEW3EoMaxt36MereOHfdsL+VOShPPV3SK8rzU68IM0FjvG4jopxgnzDG
ZDlPbnm1baLxvcpD92E/gzYla9XKbjOtjK7/wQVV46HDDHW/K7yoWGiwsvcR8Dof7dyTB2UJ5/FI
HIDOHUAfCK/uwf3Fyq2HuflM1WYHd+4L/Vg2nqQ7l0BABQCOq4IMRngivPv1SGuEAYa2CCB+k0EU
oOt8yiGqe+T/kb/ZAtYw8Upv/GKeJzS3aGszHynkuAgY0hmDRR7/IkYRFC8tkRgzGZLg87Zc0QA4
iXKXbLN++UES2SoQws212ZudyZcddmjWj8sVFqTc4lR2eVpCBjT7u1K8qC4p02LTfMP3VXj4U95h
Hlg1VBFvRzJczEqov2bKHJB/G+FQmTgcB9ifVHOKTJHKsmQzg8P1eKguE50t9Psrp+CKN8KV1oVI
lt6ZXpAMTl5XG1eS3Mso+uTsTpWTX4kq2BeBKlnqRwbSWsG7RB0ax1A8z3TXvSY39CYSpDWW0aEb
mqQ0cCbXqndjqrslqGXSb+b1BQy45di2oVScfRisBQdAiSDhLG36FO3hXcBQiEcQsEIil0UD1nmk
mPjpqUx5jnzKkn7GwqoT4sJnsXRu+NrroxRLniDgob2i4qU3f12G9GTvEtWzHu7uX4XhZq6779/f
tCwLqgfz+UQPsWTTfnzIxWFdZdRzfY3ZM57pjs86+5hIDlzZUSPv+msOC/s3rtyrOCaMBDv8saZJ
5t/iwuHKmfecKRaCFi/l6bnfiU7pV0Sg8oD7WsjP4aZzdQFPcqP99Br5ww52IvDHaKLk91EypDnJ
lCx9eLEvzR0FStTFaaitYpeZrSgW+ctZWwb1kz/KLgtd8OgpvQm9wCohYiksdgZOwVrB/LAxKD2T
8cju/0ana35/VxkfUwJAVr8jyjNWEXWI4du18P1/Y4DmmZWlWlIzRXf3A/m7vw6TwQib61Uk2uD5
HSVXpqCKqbQmENCAWxv+M1NxqV7LTuT+pcFg1CiaoU7rt79E0Z+TRfb8uGN4y6ky8nmBS1UOLqb4
3I3Cf7uUwfbL4NBYPnPSqPQdBR3NX9K9xX01k5PtO7W5q1QMDF+i9Sqh3KUh8+0SEdrdwhEm1LLK
lr0LBxqETNox+ltZYyj4BJsug4KrmMROjUzQfv3aFlGB0rWwwLNAeaHMHDxAbK7cGnYiGYQcTcjU
4n+61ujEhBa9lJlUjJTz9T1QE8To9fK8/pk9WIVvnoPTdHNnC0XiHOqWWi44W/yzdv26+Xgbmm5U
Nr+AnU+s5kRDiLp3YBE0+N0Urs3aXtmf30mR+EJ/Z4PSHljZ/QGkLJoGXxLQzLKaYJBbdFIxEgSa
HThGSyeWiNcsXNh89jFtaF6v9kqWm8d3eIN+6AsUet59vThWYrrJLhvBcxz3jU5L4GUzz2M1ZYxn
izFOhwffAj2T99jtWWfp+Bc29yQzVEQuQPB4rdATaA0zuImXLV+FFzVGU8ng7fTQ1YgRbIt1p/mH
Xp/8DU/lAdfcNyYBuktOoiPPteMctUXzVBEUqw1c5jhQRiH+BqAcdcvu5bnOc5QqJEGaulO3On87
hU+lcWYIf0Nm1X3+I1MYZLkBJ7WnK4ga9DBXlzLt0lLdd0AAzT9fN8Egu2w7kKL64fmnIUkWWwJ1
OYbsbhRF5KoD/y5Hsz+ZCW4B9BoyZMVVy1veN4BACPtwyFyhPd+FggaD52cDdV8Pq0I4U4C4+W+T
HvmJCBy6hYa8L9jgNWVRBfRUJEkWiZsB+F91x6e6AikW5ATJte84M1sXnKKM4MnYdYqhx4VKcmVV
F/M15r1JEXCHOE+QQVOYUULe/a0bEQm920JvENEW8vpzrrer4E4ffCZhuS8BODlCcED8OIa/t51W
qyguZYSeWga9Ymy33bxKaYj/sPLBiLFhus+ok0/Oe546J0W9KivR0kTYWLndxoD6EXZlWoOnjpK+
32i7CRbJkP3GAJwnsr8+jpFOUGYNUfggN7apq1ucFOBOCaUqecAYKU9AJh1nE4nyiypOWYK4XZzx
eFNxCcNGic7XOT5lNx3D64l2Svte8JiJRw0ot1cGV8osALFFy56zC9WMScoUaP3OnuQtuQD0mNgY
dXJpGFZFSU8R3gtnQwOCFIMASyorKheh8DGd712e3e1uw+jmP2uwb2HB4plUdM3C/HLqCk30pHNC
bGWQ1v8hTwEWoTo4w8paqtmPELGBC9dumOTImOI5vHuQSgDvum4tlxKZ7iPsA6h8MURoCsA5b0Gz
RzLuHcPew3v7oU2ztYaYxcsP/jzaDj7tfP62imvMWS61JD627zOeArotRlhDpdPhAXCW0foR1zqN
tzqt5HqgZ1LBiGyh6Yqg5CEc5HiBrcvq4LrokHFVOMD1xfHUltWVSzfVpJxKwfzAo6jlvie2lrnm
yxq/dR0EQ0Yzv+bpZBOy3hM9fQE5/sKN7W6GrYMgAv5is2YKOFPONwBthhzn4Jbb5l1xu+15f6Tk
kZYQ3/DoOUJDpL7EzG8ZKtzF1mb8Fsa4SjMYFc2J43uqE1RIdDo2KvaOcQ1hB7KaOxNqVHdExpDz
B4dNRaXcjyUsZbVGH3RTD/fBaon0Z4pUbP4IngaWigAcoVhdhxPQtnbCE6b2VmuNGvr9DIANzkOE
bwaTK0IUr12bHk4btyQNIQY4u0KwU69bJGfaxGfnMnb31IpLFlk7+f/5GYWNXYqDVdfyCbaNvy76
DL/cl5PKxRIZ6slU76TQgcXtp5FxEHF+n5kgxEmp7sWAaOZ8+GiuvM7CdHZbR6iyD/tcUfGAcFO1
nTpbjkLLz8XXwMsq5O0PbetL4N3ylG6ig4C+de7hr6vI0KHPb3bbDJSGZKfWu8s3O/sNGvVvpfuM
yvNkNda51DZego1wHv506wHV94fTNTeuSn6gHmWoAtLz7hX+PNybTarZpUh5CrS5z65KNV5lyLq3
Vzhap/jR3ydzVHqH8Ascm8ZYGmeUkGxHIRssC8KQ4NQyjzCbB8ukwl46uf1TTv6DJIp3M72bmJ4l
WWHwnV06W+AGWAEpYfn3GeuuKHmY9EqJthAOBwl1MglTn/Bj+b/vz/WD3kLqPsuXj4m54TEvdA+r
l9+Bxr/kbA/JiIttM06uQ0Nfm0mOSZ4RBi2+BYYgY9zsLeWZPMArl/a8/exa89q8QMi5ZJOQE5kN
HzkOb1EI+lYTOsYS9PIvUbYhPmiunNdYKlaFWD3rPAY4XB5Jy3TUILdIBt773Sg7s9hREd3L8N/X
DPU+KnpuCftzijrwYi5AeIAQeE5YbEVzuO4nIzjcp7SL65oOMqVUhE8xVK939Ls1PoQ6Gp9PA5xG
l4umLSeMPZtSMReEqOOK02uDGI1/MuC9LvQR7bIWHyMzfMhhdwXdnu16RXA87f/BoROfMpg3nkof
KTs6AgNGEsKVBhsod5oHoAlb0SeEOMrla3qOK00Cn7FLAPLZaehapwbRqdj30GBEceH+hYbyUa1/
7pe6C7eQIITXYRfDl78Tw0wDh9ciyT9/xByjTZfz92LI2Us6xrmTEyQtuzlhJg1sqtJAwZX6/gw5
X9mmsPOnz1yhud9GqRLiE1KZpJzzum3anbFlEzot6FJAVbA64WZ1uZ4MjLABPSyTtxQdy7BQ03OH
qqfmGoSydzYPVmIJ+vUtPnQlRFJYnZJ8HCd9zSn29iiJEEvlox5UYU9mJ/Ptsmcj8+L2zJnacUia
7N4w3gVfQJzcdaH/68fUovzUllofGGu+eWas8RNzye0y/PlkTmJ+9Kv3aOlAAZOxMKrT3H/5dTzw
giLnARfgvHLCOU8xCheZFIAtlLFmBpY3wwh8xtIL62iid5uSO+bGcYf0wS4YcpSoU4E0jneOLmZS
gvHIFcVfbpw3oUUmK+spaiOK6zA1/UgfKSJ+iUlhmXsWplxe3BIa79qIEBmTBcCL23+4cOpZ/yG3
ETjBR0+/QsahgcLLCoirQPoHKEuam78pYVaOWYl8AKbxxyiAa6DY+SPvGFAJ1Mwt1CLL2etuyBQx
sWGDbVFqL/QxI+WX7/Y4RHugN3XY0YzBQcS4f8hNlwIvcTth8ctTMAL6VmW9Ti51fHnOvUHOFAWT
RaRkN9Zy7IvSPXCe5xGnpQ2bdHDK31pkYfBb7FHxBuwaBnnD+VES3qC84MNMqZmkxM6ysWL6pAv+
wIv9fd5gdUGDnCa3GCfWLhr676YydKEm5PLRNjYqlDQ5rR93WGWtdTYfYJeFIRM0XhROrEJ3oVjj
OAMiS/0Wl7vJR5ypbVL2S3qJrAyPxOLwXpZuIG39/Wf26CDpGiqBf8lBu/0nvd41kbWmerCvwtOU
0X6Jh+fAO68jHQWFM0qjPDj4SzNL1Cxz0wUH9fe+SK5IdF8lCihXgXo6OY5D60ewLLUYUDx2IV4X
4rAek9hUvl5FeTBkk6iz+8JT4CwUy1ylQkku7lm1e5mmn0rVWQHtEWmwxbpRjt9OY8UDgcQ91ILk
VXUPc+JbXehYvVi7/1MF7gv1Id0md4TBN/DLTa6SzDAKENZHtQHBcorjLPa76QLL6XobL4eJ87Vv
EBJM6Yo/PhAN/+2Qy8MY8zxmCgw3Bycl/U5774d7W1mTJIxl4zJrA/Ez2LGNtGrFWdhN5J1WWIWc
hTmixZPnrDnjxTSSBuyYwQOwkylOJdD4EnXqFzn/hkDz5zsaDZM5OC5A79WsxwjhnsjOZs0S8WEO
4pvST/dvl9a3AtAhXhTB9TK121qJBlF/rNu0JYe5/KdfEmM9PvYGh6igecnwCwHzu75sjFVDgcRk
e9MhtecYBmuGZFmfsBgA9tHgNESmXt/iCvrWhnqtgRSHfwUCyflN11hxOxSC7PCANfVrlpGyGz30
qyZVqknw+98E1Xy76nEKts+XxQ9lBsVgb95Xij3q7b1mduu7Tf+R9U9Jje5JK+L6qw6nlCDUsYn2
q6Wpyprstrt/HISU63qxtA6rFEZoOT4J2HSIARp1un+bXcYtFirxZGGI8yGE/xqNOFcxaKfHlvhW
dMyfeQJxfYOcSflmr8F20efaAExH/J6NFmSDAV0SqOyA1Wprpso4Ae74eollbkykT8jjZoWWGYpZ
vr6kdc9CA0tvsTDSbyTodnf6dlfEOT7vfWE59DEuB1EXrio2HWaeBYyOMJfr8g5h1C+53TnYNrmv
dTAsdXQHttCVGewdwLsxemys3YMUyHAi8ZKpNplFh3Sg+AVz19nGC5g3IPUXNumjAxEMTXmSyteH
EBFMaKLlu8xEqZBrFTDNzOhmDjDjWfuB6ZoyoQ8j6dgnXp9RrGKZg1nM1C6GcoFVohSVC5paeQ48
siTzpYb9H5pdQaeJjUBcLDATJB/zNtbX/UQDwUPWyOaKxA+75yS9+pKGr+9JDXpFnhqzczibhSh6
mv7U27+3tRe3qESHjnFpSwDxqdMJNzmh/dwe+ARfKBtwDogMxE5ro4GJMlRJUxuLWP+sP9Owk4MH
Q0vnqp4YjvfZCPmRGYne76zqxXB7Bzbyt6qBgBv0s/CO23T8k/hOLnsh1f1E3e4Bq7619s8Abqzf
r5tHpjd5/zztqgIj5KbcKrZ021pcHnT/24Dis2ePbGp2SwS7wHwuVnxt/7Gn8RL+hjsf2g+zFR+B
Xa1YxT5hI0p7N3lYaYBti/CYr7aftdcPVcu1SaLxl2i7B9zPzKeX7ZjWpmRtid8WLkZpg2U07uQT
tsBQ9GrttbFG3Rt82m8PE16CrRRmmIuaFwwNlMApIHmFRY2Q/eUQKSjLBATSdOzke9akR9saPFsK
g/9KiZ1hp5mHctFpNhWSavXYmZFfg9SQutCsZpD0y1Cir6XPqLfCn+8rbrR9RH95lh1bsl8J28rw
0AT1GpiLykwoFBWqjq1rTDKQKzLodPOQguULIVc1R2uLzB+pPBPmH78Hg/GHNzWE6imzjU/VLlxf
uDOxDY74F3bcVfrztP4mFWoZwvqKjqa2b2a9LKB6DXdJiJtG7/vND0In4DZjwS4Kjm0vTrvXGkzU
uzMdHpIWF2VHYXXzTfUQ/5PtuPKS+ih9kxB3JhvOPh8du+8UrUWVz+qLYzciRStnKLRUR1rD/mB6
QV8Zilf2+jEhiyffSUNDJBq5DD8HlRKbNJdHRZ2xDvmE+Zw74CvFKdqWVC/pyc/zifuX8EVvg/zZ
uPZd2K7xfzrs/vuYFr07SXQlWTQuRGOsldEJxVnMZiJq3vi7LXdMBf72XDsBuAfQ7fb+iKBXCQi8
MmHPRWCubfGEeCkYEzndpQYrYjiXUcSjyAnPfazlcTwWMzA7Ds8P7XCIl10hmLox5GjKP2i7r7JM
DHPtNUmFl+B9AnmsBF3wt/rrSAXEoDqHGH3haBFn236FvYcHPhFGI4ReqiZAUaUBbc5q4teh+ida
uPrJfVe/ifW1V3PezHUSVxKwoYbpQswu+MaSQ2j8k/WM8P4wzyoTRKTctRzp9QLAGs15u5fGIP/y
UnJxoDiPQBAT7pBkK85hq+SRd93LMMzVNBZudXlXmLgmlTb4WA6V/bvTOtnBsNwcU/WZMBR9/fOr
7lKCgnbCiFB78j0Dnz92Di8zNftZeseEHPEz9icgrVfY3+sC7GI3l+dFqVas7Bf3FljNfTPOHY3X
WR/aZrdTfk01VKzVtQ0KClyLbJj16GYR75cgdfGJrZFBTSLJdMEbXwj4w3bhsW3m6r0A6UcdPE3A
HLQUKPbHUr8dp0ORg4+M32E8xG+cOmJWLuK4+fshd+GxUHh46st6E/ComH09OZMRO4hAO1y0B1Hn
U+AaXtN/qHHobiPSmN9FjMcauRrLy6CaV7ff+6Q/w0l5GYmq5UITU74jlePZXwtP4r3Ca5JCOm4A
QtrlrWoZptVjI/mr2opHQ7NB0HY+VGq5mBQoHUJNWs/967jZvca4Oq0qvhHAm54G9gUwMjKXKsPr
Fy3AwZNkr9GHOdb2p+3N5Wl/Oaa9mHm4+BLo+tQGihEJ7yNNWitqL3J5hL68oPoKLbqEP9WGaEjn
TndDWU2dNfXeFaRujDZSGvVqVA3S9s1pom/py6eaKilSAegsKHPQy33OWT35+7yWJyt57UNIcrJT
xBFnTc7uh0F1eQ9OuHVUNxYMzBEvxyNc1B57xLDtw/Lr16y6invIa278CyBB6CGt0lFDp4ZZ+Byl
XX6SOvo5FsUospqn2e6gcnOF7dpvvYU9pjIvKh0Cm/1GksbIHM/7gWcI9mlBUxoJtDT7oXNJzOdY
XiHs/73fJUO2Rz6lfpRnmILgtKPMLGqCI7scMIqR6PmlV6yQPpuldvFYZsOJBs9sbAwO8wI8yR/Q
ds7yL4f4J1C3zo2Lr/GNR4dB8i+xSPRLpvWQ99gRFcPkeJzITiGlhxkeqmzYaF3MyLrPbjdrSZet
sV+RAVR0mhfgVK16cj7iBwyPPs4K968A8+/IWq6YqxcBDV5k9I+BJO2FAPLjyzjcgBnoxTlOTHqH
Wyf0VqtoITwLCwQui2yXyMVjXzPvK93f9RnuMmj0CxmnWypedn6rbifj5zjoGKV3TZcRscGumQSg
85Z8K/beWbk1Ts1oEyP9qP63ZnyGsJ+Ic0g/UeH4XuNJ8Im7aGC7NPZHz7J8g75r2ZOi4sjfahme
Bi8wVSNf/zVh41D/xAsf27ioCCeSkApKmUjFZd3R4ZRIs+RN0Kpc/FmbwO22DdPsp7TiV6JDQakP
GLorHDWSa+DcEj7OZiM/2fm2t2jcPBjjAWrWgGmFIZEXmP84c6cixOSemsBDhXj7AZXWC+gMAH57
jirCU0fpSZRzkU8bTSw5T3A+HFTSLsFU+M+a/BOCnFvF/zZqz9r09fEQbrciQK06CwAPCKZ4N0tZ
DCF/fBHZNDx/LuBc8VRDkovEFXRaliFgMJXDha0PEqREHVVp8DonokkYdG2XWMIjJae6q1BfPe5A
4onp9cV1h4mflXPfeiAs5oCRiKBQSMEpRytJs/Wt18mHjobC+Elv4RNljZ9I/Ewydqv3Bxx/72P/
JPDuBKatYBoRV9VtGej/Cpo6Fg0Lj+XpZ2aXq/jQ5lfCUufUFTJE1c4UZHlCgQoMphlnrLWxHe/p
6t4XkINrWEa46VBJD9o+0ObYpzHCesGtTW0c+qxgVSn8zC888VsZZjYgjEf9R/u/mLK6IzsKfMrK
yu9o0mKMnozIKUYC6wcenQKi/lz6CppgBKBSTWE1ZB7OGW7yybvNQb7lwnGPcSbUGXGcviV/czjw
UJ2rNSoKBCgOz1EXKBcXncTbFeHFtuxKRMXgr5mR7A8tBGDs25js+KIZbtmw0Km/HL+9jcmA9aaj
p+WRml8DI2XCQkW/Zvl6Z3bzmY6VwwlssHaFLVbLaUT3rQOZSYJd0elgNj9l9ohDxdOB0Icq4uN4
2FlzwWT7mRawXR+FKkDLLIy/QEi2ILKnfEiPsJGoXN4j8X2cHZRGYEHO8vi0O9UZVHV0StD7KkdG
iPKwKwEEaPJpjImdn+4xvOKBnXTfOtvc1jfprxjLyBX8jS+UkSuFpfdsxzoMZ5PEqdcUiaE6tssK
E40nbyKiR2bfpW0McxWLJOl6H/Vk+Gcwe9TFyy962lBkxB1OI/d8sLPTkgk2bYpi1YtJ3S392+kg
A5dFRV6wU0Xa+JJfRd1P3UWrAh/yfJCVE6AGY9DxWarMIeQDRxdvSgOAE9sjW68rPbn1PSJ0ofIv
AAOvEJ3olzBy5MzEBSHmzdrmWljf5eopriV8RNYaFmtmMm816QaZP6iWG26MpeTohLk34o6qULWO
VVDr5o/QH2NCyRrzv8vD6pNcGAoqhkcpTVW6NBuxN48IwWG19r4Bk4d+0dE6Wu6NAECQP5JZpxZ9
cJoJ2I/ByhVOgRVUhZWZ3Uihm+MGEz0bAr74tdVNgx5dEyY+XdPHl6s7yoSE2HKYetsb1uYAwfGU
d6ro6pSJTTl7LlOUZBWCtFHMuhWy2gErvl4frAZ0CUJ3q0ppP9oTUPDmp/JOyS0LU4m6JkmoN/zO
v1oM0E6qJhP9MqC6+f/+q75M3maplrbFLwaWCyYALk7igcCciQF+tArnI7uijvMzNlxPhdofsaNN
+TZkfy/ekGZw+CMkudFagWO4IFv1GtCHCpsG+HN4myrRnWlGjGuIqcHf8Ii8d9KXaLoMk5vX1zy6
i1dj3HkGuqK0YeEVrRo+Q279ksk71LJ6OFRJLEHElQUIReFRb+WO3DsFHEiAqPB54hqgvTtEDBGB
79r2EBorWaOVnfLEiDtPEmJopJ3m91OcbVkrkE6BHt7HF9NqMdcwpke3mz/+VbQ1z7Ls8sP9WdSn
LLNzPAcFlYZrDlDU31P8csDsFd4UGeDf1T50MyzldzjC/Wxv5kJ2cjoT8dQwgCOCigQPQNAPZphJ
s+8+Lt9F+u3JstwBpLbS6xxC6m49bpB5+d5+c+wMerrVJUdZ02rw+aikOCPGXVcWZngVva2G/2zD
FFFTeqC3cjAcIIxsVE0fr64MhJyfdXl+bvXSt3335NRmiaOncy/JualgGH2AV2JJ2i+Mvf8RKdJK
VO+WL0wCwrS04St3UtjBxIEnoLTk8VF5owl+adSBUzU6cM+XMyMV/FfOkWY//k2pBjiZoaGOwGZE
OaP1+JXxXi8d3JGixIN4XLTvyvC/xEzgntev/qlpuTp+DNpCnWWNeWwQAvdgnAvsjpz1/mFPJHs5
HN+xIyTEhGri3kFs+D37Xxja31lNnjSGxuq1M+z6XWLHj+I8oWhE1t1uusV8+eAnTjoSh6G/dCa1
sIkxnUb2LRdZ7AdlFMjkAEeGbTY+YP7Jc0bzXzwP29zI+Dws856gqBxnCEdnEoZbNIiSATfwF0jo
uAW1c2GTfS6BDAy4IovUV3l2zu9EyieD+Ve7idZKooJfc7xy4O9gU5vQeEVRpZlj+pAqdogKioUQ
i8HyM9kqakaNQPkCw/ZJje/sTcKnNrn9Clvc8m0h3Q+RF0GJnEj17LxuSVighVIrmL8dx6jsr4/7
VE++/D/7qy+iAaH/iIdbqyRHWVUb3cbZRpQoH25I2CMcrFG6zwwZyM00bXx3k1GR4GDkLKVQvQdH
hqxCNYRs1wPnOQuw79q9UL4sYL7owCjInJG+eRkQdn2LfEhjeppJHTzN/k+nua968TevRm8wS8Yu
wUkEhIPPKd/uaI9bbivs1JCPjwLe71i7GbDG8GAB/3Y1Pn8bti2nztEccwC3EGdFXw+s7e8uA0iI
a+KjARxphlH6fhNBq4cyG3gmG1YaCNcYceFVkzB0YBEhPuNVpWo/sVCJ5i/ZKxtvJ7C9nnBJuvrS
hMJzl++csx6pjlzp6TQtyqM8MEd1pZl94YiQG89A4toK9kukR8FKwOObtHLyKvomExJMF7AbxWXa
e6m/S9R1Amq/9EsJE8eyGA2IZlhWaTg4s2f2a58o1+bA2t0GnWdHn73kBatwJE3ELEwVQVAFdvJC
Elg1hIuugaRuWqOZJg5M29g1n06cTqqbwuYooJU/YPPHrHeV2ShEGqhNOWxUM90dl+yiFNHrpQbB
3oxHDNbntpatuzH9jYw8q7J0OJyXB6TeMYWq0qMjSvmalB5+MHCAbMjSf07nF91FnUkGnmuQY+89
U/k9iGbKZqi5RnPJaPavanaaEkqgD+RR3lndouUlE0eKgCKa1BNk1WIC9x136HRbvfs+HFcx7ry2
lKcO4SDizQJ24MARJfvke15F50z5l4QFkCYWl2gqMw+Fou4IRd1sAgZl7qGQiCwEw5bPcmOmPHDa
aZZqHYtFlrxDwV3hnKZwdGsuvga/M1rptABgnYJaK2Ag++AkfaqldwgHVISPssqUl1uTmsmBDh1Q
ohK0V0SPkSwnbRrwL5GGrzCGB4d8wUCSuW4w2BhiIXEU5vxqq3ZIVFPDQpq8blU/uEKamuRXwS4k
OZlXb+NxvNpqItCOSUXVEwR1P4MWh4cVytUmwhMSMCGMdMarABx32Qdr31Jxk2ViuWLRLEAaXMrV
lB4L3SCpJnyLz6a7BFN6B3K8yNQJBbC1Lg54yCzKSKBimOz4qpChtVlikVPslnAH7bPpFJ1D7rnY
yqSJwP03aPCg03MPtxpjj1Er/rbPcxk4SgZR9JRwJ4SBCclEYNqVFkGhVrsIza44d12+qU9p/W6g
pr96WK9y3OLHxpk1n1yPTVbfbObE1JdZB5+jAxlG8QDo9EFLKvxALdTub9ENjn2ivfP6UY2+J4vd
QbA+ZTlUu5ULu+B3QlI/mWmEBjWF60EMs3Dfd4qPcmWjmG5Ux5wDl0Q2d3t2tjJEAs8N07Xws0ix
mARPxS3uuOirMuyLaDAFggxbdYqf7MYrj7NYBJ92GTqAkEtRoeOeFYXFbwITDdYzcYFSdxDz6n7R
9pPSQ5pTa1qf+fC0J53Li8LbIJKi35+bPRQcJ9Pum1ePotkRx8RySkf0JmYxm022edj6TAER8T4b
IWkFRilqMVf5InIJU6O8d25/nDIcCF5e8saqxE1+uyMWl7yiIArWBplG5sQ+MsYFBz8hIbPtzRKt
tcUyRYzjiFVXZgwka22BtNh3AJcvgEJvJ3mEWYVun0ujn3QMPuZWDKdTzlM+u96K8DHWLEh0+ajn
aP5DXhpHR8XiRMJ8EfO3Yj9Aoiad7QqnUlpBikfv102mHETC5eGM2/2V2Iih9qaJKhu1A7izemqX
QBXBXVhhxWSST2HxAgiE3c5MqLOcQmBOWvTbErAxLfTt2MJ/VTzFS2LQHn8tmoH6od0T/qleU4+Z
zFOyt7Fq+CrFjGcd8L03pB01gv1m7X2UAs9fXaUM030hjsGqKSywlxPOR+nsm2IOhWULO61NWOs5
3RMtl+e9uLQgBtMASJesEor4OI3DIWcQLpe1MhUbYrDZzNC5Gf+M4iwUHh0AcEBj0cC+qbjm5CFM
Ov5eQx41Dlwj0qgWJsKwv4C8tjYCy88AMoeVUWrmphxbld/LmBHJBNwUwwe9rGAsji5tIugJ4oAe
CQhYUsPFaAJMD7KXccugxMDJOrs5yQGuy10R97IF7vjU15tp1N4uuk7LblZnFP3/IWEMBpGvCIlg
u4ohmShOxnhN6wC5cjN9hnWMM8N6VrXIrCxrrxUy8rl7dGsY6Jrye27G5X0rg3AKc6vrr+8T3GUq
Y81ca3BFOarEeK/LdKXyJ0l+arIFuJ1kozMxalPiS+qlGVH2pV9EfJJ8OI6sJZtXEQpylHOJaQz2
ZisUIXzj+SvmFbiUH2PfZazKjPIvgExWPg/F4Rk2/LK7guAKpNi94KbVdf9SO8OrzbqnK3+mVdgh
mRSrh1fivsTZEmeljnb5pwduKNQ+j611NS20AnASDAWSS9hB6nFTW6OREvV2it3bkxIUwoauqb2R
USyVHEx0Gb2JnO9E4TsNEs7SsJsRSgxqs6YxY15XLia6YLKaMTuvdGz8xip1pC/yYYzsW29Bh+E1
4lPBKh+9l37CsumSW7bVpe+PRRNfcFN1bvUHx34zsYI7hiW5z/IWLEPoj4DMYovZUzyVVzqVcLrR
KJFcXi4jpU3be506chz0TuPeEy4RDB/pDyKFe7YnJokdp9HnA2uDLk5hW8B26+lEZcXXuNFIibSm
5gs+gtlQQ2jL9vpHBunLxPRzWRhk+rBIMe8Pbh8Ti5W/QM+GTVL5pjXLQ8e5qJg/6mQV6/SAkEPe
Ub23FsjcKLRdkf7vxLQBGhHrtTpAViAVvk2wHNPjTgyhP6HWxYvPHEyBxskjj8lC2eSTFoks7pqf
iEcyjG5Dk6TCo/87WOzBB5nrCLMAIWISbQwIP/2aJki5iPTdRxL06+UgpMc/piDZq4PmhGCA609r
LHVABz3xp1ZNWoJ8tDA/N+n44QID4KB/t7x7Iqxilf0UJ63z9kwp//F5s64Nbmez9q4QeF+dVL0s
N0/no5gCp5t9JVMseNueVaL1+FagXlOtn0bjmtf3Elj0RGRIn+5XsB+XCYL71Y9Mp/FKv2FvYkZN
PgzHINkMCGvOoPlPkwQhc/vE8h0iaElMNcHk767R+PqXaE/ETN0w2krPUfumXSlp4iKO9hV46Xst
7OlEG5fD6CfhHrYJavZUIjgqhyoPmoAlxHlotW6mj0I18qDfN0mFwQkw2q0RBwCp1DDWnnL1CBvm
BTZ2a1j7fSRLHAjfHzxb9AT2bYDGr5id+EODhymydbI0W+K5xDk5m+qFG/qb6O0eKKW7FkGK8Yyw
u3pobedp1zYOI2TI/zXg/Sg97dftjReUypROWKqXx7wrouxPC8ZhPNEatjf6iIpm4AKZb2XMG2Rf
TaFr5yB7D1Ki2GjBVoWtNQ4Y5mkyiHJk1TBPfBShOhLyTS2EH4iOOHDAmWM2yikZJaSfAKdsoEDk
IsZPpp99NE7znsYxB9MygwgsozcblgTJOMATkDWtXGmLJ3x9B3beGXAGSHRAKpTSuI4RBCSf+MB9
9uKyGxUVPYfPeabkVl9P9nfFLJ7Ny5rP0RazD45f1mIeV34vOi2C9w6oRZ6ed2MJXBpRoiAd4WRl
PwcFU/p3JpMvqz/VAVWJ451aWi413F+pMUCYC231M9Kll1zk9mzw5C5Toi57o2cz64Y1Qsye2z52
YEyQSb5d7yz+LDDuCSyvaFdRDVbyvdOkuQArf6NNPspOLhVIBWAsh2XnK9LsHbePr2xfI6JG7sLi
lLP6FyB5YDlgYdKE+WleStwHyj/V1BnDJC+V+1No6jBkdHOoDb9LXJoYRXgSo+2UnKOfcwSHHz6g
yn43IUoq/PXE4tk/xPbwVhYP0r0GmZ94GhagL6X3GeZmgWajCz33rtroONeOEHef1pVLQk6TY6Oc
N/S6PUPwrkLZIFTinWIoDy0uHUkI20YTiNIoq9qqHyrHqh+QQ5M/WBMyMikCbKSuKbsqok+UwfTm
B7ilJ8O7Yt/eGOio+fCDBBv4eSsqlrcKeCUbL0qPFCfzI+56M+uTf4ouc/W35vK2bdSCc8J5a3GY
mBmKhp7yUX80+F0ViXMfbQYCnx3phala55WxKVrEQrAGoqs3CacrOQl23q24n0/B6qa6F2ZhPdVS
l3QNQrqEcYLL7SzxA5le03yGX9S+V0H+0oiS4JFzxb/QL8nS/bVc5lmI7k9chEAuT8QMylggdBgO
x9pqBH+Zf3mddrenVRCYCLL3fRCPXVkQB3CqynbdQHVt70wbLnZniokfoQU0Eh8GDAXYwdVpChJ7
gWx6GLsL56zGNm5/J2AqLnZehIBw46cA9z07hH17+LS5Rh0wJ67mnca6FFjjxU9FhSgU48PCnSoa
DmFPfzsZZHM17fb9q8hQ0FOgPSq8OOj/2GPJcHikCMH3wpTeDeWSBUWiKKVX7FFek8pGHTkXGiDj
XLtmz39SRyTRy5Ao8higefF6RpMF9Rqhpsj043D6Yux+WsvSZkdjlIYaFHL6tx28hno8c46HEnbW
yqCOi2RB3bxTpC240KrYX4CyhJtiAvh83UkbpDzCAeFvWSCek6gvIOWQlenOsuHK4iy9SchTeIfb
2k7nV8XzsGSvcKobBV9Wuu3xfVg3BmJ73ZlkHd1MVyBbWH7x0xR1ugwpcCiFmXcVjCNnho6oFSf/
75ChdsjilSsJZE0+3IGoV1Eh9v4BdSd5NatGVELtOEYtzNjU/Ccaz69eElJMC5FmdjHBP0Iz5Iut
veOlOMZAMpPHL3k00DPSvhjhMX6lZ9czkQ7GSICb6kgA2KsLnz+ellGt0Nw+ZRVBFTSS6qBCQS4Y
9VekZErTrwzEYuplPzQlmcf1EBXICQN/5NrlL9yHWRIfhrYbCSKockbYgPV5/GC3hREgIAJTaa7T
1UCRObqTCeXDc7Fto+jIdC2SL9FbpGQGABdAKdNmvhBdWg0jVN3YjHi2ZrOGzUh+Tcd1+ka01/ri
7a/iv038YrUEc2pWCPrDs/2uMxi9SSl/07Ty79evencqJQfMENGJQHFNl7HaqLr/w1e928EXh2gV
tWL4lO8F9RSgK7jKhiV1AONPDk4Z4Koiv1mWqSV1Bh5B1cZ2MT+UOV7vrMyN7BfflfriTl4pfJhS
gn6jbsCqGNyhM4sAIKhUWoyuqmzHO0ovPkAiwshD7RQIzrlNSVdh/uD8/9ST+b4OF9HYOvonq2Bf
s9C3YCTXoVKPWWHE3L6pnz0UwUmukLooJNd/NTN2L9AOBqAMbglMVhv4gO1RJ+/7wio3LXwdzGoB
tK4977NJr2A3AqvUwJOQwEfddOyxL5PJClxWgzgJ/N+zvCQSaltFK9grht/bFAKJaj7WOIh3FOnT
HGkaczX99wJ2snQusv28VbUxF0b3nM2fnbiO+BawNnvz6/MLOucwIlJDxbg++4k1JwGC7Vo9VIwj
yXgmU1Sg+PBksLpW46quWuLBXuHobAPtpGw0a5ipKeavUmitfLF01/ZtSn8vDDPgISswRqcmHPeX
Vvr7c1OCiTJ27YUlGqpP2e6J1dconI/Dphd/HeFUFHalK/OoSSZpryTekouyGKU4ZDghIJoMoHaq
CqXvf7FrtbZQZGFtdNLKDoexTBOP2pPWjveW0YS5j/2rW+hx/ReKNp7t+A+mw970E4nso+1lX8Uy
wT7eCadIznKApqELmf+0gH1N6UCMybJ6eHs80VL08rHQbUTjM2JBsHjowekzMD28BpO9BVdKKepM
oTuB3c9ltX7ycMbLSO0dkrjCy8XPIFTM6gD/DAeB96kj/Co/xNWPkx3f38pG/Pm5AbGQGjifpp9Y
w2JRA1yVGmP/hhdWn50PB8zhHd3fXEGGwujXIg4f+n3JQ0ARhX5B/Wg+5QSutvELbjt3dL91fpRd
bVhJEjgxCX/QBGAaIX4DdtmCwNytQTu+JSdv9ClZSBW9PsSBEofbd5mVTGpN5qKF2F/ZbVI/5OmF
hVexb+OSbwaEUdSzXRy8/3Ic8sIThFk41a1LueSLoJ2BoGxdLp/9vA2vbBvyyKn1uNELSmK56xOC
pTwUhPAQ7a1Br4cPavefAawjiMXxezSNjJ8sGUYhuFidzR67J6MEOob/fXsW1eOFXZWqXnMHIPgJ
a2PGbpuN1eNNf9rP76QzJxfEl3PP1kYrrQJAKRY0qrVzaXTThuZriXmqGHZdIcWJsFg+uXAgqQhy
+xa05zvU4DG6dUCmKVYyne7OhXfZoHBm/fSnkovDVfkOeXXf4QJgn08fZl7/6uW6AyqU/GVoHBv2
grMlXRds69ZtBK+FAACbCbZlMYiRUl662jQGZT9tNiSmfQ0BquvikadmTEiOkTe7g6EjjUxpedLb
J89ADAHDzkbHNZeq2Z2SxyX7gWlgbCIOqxKdcLgW3zfFMh8UJDWEEITirXpp564Z4gYfUqIVmrpG
xd6psGr5yH3trHI5+lCK8GU6FQ7dmTh9wbFFeEqUOZ7QhCKSFPAHy2NGbmwSQMwUTyeGl/vybmRx
8I//N1SCtUzkgi45qwsV7zOjfbJy+yZp227EpzR8KQ26wvz3keeuBFbioV4pmlfc1yQVlBixySX9
YJYooNoP0ln+n5bf7dwFahxygPvKd1Aeh3LCeDN3iAfOG/QIQksP7YNr03lbhzBkiwwm8xKIDwOM
VlaTy4DahXSOBK70xROOZr7KnbC5MiLMb4HENlsIQvyyT/OuYJwBiOR8bFqBy2sY6jvjCaejgAdO
YnYHjOMxFfTqHiDpc5ThAFJtoqy72blYLJsbZeMwPspulAkAXPqq68xWjffnP7OO4vh3nm05bMSb
LIbxr/VXLNP64nBWvdbOsHaUIJ1ZvoksU05TvEuNLxaVy6k5fdPaQsrUYhN2TkErCPPqJm7q+Mw4
zP87ilJCNfpsemwYMTU43obcC1eLSxPvm4OHuWw28AlkgIugxXz1/2a8rCr9j6bOdoarH8+1CMVc
zmHyEBqUAT00ZByUdi5HLwviHoRASUq3yMoRf4gKj69xs3SuivsxEc4UHAaotJYJWRPRQONMGMsy
rWEH0sJ6n05nslsgkuLVjZNPKeLxqinYrgWrMHtFzHzSvwqAWqxzXg6Uobdai1HCMWVVTh4Fh016
CmDqk8jO+O4lLX61aF5eW8CIsX3pRiYYs0togEwv5VSQriVgT4jFNFPkd4AVr8JZQ8GHX7jqS1sb
SKJDtw1ouenu5MJmTvX8CBqljBY4iSg1PmvuryUK5zqrBroWCBm2oShbzkYudUsj6J0HdgD8jRQx
AfMB+pamkFI4ryUjWgFY8rlhvtmwosv2sa5Rus2HPHwjO1MiJLGHqkh/FL1KIOMPbGkFDdNJ+ta0
32n8khBqV9Ljp38aC42UOE3cuEA8T6ddPpcEHVXVpdYkb01rukZT+cie2BOCZRfNSslpBZ/FDFCV
AEvuQdaOt6GrmnHiFfruBRod1ixJ9Om+kuCuM2LC8539ggvf0VuJAQJVCkibFh7on5QibJ19+KBL
t+mKAtZu54VrzkhkflMH6RI+XwQckJDCW9DDOJHIMLoKo9GnG5ivmleXDdkAMq1Y1RXV7LA+ZrwK
YEdmDT4XJqiW6vYxRIV/nelJIplQA8mSW8u1y0nfBxs+PJ4A+DhjzxtO+0+EjkKgzOzD//LztUIw
aUjn5cI4lgVHn93FBJx8e+Xbj6GgNKGgGZTgN0IFO9PYBJ+S1/HWEJKtmujlTH7ceMd08BJpBQhC
XG0q3GJnhlszl6HcHQnsonxe9painC+SgLZtS94gl/2g7MtErG6goyFmYFZRoGELgoT6NB997ErV
bSvH4/Dx1bcYYpGqakAGhtSFums+P8kEY0Giw3/6prv3ZovYTdeVg+wp14iX6IoMIxLKnZHVhWrL
AG22I/u4wiLNwvQT+MwyCZZIR1N2bl6UhQe7JhAR0iXiX6XldMoVGPc2it9V88KXtH+BLrlTMq4g
tEUPctOsU8Atun8o3mnn3MdTFufRKp2Pe2qUmzvvUzxMjUS1pv9N4PSt77bEqp/AoOdRO77nKrZB
qHZeKJ7l2zo1zTQ0dLpZS9Vd6GhIJZciXTzKWaYqDN8xeAbJfptoGf0oZOkH08bHXSYp/c7iiyKb
Uvinvfspml07dx//Ws+/mAesDKbVtvVB5iwArKQ2mGCFcRHxv1VPrMuqVr0+dkqPGS+Yg28nyn6y
vvCeBgTH+SujCtU5/TimmePv1YH7h3p3L6pzlp/8iBq9N+0lwuvDBKyPRNXEqhNyIbnEZv6Nx5iI
y+HZ9qq3weQVWqBNiqy7zBMzd34vCr2EmDtKvutQQol5vAiIgurwzTNpRNx3NhOQ7uPmJjEmfiqQ
oHENuNayC4/y+jq4o+FemQgx7JkedoWuv0Mul8x3NyihGx+UyAYL2XstCJ9c1MmAF8a5AKQVc/hT
552iTIERDZcrHfyqZojT1yK8nqcKyiqlvk34e8OoRh9aAEFDx4cPbZF7hDKXUomx9drYzz1nqEQj
1YEXmMBINZgL8vlLEGHnoQw7eA3Td/VPCJdoCoq5PjEkBLIhD3W6BpBm1Q627z5VkTHZq9kuIMKh
cBLe68YqwJsPi8VrfhsD/LjDG+PM2aE/3jWUAyD93O7a5eYB5c1+mX+Rtwj4XNQPDrkuiX2mOhHS
qAkfQhFZnwo8A36Jh/qPuOh53FbnUAfQrwcu6x5OeLfKpHhfqtXs4wghTwzjR+wtRtyQxOwgahvj
PZWNp1/C7SbH5ZVUvCI/HHi+Yghw9FbdgMGtVrATWTUmQcUV+69mSWmS4DtTH9RU+fP0LIV7T/Jw
3lJ3HKZ/sQxgazAlXBoLORC6O+xRdN0mVpLBv9sZ6WItdGaS5sjr/yCec9HyL3i4cehVqb9x7WpX
/79HVRCS3oBhsmdII8biIwhi3vXEs/1gjn74jgI+u4nr91xTT/3kxK2/fDCXmYKhq9sA3knJCDI+
D9wXK/VenuJowKQeoyR1mDircODGEjwF/WU008xWQgYroDd7kuBbkOpdQBRJdsB2SpXnbRK2YKg+
lth949EubJOhSqOcYrcIf9Fv+EgbVxzcp/RHsjnBxv1AasV9D2+/0wPlb6HSQokCOpX8v4lmUjlQ
rl0cAb4NiReIZ5k6YtoLDTPnE2FeTEkqNPrBfq4x7wHX23h7SuLJ4C/Qmz7oe6P9ehvzx3VB/ee8
VYEGSjeogAVzkl4NjcPqGNsgNZo/zN+Gr3hZgpZclrKN8bxuNSBVRtGfyixgS/9pMUIvx9iES3qo
SQlobM3iNrTtiOKDn7+oyuNymUZKZvZ/wlxEjebaXDJ0K694Hj41HmoWaqIApunBing0dHH5bKOV
8XKfNYKO5RKVIICc8J9uAaHCEXkOvRGlwp2IMHS85GoQ0KBUFHsplrHSLuqS+bNN55QYruz/xboO
FtTCA+7OCjw9QN7a3nv/tvpq8ztb+52twObFHrQ2RoAmtjofUq3Zrotq19m3YKex+yCEPba3/oJk
hUcCksPzqS0kikqVthKVVoXfdajvw05QT7RkBLopAy81YCqc8zju0WGN7az8jSP+JQurhYah/Tgt
8vmbwJv+gFQxD6CrYbSEPS3z9sxS20BxzEbTH58e715r06KSmr3VNYN/S+WW+o2AxwF+6e2FPwza
PP1YJF14uroakslhgv1tfOEVYcwjj44ucexpsNKazd4jTcFPx9Sb7WnQlData1wnZ7e346PUOjxB
WIN6ETolFleaUDQI2BMjaff0mj7acAB7ISiQGYocGDy2FlxrW3Y8v07ioos3wqKbItjMwH1BTWeJ
XYLhZxB5YnTdpSthgLdbbboFFu4AO63uHKjThYLN/mcFqK7MyzlU4kPaZAHbQQzro5nnoZ6JtE8j
2Lo8fe+Hc7gKjQSoXsI7x3/xuB+8Lgj0sLG6mk/AlEzxF54Mq50+cBSHkNDochb5AEnazai+R1jl
b+kpZU6QYjRCqKM1du6Cpak1HvEmpoHVensMbF9cKJZAunnbEkevjACIBMrbBAbqJw+O9wt5PDmk
XLhV4b82oX3VpWWMOHt0mun/fP2ycRCeXQP82vZXHFi2snZxfnaDy8HXw+r/Zb+9bsXErURqrCe1
jD4x+8nfS3OTByHea/1Y5Dd2nJxqJ9hAGooy784h+G+bEt9vyQE4hQDu7EiXuErn1YkGlwyjJO5i
pOmOPHCMKgfa2K3bLrmepXFp7a11a4DKA/khaDmy3K57mqn4NKb9ehlQDHpHCBD9yMTuEEtZ8qbh
UjpoOzkzuiQs041/biX/AOVyZosfPpePOCObMO4GgpA1xcAsEE1cupXuk+IMgW0nAnP1TVqjmDGf
OaxlavzFnkqJL964IPOFkRYLwazsDz97QqmubhvVjhgh/hDhzuKak+fi9JVTmCgJ7m650zi9wcyr
dXS0BGRoSBdNIhCAaqB9zmEJCiwSdSm99C5L4xpLNOy/VGhgnVUmZWx6EtEkbFkjSOtzbVIB0y7X
MB9NtwEMAxbMpNFL8sRT5UropDG2Vre+PS+orsmfY1QkSWhlCpVrxQrgxT2EsK/QI+XzgCd8m/AI
vGHxj0YIP/Ikqh5M/20NVp73XvIG+unUY1eOcMSG8LAavHCWPZqavntEN5GnkqTL7pcoIw8kov6/
xeUeN4t4SrE+2huNj//oD7+g47GzWVZNGof3sDm8nlb2/f18DaQXR4ZcNiGxeZs+yUwmVFN1msj8
dMzUAi4todPNBK7qYx1fU4Z7c9r25SYNHo8bceXqeUSyrKGKDRFvpXu5JVz3t8LLFzJIbWWHjJN9
66f5H23WGJWCa0FAvzvbOKAYagT8r7KBXbuYl4q+YDLeFHb3KAY2/a+NjeDxUqGDky3s2652Y2dS
lD90h1vP3m3CdJg36FwZLfFLsBpS9ms/fF/7r1EEGmcXlO2GPqGunImO4L16Q6TQzjiewYwt0nui
nbri1TMaYyiTy+GKBGQJNhJT09+sb6cx1HZH5F0b4xlXRxWcng7nnNsSyle0sTsu0yN7CvvgM3tI
MeR7jTzrPU8uF4UK6cJahQo900sVOfenRoqbnlXqsqTo0mQI16ewDzUASLsZnv4fFP8eGXLJV6Ea
2b/AG1dsYBYB+W5LnzZhG+ucVu4N8al+dOp2bXCuUli8x2aMNip5HLNOzbjSlfABBiBfVes1hTsj
ERiAD2hI4Ce7cAdlfVI8Oyu/QZPBntAuR48lOiyRfpqdjRrTlBLXe5dcSmRgXDszeyqW1tZj/YKO
9eHoxzwZDhU1R2GWgQ+fA0584cfV8PjCEdWlR11JUQN2o1wqnJY4A7sLoKubD6VRXh3KIrgsqiAR
y5yLA69cbtEaXKLCrwDNa7nsCLOglcrRSmk5FzqBKLDtOUWCxrrAmv/MNIAlLhK/trkUnjFomkJJ
ThRiCQKaRRC9N0RDEbFJGXOq67g3OwXhSDDKAUASH+RrVkzfGdMxUySm7p63sN0YO7RdsmDohA9p
hEepYsmOBmkm6ityY4lm6yroCYhPDj3nX1HPLP/vmicn8Gz7nv8AgyNN0uphsj7KKULVOLvuxtps
+6Q4Fr//QP89khcX3ihJyLbpQTTax7cudspu4Y/SMcB+zezCd481jz9t2dYGP9jJAFzimUOOCpTX
DDgJJhSgveEtfRh/CDnKqFK9jG/coNZ5wJU/gfUmCCPPKg6Dw9QH0P/RkwpEyiVju0W4BAz31aIS
lBLIqqzlOaXkpuZb7O0k7h0zbzzXlRcVu2F4WSOZZna4XjdGFV75x4w3OJRFmklPuuXGf4HCsG5r
oMp6b2Gq9uCHZdFNLqoydMmVg8Q9IbJeUkCggwm0aKzuZfkjY//dSVvPuzNjyaNfLY/R/We13k2M
FlKDSlaQ5SHBih/Rgh8+g2AvER5Jo1RCzHLIm9C2c1IvatZ9gqtZ0vgqH/dJe9CckYPDS+jqCML6
QijHTgLgCKUklngqk+seToOJ4Cqvox6i9z1+Me6bq7ciIzHsuFKoIL0jLB3mMHFgWHmMumiDwUje
/PG0LN5osYMFYqSFLsYOpXEZlM9yDJ1wYChDNsxxrG6Uj1Q4dkRRdBEg2UsvezCPvxOWoiUEkXKz
oa4taLwp0Itz/gkKbdFuq5VR1PSo4PIGxI2MRkcZ9POlO880pbfjP+6tAIQRmLHIACzairHvpnu0
p5SR1qsyuJHmPikp147GtpvieLRRg3pUeuUg8EMHhvpwTVQ1FqBOljKz85vH4sRHaW0YsYbAx2IT
w6LnBVgfH+ZNKVt+zX3SBxZqDKRwusSUL7mQ7bBXoy4RjupqDnx8pW2bGPGPeFuP8t0D6cbfzS9h
cLM/xwE24dGJpEdOeiByUe2qnz3NU1UGOSCGTw23ha+J0+q5Xp9SvjTVZwopgX9Asf4II1Ks07/8
IGT9r5nlP71hFIqIMU+t2AGklK/fjJmFE5JZjzSMjTV99nyuoBz2FVsGJioaryebAnxgt9TMJCWj
lVM5Oq+EzDs1Sr5OquLlXBGdbTo1Y9wQb7eEBHxf20bTS7LQJ91MwC7f3+MN7SnQRCFTDcgeI0yT
c9K75bhd3gfovQp8nRkyVESedaeVhS596CjRYNoOC3SajPFtu8d1bE6OGNTo0+hP4yAQsH+BsyMp
GMpKRxURr8N4Ov23y1/FQ4Rz0BEns51/oJOuICO5GQt6dTvmcvwGBeS8FhDGRnZS4sYp+FNwsRPR
3a7xvpBXTa22i6zBs/IX95OW5WpWsmPX0OPNnlD97/sG7Dxa1RnSA4O9ByvDcKH2lKRi0n1MVG8o
kzA6o193FRaQ62tDQDtp74H6joRB7Olz68X/7YPp8oIKmKMhHkw6Kj4pqs1eD3yDFvW1aJeG6er8
y8huylk9RpcwW32xk8w1jMe8XL+m55irRVRWptDfbHhvB5QptWxZgR5PTxKZNiv1uhWBgpoaRVbt
Nf0Or1EVVTwiYUPqXJzIqz2ROUuwiHHkQWpfB03iLBlVkNewVepVn6cdFerGoFJP0/e0+c70uoDz
/SYRNPx9R47qBvAKJzYVj0ygSgxUl7iUorPVaV4u01qP8YOaJIVVftWWEfkqcnGKJIbd/1aQjXgL
ScerKY4LlWG9k7O8KAjwDzEUDbpouFrCAbSvIWGz1Oc2rzvZeSPdh61jykfdPhjCfNSR1isECHS1
ef8Tn6AOxrRhhIBFK7945pgyXcMENmgeleVwzfKajmIk8T5qzrhCkX9yD4at2uLTnwuqP0ByLpAt
k1vSNDx/Za7iZ1gxiOibbbb18RaBUBBDmjl3h24myQz2lce3R4QZlCvTwnKKkko0QueZZd1EbA5Y
FHKA7o+UiMWYdyuXmbZqsd7c8e3ByAC6zPuQwj4CnpoTR+HFTZzw9uOiqBw06PcJbBZp0yngI4m1
I4iYuBsPCCPt8MV0x1+/RvKTAHxfOVlVVzt+ULmfBWf5W2KIK33iolghkzwzR8ZYyZgzS1/v2hci
Kj303ltCrRj9I3+0PIQB80550hHYLZc12T3i6OS1n+OgaXVNestIns1txX6xfuBXVlBfaMn5tUkL
pzufYTUxBVOzW8jS8A1BGRjeze61pOFFjRlePaBVHzq+0uzHGdfbT9ouxip6mUPqLaQViPzL9YhR
/iVETsnPTB6ZWDfcwcHFhIAvKoE/0+sJi3Im2yRUr9oP9cp5RXKFAv77O4bzp2aod7dKRVUKPrRP
SkzdaMogfxvSQwvGGZUEzQr7Ebjv2A9EdbQl1DgdTCRwH90bofAWxpoigEzv+15Lhvtug31qgfTS
P8NjctYwe00g2GEVIVEHe03l0ndpE8A8loXFlih+JvkKG8IRW7GimtQYWqFxL45ifm8SdoIAC662
Rzb2rUVoYuzaUjfie58Kkpgu5/ODB0wE0YiP6GPOTp6m7zornqHhjyEDjiWStl1rafpL5cwWQSD9
uz+3Wmxiq18dQK9JnjQx4EaWEtka2nis3IdX+HimgVk2FBcNshz5X0uUPdGhuNQPo/xxKq8YbVB5
ZvzNhzbdzBE+4pu7HAt7PMNtjC2zCu+nCIuaYzNT8VTFCiUXit43keZPoP0/G0mLB+R2f/dhy7SN
TFvJkgnS6CzfpBb/hi22sReXvJRXmArTY820QftB9cUifRFjkfaMgjQvVWOfTisNnH+jRvOe5LAI
uUwk3oicAkstKYt/QVURWg04D4Yw8Ge0Mcm6QRYt38ouZiIAzwFRYKKX31ptQ3yRqnHhX5PjOkXP
wQoFWFKMf3PhkTsYC+sei1OxT6tUE5nlcPMZQOB+JeP/JCa1VvvlwRGntBaPjrc0Eu8r5j/7EFWa
C3uEcgTuntSMFIvBHi8cdy6IlMi+LXC94CQIzBsmPXWku/VJ7sQovBtFA+qAqPEtpPIQSpxVtRcc
9OtJijDCsQNVl5k22wYNLhejz0Gvi+zFTayvF1/gWQ80qOlB1dmUxeD8t1G2tAAMhk2QG+vwwgWo
tXK0r43BshJ9iKFFvfBVYPrgwiYTNR4YHvvDhWPHB5S8ZBxMddtqcPwVoAXE+5Uc7eYvSEjzyjxG
R39SONDsKNMrZa05aP3jaQPzDR6nkb6xT4qXIJwFPlGPPYvriHLLk4S8G2ywLDhFX1iNJ8cYCdai
hddP7NrhU5bUCVcAD+p7Kna5ROhslXOeMpDoq+PgWmrh6SyOwtrdWuB4uWKCH2cMqGnqSBrHBvLd
dLS3raK4cfQXQOQY6xLQuh+8mihJTlusHENes2gBRKqd4xOYbx/p4MOBSgNQzrgydE3dvgKBu+XW
fpGfZLqZTaNtEVJ7L+dp+bRCY7eUIc5Nw8xMjF7fKCJ17TJ288fdDg7e6T52SYSTI5/6DsHcv67E
cSGzNZho2k/TPWu664JTABTwPSyWNlVtTbcNZ9rx6ZoO1/y3gulGRczd9se/H5G6EJ1hliin5kBg
s07Ec1mtu8qQCPHzVid+EmlEtQ1O17uSS50qZYoQoked1/U2+GLqJSRNN3ilprYPRfrtz92klkP8
GTYoMqF3ueOXvQZWNdRLBERMYOmUg5/eNzMdmOegsuJf4CdC9Z7OaOky5bkx/kyviZA2YhrXkWro
3o2Nxa8/J6mt8OpamyY4F7sJyo7cXM8I7NooWeeSeStb2jVqBkY1wOfVuFUYXws9k2UxpHGMY37A
q9sv5eZAEJtMDBsi539UFZSaBgmvw2s6KoNMv5CseWCMXRSCqxJnh0fPHRCa3E2v35R1YhGOtPMN
bcfLufTTb0m4B053o7JBhmFXuKcUGvRHEgia9Xflfn46378If2iDObO9topz9zd7VfCJhgm3J0+e
JJ2oGf+GDzzyYK6D+ifgwVd+Qqxkw0LT6WLDunWpgTdYq8v1e61zRwX16pub0ud/QqDfO4BkOQxj
ohgkzrPx7sgGqA9AS0JD29kRGrUFsEvPmcRCbDJgZ9aWD1qgfrKGr/oXYG04VpC3PpkPFbUZJleI
qDIHkpRAv+Hoi7rV0Nh4uye2L4C7uw+blrGKNRFz3ln44zVhIQvVEWMci1OcFcCpGPvLNwD/NqCp
dfD+joKdRHS0JOYVhRVGqs+UHAUJuFtqZ3lG064TFmkS1MzkTwmciPUMXQlB7a25R1MUA+qsxYoZ
XaDUWDihiQW29lgqDuQUr/XKpEp9eBwt/H23vw+3E7wJDgUdNC2y5991LyHIiskzutMNEe3LzE5Y
LnaBw4qAaeo4V4eNd+5CQVh+CndxWj/QLlHwhnLWuWA07kELwJUWlE6OgqjpNxeLw0a82OFIYto9
eXIkFvpzX70lrj3WanxJE7+s6+MZVsNecqPTyctblnL4lCwjtOkkIkmyL6EasGT7qjaK69xAiaqC
w1hTkAee2nMEpuRgznasuoVdXii8bfTznAKK6YqB93gD9D1y6Fmc8/e1NmdZ45YptvIVoAMpJij/
nL/OY2vWxqpUsNXOqWKGf5V8qUYXFnocipMH2N5b6ODTc+wC///nB8q91QJN+ZmkVLkFGBgohxwF
H4T5koX4l2BvyJcH2/NlMRB7tyK+dCcNB+9mydIcxxOfN/AC6ksWAneh9diW3pWoyNEd/mNGYfRb
wHpUl+Ntj6I8SAV1Ma096eNNI5zGuq/LcO9IbMQGGuW+WdqymuYv1eemuAMi/ZJFdmX8t55ImoK9
mQFzeMRFpYYfncvthtmRwYpBtj8h5nNvsU8io+/OCoMJxZLPjaj7/+qCfon8zT/UKPmO5idl81qn
1tjys/UXGa7om/8b3lbEDK4GSnIsd68d7nWmObacMIxt5+wINlIzPI4EFr6hsUbw+H11gKgBz/it
X1vfWDYvuLn01rIwNIEJ/1OjPXzQDKLVcam4kSTvdoAi7Q3DKApdoG+kYNm54dqrfPhXaQC6k2wZ
98QBJ8XwzDR2JQY3kW1Xs7h4TL+XKqJyu5tQp+d0jq2YD7oWFZebImgzRYW5Xj3dKmMbd2ysqOhH
5q/uOu0PIpxZX3PBZdk7+tcn82wSplobDCxcjst2xBqbqTTwD4vpj2QACOdPvOBcSlq91NXfuVun
WXVklxjSmH74KKXCJjLs8FgJeu8LUZsQGy0YMMyS8J0Ke9aDgkHfJXw/VTCqUk0HV9ztKA8XeZiH
TJN3ebkJBOqcKjQGNiKFrliEyZYUvNl7NWK2hqjrfHeAkTGf8X4OTx0shAuv+XAfcJJ7WgNy7Iua
XOfIXmg6bRqW7sKPOPbuCJDI/6LUaZVoUm0Z+msREO+tNh4Mr2avlbunlgLPyhs0StknbXFd1tJx
UJ9wVkZkAsGotVvfZumRF3DqpXRN49v7ZUQtWCzQZxE6H5upAESYSCeci5IbYaX+rz+K5O4ck4K6
z6eSuhJ0wH6Dm4OIMsWWGuK0emsdZ422SQHqBO6tjc6dZFiCH5jMJIb7oJFIFQFvR5KIMJ8tKEXq
jVo219VX/81WaNkq/A0VG82lMRYFbOyDbk+riwJyd1TaGoq0jAan0tkOgaNHAM34tzZs4f/XVtLS
smbYZbVoqjLJTEfCNYjK/BpUzABEE9SbaX/5naykI+u6IwtEMEQRU4eMYsdQ5zarnWoSLZf2vx+s
qxhEtVTrOgvNnJnpCyq7mYquZZLk3egU6twBYctqJmwM61GUFgHou7MxN31XnepfdV39llGQlmWD
6p76w2IVauoPr0Ln8GnQObHitvpf2rn35rL318GaIqGu4PhnCpNFgxzvnfwIGrrUeTyf7Dc/lLqb
X4XQEIIyJFRn1LPP7Ure9ipn3LS/7HklyEky1sfbqZmnYzdhaqhBUHZuYnE79hYUQNaPTplL1UBw
8JzujE1DZI4uWnHdIH4iNlZG7fH2hAmELHpaBHYjNW0xnBDwl0E4pl90lFXTfbrbXhTsa9eUzbWJ
cOoIWoTWgAKZzuJfWhmY54RwvrppUO02FqCyjtygQ/TofzADgBWfc3+vBF7syDicehtpl7vUtBZj
E8f5+Us5+vSvZZxDJ3uYEv+GpcVzxIa69WUzxhBJ1YSdu6hcsRkNWcUmS+kPdbSsDww0ZaIfHOjp
EM1nWPh3CL67gaAQ7i7uI+oOVt5KZabdM2CMV26gjIIsgGmsKBvjau/5RQx/KOdAz3xHuftttpeA
UHUmuTrjpwMlRrWMYfocEnlgoNRpjplJ+ep7h1YOWh8ALV+RxrENhTxf/vQZhzKODpnMVfkZAxgt
rL0uMj9xPt3EdGL45ozmMU47zUCy6OOg3DlEmGJaVk1mrX+6pAtZftQqWaZZ9ThRY6ucsW4gmies
zBhxMTMCch1XcF4Kcig3CILdGVBJZMf+b/t1LZj5SZ3i0CTAR+gYVVvJz4fN3ZE82gTcAiS58K2o
nz4uo+ptorgH5a2dOVRfMqQzhc3ZP5p49kdA1tR6ujw0XH8lG02yhcKXB20tMttd7tlWvR3v/ck/
YRm/WQb0gFMFxmgzvEwfGbnkiUJwGrvfbS+2cpB6n4c7c/o5xwUxmgdJHbEcDi0KqSp47CByn+NR
lizkp/2hBtLgvTRY+FR/rgOGLh6GNZJ9CpjTLHY9Uz11Y0/OOfEM4TF2WVOQWso3mAfEqZde/iow
6+jmQBxOg+Qa4vbtLseeWPa1ksVTHRrImNsMAf8II8skh1g8+VQQqzU2W58OyuD8CS18DMR5c4ZC
aE4rYuW06OaTLW00d5Jh+Rfrq4nymJf9gKHOngaUtQruQR3KVIlEpxSwnslnUBfFDCc7fD4tai7C
FP/8xhiXSzmVxdNFNzCL7t1tFHB91/jVrpQJbZtBOyFoK6hYLND7zwGPqr/TQGJbsAAfvdm10crM
nZzCrfMmgaleHqocbg7cwYyKu3m0UB/xAIYtoKO7K+xZPyS/2kSoFf9Ma+fTeV6VP/RZRjuh28w8
Vd34tNc4mhFMtPggmPcnikCvXiLphoyjk31dnCD5VB/Zcwfgr0+NlX2EGGJWOWCwQuTk2s+DTWd8
fpYpgeNXEuE3iCYe/TF16ZwCqPWCXJgbyJl/wjdsXE4C0zajupJBrnFj+keLA2sgVyVY3vZsjdtz
C3Qs3tYmJKbew8iuuVBVB+fTPiDRPMyqe2TGGUyXSVIgt7qtjQEyjSRYK9mqSkxCzQFSDptD72/d
BYzB44e4AB0+apCmTJtA8kH7yFCgJ+QLrzJHjVcDVwgD3qKb3tbnnbR21x2a2ocnimT8P8sbfrCI
+tFF0Al8O2GtsnEoCkvHnq51tuyGoCg6pRpsC0AUOFZDjHfdbIHRozm9tvSeoGEnBGIpAQAXJde9
6SbvHR1CJRTBQvfj1Sqx+U30+zdLAqqYeO7mMq0lnOcQPkPyr85m+5mHRbBD6MHC1oi8ZTlZDhaC
MUQ/2LNbBuN9s7TiR/Fu9t/QGWHtlb/589aEq01etF5kcd33qYQZiauC0k4XjJ/9vcZg6zGaiiTH
gRZNjy2QaDwEQ2SRdUf/dI9NlTJLas/TBjLaFTvo7jxaLNeW7BtBuSihnErFisbktuvUB24pjFua
3KxagnFDa1zfCVjUvyQ00Q62N33Wn1lWosByHxXMNQidTwI1RJenar+hv4zw76o7PDv3pTjhaPkd
9tmxG+ql9RZzys4Do5TP1CbTaXqTWnpWLalpz+fbq0csGMDF2Iw+kYnYuAaAfrhhYNl71dingIJL
oIE6y1xNu6HKnV0GeZtjkcOZ+loew1VlkRBGvVsn7zq97TbWceGN5AZbyeVgdHJwZZ6xfl6XqV6+
yZWfHNMbHY5wuikIPrYrQH/JnKj+v63IocbFNZJBSucve+nZ1g5sNNbgzPL7FJxWQj0As/p+Q5xY
ygfdSDovMp0BfBMBrNSXofGazG6sDUkSmKn1iXrIIlQ9AUNQ//Gb9OD7/dNl7HN5uy3nc6iUMr8s
F7Q65L/3JEGrbjVCtXEJuxnjrud4dmiroBGmVh8sq1xyeIMcosyCw6ZGazfDx0xCrz6YP1oK4Y3B
5wqj2Fqy9FG/akhtSXwrDlGNOQP6nPTMmGkOt11TIrWBFrExk8MgwoAmtxYQ4/nqfzD/E8AETtuI
6miZ17bcVH7loU1Au9JBJvMF6DYo+TFiNAHyp3Dxt2UQ4v1G1Dp4830qU/lfcDmaYc3j2VIMS6l4
H+CzoOrDRvKdxtxTFocUNe7uAvc3KKyRM2qrTK9fag65mJQ9sirdUgCqWdBdIDQpRg9+nKUFNkxN
1s4wqF6lVLX9nDz0m51yOQHkpkpCagWJ4zD70qWT/HUw1Msy9tI+46SZhUIL28oECvfXdpTPvZNB
QTNV+9TqqOo7ya2J1f4UGdrqd7Y0nA0aAqoROj6KcZ07SU10CZRz2d7PC9jSq1zIV2qwSx8yr+ZR
LMIk3QNSoGZ2y+cDhbe/D3lE6iAuZ1YbUdcjLr0NTbWojLTaQfq7c6fjUM+YAvogr+y/gQTNTpuA
QmC8dzkdfsiIKJiFl99pjFQluY10SHc5Tqk9FZAYX31DAlPRvZyTMDax0/L3I3w8rDtgQmKCMXfy
AKTSZdcCXz9Y0qQjkQiPv13S2WvSXL9RnFy/6qdwCdIqigvoRZSu0mnEzxGxgGuXbOp2ndh4bl+o
fdXs+CS8A1dsI+alDfjo8+QAaGqAGemKklPioKL++Ct6V3n5EaeuDBIPWIGHC3DBF98sRkMhkQQG
8ddpvY9OJThBwOsU51rsUAPu9Zi9oosJr5Ms313o9ny+qGECOoO3Gp+9mtHf/uFFhf5QwiakNM1/
apEiMmb+d8uloY8PPPiA94G1cCI+n8FUPF2EmweVTOHT1QKb/SAflbrj3SXfrbcd/wWv6egWb1sP
d8uQ8GvAqsiz5yKRsaZPIlkKdidd/1QlCp5XnRsI+3ECnM5EdNvtwv4gxlS03bgg7vIMorEg1G/A
ZSpgueVqLubjH4Xyx7Iuna6UcOTIStRbcmojQzDzb0Y3HXp0PY4YqVOlQy8HWxusJTTQPtz6vnYL
3iF6od+yIt2Dd9QSJg+0pxitwS/PF8ZhsaDdKARiS4LKtiqwT2RFOBZAF4l6FE/tSsoIbmI1ffMh
If83vmYJ8wOUkizn5PcHsHZL72AnFKG8HXLodLHO9pHJ873LBsNrElDZlBCBJJn42OrjuCJmyBm1
ZggUQlSJSbXi/dV4IGRZsspGtP6b5dGNGSKWEt/NGERiK20aZpnv4N+DAT/s7c5D1TfRu531MDaG
5fE0dPtcxnWKV+mRUwsFLQdMw/EcAAKDB/H7XiFBJeyYqAvGBTcqfIq7cszf+w6YH2tKc6Wk/Ov6
yRHdc76zHjuawvnCoz3mFESpPGI9O7cvoGuetQi1sNfJUcQREbTK1A62Ypq7+erYSaWmWi6YdaEQ
Nlc4Xgr5vLFAAkohDGxUeZjearOkINjLCrjsiu468IZ+EGtPeEdK1yATzg8DFtP1A5g/gOAVvH7a
amBHMwbfNg5Kb+ZfhPbHu11PHgXomXQigprcz3q4pcnDbUYOCgPld1cz5ST3Be4yDJ0pFoMpJA+C
pWmWYlnCO9M2dGG437muC+u3nc1D8SDXefD2qrBAV3lbOqdAU1AVwV+R6OgvAbdMi2eO59rMfGwx
Rcd7dymTPvJzu8m6XVpioteYdXTCsDUzF7XbOa8zeZsQI9ANHv53uPByLyS5wkYU1VA6D4/dRgmm
ssN2ropjGW7AXkgoeD10tTsa6i5Fy2Q+xUPZx7QNw0c2Xla7n9WuWsuxMCCGwauImwyFp9EVq7Vr
1zME/EqxoqaHLVKdN55HnvykFNKqMsckXtZzUqSFLJiMh6aeoONFX2ACJqK4QlEzaPDhoSUq1+n4
SoIhOXf5MYCWj4rUbVLzvfuVhK9ba+OyHF1VV61uh3Ma0kBAVuHYLAeTIRYbHtNUUuA5ZRo2e/QM
cXuXSV/TfqWTR3c3ckTEtinPJKfmZABH2J+mCIrdqyvM31/e8N4EPR7GQIlPto4HIk62wwN99Ma0
Q3+DT6ihjPw7uw/sAhBmyxmP+IlDRibvc5z3MvrQuXpNQ3KVD9atma5kmDFXCS0Q/KWZDxKmwtF0
MWf44gHrN4yPoAyuGBlBLKpgMVr03h+x99vj4FuM58Xq73mEBs22YXxL06JSHkZDXZ+/rKiDRtAV
6RuQtiJd/y/Pk5E9a+z6wwbAxHGe2pjjexVq+/5oKeH278WKPOY1/kI4lpzT1PGWL4zVwl98+ayt
vPE910/cn4giI92y9MLdkaAzT35dx6G1zvapb/puPXaMORKTVSyB/o/HEqUQQTBOAy1GSSQgYpjt
o0CK0j3zOqD4diXzdB2Z0viwV/dXsxpCXfJzb7dIFCKtgvVlUGvzLmcbWpYpnlw8nsK752ayUl/C
K9egFZjAtpzPVrRf86qENM8Kn3QImG5S1XSHMQqYkMJnPAV0B5cTa9n3EvIQ0u4oaQRm+Txx/Gmr
Ti2SxyQI0OoXqOsnpj+wWdAdCaWShQ/NhWlSLIrtLA7PTAzKbNuBqepE7QtGXCZmCifFW4YgyCuh
ag2F60+4ok+0CCgL7RJ9ZnWi3O845cDfb/7Nlzif3Gj9Kgipx5O/NJW9Q+H5xkQJ0SMwiv84VnjK
KLr8qm4XCUz9pjusTw4pG5yvFzlMcS1Nd4qJ66lq1PiZVCmFpFNan5lYTWy3aOq+gMYMDiNSSWP1
VJO0SE16Rwrrmotx6XIY7FUdt8rxkhyzK9U/fXMlCTbeEGHjEMh5JmluTNV9JxiJ+ak0FyNx/2eU
eHRFhW6sTYbH27+O65Q+FgLC6lL7LnlH9N0wjZGQVZ2TTOUk1smP+5ZXqyxoQJb9qJDmccjAYzjD
8qYrMuzJDhauu+kjXb49t5FyEYC5n93kdfoTSugMxVdKu6MNEmJIt+HOxOzMPcb4bv+SSYmeNYIt
lFAbDljfAQBf6SdAnHlnCnBAx9IPtrQvaUcas/qMTh+kLJyFKe9XdB0cUS/ftv+RTY24WWIJ0aV8
2XYBuP9nIJgv6nA4deBNOp4iRiSBqJJh6Y75Yu+tsXdzxwI07P8OQnkvJOptZJ4OUog0pY0oMPP5
KUks8/TK5nKnp21r6PI3bj6p7P1GBt8tEMNBlRUOEg41kec2asjsrW7b5tQ9s/Z1f74Ueqw8CJ1z
ksNy9tg6fEdmo3V1+u7ez4hEhuaF9A9lhW1F5Iilq9Bgg+5DmY8zjEg5wAIJHL+s5lXQN/+4RfQY
0QdtyhDdQLGXZIe7yl/WpanKRcukVc92WoM+NiH2HTVof89ll+vXHbjkmkxUyn5D4TNwBXWWBJI0
gL8ZYyeIoahtwCz1jRsmIINnLgSTSTFU8PMk58hx2O4rOy7n/fpCFYjG8YPUwuckW1rnPPjuhaZc
OXTaAvDSomvo5JiJNA2awO5sMZJtj5pW0vaM6Ef7wdR1be5UDYMyP1p451LmN/eYk30msCtJIglK
7P5ZDRODyR3ogZSfETuGLz2iaOWwT1VJNSgJeho1PaoBNXdpUbv3oBQ4eDRGRyPqtf0MTlYH5GrA
3qi5+hxUHCm5YzFdK8YWkXH35MPml8WwGFflVws7N+FHwI3+2ub7zQa0EpArbRoyW4e635CQk2b0
ORtzhvKjSzU+9VVCDhyYqOahXDgl2qqaf84+8P7jr04jFBW62Hb7rlUbSxhZmXG96LvShssAepTa
8yBcBuP/wtMJfdO2rhhdgrTs/IH/OxPqbHpHyDfr8uXGRYp1UvsUMbdXJmn5OUXnh1pwxCcXZAtK
T/I/03nFEtcCCTAe9Rsl8/wcSHE7Ow7SvoGyzLcxbyi5cEiDbb/STLC0JQTXtwuP3j8NukFIMobI
5uPYfd2PL0HHBQVMfVzRcyN+5k2weU4243G2j07s+6X1IOqbjLe+toh2lBRxeucyB/kUKsk+hidn
dHwps0UJ9Xyj7wULISKSsuEAHK0FdFE7s3z8am44b7wSP4ibU6mH2k2W33h+jhFVfRghx+tnuTwf
NdqL8Cd64yGqMbJnD07wO/Yf6ruGrVIEoB/fqzivbqQ5U1wtxs21FgEYNNBy9QNysneWWIwPnU1B
cMFm4HsTulyClJBs1b+pWH9paJmwDu0IpXUjGzOW+rMddNO7N4JaszoKN/7+daLN8sxl6Am20sIs
j3yH47DZm9hMONUhxIbvBZ19DA4QsfxLti3sbwb6abysQky3k+0fG1nkHQgHqWWCs62rHvAStI7q
DYSbOCSRYBG2rJAAmjoU1O69j3nANVpEEUN+G8JdrWMQkRZGU2Co8mdnucT795L/nD7vhpM6/27S
k6yEjoOJ2S/5Xbz5pMlxLyKCA+NqR8USitseoGxOUcmdW18Z3KwDOJxOP+OJM+9yBhzCyHmcv8zC
LJ3DA2ws/mzTDER/LC5nI4mqbhe4vrPk325BuFyBqu6/YCEbK0Rfjj6ydgirAOhkSSjdZbv/bGgk
t2n3LM32+LC9BrxevWutyti5QOhh+w+gRvBrpDLWojckny9FPZnZIQAqXW7LHL+fwMFoGOysFQe0
rdGvvWP6wghF4xaXdVGibi9/eUpf5JlpX1wfN/fRxN7+7uMJrVB8zKJqyfFGfPxUhKXTiWdv5Dtn
JwGBgVa0oSFXoZOqwwpmCnrNY4KNEWOuwfiF01gdDu1F7SfD0N5fWDqh0GgCKhutOTyO2AA+hHpu
8UNce8qs17VTKflYjUjp/x8cviHpAJc+hCA8IM+JhoIV2zkFcrjBOyzSmWeW94N5egFfbTMVxjMl
2x/HNIbdweBlVchg/aePVBi/IlOqK6fmruftvICKta93kSoBtzjHMqukYwzVSOxJkqMORwI7HKIv
N2Wo6luN0IBNI5vMm3wDwVWqpizpbUlrZ/BKiasd9quKFcbo17kdr4r5ODLBYsGvgkmgU6qRore3
t1ZOAvMPpIAIpAv8366/VBJQkORjQH2NdDJn7xqdVG6CqeMElDuAsrjPGkb1iO/sWNnCtsgb6gx9
9YsdhcCPjPoew3iXP50+kU8qMeT7X910fmiFFjMQVA/RNnAP81cEwEpaNsBqsU4YjK11hIewZY0V
oi1mDN2MMTVT6bEOGWSzecLjipwMc0HRmhMqpzLBNEjc+qq5+ZZvQjc0I/ZaghDbSYk1pEk2vf5h
M25st34D4FgzU+3sRL3Tfnalxlw3khRdDEGoLEIbaM7VXd3VqHGAXbri0M8e1wgW8F5h0cnroJU7
mWgekWIYP5q4Dq7d7uufaypZ5yZ3WZMOoWbOgSW1SotOIunGrjUh911uomEmFwwWyD62R7DCkB3n
HBauTh9iYxh0hLkMj8OiHQly9coEinnibwBSaB3tdWeui05aqjxk6uE1WqwUeZZvvAYeb4PmzSym
zA5qtmrRvQ5iNFME1XRW2AAvtVbZqq0rLbcqv0ZDH1C9cGfl536ro8CLV3ahF2kC1MStd3hhheEZ
TxuE8ai8fKTTH3t+Oxu2amXZGhMSVtCOnfSiEekmojxlfeXcqATZykov9d9sEbW427KioNi+VPbg
7U/C40Mo/zQntqRSeJNI4hYd2Ryo9/wzBMKqPcCwuG+sAgWoR2xASAqnxM0HtZ0+Q35ZBbxYOySN
I7zAuHPR+Jrt4BONApfnPwv67vgjWXqrafk19KBRw9VRf9vY4b6aXnPzJ7kdHf9J3C5n3QHQKZ29
aK2m30Yl+ePGOU8zc41XrAAeDhmI8WC8XsUj4xfXkRNFWZd3Lh4RHT52c9jbPJzha/LzxMz0bqdy
Bv12V2WEj9/ajIfn5I+QQJB3D5+TQB+o/WSyCEqJIUC3LUDoDVDlWP64T34NcRCZx1TFdmE5T2VP
au1gApLYMUI/KsXqiCCRDHI8OsCKTAX+GXQ4xL8nfpR6DciIGRhRL0C3Uirz3Dm7/bO09w0BI8EX
m6icSljreS6Sl/2QJKABRV2KnKo1EDwB+uWcT2EdEKAFvPHaIQccw3umEoQabfIFaCRQ9IyoUihh
aMQAUS/IEKAkPPRIlRQ+/mzjE3kjgrwrVmNfb3oTYALcgdtMCUSAivbQWleoXPrQIO9M0+pV1rzA
P1om8braSCPImBdp5rle1O2vT3kXMap8NZ+M4NxN27mHvUCsBNNtT1aPc+zQj+HwwiNPiPiW5z5M
W+4uRxbOIlOTZWx0tvjRT6eBGdV1RoCwQUDj39UzqkhJORsOFU6OLQNFBrcneeuaO+oOtdkVAZST
YPvP0qoZZ32sgOXJyvD9G1c7E1iBCTD0oeHq/DqAOZDrez0lyUPyFkbkYf1OtDzAmA0elPCnm6yD
UANZiqWDuogwITRsY1a68B4b+I40W9bz5YY6M8Zsw4gs7rDBp82WLWWIrHx7mMI7Bx3JXTwQ6+R5
gBHRrIOhq0oy+sH22TjjOYb09CCDDIJy9PhFf4XpM4HiuLcwTT0hAypo+FUJl8q7a6INn9+Z7+H5
BtB45pd+GMEHyI+PbAXra9w+RELTTfXfkEhA9Ui4UeJCddu10O7/Yvh/4JLO/uiOi4twCbZhaP/1
2r9IkPxvoC81UZMMUhkwBUWxEaHNHoMusbV9xJ/b8CwQW7YlIZ24fUDS8iovnm7fQAtvmVoj6sGT
4Wqy0XBbAAghdLRaK5+la5cRjULSP8m/RR++sGaxXyxhspUxOdqK/af0ecebQvzlgBbqB7o5KRgC
YKOFobYlI8ywGa+UY55NdY35my2bSmgxhXB4wk1RY99RtUEMomziKFzOC/pxXi4OXfR8zgE40pUR
l9uEJD1dlkqkAH64aAl/XvfSYCLCEOUfe/JydkWysfPdShnAuyaZuanLMrHsSn7sI9lYZMN/eHBd
Sv5DDbscIXb4phBbYCqHCwX7MsUhW/sw/qbWcbp4PmbBfeVtyxt7mLSXpawEcZZzazJgf4aqW9cW
K7ndRrRZVbMZYoRB4f7C92dK+jNydZ2acRSIAl8smKq8fb9JbPCzL5capj+zoLD630cWU++EByNL
h9pVhjNvFbhAsohne+cUpIFRfJgyY1gwpWlyOGIvIOB0dTNRMaQP4pmdV6/AT/EnPhFAQx+oRlio
2tUbHcUMIdV9ej299aPG4LS2MbqVCggNhIsmgS69AdYa373CwTlvRUuYDDTWx4vO7cjyhyZ+GtYE
bxelWlUE98e1+Tg7JmoSNmIPp5z5/hHNMMC7odoQErmw6NaSlQZRzF719bnDspAqe/z/eRLTD4Xh
GB+v+h2oItVRUZyqLTMsuPbKQg2M9VmXNPx84XoRoitJcoFXydVZS2WYgodfOKYTrYpNoPTG3heN
hAelXyuIT1d8JZ+8hAHgYdklTUPmhdnFO1ZFJKh0lYj2+qcPMQ8wnd23KKonxrTslRkPezEp00Qy
JFLqqjW/s0H8nzW3FPXV3bBy1w0/8OmDfUr0jWASLFnGBJqvmqBs3wLwK+BM0y3JOLzuygaNQyyB
XnrZTiArKb+vsMuSACajrqk3BTTTtPe459iv1AJxUjxRdid5zmM4GRhHbWQVCYS9DWFqXxSqsJfi
VUDDfJ/oLSSCfnBPcFHiI6RfqEntUjLSZ8xVmulVqYqubcRSBJfSxi6grS7GQIS9IoiE7C2gIDfT
ggP47IoNGtwwI1o+0CWANJuf01PU4aL0lAldae3xbmP5vaADo/HP7zf9e8ttZYa+/je1O0OXP2FU
zFIAsTsfSbiFbIvy1rtpm6nZf4epVZXwN91TSUWL7U250aKYuKbtu0NGeQt8NY9oUada9IDHo1vC
inZzp1eo3JzGDGyAxqD/duAcJBB60pXQPOaTVYGGzs8kRu5HNLJVGKS7Gsu8dMD6ojYkoInOUaZP
XBrmWcPiAze1vvwNoKfjUEKZNnOXa/quVFe6LLUg3CJhKIPJtDWVawMP3eWmc+XTlfxtSfJyK7Kj
j8Mr+wF4eR20TUMCuGk2Xa+4KfhbeFg6OBprDwgf+QwExkdcqj3p+qqF9w8o7g0e0Tu0gt2TOf4a
sdtwTIWOv56E9o+NJ6IPKzDTlfK64Usm/XPcd7432KWLlp3V0Eb82CxFmZBx0JoLolWYTP4A3w3d
zwUdHII59WP8c3dA3tYwmnnYkQA98TxixWPVnPKKJGOZXQzia1nrsB1wozaZdnBir8fS3tBvWIh0
hO0NxcHhtcaqth5XTunGmHMTx/agLJSk5A27aoanoz854M098eLM0l2zfYo/L/Mnmc995lo0YvWl
QJKqj/gts/HzZl5kNHvni0IdHXPRvLbqULXp8fRnNEc6zHFYKfJajOKqv6/9GzszVVR9D3avze3i
XDBX2a5vbTTgR2pO/T3M0ELOwAt9EPF8cWLC2auoforB4mHHGQuLtVP9hGjSot7gBwQBmCIOsXRl
VrmrPcFqM0Qg9j/xHJYmFg84Lhl97Vpf5AqnEz3zcJUNhtwg4tkIEww+5Bs8wBzy8jRL1Zsch/89
eL/X3gxU9lk3QIHg9z3I5pTglRlu6TieK1gX3rOh4Qn8zqZzOrE0AF/yt6gTvtG0LLQ8SyVFz3ht
B/jv83ENNulzzoX6KUnC6Tqvxx1cZkR35hns1ZdoZ7lYay0QQrzXlgmEqGn8AGVYv4CCyM7JZiuq
vUJ6wRK4cYhgyH72qu/QofiDVeB36LeXhIBSzssK4S8uG6+QKDXO9CdReo9HTr2gXNLOdH6lUVNU
7IW5jxJFBoj/LqFnkC0nLqUTJzU7V1CZWHuql0Xc+B60WgaA5Vf944oatHBR6kautz1E/OfO1QQD
ULDnky9rLk04lsfe9AmiVL923uV/FTK0WONVY//D3BaBdaiLfKl87ee5VarvWZ1R1Rh9K3D2tM7p
nT+VBesYlvsCp8FCaOo1PkYws7bytpPFPQYzM6csUGbi9wAxkurJ9zmMCNYUcUseEZORr9XTi07G
CJDUlVQosTXFireJ5IxCJb7f+yQrxfurB31QUbD4si3Frd+BMcIMCa4FQZyM+wiA2dGPLqZo86/N
oYqKfMocenGTj44CIhmGG1GViJpZPsASC2qIO5tElPlBWo0kVXqaTZHaS80d/9H3LYRF1j/TlRdf
pFiGkaPKsVA83i2/azc3G3OLhYm76OXlLAZMzrMg3/uM7On4nY+XtmtFqMA8KQySwrhflQl4FkOA
clkad1lnVOXm4ZybFnJmkr5+9CnAJFBdpgSMpM/kltUCHatjKhuaTWZwkC1u6JLstIjpAUZTLZdo
VHHBs1/FLj7RmYX6uCj4mB+j65ELyBImlb3F9CMDc//f3GqZ5rSBjilOkklc3a6Wl6+Fm3kVL0lz
ooaD03rGUJG4DryqEv14OHWUBzJskmEa7BJYOvDsCgqMrJArP3fCyYI/fakypkx6fdfnFUp3TlPy
VmMisYRfgq/QyGoWpmQsuvoqFxGG9qMwIYULbzpAo2OEkBVe6gGyheRNxzZtJwSzdpm46v1wzYqf
LSE8ethYd+p0guiSvsNCe/4onWSXyMSKiqYivYLRMi+dBCHVT6uYnnl7OPAJ5lBuW1J8TL7v/L/q
rVBZMWGN7grarQ9PmxA6YG0lXEqwnAKfzhdUqjBXcx0r+sbY3R3/YfPudjNRF0y8xH9vX9ODR+EU
4ZTL9oMU5ibBZSrhktuiFFil/EaLFkHvH+ouUHZF7faJK6jndhSvATxXkgIdiSpOP4vjk04c12j7
KeGSbV4kjyHB0yAEBTx+95srvXwRld4WTqfCoj/rWjEvC8Y1B7EE9ossGZnSCQTy+T3wCBZcumKr
GjquIhe59IHZ/Cg2wdUP3OGajwWzPqTJryJHOh04zxbZTlK0JEOKldR6l1Gn++R03M48e/Yo7h9G
MbRAj6pL7ZerJBkgvZZrdwVsmm2CUyOZzt30JrJvJeS2x26bWKYbLajfb+DJh03CItMDUfWue8Fr
2XOlCo+FqnnYQwciTJRdym1/mGT8wvy1e2pU7//xCbyp/L7lFckdV/PdSJc0JfqhcdeJnZw93PtJ
ojA3m/y0vx0UFhaYh0F/F65wbzNDUgTC/4STKH3Y1Ol8orkKajprQuV1Xc3xNe9JQKNjLKo2y7lY
Ag6JwMYW/CWOvxPzcTrAlY5g0QpaMP+R70CBB9zKXGzdpyeBQ08mNInRyvtgrgQ/Ki3IjvGf4YtW
afIuxOwvan6R+90BSf2zD6YTskAtA4/hbzBtfa/1F2j/F7Tnl+7gdTBA2DVSqsvJFMK7ueMW1CJM
avwKHXv/j0GLkMj6LntwI4H8dMs2PaGKdjgpCIl1O5uAviDnzMk0xDKRpdiPBtJEpo1ztKCXndvk
mwW6EYimEtQxw1gRK9KjS4lhLdbhZnRMZoTaG6jMuITC3wqKIiHApS+0B4D3bYolAM+d51vvc85N
t3XunPD+AGafk85U4GDk6+bYK5UPkwow4qdx63riB/IWk3U8ds8XO8NX0u/ajzrJ3f5Giud4L75r
/yVtqEUzxBYs0cmfxdjMiHdSMf5a+olLZAoPh3gKwAq6VR5GyijrJcTF/YIMMjkIAmnsvNPW9N22
VMJ4qU0qkgCf5V5Ypwn9fdg2A8ju330FW6PBlRCrilOCBYKnIyJExQNzSHT3OMzZ2I4FmI5DtEGE
52xKE0Elri1myJYK5xykkMkDn1Ec2Il0Hc+hP0f9p4Bz+NLEogy/98m78JFQMKjS5jk250LpvUBh
CRd968t87do3CCta3BS8hfAhZRuMFIAHemzd17NN1RFXgxfB2r8Luvlvyu2koHEm4QHe6ixUB8Xw
CVIdA8mNfTQjlW1hjDtDrZRyznnjvut6EZ2VNhqx/sKlaykDuSH8t7Xgo0PSSoizyCw3uqnvutRr
0fHsrWwWLj53Ol1MY2KR/ETBQok7UMrnuFHN+9t6qHDFEoPpaee9PGPYgsjP4E7rcAhj1lotXjSe
U9/TE1+PQMiosp9UJv+f/Kvs5AR4d3LqCQejS7FwqtGRzyQg/l5v4XPXzX5iDk55dxbk3cWHVLkI
KNCmlpEJKo+jpGgqfxUYUFCyK4LFD34RmaSg2xYuCDrw5C4Mmf/CvMsbmSxhZqt9d40+i7G+a4EX
+xW7yPJwRYSbqIst/gCREwwiOYAg2pv5fG5ORcux1oK3OBg+1gFIIWQrV0fZQgOIO49mFedOPs64
frPwYhc3MZ/HvIlqshBuiT+pC4jnGKoNspfcuPFryZycV4oxO3C1UR+cvwQhDjncnGbvn6Dl46oG
0I5plIFTe+xC2cfse1WwCRo0kNXdWmHdhjEBAUSNi2Ba2ZUtQLvBbhFeiFriL2ZaNqvhkPgMx0vs
T6D2m8O7UocJjJ2I2zcAloxfdJYazDW5eYEisRqbnQojKNO/s9IeqEGa4pB6X3VDtCmT+Vr5SJRZ
UwhhEeZon2AEokEkzB2mw7+jPZ037HF701TAuTv3rEnaEhZ2AJ6sroayYTCa3l/MlrB5qeCILv6z
zfffgfh20tL5A86LC6RXFYQXkuOHYxVkPOg/ruS1tNZO0BpLVNxoNdqGzzFNAsVLVJFCqTgbL0Kg
P63PqhJCsj7MzyCs1TG/rNMkwtQVzeWwdfg+dACbbwnPOicZnz+oBshLpDsI2NoSDfMcIQpVRCSA
qfUQLI3Kn/CKNobmS51Wrtvs29APogVPkPDIfjJtx+KLxGxolcW/P81MlNN5bOW1tMwaEoqHx4mQ
BkfZ5sQ+eB0iBF+aDAObfC7rqNNyItur0zNOou/0KPkp82S+WIhR5L/2vVk1yP8bkPxoZ8DTXJfA
7QxB3wMmkZwYg//qWBaS1kI0vF/fNnPzNWlxMmzIHHcCv3H1hDh2LZ/zRW9t/obzmxThKd76jHZl
54l45P2pCuh4sI26Mz1kzYC8fTXFr4qy7uP2zg3p2wDNbJZGRnm5Kc6aMn8U80i2mfDQWbkVXQY+
D4250YcX0GMIcbWtS+S7orCPkLqDL6S6pVgDkgCD7Zlh6+Q8TH9R1okReMufzcbglSM8sC1LARtd
UINjA9FxwgEj3uOQSwPH3xilk51kThahVDdjY54iUXR8AmpONUwZo/WSL0ANZRrAFcYuVDyt7Ty+
JaUF3O/t2JYWs554klnljOXsG1BdRXibTLM/gjnu/BQe76CoOzK6ppyylIX6V3iBPaGxktIb813d
8eOz0jOKFaBrg5JBAN9Fg87N+RNZm669CrmgDaw1yYjEn4n5Lk73qA+frnhSQkbjmHQPyT8YbNfh
3IXXfvInm71G69cQWrHLoymxSNHMhYhMePqLp0c1WEHWEHXCTrfeVdYEV8+PYu/aM2g8Lj019ecE
LhWS2cv9EK5kZYpWjcx5ZedegXOWS5QyNnZvRuEUXGLgIwB3EDojFVqWzWKiWPdvsuxPExfF944s
x7e/4V+DzqCS14SNpKMQoxklI8u2Lp0yaVHMgaQoWzVxB5muEPZR4MTwL0Kd25unusCSMSOxl7IA
GK69EzF2a8Hns6qznlxIhIoxLhgNck1cFvkvDPl/O6xno82LObUQTpagXeITTAuuYfgl/aj5VSjm
LZxpvS2smc3UdBhHQcNA5YxVRS5EApbS/TQRvl0LPCHiWQ0PdtGcYeoYUISTrBQWd+8Q1KnJOgb7
9o+Q7aSihYSXthZoVFu/nCXvrS8gpK6zBF/UPKTh3BOMh7cZlVu3uc1RfeF84xuMnZb5isvytJW/
IY9Utb1rqBvMqOn8WNsvvsSTvcUWDQDl23RLzPwhkN7+dHcdb2UUeGc9nqNfANwNhcxYZ2VZ1I2Z
3Gvo16MRdXEJGmpHvw44asS4KRX5YwZq3grRnlgYWna023KgL3E9QPCzMSKgpfvpONJgthh3XgqQ
E8PKKHNXIuywPxmKlbXZiJS02SW1Xl1YmgHnMWn7N6ZLAUb7SJroO1+xerNKB5sObxpHmySClOTg
k6V9fNH/Zyg32T5dEwkTzuOKtki5wH7A5yCjmrnGzMZ5lFju77hnvp8Qd7bd64vAND/Z6rsYPAko
k/iRK04r/LTeE8ZLnT400P6mO5s8Mxu9OiZjafUjXzLcct3+0CXqTb9J9bUnE3Vb4K28A9+861bq
MR6cSjZedzhcC/GB3qYpHZU/kEg/kdAzLX5tYUp2PSZKWPdrA0Dd6tmM676o+mzaV/UIYGmLQFdI
mzHhXp7728my5sRiNkU0MgRNt6Wt/UYUZyQXpozogX4gqqkyj80LAIJEqEbk50i+y5B+Dv6KIC91
8mtGEA+KKIgxVtfoin9T1zpHDmvtRZnNFpa/9I8Br02sBWYKUC9moan+QrOk/3XWg0RmAsgoGp3Y
GI2tEy8wriI4rX33+RueKnk6eGH+5RT/jmjRPUB9vGqMnBYHpD66DcaShe8j7eUUp6S4H+6Hm6xp
odTfJXI2Kc1yb5JKl4D6V5Pe/2IrfpoFt92iiTrJj+ADl3DtXvybUlt94pvFWQkhGppb361jRw9Z
9hv3l9KWPiqpuCtw/bph2L1M0sSpC+YipFhZ0kxPTmSsBpl2VnDWNxkvFP6ob8iklU1r+zCkgQzx
dAWc3LrOlFv4mBJdTMk6idYYyvo7WfCLfpdA3X1Yn8CGlUHEIAwSmZFTdA+7dylq65aQjRA6fnSN
TtcTxVm/ARVrP140dWsN3m2vWf389NDBbsv/VK0MPaM/2V5w/9rVP1wh8iNJA3goaW3qiAo6a2ik
QW15j4xybYrwk8dj6e3UVUJ2ZWU5SD7n3CPQeX/nlWFRAuXsPDEtI0kkbvMwkV/33RsNgPqCTao6
3BJtfuFwDDHAgp0IBZPQIeJbG7xSO24zpYKccxQGVziXN1jcVxTUimvCfSk+lu5jraHY1ANGWiHk
kJVJFpwXNdyqwQo9INln/yLxdbUpFBdAv7z3UC0iDQrB3J3z2P8n4575T2R48xxHEhhDo09AnfNs
v9MdyAm7cftHa/ipfWTCwRPBHsyNK8RqxeKFYGek+kw4X53Lrp/I7wFHhR9eXqeDOsCGg/9I84Z2
O1BOHcbUPG7AaTT+Bt8G2XYeT8aVslTrBpKc8w/72X2xBPh3/2GE7PX/0FfdQwA6W96R8NMF0IcO
CrfYMX4TvhwH3iGOyY2hokCOj6yBw+GqrNMgGZ2G5Rf37x5IUH9vnVmRvEQy5YhYepSyCknsTvzH
9/sYyDCslxCJRFU1+b/sXcBJEfYhl9uTFv0DKHN7vXPf1JCICTcWNaI9113iyzTI8Btdrnz89Ikf
gF2O80o/SOrQ6fp8AZl66bYLP4MgldnchmOITND849r1mxfD6k4ZDdSPOb73hDk/Qa2b7Px7kOYY
TgtusJr8PwkPoHCb3oZ/q8kKi7T/t02L39ZPhBK1QmYQIyLii/d43ybnkTQD5SAqdNKsf7hCO629
wiwoDFEJeihVKihWbrt1BDU3jwMUV3uz3AO1jIit9JzuPzZGLcBouGGuGOCAEDLHq8qNNXKUe6wj
y1Mv+cuAQTVYeHn0OnnotW71os1UBdkyJzGF1GIN0UGGp25cVxsIHoc2WxNl59m3VbbuoTe7z4uD
F69gpMiVP5ACYrdsUI9AV21d9Z1rAOM2//WFOyVnKb6s4NIa2BS3oFh3SVlKw1wkrh+fsKx8uwK9
9XO+IUjtoK6YuWc+6udMrCtVgFvf4xFiGJdvk1NnRqZ35160FeNw53i3E4F2hNXsOa+B67Zggv/b
LpKGmDq32oe8g0JC4aNeae5ad3nMGI7UuubQP7aPOT20vxsCBckGX+71cpFs757inQ5P+b2X0D1T
yjYS4I4X8oqGe45pBKYyeOxrBHCF3RPy3ywYIChMpd3S6IySoBMf9Et1JhSQTNID+PgA3xMN4CrY
uMzDzmMjQIKEm4JObAtsDwW/g4Z38H7Wi5L8H+FH1g+GUz/L5YmFpAZkaRKKWYnX5A4YM3MoNetx
H9x8XpdB5T1vK+O6hSvjALnb1UrrrvQ9/6r1tXNFUL5cEpPzJlCSlFCDcKAnHMyJz6DUimRpj/q2
XuarNmNtZFeiVAiszokgRm0YfHd8Gdf+p7ujiCT9lSQQnm00xbRIDiUwdRPASzKuOAgr8v5fpnJc
pr/HQry8oeJei1Jjd6qATEzy8gX6OVKtB2kIDf8UB1yqAdGuaHtn8ypyJk6EGxkoPP6pL/2NdmN/
vjqNM6DoHI289jj0tq1Xz14oHlAy5vvdKIMYca+dDIy37rwJj2z9Onz2x8cJBBE3ZrwVknrrXZ9p
11n9bMKbg2md/bDdZpgtF2xkI/cVYLj0G700BtLYaZRESMIJ2Q/N1aCSAP1+KB0UgTwvXS9H+6+Q
U7yhz1M/+4j5JSVc/typYIJD9Mrox0er9xUUaQE0xsGCMxklAvFeLufgcwEhRENZsz6JnXIDLalS
X5QO4F4XBwSNCDYjLD/XnDgC+mmG5i6JV6ytuC+seyp/+cIu2L2FpeNC2Rhg/RPVY2mHWOrkflFY
P2uUZawpGfx/3sRWvvUA1UeeU/Eh20Xqq590EBVJk3O60U37Bd2yZHFJ5NzQjqD1oduVwYI0i1kY
yOc2ZXkj4d9phfEr74F1QtHGFFooo7IgUvdHxTJpAjUcbsh6uCe0Rk2B5yPeEJZdA5sbFFrET8mt
18fe1MeApTy6KT/Hj6rOKqYAw9fG0hd5vYzDmEZB8VU+GOkdE7g2gsVfXexQFhT9iEu9y5f/la6n
JzKU/EbTu6OMYsyii0XQHw+nGszdyAmydSqooXj5ZFf1ITYJ1oX4/G6ExRW60hamRDyE0xz9/Lac
1vuB5RwsLZF1Ne0gFHKuRlKo2dxCvAqZd7er+rNEIUN1AmFo4YU9atwBe0kXvcC61sw8ahiA9wjv
ZHUVJR2/AH8Bym4z1dP2EHvWNFHtmRVeCeMQapxo0FQqAwbvcoB/ZqyKHiD3tYaC8ylJN/Yw6h0k
E/j7lProSju0A3G3D7mYd+vd0Dp1peg72VPvXNxrtt94VjFStrQIaMWa/iwh8pdsbTB4h+kHgk7L
uDeVczutbOl04/GCPfTr3psq1xMePZpCBGBxnaGz/EpLXA27AsThmGu7X/URc59bLEARSij21kc1
oa6IkpHHBrlQj9qSrnks7wdzxIFqKLTO6Zht18W6OarHnAkyFC6o2IE5eALnjr2cBTEI+P2hmjbm
q7fDLg0UojreBHP/Y87rlrwII9ErK8BnB3ftFI8ZhuaoWrleUMolEyA2k7cKMaBXl6ZcA8bIS31s
9MHz23oj77uW4FXTqsRf0nqqEq6QNLjcu0wh7ijtLYnSn1vMcD5RTqXTH6dCY2HIUQ0k4yDLFGUS
aTnZTZAXGfMa0wzGBLyn2XETZCPfHR51QaOQ6W2/FVm2xmpfe2ylLIeeOG3ZE37aZCBbo4FMrR0E
EK7k7Oez4JBlAAOqvR77O15korhA8dqTq/eXgIqzKdjK6VwvqLkKVG7jO+6pn5W0m7gpsLSDF64l
4I1MBrPHknVjops8NHv+UZpo/YdQc0OxBm+FPfm0Czrws7x6Jke/J5MZ4+uzZWx8+7abajJSS1Z1
du/3ThZiYJO6rAXZJnQn19SgSvPHOP3jDDz9Op34eXLfHHvKUHdzSBCu3buc5A1UNYdy1wr2i150
IF0/OcXo2OsKIj2qWCJiOhz7+aONyhwjmQuTM3ETcP1p35e/GrOom7SGdSH0/vJ13FPn7j22FOVY
AVjO39c35QuoH1mDISshqhFaeQYLXKI5CwByR3vMvB8x9n/Tnx/RxjV7u7Z+ft0H7YgpaoFa/Fdh
Jfbh1N0vnrcLTDIciWcdw0ylmZ52co1joueTOtBmBltEYKXuTqDNVEHuZ76iCRdRafyz2mbjZLLN
F3gYQZqbXO4+V8A4MBb5l6fu1/DrPiInG6UMgf4C1509LR1Yr6v5j/gbBCk+ocivqRlvCkxLyhlT
elH8W5/xao2ZAC6hnd2Zv1ofMC6Buu7l8TXvxhGfsMIhQLhDMwvUtw+M/C3Ve8Ln1cgDSc5bRvPs
p3kbyVI8uj/5Pv395J7foIrFLmypwUBZThSsi2bb8uWP4fQXoDCuzZYcWNIZ3l2rfJdIjFsUhWWr
hQdiX/VLstoHIWYqjZMhKJ/bfN0iW0NAnINzfl1zBp3h4nUegM16MekEJp8YMUIiPHE3xuIaBIea
Cl9kwGUNJ+q6z0AOXkyaDlDQcETnVx18pQUBac85uIJUsdGiJoCYJi6kK/woBxPKAjXBDclt4HPM
UiRTWhD2EF2tvMegQ6/PtjayXVMAuYHu0XfkIz8leu2qYYEoq5+0T05sufHUCYNCtSVtkuCSzBva
nGbDi0lDA0gdfOcREgsB9aUcDTxJ6fS3r1BNx1OhqeheF+3gAePqag5mZ3AAkrDP27R1AgzXmzEn
a0uEw1dO3hBQmxooTaf4TmYn/UYNU+sMcKOGwMHouiHdZ4kGCI+ggXUTmjrHvQs2M23KyxzhoGX8
JFDs6oWFPonsJ9/RO9t4eudGckOTXNKy5JZmXdoF1riHkrsfjAdR6j6Ti0rP4b0S6yUEJ+crnUIA
v+e9ebfIpq097zCi7A51iAfCKsHeIV16CAJMFJgy8vf8zERVwzlNzb6YLy6o9Oul0+aZL4f4Bsfd
YzcQfCjQS+zATRNlhtq1/Pt+JfOUKP47SjKGM8GgGC5hfasxNf1exOOBLHDiKkGCcOIuRWMHp/iG
1M82TFti2XBEF4cNXuHbTdoqP+NTqkKOWUhGGfclvzOAZu4yZJQRMRTt4MI/xiHnkdP/mGEZxlg6
6iMd1cIPpHPrjevIg6Yu1xYd1sgp/RjEiFkugs/lrGDmvWqRmYn7qF420NhMwTJKIL6WBv2ZNgCD
Hwo+hObRZyVBMcC03nOtHjQ3RyZgoRx8qS4Hp3Tao7ypjww60yJrWurpGKF5nO8mZSHFs5IPPS24
gtJQgrIZRQTsAY1yGivj2kDTXLXwgaHeBUhbZk9eRnvJg5rDhABR3cCdy7tWwisyXmYR4sdiwDsa
xtcsglo9QgIwdf28ofZ4cPXSDu8ZOtBCcRD1Zmp4gd7huHE2e080KJ18RKYOWGHoggTS5LxrTdBv
SoRbgOkOauO2JiHK79CuZQfZqpBXHz3mW73cmvE3SVFWlL9V9Zklkp8MTLTzJufRvsjMIiw9n/p0
o3YZbnm7EEVTJhVa4fcjZjrK5cxjT2wYGvd/B8d3TgR0UfBKuTsPsDlDEKlmB7/vNW/DC7J1cbrX
G91YYKNneBum/48Hf+vY03dspcKqFR1rG5fPGPgqZ8PBpl8AnC/xkwVimrC1jx+ZlU70Nz7z197F
Nhy3BRAN3J/TNeUVqYdjTMInN9NMTj3MBCs8X6CS70lVNMiAJlQuTBLGNcugFfsKT1f7FSP+iQad
yMs4+CpZdblkssw6GE3HaeRKVARWlp4njKxZ2EbrQ98z6YEssMZc3jerK66k6shmFX7OWI9fejUt
LPY6PaM4vZpYYemzv/ko8wQ/rab5muQlf8QM7MSLKZS5keO8XEme5R8IIFhG4MxDyc+SALCkXvI+
ImeWovWVUYQDLd1QJs2z9gf9JKbpmFSwEW6bUdnFcF1IPPro87JU37mnK9jv84tBhpgMuadvyMJN
bFRr9sPbBTd6qBDkAmL17wEnJKknQjAKevgWhVtAN1SYkaUp1HovzgYnDBcMmZuRIEDiMv9gNVJq
q7XE6ZTlmJEQ8dThpA67EsxyN9OesFBBk5LKfG3ybVUhEp/q/seSROu1CqVUpBxdH//CjwLsDWy5
0Jk198543UN2is7FvScglyS/X5FFmosDWW4dyRlPa8b0i66j6/Pv0lkyXd4F5lMRywDFCZkU0By1
IH26uThcNxMA10Y5uax33BHFpPGHtmg8ErNuBuzGnIbRXZiX0C0CbYN3NgQHuPNDRTO+K12L0hyZ
sjvDGgMmkoTxddo2F/ZXzAiWdMqWRnrOID+jmuZpZqC1XLpoPERYuIVq4t2RpZxvWqn8GwhwWC0v
CXW8VBSHX3T8ESYAh2JmQsKffz8KHC0aKipWwv0xDBMH4Uuy3SdYZwzNGBCkvmA1l3CWiJWS8rYs
tV8CAugZFks7xrpxwdii80FiHlRSSC1mlLMGo0Q1NO8Z4LYYn3S/55b7TNxt5IwUCddZ5U3v7Eu+
UHIVmljqq8M+QAfCP5dVkMDJVdBMnEOTp10P9skkPkdSIUObwQOPqxf+RzHQ+Q1tN1U5CuHqYWUe
2qZMK7AIqr7Ydoj/V6kwomIuXxY/Mv6+NoymOiJmiCy3GReIVGimUO6bisDE/vdxCyZH5RtFG8rt
P+IgLElBmwsuYC0qtgbTm7DG3zrpCcO58Bt8XcIdn+XgeMrJSE+f0otvCKqDdvkiOJrhJkMIPMjE
qdSZTsk2104mXtZiPu4ypDl9zMi9qfxsz4ImDwLSItzqviidoblebrCg2QnbZu0dLKr/JPWXI0T0
EfIYUOavXBDr3LW/y6OBwPKAzZ0dV/oeIjF1nfI5/B1FZqhsI+r7OelPh8Q1ZDYmNvfbWpRFalC3
5H6wBZDyZA9QsDrJu4vXSE7nng6ZT+GgSd/MGkdaFkpTpAPkLXpPHpLGxivziq0/dPRZRdH6yhMI
5QOgaachYuuGPs62TXxwDW7k0AG4xOkoTNaxI4bfdMRssX61IldeAdCIX7p7suk2Zadi+YeXpnJo
rWeP6Gzx+AtmaW1r2dGsp0CKCTDLj2GNHZEdPQ4pyQ+Wngn+DZV5FvJ691MvKLxS9uRbPQxOeKMa
GztE8VvSHWxaMdV6L0sk7t8MJN7l3fQRAh23kqXHxfhP1jsmjwLEbNwaXowcO/UA3vXeNTrJB8pj
+vLf/mTDCiFAvMai0Ibia6ZySOmTEjuZh6BdZFIS3H5n76zioScSh1q1Kfs9Juon39u/mJdiL9RF
BUdaaAOMtrTZl7dFiBcWPSttBC9LChsdcx29UdL3EKNid0HfHlPy0p4EM3nwkFKcsjH9HJCFtSMJ
Vv3x5D4r1cSuw6yS7g3VhxipkBz6skswWejpWa7UgqRt8rVLNmJbhZwhpI+tGXIdSG/5q/uwqPVl
lUrktR/hhRNvTie6cTRl5M3t/70kW8weDrsn5b0eFa1kEYTOHDt2Dyrgt1+7/a7j3Q0QV95HNkiU
M8yqSbP/ayVg2qSu4TwBimBRu2lRzg8+to4tIKPbxWorWKSB/xiWW6vfYlR9dVmZKHaIN7/qpWX/
VPqRzk2/+wm3HamcvGJc0iHm2ouALCi/Inhi5+48a8OWQGiDidad6i3KMwHZD1ymzW0nReenxatI
xv5EHKTkx2s18FELih5hiIQFlrWZmGEV5Ay7J/dC/lbSAuBcZw0+PvZ9UecysjA7XedGlrLn8UHX
R2N0L54TXTnQaghy8/n65gUBnrN2U1LyafsZUtBkM3kqsvCr0GbTikduzz0K/te/kkcqIrft3ZUQ
cjzAfSymFwi7WjK9bd2p319E8cacTDdTKi+mbygNBTgWZb/A64JJXBYlKxbW5Q16mBc1o/N7Zc2D
Fl+m2fPYtRWBqLv3AFdmuNE1w43wSLBPBHu3+Mf0IAlat94HnXbHncLjRkrs4TGu09/i20RjsMHj
/cvJAenQr6xwZYl2xoT2upqzlUOMofexUClxY+JRfgJ+HJHYSl4k0lU3u8a4eZfXsC8m+Z6c96Pz
yd6s7qbGbAJFG9xSoYsMoMVvqnww8csaeFO8vex2GWJC5WzrrnetJLWRhzk/dwkzATvZ3t6GlPGr
vwtnMMlG7Dh+c/eWSOvgNH4RoNW5e/LblgUUcpPYLI0P29MD43u4dhP9i37tXIbgE/bq69/+db2w
4V080IAvdywNtnX4wZ2vOtdaH8KCcYnS2biuxSm981nXWALkpJ1dv12VIz6wkAkjvafRAKmI3b8l
gvb5OS4Is1sdgXmH31g1hk3kQ7BHCnq4QBruu41T0EPRHcPvMgUr+fQPsRhjQF/QwslibHYzCnEs
C6yNVVpdvyMpb+PA1hNglVuH5pcj+IlFZgH0sxSeja4yA4iTxxBQwrkXPJ4CcygmJgMV3HLQeF1h
OF6hM3URzmxpBP1ArPlpLDEDUO/s4Iz9/surRwSG8ZQn/nh13U80DZqnBAuXqKQu5Kt3CmMQeEyt
UTeVKh1qKRTR1YFZNsq0ZQ6yHOKA6VNnQ4lfrE9KtD+G987gLQRDJldjsnuKn48dqAlRIY1Psv6o
+ML5JhDiM0LF8BveGXnZ5mGviMm4EmYKW4Tu3hgcEg5BK98HdDfzKjH0vXkpRUn4y94WM48K9Qhb
hS34ksg30bktVoIhzn1oTAxVoLoUHRnBX8Uav6JIBV2fFBRfo8wxgkKZI3jhTLgG1n8QQtGoqdWL
YGfrmBDuej/vBMdCxIYLcYh7E0KWrLRZTGe7eLowJ0TOk6Iwx8Kr90T9LXTbSMhsHo9P1Rfpz8tw
gzBx1Tp3Tm7sgm4JjZp0ihPenEKvHiXhZbCSmHWrrKvsvzRMQUtqO3RMrciVobUZ5kWURWWr5+sQ
7v2nhzOX4JzotWDdTL3y0M8s4bVanRu0xGrekIMv1vaCEpV3OuwdQhIKJ4uFxIXLGvm3qBesFTV4
zb//lcDEl0Ha0uO1TyCri8lQTJUJsrsHt+lVfdORVacOvyPT/7XZRH0cx+O5os44DgSqvC9PKLBL
lavnBvWF1ipugZtuaA5pMxEBtoTsUSwiHX84eG0tPnbbOBL3vah32MwOA/w9MCLo1AB3b7Yey6XG
hikJKQePeZqSYC+F9BwNAWy0iC3XORewFBg2r+0A+XbTVwKqJqJnq+RqcAGouzMf3IJE5uLzj8Jf
h6515JsZSgZPWJOuCddi3T7lWN5M8H6ZeJ4PQg4DdUgom9fPKbuUy0hzVfsNk8NRXQZofC35f6qM
tdhAZHT2q4/GrWXNujN9urLkIadSEApOD++Ww7DoldBCRVnDkoLzSxhPasXLZ7eI+AiiScNmxuRT
lG8mf4JnyoV0qQMiepNInkQi0I1viJdPtjIMfLRld+l+1JpctxiGiCR78uhrXZpI1BKOJmNHPrr/
IFk/XplrTT7NmznT+dLnBZwA7lBXiZ2QmOlkYQOiqVsx5qcxsO2C8zRZvAFFtt5IgaXARzx8JQsX
UxlnlniZlFlMi8qm521fqMXm7nhofVY9/wuZDmgRjl/GHEoMDpg3jmEutHyzhKwSVdRCijWJIbZC
hHfkK9Y/0aaIbO+rJiqJsT8f+tNPyPBT6AODoX0hWBZUd5fVNNskFJKHFY3LdFEQHRdxYYNWaVJq
D70HSURgAIiPsYsmcmfD0S4CrNqB1pVKt24QflKrujjKgRCYpB/Nw3MTq7+yAt7sEWayN4EQQNB3
wJYZXQgLyn1faZNN6Epl+ZVmZrgIaakvGDiZqsg27WhDpHT6JpYqZo3rAOZt3cyNhAkYZ1lkSf2d
GlRol4RYC98bLU+Q0zj/v58BuIZZFTbSg7Elzc9sL5itJjrBOXFOE/iqrR+w14EPLrifMvoxYlsz
peGqxPeRwpCUHz2lcz49R7N8bcubGS3c8shP4+dwCtcxxmlna5X8/akQpxvHGRFxABVP48i7vs9m
w/YaLEBtXKNWavXMpe5vGOeslOTK1zbseWRA2UQ+FcugsFVZ8CQehyFO5eJdWWL8xgUOO6381SqY
n6bU9j15uvELnaR4yG2cjdCtb3nWx8QRBmhTTuFar1fyjVd45LOBKS+QLp6MjLmeH879ZXpdxhKM
bbTLNdqLTbnmyFbVDY3rT+CFNAVpghohim3+RRMOaSYsPVvZPNOYM7tdxhYcgL+y4TKkLa/N2Na4
SjS1L5Mzp8cKEyFiTSLEZptFQMr/NRvp+3n2Q3+05k4YeK+oCcWaiwqFi3zvMDbdmIWre6ETTxx2
YnCL9ZZUe6b0KRL5TPPHswrZBZRZQjmhCUrp0dQuWf+1KZEvGd+AaArylP65QYiKx3tIzaS62Ann
Vs8VhxqVE7NTujPQzAg9Y36cTg/Yaxx41bT5GfT1FopDRmSk6AdXWiKcXJTxzi10/YsxK1tMg6Yu
JEZDDoXRbts6nj2pHZv2oDVjqzilW9pKFqGzLPGPJxRC/m9pUuWXqzNOH6zTsEpMUumKrIxO5YED
G+Ai/S0b+1b+Ys+mTHlHa6rBTocWYEnDjng7NGj3YN8i7DNmb8xTEaTgBRu3tlt0YIWSMvEKlH/f
2+2/caJM8XADkP9HDns8NKYcmr89IE7uYO+1RSM1I2rqOlYDYwOx+srQcHHwYaCqX3zmDOWHsw8C
x3vCDE1t1CW9NdSfzHMeYy44wjia1g02QtOfNdD25gRSAw+HeJ1hma/D/7JFyfAUUPkzHNQFJ1gl
188WMzi3d3pASo952uDu92Hjv4+msiZB9G57j30MPRMug9PfVHqFV5NnjlZO+pU6wNHV48FSlEPo
z/L5L0Y5WYQ4YJq2F63C6CqhBPHAcP3MptU55kd/u3G8oPB118sIkhMuiG1kyI8rdK5taESCOqM9
je3Zjsf9ynssegeWulf/TZEBwpjiWk5aUdBvnj4bFKk/d6WcHUA1j0k/bisnMAV/40ZMIeZYRQPf
x5zNaP75O1OjLy6iKwPrZy+b1mUwP+eI+yJJEFZvOOkDFEgOO9faWzhJEv/c3Cr+uoU3SblpLMtw
shErRM3aoct51HbG1W/m4ZNxHN/KqmYWWuon1uDoDvzD6b5RkshKLHO88NCctmITIpdJcsnIBiKs
vboPCrumrvREc2ArbHZTNMCO0xlnEvFLIcGgJlxg7vkzi5btZG0P2yRyqkzOWj6/rkKn48fEMdmF
0neXFUUkfmD4oh+KAd+1iE+8p7I6njcomSgDkOpH+d6ehc39+fj/9Sz6NKm5KuDZJldRtDXmTN2s
AWiVJk/45JWvD2IEo/dGmvT/0OaNkBikxd/jKiTSD7gu4YGKoVKpwpOrj6g4d/QUXyms9hKnjji5
95Wo0r3ZfsPZxGrqyiCMWhWT7jlsxW4pGpGlmQyGUNmo4xUkDHGJpGjBGSKHMXOH3rTY7ONQMzEE
6la8jHLe3mD7ErIdHVZKMclxt/hhwGTALG3mgYj0PTDqmzJ056Uwke7FtiTXrJ8bdpEWCOWdnPef
E8i5IFtWeeeXA97PgcPXCWEUWTNnN/ZikN4nVlOq9iq9Khm56y+JSkTPl9Uj/ldplZyl3E5Hn/NJ
G/z9k5wU28Rq9+9+hfqWeYgI656jJ0CNzaDbYqIM9ogUQ+qkV3gIG7WrTCZvXzV30gypeekgT1rU
jR7+IDGXaNtOanx7jykzqWcA3sqNtG1Iz5fnzAtVRelKad6jxPLwrcHlpul642SZsciOkJElZKA/
1jEMMmudZzQ7YTIbggVoLxYDY6+ZUuSmVf1b3Lpigm1wjpdBFD1d6Fo4t1Iu1Xq/ncsX92zNh1dq
PK44NdtEi2a9sXRuJQYnu7uHlKRR2k9IeBoKKaxwpJbAvbz7D/Jx5HC5ce2zeDKRkXaOK2hG1cy5
s09CCghuqklh5grvmzE6Eaoi0WJIBIbmXbYS5Lo4vQMZIeKT33NAV/JOKt50kP5AVGbwvIJxTTNO
Fsbvr1hEkr31HHYvCRkYL8P1dbwV9gGGqozU878YF0oJm42glOsNO/rTJ3sCcCLe+H8HTHOKcTdS
+Q9xj8RV8oO4mQkAhSvseJGgJrTt/iosn6SYKk7Z8uYZz1BTzu3IXHFM/LtzgSLG/6TdYM+Oe2zt
uGxhHZYgb6Fjy0hDMRfrPDKZNA/ZEx2Z+BYyd6bdecwxcjq7CVGs0GR3VPI3rTYy4DsN7B+9RzOg
3jxJIDctbiGhJz3iP665CRuJwB3s4IPj/A7TlLosUh9tc7LxED6q2yDK+PCuIdfuxuMe9P/M6ApR
f8FbcE2Xa5AP8pRj6QinH33rcUcJnT8+kQ5+7excb5U0fklQtMlInUEg6zslSlhdmZpk8l1N3ZSa
xFbErglG2XAjbVRNm4ZdhJunwbGbTOy693Ym7h+jXe1OZbl51TgYzQdA5k0MIaFJG2aGZk23UPs6
IRB7l5GaiFnqgBbAd6AsOkYozOdmQ518p2SynLNKPI/tDcrBAVsz7Pbh+MdwCF2r9wDSvJI0iC/2
xPgMKe8ak9n4ARlOzPbPo85isJvjN34YNC7e6LyoD+0Oxm4J0fqqsj2JJX1PwyqAgyBiCMw+mreM
kN3oWNpOfm8tVYEKUKveQ388RvKrjLUd41nJMDjQ931Si7OQAHEnKbXFlRChGoY5x1SIS34Aat8X
xQWwHqJzDJ8vihnT58rGLCyZTaWYnPaD9p+GmUXMS18pMK7viecEDVb6MxjjRR3drThQrpqfNX0B
+U1UZ8VyuEIAtPKj5pm9RLQbGowYBxYVwNnFOyCEaCLgwVTPVN/bUmUy94pnWYC2CtIaIEy5yMDu
rr4eQ0Ng3jw0P7z8T/BOVq4DipT1CLb6myGlrG+mxNNVADt2B/O1CkuY4dtGk6/mNFlKcUqRv5tT
/GBZtpjCgIF8Xs8O17y+vh8L2lQYmZEPuOCIRQw+CLPxl4UXlP53QaVQCR4nG+lOWg+fvIZJVDfR
3YQgsWSI3CXRUMf50Eu3UBd71ZiQibSWGnERIZFGp3zw/unbUv6p539qAH9iq5Qg0jQoqQOmd4Eh
qI0GNoArBjbI9caUAp57ma5ToPTbtvTFav/m2iMPtJbgxUXBj4i48UbGaMECcxHsHNIq5QedgduF
eOnpYICpq/qf5wDz7yfqXhIpt20PpVAZcVxT53S4BYOooIv+8ORXLBQKBd4aLtf/5lXm1+KYtpnW
M3FXmLSIt5CycMKMvRovU+OpzU7f4QrpPp83ss6sd/tz58tlZ6ppEUzVK4ce3tWIAd5knYMlq9ho
AakhwMAvViyxEjTnUm/8WupWYLTO0pwLhfwVCmrP/PmEgf2EBJTD5wfKUYeuNvol/kvvA7UJt+AP
X8nf7kqKQ6ILHimNH+07AO4tG61z5QOQ2bs9iaxqkCY9KF97F62wHF8UPzkg2qTSsZYDti3/QzoL
6n89Gl9YdOl+1R24qSqTIxbUhPAXecPY+ceg8FgTQ9XXCSGwdk4VqvU2WjEwvlK2rFQddjg7SG41
ka+OIwTX2FHPoSDZ39KZy3mnBhoW3zl9b040PfME4RFXK8cpPDqdOMo9CrvSzohZSW/t6bVZenyo
MHN7aCRCyNOlauTrsPrbVk+qIDo6lHke7I8X1NHperz/6LiX8NRPB+PLCYP/ZtskjKMwT8FmwyIk
mUtz9rhqhZs4JpXycaZ2W/1d0b0/1XhxvzQNdV1fUcsII0Uh54Bos3UhBm1SGfqEaR5TizqWyFO5
l5iSebKSPybDnfp2LdZPe9NOIrOzF5+KSbk6dC7ghkQap3qWvLabTXivCFOS79huElrtP7IP1zww
2vBrbHUxCK08shfqA5akUtHlqTKfg2coyOBDkflFuvckE3qaK9scQ0/4wlwcLjpZOX8Nr9G8+Y8e
sT09/NDNWsdrUsWBiFNpd4JmVhzpKLggXgRT1V/ZU6tWmkzr1M9QIyAZweKsOiBwJMwXz/WapkU2
5H5OizKb16xtFWFIHI8kgR8f7c8HYwrfjWh1ohqRb6R9xGlVUUY5DCHYU9bmfE57xt10l2RGD9Ia
UFJvR7Tbfkt7oMY8u2N4s+zvYbuGRhC3CXIV7zCG27p9rJsWAbvXMs+7VlHhvog4y7uMS8AMmudx
YhGsuiIoidEfPqUTPAo8kM/zLEhQmAtM7whRQcVTHqPl/HrLoNPsUG7YPKhT+SmMGzehzBgBnaVH
S5k89DWF+NVS/JUgGiSL53j4gAvIah+gJKnF8sv7ICMfat1wy86DNcm7OEjsH3feqL9pLoO8dmsg
unxEvhbT+vwTt2Eur3fiGHd+aSJ9vPCESbIEj+Rt63kPoiUf/vK/cARI8jz4V5dRw4Xkn9+TE9mx
uaq5tW686U8kxslQ0MDExr4JXKlQm9TdgolxEzuNsuv/f5yhVj9DcYJgXep1Ycoqv9WesiFy6fQX
qlwe0YHhsR9t3DiD5yL/P37t/oYy2jN3af9I+QUok9Kh/pZ7FupgiGdOv7U3bDOtWaowND2EvAbE
NLaxe1GmTRrAg+0zunC7SBQLaFvJYFOjw2qtq4+36jwZznHdorSJVuYlcM4MQ9zC8uek6VL8GYnc
hnZyxsN4XRHvne/WOYCo0cq5WdyhF8gQZkMOVtYY3sLcpKnzLYZdCvt6O9diHtdgPso2XHY2MYYP
ozlJkE28RG/bMUUhZ+vRzoNn0r8+MiBeFoRsZbtcmSVZDnpisJXDmEwmNQ/Q7RiaPkYW4PQ76Fef
oW6/3KgtI9KClBZAQwqvsLHOeLzhLUx4Su0zfKNrNjaGQFLjL+jENKXGWC1bISyAKgJa2ETTnjy6
VR7uDEU4NrOYh6K+1dhpAJPqpxPH0DXPC2bI5rS1h6b6i9Z/obr7gaxURfktc3yW67c2jlz7Ttsq
B7rxq64wmvDOcYaGr0kP4NWu/D8bU1ahW4Oso2OLwhUV/CNa9nehjDMtfsaeZAVMVgueORtNOkD6
/mmxSs4dIyNv/rrQaeE06c4FXudWaqYp2xIlFd//gZF8sU+sIt42J4wZuc9o985Ojv8eos4KOiAN
Ttk/6f2xO2/sq0av0w9PZNp26AYiFLXDLb4xlGZa/AsiMNKGNt/GMWUSVfchQ8hZnfZ+Pu2tGK2S
ret4O9Foa6zlqH1bSyoFuwUyv8EpslFq46u/EUNhxHQ+ngjwsXOGWNm2lrqHWAmqwa2BN0CVCIBv
QIiU8jACrxxOdSdHm+wnYGr0LvtMq+MTLCQUxVtagU3rRP7KsR0T4PO4aFy6hn5LKQ/6xCijI7Tw
mkrlPWscOyI3vNjXs9vkkLFcKoXPHppPPVWOZkA9zE1kdjzSy5G0nHlON+8t9G+tj6Z4HOaMBx/k
HHmcL41+0lzUCtqs67XSIAs5MFC9Bm88ZuYg8pQNWyJFRbFiakqmB/SXEEaNe9uXwWPEtM5FtHtA
9Rc6wZz6PZKGSb6hqci6IstxBCrPAwxyXyX/VBueGP3HxD12zDP0h7xdPHwwAE0JTYWyxTkprl4x
hMS5BT7LHpqkeTWrVhSN++sGupBD1jafUQVmEH53Vy6a2pZ9+xlvfo2OChh2RNURML0BxjyNU27c
f6ifNEuCv9jipERFdoZcDcgBl+UpePycntioPel/2BUVddM6AMxwzTdxDptjF4wKevPIq0ZybzP0
e3it0UWtDn4g2boVNiAKEqY7Mt6O2VVLhdVurYBMV6g05fyAjdZWK92s50qPPGLBhPZ5Pf7EXEhi
dEduxlCR32LnxkrKZzbwGG5J39H/aHp999Z3yUCDTzfipN4HfuXt/RS4lRV1WNO/gAy8mIUgoopU
8k3ihvQfzxczRfhSgZuY6cgvEkZJ7veZkfF3Yh3DzuI9Fm0e4QBuCz5cuq2P+4GX9vFjaOYKYpvU
T+QgyjpLeUqIPh2hATS2GSjQ9Cb74lXscjuylAikd/Y8bzyZ1LqP9sbdLcAfVsD105vp0xpnTpe1
HX0l9dy01uZ829nx5meWQwWtGRdb4DKvCpDc27dsPoNzEydeh+oTJiIK6uy8mx4IXwb62ckZV5do
+nR+qmp/bczRhP6BRgnk2BsMmNM7krmd5gc4sZDp8oXlDuzNmEQWgiaAZI67DxtUvWdyWAO37nFg
k2l4k+84is+wnFYWZlzQ0yrgTo90Mkd9Vtu40KaOOsSmLd4oR1NcoUsoO4n9fzAvbG+Yc0zpPfwJ
FmoSSmAUiO6AmXHxJbidDF5B2esPBbK8PN8CG99kwzcd7HgQIox3co6puEfrFfN5d0ysH09v0/oz
s38kgERbe8VjVRi6JfTeLI5D9eoK6x2B/9Uyas/lQEsqPkNB7icX6kGZncdpceaCOMJz/ciWgrxg
4dj5FHexGfGjqWZKvPE/fOruCxCT+dHuz5WP0kWpOncgkmUIRDQNW9XR/npQHsrf9L2K3JJm6yIE
4se1d2remysnVUgv4EBRDUccxG37ZUJ280o/twIUkcM1ShKUgXj+Yc3duOx9vXs2fiWJv0ygO2iD
KefAGqlc9E5mVhzz7nZzEu0Arpm0gIbTHaWqumkig3CV+0ZuNR8ufujcsdQlg7e4VkpipOBFOSG4
8YhceEOWLVW9FHW5vJY4hxqEQeIKAxJYG7hvkMX30LDoBW2Row1PAucptX0jS/rV9H127SsjllGr
0LNWIQFpce42YAhyNuxzcFLsJ7b/6km1Owp1fXSGqNWMUC1S0HggL6JaEAmq9dSMzmN+JXtH2eTW
atpOiRBujQFU+pXgqktaxFBzXpf0VOROKAtouMKk/4P1pNH+PuiGE3Xli+cjFxHMFuS6P+54OWy9
hbzE5CTrd6cxZ2tEc25pOiAxi+6FWpifo5evofl1hfXKZucCUFy275BxkdOD4dof5IIfFt35V5AQ
TqI0sgyphd9+eDSMn29NB6YHvr7dhCM7gc4W3HIA/8sZ1bFlfc6hPuX+ivY4HS7PktXe9oy85+0C
VR/KVm3tSa1kbj3T2yGdLbTHBhVm780a6DfS8+iviqI1SNz2PLYWGMn5MOAZpoGO0i0IFBWaEjOR
fJEjHeCbMJuF+wjBrXeTD9jZVCiM5Ri3JJS153wbGd9WyAadcUlS2cDQ33TCKRnFmT413HTZxJ0a
zMkQBqfUGv2zT1goWdYSrd0RZ51vVrXYgY//5rdhmlqo9LKgPdMWOvbl76s4kCMpqw36fQkneP1x
8Vbiz0lpnr7oO7Wi00qzLZs7jds2gaV/MWWFoP2BJP9rfwGe21r6QoqoNVtamb/8jZEhq7fLujDK
q4zQ/c+k26uLstJL1AEwR6Z4uWv/n3lcWebcDNQ7JytdNNQmjHPLIV3ZNhVEKwFM/svWD9PEiuVj
NLeMESc9JibudNw0p2vW0eQMfs5uwrB7mu64zO1FbgHtezcQtcmPEqgCoHzJorbbWGiu8BKznhw7
J/270olCpAIhfC+WW/PfvBQbsUCgBPdZEB64+PNoXdIQxPUMqO8oFPvQ7Vq5V/2KrFUQb5kFGfyr
KTLsyHjy4u5HRZzOaFVQ6feGNxfrMDjivbhAhszGQb1CiQH298cHtRBK/BgNWL9ZPuDwMo24NI8u
qqhBTven/Y1dPm9Q7IlhK1oAKiVhiIsBg976mrDS7ujqC8WcTOZX4gWxMnNoC9uwz7WfbJQjjS89
7BkCkYyK6oermXfOtAdD6LSJAbBwe/SpBfdYjR8CBmeO2mk2D8DPgt8YbZgDtcCE0t8VI2i1Qf+h
dsxErniotzrRS8tiM8av7PcDva5N1AT76E2r7ED5jkblSs5fbTSD6sCyVMCN+3z2l6wFjZfDdytR
tsHhC22RWU7kmeQaM5Bxw/KLL/4JSk6opWqufEB/JnM0fL0Cy/VOgENv3xery+23btRASCXhrjlK
uWvU3UlJZJXVLghvrWHHQLKoopiNlXX8BEXFWMmmFw5JGtqGSGvhGic8MVeOpPiUx9RmNkzJkmsW
t0Llmbi/QPp/o+46z2CYL93IMvwoEYyBNz3hEw5nH2u3srFH9I3p4pRycdMogYKBuBHF7ACF869l
Axh+MN6hTJjLWsCFefEAaInujHZ+CYztyrW32tynOuy2trZoh088ydpwWZyoJWt+OuDEBpFXBSnQ
IsmBAMhpCkXXBhOKVMDEV4XXMuQC6dXrqVP+z90n1jhKnaocgeE29t3y0EEuXSDHLYnh7V/9tn5Z
YGSksAhEeDpmYMv4PE1I+zxZnj8GPCT+VKt6OiD7+ziHT9+9lJz+XlJiH0ZgNamCJGUQAwFCCW9k
YhjP3IYJWvJ/MSpzOp35jhFTHsOn1h4HyjS6JboHI3hgNEsgdR7Do/zbLPwHyH2E9w5JwbZ88AeK
s8uKaU6wtWj3LTWer2/ajRAh5UM3DQYf5oHi8jApWffaw+1pq2V2gKqwGI8nK8BihqGRF0zs6XXT
WPoVjawgeNcNuLXX5XybP38tDaboL5XCCALby3Fpf8iqonpfBEIjTUAcVbY604OOV9cYGet7upon
mTSW0domVBEGUzwcGZRdtyQxM+NEeU0hr5r7KxrY585vxdgx09yhyuhaYXjR3gcl8dJ8J5osLkeB
5kHLoVo0F+X2X923pCndDxmISVZQoMLeXkbkBkjhMRAhLiRoom7RHM5dSb2A4dSoEWk9sw3/rLBp
PafqVD37Sw89NwCsGNg2GLVmsestkpFcnQ0RZojgJcxGLfe+aszM830MwYRKO7WU8lhtyYbXw2Ny
/Fm1Iixg4YyDOJ2wafdchZnU0ZQIpC/bBX74RBZgr2D8gWH7Hpsbc7sat4vsOOHBC/vReERDxBoY
Zj+/r+KXfNV8LuFjcmAUXBH1LX1O/GK03XBZQqhUHGho41FeIXE4tTpmRW1oYj37TRufmEQIiud1
3CA40wq3V6opC8dcbPsNU4CifkF6LeUoUc8cQ3cdzED9jnaw8y6NMX4prv+T/1WdcwYn7QOOIdLs
MM3gvLjE60jbWf9JG7J0anyWSvCpBxchkERbLBsbePK1RAL/NF6K1BW+1Q94vGV/dJkDiVCzw55I
q4t3FQHrg75ox1nMBOHLYm+XdfnpLWwcdwnQ25oDEr9ozxZ9VPx1ojgd23gliR9zitB7wR/3fu12
axfIJFCYNJihBenCUhnMBD4l6zanYLgkVxgB+79UWJlJr2gLZ5ap7lICm+lCpKPURNYCuKqEV2hx
PxHYMj4IN3e/F3bPgvngD6CqgTqg+en0p0eMDN5nj9trKOYLpW87Ncu0xadwAAF33iD74WOip8y2
FxD3mCcDiPU6WPSxOnmROXgsB1Ls3s7rkQgLVZzuWlwO/ycvvh6g5veBWoXBLXBi1yVynEPYvLNy
U0iwgmoRSJh9S0kdb39Mxdbe4Vmbi8HxvvLax2484BU0gTYCirCPr99LlIr/ixqVoYroU0dGsSqE
bIHyjl42iEQ1pvHEOfy7ICP6gg8YWWzHg0q6amVeDnCeZB/4EROdBkEuVd1HjnEk4D6yjbWpm1lp
Kc0g/yioHv+v0hn3G5u5Qbqxf66tPkUOcfWmXUc3v3Wg3Bw6oEJZrJmKrfYH2SjucOnSb8S3ak5X
0JGF4JzOQaz4jpmi62Xhr4m5qViZOmCRyP3339M8kHbtRmndjQ/TyddDWnqo5da0IYI0Gsp2QlIP
eFhOL5kHhEidwxWEUJ4dhQgz8rgP0MXLAgrG2nK+mKZ+T0ASX3jSqGimUAJOri8LxetZNk9BrQmZ
pQOLCt+i5oGYucbI07qBfiuuNP+OPTzjQsscncEUQj0r/1w36Jm/o+xDW/j41GknkQ9kXblBHPEx
/LCtzrIp7bMTbLDDqA0tfLPzBkSLDOegKqK53aJnZcwNjTykGeXxXU0EuUbmIQaZN9Mtb2tDEru8
dhzT2K6flTzF4uxnWlov4AKAO4QI/D9XzOA06lKTtKMpmIgtEaShl6qwGd2c3Gm2jk+UB1OKCwuC
qvom90x2Bt3T0LskE9hNwn7vy2G/ik/I9XaK7GJte7W27QAoCIJpKk0I1OT2ATmCIvMc6F71QMbZ
ZKxk/YVCZPFsbzkryIsMmlSTAhE0AvmEpckqdwXlbrx+PlZIzpIt0NA96U/EVrnWtma/u4yjd42b
UlpZnj/C+niJPo60Nvs3w91Ql/Acsg71jX6y6gU/oGRz1dWte8vDQdNChPJoaRjds8tU5xdbC9bB
MDlHGdkYx8sRRbMLuXyz3B6xav2kAPajPA/T+fxx8q40WWmeBe1O+Kgs/ViDbDyV1tUL4xk92VUS
eNpmYNLOQkzmKyOWtxVOALrmCDdz6EMf+OPYWkXETzFhBvldxtYr1WokG5oCUV4BXnhy9YskyQiK
B6OzuUQ5eR7qaCNOHvA8arkHDoqADU5uS9Jt0YtZtbDzR9xSHa4UrE7XMTqsVEhL1zc/72zyMqs+
3gFTraAZ/ldVJlmw+vipTWyvj1gstgon1i2Cw2vZ3Io3Njnp+qQjBgo4benLYLn1bRA9P61CXSkA
GJukY3DVLEMpIWyr2k1bSVTArEheTLxNvzVqV5+YVBxLsZ1SfEsAqkk0IgLC6Kcd7mmNx7G8YjAn
awxShfT8io5t4H/g/4Lz/kJVKfg7MHnLYJRhxoc9E/30Ecf7f3HSZAyXz8Z3CE6xIbAGFt8LUc0w
PE7LHG+xvaZyRLDjxB92bIsBASDmBeZlQ264eENR/yfXs6rIW/RiC8TqBlSMDXXMYOMGmbm4RnAt
/a2f4txt7UhZcoCmkWtWgm3OYN/7lZyBHN8RmegYBWePfFiTRMuQGeR22F3uQWXKQcqHrph/P8Gw
kMYWMan/TStX+XtCRJVcbit9KMxvZndsQXnLBX/+I0Ae+VaGjbc/SnJGJxPyD7GVudLrJbNyTUEr
rfitCwdzd3K9qmUdqxWa0AHXB4+OHCa34YQzybZ7OThN4eL32dA3e1EM9tv7UMIBoYlLNEO+N7YX
92Z7BJqJGRIz6SsfW0fG4M+woYe0qylPkC7I4cJTHptE9rSZmzeOUNZha6Tl/YgohD29qcQUYj4d
0WjBYrSS47cvzKIOixrHNc8YAV1Rvr54Fi6poBqAlGZTRe7qXrbXYr4DJ50FsEf25eC7fPNybh89
Q342oa/wQwhrwkS6imgP9KO0xma6AC5ECqUbMzqUlRQFpSF3StB2KQmo3G2sTK975oQiA1lKrlig
cdLEIF2PSW1pJZtNb4abx5pr40JqkVnOJMaA+kHPKr9udc1kA/8dICudCdlxRyrvTlcWLl7m34HT
3HJAwjUf/a8kFpcb0qtn2ak/qOIGw7e+bkq4O58lXCxjPOz0rzYpzgdNuAy3mrR6RJD7EzmWDxEt
5DxwjdWzFPpFQRdyI3Or/VbXsbRjF0LFmTdvQ+l2ke+eJnFaJTiKSZRUVgvgL54m12W+gR4FKLio
o+IuHX4uuq9RXM5WakROW7pb5of2qoOf0z7jnXZli+CHuBqyZAtQU1IG80MGvTSWP6ulOsLC3NZk
Ujyto2Y4aaIU+hXYRd67Xnv5F8Ipejlzy+weJfwXhP5UR4MBKOwAFdhbJA4Va4xkRlzcmfZhxUEE
ZVNgTX1dW/TBoFPF1qydZEFdNGs+mCuqQgPq4qWmCPdiOw7/5O+gLk3wEGzFZnjuxy9HNSeuECqB
cNxMtoK5h0x4jIIOXtCgVg/Mhdha2J4NT0eUZIpnXr5F66ssSpQTj8a8ZprY2WKcw8VGWu5cU0S7
x/M2er73jvGGTad3DviUSvWPlu9JwGVJTy+/xj9PhAx4jzbwJbrm6POiWNRwD1h9yHqjSLcyITkG
TOAfEo7wKhrSOXkcYYwirPbL6DCCHHtl4xX+MAQYVNItLcpPxgF6oRh1wAUAIvE7FCx1GkQd9nc9
2kTo1uIvKqTXtgTpZ92asd2oeM0jjrI067bGBioU4AKzi6sCq3W2humysehF7VnMUpA4Z93uwRTD
YByUuVhQ+wGXZapR/pjRnt3y/r7G2E94BlAsPUPpB+LbFz4znwW6OEu93t2JNxcagA7Jc6ty72nz
BNMO54qYKNr4o0K8TJej5W6sry+fJ5K/toYcG6EEjbEIUOCcv1QaBTrWk+fv25zZMAdL4DcnPJtj
3CN1HtjA83GT1p5q8u3BWKl9q7/dBb10FcBq89f8hde5HdCHfTcLqvr4UShulY3b5kHVG8pc9uUe
qnFiWuC009md7Zrwm9L5XwM25puhZkvFMb0fWNU93WRDdy5vQyZiOc9tSweqFqY+Om8qjVPJvA3b
nKxdrlY32ztrAqN+TLM1BqopnUi0XWyw9D5+zpQNbPfDm+XDXSdbFNPiTp0LjTl38W2Ee4cJDjLl
mwvlNQxEK/IcqwMCbBUJ0ljBuj4VOimQrih8p2szAkc7FraW2WAtMnoQgg2mGVQHg8kxeNw26b01
0augr7v4cDQEu7nDqmgfK1C9fOX72MbZJSZpqJrQpWbUBf3gaqoqkBtV1tS52o/MaNJDjSYk6p+A
DS2twz06/oyIKiYhPKE1uDw+5JA59xtMQxwcFgYeQNLRd8reqv3+0EiuhHFGxocH+bjC+RmwzpIH
KV+9JuDBq/w+hdwG72LMz8yAYV1sDycI+XA/XHHKhG5QckedC+ATqUleLJwtDUGKZneVRonURxYj
Jyoe4SYFbspOUJdzos0W8HYw6Gc34KNX1XuaXJrlnU1OSE+Op6r1l51OKuOt89EVHo0ROaTJc8Oz
8Azq4rCUmVejXI2gi50Urs2AahMLbFPqRIbi+vSGJxfoxZd4V68AeAAjkokcwumZJ89HUyTJa8Z+
0zX0FKvxdXOvpO9B5mDT7q7kqhBVmGKnumot8R9nIdN6bV1xxsqwpnE8Gx5ZKIv0fM+gDEZUjn7+
iN/6yWgCJAPFmmK0PLYG//L6l8PmtaBexcVt1LctxKsYtaH52EAESDkOREUFnih258NBOIk1+qCe
/+vQjLyrrBugJaok6ikW2EzpuEDfmKmhQy5mGr1PlWuitZrcB6AKV4q0cxQsS2hKWJT3hlIRzcu+
u0vDGofepKUpBNUeDHn9VlzVR5xBY/O5Xw8mYNfmIMza6H8c3kzF2vHVE9dkadWdpYjOoNutFDh2
Zzw5lasFXZ1kYqjg4IeWwVaK+fcmwO7ZNJh1EVkOOhLwLr4BelfzEjtLmN0dmKwJZoBGpxQBasbG
drcGco7ctWYa4l1nr9VdQJyBMkBYDZOQwYMNEiA4pwAFaS93bfFmIytELYTyt+Y29F6by1Q9Srtb
Kt4llOr9eAFUjjsl74G6k7TXIZp/TydueJDLEpXOGFqWgCzR54IL8YEAbBtODWFmb0bcRxiergKA
zHafkeJadYhYKes1q3Niqp7e50NndUFYR5iB40llm6dmqsDEArmu/IRMjUVKq4s0w9wqyqLCQYVC
rjS8RzM5bnKEmvP+I1zEkGbETFVwLY1sSdw0aaCErXQzY7JzEM3DqPniAomf5Zc/a8X7UxnM+VMm
w7oD+b0yc7xvSTGf8fRs2ahR8xBY3TqidW0PNHDghxvDY/zQLMIK931d4KHAJ2DOoMjvTYuQthi/
FN+0O53Y9YipVKGuzudQKFmWISGRTQCtQzBRnyEoKYwszNkU7cXSMtZfUGztPjtycwuXCJf4WQP0
AiCDiC6iP/UwIFkr9Tr+nhNChcI7oRi00E2aCHhNMX2qqSzPyKl/84n3YUAn30EwFmcSIXsVttNE
iPWqhjHGZJ/ZWyLwnVc6X3NAcIhaGpI2BV/IlklREpFBrWMSi+HxKFfuw2TPeKjLhDg7Yb/0qZcS
wwOK2wrYEo/P/vHu5YE1U9MbH7LMsOJAVvN3HpBY30kScUFSNxzc7PB9mvPr5KsxuR/+q/EvDOTC
rw3RSl2SN2D/VzJqat7gDIU2UDErY3UhBC4VvneEyCf8Fr8p3y86hMW9p0F+URyi+/hMZ5RR9pLO
mw3xGDNclsmRMPvCueLV41VG6xU/Cf6jqm0QYsw4vNR3adiNRT96aSPHEMUIg/4Z9ONdfuzZS+s4
FnlZJ1MOsO+13qvxVAwJH6WsjeNAjAoFJgXTpZQi74eNFiKjpsXcKTnq3+nzgeXca42TCIPwbHxx
JgoLR1tGkpXgrLTYvjh8XD4LBNbX7mK6aZJRANB2lklVL0NdNVbpTITjzLTPdSre6saRLR+eo7jF
kdzGtDQJ2/J6WVufq0MA32QwNPSS+IG4MFxpRv61NKHzmzhDKU9xgjoi6ZWWEYuDbeA8ahskUlnL
7nhHFuYy5CNjpusHPXyXHjJ+s2BNBTX8dlm66lRVt0Cp+8hdAegwtBAt8ngS+3Wxv1FMGCUGoNpg
s508Qznksjs8ysaEXcRyBlrqh4QvSPLNMi9IL+Keyjsd61jtMfmlRcFwOb4wB/IhnEP5ruBOnxaP
TIKHjyYXxQSkoUmBDe+pOiw3MmYgyWMe92a5zbFfeVnGYFWXDzy0QdhfWVAQ66VzOTNNmByoy6jN
m0A9rLDROpFiYLcCPQ65eegxgPdb1W0Zt/KLtttoi2SjJOsHJAQ4FosHNFlYTbVFgsr4CIPCMbIE
nlGRzd8SFVb+yf5bgqbdUARKM9JqITt5V4K2WbOQjAZceTJy2METdAFXIxnKti/FLUXJ7ioyHYEI
XIlMceTwnlt9h7VJFAcvX13mfYeE3h/qYYQpUIbKAQ2/19lI5Jlg2Sx0ARB7zSxUgi2/0yXtQq3b
do7yI5GddzG6kAsPZn7r3v/RO3A7AVvTKlb7ZRznx0NGslsVJ2zKxSvaUGzsJlzu+p/6bPZd+Xmw
C7d6V3TVaR/TO7DWOfJGir1IrMsUEUGsynOs2wwT7Vya4U68bpBdoxq+aJrBK0bkVA26y5KPjV/V
kbvQpPHttyT+uoabiwtc8Nhnm2/Clb2R10cyav9ToWApU+i1GUkoStYS3wjAL5Qwf8L2Fp0aPqPx
vqgbPw+4dHZYXNM2f0VlMsbZkZtZrfYMewLIvqL+UGGdoeFpJr6oVuscMZlhu3T11EAQOWK+JARM
EhzC7vrXdHSIdZwvF27p2W/wxqiN4VbktSBb0vDMS3PbTBbhFbbeEdwi+QIzsDRNKSpIHvAw+5l9
cgtGwXphRJZ/shB5izQfCGev2QdZA9uu07KOaHfaii37vX6nu1Wk2AoujsW2tPp+X7i3EH0y7TZA
a/GQq+BSVs0zEeadIS4y0wPoX1DPIlJTIriPa8cvypAfWh3Bbi+9N0VEB1nXTXPrqlHV4rLuwTCD
EXXI5Krb1ieMTNxpom6XpIoZ34KmmguSZAIRg6EhjU0jcSDj6mfRhtIspL7TyW6H2CN5Fv6agOpL
2yRscOg8VW8RcjsNCNwhfESI534tu3lM9ZRF9JypJcoK9ZPb+CYNC13Q+SsTs2v3EHd6SXGQrFti
MHPiq1JJWg+0/0VrS5iM65tBw/sSuIja6aNQc2LUaJjBxE0tBeIMHfn+yQgBbbARvdyQOuqjiE93
9r1m1nLzGiiYA0wjZzJig+DDRidswdVn9pH2gRNIQUF7cice3kDb2cJL3/FN4GzvxOtGCmsrb8af
mYaCp2Rg6g7cEji89c+DBipOsl0oUVieXEgediveMkO7PVsvTJJkbDe12mhwsXucSJpu3h+7MIu1
5uvV3vYbA43BvhSS8um4qcDWB59PwSPemfztVGBjpnQ/44PIaxAh7xAEXSlw/RY/pMO9+/EQou+2
QuZFOtJIlYnRIWC8MvblU6AoAPwWXHfnrn5EuDbXuwR2h0J0Ni8lWeT1RoBih7TjgiHvwC8Q1DHv
n3rSFmijrvFP1jVoOcYMLMNSPZkQfGcQxcWw9nQBofm9F1a54snbvGftJZrk/0ppyA9No0jC1XWp
wrClYgD+eCvNifYOB5/d7Jetv85mssVfaQvypjj6l3VFJ4mO1XrX4m5F2o/xc9Yjm0MQavjQnM4b
q0xx+d1yXME1xtqt23iA/i8dK3Cu9jo8zG5C63ITWTYCzppUiOhwCFr2+dZIYzSayV1lH6npZ5BU
oC0qLn0WkhlqidKDEbMAliQFH1Cqf3yYOGoTz8OjMM9AW1hVpaaDoI2cdsRTipq1fTeWvwWYzeL9
Ju0GC74Z0mrtoLQYFfw0FiFS3mTlj1XkzG7ywBUezukCo8iKGHGZvJX1bc2NVgI2jZXNZGV7A8p4
wX4DFaMg3WZ48xLlkXqVupOiBohIe0ADgK/JdIECpFkjkJvp6H/Z7HuO/vdF/ceLd0boDM2QVSY0
XTvi2s527QXm7hGa8akrhKoJgv4UqCzCsIrI/B+LoBeiQP20k2JcTDBKhCcU+IOPYJZ4DI7As+Ed
rJk5uHPMEjAhWghv7VFsw+TkbY1M4rDR/piFz/foUAMF2udlS1Nx8y/qhIpxbHo3mXZVgU3Sch/+
bmus13PeuLT0BAYcfuf2JZyLqsRw/so+a8CPRzBlTfran+eq8hAp1iLmJKSvvTDg+RFcFH3ySg3t
fMATGPcBxlelpsbJWx6PYoIobCklhpuJxYC2rUWWqXZXIK3FoanFpWQX3xq598HlqNmhKuae4Xsu
qtetmlmlRCKvajjD9jqSuuSijE50udhtpQ301aKey97RN/KMoGYUJDHmnvsZDeh8Fzg5/+VWSint
MtJP4u/HAkAJ6v6s4g4gXmlopIvPYF8jr9/Cvz3mP8zLgyySXCJ14FV1WJaIbC2kc3xi09ozaQwX
0rwc+QMbL/1dm5p60ylVZKEQm75JLSr+xrmev23N/PP5oDEGYl97nonfd1S3A6r3PiNp66Dybg+K
oxGvCylSIK2Ox5RfCsxIOfdThAvr8C/7gBXYDkhwUfYHnEHwqmtgGwD2qOtd5N5qqai9DJmjSQa3
DJmnKKJ8htT8PQE+g7XxKuX1mGL26+RKqxZaAFGjvbouUCyHaWpUriloOLCmJNbYiSZqEd/5YQGE
z/MX1lDbzC52d68iGlQVlrydmMDNJmrwxLwmPpUwvkOUQn5LcUlRbwDFzGrhQhwWzXrg9yOtzupe
gKgwN46vxHSElyYoXDTecS0MOoC4bi/K+U7ivqSbHPtoJ5AN5GhLHdNkgK5y7wkKiwQ8UZY6SGpq
jtXTiUTiZNCdSdhh0r4sMIr4OSyayisRlMPau/Y6DPA2lCPJvrisQRd9op+nZuwEwIcjcmyhSg9I
W03qTk38j3H2fxpnduS/TKY1A1YBU/fKh86Ynj7L4iXFw3zzJNKV8iuiB8b317FMJ2HVDUmf3jz0
qpvgifXuhFVRNc8Y3lHDAqw0b4Pk0HzVt2t3PdGhGtA5ZCEiOMUVcHEVF5tCOM0ZO0prwpLVsKe3
WnkRlnpNdqvDOQCDrVqln3SKpGVdN1d+g8wXVOn6Hf95FUJelf60zzjrhGJjbgVjzMRUd3Yxh95c
+N85A0PA1VoT+JxeDIVTCTUXbWAxRQSCOaLUk5Hqfs6Ss3K+CSs5QBh76984La7nPLgcPufOymC1
0mCmxFWUBOnh5xR5UfmIUSeljG4UINGSRSOQ11HSX5g7akGQ1Jz7yU8Z0fpwfq3vYK3TKGw1i2+A
kVdahmzN+HYMsrBpG5kvEPxSinchHnDOAmVzRxMn1SQPTp9qWD8v29NW90x34wEZNaNCJ/Pfa++j
h4UzN2IbxG2u197wp/ktBuvnt9P4WSzc4Qe9BwxpW42kWZxo+JqF2AlnGAomOAEHpWiqlWwTqAEg
Fijkduj1mtk1X000AA2bxQcI2EnLpZ9DfMG8MK2Lcf45qDqK8b82BE4xL5jCeRUlEeG7wvKQfP+j
NNRYDXmq+AUtA+974DbxhY6hyl3SJDsJsI0RKOsJDVIoPv2p8DHeu2oPrTmRb/UlZaaZNeOly3A+
YrRLNFpuGLFO0/flbpSs4+y9WZBiCSLi1AhLXjmwt5NNRzKhDCEYB0sZ8PHnLww6d9PKwG4KEVuU
iwp7mr9zjpkZ2BFUYhzZNKuWFRCWegzxBLIOs4SIoLRD8HATTelzp/ZFV5Rv6qnh5LjMwE1uWNEC
VL6qBr9RdsMwaR2tUjFW+sf3vvAotsahUXG4cDleVqsN3ZhcwLNH5CjJpOpFP5ogB9RS/Un8rxfA
UkpWF0r2c9atOpKerdPP0kTlN8IqGspV/LQYVL1JlJaHR/gB3xiwmg4tyyyfROL1VACZ3ZV43M6L
DYWiTCOJpig7SbuRni3vYXLNTWKEQWClnagjZm1Jwy9Xc7SUxC9zy9COFDbctVhBzcGNPbOIsunt
bZhdbeEkkETuL7xdQ2RaB8c5mH3nKaYx7JbCOYIijQZHzq5PHVcq8xFgMawYSXjdPvvdVTozzKl0
nRz87b6miMIuS7xZDVXpmFFVAng5JcqGeteJcKp26Z0M3ZrFUDmt/VLf8D3+2J1JQ2IpCk6E+Ryh
lIwniqTYfCXxrqy0MgaovcxjBkweAwTBUViqgmmYtn+NLNcdWIF4zAfVOk+3omFX255dwk1l3/9R
bFQlswCYMV8PvcmE6XaTVLDeFr3xRi5KdE/juP9odTMAxbEP8hiw8CB0anOL7euNeO/lBr9j8dkD
m6jVaaFq5e2hh+AtT16hQJriMqnLAqnBeowKmGmcXn/Z/sKgVd0+tTp9A2epeSsJZ5VvzBoIi2GA
4ZZ2qpbS5U/3UFwwfVT9/6L96W5yEuxOI2yXlcHMkozt2K9B59/k1qaYQCtr5WFYNFiOcJFXJNm8
RCq4WoZsemS52FL5vynXv/xI4fAZwdq5c9GuHlKBzHPPnyd1d02/j1+xUN4pO8r0DdjxeXjdCwZ7
ZVXB9y80rcoXxd2a1zzJW2H0nnflLuMmfBUzMASGSzjYfzQJmU7tsCjv4EMB2oOiSZRr9W6IKLe9
G1/BnYuaYrAYtc422uEN17O9caq12cJQiKx9P0cLvB2sPfnET0jwwMQ0z0b8nqIPnd56qQKaaTdO
WmPGbVwGGZccnHv7vs9rJh/S9bgu5B1XZZ/zxhcrebtz61IkUy5Db8VBnpWr8dGNCWy09MyPVLw0
qfBse2F9Fs4dNcJ1FjynYN9y5u05MATsUOxjng60eXAvoJYevM8xzmFfdxFLIvKryxC3p5v7OsLZ
JxTKn2icA8ygUrZ7TEjiVY8jVlvtDSI6ug2Ix+/bd+UyBZFlR7KrhzxFmQzK376tgqgChxWXt5d4
Ci3NOORYrNPmpKBtD811BNofy0jUs5x5EqhzKQCExedCg6WWAkivO5z4riV3IO46tTWtBwFjGN6K
5B+4i/8vhjPqtD3hxk1mRUFPhOmylUwI7HFJ/4f//IcvKmERfb4DQkqiAem5qolG5QgqxAc6jGVz
wlniL4He+TDzuCT3Dx5ofojavck6gmxLnyIsZY4OOJfCj/yY9/dwKE+NyaUnFAAWdPjHG4+1Ub1G
279DAlVgsAGjpn0eAmMCleh0EjV28S6TO9z6+HOQdPyguJ08squKHsMToKO+ZdjfV2DJpQrENuQl
Yy/jNSGit1x2wkKxDVCqiMElqsqfDEBu9ESRLgM3geF8DyHyJ+EoJPmDUDANh1xUGUfAu4Xp9AEW
4Xv6cHI46/XdS2f8hG8pIi0SNGzArn/aBYdbwkI10kmpBpOcxsbBerERX18ZqSOeuWsD6540aHul
6jTEi13ybxZuVfAqIT5q1DEWfGf01Ing79WE4FR8P69Ex4wd2ZrQTFBFD2qmKAMLeusWdzZEt5b0
Cecgqxnr7jO+gHRJgHCK2CX3cdzI/FgWqQYdEe/zgu5qhVs36WTnUCImCdDFHDvtOUUJQOUmW0xx
zHykfqX6Ns2tRFV+UJEQeTIb7xwg425xgFR0+3auiiTcxRwW8kUkuw0q44jJ0BShpW/K+MPScH9c
SC33/i3J/2OcQt8kMQMQFCJ6vvk+aR066ZK+PbYBtckQSMeLamMpyoskA/r3QUCjYUc2NHdryd2j
Z2CCBCvkgUNpl4nFtK/3K0g1KTeOc3XNbDfaCn6RsL5pkL7vGRV9PLAvXGLvFEqIiw0YJ36ScJhK
QgRra7dYTlQ0dw1GtY+VkaDqATCWZMS9herTGPQgWetZm4Ky42hfJzzE63kLXxe4U26xlBtefsda
Hm11DSpLCiUPINAuxx0YXpDBAfFvLG5ZGxHKzWMlRtSNvaetnK/pC95X4prtAbtQMW2vQqgcliLH
jdG/TX5SHGguOdjW1evREc5m6vIvZ5mzX2paRQSRQzhxFeB14jwDQtJ8rnx4AgRNsmv6CpuwTqtp
n86zxd5C8E07tJ9AXVtn1Vu+Zc3IaHu1xsSLXvslkv1ZASZGH1TwF5oHG9MdsF5cFpVdwDOW0tHv
79yuaU4ewX+QUfJqTqdFy2XaMNAI6z4U1wBohUaASEHE5lT78O7NA0FqjRQIKkKK3kxsv/4gd7si
ss9fcuz2OWk4Kf0YQjrh1q8RJnp5WhmCFF+/fT4xs0BKXsM49cjKD6Sq0IHY1mlLKy+SDjKEnkbU
etB0xB/LfrxPohJvHoy1F3EDSVrHuUbf1s69IbiqdqcdtgMrKrACDyeVXvanjsCggURAjkwOmUTJ
Hmd4BoNK+QfcVAUAW89nL32d4jo6quZlcyYkZ3aV5LP/Fs99otztROv3spQtqS2XpOMVmbRHeR/H
ZNSoEvOLx+Yu8tmjrfWOF4ywLtDQ3teI3tFXQULVOLmU1fXxypqs2HyXN8dcfBeUNVZsTRrxqlHL
fLVUXGh6krmPaZtfSs80vCEmCB98iMIy10VtzMWu9lrTK1IgmHQbhC2cW/g+K5y1O717Bxv4n8V5
bdLx4ffZQuX1yKq6D09ykOCOQAwzEeKTcvHp0fQEn4FRJwSWIptMh1rxj8OZK3C9NRCl3s1CulCo
Fd6U7xTVnDxkiCQUiDvjWZeImA8qvO6G09aD5BDmEtmRfS+6c6GcoCZX7yV7VlnlF41oY6T/z9kH
J4GqoYAcnq3Xo90K/Spvyq3uLaVUsyexcPLOV2FCEOGIWN9zPI2qaC7ipOaG2E8DRuz4976KIB13
sHvJohpvrd8RDjvwpdUOcl/bBbgP/5ROegoxGze9rLUFBUzFbxUF04IgH4AYZwjWaRYUps1fv7t7
IcLZMYo80nZmA3YQHzAQszky68DCRCA36CjyEg23fe12vQPQ18NCNB/VNxWtIz+duNgS7HObmKEv
3jk+7S3Dvt/QbieX27vHjRPhpDgMRy7Odyd7NzEDBrXdRzwHFo/ylKCcVSEjSwG9h8oWG/ye8Hw6
XFX2MRk7EgyzWhFmUakZ5XYI+QtSkFSkBZtI4p6qfxKp25PLmufILqrZBK1elFlKlXkcob3hCFNd
hEQNQYBur1+8Viu4jd3iac6d1tM4WBGP9lTMjGmaVH7CffxoDcD8qJ7ohmHm52IxkT9dTuiONdHz
4QjnI5jg+DyXoj9nQvOWsC+LAt/4fb/B3uOp3huNWe5ZSYmV86PkYjwKFeE67wUzjUew/z67X9oO
Xv2OxICShUfhLHJo5/Zbcu94uSAw6F5KnCpTQmnwIW4w9F56HdCCuZ4k1IB6Cg6rrGXCuNzdl8HE
CaGBgQJrRbQLtGost+c5vNlm8/P8sxZs+Nv80ISVD+cPbB9Y51cIqq4sc879i5VDK21vYU1QM/Sv
oSx1VLKhhFPyvDWJwmu4n74tCOSnIOOZO1qVhOcwxzqUWrhh/AbmOJ36Vz9AAAkQOUt4TPJ2TtRD
BZyS27RMlxPd82Ds97FEnmLpM4MLHQOgCPiaYvw+K0gPQVOrgNStTEKWqmq2yuc3vttyDNRuZFTh
PdBdUlcPXTbSu3s4mhhHuooYRQospHgLAyInLWrBv7VFa8B3+ItGF5zdTzBLyZ08wBMaWZvnvyq2
N68GZD32OvrIbXgJlKqNyNw2xN9WoAelWzrotSa/XetlXNrGppe3TgieRQVo35aWR12D2Mk35TS7
MQ84EXfqkXuwX5bWHuYq4KHd70mw/AVit6DgTa8ifaW+s5PleMhZ/89yC4EwGEaZ431BNVUpqzsw
79hWAabdDf/BdmglWLmNYI588Y85OBJHeDGuYT6YjVauVgQ79qDZUwGhtBX0KchPJyXHkEjEnkQv
Kj3y56K1ORYbS3fbmI5pLwqzG5YhxnwQGOGJdXXWfHM8Fjpc4nAV0Tpn352hW3THRH9B6Sr2h2ze
lmCRnYsYaX0mEteMg15k7FvRRJEhdkS9iV6oQSoS/NPrN0p7CncKhY3wu9dIx3wrrOQOcW0mfVeI
lrHESt8H64kZveSJfmM/ELrMVG379V2tSmtSpfVRmPzkahlhekWM2gk7k2rXIQsBV5pdFArPJdSV
l5GPm9hH7LTxxLvkUYKdMUV5nouc3JUyzw7dNdE5m438t/RzDGnerePElG895m3dXFx4Ny+IrbyF
ktkhQv9uhHUQd9bobKmQxUp0gQDO88BNAFPXVpvgS+efLVpEsGpJgt7gcaert6gi9JI+nLFgawbq
Hk2TJuVgFAEodtCtyH0garcw8/re7hJs0RlyjnMrCDbnKo7TdkCo70zH0Bq9fElk0TIpLYjglN0E
wg0mxxmAdZ/RZfTMjUXSzg1zs5YNQucqi8Biv+zn4k/uliEnpLF5JCXJfPjM48u8UktsPn0o3hHv
Ht57vVHn4WAwoRrAohyMKX/kVJQIV95kRtHPGEf8ZrsWV43QnKhidyDG/fJxUwgsRcHQNSxZ81Lc
4qwd0Zal2Ysbn03WvMN1+on5QEB52tlEm2hgKlQkCRYONhdyCP1VsTfJacBYp1NJv3t9hTWb4iNn
zSXAoAxY/kNdor/PqlocNKyRGEHVcfjVeMVbxvSE0DOsZ5UPq2biFnWS4oTjaZIUGI1KgS+/4nF3
cXCd5lxwKQ8d9m8Lx5wBj+r93weOtnuBRYJCA4+zO0Tb0Hpm7gC0jTNQb9a3R44CPzTGU4+XhJbz
iQrM3wODM7IWCmpwYfgzJ3NqCi6RXZUbeb3pmjVOQB6J1qEH5DEItmhFXb+uyDN01XVSqa4S98CW
eH28eF6g0S1i4a6suOwQNGmqYznm/1l5c8olBICjEIkks6QOca7Gf0Qz0h4fh4sWoW0td9goBxf5
SyNOEaeMgYgjR7zG6y43QiLBsF5FTaFaNi6uGgFvOVFeWutbPtAWTnbcIJCAOLgiOUobFv/ntASR
cCYqEsdXb/8MsvFsxwM7/jnr+a6TmRJFJka8Cfm4E1yCyva5JFAOZD7HOvZP6L7X06f9f5+FwpcU
7283gsDjqmDGZPwHoA0bzqvGw4Zk89zX3DB5phb3Ye53D6SPhvxns5BfdRLmXo0nzNechh1j5ZdO
GryeMsFNyxGY+DVhwEYl81DjM7EMPrgkAxPyzOGdqgtC5Ktl0nr0eNd/l8SDSiHjt4syquvhrwN6
hhfOWXDYLUjViY2lLVRTeIOF40ODCgoddFTL216p4zNIGVft74Fj0boqMDbPegt5axnMYFCJLTRy
0JSeU3Y1GVl40IWWXnTLPd8R2SqViTdDFvpdVoNo7KZTSnc/GQNsBVwbwEoCNIrJI55jenZt7uvH
acHKi8TVxzaqPjQ0fVv5E+fBhhLFApwNh2CYAzyvZtlNEL4cyBdS7dmZ6ekfGcxa3bOksck0lJzG
CgI9svvjuniTAUSNkvs/WF90XuEJJrjvs9pEZjPpum4Ov3SoUmPrUP5SKvmo0e4sRcHhFjSzDyl3
tnpR25Xcy/JEuxgCKng9wzPTrc0EcQoL0h+EbUhw7Xq9z2DqrvwfqlLPFPYYGDZXmCtBrDTJ+Y0k
2jBR1j8BxMw4NsHizIsE0KkrvRb2MPF/mQ44fMePKt7n4YU+Pjx4HdrZALebW5hIbCCUnVeAN3YQ
wSm9hbbjEiyCpys1PFdPkddjcBG7zldxeyEbgH5r3zN0y+mfIv+fIfVQUuUSqsoLL6y4EIm6i1ok
S6TztLWFFaej429EPBnmqO7oYg1cCpaan8FkORro69GMxultST0anSh/gWvP1dRrio4OiWn1M8Ep
Go+0xMevI8T72NH6IyscTMDwFGjzaCPbP62wJi3FuXtsBv4BeTwMcIaAM91VTqo3sa6A3nTaptOj
XrzQcK99QZeWZyywTVMcvAKIpEU9+XleH3K3wfxsr63GOIFLq8Ud8lFDRNQRNH3aJiohivU9yiqR
7m7YB0ZL0iNOJhZKN/iXYJI8bQnyO5cmWctXMeTXcxJWX7nde8ULO8FQjTgkMwAZ2/bkynQKUsDi
OnwiOnjUzH4cbrFGdat6fXFjRb1b2N4xO7Xo4hih587v30hC0AVSIhJ5fiPi5VdvGiVPDhXoVu3m
TTxRiyaqn5J0bO/Dim11WWszeEC6WQOfLY8GOO3O1yEdtR4sViUvqqrgy4OLj54dcRcZ51s3ZFRS
jrrDtZXJAKcWH0mg9HxEZcbHhvRbf4Ck23DM3zRHAiYI0w60FFSzdUAghVK8LU3NAEaaVHNW8qmX
vT5okPptUlO9jRZN94ZJ9Yd+P24mBqy2cZtP3yGGHdfKWEwZTzGASRFzpRw8PkZmrB8EzezR2jW0
BiP/bKluknkYVbTib9mH9YInM9qnwTRqquq73hm4Dp6Oe8JyL7VGJHY2YSz0xmUM1sdoQaNcV/2d
Dmqa7/A3WEl73q/6J4DjZ5TE5LgewCOSyQ4OjuRa2dkc0GlRJiVSAQeH+xZKcK9D/X4e70/rDCrc
aJbhXb5Rjtjytehy5lMv5ySLvVil9KlBd47QGzOWXo9wdmRshc6ER+Agh0HctRjHza0i4458JpBL
LpJu+U1hbBqV8A+AQDhaGNQnV2KqFLNp/lmmr6y3awRt1IvkZBymfgHQbw807sSQaxGyz6CaCZqz
9LdqUUIt1K5KmpoCPs+IZOY93j2OHCLfwN5ZC6r+xdHhPpBGnqU0Soe6VShDpTi9clTL12VQ/aUK
2abyab7lRaVIeEsfhJSzWXYaMrwLpBkyKoiEu7q7rnjOLyVQkryDDMmI2S5gzJjZb0647qnatTN8
Y6MMMzrpxPw7fU4pkTZhMFOU1B15d8vnmLGZo0/AjrpIfrYpDwkHbEGAd/xf3pzQdHE0gjAVFRYh
nhiauM/LCCuqFGUNpbTNfPQxa3JHrOHeC5WjON00kRAzYVyAwYVtd8sm2eMMjkFMRdWpl3D7oRLl
jOGpq1TUTccriGOIFDjHqWAeQkOGReO1t4UhzAIzQbyIeQ5t1xEnP1ZAFooJyw/BgUB+E9CCdpoD
L6eJtEag1p/B6QTDAKa5Rs5RpwFSv0pxXp/Ue9QVoBLKYuDeUPzR5VfgTzvptdlieChfEdaK15VB
vkry8m5+FDNJruePrNCTonJCDcwV9Csq4HJkqqedwoYaW/EuU4roBCGFmFyJkoqUseljJGqW7SyE
d3hlPYEDJ8SQ0zMAednZu/ZiK66CMXYiqQCEtpL7Nfv1R61Y2ZinL+cagzI+ib38IbHKt56ODRB+
u66O4ljHS/eI6S9UFjloEVepgz/LOOnIlADyl/II+F5R/nEOcmB+dp33ZLW5NXySSuUADjmQFyFa
XVOQPdJbyH1hW/KKpfk8XXstf2m57RhemfFNs2JNi72sRh+fBMvBK526wpznD8OvgcuQDnjBafLx
1BMaVLbrNP2VmAPOs01VrhjY0rneAuAZjNgEuKghnBriNbxc3cNtjelfAaFeWE5cnCcQRneu35tR
6pJUeNTaizElfrKpksHZ6G5w89vZfR3fwkZZj7nf/UAzoBh+h/gFSsPj+GFM50qJDd0F2Od3uxnf
r9dB+XYWxsfaainSN52l8ZcDt6wZ4p/Z1ctjGxKq6XYLXttrmw99L561acr6+JAKMbdTtHAdf9NG
bWR4yscOrPOsCp5W6E74F2lACNP02q9nGlgD+asxNNj4QH57CCQpHCE9mX/qQaA4nS9KLHMpoF3+
zY8rUOPV0/yvbzqe/A9hm6rd5G9qCUBb4nWvsp40gBUqIbsoGV3Br/zSvPsX+BpVND/ElvBlYWJE
aom/KrfQfMkf3yqkJZI487rpsQ0Jku7I7MyYHBm0pEvU/+NXsuvlNOaIRWFanddb3FtV0umrxNr4
h9JDJypMp8lHHOgPXLfPyy8CzLroo3CqKFrqyFokZzfdRKkoqama0vGB9P6qKR3LVwjBABUPrZpc
I9dboMAs6L5wdRnh+6U0qoLiEeTi20eipceHvVR0/TpiU9p4bZWu8h7Yp0h53TKKgHP0KEBhQhX/
0DkMTbN+SRlN3QKI7XOKBp8HleIPFy/TblhWO1qGSU6/7MWJxkVz/vTRImX1WQcaNCRLvpATMUEp
WfQeY4TqpwhksBVurgjx/d04haSDlwpw2HBCKAxjvn2Q+WHJ2ohUsBDbMoQTpW8dNpwx7AdlMdiy
9rHYEl9GEBDXUYr+CdcgQqw0NM9DX3jeXzNqa9oDV6BBG7LowMuAlSojRmqq+yYEHp1eXmHKoQR/
2uDft3Ze5rCq07CwgyC8ZXPI50w9cbZ/RKOvmHkj5O90qBIHvLwXAorSnb3HfcVvAOGLi6mNfu6N
cfiT3VTBqjOdAmIPVVR4d9RVouNo6+vv6qd7wSZJavOT4uU5eUnlRZlqlElHdzVr/frWRYptarcw
K6YVDQEfJrcJFWBRZ+Nq3hCqzzREhrALd5dYlMColy0/QfHKx9wG6A+usXGx+YUwzAaEuS0wCHkA
NMf1TLNIikeURaruH8w5mvDz8tPbLwbsCiooUge/W+VTVZ+gmPV/yD1sn0+wj5pGZovzIzKVM8Od
AAwtDnS9unw4vqMKlUB27wTxon1VKuWohmmDSWdXuJxRXaQmiKstyZPXMF4fqN468kred65ZVjGV
kJxB3Ihok5blGPrrhMFI2qxcZTQfk+6GpzGdVD2mHEGxryAbWVeosjfj78XqGWeCi68UVU++HvCg
zHxz62IxkvTNY/DIchEXcccV49QpTqSHaMuTcPiqMwrWzOLvZHby7aQl6BoB/dZgj8dAwsRRDG5n
HOPM2ffcKBZ/xCuUBT0eC4pCyh+oxL/y4C8Bq6JxePNsI9RQgHMXXkbm6060DMymH0XEqcaVoRl8
DWH2GsMO/5t+a2xeQ5H3vuepB88MUzby8dPsI1k2mCPky0/0lZOTBc4Zf7TqCsVj8LzMPQaLSuiS
L6qqSKx9rfxaxoHSSXlYvS++/4ozoQaF66ZtFMcB+8cGR+Td6zG0vwqThuf0jIBBjssoIV3SMHSi
fckwaURcp5YpjjvgHEWRwKb0xSN86JakSXkE2ABs8kAxf1WVbUz47SuIU3xK8yDpT5AMY+7mg/1J
EKSmKpjhYkIUgCoXQkGuptKSwZVFVI1q5vd4Sc/sHql3PpCeAu8YIdbnLlLiwdS+MgWoorK6/GnA
aXFCGw++A+SGDDmwAsjyqPvsIKqVkwqUhlF/fR0DJxUzm/ZZUjpVNxkJlTLhhUZmc/BdpPpYzUHz
n55ANBJth3r7ha/WybsuWpoDuWcZJm+2ixOl+wmhxI5N4M9G1dD3mAWDhW4WA8+SGAx2Ief/9rir
fZfTLRAM4Nc0e+I8SQUMB0Be+7CyW7FqbWmWYvYuZXlNRm1oRbQzlurvHXSkoNAR2KLuf6zCU79e
RSS/BMXN+n2OjUKxDhhFf2Y7Ws0+ZWYyY5usy2j2jtFdiukRxX8EC++Anns6lI4nCrURnnW7VTte
6iXE1qOKurn905ikPP13iExPttyYs+/b5ZjURDF0BTwzoZR/t0t9kxxifPAVAyQs/ndxU+KwVzGb
hZKC0sSE9Rlo4UMG10mXJpJesc0GcLdt8wl18J/3Zx3PCBOSOQkaX4C/cmwaUxG++hGjaMCl7ZLd
W8oWqM9Uq1Ssf5TOSqMU0rtf+TuTbFa4KA0qrvSucP0vpxgPMQ7RL+vXFqsTdrAUgW5iv8Z5+YRU
hWsnh8zo1G0Zf1y1r1l7wwokQMEaNY3za9pVKmSyD4ywa+fFeQAS0H5R7O436C/YwD/lf/yWbNWZ
UA+SpXs8cAhD0pxrH3qqhGQ6sLfH5uLMswk02DAKdfGiZpEYIy3D5Wg/F3s+G4NCo3c5KHmXzhda
hv7nM1MkBV8bDLhMjvI6TFmV/pAbwbp7krEubiyxoRD7Je/g2AJ59kwDOKB2FYGsMjeCfhCY+t0G
cI48TyQDGF2ag0GTTQhrlgylBcnEKTKq8mc5KcEHEteIuezE9hbUkGfFJ5i31zbjAyxrT9vttBjI
pOMHpDhA99yt9zGAaM/TMh0MZFawhckoCMUnliXpj+tyybMzCIpRb44JpNl+d9EL27RWqdNdIVFP
O3uHUAmVpgzZSKugr6gDzyRmPIGhEYPeIBY3BosN/kHjJB1I+xnn5JZOp6+1BwMKA5hJaR7QAryo
8GiGB7fMkLN3G1tHJr3KhFQ2++YLopyR/PnDbgW/Whklp31+AdvSysl882Ll92pXx35GCWjKSymT
639erMdbfUzjIjgq6mr57zK2Zca+flLlO2mt4CsI//woGHUeLRr/ENsloXj8cZ/U8oHKomIL2Lhb
NL3S2KUkq+2X/HDPid+kQ3TGm57JrHr5OYfCg0S5I/9SH563nBbHOnlXRmI8xg2WAg3Bh7KCMwoJ
9Om1zm/HFPeXjahCmrUhCaMdQVKMQE9rusOKNt2sPTHRMek21cgT3FZhobcUBuM48jrXletc+7L9
cnb5N3BFpD+sEbbsbRH2zPHhamXvMkuPlJnqf788shyeW32eqmQ9DgzGRDu/0YMS+lJzgb3HkPej
ptJAK85lOdPA3FfvSvuZDDGcbBtXVIg2yk2MAGtU7zms2lnADbHVmXPycv41xbzZgpCAHp4CiWb5
i/777mB02scsxGn+aZb8XUqS1MBZ37nO9qejlYuNWlk4ii+tcX11iZFi90LgjdKyxlEh+Gm5O4BT
98Mv05uLnxLlEqn+9FrsflXwJwm7JnrolVjv+P4AW8HVhBK9LHx51iROC9ed8Yzmy73AT2k/c03Q
ygb6dwgTxJOtpxESuweGOjov+zidsRSQtwr4R7Gw+wN6enywZE/aw0nWSqt4em55g32oxgng6JX0
g+bLeQGl5qukf0TVdJ4IwSn4RXOpOj7TGfAORMJ2tKKAgA796hdY0J45sRPxpqep2Mp5dxdhsmtx
bhniSKT3MLacl3ua+c/dGQWCubFUS4jtG53Lxpr81x8aC2p/7C1ac/n801weJS8VhTx88yesDgmd
Oh4rtfHB+MX+rM4xTEv4zFKIwzPcG6cUFVidh6m8aFxIl147n/SCKZCce7yZ1hQKWVJ3dIdkjlYX
8FjUpgwz8oKKHKBFDK8BvN393ii/el0i/4GC2jkI0zQ4j9s0HYM97TMonbzu3xqEFussXkZXRKU4
kTtsUUJn0EVm58tJ+z04pVpA02ZiSjOZdI98dNTn2S4MJ4M7kj0I5F+KjvXSjpFXUTY81FN6luw9
NV4mlibXPoB/TnXv9hVpH1TWOzTUi0yghv/EjWiupmzBTqwHMb9BiswjtHqajuogZw+qieU8jGkz
8xkS2vOlyHr2IqwxQFq29pF5IniJ6xZ9dvfwso929MB/UXBnR+GIGLWB6DFN5OopQ7wa7QMSJqGa
s3C/LiHX263E1Nw6ey/Ee+NF2V+7RBQ/SfkV4L60r5UfVXiSlipEDopVTNRN7RNJvGwiZs0ExmfO
5EbxUwXJkgReJWW0fgMqTRXS/BiH1MeAltPQluiAB4yhiw/f96R26iycfJW2ifmHsLwfIerBOOdQ
gKr1PQKGrQOIWeq5i49YfIpWmnWSlvDbFhwjamjcSNPo+ooe8cu9Et9k+8v8zZRhWyIwRBkAz4Z5
i4N1+HtiJ6u6GYmNdMR38iPfqpVAFbDTMALCLf1nAdP88WDrqW/qYbi33NNkBN+kbF/r58tSMFIA
X7bwqV1FPgCvwywSD197sY1GRxUbHbJb8jMGAUfRdL/sOvDusZuCUYvdN7a8ZvV9Gnys0OqeMK/2
7cN+N6HP+4v1euidzmMr/pddtVph9bxNZnU2z4iGCC7YirEZdlfXbSwCblWtSumYvpQDFgtUYl5n
bGtD/41ZzvhMlIGK+8jXtyGYOtdSVp9xjGXjEex+0CumAJr9c4SNHJPSprfoCfW+eiWhTRPmXBkR
Qn1hQT+TmW6rcXLhqbQ69s4v6v0zpiXWZlGdZ1KMzg1brJqUSfb/waoXQM4XGEcEygXBgqeSDzXM
4xnCKhCx5/q9bgQrqEEDJKLWdm4yEeQbghL72q7XZEDTQCBipZ9d2eVLAa7111VnZzd0DSgih+Ft
onCRA4B6DoIa6sfs7k3MaCSLyQPYtZy6ggD8WU3BnCIPIPLB25c9mPxogUv30M23OWYOnl8d9cuk
S6+Uh5RDV2mdLfG22CfswvuPytZtjvBYxvVDEWdKTEYJiYTzZ6sRzBIETYJZRBFyapeC6OPsDZIx
kQYdpWfLnilRUK2HOLc5NU9zxn9QA6xy0pCZL3IGaqSuw4Q2glMFBJNIidj+mIUf9dTedIPldMfF
5IN+5OPASm/AJTtcwK2S6RaVWYDgn9WxhYjxA/xBJ7v6XeBI/JHUyVmb/xRt/mCOP2alu9ic82fo
QqF5pIyud7yQUUBftULPsDYbr+Y8m3ejpagReyqE53ZIBkTy2PAPFV9mLsYuIvt3c2zI+JjSjAWj
HnEkQbeoURntIwDWMqUmXqYyLbHAikCYjUNt9wQW/jwUyBhR39z68n7FYyHxy0TtoMu1NbpKoDo2
CWlefXIqXCn9i9AtXQ5q1aFw5yc4URy5Fox74rwHLdVfPl1deoJO6MaGXTbrcIZK4tBY3lhUuAUo
2cSa7cim96p3PDOMJvV/rd+pwEKE+ywtzx9yuiF6gy2O8OKw/d7pjRnGLgPTe5jwTZYwJxsdx0rn
5WVgbSpbX7rrYdh5yCH07gOmRROEc3UE7VyCvrTQSk0VEcDIMW3/J5FJylakH9iAsCeoAwC/ocGD
hMZq5Hm9zNvwWUYWvZYDPpK7+mDn9T8fwezpa04BHlADNS1X+YovsEkqWgkJfHMWKAorQD4+EDgy
gKm8kf/ZW6lqensUUPzLtGdi3yUikpFUDYpRp5rEQBNe7UjngHR9rUSVlGidcMukw78VNdWYkpLe
XrFRhpFStOKHAS91CKUKp0L3rRit8+humDNULb4cb5qx7fjBdve5iFQYWEuhGgOv6aVz+uib/zcj
5tppKxeL2s89tpYVsJaGBRDyFTsoPWKbLZh3WA/CDUmGl7jl7mwG76P/lN/7uZrV97YRHrIE+vMg
qBHx0zi7yqiBvUaInQc2peVUHkFfikLdR/nW79pFzssCj9YEydvHm+zK1XRScJKu/UTqxkWATjrK
flxNx2DKfKr6ac4PB7i4zdrze9mFlYdAnizqpGScOYWG+e6udZUZrNxQW0cEQZSqhmXnCt25Rk3F
UQJ70Dlj4XqA/B0F3MU8W/SOIsQ4jl/iNxiVuUpjV5UqqEGwsbWiK1Mlh3BnDwW0FSIV8ihtJ2/J
Vbdj5Xxt9CpePhapKjyaqwC+WYgU07x72fh7O5FmaNT7Xb/FM6bK2LRIF6B/rzBEz0iRRAourRgI
SVJjNDOhcjUcexawMuktD4K3xz944qiubR71uW0MGsX5yyB3iPxI54ASE0jNB+Z+6IWSlt2r0IZI
oiqGnVoA9B8YYViGDsFuMs+84WNS+ccVZjpnwadUKCQ8nWEIDsS2N+/nNO8IaKbA+7FWnzyvUEqB
zM8SioJftWZocgcsdYopqczovm0EmOV1FjflXJzFAtVWKwUwiemv/XUbFCXqmFJNwxO9zIcIv1hQ
JR8SFfdWEV3IVAGw+KsDFX4JsXTayUxHJ8SkBW51kCrERSe+JaqhT1bU7MbdBDCs2rKekV+lPfFD
O4evVsFs89iv0N3+nBh3a9l3uNDOewqkGNmlnYwkdANsIR4t9RfPI4rrOPCmDWCkcNXaFcPF29EQ
Uc8ao0jil0OVpeV0czNvg79vY4Who9++0q517MqqYQQYxeq4/WMNtMvlhZKatJxLgPXgX/dOki4F
URozQn9Z/t1DeZrJghJ7ExLg9Xvr5l6pJEoW34RN6AxaINrLBLVYI6BGBjTOG23ohf1OtVkSqkWu
oJbS9UcDGjJ6TXLpXBVsC2jwOX9UilZWwpnNLyaZHXso4LLVNJZKXhG8gLPxxnjO+LQQB2awaCW9
i9OE5P01uDcp7aqYhuFFBfZ/8Wmh71bFzMbVg2eG5B33p1gyXMl1rYzC5uIJjhQJdsmOkgkdurkY
QCYbbAKzEjuWcOdh3wXzTAG8jbGf/VTvrLtZ+21ns1cTxK4GpM2ZSyKQMNAX8b9zGKZhXm4fqhSS
gvmKF3uXwGGDHC/EdBEiXfH8jmWCLOWewxPFBp9TZWYPZDjY4NIPysbUsw1pUIqFKUcRb/hobXm+
GOw1l+PTM+gcpsw41PCNtCijmViF9VMkS2cZFmxQRGE8UGOKkOBFcFBRMOt2JfwY3BOBPNVYheZv
IK16TUcBPhTYwg0i05aaQl+DsQLlzmJ0er+lNtED4farNBhoJvCWzVw8BsudFO+2g62pXnBonw1K
/XAW5AhgDKihqpnkO+5QTSmfjPqW9KBPI6DINLlJAwtknBLITnRXWvwxDcnXiZFI6x+99Cy7wZdp
zzyB24gwdzlzN1lhCZji8J6kohWSVWI93Y80kavaCGbpUY9bAytGFjEt8T4oLTcMpEuuperYAAR8
LdJtrAoxdO9ZfqQf0dBLAPXSr5e4/6Alb7oI6wjsN36EiX70I91CydxF/3glTinpT4c/48KZVslT
VYM++AOFP+/T0zkc4038r68DMMVJAtr8lunwHmdp7b3mosZhgLYfmHMCbHdPPkDOcYyt431JUlbi
QdL21OcrTWPs/nPReB4P2/DRwBT4QNUyp3rsKWcAse47waC6XrM/ttRtX93Mfwz2QicJaHaIVpK2
gnTkW73LSzRAFHfIvQN42ax4MFfGgF2En0Px0QcXny/ffbv1G4EmI3DXiA+/BtF8yv9Y5ZU9BZIp
rUgJPznHPrC0oiXXilHln9g2oTfE0Ra/ymXHRs6qdDke7vKvPC/iXKVUMOI1LbP15KPCrTar5nBh
+YQfC4t85BC5Di7BB9jURpKQh/UhRvYxkZkt5F0XEg4Q61VWK7nDrD2nd0YrYBw7oAo3MasKJy4A
Kb5xe6qV5q3lo5wrpRczG9Gr0ZQ5YHTcd8dLsAbTzh3K8mlgTVMke40eVolLt7lUzfjPRM6ZeeD8
AKB+iGVl1/paDhpa2eR2YkwUu8AlvMZ7UaaoKI9jnlRFh9Bd6pNFszpCXG3PdY3pA7rf3JVtHOxX
Yx4e+EoE9oTCJ5rY8HeHwN1rYtU53iF8PTDijvSw7L9rCr4ugVyrUGrBMqNPzdm9jndnbbdObBmD
Ctjz7l8of2XeVOutPjERWajknse9Emk1qqIpHhAInZ1i/J3sxvf01xrTP7fqbhacphHe0lkl7nKQ
yuukzkU6joXdZJ0lOKsea8hLCi238i2qQPjPyOPnya0h0MKhGwKrS0jTaJKRXsH0LWzdgcYO/IU/
cWkQyMNDXz524is62bz0bBSAST1ci1WLlk7fTyD7GTlfwuGtHRyXIARrTzikPgz77vJPy8yReRmc
ZVo3MGvvg0qT7w23bpwY4XbWc2sVVayaWxgfC11UDGWZt9i/VJhX4FrFGBJcnjakgvZfb4JmHwBO
ASUvvu4AV1dDNK0dnqjZUsiEeaM5/Q0lN1Yu+rDr5YC1yYIZMr9xQFjWRBqxnkdk1fY+opvelOlt
mTg8RGeUAcuGBRcRG3jROfH6zpfFfsQNlAK6ZMGaLaOLmo7KqzZp+vniowxX2jQhUZqlLvjO5QVS
I9OTHNLreGPOybuVLjq7AT62TRgvR+NFFlKNt2EK9RHo/q+/beqZatju5w1Ha3kgvTECgfjk4Q2E
jdc4NDFGbP7u/uEO0O0uFOq3/izr6UfEXK80FyTEVAweFaFONKDxrdFTUGy6TsxG/5kBLheuCwPv
2sa2ymczgcFIRq6dyNNg9gFPEF8+d9LoTAD+6FdEMEjrNDAMd43JAFEymvsJrJfbPpH0dQoT0drJ
Y7ySDrfLPxGLrtUSkVYzr/ohV9IswwqkCyCsqBm0l3OEW4hBnQAk2R28oWefPslRxHNfhD/yHSwr
/CPh6IGdE/aN3tTwI2hNJjchK+8Uz57n2wgpsYynTu4+K1Q2H/SHQXWzeZfkD8k1MD80FEntlSTu
J3xU9mEZApyS1V4z3OVyM4kkVo5oChB4cZ1d1w8gFFbyQbAOXirnLga6BO1fE+739KRpnXl7iXLI
ufkNzakSSuntrPwaz+DR9hsZSUXF7/rWzLW9AP6IezkzXeFLRZMr3nrQsS5xu7RlvW0kGuE14PnG
y42l7QZiuABswjMuQNU5gktce1x7WYJgkQiWdam2lrIM0Dv/Jsnw11LctNn8RpXIqBQ6m+soeW8x
DFujSoIlTrX5gJw7rhfhBucSfsWkXzR//n6GMO9TR42BbfyPtF9BOBZNnzX4JDOV3IGEMa492AGB
Ah1YFwml3LK3EE25cuNutrfs6h4z4sPzmNvYkK3VGIb0Vq89QOf6okXDVAYGyZRD+eR9tirKB5Bb
0XZQ/VJsDAkxADaMSm/K++RCYrZpn5iSNLoSDB3PnQBtPfHqHp4H+EYo4eAAWdqvlsiRlvR5ZsBO
724vkpJxLIhlvwuOY+hyxznwAHcgZOcFoTnnPt7i9oct6qlqTplirXpIKKQJo5iXGQzFSUvkj0kg
MoEUhlHcjFAchi1KbLs3sBMBI2wdCHaj5qQSHfjNxEZqt3VffwVENT9LnIvb+jjmEM/0tkUhRgsk
MChznO8iP0B4tsHLjGom9h0BzEjcMSD8WgDSa17nE7uDQMG9peZfd3jwvTrRL1hPm+xr0fgvAl6Q
1cPC8j+Ir5jXF4lPn8BMuyIOVbpqZLuEfTRQ0yuxSgwr/la10W/w7PjwtZDCr98KWMnCWDZDrPuW
EB23ZVqr56C3PGpqR+kpjwxMKtInz0sbkTiAcpnqPyyxDYNUhoFXhtToo6co+rabJVixnCJDiTH1
byhv621xEFB4uIGmnDNPrnEsHyfDbHeqLcQriBtgboUWoYFsDR4U1aEMMrzxGC47MhTCqFAXxgW5
2ts/ATnTovoVtOT7I80IUNZHq4Oxe1iC9nCcNCClOXo8CWS9WNEvKzJ7XnnkQHEKVO7CDKWM95lB
FwhoE47QFWtMyso9C6j7yixmm2j2J97TGA/Q8KJF7zWt1oF12r6EHU4H+kl8L1s8ufX9XgzNstpK
+lAfvvYY8GKVz3w2F34Hwnbhum2RoatO6JCJ5f0Fdefq3fmikSZKU+5Ssol9miu1CuSWaMevt1aX
dfw0+tNK4R6GABKiBTsEWi0GNJBwTSl112RgN7R6321JmZ1zKafvGsHJmolG9PopdgUa+Vl9CfH8
JK5OQpdb+FBDV8vOi1mnychzGI+NqMdEU2rMT0AAIVRUEPcZWQfnKGcicJtbdiRAvxPM0eB267eJ
ZeScHcSlruhEUi7JxcRWtd2t7Boom1e10FDNArPZsgh1vNVedJIXbgBEqAgn1y8dAJd0pj48mU0J
v3UB4AYZ6aahm5gi7tmNNc7aLpzVZ6+sn38RpC+Gvo2Ji22iNkuaZJunMhC0eHChhrqQI+Mkm7sc
6rFlmFdh/yAtYsJ02WbgsylUll6cu87QLU8CDf4wQho/A9iNmJieIzICLMY38gkxu0ZXTa4uhdci
kj5FJDJQCfC/65ZodRCIcmMKj8/ItAkDARvUwkoNBlvqqNbR+LbJ0vDGrIdHSUn9SeekTyX1IO9v
XW+EmMuYUo0X3td+Q+y1lV4BHk8eYzrkD3SudNHn0WfMa/J4gnUhvjzMYS9wfugthVlTFXBl3hhB
bJS/f8BEYRm7tCBIbGRQ25AI/Apwx/mkO2dRm7SzRX/SOOGbbu1vb1cwM+2lJJ8/eBgIrlfrS8tv
DsZggso3kVoeE8YkLKPYRA41k+jfpErEMZGBVri3GLZt/VJrOd0mYodqR8Nk/Obt92xXzW9q0KZz
KJcZbe+HSCNX/rr7JqliRY+KvqqXCad5cDTXjSK7hGu3LSVKYZzRwU9ZXZfWscX850+2mt6L1UYO
FDdKjgQp7iDXASmxqP3QfWR0oV22m28gSrNfr9ajK3kmCzoN03v0jXkwYGNzTDcPkMznM8eeUHQF
D+WvwYzowoj4SZH+7QNro9uycvjETAe8cgee69byMTHb5iICY2EUK3g/98L2u8m8vLrWzJiUB1HH
6CxgxyHfZuF0/0GksMNfAQHfEgJJ0Cm7xPevgfIc2oGX7a7ShXq2tWIIqUEtxVAyWAO6GPFBS+PZ
sB/jkAk9d4dgKT8mipaEgk01Q3Zw6AXmIym8MyR1bXuiOnUa3xWWICEg9avEHkx7nSOjQkY/V5cQ
jYJX8769/tJSNw14LDQ2yVeFa0gUQCom22eb8+fvaFQ0Zaxg8fIw3Wm1MO5Z9GcuAX4nPAxHKVRM
tBJOAkEw1eIrnMKAt25HHeUVQfa7pDDBEfC8EqMV05b6S1Ksteu5pacqNlcY9ljqrQy1BQnukPgS
ImNVuIOF4KkiZUrwa8kOy3l348st7bi3G5TzjWtWeNJ5dSvTmymb1syMKE+Ljmom6opixUrC1aQm
+ZfadpjVfKTqZJcMxg1JEPMK8IiRDpNqXwCcdJan4ztt4UPo48iSYhq6PGqol7rvdEq0S+IYXtDw
3HboWitz2gOGAogmqdM3FkZ9vD9y++mrG6v8fRBEVzN0Nj2axqSOYE0fTalrK0qt+Qylyoo2avVj
a9jHZT6H2sIQkYcOaNmGXPqEea7al7gznmT+2pzucPD+FDo6tCUqPwyC50A1cXEhOL7EtPErtnhO
qKA4bAoLI24iN4X2phqwJgrvqRHXqzKJa1VI/ezXS7Va9chGJnLN5HrC/x6WpvtntC4F43nVZwVr
VUPsPYGDIhIWZpkBPaNjIawY9WNQjXgG7q/HmfjaJAESWo/T12zRPhzkRhMui0RU3idiBcUMFrYs
i5qpbdOhao2x97c5RFl4IsgSxRGKBhzuJL1OD1quufh4gTJOquu/ASqrz7dOrlPHHxS2evfGdmKL
OZRUKW/fXDgzMdbetBLk3Ba/q/MaoqhAqYkCdVQh3G3tgnCZSUZwvpfsx7oZPo61UcDzVg3p2o/F
VfmFzvFx2YU4O7FrvPHd7YTyM7dAG7bAaHBDKy9EOTSlVqQxtp8JIV5D3PT1mwO9TWBmsdJkIB5y
TSvOplr7prpxj8p2zIODNbckJo2Vcc4rsdOyLi99Y8p38d4O7bN+Fh2DPoaMxs5IU6/HQm2sAjvn
E/P558EYc3UP4jUgBgNewi9FarT8mGk+y5fDjFCZy4RXF2DR6vVv5tgOJptuJNIlgeV/gB61HEzv
UMYeU/Axm9SpGWxI8eknEpMBukDsvApt3VHZj92t6sjw5IpQeBfZbiykrnr6Dv8lYxH9Oy2BbmQp
x+RExs402gS2EafjkAlP+vx79qWQqlO3yiCCOzl4SP218otiuo+OV0LDqutY2d7qsHKMZSUC2yvt
ivi7FdQkoAMKIzbyJ/hn2aqb4vbqFlz5O46oQRikcLLxsrznbf3h4dg/X0tGcwVzHSNqUr1smVWC
/SjBkxzjSZ7uiviQfoxO1PcybZWujvcAGuNi8pDSGoqlCpTW7qhCrgweKtCMXtCq6YOZb72K9DdR
9+JU0gifsHV8JThz7Arw/PX4th5MW/NNQlrnIQSLbY71+DhQssDqQymnbrZMNEoNuBUk35dbrf5K
JCh2kEIw+3Ow/7jgNBp6VYifVD0khCKYCt7QRcw5xiC2/3kmx/FU5Wwg7alBJ/ZwFNWusrOzqpCq
hoj4eNYhBiCjEsleGzB9dfKrs6UBwCBbEmXWvaEZ+ZyWwn6+89h2kh8fAgmd+CGwiJf0qUjB3LVS
uPFlWttiaDQRxnTRtHaBjLT5Yb/2EqJe7xXy6eauYubukQM7WTz7WW/S5h8yw78owk7MiD9galJv
QXiYCcKAbI3PGrh1knGuPt6VsGMM1NquYyYsEdMjqa/v0z1Ur265w2FUuV6VR4WKqdlDznc9mTl7
Cv/tI+OyCMzlmzZrE8De7uOXdZG8cU+cHCjTGh9J6hqxLlcbHd6cLt2JNEb7pGFiDKYQ6FGhI/2f
D9c2zv5UAu8bNM9U2PV9Qzk8j7zLMrKU3QBFaUCNQWc20uGy5ccviSHeMjWhxp9ha0TUgod/TBj7
zAw6//D2VgLuVyzCpMfIiTDtTdPkALCMXHvlB7FCOHBeG+9MvoGTVytVCIrpQoZVJXmDou+lQDEk
s2OJ87MrZn2OAAxz7uM3q6rzJzubTrWrQ/HDsCNWM07/AzoxEpNK9aC2qyOxe19TpN96ubuZAVNx
UnetxT7uT5n64QXWaimRSLB4A1ru0K8NgZK5x0q4Wsb9m1KNVlWfh7WL4aouP1wkFZzA5vbaEXpJ
czcqDQtJnelFqcwYaiIaJRDX4qZGHrW9dBANuVKjiVlxznP855m/QaNq9orTYJvBBydjCRqtyMpJ
84mlV4I34GVHriLUVBpDJlNcsEuTuPrJYkDepE27Rbuj6H6UkJwuxNUbbkFtGQ24aAiX2mPVV1od
JEsy8PI1ojSJERGtJrJ7Lgu6C787DjhEUqU7lF7zQrtMirXRBsp+8cZTE8rQoKj/YQ6BZmdZcyZ6
SetXhhlCcRvqTby+iu6RnhcOGwtq118cNeW+P2wDa8RzhInHEv6fZiJxsXb5P7/WoKO5p6CGSRR1
//1+Fk6/Y7lUVV8TeL1Q4K/QX+ABg63i1NjqVzNL2eLiqUHWH8Uo2ayLx1p2o3Q0Zb0n87gcRlCI
PHbhaAoQp+ONAl0+4pnxkc1PF6urqtxEBVTOllevjnASbmogo/3dxTufB0wXBqPSjhuQCj+FhvLf
elWsyc9ZK0R/vnH5tBf1q5kClAhw2qX02iZ+NYAvzoaP34kYj/LnFahCX4dhiApCfg95AtCyyoMS
7vsJ1+xIUe6ecBfhMEsdrNl8fyeHBbqKqav72kzUC3wCRDYNCPKRmR2b/umeN+Pu6JOJUdTNSSGp
jHkJBnvlL+8togS7QTYAUnC2pAdTrATE9lzEH/QQfw9x1K8768+A0iOHh8Lb0ddIYjH6WxCqaTuo
krhNyowHQzSYYDuamTJxBR0VTDEsv6blA2BhX0HlX+ydjDRc248i0EnlyOerZutM2VpI/oUYh2Mx
AzxxoO3nmfBb1WAqGmvTpKvoISjqxRozzcv/B+EObw/CZ6dpWocHmIhgLMIhFZf25dBTucNO0v5A
UPz+5tVB/DK/JDW3rKx2fcl2mrEo1tNkpvXFIj9dlpcz/i0lTsOW3uggvYUWK2WbPvcYNQ3GNUmN
I4LQ0bYPO4cEG13pPfum28vKgiQ3XWrWkI+KNN0XJvJ6voJQ38OqEsqPgoy8FznN8g+Eq8KBgT3t
bayY3pPV+isy1dF3TlEvEJbrLPh7vXc+9DtSN4zQKAyvFlLx3DRADWYQxrAFJCBTy8WCTQGHyxXv
Ow51wzeT4AoOG7DxWW+fIrT7d4VLJWQWOfnmoxEjOHBL/AhmJx2ML3Lnv17sR1iB4WBnAyhdw9Xn
4Eoq24BgA0+b3ZiSoIiortjNEkPV8KLDzs/TY3934rDKauiPSK1MiEdgM7/xonCbheEUksMxiFT1
oiHOIecpaZrxUs1idrWlDRY1joiK929nCXtMhETZm5TuNczsH7+eSU9tTBbTeNTpGD4DtDg3kROh
CXeKLLNA9wC0oE/Ox3kOAnjZUB/jMz06lYd9vFIHF/jEXS8ui3QZLL12ouUQN5DXxnd0coKdr+rf
SskoAzB5kDqmHWG2JYqI6EZwlwEk7UtXYLTs+pkG1BZMQhLostBGi1EhlfsNhK5yFP6oC2N5kV1H
pZ7r+g9iXA+S+qQ1cvCE/AeV9DgLPXR9NrdK2pghvd71nJwVVmwfR9V/W75v8Zc5wuPIYogfUN7q
A3xbI9L3aM2zGGXGR+qXzdK8inzJccW2Yy5kMb8SiRgnPM2vSDXO9XyQMNZ0wcfMs1SvNokctqaa
eezs7qjqw8hV1VqsRedCegYgNLgPEftZ/+nUQBTR8DmYWbjizZ4hTS4viJfJoawQOEHvqTwAjC9h
EZqbDvWZ7tl5IOTjvkNsRV90ySGbNvqll8Qw6PoLcTx99H3FiyB4PbY8b04NNrMU7H+1r0PqPym1
cZejfL/Z3LDrgEIp6q5YcXFdq4VKlliBl3ErOSFYiBTNuVMMmp/w79EKG314vyCGI4lQKbAQyar1
qKEutDXCjhr+lQ4XqA6TQDgQBKNFUZzTio2oA/TmB4/PxisHeOoXi3ZuSEIR7IR7iF3v2TRHCdMu
VfbNtbQEAE8E/FjhTPplcCklpcnMoUaX9dLu86qdpOQOLOKBUuyGthLWlZ+5QPRNV06+xOFFVa4p
QxaEVTszj0UY+TC1IyH8Scti2pIf8C7xp+Fe196fb9CVHFmMYb59exzhfwpEC5LD7cUWmp/SA9rP
krZ3QNDVXtW+OV597I9obWxyaxmAjW1h9ptONYjeJUmDBsI3iJ2Xg3Vt6/sHE12x26umCpCAMjMj
jrrCiRL0AK6Iscg1UZJFHKC72MbWBKkuw3ZYLXucEYtJGXuERnKHWHUkUrAOSatlPqJ1bjF6NdMc
wGE37/icP6eXAf/rGAfDICuKP7p2t5wJZeShNRpJ01QcAeznwZZ0SGXBKcStDEKXxTY6L8smf4ge
7Z2/qod8As5eIPd3L0j3wFc4azCeI2SJBlV0Xoo67iqAMSpDeyTtVz1juWSGMYGDaxD2g6c92fdn
tXZa/a2p6JioHOIwIS7+QIoCCnFN4cDssz8u4+xBZ/qz+Xt3h1Og2Z83kos02cDsw/n8LDhFpE7f
NvzFqAPvq9xEl4/tIPpV9ji4PQZeXv46pZa2weD1CyrMPnHEgEHwr692ORnr7ieumnw1daGc1KGi
dc1XayiX5fhZH/43F5YmiasauKhQGN9eo2Dv517UWZ3fq0I7xM2wtTpFEHH0z/WVsTzkGch05aYC
67jEmSed//xg+ckoIjVdLXEu9KR5qaFTWZnReTrb3+VEYJ+zstdMC+aY7JwABKnmOVo+qkV65WzF
WTi1+fMMM6AMgG3MmIWH9Cw2RV66wZbfoaKf64TBUnubgMZOkbWIBcP+W0qU6SRmCjlQ5TPg9m7b
AZk6jEpP0cn/7mqmH2VJEvbYwa9QkGJr32HKmMXqkHZaiDtLcV/QD93qSKQe2ZwqOjn7a25AIBZt
rRDwY1jBszgSIokkz+LYwwUbrCsA4rLNDgAPWyNxHCAG2N4k+KNR/aLe+qQ0j3NiyuDmrz2DIOvl
1mSwBa+/uDnLEMvmYDtaqDNWsN2t6CkVgEz+rBjTiNJsdK3a54q1JdNH0BC8CU/Qyr8pI/RpY2Gn
G5NXtPYQjx3E6KOXGw+JLGSxvQKhnSfAyuWh3rgSOPzuQEW66rmB+yDdI0WmkV83gl1bQDF20e1o
3+U6C6NK0mizGmHx3fA09S2rYUbLPoa1lTqypLYI8Y5lPTdcaD/mEwPERHJuZJoY4fMiBrZpJ2f8
CIzZ+7Sd4OGswEjwgDE/t3XeJ6i2Z3smPJbJy/+mnODEtiexW8iMklf/OE7ID6FvyaBia4sysUg/
nMkwf8Wu9wTiii4wsvY1gs8t2a08SHU+TLYpCcQwW5Kld+8OkP8J6ITzc6xIXdeTk2542laStSSt
vVby+1HJjpUaUd//W3N8KyIddSY4uNdAZaixXPApg3cbLVBWr5Kk1c1hDH44gL/kGi1V6b36HTZ1
ujfCNALE03kW+p2wYNfZoPO13VO21bHm5kM7DBeo5GSJ5EN8wkiQ3/LWDUcf3atiBGtJVoWLa3k7
9s5K54cBER8NmalIBm9jLxtRGxKb9tVguuxVyGaw4WNyPMxouyDVtbVZQ6JL70rtoY83f3G3Qk8g
ArEXLi4p4akz6YkYvSgAF40GJ0/0hqUIDFZB0vw+kqPx6fMc3GZnv3OEndcqN9TTplEmxf7xmkFL
8/2cBaaWpwdcg5jM9aaLtnT+oHBrSZqo/18egbcjNuSZIKQr0uh+stNGnSkrzyTzgPACel7MgRUa
mgkiodHDlrpRnHjJBCTQV65gH/dzm57+LDGlVLjWEGUNneF3yClt4YDRMRDCcljzktZ0UJ6tL0Ki
+xAFOpG92KBE5XQA6SFKOmBE9h7Q1gu5Vhfgaxya3pBGLdO1x9lUt84AcprYcG+SV+Tp7RXmtdJu
4gAMe5i8IjObPonaR5Vish5T7lKpkq6JUsZvRBFE9nnFLe1gGAkyVjUi+Wwp3h6MLWwwcQzNBhoR
qKBHHd05zzfoFLQnevcjTMVE+HYudwxmH04uygKXZebBUnwPGE2wcgEfhPNJSnGC9tFtcHZ65Bkz
69TWuvScIjgqdj9m/l8Oe6KJs2OGEXNAu7G63BpGObQsXrBnbsXIDPbhUuMHJgT33PsNKbfcFaZL
Cdo/0KSCg57JdNJoy86wl1rhCZEFdNxH/ziRXhwfeP2/wKQOh3q8kb9nOntRJuYJMzFJc7v0XrZd
FzmQjD4XSUSvtkscgQDJ9wubtAwIdvcDTbK0YCwSuu4WvFeULI6DbtRO34431uz6Hc8I/FGi79Er
T4QvNtbfU8xLY61F/uHRSYvee6NSFhES8yCt8O7SmOJkaDwWuoxfkOjg4fVXhlqxVJJzGqt5CSBi
/UBeM0D/5q75wmSFInVOaFwM8M8OrCSwUS9p8AecVHPHgTmEp5BzT6VtVliBjbF/rt2MClg9XF3p
BG3nIa/kDyH6ubmyx/wqt87q1U8lh7CO/fOePl5mL0hxMVA7s1QflxCe3iSkbBv4IQl80wLmeMCh
1ES0a3b2Sejg95PpsCrIhkWvJzAn2zA023SX2C0zwZvRtJkrlOx9WQ/VSkBbERPIE7NirW6g3xFl
m/KXOaxYB0hI9+vhQ/oIQKsTf04VO3sSyaF369vMyIpW4rsShHldtOtDUd0kY92/73dx8JdeNSTU
TRgg8HAHZ+RWGMOYeJ5Qltt1fwKorCc1EujS9h/wcT9upokTHd2LqHEZlOJcwLyAYn+83w5OvrJb
/qyOz7bcLbuqpom+1uw7YLam6s9Gdb4cNSRMF0CzhtBUx3hwex/ZyYVGUE56Lqtnqtt52d5pL3yg
V7i2K8Qv9aKt3u6Zfd2bY7yawW4VPQIFL3ynE+a3Q27aNueuVvVtb7tN9Hn9DiPMRefat727iRto
4MgxuUmnUg5mC81DgvghnVTZD+ONg8SUFE1nQd/rwbM4Ef3DPW9sD9gK/NPMn3Y/nb3r0O+SmKqm
fJVFgBHnxBHT1Rd3Ohsk5QtQH4aP6iyUn2Z7rgafNZfFSjp2yomtrmC2b+om+bOPHC+tbKyF9kLe
S39s8k6zESsTz8ribsr7XJd2F2BekyCnsdKYgTWlS0Vjis8RwZPHY60CXr4/CV+ekcMU1Jh6jBva
YekdcSq7D74Q8E0a1ieFHtLMYVKWQb0Ovl+ZEZ059HiDDxCsHsnV8lprpb9p0NGrQB3xeU93CXht
4xEVCkDOmIIYAH1UPuQ+Wp0YSbEGb1BM9zGM1v52WyN/2TKXY/VpSIQslI/0uJYs5cjJyF0FbiE6
wU6fV6mtJfyk4sZrovNRSObFkaEzvE8539xz3SdhiuZdPIPqzoIX+qZf2Ed2lQHn38HKMxuP8Q5J
u0+rb/cDHqp9E7Vlud9yk1kWFrupWWT0CXDprTrxELDxKx5jeRsAkNdAnQkfH5eTwu+DysT0hUKY
ko24USdGKjyt+EGg03mnH9O9B3YSMP4OZH7uUrfgP0Zo5OH0uIgIODlyduOXTv5Y0OKrhBx3dXiG
RppkOfXtghMADkWV2sbAXmzyCGeJBy/GX0Y25i1ymZS/15C4qY//XX+OBuYw5luMEj4dbaf/J2Kw
6MBnnTd6B7B8Tmd13n8Ct1wx2Txdv20QKyiW5cPmVPWZyZsJYp8pCPIxS7f7E1F130jL0kly49qJ
IU0MN4ko/bf3cRF7mbhGtjbXq+y+YlWen9MaTRpLVMA0S+J3x9SrOA2wz30IUMaEsZOTDio3j7Le
5YzqJjiLjk3Dz6Dmp2ApT38h0PcihD83tNWIVnoeud7+IKSPj5V/6/7LEwa+ec/pe5bpwu6gGYD9
2yUVcvrpT184+/B6sACBiUTdN/wEYnQGrsOmTrnFmxvmTkvxh2bxkqNEdstVJGfsm+GRlKv7hfQ2
pifZH0v/Vw/yhi4tuOgrE0xL0Njjg+9soFYO4MlYZ1KPiucC6guPkUt4qUwHVpZIlfM0TgfYr12o
eKDtWwpSxnh7yEBteHiZKR5B2z5sW9gjHaNlCzkqt4MhQHafePB0DGX9jIFI8wQOtSnuGxUhRn/F
T3bhege0XSLbnFouYuQ07GSo8CUoNNdo6Y8Qcg+KCJLoSUuuXgA9c2lRVccG5xLIKpYiXOrmGV1y
0BLssGE9wnpwBlOQuSdgCruJw0zSZ/Zvcuf/Uz0/c/mMTCArZyIEg3Lu1aIHtTXcdGG9WU64/lzX
ia35lsZZ/2/STu1up+oJtnN6uYK+7VCaVg3Qlvkb9xxJY7owVVuYK40YNklV5djz65zMxJHbMFbj
K7Ydoj3WepYuZ6EfZhdVVYU4N01GLMYHDiAwjJi5On8xp1OzqGcQOzyuCZtvFW740Zek3ORY56uo
FMYwkrHlXU5Ffk2g+iWSIkCu8K3qwDtqkMqi1wrFvjnLGqha/Wbth3g9fX/N0OIzyJychT7wU9kz
qTXVjimX7DHTID8aKnr//gDciOTk7SALfkYkwPWgFX08Qd31EAT1D15oadDfXsBxLTaJUC6qf6ye
AD9OFgHvFnLx2hxSWXIrNjIT5Re5gNltaFLLhJo68E2uGgYflBibBLrYFk820rl8dbe2WoyOEhVv
pRZRTKPzNkwPJvD3lrlID3jzXsQz1INnjepo5eCke7ew7M8Bs4N+RbdcDw7zkAfe5DkTbkZ3LMXK
KVQOvr9CgCFmwS7IJXTHUyoe/sJz2su1Jhq2RVa4Cifyw3bWNnPQ35HvIj/lVtsUKCX6vXqjEmFc
PFKaRwMzTUsWi5jV+/XQLU4ssCA7MhXGTWhcQfp4FOZGvoo2tu4MJRmQTzymt+j9/wyKbpJsZx+S
OsWZcBgX3fK2qUJF+yVsGb5+rUysUQaPffAXalqebySG5s7AZPBF+fdd2pdenNBhX02kxUAoCM8O
vyTpflpQl/S40Gsm3cuhDYvPZPwazkEBgQX3UJNT7EWAIXABMqH9luaqRvNk1K/fENA/Xet+5kUV
qnE9CG9Zybywmmjk/GE8N9YZld6eGbXnGfW4KkkeqjCb2N95QUqgZumo+Jw2mKgfnojXTRngzajy
fUeh5EWH8xT+IOzoDkjTTZrojiB9hY3TNTPtqOps+qcCdpPCyteJy0TNvuwcAQdS6GD5TWruZ9Cz
R/WDwBjPOQaOpQ4ZFZuvmSRHsxiWh2pKE3qh+Gg1nieeTrVn51PsQHyv1iQADiYxgc5PldaAmXlZ
K4ilvePAMM9Z+ari8DjZoncJ3kPKwD/22tVjbv+qU+Z4FME8mKTnOWvlyy4Eo2/0Y/aUSxYMF2qK
bB4+jyw4PsUEtcEnqw9aSK8mDQVe94tBLg+eA42WNlYEGx4QP4LuEQMZUnf7gWDIwSIr00saru8z
kdYTVBtblQVvEt3X6McGJ9pMLwsjXrJ6yNfUAUSzDZkFoljAkLTSCXMtT2WZzr15oROPL8HHqbUq
5ARUUCs9qYAVYXJ//aCOVSKOy1RIXN/0XI7mQozgQdaBp00bA1M9UEa8Z1BgkKWDLwUeB/QKjAHl
NtsQ3fWQKjSi3zuDTe5Aw2RjfMWvFxg29Lp8W1WLZldOEQ/kJtcwHzWxDBcvAQlnf+E8jnkzurKI
qpHeA45GYPa2LD7xwYLESFC1rhSorVbviXi0uAfL8St3EfVrz3tPkWyX3BgATUlR2QJNG9ncWAZi
nhEJfznxjHvVqJSX9Do89Zim1AjcALYXAdG9ua36BRL0JSYLZ1kA7+KnNXV0TRx/5bR/V3hhzxVR
HxMnmAyg9xTxC9qSvsmCc/ZuBQRKIR+uOzmgnHHgjWi7ibY/8WPyE1ikEf+AkKjSucx0TXG3G6lI
BWZtW6Mgy4oR9yx877GjmaXT6Diuztz9kBFAupW8eqJPLkFBbxu9sjVipj/xa6FzLzECApt/GSiv
SWx3PJXX9RuX6rTcIMS8EvS7vlHs7xPa+eXFOMXQkiTX+crrR+KsvXoP67rZT7HFehMz8cknQeNk
jtse5NGu43bO96+0iIN41hoPeUb4A+qkujiLM8tl2iEgCwTboIaAyonxZr3RdlX16N880uPtBjiu
fUN8AqA8WIfFf39RKWDnDJv7/8WdeIN1V8m/9xfzJM3f1z8v4PgqKPIk2xzlhezp3n0YdcQ9NvlU
sesaoX3YnbjxIFNkXJTRypMjaXlDu6c+TtIsTEBH7j6Z2f7yRUnKkHdz9M4Ptcyx8y/Mo/4kSwSH
d5KldOiBUx6j5OfIUjLACDu9SfymdKD3RQZu8heaRu0BHaWP0X/ugXzPSQdOLckhTXctX8BtnppW
vN4gcAKHBol/SY3dHTKrm7gO1osnMez/5UCtSvm/gZhuW+E5By+f7UYs/zJ+67+d1MSEaYOsP3fo
B0EQ4eV7NfYFTEjZnwBTunopNhZcOaz1xPfr1tYR9yiLLwtRYkT8V9MQkEp9W6wtwnMU+dq/+QZL
ckYNXl9CDBBUHduGPbO6wgJV043t6o6NUwcGA6A60mVq9b6auBO8hDpbhjHt3WXwkue5XGSNNr68
hEZ7FUtTvrIzJ5aCEQBZ1Y5hCPOwyWHmy31jqnb+y9LIbd5vWzTSl84YvmN/xbHHZsf7H7tmwfJ6
V03wz7tWeBKCKmdE4Np355ReYEddM9B9Xgq624dqiy22IpVmMy5bVkvdsLZkEZg9+pba8wEaIUjk
QJLjWm2s3yeMo8DQ01wdxJFlhmAKS0cokJ83snGpCKSubpiW1uZ/XhPA0LiQn6QgLHtiKoLji1gm
mlILYuGbc1AfNVzWTjZVuBEgx7TGkQC6ymc5le7zLoIfGx1Tb4WzYKo8CQkuZGOgUY16r22YG05g
onEBEKDJqPyuCF9c5a5n4G0AWEl2sBSr+QYqGz6iJTQXhYQ9P206XnSZ3Qlr/Ng8HDlMDqLirfPH
T1X5avll4HlmtQwCv9eJNrJzy8zbPit65ZI0DGfc+ZtzsfWQCe9gAgk0mkje81v+75UkjbHY6G2j
6ryTbkjxdNcRTKhM+YL47dumB+F2ta4ZVBhVoIzbUag0O19UsaRRVLnZIitaN4fNmZeVAHAhNRUY
/3c5E6HpaNV6tLgpOR5BTtCZYS7KxEyT8VLlC9hPo3V7SnREHCcRtkKUWPpTr85cIJFQ8p3DYhgh
94GdUf47OWLvHzGVTxwcVEvt37kv3ApkU0W3KBq6aWMKXf8IPVmHsbRoVLo7EbJJOxPZEKyNMuZ2
lCDj1c9fgFTxdx5QyssaCiBDFvlqL4QlSlZeXtWVq3FnxizCwdyWa3AvntfPVPS7ESYIaL3tDDjr
/rJmOyZTg6abHsK9DTPONU2p5XFK/QYanbjKcRzAaEz+B7DzSAh+RjZShHAQY3d+XKcF2dhnotsj
vUEEIhKikOLCWqoyDsaJ2OzjmpL34n+3Vd0p13lvRXnbJMIVrry2Xdmad7iLeGJeSRDaqOM/gCIA
fwRr54C6k22KATHze63tqoHPM/Gejbg3PIMO8P8aOyafcg7pRYYQGUt6e+nwOS3YPkuH7ezgPrPS
OhrmqNBSCOWlISL8pvotBalL3duwa+aA8MpU4kPW9+eqltjMykzoQ2cCn8APo3EIXctikK3hlTEg
7aincZOikPjgZb8LHpRV3ZMmHzl3jlqUIvf1YVnHo4R6TxUd85qlOHT51EOldqh63k1efmni+XaO
fN3YAkiTAIUBvxaf6XBl8+SRzGxCfD9FxPFt1xM0lXFFEeBRjKUlLyWwVC9d0r5+gu/E+0+tPGga
8PPBvl6U5TJ3iF/lkCprt3r4Kymr2qO/pK68uggKbbeREQv3gOLq6naD5xsLuWA+apS+Y7RHsUGn
wmF9emXTRQ9czMPMqQgghincoctI2IbUg3Dyse4d99ljTsMhwRzSfcQFbLaegqcG5TbZ67haWOZq
hM/Yj51vmuvPFwnaiVMBttf10hlQHR0iKEc3lxaFV5ase84Qgv2/3LEFwwaPfOPEOg7N3VkHrtQf
dO2BWrZFsZorx84wZk1Cuagb5FYxfUNOzg8i5A3xkaGIvGPg43LqBuzdRuXNG/gV46/BK+UPgkrC
4e3gDdWsDdR4XGUJkeAHPnLXNUO8opNhEqQwex85yeCQWv+TujL8FjSLMDTkvQqn9d1ZIsUhWWTH
gebtOVGt5nDTkCv2fL3VAe7ShtCnGfrwyi1KTdGxbSlJfiLA7fTClUOdHphky9swINuThSQPmknw
GPy9qXv4mN0ETj02S31JnULhNf9iR5JmFMx3oDEIdQHRSiua2FR9LS6Y27SQ0qpvulzFOnWModSe
lfjvKju/22MVKQoDbbFRthcqKz7QAQP8Y0n8PaR4rXjGN4hZDtn70FL+dUzMEuF/4/IGejNsfo1Y
9eqQU+Ax/LHdrdJc+dRavKo1bRDDXSzA1BEHzdxlTHhv0VsmgO9QtI0JziPNUKHeMzAdgsd4R/Ir
Hu1BKymE84bjCok5Kk6jfvhj1QvfUVZd7Qp54B4BQ+fhU2YTJD6/6BXDrlCaCUSCbUqL1IDxbHUP
n7gId0qUCLJ3eQmsbWAvUYHo9Atm5z1hIEYWtoDhKr5s4KolYKh0O67Olx15WVfd+hzSREU6UV97
7oE+WGXnmYLmOO41QJqwI7SDE/PFoUDLv+YorY/QlCqQhjYBy0nfLM32cIv2R1WixTtOzZFUqn5K
Gg4oOfaZgqVzIBUvq88RFGLVZJh6mQxJVSKwflwYDcn9ogKBYRI8YRR8jmAnruLVpf7E5nUnCcUF
KJ7NWw5GLTzXTalc53h7sRFvkjRADczLm7PKYAbs8CZKedkvdT1c+0UnToKIvzSyPoMBxynr8IDR
iFOEeU+HD2g4SBD+l14bLnJ9eyQL2eE9nt1cUhbaHu9ejeqP9afpfA/upB6gt3ORi+gf6lYj8IgG
QhjQNc2Ml3oM4IZ2Sp6pqXDmzKUIICEZ5Xt48jO4cgngNOxzQZGegc/btsGEtRJG1PEtygalbRvP
65XdZY/8D7oHtcrjdotrDN1xngvaNU7q7uW4NDIqcgsfw+iAy5+G6ekmcimb+aMS6rr5+I1ghXp2
BpokMIynE7lfjJN797OlhS9kVn0p9sLwr9XEiMKZv/G8qyH7GtpiAjJkdNri9KyeOgxwHVf8tyS8
5ob2H2lrgi3TIxQOX4zj0tV/Liki+qBCv9dug5WojEJ8l/t0HyMffWai5a6IJYevNXaGPz1dKcvh
4J2tHlsYwjatx7eEwyPeQIVVC/nUeFVGK03cF1qUlh/IXrESx51Png/pHlzNUwoMKF4oWRS9dGrQ
MPnfJ9vNYtQAwWpDWBQ4pEOG/0qj8//p0DwMjDO3MXvzUqrdCFC0ZBOSBgdtu23jl6rY2B/TVsmI
pG1XwYcS82pTdoiPkm6qq3ySU1JzbmBr6NLHAgguzhOo/bLVWmNmsP7ZmaogUg90HYAOOIhJ6Y3q
cHcY3qt0uoBoy5EoXsuwEaWRttHTc6HMI04rqIMsysuG/1bYCOgKW1x9dTy1AnuK54T2M8dpIZJU
TK70WyPDjGGOI6W3g/kwSpuzKDG3pFVIoZkQZULOWznakWZ77A2vtMlX6bCZvdqynUOn+MBovLKY
0d0JNktuWjdAFMr0gdHoU4AteXs05ApnCo5w2qMtVD1JdtNNToWpnjn3aLQ3WMTNBTUvh3nHe/F+
zQCmKwnoSBcOCllP7DLqp6/kuAFtTfnvTnKPcG99h971vcE5Ic7pCbojbqpN0PfUzMAF7sJIE2gr
BA3mj6RTfPD4iTMrJNWrLNWuvaDfB4yrmsyUk74s9lineANI4sciRRMTm765ffdqXXNFajA7KccE
M4ojEPyxs+77OrdkCMx011go5thYKnNNZykvsUgRdZei//bFc13MdWqBh3ZWOYxR9ai6IJCKTudd
+nnqBmjIx1Uw63cFX7CAJPl4iqQq0q9gkN0lC3OdU57tcOkKEJJEfukN/vOZhzj/JHbsGN+EOe5D
BfIQXDcl/1LvgFjqU/oYMWPxqehktoX3os/e90uw7HuYVVChfL44RjdIQ41K0E9nnHplkcZnugbb
hGkdVU7ivsKXT74V5NK7ceW4Cz/y2W/eDPFyeokdD3nPMBzBdMcPf6JVZT+M4cSUxh0e5KU1w4ss
CmGCggmt66qjx8YBTV+rHf6mnKqxvIBXWxLCbBKWpLriEo3RnN4ztIMEluiPsyWuFBGAh8vHZmVf
lUiuF+1oc0Ol8L+QhOq/aaWTe1Jc+KflwO30GVEQ2T2IIyxZ6nSAL5XY8RCe0vk5tZ+lYsO88ZD9
nclGjrIEeinZyt87A7SHFqbxz/NJLH49Y+Ih+Jm3InXjaCoPSZq4ruWekwWkuEMeBs7IQH8fQ44B
uVQG7ahv2lW/E3zvWEZWxYWpgZezsaN0Pc52OhmmnYLhie3O99aHr/XglWXzb5e/y9kKIeUghQQi
sA5w8h0KNZmvsMQ740pvy8pi3Z3gshLvTfrge5AzsrFmGg72d2iWYVN9JxNDrYVuylZKu7cXE5Ik
0YiMTaJXiXtU7bivglDB1Im0LizDGt+xMz3bPfslKPzYaQOCBlvSfqlzj2W8AewcYzYY1jewhXLJ
NSyJTzv7EkhGRimsbY62kjCzSR4SOlJC5SetVVsJts/vJ00LHfNjOBy23VC/e49qQ5pexPc4wqsu
lHUoZnC27NwDvn9lknzOC2oWAx3E2RgTAZoZNrWKIZW42nu3Ph2793q0IoBJ4fFO3UOYryt+XN+q
QjD5q48C4x0K792aO0Kj5URNgx11WOSKG6x4lb2mo/BI0pZtQoVZeY0WGYRmiOmYy7kUTRD4d/zM
2nEHnOJqbd5ghbsfy63mN5s2CoadCQ9owHLVmEO2UaHlz/a8FzXsJuwvoRmzlhsPxZ58X9UTQejI
deBTQLOl6nBZ8syyJTyq8vGiK96LPyKqcENObBPnJjjasAgxmMl18b6fH2HgHXiCnrbR5SWQF8qZ
J5SaEte8tP0LNjxNfc+A5Wxs3HlCVdYqqvqXYsyaM2KZAGzVKl0DJHflMQXgUeEBAyRxMR/PvJ9A
BnCu6PbdHgYwL5tiV9QVyJpBfCK/5iS5C7uMQyHeeb8hZNamar7oaLnKVwYEHt6fPLFCZwZnLTCw
GErLoBLxPdyeJjItTQ+SoZwjpqpnMJ5Dz2L1eINCcgO5fIhUob/SIf6Sg2OZH3YeuIHE0cf1izCJ
6iE+smavK68+nHprSvUiUgXsfDneZafCtgi7XYaGYGnqz8wIq91vgjKCdsD1RDOKpCwnKC8sNzzC
yepN7NY9TSNG6k4OMNxkWlAafBKkKnLVW5zFF0Yddq0QdVVVrL2hWri2bNA8soyZxL1X7in0wf1a
Zu4AkVJJj7OSKEnTMRxDkzU7JZJH8WdF79aMrqcvfhpUD4e1OkceE1hZCK7gdjUJLRviEyO+Mz1X
1c3Hthuo4qfh9UpIKxr/ElZ8ERNgOMi4luzd7md5a8rnECWu4yxztZaT6rwI3VcecIJNbmxjAsuZ
+AVLlPKZaWKFk+eKedQr/UyWnh3IkYYKOZi/RQ9iejM67rCYZ8fMwhicNDrt2fEs2pXxLMVImcN7
zO9s7bu4+w4uBSgWPJd+e1uXYEXyCreexn3YTTY0kSDTi+zLz+6fzHANh/BUSXZNh/YFUR6KcKKw
SsMOPnjZqzD5Qd0Xvh3Bfr4b02UQMdkItmrsliea0URTxWD/+0HbCt0+jgE6xCeTIIZc7mqiIXuk
VYZTsjUpCdBA/kWO8VHnNZA4rJCJKa00siSBQ6/Gf/M3DuPbeXawWlt/E053OXBIpHn7wcsseEQb
AAAqp+jOhADS+2WjAqM2xwcsxxeMdHQgwJPQz9wFnShnIvVaUx9m4XGHUZT43T4fqFMWQvq1ZjZX
pt/x1bHHmjN7pg/2+lJxaPN02ZERw9SzmfN9xCVcn/IrmA/F2qmVk6m8T9KY+FEvuldDR5L0PIcZ
mYZj4RoJYMU5+7k9pxhByEc8NnT6LqLEL2evB86dwu1BgtuCb2Rn9+o2dzGi+RbPnNx3NDkdF3Ef
hheZpivvSkcV60KqdOKma67hmZSJwmACxUemQvOaVkbNVEjTIJRrdg7KRo7s9Mi1rMCWHk4OmQtT
87FZndEemRsSBPVWwo1HiX+VFxUimLrfs96Tn1TjPbZ8KDxmOE95M7U9HnfXqpRYptalAbZZd5m3
OyLkpa/Xiq/YD/54dkp6UoloeCJAjeZIDgyLBjajkkX3lvA0TS7s+VhI+2bLvu+4siDy+I03A4NH
U5e5R0f1kmZ4U4rxzYgK13kAVTX7gSpPwVimrI4ciyxsXo04PQFIEkKYUCnbYHzVSJmBHLCCAsYe
xOzePqJCMXHhOp1GVzrdl56pXXxndi19NH92SXoKuPoWRX+JWANbbteL1WeEdgBdS0UpzaiESqkq
Ahe2Y7Ayr1ZCSv/j+2qQPdq/jCHNetPpkjIT7nfYVh81pX+FxjIe+Phx+4OZIvzNPosYQiiNBLhS
OWAIdSRXlwE+sHcMAxKj/uu6W1wFH5Ro9jUoRHckeDDzetDK9pTuBnCUlL9cvbGnHDLBCossirgc
2b/UCCNIlN5sRjVwd16nGJ89kPZvwkozCglBx4r+YRSRLUGOh8L7dvqZMCnDfO0qA3pPojYSx7fR
E5WbcFBYjuaRz/KWHBOLy1QnylL1IwVgI1rJZmK7OeVDZlhRHjwmcsdTqcEynhaRrNR0a5OxdzcQ
9VdZNUfXi+P50IrAy1hSZbOSMv2T1wK/RqJrno0/To5yH3FiwZc4SSkydJDGk2WI1o893TI36KgN
8HsbrDlnDN9gdP8qCrydcavlEAfAYUE3W8HdtcQjKy+nMr+QbXGYFsjJXTyOgek1M1WKX7VyQaNP
gZJqwpcR7ejfhZ1yfO+JD96A17vL5vbBxeMB4isUVTLHnIJgyMdff2QyX17K7T/WHpZKS7p97iEf
+dUB4e76YQwJljbZkacMP5ss0YmCvPvUBB32dkYYmTzYFLX7wtxzPyFVbBlmRqPCGsiXvxzffN6C
t/8mBQWgGfNZrIBrBQb3IXVeG//BYRueEWigJaxhderf9be0KC8Pivkco4RpylSMp2pJxaamCVcv
bvJ+qkwOi+HR9BVcwgNy5EU+2J1ykLIVzoDOAAqujZsj0yXnqjlTO7y/6Sw5G230ThW9ScZk7L4b
YDN0M3wHX3Hy27FGkwbM1/xPKyyhH1PoEraQJ8KjWCnRvELqmvbVahtKNVpRS4vYBy8On+AlwLn9
o6pkX2lqMs2L6YXHFb1E/qYSPVZ4I0XHmeUX4lpo4XGYCxFI6f1wt7JNDfigik1Yzm0uRDp6GG3c
Pn+DiGJJ9HRl7oUq4vMxBeJC+4fU+KGBPjJaUUvk3BBwAUd6uU4WWOB/do5PDjwjmGcbvSK1DPWU
U18z0ov+fwqOuyOoxYyN3RPrRck7Z5dZBXbZ6Aq0ST1oyBvOvaZD3eyxlFQYIxR4Ct4IYw3ClaKd
M2SQvj+PA2wyaH4N7KtL/Ot4vHWPV1P681rrm/rrRJTvAWWy5qHAwE+GhSXkTVgd136FiwzRwVgX
Qm6AuF1JNujRzOIMSCmKSBYWs3JIck3aZoZ9PspQ5ht539r0EVyFDzLzdfgPSCcdBCjXAmpxZ9NN
1SM98QLrJeoY2eiquvUEMQpyEOqwSFyyYStPUlL/jCV0bJzAwkjIhBZHTFLpKm/oo/GWZQKPk1py
yPAkl5srA7DPeVtYxChXqhDXY02F1Pez4pUvEU4hvMvg38/eF4D0HBmxMU+UW4ezceR1Wjtj/vlq
Z5Zqj8ikUpEZagVjI4/n1jZdR/lKYMMHHoXIr2VaAx344GwxBdABIvZQ1TuvEe3sbII6ox3LMdQE
LtEEV/qzKRvgHZH86aa4fcAOMCk0VGRYb3A+0Y4fz+4JJyNxCFYEbSJWJkDkL9cuOKTu4nVBqogO
ZXvDyRixbLYJxIUkFpTA1RSu052oB80YUCw2VW8KoGPW8XMGqy1+Deluw8Vazdf8y3WF9qoKOXPN
GasG0qTP3BPEaiYVCuy8MXjpy8PZc2FYH94+GgxIy4d8ULRL/lOuD7S6vIpYyJf4+/C/lvm0sYfo
aN/S/HE/Cs3ck4qGiEYemKBN5umUXfi//ixR2wgQGYRgxnYo+s7AvwB/FPTxiuIaXyw6l3fI/5qC
XvBfA7IDV8018DPtHBk1n3Xwzyiy3IsywPy18Ws/WPLe/Xbvbu2DWcZL0cpYLnfrFvc81snowVnQ
VEpDgSx3VMg4YiW2T3Gpt/E9xNUc06OJCNvGNcwQa6xNPslcJqPXtB2i2gK7wQJPDnVHvcxtnPIr
sKO5wsvKx49uQ2LAudrxvoJILXVTdoIiO4MhJ4eW+CxfDzcP0O5nCuoudy4Xy+i88wgSgOLb7Eze
fWID3OOB5Fpcv/YYXXXkwiVLAbWHSlRvQ47UcMqSgYNZvcsh1/vm2jXrkmYkIBplwMy6y8YuwfiG
25BpfptbvaRo8lbBiZwDlwVh2C9DiDavFciIZ7iwO0BSMWnn2fkZ0Q5Xmg8i7tLsvs8eHcmuYGnY
boZrAUeerKvQjP2x0Iwbvs9SrmCb3NKJTMSVFs0znRgXyol5WP5ncLUWnkr2wdEhV2RPbKOzWFPZ
woQfL10vtX4/NCAvZ3d5V4Y3fBbHqWtGUV3sRyX4vpfTvSqPk/hbSQNjPM3Nn5lMuhp9nfFkmv+x
xTaXdxsUhAP5WLaS4/pMj2a54ucIb1rZdasVByqxYPoKb3RxKcF8HVglwWS38XI9gnb+J/OGi+04
iGSQStmxqSpoR7d0qF35RPaYjYWSAzLqOhY94fSCM14gmb4z4Slztspmxo8Fh1J4DjbfbbiIHZ1c
tcOikAGnUy1lo0bbt3V9mh3Uz5YPCBAg3ILauoIy7MGi9jygvswBLhzzHwsBYdM2anghQ0tzNswC
GlYfA6WsnNqia0QlM3lGesZW1SLqWu922mgf2B6Ncq3M1anJByAn7w5KzI1JHmfWA111rtKelM81
eW03nXhAm2lcjCzVLC9NjQgbiR/eO8k6Zp0pPE+QLbHXnIiZGmoa2Y+/zv6m4ue2VdW/PeRwkdCy
BATARf4482SwlhZAdEx7oL/Wbqsb7XSHnPU16ZxaAxwWHnZLVBohqwBbPiVusVOuNuUMwDzPrXnE
o5yxCt4dVH9CS5ZMKkp1cO25b6esvTabitT+9lovKiLQ436FFIcoPzGINX62uCBFSeu4AvRGQA5T
ZtkIMHh1Q9uSxwAL9HpgmqG4lBrWYFeWEzP/iJQzCBh5+GThmu85NiADpt4B4n2PE9j3Waw/j7qz
I2KVLgvOX1dSdOXdL79cNA75g5RJ8CN6IHaAWWaXBrWkcHvIRH3ILJopXgcJZgEQXQkmpRZdBEP/
EVWDpkhO9XesTN2Ei7INOq++VKKS33pHJ7c3silPmy+InexmIfI+rvWdtni/X9v7MTLi8q3B7Jr5
Q0aUx07qYjcuyT3sgwrB4MH4IzhcyPrJ8Ng+sdfCB7CM6xuyNEVkqWKEW+y2DWHOs8FTFp/pHX5S
HxiEa7xIAF+rmA/h+W1AKLwMRe2GaWM5bMFRud+TTfylhCbgvKVSgsXhTyhFliebsBk401Pstux/
61dB1FCXVSO7hquk4v0h4+lBWw/mjCmPBuBEfwV2EtIbKOCt9YDWr9zyo/lYnH4tfLl/nEsQ3KI7
lF2Me/Q84C0ky7rO0hIGTS91YMvz6rD3XxtfCnPabRMn3j2udX7v5+TjXNvt0gcPXlxb09/pVYvp
X9/O991FGWFs3uctWc135hT5j7DapfQz6pIhgHxgWP+ncNla3ksHfgO8a0TgiHNA2Lj0Vdeq5jab
OXxzYf0r8QOUDlR6noRC0LNRE5lrj9QG1IhCObI5RklL7w/I5HJ7sgWav71KT+IiSSZIthPn9fWX
5r0hUG0E5Bn4cOBH11rjrDXkX3xjQhYwCXd03UdD5F19qtlMSF6VSaCbmvD0GPuismqY5UjBnv2E
Ns1ge8hmVrFD2sgRl7du+o/Yl+itCq/njxhL0TP3fOlA8berhRBqI00zdxcDrB2NQLym86eR3/kz
02SCje8QVSNCUiI4Xrm2GH1nC84Uy0H5YTwsETT/JwK99pueT68ab7tBft1ixZo6nHXcQ7nISzhS
OkRfCE/WPbyL5M8tHKnBWV/lAABjQsQgqzl85ImVGmHp8FgT2pyyPGZX8L6LkH+cvYxH9GjbN7JS
0zFbPEnJ6VN6ppnKddO2velcFYzfazvfeG47+gW0glwNYrVVXjz4a3sTSWGYQ/XzpiECPhJ3V0yj
zbgx0ifFFsAxtVUcG9ineO55DymHw9SnJGtB6iAKs8MlrAe/r7zB81fO01tRpTv++dlsbNje85gi
dIP7yV7oO0U2nPd+fhZLWnXDknOCktMJFY1gG/SRui7vlnJqJLSr5nIhjQfYcqDxbN+5MVg5kra3
RcqM+MtzZiG3SYhB/9nc2wBsu1a6TtoTvbQH4I2ywvlbXykdGRPvoSzv5cGyOv6GMQ3+9h3GYTfm
NnEUsJOJj+R3LRrWQUl9ZdzZYKUgD0ulk9gxL8EQheXWD+we/p45O83N5oSfYA9m4yNJqOx5Wyg5
7BiRzdkmhcWjd4u9uamphKY9sKfsc/9eMiLfBwXMSWEb1o/qDUvIvR8dv6J9HNB1zgtQsx76o5X/
brzpWkoJmc9RqC0+Bgj5mw5IR9KOL/2RNX+1jrLFoa2BfyBMLaliUHUqp/ayj94Bhz3PI7NWHRCT
MorCqzd8dGcBf6a2N4Y/qnR5FkrcSBslM7FwH1kJAjegiyg+WLWo1CffP8FCIr70E8jgBfFEVzHn
d+0UawkQbZVctvzPoDaSFLYI3nT7vwEKZe2unmQkCAE/tTyNAt2dc3332yHfEd8b62vVR+kW+1/w
PjQGk1sihZUAO4CQTezCPjwy4qiPscuIZF4iKraScf/VG3XM11PaHJpwvcA4V8jTh2zfNrHUgeSa
Nn1Pv3e9zpwTna1NsFtC56MqhmpEKTZjlAUSTL1GlVEpYYhlRsPaWV1xAaMQaUuEG/yrueuykE+F
j5jCTGm9hdeBRgm43A4O87KIwLWb6XEMToiMdCtmekyz3wZ3achgRe1hs/YYZoQWUYh2sxkikpiu
nB4jPsObtkUIDsMzdUaQuvhzUnnoQJOAuu1UGm5mIzWtfhBJOOP2T7I5J9zYy88BKuwyrb/kNccf
ahergJfn+sLsaDvOs8cBNPDkYSwxroKE/fEKFa+DKngyxq9eC0mhL2+3ogvOLUwT1vwhk5HFeW5a
k6mWPimxdqdQ8AObZB3eR9oqQByOqOdlaFZ5JjMuoKivg3oy+jAmCeowJ9kJjbNjzFssKB8knGi+
JvMSWAktGn/mChODNndsgxbs+vr8fw9DqdFWlRf3PZq254THr7rV8bYwaW2XTR0WFm3zQXA60VG2
KIFSITDn3/M4CuxGhRsXXeynTwo4g11fLdVc7hsrcEAGHsEsp8nphUWwGRNc8+Yete/pGjJ/TES8
PlD8eptAQlR/cA7yLWitGGiF2TfT05jxGLuIdCGP1bEwn63ehDz0FsfgpOJJTrDF6YB2dO9abqgJ
MlwdPA+v4Vgchf4rxS7l7A6n1bolIbMDBsr2DvvGgxA+DJxQuC9G7uf2St6YcVCLJJYarMnK6uxQ
y/8tj7pva5HSM3v5yZZpHksBw5cYCquANsT/yl/Q3AW8zikL14weWRworIGZAkQBNz/6/ixpXHGn
PyVRYyCEUF2OKjx4Ktqnnp5R+emYon4xrfPMcF41gMoCitGAj+mEG7LQL3rfsZF8R2t5KaHgpOf2
YxPrgEYsi/Veo3nL9h9dm9Swolv2GbUoLH33ZMQBeLRRIgni19/SsGjT5DJqF09FsZX1Yfw+1ucJ
iwqLl19V3SFlEN/olhsQcJke8K9/Ba3gRCa2WNDVv+fl4jcrdYNCbrn7KlX0dSCuS+fAz+X9x/+W
rB6izTvlWHj3gxXacF0X6Iq+j5I/FRkHaGwMrRlSvmXfPSP/nFnJh/7I+ZpGqWdigcyLM+EC3YZo
TeqkMgd7mkjbxGbNKNCONqavImsHKw1e3pMCGdeHIpyeT8h1hqOsxOcQOO2HOnYQ1Nghcrr+TG+Y
y14gcJiBuad0TBfhrNfKUkTx51UpMp9yAYPZp5hGUaFWQanVQTUoef2dP3r3Av93GQiE36pdWXQf
XllDUc9PvLbTjbNIr7GIuEFpItAUkoFfSyITHUCJ5qn2bx41moynAye6T0AJ1SnbQmFQ6KgM6Gq9
YGJukbm4+xwX2xQTjF2jQIjgdcR5EWxpTU1MkKxEH2J3SWKYJsxSCPRFLyVSwTSsyVrINGGwE34w
6nNr5gcJEWMKLJ57Paj5LXP2IyqfriEQEIeXbF0NEzIYHPOgqEn7rFTxucH2AXgmqNgsoprr0bfy
URBTlA9/8tc2Fy3Oh0ba+uYxIVXMIPYOyOAay4gbd24Jbu45walecBcdYaJktphT6HViv7fVaTfh
TROREz97FWvyuOtgrmLzRqbxKMb4JhM3o6kbdmQiH0KBaNPIlTq8LrlAoCRI8AciC8anvJyoaLGr
edH4jSQBKSkColQE7mJOhQaF7WEoauAQCO48SwgOSWRNgd7tboSWiJkVMiljsPLeNyhFVowGelzn
Y0itV44Skjmd7IyQBcQnGo2ywuzmnwtqow8uj812zon5LwIIpiNqS7F3kftRLrOvdco4waW1+N+G
WxEjeuCDR8084Zpbjo/WZRAbAzfvym0N2GeOYHJTJnPu+I+iOQYv8CE3WBlV6BR1qj0lcjUPsYwl
4ZquP/kjLwGJfvO7O7gTcuTEPb9bX+3l6PQh/osjPFgvANbyKMPUYUFAvuUQvXNOUqy361piK9KV
0Bz7N9E8Nl5P5WhAzUEGuLIt/hIsPiY+D9+9HIN3STfiDwb582oDojS3lmM7GGB5Rh1yzYopU2dn
AXmksuy87WMKzfFOYmAey4bDGUQzGCuz9pK6xjxq6GUrY+600+40xIQ653e1ekNe4kZjnFZTC1Bh
5FhBL/r5jAsNbOO9AC++Yf+41XNsfSgW8pvo5bh2UED5pJYxngn2HPtXguu+nv+oHVpgVbJd+LAw
bXYdarlRfyslIAEijZJQH4rxvW8v/qQHVm3Aq0iDyteOEKQ9Kl22FYimux0llZeDll20vLTBBVY7
TD+3i5GohoDCUtAHsSGtMWBdi4D9j9F0/GVKAMkGruC9e1kgW/GzAEr8cGfa3VcpAMUF3Wt3oIuL
aHQ8AVWfNMtCDRYyLSxVhusWnE/d7Yx4I9VtU+bt9QwJk8S1Zzl2tI3ZPHSNRVob+ddjMepX3tWU
MQHM7NpP4ZPoNor9mAYvA0PrnCJxEtYVyspAaIoZaEKciEaAMCCdrsH0s7i0xfcNyyH3sKm6eH87
lpQstixbpDsJ8a8pItJWnV0gEp9LezYKPc/4WNR7Be/enpxO1DLWvAZBfv/eNmGNCD4+wrpvYXs4
twsvdaszen0iDBZkaEoURL8f28gzx7lsq1qxRHiyC2GEcVnC/Fe3KO1ieF0pbFn3tA+5uOKkwCV1
hkYgp4oLERQ70DQiq2aVXtthR8SQzk5hBa580dtsgZeJVQcmpEhSDxkyPS34wEcDYPwQ3HDv0hLB
+0JNvc0+9vVt6kF4Uo9Rr9whP316/qGSj9Zcj62LImHrDQskuebHXtXxE+EesXHsXqmEL4jGi5kR
+DK0l/VjzMQrfwfzUREkHlBGE9ImIvQkxHofK1nFpVRWsIBIJB5cJateYn5Jz7ckYAO/ZELTlup6
LojkjW7+swpInqEia8hc1RWEZ9CV9BeAzNKNQhqB8Ea2Mtr27u0PR5Lqsvs+FL0OxfECEsC62q0M
8HxdXZ58yJ4dWGj21zqqhncUGYtpCY3miW5q4tGWFyJBFclIFu/YHXLHnvLcVaGS8+Rbtba4n2Vq
VtH0fAjCriIKhWMzgjjYUG7/BHXSINRL03bxl5xlFQWM7HJa3bWyPHGRkEX9aJPq0UvfP+HqNw/N
yQ0yVUwfV/cMB3RCo1sevqtyv00NuGhmvRVH/A2xN0rHWIeaYcTtXMAAlrUugmkP4Vex5ITO7p6r
9pI6kSjUeLav+HPaLW+HBahGpo/ejRsQWWagkS+Fpa5bFYny8ZvcdJHZrep5PGFkzWgme2KSNwIv
1v780G9WRuU9RxtpymrkPfBR/XyWt1N8w5s3VbEQ7tSgUPpcGobmKBI68sj3S6L60+bHPQ+kuX12
WqHMznB6VXwr1W2llw5/bshLzaUpqcwL3LiEQSfkBjxquBbYZTykKVgPsFIl5QSGrWKQQ0PjknJS
LpvT2XjfXNFTZ83qNDJAXMuu9mmDNMNLz7fYciQWCVhK1ZIOwE70/0kEPd/EsVLW6oVwIgnl9hhc
CkBuFTe/AA/8naw/m6c9PSs1veraLDt5D3a8inE7SL7UTHjvKPC6UqF0dTXRRY+tooOvsoNeAKgn
/0vUTL0PS99LwRl9vL0bmp0naIieRTP70uJ5Q1jcGCBCOVpxcJg1VB6lDP5YLJizIRfobN2kOjdb
V3rjF8e3XdUQ3dg9a6lkZI2XpYyW4+oWycgLAAuzSVbivtAPdt8mWNs/bzXch68Fut1bL/Kpy0s2
oV52E31o28F2WZaqrq6rzGY+QWhxsKH8VzEZM+IYwkEobcmc7ngtIJN7dE5XA1Mk9R0+D5ylV7LH
8tVL6Kh60UmVqdcJJSmrvjMziSjtUrA0ANkwQ4CxWcudny24eeFit0hLTezZWHzM1baadqN4Kel4
1w/g86vsjw2Mvx3lsTUKxl7cBVE4+D12kitmLqgXp57z+NnJR2fl5o/d8KfK5q8ta24rkp/n9eZ8
rUo0T4tV6KQZIkrFB7ZPXCohZha9Vfi/5npBSmk9RtFMY710juTRceN3NoEyjbcK9mKrRe117Nxo
kTAWaRKklK4N/LPfHFntC+vdspbAUCnUACjrbm3J/sJgHoU9qxBOtQGrZybQJ+ZlYXBue6OEGGBB
vjoA2g91D6j9/tPQYR+Hx1B7RuwQjogclK75c3zc0ANe07IFkuvPem9iLU6KSFtRIbZfEXjb7JqV
zZoeraho+obZwgHrCh+MYeJrQzDK2DDyxTFAc6Dnp8/Vp/bk/38zybWwR5z9iNmHFuqOq8FFApNo
sxIpVcqmjt4uPqjudgO0cwWLjp0SzuyLdK9ZFsTmalD2r8oj1TrBFRcAHJohRXkKopRw/5wW8rUN
Bv2H85UZoTBwleTgFUG9GI5Hjwy327N6hEXQlmr0Jjmpn3yv69PJLbJIURc+Lf+0gkmEHYdC9bSW
l9YOpdHklDuG8sAGSzNnswb9BEzmte5Wj830BmBUQhtSaz7DyKAOS3jsVITpqoWihLQR0QbjdUzd
bql4Kq2Fgn1nABxDtPfcJHVcDckqQtH1BAY2MmTnw8EYj5/+YjlxlNcmSu4F4SDsbwKSMji0CXyb
+PFWhWNf2omfLCDHHJgCErqDFyU91DJV/jR73+hrb+rZ8g3CWu9US8PgxQUU2HAk4hL3Fh10HYQC
QZ3DWjcvKwpuBu1O3df7TOBQMBgOr2U+kq4Tt6lLQz8i4rb9RJs0H4KyA/ZGORnDQnSFxLgpzB0+
PFlAVH+uQU1lbrwFVQOHP2rks9LvHi3VQKKF+zk6lCEa8jDhuscrlVn4JY7G6zRmAfDF8QxVtbk3
glYbv1adJhf61AL/6ds8JDJoekjLgt5Jn6GPszJuSCoveid9N2NBAPo8ZgwtKtVsiEb0HIBilj/v
GvsuUlmxrWTwRQXqCOie9xLUdEWDX3Uu9u5n0pG7Mtxs495z98RDS7/Zua+nJYRcWxJJAQTW3dei
fds4q+Q3m6eHPRWq/WBAVbfG18jE8Ot3oPv1Z9R3nkYQnzzivsdTBwY/k6KYB+dRlRkBE+QE0AMf
4/S4N1jpwP/mMSkHlHeu11AwdQrZ8rk+8TeZ9sR/dbdUrrG/A/UDLFSSCJOxczkdK5pQhg5HZ2AV
tuYus2/I63bXv0v364kyvKHvVUriEWsb9lpIU+dHYMXBCRqHmeQ9Ae5tPNHW79tDwW30eE8MehLt
vDkb84OBKErvfqY2TtoO6hXANkGhIDsAeBM2E7lfiIeKEo+ivCRsZOh1TvrShgmenWJhL5YB2Q4k
pmfohCL5o1xy6j0G5wu2crcr+VPjzRr2GUHfID/FM5k0B/BRe14qU45rGeMNrPDJ9gd0eLg67dj6
vI/RN/KLYRY+ytLzfJFm0JxK6NRmxD6p9VVoamMpGDN0BX4pkygHrjsDVVbMVS4GeGDyxRabFTuc
kG1G0Wvp9yXYL1Fl+J0+mrE5EhssVfAST3e8yOIBR8Lwn4bSetcfMTf7rprPMHXZmdLaTuQsiHxF
vO8Bjvl6XHCxYikR94hnEWvPnIoGFfoERWzFQ+V8prwUo1KtVIDWzmrZZLusuPs5w30JYaezuVp0
vG1AxzsB+IVFZH6JrSWwiWf4q5paO5h4AW717iGue8FztYKFb0PhDJ6kI9UrVcVZhDyfBxK2Sc+h
kQ1nJ4zkq0Jvl8aqEgZ3Rbx4e/oFUqcQTwGQS5FeccYhkO+f73DidswCV72KZDpqJtpQoQcPetF/
a4r+GXJ5ieAc5b53haM5B1NdiKJA+bK/z/vA25TpPeTuyfYjSPf3ua6E2tt3uAVowng30Qs+ItW7
kOloceRMAw6N2cntjKbJH5VJBG3cp0Pj+lWgwrMcbSAL4Q/jtaKjByEvTdHiBmu1HiW8iTeb88eg
/qO8JTiuKA2CAFaiSkbUkPn2IXX0EbRxL/gXTT1KL5wbmEZ3hEJcX+ZsblxoMWgQXRAvRgvUF05i
VgRymay3rUMW9KojiZBrgPeqiyfqSKo2pNgZBznvNpNbK+Lo9K4MPgzK6vB5rupBW0KBX6GhWD7h
VqkkMgyhbc4Ez72UOQmc0sv5YD/Zf21Sy9Cn45Z21T4ZTKKyDXAxnFFWA337RuimzVjXugBM3uDU
O90XkyqZ52m/AItXoVBQdokXg/J4lMkTyPYdNNNHMEP9lZMj0YmV+4aGQqCcP+IC/ZP7I7gfJYmG
IcOtgSnA2Oef/TnBIoaEx7x/c8xoPEbu8mavjHmhj//Hhdl0f/qsXVcrvtKE8pyJ3Wr2Gb8Df/CE
HtHOTp01bGNkRdS9635M9cd7x5H7pUkcMVVulnqs1mOTAELKoEq7xCmB6nWGkl7gwE1FGP9CkNPr
+DLPQI0Na+H8nKLGEQCJz6Fa8yYw3rxEXRlvIM0pkPxSzY5r7T+uA9WAy4UFzI32vg05cTBVvGEZ
CtCXV3yZMYXuEC0pkeS49oxO3Raiwv1HOwM0VsNuL7m7XDp8FHNgEav1sd95Zq/6RUS4W6KUB3uq
rHMB+t+uCLEMY0k/OVDbb44uE3KHYK7W7jVZSPPb+BVr43FUV44QAvuNk/gptOlPcS416g3Lu+m2
kgM5IRG26hYCfuwuMZTefH3VfgbQCH0gNVJva+fQrTF2TLuot5Ogugs/pknt6Ci3ANh2dTc+EXOY
RHV1+vErmtiJesuo06hrf3GdqPvfgsgZ+tt2F5RhKaFaF0uRASJWUNMxlJum6ZvAYkeowXjxrvCe
FKQZuVpHOEyarfCs6bcwSfJf1Spgbj4gQx5TctJywP7MaGvDzSmUUa0VurLRuCuqgvplG+cxPwLi
CzlisuSRiocdxcrXnBkPOte4JQhnEdqtfwkh0q9Fpzj2dhpFd0aLsAkP9tQZh0zMN6c92QYDh4ep
IfuLFnGNgXGSjmxWPC5ZXofBCU8a7Hg9YL3wWHF8me5j10dnX7vhbxo9Bzf5K0g+QuM6xCcIoQEl
71atahB6mwVOQ2DIkT1wE62BKdd9k4HMPXlg83z3382kEnjIh2B0Q7KcUjnPAsyR0FMslLMY0XbU
SlDa/eElL86YkX5/Nfw76fO9U6PykMS0HemF1saxNEoSYzECsWrNyOCTGlqDVI3T5D2SoRbpjepK
IKOAhUiEJltGCnFT4/Bh68k5YT+lui8Eqs7TggK/WUnJ2k5JUTzGCpIAGO+WuAtzGBrxmwk9K4tW
EcHTLL94Ib1nAC0mMPI5FFX/wXTFRE+1ggjgGuDwOHRmCUEUYe+TlSx2eV9XG+OCyKhcnYTFqjN7
HcWzVlzn2XPPMuAQdpiRvkhXKYQmezs6x0N77rqQLhjgLCgKe4kQKiLvnBjU2HF9XHgtPMHSmsMI
kzi5h/mouwWKfFRwTkucy0uRVOBau0R5yMty5tFgGRqhxiyWSQxXRo4XNoN0KplSgMuCrQx+L4a3
bmS8iZAQypz4pEHGoil26FyFzJLb968NLaCBMZQRD6GK0CxtShwYGOfgAzYb0eGtFEoFzd7EVLm7
qDdkayx18JjyBFZO6mrNirtasenwYkuvv3cramsG1T9X2Lx5Jvx3TKl93J7cAuFam0PJ+1rV4aOk
Ec51WyU5IK2QMOPB0USKuM1471Cb0baZ+Zs6udM1VctZ/42gV74w01z4ofWFX3gHocoeDSaKb66Z
KAlOrmnnmzXnmgXM7hFWE1vUqR6Kz05mm5Vf+CaxgANu1BcPSxlDcG1y6FXeQUq6jAAHQoGUw+Ad
ZP+1Q34JHAXm5SsKJ04+Q75H8o6O5vaE9nobbvkzCdjnFeg86Rph754M3l0deEx1Ebf/VwkZSpR+
qrY9TfKo6NU3ps/FI93DpY5GXxVOABbpm1PE7fATBS2dat7xRvydbmh8QyT+UGWGudmMQXQvKvrG
c6AE3pLWsi1/VloUefKKEBIEkmkXTrheXNvWEnkhts4WjX6wqkWNRGXrSf3BwUEQSyikkyXzFZws
MrWSpxC5355RkDjDvkNxhi8LsAOmvRKC6mF+4Fe3/86bZsWI88FEKh6VmlQyhWsC2SuG44aePFmW
UUH7Q2DE+aJKAzta2GFif/7aJv0aAKzqEJbRJ3+pyrysWB7iu71cBITD1OwVvn9WunxrcF/mNY+S
pa4dj5uCSs9v+JBpDzOpb9xr+ZKT24BrK0wsg4l9YmhAcc2NINIUTjngpEW1vzX1+GjRxpbZ8vnt
w9JD34n35PTdE8FXd4WS4l+1STa7SM9IML4T5CjIBeGgbuCERxhHqWZArn0M9WmG7VqWYKWopGCU
qTGOtx9p5R2VfLyjbnDNvPVLYs4LYS+k+OHgjJKRmZ1GtQwXInwuXKjpk73s5BhAzsI1KFZKai5e
hglYKOZptKMeCKQgQV7CAM/vG5kqlejDKQIFBbVpCJlrUgg+hxLHTs4SpD9tL5XJW/w1Rfssnp4o
d4AmuY6ROsbqj5jgs4MhHtAM/1m1VIRPaKuKvaC+93kYjJg40//K48n1fGAme7NjLz3ooVYehKzG
DNbGLIWbH4R+ea3zvHeze/mRZOKw34OMSsCBCx7FW9tsG+KLw2zHZB75L4sd/LDGLnOS624Ewbyj
qc+5orVgUvBWNxrSSDEehV/ahYfZ9KedNWKvfufL8nzvaO//LFd7AQih2HSUfP9++hvLUxUWe8vB
zscFr1CpaN+QFoeoYBk7ulDAtpQTC0JGV6wzG/K+Ng9s1+bPjloNvgJGz8QuJpNXxM072WKnH5in
AgzX67RU7OfzgijtK7vdZl84m4srAw8XxYUOV9OMEd9LqMz5WscvGWsaDS5qPUhXWhrL6yuhtkFN
YMsRUg06xkZ1jHAkuQPwt4fYDmL8vbyVUocebQfpW5cRYFTzxppYOFMyREQLWVDhgJCdBHuQv8+x
SZLHAfHm7jWCvB/1/EcYF8ComujF4jmjOqG4XBRy+ji7AJ8bCvPDhPW6IaF0Y1ZzPHxh+0Y/++RT
7YH/ZX8HSAaNRna7PZTA6AAarOybIZ12fsZnMLK0nGuYAenMnPQco6z/6INPh0xc9KjXociYpJbf
Ecgtwy9sNAyPZ3bCjU2TVPX2jP2GiKAqc4mLF08I3VpLtevzJejTAPMlR5pXrtjmnnr9mumH1R1I
gl2EhGhEgyFYidV0LlqLr25rtqV0TbHYYr0TXdl7sBrVcurZGN4nvAg3/OU/q0YK9s0iqA4PP+AK
kHIwxge47A9AS1xrQHa+Sz18XsthDd3w0ryIwyw9F7MTjnHZEFK+7ZErDt0ZxssQQ9w9O/FH0+VU
k0Tgb9/zSLtTU6x21LIhksV0LVMLGIssz59QyUsVqs+IjfkB6IJ8Ykh8MPJs6IKBeko/b23i3PI2
mqOP8+qf2Op+DZ5unb8zvxLUdkiSG70jV1VXl6OCM0ej0dgqdts8sUVAM4Veu2jOb/WtR8xI0obW
qtuzBVxvwqhiIAEZfn9ZhdFziGyaE6gQfrHsmUg4tbN/EKZxt6cyBj83sjjW0H/y1PDwFXQkIQT/
qDgaFYpOidwO/4hCP9RVgrpJ9YNnokGa8scoAqpn+465Jey1DSbVyhPdeGaWoaOF7DwjRsRpG3C1
tUl/uHYd81pO5hICDVQE/nDLVY1I72XYUFccp7YM/8gN9gkf7Sp3dWVhq2AD0VB2D78pLyLAoXwj
cu+ViaJY+gIp4farwLebFP7Logwo/5Dnhez9KdKnICa4ADzZxqVxOLnjrBqJL93ZNqYzZsYflzE/
5e8eTN9vOQOhbCbAY2HiQuuGwRBVn1OVTqancfUydWL8+TNaoVmH5r4OJGej+XQkm3d9//iRmJ/c
ECh7Z68PGC+CERjOpJko8FLh1rvYXvkJoIyh7zyDGDvZWNJ3jSbD9fT18aUyb5PROHR0dRhPUq92
6qunpRc4hZEojJLlLegURUvVH1UY1KXRmEX9BtgjDLHXG0RWKfS0VbmDzvWLJGsf7ObGruW+XGIp
sImZe80QlJPacVnacG0lgMC2vLXY/haMJsVXfQeJ14w/ItYN2qHuzE1/Sy1jgPRtlofMhn69xpSd
9UJq6riNZC8W2+TDt2up/LvuZW7WqxncKNrxB5f/P4PM1MJ5HFtY223g4Qe3hIRM01W47KRmufVc
5W5yNNyAVOXg5puS734f9B/lOeeIFBvy1eLLtaSNwxQ6ZdN3c5brte0E9LiOU04gUKCHUCC2twEu
LPxWvCDVLNrZlqibdSzHYp3RG5IVJGwY8f3Vz1ei2OeLh0joDrLAiJLiRBl30UJEzRwfUpCSV2Ds
GlxJOerF+FWxFCztCe7TSjbI9EC7jqqmUrfBHgx0eURpjwPaD+OB7FDiJwgRiVUxSjdp3zXd+i+1
2ybOA9bDkRkDfyRGynIxnJGHQSicC4gxNI0C2IOKFXcspjSke2qOkqqQcd1500gURLuTjja8bkhQ
5kT47+EojjC0kF1j/+TIpbOQ+ixy5ISdGILB0ocD6s2MDfyvf6HY1kxjeFsDNacHJZcRZpzViY1V
OvyYn7rTKbJ6QWrTuNke0wPii0G/DCR1t7+yL3WJPgdPFGOnAuJZh2xcB6HaXA97qlZjbdjBA9dU
6407OntzIICqe1aqWxfT4+HvsqNAJuHaMIqtSuLwaH05pmTCnqJGTDFDMVsiMChdIW4T5KWKJ2LG
ofRPGxHV+NIwq4dows5ZcFmNMvUMRrp7TbCBFQTyTXLrGBgOQrIWBW6PnWA1kN3qetRinli1lmwk
zn51Q1mLv9eE/Fym5Ad+CILnS86llojEDqnKY3SFSPS8GLs/jrfH8bJlCU1vcWiJ/rLYWMp/sQwx
DqQLx/JbMfWzNFk2S+/TwkuF+YC9qtmApcXju25qJ64iWHdXz21PgDpFlFj6+uuT+/1WJwlY7gLr
nLcrw2aojG4R2kdeCjRuDvI1ZwLpUJe8AXG9P0enib+1DwZJrpLpAc7v9ppV312XG9Vc6kkp194C
MRj40QPYAcVmkv/Dur36Nr2sYfojrxH//K868eH/dHN2MxWBmiXGmskgngmeBGasnVBXtusBzPJ/
i9jQbaSc/4ycxv+oyE0c9n+1DSr45BSxXKjYZAmF/bVM8qjVmVqrjOjm1EFjd6jKsjUBO2ZiNg6A
OtISaEmHShOEOf0IozaXtfJY6n+5y45yXNU9lv6+UIevyKtqJTAwOrt5ZvmOSdRBqzvBj5WtGNOE
VoEhGFFbm9h6Td2tPTay+PJsgq4cGkOl2u/Hyw8ggrsaKNI6/tvAnr8u2xtxgvdL3iWICS3ZQCaP
gZBeCmb8rI6rJrJ/I8eNUrEpQ5sFHHqY5l1qUvcWxhkPjx/PMBODnjkn+DmQBrWz4I1Py4tIPYvH
837yY/v+I9Tu0FYwf9Y7ZmelfbjFuWTKDjSFUfZaZI5VdHEtMhEH+zmoQJIzP7Z+8kmGEGMLIJxp
tIdVE8YGwhJjrxVojlHQ6cExosToSykRulNVEp+QqZoGmGfinteJQyq3vwQjX7CoQAvKGdqaoA9n
IE/EkWEe+NYT9KdceRFKK7upaoTeL7qz5KEYa7bbDMC+zet+qi3POw+pnaqv5jagXNb1U1JhU9Jg
9icZHkHtBSYYZ8gH8I78EgKL1cifPPhYXpActtCbCheLeay5Gtpse4ontSWfsQIcR7BXck7X4FTM
/FQddKwOKqj/4OiryzCUR6ThWcFV9SznKBbG3CfW2/1zHKQlf5OVuZ0ZbIgeIaLUod9HOyD/EHb6
keV8XwWNJpO3nZlf6q5UGw9edo4B4yXtd3oFWHAAR/CNZaWNxBJr8/Zh+Svzg9O4LGoRTSVCzTCN
jqp+vORbgNt+3l7pTpU+XeB4/JQ1OFsIf8ysDqZRBRXTF43uz/0cT50rPAuHgMpfZc6fUoCb+uff
2Bs2cPPsVnL+lq8TYV+tp8AzSzR/O7X2t+j+HYRbRosohiRosNcFkbvdFomAxT27+bP1YiuJg+0d
/mMuX1e8USW1jBEv1/I1HMU2pGIEyYBNgfOOhpABvzeydbgMgjQ1qnKrEy2PBGOVtyVXDY/dmwBi
vav5pFGljGBoh0kNqysUt7wwPe7B/rBXExmMr4pUhU8R72G8OMA4H0lIKFWINo9VtDQXBQ3VS/OM
ueoEU9VqIWHTPuuofDjJdgH2XP0Gf0UAMsViwbB4KtdlH9J67vr/AekUKBCwjWR6K47KqEu1dVvb
AUEihBODRi+LrbB1XUc5FZfJ/pCnqaEMP3DsWyOcknV8hZLKTBu+LSLBgo3Om+lBPy/ikHEGiLfS
rgddSYkI7QRoexth7OaJkSi3YHvSHsd751QPv/SPToVnYV9GTHzF4aQeaJikOjk0lu7fUQyyf+d3
SFL0ll/n2dkJvcpSjuEeP/bzilZXBgCeombmA/FsdDwZmGeQgAwfyCazYEtmh7cN+OE/2AUlU4om
S/4UsFSHZ67eEc8b2GMQhN/NbtDuOOd1qlWsywuxSqaV/3Z9VHxuKAUkOFbn8PEj86p/K9RoJyBg
PAjPjVHqGKVW+4QPnrKaaW3M6m+ML9G2AufCZ5mW648YO9fOWPBgZ6pIlz1Xew2mrhAmgkmhYo4d
rk5Tz2HpESsNGF6W6TYCpIc2eGg0HKjD47rpJ7QjIUVWH/BIC4jKYjvUDRBZkX0eBoAkXPo9UoWD
Uox6IVppBKBiVcaDGf0/hLi5gcwn389z8ml26F+4I443eh/xWcw/JxGNB1mUDv/9CSXqiNCgezUL
oO39hz1wYRQ2wO5AU2shsMdCVr2eRqBIY+TD40g9v2n3I6+SD4A1OIAnlqJo0TuKemqQXcODYAMJ
0x9gJJ663wa7pwOXGNnEnR90OlMshiyXiK5it7Eth7ZYyUw8aJaD5cB1yztYtiTPnmGwExKpT9Vt
jl6/aSbyotDidS2aKYXMOry9Kat9a8zfkafJrZ57R1VsxwewH1wqgaeq3TVumPrHDPfsJELSmecI
jsOmc58DoZ++A07+4B6lNWg+31f32MW8UcwgesQC2g5j3Kk0SZdX4mRElNvhHAkeLmzY73a7X7Xf
ZQO/MmEZ7HMCS8FPqr/ivBS+qzMLuEKnenZ6/zcB6rFtSYM/6ualpSocNk1E58B5XLvrFIl4PBZp
n+dxhx81q1IQliaOm1Xa9rWchVEvw1CzNixTeuJAUQKSanSrkrdwueetQourfXq7DgpE2zZuclnq
47d9anVil5+uQakUkSCke847tZmCRLl+lKMwoUdmKV+ZVX37QyFM7Wf/fNnVZJqdHkQRTZGf0U77
OYwvBa9nHgPHgu0KHzF2EXTAD4OzzCm154H3XcjIimgWXtVJmPs5qAyNa5XgR/pUG83UGfskYlLf
brTLmoLTt6rhW1/NvsVdcvX6lxPpjw+UzwZ3oZCeFkfh1yytWWXc+mTiiPSQ6qV4YciUo6jYFC3l
Xe1OAafPIbNP2K4iQytIa85QYm4Pv+lS4VWwLRqEdt9PQFg23S/AdYT6Zj71WyOdAmFT4+Fy8fCt
0DywcwyURoY8RapA/vh/M9I+wD3LuA6dyFh0wTUa1Jr6AId7rk2ib8N4t7y55tscygqbv9kD3KXQ
cHTCmUCKgbhk7kl6M284ihoCGAEpZHIcYGJjOPV2PLcDcoxFT3kYJ4ofhuv0cJW85nrTIcV7RBbP
l1XgQ5g7CHXTpGHxaBOAMuvz5yJpfKRis3bdcgZwWm7g/ceJbmK85cApGyne6hN3EDfzcF95gUnE
IJs+6DHi8ZG1xQGUoYttLQ9ajlR9DydcXJrFa0y/XcfeQoUEZ4fH4HaXt4728wgPR6AY2T1hbEId
bNnyiNvbBtYPtd2YOAGZsHrlHHDTNwR4YqEV0+afGJ/3rKHcc8AOta7rwucE5/Q6hFL1RoYaorUO
V2CJbd+yaYdymD7cksG14fvja3lGThww9+ytvEw0Pk3bZbZYnbooAfPIx4Fq9qwzLJxZye6ZOhBs
oGcVAaIp4qyvXkNIQqmJhvw+cAejc/HU3Y3guQRrtVlYK2uAI6m4yM4U/IEFGVCw1tQnrM7B7lgY
+x6fCBsLOumt5zppWWdw3I0cno/DxxQzbvdGpN/oiw0Cc4knPxdUxglUFmwTk932OWbjJLhTRcf+
KJ8q7AN2mp3jHn7Q3PkADHKIdjoNxjVjQKAfTPgxVq5aseFWo0dJdWiUCWL/Npd1CqqObbk3VI31
/j9EeLurW8uDW7VgI609yci4AeTy2lDHi5PxjMQ6GIFQHuMfGGZ8+xKwoJZ3DSF2SV03fUJJ5QL/
TJnibN8NttI9D3uq65DV9ZJbvtGcy455ANCLVQN2oNP5JsbSwS6pCqMxVkpAjcLkZbMYwK9dWBJA
BgmjZgu/2Do7muOF2qnzF0UAtPfuyB3tL9+V3ZXsCE9ce4ZE220H1PwGTwEyaMncNNQ4RVFNkRat
6PjEQ9Z3XqRjxdSH1wdWgtO7KeCYEQHENHyPlSIht+tH4EBVGo+oBFHo0hsN4HH4PF0H6dK09VAu
21DggimZjHGQWoaAXJXER0VrR9mK6+Ce73pvQZ7i3XumZy4MAWxG7UUKXP6/mDrMxZG3jIzf6cYq
Ek9zy50a7dtJcTmXJeo4Xga3sAVwprk9RlsFl7hCoCsx0BWY02/9ArwLy03vJheHHpTfXgjSKzT/
ECItdsRKLoQNF3XIwMC2GQh1Fq7PlSks5aBKDdu+teFkyxw8gvcz2P/8ouyXlw36fxaENW7cThCJ
kFOxPnwz8iHCiwCORjxmQ4FVZLpVDcAvm8TC0yyy8GfjZQfjEv/3JAbwRCSYu0FGz37Vp4z35l1q
fp7ZY1EuEkTJneolBM8VQlX8/l/DVH/72kk+NRH9UpMZ2TtbUuYzY4hlcxE0qFhNowfFe3ew52Xf
eB4F7y81w9FpIMJypDbEb0dXBdLhDurpJpvmz1wXNxJm9lmWRE6WjZ5qD9oUz1hKzdsjw36OQ+Ln
BpHMeuB1FY92vWYzIi8A3QbDhXD/Tb3CG3VVwFVTlKReH3nzCgBb4p3kPCJ0TyKrEydZGxpkuRme
W5hyYSb3kUSWUmyzQv4nQNLVBXeiQ3DvwqdEFRpk7znx2yrpq43J0Vm2WRIFGVBK/BpDNZB34AAB
idAEanuYElNbtIf5LtqSqdcyr8QTRnXNrmlOB+uqwfZxi1KfUkyh0GwZkPQze98rARQ7ia4dIjCC
sG+f38tJ8fniLLEvKjeBUdztI0fig5B90uJij5ZJReTLpjRVARaz8hA7cFQ4obRCmiosfHSLHr/W
s/sS08YID9OYVb+2sojH7mnjGTfpc4eTZUdkADx1LTeE7mQUiNwnzClrAuRdTWZd7wqls7M7gV6O
Eue9kU+oDRdcmCY0vBLCTTORga6eADBz4wcTaildtbgn+ZuJbKQodWnivcrFng52PPKOunZL/EF7
z2qfbZYrVtycLtSbWpymplkucG8qzxvFchDAkVq651TVQyDNYWbSo6ktXYyUn9dXd5nSyJ76NMHA
GDhyzWPJ1Aqm30WYsCY1dEOTJBHlTMcmwzUDzUSP/WNhQjFAf+rhlZ4VjvsFHxSgJGaoCHOkOe7y
WvEGi0+4rLLsMEs2L7/kYQplzd3TINyjwiVP25/BamyffWndBmPyLjZyeROF2/BVJZRaNuppAsrk
yfIpDxjpDC9aU8zFJEtt1367t83Y+lWD/zEAYl0gft+MWte9tYxWHbOqq2WLqWtR1IQg85lg8HMO
j9QBWBPC6UjHFVnElR3loemAZkg8/qpDIFMOPo74aYQNdf795LLjB/D03yxOu1wqBGpA5bob4Ln9
i5K+IxcrGz0XZGzxvDPxO53dn6Yq5+n/4KX/pbyqWGvmOqcy3MorsU0wHRXtD4GumvaWF+9lTAtl
diZ3OOw+4kv+UFeSaA+98Mvl71PZnpG3Xo9y7KAv0jv3Gv0MXnC5yzMG/9bZ3eHd8jIza8P4zFYT
sA0TC5GmWmNRoOnUmNzon8lnujprt2AhKvMlsIMCGPQtiGQkSuY2N2zquTZouZBp1eoQ8dfUVIim
Ft1xpvzktMKwNHJkNTDKJfpIV9r/L5g6hKIZkcxWcQzbQdjXLzuh5Lj+YbZ4E6nQUhuGSPVpg98S
TsxZu6MBtiMbdBotBTAA4pPMRwTppPvOfFfmLLuID9it8Yorj2OwacdShpt6LNw1z3GZGyoPyHmn
H5jNLq78QR33PuPI2jaBvEm4MNw6jAhjq6fE/+Hh5XyXFWaWoik+uF5MPXk/31hStFDS1t/Vdaj1
OiTJCkk/pmCa9dBB8q5WN42uSCNYaugP3IjC1sR99xtswAAxSE6RM8ypteKU2uYF3XGwtNgKYjWP
5tM34D5SiRXa8BmXzmmXRsozyz94d5Fqv8A9BMcIrPkiDD2M/RuUmtVXmZy5ZKRcweJojVFSyKtq
MXAF5I7ir1c++sonT19tgwL+Uswi+J9y49VVhFRRKtSsDVFzWEfTWDkZHfnzeMGJtDGAY/dy1A2r
KIJWsqJSS9o2TTMYsCPcEQ1eYWKRhJBRg3Ey0A+sPLkAJcdqCPFkWmkCEnY/XQ0B5nUGjdSuNbES
GET4CJorSSXs1UBPvHt5Bg5cBiiLAjBO6Ps6Ghfi3I5DT8SU5m23yaEbuL+3NKOyrVUctRO35SFi
9DnkG6+2QUYiKLv5JgaHduZ7VR6BhwkMnghSUrdkHCfWl6/1wfVhXgKMcX0HiWbqUGBNp0u7Aeux
1zQCvRaqbRwJfTxpWk/tq2dWu9rwHo2hO/YZ+zv+uyIMr6YeqJwQuUTr479D20I034sfJGrgs+2n
K2TgWOyzJKiRBgxMAEAYD78K25w/KMtmzOndN0O7ClyLCm/Q7JlRLspznlzHDOzuakWfWqMqdyBA
keNPOfqAMsaloGa1Ww0Ce43uaa65VtoirNjNrLStzmjOWzpAVsBynoTjyrtnva1WfocX9oRJi85N
dhMZJiQeEFEgn9vV5XYuCwci5e3UMey2SumvEbeBaGBtxfoYkSAX2KlXo/tjf9mvJYgNtdBih6hn
Bf0UtabvVRx3CB9vWXPjNWjLSnAfWCNKY0C9K8q+ZToQkRVvndD4pfx2+xLWrkljx19lH4f+ceB1
Zao5TnRsgnkDMavQFbWDQdmC/fH2fuwzQNxb7bORe/lyaL6MVyRXRNRCh0nYNONO9mOEDHQMcC1+
RPRL/ZA477HYY1FydP9Gv9bilZNS5SCJPMJ/up50MR/6avr0e0BUeT+k1oS4/zLVqsvCy6zGHvPz
UqVm++BceB9gEx1j8V8IpYRZy4UsH7aJT1mNjceprvaWlgf0HVdDdz5DFKZOdkcimwIhEZCqgYkc
Lrwuz89O6xJxR41sWYhaI+NBTxzjn9GEB1TRvWq8Y22rqffH2HbRVJ9JmNkdYJWiUEch7moxWlBJ
NOQyZwWuCt6ncPnJ8gy1ADqklQO2HWWasXtiTZpqZqnK0y1rMZ/b/Z99JHmxVDnr9rXLunsSVJ8v
AngSCYHhS7MJjV6PmajLeGkVOUzkohTFxSWLkdGHbhCmUsrCK9xwZFa97jYhxj5DAWgPeae0YALq
7lZfnybvKR45fn0Yj7hrLYFWfijxo41dxU3dcT4q0yysQ8/zzh8K2HoacexsJQXvWgrTGvdfsp/L
C69SHDGuav4CVat7BscIpNwgwFJJMZaG3vAos/HxVHSVFt/WKX/2Z6Sk6903QpKqK12rWXR1S+Io
Y1oPIJ74C/J9PP3JToFgCvcVUj2tl7YFamPhm/9ka6Buui7spp+VPE6RPkgU089ck9/g959W0qaB
p8MBywTZjC74wOH8eiuphcAOZ+PTV4dr/5XSuXEYT/TTmkhYKrGxV0a9oTGs6c/HndEqP7ccQjHY
c3LAFGdyVhMJ3/0FItmvWYaoY/xieqhV+vDS8AqwPUOPQ35/PaG7shVZlr/PjDCNq6GRI3Ddqzv+
bnutLTzPrbGRP6nQ/iuA0tT43AlbOtrfipkz17Qz2R0CqeCAkHqFBd85L8dpxRdlCH7tPQRdb/IG
Em6MZ1O+VW4sS+Z1gAl+kvkwKEwlLodLcI1WgEJ+k5h3UtlIf02fo++uoY5eZ5/Ae60vzSmz8BV6
E2CEp0256+4541IB3I2QeCG5o9SATMrCl7tUOKpiTrzLey+v8e1s7tsjrohUZ6JSRqSsJzkgV4pW
IHWFzsloE9mi1x+0o2kbIdfRt3CU77L2fOwL0SuMSU6fRl513zOuBvaVnI92DyYTLkkUhYLY/qWc
ZGbCUbwHN5U0Zk6ReAOwb6d3vtUSD+KKT3VpwlAam9xQePOfmMr9aGFgxKi2ZBAS/LUz4XnniOMj
X9uZS1+aZVHsLxWGbdlFJBX6CyvJOavZ8YQh0COK97jstvrcRU3ieQxmWw9c7fBCdM4NMyWHF2zd
c72IWm5o1TIJOs991zNpV6gl4vCrGJ5a4xGV8aneN31Afy7ZcNiQ2Fv+btQHa8qaPZ/Ib98YsPQW
dT38s4DsFkwqk2Gw3IPUOMedSZG37jYXMh6nb9ZbATMcdIwrZykQZu8NH017+qMDh2ESwyXgERYk
MhYajygShA47F1xOdgVfcM/X/DoQyd8KDJILy+5/eROkzbpt1D0/79CbIiF4wVrrXIBf8Eu/04Gr
gZL1TStwNeC0UypiFFnLxlLNh6S5GsEN8JGC5DGzi6sjyJI2RI11Pqsa9lnZicQ2RtYg+e3cXQcy
+AtaNaYKghKUJCAcSOyGX38tmMuqkUUttqB5ubEYNZuUmDjypb1M9nK54q6KVzAR5+f0MdLu6ONP
pvRX835D++L3bUxQ0nFhk+hIXbWEZVLwYbuMCaY7btqKp4N5VRBWSfatI4x1ng+1wUBitBBBO2ku
OO4ZB9k7DP/s64PNXj61Iq8hEZ4Ck54PHlpWWHeE6V25vhmbSjlN4wezb5tfpDHbzy3vrz/N9WXh
aDm8Q8qlaxEZjJP8+hHtmly7hctSpQ6O6Jmg1CaWe6VzYf0ZKLRQhBXUvPGfmL1uOwNfRv+E8ThG
GJ9lW8eeQyVb+QcD5XuFtScmxoUXH8GC+n5DWV3uYLz8EZ+UUOCnnnswvKqeJ9gytqoFTGspeTM9
zEtPnVsIfjYRNmQT82U5D2eHBJuQ5KMlRdObfwxSfnQIc8cvHi8YIElfuK0rL737ObDDKOlncSJN
Ik07JSI8yrreVvQdveoFFT63oe7AIaE31QFe9hfI/xwG+9t7W/QMi0f/dtQ3c9Lgu36/kvFIfeuy
bTCbEn/HlzGtHhJQnM4055xMG7M8fwM2nxAww/w/QK9lGLMa1NLODm4/8noLdKCMRjRZN7Cbs6jY
fcq6fSqiVkNc6uKcwAKCQeYZtdypMRHN04E+rt6N3DRiyw6I5tpYfDNn7lABHsKNxwuY9n20eGm4
MrcdSugupUY6yx/AisxXfmoUucJWMkawSEvy1cXo0w8a41p5uhnO1vcjOfH9MJuNKXgYv9Ugkmaq
SRassLeKQVgUS+8OjP5PGPSjAL/Dfr90R/lFs8yfsytULApemCYWmm6o7mr9LOxrFc0xyZxhEmkV
7zIBff9ppP7VVmrsLwNN08w9XSybceeH/hr692r3nYTkHrDE8g8bfnTFS/8yTuIlrfO/warN2CPP
rhJYH4a0fHS4mkcuSsbCBXahy2/UCgJ6tp9iTYDZ2srj6+lpMEBjPkvL9kLmp5jsVST/ktjW/x4i
fMT4YPHztUoBQq0+ppNSjSax0tVEB5nQ5K5qrLEtfJGj/p4hJ1wS5EIB3m+0+XnsgLZtBHmoNnry
arCrfWJ03O87zLjcR5uJmeuVj/Ts1XdVej2nc/9/Wj1xLGImKehMLrJypsh/fDCtz7Y1GBooIET6
yg+VakIGMVUSUkOOCY/wAZgF7aanGH2G4AZdDJptu5PkjP1tQ/R9/qF75pX7tquhRklQAIphEfrH
mNntqONVP/oVmhJYdVn8mWKxcTqFuQMpkvcu3Cv095K7sUFFrNy/DAykMr4gRCkwD3ebLXGcevK6
PMrLzfxLUYZKxJRInRLEADNXVzb1ktIuc06rccrDwJOYEiExOsxzwL7nRFG5bNMiaLhR74q5dr7z
LUt2VhFLqQ91gh/SZ/8cJViFE2dV3Byjd5vfzFhcaX1g1lErlKRPrG/V85jZm2vYOrVU6N3S+ERx
a4G2Dxx5ogPtqr1CBykVsm+eF/Uy2FU6DXQv/sCbiHmbtZOlJaz7uhmErYy7C7cd5gWyvOX8HTG7
/YiH/M8dSt8y2VQZjekWRGaqccR7BKNjKlgRzDLBVZFGzO5B7O2pblI5aBXbbUNCYHO+6cO36R8H
1jASpX004YmuYBNOAHDHdz4nCDkjpIpnVPA4vd3cDlwzpDhBg+y2E94FhwzczI9Kds158wvuVy3O
fsBr2VorvnLy1rZIQicgdFkCe/KxyRMGCBBmnHjUzqafvqNZf2EzIif1xdiOTD/whBcE7pm6muQx
aszzD8RRbSFTI4g6cJTf21huFrd3KhxiDnEWdSyQtEdE1ewRB02HhNcCnaNZ0axozqKlv2wKxYGa
/9UvJtJndc7DZWdSuBJD7RAMkSE3GGLsNF0PgovhnfrWxYsWAWHzuTZKZhJOp7eAvXrOrgSyvLP7
9/qGnKKc6awmACxFjG+kwLMXWyGmm2fngkuHL66CFP6b/ihvrG4B5UTrKlQTFuD60oLeLgR0ZUdC
sHjBeq/YbW4GFD5ADb+XNolBCYp8XsRj3Us/+hVaAFCMjaaFF2ILE0QZC4Vbo2poQe1RGhPKIP/4
EKkCtSkwfKDcWEkKJpP/AvcdSPWqDw2loXFj0g0KpT1uZs8V3m724w6XQSkwng//R9HVjV+yxhcJ
eLfaRIYSqsD9H/ZatgxoJRm+L3xXMc+IQc2b2LxbrtBwUEGPM3+vlcNCHpTWd+0B6Ut3HaQh9fw7
QbpquPRSaZWHVgRl+RvBjRzVb1d93T5GJnaZYEgyCG5zoROET7bnvJUO8xhk4Sbaw36+JcicKnrE
mFiQNda5tfLySAWzG+3ks4LXVZBEx4E5WbKfn1XeHrLG1FX7nrpTFwTkU/LY6gQqHC9DfqFV+ZJv
Eblssjh/w/ipmMlmfs8n00fWSKvPDjSEN1gNdWb/SGNp6XJs8lnqUV5FoJtoDLXR201uR+cQAUVG
Yv96bINQIRHJ3jO8Z6vsd8agNiO2kRpYwoYci518kcP0SvyYAC5AbBBlnZEIUmrNPk5z3wnvxzbm
aP+DryGzMmmPzRziOok/UQOCvLXXhCkUh22eREhDjXNgiSQltUwNl1SS5v4mqPY7KWBBV1oiye2t
cwz8BRa0o5SZgqTIpDjxHEnyj5Mdjz0va2RuvuOZOhI/Yq3x5szKRh58yBOp7pY1/M/BPlF1DHcE
6X5/L3Wl0J+EbIADH3HUlLtx7C9CPiT/QT/hWKCm+tta6lETn9QBUzrR51+lUHOO+7AkKC6e2uu5
wVfFtfs/Jj+gdULp/iHUdNCyPfR+wu17sZrxFcYXH6fruQF09OKjJP7rwDj9FI/yDRXh5ilas01J
3VfUi1DjpEA0Ra2VVPfXcEA/KxXUOQ+3+AyNorni/+KzFUmCS5+NRS/XqpZz05tz0K/jOV9C9P1h
snFeIHGE1yE35CjO6mZrGE0/6yn9jO7vhNiXpIkQk0ES2anO0JN+lgjBL6uxcxS1AgH4Z/MHhb1p
TGhD4EwWFZ9hk2hEecrdKpbfuHmimf4MKkyFN0BXPYaHIzYV/CCMYbA8qlgn2CvUVeej7+gBUVH8
G9qNo1mztQuWd63Cd0Ruh1BSWuZFu2QhLj/9weM73GXLcpteWvq6E5L9lVgdGdWAG2HRUY3V/z46
Uz5B+7C3BUKgZ6ocj4ejSqSKgXU2MCs8KXx4obE/EZ5ijQGkV7GPnHVFHiz50GhI6zIdNW20QyLZ
xwoJE4c+kJvoBAyIxVoswq337xv0wRLxOlgNCyvWkx4sFQRZFawKGES7HmnmBOuewdHBtyMV8KMW
HYksjlvLJNbBqdmIdKspUfdHDtpMDmEBRzi73J2Uk9gDHkCMlLk0Kghthm9sO5PsDtXTVhJQGNVr
4chedIkMrZqvDV+YaCAiKV/OeY9Ackgzn9JNqddCQxZjvbMORdhmQKi59yujfijFqEN+Q2Nv7x8A
A1vuk6NGD1q2ZhF5TqZNZGJth2ye89uvvjV0jIN6Sv2K15+dP1qlMMsPOgdbjWIO97GrCFced0zv
0JOiud+BMl16424GDptSvGYw/YleXDF96BKOIdlMNVk0xdulVp0u2LV13KY6xM3ftfH0eHVCjvx4
MB85bYFSCXmuBIhpIPgUXd90SW/xUrfu0tL+aM6Y+sNNHBVuxgBqYfncmi/5BrPR2TcNsmIgvAFW
0xuME/xYFkleUYFF1HKMvwFpJ0L0vhHcfvTla9wuRdQ0osjQ6duEaXNjyScrjXOMOFWQR4GF/R1T
V08fbrvAUm/KBjogNl9ePWAFtxub2cvdohOivPnYNFTmBJX0CmMfPaHhQdhJvZI6FIOmrmUbsgSC
/UdUADnyoNMqzXzM8yAwlqc99N9EbZg2GXbZ8BbiY7o9VogF0ZVBbyCeD+lmOLj3eRp8/VHvSNXt
UCzKBzF59gUPsGMr7nf5oiXHsAbj7Zf2omfHQJb/hpPNQeYXHJ2gLOashTpjg2xl/1fg8m9qqSZQ
FZfMW+xhASAV1Bex8/WG47t8rp+oA9CRJDDBJuQFAuTFWRk3aknrsry4kq6FeAwYrOWSp0Btz3MP
la3YeQHfm6wHCFyquVv/5uX0uo3BbgO8wTQQIlqQV/HgEKtvzybw9SlYkOKNmviyhkYuPeDd99Nu
xzuDy2xeVIMIMTNbz6O3gJ7inB44f6+iSDc+f8mkcajhSUcrfZ80hgKyuQrOqH3yxtSA4E7zUHzw
QfofeTcySUp6B2rx/vtaLvBCxLHik9G+U+ek9H3NEaCD8+wjF+pZgoUk9kdv64/O3kr/0Qb1AEtJ
2EPEgMfcoKhYsxewuO44MXAB3z0Tuq9YkjJK+IAscKMiBtZSVgSqTdR3nKa1PMqjCOt5MjQNOSfj
9f3IZtNrDeoUEqQLK66nbfKWKwzVqIxUr/dYrxP3PJ6f5KHTREEJRm9fs2IzwcZFzVOb5t/v9qt5
BYaeQIX917FCySQ84n79JnmWjYZVPiJBf62TkFiWiJptCXEN4GbcPZXOP+HBRLGf4xzGsSKhRsOF
lPQ9sC18/ZiY0hr40SGbkkjUnBAuYIj7sU1Bv0RSI1dDnGnvlwqpWuRfd2UKilDtWIr1Gx7WuF1N
MgvsiiIjvJBXTAymE6EjThLuf8Yg5483s1eFxlv508kryNvKb4Vin4bQiOaIRm6SRCxdLmNyJvZw
DCdYhRtZtElCvh2AeCSCqCQqmgZUSCd8cpx04isJUwqnn9WcoXmBjC0K+03y/ZPC4Tq1ilU2HXNT
vds5qY0JD/nxoz3VFfBLFiQJMGB9ES9VyDwTV5Ck+lSMbeMPOK4tjP5bzFiAzjnzrcUU8gpRpq6y
m45MrVv+AfD2XOqgb740Ij2Uf9GwHxVTbMpMf4c+lMwO8YGkPItKENsJrl5zDsFvNR3cSBVqviMx
tDQanRmWVZ0077m+Usvnvw/hWaflogRZM4TB2YOkCTQZfKhsJwPqB4XptbbCwBEiw9V5zFGFQofz
OvoxBbLCcOSh762hOVI5eey0jvzN8Se4Y/pN4GQfYFTO3EqtjcfPeEbVfGvWOS3MRfw3HYxc2nMj
ng3dv4WSYkWcU3kObwtZJ/mDTLRqY/NEZcw22cxohIireXL6KJ4+JuZmGKjSeSkoxSmkh8WDfBcs
ez+jdODvIdk7cSLzFJD7lBvKKRLiudoFN4HalJ0p0NzjXoswKU3+U8ek+n6Qd2ZVwvHEAYVcAAEw
X6AFg6mRQBvfdzubZGTdsl69JCMeK+OdAcVR5lt1yBBbF/pEa0m1cv4F5Eo2YAKA67O5aQBKeevT
AfGvH24BKFw7aldeE2ckq2NLu2a8NxvS5T6v39tg50NDJwhenU3Rjg2UL3Di17DPFN9nMoRIu3E4
FZxVzzlW3DmYqcnPx+DJf5FkJ7Y2sjLm+zkBrSeUjmtmtrGW5K/gADfMs8jvYKGpcuptESPoXhx5
tT+udPCv4wfrRnW6BG2Rmr6dmY3ecJaUuyJEoeoSIlo3ppf+d0Ync5ev6eRAWiH7vCqtT9NzM4Id
Rf57Cf3HV0KpIcdc8RE8b3FZC/xG5jb2YHC/NPCwpIKTuCqwKZPY2pSgkndppK0ZeZmsxqLJV4Eq
9FuHZw5OuYloIfdfbwHxPRPfc4S/HJguXClVzj9qzpXUYWxJ2MMg+ofSycPNDEbyzy0q7Gg6K0dA
h89RlQ8I7SpVo0U4N3kd/LvKSrURVc0qQq/v/BrIPPPsb2Kvtch+AjTyuM1TQWWY3V1W1JNc0CxG
gzjzMp3v90qrAuUgPJdElxi/jVLrvf3d1+Qljrq15dRb7cjKyf9/JRB4P/4xijSeNZ0mJ5NH0c+9
nQ+/mA/AkQPiRGhNsUvmtw0+9SiJHpOHtj7HkzomZpt/tP9Bcq/8Pz7gRdeKJE1DpM6/tOa3FsQm
ifEM19WJa5edep6NWMMuWfd0yAqaVEq+3aQ7mNx7l0gKj9R2R9dHMpGdThe3A7O67g+wZAUkk9LL
ekW+nnvUWJEXCNVfZDkoaZx+v3zIUgM166smFyjiqhc9NlUvhU1UNo8FZkvU88T4f4GdU/bsWVha
Ot2a0Z1cLOIvSrvavm9eoDYrc+jRLUn/xtFpPPGPyU0zj8uEDGyrPyS9/RwM+6BH7Y/c30VkorsN
1L8Sb1bYpQj6LDCO1X6d3Of5ThPASKdtnqRZ34nAh1TDWVTXzS1VQMN7pKUSREzNS2+l8DgRMlpm
Ld0Q6QNkv70hwtY1TwZ4WPQk+ePXi9lm9GnvbuYzEGTT24UT6YV72VSpo2MD70UgPaM54hwtqQbu
R8moIMKX2CYp0bf9OmPMPFdPccQKAKMbjzEfQlb/nbRkn7hkrjVkHyPIksD1KdnBSsiTfTcdDl1G
wouB5HHulLrTgz36O0Y9WzR1bANdBh3XeufJDkraYu5MU4nS7CVEvwaXb2FmkM8Lfr0Z1ojUR5zv
RaIDAsgN1Nyyrw4BJ72G5/B+7hcQMsnKH13vVB6BmmOph1tw3JlXUaNFqOsZ+o3pjrIRM0t4oMWj
82iqvhkF563Mdj9laIpgIx+uBKQCJ1hUZRQVtNxdhHw7IrD8vf5rAxX44n5ppVFdKjqoODmunnp6
DI1f/+Xz4A3jorQo0F47qTpte1UL7LHH+Kdgh8SYjPk7HES9Wnh9AwM9Gd7gDd20k7Me+hthgyp5
R5fO0H1lERV/iiUIe/f1cTr1+ufoF+05udOezk/ZisBw2AYU4X/MzWUw6MrVcZYJh5cfpPslYbAY
BG4YApOv2qBLjmoceGPeAIuJRs8mcGDu0IGSXjM0hkeZv3kCfzArPdi1+jDP/ZLJF7sV/I5olvQ1
MbUVrP0C+IU9Cjr8n2mpbsvVRR7T2GwxWbBtlmYiUknYwYyTjyAFgolmLNgp8VA4CL5Ju4kthq18
aruT0mRtGjJcfgKbOoSrlKZSRpdcvQtiAAfAEX2qJmbCAiEp6lvrLI6XWNjivkzqWtdeGBw0pqGo
boK1pqYvJ3A+HL+DpvIRAOOK8HpzHDLX+v5FHni+BXdJKJ2DhLVkhLa4TS2WnCntsFfhgDEoF4Mq
jIeOA46kL5h5rJ/raOBkWp35OZjPld0XjL8DhnRdm6Cqhu2gmpTGy8yTSeF/VESObhO/dyBWB1Qz
/nlvh3uUhCV9r8PmAGf0y459ivzvngfO8AhiUFOjZ95qyYax+wBJNlHto+WSqLpjQhC05MizhMzK
Hiv0XlfIC3rA4ewMy0XpUZwp8eqbZamIDDwVGbdtf7iv3tTdYTdx5Wp1e9CJO5MGcPxuD3yTUdLZ
mV9ab6KSe1owCBMIg3y5QTO4uvTc8ddcErdIoM8dU8ijyo8psBGe/lCZ5OVoykhzkGaCPVGNsqei
nTdSVl6ChJHsK2QcqpwP0ZNuU7/K425iCqnUPFIBK47Nj4UyYj67UCYHkxEzEUUfRHOgmUgym+Ys
AFtDq5JzRvWjnLPbZVFe6QkN1dflpmBw20ciZdk6DIwl81ovkw5yohNaGcBjuxne25o0u1Hu9eks
c5Kruu83gAe/Ac1f+l4aYXPZ/AjEXso+3cavqLdoSFKFYkRQHZII/UAWzv7EYpcPRBy9PokULOGA
O4d/9A3zGylu9lDKfhEqkvADhFO+pFjfYLFdY+5eKZZ29nWVgtaNfDncLLC0FCjMoEeVRNcVjRgs
BG6sOjynXcVZh7jGR1BFDazFNWYhly0DcMrd2QvrwngKfYOgPHr2yapw9DcNs+wMuX4qIAd/EYHx
R1aagNPPEqXROgJsIMSBFAt5/wf8LTInXxS9Am95Cv66zs6KfunxldAqT13es6pQAy6TenI9t257
H9dWmFkyjUZJB/Fkwo09Wr24tX0FDgn7P4FLOlRChngzdMVmxTRa2+Y+RuPVCIUWgGc1R7VMmVkG
s+16sGD1k3rf4GETGqjpWG/l3TzkDkwB5Ia4+aqDyBOf/4SR6iW28ziY/TmZYFUiOPU5ll+32rgZ
Tr+ork5gk3f44s8xjeTlz3x+g+mtr8Zof95lpnU/BvEh/V+GWfCcqudSSokUAy7vlPhLt/mTXl27
V8gDx9qoRFo5Jb38OlE3i3a3wmFmZLHq/QxZyxugHSwZH3268Sw+slUjKimmbbX/2I1rvYy2wHXJ
sTxaqY21jCfSdmmvwV1LuH1udMvKnS0JaELRYCqDcvBqCotQ4Z8RmhJMU+xK7MCsYbzqdRSYGU29
S4Ip2KeMPr7HrNp2e4YoU1fIFNslJosx43LJ/Vu1MIFzj49lCNYaBqYUQU+Vl2F1HYeJ650oBdnJ
9vs+xfkfgoRkgrURdsmovGJjojWvXquFQO0IFfsxeQz8UsmHW6i3VCPfii5luAAmXDMX1gukFETD
gCKA2PVjxiN76DnID90SfkV8PzUilzdVnUwr3IBSFUHV5F2dyEeLeukRWk1ceoN5lC9qI5ZboImU
yuG9w18ljgTOU6gL3ZiX00n9t5fvk87VJyScbXIJI2O15MQ/n3+3Uh7Opo4u3jpCTOotZy+eA5Vq
ogpTCDc6oPtDJ9yciIU+B0QiWipCy+Z/jNjwbK0KLszoAn1Tjt2uYx2GtRdoVCrJ1gzNyK5LXWwY
2YFmQ2ydLWfZcrC1Bk9m6zj8hYz4jBN9lTMpLN4jY1psumZSh3FO0VfTkdmzSq16SijA0OXYcaQw
MVw23m6s7f8Co5B0zdWVyf44lPUdH/WevUpPGSHItWAK3IABK8z7D0B0pPhhN2erNZVKw8DcVIbN
CzPuorQQr+bSE82AYLfe7YSeI7HMPbdhAU3ZxI+T6MlLfOCjewIHFNyqEjxgTATYs28Y/xozmwHj
rQJ4KstAHmTxzuFK9/+bNDBdzSUFELqPN3cnHbYGIQyFGrrj46N5zfXXK5C/kHAggWPxf3dABdjI
fZew9aiOxPejyJl8Ibh1dXb9ZFoNHWwTbEvETX4Ee4vp/oaYKm/E5K8BZvSjc0FwR5x5EJDHDZiN
7RYdtAmXj5JF+VSEYPwM530N4R48jK8nUPT089Mv6I7Uj69b0Gx7okoi9v/TObSPplhqsGxIJwaV
iiTbuNcd2g2yGx40ANmPQ/Q/ZPxtEQmmgN3agGrnclKHgCGuRm/NWT40uV0psRNQsEn+suDffmTK
aLZJkhdT/lHc0PomAz9gPsJSpv4TxkS5qB2oPywNan0uaoG+wnSZPGRV4UmYbkiAt4xfEEwKMxBE
U6roNHL7dHoCoDA4k1vvrbQIFy4QBTt/+da0JKoVE/gjI743li6n+80xATWl1+oY495H6Ss3XQP9
0o+xAQYxh9QkaPhEoXHiMSt68ho27iOmDEVRjbW8a6wO1ouV9MTgWJO/iNBVEviJSlZoa98qE34C
TtVoPOOaFbiEDjO+DP5P3Ag8jtoscpSanVDTA8jAehxlq0jQQ1p/P76jSf/wQzM4NlG/BWdNjcfC
jUVmYrXtU3M65c5vbCc+bWVMK5ysJMdjL6aRsZ2Ug52/ZX2ON9YxnlFYYPelIdXw/JNoufqUlX6S
S7yaa2hdlCLgU8pFMqGRrqAgnlomsZJ7aUo3bUP/cJdwgrZbctL66CtmHCFZc+wKk0hdfhHj8Dy2
tOTkJ+lBBEXWhgMOCEwsZiTLg/SlJdnOv6ZWlXh9FkO81PIFwrAvV+abxzhg95O/R2katYuQ+QqE
hQpxKFV/3YknA7Pk3gdYQd0VdHxSOn15Hr38y5AmBy3NjJjqDzJePQIebyOPyY4bxzqVpb5E+CRD
CfvfrUTu+jk921MsZ85kchX/aSMR4DeyccHQN8SJfH1cEIXSPkn3CZUPD/2MQbxeQ9dZwcf0NCji
ViWIT99OTDoQYZ6TNHvRFB0GcZtGE9/hboyQPv4ghC4A3on5esKlKKbChCDlcAnr1CRWBge1yNrO
dFMUZX0dB2KgHwD4NPW84ow5RRh+QGFvEjki+yt3j5Q2hHx/OllfnVUv5aAVnVTagCOXkDajWh9R
WCzaCp9nfV7V91mj6nb32Y+5cqoHwAuZjq8gGIWSRXdKgSnCENmP36MRLOA+QnSdsn5RRjWXua3w
PqCywyelyiqPIgSn9SjMVswbx9+uJxGNrzpVHUJa7zQ4lv6amc5OVXhleiDfLor/lm/E1rxQTMuP
It5D++7Ph+HnPVLIgradiySfN2qVwiihr+DGZ4ypaDXcwvFa2VeN2Fo6AqYrF7Q8w0bnZwMRbhm1
z5HutuROZSYfRjP6BYGVyuqdEafmyUZPbSLCiKwiALwRbOwcWZNpIkqFt11fXJxvsx2atTJep9YV
Cghzxnx9zEflvzB0IeER3a/xvO54TzoFYN9haX65R+K1reB3WsStmB3d164RKUu44wScc8LdQIEk
TnHwGaVQyDScZi95IrK8eDl/idrE7aDW9CU2cNgz7EQ9UP41svq+aRL3fMNYK5yB4Cycr0pysuhx
tBdDESlTC2ILoBAv3FDt6WfVz5hq4iPCf3ddF1CDsSODt2HejkCXSjvFiRs/vCSf9VXZy0gGVVXS
hDr3JXocETCi0uv0c9LEQSCdZeu8MlvqRX0w02BUcV9CB71y3BI7j/+NVhQfLWS96Ub3IRI21ng8
Guh5eocSYmgbRZC15GE6us2pqAOzbZzD0bHsAwoce0qi7h54r7WUUxp9Jl80280KId6+KoA/ydHz
HYeLRdaDFRSmt825MbmI2bGBdDyE8xWtzy8DN0fWEzpL9rtubeXrsU/dkgqDR5TGrftKFTYK8l6l
SW2z/vYQHEePr8U5aAZB9eWogGbfqj2RnHjlfPpV27voL2EmNquGmF5yvr5iQW6uZTVeo9Xfvc+9
HOZh5qTsBs3aVD1x7SJRAbh43GB7on15nJrcJ8bqeGHt0eyTPxdPoYJcp910S/AGHvEOMXsRdMOY
F9CG1g4R0lDxtjSQQnAh9jk8mIq2SUNa8rG78mHFxzzBvdf8v3+DWSebMtaSqsVFuqU6SgBQMaSZ
mDvgcPMg/sdPiTQR0fBOd7OqeUziRay6vWmNY60sprbdzlkM27E6K331wA1xjZNXlZiEgDurKhSJ
DjvPASW59L+TQGIqxcsbTLW2LcT8LH8hNffDy5pTYu7pgQG5VLHnD0v9ixrJX3MIYSPdDsJDIsov
jyRhVw/X3w7q4eVAKRZlG9ahTd2BS8Oyr+iH2eUQLbM+YyLLwNi3OwGHcsAeVFQkT66fGQizWIRz
7LWw5EIMUVVijrSy2bf/+Jgp8u1oPOuemakw4q/dPiCcS75dQTTL6PmoiF1bQemUz0ZBkScDTgBo
Y/95Mt7aGW1WmVbHK3i3+E98UhCNbZ3R5JJwGp6GAh8NHYQOU1JGoQSnAOEyulTxMHJ1kNrrBUM6
8Q80N9clpPt5q3OqJU/sTTQdL/xSz1eenzfiYhwakuyX0rjNApxI47h023sb+WeWQNDrvwZEIvFk
WFHjdt3LaYYE6CZrtPaokZbCv3JZWKLDIL1hdu3vyFLTNUT3uCiock+Bn9TaQ/VXgTRdlfYHukkd
tVx+f1NOGLpezR+i1DEFaWcZyk4qPd1Tax85tcbR/P9B/+bANNiHiubYARfjZ3JericbxM7ly2PU
+LRGScRX21nfDPuBI4koZIySC0EmQd8QhtgnnxB35/IAS1QxG+E0sMsy/8CM9SIZxqYhYWef6Tct
c4PDuHvytDUTHTSt6qopiLf81wXcQCgu4EUFcfgfINMdgoC7SL69kTrhe9PddY3o6zs1gLQ67Z3l
bzTiokZ5hP+tHh0pip6A+p5bI11HECvfTyAsfCqOW0J/oN18gtgALaU7D2JSeVoP50byey1ER1rU
HRAit8uAff92mZc0fLz0eyalcpKPpV0aR/Tuog5ximZZMenIaCKmWmtD/8OFgGO4zEC/eWOv2mpH
mMHMQJZPkyvNgt2/UleF5q/7/kZuE5pDBpiGeBITAP/9yZWabu2IJs2131dNjfs/Ry6qMwJf+y+K
QxDKD8WU0S3h1sBEP9/hd9pz3kflhiQEboYgRRtZQN4LFHdn+Ih6YwzN9nOM8McJwCkf0/koM/dR
AWF5cEx0Zushm0+iwVMbKECBgn6wE+Ev3Vc1OJPdfXaTo06EofWKsS3fUJfOCJ2rFPnTBe0nf6/K
sIl9gTUz2TbotQqK3n6ovDdTzEtVZbe/BSiOtqMDshRcQ3nEnKmV8V68/OD9virE7HjPmau+bep9
osou3HS8g6kGLjoSN6+cVMeqwfcDli6bbJ3xJj3LK3vVXy+H44mLVkivy4zqIPpQ8y5N0zJjf644
wfF1PACE/P0KLj/PwTMzYbSAdz2RSTCZYxoFrWoAZhq/grkFAOK7EsIOrS8m+P6XQvd2XcL0pw9X
Cf+asmGRK0kA9Ef6Dn5gQAH5B4PAZ9EnasINAVvjkdfy4VU7JeSHL289qq0PDttOKHeAhydkyn03
pkSrSinmniA2sz1v4kzJGpRxdRvBO8HdtZ4snFac6oZ1xjoCXNegc7rhppB9BR+nPajcNHE9WFys
+HLZtx4v93ZTF0QALUutg1KoZCZJmvSHA6ziY/9/TLQn53g/bJWLaKTxURdUWdQsMGyNpV7TTm0U
cGl7w/F9Q30mMRD5Z8sTMmfjSwlIlTIcUm2Okrjj7TQBRWRCBovdQnNvbiF3Masm2u6h4Jkq18Qw
WSz8ja2ifabcBFQpou1/DYlA/DAnxRSYc3D7BVZtkA86ZXKyQTqqItqN8obVAUsKy5Y8DJlaHSez
5qV4a/bV0G7Qbvx7RcIgxjhEf3Q4+brDlzUsYwEIugyJtyHs1ilTko4H1QGV6LR8JT8awVx+m3eW
zZvXHZWa/Km13UJ9zshw5cT/n7PY34Gc60g5ED5tgQb/zpconvyznxkBWjAPiLoymDzALuPChQyq
yUlOVY0J/vOSp2cg9hjociN49Ho5DXTD//Ylz9xSi5OYogGGvu+InTda3CCp1Hsrnv1z9FjVS71X
RMAXg89V0cdhDOiop2um1a1gCzCA3tdeeDAc77UegI1n+gTsF4m9HaJgO7hOOaozkCAxHureyRw2
ZMSY5LvUgfQ+KLBn8hoi61w2wQ7gZrvYnSAKuBapBcdVRHL0RClyqlhRfwI2DykuL3ezu+EAzjnM
wPs/Y4Q6yGZRTIOFOrvAnn5A+S0koZ0ugsqqaZgdwQL7l8RtSkbHrAx2tCQA5LdBDu5x1UXaFXXj
YFchyABL38b2tnCN64knumxkmL0zt/ZxOryfFeWIBv/s6oEdQkg2SCwxLTx/677IqzIZ6xal2Ihm
LtNMaA8JkDGX46XEeu1y/ZiqnMiBnjUW+aMa6RCvbJ92O2eoSTJpOWo8uHlzfCIob7jonZPABI/u
AnY3YHoRrw3y1dlwmDNVglzXs0kp9UZTxsfUxlK3Z2x76SsY4rZwPbaQR0GhlrC8CMWVbmiTXdXE
mL43Bj14X1UecIx+hrqoCf4cZB8w0QgSauag3jjfj7MeBRKCiUGPtklAOgDMa+SuEtoKJM4SfKvS
22fDpvA/c/UuQsGlRkf1PM36+FfC1dyWJ6AHqqrlxD1WJthaW2VplEgDkoNyUEJaktA/8vKWq4RZ
IJXoTGK/fPin447eATTRbkZMj76tNT35plMNvtQw7nj8bYP2B50+eFlwxti3raVxYpS47K3L7Cze
ElBUTonMbtRUxUpTKtmDV/kytkKY1xyDnL/wYPZzjGdYpL62m+XAC8IYnAfKS78Q9xY9X45IFWwQ
txIMAyINPCB2htsIOFfpB/sfr9Bj++v5qP8VnGwxZ71e6ebQqqzIppr5tEpbHSHR9ytaP40pZkNB
4wrYzfdZ/rnw/HlhJ9I8rLBpKq38nd7RQTDR3UR7phnOdoaTXRE0fAKo2xIfZmUS1I8LMB2neI0y
QC8RPekvq/tKvWeciPztRGBQl1AvXxL/Pu843p3g9fpEIU4tYBnCJo7Mf+Uid+pOA8xho/LloCyD
jYeoV0yCj2oXXK3Ntwfa24aFAK+a/eY4V+E6bcGFE7+nuwm2pJiBf/PpBcdaU5x60nuILc1X7u7R
MXn7YZtTYSdQ1qRz8FPyIn0TOwCvoWHkwFjKeJQgTLsfbpN2XfzZj+M/TAIgDBgrpOJfY+sNv1sh
6uVLfHcAD7YckwCGtTqnY0ByQtu+rN8ZdfOxG0WrrW4fVaThWxLpe4ZKVUBHKzepZGbsDCMqaQF0
BTzeIPqgI0WM43yTDmzvJGwJGiX/UQJETowuHtulERmINmQEQkmNFBXMj+KR9+KKparssaxwCGqG
6VJh9+qSzB2eceEY/C2VEJgNdb58SBDL/vrjvPyvYbpSuHfJEYNoC1QsFwgFrsQWNzFbKB6wDJwM
F7kvZXKshR+LqERDgLpXM5mVNnBCSqhUsVZ0dF4bGPRpirfYKUa/F6pNDsqqfiSIFJ/ejpKpPIe6
a+DhKI5kMtkbpnKWrFJA1VLWoglQomh8T6Trv3/ubBmX+vv+o/5q5137ON4RafZ4daZCD2/Kq84s
pCsvMuqLd9goUd8AQk3ZTUy8LG23WjWqxDmqyCVkEEspZMFo3uSgnUucU1LXXRf499/b2cGrdIb4
AzuBx/ZkR7jIT/BQddw9YH7Apc+LvlPXdqz7fhBhSE0hJgiKWOAkYD4g2nbtuam5pMbefOzg26+V
VvsfYBGTZfz5Jvu6iqZZGU/JrskZJc8YVofAXDjfITm5ge1Gf4mTf+63yYGmDbqr5mKTzIgQVT5F
rxhh5MgYriqGwFzMwW65Oc996lXsnq6DeQ3GMxPHlMKpoonuna6uLmvtAoW96H45EoQ+KgHSeoNq
D3ZJTLGHXmJLJlB2tF8zntj71LKYliUObKhr4PUv7re6rEzthKyx5hfzV/VW7xrKdWOAVbA1LW1N
ngnsivSKFCvRH095wVtD1K529Nh6dm+w31o5S5WRytbM8ZUa3eZ/7wl1VBnIt2j92316xW0weHfG
w05g9PFUr7Cy8GOwb0a86PT7kzZwHtk0hWJjHJBd7dE3CE3D88JQzJ8ZbgTYajk9M2yvCTBn9sUH
ftxn5YZadOYg6qhuKzUC3zSgaAOO5BtSjsJeOGMrlSrKi0RSXcQhMl0IaI6/iervOGuwYgbCd838
gBVL1zWlyFHM1PpBMH2IiYdbzEkzp+5Qmb9iJtocsFEUB5wgkwfjs8M3A66iwiwP0l53dujOcYzY
WKw7ikZYEZkD3uVNKyMIRLPhN9XbL3/ZQPG+l3tIxvBsJFqD1fyVa3VUKYUKugxpfRdtylU5p8b1
6WNghQusojUz0g0LVlHg+EvguCicCXScGqj7+bfxucTehDfdgO8LOQsTiDGi0tGiUDn2n39VTOmW
7dLWFzI9FrblqBrTCJI2y6GjVdOSY6h4RlJxXWXGF22yChYZb8brF4LG5gulX4ddl2vhgqU3I5Ft
onY4uMMej1dY1WMKbf4GdfTXHMqq8rWrT5MH9s4cXahldy+dMW1EbkneP+NOCI1xP9hSDoF8Fc+a
SriHo8cCQJjDpzihr07dGU6CkkAh9JGbG5o3o9XfFAbViVilocrVtJotbQ8M+410ITtcgQWiTk8l
H8JQPKyfzHNOlyPkdc7LAW6N8oqmVPLb5+S5ZvfxzMXpyN4g48g3OZcFvtKxbkKwrVoCBuNKdS1m
oHOPL9Ly9KwN71DK3lgehV/QON3YtKxQxUX8yFq7jHKMqVZyYy0PLHPrjsT36qF8kyLfk+Ucm7rD
iMeJhweKLSj0FqOWZdtT/kb96X5s+R9FhsACYMVbg/A9fqmHwmCFSd0BzB/VFkjcqO/j/+qvvXRM
Tfud+gyovP2UduMN0gdn0SMWH4dBQw+jIu3MqDQMHwzWDKu5Y7X7HwTboqtldIfWXTfl96omgfo7
g8LIOC/Doqf892EF3YGF2YfPb5DEavo4jXKKpA3RyCm72ft+9QYPiXRb9260Cb3LLMCFuVKtQGyi
jnDOHRqpCrfl+UsuTVQmwrsN5UU12wCBe9I0iiHIO36or66m9YU18eEDylVAP+zwIHyeDUCeMAna
J8/6h5SVGQJGA4fPLwJvQY8jybgq7bUkepQNy6M2JXY8ZNHO/dsUBISDflnUfvJkIEa7HodwSOnQ
+8hEHOPqyB5w2CRnWHVHrLMeOYbCPApC/9R1/XLRIU3IHmEpr0IeT5p2W4QigWdoU2A4Lg85zRDe
/9mCHxeAjcS5pWObF8CtYksIzcor/naOKq4sPHWvP4MOd9xbQL3m+cwbC8MEWGxCZ0u7aP9EFy54
QrZKSWljZ4vebkpBVUSQXmT+hBERCixZLMx570XEgTMl2FPpJFpWZejqhuYGno07xTrMdnT5whSP
xoE9bBvYHM9/zyBpQSLFm0+wapKQfoP85+Ry7DMFkqsRO6blWx72FCZqbLDHetquWpWYcIvXQOwC
CCuWN0ofLsL6Y6wtVP4l2SdqyzVq9iqGPBkpxqm47iGJCh0ht9eeo/Asu2Alk7WfRISnxBCyozOo
udmlYsIINef3wMkFpqUUtOvSrannUUCtU3g4BuPfFqLWXOJKQLx3/WS76/l6LHFd1Va1KeF12fNq
+jOfVaCmHM4LvveDoMEFsnHwyzCrOB7oXMt1IplmaVwTv5+H9sQ37Zxp53rA49p/PsLwwOalQvRC
zbq6pDM+odQOojI1QiUgOzKB8gD9Vgj+lre8HrufMTOeWAOLQl/EaJDqrhRmtZ55A4oI9toafH5B
VBbVvcJUN5QE4MSfekWXKCvZXMIF+zi9ePkys5ptejsvDy1Qfp4XfKWXJheGEj/aypy0SYiOZnex
5hs1Pek0GLKTLo5M7PvHu1BViqXmTIRbmYzCjCuX8pRQquQCKzHWKlmdDpMzGnU9xbbnOeRSwVeJ
wgdrjnWRwmzVuV4DenPlRwufhzQ9BGC7XfDkZV6OBxauszOSzv475Fd+Jh5n+puSEWgcBMxDco4V
CxvsvYv/04YCkiYSf8PVJX4BM+gQwB9yjcq9+AMJhegoaDyTf5vud79d3nnZ6EmNq6+WRYV+qhKj
dN+/ySZsCMLJt5O/dh58oPXOnjNmPvFojYzUINijU5RscFN6s1tHdEIcigcXF7/xUAV201saee4/
A08s/5uEcm1KcWMzYQetqwSHbnSR/uLpEea5bbn74dBbNpoEJWeeWKmfVFWJchyaLtqDuiONUbBp
uG4sFvI95oLdmaOikynomfCmy3DS/SmcG3TttSvgkRnhHuMH9ci/w1a4QTiOBf/BGdLQeESGCjxT
RWabvSQ6oYWW9lkPO3/QVZWU7jticmSDCrQZk5bXPbM4hYcsZTxnJHcexOF0GlojLJCaYCvcKaav
e/5CeRocfbZnzGdbIK63OGJgUQ/1S5VmoxYRwiT6xfaeXFMhMX+X0iWoeaMa3zOF/eDkwA/xwYgP
wMXA7A7uYxqjHrDN118RVddWcQhp0JY5xaM4G5yHE0LjADB4htqppGw1T9IozZc7WmvuyESpKbfu
Fvdaz+HzGmb9kR6f7I/I0BLOWhv3kmVD9AFB4KSBP3cYIUuxfsJgk83lwpFmFdYNL6E13ZzZ0Z89
a3RI/M1G2669u+c7Td0g8FgBvp6Hz5imQAbsuANuqL+8Jt1/947gd7V+QLQy5tZOzI8z2gAl1fKq
nq1pyr3phM781V8SsZf6I9R2YLWD7njdc0stfspiLWcF+MNieqMrqJYGhXYHuE0t45bxZ0bVVYkA
lTJrBc2I+7VzCy7CU8rIZD5uFfYXKUmMEqfbt2+iCGzu5nL/YhO3iXi8uBiU1FkZl/o++rEax3MG
gYpbqPj11GdKvCYOZC4tjcWn33fQpQs5OVwJTxE9e7z777h5O0z9s3zWJumbdmeajueXLLRuOgeg
CnlqTmUJ0WnjGmdYeWzYSpWHvMxsRhpiO3M982AokVuVEqPDyDwLvEr6qbYGH1bLCuZeLfAn6VR0
z705RRdAO3PMxsr3LsRQhDGK6Kzj8sJsR+KOLtZyijTyXa80HW8p5RlZWnYwt7us9/HxqKnJDVeE
BlgkvtlUN3Jyyxb30CPkU3hI+lwIfaXl11Z1HIOn5ZpDRF0NxPpumlDTesnZsuRwcmR2EaNQrPdK
DY90bbT97VC1zCuOh9eJn2djwr6lucVqtOCguzMggkRsq+P7a7MUS4VrOea/WXXSFmUOC1bpiugs
8+cFYqksq0uV1hB1TKzVOxozCB8HWI4stJHy9/yL3STVBb0ZFoXAgp7jYHtOck9bNQO/c2Jlu7lh
nYE4nRfap8h/e+1fiJxXjuo/yMJtLDHb0TCC0m+ahAOOYw2QynL2MVl+RhNgEIIveEQQdxMQbSEM
gs3EZWvzGfmzcdLdqqr+i58nDjeKEWH4MVkUz81K8bUDml2otovyzVxNXf0KTPKRsdES4gPhWcim
EXA1R5s0NybZauj35i0Si1p6sCBOQm4P0MNjQZAGvWMRerg1Rkmfnww05a8MdQZugjJgu3Sr2WPh
iGUkc7Mgp06N07CjOLZTXqbB25Vawpt5pXKIDHB4jbYa0gvlUnChNOEtSpgapGeNczpZ5JXgUlE6
XTwTZQIkngkTJPo6O2g++EETFCgdk95KpcrTyKXKp0tn/orX5GaxFhNgK6YXxhN7qX1C6hYfD89v
vqr1B4EAUiNjUW15Aj1QQxhS0tOEYLDxwScrN29yhoVucu00kQZF5XjVnSmQxjF1igEmoGc1pBad
6zFEkFjpU9LJKJm24rtuepEitdby82qV7zYqR3VpOY9Y5EzRIeXImITeumsLHmMsgwfTco720XGB
C3IapPV3B5QSiV7X/Ow+yXzdkkSUYZBx4LjcHspX4qOYpPncNEOBp2nZk6K0nCNsutIf6ibzhaCx
mvnwKiylGgn4SZoAygznQTqq14lgZR8pOVIkSP7KL0Ktcy53Snt3oX9lasAQIliKNIreX3M/WClj
A+YCGdPxG4LmL3492vF/b3YIzO3aKeyMrz38G6vBzdUhFeaXL8e6B0lmMjH0SFwUpBXMWvDxqCwd
GAfTzZu8PN6sGQLg6ZZfcTWgW1jbMpUEvqwN4z+LsSBw5+ga7CKiz8KN6nMTCN6wHOLzxlx7QaBO
oQkKb7K/qPu9whI3nJE7zXl65BWINEtRLddLu5IfaE4ndRFjUlRvvmmyLm/Tw9o/mnIk1ITG8YwB
OdW2BzUF8lTfnXYHkWVH5ggKHmbILwShXkq4pkHiP+T8c5Y6XOL+/p2p36f4UHGjgE7/3HaPAWx/
Czr7zZGE54uj4pJeSXDqDOTY9AcngsETcZeGFSq6TY/hbS7HD4Lk33pwEyw0/JcgQrWrCKItBpiy
43i3u0U9EbRrKmzzVPc4JTEHDyvy40+gBALY2YKBjsCjN02h+OmdoHoea+8S0CJHt2ICPETOHmdX
5xC5HGbfVw4gN9frYKn4vfQtcTlzzNtx5gmovH/Xobuwy4t8SBYV3Ef7pAcnOXxWMP3lzqkONha7
19xnOKlWLdMaY6JyWUnp91Uio9BNYrZeeotHmIlmNseUEJpzWsFOl42bEUxW8oLBMsTHlsbrglZa
k4jVj++HWsvgUP3KQ1YXaT0gUXotOsgSlMhdsYH5CInnlAWWrLFy2kHf+AYP+E4hqPpuS2ivXJBg
G1mcwycui92kTzxjyYNUhbGTOjFXBLNVehs1hdyjs1mdxw8OjA7vUNtDUVPepD+64GmeOq0/gg5g
/oPPPkBxZop0exo5kJz/83QRGydeMu9R6XWdnzfyg9LwMeMNurZEOvN2HYfUdWNbQ5IaGKHCafUK
G3Uy6/DTWATb1TH/5JoLErHW9cyxjJPuTmztgCY1z/h5alEqsWQ+Mc7qffBfElK6W9Qr7UOslrrV
am2eOSbpwOOk/+6mr9p3hNwcqOqiEDcVbZoOzHIa3ItRwxmnaGCwYJ37+xqLdSbTC/I3pBMhRD+c
2zgJwRc78gDumFj2xRSayNqDzrI7uHuGuQGCXYTSFqEja/iOelQE4+i8TdgDo/ZlXx/WIZtgUd3U
4/cSTFeNAlW2wksXEowRecSb1pPqT0Yut1zhf4SYGoRCV2W1if58EwSxbeodFm7VB+rdftY/b6hg
s+SfkJyk5sbCdwjUmkV4idraoppdfq3WjaQapM4bnH+0HQmXBZI1GtR78YbJmTIXbXBTl0bgUGuC
5vzjrseOtfzn3UL9qI02Iy4U73Jwb9OeuWvDdmgj6OEjyWyPwkb7v5pqBCRmywalsz/BlW8aiG4q
p+yCToVC1hY0wctiUTW6pxFGXdmeyFWEFuDQU6L0k/n1RBratpzZAavYxtPRjRD0KbqZnzf5yWQO
+1sA68+R3roDvgcUME09JAKtahYvPvKs9ayk80CBm5+OmcoHLnBGE1qTQCnoXmdNSI/KgN4n0nc8
gpaGeaGSXArTOjXWXX6pMTb5inls83RBGgJ4tM0MAmVnNPHc27CZn8BFfhnWnfe87CrbHhYPO1nl
sODulrnBIPRB1cKfMB06y7D72nPiDqFCw2+UtmiGsVWmpcNI0rw4ffrB6gN9oMIKuyC+Z9HH7CIM
ZCXuo6fN6AECx9BfD2yB+IZUUNtYOiuJRluhBJLSB2cf9K/p2/BJi0596y//+97ADdVOCMK7HfYx
uLXGEdYc703vUu9VrbMPmq0iM2zriApQeEl1XEy+f7jbfVz4TevRvDf8pJP+cXn0aj2o943VKiTv
Zu3Ut0+9sxxIRef6ySN8rJPXBgQrAIwN2vp3umsW6ENXc7JQl8DvqckLzOxDf1Fb9JPAh4ZhcpHi
YvEqYFSac70fFkifJ7M8CnXYWrB3kY+iNTCQhRpsTjDLGcDrJqEJ/y4mMlFMKRXrzSM1Z0QBus44
xZ1Z9NXVVPr7AgrDaEh7nfCB+uy5BIKVDAHPGmx7BFUjDOZTGXxyb4aoxddxoKIX/pkGdrt20wZw
lEBQfaP+vU0trCwkzd/3CoZG5wh1QRB9sUq8T9g676G1X1waG1KwAYF/qZAd/Pfj+fVNUvxrIBVc
wbkcZOuTUW07puLuijQpSH5K+YplVeN2qk3MYzEbLDCLezKVIKEGSfl4DJjNnwRIGL4Msy7TmaWo
KDiD8/B3Z10lWo+1mJl8dExCXeQQhOxkY8ZuuyDomN5waVNJqSG2Gz5pH2tODmy/EP4gsBhWAwIJ
/chV6mNt7CXOBl7c6GFqyvIPq5inSYxiAMsqnQp5N4/PBtPpkUTLxRi6EOz4EfIQT7Sf2cmT4jlo
D1gEbWiOlA6q2L8ikOmFJulNEtlYuJk8yGIyMZI/Nwy9d7E7g0ImpXJDsO7HsB+Rt9v1apra/kDf
Txe7L754Qkiu9AKQhPAyLAp9NUWYq24VCbIvhdkTKuNcBqL0HEho78Uwqwd9lVbGh2ltj1i5K1fI
5wN8/MVVsdeTDxVn+o0tGy0EVW8nHvZjkX/A+dY+fUqdkVAT+sFhuv1uEYm5puuUnA9mX6zi9/cV
mbNgf3enrDKon8js/mZA2TVyrhg3C2MqRsl2AfRTjUAbuk6zWl6lWwzcmDtbw3odfzvqmSrq7nGl
3dHE5s5rVEiLMkSvL98XogSKEy2Qi4f0VhAfknaUhBFv7IG3/tF36JKKVEjP4EOt5Lp4MTWdV821
RXKjZAMgCH/YEtL7Krfm3V33Cqa8gUPemkSqYQTitP1epyVhbWCCVp2gM3fg1VEMVRvqJXbtoJXb
/sTFVYG17RL+SaNNjFugVViReVlfhun0UbhEd58cw6LWQZqQ4mIDd1enQmPZrGbMpbxRqvkJUw88
r9AOIioPyBmlqQCfKPttAstC6awkXxjxURI9warMmVeYdDnkDCmTjJtt/dD+7Fol43I1e2t1MHgT
8r2e880e1EGHKxMEsfPkQT7TD+MHsrFLJrGVv4FlA09hfyH574Vs/8rMUS/XXatjpy5aPV0Brsfc
yVkvFwusT42QB+ifIi/wX5t5jFmXmI6JK1/bcjXiqkoPxZSYDElqJGupeyg8lTJQVc65xa1NcWng
l8a2o3qrwlePxWTWpwluhMRQl4wbqorseOwIB89AysUZoYzBfD4rJFa31epSEdUVOpJ7Ch6+nQgd
C2+Yc3Keys0AvAXNIkNpNzD5qgGzUHK0mJVhB1KWapoW4RyhJpYZJdGABpR9mMgP6p4TDs6LfLhY
HA0M9TUccyI/kMtTvnrQ/DYLHKMLbudlwB7eNeK2q2HeqJBpB5HiNYOtitL4D6fFcnkKOZfQwKSs
EY8xKHSWeUGJc6k/84/0X/EHu+8sRlPHJem2FQ0FpPdCrieiCMhIWdqPQ95iEMEoH4DaLfx982hf
OAIQI+oE4PFn9bu/B7/6a+VZYG+67HWHSBXMlDaDYq47cOkazMWuhlOL2Li1BpT+78VPbRnSbDma
lpo3ZpJ3JNsM28v3lZJxyqV3t9MEOVKCIyM5oCJGT3yZTxivdI3OTo/jsBY9XIyY4RI8KpPZAwKo
3Ldd0YOYg2Koft4cF3oUbswDcNhjq3oPVDFrHuirsbMWVO9VDU29cee8V0YL3wkTS13XM92aegUJ
19kUrB3Kx96nnVpr2zzY1N0lr5RACpnBLF2bPkYy3LBk46No7S71iV43L41dYNGrqWVQO3XMP9r2
bXdETu5h1zfxZa+1TtdfHvIgz4hiyfok42g0b+3ux+4kqJYdk3PIPN/O6ddVH3ZSmTSrFhpOMXUc
y1n16nPQcksl4Q5wQKE++wUBTfnmh6Y1XMCwmleOhlqdKsL2bLaEuhiWWykgIebfIRZgu01pmaZm
ubuK2KqfT0i3kM1SjM9piG+MWbbEhTy3TiOkQGb6FOnxQO9NOJsH4ef4PXbNV5hGjoGi8IE3NIUH
WIWfo6OZCYXsg2pJYUrgvqhA2q4NgD6PtxUMp0LD/qZtijYeb07mmGSqmR2d+ybQGFQd4zWqU2HE
cdyVIrySkcC9HQoSNyB8Vme6KKUTOmBNAD18sF3Pkkwz+teD1deImSy20FTO05yjSwJthYgoizya
T9D4aLI+SitUBf7J1zWBqXYNJWVMiVxrwEUmdpNsvwQODh2r6Bx3J0emDxC8MlTH5HqpgEt2Knxe
yBqMzz1TUBo0bOKgcLqhAnl64OeZPy8dl2y+GEVbdhWreShbFXAc977+b7zYBF5YVzhcDo02cbCY
pA14NKToM8sqRxMZ74CW9nUumaZblbzBdcv0YpoqGPo5UPBQL9F0xJjELwHcNJYsuCCBArho+lIB
pnSnEZHyULbH+ycDPGTvLRHU7WSI88JT362DfEN0eZLeK+4r13TfV5Y3xDcaAf870QhUHHcK0dNZ
Z11FXTSKwA7mpgZw1DcBInJiSyx2sfIyVvkrshBdUxXXanaOW8mBkcJx0EGeQf7VmJD1rB9szuNo
Lr3ZwHseb7k+2sOILQ82POSJYw6rTC7gRt4CguccWqTWIHZIvagcwrJyZmwB+mtl4hZ5BeSSl8zM
MwHAsJW7iwvaMMDy9mNl2ZtOSWrPD5gM93/I6UHJOj1js4oylBORDcud2MCTIEqLkpIAxm5t/A1I
LqFG0SvV1CNKX39fjSiwpLkALlURDnCZ0zz3k/143oMQKyGl1nUvo58JE5C5pHbdD6R87qB509ly
WNUlwyr49qalYwZWGI7HCgOTeEtxR3smkuuwvnAskAK5FRBoJbuV1YNZ5kVP9bUSWE46uA8aZBR2
z+AkpihAEu2adiA3MVnO1AJchmOwx1ltLwYlsahsBBbNuDU5FyqMM5Ic+8hOPvIra2FTTVrkQaWS
uq4MS6xL5x3wPyB4pN9abd5cb4PphIWz0M0SrDXxlMZx0zLs2EjypIJAYyh6s0ZXdSOTT8hrebts
0EOMy4yQLdCf0ST+TPhrbn5CllNy380uVYb/C1VL/ycb4CNg/loDzoq8dI1fzoqVOlK2ttPPmqS3
mh9L1JKKNHA2ES36V4UJWVPV6sQmEBk9lp3Y5hUk7ASuWGG5ald3Ss284ny8IXGVi+uv8gB07wLh
jXhcwRKOolCL6d1SuA3hRSlbYgazP/4pfPhmAW7f4ER2fn+ZzZG+fH5ZeIqZrfkcFRUPj34nfWl+
QY1TkKlZ1EOeKoOyAIjPZ0ne99btmYcY3Tc7HbnQMaJ9J68G5RICxfZIQA+95V1hPipKWxSn8O5A
5JZNZCSTWaffyMjoNVzgXeRxCOxERgYT+8+8EcvSVl78cHwL29jJldcDwoJQ3wdjEvZvKgQmf7M/
5zK1KZVDxP4xVpG5xM6zGXKMNRxK0AXujdXBOSAQcJO+Tq8GQOWThJzCflvUulD7NxvCl64uDyWc
/SugRsoEAgUQ16RyZr5sOwtn1ZQaPmqgVQwpy8j/EJoN61SdfhTTERXE03o1iXrDP8BUl7AlNc2a
g+34PCeKZdhpeyOdwH8fJGvggmQt+7gaN3Fx+ItAacFr9mkXqA+sYNbGBUYzLHLLZn1vFTpXmDof
7Z7H4ZEbFRUWvlEsm5F1PIVqntPDBzfTW5EHwNwqc4lQpCCqd1s/6grrak/M3jM2EzrJ3vEQu0kF
zKuskIEf97gnGA9tvQIwx0o/oy9emA3YDPm1J4P15YW1iq4Cjk8in604SGB8jm3d0cnNrFC1x8yK
0Fd1h9+R2vnAUAS2mAmaq2LZQehNbbXz/Kd3yBaN1VUyj3wOTdVFRXE11vJ9FnaDfOLXg339wbO/
MDwsa/dZVFCcXe5/ehYItQ3Q1sEr31u5E3hur6PMLe9FYVDsGYuWnXlOAkDu7AUmn2JU5c0ntkgk
PhZtNvDJIz8q6sdVibRZGmf5GhIcLnzibjjyfDvWYaCNIO5gVgsBn6XD71pdTTLt0d2HnZNBH8YB
jzwiyKk6Vpmprg4YBqXfZWUmbTD3tIPsB42/JdYWAIN+FeOCmjnZoD1RHbACcKIB6D++TSnS+2Vn
bk0TB19dytiVQJPO9126lIjYxvNLiWhEGXwzYnuaoO50alt0YX5cgomOe2EamZmiSiXhYJv8rFFC
aO7vwWdtpfb0kOfeQ7SToHyagJ72s3HhGOtFvX/JrU6JNy3ggWb0fEqwwX3+Hk9WHsaX2IbDT53w
gPfgSjCXGO8JjmpoBd6O9s8v9wnZ/wsCStuNZyzLrC08dSzwv+1ijkLXjyGV4BwkztwrVHr7cNMt
tgNAtUkI2rrzqCYCokwDMkdlKaKqz5jJGwjuJH9fc6mZJdEtGVOIKJQQf9umSC6wTiSm9O0jkd6n
y+oiL47YLNK+1YvHAFzfZLW/Vqy2vriCj7jNT7/5NDBZ9v+s/cVwtCaCT+gQu3VMdbzb5emo76/R
z1e5PXNdbuYdgFs1lANnljeHt9O6gDplnFYQd/FV/r//4IeGGJrCCo5S/ggGv2iNlsdebjTG68LX
KXtu95tIT7JqG2JQcXs5Ebha1N/yEI3V7KB6KpY3FLG0IiakV/0hFAjKl6TLcg9r1PV+HMAw718l
vFA0FweZxFmdTnOKt/PqakgKylxYkdnq8ljl1Az8Ha5UqmYPp0BJbAfFgYLwOD1FycKApvc5tZj9
aWeWW03ltzXmz9Y0TJP7NclfE592bmesx7V8P4FEAJ5IVg6C8blNn/pJL/yHSR6EkL90LlwQkWzA
kf+fcD8COPkOWlA/XG16w246LgUG7HJBle5RSVrg51mk4uXm4XL0LGkLBcJxVK7LxBXJ5OAKY4gP
duIbuj3XG4A98CAtKq1pv5QvRnG3mMN6mIH7VRpQy4xoCzzd4ypUHzZH+1P7sQ9XWi+8H0sAf/rp
wRAtv5mvS0OOPIoppW6B6BwADhhV22JNiechxh7HHp3oW3SWOzsliXLlMDd7F07sdq8iKmFx1ZmU
etIUcPS4ikvdxF1d7Tcch7G1obxHO5q0tJXJAnjAIgQe8pBuutkfWo/VrCsxs73sV8EkpX70TzwC
KFblY4RWvKhSSmtjnE5YQh3hmyHTJaE0BMGBK2mcHYjzdJzq5sidnVNyVLy4u76UsSqgPF1MjebL
ZSQ50Agk+PqKQY58VBO8YbhQzOO0N1OcO1U7ItN0rB+D4Gj/h2eg1kyC4jUR1Lz3ofix9tc1MCkp
hQOU4BfUFvOHgZTsKRHVR2D2Im9X6m9OtZgy29dyrUkFmtcYO5HctjSzU2UAnH4sSXyi9PMtctNF
4fQbBDNRhJdHzSNUTSbJWiSbovmLz40tNKPvOLFtay2vCsb12NnLt/nb1pVOsa+dKne6pm0UhE5i
BIe9+sCz0jipkxhDAWy+LAjcgRB4mGm+bgmC1cG+lMLpECu8d3eJ1ZO9ihR1To1IFTJ8inRoJ73I
TQsXkW9uhMw9RpVX2wMVMV3fWyklbV5vc+ITp8sWBFmvhxIX738D63Ex5/dkDYj07ti1xBYJb52R
LZtoSL1dsvT0OxLL/ceKDZcw/nMoEFHtrWjiPvV6gNousHTwLPQ2yvwwPAj1hQV7k7cVBbNPgFcU
Ibqc7xdDwe8DTYjJ1Uj11YQMM4XqJLv7/XrVCvtgYbLffqHQtdzzUbY3R7W23RrrwwyDeyU95tok
qAtWZZ+wBGahbjn0Rn0AXbFoADduF99PTgjLnNvi5b1yhrzdmVEMTxCGA8xN3O3B2H1xwgWDceEW
4kUFo3KGPaw6SN2i9oVtY+TVJ7XbktdWiwnuZdM2xGTSAkVO8IcbTY0ctwD/NynuW9bMGf/mjacf
VT09uEHpVSz/1Lc/LaVowZtKtY6cOp/9wajfzQ21ZOW2hKgW5nLygH926JCHdKUqiBY/0ZfGz9ik
jpq6VGK9ajommiA06N4KQqpEOQa6SHcypBt1uCJEYjV/kPwryRh4m7KB9vYiAXkxd0XnmFlrrMq3
IG+3/WCQAOlLrNYZEcXG78Sw2zvH8O4YcUtjhgN19TnIuScxLHqNXjSVS0eOdcNcIXik06C/BQ6i
YC+J02qNV63WZys6LACU5pdOZFUulhXM4IIieN5PKBH030igCUDZ/x3Uyu7Cx5Ide8qmkbG0sCQS
kE25L4Y07aAq/EdvOuPE4HBKVUN61TXhC4YxS9JlSdhMQevfiC6hGotK7NqJC7izCLNd7ErQyqk5
9U6f2Z6u97F9tZxBubXTWYB773mA/i+K0FXN2h4sBZ4xpCjnhdzu7/iwGRZlZA0Jl1pxxn6jBebr
8oz/2xmGxancqXXKkhrgJ0a1m+bWCHs94DShvYVr3ha8WqALIV6JQa/leFrm/hkRbbeF4dgWE3xs
+VaxQp69B4krFBiDdtJP2vcgSyXVKMz8/KJIIjwwhlpIDQSWvQ4a8zsVJ3b+UKeBrPgJ7gdRyIWM
LDY9ac4BUcNDAkZO0h7SlL8ZQw4hWcJBh+R3szJ11BhPIpUs+P+mKYFcKjcfQCfyVRjizUiajS2k
4rZU7RN5AoOekWfUT3iAtIwRl5OwZkUgK0bJRWUSmlywmoy3XNzuEgkd4zhGmbTyVuuDw4n7gwxZ
1ph5i/oI4fpa1+otR4t0uJi95YePJE6GdOunBW8RlMBf/jGCKlX9hp8aXmlnNijL5kqWXHPRfxvI
ooEiKklebG68xIzTX93aZSCMG9IK5LNRBebmN4HNO8iObgdMykGWqSPckh4fFe+T86a44kkykUvK
Y+gvqdDiT/2GHfJ+WAQM9bC+ZI2kckp71oOvEsRTEOzjuKQti9aPe5zQhjUt6Pb5FUvn2DOzVgCu
TBf+Nuk11aZAYKH7G1BUIF2KO0dEPnl198fCV9gClbl8DruboloF5YEPLKhLDeBiWC/r7V/w4D4T
Aj2DSmP2NAiV0Pl5NlcMnRQMn8ato6WbJ3TyragIqUi/ZiExWbKXxRAza6qlnqd59an3IVOmjIGU
hsHvWA3nslvHp1Gb1atAj/hVlC0K/y8yBVD1+OFJVbmsrovfAdwGWiM1HnKIT4DOGynlxYuTNbMA
PbUAlnH4HwFdGLREwNWUtlKNDooT1HN/Wbbd12O6I7gYARKhbNfS8uCzVXM67OVRrUZ1JKXKCCZC
wRNw0f6P8VMFyeJLFR20jsOqjMVaP8X0p196QKxpd1Ke4gRYrXBLypXsmw05MAxKnBjyEsUwSaHK
Kra0x9poJpDPYMpG++UsNHcv1yxpQFHbH1XOQoPbaXVa0EJ9Xg/FFnIA9nBgD5eTIzAgfxf1LVf9
DvDqnwM124ZbLWBgNYTtDwIv2ElZJuGp4VnsElgNtNOLKqnAJgu+cd9TlYKtZwgoqETZQ0y9ChrD
VG6EUrp4qIBv8CovxWHALOv3dnZ78vLDwjdI6iNhBgfq1NUbm5IeRn7RJHGYCtEHOEF6US/NNje4
4VTqeehWA0xdeyTSbiRD+HHBuloilkxVq3346MFNPnf8pkqj5F2B6//9QOYeb2pDw90NHTDJJ6Pk
EJP+XQw0FFCoX1V09o/UA7+6713cJH6nQvaPXpAjhUmu0YiKbpjzDe4g0BNF417z9ZLb5lgXAr0h
Wjw4q1MkfgODHHzS6/Wayef/NmA5fdrtQ/AyUY7DbemXJEF7zlfuHeZMXnzzpBJn/VqlACCjiL7d
JdolyjT5tahgVsY4KjqU3K6pmSq+Lf58eFG/BIhBbjpmgsITmJJ1tlH35on6dTwru6Qm7EWV2miJ
rJasrfXrCYyFEAtQlF1pcS4jOijiGTtl547Xq3jZHEXktFIWfBX3cQNjDE4rEiJXxXh27AAqb/pk
XtLuIVAijPIEHTwiAVEcqxN2dHm+SDqgOI+/vm/FiJEdZG7+7UccTXT+E5LVub1EzLeIQ40uKwim
xvhBrRpLnxYrtaijnCn99K8oczRUqVK2EuDt4xi1tQ3g/mG+Vl07sBrfenT5MAJZJbnpPNuSXVrn
s4/ApinQRoqsSu7AI0L+eAH/qD7zxAahhY2zFjWr4Da5gYztCGyxfkiriQxthUw2TeXBseAjha+X
OfCfPF7RLwBcHD0olHpE78Jap1dhrrwBV4woaQodED8N+/+pfpIsl/WW7ChdGB74CUKHNVGZWKFy
R+svlf4WBnhLszeIU8FZK44N95DfdOrmqFC6+XbgGa6ACL9Tc0LBoOFgHHH4/PxFG4VvN1Ip15IG
RLOwk7b714XBCLYjuDzFc5rDIeq7J5ah9C4Ao1B5Dt/T7n3AHWqCbEQVNvWq/6DIeBkVyoGfg9Xd
frPSYPYuw90XUT+H34AIZWPud+gODVARDTonwvawY90TRC4VTtSOXVsCTMW/sMuSLj991m3HhjAn
2JBfkmX57pDuCrf1Efjp3cTkeYVG9peWos7vdUx8lDdgVU1lU7P476P4tIKH0VW4TFege6CMPtbU
MXrcJLai2E29fTk+EbRailF47e6QuBhXkt+jqea4/joHvBczDwZw8lazWEUmz5OGOQoo1NAMcnSw
HxiTr5Knab/lnwgNeIoGx8UncN2x9zbbJbBj/OKDFXpLctbk6VFZDt+15wwDpJxqpdj7ET+e3rQ+
GJB5Qe6RUjM9msCpoxp0eRxQ82Cvd5RtdzIXU1+K9u6aPQBU7iEoy20VzleM95NDnkt/yhZ9mnsu
odmnsKejulnZkcTNXDsKB7nM4xhi3oeQioSDcLW3QkeVScOa2bL14w9sgk33u155xQGVTgCMex0k
MIcTD2FI95+jQFOADAofDDjzRt4NaIpXbShdVGi3u2ZVxYMC+dZZb3KHTvPAgkymOhn8lOgFCVNA
htGdZBaBiK3fKKSBe1MV4xe7y8gCfQOHPFslYT+RjB9Ks1yO+kF3L3Ql+r3fUQLFALiZgCL9KOY6
Rw6YMnbfazbWCkPq8Lq9G879qCGKGwSqgnzueZaeKTbtgTtACLDO1rf9XDXCUocvHPUr8Aac6tWk
b8Lj9TkmHvKUd3ritECzwLMTdmRRNITsImnlCN5z/lOUI0kf5XFvkj+CA36k447yT06AnWm3/adG
uPuG+ZpGFLW6370I9bXYqypKC3t6kNyoeGt2DKrGqxsrEmrz66FYOrPz3I2cbt0VliNfxPCf61Xp
TuutgpTLeWzPdvoDPag9vzRFi4xR0SpNDD015H8RjvtPraF8VU5h+G4EOervnWsl/ncfaaKQynx8
qAsb0Q1QPtF4xkQzerqCuLafsNifoxm0wxz3qD+WfLkedMcq3AzTcPt1Bp5LZ2SJ/eW3O7sxC5is
FygIBxKXAJYKHFeNmIaXjFqsLgqV/Int70zB/E4eMgluMQbfirhqoxTIz2dOw1u2bZtyppiLOWEN
rHYzKCzHgSbdw3Q8RC0O+gbm9H3Mj4A9XaBxHKV82xmunOyUGiEg5ohIgykip7uvg9GS0OUQgGcp
WsnkIqy7QDwXDUftdAn6E1ptinSP3o+2fgC+59iVX+3tnBV1VVWOTqcC+8V1SmwGxSB9GMZrYuZ3
rU68zgP2LmzVCeS0yeBNWJtaECjspvcvv2VUMKPgOv/z/HMbCe+8nuALlksXx5i/if0ABoQxpluI
sq2zPe+8QdFdgb23LzVqYEPeRPDyEbU8zWQHDHb00hqgwRkGwElxlEDzO45A2XJJcry1KN65mPqG
PTq1IJFI6PQcR7uxWYLt1G4tmpRz1b2r2eD/STFSo4qDzm8kXOTbL9zXHEcCk8SFPkc5lLTaG4k4
CoVKgoINkyS4yHox0aQLLqQc1/x/CC4ra+7LKY9rFswimWZDWOnc6QOY2MYNMT8a23K4QAkDQQ3Y
15pozUkMksCEpNsiNtxZPhXdbw5CRnwLUEriJibT35BE+lv8FvmpAzBnp6iOnoanGhQ+uoZ13wt8
74u7jyXS9D4F6xWnOEavj97qhWQlb+F8QpPjz62uEu/ARUST7mmNiQx67HfrsboIcY1vteQtoOBZ
+Lf/X6742UkeASAnwFvcZoJu6/Pigc+pQ9tcnqZIOgAtsCqBTui50RSDQ/+HKcIbo2otBhtb/ssh
S5EuTZek8LsWlQcoC6tfjLm1zucDbO78/vea1CuNd5iePA6GwHf7hJVYYWlnZw7xdDs0F+MDhKC9
hy1cI0dz3nSDrW8YhGCoFX0VlnNCcRC0k/8EyCWS0M5H0pq7xhzZEcyltKaNugrsBTUuaw8aJtmc
R0RS9OVheYSYbwnz2QV99V2WoU+XxOtzvzrPW5ieOL2l1Adi7f5bTsLJCggI0Z9f4OOrOturvgrB
wS1tT6uyyPFyj1KMBGbz1fUVP3JPcbLeBvcAeiDA1BofHCeiWhvlSTp9npLwpYdzyczU0wA6qYrd
qrj4stg1xlaAhF7JmR8IquNceiPkXsqPZn/ZsaoeNrjDssq1MV2m80jxUsLHtnijvew57mM84fi1
l4enxhXHGHFddxhVzPTpENHJXX0in3Vy+aY6feKizTaKJh773AjsMlqp/VurHTVNcI6YYQktsjOD
GpuuMLD32/1jY0gUgwlcSkiArdEAf8IgxUAMSh6qoMIxPYh4Ky7MPDY7UEp+SPVSZ7R2dlusZIxX
TpgbOyp85rrHSMhe9Nmx8kn+Lnnml1izoNHn8EqB97bZbg9nkgeTE6t67CMI9f3IQoH2q93S72ze
fJK8VjWsMd877uNr08eVOkc25vIeK3fz6bnWsTNBkYp2GvUGz+H7owT8HmOlpoQ+INsffgBnyomG
zuAGKqxGg7Xi0ybqgzFBCZatQSgvargmBpp1K6AOyH/F6IA81V+PuDYu5SH53NN98wLfrZQzHi9r
WU4Yj0+kasRGAeUqsgjyneycKb8pwDxDZfrfNcM7EoUo7j26E6rRFXyd5Y3HWx7HGqi8QbzjeHH9
1L8PzxO/iLfgdVw201DsWkMRL/hiIamvDNyjkbyy8kc48jgDZ6sUZfc3XuGDJAFfEHwCy+4MV4TR
QzoWt5qub+EQFOiqP3Lks0tHheOUU/U86DPqoCtNFQkaGEYhxggnXSCVkLpiipN2cYoqHmkorO00
0Zjt/krvkqS+b5tB6fOK00AgKn1jcD+5GanM/+lEyYI86DTP2JCl9PPi78iY4NDYfRit8asPK6JQ
rsHbXtjW28s47fdLID9ENFZbd0V9seqsIhRcmOiC6xUsF5ZkTcIJxwrSiQ+PLne8O4gM16P+BMkP
Wte75hHAfvf83ZTTLWl9bGVt+upcTci0uVpuTqBN7aCrxg18FMkIA0w4e7QmmF0UdOww+qhKE4uV
qAr7wLlITu2b9qmw+1CL4RdhsHrlll5Zbc50w6byIkKGkkoueExwGfpmBNhw2vnPUhuKLymEivH3
Gi0O4zG9kTDzNvMWUELqYU3/4mDcKUCEQIS9ivENrUf0PHuDcCEWMywU/6/G0UDFhMYef37E3z6t
DjXfYFB4G3zddBtW8KuLZovo9Tdu0x9COPRWWHg9nxjjgKDtOEwdY2/CwTGixYHUSNyYqjX4fyny
nC65Ht5k2w98b1CNpBh47ebF2noikdTyz60WPrMoRZH1rO2ub26sG6I9BfgpUNwG9/+JetWuSrE8
gGzC+ycUjP3al9esIfXlFohwQ40017hHMBR3xavSYZhZH1rS6XdYpM8T2zWm1qftWiIPg9MQJFh/
IzFwzNoVogqZN3Ry96y5yIpF+4Mw+8WF7Gs170UPLACv1ZO5/6XiHVmkrhRw++xNIdVowmnHTmKg
3IAv/sELrx9qOkJOCK09zaW+91tw4nzhC64O/EXbbyHd1zB2Chky0IXXqkZ5mVmemt6ln/2hquqV
Usi3RsRP4ydckjzBlfhrfnMmJBE/GF/OFkvJfAqMc3C1vkeceK38bkRAphzAoA/Ctki7qlhSFIEH
PIeOD4+tpMBKcQkKeK8UIZxpVh75xV5ahO/i+MnDnYQydtWSu6f8P8CLNtWbhR4fztXdjjoPSFaz
Wrt55qbae+8UappVD4UuAsWQYhMcKfPqtEad7/rZYFmiihKPIQogaZPFdiaIOUOA5ft2Kqsc3awe
5zpdmRmW0hk0pVc9qPHWT8QOiethPX4yn3RvR9fgLCq+DhwLCbrKO9sTgk18B2zFn8neqelXuBsD
sRPW+7r0Tv3jkjUfGaBK4SfvhERi3Ja1bF34oNis6jx7MeUM+7jRGViiitrTQM+IJ3q6fJIcIpax
mXkzmP5aVY8mOpjLgky4yKdxswUwYSveYecyO969+BYvMbEhmi9XbuxDjr7JleGwuykJLGa8I/Te
XaXRm1xPkwh0EKZY0mhjHViYljXi5cbTWK4GZY3i2yZ45NE9mnFeDvzfMSZSENmBOC3u17NKxvaz
fE721oZTOS/v3br1xzQtjy+0CZgmhycR74uP0gepYeMs6zIHFZb9Y45IMPaeqroUNb76mQaDmAq6
tmRXU7hNBlkmdHSd7jxAxOHViyAIX3Wbg9Wu/rViYQ+6CyYPgy/3JgIHWjPdd3EUX2+eoexcsuUH
LQdoQPnZ3enpJiog41WFPbi86V5lCOZF1ckCdGtFMFmzjRGcakItTA+XQYRYafaGhx4M71ER0/Q9
yolMvUsjIjZ7u25l1e/AlveL+WVuXfMQaW9MCCMH6HN8Q37cJldXPlSLMyM9DK0ZVMMYQygujrk/
Gm0E9beyPovOIYaQ4jNloczu1otvHoFucHV6UIQuw4O+rw9KbX38nVTbDyG8o8BJ9lsWBv5SPcvb
/gvyxVVw6iIdyDbmYdzxp8LNxHnA+1AhhzV+3/IgxbBVz4WUCFv1XVeI3P6ozLp75clj9QYgqaCz
AdeDIvlefk/ApsnuMTYnfpLA0yrPJzx6ZowNezEE8oByxs61QbEBKHq3Z726Tq0/u6CX4oiG8gGD
LBTuvce019JbgrhQIMgbzvZQDbNJmLI2QBqVjEMKXfzv5U5qF+2aVBwh0HZgJPBJPlmzwDSG20zh
bR68euOazXfJFhr912dA+fUfTQoAxXJ0Xv9rsLedMQ3n3GPkFfs78nEIfVu2NCVy/LnNx/9f8WAG
BG3RuFoFm/2NJBqs85iyQImD5YU2d5WW8dosMNDnNI25NaxCBB8mi43CTUeBOiWJMKp5lRj6tono
Yhgj8i+ZwFe/mbSKK9ImX0/qXB/eCsRHKAINcStAJMg4eT1J1xYjIxfPKKtnaYon74TRCAHdN4lj
dDdgRbPqfOjGkfrwmWIhhJ1ZTbaJW6ze36pZsALFQ8KbsiZtbAsobEaQcxuZYultT0bjtQ0H/zn/
oh3L01uekMBAojJaWYPXHwlYbzthZMkdcd5RRBJXJtsyJsmhNnsHwEaOOlgvep0UXo7023PZ0yFO
nNI04fmtjQRyPE2evsAaHVBHmbdGpBeXzbULlMPqU63NCfUek0wEQm8ryzB6mJJaB7sTcJFI6wGA
lv3BHtg3eGHYnBnPvN5mOG3C+G+/ZdU8PUyUhKSHnbHmFsLiZfS6NU5ozZXsRuFjqpgZMTZmwWKk
PfShFH0VsHRaYlG0EaaxXae5EEXS+BZheOybui3Ld6+s2O2uo7lbQGpgpnaZao2n7mHoDxuD5iu5
trV8teaMIiTAH1scTU31jeos7Nhg0DWwTmbUmwqfz+aTApryFCoQEd+5wGF3uZgAyIaWOqBn+beD
WeRLF+utgqiYXF4HlQTJdJ0odOm4xjZp6pdQIF2i1RMkSxj3vwKaCiMYPnJjt/v7lpjGslHqL0E3
BOnXgiUUBkgWCMRcivNbngpGRhlduAc0o+actQwOLyLPYkyBQU5rBsP1FdeyYW8u595FtfN0dwQW
U7YHleTZY2+O+6KVzB0SpENveBqThR1GJcppWmXQjHgD/Yiv7dsRHeJDl5YG98COieMGdXRASsRc
iiU/TIPRYenX8Mh4weoYnJgfLU34za8gJN+aq8B1s+K9jVdUFzGpv2z3KsqnkjZDYHMIT8oMzE+U
4Ua41MtBwbPMtFoYYPvMH3zpOColpJN2t95V9MxNJy7yARf4xTQ5bZjRgHt4T8y4UXzAVqKWAE/9
PQOqQUSl82gozapW4CXgeGUsfkiJV1Z+eXWq/DM4t6vwgnwZ9sO7ql8gHZlLL5zlWeXqXZSdc7KG
3Z/m4B1LTY41K/4kpxz3vCVI2m2Gaxm8O3NWC6GFXq7pyO7jU1ICSihQksPJKUwwdOf7lTdFGEUD
9/UW0Hd09ZaURNgzBJuOAtPren+N2nr7giCTEHzIeAXWuE5oOMUW/HBxwzwDb6o6M5Dk2zqSvSOQ
f9Vc1Q90BxmyFwcd2D45/OZn5jPdBbvFLfOWJrabLC4YIw6B8BaEhgJ4lguOzNbR4v+N2v06v5CW
RF7zVeqvE+ELF9PgW9Pgw2QJ6TUWHJM1RIJTDYpBNQw2UxgZktOo2kBZPBvzUTVs++sBg4VkjhT1
ZNr5NWYpwAiBXZJFigb3EpbxIHnFsauKEJkw7mCtA0AO4RhgoZ8AkdxFl6b1ohS5Zb2jZeY+4dgl
qBL8AXjHyJ6+6CW/B9ChsxknyjBwDr8rLtkEzoH5xu6au+vj03HtY/tnGSrB1l+9Amt3bc1qWvnl
wyjiaWgZngVejaJdo2zayt+LvcHA0ps7ZHHRILgU1vg2aOlpwqp66seBlGPfsnGH1rPiVQ9gisRV
9p1GJ1nleRNIIK+S8TKNus7NhU2yuDeB9Wf7EPlJKx7VhBtqSTtioYolx+xLEKBzD4Lj4RtDYBfs
SuVdiuFWeCkBs3vQQBXAcXGMbKeEOsvUm86TavKWWeA0T/dwL7R/oyxQp59rwW58cURzFfle8rJa
TMtY0wP5WuFZprKsH9xRyghf13mDQFkxK5nLMSNTQZh1akqlES1TcrEHVGn5jV482okEgZlRxkGd
BMz3XysFEK+LL57QOkf4rpNfgNi+1akQ+CQAgR71G0nVGguRYkFRfw7RCzLqcTYYFw88iRl5U307
HCitE056eJGEA23J/FHwp+TTLY+xoJ2BnZEF4fdqbkv8WRGKcHzqDRsbarfCsfJ4McUWG2Jg95FD
0R24OmMWS0FTUVHzuoPgHkeAB3qEducmcS32HfokGK0xXvB3UDhhCtNyqdJliPSQUQJax+05Ud4L
iii37l3W0dKRRySiBetsYe+Dw0wp0vaP7Cvt+iJBomucRV2KmdWyQYSUQAiq8dINCaCXsHwTWhWA
wHBHmJ2bQXnXGPC+8xXKn/RspDy9iZYsxDpwVBs7WOPTnc5yQVT8o10kB9OeCd+OJYvWkbkbNUnL
Ogu2hpbqQRPMItnWTzw90zReuwVLDI3Sdohf34/J6if1RqaUg87oZ0ibVh6Ivmp56r0Lfe8D+r2W
h+FqDHwPdvNTgfKVLRW7t2FUZV+bpxMRaJvxzVWNJSSqispTTEBpDkkTGgXRvmsVRywBEewJ08V7
kn0dtP8LXpA1Uvt32YA51DgiIcT2ym6Z2qvhIVt0rcTQUshcJCER4QBvkx28Z8+T2QqBquMVilbw
roXU0yw2EXvBaCF7ZY1Sc7bYsIkTQRSvm2cs9akrfy1FzhatohwOjOb3vac85HEFzUrHIHmV1t0A
E3rplq5651J3gepuTntaEYYErMhLpKzB/e8xZgZ/0qZWzfwPMKPr3Eu6NvsIIl/RsZTqT62qa8aP
4MQINDjnKz8WtGM3kSyjzcw8tR86JkOqNk5Uqvpr2H3uNei+r3wySbNv2RNwhol3lrQ1tIXYp1hf
WG3/TQMl57+9jkneH1AdyU91aUpFaiGP+zytsWgxLNq8TJG8tt6/vabVasCO2uikUDU+bXSqr2TY
OND2wKN8dM+9Je7WY3Yk3HyO9pwK5/tt3+mwETQTH/639qIZgH7V6VhW9RfmDWnb3gcLXBb8Ydw8
157vRV8hrFbuZvqBeA9f+w5NMQOV8GFAFtmrzv0iL7vs9GpVHVUz+z6UBrwdZMiJYbRgfSpLrCAw
dW2Sn2btQZpzWTWHUWl5953P9sg/srkilfjjoPLW4EoO3dB6Wb19wgCUx4hi9+vJIRmttSPi7DBR
D4mHL4tzhYTr/EfeJVtwUvCDHyYs2HvfUwMjPjWJTswzO1tTVi7RYB0RCEU8zpee7RIDhRE7RZfW
MCNU9MSEBFNNn/2XmxYjz8a8LyDIG7yCQoXtsV9DZB9sHUh90t2gT8v+i8RiSawrJ28hHx7g32ei
EOe6qard0rz+tkWZnykpoXA8JIEcQEXztM+jLPXz3SUTl0rS2wlZ4YghqeTPXMi0UANHmJqpUDJ8
K1oOYDp3Vts+RaIz1+1cigOVZ1SJ2JYReCeHuwLGF5B1Q23l4i2GuOahd3BgZRa200X81Ep2RR6y
mBzJx5SX4Cwp/01AKVEx7jvvUfruGnJXH51Rd8cYqjceW/yYsX2GRyCYZMcD2fK1verm5i19VSiH
0CNoINNwj/G1V8qEELM5fmOWzgIds1VInBhv7jdAmo8B9EuqFazdRsJ9RnTSp3Fj0FZiZc0plzgE
vcGAdeI4ynrgHfcyzFaZNvoXU7XVtMR4kSC2QO7WOGdSVjpIho8py/Jk/1we5pAhI05WlEalqD47
S12kA1y3IPN1sGcTq8rM/bpQnN0VhpcxPzrcFyt+fwjptlAfBHkschSSSNMvOz6k3efzPolpcFFc
7sFubTj1z3fF2GWE/ojxayvoB3Y1aY76RRKkzqy4TLZzf5SsJbTs+O8ppRwZB1/CvWKE8GZSiewj
GbSZrlsdQ6VFZzLzNzxXkESKrp1z3kriap4836RfM3iMCDoHhMSynluRQWVGwkImEYTg25mOn2yI
t2IoxpuLdoH5MSA3ZZUt/l/JRyg/TLBglhXdNq99fIMJa3DCjmFQtjTfMJharFIRadZ9fDCHxBvi
6rx4LTwkuEZD6REwHS4II/sTTk69oiWZtOYOIeRLszJk5O2S4Oh5IVlhlO5GtHv/M3GsN4EYVBJK
/NN0fVCJLCrup8lr1i7vHaFPC5XkmP7O1PgpcZezIXnTxk+U40MCn7GvKyWPfW3gHDVCaBvYGOGI
mYdD7oJKWztdLNKMs2PmuDlmCs38/WVeDKmMRffMkSKrP2C2Fc0H1f7mDbNWrdHBqaTHLesKF9y7
XV/E7yU/cw+7IPZw7XfVPsSusqCJyfYOIkgD5YlPJLfVw1O5L+nu7z0uMI8Lyt/G1IN4mycLAAHy
bJ5+S7zIb4zfh4ikdCkrdqqJO7clFmXWBxliCNMLcMbXbyppQ1X7gJKjPguBSOJaThqOTkeJbBru
qyWcO/fvobkukNRh6xee+opM46+RpZoOsJNadnHLy6sD8b7AGhZ6kcubuiQm4D4fgTIxuYGDwwwh
zOa5A0pO89XGQ9u+HBoScgwGhMdQ45Hb2SVx3OS4YNGp2azZoSmMqO15IzowZCPho7JweF/VUol2
L250cTh790uGCH6aHRGguLZbo5SDRUyYrkiSA6KSVrtCzEh6tfJPS+JxEna7CdaDqdbQ6bIFVy35
Q74GK3+BZLk0VT+XMkluoqsvasmBf6xozF5/BirhLI+Nf3rpIeiY9gwECbWm3OH8JjggEG1ZF8DA
3hso0IyDeilLZvcBW84LKHmVNk5DL5tmBXH4qSNiJhhMcgsu/MzxCHCreDART9UXObzqf/ES/fi1
I/C36vyCBFGQn389NVfvJj7IkbBUMbToXO7PPj82PE+u5KFkUJNnC1emcXtKXRbQAGTVgfvDCSWO
NP23i5UBHMzCiqi33nN2FPCwuRq5QWg6+20XDbADUbED5qUKXoe8wBplC8qgkaWYhCncxBdh9iul
hevGYAFNek9Jim+umWWPFSqYBaxjE/UcEiyFLLGanqjP6XfI/BarSX9ep9QrkWKvcYaEZs3zNDVY
1Q2kkhC5fPdwl/jagZQA64tYQm0+jXYvJRuZNnpinhf8Kh4rZ26SZf6Y3eQUT5dV5y9ePgHzbjAg
VC2XxK3Y7DRLoDZykk/Bjd1NlbEP8mLDUMAIkz+yn85CHF99xbNe5oSDbBNsrDRI8yREBc8+/yCH
8ZZYJbONKft0QpJaYVGl/qoSjO+e43UJGqzsbyQJVYvoDKBFLoRjgpkaMP0WYcWYb0gLIe8opgtM
7xy5Y8HwY0Cbln9RLp2M3APJhZZbr0SQGOrrwEjEAilRw0udtOC9rEHNGHNEu/Sl3ZrxqDwGEtoQ
JM9v6+TjsYvCLkwzuTWbocNmnJQVOrzTvGL/j0fpiK/xWBL3GKRgFtYty67RpjEXG6az4g3hW/sj
ldfxqXa+6VW/WTJnhwWiY8d8KmdZXXkR82xOzFt6TcSXUPNIs2U3d+THqZXLtaOcn0W+5UEw8CpE
VgY9F0X7C+RrLKTjJjYrx7VKv0qddTYtPfTrAPhxx8BTQ7Qx0wKKJrNEwi9doYSXaAH6cORxU7tc
eqGSdg+LZ31M49TIczHiwZLmjQVaCSRoi59KiqXW8fIy9ddluo2xXOynIBtq6UcKEdeD/edZhBO6
9bEWxYQ/n4J/OpL69F7c2LhtAuwbLLTH82qB+QzdDaclhteBlfQlRTsmhIhozxSlpDGjUJyAtQeQ
ebfIUHC/deF4tgXBZ6Ot2OqDrNRxyKkpL6uErhHhfEGyOLfsqLNuJ+HDSBZS2k5Q7QJuKQXDM2Wb
BBW9gIyKiyfP7FhNWIBpPZJ9O/DgpExd9uL5iFS33FloogGuaFw8DiQcVH80JflVMzdiWO4LopvB
+4wJBwzVZII6JcxcKXQ3JQPoQMbqathqJd2CgBfqPx4APmaV4ooKG84v8Qe7fSXzb60t7Es7XfSC
hveFhPVVkcHg0qS8sZPCbby1PogdonWqoJaeEUt9dmZjqHjnH/IcHQ0uSQT85BSiQNMUFn30p31q
JPYQkOt1NNRu+QTIIoAwXtxwk1ONW+7fZlZMb39YOPGv5Du3o/M/4gaNrMwJAPjws619K9pVPKqk
LFQmNSfZ4jXqlvR27oouKvl+G0Teka5U7RZHsGGrUjHumy+laFVzf3fqx7DgcgB9x3ZC7E70REKV
nO63sXhgHDEd179npZlQffAVMEEhAdVYPd8ECPgKw+mmPlfPHQPF6Ya3ry5ooGBNohHa0aQna5em
W6a0Tv8Q5pbJVwDReZZlUh1VlfnaD67PPneFij/dWi5Z21SpnjHxAVTIdlxsbqxWMEz+4fb9IedU
iaHyyLs9cbWjhf3ucQklIbrFANxPybyQJcz+TtPD/Qe+6pvn26FXpSBdT0kmfODpHNIpvztziqw5
OVYFy8Hs1E7pp9inioasgyv0ALOTZXJ+rEmn/ue8p0VmIAmk99aNYB/b5NnLiDBqQ3uvco3gPbXK
e966rf42CzeDbpJRwLg8+e9AvICUAbrVwS7++ljoUQJhZjhR5CuWw/InRkzXQ/AFD14JmE5wl/RT
/RR2TYEt6K7xmDlxTNc/UlUiRz7NQvhAEFqQU89ZchfhAbEHmy9GL6p4Rp8DwHokqaakW54TxxWJ
464/5v0mEjLvR4xhgXwH4Wa4Q/7dmTadwVfS3Rus2acA+2zqOeAQWZlNmIvtVjN2q+xFLM1JNteg
5LI+AL7kaJdIxcK5Mg3nJONkKSEa3CmxruS5cNPpaTuKvRLR75jKfnidP4XyLRqeXMn0YdAcR9vT
Yw9MmUCMe0n6hkeqxLPewi3sdUq2Un6zWCpu/BAYmuK75kSXPoqIQt0DwT2x0yCC/B06vpLTNvWW
uE9c0v7eMJCm1xL19t/fd6D1a8a6iITkLcafdZuJNCy3vgXQ3VUc5sJ/rvYag9r51/6Z3zhVAht9
vO1scYf9i4lyo38pbFm+xbUkv21ax/Ppk9FZuTVmHiMTnRWIxeJyCbIOSlgqNWGtts6oaKi+8kns
6fl16wNPAwbefba5Eei9dTX3fdd6huh1fGYp/jX50t/pPtPKwrRJi5IVBGsQfglWxWWTvdAlnKYe
S035h3lXtKnmXUGlltzi7v99S+hEHR8QS8L1WFm1lO0IRVhy6eheDRd0XBLM6VkB2ppyfm9qnASA
egiathRWq14N2tfSq3bhPQoieMpRBGIgJEACrFfiV/3exDivYIsEeQS3afEnjfdazA1CtsFsGztA
Piposx1OBCU4cerom1WIJ4y5PjrMvxI+oIOt3HnRgMOasVODIl7HWUMiQDSQNaQp4Jp0sFfYnr7h
oXFUasUYwcaFUu3zpZTH4ZxvLDPHwMZGTaTOz6E/mgcKIfPSfBTUEvTqF+WLYbJbdkLfVGekgbyW
7gEy9/tzfKUo1CoQ024IoInbtRewv+Tv5THoQurCa1GrlE8YJNuH0ZKJPDlthdRW3AgIKtfWJ/W+
95jp/qyQj3O4s2iDypXPEwrU3RR/ZFGMAGD7yzeYMed4D06wDuGSGc+rmFYu7b8Mc2DHL45m6/f3
pvgDPZDu7f/VqWHgUxCRxVdTU/0vK7mGrgyib6EtPOWTCUY+xVpgfWWp4yOWS3n22/MbALNiLv02
ABmVsj+m3q9X0r04qiDhXLMUuRAh76cZZTuHnqrWDMk1fbujQmKtcxbq5rzEOKClf+uc6f5G3aVZ
P7zZK3Kkk+DAM4uqwYcpM/8pSRwOZXktKwA+QVF8a5e7y1Tu/1wJQ82ga64j87itFpMkKaFZXUcf
N6TGm/52uYNpgevnQZHtSWD6vVPOgdNRIkTHRhPAMpEQYMvfGgOiuc/SLiGOcaV1lxz70q4HYk4M
DffHKkjvshnE7YqqQ++89r/F1HZCZx58/Yg8hFY5VVKH5torjRhOhV8V+4P2BV9zouQs1w46G3DI
2WcHl5UmV2/4KR/QFaHSjRlx8L8b11rY3vDREvG936DfNIVytptK/SM45gfoBLRVuoLOPqYQXVO2
mk3v4dw4tNR6R8WH50Bs0y4H5P7xulOAIMMc6u6ofybIh41BA1gJ81Kayh2r4V/C2LifFkA0EN2E
w6ZqTECgjmPNwyNS/kwMyRV93kjYbhziB036FPjHCn/7YgiMjQjHbnqEFva9DM7TJfs78QqOxPva
Py/Q67FQCE1Exu47d+7jwwW7z1fSvJoJAfdZlluJK0kFLWkb3+rPwPFGbhI6pCgcoAG5yOCvSYOY
ObMSdGcOA3YN+iaO4JSx86v1NFBjfyc4Y+UxMaARk/jZ7qSZhutdax31iEPs0aQNpr2xvd1scgnZ
N5MycMkVjGqijvPLVo0+SulTDA2nGNgImfMjprrTeTyOLBgpsbZ5vLwOIpf2a2ufFlPACQf0a72M
Ws8ec7bfnVRGh6MRYjl2Wl7qSIBp4qX1rxfDtvTebT2hzlh9LJr8s0INfzPkmeduxecDb6OZqSFK
M1BuEYykMJ9DGUKH6hzlzE2RSiYwix1641W7ikDqot7fMNjXubyTXpQvwH3JjsS44CnHbgW7W94X
Bc9kNLn4CK3wEE7xB5UpU77JDdDeuFTzNiTrtodLbd0DxUKs8IHUXOBTv0C0op7whmEfDwwMfOv7
RRJ2faZduB+Ib0wA48u+2moApLbzSVz/Mt0MOwnM3yoCzgGcca4z7mWg4m0MXqiICwY9xs6PPw+b
dLpY0n8FnBuvU5+LtJv3QiXUR2bMub5hSYIYEErinZyjaWS0aNRkgupqacLbc8Zu/nSjoQcr14Gz
mNfUelCvxM9O2EGja7rpfDYkQO9GTE2Up1sYpUrPfm0W4AIb3Xq9Z2BuYNL50IdNkIuhhRkRZlzJ
OQxZqksgUNCphnDSvrWa1kRS/3IteGzaChrB19Vc8Tfi/UnpG32q4tUNtyuBFzm8m94TqrZ3wwCE
TPe3KH+U8pEGtlTJPZlfws/pa6jHj8lwummLYSe3aQLrWUfV9mYrVxxzJYpIP97He/GuhTOgnOF3
rFBInXUIvS20TBGFgX32IWB4yzMlk6rNnfKi3GtQzB/Y/AoELi6WAt+fO92B+DYfMYvThXL8b8ay
Hrf5yG0vnVXrcitrc2Ls4mA8Hpfh6sBAJk0du0z22vTyMLBasD47OVCAVtPAZkNTJEN2WVkxWLiI
wvP9I6ovMQjTbKMw+SC1dGCkrQiog4dSXC+T4xjhrymcE1Vuwj0557nqVz1OL9dpTcGMzSFXZXe7
maLaDd5Lyzx8endTO9Q+JOJwD2hf+GShsrc7+mWXNHg6rw+qPeYG38tTfNY1C7fHs2NRnMmiayU1
6Ghv5CelHstNuz/S/3KsZmdvMlefK5AGvdrsbrtU7kqPsO7gh+2xnnDSX8yuWsb5i1iWVwSirKa8
qfTbK50fTybkHagWdd6VLAtytFRNUdGEvMVp/A7E1J/6a35CKFUIDA3UllVk9ApqEiveDIIxL+Of
EtXAhkqI9sGqlIp1SIwB3vw+oncFtpKVek771UPtN/hyOoYen3bRplco2wY4JZ8Pkx1FAqZaYBlH
ejZ8KDsqx8jCVKKePaEsEHM/qhd2WQfePfa2ORKZ8KKQGX4V+l4qrT1bhDsZAEfrPOL3q9Rczou9
bSXQGiDsikDdk7JYltYxiG+R6ToddARwn+gMqOECF76pNDFKM0e7B+bjxRfgPtm73zfZAhHymn+W
Z3jvIVp5AiCfEmkRBjzGKRaeTm3gZZOCNmfPOgSXnJ/S+3fvRFT6mJJBbsdWUCTDdWmLW26q3m1m
fV06LEzF3TNTY8EJBg03mdpidGjHWcJYCQuzhNbz8v7VjtsIQJXb/wwZH946tEdHXbg4+Qbuf8gi
lUASEvgbhZPWXmjY5Sdy3cDUoniV6hA0/pmVfpoKmMRWMwbLVYkFOyF0KyRo8kbCVVv+yRXvFASj
NWPUsxZx6Pb8aJBbK3eo7esFGF5WUEnzbNP33hezhiAUqs+9+eG41RNOudkB8oPS8P/CAaEbV8Z9
h0UZVe9TdZamP7dmbKHwCceZH7tGqAnDdhlsQFirXCzau9O7NJLmUifgp4Tb3ceQHp48Qxj7sGej
+w6UPPTGg7RE7QbVZ3mNhuxwjBSW3uJBEdgZl/+S6WcfUtazKIpgO5UGvGlfRKlEIMxDe0OLrbfg
N9T/hOHodZ1GtgL0skZS11PDoHek8ryKkPXPKs4F5BwPY+s3xsUeHumkBflm2y6bg1g/xVZCGL1D
gF+lbzxf1eVFexQvXukHdMpBpz3dsg/V0NlXXTZI76tHhebFV3qU2Ot8lup40BV961fkAa0NIPEa
ITDCnqqNBFjllPiGdpsQxDPQAYVq4gqAJ7UoTnml8TghqG+8ZVrTkSR5KafVhX8+d2WkYsNDVDWA
5a+jdg5waxNBFXcY4A+2eZizD1NRamX8U9sRlXAicBnVoBHrfu5c/TqtvObTySak/jK4jz4dhGEk
luaomM09Y34FTxJL8yFHd03a0T/7GO1R3e9eJrlXXLXETjJDrLHAD0ed/mv7/lU3LXo5gs7DCAnB
0SjGKBTS4XC5TEXs49t7mPLU3cVJL9pryH35By97xXi2cW/P1H3FiKHZb/4Lv8l349ILXRFTYgjy
r3vDXPfNRhAcx7Ag3/VT16SwzmHqFlTetHQ2P3tyFbSRM1pQRC2stuegwVaZcxClOhPyiZYhGOZ7
9oHuCPTe4vnUFVgiCenLEbkC5yRRxy6HS6IAaJrZzjWD5Pqu94ITPphf7cRX6d2s5CzlfagdXnx+
NIlwJED7frrzT2TpPUDwnrX9LSdMc5lDxmEevP7+JMM0SIyXNhRPVhhIuQlM8ZRjBrvWxXvPqG0l
VMopmJeHFw5FP3KYjzEb3EtE5W2EvIF/l3jIYkzhYCaw5V0ybAlnT1Px41GTcqwe9hpprhIKQRpH
iiI4uG8uZ1SFiaNBx/iaQPRMBDmXaMh+uIU3OjEUF0AjLrrsf3HCSGJFg+c+FW5fIAtBKU9r2XU9
/aqqrM5CeJLXi/QnA85q0GEeTtvYVrFsD5nPKAj+OmUwvGK/YBUe6mQHB7VfYosVP8mgCC0EYx/L
0RN4SAZJyTU45cgGN7PgUFFBhaIdl3IQyu+M/BZ75vdlP9BRm0qfTExsH+wDJN0PPtQBWgm/WtSQ
WmMtQy4ouhJTl52LO29bo632tTUPeNoaSxIyq0l6MScnZZfE8+lmcc175v+FBf9SKdxxBTTI0U9f
RdKIfLRoAVZq/wVdcNss5JL3DrN4DPuqiFsmoDO8aiMxxPjbTKjy/f08u7TP6rWKmEroW2KHz1dN
pGmhqpcgxe8oHEAQ7VU9TCya2rQg6ktytTJNuuZVZ9cAgTr3by+RkbgttbuvNGXHM5UT7AziU6iQ
44VKXyk2C9Tr7fStkfPjJ2OdDRFCxR20USLVqPOjd/jy4KlXGv6ePKoVE7b6QKoFH66hwJ2Gepi7
pXnGcFbV9OeCP7cPfQhtqUACcH+cHA0AbrdOe5ig2zWK51ugWmvNFWGu0r7iz+ia2GowduBQM1nM
lDRtg5E+wIg+NAMKGYzLVrGkCuLOkvQsp/1HqjSxfq3/1oDPkfHOyybQZwNZnuxEzBbso12aUyA4
NatUZBmVOOQVGwAgoCMryRUi6Yw0RQZPv5NAV9uhOqEeqxcqDzsoZnd3zzkHqluMpCLpd6b8WQxs
L4C9P6qUVQuYlQGtiW+WsuDbR8CQ6GfAWvgfiqI9gYSQa53dCiDHZ+twLaK6F/xQgVPyiBMWNaEL
PZZMD+qPVDt5LIr3zGlQtUzvbEZovE2I+JcUEbjZh5XTY2qLjBglqgmEs/+Lkr+AxiRzAYSe71Yg
b+403zZz7jjR2yB686FhBI3ytXjOFN63rmpCu3WNC4aeqsgNLIwP0GB4xgx70PSexrF51YtHqEyF
iHE/Ublc7qot9j0o0R+wDw46KVPYV4xQVFBqT9MTFwiXUJW4YoGyZYs5AuIG1jBn+e1VK5oHj1s4
eaAsj7KpazHS4t+WTZ8ADjZWCZRupe0Qk600MOqGGvgHvs0exbRt+SD9zN+gwhr4NVVLNJEvfKwO
pbXShYspcHBBwTPE80Dur73tint/1lkkHgYGKZVGD0/nihBLA8uCsCo3ZSMqxq9P3U9+5K8CF75N
5Yqytqsb+4ym4g7N4Fcx4LbwhqBkH5EwftrguxmNj4jC37mYbutLr0Ue53Krw8QWUBkAkmxZV/eN
MPTjDRP5YjwqZIiZzpSqJ4qlSZSASdY6eNsXABUCB1040l2z6f1m+gIxXcx9Jm7eNcgtuZatYye4
U0Z8E8yvZ6t45Lw8de0WasUfNpiNaArag0xDl1LX9yeuNAH7NA4ABMaEAAlo8ywJyd6CoflIKA1R
JxtDoRPHlaXUBnyFgduSl1at5n3r68srBuVAlGfe9qW938Fjm38CUE2XFyEMm2XrTljDhpgbVzr+
HjeQqW6wiVSRJBcRZzxFsACIfVpmJbb23Msgg0ZA5jQh4I/TMRusQtxQBAnnxaXm7hzVqBSpRqyF
NKteimvVgd6vcXlZnRND0NyGpUvZEC7Whd549j/Tw7HIDtjpPPBVxGNtekyULw5IRrB2SATARIJK
3kUqxoZVeHWmV8+8UL1fUNSPsSDizoIl7QkXJ0KpjeJjuNNSrXI0yXILnxBtGUBIUvK+8CroY1Eb
GxXdmQ23ySIvNpbaT2VK+EhIDWkKu1Khql1U0VGAOHRIzqgLDQWZI7mjUuJZK2HZH9yHPu5n5cWn
jmEHqAWtDx3GYddjZ76pA5q7d2Un0fx3RWsNeJSHjjhf8jibKsjiGYSZuQOmeEzAy9W+odoOv52z
MXqsOLZbvY8lEpk5U+i5wDij7mgLZoIo5uWHEqxKH9ubdbo/UbuFa4yhM/sch3UTIQWvZT/FAzRR
YqdCwzKvRh/TT01jBLQ0nC7Kv2vK+9vbrY7kzy5vhjA70bpUxFX7DI64qOtzQix+NqsUrZhJsRgz
fwU8RTUZxVHWedKdIi8uw49dulFPANZFYh7NzRbR7VocwhNKOztTf99Ht4TcWZm0mEqjk9++jGOl
GpBrpdzJq+qEx0Sx/d4n91Xk/lgiVNrwbD5s0+R7MP35PDXR34yFr2c/SbCvBjjxINMd6m5Ef+R+
gWGimlS4GpvZXbZdMITCGERyEey35lxdNiJ01omfu2TarUVTTRnR9G9+WFUfdyZ+UgKsF0+fwD9l
vH1OBRMluThuSZWWPdr9UL/IFIH9Ed+vf/4mDP7fpybuZvePpiTvynhZDDDjKwn8/G321VT4rUvs
0zriZe88aYng8TGJsJKbmyvlgM2COWui2Dgz8fVxH2oOyUYNPoM/7Et+hQPbiFkvhIczUId8Bat8
FTx+NUMUoqpKp7NdFE+7UPhzeyPibZKt//ciJbRYMFjf4u4HPlKMvr3WusirW6zDZyPfuOOe+K7E
Sr6qcVIc159w24aKiZul1GWNaCg+zL21iBwYZa1XVOUJDNdGcUu7Jv5EbvOI3lxwUJQpRlnZB52d
JOzFrt4zbCS20Qoeoc4RnlD9Z7dwob98ffhEb2bmJNfSeaY6IJMQqiaXR0fZEKH7kRl60AIxOJ5l
h5HDAfcPAqqLSZNyfdwPNH6rHxEkdwfdfYxXzckLQeHmNCE0ERTIIqGJechPU/lWUDuUWyHKmdxe
7D9PK6uSWs3UHrh2bRnE4QdJbsiH/1eP8LxrqcoYOIlZKComBCRVCVhRo45Mdv8e5YT1dSL4qaYH
6Yq+Z+tKK8VwZ6GFy228G8tLWFip5QmjnCXGlfjMz/khX/e8Yr/suRLVHf/pdYQN7HMzS+S/Hiaf
iL1zQT4WrCeH73Ulh9+b0dDjk+vPQ1GtZRUvBLQZv2JmTHC662jyTuW7FegsDX2DvI/c4lpgmco4
QK//QGJ4aH5xzqfrMvlrYXP7CwVVecF2w6N9rT9aUNZoS/VB0oxjGzlLG1hXtJKyUsTh0Gg1dyJL
QzlneAuWxstrx8SlCoihRBEEiNFwv8v4uXoWkf7VrUKstMe6Uv0rN6XsAKYE3nOZUbWh+QhyafY+
PrWq9SjKa4nQYtmIBogSfIU8qr8XXzgi1+XVa/TfQx76tX2xIrqs1+TiRD9pfRSTcjEqSmIafjQn
63hqv0fDYxCf9/BXP8yF6I1+X5pcmnHLu9t08YClahD9K+uiYlUZUUV4GfmunNC5pUqG6Q3DuxYh
gLYkoF4Qog3KE9EgXEQLveUJ2ZzSNKwa0tcOCSC0BsnSNM9WLO326vi5mLkQlN0eMekdPQzaDME3
1XVKreJzv/r0OPZqg6ASRXuVv/d/MY9y7TZ9POtuGWq0wQZbFxPZeVXlFoIIgzNP1eOeh2vCP7DA
6ScAETguemY3leLmSlHjhb73wMwEN989SgAg5kMRvc8AawSuDIpZa4Xzfi8JuPqqX9eRZsNiMDRL
BOeT0w16K1ZTAl+Zq3PBDYlpYeXWdNr1cnm69zUbyXHBRkYOKecnqtZheqkGa6cxysf510AwJJnA
ceRGPdpkawO7A3hKOXmNy+7Sm0Pju+iTY4k2iHZs50aPC8JNU1UFGTXPEysGRtyTNyqJrGJwJnfE
8gSPVZIhW/lTBYJx+p3Xklbr+4cndofwJHHtsKVK4NBK0xOSujPIEMBd3+SKQAVBEXnX2QmueDPQ
DFLyaHx4kfQFPjnJfOjM4lrb3JUZ+2/c6v6PYzDNLpX1HXTCy4Cbu2rkE+plkY4FAJzy4+EFxRa4
hHvibubpGJigMzC3aluHqC78HlUSs+Tg60wW0NeyQcF7nblOUY14p0zH/lPsXZwFpyAgRmhbB1Rp
NzOndExAymw6iiJ5Cg4kPnggWYbS+Cmh7G+FPl8ChVzpUzBm+dTQ4DPjNGJor2CeddgODEP07+bX
buo25DrVVn1ZvndmfJGqqrwdzsABYTvxOHi+tQJdGCbTPHMuuDEe5dN7g0MJh8bxRjblJrl94c5y
HXWaQKKhAcu5Q0qLqjOjgi01+TJj0cV6I+/ZKgmuyH27tO2oB298UmtWqMpwl+/AUdXbW9r2tRNa
lTFtKaa9Ro6MYxLv/0cWifkL4txmrVDYXhpOek56JET27u86NcYSFZtLmZfLSQ0AVoLqtW3d2paD
VQvMISChEIHyfkCxwCNqrs4EiXGcgpjBNsBHiDbf/MIbXeIrIP/yWa5lAEX8gFxmaqUfrFqu/uY3
23bDum7WrnTImVGG+LBlKHkQ1HsxuBsI7fnaaMgwo2rZaDxyS2/7o5Yo4DyBXSSmfq01lsxqbNdn
cDUgMUgZdrk5NuQVA/Vs94zqqucV4nKDoB4UZNVoslcQNt2gto0RWyvrog8azmNmUR0vs25guQyK
3wVXx5jkQevj42UPGqOaFun2cUtLthjqFM7RH76RoZCAXTnmP64SW6rCX7ZML5+vD66fNAH7gVMk
UV1sLVU8T4O3H3QuzPhZof90490FaEhJfmz9i5VdtWwBB5EdnJMYwkn70DRQwxf3bT/bX3m++m6p
ieZZqxKgwhS5Qcm8s25LyHG0LKG8OQMBSbg70Nc6BdVUE8KP419e0NRDlPcdeWBhE+A+fijKT+it
bMZELpzULq/WAe9c88uCV/uytl8ZP4OMusPT4RrysFvgvX6unBsvtum7alhZZbZm/G6OyNS/wv10
6G1aJoiWcisIQkbH5sLqMo4/txwajTpEhuww3mhaQMDjm5JDhbypH+QQ/FsNzZwgDgYXCPkfiMf0
kNXeyQFcV7iKQDqCrIQ6Gb+CQ1jyoXM3JYupTJoqJyXLkCJzoW7eGZtBiWt12dZl4QzMKLS3H2Qe
zC2yIoi6NQKAgzp3B0kEDpe97STiZuMsqsIfanDfRAfY0CEEeFr+uJTuPsou+Rgnw4cEqQFcKau/
8qx3Y+78LhBz4yr0rMdcQ9wjqm4kS6FpR1GnauN7wZzSWaVwuTZDey/iZnpe6Ls1xcS2w3w9XHoL
TQ8n1RdyEnSUmZzSmOePxMV7mSL/yDsvEi6Fcncm6c23WkHqR0GTnWilxBrhvEiLGm9fsc5dYH11
wSS6tNKKDJV9ET1iXiXznXuJxgtx+yFKvQbY/m7GtZVOf+1ouMNUUnK1gjVUTsgG0E4g5t8T5Fp4
wvsQdSBDuJHukieayOJyjhzInXIoWRAWioahXJS7BC59gT+z207h6EaYK+NqPBwy71OU2UdKChp7
WkOYe3xYymXJ4cc21C80ek13AuAAr68CaaL1DHbMOKdZlI+E+MgLKLFVGQ1o5t1GPh0cXgrbcoZo
kxvlLfOS4CIYlXsUNsC98tkEGTfPozZLSkespe7ntnT122PV/Tfs/85GDxBbc3sQ8KgefAT436Fe
JwYrJzwsx32DJZIYdCTnxcLK/FBB1O5jNt5cvq0vc75/O5ms1USybtx2n6GBtfgFzSYrRblqdvum
WCfI8AVVkeT9CWwg7bA/Uv+pklTfsHOLm93nXqTZyquwWpPwDu7LLSfKU1et6PjoJoanR6FHPTMM
BUpfqVyyafCWR6GHJZ22bDWassq5JInYB6a8FX15NsgSoo3NHwl3c0ICd21gZSt3TGmtwGrycDoy
oDZXSGgtHq1obqgEa8RN833pEOjk7ziMboQ3TUg0dyRPDotaYt4hEJXbempd+N4I7sqYq6Fs+dH7
lsH3Afk0AtJvm3DGOMxjRc/ht+/ApTsexQhP7uAyaJeKLbD4LIiIqJ6Pcfdw7u8HRuUaNTTeuw2G
Uyxw3XV+rnbNYp+f6P+QgkaV8mQELUT1LyTt2UYlGLeUxCDLFN8PdKGunpfNymIiVXjUW951TQAp
eG0/QIf0Z8+6r95GFpumx6f7epag5MTS1iUO+Hf+nDKhI8spSI5TqaTNdqiYbSIkB/rkmsfmqDk0
Pk7YhFkmzGegsX8a2fTJhg1XgXKfxeqNxyil3bOQD+bYy7V52pwMJdJMCyReGcP0q4Bm9E9BaWQN
g6YRn3qCiDUTd08tHA+wk5+V5TrEfgVvUdiv4p1WcqpRSWN4JEK1zLfiuS2hK+0WkXyWfdYxNQLB
dG6Y3xNEM0VpMaH6z2Ee5Vrzxgy0KXNGk4j11ooIpn6koZMo4Uj7CoaVNS7yt2+HYhS05bSUKfxe
qL0nSYDQ6Vlyj+H59kGdArISY3+nv3KW92rgGpfVBmTYpEe/lr/ITFxfcRSnQqy2+sbjl0vZQ7fy
JM3O/i8UO5PBEmfN1i7QHM1BZBMh43MHHvV0W97bFbvrZWcojgdLZ0spqJfg7zqdEXQ3XTKfYaln
4SmRifsk6+DWp9rWmSxfIY9e9w4zm5XYCGuaZ1si/zUpxYgcubN2U64iL6IjxqLn+ESlfG6GQ1iU
XOe93XYYgTDdM/XTPeDFY0sJ9dLvZSa+Tmy5qN4qRBRkCQFuxudVC7MTGkiZ2qqZMbjlxvxQrzn8
Xd92gsSclTY7CjGZaENiyYCL8El/5VVvK/Sjncvsn/DmyV7MnT3SJSu2PsB/EScqVJzixwylnAkM
qYFFxTH+QWNjAFLxVGPf/kWHneMUIrc6zqRxn5uBrc8HX7cz55TQ40/SNKulKiI/EesgNNpCmHil
7DAe8dslVi5mYHqPPDndnvC1jmUb7kPKvDdPuMMgGHlidzq4DMB04JeOKN319JunJFOYhu/ZRbGv
fFFhNaF+Mg2hvJepGvRA2ha0ycG4h4/esZ2StoWrQlf7N5Ujt14jRaQDAZDqQATSLuGspj+v22BD
C7xOxQXmJG0IKAir9Og7Pq3LrJdnlb7oedyi/W2jfOD/CaVi9OXsWdJUb78BiUUIHQZyH4NTR5yd
A+gkTz7EGsVEbcyjXj9vB4EFvPp8AVMDtpc7ju9ik10lpiIG9ANGVtGRf7R9lTfKZc12GCg2XS4i
+36qYfT98Lc5tEtyOhsICwiVLExfh/RMWJtXPHgtbb5wVnm0yiv7aRt10HUJRqKW0vujtVKMGKPg
FZBk0IkznmwkPy3uMxaNfNUoP27wz7XVrEhBN4xxVUsnoU14ktO4vCT7bIbXdyPrKVbo2qDndziw
ALfcevfseDr6G99H60wW+C2bRiVxpUpvAz3u4fY9MsfvATZqIYZ4sHV2TPE8JXseeyduIWd3xINY
J8ETAk0ot+J+vwx72zCsjxWhGaMxwFt9Ahs7lqM/vYmmrpwgoF80JO6VNRUuJ2EC8/7832cwgbzc
GvKZBIvrUyzxLL7I+Qkfm+8ODw2J9nnKiEf0ITtqOFyzgN+mtB1taTcgEhOKWyWpmPtlbBFOfjDn
/QF/r34PMfNFw2ki/d3dIXayPbi0FkGyHI/Y8+cfQO+3Uy/LOG1mk3EgZ0M3hu9QvlCesp4YUC4c
8dO0P6xBUrH4JcXZcrmec0fORRv1xREUxoq8SQv8GIe+kiYD35DGzJG/Nb2hsKNrqATNInHDw8j8
Rk+dKzHWxLS2ktqh44J1GIoKPQmK/chqQC8+7IWzIGC2vWex5CBRvN5nBEgh0ilPXSQUqeAUJDhN
rUjd9U4not2lEKXlOWwOinhhvM45xspFnjooRo+OeDFYNnkAsBGzqlG9FqVl4aw+5AgPlhB5drO2
nJPGsKai/U8lZcnv33BLKk4VqOnMEykeFVmQo1NrLHFcU89nNvltWFA3gpj+NltM6vq1FVmAcjP1
pRjPfqSLYUIcTAruj1bREG810NhkTu2wfoiaFFAEm/6mYGuyeXa6qx8vnSbv5A9wC29ggzRbiymV
l2SZcOq6zLopUBEEgD5Q8BMCNDfnV6xzQ3MdQwS20nWdeyrswYQeVYXh6A+pSeaksjqonczqIrxp
ZN624j7SFN4Et2UrHFIM0wfTXIw1EJvQoqhuMoEA9MeCEFuII1Ri2h4adNy0qRDKB+nf6uqTGP63
mQ+cj26naXfdqXHoARcb8zQi5cPxOmplGwuZI3phZF8mJwBjDLE30ReJVAl3EB/1wR9LB9YQWHjN
PKfvUxTLDtxWOIwD2IF0feqREVwNDOeQyrHL57lB1LN31KM33UBhiNPiwFHxCyPzS6PgK3RmRl0R
8uC9np/lSzvUI21qGHV0xMJkOOBUEokNsf38UHfB/1Uh5WcGKrFmwKGywS2ctXBve1zrQbYcqkXe
zclYWdCsYw5mBMGcgGwbVBVt4RJwkyFNgpShEpgjIkBwLvSMP22VlrJM4x1y+VfIyXQiEUV7CR17
N+58DUFqNY3bF5LIfLe40e/5ggWHqn689QrFqTmyB9+N/rh2VjoqJT7DyT21D9iWpFJUyYKi8sVN
lYttqYfq9Y/sW6hIRFdxqPSM07g3coyFvHP9j+CHkAsBr03aUHnQ7QhH6yCE8SbAqEKPO1PfRXgf
+9fUkQhCliXuCY6ngNnjEUvqBWJ7cFdTR9sm7/2Hd4z2fUOHkCAe0jrCatevZiW05LmQ6lP3RVkI
sNLd5HbAUhYcNYbIb9Ay5EN9Ij2Hz09fJetRYwhzYCf4SAA04s73xePOxe5okLS+RsK3COvClVhO
h76C67iHaxkfiuKhhKyNea29Ox0aWz/kJXWUOgBfZBFl17oIOVDHhpOL5pieCGiE/voJet/W/pbY
inyF1Xs68/Y+rvg9KXFN3Q1I4t7LVkIuOYTLEWr9d9uL+jlg3NPWEcc1gm7dPcSDBKE4yM3GdQsq
RlczvXKQgfDxISoJLZ9lHkYlfQ/3cbE2hR/ljXS8y35DvhEl//shQmo5f0Go7DNtGDcQuqKsbZwH
cIpeyb0jy877IzK7Ka9yTwZY4HRPCTAADLMIp90G84gfyYQd/WUZV/2rqyEeNHfp8m4NUkqlF27u
7TstjazXhQDIcQ5uzeUx7MVijGlzmjWdvLFsLzR74727pVEmrfzIdQXX/nTrooMS/O1AGhUSg7+t
ey7kQyvfkycamPG6DtCg12sLvUDLuBk/oRGfvObX7srVsdW2I/lAwW9PpStpe3JfcsqyKr16DU4I
hmsVJJFHJHPv2igbo2QWpo8McCUCX+VZg8cVZv+BnDa83DVVfjy2tLvxhFYQAfqzw160UlsYV31/
zIhp3L7/h5/KZiwjPLeQzHG15GxK6/BMV5WI7M5yGfQ3QpP8dGHbV1BOcDM+NHym9pT76lcKUkcf
m1uy2FFnLeo+djL1iitnFlP2Npf+EmkP/f0pqutdsxDmBfhzRuIUgybiDT80mV0b40Ci9f9UxaJD
WE6jLrKXWxVrro6HpzrTwpjnouw/NYXrS7HF/oFFJGE0mNZPKqnH518iXcq+i3jHhXnK4+wD4OkO
loLd4GxM5EzOol5wg1c8HEiVGGqxOoVa3ruJyI/w+zwyv9r5ygf1lJZgtyLwkoPypdkkmxCLVv5g
A2iBGP5eceV1YaxnZgzU9BvcmQQWftr+LCtY8XkclpFvfbFl9aSGUNOMP8A8nCfYcunZpeN4+H64
Fhd96ScxwRt7B45oEuIEG6QB5BcTcw2lLLGyXMmuxg5pqtkbHQ+oFDzkmByLIhhwqHPAuGGHtVRl
j2Ph5yqolXyJQpsMRBcZ56fN2c6DoHBCk7841DQHolsMpYzozk47AGT2Vf9nkd96NehepXPEHmH8
u5lQIw+1ocOOKeFjUF2u/2g5jJgc46YrQIKKmVaFByXFNT1RBslosvjgNI2EunAA5F2GMPlim7uM
OpjiSu5MhyUFSA+VX2sKDKdUTbzFBbpJotIrgGAp2X8JL4/cShd3RzKdGbE7Ub2Gi10NmLtd272i
tX/QJciM1wGDGavPe2mnfFnFkF2TPcvWhfoYOoj0QZ7s14ww9gC2xxDit6QXFSX5SQp5Wy13FSv/
zcdXl6JANQFdswwE2caxF1bZyNuqjiGpHBPmgCh0SspuB9qP3C9yEriHs+ifq6cnwhAOmi1IZOes
1QBbsWtp59wM/xVT+h0wjN3DzBRuVPeDCAcoF+fAgSf5z8yTrL84L80bzUJbCPvUscBwVgfUQj9+
OghuvBieMS3x5pGc2CNp1wmW6V4YYiAdd0o/SClkManjf7WWiqTTGK7VRjt6t3fqvrHi/TL1AC51
a/0SxgSPi73IWO4KqP9mglIcao5ll+EGSz1q5lLuKLV1SzYDdgTZ3zsx3BzvRG90oMXc59zfykK4
HCww+yZRikAuizS0uBEhVUKxNokzDHwnfGbKs4D7aX/p/b8gBcK5KebzMClc6xFLzXME3kyZzKnQ
Wk7wpegKA24Cgq5xpnn3HmFznZ5Y8W+EttWqkhWVgN4cR4MWpTLhN6tsEKt1OsiqLjp/8Qh7Nah5
vgHOAFZE48xgTjGqmCxCZ80SbxQKCZ/mGO86yGZZPQyX2I3p0pAYlq/8b3CGOZLwEUAsLPqamBGo
lBnHbxx6/1Dx/AGQpJYQBljKRHInK6lWtDgRJ45cC8ZkUCT6eYqS1oS4mvDxOiwhgs98oA9BgCNN
CccFFRh36DwC2YTttUVEoBi5+02sk2Mpp8Yg5Wqm9hCmVOD3oSPV5LycDDmo1PZDJrXIBZ3fBD60
drDZbjOyjudZ9gs9uCYtW/kQf6DUsVYUCQjS7kYkvVOMc7ZhbnSh1sdx3IgQszccfkjtxMeX62a2
4cCGazNVMSYBsZflxBXPkabJmhMozmg+Wk5ljtoUgkzh1y/1wZko+a+LwsXWfRDIac/zZ9+6FQ9k
cpszgRZdNhcOUa/DTm+aIioMUG3UWiuJf7++qJG4drb1QOYJALsk7COVJZtyPUbr+BClej19xDu4
OYafRYj1bq0ENW9PBcRzKaeMs3kfVGEeyopZvBRmYwWDfA86IvhcjE2wqfBW2/GHbtn95M0Exgmu
9m8iRfgi5GkHrX7BGzx8w29OG7E3uxmAdLiEA2xaH86RnDZ/pW1AgC7JYnW9swv6JcC3VycZs894
KCsyWv5ws7zPW1q2xtwDW8IAFThnyfm75YcAZwrkIGU3ZhwQHXZ5zH2WWGPofPUjNwg10mpFAUlm
bhjb1ATzJZ5FnJtueGgVSd5O+RLThLKoiMO+vr5L/qy8AiIsB1ICs5hdkMQ8g6clzCn5ynjlpRfm
sgkEUXrsG/9AueJdxZwugBQmmi4Soz5UGlgyBEjWwNXHQtSM+SwmsVjPUN0LmxEdz8QU5Plzopl1
e1prydWhAARtos7LE+9HyINP0Bs1bkcACEwiJ0POT5hQCrCDZJ10AEofnSD57b3+Xu7Oi3uHq6jY
k7DTwuL0+FeBBiS5CKtY+s43NVd3Iw+q6niIV1lSPFfu/3aCW368SiRjD67kyGj3lm+g1R/vwG03
dY9NkPYYbykxYGCOyVH/WXz7+oh/5QBb6FMcQB0DnKAaUAQZ29npEIS8hQlGm7Fuz3fpCWCUIKsG
7u0xcRQTelBtassQVvRu9AUesvtiVGtEA2F50GTb6pyWrAB1CoFzaHWthROfhlYosuJ2zcROI2m7
CirbtyiWNOIHnlfEegrj0PLJfeABNe+1+71cnpZFjFTViVMKj+SKcKdgoyNYTitsfGZGlNO/GJes
S945xg1YGNkdPf4I9n9CDGxTIf06inN12z/UPQT7cmzRvIhJlKMzXT7sTolpygOf/yspDVpGcKwC
6a+qg4p/Q7x0mWAZtKg0wbktr/8m7foLUML0cb94foLjeetFIxmS/tk0kiRx4KRh5wOyWAhRu0VN
N18dB9hW4WsnvvEnVS3v/3K7tjejox2hv/cvYMcNyNIesciqZUOjhaHaFrAuQ+UnjXQfraeWJqz/
0ySjZ20o/QIYvZnQOXrRjB1lxPN7c12zUuTxQhlbCifjI2EikMN396wZJK0oRtcjLYuqQOvRzX4T
rt7txH0Ovc5+UxPD557yCBL/0TXNu2GRvd32vCwTQHU2LwlG7eIlWebhUpCQ3f+/cvDssW7rSqUG
ZBAQtHI3TE2+eLao1dE543H3rmAOeoTxfgwCcLdn0IR1iBHo9Ud/l/epy/88uVlcBpeJPpDidV7g
THFE5NW3xJ3IfYYT/aaG4u5r3LQnNJj2O1dMozAEDmkkYEvvwrTQ8o4Rkj8y8dGOne7Cv+KV2dO2
UMVv2Cf3Y0JcDdpsZCB87O2O5fnaY13OnZ0OxcD3NZPSCTFVcyr2UN6+ekb9dN9q1gycDwInkOHQ
hFjhtMRrUcdjCaHSvovAT+mchbdo1buWU3H8ki2EhvJvLI/4GeE0bEBg7GjJOs8KsEcH+D++Ci3c
8dI9Vhi8HFTm1asNTPBocK9U4YQ+69eQGalElxGv7+/zv2PWWkQkaZcUaWb8dxj3V3lZ2uJa6L+4
xTUD4QRvPVVc81UKCufC/1PyMfqE1UwNbGmRp0/y0SFe1gg3M8nfoMEaMUAlEjvU/pqBUiXyk+h0
qaY9+H6X+mSSeqQivh4Ed9TvmgEKCQUWaS0Q9X5NhRtXeTuxKqn3mPJAdRNCgoJICD0b3xL+FQ62
uOqB09M0fUTSvo9ktgQN0hhKqGmhMXbf6advRd8uRWGcyOTk1NOovDvYVH0A9vqONIGh2CGXwWTm
RJOmdbIWV97oAghtekDOm86DnidJCKujYx9RhZm2vBIKoVrFXePBCeL/2GAiC+p9jZ1ztby0jt9S
0/Bq8VH0ICAw0lSrTHrhhzX6pJj9UVxO/INFejHn2Kb6iPNqXBOysxCK/gY0c/3Td99pNp7GyDGE
3ZtMfCHkc21qxjAxH1lXQEJSshRTE1ipeSjw684PgFcHTfitZG+o3U9icflca8mOLR+HUiE6xpYD
5SE3xA2/L/nFad/ctwRc3T553JBe6/8K1Als2QH2AxCyy/PSaLgMp+C3vpA1B6sCYmkd1EPQBrdY
NmVwpOn4PdOrWDA0XcGp5d9oiWagSJUzwyaL/PhUKP6FnWwGF+64oXFQivmFebUsXGJ8S6M8y/RI
HLy1wkFDOcOKpU0DH8Okv+yKB+JifVR4QBLreYaWim2UAJkPeDisGhRwemWat8xlnyMCrVFB+6BY
q5BZ2Sju7RMgRMB+M2RkjZyAK4BXIm8LfixKCmHyvg+qBqe4GQH4HdKCqXMx9wEupnSXNWC9l6nT
LpTFlQ0XfahjkQ4V3qd8G2v6e9aCsh1lbR+Oq6/sRFw4GKcsgVcSCwQjDZ4epYYs6y6BAVIrgHuF
aH/LXK04LwJTmzocSj56Nzce2JB6568Cy/3uRsEXW0qy9pOOvbEckzlWfsGhkk9M2wNBsXllKI5o
0ZJOPPs3BT1mNAZT1PSyWFb/gDupEgT35DKjFsBfE/N2OptYWEHQjP+dHNNKNORAmIsyZmNQ0AqI
OFkAqvxH8GKZI872cEddtDyNVpAvVMXsiXUQxDPQyjOSnXd3QZHRQiPkbzNMxRzGS9SLYB8K7QOR
rnSO3iT+2t4Tne1MIuoY7FEH6ToYpVcTenUtIU9n3paAPP06leol+IZoJvf2CUTw9VNGZYjxjw9i
yrLXKkt8tSwmC5n7mHqpNG8DMQkdhBr3EuStFqr1P+GWTJvrLl3e40YP8CRmqqFeFFXrXW+b5UqL
hZfz9Ef1hEko4sXgcYcUc8dLniQ3YObCShEC0inYVfBtCb9FY1GzLW53rD4Z82pmk5u8xH9kSixw
JfVB9dabgu4cSsoGBQn3eVqJl4BfUDU1GTYvw4vZJCKaWTLAAsW+n0y9Kv6D4MwwRforl8RHsjdH
sd8wPWBrvFa6lg3JAx6TB1mIDD6dyxFW+Irr+AOmnL51AYwYSvJVV0mJz+vo+pxmPOVZW6ZsvPcr
Dd3qMHy632p1sptVovAAxHbWs25nwnq8Y8VWqT5LyzI8oc0fpEysAtPtn63iwmPMum/TEdXw3hlh
b3p3YGq71Z/mlN+ozhNLTz4D1ww+540lV+PLvBtFsA4uqDvlLbzAOJwNkgmPpcOtuhH12yetH1wh
kat5r/WCvReBz33T6h36N09KTtXCXb8uD9SXmovdQe+TxM4NKhqcrNzTVyKTib5rH6PImLtlwQuH
IGnExEICBX43MnF9l5lYWjTFNRZYqsnqj5vddonu9JsTbPR2iee/TGixnepwXxEwWI1jPGuzK4tP
Up73+8cWsrWa0kpAXTNLEFOVRtuA+jF0/CsnhyKcTMdG+VTBEEXw0Yv/fYbkal287pLgUJLp1oiM
CdhyJG2y8Ox6Yh4mzY7onSg1k/Vva1vUJKwnVuVWGU4gKRMsFNs4hLvE8Xg8hchNtDaalt0XhoDK
XPddlDaum9bsrfMGVTLI5Ymat7E7YyZPkx/U00xoyyz5cwAGG8nbiaC4o6/e0Hj0qkfHgffoqnfM
5HILdd3o9UR7vY+pRHHOXbBwT+K03Z0b77C+bt5JMCJttbj6astImph+1WW5D7bZLCvgE8PKgIYf
impojIUsBowb1bUIJo48wwcp/j2cggGn1MBSvr6MGBkAiDKA3Rx8jg7OIPKpZvEfO1pyiAlS61RB
03WWKfNLZw4Gkt3o3l38QmDGaPRBX9sPf0m34ygrMeEWtHqrLdB20qUK5aPeAxwstzb2wtSBihku
QXhJOCwfRVb774aryz8NPUlsNdDm5N1KIzd1o199yu7xPxdUoJBdNcNDLNkg5WVSZ79vqKpujYnz
AQOKf+TweaBAnR43gxyB5Cj/6DomF9pkF8kAsFk7rIddXtBnSfFag0WTcyzaBHC94b9SnuIBRNKV
a2BpKjF9HzERqSNhsu+5sbqNwCIGpHaQJl1wRlzaq1r95jAcpo2XdYfhDNOcjhXNd+OUHHwGbN7s
9J0ex27/dqJmUx4EJGVtXrfgVuUevJQXa3FmolAGPW0aPDEKc3v7T+YLgIUAU9lRKjT2Mq4400SY
Ag8PCJP87duOTLzJonrCuhd0Fp0T4qqXrjT9tmnPpct/wvB/tf1SkCd3x/iPKBb07p8gRzV885fP
2hzv0uhmEedfoesDmHCrmNwY/iOW56EAwqWdHSO0/A2XG+wDKRFB7Ggf1JLPKwooYMerH//Q+l4D
duTH9U6GGBkEDpnDIZOHvHHuk9+/kxStWXUkyBQhF7LtrklBx4xs/woRtylyWw1WzI7neV470idM
d4yknNPcEeuthaMT5WDTSOpF3UDb/nD4Q95Vmx5wmthvFDWRV6IHlm8hc+BHzGLi51VOBCP5XLrd
UViLbR14nX6Ih1vLgw3F6UQMZE9Ns5UeXoi5ESZ7f6dDKUBtv8OUtc8/ObE89t4XeKj5aBbBRDkE
AHcqLRWjRjsxvW4zhb5TqvDC1MrwcPBmmOQREA+SVGBkRxPNIelYKhVYrlkoVWmUFIWvupzYPR2H
z4nNKom6M2oWH7dKC8jqX/3Vzk3GFhzU2zb4hTWuMLllzAUhtL2aBWGPkZWmeooUGEdh5zt6/HrZ
+4lzwGLg0xCsVdMGvh0p4tscro4TGmXWpw2WipEUjosU1RcRVf0z7tYQowFUTr4Eku448vIoCNKM
NvcZVTzyCL5sJAjj19r+ZQFUcnq53/T3HcAmkZFvY54Gduz3IEGGhAcRYhk6L+8TFXuMBsj1eCrE
NwMXSM1EcUzDopn4rboTKRgw2dURVAcIsCN0D/otwOyr1Y80N5pudnBKvreOcFtXQ8mV5pVTM+Ly
tE55szeU0zCvMnqfefqb8KQGV+xlLx2kFBwkSLTzUeRFafUFKY0cS10Vb4ZLvNK38esvJs3lcyT8
2LZvegjD119jts0nV2495uEX4l4GI61FDOAM74++N2ip77/hyikGQ/VQjaYeTbuGLQlQz0GhBiGe
FzwhDWhPPZF5wNwdyUBi1WkYAB+ZNuRZYZBYokMyzYUlr0Rb7/qRPAo+3md5iRDvvonMWx8wBm7E
G1Nz+9rzNSwGHNkeVdCoN8S5M/vzybv8H9PUlf6J8QYgg+nv7lj7QVp8TbwpgIeCp+BXPbxqJFpY
kL4BJRSAYwjVNAGmB4A+TJtzl3mC3t4XF/0XtOLM5StlF1hrPfppGRhlTAQQuYCMlZXwME3tUswO
ryiC+Ml2zqHvFHKO5xnELOHaPY6dw0Yr5y3AX/HVgynWbJvC6QIxymOm/YgB9BGjwwuIHZdgEWMo
5Z3N5ggzZ+8b80Kq3lmZm4kyrY4MluiLS7cG3fkU2Ma3LJXIwyBJEsBjJCxvY+YlQjoHkY6UMoJ0
QUGSoubikw8SyGFWY87X9EPQeJVoaAkuLBw8o6MLCAVeK1f4iDKH+z+kwnuMMTvOzNcm/FDoY/k0
QWKkDQWQl0HgGQdF5c0dyRT6IaTwbx6I73tNkQR3M7Y6SfnmPChUIrFC3drAc6VuAyLKx/Rp/1Na
DzHuhST6xElFIRwiR/ryxVx/657frX2teEppK9nWXkUZgaGsIz0tnIUUwkItYFTgmGJrGKOu1aYQ
un1Csd/FHfpKi0mn4nSRyFichsio4jv+8FN63CKI54RzGCxnjljijYWlPZ2De46FJQuZYvFDTX+e
pY2MuDC1PK4+lmU7hejBHzXi6CLcmP/QZar2w06LzWT72JohtEJuOZdqRiZjCRFKswRnMZoFUZ9N
O4mzwuVDqaJiujTHrvyY8aewufHjyyZas28e5Q8uq7J3UIxJS8k4piHQh3AflQl2hNio6Ro2WSJA
/cYV4/dtWa1Z9liVwv0bUszwRvffvkciX2UrTr0VpI/owJCaGhFjrIGFXl4VC/ohv0voqV2mUhnt
inH/o+jFffJomZmJS0A9pBot0o84p41kiNvg1VVsFB8OKyQ4+nziM2sRL8Z+VYU0Sd1RWJkZ+L34
GM+E1KUTJjAItZMAEkVR0JYTrZx5k+gBtrYfpmjOc3A+fEeFktzH3fud6ys8GSP0+5bQ+JE9zwkG
/s+EzkRgKyr1/rAQAB6AsXoyxR13PxWaznq0G41O+QBrbu3IEHQ4oTysBXLNcPJ3cs1CRawoprjp
NXC73UV5cQPq/7pq1UjO8mEgZcbGJnNv+OAFPey+6leks1zBKkHCA1NnV8I0FWQFxN6HuiXPxzij
D/ZMTp41luU2jy/Q2fayeNPd81U2XuBlU+lmQGgvFFdtQVcOveha1lo9ajlfmWrX+FZxT1GL5O6X
J7yjfJxv8fKLPGXMKxSULqDOTypmxi/Eq7Jl+1cLgatK2KgU6Y6eaZLpR43SIUkzDqExnmRs0o/W
yzWUWT4Fi7q5yEqp1kORRnrVXWog61iS7EAScctlDqBr2k7ANjznjWh7YhI7uoTUP3IHFUsJ6IZc
jlga+RSSSi9isDNEkycT3mUxP6aHi8ZvEW8MC7eZAfx0+RhmwHPrd4SvlwUJjUphGgmIerEq5ckj
5xEpc/yps/kViQ4IokYwwcOy133RnZhceQWow2dNE3jRfV9XJZHc5H8gG3T0eOmbcAQJMzm5uwgq
BvL5eAcZsKtlxoECyZzuzuIlbwDapn/j6XaMT3X73ySoQ1zgeGeIuaOcvKf+Vo/VDxTxb/YIVcCz
H12j4snTzfcpzaKmiqGdZafu+F1uGe1K//WGW2dvA9JN6n0OfmOnk7pYaqhukFXDFpgZMMzY9ovY
QVQTWWvBa+1P4vOd5WmRgqzBqkAjZKHOkvo9HXgnVEsTNhkD8f8afkVP08hRyL0QV2IjXQQ6WEUD
GEUNqGiIqQItooG/so+sJKRkm6gIYP8Ekxm2fnWXkcGKKcsyKV0vpLr7xstiKnY0na2ZO7w1xLWe
zNMRMZz0/ZJSRd6pN7JbJxRNCiqMlcF7Ts5NnNxHz4x/IILX6ROigq9t3VWHkmk+yrFVNmlR83r0
z042fI3FT4P9i12Usw/LclfsOgMT9ma/Qdk20AJW7KQ3U2vGQ/ix23ud1tKyUkXNgQm7kAfUuIx9
qjyk+1K82EyCc/tZtCVBYiritC9hxqP4x235atA5M/je9nmdwRgbTN2ma8FOUzgsZRUHbMrCoKlj
lBTvxttjl4gpNzpIS81TUFPjsogtLU18bDwaHwsgpiaYKYh5GlC7Cp9F4/M5V0XsIk4wq22Q0gvq
7UOqqCuNOLyE+gzZ4y61A5W/jeJMNXzxvRwRKTqMhs1odqbLBdlWQMKsGWCPG3GsFWCH2IRuBamW
13sBEKUvOZFWQO5FN/BG39N628OGxli/m8q3CqrQiQ2AtG7MhJSoaEu3IIunzgYEzWFDWoiciaB3
H9BzUOUbQrFyoVUWmppQmKby5JB8/AnaJcLPWCnmpeW12FeCDg1pt2eBQdJETy9iyBaUE9py+L4D
ObX8sNbl+MlvVEiZivWGCTnpQIlaJtrqWN+5QnqdphTimfzylwhTDtwyUIMku0PT/3CgKwVHSqCU
/YpmyNyoSi09xt/K5NeMXg0OV+c2VJ4ezUCp6xvpn3XkQarvIU+X7+Rgjqf1DG88AGYrM2rS4Na6
X04T1aKmZOCW2tmlNz/LXpkockd3x9bVTm+M0taguMjYOm10n2Nw2fCORKuDcckHXOfy1CTCP+67
HCLPOJo6XMsxBW0bnEnRRUH+c+6Y7X7g0V/7UPshXqmESHL5pVp5v5PxqZSzo90AGyP1S+Artpp/
C+lHC2fv8BSY/yZY5gtK0G/9R8CUQsPa49ZDK/4jLnhfRMewdiyOcekI5U1w6M+qlq9lnhfzl+Q3
X6n6qiTI2prcLnmi8HV+Im/R8Rqn3AXzs8H4DEbUmoPsGaBTy/8geAWkoqjnzQ0pQurZNNqTrHAK
VAv+X16vWamOZDgQgP4SbPwD1D7T+WvN+r9uz8KI2U32oZ38oCITicaZvPSHWd5HZQlQNvjHuYT2
ja/ING3GicIHTvRaZSc7hwX7DUdGKmAX3F+H+s+54vr4zYrtQOfwCF6BiJikm7MYdv2+Ejx3baTI
3RaV10e0V6fLSJo1flvgLDagxGHMHbd1n/LiLruHvjjLai7Xd7uULxHDXetm9vKr+1G/1I4Z9Cfx
Trh8dDAYnAo0B3umMFLq3DV3qJwAhLUAdv4E07R5ksVgwzV4P+LvWoqU9LU+9zBnNpGkaaOpbAZg
JWVR1vJApeX/iV7aXmkpjZ3+6FWQ1L33ilFIE4LgF0Hupc1Zb7FXzkDgpohUP5fSdqahYk+WmmI3
bwwE40o0lcBpmmFJuoFRd1sHDf8btRkZaJUAXsjnMHHrzmEv0af8Nl+sgK+cgSJRTGHBbRF6U+Wv
ne4BplNO6mwl6XijSXqy8GS+qmO6trvYSc8ePilEmN9qvNt0ylxdb8pOcxxlYOU+Oscv/KJ+nKTY
Ciy67IpuB9VQJ2J+Cb9zplfboeh6u728LsAyvq6+OHzSt6tEN6N5GhTlx3BY21L/bOrosfCq01hX
2+poDah21qBZ8WJp5/nZGaO8feEeWsFoNPNe1y4kGYZb2ee1rNKYFoo33tCEgOSTo5BAdkgBZlaj
nvjcI2xWNoWjV5RRk3CZdxGdfJKkIiFy44A/QACJKWydSuruZ24/cRyFu3IeGClUGRJxUQBn7gcb
hh84t9rqHX7S86rulgkKQebKPIUseolg5ziH2qelwo/lobo7lAjwwVeVE4haZYE+l4ZWxrzkc7Se
t2paULb1jt5eG/i8Jw0uIWMahspXz/6iqyOCl2nol+h/LGxax/XxnpysppVONjm+UPlXIDnZhmXC
TqMfc2DN1kazdRn84WueGlBemfO+Ze6AX199uJgkEbIVKfB0YgosJq90DSxc/sHbG2ISanMN0zWe
u7sFbXfBXtc9es1kBSaJUpmjJ2A63j0wgSPfBcQuGXlP37a4fzx4uEE/DkXLGdEyN3iqTULgnQrG
bMnYjy5865BdN8sZlrouBmZAjufJDod346AwpwyoQ1S4hd0fi64gU1nY4KElrjxpU3bFljRUa/Fb
CkDkv6DrLRufekokfE+kDP5AvG1bF5m3ReAX+3OEgsUI4RPDbuqcmIU2lsIULN8lwUrIkeX1pyby
pn4fxNfs555K+m0yfK/gqpuJEUQfomi4nFS2QQS4RaaPehXLYMofgHVDBZ5XvalEPib6yft3fih/
iQ+obX6OJP6rqJ6/9WZ/usq6iZR2RIYBECf9mge59AZYdxc/EGf00xa0kYJwzifmOQaLA7YsmCpB
i/97WyfDYLNkw2u27mlQV7gnrDyYzLGYKiir3QkwSsCiKowzKJ1eFy4nHApPtPBwfPSnyIXVjM5L
tCegSLAIaC1GUlFeyPgY3tdgw9fy/TcVB5FIrqt9c13tdjmx8hjcVn3JwApU9ckCCPaW/MV7x9kk
Nl5VAv9CmE4XpjSOVl3V3qZde1UbJQZKUh6XnDHRNK3nbzGgvFML3tuZBPzX3A2WrfeA9wrMTc1Q
rG1GxaXCX5Q3X0dyQfuWofxxDb2uSg6AywgkWCxen5xLp3RHw+vB+FlFfY9X9+lfnL6IGV17W9qr
aU+GFH3CSBeW9i5ETV/FZMakIEi46DvQW7yTnwg0MKe06a+V9SWPvQ5Iu3HGIG55DxSXmXQ1pS1G
LHMTDkZxxAzPQm4erXLiL+QSKVIL5A5RXmPa1tjfHEQNB/BmxtWqoIkyWEAh94F/adDRejoKu2gX
lVEBs2Ca/jmj30dLSvkp6wwuPsdzjzr9c1z9NoYytPCX9mJCw8H5LkiLU5bys0qzTUGPcPljVgjN
PYI7fNfxCycALXOwz8JK0egXL9j6JKYzpNR68ZHYbXO1ssezkvg1+gb7TNHNm7v7KzceInBB+yxj
iXOXVj01JWBj4vmmIpC4hy9n0NXnklH/KktPUZWpOaDS1olXbrcGXuxuOuzppyOUiObTeUNpmctw
h5pW/Emr4moplsWAEQYASHF6vuO9hkCwoZxhc6J612M2+sSqL0BWeD4b9ir4toCw/X6vMEyiinOM
wMCaSCPm6a+8NvsR9tZB6FDtK8QaXSsoesUCqSx8AKn2c0Aj5dt345qPAbyKJ/B2nPXJafAML8rw
S8qmlaQ6UpY24B5Fd1GqC3cbM08XHQKQ0CAP+lwvn+mDDQwTkBRevXb0uQVUuqei4YdnFiNV9I/3
wYwaV2kiqrl7k4mdL7JWDQAzz7HAtedb9DRYKc4YdzpX7urwe5MR6UNpdt9JbwJc6/g8U5sRl6E1
oV9bosnf04ehzGIrK7lpT569bNLkfYKpLeem8oZhP9q3RPxaetyngkTwLvUQaPF+SEraLzFIyTRq
GrpmXk4qhBwdFE6eV7Id0fjp6sMDpD7OscOrRFdq5aV0fIJakBLBuSGkRahf3Nb6bUunW+OnXzOf
wtYvZgfjoY+lqsxfFRa0Y098XMvhpM+Xh8u2ztTGf2KKKjTDiwk7N0+1dKLk+6SGXPDuym5MVGGt
lymMX7mWeXiw1WXsyVbhSExKK89a/WVjk7+4hScfeVz6LTY3rMrRtzwSS22/GR2cx75mC9/GS8rF
yxIYKwMmoj1KW2og1hrB6PTZCTiTIsSGrlO299kRosVIbXWEF0ngPbA537JW+vemggjJOF9dTXrT
mlJnnVhNOu1lZFT/C9gBT5Pe9qrtD1Csozh+iBxeHBZpJN58nL9cioJPJQjOCSkRcesAGEDo3jH3
eIgT/RgHNwe0xJ2i23xJaCEoZ34LNsp6AW54cJo1SHOonLk8jT/fl/rBS3AA9V6G+o9RqzojBZFk
n9Di8EdZUHQSsMAJeTccR79Xs6N3VDxI5grL57d9esUIfAh9on4e1ys90jEVravWj9Xbp9aQePyc
ZxwELTuImAxrvdPATGLHQo0XL27FSnZ62v+sUs/le08hdmtXBNeal6vnqA9oTkX7kjr8CH/fDxvX
CDtrNQ4JK6OdIQQpKuBb3y3flHkGZsu41SuB3VCeRtZ5ERrS05SfBeixlnddg75VLWDROqW4ni6H
SbjI45vbwXs1dbqE7nJxUzUE8MUMefHPqFiYpDvLUvwQuvOCGEMCudbKMqN3DlZTq1Lk5fw8ijp+
N3WyvFUU6ma4AkvXmDgxEkmMkbySsqUSZBHKm+qT8CRRtRRHGJt2Wp8ajBxyuJaUVFqUmz9TMPCP
9sztWlFltQeESgGNZB/+SQvrhbDeAVKKxY9Vzq38TFUj/PJjmpuDdGQxsiB49enY3S+jf4ZKY6Jl
sP+d4rc6q9q/wXNVDK/dN2dF44Y71FdtRwpxsuXO3kQFNWFat6kGxL3xzIpq8M7M0IKiGAFXHhr+
Lr456g89rVdysIbVfRJ+nu1YdkdQ2/Fse99w830agnjv1xCPXzwwTab82MB8e1+/ILsKoDYbQBg0
KeSh17QCHNcurceMU2llG3oTKZE1cBKXFEz6DiMJS0vuHYdDIYhua7NhUzhxpmJ0/37xs6Ml4mjT
mpseJz/uQuIdLylCMPyZvxgH8hmWpwa4d1BnEgI6mx35XfC2BJih2oTk+r44+3r6Fbrv5iDg+9hL
r/jo+JTGYiQuY7yGUkSaBKXOAuFEcI3m31l4jfYnyQrRSo4cy7k7P1YtZPmA4Q9pi4Tnm/I2Z3br
c4t0YIrAkhXFBsk6OgZ3XnYkJvlXIY2qNfesb2rk1697gmo91CFsPBMbgpoQtSQwnNoM9a1/hcW+
v82rCr6JT1DaIfs2QT53T106beQuLxUQPMNqExdpQSpHjv5hP1NdKhDLvL6I2B4QIc6yJCI5nJS8
eKPbJ4Hhbl7kTZAkGv2UjUSGLez7jrL7Bb59CnYwJNc4b3p5/7UL/CqDFDEkFPSoDceT9pRySmuL
HZ8esIs3lxxTno54wsvhPQl77sJ8lrW/cejcLQflcVl8MCVydclJTBnlR7tTqK0osDrDD9mlikus
KUn8AhBJKarCJBGWoOZvq6yn8Ajetf49yBJyaI6oIVQ/pGKHqiyxcCETIBEfslOp9eoCojncRSBX
k72S2bfJ9x6ObqxDiJkv0R0KoBvUGoYmurrE7AChvsFBnIICk+gcoOhK6+aUfQd1aeVTcpgGIFlP
IrIcMh+Zsg2zOR7dF8KAwnq87sL0u5sqie0KQnROY7mmw2cbjcD547TqlmQ4OgCwvVdyEtJFF5vh
eSCfx3cYmeLvBwNCPz8v9hQza5M1j7dNyBP9EoTf7iZBNAvgYqFvNMOSvau1Z3I4YsLgJcIDtxB6
sw4lo3Y6UzG/ksUg2xUf2OBaC2/xBbW+8hkGzd/k3OhghyS+6045wM0mSuzFn7j4O2f6O1CS8sBl
EhBbKJZtPgXqfmSlucPPEx3RPKXEr6gd//fOYyfcKnI4jnGlHC+0JJUZZ44yLwoQJ+kladCXNM4D
kkflkJE8U3o1z3HalUyeKjPa5B27oD+fNjIVnlFWlYIxVL94DhjMeeZZ5EL2UKXDv2mokde2Q1As
jCkqG36mH6qCb26HHrcZYesw0MPCqwpMaestx/Xtq4Fg9EXnE6QbPJme+rdlPoY31dNNppGCzA0N
h98D9OtWIS3MiKaOSdpOq7BhYrzvw4X+zVKjAWYyvrnsvG9Tv8n2UhXy+9f5uKs76MaKsev0TZvp
rdOs0AVmnj8z2SJjVlqN+0m61m9sb1hyhEH/X+lApf+sHYFwU9Zg0fFBKDNUkQpj8YVDXePeRcg4
Yrzk8xsW0L2XdT4XgGlwTnCv80nUOsidL7svQiyryiJsP0elWBb1dT/3nRzVnzgvYmDLtgpgEes1
l3UIIYl/BCVlA8jHJpClXDhI2mw/kkmozL1dALIA2ynWweea5RHzrOxhGJ3HBY1CV79E9MmbWa2z
EgaMK1D3V2rWYVP15kNnZNvCDlIlPteeLSskyVad4Lac9O9QkDZGnGlB4L5ig1XN5G+rgg3qBYT0
iApxG8cVV2zPrp0PoHK0XVD2YINAczhztxblj26bRVqcXRUWqVNoKbt6x9iC2yk8Si4LGF4W5iYA
QPHwp2BFCXdOc2E8l4r1kCajsXzHnMIZB5iHRifdYgbxPlU7rkgiBmFyrCjfgslD7HYvvFjHcoOH
QPcQ1saPTdXOjTJzlNH9Q5sAKmzTYuRs8yBGGy6DWKCFqnY+ldEs1ovKJimPxmTjbIGdjpnWrRoW
ncP14Fbs831AIaCOemsFMArdJnEp1roOCyvEO3neTQATvudXGMwbgjR1v1cqglvlh6OKAyR/rmcZ
FCJeq4nSsmmH8o+80yiLmj6/hV63UUVOyJwOnfAEENwqQ8fjk3Ly00QuDCRKHhJJI1rVoCWw/UaH
uj35o6/KuPqYisfYY53E0mkuvF2BKn6Rbxif2Qznzf9/eeVLJr2q3LbdDbnlX6QlA8Vx7gnvISWu
mrUxgKMwO5j5mS9LQ3r5Mw6uEIsawtSMba/S46j8glQhQWFYDn/dseR/h1W1RqcS5Jxz1XT7Wk41
Z4+Y72k5XWgzmDeoajXrUzI6OOmlJkdOfmjnVTTsoloiJAO0vIkVJ2e1+yQoFKEIZqv22Y0YLs4D
qxf+xPSYY4MSq2XGg4Efqm5h4mD3e5I8fY94kry8QaFj28LMFal+Q8w4Z0GHub0+jKw+bPF9tqNt
7RdX51XM0A6mSxvDe6pKQ6nFFaUg8fIPBrkHGebtWmlk0ima+EbMFg+mfMkV1vVRcyyx9rUBDAox
UfmNiG80Qnco13+GqyDkNDIuQVsh4oQvXJHDN3wtjI1WNcmFEttmMhL48E9qZcghGwSUqAQ7UPJv
gEF2b5jT7IDrxByw/yNM9p+Bm6zvRG0qmH440saWC2EOqt2T8gMasdtHswKmUNwJVZB0wWmKpIdr
tBT3WmjeUR3y/x7xpUDIM3yC3ZQnk72yK4/K/qUdAuumXtZz7nV8ILT58oevGwsP2v8AeFTwfXQ/
03PFXJ+WpgeDNlnpKHDD+og/rclryJvMvOOnGDPfHsYxFjFXFTU9sFLxomtwWoz7fssgBEaQL8N8
dTvqC3E4OqY5fqFaH3htnx6/E6iWPq9LjYhgt/SBr8TVDofbAqA0BZWdFuTcLNZXnBSvEj/7JpGO
DcnOfinNFARz4xfiUyMEQV/Ci/ItYrOlEYMkSHbIPNKTg2Y/Pz7gMyzDpSEeKPCbZ+RQUJtaDg5K
GI1xWdrmhOamzH/ypzWYlFCecxkRoY7vbIs41iimB54mCQFLbs6ihIAutHiss93ylqvpnW2tri/W
nvryAdJ16xLr9fzqfZh9vZIhbM6p1YFpLqUsPB+ivh48boNlH8G30CipJiLcLhnkgpDXPJ5BxtxM
r8iEujvLOAK+WEow+dN0uIhySQZ11png0e7Fw1EbBL3gAFfQLr4lVck/VQoNwS8LuR3fjcqDI3LX
UJI5UJfQETuJioXR+zh2/OPfb0eeztJ78y+AI7dQ9RfRRN9n+DZ+A6nyBHgvndkGfMvNINux90JD
3rvefhOISZ7KXwAIX/wfnCX+oKtE0XQrqS1kghkGgeB7V3Xu6+N3COf2BFJolG/V5JwofxuNWemx
vnehzpStP4tSPAQ7Wa8hxKPMD6JOWp2j4kwni9zIEosn6XYMir6//zSG+U9QqQ3vCuV8tPpX2+pH
EWy39+zHGm+FbpHyWv/4dwm3P5qra4m9UWZQpQ7zfZQwwuXvpTuVYd1pVKN0nY47hGmgK2iirexK
b5Ci/afapABt6pX3lXNQ8QOScaBqHIuARIEIsKOu/p1Gkuv485dZ1idE4QZ/pHtc0H1qLZ027OL2
QiZRUMEGiJdXm17OVT54XKAjyZibnoAl30wbxmBbIQdUi6w6zIdoeJwRQjckJXHeL5daezYzv+Oi
y6EKkHAcB+K5q4D/5ghSjBfEaqSgqKyGDkHlejZCTvktN5ozqwY/d1pKkmwdMqLQhsvCU+0OXo2r
WRpz3CPHwttGiOiYVR0CL38fgaonHeli0CXVWm5VDzbl7lOAqxFM4jhOP++yUAh9aPWQR2LfOJiL
XxVRjd1ZJEJforQh7hYx6NZHc9tlfhpLZCMkuO7Vs4qi5zjqasDt2WcVaDG/2MKJVceWcnqk4dPj
/xEbs6BTNvdZ+jHds30py4DOv7P1ndNWfeBsnvm7l8TVo5tPFE+TZFk3OzVlzbTmCtqKkswkwe1Y
KN3uY4KCBNqoP0VKNrugTKsQX1dDibkHHE556+zk4HcnrRMNOyL+h+jw/0UGHuO3W4+aC2b/yKd0
6+rzTAl9om6GNCBHqz7z378sAnfohzlGKDBhLUeMfVlOzOt2yMVkGlJIEvI06EtsC8nlbByecmQn
KdT9b+h1UOixcLuDMlapcHTcevfaW+OxUhF4pgIbplS6jR/k4xVBZL+avE69z605Id0EDqEziv0X
tgWOur3+ULZL8sbj8LV1uZIt4gXoS8km1amIkU9rWfCbEkqeC1w3Yf9ujHgQoCumFGHGOxU6y32g
c7EGsLw48l13cllxne4AC74JwcpLi1zP3Q91ML1cuqsjKOBR9MJM86pWmVSBkERd+KYcHjbD0CZl
MnBs3myelBLeccBQopVpo8IorHlWbjka4U0Wjne4MdqLoIwvPhAdC65Bbr3H220LUBDg8s5LDIWh
CEBZ4Gk8cJ4jlOJlkoCHmDXWaf6+vOgvc2+TusnMUzLUEndvLBfoJBcKmd2y8QNuqg/RKUKuLCZ6
DOaGfz56vf/ODN7K+7Wy4U8XQfVt6alSDYol6ujzqABPdqvdRr2bX13nCPIqlblLxW93GZb+hjfA
R0jz2mRbVtiRvXDcDNeghL8FrYIc04ybE76Ed52fmYtnfUnUDHcPdQ3hhQkfOw8AZGyhAqNh4stb
Akn89/bjXLsk3hg1c9ptVbi3330VayuWQ9QTEn3S3AflOOAhHvc/vNi/QRiL0weO44JSU8JLkLPm
ULf1xC8S7ZOI5YLT3ZNhDO+QbOvPPX2IXh7Yn5x5DJJs+4dPlFl0PYezEjmpV5ZwQ7inacHro2lc
y/QTTeOk17XkH02TEO+6INiTsjAEjiajrhRLCYaD99J0ovMtM4flTX8HFwxK0sq2BBaCL2YAMnly
o3jXtvYWu3r/VRAHTakwWV6Fx+mZQNm7DCSp7W6E3MjFDVxLiziFdem8NnjNA7/a/mPNHtHX5WOc
ciH2ndOb2gaON8L5AD4fQXygO568QGBd4UeeapGO194F4CSTPD+Xn954y5V2Gs9VY+FcrpYwqS8C
GJhIZl6IQpD5KE+pNEr+8OYfdUrpz0F5dCuB/36nKRBSpSMYHsuouzi6YN2GtNJCP5cSue/M+yI8
+RxbjacIAxe08h6UXUzk1YP98DBXGx+qBjO7rOXnmC377yE4aW1aeW1P+igwAfS8wZVhT4dclh2H
s0yOqdG7WVXw66R4V8lsyCk2LRJS3QRw6YvnyeVIjOPG9iI8Cw1erHxtt638EXRRhhXA28pepGVc
JR8PUHPQ1lItrruhvW3SPHQK0E1sxduX5KazZl6UKsEHN7KgiUt8GzFvq56fXd8IAPdtsDa7uClP
IyXzpdR6QUNfMjTu9tp0h9hhz8wU/o/9Bs5LpuHfXn+qMs6qIdhlcuYP3VdwlqRHGYS07mVEdHxn
qE3NOn2r43twok7tXnVAC3557nvetEgBLlInJd41PWIOrw347jsBEhjbA+BB/ShQqvdz9fMiYKnL
b+UP5p2Pd9YWT6D5kM/tIFsqguyE4G3uZB0s+XibmgsGNE++Pxed1EdWQQEod+hVCdSr9PCd4yNt
OlAacwkZuiWiwn8zkUefNXE5d8OSRzXxdKYQVaEgtvLrT+5eDvT5mEykwxNhFXRDeRacoi84G6Mk
jOyVuR5xpFKeZXX8csiK3L2y54eoCaFwYv/fn9DQ0mNGTAmleOSS+nZgRElBGJrgFC+1TVFMIfYF
BRvNS9xREaD2Z8hWBe/CiA5CiyQE2CaDQINQDNdqwBl8/1tbHWlsK6miOLHOjuaznb5YcYqeo6rH
ItqXeedS/e16K6wtC2LmYxIGA11MY1VvRUd8W4p/qL6g9/edFJCNgo8hL+yd47CPFHIiImvAAmF3
/PlmIRDcfu3zztoI+nB56T6vQhUjgQqnOe3hBJY9ZqUxgPqnw6rz2hw9Vh/1GqSRhPS1hHambZno
tfylZG0/+ZbfLr8laRq3BrpsC1ItoMvfF+yAejl0HI/f4HO4uw1OoSBc1femtVyrVDxps4xaTPve
giNred/Z0rAHX2PCh+SsSYXK5XBFJS8DVbkgjHBAxo8SaDRVmFbrzo6hVjYWG+w/lfEKpIcVYw4h
vmSh/DHTWtzEvI8zfZdLEmzN8uuwatoz6OLHQcMrG78gpLcm71Yf8IfLD9goqqJNoNX5HRGcIcoc
zdZ2LrsovE8FRwFnA+B80Vx6jh/BVpd+WN9+B24RHSmJfv+OEXIDQ0GC7CXFfXs3rEXTi054T4DN
ga+gXKjBhUJYAQc2DJQpiYT/X63f52VaFaCmvtE06p/75ohzL0iFac1WjSXd3FUyQBF6rt/w9Y8J
2/93oJIv2Jy2XcsFLCtbLDE6Qa2e6sPuhnVLYZ21j2ok/blHoFEqqmglhnk+EgIJDCXgJViKbjoD
hP9+AOV4tFOYl5u9Ghh7BkrYvQF2mO2ekV7E7bM+QRm0E4ZHJFWMo8zXZp8COlVjfTrEVWJBeqqW
ZiiXSJVd7TIhdvwC0IZNFiUoeqG+DCZDOHROz4Ijgp65TwggxqZppIPYFwgssNJX/1siVfkfTOwO
FPm2kTB7LPXQFvYyn4jUPNzRMySCTQSB50ooXepo/yG+rTJy8/PPkYyLfoZqE+RyN1WiW4HEQivq
YIQ7ASgu6tKQRhVSLHnad3mZE3v8WJampj89vR3SorOXhLrQ+b0ZwmRkxz4+N+2rO6tgtrmSAGy8
ocj+qGuUeQOdS0rV5htquSOLA7uvhG+fV06KRXCDsu6ApLndk/Xxax3lo1vdWdz2ffyj2wCzvpkE
c/xMDYIkL6R/NJT0EqctG3p5YaiPZfY8GqUgTKc6w4GTMFDz+hrKFxsJVQyT7YbbI+nsdohOLB8D
sDybKVBem3HnZkepbyT61x6EvmVvHd2IEgMU3pN8R/kVtXH4qRIDn5N4g8YCT+74z+F9w566NmnK
86Ucx4ebrU/5rlj3KyRGITepG6iREF5bi7xdH2sWPi0lXXXLf+Je3VyCj/mxamA2ToauVtcTH559
tw0b4dhSdMMPIQes43MigUF7YhYM3/Im/qz1PRqFbu2GKe8DfnGkNF21CEfc55Q760wIB9Ln+vCe
xWK+0lVaEehJMQyFntbSi7/CEYDpwZNZhFA8KHA5Ld5tuSn7AGWnO2R4baFQmfKgajpPcAB96zWx
8HqJaqDIiToCYky/JGs4orUt+8SqlKcKVIO8dTPV3q57Xxoj0xY1dZb2neJsp5XQyo9Eo5aEsHUV
P8xIEoEa9cz1eyIt/Qe4Q9zmKVVfTXVnHDDn0z/JsCctDeYrsO1o7YN+k8iOxN5japOE+iYOopWM
qsQzlRJJ12bUEh9DlAifMnDAmGshONPoSeOvX04mlB4w5jahrKITVNQPa561SH0Mff+R4mezd5Lm
bvtEt1r/taeY/OO7m+EfF/NLxQDwqXboBctVRE9a4RhQrMKBeCoSVyyL/mB+1/QQXv930NSkqB6d
ygrHyBEPoRL2o26Wr7xof9EEnwG03/CgmgyWMLQcM1o8u8WSm9E26V1zJGqrof601cXDVozl+N29
m+iGQm2T3XI/abu6fUMwsXaGtxMF1HAbkJiqreKtm1tGsyFFY7e/Uo00IS/RtT9XhHXJ7YrGEl4S
b2NKH8Q60xGCxFj3ENviIx+yOc2oBQ8rCEE18rLNYG2E8BBgvs81kfNMXk8WW6KLL45XaJ6EhxHS
GgFnTpBgCkcaUoZybJPApu1zZYpt4MsK96bpptIwWK20VHpnOfUJYJn67qE/axl/FM//SuEE9lxi
kMBGO3FwAF9BT0ojUJLHhdk9XeTD+TC75ZkPa/DlcU0hDdbWZzQ/f80JYN6YM6oRUDiUNCO9Z5O6
MJKifhunhRVghe9pvmKbKHsoCY22SyiZu13mZRYUMXMLJDMTyw9lYC26NlCeDz8XZgG4U5SBoYBT
Ka4XlFRaA5L1tNRHTXKhF5bVFQ472M5KWrk201AfSBQkM5ZoEB+bvRfAHNCYf49xnInGAdxjvPWS
I7Qcl+3yHtBbj3lFm0Nv+Oyi0clbKEh6w8whboOLGWCG3uaAZOXwGXAZCWZulr7JKuaxvZnRfgX2
b3qePLfc2Yk88u2TY6BHW6CkJ6nfRz34vss7qCBD9len+5ODBuQ+HBllC2vd2OV+/gABKtp4fhNF
T2cmZX0kOJKYxI+02adb6ZlUc9fkJ0CtDNH65JskMLnqOyGrP+iUaAz0uWjCCiPtAK6Zb6uaOSEK
NR/uDN1RaOyHzIC4imoDsBF5Mm0wBctX5MPoBr59F775h5k1gQr8B5pOjoqYUCSTD8/6dRCZrMMa
syKpNQSd1SMUh4a95IHifHmDfqQsdzNyKxyHNdy+wV30Gy8s6txWwNLAlt3VDgij78nVtHmbLbk0
AQhEf/zTzdlJBvYhtssxkv84MD9CYjR3rnvOo6+S2AsVF/jo2H4GQww1JdzYw05m3cTLU8cOSR/8
K5D24mTuVV7CFdBsaFXG2Pi2YI+/2pwry0hvU/DypJv8Fgw9KklanaiyVjqQSmWMxkpRsVLvdRoT
68MSlq3pIfE9npbA+oEC8Oxgpoc+s/fSVTYJ2vFsTWi8sSbOj9yRh6pwUoyaYTWPnl362IJbSg1a
BHCCVfo0w0ouU9zDQm+O/n3a4Rourqu5n9qAPKO8dbuT3MmEC/J/Jfl31Xhv5TWI0Kn8b5qz+9SM
uG8g/0zRIKzIFDuyC/q+3wht2q7aJz6r5tJ6x8uAtwO0S2tIP4e9O4KTTptZSS2ekdbyq21PuZvZ
z3/HE1fFsnNk9qCJJoY5X3lARS8ueNFuo8HPe+W7eqlv+LC8VzQuLZN7AgJmwJ23a0/ollbLPTab
CzUPsH/A3FonMBjtUL7od04HAGMHyk603edz8r0XZeqoMYs1C7o19PZQVACYk4+1cxJEPsoES7O3
sduU1OfAZPFFU9eZTkSywiCJixIQobIa31xJFngF1WbDejaGhF+1L28oFuynM59ZVImhL/I8uc6f
i7vBgMkgJ7hchhjkfKswKT489X6LHQrU2KLGGuLIpIqZCE0pj/5QGSN4i87oYNi97jbQ45cJaNA0
P7zPRV8U2JgCdyPlJYsyLuNsOjh91F4iy5pXM4GFNy+RisoduwjWoGrrGQIFNTz/6vmLUpI9+XoE
VCGLN+jwhfTBB9sC+luwDtU7Iac8Gger4SbBF6DZ3nNqakeOlLvw04EiRNoi+uIbPi+oD7c6JSS3
zZi5ytr9htwl7pnl9++uB6ffz/kC7SSjIQfWt3S43Ii171Uf4WrcSa3R7fzGkWjYY8do240pYv4q
/VvMyMphq2InZQmpEwgbZ327J8spmcreRw91zlGUA23An34ywUGG6MElgaw/dMzaFKWTGP0H5T3M
QikkC1iahDEAPUc9hkx0oNvDSj/tr+HFD6dgHC/gsltwPkzCsxqfKEHv8WJWRudNdRP6jOd2xNBB
vHt2bAk3+VXCbfwsmjt3nU+amCYNe9oUV/77w9C+FgffmFZ9kGkQb8LGVdbJp/kQrhSzJbyFHXqD
k8woRHLTZpLZQKLHCzwKX2+iLgGRbZMSI7dkEqaJVNkyk5HOPPqqbqfV0UgEVmcm8YNwpY7OY1aR
+iWEbrGV1v8ZPJo6GuB0NNUJGdpoRqJ+whZ6AZE1QCKSAk0UWd4wvicext59aW2kx+uufE4vnjcI
eaJDI+9hEd9PnpATRqvY6IrtRnEQ6kkTcltvRKTttzFTQZkhVcsL0dHbwWWVvchNewQ3AJebok0c
nImkvp93Cs0JyQaVriTBfuA0Le4RwtkuCqSr5cE5nVnGmZPnhlZXo2VD0Pc3/ImlM5cVPoSixwg6
Fvlz3azX/Ne9bpyeyxpn1ZYwqs+CPM1mD0NDxsaQ6lCRH2AA0oyK0fMDoTQtULGArTfitzsYLett
0N5XD4P/2R6rrjvE8gPV3h6r2JxUVtEwbLOK4ubm4xGHutjDuS8s+KvDx9BJDjI/yZyVJEpEg0gC
Vf8ThJ/eQc4vkwyhUAxBHTSpCqOnP4epCtF3aMsRgANX6M19KSZZ9GRBY12MyPQ0D28+9s5iJmTq
NH22mo0nQnDCRpa07VkombM4ldBjKGnZkELgkff3mEwicLTV7pr3Qu0aaLnGZmN0LkVEgsSVIOeR
fR4XWUmMrcDLex4pHNnOS6dz6g3m9TjM09rm80uTfUGonz4wkgxM+1VBfEPWemuJgNjE2rhbypSs
hTE4SB/lUYywSSr7iPHdQXKHasA07Iq27tD55zQsRsYPdsYPVsDJ3mKNnrGYlohcAPblJbzEcDMU
4TvE2d+pQSghML4oPhSVEmdA4sGbWhWm+QzhmOnoZvZVf1P7JcRCfVDYh4KRoa07PdYDN/G9PVvW
OpfKzwp5mnvdK4G+nampKdnp79CqjhDALaXI30j+5lA4utC5YJVXe9f5zSWvdrd4tI+W6KHAaLuc
Dfy4C8+WUprBnj9irTQtdreha7ab4OdJRJ3XEarN5Q8UuLvEanfR6sVbNoon49hbv1L41AfLGgQp
T/zEC2Il8nFN5CqJ1pGOnGheALoWiCJorppmy4xeSZkmQlNnRYAkDSnPA/rDajxmfHnNc99rpw9Y
toB0wcfwtSgPBKZwqUnJPccfpBr/AhJWmEOpskFiwlmjCIfJUP9jK89d1E0ErMqMpP003Go7hYga
71q1kSikZgi8BqlnCCotj17S7Fa21Rmk+6A3fnX7aP/gP7wYBkH+2lYuHJzaiOJv+99rtKS3G1M9
FHh4SaaqIwErDAttPg9AslubtDrcwQoPrdjlEm1NFB5HGsi3SIshnr8Lnrsanhc+rt+GNPPpkS7M
r5dd4fXTPv+5X6V2fhlvEQSdNbik/dawI5uUUOfG8dz4KH2c24KHa60T5RXG2Cp2aWXYPJDKA+jV
CkA0I8YHSjVSzNM+JwYyw0M2MLmvRcdxDwrKTg/09ku8nDGvok8UE5PkZe7EPlEtpv5C88uLI8np
iXamAx1mP77zjwlgce8XJjiqtnKYChidH3c3wKOHOQv8OOZawBhcP7J/usT8dSjakileC6IUIm5k
QOfX/8xo3S65b41CiiBEGqLTPHE5yiIxfeg/xgaampE4Nk1tfoRL8T6bjPzbvwfjJt2X9H4bmN8+
pMOJDtbjIqqW7IuMrpS6j7zuvsXhzpA8dNODFGdkrw3cbgkj5x1qIHoJ0BO40L9VA8nfEiW2z7S5
zTse9nqoDBrpLl3eHsZGVibSG/vkhn7nyXwy8/Bc+6We6m4c7shDriFjoYRN4PIOTLzjYTxPHCt5
apXEixeFMYRrqNFwQbYaIoGWuwmD00lsGiEV89FeMH4Q4sjO8NQ9DSIGBtnbgp3+sznZJMdX+85K
D38RO09iUt6enCr0xgmn7l2ueIsWhHqU6xEYVW+Yw3N9bV/ZHjhItwEe7ZhaNvEL21tRep/UQPov
m2imSmSxiddsyfT/Pu3FNLV92eyYseU8yJ2IQlVkFhrC/YxveT5pEljfE7PKrxXybcmudRhH1rwI
4BOSr5DrTXb/y8VeEUhZw7Dluv730bq2GRFHljWvlBZyUOnMB+IzS1+SGKYhRi2RJ7FnaqiOVCI4
vlvyl8vlQIX7wSwjAHPtiUZnzqkrfa1TVZFVzDnFZwAqaZgDKi5fOjPulcerqYo+Od1IFLTvbP5A
TqFyhVfjBbSpPxcGuzwY+v+T3HKoVOz7YufvNYFlpRkX8PtPGeWbCHy6sP2IM2ljuYXET7Bs/Kd/
7p4wP+FnN8gxvQ+OxMKsNAOlfRRKWRsacXa/Xd/XQKBKtx1hWKVcwL7An/EmpJnmgqBTRVZ6FBEO
K+NxiKOn/N4+eLXZ4iXQuHCfPvvUzL7aDHDrLgdJ2qCxlW+T/+cBkudeYRMFpvCAeBpjkiyzmSFL
5CuXOitb9mEBEjEuzEdOthKZ+jhCTnIulZVWF+ABcGtRdttL+RrlRDlTvrS2cQ0N7vkxUwC6zkya
vY1E4gQjLp0Wj7g4XpI4GKxhbcLZpHXew5Xrdy6ERjtiA1A8yvJkmXcv3mWBw3/BL5whYQNsmlaE
L4hM1pqAF5RXqNP1oZDZEzzTWg8MYXD8z5TtuiLFm/xnGXln3OafedhaXU0uAhCGpIytz3pugcWR
2yGHebZBK91YQcr1vkCrjSQ2U7vl9lWU5+55miCw2qBaFhu0glwYxiaXGQEmvdnmO68f1kFZeH1J
EdWrAehlJR7MXN+p+wsW4/O35+t3QrFNHQ6ISXLgoh2HBIcLCzjD00dULmkV4+xep9Rn/YUSVdQf
fkBvSESZoLEd2LqEFE9Pyck7q3cj85Q01Y/pRG1PwDUL1loMy4LjcyPp1ZHHIhVx+n5R63g4zQyl
3GeVDUcWP139Kbjl+M6vV88Rp9XgDHC+oZ2nO8n0utsZajYrufNYMnaJLFl48Gm2/HmfUxKOgJWg
oPImpANPTEwwMHuVbE4r1VR1pZ6IP3mFtqsSNx7xL1sKakoxpk8JvfVIU6DfylBSwyza/SQpJ1+y
5boK+p9ve1ppGa60A7b4TTRVCY8wvJE008LWUQTiZBumn6fUsnQ9RulqHItQ3vSTJpsPd7vNJP3H
0pZ1hh3X0EV33cavxgWfREX0y7hBSQ/NFpWQLspYlPs+H7SWjD0h1OxgeG+LzT/tCyVriZRJY/RP
cJomnsjC7EvX11gID3o2i7Ap+DFrLEuB8ql1jRSP5EJ+RTYYN73ww+8P3G/jtqQPU6IJzbKwXEdx
BfvpX/oDV3JSTDjWA+VMt7HaC4B7/3wpiP5K4lzuqIJUDYZUQQ3J3kcpS3TIATmt/Ay611SDHy34
eAXj8v6GHZ2iqqPv7QHCp88vffiMFZS9nYk4UgYXctjXfCdlsICZjsLoR82oh7HfCxv9JECiUM+o
kear5hLuAZapnCOWjzF3Ka1yTrI/JAwgS2NqjMK6T/K1gifLWK4UlsGsTXTFFQAH1gs4KJlp4T0W
5UxaH1Hen50Mw9mbHEdO+AlrEgRHCOwibKMxF0u3GuEPPhYWctRs0omt04vtafI+c33XdAZQxiR2
H0nw8YpvZHtj4XRtBs1u3hF4QBfiobUF0mRfEVCTyegp7aJtgtlY0cNdeRrAYUZGWLPncw0sgXXT
mjKWKmyC3H2+OJHUDWZWLZtS82qnArALIq9Vt53/FREx0tazUYjTX9KrOnx7FOVXH9h6hvCYBMGq
pJJj+lrh3dHX8gSVw5JP5ij26Ro00PBi27KOcsIn1GJFbftHOp4Ok6D1wS5hJhwGbiXPj4Je1TRE
hOk4ILd4rVIcU5jKfi/Jq3NKIvnyBHb5QIRLI2UMGZnBPfTGcX5hFZv4PP0Q7ef7HGuN7OusA7LR
0k5DjDbYF+bzILn1vkHjJzkd0jzkxNVzwI8GdG9T0TLdbkg//DtNA0PRYufkiUmfaFBo8+FZ/5JR
hpLh22A091zl4i6g5m+N252Fzg2mtDcMXyoWgwRkf8DJ6qYJfkESCON/pB118DYv6uBNJ3B/jwXy
pqecTv1qCLdr5rW+VAv6DMhK+UkOyuViVTJNkL8B6ecxBX6GByMUinn2Q9mPbn8mcqOoXK9dEn/1
Ss5XW/Y5b+tBQpsDvr8SaFY+qS30MNeOuH4D9WXCdMpQRWQVqBPFSFoW2+T8x44p7UOmp79TjlCA
O/dt6xooDGAMuVl2CWXKGZgrUovx18QlA6ngwgSEqyYoABMH7wEsVzo10/3aYvYVVvMpkHJtnk0W
JafsW1sr6r/STirIZL6KPQcZYtenHhRvIMhNZ3dRChoXdYUX9dvqVGdTorFPzrJcFv5GlZ/Wao6S
M/k/V9Gt3qn8M8w8Z7lf6St/zQnNVExm86WHOL5pDT44log/Exj+CF/aq6FEu0krgVMld5ojsGBd
7ceg+pkRyop0nmVN5tpqgYJLJ/2971baylnBX3axdzEapGLzZLKqV6LMeyeum8otVdND2Ki1/cIj
uaKuFnwIJtvyxxoI0eLFmGhcVFbumcr3eJwflK64A3VlbebDZjyOWR++rTHczbmNbsWgiju31IyE
HWHBppN5FgN3eUNH9WO+odlgbuxqU8LalqaDE7BuIfKqtitrp+ScCzpWgdOdvMA039wkMVayhKkS
0d7O+iOnNOMT1BgQ3GLB+LGvXoXWQmKvOK1H6b03BwGqXSq8p3MwLU3C75RrYtkEh8cw7x7r5Dnr
3huPUNTmkf1yp7jblwm6PGuCXS5QbggQe6RQJWLCbvD/4uZy0w0nOdMQQYBfjsRLFCrrXwiw7wTB
w+oKSRDVBnBF4lDNz7mzXKRnzVDLcxBMubLuC7ToFkH9ry4FFW+F/MevoRn1999bFIEKyvM0cpJu
JlbX44vMv+GNEzZqf0EMEvvrTuYSM+AeE7HUZeesK5lQCn9ugJrQoTJhSm8S5Pf6gNXPM0uZ0U+S
lMSDz2iVIUdAEaq+o/OdXOBmicDtWyTideYj0W0ZrvaKm7oCXBh5BjJxyiYQ5rDO2IzAJ65Jf+RM
nz/2q9cmhwrRSsme7i1Hi8AtYTJDAyTtGVz7OKOK5s6ihRYOD6mnjn53yItmpD1hXDvRv6Lvwt1x
lwDIeVB5vsGn8amgcwDPGunmVinMqDl3YuulPOKrHB4abU6i9SiOjE+KYKsyaVd+vIYcNL3dXoAk
RxP9WG5cJUoc7PRSX38I7uorD9A8EYtWqGpTPaESEKssFC+dtzUG+yUbUUGKrXNMk2zwoqZpgaDj
tV6v2sLZITEombPvsC6uhamJc8KHGlxubyTFL1xExMtYvw8ZEiFV6ZbZ/m00z0Iy/xj8XLCv9ujx
hGYrdbvrx5TKYS18vOeb4y0SRu4nC1stEpJuit8u5dL/QLLN0o+jHLkj3ZyQSOhXTkVSMc2eeZd+
h2rAyQ7DayrM0mDBzL+jHwhTiyJgoUsQSqbY+LhXHfRmkgP2uuwFS9MEDU4iOqH+GW6rG/28Wuhm
U+vhblGKvegoJVTFTjojtVUtssYeEMtVN1YYdiihlE+/UHZxYH7eumCgprOaUDuVWErXCvKn9tkO
g/CathiOhk3PasEN+QZ/+IYJU5kfiO0h9TAJN2TVALfbHIbFs/r1C/R0k9SZJi9KcIPQrI7BfeVF
O1834fW32i4b94BMXcOiasJM29MMDOSTNuLtmJk6jzP77Cx3KjuEuWMeTR1En4Obf1NfykSZtqH/
jV4BsRWlzbvIh5cc2vjCZlhk+AM5JyKaOhVhrRqgklpqlj3sko4A2cI2s39Y197Uhepl8cFGl68W
aQQs22yg2KZAttREgLqcc63aWzQqzwlzLGnTHXPL1CsnYS3566RSsqHLX2nwRI7eNHI6WRma75a5
jVd+lQVLO8AFK7XRSqvlz/qENLhJ58flbwfptw1p55hK67gJUhPRfADyMGmniOrrHM2Thbi9GFee
svCqnl+/MpkKcg6zfZ5roHOtQL+KVf+YBSeRh4Yda2i1zq470P9uvR7xxegII2HL/OWBxhnvRYpE
FK0iqVZKTZzigjMY53YR3kX/jDCmnzzPerBNWsIJ2xlxNsyratomN/YkECEVU0ccHNwOM9n6uVLm
m+VLIr+XWzrxpArvp4IjCkUcALG30aoSG4jHgLURFOcTQ+E/W9QN48S5VEPnJiDtAQWhfpCrwkeL
jFTygkqxJy58AGR0RndG3DfYoPXHV5r6LghnnZ4VIjFdl+KZBu0n3MYmVcP4FDDbZH3zesH/39za
+LoXLqDJGBCGtBT7ZXUpmEyHbajqnY0wWJaFgzG7hLxDFZq7J6CjlwvOdqKIlM/+2aAbSuanAiAG
0ivABBfri/w5KvzJP0yEoYFPdcWbYLRbZ1tdxsXwilAc4IuakSUaJTlL/iuYv7/bcDU+PNJ0BOjo
lZ/+80cWQ4zbDyhPtJewOCk9ov1a0bRIVrl+x7KKNdm3+d3iT4m5oGxF59cssb0WTWOTOsPyFonE
lzZHqfWusthwiNqWUZBnZbrIFOW21hLHxgpO4GHTyyPrPToAHpGeMCjqJ3OCar1sqjNLPN8vciAQ
+2g7sKIupr9NrcRdQeyevXVjFybzZySBacF5ilCFgeMJrEsZf9jYgBYM+pnwUA6CGAkwbOxDo6kj
Vz6eTwvyOw/KafRhNODFKSrXnByKuki37yMcasFeFz25+HyW+yIr0wbgj9JzR8Y1cE6A5KYJ4wqg
qAlbyC/m+qSs2k+1K8mjOQu/4/q5Hyt/OY7PSn/6WlNcsqQ8ZgLP/qi6qo5PgXAl8tJOM4uAqmZG
LTd6y2xWmIT1jkoL1CG50UWdKulq+DP8YxctjAWliem1C+MCE+P/kSUltnu1PJqMuuQD3MLO0dTr
/nACeLGlDtub46ewnaqBUpfcBueGmMzmm7J4k+izhICOH3WnAoh3AFcx498WCyhSlLlYLlmVWtnV
kyUa64IHscdyugOvGlkpz4ww69XNfLaYubq+PnbNHIIxujQl14DiSwGqOZJCG/6iFdof9+5W42iu
F8B9bcBaFtlvgXu7bb/dcTBfgIJ0GlJLlXJSPeeEKbSQDvfqV7dUujqDfjV0EYg2wjr4K3e1+l3f
/6xNopCXRoKXPosyOQZROC5sInqW5ndnY7RJryiG+k1QCss6oFO4KsUNUSbd9gukR0iZBR4QYnPj
P0ypX4A3p4rkKjaCv9HR2iyWO+TgVRJ69cjFj3y5VsNwMw7rZoKsXQVhlO7Yp3IxgC7J+Q/enY9/
JDQLHjLYJe5l12Jzrjp7WK0ib/r9yEv1dxZiVKozZQrM/Sr3pX49Qs/VcBGxPJjYqd6sYSTV0FPf
yHFbPx60viL4RWTru0rPVZSvLSnRRJBxLR5TfO2rt++Nn92WAqSy5lIlxJ4TtIZcPa6kHvXFtVl+
IGZzHdv5hd+FF9DDaphgzO8bRU4/G3RLQDm1s/IszudhdTg/y/tpfQP4DM9fVUqUAsKaM7BdWl2a
yM8DbDPoWiqkWwevCsZT50ox0eIIFYb9b+mXDOCJDi+9nCOll38p4pGjkA142nBY+r4aFvFXxnjF
vM8yCg7ezk8tfh5cO5QYF3G922xDkIbydQMc3XU6DNnrnfwq43aLtQ3w4f0cKuLUSvgtXbZ3izjT
gwU6O5s3w0zXhiRoZzMnuE46GxZlyouMeWHkCO+YeqLBZnpggQYK7af87e5PVf0rMup6xp9uGapt
14ph/+pRio6DHGKxtW+3PcgCJ4BUoeHsaR3UFnZdvwDxQJ+gPCx3dZoerJIBZMMFf5ydhd5P4GPc
u68UHTrHCmXpJ5LfoK+sIJ8D8r6TyuHq10N/Yb1JsQy41WPYqdnYT170R++ogNWYvL7JuKDIqDpS
X8vyHpveQEdFIK/PbH8fmZKjPU1q5qLJezpoJNk5RWc4ppxg/y3TMopRDWLMTfh15sPz0sp+jxSm
49f/eFuSWr7lfIqg0pahMEFaSTb/BOK8Ai70DrKMGrrVS2B0FBeiYsatBBLGcZJXLqtq23x37xBI
4yDJVXUHu4JsUwFflSJ1SuHLx2GpAUbRmS3IEDSg3buhCBYenXIecZ5zUwdxVLDaCHfttk+vNMcM
ZYL/ppSdUd2+X2FuPPKOcXCNVp3MLekHK97LwzhEzIyV6OUb1sAo4kFV3AXWtY874PC/8WZy9VYY
JbKavqyJjJuNyFokq63y3PUadHlZbyqJiLoNiDdvihlNm6O+kjqfBiXthIqmoIRLzUw+IqyB2wak
cL3XbJlY/PRzTITmv8ENp2qyjUGOVP32/wzobF1yNls4jvaD24qcZarQkuXwOdyo5oOMjCQW7pTH
tyEXCJzgNW65Xnf4C5bsowPMHR2PKwoGrlPsDlXy1hwgtWz7n+2aJPTzQO4BOnukm8xX8ZvD9P5Z
0TU7Y5IOlcNuVv1shugJXr7zQu+XZ2T6Rw9ySqR3wN3BNgP6abcLa8cD8R+H5ri9OkoiTA6P6Mbe
VCnv9dEr/f+dgSYGpmamU2E1WeAXf2pwForfFOdXJdao4aE+FGq2NVLdkGnu2UYJMXMsltZ3SSe7
lJSPUQIirNN7TXCwsZUwG0F0fPu3NPrgySDqk9TpIkobkwBeN4fwXL10ZLTLxxxGGsxEbcDr3krI
NtmquHYmjdD3i1YCO8yRGDJ5EZbrOkNOJm68dhNb57S4CKRS3GKkzUh6Ac755qdIU342wHIQj6tX
u9HoqtX953r7LY1E5BVoOskWkzVsv97oNr69bnwKIShh7tNYnoZsHDM79qePr6tPfuEAR3k+SDOE
r1V9JoR7GGCe72UZ09xIZH5L1j+TMj7pu1xACXpcE3dS6KMK2HgbndmgUoe5Zw6hetIjsIrfb33U
LOlL66FT+RHJ6RFc+P+q4WEMy5IOC51AryoiDX16/TbfwOt3DPaDc5O7KarLl9m/V1ZH+X+IILrL
Zuigj2Udb5jR/HACoMVzRtXDQqJ/Q47vuu3kk5oE7ZfwJHnEZ+CqDaBAzZ/QFhmpiRHvSmUO31tO
4jBPgJHFb/jEoa2HF4QXQB7KbW8v+YejU/HMlcciW810/O+gZ7Ifk93+Cz+z8/2++0ornGAhq3G1
v2rTyt6duVqsG2ySjnS6S2xvOaulFj3j5Ge+205SdtoUZnCtV+LmdQedKDKeYZGXOI2Me8E88MHG
lG6Z6qrGf9Kj5PdbLRX17x050Nh7VcbbiEJhpAOYq+u4/I01OUpFsMDzDHdGDpFd/dVi6Ld8EKVX
PKxCQV6jLiM0pI8pALs/3NUiRM70EabrvMwRt2Wj+miKTjIkijOftbsMIw6QrQsGlJR1ZnBYYtDZ
v87mRt1+XqusFk6bEGVS+8rdEtngnRqE24o6PRXSDE7a2jj5dJeE1IRd5Zm3azAvYfzBpIznApTQ
tNKQnSh9u6urKFXHYIFX4LcNQL3bbPSq0uw8hY6PffZt0rfJ7y0qA6WazmKsd14fm7ahvNISg3KK
SELFtGgE1v0q4/0nbTLnNGjKqX/ueg3muOi1KTsxRJPsbYxYT6W3B2gxfI+Jitq7QowcohzfxfaO
xHyNZy6guEuUZINrpx7cg9ZMgIUPcjNwSOSxJ7EWAyV8IvFXUarlJAnnfm3GUE/RRIZdK2Ik5oGv
FOcRJ7E49MvnDJJyF1NnSrccCs7om0SftgzK3v/TGyJ8c6qInvcYiTVXlEvaAoUK6FdZ8M6MMS+r
y3AYe4z0E/eCjrUTeaheMwddLQY73wsXrVb7yChA++EVILhG7HNo1gtkiG4GdG0uVhmcE+IB8fyi
NdUddp9T4lSzdejasMNUkzr8JjCmJbjNlGkpY4vgsqJuR8Al6Ax4ZnjhbIAGU39XXAXvyKW/+HZ+
Fz89BFDjWBfOhy5qkoczBbgkKWQl42kD1sXRH19gsD2+FRMNFtJUysw/8krGRwiowXJ20dBN6Of+
pRywaz1+go7O0YvZGgiOQvOlYW+cG/sSrshfsN7+WCApns8b4Pac4Ic4TiR81PZlAcn2GQ92msAH
LvQisgcQzSXvUmOHmZhIgMpEcK19o9hkH1IdryZIsgVjjjVdlh5e5lGY/nyRp/mXKIUpq6oiJfua
owLWRmxYj5es/30OJkaFQTV0fyxrrexllT3kzzwpKXWbSHZbwnFHKndvLapv/OCJ3K2rzY/rK+K7
v9foBZMBRY2mnDACVI1zQTsem60UkFXZJ/+8yMdkfDQYkrGCHXVmRispikiuYincB6N+ISatSrOT
cgBcX5sC4XWJWbEPExasVLFM3uLciM4UauU/Uhi0QRgXJzrfgnS07jm0HS64rLw9R/vi6F85gmB1
O7PmMBH4UHTq0GAMHYtmPQAhyA7n1YbOs7pIl7v8w9zM7oo3Opdwxel4zkO9q0wtGFOe1Jq96Lqg
lVnbh6SDZjg1no4SXD+HhhUZ1zeix1KR/uqUXS8CTNxVL5Z+VB87DLfW7Yx9rl4gVGdzr5VkYYxS
UANu/LFfAb2c29YBq3Hyo6XvFHP3TNkSrcKEPEUdyY+myBDPVipyktd//vaZ+xa4myg9ZlHZXMcT
RNzoBWsuE2eCDrwZP3Krk7L9XudG9mgHErIvF4BgKu9PubCD4wlYJleNb3ZI3g2ESjDVVNDoc+NS
1PGahX5Xko8yYa06yMrGd9V9Kq+4KYnkbA1kBhkPGszPH3LdD44vREsF79QOJ36kJ/65hbZRuJuW
7h0QGUDBdBSYRwXYbtfeJkMUmCLzF8/KyQfnI4Wd0KgIqT7THsOkRPtW8oQDbjIRQDHMGhjggInO
DwSlom5JLBuH2fLfDxuZqRD0fKLrLIF5KZ73gMoEjOPhajM/z/UkQcMjcpR60A9BdtoJa5e+M41J
BgWGERwcnSqc3y2EUtoDrWe6RHN1n+K7tJC3lcsJqAP5GbVhWJscgwAgvmGqn/RScLd4Yu+IFbUd
muymuVPvkLp4hS0eqSVAePeZzqYj06SKXXuPyIoGcxLcihM8vWKRK4I8LQrMoQ4IIe+H8NmsG4gQ
IF2WUBd6xSaPES5z9v8uOrrc1n//J3QwV6ByJgsdkvY1acBP12Nl86jvL32eYf8zApWiZDwIhVbb
VkPAPallbjevL59uxeYtG6mkyhpPfj7SAZlotjf02NftSXXaaMzIv6aRxmf56Jsxt4UjuBkbU8BC
/Se9xBkGUAiyLhuhY92f08Dz2t1ruYJJ7EuMCTLJv7Tf81LMlC2VaFjSoea4NhyZJqkN5MzJ1VuK
HNT4oFiQVUnNmIDFm7dAJdQGEEnLmK5TpMzAIQ2uXlzva4pfzfzNR2TVY0s2ZhyJkzloFCzbE44F
3pt5pvriDmcGKCO6eM/4s6iuKLgJbh2XV83vBpuljB2hAXlOvwx8EWhZ64QCmxS0mwaDWzWoAvbg
13XJ6S98vI4kO+bVJkC1LZvQU8EqJclzKURUdAppbcKVZ+M9OXkEAK5kGYNPwo/lRd9MmCdggry5
WF/ERS2fNVkBmEaPGB8htqzKLnHvkjINY8wrHhFuPeo3yoYVK6b6FXeEzEvp/xcsT06BHEAaf5XG
+MwndzG1k7cQZZDYTajBdljVsczGjX+E5dYLa/6FTw/0phoVmwPklbDCM3iV5bvr4P3L31m06Sie
6GPFsGvJ6C4pzVbPJichdauGli/2UrNY9SrGX6TKENlY3lQRbMfKi89ZnTZWCBWuJclZsPDqLMdl
iAlzQqvpIbgEAUT7GO8z+LFiMkirGoFy+nQ2TPwOIuxktZDR7N6M05sIdM1COEw4hEsnKrtYfZnT
320HWo46s8U2EtTptAKYyv2Vj1pqZKstYHyB45VQKl6bO365vw8pGkQJ706V40BomU4Q0o0v+GFM
PVnlrMrF+kyngrw5blObX1ASFcYS4bSxF7FO0x8r1vAuU2O2+UWRZUPX3vhmtcsJH+4S94RIr1tE
E+4CBfsaGPTIBUkts2YCpelRnCFBHnd7AGUHhQBXGHbEIqH5y/7bxASmasdzsh8PEjcG5Csf8WDr
qXo3uGwdwS/i3KIKHX1JQOZidthkKepKAslONHfRYlXHxH3BpePC7PMrE6/RrTBsP0tEReq/VJgp
hFYWXX3tArFYb0hGDm4gT/sYocOVyESGn9+Ppk53PRF+pTzY+6LEIL+UkTbPz5mPieZl/qdqTI10
DMgKkC+V4DgkVV36OCO3dfqgzYtA21BHJRdWrgjjXADdXBnKJVjKx+pvyRaq6gTXcItqQI5zYkB1
Z9XtLtACHktlTFhtMDug/cFOavI5j9cxyWQYcvWegfmOOjmf+ma5aDGE65hxNAhwCYI22UheDB5m
XxelFNMUCS0maRl6IoU9B56jZRb/4Esm/HySnINmvVejbEEiS9v9RXgvZ/ttwkVitj/m6PgOqIhN
ghqra8Ub3fzt2kZpaQoTrC6DwI43clNStgQcDtkQj05ejSeV7Rw37PNbZwMhV+CodgrcsqmsopYO
/60PDGvDeI2YPSyQKGloHRPoUH9Y4TdG7gKd+0tGDK4gCzxqKH4RVCLcFygG7xsfjXBddX2WtgjI
hP+9OFqm6deqp8PCxVPuTbh85lGZcPXBJdU6QL1mjnIl51TmYMmmD6xnLtoGQH55RAmO0L6Pqhpm
lX8KRNcc6EtYJ+5hd7X6N84UQHEzddCu3LCXZC7797U18xLY/AIfFuhqQG1WB3ftJ2YCifPQlR/G
fbu4vDskoZ6RmeTxWWMvLaGawWsQNhBmo82yfKQx2mS+WvaTX+8yBAc+I7fVuLk8B7hIbSv3+LS/
mhXA8CXlAxTjz1oxEphZdlg+eQ5XucXzSADrWrAR1iEGWGal8TtJ5v7S2x3ePP4Br8cz7Leyn1rI
iKvf1drbFUx92DBlmpIGsCze46o+f7gR6U80Tdh3wFYBwbV/gZf65yGl3/sW3/Bdbh/0vJFf13N4
Z2x9fNcpx7ufjKbmOcxALh3huWYckRtmYSFFKBvpdAJaWIriTW2m+nI3m91gsZjwjzX20KKT+Gxj
EZBugVzIYfqNThKGwxj9Gh+Vi4RH4ma7jECDaFsaSJf9G5EYhoKs6TyHqR+iyFSUtQi4bvAmXhbj
PrXMAu1GvWT+zUAa9tj4kPBNx4ELXXLF9N1iSU+lXioudcrbYrbXZWBZxRI4QaLidAJUidOs2Y49
qXeUoR0WbAH2YANfGSKcQ5GqB8AnXtiygjHbZGg2GeD7obxkp8LrBPKmc94zsJ1Y/yPz7ku4DhmT
A/i5iGbr1ZK0fpbf8OOwj4vxBJEk8UHlEtjuuxgVASQ8Yhr8vgEKbGU51ZWNb4p/lQKHb99kLMl6
FENRHy33t9sr7o15TUotap7RqWHULffNs2sCewmmcO65bN4Ut9mF57iNgJu7CSngIESYreBXYqvj
tyDWG2uP5zc0o7qHzi1DY1bKtWxcP0W5qg9rJKN4p/4s1zPz3+loDzsG6jD0VsPJBv2vFn3uo6VI
ezqlNK6o29tBEwaGCO40U/eWrlJ+r3ZLJpnPkD5Ev+M3BUdPVppGjcGn5fJbYFcXRPvGDF442Tw7
F/95NiBXDEckoNcwWoa0sEb6Hv6eApXZEG8JGtDWIMKMjNONdFLsPJSVQA1JLp7w9cEntcq4COct
8dQgTVmyNvgBYhZwVHCQTXl3DiuiMJapTFThFhL6ZJxMV2EoWlBHOX0WBEN7vHKObzj8DOVMslPh
eO95lq/S6slK2huKGf8FGfFx0326cj/QEjTr7XmIiYPIQad793JcDdqYe4wrsVt5bBwrwzXXRSkd
zDprwPByzGHwVIj8CZUhrgncHPd2StwZuqXuskFEQIe1hqlxe25Bh0iIPIgh0vPntrYJ2OmrBdFq
15IbL21fgGybjgNqDKxpnuVB4lZ8C/U5kRZW8ZvuCjVIC6dHNmIg8WwneXKFkgsXIDbD8vJTJPTw
dDKnqqfF0rN9ug9yD2TsIDO7A3TWDYATzHtjUAv0MBWD/wnFqKPlMKiy008qT26dwmeYAOdeNUG6
73XrN3EqgiHdbIObzLGac6sCDHiKNkNIp+leEqh5R+A3AlwBjKD7YuPlFg5Z0xG71QLATa9GiSHW
5RtPiMWmqoDmDBT38ViiYtv79EsSU1lbfT1BNhzs/dvFgotqpVVjEGz5RyX23YnuULLIG/KEhM05
2QzDqFIsNPOs7eh2Zsfx+KTSSJoMfgsmMuauokLtI83MG3WBjqMzibOFgfSJmdzKzPHvOgMrtztq
xUXDxz/2jTOF6Ao8YCWV87mTpj/YATRhkSt1UZVQZsQtRivtbD/ff9NKxid5m/Aa4FrN3MPWkQoB
54UTWKJ9b7TGlLpZ3O5/hvOEisrh8p5ymc9IRMtMQrK4BSTYL2fNMrfdvnDNnRt+et3qxodkHIC+
in17mh/HU5UuTsUsuyoK3eGNsysePgb9FoQg/kRQeueMhPWE1TXcEqIAJLYBf/VnMWsbqsWZ9ba4
XQ6JtKadecxNBgpLYS7GSdz/wm+qlCLoSvBCiXclWJPtmBqmlj+PsJIlxY34ghzZfqNZZ1zDOKL8
30ldWIO4r0zWXmv4ceQurW4HBLXPv+sHA200YWpXqQknPFZUF0DlZNEo35ULxpgWw/piRZsZK5J8
gTOf5j8mdlL33g18FBOo8+dgFSmkVJMuxYSWjlQ5ngUx32NzkDspkZZ3Vq41i8gfBV0zxKLyAROc
8DE7URMXc4IWvHuuRN/gmNqDY+jayg5JCkrJuNNpgLrx10l7ABM3evv6QWzhgaEs/IEc9xZldi3s
kDBIyuleY/XwbnFSxgtXXuyQcOYWLpbWxp7/0OZpuOOhk6EzfcKk4Z6UVfJE6jQihiytztyZZX+A
8gucIroxXN4TgZaSKMWoovPGPhqrzwUSSgm2eVcjrI84QqhBJh+/7dVu+DNrK7ZgAkCbRyz/0Fi6
z+GQ3Doqi6/WfYcDYmJaCcqxWt+bckTm11Mjm4JOzudFCcR6TqGJhX9gwrp3V4Yyam3tYYoYBnph
sJtjFBOZzmHNis3DOxSwIFZhuQLrp8KavhQ/HSJiSqQOJBgbP8woMPGa196s+n0epY4l9oJVmsvH
DRWoonaIa0PoTM5/upfHiVldD+8uqhbgzzZwMO7vCSE5jILGYOI0cshCI6Vcf41FMd84uFb5V92E
SBpE05j0CPISZC7lBD5LR+3lyV6wHeYcJZ0MvQICSLY3c0m+bjDTIbU6r9EYKKwyldd140t+7alD
ptpHw/akWUf25I6Vr3WASSy1k+1acCFxaW7Oj/GhH/EGPWQQuQO7a6grAiZQ2Px+OZ6yqnvcYOHl
oMI2igcd5b91dKTO6WP+C1nyPAMzL7AEajlOGgqB3LRjkuzNU6F57/vS5F0+x8siPckzknQpkDqs
X6RHiKHbmXKpU9aVc+B+zLRWhrrrhT9PlcLt2iDWv/yqNbeu496v+wc7XMOHvkq/n1sKxRnsqaua
7PyWqVwZ34ROsNyKi5MYaRa5qXm4+zWiJHSn8xLw8lnim6OXdOoTy8JNscPitxFl5MXnnbqu/9H3
U02j72Hi12KIAwSnz+3Y6ZLg9jdykqoFJOZI5U97w5FiPixlBrlgHHwwWQ6byYS/HXyt/ZPFxlSS
FhMRLRugfWMrVUnZtadFTPyfl3/njhJN7g4OYrGUlMVC9/UJkkhHd/lhZ+VVAXvv0qbyZHfQvQI5
/U76YRz28PxagFttyuSPtwOvTjvc40/qkqHre7YFY6pkI5ldPQQ7yiitQaKjAaqORXYcjFO++AfM
8/NmWJqpnnsZlrj1j4NrrSHuWLn24Sap5Emw6p/Lzam6SVSaFDzocQBlLUJm/tUjdI2W9axCfGON
tryyER/JQKAuquUGrqOJgnA/rSUtPUPHA7EE17FkEWtsRzYXRsSHxRqf+7XiBurtNRwwlCUgiCAq
cOLZTp1CHb8ZG0YxrCrHoZVA7O4pM6qc7CCcFU+Tft2BZyyTKKN9y4puPVMPxg8i72VqpOwkGED3
XQHjvFbzkaY8ysVUc1xkuBI2pdUUdo5gT7DInpc57vv4kFPGbQChp33VxUFYWz3PwJ++TzYAShPc
j7PuQsGn3rdyOqhjk8oRUDlCzFU/7emKensHxzu3vXUbZaCudo58wwJLbjoL2lo9P0H0aAIlUPLo
3D1AEP2r3x79GDu7GR/aRUowcStkHO8Jj/hqQY+ovxUn3QtU27hx/RHBm+rF9rcHTF2uIyQytFqT
w7NmLmHOz2Ip5d0FR5XFw/mmnC/HoYRkTSIn2SOLGRk+aR61vSfOo/v8R0JJgjp4EDhKtNhFmTYo
yAjDGf4XCplaHDsgqXUJlLUQBsUHfF+AWHjlS8YkU78OuMO1o0rAyJVB3wC3vL9KqIhXuIM0AQBa
K+rL/1XQiDUi5U+frINzrFQGgUjXLS8qzGH0jjhG0mUySsrYuH1D1vJo4WDpvYhYX3DbM+iS3AqL
jultcSG6yA+7L4WrY6dQuG4wm8SDORFMjidt/edWdEtF0oFXN9Ww5TO58nN5oKEZMCqMUsHVZvA2
3OghGEgQt8vDYQKtV1Fe9t/4ydMoom5ccm9rxEbZgN6kzzdrZ+/C/ksMorGX6uSjPnSnW+7bmUiU
gn29Y9C27ADioMiySU7zTzcmlZMVDL3dn2VbWLkvpCyWZbfu9hM7HelEngUTx8J0wTVU6sTqUdQ8
EgUl5DJS4v7gQk0Smke7506yJwBJQrC8GNXK4F8TdoQNAOBEKag2f4DRbAYRbivhxbXzEC9kkJhx
OKeWhrPECnaP2ObVzRsXUuA2pskpSHZ00o3BJOQ/X67XFd3aL4l/wiaqbwm4w+RLZmqaEiHJ3MPs
spr/7DKX6M7A/Hhnh6yHyVuw/c8xPUK9ZSrYG0ikuXxjfZZHpo65Y3ryKaWzKwKZYuOcNWGM9/hF
N6NWc7QD+Y/kJzGMwLSt1m+B2qsW1I8nxcyC8EWgVpJuEswLS3aOko2MzKjWw90uQvW5zc0yDh9B
GMGaSOxR4LTWZO7PCZyMs+g0Vg0jofd76EoWCQfy8pLxaouFjArRcdV8d9fJt1l0MeF1XA1jWRgn
tHIeaLvuZwqBw17DzSjst3mL67wf3EAoyFeg/gawAwWGNM8KTG1KhhWr2SFWhrp8/JsOBisK+Y1Z
DKfDEJmdRklRuBiCYrr8RF7d4LhWSccSMBcGjEDXKRDuFG4pGr7JtEpCBr8DmE/MZgEVf36xka4C
Voz9fT59b5tQ2v07HH+kZidZV3pXvn1gY6dOFCmirDx/HKwsIJs9ENtgYO4I1+b7BvbVrnSpGmHR
P/QCb6afOyWECbl6xfD/uagywafod5gTjjc13/WDNJFdH0vEOA6bmXbsz1SJ9kdeqvXEvDG4NucV
Q+bv6nf61myWXElwaHw7bnFSSRzvNqZVbxkJJ1g7cBLwhr+azwwjH3j66Gsncj7IDXJ8dBMcFmm9
tW2ie0CIJhKIEy6tRmbL951UV7eFRFUv/o7Rqbo14Ubo0Mz7pKtUMlHDQ1pvsokR3lBeZJ/mF4tI
rTMYA9OvlCgWO3iIH3VFz8FVtaxmPXVCkVgM/0vYsl+UYiNNQyPDwxrIUXJ/rWe/JIbNrjjensdW
vSYh9vvj9NWhECZOSFnbr81IG5tG+JKRQyVWuYfAOaV/gSjyqG6tIZQT9dnaVN5v6ooMqToNOpXn
bDSp+5UDCgezvHt+huuIKLmZj2BcgJ5rD63xx06L+UU8+pDje0/Rk89hPJaWnebC54zlgMty0DEf
lu8PObST+OMLIe8HPOU4zKH6Qyw7aXUzy6CJo20Ptgw63iYWYRNReZIWuCYDnIxdxYAg6mzzoISq
tasDp/MososkYF3VMmiUF2X6dxtaCfxEndZH8iPt5hr0nJLjm22YfvEvq64DVL1A4Pdw0z3ERFR5
fqp+brPD/aCfSzOP8tGeCv+qgi6hFPOAGmlGsIeSK6qnmIvPJMb6vvAcE5F9VPFLuB1bqP7MUedS
OIm7ePBnzaHj/LGLJtw4U5x4lweLmf1H76NXmkryYn4l9Gg2JF0REA381asq4LNQZOHb2JMJst1Z
tvU5CgwcYY4h58HFE1jmcoLb/gAVcgxjgLHU65Wtecxfk/Non5zWK9vKEVQUb+aDyOelHZohmn7N
bnlxGqmT/maIX1ML7rVwcISK7h15uPkTSwKTK//p3CLKkR/eX4G7ozKxrM89dwcmGVJtLbnPU8Hz
MAshjvF227+cmL4C4s3Z2A5/C6MpXzlDedV06/GPg4Mkq1DjD8Tq8VREH7cM6G+iAIAav5vic1VF
SNI+c+FWTme4iwyNm7y0pynZbh+WgWgdBoZEMPnf5ekMnPC0JzWTZRB3+t5NPM8WY6uizBSHPoc5
ac0IZNpsBYwKagC3CHQXTwOCLuIuY+h5C5uhpAGObQHXXOXOsT9hX5mvflB43Q8i6QEveUp76/JH
ZHePrnldom1iOl/xZ7IVneOWq+Huq9k1NegYMZZGYUWD2UcuLN4lbu7Mz5X9vh16dqfFNTppTs9w
T62GIuR8+vyRF27LvEmdX5pJsizY0oStF8kigDgOIkU3pc5Rfq+eE3lqK1NtIZs8bh5OmjbyeVSK
twt3KYSVTuUxYWuHc/kdz2sYKnGatMFrLzpPNdkbk6aC6xoC7mwTZKG7I0wMwV5Gh+wrLfyvW4P7
THRp06UKY4iYKi5xiW3a9r/ZdY6MHO0RsGPPjrjzcXyfJ16X0DiO5IQXifBg86lkaIez27sws3ZF
BwF2jxzMfGfGG4mM6EgdMxrtmVl7jKZKZ4Y04DxixP1SdOO1Ze2gSFarN/t8Qk0ex8tkOql9tmSd
eEPbLGcK/sAwg2jBXqXMoLgjxZDtVGjacyTvR+ft3pin3Cn57VT6HfUEorzDrQimtWsFSuv6AuuJ
NLmY+g/favvIl8iZRkniiIOzRoIR30oo1480Bzm8vz7mqH+TBKDOLNtRTvSmxgcdXpsF6/xONlNh
dThvHbdFUL5/9KUh6ppyhIidJWxh5UttZzYdx39WhnmmmMh1TvPMuyZKmDg8wNw9sJ+Jk0m2ztuk
FHVwy5TxZDwWHr0naN3pPkN+3MrrHhyCBfvmHpfdiwiRDqZHrSwkpXSHuuoR4O6uLaw94ioP9aIB
D3WHWozd4MLyQOkp7iblrVvlL/4VUVWZPkuZq7bii6fb/tEewrJYU7M1kZdEymcVfj5wKPpFpMM4
oVWEYQkkLqb1zLs8RLY7DMChD71bbKA9kDzg/qaurBbq09tKavGfLLualP9U1vE66jc0s+edK0En
Z3NQKtgd75vjNknHW5XDSCeV01J9P0uUbSwccwqLolQ9pvN6BbJyVmUzeIRxmkSib6jRtydMy3k+
rFH1hHt0d9Xl73ePWUkue53TQ8q02ibNLvihl8ew6pxmbQFhHseAbAd5uXU3jAzt+U//p89OUs+0
/wUDg60pTkRVJfv9rbalWtPOZt0bviEvg3IH8QXS9IX+rf/dc5ZrG349nZgzK6KzODNrr1LzBhDV
MTf7CNtMjEY1vH4W1BVG42iG0OaUI/ZnyhnTwdSVrtiX2oYlun4paZ1iYvjS11f9pdtRbDamcQMz
A77UfuWcri61e6I4upQ229YNAFEuSHDD6mB4XRFZ2bOACPywxiKJ53+KXYpHfV5yFwVBnIlATMhZ
HgaEIYV0HplfK2o5w2qugZZjXgvpDaIXiyR7EkMreapCeBHEPcdXx8sgk947P5pNqenIf8Y3gFSL
Rjk2air/djtbJaVbdzqOzj2rkynAROraHwVb+sQ4ytc7vZm9NdN7BtHJ/21dv3/5EHAHZHmeCW8k
zW5bb+YIrjQESWnYg+CIpAu8yn/lHWr4n/3CLtdQPFt+w2eBNg2CDWymHmiaR5Qal4tD5NVpa1lV
3Mx/qyh08bKL6klqc4X9I6D0KqNHI8PeA1bsMzbPiQuilcPCdYqFuqPkLYOW0Ir3cv1BJ/ujsfFO
rPVwVcn9jEnDLlWKzlI/v7Tu1BJqXAndE19fZqNcB4J9Af68sTgsRGBiuWMxRmdEbGycI6pgjvi1
6MB839t2MrdNQ1RJH8g3x/teXBWPETWgBdUDzLiNi6smap+NVxnXoVsGh/PWSKfWrg7JEA9caO2v
JyLyNiZbrd7B/cgJNXTNDpaGrUjZyLKv8buyw2et9OTmETbua6Jc7yXS8ac1G1ig2aX/HohoeX8W
2fdINtu2MgvA+erWG7Ewe1SPx5EHKat5WNw+B95syFEzBjE8obgPuLSVe7YwrR4TYBo2OAIOvSO8
RHJm8qHhVep+A3BOr9pkR4Qzbc8AWiR8BBLC1I1lUIAZxr1SaxktMqWCftqyyL3W27LOpeAuYzEE
YfYJSEwPRD9hlrTCLeMITIK8B0XhrSi8G3EfaHSodZtszZu3rjh7CGvKSADCLYjT2f4tLR8Pacat
ZzyEPVhSistG3zOYo5ohAX1VHhxiEFQABohfbXI48Z8LM4QrkQ85ZEE/7FRP6VHii+c1XzBMVltl
kdS5pSZRox/cyKg1ecoCHok+nZhCBdIbsCdDoFPvJjyU52wA5uUWfcae7CP4ioLsYlzMl21PlUPd
NPJISA7JTy7xjA5JOWDnFNPdOQTNY27V3PzoIjk8SqDHWQJoxeOx/HA5UlsUDH5IbxlJ4VcP6pP7
pNg/FgTURCRw8G+cEhC7xImhTbhYmVrlh9g6cpxl8QFj1xOZJ+pOeLBsu7hIoOfnuwpcI5uJnNgg
65hkWl3Ay1t62JU4JPKYWREuuhx8vdtwhrOmTB9FZhRKZofAscTFbP6BHV6V6yfyUXRo1BJhK+QP
GSsJEkJ5XYpXk80f8t9gpooWnI65Fuf3npLAyCKjQ3htqerUTHKSUmIM+smF7seVyuEyaMCoS8mj
vPIYfPa8oH3vcvZb/1RdnmL3nnDfhmdj/NcNPhphaNHu8/qTNeS/5AsdbCHYAr/lvTjiOlncAsz0
J4lOMnOP59Qr//I0uQ0/iogVd7qTr7sdgm5w+Eg1c7Y1gUftwUyv5yVBjmnq9FCzBo1sKOjo3GtU
tnI+cLmOdCCN9jAdThv40OYoK1cj5ZLD5YE5/HzIYEpOfu7n7tJDk+vm7KTGmIlFxgPLeYtc+FGK
DYKmdBkNzJTB7pH8Yor1T2Ajuwnxu+0RmGiBcEp/9Xins621RJkrvWJY9E5cKLQKvSJPoEPNjI9P
O1DR4JOtof/Uv92eHiG+7mbfR72/RhFJCM+LsxtQj9tWasR8nnktYN5XinoONXHRdeGc6fMRA1tx
NAveUekm8lwlj1nvCYnQhxrK99MFUocgwQ8eZ2EyG24fhzOxVUKrsn4mgQMgle92ozx844ykCHZg
ZTZrDVn2/IwsgOG2vun+R23zb9I6eo6zfiG3NgRnRoyjPse0bn2cew13p3HP79eWOAsl8exGrLB7
YhDGHlPyA+3fFRWpQz6aVW37seooh9Q0L89lki5660fHBm9dElyiw0LEKbVAbZKZ3FPS25k2UwwR
IYLZfpKdGilq4SJ2Nln1vnp0gp3CxFuV4iuYx1NoAufVoN8G4LeyrNPuJpPq9r1GAmyAp7eTAdXi
bqadvgJ4KsEur4iFudz2O5wjZv5qgW/qj8Igs6N+gBNQSLeofffUAHvzUSDA5FmUzI00mm+zxvRY
Sx51AwxL7x6yqSN8xTKl1BVzcUU8vsfpTg7IGU0/C1hSM4evX17ygt7osxFxJE1qaI79GCA1pEcX
8Sss24KTvJDv7VPS+vzuML/b+D1x4YFDi1Zy9Q1hsU79dmAzvKtdLWBcM6lRuYtm7hdIQ4i7sgAX
2R2UNoTaS52LQ6GxQaf5rpLyUHrEiJeoo1I+yDPDmnB1a6qNsRoZ3JQaaonYYOJfdak1mlsadFHW
DII0zzpk60eTJ/CQUvcIR3533rwqGIPej8VojjiLJY1dVxvaJ6LQ+o7VtzVD+qKe0wHEaLYbJlMe
+YxQtstZWmOuKyFxbhJ+JGOZwnlQVd6yJmi29PWtdfiYkOC8cyzukPgr+tslUbMdj/YMgb8LJRbk
YpONyhG9nP5g8Rcm6hPqppDvkpnhKXbDDjkWeXg5I2BR+uyHTAd7mAERA+G/ZxZiJT4AHeIZzknO
1rQCk8SbDDc0adHBHegTHu840aufUaW5otojBwMNXEOFuVBuqcLrwmvY1JFj3u1IHYeo4QIsTh+5
2x/Td6TYvnAQglbyR4zs/SjHsE9FFJNMWLUdMYcHpmSZnxPY5RADIgA0Y0fL8VtHYt9sBowhjINw
p9bdzJZ5D/Ri/l8qBl8U+XLL72uEG5b2PK+b9EAXfaMgLhbmMgWm0LCU/SfCEq8jq8sMOYqBTLhE
BcuTsnf7BVilwGh7GeveCF0mRq6T2G48NA7Nf8u5xUSC86fR5CnNe8qmjXleb46UVqSLONcrj1RV
ptCTuGfnfl+/P4zm2I5uzMRdk952psMX+21iUuUuhGnD2qxBiDLg8oN0+Rz/FuVmXLOfORWhqYOT
ojPSjXZoeGvLAXKzDQmGPKPWv2Zt02MBy1qBXGlGggC0DY0PO7gT76zGA2wWYMRuAjB+wl79pzOd
t7cJbiWp8jjOm0DeXT7ZUssDP6sMqxMYdq7E5Wdotrhl8U+IWJtL0ejbkYv4uZ3F1noKklbHSYAT
tKi1vnL2j6u2N1gr9n6F0cllzCXR3P5j9KIrPPWk662JHzScp3QFgGri8fEL9DGK2ABZAABE+MkP
+Nlv6vu9jtJwPbIS9FMo0tkeNWbEib1/z2L6rlkirKhGqKMaQ0N4trT9rKw1tn+Tp/b/S1ZtH6wZ
Ps1VZz4YM6PPXIjIuzUmTUU2975DGq0jiD2HOhtitJYtPH6isZTZvyv9OWKMfn6kEY1tgk7zKRaC
2uk6K9RKNOMCa7ad69vDzUQiKSB50QGG6sEhM1IO96GBE1oTdaNx6Zc+Cg+nGMjRN876O3EU6N5b
q5yH19QA7XN7/ed2j9OzE9owFhc26CQWPIgEHyp8Sb53IGP4xwnDHrpCrQ7GA7MngiKVRGb1UaTo
tNJ6OYcSpVeb3aN6bPwx9Kgln8i11nN+WkRZkh1Y/KJM3iXxUfNFd2agQlAEijxC2j2XM+DFYIKC
eTcCKwjT5fYt/YSTXoNsky5N8WO+OdUCeOx7Gq9OFggqyQttGNceTZ13lAh27dgahYjbS8eMLUYE
Cx293zyTP3vfj3MTzVmoAEIV0gOVVFQCWHhQObXuGFUvQmwmVadBXulsAKYaNEFgg6vIY1jYfZ2I
/NeygPOVU4W0KpxVncI26do8SSBAA8AE/vGVCUc6gm4RtcXhJD1cTPwbXkkC+aFPbHejO7MTJXpP
q5+WDLO2I0sYPcN/SP9Oz6oLbRCBgK+m306gxNmCw0eBE4F6AW0XPK+Po2ZsTHVT271DguAvggAl
A5DNXFL2y98e1nFe9H7kDPkxyraPcDVBxCTwctL5huPNNKNSgzoQURd3BzrZESaW7+9hG+FKdl5K
EQ7MAOAOwanTTdoi2Sj/+T3mdBksN5AjUxyBH5zgBpihyvZtug2IUCeYRnW9lJYvUD487JAy6BLM
q0OeWvSd94U47lDBNzTSNKM/S+A2U97oyuMCLFavD4tyXkpJw7KwxosrmSCQ1J7OzsGxI4V7Rdvz
1v37sluOiQ5dmKy5dYXeBWWOn3AX+0F2kqvw5JKDBns2Xb/R/Ny1So//dlSQ58m0gvj5oHJoNToJ
/ttqDXIpMeaDarTSINTgqq3oWz5s/Qm2tT09+QThKb77yQQM1SDxnlPu7QCagmG8T8JnKlSeN9GT
ZExRmtAcpS3/QadzLGL9HBOZyXx9yk1ydvVXxvS2xrTzGc5iOC5g6v2TnqCOSS42ec8iSnJ3J2GF
UFOHcz4+q+3cskCzCwBjN6U+60TWmEg3RPX6Qmc54t+KjgzBGqhuNrklspKEVcwu9JU3KevLmzU2
y3vr2OZ+Dwpbm8w7EzHn3FY9YgF0poVFG8l6oiJ6DKdKSZnKzdYYbZGQMBlHpKkCD7G2estHYKmZ
Y/gmvYeRYw6Gd/do+7ZzhT5TI3RiOtedNPQ9omrBlMRnUYrMm+TTzPx9+7nu1rEU6fal7y5aqaMN
FwEN8qViRukAZwPhwT+/zJlYzD4WEjT1/EkUffKo5f0ECPl4zm8yfhL66xrWe0EMN+1WcqWmwfuy
qdUakQjgkwO91sIwXGw3rjg3H0VVB7eTNamh+EtErmCcJlKDJJux17PzPU9OlRX0/86t01KGvj54
HtVSLvghf+tcjdcuZmWj8XPuFSQpjmlQJwBA0a89xc/Is9CmeRb7MO0ww99Ov44VyfypsxyGIwPb
xo1hwbGW3mVuxJi6Y7O4tAr6QaSUmIniuc/sh9LZJjHdF9Ac+CX/XJmZhV9eteH8t/SDlG2cI5ah
fgsyXOjXzH51z+9nWrqc8CMBTQ6xbkbftvXFJrOIue8wHwTDkIF+Hg2pNgIfbYLwzg3ZlD4SBeKy
3KlcNEmJZWZOIRinoxqyJyZGC+tkH+uOAHg6D2gCGylWPW7jO/tNS9XI5kwhyyY1gmkr0eGICH0H
Ukfdbhhe/NBUux+gecrOFJA1Yq4oaVdavlAAIZb4mw139caJaJR6RgVojD+Ardx8QLywt/oYQJ5z
AA4/Af1bs/12uucA/iQ/2X7FPORw2+ZjDVkR2VSMMybSd1MOpbTekQL0iHwwDX/zQtw/fM4gdiNg
OAIYKeJXX8PJwndbAAF4lVAr1OOO5w5bnKYW4f2t3v2PFUxarOZvS/3rv9NlvEwfEXkUdIvJEM4e
QvYmPXZqldcht7nhSUeO+aCzUCDRlNEfKKUScACUSiHrq58ZG6oY3WS/VDMxTuoK8bwBNYOJ0qHI
foes3ttFCMSu+k8F48QYbhWo3MdX6bS7PD+7WIaAnvg2KwTiUxhLRzLlZxIwgt5u+c9znExuZeHK
fXcDQdm0not4mUBGcoRq3AQlu3hAsxQJZa53MCD7+Tw/XEw+WoBqtTLIg44BDQGdUyE4EJpU6aVn
EOlSqp/SwB4Uz1Q/xZqiqtGD+rH5Co3MFx1hRS7G+01fvnWNuZqq7gMiErKSegGrh1Nt4tALECj7
C60u7XnecPP1hXffJTpLwHdhYNqul4MTD4SbUjDNA2/Hb02HkgGYbMJ6OQUt1Bic5s3cY2pEXTYR
UrItuDlE5Wa49HsGTJrRgc/HkiB+krhtHv6Gl9+r8LvGuh8mo1bnmEQ59Gkc5sB1wV8sLK8vax8n
pTqF6GpGLD+KoS+RAhqRd3QEKDbvDxA6mGmr8Sfe3YPuNWV+UQcViKJSeoXcaApxxlPGDOsu9AUN
xFvWp4h9Hl69HvLh+VBxnMfpkZLvq1fVByGmcsXZsTBfXCqCf2DnWucEinU7RzmMk6097Gf0SrgU
YY1BKRJqAZyHXjxhcdAvZVVr62ez5YFkeV+fZL9mDtlODg0Zxv9V0r2kYeg7aBooTbwmJ09U7Tcm
+0eWYaq1Qj86B2znWqeQDgIl7YlyLtOm3lyWPB6/Gl8IogDsWHkCM4KFIkQosg/eeB/+cRcEOZjs
pnfc5plr27dnq1KB9hDIQnUJqnxqOcraV7QwXXAYJq7T9RNcixCIHSZ9gTOz7SLutwPWddbRuo+m
vMpDEr7EOLydz+BZFAabElYr221F2LeI5SpNB7Vvx0cWDF5KxIpbz/RbW9TcdWwKvCYvAjLjh5np
RxgkVRAWpT3E2mLW6xEdu+mlV0YMYAxHXWj31XmCGK7WrEa3Fc6klkhNUF0kx+fkbExHIdpVHqpo
F3otkefinEbB6wuiXVgTJ9HSSompDV7Ax6uQ7aNtmVgd2KDCdx3J6fRCmKIb9kAUCMBb0P1dHgLx
iY1iTYBTOauGudIdDbJKAaQvyePHDD86UGUSZtbSniA7FLAKO/RR7fb11MbQqrcuGBEc/UonotmL
DN6WLYPLFUAba+oTzdx03ZqeF2ipWQ6z79cIkw5lH9ewAgDEMKSDZSXdEOZYl4rtp3vunAjSdRGJ
C38CwvlyElvBvvKMJQcK4RPxEd4CvxcU2BGRqdSI6HGKW47zNYNQh/uWbE3cvr0edMTwbecnwQnr
qN3Xt960JwRe55sOu/kczgxJTWwtITbQdK2Fu0P4rmZFhIxoSnvhlmoSQWV9T5BHUB2Y9xhsUfEj
9VWjaMJOzg5kMafIxtWKxKXMniyk6pWtytXA7rE1PIevSwT5w4bCbfYxmJSopR9rTHXBhLlLgjYK
SiLMOdDJcBYttQjLqUCS9bFXf4nE+UL3l/F3Ot+UqAflUYltV2o1L8/oLTan4E76sBogmza9/YD8
MPiw87Ek1/7ex3m7cQ1evz+UvPYzDTTemPmZ3xVMFRWFt5uwoImnShzm/JxpoKbkH/J3gsHoh8eU
70a0bWZOdL4la8Yx1Oa0Ksb+XD1egCqTTgh8dJfOwOzTXx4NAs33Lm3nXYlu1XC5jWiKW8O79sFv
XBQdR6298X/JNnbyOH7hAxWOrfTStBCCryoNCUFQT/L2ImHpcUIdKAkGFK/G0piL/U3+nCv3CpR8
Jjc9VV3QvVvKN88p3y8Cqrrf5QJMjejbxpITutAGHv/PqrPzGWYZxF2aY/j3u9DVtX67jSImHU0R
9cDkQwtx7z6zyv881OjEb/uR0gXBIK0xHbUPra/bRsXN0WHltg9Ubqn8vIoTFjrGmnvKGI0B1oPD
rWCdp5aNwzF+KHcml2bld2wMWA1QvCsA6lCf350kP2PuEh6SzT7778XCL6QoARKNbM/D1ALoYQPg
1wBkvGuimo/YO3PrObSFYh+1xR+BYlX+YdicR0d1fiDsXz23OFbPnGoRAaq9gIlDCuBi8uAxycx1
Q4BnR4guer/S2czb5mvb/oLIRxEOeM7uz6rD9HB53iaWyD4WxpkMYwYKjLbpXAKCL4AFw5TBWTiJ
D6sms5fe0FYXnQsuKTPEwUhOm9bN3zW/aY2kqJ1jEDoj1uFbZV+vE5ZeRIo/5Ye0kdQJTRVRHZFW
XU0CM6ugtLsCj/HihwWGszsfGaQJPMEbiLZtnQa1BcKlBMy/jp3BKCkIBaOnKC5iNkwn4yj9AvFt
2rzSC66z/cQbp9Tdn7PXxf1sib9fM6RXFbuxFepsnK6b3jfH4exMWr+DeKaed0JY6XaPl2L8RiUe
jJlM1Mxp81MV9f6g9sXUBki1+RvBbubNCPPJy11XxaK+GfJOOgstI6/YykCFwXShqMZtmRKMx1ql
U8TdM9SC/pfFlGfm6BCZTcNjmjirG26WVjOwBYrMevHa6JIQnIRJBXn0bmvXNfe0mDIqPwhVIYV5
DOE7gXwVSCDtAsx59mTZpmO43AboG8Ni/RzVUuHOz6F4wwxyOI+KU879cayABzivxjy/X2qZJ8Ye
UbYKaR7HnV6uMya25F0w/8Que9X8CEPl0AZCxIKigoSiCAEq1tzimAsWIN68eXBKaQLi3PZyUJ2u
hlwftVdg11rjj+hMbAHWhkRhMKiDbgZpRMZNCKk08yQxpbDpRr2za2T5ni/Dnrhmrl0nW3N1+ao7
C55OM1Jime2GKFTkESfyeylURkdEZg0wrknmLtYKaw01MqLpyeRmBfA0jRUqZex3/YeiTfwl8Yre
k0u5cPJJyQ9IF78T6SoL2I3tg2H36NDrg8dJaRVip0n6yjjoT8sdNA3L6yqifs+kIm5cfSmt8KlJ
H9R8Nfi2V/B+lIXukoUt3kSw6nPADJbJ09ZtdiHDHDte9O/anaZmpum5Sa2AMPleY8xNxLGKvO7V
WwMy17GdmJ6d/HtyYpTbg3sXMRUOpA8GyHzwsrIPkB0YP8gj7VHcRcKKwyAJYLsrXNqAhNdAKPQt
RFCcAPkIY8UYBUoB0zoaHzAzRcUWM4EysgfeyNUIygx3VEUI9/H+BBU7NETc0KPjNipGBDGV6gZA
HEIb4rnIitJAszDfrtMBE2TEmdlC08KDpoxRAwMwrrNZEoOMtdIpg8/b92P7Bc5M6PD3PLqkcPfl
zC0oDXr9AiA8n74oLk+Qzu7Jyq5iWoUsAj2bWTqzX85qGR7f8jS/VdI8SRo9rs2CYBROTmgmwDqj
9YAn6d807M4k++3NhMBLGyXD4r2Jl7qQRhaQJe8pcCgGp2j5b7Iu2+D4fHiGGhIeua6G8cXpQNyB
pZxMGu/ymafi2F3C/ltwhyGF0+uu70un9XPhdG9jZkmLc2ED0Qa/YykiH+pSjGbMGrr/drSl9vcj
YKAuWMjaZb7vueaSLJbNNxT95okk0e82CWFpMfJ1eLxZOpYcR2XBxBfSIb3eZ0HwPVvIsRL9qrxI
OV6s0DuWHOxN+odBqLLULqEenPgeQh5DQ4DoppSY5Wk+ST06bA+/uVQ2OSdTul5pjhRht5tsrJXB
4R4xTWK0mjXbHUxoNxH2iL9qmY8yhsjPMp9iR0nGiZh9Obid0hzNB2IabzKes+e6kEYGjOdlEJcD
XCM3jX7bKWHo8ymIi4cXN96ZndGFFVk2pV1hQFtwQok5iOm2FW53TXZOIwMup5YC401uZaFvLKLa
D4L0E/ttvMW5NnAtCbkGKuaVteGy7YkuHvBT5MS+3oQtdANOurVvxnz7s3VzLoiEUwMSo0Z7L958
t/ImKRJuMi6OozR7Uuqq4Tr8dl2QgWetvaXY5v8QJKMT+RI9IXlAFR9+kXJoWBQvkarDOvkLRsz9
6DQNM6nkXI4Bixu8xH8JU+4e+ckDbR+SX83ZFMfRJyB5pQMJewgb5nSkX7R1T5DSvUYpuP99WygM
pEbD8qlHIkMtRbyYvbvhZ8DcsfAHlUIiq58rxfnpfVgn2M/+Y6q30OyiXyaUApNPrBJOUyWekBby
rYOHRc7lnMYCG6/SfVstqsuHTxgmw+KhRyrlevOeVIkQ6x1tMPaU2r2Tx6CszB3+AT0DoD6AyewG
+ZqWgj7f/YENsiiViG5Ye/sny0yKvVlHnZwbHgUJ/Ojd01DE6wOhjFqDYsTSq15q677ELYvWEmGB
DbR/TOn14J5To1ZbXH7I/ywh2OAMaFE9gPpjMtSJ/hxhkc+kmlFpvryxUlxQbbKhT68WT4kIAmBg
35owV+O4c/kYwlb/OQV3NNgPOhihMp8V03pGYeQ27Az5O9PVQeT6QzD3yHKbSgr9xmVBolKb5cTX
ub4yjYnzVwyL5RTxUmNAxdTpgrm93xXOM3MQGFbz4gGCVZd/9SCbyISltYCgou5n9245D7woaSht
TT+zKwJeh0+BV3ZfzmGmai+Xb3pEnIc83q0ZGIE9O57D+axGOsifcjtOh5cLjxpka7ZMu1oiCQvJ
2fgySBkXk2C+2IzNBfowAj/B13Lq0YqR2CuJRAhhs+txy8NTgD4jpUQmxphP3yOOtMugFNzHUYhd
TiNRmwlFl4aT9kiIUwcXB/+QuZZwKX6C62s5ZsucA/PJQ10o+5ItdbrIRX8/iBUW9Ka/4rLg2Xi0
VO5K5E8mmjvJeH7BSRkfyIo+l+TL7gJxwjZ1GwOI43TNR4+7m9lRGklYBXEPWy4BTnr+jr5tcdNo
gJDtC0d4sL30xHDnkNbrYC600bNXUDB8vhGIamp7C6uoVHanSsnlJ93/Zr12L6nTh61tx5EFEtIw
alnVAQKsXHXjKzrjINUPjSBnIxhKsrHihQZdlC/uXEa7PuKJY9CpM8lfS75uyyuYK2YhXcJuLiiX
vCevPdfHX8HDT3QYqwiUe3qit/NZRFkHD33Uo5jTsjKUYc8K2RVrLEQlgVebUnhErLygQlYihWJh
9gVDeDaGPXzEMY9GF19uY03URIqlqy9+B6SS4ptawlD6+yx/r6NLnHY66xCSWWnIMQEXpN4hl+7g
4OzBIGtzJBa7HFZhZtCgkBL9mTet3E9nR0V0aG2VumsPB57jlM9UL9Bh20wR70ci+KMn1k7T4dcF
VUGfH/dKiPztrz5mkqh2B/jZIC6vbIc7MYZXmnfYt95MoLWjHfcTApkGE9NXO9CsqO3bp6T1wYJn
BKNI8jmx/d+uHrSzhT6SwQckobuXsGg3NgQlENstKYGl9YDH20bvtD6i9Zgj/P2DNfEiyzx0d+30
lSK6X73CAndpcX30gHCRDhWP39cbpu1i9OvqPPvmCYCvOd6mr+N2U0NLohQ543gck/v8Pve7neOs
xFGGa0LNaDXJOT1mpqqxGKNftJtVcP1JVT2c4EqAu6tvX+tFC/E1nq1sOM441df+l2UhnJCt2EFa
aVy5IKjywOTW+6aV3AhiQhqaOgC/VhXmrKktjzmchGD1Y6J/Rt1Ur+9FLrOPViaWWaAn0TJV5jwh
TuzdbvzV+0kULtgqyCpTRnFPpoKs1lKOcRWgnxLP4I+nxXCc5f1qIeKqJo5uusmOK+PKgeEAYfPg
KRdJJWsVkEv3gUtXhjyN/imHapdfHyfu1UusP6UyMmasmM19WdvR5wEbMyLsczlH6Z2zAo88+949
V8jYxDkiVl6tmwhWhg00izgy+ndplecKqqb6Rp/IuHaB2TR2GHLY4lzVW3O8otbQpDLeKUnKZ4Rq
aimQLlsuWNFbs/iB7Qgw0n67ME5BUBB+/MnOJ3mkAxbGJmOu8OZqzAZ+0xkYm7emiS6ArzfIdfss
o/vWVQHcWq8MvF3A9gea7xY6+/83W+4v1/Rv2ovW1nvyvtK3C0r3cVzCpzi8OYpM6x1skxaGvoBg
A8NbiAmfP+p3W68BowGZKJCIQ33DaQ/8fHv0eU02oJkD7Ynr7h2rE+e0yOQ+XRX4QT5Yo/DkVlSg
BNjeGXcqgbSLMA8Uq+jZtlLFSVjQdXkfOM/JLdTe4jogT3PiamNC82ntNUGtPgYVvfRM7+Cgc+Qu
1OzJNj398M9xat8kRTYThj0zKanJOzZIdWQ6v1rWwSwp/T0VX3XoUvrvmBDW0MX+ue9gGnG87bZs
UVQpGRZSMqwka9TTkbf/14a6M/GGvSP1s5XPPx72W0uk4zKlo8EoyuQezAoN7k3f78vOYBDeFB5K
UdsxxgdcjAnUQ1Ox6aVauQFAWiHPj4KidDfWtrzi6beVpRF3U1qzf4IJnQJD7gxpE9zO5kFHC5uv
N8LpbOGnJF3oUs+rvVIQzt9WF0nYfqVbD6jR+lCdSvZcrosqYmTZvbq7wEBLO3l1eHGzX9Qg6uU+
zOCqpls93HOV8vpD7JHB9qeKGnDrBP3DsMt3NMVjuxAtiDvzHJy9ix9679HEpAPg2NU4FiXAy5Vl
faIzUwlFkAatpBG4fo7vxCgUs/tCcgTrZ9KHR1QaLZcHmt7v6V48aMp/qVWfYOCVIF8yWs31NK8K
7BzGkOiDa6hw7tB020A8KghHNTV1Wh0hnI+vOidttgpdM1ZQhZS7S6Ys3VKyTMz9Uj2WM8zOb/k8
s9SjA5tdm8OvKkeCUAV9CHDOIVFjU9iwrhFvG3Wa9TMjxJvp1kOTdUH0kMrnvp6ADuYWsqsb9Mdy
ncORiTvB/c76fuITqm9MWmL6ZXYZKs8FPjU3iBDYDc5H2MVUIF3uGVw82sBGKb0+aKqu8o4B8fje
durVhXwn8o3zvORUXDVOi6TWWFOT8oaalz7rnhApI8XK43YV52md7e/qjWggQqXfELH43/we0lQB
E+VUrGD4i8AJVR34+ajHrD69PsfEUlpz0oA4vmT4oE8wTQ/ILFI2df02Gkp1r8P9PS2QAUuG6ZW1
Nh6tYg8WK8FT306DiPuS1wDjWJSoR/I+tGKSzRqVdvEBFt6u0IOWvuo/cNFVrJpCieGD9hkXkex6
y1/rlZgMmFSd0GkkM9ew0EayNg8ArcDFkxL94rDWWuZR5u/kSOr3iLOn+BrEoKRHeiIsz9LRoeFU
aJk1mWfA130xwhgJ71E6Zx6XV/iQCHaS46lOyCu6F3ddTgwFd7d0AodwP3fpu2KE1wsr8SZ/beFG
6DJTbDDAEuijYfSFdi8p4YDzAOOGCB/bGAPgK1rKpK66j322bvJaIb0e0/ZmjhdLiQ8useYfodYx
+nUVkEb0OrwZLGBPyN+334h+ffEAIhxbOmfiLiYLjIZQbvZ+5hIheE7aQ/gnX8+PijV6pjdqDjEg
raYUsrgO/WHGnv5XwpJTqTMfceXAT09Z5xsy04LIJhkstCpoVQNVCgBgxHld5YXDlGDFsruY2FwW
U6zkIf2NAWoHxJ0X3o2Spa+cNYf2D16NdgdGXCCIk98hl0GuRncomQIA0kIY0WYovZP8XeRmEAbi
Vdx08wUOTTu3bj3DZgvHN4EA9josbTgYSmz5nd8DReZ7wj9Sv7mIC7I/o4NsBUwIrnyOFN5ixrYK
hayLhGwZYxUcNh0nOjRxe8/9N7P3SLcq2RZURcdlqI4X64vnlem3PB1c5mteBuDPWerCVgUSsU8P
7ReyciHz79fGZOL8475ICPEIjB7p3NhynmRev1f8w3AwIG2MY9E/k1IL+P3lC0fAAkRwrX4VCYCh
qDIKgdDBv2SRLyRxoinYCqiw8Lo+egJWamn4xqVM30Ot37/XJFVy0oRLwIX6tETisr934kuAcUsd
e+gfEvgO3rgqQGi3X40yFkM27mKC+0pka1MgwqtlqxPzYtoafjT0+3cA+giJsw3pUgeoVJMSmZJq
wcbY0ZOpiB3/SKXXAlLtLEnLXvAOeXFwf6HVMkaPo2x5rCeXgzZ4vuEjGwz0VaCw/YmFUgbMh+in
HNSoMuUS8FJde/2+8AHBaEhz2/Ay8vVZMdnccOwoSsayfEbzYRcSLdiVdRBCc3eR8ApTsg3nTTtl
vcNpwhCPwfiIl4KLT1Zit5TGfPw9jfepnuzfHWpBzxMPf6j5mHhteSCzuK5Ytbcqcsmb9J72XjLX
3M5aS3lIxceh3uihm1vKTjpmDeS5icjSi2KC3VWRIXMdJd6AYQoQc1D4fsP5/VDv8ndmZn3XBrxb
d0uJcKcaktjUmaSoqhuV0jBt5EF0UWwVe6o1XqvvZAezAo+RpvrU4zSrEXFSy0WVUpxDPM/6RztW
T4RjCntFWz+Qw4xJg8ek8D5XgIXmhK3YBmkHqdAYApiCgah8lOS0KDj6FFLhcwUjIRVDyE5TWBep
2m3jmOSoivsCFWVQqevRSid4aq1KJBKnzjFEOo7L6X5AcH4NB39b13To56p73l5ZKFEfAm6oyTz1
qUq4JeCbSv6ya4Igti5FLOcxMhnweeSg3OOCQvhFNGNpSSKg3rRev0xX0k6KPz+cEUeqrj2L6pNo
6cZ6GuOrnD7VoSCRzCtoHB+Vn1LDlT/bN8yGxYASwmmPE8Wh1/x0n/v3sqgBPwqyUUl7IiUhXUIf
p+GtphU7U2YetGnFmchyo/FsFvphrr/EJ0uNMVM0akXpyh2M/gkQ+pbcXzNs2e8Fg5SWI7AURLtQ
2ua65vyUsJKb4qVxCKUquqISdglCMmnwPsOk83mgy5O5ubAxPxwF3yzQalE5MLk2fU2qX0Ln4Ls1
9MAF+6ytU6gn1nlCHPQzPgfSmERb9KWQ+02K1W6kYJIOxGmmOBNywyY3slyopf+cc201Wt6eXo+N
u5nYj92QfO/MFprawuXEDtLT4VIZ6Tt0l3RqlT148Lx/qPlps0zPDHnKiT6ONAmIk61zGtoeQkSU
bLrpX1AKr9ljaYsxGklMI9BsRtLxjkanCJXCw3KbobCvYjYnZiXhMXqv1br13kC/NREQtiHaMzLI
9oUsaUqaOZvUUz9HLjNDr8Y4PIkgE9PKeuELC6qyGKSNokvxCAq1Z3TIvmlAdhg/he9zFHrgOaKj
zcvcsdo5A0rEpsVjcL7qJ2nW51wY7QJPIdVGXvIp7+UMyt32Oyq4zSOkhEo00C2+zxUAPXbRdAL8
vowsselrcde6rC12FVStXX4PYiPwd+8PXGJ8cYHFUt2CNJbOrDJiusYdNxnBqmTvLJEwWXnpF15s
XcHPdGqg44zOh6thRvhmIDWot6FegxFWFhqqetK9fVmf+ziv9BXzfyTVi6LW2Y/NsP1EvH9YkBxm
CuCNbF633LSmRk96VJEF1OQgrHUN8j+WmjGbEt0iFKkGcOZglitsI3i+RRvQA07wqLFRFj2QQieH
S5sNPWT3Y75FrflBWLzo7f0Z6YrllQ0+Aaj67a7UZYx1inN5/0OJEUPsnfXb9woLtnp9KqKSYABa
5XPYXr+tNJITr99oz28qos+7KuF56TXWhDRqM2Lj2xzPecCK4b66UxpZoWvaM6SRM4PEH9Eo3GPT
uBCG6Bq1WL6FUgJ9qahJhpPuyOg5Ghdjmt8OSGLwTFmICQ4TiFvncrpwMqxflvdoWqHf5HdY8b39
f+8bQ5J7NTX7McOPCtDLRxjIZb2dCXT5GaP0u3mTQSf72gQl7pnXb8aPEoLWayMwZZAy5ZIfTfZ7
ShkCnIHxkBS+C/eKmXIQsfe/cX2BSfEVbU+iEfksVLjMoC4Szn2aN2mxr4+3e+OTlyTLxFyx618k
AgSpwxECI1OG4BQ1q5fZJ18IYS33+swRwr5pHU4Q1mrk3m0r0rp2WEhvfF9e9si8vqKv9lDu9q4n
90LX5dZtZccBrUw7gwwf97KFxjuW+MzzaaGdh3ZU1IB1PCyiUL49jyhGGTNkRiHf+3JCEfV3hROh
NcRxxLs60M1faFEMhLI3nHblCgNMEt7TuWkplHTzgO4JxzlwTkFEQQTeN6bQcM+kiMfnjUOGWVbA
IJA0csX9/lc2e+sCgZfhc7zOgzKqbBH3lx5Aueubd32xH/AnLARHtFAFO1w3v4nP9EX3xp4xCTW0
ZFra84do90zppbJbLFoGDVR/vA8zQvEJo/tgGowlmEP2FceYdm2ymGRTRgfo6flAqvhVQxbhNbNT
QnXm9xg5wQahXxJvLyOPbPB8Hw4PIdGesxA8e3lY3Oy3wR+DbXa08L21H7ED1Udsva+2pFaPXcUT
UqBHvfjTfT8zbIsb1A8qdHnQJweADhQU5CH2LH+4wUQTmRTjUI204Idi59I2xk7T05Gr5+e9UU6X
OzZ7LRo1dugPhT05q3DE1sbrRmLh7kEZM+TWTfCx//GVuzHcY7B4cvMwT3XSEoVRtmpQBoHIQXTU
u7L/38ecsjm/IzzlFkg0oriCeyBVSVGrr6g2rvXCCz1VrAirI3ZghbeqpydZHSlCiReYvzV6iG0I
lLxTtSj9w2ZStuGe+0lQy5Gdb1GZ89LCed8XXi3KfVcSKxiAM5VqoTKL2iMlaIBFU3RbDosPySQx
4AnrV3eJWdCyX8BAoNAontkuE5faA0uZUgAAZ1t/PurXVxOieRZSTPEI4Y4nytLawwv82xpnAcAv
hb/l6PK3Xup75xef00m0ETW24ek7DAZmIHinplOBNtJSxarMGkUcLWwQEiUtAbDrtkbNFaTE0ML/
rXaLlznAf++d9l6ZDqObSe/cFi3xZEqLRJoU3ya2h5aZvcXK5jD99JQXu17qFlvhvmSNihFlGZgs
ZHO1sOPIoI19U9eLhgEsPtdlqjlK84CbvVbM6k8TMCSwh9pVhPWeEFUh2AcJUKu2SB+LiA4MqsKj
eh/JebXu33vceud/O2v9dZsjpOrPtngeq0D65rdsv4dXxG5vP0f5JrgjNP1FAei2pc3EGMdOGQmu
jOxJkSASuADtuMahtL7JYhzX1qwXtVCFKueYEpICDy5WJWl25W1b66aUfHi9mOKObTf/GFBOINTi
cCuKlcXaIogjsnPbiNswGtpJSE1YSIhOjb7EdtoDf9uSlnkoE8kHyfTj+S96pnvlQ/ciW1V51rG/
V5da7cars6vhy9HTaadiswGFO+NuSvwN0cdWILR6+MqkyYfi1vn6jFKlzaQ3HTcWBqIrwZL11gbP
brAo/IrvfN2gFit9weetWPGyQ+2ou2Lv1J3jOhnjQHkHFkGC6LoHtwZGY244eMjM03MRjzoL6qrX
Ehirhy0vpszy76zQCsvFn7+opiqmFxDw2vqVu+9xVnhe9/yPG4VhrKWRE2nFjEaF8UWhwnPzsJqq
Ydx17W4jam7QTEuGdBmryXuxaTAibBAfBOmzMJr6NK1RwNv52JRZRYU/FgdEMs5GZKd79R7d+oot
Z35UhEcR51rBIVIZXq8FUoHfQGxTizU4admUcpfjCGsIXaLJCSSacUYMq41ulm3uIgb4aryIW3mR
qAecPbDBZh/e255G8tdJ5FNPwjgmXK2bO04eyS/8MxQ/Qcb8asJjfAxxStWUhp3kOdqd5cd8G/6W
0MdWfwz1IgW/DFQmDm/tX8sCZOlI2IqpJjz/i6Aa/OnBgOXumwEt+G2XhXs1/MLia5bs+UUdY9EA
Dtbo9ljqjQz0hQOkqIHfcnzppg4BXb1eI20JAflmgRPkgmeXfAJrJJp0q1N3TU3op8vw8V2mw/62
9AfwXgmvZGdeQDdjBQYkj1vMN3gB4GbP8CaaSzp5lCdfbt8TxhBFhGgXrEeOEP1W2ppckL3wwJWd
P4NvwfrdzfIiG3rnkwJ/VEVkS1baTgZ5PhV2dUaxgNwh8HeevJb4vNYVB8jH2wkn0bGOygj672DJ
BrEeVqPFqNQ5qDMflKOm9HeWyNTFEb1WP6w5mLwO5f4boAs74pasaI7QnXT8FoCzVtDmFDZG/Ste
JOJs5uoKyVLRuZ2eA0sEiZZLmF2wJTZbDm7hd7/Kt836l+DQTyooj90Jn7kUhQWXA8Rm2aJ4pdUr
5fFQ3bBZGVmL/k/wfWyhuB7GMG17P94G1Ua9r6sGCArLXJBQPcH1b+Nb4whOUtpLhH/jqwNmHqQf
k7hVCi81AyFYK6+3y6FrmKWGqbnGKknNF38J2BQLiYi3vSSZjgL6M3m3zKRyX/j4+I5rdUlVMic3
D8rgWIcVpC7wJLL6osZJJQgzNwUAvnyMvDnySJkh+ZczhrvYq8JcOJoj+pf2pEbLiI4jQEEEuUZq
KjMveHUVyTdhjLJc/6dpQlvWkOD/nMFhCDe6IhF+SzAXYy2LCbpvrHH4WirZ/Nab0vKk9qnYM7NO
ACHYx1jvzlGowy965lOCUvmJRIr79R5T5d3xOwDSl4EHCDq4DbZAP0/saMdo+nvF70OEtmj99hS5
2cvPPpCl1ouLb2qyW09eWkSVM56sBwq75eRECtLW6xZrGuh22y8hh36RIGZ6N3mla9qq+5wiW5Ns
QlCkb+i/Z1vxDJHPJBlasyMxDQ0IHVMLJynYibCs8hcD6iiemK22MpFsFtBFuDE9ht8dXORQIR4/
hSrj8kMGuHptz3ybNYv251RnQhSZr3bA5sE2GK/j5MLdCFmHnzWaPKb5XgIobAwKPv6y9fO6aKJy
6NxG+5auN3bJ+xjtMZUFj+dsMq6C2zx5UUVzfGg+98TMO2Oiuxli5DVS6PYhWy8KdIe06g1deeXm
qhWBKzzHgF6YBgC0X8cO/gAKlBAkL6WtHAcgRlhx9bjMUfxn0oxPIe0dkgFrP44Qu/lWH204QQoM
r9d9umQY35QcVpKK7ZTSU3ER3eIpGKcvqZ2E0alxeHcvOraIpI1Wj1dvmZkuomLw1wxlPvcsO+0j
jvJwB4PlV4qVT52ik9SwR4Hcfjck30b6i+M/bogs/c+Tn00Vh9OPwE1lXhADONKhZMdfjfrjVpme
ksJuwwYTZkblpecztHfPv4jZ2prGlogWECwgvTKFv3a6k72d5zCybtg92mP29PIooNqbcOge1UOd
aKLW2+4MzctkML7CpKGzElHwBEhCvxr485ZJ3TELrcv1cLy/u+SVgY9QlJGXIXK/g57TeyGypQx3
aHjKqdVAzIBcMs13wj0centxZsI8ksvjdQaEZcHyzJdzD97eJSYkWmt/7pmeQR0qXu1hvmB9GqMT
TRNZc22YB793RnxxtVIsCkkYZR18OZ8vyNqbQitDQCK5EUEhl0BAvyeKVQ9/SJVl3RPPX3t85SUR
3pd+pQ4sjNmg1G1VnbYJw1UCfYJ4BSnDvTS95x4aJHNVM/spyWNM+Twe4Sru+EETqtehZTEZLJy1
/yXl8pX/MQ9njIklxMJA+yJtwaM2NjATbOd1jNzdwiioVvGJF/jEGS7K5goM24TpaLtQvgO+kNNl
H41rPdSECbB3E6zEwVTMbeidLwiSdgVefcB5qkkXhrker2DrmiuUCRAW1MOr0DH+surANXVcsrCP
YuBtsk0ZHC1gN3PXpeBn3F7heOQ9Ozf3HV95ELkSr7pB832g6VO9/VCmRB4nFarrE5WEOyCx6EUZ
J+sdsdCrqtUnWiQtMzOo0CyFRsqzM6bGK87bOjlW2AijDxILJ70LdlSag295jNWSLEKqr5g6oNP4
nBokN7fq0I7JHN+Ygi7xBIVrTENZToGdPrTHXsN5ERJ/LdueZjExXJcBlkoE0UOM/Hxlo0wxexWg
wA2e4oma3fW64UtgoGMl3bliYDTplCQ0gpNkXuX7lqz2SzXpttixDaPK//TYNUhZsCeb1wz2RjU2
5IcWAqz8hP94zoUkT7/esbOPdbCIkXh74xY5Vqnc3h6+FkG87jFCzpMklXMeOuuWvKd3FU5kqc0C
xfy9N+dCLNGzlZawa/XM05+5tX/sUxzUSxxZ5aHVwTtSw9F0gT8GfM+7Yr2YGhqpOOEOrk4pa5Zc
6rjnnqV3jsnOgK3/nJHcjjDOb++q5t+311qTIpcZsEV8IazRC0tg+6z5Kbj0WDpwAo2Imu54mk7y
eCg+ZmvgKen/SvfkMAKAUHWOcvTixJNpikv3iPmiDcTOxpkegU7BVATlGhM85XNWIb+rCxAkmziQ
s0xMIIcV9O870oH3mOMCU2xcRfwbi2XsRkkihrdsN3vPy2wPqwEMwksIfX1+zvtjsazPaQD3UskG
muFWaT+lQkXQR/CTxaV/r1DMwqktkhZcmpOyCUjctGLXMj7hKW7ySrtvSGcs7N0zqs/0Z4v0nbnX
k3k+uz9DgUFfa32/OWlaUQpcXGatRuu0zTG86+dXIZ5Cf1VLwDvGvumbSKMVTByMJh9tPDw0LTQc
t4urystkDgaqQO32m2rpYAvxOMm1srJQZrNkey11p4mLGopI6+ckYTBCVH8W9jpt3fdyfQDoFCAq
cvrjiuUxi0jwgFeoLPbwbvAF1xNPnKIqE2fedeMdCKMHViprhWvarSdUcxj3jNYPestZ1zXEKA8d
dIqpkaYL1dspc13G9jZRWMVJpS/fFeGtGB/MQWW3aMwwGIwL9wkbG/7pOZVOpk94ioOApWaB8v/m
4oBiIgtS2v39WemqG36aH08X/0wzSWgu7b+mOdk+iUf5KETiq0zkfIk1zCUJKXzZAf/CL6bngslu
owBEfYLidgDBh/rHztVrdNcrTSsHR9Sf4I3tGu+Uoxz0UZjfddel25v8WkeMKRN7ZfvlwfZNo61o
IWEilsQy4ayws1nhsDUTByrV0wZmrrCAkGTbZFZn0Cf2eK2OfOyn+On+FoIUQko1sKBRsoKb8RHt
OcFZBYeohL3CyB8ymOGr4H3ZLuVovqUdULApOSjzMXhhXZi7r+97nQ32hfMDlmiIYsFv5dF5lfc/
vHYfs5HiBcIRU3/gFj6uoecXTZ/p9qFm1544lp8Qf+Zqz+GVHWfvKK5obFMt3ZlCmyWx5ejwDyrx
t9LkpWdu9LFQXKA3eO7VFezazEJTFjGoCo3CqOpQfbfRTPtIqZPZS8TJk8UnUoTzoVPZ/ZsN9HQQ
GBNMa0X9GKR0Y9jU0jIh3kp8w8aFuMDgUTeX7lGXseQOW6reqbDyzCQCLNTt+i/+BedWju1yQtFR
kE8j6StCL8WzczUTwWg4MysvSiIRM1NkMe5/azZzC40lfbkzheLoGAsUscqgXaytuWCG2iClMnKh
lnE6yA0gSoURl+EaYcJ00HTxgWMEfly6p6C16JFFrfP/XSjaPkW34bYt8ye3t2z/OhooWZ+fy8W1
1lSSH9YXlXzR0o///cAkf5wu+5VJSsvQ3HTxBkiNKzb5P5MlkQRELrHVNyUe1jzOIs5jfArXAmP8
FUNF1kdghR8AFPRSBQBhYlyKb/Z7EJKMpIVW/DHEsjrfWed3lFaaBY7MriUZISujFeu0umjyyMrk
jKF0OWOB1KPS0N4y20cy1Ku3Vzg7CQolxgD47ZUrBiC4trxoTXXdS/xKqQB1RO+G+bDmnQfOVWM9
fHpOU54kBpd1iHATtzh2Hf9rEwD6x0UKjMIhRQ9wbxiFs4bc/QMOAX2HK6AKt9v3qgbeRBXFp5Kz
8FFQIilKLGkBUtJIsOOy22tEb7Q7rSOlUxmi+daDHJ8DKZnn803slTYjl0/BYrQbCMBSREraA5PR
wTbejp6oiiv5lAvMu+O5m3jGJmKkaynHxWzzV/55edglkqXY/tmy/HjS8vwMzaV+HGl8lYbJ1iRF
JC41S7dXAGsM4b/I2G1PqtwEg9tN60g4msp1/sXGAzuqcVbJmeY9jU0NCO0Erimer8OTB9Xl8sj3
JIZPmr4Voiy6nKnC2ocptrJh3NUbT0j9riRUMjK00Oi6+vLCPG4kmD0qZkSeiM7Mmdp0rBb57PGx
rlqNmrG705AsHoVWmV9DkXaDkKPy7FUFwPrbZIozq/60+T0hFsuwkPIdzsrnbLJ3vVFdKNAilFWL
XsLT+gkvXJ+1bAFFerPhH0UmPfU5iuSE00xrey6tTY5tvQ+PtPW9dGM101NyGJSoekyDqycj2Ffg
GFyPwrLQJUdfcpQcXnY8VzAgWa1nVjNccBuACWDB4kLYLiQ56O2Ubpl1JIl779KY8IuW9d7bGgj8
ZgogCdr2fFqAWEy06xMN/v//vo/hiFnDalRCuqygTIeHOvCQyMJ7oN30gwXeqij3qvlbNx75TXqE
m8hr+bvYvP+/H954MUs/F74ASx/7Z89H3IDzGHVNuBWWePS1jJhjKB8kGfSYXzcE7k42WLuurf63
q4TNifjQNrTRiXbRSd+2cmhTB06cJoJFk9dlkIodyzuWLPqx3KC/SOHHe5+w8NYV0rFgH8unukYw
6xAxfbxy24JZgDUQ+BuwcS0OHpNKSb0M4y6FK+Iqf8Z5mENpGn2rrylpYXq4rE8+W26EtEm+1uCJ
S3IwYr1wWZmLul1hudtYHEQ3ha7lOEO69V70s7sChO+m3gnMGfUMynxB9r3eJHBCwvhzLtCmAk+m
vLwf1c1F4RBie7LjIlqUykrwkwaI6Xwwo8ZIhJ9BIye514d8ysDhn7JWAxyeIh+km1ZGnX1HxmKP
QblAhWtF0reQoXVyvYR3wdxAGsgC3EF5gEjdoQUyewWCM+i3yLbA3WyT3biw742yxRKmh1FKNwcs
zdZmyEWRtzyegATOj/Xl/+KXBPVkZPws7OjEqqJVAPvj6ulPZcnfN5EPkbOC6lnq+D160SH1csM3
pKxJG6B9nzo4guuNvksvvdZSjShsbY86b4KKXTtJkupNqwuHO6yBpmqP9DoOpBUWOiw64xLEQzZu
VTwoYxaAVJ/lOZ+cl8GAiMntgypJzbipl5i7iLk4vvhHUowsfWmi0P/hxVinT08hZP6E29Bc2K8d
Y4IAb6tcEUymMxj3XwJnnVDArcUrygbni3HhCNARaE5zKl+7BC4trcC4sR0QBWQgXYyYN4JAu1au
T+4yetPNKwC1U2cU/kj1jxtPiJTD5m9ieuQyLRruXXIo7BG3N/+CukQ0/WrRHSxY2eRPHuq7hYfo
7dRQkmIlYhYNBOlQAznyptEebwApn+CgVMTnMMSxJG05JTfuXtrhEna8KLiNSqze0Srf6W40y95P
SQXB09TmNuHnO6SgEYslUfAnUr+8swrWlNsP8LH2ATjNMzctA0GHX85/+28GI87c7/uLT4gG/xz5
MruCnXvESrNsReYgQAzQKlT8+VRXHJTrKiSwfB2+wcrfgPbFTkkE65mKu3c8wwQigfMa/VclJQp9
ZadbLRPLr/8a087f00jXEbq1bJA8r8LZZPwDhOykjmWqv5qWcxNzI+yeRASOtPBu0R6hVNrqh1CC
0bRgLZyphmtnZdHBxssAAq7EEZkhAZHEstFHSEz45keZaMhddCpDUvr0nZsEUeqfPHav53kJaLN5
w2IzwfyBk3XBjYCj88BAHS5N859W3hX+LQMcSXwGNNYRiwpI2lH6uy1ysDHmZyicpN//O49IgjSr
LX/YDcFhTsf2XSNmk8W3Y4Wt/SIaUIUYG6rTok2SKN9nXWdRfPWRqK7uYRjC2XbEFxUdvh9yyYVR
uYYkkNd2srd6TfedFt23wrNoOlDS+wUQww5U0aGZfLk0Q+abItAnIUQZhKJzQPYY/BUUGUn9kv5l
NptU5oEmNe+nLdl1Z43kw3gAAPx75RA+qUJEvr1F9ZKiFEYGJq6NHBCS7goZ3e+OKASvyCHw2vKM
4qUmT+8yMcfJB2/IQjbzQOj7BZCghYkJN5LOfdGiRY1a4vGR6Q7kME+C6EldNprA5PjsuJKNGs/4
oepgCIRsPMr6n6wROoYwGm/3oiukchg8oTpfseQlri1b6t3NNoEnqkZHTmx4PxgFS3NX+M4Bff67
VMIjR+i8epAbC9OKixEF77/glp59oq0XXbG+vEfzv8qh/riYS1pMNyN/+8FIhk+mT6jQ6gazGOvS
kuO3/rryWAAkGyJgBRsBMJZVRwugLqx5lbDX2Hu2aFuC6Yv+IMJ/xfnOAfyEZiMnJzOifKzVMH/4
VyfZ8QrzDbOUV0HwjgDdpFiNY+TrNPLxUhFjefTyU4uaNKEzTg2xhd0ie8PiXROtA5zvEFaWOVKI
9P3xHtXgp5JyF5mmeh/5bPeiTbx8WxOmCRcCCDY5Qy4IRD/ehMHYYgLKiGGvODEKw0fnExibJiC+
w0mSrb2QJtvjPI7htE+scgK/pR4OeUYlPo0YrvrHyxyRccX1Em8S6Jn4AOJd9sH1hDqVbdGMR4cw
f6iAixuVFYfcl7NeKAmZqC04iMnc+E6BhKW/LLdeKS5TMEpOcIALKC6R+1BxteOwP5eA9ruN2Xfl
Er3F/DK3Zv50DKLS5HQoMSF2x9TXKi97xEf8wsmawgQThTO3UxmU8p57bh+P5bt/EcFCORzBxMiu
tjQ//wgEcjJw2NCSJw0Hoi4Rx5jbG2VNqaSPykB9CZnVSQO4lQGe4l/kUdqWCpXPFfJygZN8rkky
Jw90xKo2M32759VlpVjJBcBdSBUCexyimP0i3RTL6HnhVVKsexlBsHe4oPTGB8kbwRv9qM90hm66
tcNu4nI4yzEY9rQ7wNd0n5kenGpQKVjErKN9Rhd6CGNhhSPGhjgYea9d8JsO5vvVRnd/W+Zayitt
FOG9InKjADE8T84A5p8PdoV7sKUf5ev/uvSXlOb3ExcKuBVCnCylUKbnkGcmqEg1RtKprDXB20wp
teMqcYe7AZ5z9TiHd79U7VeeCABDFHEGwNl1BJ3mABxBJLXNKU2LTYZUg+HdYf0o3zPiP91upio2
DjTZFtsu/6ECVCS0ALV+Ckj/zA7fZs+IG1bkWWE4SIb4SzF9EtR20CgBQPaik8D0X0T2mgQDls79
ijHeYX3ppcrqcj7giKElDAVmo7EbEjKq6cl9FKkxvVIvIk/WkbZeTITxHQlLdAQ5wPCy1IAO/K+P
yeiMxTtsScLgAfkENLikFpr58VOgHY+Bmd54OlPVlUvMCss8Xg7j17JOQMECQAzwRuzMAMLT/vXU
BDmF9FsleNRlX6/knXzFCAkmVcGLdO2u2LTlll//Nz2lNRjKnsXN/GsuWeh054Y2OonXSqhftDic
ORRb4aQ3KuPL3x1ZSsOT+9FrSwhRXBuW+n1S2zVEJCayJEhFvrPZl0Kgj+A15qyGsNx6p/MwTbfP
ee9rDESAmx0/W+a7lW1nSi6KckP9PBq3UXxhNV+ABOmSPI+pujyqoMZeUnADqnyygIlqT/lQhcl2
wgFJt6IAO0hfvqHNWiHd3ZXM2LN6fWlY4RVNNrmjCIZi/Jd8fkYQMUpQ0FH/DPb74d8I9TXK7LTQ
Xpi66BEe5PaCDOswKLZpiVnShY9jeEwXrQ3zr8ixIGVSpK7wJubVOZNjjOOl17S/zKFWra8tp9oe
uRo7612bj1HA+RJ41OKQGPEh660Xtbj4eG2rPf1dJO7c9XG8lCKlWCT8TZcRRwc2+VfnDoPoWWck
2yidg0CFezRKVkYILYmAWVkd5Qq/3QYA4B9T4kqUvGeFJCX5mIujGsccbt+2zHhKjC+dI3hDw3qj
HdV6kz24xs5ebdKD8bNZas0PPAtqBOT7j/NV2bYW5pvDcNxtxf7uHQi7j87zbcy/OvZG6PwKr6EX
say80sO2bjuE5HH+M6RwRycRilMih5yCOE/9XY53U6NXsU9eqbX9r18/aHz8TSv+JNKhg/szBfr7
LCUC9flT1NPIfHEOvRBSFBVnXausyoxBagHESJYVkQLZnuqY9pnJC5XNQy/RmvtA8P7S/Ai/4joc
gbeIy+7PQQ0srMvRKBIsX9lTgPzI2VEAawKlVDeK8NP5PPTdpuoygJdIQRPVCdBpveBnyX0Neh/s
wO6mBa2lHxt7NP9ffe3hm6cbt17ivb31oqCUD9cWt7+bg+qUhcxN8J6xqHVzLoiGQb4mznZJ0OJW
lnPHHa4zAW4Uo+N7Xr2aB1KHElMWOioyfhNIKMMouE7he9clWhUDHtEDbgHjfJf5A79WHK853cSA
yr8ZzGLuchYO0Vqju65mATQy4xAhCrTQFApyoYdSTKMRsFYYejLD4lZ7ByUjfvSGm8MoP4YMmU+e
9Co6UDmFk1uSffczjz13eCAAvl4OSg3STCqUTpFlCvpV4QuQiOswLcu9tijjLGaUcjQnip0919J9
j+2ncCwqn/qFfoRCFIeakGn9ZT3gvtrgrMT7GCDZj0KCq3hhJwlkxkySkG4Vgjzy5NRDMM3wYeRO
hdtQRfBF5MRcdOMUler45xi26pJu4E5x2DgLJt53ybAV87ZTuPJLOgdnqWZ7RrEFNDloPlqbimyb
8a6ncMQT8TnVWV7095dT8JqtYE63wbxgZebLSuSIDRea3R0jzWdRqkT4QWkffu0rcUkXMm8LkO9R
71KahFdPf7jOE8EceCtZ8j5JsUwv0v6lp+4b3+L+H2e867YLdKd02bDx9sJoK3oR3O+sxqVzJj9N
XiRDNNxWlkb7kMcec77JoGAxSrNy3mBxjFzd95bP9iGHe9rk6Cf/vMVB53U3WZFQGPxEdMf7QgOg
jm178BZcvLXN9S88Uf6N8gbWxhbNaUwDNpO2wR5whCHI8KZdpwtmWTf9aMiKzQ9+yFFT18KNN6jJ
WONbHDG/RxWW6rdJOhiZ+cCTc2dlAuLOTcfBmcfUGQyNaOxScN+I4KbopdlEoRlWYoh+P4Zofz8N
VY2RnZzY6vngUJQUpTcWRa6Wi9WY2MKf/S1DAp9RCPbNvZM3wRExn2X1dkU/3gNiV0ihVhPcTFR0
q0lSc7QN76O9tkcDtGVKmHqm1g3Rni5UCd8l5cY9saDpn/WfcFQNAY3dGDzN3zkBxlS2NcXQ6WJn
AX4wDlBMTr0XGQ/mrtTYUCxL+P2XTmh20z7O1ajXUW62Y1KB7WGhXw8BRv+elfIGxGuGaB0KZgrT
K4kHCnjz60f7K0oGPJ9/ZP01n0FWZVgj+vzTsvzeejifCugJ85EYqM1Yz8Q2hySvYJnLDlmO3hxf
dGyJ5VuBc8sju5EoPv2HlSx+U3nJiiCj7brYbFP6hw3mERhEmUUsLzvP3TvDRQoO2Y9hGFhrYy9e
3MrO08jOsEN110jmA+5fOj4A+ZdxxlPsHHBpHUaNJcKxcDPj5pI2dJoyCkMmIp5sMZLqdgXkYGq/
I2ItBEGHraOCMYbu0DIx9Pf6RUO912co8GNcBg9U8o/E1q+gaEkP8QwggL9AUeg6I1OFikFiCYih
Zgao1kIpw7pm0Y+IAdZAjHMJspNsRdNpeO2AOnH+aujuq2O2ipY+VWneT4ZCms9ayuYtXZDJ5Qiw
i4/y7Wa0FoYnYjyySQceXaXWd3cpEqSB+r+wOXkJMxM6FdJ2STI5CzScMvQVIVwAbb4mdkjl3zds
0LkL5rT5dI8V6Ez7dXAIUqPiIv215J3kyCEyZUcbTtJ7mfB1V2gXxKKkM/elVOwnu4aS5bvfnV6R
f5d0tR8FB3EEeGJPzhj1mbrSAS77fTX4TCr5tbgSOqaPu7NXCNfgP0k53EGxG1UxxpeagfHSoM2k
4T8MmaHNbtHNHfI9BNABJ+Ypb+sZZXEuFdpK5q3cTWqBhwZvCdyEUVTscZ5PDPq/gUXTGZZbRBWQ
2IVUBmMpBEvvIpQbkncUbRMlX6rVO6M6sMXVfoWmiT59RE59LmeQ3CjaTejyXV2DDjdn3VcoB5C6
i6NOTTpScz3jGm0ZKfsy7+5n2rPV8hQAFAJhFPeZNQEbmok01ulMHrSdP2oCnu9C/OfUgRJs6Fb/
wsy9acb+d31llJv/Awe9IBjEjMrXXOrwTpm5hBaGobkCKgkUrpqPs+MtktsF2OnjahcVvFjtdpx5
3GHp2Agy8M+izshpYNrwMpGO+z80YTx4cdu2IntuWLeKgGLQhuYb3MLsOPTOEluq2awSa7hlWVU6
HcKQhPiKiD2qMmGNrYkh5jWd32NQzMN2uQvVZ6pOu4PLbEm6EQ9kArMZnU0qxfOYt01nvRx/L5nN
mfy4V0BTceYHHz1cnZVJKbHJFct/nBz/vB+ESrtV8g4WpwpgvcUI4a0bRv0aF26e8lhy4UzHucLU
SEiMC1BAubxY10/jLnusfGqiosYbp1dohd99wdlTNiV55t3+ZsqDFH7KO3lZv47rA0vdc7RpZoT5
3uVLaOWpN2J4y7Qu+SaYo6t2l3W/prQPqQGP7Sdk/nUi4N/smCAlYtXYRmyOq72PZ5PNt1UCnfHP
n/3LbxuwImmZf8z8i9QYsixKeeFcWpuDrWAgB0PMYT38F666rle1WBnpTEMuWP2X+od4j+Y1Zq8E
6fSRGT9Wqv+vNskSoxseSWkMLewGYM7LMIv5mO2ZH7mXkiWtfaJh+CkjJBbEa3xTMCHpz9v+BIx+
AFZ0PNxRotoa+SeN2LqptxX9QqK3bXGxrMf1pEgNiQeAQ/ZdH7Z+tgGzsUXvQv4Tms8NyGNI0gxx
vNUwhtOy7U10XpCmm8yvxvkhHEXYCCLXB8p0aSyTijwNpFjDuA0yo6MIZ4y2H04dWgix5jAzEsJ4
Am74YCf1/GIQ1UWX7oRxKqszUnZspxHTH8CGhZXOYWu3tQn4OpagxFlzthQNMtdVMZnS0O65nRxN
2EyFNfCkW+H9TqcP/UIBp34BWwHhvvFXZyAE5qQZkNsM8F9XdGyihYbqpGxYw+QUsX4uDkJv3zpU
kvRPRpOERc7HmcbhYa/dSMB4rgLkQJSviSmC/81mWGYhwLIPnE77ETWpSt/dFXVYeW7FFEAHqxk4
cFexNJchH0lD8zZqgSmuHo0sqSr8LTCs1JKlqfII00SYn5acK3CzY8geu15z+1VZY27AQSYGR3+x
gHGf72V4thwmn6vNYDxXQs0RjF2BY5KVkKZUMIZ7edebC6CCUuZsl4ccLJLGZD96UTgFz9qDfVY3
w1UmIh2+58p5q4vQYpgczjf4sllF3g3i+aQejqsZHtn+wNQjTFJ6GOX6ig4PoZIIYcyEAozseHR7
TklBp5BoE+X3jVONJxj/6ES5OssQgKt81t/Djrff7xGxaBeE9q8sZKEd86LtjMuVEjbYe+M15vNC
5jCYnDJaKtqSNBoL3J0Qe97qm5kZKmlkWNonmR5d9JrT8JxKdC322MpLzGc9l9pAdUjesG3dbQr1
JqmUud00YmSKIcUNPRE61J2Pk2alAJy8+8bonC8URNMoX1iT6Ec8vUXmL6ZFCbQg2HHn2uKCEGe8
MVSM7I1Pgl/RAA+tjs89nCEr2NkprU7naKZ+jr/Ba/wbgi50ojXypnaoERVJyudGK/IqUQ7kw2+v
Mc0Ydt6wvxgzeENHv4WfpAss590D52RYsdLrzFoG4Cx2gbmOiObmMmvKDrBbhC11JnDFhwvUtAr7
rG1rJsNZ8WTD9jGYt51aOysGaKLL1wGdAXCjQMLRN0hryVprsnXBaXbqPyXSWB3iJv47lbCh6lSk
72k4G/cvhQkjqZAGCZQLE1e+5UTsWc342r3b0bCDqWDhrWsw75iLvhtQVaOJnXsFqAgTdPrtv8Nx
AaDtaNlThXl3rGNZRWCYXdxzn8vPK9/O6ACkxHj9foNpvB8UgcU9WYcWjgaGEYALcf4hNzpODpJq
FZptjkhVkbz28zeJevj56sPzgdbHcfrjD1i3waXw6GjKB6e3VqGeEbrCwhQFaN4mB5HeRruFbR7O
6Xfdp/gWVwqBNfDYlCopwg+GQHSpEDi0FsPKfb9OtluI4jk8ZyKVRr4rBi1B+CfVNgM9NSd9NGax
npnKAr2OTgim1rFr4vujvvTYM8ugnXwYeqRs2Xq2DCIF8/FjzfT98qJEVeYzcARz62IkXo5XyquJ
fuvzzcK8l2wTC5OfMFdzByd4ATB0qiS6JR+q9Fam5kN8qQ1wwI5IEV0LcdB8IutCQ7CjNesW2S8Y
0vLDyRrogIR58HAA8c8kURJFw3W9Ybrbe+PoM7zWf7s2WeJcTUqglNW2iRLMkqj7R4UcMxFp5rEp
Dfa3uPUXfiCnuFAJk7qIAVM0GV146DlHWDr8M71Qh5WDWttcKKBMSF0Sd2vXE1WG8fS3Bbg/6CQk
g0EuHxd1+DBiN4yA7G3OahVsjXLQhrR0Y6iGwKKm4dNCmNuMrjY2UC9UyNr+VtAkz9dpjsZUjpIE
zB0wNpcqsEqX3R/6qPn/IcjtoHUybwHzWnLXIpGvcb+r22BljIPn6L3e//Mg0Sej6F0gnL5Agft+
ZxAUBn4AADFweUfrrCDobxjQBpG+ot379haPS5UwGDgNR9Ua5SbVlNCq3YNF1qCd8cfY6UXESk/c
OPN9811oE0ZXtyFtzQiDJZ2PPWAQHAkyo6wNi252QD/udy1XG7l6rCnJQ7UxD+4wqdunJ/y86O/K
w++AH58OaAdwgj24dSNwGKgm8GVa0/WFC7FaaiKEgxgoMeRqjfM/bLP811aO5MBtK56GROOtI4Kp
JtD11CHMbO7FOdC+HY6Q9943ln8RvHVQO7P2MeSSKQFr0AbtC0wdsNg39S81hwvTtjQXjidVAY9o
7nrjeBT5wRH3H8WtuBBG+YH+vWTxdGLcKpTX09Sm5W/nb8PhwBwQSaGqK+08ijg2wRtHvJlMuuGP
fgrkSoSpEs5yyuBA4Ecq8C0p/K35o91wC6JBQvF3ZhzyC1PVLV5aDaC88fdWPaIiOZfJVrUGo2u1
OPEco5uT+GpJrpWCjTuWsY2UEVCtOXi6T1GV2TN9spgqyxCUEwJrkXf1SADu2IZM+69EfiVf6Ep2
beEOGGpCJJKF2MNjjfJUG4ayfNdCYn8YxmdGGe13DkFIGf6yLIm1U7YJBLcH49gVN/MskOn7HGrR
bVuwfDgXpLtZ/gwv3HPsG+9DmbXMrqntCPK7aPOyaa37E70cqk2ZpNw+R3XAVEHCZLmyhoE8sNjI
YLSvlSzqkYsY3nD/aHvtr/jUE/rnG3kNjg2vM6IjrYXpePlMtSfF44IY5Rj49YheTOh/4V9L/yUg
42kVU8V3Z8wYMUZ/Eh7p/SMS3DZjp8aA+MCXtQydxwfQ9DplIFTQ4+BuiyQzuxMq6jKI6Hw6+NTP
cubuiFvQ6YgEZyvPjhqka3JzIo7pHfD9GgnCZWBwPdq0L8Ykw23aBiV7Zp2YvMI9Mt1TZ7+5GP4s
VMRQ/19TG2SZtE4n/ibxh91zbWFG/7uRJKNujS51PnViEX6mxnsJtouJum1QfqmfzwU3qHeLcjJw
leagEjTCWZhI08hYDq3mBBbUXMygk10nACb1ATWD0qYqDF6qZroqHQodzQErUhnMlgBO7BbfZhB6
oBf0XX9WYeEvhskVzn8hUt42aPcfNicYUssh+C40pXslKZVsh/YlA2cDJ8EaJAKXCyjiXCoqI3l3
fB+HrxhKVFZOsinIU2NBOQ8FE9yVSGoe8PmC81A6b1UN7TGMYP6F1xH9iwe6YWpPsk7Doxmi9CqT
WI1fKFCIzRvaEkw8yCgr5oinKxO4aj8HB4RLcb66N23tG8443wgHzDWb1FidRZk+iyrEuwRgqKa6
/RozU6thRURH6Sz2SfelWhRuOfqosRb3szlSqwWkxR4rvstVPTvkdqZvJcFkAOSjly5QdCC19K1e
TzJgdv9KYGlNIhCmh0KFqnYLlf5ufIuCpMnn9vNgReBnRVb8H56vjtzdjKbMOu72wNXsjYVe8htf
yHQtUY+33i+/fEQicKRo0pHnYPxsg/7OHUEmDSQCV5IiZWPOvY1BdKXd9/vFbZHwEFKEKjERXHm4
bMPXN2GF5i4F63SC5S71eeUnx3xP5hKyjlRuJExbe5+alTm2d5+U2Ih+1Sn9pZqFj9P9U0zSmgD0
a4C9kbmwG4RXCz0jJaOBPXvKKiwHDcF5tBC+JZmN8A45/AEqRRRh13gHRbB5k+jycObdrMVwfuJ7
ZaYW8mSPOXkR6B3ruKf5sO9IZmvwa/8SgG6mpgI80vfT7GKIabgMSx5dqTUGRF+6JGkkalaIKdOa
1SCPrasV0ERxE1inFkDzqd8USzPpOuccb34I6B92j1aShXM2G0S3PEpIx7K9y62dw+CewvJQHvkd
B3p7sPMqdIVB1Qhu5cCIJTKm8c+BAluKQAH2NhbgUmYirQA/6jIV8DbbUFCCSHhOMA5MET9hvhyy
impq5hiZdVq5FcmPGHIrkJpYPPEl6cb+LAxHRCI2TO+kDyvaHgV4wgV7BSSI8Hrpv29wDvnIPHQE
/UuiC8Dht6v24j/vMI4G1yda6MXihM8o4jHqxUtRXKwhIrYEXNWPHhYzMNxttZuJ9knnezjs0Zxv
Q5pxmhNOW1pgJWQEcNbnhqqw4k4PZ3XZT6BNN7Hww3LofuMOij0FgUOb5iq+Wu8163+wpAutPkct
RxBt3sswOue0kRdlze4QXY88NJJOzOW2ozGF9eNbnxQKrRyH2YQoIjZy8N3PuQCZ7khiyTfKd7UJ
Nm71876bmkgR5gDPN1qtec0q5LPlLvJBQRMR9lEncarZXk4IiZG5FgLwASJCvrrdTuCZ0tMDG+l4
/tK1Ddvv2tIfjdwnCoy+UCuCC0M15xQGhC0RdSNpi8FtNGNT09+Kj1E+E8PiOwKEXhKq/UJnkdsl
04D4Tvt2OHciW1LfK9MJQ2UQB8zuwypxY3MMqwx2Sg6iDvLCAIjueOZ8DhBTUloDk+LRfj5QsZax
m9e8/7JW175qy5ofG0ZeCcIzbF1cA2ANNodzqA+jqCfont0EpQJR7w3a+HllwFdxLRjIOQU//2wu
H8XmQPhvN+hxaeJgFNw8h58DUm3/Mt3BLz1K0QKLsAg9xULe/fdpY4jS0KgVo9BNcjv0UvFMbOb6
lsGvIJHRT70zwDZST6dHlbm3pDytYE8DGrIwPkDUZn0GxNdApd7q3tWeZk50MAJZVagd1GLIp5Jn
aV7UZm6V8iDZ4cgayyn/sHo/2lmmBQHipTqw6RMQQ9NXGIEdSYpQnck7dSVoSCjQlm5RaceHppzq
4BCxZtCVTQl/xuBbOAZj27ZolhufSE/0Rdl4d4Ug4Qswigrl9kILr9NCyMLWzRLxXKrFw3jRJnw6
R7waRAHfGxWzvM8zUBhdwoF+JNzcf0MtMhZsb23tgzFP/NG6F3q6+FEFSLWQYZuEhxG0GmaELC69
rxnePCFWtmhqPIupZkit8yhq2LyrZSKFEexo3uqyLYGXe2mXNLDxChMRo3TENDz5DChQmcE4AU6k
fshFyl4lH41V3t9Kn8p7Srz2HJGx47udXV33lvQV/KLfKOtlrzhp9Xf5GXO1Kxx7QK3IiPFJ2rpb
iEu4lMZY0zxUE9SAUKLeoRu0gXk5l2YrlWKV3R+0m3+xadpDhkQVfo7NR1uocS490m0LeIxLaA0i
Er8xFekz99EQV+77WV1vll0safBonYTFt0kuem8F87kW7B+6wCQhacAJDpcPNEntzEmjvuzhwjq8
tv7JrCqYudPLReM/ncP0pGE0Kor/6+EIBRW1fAvVOhuJn4TyhGZjZg1ogWBhyYvdnNkUMC94fWFy
sDttWSVD2vHHbcEWq7lql8IL6LLJdFYsju9LNdJ1xNQpQFzH+ABRGzdovQ+GirkMOVaxcTYIk0NT
wbd5Pf1ssIML1bn68ixMrhewTTVd8fHhXpzr6M6M2LFAZ5SZwZXM/RRW4OvJnXlp1FODgNJxyZjN
RjkeLwqKtoszUEggGnXpFl1VAuuHXrlLyBRQwypPGvf8vKdXEV5yIBFWY+c2vIC1C3MPArpV66vz
1KEPD0OCVTtkIjtRNFyOi4pHJ6FNOnU+rmy6P17D7BDsr4DEvstmiih1kO2QoQGwDiesgrc02l7A
PfHMqbcXYMbagUgGEJrq0BtIJWvNn/cT4SSf4vvLtTLQlTO/NXF4JqjEnsiFJUdlm5vTRj0x66BX
/smyW8zvOklFzZ2lv/DQA+pUvlQqpeVXS5F/rfyYYq65d2lqQhM3eLBVG4gRAB+9eqtLvMDtrB+c
zU9jFFDsgXKxDRneeXS+X9miiJpo2vClV7d7wOhbTFCB+6+fIbPs9mmUFUfbOmnuVokedIyqS7Yo
I6/QPoSiSIcqrSYDEe8LrTiJY6dvKXYatGMjCGePHE4GinZ8KCQKdOxepP3QHCbABVSMqYb8Klq9
FCwteEJjVyHelmSaIYedhPz4zIMXcOkgoxfMskjGgpjCyySR180S0brIl9SIitWG2IWKHbCiAoGZ
jPXaV0D0r35T+bhsnDkjbnxQX43SV44JQv7M1PBdbQARzCCoVx9fIoEHD/8tiVBJHlvKy84LhNfP
PUUgsT45t6iUnKH1tnQSuCELrg2gc6ToieEm7iG2BvAWuKc/4zUObK4cBiOH2DUWWmI7+PiHo/Ko
KfT1soWxVpMEjxNjPKFgVSyyL70Vt8G2IH7Ru4GwKK049RPMFJzxk93W1rnQ7VK4RlUFnsh8+liy
w+Fn26uD9UNJiMO9xwHXIVhqk7z6w1JsP5pl9WlwEEh4ovZeV83GOw31uMLdGyC08RILX6g79aUv
TFxrmFBQEtyq9mTFa+7/2VxXk50zbUgpBSBFmm/dUxnj+XDMRbZXRB51T22eAvicypViCNwWjemE
RR1XePLsArl6xspaAl6Slqw71Xc1TfV0FO7G/jHD30EGNkzdmLk+qwBfG4xhXNEDwQ6GyiteJskP
xc8ov+UQyihfSFDJIWIvghsNfV9iSpaPxVjlH945iOWZHZXwZoBuiTvxnb4GpODBN1oH+CnIV+ax
XcqcUfmtXSfNNNUXCZd0ck9CX2P28lPUoJsPMecky424J6FCKNRLt0IMzQNSbvM74Rz9ZqBSbbgO
3Tajs3MFAhyaDn6TgUrWdIGPz2igc3PUJ+AaeoSJ15n8mwAyT++K9TNcjC7jLj0DS7uf2ajzH6ir
O5Y5IdaOeW1dPUEsfXvc+tqtEbCpEMubIl8nfPRNVW73HB181J79z0qMNxTBbI2ywBtEd50ZSfML
sIWxhLSLvziA6zeT3VpJkb/Qy/7E3joR3oImTrUjxFv3cgSuBYwvD2r3oU8++p9tn8WPoz8KSqt4
DoZvzRHp5tUmHG86nVcD++4MPzMq2OoCM69D3xko6qZbBiPfBK6cxb5jAeeF//Is6T4tLRI1kmcd
DrsF0r4GMyOpB6os/F+ft0/nSJrHE4mL8/I8lY5GLN4i/4mUt/5vx4gnA6WI3gosPOrDgnj6NZN2
2XWRJ0lQk+MQZLgVG58IsQ3KT9FSW0KNCE0sZSjRyiRxpq7FLigssEZsTprifLyfCou4hOdHvT2K
WDFtLpqxnjpodnzKAV3Zn4Exq0N0BaDZsGuuoQekGxPqG5nh8DmNL2qLWN6Mu9St3Bc5sjGgbof0
dKBr/JjAgeY30LVX+yOR/6Cj08CJ7bK6eoYD2mHuKPuDko+WomBOXGBCLsmgm9GyfRsTpQJxKxNS
DXW7+HCU51x8BCE2eNyUu5xHHnYPwknmrNgaL1O7G5vFJwQ6XmmNgH9fU55LNLcKMdjUa9tDAhY2
lnb/xy0u+9LGVmj0YSEV/3W6dJHbgqZ6zT1usAuMFhYX3InJLinhIjbmbbhCf6OutXQFMMAhpo2y
SVN+YfouiVPoD7One2MnOUat0G5SVt1P+mWqTdBdV3UHn9B69w5ZQcorFdyggaZX1u8ABY4gfxfz
xAcEUsRN1rUFShz29c3mnDneCkd+DcBhTia1vbLggw2wGAuF33rE1Kt5He+xsl99hMc2/WtgqUJp
gU1bYKoVkN8AomZfHN/GDa4+eBisx1ixf0OMCcP5mEIMu03pkzRXgxELM2fAV0CSg9oY/+YYCSb9
gzBT5g6S7BV+6r3bY4dblzeBXVDutkwTXA7V5Dx/fMS7SlrLKcvnyvLMtAqrX3WiB1z447vuzkiN
2k3Phb3unx4SOVWaqKlVxaFmzzjgCWTw7TjP8NggtdOSa7r11I7F1UgJw/Rnu9itKlF/hkUmCUfq
vGXmtNATT8gUbqRGcx5EqFbvMxQhjLXCY6GDp3LeWqWfoYjjKAMKIWxtJbr0nb4T8DpM7fKCJs5V
dV34m1X+IP4Bp4mK1/MGrmTcEmwBWL5ZRaWXSkwEo0/u7bwcGOjs6cYnyziZu0hoGtowRDWOgk4y
mIEGlRExdsWC3zyR5NbYnUNhN6nZutbT8Jxmv2OExTtHtaD7zt6z0FlMj8jSiYx4+bUTURVB3LNq
QtKQzkdGNneZWdz6tNH4XO4EDOkjpbqGL8anC4SsElSRF4SySbeNYhlE029W70EBIt73xKtM7Dyr
y37od2FeKfhfoesGSzCnNVK3QiBWtRPnQUOqBGvDHwwIcak1IqgiAqlo5hMG7/kDbySzVtwVHxcz
8kSKHRl6ZWe9gJYfOvnX2zHHo52nJQpbIMklaCcCy0TLZhMfyYhuitKRt9f0GXvvcjYLs7eUb1lW
CjDWVC3GNeXb1w7Iiw8QTaSkM8Rnu83bzRhVZM8bh9Yq7MJLmycHIsleItd8Ncr0IVOUNvBjZTmJ
cfdqdh9Nzpt05BiOsjq4bgfROhpI3P1MMJZPRvu99pWSvTDlCPSr4P199rILggh2tu4H9o2cQvLY
6LJYFlpY5gbTgu1SSObvsjFNPjB/t8EwfCVg7w5Q1Wiii4aUJYywQRDC7dbMe+kcGh4XsGkkuxVQ
a+y24mY2dMmg2m/rQd/6W1uY5ipJjCxc2kvwgl4bE7hhaZuQpm6aUM8iqiXqgvYxj6X4hPyCFq5R
zzX5pYY5NfILByXx/aT6Jdrsh5vk+V4JUYw5JqFSYgQ6rLLRNETeO0CI+FL4g4f7IQrpDdkTwVN5
QOril7YNHipsnYDbt0YC88WYf3ZGvmAVW8RQyEnGb3NnqsQlEVjGEKlNq1m2HXumq0q7dYfI1SGL
iU8VSkAQe0I/b/Ioe3YfsaHFbajZnIH3PYGnDT8/X4prBBwa8vxQqE1eOq2E5D8qj6p+RnAd1uYd
1tANlMTEsQag54zwWRKzFczQ8V3vjcqxrBjaGs4GjtpJ4LIHtVlSYNxpmmcmbZW05BH2IfndMd60
WY5lPdKmIEW9Z6xZWfA/2Pa5pEI2LZdtyH6NzvpUOMMcGmcc5m3x+XROVm+nb/4bEprMdywilkmE
ZPBRDL0nsXmMO1+0rnWIo13T7d++jmQ94f2VYbnRRMUPbi7n08NZv2sUhnfyhVeGCh1BxuUwftBC
6BQlzoEfVCHHkvI7m1gCwxRBOfT1Hkc3nU88VPfeOJCmLzRFh5esiRS8mCfJwCv2HnDRy7xc40Kn
1wLbMO7S7H8IBJBSjqlihGuNWp+gqFd4MiugL+ZXnN5b8vaonhRNS1HhiZ/RNgov7jWbiO+4aO4/
+Ks5atAm3WOP27uNE46QDtBEUQRIXbfpXE/kf+YaLFd2pT/g0U+Ootk7DYBgQgyfcuZyROMOo0ol
goSmQObUW5OB86q+o2kzCKfpYkDTix4dXa70tHQQWpcua8LC6jszI4l+/23e9iw4gZUhArv4B3mZ
2cl9SAndKq2e+7WKsk1OOxHC37SVjJ0N+9weKcvI4AB1CTsHLZ6LcR5+t+Zb5FelPbJVQhxTWtvP
tw3aL0HplbsACJj3yngfhThrLwC3AE/FQay/DqzkmvY8MFnCviSc/bO6cbWYh88IIe8dtZN+Wchf
2zMMfHUiP++TQXZFndWe0lubDTcZMdAKpQl8vxi/in1YraFL4O1SDAKpXEw6K7L+EUb2heq38acH
myogo+4I9J3fLJx9njeIzR2zMtVelpX4McHyZdUt5/pBUYE55D4o8mHW7lDaQG52/5XL0A/MfIbH
+/OC5QxZsJeslMK0aK9NJTOBdfa2yf1yMePQC/iwtsu3QqyCX4vtiPsYfG0wHrd8bBNB5jKzMyeD
WZ/LgF2o98AidMSeDg8omMSFjFcghR1U8xm49Eze4mQoFo1JBAWxU+fKol9Lz9y3Il66BG0GSJWs
rTZmOM6PN7u321l4tnau+lbjxusxrP0oNZqdK7+q12Zq3ur6GvH9yDCs13afAwWiTqKih4J4p0X2
FBw3shR8RntHwHPHMYEZJUZMaCZR6LbLtTjLAiOclxsy/l/gXbkh5vt436bKYq0LnS+B//rZ1iL0
TqJqq3OwP0zvcHY86vVsUDGC5T3oU6x9OJOdFa5hWANulNgSBJ7G7RDWewqUn7hs7zrtcjQqFdWE
H6EBjC8wblJaZUIIc4yabg3J8PgDP8WYIcIAdPcSFLhBV3Z+DtOd3ZjtYgpfRwi4nG2UplCF4+jd
nS48aQkh9GbaBlz2KARLayaBzrgoiAT4SpUDBtW8C9ctNPq2iKmz/+NyLlGt3F6ZCcj7y5b2rLJe
T67wJmNYtn3+9NHa4fNtqbVvk/AYxHKffySJO/A0I8EYgz+bbMsv25TB0MnjhCoH0CnTGaOx/8qS
EsNQ8y6rIxL4+O9dNytinJcL43XDTLs3jP1m/Wj6CqaswH4JlIHhjv0mpZ0qyP104u0R1YWtEcve
/dJRoEcMohO8+SxrCLjMO7zw+ZjXWR3MVUg9OxEcM7rf0PS2ueuMRc9k/UgvBTOrLKSvAaUT8vEQ
nkHkvjMF6aM1nB96a2PowCt+SfLh21P1S7cdmZO77Ie/aksclZjT+ADGoJiQzeuZmewgTLw7p5cP
B4tuRqnTCRQbTkz99oDNvCvgj+VvRRemaIeEIq5nIqjsWh/Dc/IobTsjR7P1jZzjxSKxbrbulwzR
APMjgxe14NPRrYymL1WYbPjXrNJr62EUcYJCj/KU+zr/yT/Aia5S4OKiygZRZRj/VT7BW5Z+ZpTV
cCmmSNd2hInsFWFXCCaXDifqtsUOWlZWLevZnSlI0CNsirPLXx8SPksSGcq1WKbphA1G5VLYosOo
G5vcIBS8I/ZYKjWCC1CAXnnLkCHzApGiMBURGrjX20SNpuHW49HSfCQM82WYkZdSIsi0S+ZMV5s0
Jo+ka9izHXFR5G/7ht55vPJSnD7y09Odv1CESQpZVkPyX/ZAOEEkpdpmRHXEZuqY/Y7we1oJnCh/
1hfWfGZxTCzEdja3lA5lYhNLil4ceGJKF1BuVMySlQbEL9CM2/jiZV1Qf2VoN7Ws3VvF0LCuL1JV
WdDXAxWPwOrOK3p/t1bPkC/OFk05pmzf0lLuy1o+/Iyb5Pm/9s6VcI+pqwuSg8Hqjnz8NuLO0m3U
yKxS9jj36Vc8j1mXo89Q+8KTxTapyXBB/pjyebduPvy2sTYRhOMorVu0p4PVrhI3grnJEdAQVP78
xGpK3+j5q+LQhwGgL8i0yH6PvSxZB7PrLSIqjiL7NU+zWJlWUgjAwBBlx8jv86C2pJdxir3VJf/m
QJ16ZHwyAg2PkR2S3LJCvt110tSI2PIX85lq8+AmuGSe8mD0//Ci9s2u7yJ2DrQKvmVcLOWbtzW6
ualehFDyhdOcfgmUdTwGgnHMG0Lv/tHLfdvEctAJoJSp/XCLIJME641rolak3RYKtS5Ea98D1P50
WsrfMYGYJahtNjveXl/Yfp8Rx8DqvCPJvKgOlVQhY4WnsIV3GK4kjIMe5COIxXP6WVy8cPQ+4Wzw
tgJ2sP8vcULPdChIDG3bPUC0FH/grMtpUvtHqm89UW5i8/iosJzNvtOuOehRL6l++nfqULI5CFZi
4SUBrjwMFBJtH83BkiQcxGcSjeTBhS1RgNmAC36VMKfP2VIhPVp4verGYyIq1Ktd7DzulrpCGyA+
xjcs7K3YqxDKRku7Zvqake1X3q2CG2IxRV6ozM3f0JX/cKcNKKREGKweatlN/4aU8pU8+oAEXobY
AK9xJuvw87xeUBcHu3BlTtwlimbm6oj01wCarHfWA3tRbmp3LtQQM4/QU+DfNnj2DuS2oy3+FK/E
s3ta/u0f09f1rIrQcyOmKvFN3Kp77kFfMmIRwd9qrZMRPAzrXZQVFOCOOU8QZ94gZ1lQYuoQn4fK
XHiMLR44n04h5H4ypgHCby+1/zP+rhP3CqpM+3aLQ2a2QrFbrXRrxTk7HnVlprGfGQqGBZfiL7+D
goIJFkW2pJeR6+6R72Q4mP/n1GG5N2MzhS7B4OiCTSJsgrPljVr5v5RBJYW9iqvGy8ZphzhrEkut
RP1LNd1DEnleEvPc+hGMFKNd+qUAaCMVMnzHKduwDf2torcwxGhN81dvegi4D/XLaOK6OrG3ah6m
zrH3XcMMHYFZzzCkCMYxUGJqumCXGg4nrNgu1BkXzSX81NwKFLSp3bb6W8N7PbboL3HXTTVev5ix
4seqLS4QXOJYIgVlgZmxOV0V6qHX4FfaqrraPyj62kaHEzKy6wlMIaM+c5m+ui/dO8EDmfXrWVOf
Cg73q8TrzemQvVjevLhb36SucklgF3q4s3c6D49zUfCy2+qx8kJaQXN61l12WSuwZZjdYXf7H+UE
8/vwbXFUpj+f7+9JgOMay84Ywz9W2LamCErtATOqbuEfPkUdCWjyShaOp94/s3NYFWjaGdocw40b
qEoi+RDicgrsYNv3FH2OeEZOnv6eIk5K/mC5WOkjQyDxyxq7XqylDKW6UIdyjvhJENQPgo7/LyXY
88TyCBCEN8VIhvCD7++oSZrWiO4ZDLsxCnDBGPrbk73hJw69+T9MbyP0zi65LG8xZiUILvhhFXzJ
MsxAwspkswTFvFZa7okphLfwUXl/XzhDzynAGnbjctJFyQA3e0ADcAvC0XoRtqY3sQi2FYwOyiYl
y6nOZusiE4yo/Q9jCn00m1tCpwboA0tGMEAeUvW7Zzm7l42sUIBlZwa0Mu5nG/+ZLktbi0re9JUM
1DXOdnlyy92s495kfoXYZtgC3fEIiT8EC3SFPuFndnG3NPVAjmHjk9EN3mglJP3tGeVdG0HhuAbp
SE81u9CpeaJGct3lD3G/tEzKgPOLC0Qjccd7oZZ4WJ/hrKpLClQXCpX2GVPpZKRuivd7R7RuPs0Z
adDosMvkmvFYTVqlXxOTp2q0JOyyfOCe8nOG/rHi9BVWVEhQxpzMRv3N5P1WvJr7OEnQsx+4ebk5
YpMblYFF9O4l7PNK/PyQnXxEoXqf2NFdeEO0J5/eo+UxLfP1dW8UszzkgMh5A/ILb9VbIkPkfhZf
IU9wCFpYhfaS/7DzUubJT0rh/u6R7PBP6npm75oIsNeOQa9HeOFZZxvYp1Ed6cni8XvVI472nxjJ
HEjfkDSKQ4ff9XDMi+twld8vPzD0pn+8GCUg+KFotnD02JqsBd//9VqCfFPfffdDkqTvDjvFmsmE
6H8QvEL5qvGC0QCBUnvxXE+u2DAggJ4RkKRUNOq7Ule3z07G/NQjLvy8+8o3VVCAbhsmHMPtefHl
Kn+bvJi9447b2HcMw1AKsytBvzt1ZGcmvYfytbvxEJrNAGNzfkPEQj8WTTdEOyebnqLBCU0+MyRR
3ebWQtXqL9Z6Tv6QxiBfJ2aLhGjCmZbCwuFKRbEmet8ySAMFRR8q+udaFPl06NcY4Xa7N4tdOcHE
JiP4lkTW7HwT+GND0Lktk2efwmdYUR6YUPuXVzivI7c6LZLLjmT40HYdhvSustb3S2kzyhE3fz8D
hLX0L8rIj8j1fqtHdfYTgfcXYPgArNEUSBLSiYoTXT2MkEJ98BSbDRjtxtSqh/scVg1xcZOdQeE1
AGLXXDlbIqtQJwy4S9+uD3ekQmX0zt9uJocdK2o4Rx7GBDaVflyQaSGtiB9GYfzUjzuXtnRhJ6Xe
BRu4KIUWzdAvh39TDMBQs6S5GE5oOX2F5p/Y1Z1Q7fdG+Y5ME+JInU5UFlKGU7btwVD1St1KpnlD
8MLjsHlWnrHKKgxvyRjWRbmRqHoDDnrVbPkG8uWHyFrcPULolRkrZI3ikQLNhTypmFdwrljOphUi
zhdzdCzYJ007uPigEU6WCwTc6Vmi5PLj/gjaep6ODJx5qZVWEnCNwiVKcwPP1+PYIy6wnOe+oDtn
fNMXDagG5sa2zM/LO9HWTYDy8DtrKMidGEBHiy44BA1B9IaogsfX59ML4BD7prTbJmstmtUdYaqR
0XTPU0CKtHOcLVHrloWyZokjpvRnHigYk0m05Uz57tZ8FX4HkcwudxCU+P8NJhCtQgQP+lLV+2al
1Gr8VFQtGQs2PFlG9OF2B41rWvhupc2Pbqk3hSKGzBd4jFGfzFWHDwgKhJlh3dUEC0iw2EMko9EB
tB33k3QoV4mhgDGHxVgnkLs9dk9huRNE58ob8E5x5qhP46AIxMtKe+UJ9ZIT94tTxAlRiIX8xIJV
1bQwM8LepwQaQIwSSQQ/D0pt9Grtrc+J8wrSGOaIw0StTWGF3L67fARC+TLo4bXY8cfuTz/o91bh
46rp7UqPCAWuGJFIBHSk2SFm60j+7kUBnj6aoue6GotjkaPdMBP2ymy3H+hvySPAPew/S9bMiEoj
e7Tti/rtSZccl7P3zVM5x1tT4XHgH3Nxs+xHSw3+mRFtku8BsdPeePydwB/TtgCvYxeTBx5+9y19
MIW5TvsZQPICWk+WUedHMTCB3v1VHiWa2bmN7LF/D+nZQtLFok9uL/511fJuBPIRumfFTRGK1se1
0wbqyn77+9c0G9nt42ID/EZORgJjqyY5s7X6pFkjLg8Rfz7e2YxUkXj6uU60K28/8+1VAw8H8Igb
m1xIZYdyHFB+6tZWPEuUuR7vMpEj6Vgh/a+Mx4IdYks3iPtK+uvfixWv1fCouPxh6JpXuxu25kSr
p4eIWCUHjZEKNYrM6eZ5crQdh6ACdhpbT0s5TOcL8UD9+xWXuibbrrLXaaS+0Bq8/l3gNUn/0C9d
eWoQpImGFeMnQtArynFLS7inWq7dSrtwu+U2K8Bu9Q/d4FNLDG9GbkY8ngOWIgd37Oe+k4DNTCju
6bMmOGULfnqDWwjM/FCvbWui5lETVOgk0MerQVIor/5Q/5P0xbN7B7tDZ8uGvVqf+BGsJoGcvwPG
RwTHkM9wj3l6FBNGiLBevakQlSgFnEmPrTK+dlAKhs/X/8m4q4jy0F9/6JVpFFNBBLWr9d9JivUp
8yhpIQ9Nijej9e7goGLiJ6MYJaifqwCrR1AI03ILH3QzGvf3APBbB0sxRl0FrRbHX2Zmj9Qdp737
jN/jT3hArAAPhi4MHlTghzkJwJDSms+PZjTmOdOq7eifv3pHYSxKxhO04c9bqDhIIqhl/C6SyRfI
q1d0q+1PhgIEiG+Ubr92LwmX4P9KqZ9iIgabwOIvX2kwpi7talVRi2wtPxE8leC2z13ebE+riUWb
5ea/QhmbK4OomSm5xFo/zhhOB3vkPcnJRWha6UnvqNZi8kg31DlAdXVBpUQ9nSwf0Mb1xAsIOp32
Mxi8q0/3fm7omkrmMKfcbvjyRgF68jNeOWguOkvV9gvmAJyVGCgxUgSlm8Zjr5bIvlEBduVgpv4a
ZpTX0TcoIeoQ8deORPWCUJV7AH0orRw1p7XJUkHd3jIIRdjF+dZyy6Kmef8Ltj+bfpmAKiTMt5cj
2e+4xHeSIPr8G8QKFoRvbYR5e/XwI/KRcbQU0abA/eE6UxGJca7wbjaLauSXsBEgvY2948aWVsAF
NGSyf/BzCGHkKSM7hDQ2akVMEtkiLPRBWuUkzkX7/7dcnaM8TZKp1DIlIBBL+efyJPrUUfjrJMrG
MZH6k/e35fvwwZFDYx0H8IrXzEzMME6xGZdMaTzZkxZ0I/aGnIOiBCNal4uhrbNvgD/A561Be6XX
gf1GHFUs8HRfDouOc+JqPyIoDBFUu8cNuuQY/hINDqRMvFJbGxvpO2heq8KthvdlSeGsJE9nbzos
SlF788VxwwqUZXIPcd6GtmS+BMRk90rj+62K4x5JBZl8NRY5cWnk/0vgih4FFW6vZM/07bnG5srj
F+fxTKAFWg4uAga0/LnnxhuqzEqUl8cnEY/ofqmHUApe7gJBGlpI2M+fjiHn7K+fIFdn6ObTewci
KJXJIhM6BOtCBjF1d37XzqwO/eMRD77PHS4J1lT7rrFIppLoOkco2mjeWyjqVABn22yUJf/rFuZ/
8UeBWOOkkvoZfjzEOdP+8oBLM4VjRpLxfItUoSO+rUfsJW6ICaMvho8basMTf+HVO0mK17PEKo4c
qd++gfJnbzAnBIh9lM+AacSOrekH8o2OdN3L8rzTfjwYqwAP8IbXnDUxeFnyfe8YQ55/FzwrYig5
KNrB9zlU8Syb4nXHsmXGQBCzDTp/KR+XncWseKkOuK/a2ojzonwZiO7Iz6S2NnVGiOQXpGrLSMFk
Yt98KijuIw8MOJ+hMBpfOtmciAAjCZVfBYy6cv7AN6j8Opdy9TtXuLKOEJkjuxLhrhBKHic2imQP
jgUzLZNjI0Tt7BkPkJK81hAPrKWP+NDvhx6UjrOJFc3iMe9DWF9eWWJdmja1VthiTFBoPY4+E0X4
vVTsflndUBa6nwguM0/+gffij/r1t5lRnrFa6Mya2r+AHbw/mGM9bCET10elZ6KfAHOuoN3lde2j
TRfpXn5CFOX+HpypqBhBi8v50GZecDollUoTJpQdQ0NRaGuSZWnkrhxDls79guI99u3mXbXw1CS5
xG/OKqHxZUiF9moBkEqg5g0HDTV1fyrmx/KZ0i8CD9g7tJa0NQaemw4awc2Qt4yo2gnVUvsr1NY4
Ytmnut4bncTkCEf8pDY9MfsHGkmbMuaXbveLXZXdayO9BoCXJnB6JJotSvINGROeDn/PvfM1W9GE
AN531enkhDevb7LwwuXkErDO1h2CCbspCV9ovW9tepLNGi9TVV+jZedM2jQTjZXpeaRJTlAm5Gmx
obg23lmt1H5LBipMOb2eU7K/GDTvatSDLki7hXb3hkME6/E0T+vc0E4dywszT3GRzIQdyc+Xv1cP
J7NGVw/oQmZp1PEdg8vcH0rsQBYKw1wEc+/5Pym2BSDSQoUWMpkTawkJ3dpLJwjvuav54+m4CqJ3
fStFJ/qjbsjE5rMHzJXT4wCDp3Tt8G/+cggwtfb46IFHu/OGRtYrRH1s5OtehhEeJrfohu3Pwpu6
2W6XtTwGADL4clegsJonznti52aMxTS4okINIZJJBHtWpGFbs03nwO19jRYSU9kZSlEA0oIjKDwg
2XaOcT0zY2aVA1UeGvXGsQHQoNL6811QHhQQ5OwOSYfZw2rJTcjm4A4caww3hn0RIry1vtF+rw3A
LMvu3+mhpaRsqx5QqxzhEh8rsh8r3ABfs7kPtECKF3mHvMpuZXtc88QRGF2vgFjPwI7JaNTzKQtS
UN4S7QKp2mGjHRyzGcTSDi/ntIW3QiWvi7djQt6zqGFC1g/LqwEJxXaAioXHqN49TkCGPASnp3nl
9NMOSiS27OzK7MCa7jokIXuaKDJBf46xQ1Uh47/nPs8KNI+3ApDfgV+J2dklQe+x6Vq4jbqpTUBg
3bX9jg3HBS9Pw0b3Lz/10ixxgSlFPZkFZdtvxomOBs8ehQsXHJMEYc32dh4vWdPayBYVO4tOC2QL
e8MmxEt5A6oWFWqfZRgV7E3X0UO9LJvcMoT/AJUPOZVPY9hRzkJHTMxhRBD3we/9JQRbns3mUVxE
NiFeaptDdZdxhEq6T6jzEm8hZbjU7czqcRKEzPO7O29Z8fOadfp6AHqtNm3Aw+vvjh0jE+09OAxW
fAHxqBTrVA7CP1rF5Sw/Tb2iueOyJ9mLRcmfh5TTMWRIlvZ/+lIQyKksQUv/R6ksurMykaixqH0d
wcjYLJ/Zk+iSMRceQs94Jz7p60UdqKXy/O9H7+MxUX+LJR0kMeu2JcPYXHE5E1FKfbf765uq3no0
Ssq4DTJfYMwBI+oPSsDVlAAqFfo2VsPeoySYPA0uJmliEpRL7WqIK4y+G7xnJFX5DFI3TrM+AjOR
pQn9fP68z2uVCiIc6jIyUtgnpCvrGyFbJ33LNQ3v1oEYI2HPbT7foqZwWHBUR8P1pUmNAUqMf9d5
bmXd6dpwxuPWInum6aUiv3+fVLYEtrDa957BKXoJEFsmMZ04OqqwaHbMX4wUIC3ePOpSFx1rwj/k
6VSdvLktXbek5Mzg2qrMVbLQRZ4DHOQvYb0SLkyi4HOcigZ5oG7m6SMpCvV9xyGPd1LWcw2B61NW
L/uSqQXjNGmZUO3bda3ue+cdno5Qvvsk+P0Non85czSDWhBoBeZb/tLK335hOX6BkmNUsYcDur4K
yMdvcNBgLYQj0eojTIdMFXLorbvnMX6r026oyUxCgylYrigaPW53pStwWK4scuYUiV7BuU/AAQCL
3U6Wl/z+D1TO/5ZVuwVkw3RlQDoplkp4F9UI85N6EJLOzCLByrLKZYpUOEIhjziE6FRo1Ok1Rm/4
bebKdLbliqHTwUcwW3QuqFqI33tGii44L65AuEuQAcK8njudgG3+XaWgStXFHXC+XjZkeej8VqJf
OM5PuVTPn78Bo40JGqGYICyJevERP3d9Ywd8OHx/8hPMPBAHFs6brQxZOkZ65IwayrnyCpQ9+nod
dLPi4IDdq718VloMTJ9DNBhRpKrFPZNtGcHRSSMAkpOazfq1YyePEhabn/ePhHXcN2Y88KYHD4Hu
5c0a+IrvS6TxAhobMVmkDDXBPsO1vYWnw+FuzPlBZoxtLnju+cVbr6AE0xhMGGirHQkuAV9JR6Lg
TrT+DaBB081dCMV2CtmDlF49s2mRFHMCnwjxOCrwwcDASeALSYWMyGYi1mUhbCsiXV7YVbMR1Xo6
zbvLnzmUvvsN6zn+sZhQsDEMSBOJMmddgLS7MIiCoTaddGQzk4fJPOCt5yvj23+ILyqFmAPZTbyA
uygcWUmodJavuotVfhNJFsBt7zSRhzxCqW3Y44hV7oWb0S9zX+aGF02pJGxpJSgyVArXKDG0oUyq
AAm1GMbKS4k9MBKcxuP/aJGhK5tmzBFx/BDJyiVtPvtK3g4HVuO/GOkwJlIPxG0vmbrQjg5hmcDF
GcTvjkD6G8tx9GppDS5OMs7H5z8SPjzcmABZjArAkcmmQ/jsK1qw7Q/C6Ss7qSRt9e4itQ2PbTa9
oyxllRWaan+oijhgujdvi8qhrMcpEtgKiqSdr8p/Sx0XqWk66X6gHRAKgYRQEYbeJoeevBwnsEvq
5ZfAESA/7EsMsrLaxCCPEsNqwWQknPVeADvpWQfeVQqccEKSXJ+28YjPSPtg9ckAiKIHg5uuw3Xd
09lzO5CoMgb5XqHt+h1GXSMhm3dGUi0LbNh/DSZ61QyC3gcwg9Cl4VP3c6Lw5rwuEL9oBZLb3pCU
WIGbRTbsfLRVEnoIet13obW1kOHtkY3x0wpb02gqm5/elRRO+IlYX7/xVUh+0WAJW50X0GVHvxVA
MNzU2d4GigfZ+cbIVTPlxxdrbsVZoSLCz5EaO8QKTA0ss6vBd2GG6abJDkvsc2+/5AijYk+Ofqm4
5avZmgeeMYq38Miu9afp6v7iAtQoX9THfUpsNOpqXmRN4B7nLwYkRe/FIetkusSTa6++lRcSUyf8
XA7y4PslMQMKgHXqzuugQvGxwwUezwNPG3OuKievKQXx6Gn6G0sVBrMl3731DcD0xQ6SRAx1+DBb
xtu4hamcgpqpPIfMkt0d4l6HD5A3lqjziChovCqiY+D/jOtY5kcPKfvgILRz7a268GYPGhrlI2xj
plI7Nm3dgrLw7POX7Za/VpNdB8z5J7ccdIY/ZBVsgm7+xb6iA+frLTJ46XqogLwpa5TV2UyLK7Z4
FxmG6B5hMCtVXZh3i8ghyspSMN9J2ro37C15NDplULr5VTE372n0QMDwc/Y4I0vQR+w2JWwIDPuZ
e0dzwKtyLDe0JeOgtcBo+yApJTpBP5kO/AqDbQnCauCZG2qer06CwUlHTva5E48QKX7a4C/AFdF7
82W62Obq40H2kwbh1UTgHe8sBk6aZ8y95frCBYXKsjCNwvaxiAjWr1TXSqW6vTR8N9h8BDy0lWar
MeyAZyunZ84qBLiEPLQdV6XtVD+DxmXwldmV3XnQHgfYFBTDhuRqtwvPvmwKSqeR77KEKKs0v/sD
VnRjk4FC9xgNg7uBJdglH8rXHzbvetqv9rf7k7vl5Jl1nHi4yjJQMHcVo6HEIw3+dU1H486Ov4hZ
GpldSABqC2JqaGzU7VgQQ4gDQSViSEZTA/ylg4mZg+sNdcVZ+xGSH6GIXRebGlnf1bDO1h7xwOxS
VDvR8iqvQAp8u8MKBSa2Ry5MmAYF+ZXkQaX2/vWe+CoLQ/Duv1iCmCrV2/Lx5a2vN+GFB42tVltH
tfTjdGTM+P6MEB9HRMeDbyqw//089ocQz8i6AsZ846VWLsc7ZnB/MXRJTn/O3dpDFZQp0+jyLDK9
sW/GvNiibVYWOr0yn75QX5+sJSZqaU9pgnalac5x8MdrSepaU+XqNjXzHRGuG7V5W7w0ZgfoOOH2
xXohpvUJBNRGGFFR35NH0xLUSNzNE7zh1ErolHi2mY2P/CskWeWRJ4M8r2y22oM/y397VVDy6SZZ
VKkSQE1tXmzzW43FUtFCtBTIwY/JISNngAl+VVmsZjDeH399g3kuRci/yAWBPQA4Sp6rvEf3ni2s
MrPHXmRgenWRfUKS0D5/P37lv6N0nYxlNCTpbAe9Tk0BdmbHeSKguwNZPfVO+Kc0pxbCuBxqZPmp
A7ieA0DNGRrrfpww6R4AgkHl0snGFS8Ay9xZuC8PGHAs9VHd6zGkH893sHaSnHnTmgK6gZjp6/uL
ym1hJb3zTZyu0QV0pTy+YOfq75hfmzI/qP3FdTBrTRN8fjH5rSu+AueECEyRbZozH1i+Fgd46sDn
0E+rDJGAsDONn+Qtg1AKhKVCVYa1Hr439QC/KLnWGOsYR9/LKHjqBCCsQKTXa43ZtCBzcPtpdf+0
rvYvWZLFPDk3/CTRHlGKjDYtzP2A/e8bI/Znt8xQK3mM0xsrOcYkEwtLKqwNfsmJdkoMTwLXw9OS
/LHt0f4oZCXl4pe2sCtcfWqXxFeaNBEjAO53SVR/sVk/B7URL3w5EOehcEzCr2doe83VI2SUL4S/
6kxuerci3xNL0qCDxwWcfOoOa/zW5EF0yggXbePL37Og/oEkRuu+AEYVD2wgvF0m05Ko3RyuU5Xt
4dGBZb8DR7AKS8yT8EUSpEes6Tkb1hYHZrq1A50au0jQsLUJuB6yQ6RRtXTkYU5E7+2/uEkiJ4gg
Pn+JyrOrj6gbG43Hrt7Q+bapu2zxeMfmJxJnU6QJQaEq6omN4P9ueyezSN5rvZS4LPdTz+YZ/J80
6fpKL3kUzoxdhPr56YloF+bv/hTRQAQDLZ+jmFH7AOUNZ3gI6wz+5FEnshrz+ykAkBfzNUsJsUme
IYdQAYvkMRFfhzU6s3REkWEdohNcXxV4HuwkxcPyttOFbTWAwe4eER6rC79pHglpdNfbSMcKVx8b
j95DYdrrB1XEZrfvJur7W7JMi5JFlPHRCiqpUOuCWjWg0YyZ5BZX4aDtlUs/nOwaxqT6xbSY6CIr
XyiZScpt9g1Y7V8LP8YBBQ7NWZ9IACuuJMDzSNmtDi8nCvJMAHv9IJNrl21wJ6EOGDo6cMsC2IMy
Kvblrk0zfa4iXGc5jAX2OY2wJMMPfWD8Co1kHgcsgSA6pH16If8+ZGY89IhsO4fkeN8WohUi32sv
1UFe9JQyOZMcjFmfA0flhCb40g5MVWUKH3N9HhdHmmY5kE0TwzhvVFkL8NLeHPZ4KWfwnxzd1evd
lrz+Cfgni5Ku3S7Sda+G8dSuIiAF0FXt/jVePLDAba4LLKhDYTVyVhmEM9xU5K0zPYM6uSHbYpbE
HIFiD2WlQsiqPzUEY/E4cF1+K7x4Oa8cdwIXpdUMU5IBoaqOlC6O/iSRl+prKA7Jbbz14pvXtsSC
/4UluvebVGwDkLyz/Qfaz6i3Lq5FO+dZWRBRV7leBDJLloJfElzPcCZHdWHTrcd+MVkKQpkVhQ3E
Xp9qIQWExMLbMGxJTN9l68TuscDtLVlrQpAPVyNnsNrbw0anfidS89CVAnLz7/cbi2xH1R1gGTtX
zDjyNF/rj02mWuzqsagzsCB0g+qdUfgr2XYzj+QKbNP10Oe5tSnIsqraXhrAWPQuUdKzrs690rsk
xRxmsqsxQ9YiFHE8KzzQg9HyQKIy3mKvduSoKVSraCW4WCFl8cWuOEjPtMJxZN/nihTgs8rjUJJ8
Ore7Nalw5+MHpvq+2CyEgUDGm/Sr5kxgFSvnEQVSAe0YyDh3PCr9Ed/4XFgVD6RLQamQSDSTdrUK
o6J8Y/WEAOjVx2gV1ID9FoKZyPP6xsrWqXpOxzXt6ELAHKDLG5cbBdveqWPTpAp2h9/hYCHtx7r0
IT9MStkIAnrpMr+WI86K8bcUYs+pt9QJQ8s6BqHUdFECQTc5EQ7EdHA+ya5fapjjdctZrJhDgn23
uzDdFZkAn08aPLuP6/MbPcNAmA6sg2OD8i7sXJ7aaToGmmyaeag00yZu1QX3T8wWSpxL+Yqm3MzA
T5r0pwieHEf0jjo6JTkE2s3oBBKPnf6o9K5UGz15T1yY//I+wuE14UYBHTQvvSD2popIzKKqXR64
zbgfB+QF0qzvdyJdMT2YUR/lFPP/104O7WJeYNjtm5kVvH7xYH0megKs1ljbeKwch6ko7DOf3L0d
1wi1aGHT/7YjUkM3rnIqj+axWeOck9pYQ89zDjYoFyZvIf612agzejbx9gRlmCsqhwn1Qr7jWvqp
zJSvCmSfY4EGvh8EvVsgFnqG3zY9txrYvqVgd3+Cs/xrBf5Vj/uOl/Yf/iaHXAk9Bpc3PNTvIEcv
vSHapToKLvd+AYDkYq4NqqZpUYyTsxsV46b7MKjfl0pdYnruLZ9VFCFBoGBkStwNZruHlSn559CI
QuSCmRdBiLo9ZbEfYcGMPQjWrOPYUt6/YbP3VQRRHoV0AyXT8OqHuWsicWK6t73vXY+VE0QPcac7
knrmsvZLQ30pF4BqP+2HR6HbEnXuLXKw5DJbQAkhQ4m3n//EgTPPe6Y4lDsrUXoCK6WIGP2LrBmi
4p3reNiKZq6rW4n2y61Tqdn4jw2NFXPdO98Zxz016gaxP8JLWhul+kTgGCKeajE9TxfaXtyu8i6N
DMSwu2/ROUvGa55bo1AAx4MiM9M6T7os+vq2AbsANXhIlsreU2oKvFROwRMiF8/2qPhajR3if+4f
UkNVbwWKLZdApV/yWMytK0LUkEWoAorLb5o0LEczDfjE1BT5aJOBwfHucGOZNN1D3jt31m2poY8t
85ABj1mFWAwVWRSHsP0ygdV/RPbfcyMmLbUUyKoIWb12GB0899sffBt9ymEwVr4WUk73HfKgkod3
LitAoCro7oCx8qG27k81vZjyaWbBRAbyTRcFM2uEA4yniff6DKZzw+00AA2uw7j4xLv+KRFAlKJj
R5U9BDzDUlWIUGCsyxP9heyGXwrObCCa0wujD1NYCBOCRlQBK9hxkjiMfU4fvogDLhQKcRcX9Wi4
YkQ5R2WjykZvgTHrgP13hyNRBOVcv1WaxvZo1VX0Rfye0uP4TMgZq+4rNxWRMYv2HnqepsUvqNS7
pLcL7sItz+t3/0HokRQIutlZvYp5ihbx9mPqxixokx5SW+pKgFFopLESt58GJ0/gqcfmcHQZ+acT
ItNAEU+heFkErCCLUICqijy/OWvuUgZ6G6kAvtn97r4gKn8vxr6tgAt4hITchfP0ctWNBhyp5j6K
ZfaZkfBnm2Uk8/nhzHBUsub9b/fM3LXEvYG9se2xERO0b9icqMy0HAGUHkWoqyt60HZcGSc7bXL0
YgCK/5TvHFkf4k1swd/toF0ysMkIv1CksR3CRi5fOxqnft0qr3UAHNsvnhxhO1Kj11P9r4E9PgH8
ALXBxMXu+URupeIT1kCW/9/Wdp5ajOdyFCx0ITVVh9peBTiAee0WJVddj5+1pVtAjYpAAcmobo2E
2xUKe1RLn2s7uMM/bj1SA/KSCksTGg5UwqJpyIYMbwf0AJ8mxjm2WkxlHrnjcmBHo49anCyNOniO
QwgV0ZIiYgkjLdVTsFkilY/66k5VFKSrRCMOWVIsVzTA/c2QJlqpvXeu9DSyFSq3ATM1pYz70YAe
N7ZqLOhVCJ1C4xw7QnCjfHAQ/Y5TFL89ftgGSMVhl5FS+Vhv9cCPjW07WWTD6lgH7YlHsug57dXj
Bk9y8Pxjsx1kVZJ77Lu6LEbZTiqiis2Tv01i3Ec0G8dbWXU2+GxA4QgTv4rPd6KEJy9Qvp7ajKuZ
uzanRnP2Yat2UTUnQul1p2t+dQzW4qk2nj3+CPeZFvuvDO4yzgmLeb1nsAguyqYt1WJcpb6DOSeC
AnvxXGdVMVBjQF6rXXOQ+GzHixpHUaNODdjwnXhSwYIEtLOSHmmFGbjsM43h19Ba4em/gzd0kdwP
mJDG8oy9fO4ozQ2l67wVmG8R3YH6Ycu47gfBMlP3b7NYarZ+MtloysolsA0RAi37xey4k9mwMpXV
cG8IOlicx4F+icA5bL21ivlKfwpYsXgyDS6AYv90uVX8AmctRIs9/7eDmkxIpZWXTr8vEYBNhgLj
L3j/KuWRp64gV85SvVDqSYu3SIegthRuYI+9WoLjVpxZg90EUKhrG+xhGlSPXNa+5TVxdCQjrGw4
hfn8/NcVoBjRhkJTnoq3DIGorNEp7XopYd/t2pL+rtBBZJAYpFa8BSfgY07XlATFExqu1Db2CfAb
x4YE9rJan7Tt8X1p9BCf25cqLrf+IAvYgwRloOEshzOhP6LIe3qPSmnpmu3C/72a9hS4HoxlKgP5
vzeNl9FV4bvCNP2dMcuFx/4JG1QPrY0bUY1qKSySWIu8tAjlFuMP32Y93v8t/gJQaM/jV+fTvrx9
m6qgYF704gpJIXRy4nF2otrJ3XLx5IPaBxd5MoVZHDIY/GhVhS3mQkl4LI5GFOTLAwhLmrM0UHJZ
Hyjc4MDERfMAVF1d0LEuLd61CZWUVEo0PwFWzLKEOiu/FvmdUIGwHQjGEKuUf2G6sIDVGbt1L74O
2zk4M+ZHHpeDJsohx8EYznyhNhbfv3qrtatBW01QHLFSzqZeeKxEf7X2KQmcRTuSLdb82TYWVDeM
KcRB/sOVd5hkpNYionkMQVEsroHNO/zKYXg6vtSn8RmmSJKtvMAKtlGudZnXRMN09khO10yc3/nG
E9lsZlHNxIBKp25Tzrr4G/HhtSy2BprEZyWKzxhpKgMrJYMsTD94tFHD/l0kMAZQ4W3NLonDf81C
aTXfHlDxt9NZKQ6iKIuKTAT7axnfILe1/SjOWlvCyZ0gPwT5LhGP9DrF1VSMuZHFu9A6BaOQvEzn
Ad6E3GZA77qS9Bjuff3hLQCni4UhyyHzbD2EusIC+dxwsui4k8OnsxPSTVoV+kK1fcKZ7RnPwt9X
r61FNjG1l7YnN/Pl6Y2SPPBEKD1bqvvUeI5vLs6C7PSKLKFh44aYcvebNSPL5q3fanleO4ZkSsQ4
8rjA5HDoBJGTFQRZoPGxt4SEaS7lpYHtFzIzKN8RE1RTsS52RXLJoVPWTKUtLb/aBrxMR7xSvKj+
4mzhSXyghexS/YnCqa7sWEuQF5Q/uK2AjvjReHMiV/7Y9ELppraaH+eNe0i4N7kpYNVIrTxt0Hi+
JXwwqrSlwRBt9tmsFmTehHl1uF5g/6HBamJzzi/o2mqrTGf4HlXWgrKl2cyZU11JVJBAb3omYRS2
CFRR9IK5AnYxp/PN6a0y9lkFK5DZNDBnVRtJJma2g28AgohagyzwRQ7SU1tl9ak26SWMoL5wivq5
/lAWcbTNUEre5SxxhQS5JSdeeNi8MghmG6Ek4UggPBgsE6265g5HxItDYRBaTAp66tge2zvSlQWi
HvUTrOWp7mlnuIfl9dJnIQl78MD7CqEk8DTJCTpH8pDGAUFh181zu7Nq/xDM3jECFju8NM0dYDZU
t5G8SZb6x0cH76RYI/mbqmOwti5TFG68BcbpijZheBKy/d2vs3z2shx+a4YniHBwfHMWEb4IqwW8
cHiUExmqPAs8Pa/L/MevkqROWWxpiie5lZBq9Kfr06C+KbiAFNQgXExJtoc2iIDKl/CcaMdTI3Qn
0FO6wEX8C1Gm6Ec5EF2EvVSUyMcUw/Y5WLkkoaHEONicaQPHBn5ZBX4C2e47sc0AaDc+2SD6PuNm
zajpHiWd2wwnkjGw6vs7+6s+04eUz5uOOWR80BtcoR2HeybDbjxDG/qo4VNvjdP0ddoLUKznaL1t
Gjb+GokIzm7ru+lkcjcaur/hVT2PzQR0eOG7tIg7U5h6e4og1Oz/f6GLoH8mXlCqAm6n/AT2djNL
12zWAxMmA8vsVF3Vfxmjq0mU9REuu1jl1Lsn3JgKpbT0okadjrH/G/1R7GbE3XleT7vuOW5xVb6O
+hCvMSypgGsdq96ia+yFepGDWYa+so/nj3E5UNiaNTZb3tqcp2EvoL0ZNTpuhZo+XHkuTubw1NNI
aAzl3yrkME972iWtKxdS0g71CwigEyTuZviyeY6gBSQFliUOplOkVCVAfF9aA1DYyQBwXLrwDP4D
utUcqPfQ+XWSv5OkJB/fMbUHrDGFpAze7Z+1RFHHN0PYERGvbde7L6Iauts7epGgECLbfKuSjjaY
5oJnHYLBL7/lmpKLChiHjtnLBU+uOtYfNo6hKqDTpyDVL3cSVTknCYUpNN3Vul8U8EWoQBlIyjyd
APR/7R9hNjHfRpK+lYJt327NTbqxvLibdJg3l+haxOixlGDjzY9g0liTtFV7icBDOE+7ypfLNH6Y
PJBWfBanl0KQKkMbaoQICnB1xqIfVoXyeH1cx/bM5TP83nPN+4oNbgKqCtF6Rjo0OBDyyDvNcP1c
NdYgF9I2FwTbDBOtUT7A4V4LF2kqkzoX9/pzhgaUm0t80T+AHiaXHAHCFdXVDkMQpbIErdMCznO3
UZl2haxYsu4oGilp1rGegT2CEjVGbOXWXLvx+R000w+tp3uip3RAERlQk75Km0vUCdDTZoSWga2/
kV+wB5Xiep/oJWih9Kb3Xc5cQrFPZ2AA+B4fSDAtTgglN7gpmUZTUoMkHQlnxR3+8qrN/3lxcvwp
7+AeGJcZssB8/7AAXNSLPRZjKGawPKIgGrEAiZ95UVjAawtf7jV21w4iStKIAnBW5XIvhWiv86CB
j98+4Li+TI4NXL5scCi91vbuMmNYOqG/UOcSEekrl+votny8ObSdXyvDxnmb2D6HlTeI4aZc4xc8
WLvTjQ/KKje9XAK9/5n4jkpvcWUByEaGXcg44BxKoNqqTkF+wusNkbNsW9Z+Htkd1KDFzbH4oaOI
WWWsuRpNOgWZwjTEbvhumXFtquuhjRU0159OftGIW1oVze8eP2yBRz7IkPOu4XlaZbqTOZGrCeYf
8CusC+Cp89gqltZlZZE6tm35GMaRb3ylwH3n2Hb2IAFsUl75oDD8Mw5rXib3aY6EAfbK/9Ey2zGT
qQluc3+wQAWbuXfLEJ/m6L0PWxAAm0ZRqUNe25AacHvEB/1qWgr36lrkXRtZYMAEk4bkfQRUMZzI
Rbc04pWHrPKnx2GiG5sF6XN9xWIo6vZEbshV64CfbOXMxfb+PK61fkWr1YJvadRs0ULmlMLA98no
XXE4TOAECd7ye5/nz64owljp9UG7GB+Z+HqWuMcBQBPgjmthQ1EtpCL5t1p9vgTcpoL9eHCUQX8H
bwqNasAJZB2j+VDiOJZ5dIXnE4vG/MA65peKa57J0qXKgv+FdCcOli4+8m+bq/yKlID00M+jFn76
/R2AOHZL8fCJeIJTPifCCW75s+6nZL3A1vRfYoaTvmh9iZT0xqJrUqBYooCtAG3GWiL49xai7K1/
YP5Ge0kxiXdmwOJKBuP4xz2b6vYYSMLXH+dMzpa9gv7MTaFQzPr6QmZSNXY1XdxbmVEP3XV3R1vK
WE/SdXCrFGUgMQZ+jfy8r3LCgiDh/LmWCW/f6fUKkO4I9Q5F6Uu2rDaChl3cOdwiR5bZDu/Nnxso
YbuD63GjH2SB1LFPxBtPzWxwNEIIfMOGjaEkn9CEwJfESeZMVKas/oXbVBqNDkOPcB3zgYwC2XN2
g4DmA2sWMx17NdyqVOlfNXsCRe/1+usC52jpcI4/WRdQbq2bgkvrBukNAcG5BRSortP9IXOLsFps
NbkRw+DnIBaHDOL7c19Av0o9i5Ilz/1Q6BCWi97io2jFNM7nX+I2qbqSiMncmn94ZJWG0tfQJ9zy
enIhR3+yYsl6zGLKIC346NkYOmIIOJ6wkVKORiGk7Tcow29mCPIDWyLGjqvfwv7drRYAxw2KUs4L
6LoB+SITFa8LcgaV63F7Gdgl2M7h0B08kE6bO30RSAyNH0baPl8cFe7C8kSBu0231x0ivDiz5K6v
6xwccb7PR26I7fEFEKX2/JlYFkxlLdORMKFNPXNu0P5Wic/0wzolXnb7mcKp16a8TwS1aHj6KfZK
TcOh5uJbSQz7FRfzN7ou4B8DjjQ6RGWDMbVx/BL9NpjdYaa38eTdABSHjvm2YGWmouaaxLPYARgY
R4nDyzRd23mt7yKYs5trbaXwZ80mdHSHUpwyS7nBcdpAF22CIPIKWPixybK/1dSjJXGd0DK2iTOu
gpNQNlWC4Kf7uulFUR7WtCiLianwai5HbuOILXo6X89dzz/KfrTq5QLa6+W/tk+zJfSlgqePwFwy
ilhW2Peb7RiBh7+NMBYY4GAKY5PRcz2pzPKK3NfwJLQ0YUJ7ChgLITSYkw4HINZjAelGFK/oP6pL
TVO+aG1LkLmd2tjZh/ZCyFlFf/z4+IqNGlO2/0xDv3LjQAjYyHcM3nG5pIo4fYBkSgvSiJ/2tr68
XDRq8+jJoQNnLBstLC2mQL/vaekDctCfpG1wzsrljgqa9S6LzNWnpLVNVCqT+96ag/OK+oVDZ/Bc
W1yPEIDf4QGvcXcS/DlFffEmAYTwcT5j+gS5+ydmiwE8gOwKBCo+kYAfna7gZVN5577bNnMoY3Aj
3c+JIYtfwIqF6TlezdD7rzHUO07LHSsuY4BmBlbetNUbD4pj7CVCyDQA9rr4GjCYkN3B1cJblKbt
Ny7MLfupV9aa+FhX+2ozCpWk0tIXUNCG4s/nFFGtssxlspQaIoAGC0es+WI5uWEps0P8TtT6At8R
spvjEUUCeZATZMV1NSi4BOl3jLDF0aPQn0lipEGy9moav+bWedRr0g4n+Byl+rg8bVqrc/nnhdW2
E4338/id3RF8uC7eHiGr+18lif0I/WeyCexyTueG+AIPR7mj21ybXD8dwU37WNqEfsa53wtxpFBB
txQv6g41f0THuiYi+0oePMDvLloY49vWcZg2/bmRb8Dke/L7JX48eKtjWhA1mW+Y4Bx695b8DwQt
lN1f9+NQMGdD19AWwUAidShZh/XmrbOzngCnWXXWH/VRO1+w7aEEE8yfHPwGlA+N1BrWaQwRs8Z5
QXzi7bgzvwrbm1Vauaa1PC4Kz0AMvr7saZFVWhjOA7T06iz87s8rZxMj7VF0HSV5XFUm6kCWRjpN
pPGnFOuYKm04nqedleSSQL7RBJXoVzTzCLu9xJWRAuiHO21+cdKce/4X/sNQpXXs+RDW9XkrmL17
wy37u5Zq4UrBGqFSYjs64QxusXPS3FxmhcRkNN5vDuwoHGA24n8A27yGyWrW5MZ14GG2lUVzdKdj
KJdwIZgsF/0l8I9JlOh3VDtzKxzzejDaAtsbVazEAnYHuQyBsPNiaiGfGq7/4oQF8XLCmj2Nt8N0
caP8ewLHJzCRw9gGF39EEONuuIOWGYOCqN8uqEJVbobOR+vAJ+0kIY0fFgQF5z5CpRlcjyJF/dly
gXms+1ni2T126X503oY+NvcEZBWhff+FRpl2k0mODCz7v+Ty5hT1goECXpCqqFtxBHojqVmMoatM
3erhmZiR3oUz8NrXYhHa4B33al3Eoa6i+Pb7HD0xDmukGPseVgDj0u+e15AvMPd+OeTi7O0Q3n03
IqR/ZfXSph3EquW/nxmm9eZu/vwJLP/mD6flg2V2TYx5Ck7mpjmPa1VBvDL+luaxDZD9zwuqAZK2
djP3W9RyV5rB9FmBubLvWekq5LbIFMvKKl5TIvU171hbLEo6xLCADPFFem6yeYIQPJVG9UT0oTLV
w88LuZZHEqv+13bBLGtEezX3G//CQ35bM6sNGvKMJxwmohRRRt0aqrFy6reerLOUw+zOcXXzSEsF
12AGkrbFjkojRLBT04yxZhRSD06hcQNit6I2j+ShATMML/9Shob1UyFOAGdp/7/zVXKKWuqfzrm+
rB4u8Mb8q2++GUt1Kj6bcNockrqP0o35rfVc0x7KDhqEkZvI7nZKsH6Q0HmbokfcUafQYr3blyHe
dUaqbi3nq0S6TZy7wFrYPoNoXvvRpnC4NszrlMAM3AWp+l/uk2suQwqLCg+h1VdRa/+5mYSkEgp7
MdnPIrjc0t9a+mDz7VViyEfVAOp+ya0XsFVkjrtT1Q4z8cY5s/B+meTrWZvvd5KYGFL4MhRf/qrK
C19ENAH+z9Jq0DztaHEenOcWDAx83xHxULDXA5fX7LlKwCgnZHzTyaFy9O9JlzLRbrg+zhFkOxdt
DJk/WvDjTVuW3dbb7ckC4N7kj8MHjkWliskR56VWh0Y4bzGowpSHVXIVmMkb+13gitD1kUYQtbw9
nZwaOvVeIY6ZOY7VxBOwn+WDLjnJDNVGzom+SZe+OMB3+6zT/rBESnoo8aXuq/9qqUIm8dXlxLeW
dmVNfIU4kUZ1y8zBuzQ0R70r8OcsdRBkxWDtYTTcwLzBDxc0IMa/84FGMRXrJIuQCL4M9d37OUdw
pQKancYkcW+Cp1ZqsDuAxrrbqGee+OEfG6OsGUQ97uCZ0u9fOIHZ9gWfG1p7kszD97qa/yRXgcUi
B/0MWrlrttPW18fDdIAiM1LBBPFknGj0IpJAxP6BlPE5g9RLnvQ582vcH5O4dgaRtMBWsRDp9Yxt
elupw5we0UkDhFIOza2Q2FYcx8WtA/BclTb57XbI0kgG7rfaIcGZQE0WyEL6VRo1HWGFdJn2m5bm
qLmJ+FHFgQtOqQFGsk9t9NQvoWuGS1B5DiKtAwPQR3nEi9jVeofoEmS+3ZLxZ2L/g23kPH3rIa/O
7wRdtvuzBfjkmAcQepqG9SZrK5mVaEGVRbAYzylm8lA8Wej+QEqHcb48jZC3rkgAGUk9le+npdeT
83SZgrCeH/MxaR0MViQzjaQ23DNZ6YeVExkM/Fi1vWS0CkqtF/aIoLXE7ZkCjCgxwwOOkcmi+AsN
C+6+vx1P7ex9Jz0enKOq54G6tvyvkE6htJnrNbTYOlEj3ZiwfzGz/pqpOfnBIaXkSg2o4s/DHRXN
f2qkdscNfUufOVrhoTf7nJUpPcDkn/O0e1ED+n76N8O8OjWS/3d1mTPqli0NfxEuyEqvFhUN7WPX
iCZ09LMFdoO9UnRyEiCOtSK1DXWmzG3GkvBPIFGbQTO+C/chlDuhibTR5ZlfotJIUHjt0EDU5MVS
9HNfy1xomphbxfX4jiswiRYcQMMOS/ThtbTzpNU9me1ZmgycHUhByOoT+TdPdPuXZgiGLRfkIhy+
dE8u4wst4dmibzTRT9zH3YD/woLRZtq8ic7njN2OD37g50PURW8+Iqu1YQZXCoo2EBwM0ZZVvpme
HYL5YchE8Amakt1UrGKeVAb3cFD/Prfw+xWIIz6sw3r97b/yLr+bJh6XY8PkepwrFIANw+Pqwp9C
MsFcJgNuAa4QCGGQGF8VpxLOzn5MMJjPLUOg8MJohLWYcQwDIBNwpBI6ZAv0heB8W94LfciNRLgt
BpBCghV8eZrLJuI7eDwIjNSW5ISyp6Ig4kOGImV84lRROsIvkwQawVy5yHHcMYrQYhxk+riitI9q
RqjSgdejDcC/JmV25/V8f/u3H2WQyrNdudEsGDjH4oa0536X8UeCQ385P6kRmFLohsJI/dCEjQhO
2xDHs/AG/3B/0UEuQG65CVgu9z6EE0jdTD68JxnHQlEJnq5ShxIVFI18hcwC4Gfsrgfrawv86Qe/
Si4noVVaOWn+x1gqCDdpjgPFe4FX2IrY41nQfyuMiBbBnmfl2vDzYVf6dKXXk4FrYqD99U7EssLM
1r7cAa1at5OBvV6eKjJSPGuj8qGUUoTRwqiP0A6vlThbGejKjgerSk4WdidWHiJ5dCSTxO7yNgAV
kmAL8AhZoE9qsPIcNZ/6yjh0lkmhkLPjX5/wYb2BoBFR2296OKBM0+/qLKMVlH7HVLguljCzlNBm
gPWv99Nw1hpVRZ316IRGTzq/jNU6NvrpvxcIrxinUop61TzFqxUpqXmrHjRgeu64SfMgEwm8Kf09
rqd+2N04kFTLg6nr3yowwSc8tKVH9PDjVvjhY3sY0Cv15dy0OR4aCNu0UNxtfanGTiu2HLS4FNH4
k9wgmPfsD/kOIhEPhPEVZZKmtt8nL03uZgClIbHBOKv8q7pZkgFEHwkvj56bIIqQYApaYAdaByFD
di+ex/CUi2MYUE9LHjpjxWIFttWSr5wEeoNTq15rhE/j9/yui4Jcdxa/YuSFYamhLnFjWHPrMtQy
Q9+V/2Rz72FpSglBITgMzJMJw3pKpFWrefSZQEwzwnnV6rTqirHmXBhobBUw7siQmvkHYIrFB3b+
I0fv96g4eqH3w3+krljqrOqlhR/Yd7DT+3W22AqKabmPbpovf35qASWKsmieNiomylxgIrnsIuRe
DKKokeZ4ZLPIihyGtAc5Jz56sAU/gHygkNUQBqGXbGhd0jw7iFNp/GJt78moqvxpa+4Xwwpkr+D4
EHhogRPPwqloi+hLs87k75VUiLkkF1N1S5G5YizO8eJP3IFzZ7CMg5oMocK15Dn3KuaDMzFt14yX
NBshurxvPNQ2HV/v4h53k7msNFJHzfaUVnVfkQ0c2tNQw8Drq/HyqjiR/tK0qPUhKoCT4a1GplDS
ZWs4FrKySg0694RjbQf8+hcenzPBOI60VNCWzPeEdYdmaaTJ2wohIyIUPNt8yv87g0T+BKXB49V1
CtoBG6tS5ICWpxZ4pdDJ4Kd7ad36G4/tV9+PD31p11fKCU1ZIY5SjiKMb+N2Kug/45K8SRi2/J4c
jftKWfRqJ6ZryDFKe0xiSDzz+ziLsekpBzOP4illBRJQktXAgL1IxRy73coOgUd9YksNwSO20haN
9mYeD/4L1y8kbaeqT2BddF8dFE9fDgBXj5386YhzpJg3pTYoqiXFDUfjLvwEr7ImMrvjbSPru9Rd
TpBjTdiha54e/E+cPenYSSezLZna+GgMn8gRezHM107i/7n2giRKYjqTrYKJPu28aZcBmwa5mdhn
bscXECwlgN88Cg9oSmhXRcKWB1/u5/WxBTkad6T78pVprchb/pvfb3IuDFfVBKnHFL8IKN8iVWpX
vCUMNrPtJZbA0DjiU3CZlGe6arfrfHl3KrI4xm1Qv/fP7TNkv/Vwbkv1KYLZPImxbZSBumSKpgFj
qpGotJY2z+2jjbyGfn1QPupkVGcslstB+D4F20GAvy0q1cavm5zaH9ZBvu+ZBNXqlvb+klHtiq66
3AxMKaa0pp42WLvUDIYIBgs9jWIPT3PJcpiku/rIv6TJXld1t2WRzx+t7emjSmbT1wH/zrs3jn8x
14CIOTDC/cGJRz5+kwFwBNwAUFc6bMBg9AacgngSNM0QJey/6JYaILqgzxBQqnBS14DgaipJtn/N
p9uXgdJQ+R+sCpDebhN8qvmhuaEqJ6D/pbwqDy6tSxEnEo+sObWvU1W/dwqiUOAAoJbivAeXc7av
FH4SSEyu5Oag3TaC15DMIuZ1K/igbVhhnLSl//3hMO2ouOrbGmbwZ4kXPZxL1CeUrXzkgada68Oz
gSRSR2VuDtcCcofufVrBRiemNgl7nPVPnAwwcHncezfqhtapXLO9ItCfmIbd5jW2MHf4c0ViixBS
711nZsp4NNd6byHdoQFIlBU4Br7u2jbz80Bb54KmKwQk+oU52wbb8GUduComBzw41V97XjgMJNzO
JW+NRimVP3LSD1oI0DWF2Q/6Dv+NOw/JWoUBq8u3D6y5r+Hm80v0PIs9vrya/bsmEjSi9QGCfw5b
Cu0v1VMOwrG9d4LOZYiIhaayMkeYF9Q07gBybcEYpsMIadgXOpR1AjuLx4u9ZCoR/mM5GP/cCFUe
Q07/0ONMvZxBjer90fKaR8pH8OejrnXvkbmlRT0mhHLKu4GAEH3vcLy3RyAxuJs/eko4ihLvQ9sa
Qib9SOC30qi8P6EJ/0CICEg/Lfvp+bbZQUW746IOcbCugl/WJa9etEGkPRg6mEkVMNuWMPA6cxnl
M7y/egsyhl+d0XOi9W0gsRunqtcbPgPIG1yLEc0MZufNEXhqhKo+PCgbN8Vgy1uzOCZT9i4HRwX3
QEzTitJjVCoRb44JtUCbbVF7SWDcCtIMR9wx3WRjXe3ll39jA9aiLGk+ZSgIAXqRyK9+KeYxhbvS
OIMaCaTLqxYRXl8OCVSIdXJ8qT0yZ0TKkLN1IwKI0MKzdiaF93Dy3NvAdgNqmnoxLc2aicmme+Cf
6qxVNshsEUy+UTBBwOqUUxdHH/Kd5yp287ocTWsKir9zlI020AuBiW2Gyk6xEZa5vRZy3fqjvbVa
UMQW7a8Pe2GIJyywqnLR01MEqfhiXDt2blXSBB0XMgg6q+S91v7IJrORfGxiHU5DufZbtiAF+gXS
nZtluT416X7eVq/km/WOY/w2eOUx+58UrBeS/APd6bv6cDBfNI4aeAQOYiKkODv311/qGo6RxHeq
5MRU4Wc6oyP/PSwPL83AaTUB+YAyKBo3isXCUiPmdITrtTFlaaYUB38XgaLi3gSBwakpKFWYKdC5
k8tuH6oaEAT/arOiW44Y2yNzjDDApsU+3/yG7ejYdAgXcNAlcemcf2Y25AM1MZ8/mPkOkVJy4m1w
09u1HwteIzk7n52xOdMs5U9OYqj8hpd5HJHEbKKUSRytcui8zp7QcYlHeQxVC4/Fr9g8CvakKj5I
nXi5h5I2Yep5+j73sgO6MRhAPL/xsno/RFkgPKHudeLAlr84Bk+GhzpElP1xzjO6egTrUowxxJFK
RgiHrZM5yguDjLcYGj7ONLduknn5DW57tRvy3zJbijUaBpuSlpTTIQvZ45L1bxEKviZNouNC6a0N
aTmWY29p+yvTFvW6k42d3HmItd+DbuCLrQ4Y8nnffJhxksNFU73eECn4L0jMVvBhPzCVo75At0SC
a3JaFS6XjLo0C1+MfV7OH04bdny77AvaKEyPeOJNJCq6Ml0GiIT9ZTi6FooQo7H7qUcI62cIjELG
cYT4eE3w47A65S4H/BWDYyHaScoUjaftaYf7OyaSsteedkvYFJ8/n8s+1tUOTCKh4HAHLUuzlaFk
41/+KUdhLmvXYQgtc5yjzvJKOHekorfVsVxoqnCfBVPgLsWydo1drXPzqJwnZcUOLzRXjoHVT/+O
mhIe/i4VN4QHrlp2hnOgzMNDry9IiyNeWaKPmLL32a1SNS6HlFf7bwmBXbxqF0agdiaUbhRZCbiM
YK5Hb2J2OL0JQbL/fRtaJBCfnSSg3h6rkLfFIVCKb+lyQBikAaGXR9pAw9xD+MuWGn1B1jn3tF9p
9hlrXOO15Sochm3PM7SC1UuqOXvyBPcDUxYcMjOdaSgNSXJ5ItXpHPEG3WwAT+m7G4nTFz4Z/Fyw
4AT4uD7nQE9kCXLwRbrON8lA1AeJq2Kuk2rws6m/dFDlciStJyMNVaQGFwmNYJJeY+3c9orYGNQV
BuGJdBQWB3wHGmEaakURff6UmORuGrJ7eSpKDuUE9bR1RWXRfoBrMpYEw7NEtu5cv4a4HosLNeA9
0wLvkoVFMUtbHPxmfi/qllr6LTH2fAPJN4yaY9XTA3yudHo9NGgIBwC3caa9M0icP5fOgP7JxdRL
D4lNH/u4FiYAGrtY5frKzwAbypFLLzshJ+V5AK33xhFztwipvAaOIlmvKOEkmcEGOYb634/qn6x3
fPoEjSBgTnDj9WEPIlMQAcdD+75macX4V2o7mnEF/oiX3m/RC4DUxzG5NE86tRi3LNIMWPkM8svj
BHd0dMRHGjh2kOP6Ucp1/gtNFJKVKHUSgwA+dP3T89yEbFw3PtYrha4z7oupqXHfZc+cdcYDBjAG
TgROgVx7q3rFCmvQgUvRFh4oXi4H8M9+FS5W1f1nSRqlBVpZfynoBbemDdMwCsNrBWU3M8VNNICf
Q/IXIfE7jb3l7DGNPl55sV4f6nBV3gP8p9VDrf94P3GtX83HTlJ/kwbuebK30yatVYjJ2jb4pAED
OQPh1FyyMR8AqCYsWefoPWQt8qpuL60HQ1E2JelksIsyHbxhiFQQrqQIrPRHy92wODkARPCOKxsl
1bMoTjSZlPCr/v3SUI2I1PGZzO5ax8EkG4P9Z83PgqwRvG5oV+GFDHtK8bPBbTHxj1aqjvmqiUcr
7XBFprjs2lAFhzJeWfkQCe6PPmbQKz/EXVrULQAJyCRc2/Ki1zrfSC9phTqhf2qvCMhF4XZqipKI
MRveLWVrdQ41AT5iYF1Natj81mfOSPU2N2Xq7O7OE6gtS6ZiIKPTnKeCrvXUBLGVDyZm9REcNfVB
Di3iiclWGzBA8P6Ddszt38eleiAQ53CpI81oSQTNlP+GDFA5z94nFqmiSvBDpHCcCken7wO4BriF
At/MGPocwhQdhc3JQ4Bz5COCTVeWCN2ViuwkSuZToNFxJ4XnAcuMG3Ecrv49XlVk7VV0Q8XGwWVX
uelai1Jb3HGfIMjnruX3RWEvhU5JIW9el2+XBpgpYPeZEKwVWXtBmgksMR2kr69+S/VripdZMVyX
rDB4KLi23c1deKe8GWMd7UUpQjohiLYVYVk19Bz1stjddc4UUwhRDRrXnYoszfk3QFw8q8e/vCT1
q+Gm1KQiKgp1t4YP/M9p58kjHhMyHPMUYluM7lA2CW8pCu+7+9fLQFydSUNkPN+YajbZgVxyfaXL
Z9xfsGZLlyOxZVV3sFpEJHd9uikk8GAX/WGbfZ4TS3gAYuHm9lHAAMmhVKeNh8cA6WzqsvAKD3Ai
k0xTi7OqXZwdzQ5299zqIaJ5J3iF5LP/nV4HKFRWlAO6FekoLXeAWRQN7YFb2RqRLA+qq99M7tm8
akj7/BJLGdfq/5UPkuTxRjLL0r8JXeK4yJojW82bm58stPqQnSxLXb2DAhhC8phqOHynQ9NTSGlZ
LxmuZGeL5bVq4n1OV7TvcDlbHhW6AOgbMt2SWO1cn6p1SbkjyZa1d8oyz9NOaZHJ/zhrWiIA9qD5
rYXR89inHpeAsqg0xf+Q7D7mxtQ3pSm5BMM1TbMNVsC2MUu7KTYnHTpX7/pFm3b1b+y1eizV/wxg
iS5r/P2DMvo0wgglJOQqCrVAmlZYs3IOPAE6t0NYoCBXDWSrfC8GH7e3pA92suoZSub4YHBV46yW
Fdu1tO766Y7ishGPOlcNqmEXFr+JZiuWVGVC5vAW32VCP74j97MmyDfIioqEZp1laViqAeo4BYyP
CtZ1w1GHKGWGdbgmzcm6y+Z5HLs8yVCgRg0UQ7jKeLWLsKgMlHqn1RIS4hYl36VTfALIJs8rQnXi
6f5qKOoP15biOZOFHdBGoYTyvoPMoKAUsv0jLTE4o6wRz2aJ0akFc1wwqng2SIyS7EyY0JT/s9Cg
k8dunZ/p5O6kdUCUudbqKS/sWeGgO1a9OUpgcPJRG51z3edi63TK5vI1T3P262HHJJHFYgOQmzfm
ANPYN807J2Hh5e3I7vPe+27bdVVhdBJG7yQIzzA5/vvr00wgRpq+Q3Dnavqj8Jeg2fxFqFllUpOB
cH/b7wthJOydRAWp2vzJalfoQ45jV0so5xUmm3W5X1kJ4NaFrmcCg9Tz7NV3aWoe3lYRB7dwcbOZ
KO4/OfkDsmVAQCujTtkNxF5G6hqLtC8XfH7tb0HU6n9/J9T/n1mOaBoTlKH05EZ87bETn1dA/ncB
UJShM0eMP5erPyAB8Zg0ZGzVnXNIlK2/qJI7kkW/rRz7UkYoHuOdcy0wNUIIyVpAey4AKgBVSv8t
o04ykqSFzB/gLrUgzM+r0AMt4OmQVJ0EM3w4yWtyYhHvJGy2YNuIeO+nzS2XEofUuwIqPV6B+BNI
7O+h/HODxjghMC+xtK+GlTB1pwDrqWUc0aX/+/MjaCrKYrFELUIFs1Z/vasBVwHmK0BY5Q2Bih4D
qsCSzaYAIPKyKJkmxov3fx9ZgXl8aXaSuOkXLws5qZsTQYoQrkw9F9o2Hq2SMtxaXna13yczK5df
kXNi2FTV4e6nENv1XgiYtgz7u/dwSKZpn28IuxkWNrIPJH/XRmFs231C9epa8OEiKycVIgZX7RZr
scvpaNr7XxR5DyyenZtTbgInab42WVPyf+/xs+b4mpTGnXBc3Q47j9bA4RkY67UHBEtcYDNpEK7n
JX99K66atZLtF6tzO8CUl08KsHIN11avRtsmPeAWfM5BOjE5G0VlCmDD9AL9wCI+GaiPKyJGEKCy
sL+n+F6LsQqAUh6ZB704bh3JdTkuqEi+TyGtcnI//c+j26OLmjmcsHT5WIXXUMpcuFaqoC89GtGf
YoVX8iJdGIAI4w8tN8VCKQ/gWZCMipcDk9cRy7Jn8BgoGm4vHmEC79vgeI+SMJsYIILqSx/Bcr0i
g+ZPeqk6VWlqF4Bwg5IlaMEwpZhEj2BQTWUawqIl1OJIpxi49xpdY2jjDaVAMg9lQaPl1Yx/oKPr
p/4LUGTpCyS/EgqIn9UmcMHQV/cpSCIW59WdTyTqgvKkPR2rSbvpGIhoStETzsu2domP5DFT8haM
3sZ/dTUqDUoMV61tbg6X+F8uSkvhTgkLAF4ynU21IKqEXyMorNw/8UmGumjkmonWDiv5iiV6qYQA
8VAWH1DzCNrcq/OqhAR6fy+3TumeiTUiiSbPim3IfbPVOEmXx5V3cJDdRIHtGfGjej7tnOEMwjmu
10Ka3vM1I8WZeueXCEbQtlMFGiNmNLhRLEBvK7fQPDrIyp56Jf8VODBBKvxbd3IhS4UdRUgGL/3S
YkptoAxSF1rmzI42jayRp9arv3cFQLtOCFbFfWgFewCEZ8c8IdEe7A47b5S0wdYfUAlMyJ92W3QC
Wzd/UgrGAqGuo21WHuV4Q1N0M1di8hqHqH8X58RlYlN9OoXBsSFKbkC/LjL5Nxbh0gi+SlQo3g5G
CxP77LOwgn8L2Mw/bZClnG3nUopRtoKwNL6PgHob2bDTMzwBWROOSllPTrqc8lSRZzXY7vO42l63
iQFUPHbjLTBQTTqpA/rTBv/qzcL3uID/yySOZsELcUCkNf4kgSCRzCWQ5AuoVLQ+bhK2Yeq3Iddt
YFkIrqzhGgp8IchzrO2uTtj4B8DxkTHAgKZH6hLyC83haQX8q/hbkoM+JWceVHFsBNR6b203z1rI
V7wsi+jMrzQ1oulkDIIo/i1/LR9vrteXRRfcNfuSg4YZYYIjb5pv/ABE/6LsL2L8O1duO6IAYOiu
kguXMT9EVAvyyXXp4tIQC8wdG/YyTq/QCN9Qe/1DqIXDs1mvXtzqeScOjextmwpq9rFi5ORKxDYT
9GZp8UX2fsNd8FmT9TZ5aiIcOOnHN2LW3FEySCgM/DWVK6NGloM+PdPrYq9pnOehbU7a1W8ZWNdv
PcAL9DtIEyOwnpQzlNep0Lwh3kj2cyBBpukyu7NRkDN6ake9leUqcsTWcVA1S+RmoigPP/BIiYfp
HL/ezmh6cKzi70lM7rqOc1gTZ4AAeNUwGdJ8cP4+iRuV6771d8OaZAjKNsxkHxVVGJl/whmdVty5
4lszat1fcH6Qp094rXvnNIajfHr/lHT1Tajsbl05IuWP9OJJm9I+eevYY5kfEIEhqI9MrGXCFJOC
iITZ74d8WVkTm/sJ8XSntjJMZa1CWQAsS6wPbKrHOBQsvntY63fDHtdDCC8vdye6pLMY63DP3Vt9
nzxBNzup+tYAJDev5tdBwIHWjl+Vk4wVjpVhDM0qJdwA4Sfbs5KfkI76c6d2pJvtsYWFEg2Mle+Z
U07+S374bh/BG08tyX45brNBi9BqiJg/8I8ZSRHE3Prtz3U4FOBAMhTqU6m9Hgj9I9rMpIYRlUd1
BmBSvoVUy6Z3IsvKBOFjQ2BD5QWvBhKZ2eugPNidttlskTbDucN0p6z8Fgxej9Avvb+H+sX08gqR
nJTwC38OBhTwAxdc0R6r1HHI1FNRtZarru3AlVvrV3s65jZ52saDuEqDDC6pZby6hJEEa2z1YmvR
s8LXYj+4/YO6P+IzxIJRGk1GroPQU8Lq33V4iQnQt2p7A2xUaL6Cu6fxg99YOJlWh+5YWqi++spC
W7MMFE9Jn+cCMBB31EoMtEw36roHkPuTMzFjUeu6d7IiqeiJ2JT73XsQHS2zPTJqvUnrFfJHq4Pl
rTbv5itpeaC6u5VhrZrVDQ8NFFHAPslarEVPx7yYS9tSwUnP0aTu4nvtAhn7GddV9TSltv0bDDZJ
964vsOQmQst/ETZlERrdPXT6jWCxoJ6mxnmYFez2Iy2E6HqVKR8aWOBNR9ERas5P9TQk8cadanDF
d41fXs91urfLL9dvuCCH/yETrBJErlEzGTBMo4DGqWmxIUuafv550sjoS3fPkf6E64vXylPWBAa+
d9FWPRw+MDWvywfkyDD4Q5yh7Ge3Ch9NiZRlBQOjS5SznifDGbbwjg77uCrvISeM3iGzIqFlT8L9
9x5Kalf8CmqmWZXIOHFMh7oanUpceQSIDoAC4qoZ8vbzOdDYw9PJIH5vjjDaA3NZj3u/zfU4+vg6
XJF7qnwfBglMwJAixGZGpfU1dEyD8GldSpWH2FULF/4bKO87BRLAfk1Qs/Zc0B+xOdAbbDB8eoN1
mK0DyYzFEUpPxqzv+3817DufHds0K/6P23+0jbZxAsIgL7yRLeOoX8kMI9Xhn3uv1ZGx+n+zOtpb
lrAkSzBLI24bI7ZKUvy6yBRDopijqjQ8piY1Hq5OiVE5/uHJ4qtnnMtMRIP2/IY7rGjS/pdIMS2o
vzxTglPYA1EjhvFrnw7zWcdCtCrFDGJAihToJ37qKJw08f7lRTTzgKkGADve98rvaX+B6GGpR47d
yTRJwAHg4MQLLH34ZZMN1vMxR8vfPv/+fvlAs+sNMSytbtFjq81XpuJAzFwHsaH+49g9BuVfvQh8
Rj6m4zkYhKNUPuf7SeNB6kuZ62a5VPysHodony5DH2mlGU3YfBW2DhmsQuoruzDN9gqssCixdysI
SjKCnM31hU7nYSqnv/xdA9Bw+FVe4Yd6bimJ2TSAPrpLNJ0SPCRfi9MBmyulSEcsIAcTjGHvpewV
EfItAzY5kGkVgJlFFhltrI57BmolzOBdTrJMpqsRrX71j0KNRRgT6BeiVwa6KT/UnvP7YtpSsmm4
d0ZKAUMHeC+z5BZTBGLZUHo/T2tLY2+ML4ddrDmTMurPytl0QMis8CV6mHQW9ib/0NIZF5r9/7h8
ICckrayEc+DW8lsmgOlx/jPzUmpCg5pL5Qtu2RtZIdfLnw7SHfT7342Qqn4Mm3svx5CV74tAYnAX
9KNTw/KiQZcWoFeAdY20rYlogKlo07l+0Vn6LP11pVkaHQdw849CCeZCeecGPbkxqlqZFx0PSFPO
v5lYIl5rJhIVSvEKwDN6ZQcXuDwTaLBi3pry76B+hnq2z2ziDcyk1AqEAY3aX5Xovvoqf4NyELdc
jzP/FVBnS7Bkfa/r+M8WqO6SyCPWlI7HWmUFLK92NszUtTZrKwrj9yMTPQfi9ko76z1HT5pInGrx
abgmAfS/PNkoBXzTI5kLvLR6j3KQj+T0lBn6YRh2wrnlA5H0zbUA5SesDRHC5OY7UeeIbkBHejbm
1jtqExa5MuRq+QzWoMTWViKXjWJZQ4sF2O5G5wvIgpo9xQC4I1eo+ps5RucJ1DIqsi6p5lnauqc9
eiHKHFw04EcJ6Sg9Do2d9LBixn4XPYt49kC6ZqtGXoyjeL07+gu82VcSLjqffCHUI92wodrlV3Ys
N9AAjipRQtPRmbWWj0lcCvSU7sPuBLN7GZpqEN2s0YWINxzSn2prK3SF5In2cmkx16FcRMCTh+YD
VkCd5hHsNSsGwvebu9SxT6GNDzwE1nFSYkCJ41Iea/8p6VuyKec31Ja9A1MLLybfc+ERQwOELgri
eNZEFj2jOynu9OIdFnruIzhJC91SvuphWx3ORQJ0h5A0s0hWg3vdfzkwb0sIEjjGhNK0XoRNwkmd
SPVOpXFHhbJ5RgYkQku9Y+JQQJNOKG0qgmZrpx9LIKiSBr9BqvR8dbSO00NV+ku31lp1RmiA5vg/
quYgAAesmTVsIFCpiFfnlgy9odK6Eysq5WExX0bmEb2jX+sBybaAKN4Ojwh2wlT5Cb8jhRq4ISwt
MVj0MkB1G85yJbVkJ6TjlpljEq0EOluqLcH+OLTQVzEiL8k2IkEdDwJ3Ujc4xet4eG00Pr3DF0NG
FK05BseMUhkNVA3h/Vb4nTQsNVhbXaP3qTNvSC3YL8P2S3tsS5BIOolNH8HxeChfT3UdOYaRu5Rc
smebvUb4J15eB4c0482OrK/zDO0yvL6lamZ5RQ60mvdAt/5Ol8hi0HYeEiGdnVhqr2m8XIMWYncD
Qbs7liRRDGlVEr9fFt9+JldIpPnUKwakVgVydgJcwID6OU9exN1Ncq35h3VMPU4V3qx+XhrzNzA1
8JniwQ5AiJq0ldFdPen4U4tNVbOq9agF2ORgYMeQlh9+MOchYq6VA37BqoAblTdVLaanyxsViPZM
5nKXn70VUmR8w1Jw+2Tm023rTj/LoJQ19ekvNRy5h+12yuj84TGAdyWaAewOmE+JhhJfLNmcMrkC
LwMNVj53Skb27xQrf39+4DBN8Foiq884gd9GDqOZn6+7EvW8rJBrGVxTAPXA9dBt9RxWoun+PV+F
hXFO8JHiirGyuhbF3RUTKeisIiFSuzShbiia1uM6LxvxzC8Jq1DuBevsml942smIWm4yS/p+OYZZ
vhuA6aYM0tnQQfG8+/23+xA7KPYxls2CTY5QGm78Nc9+bgMqmAoXB8gQzOlCgikaOHj77hoBaBx0
UYMGG1qWjsGV/o7MpC3ndFJVYMCBb023AeI39zz6mFUymnJ2zIN3KsoNP5WFaTwxAHaHI1XM09PG
6zhJnuWfBT1loKBUBVcf0WeMCdKUqY2UH3TJC/GcfLGL+abnH7oKDAxsO2Lcqdp3H3vBlVg7+hoD
LXGBGOhBMW/Fm4NBLCRhcCCjDv3QCwfsxinGxReSDH/n2tDFH0AmYnp9+VhlNuw+qGR8R4v9eKm/
DMTkKCXz/1u3n+dmFNd1xpQhc2OlN9MJyPq4kIIuYSw17m7NKhvS3GVfg/SuybAHm8p1SBMpZa4l
Nud31cLaOmBwt2N2HHi4g9zeGg8tjd2wAwGGJclSClHwzWdtTEEJ7zmo3LWNp6Mbjo9ecHgpTZ0Y
SsT5wTHPbhIsndRwHBR2Z8NpIEvydPqqPWcDb8LaeeMalE1OnLCMyfz1rNixBLUWKW2WeHv8VLiI
x9SFGi9hnKoGrQtdt80pjxH8FYBDZ0qfBhwnZ8+eylc7/5nn+uP09hvT6x7rWOI+iFkVzr4xpjmV
gm+YvzDAG8AW/k3NwVl24G3+y5VyU6MJRH/FqNJ20VNy7XOCb3y1Cku2L5mbaDmTsjr+kcvhO5vB
zQcQTMFVdjrf+PzT0HbFY20K8L4fLJ67ll+RbL4adCFm/tKKyFEVXm3akv7gTVxTXjODpi6NUyoS
RMKYUc6GmZGOuluYNegmjwNJlbCGX1N+GQa4P/r8RZ5ULmqs3VQfvqmc22CYLqrJWgMmfsN8QvJJ
3Tct1pbYBuaqVizqWsvihvQJjUrGL3Os7NZXGjdgQRmlj6y+FdNgtEkylgFuskeX4KJqxbn2K3Zs
FEHbq94/tQNHTfBH4Pxn8uGnMvW40KZ01bk3gqekVA+rahHpRy6eIJxzuwfesQa6y41DbEJzyWft
5VGE3xw0Vu77L+4FkDm4Mise2RMSIJK0+0p5PvAlIQWMoK2FULcY0feAJesQW/YZpE8mGqhUFkIR
cK9fBgjQUcwVUq55o5vLV1fvyd6YQgOWUtoNJmEcqYtD6mqiK9R9IIe6pUbpJidm++rnvbpXcZvx
NIW59juqaSyeQ/xnckOdbhUKcZdPxxDwt/g1wF4J5ExXtGP35jwSaWNtG5NV4xvJTCbFX5EMQ9gA
E0nMrnok5IEZfy4tsBA5294GVVxQ5nsX/omNKU51bXW5NBWJZEqNtC4iJhQK4pz9JnH+8apuA2nr
UmDUWD0wDMOUSmuN7RrhZTjgtcdcKZr1L7/mqYfSZujUng5CQUIOSAzVMTZGdNVWLJdN1TzdNxS3
Jbg0/l+reNy5/jI3VFZk4ly/E0Oiu9+aEZgCCSn6aeRY3pRmV2tk+4gnId6Qymn/umRJ5B8NkvTE
bi/dMQbSW517kCcIQrm/rdnZaDIHDL1EnW3Tf+3Nnol6ndRZb65wI0QJu3KAzgs75n9NinncSjmm
edP2kE/eTyPCASdY/4xF2Ga0vvPWZ0RK2WP3GjIMyE7NtpWt3x/1Pz+8NM8MD+blcnu9jWVGpYS+
xFZXt54SxtVbiHdr6QcXJ2PQvx5yHUh2RV0GmvE58kaAn3zNThr6SxeQwPi3VMBX7SRDuZGr0xJD
0yVeUQF6BEThnMKwLVQfkvUhH8yb6OpbGi7nCfBsZLf42uBp+jn0/qrAbtB3PcsaedOe88ksCqgL
lpc73k5BSOsd60yZ44Z6r1sFN73PAYNAcuOUggesvRDkxh8iwHo/d+rCFQg3gaVmIqGViNB7/Vsh
6q6GwJZ+RW7nItoKMLmycvX/AHgZwJU5kCZaPdkTKBhFO7BxWKCfLeKya+KkYQi7ig6KZ1t7mNOj
2bKGYgd9TEfNSof3Zu6lYTvRu4uf7Pbpr7ijD3ziQJDtZsQEiV0CC+s6wEYy+QvqE9mnLyrnfIx1
XeRy36CtRST89J9jBo0R8qfuJF4soXMWQzCVdj5c/i6zkjTgq8tQhu90OnCOmjBGHW5EOdgLFb/k
4uFKlVXMODLIjRgxAvTJs2pY2nOmmzE1hIn31EYKnfmeNbvGQ9ybQ2GKnq3/iB5bXYlS7mKLHh8Z
Rim40nS23x9SXD8U5aKFdv308v/AoYdmtbVVrD3WxGKHCmI1Niec8ZApnWo9k8F3dQlWDhPKSAjC
pNsKErlV1NMGzdlY+iwH50tGY+DOsl8SmDWT/G7uQeuUAtasQ09FvoPb6NBueeXGNiGy4HQhfUwx
pFxppa6sBvXA1/t0q0FTgudX4agFx2UzZpoVBAFcQFK6BwyXg3nUEpUJ6+0DQb2KvwmksDYF0iQD
AOhs8Nuqdk3Ixa3/GEHI/LBIGKNLfFoW8CRfU5DuM7fdRjduFoxUoOQLJgxV/QBwrBjx0dVV8W32
jjppOQMqQZv7lIoaQXgAc8SdzwNHidUXCBHnEfECTbG0ktLfRNXCZA01EHAD5F4SrhaJLTJqo0RW
8RRvxXyc26noZWegqvM2+8wjwnnX/jpoaNV7tN24g71EViR1SlJlLxPo1B0yJJuCa8q16yYrmAYg
Qkm7hvQuKsVSOu0LpY1NmUcZnEubrHcGcfpDSBKNhBVLNrG6IYtxGd6Xe3Bf9RGs1N2rqJx23BYZ
WR1ABgnjGljr7LghrG6hGaMVomW9+qHsYSkux+hPb4na+9VREA8a8Ay8yZitrULXxRAzvuG781hi
FW6ih1vlfJqIBxhp0vNsFDCbeZwxlPoJruddB4kuN5o5UT0drpmEFBORXVJEqLnwreixUEkxIfjF
Tta13jOYVNv4H66NuaMOx103QfODRzmVqXfFj0QcoZkpBTtjmSM2/mgcFC5iQcLgPoPfjrzHx83j
JlC61qZ81ahnjHcNHwPY9LYHJRQIY3iV395aSzUEo7WDBzCKt9HjMtXD0E+9ZlK9x7f42ofyTjil
m8hBEgOW5I2dpIxOBFieMrHwyMqzKfSyUpL9lMOk/u9rYeirNENdKbDdo6OnwWuoZdo9lnFrd+hk
gePSrX2NwipQ9ZGwAmmrX+fI5vowjtOc9frCTPUdphc9YcNJXThMb6GvOhCIeovGDbUaZJgGBh3K
TnozDpFjKM6vxfUmXWes5H46dmWZbxyp9LdMVpVE2vP3bDg+bI98G53vTifbvlzzkCWXWLuVO7tg
uPTqVPoiBu4Thyo4PC9mLYqNT5KrJgp8B4ZTwAZw7PSADtwQVdfQgXfqn9SOLRjo18IQh6nByJEm
Q/GAQzag4XaORCaWUSGf7MtD+d+cu5CVNVx8Up5AAd1hcazyIm498soZFfexS9Hm0LeV6ga8Ptxj
Z8KgN2ZjEr8DpKnvs19N3b7SCrHBLS606X0eMx8Ul3UhnjHmDw0yPF37JGcsGbg0JhccUztXuznd
z8X5Q1FYNxyMzSUzF4NniArkCcxT2g3ZlhJh1bQ9JTkUKZMS3GCn2ubOWOyc589uNu2opAPJ1Vzf
bULjqEVkD5pSKRaj7gWifGDmiZnqc78g5BiL4P4OIXo57+wCcUK9W9noElqYxAci+g6S4xSVQ7Iy
nPx7NlkomXKNaFYCMQsli/JGh8W3r67fZqroufQ+E4sIjqj3YbRnp31My8Xmxett6jf6qc2Z8E2Z
MsKiMgNC1Sw6LaSKoS81s2NDSavnXO4EPnPxIv+/W/+VLAjkJSNZNspk8aqDNIheT/oE9sFHmwIq
J59gFPjr8Ny4Sej32xYq1V59HYcN34XvBODA55jgF/z/Cr02p92+ZKsllXYqGbligTVQbESoUn/B
aUpbKf89jRbYyQJ7CzR33qo4mup67ByceBK8MgcXZEK9ycyCzPsu2O+TLHKFJCtQNIwpNOTHmJPw
op1t55HIPYuydFHpjtwdsg1g6cl3+6qI4m/BtlkNuIE8Xkei8jkwqbkGiN9sk7dVICSQuNYwLhjU
KPKpa1uTz9ANOoB8EOdsYFrD8ZXJqtYTVDMpGWdjthN+73v5UAZftHkwgnHJcyqUZU+jRo6LIfo4
z55hPu+Lhdbwoh7jCDdJ2Vs/m8kcNawdSqRymwaw1V2No9Sb2FRNZ9Ah34wqcrYqkdS0iaWdz/Ur
tQSucsIitKL56zPZWjvqIMdfKJVrWgIhxJC7z4hM8MTfZCpywD9IVXLPhb3f8O7K2aU00OSpVIy6
xBSSmlzOgqccJcTT/QYBZ0VFS4gj4J1x0JyjISzcfLeUApQmf6NO06Nv+JliwG2NUie6P3ArvcoE
dbvT+tG5TQIeS8I3d5zC/9dd4fE8YntUG4iVUtsN75LN7U0/U8GK2tX726SopsMyulysR163zTEA
WuqNymCbeoqsXfL39Y0eGD5TJ9U+boJOT/sJjhO9knGsWJbg5smURS6dcqkDMK0pNsW9Mn+3ojDI
/zCd5vM/W2y3uanJSbGE3kwV7mZFbdcu2Gh3nCV7qWvpwhab63gC69TiIzkTnxMiJOcnBQ57hCiw
ZHl4X0M92RNfanY1/wO/sfv1pi9pGyZU9QLKeM3IJ0L3ImBZeV7tZ+CvtRAVIcWDjh4MEj5NcG+b
rSYLpgM/6tJA6XE4AU6CWQ4TOcQnIY4fkM0T0uqjOPHg/cq1Ud6Tz3HrmnZlwFW+PEqBwskLBUow
qV7p/Pguf1RDeQ7YlEV0rtGHWHiPYoRXDcKdtj4eptJm2u4iymR3eNbjlJpEOKavC6QCWp8BLdFQ
U1BpHOoiL+ZE1d0W3+XwvCLfniRk+VkzPumbiuR6lEFHteWbJCKc2exEory4uqDJbjoIaOd4L4IX
4WeumtbTfebpu1yeU8hOuG5A/ZoPL/sRTblJ+tfehB6LcSC4UPWVrveywklU6JLUxfgvkmK4kBkV
Vgj8VcRccVaEWjPnX4IDjxHlAc2tg6+e/F8torNxcJJ1gPoQGQXDxqFpLEm/NAd6tNJ0eVoSL21A
R7B5BDrHNlrpxzhRazA2sk3ScoTTGmkezSRRbDBZ3f+wBI/J3qI0uQJdG2R87Jlc9uosaBQ90vwM
WzDAaugOZ6uWIlCMib8S5SUyop4cfDtxL3m0Agx8fEr34uuDyFNADxvd87uJ+WvtdsOaiJdcvA/e
3TzCkHPRE+3jzP7VwYClH5tQApGIqu9fw0QU1i/XX4tY3xmzk4UHQBaM4K7wefM6YqKQP5AyhWXm
qPgf0DKxshYuhpNKq6TVlhf8D4P2ZGDdHWkHeexH2W8T2zfi2gr7y5K52cHuWUfwOkCB/tqZjT9Q
3nBF+Jb4PxggcJEpL+UISy9iAzy3wX0hr60amRmKwkGGONFm0yQdMPPhSC23UwIXDWZErvX+ar8+
fLAwj3jJ5YdW9Pctg1g79UssoN5otX87vOngN0E0mZGuZlLwFRpeIPppRilN7WPrH69sOH7hQJp6
uEIduInXzaB1PCcHHiZkEJC5aWhbh8MYiWbCzuODCCUQ1LYnAd5n+Z0pk9qeqc8OjcKGf24HW+vB
pjPM+oi5OVzVpUE8e4uBjpM00ILf4wm48yPDEcx2GCX6oAQwtpK1mSMX7ywakdCqyEU4AFGcoZc5
Ti2whJwSG5gnBD17riy8nVgRXpWf5uAy8RobWrvTyIwmoFT9qJ4xH/Ye5sZxrBy4fRaNx9nDt8wf
NOf/nBHq7od1RSx9qgy8zOnTnlhAbntRU8qcc6oVBUX5IJxb0CzNgiSdZVuKc+j9tgg4Q8BtWVJ6
tct6/+KInv5EmxQT7cMvW3MvzMWP7+Agj8O7U5KdqjUv7XnmZLPPADsjb+UqQ8XvVF9Jfsqt2V04
bTDDrTxDFMFMikzp7YJkEyq+UUVY1JN5ZOlwp3p656tXrX/kaBdmvmuMaTzhRxwqaIG/PSKmMa5B
q2L53R/j1epBQsVo1P5w0O9XSAri5w1gX1yDPWsaSagf6buMx6tPcTeoFc4nG6v8BL9RIvcnx7Wq
uHwz6IqKMi9cK1y6tTO6FbzUPB2ww3iBPD70TZGOsrxNZAkaFwahEip3kDR3jL4dfjZf8TA21xkj
teDeeFAYx11eGX5xFn26jzESuwcatnc54TFZegVMxuAoux0hvu8JyEKjpZukMf5nZN9e/XJ4nDsa
6zrz1FpB9YND5HP85JJNeW5uzXKJIVKZMI6ClsZXvwhLyOrnm/swp8x45PmhBMKQIlBbpYEXtTZm
eSMeWoknhdOq/wQ9gXWzxDhrpGxIFYC6Cz2Oj5k8io7u7IeAxW1y+DrPPHE2AY2P3vMHB58Q6s+5
i/ty1J6Dw32q0H3ByapZC3T7z+pCgt4JbozGL/Hp9qLWZAonqjE9OX28xvw/bVvF1hcRFSVD7evn
shKQQVd6gn/hsHP5k53POQve6D7T8dLGxJrHoRZpAlDNXpxhNw4P27mh6PWay6Gxu2gRe7/0UNOc
ayF+AQFWgYfuqq3ypKO2qP9jIvoi61pbVzlBvHs46dIAc8Fb2ZKVZCfRjHzv0ChExi+7I4vTIm9e
Y4XlEQUw+S/9xd8MgFaWpn/uZ4KzUryyyFA2RDbLN7Efxrk7NsV9t/8oytOJA2xhoS8bq54VzZce
ecYlHrGfJIx2OmOgBQqXJxCCU0Z0VPTp+LTU28b38WJSeY+gwS+uNG4Mqn476I1sICDZb0qK1e3M
8wyuHirW8+BXmsNIgc4lnOXhN3Blya0h4g1CjE/XV/a8/1w44Wpjst4RAcwLw5GTdOXWLd/FodAf
N1c1cNJCQhr9oKkHCBwSD8rfc+wyTQJeUfygONBrwjtO5VTKzlrqRVD8SPF7iEnztQ0e2c1Q/YH6
v7pPqU665DH/w1ZnAbHOGQeL3dyR4bF5fItSCwwi3yeAn9Y30IyE4WBJQ7bUT2vDl2G6Yz742jWo
x73CKBsRZY1GbuqwxmExxW65q42kmN3FP7BJtlCQLHIZUtfyaUbpDRFrp3QIh2nxOAuwIJu+FxcQ
Ca7hteHqkHP5bNP0rl+oOpM88yIpUo9631mpCRK9xHElxQGFqgkcu6wtPz7zMS2XfNPgahGOQqaF
wOWFL3rzj3VfERCDWM+Q04xiweDbaRAnIfUVDXDrY/MSubcW0KKkUn5qo87DOkizY4H/hRiZ5pKc
04G39x2ovAqKTnUzQ/q8+1SyspWxm1oGpHAU9xpUCxfQBqPbPm8gwfKc6j3+/T2PIRp2YHIwk0Ga
pzEltmlFtCm+gQACFdyYNPaYm5uvMmPvfFC2iSpcKlmp/bgdDb46BfbVGpgQJomW2gHjcPMXMqon
hlif+zer/LxjEcWP17wP2ndxXH5zcUvpQ5jnq8L36PIe09KL0ueS2+01Ex6cXI0sEqnO5x6zlliq
lqYT3cO06mmQXdxpWwhjGTpRNgCbyh+qyTra5dIQLc2mLHvMOtWKZkvaiMiHgGdrSgWhi6aFYF8j
EVHZNxnQq59u6E7MAkRl+3yWtBlYg7UhazN8Fp246BnImOS1vriatS4WI16QBla8A45NNzeveZJo
kmVoy/vDd3anGZpn+7J9/T+0JKqcv3ixv4kwwcxUm2vnO6a4i50+HWEkSBULuwWyN8AXVTGaq8dQ
4Rw2Hn0Qrf+6mdYfXvMNuSX5yoLqGAx/GQ19tOfVU3W/kZgkOXdAcrTkUKSNt6fXZO/30AQE2mYZ
mtabjf5mxdAW3SriE/kRqjwXEy1MP5+TUWHng6QdXGyVPZ3DQLtncv7Hv6mxeotBMfE3ex7wsqQg
N50URmXik0Adud4WbpRuxy31PI5MTsaERzQ9se1UkbZ5B39HglDZbWMVyIft3+0//hvfu0RBd5yJ
SIUYOuVGAUJlLe6IqjQh4Th56UKMlhWKQX7QxZgQ2RpAw/fGM570a+eRqsGRPWHq8x3hIp6WcSjB
c9KzdNoGNjn7sZB8dTFjkzN1Kw++vySpOL5+/sLxX6D2q4KMAPGkivgNnqOV1cQSSG81hQBGYYOK
FMHsPIew08O9pIe1ioo1AV25NP4U+LXhJf0jgrn9iVONzRJeaP0m9MXBiqC1XjXdgu8GDAAtE+nI
p+JeSqiDXn0SjIawxyRrzyyedD6waMsNoI831+4oP3ySUnTV8992eO+stxAVdKtFOMeiWPP/zrsn
qMHbkw87fihXUsTAyoqyCw3p6UYvzwHs8syvnQG1E+DzGa3Fl3KNxRIKe/G9T+RJwievplP78848
R7ecmXIe5lEO4ssIIHJ1lUCdxf410RzCBteIquNhNAXywU4RXMLcHN1YJYf5NcfMZhperQk9dzxD
1KKXMzodULuknyhVsP6fI8Q+0709aTVoXdAeQL6JwG01QI8bxJ1S11ZIPTgQbY2qg9pNKSVmHEpB
zp5d/mMEwcU5BdkfdHusmRYQWdEP4O/ktyGiYNfvQCLeMFj/bIkjsHFp2yTuRjuRCOBIrmSfhbTh
1EjJ/qBjpsGNfeSe+Lt7BO2zhF8R44IhDb+OiVXCt+7QSX84hKBOWfQ8/I62PBe3q0v4G3Q6mmJ9
Hr21Wr+yx5X78pdUXsKEUkGRUbPBvVSrOGw3HX6Sy2sy1j8318qzK0sJCmx7Qk3XVYGhCc6YGJSw
LP2oZQJ7cu6lYyuayBR5RK6m0SzEvn+TLJb3azHOAw13LswX6wOZZNTjJxYfLxEL8GOtGPXuirDm
FtwBu2Vi9E7IFwj4QTSJOuJP+JcG7UuZFyW0GMC0ivFUcF50qGgBbEC9XAs5wkYMkhaizanH+k7F
znzjKZliJJ6SUCDwV1+vrkXJOtl3UK6sQECcpzJYM/Z/O1Jyp6APeTrBem38lp031ZsGhMAEIkqn
IDP5yz/Dp3REQiyLV6wbRHRsh1ngqr1kEUGF/gLI3yTEml4ehaRWbXwWR1X1zeDSzEEveyK2u883
r2kATOPlE5cVEdYsNt6nyLWPTMAvsPZy3hk1a00U/z5e0jiDw2qje2l7EN0JasKoTkYlTz5sEh9r
nXWuXr5uCQ6RBS3iic8U8S8CyVJvoEMpiJv/zasfvy0vp6NsOC2BspYuHRs42VfL3zPfJfUN3xjI
5uh8KmIp4VhSIDrKW5ooihSXMGcIjiM8LUY8fXtx73rO/kVWekbL3E9SAcO2UYlP+s/gA3UGTXpt
t/e9uGeEfC+rzyjE0yd6acR+ak9tb6QjAnyckICJPVlqd1Ho3gDU2tY6dQigyHgE5kuKc/+ySBP7
4wk+rzV0p4a22AISf30idNlLJZuaQQJWSu6mRzHxChdZ36e1bmPEL8sd7QS9hwEk8FNL8u1KVTXh
WTensQ83ZsQMoqFmPvRKwiarjI3pVErGG3w93OX0FiuEC7GSenjfKz7dBRJ5IHI1m2EXu87LVmqU
nSPm1O+01ScphSPJZG1TxDGTdlUoy1P6yqIn/+XOk4WhICkF+DNebIHS/JU5+V089n38q7472pRO
oQxhRppD77cxpYYXQGSPhtAyjIGOPouEhhzrMUArUHwXLmHjsCYomQg0j+LGdlRRbbjb3IsEh3/u
fbSkCKYAZKul3LZ7KvtpXVTU3L1g+eU0fyvdUr3zlt5tohmpKu7A+hfsmzZwsKxVsnCbbvkzXUif
bjii9Rb1KtSXvgqG68oP3bS4BRwfmtsGpOr0V6q0ScuDcJU0k0Jb0VhStm2EuTWZl3kPBg3RiOz4
dEDbXaJeGF9P/vYXeMCcEFo9dShqSoUtq0eutZ9UcIzbNbjceLnMD8hhqk9NTgRWF9cOej/bWMGX
wxCF2yV9u+DK910Fi8feYv03r2yaj+GeCABm7cCS6JzJV+JSTEQHGnCMQgb89EW12+z5lFffOcGN
eIDPNF8YzPRWk7k7oeDWuvNGxKzz9vP85npU9DYaQCA3AiyY5IIRIZwpwqgevA5UgHGrJ1atG9/P
BbjxWJI+Pkqoj22Jok0q3fELNMxa+S3Wby/nzTxsBhdLGLhFiYPngta/QHUxhwjRzePtwNhg3f0Y
cZQYcj9iABR8l+BETfKuDMHW/6KhEYQIaFKhEUFEEwN6lmf/VT+Gd7FU6+xA+3cIrAdSbWBqCIhW
PiGb8q1/j9XyS8J83uI3PiplZOGAJf2EEK5lhWB5bqKZJVsQ74lEv/8za402cXiSUO6fWuYJx3kq
iLE1pmnY19jTed/2cty80feKx19S4Hd4uVYvk7DuLrLiT6IpcCtc37f62EvSUlER4494GGJ7BLCW
Ky8vgj9TrYbMyFoRbtlqG4funhTc1y6G8bolVEiZNQGkQUUGhrkR+Xxj4alb9+0V/+EbcDZNLcuf
MGrPQoa1v5MR53ldRSMfPvVZCTmwKr5Uj+gumMcsP0tLxNhk1qv6bfDoU/YfwQlILEn7Q12ud3ZQ
9G+aYACaYschdCyQ3ZX5roV0ombYbuKCWpPHwVr+U0QPrJHfJhBz3ETmFW6yvozUuP3Uu6TVgD/t
TqIHhyVBPfJnm9GmlJM4O7YIJMInQS/fiEQ69H5lYT7ZIKBeVpOpaaEGiAIeUqJ+ErWlh7CAiVbF
6yjg+w9FOYCP8rr2/AfAihk6/cXMm2+t4znaEyFJw389hXKXcZWPYhvNVy4NJvGOqHBjoqFsS1i0
GX3oKKt1veEvtKTc7kiTxbvXP3cEALaKpXD7O/JWS+OGN8twIE1psiw/H+/ATiFo+9qUVd/KO5uX
8B1hMfZ6TUw5HVvZ7R/paKlV/R4l2Ef4sSO8ot2HlkLq5gepx0n8+CKJJzjN9DZOJjK7eC9HWP10
e9HntOmpS4YkCotWcBjY2VnCLRwuEHuwII5KRTvxKQbEJKeTXxzcJB5l8MVwJk6eVfwEb3G48WVQ
pDDxgu4iAwBJqgBt5wpgAgmhL4C1AbN5+XUVTVCohc0y9trpPQrkvZpJI5/dkAHO+C+R1A+3CodD
8cCuQLSkhPkQxjn4SfpV1DnrLEFqxauA6sew38NwDjY5CzCHgcfTPCD9jEuaz2jAty/zIm9nFM5+
7pYuo2ZcylFiq22exGYNH87yqOD4QHqcmUQFiyHK9GRChKXifLt5PPfAqkJHDdXxRs7Fk1e17bu1
4XSeZmUbS84iOo8V9CwNYnA0mNpSyqV4jFENji7/FItL1DW2LYMzsLUlVA93/cgDO7CHkE0lytxF
IfNK/wPnL4y1D825VaI8e25i/3HKpYA/JiKW/CWaSHb4Po3lvbQpmOTWLAeqY7gFlPC6aLON6Ab7
unpG6uBmnOIZQ3kCV2XQWNHiYSPekTtJAwXRimfQh9FPnoAIUro3cPGJCghbWX3ex+Q079PyTDqK
n2UH7000Jbh72B+x6WpBZSms8ijV/ElKQUUMx+LzozxX1ZpqGRzo2P3NONtcXJiiA61GweHcJv0d
76l0xknr+lBix48t9dQM/XFg/sGG4fQ9RxFJmX9YgepDdiXPshGPWWA5o3Ev75vEVL4feopeQqUG
s+dqqAQWkNmI/cHFugZ2RbJ+IrlzU+UjJkKQ9s9gYr5W+jBV9Phdtl7Q3LPtKEerlt2fu6jARyaf
xcGCMVfAiQ4MzaugiIaZlWlX5RAE1e69yHyg98lNUe2qDRkRsrt9vcff1hWKTIxTwTQi0dK+cWkp
wpm1TAVguU1bHZa6j0lnFep0i4fDwPjgh1oiVAUDJEA47/dZMdEprXgxJkBTjoa0CTI7YMN2kDgd
zuJ7Rh8ufNAwDjiNKsVtIYiPF59VUB0FVCiFmFa4QK89rZEYqEb88Lgq3FcO/WONtNnu6XFafyjR
E61ql6g00aCsq03A6jibr8o2Z3qoOBy7udYejyu22mk9MXrV7Mw2pgZwJI3fOXJYUrbcby5u0XeF
2F29aHmEIKFYcsYKqL6nU/UDqiS4yHsurJUuqpWiQcIUhmoB2RiRZPy1C63vkZTAjmZ0gFSttAEQ
8uGuBtyEDb2ZGSY+8AqP45wVcc1lL5/Zp29jPeadq8kVw4B97ZbFcdtath3iva800EcDUyjLxCfW
tET8fx42vANeaIQOGFpOHDGL7ON2xaPlDxucjQqWPJvqsrQnwjrUx24dy7mPt395cc4Rl1Gi1yI9
4ZD6DL1Ke30RGb/gR1n1Xnf76oUP7CsSECedCWU/GYNZj3VNVT3RDJXwXlj6gdUrq70DjLRVJ2ZE
2QUKA96TEd3aeEWqO/WSj59VQ/83v2wUrCd+yM1ZpkPXmDLdvrm5Ah149meIStGLDkMVqygSxbFa
S+7bZ1UiXM3CfTICPBCTCp1Q/2hOqqvZiDvz3s+hxrNR/jxkiws/Kr+P4/SBeWxkA2YlvdAs9F7M
4xvaWUG5PMBKT1pff2YOB/QxcjSszIee3HrvEjt6RS99lluZuLPRKXZkoAZwJLzurJm+OxgSZDEm
4v8R9+C8y8GivFniWbSW1WuoY0BIPEYIiDxxerI/0LG3L0ot6TyJOkgdjyI7Sa0MVzg9Wa4u4QQF
mRkZ/Bzsrnfz9Zvdomgzvz7QDTndb4zRHIIjFN5W5NgwmGa4LfZ331wmNcIdPJY25CiC4L3x8O4v
RvBEbX3mBIkzt8D62jhTJSUkDfC3YBkUPWqMabgkBghzW2IoojhxqpSfB4Xxu5K2nTPJYnguj5PG
6WlAU1DHTa5lbgsXGEi0Z9h+0XwdmBdJo8+oM1sRa7Ix6hTnBpSxbW3iGvrp1l2DAmcObxHbvdyM
jlBqzUeLyGNrtC5U7FdTAhgLMecFjjXvr5qk3jVhFC9ELa7M+X83GlaAgjBXwQKkhuDenGCexb/E
ME0S2fNl7VEkwI/K9lPiaFIGRDCcUrkN3TZbo431UwlTULvdkW7OdEwpAuDULPOM30Ty2/cKFqkr
OVxQpCbwcKAuPWJn41y9Amv/s+Z2IxJHGN4k8b87u0ceZNzJLEMKZ/wcpRZ+CY94WEap9TNy5Rnz
GVJRU/DvSrs14zNVKl+g1A9LyLkKqq+VYL/889jCmfeHRHPdn/2A9FfuWXs++UANQbpQWTvGKDhg
LQb6tl4dyGzyM7BsfJhvqj4rvNRGhvYr3EMvsyRcvLlWXiyYDyqk7ywd+P9PzlkVVeBZgorKQYJ0
nhZY3j+mV1n3zp1fOgqfMPN4XyPpr5T3nF3rD28cuXGfKyDIPpU/2T6Ox+TB47/xVa35iMudzeVZ
Zi2eRWk7pvCYM1V5VGjKm8i0Gz8Wch1S8IwOcsDrZ4FyCbMArDn1XIFfeKPjfOeju6+5Fv8ApQ4p
m43GAomyHxB5S3QmndRhNZBcQ7CxPRdOotociPztl+whEH658RtNfEsSamBDsgKamuDA3GD3bnm1
tlAkzA71tdZnc6shmQlPOcMkWKqP2p+LSHZXllDJ+gsQ29UcC5WPonB0IYIwdd0XHzBLEuRxhNJZ
GcfvDh5/rRF+EjN0unfOFWbhy/SOllFFsY4JYuxILC3m6oJHAK8O1o27/nmnu18pTe4FTyEvrhko
Kb57l5XlnyPXbtWoZGZnfqod+Gy1DW30OqI/C1EetTBsRXxu/ZlF+sIeBT7iVa063A/ensnWHI30
glPvusKwM/uaaxDVb6ZhBxfcJedB/e/QDl0ShHVGb79Jvve9JRob4WUyNMcNgeQa/PceE7M9URmh
hSDG+aycyZ4eFxRjfDxeS15TKlq8iRAQW9vbyYb7UdwmGv6VsDA+0r8YYQ9ROV1z7/Gw8g9NEWza
gOLbJc8lWktVpNsYvnSAteCEYxmDLxjBHgRZPELTDc+wY0V+xesO+zVbaX7TMMYw4kr7t/nNBqqR
dZm263IaQiWQx9i7VeM0ec4mA0t+bCqoRcBo2VUC0oW4C4u0YWlPOVOfwYHegAvlYa5HKi0MulIx
Y8M6/xNhLkaXcWKodtUgRod0cWPbrXcn2glWLdQWuvEzz9aRo3PYcbF7WTGcMLCL9VOsTIZPIG7/
TNklAbE6Wym5pAAvnmGeDA1+L+PSyA4/gWWI1JGbOdk89Nwh8RYuRfcppWBCEPUVPfkqh2N/ZbTp
UqiP6OdjpMzoW2ssfbg9valqgWEyvUvVf0Z4DBOJYZHZ3WJ5KwQcZ/YuxHn5q1fuqFqdel2SGX+S
pcQkM9nEEs7XUqWTqCcjgKQAmHvhLwbezoCcVM/puEsbediht4EHYYfNfpp+0idzz7wYAy9y0xNB
e+yuW8K6jf0yBhUNsRwZR/FiJUqXdvMgN/EgeOP/fuF2yfsh4W1jB/RVp2FNwqO+hTXzCKRqAM05
jM1msflzHcsQuW0m1DNQd0aoJ4H/82Do9DiwNDAuEvGYDE+5bEb6Gxs1T/p0m+Cwc81HuyckC9fR
QoCMGpjllixADiRVvsUBctDogPrYnh8x+Lp/cnd9+P+YAIhZpN71hh7+CctyAF0cIY0y5h//gcSM
rrFbgLgi9A9iF6KgVZrNaBtAaSOlerOW3pUpRIXyrXK0bgfaVGmiVrvw5lVE2kuiEccHYnTp6EJM
65gvxnwWaQnvCqBAqBfgetbSrSrxLSLnwBq0urrKnKpTXWCEz1sNW84L8RdBPuDtD/tuXgTdhybi
Sf68Tbj2Uqptcn+MbSV/0SJgF3nS17U4r2Z5/+BiJ14v9vpqUYq80nU5kha1zJd3qAnMM/D+UMfX
DNdAsBgGEI+rcmz/iBTBUZo/OHTPuTjaOay61e8vjA6q/JAQOwoS8zCE1GGKM8S7yXUgLcfkhXYs
6pbSvhODjTMWSgOL0baWgRyWiouN6W1F1GaCbgZijO5HQA59n+iYck3E8KoBSXNqYfnIDIDW6git
q87dTsY5YzDEYWUeJKL1fEbvEZyGrEx99tcGewjxchFi1CicMPffW/+5wkwoy3R0kPsaZX2tZonl
3tp/wfpp3TQY7sDrNwCIoxCAPNLVTVXi8xY3ckJPTH2WYkvbLm8lCxk296xieMBWQD7ORTo8Tw5X
XoKAJlpVOdUntF2W521Df4FURggyMp9WCFBtW2NBaEhIpeKh97CSAAr7ghWL9NBHs3SUgBZpkm5e
HbGO5xrL6Df9RuMnyxIerLUu9KnpDyCmmLoZVNKtsTUKkx0n+nnTXUUpwUZBexzjmPpGhe+kmVgr
00APBnNSIspO9DKGNNQq69O8/ssGz0JULG4xI2BvFdOgNIcSgb4hqPkaL/J06pQ8vJRiUxZXjAxn
dt91ADH/k0yi1eWVB8f12cCSh/iZRy9mY2oO6HHIoaQVdIK2jAmi+kuSVYgnvgm6ZOrKHiHAYZ20
sAFYLdTENGquA1eBDGxsASQV5vcMNPowLmF23M43wFK/aw3U4rjHWP61cM36f1dnFPm2CPwaA0lc
LVFtC7IKVmDVfsymwCNUI3KZKB37ww5XJFkEawqDlJDgOTtH+J7ZxmtqS1g2f7mF6BREy5EVqty2
vHa8skrsa1ZpRQVnjqbn2sLt54I3MstW4hoAXgL3oiDxQ+4u3wUMMLH4fY5KEqmh2ggVsfbahps3
i/hYqGXxaqEz6PhNxZ57y7HN5Sh+7hSFojfaIM0mP6SCqZ6yUxEwS/rXzNsQuyn4HSJfo3ocqshd
ClvlCOiQ16zAeMKM1daVBwgiHEyqyqVzH10r9/KNlpdqyx2mufxGqXYZ9/9bNTat0pY31+Al5SBF
3n4euPhzpryLDY115TSzMSgSNfxhFU0vCvZe3lpdAUZ1ZmPV5syJP3m8ys39zd2ZA5gHKpQwG/gl
Mk1e+2idAa1IKO4/7cpekdaL5mvylkM0uXo0d1M4NpGeOY+pDTO4JuElmgvP86t3oacGppZ7lkiS
SGT7cBYejST8KraZmwoCGPMD5QWPQZf+PODGIGLNssgUO/BZJlYMPqv+0eCF4PdlSwxbnea5a/tc
aGWla/IrO07FtY/mEFi0X9UG41qZKuCMKa4sHU+oAeczHfDAKXEtKwP8GY2kxepZqf9myWQjYRwS
Opbq4ZUXoShcvIg39ex9PmklnJZUWgJYVrpGYJGau9RGkp6QxcPTP8TFgzf3s3o5Ir4lQj177z8A
vDPVZsN+p1frXTxDAQGZeEvpyau7Vy3UuLSosHOA1ciiig0CBR+bzD5aEG1ltULA04dyPUxOVWUI
vN2HKbiyfKBau5UBQpteos7Zuw5vF1rg4Cws8JYKeZ+sNjKqyqhvcMKxszpv6TiljLpZyEq9V2CA
Wrt4rK5uzXkyeJWqrLWEEehYuFJmEHlh6fVMUP6N5pbQeWlNT1W0oLxx9Etbot5rjSbpwz3daENm
VKqNitgnbxAbjmx8tlpEqfgF4VZLG5pmCobWKJs2j1yvDP830UOrr1RnwmW4qFptXLec8Gmg6edt
fGwpipX5hfGAwYb8j9pnJ+0ucnXQ77whWZx1F85CDBHeu9B7iBiHNphgKUdRD8YkI0RXsVZnH8XH
GDAgZ5fdpd5LXatZwaVKrT7M7j/alljZpxRdhy8lkHqOCXXbewskcFt48EOUZfvecRcFfy1cYjZG
ktfOj/PjDd33n726KW9KLlFsdyzaC0q7X1iP+mza0ExUTdnBPCXmBrdfvr3DVW58xs5NLihyHOkb
fb7obU4p6wZ5VXWoIgobBo2pgrlDKzmnESmD9/66ad+KnUs3lecBU996nNVrFBZz/oezlaljmxw6
p45llpfTov56YoW6Yl811An56JYcMFKPQ690qWwgPnkgGKVOICQMoLBPPBs970e8Fi916UtCq7jW
mPMejEfAILs5wRDGEQtyWHmxslgciBgveVpjnlAVQswbtEaq2Ffn9BlqP7Ocq8zV0VJoGwrE6Dvw
ckmp3acTaS6FXH0euRpMT9Tn+o56NKCw7gBl2w9enPKzKkFjl+z8lVBp1CHmBa+yp/j0wwhsd0RZ
gsh0NEuMUrFEwNvOiDl7PxVYW77QlYlZQAISjbXUGmKD7FDaX+q+fvprfBjlhGcbbqcG+CdgC/RF
lm4OdHuBe5yKEupqc5OZS34c8v8DgWyiIUnUTnvimbCd9ATFh+TC5/VBQ3NTxVydg26zhsSx4n49
6qRCNFCQdXrSFNeUpb603fEbjccAO8H/qs1DlFYWtrgnAtmOQ9cgZS7i8yocG2Umev7PPlYlU5hZ
nLkofrMcP2QkCyJnPHW4Q6CVanj6A8wajQM01gu8cCGfDV8VfS7X/3t24TI6hha1tUoqXmlf7IQK
4sZqHeMDk3EBxwIJY7/NvfG49G9YpJ9rAe8XcsB5qGKVCCknHVdOSa/NYSOeM6X4iAst0ggzEYWk
bWzCi9yqfs0MPY2avEdiU1SUR3L9RMbcKoOgForCWtQ3jAkXsKMIQ0lIEnwWnV+KTc4KMcXdfRZU
arlxQs0EQE/IL37BbEpCadIT+utAM8Fz0qusvgQtv5CQqwEQS0e2CjSGrCUcMxTTdf2uM1gjgnoE
aVaKa/TPyt8k8xuLgE1UrBo4yYdZimSETPe7ZaWej3cehOj3GpiLUWZHJCQx14pY8UtP/EXy44vh
R2FhrJ1XkrA1AR+Iot8s3973BqMjPUk4isxftsFTTQB3fKWEf0d4EgLjPadEzLKQc2ltki9+ed79
ahUDTGfPRDOm/d5IVdqueyQuYaD2+5xfw01reGs06/7yHh/EfsQUj2gDozVlzJzlhvqx03jRS1fS
GK9OLMyXb3dBbLqxtj6o+2P7C4tAzYYvtr8dhP9gCV1IFSu7o2eKukDAHIlyop8zyxvCfRuH3o9P
q8QDbM/LM3cyLzbKwMSMjrLWqold0nLBO4U/OfUqqzncYNqCXuqVWvdZye5isc02KakghcsCSuCa
y4txyloNVIm+UQ7sGrHk4k1DZCbkV5JO4wMUP6mR+UDdcxIIGGM2qLwCouwI1sfg7SBdZWI8SENB
pxdOb0ci2ABHQ11QAaZsrYKYSETNLuuG1PTxX/GGlhwrZlCjZqBh6OCAGNCEOP/XMXYSmtXuUzVX
7bbSxFDDsnSDb94FMm3kFuLYwR1O400XUY98/Gb5DpS0pxTj9t49I8K/sJrVpS4yq8NTXc8koEQe
1xCBYyL5eItS1l+HQjf8raHadBqgWcVnuTWbOfsCGzJ1kR2+vRXcwaIa/ZgMxNPmxg3TC+NTY5lP
O7CyQ99h2t5rSDqjd/Gy6H5zOt03BLoBHyfEuttFV49eQrdmI+ytcdPX+4O98InRMzBt13oYVFD7
TRVsEgk6gOSULoyXipxDuqB6h4T7kGPibGllb2tNRJYX0FYVDJusKArm1IGS2nTd5WKSlt/G2A/j
SqoUFwnUepBIK0HbFX7DKOEZOz2CTamvYdTnEr4JTDRSPwr97333HWK9diR0k2u2Lg9de7YYlEYh
08x4FP5nAdhM3az+DDtoIoSy2oRZUtYqc5XWjskDrTW9e4hy5LJp9YP2CpWQFXX3Elst50jLBQhy
VlrZfq8Tv6CGeFa/eDr2qztLcthcV8mYvt4PntfneM9zG99baBbcSx1BzrWTskgoKQGjhoPlq2/D
9hIHEhmvh7bGDbTBu3kcqWwokUZdvldewqofqF77pscdigJaRWtvWiaDwrhfWzE3ycemhValshWS
2fDCqrjiFST6Ab364Evc/UDlJtvpWpyw4601K8mzg4qDp9R5WYeE+ku1q14FIAXyri79R/Jns8uX
vzNsN6i/iGYm61g2/tVL++Etcu1jdxEaHRwCCpG5GBNJdLj//HJBQcQHefsqEOVq0H0WxrE3N4p0
cTqPWu8iewK888eGd+j93R+JtwHh1JEt2+ydtZ+cnzABHfiODnWbTlz9wsl3bIpgUMxF4IVxfkFr
F/EEswA5J+8JinAEfWZNrTB8rD1fLmeUTIoi9+YICXYQIBpEeVBWGdZxF0cG3xy227nmeZUjez2Y
G/Xi9Vja9m8ROLiW8kcp/3aleDSty4q1st/jK+b+/Hc2AH4peGjcUzvm3/ttmawK/0O+1qjQ/E7T
oYSVtGxEWWQ6xZVky4KCE+k/Y80Bm1PrFQOJT1umXtF17U8zPa10XiAtug/kycPTwowr1bptSIjN
FSN/u2CExGfthPUgOaMtDiyh9w2CFId1UjSxDECX5BHT5uaphHJe3n3jOaZjaczofsVDISTgfUiy
7uT0BDVTSkUH/i4nz1WmRAVUXOay7puDwdzEqVgHT/zwVuw4CvxC5vKi6+Zr7qhOfPGCzSvBwNJC
NzstsQ4ymBcmxVd8j9eGHSs8TM4f+3BkCmR9d7RpkV110Ct+18d2QY+9XohQInwQVKDgSBApptyg
1+QCuz9XHC6WgD4LxJ0xrfj2kNM2sfjEU8My8X3ydj5woIxO5kSmRPPMpb2+R8h5WvKITEpl7smM
6rN4NgiPOz4EeLO0DEgXccOwJ7A7htbifjEwr24NFa/RH46TPcMvE8tj2PjULuOdLD5dBNqleQK2
QQa9pXpI+sDno9oYPwYoTClaxgmziWhEXj16ObkDPzp9VJiOkR4+zrAemLwUTaiqN0XBEf988H5c
6npKeUvWFgnHoqfgVRHeA0nP8r/MUAhplN7vdlmikcT/RRIKiaYy2cOgF5c+gWDSt3eKKgjbNDAq
xa+dg+9QMclTrnqEci/UNunSqoVq46Skhid8554i9INj4PwySZMZx1Y8GVO/+f9k/iRTgf4PDor2
1lkEMW1y90TeIrPzRl5YBTqV+S77dMtADYGSToU3dlwnFTdGLVHuPx5uqGeYwOIkfEnakhPOWKzx
+Tc1L4QkZO744m+EXyxQ4okp8eKEMQzIvQyeV73I4oFVxwz+fcpuqw1Hg8uQ/OsQaEZkrazRW3nO
zU19sIPk1hDw5vUwde5QicKOT13UWH3w1DPo5wDyYJlMVekP01NoCQQBOdNV+V9WX8cCxU1qN3ce
inwBROpsy5218Yvdfwy97k5aYaIHuPE1x1BROvPLD4DHrdZl/87+APmsfpX17+QyX4gmX0b7eqyY
VN8u14hYrUbBco8qo/xRFPfrU2mcesI7WxjM2f6fP1KeHTm0P8q8jmrOa8ZMjBJjeHMRzOxRGoa0
NbF40k2l8lVD8aJ15l4xg3dem3G4HPchPsr+OWOntwzzrbbk2/TV8tgyxw26EZlrM/881Uod5X50
cR0J/4a7NAGzl0I/UH+l9OPqInBSqgzkggwYrwujj2v4UPrHpPtkHA0UdlY/jxvZenjSqw4VjcNf
MkISq9OiUofWD7F75nv40c6zjo3YXirR07df/zom1IIjAoV94u7A+JdOqekAmgx3GmNviyvHFKMF
hTYRwBmlSkSKDd0lpRey3CE8MkK5Z24HOQaWo6K7ubowvVOnTNnuoOyxiUnHpqXxKrIiVHAQPEo/
2r2o9VNlx2S0gTZhBBPgeuLcNTuhjT2hdo/8MjLaiqbATMIEg1X6ZrCnIP5p/sWfbFwLB6zw2gpn
/fyXw+CZuTwlE6y9r8Y7sh8F16/feuAHjm5R+KTTNWWpF1bh7YcoOpjS7rTxqBNuQefWpd+8N7Xy
hIWEu4XoWQ+X/AU2/vn3ZT5SEel3dvzYXPjnUP2I0ZKH2OFu8Bt/B4AO2N+GHOezb+t/9GqAMtIv
g3muCmaTu53bOezmhq9AgeVb/PYyDrhw46ulKS2oqm5qDTMncbPVNxEzw1WjuB50XwSfMgFIfoHm
1eO7klITm3jQ1Zx4kr+edCoJ077neuXOC5d6w8U7ZbV95PSH3oCDD42IYfGVALs4bKsfUmAdJPJ2
XEPbOBqCIFmpxMMGwDcJ44JR1mR6zhHtyt1WdtLR62JYvFlRQEyVLzanMqUfeOU5jSsqm2AWZMSM
iA+UYIZ3Lk7kObb+IyELYWNMDg/mzkxRGZI9wVjmSJF4q9pb57/c0WeLqVpsx6VNIfoyosfipoqT
kMe2M3llgCcYAVYxu0jB3+fT8BVq+423BvXkltXMxSLmqUNQl2D5JikJMKhBA5p2AXLjZjHu3T5Y
Kw+qNYFei3nhcbIgiMl2GY0gpCJYgGXNlsOzAXmXlnurjaFdKke6P5oiTWPsSTOzCh2+rQxbEWmG
nhNApFgv+B+4r5U/oMgUHx7NUGsj7OdHU9n0wg1fapayYnbEZy/Uw5+Al6/Je0cg+h8fuDPi3nlJ
sBYceiwfxqb9xVfYdGfB1Tomkbensw1c5/YtYt7SP68mh16rVY3RKTC22ImdkYDrqOutK3w691cN
PAbyXi5ORi/y1MW1d2g0Wrr+boyAILHs0y+pAD6coJ19UwiiVaXLO8irff3+Av5fv7s9G61WYRsN
IbLSWR2H+FqytXmRz8qWnaqgqVKXuA+B2iTSc1+xtwNCPxZYeJ381CHi1JaDIxelI5uaYYvhcsZq
QeKXjRJlLIrfJMw3BQQn7cE+BmlKLfFUmG4lc3QxYk1NCeJWlBP8np8/SSTVw3faFZGb4yW63B8e
PPit873Vh1ToRkLLGggmHHnqrzpl74wHas65w33KYOggEq4mzUhLMeLh1dohZbf+cnjabn/8MThN
uzQRyE1cGg3zRQxn1Ua55+jNnr5qxueFIPwGzeSJm+gRzlKc2DJS1Gby/vV5zk4hQL653ICh7nwx
vlSDBzIgv+rL+bGBI3/eocHlIRqKRL+IMz+ayKFt4Cv3BjnPBx1Y8sUHcEc0n47OKZfbl9u2rH90
F+6pi4Fjc4+Jayt6P+DzdZGIro9nOhrojzIKKtEfKxVeuX+RooeFqXWBq91FMAiVUZajKsOemr9O
A4EtIiH2xYRty7rvl2EZfUPQiLerM3FrpJgaNRtIM+flVLzouid2wFOZqLcH35DYq4x+alggx4Wn
gfQwCeKePzLrEUlA5EOQoUhk5u71YM/VoyWz+s94vDzZMNc8fEvFJSeUHe3t0KmMB7ei53tcIdOc
VOQo/1H+KKOFG1D+DhxtLiaFp+molpinre3BRuURiRajqh/WSl2L9aIR/1jNQiF+ETF3LvDjMNyz
eQtgJRcQxI05bVuo4mW7mpETx94vtu1kYDY2scpiEoXHEw4GUvQexrb9JAez0zFO6vuF0iQTEiXC
5Ooiom4s1p91jikmQnfQJUBap4QdXpYB0pRAM8FlcQ46tQFP4tV5L3P0mBrCMIGkuWbkB/5flXLS
XEs1kWlfSuue8D8I945HZp7CywrWJARjpiECBfqS50i/fW3LBru9cNiJZYJF1u2hxdVEpxOCpDBO
wWp3FCl+q8HtZPCWoH5AiVAFfHE+UZAbVRFk9tMFBc66/1x/SttMoGedhW2Wn2wmHd079zt1jh77
bFu3z111f3L6PmRCvlaFiG6mf+FwTVFrQ/zRQuK//q6CxVW7WYivWQUAYCZpD3jnlsDurRby98Jh
7g9fYYpS5FL+24XplZDCPN8g8EYX3QaurvTW022jzvH64OstUh5UYmGDHbmuAmabJlEB1TE5d//9
aNp0hs3OzpM7dbnh62WNRKTYMYYZ9f5J+AiRT0cmnh366enbmIohNR6QB/UwcoMUubsgDufvGTXn
x2UIBqGlzzvNgkI1Rl1gS3+07h4KIxJJ6j3XWYxxr2QsXQEfvrInz/c2HAKWUac+Yv8m3PqmXALv
fOY7QaLwV5ZvSyHEmLB8FCf7ECPQeU3jl+GvOD3tYRAPFVT9nCE02r6Rps6n6ZqtMgz69qwkzzPb
iMGiOsWYAQnnlT0LUPzjUUnxS+uTmjuf6ed0PRLzcw9holCi/hD4uv5zE5JvGe+qr8UralCIYelg
0ESp7Q3FdX7JISeFPoTDdL06p7lAT4SD5aCxicgjghk/owRy/dfSxPAVn0I2RT86mjYTtOpjqiaC
zJ5+L7GTGxwreWXJwnTKATBZz7w9OiThCN8ocu+t8f5RrO0FhcxSx2tFy9baAI3wfX9VrWuUWDa6
8tUMrEyY1U9ij/pU3TLDetU93FxiQ8FTsSAjG9lIJR9KxGMbKNLULJS+fucSZ4kLltS9m+Di7//N
ibwwjd+GXFqHFJ4WPROu3/jvglImLpQwpPPxiwov0C2aWXjn6Q+txkPcobAJ9+wnjgOskGNOVy1R
W6xJtwBliLUSZCn+yzT68JPSLQCOqm61KQpptF09SjWjs9aRsGedSuIEJkCWEVZt8p4DSOcpHycn
AvrHrK2DzTMZxd2In6RciqlYi8qoLkWWC7y706AvsLb4PyIoLuReo73xEaDEgVl5bf2JSdCO413+
/GgH8g0HjQEmfzfbErWNUqzYpO5HWuv+Wn3vvNOOOTyWYL1DrZp18kn2oem23oUE66qsjxycPrOX
TuKB0hgYblIwfOsLfQdurmqAHwk2EpwXjmrDl3Y4r2ezJA7N6tUZaEMb5H3VvNi7ynxhmc7Y5wct
Fu3suiDvcA40NqiQAru4jYl5k3D6Dljk8NgJ7vu89GDwBF1ZCEKojR93913w4w8wM7gz7gfQAFEA
SPYS12IVhsfUaB86lGSrgtA5NACObCmfOEvpt9SuRaPfHO1cgGj1MCxBz/Querno1t0q1zWEItfC
UOz+BP8w1+LNmoOYohcPBgA24WNvvM7rtrXkQTbg07gWi7mWA4aLZhCv9z+dMurLeQ+o7prJe+0a
Niw6xcTvn/hoeg2jfPpdClF4T0WkAeUlJQgHiBg2TmGXV/BcnUwL7VbQsJEqnr+g90RatFr8G+lK
2uV0MrZwdiGtwZ745q0g1+W3RmMU2s0PZPPrPcN/RUL4ycIgHwz2m03XN9bJba00B8mD6lufCKZ8
TVhEB6AAD32Epxw+W9Ik5COduKIjPLKP7cwQ4JP3yZ79HcHDY/1lWmImn99tGyONvYY6HEdXbCEc
0v286xK76/ImteoFtoiGvRUqYHJaAbP7K9G5afJLM1JsrGjEai7jF9EcT7xyd9n2uF7h1//8p8/p
ABTynBgo+ka2BPxP//Q/bPymSfXSSs+XOMB7PSehuKSBYehMhBQcRMXuPQlDejEz/9DjIGJAssuQ
EBdwyVHtiy1EiGwYQJFX4FcT4Yb7E/8v2Et+l2suGlQYOLQUxuBI3sVqLKpRQpg9TcYRuILvwT9T
ifVZebgQy2zTezzvk2bI+BtH6o/mrrNaca5QzBr3awJlGfRiWsEeJAmWXHJ/Q+SGNgeDiimljnjS
eVAHKIKrzMm8vwe1030db2ps1R9e+XCtj2p6h2otn8ZNO4x237EVdMhNZCJF3h7R3eNzssyoMaxc
nCwMpyEULCLaIjJOXvul4Zo9XpVMdI+LKpJz4eOJAkK7M3qzBZ5yDg0q1k3xDgQfETQz7rSIkH8q
WHd1guBZ/uYiDQA+U4JP76esUyu7HDE/gTZvRYe7MqDnk5FPoWKFEZHXbWApRVBR1olgCV4fxtL3
XxpjEotnsCmBHR4q86tX3FmkeO7YnDkFJ17msCliQ5OglpPeBZggPfV4Vs+Y9oxxuI1QVfgF0Zp5
gS6dxomwWbsR3qdyBbzP8MVwiR/Un74nI4n6i6gb6EbdMXtUXlk1wr8FP669VS+xkLAcWWB+f0lC
wWa/0tU1rx/q3+i4WKFjbqmTdouFLlI6MBwNF0su3Wx6sUxPn3XOtaIFYE75VRIA64J4jz8bOtcZ
z0JRQFaFPMrTnQNszJIQDQ9E64JHLYr9GFiwYyFKOT1LpBt+Dd2IuMI9tpBAY37tij1D/aMb/rbS
AoKyO2zfGNmULeITPVvrf3i18b7ZVZ5OLxSTWJoKekr2zEmiAsNsErZA7R9EXezZYbXONaWzaOMQ
96RYMI6XejYJMG/JRBCeDgGKvNBFgzbH3RmLLQk8zZKPRJWtnSiHci3tSkuL5jkNys7AAUAfW9Il
GSd8Ih6OAPPR34nFuuuQHXY3WyJrshFZ29zyVQLa7Fc9R57ppe7uUu8AWWoWx2AWM7taYj+H4Oiy
AvBOp1YDxzljs1DfVrcHTYXfUxeSnsG+vbiB9pb4cDQ4Yo3om0UBJGNoKJmERDskf1EVEek8HzK5
3zK98RJpz90pZlXT+eY9LohbQ8Tf4n+2NqjmCHja+1IF98tUNLoR0jWvcQnfBRnMmYxOQpwQe7Up
cxTIxDY2KOjtAPay11bMNdSCYaMgdS0ycyHWQreAtEnsQVCH6UfEQbs2ifDAmyOf4mydRD90wziz
LfdMElXwyE4NPkjgtgS/WwE8vSOt3aY1XRO/9i45k1xX8k06iumUFOO9nC85PkcxnSFecnxmsD+3
Ces/Hh1a14B31UGkSCpMoIq5kE7P4CT1AXHzXVeb2piRFeN8v7vAm2YDemIuOZSe82Ue1enjMvhj
WZh7P5co7vX+TO8FMAFdmAlbkC5PVxiMN4B+uKJhO6ZhjdsVvFkAgoceJ3IdG+uB6BtTjewkkrr+
5UnRyVhVg650mE21doDKmm8b9yQ8XqpVT5auex1PFe5YdLmmySnniF5BXHziwNeQjVPdmmhafpDn
rAwB9WsyARmyQ5Up4miIeZ3G99i3ut1bxdwI2hYzeM6zDNA0adQcBJxTUKZF6D5sZ5znEWhOSp+R
0izgm7yx8NQRTnyyNhK5Gp1hIY4aynXjDxk6Ts/V8lsMOxncjzEzJ/FXJuIVEIgGRO7W2Er+UNUT
lrwB3SiIiyIzb7hc7/wnPfjn76VzzD3TWw8aYtIBgZVIXgX0PpRtb1cuu8UjDHwxgDRDs6cbH1qF
OyE1gHR+kOmrbvWU7CqqgwTnMfh8Fav7qBXeesLyuesqqBu7NGgWkfKEpaCHtmti04KlvI8zV2VE
iDadtZ7dHHmpOLUlMEDicmhBQnpicLD+4n/PMbL7mlwoYe8hKf9kjmEXeSwin5DmpLfzFfP2OE8U
kcqDRWqxIK+RvX1dJItKT76RzyaIYLyk5W/i+uax2w0GDyu7/O5J11igZ0VbyUEqEkAKn2M6V5o+
J29CV0B6C35rEeR788uEkdKClh7obrQzITDAN42DTJMJPxG+RtLnzuPIVPkKS8hPR6RokcxPuIgS
0wEjThsn+WPgF1agfXXdz7wNyUTLFw0+mrIvZeuvNNvjPkefVbhjC+Zg+3vJ4efsmeAS++i0iTbS
eZSTOs/dVv4aKYoNcy4j6jYO+bSSswZ/8dtN4/AsXVlyu6OUCj2vCCX0P9tOw1E4B9Q9yFiPN5yC
BJY83L060u6ihEppzXonXCVzwUV24DY8GTtKvmeDob55D538VVU4gX83nkYIwslGJdiHgbtOtbyt
1sAfVwiNVtRL8eI8U5XOms8i3K4pNyMb3gsTYJhTucso5eGqON3kVnOZebvcesgbOZCQRwjjCKC2
+jLujSmzsdHiattHqt/bacK5JXQdD0uYxPueSKZpO0je69C4O1IaKJRhGGKAvsBxJCvJOxGS5HV4
nnZMZsTZUH0+0Wpzdlvu3g99rqCt73AVR1AxDoQEPP9En394NgqGkJOvWABqyCF7vB7OS1WGPpD1
JsCyOPpvrQArnCJS/ZyHqRS/fAQNVYONJrseungrCy0i2+JhoS6FJDQoq7WMOaxosT7lQbZKhSxw
KSVTeuCcZTMHX/NpWdBtguglEU+BQPBEqiArLMcLfRiSDmTM6nrYKW7oo03I61TzQPXRLzvFzVsQ
4B/bAPTFwPUVM+rBaYxNbwJUClZgtnPoBbNcuLyTS7pVMD3e+0bfsVD/LZ2KcyjTx74Ck9eG5ciA
XQmZ603KeQGyJ8SWtB2g2HxP9p5602iRXYdFryV20Q9HiWwD6r/PCEIS+DUgpnbUQx8Ss0YoQu2U
LEmHjhShC5yToLjU77O+/fFh31/DOnuce7DTvlCD3zYqaln2/cU2K9U8GShEWo0n9NFAPtOfqb3T
YqKmoqE1pax73zBZKofnmcB0jWIQ5L6uIBs9/e37rrOI873kj+G7x2IRyIWLqAY8ZqRZVZkqolm/
es7ChkrpnqKGwyrSTSMtRP7rhXgrCH6c+QE03adtmDiM9xVsUkhHkMoZ2gkx+tFBupphDqaGHode
fc1CZYOfqkNCQLigUVBrmihNd1JmLwYAmlQ3u3hG1EqWm3sRKxPoCYD6TP7hrfEzU+VekAwq2ytu
vPe55dgP5IX+FbHK2FDiSqTU9mNGL4cKaZ3EY2krLz9vB4oy0l7IQ4BPYoDylGfDWyhistXfxyUD
9kYc8YBs2bVmxIJTZnTm+ISmnSpep1yiM92fT3rQA2/MEV0yuLY3dsmZ/dMCmjqXsU3/kt5PEh/r
koUdjb4n7cif7bZTgqRwHDBI8No0hbmP6IkQFZTO13QCh3YYOeTZQS6KAzbksGY5dTMf/aJCh/vi
8oObecG/rs2FecunJLcA2FZ+R7mUOnxFXrHQQ2pDYT2QHzUXHJnhsxpEulj4/m69lpzuGEZ6RKLE
iKL3v2rl0f6++RfLJBeWcRZdjpNZ5vTs4qEydnZdQEGUquQLlvzBgV/QVPO7HypAucw77XL2ZWI7
HAfQFsu6rHbNhgj51QxpRmOwH6jRPdJv6xWRmAFpc7KHhfmtkcdl/FPVHg5V7LAYGWLFX2Hip+wA
xviCYgmcwNNH7bgZDBufRoTe8v40UAkn/F1eaM1aqnxN8d2vdNBTYnDqYwnVcjuLBz0kpWo5Y5qW
OVjqm280bRy40C+LHWMEfFRYBpZbO5UmnDqlXWKozZ/PTuHfF9Wl7G9eTtKwgSjYmRAtvxrF4j95
W4awgKjwZ3G5sD47MLxvaKvEmOBrH/Oo9ffvpfCUdlf+bxqiNMmbIedWIuCnX2DBg/cUMhl8vUWb
gVj/B3UyFEozD+Z7h0FcBanOz4uK6Rq94e0DW7WgP2Z8NzErYHgZw7s92GN/sxz7ftCg1MgGpxzc
6tBNL8e1IYGPHQwFV2mM/HZwYv53CDg6NhWUJ1J/q46UqkFcz2UFO8d2TkWV5rayxf5k/rr6e7/N
Apm+QzS1Joaf52NLGVoPOPO1JMg4VxCGAUBXQbill+wZ2FnCeW+lr24IqANCOjdGTsV24CJbfuCj
StQcNycP+pEMeaBz6sV/1/5SUyVfcuRUfqya3T8UYi0bhg4lw4wvL6xwBlf5DZ3ytHDqZ9wPYHkw
nhu508HpIQHrGnOvCMFvfyslDGEcQRolqRcJ2uz3yo3nOLbAaV6vnjhLtfF9jaYrI1yG3oQYozSt
ClktZo33ZHB1oLUUdiaxv9cxzdVq4Hnknni5PYWvS9TjgfSAvo1oFLq/nTUDDTWrKRZw2BzTRjUV
b8Inn2Xl7fz4fw18sEKVBYOHVwNklYYyju7zvs+ZItPgJ3mIO48IpNIF4gDmV2zcPFOkI/v7r7lv
26qhSTddX2UfbcSLGtjNbtDL20onFI5fjvX5TyJyNRoSNZ2mfSGkqWdj5nzw5eil6FY+jMQSSXPo
w7p9KT8pwPfGfbyF5u2sJBsXc+qbL5KfUK/NntmVw/O4Hk43fq3Pfk6yyP9uE/oDMiJ4p4OiXv3O
MOzo1HwlUEkk00U4ywMwTwIAJduN+DBbHSrfGufBj78G2CXvvMloDxmjLrSN4ziNqU/PP9ZzaewF
orNnoop0flFBj5O3/Az1L84+xt6k7e7LRqw06bRVodyhFwcNMUY/ZzM+5s+yG6+Df8tTGhQDCtab
vJpOn5a8m2gQNDLjE6muYD7/nEu+9RzHUvwGewGbKS/c5uZ19X1Yjlfbl3I6fZ1m0RqH/7nZM68B
xoboy7XWiwyxvRIiy30mG3EFpBJu1I/VwG9FRleN/o8MwIDiwPslsM+NNpVShkI7zDq66yx4FVVn
1S8CZMZH6WqPBzK4ezx746Lit4beNZdf8DM4/PKa5NPAls9Q4EUikU1idXV1cxd7Mk1ffS4A4X+H
NecbdRkeBca0rq6PDXfDA800CAksJbunty5IKqh8s0BxeITl1AfkFF3vv9baH8b+eTy/PFxgtsHr
BUg/HSJ8ooX9Kal43GuHuyV+SIk3I4cWY/oFyFVd5ixT+1zhknBYxUmXTUT1wf1KiafsIqeX1T1W
eOSNXgelQth8ZKjEtSgiPk0xzgeFnFbHTSG4HRCCiXdf4+LYjwFdS8R62ttdKl/Pi8ONs/Nqjchl
1Ph2vfzHijX4SksaMQsRjKqfMoE0Ezbh8ViAKXuJjoW8xraFmTDQiS9XoHBel7xE9S6axxv63x7b
o3eN6wvUK3PWh+1t2XdgcEMczYpSIKqoKJGKdaHtAhD3UGiiuUVRhAmGa3XzokciJuqrHn9zDqWS
wJDQW2nBwx3/9QnYvbb9NY8OOvqL/NqfVfb0HuzcQJrENO4hLfirSMomObMsJ8ixh2j79PwDQZv1
Ej+LGyMlQ+RjSwKWzIc+0j4aQqk0e2rYlWdiRZ1Dur2cM20JuYY9BoKCiTmjxVg6EAjhm6yz3HWN
5fj5gSwVhHnVKNg6RhAlWNnBp/Br0sJtXjV1/4mcs6P6SLwWAhw1PigaJA6ARekYm5Z0HrVaR3k5
fLxXofWULWOAQ2DevUIiloMY5HU9xpLL53FcOvJK3s2ILMkKZAbwokTQkkloM7L64Dd4WeGg7Nm6
gxpkAy6eD3ybqM6S7+luNztpcbTyqwMlSrcyIctXDcSyrI1ZgDtxIVsW7Dz2+l3Cv2KBYS/RTqr4
pscM29wYWjA9bWHccHOCNUaWlvFDbfzN0RAQGagJ9X1C3wMmil0SfI8glKs3vhVp25H/nw/R1sz8
E9wRNUCx3GLoxzgEUUFTGB1I/mdXQQlye+I6FuQw8V3ofLLATU8T8F6QOvt+DfGQWX5aHMMXopkE
UjruJeXeN8E2h4mXsRJbBzE/SOPF95ldr8By8PKykf0hNVlkbrmhgpvlgZ+Xo1VNyvjsATRAovbX
miehHw6kqMVsva9/SMf5aP1v7Q5fQnQAvZuQ+KIfY7fZpHIFAnh6DbmW9eMO9glk4HBSNKXWocH3
cWFIlQRTtCQ0iv8TyKUN4buHvWTPjqIX7zFlTN8k28JrZTjArsgVJ7xLNVkR+pjTFgZLf7fMEDfN
PPoJFDsAJXYX88iCPcq0ZnQth3CMLRFKMNEOgRuq9zQ6UInIXRJn5TAzDaM+wflQp4frBzn5JfYG
oZNI2yi7NzzKiJOm8Is5KS288TlytCrmr9jCrjBShpJbiDX7P6HdiTm2JgbJOmiNX1K7l15IXJho
i0rZ4Y6xr6B6aoDmacpxl3hcjsQ3Mkmw6P8zwKb9sl0cif8jBzW+LdVLQMMjrBBqyGWCC3RUbuBY
I6aVIfmV4DttAnnranoR/hoo+cokthYBRz3f+XRSRUP0adIQ06ZlwXUFwn3P2nALrt4fRehxKhz4
p453CleXCLZP3DYSP7pc1WO1PeDXamYRSMng9EpCO8oLQXzv1QNwFJ4dAKT3iewVEzv6oU99eUPP
bbGaWsTwSV9nlA2s8o1ZDE1Og7V3TYRTIYE4TI+LmpHC1ISMQcxLk365CW+e9quvX3ZjZzOXR3NX
S07e6565XVDadkUXS3CaqmtAGOVLoVo5cKtruwkr0rSq9Pt8rJxg2czyH4yzKX0Pj9sz4WVXCRau
EcXiBXqAet+IkzS4wV9PtTXfpwwsuykIZ8mWM1jWnurLox9GzOSo+Qq/AoVJACFzdWDnXD+Sce8Q
sD4uBLgfObowwl6lpEXK5MsBcLHDWxNGuqjmqGCKQWN5EWbBBwX2gZM6nKR4bVTFsIDwKBQamFJL
tog55Y0DG638lG/Kitt1opEkg78AylvY61vLF+TzfGhxkT5Hee533T2WkoK994mL/ZweM0oNi2d7
CFM5rD8hUzv3MBO5zJLXkGk4GBdpIHun3t1obM+NwiQVJKGjYWkg5LXBtjmO7Ym6/yuqDPiXd49d
ErEe6MgHlPJ7H5O81E7rYUoz+xGgsTTy5VvloTT3cJqhaRDBGtm3Ok4nTxeTZqfqyiNMnlfLdTj1
rsCykzevTVggrRlnyhEP+HOh8oVdb11KYNRatb6Zsp6lLP9JbTm1585CA12LxJmW8jSNgiWU0pX+
UbNDH/7QTlxWw+VxUIRgibp8zY7KLJZ+rXcs/jql/+/SxtOArRwPxExECqrsO4U7UE3hFLzbJgWA
v9SlS4d5R8Ag5F2GFlHbGKPOLSkTgaEEj0+9RChYTPnWG4iiJX79DE7aAySBSJTi44xAdU1qdQ9i
fOdMZZgj424oDBi8FoHsCVf/xL8SbhLBzczp3qnGoaXiavmMfAUvCPa1ngmoIaSIhs5ZzerkzX5u
a8OFoA/aFvRmGXTZVt1EXx6fe7HylNZg8tbtzFat11cFvGOqB30VU4G7R0OT1fg9V9OzJijguvla
QHXHard9ULmjB62GGYf7VGc5QT0pdWctQJhsSZ2hMHHJP0fRRnE6RYBYPd//76d91pz2tHsq7MaS
LZ2ASMpL6ecbSyDp8F7+oU34SfCgb82pcw/Y/TR8dMEzoN/p+TvUxnM6u0M3D3Id3VGLD0gtbX3M
9Ca6+hPnFyhnVrTyEVcxTWbaq4hKBSIbTd/8wRZIY4+D+zu5WaOVrVs/4zfwzY9ly8oe1zE2VMbZ
qIap9IhH01ue1aCkV3JCt0u9VoYij0D3wRXhmtSb/mK+IXjY4trSD6NayCm9vBIW03lBuH//RPq5
FOqAFS3bGKXHyMDzi4X91XopgAwcHpYOQOQtNqKp3vinmS9/c0+xhLAiUG1S9Eyu5+jCXzG7BMsX
HZh1ZUliDUXaDR2qkF7Nzv86KIulFmNjMVO6aPXUbGbAmcTd1VpWJ+VDbR/7So4EL277hnwabS1h
5BFMGmnsuIU7k+etpTqg+gFfifLmtDN5lp1MLT/2juoKdiP5Iofh43SktH3XqpdRhgUEL1aWXb9C
yM9yX09t+vR20eQYptt7NibxHBTDHDgujztwVeASBjwJ1K5L4JT30IhqWlA1qrd3HhDpXKysqCfV
0Zr9ZxZf0q6m9pXq5Bu+32RpaVR7+uGZE/aGdgmWnJ6XnzeS1IYsPPCdaMq8uL5jwhxHHxVGrwMN
pl9jkDjC3UMi97DfQDsNbb+HUGnjKCdIkS3T0/0ciooFH4cKEdEWZ+RBPofEU/aTlO0N9m4rE6Zp
VJW10mnoqHlCBgf2yFT0Nbat5e7wvNJKd69/nIJfEQ/pBb/QiZwhsDetvASmSOkzCtQKVVvKt32F
muBjSc6UrNCHc49dgVhDpLkFsPzDv07Q0DX+WONmVMJ5qlLCrEZi1AZt9NNnPTHFs8FUBDbqvgcM
NOI2TqTmZmtuPITELmHjCJJGaMzCFiAgBKFYP+akJAdXPw5mo6tmRrOH+K0L/0Cfim+JHi/SR+ly
d9slESF+7SUXnbzzjGDvob2zUJVZzUakSKUESvUWdvWgcHm+baf6UMuystL0ILuoxLQ01yl8jHO2
hQbmIg+ThD27+62MXv4glcK0VpwRurZHLCHznNbrKrVydxX/LPjBFjQdSDCjamLjliy3X+z91rME
KGeKx3Pourw9qcbWilhJf1RP/QaTSWmDTYa0Ggohw1NPS8DrvQJuMDRaU+nWkO4x9FZG7jMfYfyS
q82m62sjcVSSGbFviMAQTLDEkSVmX+pS7DanL0cnHCs39N3ao0V+irVt+7nfDRDEYfn/S4GNeYBQ
gtMvjsNHQRaPTztqpJaKG7rH8P1MqGiZ3lBtODARt6UQTq/noRKb+cmqbscKXWtDfunQhT8ppco1
exbbuTkV800ui1mQTlQ2RWtuBJowZMPkfoAQ1Fu8AM61sXKngDx4wyMXkD4dNjpMeS54I4NOZYtF
U1AdqrkVl33EoXPEBgy2/pp1epzOz7zd1YgB57//uFvyUInNLC5KgTBX1RjR54+th5vF7jsKMET8
wpNFYJKWE0SZinHHY1n+1eLGcuxF3MYNzAnxZyXF+uOVquLb4eIkpMwZmoSrklDHnlYExgfu/+iy
czbxQI0rRSgceViEVWqG6/br3S6SAD434xS/3zCiiRtrhydQQBOiUSVEoINHSTeVvE9SAZmBNXnD
Pk5L/mwwGatOI4FigaSmQNMZb2DlqejroyMguAoiIrRxZvxMXRKCJ4N+KzYlO+g+U85Ti5EDXRS+
VFYocJ6iojQwJNtXPD2QKHWsfY52CU13ed0Zw7LMwUT9OdOANKGMo+sodOBlAoKn+PyqRo6nvaX8
7UwmdegrdTpbhO/qcPTrUIkakYR762uuZiVne6ylBb4Ag0f6ImTlm+pWizAyJoTfMQATfxk4Y4Wg
PJ5q90/T/KG1k2x5b0eXwQsHzYYdiVyEa81JUWCTdY2JGf2tKPmr8MdppmqujOjTfSytreFSDCKy
kBT06Wu++hWESgmpYrH1AIEefbakzCD1UT/TQEHm+GjEs8IlOuP320Iet6hILiMUP194FI9xTB6Y
JhqRlkElMKUYUElWGdRDV83wIv+lLzSdCQHDib+k893gxFugTnL+xb28KDc6ESKb9FaM8LXtcWTr
WzxbvK9V1u0HRg2DlxO9EzvP1d3Gh4xKqofqdvkgUr6Z0as4KVgsaOCxg0kfeqvjWGVVPEe4Pe7Y
9hhMqIDHXO8wR9/LssaKVJSn2vplZ4a0FxtaBl5RSnwNwtmdfuFUObgBbvmtjhn5P9E1EEDyFMAx
TcTHtaqx0KEzJFbgyDfX8lBgZ4xhSeIMzVnloNubn0Xz7KwNCEWU3EDa8OcNukSoqr8z1MSkFstl
bJ6TI+wgdtiot/trFVhVbiVI1WPOLkXwELyWQeQKh3TJWz4YGQkB4lFF6Kz2bR0+QOlFLzJ9m08k
7c1YB2PRMzbS5aM4nLDCpt5Bj8rXTkg/aO/t6B/MlSgzuk7wjABYLTrdLUBkxRJWnegJGfOJ/O0D
2rJIZ8DnD7sZ+dzgGUGb+5Da58yO20IVRHqS0zE5qLvzv3ScAVKCQIrdseBbVttGV8t5bYvZUZeg
PHGAZ06HgfzYV1sEn4jmU9eSRaAYq6V0PDRWKsFLIHHoTBLL3B4LhGtRkWqqBgaXY/51akOBPVvH
C1VJDG5/3gyoQPghrvDOJzFWKxBUMjiLKQ1E7o4azqLLfe8T3t4bvbaH1akF3ReY+vrmfL4wKj2r
fT2/AtRhcuSCK21k8WFPdTevo2lvv0qK2mVdgHKxGJRgd/MPH66UG6epaB8W1q/uUWbErlTzg+pv
HqjsyXRf6QnLMXSxzLFgm1B8LScCXwosTv6m27ao4XNMqV8CFw7dPD12po69wTKvhIZL5O1dcnVP
qfv9e1eqPINb3Cp/ERusuYQ36cY3OZozkuVaPgzMI2Flj8ZRQ2LMqiMV8V5InMikY0crlHsfqore
a0yRpC6Sx06Rc1gwGlk4yTPU0tbPCMjPoUSAbCYgMzJugC4+8oBBAeSda/ppZHggzBHsa67cWSpi
tpCwQJkqrVHCNlAnwzvk+CZR3nVOQpiJhoo1e3JKWca1Ga4bgp1WyGqJoyX4+Ee5dfsEnQQ+oXMs
RYmuvV2OxVHt6ikTYMVOCNirphp/KMZeKuP3sj/YY10htQtGQ7KX5q4Btdl3+SOwmUybPwWOBy+c
5oGjmzssvk5b806fKdTUUDn6rRCR6FmFMMbzU9eOkXO9t6T2TtMDRbgBPR76eQtnB610n37B64rv
5LX2h4Afpob/AWjWEVo9vnr/ZmAd03MGHw+BBkaVUD4L/qSvB0xA7Be3/2PE6cqABci4CSbB3EDl
36v3dK0p2pJVw8otdCGLlJIfgKjEgEktV+MTB0jsJk81piHoAH2uAH0OUJtUmJxWeUlUouo33UGl
HEjLmkGhUvJt3TjL/ab5UeuczSSriWwXwIB4A4DfIgKXRIGpxqCxKfqskP9masABqq8KAMQQcSAH
akUWATALCmDXIg9RYhyeoh+9LOWGkwQN2SRIgrCVDID9g4bGr57Rzh46xlkCCiXHqljgsaCxk+eV
rfPTRipSlkfOzS2J2rvMtsvfXcA861eS9QAvjyWMuh5pZIMUyN8hKZ4bgqxGYP3DUHLpE+jjPYO/
KtfBVGKHIo9WctRYCokyBsX/rssjeduxRR1+ttC7hWx/c42C/3vsOydTbvYkix4JFFRdWw/EaIVq
LRUnj8FGhiM5PRM23nHVO2guiXnBlbDTdoZnCF+BX6lIc8ALFpgKW2vqstc5nOYCs2HyitKgl7Gx
5hxZwhTHzs/HV+zJEG1SDC6rbSxXgXKo4LAoH3qP8YHrmuJBd1EAHXftE+6MWWjKA9UeBJeAEIPx
PmOXPg3HockZIxuphdu8H51xYvPpMVSfE16foT3lso6b8RNmg5zSjeEQhmVOMxu8m4uV86EB76b+
5vUMiQAuQ8szD5+RbL+VxWQ5LCYMAenaRHWSRdLNMfr6bQk+actGTF8wUNfeJv4eKOCkVwMrFVP4
5KD/OwvKJNBahuwCD7mRibe/y9nKjuDL1Uj72/MuWrG3ku44En6zE5Cz7rkPahuI0BuMRw3crEfC
Mxrzfj3RZ8jDmlcuwA/rjG7UstNF34IficYaefiB1AmwYRm1q1LDKBEqxNBQHrW1NszI3TNKgXXq
2qOBXcd8p8WAlr8tFsc2c5CNfuQdDwEZ6YdsZgyfLgDE37mLFdRiHxyleeoIuDzjHbDvQ0PmzV6v
ieYbgcWenZcAOQcmb4r90J4bqstCaER2XQBpPc+DNwoYvfSRbPeuQscF9Z+rDs/PWTU5lCpkE6WG
yOfGmVA7yiyeMsV5ylo1cGeceCTfgGU47cmVK2IptXmH6OOTQ4LqQZeHOF8ioZ8+iK8X9SqX0QlT
7Oz9+a0zjvt9+hYSFcVAnkCDRrsRIEPpxVYaLtyWxEB+H8Px9VuiAJZSBW/5M3BpDUzF0Mr98jc9
mmrcUg6+bSDX9GQABsZcE6V4hB+5d+0gY/2cmlf2kQ0Lyb04JGvtJbIuoF61BD7CoAUQEVMlFDSj
BvW9TC+c6NZpZLActWRICrefXrPlqLPirjvQr0i9HHci1fwxQrhUixl+wYRAZwpmyxeNj0SPhTWd
t2SrQ9sPn1JRoEQ9xGLBxUR4ClMtbQG98w3EkqccBjXQJOll7Ysn+YGboxAdF3T3Kb6NuqMkv13L
t81h02TXtyxUgXa+IbQGVO0nfxgNPO8S6ZmzgC6IjLkmVgWDFFZObXy0h5BoiXd2pIeKIKLCDZTa
7w/6olwXtXX/Lh2CtxYNPfvRUraJ8WxeXiOmGpsa9nZVJFpEZ0ApWICnC8DjgF6wF1YBxEOGq6ZC
afPxdq2/cV4SUAPCFb2QWKWHZLU/Tq1bkn2hcsdc5SjcT/f9M9DIntwTpjEzS51P/i1o1cxAg6JX
DzJA85BCkGxeLA9arRXHw/IPJ34NSrepQ4stuMvUI6Hk9EdrFedZRTc7LJU43EaBEx11hDmdABIQ
fYYi7I2v/9rW59rZVkAnDafB8JjgEmkTfV0DYmXCyoS3kErACcvJhNEfVJ8KOQjDYFQIAzaweatk
hCK45IpdbA931F/uYoVzv2QIfmJhRbjgjvXQx8JjTem0mx9MPbMv94Ppf4hbE60avFFVkx1r8t3i
01ITc0OQWDCGAJD5JW3drQFv0/kGpzmbavC6tnVankWL6n+UTEc0gsnx4rm+UXM9nLv+s79D4XYH
ympxEJCNOHf86P3nA7kSZSpSgJOEgre6/n9dW0HGxCNV9GOye4UrjFQkjSfz9scKdzyX8IoWgcn+
6XxwFtgjUevokOtm1Q+LfS9gIDpUiXwgP/BBLHgbMNw5Jbv8VgRv/qzkCyxJ9A940EnLWTwT9XeV
CHWsPjoheje2QiI9bCpCc06TOMHmVpDAN1j9/WF9osDAl0QCKv1ce4dckiPPjaUlvdBR3S1rfXa0
yFoB/mxI9l9fFvWyp3mGGHwNkna9wX3qDLV8PFuDx3aVObw1/9Ab2Unws18g8HWVCkSnrLbhcOFk
rneEEKc+GL7eByRT3wpa80FOGkZN9lxcGLKJ1BWxLe9u+EY+P/RPy3od5jro5ohNCb+iRseM2ZJD
z0B5s5OG2uz8bFsq9lk0j+DauuDZhDDgnmnC1LxGcqczcxci+6GQ9AY/3FMt67WicUJaziJx0Deu
msdVuqDD4ssKVaHKdCItFKxhCnVGnjqsxJnc1txbAnbbcxOJVP+A4jVUrspLsmVYB52FCpuS/ncN
J3Dh1eze/gRY6RhJAc3cpaqZUsm1Ivd+xH/TwPhi9bWkOEM2Wv3Yc88FQytnAd+JDZ6BZvQsg8jT
Ur2TB7z77nPK+yV2Ny+npSYpQlblnwfvGVOJ3aYICAK/eYZx4TzEey6r8zBGbRyjtchgH1UuqwaX
D3ktBrcpnh2ddSjwqb9n7IiNp6Ue11ncebydeNiDT+4FT8BWgM9Gw5jaNpuwF3WlRjJEG7Na/K6h
9XtO6+QInIv1x7ZxvIx5l99Ixcdnz9P/zS9/Qt3VOR8ms3eM8F5/um6TeHyv3yN6XOA7OLpYw1iU
xDhaSUAwcBVwGI/kicQtDPXlLMawVo07UdfOoSBeBIonNaAYoKV/kS1Npm4c5C6H7VNIw9b+XDNs
ki4e02NU2lAajEAnknzchpJYO8rdpGxoYkeNY2nVYhRTkyJu1SjcBDrf7rC1qLE4BHQeHkTeO3XI
AMvI8D/v+e7YKtf6APFnODctRVGw4B+Poab0is4+A167dU3L1CTBRhZs9QjwzRl20azLUQDr68Jv
rhzXkLHuHgo6nvHmFcQXDsJcfprChZUf+DsMAZsQ/+Kk2LLMBVL3C351vVt2FuWO8+PJZwbF6b9a
mtbTgk/L+V/cfEtx4EZP6EJnpEQmiAowWdQZP5jxqwFU1Qd8aPHemeNddnj4o1zRBXSHcbzG2zcT
d8KKOvNmfx74CMnZqT4p5x2VYQnfXOMPapHSPs/8YWRJ+MJizUc7P9ayhhh3cWSWqFjhGWWlZRro
RcF/iujE8wTmBwOM2wC5rhWqtTMnTaQkEiHv9NW4EzjXHnPB4V0vo9rtkKtg7xM7nwH5yqj1F4U8
7wLW/qbnky8HAiObSXv+zk2+co16J3MJM2N9yPxKXQxcZQ3E6dKy2EPLiO61JvEZP/KV/LQaD+wg
ZP0aMIPlZ5gWryAtGsJ+dAdp0r7zrTSzsDQjnRuy08UDyILcDfd8mt83pyGWoyWzqErTuiPECKD5
gsJ0TWf5LZ1VbGBl+LKO2mRPosJiyZcfAbwpoZFqlUyHOHfbfgYjf5hLo+lhs54dVIcdFqOErcRK
OAdJV5Qc0d9DCZy84+6iJmdnYYbdBNG0DLGcqbFJYsQheDCBWwR2gzO4XQV9Kqr1A8+o1Y3uDJ+P
umO43RJ2t6Iooyextv4mmxKir+ItuAi2+Y38sXxzyCSY3p1L/3FPJJUDtMtBpHSJ9oUALj2RXtsD
WJJ0rBGJfFlACzuwLzwfQR8gaAxWqU6JiNtzK19BLuMfbhe91R1yjCEc/b3niEMA2j684q/CHo7R
5sDV98mq8eHzRwDimkrMGrfyY03RWYJgECEqR+8IFWMyf/MPj6GQf2JILz/Qb0Di9FDte7BvWlEL
6pRdhUdGjwwAiZ2tpDCQQZm+j3K5pUiHgJihx49iUDRllXS5rhnbc3XdmqdcbfQMrwXTxwDIgcOk
zbjhqClEjUKP5KWCVN2d7Z8SMVZHpW2YVJ3lUpCDJzWxfRyPv8+a3SQl3QG6La3RUUP70FOZQzG2
YN16l950kbgQrCVeAx2p8/oBRfMlxSrYcN6LVSlQ2d+/UCTXuNJQ8duzohbHLgjRWskzKhtqshTt
xD/SYqrEXUcPTrJ3KOPuBJiA3qC4IfAXVQhN6/cbEVgDxju/uieUqibNKYlXez6/SaH5N852V/eK
8+0Seyev1w7RPrw9B9cMBuhkn2rni31VTmlYLH/JehvUuhRxv+MMNOi00wIbueVk0CX4PTlH7zzv
UQSE70JXSKh8GWWxQGldnf7fHFfyie0JcgZDFjVvs9h+Mvp+yxiTcp8rs9wT5YmWLnoFFaBSpZo4
TFZqDAqiF3gq5lFo3qahDmwOj7y4lyk7EY9BNImszsT+c8+zznjDGQ4w3m+jj7+81DwlsIbqWyFf
Gd7fIG2AZnEwws8j1RQRMAFGWau0/QUx6cRwE3Gg+T48Ovk/LwJaLfdhgfyJqPwxkxIQREf3CLdH
pqfrPBmRIOuXJBcK4km63F0wFeRH5hth1XR4D1wky8Yyn7MsjAc+mGyUjNah5RcacRH+XUFMQz0l
Ts+6317CQVTA/NmuBwV1fhfINa6evwXWDjCWdV/Mt/18qN9HC6fYOmsnjAzCe1h7mWctNowzIyb6
Uo7DS45J1t1wUzDkl2VxnHwEG7lIgJp2wd33dILNW4whBduQMFslncbLcSKYTUY9NtLUhQv9sZe1
cOPMpmENhH6CK1bBWVHV5kjcub2eemtiPLvM7Td4r6hTryTx0EcHngKjOi9I0YHBtjZx3Q/8Pp2v
XWdFyVhcoxXtceHJYDp+hPv4Cxj/JTgsqezS7D7F4zFPmVz7M6Ndq5fzMqr47cCzOhqztte7Hk/i
0YVx56LvgiMRGFGhSE0bB4yq+nd2hK5yh7gwK7kXsXg/+Pl0vsrYMFCeu3B9NqELooukwhUea8pB
XfeSFkweNq5wkJE/Lerz21S9ufTvhHDMgDw1nUZRdMhexmAUMIqCGQsp7w13CyHcK9e3o+htaGvY
uNsORWBtaiqrKniHLw+aLgngxLGvzn9NOlXHwW3Eh8RzpdPZmp1RFefreBGzQwb/XT/KRxjCMtz/
40f6c2bX7uLlnPQqmhNlEzpOJBjJBELZuXIE52DgCACZz6UBxKPtiWkhjE62G33Y1u77hQN0WqEZ
UFXi1hIVoyKpVWOaEmiruMPt9ZYAj6YYrDDMmETS3TVbx/4vx1iav1x1zGZ3eI7T2o6kxT6t0A+x
VYeFtJcDzn7f3sqpDJGhFocUILGiEmV4inQ8NMRaXBfun8gZ1EHS7AlWxnxsvIdEUZtzE1tTjvpC
KMXiboUb0yvL91lKxLJUWKcfnd9mHD2Q2d0c6a5DV0AbTKVFH6jqRa23t9cqxbIIvXdUJqmIUcdl
bZimEXx/qpNLMYMESCGfREpdo4svWXfoKa+eK93jpzU5fg5Nu0ZA1zwr5ugQHV4xY/Rff2ZzVl6S
p4MkIE24A0Q0VFZ9mDy5iPi+mBV+YB3+QKTC3kypx2WFhXXS1ucNeUhkQhFHkcZ5Hh91gk7n2U7F
LS8rhRuKcPr96nsQ6eYZr4iHyXTjGzt7uXLruyModnHQWE9bcq10t2YTqybwlCVj5Yxvpl5BEpfI
/qk1xgMzmgEbdjKza+9fOH7eQtqY/oY/gofU6aDl7GlLeUoVp0GmxE7fx8i0tBfTL+5gD59AKLKR
jMZf7ozAoMYHb1sVTI16mSlCEqOFEuQMekFXyW/FeTQWZV84gDUr2rzBMAVc4VA36i+O67pNi4XN
qQiZcZFmLyAZtAsUUxWF+Cf63gvGXudJHHRNNPUmyov2X5VGXvQqJoql74/KM3iqH3XN0j0hSVc3
pg3Qq6exMYlJ+XuvItCrP9kSvfLUjX2EedxMK9F/UQomiqifFLqOE12YOLXynpC3h/3PSDm2R5zE
w2lJF8qecOjh52uWjsx4+wDQB8rqt/vvTJhyg6M6LoAEfXbviz0pnUmdTU/b4hWvROBKRzaNrlz1
jo5081zZZaS7b6nA4mg12VlxaK8ZDl7HXEMnLKp/RZnjBFK/+E08htSSqnhdvP6Vb5GSJY4jtqO6
cX1+2VkhxN2KZqWGN+tKC5t+ptuOyJMUb3WpOSvF+RwpVjSmdFZ0jbwu4BT9hG/+HyPiDhddKduU
1vJmyhNx8uW9z/of2McbMZl8c3Sco56kzRgUlkTofX3LzQLeHU8XQVnXlA7toCy556LfOlZ45rIe
UVsexFjPrYwZvNTd6omZ4Gjaw73fjp6dfJbTz7TFEShETE/j3xCgXTyJQQgDSAB9QwVbTEOTN37h
3xYhuUilHIsaCHWJd23bbLoI9qbeCjnpVTNPN6lfKqHP6N7RCQSCMRwpCEpPc7N6gZk0k2YWX7lg
rd7rujgt0xWkjZU3P9oNXubA9pdsJtviyqaLu5mj7K3/Q6w/V6rmIUKswNRWGZvZufiX9ovQQXh4
6wWT12hXZJfh1IffJ3oj8O+3Nmu2Z05MaWCM74+URgzZLzpR0s3H9dM+sR9ciBueP7qMRxtF/n45
RFXkAtpXAqLlCMLmUL9CsYl0EALxZOeVFVM6nMh3QiZ6uMTKxQ9NZ7UjV/Wg/9FWyYH2D9M9uaB0
BaPx3wtZaWoXIP3q5mAXlluCy+vM7Luvo7ZNjv8U4TBpnrxWknKXa/UWOYA47rNwqA0yOl57aHvb
fqBcS416d7CGf/ZpxGkaPlUuOTRESeMh+kA/aeWLGFcHNMEbFFlnuh9t7IDxjHov15P6mvNASD/l
CXWM4ApbmoPRgrzMHFpCuQWSWqR75XQYFzupQz6QeEOyNbzb8G5PKdLas+HqG+B7FOSbPcPP+v3O
SvAZpn/QypFS13nJzAH2R3k8QZY11b+IjDa/pcLntjyzbCHhXn6dQEwj7ERc00YuHwkvLWU6y34X
APnW2y9OBsScz6qbo2jd3v1wfDFJ0K2+KwUMSyfl8kWP/GcpYgGoA86886f9IIove/S1W0qcE5Zz
dZoMx1rWCCf+Mp4GsdNi/p/Hi2se31P7J/3S9EcDiUbc46Emj2uqoGrIxqUeFw5yEH7D33zV06x6
aa5TN2akiPnMFYHugBYhwNFhHKC6642uJtEO6tZS4cfs65aUBlYyRMNNIn42nwwnUACIr3VgGYQg
Wl/+SagcVzOn/cOX+ESZ+1AfwOhSvfkDV8a9inAhOuKNpO0Iulr8H29U2jKXR/256BtwBePH53o/
auJKlzwuG+8sWCI+NBpAK3KlixDRQ9QZHSe/Izs6PhKayb7LegjwSLChe2wQ37jHJtdsARvWS/ya
3CB/SJRABdghX0HXL8noYanJ36FUbbz1B9/JllKRHM/gtba3aYvsqv7OPep8liDBaZeaXYVda1a7
edckyiGOcdogYFD6+BjPvLi0LjHSF8FjrmY9rwfbd72FB2BXZvLWMcHhlzoY2R8yZStvhzyjJ1me
ki89by1K8tiu8q38OjjQKjp2g0hHKu4pRot/f6aN/GbhjM7iqNcCBdsph4KD9mhemozQp4oSmYz7
8BCnREz6KzuJ4spinZu3q7d8FzCSKTQI0uZ5aF/I4Aj4vCIUXZ8f8gbWhV9wSRU+8RkAm2Vr6ypZ
EuePY4YIs9Wv1ShemeZngpvyduWRI0YOsMs4H4drYbKiI6abkSdmBxCQFUpi10mCj6RMyiVuLqDq
Zd9GxzwDGs8qVsBNMaLLL6wdMZOlQhz5GZBa1513RooJGXWFeeNak5enrQVTryRUKorsJZczTh1b
KzNXb+ACfVNXZKr7j8RHweXs4FyH4epzD72BWjDppbR051isi09IvF2wEDYSyCB3AQKsKdaIHrVx
3ZXaSJfZiC8FyxFNIIr8LuyPJsldMYwYFKA+c45pwyVXW9qTcmIKjxCIdLz6aCfFi/u5upwyqXFP
5SgCc/wgqWz73Jmt4DJt/fiyKkspvYUZ/9kA/fGPO3KYYCM9mpOJxolb/vCs4ZF2p/AOxCrtEQpW
OYRlx7Uij52IhGRQo7koq9JstRlamxXH1oLpEEaZpQS5IIcJBaV7cZ6UB6a1BrB4uEizQbm8lUb0
pMMgDkgwYypHtyV3kq1NJYiEwoi865k1L523/hxFujbxPypypVPDKS1E0trnv1urtGucywjcQ+2J
N5cRu8cOBTLJ1PpDMXwMMaWUO/zO8B7TuI0ngJJLQyPAmE+cSZ3gMubRvM/v4zHKKGZdDdrjBEIu
7Ub/yFXVUupH2GPuO1sjz1bL9o85JxbDWozHcF396LoaCCl6HOWmpX/Nt3Ut7/2y7Zt1aKkLcDp7
d579nxdOo6KPu6FjqcoMOUuHBfIrAKwue1V7iLsuy5A9Rw7k3NebpT6vB/DE5qtzKupCsuTG+59/
aBEzkXb3q+c4amL7OU2KThcVEhk2I0wXUZ/wi03f4mNE7MaWkwvlOPhCnWR40vB2L7FHfWnB3j69
42VjSj1kk2XHj5omtQ6cGMH0NSAbDZ7zRqfqs5OQBAdbT+z/WoALvX33d8aYlYez9zH6cB72OBAF
yd5Mi1BcLJR07Suikk7ZDztcFXG3FVmvDePFLJgrlNyLn/sB4Kmm5wH3itbzXhfymcDgbEHnRZ0A
WTQ3nVdZDAjOmI0j5e9QDldbZp+YVfq7+7u+luhl8GBAegqjbvFfIJJQP0JI3KiIazLQMl07W3tf
Oy9hnuIwOCuJy5VrjUE7d8wmXtLIyL7rbHcOfaQixXFVDExD+tWfDdP5KbyVxFl7QExefa9GvERr
uUnfVCiXtJJOdgNCftKZPj8n2jXRy3hzXk7kbL+KfMVlBGyFvXiI7T0GwoHJktKDD3DUazS90Dwu
YuCJQyUes2pcV/enOLIUkIz5DEOLBLthql3tzcPw1XU1Ju5HuI8jJOSyVpa4LjQT6JleY4zvHWjz
IJ3+9e34t42XYVcfUt1q8YkRyfBuP+5a1j8ClWaGDVDKd0ad1tYt0YU5ZQ8dKDQ1R7VrQDp9zpZ4
uoyfcvT9DOjgT73i4m8srKq5401cHy8/p4get1O6As4DKjXbmiqbCRYeE3FEOtlBOlkJCxMcQfoQ
24Dg1gROTaVCP0rBWzehy5OvCZZIcyDbTRiFtknNyWvbJ6RblpTJ/tN+ZjEt9Xx398KjBoImI30C
2RxSHhRbe6cVxWPazbSqaFX/UOFEzQ2XWeP8pgJht96GYzGvsZW/UB6gjEzteje/bXIdliiGXf/2
rxSRm/G+Q14uc6IQjgIYP6YHUUVX6kRexWLI3KfF0ihw2/ujlW892fpfyXQ9fjxH88UG2eX0R+3f
mP+Y3RbwPCfWvECoV/3iVNVNhTV/VDu4ASo8gf/Lx7tE7PJh4iiHyjXhkbPj0uftF1yR87eghag6
yOUntpPv4nEhws7VOQOXmh5feuD3+grLUr2bXK0JsKgIQOLcT70uae7c43nbOTcFbNbtNAN7dX4U
qx9UHl/ZXL8y2Kw/hJsJcvnyUhjvOF2AokxlU6ExLqOSJllxpiW0RGNZ79MPocfrWCbWQc+48xtv
nRFb1M2gahKRI7hwzQi4xF1dD1z2+21zU1SscEkByEMSXBwSqHymAUBBvE1vFKoVbk+ft8MCe7eA
jWmP0Qoj/fyNhkUydvnKOYOtuSUkeTJiTFW4zNhTOBa5Pzfd42rxFF/NIzJHuw/z0e8MF0zst/sJ
imVpswSj+cuADmRi6dojB0a+vtmvb7zqE688+lUNyd2vxB67oImIMo9q1ZwJa0igJZwj+XOs5DXS
6TBkMP/AlOIS4fKboa8CuOy6GvCd8LkHN4PaksbnU0CuRt07a1V+GED+7fvAvQtFBqgQQzq5APOs
NiscJlmYjiToaWq87s5F3JaN4ul5f4ha2L2WrwdOUqmJhWslC6KGNBRMq+0zQv93ZJGuknEUbQea
xCwJgPC9VKp3eWzfB1GRa0W1seK/u+EKOEadOnfh5jNE88ohqkt+pmy0p2JMmz8c10YcpLa43XJi
ygRAYTUsuyGxbF5Gz+SSxIDyv9Pq8qsFmnGxuor3dI4A1dXOCE96HdzD7LP1d9bcas8ItwiFjZ0u
ZK/k7J4m/hPNDoxy/g/Bh9Sn8sBRflKz8cJ4juDDrK9lMVhahjLVrqvsIg54gjotv+ZL+J8IvcwO
t/9RnhBbN2WZLEuSClMneOs0qZKlSNnrJUvS4Dw790PPFTtHE3Oi8JoaurtxJwnGf4xmY90nx1fq
V3R+UIeq/X9nbCdz9AHYMpM25ntNKWMpoGbMTKUw36/n8IJHdLpHsO5cVGQB1RMdubQIYby0x3f/
mH5zEd1ELy5nuFZ7ewdosajTJIvcFxbNRHOgkzZtNJIrF9i9ukHSd8ZCViDBxo12SFKF3pOxakgd
7TMQnRf5uH+G8uynVGMbeRebRopvA4HRYT5gS5n9yBNVrX4EQRDpfnfMnZuVDp3QKhA/Jm61hfEB
F+NNhCwD5QCUaNCPpszlyxLMR+plSZv/37/MiJWEJkKTVA0ZjWOkRPJfryogMhkcyMrD68g47C0i
ZCZPYnOqUM7VUjgaAVdjZRmivJGZsLP/twzYZeiyWqNVjbwLQgF7yJFwRuWqrt1q9bskwXlydqtJ
vYZYdGohdbk9QF457ns01uUrN966OFnTb1cjCyL4f6Alv8N9h0wEeSqqTnClpOQrM54o/mtoOKLt
wK1LoqUYOHhipxVScBEaaazBEAscYwdzmWf84pprl+uzZd23Qs10fv+O7OpB+rnBtHKA72qk8T3u
cV/oRa0fwgR1L42NAvkqLDxwIa0Lob+7cH9vqddiXT1vNwNEqAp6x37E8jeLdS3xMwobT2JZkdiO
M3x4I9/MRsabX7EUlE0blUfJ5AFpTxQT49TrWq4ohJWzLnIFU09kA2Laa0sKzFDS7wfu8qTVbN2E
Hiq5JCG/CdIIF2pvOb972EaZvSSnMuHZsfuO1e9GIZrdC2k7OS85t+cE/Eib97D6PHwUgSfDtH2J
jEuH0Zt+dn4t+JLvoM3D/w1B3aN35QhTNZwd0jMGC+eBZ0CZQ8Zew0gayuSxgWfmVw93pxfavBK9
73vvJw1/B8gBe8nykOgH2lLRuxf2yz/rKTSsyTeX8IT9y7gJMy6xB6GzByk9FnRIheTVBb7tl5vX
TDPm1+6E0CgGKXK/75lHK1UNUsJ5T+t1n0vYS6/Z6z3jKGsV5SRdGgbUL6WufpO8Bs6UknLQ18xM
hI8leyYOfkwVLdopWCneGYTpB41NvZeBMSneiCXTx0vLLNJxnmV0aQf8VoQvb2/hIu/TQtGN6Ue/
k3C6uwc/elzbd90H1iXp0giBaRG/QFfBDbfQdp5TUXi7uY22uVldXMUhj27JqALQuR3bklUm/2YL
Dy2An8q4/OB4ruf7EiEYtxuzrY6DTS7xQuwhIzGEk5US7B2kGkZFxVz3Dya0WuUjgObqEp2m1n7W
CqrLVAH25VmRnpHrxbzECIkESVlKKa/Cuw4NAapGXiAaNJHa9HayqFwyrP5TI1DioUFDBta6xyHv
XFhq5Q/XvloBs7KY8LY/NdEWCwMv4o9YxaWq8UoXWBqoKxRBIoL+hTKpzG/T/msqmY3eb4Gm+J20
JTQdO18UwOOK16PrXzwCCFeXZq3Vzs/FNOCyhmwxIamBai/SZLOW8MPPQxaZyA7Dmlrsk8r9Ud1v
+7DRet17uN8SSa9MvQ2fPItBz5PJprgJdAyejWGUM2fsWBEe6oD/G0Pkurxx4pVBqcb8pu3NWWPJ
mRG1+Cff9c5LJRZKvdG19K/Eqsv/PEJy2tlqMqQVk1m/ikWfMzowgabcZHvgxP5drwUNqzGPIbht
0/9HxrTsWhjaml/0wE0CXsRijc0Wefm+IzIOHRN9ABK/kVfS1mKjlPUekfBCRfxGlmxUP/4y5i41
E+HTqixoiRCnYCRBHXNhLclt5vK2b687ZRgqw2UUcomJPC7LcHOAfAW9SRiikXlYB7zEXYj+HRUl
JbJcRxN6jqA4uysg+d7tUoKWnG1JnPiR6UsKGEReLsVG+rQ3G4Tk5UsfGAKib8Cd3ONEKyu6qhsg
/tJPEITzH0EO/3t901itb1NKn2wxhSEH/IaqYv1szZCq1iOpNyWhguNl3VGB6VysKMbGEiIh4uQQ
POHk8lxqEMJBwSgLR5uJFgWZf/iO14LeVItqMOncEqVvp1HgMbYGrjbybLD8YAKgx4mkhIoV80yZ
wfZFNY6+TNs00CYOCo5TkMk87UzbycQW5dHV9XH9HJI2H6AonVTVfx50LGmPVmGM6neyM7XnEltT
SvWxAT81njXmLG21rSeQtEhpXajoTL3mU0o+zwOljG297TsLl5uT2IeUMJVtE01+BUJgBo7MA45V
y9g8c8zHKOjY1OW2vbMBB3JH5LXd3zcxVoPLw3J9RmNNwPgJs+Y/9Zqo1oAPZkDCyqgI+GiICM0a
Z1o6o1Pvt3YediMl/6M1c94i0Z2OBMcGpUm9z659xzIH2K1RyrPuWfynjtJNQjwcNa83qNEem0hP
cDb9TAJm5AwDNIAqoMsBVQd6dnWMrK5EPRq0XzG6YGgMi6Oh9v1CoklSrL89Gho5oTch9bVvDexs
Wht9HCl+Laz43t6Qs48jdpUUS+13stXebt7bFFbY5HzVx9Mql5gVwenpt+8DRPAf6djQ9dyeL7Lu
uosSh70dwwDDX+WrmwVjUNnx3KagOjreoj0VZtLFmZfb2HTJGbkkN2nQDQsJWRfG8bX46rQEqDiZ
0zbAYCpu84t0G3sAurBPcuiFv+jEZYCcvypv32HYRxta84jyuNW5o3/Qs5r49z9Z9Z+50/xsI6QG
TJXPSpzaswhIOgU4Y9GvqA5IDjVML42gHwwgTRpan22jLk1Np0wtLxPN3QdBqzowQVhUAsxSKV9p
o8UI5bxw6sqD94eAxzgP4aU/mbsQM4Y/bSfQlsb/TN6pLs/iY8ehJT1mS4iJmw2qhOFgOPdOzHCz
wSBiUzzTbGFGvngPn8bNZ5axBJC/hDFcy0yR5xqyDCpcz3N/AJUzAR8+hIKvG2pwgTcMIyBwj4w5
pY5Ih1KkouR1/GLgALvG4kwu2A4RAS1gvMx4SDZD74GjOya57OYeroA58TjkGQN5fZJF57DEyaqH
JMup2BeRvuhY9UehYSOsz6SAubyfpuW40tcGBcbA4W7xBB+y2635wroKYKBW2T0kaYTlZY9EAp6Y
UkzfQdS/Unu+e+bHRcQErFwvKEcEzFELWuzI3/+6eB3XD8HQHC/DfY0hnbGUHA2VPhqWIwkTjF4w
hHhiqc+Fdby6A9U+4r/oev8ukOGXLVE5+/1FiIsb9a0fdgX1rY+S3SGQokt6RtE0QlzL7bhzIRl1
iAq/PzNnKVLQBci2z0jhg5GSpux+Zi9VqEU2v24qAeCvXvrdX3WLwsuDXkUT+ZPeD0SV78/MLev6
xLrubPsCaiTVc/6uthmBP+a2iTAyHWi4gYVkYtNBAFB1qiTX00ylny4rklI5mNfL5N3Ux3wzYjuv
Ql6Zyv+5ZBunG8P/C887Vr5lEqr4StZhshd2QAJJPzLDNlxpVZh5n+tLOst0fECnkAXfUijeeSAe
KND7rPomRiiBR8RfBGAwdoQS2a4k8saRHe2CkRC/Exlog3junDCT2fsayHe1/70ijxgW9u+wAyrJ
lwHWKGBg36qpGaah2ovQw939YLNcbvmiNRHd3qOs0V9vMSRj0o7ZTDiGIZqR9o1hP+H2kbB9ndef
B9U4MClLHmlOBZPzna9/IXu4MgFHUlDfx+/R7CE7bDlR1cbOeCusr4zRocmjUyOIBXSJdLPFhexw
3ugm4e83gcuWOOHsuk686Jngnmv9YO2YEeEgEH07HUBF/O65ZHcc9Izz9vcoQFadY8QvOa/OoDj3
S0WSHSUsKiN46zAOzaxH+Dub3weH5eqEo8UxhjUgOZF66BB+4/hhkfQ1O6TxTqrZ3w8A3Pqnwj4U
CukcH90415YUZFmiTiPvIUo13pgptQ3YdRZmqxOTewchkQ7LZwLZlx/gYy0wMp9MCE0132zt4E+Z
aSLyBTXpJES633FZe09PT3L1UGyLKh9lIGFpTmBNDoxhk1lTtNuNNNrF72nhghkdPg1JwfkP/yhn
q4npvwGTojVZaaYN/DAK9MSJ/defo+MlJlUNg6TInA5EikeCWzFeS3y7RmqHA0AEWj6fjHd6CqVN
rJ3C9ITwnToLMQHFiyBys3rzmjgJZ0T3FH0ag71zM8wWdOMlVgztGoik5bMK3euCcA+o00cV+xjz
ugOYclcD1dxfbbgl2zlnIZapyb/mKXVq43ePqZ8LgL32M9NrkGsw9yWGckzEau/+xzpobYpZD8P7
VG3Ns/5znZNfnANdRkQcjVkBNK/2K+8z52aSnfwy6Iwhhw0pMY4HfDIBfIfmSWyx9NLhmv0s/43p
AA65myOTn14+0PzMNG95nhzkoi2QtTy85GRhUOnDk14GxYYiKcMWzk5M6IhXPl5uOiM2FvWNdKL5
VSaFhdWyPz0zBN1IiDCg+p2AqVWtieGq+v2NzG44NKQDbjlnhjICRRIrPNgMvLpZDGpB61J/6wdG
J5BPA/b9kwmwELvXPfpScOgXE2oRgNbu9JLHVekXI5iXR+xwWOMAD6xr/2d4svPK+K31/HDLnFU4
lf8I+z9+Bs8ayg+mmzgVj7fbT1rx1l6Kx9djUDJNCYkvpBAyKTxpZ3+wgU9zjnPzPdSkP+KRFduE
uP3gKeyF/T0ApS3JhUol+wV1BaqEGvq9Iffelxj4WRuFwphLbe+f06FWtW7Hpd+SBqPXesAAKPYT
8XsNlkshXkiwmEo5o7iXkonW3aQrpaaMO9Mn4MnXWAQTbdqC7MMMdqPb2WoHTbIgtqzmoKl3pf0f
8czMowc6Nm7CZ1QzXJqvLufubK/H4IUKXpMVa4yp4sHKD3eyeiJlZswQydJi0DCoS3HOV7h1rE66
lXRcIXgIy6XUhihapRgqhIcwJOoq/so84gfg2SXBujdazA7UmfkVMmm9rk0tqZEiYau41NT6QAup
CyNqXwCjGPb8W70RIJx9G8+6PWfw1gNPqK/xcFezMwwxNjrfEwsqOexeVtCTWt6UvRtvRfBoL8cA
XzP0giy9c26hAJZmfYUZKOrV9jq6EkBWQOfC82RNwx77lZhfKqSYK0D5g8rAN+sf1CIoqEom7+Jy
XT55yvFqXE10sXobM/ej2glK61JJpz/wxqrfXyh6+MDwl7CCmNGqVee90hFDFNR+O0Oq1B0ipzfd
gjdX2mIHwT1fzZq0q2pAV4C5osURJFezDnr3fu3GqZoYU8N0hOO2kqUgsw+pALCipYNOBa7d7ZIL
X6nwnud4qIL/r4ORonv63PMRtP2vGAQRSYaYFzxINSyb3BXSTajDyRwwmK+vEE6vmifuGRSoNhvh
+EMVwUgBEZussHIvBVkBkBWtvNBGSbWc0Wn95Ko64PMdXTdJeXUQOe5V6ILIB3AFNCCI4urAsmJn
PSXKVdk/fXlzo4vkBFTz+X6mlUWyNkpxWUV0Ew7dCRv+Ae9HB+aZXDeTXJqUNjEi6Bl8Chmv63hy
NbVixHtGZ9nptfRToiUs5MUFHbfRnhHzk1N5bVs1ntRWL0EosEfO7p94a0ESAwVIY0+YLLL8vt+E
J7imcxNUflvSyHAAqU81kZtW67FHajlwlmYELSzDSeZBfE9dDp5VXn6tqg96YIOe96U7O1bTKbG2
jrAazPHYKoMR+gVvxfa/NIk76I73b2CTiREY89sgdObRTokNsehxtXPTFUYbezQsPkhkjiye0nb6
yUH4hum/NsJzVvqetb0fr1sLwGCwRp6D08kILTY+BBfkBBSVMJA41tqH24Isg/6XQ0neiKUPS7EN
Ya6JQCgk3t05favQd9ruNC1tn5chkMEJXlHV69kg5tlVCGyPXjrZZpi+QruQtjNNmduVci8frezY
+HeCvrtBExJPtYhMvw10hWsYR8gwj1C/OWbbYPcO/N1SYY2Lzy/aLCo6gFJlgPsr6i6GHEfKIzTE
VzQTt/GHGQXI7QDr1DGqRQf99oTnViRt0mpCDL5ozisnnx8NDG3o23TDgVSi3prekcaYJ2eXBYvP
U+iGqNIQ6u6x8km4bgbhSieoNBAF0oX6Hf0sCuURzBTYhghRyJT6uroIM4leU6Op/Zrmx2aasg4H
fWVjRECEJPcetK8KGjtq7/bkeKHvXlmhJRVUKKefRu4NJdjhIlzG3NTz4fFFOlHmwiazmP3WbxL8
/R8R765j2J+QntmADy2pzdF3LwrbNw0N1QWuxHuH1w6pMYcJxil9oPy/QQZOM8JblGjzma25Kol1
URuuU729iUpytIrpCaInSXUO1QcT5u4RMui9njHsnbx4plCpo2B1nlkL7kzIgHdE/hxucikPEhsG
LDyON1cDKhNu6VMPFNUX3WAz3j3oU0EgX9qg1CJasFDhseAxRS9M8SJOF4pnClVsHWTvL8nrVR5y
seUkV822tHhvuiWqW88U9/vtzQvD4H9D1ytSRKVNann9Bpzbbf+7itop3jhWeSKuM0N2AGBx8rxl
xJGQm/5oHSEj9lxNXpsDwl5nytgTO83cwBS29Uqd/vDm5oosmJTv1ORaioKUsxFTZBiOHXjxCWXb
FVMiFAUUrORbeGhb52O8OS6kLM+HrXMTNqqns/6bzlWgKClMr7DKQCt1m8WQLxuuYq/jWjlaxRxB
XHcDHLBWdmkNOilmAgJalngn9is9AdpPB0on9L+6dt6ltZMW23x3NPFDYgj9ckk/q9YlGsunwMwX
7dssClTyyY9QhCUuzWZ9IHZ91q4VoQXC6Uu0nSPVib2KWSWcNs+1mPiGb+1/ud+QabXVR8tXuAjy
OgzShvpP0b4vGUsyGo7AZNUZEecrCqdZLtda39pxH57E5nJIKZ3wmTJ7rhXrYetIJCrdZpyqQl0G
DOr7wuZ4Vcytb8kFLL7EnObZZJ7gM5RySSfU1eXUTt8rGD/5+4azko+hObBnvsWws/fJYzFLX3D6
nzMlHHCH+OCwHiCRHrUa/7fI0skSYgEKtDtlI+UXSITBsIZZP+cI/Za1Dj3CyccZcnwBoTyeDDJh
7y0/J4O6FDxrnC58J/QU5rwlTkOaxkl1MA6nNEasNlxReUu0gCUJIDoQ55RfRWrmrUsKhBHMphk0
YXxRrRFTqb0UY4QoQIVv1H0vetrATunh6q+0APvy94SxzdtDRbIg9i6tOkEWJpRMhNZk2trQpMT7
uo44Q56iIW2pj63MuSjilia5FHFCPxSR5N3zYG1xEnankJ3Ty5qDIeyL4KXXx+xkGo/Xzvi3pVsk
333vlZ+WMon5s9N5PaPmw8LXUrPetAA44dA/dWtgmqqwh67E/NG4I4uXRKazbhwdEye25e3XQggW
lu81XzkipgtuOHU+VXP653yotP3awbMrSUvc6sruoVt1sKcLChzEiZOiDMzAYSiCwwfHIADhVpmY
bwC3lG6hMKlzgD/BtXEaXITcGKcO5ImXMRyE7w8S8EYWFrs5aDaLsoz+XyQLDs/KAgcGpbMYyOM2
k+COAZsDGCEkjMyT/kVYcilzX+tMIw8Q8S1+2TaFY8QbjiiY5co2gSMYxWFlS7h+vH7k7FoZrPDw
7PtKGdtCdhfdlc3b9wFcEMXCJq5Z70NgA7e+3XeOdmsPkUMSz9zaKTOKPX4Fp+pM8bovDI/vegTX
D9rE2ZC2mPrDPtUvGDNYcpGa5luMrd0RlcZg2hGcnfOhV1F3P9UUc3hneoUZS3qoX7RTyA/6QiKc
JgxG17iolvRKGbfdN1WPNoB+6sfUtwFwY0arxRMgLxFN+rjcrmA4MHAOwUjSOhvFMDAPg8mDN70y
gvnjXQuh0CU+IKI9pJWxWVutaTIRUBWd1uc3SBsZXVhz0EHkRogO0F1WEB4pwXemQjkO4+l82RVr
j7wG7+Md8ihH0DZl4ZLblKLxjWU3BHxZPih2DfmwHS4mBdfbIdM/FoGFTvf0StW5JCXwfhiiaIJz
zRDSF6T2tmAdvabZnt39Cue2o3N2Rag69VLMJV6vzh2H/plG5oOhHc2KZBFGirv12tQE8O193HPP
2+wzFGPiRt5JPBiqerN4ZbF+kr/aObgHXpSg3fUy4D668mtDlZPf+yLz1Jsl+tK8dLzOlTFh21eR
maU+azlPvEMzVWGmL6bOMtaD4qmDkLTVwuIDa+hZNXmu/UHw+lrGCGAFKDun7ALzGpR6mkw0yeTi
kRBDHzv65LL65jICxOTl/Iiz4UqW5XHa3sUHeQQNwyXLBAV4DllRYkDKBLaD3buf+KBlp95HiKgA
f1MJBoJQIbuJjlhXSEwPgoHkqfQOzWzCqDAl5eVPVRcXeDPb4+XhLbnau1CWqZTAyPtyLVbryMxs
mGOb14zieD35latnCRavGFAMBXEgsDJwivLMtUJEWhxIbHEjTDkQjSN6yyR67xLX8DE+aTiflRYo
vsOK2c6PYMOUEo2Zm7RbBzBtX2Y6fnL2T0URevnhStiaJ/S3UOTAPkdq+SfPKm3112vRtAM+RWI3
Fwy7mPhth/cUcUsa1UhjO9UTB9K/L1tzU6rEYr00XEeGYnhWK5U4pg0kyHXayeVvr/dRXzE0wXOA
bCJkN+YdAM8GjIWcDFpQy5wCoNuOL1lGS4ObIVlmGBzcKKpocz5tJRJuJ5LkYCpnNpUv7z1uBpXx
WY8ZyH4U+zhGv/O/yDE5A4qM9r59nvj2QBoBU8/pqmJd8oHz4QSZGaT53M6WU7ZIlWPehL87lw9I
f7jfjc+X5LRenzGP3rJUQ0q7ozX2EJN4H40j4TU0VOOdUKU87rkyRNZCP1MXGeYDY5Oa5qi3pleO
ihwnOHdxsTG/z+nXPQDNfTccEyCAqKRIX7x81DRHA9slsuv4pSUS3UkOP2FJR9IQNN5Vx3Ulmk45
Y6M+2fDnuosc0HPrX2sYVCmjVQT2Y8I9/ai+o5ve4gqaa3Ntp0MEzkDrxePPQfJi0Na2iSJsyZll
SMO5p42+7P8CjC6T2EDhjwd/vc1y4eG6pYtqzeekqyawLxO5l0axbpAEZUWu5au+WAu840WAqmnS
bH5ycVnIKbHGIwCIbqBfnqTMwo3HCQdMr7cSMwN36w4QTFtBV1Jq9804MCdH17bNXSRRl+c0K5S3
DR5IgNImhV20xhsjV2dFURf/vuedsg3E1UGRzLFJzsiY0Bd5oqV4ljL5dLnRVY+uqfZBSZ+o5UIc
nH4eqjXI7iF4//Ma+KBApBI6Cip8OmQga60jFkGW4+GAgLaDKkUZz4Tfxp/UMLVuWPxbGNfY54fm
6rzuPzZ1ooHsQP/fumdOXskFZqT+Zp8GLnizrhpt2igheXyOGWtWdivazYnpZPGOH0nC7K4x3FoN
X7r9CjkMDLrnk1BNkQzBlJRLkGomH6A/c7tjDV14RkEzVysOzUeUj3TkIWa7hhBzVXDqkgt2Hu+L
uPd6BaCEN2ZZh8QGC+OP4SMjhu0hFIBtcgRoT1EMrH2pngDS8z8dknQr90vTJ6gyjty2qnzNDwfB
20ZWRq2kAGPwcH1+txJlU51OLBIti86zMQfs0ta8w+NfVjcOE2yjap8PBXztV0/qtFBFQ0wg0AoC
kFe70Kd4rkqiP9chBKTqzyux8xC8aNp5HjPhC0U+3t4iZ8+KPd5PauWt8WKNsqRolf4bXiuN8kai
m8aWSso9kovRpHmUaVadC3Hx+n8/pH04xzs9pgUPBDsjPH+qhk1p5oV6GQ7YQF4b6M6bLowKtDVD
B4fH/xKqCWyIJT9uiAHyg70ACJrWZ8VjXC3D6dBUB8M30ICP0wBOmWPkoonnqFOVgc91MywXozhx
JEzpUhZy6TmGUaIBIH8j5QxZNSTH3xpq7XwMpaEGU86k53YkEVNwme0RnYzV33nCekY9ptKHNKTR
jsoqMmlTc/EvSSI53Rgt6EBDa+OfFVlWlmyXtYl/snmHiXsg0oO2rU/Wxj0bIBsgB0+WWSvMPEoQ
QVuWxTHZ/ofvQhsuD8SydxnOluxuIDm+GGNAmfILtLfuTxAalPGXxp24ECw4WC4vhMhE4QIPJ57v
IFSmi9tVtR6OkSHekjmcrD6n+B76gpFC86PqxmkQUs3UuZht4b0efHwNUaPOS1icf4LGKhhWLMcq
ogC5IJsqknPZHqbVoVDAUABKibeg2YPGKaTVjfrH7oCI91QTG+SBwhnS4XqkoBG4OZZwQ23ipw2M
IlXMe3I7+7ETmv20s9jCvINxtihB+7kSPZ+P4jMDh/MfY6lWrrjx2kdgbdO5G7S+udjW5Wl8IqEE
1pe2uZTOyM9otzrIjKlK0b0A8VyIuWzgmeVn82Qv+c/JnIKzTUeyJtpjK2v/6Z0wQMmMjA23o9jV
ACMZejgY/7clkhQ+8glTg8LmmP6W8pHvPJDBrUxkhJR5ad1LFi3xuVh3BueVZs7zT8joRgE0l76z
usN6vEhGzl65ovu11s02j7aGJ8nQvDJCXzK1gGD83reN9/Nq5pjj0f1fuv7sWPm56Bo0TUccACbo
TspI2lIVhyZbaA7KADuT2biVNKKgz3virvWqj0yq+GMhMdhJGD9pNeFq5FyIGHXDTcfKJ3Lcy1I+
V5znGHgJxEkxlbw9qLqaibchS631V5vPpKDASJRTM4hXGnHZ/UTr3F4lLvlUG1vE74yqE3gPAAlm
yy30BwL0tKNzIydeGgfDxk7lziCaZbpcHLyzHeL/wrxRhTEC7+pe7lfiXakCroBn4kXa2g4YBpbp
VpyqhN7FHvdNkTkxbx2bSx1ZgKWYIsCkN3Irbh/O304K/LIJ6e2gBTm5O4Z+6qc53wpprYLziZ5H
9O5o+z3i2GhSxUkRkN+Lt+VZAaaL7PAIoUiCHXyDDNrggdvxWDzg4SBro/P1i+TH0iKYzrFJm8hi
UkVT6RMU+9vPkrqgeIYMYyccReO/SJ+10tvgqT87/kg1pkJfRPyWf5fMi6pD+ucBYY16qKuC4Za0
MABc3Jh0nooipDKxg8xZJzWPy/QNI4sItHvAitmagZG9lvDwptQHvtF+bP/mBRzlQpyITyopXX+s
NvrytxrArhYzLH+u9JqXQ+sxpv/ljPF/gm/xGIVGoGyMYZpSjFHmiCNQle4t3IJJrMjJ7uCAlri0
/ipDRRQBdngjXgtORk6IjlxKAYiTpbKqfz5J4jZaJcxf15JRQcl7E4f2gdBYBW6/CxEoW3T05Uxw
N7ki3M+ac34k9PSdLWFj1T2LbWOrGve4zzpvChhMfiFhFOwu2R+Kb7lFK+x7oUmnP+PQaxCXM4hk
cNU8c9cKIKCERihjcuQPptxyAbnG9Ccw0TCMbQcELWfXNKcCT2UuhJpVyAP8RPWr2oXpEQ3mkROZ
TYTdv4WdLKHbEjwnTtpj0NL2vUpQgtNWZNuqNGX3Pl2wMwGOCvx97TSfVzeTZNixID8hN9nb/6Yz
wr3GSsUQdAXpKOW36Mvtsnm8jyKPsb1lElkJ7YIOyuhgQsXyXPsZHaKdQbmWq8F2RCy/pkaKM3js
C1QLILJlT2dx1tYGjmZ1IZT2bv7I0NprQq2we1y6qLZIoao9kWaEptRj1fhY3DSiMAgZQ1hPdNO2
9tvF7kB3MfPehF51/DMiQAY4IfPdOkniV3nXyErITBNQlF6Qn+ipNTZtByg5J7BUXqij37x3sk3t
zxgJLss2B5owoDOFmu9twhtLE7D/mid1VvqpVLMkifwVJ0RaaXgD6ZeoYei69SQtp6HgpXhwUaQM
P3as7FGwplarShMOzu+qogk4r4pljYXwSJ0QbQLwDjiUwdPCA39/Or6ZJnE1EUVXyQURkUwvRW9l
GstRSvfL8D9JuVmzlSdRKQ2DrS5KkA81mWbolsRTP+qUDAm3c+KoYGdUdwM5ZxNyY5hOat2e801B
hE661jaFxJOr0fnFVzq/Qp5RyJuJyklt+8jAugSriIqHUPMxD1lbfk1rRMcK9vddFfZTMFedL54L
DdkGpyre74uTO11n8NdfK1FXE4SgxUTrkSrQLrxuP9GMVz26DlLm46XFkm/WCctR6pGywl6yvxTg
b8KQz5xFscwpMesTc4TfJha9OFw5m7uN0kXxYK5uZ+A2Bak84vlinBu+owL0OvPYyaRWmFhWYrpT
v5rGJMifwehbwE0zJFVt1b06w6gbBfs7z8wF/Yy5rfS+J+gO4XNYxW34zn83mRxppFDbfxV6JL/r
RV0M6zNqt3cmiF/zKGqNeJUvpSESf5gwNlfKrrTcB5udYcjvD+G3Pzq+kdXJVeCErwn9+3Aw8gAu
t4A56Y/HEkFVT8Nv52MensACgjS5vu3FtVmtk+B4oto+UljD3K9hiShPuEoIS+T6Jan0EtLct3qf
HnqxFpV+Ei85GelhuGmtLd7Ag+KErEsKwf0/0ueMfMQHGbPmDqxpog4LLr5+ANEuCbKY2a4UNMCY
azWyzEoWPyFH3mH4/tkgSmIMtk3HUg5CP2fpr6nURvbbA9n96a7rm+K6PmgKJWgpkF/wvypBTg92
68gAhQ1XZRsmw1xzensEUxA2yLErXHeZLU2oGMORYkNntO45it2tvmU7KNHHPGRMrTcHB6HKCbgk
meEDkI+iNJW3GO1pAp6lvVQHle+lASQlef9ZiSUhSKmU6aH8xxtr1Aeu3Gm0gdKj/pEDZxP7TNjr
z20qj/lcEUs8gsXEiZ1RLzC+pfbQuRyXnvlpnYkA7BPPSd5Urh/FMg0vHMceNFBkxdSYXncEmrSS
iHaTjqroIEbZKf4B2aqh1xQBoqyfnYdDiXlIDTnwy5S3QP0EZ4HtQ1I+QQ/JHAJ5/mt3GyW+XdNj
uzfKBCU5LPETokpXBEdqvLkds9y1tOQXW1oNXmeKFtddmiuWMOyMSh09755Pph1eN3EJ3KjQ3Dji
cwFoxZGSBa52Hd77jStmhBq82D6Spzi/EsLBrLNG3SLqCAY9yYid5+UkYFs9C3eAXvqQj/APb1n6
lpPnGxkkMj+Zy6Ok4VUgeFC4/sz7CZzTMWL3OqWRt4sHOVTQVN3Fcsd1bohKyHEVKa0XCasx21Ew
VD/ynSct7oMsk5Ym8ElzZSyT6+11c76a7ukPF/ix1eVSJjV5ZglsCumTt42oid1wc+paqLiLXCnr
VCItANmvtvbxNLhqJX8UX6vMj4WlvJgTLL1Pf/HT6/DBkiXWLFIzBHqYX95Y6Gmd0zBZ23dpOeUN
HTcoftg60AAkqF2080rIn4a29TQuVmD+20lExxFOYHdOQZyuOW7T4YEpwMCoxzAVeRieF1RodY09
x5zXEdiksfu6WTFmHwpzUt9b+MkbvJnn+u/6VgYXKLn4+Kp/FOi56nIrMjS4vlADAWpDFYUtHUqN
VdkBv+h4YhjDnwzzTc7tA87bZV5fgFpQY2PoeLpEI2CqlaV3Bp0Bd1FOui9SFxjWfrjn5M2VLbUc
FZy4dKwk9BeclIrOuDoiUdi8g5j7AHan0y6K9iilwJ0+XWssLCY2H4Fl4tj4Nl9GnrkfGjnWoG62
IgoVyTsYyd/HhV3H++CTQaBIVMIR3i0WRd2HJVg4lxyyrZh4jIvk9GuLdonlwqsvDJkh1MANFbdB
DJkwE2Jp0F/GskC3okXfgqMqKnOsa2ZzJIVpCzQ+2U/jGZfeZzSqHlQMGbrzTWyk9ccxuSZlfWgz
bnj0cEX61q/+/bQuw39JAYnclhxvXzUjHPQPVURAE9ZRL0sCk4Dk7HpRLvDtH3Q1WsCVDTYk19Gx
0xmN19imb928TtYDvm41olCvxM+tV6+KoJfZpHiY1cypeFRfT2ngIOV1Ou5dkaVQJ3uhy91UM2mb
81DytDiCpDa3P0AksxPcXxEETs1nXyD4bANFmtdCTHBfhAzoHeG9Oh9kMCsUJ3l3kz3Mnu0+7mi0
LbEm04XWZ1zLsPfE8gzx+qmIOcHlHqDumsZ9JHDP0Xehexx3FAe5piFadBWkI4QHp77ggDTw+hmD
j7MLQ8KA5grSQ52Fn+RQ5Vd0GQedTFQn0njth7PnIMoNk/PjDbWc7mOFBzABR9RuzHuoUoL6kRLe
8qkG+OzhtfNdYayf7krbrQHoTSPzN1AVM0qxi0i5vl4/Hv/JV+7wtq7sTbJuPJs1+W0KCXgKJvTl
xoVIwPKJBw1LwuDkaYiyS2xRPwlaek5lr2xBgwq7VfxEnG9ySduYpNYbFwKLjMCjygyIETZtgMev
Eh0UOJ3R5nd6X4LjefXUy/EutTS8ospvC+xTTAgba3wg/yApPKHH5ZZrt8xt8ENbH54MamNDm63b
vYW2LqeE4U9Vz+n4i3wPgdoufFsquM00FrTOg4rHk+ruZLGKgei80c+SXM7uyXo9Kv20RULKrtyy
vmsvdN9fZK1ispRRMv4453ksqqDgyx9aVha5FQCaAw3czrwpVbbZnIkCI7tHztG1QcTFAfGtXaG9
jrSu3jZsxfhi5mhOq9EibWHD2pgyT/2K4ZKg3cKQMjil04a8Zzt+ELW8ORM9vCQHsP59nDhGnTgp
u7kaTNSsU5OCtCquicZBDznj9yzQQxNKEWUrhF75EG72KqVYrCACdvZGbsoLRIk39LQxImeUeJsJ
VdCmSkL1hZW4c+UPDgH9TQ7rRAGVFuKrW1Q7aI4Z28u027pTxX699v0hfDZrCxgRbI14uwkjyt3T
RmMa4ugDllP6BEmTn8gfO9w+UcxIVrkXF7kdsfqMjZVM+wrz4x6+r3S94R8J8sk4nS+syrf0N2Lw
4kkuZFimSFrtNehd3GflvhFgBtg3+HrefKIMyIH1Xe9hHUL8Ouf9buFVikfmxsSxyWVH44JJ7YPZ
QbZJTRn0OWQydG/sWsydOXTTmkUF2htQsYjx16FjSGGosxV0VzorwDpNR35fFI1JB+VxtR52/32q
qOYEZpbmItLNe6kXrFFmHpJi+8hYO+aVfEpbY2tMDE/gaUN2+IkwXkyvkHwONsWd8R75K/fPAULS
hdw5xtIyWKteURr53vG8dZtvrfyUOE6GLVcqsY4fhtVJNaQ/J/9xQvkMGNQN/fS2LOEQz/3W2A/h
qVnU/KtIgiYOPebobQ9FMBp/lrgNJzGQZxdbOj9iTc3xFm6z2NQtRvIKFc6wnS4sUNQyNbZpVEKJ
YT/4RZmfAQCx2EIp1yLI3GmfDxXcPiElFsuwmlAZWCF/e08FV9BKrGyPe0IlcpHpiZQVQI19la38
ub7nHNX88HG/yFce8P1HGNPknRalV+GKBTiZfCAKNqwAOYbkz/SBL8g+/QojD+yVh06mUbHM8DSh
4cYD5p2GR5LQyh7cHDNQ4ZPOl8AJKUHc4ch+faA+N9GgxOm74Vqbl5kgJ1RMGc+ukGNOyWe9/cRl
iWIddXQ8nuIbCq3DwmcIVZBQcBVfnMxtnOLHAnVUKy33z9MoxaGQp1N63g+rcyGmr3Vs5cCh6nad
RLRN4aEtfkp9v32wOHCjkrSuB1tRfIkm8VSduH2XM0uJ8PkS4jiNwiaBN1Ompzox52U6aHb6CTAJ
O2WWuI8tPrbukdWzF+DiExGLL6B5oFcPTRYihFyxXB8CkRiQJhpIHuQuVBQT8maPpDU/MuzNYdZB
+atlfuTG1ekgl8e5hrZRXbBZKDvphXICpdW315Qq+oYTul+Bl7XCWWs7mtg4kc8zksho5vwYftsB
7Rr0RQv39Mc0bmYb16bhaLXICZyz6AzY01enrYKSWbPcx2zXzADMMigjMlGFwyFZXxd1xDNTc2Vl
+QogJaUpCmLUpX+LWQlv8qXPvgRhTCc5/IJkyA/wLai7iwxtaczFsvKHEHyWUW70HTVaS/bHNSHm
a2xPdeK/X2aSdTUjLGBv/M5c+xSuWRcWg+uq9975M4yPfh93fAkw5i3EBFNg3Ag4jIz1Y4yPFfas
c2LuTHZWQ59SkPb0f9Kxk6ZpLENH1EHFzedQtojwpW1rA9pVOn38jymJyx2JAhUT2YOsfajDlTnQ
1hZueUYAk2rzHGiKmmBulIdaxU8x+jSumLUsReDqqvfNQ25US/mrK3KOfZyOeHmtNImzd1gqzdat
+NVf2t39bR2uMrA3UDtzTgLXDutgln0v3/KKXVtigpZjOsE7LTYEucPXzNvwCc4GByyPVwa13yDP
JcBcWEPYdgmHF9sAGajFubhKxkqPe0F9Ph6kOGfy9xsAR0M+23PfqUewQfsbks1TbI+3ZmVwNVlP
XsNlkqhK7tBMhPvW8dSTdd2xxCtmo0FDFV4MhLDxrakybyBYEpRj6AqUBiHmBWrEP6BJCUNLcfac
wH6VCc4jghCCJ7ZNyDAqQnWUEuVVqcw8+dmqAIHPFkpvcJuhgPpGCHN9Vg1xDN838+KZDtRtrdwN
qXEj6J5XWBnlI1tTVZskIlACI2JgGO+kt9VzydCIKebvCLVOyuE9032Tw1RwefSrwZFlhqP4diWf
Crj2C7K/CXkqW0tMHvnMsBRTA+mTCxfkh1LijtjM70y3FJZiebCGF+znST/UOvoNG5qHtf71etqk
7mt/rhOCjt3jB2EZMHImCEne62uyVYDWMlcVjapKJjm0PYfidLIEvAoXtEQw+vXuI2+aFBWf3Iwf
d3wq0O/SnzYnlDHSNzmv2OcaaLQn3aEx4k94804nHCk7S6J/1dzqJo5HKyF+SPQwQNOjTU+pHQPN
BZLes9YQntwISsTOv5sMjCG/69emL8j5s6GuDq5TuIAewnSJOSxJKu8d5J0kUkDETfTuBk85GENT
gROFOZv6s4X2RIpl+GckkcC0qCtq8hOaCBnAov+kp5Ff+8NxKBIbSL9L7kM3HEXhvcXatI5tTXNu
ZwJPuBaKoT7qjrnmRETF5eAL/WDbbsoP+Bump0vdhDwsj1IgBEOSRv8cODdUYUxGLhZDk8TWOx8A
g++v8SdVZ00kItSZezAY4mRs7GlhfQSX75lZcD71kaNyWPLU9JwjUlLdWj5eaCw12LKn1uDmmun/
NAYIysn+wGonX/xM3oDW2mCmg5qLgSXqY7wMGBHEd7R9s2XyhcMkrgClVabgX5AXWRmUY4FXBLaj
Kt7SWFETzJ1Nchy5gPOhXIfzwR9PM6cxsQoUODFi3nfpC9YOUaCsIcOB69mnetKb1SyfRUBhlmoc
ag9BufZ+RZRT8gFcMsKWShfaqD7UHz3n7LAmYVdoSzHfvD0uHxf66fqsRyHP5kEJ0XxkzZ1elvTs
JrIH543QrznZjhuPtKIoG4C9b3/Fv6QvneYds0L/J9D3eFM4oJmsvvQN8HSWxjSlS/+xCG95la3a
n7JuDTYw1Q9bqS0sBFMm8jJ3XvmAST834H/dyCLTAQowGL7WNeEMrzZpCdBEueauYk5x3vdNGy9c
GGqOQwkkoRawlK8lNGkFUg/7c65O5HalhPY0zOLQ+jsOJDkDhHMPVjm4BaJSBsJ0hsw4QrO2SCG+
5QQC3Ew+YJJNsMceK5mq6xBGvhEGlo30dr3cU1BQKlHKZTFbQ/wQaGj4+urpBrVTYtfOj5C0vj+E
0fBSrWDkJhUvY1f8naJmUVHQJtVJ+B7qWJp5KcUBuJkNa9p3coRRa+WpwF00YQbseKH6LgRk9+n1
zXSv4FbXevA/eKkGa8YGxdesPGvpR/nWiAU9rXDskpovKQqqpeOAMKQhkKX8Pvcr+vGc4i5Ibqtd
5CSlCTzv8/kLN40QyGY0G174JynhbnxyreywPzac/Cquswt+mXVLr/+P+FpCwgoyA8BKEqJ24vjB
m9PilU8dQiC+T1k/8puTTuh7gC1QH921Vz9eXwGNrAmrK+iDK+To23kUWvEj9CPZfrMhklBrdoRs
MKLu2AzPaSOZux3tG9AKR/O9ZLSb80V5v4VQXh977GJUxgEtoqDuz13PLhl5O/6++cjwDS7N5xia
L4zTDxSe7yOHAmW1bt/Z0V5lzF2g7DYfCfbtmLv8nvk6lZheYhRE5qSVzM1VsKhY8LU0myhn28eA
9Ompm1mcgeP5OSg2GLuTAPhk/7e+LTR6osPeTFYw1L7I7JOk4pXGWnu3qAQsAu2qvO5EzD6VrBET
rj4k4SRe9LI7OU0ljx/TK8ovYwL8eoyt0fgixlP0PBGFwSe2UpgzGOTohkBds1YjsJLkjZYbZK0S
b6vOBGeafH4PWGGhh4te7ZPlPhnE8xHMrIXoYxjkNTD94nQiKpTFyzuBfVLQ/odQBEXku5m2o8we
r2ffvf/Zj0SuDtsW2ZS4cqlSEps0eZLkOZ4mfGCQFT0KWjPWe6tXJoZOCDrqWSZzNZPx83jZyAiU
njIQGoHC16+3pe6QEv5pCI/OULdhiFakC6V43iE2EiPr5Y3YauWhs3WqCZ1sySy5k5K54aaPD/T9
jWThsvaD61wNxhBj7rz3O6mqw1BOOXb1M550ZhudIy2VIpuJCnCeW/V2yf6PvgruAHK6ZVJeFglT
PRCHFpC5CJKXtkJtC53izFzApUt7Yq5a/Ff1+c7UzkmxvXWKwFT7tgwse7/mkqk0oRAmAq1m/rf+
Ei9fHhxAVVIEp3B5bylWGRhkrzZfi9o494hWX+dhijrkJvXoffqiQ5ZA+234nlcHZqLE9QkAHDqC
nGdeCflXklgXZrKhbv5c5IznxxLCxU7dtb8nzyiUhNc57WwzziluxJHGIdtF9fPsX60CLxURITT1
IOI4/31uzTwV53KnO/BLCqyEiGTO58n9O+nvQvJ5F+ZwKnqDOze8jC6OpbScIUhuAJ9BeKG62+HN
Vsm0LbwlETOXyPyox85v7LzbOKDVR+Xbgyn92iChP+c3nkxqhUOBsukrG2FrptQOYuZ8kp19QV7P
W0JI40w9yu2mvRO8AuIrM7ZJA0+c5nr0VVG5KBK8SMSlolAk1S90GzN4hIl/lrLSbYWv67rwveLR
Z1ZjraMg5FjWyfPLXZVqSsx255m0cIbgqMkCxaGAclGs4sWxGwO3Bj32zwUxK/oTUottclu5jYe8
84D9dVH5n39t7kJVZinl05RWF7DJDCKQ2zNfE40xpWJY8g34kga5WcRVOT3hGBvC3KwDICZMq4am
5nYYeuPBb0f7httuEWx2nNJF80pEC/wutN8mgluygWNhN0Tf3k5qNXjrchpnp5P4ZorKqsfxhzdR
1U2bIk5y5N69FWkuNbiVQ+rjOrraVJQzeEgyZuporC6d0PL/h8Z0gfiPnCHQo0aZujZvHEYCtLQm
OLM1vza5/g7Nksx+NLFlw16Cgwf7njpKeebfShHHwBz/A5fL8fztePfjMr6HDyfqSD8R+dsXD5vg
dSuDOwAjpAtqCUAFTsObPQNUMsRap23dYgk+YyEPSmSiOt9IoXdF32zBDqeIlC8aolV83QfBxjE3
eM8YfnPnWpCkmkEXb/b+1bPIeG5J3UpyBT4u4YSR6YLUhdTkflQqENTxVtvhnAxTPu3iEsjHzPmt
ciLMyALvWDOG6BV7zD5yFRJCm3GL4QD+ve79pP7TjOaXaSixbbY3J5zJckNRgYN7tmRr3jtzaQjo
849K8lIGr1NFpod1CVmgQhclYRm+BzmWlK+hxzgeDa7cGm32LOuuMW5E7ZD4r/7SCNEgeuuUYzt8
8sD/6EyTn7TZZMIFgDScOopuOT5inPAkZMuG6VrrcsVLBant5STXKUvofL8FZ4g8/8tYbyEXnXM2
ghtRqqmISDofv3OV6nKMa0LQFe8qXl0UhrIyTbmp/kc5iGayw5pWOXt5jnm9sBu2aJ7Zdto5zqpE
gQ7JDAAUXo/z6IR6eJ6IwbhKtgFDZzgSrLfB9TUmDfI46aMXQ97R38TkWu2EoaKS56M007BpNINL
GdzoSWP3o+mX+7tlEWBkRLtdyJNNgTGGk1lk0t8fokruP14IKs6VyjGGVJQcEdABSKyvZoxF6ziX
XNg4gJW6VUan/K7YoIu+7zzJeJ59CwPq32t/lyHALZaVDID1XwIaQ5Fp1P/fpel/q+NKD0CrvEQX
xWXIHQ8HUMzfjC55Anv4VQGN14UxVVfmxhCTkxZlbao+qmEiS4GyKONs3tARmizDs0p/uvP6n2gM
0SZewwpOCC5k2kX9DllAzYq6r4FE09lDBLuCYSHFxMGjpt5zmpcKM+PFMjAbwIXYl2sOVKZyCpYQ
Vij7ELXsdQJaPyWv0oElib+/zBAN8K5o+RI0P4TyYfGk3dJ5e+wgH05FBPY+l+g19QyjVPUwYpwe
33YKDW519RPfX+uh5F6x2TaTzyF6V43gKFOUsnHBYH1KWgEGZ+g0kWufggBLotPt023kwAFpXA9g
4xdeSsYKoCw4TCgbDdNAXwgobWGHY7YkoOfpdXwdtSbdUAye4Vd2jbK+N6ODy9IezfBmxAkQfToh
myJ7MdLCoKKGz/Ml5KYIQm/XQrwZoxxUrT2yO2FtZm1rUdH2XcCnUue5TxQ0+O2I+H5OpsEMZ4b+
DFqO9T4YoBuOi4pPNFwYe6rOJi2CM40Dvtpwu1CKKT7Tnzu1qYE+7n3llRCSRQvSKgi9OUvH8DU0
NyvJsyvIpCwyhBDcEy9bWghDMQPtNNMoNfXry5qWhDVqs+HAljPUSrmViJoPSfOSv3Q0E5igIiWp
x1kIrlc1xq4N8BqQCS4xrZD7Ds/nInPgqqRG2JTKPGE/ibxniUtDbwByRiYIfuoUiPNpt/LNj1Ps
GFy155Wlx3w9p4N0MmXs7x6pOZq6FTVXzuD92s+IpR6nbEPWW6niPxhcESzZFbcEkFqfxXtoDUps
RYSuQakjTzAUY5niKSh+tTotofDqTZMHttIb8xMsfVvfsxQ3duE9xoy7HzynOgYJF26ATGFVOAtH
ejR0gqaWzds2PPcLZml32M4zL0aRCZROvBVbnyiYJmRhwhzMLLp7VsQSe1iYRHb8pqqY8zNhGvto
M4+0iWFhfFN/CLFIE5A0oiRevg2doh28dyepg2/SULrdwEVWGcrpUN7uXAf4wb8ZenAE3/sR5npE
uadioo3fvGfzk5VRrmf0Xmg3ZvFMjRCuPiDoNf3yW2Kfjx5GRhkSDpA3/P7t6uzLKCXr2L9DFI/z
Ok5dW6dghDsgVMJWWhfY7SCZxul6qZwuO00sAOkTPsX/JSgAJ3F41rlUwpmpDhwIoa0OXYSK/HxU
bOJ6dU9jkXDm/W5PTV7r+OYJIuBTa8/h00BZzkFYr4Tu2rhTX/lHc5GSZRZ882O7F4onyoHIEWNg
Sc4htFNmoPjq1+gpvLQ+afZuSt2LvCgFFVPvFUAbHH6KPVjSpR5ZViD+djAJCJyq237VJ4Pp43VO
aL3a3DaZ/4lsvxeiAaY2qFMhQmF3o7ihtgbpBJlNej24ZSJbvN24rSw32y2n7yhde5stT1LbEu/W
uAcG2/CmtyLqb1giv/3o/0KTsg1WhQvqyQJNWP22k28f23/ZfKHSqi+Hk2dHURMinAOKQ6+MbGWK
SkTZyZXE7PHSKPsR1yGhIBwP8zzYZb1vB2vnZRrGbmpC/0AtW20JVR7Zll2Hy8qeCWq0OH4Yq5Su
pvqfefSAH8NXwJWWbzyHLb5AYtRvm/lgViD5kxdSX9lfcVhiISIZBaqQBJYGz5Oup07ooDQQjKip
JRl3Aolg9PPsV5qjpGICGhDqA0qfaravZ8PgZiiGlmBFk9BwKyXGO4xZh7uSsiw1MMB4vD8qTP7I
xw1QJDqaNc0ufMoO6MCPYB2yfVjEQO5Fmz0mAgY/r13XY8/szO8LMfgnQp7cyAl/rfgW0KU1RWMe
eqT5qCF778k6+0YaqkDTjEwe6viHgmOEolVGWAQgHlfShS3F70kAOReBVIx+f7TlTtRJJz33YIdp
3T5H6WSURDlr25rrByOgiWDPNu1GBCzOMV6mwT6IXIalDVRHwF0DenpNUaaZhSzDky4KZdsRkVFB
DLLX9n0ccUhBwRPEBzPeyFMJMx7zDPQfz6jz5cv67ESAHYZ+bNi3xXpbwJOnkXCuXiu2BnSkmdNJ
eo5NshMNx+UQ6Ih/CW7I2PeCChrL4qa9nO4HuCyfMP937UwQ3Y7cEPytW+DD2amXlaNFR52yEgZ/
l4TEGf137/OJPmOF/iHYW3qucNgps7adliXUvly7skDfKClh9BeWzJbra4ULzjfyaRrF5iyHFuL/
NII3o69VWrq0F6S2K73jQFntc7a2Uo7cZihq8y2i1LCpkm1Tc5HGHtBD6YnQFDf1p+bZ4VSCx0YN
QIewJi3KCBxV56tSoOxr5AYZUc8uVpjm+Djt448mV0Wm43J285i7rf5uuaTIIJuv9xzA2rze8qzb
ZV/6g0LIkQ+LD7cVM12fLpgQ+PDVrRS2muaWsxtviVHuvdI21yY2OG7n+uMLmOzeeAV1LpnE8jIf
YSQeZi9lz79uzMO5FZLYo3tpjsCxxZirkQErzI1wrBR+6h1OXmOkHB6U/aqOGv/2jXKf2wDthvB/
7FWv4FasKVvm+Jo4/Sk2zjYfMFhU0vEIBuA9e8d0CEQu0QXjdZLUwXUnVpSYesh8wCdMRA0x3UjA
hXukxcq7QHmgiL/DG1wjmmniXpXw/K86nbyORjY1tzUKrqVstx4Em8PNt11uTWdcdYeBKsKsS5me
vwq6VjUAb24SP/wQY6cQLmrxcETlZsG7bvw/ndW/461Wt/wNXci5xgdtxy7QJa+kNsh5+Nd5SFBv
ANtOZoIxLtyXhtl1yBV7BRvCerQa3jU8+F9Q5bpNDl/5+9L8x9AyWy6+nPJuYRt+gFmwPBs4MTw8
bdiT0ADGl45GYysiw9Ku7P46iGfrmNpo6Cjr4qgKkXYYBjg//2PlnUJkOCVIOmeN4f+6D+QlIUAh
D76nY1+IsYT0ByNzy8iJ2AAi1cX7ZxgHE8Nk9LXqTfStwTWA4s3EC7rQG4XZDZ0RpwOIY+on59Hy
ttpy8fc6A2+gCN74DCTi0qWr3Jvo9dkQRbEkWBGAE7aV2MMd3Kc9+00Ns+gtE7SUFRn7IzI7SsFr
Qeh9AtK6wUJt6RRSEgFvuJnXE12zG7RjJZNIS8wZgXRHmTEcjaa4jy8oj/HTGZ3kw2NRuhdyztEj
JjVL1OrTUFTvOy0Ws+kPuVF0AVkmtFWx9PEPWYvoWaTZs1S97+kBkCWSepA50Enw/nyVsQUvR+Im
+8atvLuZhpkCIj1B6V8a+ijmZpwD3uDBmeGyYxOuMNOdvLL+3BQXFnUqUCOXeHZIZkXA0/VdmVek
26/Sv63xALazd00foeysB+YrQzdsuMcRow2QjRhkchsOigLJ5pgDcpjZ9zZ3IQiJ+pRTzzp88GsJ
bPyIgjfWVafjOUiid9Ip0ThhrbXrJZXHBJGzK5s/VKHqaWL1VFgl96Uc7prkM8RE8/3bqCsaNi4K
D1pbkLhPIMgO0CtioNtkcWeGAqYusXZsvG26NefPk3IqVMuexujABmCRNawG60WgwpiDOWAZRLeT
+owR5XmPtPeQvYJhKAeM2sTC95SwAHn7zLKrizDXa2x2zVs4hZb9yF2unkwfyUthGba60kOimbl+
/rRjpkzbt3jfZFzmAoUbX3sCwGsHhqVVZkv0mnywb7xyxZ13tT1KyvYG1KHYhVj1qggD7Tc4hzXb
q2QNBp9tbYdPYEf1/Ek20bDhCFjpnxC8Pzh5wBI4/vJseQik+5BtnELIYK9034T86H7WpoMHeQnn
Tv2kkHPjvLfprATUDaRZoP+WmMmZZul8cRv5MyXdjPSkA/vBH/99bMVvGcxYspGdiM1rkKFn+u4I
1ATPEXcMaTKtB4rBY2wd+N6oiNBQpxSs2Md5WL3MlkxokWVDS7a3mMe/xPsyZvzd5ieAa0us9wMR
hvA+cCkvL6mXKrEhKTu6ciswfUz0Y2F70UluOoG1Z+zhEfot0nBhPg/0/k8yA6REMysp4G4GMre/
fxSSQ0CqPQUcL1ye/Fa+Iq3X7ske4bGSH7INmLkjgJkaUcvv3E4WltljBpA7BsZHPKNb1S6FC7Ew
jIt+jq/LkR/DWwl5WEEv2rppD5ZvcRS/gbCtvrouGOq1vMGVDD2oAzgZE762/iNThBnIS1yyV+xh
/6qEAOAaguwQYa2PWdqgQsCLVHDNfkoxRGyMqZfzq0EOxiyADRWE1mRtOk3MDCqI57wJa/LCDa/3
t9FjlPduAXx6AAW/wxYxM6cNIEq9Bdwkb2obdT0YoKg8pGIkby1FVaEmPMTf/RlKRnWmcrqlqqk2
CIXILHSpKdVj/LhY0zmj0s9BF6NmW0SWsAuMEczXxfLllSlNB9wgQp4nQDilrUqfzUZorxtch0Ti
papYmj2EMLwm5jBGRMSCTNc1g9a4u2J+OS/gyNFw3hA7No62MKymIrn+NlJ3LEdUPPhg7oEyUhoa
9Iel6rR4mOPpGI2fHlUBGraDfRRjxU+aWthWxlTsSsH/yY9Y4f/o3roIlghBoVger9NLbovgitNZ
tcgRVaLEKTy32Q3+ss/jLTle0Fq8vNUzoPv/qLWogQLLBgQ6epAWTjfESL0cG3lREYmsGWIimK4k
mJ+CocO3yvAQudanEA4gjs+5ljkFcJReHQl+dQvN00TYtTc/DtTfI4vEAd/4FY4yhQhI4EZ8cui+
58xSaNzqlhfc30kyDxyXjeu5TPLzGevTPZZ9U5A1Iv30b0qzekH2Xd8/NIiSEg0vDObhJ/2VN33z
1gRZ//JvEfWhpTbmCtmfvfHQAsV2IwZ+EK+AHU7CejW+vbr9fuiWiHThfnRkbWUk9BzB2kzAyitK
oxIMx5gRRRkNeX2+EqhC0w0BvUmtv/1rSpiFrk3atzAwPp27drl1EW4fyUyK7bnDwOD27JzYPDBC
eD4eNaugUPiO8nrTF7LVCfaXndPRHLYvdupUqWFcJiTVbot2dcMWEbrpVvADoZbXieA7zDwQD05d
oIvS0EcY4eSNxOPPe16JrA4TjWipXzW/wG0t1iQW7jhKSKUeFMIQ+uzJpyjmJZQFhCDZyYnm7Fva
X2+8y00LTrau2rFh1i3ZPce4DU7PkOoWBJ7HIwtsv/N+UfGbxa3KKw1xnuL0Dz0OjFhJhtFPisew
iA0/deGhW1LuGPJD+6yGq/O6TUIK03sPH93hceJIxvX+IdBrytVHlwFexE+Eat5RHNIsKiqCQ4Jw
Z0bpZaoE4JW3NiBUe/xdFLALoRfavLoDuZeffrOXTCuvp9KYg6SBFSEl9SDSvRV6Tmh3jetmahyX
BZw1zlg4LQZt3Dim/GpGzYLR4EJXLC4VIbyuTO953NiftyYV2QvB0LCplcC/6pHg9eObZ54P2WYe
P8TCq5A9hVSFGdoVyp3muuIMAk3qQBlF2RaBzaMmigVTKEeI3asILOLCKbNawgRhkJCuQXCz/qqC
s/Cz8kgVXPaGFsPIw3Jy3bi2DyE+OcErkTLUxcSiobGe5fwSlXWKE3eiDemNTdn/X/pVGoD6zO6D
Gd4fIAMGbc0M/y16hpAexXHg88w2mDOUW5f6/oDecepnAXLlF4R0GZiCunenEwjw4n7GYEBBiK2x
C+28SS0yXOOWC/SZQdv7Kjjox7p/whKVssABikXf5VEps9/09aTasIg0XKkWT8LLWbokG1x+IaVp
Ylbt0EN6iQBrYbq1yzhhhDZMbSM4eiZtx7IvRq99rryknCZMxTs38hwS2Bs2GFX2x/B57ca9YhTR
Dv0RZexAfQ9pqR4+i1orzXREBTwUmiHYa726mju5bUuLhv6WG08Cc4bb+WDkSYUJFKWPRzHTPYI9
QLaHmp9d0vgfLJ3659NDL9UY2H/OsmhCH8PdOvINezfKpnX4iXUFIM35EBJZOnauX7HVvOUICTcQ
Bdu8x6LGG0AmITXO7GvlRueP0gBSS6W+N5BnQP6Ovnjp5ZgErQ0PfaWWj/jL5/ETy1VwXUvB8btm
cujo9bRUZrLKS44r1DtoQjWzf5XfO491x3r7j5w45xkQhXJt4+3LYbNI83Gt/H02KywVFetYHemJ
F1pyOl7wy2t/BVf3qtBNnl97ytXqnXI3ARXRhd7QIg/sP//UZh21wxARnh5hGzh/mN2L+0RVJnI7
xQg7senk4WUQ+B43zC4FgbmP55yJt4Yl66Zjt3H29toyx8rSO7j8ejPOAWJgcM3/iFuwP3IjylsR
+tiY6OzIeZHVlwMSPHXekJ1DMC451tnZXRKgB0dcHg9dfiaRRnwre/FCFr3iV4mK46G9yLrhQQqE
aotdTmM0sZFBN4EiZF2kSfOltg6P/2xY7KsKfAvbaY4ivfeWtZgtQz+bOBOEZLY9Ag9K6GllL/eo
9xSpPgYGTN2R7MTanXHyXnohg0WSf74pRxjTNsIWrrazFJxOyzRZJmOkRemMU60+mDT3nelntYfN
/hm1IaKuYzYMIg59p+qFFtLv7PcIa6rz66L3vSpDhRKIvgZqVMcSZKeykMfatYkC4Ex1FQfTddto
crj0c0bl6+afmeBgDRY2eaaoAoQMnIjA7tqX08HUDO92uOqmkQWJrxVWSOS3Zb3CNBWWWSqs0t1t
p4k6taAx/q2dedLJlF+HQjUlqY91kA4J2QeByuxD7Lf4v4tMTrtHETnz8tJ1ClU1pkuWflmpPMWB
XpCdSdq3VwU/+nM3thntWV60vbrtDYdV6vVuUkCCWJKMNxxTWFgwBszFCCzD263rkXWxDJCv6wX0
oIDIRL+br9kIjEZ7EBN43NWP8VjIrSJTSXYnSceBhDVzxgXfbzegcpHi+ky4ap/1a9R5iZMFj8Do
j8wF6zbA1+JNiR0s1IJskS3LwYgLW1mhlLNwka6rLM/nnG//vDCsIDdyAcIH5ZCKp2OtW3EP/ZyX
oyTRxasRtQ8I3iV6gSur1CET+A0WQVKUiqJRBBmIbHZQHdXyOxwkpEuBWbY2UsQ3C6RkZ0ddTXQl
3H02B/eaUv4BPjG+extWDadi37Vi7CAcDl1Zv1srgohq05lgh5kcjDPyz4AiHXzov7oNZQ5xgbk5
iCKvkuRymNtAIr+rHRpIVRGEE7tgwTE6+tzWbBUVYMo4uMErQv8mZ+ZsQVG0EQM9enZKJ31aZKEC
5YAe98dygqZk4Qw+gDeG5Qra6KZaOSJgwrHfqPf3L9K8sTdgWCJ1eUrxWjhECw/lAQz4btLqeDhG
USIbvVkJQESmdqoN1SmRPUHhemWeVe049vFspaeQjElyBvFBXt+Uzzi31iFvfyQsXpE/kbCE2QhE
Dj97JJgSdg18wL38x0p8dPhZgcxjTPB2+Jp8p3HAjvvjchMbrDg8qkAAyiuXj5svOuH25igRo1Je
Loa6ruz8hVuZKeqcNFoyIzUpsE5l2QNmywMCxreh8GvygdrHvdN9Ni+U+2C8AbKBYXXpnX9oSKrP
1n5SAvgpuo/dde0YvRB3KALz8MS/Wl4AZwv+oKolMOmmADBiUe8hS85zvTY+N0nmw7vZF2DtO7kc
2T06FWRx1a3xzXe+5zwdja3QoEJxMCTpGxyYWB2TQuOWiaoFefSQKLQomI2ZX4Y86nZ0CbAIzUnA
GqcA55aRfYfLhNsZsqHn51O1lfDDZT/1EdxsRBgN7/KPq+5ibnQ3bSn9gNWArlm1qENIOBGgtq7W
kv1L9cemqPsNxzsUhgo63dLZQtAAt3CSLu8IjV/Mc7yn/Zfj7h3H18Ke/EbLSnOFi+/i3ppCIvb/
ANUiyoZHKdLX55JRAYVVN5pDK+PEJdDY7MtYG20A/ewhmEdhBXLgeet/fM+1/FSE7nGfXJZWC0q2
4hn+ufslAvPyegtjf4p+WRKb2tdQuicol5VTHSVNWRl9j74LMHSzusnnCPtSdg/0sLuTDCBjeL+d
XzXLz66lQHQe0mrJPqJcfdwH3IAdyYdtiNAtm20WBxXfci77/f9bCbTdGXqGcNNVIQHoifBgc3/Y
ud8SwzQHk/eUC8qyQkCqLrjNjbCISSjT2eAiFcTmvsvz67E401WC2zUiWXh6IAt6X2jhIZqJRc8d
2Ot1XdLhPBj/5tcK5kdiPa934xZOWSBGBGXOLlZTIAqLlNtLNRzKzVT0f1JPgu9mPtuzdcFPfCE7
hhiBtt0mOG5VWg0GmYfrI5wtL+amTtMUVScP8hAsSbnjNLBUg6WUk9xOawQR6RWiJwSBv+oa7uc4
SORdM6aF8+TLFLUKWfkvfbuHr0pup65kCrm5wNpgo1rVV7WsM9AhPyZZf4o65lJhZP9lwYLdFFog
wILV14UnHCJXQyEj1GVA2TQAuPU7k7qtDGq33yc3wNLp2sBJzQ0zB+HFxc01bHrXd01VMrSCetqX
1o9TraEpci7oBPJ3gNG9/3CCgdG9gOqcBEEiWh3wy+Enc+90cejVTtKPC958fHoN5XfCuUfrUkAM
HhFLzux7iZCnEgg27qmSJjFpLIGGY9UW1CL8TJvXXfFCZeaXvycH0Bk/sW2nQ2Am3kbpfGwh1xtH
zaFQe1aUJl4GSWoKAK62At/T+DhjZKsNiCm3hPxCg+vm79rHcr0QvsDyBfCFfvHLQeD5vVjOWFML
enhe2cvX3WhNLuHY6QbEAvWVCZ6eBRKbsrfIJnNtuPmhkJ0zFA7iQQVFUqEGyws/8WgqhGa9bTcP
7IYMq3BUuXH+C6dmOMA5+ofMgJ8zdGBbQLrGjSWbDCGXvoECn/Xv7/X8TCYqn3hi8shR4OnFlEZg
nO3y7ayu+eLsm0F+rYA83QLaghe6RgWL5Y+Uu8ufBDFogGwbX0ioqO59LUwKWnAlRJDgwQhrplfn
D6hYjZGOYD1huFDYsMogLUMQFnhWqUDpc9+TIHP2Uov3JfoLKjGVO1NL2RNs0ji0DgRdGI6hbBUT
EmRORzezbdriCmQZWSpNaVnpGFbujiJsVrzrJIRLpJvkq/JBBCfbCSh8lfqNNm4kV5jqm4AD4Vct
xa4c7o9S19RD27a5OQKvt1fwG0UjbpoQi9abbJAjy79SmVf7y4LEXWNRMkFdIKco2WaoG+9X4z20
9HkZsHLaqxeeKD7v0riJMbZGJoVoi93+LisszrOXT7PiwRYT28lcSYoWM65jKZWonOL1FSWNb/3q
+gIzoGUs+dahec91ztqYd2Vk9k5UZ9wc9S6KFmkjYp9py3I1f4Sx/2kB8REM+ddaCmwJjTgow4Mc
3jghAUbV4V1L73n2IjIXN+AyYen7jR11EKshyipyupBkOYVfMVi7CQDn5gpOozasAsoXEcerXkiL
a8JOfxp7MstD/0dU9UrCkTMF/rjAIanCoxlotmR71BRx64gTx0sGwWAWoJNwhLku99k1Db8+VJHx
Yr3h3d8sdh4Z/xFo8BuizWiZj9qlivHJEmkmcWetOONJu56VMN9nHStCmb3hX2mKCzrn/EWSVaXr
RGGTWXHmHrtOWQMZSU1C50Dx2josZnXOOKZAGnH+8Of+wthZ9FNnXYkgvAiFmjdIr6HPPAv8k0wi
pKlvYwA5qAiu3NiRCSFzyVJWrpGXJQKleOM9JTl/tU5eSW+4BX4i5l5vo2ZDTMFb94CF9Z/WchgZ
Gm0Jl0pXX+CNdBh+rgKEI324yfIDZE3/Qolz20VFesEtx8CkQzReUeJjef97UM696ohv4S1R4vwy
Gd8zpjovgftGrcMRcrb9TbW6N4OS1ftCA8g88K7cxMJSuZJh5ZNC48aJ5R4LOxAz25nZwb6My7nA
DNm/a0zJjYBU5m44WGkLI3++ZjxiuE40M4aoTHepOl9gfMZVkjM3w0bEvSOBJgucWRi8E0l+tALw
gr3G3ykgT49zJ0mwczxb+QZ5rT+2YXEb6YwUBZkyGkdbx96LyDR+X3c6NQJcdWpajDjUDYIsP7Lx
+tsDOT3bXDnBrKZ1Nh8DmbggccuPM1ivGuUYMnpGzMwRuEoURC6LMhKmScI0xmLMWYpyd7+HZw2q
JXWFtjdALprKiNXfSh+7XodGJWIJtpFGIT5wIzx3uod1MkO9kXHRBTmfWFhJUPG6ify2so6kEC9r
LZAk8rJ0E0vCvE5Mbq6qW8908Xxo28RMl2gmkrQzZRPQ+aBXxs9xX6y0nax4IVHSHMukXzlR0Ojd
6oLy2qOWWZFP4AYFEHrx9RZNEX0RITwUxVqcGOflmEROOIh+aeiIHRLMbVIsNKsjUwGNuCnaURVI
xooUeeP1K1WVWEyCvT4f7NOnFfWZs5Ee0FI3J02HB4gxh4XB0aQsDavvNHQINbg9so2YuQIc/BnS
ENirMAXaq7UJbfpSQBpeoCm7JdAavd4A6UBS3NFKUrZQR/Y7b1rtmD24EhrTrH00MjmdvT0qe1RA
QRtIUZGPPKgyE0ehndAGXx8XD5I2jZbpCDuoKsa+zzxAylQr0lO+c2SnVVSR7K3oX+h2ABgtJ5jG
oaFL0IS4pXId0bDlt8kyZr/10KtiR4UnBG6EyVcpskwGIVL7PUELTvwpGWEgQNs/P4doraHt4qTu
Ol1qqkdTugz+zQRPxRXDRNPP4iCUAgtpwyuWrsUtBc3RGwknP6JTDhu/a8sUPoSiK6yw4Ce8aGgU
80fIq1Q/UzzPOQIKY3AbGTt3/eU3tz/qzlyguEH1ju/hCe+L66p2zchM+Ce4ZpMm1N6yN9Kq1ZRM
o+xkCflnTjTL6BJGmb9jgAZgGOvLmSdo1zz+qmG3BmvWUD/j0wnwOSF99eZiQbKaeXEZe3ziXBJD
5Q7Bzq408R1bk/yUtG3m0zKZGw9SPPRltUdQrfbpVGY1xhfMjzcW405cASjPchG0+hebnM73zhYY
F8RAZPKL/6wdeJXU53/7ogjjnW3zi5eaCmK0hmedQ7a67BL8/6OybtDGtliolqUJhRxvRqSC/+oa
n/0JVqltjj1f+oIpLxciAUeXRpJUgo+j7+nX6+a6iCKovQSrUupEGnMZo1MzPhQvFaOw9FeZGogu
FWa3kVbXL/F1kqixBEc1FavZYQlOHGQGfogRzo/ecz3r5S6IfYu42h19YNd8YXFh+EXsqDicK6q5
jCCdFNkgcd5LZZ8r+xyX5upugSjcbGwiiIEhddpkDKB162Zv2g26yWBff093EvHp22BEcOJINWDK
XAV4enMdt3es1aJgk2JOh47mlcctMYbE2P/aF4IcXP+maj4J4HZKpRGtxVSxZSZOtGFiDM3vPtu7
g3VNIx/Gd/LEEj/mIFBrgXn5BKCMKB2j+s94kpS0zCqRvYMd9kMuUR+xj1Z//rs/6gIRQlTKvtyz
qzvRWRcHFMLdi38Qr/3LlfroOSZVLl7cPvJHPEUo8FgfRyRbZiYEV3ttukYHmKzqVqNmseytnWKZ
HVf3DT5pOVQUH41TnTtD4/w/op/4ZImOKS2AY9bsIC0HWxYyEF97k0BddPl2bQ2IhxrcRweBCMJG
XGeKfn6gCrtpizQsY6ZNm8pQQxpmakmmUbVcg9ProhLFxTOlS4af5kdaUXZpAaIxpi93NQoeEPnB
bnGLkrTVaFLwAfPA6dvQcEeMS0HtXqYDbgn0P02VacSwEnRPmPuvUXIs4Ezc8iAcceojN3I+JdUU
5ZIDXvAhiKoD8lb62xXFBJXqt+nL8BIrF8WahR5dPOlC2F5UPC/niDJ7jme8yb9FCsc07ybK/KGI
N0s7emjrqOI69Mz3urU5vHyMtyfJxDcL8i5qk1KTPpdHAN+oEHNUDMfn0ga+n7irW+vgjjW1TwdG
qBeVD/wCQNzhgBZbRgYi5ZuU6pzM8vVkVeSk/MujoVVHzpU2jqoq6IANB8gqqBdXYJ0T1H6GLD06
j/A05kHDfWUb06CwXuw6YEgyoTNalz0DxbM/NCqp1y4D2Ef/TBX2aue7dvmpZV6PkdwLnzS+JXqL
LaotRQJdU38ROuBgeFBOYVSQ0P+ITpT0Ns8z0AfvEi7sGQoAnE9izFbKnZQ+OomWARKRiynAezHX
OZ6Q+apQMhM/gV03OC/0Twi4Dta/ykDc/l9JV0z9OaVYNv2cmd26M59gOa0AYM7wbt/em9v6Be0s
WL47oDBKrcRM9onintuS/QS2gUsnFSeq7/WsCPykaBheCacC9LA9J/ufKg/6gwc0Nj/VQAI4GUnW
ImV4RKDi0sYfg9ct9Zapo5slXX7VGgIcyUNjoBPs6MjjljDFUcPO5H+n83kkDUtrMt8Ze9sP2m4V
xx5JtZhnTMrDEbPZFBD6a4qjwXSG62okmf7zrB7BH498lSPDn4SfnbkJCOF2Sh1pefgyeTrG01Xh
q7IPwbsoVncRDrMivwkI5q9ih4UTpqRnp2sPxUz9hlmbViX6VDDmgtWwPbHrhV2Stin2QOUOOW1X
bVuPM2VSw+PiuhOQLg0gJ2TxLOnFsSFMmyfXYCLV1PFNSILjrrDiZibcIgi31ELNxhQ5X8Pq6KS/
efIC1cTrAAmAJo0dgoLIFHD5qVrtJJ/qKGoQJdy/euHWd5NpVTFIoHleW6Asl502XNgWeQtbgm52
FMXs+xvia92sCbSvkkG51TlQu+JXgvYJaQLa+IDzEkJ27vmC9E+0qbiNczcqpelF3Yr1YOMLKvGR
t92OmeLy6BDl4tTTUOpwGwJsOVJmL2IYMAPuJtgIgODPJqfc1+G1ZXUnmjyOxYwmcccnEnYba6qf
oSCBfH2UiMD/1AUIYLcFBZxZqS1v83sSDLDYK8DFCoL2gG5MXOsbmgNQd5po95ggVRV2hMda408M
mzulx2nPU+lJVIV1xj1adsQI35hGAz+LPZeDyXU2OmyStT3oyJGu6jWTNLj18IU5aWAX1RW0hj+a
1XzRlC5dx+de+AEQib6V+aWYn3iLYqYMvHTviZBk6NqPuGaK4prB4jbiGoZdaP1s6qngtVPhgPdS
E63nnPegIc2eeEQ+GU1BBsLuPNd9ZfuTVjObfZzko5of7qSl9MAQMhJ+uqAch/GHKbLqEimjvARq
LFVmAipUsoHddrnfSU2ewDmb7bXdWT0sRhecDewSOXPZuayj7iAp5x+A6pMHFAa6AuUHDWTUc7pv
8jXzfktJlgPVX3PpvW6QFasVlLWbxMQib/W4/7xrwd3ayQAdD71TVtjmddNmymfWVPV4mFXjRb2p
MT+OPdiVlISzXb7ZOgvg/l1T+ZXfVv2+LUkPesZp9u6cbeXQ6HONUEKuPcRN2Hq5ksF1gz42Dk2s
JPn4FbzgYhazHjLVJL4hASKeuJU/Il8Prpsb2z9kl/Xs9+noML/z4Ksl2Q0Urr4ao3F2JjInlShe
YpkwWvBwWdxj3R4Wrhy7r1ZYV99UBPq6hNbOYuY0KC6MCyaEs8UMvmAA3lyxFxHJp0n1k8Gy0Yfr
eE2BCNDJUcSVTBN+Rzol/UrgMkkQbQCTC+z3l9zcp7xptqNIz7jEb8Mf2NeipqmB14Yf0PqXkKr9
s4tCTS4qdOU91nvGBbRjlLKTx6HjB+/6gBLOfbePd92OqMuZ8w+tPWlocCwM1UHTc4xt2CS6AXM4
sZh7VuS0CU3TQRCSeN8xs36qoT2ZD+hXyUOUSG3PKYv1kpOGlg0LFdlltciocBnXmjENBj4tWy3R
p2r+G+hJBm+k+FCcs0ttxg/vULVQit8Drg0VOZunym4si9SQF0WWwcFh9R4qchGUBaqKBMmwGJPE
Z43sfIgzmmTzG1GI55X4AVhozEvpSb9/g0AuB++FO5lyp3i8QDyi9l4CoKumCOnqKo1A0jQ2IExT
suSOFqNPBgDRhXDp9gGYd7G4Y6hDhwFqFV35K/iLWOB2omWaifcTAt5rc3SCxdUmaICEkuIehAaD
+SHyFHbTRJyPxVpGnIgShWEeeD5FySWy3OPT49HYEDiw6TQRKZYamlbbwzzAgoUgOVphJSmrsirU
s93MIZqP7JMnQjZvf7vUyPh8kpzVhs1cYnG3pADtqL5lSw+XQaW7vC4OXuQ15Y4QwiW69WWaQnZO
5IetQpx/g+AHKb+8mw4yD+UXzmTHSX0Zu9mhMIAngKb1DpgV2wDk4mg5HOVvVAs/3jJNniUPakey
1FkMtC5nMYK17E7TEz59WPBeGZZecLP3WeOOy7XPjhg8o0QwJwddzIknzU3U/p/JXr6Bj63Msb+t
WEo2UjJSnn03KIHZth5ixqpph0pCjbACjVpwaoM6ksOE6KvWcNiYTptzBi9StQYTz9cNO56UrCN6
hdCngw9eOxlO9NME5VjRFpOfnjx9f777GqKmcecS6FGIa7Kvno/yNl/g8Xz91SDiJlqepdGhqWYh
y36sOes0FRLNzhN3ChiSGkOyhq/0gIQdWxREWe0l+UmNbc4rGz8tulxF8Veshq5JP0e7dlMhyStB
95A2iVkrSvZVK+GmK49nrunNHtt6KiNsuTAjaQuPrY+4Bbd6prZQMcbEzQfmJ3jxWlmXXdymM6uG
yu9XNA+Ilb7qtPTQJdgHV7AyZxbirq1m+UhCv4ooUlZWEQqs1kCBvh9i5aY8C+r4afG7UBYlHJUi
z7thxmhvioDY37mmI7ByaRukA45hRiCvcCbZAeZ98dA6NHzsOJ18kivvky4BA2GyGDe/XOt8JOcY
2PdLo3pOz/X+gJQi27ovEeyktS6hsIMK63qGS6BznU8x83iaNyxRrFG2DaDTNExL8fcex9/n56bE
wi4nJJEIxkhsfwWKg1wRv+SWa5QI/idtPzsqCJhlQsCYhqmhfpLpEuzho++5GDGtDtBxuUhlSgkz
85EKDnAcuzFNOYd31QB1h83TI100tUUiVVzJasF5M/caizxWtIxOOUs8KHZiWmLteAlYGSTegG7X
n0K+lDANFY+EoA7Ul+7o+HcT2nkyud+dMQu7X4DJsIHtkrrRupV6leoQyMorc7KLJua1OU3sDu3B
Hthrz2Q6Y5mdT2QZjl3jV3hIcH9DZQz+XOUMI39/+MowbSv6PiQxmS1ukY72c+4zbCQeLwmqXZuq
H835sI0kz/hAzkDypwcBBEUktruwPA+hfjN2UwiaoaNHVV4f+C9xlFetVUUFgiP5RaJTjCFDvuLy
k+0BnyVgdREPbYb6X+77oHHbTuUiaMVSyD/gIbx3Mgufh4GNICzR48HpDOUeH56gQxMvv+9viLwh
UzU1QCDhlbl3CpjE+nohY5tf9IwFawYW1Trw1xbAhdhdljQyzZ2gLvIjkGtSiztXszwWHO6npBKd
H+GZbZjsTavUitfZ/vbBag1HemQsYN8D8ZBZz+6oWz3b/0yNQbPM5ZYACSuQVZwA7godf6/ZqWak
8eggVU0OwxfF+WLZSSaKHi4nbuDZFltd+WBA7YgfXLwII5FnzO2g2UCfQklhU8QBc0tEstwfmqZB
d4WbgOx4tUYBLbk/bPE8b4jHsGZc0I5MYpwZGCc5FE6XVzZSNQsS2btlYUYWIpHd9djz8tJA8X7t
m1YPzlc4zTq9inugFk4ml6W78hx89s+6WZBDz//OVHH292yZN4l0xxSnqNn1GvkqCD0zovHh5YCA
gQtxDEM13fzrgULkEq8kHDfcrwFMpv1NA1QUvSUn4JLwiq42biPdEQ2StzdUzWFoCDXg2qvyNYrI
lFFYHeYJSxH+8LLxieNGbKxa2R+kWwz4EJu/NOKBlpMoe0ZKr64e14aWhGadFssO6iHSGv7f+Jz/
sJTDzRXHNhci9VvzPWHe53q37GZtQtW4kJNlkl5UWEb8WZ11TBtPXsUbN1J7ZnUNOB6H5Ip5r/P1
BJznv8MVCCrprCHaSyg958cvDmRzS8Vez3PO43PdFURZArekidXuHSBz/CAYzFv1SHwM9eBESyzt
fgQFv9u1WnF7sE9h9wUTQOcc/6hF78BII+C9x2wU6BVYvYZtqac6ffnmVucuiwY7FDAlqPA8lT5r
VHDTj5PjcK5ij/0uUBpQrCKODMiZ8tsc4A7lvQ6fBTrMI6hgEIfQwA07kJMaryI+L/Womwo0vrjJ
IlOaMqR1YBQL0WAcgsG59933CFuEb5HpZ6raKIJx8T809v14PJGEO/TEeOZecpwxnPKyAQ9yS6g3
ufywJtNaVyJwxhwA1SFl/9mdoSCeR9vWMnAU7Eu2TsvJAFvYLLcpeXqvqkXuZoSOeYZkfVfF1om7
VkIHb4CMC+rErl9Zupcro1dJRyWkLWmsr5L92BsoeOKGZLG73spzMiyDVVAI+VnMmexlkU5bpx0v
BJEGkRSqDYkIe57eH8JGdv55RF7uQ4kly53uU7lJIa+4Tdlhezh+e15v+oEs+xNEp4dbWvej3G9x
ilFprzHLao/GxOQkKLSnTV9BqhvM8WIO+x89fllM+y9Ylo1urqohFmJz/1JuLYMtgkS5DZBJnrYC
BYmXOT3/bwZVMHDCrkrWZfnMy+EtQN1P/q33OXNzZ2xe41hEQ+TlpDt3IcCuhJjIMO/ySPAI8CuT
zI/5BNyUqMEQCBJ08cKwpbzo5l6AT0huqLBOoZAL8FblmgGx8iZDdqUeWGq9cYOQYVpSQo4acMZb
GSH0wbQAvu9hTU1nwM9Vt0Yu0aUzVmeeaFpgyP3PniBUZjMBUgs/l5IJrGUubBNh3E4V3n4FT5g0
vZy6JsYHxBWFD0DYFqGt6sidn1x6ebCt6ohwFy+RZgvHrjafsFpiSJSngJeR6s7H9fJ4BE9QCq6f
YEUDxyhV26bMCmBjPi/BWZ55j81dwiwSs8nuVN/CL0Yb2RTLmZU8OOtra1rq31o4Td9WkOuxy7kq
waKqOneE0ef5t2lfqg43O5VPfgPOEc2jZhr2LHnkRdrMviLpcpCKrv5DrA1+1/GJz7XcM4aJP5UR
wcPdF5Ly4yARzTJNHvrLSoG0owGZHdlrbdiJHMp0FB/Gw6qMU/Pdl/XOk0g5pJj3VKMU0MokHSMS
X5ljnwe8F5eEriVoDLuvdDtlZ2GCcHrOmjH0ljRPzUb5sTyey1CuQgGBykXrPiuqXCzGA3QZWrSD
9RbyF6zY+JVHcuq2pbsrDLRg9GFXZZmaili51fMfryUmwb1GM1uhAWc2nPUAPZwLxAT+DYgv0W3N
jzVBgNiBcYKKNkT6ZOVSV0DcPReYnMVeeZLQZyWbLHRaHQHdv0ykTknSerma5A5asmo5HwTaaXT1
RlC64M5OOHDG2wVAD1AjzrVjRlZHIEyvbLHkCTSEG6mwaaWv7mYrIddrAC8bhJjE5jXG7ByfFHI4
Kcnjc3stycg1bg4icNY2uFrEWxNs5x/yJpTeHn375mzzWflZJZSyB2LEBPGUgCEHzEAbixh1Rzd2
kwvpeXvtmucpijBoSwcvVgakft9UG/EqS0qDyDgLB9UCZb+jN1VIt4G+Uw5z4VqrB6xh7Ql93T2I
wcg2AFu9dqsxr1n0+XG+ZXxJo6/CC+Ni8imMd1t9tMfSLeW+K8jNkbiTStPnTGegvCC5bitjC1xM
J/JKytlvSQhrdFc4tEqeMgj2MPxPeTI7Y9c5XnzKpMQcrrJyDB+GGbwiDoY53lGRwhVr0A/RlHA9
ulseMpEuZQxeUKc2ueYXrfcWRDyDhH8H/2/Z5ZKzIt2e/cnwqxvjjUlsxtF63PsrSVUNGpnTSlbd
KLyycLTypQI2V/LEvM1R0jRKD6fnGZ3uizGt0o3HyYdYxQZEY2xzS1SYnu1X0VoXVB4JXDi1Ccr7
ZGBb0oq+y0DqwgfThDvq2827TR45jZr5Osy2w3iTB0fPlxeFHm5cEl/14BM0xHB9xJLx6EBcb08s
WfMk+XSEKLJGRPZuoObFz/jJ2wVtEW5hzt2+xltPl4hH0reKy7KzUvyGWxoMP95g/y+3do8sHXad
NlxhwH9Fx6GsPJgq2+DyS6GWCiEDNyEfg5HHC4qUP92lkWCuN26w2mPhcy2YAeqhr62RxLJvAXag
XLylRtUlNTOzzbliRDES2BUq87re+Muho++IK0l5+7g2zLm2gzh7c4gnkr2pdYObWhiJyASQ0PWq
oeXwEmvgCUzxsdnThwf6sd5lvkYTI7JLTcPl7aOX33tANfMHOJr8eAa9tOQ1yFWAW1BoAPJS+wMJ
xrLsICLeimraMcG/qU1tDW/uKrPlWPdc1vtAR48CmHxlp1CEuexKooj0g857THvVRaeGkjS2b14e
TgnNbCQKE9dfXGnWV9wXHCrq0rtjT4On4IzHbvqyYHreA2ddLSrhQcUQOBaSHnsGppY6kYwh+WRd
q19R3tYNXTpUBP+ktY5zJCgp26jVizWJAhO9b9HJ+5gCaESNXOS58hqKc2oOkHJmkDC3eiiGogZH
dHCwDpMNeuNUwSo4UQ8VG/yXe6dlaM8vQfAU+ompfr3fQuvtnfXDp4Z+kA8NgknmMblkgM7DQv2v
3lyl5ei3URPOYV6VPKfbOyUmD4Kx8IVEvkim/KaZI7hen3bTt2YpgSu3qeePEGMjWuvEx4Pw33V+
p9v3oCT64jFY1A2WjeN6HiZf6N0Ho4+4nVvvAy46RQk243LN8lcgG9z3V1exYeRDUbd10IdvF+0l
Bev9BElfkUPZWGLiFR8E+K7/Hzswi9u3xHjKAeQDCsDWxKNwyDK/dRQh+6lrizDLGNW+xrQhjFtg
b4qt3HXFcT5u67VaEIzdxTR2/GkL2ANz0TdFd0n/e4MMdDePPWvzlmguVM/lxVxxwDMWxkV9IwTF
bscecQVsn65FUDD0WXk+mdFNM8WGftidS5Qw61K5GDkTFsJAuybhwVV6uYe4SXDFzM61Z2up4VXq
dSuznsp9eskSdA6BBgRZigt49FMs42NaX08T6quftrHbZDdoJc6uf3tzAzGzuGLgs6NS0wIeLCZb
WKbRVfFzK3gpQn4qpLsnU7zKv3Qf1CHHBpxEfjsZqInSfVtAOmgnipdjERJ+rK0ubGRBVhXkwHJ9
cvzAwoTv/tlLoZCYBSr7cJVkhb8Vf6NmiSfKRTHkj0WV/50a/nf+wj6QLmg/dauqyKKl5q84kE6V
ie2vrCJ0XEbrltyxeXsmrPZG4FSjsn/Yp106cBE3Oqp2ilBzPi89MbIHm1AJ6YUETmwFaKzy5Fo4
ldv3VCbM6vaIUBpMN4iOvrmUgTgZlEkbruhAsfFegLvAtM8ozA+qsznobXaRJFXcA1P0ZMpqKsa1
9IuW1T0O/VMxTALMPM7VA3Ixesv9hFtPzbHoMq3/yfeN6yjrfFt8zeugpQWBUoH/IW8RG3xuoU2f
4xeAAWBOrK05lQdmJkVIsEUg9acdy4H7QGXU39cSn9lUs6jJYityLIHZnIh+RNhkGs18aFA4xe1X
Xk3q2ubaG2yjjza0P+Y7/Ikiqts+tcWHggOIceyUy23sa28uY42Z/bdvExoEJslS3J9Tsj1/dFBn
vxZFzJNWZvuN2gIxcc+PzR75BHe5RiyWDMfiOyWVrEaE0L35eswmNR7kHakGrNuz9LD2EfLiA9pV
nOUb6mCPeh/OMSOggoHFSPNh3SSSuuZSyO8S0WnRD+khlHb587PeaVcJ/92/cDVWR6JpmMgKJJmG
jdx+fPvj3IYTG5kT+J3Z98td1qEvvYB51xp32iPdmHsrGKsSwy7JgnoijgYe+6jvB2Z0tkDZETv2
CyXsSDk+tHaPs+DpI7yyVwlNx4tn48eM93IFbhBwFudhzpDgDleVgHKEJ4SPLF/tp+nT9CpHu3FQ
rcZuFxCFPtsBUNLyn+J7yREimmq+I1Y14yO/MihHCOo+CF9o0R+v95xA4Al4xKeu/2kakDt3PCX9
g40jz/FzBsecVYjToBzdxgDZpPiKrqtg0cPtBo8zkggPxY/vup/NfR8rvE+AtUP5FQ69bbKSWKLJ
VR2qHwmj78aZQ8wkdhy3m8oMY0HO0FPieor8cUi/mTSc+d7CGay879rz2VeR5qduQ/SHz87fj3KM
hw+h796G0+Ol6k+gNReH39jRRqu0pe+AAT5yvek+wnWl8Ngr81qPRXaBjPWC/DSBEBwiBJ2iO86c
cgSOoSQR8iXK+5JZManFFF3hkJo67mNfG05kKx51WAIqDgCrQW1rlmgje/+b0BzUcYV8Kh8lK5zL
SgTw5JJa5qGnwQiLxCRnaltVwHrEJYNcVfU8poWb5ezYwqu4lSiPb/J3FeAFQWwVSU416Pia5Lt4
wrMPfq2zhXPnjCR6AV/WPiPLJIwIMe4SRdZ9NUvcdvEzHcOSkKDfo4tPgKX4ZdDOu9ZVAo06WToi
oG53OSD4qCDfOcgYwuhhwsCFlmc92xr0pFldTRd3GJktOCf023ED0rCLBbmjRciJEiR65JydTGpb
XLe82RJZUpnv/beLMbeH9lpWpkAlJyqmn8UcaXwvC2rVkA/1eK/DUnQgfSovOszKnCYc43nw6CGE
ejCICAfMJw+P3oWciACDQTjP57wLyGZdTdS9eYTabKh6ZthwI8PRiNdbqSdlf6p0GBrX8t1LmsIG
XMkZivHI/siOnlPHPLLApjnRxl/wVnDInrBVJ4nGV0swtYzCGARvHUEAlzyD8jxiQljtGfjrz6yJ
1MN68xyVQjp6cm0nD1IiwrPeo/TPspLvjvXcn3dN2ox959zV2z17kezROrX3GwtzFKANb9rGyvDC
ufYbi1U9RtaMiEblrOQc8/Qv2/s/Tp2JvR9qWwwI3H3cvsILr9exILRP3kYl81gwd3svhqxMZXGN
BUHw9LpHTCMx87Xpz6WtuL87b3rje4HY+2bcO+wtBYoico02KyiEm+ev7xIZ88OzX21Otqx6C+1S
EKHCYd20/iDz6RIttWA7+dakEHtuVLYzKwyvmmgdQgAS1OT0xN1J3dzPd0TZPrUW5gh11U8PNzIg
WLMD9EErnI6E1YVMPegc3i7mUsKWsncgHloq+WAbKQTdzLQ//4O3AHy1VkcSGvsyKrCJdDExRW2I
hZmI71OdeLm3WGOCnrwAPveENfYjQYhav9oUwQsd6zpf2S3zDIn3swBZdUQMjd0+QXatKOrKMGAb
24v9H1Uw5GJFKSyohXKTSss4OTC5n7qJe17IZ07jZxio1i2dXTNCI759KPfAmTzv3QcinmqK0Y2T
+FkiWJKBUG9iNyz6FVN7diDQCtNvcb/aGQ8gtOSrgIhDtif2ORoZZu/cHa3Zkf05aY4qWejGb76m
apJnrZlK9Ky9Ynoh3dCMPE/SEjaxPUu+v/VMoTR7JWrNZgw7vpdkouyXMzBQ85UFENn/GsasYWNS
JOfvTt8QskLRQWAJZOLlVNVNaI/KiDewdsTz8FLnA2kEzAaOac9weoQLeibnguBz0caJhhSs1uav
+IDcUd9nUXtDEnnPILspmvG/X9IAppnveeD9rPL6RRyGsZT0iDnZnoZ83rZ2Uk0YNwCE3UIj8jv1
kOWnUnY9N4gyNq92ycyLUV9WwiZ2RW3ECeK9+aNl9xPTjMMOoL53aX9hwAZclCAt1RiR1JWbQ2u0
i0fDkOYr6akOIgyJyrNfQ5UpE3lgHMXZlpyft9aJ0cOYWgn+2JKWTtnifA2entSxo9X0DeA/esHc
QLHujYtpRJOF7YU1Dh1zP/wmFGs9HrVyCjBc03+yIeQrAu2+7tnsqNEVDOX9WKjnIZ2bKnHKnTrM
yGVqp8PSemg1Sr8xNDT36QEJTRg51XrLkdIt9bU7H3HHLfw25p3i9alDfiC0nEmhlTpfYf+UAOmI
hKwC5cKrecqTr2sr/G/b8Wy99S+iw2SsCxRECgyJQyof1ejAiIhsGaVzm2877sCgDeH6dPIM78Pa
E/utZ1Goz5CVPAPHm7VoeGC/dojWU40AtA6b0+8JiJUzdTlRXZYMG6JmTY6Fb5LSEaRtxdudB0F8
Ji0IFHkCmNOu1ITl/vxxEkz1bTUUPkzX6YCQ/iVpjZkQpy5gD7VWoz3Rd+tsH5be50/g3Iy19S4M
K8EtYWskreDjym5QdtIfrp8OFmeLS44dAmFin9StWYPgjst/wU1Dq+ICCic2ksYHLQNIQhIwJmav
f/yfAxb5aDRQoN8HkddYVgZnYv184lRSoBtSk/Uz8fGQUI7qZp/zgYTTrQwMbAAPw2L8a1ZB5Iw0
UTsnx7OfUzcYnMTlF62eFNalshRB/BIVpOC4leJsYJdnxvRG//EwyQSy4w0M7S2nhJaVXkKqcoqc
4p7K3qVOBPEr+zKMtu+x4WuxGF+yliPCXt4HjNO9Z894gPDA4AtLI5P85Z7Mvamgyczr+6J/cS2C
Vwd8z+3aKFr+wnOI/V0zXRK0g41n6YZHqeF477t+E8eWEG9p2/nmsNFqvS3kXCCoxh94qmYljutn
JYuOY41SYrhSure8T9f6YFaB77cF5OHZqkyry9t8mwipCzpXLUKS5Iqi7LOhYVHeN44zUYDAYVYo
d3U2RsbjGH3M2WQns3MW+foGVjYiSsGsyDeBw9Wi1ywd/gr8PtXSau+aLAta/oIohSLscfxzpUg1
FwcD0A5jbSW+yy7RHXdcvodwcXSWnHX2bQPzJfwZEbDOmjG8bn5O9sYv3kqlHucTp0Rs3o4EWZ+i
kyCDDNXRtV7bWCc44pyCiB7jWGhQXmqlvr5N//9ki50T4r0BLQnwMpDLMZY8g9OjWZ/8U4ZzADSN
9OWU8oS/gs4eEh/Z/6RJ1kNrmsSsbr7Y3xa6ctSciHCtz0yGTF8ArnWd6IlBLsfZgG75YIhXoYVi
Jg0YRz/0gq5RJQAXHi1ELp5w8F3Y5Nyc4Sk7ONEaDlv2hnbzuU0ku4G8flCzrBnapGsC46GV6nHf
R9puAjnMUcoGYc3yX838TS1qeU/AhS5MJlWZSHpjg7K1ijX6XnY4DaSVezU9TOq2p6kNmeQY+Yqb
c8+iWIoWxp3SdgaiO3e/J+3Fc3Xt6WQ4LlklM3WicUORextfaDnytmjvkp1do+mWLX+f06AkFM+T
Qm3BbE4Zxi/oc92DmSXgBCIiLu1jAtPFbu9z6PwAGPcNuX3Xf3MsAA/R5ZzWLuk7eVpPAbFzqpw3
VYm6qcIbUs1M9H/vxgmiU+0J55CLkVTiUDtvJidSCzYWoOZDq/zFbbYsb5WQlzjaxxg/RBmCv991
UaIZSphJNnekRn306vlMEuUup8BTCxhAASghGK3SCodZ+gfiMEnUwXZ4rpLYNOV4fSbDs/n9kxDG
V13bv2u5ZeyqczO/Al27v2mNwrMUTKhLNLVYXRenMmknqvJLJrPZ7pGDJKOJPlcDkVeXui9DOM0w
lTdhd2TAVYwRGDDIWJM7xvo9KrQKsG36EwJZpQAECUjgwtS9wXcooVzQE0S6K40n2GIYgsHCtgtl
yWh6DPKB5du/AFN7b50KGKiUGs3WdblTFM9EVPozIyij3YJGIQosgDBI14BJoNggcRYeGIRn4QQI
oUoe3Q1jdIVPBsOXEBS1qqGX7eatDF1RPoDqFDOGTeCg89ERo8/KbNhp/OqteQgTprLnRdDhkyEg
8hG9YOGTSs6UdBJRguaUnlhY1VR/Wzc6siX3VBf5+99OOTp7U7uqijF19BMJJFexHoL5rGQwrqPm
SQ7heBT1i+1lvnsM5joik4Vzm/suyNpWRgz7ArG0JO0UTpY+L25piAkTLQdfsTHwdWa7pb4KPEqq
MqIyzYZprBVcY7gs/q8trIYiQJJ5p1a3ys/WtGAhahZxALey/hQUciSUCKY9Mmm7y/SCvBOTehlS
uXy4syDYNxvpVjU+7vHJFuHH8nTN+9QMANM7SPejIrOmj9WfBtbD8ak/77gqdPq58ebkb2uF/frp
nGC3Eqm/4sSgPfQGEHJh9S8edulHDcxPsjdhxfcbt6Fnuf4HCCVHUJP+7Fnrfw1Vk5+99bVDoGqz
SiwotXrE9gX9+euZt9jMuiK+PhvClOUjs0Qq2MEuzOgtbsJy/qFQ6138oa0m0dmCQ6FurxqQTUT1
GjjrAOtz1I47+RiqsZirLVh2F5jAethFU6/8oXKfojMapy5QwstEVLkDtVxUSNryD48Z+JnKH2xE
j/yOB1iZQEYj4PxKm16n60q31EBKruvwoFsZBRP2wuoHosyjoXD3HGpZGlaUycqK3vK++fVIWi+a
TAvCqDsveMh3u4RhpalT6qCke9mNd2n1p+OgioBmMmSvdaCF9Xq89WZo8eBFXAbhyzBsUwOHjaZ5
XPRi8+qlWoH2SEHHM4rVQ+EpNIR+dgBgsR7hSKTYhKYrBkc4cJZ8LqqJSC0kFHli4DD+cHJx8pK5
vwhrXM72vRJ7AgDYMW17JqH2uTRENaQWCEEXscYGjp9JA/LDmOVj9BiHlDnUcqQPev94+QaPUvYe
vdxnbYCtxCM2VSf+I+T3NZh8a1L4Z7Xm9XqFJi17Tu9IiQwqO8hHDMPhHgMZ4QNRrkJNNPRBN19Y
CNniApvgNERqKQokYzAo/bERTNYD5yqyJ2tooBq0nEjhUs4NLbSpfs1PcErajakKYAawI7pCgqji
NOT+j+EFD7cNtV0WSbNIIiGfP7vAfJE6zL1PX4rh99q/9acsVlkJqcSTBwHNd2LWIoRjx0SmEMDs
OWWxYbSQqypEb4Pe40ObABnzT1x+U/Sy1XwnyKPDb/kTP9cvBzwaRKay8ELipXbc3fdEf1BMofmp
j050Y8VhCd0GMVC1k0yhYkH96OUUCoR8NMG6X2srtA36CJmjD6+iIdF2gWOG08xlz4+5MugPGzgC
FBrbwRrmCpVOXGapT2897bxotXhJd8bVRapcEVKF8YAs1/Cmzpb9xleLQJscnhtN4fO2snyyunXs
PkFMictt5VTiilXkFiDZP9dptgCAjs1rTKeMmXZC9F7s8Ips+d5LiRu4AHUJAqNP1RFWOBwyb6ED
xmSSeHLTpjTvlf93+p+6epeyK6tAXjtK0YOYFF6MJwr+qRaZDfYGgXirQGbqdSy7MSO7TYESsU74
vOO9hnGceJgkmoyn1j9cUBKNSGxkbXS3HAxlWuj2kZmrIu7WGOtJnpOi83HodwsZElVlkzq2O1EQ
Aq3tp/nWOymfBgCN2f7La6halgSPeHZQYr1CZo6F9QAn2S3ogXrib8FMLCaOhwV2gof0n4tmYVMq
5QIo81sye0CkXTPww/e86/QIoZY5W+0I65f4KOqzqzCcupUCbW0AWhovSpIOEgbdlJ5mK8ikhExQ
+tNPJLDiunmg/iQGE+OMB7/eAz98agGfq6YJsMtB6yqmKLvJZI5b23filUW2BgCmo6CET2f3hpil
uUE2AdM6sG2ay7aCFLHzTYZuzAA6DVbnhqbeYfoUdrE8RozJWEm7ZWjo5QX2B0FRuOaxDkBpybIv
OgOW2d+2k6eHLGlOGOlyvx90A+Wg2QEUm8DiPYso3jD9VuntLHX/BW60O5oHTKt1k0MNiJOyqr3A
OV/GCUhhuqFHFyYuCAmFYJCMjKCS7DiVDEEA+vIT6cciZyx5BWPfmeyN0KjmPXD3XlVPyhqFwT0Z
Q2DdAa53JenFWqxr4FHSOBuJdPV7T776R02EoEiO5rlCEy8Hy3v4g7HecZCJMZhzCTZFISe0tCzL
rFeTDzDePHXqYKmOEuR4EB+3et1SP4Pki2k5VT9mUQJ9OqA9twf7zQh/2794FeTr2tuozDJRVRmi
0UgYBQ2XzyFOlMKEbV6Bjm34ZDemx453VH4IUsNEcgzXzYSDqj/PRNU4VJmn3TeoinOdMiVUjrSk
THKBDFa0jsF2m5jEbu1EwAK2dFpeSHjiwX4dj+flBTeiKhRytj7AGr9AL1wWcw8yoFuGWjQosZXG
upk5vIdMoT9Mho3uoUDskg6o9+O8Qt1JBQ7TJU8G/JsEl299WHuWSfPCXZBxdZX/7Nb1BlW8HpHr
2pQyIEqcfkIG08+zVa4T1SyUcYq9qdOvo8ApnyshHRen9EEIJJYQBTsmm3V6yA3C2HPayymGBvKK
/7wOA9yLWOKLZbPo0lMbzS296homnypiZ9JVoJlsl6F765AEGG8DZzQa/oFZyhaY6gwZS95ih+3+
J2HY3hP/iNaUNTaQxZhRUXbWVHodIN/gcsBvlqqu2CJVcqH9Ljj2TiWHwxtLXdyq1JLuksdjJX+T
pGJPIMcoXXXVoi6eIp5QmYQ9hDs/zzxmkdEeLXm/bhMLDpvzc8WY6z9pfUQEn60zyCYmbp5hzYUd
Nz6Iq6Xh6bGGhYxRp0hJP1hlgfUKLEUqqnHi9t6mEnTvJBYluainlZJ4SInWcTVFZyT7zIUgNvP0
AXaxRjo6CE5komNlSRUDb51JATW/UFMGH57rdUwXifxTecIPG0Q1H8hhHjHrQ88ar/ztiJC9dD6C
3n1oCFKTue/CBTaQwOkEDNf4fg3ILSTp75Ii33c4FR4S++dmNk39yt6ngOcAV997jMqTlDq1ACAH
Vfg/qB4GHm6eFa7WqYwmxREHMNP4MRjHVaYctESwhZONyBcH2SCVcKRedJ8932bD14z4JX6Xuons
G/nMwhTpMShHwqhARKseRcnYHuGxoKxRvvyoF7qk1/+1f255l6rL/hTrM9986syLQuxdmat/TLHe
dI4iqxP8o47MVvrwH2jbobY4yjZW17V2k0CoVo9IHRZTv/6kV2gz2fPVsQAc0L+DLm4gKmXAUaLX
OXBB8eeUXxTg+8Awt3SfQVi/jUxg5GybxEFblLb0WOPiuXqlBCRhNAVHZ2/C/lHW9Q5iiSqhINHi
n0o88lXDB5IEbI4FDvPj4tX/J5wFSvxNjmAfUNtOLtdLp5m4YVXBpnwdzxzgMdUAeDQBH9yUp1di
XNEhh4/XyA9Lvl12t7liFy2FtfwuoLGpnpJy365ZUVHyzZImUvWOqyhNIdr9gxV3k8fVe5Q1UZR2
qTWMFflau1vQfUpDgfEQ/UWhqyvfJ9QVBiZqJfUAVRhpJalvL8Fv8jDAVpR7dmzIEQcIMOKGk+RZ
pE/7nQ/oC7V0BDWDnEA9BT7zf2aWJdXTOApgdhNmnRew6bGDt8EDimMQeN+YhxMdbmTIL+eK8ztd
Fij/C+WYUXurgJnAczdODoT/kVgaI4lvw8oA/dSnDeYQ5+Aq+BBpjNLj2eTC50lRy/u7fMcweDRL
sxuDEuy/qCsklITHbHA12QyC5/S0obR+5rKUzDPoDxBt6u+A8dyYv2Xvcze58fJyX8YKKR1iAUCQ
p1VJn+hyync9WjVrdef6sLq4/h4XFKBBo1PJTG0GKuJqg4MybI2JTO8FZ0W0VwLKtAZg2yvUz51g
VJsE6S+exJO8Xa+ypJ+TM9p8aB+gqkbWWa0B3/DiJgHOb54eWKBR0owXHbvFgCBIhAsSHhj8VRU6
dUxoojXmA5IBKgj4ncfHlJVFByRtTzT5XKOGDfKO8oosnKeLVmW2nTb9zStDvYHG2oNPBl+mZPQ0
d2EUSX2czRpMw3CcmUK8nBeVNm5yHnqwm9egm4C2+0T6Q36YUyvyypsCwATnNYAhINnTA9OceN7p
48CWT5jIvaIRm3zBkNCGsq4NNWBVccgmSBdEUQkZ9Ue1KmYQRM0TkD0Bp/zsa6MlFWe70j2Z2Leh
5q2f4kXs66VNCNSerjABTWWa9UhE40Iu7HvKciy0JQe/wN9iMzhk0U9FWazx2NzPLHxuuUhxHNv+
BJt8EpYklg5rukUOEysbHl/dVkT/ds4C/aGsjW6QN9m9fdXlt9+9w1RCCbywu3yovAjMVE2lePH2
HGAxyiyh+4jtEUyaK/QOvHFCOPNU9Xv9e5O5UQAXCQbaXwlwbYNWAVer6A3h4G7nrwwNwXy0nGT5
973Jk4jKVF+1HYflKqg4e25UxPohkxXDCo8HiUcLG1JDwUahjOLWVU8lXDxnaClwSuYdSSa0HaDJ
3b3tZC8Eghl2QTJKZMcRVEgfCu5YyceOF81mfOpFukWFMElYMY61IEUzcT+JwJXwjf3Gszq+Vei1
i6IVxdXBCfR+1V6fZzwgp5DkkjEUVVHoWA4fqfv07My67bYmlOY/lWHE3BffzjCVYYnfVmoGF5nN
7UMloQgN+bBzk6v3a8wOcJ6gPR64GCPQjEouKduZfbdtbYavuPZfn5keO1ieOEhLBXtWqCEhqFmU
23gbShKmuo9/EHt1PlGTmBWdMzEg8Shljqg/DfevKyFQK2F1NfHq+Izjhorb4R3ByEzHhFxbg3Bb
nb257wbSKXMIesiaE6o3ksCUrteyOPgAGJMcPIOuIMQEllWpg69+FtNtX4cNot+W8wc7wmJULfHm
U47RAHSFFVwkz3XETrGO3Jj79e1Y24nBJP16zPS5KI6H/tqqxnRiy8BlB0pg0sWMoVU9SvsAaEee
wcdTLNdMQmSimH2skob3xFgiTg+nD4E8Kt2JJgQoJCQ/mf9cVzPjLtDVzkPVMPcBX4gWcl/xU2fV
jpOKso+ujghWU0ho/6JkiKcUD3SwfQViOwMpHqwYgNhGYYxhiosGl0+hMeXgpxPwdO/QIyuYT8KV
MY292sJyyuZc6SDb+Wg13e8oxKyVCUEMwRK9cI/pAwcJO2Lxo0gdHMpVsth29FsdxfOoKSLFZM94
CmAHX/5Nzu7uu+Zoqki7gvByJOdd5o2Qt5kRtpGBWewgt/bhxoMWvCfwZ8xigfO7VCMjDB25V2sB
yzhBxGHfGCwl1iWUvjmgQUl32RieuOWu/aFPi4Y8E0h/+LJ0e+pYsbvYRaXYhknmeQB57G9OroYW
ea1lzy8wTQh66Ic4XVGw6wb/k1yozhHIlSsXEGZ8JQXyAWjm4LMygg2z5fMIx0OkCPzk96ZXd9TJ
HLJt2Tg7RlsMIBVKH8b8cXjQPPSm6Cx68AhPFOgwvv7ZLWwvVtrhSVyA/kg9qtx93Ci4fCo9k0rr
VHGqSFu5Lq+Dy//npdGiun+fJZEGfsUeWo4kWwkqgkEseaWv6iWiecrKuVukRQ6OnQyrq0aYhV3Q
7mIc+11tvjhNZiJ4t7SB9/3cXF05HeC6sLZXVcDNmfhRnF5i8VPuHIuogH3D+x6r/qeJC9aRVaQx
8+cMrSD5VwtqlUBgbttcBDkh4Xg0PNE2n0239vHJL+RcbN+5qwqFJJXEopx4pFnfs4t/y2RYQknr
0dgfQUn2luonw8DS0S3A8x5ZHKxY0uXDb6yDPMbB0CJziypY47xjKo5xdCkfkWzdO65AOrklXpDo
oU+b/nrm6QJTs3Gzr1+9kEH2k5HoPa//J9+ABwJwut+ULd9jX80hpfIix17DEOJfZfXz28/1fg4T
XuyMSqpumwvNUK+6JbZaYWp2VAgvd5WB6Wekn3bgTFRGSkrCl3/UgR+z2nutfcJNmTAeXXaxtgAh
I6sPf3kj3SwkPj4TNlWqVjNcVepG+aQu6/GQMin+xmj5VP1mO9taqTbIU2LoUMjT7NmmXu+vYh02
LLWYsSj713yptIAYk1LG5kJHfM4LlC2c1gcfLNoRNL/HN3NJKrr57iZJ/CX6BgBRk8ttfAFNK9Ob
ugVfnM/x8iuH29Y396oIJAvzjjy5EvrBV38FcrFNJ50861slX8h7Lhxl7h3YTrUEAbMhFhmtor4V
nEZjTXl1OqYL4tzL5LLAuY+xIpk+hcBMGT0CxbH4JAU0uIK6zkdkxB3jtne1YJltGlid5IhKaVq0
HxL/hGjfk1x5wDBhLJD6Jqnj5vVw6KWC1a9gidWmEsLvuXzMmExs+uizb09CQEmUqcSAKMwr1Ye/
KdB2RAQkvaV++2fKUZ8AempT70LhFNNrHkr7Pnd168BknB9+nRl96A7ZIiZH82F2N2m0GoOKo8Y+
mZLUIMWGA8iyH/9IVs3n6OjgaOOD86vRxCVIoCZWDUJejEAp3tgmLCABvip7f2cpxlUmyeqxFFBC
vfKYZFkChuYnBjWbe+Nj3DkRrWBrkjLzGTI2kwnENopiwY5RVQXZDTRZ5sCMyWPkvWimZ3jVl9/n
QCl/gaNzzrV85x2Sr38jTOB50IdrGY4F6w+5dMcZWC1I615cjxmCC/l7hLaMZnsf2Ne0LjJk2ILL
yt+ASFMBFBAIaG2jYRVsTUlg58lNy90AFiGbPdBSwWsObZj6B50XjV8GWaxyrtY2XHYyB24KZqvV
9SQEkrCDpkEn5uKR56jBK8tu5QgJsIcg8IXDgS3mGTAjlgxj+RDx4a2cM2CNm2P3zLp47k5qt01L
W31/s8GrEAgaqt8/0NNVtKnta83gk7sbng3DiKrAAVKHeBJCQ1RLxD636IZg1flR8NFHXhEhqF/+
94aF/e1ySm8roYbmZHEEJEhbneiGLEKSI7OGA+53o/cDCz+U33nDLUAb4ewg8JKTy5Gj5HIDRPaT
49G9cajMpU2SCwHq7u70YNCEBnakkNeBrG0FDr5ojPiarXKnahUcRPRM1T8CfMktDw1f/cgLCsHz
b8T9gLfvi3JdVQqWlUqTsUTsfuIMM4zUL+ueeg54Ac102nCH92e9sANBfHNrAtCoXzSPKBkigxC8
TL4XX0y4etVuoePJ658NUsD95j31yy9QofzCLOKMP7h/r5vV1FCnw0e1P/SMHbXAJNm4HO5LLsqY
zNL8qm/DXXj5vFY647IqmhZvFu1vijeo1w/QJ8wBSGghTMc5l+WycF04MH6cyIg+ODPTjqmyok13
ZmIdpP3onSbDh9RJlOXZ59IpSnAkcFjrPQcuD9UCYC+yAl1EA2uhCRVmctNrAgkKQH4RVIkudJm6
V+mlbCbBGyKr573xSi8kOsKgotb76tT56adB3wJbgUjjqT8CBcPpIrsyr6vAKJaHuj3Yuodx9ILt
23v7mwkam+GCnlH6g14nd+bxrTCQ5eiDbxMuTnOD54BGOHbRLtcf17tzzIhH5vGH4k7SjHxcyyEy
Y6Cp7KH2hAaMNKQdCIegd7beqJ3mYsTR0LpVXBDRzHDsr82aBVGgpRT8xo7+adX+/OgAjq6Ho+5G
vDPzJp5cOWfN1lJYhPiqAf3qNpDUT0dKrSHYAO0fLs+rlAQAg5ax6L8DRn6jgLuFFz2PCZnX+u+s
ZvfCw94rSv4lBmYSqPN/fo1l42R9XV6ENb+X4J6OeupmzcU0SDO/vgjdCAxuWbQIUjJHJ2K9Qbp0
kYNfQsgRaXraALIicXoia9bdMJid+lLmpYEHHTVrEJUp0HNgFyA7vc9wyNrxRTACw0oYZjd+BX13
If2Jeh/EHD70Q3dK/Q3EwQ+G2aZYQS33bQihkqUSOpCGfjzQLi1EoqYlLW9x8G9Gho74MjAfO6e8
MWpXlv3v90RYOlf1VgLqe2Vr5AlowWO8PXi6tBVunWPW/14KQKpXUHvf4VHwUswHqg66ih+WOllR
5KHo1fvhRh97shb9o7Yfj0LtBReQ/Af/rvOLLUOajggeRoQiyjtBOHM30b4CZAxLH0eQm1kLtUjA
A+n6xKMNo5iBMwOqEwRYsM7uFmkdfVDd/utWb/7fj7p3vYVSmne3hTnQcwvv7i3DTM39St/LAcRd
HY67lmPCk3qKVQA+ROe1h3OwZCJ0Q2sUyfX+ribR6ZJ6FmVlzCEX5IsJAYsz/UwN2EpFbqEMlucW
ZjQn7bwrpTWXItUhVTHSrphMOeYExI/cIgLItajHECBZtMegeQPn1Eqd7CaA/A7pcbPqgiUxuZMA
/KtVjch1YC5bskFS6ILS5HrygKJVYSpD8MFQ094I4g5ZTa4IHDaZ5x5ClgIYsM1X2PK07A59QqhR
Bavwq0RYTElvh0uzMN213oqk5StuGw4OGigMt4XM3So3cQNnla/L+gZdfYraXyb2dI2hbKIDBHfa
ySOLNw4OXkcL+zsNwmfNquNtQLoAJ+iXqS0rhVcXbz/u9JyGK4UXLpfxllY3rghlFNDmaEAKCzzX
a6YiN/XZEsVGYJn1NN6+nDJ3pmyQQzWs1/iM780Yy0Yxk2bMGMcQwhGSEj8UCR3SjCkIrH6Ceoqj
Zsw9rFQQtAChcEfg/ktKY0Jm2l39p6/OFvNPvtYo8LDWZn7Z2Qim7R44Tt6hglWTG3hZcPgr68pe
lMTic/bg59BFn0D5eCKu5Ipl1pFLY/ud+udwpiG//jkh4GBrq4hLGaMooAziMcSaeseq3KKiDZuq
4gzDiSlf1wWgrlFiP7GyfhUfjBSSghyNptI/D25CEzfplNsbKqdmgbEVop+KPEeMmYXJnW4+45lc
5x3LsPF7yOYaU3DgcezdQlZphXzYZEdb/YbZl+YzBfODalT5S05dQ6UuvQioDjbfZUCDps796+Gn
73IybvOur0Ic9WTglgicq/ydeg/CdcNXbo3/uli7Tl5OP3mE3Cd9O65XGXCmo+BY17AI6HhFqd8U
RG+RVlhZVjfnwzTawy8L9QA0rxIvkTZoBgrrCODGG+YOFFV3M9k9hOwji0AQahb5oRkXnX8cR717
6HytZo7WACo1yhyg/0wdR/3M7NeNEbFX55dZYxfiGKdj+YIbSAfOvsfy2BRHHYwz9PAjVTQcp3O6
XBTU6lYJUwDt6GJcoBzMQflrwaZ0uYpIe6LSMx1f9az0tITi18USt4igbEX0CD5Xha1pf++WAlWl
w9TCZIzF6VdEjmtw9wuiMfGe4kQpKYnGEt0YfgT2UxT13UVwuq9akToFy128hFo3jaD4U21x0O4u
nMrivlkpfJZ3VzTR25KWuMu7aDLUjm16pEYa3blEhKDkqQYvIaRzFiEUbZwlUaCkMQwe6s5GUCuI
wjcH+LjFfuWM+0ZiuTkNPojzTiJU4Tki2Ap/eHi/spZ1hruuIIiBAxtZ3+vMAzwGrXEI3vQlLnFW
THeWFMxbmUGI9a2TBNG4nF0VqZUL+79Hmihl7WjRoyJW2YyWv7oAu8uPaaGx+Gb92G5oRwZtnftg
iJg4a/28DdJ+k7NV3B7aMS1r9GzItvjssCgcTysd0p0nlqAcZZ6BSeyB2KyJExvW44127w7UkJFX
4ZmEpsU9jXODmULiKCwYnhfsgCO1p++Jx/n5BmkTlh0aE3+wV5bXbJI86RK6KfLg6LFxPi8irboU
UkwjA5u1L3a+DAQYer0NntAtkbScm4FhQk+RqWfOkbQWhVyUVOfXMI1GCmKFFIUlGAZ0cxs+Sbrk
Gepe56Z1wCL/9qqfBugkd128o2b5COjd6Bsg2KBLKCDwLBeX15qehJIyQZ7ppM1sh/nq72V9MZTt
I72RyciECIxyc6TItw3wCG2MHhrfXNhifrTMc3QsOwv6h/T50Bac1fuxKejqDZw4xEnEyvVdF7qf
Idq2zMy65OK2jLQUgccg1H2Qmr1p+e5DZOWoex2GtIppRB4DLEuvQMs0LBuHcRvd43mBC6JBuOMb
7IVIgS75Gwd/DUIM9sLrT1dfCnvNRFglFa7UTMtUJmxJ5CooSVb2A/QgKEWk3pOMNpkDTtsZ9eqj
X5+d5/Toe7wecf/J7hTl6uEr+8yZtLMdndP8HLIEqmUSR4T1E5OM1SW9NN4gPvscob4OdXSPBj4v
vyjLyOE7QH3BUvJ4OcCbMKG4gFR4H+cu5GAFD/nJeDOcCDTTPLS27I45LycHjk3NidBalJuUnDPH
jMPjI/NKfRGTNwMB13hYtWv336uoLh8zQwLIdVic/qdeFPwFqyhO5S7/sMLFjrbprQZAaNITArHo
YHDBP57uzLcJ4/0AKv4SvkGHRrVKidP/dPzl6aG2wvWorDXF2dc/MwpxAQkC8VbSS8xaFZv5Pn/L
+GpAVti3rp6keyge3n//95rds4Wm/q7xp9XbfXexrjjQ72rHB0lk8OzAbWsCng5Ds/sCTbmQIovh
W9irUatSbyfeIqGkRhPzc5UlNhfW6J4PqW3QZcyPr+umqyY6Tk4NoFBcUfqC3IosvN1nKxsgu3qn
JoG2oA+i87CvxfXGMTgtd3PWAihXtWXyYLQFI8BpAdLiJHVx/5rQ7rkTYvWwTM1UhYzScoSkLsPh
8qWDbLmlKKGTkJdQqzE3sJjZVQUvOQfhKnKT7tEnY15pXe9AoZjphe5YkKLiZRaRXEaBZfw0VqcF
/q2RYQ80W+vFVGes26cBvDglGG95ifvoLqUSvdCT0djgRHPiVwk2d/8azGKGNXm0j4rze93MGYbG
HcqLNQ+OsjiOyXLIuNQLq+wCK7FcPghTBJSgJ4bc79KwQauR+LrpSTxvzo0AtSQw9Rpl3wjfEHJ7
vYZBEgZ6yW7smPbje0NsanHZnEnYbAb+vit5M9Um1DLm0Mcwo+EylM/fMYesip/6eDN48VZHPawE
oUcA1ZbYiGFJ/ql27B9lmrnqannR+94KTfn2R6xJPW4YjAkYWMt2vG2DVC0dFSPKKcSlqV6UZN/a
RtmFlNI4Q31CSAgRpAlZacC2XjavRAhmaX8bQtojzysqD6hMfBOl8OUbODtjCt91Ia0hRczJI49c
FDNmYoN1k2Y41lAOsxgCYIT0iTGxuFUTO6eyzhpG176gwxL89vkSYb5y1S3oPLjosjPK5mvArrTx
K9ER+GC/Fdzp1dryQNuDJBLQPT6eMZD/uin/glvIqupjC84QNZcWgaSSqPzClCDaF199XDaTmES1
kEwtDDe2b08H1WVfnxBNMjPH+6BjvaUtf86wFws61gQD0BSoCSF/7tbzeWWgFGXrliW2YutzHwpB
ExkKW3HmBbPNDbGjpdc1TWpFH+7Twdx3JADzctH3+aspl6FwkTPPji+TxZlS7ia9DbPjPMNBzhau
F/FLubWAPeZzoZL3txYngyKpY4RIS/anV/yT05XN9HEb3PkhqyP2JYTZ+2puuoxuIhK/vaYSHAAj
foFboGPzPjETzu6RFpG/AA3oQ8a1o1owsLjOvZ7JqRCZrU3d3MdYVCWiBXVJICddcSYZNjcuLCIs
dQsCOrAChJQHKpxYuh7XfeVOrBRgNSVyjgsw1hMjEGFRUjvuOc6HVkClaI5xGfwWQdOu4ZGt9Dzy
iG7P+VIRRn6WYUxsiLsZ6tWg7ynu+I6sKVepb1GQNIgDJHtPXD71XO9Sa7hLZ89sIQ97jeXniEoj
dkmR22JyLgVdNSteWiYJRGGIaYTlRFkxRYE2/OdiUVtdQwD1qzIvIl3cZxx4uz78NzEuAKqCA9fS
xEkduxPObpgp3nfX8IAFuapZWEcQI+vnXLfOL0Kuib1yZNsxbGGGEl0YE3dgkyouGT4KnhCkuSHG
a0spsXyts9uTEU7B1cty7Riy/rNJ3td97I/epZNQYru2ZSVza/XlIOzJqm/1aj7wKcvMBpOmGqgS
sSmm8/7I8tBX6zGhhmg2tJAuy4nLyIFnjJOSx/KikNGa+U0tijU9EFR8gQvNb3y8CSUmRkDEytdh
hU9YCQWPVRzudjLpnv8VvK/kRKznmepJdh9GBW1zW0w0CsYbczoqjL40WQVcDqIz+7pJMSxpwWBF
4reJvvc7WrcOte8sDpXZYGClrF4S8O5ehdvQy99tj5aM6eK8PiTGTrUYMBNt/vbAPTs/ErE7M7VB
Ld3oGTiyy6U4+hxs5I2yVjtjqzMZzXYGPeeSWLefhANbkSgKM2K0JGhfybhIC6tWONvobBG0GA5Z
ai/PRx4E0RiRFPiRiiHZSC/5fa+TuXy/KtXN016M2uXpEcGkontEtUmZbcj6dPZghQ8hq8Df8O6s
YieGm8fbV3h5GfMun6qWg48Dbb33PYLje/CbxxXgro+tj30ZWNeva4M0tsLJXwHBYwUITZALhx3c
ncf9DyyMiyQZo5twMpQXV4Z6ZQJChLyIzVCK8ZN+nYxPQORTd9CExr4yTvv/BPeLaclsTHXWmRd0
gGuTKgYTJ/1vKVznqW2Skab8ASOb2YzsTseFqNkOI52eU7zoVpV91JsS2Br/RyXiZampJPo+TYRG
jtEmY09xprnbLCqoXrvAvXtmaalA7Uz0l0B6Pxs/AdSFJpiuAYmxNjWS5IbZ/IhlLKJB2nW0F5oq
4fqXlVBpFNnHuxYV0+tkN6KEZdovyobE02ehJW2XMZgpjdVA+d2/5BRFyhu27NYdee/Q5iz/nhFP
KGSszkPHYnrM9L2/WTgSwNsu6AdTK9eitKBQmuXTTgNVPykK2+fBGCsqLv77DATCW8cG3t5SXMGF
Baec8MyRKSyMaR5Hwz3jfPujybEllDsPLlu9BhDfY0r7e0jMxiv6ESrDBKFIA+mkPn5otHRtlbVS
4x7080LwR+tk9wC00WCVftvr7KKGmSMOtJ954COcocKMtxitcarLuy+aHeaY8nLq2R8LwNQYwVJ8
HUk0bdlRCR+0cHYOpMv0y/exOISLn73PbBZRi9Q187V+Rimk8/oCSut8uK76Ze067GFGh2EFkSyK
1eU35xQie00/IreRoXhVTph9OJW3vDHWQJt5vx+VESTruEQyIdzU1Wma4649ywvg/VMyWWrurPLj
LUmZSRJa7U5PdbSwr6sW+OJrE1saawa7OyNdO3VfIlHQiJva7+Xif5g4Oph9I1zPx6HYVSzOXGNu
LpcGuFQ90TkKVcz0pMdiI6K8H7K6iW1IBPNLvowd71V4fBpAz+bS3jKKMlplCVAP7M4rqZm9VJXj
S1kfxBU0/aGUOmdGNbnp/G86b0scTNlQxbRE1fCgAZWUVkDDs/iR7YJjkS0r3qsvuCXl4NdO/mTw
V6TxqWpOLtbgEqODQCPTLzt+mg66vJ6zYWebZBI4nqnuNE4Rg9LYQzlMGtq1w762ufN++J0d8i21
jkeRXYgUIN86Go9JADFIiGxG9iZwKpjU0mBqIMnR57nENLI8RQhZ1nspOHjyvEI2W58e9PEi8Onm
av1oK411GGsklRXH0kf4G5s+JQbMhEponiiG7++XIWjTDHTENTBUzy5u4cp8gVoFhPmlwyp7aOY8
stspXOSsVgxv8aUWr/XzRrOFxTL2TXSGcbPD60quJ48K/2ZoI08olXyHPJJ9zian7eTgiBqTvxHI
1Gqwao7Lu18ZigdCER882AKXDLh+FbOW72PwmgXgjuarGox1jVZhsywBl4ZcBbiWHrEhbGesiCqw
A/2y0jxoEj7Va+e4ib+cFOGxPoATx1HbPHkc1o+oAPhdAAOGh/SHtfvBY1365bIE4Mh+CINo+Rjt
70HFRr3LaUsWz0NkHDMura9C1dlTCN9o+XYDxlAjqqsHJLkN/bwveBtHQDXaTXoYkfFKMWmvp9Xz
rbQz+1yxbc5QMTzla8v80lGU8y5UfzB/YFY9cOcmkiAXGEYyXqTbWhF5t8eIklKs+dYrFrOjRxPZ
xgTHBv9pDmzyJWICYNy73xShDuyWBIpHglBRU+X5FL3gvw0It48cEqltPkOnWSelowysdPJCc9kq
70+SMhR4woonOKLhOzLJzMJ+yZSNUZPLKMWbEt3SJ+iP9Mc/o5Lh/eHfsYuIVLcGCVomxUKAP/1J
XRa/4XSNbJDW4knNFjjs7/WI9YxyKwfBuDbk/OF1tjcD9wTjC++8wcmxvQI8BvPKIciT1GpPbGfJ
yH5rOsCZpTFNlfcFsx2iCk0yO+NgGfYCq9mkpmtNAls5ZtKCvAdY4q16OknPLgyouLejvBAhQyKK
G3Se9ty8XwWUbbVE9x+pkNLio4iI55URdYequwA6FFpd3n3DF3/vyuzzFNhMDgOQojpcPAS2/u93
b3bSpAh+pBnbLxAcv9bWNv71IEhyRokQLRPgPXnsLrQE4bdIuke9UJq4zZSNw/ev0G5aHdyTPV5V
Gx8gw8avOuJGtV6xroguouNXXCWZckXtuvsKrnSid5ts8ZQ7Gy6LZds1wB+ZJt102G6YzUumzibx
Mb8HIHUIZ28jzYTMyxXrjzS8nnKxKIwmIck+6UaL6jcKMQbE8ZQGHKB2gAvllZDbQd10cN1DRoT8
bVVHHEmL/STv/x5r3T5muJOnzmIjLbnpggJ6V42NHIZ41CeyBnNuCUDzJL21Mvqct7QNc9WckkkT
DYNilpDC+PFzGOnQJeIKj6uSaLLWEBMpphvHtULq3ildsoJQKv19zarJE3lY6WrgsZTXhm94SKtN
a/aS8vV8HwTHHf1Mabk/Rjmukmlj3omd1S3FL4/byoAY98Qalvd/mP48LXxv7DD64XdhQD9hDsVK
j04UX+hGqEo8bUsqyITCHFhNz1r8pVVjHSSF6ikNEk9lZPCfB1Xb1ktaFez03Tq5bd0+Y55cn87O
82FwZ3krTz5yfKbdQ5OBZAaDdLo6wD3R68u55ESg7JlsqntmTpXgpbesmyD6UZlLyIjhhszr0yxj
EurUBTh0gNUREJJK/UWk0kUZqAbjc1LOiTAQGaTtfn6MYlaBK+uWRftyIauFxjlf7aW7ZXOk6fyw
OBltst9ivOAPcDamtVmXesH2Znn8/OEwGSeTNfXfl13FdRXPIqp8psinTe2JjdTLRswmOniC3JJ2
rsi0NuWp0QviggVmIvfsieUfR6Ltp4v6UBJWkc0sxBA9AXUr9Avg3KuV8/XB0ACKsYhfQVD0uYWa
L8oqWlGg7vT0vo8z0JSlCtDAuNiz00EDsLLr582Hn/t8gRb2adjutAZbaZalJ1NfO5EBsEcypMZR
kd4gV2UVNLptB32C5c8zywf7YLVeAnLTwy3CNajm125KSp/GeKPGmlCK8lcaKecZyOhwg88wRhr8
zC2BqF9qQhPHX9HvqxCxnN+Pop0gg13UoCtyY6UUcyaOop2yFUlB7z7qeVXZeCUluW/rOjB9z4/r
tmsd7H3Xoe74k3c+3rhUcZkRM48wsODc1VWHpt6bM+/bXyiXxwC7W83XxyByvKZOex4XoFRJI/3A
u9Ll/O/OBsi+tyK4fX7I8EAc5Iq82mAPTqWDUyWzCKLWKchyw7d8p2jyGl/RMyKoFiidZhzXkJDK
nu24/frrcsE1cSfONtGk86XvtxRXA6gI+AbLQId6q53WuDdlEO42SfSe8CWTO1kKpwpM1mNk7hr+
xZLFEmeutGxm5tbdX8PnKBcv8fp8Hbkk1b/xnZyMWa5KUZhfrTmhG8Lxb/tnYainATLnaeXXKUsD
5UTX/ft24Ct47bO7RNx58U1dqrDVWPIupuNcP6Rhed+4Zr4kXG4Zi9//D/mX5E4/6UzewzKntxV5
L9kQNad9dWYW8ayt9cZNlLDOMyraCPyjHu9L0/op4F6jJMd6GeqHuAmTGgNXjVHLUqDrHMQT1xQ9
r9wh/mRmIF6AO9IZ89hCcrLoNVgBxqmy5PTyPnvm6VQlpV8M2D3H+6/IJqQLEX8Ypz/Y/YqgXk3y
f0swY++Mc+HD2o/DDf8Wpppj3cpmpERY635CUZDJTgdOnaufUG595cF2haXlcj80PqJVlj78D7Q7
MTI4ZRgEiqaHwhCADc7nJLAjf5qUVDdvK5XLpWu8PWsNcdnpIkDySnVDL74k26ub3JfdtpsKdrM0
iwTQJyAgN0QSHYsYC3/IpwpXEH9M03ky+9SAzFT/LQwcOHHmXdM5JC2ErMI8qGDs5ZPbq6TXaTb3
AYE5myUbw+s63JyyWI8m3EbRSSSVR+XtB+jEb7KVvlcjbBgYXIgqUuqGyMv5DDNTGhcZLqj+zr23
s/btTKO0wdoM8l8Exq0wUDt+sF3nM7BFskTJ4aP/DMOaha8wBs1vj5O4TjyCk1kxclafRRvnzS1M
TMufSIKW+msObCt2rhrV9TLGxbCODAqq4adS1uLOTTM9NhzezqQDkgyLIs6L10puoQhc3g/9Y2R4
mBjpQjf9AbAgRubnKKFn1ny5Q5v7XvI+bHMIDzq2cPItrsKkTdc4nk3wRdsPCenkGbyTJlIYBrCh
ONb1hH0IPw11ETaVH42nNFHVula0FMoKU6SPajOuxmAb/21Sw7DSfGACwdSKVrHSkIkO+NDVcj8n
SXBQyX2mxpwuk5NfaSVi6oXOusC3Sn0vKtH0dwwKpOPuEMA9k1JInK8w9XoVm9UrqlcACWR5+L2H
0ADzsa+gWWYhEzEKKtbVVaRlC0/VDBew2b3WjqCPJM5ohLQvPMngOb+TPKxocDpnlZmLwlPe/Hn4
l7YLdlxJMB8IjyxChN3vju/+VYvxlCM8kLBhKqUsfSpFTGB33e5LVvV8kJbTcqU7FDJz1w38IuQL
KY9pW9KV2SxOxqHFS83Pf9E4NmHAz7MYJDo9CM2JY/aubK9dY/thF1yw0vsP4SXMfeHU06ir1ej+
jqnwXGlYI0WOe+q/XuwMzMgjbcl815Aby1vLqpq94h2Sx0fmoFF7uhui2+gOiftwNlw76yoe0BcO
HC6Tjww+k8UwIDTKmi2wfF4R6w85GxGAjKTzIPMP9/P9UNY8IiAXz4e/9nVU2SR/OhFDCLu1VIA4
vgrsOxz/7qUOwRAoEtf1ZLPQlaZKzYitceAwseaC44sJM/oxbOKgP5VCCK6Mp/YvyulftwhdJLNf
sRsYWwrW73jZzRWVWi0AQOSJEN/UQsYWpPmsqo3N+86KM6jTnhDX7n5ppdm7JQFqSSr/cRm1aEMi
2D6DSbwslP1AD9UoKMG11zqedLhc0pARiD2Gqw8MSF7bk7QnLMNNyVlrRU5amF6ZpLJYfXJ0OV8g
+zYYWwi5vxBNeH5LNJDvy/cqlEPm0VAY7Z191GWyVGsjFEfYkBS1tYWcRo0gemYmqLWHnRJsvsFM
vB758LaFzpGpvK1+fHIDFz4agft/JI+uXoDxAOLY1Eu31i+taoq0jw9gNG7vnFz+0fVxZ9263rSr
mMRKAKOsqlr+KcrGkqVe9yqOS5qyvYigLNhXjjm6R8pZpWI7kSHNs4oYRYDbqxvP4SEXh+D3EXR0
za1rR9MRJ1MMMpmsJ9ENIPiQUl8fmDzOj6H5KFmWykpz2+N4t4m0E32WMgnrHrHDRxFiSGGpn7J4
7qjFoArYI+sADcoaoWV7FllISxRxcDJK1TN+5kgWGEf4Ki7ZRB3iyOHcsgI23yKbPeE1pmF+bMF2
WCKqeRNqoLXPxylGqXZVDNuTrLCHaiMdyHHjZFvqljWC41TtOpn32YrppBghMG3SxWT8/xKU4S9A
HwNO8hTrj1IEfcmPC0jl+xYX3EZRdZQlDZa+WVx+ITUp5rs95yQD0eRADAHCsSCyl4JnzL81Qwgf
PbHuLLKdrAOAG0kVufAgdXDnljxqvcSOTR77a7YmApAl2JeHgFcwqaAmiFoSCrkoDrkZ8Tb1oy6p
UculuiMPWejWKCgdvM7g1wnIluSgi/rrcu4c2U0t7uW6Vfe0T58AuJze3EIZq4BvuYPzTcL2AdUr
RVdvQv2yTLdfl3iAbTZMHY8wdNHfOcxf5KKnuTQphN61qqFkSJbokxv2mqmjRvA3WBxWMHMPTzre
R1v1HcALmSwkBIenLTBUHKnlPxCWxdNKSR/yCVoiZTCi1wTApvE3qXqB30CWyAuepyXNf23uung8
rWgykqWdmGtOIu7ANyHUwC4AE/SsRrgcTHvAHpDtvn+2OgM9KmK2irSELrnWuzi4daZ/SsXwCyak
RaVZlse7n9qEYqBrLyTVh0IBg3RuCL44oLLyEdKvPJ5Y9WwncF9izfUf0jnsN8W/R8D2GitmPXvD
rl7uFENayVjlp5NLXAWCswFMqmjw4BnB3LM0xytC2tV8qBe7ho6pTaxc10qco/j+JotMl3TtxFrb
5R3Laiun/VOCWw7rQK//jciefGbA3yXmqKwob1PWMkVu1TYH3Q8WxzXgH51z/lZWE/LwwmAk4rAU
muYro9p3rDy1iPP5mKNncpwL9HPa2AJ3dW9jvRUcoNzythPqRhjoaSgmKQZmclt57E0G/3IZRCKB
skqrCPxZlbbdQfEk2gfJvpfzHQryPw1tkaxJGFaHT97YrHlu6QMtcnQg83pTrWTH68LUQ6WxUXNK
3L2fcr7uHlgyuVhpooW0a76Dh+ie0j7DkbEwHDoi8858wvQ2WFISj+joJzzkJnkJNvXQCQl7+8+v
nur6XVelVraG/1RmSojAZfJnnYHNww+NM63AmGX2zWsXL8AyADhtrohJBAmCs3zf38W0Y3tChvHM
xn4sVXuw9GHXMhiF15MTUUePH9vXmtt2YfQ/Y9sRptLqsdI5zeNgdn/D9WCvDKsX6x1CfFJFRy7w
9WK5GRivXJxuyeVxEPYlhAyFjcQ44Em3Q1hEi5Eg5/z3J2r6TMp+wFSHO9UMCTp5+tWdfnDCpCo9
kpIVFUMiLKe3k0tepR+mslu6WoVRq2ts74/6vOLM3VrOj0m0G1tP+RrsVKK7oifdnCezTJiFj1Fs
dl11zYiuHePHCg5LbcibHUaZ51ntEy4yxT4Tc83yDt4zeSVyoUMx0tIXCt8pmHYxqcaTL2BGwn1i
cngK7HXQddfsEkYRBpII6+1fSe1UlpSEpXStY1VpEkn67O2EiqRdubjklQFY5s5D2tz0n9bEq+dt
VnyaQORKUIXguRtRTghtZbwx6AQ9ZoeXyWJvzwzwx1qpsLYra4PGXHPpW6JUbXC4sN29r5D0i5va
GG29/Sncy4O605MdwmqbdL4SIbEV2EVN872D+zVRwG6RKwxcoBsQFV2sHZzfoQAMbqvQ6GAyC5FY
f3xH0Yw50+Yu4QASRrGqJyd3h3DAihj0u9EfSrNVHFBfCj44fqMMLbgoOBfyFVYlzejtdwsLPi+s
6BuUUifdW9QWMNAjLAnRj7UGiAAGTyVfCmQstlXFEbz79wHUoNX83zgJBic+KzyHQmhURe7XLP1x
6e5/SJPDgtLmqXpQ4PUSxHI9WJWroD4+ZPgWKniSoGM4R+30fMTof0TuB+lC3D5iUPUVC2WFnZQv
3GF+eAPjCGAwdhEACCdUCiRWjYOKCqgEo9lHaRMOsUmCsKqjTlrVFIJf6KTxufZl+C1Iv3wtdKo/
uE1xlFSTnM/9umQpfug1nH8l6eFMD4BalIQGe26ninlNqtTA7YmS3O0DqEtrG7MY8YMJcNU8UuW5
fSc3eXiu1ZEjXXouv8dmKj7PWV1JwVfgHfbR7sRwOWOccP7/2Y2My1MLyZ95TTot+aGppwprOLrl
NK3P2K39PmAzWtBSi1kiUNlDnTtirs18LD4rV4g762sL0Y2ILVL8Waa9tvnizo22l2z5Nzw6dDYH
Z4OkgRdnajDG8QN7c0QtYD0KpYf0SyvnsJhW2vArvRxd5uoSAHDWvW1BDJwi3mXyNkPL7i4N/qO0
jzTcpbC6LHoRIbPGsHDPi8hLh2tEa5v+oz4GuNf3Def7ZsdNyduZED7GZRqE1hgyxYAiAUc2mevO
tI7Jccv60giG4M9wMxnuLcHDcDMbxgO8y2bIiPkwFj4NTPVQflXtnt7UsNO7eG2AaBhMqMM6rd02
W+2vLrg2+2c2hSMTBKoRQavKLvrWYS6W9MmD1msqHwxePrv4qvfhklqhXuuDn6k/eMH2ICFZuu5O
/ASQFI/j1yro32js+66iYm4z2DA1wGhKLL+Vl38H3C92rrJZawZ/iFxiF978Eg2BkjqN0USwPbBX
2W5w5cUSrfj/xCbIHjUe5H1t+XNQATYt7xOTU/LWiSU577YhdYuElovzTKnBPfwZqcLAMkMc8BmD
OiTEVPeb2CXf9fMHrHGHrIu8vXoSJ8hZt43l6r31CNhXExKvYItfQ0KteBW4jA9Kd2rnc6xF6bxE
lawIXD1vZL6MDTbACNGNuGKdkJiX2lB2BgqvZe66zXQLt1ifPsEn4NmTEj5WUwqpzFGOkVu2u169
yXYmcUAvZWSwXlmIsyyvzQDRlSS/2vYsCETPJf4g2dGAM1I6iYLaAQGIwQVUWbJTIZahh6Gh67BQ
i5LHDfW+BoXu2ZQnt3ZGs3/9CfhWrtkX+mZSjHfPurVhaa4afrgT91xJf7aWl/IYm8GcF7ypzyvf
8DImtQ2a+xFUZbmyhMvFXzFtTyQfgT3SVNHWHlowKYUJ5eRhUlgfsaga0ajyswiRHWMq0ckjnq3R
6I0BnLjoteENJr8iGrMzNRZ7eVbTC/C3UNj+W4HhWS3HZjv8MiAKg2T81E6j//Z4uxjmOILu8dcL
vmPvkBzoe6MZp5Otxen9Z4cqaq+eLBGFi8s/t2pWmCIXrzdirCkuPeRdpNJdDAhNnLwIcZCfAHGW
52w2coSQBpuLkG0fiM6X0AUCUFCArSfhS6gDfIFmRbi617bEzfhKFasx9gg31ikwB9jRq0wKJhGQ
bcCkgAfuIYsB3qrYoILRe2QLO0+/utG0RGU/h1nDxJ9DvEOSW5XWDiBO+Lhk/g5syS6llaTIBbXc
EUPFWqNgolABKGZRU6XuPvAEitKf+xTT5/mXs6HL85hRkpEdfljmCR0tJcug73PZ9wNDU+EfVYLq
eXPiPuIKvNvIwAc/zknRTfq01WKNlDXA5Ekn4N4ln3beU2tegwAQceX1aMdUP6a+3kE2u9kZLz/J
wH3oG5/a58W29hfVq+JEyIrQP4tvBebFuw30bP3X0TdcF6bmwixXJrn8dVPU9mKXZ8ugJr8VeGp4
TVZfnglSa0/Gfu6MT3vIl9PRHHPRP+C81YS32zN4S2U/BHAY8XAqVLbWIQ2V9uKZA+fwn9kTb6k3
tnexwpd3D1P7VzQWrwa2vzuji0t56mo9oRRJ3MXeux5xByvYHqhGyJ/GYy2KLGHfgJTSGuSfIud0
pkIDHg7xpSsxFKXt8Dwi7rY25UFrWVaQllR8IWCuqUS6pjzsGoxYXTF4CWj8NEbBENePBPETM13H
xWDpNtHlyvdI6N4rDz7RTMt8n1wHG5SRd2TDfHEHG6PAqZ/sYPwo+6y1v0jwizQolWFX0RYQ9NUT
p1TiWEp1LVhAiyydqEkieYJCc0bPXvLeNqfkSWe1sXNM/Q9oyz/SE3bNqyiEE/XjoxVqbPE1Sq6R
FyiBMo1UlWRYnv7+vcxPaYD0eYjOKO3FvRMsjO7Sj1p1giaU5z9STs+JuLHMGaklw4teJxTPoqKT
cTxeiQWsxa/6fAGlQStIcWqNJ8k/DRgOBNXnFedzeyDiorE1Nw0hbS2drnZqOgpKElonRDts6yun
7pS9txXMd9ngdEQ/RiUXOs3TOWuMZBzJjbs821u6mv/h941soQucp3FhB8cSbNuFFxpMz0tU7hsw
POZ8ohIuCpb2ytkiuhvGMOzgWNMakcjkhGbT8HVPQRKa12T04lRguNFjGM2N3CxmRLTOCkmcu9cP
3PwzKyU9vHUYxpta7KANZizF8MUXtvaBZ+yS8fkyvvtbqo4arEQbDHqFMmmO8H3xac7DgOizzQOH
G7B7EYSe4lajOGlqrkC6Y0gnqwd4Ll+zqs3QbJ91MOpiem5cSxWXHUh/SjJgCwuObAsMUttxpzso
7/0pz+10DnXTQRqa18nzdghWwd/F8Er/FUJ7U36TgkJ5MsNJRkveqVoAHOZrvedoNiOuBELDp+6A
LETszWN5Sw/lORfKIfdcl9eG4FnLMnNmS/d1wMEaRw/FrccKugIPhE3vbvN0AHb/NMdceE0AeIjg
0ZPEyM9RqH1GUjDdGXcX7MyQBT96YUfuLciH7YoeWSd20RN8kryjawFXVvLcXR4+BUYD987GKS0i
Jv+X7Ns4tVVVNq+x5gv8cCCBXYMOvcfwokObdBZveH5HLMXOOxQlP0ellPG4xwiosNg8oP5oFDn6
GNFUi3At/k3/cq1P7YSbc6qcw7gq8NcPL65gtTlcFCkYN/OBTNQ6K5ptiSqkD6JqY52pTi0HSvAx
Ru/78o2Af+1SnO9EVBHav3Try0HSf5j49EvydggXIeQ/mlHrPkgEkwijIYOV5vlCaLl7rVRVFR2F
d8qXyv3IsSijmnD+4TkLc9nXTJJ+lAL0ZSDe5KHByQvj0sGiaQ25UPtHXRRquvMACPF2J2KVp6oY
QJHH8USPSAbb9v4RFyKtHHJqpZ2XEY47bGorZTX8WSremTlx9sHzgOa4OSiZxYJ92/JwjI9q/jT6
Osi8cK8gUOy9YE3dS2JuafQ9C5N1JMjBFGSnTihI0yl4FrYlPLbwWZbgg/Vbhu62fmEALlhhSWev
74E21RwTIIGIl4tw3ddSm1Akni9MxVGCb4EkoH433necoJoQTRM3LgiALHTeT3KvBvFhIKDeaER9
Zu4JMxj37GH4f4Q1Ta43TpWpa0l+TLX+YTQGleEMYaFQHNC5+brxvERaBHIgOgw4gzFQlK9vS+24
sxrsGFC0PsaTcKzIF1T9uTmuXjnZsnxZtaLs5z7Kfr6sfvzQ963fDk5cTP3rlqV3S/2b8jpZJOws
NlYQLR6oupdEOKHUxD2hGCcwYE75brJy0aRNy8EgdtqLtVxYQ/2l343smj48WcaoknT+v9R9fMCf
XttCPjQ9pmybDIDXiHegFTrfDWGG/YI+nSUxhmhqQP16aBF8lcB85xQcwlOzqS2WlkryPHyi3v16
/c6qA51yGMS3DDu2wGlT+3er7kmUc96MZQR1IGDRRRt44C95i6nIPM5CcTCrQlQ0TE4Qds30j5LH
jP6IZ6woru+8NHuJgqJ1l0Jw4lKtP/Hd32FZqJ8MnFnQH8P5ZYcgN8vyaiLHUv8vzFPKSLGSCRKP
vULRbQV9MkFEMTuvRNDK/TuoMTjMjy3Flh+sLmcV2Oh3o8ZJrKylod1VdWyMxevhwG9roVzZYUoC
o1gNdu1fWXbw7pbdgl3Eh6Fjb3QAORMWlVHXkMBDv8nOlU23ZpScFWlczeBaM60DeT3fVCNOCBmJ
dxssqUuBC36VQc/5UhCcEIwo5slUAT+fKXYGoN+mOt/6ls/fZNG9JebPh6yIndEDxv7HwR8qDgwc
NfAfdO1V+z1gGM1/ZBDOTaEsZ+jVezFpsfgSj3kI73KYrREfmZ1V20dUmi/96r3h4YqX0ZDxz2xQ
bAqStvaCLiKwANpzJ9I8fINtev1abIMFbVS5pAJI2qctR3e/3E9ip9TI6zD/4zuRTqxCfcjpDdFE
cHPyBBn/7ecZiPgtzJpXVNoPJgOxQ+My8sqs/5Nql3bjjqF0fxGe0tZO9mFbNxgG1legrYAj182u
DINPcK5BbaO/38MaFDpwGEsPtrJcfMFo/Kh8R8fFmtg6e2MXXWId2+rIRp3gPgTBnDU8OGi5iXzW
+dNpXct3oqfvSUL5rtmek0ySYXYYQYAD0z8Hv45zMttyWWs8mRTOzG/3NBbM074u0w2IsG/RhnVz
/rXCVAsYZdWMCGPjVSeR8ybD3s9JVMbrBYgOg2nTwrX90Ax9OcwxjgPtfvp4SycSliZHcUnjk35X
VLl39HHNsaq7dO6LZ3QVYTr5XNNwCcKI6v2RtlJmkThdsUItPzS5NYd2fsGa9gn7sK6SogTtF78n
iC1m6Sm++1zlaBuend99A/RawPVRUdgMtvDmwHLyjiivTuU8XtzP52JW9tO1xUITZswBkCKIN6kz
wEoEVRNJmaDR0MglNMPtrynDv88pH7XRE3mg/aJ+tqwzMM6Iq+br5OZsYHRNwyP4Gw9iJX/tr4g4
gvc2uVZ4Ty5Bt/sSYve2a+f5UQBD5TjzPctcvE5LRoaFlFdOjei1zZFoRxifoLd6edKpQcGzhbh8
Qi7ED8kKLfRL7QZ2VTz2N5jyd7r1j7gZ5ZeZQoKziQQRPeFcgOy40DnrwdKeaLwLx9OFTX+F9QVj
jAL8SUspnH8ssTEHhjDwBTckD6E+thDNLVuW8CH3PnaPigg1ufbZpljPJF1EoxN3dUaHvkEFLIDc
oh9wIVMdze6topTlD6puQhFKw0KaJ3lbBUgHpEdHV7Kdcl6MjxtW2rStnZTVAtVSUx8oM4t6hXid
pGpFxxuTrYmjV8dHZNHU+jOrVUleG6BPHkWvRKoJuLoZG6kDp0MNLWX4t0MizoFFaoCq1MqK4CoY
9zKey7bfj5naf8NLU/40iI0RoefszFhhR9mByN7Eel9zLCZB4+X+gHrURczsegsgBhb3bmJuP7dJ
l2jkIAk/7T6JpiqLnbUuPwn39Y6jYhsNYqiGr/HHSIGvGpD231tsyM0+kckrn6N9wQvDOR7pfqzJ
y6k/vrUhu9WFMJTH6n/69KC+Xjg8DieV5ARxTbHfPaYoN1msgmNYETIbHp0x22cd+gzugcO2yyuX
jTVUHc/rgL9fVe0eWIOjacvHm39MITi/avlcyHtx+uBQDGRFYjmNewyNAQbKgGQFV0hF7R3rb9WO
VI/L/uHcMAkP+rt3q1nMrX2xantDe9gI1/8e25/etoCQlO5Uj8hUQ+IGDMuRZMxu5nsIvvFJKcjk
pJ7zVQawBN8iiAVg1yxlj10DlbBHj31hpjIVrhVRyP5MWPkq/ETRPX6T1pgPRjr0NYNd0cOkdXZh
6OyDquCPVFTvYcSKRX9Dcin9EbdgEFSSHjaO/2i+ZH6hxxHjg9oLEEZqTKDmxuq4ldHVJ9JvnOlz
b1OOwmkergtG/C1M514x4QGzq5KEUqmRX8msTOSYdd6IgspnRq3MuiqxmojeyNYywScK8JL84zW7
6YDUTwXjBaSUl1vkFgelIecyOMmIMAuCkFRu4tZimey8AaK+kflAuX2vEXzolqUjkOWB75/9uiTF
+pID52utUFQWso4KQJhsnTqTHbkFI9hdzOsBDhWHBTcHVUkHLkLFOfX/IGOqmu75OlWksN/w1EAy
apC9J6GtyFw+up/xnWC/bzCF2mbPrXbnzyJkSeKHlD9O25zo7srjhQH3fUdO1CB/RL6hzTQAFAlR
ds7c1++U9bEMs4YsmuVT0IsSjD7dd/dIHS0YfbWc9lk9ivgL1bJy7PPWugatrKR39hdku/IV8geD
n6ZoxjIuEp/yq+TzKIoJFD78HjoYdn6mdav12sW7Z8HQCWr2O6/0ii1ZGK8J1kYaRUUZl0YRm6xf
60QLUTOK04IvpweIBYbTlho8TQE8HdUbOjglZ1njAiNuIvvmMPXIcvV2cWY2ph47oL89wG5thGx2
kbLSD6MHY8512yEXIyaLYBvpzhTGI0mqYkkWUqWjF420wGB3AuzKFKOSDDFhdsKu3ybUZ4XFS8E4
0zPNlk1zsHqVl41hSEj0S+JyQLrglI9fgdM1s1/82kzzhhCIR4HVj9H5ENeu3ODT5YaI8+91/yk9
zMIKeXfz1k97y5cbampRMpWLrktpkYgHIo0ojoIO7oqTGw2KU/uv4fAY4Om3ePZbj2nHg2OX4fsx
H8ppEw8y+Kcfh/oMtfOlhltvtriyN9NrBhhY4FjxnjCagxtzJy6DRJMU5v8KOXFUnRPoKUKhhzoA
rZLJdgk22jSSnoYb9GEIpFn0+wlmY2VWdpt4l0ZbmTrJNYP391C+60dNEURo6ALdNCbvDixCLePr
YB9KtuwQtIkZj88w2bv73U4YwfD+4GV3m7H+ym+ZSg5Intkw+mMdCXVz+kvqWajnrfMN6PUBp+rk
DKpIUTLioLS0CyT3DqfTrTAMnk5/ylRxq6ajdUiEwkaA6IMyJD9ueUA+74V5Vtk6fTSiCL6DHbuc
gct5oQzv11Zi++T6XOsQ/zUI+waPYcmQbo8QY6lZU+fCUoexvqkiHxwEiSf5MIl9P2jXj2dkEPY9
BkVFAHhphEXo7gMdLjaPwD+M7B7qe1F8xIKTmrvN5LKykHFimKzuMXD3g2Rd1iNUkr9ByviQYDz+
p8qS2h8I9zARP1BBD94qqDiIw/U57joU2oRBYRuTpAjbGppGgbjkNAuZsi1dAm7Wkq1fgPKPuTe1
zHpRt+zpHt+7TdiYNczmVUPjW7hOG48CQ4mZYBnqRpo/HTbT76DE6PSaCp9nZm1nK5cVRZ3/2UbC
y9hd5C/r6gzMuox4LPq+0iMdzluGEyWkCuX7/KosR7PDAslOLz/uwHtZ2FYwOzGCrJBalq1xPtMi
urwaknKBavSoA4/uToaFAoPnqfcrWzGeZ5VVEqqfTSkAm2tLY+qVQlpY/QNDuf/NwsMOGi1DHFYt
cEEav3kAc+KVQSETgmeaw1Q6WUP3o50FCDwEKcYL8Wcaaafe5Ed3pJ/K8+bI7ZWCrofxXl2aDVVB
8F6nmK+Jv7H6KvsZlXhrsw0zzna5HMX979GnKB4lXApnrWN10i6vUrekhRr/jfDy7McJ8yjJ3iwG
cPjfeia/mjp40UhmcFt+XTIZqJ9pLshUZAF0oCTepoAUhELSWf1PKd6N6zEzgCN2pRALfz2diH9K
S1PVfQHsIliYrAhAh+gXxJFlDercPNQHLqodBoh3evIfEFcN+n8luGInACc7uFvlCPK+wpGfFQbW
o0Ih+0gAn9BIWesieJcy8Wm6yubs4QtvpzzyX4dy1zAqllnjk7GvU9AWpM/MMGfO6wXihktXysHX
O1+1Odi3CFJL+FBvLu52JV9cQ542tlEWW5srxSr76ozrrXRb6TH58uW5iR09QcKzy4sx1fTz4CCX
X5NIdn1W3rdiLFLfXtbkrsQBdDaGsxKyuf9zaOoW3mA62M2J5px9NIGuiUDOJpyOi/IDeo2to3NU
tLLoKzDIcHnQRa+n0ctA78Lhps1mAfJFixSwBJMgi/1Wn+JqN5mJIRVw7F009wNx7Im798gFptpt
OJfEa64dutP3zPIeaeIyUeRBieKZGjKsdd3YpuY1ZwAvGlgiKX13zRG2AGhHqoLDu0MHi6RWS8Mj
lQNlOolk8iAwDQXqHoTptH61Pk1jlsQ/uMBxHzl41R/PkK3P/9ZlGN/QYq9ETNKesQe6aMv/4oIb
+JEhBp5ukO9BrTIF9F097uPSxkOugtzfO9ocUoTxW9I6b0R2/h1/oHe7yRp84c1K1dV92t/kX0lz
g8qMuxwCEt/S8TanDE84ryxahjmm1mnNZGm8Alk2BjTuFrHfwkZNn5LYNpLURdYXaBHyQvXj/ENt
6g0zO9ekVfMjmTQ3oc3QTgQzCFHmZi+/oHYe90isN3PY8KsyuVIPXn7XgWTkIKwxqZtXK753HW34
eL18NNTINlv1HkVeR+jvH9bTeeW025RfoHZkJW5tDf9hCRAYc9EFREY78qHMiKiXZ4Kp6vjsuS3O
U5TF5b3++48W/tcpiIIlBN4xqawCDdD21IyN8tdscq1RczQHqxHihjuYlsRNdF/R3DhkrCodUgeq
bZjAZ13GqcF/Yn1VsoQVZglpxJ+A3J3GMZRhxZCuf4ApHf3FqE023MTvBD+yfXPkUZL/CCZNRDj4
VjHwFOdyYCsOEn72IiJul7NXNQAMtbHG1kPzbuj4XsuNiVCN3b2Ty561XV5Mv7qfnpbppcnrb/OP
xKWQXYSYZSsvX/1bLZJcSX2rr5rMayxdNchXvoyIKnM7MNg9/w1nZHNpP5N3Bptz7/rmJl6KyS+P
diTr7O4KTgt1dicadWg/3mRL2NnIsazwygC0CggrlP0skJ7nBOArf/VHL20rg1a0MP9z9FIS/Cy1
h2J9lk9v3lPu/Pox8N2wtDOjo5dOsleKeCtQkNpfizHoWgw2vnVZw25xAe4skyef8LOjm9LiYsKZ
9IcMOXY5FX87Fm4l1NhiTIuF0hGwO0pQ1BOBSZC9cxrDXbdVxWxKolq5MsAclE2g4QY9rVMwKbCq
zSOiAs6iNv0df33ioIP07mNiWh5PJsRyQ5HwMxtY6nu6tFrMG5ElRSvEVYzET1dBj0fAiTW8utmI
YFRl0Hifw+HyCGNMAJoTv0+SkFX3kPNuEKCddsAY2q2YNnXg4gk8yMgD5GRxJjEt5KP1Wp3oWoNh
WozF6Q+kVoIr0yHcVCm8AfJggJ8E3Q5Y7SozrmYtwbMN7zKygXeMpxWvg+PeJphrCfwTdJZFva80
BMIh5xYrc2BdAk0p9Kgg9tMizTjuFEg2XVx7eUvIToVPaR6OVNo01wm589Y7cGd+HFjAkCgtp2DM
neqYmIh1rjbKiR5mDRzY/7wZogrj4i5E9SZ+1Zyv28BkHiDbpmK0m1cAE5RYHDKWEjvO6xK0F+6d
cEvm71jjtQX8INmx+sSlmZmfT0njJEU/8jgCv5kMJFi0qPMfIfZb7UlxnU0K87x1z0QAyYjL5w+W
EuoYHM38nx5W5Jz58OVigRm+NB5ZoPtubpbkl55G7nX7bAQ9Xfkr+7QZAJ8aWjRd8IUK62JBMiCW
UQuoyydiB2A/pDTIsjL8j90eCw3MGxoclDTeyvlForXo8QtuGn9/rml2O47VvmzwJQprRLpyyESP
qCLPsLl2pE0ocinth34+jZSVCmgzMunJ8j6uZ3kt0+SjNpF5rg0K5qIrYJ3Cu/BEGRk6hRsYWnOi
+eD+Dur0iDe5QPljiD2BcGnOEFXJHROrvioIdlztw5EoI76pXLGO2yCuXPnrX7APAlYrsUpO+ahI
ducl91Ieb38rSVfBWY/X6LrdhM2iBgKZiccyp2HV9xpPPmbHvVETyWA3sBJFvs0HOcv2pTtPDPGn
Jha1j5rnLIXfegnCzjKhDex6WPY8xfRpAGLUi3zZ62w+JAPD1T2GErm/y/fTRd4QJqQAvCE1bvNX
00WwbmRVB59MuH1qowsB2hCFPzYeErYfz6HDTKYN8Ujv/Ysj2wJh6ud7CKHHpEwaTLbXX3cas3Wa
ACp5OK/4O5CfoCGrURNfYG3MQaur9Tix0J9JskfTroxQ8hHLBDZJPv+Hxsm8lVuK5aOi1/nkrRwL
2POlDA5kJ0+w2asmiSG+30L2EPdxc4Kjj7Hdpcp0tDvEi+vjsSpfKoTYbu4zHtu9VRV9kDqIrs/z
1upzauxyxtRK39rkmMDLFZNxzDeG4TnNJTzSrJZXwafa5VQQQiFjNJkVUCAs2FuMAkN9UquC61O/
RseBxMT6jmeY5JW2RCot9GkkmcJ88ElckY+2pMxn/b+vfGd7pGGy2OXKY/UIvpgHlhbnaSzGcq08
WezAbIyN/eICPZuzX06VEZlh5OavH4p5+QMV4bdPAb2zfvETeouNGKLd7rEqK7EVrGJ3YGEzLvsb
kcaRRAQy2sEYr3ijTcjYpXx7rJU0xBBOkRRHZ44B1wLIUaIZ0Vjs1RaWcmBGfmy0Y46/DX0wbJ4d
tauP8WJqfOlSx8ds7lT4AEgQm5Im1hx3n3bV0Dy+f4UscaTiwB8f9QHUqFF6j3e2PlTDHpnH7WOE
uasv12OTvz0ttY29oXXRVFWWp3GcB2KD3yP6xd9fbcKv6oY7dUPaYfnxrble4MM7o/bVl5JH/YmA
nSpWbLnR46znsdZQVrB5pD0vl7BM/yJ/NGZQ0+OY1JYR+6j4gPchv+x7RsUIyKOoLKGL57t0B4/i
T6oJLP7gCT9KC8EIZQgwpZ7cP+CIgUdi7Fh2IxnNzrvmUKwUIasaGLvKwXKWDePXe8Ukmdl9dufj
PIpKdcPGN2AvXAuS3uIvMTDOeK0nozZZa0lYKGOfly8Mg/7f8Kh8YJ9GlfcdAQx/A4gDoE1TfZUI
Tj47bMn/RWQnq2swC4zpZXbAAy+idEENhpDKMyIkhKUDAWPMweLnkyWtxrm0DPGNlKvNTENtfzt6
d8LuMSdJGJyk6wFKzfIdrdawaTEMTquhX2nq/kjGlZaCVvUbKNHnJN0qGGbASFRP1TUydV3bqZGm
rxirMc0QeGsOotsbPPLfNQ+OzoPLMk+8f54JzHc0NIvJjO+Qic2Xw99gCXkM5KKrO0DFQJACVyDi
0Br1TkjkrToqZBhB4ZkoAtI5oZpGF8bHOR+KukQgLbxEKAgdvS8tyzH+EEAsdQlD0C6aglPWBULE
8w2YZkIaXWJ+Jx3LcnLfqQyTsQTL98lHTKN0O1BSHzhbvSCQQdPkTjAiXtR3c8KphBL8M24Gn2MF
HDgVFMIKk8NlJLkP9CFu68TzIpE2mGg0XdfiDihDVlfH3XxDQCpNEFI7Y/GkjSG5RSJLLSuTYidG
8W9ZsWFji0CjA9Rw9B49l3w43hlL3wpICKkV/D0kIEeojtzTLEKKcDq3oO79pBUkPkCHtbVRY/O6
rFeQSVjvC8jNvnY0psMc33qxuOfj98EiGsjvnenJ47aGzB+mtC4nknhNS/d1QrlcDBpPJ0931+F7
8QoYxHFXn7U7LoCpiLBRprum+UKLVn1bCtVV9EdQIxJhruAjFNi5joXiSgWc+BIdizV4bJYscpQR
qzy9vbD46HFltEYmCZdu5FL9jJ97m8Cr1oi3M0tDdNh37mkrBadJ1lniM6BsYrZb0UmQr5FAZtVC
qD1eCBcA6ul0677jcrpR8dBDKJ2w6jK2L1IjOYv6fAoBuDtjc1/XUxGTjfAtR/I/9ZNY8hKl2aYt
tJRQ1/JX4VmlsLR1ZMcdXRC4WPZ/eZ8uTDPqd/AwKTSynQozIwnH005sIN+ikb+L7pmxA8k6DGH8
cpKlmCbWdK+BdVEII9qUFUjca4YWYJa+ES6UhMDgOd+aZb0dhlhyPaGTbBYuszrozFxxfbDT9r48
e6/rppMFYqTU5xsRmMRDPbD8rPPnTvJVG1B1+o7PD+ABI26dMlmjXk3aVA/Qewd5KH5AiO5rpjut
arPfLBpkCX4JPfMd0u+LK0pFQXZPYU4c409MKHv5e95sGB0S83kaN6nOu/AwP94QVv98csk5smz6
v4nqk4cW1iRideiJ/9lQQaLT4wF/UXfLvoAD2JJU0BO+e4mhXP4AXrtL8lsJ5yMFqoCQwZx3WzTv
6LOy+aDR7zZBvhuXV5IRKXcWjsohg5WmQHyBYUUJFREx/JUN63Fc8GneHitNXjTNhQk/EXge6olL
hMIXGWjyD+2O3vq1qxRM4dpbkXY0Qd6U3Rr81DiGYd7mM5ydy+txrLkJSExCM/FaGgu0QdnC8sF1
qITyNJSoUQPDQFe2ablMJAa2ITFqT9ybdf0PLiqOVIWc+ndCnsSQKtPfVLJS3V9mYSCLZePapZ/4
WhPz0nF/pXTCckx/VTsMZ/gzIQz/BN/ORxdyq7uecDuHDMRBoWygYWjU95AKNyUj0CGIP3vjTl0Z
zOvIARAohQre27Kxrw0TDz0AIF/aAsHNBXTtkzB0bIGt5L693sy1SO2KwoBq07TUnbSm14yn0ndG
HEZoDaSVqd1wUqsgBFWpMwW0/KuMM2Bnwhu9jGSNcGBdMVvJlYYW4+XLNCXyzRR4kN6TGMTKCRT2
JdXtwZGiblBj+sOSlBR4Ij2UUxAIUSNmq3q/Rr6+u0JPwM63blFvmLTPhKMT6/YP8gZBu3EO4OLC
R4H0/uQe4bTaXoGfVdkvpEbBr1HVuvgP2CDz7H6dRTHKIeal6zJlKoxpakqqQoYdJ3haftYb7Tt3
J2HhYUc2NZ3OhlbF+iwGBlVWlfK1iJUqRiFSryRQG7g+PmdZeGU08h8nRj0B61UXUBEO9JnXxf7W
3/YLZ4KKlVHQ+Hlfele+AsmlNhOeR5Y8n3ipkoJgz6vC664O4F3kbWN8Mr2UKPAost2M+ksS0oSW
s4WFR2WnCdjbvaIVwF7IQBbRX7hrqzQZ26eDun5Xb5iDHqy/vqj/Iineo0mhQG04MkwEcxHnUxMl
RnQ22S5UmNgklQBhm3/Bmlf7J5zeqHXei0pzx3CMvrUbw/tESmmgsiqhXbf6nulNpIA3V3z+2aKW
4DVcrvt4SivVBFLCKN9n+gldtAFGT5K0N5uIaCqgVaA1kPMh9PGLFPVKLcaqcWgYDOOHXvp7H1j+
DfbTafjMNNbkVR7d7+6PBf6zqoRu9YVmkX9pAkTg6BtCB3cFb5v2c6bI8vAfOqgtD2ay7pj/M5TC
bEJ0mHevdzyn9lXiKs5VPukOXGKOyElk+vAdi5cKvCIXOlcvt9fH+0eH4UbK3oJ8nyfNgNl7asAu
mCahWdEqfh/OTxJgNeCINtaVNDo0KBLEspxjb56r0nZjd4N7yMEFPsj9bXFuorHc32jvD9U9YWcI
4rEb1gyWQxTHZuhQr+lYbbS7X9H55iv2D1qRXJa0IMu5UBsokIra02m/DYyh2eLzCRXDyeep0ewU
kuxYAuVTWX8BYFC5aqKfKOqKcMXnn9XElTQAvB2jTBM6/30Tu91CRQQteGZ/r6red+83LJrP6Ybp
ljSmspnefMKWcS5cXxXj0IzJtdo9MUbFNf/dcM5gpn/FdHiiJeKuHSdhJSVA4Hq8ghpL6SO+c0ox
k9LZ9h2KdM7p3S3WcQ/4BFP0yotjTZAoTn5e3cdi3w4nUJAYRX5NBK7bbUjpNaREx71HQ6MvniL7
Q7vnxeDQqs1H/7OGpIcNa7NzxyY0esuaeOgu//WQjOvQBOgrqCg2Uv+5269D82OSmELQxMWhkgID
oaG/+SVFg5JSX07/ZZLVuWulJdl1lQ7HJP9eaJBBU7Ub6KierogKBwF51rmiyzXbxVV0CUFBEliD
+d02WqXlC+MKVykCkTSyCViNHGxHOP4UJPDzCibkF2keweOMf0pPcyf1hC40p3WliPTf+rjAWki8
+4iwLyLpZTDwLb8u1bi6jcnEvKVn764bhgD8TdaOzYfUdchrmae3+ND82fyXvyXXlf7xWGvi926G
Fuoy0lCU1ovhqi0elMpWuY9aQiE9ww0xqrzz1YnlvGXrbtxDoaKRMhi9YzbslTTW+KfmGCe8D+Ae
QV55to4YbPRugI/EXQ1cL/rfE0zKLTHGo5MpYcRNI2nB8UP85dw1bJhuTi478nQAaxIfTsrgBL2u
lzLApII1B2j9m+t/CorsVUc+6ZKmEf/6fb1WnNNo0QDBY4yMrxnLwFWKL/HESoD9Mjf1CoYpFXDQ
iWRCL8CnxkJHnUuGZm57lCBNzvi9NC7wtkZs/bDfnVmN5I707VmdPDwWme54j/kXlpfqWiI3C+Yb
Wx5cd0xnJIbAkvfxTfSALXTSy4vk3fLQh4d0V8CkAnw4ncwYcWtYRP8iGkkPzTnaf8wGTU5/yiq9
nyBJ81W84QueBmyzqAgug3fjjYVXAGCSWF7JpcKI59Oo633uWay5lsYBPNi+OqXJYh5+F6hKAb5g
JpSBZm2684nwI8bTgfc2pFvU1+MGKxDVsA9A2yEzV0d6iUMMbLZ1Nzz1U6krCFXb6xkNKXfPCeRy
ZBH8Nq/1N6XfRKcmVCNYYwj73ruClFEhW/BMGtItZo+BFL9jHncEMtv2BAcRTHyXZGtQWy99p78M
h0FgkOfFjWE7yruoxHayPA2PlnZFQH5AaE7GaShYJguk89DhoZjILZFtC0GyXZaJDGS1vRkRtdtc
2JtSBwHiWS+omsB949ZD4F4M7ZgX+WvhBGlMv+p1Uugy1vaUB++0nergnWStwvcfQtO/ZTuJqzao
OvRppfvff8BpJTKShEMENSTYGH1uA/SoX7aHsSfWELGswGXcpYBBxp1jg+4/W8mo5XduSsePpu2z
bq5NcEI62RT/fKEHWCyIoMYUBT1lD8vhtCTklhzPYu6w57vVS8I0Ref8JqrOHj7nxLqbEPZQF6P2
llBOG61f6SOXQbsNVd3pOTSl3PBQIzpvu62Jdjhn3iq0Y0PnNPMZBD36sBUN3vxTJ2GWpVivJ0gj
PfZbJix7+VpHVC0lw5Kjk67DX8scCAkN60xwnyCyZZB7djjaYwQcm6pA1hq7qPMP83f3Aur6qADY
f/umlGD7Suz3/N5PYUAYgCLkLOpTpnUUmBnjxfmG2erOf6OeCVrX6/3rOFnbD7bJfFk1X4GF/hTk
xM3QR7kyTIqtNA/q43G4iQ/7afNm3VkOjHcXMJTYxc8HQuBM8XH8g2cZtbINz5NF1g6Pi5avvFMn
zWBIZ0bgvOmySKqODqbvcWVsXd6Tgzk6U1UQuIuScObVIrX1/PXoqNMjEdVbAJt8mbfxr1fnSjAa
+5WfeaUP1N0vHI0kB6H08ilrUNgO+zQfUgkfgchA26pIoyVhX2iy0HWbVeS36vYo75n9VyHPF2vd
mxbn5DtoMFSKkq6Vq0XOp5tvP1JlOA27d41CSNYnI94mh8WuTkbGiskbBlnuRv5cWHQeSWIN/T7W
zYidH912FErkJG7EtjFOFT7U69nt9VtkFxBOT313y8I7ljKz6GlLS8xM+VIC5nApEp1Zr+6BdMA1
ZCJn8uoFQG/hoLAz7i+7oS2WNFdBJH3qCtfOI94uJqUhXxNkk/MUMmWVQJYTnlk3WQgO/GSxv7/T
MbkGfxsfwwlqwVp6M6g5HYrDzEOs031iA/im6nPtpUIJJH/pll37KJ2hr2zh0zwJKNjcIo9sR9nk
Tp1JtjdAVfgXPXuGv2i62NJlzTbtO08Ft7VFmzBwciFknQzPkXqGqJsTJ5o+Hw9SRcdxGszNAA4d
t3lfhe20OXbXAOXdE8nrKfK/qlRI/06yL+2LUchtcb17T5VZHVQ/Unslpxk4HuDdG0YSUvZbYOFT
eKjBwz5aOceABG9wy47ZG9iEHzBFNIirSWj1k7KHCoOBfssuM9Zz1RX81uAXRJjo1VlucknjIcem
fAyePrOQfwQ7w7kzewZxYMqusAX/P3U97qZ6EMp9S/gJyVEHRJYdXrFCMnyO3RLSSxXHJ3aNMmYj
LBE7eEOtSY8MhPqJOd42kOVchDmaPf9+ag3qhMcZdvF3+2jnLrL16HP7FTkLmudzIalURjc/heGw
8M84VJLj6AnYgHVq2ISDAZGzREVw9lOQwLgubgfT8/KcVewi/HqehnecSMrLmYQEvZE39zZfRSXW
JAxLDFpmMSwGLaq5xdltRl9zMXsrB6QkufjkeDnK4qalmkkK1k4sAQ+Kn8EzeIczOcJSCoFgnsx8
UZwOOqIrmzi4y6yLJlBpaE2oObXFJgLOFQq/B4DJj0QKBHfbjpqfzhV9xINKsrIUsvX6fUs7MX5F
/R+QrMH3Hi0ze00IWSEiOmTdK49WivmTXAeGm0Q1xgR+vIrQ5SWD+hHJDzoabtK0WkHS2rxJ91zp
A5+QORFExZxquST2vl9k8fTmVAgZledKx6ttckhWXRdOgZaBmKAilh6441pWpEImHSruWZEijsaa
dtp99k8iC7P7HXZxAnVTFWMpGP+E1JJljNDzi6zSxcLyZ5LBjkRGQqIyUl7J1H1j3TGse0t0+/rn
zDzBwh6j4tJbv02DemoRuhJoM1EDdOJbpHxVM/z+4nWVbA+X4DsjfOVzCWD8/GlIR0sKbRM8qI5D
S7WT/CzUNqHbot6CuR1tWtH0hqj+slRQNYR1DvPkDmE9K8DytHcznXOTEvbP8R83N1A8jYNYSkZ0
wCD42mURhHbFimIHrs7OwhH5X9rQcV9VZus2XX3KT87Tx9hXEgSHxyWUM83MNJwjdbDMnURvQemk
o8Fy+BSBqnjsf5KJxNNwV62+POm0Oa9oKMQHQcJkpHjKe/9MSFY7jOy+CXn1yFa6KarkBTTRwHF+
mVArLb+NrmOM9gYnUKiB4IqmFBqLVhuFW9cQwZ610rgt9MNKj+GK/5kfIGxR4FEABqAyGLm3ZWcs
0hIMdWuilRwb5BSIxORYMbudGF/epIVq9IkHpyCCsJi6CQQNTr+U9w19wr0wjzaTkW6jJgG/VVFG
hkZOlZ3aITuudEiKn2sMnhuswht8QyiJH6XLNL3bl5EuWLpZJXPRIOFj4uPaa/sjz8Uqz9ZQ1Lac
swDSY8K1Q7H0mLdi5gugeLfJjOjdMCa1LayqjZXEDbDT+xh4KQg66k79LZ6pSTVg5absQKtKCjbt
NsFakUuMHEHB4x8oh44jYb/VYf3G+36e0tDFlF16ztrWZt16xwcR6Kdgb9oJt2lrcL9UPwaoAClk
E3aViOsImNpAPowSX+w33araxpamdXj9SPetbWzLFQjdhzmm/tmJQJ8KM9RxSWnQUaAMX8Nb7FiI
PaeU+9mQEXfUZZQB6hIwsrYrLVo8hmjYEyRSagbVlDWJ9SOGzXjMQ6/CrAUlRxnqGKXEqchfnP1e
VdNLYEPKQ3LbVDovAEL2laACxr3j0enezPxYcBBM9GhGcjT0RkCV5F4EcKQD4BtjGrcwn2+Sw0Fa
iPI2u7ZTU4iaRlswLp1WAFTu3rIP9zqTJYbSnBWjTGPqmjEH/7wS8b2EmMqyuWZMEpDPVOX/uRgP
KfvhrvDt6xKtBhUKeR1vO1ulySrErsUUeV5vQlT1UryXc9kjaWs/Lx7LRXbxVvkxjXWfLH2qJoo0
UzcLzm9GnlQ5p0O39MVpdqtXq8NgaPZFaKXm4r3Yuj2NpoK9/Qn1+m3hfv41YJpiiuijfW9S785l
NPO2pYgXTFB8tQGiv7a/Lkt4SljvEiQ9QnVRcjl/8MwuKuFw8IPt+1zZIFv155+AsGipCizYkRnb
mV2onKJEVPsPhYXEksQOvtYYE1HDbPtO/OSt1nShuly6j4VWgFll5yvNyxrKSnONsdcALzNKlaxQ
/C/uwZOhF5uFIGE1hI2Nn9Tj18A/btrK3cB3WbBd+/9r4f7TzJ6vlUca98f+iK0BjLDrDuTciKUv
8wPzHHBszk17gZ9U0UZJoIi1TIWlC0z28aNRr40f2GEOQ6jcPXyxNtJMyGzsJgOGxEQiCB6J7aKG
dqoayYdqQXi2MZQCrMadoMeXULfPqcQ9nDthLDZOkTsoXXe/JEkaQIUOq3pR59b6v/GnQyhEm46L
SqII0yVBWARnxO9M1u+HHTBxyc+19qkXIHmDLuughYYAARMqL3mhynXb9GkD3BgJNARtORN9fJ1+
/evjDDQBN7wdPuCKShlJKW7FgBD4RnTP3yGDBGMmncHm6a0Cg+iHTIdlRRSHH9+WBPva23Kh1xEB
e/0oIrn+jDEStUsu+uXKerVss+iOda++ZNRpkxmM3JjZmV6inS5rcqUo8dN6J6Y/+5evzDqF10BE
HKiH4ii6tEUUEVszCctNbfClJbg0/ZLwoejLbD2nks+NTrA0jpHN2PZFDZezpx8FZtE/rC3DRsLC
SZfLW7EtHRAeV8TVPt0f+eokyeZEekWjIwZQ9ELEMbxtL6Fvx75KgMQrFVPU6p4sA4dMcRgYKnAb
FU7Sn0PMx5RA8JsjpC1yU8/a/N4xeS2rLxzTYCeWWAfBI+xmQv77RgpaKAPg/2kDiBzib9CedFlv
WIalpKZCzG2je6DuMyNZyEIFsEug4rcy0lfHh4L3lsT/EVX33D/S9gP/ElHLHlz1ZUW1onHMXgLj
eApZAWG2s2XxNyTL3gHbY2L444BHHR8Px98+0oQXxWpCRkyDzcFpkcmAQx/kEd5IjXA+BUh8JWP4
N47ABykQ93KLPuYTCDqBA32Yxew3XG4bsPbUTpjv3duYL9kO6EDQmyv6TojZ4f5WaqWkUhVY+AH5
eXaELtFt+BcPZEimr4i3Y4aDlCQDIOxpsokcHegzAe9CRWt5px2SwQFIJMqcZQyTl6w2GrH0HPdk
VKLx4xgTh9TmRjE69nouRK8RlD+u3WDWcEkjrKdBhmrqzumDpReIxvLwkqmS3PXdfseixiXLWWkO
xzztujXA8JhIuSVwevLM+FVznZTSP84MjdaRjwuRDqJB1Yly1G9EiPrEm3imFJtqdlF1ScutTVht
7Px1ipbPLPoN+ifnnHTEAR5kVj8oG6pxN+0NLRZLeEFJRrsV270946tZB8fV+d8bieavgjstbt0v
isRU1tLAJVoJWwI55et6Jg8R2Uhd7PfllON5I/gQUvFKIWe+RwtoAKZx1ewD9W12fqn3AqvHl7Lc
Nq9Vp8wADwHGdNaTHz0R2ItI14bfOlwJeZDEHo1CSMHpwfhsALnf7oN93dr5yfdJ5zFaylXa8nFG
tDfjQGJZUvuwGSFkk9ODvStj+pOtcXw9Udk5/xWKwYxVeUcJ/e10v9jQUr7DKdxZRb56iHZX6m/g
hvmb4E3klCmq6xCIqXpTHHOm1Aa1u1Hd9fqzbIypI/1yuD49my5plUHRGC6/D2aVF1FxiFLtmJNc
sfxCmRrKD4fq0lKPgycvjSCF9qxsvjZJEeaZRgClTAb4cbgLgbHJaBivPZgK8DQlKIwkgfgO7aZH
+pe9Hut9/XIRp3BmCLoaQmbnY0gJzoxBJTlj8t4tKBBGa4dKPyc6Z42tPSJyk3C1ZeM9o2CZbK34
ZKe8l9KoLgRp0jf3B7e1hPz6h95P87tiQqKaEfJPE3b4nPM2ySZozMqRpx3u7ycP5/Xtwbm88M3R
XeqnyxytF+eSt9i3+zYTa4dvhz9mwC+qSD7zf2zYkqzpQDP5DdojlxxcHykl8BT6dZGxbJtMNxPH
gsDefRWbf0Zqn1ICxyw7PE6/Y1iXVTlGrV5K318fHE4diBnAl2JY43c2Mpw5MBpF39dG6W9rpsgj
GxB6rHoF+GeRDpugeCgS9+xULD1bRsMYdWMd2J9un20azQew8TqtpzVdDCRXPyHw6VRBxtYtnOc7
B4J6CfwKOzOMNfpQPGMwtd0pL/4XZIhwN5b/j0PqOACQ5s+K5sL4vFo6K8iTOn99twNoV8qvTyok
jLtkWZOAH78pUpczbLRWeRYO9f2S+eoGSAb0iYGUdlqoYBsmAnrK+vfpB7Jiuz3Whgw2omgVpgyp
PCI2hMecx33Zi01YJmee8pDCbuc7OyF+F9uNZjbUBPknvXsFmDQwonAZuSBmfdRz7F2K68ZPfoG4
s/CmNUrAmH3i5p6b0EzAa/v38ggjSuCmWVe7dNN2ALVFuSV/TEgC4VjU8bb9+ebMm4X5/urh6hvj
RiHlMxMh6UtDyioN0ZDXrVFDN1O9QIN+8VAnB08WCwBzRq8HwxBlL8Sjp9mBkcQXn5KKl5IrRO5K
IuVwmbOQRgDmuq21YIGIP7YjgWgB1/Hajxl90Dz3p5YbYPLDMBZ43HhgJEzqIGpiFiHbzhZq2KYj
aGKDZIMN3whnPRqlVq46tc/IBwlk3xmCrXgKtXBbUr104gt0W2LUp+JFdAqYIkimI/NW7Z36KukM
YB+bJu2tpkhGzzV+9Y7gaxtt43R8z/YEaNBuyxMxdOQ2nR6y8oRdeMdVS336pbmSC9vOQvSymIFV
/8BbI2zXwithSQsxbndBz0sFCGd0lPoJp9O9ZIXmhLTrWb7wZX4N+YMaD2YMz0Iu/s5SXz3N2wZe
B8i1uvlJCjAYXwV/W9/AdWSUSlCjEBm2m8JTD1MZjUri7jUZVzwcWaV2+euh6cXylMmmPRcQpQsL
p7GHBNyvIYR8+Z9zKL2FJfs/9XlybcL8xxfuz4amyYw0jMTLnrX19ELOz6dpTSi9SbeaZAxK731Q
BlgiFwWw2wp6qu4UB4G1opqHqb9PMZNeVJ0qHsBvdQLhbiHbVw00CzgiNE0FqxJivxx+i6PvpRk1
7+mc7v1Br5wr5QcuhM2A8DsBCTgGJO2VLMWnKEOj2uwAjDQkwXwLsIJ0+dCYh59b+9A3T4Pi0fKJ
Yc7aIHdo+ogBH/q/3rVnlbt91kqD8J8NRqp5qnDMz/gMYWVnrnQqpCZBrjvO62k5bCpZNtGW2NJ8
7+PXV5jmpycvVztLF8UKsGGayUCHqxvJCXd3RStW2q6fhfRqB7NpGi55ju+CYpwmkMFcyJ57D2s4
UNuKz7yghPh5hD6IHq3ZmBJo5msv3Hd2fp2Q+Zi7QSbNFwhxaMw9/wrI9YBOFSwAoNKVPcX5NOoh
eqksELap2TL7oxSDh4C7ElWncLElfbH2fMg2pgNFtXiGkBdRMsjo6DiJdu+Xg/qWFFeTqFrHaQDp
bMt177/MbPWc3hs0zLVumkyx/9yOmqLsaI96uwxpATxcwOJf1WrXYNVf4P4xP36l5gD7tStzyLEs
YSBAOkH1AafXEig9nmoh30Afvd3YuPEUMUrfjqzrqXndUXALyau1VrkP2Mde81MDTx1Yn/E+2ax6
IfR4u4MNkdm3kiRUTl5yhHXM3xJHWW921J/sdqPPxTY28neVHqh3UYFcka1SYkPF0IKdN2+zHqDS
PT5aFBIrCdMkvwd7IJivyFt7I9GMlRNMoadxWliG2TfaOHN+dQOKyJIcFzX85eyjBA5cvmKqBJ/K
3us5poJybGaOJDC7IA+nYs9TmgEDJApuaQBkiLM+EciTOnwex6B2RSipr9is9iaoGPBqomWqSl/+
h9vsVcbH8btnjjShZmlczqFsD5OpMfDM3n7bI9SiWnFjX3+hZNqL9iyyy+wYu3iuksxZWtCV9L0s
WTur+eZSN/ZHjo9GG6k1GHuOlwtNR1nZgaiptkx8pkbm/atJDOoaEmaDzSKJiG1iMG5WKUKTaXSQ
PfKTkYSKDmZfuulfmL7JA911Q6iZ2U1WrUVIimyyqwzsh2cy0twC0L2BV80bbGel4Wzyjvx1gcIF
n0OYQIy2IAyjVg2wOUDcsVV6Ts5WmM9XWBrFKHjPZmnE/+Y2NhBh1G4AOGxWOUcaVtnzLCyWZMiV
SM/FirKoeAfBFu+Ei0DszJ1G0NzVqoWBqSGJ87vRZbsnVXGMyzc+V7p7AGIgtJ5UydJpWBh/5N+p
hO2b4E7q7/mmus5H2P+w4jKFiwmE9C7qYcNcs1agpO2d2FfXmt42iLmBoGNnvUMJpGOL1UDcUPYb
p7f2nsSJYRnnP4lR9mq4KU4zNLpQLZTKGSmNfsK1C3HmALVkj7OVniYCn+j+7E+gqbYZvFa3vBxm
mmHhjiZvoAobbw41pLh/YduFKpthz7B5IszkygwFzQfnxT/PS1DC5+4hAXf+Xw5Hv6inLgF4bhlr
FH3B9/ucQAbETNIW6jVi1/mVnPB7AegypCGvnhYAf6qYEwlopl/ne7IHlEKIY3fxZHt6gfuheX+L
ZdnB/i2YgeZ/9NIsJXOXTf38SwhVJKhroWvhAMXiaUvfet8C5J0lTWU1IL/f8cnxh+Wh/koTzXVZ
Edn4OPhB6dozx/Fju0X5XFN3gFij/7R9qPR0nDnE4nosAKxunlCkqDIxSz4wNZvcjbhS+rYDaCEk
cn8N41TveJrAC2CkvtnkEUNUh5c7kN3kWeiR3CrzWWgxFTHe9+dhmAWLevbeV4BnGOJ9mW+SXIEB
SEUfVTy8dSDHTUMHigVl8oMopKwNO/l44dZ4mfsKNBbRTjxlxQM9Dao5SFlKEryAl+FoQW4tO1J8
Ws9dNCWnwnU/xEamvbpmB5raASP2Y71IBUFUVTfsV0TTJrtw6Vkobvgdf8gL+p6j8OeNapMn7wa+
EIHFVsJmRE1UFfVKH5b59e/Lo3QurwbiYm78lNa1Y/4/Nkp7EYpXNgVzDKXbE9RiVMccRB7aib8b
oNZs6ovJeVJb9kLHRQYehKGr89dhXuLd8dh86rdPgN7iXakM7xmbTHtSW3XP2olzDzrjbBMCOyvq
9/zcgZTl7r39+1aqE6i94tP3UkDoo9V17ApugtJZATJmKMk9yMlWKCF8IoZHq+fzJI6OS8uw556M
3BWGpBeKmTOxAYLrzELbE/AMYla5EWELDTQn7Htc71YVSXKpPpGjH7suNP+eAtxKFKbGNwEfoBDz
HxzCr7zxxW2UPZxZnjnFrvQNUoRgSXua3Hav82mbYCWGb8UaiZawHKY00FcTbyEnqHK2vlkvVoQc
AHO84DFm2+ybW27yEjaLnfu/XtFAgxHXOnMRh+tlpAS0pEYH91qE3JSB2T6jx285jC1ZuDJOvlfT
1iaJMAy2GVy+c2Mbd3sXNXRw4HIgGDR6udFpDLN0iXzsr0uQK5wgkQM8j2yAoSaVc2orMPFfDvGw
F8+rrXC9mgm+MjWWulBhMdybzKRsd5A1FjzvsOe/YQKCBk+VJa3Tns1YGmUxTMVXjxYmmGFrJ6NK
mUfUb0tJUR/P3T2HvPrdY7qG5QYGdiBd4TK2hOcCwcwkJMwJGPrm5LO66jWNFEspHGaOjupwpIXk
7camLjr/v8asEqloPHUsUdEAUQSBJcJKput/iEaEClXg8ut+0T9kmGlUv28pFP1kicPT3qXkunE3
qaUe5IB3Z1+LyU93ho+E5WThKY3kF+GvayuA38AEtPqbyfyzSVxYcRVsSOSCFI9W/eFgpOTpvKr3
MBORzqgVcJm8FtEUNtF1ZPs1lEQaAxM5JDBlcNUYwDzMwYbDhYW+RyjXcjzN8Rc+f0zuBVxFYVbW
2Mvocmql9ceBMp/7PZEU+wk3zouW4IImntpLey49Zojl6NjmEPoWQG9cw/xT0FbUEWMCE1KuXSgG
moCBDA8PUiR0CMZGWS1IKKD5xKVeIBVZxPJvzgXQxO4USe2o4xTTY/S9dJdH2xwvLsbZf6TBVlWW
5tDp5I1dOxrM0suu68MJB+YmzzQZ1F9bsktmvILN+topS8a7cttT7AWdTuqnhT6y1towm4T83NjA
LqqEqKfMCPPN2cSTj0Nk2O4SOX1XGu/Slg03uB4PQewR5aumqdLM3KlQhILX1oWxosz93Rhc2Ivz
mz/c6phG+40fPSV3+XJAFhcvyRQIGpVz6DF1HZC+XEIsS/nr76LlZbucX/FWvKmLT1VTc5pXG1gQ
nlyZKZjRYA2n1d6M0O4Jag74YpNTSNMe48vrVBmH6b+7Ii7Wa+74dGZS93tw3rlitI/9q209aPBr
6EeXaoIUFjjM+zhJE5AgxWtKvWO4RnGovdPuOvwkh/Nzk6htRVJf6Ss+uN6oTJHbir6PTWzP+KrH
4R7JDHwmvqLJU7omeWlOFjaiBmIc2Ipm3wf4T3qBPmDi9hwcUFWNA6ixLfR33ao/d3RGYCcxdr9I
EYb6WERN7gGB+x76RxIoz7NKW1CsfgfN8X2I9DZelS++n891PypbC+8AC3KbMI4vDHL70HvBXWVe
8Pnxq73P66b+qgeYBDJGoF/FMsNpVP5gb/WyX0PvJJTSgIj+PbHF6Dx+7AkJiV2Hi8Y/4ynDum4q
9Ugw7UKo2KKiGvGdy6wqlIRC0O7yx2M+GTVPeuW+HPkeqr0SKFSGxj6XwOJLa2bDxIS3xCx1fc7/
rU3X0gq97xHOB+qnOc9VqP6vcVVoeU1TixrAdTuo9yIeOYpmMFAOnmcr0kK1OfmqunPVIKXN1dXG
90TpzOV8HVX0P6XiF1vUAgXO2nV/UTggveGUD9JB/oeKlrMnyQ8VV1HpkoLBrOrUpim2kNBgCBqY
EZfm6BdVJSzAk6/ixFCVtvbOEeu3duBr3FFzpRuQoi/VIb+I1aTK5ctT/8XdNdVUIsNNvrhmL+0k
oeBG9CG9Y8MdiYQvK1rXcmW+IpPDbjzo5/P0Wdq3SpF0tax47r9x04ib+1T9GkojO8RiFud1J1We
b8uyLuB2H1J1lOll07OjXjLO9kPahc2tiiwmZ+ffoNl9nScjDblAbMBKE/pw0ODV3eww1piokiER
WNQwZDDHVrHq9ZmhXR5T3ntgB5k05CYI6zS83pZA26hB9CzO0woz5sfwU8e5J4NZzK6/+AlkKjxo
o4WAVMqtxlCVyxc/DVJLbbM1jRSRxtB2ZlGbzChzzNtooHeqxPpkACWCmgsEsWK0bsO2BGldQVD0
ax2fY5Uc+2n/nWo0uEPUAvU4VqsrbcjXJV2ONwLLQ6Ja4brmPiCph4EgOtYXddmRpjXiKl24t2HT
QItx19CtiKSzYQ3wEwrOwriLTMKzvA3Y5Z+iiKxc0Lk/prAmp/kZfkCfurYQYwO0dh66o6DeRc09
/TNESTcsRnEXdzkcIWLMNbRIDTSoiCvnb53Akmsgsxh5kPrOhnJGcm2syktA4q9xDOfkoilfVlQq
s03crv5qqHG24vdeUr0we65Doq+12wB6FKH1doTHaHLjNpKReJ54a8bCB00Wr29yuPy3+i81kvdD
/ttx9lRsnUsZWPxXXX8KJwJX0HzVgqqpE624aoPa/2mzSjvB4PGWjP3DjCGUEHYtT80IQPXZTpse
nVQbF0GkwFlaLZX3eXrTkYe68uBGPYaPc+MBXrdtLKeFwsI1is0ieCD6ES8qQj93wpmxnqIcJV5u
OXh+pzIJVmQjVPj3Lq1ZY1p+brEeq1WKcU4zaWKk58YGKb1HmwIad5lk09HJW2ZxHkHOzmmcteUt
+7z3KRiZwU36iLiUUYkJa3BRsS47Xbl/0p04Rm3xeC2XWHfosVILXMkzKdT8te9IQbjvB6O/qEiy
9A4SJjcHpJ7FfRomS+VEivi+DPZNQNGVHTKZISVn+s9+uO880teUsezNsp4AT5tBENfo3MHNWiS7
Drw6gipdK6moab+3S+cw8al57O4kzQXnTM+jpYdvlaPVx+BCl12ySkYFrIE0iR5MO3T7DJAuMQhw
x2gAfOm/8vEO2rGcWN0I85N9wKMP8UNIzC2Rappq+nthgVXkL4Ly/RM2m8Ti92/ZXZnQ/bRSWjbL
7ECidydioWJ/MdDtUfTS+1vdBBMfrCOT+Yzj8S28hDE57KbKaQUY2WwID01m+jJdQP74pxKm7eNZ
9/8XVlHTPPqzEhoiVzknqYepy2vxu/thFO8KJHITOLY4i5zfE2HfZfckSjEMsU5RnrWTf57hq3KT
vUFPA6L+rSe2/7rhBJUVZ/0dKkwELV1TmJKSjoP44mwY7gR1Z8DpZQA84PWMpQsbGl0ErJxQu7Qn
kYktYb0J58QxPuGk8Ikj5rL0ZlIkBkkvvN6/4RPQ6hDvXWeaRCjA8uDPvpSrCHMDc2zmebt7YQTl
XT8kzxdo4eSziIe06OlvvkqExpkppoZmWDCXjkREuUuC/qwmvgZG7ck+8/0qzajEpqjP1dIME5KM
+qgk0EhXI6+yjCFeHuK3cuef+f4hbsAdsdnVCkWZkYr4qrvDbbKGDlInAZZF3DItauXrkKP/IwbZ
Aen2QmhR6Gor8G8gOLeaDdLmJgxIfpiWUnqdZ9iSnIhkVpeYNNAalMV8tqWpe0XcaLdScMHPumQJ
Q0Tge6A2n5AdWG69YG7aSkf59c8ozUI8+nDG1BtVqlLLcomS5hnJjjPXp7bHHgB1ipZcM5LMacul
jfQwUTwagzVBeKUnNrdlxFHb0EoQrrbP5Zyqgs4AWbKw420+i7rFXF5uf9MvTZt4A45aZ8hS6nwe
hvjnlmMdHklUqj0qGsV60NZLhj8+u+wVLkUxAk9xWmt+q+9p0S/MamW4PHCuV83NVLPP0rYa9SX0
ArdTXhkx33ND7AcFB+kehhQxf3tPIIZd2QxU4xhwMsBpw8ag5F00Q/K55cz/HeKGyYqW5kk67WKr
o3Uou+2hbs9kaIjtzYVH+6t0EXzLVEI3R56GY5ux4nkYyiky9tEffg+C/LMpP3hF0NeoEpQz+Iuh
LKd6NS1CLJ6vblvThs7yi66VU5jyZ7mY+pjQ7c8ifdKa6cJFUdSmBdcbBRxvC6EpeFNf7U9pmGFt
I1fBnmusWdA1mfEE7tZ3INu/rBIDV2ue80VQd6l5V+MM7kF+1wBmT2yNKWNcUCVR6GB9ePk1wWkf
SkIOgabHA4Z7RXY2He7JmNXF+Y6AYHw/QQx4PhBBEWutrR0u2VieM9gUD8JhSU+HfrDyP36QChA8
n0W0WyUY+q3F1kfYIxT8YtMpBOV3jXABZBTYZa3pR+hs/UiFfqQ3sAN/8/PMYLz7oN0Iki+ads3n
AiNs2JDhI/70IMCRXYtOG8HzR1vUat3xfjg/gga90IAMANc6IVf+M9DE+cdtEwFGvn1ONssxEnKK
ryMlKfwwihZOCrwfEoxKkgeORGYJRePF5U+K6zQSZywF7uvLeV5hnOUzuvz6ZNlB/rZz5fkLiDy0
GzkdoXuRSPOesruriiCubgqadVUnLozCaQrKUWzmEmAR3kb9EI+XblKxhDUTcyEa1xE3E5kS6sVP
6b7yJgFd8aDCiLj2l00k3Z5y4eEqVH8Pb196mDIUUuvEn6rXDhGWzfgG3fGElj7pWfZ21QToW7MX
vPsLUtAt1t9xSikCmb47KSA1ja6nBm+qD0cWoJELsr82b8Z/iS0ivtq3Zac3GXrJ73QS4fRMi4Jp
UN4t9wxoqQSbydWLrj9ANbYfpwodWmvW7J4lxQdlkPwzoAvK2aF7GfG+qb6FXyQZEzCdnU5z7zuM
yFWltJjz9Qv+eR5tBMGTLbaFRTcYoX6453v2F5XtOI0sjlmsOYKqsP9P+/ZCO8A7mTsMU+Ph3XJn
8n9DGnC5J7R4RKnGGhtlTETmJ00FI9YZYZCVg2pgT8i3gDzqp+BcGH/Xi88gr90mLgFJ7Je0ViD1
uTM4Wq2CY6nci1/SN/6CkGzRS2fqgcXf+Qpp6Ubzim72WpA54s1VGPJvNXM8d2nQQBxYndjUKj3y
TKguYw5G+GXnejofilYji0tob93wY01jxcBB1h71eaT4ZD4ulhTQJ5wQry8glXFlBEeumywpGV4b
cJFTiKrG78VyjHURmFuMgKICAdba0QMAXyd/hU7sUuDQmkXuqT0bEvIGE2lgKjhBJkHLh1zZz+H2
IQoSMIfmg+zKOiyciJzF03EQu06kJFMvGhQN0aFgYaDk/MhthVFh3HEMIONMxPcEtNqc3Ozgy3Ia
jvhScq7RW0FYuxxbNGx0/QZBqivxoaCvtwGaCJNouXirGegrTdaXJqkAB0S7WkW70nlBMEmZkloV
c9iye+8k9vcFZCpWmc0ZlxMxEARE0uiueFRJyt+cFfYmzTCid8GCAsDvRXetqdxZnpTs03yJbByB
qWvbh45Qr19gpKp0PYrx4U/jnqI7OSoWpx6H7RUbToED4o8CkT2RnZmhDT6NeVAFEBjxaGIM5TQ3
bHur7xkknyN2UjAiWomVXVEEnYYlhkWPxCqBxcmXS3yLVUyM9oD03fBe2bp0BGN1GJpXm+RWf3jo
tDHEiQ+qFzR5azCkH/fHkFqxUW9vdEvTQKTMwSKRsZ0cDL+lQtqzdSaTrm8Vb6x0W5zxBjCQj5ag
o09xRBTPllbVYHQst/lZ1wnoALMWnoA+Op8V/PE3gr1uHzJy1yL4UP+YjAy7S/wFYnrvCwKYW0NX
qf0mkDCn1wFWKgjTXWBSNYnzTlvNgVWG6zS0pWUhS1T6E3nC0t2mzP+4JaBqKyMPSKQrg9bIcI9D
1Ut3XqExGPreXk38hlWw+YZE6I41JGxLfaAoQanj93gaW6ZhZQ1sBI1RiK2QhhmZHo3079vXakm+
Z9kAbUui4NZxEvxJF6ZaRoKAsf4whRD1QfNew7AFZoDa2gxEccxgV2EmCHaBXunVFPBA8A8YvveL
ODowM6YxrkoGz6Qfa8RpdSNm98wsKhnKMg9n/Kp9E1htKaL7HnLPaRQHydveTmurwA8gOxd5OKWl
kRsiKEIiFdN8r62Q0z4cdytB+qdRDDtdRscWfFp17usXw5tDu5tStGl1P31p95MgykqlyYNxjB3L
bKKDeLNPCbGVDyjVtEh0yK7DFkchdmpOZUiYpjybgkOyOCc9sW4FaVse88O10Z7ERJFKer0aVlSy
6fbEqFtEX9VD+MrWcyE3FJRhm7M9KXIpYmOLRGxSRmSPD1/7TQZPNYVr13wy8b+/P5c4U+DjIH1V
bj0GzZpkmCLE2WfFted/W+Grfe6BGxACUtc26R523ifcCujritO+QK9eD/hSFXfmHCLMFCsOWBPg
CmqShGeGahuGHsvY6TlNiIsNLB2QeT0tmpl/qVdeb4d9PKW/c1c84FtRcHFoXzHzTunTxfykQl91
08BtVjhCBXD0SSXdG8U1JhsaNkXC6kCVzPrt+XHqUE75XK6OX4jmCxYf7o6pB3bQiS3R3zH9dPfQ
07PY6TF8gDOD/ctqG5xI5/E/Ib/5EDY5mpoZYIz4Zh/nd43+yYowoyWCce5BLOLz7F1rSYDivzOF
JH+yYF89h8s2WlXnmDrMs2EWA0oSNVuTV9ow5fA60eYr5o3eYescctiFlElh/JxgnD1tRkQr4bjm
kZgKgUqXnTRTdqVvvpcMpQjIDkmkhHfo5kyWng+IGf8yh0ZA9taabJ66oKwHeboHARtPru9Ga0dA
vzxV3p/Vtt+htJFCe/7yZ1E88S2u1xT9jc8vW+dkuIcYqpG6wsXaG65kvrQbIPPPvc7q22Nptsz6
ARXZXrcwy3fbn6dOEXN1HcbCBehy5Gqmrfld/uwf3nGLwtO3N5UbZ35p7a191kBZpDKlJ+aeMJlY
suoF/3SQB8jaa1GC1ZYyAl/XySTih3zdfYUKZz872LYDr9JgTKJShlPcBrdB4qV1v+fvFY0oST8c
WKNHfN+7pxqTPog1Jlqq+V26mSISBd9TWy/1ZpsIJinBNWBl9S6caBA1drJtsh5p6ORtvPoltI2i
a6UrGhsvs0FO0YyDkeX/mJxT0d2FyLWvndbP4sH2WpTxwvq6zUuM/9qppxDqjWv8PgmBbQJfiFB5
54rdTYwYfdhaGFn6uf/YLjCNbflRZh4bEIvfYBJAyTTJFhRuiPLreaKU51qLxV/lRz3M9vpaVb57
XqxR/e0Ew7hUiKNa5mrAh3Egd4M4T/I6RWuD0qCF7IHAXVNJL58D92HYuCHxLF2IpL/hbzPGEQj5
P3xdmOR6nVAbgRos2P3aMG3nc6MHf5FeNNVy/CZyQGaC93C7CuPXgnM9cptjL3+YI/NgKWwDhKWj
4ToXz8/Ethj9OxNZ0EG2Nt7Tr41DktrgumaiTX1W595P67ksLY6fnq71874I8HLtm5x6GdK/WRje
+ySpMEW/Pi17yLVCPwjpHaDWK4GlRqJ7JjtxJdiPp+vl0aHvYu4ulg4vI//RRPeMZsg3Nnza1qbO
40B44hfbBThEAMaeEwYzfJ9OjWEtho0qmMyZXAN39pgMGLPbAiBsGgAhsjnbMvYj+tGF21ZrukWt
gz2L/dddUBSmH26LmN2NtC+C57lmDJBORelDu2IgTwrm6Z74YHlcUZ4hF9JKD/5DU8lbBMt77Zjx
uxHjSURV7UR8GYzY8mxvQdYRWyQ4+rJjQNJ8BjlR7uGhniqiu9QJynezqzLFl8HOfQz/tuTcWOyV
QSp0GFfG+49lYOjOAMJ4NpL9+CRdcyPO2pQ6G8xdcE/R9Jt7o1bWIePzoVy3B+XitS0NxKIWjBce
9CnAkt5zZsRUnrf3ZUDL0vULdRXANMIme5eVSjRoPInFiSjPUum3v75HWKUql2fRGVGvo6aaigfN
BmOZJFMcpqO58ludlnuYNyhKo7iCXKjRyChN2yaDkwnhmurRujBEaO2RJJXSXXXWHjho9E9kRQ6m
Kyp6D8dxzP7JNoWt9F6B/aUuC7AzSjCzIHMTvqDZZQegcNQAQPM6Tokd/Ynmh0ZkvtrH79PYd/qw
F3gQfQ0DkpeHTvPiA3Kg0tbRKikyU8NumrHDccRyHzRkqeSNyO9DuKTo0LyHCCaP5sRpzRnIkN2N
qnI6T58HyKrDZi2QDPV/jna9Zfmhwv/7cQwDOttq3LF1EbMJnnG0BIp6E9ntlOLgQlXMERNfzSi5
55Kd7ljKX2NFwwrVPTqq/WFeVe5JSZoAYX71XaPA23N3Zn8+tqFWQHJnOVnmddouy+gY2hZrAhJK
QNWEUszSSE81H/kMdrRkgyiyG2jCTTmTADCj44OOSgKzxwcINrEATrEP0M8L867VyX97kYsTjV32
K3JeUrBPHbfqoNF6UoUEGRW2O3C2pxnXYzr0TqepOkumYG9L0F4RiGmAN4YXnJjgmvxyrOkNqArf
6YF+yoVHeKx0mosdctV//Zx5X9pHXtu4W0sHx4oHjm4uZjYp2XFVc7csmstNe34TnkYKi7Uuk6QP
JQqD6Z0n55/b86sMSojIUac1ZNQ7YLMkWWyHb8eVjMZjMt6ZHj+ytFvZ819M9DAWPQO7P3+rYeZT
7rSKLkbtQysVGzB25PLkhzMY8wg4lGVvngs6pzpVekn1lNhycGbnJnn+I0zoHibLvTWz49bA19P5
FwIuIeo5/4gtIrvbeKbNnwQgPwvRpiFmJkAmglTIH9WP4Y8xQd8LrsS7CQp610dOU1OOHrirao35
e+j3QN77Fa8cWNTcFnF49y7DS1bH3YPVDoi9JA2m2HK9lp3csd3Nptf9CzaU3WSqd/DOeJCYJAHZ
Hyewe6fS+X1P3o+ZxBFlT7M/phDPOdV08lOoQ06RkHD0sIdS/aA1UeYvHN06VVvi9fEdr71KPIpe
qtf4+gSqlmonDMsZGN831fvIhn0Oi49hrj2Nzk+eiOD7M38dtedJMUg50ZRfAKhe41W6GoJ5Wg90
Lj5q0q2adkgh6nxpq4KLFK4R+Xw+O3I7rH7cQJht+xyPpRBhVpaccPUxlaB9lB5EiuGgpbDV/wqn
EcaBxoxWo4puhpYF+EUhxm8/HAXnOVYaUwXnBZYWoaZH8l8JtGF+ej14ROzv/MCDPQxZnl7cDp3f
DbYtlHt1lwsfkaGFUPusoGW+N1Cqfp/ExTLJUJLSSmIWzu+h/CsyAqrfUmuMZAgUYsqyKli6WtrQ
KY6h8NA8jcqAWyqeVPo7DJlrBVQLeoJLRWtaIk+1CoRCHjafeGKIfd6ebGu+Nv0WK+8nNshs4T+K
j1AiUwM/p03BfcYaYwCvCxBICzlgLSFVvnVveBjGQVkT1RMqPW5NPamE2plC1uIMYBmF0V6jAJHz
lJKZHze+l1ZMXRc8Q2w46JL6dw+eCcDN2VKZuc7/TBThXlDUjCnUh/Z+0WJtJTTjl8jrd7PGjdla
yXC4pWhTN1FdPiydeJgfknAKGix8P02WhqQH4jDLSFofl1scOs1biPx2tOgMfSVLdxcFLqPlpc+K
0bahulNagZMYOZWzjz071YShH3BOWwXlc7AT0YUh0MlCDiEXYzSK2Y6p6Lul6TiSKwyLOF9YaneO
9ycEmB1KgKZrSDAYmq9QXImlKWd3wozIXVZ+ioBtVbXWovvFebPrHvNt3smVc9nMjVgU+BvY9MZC
A/y7UeKurU83m51Oc+izO1tC2WLPveiPEDNxnIwVkrR9KXRWHwIZ56IoVXGJE7NVP1ShXTCSWVFY
DABpLjDm5XJaLcA3fYNJuzbRbPFo61x5NcE2Ge3J00YkuRvnA8smchrsmPOpbUTYzDFFRQ15uJnz
H0VfE0uiILNXTHcNdZ1fRsM6OwNQCUXnxcnTEP53me9qUe+DHzz/VNQo4Wz9AVg2gaj0Cq5va0n6
ux7Ob9tiLQkq4jLT3YkQJgL1MUzxAOz6SwzUDQeRl/wwouz0rLvzYKCZJ1EgRlcySUAaw+H6/pKV
jmjlookA4F9tGNUoCiOVAMN+pGpsaoqjNAoWXF+6anjCqYDYzsddwju76HImEIxZAHfOYOP2+fJn
eyPjW6GGrnjq/iIg0V0HptfiuGsHprVvva68zzGDWiRsv/kwXUpa/l4YkpmpKhSv0mnjjuyM4CFd
w/VOdfJrkX8TrYKs5nzd2UdW8hi2y01hfD3nCdL6/zO6T6fnPpVvxrfnUjZZvCtMT9jX6oaLaxhT
a9v2K/HUbXtgUGVIiLvEVbdJhsQrQlRVUk9thgWeQ2k3gjf/5OS0ZPnSLxD0Odsxq78TL+3F6v9s
GY82zrNCcb5Cu4rwWoM2qHY3JkIjHKAS60+RzNkN+MhyQSOXhwh0JKvimPSqJmxjnevTK1CUndq1
v1bmqYXxg9GZu+dfgKotB8t+spOzZRPX6C3Fxp+JEmHSyo7Q1v4JhvBw4K/Itemv0c28j7XBkTMd
N9GyqK8OB2JhTm66K5lqL9QH4vWD6wrkD6rJv9DaTYCGYeSz3zyEkJGQkIP/RQby2ANyouqEgIjI
bFTgkQphQuzeLoaVzbpCSmyao6XZu8ufnn/Wl8Y4cXp595wsIUbPm15RYLXTSAaA1ZF5TzMiKR30
5/eFQhwwAOvCy4FWoJH7OvI5ctzK2Vt/TVXyqxDVER0ciM49d/vhOnaIQxayDnq5G9jUXez8M8Tv
vMJabVO/lrp/0iHt0pXRTGAi9o+eKrb4Uy5Q3w/NcgpqL7csGE4ThxGAIvvgyQ3ZoOQVaSh2sP1O
DWhU+N6v9OIlNyr6fvJl0TXVcr04vPPTuH3eDmS64ELp9aCPzPhR40v/X2niAsAeCYL3gurVqkQb
ybVJk7eQ5x6zTsaBkAMt39jkPW1TqqD+mgJ7dxjbYvhmwlC9KKpwGrhdM2RSPKweFUmT5OzfABjE
7O2YACakZy8XfH4UJK7PJwKPR08HvRJLFJ2/cLbhOI2BkzSYGBG3T3VQJjws+wF/PUx66vK7aQLl
h/CSTBMT+h3hh2SbUo5zKVBUVdBffppLEeZl4EthGB5iZpHfQKeveMqrEepcyKTexCT5wnunuety
PBg8jQz6OjSYdZ7OLsCGKsLpTmvCUfBa0vvIX67d8SYFsAaGUPTGloxAFwmTh37KkL3uc+fx5Fty
WgUlyxgqBrfHYF2EM6gfNdak8tbGi/zpeQFajQ0IRNIkGyYSvBEf1+oLwzRA61bVMHEL3gWN5E7n
g3kq6QachUqO/MLPVPOPF+ya11DcxC7ste1Lvgt3U9rhgQ1qXFuLGiuIRnVmXgQGvXVC6SbhRyGb
fnskdRjIHLeJ1bGuLHWlAQCuXPwxkLtep/9twOY996VZmZOuTYIqMKQvtRUa3THY/17Uttp1LjN7
SQzpEyKXRU1WBGptJwgq4zsjze7S9OCxOH/Dtx12TD62fdAJsqMoD/we6NECph+CeK5/HOBZamWI
kczGn/+b0OBZ4/Budk5zKQD6LNaJK8GGgI61F4PX6eHk7vug4xEemBYV1eKnK/OUDryuh9piohwG
q+zMqapihOvHC3o6CNwtJ44kxZFvmSOuuLFfzQy090Ndq/rLp2hVtk2WrElLs775KxLvR3CVBzAc
1AXwFoqzxGkYfI7TEOIBrGFqun7gde9k4YBRICaFn4UeiBlLeQgqnmTTgiVL8UZ1TVW856E8yYk+
0JQ4zkaBXuNtgC/zBl8/IJ82jR3qd0Q443Eseug4BbigGBMQ3RR1Kw4AfxuL8exwAQKmbf94PZ9r
NUp3/O+nW4UlgO/fycSEaasNzfw1/+McPkA7GNuHisO5YUIGcrISo0qf2RxajXR9epVxOut0i7Mx
bA1fwiMcIf08aXG3RrO0RbU4IiQS9NM9f2aocGMpQhYqS1KH/oW67lvrom7sHZJxogsNpO1J7UjD
OgzK8IdoG6owG6jUsXW2J1859QEqLBRT9gzacCgp/HJblw3fi17TlpUMCTjYjg8ywDw1BrYsMcQf
HXy06ub8px9wXNVVBfw1nCepSroAyZfzMyEfsBtnMJtRQTyM4C5JgkIZcwN0RaQM8NQS7+hNDEm+
doKpkTORB7syupdC4Mxz9Q3wKlFoRlXcwoDPNBD+2Dl+qb3J/mCjFlEnZEe6LVIeocY1gQCzABgR
pOYALroiSNu70ShbhWIHQzBX2HMWywlJoXncSZq+/3x5MS6mkrcr5TyS4tLhGf3a/sKBo5c90PQP
Sy8NfTmdNgLguI+PdA7PW51zzm9v+Rm86A614sTZNyb2PVHdOtXrA8CzehDI8siguwR2PI7N03IK
2Dw6HU2fNQ0cJVQumhdJNXGWEGN3XkFQT8w/naEtS87dgenlfvTq7bO3v9Ig1mLJE8Qds1000K2e
aWW9DsEpxqIB80aOpcO7AoKRQ90vQsP1U0XrSyE8fVcCe9khz8E2PJvXzc6f1lrIUkJSWt3xVXI0
XfRxn1l7UejJGghdMF7kOxLRtvfHH6md8Xh6DRDyzUuI/zbg3V0p/EkPeP0qa0gvzi6vQUsm3gco
MoBSqj0m1alLilNZsXFIa8YOGsmfA8UorW1FkyCCRxZyqYVbPncYyfgumjqa3byerf2YLlh1xJNy
13iEJdFxPI/T+aZvzvI4oDjRPG+DQUniLtdOXVDJBu3Jfp2D5EpS1iBCUFcVoPU6QvFgo24ZWNBr
RMTVZTR8mXqcsy1+btNeX+6qKX7Ght873wk2KJw+h3aNgGgaByGpWvkblEqq/AqMhZdmIZuIN88+
e3uyWPd+kepg+lSa+3f4ZeY9UF2VPWCg5IIf+fcz/d6mWATHd0rnAPvw36JPvd3Y+UvVkyr9O4/R
HFGOw5wbFsVgNj6O7qXtq8eVx9OqKdY1CWz+yP73xcmQJCuO90jxgQ5QTL/CduF3ij+RHM9igj53
W0165QNMfPoq/XVwMdu1Sb4rBZsiks8fBSqL/+7oMt4orNd3KEEc+sjdxgUi8LmN+WJmkeqYUg9C
x/FeDT9tQ4x0uUuFalImqAuDJUM5F5TlLdxuNs4xDOUChswRha4/svh9nLAm6KIHizGMy6EjmgcZ
u5q6rZfmg+RnwsLFnMQiXwQLeBcWRJXL/McyC5+QRKb793fkeJ2iwM1IXsEDMwoi3QLahkN9d1Jo
vafMH7PQUwi1wbep5uBwsvOaU+owo7NM1PfmxQ18EJBAGpOONMiWkZBXJf34C2uK1Mxl/+W3rL0w
OzB0DyCICBQnIJ12009/7juQeVjM53vIGUI60Ib1g1+GmKJhro9SB5Kwz4rrpsPRu+2h696iXDcu
wJgjECzqHaoeNqcgUy66NyfZGCYFxPvjJHH3yxTADjwQOZ4aOnji1C6uZbW7PeGiJfphPoUdar6d
SPed8DGdJi0bmsa2q/FJ5QHLL6dEgVce/ZcaawqRt32Sf+aABjrZsqeNgGo/3HyrzfeN+Xr5HvLT
fAFjlAw9vE7DQwgN//xYnfI2j3iIkoaBjelWkj87SnuMOUtnGWS0sR1JdW2B/aJ6E37quRicf8vd
PaniT/TijspQBMAlHzBsydhuqTCsORtqQebZo+J0/jVDgFK54md56rG0JdLdV2h3diNOJ/7HEpjc
z7+7VabobliqRyJOJKaClYbpW/pORHmvcNr1I/9RHDMwfcXr9X9Gea7wtVUeKBkt1k7ZJpHcQmG5
UcCX5aMg6ASqncBc//LtcvzIIR4UsKtOEWPJJfq679LZRNhn93GiPeoR6yz0FcpAlTb0Uw1ZGPfx
aShu39asO6Xoy6IKlap7/o1am7ZD18GqVClRIZ2t9CBQfgWzsqXQEzIcdbHWP1EHs5czsIRUq97Q
YgS1HUwqNcApETFcHyP+C8IeUZUPGYrjvTgxmLPOV1SYd0BpLSZHnH52O+h0O1gjXO8t3gQRZbMR
J5XaSbQh8c1oEA320Bw0NIWqre82pcevCK/6MIkHrDvG1prTej9kay7jwkka8L2AYasFXHv9npj1
rULeYO3C5h+JI/KaJ03m/FGLHhnXU2nUzXlEoChEowFSHFnuuuNeiKvrNxkPAGhXA+apIA6TmZhD
nDDOEtOPn1Oxj7ghWgFpYnsPVPd6yVKYjOOQILsLaD49iKhWi/16wCJmBrXaRpm5b2znxHZ2UC+B
j4OnB2G1kCGAQrOW16yWQpxjdIGLFfpAOtEgtLlukc4BD3pgIyorvxNi7P+ITyZPc2rY8ZGFzr+W
DiAMWPU9IqD9YxO3LUqjCsSUknWwCLhtOKFXWoQoJfSktmhBaTO1pMLsCMlzLpZKpRhfevIngTJL
/AT0+oUNxlfJgmDXXswBFVoFOM4YhP9IqAGYkL9JLu7BPFemlIhPcB4Hz+4yZqpsGjK+9EzZAl2g
rE2O9EtwmT+hTb4V4GfIcncnKxku5F/m3x7YTowV7yr7b2innEbxhrzrS/QAb1WcK+puRe/cwZO5
lkHwLuaXcgPn1tfoJpztVIKy9Z2anSRjKFu05eZR0jla8fwUozSoTb/OVfQYcGBS0WfuQ7AbuV6i
tOl9QIvnQXWjSylAZNoHcMK5/AdiHAqYVivYetZlrK+GZ2lCE/0T4s8+xfpvlq2UtQTPRkz28k+9
gSP703S4//jApQi2akBkyTlaYdZWhDevvKHaBJ34GFVU2G+v3qW9xhSMHd+/42aaWVJnIhYbluNN
V6lQz6nDpjelnLdvRh5oDfOzAElLSwJtWwMZsORC9P7Nvsnd/idy8JxnpZNn5oMCafPMT82TxeCM
VzOtRkJbKx20qHUpvmKxutwvueyNAFS6tDjEYlJaMWmCV40dX9xxhod/8RCwVjuCQXWas6emoNHo
N39doUll9AnJqoUrIIaMj3Mw12IZuo59MGGKXdTGj9rbagc0OBuaqCVBQRQ6P04NdCOVRJzR8MCy
TiXHdxk3oelk26t/HNWlFBPJYpFQkfS6sb+fH3Y+xCQiC6s431UlPk588Mx4pUMI7ouGeRHKaSa1
hPMTQtrrq7PpyFu9W/hO6Lph5/96sDrr/46DuWHK1qtg+S1MuEJTfjjEPUCnFYVyxTwOJY0c7mhm
VCU9Em8zyYpWhwWzAT2E5Ga0IT/MhUgc4ID0LNfk5WHOvnpb3guu1MeuaVCLm77wQ7fDDNJaJgoT
rGbIco/gTFYz95yBP6RvvtLZo0HqTuieEiuxRBtzIXbWcgNzymmhDzS47Z4skgr1SIgKZrYUU6zm
ClObEhRRf4n2TDlZCabcVUc+wIZXOVJrR0nam2kmQfhlWxEiRQXXX7aSwyyXO1ZS50V8LOLncDdQ
REmqGg4Twdve3iIfglP37SaBEnlzXsNinWqWDMhx52/nEsAK61cdi2TRMNzScMjZG59pcCtnYCMe
7WF5WB/iIE3sffLePU6j2lIQMpfnGpa4kU3I4dtOokgvENHTK1SwhPTnNCS2f6ja+ig4xR61QH+d
eIJHmKL3/H/SWO6kibOpYO6wLeqsPJvY0eNNQldLk06Ex72eVpY/uW6UM0XjEYRlJ/3wZSRVwmGw
9f+oSuMETeTnZNSnrmxrcj/JhnAwQrI6pUXQ4LQErlByja/Lw64Ry+9XQtmj7beV6nQGvpe19zoC
eh0b9bTY2iHIYOtcBI26Y4q91XbSpJy6JEIqAVUo6EhMGZvzzeuSpEdTUhKqMuDPH2WFNgOBxjG4
mms08fVlkZMLqjkRKdgPxWbZWbQW/Ipi57qQUn53TPfdRHgPds4gksyhHj3lHEE+GF7LFDQTN+9n
jeNGJHzJ6G8Yjiy6ZzGIyVhUi6MGcQePyf3JoNjo+frD3gGFVwZ9O3BHRWtBE9HoMFER7IUoVHQW
g7MFWUJZRVOKgxMGfUTD6KFtfUsAO0GLdCmTRhhgFdUhPG7xHqi1CdaIdBrmCaZcQBghcGXss3to
Pc3bV6T4vdeNGQcg/EaBXTW+zo0LKZUJG6m2+jYgSi/Qyr/WqQOQPBP3sioccBYdciAcw/kb4UEs
sqhjBa4wqCpJcc3vSZmCLvVQSppMCkKUU8nuRA6QqY5ibOodku7489/vZ8QkrNO5Ci/iTTJjrOyO
KLWMdsjiKMOstNzHkdhdD2QdRLek1c4S160KzUUhdiGzIo9b6+INmVCI62VEpbfz8H6U/gd8GZVU
4Vt4Sl10w2aePoQecqVctx6ctAddahAq5xatRgZBFJH+QUbvy192DmVvgVUmyoqVXZTcuC8MeOuK
yM5nU/DI4reqe7RU2mZmJF0ogbDxENcky0Ni6CKUhC/FWidY5Jl22QpuwJlc82DK/Xa1JKzuyUh/
N00TPx13NUtQnicm+v1lxne9RAgd8XsHc0t2JZ0XTOSfeOGb1nvfPlFkqD7KCI1IL43/Su4Ww0B3
WuUBbRbT0kKg0WseQ6JUOKUf1BcQJx69rz/sgPDdN71yRFRPyIAi3hC3iRikOpCeMbwGoohptlBY
VCXlS3KWx6w2zL/Z1JS7zaTY9DBAE58suBvoIknFeKUlTYmJEwv4fI9kLL/D8jCRCwMrVtTz+Z4e
yGdUnAgQOut0aXrkVFpMwAB6jjiXwOLnO+ww63iI3gg916mOyrE6FUlz8x20TD7EvWBOhFgvU3sm
7/M78TMgXmfdCh0SwzQlQc1wDqCkPvU2ijHGsT5OVVnL7OehtYvf7Yoay1n592CNZ65602VVTNyn
vBeGZM6m1Q9HgzioFdHZiNa8B1gCN9zzjbZx6/LgYaGpHj/j9dI4lGsNDmwKNXDm+1HezCt/HoSR
94CfJnxKs3zj0i4hzSw9Vc3ePrsfm+Sbknm37nbEt3SA6T9JiPru9BNcBEcwPwhUJ/EuyRiWlOp/
V0mJ8MYRXtHucONQBtKYl8plN59TT+2k2bpvFLtO9aXs3ceNFGReo4DQES4YQhdcIffRW5U7BG9O
OzoL/qX2TSRxe+75TfPyringEP/UydZtzk+gXhNBAJdXKbG/leY4ZEGKQIl5RNX6ecCbpnT8IP0W
2Vdths+wlU2opIzfOiIEPOhcXf881n9b8FqCmEF9fMtYPH8USQPZaVR5qKmvNF5W5/8ZWrTh1rNg
ULBWBlU6E3OUrB3FHDYKbrd45Iw4ntOFsHbe+Aiz1Pfggw/Wvf3RD4SRxppetXg8Oeziu4GrPd3L
1IorCGWHfqZ69UOxTijIEe5kYcNf/x0EXNMnGLKj6FRIXcwIpN2nUOGP4cZ59UInlslqJwb5DTW/
7Dr8NPltR44QmsHKu6Elj8OxxkC9GCMwD3CYvjSTulxAi9/wTgpNEbjRGOyybD3ahPcTvc2DbD6f
VjW5Od89IqDzYawDEfd6ZCTdPSgX+xAgCjN0UagTsHrX6GITYDhoeOQKxseN8NOsUusbbS2fYsV+
BOcEMrtVXOAwDlCoF3Lz4iFEKgwD5CqNlZbVMsi60bws1cQPBxMhBAwLyVEU8mkwMWgRctYgIGq7
BbUgoCGJLhrD+DOPSU/qAg4LbiZaaMojqxmPjhbkGh7lNGelcujjGVUDLTx55f+QWrnQ3uleVJ5a
9dyrY4bBLsDzpXGrjlNjoSZ5JFVrmvc+JlHgGNtt4KAaKT3aZ19S5k1PiMaWOPCyVo5gFqk7hru8
DSZdcUxfOyxnClhSA//JerRCv5F9VIhGxYXeqgvqQ1jnjYRmbtyNpxmWoh1qTVVyAJePkE4LgTLR
vQp/u6kbba5QgRoYB+o5Wkn8Uo2YVq6KRb0ol1cse1RUO8h3OcTBZI0de0JZY/cMXur49ecdGfGR
W9jIVUEJ+EH2LjSy3KR2cyAcSan6M9DI0xdtm5ftdoLKJsEmQGUldvaTZIYxD8TQzUf2ZXTrMSem
zyO7QHln++TznbQ0E6kDnHzRUdQxzZBzDmQJ7zctty8TDX+J5ZqcwKWwOe2PySirAkgGQKD69BrV
CTtVg3x63HDDbMWB4Q/tYe9iXqkwGTGXn1KlZAc10weV6eO2cIVUOhWQGBywAzT7nm/10AEy5e8U
vPQeYR6S/A4/CjpDbQ8EtTsoJnk7dy1aO9YXvwRI+nJOFaCtG9Sfok9XsOh6CYurZ/FaVLQnFBlL
kPlIlgyiixpzy3GcoVdW4litui+0byamYkCATB1cOmZZ6vpTtQm5W9lahTdjaVluOjbi+oshaCZB
SE3yL5ho+jsLO32YpJrYaIX1+Tej+mT4h1xVs2xDpKongpZ2pDhHZiXrccEKeRO5NEhdzk1KvsQf
Wn1ISDdac5VMFzmVWdN28dTZ6DnjkEpGyjXmq1CWOO+1ntsRmuB1Y/FknvR9qUNGDkMtxrFo/iWi
UeJQP+KI26TXD+Mro1ksAtxHi0apJuTc8GfsBso1Yt3h1x0k9gQv6K5EJ9Gr3LVGZLenCKuJKt5G
bNL9mzGbJknRlLaKQ2Ff8KuYlMyrVZa0gfdnTeKSAFsjQ0id9TC3S1hpdx/mIIJZP7FXPX0nY7yD
RlFeRiYktH2MfOmD6UOoRjEREM7rQtXySO3OQ2cTXawimD+Xxh6uy91N2vdi97NvHZrWpesiS3Cs
Fq52o0og0ozHJTsfA8OZVprsic4QVDGG1gLcF/lcadBFyscd1wJl7FNRAmaPjC0gvc1JJY01/rX7
sD6mYlVcPvXEKjMu1xBKuuZPP05/FtoDJALN/u8s5VjkCuziV8TNGXo0gpWU94uz16PlFcX2yxpI
Eb5yVmC0OSKdWIz+PxaeZBrb3jSf57GGflsBjGigmabAw1uzWfdV2NbxtsOUxyrSu+RUEE02MVRq
4OByGVnAetH2TqIMajqjvBSzx+jq3xIeHfwWxGeONKzfylHDEZcS+nBW4o40NFoHOJi1R7bnE7Ud
zFG9rve5YcJCcpHTEPcrNqchaE9ypgbmWu4r2ve9MZwablG2ZwQaNJaa0/KPgFosAMwd1+jA6++c
uQsrbPS1xVI3Bb4Cz78U2s51ONhxR+aqmuluSQmzjr42QgGY3HUFJxkKAvcl++enmMwQq3wLgkwb
MCkPDuBh8lQsxnDlBtVh+9HZF2Lp9UxpSWxDifqPzgZD7c4xD9LrkDwecG6W2aytpVWy2kSbOpP5
7fsoObgKbpCibxlfR5jIVV+E9Au4SdvDpqesV36R1QOX/aOwJodQLPNDewBx9w4qiCHEFwajqrQJ
XfvU9H7/LRC97r3/irEFmPkd+3B6ti4Wq+eyzxUhOLbhUaAMeY9B9loT4p0cLfBo/dLfJs3P542p
/BKI1jg4OGKHDfE1lp7ueoHekOqQIbVIfx4BBXMlIF6aUwbGnsK6s+JM3CDUDzwjJXrujBY0WtbP
zKNCDrwXJf2hv4ToaJxlY1eaHQLIpHucdN3lyeQoCEJeI4cavdaWvDH6Ibkn87h+6AITjcOolFkT
f/j5zUTS1b047Xld7774rWo/3CNirA+yyRB8w9eGIj2tKV/zDXef0Kf1uXovqbfwmJeMCdN6x5A5
G/Z3ty+P+ZFP/jdYkaV5i6dGD70OaN4hiD80akkg++WJWPaQhrTeTXFRWx8iSnTrdirS7mcp94kN
qFysJj/4mWeh8WKc8SDhRBXR/EScTT8KFI7bezG1YNx0Rd2/GsEp369MmbHHVNAmBMHKP94tiNPI
r1+JyOoNLUz910u1m2BdxlqGzFQ67+DdMO22SZ42xSUhKbAplli6UdcjJ4GaUOo0Sy2lborIa/0Y
YAOjZtBwe1VL/Mu16/voROQGbzFD8QD/PleAKlKJMiHbdjnQwRSosNP3SEvgnL5y+iLituryemxq
qcXfgs5KO5Ca3cnvTTDVMn5V/MAep4XEY2Az1afOUsXLmFmLvQHoGp4tUzW9dXpO1uwBJuUIvSyP
uzO+BzH3LceyirM2dxmGjm8ioCMWZeyrGJ1AzlehpnGyfXWZ+HHP9RVceawFR+M7ecDvTvPpubbO
kADvx3d6fJDy1/dNM8aj7I7arYT8zuPsfjbrZkzOVplXP2HtGWrP4r2zh93YVivF/hB09XAn+I6Z
0+06mDYBkWF5+niT7L3cRTampay6G2ipxKo21sAB252EV2qWYTDWLCJLwg/lsG/TWCbmJzwu13oF
W4tYQmwHXT42RzWghPc3fcQJeTzYVW15kJMFdSwutc9PyTyeYkHHjRNCk22BRQHGHmnrAeR6eXDo
fNqwK8jvAC0bOBNEe5gMZxvyEgZvekR3m1fbbjUTvKe1biOCVg8/xavN/N6DVALhT5jz42gy7txA
aOWhcAtfd6NvH43+Fu1SEraNSJ6/2Qd6K3YaC9YBwvq6ymtqwJA6uVoUp5dEtQ03UI5waatBZfFo
L404AdtbPgB06YN5Pl27cuuyqiV35dLkRBX4g9u3aX3WImGJ7dxQEB0YxrOjr2hRWhNy8DNOVAYk
Cm51Fvp9EQIGcp4bWtbSng7zNm87cE8boou59L9jqlLOUy03lLPoDIKvu7D/6NjVU+QD2VWz9lXS
BjgrZc0t3uIDB1f9CaPM9PWyGQOnawO3ib/GgJNwBGeNdp1zCqYjSqLWCVyM/SNrE2hzJl7bW3F8
/SXMiaaxhWiNQL44NlbqhHKGNn+sN7E2FEsG+WbxHpybtAyg1p+IBRP+/xExY43drY+YHlgL8yAD
UR/2e7iezAj/4itfBW79+D1MEl+8PWlJ5T33pVpwJcflSJlaEFwDSCxbpVnhR17liQUrm7U+URpK
0qqVXt0/jgjU36LhwIIcdFSKRm0CCW1NQs61hnOogoHtRY7UVa3FEeqCLr+pGlD9cOvOCalTSYf9
ttO7rJkK2MUfq8W/Omqpz2q2J3HAbEznNsyCLJflFdhXbgvsFIH5bw8WPttdkZHkU/nzQmcjKnrW
GsvjfeNisOf7pFW0Qawa0RuY1i/L5mJA7oV5gPaOsOk6F+Rf+bmylRtNkdNFoGjJqjuGRt8JTM+8
YhO8Gl5dcnC2Axl52rFlz41mE4EuiW1W+ibxJfSp+vt+qK2x7JFWy31SFxEuUAcvct3sDKYqwK1U
xeOo5J50u7y0D4S0wBuxAiiFm+osxKyGDm5PHBOKAeH1agFolPnKSLQC4n8mHLzzac4arKCMPmxX
PPQXppG1730B7pe8awppzJLsF0940ffToyH+eyk8wVBmc+uhg1LTTXqp5vtMN+f07rvM3ypLYVcm
WQnjz/M/lpXswoFiyKh76AmO9AyKjVQI4tsYIMAIRijP8tGx279Hig/gzqUbZA1uHl6ASCyq6H8L
G+yhxlvOtvVGAz4Jdqj1+HIlbqHBvpTHtWFbMJJV8TwQl1XZzwL9Su2vsURRUBw5wR25m+Ui70iZ
INxKwA20VmzfGdMsxpHmdjvxVyg8PtVnUKUfloABMICsFqMaGwAuawLmqpHkTKwAssWmpgip6emc
k1EsLQxJAOpW7swvoy5pK64ViXYMWyDa/bgWyLzm2o/O0YtQdxkpU5gWuTwbiBLzBh3ImOG+wLdV
vmxDVM5Sn1IuZyz2Elvs1B7tlhn14FOsn41Vs+8NzFOFg+vGEkxhHcgJk73r5d4BNSWH2UF/ES1k
OmQ49aduLVdFlXXMvQmOpPj41CZ5J0SCnPgPavSNyhkgaICIPkxCJqxU3X+0t/ZhAt9yTbmsiYxV
dT0SLxyCZcBzWTcjzowG7bWI2AQ5l7CYfil5zYefPBphglZ+AEVsgVCcf3Zm7sID5Lv1GW0uknO3
m2gnLkTDFD9opLD8LEs1Cm4tVCoRth+sCo55bPqgOF+NffWMbdU7g9rktyhaFoYStLBOH3NrkyEa
4D2OqlejF51KcMysy6x9OhiG2B0ZXUf2kgfsD8U38DMVF5/iVdjgMG0s2QP2Txr+SY7YgRm+0YdD
UJHJ/ql/q80gqoTsCRIwk6oJwjn96mfobrX7QzoAgFmSBccFV5krwrB4RQZC69KdG5QNZe730t5n
iPI1WPf4S0jAOE6TQpo/rXuLPdHugPnCpDgmXVF3k1CnEyA6KiF4I2rvhuwQ8oR65qfYVMyG+zYS
FkPEC0qu8MXWD5GHIzXas1O5+1Gq/+8Jl3a/R6TU8MOYimnusrFqjZKqwll++XY99WOoM8XrBBCy
Ih9sZTttqi+BZj0KHwUX2L+0uDA03Wefr6So77JefL9r3f8y7dez4Rklq49awrNgnzj5mxbZmD19
AP3HQsfTlU+1d9HzkGXTA28zyGyDnW4WCfPhUDrbBPjmS7IZlOtMjKzUYgKdMM6c3Hkf+nC9/jX7
K4Ga7wmpK3NcEuU8L/Q9VwjZA5BUihSUvXswI/wYbs+OptdiNVytGGZBrhmTn3mxOMZPzEG7tbV0
uwE+d4nlB2SwzST/B/U7rWX6CEYp1D4tCvMONGU7VFmdFN0kYGNSKKKr8lqBHX2Mq7RxOs2Cupls
mU3yxuNMo8hahpUp8sxOLLSRSu5lhuohZntFZmhuciycugJ2+zz1oWFZU22tQG0po9fArfqVjTWY
8qPW6g0DckhykK+kT2SrgtrzagHUOOb/3yzBqOSU82wIgnICtGkvOckPyhHPdZs+1eo6oQgc7K6a
dVfjTEKnindt3VNIkUDzwp6tXHHg5z4lTMlTXcXdSk+2k1znWrIVUxIt+E77fxTJlHHOyht8g2KC
CwbfsBQyJweYbXYM8nQELmTy0Kv3KXnHn1OAh0/vs3ABiuLXx80ig/QZPrJnmnX6HqQ0RDLW7+4w
KZwDaks426JD0BYeF7HVy9c+l3bn0TuBuBTR5xMSi9T20A7Es9esk2oMXSis+qGbR1s9ykOk7BXT
kf+cta3efZ2GkZ+vfRNZAB3w4Fc/PK8q6Qykkr0PxTcl1cJovdjYq0aDopRldzHto+i/TqlRl133
XsFfxdme3lOL4cisduosR4Drv/RQAd6I0K/j1jJy0w2b2AVthS19qxckR0L1K4gNLojXCs2DHdV4
Q2/UeHZnxUU8pZ4Tm/jUhPpJMLDMENneXGe/PKYkrA6lgrlMfqdJOeS+FlXE2+qQ39E9n2aJ6QlC
k3ZipHETDbXYsy9U0aCRdd9oMGG82tRSS+fOmzY6LU8DvDFBnTHrs80Kxn6FDD9PFgbLXxypbped
Pbe9LFYCvhROKGGIBLU3+O8ILAa5jgNPhbm3YjwD+CH6CpYF3ZYd2GweLE32mQTN0buZnAotxVMG
0WYi8gjTsx/dojaPfE5+ENDhTkLvhG3SP+LbMsu53ZDaN9KzhK0GI1t9INJ7L8FIXhbT0HSw0UrR
0Eq5fg79XkVCOMOJoshc1PwMdqQvd6KKDGhH+73NxXJJXHrsAdWXLmYzX5t8frCtxCcYkH7Wj6WU
7FGhvYiFroKKCdTp3sOMqd3kn8bcLt+dHF0QADPV0Qat1/7F0FAgc5ln3Hj8MW4Fai8PQo75d+1t
gyWr+uiAZrYqoDQt2kd4ooUTmAlbyF46+HS1aCHRvcBMNhsZCklcWRMrkJnjl/kRfyj5GfkJgvmE
N1EH/EJQFyRkiGoWXSHUFBi29P/6VLqa55v7SK55VsKOKadke2GHowrFqrEVseYAnpY2bQb7x1Gx
rTLCYpPMGGqg+2OC2BqtaUb9lu96DdDZka0kM4I/VJPzc5BRK4E0ptqhHtI9iybkgknUaQd7LRwd
w4pcb1VgdZ4JFMz0jgU/vvymvaniknM29yZRpjeW3DLSvZZrmeM4+6ox6q0dU7AUvsjG+ddoNshs
5WmBJye/kTIV9lSsI+c5YZ9qZUfJxcntz/U4HZDGQx+FXej6rmLE6Au+6pz/RVd8Al2GES93uHfS
D9Ln/pZjB9W2gd9dwIoL2pN88+H/Cd8NWCzhLPrqZFtPruLVxNLopMvWuSSMo+2PF83k8o+Wbn3h
uVpiomasYjSf/r5qMXp3Wq2hhrW6wiwmiM3Wk0YF3k5K7l+F+5n6GHfOg6pd9/Tj4ODNHKeQDmJ/
1PoV9UrL2/zr0rFyEawUrWUf344Z20VOt5p5zWrtQvDNJpCWOtzIZ/q0Qd7OodsIILwDj5w2kIud
QG9AP9v2G50zNwG7jSOXhe7J/+mCf6k/obtOE0V6kJqemOEDYDALlbdQ2yQUHdN8dkXj0HvmmPc6
rIPiBHy1ikBkvuyWIDqtFhaDP+s2ieEHiLXeSBXl8hrNbWq6X9AN6x3CzvY6UMMvzGZNc9rnDR43
eeaYt1FnvmZiFXNrnfZPZ83ILVvNc76ecTiLZy+q0pwoEyJXeTJUftuo1zVqf5XfNodHKdCFjBLS
36CXkr5CRU8giOzn0IUHGqpzQ+c3pksViDeMxacp9rcx6TijC79HKIKY1q2Bp9+vwX3fpEKIbmGg
dx9YebWg0Vx+st3H8bWDijOegfDs46aLbfPtPHrRkP3Bsgrm9TUD/9SoehaV8jwMsgV1v3YPPia5
9wX3dfcaDG3xStXrGFoa/akd7vofrjLrCW4nMQXoPNaeFOhapdIv6Pj2u8VxD9GSPOWtrmehYVS4
JXS0rnalEwwcOz2EnJvCxwEaF1L8hi+5X4dpHpADWVryTpmnz1uv2/8IBSXjsYoPlq+rfxBSHmBi
Cd5DZL8OZphcCr9HnsN5BB/K3XsYVd2/p/EB16vU+1tRFOrKSopfYDhTYZrbETDMZ6/DFQIhQ4Zv
f1sYlL8SYKlzN37OHIVS+RE/2cxH3mQJXUT9frXtR1ZnMsBicE5tudAzKY8x07Ubh7hpYUcIjnE0
OmdHuVsia/W//tLp1X7BWLFOLDzDC5dk24BNbvMIcLS67SynUnFw4SiecpeYvpp9cG3T8ZcGLsq3
vZAwS3HvR642l1guoLb2SEZlR3Z2ZJ2M+RejAl0lfDz341ByyUsUBsmm8f6D5sYH/iv/5QsPRzVy
C124PhK8HHofkdhtJrBHoSxHuIlM05m2OCcz4uPPc2CTHaeWVq8yDb5GkxyYVxmTd3YM8SMm0jD/
j1yt6HCsgrMByc/slZcWYZWmEZToTq5YDNMweWQ6oYwA6xhjq91DIaU0ygNn1omQanHvdPk8S4A2
r8F8cdwmg8ZwRYNLKZqvxxidaDuu7sx00bRlYRoco8GDHemda494y/6jR6CRSCMAHeHUmqBs6WjM
VePJWHg7qCTH9MhnNB+M8E6k6fbIVo0JVjjEpgNsjyWjGO1Zybf2n0+9AsE+mso2WdbRYO/GrU9r
2DEEh2VW9rElnIouTjWXuQVXAg2PvAozByEks8+2Z4qWkp7g+eHENbhMu7lUiZ6AaowuTUBFg0Xi
mVLaW6RaMqAdhC4fR6v99GW2S8oss9joDV4eEEJY2YbRDCeVIa9bXfyo/6o/KHWM3FA+uN3I4o3h
nBlMFYj/Sq90YR8ChETnZBYoY0w52J4Spp7qGsAPOcO6jrJGngx/akrHDTo7MW/wR6KDEpZgxGXf
4SYTkOUicItaH90Op9unje+9gY88XLJl7nWrOAiWRJFs0eDvgJhYvE5yUSAb41HusSZj4cwi8sjm
Vu9wKZEDbMU7AghdO3EL5cKtkrYT4UTsP3StrxkuhIGSyJqjEx1U4gEvmug0dOJ5qegqt6Oql9M1
h5bgnGIQb6e8K4CcSE1CpZT6hEJaNO16JHpFUJYUvky5+CneAkdas+b8pIKncgcdDxlAyoxpxysi
yv3HI8mZT8ml4m0jin+vK5H53S1eHgGg/xaFV2bdOYEtBt7M/fH7c/zw1g0aojLdD6hgkiC5R8X8
AICykOt521sx0zvmJjPLJt+T65SF6Vb4Iy9Vrekrvs96Wy9lqDkqsP++sAryMdez51nhnDGH5Q8F
2Z1BMV2Kf3WVdxc4fjSWxBGcpfFwjAXmrg3rHSY0RjpV+mAAN2DzRzbOFSfqsL7aHNQGxLCsR0ch
I3Wh+ydiimb900j0AlGz4m4YlZbNduHBy/0xGuHAd03vMCM8iBDiHPa9+DlmFeCAgaugC9hseSmV
m48fTxDWec+18h7cSE5fzH5sAZGA2bkkUqNThH/syfi68VbrWeZxu0+V28V2gRtYmIT7OhW9EIG9
zzbD1egA/BbnF0CrCsOlNtnqFu537/5pzOyGdPOZriZ5TfMxsgloRdWbMODrwKrNOTcXOpG0Bjgf
k9PakvAtA1J2B4JgNkeDK8ogZT1ENBUD29vL2cH6CKD5rL98DypkmX2ym5GtFfW83QiehtK19S8b
rlZUezPXmCNul9Dkej44mDq8USvUUBp8slD4gd75Pe5rSNgHbJGoimit0/AioW2nZDGoi51XbqBs
oXtuto9JlcsaCzHE/SzocgQlUq5FmSW5A/W+YrSg0fq8P7aHT81cHBN/kA4v0IrC1f9NC/dmNyf7
JlQ/FSlFFwLm7rbfKsO9sgSGcHUqPba+j/CPKzEJzixaiYbKLxUlYhu53qXtg2CTAljYJqlE1q5m
8EgemXgWrbkjSwIw2MGHmbUlh28A+tr3bDvIFUnWumHOZd1ckISjk4rAVglc301rn/+8JLeXU3Wo
42L0Nz8YlQc96tEPv9qALBAp/So/GyoKkqgY2u74N7henu6veA6b1kQaWT77gQJdN9/FpPworL7D
qSPflR+Js8Eg38bAwsGHj5gZAjgY50r1pzCGM9gtlW3/iq5YftomnXcGW4D89ELEKmcGnM4+F9Sx
K/QdwO4bUBdq8gP8xcFrBcu2b+BxMJ5ql4HLV0/GJpa9MlMQyzeidxCq+/i8ZzY+vv2tdSt3LL+9
42NbHg7aVUtSC7CRTTUol2dwZIu27AbZsSUNXukFmTNiTEYUrcBxin9VthkNwN8lUbB3os1Dti+r
vW4wEnFKImXuSGrWJ9S7cPTLpDh0ic9r2EHDBxQjoWquHnvWwAVKeCzqkiZ/Eo/jGsm5pkfdrZSP
Tvf0AI9tVZGOVaOvVOpHthbzTE47C2ARsp6V4I9P0FP5ixEl1qIiWyaaE/S1TixI5gDM09ANu7vx
muAKOjcZeP67wALH7ZzXHqqRSjgqPprcbLMTSUfHZCz0y7CcYWhZYj/bZ7ZM+7avge2Yq/CCLZEc
8tmpjy66xIL7dbK9UBWmzdnVOuy5iQc9K6lH3tE7ZzzDoD0RV+ST8/2XQqttpBGFIKlnv90FHLdy
0klDdX4K7i4AP+Jq2GKcl0pvfOwrr9koqQucql8Ou6lti0Yw7BLy3zPBRP1LXxYuUco0DWieV4N5
rIYPQL9P/9axDWf3CEq/dm2oNTkO8OV54jpfrRZxOepkKJdIZUlYbHYCm7j472bncl1d3Rd9jMHS
+sj+8EnuHntOnT21n2QtX+1ThJRUxnPtObSPDjrK5AcNzlZ1RSxqRav9Q55KAbs46LOPRozonHPQ
ThJfMHNn8mswuXtRIjF4YDcLsyk+WjQCrwdmjay/BOhNwdnKeqT9H9B5GAEl428Hy3zPLjSgop9e
xBDhGkIRWjlvFDWLO1/Dcr2gCefSyyxEKvAvDdlSAY+A26j3XMYwXZwelHHIy0q1oS31yc5/dgvx
Voz4dIZbcTsHsm8/eA53nBo2XsJYICTWM3ewhGmu7rx94gE+Bzgt445Uyqc/KqFowZSF1JOir5Kb
hI/jHJPwrXXzhlCl4CEJ/w4BGajah2ee/zcLB1O+rFyzn5Oxmrz3t3WgtlYVrDDu8zNlrVfhtPbu
x+cQnW+vUU3mvvkktDhblbEYJXNMw7qrnvTWGV7lHiQprUM2t67nyDjQcu46kM348NxIghIs8Of5
xjh04Xb6xZNtcQHrpFeO/KNdEVuyzoxfmOIibzpe1WnlSxHpJhNErMUjYnGlviwlI/KdpvkSNiV2
6Lsn88xgodqtQMhk7D0Lr5jKllRkO1VR7e5kpzYDSxBCNjfckXRWQ7bhXmvL/dt25vgKbKEmdcAV
7kyNQ+fGQtaa1V1W0AhH834bQvGZiYpjnE7NRqpRj5V7B7l2H9PYATbOr6GfontIhptVH5VjHSqw
NUu+U/+J/Kpz1iW6XvR+jpCYqkctEDiqfyQh+KAqa5qvSoIRjs5aZBSvERD5ub5Z/qwDtepp69Q2
mAZNkOBZX121lZWT7W88gT37yNhxwMBaqMkTr/l/yAW8/I59JqkF9hRO0JCZ/IAOsoRKqsawnggw
LpwDdSpznhQae7pFuA6DdFeedQf0RbnObP3rqvKLVyaXJlTG1M3BqW4r3+A+6kNOIxiGyMF15xhh
fTY1O/w3pHTktitZhjVR6y5oDSCdFodC37oTtLKA7oxBnfnpbduYQ9BH33d93zuj72CBfn2odE+6
hZmD/V8qIb5SmFe/EZud1Wgb1Y7LF232DAdpK+495nJvRd2Q0q4aZ+mJ2blGNRUMWpCiLFBU5HF2
jZu3NGifdeyRU7gse0oWEun5F7+1OPGBeXxcnXS9nobNz5hNBoOJSoQGYI76zefgGZyuwx8gwVfk
uBttVCMCrklWLwa1R+4LatL0W7Yf9RbeHsg4NJ9eesQm2WeYFRtgBhT5ngIrVooNAs3sDyDlXd96
j9MbwIBFq5n+uEYEPIDRqgoiZfVR/uTL8rBb+BfGExZwA7S2d8bBDd20uTiumVfdNMc/XW0nAG0X
mDKPhj4WY2/iGCIuzMZ1LAt4buarp4kvMC0hFPuBR7xU07aWbb3SEiHsUIQhwhVA17xvIHLFNZPA
oYMtoFJ0pcjMZtBNqSjAfw73WJFpC+canZ7XaLqYwwrGKv4krWLM20tBIcdsL+7Hli5Q0lF1NN8t
uAQr6VNygZjvsXoqsmuRfMj9+UPqDuoUhomAKV6Rpepz+IHdlY7G1H8fWSE3UyIxD8QImDWdk0Sd
VZkVS0lCAcx7oiLowR9mAWGxzDXcJj9M5TAJvqQXhlOG/tYNmLA5WIUwaQcpqwnPR04SBu88sEjX
WruuCyrbRy4EuuNmwtLCv5m+IcAcaT5SZI4Kf46ndApOosYX8Be2922uIrMhJiT4jSYj8tmW1vLs
+qevXv5W5gNGGpBYrVIpnfxWwE4yoIs0iz0W5zSAXJNNs3GqBdNpxwUAiVdiIHOf6DIyB+s7gQmW
Q/RTLhKUKtw0UEAIO7PJks/GxD2KxeWL3oM5dY6T4j/WSTiKW1/cJ9ldNWzYWRSNC7SDYUC7NkpP
TECuMoK4J8NQh3c+jho+5umearVTjDW91iYcplzYR4NYf/T2F9/Ups8h1qxQI+hCRQUa4yEOcXXo
poX0zQf6GIFx+XjDVJdOpo0+plDkHRKcfQOV3aCpu94xQl2ZNZnNagdFB+na2Q1vkl6Sq/z8M0cI
5e0s59SG2uHoif8/X/3C+J7oHjEsFA1+Uqk8Bn85Ejp9oV4xuRFXxudH/HCU9TYZ/LQnDe50/Bha
1cSu4biyYEb5ymYxetL7sTFFdeTjRW+EsvjXNgv5la7bXl1DhU4oxYgyk/th5tZfyd/VzkRnWWax
sO0FK807yciMoUr0mwMY25XL8MjH5cVgIckFOTGVrwdprOI1NHmM5fcrB6Qh9WnV3s3EYEg4VNit
sIdxoEhGj8EGwePb2wDRpSaKJOei50gLfZ7Dq3zyFK+7KHLfMimNgUug4YOragHA53PnlljVHPGF
3Cnd61M/rPr4RP8G/rP5VWqOwijCmpxvwm2ZxMslDXz+OAyZE+x6YpRn7nolwvdbgG+LYoOpeLWc
UYX7jtA19bS2Sj4UwLUb/o4bbV6iGIOjRfpY4aRCZI4RQgK7ROADK5MNODjkUQ9iPM5zA4ekAXlN
LqXk95/V1+OIBDfVkGR9836KYdQTAwL7Rpt06qPndeOWgwHLeZQa6fWotW2Dzgq+C7ZmeJpj7iGS
VSJZPRKOYRbvA5do+jz6iwkmW0zYAIp8vZ/5L/KZ93wDGGILfOGdv/gkm5hj5DC3j8WR0iRiBZQy
ZDPR44be4A6/FWy/25p/TPJKvyHnE1g5E9Xit+dC3P7PpktsJhqkVpJxnJV0Q8eVsRfIpQuwzPkc
hTROTA2NOn+AtyyLih4O29dJR086+59NmXza3dImA9nM7LCUYezhqHjyB2hQ7uwJMVWA+jcR+1K7
R85OKoLbff382CBjVDxpvhdLwBvAh6aRum1P46kidT9nxXQRJpwQIRVUELcbYi98/LckXzLFI18K
Bk5kZ1Q6pUGpAY5MCrf2UttsvLvR/moxJd3q2exdB9wcgSGUxbQ/EEI9awnTKHZ4ntqhpeyBhLm4
6hlpHRVUVD79CpEpUREn3+pYyTczZh1Pcu7Z0NHeJAsH0FyxW4aI28Y+P0qdnEvryN2ez3AduTqD
E1c+xVsiGA9Efy5TewR5dsiFkJ9MYl37M3GY9o8aHJ9DsR3M+MIhUXtCKBg78hP2YNHYBSIFjJt8
GpiKlsqXYcZndAMgDjOLWUlmLh4ul3azfvdQRwXox96Q5ENlb4OdzmAW4NYgrsGZ2M0wUL+/j1O9
K3lTka5RqCdwoZR1HPPxlYI1VJLeQs2aN3ShGYWo/Jigzpb93lKFeqTj9ScEBKziRGxf7b3NH8lr
ZD1RCPa7Jfa7wlvdpQv9wtb+s59zoC+uBBXj51DDReSpkD3kFGVHPVT1TC32CAl60KX8R9soUIUA
LGUJu5MY+O/hyEmUrH+5w8Xg1nBjq9h6nYzEppkYR/OFEfUjzBbMpnETVMeG7EXT1DPrONCI6IBl
T5A3cjd57TDFj2H1mbjucDBrgK5LcDcTJs7vorViCVt1yYpGfZIYDbtiC/4GORL2fpXBtYmbHHsU
r0wY8tMGIkHSMxcGGwjbIMXtUvzq3RoOWgbNl5YUVLJfGNVDH+Qxg7Qar0vJo2nOgzK1id3iWNd2
PQ0gwYAUIZP2u4R4CQR24XusavIH6G7ymivGPATS7ylYxVJ2dJy3b6BBM/AYGUEQgQtiuOuiqxS9
0UwuO3PMArdXkxtCUskSpPTYWgH05Io8pXfW5yiLzT1CZPUDJGj010yAuZzNE4F4aXBxEyH0aP3e
wke/DmWpmSDbieKeqUXNPYD02N8gPAtHQzA9wyIr8xfKIWhuZKwwVSCb42GF3BZLWrsIHKkyTU+F
VFBSLM2mpBnrlIuQ3DQ7gIOjvVehHgjc+bbb1VUZoEEXIkIDnTSMZV2yrVrR1e4wR2hmWRUkVRzQ
29ToejOPsx+IUGFwFPOkVwftqkoWPtJDXwsGcOVUS/OxsfUvRmljFZSYkLAjIm7oT15wVA9acCNO
18PX1LZthXg0HEu9dzBGCx274WwgU1D2JiqF6mNpb6zDYWsWcyLGqsctKSrCF1zMGLrveeb4yrwJ
k4n1Y9CxWxXPN3YbBQ6V1vFKbwm+S98KFEvFTgAWXKLJekcPrm+vzJHyLzs2sWhYwzZBCr7uVqxL
M39sjr6qZcCICOO/74Nb3hvqfcw++MepeCMIYYaGu7Jx8Q742tGGGnn5k1hxSCWUy2r6BZ5+L24u
zM0HbQ4GirG3JBrYwwPQRzc9fLRAN+Pb+LxbZLnttrT66nKtxK20FFAO3q3gX/MwoZ+kESpitEjT
aaXeTxWroOfNmOUBVIaXXgDDp/49QxnKrmuQr94wsBC0Hj6TN1rBBf7NU8bSj7tkMiGISCwg97SU
8bfOkZeeAzljmrTjNSsSstcEjOHH0v1gT3ElpwAYYyWToA5XSyvOiWrjC4kdaESWyzi79qd/Q77I
KePnXFQQLfFqbUjEaTA48kyShEIkILZXeTne12IePQD273uqJbU2Dh2T0swaKUbZMDWFv8MT9rqm
rQHMYNL6s+w1SBuCBpttrd/V275l2hF+PjTC+HPfa0JVEaaTonaBRPzErp6y74h7oNh0fHE++1+G
Xuyxc1+rnnx6PIQ0Bew6DMhav8QHqKsNcK43yax86TtQO+AdnqnvazurNcOWetEjEyHVdydKWufg
bEJBZSTqn5cyLWGVOoNN1nUjGA0rQZpOpBuDHnS1Jwx/DWl+lOH3OzJJkl9DNtQ13/0kCTs8bSLk
Bxm+QHnPmFdWMv6lqy25eUi+gPc231VMWiXgk3dWNEtW1JkjqbfvOeUxbAN5iCTa/sjQK4FL1V+9
OXYw4g2xwZ93vkmFLKHUexpqa9oWWTJMMRFsPQeIoMUjTr5P3P4x7BTz5D3MIDnk9ieayxeIA+Rs
KZPsHSqKzl+oJRjdF82CUK5KE73iFsJWgPwHfpwd95ugFZQnwuLBTL8e/yCXgh/od7LbvPsJ2hBf
m54lrIVUp+GfT04ZBuNLrXjDla1uTKe2DWFkyAPGT4c/adviJ291N3oMOR7wtvMr8TZdWE57dwr+
q58pLPA3gHKXS2AfPX0Jl9rUA4O9ouW45s8CT+M8fBYcWWqzpdaW62WK3yYSNz2x2JA0X1PJmhT8
w6f8/LG6jHNwWeX92ZZcOtxQUFxMtAQNiIwdtud1LUsJExcm3q4RIIP7sgKPAjamDpVg/WuSG4ng
bukPkiOzbYWbqaKzzgkfZy8vAXAiNpr6FKblsFjxRIZ5Yo3GoXXcs5GbEOw1wenVYrt+KmCY0VNo
T3lxxa/AAk8KP0VtOb0nYGT04LTJq3vpRxFxvjn6SY1d1q3s2F9I97t7zAIj2+AGLssL3sg3dLO7
p5u9uSVOe6BpiaAr+PEcVnKlU8/QuSQrNPjEn410Ry2Lwy65mgI6ZJwkJ+MGP/z2GaxydxTTJ4yl
vW2uDZsJb8UxxF/0eUzGqis04joE36oNk+saZPSjQ9pIB7dnjHMzhkxzPik53cLJzfVEuzZpYrjM
aVIz8v2ArySbW1mZ++eMVvxyERZE9jmC2HLdLEfmjdT8FBqYAKTNLt9qV0lQ+LDqFa5Zzpw+MzQM
GzuFbv7Bk0vetJwfcYRNlKKrYip4eS5rqgOSHOP0cyQ8zR/s3WbFgAnM3PPe0fUOX53p7X/Fa2wK
dQ2QDdxQnx+VM4ax79oQkrkkJ8VoyGs9ZrrSGldVnEXiUS9TpWu1+OMI6WiUNrjlZWY3rO83iToC
kuGWly6F+FjW+1JDN4fYTHheYEeABoqijWazTZ763rFv3cuCO1Z69iH+I9VAx1Vopt0OQR0KrOjy
0vzXE3LV0CgvdaIo/bOfuZ3S9B4KcOmJKU6Sev1XfUkrg6aMivRAQgUpyj8P9UlpO1dLwGOM0VNf
IlP01T7zBwJ+hhre8ake9jGCx3xOXvQLM3RMvm8lkgSHgXjLilkF/Ngef9W7dH/D5KkGNt1nAhQa
VncRcdEoCor6gqfXMvfmB1o2P1H4PhfNSeR/h3GFE6wWuvJP01SZT8YR+NJCQYSLow+t6Ppzd6eT
Dd13X4eABNqWbQDkmzPkn7qVkoiLd/UvXg53WaeCc4S1eMy/JJ7nUFowijYTTXoMzwUJySobRXRA
BB8WR/CzDvNfr+ewTzbfXM7ghVlFzgAXei0N7nPZ5ans1x13TZMX9md4lsJkiStkYbHRFNMW3qd8
CIpp0J2IVXexHR+vXrUoOqxoX2retthmExT4vKn51E6s7OLVE+DgFuxw9cT+4f/yy7TGG7w50vEG
t2rxmvrEaE8zHzdGRhTo2ZEyEbdNp0h1zGtFwuXzr3UMqXtwkv/L/QRhFyZsGsRbwBG9scs4Brrh
gluUsaAFjco13tR29v+lZzJGZUsDDpIJtBNYgA1BFy+K4yGHZw5cwG76Pia4ZbLDXckfLxU4h0P3
ncHVpEG7cWowBRAF5r2rCWxoIv2N9kdTreSCXM+2bPwe4k1Wks34KzpqctPXsmhWGTObwnMbPyHE
cngDQortCq/D7PXWCCiKau62ZBifMOPaEX/arLccXBodaDOsRBJ0vB9QwHnSQfkXG+8FbMoCfvQM
5+iTgrv6l0mYyXPGTbEeTIKIqjS+R3HEN/VmvwwK8JqeUbwMd3gq/PH3xE2xSw6zHckuWOPfevZq
YvpoH67HaR8GBf784Bgjw1NjsbFwSeb7YWZpWTkWIyI+oD6Ji8FatddO4M8lPx3qr2N1UsO8cO1b
lXqMrWHtH5B/DvVa8fEZCtqoc3Z+0lUkREpz1dcxBJbk3hoVlmpWfdQ5nsnMmGHQnaEwS0TIThV0
CmistaqZy2hgV5PYJwOts2wwWyRgk7ce0blKvTvFlaWapMFXO+6y5X9Di5Lf8JzfMO5IdZmMZhw1
PTugFB8GT6kwT3W0UAl8Qux0jCXbnZlz5COvKBjbCDoiw7S9wnMx/Ie63ikQkVmKWeDmc7QYqfOj
aN0cm29iFhljy2UhBIWoa2pYL8fSrZaPGoLvL3RAD9xqxjNfH1uUMAiVl1P4dveb4haWMbhN8JbP
swlBBpFEb9xioiAOwcqIBwaE5qd2wexGo3bqNSm7767fYhOjFg1wqUyU5Jivx91mRz/j07VfoAdM
Jc7Mt6EipRKxIcHJ99PCBnOpUMqIiTE4ghs0+0q4iJVW0qwvJ9jCQGu0aOeoZHcOVa/XQxPqDcfU
Gu32JPg4kWjrOGJFk734+RkJduY/IH2oCaCHkxmZbfPyFZ6A/n/IAxFPH/48UWg263vSBKmxG2uK
xp+28l0mfG6KE4O81f9ZnRU4jiQpmXzPr/CJKclMIbCWK5f7Lkrz/GEP67SMPQjFm/V6neyXXasd
xJdB1Ok7pG/x7sYaVg/+XOQU5ILk0+9y9YTSXEpPlMFQJSM+vLhp7HXq5J2f2XUwwpf1w1xhvrwx
039avfjufNhAcJAAGX1cuFuzQEqLMIL2x6nRJfA3//x2cPmG3Qv9G7TZphcJK1cVAHzvJJW6N+Or
23NPr13s89r4DmX1sIRw1/K11jC9mwAghUdeoQwO7QeLSB+L+zzyTiMrvUhZ08Tl13LVvcQU2RP2
BRQvfD+q+cNEfUm1xVqbHP/0YkaZncegscs/AuH5nyJKHqaWBzJ8TqnsJGj4Lzubmbxf/4IC4gR7
d7TysDjRQecVQg5LDeL00ZIUIsT+MwKVq90hDeQh59Cs8FFO1om5sQVTF0cW8CxKZCKbnEVYPBTU
JwSvQ+0uCi2YTwXYgRptyUoP2f3An3QT/H8ibPrpslu1xo6lHiwFY6jP15oAYDjq4vFQy6w4/4I2
mRENTZZkqc4jrmpXo59vb0ZRINjFT/FjZs7TD9sTu8VFuHBRkmNb6lRGcN6GsH9JtVa7I73PVAox
DDKIBhNgWlcxcYZitr2omiUFpNt/NG7vW0683ohqMSEQAIvDwqn66VsSv/PPHXD/LY1l0lnk2iaJ
erAPExYHE1W0PsfFMCC/Ij/ON8KbT6+wrPxlrOWzBysITXStKZbavz6ZIMkP9N7o0jneT/ox4KQg
iCdGM/MFvVaKbKEX/3jS22XIwRneQMp4O0DqvzWuRcf1hqVjzupXOYGYad6ozSmTK1pwHKFoFuPk
O2aNIddepZThNnnrBUx0g0BNeQvmsYjaj3DLVZg+fPMF7tu2OiKHdBOFGpOKIg/HnnfAxSKCEvrx
iP3wHTB37pYTBhL225myGTMKnNFFeSX+DZuFi2FGxuqv4fGjSqHQ0zQOtFLezjnlE97slaOrOtTP
tP//a80jtAo2lve5iCIHwJr+tis0HR5ELDef0tsuXdU6t4y7CyTHatqqNkdgOJCaYvS39FDkEtWX
4fgp3QgUMKNhtU99pdBhIgdUUQ4skS5mQj0YyuVQ6fcDw4MYIqSmzy3wSRt1k6wHMr73c5GHfVMU
Iq3vAUR5oYNdwgVPAy0sm6nKTWHAhY781DR7DE9DUR8W8urrFFrZD7SRGyqYBW1Nu5sjMiBejsQK
yfUq4YN34di+la20FwZTGKKhmMdbl30xzYKLLUs6wKMfrjZs7SU1wdjoq/+BpSUJNS+TB/YdDogz
EFrJye+4o294ThNIWkFrHtXiyl+rhzABjwvXqY+iUWr88QXW1vjoLz6vj3/8+gjQZki+NRDxu01K
5Q1BEg3uBcdBJS1W9kgIpSgcNctN9r6AWRZGzTg2vn0WIueFagX2dUMtq+lMDCx9/9u+XpvY7/Qc
BGd3KQhfn5WgVvl9fG4tBbzRVJN+YRhJ3TE9K9JvS7/pv2mQbYK82PxJgmU8CPR4pHN210PTYLEG
1R3e0OyN3tayEQpnmSBc/tVSHHmGHAyTeEh108QoWWVZmFniFmJ/w33u4FNd37hAWW02q1I9mhS5
zQxiF9raXrSzHSZbQLvyjh+mcppT9CTZaSQffz2BGw1dStsjyUxOzE+t6wokZfeNFgbC4v18shz0
K16TKL49d8MUk1Aqh3s+iVXIu659ABDkJnMKDhwa0l7tQ/8hMmWA1czfHMu3Ij9Y1x7W/BHu4KYv
b9QdGw+rzBHidqMDwe/xPT0kUx94+ovAJxpYGeS7ZgjK5gkuF7bRMoLSYITsnVaJemJJ+zl2jQ06
Zv01HXTYBhbVxhceaTWAZ2vGSxeJNKMDu02Pp7PVOWBnDW0aLQC/wh4EKMwUykBJwkGGT7zK/XKO
ZMMSQ9OWyCryelP8Hkbllymm5wt9MDrAW5+YKKCTCUr+ZM4vKRDdOl//m43VUUNfGIeFqkwWw2Og
T/uNLmFU7IzRQKFLl9QCUPQAXiWACOqt7mbvOgzApSPerDTv1Aq6yGZIrUXJyE5Bg8+9xTn6CvPn
kYiMDvgLifiYOSHIcP9sJ5jh+XhuxesCfJO/5QRvzb16Y2NUZgrqr9RmBmLH9AF6d3jU03sUML3k
H9jyBXEXnf4h/h79schcK6JzzbZ3qaUlCwigwJE9TLPHv2yFlb1WSrfcn4uUMnNScNQNtZEQ/F+8
n/vLvvrdPVQ+YkGfdoB8dSpSMgx52ql7yn7d2rXgbj2HAkTV76yFs//gJHDLxTel4mAKFg6z29Lg
6wzc/d+SIdnEkSNNEjriga7weN5/t8tZFEWk71te8fG+1y0brBe8gwAESiDMYRJicAD+htqpneKH
moK5oMugqvTyheVEzBamDSiLMVAb/vVxkCTKpzKE+QoxOjHcaHDYU+UiyK/rJoQqP66n1jefgnTj
drcmTOkoxvrzdpONMcNIErtEWKRmaJuRv0WGVSnOJznd2XH10Y4X6uM7HQhd9CyRTTYZEoO++ao3
f2P+NtZFaqG/oPzr62BZS3OLh50En9coa4K+OA1IALO9SlVc0cNSJAcJ9mFi+/AcGBxN20wxMK8H
1/sspIKOomRUlzuLlGNGiLoFlAYOjSWjjT8qjl+Muqj6WhY5pwEWebJ+F0YeaBz6PqTWonk728Rh
5Swq+N56tG8R+FhUvlNr/hNxUpAKcWt2fpUEyTDiwDCd4lpQrAMJ0kqBQ8bDHmcEW4pE29bw1cEu
Jn7ytaapMA3y/G+fqVlaNLaCPz9CozcFjULr1EUDP2daJjDstvM4Se+7OmAPxp+c+HE3UghwrIBv
VykhTmAEmcnhS+qTyxkVAuXbr4IwZSVqT3QIAzHJKZI4zf5eL50TTvWMPVm1h/vV8yw4PK+go60k
+JFAiUWw4+OVDn8GoELGIdJlGVW/87hoS67MiarMXfeJF5NkDbcKZ2nf9Kk+zrLsJit8K227mQdZ
uFejMjFEgj9CefwuRmGyX4VaLvAeHCndbgmD5JvjYXZ44WDGm7S52FpqOsqkQt/hEt1IelDA8Ltz
0jjoP4CdvLKQZRbycb35JEl/ApRFYRUAVIsUS3cwsxHqwEDJnQfUhQmviOyJpLjL2XPBriW9Fnt9
tRFtbWz+a9FdgASAUvIAWBWC6YrRrj7kyAI2LgZiMUwQExjCgC5NBpnKhqBKkkrzaOBUwrG1bDUk
gdwU68zQyWZEvhpBG0G+hHb2DgrG0xABMAUk15ryWsoyQUL5RN/Zr0uWb8PLXo0GSztDWFmqRqTv
ClVyccvYBa7OysrQ8NfAQDYNTHxmNg5plcYrEMOQ+aGXbgRaH/lPEvH0WW/Lti1ZP7ZVZhlrxNlt
LVC3P7X70iu7+o6aeBipJLFtymqx/jU+MchbJRtgNlhb9QmOoKBcXo0FegI+RgGAwUGTsV7ocpM+
bNEG71FI7pdpXq75SnESmOaX5C+Add4lEzm3qurYYAgHIgzttQvbsQE78E4Vw+9l+31CcLGkJrrT
jWQAAoz8EPb9h5Mb3ovVawDULK5WQv8ZtI8woIbhoehalN3wIG3cSB2EwzTIWOqzTUtSxJkeFptX
U1tkuwrusga9AO4MPFcJAi3OxYIPnC4z2Ad6uTOoX3VZ6SstSM+yFAVM6t/YHej3aU+xwd34Lc+4
B8ekd2rQfdNAaaD+rhzGmqSzBENJ+K4lNwMrgWjU5ugPQwXSPHoZhfv70AikhMd4mz7oUAdta3if
ScWLSUn0dRNgGE/4PbItpmDaaxOWv5sClFALqLtdpw8Zy/y5MxgRB4OIdYakytGsohjIoTtaW8wK
BzbpRr80bHzfnxATKXmATQTFcb7UW7Cmfi/CJIqmmQg5OfL66Rpvd6c/rYUNcNBOY3JhZDzRlPiO
OnVOvyXuOut5IuoHzRkSGmTT0vvJacbq7Z+CzrbU8109YF7oiNE23ihcx+r9bYZt/yRF221PJauo
egesVT4vEzT3Cgbal9/REkGMfspXeGMMWAFpaiECoRv5y8MwJd1DXmCrF/mSBIyr860xr3c5jZ8N
yc6pkqlaB0X6aF/U+eGzie/Y74ZiF1u0Y9Z5IAiTDrMTIEBnuWPwFLMLDTnuRKGMZ2/EunSmN1/3
IGhnySqN6gyc9gwfLlj6pJd9vNdUBZSDbVLazaYZlGo1OjHC3ENihl564YM8vvs6/coCvYvMaUG3
qr4g/jBklZdPNSorQnwf684zh+ITMmrah1N/cUUnPcxRb0T7ON/li+I65L55I2a2VRSDsSXZEyCi
bQsj4ECeO7/WbaNDlcT492hPhlUqVXsw5roTAH3Jd8Mw+79YT35R68CfSM6h6pqQ6+dH/3m7lsfA
DJg9DBUB80j2SQ2ue+YtnLbVxwnnFxDwZ0kcRvvVoeQoJZaTLuHc2BOeAgPBz/L1xn60D9AH69Cv
gAX3TbY/IQRs1iZ7NN87SkVngdK6VLHAPdP3Hq0mGOwphnDtPean06T9is/oyfa66H4pc6eWuz4b
AFX5G6K4rU5dAc++8aH6z/y+sixr1htRghmULRV4mAhAEJfmZ6mncdEmd3YCtTPAfDrvZSBIJmU0
uPjo/PRYuRMIajz3MUfcxGqDgq1iDcCcC4p6vMOCw0/ArQtKPe63Givd6insB9rnZPRnuwY2s61X
nnOyCalxZKoKEX0V0igOwJiAjPDbjIPi9bBXte0EQrFfjYqyCdwB/JpzuFLoUbbTrWQWT8G1UkQB
SC/wiaM8V/CTo9Zh0lMf6HFocEllExnySRlNYhGUAO5ZiX7BGJhKZDYVYUkNWlk8grzsva0d3VLj
kiWxog2afQiq5eHBRACOJYRdIHO9moxznNWdwgW2hZu2NUUhqLyKIvWKOu2Iwee7ytLxZkgf8p+P
7v/G7bfUtEzGVbDgpHKf7ao/TsKbAhkl1xEGSqZKRTs2yK9eHHDUiUUumlZh8fYPKeqE7PRduWCG
0HMPeId1AxESwXcjRTOrls/kWAiv4Q6NSjJx2fOztiI85TG4lUDhPG0kEY0BSMkaqS10FO4fdNyX
NxHKRFj0UVOgRpj+xohiC94OIAoYTfA6opKBBowdFT/sFl0bP4P1U8Z1YbOIK/ZEbcwffB48uBdT
BI5pu6d8d/UDUY8iHqaQ3f0X5nuvC3glh4jku7KqRWL3OYknL5yZ4JGorAK+SOzi+R3CDr79DsXR
viSZperEJvWzQGujV26fmzjsKEdolI6hr0cyw3bzl1BYfYJJcthdpXi8icKEnHZ7VC8fcv3s/NhE
9A+CHfQ5dQs2qVbwW8E8VG9jvtWoJu/G1q/AELYIHff2+b55OdsPlR7NK3r/FML7o0kQ8icqdTcx
j4Y/XEdNyQM223L2/GZl6VOTfzpbORth9ebfy/j4MXYHTai7fuleOW8DTwOEhvhpzc9ozsn8Pv3g
BuN5ao7foZH0jJyyiqX7BqGfKd+i8UWF24yI7OVu3mN+fohHOYaZrjTXheSp8zJyVPlcwciE2mJ9
eotIMZcVGxlZ04lU1isllptlVLWGq8Pk88sNo+qKUgV9FTObZBu3VZhsI1s3hFcrHfrj6G5V2/3R
eaxmSwSOmSilIPnSfZ9FibhruFed13EyS5quZD8Y7gvdWGH62FOrNc1xT1hOTg1a3LYp3YMTyDsA
KnZ5yZVSH5H5Sgn6mgEaKK9fLLJVPPobHc/puhyR6+xGHAp3kLxo6I66ewB42mnuBeOsMIQct+ju
8RRi1CJP34kSlsVU/IgV2k/BwJnk5WwroVTM/d0WXQTgYkOqagk5HbRevThKVIb4B2iHjxDWh814
d0bhA5tV5NNg9hpiBQaXyIIO/BW14Jy+NcMjRBZ/mhqt/WhEKuex/E/HldaFHrnCDn11VWO5zc+l
d+jFKhXQ+1upLDd6Uhyb+kTJEnpMMtGsy644cY8qI2n94Vdb1BynNrMn9wxQa16uGeHsuBthwv6R
nA9mARv00136G+zjm4hKYtDLlNX7zi7CqP/oDjdpCRWztnuEP7cfnZFiRXbg9DHKPJJnQaol00V5
83QaLevlVAgLSEWKyqPe6baqfnvdczxJkvdgO9AO14wH85xXSJiM8GGdnaAeHdAbcHO09OWLBNmj
5WaRJ2RcnqlwK71kdlfuY7dVJmkMAwG4pbl57l86vhZSJCH1Shj43BG4ixG4TB4dC7hdmMR1Yarj
rXu+G5sZuN8XdmySKm01m8+b68U2WxGTsnYxl5bWqebPc/dO22VIv81k2taLQW2W+k2MdVWb1FaM
TIAIGlB7V9CGVl4FZ+I+tS1vDVySZZsyOlSKgAlljGHozJ8t/B8Ymg6hpUC+EKZnGZBOo8iK5eeB
aS8hIk/oqoCgKQdFA2Kndzw/l5m+S2pmvw4sjdQ3K7OjDx/R7k1ZS7m1rkrFb0sWi5R1ED54Mz0Y
Q9w9JZlCMbOk66oQXlcauposhUqfuT+TdTMXGrP5wRQOnIS8HsuSb2/d7eWtkA1m/p82sOxIZZjm
0aSzVGRA6BnMYYJfCSpq30Pc/q6eh0CERXDJ6cGJ7M1uMm9/u1DlqsbLO9eFlaAoORT2l0wbufDF
x3pSEb7C/DqcimcXe1KGf3j/PThScSWidDZiLSzAn0UPYsSu9Ny8WZZUQ0jnoHQsHsWKWbZc7Q2P
ShdtZtPZTEqsmj8qC9AWtgeVsGrRiAX9sHqZDpK/PCnnKbBABpv3ndTzSV4EtkzS/QSHDZleLVBX
6LsyfSsYvXNr7G693Ee4ZjrbxY1LBbsGeVihPNkyqzekgCtTvKCZeMEmndoCUZXSOeiLovIrxGm9
IstdjGzE9C7PqRu88FxEmLlWKr3Gi0zH5acyGy7zEgiC/B/ofM6LNtuDvVHE1SWTdOqBk6FtnscW
jFXj1gXT5puMrbV1nwIEwh36TGEBTXkv9meaB7PUo9b/94w2zlwo7XESaL6LDmsp8PKWiXrkdaRZ
+iXVOoOi0PhaeqnU7bcbR2CodcCvcT/1ztTR0juEAZQ6fSaCoF1QtzFBj5wiqYhbxige9ROm9sST
96uG0cWKYN4y+BK4fyzfhq6xFtzmRJqBW2C+R/8mzoaPCa+h/e0EASLdNM4fiZMVgCJxDNWN5tG3
wZf+NEnU4NO1prnTVQQItD+nePAmM0kmXDHenGA5indp82DYpbFU4WyqvdcwlH2X29HOdrmdhqlH
0fwTAJ3HCN4sOMi1RzttSKYjyK9+54jUSn7k1QcQ4Uo49N4onHoKGVLn4GdLHNvvfpwmtoFNgS4M
51shRfmoRO7DcKBKyThjkKX6EcslBzfspGqNmA5I8uzeN+aSZhsUHsGk09iPw0snoI6XxrKAigcB
5/SRA5ZG0CgqavtzCKUb7NnlwXrMoVVN7AQhO6kERg36KP12BLA2X0ayaTDmtyxLZHIR2E/DFn1f
VqHjE+zIdLvY2B6pJQKi8X1nmSFxIRY+wM6CYElerT/js++clqvzCuZXk8pMavSKmaiKjxCGdCVc
iUbwoESMbRlyg6yLcB80V50brjIrvs/lf3u0Ib73178aDxwXlrbxfSSr/y955D5eadMpRiE20rTw
QXdVhQhGdnNuHk2S7jO3vNpcmQM6UrPTIP94yB8wYGUKAOL9xvx1BLVDq/nzi6vpv5y7gTpyPviD
uF7CBMZw6PuFzP9AEF932Z0ivelmEGRB3N5r0l+CpyT2tjeVtXeuTumCf0Rfgv+YUZlZKJT/0KQZ
xIh1gYDDLFE3hbEdbok5rd3wXkb6BPh60fiOQc4AuG6+sYxe/O76bI2g1fN2Ahbggsp8n6n5OSnh
ZQcgLBtMaAuNh2v3EQcXHLNsamSnoQ4alCJJBq1PLg2wp92H6xr6Z8BSuUzk5ev+NU6BkFlvP7Ju
6biQlMxZEvHOqZDKbI029/NAYLFq8TA0IBILXpQUVKS9XV0WPTwqlTpFqGlykoXrKSuuS4IU8ykn
Bf7CyOHB5f3HhRB1AH8kBI3tElS2gs6uTU97pFNq1/AnAi+a8V2ETG7bOVmAtEVc548cYMmwyJ49
y6Y0WIDh68APzs9a3tJyynWY6jG36H2STkA94ftk3SzrIfBY1wsL9oVs1VKClZiLXZqP6AzUmzjk
xoUKt87+98QK2b/fcQVJU5mzdl/iBcHVeP9hadsQqIBeQCJwRCfEB1jSBpuKMcypYf7kV4bERmKu
NRlmE3bmKk20tsr+e0sBd/IhMK7c4OD6wNLJvpQqmKiXPfXnUA0efOf5Ue08LXA5s8/Vhh2oCUAd
wlhB1TzLkH8QnaHDmRXFwJOF/h+Sb6HShB2k3cVhNmNIFsN+/Hy6l1yvWJecIJF9T5/y4MRdiYtK
UcRlS87Sdtcvm2feKQSFZUl0evUUPeI0Tjkv4chwedVZFFVzqTYgbfKHbNUCDKKO7amalyFSL6ka
hyxISkVp45tXxZ1Yp3xW3ASs3Ru0hZO0z3Gq5W2OHxvx9J07/x6Ts1BHBtrVJEY/kjqZNwDMlQLR
ksJNxSm/gvHCaQylsJEad469EcPrTCWxljcpsJuoSJ+ygawP81OroITs7h07vcjEy8acSfdEyAMC
Uhhd8PYJfBOIOMj42jl2uVJW7/JCm9WvC1WG7ZaGh4OEst6+d+bGO7gGsHFIUTOd91U1FEod82i4
F+nCnIoKphgWwE/yZ1Rdjcqld0rbdrFemzTYnAvJsefrTYNhLXdJWfJbq9cIW4dtEv8MkC85EHhb
0rrG8o9lWEowD3ElG0iZlx3+7YDGSsjGgikD8O7lwjoOlgZfxVxnPVFNIoxeQOwAOuhIJZYgQA6e
Cx4gDvFYAxcqXeoHJVSu8OrU780Kr5NfYiF2edq4zd70QMBhCE19BV2pY7Z5aTuu4HzQDxsrQpa2
ARzK6NJ7Kh2YMyJ72dRP7iXZsouQTkM1j3A/Oah+FnLvtmFWMVUfWC7M0Ql/7oikuX9inYFacuB4
KmRgknDvMgIr2AYYLVaD5A1Q34k99yWYW1QFJKHuoULRImHwt1u+Tf+OPYyCuMxHZz/W6VkHRP9z
wNiEE9adgM1EJuz+VPCszLJtbvguTwTFyAYC2um2YSmLx6OnUUMBSEV5utThEgBTlQVGxaJheJdD
joaqVSNLoeV5+uY3gHe8ikxcKXeVKQibz58Wc6MTJoxlNxR4oQHXjR5ANbp2NYaONaijOhHfqr/V
vwh2bcS/Y9hydQImOtEPDqmw7vRruQterkIQ3k3ipz+RT/ZVkwbqeJ8iLJPVl1f8SQlMXUSqt9Y5
9RDGt5gd5ZmU8dpzT0ek6wg3luQm05nEgTAh7Lo4FKImcNs4YYefwr5rkT1A22D5e8NFYFiwhyvW
ztyRmnGYoVEZG+pMFd0WPkQRlG82SuKmspSdwd6Q4Wictb9aaZTcy4/LZ+7kSG31qnwleeyj+cXi
W5nkRXtRzoNFsS4vUPNyjK9VJ8yuTBv1Ctd6zVJg3X77+Gt1AWB550p33mJmdTBpXOftPp6fL2W7
KIRVO/Ws5B71R7tyR3wqrx+C0ndCvOMwmxE3XQLd9P3QUq1cNRMfWMbqm9aKwIIDtRnNsfyqeQqB
ZmMKkadLH7fkKgHnBagJkPycy2ySpzH0zlPRCScY1LHtQJlYxTQ6OIx15WS+C9nRtnvsj98/RtTj
ERGRcMjEk9xbbLezuRwzj1ABG5UeVmlaiSSUcifXf69nCLKkceN2Uv/gB5723lVjnvpUkQj35bIb
t0rHg/CxV29h/9AxShKWD3ZhDolvLq96NlCsyUWbKV1HOyCu5iqI4HE7mcqwXMRxW0ys/IEIapJS
duk1wnHbE/LOY2foK7icM/sBI7KtmFx4aexITgzvPviGPOdVYPE5kEzuVhNznInJ2qjeypD1E8o2
GMpY3zS+6nC/pOqekjVIgu9Kx3L0B9Xzo9RakmHvA32C3GZBz8KywM4+x1RX9uj1E5EZsJlTPqzT
AOf56HSvlmffbhj5PZbB9IMXKjhl7T8udidlTcgtg8XYvStH/o3nDze103/G599mmU4hwKYkDjXx
3wu0MseuXTYWr7RqNgUdRUbSO8qsnxWmGehqb9Vf6W0sYECJBgcQ6a32rCNUGq2OPt1YogKbdqBO
dfCnOx0UuVtqt+rxhzUg8gx1gTXGokKKH68IA0D7kMlCcBJXEnz6qTMFwm0b53Q+sYnUU8miIQBu
9yoOLSu5Ah1IeLUGqCSQFPF2ORek4zJJOYVAIehs4jNE8WNsD0HuOCtg8fykv4GpvIYgmuXbrSIy
uPzm+4cIiNye13k+X/lz8qIQCFYl/GcaoDs0zNt+DTTDJ4sEeasaYrLfPv9svklOI3ZFwlzeszFt
FYLDEsH8550g1fgrJQsgCno1EmEf7bwcil4XFnxIZy4dLMlHvMm0TeuV8N950V0fVW+zrBKFuDA8
REpBK6KMqdF7otaP98YpCIhShzaU79kmZxIP/B7cEGHnBHIsCefXYjSp6Fpx6+pDeiTZJeAjjxaa
OHX6XPA99PbUhRkPoZLtmE3DpDx6qm2ghe9MeLNplgsrEkylZT1g53Q7Dc7EYybpBARsRDDi2W0D
SxjsqXDswVPGd1WP0Ew3JAxgT+DR2vmho39rjmcoLQLoyh8o2dugLpXCbCproNs/dAmBcMk1BCxg
PqazAKU1CCxr+x7FmLEhEWaI9/PlEt/zrQfkCJzsDG18xVtZI0Gk1PN0DSrQH86Pgq2oB60fFJIi
aP1Hj7P2NrTdc/fgsDztry7lId0dxUvqi81/tXsHmxJWNcPjX3azFxjdye55UF3CFwIZp2NZJbCL
tb/gc+xnUDOUUZomSjfAUsAjRHifh7lzfrQYPX+ZBkVMALIhpT/Mq8TVuyhtA347IJcf0yk/0zRq
/ECmdWFnP5nQykCansj1HdsfivEHVTM1D0dxNc4TzlBzFKwYOt50vQaA2Jqks2x5ludmZKyhMJq+
pWS9r+IfUWJHaQcGIiHUSDGOFiR1SwsG7Np55C9AvwMReDDAB418vd310dMqkIRP+QZuwsad+Fnj
ubW/00XwuaAEhJGZ+HLbbR/5R1TCqcxpjIJM+y9Qfv+ooloCksKMJ+x2dWriQAB3LCgYNSH9A23c
Bd67OZiq4zZMvkPJTv/k2KXq55vO/S92DtW5FP8ZKThuxr+1ohtdGibsITfJrvuxBjoNmkjVUxe+
X8dfMeCCl/8kkSZRQ2+8DiU1ZX/FW/Hy/yb3+NQDWddiNVpF25amiyhMizct80BMJS5RjocPxb1j
OSd/su/r1Tnzyw9ZsNcJu80kz/h/7ABvaqdEs02ozy+glQobYqrLImOufexOsV4YBVQRBBh/1IE6
dIZDpxLDJ8bkvZ6kSxY1OtXAOL+sK/pwXZDUGEwRWtHTt5d/KH8QxItQdYvtadMPSyNW1TBEy+1F
t8wjy+HFH+zcuHZfbgEWRY3DoS/1Z3LuMcUCTiHrwTSQdneR2DgvCUk+dwkQTiPk1hAYawF8DoBU
oODzk7yp30hr3M6QDoklr3R1wPpCCEpIusJPdyMrZDGrOC38kTuxFhmNyqd0jubadDTG1iSP63J2
S0nAApa7E5Jel3qwt1V6uc5E/jDK00oTK5+3wGKH9h5NHfGVIcZvSuOIqMg3MMmATcNXRb7Yweyj
dcI74Ev9d5Gr9pTqgL/IrnFOHfwxtVxXQz/KCkIFZWWkbj6Y8MNqFsjWfElb8l5F3gsERw2NEcFT
/YwxB7efniloSacBOKncjxbgfkr7723gGf2raJ4HAeHiJifJs4bRFF1qKbM2kh2hgPISvB5fK7cI
fkZ4pkLs+zacyB7yE8n8prYBSkjxzgcsvgCc1cVzTJ0+ezcHAJvS7jRWW5sPlcPAyO+zWOfSJhOe
1lVVk9OH1vvQnvg8nlVaQDSNUXRxU/kI1f6TdWJ0c0gMfP6DH3Lg9xZt6ylN2gF+cKVcP2jG3LIm
+eXVSBPcIwGKT1qN6AxhKfc3gjZoEVAyYI/4OCMuAsK/uzhZ650cfe0Lg/op8rdfh7f3P2cYcWkr
Z/LV7P2EnjTU7zM+Nj7XX2RghhlI2rMeZ7ZKDIqngjJTFdIiNQTVbxIEvFIyjy9RTqbzfCSw7YLh
1RWPC9ri9iBrmX61GpTiE00XZp4JEugINMamphqtXnF3zrGP/KAHHrgyVHgQ004miaT5LJ2wZrXV
7b94GvilsQKr7TYogLvC/ZoKqcDYFC9VtE1lxHHLCrTPwOThaMNEiDi/UW/36Ofp3G28OtOK5TLA
TlwphPZI3VzKVkEmkAT8bjxfgLOMrzH2QtQAEJEM77F7bfsxQR9v/oq1EDiWyIU1RDvBllTaR0U8
g8RFQpz3CyvoLigCAdjeKZ3Tz1Y0kbaSfFOtEZ4WoJQqFwBP1hcfMfOwHGTAKa5s3rAZ00AN5kqm
v3kXAMWwV/6Zlcv83ukyuhedkBG58S8acb/7M6h3ITtI9ftSMtXES1ufFMLgJt6DnvkH63K4oC01
GcZHbhnF1NH66/e2sqVp7Gt82YwfYLrfbYJhafVmEK054lsvSDZ/E8KO8/ZUyqIlb7BJYE3IuleD
VMekXVNlhFW7Tk4HrZvaqJv9K0aZk1Cibk6WmYG7aK9aEc/3QrmhZ9nn8FnXEK+Mq21eE21XjZIT
JkL6nDYbXZA5CxLTdRfsLhSDJKkHIlbsCs0VmTPaz0piafVm7bTevV6vY38kv82CvrGkaC4oMGcS
iRt+/TJqUhZk6H47N154k/XzbNon3BxlL2+3/5x/OMX3nVldb1PQw7Hq61zlaDKFX9GCihWFCnVs
DvNT6I2+RHTB8LMu+Gg0NYF/ejhiR0y18HNDk3PAKSTrfdf++nY4FheYQb+y53vCLWRpejAlsLCK
kNUs8Pj/HuTEUcMMCmzyBsHhtJsbwo4cdeNUaGKxVuxzBSD8YJe8fiRK94LDSHqqN057UXlqBU8T
sTkPHpQqtzWlz1+jmcnTPOQxFTB3NjvwDAH1cXZm54lb2tTiC0lgfJG7HVVp2/PXke0sOY9zdzPi
CAqCWXr5u37LM5HEOUWwDWFyx4EQJpMDS/qOFPosVBkeRDTp4TFdusq/B2A3cEG5mqlcZNX8KcLt
0tG706lBjqbxeKgbZPAIk6CY/al5QRZvzDGGbe6tyulu8tt+3W65Oi1JaJC2kGxJi/dvaugUANxv
gYIUSuqrwq4/LJWBpH/oTvlJN/k5jcK0ZbeykFtCJH54hjd6uzilBkmqjZhujLQkItEeKaVwy+nf
EZP0CJ2uDEda7guc7wDwLBEynQ3sVfY1sAfp4T4/USHHYIWpxj0gC7KfJdT2+048YxnwP/mushIw
l9VpsRT9+KX2ZJmSC/zjNWF8NdEh5xMemBWZrIV7yDP3paCPBFCmEfkThY8r/Xj4Y/lFBnXQ5CFO
MRXis0iribbFI6HyaorlC5dlMvNc1jrHEj7afEx96VL80i78pNUJtISGzLiDjjknw4cvFiwO3IaO
q31Qtw+g6rMKtKi/ZUCREsP7y+i5ZsHBk02Dff0uxa2Vk8hrfXYBfi+RJdllxyK8TwF5yDNJvrDv
vU4QQRjxB57G2WelPoitLR9UDAX8Fs5kHLLnc63ebrBT6nxDqg77/P59B78vpI0sQuFiLwdJ+Bc6
VB5olG+VCxP1xBwX6lyCk+PpJnV2Kg5y7naZ0wZshP39BndDtkf4Oc1bLYo/5SF8gWYWuN38Rgy0
XFvnX6GwXk4kW7GjV2TUTKqPU5qawtVkTMXrMzm5Kjj7TJhjB4ViiOp0jGLMWRrAb23vSc1uP3mw
sREFheGiE0zDQONC/3kuN/pVjC3RExoa891jNMtxHuMEpc/XBePaJJzR5rtQawRv7xKk1YweVf0Z
5+y4Zw3IvBu/ZEngHs/HGsGx95v4rax+eTElhrz45sk+cBu6MOk+uqTgOfZyhiCD80ytys9xwrWq
NgydFS/Ozk08LOnFEtSLNgXO7JNt+UiAMkzZZSCL1V8YSUZzvaWOUXs3px8VWVhVuMXzm+GdBUEL
J28Dfff/MiqX5W7TRVqFeyFLnrGoarexuCfG/Wys+1Z0gKqfW/daYqm25LsnaRjXsQ9vTVHauTw7
4SoL9AP4qLUZiFCur1H8b1cGL97gbk+8tgIxLSH3ANT9g/2wngKVRWzU4XFHF5nJe5zN8v8yf0cG
LB0p2hGWpCrSIrg1mrrzUmBL6Qfix0rCvKZDSMOZoD/rswSL3NaW75MUF2Bwpnb4STAnPmMMXqKH
YaSmpSdOKw+ebDrbJPnfzQ0g891jwfHUjKp6/D3XLNAOfNUlKDPcBsCnC2joF6nbcKZtt9zKLq1U
Kh+E7G4UMKjbQsA8dwUtsu2pZ3Hei1m3L1qDnniYuVnfKQNp8n4L8Si0KA6EgH99KccJq29HLNbQ
GN2Z4/U4/T8XnNLWCJbLRI55D2Lvd5YsAiiynrPXBUtSLPKFu/a9yrFcTsOnFWlFxvsOtgDEqe58
lZIwvrOJBtNip4rq6kY3CMUo7+mYRaD4SV2RL56obLpvxJUve2Izi2tCtnhWRZxVg0Qb4EHI96z3
GMID3ipJsmOO/s315Dx63ZJxqmdJpL3Tgfi3/UirQT/QyG6PodsQeQGS8SHHvUyWaD6tp6ynysZO
zFFwpeSDk1jav6NYLoAUYy8Fu19dVQHPoqMhstm2L8e62Ul8CQ41hXclT4Nei5usD33d9iAxQo8s
DI4NKl7DLEcUV1oTr1ER3ZI50V+RQdVumikFTW0AliaZyD/C/NEt3GArBiy5Pg6PNWch/ex8Cna9
Ob0bWV9QF+D8o/FbC6t83R9HeT6ZKUsJPlE9eqMsjEqDorgSsWGq+X11RSerYIhm+gzaETTP2XA6
ZDJ77dBHqcRu4QjZy40lWOAd7Z5A/3s89vkC/EnyGmXfYiir3xTb/gg/Yy4O8qxe8VyRbg+l1Bg5
xLd7t5FaHIwJBhrHBvdulB3nLnORFAAYXRNxuIL9SDs8eNE/F1AED3/dtZFkjDZdpRigrGvCKEAN
U91XjTwvHkU1yarG+xTzUudheCwpVu+vTLxV1y2BTAmnF24mk6vWk+OrxhvmTvdBLOtB64sb/B8m
vlTQPTskALsAn0r69QeVxpvaHx7cgtFsHJ87TVdDm3QRyYYuT575aaU8KcUI9LfddewICzvoeDY6
9OX+FS+gfAyfp03SsWFpny7VPxlxEBUzsItaYzk0CalbwouTREG1NaWhAJ59XJCIgWuAckHxScHC
li0e/aS/uSkQeJQ6w9vKLIiu+treUNpoj4iUjnjls04mhYhZohEDMeZtygXnfD1WLXgEnk9K0N9a
VZbDTuXRRjpQI8mtzkOEP15GPquuZ44UUqFD3ln6eUEGeaCSJkWX5vGLCGmrPNcPecWQ2UlZcjYK
CeoWeOsVK1WE7QwrDdX+jGMTOwHBESHqzbrwq7FAHMS9j3DBN7oVkjBgoyJy+Zs9JK/jbiTeS2gk
2O2So6aictyu+TC4MTgufHRfaiM3/frmoEGJ0XRWbVu14hs1fDd4ccH0xgzeaPdCFrFiV82OE9oN
Cn+QJy9+YKotCEVbEToCxSQSZm7AVrepNtv23zQ1wj+cJqEKx/nYZS0UnCTs2Bk6v8OfFk4tecKv
VPciehGXfzx6Opc+sfV5lZ9TYfADvxwaCpSxRtNicLWHI3w/8ZZwsnvG1sVEpcQp+OSZAjVt3Sw+
kFePc7ayvxEun+COtS2J9WbEEHdldIuWrBfaswsdikRoSOyVcBE/aZxPbL578569vJj4VIe8I4nt
/UmASNLbLFkaDJw9vNhAjPsuShbuRqE3Mcfa9UHQ/6TJwFhKqHStdHN9e8MP20r9sev3NB7dUhs8
5Xq5DSe/p/Ne6esi4unuL3r9Hh4fTa2XbzeIQlB/0TzwQNcwF64c9yiLIovO3rfwaGxIwZ13d2RV
Zegmiy0JgQojTLsVieOV896OyJFLjsGkhIj73DM8uox4DUcSEY0EUKP8VymXusstTZJPcAsiU4bM
X7eaGo0LFwljrICIMPhSj+1UVYjpe+PTG+Wtf/WFNt0yLCyrAXCTglbYuyjbErA2ut5sKbBi4wul
PwPyGeg+XgGCQiQB+R14gXlIngyRzueCGRldD06jyQZppOYOdkwkXPFyanrlhbe3pzrh1Lt0EJQJ
B8Y0B45CNOnfTxZKAM2yCGrh4zoE5iY3thtv7zMXxQLL+oNChocuDUERs5hBeqAYq4ZiSoLy4JtN
1a95Fp8KN8yKiUvcoCVS9U2w58IYEc5YJt4kNPd5iw0GJNWwtzu9Nlg16O4bByWnGvtt6pcYWknQ
EoraKlcxXg0yPE6FjIuMsd6logwoThJ0SMAYtfxrKVbwMumuLzKCFY7HbsWkizrCtTc5xHJXkeUH
AHABLbvQQaXOHRtKRHX75RIirk4te49Yycm+9UPKqYN72HpMYvLD2zPgrf1Zh+JG/e56fTF5vcP1
QU+hN27usWB//KV4uhMQIQk1I7GWRLBT0bMl3PQXZU8iNeDSSF9+LYC0sO+i7DaDxRBYtLd2AeHR
8HdG9Qevo9kzM+Kt3NenYg2ffcWlD0iKC/D4hDWOTiRGHcsxOVtgbKDDBOf7iXWisWDRTvgEcILS
qG8RxXZKjLhtfMuzxAlt+U+9GogR6TinIq0y9AbB6CMqu6R8iwsElxxPk/WycYhFZ+9vnagQAqHJ
yB1gbqTGa/IGNG1AiBd9kpqDbx6O+YDtvsmG4VpeJRD5ShRnkTcA9iocYTF0WxF5nbtoYQcNlOp2
aOdITCXcDC8P/Hcrm+VeCq3aocMaWa7Wv8v5yjtmIipQov8Rw974VNXV/fUqk/GNP2gV9g8H7fwg
iDPXx7lvt/wJvDbAQ5P6TPmJoiVK4oAAauL23BRu3ELTrpvkRxZr58oOPOJkceuo++vwCSGnh/Vi
YvK6w8Y4AMVvj7Q1IoA579l1b5rfeRftbM7C6HvxvCA8dJLJX75qS/cqRlNvS+VUdCncyelglVF7
31vxu+HNAhCUy55z0KEjJci9VolQ0KSqq//ZytBdxykLMbcMMullycxFK/0VSU2VhTgqN471YwVv
Nrk6D/YQpGP4JjnEjhBqkg3LVyxvIPeb3mdw+b/AHzLeyY7H9zAE27ltJwsDxdtgwE3LFnWO50eV
0UB/CTB4DXySslNjITW27nV4hvyAz0Qa1Rf4EyeNXnoH1I8x4IZvoElgKt942r7JsGuPPrdqqxAZ
bolk+zrcT1iaLs+KXGRG4KmQI5AC8wvjm1g0zismdfSfCXYloS0/lt3oQDAr33ya2RqN8k6IT/Zz
KVVcKwFgP+8cmU9yq8kdN8CtdCtrdFgIuyQBSOjxaqHQedSRLFTNlwFnEqwBsFI1RphvnehKIwIM
ZzxVh4g7aehcGBvDA0C+6d19xDhdrsahBDnCUvDGqrGVgACaoR0jjk3vX+khUexV8yKakkY9ozx/
gYDlJB2QeJ6jKG94+HPDheTMqohemh0Qi2muR3YzUnRf74B8Fm4kMrm6aOHU32f0rW1U/nUCcHWi
4S+XeYv442jbegvykIm+bXfq1ksP3QeOxsBkKqgFSxPNNYihb1g1kUMwtjGGKcv9kIjQmKv2UeUR
Uw98JfKimLlczF0IFuUYyb6XRPl+VCaVFrii2Knmm65jNEqd2rJszfU9jrWeXQ7zBzopDFenpgYi
iphOOdDPlET+uV4OeVoBhjwkQQIlPq+PVKkT4JEuKu/bTZKJqVLx7nNCViDCRIBz1yZZyHkqGE86
kZeKlgVytzSWmzA0FgqeYkSi/WLkXg7QknDoHbh/9Hutkm7s8hNjhSxuSGqlQYH5TsbbZDGC7mxT
7Pu7SZjON5BNUOn2G2mEcbTK/xNhO8wU3NV3iyW4q1E4Y+csqDq3zFJd55pYKmxb9GVjtqbeUiv+
hDEIluXb7mVHtSwooksvzv5lw2yVUs3iRjVTYDukAMF18FFAbR5J5/j3gNFlhRRn23zJ2ZXnQht+
w7p5F5cIAUBmDj135WXg/IiLGNKmdcpm7y3HJfrolWHIFuXP5OM6W2F477+CoZ9zV1/NbSZmvcWO
JoDIeuLoXpWL75JFrzwg/VfNeB9q4j0WRswdfAF7VYSpLPYmKSAj9o1C+rzWhrR1125YpvBl1TLU
Hemq9BOpFhHHgzCz0OkesAiQ51iFqPSMlkialNKPyGM/VprqfJe3KeBtyBBotEuQAkPkhOKXL6zq
chEWazV2cB85NjjfYNv9hNrRrYUh3N1k5xt0dvHquTn3a00xp94UM7VEvEh3fnDXBB9znD/+qztS
YcQSp2ojMrmKZoJEUZIFrOXY1QsEkxHoKmNYUkWvjnjzvkdL6NjMFlY5putw5Dh20r4R7ZVPNBeR
2uAJV93r9ql0tOJS5/qYLI+YAbqG/TeNcKKEQATZ+bubkccEPam/2EyT0u0LrUDjLfcJrVQ/HtrU
KKwOA+9XXTaKEEcmLNrRD+ML2PFkwVbFQSzjlLFdsNGcGt1hiqzu/kn+gkZ6OCCB3s12YAb+u6cQ
6yu67caITYwf1yiBjxseKDRhYEtQ9gS2M2if4hxs7/jgNqs+GqkS7dnROyYYlNdLBZUaPvUEYuyt
ziTUJMMl1LqFsKNXDdGLAMIr7+EYWmWwqrhvtI9eTkL3H6BHM3n98u9MpOaQAuNqiPTw6saWj7QU
MOiYTazrY37lcEQehOWZW1/FR/JV6jGOaC2X2p5MPPMbuuI4nwbhGMZ/KFtKuXaV2JtMu40cO9B1
5ISo9lNBHOv+pue4oLTM4PpdGR8Nd4vPvrK84mXCZBkWKPA36KK20TWl+PS2rXsHkmqsivQcYxNW
DfAdABGrpPZKUQrdsaSA3ywlX9nPF8IhUqrZlb9zHZAqFB2Cw6NihbhxA1DIrKFfB1wtiE1h6+sN
Z5dZb7ALI3UJPU8RvTSdwKbar8UUbrUG690UOn+O52F4w0oMvNUzbTiKXbxEONOZpA2sCLBV+ko3
c9oe6EX429ZZZXHIE7ez7BSgqGosInDa1sa6Z/C15HdcrMiPd/gsut8l2a1D7D1PkoZgerxa/NyZ
D0OZ6bqAO5fJFFWWCVZY9kGA7VJ4K/GuS9XLYIIndN1SgDyNW1KGNXiIdNNic/nHjOsl10Ef8K2a
3MN9SLUfido/XAAYkkUpTuBCRhK5b7telJ5hOpEac3bq6DK1hKQG2jPm90HEqnooQ/kvnH2PExqk
B41B7ZBcnxX1+3eDGWuAiQYdrUnK6egIK5Lk8H1MIg589O6Nl5wTmUDE7SEjhgoxnGuvg9k9xqFX
3p+AC+FXowue6D19hESpa9ZBvbXgNi616y/o1vSfD008j+c/r472RPattapvRFKnTcGypLfptXCA
dd1XsRkLU8fOjQ/Ub0rk6EHVQ6uvZABlpl+Rt0U/TreNY2Y45IAGod+PhwiU/LnykCU/K9z31c1A
OCdkHbyC3UvEbXT23/oR3z71dY2xTiixrjThshQrI6cxhlW+e45Q6PvvVLt7VrpERyIo2tYbCx1K
DjNRjzvsCsb3UyotoABAXPWe5aQYyOBEHKZYp4zR1KlqXb84a8Twe2DGG6rSalaQzBJOu+KnOr1w
GdRdlwPk27isIFI/VzLzkAjYTmaF6xwFAmO2HBbfKDMtq81IlQ3HCzeR96y8IMm85exCmMMkxngH
26EBywxJNJRB4U/IObkAdpx7OM1mqvifMyT5KEA8IiM/26mtBDSOXQWPRRISca1HK6XErSqzV/Zg
QQRYVidA8k5RLMI7cE7CcVHoM0lnicycxmxi6+Va/SluwXbEBZOns3mVtd+38HwHfAMu/HYyjYzc
NTjVre4SnIWxZlnps255WJKQP/sXv1u6JzoS/XQfTQNRlmjuncLRyiDWmT6fNUldVNbJTjl28VnG
grjC7IaZz+ktwKjevMls0GclJRZ06MfYz4ToxOep1c2vgkWy1D//AndF8g2ZjLb5+EQ5gYqf/2Da
rFgUT1+XN3iySf9C/uxW+YBt21EtjZjb6gX6IKa1pkk8h3HEJjL/7xmgT6ZDOQhbBQDRe4UBkorT
l3d3tItTAOIivBnOFwCLK3DKZCOX5nxOs9Tr8IysYAjkxz5C46uBt2t1HfjdFybtg+VqzR8KMnxR
5g5CIliPUaO7FFaAn9PidwJfjgq1/84FA+4J7SQN10pSCzrKs18p/PytSaEHo/qBGijJKLbnvm3F
0jWJD0Zuvb3ogeJhSRSsocZvo3mOiwAoV1siUhjE3ptdHE02dCmWfG5DwoEG4XWVHjMxfGJme6Y9
+ZupyNBBHWvfMtnQKHjZfDOW7Nt9RZfHoqd5bRU2fq563TmtiNw6/MosGK9pkvxu83CgPOo5KJMD
8VhqW5VZJAucBFjhn+NQ9NP5AxiuUkQYfn677oNRNhfAzuE9fZPLtnBh4aQmE8wYQq4k6hY/yIAx
IsKhQiU2ShZexvOqphxqQehpR2FlRtK2JkX5Od6TQdTb6YQh8rrKHGEil6IG3/c8NXsVrGjdRe7V
5+S1CU1vfXadI2ofap0ePLgUwyGtGiEHNLdCdzhFOpXUZE1uG2QT63eFbJuT59PM8g6qi9h7vRNg
0vIQ3Z82izs0LLzQcnVcEogwjd5Jwe4PN/tt45yKP/NomN7tboj5hwydfpqIurupRXnbq2/VtJx2
EIT2NWoK87RD2a77GNfteOmOWQi5hY+VQp5TU3+SDHdkOSZr96esji1oaREkl6uCe30RGwnjSG7e
HI7iUNz3Jg95HEBe3yj0O5YpZIPWQe16T7rR1/O/qQrM1dqvcgTVotsUPJqNrRGeiY2pUt6/gIED
lhbWIBhj7DuuGPZk1STvFGkRLLxyq/gk+MmS/h34ocjWHnD8+xBQqNZfC0zNB09D3UygcAoaSHjx
lGxht9kECYst/0mvQ6e8y2FSpjDxzlyHEel+N0QOMa1bWLFKVKkxX6+WQlgIRTMWGc/HydW+fOuK
y+czxfejLDN0GgAIM0z85ogj3EyWi72slmLoaiFT5MhzDYd+207JTXl9oIjswhc9Z5y5rxbWLnCq
IIwOYjfN6yPfVitAOLFu6kMUWQnAIk+UcEZBrE4fpESNAiPubKlE8bnOkiVFNK6xq6zTF3Ybfjvr
p8EYy08cB6QAYQ2xzbybAhAEnI+DRlNX3dhLrSnpA7SLDDiMCSiDZ00GzTpUBcq9smvZcTKnuae9
uSe6VwP+B0546EnemjidH/JRDWgHNmUO4Zr0TIBtu37PIR0iYTOcqQVXqMwtFUuKhD5XU8UUvpFw
+MkrW1YMZWzTZxzN0qygzKk0+HR7csyU6Nw1OLpWcC8sikw6zg88caOvmuEMH37xUb2Xiy20/NTO
rImyk85iC7Td51dO2cNVU/pg35c2AWJTzrAunw3CfWAFaVmBb34uduywYiNRJsfnEbDlr3CLgv7b
sie6xb6o+edAklOhjrV0OtanUQ4eYxcHkPAFx8SDqPr5MTAawMt/tajIio/KPFA/pDP1ny7GYrn+
8vwjZWynigcCvn0cabk0SvNfXKoqsXX+skZ6/cb/yIjAtv+u+m8ICO8PKQL/bpELx7dTo5WLRUmB
Cb5yIPEGqSsTqTuDOdkZ6qHTOlmoVhpO5zRUn38+N1GhFUjEOSFqu4hajeYDHg9blLsnOZO6l07g
gikV9uWItJUzvBTYOSzRML9odiZbw0Lwhu9a/bgUyDmWQwgSZyK/ywEq90GHzOjb6pZDofWVL15d
VNeTTyKk1P+PwmL0ZHvshk/ZEO1OvXq5KveMozOJtjwLZhzvV1/0GPuAuII/+GQrzUpQj0FsAHLx
VdUJFj9Q1lInwgtj55s5/lmV/2iS/KHxcK2peyJniOsPhqeyUpwQa83+sUefEiNT2MGOSSyGGwHT
c6qEh0g3RQkFHM2vHEhq7xWxUMpXMELqNjuNAh44CO3LPVgxPXtHCpPKxIcktO5IcZB5K5IQ0KBE
mntgb3L+wowXKoTFmmhGVhqoc3zCOM1HpkEbgUVgFIRZm092RPEM15STG8ADQSvxvnzwEEKVtfMN
e77WLScoO95dxDZ7XL7oHL0dgeY46h669W5NE9lyXKieBviVTa+06M8qcauRvwwzPuYnbf4W+GS3
ahUFP+4p99yysu7VGqZ7TmBjOljnBj0+wYqPdTGQqu19XqtkEraZTfCk4ridRMWjKCGT26xAhqrl
QMZFW4v18yqX3RXkKeh5/yUedxnK2/Q6DXiEpZIKMQlIfQf7NfwcPQfY7NGGE+jnM3qsvDHrZbWn
k38+6Gl4wb8jptYSCBWFwSgm1qCRZbK3Oxfo4xt1SEInhohn7IendQhIUEGIg5fCMrNgXdaWjEot
5aWFugyNv3DgWs1OqlEk8fEMxbW7ug2fDddq7cCDJgYh4z4VVw6D+FBjvK5Q5Z12fl3GmabHQm2P
zBPnnoDCXETCAVaYILYXxSLfJRnkG+64TJj8u/Ng+SSMuFiEteKEdpGNnPPLC27OTm0LvssBIUNQ
iyN18oscNHKzEV1dEers0eOE2zJFqz6LeG9u4H2swo/DMemeGtZRBnYwErNjAThSnd1nuK+xVWhH
H86DuVkLUPorHu5zpDW6Sx5Vqjq/je72ALMJmK3OPNVstiHpPaIikpetA1djbSDnM0UIJgI+m5Wo
zdq+fCoI/bEf4oAcWEtRES+4d1xbMuqgGxoWCWmqHwYP7dM+rwLZAfh1dUcU08X+o67uFxF9Ud3G
uTuWkVBzr+WGO6ohZAe5dFHuwqpgNf59u733BoKYUP1q8zew/0lI/O3lNALu8MfOfD1JnYag1SKV
p6XsivNXR/Tf9GMmqZF8ZWZBsTsElFlMA11XZxw0l6brwaJV+k1UT/6LqduBlJ5K58mpET9VSzoQ
WpSYrwrGnHacNL+EH/rvDmMp/EpbvGBZOF3LSPFwayKD/q3DtYYsecmG1pXJFUh5V3YPeqk3Cb0E
kRjoVAVLo/sbMNSHwCpwx4rrva4QNyMdih+rD25BywBTmizMk7guvGYppwMPTRZ8LBD3Tvie4DO8
qfOyY8MGJ5CPqmzSyIsJmdulAJcdiCBDmWwHxg628fd1glmbcA0kyX+ixL/zSZXB/9C6Sh8SM/se
L2lzdRhTjzYnaiG4FXKyK+R31UVvzQvqeXLSoLo4yYr5Wy2+o5g/tQ/tR+lGNCQ+IyXqc1ds8zGz
OnioO8/cSxPb9gqffaRCxlNYlkKp+HhVBnNmr5SYedwid92pLQZHiCWffo6yUf8XHtTglI7mTm0+
3XpNOLRGJZo9iXZc/Au/yy/Q45tV+Ww29MtHRNf6+JuD1lnTJ4+Dd9Xjq2SOYTI1xXZ2GY/821gf
Aie+gYXofG4IlXl8xlL9uVzzBP8PICmvLmFytsOsF5tQOLQZEgpgGYyIFRSVIOOHEd29HGYEDLrM
/7IrDnYMXyYVC/9QvEKUfil6qUJ0GzEyMdXsT5Y3J9npu7xggmSIOYhGOYS6h96qlEF+5pGWGokZ
j8ZVRsv7Q0ZhPZ0nD+gqSYbEipxnJTyvliUq5rSYDNXa60BX0jc8hM+uDsBec2gTb5PV3hYUCPWe
ax273Gh3WNkOMzdRar+Y2ZqfHdCtKHyCAA/bOApvCPe0zeiqNb2V11q2iTVANcgHYUD3g9kKBJyi
t6sWf+GW2cS9cDmJNCM9GdSrO7XfLAWRuyga+yIwPAR3lTXcQK3mASm+ldSKhz/2K3W1JUmqYWVl
2ewFVEYZdQ1IJos0gsUtEm5i35UVQ6bUTalpcjC/kXxArOTePZ2W0+rUIONzYmav780IsDFaiM6n
HzfJQjgA91alcMLGliWnvFcGZ+ew2QUihR5QN2MIHW/BvO/cPkzAFrcGMYQtHmH38DFLTPATe0we
V1kVwPYzq5nAwzZ0cj5X8GJtJWFu5qP+GpyQqICQw1W5K/1zFUCj1SIx4Za09VexFFJFRUmAmTj9
qgiCFnB5Pxg71ARseQqMFmjgsBlxi4YHtXu7+jb/NystzbgH6Eb1Bl2IHR6nBH7nmc1M7Oe/CDAk
ldWiYneEKrWAXHurKJOTvrpjO4w/5a9bLs42JqpSv9psU6kWg7cuJeBSMid9JsOeuwPUnCYqnhlK
T4X1Y7A3acPZqfxdRYaZPinHYJVFN+KWD3pEXpspXOCXFbmlVl+fV+5UWkEhizTQhBS/t5I4jroI
oyyYduFXmMrZ69NNz0XJyntr/80kZq6tScgV7gXx582HIoF5HJf2tyFKo6Q5EHE42+1fdvlWe0ju
FQuaIyyeewfY1ZHNxt2+xMkWfVhaDJo3XCfMTftdOh2K/U+Zlg7dwMvJPyIZSTwDQJZGgoB09Yvr
Wo8J0D5/sbd6RiJPNS7BjI8PmkvYcMo86Z8ToYf6jQfST081PrhTy63t4GMrPcSHgWOsvvlrNUzF
+QW53JkgH5Mhhv+d7AWTVn/MlyYSuxislpb3g4V5cACaOpE1hKArOmZS48xUUYU4VNXdlh++vTeH
RKMR8kpmm15AW9IME0OIEIKxhB+eJt43ym9btbg+14Q41DMHZuXZdzgW6kvgmadiErVtfZIrKlhc
jbu3MUGS/uK2dp6vq+ANvwABKWILCuvb/dP6/qjB59lbOafvj2UhOEFjPPOfwZupCmzqnbaFujUl
ya3whpQ+1q8gqfgIO9frHdyJpxVxz50WwwYbfhh2KBvtKl3jRAet+9iMz+2JKnTCIYpkThchMpys
KDLrBpCeTUJs7kBCCDTNOdtm45/0q5t12u4z81TqvbSYQbYVp5qVdhegrfbvfZoPsABUnMfLVTJ/
eXc8HXYf/euaFa5s9+0c4R5pRNEtdw/P9qbEeoKYAub011IIQuj9eTfcIN4GhDY8LBSkywMroMj5
JaIrX5mE5lFAtzfzBHd3/D+5UpKqAKbnSMXc0jjOinqv9ZW2N4xoH4YdPIjHK1bhm7zq5ERHx54e
Z3PEl100RVzkU0SlwSchtVr5bLf3cYtsOdXN0W9l+aRVnP2G7QQP+gzXQOKeTJ1ePZCaR7Q2Y4Hj
dUnqEJVGEeYQIwAt2f72q+xpOaZ8oM+3CTnqanq5Cwe2fqMIBUK8B/WUYLSAjOoT0106tYI29HHc
0kKjyis9wL/XwihulsZnBXF4AdhgOyq5PYoQBy2krrJPoJWxmp2PahhnQ4rBumn9f8l50gj0xkuJ
jzvKM4Glwhrjlh5D/WehwQAMPIAznGMG/iujPjNi11VzlFC/tz2UBzM6J4hwKKA9sRFV6IvhbIna
m52BplmUJMbin2WL0pOmuGHioYIgKvvv92unHSqKdxUOxICiv+by8+kphvrtAadp1zIfsX20U/Y+
fFHzL+JO5HsxzkXI0Hb7LSnRIzpqMcI0qaHoaV7JOgxHFhRa3KNVj2nRr+RA62aySONYmepCKssk
WJt8sMQdwWNDfk5HESZ4j+FRPO4epVofz7an1vOiQMivKyJfFBHO14ghEvdmZ46Aceo3Xoa7VYEK
uxtwxD2RRa2CJeYRg9g49leIrJP/opsaUYgF8p5FKVISXfDh8f+GsX7nB7vWY6xf3IgmJS3sVq1f
KBUBghVtB3GKZcYPf1UjnMfN28XbJ41rqB7jWjZKWbB/sbga5dlj3bdk/gDhWXgjBOCiPOctIwCq
l8QdGPUMBfCssI28Fg6V22mui0GMEuzRPxpdHM6XD5E5L2w0/iULlHVArr9ASmXfd5jDjTKnJ9PY
eU8y11BPoAY7G6jkqbQVKpS2t/dYMJe2Rj7TKzCf6WZlPBQy5urcmd6IAg4oJ8VTIi63homTghwf
FL+I0UR1lsGGA+u72QSM4MAScVY0tMP0fPC5PNHo1kWW5iEMQLbM2FoDRWVh2kq8qwBQcjmK9IyP
AfQOC3IZBXBJsJZrJFh41rEul4MqcaWL4GltJ/rB0t1bQDcdR4zeJnwQRs2yrYU3/CavnaFGqt8q
j3kH3uZ7veS8/GfPWgwHdksRNDup3tsjZ0HkT6f1BJjE32RBy+aGsYUFQPBAHX2qNvM2QR3+fQ3g
Fes3yZwPKjkmeqoHiJTHVxZbrKfoVb7o29ndZFd5QeMOaDCIn5RBZgv3XLOK4MAoO75TChIl35or
Xd+nY2uzmzrtA93BFSt248MzcpM9IbGskcsyP7+KUq47scuATT7m1WPjZOTg8cghXl2X9GQRoluA
0Tt0TR0de0QEcftSVX0Bd34ukJ+Ktn3wY0fIXbDa1iXj7ClZhjvrp7rQFzN0uL/Ys/Lr6HMPeofm
ze8lR1iwAPVs1xBSF0xRwcAxW8a8iJunInIXHz+8USsVugyWzKMsEvTdvrrPe+t9pRTcKTvUo3N6
9dhWYSKYfEd1Mil+/pNUNS3Z/V+PY36DREU7io6IZdnqQdAa/TZPG619R3c1bqKx4o0AgfM9OEgC
px4k1cURnHZo260a3TUEoNc+bZVNFJL8cmvuP8WpSf7umiVBaV2m6Bm9urB9y6PDYVZPiKRRixvC
vgFUCVXvJkW3q6U4kpZhtI64z7l0Ufpy1YzIV93cpZGIGjo/Arm3Wt1Ag77xRwpzRUArJR8XlIM4
inV5X9UMk/4k2F99q29eWLCED1vRYI0wFh4j5Nw2dqlTWBvZ+HY8na0u/p1coEPj4W6I97K+hNC4
/KQ66DFjiCB97UbrvMBDuYQA9BxVM5h9uKAAibepU3nVvNl/JOV3rG3lXEXkrh7+bsBvdmesLp7Y
AZjH8nq+29hul+kj5b6yzGoJG/Jo06yN8VLuq8P29LM2mO7snh9WRfk4DS8hlq8EbDpWnwjN2G2t
FR2qMduijGD2Fc2+cT+D2guv3hvKQLkyPKpczbVn2tpVchQ/Rg8+TEeQxcrGgLCkaWV5pouzJs37
30+hVjK4pYQOsbeKWUztzJ5ROMPjH8x9/xBye6NNP9tvOyRiaSjlyv0C4hj7E+nRmkNDfuSgJQTQ
B/er0wmAcmSnc3I418sZOfECoRMGH10/5o42J54cLJI73gtdZyqt6DN3GYUark0VRq6OidfMp6gc
ZaArrGpk6J4xSsg9JYhWRwmbubygM29PGSW2Qo3w0QHEXs0Xe7/FkE3hT8/XNWBtesdm4ESMLEMA
/m7eubQYFzLwSqYMYzuc0zTU3z0IOegpDeUsfVl6WkAU7sqZvJmPQMvWyG1nx/3k66tsJhHboqBV
vkyeGnr0Jyt3iJH9dNCukcCO+twscsD+0ohqwXC1yc85fCWqYKt2TAbFVQCa0McH4mhEmD0vHMvj
m3faU4Qyxm31aU3EcXuVSGCxe10Aj7hbRs/r06Yefifzbd6H8z2QFlzwK06t6rckXCtp2MC+lTnc
iYpozL9bALXJKfNfj3/XKP4qnx4woIsfAsn9MN/s0KB2HtOWXJDsTNzrVucy0kkX328cLFryPw9A
k9LEgTocVUoYNqAoPd7wt/3bshEq+1YdSd7PCFgZCGLlQ7v8xnzdVohZ1a0SWiGUfn3EZfuNVkH6
FKzyFKxv1EC6nXi2UpcMzRM9aVpBtFdbgl+xjEi0zjRew4uvgT0sqYSX1U06++v+rW6Sjmu8qRN+
199ALm4YA3u6529uYT6p+e34ZEG9ALvp9lI5IoAXd+5l6qUzLmRB04O984Nqy0gfaKW78SO8XikY
+w7HkE3DM//Bt/lUEWcYz4I/2f0LH8ZhUHsgEm7nBa9H7JU3Jw0nqxI1wC8GIEO3hdQmT0DlULGY
pwupyXXT65LcrtDQZ2QGZK5b7yG3AP85w7cI/EgJmHJWxgiMIKwv8C0E80AfHPj2DGPydsDhO0Vt
3JiZpHa9UYAub+sBYa3slZZr72Af/Y6ibOx5lLGRYg1yRqXfwx+7sbcXVp0j0uOqa3z/94Q2unfs
Fp6UMb2IBWqL59YT7ik9ty3QhxTICM2CEEB85Iwu4/t2RL9uipU+9UlTGCCG60RbWeV8/1bKht1Q
gVWSW31qweaaVnosuRuumGPfynrNAicHmeKJbq+Laa7X7A/rTbxzgk88wchxNL8LUZAEb15QvI09
vCknf72SxYntQOx4rjpixRrvl6Atp7anyjj38qElVl4ttjq6PuqkUC21ZAjxmBdx3oS/QG6zlOaW
s5SWTcuEDFKb3jBhMofZ2BE83pffLpLGd/kYsqC0O+MVcOhwr/b6FVgFObgnrd9eagO9j2iL05wx
lFvcpcMsXmwA4cbPM1M/gWFBfyFgOMgAlwKTs68GR78CxK7CBvMX8H7a1xT6TOqMxVhfOK89147x
3WyhWdP/u3JpFbG2ScPUwjTTBzLflqtUYgAqyY1AD9KD3grHjTLpim/K6rOwlDuIkRqQXdiwtwTR
kSYyB3AFUVRelnNLImll5IGn5VLRhg4dUzDsK+/UQdYcS6VXasdPs1b9dOHN7ud3+npAoqNHgvFT
PJk+QbrE1jJcDsDIcPjf23VsjolT2sZfgPvxVr857r9CzHFNgo6pbWuNrKbULUeZVUSemEWqnaAH
ygdS2XUHbrcuwknSJKg2VC5JEi79WqXGFGsq225fD50+ktOodBP8fWO7SKSJNyq9MW2B5tCrWFxl
ewcvHcsml1TdMrxS2IgUTmPJbvEBKzSG61KABr1JXujdCQx2qDl5adLaZ/9IdmupMayA/qTQYl1E
1ihaCex9It7YiyVcq99rmsz8CaOi1LDrrosP2SxlrpMiMeSFT6XrVpgPDiWpIsdLjEEkteuwJt4n
39fNxBic6X016NoQsJdSISIT0zvdoiTx5qO85YuRLKzX5oznXxWSupo4v3H9RpkZ9gASxn6q+571
9iXS3CaqB7YNne48jLGME9MlRZOWcjq17hk/FV2NpOxJ4fnua96e8mojMYffAxob9jD/Hb6cYjvs
4S+Fg2bKDI2q8XbY9WPnVKt2q6A8C5ePli+OX8KdV9daWLwq7PSy2WWuTB7RuL8AfUFeC3z+nd9a
fqoG9RcJye8TMIbnsiuVNf4KhT6V7InylOSen88XKleXb/hlvNyHP1svP2XityB5fLVu5sJZyxyx
2odaYNg1sFb3j/R/BeKbJ3SO2CsJ4d4YoqE8+jdOz1YonFUy7qeqthzX3YD5Bs/IO54Wq3NsETgx
gq1swSQ4yE0mt6ANKsOTcWCe2RzaQf4aAvkRw9qBUmpNOouSDkj+DTltxQa0sHFjFNRTxPDgpEZZ
NLBOVRDh5GdwrXDcgwAK/G1veggGOBb53BriVDzydDEkZmxEikoIOUVm/bvXWI+SLPEw5dKlT6IK
2aLK0ETPhH0MeCyBdzzIsnuh673/nrNYgRtlljzKCdJejiAMrUSrmRmj78VQY9MXcWMiYFbZoTYc
A5sqC+n517WsPW+r8TnjPjT+lW3zhVpz3ZSLnbHtDrpxSRrTa6yrWrGT3gfp//SluABLta9Yq+fs
dJu2Cd9aF8y5GtAwDbe/T1lB/e7xRm7WrjNahMYEiADAJz587NGqZCtPlBpiTv9GIREobvmtADqV
re5NMcKa4nbvM4jkBnPIIVnfkEHuNn89gyED8f3nF5BwiMztxfKD+g5VZR4/MDRA8y0F/jN0yHZ/
FxPGA4XlsuKe+eH3OEvcbcvzVNojV749yKpOKHXENTyz+e/U7rQIURi6CrLZ5J8cUOZrPM39Yimc
8j4PPUFLrlnxOTeUEnmlOJbXh5DGptgy/2Y5305DFxz85Rk7FI0o0r0MccVdYXWGMzoKoemjGPfd
TJJAbamlVbLIgx+10QmKIDrj2AeHAitYuuNpSEl3Dh7+1IhFhwPk2PNZ38+Y+mhOzBorfzol/nc+
PyfXUcatHrw97SKLIk5YxlyOAJwLPZos7/fNSsBtGaA20NiSw7LI0J6WPzYj1DVoCAQPYuVLi5IO
wyyq31iVlCPZ+z434DDAqG6YH9dSdCdF9A97ky1VDDsrIXxJdj1/1G9DrbHZoclDvO5BE2rk3s/D
RBhawAfzLQs+02GdayLbOiCygILeA7ckFoGqZEkrPWnmuc2+mkYxbXfqRyKaljHwQuh+CpuCCYhJ
poTXb3kDCB9X1gvMV55oTmOVqw+15FcXprw9a016D6Dbze2kVsFTK6qoxMdtnk2iHzOpquVVLPan
lCeuvGKD96Apl8R+jKaYP23JoAiiJDmjqMd1Jz0eW0ddzpWo6zEEisMx+YW56e2MkKGWhqhmlTXk
gPxM/NOl7Azc9sOCQI07I5kwwjIZHfSKRVIf6lC3SAie1a0GLHqrSQvsJHnXoHMMUJl7EC2ozSOZ
6RviRwhExoFQf/EGQ+emeuVkpqsah/xprH5DqJwxnnWZh8rCBG48FPf0q4qX8sIT8c6UKC2jUfkP
MtuyLlDQOChC1jncDt6/OjWOQjQWyUEh+T7per4089Tx2IwKSZihUfzXmi4lEipxGTMADLqaTgZn
GbFvZFnrw18AC/GgcdLFBexkKabkV7vshKU39yFLsV7xvLB42P2cKEE1jXox99umwBpSRTd4Qgd3
CFZi9bKW3FBHYJp1KUqH0WxXj0fueeUzvC9UGWrnXIXWXrs7x/P04isSSEH0cAmGe7T0/Ekq++mx
aGPnQwUjTVOe2soWMNmefPGuDRaTCIr3opPqUpmip9v4lFPmGmgv/Tstn85EtW7uGM7xAgTk/4rM
0Ftgi5UkTXTyEwa6QKQG2x9a6wh6S1qGHaJaVViFV9jXkPHIZofdU+YN/JjHchwtTHwUyMdIgZFN
NRvwjypkyuefq87MpgX5hQ6zFwrYoJk5m/d2w2An8VPitd8SOPvjNbNTlPM+ZjsiLT+AJEd5UgzS
7tudrCQ6GZIfORbujDNZ9zDsoLompUZFJD3pSiDwMuIwe1U5OPBAyUV9Ous6LcqOdWT9WztijYer
TVruzA4RKsrXiNwU53k+Rvm6fNF/QxwwUbQvtscaar9UeZcwm00ZWTlNFCL0e6aS/a1xB0iGVTBH
UA3Dvu2n6MtI5DoctUkUINm1vm82BK4pD+J866gaTUsdHj6z6r5PUU9BdxXFpW9x/pYUtle6dyDJ
MaP9lQ/zZd5EDw9snrDoymCf0ZUykBIghpn231n+oIqHQ1Kpa8i6669tz5JRvnu1p6oEmejjnFrG
nWGTCNYOL5DNceDTptPRGd9Jqk52RpDxmjVGSjr9Gv5lKudLcJ2c4z+c1rXaUsgi2J2EOd4Y4ghg
EOOu6xn3wZ2UsSio9tJoty6ldDLOTbiTRlxY+3EE1cMzYCAO4hGJwLtZA2PO8PNrV/Uj/k9Ushso
t+qHRJXmkuvZ8gCLCSJ73ezogbyAdSt/tIyfu4oood/g1k1x3IsNPR8wN0+44iP+hpmEB/MzDnTW
D2CWEmzyOPt1Ug+9wFSayB0JvEKjAbbL6pmD59xVx1JCLDMhys/L61iY7l2CCFWppnCwZRoiyaMP
YTd+ozJBzSCw3/63t3GgcfAM2JtjcJkzSlY0h7t99NFySJQ+IRTChNVulQ2aHV2I5Eld7S/aODil
hMzXBbCpiFV6xf/6K7iXxakP2rcBMYvi3Ti8NgkwXu/Gi/4kT6Hr4QFkpa7m0Yyno/89jY+RJCVV
Tf/XHTxB6v0XAQB/r3wCWtpGqde+/zczBzZt1Sj0RdtAksPy38vYjHDVwQeFV5I3WfAeDvfmfHs+
Ygp2ljT8YgZ+3ct1ezNnOC/7UQnIjnYgfMCgrAt4JjksLi9QTwZ+G2CEF+pgH96txuIITMtCtfS2
y17+vC9NwGqfrldRSXzik0tSyBNqkgeTJWVL0Aa3yNU/wnOI7IChdwsvVq5f9CwvITpBN2wKTIBQ
S9x+BysG5j1/+wObt+rkedsBSydUqfpvN+xXhd73oZYOq4rfL7Qcq1bQz9CKkCoUTZ/ZOpnkdnw6
WznwQMOxy9I/VghCXUQWJmUrKHUcDynQd8I7E/f5VnQ02u+dMhL+mmr5m3xAX0+yS3+TsPC0+n3F
Oc9O90/4FUvKci9XMwogE/OQp70H1AfiWNbRofRO9Zf5NesQ5IULrec56q7k0UDrIkFxbVhxaI6f
nTM3m8e7Y4RHxFGuFQApN0fITR9lMFaZln8VL6sMVARlzHKbBEIE8am3vHFXQQ1qEH52DE4E8Dn5
qGGMBoNubuEdJ855aWh/LZp/ocKCt68TKXp8PjsyP2+QfVNl18YxVxf+pfgjkF8zSTbGbWAzlYbU
GzvtsiWPqe5NZuVrNOu/rnVr3byf96+iaEMOV05jxCVhy4atkfs+/EPerk0Zv6giF5ynHrGby+iv
bQ6VwBF3GxUjLAhG0kg8aV2ctsmaxn7eSp8jDfPkxqi2z6dLA9gwpqvlzYJ8WBcjotB4KX7SdvcN
kgmFlSxIU/cuEw41YGPk7jmfG1tMfpecz3fJZvACmqHVrARFvQvBuAfGkdnN0sq+bsXOWrcCSI/o
lxIOFdKfhfG0ja8qfO3NhRhEUWlxdCIqoCkbU99mUdqqIzl5e3Du3c1uV0TXt+HmZa5SD0Wi+f7C
G+Nmwr3YxwS8kwbecVLUcjrkQ7aPEJicHw6vcq57W67PzwEqbj+5r+8g1atzchyzbvP+kTj0nrg2
IuIJ9Kms18A0okrDzFqWwB61eYQyT5Dea0taOpDiqFKbJpYyclQcBbLnq6tbDxIpyu5l/2dMbdsC
tphZBdXmLinarxkIiqZmXdErxn1bSquMsZ5aml4tDD5I2AZDNtyjX6d91Fd0TxyHPKXM0RROjgfb
sZGSa24xTxh00hHirUNk1UHgOD72yc5uGMd9KzbGzI5NWpU8PrNwAQNHnRQkeoGHXGKn2xZHBj1o
5FV+AjPTLcFayLtySSf0fRFD9H2Q+kQaFkxpdx5e5teO5+QO/30Z9KICz9CQx+Wsfbc1QUttV2Jb
z6vLNBKtJP7XCTcDnthXTqmK33BMrARaGsKPUPvt6nQV6oHD2giJLcmcKbDoeo2i18lJbPvrnbwb
NkJqJXqaju9HtSQoGE9L5sO6/FPjpsPlxsXdAVrGdFyODaWZzYdEMuL+bgJloAhQNyoDgVJe6X9L
uWZcMm+rSyLuQuyOPaGVO4F+imTZjID3ivrzE9PXIpvNiZ2nZGKV93EwwpHbfGQx3D78jbjdcmrr
RmkE5Hbzkk04YKPv90e6P6yEqcW4h+yDDynWEbDLv4zotD4GKRkQCtLfEKEM01Kf+vDYxcQ+HIHb
Fw8Edf168mMZaFRx8Xc42q2GU5fn1d4p7+4/pyq6fCoD9lKdK/Yonu2XKY0nog1I0AnG97iInVeU
GYqaLArh+JM9vk5MWPBYNdqcHMu6mAJ4UNwxCLCTxA0g29U8V1av3vNievJ9ZFLLXmj92OZsUtE9
LQ3pgT0CwlC0B4IhdZeg28UwiQLPuulA+V8WDO8HK/ow4GpG/Hz5pfGLDGlSSXUUf9zx1iKSO92N
uz/WND0T1z8yT7iRMu9tMezjoXiKYCUF0NmBfx1kAC8St8e713/+JhCrxbz19Mk54x2SD4CYaSU7
+J2FdGBJ1AHfMU0DkTbNaCMGcq97QzHx/PCtXLHxzB13/egKyxiiZsBPlz0SN0YuXr0a7WI0O0MF
GqUY1ZaZSxBSonhZnrgQVfBXGsCOII5AfsnMlZVbF49EYeRTwQszxdeyl7HD3ABaVzuGSl74rt3Q
zW5oXWFZ84Oo7QZeyJJF51esua7BEDGlV3gT6PKDxgR5XeNNDCozWhoKGxNVqt3JKGZFe7xgjNI8
D2lwDrlNo2jnZ+MSNb/i+CeoQjGFJqHeXO4e8tI7A9CQxEG2Fq2jcY1zuJ2AryIkLxAVpSdaUEII
bUXK2ZoaCSgva4l3EmeelRgtuZSYM0x7Macb0dRZFcr7WA36XJvnGROlUI9RUofeVy967X+mGGaU
hIBmsnnDJ/vub4bwMMufGhkeRox4BW7s8uCpbtMkTHimytRqRYzJiQg7s7+VzqPo++B4igphqxGc
WMADvWihrUqp380FyBgmlLYNbmgLRGfYKGSAuwtVWMg8CkeGlytRKsp/kA0GteOeyW2IxC0m/hmk
ZyvEB3OIOpJhqt9faw4ZCqMj4DVzbikbyWvY2bZFdDDSMU8Hlbbj3qTlnhGu/KGkU61gXy71FimT
XSX+8zNxTBgKLdxU3xw1bmAmAM7Zxylx1TUzsHqm96SfA7zMbnN7jEk7/l1pd39pwzlRswggo9qY
eegWQVkucU1B0Ku5usHPpBIpLyo5mTgKJU3WVBkgIppohP1wJXMgNrnLiRCb7OfXDMNibntKBgq4
Ur6q59uBT+clJ17LQBx0k3OVYn+aTxIQlzbzhg37XzLAYxPIp6toIkRLavfHSUxEaxynZC9pMV/l
f/HNSkDLKWJ6wNXUZz+1iA8OS0sk5W4rZBKyo2bbyim9N00wANc025JndwJNoeft9avgWrdY8zCn
ankb21DjBkVUMpijpQKrk7l5gF7OdxFJ1NM4Ve9kw+UTSq0ywrFUBadKSsYx89FRN8dDTlGb6Pf8
rwvEzb1EjsqwRLjJ4IR/De7MVkOm+TBVVSh4EG9H51FBGWgpWelH8J7AwUuBpI3XRJnghzdwhzAY
ZYXEjkr5uufWsqqzVHIjE6VKeeSvY5Z1+penp29mWIDr7JH8YFRwGXfI3SO+V71b/xkwRSAS2UsK
iR8tqiP83VXwnAFp+ypo7sX3J1V88MEfEZANn7T8PD/nlJHV/P2oU3kJLb/JmOhpsayEItNHl9Mc
If3cl5JBbiPwaP+s0tIw0d5Go6OX6D/4rFU9FuIBdn39TYCWtfw3M5MJDYAgHN4z/YsZWcAUD4G0
u1d2X6S94WfKioQNoVMY2boE/s3wZR7J5sfH+YmouINqU9MUFBZCGu1mY1Nvq+O4Xy+iaQbTnde4
Phv0myX6URqsiNIndcUjosEAI8vGA2t53oMS68So2OqFY9tcR8hZIL6rJWHCQFCGqCkmSySitTmi
Da2LoZokA+J5wIv6e5C8kTvwCNZDmVFq3RtBjmFmgIEzj2NVSvtx3HGRRfKhMU9zmjbHmFJR1Qay
2dBoxNtN9h7tMdE4MaBN8KX8ABXbnxDvRx/GEeG9IB5OKh7moiXT/Oiq7EYBWDu8/Zv2YbXCwxfi
Ajh5o3eSI+vkKIb1Q+y6z9Vo/k/uO+smxLDPcoI2VXOg9spPmyAv+kAIatVebZ6QMMTzFxIM6yiP
Cnpk+Np1TfW17hex7ZxzgTlK66emDukgF0KwwizKfBayzBy7YfubL/2vRe7pBYw77I4bnpJJhtWI
7V/JiVmoTz3CUpQHy2pr60wAZqvzAUE9f4QaJ4H7kvLVl1/+IDPdCcIHJYkiUwKOpNiMSYLAKjmj
m9L5Mi6vsbYxxH7lGyyZb4U9QuzOUZEz7Cwd9PWqA1wfG8emsQRB41Gcu47SG5Xs0FkxchuWMSh/
8Y256WZ4whkPx3Y+IbsiAXE8qEsqbR7ZsnGdO/IG2xk1hy7xosYZ9pAJg7GD+wU3LZj2JGDkMwng
fnuJuNCXo3fum/TavKqtmiMvHqhWP+V1EGWIgBmhcss1JZAVXroBNlj2ZTCcBYmPR0H6dwhwICem
8ipLaw5AC1HD3KvHE1e+KYwzhIgPhuW+kRuClCwK/Zu9HHNRedYsofgA4zpNVe3q2rKqbBtBx+ZO
TOVopSeCtO2zdUFnQwEZK+ppgujfP9dM3tziTxWQkLZpKYwZd6uvTBNV1ppDTmQO2GJoZ/Fg8YjZ
RFtzpS4uE7KfvTzka202VG33gHKH6gJ1SXc+tmTW1CszqUSJ471fGJWmBEWwHjbMNtTni4oY5CEp
Cnjjk2CEp2VFH2gynx9EYgzRZ61k9JcR9m0lKfKPS8gf83cYzhC6dP+6W/02zdjFVT54GLE/527a
rKK/ZPDnlHNXwdwiM5cLmvjsdfGQhXQ4tNkWRcpLl6ddKnnELSnbgHCKXQ2lG3/DMUgNCpAPK7Bq
wzZG0i8kOvqtdYQGWLVaUPxHl/+u6C/HQH8brSdItr49N4naf2jUzrhppyoJRQRc+yI2ttRy9Rep
PkLwaT/23ycSyNhOoe+F+UJGqr3WhXejQFWMEE5GC8h6F5gT0Ngi9kIqtpzoYyUuDzU36MncvWb5
GswXQpF+o7V3Ee/IAQGVyN0xzq8/2TX8Ql7Z1yAK5PwdWwYpgt39Rnj3Fst76JBguGYMDzkcipio
EML1nIyYrg/kJ+ia8DeVSDmKQ2SiwX46xjzSaOv5dQlFr4IMZqoCnf6mr6LilWam+d5q7G1yy+zs
JIQt2mbwmjuR/hyVcJACizP0SdhR7vZOlrF6g9uCZh0AxM8F2KcMzhIZiBI01KhKJKXEeUermjM6
YZDyUGEtRuR77DffWL3DA9uwPcygESai9Hz7xFVBQtdCnMQfRqVKcF6+OE2cYp6RqMsnPPRsH0Kd
miQIZahuniXU+K6CJGbq0DJb05R+Aiz/nbJOr2jjFj4kPCvt3jCxCpRcHjFzvg5q+oiR96kSvgW7
6j21ggcx9CbOljnRywsqo9j2FYEuR9dw8/FjWWl5vYM+TZfagvEagBcqOqKbhVFxt3y50pHr3gPb
5qof72ykZ4lTZaPFMLPCzJ2lN1/6m/tKmXTCKFqeK4NUyfOj1u5Bi2s0LTei3FayVUP3yr8byTFh
0mtWrN2q7m1EYA46HTWKfpsc8KzRdzBNfy7IkrMKdF2tBWe54PLFgGkdV/j7pxGLWWKT7JwNFAsS
m7KCYH8ufEoqEvzIb73+uY7KuSeQ9i+kEtFrcsyVwN9sJbKsUi7Bsg1upH1GApQePcZteSXUxx0l
MiT7RH+/fMQtgXQ0jIly2lBfL8oM/CahQA2ACVsIBT6LLkjlfAbJc97NMiEIVadW73KTBaEnui+R
Afm3MZ6RupF7Fl+7s22Hu7sRHCmpVtSQDzOZ0KRczsSupppM9j21Rck4kFdrK586VsnX8dYenl3R
YsKn5jn0EQLOt1fAtg2oL9DjjZclu4mNfl8wPPRGglh/bvqF1MGnQ2vshC+JGsvTgJafZ+kskbse
FtTF6KGmjc3rXn8zgthQq73eeip8Io+E5PRUNQbn8p2446IEsW5IuQQHNmvusig8QCfUlR0FYiMI
xt9kwrQAwpmt/i4UqKUAhWEgDvr3gNayiGjXGd++oGZPGTq21471qGY2e7wNeg2ugsFom1p3cArU
zdDMu4wH1EcMhacA5oS7wgSc4+seddmFYW6TsMFMpYswThBUfUdURzaKpP1dY4K4B8ng+MtGcKOk
lfWkA0gXqUaiVJBABSERbzJzEgPd3E3eSipIH9zsvMg2BvZYvrQ+BgHKiviRAiYVdHHk9h48uCCN
6k5u8tKloCTciHaD1I4Z66fN3+5nDEzE7PcYMYRxG5f6zlqUtxaG5+JPsV80GdHxBEcyXcxv8l8a
zpfsD8w3259fKNMflCs4o4W7BB16mTxAsQ7sXSDo5693zoOic1a7Kus04UTWJHNRQBW4F66UPfRX
j/2Tki5dEiICi/bNthLIGXLeOdVk5tD7lfqonsG7wq53vEeZ3VcsSRUwtn1+ZSrMLKYDsVIpTzev
ZU5iT/HeEiAsdscr3RCb1o/crL0rTc0848IN3hx295tglabn5w6YV0ZzfFdbNHXpZesysyUJNVwn
Jjz7pK2UK+sTe/uNwFTNrS23TedKgy2YYNxcQXEGVUQuD6SS4OdFZV7IMP5/grqQZp8dU3mB3nZ+
d9EW70kDa3g15TNmGQH68RN/6sV6wGhgU5fq/E+AUT7aEqcg0xhcJFKZKvwn5Wfofcz3R64j/Ik1
m6Igi21iQkeKRlQgzmeQWcTxF+B7Utmgx2l2/4cv6P27+1V25efKyjXA2RMmbk3Ln47QnGaF6rj3
5Dw4SU8RJkENmAR5Z6e9qILF6sXhkb0WFmjP/WT/a5LPMrrIc7bb50OXmZrP4/UPHnTDy3Ya9eLc
ijBe5C8MbOQkHl2TQL9tHV4qBwvM39t9cg+objkqw9Nf0TZGcbTiukzy954gNJjObuSAH/33BuVY
r3gFBsOTKHBeLZ3xIZVJHTdpXsDTQDlbiPWYr5njvppF5W40eUWvGsOuowMWNyy2dCdEz352//2L
N1S/Uz8wxqcYGoU7kt0m/pwjOk8MaWVQhEhwhWUtX2SiVEor88tPkIKDfRKlhzaTmiDa1t/YGno3
t++APys3GBbDWmdRJR86z08vL1Jc8SY1p4VGxwUFetEDMZhd+AQPOufEwJ9gWP1KwkQ7y8YyNoPi
lECw+umDuA4wdPeFa8CttzHkNEzSsul2xNUyPG5PyeTYBUA4yQC/R+e9/WWej5qrbvHabLiLcuQN
2NDdi9Cdg9DVXzgqumN6wZnsZpp6JfM867/M2uLpAbbk6DGph7zULlRIUdcCmuhN2ZfFdjTX47zb
neaO3fbYOuykYc824JAilmTixZoMQtP/JGBH+pHAVieNwgS4xX5Mc85j6yfabyrV/QIO6hGO08aW
gf0eosN+7R0i0CzPTie+BzNprzjdcbhrrUZiUcvdNyCc5a3hqqgefUFSBFoRh6OQKnO1sFCNIUdP
5t28uuJ6qvP/p69+tkW6dyftXw++KeHsqhgKAa0k+MaHUXDdVab373ic6nVOClZrlxVqYjIaoYHp
xCr68ZixTz73QPa6X0Jv1QrkVenn+k2d3Swx3ioRH52aGkewJxJCoTMPUBLUVdfgeQPvqMF6swu0
3IOV9+b5bNd2QjfuxGRvGsgwVOzPEMcbsgU/JYYUvtjkacqCtLUUq6wbdmCCrWiIG7gj02Zntw94
L88aAsUmt/c5h6wv+l+ezNk8WlrWc3FDlmFvx0MvBwEaFYH3c3d/nTa/R0PkF8tQwHsty34eXpJd
ELfYH53VL5kjRnAZV1dPQp89vRZDaXaad7kSvfZqCkNkt5b6goBmLOgNTleHUOKaNFXOt+gS8Rxj
n52Cs3xtdLtKNugfSSiZta7LztR2defxWX8uA1X+Jc/qXw9wEjCnrvj7GFqi1JefWGtGKXHkRDVk
bus4cLUf9o+xAs7rJ+djNKFyEPJJeNlBYtRFC0kPXMBEG13OUdVg/BAwgdx0T1Ya1dKE6dyCA1dv
XkTo3ufdrp266XTbz4caEn9lNcF3ZrQwx8i7ACFQLJx5okUz9gw5PwNMhbWNSCzPZKqY6hIUnFY+
t9oU9mNk4J48boZlkzF0RJFRlAgb60/Iz9NFjvesHN++WdqfX815AoiYgvUobYKT/HSVE4PHIbvr
yMyrZPCBd3zpYLVWdow+9z0D7n/vjo8dDGJH+L2eeH4qgauPJbVXx8Yu1AB0kbxjXfxmSzF9jjrr
LXxsecdz/yBPCK404r1Ah+QpQVWJD+F59dW9PZHtfTAfTpSByv58p2TkZOgPPhtSddRh5cyfM3RY
uvIwvVf8WNfycDMBOhk4Y+zj6TJ9JY04QGVISXRJIGizUz9bSOlHzMrooQQX2qcA5ptmKUMaK3SW
daDk3qG1BdnXxQIFq/pINNlBn56kWSyJnr3RoCQWRHZapFeDR8MLQZorhy79ZH8iigAD9DPkDAKJ
9lN1Upjj56puTOl2E9y+9eoZxQsBqQ02yun6q+9rL6Q8w/03mPrFpkdJiHgbaN8h2CVtOelI+yLC
MG/hKsPJTtM6yH1iw7OGOQqQXSx2PXSaUG/r9DeUjQNgiY38Zz0W9JIuSE8iYgztVwC6Pmz+DLJ9
4P/sdw+juPPiGOWweaQUiCnNiBLgP0TWByolAFRyvyEs22Y0fYcyvLWDKWPIdI+I8WLX8JYb7kB4
wqbyDokiq1k0FBsiV/j2yyRq+VwRJhqJwzkVRDPMuXVRXtaFY+lgiJ8E27CK5XpS+FFMR6I7Tzzf
yIBRxznXGNiUYKxBAR4UZOD9kGxcOZ7lOyxCMHVsDJs73CfHQDMrDQV6kcI34m2bUHBkRBsAOUbu
AYbnzX2stq0FkDz3lLS1wiBMRImsyB5FyltRfq+iw49oO8xsn8WXelZbZAGTqOmeFnKKtTV3ueCr
TREpARaTkYDgQ7/WrUq4ryxoMm60fLtiu2RXJWuRMDEn97sO9O+JWpr69SvnmFXIe95l/2sqXE0L
GrtwynqgYFxn7B1tw7iZSItiUhP5/8iqqrWSxVPXvl6mEHJGW91JZ2WGSkYQp8bsg18/3ja/dwp6
8weIK33faqQ5vmav9PqdeBl2X27zN2F7CrWVXENS1BmDuDvO/9LMkxjSKF39Qk5VNMXowkohH19D
VVQ+qe97hrzFiLa7V/jJ2+sxEISGhj5wLXGaAlfxD0EsHoODfiY/K9isZzQjLf8OxzQWQZ8TQLXV
tXWXRUjXbG//pwkvYRIqWqLg/4vPEU+/8WjqNucUGPe1xZfYpMwr/Ma1KxpFiqhRX0CIpcGV7EIo
rmz+cwyjLkf4wRfoeYq2/1M7IGeuWCP6PWe0lCRizKlHf1WqKAJa53pkjpKphhizO7hU1Tbq2s0h
lqPf1T4nOQItznkjNF/IgUtJ+zSMpVrHhTgsZa7YLa2JOltiN4CxrgDZyjkvvYMcEKP6lLHkkqef
MRB28PUECcUalaLbP7tVJGb1nO+Yj1pMDuHbh5iB24stTzIGht6ojEnht+z75ZvMBJ0kGxUzExMP
xdcoUEgwI+7gStd6qsjA+UI8B/JNp/4PPRENocsXoszxiStiGqFEX+sdwNNdaJSXNaOrPs37gVji
x39MgRwYgiQvBlMxBiIMJtW05wkqmJ/aRydDDprPnJdE7685t0Wfo3H+y2RJol6gwXei7WZYqQGW
UOuNeQn/Yay0vP/i4tLL80iAxr99A8JJEiMy4LEEgAv14gslTGB06/jqmT8ix66sSPJpMpIDq8WA
O0Yo/Ndu+ylEY5/3aJDkohnIj6s5qoD/ZLFhvYCfc79GNakU8iQGfkHdgCubyPlF0A4mYnRLCPLc
du7b1msx1rmH8M8vQmizh11UmN3QMaGt1NcK3ObmkpcSQ+9zYOjJQqg6T4cPkppKbhZGInZAutvk
VEEXNlP0V1s6120Bd+ovbr3bTDbeikb9eZkXGuRKIwBQ9kpJyQt0NReqmdpDAGpBbVmCZOuf1MeE
ffY3hRZ3LUGCl7wJ3nV08z8Ba33MrcIJxaYDCPDu8H2nkYx1ONr7/kCHhSvqwDfmSRCqYe1ZlBZs
1jc4XXmZNVrOYg3tjIDwdXGoNerquO4GK3sQDy2TEncClzYZ3X48DQQLdwJ6C+dGHg7JKmjskW5w
Z/HvvBnvMGoWJENUlRXnfj7kwvoJO19jIXuPPwIjt8hJ8J/PUUWjgWueh9cOqiOzBV2d7W1tVaKV
IJHGN+n8dnQ7HedyLwZ7cyYWNJiDByiZpDDEKB/gmvNPIftbGBWTphmd/Ud3i6GnTeZiNlLYpj7i
uyfHiM4LomOnNJXoVQxxaohQygii0w4Y2122TmAF1WIl0KwETwsqZXigNVASrhF+6Q5hjFKsfIIq
mJs3TLtTgOsedjNor+WlnNfQ1t94DAt+OWrlSZZIAr2IDZzmrD0hmL8ZASB+8O3NSHxVD2s237rO
QFZ+LLUUJWVMrE/ftzVfrY/Xf+pR5u6Ts+AFS9xIYvPxrrdIBXIZO6oZ5RV6+tAFtxCxoU7l6M8t
WYsvUlIVuUDOjauiLSr/VAXsd1vUq2OzKq5f4khqHz5I7urDYe06kS3fs0NKN1Tonyuobu96392y
tGBRhMxElGjPINrFJSkZhIUYHvTx0N4J4P228mPEGQQ+Nk9Qa46jd6u1Ru45OHmYCxv65MspbLW9
yV4CJ1TSHgiy/wZwIqwfOrwwfEpNLmvijSoDCkrI0eAyw1RUskllYbByNtgHom6045iDK/7pdZjn
3rYheoaHTbACOa+lBPCQi98UTF1L8LT6iBgG48enlwq2j+o+9iPQSocZztEpkCfg2W8U7daSv6UO
mYAtw26I/cH0733wnKzeKJCptrRVTXmmqCdxOIBILF8ICgED5RjdFXgUe/nzfTLd8nc//DnXYeQe
nlHKJBy4KiWlihuWZQr0UgEUoFy+uLcfxEoBHeAU4tafmvKwh8gGXCRKcm/ExchK7AUS7XBNZDXI
IPa6qp5oPOOqddBfrwKmHXu0xhWZRQkVJv5h/MOG7W+FV/zjlBZQlET/oiflpFK5BJV7YFdh3BPA
DPmMvy9DtcyGoTE+5GMoSZY3BX4VP9UiOwoWp5pUwyNPm36aSbnhEA1cUmiy/3T5tRKmvvFqMxR4
5Mh9zLRVyyAG+TQSXbv42v9oUlWrBV0DFGSPJJ9TLbYfDhfSRCyh2Gk55Zqhca4mxqLPQpQbH4vA
NdczTPxGv81HBEjTBSbYAqw6c4wulWdMxrUAyU98IQxT+M58zqEdnrnfvMy8ZWUP6YHlbXyq9qWM
5wBCZ7B3lct+ngBQc8yW8hainz8zOeeRV33YQ2+bYc0yvpuZ5I7qR/9LoPMY5JHaby86I3Xr4Ckp
UYA+QgY2iaskDCZ6uj7PVhBUfDgxu9Ya+1q4TIuU/T0J2cb3OOIf2wJX408V3S4gZfmLKiq9m/SK
9sE+dWQYJgEnMI2gOKnpnr/dYLalIhjGu/DR1g5T+Re26pkHMqq4eEnBqBnAIsXROdYOKsW791AC
epwc0+yohdgSTK7+FmaomoxzlXEIl5dQ0cy2TkqN9fbfknfYLHRdC8pKOYFkeGZCoO9vbBeRY/JF
vx3cq1h+6v2GqYgIFTYn77okCxoVHJ1b7SY76LOA48+iUedt9PIRrisRR6Z0EBYeEHvpdVoohdYL
Qboc7fbQo6Rxan1o/2u86Ga33DyAQWOoIb6qLLIl35cEIHix4r/tzbYS/PpEwEt4WTiAHdgy5kvx
+thnqy00Vd/V8rHf2wxW8e4s5R4ZgeAuaOs8tvHaPs8S0jpQjB6xor3G97jpLNjIJbfiTR8fWqWX
KElSrP45Sp8O01zc10R5uUOgDjd8+jSr18QOhz9rx8UKQB7lIA+5dYu8Vtwjqfu8R7RcpC8a8zfK
3IXXkJ8Y+ILc8JzwBb5mMQPy53HL9JTFALqj9vzXilBr3PbFowdr19rnsRIkudz4w+FCGqv9j/07
LRsUqSYhzHczvX50tv9nFqzlBswjQBD8u4m6eyT5kXXhJHHEvTF/bZQvH9M7hDaW6zE9/9Dxw1nD
dyfLe4av6GQjUzpQeMRm/UEDlhqI0baLE7dXnvM/GNdyEsff3FNdaLOM1cAOds7KolsBlRKVMtJE
C2ZPD/CVoxN/E3zIR0pZ1StQn0R75ZYQMLmg+7HHkfjghYAWRaCtf22mRMlXtZjeryYb9qqEY0pK
xpj5ItVGhJZSfeq26TPn3p6v6zurixPVub6t6uZs7j1Sv1vMk2OOezG3B2p6YbXH950AVM9zgDqD
+uMoEKmPFF5StWqJ4nwxBoj4iFh/h30lCkLskIHkOakaB5jsfO+yDa46qRqJCfZGCqqsTkt22LF8
lZfO9iwXrfMNnC7vDcHhE1Z0d9Zr6bo9Y/8QvM+zDBcy/Db51QjbCoHYtjwWoEAg9nA0p/wiItw4
j+b+B/kp4o8lgF0XdUxLwUCm1vU4IHChwJ9eDXH7P/7dkKTgsoaayyOrHoR9vjG62xMI1JxTWe9h
uvC8mAXiMGl/V7M0f/wLQBu1JvYHIab0+0CrdZ6OOAPfF97Rfb+eTLqi76qj26YOVTe50gbVUw15
qhHqinWgh8O/oqTgJ7WWYmo6RNlseKqYbKSQmH2ZWS9FFWwbqkcDP83cNt05GQpRSA5/BIRun1vT
A93eEdmpsqhc/ydeQZikiQ+MvWWC7D6yCtqY5LARdpI2zdi7sgJQQkl5StAeYRB7MVS2JbDlynbw
xOzNaxm4OSbESkIj4CsQIw3RN2IqbOA0XY7/mBjuBMhASFHYhGLGEd88BygF38tDAFjlL4p1PPNw
dvYnh5dD64z1auZieqB698ti/i4tidpg2A4ozxav+CIZIXHgK7qERqK7IcFN+usvFSe6l368UWhk
PKecJnSNaP3waXxO19m3ua4IXFLHNZEtKRuY4+ZTFYLE0Mawg/LWaz7t7nHPa3JVfX2PbDBfec6d
lhJWN11SdEQLm0y8DGbS9y5Ll+XxR8idsyJ6rr5l2+N3lMFqYUREx6Iwo00kC3So8njdulPgF/db
EwD3HNHvNUs/dAl0gYqeM0wtMtWjlSIeQfAfERnt+bbCOpOmEejUgCkasqKlfBfd5ma0d9R25v2w
9sgjn9Bpo/PMUi7CByNo7R+JFNxa5aIZFTsrCL7xixF34TuxaoNz5IF64vzoX8WB7i8J79RrXX67
ThqdS/Hr2vGebPrY7N2u7R6BvmWA7LMP4qV6smjDl9WdGs4QJJnZV/sKohitczrxsP1/ErF5C3Y6
u49KOloq9Nw9Xa9Ij2S4Fl62NcA6lVobPNQMc9+r2DwMu0nhQE+eQU34gdd2Keja9LVUk//f8zOs
cEmUoZoX/ySj9QcQyHQRvpkmY6qTyx2+cCS5322ldvaEXFrZvrHBlN9EsF9N+xXaoQRb9DNJAt2+
6xwLdaU2zaY6jdTXdG1Z82FJUkCPNGTph3LYnTpNeCYwBo/Fzi3r3nR7Sgn1LNG5d+qEOZFKoCao
6946wNkRm5RbiLt6p/YkR8bmLaewoyZnbfAv/h972JFvXcqijRVbhhL6M24UC4R7t0W1eDngmxAz
TkVdA8965vBaP2GbiX3WsK7Uqsz+ZJFgIprYkghx6IUtVIaf7BXJA4gLw+OSYuWVnTErkC+UXVo1
WcF1ICiP3ij/Zu+WtzVRhHpBjmPv15DG6Pr+RF6+gMfOSqrau9Oq+Ba2v7u6ibR/puvOzk3reVg9
X7LWkNCkiR2GSgWrg164yDbp4eyHXT1wzEgrHNtvr7OhiVKOKBcA7vDVOpQ+Z2F0jstHWml3UABP
Dn81zOP9MvVWUaFF22GhFIuKm+jTMRfjp+jEBoDGdhpzvbK4/AASG+bwoorvj8aoUPOfM1FrLxr5
30CLcOw4fl1TuMDTZnyI2ic6msRAviT1OHYF2NLnmi1eTqF+XPmI300DOUTOPOu91BfNELk64fq7
pq9/3lNdltf6Vu7+Y84kYRzBz21Z2r4Fkss+oLutrvmeW3UAIiXzqxsQOZNYc2bf8ynQvZiRx9EU
UY8EYku5/kQknlxC+vLbRSq7ItkoPfyt9pHIbEI7317jVXh4L4ReqG9uzpoa2AfgoO2UBxNZ18kg
338iBU7PeYtdI8Q7TrgICwDgoGZD9WYL7Y0TImmw1RTU1wD9xgEwonmbZ1Qh14vF6VJuXlOxi0Fp
Xj8K59rnXbn3QKQdkiamEa1pvwxW5mQcWOh+szTdFBjC7RCSFK4Wwlsln3tRCb1GRYXV/8Ei5Qk4
jIkt5KhxQryiOSm0V1GfpxMxKjgHbZzw/gzHrhQ2953Y0M9DGTW1ZP0a5U2hUAyFxmTejSuvdOHo
SuzI0Eg/s/quf8Qx7kP0kCZLVh9dEBc0xvBsdGK2KD4og4fE5KAwA1Syg+p35TSwxJ+e6o+NMlj+
9WbBMrzsYtzOgB4datSjnvCabB0+bVLPxxCmHAjAouj6P/HhXUxtKzQpHSZ/Ff/6GubKtDnEb2GY
CPRStCT5+hFoSeRYwJIZr+V4FwAbIj9jDaGF/mwAohLpaAzWeN3K6pRzDVpKhT2VOYXdYsgQTh7i
POAdrxobo0AJjxEkG6OtakSWCoHxvgzlt2RuKNIpMiaDRQXFpISaW2BwZr5l2N1R0vqGt8aojQcg
CYQ/hIwo6fst2Kxy2oSh1lBUE3CpIrbJu79LLpauyC/66fty9qxb3uPetDOTAvEtxp7wXsxhoHSR
7h8Ki6Ms7gfRLSjH+lRDZBnYBypKaXU1MLFcGO2WaQ42sW7ERy7dm5ATPx2one8civLkmi6uwnxn
khZtMwoltS7ruTK+5eJO1aPJwx8jYL0M7Epm8IG7GVhRKpdmXyc9Xv65tVxPpUSdyJWR92HmwBPc
KV1yKCWhxFOUp3ob6DmRtIrMPd4p/XZO/Sw8hyxxtRIJIdvn5bfgpFJZ7ihZY1pJSI9LrPv4itXt
9ltyTDkFYm9UvWRdN/g7jf3qxP81sDCemMOA6aXVwVLhrca2fk+GdL2KshhGdyOBuiOEp/0krxVW
VGXeBQ6QrrwrP186v6RmSdNUPXAUXGROl6q2PID1JbZ2RgC/YctUcD+ftkN2IaIsFxYR0E0yf+42
H9tGomnjFpGya6KlKj7CkJzpEiZjGtnQiY3Ux1wBoxrgQAZuugAGml4aYJv9J5gTtZQzV8yrYr60
l1s6AIAiYj4poI/57Qc6ktI4kZ8ba0x0CjQip185yB8IzpmPK/tvIQZkQaXChXjYAKRVwl4DSs0s
rMa4Z1hnO6RNFkVgucID5tFwcP0mQ0/fOmUrPQdFIX7JmKqf9D36abpsVDd5KIpLmcwMe5/f58v8
T+ODzvHY1Ww95HDLIX2E5bMOzj/UeGQe7cRCUWqIHdNgnWIQ1qb01JzD4FqrJPq0WYJDDxFQcbdS
lRg3izw2m56LigcF/Pl+PPo+HU4e3dHhymqXbcIdH8WyvSreOyzQAUf+lJI+WZFVrhEt4oMCyoE5
BkJbHkX/z30bL80tpYI30Pq9Woj0HzeMmScIlFzXdwDGxI85OGpMH0kTUZD8/yBwpI1uxn71H7gQ
O6jDijUfno4V+TpyUorOexQuy9vZ4gBqfeAbR05/x3yrb3DRcTAIEVfnvqK+aXC4Vq20e6qPrGoq
0q8f4kTwmlL6sWGsVxXvUrOhZ9JID6h0EGmqDV0+UiPAOswZLHjqKelQM0OclOr1i5xZ8Tm+XXJX
5qZn2kidM6RmxQ6Lb5GCXfDLKbUftduP03qyBUKsZWyj0/xnjAms0b3863luyKoVW05p4Cd8KgMX
JScwTLlJkdvXg7wvHJQUTSZjdf5Zc58Kkiz+XIAzC6mUb838sKf3txg7jw99JaxeujwX75gtNuSX
TGyMzcNV0XU1/3JRW1p1uSEMOsBKLh0e1qNnMdGC1NfUckvuWra4BVIUI45lCAyp93o8/TvGlabb
1Es1336cltTiuqbt8DGsjwvfsKO0C9IU7eta4JQHN9Q9Dc2uX0xq85n1t93A01iSJH1E6C2d7joq
87QyNQoCJ3RBB1GNTTaYxRm6QW0nnK6nHvHkbMoycrFUkX+FSAyINtt8FuTqNxa8EV7uTyhdh3ip
TC+hZFMbIpuYyxYJYSCwQ0iBiahv6Yi2ZW8bJNtO+Z6ByxWBSkTBaq4qjJYHwm1RMS0ii0JATy0n
HA0ymoXfOvzokeHz14xMBbef5+PDm63oLgW1rEYdioRH6+a3uqpiIWs7UB+fApIv5Zdya0MoHRBP
JlfVc5T84U2Q8VJJlHTRPCWiy96cg57G8cZl1iOfHzcbxmYlxK/BDAZ/m5S4jJmszlWmghckdzqR
pw9We1Q3tPt9KBnlJvKYf2p78H2I855Dh+dWTkpQ5NwBASCpvRr5JBZO7m14zzovlpkocikiOMIj
8m4inuifmHobXRYTBuxAPe6CoA0V7wNc9aixsSe4Im7EHwgvVARcZu+C3KsnMA5TjQ9LLuG9vxLa
zXzfFJZTKqsf4YczSiLZSCnR2336ZYaQyVIl+2jNor0Zh4GNVSwpO5gX2GbK3sWKEkiMDj3gY5+A
LCd4F1z9/X/SY1n+zBDio9CpKJVlW+8+Rsx4LUSndIdv+ptA74btWY/paXy4wvLDHuiLMrInbUbL
MZBC+BGkf5ewqIYlsTfSyqjhhiACuuqjemBP4/KRRQ4bec992kNg/PUTzMzj24offt93TFnwEn0L
aPsuwTQgv62fZ6yuwHyb/rngGBpqanWUn6n1hG/PbL9TV8oYePToUiJjuVZt/5IjKgByKOYUTB2L
1b0aKbHi9+ShHAZ542F2AWh4MqpXkm63FEXiEvdooI+76rWAPKiSwycuicHJEg2k8ugfU1rKakfR
Znv/UllFLYQuxLjleK5goA90Kt3e0IuGtGM+bKkztWdh2LDEWSTIq30xaKGXc4UFmr4c0t07x02b
p/ZSpoaqPwG/WgS+EFVUbBWFGzINzeYbX0Ys/xAjGpCDDOaNvDl08JhM0iCvvP4jKCNodcjBrCu3
iycUES/CQoZ1dcsjsEEtQlg7j8xGHZP4GOPQhhVDqK+iWujtH9g5enZvun8e5IEZxVfV/5rIdxoy
hs9imOm1RhiKyoym9rp90c9eosIgiN+OM4kQTnEujd9/yho84aI1MJnxRqeX3Euco4g2OH0SA8k9
QWmqxbxie/JSZz1FsN9ODNFvixmRu0EgurBXzu7igUkq94SP2EYqZhkGaGEK4ah5cUbunNHNDu+4
weHLokMf1kksFGKDXtOheb2Z7G0+MnhVlx9OlvAnwEqxX7Xr56MDCxWtreeOkG8jeruig2u+QOCY
GUdw00dUtDeed5dW6Z8v2GLPEFFYH4cJBLsOI590MwxU9JW9joM7gf/pcFXy8QNG74tzGIGXycpU
zm7QZbCkjmudD677v/3cGwUhHDSc/XoIUK/5tq2aebXPzQ/lOX3I1sHjb1SiJ3qzIyulXOQZvXQu
YAWrlZOh65uJMaOKIxLqUcdmTgo3svBkLrqQrGdVxuh0iN9q8bnA7EKjFuuJKPelj5C2SsVUfctI
pBQawWwZ4px/7n5hnILVQHUxxRWS5XOTLyemtZxS/570kUbeVsyOq/5e3u6HTfsu74XwMJ84upBR
6VpnY713X8YM84xYcyJx6RQP3IaYEQS2Dp0De9xMInatExaz7jQe+Re5t+knDTnKLZc+3QN9TbXf
P8nURj8PEhU/YSu4rC7/1+Dsium/Pv9izERV7YKCyv6N9TcdAFRlNBxLbq2Pnmwo6qxOkveOWgBF
p/PZDT0V2NzDme9JmKuR0bvMtxCogwKfpU0YWpCiGrq09glUvz/YsOYyDVz7s6bACAU2ngEuCF2S
Je4ffp5N15nO+kSfaK5ZMJud5YVJFnDGaMHV4U1YMXs6NMGU6yPdn29xeoPNz96ewS+J9hioc/KS
U5uSxMdvanDQX6HfIlur9STgdnvhrJIPoESDWFLEUZ6G4bOe8Vz2nTrTo2yQ5y0CYwkjzxOOvRgU
p9Mp2thswl5n/6Xn+QQijD9iX3VZfQPJlwadSbRmfkyGtv33YignznUaxpePEAZJ/3iZTPNo4ASy
LpgjWsj9NqkLEJqi6tbs8xHSxihRVSkTVE/VR4Jvj4AsgDm/Tr2JkCCymhmtagvWTb0VoUcWOj6k
YCy/ekinMMmfWzs7bWVg2z9wUpjesW2HWRjUcNhvPjIZVJSD8qmB2bJp2UNspvXXZnUmTUsqtzYU
8Sa/p7HstZXjJOQQoelcqUvEiVmqckggmMVFaaKe96HDo9KbM7EfCR9Cg9mRbo71+A8d+RjdSm1J
A8k7ReZAYs6NkPC/ONm18Ycok5XEqEpLUxtvdhV03fyimx4dKzhMPYU9Ep+GfPU3AXfgCBcbnnNh
yl7n4jUo2hBIXNBwYQkrfcGr9wbkgYkAAUhEW+uJU3YCLEKSjjUahKql8jKGs4WJXPd+McId53zs
lJvjJWU3heEXCsTBVwUAg4MUrfkpE+ciXMOO80PpFuyPLJIqiPCORG2yIoaroxmkiSgCXNV8H30M
xZt0N29AljKBoBOJi5e5SndD/t1phGoVMxTC2Gfo14X69XE86WSuFKvexxmy6DLLrSFv1k5gsLPu
lO/Oouin0Na416QxNlCS1um113PvPM3nSa2wlSzXfI23OJGF3ncCPBc4O6pRsH/1IZ9wdWxoBfw2
Pj1lQIwgSPcFEh2HxIWA8q3QQl0cWc88qrU52r/QRJZ7iYiMTIoctUoXvLtrAFTGEu02Btko5Lg1
BwQO7X6dhOnrcEjYC0cB223N2GEKSjZetrw8M5Kp0gehMAmKDPBAd5V8hbOKAfkwvrKk9J9QEkGc
n7aw6aAEHx2t+wxJoLy9Lm777+20B+WPaYNVl4JXO2UulKp8bUBaguFVd0X1/BFtFzklyARya+C+
4nr0O6p7qAn8lDIfVasUzHIbI2y5skB8BJG5Xuyn50DQqqpG6dDI3qrmK6DUmzzec22saxg8YQw1
ZIMVkDIMw/4CmHzUnyczLCCI4kkQPdTtTFbYKWlgNaVN6tyZjYaAhOgNMeI923/UB0T/3ozD0ijL
9fpadufOeduvMifGWmYI06avFd3+xOjdLbg+eE3QcZapHIIIwplnOHuJgt4jcOmZDCc0MVW7pnCD
qf9uuiXAosojD6P7DYEYvyqCUkzTmOxAU5eJv7LvDqJ4xifyr3mwLe+r4jrXAnaF4xGj5RuP8hxF
xDt0dxB80LcNs3HaxHM8cNKiv5G3eNZJqTM2Ukgotr/rP3HUzzty21Lg4k/fRgg/3XFA0b3nrP8O
d0zWsQMs3wPvbdyWostwHicBt/TjVzro7Eku2W5bNpbbrG1tqx0hDZnwdQmdfvx7sCAMgMvZTFWF
L9bDPy8beN/mSpjf81dr48hMg4bne2smmK4FzXu4JNwYh+8HXkMsJXSMfR9Y7v97+fspTQArsjKB
l4b6Mc+/MUzUQTJ23IRC10TB0q0DG7g86PJw9PoDMdZyBw3Vl/U0XUrRrekZdb/x3ubHmVX9hhh7
jckj6SZmrESIjWQLp2xghzCfNSbdO298wB/Q41pBA/r4YOg5R5i2Dr7aG4Pujx71e79wAIYZugsJ
kX4dTwxbrD7qU9TonfxaK+D2BFbzH5tjqCfyBqQ/nAtpc15w5Lh2BVr+fov5Q8qztOkjf3nFVF6H
d+BW/6k35KPTJtTg9cz+2zfrN1T9HUPtVlgooaZ+5ETEFmJuzQzIXcxwrfpmusAeUaBE3klZAjMo
Eot2yReM/X5PyhyRJNCtpDgocoqQ/bt0R/FHM79Ah964/Sz0/UoQ4f84aFoEmPgaxNHiJUnDin00
DyiG1i8HIgnh242PYnNF587MVRtas5s64wzeT9YrJ93f/3rDSuNlQWiCsL8yGKs8CT6+oZ2LmGA5
BJxngPLXd8J8MHqGwNfiv7XflyrJBkqXIccLcZljZngF851zm6wwXGj2lcf8UZj9f5bgau7Emxsu
yxnuJHtW/WzRHNhCCoKvM8DERzpU17sPZOQh4qJhrRNfDD2wD5F1fYjQ/6iU/0AKQqBAkWhT9JOe
7lTEw9fudkg8i0iiuerFk2KvL51tAw6NlVVllRVjwXyi1/jxzc/2VmgXtx0ObNLqde2pdEf7KLQE
BzGmJ8CI06sIFrq0U3PEN3/9SHbu7IH3xB7Oe6HA0n74N9sAwWTAEHgcDwJ8eSp+JNvedW4chYMM
9fWkuYjVQRCh/v2czcXxrev6iPQTatHc7seXrP7z74eQYkhZD1T0aMRDEQYlj/dNhX/ImH8KA08x
RQy55LqArTeTnoyrbkCs4QJ8usW4CtrI1ZmYQijqxZ5cFspNnYqY1/O1BQjWxMiFFrk+g3OZoTNs
/Z0HHs8EiDSg98PsnCz0VL+lqCYbqf9NFAomMIN/NM3REYsJ8u0ZJ9l3gdBWKlVCwidcLzXx/4wQ
Mh5OJ6ZtwcUmlUGQPV9Fucvqq/yJQ1amb2fztY6p+dPtQwjpKYV3gsyCg2oxTqgWo0+6ujieaZcD
P7QyAUD41l7er5AFDimX2konxInnx1VMX+GKP4QLlmrCJEomETBw8TAyrIcSaPzOyuS3vEJGObt9
TlHc8xoKAgZJoihQiX0KAtTZj3j68IzJevdUmheA4Zz99g9x/D4JDhNI+hsS3ixE5IWc4OmauNfS
yaaDiXuBdFW1U57/ATf4tRiS1eGEK4EQ8IyqlZkMtg1WUltXdAzturzg8f8n8l97DXzqG21msvVh
E81re+fgyPdVgXWd/v6B5uc1BK/mC0GyROCXbz3F/VKCmNuYvsu3oC7Cp+aJOqC25SmWDLGgZrHT
1MVgYumO7JxaEnEve3s+T8rB53jiqzpmPn/gDgB9KQG0Zmml9ankzog2OOzI30a7F/MKtNFOBnlp
SGgyAo2EaksnF5ADoAZl/FvGYPfmHibfwvwNU4qbQBdalE169DbVgkxPqsCVAYMZGibbbseJ8Q0W
kNZ7bCrIpIC023mZDlO3L8K2e9wIpOUC0PxdBUomt1xg/A9sbJAkz7lebQ8o/BxMYRJsN3/rJpLh
tDBOaTErqe5oroYWvC8iSDrhJxLoarVlCBYbE1QUk9J5O21mG1NhAS9sTZuzMwHFLTgvDdn7QqFu
B2e4/loq5c/M9Nj1oRr3jUhWX6qZ/V00Bg94nLZLNXT3N1cj5E67HJxA0TBFAS17es5xEDz/IU6O
IWVMFZBIUMZrWVLZO9jxH0iO426KElK2R6d0+kS2oqvooLvdJJFhxebMoSipqhuEWxvezR4xT30Y
JftgZ3SojgGhXks4nlZx1bIOkMbKUURBVnMtQlTh/MPeQPm8m+Xmr241uPFbQKYLR3h68tE+NlIp
Wr8+74C+hc63k3M9u79eWhBTz+EbUu+S2wnViXyqmGz07QAFj4wz8uQqCOaG/6sSzu+KqqP+95+g
cS28nH3A4KXntLVxkqto50hReUARSx4EawHTV4OIUkrmndn5srUcnhcdCizRuE4ShoPrRenAOR77
z8Q7tiKYybFJJj7YvefbtmwKEQxryLApF+eanMO7OYELLthWGYZU03a7ihkGQ7pBXwrWjAmtQppi
OXjKDc4TJKCClwyELqNGExIC1UTUitRi4x+i390wEyVrMTnTDuuVmg+ALgxlpq6jyanx/RRn/h5f
fyikj5ScirQdldWG2X9h0KItaeQLafIFX/zXyKz5BQvYrUwSf4fCoj1sLBrPPzGwVlL9kd82yu9D
Lr3NSl9FNOfbiaptkCdcn5EcJssjYaIvUarAka6BXm0v4dBPYKgj4GFrSaxdhIvfDZTk2sOyTW4u
OLZSPVpdpAgqUr2HLOG3xBm9W2i8kHv+L3qyHloJZlbkmBcyY/vctXM6gBFpAPcp/5NeYsfy4vLy
12PaZetqK0YiYlSUwM/wIkXk8af9WGTGjvxHML1S+c7efe+6G09vCUYB0gF2dLS8TMFRQ1PxqQDZ
eMlk6y9A66x2eMj71+megdO/MKS80MHpYZJUsBQTJ62KOLIEnioOcn277I4WkUJ1ZRkkPfatDwU/
v5NCu5zpD7HyXE/dohRDE0gnX630OPT5kuEtpfzBRHcqRhaOWfMNw0AKSiuGJxqz/cjf2pOYblGb
N/x1vXnEuJ4MdMExza8EEUCGk9tbsPudam53tkBs6I+kZfefyEcNi0zj7zncub9shQCkoOub4cN5
aVEXWCKOxkWVT8W3WNv4TufBwWKokpBjRc4KFOzxepYIr3Owh9EpfLn759CLsXZObQSvw7sI095a
hivktaf0M82eBDqDQJg77R9ghNG42hlFhKjLRF/tWW83ZbgU/mL9P2EgikFWkEWVYD5OPe+Uto9i
k7fLAcBO8LfUnNXgN66GhFD5EbAUAp2L4lBvAvO8kpATLGcMfX3bQ498FGJ/eXwKAzeYTahfV+Jy
m7r/NZEZKnAwdbulDV7mR8I3PDEOGEi5c+kDwvK5bxnj8VRoFMMeCb5KbvdsJGp2j5VVhp0bDzqH
SLoeghzCRv3ZxYdtxPqPygkfGkZ/88gnq8k0MF78MAi29Bv8cqAGqOGabLjwSd/sHn9tPp8qBbwM
bosowy7LGioTgvSJza/CwVfdaX1ktVoKrdolx9tOW/CRcZdPBM0WRBqt48rnxsTvjSI1d40i0F8J
A+FfIf/T/Jbipnh85nr7XQNYrgSEUW7xMDPHFbGTp9fGKD0+N1C6cEk/uG87WWeqLtCILdWulDN+
FLKPdyJY9Me3nWNy0Uzf9mJvNr6/pVHUnwsMwNNGf5l+H3LdyPjs3rhW3bdS2cKDu4JtEikg/+L2
DIZ5BcT5N4PrdROAHvshmROa6HzxfmS8eUJ98SNbQT/OoxTjnZ77r871UKgKrGfCFagqBziIffWr
igGiU48slg/UxqatfQdaSzdi2J/hBLuokeeYy/E5rq3KGFbQ7L4mmw51rpXv6IzUcHA66rkV8Clo
1BZljhkrnGfgQSQ78VFvok6l0fCwy0VbVRVhPS6/kdoIBE7qXVXY5IQgQRs5GNodChEAAPEPUmNh
Xz5RFM/4LyPFBvU6rUcVzQFbvQVatm9D2lauVnHojwg6a0UVvf2932DhTkPQPXfi4m9LeZBoaICO
0XW8AAIGZZnlKHLlMhYs0b80OK0bPCir+DbIlZ0oEQ5v5o1wwLG3c1QoQ/JCgJkBwX0HTpifGmGv
5hdqt1LO+0iNVCWc1gH74iNaVtXBjIpomy/XTKTfXPNaFnh6NUeg2fARpth6/V6ezoIex4yBdpXB
lLtBaWFBoiDtSg2p0S04WKu9DNVL+hPIUs3pGwGE/65ZcG/Hc8fbReSDvCs2Kfn7AJ3T0BS66bt4
vj1lWpCE4G6Fdwixu3uP+27DydgSpyJpV4Bc7ehZuIwoVbNNnrgUhgtH4xmTGb5g8cQCai8uV9u3
RFNkD2Qut5HJ1gZ2/ZhECUZJ8Ix2vupucFuTwigcLiyvUr7oHVBfRTttFhSqviRwLcamIx4A1G+d
DY1AwUMXXX3wMZEt0NuMoscypdT90bwxyROYnIjTjI+/EVag+WFu+Wn//041VYkaK8OpPip//7ZC
VP+mbb6uD4Q/wlojtdLZsfHIjk8Up9XA8pWWtabGCNcniXm0Ve8Qbg6KRAzoZw5Tj6rP3W8dill5
6XhTyWu1BBEtsvsqBEBFqjBWDdFb13JR/ghBwuvLdJAJo7Aymh8CYPCjpFAkUxZUVIbCrw+jNQ0u
2ifswGQF/8otMF41DjlNNBWOfDq1ER6loTJnPVyVdBXDwVSAUmtqY42uT0Ibd/OQyqXPT7yl62W2
cGIO+pylH2AZaVp/LF8WYj6j8QRMlGU5bDVzpZI8L/TBvJmaIruX4MNj+3/glVd6cVIGpWhnvzgZ
Ds7NqGj+s9VrvHThhTZLsN8ctp1AUdZPSngbNEGiX14SRpl2ooWSIpKEiyVJGJnU1ztunvqb78O8
dxqbZz8bXuNdkZuslV4OchHtqpma8X59nEswmZP8nh1nVAMG7jxUqfQzJeKDz/1Hvw4jtcVpjkwx
wE3cpfrywYdM9XiCkkhpXf04wDAMrkRQr7Q/0jxDtDwYJWuWk8A8qTJ9L46j5Ctw2B8CgCleWTiW
UelthmoDQeC9vAL+osRHfLiVrEox+aEQyxHZlG2sL1dkvwm8suk0mqbsXIg8z3ztny5WsilkY4e/
hz8SA4MQZF/Bczjx+NVKZ3iIicvaVe917GXIv87YxH37BRVGmLEXx6EmDMRekEj5mV6RK/2MmDFa
zV8mR4jxWJro83n+5qkmgP611qiXtbvEO/O4d5gJlREl/0hJdkCDU55guIyEBdyySvrvQn7xUN3M
eEbX8yH0K4RX5FR0HEu1G32UpXG8gxk1omJmax5+0SAPTqyfBrT0FB02rTjvMWnQN5sPel0k6zYd
kZsPPMQxEsI95dsrKhBoTGdVRco0pCdosn/tMGRfVyj2ecm0bADrYMncPJtMwkYVF/nDYnmEOKEo
ekmYGJWtgiom9meNh7WSKArO9KAFThyatYEV0Tt8ESFdCzVrv9rV6ODtagAjln4pnYBA4PC60SlU
RXkwo7nJC5/wH2OuGPAMmbT1pu9f5yff4Z3HyD2cNxWo1b8vFAkjcN0lsbfV+DZ9xmwpjb/cqrEh
R+yRpy9gb5TRmtnydL0RLmzm240KYp+9mPRJATXIHkJ/eX6+z9bMULmY+KGb4JtnsBPc+MpKcoTp
YtLhn4HWKaXRarjaFXqLfl+X4iQWfg4kwYnej0qJcVj9YQafRep+PK4cK5mBggReS/Z0is9t3LHG
ioHXRYBAaqkBLMF1l3N1ayLjeEdt3DSAVHeDAXCCQdSZNtr8WqNuZXtf0ASALCDXImgjUkKwUKNa
ymimP4Q3zxa5O9OZayoqzS72E6DmXdVnwh6xv3XkNIRsOt1xe4hfiOlpQ0d6vZ9T/S2Bx+UC9zUb
Ji9kWOVoWWdf23ebnkUbLOXmzxejf24pdEat4DQsnousRNRWvSRZbAgD3DjpsgBDSpHMbSytzY2P
x76ipL9l8o76UO6+JK+HnMKs5DneQH3e99fYr7u+zts8vWxYXEhXryz0LOX9FdWizhhi43L1Nd7Q
+FgPUdbHzFmxPt71tQUfjuo9E5B3qA2pPDSPkERuWQNe9AJgKQl6Vd3GwBRMDuMTUvQHP4nhY/kO
zNdH6bAC5chwpYHNozU02MiwvGknKFlInzvyUdKxXalZZmIPfNN4HsgDEf5yj8dZvK3XSDPRr7wZ
xoTkLdpafkKUNr1uw6udbOjqtYK0TfaCY0WAlHZE6utxcAxfWzGcXrykWH6Pee3h85iMJx8M8wfK
DzN+zu8BNwO3pt6BXjmAuRpHQzLLQ2q2vLzoxsGbM4kiAGHTC+LAwXryqRFXKq9NpiemjlZTrDVE
WresBwbtffNfYWtGIS7ryjHWikFdo7wTeam97afcpJINw99i/bn8Y2QH8DP+pg+JdbtTWMMuvtEd
7P/BFWaOFsQKNFkzzMYtLM1KNC/MQLt8jDchMXZMpxVb4+uGhmW0BsVNvVsfW5Qdm+x3PREql7TY
yMFE+kbU8tTzwOFV7bi7OBIRJejtMQT+Gk+NyboAZnwZ1DUrWQvZbFxFzbStqK45iiX5klwuuMCw
yqqMxlaQoQxNgbk0icpSZcc2zOds12bkt51Ei1H22LgbWVnGobdth91LnOhX7rCXWtlzeiRs90UU
XWDbo5dX8ed7ldQG91AC92f9JH+CLJAPb8EPN+2toug6XZ9q5+/WqYFzmSaJx+emXswU4Lbm+VBP
JSq/en0+IKpKHxVSspDy7vG3HdP45yCkRIuj1ALbaBEKuSzw048ywHB8goYP6UXUg19JwJd7pwkr
hB0RrWVBTx2eaP6Z3CvPolm5Ce4ojcvYhQUpGn4mh+Vj8Uq9L7yeo2OZFDohotxAdQxY01kHusH3
ZDaqDP5nOBbGCT26czjEZwsSznMO4O/gH2T4/dxPctzBrcdEvJApIcHZdte2qLtlckSKUxJFGuvz
8jDCrPlgUyZcS6mtXXGF9r/sbUWae7V2VqM8fMkeytL/XsoIeM/JFsc8zSDOoqG/ncFsDM9LLRjy
U4WPKqzUCA3k/jXm4Fcfkp8Nf6iM4rzm8OvJwZeiLVdi7pHdh/x/e5n3i0F3CZ2cI4NanI3kuoY7
ymhqSqBK3kW7qJ7IEahQbYA/xCs3XLsTg29J+jzsuiVxYwWfOe6k3oZLvSGgJkf1kGnPK6licMfG
EYk4MbpgH+8J1mhiToduMU4t0PAKF5d6Q1Y9xXW4KHsNZXnih8wLrDRZ+25jsPuk7ceE/iFN0reU
k0uotRi8ZZQAlmQn0RdRVr/EamzRw8yhZH16ea0F+Yg62YE52DM02fhVgiiY/o66wzAjSSkW2E7+
qQvkFTYuG2e9KqgJs0gIZqEI+ntncB4SggO13BJooAQjLaOLFGDmY5EIKE9O2B+NTdB9WlkFTVZv
aGOI7Vnk63cm8UK65g7rZ0CbDn+dOzbSONLbnZsa1r1GeYrGIt384af7iIlOyRlDxBcR2wa0AsoW
AzJ+W+tVNzcKJDniyOyWe9OCBKDA+jJnFXnjUgmdw1qYoQhtTMTU2rRin91SaNf73H6HkVzCYsCN
/xfu2fkc6kev0p3nLEE227vxN5a+8NFoXcJldYvoTuRhDgYCFCgf9s+ksK0j/VI34MVJ+OQXnIJF
hkqm3V045fyqvl6x3Xk6CPiPgrhnVyvWaZ4a9e7bhlbZoG0rANygKZRuRwqIbdHT4UuUkiHO25Ve
EMZfna++blIt45MpCV9YB1b/sHiV9kGxHtuMQluw2oVoKXUD5qFZ0UHqOYQ/ZlUuA4HIi95C9On4
jtbVQLuG7Iy2gfg0c3yJhOHD0Wq1TuJikLgTwWq5c0Xn6jiZZOOyrzZHF4X2CfNUPhZ67ctP6Ol7
tNoBjGwZDxkcUSp6fzmWJRjLX1JZ7NSfjbWFv74tZHcDexmektqavunMziTfWoggHKXxRFOhCjYH
+LGKU+GqI6vnGnJI0gNjZM8cf5pszniQCAZdHLLVbWhyS5q1Y2Ocp/kh+LBQbPxmyxlDN7Tl3xc2
Jyw+I2YgrMz//wmw+VkzdxZIVyg761TXu0luFLZQ4uK6z9DN4V8q5TgwusCSGweu0YBEJ11zZ9IB
yuks0Ob0qxTh+sQ+aKG2dffJtv6BvPh45VLm79HbjJZrDmmdcVcIYTMbEv2MlHGAIlInDt1QKReR
Wn5CmX1/LyP2p+HsgMAZ7b1WUiozCJHmi51zcj2z6333dCnn4o9iZEy4/scThpZ813NeCQdndJf2
0uotfEG/2QQ1unMksrSvYG+UUtS1Nj+N0KhwmUaOoooeQj95/TuW6pNhQhvHjf7YmWQ3YbB2lJHa
9fk8Kvks3LykSStkgcRdAQGjEc8/unVZVgoitdjniM89+UmYzAmdjDBeuiQ3yPwxEXO2fP3Z6euv
rCTwfbPTKd/csw7PotKYZC4lxufg+y1ig9DygIBSHbc/sAQ6Op2AMmUtip5UolN3zmp8IltkzdO1
+8c467XcexH3Qtu4jXbg5oc6rhGbl5V7jvvsAguzdiLhsbgCgzQxGjV8wWv3nWX+Qop2LkLZYe6a
Mn1nU19KROF85c74TKlvkIaWKhsbDFYvR2G88mWu7PFki+aZLG3vlIdKFbtTleouhYAlKN+vKC3K
y+18KHqjfDpLT+Gvad72jajbIV4Ihp8MydmAjA88GI8LLFYOJuoRUhd4Dxs1npxlqDtAhofEiLIO
s5cFAYHrBRbfOWHuNSUMD0jd6CFq0+QJxPRrwQY3qVoR2qc6/qbvSL4TW0oHzORVJDFiRdBKwu55
8ZdzBpAn0cG0d202+uW/bR8JroBlqPpb3pxtrYMtyWx3PzBACES3NsWf/cC8v+1yBDP8C0dbvclw
RdD81h1+FYck5rpUNFyMp63CNtEN+Vse6aBSQdO2oNR/V3qw69bqIfv84k2Es4r4Aq5snzpcQlJm
wysX33Sf0xMVMgZ+j7q7rr9mmED7rA++ikefySzajyUZhyJJ/I445aoFmbk4psAQKIDF1wbhOcTW
7f45dC1ceopmW7NuFLwHtlsP/27kb3yInSI0n2xovR0fyrLQe1G6OxUxmHD5sC5ipbDRQuQx9apI
F95+EWhdzPMzpPrwuy++fyj/u8/YUSOMomiz51IhtMXbtf8ZfikI2rgYxqbNkmc2qDCsVU7OEGlU
2HjkReXbrN8TZCANFkIxER6seM1fRNaze/aQEPAiRN5/27//dT0iWCCfG4K7nw1Spceq4ySDtlmp
AsWWL5cB80RD4l/2BrC1VgBj6khMmCHJo8SK8YFks+XYQfTV2LOOyPIAH/cMW9UJuK6j8EwNFESt
rzQXyhS7PR64wP0DQTOBdOPs2QrheKWLbKSDE/7cs3R0472RqEwsD71LeE9Ah4L8MHzzXoRWfLvf
RpwaEcz2BISsuZykKdXpyqA84QJWLjNJUw6QQ8zEAJQWtMMpeBOO57UVInkVaVs7jPZLeq0YUuBv
SFXBiR7hpswUztiUu1qGKmFH6lwKtV6St8lQYSs9nUibULeZiLswF3oDgzCN4R7+drT7vQZbHeLx
QmPl8m4xssVQVIMk5z3nOzlWGz+vKNCpCRGUyVY9YzRECIavqFNr/YtUShPNMhM0XRKvzX6DFW3i
nF1LGOm5J67erDOlhDY67jrCnd6qz0gfg2tRdACRywTA/8uhPTKRNbDwzyYqAVMRJ5Im9zmaUs/J
3gAFOqsOhCJ2bLZT8SS1SM6moV96LYVSmZWDXznhAWW21R2pGj3XhtgJcdYudOrV6QVGFkRjhlb1
6Rdz6GlCXDLewHiiHTTUrPkOtoLoHRfoab7al8SLIQ77MWjNEpwyOFe4a5mnW8c/Zo9iiwwRm/hb
0viAtaCTK6WtX26IXjEaNxJaGmgx7eWDwhJhTscA9hcJm6fqEJPlhHI6avsxeHl5GLTMuU49nWkb
ULxN4x70UKRWYIdPBaKLWu9Xb/DBbbQA7Ckf2/3IUnO3wyKVikuJI1EcMFmk1fawSCt83AidtVo9
gwccZNf69O3xQU97zTMqED5HlCUD/PRGPFjkoRqAEk4TArDbmZc+aXrpRNs/CM7Fx/r30lR8Hl7L
fDBpZA43Z/ghxlPeG5muABQIkVoN95Wn3Poq7N9HF0vKTieWKUFvfAodt4VIgnhmduajtI0Fdhoz
TbxJ6w8VbmjsCmUIc9fVxtXzviRrBzRo0NflouQlMkoHm9DPHQHDflX3G4iRdSJnWQincigtObrI
jnQDn8+7w0HMFba2CXwP54Ahwhj7XzjZrOP5UsuBt2TuKJqKAPI404yf1/oNJdbuES1649/dVlvh
qmP2+lc4rsv5Qt7Fg3AA4TkS/xagXfKy5xeRIkDZksBBm8ItE9k6/Q4yRvvwwliRjhH77w13FUtN
7x0KHimWYHfdMHGCif9baKvhnTN5EQQJXRytewut1VlVfhXZ0Gyq6LOWn9hOe9Lxku0UNYj2j/3N
x44WUqMGXwZuUS/MaLUoEaz3eHUbPX4aCjmsMjrk72h4isUrS2mYC197pq+vfDg/q4ywffdJUm9D
sfLI23c2tvF+tgbvK1log+Q0OiRHlrgFSpIoXCKxzvZ+Ibq29LesDn57h9B9nHpEzoW/nV6oSOid
g+FPLbhUqGdEjkVpWAiuOguUbTBYy5QM9hEeN+Ed0A3qr2XYijACICOD6KJo1bqXylHJn3wq/lK5
ndfEOLD8C24Oh7pqDVvS/IrALKVQ2+sfUAJaxxoH0qlMYYGbZRWkNFw8ggVVbGVZnLgq0OzrLcj9
Nlr6Tt3krflkx7VI/+za0XgU8kJ77lXRUMdFvUwtLsk+DAyhOigsFEsuS4V/kDPAbXQReOp0aom/
Vffti1FqeGs6qwS9NKfO14AbAqODYbaulNyc83j7TketHQwk9rKNJgY8UdWGVluJPnMfTUAeF6LU
OgM3DSaM1FPU4fS5dcC8UtMdWkrUaLfbxjHeS59zC0q/pyAILIOo3RrhlNOZax83xqFB895/XmOB
s9XP1jbkn8HtgqFY6U5BmNRexS1hgIy3H4iuPrlXlHq1q400jurlm0x+ucuXaxlETmwSpv4PuYwk
GANXUkH34x2DkT4IxVfIgtkw5glvwLu5YIZGEXRD6Sh9MLXYsPodDBZk4vLxO4Pl77LXl7nQb7Zq
6DyTfX0BT8LkSWo/yXnAf2hxfkXmjzfrk0hstaM5UvsuLcM1bUEyY7Xdm0RbYCcY6LTDiYcGP695
42AygSr2mgKHTQli8AmSoTKBAcGYQbc6E0f83Ml0XwBsLIOygbH3BzRESdoiMosF9gFcRkBpeGzJ
/6MgP8K0ZBonA5DIsI4cwagcUszzE7oDBx2FpimvaS7jcl7GcGZoxtVmKR1wt3c7JMZx4WlClRdX
J4kZ+SJQDqQ3+P4c/GeaNgc2qiaNktJxYoWoKAhf94ysoKlCJRrVUYipreXA2t9i5dkcQ/4fZ4Qo
+uWn9morZaxlTfA6qY7x1RnFhZTyWAolRKJZCzxiGknIox25bqIMekHGii8hInXl2GviYrGMF8B/
0JtJ5ADuMTjL8ajkVn7V38SwC8ruOqdtAU/HO5RDcRJbZAk1WUJg9tXJc1nihw5X18sUThC69Avg
RcrMbxMShd4zRi3A808Y0x86dXdR7kApmoNXIN9uiSQxi56cvBiUnzDAWbqlgO4DIBfh+FbClWWA
SZTggqBs+x7TtCbnC2+wQd+6+AY3zD4fkjIB6LmLEIwD0HmiFLulFNJv5cfBotNVRt4tgUPsEhLQ
ilY5zTE9dGy+hAI58Xs8ku4LWe//OaJ5P7ggsbnesMFmauy/XCWxsk7BgNNm1MFevjUjp8vVFPMf
9r/tNb0hDO6k+NsxbHgjTmX3YMAbWSoyxNK4AfA7SFpLQwvVaca4V7efAfMDvkmZDYTJLcr+Ugrc
NFeIuO7+qcB74FUdCTpGT82VUVSkSVY/RoXodLXgAruSoV3P0Y39cESvXsGfOf0O317W9gUANLFB
UHfgXuXAnzVEBAorQP+m9gTQCRMQCfJsIavfgaSTzG8wzkmvZmByX5Gk1NusRwt+JjgVSK0760Ny
BQ+FcdZt0R7yhOEbb8knvrvKQk4UV1KnEFb7n4BPGoz4ku6AMc4cG0zGlPwjue8ydleyZgAKjwC+
SwBJPiJ4Y85P2L6t3eIOnakVEv8nreBRtA1kIk8k4aljbdugjrvD89Mb2irg7Hj2rMSEa4nS4d1/
MyMtvtfwXQNHwjfYXJW4aebzcnkoaiTmOTXTdaYSPDNjwADmf6fK83VIbk2RbVgH4TDbVexBQJwN
Hh1kOJJaecML2G0fNDHTntU6JvKsk5ygT75h9wv34kLv0/g+PbQoaxaOtb+zxl1bizpNV4H+evE4
vxw/bqLNm0DJ2Pw3BM6syUVBhTNP7N8dVIXr4ZZ+ipsOmfOy/1Axe1sg0Dh398Otp1H1acBIcbcK
/UqLbaW8PcS2r5xRDI+Uv+Eqf33MzpbYijHrxmIKoyED3T/h+SUCzLM/tUjZPO1g3A0GtQ13hYVQ
K/CJJW/V4+E6kNoWWpGYDiC0EZP25ERAjjiwKqMlOYjiPxX7TINHinC4gl/DxFe5/6QJlrIjWSRY
zLMwjsSumODDGUKr8mzlWccLP0dcAGpW5yjmHqXQBEoyGR0xJ/I1nGaoEIyy7XZN522+FjsMUU9N
1BoegNKIj1LOmeLdJx3P7XaaGBx8d2MMVqqwUTsF5E+0ccLRAlriw+mUDn5QKaVtmzgbmKWlEuqR
WSbMy0i54vR52yuFmh4rdcxRi7HSApR4Zdh+uF7Scykz7YcaDV4ZqRxO3YaCG7bWfuJtRyl41gPN
D1wTN4tRPeL3AdBTXi6DQDA7ttgLdC61BzbKVkyeY8Yk3z5L9REBgLJxkg3JlLROUivZ49t39DRF
xni7pUCt658TyNeLOC36MovcwZtwKl9U4uWZ8mLfuSMCTfWDdh7u3uV0CkmgcUilkfxGvvE6pEy0
dgWz4SCCSa5vr0I1tsjhWwQWA+KqmiuFff0GAEuV/qSUfgzYf1cXq0wPe1+oB8ZV667wU4/4Y5Fh
++mba8Sf9WssMpiwfKtXVA0uSs5U/cenT08Oe4ttKQzuRGw0dQ4V3GahRsoy7v8TB9w7ISqbAwA9
mtzTcKFpERcrMsHYLTd5tPWsOo2zMizWlQOot5aJliBZVFsAnQwMjK7ATHAbsoE5ug9XBZvWQPks
6xfLEzwvNyMxCRuD1pDw1SWNFEJWUct0/bC5lUxErzfGpa1Qz9dT2NDBJSEYiF1JwlqBdJIv3xcr
1ynZhAmZIJeEbzHfdaI9VHIs1lMnz3Hh2Rn5ty6uyETx+CSnNGUaN4aP++AuM8MWmVbVzIrIX54h
NjSFKFZ1M19RISWuDK09ZcPlc3AOptl+OaZSWWJQv9JrxFFetEphSTR+gX54h1N6czU/Lm0iWWT6
i3x5/KJsBtxlgg70DgZsF1dubE6p7145RxcF7MSjqUe/qoQAb94y1Uc52CsDZb89Rnyco0qNpTP4
xAsGN+Rbsx4BRgemP1zUskzWZULQrGfBqo4EQ/m2tQJFmizB9LCowrNhLXv9Z3G9XWpRrcJlYSuD
t0/RmU1pPyCrLzDeITVsZxO/FiQjW1PlDxSxhDWeuAjCOcN7pq2gVp4GQeV5uoqccJr8p/CQFZDe
v29ydDL7I6s7THPl3kUh89EKF/gMET1tWgOZRuU8xvMcOwhAE6kLNCEzuVWW81F/NWt0b0l6SSLM
lEKRiQsddyP1C01/CnkksPpR1KVEapCRs9KCgDviqINMQO9WD9fvypsvJEVOLVRlJzR0F4QxAx/V
Wf/3Ge/JxaooISVhl1F5CwgFG4rNNBM9/g3txWvJAGW2yWfRnoieqlFrxogUcAwNJ+dcGHovU9gC
3P3Tf/bvFsvr+i3WDyDQmVNGaM78qdsglzD3RGjmkUyUzvMT6UqTiJktTqxK97CZgVYlfXO50KRI
uyrH16i4BAXQt7ItSW73sNQF1Ac8v09tYnDI5xunV5O+2Cn/VDHxYxmejhrfxOet7vkhQmdM+ing
vaPXukEq/dM47KdJbIdPhuZ8GBt5IWFqho5E1PSsVKpdsKcqWCI7ec3DZtukGNv0T35DHQW7QTfC
xtE2apxRDMMC6kSFUUHRkipKjnEz537pTnnRInhC3ZlZ78Gy3pe5EXCFzM6gNEL4u8AUfDFhNdGQ
Y4DLR3legqF9/g/MuSRUF7VAKZVgJDwd3/aHp1b8bFF7tI0oq0pvwNnZGZM0kXdow5R9Km5U8XAG
wLPok2kc2s5GugZ6xaJ+KxRYeD9Q2oN8cKfWyKiiILs6yAS96wHj3Ebr9VkjAOrnqHQ3J/bizv02
oYoTil7eDzwxMpK1tKttY5wgyOawZsW7MaVRf026Xgh/uWIk35VOYPRRnu/vZH3F0pRvSGybEB78
pcW6X7aAHOfon3XYlUldJnch9rvhGA94cqktCRc9Fk7PR85SMKj9+MBSstLMWCrAmQ1KVNTe7EQ3
ziJOWN+DzOz/8xDQKGQBsrkhy4M7ymlMrr0Z+lQL81CIknV2IZkQ6uUXNi71Mi6jTiiEVQ6vynJ2
OG/pU9kIidCP2/qNxvlJzIC60HSVKeVopOpJixd9Plp8JCr8coknkwt9azzz/XFt6g/vggLo9rRa
MuGNpMtDHjBUqaDEe2MTYmIXR4Kq599yq2k9+88TkOSvV4uc3/GxjkcywbuUiXhn/d1J9Ltr6KgL
97RAphq8Z+Wv1dj1iUJVOjZfZ+BrQqiWC1DlW3jPwOz8PnfSWDHal+aI6voGy4xHt0EGncGcCFXz
OzLdXZauW0IjlAPevzxHu/27Y5TSlomzQWY1Bi13UpQnT6CBP8ujgNWRzgdkUpxYAbhqkL75TU95
9JZrdoLYBgjTh2GFo79q7ioNknGI1BMj3xnrqZPtIZlhAlCoLMSJWTDhERl92lbcGa4Gz0kN0X/5
nc3J3GoaFn3eqYpF23SuP2PksEhG8sMQzcTuqIiDIHkaWrhNojZBu5tRJYyC7xTdOVBxKsE49NEh
mnAv6mRc5nUU7N+lXN1Xs4Me08JJitSUT0Tl6NmUolYVejqnxcIJiVVmc+YaRMlwyKxRU9DnZVcb
kVrL7Pjv934u2A0SZwvKJ+GfmSM7Nfx/HYoX10iZYgJ1nwKzpyHg8CszvQAngjprZKMfZgGZZR2Z
xWZGHvtCOskYxx5btS6U+Ogyy22k3pNHFzEon2ttmututn/o96rrLaNmGEG5ioHDFLWMxoB1kIRn
3KIdgRklhwFYYIDkE6uDkpBqpndPxwbkEGvQmXOYuYuFq6Xe22yPUs939/RowXAFW4FteLLAiyni
YK/wqaYf/tCv9+nhYFO7eEIGNRmqjY9SHJsshVkRQgRlz+rQwVtNZV0tCBp9TfUEbRzQ6E4kLWUp
sS+ddWVOmcXNDp+JnTxd3pvq9ymJkliuBMMjXlHeQcjbLbhKOPC1JEMBbvrRn7qLEzU3AIFXzMuT
fVwouDDeJ31KTv2DDv8QaFJP2F8NdxOieqDD7GvEiHBLdiAi2kIQmYGY/QFh03rC7lfkSabpWLX4
XcsJhOEdX792Z+mnQ3ChR6WogCTVRO91cHCVkfofG2QGKiIYGknEfXmE+DTbtCyisHG0FW0gMWm+
6s6Txo8su0oOnk6B+IBglzwfKcSlKXECEAUCddr3QV0bsv9x9sz83f7dWUbFzEuSR7ej+nHvpAWi
bCxZYsqtWgl8Q2kiXvlRTNQb8m1InWXv0gEofZctCG64swr7tsr+SoJ/dJ8L0hdRiAxpqzLtfgi2
ftO4bVFt5o1a/zKY1PLomY9LHu2MNridxRVv+Dqe8VscMAH9J0HD3H/bwVdVl3MiRJH4qDL8mEqH
mb4IdlYMbuhY9yWrqK7geQwkRVgbRHI1dt3mJcvl5SJMkGrcaxY9L0iq0ziT7cBR7tSpztcfy+Q7
6CacRZVwcbt5OfWkVxkqJk7daMQP5hbF1TCyDictVdfwIHJmo4b8tED+vHaNJpy2VqDiwOCWIgr1
DvxyJTn1ick7sGytgrb/ZB4Xp5FWoCi2hT94HxZOOrqxlq/29AXDJT/9JwgvkFYfXwTpOGBRj8RY
2sLUDRjENFxY/ZY/Qxm+DlgjzlnAeXTjQJOc3RVu38NA+JtlGfA2XiBl+bUoESrHemdmlDajAKjd
oRC9gUGLUwkB8US8xXxTCXdU5XGYK/GZlj2PoJRtGCKscSePtDG24clH+NWfH7Zgvv/lIbx2MuN1
JfG5cyvrqobG1qdATeeGFHTyInmNIWwBFmFiJ8wfKGnL1NV8cSm4x/8A44JTp9pYCBSgLgpKZSYW
XFitkW2Hzpz6WHMUKD0qjvMg6PwSB+4oMPv9MIkkQbDbqJfN2sri+/z/ClGblPz7L9TvpDqb/QiW
yNLKJiJYXJqDf6zFjZN243SEhGsMcx+YM4D/ikx8B45nV86Uajqsg06h4ONX39gXBz0c6uEjLBsX
BeBw9+9lYrlMKZ6j3lHVQC04zqoKcyP90LE80yUnVrURLCjULsdHAovpGQxoYIUt0NiCfM4NKbpM
JWp1qsIBGDtuBib/RmLYFE8/Uub0HwkPSFHmLy1tRFmcQzaeU9Irxl8WYqxUsObMiyp4Fevm5YRS
bUk1HjUvbnuPvKSfXQAeCEza8nQGeBqUNV5cpXm3v1DcSCuMldaQhpHvZWgFosuRd6653Cn+fzAh
b3uNooAEeYjG96jqElbvZtofc3YvZeq9ZEhn2pP3kaTLMlxnA20FBW3J79L1EAno3YlWAd8NorQU
y4u7JFnewUh4xsYzKIurTaxbr5rqKmj1pLY9x/Y2yAdnHkAHiZFWPqwb2j8I97O5NnVHkB0KPBSS
Q/uDfxZAlTzPcrl8m03BoGuoNwZdDktyM4Ntma9VhNaUIsdl21Ry+HLcjXjVyAKy3de06nZddHH4
zUbha6gW5UH7Bqd7RGBlnL2QjpBvP5D7yK9vZl+/TtOt88QcADXEQkyErxB0AAyTjWOEIKuctsuJ
C3iGFIYskyfe0LzIPxq7lvl09z6d0teUwY/7gMsuQBQGkoQNqiAl9jd1gpN/f9RzPWJqkvYuf0wL
3q/hR/yvTHzMyDehIGOlpQbrbly40uYstHh0GhdS72diI7ov/dmu/IV82hnd3w1nQ62zw1hqFkaM
QeXlZapdlE/wyr0EdiHFvkWvAdMR/IkH/gqd9ZSIJmVrmzbivNaBro1VjeMgIvY+bPoujz0raEhR
p+KscdJzFXYoUOCY01rgFDYQtkWQw0p7vgI2P/nfd9GDD4YItLfgT5iy6NJY23Bf8Z7IGRJAOfwb
cE8vXmik8hRxbHbDHsSZl4usFUWy4JnVtg0iAdGTakA02RnRFyFWhI6rHIU+p+J5l0smJ9bFFujv
IrW/N0qU/ro3vNo5vD01059CF7iin8+JHoALqXcyFF9guiI9Norbiezt/ehC/lDiRoOqIMeemdFK
ebgBDHYdBaUW4A8yY62KK/A56WAZX7R1R0ft0bmv87NJbGMtcg5Ku64C4d4eiEJyzlwexkQuN+Cv
s3lJ80DJguAAU3hQ3qKI2VvBtcmzgmhQe+dDnZ4lSXIu1vF37y9zdPkKgtjMafUQzfC8VXC6tbD3
LfMcLluZsLBKSRGjkL7vmbjCfxCxtwRkuoxX2yTPSLuwPDkePsjg02Joz8RVciXYk4TMbWnkOC2b
LN06thV0tztwWHEhYfjvWGPvlszI+r7xKJG7jprFaYwnLpHK7UoMX+WJbIz+U/hGKGlJkZcTe0Nl
0Aca0gxt6Sy5Mge9xjVTHHYNMpb1ZERAh0CDyV82ZpS/ZO9i3amdDamLyYGW+s5uyVPG4i4NvFM4
g5of0r8lj8ruEYjPa4hU/EDXt2EZZ4jVxD+rO8Ksis4RrVLXeA15hv2iP8Qz17MoPnBF8N2kPrAS
mQDDrb/CZqUb2BmK6H9aABQHaoLcGx5gka4liWxhJf7zx2g+ggPPATFCPLJDm6ruCJ9fdZH9y0BX
5U54mB9FlEyW+aqm4b11mK2f4ojewXuoZsveUK1XEYOW+ceklBwaGKhQCoFlw6Raxg5CpiqkAjWS
moppg/NUlJsOmZQyh+0xjljdlxWvZ68Rg5e+zEGNRhzopDlXbeeOQqISsLJKxLa3uX+/1ho59ylD
xwdxxuh4C1Avj8IK1jSt3Yfn2RerviO7YvycRkf3MAPd9v93fgHXfNbeoGaM2W6IdCEDB5Zd8v/J
U6cOCN3IeemsskLS8djRDVcv1cGoIBpKFXbORB3JqM5ug7Oab0FNjta9CBQsmbSxcIfSCKwwTsP5
3wTkd8nqctImeuLd/kOpYl31EJHI2+PVmdyHLI69dW7oscJFuwVAEAg+xZjPnQ25c9NDa0DkpEp/
ELYsajfdF5AHLa7XxJ9etfEcxTeIts1l/HaEaWtKRcAP6Mh58BP8oFuFlFchleASpxHF8XTEaUxu
bDcfytxxX/5wugc9fIaeDLB5NrQ/AuIizToFWKV5rQBeF0TMZuax2LT/VWCvEfomFOAN6eoZV8ZD
BhWZLzhZ2ZSeWFIvnHgicCMjOC2bJYga8dKA5IEN+MtnFcP5o7L6Rid4MIAntXnofrC70w3jx8vu
2b1ItdZt4zlSnQh82KpESj4TCYnhRgX0ixj/S9FF6mVK0LzNjNXY0jcWsy6p9Df7b8RG76SBcGhO
W+x5sa23VvWobgH4kuPZK0ya6XhJTMca/cQocBhrhShd6rv/INx9h0i4StdfYehMNUKakyPWgYlA
efWr7CGtO0fj9YEsO9sP8fAVRN5wvJ9T6HENk89+uEGqlKT15R0jSgPFSTPwUveqm3doVFPeU6TI
XrJ6xpObi28CCnnDob3v4L64l4jj57ePCHhemSaO5phYjnt0gjWFARks7ofMby5zVljigdyicQ/N
FaqsrIPXDx/JIrGf39H8vxifzbz857MoWJsaJ7/hUk38BYiDDVWvkLb7bxAYB3CQeClNEQdiMNq2
91mhyrV09K3WYGsrRTDrWcZZJe9/QI4XwZQyVekIThO2ACAxplwn3Oim5N9a8pFEwnATWTteOAc9
GTppTR+/FjprhAHcbwQmB3GeL/IF5dUkM/YbD/q1nWQqrfWyM8IvmesTIJ6nfqvixF2TZmQnlDw4
h6fjW/oZRvmJcSOjDWnF0VJru9i7Hsn77hbEjjJFYXDE0nduC6d6MuglLK1aKAlQ9tg6YSSdLmqt
e8DNO/cJH7ZxPoAz2rQ/KDMThH7w+duqzjBU+zvvDdnkXEuePOP11wfRC19nnnFct5ZM4pKgLnSh
KvRYNHOPNWl4E7KEUXzCcLUto8eqhvatJWYRsu4KKoRyaXLrhe2HhPoWLLXtOr1Ai1ZhPVh1OsnF
z6BA4YR0ZQt6MvSXV3xas0LHeJD3IzMi3fpA1fxYPsCTLYvAvNa2kHjS71jcDuFt6PxU+r2nF2hX
re3DNrYuXnMjf1QOVgdIYFG7iNYrC6AUZz/k27xSDXDUaDOHrSrEdiFBaOXoktgKD0ELN/U8xVGY
MyES6bPIHVgyIheDr4KIVzOTnJduLIyjpd9eTQzrGW4rDhd3V3vaxZnka36vnQvsJ7EcNQjX52R/
dUG4iYzt8vn4mspwSL/PFEK5Uow/RYFD2nHOpKdyYhYIi4c0e4gbb+xqDkIAZVjuHOy32WsU1jBm
jTrctucNAle0KVFrEX2FyHLrWfnuQ2ipfGZJ9+C7AhBsLzbl6Fsf8OLXdj4X35jfYiUiG6ZVIHYC
Wh6FsZusDeMtdGgWxTT1I4aD7VPMmhlcFJBKh9pG9eZf4Bf82YQGnE4SzkPJ81IkAwbqqyNwaElX
3toJ/ge4I8keJiI5QDPTeBFcerSj88Vi492MMaDujGLUt9X0n7bPLh/KoE5klwsyePjOmxQR3QcE
4m85BtR5Eu8iUolsnz9gEYTcMA8AqSpQwUec8vb0C6pJ5QCXSeaP0zAHanjGSIg5yiSM1oeCTBzJ
coguSUhF3ep8oMhs9rPRD0TXsRtG0UH3T3m4UO7RHw8nUc2frISazuBsUOC9sZOWy+zNpEhY8IVn
Jh5amWQKU6HhfMERf4nj/s/vwYxXSQ7uDurf4sswnHn4DcixbpvYCJMwQw1HHx7ooQQL5fI3QssP
IAEVfTHSEbJFHuiPGHevTnCtqYoeYwOmd7L/pavci9T74FKckYNhHr7xnd8WUk6ZKhl5DvMPUe1f
51iaXRio1Mn+EV37tp1QprF3xhoLBlX9v4nib+G7/59205YRLAYghtVS9TX89dmBHYQ8taS4zAu8
Y4vxmpvGLXpQDQOhISpNnZeSVQn0eaBnYn8Cxxh5Rc8B55zSMkotu3qxtzHxq0pcKf1NubKW0XwX
c5yRvJNUKI5YvrIqja7t4Lcs8XCJNqSYTR2U6GNe/CdfzcpaOm5I7H48+SrV41nr2k8+pDtxcmcN
7hO0fHdtMEERuyK5l71f6XRtrDzqf1hqCpL50AvHaOJEZQnC2Gf3hW74/wLWYp4ZZ5uFYb74/Nmy
WyNYagXu/jCb46b21mYIWLXFs9mcqDBaHg33PFEg2b7bMG30yKDz3HrxNg47RdSsfqG4e5ZQv7mG
ugwP4Vf50aXpSzXcH1wXGIqk0HAVwQI32+qxqSKs+dEuRWrfBpChIMibTPgnEVGHBqlbC2rtKJhX
C/gGdGqb0S0/dlkLiUO99o/1+qAUhMEPGyqOYCNoyqTQVGhK++o+JJ6gDx7I0vqAEd0/g1rsFMin
ANOE+VfRtdHuBhmOZDtjmOvSAmIqQ0D2KtPiewdnEyt4XFNdwP3mpRaD3MR0zv8h9YTxMQDv3lrH
4zZNAtDnQQLTZ1SPVS/s3so91LxOgqDVaFFBpH4+okLzI9PRaWFD41AmbXielOEW+DbOge38chcO
GrwrtppmosAqgb92tLX6Xq4gb5cIIbiU84w3Xrn/08hXXw+lhXCyAesvKVMGTIVRUdjWCmoSYGOp
zBjfU7QDOHA5iebTJDXUWOsaO9Ci+HeRQX2bjDd5veX6+zOmylQoZwEdFxwyj2R/sGHYWJPU7jPT
Gn9MTJIsnK7nyKQ3phzOON6i+zfvpu0b0SDfBzD62xIBlhzCpzxbj8IZVY+eVmMZZtYCm4kk+QAa
oGeXmRTckx7y2KiMIlOkJnqBgwopM5XVHj4u7s/3kmTNDCTlTXqE4e8ivIl7+KbxqjcCrv7biIUJ
s93xfSIf0TsAdBDPg14v3E+E8zU6xc1+YRPpFM66xPctn/Jd+9gLlfuM8ngMm5mz4yq2LiAcg/Dj
kMqva27VTZmGmNOFDkY9SuoMb0foACC4E4puLu0QMVDDxTi2wX64HJ9ExaVcKjwV4QZLDLPME3c2
kHNG1hprw9uJab4KPsrbrBD466nX4skcV901jhGVpB5kqrcLr1l0QcOZajUe4C00+V/J1YlHpc3n
GW1MziXstI5HNeZlx7U4TKCzSupDNrhAD+F32MjanWLJo2W6k7j2KqntWBb1gZt4JnyvYXsE/sFa
S9TKWYVo167wdEq3Ipor51dOAkrptHxVHDQ3SCSEUJ1feYEtQCLEjft9cOr9Kuf7EzbeVHSCfj0q
0CIXQgOfkjflr9yown2ripjtO7HsPVm5xZ39cgVYTw2jmBaTAtLpKNLnR/apCIFvwQsefVqzULaB
NKA5i94tnGPRbOASJX1JD7JZkPVDqTpUacQS+E7KyCxvQCU4GpO2w22KbP9/4qiyY7KYp3ZXXDBF
O9vmnuBZw2oIKLsT9gaW9MC29YG9wXrPuxg0ns3/XkojTpDdyfT7HyPkxX/8SFhyodNSWOQuCioG
AaTq+dQveft66sQogqmTQLm0BS9dZ8J2AgZggs8j4eBN06busS6soL1RMUgum67hFPfWzUqLv5xn
+FR2C8eBHRQaMZmhgxINhb97+NZuWxHGNdo6U0AaJ1PVo3KJ+Rk2Hud0+hQIVMAuyvLne3fyh6Is
faPr//QiE/lQkPnLBOIdsXGZHaATl7NYqihShyJKRv4pCV3CinIRrrWI/YaWqeMM270pcWfph2AC
TaRuk8L0UBvFvtjdkCfhL/euxtErH/OW3G5kx0z1oU0epF1V5l17K+1Bl2Voo7beYHwB6Zzhcb9y
2XIkSyrYiw/HwVe+WWRQVvN1IG0SIXIFbHkAaw2zWgPUPBWxPeDk+39CGibZNnY8DDDKOa/mBsYN
iTXDpv9AvS12d0rpeqKqPzuXFRMoSE+YSYr2L42Ud4O+8ZGnkiCs1KiXwEhNLEdRZoyaITp7C9Je
hvuzXm6jw/9ghFNSpgn3oVZYxIbeZGWzAAhTqlBvVuLaKUBNQP/X6BWt8TbSQsJNkcC+s+Retn/6
YX5PqeJf9629qpDWm9emsEANXwPYygh/8cUvr77T62uAUmwsLXoBJ1smXzIXwD1ht3KJByknPVRQ
tzoz6IJz/hkk7K1YQAfcjoZUT7dHtNqJyYVGMuz4cMSgvufidp8m3FINfqOdjSR/b8rMuet0Rje3
UGTtJ8XBKLCOz91oVA8mLfu4yB28hQrzbZfQSiFPXznJqEotHz1Pqj+AYEXKPJg4xqSoiLiLnfqi
bonht5yf26p8CIwbeEUyIYvZigtMM/Rx3miBcoUxk7O8eJYjVajp6MM8odaE8SVL0HTvA9kQNntO
mq7ytbV8mjAiVu7yQMBbqms8UpyGlI3wr69+BfWiFW6YpeCvZRc3c7n6YVXZ9O++yVHGf/EzcAWO
BgM8nUFbGdaIIEpCONlvH58yKEzNaURE6nTA6DQCAORiSJkogGZdAlaCpvSvA0jbUa+5v0i2o/X9
lg6iTcSFdlfSSivhIFE5islu6zHKRP/WP22dMlpNNIzhb4ebEYp6DPmPgeN/PiSCQg2K5D++393/
vpRkZ08lrkQE31VBq2TsDX4ZCSiz87nT3Ne1r/cwEUzi1WE7Shh4kuuqRZ3+4Vw4glfsvDVmrNMC
VhuNwQZtLNXU/bwhj1NLWFKDbhUOuqEMHnGIa6dZ14BjePm4FMf8US5YlhIpg78AHDE7GR2w4MEy
ym5gDkBmiP/Vv84GTfGxKEEAH3unRdjCDxqN27cmyf7cU4NLF7+CX/WkaYD+JiaPZWsMMi/MZt+9
9hGF817anSHsuc2gZmjiHTY/5zD8t/Cm6cbXh0WayU1MbK1pjF9n5ULlyhzfM3qc4jwL2rdwf7Lf
5+4lh5XJ2mpBHNd/tUVGpe2wWaenRzFAJM88JrO++laMyu/nKKrhdVJZFoPfVudNNWvx/CphDTna
L4ruOL44pLKUqAxc4ETfVIBW9UYS2sHd27TdBx2Lsqg3piLvpXmvXGubyx3Kgy5JdJqsbO8Y2Y2Z
eboAZZeuLKmnyoTFIyi/wiqhYRCj8d44dLxF2pL+SLumqZz/aGbr0mtsYy/obFVK2/SbmSnPPY6b
floVqNveSxnECUFwwZrNtrP6G8/TjdbDHJA2931uqUUU+1JUpgN4tPbc6ytFlaOLgvGwJC4aqbkS
lp867le4CuV3VMDF7CvrdWIarFAD0XXB/AKcFdKhxt+pcQLms4lj1Gl8fVk9XfkRHi2kVCJ0Ob5w
6JbxZySLPfl57nDq6wVTQROL9LaPgvpRG11nyN4SFA6r+yZVqMzFX6j2vYFZi7XlboKfi5zb65Ab
zBRhgiBYCDw67wq37jfDOctBOM3d+V7XNRwY9TDLeep2UDZdpSP5cYAoSzxWxe4K94q/eQHP4SAb
DmNoD94KUkpDr+Pe3IjilQim8JHMYP3KjjQh+o+W7sDOWDLIbER3m+vxt2p/dKs//fUq7+V5mExQ
lM/Z/4ATeMEHCynSvEgDJrGp+l3O8gQcSfIZ+NWSkEha499VIvflKBa4QvxawamMfb5duVjhV8Qj
T+4SLk18Q12sxJG8XVnhD1nZmDg9DtWKvW2fw0qBp7otI8q1K2mKbesWRvZtVb59jHLiflq7yz9o
8r71eTcdj9oHYbv08N4LPzkcBm9RInjU7l9EJG7GDeuDyPOmCmhfDTSaQafPtrs/zQ5zR6qef2z2
Na9sYTPV/NMdEdkobeVAS3R/jBou9V5MprE6WCbNVY+CQu4ow0rs7e43X0Y8iSAfwoPtkvYNW8W1
0mugsdE/RVutDOmk8/OUL2fDcKWx2qYGFzSJW7ei2U9Nu/Ve4wDpSD36LJRVdCV481Lke61FQbdw
oAyc06bhcEUxM8LSmU9qBAYI7zSWYvGoAI0ltBNRibWSXhmxCWdMrXKZEBsoRBHDqgtW72/h2ou2
0rtWVc5/bYzpbH61D5aeAN0JCJAH4HBNeq1UU+u7nZ/0iVyTCA9w/aXELQ18oiyJ+Ws6ZjKPgSpb
rx4L0S8L2eZVuk5O085uRTQZz8YSxI4A+g1hzBGBfRfCW9LhbPYE5g/tgLKl8l0bENT/hF7XA0qs
sDhIiJqVmveMh6LBz54VFTnzSS/0B7YNyT3AimGdqHfroUYLr8rOVCG5P0wCZKADCJYjFxyZ8R08
FT8WAeV3TeI1xNAvl/xsVWTFCOLIYLL6zGMirpcIjhp2SKGwCYT67caX/ro/yolHM6+ZkeWGmZSu
Gi/4pmmFez47j0+4uhtNcGca+dUqpZWtNCPcczDL9r2e88xKaTJz6+dzvSNtjT90el0tJ9/4Qf6X
TSxqO8FDiepvq0/fSBkGdK0QD5QrRUNir9aIHdC+pEAMkPuT+QcbwtsA0WyMZalWl7P7uX/b1P1A
ZJayJFDL35aB4Y1lZZrcxPhrQRqfM+MwGpvIvOWq9wXjSuvOPOL8FK+b3VDK47ha2SvBuB4FJy8L
QYVmBkEXrYxXxjcXWvy249orT3Sff1z3xf8qHFf1+DO2hhfm80Anwc7om5oqsp3HZ2wKZOUKH0xV
gGZF17GtOnXdA2U4GRqBIkvGGFYe0ZdPD2ZEbG3Hx0D0EVTfLoUvopJ62kkKq+u6iW3pJ8OOKt/3
AVNSbvY98Nn0fGjdW3ryif5fhoI7ArGo/sxZCxy3ZrCllF7D9fMmWdY2ORsrCx8aavLxRz8reJkY
7tuG8FZvrvzV+rxwXhXbo6k0PLzDB7Whcoq/bBXf8Hjvf/OPwAdkJDdQaWC4LeK/LMX3J6+2oyG6
m7PlZqjtifnSGQyJBwrbUGPINrHywN8top5UyV1t74SHqWx3nD1tYx18CkVgAoC0jX2bGUjKhKUo
9nIKcLepHwz08qDFtytxuI0D+z6tuG7agxq9kpjw+oG1TW0ADU0iebm0jF5weMuxKWMLtC29aZFc
YHzZ5ACHnC7NVSD7kx3PNpftfNUz96zhXcs4JaOM6fqVMVrWB1XoAgqHbMamjcPKW4lzE9kWaMNs
SemLTh0J0gDFZNYkQZElqTMRP2ADPXyXXeXMxl96XnJXrWL68QV98Uy7Tkfr+Jt4HADsNFQW/E0V
iLKDpH6Y+E1YeNxabpnyfhdiNaxOHbg6JGzb2bKDtj820PDfw9ctH7w2F7rLQoeUiIZWL5240Lvb
G7OO+SKxmsNYFV+KSVame8POYbWGZKM5aOOqQTzaIIzABLwRJphCffoIWYVWkiREl960YA85mTsL
U45KcDLlFpnukJbtGG5cx71bCct50omVPyzMqDDl02vpUb2/CAwwRx8oEyUI1m3ASuBaQXaHwPe/
bBKynShalcHPPsapgv24quxpXcLzImztR+t6k4eDcS7UJOilTFCe7BA9Zf5S1Ln123fjKb70EsFR
a84ThWwCseQ14J5oB9t0yumJck/ZPXzuisbKicom4Z9a0Yd6A/GDrXzwUwvnH+bh8hV1OuEz0hVy
4A4Ab0PSgMz3at+eKkAoa4XmC0P6jkARd8Zqb9yElrKhlIXV5hvMvNJ6WH2ZNMB5POS/Ud6bOxE/
lQdftQJJXlkKwoDuLgzf8PBeNSv/SdDrOWgodHingJREksdu1t06zdqq0cB3r7cUFI8Yqrv+etjw
VjISafPiJ3MtcDV2vZyRUkFiLjmRlYIadUXlysHgcaDLxaRsK2x/uomR/dBjkU/z3MEMdL7JVm93
s2qQeYTFZIIdthvb5W1b37b2uLmBCN05U/Wa06fZRP4IUL7JO6qb8t+21pxcw4oui1ZQkvQMLSvY
dC6dPrYQOic9Y5y3ZtiCFcuztHG7tHRT1PiQLopAanl7bOKhhWbzbJ4RmXwMMMUX0gA9BGqsGe2T
Ie0n/EobYb06WsXzr26jYC3h9QYjd1wHFk+FjjBl5CdqgyTpUagDi4MeTX3hSLh+wp1Vb1hir+5S
Kqx5JfNyEyJyoFlTaOgiE6AkNzIxoB5D1PN3ouHdy1ZxkxUx0lXEw8YEBvFJzypH8XRJooXH/QwX
A2pZyl8PXjgrLmyLHFvcUVO1aWYDvJLqiZagSmM3xk+j2uFK8zxnJvZZrjRmvJu2S2xBXarXnBZo
L1NbpYJN2OdsB1x4+fHOJUVxy/03TVt+tkLfpEdhVCrs43xb/XhNsSRlGGfPQPsZkUdv9m0uUbD3
8TN67poSyhU0x8k15HrAa8K4MZNR488rHPxQwcZoaYdlzvGRkaGhIJj/TFze64ItiEXQMkmv/yB2
xbNMknOWKX/nURAjWDcB3n+tf93wlhG3scFEf6kGZuO0bTBY23vReJrsDd8T6AFnf+D7XIIUCYsj
ojlO9SXRsknpH5XFXaG09kJ0lOOcLEFlCQwiR+UAuEqsjt97fyub9Ci0BlW8CaWHRra/FYVHf1ik
5WLFoXDufUKThjOZGCaLfkpqBTxdpslNNep9muCVROXF/ccp34f1BpfWDyccQegq7FugRcDY7WJf
hsK2qWYAAwOWsIQWilac/CboB+orO/Lyh9rXKSlMfu+l7IycmdAcGQu/QX7beB8TJx7sYAgG2iXa
jmcuBgYwuOwqt2+Ae+yjgbJ6kvkNLYWN0qkcRBKqX2oDFfchCFdQeFbxahzvLU0KOxN5lMWX4dqM
2TQJtl60XVljYknuEd7dSI80ZTOTKKOd45PC7HHqCNDcxzpM6zScR08hq+2SPIEeAi5k7xDraV8+
4il0QXKUuq+BExu4R4SEn1kxATV9ArNLYDLonmiQAbiIBgDe1pLo+q8deR6geY/Jwg9506lzt/Ar
6rVnHVoKYHVt6/y5JWFbPnn08MbcZAozJ7WuS6dNGxiwgkx1Y9SjNsG5YaIfnoxUHNhE1HFkM95s
cmmt4XvuC+sJQoJmzRVK2KhIUPSAHlyo17jgG1/QaXEUL9jtFpyCghyzUDyjzzQSpLyZ0wkxhRZ6
J3La3Z/bdJ4sH+R2UKzXs8wd8wWFU+hirF3Enpx37uyWoogviZYn5WnssvZhKhJq3VHfeyZENLve
i/eGtkyTvGMSn4pXnelcPQn+n6un6AFqSeGTcYD5WmrPef1EnLDyH5TrO7Vke3+1Yx6sQWR3MaGB
TChSrjhgVPZewFc4XyYJGq35SgXH10y9w8CgVLSAjf0uQxGizWfrY9uWTIfcRh2uSNXkk+LV9Gg9
6wLj+zHRRTBSUdF1UegKMipb3llj0Go9Fc770UDPFfxK2tr4nxX/rBEzClRH0K7YWVB5sJ8NK5tf
+gWfzb1Kw8RXUQDcoI1fn0I/fWg+oJvRLzUxmz54VqGR0LOmFP4WFvK8Va2UzabkQ9Y7/o2Leedm
BsQPSFQfdkS+ZAYeyfnTqvEkUAwR4NzJ93Fn+4zKECQV3XShrTw/99dZ+xx5+FAE5n9jhzyDiD4o
EjNsYD6CaQBt7UQ4it6VXcJveIrHUtfFsLqf+BpBgpyAB1BQgSgz3qe27WmV9vTYysLphttXR+AT
LXIpMw/RuWvDRGMdMQGc/5hYUMsC670amn+Kg0C2knAQPm0yNX9XbHkAEcw1zCMgNGcAy1tePagU
6k++8z+jrbTRQSWTZ8XY9ECslSAzWqQC9a8V1vg8RsqepI6Hev5vGPAMlG5y2b0La0IzprhJQVoA
asIzUcXH4YjNynPTp6dg40MFI1q/WkLZNIeUZyjB2/4QjfovrIWjzA2L3Cd1Eaq6gh6ZhV1M75C1
JtY+75UFNeJIuLrHvSjU7aBOElMN84R53gXxFVH664GZn/BqWYAzHJfZ+G9Qi8dkoOc7c5jHKZXD
Dzss+5dnP6Jc7PL4PuPUaixlYM5+rkUHlO4yQaT+5y40o2xFOU5/0bOk1EgkJgUerGGjyTVxpqS5
AfDbOjwFl8YX/v108ER5RNNCx+V6tIlO5W4IGaGoHDkYDCxy4iMxrP9SGBrRcJ7OA/4tjSF2BpY3
UoL+jt7TEjvgWe9JlHzs0nZLraXaRQWmG6BCkvrCV7TUNYYYGuH2iSO1aR7/IRLpzi5bJI9xLh/p
0EpklyyVuoIOUoic0VXenZ4hIL9B//dix/KCYpjnpNS5XdwwJzoF7Fh1ikEnd0Ud83i2ItjwGK6n
sJKwbvJZAIH+sgJ9ehUq3R3qOfwU3kHCj9yphO/h+HMS+JW+QDguNksHhYC5/CY4clKwhCBtLF5u
p/+py0c+YgXTX41SsZ3CoxU94SdvfFTLlxTghik+7pe3pvG5WLdVxb/iy/ak7cIS54q2w82+bV6C
J5LLIOBh6qkSNt9rRYJYQtJSO2C0kPqosgD3Ea/U4S8EG3zxz0vJlRDsxT6byRdZHRNynZQMLTLp
KcZw/hhkmbAcNw91FNsiECz21CwUdE3MqsTUSYgVhzejR1QyYiR8DMBpCpRECBS4fgu77qz643+i
vNvnvdSM5Q0/Lpb8AQPhwUxA0O1m3hP8pSiDs8pXF2IOSE8qmYluavNVabNXtbI93b8ZMvUszICr
G2Pr0RPXNDlgS+DoKvVrQQ4jiW3iJCfhkCSpdts9GaJzRNyduImBgNwFCEmgxzp1FLRk7uyzJq1x
m7MBAAN67HJJPVrYYFRSUkSFq7tYoror4EU8cYsVVhHtfm3+V/4Jqo/RqzlLYFcGwzFFN9fiB5G/
ry31xgmpei7tL5aBf9s9vBfQ7+iTTCKMHK3fuWApxsK/cVvYKlv3zrDuPqEHV5gehLKWfsSk0ezi
y6+Kbf5w8YyBcxVUcE74UgB9mxMocKRUKmIf3UPHU5maNppY/NjquAaaul7jsdnkxC2ku07zh4cA
QUnpdForilD4BuN5bkr9TFv5Qj2zHuRjIi1injQvoO2njYf82y/+SxwC03yFsjgGdwa3Gru1RoSO
lVHrGNhlpU3jWi9HhLcgwERJukqspCwRdQDLEKOX4SbBje1TKAkHYejfDvzgkAT4ugiMDAo7VzsZ
MoPT6ctceLSo6Vl1UG81XJ/EX/Nea7GPjmQRVhhhJdvn3mxVzSNboPfDZjJZjocN1WBAt9nkg2jc
blir/H0EMQd1NgGzkPTUxtHmLCtPRcxQUfJGyEjQEB4n5ia2UBd1Wsn6ZYz1Gx7PZRsfbV25hTIq
1/snD8du0k6e6YuCKafgcpqwJZIZo2Jy3XmmUqoj1rYBsvEycIJX63LvTQyISqG0Lt+ZfYiKZClj
dQwaTNOXCiX3Nfv/JQ3ibX/F4pkOCAlTpIJoF3gc7NO79mapTSmVA6F/3vxLTpiK+iLlCRp7akGo
S+XI7YM4J+UlkIiTFhleBGw0Rht5DD7zRlBth2B+780JXXKy9/tgf15pZQYvNIJSHvom3rSgIIbh
PyMNjRPZZvXC25bPMVgCek3u2T11eR4GgN7ChyrpAhM3Bv7RA+kOlwp2RkFpExSYTtqBQaXyz1Se
56U/YmP5dVX81URuBO8fJFsO/gAq3zXwicdxmqnUrNvxnfY4adTARVYqwe9Rw9YJDTLaEQtHsBec
2t9ot9ya9HgXat8ATb8SgMt9MEJlTDXpSXX9/Gjrd/Z3fgSh20bnqmsWk7+k48D/Jaumn+A83bVW
8aviTif0xMpJW/sQ3SnIjfQeqFApuQUGfIUsgYKh2F8fgLVWn6WYqIZLQAUl/cCkAFv0XthHvO2W
lWR/BJn7BpV5NEE2VNYblmFWFl9S6VoqJGwuWDC96jKAIUmh2P4xkAehBwo04o87aslepBrpeRYT
9LtRd4h5G/RFGc2Y7WjMXiKBjy8FEwllPogTCWRFsS4KpQk1FJSed9bxx/GCiexezj46U11WzjqL
14MR+zxvWfJsOdCBK47gJ6Zubnci7AWh2ygmf7FGRWyZXUYRzCctqhfSWOVolIUMvEH2ESszyiz/
DvXgNu5RYbXC+UHUWWBc1xhRwOQLfRBePRPE3nz//ERAqFYKVATHjAcq+Addh/KCbQreNnRxOaZU
zDAyJl3P0a99P6AXXGDcrRMmfvmFxjZGCfza5i8jJI93PI72VU9c9Q4aT9PdtDkE2zX0zIe+K3CL
WqeLCD7Z9cHDt1FBnkwsDnRHaPsQn2bbvsKoQ6Uj4LMKPv+zIt0VqTuAusyImAG4s7rQ1mFF9ybc
NGriUux+BT5z16qUWFBWt+M0eDADVix4424l19NHOYuvXhyA0k07AQ24aRvXxwhyyzX+FOUSUDrb
USkMkaqjLFssjBVoECG9sqXRtZgD/83ubAlDCuHRZRzdLRr8ADc7yfc5sQjuDlojb7OSXwspOxuE
T6pW351zQ8KfcaLoK1mB6n2AMOzdWzb1o/JtCOELYZq25KkJmt/wj9SsCBiLc4wAmrgsNMssbpZO
PdSeyetgImmGQlTgzCq4wu5UN9clMrj536LCZbZRfyShXECzSnztxK7nzAjv2QrcVTg9ISf2R8/U
c7RbtGtd1E5sVEpgh5Q9OpY45SCro0LqHM4xRTntuye2/75H1RW9OAwWgj2rP8iheONQW8vLctrn
o11LkyLUr90HKyHcNjwxo1aDx+OZ/2iwR6blx5LzjhXeA8/JtYPSYIrpZNb7b5Yi3CETYHHhnHju
n3OAYYMoH+TRkAZQgZw0ko6ymNAqY/IbhSqy/GfYY94+L7H7S4EwWrEs/K4BOSJi+oDJgd1EpmFz
unu7UW17l4cnpi7ETX4DiL5PjvVrVKwilIKidHgqfwqnJOa8M3kM/YfuVMWn55+eHGSYK8AhpYua
btwma2tZyCYlecruLCygvJyBnq6agg3GDV9xc793EsjCj0/rBgWcY7sUUHJHm28tMp0hz5CYHdJa
9fUUsiwjjDoqtavvYhX+7QTS2wIeJCrHRttUJ8jii2LYbiiPyAPfyZa5OFxgvZnu1myxYVYr4sSJ
5+pB6ZrhzPyB8oKCNMqTcdf0WiqMl5pXRjrD04KYcotRJQOD2EU3ttL8CFfOlXNHf09lut8ddLP4
VNp5IzoqFwybpocBCQKikNNnZlUCKfbBH7QvEvlYtF1j2TJX18Y4+9A6Z0R5URageKvCkvm6rm7P
lX1SahAVG5f8k1e0Vn8hPJvyLT7PEr5TGqBSMgj/g2Xhd85P9iyl6GUIaCz0oU7brbdS5Y43sJnl
Pp30JzkjM/PBMpea6qSq7UkxQYA2Q7h6wTrVkvTb7mrvA8RbMX2L4+rg08o1ID08whiXAQObklcX
JeP+aLnjJnXmvEcy9BJpcf5yP4eYlvaDl+fItA1GQdX9y6PHVyBRFVwJZ2mKu5GQHA3Chatc4y/f
x/ryJPkdd4kXN8upG17SOa3T/eAxWt6Pb2Ujcbly+sKpPuLzlQkboWOYHaWk/TjWqxhEa3f555tq
X7R8MVcoQW6laxkLfQQXrCpzA2dib7Ssb74621zdnl61O6etjLJ4Km2PNRbQo9Ot4mKDjH2NrxZz
WF7op5wy2tdTGwVs1XmtfgfDWlixzh8Qk8/Q1cv18VAXngPodGpuRX1FbRSq2SXsqgfqF640JOxn
OdZRCi3X5CKsN2GFLWVsNgQJyf5p8cMP+/Cp77k2sxBwTBXXNVIOOs3R5ZmPk44Y5a/T1W4kV977
4AjwhcslrsoY0dJzin80HEaKmMX+GtLSblQfuMuKkDh4yKD1s3CfN5c0zIawvrVO+VtP5or8XNCK
7ZD+YQBVlzsj4HAYOTU0aWBTShLIx46E6RCkfqj/poxQI+ipW1/oUo1r/AkMwW/jXqTFV6t0wXlc
aBrxb497HGgeQ4vwszTDI6LL1PfOVAxHPmfFjhMK6XfTbn4EwVDApju+NtLUk0Jev5rW8AoTO8oY
BB3DMn4UztWOyzcLad1miw8FPHZQJ2iVblQfwSMracAjC3+SFafSw/sUjj3jxIF81BWxom41lcqf
HGzf/BTciPdvwr0GgG4nX65H8LQsTq+gGuO6fF7y9ttW6R1VgValXsVDYmWFqnFBVzI5W+kVry1r
dEVaqYkN84Bag3UGGF7S9EFIYMXeqByJVwhHY9jBtkt7AeS4rsMPMG8k3JNX6pK9gZLj4y1TjUrA
jR8gSoa5PDs+Gt6tpRMD8LhNjR9npPpUO+hKzgX7zHaJ2XQp6IVawwvgYYALk3q+Z4tFxUn1UYvp
moLG0z4hRpOqkpl5fW4v8FalvVJP00y69upJhwZoFMafgRW/DJPrIHkbtpebBYSoTNFeezrvJAse
VH1ynw1XdwNbpXxmb7q6Z9WSP9t3zPkyvERhxTG6e/C0QoWWp8MUxEZziVPeSWjICG3/s5deD3pJ
oIlWtGJ/mja3kxd+b4rNq29VsIukziwk2RJJJ1mlPT2scUBbaNK64A3D1dOJC/pckCRa5uCJ6Oy4
/YHVsthy2YQTWf402ykLf74jztXVGo/kVzM09wKHBfnFeK44vDOvXgxExu4vPz4UlWy5FrpSTukd
5QDQqhMNG8CvnN5YIuhkMiROVNX2dBU5b/g7np1LrYUqyEwxdyHbWyzvmnx4i1KmgKlK7PyhK4iT
9o8Vn81CafUuajhB//I4OQl5HM5kKw0+YKMfDrGV2JhfSsi0n7nIExavGIvFslwHTKAfJAmgsxnU
3N9njkx7tz3VTBp8RWIEMOM+LKzeQkCcib8mV+9Vyo/FE4r0Q78l7V/+7ndFezhlHxdZnubaW81O
kF7J9Il6vc2G0w5vq9ZqKgpPa+/3MGaUy7GobrOA8h1hmnflOJnUZt/Ivdl6Mdo4OjuMxyP3OQok
JF6P0jTmp+NM3pAoK1c2qQ5r3TnonYZ8oUOwMQyogRKR/TIraCXQonbf+qb1boMV2HJS8YJ1rPg+
fVH27wPj+PbUDL43nT4SRw1pyJUOJsJ8DMgFy34P89wX4dy+m1xKPmBc8ld1rszxcKXxcFuOoAVD
GUVwE2+CCLPlP3j1Wqplh56d8Qs4Yt70xsrFYYGt0lZf1xITB3cmYFiX3WfHgyVWrTjNxJdhz16R
COKSFwiv+UoYPoGRi9FPxK81IjjZ761kGSoMeNTm92GFhTesR33UCDEDUngMUmblIzGKgT3gmRA9
Pgy1RdFeB1sedIpz8Fzn796+9ukVHkrt7IL9ZrZUsboXyDJ5/jfi/JZpHD6vwPCx6g+5q0YjWQhI
2Mgy/IMxyUbPsyD9o+/9EwwwiGvpc3VDkLS7QoRBmAqaKJBj9HJoXS5pfUQyGOIqroJr0JJnF2oD
NlYkYGnZ2Hx+qH1418V6KhJe99+ZzYUbBYBnX9o7RJqcbG6yIvc5C7ltn5eibqX9qd702BWXC8Y5
d+sE/XTgSBzb6ERSCOMtmo0Ejz3BB7omb8D1N4TwZlFk4j+t0bTd2owpG6YcdybR4/a7RoTE6KdR
+xM5b8MMc+W/U52DmpumuinNjYUyF2MNP2zpDmKHPI5TzfZJ4RD0Fo06wGXxzvDzMipaNWT5sF0R
dyuIcEWEhVD8N9Jn8Yr55Ddx4l6oC25FqZhMI6IhpXiyCZzKzxPRG1SniuCP1W6FyxngBNje2I2Y
knyEZB43pwBTjz7LV7SJYgPgJs/zT0rO3X+ePWphJFoSRMIi3AW5M6dvPcfnpsQ5irz0nQXgFWNj
mORxFd3ZNUmUbpwvk+ItVSjig6akgHdrwnF7/T9X4lp29YlaLF3HmxpdQWFWGw72vdDt9PkEQprQ
abFP+X1fcfc0vsidcpdbGWEQCS9Xratuh4mPM/+dF/QY89dfxg0vk2XaP/yMqbsZ7w+FB5S2CI/R
sG1BrJXEcDnqFvxcyCSWEa83bDZX8HFSVE1DkgRXGijFYy4cC6aTYG605HjwSFR6ECid3Tlsbwd3
nQjagusIAqBPNozAPSM/y/puUlVOiSKfATKz/uV3RD/31Lw263TJazGnq3GiI4fJglqBxvFMuU50
jL1BK2Y17v3k/rEyN0REPfGM1Tvud485/Bzrjg1+m6V6yQAudJCM0pBQOohmdMCG88/d6gEoeyUr
xzo2wrC2v43tml+mxJbDei5G1FqDXyA2rEPNKF0PZdeRhzawt/YLhAI/eGW7X5ihNAT1mpa/EErd
QnEr0KEPUn4Xv8HNOXJatVrCQfBTEZlkZSs3/UE9scbjFEm3a8smjfUwcv65bfPN72lgf118JjCf
6wbfHjslsj8phRKqI4TKKvpCSqdwZ8jRTDF6UPyymQdt0NIDiPf8IHgdc1dY7/eveqZ0Amp9/a22
aK8fKnwNXVeHMx3tJ+VRPZkD8xG3hmASyQnca7hDoEjZ45Mai0YwEUZp9DS6Niq7rZYr4wiKX9J4
YUJHD3dAltBOg+QqZNu7wsRi45ffTRW9LwIgyu8W7Zot4kSzCp/uNLcEBRMIBw807Y8fidf2+5ws
jpQPT/iV/ycuzCeZ3H+kyanh8O6PAWA3f7VoriXJKIufnLySw09TWcTNOwJKxZJzt83h1we2JHAH
VpcWiTayKupul+lCk+TzEGBpnnW7E5pmx6AKkNK4f3BHlx1ZXDAzJf1ao7ncptvhq5f3q4xOvLHD
xJfVj6RqvrcrxPv0NT8OCmh0wmQrJGq3A8iQCUboOtba6++tsd+P8M+dwhTESWCKoc7PwFRiEXY4
9nUQydp0YZ/Wmfbx9DJIrmRIYsAG/AWap3LKu6hH8UiFLUqTtsPxPM/l26QVpkJExp0gRmbUMt0m
qHzzK2sceVkfv7bNr/LWew/LUQ5mcmiXfRamkdcgmDDro+arEFaqww7xHnoGlhr572XpnN7LDcjE
1kW3BmmKMs8Bdkq8BdJyE0p+W76VEV+10Vbul0nd2fRFGSy9Bzt+NA0D9UaEdMckluh8MBjkBjwu
BUU66I5zclq6J4BcpPTPeqB7fWSJI36PdlFHmB9qWPIuc/LYUXq53XaVmkr5Nzd8r1rd0pZgYXW5
2SK38vFs+Ha75n6chFG/j914jCPPjlkTNV2z9z55C81OYhUFb1Lofg44VxMnlI49oyzaTOG3z7Zq
6ruSFREwXdN4vbBxsSBuET3SDPZJzrhYTuT210e3doqhTvYpt3pf7TsW40XCO5qeGXMGj03MCG54
BQ/DHoYubXnqZrM0uuidSonRQfIQJnz8HGDUFhOUbIb+5qur3n5psVVLRRkVN1UeJzN476RIbW8Q
Xlfqb/NWs3Mfj4GEjZ4SFmZVmKcc3nXWawlV0Ckgb64tl4070KfvW5zqTu9nak1Tq6FO7AXu7foj
EJpeWD1N6pOQLmif2LohcS+RAVcORZO0p6GlWnEvbzfaMtjUYGj47ujvruGTCYJK8raSiVrdkDaZ
T82CLaSsk9DvJLjohni90k/CwR7FxP2Sf6r7bhXMjo7qbIVGa2QvK8L6GKOPrGVbH0GnHUwuhThl
rjLNxeXL2WclO1R/KHr1RJ/OsfBIYCekVpdxIfvRoxHVR02QZStGv9QiqM8Cnvsn+wZ0GjRDtEDF
CKw2tL2qB2UGBqn0bal7A3ZzpChdjURKke7vC9oTEa9lpZjNBE/TjxfiVd8RB9JrVqtlUFoTEfTM
JXiC7E821a2ve5LIX2ljFkbvSUrMWNbT3W7U60Gpg3ettSDwoyqGKlxXhiGtCcE+3D3eb9LDsNJC
0g9tcY9J3vLr3mPipwoJHbjFV0va2njpyZex+oWb17afrOjyqZD2WRrlhY34oGHtTVeGe+PcvMxK
xWEIPd1St1hLcJ1r9+x0xLu73dPzjmxAjr9LSJHMVPCdqujOcLiPp6yWyhcL+t9wvzlyBhs9oCxk
C6mg5aMFESB11QVsOBoD+6klPByln1+6JHdWExluvY5rXhiBINNIHrdhlYT8Ka7DILRetuaZoADc
YR3Up1hLYFa9JCQWcieC8LqARmS2E2Q7B1nagcDgEsb8Po2Agln1lkG+8WRwIBuDHKfNIF3tD/yW
0CIF/Ol+fZ94ZGBxskHia6kV2aHUYPyeRdFwtS9zzh6iGCkI6IJS4cMcejs5SBU+6zL9+DrZE1oq
y6zJkFg71zo0IohXyOnpWhjm1CUmKtxeCiLKJsB0XEh4n13RglZK9PkCm90T4MlZWQFF9gelNKO/
IygrIbsPKYhPiAHIFdO9/qGq6FXui1+jwAHuhfaQ1lqBQIKLp/gckDDM6t7aTeiICtsXg4oMqNuQ
PVHLFBrtfUwNLM7SZgKEOTnXLPoFviHQTBqJCeKnWCgB5Bj6NGmR8nztPT3xATDJVq2+FN1TFe0P
xPeRdIALeyA+GfVc7D6GG/YP7HtzmHbyJIzkxjYajEvMquZFqeY+rAeO/k6PBg5QkNFy3yMeFkSz
TdXOZ/aWBD+UywoXwae9A0aIW8sCXNQSyWRPL37K8ptP7say06ZuiFrvSUBFRhfUo0YDskg6J9vr
P+m8DKhExbaxLGuT0pKAg8JRRYsaXg9xBmvts9VDbh4DHCZqllnQ46PFkniUSyiPjdSdPksf6Uve
68/tnnOOVKjthWt1+kA5zdgnouv9BfcD2ZuAVF6uZ6HF/u9UOsBCeNPlP9aGVJnJpksmKBawK8a7
l9tDurvBPjwMxnPq7fAFJvgsU61r+Ph3ssChQGjn7Magrp8Xv0Hgbv+6Yac97eeaW6x1xmLEWyy+
gRcPQ/vBjmG+TNdvtZQHBny+ztL9ZmFFjuTW3ephtF8Mrzl9r76cM34PqBaQubAJuGPp+yAVJ/E0
vc0ZjmuUgRT8rMTPpe2Bc7xM3cDGEZnYkCHZeu6hMfkOwWf/rxm56Jfu1RI7q8iI2E49iE1I69PH
4zDFJuIrLJUtAuW1TSmjksHQi9PZC3d3XoHTH0NuTq2EPQkfNrVOqTuBpE/whLWrI9PfGnqGr4Fn
TO6AJX0NBCNmFsxr5gPD4HrV9rkYasBdjqNu620r0Eix5tTQyNQbwKgOp+ldpq/5jy34NBs8Nn9Q
VFDYQyG9Rew5bJLhG6UjzWIG3AVWT930iQ8UYvaWed5bN4ZdZmj5fEp9zRiA5wIFxDZF0MvTj+NE
DFLasUQagssmbR46iZHwkuRnJ3TEGhMaDolWDiz4s6/OqmEnG1gpnjnJXuOUohm+ae6gPD/wXWx3
RsJAcyTM97sjrvFjpWjpifVNOVrj/jKzRbbB2nkWWMi2WTUDTpYspkrDJI9sSc2fMG/FZ/E4J98R
U30uxp62c991c1sawQ0UBl73X0GaWOZYkeAIDKRGKMmXhbZzaukgXgIMiQmmpif/+rGrjDLsPmse
QdrL86z05kWegDpexkST84/O0EAPhDr7vZX9H0sQ7iLjdJtOyxHA3yRbY3UKTc+YMxDuIRy/495T
0YH2fIpSaQlaU4P874xBW0vhX1K+iJ8KXgb/JSnEVBYbb/7ChI7LY5jEmn8seMOZkf47hdJWKRWD
YOBdQsf3g5kmHMXwj3xo3xVLSDuzj3GGWAvxHHf/KXJLDpeg2y1TMsX4mnxXLGPzlxwnE8ZS6MSN
cUEA/azgHNMs0hxErhfGzICAoKTMza7g/ClaZbuehu6NCvN9JOCqZR3lXMBsOquT1Z3RQkmPwS4p
lKmWf1ulAdcc51sb8usyJ+p/lhefRupjwn/fB3tYM/zooeG+l+AT3JI9fJhkfn1O1eUTpnLkKISh
Ym0YacglA9+ESTduhvWrhTgMeMU4ESD+TSAuO/SVpE8g/6UQqA4sMh1ln40G8smuMJIiS9RbKYmv
hFG6q4692MRG0SY43MFeOWb1OkfsrZhTEnbpJUJgQESl2DsIVdI4b+wDtrs6Z610ePx59tursajF
glpxoiw6Tj5lxmJ5HJZ7hLvqzxpUvJCYIpEK3O9pNT0fTB/yNx34Mxx+v1LQIB2lGkVXB21uEOaC
tk1Wx1VaFaBqjkHeg97N1iGEYc3fgqVYCC2ijpBbmnsj0RwwURSCmYOHa3AScrajlgW7xhk5m4XX
PYIBVKtH7XWLjM5i0R+ucncfHCJsvXb7M4wtMGNSj2txFmNkySbIW4xPKfYAuXvpB4FiGTnRMLz3
Cf+YP2HW8eep6iJGKE78rDLwoi9H9iBo2XRDxr9qCfPk5gg+Hym7k3PuDMgiOJvNdHIW9yjAmAKq
C5x+ZiYoB6DPtKZyj/NtthLxUxIIcu0DlhhSH0Zit+Y7RHCvP86L+kcj64zj60H9YU2s/wmeBXcz
mudQaiYVmtvm9Q3pjjvgHbenVOe1YTfmw4hc12/bzeE1S2a3k2YJbVARTZQCIO1ybKfQFXpOrCVa
GXJCzQGIuVrZQYY4Kq05dQtOJ98yxpSUPYbP5Kpzw9ln0OGWQYOJk012tQkn9iArYobN75hpQU4G
0bFt/oZ5OR0r6SpCW/vz/x3CVU/9wBMKt+bGcm9ulSVinEzuvSVmqI5Ek6g6XcnXr/9FJ5nAS963
vE81Fd5RzqfJ3DxF8oYnX1eN37nk3fEs1qHh7o9EYkRf09pw4AobEsBQtOcjztsabYRPcEvMEDL1
oKYRMYoy2fVm5eyL99ccDglqNsR2Qk7mclIclA8OKN6BDcqItryF8u/RGIHmY1feVJYBqrTtcbsy
JTkOlFux9kQGxJ+YSr/oGAmh+qvrLfnyL0babVsPm/RWTAP9bDwbDGDvsFUlKvE4uPKThq//p8Mm
A4EO/LEohocMxaYzRnfnuOayjtixGya1zFpndK5ebe6tlZqboXHfbn6JHZTndsNFA45R1rZHUviO
EWkP22MTOhZSq38muCNDe9+G8GXmpqbmbJN6fTXVFyS7VMETVuu/b9IRKzcuDLbMQWfNpe61aqfh
7Ct8n7PWB3LW1hLOnB5bje6BdYZBGmtRid8YFyJEAxrmQZ3dJPvioUoSPDGcSSOhOAoTlPtbb/kJ
vecgH9UVwULLPx8DTI31xYgQrdqSUjbMhxq+UUWPWM0suC89rz8igTPxv8Maj0D+5KiP9a2+rml4
+7uHjVh639iU8gSvtwCNH2VzIjsRk/CjIM8F7X3CQ6WcNdZ22bcfm67vl7yWSNfUMJIz3bArwhj/
iqHYkAN1jvBaPS9KEoBvCv4Qt035JgIMU++31EF23tVbJCFvkm48B5ZtjGM16DXNuETUWLuje9U6
M8mQzytNzWcT2F9h+ng2+i8/vYxnYbr7mplY/dJzJBozgXEkxnc2ncj4wSkrImc8ndxWb1WfOYIP
e9uQSWnQHceiU3xzF/BoSFpecg1oRcf43QOqbr+vMDMpYjaDMXGRbAShMLxcTU9hUGkiR6cmL6BT
Sfw6zkhdYC8iNjfw8fKx7//VqhmQ+vQZxeJOgZ1Jw1FoYKCy12zS1DzE19m77RpsBfR6QM0D2wuK
peL0aqTcty+G4884PpXGPkJjqH8B16Jye5nyu0Gl9rdqQsSrrg2BtDr0Az9S9r92zzU8ub40i1sg
c3QPeHAnCpdhCDawx3kTOGkJuc8+qLbAGYfgu6vddxaEMCzLcDZ0uq0Pu0B3tyygpqLhGWeGqD8r
H9c/9+u28br25m1B3QiIIkjznJTGxj1Z4euT30ISNgH57mME2IZl+DRKvaTSe8ved/J6iCFG4cls
vvwfXa0zGW73C5bJi8uf3F1uPPIaT7sldTPpRGuU//npt8EKk2hc0CZiDJU60uy2XB8WnmHVOeN9
6/qFIoNUamrWtPWbUy5UdiGicb++Ajd5Z2g3EeuDKIykAw6R6UUiVm8R1Yd3DYbE4nl23BooZqx0
CKi1I63dbeQkEEduLrSlt36UaDsxB//SpLCrPDjWpLS+1K3khU9dKi320jtD0E0CMGM2+0rJulJ3
z2uzJCYUUikox+RuVmJGCeXywAHS1Sn8VoY3qhXZT/VDyc0ktyaSptJfc7m3WOg4qH7AS1+9nn0b
xzqbSQTaBDsO9uy6bXjXcJTKiI5DzHbx+xNfxGH2oq+yU9808/X17s1dyUp33d+MFQQ/cSNiwovx
2R6JAf9sLDoYh7Ivsd7IqZCiUgod76BXQNJpmxU6EaNldjpN4//DshhfVSejmohvOLd2ttWqsC6N
LBqtAfAi1q0UncjUUS3Mu+1LvaGW/rwvpd+HcHyT6mdZUyILLsmb+SUdVpmhBRB3NWyYdvMF6DLh
ib1gcRnjZ8CpKiM+mCz8i0EFxeosDrO0Zixz5x8wAC5nyPrrnfHJGox4qxs6f9zz/ZqVjQSdCV7M
MbJHK1nukwIctsFlvX9hmFydgYg2zm/FRFVXmQcfKQfUUFScUNFZeGEuja4rxRlDL0QLZYSUX5an
AyItoJeE00gqD1wi3+/nLI2R6jWnXkOUVAyvk1F6SVqCSAJcR41gz58/GwH3GLHED0uZ1yiYiVg3
10g0RwiIx9+PeRYhaQRHSH1KCYrvI/qog6r/NvDRkDBJkeM9ZhAAW2nwiZvQGRv4Beto67B8GpAl
qXpVocIub3I3me6vo8ZDLwKAXDdF9clnVrMjQIBorhZ7/37T+7lpsW4Lz0Oe/0oO1rtUV1tCgFMW
PDH1jB+Ke9XOtnI57aUJm3DI+M7xZ9OAKLABrRARIHlbLkFpLYprCc6vyGaR24PugcFZBCKIY2YH
jOclmGcOQrbZxj++GS0oJPOJ9AnCAS8ZI/vMCOvBk9KghQTU1GvOxMwxVivASCJqKxTiMUVc5SE3
MaBivcI4YA6DpBpJXb5/92kPWOX8ieqLt93/5Q6N6k9aSjhiPNcsSic4KHwPmT70MSidmP5nhaw4
/X71Oy8rxt3w5Y+hIa0Qs2VIHAmS9FNGvDyICWb1E4hfEn6SEW2ejsx5grHL6So1+oQdeBj3k4qm
6nFCbwgBdb/sjJ7dMGR4Psf4neBzoK8H6MvXjJZyylLRNFFlqa4JL46K5M6f70pwjNCGAo8yBKW5
rB5f3dvt1yVjQwaBSUZrpyadkSqTrhEvnrSfoPeanN7luPHLc5KN+38l3cdraswL9BL9Di/aper3
hUiABNPMLm/0cBAEc27TDdPUj4klBJB35rdqK8WS73Gr7qAKxmtsaNg7CRyeDH5hjyIEvy3pOvOO
NCk1zvByftLLqFvZmVRvImMJA7KKev1WS5/ulrJmoS9Jg7af9B5vzPau5IKxWuQEHkQUymX1JPyI
6POJyqTphZLMzedv/vouS5FREw64xlNUjMJsU6HS3Yy1r2sKwybp7sodln9M3d7VuCE/Qubs812O
8Ec12LmJ81jDMGzNs4X66bISvA/Lgq+Hzta88xELecXAglPYDmzrTw4byRdp+UvcbM75U1WPSvCn
IMbwuImcvmpdnDxv9twiVxcvR+oBsuB5rIh9toIpw4cs++kjey5ayqGAt6sCl2Is45HNIvwqa2Qf
3Tzs/T/f+uU4eRSRdqCZIPCZFRV4YhM0uQtjoXaj3/us0WkdDYR+c+N9BncHSfYGbk65cbiCPgIe
+HaZCQkVnr1ODDswm/Ss8LrJbvKwLAgz5YpkP39NjdFQklj9T/7A1ekqTa4NRwWmUgEme3TqGc9x
ZS+kd7lV7FQFaKJKAn3arYnkVjKFMlN610MflJpMu42aCAtMMLSP0kLDMrF52SRy65pI4v9toTVx
TvSQ8f7lS/Nth8tJqNsaRHxZdubJQzU7OQWFExW4x220P/W2ZHKbcrEdJT3Jv3GacyISb1FhXYTZ
bKjPGCnWgxxi2fr99J8nhiHdI4DqX+cr8S08jlz4oVIVFPm4LqEEcAceDxpy33EspF1YS9Y5eujQ
O7VnqqzmF9nIyXWHpJwI1ffSbLLdoQ7O/iq2pJ7xZZWzQTYzxXgkStdFHzyguY+TC/wX3cKNBlL5
8vhtjKL1XhcsZUcZSF++V5qcTQ/drCn+sjH1anPYVDN80RECIAuL2lrNHR0YfcBtiVsv6MBMoq0k
SrsR4LMxwk1INqPwxVEsjR1FELfB0GxKu4QvFvrOu/xDCD4X/+wZn7joZqv1o4lkWINXe1qj9yJ4
BRMIH4L46nNh7npEkaQVtd3CfZe1KKcHksqDIOYqe502T5/+wHOjU1Qyrq+tFtwM2D4Xdxay0umL
wZrt2mm2xdbvBtrh+S58fMNT9dn+KVlVSuvbZiyjgXlT57Ahd3OYGBhTxCT2n0dqQ+6Vql2n4h1U
iu0OrsWumBNF6SUK5i597uDIFWkf/tumfIYAeOYCcJQcoMZmqUlek0UKDP0FE/AePqmOjmj/xp4F
QuM/LKQtrdKkb6n9QkHGuJ6QDFccTP5eGLc4q5DXIwz/ViJJx8+AA019vGHaqh8elAZz2OjEWwpm
h5enCkR4QEsENNyKc1Z6VIM+7ZIvwE8bHh+gRAxd3EX9KpilYuBatJYC7ZudBhyi1nV+Yxagfm6+
jdbq5aefDaqNpmgPBUvWmyufm6MePC1pI1ucpZDLDKZL3/eTvNeFevnbC/tuZ7QvwpMv1DZTaGXC
QPDdF0FNU69PJzwakO/FtNZ4cl4KnEaP+BzQ7G21i4iNYvwugs5/BluLX1VSayAQ+shwDuaNdHKw
e8lrUqI9p5gPMLcAAFYKHxj0KcqchGRJs/IHoJDERsa6LdKPgEuuX5eqFJlYpGeId4oCTXoqUoep
8H13GnvX7nCwOynKF4n/uQytJflOJcIw3VYwISOZBzLocWWi8YpY5A21AUJJvJzVPv12ugpZBBhe
wSyntfn1JNwlr5yWJXbRVGMBs6SrvEEjz8pIL8ub7eerDaUhCyJb/qLmHql+kWpg0TqWjr55B7tk
y7GMar53zhTDTUgckA7x1lBesoCaGS00Bg6w1MfjEEDdNSemLdJ+rgkcNqWZWRR5WJoY540Sgs5L
VmaggD4bL7fWDB50exbFKgo/mfSwRTAeum2usY/lzgCy8AXLlCGKC4TwfKVMrj9V+kgdwK06rsjt
0O6ltbztFEDszT4cc/CehuvVL3bAMZEv14aIOJIMsu/7K22MuEg2dlWD41qDnrPwAXE8Ahsf5JQF
rL2I+wooqEZEpXFALw/U/vusdHnCkZzRk5oG2bqyOj2svlRF4V8Um/Sb9zr05Yqy0e5sSD9EnJV7
SZDYvoq7iaTY5fX/dcyhW2oUPT/gToZUpTpoIttxY4oxKmBvPhAgFKg0DtyHSLgnAC/JccD+LEhT
yWmMuXYd49E+R5JXPc+z3UCfL71x42ftB9nXO/ta5kMS0TY2sUccO/reqRMduie3qMjYgBBfwzjP
k9u/sVOvtbfNEBZ/2XcarQaNhy/RoEL/VdSMzH89UEWoNSmRlsHGJ8C7QYvaWXWHZqT5F6Z9BiJ5
ndObWGyjLOK/NAo1QRR+vmvk246lxuhvg4+pdvYG9VhbxGVcyIonC3AnSc2AF3x0RxBeE5512qms
4ygDcoXo8q9C+C83wL+OG3RplMRIqSYdHrmIrUJJ1m9SX8U8edygzOHN/3ghzYOAnravxohCV70s
/reLvCzaO9b4WPAPUuvh/xyRyChrEMPkbQ8aG7Cz1ASDYdnkOkTYzmlivcMzb1uIdAIOO2GIAYK3
w0N4WkTGEIrVu6O29/un21ruSJuFRvF3f7wJ9GZF34Qsfh7fX1TC2g4oMj8R7DbJV0OeQPVJexm3
/DqYcRKO0WXjeavrs/IAxvpd8rGa3WQIhIXMY8WEed97mDPwUEBTGYDnEX8zJsRyjlZwqB2klyG3
xpf4maJFtttR+zNrF05oojVGdY4KMyYtVQ1v6cwL7+nPmwjPpTlGS5PRuGL0atFMbQwx/WgMmlzA
xIyYbQExrPtGWsEeEsXjFAy50D2XIXG6RRLnjwVOBA8UK8jW4GL76bjt4dExP65jxkYKW/LGEHTC
dXJD/rujzeWjna86m/jG3ST3OopsSrkHztwgSB2kQ3sFVR2eWI4S2+SuJFNoV+I6oSaHT/0s1/zW
0J+MW9la/0k4LkcFFMb5nNjhl/sZ98Ng9l9pE71eYGi5ZOdJtt0v7MKI60aU8RGL+YlCaRlk130D
l5T/+EGbdb8bRuG0kU7Vn4XpDpGt1qQUcZneSLgxCy8ktwiL/Rp/K2DW8mFngZFQgPGyfh8tWVKr
xxE1KcY1X9ZDhfc0RDvtX9haMkg5rjP1fASPcSwBLfE3VF0mtRPiPZSYrSO10gtef2b9YvQhA8bU
dTxrB3qPacPI2i7dDFRcw3ZE9tOe43bYITbtNAnq/8cXaGKDdLdYuPMIxSwu4Ob47SSsRz5LOgHf
i4K2Ld+8zQDVKJ8OJDEIhykI3TpIo6vPtqnw79vmPrM/IgGDeLKLryaKxgADzj7ZiMoWfteKJUqh
qsBwzzcIB2iYIPxxL1RdBorC1Kgs3eO6rPOdrIawqltKflKfJvLfUENO8BR3vPBLAxSbFQbKcIfD
yKiTkety/tGoP8nnb7jOByxEvKrTYbeIWQSwzCgnUPMEkU0RZdKngORt2mdQAG8KF/33a6aIgynJ
prVJdCzNenx/rJ6MfqPz8aJgPl0KRqeQxT/0gOgsh5FWFCJBbiFq0e53BtFEX+XaLZtAnbu4bV34
go5CvXksdRi+He/0GrPQ9MKRpblQBBybVuVkz0fmaS7Gn5SM/5FPXKc8dgEIt6KP21ImowbMso+T
aptAXQ7P80KMyEY5Z95bGjXrywOt982RCAaT1LrDbsBwyOTuqz3ANntx4zplPyw6uIVOPV2vLRFz
h4qbxegoAqYdZaMfnCaR/QrrxIhuvPzmYJ53nGKtbRvteIo5BQ9aVKqUYx/lZ+j07tCLSJhOux8S
P/o1gIhBOPaFR+Yum4Wyxz/2IjZ2ti5fFfGAsWfbdF/cgp3qE/r0Xh5x6lycX+wHGcMKc7qzWmcG
2bqRvbGhLt3toJ5v7Z/7Pjevb5QxFA6sQcH8YVvkZi40AGFER+9sNaJCvNFEUFGBqRHc3Nhusbve
CgB+dI8KtXnY1E/05ktLSeXHnkB7eS1XDMpwcKE+p6a19X+iUp4yaRcZeuF50oueGqFbtSON5Xcj
LF/YNT6JKqu40gBkmOYtO+a6iUh+2fLGW4hoPnktINC1Vd10clken0sSzwVx1VMzBPzoCKKf8tMv
8eTtb1Bu78PNjivaphlkXpo2MyEllbXfQCn8lPiMsF/QIyF7+hTZ7TzdXWNuJUnEN5M5BfCAvzuv
tcRdaGVQWIz6cnvL6rhIpRimarLJ1ba9Eg1OkeXRptRNmnip0XzXDngHjJW0aMMFJmAiMYacDLRs
WFQ/cL7K4/q6DioLWwEL2/h8acbg4F5kjW3KINlRgJQHBR9utvxOc0cAmjBQA2Ubd7TOCzjaNcXn
ahJWkKDPyYymfsQ+IGzM3o6mcnHPZy9xbKaMv4OHaRpgKtpYQ/wmKCGKizylV/f9sV3hJbOHWd0b
G4znDNKRGBn5IkFnxS0ZJV/FvTG/GJGh6t5CKqWytl+igZS2eXRqHqwYr6ugxY8ww5AcLStHrgal
4s4Gas4VmU1p+7Y1BarsrkNF8DDJxicrsq1h667R8bYCTTXHIlFVBjsepT/dKWII43T6ouc8sIrI
yih1WjTQ79xdHrEniriOWFwHc00cKoXslkVemnvnePg7Q9xH7c0+tujAUi1kfRxvT66H/wyklvzl
RniSCKEQkXe60t8rmh1KQRLnVCJohjYNXVLEMco6pu5ZeY0fJeE4N4afKe6+StZnNWCnV0Hf9v4G
IgyUsWSFC5re88SLBA0enouoW9RHK1P33GvVoyIKAv9CNzU6RTeJ7z7taaKCUpYKmalxW3jfokgj
wz7gISQViez49WdikWohJVoeg2jITgnBopLGo5dQFOxO7NxQZxj/OJcZc2n06QZLJ5x3v9CgIFNO
Wk1tG4EQQmT2jyMiylt6l0WCgOxPY0xvxUD9VxZ8s8wUqxDY7wmnoAGxn7fx22hQswiv67F2zrg1
OONVgwauJYV9bv43ETzWK+IfigDsigN5hIqlCHsL4d3z1QgwmiUVKpfOTGx2SJY0iEJmipHBsuZE
0UAI+YKE9jFnhFxV3f8ayvWt5ER+o7AVh1W0oVL4soSKuIap6mzuT8mmap3bXyxtlh1wBGa54xKd
TR3gplGcRKwLtIN5B2JLbLd4RlR/vKAdviKFoMqBPE/4n4j9pT/y097LQqh2bjUbUDYLl2bCvOT+
nHuGPBjPOdXx2hiuPjhFgLh5ICyvwtazucl7iRF/1B0mms98+pHO/S/2D7YjgVJ695aSh3sJZiTe
7SJyBDftKvkCNj7Vtwg+pC7n9V59BpJDS6xaQwIE5++6FltlRs6RSCUnvz5kQ8KbkDYJqZj8wPLc
X3j8KGYf/RtROXubDHGK3265E7G0C40NRsvMkdA7Qdfq4+cRVvKnGkB/+IOBVuVMwfUE+CI1jHFH
zWX/NbeK8MK0Swp4NKgbkHPAwbqH1gBeiPXlxJqidsVswOyiNSM/5xbUni7uYMT5KZj551Ashx2i
fa4MU2rdlOCWuNI2I307i9oC9sp/UTcSmpBjKb0Iu78EgH1qx+VvOq9MCkhFuXo0h/Gf1etCFDmU
qNKmRS1fPAlnTAxpr7QNDFV6gO4wIKEhWiZ0f0rFC8OO0gpZ6EuhlLVBdXU4vKSMOYIfOHTxjdoh
zldWCLys44OGAxi7WtIODWwO999HpoF3MdC1Moi8ExT0bJYYL6GJF9+u4TTN49b2KzxRpAqjA8nJ
nUGtMfQuMZJGlijyOHrV0MSc6N8EZ1vq83+BNNk4ZzDupGSVzYCIDSsIug6Grg9d2JSi+C++Pb7K
YELaFxjZTYWYgJOJ3zZwgP1xilVCUD94hyQqBrbeHjM3iORn648toH1JIzcBraeQ57FZaB3ap7np
xne13kwGCkGE38TfeHBQw4XJYwUCfcdPcK+XOZAeAnm2qd8gHLVyvXCJQFtVDgExpV4b8vj9B2To
FxkNY2S74R2PQmIpgi1FFO1oxqgs6iir043Vp9U/J/6vXArO7JW5xszc4UmCwYjTE8pFp/E8KDGA
/QLZzfkKgFFLgMEvsNXmWV+LFkIVPl6hdkOC+cUb7KKdbuKFv5qZM8af2HrG5B9O1n92E+Lt6ly1
YB5hGHT33h3XpBIaN1TG33EUFdbJ63+zwqLkgvqjuFqESzJz405HC94gdg3x5e/ZpUL6c2t8RHP3
lQIyeHF/hpTs4Fd5WOR7NCvR9cHnNchOj+1y6vVS78dvjeyLduh4UQQTVGmzaUDd6pxW7XfK+QmR
tMa1JEs6azXx+TC0BE2E+AlOlaw0xYvlsUqKQVJwx0Hf1jS1pLjwFn9Tffp2kN7mJcaYE9MrmKai
/BVpTLpri17Bu68Dyr98Ea5xV5Iek2v+72Xe8vZpQ65puSnd5iUO/MFOyzpV6GF38VAR97HcypdX
btJGzFaIaUYXlk/1fwODZbeoHG3dvcU65rXDRwjo8JFlfB/CPsykTilj4/LCVzPbv/CVbDuJPv2y
XrBGb/sewWkcZ908ypK47NRPOUyorVOIqIMz5kL/NfGb89BpCB3gOoeHPy4TfA/by2D8woMsq3ln
wUkvBaE3lNtyaYp47B5/82xc09NMewDRYvTL2wVEnD+U6+sWLojj6z537ON4+c+SyRt/9soylBMe
5w4xFmTJGonrheMjTz1SNEVj0mOMo4abl6bYCVm/LLJl8lzxg5lIoXnEjpAK0BFtoyctwHOA4dos
y3X6LHtd5AyyxfLPVZpU3qgy+sKaNfpHj0EHy00J33esZW/5UdVkDimvqpKUUKdypbqLZOQ2/PHy
wy7L1tg6oWaUejadJOyHR+PTDOiAGZH8Ssy4/XqXRSAOV9IT5iGMh9xfgSIPvR4pLL97xGpPPnTE
7QRqhMuvLgheCZFZTD8jFKdis7bERTK+Y2+mEaDioz6lW/MjQ2LOdVXnssBJgqkH+IO92SlsWqRa
p5Q2ziy9UlJlUUVBx+QQ6awTT0N9N2OPAQ5MSFqdQKUxByP2HMEc/nJDIz3JaelsyDlINSUcjI1X
nxGgZtFXAwt2mJz1WGQ3XGdo08J3vlqUee1wfcxula1Q7ZExYukVI/6+wwYCSdOHNAtCluXG8PKm
mkDrEy//XKrDpnL356B9Xu3HLkBNAwYONIVyztZ9c96F4dyCWG5wlcNIKSUuqRFuCTmQAzMAbKE1
M3MBdQpdz6VPrB7chJ++Ni5eFLH0lDWRHXg7sprxiCiauLcSTopWfA3mlPmBiAgl4c7ORUrKAzpF
+IAazp1iVfD5MZAYYnlXAesUZrPG6MRyZcZnW2X5SU962bH2P/VOEcgjdKKVTu9iuiJduOPAgdXW
y3beiKDxyFTZ8d9ZsFpmyhvTjLik8nxAwRr6LAziXxNoElixTeuaJWYL/HuFKY68e8keDh3wWtLT
NrZsFLIRKU3sUWYBpY2/kDzT4p2oBDljgUnYiGm6OPvPDQ9gtwrYDlsrleT7D/CPdlwA1PMF1h2c
gROumDDdlng9/uklafDdnh+Y1HyewE86zwl+FoiA8vj63sSK3DI4GWdq8PkeUadt9Vom9fcIRZiC
MVENQrzAfj8zQ4s24GpV6/TkbmIhKhjQikSfMTQv7piOJaHk9iM8xiePgrYcDmdWD3vE4gSsrH9k
qOOKt5jnfH7sgjhV0Hk2c3lJDyc0DXUK2AatYF8SzbVRwHHBgH+rny4TORTjGWPXTkDHwYKtIUBq
BesVtnXfjBKFr+1mBkTbN2FrqNvjcq+TK55LW0H1JrvtlNzJb9s89sINz+UdujMzjEWk33dNpMUt
UCPv5BQGuMlBIq+t0YjUjfP0IJPIwj8zbzJHT9Ep+C/qJhr3vVAo6dQEeit5AYT3obCsPO4v6EVk
u4wbYNxsu+SdSVpM7D4E2sqkxi61jwBP0Z/3QAhipjyDkaA1/rV0HJy5HnRk9rZKyNT4NsmIvC/v
deR4UvHWgMpFrB97JB/F7Bf3lGXHC1mrqvazZk2NKSpq8c7JYcVHzv/URvpwPPyEmC9f62gTV+rj
fjvCv2kRPGW1C2ZsxlAesn2JwEAWgaG2dU6X2hLFhP7xG5nly84SMqsOBN/sqOCOMkaKSsTFN6CM
k/GDEHBmO5mj1vM4RK5eJG4ifCe+A9eR4s9WRq4GQaMFtmWw/R+GyXbZBWvXXyOvq+R05DPF15sn
XOiXd/bvO5W4qdAF8i0+BMU4BK5an9WKL+hfGFuwQM+WzZbMfF8ka6DZ5vjnSDnYq0QtLuu3HFcg
eU6GobAAz39OaTfFGVivAef8wkE0C623X23KRBkZfjdgnLHs8Vvurx0dJMBxL7RIPVrOg471ZKsu
1ORwUvHOSHHVuOGltVtqevsZhd6gtJAfgejzK7glV/eIwTQySBK4lUxDHfc6ogJTnNp99OXfOYt8
15WRs03GsNuvyJ3g9Jf/eXjmYJwFlKl/KJjnqRKfLH4y1fPvPCgXR86cP/ohLmzR88ctZtxbSPUr
2p9o5HQzcBNZStyYxjv92nLZzTFrwV+5wmnX4kZnc7eG/n7Re1p9XZaal98jpBqK+5AYdOiVZQvt
odRAWcyMxZKKtuaELs5iX4eQlpphyZ8y0bGny27Vo1uctkAA1B8ai/7hR8H1opDt9KchGnW+J9tE
aWjVTmTRI4GkTMJEmJPPOZGNZu4E60Vy+MKJnMH/aHi05PMg28pFka9zodr82fcJ+/m9PikO+MMB
iaO6nNJWjka3gGMMpKZJpaP2jEGZDwmll0kgsZSWojKOCKZtq/f7Ec+ONI4+qlCjk3kAr63G8xDW
fbBDBKmOGZUFKj2qjmyRuClTufMhUHPhqHQeG6HtrsK8tXkBrVbd6I2U9NJAPEvhz6c/qV91eA4z
T5LfG73EuwiOLBT+0/WEjUmM00ZG1bVHAIh2DKFCiGYkY9qMATz2mx/GvZMpxnDcaB8nLyCPtFlx
XNt7uyT9t0eK7s3IiVKPqrJ91XcWE5rVix165uIrJPQEZSZBBpWYbH0+JWpJ7cfMpDgppxCiTtlC
DNjcoOXHUb1o7hh9FOdpCG1jiuG1jvI0qQtTahXyO4j4yNE737gF3uw90NxcfkH0NSne7UbYJ/0T
dzxQS02hKdiYVBz8GgnuwwBhKmsn25CKMQzM14PerNe9wL8HX35jJU9L24lIGCihVWEBz21FxoUr
46o/Z2JexZDis1+DoIAHQoxcWdsA81wqMwMbuzQy0GGriNUIhJrB+l+Z1iNBWeZ2Po9bmyoPyxbq
bXsG4bmbj05VRcKZGu7G3vcs2Hjxw2bYgesmrHSzsw8Byxd04q0h84L2K7I8U4K7kbJkh0tiYz2x
ndqgq2t8nU7P4MAAHP9Wu4Q+E8zpLesYyQv8kOoR+KELdQACpuDGODyltms2dQe6HiQVI08rLDlS
kUbNrWV0EQw+FpsKRpr1Gy9Lq/YHKi7vOFqOn+SC78MZ/P6cYwvtXZpy1MZCvrriNkUUsmLwLALX
YP5j4rV8zYuciiGgQBnOuQU4YSh2NQV5a9DcykIqp6NAyFuG14BBhM2WM4KROGbBKHKnjOn3ZAhu
iyg6uZSec8GrIS9DzvFtPJwSjzxniRhZafHqbfoABQRrnB88VfAQBa9LwoI4CqVuhlLpi2kSBEZv
xn4KVxT5zULqN7PEnZyjZBm/vn6WwrE4r+vJJ0m82IU6liKe4dA8NR0lm3XfcZjbYpjO+QGTCZtb
DAo4Pr8D916jCnqbZbnU+iYGBdV41BQ/imGQb+VUqovOT0JlsqbB0DyfosIPRB3CEpuWrcm9T3Sx
gdiWGqm/0A/TuItbvWYhXzernVC0cSN+FhLKI4KOcGvJYqtnHBAh2GQT9J4j5PVTeXnZig56SbBZ
ymexXEMP/VzlqGo+xwv40aoYpplJY6cRs1m9i/mNP/FIyb0DSr3Z+aCXisMIEnpWBlp6u/9V/fl0
qklKQDxsTCy5cGP4eOXW3y0JgzJqb2L32JUQnW6wbH4JEwDMemTYOP4O06Uk/PoAvnhp9sW2AcEo
9nIj/yptaNBPOJIUHMGv8io4l0ztKlVRbdsezObu/2EniC5kNm3GXbud0FFwMxFn8Nqp+wgUqze2
WqbV2oia640G2zsj2ZY3w61NrJvSotgsbKwd85KQv8TPREcEDFaQUuDAf6BxT4/3NUuOZcb+rdnW
hNW4ovQ42itAqvd5In6L/XdEgJKbbhWyhsq+fR0RSAG7PoQXy8pDscWPwy2qfk7I6MWq3eknQ7mk
r5yxOBxGu1ulfHDEUAU3Pfb0g+dfq+hJNQiRUhAZcd7KMQn2t3edvmQZ7rPg9rrgPWhjZSuz6Cfc
fpg7D33qGgdAGsDUkNNH52i7SaAx4tJNQfLGPn1rPq0VCOceCoFbo6ajnX79gJQrhcBcP44uacLS
ZzMl/gbwVtDi50fAdwyjDNpzhIiv3p17A1AIq/2XH4IwhBYJM76YQDwc0fuz2vnwhva5nkBd2l0X
lfyYmUPvBYyXLCl1cctcG7yBDh0ZWpGOQlvJ8gmv66FRBAj8dzelf/YmlSzMXohenEmMxLQ0K8DZ
mW1iG1T8WiHndj+UFSpO3/MKoH4P8LMAH5hu7oODL8ph/fk+WqdqxyOEj/xSxWIBdCnarHSnKH5i
c/VRycW4R6rmpLRdJQCrttkrUjIYm41PGZzq1UjVgZ8f0otqV43x8eZC5mPh3UOqCx1UL9tqpc9Z
/jM7ufycN2h7AwNEuqWjEfSAO63VMvXIedZMsWXSDR9tl6nT0ECfM0mtfXfc9z9BUSKBGxN67EJP
/F+yfr502nbdYab8GIGf/wnfwRd4z2z7pYJrGhV75aEQlp3kttVhv2ymMJbLE8HijDCvuL4Oi4Pq
m+PBgRdDm/hDhN08nS/HaMee/MVrYlU8EBWOIoJwL4crJ3PXABcZoE9Xmjg3+Tzik2QzRg7MxvIY
1TJTAMUsqBnP8GLxsOQ2F0+mhneC7ufYh4woKRq+p3zoJMVc7GGd68tRCgMUr+Kn52cySEAiqpxV
+ZUhQd92jr+FsHX+ls59jjoXlBdnXz2Zc5rP3P9DYtOfgESmKFdIax8p2PGcbLogTMumr6XtX2uq
QLEp+a8mZB3RCZPl7CC0GtJi9PdOxRaz88WOtAsg5/wmQINje41kuVuYjF8ayTVegyx5V2BaKTxv
Fu1yw1HuHRNffSr3dl/I/zkzxfKxPJBSa0zjNHBYfMlG4uQo3LSyHn/9um1iywXIrN/ATijKxAIL
+NvVDRYGXLnPfEhFoLK5c/Gj1YAP5VTO91KEbJ9/vhqJbZ19WVYC8qmFb+SiAFvedl8701h3VL/C
XFOs5bCZUpAexFYw6CV+hKcYlNmaEsFUILXYwP/1raEMVHVsxCTvc1RuTxrSnW6Dw1j5Aruu1Je0
S7pc47bJV1nwTFaraYgWGViln8uSpkif4p/sPRjtXUaMNaeooG1UHCsGBVXHZ5QN5PRj0bUlozux
gQQ5Z9yDWVBe78cwwYnFvDzyFCJtAho3nkbW1zM50eUM/2yKABwipZWJAKYg05ComELZPdjcdG3U
JD6zpBBXDYeyhVa1p4URi+/Y92sptG/7fa6IILaOu8KeUmxlomfD2JKkMQcLvusxkl7CXgEZUTlS
yNC75/Usz3un4NjM2G9Dqv069nhZR13bw6m9p+WnbfjHLaU+0yT5wff+nFq9lgDs+dHiThnt2pv+
03TcoXYrRIDnRPfsKp4Wxidvgq4ICHLDMBfP9Hn00PI+aBMml0LvR0lwDPqiDBuVnQMBZ/xKFufg
6bugvYJO64RWIY2wxZGCESCr91ptKyX8D8fgU447P753TZH4tfz7y51UMp1lDT9zO0Dd4TmaALAn
as3vAemrktAUGd/QUmBLquA5hAYAhnLO/Ll+9HLG6iJYYzUmec+zMaHZsADTLl2MIk5gWsed1q1K
LGLFdT2soL/9tWiPjnm8+y1FE/LWHhvSCpwxkjxjxsZIbZ5VfAKKLpNkCKuM4JN8M902Q8KbPJC7
IE7Py0kl6bUWwClbCaDsRDhDX2+cgGt2qGVv5dKMB/c8TZNG0NqASN0WafztIRZYeLc/Du4a26U2
eB5xYLVPFSRvkR2opExpLsrwwJGnWugmam5NrBcFd1ai7EbYJYFAOdjZstgpFxzwMMFBy2MMWEjK
PAXqYd+pGRM6PkqxG7ST2VB4ZCEq73qj7BXuaOPbAmgHVvmbBOaq0ChjByYOLdPionxb4V2gATlu
fq+v5nH0pmEIukAkhWA3jkj1QiQ19NMnQTFIa4F4pyv+iw0vTxdowRDZoJvqd+vXShTYaH35Ce7U
mhXRzKV19rCAsQ5bXmfaeXHVNzrpdVc33ON8ErM3oZLCBLs517CBOMaMQNqWEU60F9EX/7Klcqko
v4fCiOWQEP2R0nVcDS287xM7XwqbtrbkGxKITV4VS4U8cI1TOvQMQDBlKZ3mENjkhw/HcgnzoIFX
mqTELTuL9eyslj79NLw7ghAsL0CJDeoTf2OVWCwasl7zbz0ykylrHazDNkwI5Km9ku3j1c2xjrx3
DXXHAf5Fodzf0kfnsLjZxxIrtpFiUm+tOJVghpes80iqAYooJAsfLLHcIz5+npaHmbfdro+vYpdS
ctduixEFidjv/Wge0NYxSSTF7C8xWMfLiAGrDsNS34jc5g0ZCxiGyKs1hABOEZfVc6BMNhcgwk43
7AmME8HCJ1ja/LMzOx2u8Eo+XK1yBg6l5SU0YImjMlMbFrGPkR2WAy+kQDfaSIMiJxi2nKn2gP74
6yOubdFn3Q7wbJ0CtiN2LODJbig+CcgAOhzSYLW1P4nS0si5YgYFK4XRbQeNLxrsXmCHFF89nJQe
UvL4QhVRNlNAusiFcVqj4/q7yaEuXZab8PGrs7SdtR9GsqpdMtTvsnvPaZHJcVSwPGGcm5kGZ4M/
jy4zodU2mZ4ekaahQVlBrE/STjKU00Eatz6Af2Wm/9Nm6oUCUcs50LVmirXtZ7RzZDTzfThsD3oL
tBHtJl5J5NOU5njmTfS+Ee6gYMhonLkT2TWfianEuFGz3x7Hawe7Sryyf5FITYEU5wWZpQ/HfaqQ
7BExO367R1NTr6mym/0SYWQpAM0RqEv/b/qUz8w8TNMSUaN6yJP+wtkaB8YRm6qa3P63p8uRVFmb
WehAUaduLXdxSlLXY+lqUCZV+oelfYkVGn02nn6QuRW/fqff128u1aoZ+7O/eb0tTMFLmcXD3sD/
ypipXbczkggdnE4vNL194zYlwrpEqNepSbptN7t3HSu0XwxbPrcFhtutE9eA46ff9+QZlSAQF0tR
tIoNaQLAtZpC5+/6gTQZNU7P2YU/M11K4wBccYMYET3u77/80Z7xMawcu8wX4JSSHoAfR4yz3SNT
lo30vZ8d4yQr6gPuL7tHJrmSB8sxIR/qF0cU11R4G48JHflF/sREuSokhVb5S1pZAmMHRhDK/CpV
efEJRZZFOobqlwuhL/TS4Ss9Cjf3EHYCBTyfJtrk3zENda0gfuxoRc69dqLAqRlKLyHcTb1eJJnv
e/hO+Ax/cDmS6GKx53fUA01gPCPHJG6suiCT0taaX98MUhz/lDMLZDN963MWS84by/FpxVKee4Eb
k1Jef7I6UjRiYPp03/omH9qGqM2PGYKPWp+Rjq2tBQCcWB6iKt2vIFGDHA7xFCJzpGiASIECd1kA
j/C5nTTIdUwaPqpc3MviKvVQenF3eBw8PAvyKOyxTd+VnnBIT0FNXkeBzE6O56XUi7/NGNiK+RVW
Ejf9JXugk8WS1Oz5cVOhK+ccYLf/d2rbNvPtNKwOq8EtIVSQGhg7O7LQ9BCtuKjZENMVRu/wpMxT
Mhwd0HqmE5PA771aV8Gm2fxs1jkWMlquh6aYaoVsNQnzKGpLmj6C3As8Dw2oaQLEsiXAn8JhZyHZ
xPmSB5gUuEvh4YR9yMt0l4D0lAxejwDNRN9hI7E09EZN9rfRnqwDfDFwxgl3Dzi+Aag/BIThQB5+
rnIuPp0yeA7b31t578tqTOX8bKqp0f+s0iaLpW0vXxzZ7NoCv72+kmP8goh9BHhTK0NfKRiSPHjq
Aj6AasfbmkULsX4ha2XuyKMlW+P6OR9Q8KUDiAE6PJcorvhfAsDGEAhLFasVxNoOjYm1egdDZjAB
vpkl29O/xWcuuCQyX3U8mhtn3NTyCd87EdnEXtaXOrb40V/f8F1SiLKApKrtbEeytcXyeUCibwNB
uy/6ZjsqDR10oxKolpQm8V3jLfvm3gT0tkK1vJgXRhvIdf70nvdajyih7cQ/URqe6B/lvRnFEWVZ
P7laJVpWepnH/CkHpGAyKS1v1+w/ZJGwEMvbowpyEIElLeA6MVFIWlQ/8kR8uqFDsI9CqILfGIq4
upMyHAI6ItcnkNcUM3JXgF1aQohXheZjTZ4c2qhel0V4X6cmXMmbU2VAwmhCyESKpOqS9pZiXQWp
Owj0ou6tCF/OUNShOlwr4rPHO2DgLqLjsS8+e7prDSrVrGBXhMt+j23dcYFieZi02m2uKc5S+IFL
UJJY0vtiN/V3WNs7layZLSxMWaY0PYFWmluzVlDKX62RhiOOYAFEV3OVeLswORoKTbN8pKJq7jEE
gkSw98aWNj4y6JP1z0hcUADjyJPjITANr8cH7loGHVal7lCLWU9i/spcRjkxsEeydxRxBrTa5MR7
bF+CbtSGM+l0W+xJfPNZis2kMZBWszZVoU2YbsINcXnX/cpSvpbYZkPFDri2rT0TB7OdBvygjZMB
0BStzsQhx0Cxa43qUPcSWyOSX1cExNXmBC8tfiIe6F1biEm5UUgmC4WubZ2u/tG/luiaMjBvogI2
NJye8RH8ton8xmG6wo5J7Ft4W1Ma/m/kKYZfiwf4x7kuq1A2lJA1Y2ngNUiN+voA94cIbQAzDZpV
FGPSvK50nStyKKKEPglDTiGhhag6B4QS/d9ClX7wmfVa9D0ObyOS7EREKjcVNDzPY0p6/WiQ6uk9
bfU44JtFq6AweltWrjCo5+TfhZOq/t2ArLzXDh9TOWDvZYPZ1myPNfy1C9GnEqdE1xRrhGq0OhNp
4r3ajsPr0z96uIKr/yZOBLU4K+CKPxqkNoZjbVYlshH5uLCOhPittDsJE28c7mUBEmPuK4AS1Jmf
T8+NomMv/u7OzPpVBkg4yqhZn0rmestAg3j/L4pMOoXY68l1ZcoYXhm0/WaFodtDw2o+6ZYdb7Lc
2VWgcdj+uJD5rBCXdzpd7jlJG+Lk76AZ7Z2NpP/ELETHrl5qXSjpdZWqbiE0VqPgGTF0rE4VSo4J
UQJXEEV3TPOC/6PE0BnGlp03vVJUAh2rSgqrAAlzTg2NSiFK0yAxRreRtBU0ULaQeKookioX4mmU
9SgHoWGROmHvIgT7otTF38m9WBWUeGEgZLIEHZGisj/TrjLqJMVWXnRcZLMcB835wWfxxeGmvnQV
7HHZyLb8Xfm9TiBpK9W0bc1n7PqqahrSWnkErJmJsUqwGSfLtkqQqoEJn/vyK0yNGW459DpU8Q60
ur9cGlg4tv4XcmxidncUAqBD83RvqgcYvl3+50QrqtPwhRLulPjuDunON5lMkC/QqTTnb9Ajrm8Q
+KfgRTt+tefKYsSf9inmA2c0F250IiLV4uwt2iH5Y3MN8fV5MPYAbglz/H3SvyHPfL5yMD9eoMz+
ICeCR79O9WGH9yFpuGwN3yRg/lMwsFq/bV1npQ6BzoH+pT9XMLaJHxi4HemUuS4GXk6OdtZF/1Dn
Na46Rd3lucosk/QEIwUGi+r5XMvdka1M1Swv5z21F61bgmFTclyXqqWAeGwRoB6Er+clGmw4q0QG
8B4zX/jG/y5BhZOtRh4iYlX8yrG/MsEuMohizaVLRKSW2K2X6fIPAsuA88fb8K0pWi/NUc/jaIHf
k3Sm46QqBwH8tcRr2zhQxfWQUuSpGygqp/5sJmRwW3CrIQC33SGMQkyNrdQiejIVh7XYUYS5vrJq
JkU9bN6uZMEHb/fUS7eva/SUP46OcFWEACZvADDk2WEV62DLof1GAQ3eASP3Dtxk05GZ1zjj6QNH
51D47LHvWXc9CU7w9wwZc/H1N7maTuxBvUg9gL3m9/EZJY3vLjsWPm40C28KPRMphnKfrqoAmPEa
9JxuuYSToqdaETcac60+tLZeCJQpF6FNEnS/Ec4wPZP9yGW7It1ZXyQzigFrVSD6929dMsTkS/C2
yVzKZMCknvVTn9UzV170/4fghOlRJTyt1wKHKi5OwmpigAexiFoQTVmH+t8xBhfmrfDGrfwGTMAh
jtcAqjlvg0EjvlijmK1wq31rBrq+rrO9bmBakF3JfGBnR3s9vo8lzpET3IXnHsuigZr3NuRrabRG
SGPsmor/uGzx1q9zHZHSngvhrbXGye7FM9Rog4J6uzviAmmAOzcUkVF1Ks6YgbcBE2mPLyIaHpPO
0JRzrrmoHJnyGsypHOTN+Ajl4B3RDFM6k6mG2nK89KaS+1VJZWhZlChqRVP7NNvh+bIgAi47K2Yw
vUyj5aGGnnlVpJT69l4hhapplIQQ9SPi5lmMrKJI3x9xmKQ+i8w9MFnd+3prTqy4zJBXp7BsNgh1
vYJ7Yr+0zsg2WvxjYSRW3xE/W7PzxDe0WyKJwxZAotLdSbf6zTqbIUN2cG8WVzi8n/wmmuj2Y0Co
Gj5HBrKvbI2DkFbSV25FGbUa/Z/yJXa8zMZwm//bDl1faxxOimEjbHGGh4lWTJ70ZrGfd+GtGDqY
sd1VqaBiy0+gQregAGemmfq8ZLYwRPrJ9yhmxp3qfofRId7YtBtPTxHIEh+RN5JSTcaMyaiVFMjZ
yNhKOqK9olSvMhVY9jm1s6qZo53CNB5VZVJEHvereD8B9eHT3j6sgfKqsr0RLLtxdtXuAtQSQwNw
5pZgPnhVResBxbKoPS6Pdxl3VWvQRsUVFDeFRfzpfBSysKKH3+sAq2WX1uK3J6XlyfNNcWK2a905
2rl2MLMYboD1tpp40G3dJqRhxkGIfzdAxvr3rCPWa9Mgv1VeZhdSmOh5IB8LM0IdeLObrBi8jtjD
QvkBXZ92slAJZkGpL+ocHZgKnFnE1dvvS49Vup96rEy7Qaaa2/tRFLJHziYmWi2CrW9TDMHuM09O
NShiwZ7LJQ5XlBxZRLH2CZmZeGyqguj8clcqAlPqDvhn4jEVNb1DfKL/O3MmXb1kIIF1SjcFnjPk
LSkY0KeP2bUgACpLHwzaGW5FBx141cEfXKzSGWvCGWcWwCdJLXR87VcWdSMtFqTjy2k9E/VoibQT
f8fFISNTPvPhpqci5OtOF5mM++5KrRahuDrD7zQBMzjyRQOD0vdwbURKaOYZEmzIsy+JVbfZZr2o
JFYV15hDrQr8Cn6FwtjrQNAPrf82X6IwaGX9D/CQXQl1sjPRDs6Xh+AHkAcFMdaC0qyiUp+6sQAa
aYS4c1m59x98mVxFOYgWSg8NE6f8Iy+vE9B/M7dH2LQExoC5QrBIx1fjCx6Ss/bzG8nLLUFoA+0n
GLlYm2uVdW4CxhyAb0oRiQCWjnaeHTvgF5CAEJNRcfa3SmYhL4PYF1TGnGId2LeE4vozP+pjQbgJ
DBhwbO+netx/GstClK9kWO0kD7IHSZUZvrMelVEYm8+kB4R6Sps1Ho5c2/V/z8/c0irvBPFAElgc
luqmoIr1/ToRqUu1P86a7PbvNc+KSH/acVi5va2guFrF3GMlVEYTczEaveKqNcJ3F+Dm99g1OAsU
1sXaGJDaWeBl81HaTF92joNSCzIFu3nfgN7nJ3pOvRiNIyd6eOVjoapk7t4GMqqsC/7Nk53TZyaY
rQXTaQgb7YMJj7MoiXbfaeKAqSfMXzFM+ulZryWpGuF39ow0QIaugmJffeBEGBehTFhPVecHOtqZ
witvGQBpOfmmtO9qdC4XSdSsujg1mPuDpJ9RXUeZ030+MWLtp134g2a2regwHRGMr6zxn2GPik39
5kJkS7DJnLuMdyERNsEiXjLe3qd0Q56Ob6omuDeivBhlXUnasO7T4JeaBA4fJde11zUhYtowK5b3
pmeUW76bZRfmGoN6XdRZAeFFsi5ChiXC6KyJXLBWo7ZuRZPngfhLRVy6Il9nqNpOJZ4orgjepLfb
mG3eJRAsuxm+VPYHcMi0MgngfIRHXx5dSe+j4aPDUxXz4cpaN62/s6iXh6S9OjsMaL2RyALctAdL
m429XLOwIPoRi6k7R4bcTyK4n6a3oG8U6PowM0NAGB32faeNSIwy+DAkzV5q/mVdpRbzLrTaVFBb
U+ULUhxBNu7FnaL7qUVpsOOgGrGJ8SX0U+yLOun2TP/BYEaYOp1Mhz+v5MSQBownngVSY5w7pvbi
ayavQ5k0lj+KiXBZ41/J+VYsbkRa/4DHiyZQvnW0Ipbf9Bz1+X6Y2x5gMEZgFjPy/L77opXuxKQd
aQBOL/x04eZXTJdu5YyZB90swEx7SyvvWmgRWG4RbmKip/FPh1+8J8+BVEnRNXvB+ZziZ9wrjDcK
Okp8vLJRqE9lgB9Jlpm2EQvmFBT41w2crlb0J1QVLy9IbsBMNPGm0cQg4vKIupnYQDmjRQn3sVo+
MjESTnIgoQzsHwUkSCp4JV7ZiabucQZVZohSiccW2ZACLJHr3WU2xFcU8Vq5yUJQCO6Bq4p9Wk5p
Ze7+UmrT4X+p8lY4at0g9U9IFmRAeEYxTaAy9jwd/0fvNZMRtqN7tMYIrOMP3lVPiBr86Kjk7Z0J
NLSM5duXEOF0CCEeRmMo49cdtmaoekTpRv0RsgixIwoEU5h3hLzG6uEmiLbnKvXwdiLNKkdpFpzf
wa2zgeT6N9EuK5CpgQrDp7jdxJXnqvQAwEyoQA41vUX5sRn30Wo0ogjeXc1LqUwseSZo8bRyrBAZ
AON0V8j+d+VeaItLhEwe58o1SUGavUgHmMA2P8y7XUlhMDzMD1vQ96m0+CCbglzG+lQ7Md2LmKXc
xE+iBlDxruf2N+0HB8PxkcD4zslkhcloEV7mD7q5O5HH5IIfIOkvjKKJDifef6tIRf7zY2rRSGGu
ZS6kv7Wy3+2WC5dIz4UiOQohghQWb85BDOZAkO9iAXGg0zbxg1wfRpuirNZvWN8iEwRmjtyQxTa4
hSQd3Ibv+voSBIuDZ4KKxlKFv78boTgUA7+Wblr3EwA/aQ0+5h3o7a3gBjCPqUuuxaFaxOviRlG3
u6E6lfmcWa2kAcLxqlWY4xY3pSYX/ZsCDCdWKT4MlaMk90+Dp4MRQTaEcoMrskDImn0BR6Cfyluh
dTfOCJ48sTzvLur9N+B8Eyb6TrYMW3s0h8dh9xGV2Okzz4TPvtVPsCeaW22Edfr3TFTpA6ZcslTv
IQmall368TUqO9QpB0pn7fSo3coK6K7fxCXApe1CUV82drP7bCNT1Hh8OJZhgCElmFiupNgHuinB
9xNO7CRU7T70+qKwe05KaXExzOW5q5vrV2cOxd3ZgptObbTKxb1FRGaKBZxV7c6L3XoFQ41WwNAn
a1RFvBIkOYxMdYN3mO8p+46VwuOQU3amdF+RGEO5elXTWNxs78heHKbcXSRVYeshC5TsjSISWORs
13Nrw6JkNKn4+5jN0SYpcQudrVNRvCw/z9h69OP7woL4qbf0rBIDLSRtg26hbtee/1C1Y0b6P5BG
PZI4TMj4cFij1kiguHI1/RCETsBmpD8lUY/T1VkEtMn6EUOk9CWV4azNtfUrEX9Hz3YxCq52LR5j
JWkevhjYo8cOMUScy0baLg1GZ9az7NbP7lL6p7gKZBjMuWLwapW3XCpFjiql/O0/X+82Ozzre++u
ugZPvnBvuz4evTlVWtz4jen42Y09nVZaXFSDBaakPlw+U9THs273ful1sWxv5WfUIl2i8oChL59X
/9uVH4Tke8jrd4aS/lOUC/Jf1zmljwrYryjGBRX4mueFC+/6NxzmqaMdpijVuIBkVy175AK0q8KC
mzOijSC+3btmEaqaWffxV8iswXfTB8QQmreG76hMk4/Sk0/jbnWVnl9D4OMM6vcPd2MPDrYwm5dn
+gM1cG3pLb3F6BSEq+1U8vsVs3Kag7oeYCzu78Mk5XaabxnIZnzQsAaDRIgsoqkmBk+4BBgDPhOw
vtTlrEum9ryY3vB6TR80O6q2fpR/lLknI0escWom+unNpdwx575Bwe7W0VTbfenSu3w8pnc2XqVK
+6n2HvRaVDsJLf8TOwm2pbf5KLC3svdqUMA6SOUx1Mfu7fst2/YGWl+bbrWoqWfHms8KgCiflwda
RMlgYG57wBpTZ/UWQHz1jA8QZjFRC+I8z/Mh3/vCzx+EfNASeMOOcIP+NJvizc/b/phHDm9hbX9l
GVxVi6WoZMlzkxWs1OZXpykm9RgofZQ49L0vxpw5sZ2vkzokcfn2PSzLQDX/ICE3QSxW/VGEsWpR
QlKWckS/zYbl6S9v0TDSRO9QlIQUX1kDrdRavcV+zREF9NM1geiowfb0wpAZS2tQVSUt5JTMta6F
x6HRM1kkHUjiOrAhfZM+es6mG0y1Saavjw6LVk54GgCZf8DamjJaHImf0HHcj0Lgjydpn+jSUBuH
9hbhxM0HOATvMAKdN14zFO8tOk/uKiRgIY3X8Kdoc9tejVTpk0S7uedxLiVUc+JoSrl1vD9YzaMA
Hij7+O/996yjfOgAvs9eSWXr3ThZQ/xrXh2WKNrDCSrLS1J8HD0GnrtHaT+dQXWBZHg32YHZV1Wy
+SPQNxyx/gHXVdCWYvGLzVW0UmoCV+piyZTIFIwVupwpcYYLO14R4AZUHnPNBIg/pq3ijNqVWhrO
TiCC5ZSg3Cl1YxZPngH1GjB54+ILDIZ+JSvSZumXZK75+OoLKzt+H9xwzVt1k7sjt50NR/dZXw6R
LX+qbkzVqqR8+I15+UDQ09k7wDpJGZGf5LNe4LE7/b8G/CnIqU/IIgPloz+bFJn78kahjMtzfNRo
rVahtKotTVIHFLUdat0i2JThZhF/9FGy5J6kU/O0dTpEupOeNBKJY+Dko1DRItIxdAtu4dxQtue7
WPqJERbspLARFHckpxHe0CxIK7qNJgUCRJHrhvE5R/hdPIMxg3G+zG+JnjUqoFaHlxRRarX5t4IH
BfJ131141/6OtIc8wTNcX2uv1jIXjVz0BcTVHWfyJHUQsY7K3Wd88+BHsZWACqnKG/K21QV7jq+M
ftxaMX1qCmVkDAv2/UAZYKkUGvm8hZ3zYXiVClKa1MGwDNEU0tHC0qazBg+amd04YoU77kFW+a3D
bNigLWAXcScQo6/X5IIkR/DTYT9oIQXPkSuUs8m6i2kQ+WFS7SW3/SLNPHyaDA6Ijffd2utfObdA
jmdbs0L2KW1JvUAcvOMJCLUQVFK3yfS99qZ/9cf+wUXPjkRz6kVVqGZPTU+E6gD7mBPSx5frk8bf
oIBlYp1bK7UFo9avPyeCHHMET95pYMLbL8v7ylxdYkTbnYpHZOHkpKhgf1q+gLGIMAIrzVn6qxnT
1RA0NOvFZPRXmXnY77UWQFSlpomcrxSp0/YiAmws9xLILRb0PrBEw/U/tD6/0Zrn02vNb55zxYgY
7SU0sNWcuUNpz0+044E6MhnBaYu7b7GTNdixjQ1Tbukb5T5Q8tncfFEKxGVETHFRRwo/2CnOTGXG
HScqQ0ytH8c+Utdn7Qrhfd5Gm1H9FefCaHTO8NaTyzPrrN+sW8IDEmBXmJaGPvh1N8s0pTJpJ7yn
ZFXTBoWLuP4CxuuqhUY7eVCJZqsSdezf3hYfnKYvuE1kp0Nf7aWnBpr3uCmnPfXYTRsDgzgafWgV
m9SxSnscB7Tc6HmK0iHTtR5QKC9zWnu8uK9IxTgT27dz7dvoeQAEHJPBDbBpyR4Hy1/jyKGqWSi4
RSJEd4pBba6Xdf7Fx4mT7O7bNEduaPz2cOhIw3fh+SKpRqtlpm5hmu5Cgx4IsTZ7nC3eiYBZyCc5
WAnSIPh2+LdD0xUQOhpxyN5AiGv2hHQjDSg9hwivdR53CCqJmE53yR6URb0AqmwG4VThvpJsBWta
mGhjupQ5bYTY6cdB7Ib5baPdiFs7duxI9q6o8zzlQDsj+YkRbKQWOazfcGSG+8J70ALKg5WZkn4/
l1AZmtdzWFurEacEZO4IBV3ID4zKV9J0J1hbCPZTGguZrX3h7MSS+9S0hRAYlhvdUe1FE5KIrKLk
q6PC7qRZCrDBqYy3f91bbhdr+g5A8wBceJ3sC5dpDnge9/Pb+bdeBz2JeQ8q7Vmx6PFT51jcuA6W
oVqBE9vl9K92iSzDPvRn7X6qMdNwXNilJBAciUsJCCH9J2wFyU8O5xmEMq1flCIfhRj3xJbZh2Uw
KUdgkXAzB1RerEjxASu09Cx0i9J80/F/4eht2t0RDtn2EXQpPM8LCqG3Z+ZeuTqUCY83nJeZVREX
Olk41/QxmfqIV+Be1A+lhl2rXWmWlxOVS52RkzKiKiKgkWlx6L0X5+uGVR3kieWGX64xMMR+VheX
QIo3nFFTQwRdFtrcP2R64OOub9eYGP6q4Q1Mzab1bC5uyq1yuWomFMxASwoHka1T4GTTWu3dgXxl
Jyh09b63GUGvBnJzilIPef0enCOjpC80JbG9iUADVSTOcfs0pdPRLsS0LET3sCuZhEj2hS33tzAv
z3w11TsDG9EGN2GCoduYqy6fC7482TUu2QmLX568Rq/oynIK9IDjXm1r8u4F+rgt0gb/N3gdB52a
JoO7B2sTsTeHuXAkS9OLd8LZuLZp6EN+VIFmiDAFU6nG/lqaZ+unx1joAP3QTGURcqGlBPQ86Ujk
LKL+y73cPcNCSt4QBolk3KXI1cbY+bVjIiOWUkwG5QWTmej+DWQxvdkgfBy5IOSyJvHKLlEC4fgf
AntLn7MRX+nTyOxLOQd3t+LApZUflwIUtfxU+a2EoBvv+1o67ijRvfjU5fOrTGh1A4Syp3Z9v8I7
S/M0NrxSBFqWBJx3xU8LA7GWNKX5d8u9krR/p3Bg3pQGiMYkuzHAvu3KPx0M7R6XI+lhijy2P5C9
aoQcL+vxw/jQFdDEcc6XSpDJgnYnr9yQ8g/zguJb4YmBZHjQDzEGYbhcBFaL6HHKm9ocodDT8lLq
ck+247hbbYQho62gMimB8xMgkH+MxZJWj8lqP8MU9CkovuV/Yo3V++RdKdX58B32OMFJLgg1m/bp
DHw1jUoX7waPrVeEvl8cXARz7gEsPoTY+V+RywaUaAEhdOKPsv/nQXgmy1yghL3W+yBi9VHu3vR8
JwP8H4Hg2U+I+sSSK/nRNThpk68/iGOMGAsmX2105HjrDe5mnL8RfSLKlh3AfdM5//ki9CNcTEOc
+NKFMe2TmpEJIRqmsxiYjOYYZ/h1I3USnQILuawv0Gxi+b9deVTALEtFtS5virOBq9PN2G4bl6ym
nAN4TAPxbzO74OT3mkccnigjnITL1GrQCE5aV8U6BGUrgPLpMK3zqy7EzX5OoZOhETv9rGphBGfe
tCq2Io82E2oCGc/tMaZief1kFt3CsweDKtKA9vcZQV8lakc2Sew9Si3RdQcVGrpfFCw/17JsaOO6
vno9DGYdR6z7T70Pg2r01Hf0Qj7ffYxZiMfBain7BZwGXj52XdtMW+vB97JiXLzfkL2+MhLrRNyT
322Pz68cy1uzB7mNSKBaNJFr5QuINn0pyacxj53v8LnG9r3OUloqG4toruF/BKiU5zhf2UNEMIV7
2asXM0D6oepCIxpSlxfOpueYdzptzMoN36eFrCGaErG3uH5F9lSwbwAFjgOaASs+MKElviTAwfYm
Fn9CLBWtR9dbl2XVB3jbWsWY9RZmVUJ5LtoH78n2SUOjKPrgqbzNdF9hClsWoT841wh7UgH7Lv7L
MyljZHHy5w76ooPuDEybdkICUOnBlBOeMyPx/15913nd5qqDR8Oq0ZnYJFSWcKM28js4sVypcTcq
Om1JMavKX/Nky6HXM2CAuQp+aS0cNMfe0tN7K8yqNu3asx1PtJ5wY+0kVXP7QOn3icInI+imCISF
bIrKqK0ALQuMu9PyvbFv7rrRpNRR0/HLQjm4qWJjYxrSWLsJmEgZHsJc04kM/bXGjwKhofbFceOh
dm7WQZ19VfTnK1XH2i9FqftQlcGDEKvNgEpHDPfz5j7876AcyS7pfrnGKtc69dZJXKnrextCu/7B
rI96/JQrwd3zxHi9EeFJKyxeulAB4ppRXxt6/AMu7w6gub1teG2QRCovQ8YFLpElsrLs8/xa0qsn
PXXSit9mSM1PPkUpLjkgHYEoBqnaXjrnkvHlsb2UT4d095XNEgFMsCS5cSUlDC8XqqRub5PwXJrc
pfVpWwDi5c0XnkjmJXYIYrvHpS+zEUIVEi5stnF9iZI1gB2a+BNnon6GHVKDhEH31ACyQezQBKts
j/4RiO83yVEz0RYAgy3Mb1a+vgmpF2JHvDpMqsecnXVzyE1A8d/+5hpFCG/+NWG5cQqE4GSQssbo
ylcgvVJK9MIGk7nGK+bJ8m8MCi+uGa16zqDCzFonZR2fh7RcEwZr/plzEItbBPpOIfFzJopP84iL
WdXWo3oKyC2J/v/CJZ8V9zVC1q9RHmNxqU3ntpU8Yd/eSWBTAI05OkLKEXLapNpqrdtX1G5+IIXv
h853CLSWE16oS6UhQAr/uTcrZnAUloFzQ5Bu8Mbvlr1FWybobSVpX6frWRs6KYrpnMRClDTU2v2K
1blmhlNRTGTBj57zP1DyNdz5FarynaKgUtWCu9M6mQzUQXYQGAiqII6CxUMTgITfMBB9Lg7NC4jj
wk6xQFYEqNnjVe+aJBWCwm+ExTu1Mwbq9zeZP0iHgjWDjjo8vsy1biidYEKjt3cGMskOfrTTqnEM
UuE4zMlmmXi+ghWSzR6BMJ654gwbVL5cRh77P1/PcBU0ONqb7LjYt3qgqzEyg3+AwowFE6NQVN/M
Jfm+M1yaU+jAgV+r0HfS1FeK8mWRk/zpfCr8ACHfZ83SZflJ3rZt6FRqZ+Deaia5u66Ms/15wji6
Rf7wZUrnIEl04IvMsrhHl7/PJSTeel65rAy3ErooUAgeMrHT2bjXvj9Z3JlR7OtbJnNjAUm9C03f
qUNwVS3XkcpFtUeI4f+/CsAk/lkDxFMRhNO9XIhQ2hxYh93tV85osNPW4xPIrowYerBgisxFeYC3
gDFSIbi+sfwUNMAK0pxnNyo8gZv0X9LuynAIxkel0C3y/W/JJ6j0xanN2H5dC6EVzP1WTDBsc5cm
mmp3I2sw7WIlWq8hvd5rJo9JjKM5uROuizo78BOoK+AyU/foTKGKwqohQ5hDyzLmmpyflJGdYrym
rGahG/MBvy2T55mI7DJkX8YWd6OolwOOvj+s5ATpaHOHWxh++V0zTsyRnbrw22wYdHkJDyo/e1eK
BSbB1K2CEO9T5SlhXUJRh/Hf1ndHkmd/zpmm7ohW+q3WS5EN4OVyDIOHRB7SJL7V2hnQKh92WROR
wLtQoDdmMaWG/tX7q5CzaO274XS0TODWLzES/h0OZDDOErXyuqCuH/ubyWKIyhZuTY1VEY+Frmpt
O6KreydeLw6wTiq7K8cSimVMChdxDmC6R4Wnflf8BREO38z917PbLS2NwYGvaBg9pwbrxTokgiIU
VqgTcauNF3w9He0O5wiWvdl7nHCU0pdNgBP0cYCIJPBBN72hvX0RmjLm157Azp7XasNgwkAvavyN
ul1rrnnbUl4bJKrl30S38bvI8n8tRo1pdJNLy3KaAJ1TErO4LlMq/A/2KGUKsDPBeGtmmobugXcO
wDRxgaa98MkM3MEVZfwCRWvj+0QMPQ8OXj7o2mZQrCb/alN/uwp0vaVEbkLkzBi0HWmOOBqd2mM3
gYVWx0RoclQDf0b5EvYLEzLD5F1GNQlSTxdJjOEecPfoH7qM7GY33nloLHqcu2znnc1mPF2eHE83
fjx3dXHseb0zFgaaPwVl9wIbfFF6WtZ2Ks5w5ZVTSAfxCk0wvN4n+8FUducE75XxQ2+EoaM9zpDP
7nAUQdPOqaO3nUKDLGF4w9vjqcavygktT3AB7cUZik+6F4wCLCKf0g7ieaoUxhF7JdSF7Qr+I7cL
h8IXOgDhj4p9QNJ0c9Z5Er9TBNUZ9QTIeBqdc2t8ryvXr/XoDrS8Tzji9aF3nl7Ff0E92ydBKTbs
E1PO45juj2l8uKets9KpbLR9eypw/qKHR4ZceNZ49usNq3vaLyfMNfAnC7/7fBnPvCqadxe8MBDh
oOjvpsn4a/9EDqKJHA0e+G0xNkOOtfQWiukOOUe3Gb+Qn4579364ohg0ow4kdg0UWwLeZjPrrrlB
smUC7LnC+05vfzu6+LkQ6e9M0M9Q4B6ZuiZFEEzETHpnCrymf2c96Ze8to9ts8CEGo8nCp8c+u61
5A6KKmTLXPpOc768CJt6vcKojssm8hHSvthv7eReNI4iswBBiuuCz3zreinRIX7D6YwhNgQH+HTB
FYh3wC/RuoomcOWYSzIi3xwX6UCr/DumzIF4z2Mf9JMxS/UxY+Ie5+o/Gb0JQCNpxRb5XQLvmHJF
pazhyZhKc+VWTaCljS5PePxYWwMK07OwMbnmItno540dRU5dnlH4NwWxggqCA54RxLl1d+Wcomlp
OJYWwf69B1Jd1CamDPRflmST63aQHhAk3SW8pAqAM+3LQig8utFZGz3bY5h5mARMBPOww0KH9UBq
1zH4bN+Yh01xHfsB1TjIAjyr0hMcsMHYRtxsLXc6UX+dnUSO60RqSPdBLh89WGwI1YfakDKGzMJS
hUjuA0ujgDvIjbapb86Qg1PwLvEUJZ95eTEiU2+VNcGIpAlP5ANIkSNBejQob88Ap4IFb/zhGnd1
YFNVEg00UPaooRUjKOwgYeQ6v3xEQ4+jZ6Qv9fv9dlLFwB5WUrUO0y832yeLcgcE9q6EdQL+lhqg
zHY+qU7InCkk8wHDsaE+XdTw0ktk5KL2ltWW/F4lPQD1paFNvWaOb/PYc9EZhrYA3PdGG3euxCBx
edacANxCBXmINLA2aFRa5gnkA4lQNhXxeZ2svBO9IfrjTYOfeZ124l4ggacbkri02tpjpCgDr7fE
ICJWT94rIOANwoH6bgnibt2W+KucTERoPrZXN54Tiroev5dqugkPfyewGkFh68aj8g+goCEOCtiF
9lQVaxpMB9R7y2UE2WDbujrRHWsDfoDtYwsf/jm+graw+XyjjpBjrUSW01xSLzLnSg4IH25zhrPt
gSNCJPXbwSHSmLCf8QS3xl3MlbLwJVg1DeW13rJUnsh1BXCQG8IyHM5y4wh9zSZatvsWe/24TOJ+
kTUpZ2gfSM1dRALnnOrAWZc3rhRLtaG/wNvbhf28eh8TpOkMdKr3cbzjcouVdpYgQdnrNEK3FMEc
CRMGfb5SV3ebWL1xqr2evxdodKRU6eXeJkMt8cHug/UR2at9sx5R5tPtUHlaqeb0TOXPzGSPMJc5
eu9SN0vDtXEMW/0GddJDPk9hS+Oq/IaMJBAIp6h60CrTgb8M2enIufneYlrbWfRjKWRF6OqejpRq
8mz3UO0NGO/pLOVo1E2MlV75o7V8rpCnxc+OGwgkQuEozVRGbekRF8X8+Xmo88VltLHb6llyYUAX
wnlYjadecyBMi1ZfWx9idpNE0DVEzgO4KuayT/zoCQOCdlqw5NUl31ZB4QUNu1Pxfkd2pX9lKcvT
VsvGbXm4Sj9hSs1n+qWDuBmzVcrPuJdkklDmyFmwoxULJUY8upPFaYt+y7rJOhwXEF/dK0RKfhQR
lz4m65wfbGhqA1cAGCBmIrjQyr6KI9cQeLJxAKof57d/HyOpivArLO+MUzwQs71QgUw7YHrYch7o
5Oz1NWp+yN/u9gKRpEVlbQSE7xdexXcf4NyxQg2Mjf4L1pzgZZfNWVZchnufqG0rdX+JO/ryDSTP
5RUAiEJ90HoZK3x/kPemZ6Hh1tKNZv9IMb7vavmXolKKMFwGROkj7MHSTMyjpmNjZF/dvf7NtRen
BHgZWTxrUZ4z+3TEUmEIx5ZFOyCdYNGD8xbdau22vnQWB8Di16Pve6ajFa9pXF9XdesE1OKY/Eh3
4m5MrgPuMhABsl9kSF2Lma5I8dsNtrIqJpSh1RGP0TOzdDpjqxzGd8BxDBF8BilMEHoonJ6qGyzO
8AiXyKcMqOiX5GdblOfp9z9GjryrcD9F50860hHbc2rBi6uQRgL5s1rBIu8C37mGDbem/7o7jyKV
v/SwcX8E76CbaDQgAO1kGZUnH/gTCjydM2flvPNlpQzwjGrjxBqEoMeqY7Rc3Sparz2UFDWwDFQc
PCAyaxwNkTCHZQS7tAFyMRiR0sZ/lXRpbJPSTKl/mbt7ZlLMM3np5wQmERkY10CIi9Y7WEeiGmml
ustgwZ5Z8+VgKciRX5gYnl7ZsTZeWitSb5PzMDIzX81/bGn9kfEpRJys2SGi18/hpgvyC2aSqmfR
isKKWvbhyOVTMQt4/29xJPEuIk2PxJYK7to7leoPVxXfG1xH/996PZp8/NqjNmC55/4t9aPfJuEj
94fG1UvyyqggdPW7BvQ9hyppWcx2DXGYs5+WrHIP8UVeQciJhva1W943rm3xgcwIhaLXutIleWYs
oRrZqkZRPqqNdr0hcgwTn9+MaBtJfzZD87sareE3Z+BNL/bdhALRtocHkpC/n6CZvgbiaejjw1vt
YGgLrw5t1wALc7W2//2KYBOwBA306h+0D3dMuRe66htfBmyib8MTtwytkyF/rRtPhzJe9zVJMnnE
df2sK2+EeBZFtHo4VEt4IWTBXpAS+WsaR7qZiCt+WV3U+K4COmXfjf8z5ZOplGxNie1p4fZOl6y4
QpQAlZ1yiiMjiIP4oR9qxGF530LSk+mpi5KuqwnIregHLsmIYON7eHJZqyG28kklyjN8ZyooVXUY
ydY9rIUUjFTMXPS1suuxJfVqMI//ndfK3cUu9WVCvPLX3uYBS7NOA+aN0OfxJL352qkEJoIOJaGz
EjD82cJcFMObZL+9DVQ/MoOBM+gGA8EFp2gST/Doe1115f3nskgprI2G0cs5vsUW5lH9UzOT1ERs
xDLwUkWBp6xy9kEwGasDMrIZF328RKRHo1b0A+Hk8xvpD5/pokPygVc583ll0TqNE2fM26pvZRve
bz+qt8vB1uYI66v/d8d84I/+zdD5KjED6Xl+syfhlO35WuL2FEVqHP16c5lHEU87iiHVCUWjH2B8
OqcxkisxDEMHrD2XQbARu0+ND4kWbumyKztMU/9nhIIAorztS0sbd3XbYQIftQhlpcFEvdke1GRb
7pRQusSDE8uQ+wLsP6HTotvxF/l1AaFcu2/R29OOI7v+pip3SO/IgKuNuiYD5OAFx4eEyNayFuql
hs1cwwjEIF5tQGPbC1Z0MDyMKBNsduvOHnh6veZlWPAuW1sjv34w3gsHFjm0O1m9kMnI3OvfO7eZ
BjarruXZIC7zS815CumnOlp7jjjsl/VnU80FrBRiEkFc2ej3wOBtmPCmQphbla3lBeHCeAa5xAAP
hpz3tXaLUsr01F6f4UoXIHDoNTQkNLxBtH6p7EJCsXWLTvo47AsLcaJUq9xocdWOCqKcdl+lMB6l
mFlePcR9UV7Eg1r+sxCB7koCRv8M2V9HTjyewFxzcpkynBXtYwnYELz3M52nF2/Dy/yuHZ+Ky51n
2+V8Ts6F1lvIiZushscv/Y/beTTf2MjriLDU/ZYzijYGdSi++VUDo1exDoeAaSL/mPU+S4jYucvx
7lQ7ookDb0YzCRrxNYjKKhMGY0PuPmvDrV8X13qehIGGdmzVYRyH7KqbwjovkFXOjL3vzMnl69jK
8V0bS2k0KAnodbg7HVR0tgjuSwgcobzfOcfqIjlLakR0r9UqR//zY/1+FG/n3DnZHVVvzSmUXoxI
yiVxpg1+8UdhnhCTlqHbsuY82lOSHMYU6oeqt/6QZl3LwVGnvI4tKQLuCTiy0FXdxcJ4Ec66ucHR
Pyn/8dXXvm8WhDs1v7UEZDI6ibaDO0zBjtVrmFUZ4iTcTSDfSCLn4Rc1mLmz/L/2hL0W2EONkays
b89M9Ez3gGvoOSb0Z7rOePfuMROTIc1HQuZBUsxgBel2GwErK4hqvQJnyB4ddjSp5vtlqVLfhAx6
KFFB/c376jPOkEkdxz8RrAmSR70QsIVVKqc5fNeQ3/ZgoeAeDdmDdGM4x0cVRItXQqpTy0wO3BaU
M0nCwHtD4n/dCTsFDxbKOOOwpAy/yywJX54c5WKqHjuwjcITt4EWlNKDjzwLW+RoTqTEq4vPZ0EQ
f2K7UJ8DKjej12TBMixxqbPmJEfM3dYQnZi1rZPF72CPsT6mASvw0gae0D9qdI9rRQAQmh2E2S5r
Cr8QpKYahGfHutYYyjc6vP37W8qiAms1EqQv7RRp93h9qyDvcV8m+I6v/ookS0j3eqS8Gz55c+Aa
g6U/4/G6pTndv5UjCz7Woca9FeHp0lysDojpEoPTqTxRXAXZE1aKTyVYWf9hp6K9Q1+7cvIO7zk/
25NZGXYDEuGjDcH47OAeNHzYKR0sIv4Qmo0D/xL+NLt5fwEUZaSMlwFYMTxnolFbYFUdUypQiTGa
jWtlGJk5vzvSYheIgQTV9yU9g61dmtvfvrA4568kHRDpi8zyGzI34swHi7tGJ/HSnYbCmNNKwYle
93YxkFTwWW1bqlxSti0LVddB89qIPmc2vXQzEqRGRriSsur2rOJyaovlR5/EAB/+Vixs7F6o3XXH
BLGi10hod6R/ax2m04j5dbAQY2QzFr6B9hqMDKtVCrP82c/qiY2M20a59XXcLCbnn5YLi/4DInA/
lTuKT5B81jDmZ1MDzy6FHAHOj892jTfYa7XKoJLKmVlOvV3RZldJeXMHsqBPLUUrLGFMsQw3qSgF
QM09T3HYUwFvzCNGvj/RQyAfwcwkq/AACcj8WNBIf8Lm6FSnR4uA+zMS6RW3UUBZpyGmJTGg4Tqa
6tsg63dL9Tg72ZzErkEf0q3Vruyv9VYKC1jeMfBN20LQvN7BehjNsUkWnDpfIOYuopRcA1PJmxWK
MMgPJoE7V+Y9CWy7u4amWm/zGGkIikjmmstYqku3BwXe/1kkkUrZmoTcneD1DgPOmJLjTgIQlmJ4
NrORr3tksU6L+myzaEgC87fMGNmfNIv5oYOkpUC3JTZNTGzDKGwXarzvBse/lEZjBh5wE4TX2PYW
wcKewDVAqaARu1Z6GGGTZXJMvh6YFjeNNgpkeJh29tQx9xfnX4vTcfPlSqY4QHSZBgHPmvqRYQMF
aR2Ah83nzpwV4YKJl7xIYNzlqg/X9UplHsU42/AuoYMQg9oLtpHyn5sz8fondK021a7jQujHtEZZ
F6ZxosLG7mT0gfUU7D29fRgX0QwNUhmcmL9Jskk6tIC+m41sYNLmnTSQ3K62+SWyQEJfMEP24arQ
6MNc43oKUl6d8tRLyDh14Zvgu7yIh5KXwU5ZELARx1WJyK35qvyheqk5Whb2wu77R8W5AozufvZ4
W4a1CloxnyzPfaZ+VOMd6bQJ3MIjLqr5M8x1hJKW/FOnxHKBgmHStEGs5q+GY/GITR89UHu5k2RR
PkwwZ0Jv7FCgffeOrrdF+nJDgrG6TFqvdf+GiroH0CUdS1ERJ6imDknQsz5zXP0H7ggJsx/+FXB0
GkV8hcM/Euym7Xgg4a8tG/MXZIdeVywvn/2QeGjMRPlYzqxrT43EO/ckkc0ifdhGszM938etarx+
Z0NfDVDZ3KsF0Jsh/VMUWkNPTR5fH5+PAdU1vp3hjzBTIBDaT8ifzzzsg0EzJFW3dfvD15+zMxY7
S6nE5vXiWcM9AN5fwfH7yNzTHPmCA8CLCngxsww8c4CNBXqlAsoAikVWtfYFeHXX8yVOYYWINQYF
R09pzNdeBtQnysIcAFo1FLUaC6x8wx6g6PdA7mfP6zReefhfLi5uhDST2jbY0ihOP4KixXI1Z7Mm
Kjsxd6E0rA58vC0kq9gJwkVRXBib+gyYzGjlLO+E9JSHwbv19XuuFNUyT3W0YyaZF7Y56F7Xa9u7
5KZtqIw+Dn3paLXhKrKhAWV32shAp5JmlIebNAoHT6BFsneOamrNbYLNkEWLGCqaqBAwz9hIOMS9
/MYI0UMTpiFp4ymiw9MnNx45eG2UALFAD0G2rNuY0qPMGyGfZjzYVY2/U/GGTYygvPFka8ob5deo
45Tr5XVmXwHJPl9WexOVcIDZVqJ3+Y2wKuqI0hmS3viyyPsf3tVbWJUoAdRHMgjpZiSU7fSltjpS
tgYsknkHqbHJTcgDilq3jGyMKXPm9uSlbUX6UUnYK0ECmigHe3N7vfVPqeBVgvU2ah0d7k/7vylR
eOCg70CPibojY8WMgyuxeJn5B8WOZS1VCBigom+Gt+u069sP91OfUyGlPDMwnT4O4CXOs/lUZmKs
AhRc1WNlMCM7Si/FIeiiO00t23J3td724FPGk7xXJqNxNqw/pd51l8iZnmqkoHteqprNtMPBrQwW
gp/OHI+uZGpBZHDHz5YB7AeWSqAO1dhYhLEsQHsAPuRHO5VSFyy8Ux29ajL6HOH7Rs76XSQ79CSK
tqf9niEyAoviCOrK/mO5/efGZWd1C/MhgDRdApAKb/1hWDCwrN8C/m2tIBFYBIHjRunolA0eJEmg
1b7O+f6wDVUGZz4yGYqP9d3Et03/ZrRBt00Sn2EemFuw76HMa38Yyq6I48qzyj6PbQwR7ihnPA8Q
Z9u81QGsoOX1b27VnrAh1uXW9tetGRSFXEDExl+TUpofwvhbO0GjiQ4jPKJAXQjTmlPWJRzZ0dlQ
0Jbf8KTF3mUbSOVFzXa8Ag1dC4z/pHgRuH4fLUbxR8JliXxkJNSvUYL4BBMqI+sqh6RbRiG/MXSX
qA5icXlYbzTCTZtfVoOPNrg5i05ypby3cnp9tZNa6CU6b0MmXDz4CAQuG67UhUjc6qGPhPHWHHqN
wrGBCrz22vdJyEyzeng4yapk5ZARTiGBKpsCjF2GojEqNf6c6QhUofcRmPH+cpFwgCC/BA9aeMHs
Jvn7fcXcnkzpFsHfi86EDMkgDQ/XunUPR/xjqIFoTtKTjjasS4KqlQU3xAigov1vVAxLlfFCaIIr
vwjwQpg+6Uh7xveMcSKmifBedykrdVI9ecNgxNVcMAiT5NuapEsyqPXbMu7zw3/Lc5VJR3QJaVC7
2c99K74g+50oomtLT1WgYaCqG+RPeV498QHix7wc94usgeGXut9xFsVgl2UxJ/hanUNr0BlfnmR8
seTE4Jg1u6nXBrwc8hGQECNJDIGHrIxSnsbAsWbXF6YwhSikIMPFnULi8POe728dpU4AuLXS+M8B
8CRMfVcsfakqtnuIsSBhKaiZCzrZDI5b6NuOF53ifGzLNMV7vfCTMWISZNer4LCABxrl9d13QXI+
zFtaxrvpt8Y1P6e0j/zy7ER2MvngYZmAqrOKDDswdlZ3ynWVcfTfIOxzjdH2zEcx/6ML/a820rRV
EHxLAdcYU6PZ/x/wC0XeaUm5IjcdOVxwpQbIs8qT8horQXSY6TJiMcBot06VTUJEAcNM4Ry63STn
Yr9Pu8qbv2awJhv3NLvl/Q1T8JxnMIA/UORUQmAJ0oKEy1rIk1dSq4v5jPn2PtGGTadzifWH9/GY
qET8YHj11U/yaB3IA6uYS+bNOoDT9HQljLbqmA1uJcv1x4EH9w/1N/z9cRrxwrUjak8YSLEYwjX8
L+DZJg/vVjmfXxYaERDYdVnvGpfe/Yd6lUiDV92veeZn0bLSNR8Ts3b5ODjUdEUp1vgGFgQSFAK1
iu30U41hfQlL2LjX3SrRmwl15ScPsU7t9sCjH76bjgBRXGZ1MVwS29DLi95fKL1elrgsmJh3X/Tr
JzJ3FxUBoC/tsKTvepBBGqZfaDbzNAnm55TA5itIC1ByQDSzLDsJO7Lb9lIvBdJYs667Bi33E5RB
75CVkO4uxVRFIPqVyqx6JpwHrheHtHuphZJxG8KTj4ex7mtVK/BE1mr9+6i05nUtbWIpMQ3d1D2t
LhUA+74f6BwFSD8y08tpHdGQ4Z90nN5VzULU6PVf6O0cKzSkLco5vSu9tYmURRHvLzjSeouAiFNz
EjK65t6f3NJLGI2tWKbDIFTgtySP9DZB2Znr9RwyXx4hPTupAY3iieer1PI/VQPDfquiIMicRC3N
62/kN8RvroiAOkUWwytUehrAvJLr20Aw5lEeCQZcH6y3+jwu2VW+OYBQBR4L/JuUQwFonLZfwJBx
pmv7iK9V5JBb7RgHTGfjR0CvthpRSNoSzTgUWKOM9wyqAwk37DzodnRDR6iOzlxg6V2iZYR2eUmU
ukXYvJOfJ/mQt19sEphtof5XdWy1Wvmo1sSFb+MMNGO+A2wQjNnMfibt6mZEo5Ep8A1qJXIx+3mL
pHoOlF7eI+iFKlFgz9sA9t5ElRxkevn4BDUJf02Lrbhwk/BvgleG/jGZNS5F76kNje9loIawa934
nNFpizXIaHbvi0GgwNX5DndSbabZGeq+vyN8BjG5X0zCule/JUGkMS23kjSnkSfgfUd/RVPtqQ3L
DdngIfBQUxfN4/G10hGc/VHqMMjwMPjffk7CW/DCg1BR3Kjlt0s4rHUpC7eRYBCS7LEccmQ2O+n9
kNsYkn0wiBe8LE1m/1+xzybBWMvV1sUE34sttIUI5nfqKneHdYNvGwrOolK7yCAwcb6MiQwJ2W7M
Lv16PQgq67qBHNFjjwCyMGaLmDyTKo2PjWsv+9kJlA3FZsw/sGeS6Pv1hZsExgi/4Pp2ymPlT7Tv
oekQWNNjtScynLDmcjxDpLWTzl+enHoh3i9v9Xi1oYRzCtXFacT7RHtwqXqR6+wsf/JdSlUWIrNi
FKbaXL5ch2mjU0jwQ7PmCU0UqODq1x13AQOmQ58Gnzzk6ado6zzwosaoJEjU0CatGpPhvfuNKeVA
xCz+JUPMcSkvQReJY8WKnmNDbCeyzel5InhTvsYejBEd2ok6mcAbqT1/xoRdnAAGBKABPa46f+0F
lXIYmYENcbZagJIQD3IIzeOr6xDvpypD389HDJ2h3pr3NbE0UH/3svzSVLA57y5fhMslaiL97jBA
0DT7DIUMvaMV+c89DPsaeSwu/fCzm2iGcHEsiKtJYycJFCZ4RdpKSTaYDDEiKlOvWKbmC4PldoB5
i9qBP6spESuqAcp22ukciHmu8QPLMGRqndc2chW//nkcUJQOHgQOmrgspV0P5icqXdsgRQ1jHK4P
LVtsQfJPyRQkiVWyHkVGwPw0A9W6tahgV6p3G+1bdam6jGxpbWRGgbqTekisUlsxtq1nhM1n3og4
J7J/omzCbi8TJ+QaHDPwkSXrInEisB9GDjJzvVqVfyYRvT+k2S9oYVPXrc1FPMCe5OjgoHtDtlu9
m6L8nXHURz3QcmDRiSiJyLnn88BvpW8m/BWWbDQTIWWra5T0FS0UjvCvIlHePuPj9yvNqxirB5SE
7EgTSne6lur7Vth5TlA8Mzmete5qa93Hx2wRSIwcqwH/25oMfemnsh8v/ftYM5ZZQkt6CYNNJpkP
apWes+24i6b8oNlG97hSbDUHrlC/eOKrL4ERVTjpxyEAA5n238UV1OCqV4A9DewQxCf9ZsEmFcLe
oi+YtbT81M1XzUh56WgfoAmRJ/DW6jZRDJ51sG6Hnywb6LaTyab3Qnw8YwEN9EPMSTVtFEYkWTNm
jbftSjc8ci5IPieTrB8oY3kpYwZj/ApWGLvSdA1fUZhh9+s1abJmKg17x2TiPkQB9zaUTbopXr1g
tUbYpu5EcISytUZF2R9h1CbPxEaO1iGOV2nFJVZ42kVro/29KkZcH5dVFfnIHYiBNOrIiEUEFf2v
6yZVotRsQ7L6eTtNLvK3M5aQGusdgUb+R2VpUt+e/f3VbCwgir8T16XFetqAsUsCOl80I/jIJffk
Es6VAjda/hk4b28v2JnW9C31i6wMoQY+UcbH2CT3KV49RrDuhlpDW4GK2tuDltMWXyzAjid4aIVm
wxkUXeCFxYgL2FkfwVhOu4fci/HkWdFyO/TTwW+cyi9z78z7ufXijfvzXSrKnu43NiBkldSYK22S
aGz5ZbGe2mACoGz0jYDgE1QfO5DvRslwQiNNN9H0BLha8EF/+pVodPasdzbsX9q8Dx8i/yo/MuRj
WK33e5zcOyyv38Wz6iapAye+2z+KA22E87Rt2LuV/LwW2g9AU/coMrgrddNZqL8eJ9BbThvowQ4r
Eu1aUL2oC6DzyFHdgtEKp/+492VX/SwnkWtRgMCscpAKSqw8hz4WgU0jWoTcCY8jBsbdWFYE/0ub
mYGKKoWSEkeLd/zKuxurRogqjbgSm3zkZBrsOsGFxpYxHuzgO+1U+Zivwq0Q2Y5Qff+d6EZMGvYA
rEKwcTPUrOQGtf1fSRzSG47uN6wH0rmCUXEqafuoKK/azbNzjsLYW3hG4lEcWWB36lyli8YGDAyh
KRN4lGRh2oxqYMr86gv/IqZjGN1b+MZeV7taXbIC+vEeCrsZedJcHLXJ1IuTGbGQJg42i9pygJQO
Ay8xxzj94hd0GOZBeljpeNXHX3NzPxBkOv76t2KePTtu9c8db2azyGmwp6i+A5KCYrx7AimAakMg
TbWLuYraRWf8cCut3uO+L9W1qkOtF6w6y2XHl4/CIimWiVjafnfHiItv0Hkvbfcg1BKIJ+xe7qRl
UglB6qyNDqFK/ly0L9Nt7Cf75NNexFuoanVkBDUbrLnZntqDsIlelWzkcvyP6Vwdr06i2Y7ZuAm1
QRxsQhq6nEZjrXRnbrvd9/zNIDDLZGRwPHRZcLdqYoY7EateEx4pqBScs+G7yuJUJFmDBDXmjHzM
FN3W++jfq2m61kld7HDGtp9Zy/nvCQ8tZmdU5usjMSkGib0Wd9CbOc+k2/UoeZcJuB46RqmJAxBN
Us+shok5wC2l6iJWJvxT7NEg31NBOST0yTeEmaKz4QsZSAUXv2EcaN8iBM+K96wZEcHlsBhucAVP
nEzDUDtvqV4MxUllJGJ83k2kTnzaGwJL2yUx8p/04OokhdtpMb3977ANlzxdNL1Bc8+hnfyLVfoq
u4t98hnCA3IMD85tlQSJ8ZdijeI3uPpidNwZzlB8cJly69qmcT0XNd14DUkFzJt6kyFN1Geryjey
vdgukZ4pAFGJ239iLSryq0picssbCThswljpkce6dwxLHYiE27u6ZVx6eqD8XXYEVpG1+9j7Ht+e
O++oqhi9djp3JjDGzfSLqzxaBGjI7ZnnpIo1V/NIXxhVThPVNBdMWzA8RuBJU47Gb7tAGaII6SK7
plKKcmK69vJlCf6V/7tSN/4/BCxAFi2Q8b3NNXP0nN1vzCtmJ61GOHIITKG9mNZX7GuV9g/ZWLzk
mz4DB0+NXAs/atD8QKGKl4hhie/6kySZ+FEUUVe3NJrbqFH/thd1oF7lFLY65jJT7NsTOQ0sSV5A
a/hDpv9Ltmg8eYxIWMUwmCWiLUmCiH+EdQy6q7d3MCiFd/EDZmVhujfDAMYHx6vx/q81tqzUaBU2
i/fdwyt3MTsPTwEx7JvCGjANfDHtnB5EcuagoA+4vUdypFMSt6nAK65r9tbv8NDLkBDCexQxOeZB
q6OdZ/uEDdZtbNQibLloiu9w1k1FFwLD54bDZMo2Y/GGe++D5QxY123XZDKrzcSgNmEj00ct5c4P
BoMCpQe1jYq1HMHgUtNRacPDCGMnV2UsruuvjgSL6aDANZnIkaSYt23OvPFy1CgE/p3FgXEGP2Y8
2jV1pywlvQdGZvwUkbZQxashUkM7KVFyLyr82C6MGhZPSgfXIeJ/a7/c7OkgrXTBbirhT7UsDZmR
DegKUYqm7VsO2V+QUOQ3FD5p64TnkFO74YbUJ2BTXX+zutRXCPI5Iv4K4c90AzTZ82geBNYbwFwx
MySdBX6AklQL/Ss+AXCowuccAqoTgfshlYpPjo/veNyYQOZoAsVapzfeEMk6vmE07MAaK73Yrnxs
AtWKGqT979dDEslJQnTA3Bb05VQqBoxM0N+aDak8N7coVG05Le3EJNEOIE6CSAGNwTFphfKd2tYW
uxpdva5cKrHk0r4lwKWOLXfozhzGPOuES19kgBq0LmVtb0CrKXA/Z8BzFP2K3Y+hghREdAlGbyQ9
Cwbycx++mpdixYeTf3L+859JP1NHxPcg5Tw03wzQQiUPk6xYzR5xhQFS8RSQMudqq9OFVC/A/p6Y
7JD3QHvZMydIDytIuHflMK6P31iKdNCQPI/kwwL6Em4deg9wXVESM88IZLM9n2U0XAKxzydd4gkS
AyhjCN/a4MbK63J311mNCC7UMLHby37LCxrxK1YCcAYGSO7zMANnetJmDbft+tk0Pj8FO/UWcgyK
lk2K1Hnib+XOMNnIYRWOaz7iqgXEMQX4UeXN3cN/mIiS3EfMAktD5D6vYUwKTO5wjG0WiSpRvm3X
Xx5DfDtZ31VoGkUCXcf0ntKz42JYu8g+3dVOyblvH4Fz5Ul3m3aCSrRVWnf6hkrynyETZh0pA0Uf
6DIFtQpgM4GrSszd5OJi2buT7x9KteJkkFpmg/DBe1axun7MFBh9FJRwwwFkPBME0vb2k0tzwn9p
fVhf36xkz9O8p0Eymkga8VUTNpkmamnJfvdxjRn7hKpcdOshnIYrrv3oNOgbt0u+lefF6He7Lqm4
fJ7gwMySkFca9Jt92DVpVwghMs9ROSTHYlKdnCQapsL5llwXbh63k4YtZjQbEyO2RKOlxc2yTcrc
jx2l6zZd/3KQl3cGcSjiNBawk7O39/XY0npvYrR7I7CmH7BGq9BBdnFYorpDAwWJmHQaNmcI1o7h
igiQrgTMRZbMiH1IdubqGMUquj+LXe0lkiSkwZwQgWqRrm+jyCj6bUL2KMLsyk9dncZ3+iueav/z
AaMudavpZQwJ6xNwtZZRQtdyZeEFiTGFx1dNF5Ml6w5cEdF+l2tWdI3AH2NTVg3s0vpR5VeUp7b4
zQnQrpNTP+Yd4AQ+N1K4uvuG8E5DWT9X8l4L661mWg4+6Z/NzCFFgnoqkWPEP1ONI8gnsKTPcwg4
MVkLGNtfWLG+1HEjfkCk+znpppdB/TbfM/FULMLmHDI5hQb1W8MAU6l8CeK2qSylf8GuqTc+ZIe2
OVe4+Pk1jtVUi52XBUGQ+d9wCwY1Z6BraJHQM1fIrsQtGtTgO9bYUswRmbiYNSqWfxvkeluBTLRj
bQ+3ZKVtOQQxeskRV84y+FJlXx8XwpC/+7pMvgwsMhV/wmvZ6+1aMNNhICJlrsOS0iglwbIv6V38
EzT4hZ1XS1+v821fQu01HN9mO/y48EfBVLUG/pCHegLkiKMqp10IUVryyumdZKH+gAfOEZvOA7eE
tTB4UPLq2CNFQaoe8frC7TykaX/559gmm/dAANiTM7pTgBhcMjt+X+djExzbuRwXwa6EsF6j1Tsj
PaCSorG3Bvp5QGsSwpCEjo4BNWXKJCuKBkq0XOQawIo7M6UhijPm1btmmU9/5+FXRwxs9IXVfCaL
d6NO44YhBBxFUjJRUWQyW78NcsOLczg0eMc8VjPJhnPlTejRAxyV+cyTOLwo/1hImxBkKvfiVAaW
izkPUF776sHtvvkdadi4uzlz82qQc6iCh+hrYVJvpTcC0fVMnIZ7E3V7qIDsrdCY/3psNoBl4GAB
EwLvgp7bELnQzo5AILVK1l5vCQBdtQ5aeRHKPEmBKhP2Z9oHaZcZs/+e1f+03KFVCaOmkjImIkXh
rVwuGlw10qoOW9DgbCxNVUHTBuMxCWpYpRtg1TDZ0nDlpdH8Yl/SFKTZuKDhZwjbPjv9h1sInzix
IvyUxfEyyC0Z7A0JaEZkyPYmtLcIcTlXS9d3i8ZqaEUXPiJCJGCkJlENlo8aVl+rMcbwV4OWIp20
tbC0YobeyFBG0MJH09uwGt52mRnH8Psf3NBeN5F0bOYIyJsINQA5WvcN8C8jMfQAKckImcC1nCBH
66z+Vum5p2volD0pEASx2aBgQgT0H6QERgOJ4SCZiEmL8rcE6x5BHxzSRBwT/vfD8K8VhFmM2cX0
wDdsx60KJebKpLkoAEn+ee8pyf3agFxZSYkXIBN2mYoIfmS3E+Pqj9j0mJ+t8CWzjhNJ8b8YwNNc
VBX6THqIMexiFbpvbhHf4McnBrzIx+zF04AKcXNL3uwWln59x75ce9dNd31fq9v2OYNz7xhQUf9F
WZjpwvryQWfmYVyZ9ySB6/qFvhM93mkAmho0g1hW1gWwGhG6S+ZcctKHFheB3UB8mPOFGN0d05yS
NEM00UPp6Re7mitYD7Hq+3laMrMkFuVwgGJRLsU5xYUGj1TfgZsFNWl9ofzKUiJX9RO3Hpj0w7yi
7HqJZhUlIOn+eb+OciwNr3XLdndY5P34pp38xm83P6d+n/9D/MmAhtJkeb+Vtu7SSqAEEcFVzGnP
EVwSSr1W1QaCz4eElt/YNyqNx0vmgHRMaM6TpX4a2a4mApBWzMhrI4jk4sDNSGlgaPqquaQSIwqQ
7dWACwUOsFrDu7kbKN1opydlE6R3ziWuS+kWsy16BwsP+/8a5OSGbABb4vs4ZDxxSH/bXbKeLVrL
myo+Vrl1Oo99pXQKKqOV3XD74ZJfaqP7IAZznuXLcuQh0vLG0NMpmoZV+BkaPBbkuB8SZZW+roQ/
3Z1xd7qNFv2F+wq9QQNf8BPLDLYBJ9XOXEEjHTmi0/M+3ylMqDhp+3Ibvsax44DknJ6pcfLD/wRr
ld+7xmyOakZ9Q2Oqt+Y1lvvbk0OQ2AxxkQORFsN2yje2L23bX02wNsDelu+eazelwxBlyNDa6Avw
DiXxvsGR9QKLvOIKky/peJcHciQ8mH1wjj7aCGQk/jIg1ZmIIIaQLAEri/XKTqZcijYb4vehptiU
SkpRg6aE6/sc7Er5Tc6ZxYqTZXQbM+WRwLzKMGQmZyVFPyBARzChFTTIxJ/6t2DvYMEBsZEjoZen
shNxg7+0ZsuNGosv2pfEYIfWCvKS+rVQSj58EOoqiv5HDA9/Afwqfjchav2uALciVi0W1AipYLST
OQgHPXAlqNoYx3Cub2dlC2OIOibhjboticRLaHiNTbQDQokB6BrvmB2AP3ht3TmPIZ2oOoxijF4z
//6Piuc4/JUHcvc1QAvKE6SUY8bpjWJ6gGRH9mGurJAnbbpgkE4s4VngDUkLpXSJehqfdbvi6mQz
ps1cnq+DMG2Z/Y84qbtng31XopSM9P+mzzO/gXCV2LQ043Y9M303orgsDvh+ENIQxXPbWAYCHL8H
4cgQxKmQaR4HbatZTloWkLBgtEpAwANup+mZoiAvXS7AUCsssEZhZgOWT0tIZo8MRX1OS+JWC2Hd
oWXsTdqECGY6U1oYQaCgBPxnl4vR+shVcSlU3AEJ3Qs79mbpi1LS89TaNCl/eTQSiDhSMKz5MVoG
J85WAHOmCSt6OtZCfKbZmy+W13CKcq143Y+/UtK6Qf2y5449EAeNocTh0/RBIKChc9iVFYPzsezx
A3oWlLu58cOxbJphKE2FLWkAED10kg0bfCSZF0IAaabdSK67bDbgga+JZUHnD5d+kKE2Nb9rZ69F
xMLjvel03rspbZ+XWdx+aWx+zIcll7qNABf99NwTqPHnSWzcRE20PCcaNaTo6mplV3BjbPPOE1Cj
WYlJUyhf5FmsX39chBr36H+Eaazi3DtPEJPyvm2T1BbJ5c5aPiiySLFW9hDQhMx8hEnPwiLPEM/C
1vYvAfl6TEKz4/LufIbzP469H+wfopeq+rtGxPSVBNrlur+C/dsSCpCo/HjPVKguTCOEz2S+87Pg
JmFEGgqlQK3Udy8U/g2ELF267V3/vsf0jzhPO5+o3afNEHMMtHOhWQqShzo6HgF/pue4F01Gjlpc
nD3O4BqORWLHHyjMq+bP62CTan+Vlj4qEsq0Hckr+R6hYP2/9nNN41mluC/enA7a66ke4PhE90BV
lmi524v21Zq+StI9HVFSqvXJmcgTf3aq6xSn9PXnr6NN8G4hmMF3ubjE5dmF0vBDEVpJJBacMBnP
Hd79aIyPjVicGhbMpOVcMKawn+xhnzywSDITYWc/qAbGi0tkd5jxQEG6LGMvQDBTWMV6mM982CqH
QWsDEF/s/QpM79lN0iKN8jc5yFKosZZHGW8jnQVBUxZjLLtwlde3b9JTtJ4TygtJ7wRlfLJ4nHj+
fK1ZMCgopkcbN45bLcsimY1DsqnnIFVBxHtDN8T8UV6EyhIZH3p+K2hYQurKvhfbHt5bu99Wf8Wz
j1bukw1vTzjcGAywJDxUu9KK6AdXGioqkYExUKV9U3cJLKd9FbWhxGkyg8p8VFoeCKeozM9wy9xJ
NThiq6MOuMcqUk7SomAquF2ibiORugI5TGKcyWNYH4dxVEq7c5+F2fzM6fiEbEikfFGv1HeIbMp4
KNKZj0TOhp2/6aV3VXMNO5StXgBPnVBNxrLn0MPvG6Je9kDVLM0hsUtlXCifObPJfTths1qcmzYF
O9gRX69hwsQTEJIVMYtCOn3r96+i8RRQPrvmdrf5+yyuiFmgvHGyB06oONLaeyNWcSOw+FDPM/q/
bhDtQR38GLwOldjTJ/BwFd9q8TAp729KOVW5YkY4Db4uv9lsRLfYi7CaGBA+OCH91VALMjTChbQp
UT9IbdvQ9a5mXHEVnjtN3ezYsJ96m/MtTZE3KJulllZmKVutkzzQWQOtxN39hbNeBXYJp1GxcRsq
Q/YcrqYFYngXmUBaEHW3O5etWooROPWVr3AqSqGNfCVs2PQE9y3g6+RaaGdoB9lSh50+bSfQtfM5
65sY8/W9F7aWRif/bZNQmzu6i650o+W9TsEjzGnLYswPOEtGC3LBf+75rZl6ZsR8NajbU2qkfrvp
vRv1iTHwibvpxALwRfu8yAyaxoaZh9BHFHqbKfCIbkVyqqeNrTzqz4n3EWHpOHxBg69SqH+Rpgrj
J9AmGhiZdF5hDQvWtWqsJlXOEX1ssyaLTUOzmBfGqM1PAVciXl9VUGcPIGkneWSKRctvU+He3z6q
5l3GUw73tKDl7STvi47KDCZY+uMWC9ETn2DU/FXDl4Ss7ZBGbYq1rmn2wUdo/GkYXsWoh6RF06Z4
mYUbxQ5MpcnUfj4jJWXJW87NvlSYmkEOUTldJLJKr19p1vH7/ORBg1fQaEf0G5f0Y6/fX+Dlwd3p
wmGBufGepbNmJhbiyy+WhXv6gTxTWy1bvByTtJuUi0+NfD1gpEw2111jikxEAqpxVZmYal9OtXCl
49NCuqv4nMglOTTAn0cDyJEo2HQAK/0jQ/XZJ3ncDBMRm+x0uO/9cPANDp+/HsIxILHKKC6tHQ/L
OXVXAM8Ea1PtpKJLfcGH3qosgjd5Q94caMoyySHiFx2CfvOzqyLsi9wxjR6ZVwKnEhcRLVAE3t7f
Tn/Iua2R0T8BX/LLWsvaAJyoGnJBeSdDM+B++zrE603IDaVTU2sJbOjaYY2B6MIfzyFqZY0iZTg5
FpR+luURuSXiY1MHWT8F+25jXh//XpKdTrF7lZqRvHuoIyNaOWGmgATs1MTAJt4C/IL6XT2TeISh
akAux3mSCXQ0sj2005KgYgRJeO25VraFsOahhdg9A28qkfIDIf2TF4QfJaKipD6VR9WW4VlihF3w
Nb9rpBvAH1ShCKWcojD9xllnF+NUjss5J8a1ia+ondO6JIyJsVkYJYsVlChO/zjr9lJ4bfjV9RAs
WA0y3dKPo7pODMOAMpIEKClLbZLuofG+nDoc9Jxa+GqmxMKNmCDHLe4nteyXNWvYNJ8lYLDMNLZC
yu6SvrvQcjBYP+JnCieQxO8OSSknJvSFzRm+AgFcFeli5tpzTvNkaiFl4rwuGwFt3mKBKm3PjiTt
QZo9wKmezb5XFmvwTJRRSG+Rc8jxoHoPZCeITGEhe5gJxI/z7L+vKDU5mpqqTb+F8ii71tN5KEqQ
xO6ugMdb8CUaO+Wk37+KXpF6RX8ZsCIscuPVHEKk+BFcGK0PCVfSWpaiQQpkub8TbO1mwwGB7zDd
IrRdgVUa1iad7sCFvip9oCLduWvTWVTX5PfBhRHpPm/j7Nmcwd/TbIyGyJZs1e3RgjpeBP93kjX4
3dEAJA/7AGvTIzZbhRzu7JY62aDk2B2KjmARdFMoHLnxvKUEIsTARULeEQck+uw2RVGibx0ekiiB
vE1NrJmYl4hqF62q3uiZd9LqEAWUxhJ4beYeFD8ECy4h3em4Bff7soiQclqNRugloJPBK0hY10mh
M7tdb6LOjV+QXwwloguf7p2cOesxQfI+HTrYninKx9oxw/34wBAowZDmVIHDn3TYdlQuQZGHo8Iz
p/enrq2J+Xx1OPsumwQgx2G3JOQxCwEgeHT1acxpH6LSNHG7MDO+PXChWjiel9t7dqCa9ATCqsjZ
e4A6MRHElJOpoRq7HOd8N3zWfjq5jp2aUfjn5v/rY9Ln9cP6dXcr9H/9wf1+mV0I65sKigvpfsCK
My1mzcVV4xOXGoFcnjQ8Mb/hin6WkVs+JxiRcLwCRFOghuCwb/UzIL23RL7so+N1pCmEHX0s8Fbd
TaLkmg/6jHBzRFBxqwNK2DSMFMwznteG1OtokZMRM6bQVVaYRIRe+f8gKAJf5e/r2lqpRQXxHZ+A
ZQ3kveFaIcHgypdL+wbGle9xcSU2ny37SosaCjkUYZViT80YC/HBhO8MG2Mvc+XIr/Nf/iY8jQqP
55AUcTM4ggh2qq+0/xh+Nak2xgp2Oj5/GbNA1W02KX7Xr8rQpOTZP7jU40kS8Jabk8XKjANB9+Z0
29COavFupiQDrNO33rAKiRkx8h+jNqQH41xsIElr0cDQQdHRxJSwQ8OtAgMAXLbD2Ii0FjCgPsii
3Cmw53bf/uKigJ1n/VHwRcr4ZpSMaUvJD6i6Bs5cYXv/WuiUT1UvQqGQ/MzP7SP1VsZoUtT4Cssp
z5We4zPHFI/h0N/5mugjJXxnKXMElMPYR3ycfGQei/jLHBPBEHjCVWokItMeEtO5BK//ytWFhsPu
7vnDuDgjtsNe/sKR1EMmNgD1NYM/0Nauvx+ukvta31NhXc21XQrxyvKaIGupJeVZqNGJNwQz+I8Q
+MIQG3R+6IZHgz2YmwYskSwrsUxH+a6ipiCHJrs7hI+tjm31q5TGyi4cVvo81rdWMC2PRJ/+T49A
J8U8xdCe06aAnwW4sNsae9NsXlImlIQyPdtB+r3l2L0MeL/uaVT6UciEVBOmmRJOdOpZBzeDeBFB
ehc16RzXhmY4sqq18KloF7Tfy3P6OE2evP+aaxbTkLHT61H0AsSRx6EbGNG+RwLyEt63yc1KmVWA
VuYZKBqjZwXb0q+5YNKnq640txW0AEJ083lIUxSz9mLeHKoEc0FV5YGKx28IYgn+EepZ/wEMG6+N
gZQ/Ybu2noEZENTuB3KpXCLX99xd1pycZuDPyPMob/3UEaWiJBpvuA6C1glw6MEWvcY2LfudHlDp
9eVfQkUdD+F1cqsk5saor2Ta9rrAdZs9dfNYo/AuIR0fasoHdTi5tNj5n/exGlLysCUzpLmrPBKw
pj+MgguaU47Izzjdjp65XORHpqdDAUxKo6BANiyKerr+VZFRGRUlU5HQmzECq45OfXDkSUXQiZPp
/oYxzqXTsonDc4Kucm5UE4BlTzrrzIHvqAS/skC57K0Vfb5Bn21C3dOa7qIKUk2PBWY3oQLCDRIZ
dm6UrmvfYxa30e5W10AZGv4CeoV8XRcWNlfYKxKfL1HazosWGdGYG5wPP3EiZ2s2OjF8lCGn+UzM
+n043vWMVkS2IcJxMwtyU6u41Y/Ex1mZPcbfuc4vYyiZuUG8NQ3mQB41Nm4ft/KU8CwfzBZdzFl4
lDjIKVZUJJFukQi+CUSvQeAlZtNPA2muIY9882SicIS0318uPRGQait8seUBfFR+hvV7cigf+LQW
CRYJdze2BKi4llsXX90oDrbIgo6rGXL/VW2tyThSOnfivHMZEea6F4Z9hGtAQ7LIjnJ+earnJbZa
IJMI45WD9DlfS0zTRpuJ5OJVsY9zGgqdr2VR/7NCnSwgDT9lVhrAEuhZhrJEMY4P51JjHPxnDkqv
WdN0LJsHPHkYjmLuw3OEeaNPrbwwREl2urMTOKRpBkB2OVMOpRFBloxV7+4QWW6/ztZOquxPyFwb
4VkS/w4Rh6n2elqc7ivwqWm3P46DhLWsw+2Wut8DWmjjICttc6Ow2lLQDiKbmHecrTZi2Sf+AZ6S
Dm1HwEepWXFFKIVH18+G6gtwvRRHk9etE5FdGThpHZAqz8zdivjC1/bMw2vqbWraAYf33o47X7eC
RJAjHIKqMdo//dmJ25ylrxTrV9W6mJ0LFyg8j2mC5o9nUW+AWpu9eAz4Q8UkSjVutyc1ZXgA327n
hQdCAjOXbWP4Nhuv2gEbeSQBkLrtPvv4srgQnGXMJ3UjblFfWddPSF2hCmYt5mEw+Gbyw5vCcAMj
l+wm0EGVZ/3oEU246Yq0etAq31cEMBcL/YS+x1E8BIGc/s5m7U836AN2cdoOr2m9/O36KLmnVJt6
0poPHRz/q9Bas1h+3Z1DdErvg57Md/iUAaDBFhrZzAC/igAc3nLiQQG9ASMu+pf0m6mrDyoOY8AT
Ol9SeqAqi0aBG8jbleilICnFOalLqjh90P6SFhoXiC5m6A1K6e4BWEoznyx9HoHEv3pgk/hxnoLu
v0zKmXGrTQs0q55WtCc51S/M59moSjZvLLIAabMQsdXWoOeT5vWAjAPtxoEAqgwAyPrHG0S79BR2
Bq+3KPF7YXKyatEYbrOOyCQTDOBXxlIleYN1p413rbRYIh57jrVpeMHBCSZMQZstCanrhHU0Jt6V
oictUkSZg7hcq/I7NqCTbG1oBh2aLiUNflL1Dr1EFAIROuR+3R4vxYJs5Tf3AVpBqxZk347Qkilw
8yJyjQHA9TPpjlrKrpNdpsR6stMWMLdOiDfvpgYpRnvYLj6nEUyO3UnL9DJfo4MuZAIcpDpGEk3v
zb6woJBrQDM+ZOxvHR5cvN/5kXnWzhnbG8wTe9/mSPyu8a9U3+QZJjdDP7ftKN0URBD6Yc+joe5Q
HgEaPorjPTp1fX33/eZVsVXnuUy9z9g/Akjg3/gzi7fZoqh1Z8zuPAF4YJHYNfZ0szhshpfsuMLl
XsClDrU+zN/Uu8yrpcPugN21mP8eVqT+Uglmwy/Na2hMpeyTARo6KCkrcdqd+QAkV6Wpq1a91JVo
CnzTW4RAkTQitcvwLMn8JkflqYZeBuB9EtjkYTzOEJDAWK/9KHygChMkQnqjyZA7vzulJz7vK3E/
6PkpihFfgmb5QELmSb96A5N7VzJxtl80Q7oTdLwKDl5Lqq4zrjLK/JXwUzsljbgHHUAlToGG6c0l
CKiLJG8f9jTYa3bR457GrjlEcra68f8+4VoMi8C+7KaEP1jp3hVKv2StN/Fp/N4V40+6U2onGTb8
jekwZv+/GA7JKy+BhLnbwWMY0M0265pa+MTMSqI/xwORaWQstFLP33X6DGNEyFmoBdSpqdfRRV+z
LnXgC9vipi3jlAihiXKbHe05ZfwQx4ZtT3zuZtgJJSItVQX2c/gNKlpJkLr0wAiiFcnfDnDvVzW8
VrGl4IpHcL4+3o7ORFJvbwMwelRIHx5yZ2lyKsk0Ga0mwWp7zeqoeYfrrgv2XTSeHI/ghom/mY4H
1oljCZAep92kr8X8+hIEzfnJ6Iedx642ErZSamobhT8ElXHPdUuQGBWuSIG1ZHeN8PXuNnF5a6d0
YyLPv3LBrHcsaAR8AqwpkZEoSoOw4BPt+G5ugJ5l/zhiK/eKlNe98jpVIka7XMIxSXAGeTdsmter
SrjpNwUu2WGyD0E6tfUSKW4oWSKjsIrvwaOZiBDHbRur9wm6jC57TlY3gTNBnKCIZ/U2keWgZHp9
mhzjMhzSD0ll5yfgmeAnZpXzKe/h7j4sXUmawJ6Cc/FyISGRM/mYz6g8PBsJ0Q35GfGrwdqbI0Zq
S8HgnO7YRotQzv1RPjzpEvm7wn80M3yZoSww9ys1tE0HkwXCBC8Ktl9w6NFhX6pfaD7XmhQgaNoK
7H4YEoJuxb/8MVg+6qq4+RM4j0PzKSUwacPKjV5gPexDCU/nQ+MbYzLKgwpg0Nu0aYPDYygw/JJF
91GCX/bBS5PnFLgKsLkOEu+L7KNR9wFx4kqDXrQdfDpxl20A1QB73tjTE8REKPZV/dUoBDfLkQ6G
g8F7/I4eLT5XuKKzIyznZSfirEA3QCv4iHG5SmxdJDqk+mojq/CCNtEeKivYYrrvkTBr7nev0/aD
PXDspM2FPWsy12ZrsLAmrxxco/Kp54kPcQyBvnKXODzlYPnrApHs8Wp+9GB8X6CzJhRsFRp3ztbf
nCVcEguKjLNZnehwFiqZTkYmj/Kb+tqDbSbK5X2kw7sSvEfe1suxdZGoWOOf/FQER80U13EmBa8n
kiNfwwULbLfiVLWc3DvDd7Yd/JyP5BsmxbAOCBuZh/qDga9/K0OQ6fref1rPx8A2Ujus2sscmT7M
tKWbOb0epYLSqKYbSJs4ObDVQBCZPaLa/fFR7ixV8qC5JITEA1spN/snV8ZLm5nmOtw2Jo5obDGf
Ug+1JaaauUvVa+4f7HD0mgyiiN6uXSQTyef5mtq5/pT2MPLJKOA/EC9snrX9blcT9Tm6dSrMZzg7
OGv0CHgvBRJ0uy7/ccmLRZ2DCbi4qOKY9fTTey0HQFfGO6JGfnFg3+rPi0sScCgQELtGRLQ7fJ2B
ewSktK24y7lSdlAuMomvpYtNP2hxtH3X+OBGxMl0ZieQhHz6gplKDGH/0sKZSZD4XoNBkkSrvw68
VYjfmBRwfvFUFChPYjKtnrJzylr9QvyNXy0UlQCByVk82joTj+1N6/eTEi5MeTlUocCntv5XZhoD
2Yo/yg7FNK7m6CdsZfX9OCjqnHoOK/Md0gox/1vEvoAKy0B8KiBqkQzpIcCCi0/p0RRdxPK9AlYI
QlpbvV01m3vEYSjPUD6QzQ+RO4DqXCWQ61KRMnV+FTuESfwU2cT71oNUEPUQIx8WuhrsAdzPhyCs
KMfivDYClDWiNjnThwyVtDmcAnolsx0SXeQmO31f262s6vUXQGVDkRNKK20uSVF8/gegivB0rzzn
6sY1d6vIzejI0oFrA95N1buKz7rYrAJ644Rle/1MVLNCFI66ADSvTGmNjziDVxtmnE3EBasrgKgb
TtsJsdg7CYUd81X+h+SdJCTTl86e6jcNmyvTY1+a0frGu+DwBa1Kzs7zZlZ/bBgKochwgeMRkqfJ
n3/yLElAUG4/fOKKDzq9s+8Lam0pnopKWviBa/KCp+mUf9YHU3A8ZjHtu8A4KmoWGZo/MUktXfVd
wxkS9w64N3Jl5rDrYv1Sg77E20tQgLcgiMw94RPrg6ZspNLj++vHwefoZYGxzT2pK/2zT3xMVQK3
YQ+avoi6OhM9dW0X4OaJns/1sUX2DkEx1egHk0FnrJvXzwgDFDNCUpemjzVmugAIOLcbtjTquGWZ
YDmLJLVRqtahvUfOTpehfQZZa2iwnSjfNzV3NN81Qcxy+dGzJ7tUXpmN4bCeHS+SdYhvo9YHrg6p
4lolMm2smvh/jcCpbbrN+jqS13OdOAoQKgsfmt+sABUZZHh+2HNLLxgsODsIm3jOKx4FGRfkUrQY
3rdAC0LM6ko6tpg29ruJYqRZZVVJgoOS2iac3JbAB1yxVAGm/ohEf8YT2rvb8PrcJIKGUf7hSj1D
4RY0zjW3xZ63a3VTvpS+sChJo+xNvvBmDb5L8tAvOFtReiT+FZUP7pOwAjvVkaMolJSWsZwuH8sQ
Et0YjdWRVpJ1oql6tImS4mFBPWlInvPBicUE2okZRCQr2MDwEjouzzEDjcFExxPIk9IdJg+xL2Bd
KjWlAo0vxTMR4AQM+JmtEiJaUwbHgN64/gC17KaJ6CozbzObkYXyb7rBzHXdVGuZh1flyZf0iKzg
cEbxNy7AqhZaqVvhib16DFRsaD4g6hldxJWphtZcXE9mqOs9gjOwsUL/q8clnTo5oLAphNDcLdRo
nFyqgiijb58kTM5ryBllZPZQ5RZyPPlO+BziNlCQ1/dC1RkpdTMbtlfILXqiyS6sA1z9wGLISZye
nbanQW3cJYXAGg1WSQ8XeH9diHnUNAnfbUogmfQc2EPuucCRDlvDRukE/fBVC8lPrR4eERPaPwY0
hyrxMtvYWVCUGxYEu7+p1GxkYrOgY5SyykLQ14SftKdD/5eT+U/wDPGInJKGWDc8ZGXubtPm+LL8
DU9lTStbDLNig33tLONd14nzvl5tKtTrmHuqfP/rO5HXTXgmvcErz1SJR7qod9cmC6LJha9n4quR
vfW231SQYt36MUMy3T+gfhEKsYpJOVtwyDqKZOqiCrOgAiiAoGBQN7AwW0jOTSd+uTDn+k1EUJ/2
0gtPldO/7Rxbh1kUNEadnFXz3RAzp+i4p5xhW1gYsKRU+3EYYZHFhXyXfrgWzkUhTxNke8X4PxEY
Nn3RRoSsgzvqwEoIPCUdjX+BHcm52y42tfpIPAx04naILuv+QdvDYOQgLa4cSvPl/XdFdn3i4pk0
UozxAHCf6hQDT86fq9770Yatj8p/ZaXpxd0ivpLGm9S0PM1ZC2L5rAWV27fvyJvbTeakE4uRdZfc
OhNAQCJkgY8hRYK4Nf6qr9Ntrr5XzEvWUX9VTDTkocseFU9M2tnD04R/X9V588ODpW6H0xKKISL7
LZCkrWpoUUS5xJ+H7cjjcZjK3YAylGXs2k4PNd1F5bhsiMC5MWt1P0SsUKmgHcd46SVL1dkwPWu3
YunI+0zMvuI8q1qzkjLboyVI2cefnukiGRjgp026JYWEsFbjw34R5oGe8IshLAfwLfJ1E+gVqazc
aQT8UAb9LRkJt0becMilLI1xKmst+1Cn2xV8LKuoUcnTkrc1+avr358jJTYK5VdLcLpbJZ35eGQ5
Y6cEiZvVGXQDBF/O04wKkGMxYivFrzmUsPU8AAsDRcqvsTbiWxkEJGKSo6oHKMmkUP5iXFaSsDAH
dbBSWdn/CHyQHdmxLOR48RgKfmTi6a7eetObPE61p94SrDL1J7h5eMnvJucUFGuFUT1NwYi0WtuT
+0CakupNJsE/iIgrMT5MV/Pg8Tf2ndGzM8+PHrpwCHlWVW2y52VrLPcy+fRMcAN7w4x7jxMU2Hqb
S/MpgB0Gg1qU/qNqiscWfsUL9MXifE7fcSFsd4Q1K9mh3vQxEDSFcloWRQdagIpHuCpKIUmbIUR7
1OvhYfDxQIY5b0Oan2KggqpK3VDv7zgvvvEP/AjhvWqx9SMo4Zi92eX4NdPHyBtypOTPpqjb7jaY
ZUmA1caHzJlmgzUkCh6Z3XdjgJOOAFVOANtx6bJwuUCI4zth85xAS+hCXIra93Ab9AzWOXDMKpK3
gtUEZ/ujqYRD+6CGexS0RQJWUdEG5UJrwpZmdJf/w/roofHn3IAqtF9Z+sZyb4WaU2NJZs57Mbaq
O86x9bF+AYC4Dnr0RdYalLiVRDTDP6USdZynaSaKnTtAfR31l4txVBhWijs43sLFn8LuDGG+ZNbV
nLY7lQm/FpXaFLVsbY4w7u+eqPoIu2xtp+U8d2rlN0BPb18lRotd6LLkZLKnJlrzGTQp+/bBxsuo
xFHdk9bVI+mi1o+F/3tvj860g8VMir3usEyu4iFOBWxn9W4LU/svJOeBnk4hGxz3rVhPI/1y4RHL
OXw1kseHpxYQaNg5pCW+q2a2MXa7lmCvTWRdfft2ZnCBVjSRhgm8dEltfaisk1+5GJYChKp7ReLu
DCCh89Tp5jEwWkZ9tUqz/L1V4uo4s3Lekh+NbBxMqElvKyCnwM8OZ7hLb/C9zxBK5zUfHITT5GJ2
N7iYHhErNLWp5TqQ406MLhHlAKg9LwWf9gQd8SVtsznkl8MuNUa+5WSc7hzXQBdxzPqalR5Kta47
YHe5IscsIM1cEwxqARWLTjiC0EJFIGBjq/9MAXJTF8tqoVHkWcFrtsP77wfc5bJAi2zraz1YRlJ9
hObvT9pAG7bYIB4LNaucXSgw3Lalp1NTwk9w7NcYgALWDplZnE7rHTBfHPi4efbNmv60iqPXQ7H9
PMgAYNOeiI/MX3VBbbaevA3+infOPD8e893W7zmexoZvfdJuPQDT3nKAbg8mIhEBzBpBwZVjYQUb
jTLR/qQ2Oy+J4xeayR0UjXeP9e8WFCeJkMuQPOksymuUaS8ulsjkNhAevNA31CFIigx7Gr/RS6DH
T2Irr2/9WUevxKX1p5q+14ZxX7kC26KN7JNtpFjl4ui9yWIycqR7okkZ8YFH2lO+SUdnnfxJzV5h
LxOihtQ6Txt9M1WNXFDQSfQCnjaLIgkMIyh7NT9rbN4mQeb8JFO3vjl7trfIP9m0cLnzaNhcjrMl
6XiE48EMMUIJEgkzhBSdzfsiXW2g7Lf6gOjM5KK6DjaRCxB/tMLeilMjUboAkjQBxyAq0NNdd6r2
v7fwOKVAfLoU8J1UGVEUeCVh0l1RYUXYLJYaaEOsLIItYJuvbi+bYM7N3PS9JYvHpfQFLGZ46vt2
OqrVAbGXTV4F1QZc6k3vXn8cJUh3OKcim/QRL7ZWLX4jt2Xey3doNfZ4PZZ23K0Ir3XOccdOd/vY
CS4lf75HFCxuYFSxwPjbYXkjMMCzZmHpcs9JH4YyAZLfGXcEP9aTSigpbGByMujT1YdPvTkVbf12
YsPTCxCWsOqN5QpWF1gcqBqvKIWhmzBum9H6RQVUmXKi1mheRi+97Qs81Z9ec9ZHYkindUJamVpz
dS3tShzASI9iYyUUb816NnH69GQUZJCaRrz/htcvU72Cx8lVb5+aNemQodGgZq+rMu0ra2ZUJZgB
aJ9NMms+Bvd1DDmIOThKIc2/VamFjNX17qecRXOv+aMxT3KQ22qWD+SinGN70F/W5OM8/IpawsW3
rcV9jikDxiJerqugHCUntO7BfeAFbGOuX9y80ce4hF05outUtowGSx4BYWfvXoRQb/DdRy1MYa6l
Rc7kjNInl6lz05qIGIUHTsq4WCFkjVJdYpbqam+on2rO+DoF3TpQYHDPMcqwRFAaVkHUwA28BbnY
RqsuOVIBUAKiEV6+61RMqsAz35QQyffR7TUa7N5qVeBUwna5uESD2DGBDCQf1sPNbQ/dFi123kFT
Bc4v++HElN+3jk6dHJYTttyIJggOs24UQUd8zalFqG5Js1dLsDkqMtxfTwV9EAcs+/rXXcrY3H8V
vnbn78xrOguvfPha/suSsoVRj1edg/xLto0APLFF/JxmZ4PHhhVAFufU2MQKa2ZY8W3Awc0ISy4u
JPSjXR0ORiViRjG2m1+vF0gtzVkmZqS+g9YzHkEKJJOc2nKKbiPeG+3mbjz7MiFw9cGqDEbSXPRj
nQ/9PELve+UOzTznpagAyWG7aLFPbol3QBE6Eutkb2BpIc2ulRjFMN8vUOB8tq1kb6+gLAgS/QFO
D9H4tKiMCUUs70BVQDHEQdYug/i9rJNYXS1AQLpTYg76P4dPZxlMAgw0vMIAx5vn6YzmyPKhjkpB
5QkK0Z/EMFXWw1lSPl2xzy32aJq6xu0G2Fe8Eqzxz/igHoCn6kOpuqok2Xn83TFx7etPdyU1wdt0
Z5qNGMzwPIZ6KeNOSpLWdvKwz4d5iSKge62fv4LQyQ8qSDqWRo/e9tweNfAGeUbOGTGUr+JNIgJf
BRsaaf5UXVDMQf94vuTRtVfNZOwQ4KI594GbwmD+3X2N5eK50euOTZ/+XIKnYx6h73RxuoJC5CCM
z+t0uMcO/4rSn+d28DFRT/AUn6GLw0M7kdm+5EvrUOvVaXzPrpKlPbm+uZKSm0JYVrnvx/aeC4JN
ALKtsVlAtvgYp7P4C39R7mDQi6jF50M1/CbBG09QWq9rvqooPNybReAH34i8688KIyIZMwmKBdfD
UX6d6jMirupCJOfislkYSb5vDfCdl9orA640eaac3DFJZnDoJ1WDPLfOMhKJ92DQ77+4yo9FjsPn
SE3yVkTzf/zue8W2v8egEjF7Zf+xs3m6Jei76pJ5aLjI+O8HGCJXui+HO20zur/LWYSfYSeVlyNu
R7O5QRFfeHYFyekgCtu1mk5cB1zE0Gc6GbWAyr0mDB/AJNrbq763XW8pIigq8ux9vQWoIg2Krrir
g3qimsxfymUKi0KmknG+3Cc77JquJYTJ2rM3KkNdPOI6oBslFnUDyh6ZJAY0QZISNm9f1PTvNDQu
i9XsqSVZVm+ByDw2UsA/iLQhrZs9Drg4bkcJ7e3pYgFB6Zy1wI+e3Fq0wOIBK1cvF5+mE7sgzvdH
bCz73gVGs2TJY3vLDxvA+khAwmUfmiuMU7Tp52AH86GfGJl6i7F5fIkwU31BrtE7osM94j+QzjBQ
Kxr8JXOZhFE34DEc9BoITpW5F7qHIeJQTcoHKp+3G30EH5JbxjxWOmYC1vzNw5c89PSBPina0trv
R76MSALJVqyF9zeB4E4xPKd87qJWLpMCfwO5Km765AK1c+CeIKgSU2Usbwv8m1itiWtqZAjrje2m
xRflPpzBLh3ncT5SDUS3EiTN3553AMpG7vNDs1HhGnjLc5d/SKB/m9x3gxXm6olyV34pnbSYTPe3
7GCYxbau9arZvRjgJcLZLDE3JoROdSu9hcw/zfOWFp63Bzauo7JHznqX863uOYDt1MR/qJ75eppO
+MAfyMS57PPVmhUzTC2wKA1Wp5l4pewKxbntICZDmeriz3e3T5UPLRlY/R2YkvE3RzmQlYaWRcj+
uNrdi91FuoTxl//2PFnL9dSpepdEtn+YIgZNa70C1pXsQajZdf/B8X6Re2E8Ebh5mbVvBSozyObT
oM/Yh7990ftR6bWs91U1XgzcN/LWRkvHArVzxCs9Sazxa9e27SEKDcBoUSir500ccX0gs1sJSrLC
oTzzUTQUmXcCiPDHxovY1Cck+CJ/QEmwQyyEDSxKZwokesXVM58s31AW0i8Y7a0hgPDn8AfcXyK9
QPXvdbLxdS36zfpqbXky5fJ3Yjfuhmtyl7kV68+ml875jakjMa7Ns2FTJvZYrWYZgG5REVMzuE/E
ICPTl9B+UI8/tivG+PaRQawsY75fqn4S6eMnS7EImayPm7VVC857+N+9ivqyUNNPUYd+iDg9wkhO
4WSBcI/kjAm7e8Vi5v0ME6A2qML+03H9AEe/HoXElqq5eZ5e3AQsQ9v2aTmiIByb9hl+DcUP+QMV
JSWgFEKBMpZwKoc1CkzdnP/sUwzRteCuBaOseh35aBdbFBttBV5D7Pti8TQ+ei5gisqzQ1oCjAFS
q5IjNtvzCTV1x1BlkKTnUASBE8QWRZebCtqrfYkNoDjesrEz5hL2jwGv+pIwNKEpL+Qms9FXxRzQ
hJzJ0rJfA0iz+V0KE+/t32arWwGGGtNNMw0Jp7AcFeYb6LlThJRMqDL/CzePnAfIdGO5xwASbNxJ
h+U+qHC6SG2Nucf7z0Ou98n9BBgkvxAY8B09EsEPrsL5AfUeiQzQ1wfzqRsRp0XUIidvKODpcRdP
FnGMKg/kwavta0CL+7Pyo3CZNIoyYxkd+4nrxveXiJMa52BaJWGlUbsHNXNWehqqQnvuSmzpYO8g
JTeSAxD0cpR2oKORgUcj8UydiDOjGgbE/KqUrEm1ILb5SCZgBkTjr4XOD4sZe4oLikkU1jUH0IJA
3SS4wNgzX/pWotY6xwxZ4InuJWgqVuDrI5r4LQxZ3lqyYb7CBHa89JWIzanZRTwHEL4plB45SZca
HOuaYaNndXYhDv9nEnI+XRedejKukvXSuFO2lziXFDOqesbuAw4DlPbw4hzLiNPSfsXidCospNk9
aHThlfI4KeSHJhTYV2LPPtffVsDcxC2Cfmyq3FNbyJ0SVvAHrmyTtBdTYLXthhEM2UjG+qXEV3aT
UdQjq12rR3r6TRGbQ2spVGwasotVn5kC4toV1e+W7zVTnMx73KTPiO90ynXwMb9NyMmQiIxkOG9L
myJk/n6WW4dwEEnZ4gRrr7WZNZFTMjWzjhjSQbLeQl9C2/t62H8VZKX/AO8fhivIEx+yea6g3u1A
19QfnWel/hINIEOfaT1gPflGe2PuCty5jv7JT/vi9rSma831UlOUWrhzz4a94ALmGzG67n14AW2W
HqapEsCKRzGtXQBtheQfGWCv5bUeTZxC6skF/4Ty/3WEqnTip0CT9361xgIfqa8N6OEef3vlbigy
V1JUH0eJw51AVCOWiBgz041Xy8hlS1Otqfmk9yd1BZn/8JR9NojkAH98e1hPxlHDF3CDUPXRoOxt
evS8AK3ERof1ALH+BLHcwqQGdXbZSiJhLRvikMylT7zs5Ll1ZiiR7PsDjLAeugXMJzFh9XWJPPyf
/SG3cP6XMJ+MGZP5p8Y4LfLZIRxfTej8sfRRNCsWepn9KJvuoKq/Wb05QgYtJBSDwRNsR5bGMwrX
aJ7Hv4ZGrmgQXydbbyntZxFBqdrRkb9tUFNQtR7Okt9nUMgNLyffUx0H0IZjrjgDo5zJi+d21s2m
8tN7xvhOm/avrjkGD4tc+j58DrztJoWWqYF6mbn3C7EDx4QsF5ztaA82ca8OiFnhcj/293aSCVya
yZkZGXUNIB5UvaMXupSXzutThMgP8FxXwwgzOYLeYf++wydW3aX3pFmN0tqZjq+5o6cyLYa5PoIX
DS1kCLDeNO77YgsJJgJg1RlcPOJ2AzsyiPhSA+d33y8Kfs9Yu14063uZ3q9xpEnBW2D92bi7iHs2
KdddyrKUzPBSHwUMgPk2QySR7mqKdCdqA3D6BJ3lxmVbqYrh5lz3J+TUlf8j6w7S6si4NzEMvVHd
SSyBn/6nL3riuL7TPEL7esmPA2j0La93yT6PD6SRF8E4sKSGvCZhVm8b5DyYI6Vr+AWhRGM1tvb9
53+Io4nkTYZjbsUvEq7h+lF5HA5WOJ7cguR1CrnqtQq3LYT5eoWGclkQuqDdBWKW2tyCn3FbPueB
ShPy2e06unwch3ZyOx/bbSab/goi6PyboR8BwFxIHSL6l8a+x1v7q4X5PHtOU5GOMmhY3JIBKXrA
4NgYtBiOsM7N/A4aSFxUMKzo4eLEspmyjL2jaOuLVn12T8Pb/z4Sg/r0jUF6iO0L053U4ezyWXcC
bUK9buXAFK0eWPb/Ms/MEuv+ySXCZtFP5fFWZiVkO6mluTuhVWvUGC+SQsiwND7eQYhl7jJ2RTzF
Vb3aDACL2p1ePrBUP9iN0dCds1Ma6kIbUo7T+kcEzLXMKa6cs181hwBEfnQyr6u1buiQZBdUPiUb
9jQBLHlRQxGiy2ez2K4RSoXDYSsPol8o0gCtghAsG2INteoZW96Vtoiq/eAc/iLmxC8zceqLfLCA
V8cKUbzCIrd1Dazm4DAXHCZwbqMo+kVEtArBXO7j78Ky+/tE8KEvo4OxmtGcFUYCgiaBmzhDb4P9
BOUZv3POqFkBbxK2N0MzNYDH+yeF1x2QWOay6Vc252LDRBsbRanTh4jkrdqXxZgLhGQftJ77vsBL
hJ99kamIwLm7ZlICpLTXrz3K3NdrGEO3siAcN7myhAhGcFQa6UKPd4YbIyKBrZkN1Vxrfy4JYI0T
nbFNEmdevG3qWV/M+z1eEygifDlVSDuNvs4xFsRydXAtJvWS5R5V9afB3xlt+UivyWfu/76HG47N
0Ch4pgy1MwNiFBVu9/r7XxAXGNUFJJ8WjKCCrFSJYp811E+Rosk/30FU6D91y5bdSZWqZNVKct4W
MqF3Jbq1ekJtfbcR8+buBqll8UJqeVEU8YOEAejzgp1CJ2PtXSUVySB68kWrpAPB1dIMSZLYlZAv
UH83bOZuNuW+CREqfGXhuUDo4oWi+hwODjjaYYe/t+OE7cHGMscMfJxlhQacBXZZCWbSLPiMN6lI
jqdxP5/jw7lgS0bxAwfw+itrH0I86qqM2AysCi6GOinXXzfz9QcIb1XCZ8KfqLeBnndBNJnKNa4X
8q4cAe1H5aurA3Tpd+W/j1krRdvUceVRwu9s/poEBATZZ30NjW+cd7nCYE099B2BNHC75Q7ryrVC
AGfhFGMd7gCqrcfRXFi9l0Zy5/p/v7xIxuLzBJys/9CL5wizPKO5P92jxL3yHk9zT6aB7Ioqq6OZ
cWqEmq5+Nu/Qp0V9payKEqO26K5IlB9D6Bz7aWRfsq8oyZIfvPa7PldiP3pWEGCcjg1k37ZreSg1
4YwwC19OO/IjnATUvF5eq4h7ALdjmAebVaLrDwEJVuoz2Hw0nXvjkVFGtiFjD8Vcdxuj+9hkMncA
oOEV4cAE1zRc2J+QUj+KUYgPzWnp86hZBibfRHCpN/6KxcR7oKu/Nyonr6Xam9XtQbAFqzlalDux
3ExV/9hYRtKyA7fTy/TAATWR7aK5w0vtmIc5vQmqMiXEZkfxkvxnlUp/7FWi4zHfUjextb8PuwQj
BYCu03f4QEYEVX3dX7fY2jQXcZreBFpxnyROb/r43E0T9O8+ugEMPDjYo2zjGIQxas4LWwAI7U0u
2mfAnwbe8UZ/QvNrGLcAdZ/0T7Pv1txybd7dl2OYFVJTeMlCcVZlN0YqSUZp6r6vWko/Nej5lcaz
oLP+Y0YnFu9iV/B6iEFI5oQt1ED3Nk3FGWAb0m3VkVSrElP2e3AxjsvQbwm779o2nTylO0OKdV5q
cy0FF+jI7tSmqqSpd3p8p9mKpTIcLpg5fIOnKVjLAw+TNmCa40Vs1AZdpiHgI5toyvWqVy8Dxdb1
tkynetQn+3STE+jisU3bYwJfEHVHqNfR1++fHMwSNUGH4pnKXvjyTo3BRsWbYFLaDX6r0yoUZ39Y
d9zUExULexUTFtb2S7lSIGx6Q3Gz66elb+Pc/QiOND3ieZUhpivnkorYWLajMdlsr+QkAEtpXqqw
KuebOjUBQCO+IpGb27n3y5YGdlZYB2MicdozQHXWUCr3jZ8coXSQYlpqai7zrI8RFAuBhd+AT798
3Nkq/BXadvTaWrSxQfz70EvRjwD1Kjh6RJ1m602D+nyEAvLtj5f9BhcGdbSp6xNQirGYV3Ws4zGw
RcdAILtN+z6Vf01VpOtxyIHh0IJVVMrpcBcRS8W7hbRfZYzgbpW85aO25Ujg3Si5XkdvRP+MIUdz
aqupcEmMlQrUqnqml254MXoHmJQbi1An4H5mr7rWVN1x7akekDk/wj1iT7ETZ4R7N4F/9l4f21oQ
UXnmJMNw5C8IaB2QUT7PaaELF/WfLic4PLNonfzoF2VMZOKCGaxsijfi7jqQIgGpbbDc1R8swmIA
4i+IVKO0HqHAXJMPSy4VD+b4Dk+zutWRbtfIV87pKagvXx6cAZF6eV/1SY4ZTIOBcU4v0HCBEl3b
etp3Pnv5skXpPMDbZa0pERuKv6sGZGTpkTEtdVHhNEwmy17TflElASuOX8EI12z/kQWq2zTMrOH7
XJGO+rNU1GvFxmJuLOrRO3/KXA6dYDNil+iCzlmtdnpp0qltMFYOndkpgxN+Ewi365VE/7swoJkV
2b0dml16Y9iBaoUr/n5blDoH84lqNsezma7TfAKFX3NvQH9IzWoRBeUwatIk5pNfqUSSrXS+PsOM
I+ynCKtlAzWrsLw7iVGQ1fO9dk4cT87hxJd5bVj/Sf0+cUqYMyIEPn6YCBUrATxBU92RZNV7vUpr
ONxZYUL2zTL1WRbZ0+K1LLamisK6714ZKWLDNGHQC4WfKnhPMT8nt1pGp5g0A13xCsLWEsFqLYg4
QN1M2osXwhGoB5WJF6u7cf/UZuiEZx3rsWTFeKR757QOb7Tgg6WmE5cNozLpO2kad4beAqGQEqs9
NvgeFif1hEGSxhgGI1wS2HcxWkffDPc5EeDhWRSIsYRuYrIpOlub1BC/fP4lix0KWqoMXMZvTD/T
ifZrA0/a44NsO6/icCDeNEPrg4duy8lOc+zVNMtVLuZdoveTqS5i+mHSGhl5uYDEwd3ifb9IVgT0
tqwiPLjFeoMbLCrnJPv/kPMo7TW6bp0d9MRh0wzbdYFPPjzKCLdku2+mGYp42be0XnLxh8S6cJDx
NPf7IYoOiikka3TI0/36yl6KNwiTUU6Fkk1wFM6evb5NEWG+kRIl3FrE7yXZPeXxV7OSzOBQiAkL
5Jqqc804mk2SqdMXOJE6htl/RdL9Aklig8v8Erl3ESjOwCHHaWlYZ7nj4Wgp5ET12fpOEyOSBGIG
v9DPQh0EaDi5uHPB/6thhntEHgNlF9L68o+Svw9oWyudIRqoqRA1sUMyxpAuJhLLT+n7zMwIEtOr
5I9wOQb7ToKfT5SIapO5FvcmK0zWTRYBalFhnQsj8Hu9q/b9dwWVEQ25vtrOr5IAJgxheT0TOZPc
9pgaK26sIEbOUFX0/h7vZyBlFP8lBdZAZQ5vJjUeAgjewcCTmRVPkkpq61nzjgSTOoqXDjFA2WC1
dFt6jCFekEmLYxvkI0+iWjO1LfAB4VrNjwLLN5RPOfX0hn83jmzgSISRoS5vI0vHHybQCxhmKWUE
mjI5Wvz0v1ofweKcL08Uf/gDVGeklpnX5EK8EUPfCopGcW0oMM6YXHg3WECeA7NTKzWLT2/QmoI/
CDP2xP5RzZkm5jmSZqY1CzUdOGROe9OBBpLnsQ1d9j4MEipDzxS8stA+GT0Yy94JvJ+RSTH8DTqr
muU6hmzwlXOCa4tp0HlNrWHKTZNpD3PpeHwPFNE6jPewfehM0qMlp0eZKgjxHQxPBx6HR+jeQ9cd
Ko3MS5JSTK+71SJGNvVyTyLUGcTksydw/vHpoLpEQKjU5YVblxFV2BaUs8OLeXUDDHMHR7FRZula
q4H+xTCEtXspsk9dBjtveRBD9PaPMZxYUn0ogmSwHvQ7Mef3ONw4q2FlQ5c5nxa2kyNY1owhw8BV
OgpxdgZ130mVGhh3PO999FgU9B0Hn+yq/DxnliriXgJugM4dZpix6adhGYssuv8D0r6Hs+t1qu6y
ah8kUeanr5NSUcb0/TGquUq6sd7YcrMB3j0TRN9gg3DC0EC2tFBQrrpLLkJ92bAohE0ysK73i539
5kqYXcMAL8G8oNIJnyX9SQZvDCO3JV2t7J/4YTS7CoZ38n70w+GMWlKtJ289hVyTtRUiGqfCkKj6
uWpXRDgefw/SKDZfrUt0P3MoBf/3oUDhFe8AEUwwQ6zKKR16WWqDMU78tQ9yuvi0JYQtiMdSPOQ1
v4SL9uNEmvjXMhSqmwH4dexppU8qnwJhF0hBgxW8p49bemOVGSbXUccEJ3ORGlHjHzHi80pWWaD/
S28CjsHcvCGHzrO2qy6YTX6DJvAASlIbg9eP8mXnuASShSA7bn9016yBvDD0pOCWqpwyOzSy8JjR
ctgAs4+t8qmc0Ei0R4QGut82FTPTPq25X5aYrA3PAAFjndFVP5gvJmBvmmDiRlh6duqpCZBUKoK7
1bl+t39F7IeI4yI2QFKYPiWpXRUeGdjIDmIfAxBRaRXKFz2tUgx5D6HumK6mqKz5EzF7zww/V1Md
VfEoAERPyQxHpDfgSUq+9PCuxIVECZ0KkpJCqQgvOCQkciFBWAi8VQDplvYjMEsOoLPt85MVHzJ6
o23Nu948KVRxZnT+Zps5t3sSSHR2K/rKukC+7MP9UVFVYdGOdS1BZAfVK2TDVb8QpMxUueM5Fhsr
pmXqaUS19a6Y7hC1DliOKHkRJzoP5+yofmNiSjjRn4kOecKX5EM/vEgvw1g3FtRRMrZI7M63j0w4
h14R158+6gJOWtKALLD6Hmca6nLDx63mXCDwV9OWZB/P4RRCToFyvna84qv7aCPdTHhqZCk5Av9k
fLwQ/aK1sysgtrccMx0t7uskIexefQBdExHyjmmsJpE9hauQrRC8Q1JQh5UBntQZTGgFhyzU8wsL
x7DixxMTlpRSZ9ZB2cqd66w/A28yJ1HRsYJ440j/mYcwuQa98Wjb2wOuL492qtKWbIncheENef+8
mpgG4rVbuWwyi94SouSEfeeIX7nEvSmDo3PwCsuwm9wyqfgVCI7b0Ye//bHZ2oq4/xEggHGOUHJ6
TEFwwYXlOtxOSOePsXZ3eXEYNj1V7hfsemLBsfMR7RrC7llHe++SRS8sL7HWScpxS1jlJ7xhIgbg
H4a9P6qx8R15so+sDJjiUY9zXK9odqqhyPFCwxiGot30eJs2VKZufF/skYwCxuJuaNpzQ2rPbmcs
PAXiWE03gXIzR8H5Rpy0WigmZrVNMBdr2VViCkNvO7XaqjfF07fgBVnLOiB1xR5aqOaUbXqGUFq4
v6YQZcWTyMQdffaZuY9eXvBUarrqZGCnV9F8HV6PWEusNWrwjwmIRKBnoUdEuZ0XSsND+QxWeHlo
Yl2gbGujvwpsbUrQsfyUbxAKN74cEJFUYhoFGxL44SVDLcQNIs6Mv82UDLNQ2jj2fBbjOH213uje
2TF7HHQ70esuEirKd5Hfcjv3kejTQWViy+NZbkP3e63UcNe4teK5GyberCN5fTzZwktrnFtxhYSE
Z5WzL02w4Y5lSEFRSDDlupDiZpv8v9DvOj8TOeQcEiLqssssi61bjeZMQO2PoGm/j4ZadMpfvl5C
4jlvi+mFkeZUNM5oGZ1TofeXVFqktlBp9xSe8q3awIJc1NxkV3Sto6uJ3zQjIvs+nLlfRUQ1l+bh
v1PMPqCM7sl0Xw77wVAIYho8t/LR6Hbg6uJLA8NJvKSZgMfEyiFPI+YTseRDVbEXPJ6x86hf7/6Q
wf9AdrtVokgzC73M21QxhiF7m3P7skvJ6+tACUtTJsSsZ8hSfkWyUQx+QaQzlOaKmUsXXc+92TqM
QHRG8mdXC1HFMf9ptP6YSgZ0wPidTLCG2PndndE7VTsBKIHGoHyq3F1J/Rl+SN73z/iCs4SKoL/6
c3/Cw28uxdCvnQTpbmXgbntO0f4ijpVnOLkyvA1ybizvsRsm5F2bLEB1HSMTzPoGFto67A8FdUVI
frsC1YmeBhx8kq7LDvTaijQUDgT87kLAGG9OfBdImodLJz1xMTpzyDmf7faX2x8zbKvfPyJbgh7+
UUva3IhiBqtgnF4B3NisTigjDavkqLPHZWFisOix4poThk3orNMXJRpj1favfdB2bZMjBuDNhYTt
M31FBDGQwOUjUAP9cHyLGjvVxW+8PRMMSBkDOlVMmHQaWPk/yWr5cZogzPcAG4uGT7scSSRCtJR2
IqQx+gk9PRmcIcurGgKJfdyAQ43g+wiDef5kCHmUwxo4wnKBNwC00wfK4AKENDNsBdyKLrbk31MZ
Iqu1tZbks2NF8PELpL5ZX6weqmEaQCCOgl+0/BCUv1yw6yiIHBTmeD9dSyCPsY8xRtxv+C3zD0HR
5Ej5pGZYtpDhp4+O9ON/3txMU2LhG+urSO82Frwo69rw/EaDs84NYjwFWINzT9iV9eG6c8XSOqbQ
faLqZhMPJALYdNxdOMFtOPWsvoYk6RlCS9q5popOkm/tpq5E3WX+2RizDk6nIjRuZY1np2jRoY1f
ibei+WDz1HmxdfO5cyBmCP8ev648oT0Q52Ts+RlY/ZhKR8C0c9UdbEJ0VuTCr7v8s/1P53ImrNrL
XjpfC6IUzeYjheTKLdz/RoOuAt1hCuG/6j3qPLvKI+yubypO5dUAI8H0l6NsfCrLn/XtG5PhNnJX
hLuL/CqXITq2zlT8r1Xn9rncqJRcAR7IsiWZg+ihIaz/5uslVC5TGfqRl1mrd15zD7Iudh4sfStM
7Ui1NIhkEwFhB2U2V3b2MYbLsoGl7tbprpH60U0s2mIte4GHgTUbemTul2urd7dv4OrQMjEctPY5
zEgUPAJJYzSKGN90P+aeqJ7DzJreBgu4YM4bcZqjWBZNte297AEg3AoHfmn17TD3AXBarGZs2zKC
QWNbPc1B14QOVQdjvsfLiIoeAFu2ZlBPjestUavYofjRssQ0fl3G5jzMDEk12IuujcM/pGbLuI5R
KUXorg9O9b6qmB3pzqH7RYB+SabekAHFMB663JcNi/R73z3vm1VzacTte6JeJPoVAj2cf0NLQvs+
xUfh3oCGcMai0K6Fbnd6rbmfL30/LODHhn+DapC1zKWnlM8rjz+Ry9Gh2xzqq3tuy95RVjODmMYO
hYQhYq7zLKX6u1ci7/8Q14SPb7c/Cyy5TO4M4rJCsqo7pARjqoXjEfFFM08L0dcoR0OWBCMA9zi6
QtjN3NcZw155NIU1RDOBHnf2iGmo+4I2jn5OaYjeTQCYcncX4IRqywm0dJAg7J2Xr/Rjpn+n2Qxb
XkDzrwhZkTrIjS1HM38eMOfhJtK7SISAWDgXF3rgV8ZZvt1Zh8CdUVPTS0RHFKXvMVcBbwms41V7
gL8FDfaa1CDZuJ+8BrzkmlsnK9+XlHS5fS96okEsj3HrXloJfmnGHkewUuzLibTwtoadaFVa1dCn
v6aU0Y4Sr4FJMwzv2m0gku4KxBkuo2LU34ZW8LYFIkgnsWIl+XLL1AhEXFMxXWxk2ARBR13wxmgs
2IsB2OpnMt2vc8DljOmCbqQdFoV3xWqo/x7AhMGULGOoGEQz1CCSpKOYe2VpswiRQmZnmLZNygQK
DdIFVFCemoSJiXJLElP+QUn3aeP0j9Vek3MydZYgP40/Y9VbEKIjZ9KLnOFiUMWaroozFMYhCrEN
iDt5gWkT+7pr63P1r40NW+fpu71k/LeurrlJ4A75KDVUfTJ9N/SQjg+V7/7AKrOjX5gF1k3u/+Ud
+xYlzsfgPHRJ1rNs3vgvgvAL3ZHPpCS+uDAm4Y5xazH4PiDTmac6L1myGGeZzG7by4EP0agh349H
NC0CVBtm722JiEsE1vMjbkUrFTMs9dzc50E+z6U46F3xbDqWVAlNzqM/83lImqSlIBjZdnYEPCvE
WV9MDyZ+D6dPX944TSNnUH2jdBEXqV5hbwN7YCjxZ5b9WNmmbPONc4VXs5VhG//SSsH4FJD+M8iR
TH20ZYcFOQgHYd6brnfoePZq0+ONzZI1LAuySFaHqatU6vHkiHii6HkAH2FulktJA7a2xD7pPXnL
WVFNprmovJ3eW662J/xWE669XP8JDIZyidgee9OSEB0Y2e0M54/QTDskU+8B5BNrb2eYVjqoQyct
qpteTuMHgr8FKx7OUG1MPuWoFR/ISlc5pJTcgIMQZsObtVyReo1WyxaSVDsfC1moV1qdNYWGGHnT
AAAMt0lWuh7NzAGXirMMEgcIHU+BfSIVbpN9fbdNpoEkJwIcij/u5O++uVjI7BmLJV0kf7J5yKaD
e5O16HVTQuT7YDCYYqtohqmBOXgP1YKES0fLbFXUolXnwQ5CvlBu1Zfg9duBt33pcFroVQ79JszC
Rzx5T43+3fuZ3yB6w7JYUQJTXsgbrJGiBWFXNqroCh7AO2EMLi+m0iEB2jd2MlhTX69gaJHet/cT
/BTeLS3T0Ghu8i1eTjb+ihOE/sL34z8pPAku6eCEhYSL33sfIzPJLBDSKQZTKUT28+jhUi+rKuAY
AY8iTn/NGkzov0llr6ghKr3auy6Y1AAvUQMplP9hiul6uoJ9b7eaxqY+J+5mNok2hNXaN98CTOe2
qdVDP4DbCQQI3+0G7CrAKvqqpJZpSvMJ5v5HXA7hXSL47fZMrdM+Clx6EdTiQiqVk5cr6V44kMKl
c9KX/W6l7yZO6wIE0hsnsXDOYzsL5UaMRLDGBPtDwG1bKxv22jQQiNsvsO+yu0T2jM0vjn3ThgP5
QIOXjx4xjuQASrzmc/g0bkHwiGsRx7ncLhKF+/cO6Y9ZUlUzVQ/6xiuaFDCIi319MSWVLaxDxFKr
bLdu0GUlEEshsBKCYtcQNeU8gdNouVIj1MBYwqgOj3jGDzPx00OPcYE5bonzzMhrla+cdfiFEgXs
0AbopF3J83CF2fpHZ6g7dvDMWY5NXdww+mHYX9McmiNariwfUI1a62PXq0rsTCrlwfAoFYvfoWgu
e16ebpD91L9S30L0N8lbx+xqK2OydRuQLjMLrK9TZD2PT0MYDSi/eJXEdAmEv9WC1HL2H+wP7tFM
mP1EkO5EAhQFW+VDxM0ZqUcJV8Ut8x9Bv1zT32fJM8htnQAZTx9dqgLElq6Kitc22OhINRvnzuuo
JSL0qdmjuW9F6ULt7xz3kPaaxOvzNAgbQolDjOygetQMZxwc4MUhwMjU2KOXLY8bxdUUhnkufJl8
iV3R96g36+BUXsHqzVbzwFLOw0w4PQ+390oah0mtxqLbPI7UObBZs2l3Hz/GqHk/c6esHiZlr3KR
Kp7fJXY6Sb/UPluvQwtBh80HRly2BpoGn1WIAnxHqSvygnopLCc0J8QArQa/SMKEx11zpUKzjFpG
/YQnF8+eLEUMgv1uZIARr6HB90oiWue3mFB2EFxGWbo4NDXsPiWn6evHGCpHgtx3jO8H7+S3aTXv
EnUwqE78TzHaqnbY3lSvfZyH8gPOwUqjPqn4SDBJgQx8HN08MEu8+NRgYFtqmTgbZVTvSoV4KR0g
QtOWmZO3H2PGnaCBnrO7MjtimmceLptUSOkV7qnmNMU9XVo+QWnFKG1euWsOHtUGu/d04pggNAZj
eQGTpf5j5YdKtVy6Inh3gK+ifExRjF8wu2b/SYmaROFwASibpgbLaZ9sprteK12W+lmibpsKwV05
J+BbqR9xxXaJY95A43kmc0gm6rNRMZHSJbK0NqWvTEPVxIGlQX+E6ZX9cjQeYVsUAcx2kbGzAgpe
jSiCrJnOpjzWQVFMOrjjkFWOClV7adCQbNI/U9IBPAwSp9ZjIg23Mjr/CId0Bel54CpzRE/hqZPl
PjzzNS5Vxx0z7gV2lgM4MxPkXM8gbTinEYerLM0VHUGAhP7WlBQDSH3WGhWCZ+H3I9DuHmCJrjAr
wovITE065aQbBj4c0U1fyF7hMqZIXDzXihrWLtCea6LoeYCUCbK5fFS4l+IuQHnnKGMQ7/Mev7GV
uxN/42sv7A/rCa8cPg6mGZ/TkW8ReIOtVl5F/x4gmKIs8zXbCpDVnGjkO9KkVDyYWMlh0JQS2C63
y1b9z3ddgW8jsqgqG4eHk7Vz7xdzttUOdwXdhCTKEO64md5kFTG9m39zfjQkt28yVlcuHuCRvXSV
q6Yq1fPK7AZRmP82K2PNFmblQHS3Df8MUCFlpgzWriul7tj9Rwob6YfAA1TEVYl+B1VrujA1phhO
QMWc4i1p89a8PNjPnLH4pX5ju+L29cbsbKN1uoCsuFXU+XuF/Y6iNKUzdFzBrhQ+gaKDYxFNz275
PT0rPFuGN61oUehVXWc0aSV7vEDYG+DfVfn4e1PdylW627BrIbbJ2/rckVUqrkaPZFIoXTNJtOcd
eZsNOpYa6G2Bqxl85IQsJ38ZcUwMJXqbx3+H8y4TJSx9DfwOBpSf8ik78w6vZCTTJrw1nW2PzWyF
GE5QJuJcz25TiwMAf1oS1cyupZ7n/18sSBrJA08hkr6iUlwVTmTqX46cGBvF1lofrapBaMw70BNJ
sajz2Bj6hBMZWQ6RUyMrc8nkqkU5NIiCwpfBEG8y/q40y3CFHfZ/hs5sfx+ptTTo4Z6g8wAl7NWI
0CIC+IE8x70/HN27A4nypUcnRqzKvHfx58t6N3d4NoZ0Iych+NiftBdAicqykDmxbZDnMwfLo6ET
dqegzvj72dPxnHckfOs13ixCFPi3RBCKyUX3db8ObHOp7nzcsItzyOC6qOQHlprfO2EnvLpNsM4H
X8s5zljtlQGyw9IU7L+/VXgp7C/VOiINAn4joN1eszEzLJj3AqtSKMq3f9chE6cM2m49t0S3C6Kh
gfCSE5DPljf0H58oJyCDk65qogzg85jgzlG9dzmFioNmp05gTlNLmfRlPT8UX7hGBSCn3xoX5vjT
/7gFOvcRYBxW3HrzFtlJYkSGtP3YnVtGXJoDyq/Pmf/kv5/auhTtPF80d6TG0+JdDQD+dYAD/R3D
u40sZ7qjKAEn6q541MvXqs6ciQVEhM2hA3va4Eq1nWxp7nKeLNpTM0DLsacFbozyAQGktKwvCHv3
70btzlYYipjGYkm7i4ACCxKunLNcPMbZJ92MAc2zvgnT0+68q+rfK0oXtRH4SCedzyNx4mHy4td1
Pls8DsYEBcWOKnsBvWtyGwajuD3KZIvOE7e8bXEn+1ushepBgfSi2NiWTtBmSyd6pu/2dXFKkk68
B8//+ABKlOoh0qVyJ2uidqLsrGMGa3wXP0ToEu02YlB/RbbGSTlmoAdncqFJZc38H25Ft9IL1gxE
P3hbkoi7Nu191Hf11HS9ZltcwPh0M/RWz+HpR903vK8oBAADFV3XKG0BH5LWxUD5w5NnvRgZWb+n
e1VFzzwtx1+kztJUXi4vXmKu8yunARDvNWusQzU7kHdamBg4n++aBT7pf9TMi68mI8XDeObP+FCR
OphJOxPt5NrAD+Y/tQTQNCg/+LytOrb3s9rVjJgyUb1Iu8nUVMz1oNMw3xZYPFgXsjdfg5nxlqVg
o9tBeNdK8vGksgVIKm+rkbsh/eblnOJZ+4gtyq3lnyWq0nphmj6ctmjBeXa3MEwRxot6MnYFDClP
PIZzy9fvl8BzSuH9RRpQWUyipsk31nqfh38PKEdGalLiZcbBhHCWbTLZ2FOMRy7+Rq2Xpl+8euUW
6szZ2K++1ITznEELRZwP/P5/ljUCDzxTYf181uEcoVydzbhyuhBlENIr/FaYeuikHr0+Ms+KwLNG
sMUKGklLHOO7UQzMxIvKTMtl1EStd4TAoXGuvu6XpUhp8q6Nbs5gXyDakGufFvAVMXfGOTorYQp1
EeNJkuyUo8PiPDJSmtrPLHVL5H7BQwzfZvm6oC1WCA8Mp8HfVQANWLOyv3M35PXYSSjpxxY1on8T
daPdREh3X+lNZ+URYLpRonox9UJ/ogK7iroGJ1WHtT4H8QZUeGmxtMbE/SR6AFClgvcuBcXNeGCr
fvgxYK+wNvRAQF7dxF0EAf1NuuAHVqac57DwlWuFn8C6LWT+y1wJMFWNTqJO+8wGvou1MPq/15Yl
htrDUDrDrvEa573sKJ0XZ8VYljjUjxoXg2Woq33o639D4w5HIf0pwgf4mHnH5A61W48exC49LwX8
UQeZSWqDFH1muqp5ApuT09Wg4fKk4ih6j89IsBpsMjn49vmZRaBoN/+J2UdnemSrMERP5190K14g
2lxYTvMJZ8lh2ERwBoW9N0jAPEG1ZETli7GsGjmcVBLqIz+MyGUVYOVePPuDfff+aIBnqgo6gxJx
dAI2SDcRDymTFr4X6/ASTYFe6K/OEzHOSz+4SathQISuc+JLwB16hjk5WLstcUbv4YiWbNznyjJC
t1nuKfuRpSLHkxRnBxKfHXOCeCHDq1DDp1oOBu6rst0+l+4EG9Szp/q/2T3MbT9lG8htCQlWltq+
lq3apvmQev9BQdzsqB95SxE7MNGNBbLWTAHt3xUppDbrl8X/Ox3dCOBQRSLLk3rC6vvSZNLYevxe
WEWO1i3tCEsQXMWd4Nz0deIpNFhdC2r61HItxPaWVXHJcGuTtjeZxJ3vi1zlIfRfFwzsdHzND2gc
EMkkou3by+eaDwrDkgHzqnU7v922PFFaS2NZnGLjXnSFc7skydYTp+bqGebuOmHLVXAATd8p8jOA
wHHelEQdZOT8zr6/g1TZ4NDXEfULAR8SMkwEGEcTvXuz9b8P1GjgBoZRUieOG0xpBDtfI5clqxK7
aepkUTTEERojutuQ6l43+6jsWx+Es3W8Vc8wZOAqK0tm9DizFQ+rqwbrrmOV441Fdxmzdl/7hUPz
nooIvZ2A1x1vzdWTCV5qDKJ86c0o8qMuG9Q78CM13qlM6MuwolfPWWO9c9+g87kcR7brVSYoE7RZ
ss8nIE1M6LKZ8W2OI/Vt3jZOsZpQ1nVD/Ra6jEx2JEbMV9wOWVPCocZkfdduxr/nPWyhSjDckGKA
0p6nMzcARmNHMLLtnPzRIr67XyVtC5S8xIcHPCg1ZV2m11sm2meEbfiX9pXrQnEZbtLHEvAM77IS
8FYyCl2rz540Sxrji0RURWN4re7LdzIGs150CwS0ibu07gmWnisJ2YlKfckfNlWGW47m//gSkTRo
skl6+8rEq2tRlwRT4XGnrbB+Jbzlk+LnM3QIY+SeJY4vUujS2XhHRYWV35qVsKXTInZwY9OZ3SHp
ZbmxYWTb9V3tQuwhovLjSUnU4sbVmAyHshxj5hRmd1MTRUa2m1DSXwXX5p0eHnBOqaRJFFAn30Yi
YHQU9cihLJgwLxC88fg9JCMgIsJInDYLwUSlljIsm5Nmp7owjByK5y+FLqkqllIPOJIH+Fvoy/UE
UqbiGAB/Ex0qjHajOwc01UUs+PbLNvpBYwor+AODjrdBSjBeMd0Q54TRi0mrlOABtfHVyVuPyu/K
adHHSXKf5IzUl+Lt6L5NSDUYeUfoviwFtrahJeQ5E+F2+hLos8CfAJboD1YGM3OCEohrCo/HuodT
SryxjmrVkvlXGWeSLuTXIlDO96iuz9qXB76m8DguFomHkyEdVeoVDWIeL7Dm0hz2d+u4LFF+w6ec
f8qjPPNJ4n1w7a+QGOAw+ek48usT8mRP8LGZV1nFkEajmclxSBk4tiRx9xRf3HOhnKpevfCHSoBQ
qc7n/3U5nHHKxWzUPyfnT5j3HkhXHrfqSfj2EPpgoVltXKC7WYn7jN96KDag2FLvj2mRGHBJVRnx
aUj20/OgJk2gujVau7+QvLMWiU296RtRkihmrdYA82+l5bM2jWkk+KQLqC8N70hFqPNiiF/JijpB
j5NjfDAdHwGZCLjm/L3KyGBRr4+UD8OsK2AsbgpyQPTZsTkHH3kPoaOabzorxg/P1f+UZzerp3ox
eXOkG90LGxSkgHjg28+xKgGmk+IPAjl3aue+bL8JRRauWYZAjpwsu6CqaTCW50ajqGxDwIV23pMS
T6JciPBYV9Z2+HpkPcgImEj1hFa+RkSXa6k+EIv8YwuFRhZ7xg1iQymeyQ+H93AT46VaweQQOCnW
bzLVPmaO7sl1fDc/gNRNK0HXaiH+2TSoMt+doZitCikYMhRcX374I7hY1nhZdVXT6FHEJCTgPa1I
ZW6+HIG7Bqp/2bXWROLB4if7SjztzDu46bVPYwqmt33j4MBT3MufWmXVMVfFZr3CMID8IbtdMBb/
r99sLd2JLiI7OcVzIzyKHd/7NVL0CouJfGG8cW5iX9KwE5HaRAP5sdvlNBgnSE3vHDYsUunWVa4N
DRMHB/lMKlnlWXWGBG+LRqn6zrhyhH6SXekOishbPp19Egey51n38bp8JG4qQfIIWKPeUbLQ4+MM
AMd7MiWlip6Voc4Ct1xrnIzo3nwY+UmhNDCrjr/2I9lT+mLwbpxC8sofYNn7bVkEa3FuyEJLC1H5
pdBU4dBoeHhOW9Ua9+pGo101EerYfwXm+jNOV56IUwizpvpKkfxpfqX1Hdlqr8WKyHUbmb1nM31a
XrNyO2pk4SdXgika8w/DeOMW/P6OmkDhE8BUGYw4S2ilsU2qkfzTWBcasyhKGxDkPQjYUk5u4fWD
is01w8qoQahiG8pGU/qw9AMFabs7GsfrEbPBhaNN0MZZROXZAysrz0dVH5NIPqaV4+6jk6jUOvuI
NegksmZsNEUlnzrKplYYdjF4Y1RUO/1XRgbBzydzow41uLHzuIblDVzWcsMu6iMk/aWWl8mAgLBG
nQby9VlJyPcJ8ZVmAmA94f7QbX6YMZ3ab/GbgoWy7X93ro5ZbEAogEC/qmebSFLDJHaGfoV2xTjZ
bSG6Lfhbu8hrW/Gv+B4+mOAzN1oR6x8qfREGqtFqIC4pZzFv5KebyBC/8WLacejctSRYNCjR6SjM
EZ+eFrt7mHZZ3bYWJjtvFDDQfSVj5Ueq4F0Eq0vAgnoXm1WQ9FuYwzaBy/Li67iIn6lkvlZurzKO
VNoROy8aorbIIaNQU+G4nUGIh1CT+HngPI2bUPdRO2exAqHeknGv7GfJ2yaWd+F3OgYEF5u00wdN
kYIhbwE+frRZewVrTugFiT7+f6425N5PEyZ6IPKWfq5eAIKCErv+sgx5iH3k+etS3r+beRDs7OtB
AJ++PgfXD3SxH6YNNuQh81fwOXuwig1JPRElcSZpc4Ot+wOLKbDzGWGnF3fxUiq69Ot0xuswQX//
E6P87wJSCTz1v5LboXFiWIV3qZ0PfxzbK5+8Lup7GG/DbxGuYhjV7o4HXPYuUdU7dFZWY1BYxIEV
l7r5lM89d9cFdW+VICbh+4z7gr4sCrWPoP/R8WtunTfdOPnflcPMljPW5y4hUTcA4fNRRHBSavTX
H+K8C8dQcj9IwDRbpx2BCYWjSEXGlWHTOc3sX7O/N/hf7RS+//E+wTIV+NBWHFl5zIDEX7+iPdGg
DNaMNdqzFlbpOk2mvMjBUztitmxGgWxokOER/KwG2Hvb1uP3P265YsGSo55smXeWU8BNpvhhO2b3
LgW8VIdwhDht+hal24+vxEE/j4WDr0ruad5fDM9oGgL7zUiACVf7XJMbPTLOG/VFN6pqHpUaS6Ng
ag/AhJR5L4gShvz3xOeVBsoVx7XDfHPWw35zaTeWkNWIyQxvmU82DJuixJYndfG1d0ol4SmETdNw
g+emeeXVJ28FRpOsOiD9pI3hEyRaZPnWm7rLQefoKGfrbHWQRtV9NEq2/upRRjeHwUlt32P5fqP5
s1PGbYoNqBmSZ2Zhvvk1oRzbvEbIuGqmt5UaEaeNvcIDZvjM2bGATYCpqvriizlgPRaw88SlpWMf
MfksaTFbzcxWm7jAwhB9IZoR4d5tlNUChYFsDk90goYJ0QDYpSHf6kWNbKp6Z+oB/fODwoUvqgX2
dZptDKVB4yxyKTTeSKQxqLu5CKK2mB2ly/M54AcgIogpqy8/CEfyj1Fv1yexV9eH/iGwpF+YczjV
Io2+xmkQMWn495GoFdgHxA4jPU0eAfa/VGYSk4+Rnwq5wJ9FEcydOfxZgQUKSgIQ9fqasQkymlGu
cMQCS5gBonezCem4wV80x/8A49W1YzSrevIEQN56WXBzteNzyngHw42SWwrHdusSKcnIqINtI1Wn
MzmiRzWaQoKXovKUP8Sfr9Jjr5W4cD6yt0izHW7Va8ZKY5mCCsy9SrgLFfk+QusGgdRPwd256IxC
AF6QrG/v+JPHh3oznk82kiT7zD7gdJ591nXPh8bCFr/upPZIeYWSBm7Aa+disNpV4JPA+tjjKj4O
cbxc62Ajjt4DNoZeacIUk3GvkH4yTOiy1oyKS9qrrFZEkTvW56ZwhKm9KNDfSad6oVOoz8GlkftT
C2wX2nHEF/QKp2isqkTUKks0Sj91zanvGoN0AHNvJAqe7rw51+aUSDq6AHyj6vbZIQ8Wwd+Kx/7K
IYBtsDWdhhmAQ7HhDrQ5EN1Dx3hkjxP1Ahw3CxOKq8oS9DPolKJVWYm+sVMP3SVi5OhO6or/XV7J
015A+AayxRuqo91SO4GgEUytLrOjb5cjU3ieNcmVGcSyxIGZo++a9LeasQ3Mi8Jmp4cagX/bcci9
qZ4VamoZu8FDKmXg3sCu4sx6AIwewEurb0vvpOtpjQDILSYlDPbYDoRskkbmNYPC3zH3rW6n8jAm
eCKQsjDaPoURkTt/h4IulHKeEDEaOUxcpH+n509nPrqVsltrukYoIoM/xfLNWF7ab2TKdHvX3Rmq
Myr1H3WFmRrWqDqxkFjQSOnkCVg9hZJAchJm2puFTZIyiDx/bJdF3+uNSUyeI3jbRuaJs9HLKkX6
WWM45ppXJPi1UHGPF8e4YM8o2Y9hohSXAOWPFRJiB4/VDp+njq6fEcJh3awDxc6Xe6XRdydhtTR3
YWNol2WyN+rlKCBM1cgWquNpwjqIlItJm7Cw4+hHJ8koulc0D+LZ32vdfpdE64l57JEFi70SgCnc
2sfsMSuJ9G1EOmwYPUzJhI4Xow999fMr2vKRmxgM+IFGk00uSYONWUbgGD3FF3sRlueObeedvXZc
CAjcyVqq9CP7ccH74RY9M9Bt2jDW8WZIbP81SybRtz47joWCvpRBfG0XSl06NeC4xQEmUlT8yfWb
PwCTGP0KveycFquV/1QL6e1lhpWoA4ovQqhbn4sjn2nwASxt+qCiYeoW5zc88b2USiu4EMZd8FOs
Ce/Nm01+yjzlcveL3dktMEGPqLp0YO6FAuAjhuUa/7tgMKUvYOWD4SLMR9TBriiHkqt58Aqy8VHu
qwk8IM+veN1BOfoufo+dGzBNeV+JI+KFUWD1KKW+8IkRumx7ufw/thM46A4oRYQWN+QC9y4qy3dU
Pu6LHM+I3ziKIisnrT7Jq0ZStxidcfrWQrIYjgSfOfhp0D+XJWhBqcuKVlJUbol4iy4yv1s3UQdr
pWuXp+fQVIo39l7acFaddGcPXfswCeSZ71mmdesoj8QqCOOX5ya3kEv16aIjkKXfFGsOu4soeO+6
vuwf935BpdIgIl0yWIwPzb1v4asSoChyE5sv/pR3hD8pB8NA0m5Er//NVlg6Z3Aw159qxBPl+RtB
voGYbbIfSj14W+aMaK01Mukj1mv49RQr7fCnh9cqubHfR3+eOQKs7tyfsLynv//64QS5m6AaBtqX
b5lPozqF+zg8yhjkDkHyVEAK+1PlG9q3Z5xPKUedM6pDPORCJKJMCsuLhj5o/dt6WDMnyVi8/Ic3
IM2ctw6mKzpkPcn9XUUJAappS7gsdNarPhuJsI66iBhJN8Hd71l5On7aZwPE6Hz1LlaZZp+p/TrI
aFDvvdjz0ktyBPFnjlHtFjqaUYQWnF0rv8++DHy+z4z+ZmOgSfAlPf1rgcTCvgWE3FKAripQ1GLy
8mefjvfWDNtruAppSyQJwqjv9JXSZQthghvM9BkUC1aqGB5Zkya0g8Pw1QO76S91yArAySm8aUut
cQB8daNg7FF6LpV7BAees/1kIPc95mtNqROdXdNxMMXd+SPrMLvYXNancMPu0+g/tD9dKojhITuw
+LXCwk5r7Afm+MJP/e8SSsPxCA27hShRlYHRAGb0ceVhi95Y8md6DLZlXYoJAo7LWUSvAXkSWoqu
K/Nyu/JWUoJmmVIIw2BzORiPtFJVUoDnpKTDDVJzvqL4Hz9UoQESXkILP3howUKE/FKVPhXeEYdr
U70GkmQ8RhyqCO0qnoFRnt2j9THT/+rbKI0S6Ji3AJcbplFa2bcxiLLtEVLi21/BLeoaTJKxXZII
D9J5r424XWJuEhsKc6KmmEBEDWL7jtG/3yz+IIfYulJm9umRwPYg9V8v9+/PK3Bg6wZl1XPBQKJs
BUy/UALtBLwAXEWg7iwaRN71p/a5K6S97+fRhy+XdNej9x+Kh9nE8l1AJ+wAAoLH5sGOzolKkYPj
gH9l/BGezrT2OynCrThzLDK0kYQN+Nbgb3OIZgzipo0IBJpUroSbkzRJNSOOtGYKQwWWSSuejRg7
w27pTGAF08gMMl5t+go1J8PdhQbGGaemFXJ43ijrnzV3ECWQ8AOaoR0+G+vrEJ/4zKpbwNfZW3t0
pWvSRrnivaS5eA2nxfZyDEWW69BnnNoVlvnzjSKu+i9bd93SDFDXUZb+OIH4n3i5uDqjlAiX1QoJ
48QWHBVHPooaMHGY29QOq0nl9nAXichbr29cQBSkon74o4E6XYZ2VJZgeTABrCDM2TzA+zQ8OWzs
hq3iCLwYX+fO+f8rlXGdgm2qQcE5Orq5VVI05gnija83cNkoxcIDtEDlb4X1h3oelysD15MsA4fI
r86px4kNsOf6YraO8KSnBplD1SjmsIm95DewbNMGXeFx9dKVqwx13G/OSuXYeLsJBAOlu0t6HpX2
2/UIc8H4o8LAY43FIH8FfDNzHSplHPIjlNxAJab9rVU7KQOXJimlZ7l7UZwUGqyTQvCMbdNiIta8
bJsB3ndD466tjf7erkVDLyOpVXK+53jZGvAJ7V7LCyqFXx/+OWBkcTHDYbchcY2hx5YoRhHIAHA+
bKxwQUJjQ5/xutA9oX1glrwY3O/g8e/67IAIE/s/eCmUW3apyjxxEWWhe9XacwclejFFE6H7R80y
rm/1cB3n7OGZPf7DVMUxTFoUX/UTdmvIhj3jaftUolA7OaduK+elxgdWtKynKvJ8fNuNXe7mCpCD
TX2/aczwD8L25EItH9obOYlXSqZNuxf/dByYJZOVs/W2gZSZJGbVQaYQTL/Ho8ntHFOSg+kj7wD6
+10RuNdn8ETg3Auo7AF0Ya7xaOQKVHNvTFRkIm1g+SJwFS/QO73Du/nCOcFjAzb2an0jJuxDkzD3
iV5+6MjN6G66n4sIdU3JIYQRvfvNZNlMyQAzz5B4X191Tr1m3VIF8qsXsR4CGfwsvZyW2o2VWwZY
/sd210NasmuKVGeWdpTpocHGpcz/X7uPLCx/3YWfHzzM1ygh+HZex6Mfg4O54kvcIV2hlXSwmpSd
IB++ZECNhP2DmziGAIbXA8bAPid3cxHuhAisJGzRPMO8MtYogGN9/tm8X0HHYyRoyTGuCgQSgYaa
iFdU8h1Xm9nNGFESBpCrzsXM4l09k2S54O//AV8GBaprs7G6+9cW/wnSCazaByAzzVWFiUdkcV/Z
RkhyUdbFF6zCELojH26Vlh4Q3pZbS0WAokT/pHW9ScjUOKDqdKiULsnWuWypAKh9mo6fwLocWqfp
UBJixvVUxug2KZBnU4adT2OqVKkKCHMuHw9pQmcpc2Iqs7y9rO7zElrrWQqWTqY3+oC4R3L7u5mX
7FFDucFTl7ilELgNSxgPhs/OcRGlA1JiatRAs/ZCJ7Mo1eSYDUT0JgC34PUx0TymvUeqT9sQpdaS
GfeOKvhKtV4p6pcfh4yMt4AtXVzfQyd7LGvdR4M90sYgTpuTco1UQMXk0Chxf3ya9O5IWrMKDUtS
0FPqhBxLbAVC9b89cYsY0qfFtodlbtQNysVQsnVNunv4cjkWXUhnToMcdh7o0VvKAxSo50qnluTS
yavl0fZo0n7KQVnpm7TafZTyNkW9oRzWbyeURY2ghzivCJO2xngYBrTAANiDGrNL3bxCEFTytuY8
A9b6LHQLPm70wKNFEg1sRokrLlGy5ZMPyHZm1XRc+RPDyoUcl3DRxr3NS/SKeQ/Hgs7FSXhH66fr
A3F9OC7ZEFqY4glDMgNtUltWrDy+arS4sUeniESG0sCPRYCuWMg5CoFZqozLi27uMV8r+ZRMmwBq
rapTGbG/2QZ3IMzZCn8/YA77tawLuMNTQzJO0nmTjpRzanPwH/l95tYiBP+Hnbgd/PkvRWshAeUp
q4v+4CSUlb+owoRLFbYWij8DsgD50bD6YVwhNTRPnE/tpcoZBuFl0NjyTDarPb3V6BGHrvAaqSUz
QT9+YYEjU1Y27wNvMoq0rAoAgHn8+Ch/D5DaLF9BkM+riMZfKdyZ6jfiPfn3lB1mv7grqP6FRByx
H3YphvkIx67PK7d9Hkv7LAF1VJVmTO9PF7pg0iR2TCTNzIJAthNzyjHI54m2w4yd+ACdqe5N9zem
WBgaKKS7NhYy19Xvp8bR9PZXtIL1NWAGYkZFxkjF8WsKzXLySsx+mHciRiV7iGGgIUlmRfS27zqO
jRrO3ONuwyGtcxdmSbo+quJMs4fQstYBHFLkyPiMXIVVFUUhOX3B6rSS9ysGtUpkvGKgQ1hvIrSf
gHHXtk5vneqAAehe2ACSUAfdJcZy3Jm+88MoptuGC9n07D0GB9yz4MXbxa9YzO97WpKvROR8G5Yg
YC1iYD/MCRxi0I4Coa2JB0V4m6b3ahSbkVrjsu7yBV8byzP7jbDuSVXLfEqFR6IurO6+pl22v5up
tvi431wsHIdkhT372pg5St/bAMeqeqjm8I0V7ymzVk/mE5gzvcfpWeWxMYREiMqbnGresB5cXbvB
80Rdwm02NGfktlf5TeAsIallsfJz3IBXu44VfhJx8c8WkyTd4eU79cwNDrlIgXVc2bosiF4B3NOf
OQpRLlj8wRshWFOt2rIy7PZrqR56bTBDrcZqsfDfX2XfVa/pDYUdJx4KQTfuafKOc9TgZShjYP0H
3XXytKBmInfrv9ixxhGlBp1CsbOaq913kbsbR7NtQfeIV7qIxts6kf3JLcZb1QB7mci6ccGsTWO1
FW4y0thQxXBtn+lY57iq0lME7I44W0qWOgjtpbpAsnSAoNYGkGCcTPsjttmSvarIqJsm8YbGGrGy
Ks4gg5xHURR1udDBYY4OVHHfqjtwDswqqK6ZgEgEHph1MBIasbVqwcgR6BRgMrngyGqsuGl8uTxh
31WxBwv0mNnsz4TJgMMjjHC3J+E7uAav3rUednEQnwjgpaK3HF734KaN4NH+w4JAwhWK7PUwMFGK
naI2/NHPny5SZOXAYRIosXlGZ3p4paRrHnH06PGPnNljQVZjPHbe3XDtHuF/dJCOHyaY2OVkACLT
6RkH7mIW8R+Sh7vCBlG+Cqe5pK1p2/I7l3tRWcZsfhKyBOtGDC18SPGPp7ix3BfTOFOjtfjSzJTO
I1ClbGZIYlmzORO5IQ9WswwyRIf0ZHcACkJMcVYDOsZRbQl137dazf+XuRSDFr+MnScc99kcldeH
WxCg1rnq+wgYxmKGwzizXgBvcpMeYKOUbLewbLFS+7c9vvYLPXF1PvSO/XhuCG9lIZeyP866ru5c
NPBJ1Y5ZVX1bb2Y+NHuxerBsSiVjjqeX8tcg/CI0TrrqbxSatVxtp/J0cgzoqhGUrC82H8YQhBf+
JrRvtDfgFn7f5AUYot+gET1TCl31gzQJyT0d266pRK0j3IaDS4LlCycVQDV1k/PzwkWBGpvKtcbi
7EDhf4+/HRcZipx/zHzSbODgoX9PZEWFXsWQdrASzboMwsc7tVuepiS3j+2U/xy7xmZ/amemu2Jk
rDbSA/MIKNvWHuGQD9dTxgl6cv3rd8Rz32hNqjJPAzZQRCweIK/YfkrZOqjmm6IkKp3Z4Y6eath4
83xE2T9VUnxKzLYIaCXv61jTpQagk8XRqXpPZ06GzJ748MHlT6sRp1WdrVWG7dOLgywgIY1O8j3X
lVtWoagdoCZDOuqGdY22J5lfZjeHFblp4hleM3zurKFRT/v79Q7wI+Qinu0h0hIom6MNXzOCCGkq
bnFfjTykVFZReN6rONiNX+op5IpXkrfsp1y8UsXWwyXGhMqBFkFMLtsEN2E0ozvCZuMzUMZ4BoiR
j0KlByC/VaK5y3fJ5YtZq/cDZzaVp2VFPDvNjpSCQEdu/WN4ib0P0Y53HXv7TpWMCvgD35aUYSSo
ZDQWusaV+sYkq+tph7hrv9mALWwBESFpWBh1Dlz/fFVCG+ZJCdDMYzzDV1QL4CDPhgQTJLMGLS45
3o8AbPJSkATTKnQwIrMuM1Pdr8JICKjVHED8pXc4QxevjU+mmcmTJ+BcwFHxqPyeRDbKjXtCd1nR
sMlN4mDAGR50EDsfXS4D02SQvYAJd5veKVh9j7peIQY+00HXrAel2x+UzoCrZttG0/hEaZepXQ4r
MlotjPw5d477wgUxx6Z3IJX238X5GZ26fsNZVWvE+uo/A0ovW/UfvBConT9eDj9D2XObPrjMTznd
PtPmyIEi5/Qq/Fbif5VUDH1L4jUXAQCiGfqEJKbvTmRUO3zvk1i+VkA15D83aA5jCkp3+fywI0hZ
SD5P2sioT7yKYhX1dl95atMKS4gETDnEzc88XeQ2fMb162aet8tHCiWDAcCoDZGqrl18JlZjOb0O
fJxhMq1pXbuQd4JQKBN06007ek0dNHDj8N0SZIJsPN7bG2cav57oB6gIOsn2dgiSNvEXqfPvUaMr
fIfbIWB4AGwAE1DuTFxdYvqyQZdvAek+VJDNwIh/fm78V/IxpGb0/af75oudv+dV2boDNK8oY4Ba
4AObCp7j1+7G9bc6VjDaOD/Y+gBJbqyhTNwt7RWHfawvYuCb7Zkb0F15AhbTESy1GZmyuYlc+Q+S
OcO0xm7iLyUm0YxrjuznYXE3dZaM3rY3B8FezKUGdMfqmoGpmZdjm2qtZANF7LryzMXDz39tE8fq
N1yJr//ZVhkC81WkYZGp5XM0dielr+Ubvk6/ylLQmuUjslRgc/i7LB5VUuNLRX+RK5HIemkHzYDv
J/S5IdAdOTVAEU53iio6YbnfgThjxf51wL35QzeuGig/EhdbRf3ucsPBrbgKVlzD1G3dDCTdUgrg
H7kLBiQyWXy2AJ82whlQu8n9vkJTzOYhCki0mocCcfv0KnORVXt+co6rQZyf6R7SKSbZmFZBLuWc
jVAyHfFEA9GvsZHYXu62y4/RGoubZdcP9wxq9SV2UNWkTYmpOB9Gb6YR3LoWaPVbFSGVigbR6k8F
M5951WrgOBg8Z6KY/P/LlUFvAqC2a7oGXGsqqi5RsuocJrVwCm5TzsQQAt+Dts2OJoA2fXL1be3W
790YwpbAtWPb5JLgxL66lfXDF+vBkN6q6I4BXzjFKgKxykSD+AFf7G1ZJU03kLErnv/+ybry6PLv
IDMfGpzaMskE2JxkvyqmZeMF4PYZplgXpI2u3Xc/MhLS2ksUQovdPJZ2+/AeUj5krouKpEZhMvUh
uvQ7EvpY+whN6hIAGbHAveNz2+5N3N5gCCpjlKDaqTD1e6sqoYtdo1aqq2uu8Ek6Kn7MUy+b6BBt
rSKipuxksLl0cVWqM2E/+D4N26BnyxQaMGXanKkRBnHNIL3PUK93hPIZPY+Lf4DOFMp4svMuH1ua
R4XvQfK7Y40Odk36Nq/ybjpB0tz70jtuQJf+o0nVHlO6WRkfad2EamjxBfI1mqpIWkDICOvP7sOe
/F3Ym29XGnoLfjDfByFCsQt1D9Z+YpD6FZjj17/T1S08jxFanKkG/dVu1XAafEq+Rfz6QOVUjCDA
WKfhppEe+Wadehrd63CyaHOWascjsdIFY7s+OuqysmOpECnFJ0iSTwihtN6Mw9H24Bq9YSUp1eDG
IV0b2bPooW0ovqgRmXfAPL4tI776ZOkVkcS1tOyZc/36IAJI20zS6xqlsO7S3O2zpa/KMjIRTP/Y
RCBUDSKyL/Wm0Eey4+nxQoCDwtofel46hgQzlKbpaO6PovtbPM6uKTrF4z1WFru+1HN7UsKZ+Dpd
ysIiQC3u6et3AXgXCWzD4whlCNSbjpIsRY0CcrSW5G3Q8I//RLUgIKoSynBKmKJOh2cvnku9bMUx
AhW7SU3IkdTJB+F5UCo5mJikKt+gdqI5iaxyXkISSouAehYM3zo22Awemu/1EhzNlQ+bLG1YvT0o
z/ZJdNQjw6ucsDeHsXajVudJflGghq3mSgs3CpMSW34tYsmFb+xTZ2mtnvam/qaZ+tXu+WpGgwkW
Dr/nyx8jQslrim3i8IfdtN7/mkl45+ieY/FiOj03ysspitZWaG1zGohR4svQd4dK56sgHgXSpT8E
qnsVBwIvBDEr2H0n6VOACnPPWDlzClUK3NcI/Kp8dbONEzRa/W9ZV2/8NWdd6QdAIBDLf0oSHsgQ
zqsf7akmka2mhXNIDMRwTk4JvHVyic4sWXvsr4PLmp1aTZOzwqUv0oiBak7RRFElEgzxpp5YrXMe
C9aMMYdR35xnnFRCLOGHIJazGD5/fn1CcviYQM9nG8fzj5QLV0VEPQGECfTwDcrlp7PGYHXCd+X/
t1MPXkbefBYVFoafFI9G5QhYKSrbtvAe6/+znqbybb/q+DZaYkEAR87tIAuEU3kRaHr1JBR/gDNd
yHXwo0lkzqzRbaY2UDXWInf//4iuhu69kYdZyznLpShjd7Kx2LaLbNKhQdJexX1xGQxTO3/LSzvn
iV/w+TyYmurayXZVibi6jz7FJjkED6x0Kv8Yn9RrFcogQ2VuadpaFjeWipE3/PW5q2f0ZuzI4Rpy
XKTElEta6L94sZwb6iPTCR423FEfmut9qac7hq8bdICxtlMXAcdsOvpkPOQvBTSgJi41wEXm4N8S
P1X2KzV8nhEDGyeU5JvI/uxBX1JOdlSTqPX8uWZPCMU1K+8KM+eM+NuT5WgeHc8XBj8DYXjDnWNw
8qHaubUklaaemmhXjy3tp99lVgryVMCu6pEzzHUIimc75zsF826u8IbDzmzefqJb9tZNYEgTO3xF
8ERFItS19J1gsh5vg6YCgXFR8Jj35mf+bvOdr+6pUM08Y8qsUILyoljTyhmi8vh3ja7XojvkMjOm
zWEaFK/MChD6ir6Nq/szWLSqx6e/4N6sWGt8gyWK6guajNgTRdYcQZBGQlEJlni7GdOElcPHDR1h
v6B12MmcVAVhptHzHTOkbC/RduK8krdo9XfHof7QxPwyqQ1fxygxxFdUnNT61EPxTgMeOpmkpUQG
0PDmr8YROPAabnEnu59TkZVPgD5jJSeVDewl8HNsFVq8acNMyRbEZOdVjLZkHc337/UEL2qBDV9s
j6Rzfcefu0kwNICjbNp+wKQVh5nR77EanLqqk+P4SFVDyKV/uSI68QmdQ9svaJTSTurOdxsWjjuw
yWNa9LDhVr3KpN/RynP9ihMdL9Znj+BKnb5NSb04OlV2LjyYXQirWdXKz02Sbz6OVcHQ9p31jVgc
Vyp61g3JQv0tYbZqRJ543l5Jcu/6P9iQdjzqrw5b6ex9PZ7NCRx2kKLLGhw5Gqtd4R8kwH/jLSpa
Fqj0XlWiQaH8/TP6gDDvsh4/BNZUgBA5Y9bleLOTctfwDSiclKTdtiepwD79LsnyDdvjxwt/oZq8
6o/A+EZRi5YcAyPBOpSukBBtCexBtrntuMMVF/pgAFXMnJNDikOT8+3Awf5mvQcAaZP7nIiEpuDG
0wrVUlE9lW6LAsMZ1e3TV8oSLtQ7hzn6q8GICHeU0alzGwfaQCXhlc/+W1GH6vTYwozQNSpkMkAG
SV79566StupacxmdY9CF7CtaN7afBd0quX7wux11M3+oa2HofFZVlMmL5rYeIU4wT6tZdXWhr55m
9lpSFBswq0G5y2/1hqQKBhTuhqd6mBZLPqa4HtDVsUiaTPxoqQlo0frEQr8MFunjB28Cqh9uQ/yv
/XnZC9t3Evadd65DJdTSvOU4cT8/sSC35PjYDirIokO2XXxn33I/WKMixE9tM326j90lvBc90eeB
Xr+bD9fLrPGzus128s/dAj6o0VkQPGDgjAJk415UcPC3mbDJq7+FBtJVvjhV+95JLAHtN9us+cTt
9TJdFVdqxW6VumpGQOttAP4+D5Ga0qT5Dao/4onhl8gToDTyhAryR/tcPrph56jLRMWtStrFtR45
Qnir2eXOZRa/SmTUWh+xBIC/H27nzW83D8mMNlQG/JScPxPvMHRGz0U1mc6B0JaC5OiNzDpnp4Jp
oBqG6PfRYLgtHD/eaYQr9UPB5tWw1KZuc2jfoE2hnFC3MWT/eD8bzdGrYn8F1vV87HlqgFG98GNT
WXhjZctAVmLa7qDzWJO2PSyEyxHgaJD5PYEHilknIP2fyLOtmhlWdBdXgpkL2Z2WynbJMExBuWFN
5yNPNxVLN24la95cNujTdfuVa3BC9NOxU3xVCrOCnsuvnbFionaTQ1sYI1WINMXv3kRTXILO4jcl
3dvnhoPouxEEnZ+2iAG1/pYV1vkri9pAcUUzAZihc37QkyP6AhhQLRttd9rGds62hHb/3APES0Ga
QpkFgDgjzNdCWYYYChz5md76gE8GFsXn1bOY/t5ZgFLynnOD84CXmTXBwrY1lgnR0CwgfkuOpFKI
Trd+9/v1s+m1CHdYiY9ZNCH4lxN/Tk3v/EEy4t8Ftgysv3U/ciVNnyGkpJBnK4+RwX9eEOIywKCd
lARItxNj9LuqLQQ0xB4xq+F9Zz8frpaxkgRpRNNGA/8tFnOuO0KVET3OljFWx7d/o5Zo1CXYqRwv
M4cMif9kvkrLnn0czmUr2zgVld/eY4R5FywW7WUOoSul7uA5yDF/H3NnYa44frpDd01aJxl54suT
JZaIr1SgG18gf7bskzw/JejE5XUt2Atghu6HZAzlGRsHEx9nUrvsht6mBB15k2Zglacq+FptdkDr
EYwdfZf09Wk/DVFT/L2OKhDnAXFT355GsnW5LQaAgAo30OHlRqqXdwdC/1s0RhabJsyFMNx9jqJk
SkDfbdz4JG87CYopggyutrkqL5tkGUz6fW2B0sRuE9dsu59gJx57YjWb2VpR+wj7IyQ4LS8KqnmG
zgEGaCRGVr0Gaqnar7pInU10ApUIG5CykC1UBGxg7wx1pNK8tnFB1OxEjBEcm75govOoZGAgihFn
+eJXHxt38Uk9kJP9DFJR7cEWmZnnOmSYyUa0LFx42EcvZEVu6NnFCtcaVWE4LWHvVoSL0YPhWvp2
QDGl34vok+bRv21ZCnojmiEaDjpGnMYNPLcIzEX9LQCNU+v7DL/ZtykJtMH/bNrHx6D58n4wJwfC
xKt/1vg9CteBQv3rtWH7uXvSq27RjADHRQEk5kDhuNFx7as4rLq/V8ZEEJeSMcQYOOvzppwvIVO9
Fjo/7AR6qvDxd7dKMA9XjbP6SvWbsZmaSbws12n+uGZp6njfRf2h10YHdxd2b4AM55w5F4vp0mmL
DGGO3IGF056n1DONMdbTodG06ECZYJfWluIpi/bKAS477AIrPY7mBfgTG4Li9ceS3ZHfL96zCFnj
IZ9b8ZovdnXIfaVbh0PRgJecUIxDddleuH79mpsPYL/7ebC6DXJyLkbgwnHuFCq+C8AOT79MSja9
5ghO3aNGd711TcIMWCxPbD6LqumBF27yWuOH9gtD3M/QL/12G5MT8RoiX0K9XSvrj+7rZ3RmkoNQ
80fgIv0eqGUs73SIR1dihmLxFANNK8eoBKwueSbXb1X+NE9nOjr43n9EWMNYXbiA/1wCcB40oak2
sWQ0sEOBVZf8NHer5QesNY0NOu1Y6ghaunw+rWl3HAEKae3tB+yAa+1XHadLOtISmOaquXFZcCrU
GFtZW6nJaJIIPgm2F7TmU914z2xAeFQUdtBA/ZxPWlKU5p1E1MRYTJDjpagl0opVEosUx1Gyq2mP
wtwoydXjX/JBCbbdK+GQYEMtHYcfcQZXVUWAS+90yry4O/3vMwIUZynHHV+zMrDMgCsRqyBDbnCF
zrMGoSiNZfhsXNJQ2nvUXoaNW7J7gYj8wMl30mm/iCWegoKZXPqi6f2QsgsG3kf0Omp4UERtCtKU
WZ0jWKHTMQSy9PNr++kCdrPykm62lhsy71IBaDxIIDzAiSIXo9UmHNm6/xcD8Sq/h4ZoH6NH8VmP
daw+Uae9mifNvtF0eO0fO4KpT+///mpYPDtj/NOEuBBCUqln/nmr8qlvURccLp1QGZ5VFP38PK22
UagC4jSlqEwwWxFBZEmP1BBp4AAZ2xZEFuPNGRvh9+xXJjMKFA+MGXAlDucI8TKmnqiranJNxk0C
OWz1uOwPUeFK3OsrTptviP88J1mjwmjDMNn9z/OJK7Sthr1YHe+74RO2/J3NgUn25CYLsOrqVP7J
J6bBli4OpF9h0pKwXhr+iP8P5cKVtj2lwFOQXHzXdqbTCcC+/JO688m9kNVLK9vnP8ZYy+6yzBSe
WX2WI3rhANrSMVUFgZR7SXy+lXQZCnbMFNwRHrtqrRl9fS4us6f0mxqJLtduavsdLW2ASp1hif5H
xE7NIzSSSesJlKaZl5WKx6HwFRAyFCWgq24Jvp9CXpSSM8mrpJD7m/5vufBwWJX8eWOt3nGLrF+b
cK4bybo4BeDAS6RbpdoRZUTVpgSao5Z+7Hj1vtBc/QqBmM6y5znN/QMLZ2oDjsAQKnSwxy/3RwyR
F9z5BKhUbReLkGoGSNoSfclcyD8G31aBPF0ESH23Mv3wJvpVeISlpgJJXltto41p/pcCbkXbabPF
OLww1Kntd/ppWq19JtVObqYsrWzj0GC2j4OGewU+be7c9y5ThTZaCEeTmnuVLkzs5B8tMLUnV33h
hcZhK2YqcJFNbv/WccJpT3TuziQC8TjYokt8/373lr4+XZy+tb/IjfG0XRwqL+DZCuklwmqS2Sbc
HftK9AGeqmQqruCZg8472JoPOqCnJ9A+qO02Xb7zVzX31x1xXd7QpW7biOQaJBcZheVzMCAiPyQK
AGCtTgFlp8WNq6EZSyU2TaDl7sI41Za6As31No3urNXFTaZxrA6h9n6N4qbZcTr1l4O84uq/8sgQ
Am3+xIYwZWE+L/een/xqa8pCeodnT+fYwN6MLyYJX8rKvoPF6E2KLYA1GI/091SMztF0QJLjtShJ
FE1uo1/ughXzXRjzm3a8pxNwm81rWNzRQtYFYLAvuJE5WhAmEOjQsuSj2Y0MMff2f8Prusaz+DpF
9PE6/FPZ+mAHGZ6YpShgPbQpVyyTUFRd9czvDqqlsvGgYEibjVQSKRz+C7EXoKzioirgXO2FSGML
zenlfhjOImazJw+ce8Zdy0161diUl00FqbgEV/PszlhFkLLeujqM01zRTR2NpbvsWXlZy8mLC58x
0nzUmyt+WQ9gVga1wV86zaid2hnB1jVTAoEV/t35USEAYmJb211OcFCHa51i0JHkxAugChBf3Jai
X764OSowhPJnpcqYS5/l9h4F/15oHyG+d1ll7J5aA9jPGUbmjYZEBxP18OlmtD185rBx3mA4/ld5
wcBQ+CAQ5mpK0eG6l0H+AsqA9iwm1nbtYj2ATOEEK1azCkeAJvOypVCHtXP+mVV6BaHuTESis4Sf
aQDranekShAKHdQt9bWJ2l0tMmmeSotMniKxX1gUMMFKGArEFiVZ9O+fNut9h8eRDBB/xsaKKuVg
pJn4zjwt/QGRUYPF4DXqActZZhPWNsDDyOii9bPtbPLmAuGalEMgAeyQ8sBwLgiDfQAJvu5JtP5Y
sVdzVTcDTwXZOpNjQkFKvNwpYGLn7A6ZHfVg5q8pz+2TEsLtsQSnZefjJj4C1NPlp8oqhkPatvQ0
h6wgEMpWsmcQzeLuyz5+MM8OcX7oCEOPwU++Qo9AG2XJppUVyFd3Y/PwezaFmrzlN6FSU2VF04y4
Vnb2t2nTYSxTNSCJv5Gj+efEDEG4fVXR++18GFBCHXbrY9h5xjlQVdBTt8X0qtfekrKUx8N+psHa
c09gGtj2JraiKofYXq08/Zt5TiqkZF47vZPbj8hOZCIDnCayGWTHfPvu8KxPCjq2frWSMEENvNbP
zwRP6G2/adSgWUO6m9hlZ5wZmuCiFeprOJ8ITd7VihjFkIPxJwYw6aCgN4HvG9zNBzXX+9PGKI5Q
9+7S8YdbJWSf7eHWdpZ4udWsTv8vyPPjxxtYo4GkOyNL+BoIAL1HX5gNowYB1scZ8/p7N9loVua5
KFH8vhE9N4qydBPoamyO9TYY1pQMxF/Ab69vAe4srjhEOPrnaa0GQ9Yf2YU8CO5pQuW1f3raMBvF
iGbmqEsYlP/9txL316ZN+1/Dvt6SalgoTjQ8IU/JC8dQMGLpYFh27dQUw8tjkhBlG8Qqdf93Q+NK
wXlD/MHO4zo4i2Efuo+HP8LhVGVsQoZnceMyQvP1Yt1aNSMTTU0JwKV5ICv+EdAuRe6UYmgpx8w9
/zSd+/W+hyYsSozUyMwJet43v1wRhyLn0Txb+ApDfN/IYtF019wqUeU9Uv8kbBKT7gmYiZxgBuAH
hFgTyLMrIT1H1ALUQ9xzeoBxiTXNqx0AaDASvB5duSa+fqsFLn1xI1YjFE4pZW1B4AI4t+CGh5v5
rbuC8CbMHU9GNgom6ekvnZlE/v/XI32i80EeOUAmGIbtMgiZKNWGsaP1q5LOXWBxRJ/dbSzOGEAy
HAhzqtbGY2HIJeAQmnWgKWzm+dUCex5XMkz0AOXSFLKJjnjUHtoocm0QFsBKqJ1tQAYQmoPpMJ1r
7VZa4CXKC34WwyGFT52/ydSZIp0nLDPdpXdoZfV1dIfTQoox+rMblcFbtDJUfec92YE/caKqIqkj
cXLJsHpiQCRM9XlG5I2R7xf6E1yqMvOHR6v2FJOM53mGx5U25rTIwmLGiSwH8i92hhd4hznxUvft
BEE9luQFtkFY1NwoATAlDskdaErwlJAWvkukPmVWAEyCMXIfqG9Rz2TV/tOvf+Tj2CFvYbI9JbO4
xfjyLiE7Nk6gvuQaTV7BXFWfEZbsLPtfW5AdTF76avtQPl3n5w9KNgh0S/8ukyqA46T8z9cdIjUj
9Ub5ViqsWTxPbwmushz/YWPAbqrKCxpVe5l+THCFpX/uLwifWEaTZ0H6TPaS2mLnXurS5zzSScov
FVsPvNaBt8M80D8fQFKvkfEUXbiFgsJFxe7I8U6Vkq/YAlvv5oH4au1iNsc+I7ZbiznVKzEC3ZqQ
SrnScRvAoqCiOtZb7MFmYxnw/5Hj2Oaoq74E+rxVVLdEXzdbb9cuJ9i+LsX57EppH0fCKttnMZhk
/nShSVuR/AVVHgU1hJgw45feSojifcelGAZXgVr24CWVt6tgJcOXIM+rc8BG7ZdBDMQhfI7p8VWv
5aWk/EEgCclSLFW9ErlPPyKdMqhR2OM2V8fjM+UsTSIBxXmML0uMhb0PeuS8cxYcY/B619oCT2cQ
i7RAGcN2z6oVcRY2TAR+aR1BcY+DpYcyGznRWwq3edBrIWYc1WtX/DCayNBWsRpr2J3k2yV5Zfin
fge6pPsZ7mLvsI78l9XOl0IGMgS/FshIUtY2PT0Amv9m1XVP/Kr4oRR1roudSwx6wESEzX5QDvSS
jPFf3WDE9MmCMlcVGnH6Prw/wVVIJadHPKkrYdGblXB0xqA1cykW9lM02ULFanFHj8usWuwhqqd8
IH0WDDl8jxVIfJYOp28tjUsGhmwCfmzkZooRW3tZQXk+9nhb7ywFIfiLMIAJSWWK4G3TKJ8UEypP
9rHqiPxQNqBZDsMw/egKansplMGn99jQaXUxjPIY1b331Tosh1ZZGXtHykaqb88d11QFuiYWnfC9
PvJqWHIO3VbhZ0QRGNu0CKR7Y+4w7lrPY25gZ0lXD3Jk70zlS5JApFYJlaj0wus+t76ersONdCwe
lgzNhbKMQ5AM/v4tp8bZosBAkpZu/yorkY3cO3ifGSq2goqG5IK59FYtb1k42XqDlLyGjb4IB0ko
iVzBF1wcfbln4VaZF9PSeBCaD9kv8FAlwLMyhZtD8p6xxB9dafTl1mg1mS1fpB1GWdi3gOnXxwS0
PhP40n44+z0NN1XymGJRVmfg6YSNRjFB/sO1ft6e5PRt54W16NEgoM1k5jQmY3JQFj+ZUepW5brh
yFPKnHHTij7DtLzt8a9aWAzz+REUZnyojX23qnEBgcUEpG65GihcsTvgSKwo2TzaTjwZRdzJSYds
c3CQ8jp8aWEUQTdhw4AL4jn57UTgYH6u8fvvUszEKSLgTlfq8Z3FG06hWU+Qur05/3vrt8m8oPLJ
Vku74SxS+u4RXEmhzrPi+LuZnbJ/Sg7xm8ehXh1TEkgaleewe5gx6rUj2i5Ddm3b/r1qPUK3drr4
S0CxzHiA9kUhk+K3YhsRHVhAcrbXlgmLoSjnvq6/79q/JsriFm1/GOzbsGbSvidilluyTnZ3OUkf
qvio2hAYQKGF7UvDQs14h3shI2ym/Q6+rZNlPT7+CrhqpJUo27zZSZe59ycM9Lci7SdQR82lUWRV
w8P8cD8T2O7s3OoC9KJNr894e/aVru8aTD0Rnzzac+3tFj3CraC4XjwdvHjZdRSe8+OAfkBtEjqe
CbiWSTknKXN++EOeTINPROU2EVSlo8lEHrICKwo559xwz4C4pr/yYm5bwS389f3LUpP+ozI7jMgr
mPlS5v1/5558jjPSd5qXqpc24GTCFDnsoDn0VmNr4j7A7BVcEqUIst/3BwmHARZIeAcOt9A6GhCq
tivIagWj3kFU+GcyvcSYQY3of9/YgTUZWqqyqwiS2DWmrg+U8IhuB58+EIFm1eZetnOzw7CjOPwK
Abw3EFUen9QBcDo7MifJDnlPHvauQ5x6oOIcpFTR2tEeGn3VhLgufk4KL/bY9gxCNAcgZxebeJhm
/SGkkJMneuAU+qK47xQ5bBxLFt+PQvhRtGzMc3ltnh6f/7rJOSd9yp13KE9xV1B1oDitS8PhiPeD
opMCGt8pEf1gx30VS65kYlGYAn038kZ2LxJxa5jTLl7jGb6FCG6j7P1WZMhYPfb2Ft5kcYdkYt38
XXUAcug8hyJy4HYxUhrgTpP/o2mjbQ0Nr8GEbGwUYLRJiNzIvkqAL2IIVPt2sJeTCG2y568tItA7
TeVfRrNcKBzaTpmLJXY86VlSnjk1yQ3FRPGNl6v22cJGuL5d3mGjn846LoNwN2IO1YytBKTNJ0Vc
Xb6xYNWIqGJQJuUWz8RxPJ0Hd4p+Oz8l6LxhNUzRP5uvT2wqBQmIQiTtSEU0FUVRpMU0hT0q1UB0
jaJsh62/3PnLSwQ5vi7v7Nuwm4vEEoYJfi0Bi/BUOd6VOvP727mqZrCafzvugF2tm1xk2tBYfEgY
IJ/n+HM3gWgEjrrTig22CtKjPBWcLGAc1yN0lBMLAaowIcxHB7/XdhoO4EAGSOLcA6Gwxd6NbhaR
Swkuw3s47rxZYBNDlCt8g6mHHL8CjF9+zQ6HBkqV5Jwcu1ct5+P+nXqYo76MDOupSM/Xrz/LP13N
i6DMH78106IpTH4E7WxV7p5jpksa2g3Krmx5f82/+U7uKjOKOp6iENENz7WuRIBDVAU6BDp23Vv2
pqvXnhNQ62tRrzvPtlzbLY0FtBC7W2cLhAnhiMiebm/zdLuoYOx0hYff6u2wWZ3vyE0oxHve/mZQ
xViTu687TwmDLoJOMEwky298sIPsmlpfup2mHA9io7PwXdSl85QoLFgB0Z2btEce6/llXYjiOPEU
nd0+/blfW8meY+9E+++UrqBRV9VjYdkcrmKY/8/bXeboTWe9k6oPDmD+TJAO7ZrQSx9+InLZXL0H
XUoEdnEcMjVu6LK2JCpaAFIqWcevXksEImsjcgQ5A6bSdP4VTZDNwrdF17BoTpIgHU0eUjUqdbRn
bIXjsVKSrdvZBKnBUiDFl/iisiDVl0FPyuwqlfBK7Xcyhm39OWUOR+rAjStGO9GLdGgPcj8n+QXA
JVz4q4OFm8QbJgyB56Z7gZoc/blzwXO/9ugtKBwOgxbopYscpDBlKpWTaVSR9L1suD+HWV27PBwP
IdIyjxfHkTgnhBEKLD5C1xGBnisgOoRurpUuMR/FSWgaVA7vu8G65USW4tYrJ6U2v3d91HT0vfMM
1ZnWXcRLd64gHawQHHg5qjCl3DujeSZFHN2IOZgcr5owgZnVHtpw9X9dGpcqQ9+7ya4f9PFsYfLO
SCrK0nrmSd/0TXRsCexbyF4bQa8y9X04WCf1XoTFdjA8Ea24emDa7FJIES0wXlT6ooJioQLWjcxe
7/5oKFMc5WbogMKYYyFvUfiQTmTyNh+3nwCbIQdWbEnQAzr3KfFA3hgGCnyDyJEuoqQsWJ26vYwk
KBq9EeYIIv11sw9/fbIgbAuixm0/OUmFuubYIKagBUJep/wieUnV6PFl8Kspq2gWddD+/1coww2x
2xUhg55NKMWfDNyTvoolPrMHxZ1/pFUQ7LCM32xfKNv7RZMCAxkFohG37c/DRlVHg4lTW1f246Su
v71gPu1z3NzKfDRyhNgW7OP7QGdYs3KDt4kXV7GGunSso05fv5+Is7wPvD9K5K3eJ0I0pM45ppXV
fZUDJEjQt77DXtp/vJlZZYEQuERXS3m6tvScppK1LWgzniP6Sla3vbnBStvYqYApgBp8vrCDglno
1CBGSd+qb9TQWfN9X+LIg0UMXkxv7pZ4uOggm+SgDtAgdGst1jwzt+09nBh6BjdnfwRZJxxMQ2az
MESP1qayef5WfU9C3TRv8EWVuW3FfEkxaXo9qF92edaOuSX/T/loah9Oth+AislaeUSpIV/zLh1i
91q7jOCrUY2RhNk31oUfyygrjAUQ0Aai4o4W3I/6Z7CPpeqjwHax8w3iVFLMvplYVeezdRBoy8mM
A6Y3yX0bedlXhUNKj3ZJy3jfJRdPwP9/bI22DmhlsSFAHzglEIzwWl7glhUYR1guYWBRpsmtz85a
n+fygSQQZTctLbwybEd67GjET8eDKLfhumFbAF7bHyOxra+3hs1WZuw5REJ92yqlFA5+mTA1Eduv
CEqaV49CCInIuWh2LmDOTwiU3GgpDPINIZfwJXBHNcKsFse15Hp6NWm10Bagiznk/Ym9KfrE+bto
AfFoK/sQBVYe+aQV5fRpTUWKbFKoIT31CY9df6jF6sflpgSoF+p1lKIc3+FpnEzJjuxvzJIvmepJ
vAgj6mASve85PELPSjEuC1wAq8Q3eCexYS/WnN62XviwObNnsmGgQxH2p2vTW1D8xe9eg+ibe/Ao
p908QV9oNkDH3TArOf+eE/aXwrKahxGZBFUWAgyMFVzATmwvPpbf2m5/7jLgMdYYikQ3naPtMxUR
f4qRdbtqb5SmHaXQJI2cuP6/r2u26phetGG6AhstsMgmaZxfUT0rh/qmMqv1jXML8QEZMMQpIzZW
c9yCvBz/hUwQymoUULZzuZ6ml6fWDVyhyzWNa4qDRt5GWlcqvEjDQznRvriibeA4QPTI6H0HC00/
QZo1TNdLvm2b2GqIo/CubzrCuevpDJMZyTO/bIKqqb9L1bbwhbbZEF6OimEIF5YGTYRLU7BuDeHk
smpNcfZXf1YaEx6mRkP4g+iWQfjbBO36Y93xPR/VjkJHALCVt+3QyAaVBIi0ntcyymZIWT8zGZYX
EvQ+WKrTNNdMdljXJWCMxaza6XMWjCzFg/3fcO9AoxQ3D7TyBdfPGFjMUSeT+a0V0InGqdWpPWPL
UDKrPN+VX7FaANeYhEnKWpflWRUKDiAWDTAb+dCEyCssbufN2yJ9VoQH6JfamysbbuTP3MtoDjix
p8IXPVq5fUrRRaUVxIs+XapK88sWXgqb9I5QAd0DArla55JDeJ2Q1GGgbTD4du9rnqAoK6oAIKOl
uaDC2F8izqtQWhl6Z8SDO5+Av56bdkmAuFoRsUJ2Efm8uyhzuyBCD7/NTivxIcT2gcsujeNQjRok
DKoD5IKrmceN1/L8XuaTdknlSko/u9LM8D1A09TTZyfuEd1Dlnb1EeDiOCn8nPpPcTymDSZU6mPc
TFVM20XXyNRVWdJpcgtNnvYHrBkqqdfU67KpRRsVVFj1KKPQUn1LD/NKWPBiyskKGtpiHsYcJ68H
knaJSdVeENW711V7TRE55uTX80uMfAjYXqgx2V9jDF+e+TK+tYK6fycsMrxYzQ/pjqCfac4tE7wN
ItSeocJ8ydJslXoGcE16eGrfcnKNEzE5sWItxINlhKGogFbYGNNo/Y9ZB4lVDIBBj/ZCtQ8+ftqi
DqYftL8G6+gvZ+20PF3Z68GdLNG/ymcuRQVs0kT1+tLJmkUHf5k+CeLnldJJg6QcfMAFGkMl4bdO
tIAnu64QndTxqqlk7NiHRthqXuPyckIMOrcV73iEJ7msVBZKUz2fvCCyoUnxCQh9LPjPBexYGUCq
F5e3cSzfrdtHrru1sidfHXClmhYnGvv9IQEBXhjlqSmYFM/TdYpIzQc/BCiM61I4XGlT5RkFAIue
wxPkw8MrnvhrvSOX2GMt7xn16D92Cr6jlDel0vQFm+D62MWgg1PLdNCx2cnkzxYDABgJqG9Awj3a
IjBgKeb0db5EZya4zzBU+/ZUU9f/wBNDdxsjuV1a0PR7LcpXoE36U2QmlIJ1lRZhwWgNcsSku17Q
JOJWLaqXgeuBetd04w5VM8WJ2yP6AR/I9GXbrtMkIpeROAbEFllx29uOfV02SBVPsS+Q/O+bGJTH
Gk/ViMcWbyLGfhRVHB6IkoHGE84tXz2IIZoKj0CxhmwC3H+BKhf/O4EIoFkevI2aN/Ay9xFTVzJc
f+SP4kPmjmIvOYWaSFayMR+5BywbzA6BxF77F/kYGCm6ZjSLAHXlll6oseW0APpuShI+KJvTeKIL
Ien/WqNH/FHnifNiLHdi2CmHrW0l7iqN6vZtFnBJYBycrPIMxnZ96uPoS5c4Kf63r4kc0P456QJK
wr63aVaK5mtgwYvXg3VqrmRjR8BzFKEWV9faatYeSpyp6c79cpUZYErF6Qu9FSAbNDQvBJ/BBDYx
jydtxRGMXumaR0C/HR5pEVj/+gKZsOZQYQbFu7e6z5Atou+wJh904bJPKl6MDPnc4CIfcxDIwuwP
u6ELn9TtITrQD4LNENqOfkUgGMNqXJP6sMiNiPrQthU3mimwV27iB38iJ1p3s795suGgw9P8CJH3
XT2altnlMQIL9nDb/hrJ/0S2zpBwkpTJLRCvCNTyTlRMsu4OcBLDZYMeqD9k2AXXzRkhC5PCT1dt
F5e4zoplaHbkEMVXMPInchVLzj2lGTD5XsggGKKj8gvwFYMh9ieoPGabZ8Vh7GSThahdls8mwWm/
dIhKMW/3akcZi5w3ww5eNCqZ5v6a+2Qe91akUxvsghQxbacVTqMjI4G7YEMksaDRwoZVHfqELrE/
8VLBNNghqyjjRnfpiDI+AIPhz1Yuh9tjz2zTdJ1Iuot86SQ1Qlg/RR7f3ThQJWkPe/18rQ0G0CpI
GlJOu71PIB56zhMgxAzhbnnGWaggiykGQiJmdTLlp15T3H8SNd4ABG/easSuVDTIpRFhu+fgV3kh
qZkK5u1P/+T4MRDZXBxkfsCnC6BIva6h9UqeZUkMW9oPvvxOCKX8GHrthfJ/A1LHa7iAp9jce6AF
KaINfq+sDpJzs/EzqRJZobJQqxD1frIo+HqzoA45Wfn3GOI2n7Vpeg1NEPOrdnQoZB7vchZkuD+f
6URPMU8k/lGKdewnh5WaKMqql7Hp9vXQfMgVnwE+CK0ugYahe9EZ3qzyBXVmncUxwKi8QvgRyNV0
DCv4KEO/91hfJFdtFSG5jK6fJCfzgBHuxVypdkuTLAOY/NJ8gtqP9vCP+vK9nQn5en2NCsARyJcK
7ohqrmmSYLc4AsnwYcMoeww8w3VTc9QnAmA2Md3ooVYIGQk1IdNE0sKNvg2qV9zrSQQQLHBQXuSa
Bs6vPIJDt4WFJXTB1vd3bjHC1sbpF8sY/4TeGRfmIeDZ6dGMTMlrySKqUC6JOl+IyijkbfVC1jP4
co9C4upuR6fO/SZsc/xJAZST9np9luu+YoT26mb2hAVMZUgIoYhs+poE3cT1ODjh6EJpXUA9oPd3
u6oJPcz0XUmAoCfL0RuECG5w7F91BkP+yDkcvxDsEwT54FY3S0VlXaOyKsvnbsk+Du6RliiQ45V6
730fF0uvA7UT9jsb1jmcBvm149sZBRnSf7UYaYHgqYIZ8aP66cBHoU7y6fjDxLbNva60aJwXwal2
+PiBeDYBepDQ/niNLkoAs8CFy+13gr9m7iQP39VbF0NxQ4oKC7z7usbbMwjsyc8FPr23WyD0OuEC
4wbNnmNpiZloJ7qU1fIpIjC9SlZaA/7OTGfd8sQv0XAaPe+7FxVJIvbFP9NeZFd0nFuC4IVmMvv8
mFw7gVNOvvLRDYnyHtL241iM05fY8JpQ9Dnu9YXG9e24ZKdz3MKcL8Cakkd53altgUBep1QU55sj
8QCpkBM/wa6amtaGEfEw0wAX3sY/HPWx6NkufswgCJRnWrkh6Y1EzlUyv4IBlIYRRfK3+vVQJJb9
T3BzBLD39ct+WLwcophdubKawVxBi/YMm6mzlrbBFtcJMjIj+f5SRDncSUI07rlAJHepqiSIpPXn
SpiAf2Y9C7Af+uN3aaP1DT5YAk6sbkmJaxwOYbIkwxy6V5HyFHnAXnHaMBULc0O2lrkVMZkEt2zo
HUBE6KKs2PWWvNXp+LSn5yevgeF9J3gx7wpgrRl/hq09WpA62Y/cANZqH8lB63BzuxQDjCZWNbOy
ntKo3316zApJONCMOVZxf52fym6w8LZKqJvdZqWVu8Qw52bWkzBsF/ik6XqfofFOUdPQnAtWf/DI
iPGIlkMFjmeUFiEV/akPs3g/E6z8ofhbadvt29Rdj/gO9aXQXN9+LcMKMH7M7qR2BTi7hA3FLvSz
v0U/m6wUqwCoQFtb2gXQZJin0VaVkWKJh8KHjZ1bnCD4UJ4OLY4uBBfjP0j+l51zEe9soFFxUNP9
iESSlvaMLBFVjM9XI11hjCZEB+kdyd3Dc3q61FJvyNsE9fmkeRm8rMvJi899S4P8/ZTHEMWbJ2GF
ztORc86u7ONqRCeCQd+z0IVmBDZg6r6q8Dpok4fXNiArMhIT5yl6afFX5fLcjSTd8jL1oiIr4ae7
G4kkPAPiqQm0fTZRkbX94vQFhvYjyQuIltESUm9DU7QWfKsFy7Sbq870YcmVa0/xleM/LILme6D8
SQXDTu7bk9Jv2ILYZKUvxF+PplgJ0MU1fpD1dat3GhAf25x0qC3gwvcEbWcTUejTp1MwAMGztmh9
YzV1EW9yxHtpPOghQqu8+EDvitV/EK+Yr6R4ZF6Q1W7ZhCrjpOd6/c+FCmb/dSF2cAskoDO0b1Rq
SxaDVYnW70TNuiqsbMhJeMruD/t646YJXdJir5KtiQwEP1qSBIDO2NJcpCj0BObFtIrtjeiL3jat
zmYVjBriONn/qT0jgWwUPdmFd/NSG+9GxIKYk+VcoctEppqeyijL07Mpgt8SBRDp6y0jRjdQ+cBR
GwbRR9FtgyQpvxikDxU57F+jNKxq8ZWsXRqcI22WlnOX9U43FjwSl53Mb3lTTnSTr8a9Xav7jO58
Px3kouCeTrl4BCu+Ic87adg/phL4qYSjffjPxdnXQD4SqWhFP46RqWjUQ05S8sXaaUXdwJ9j+Ocm
4QTIOSa7KGxNImsoX+pR9MJ6P3FKKjvBiYP2l91UHelUC8LED7w9cLMSbdnIKlk+smWroRrZg6jD
RHdClKoWD+519d+kPWJl/DvLx2GqVbxH/jFfqx9SwNjLtLK8ngUcubJOb4BULuo/SdLtYDH6FM2o
FQXeEk+TVsVSxijT9K/BXQashr+Nfw00vbaa9slkeW5gn5lBJvM5T0ag02JoFA+sPzJ97JsJLDZZ
XyLIzGyQN11YwJIxAv5OMcq5BwlKhI50/UE8SFU7N4p6i6va6WWtNikcXDepPsbFEvMB3tH0OKjJ
U2TiKjY4Xy0Wla1G4YFpQ1YfNiLD4NiFhUqFx6JENxHI9jdydvbUHnxlYDJxWNazvJnNvezcna7L
/9BGh+07/v4tMDzjPUMAqotbv6u/nQWYE8sPvTnSoVP1sPqx29wgJUYH27XQKZWRwOzUR4wzo5E3
U3OgRA1DXF1sPILUhI+Ja0pd09vlxOTa+XlV3d3m09xKQCoWUeH4QCDhSI9qbdWKSDUolzXFac/Y
TinCSo0WvmtV5sUzNna7dRhd/HzL+DRNanjN+dzOslBNIA4Mh2mcrSdra+Fld75TAXr3zStEEjQx
/WLD8s3ZA2Hjh2mQxXW33gjPkdnRI8wlKeuYmKsciOKVXQXRkLtGYtN0eSQxzglCoompoQ1IOz/V
QUgb9lz8kAz33E+yv4fW8TAEVpdoo/7BehKt9BR2RX42rmHWBLkli/0hE9FLrXlUIyq0OLtoPRYM
SQSDcTMrWtSqhBAPrLwer/KPzoIcLI1XzkdlZHgQdMwf1L0sSDqmCRLtrZ+raF8rtZIfQNg9SgBK
oH/hLQFELWfmolYMGeKEVV7HKCA+qe9wsRrrnVJ10uJRxEPu5EhwH3YsDXfjJVk/8c0kfqfAJJh2
vM3Yzsxuvsg90dY4+YffroSIRLiAPOlr3spjIFM61dTKUq2EzXCDfwjXfkfgA0wqAqbwDTmn/Iaz
dY2+7wdpTSSptag52jMH/aA3pJr8vlhSDBeQzmkKFHgAObWwrGUa7FE4QHbUgMrsWy4rdxMvliBv
ywMU8Y6P8hwRcrXpMmKXJ+esDJbiVU74emKmkjA0YKGY/K9mN1BvahPB0MCo87Q3CIg/fS829dLf
aObRtKZnXuf44JMAPxUsB8l7e3PFJTAJOSzBMRapeh7S4sYB3Ixz7MHA3ImIPnZ6++PCXNYmTesG
G6IUs7BQWQ/W1djMPc8DBSw/w51D8rGvqD18HunQbx9Dc5IIIg5QuF9gILHQ3wrBMvY2KBN39vW+
2sTagRnHg53fdBcKHVjHPXfbWYogUcGbWUWI23Hci6L3PvwYqflWrFruMIggCHhS3PRyDBxB/y1F
fYN1USLSCfSdhSwCNUW11uEAtQzYF8miOBmw4/nlNTkxfaFGEZpRJlddkdEnYfe8FS0kLve2FUGy
21qMvzof2VUv7WtyMOwg6E9qdUtjUvA18G8UMQ0VQr7NC+GkfVFRjoUfc2QIGL3S8qAjIsM21XXB
fg0SpYmuTze98lAiq5ZIE3P7RbHMpO6PGm7SjN7HD1FTQOP+IWxCFMi8y8seRg6oi9IlRv97AtDi
U/2xB+sv6iILNajLCrqW6IuB1sYqhnLrs4EM3AtACLWlx8JzUQGdFKljQbgRWX1Lt0ceU0DIeuf0
a2WpvbRc3gWsWTq1bGy27PgGNOpTCKNA+qYpua6bzEO0prk33cxOkyBTaN86/4i8TLePt/n4N5In
+sodqeEx30c7s6jNM0BNV57LjA69/VEx4oWjltTBYjImq0FXltdgU7Pv/lZMTZ2PnEzp/upbA7WB
llKvCEbRRMWx5M3bhzpPQsVM/IUyabyuLiw3UkLadclZA9MbRIg7Ee2GT59J7EdN0qt0Qx/GfYsO
IMIyWQpaILo5DV7rtDZSIhA7clK4jOrsbkV+suHTvQvHJJwCQ7c8yKumYFuD0Y3s2PzS6zZhAQ2B
siQmbSiZdaf/cj3NWVa83EB1fiyxpf7KKEAnLntG+n/YyH22yAUWLBpOZXEYW0c8SCvQZVmY4Fnq
1Rjg5lAtsqS7/e4gpox+YQFJjQk3pMPVdT+gpPNZFAkkDynV55j9qBrF7iH/LsZDpmArI6dfo1CT
IoaO4vMTJL+nbK/KfyG/4r1BieC+WPK2ABAEICFqIwsqC2qCzURIJquFCUnO2CkSH9PsazRmvWrN
Uy94HsWO26aMOkErqPKjBh7pbVkN5z7NDV1+NCDUJ7yNAgVX5ReFB9PZB4qVERLpWf8gT1H+MRYA
eIY7eP2OK0tCQN2J8TlnD0W4KRX/sZUxsv0wwLL9Kfuf8L0JOmikVlevi9xbX84/p0LngTo7VeG7
0BxIOU+033NTSJ1v9zX6pOTfFLe/pTdJvhHqpAb0i2d9gzHgJd750b07KwGHYyYWZ8ns7aKtShil
0JkxFDPDUi+MYQMRN6ahp1BLAyU+iAcPMFRNWbf72YRmAV6hIQuJ+YPERAi66ej4ehr1wQqsVyCJ
PN1olDW9YOsqUVi1SoOLVMTU2ryAkkPECrszzoV5WrDIzBcL2x/9o6/MJES48YZ5NO5xZvEC33Qq
05/3sJe/hbrxco6yiFmgvcPyAC2CpQ+fr5K58KXsja6Ew5fp2vmTdvXyxBvdyjKHbWzJX1lhUYv5
WVtb8Q4s2JRx6wYY2jPUsdArspOKdiuhhTP/R1XQ0oiQGVWVMCqoUn5Myty3vqQeo2CJBF+Iy8gA
yewUZ80dfpyEthoJs5KmWES+8VjXlfz8kVPx+OjZTS2g6US23An/lXpk9Skpt7V+JEZY4XJGfXVs
c7wRkkUMNozHicKhg2D3TfPH2yROtxamWVSHzZHyKk0fzqe6qAxZGLIfIrTwA3KZgG8JUEHP3GWe
sRLIbWzUevjFXGcy36KFRDyqI3IKb3CARdgj3t6AcxitOoOnMqJ/iHQfcosj66DJzxN0DdqwOnTR
KvXs4AYxHC6+oj1OBLmxQzLRy1aMRg2W+lVViz/Me3GbPv+Hx0uqDN+DYLYw5TNHJvwmZiKJN9hZ
SWp0Xk0oofE1IQ7r/37l/4zk3Eo+FZGD7IqBixGXSWzKyBFUXM8DQJdUP3vnxRcgQYB36HdPe+qN
ZTFuSwRm4NpNR/FGBR0SCoZUKJ8Ha3FBa9sh1XuyV6mT7rKxufeBaui0ta0FdUL60c5Si1ibruE5
3Ji+ALHN0PMzSDUuiZz2lsiGj23mJPcba31gYaZmHqhip/9WBqSbgI5pwCTo5vqtSVyXML2JNbma
VyxmTucmj+Fea2BGUPq3vzVAnzGxb6U/gMuYXeV0FxJiDTwDA537WJzGv0q7741H8X/RxVUsuz8t
ihxbY8fNNkBK3dd/xLMBJe2jPYXPcuBsZpCNH7xv3niGUM/Mi4gKYf1FkuElxWizmzRl9atY7uAV
Woc+gILRrYPi22ydPw0IWkdPmhsO+KUqEgpkH1TE53hOLUXlkpHAxQmmnQWudbKmDS7OPoAtBLtc
L44xcb8OHx1/3T1QI7zlayVixAVitYCs8vZQpj8RQJDI6EUEE+qKEWjnRZVraPsgpf7iUnTB6qaA
7oagIpxm7tytUfDt9aETW4B9fyHNbf9XgmCgFdyN5V7CzCtsndZaXBMog9kwC47h0mSEROYegQS6
1DZNj4DPc+PCT5m5jmYIJ5xTnv0Fl2pUmxoy9HBsptVLrmkK/I7zfC50if/WDW4f22dZW+9h5oyP
lY1CW6/Py0yn2yFUMykurM4Sw/xmbBeKeShZeDJwyhBJ+sXTBJv2qlCNNp3fzg45K1HLD0QcIfML
njRod8OZZ59JcGu/bXxbiPFR6AsDCOuHIjrqmKV44+ICNgn6fUOcNVH/X4Tz8fie6/HQFrmBB/SN
AKoWfR3hV52E7axt/fOk9NJA0JID07Yc6cdxeMc/UVskm2Rh2jNtWRLJTMCo6QWr+J/IDK89n7Hf
vmPU1GM8eey8cUvoeSilIKkY27U+vxdWUEuBYTE695cfqSorCKkFNDa8d+SotlolR9y6lOn2ebG9
e6A8P8YZ2qbx1/ZCuJxfsX15SBy6Wu905IbUdczAicd32Gd+rU0Sac/DVAonbA4ASYTh8zbgbtoq
+NRYKWvybwE2Myh07MZ8at/ndYcx0pSFXYcBwi6W0yoU8Ffk8nRHPxgGJqs7cWSC/u9uw3nLWu77
CUNx01UBT+hb/RCDLfcNxu8T/lJPfz/d1/vBUr3qOI+5ATXFXLKSBNW+5o8FojiOTzB1AzFzi5ss
NByx9n8VKL72KBrZ/IkiFBsXFwFZe2///GtAfeyTHhrlZqwuwi6gMdTT4R+5zF2xfDUAePlfQzhO
jeYLY028DuwEqhRxlQsw37spVzmuUBH4O3Wep6AE7rVGxENJ+q61wld5U3ybj/HPtkolL2zqzZmD
na1Dtggv8HQSMDTQ+G4m9ZRKz9x2jkSDkgAGcgH0Ot1Mi8Nb0RSgJXL83OKcWj4e5WZ765OgnNjw
6tWEAK5f1v1GjU4fYnhAEBzx1oFfyNMVTIwDHnmlUZ7VX8+99s3lnVmUMiIi8wshraPPcLJkzrv/
Hf/DwAaWrEFSkiAlKkG88FsMywiVfyBdhS+1KFKCaskOHb99WbH4hNc097lUaVxrkUdBvBsDizYD
1+o4bh+2DMrk0Jw+8EgNctLYeU8+KMYTmDTJeWX9wKyILtq4aR+1MEPiuz7VxzP3JVQpYMLtmYRu
LWGZvvolQ4TfVhXYoUnL1HYKQep0hG7TLdhmB7Y1VEZpZvqoVSU6tcoo97Z5g5d0fs1vVm7MkwWw
2iRPAWTEmio34LJH55lg/erOhoXGLIeHNLFQIfQYU/LHIVe/Qy2lDwUQp1c9xaJq8XTJhLcDC3OP
4y2hx+SUf20jBS3XYVw/ANhuwcImgNfEfCEssviSt1c4QTF+hXulcrCOM7axyuDFgBs+LqbnM8JG
Tna7w9s2HFuRKMQXbpmtA9/6GdHNxDNuSk70rRDoabrSc8QbIPhWE32Ay81rQSSsXlPeOjeRhXfM
ZjBKVMhnG7Y2cIf+KtBjAq4vZ4xMEAu+l/0emYC32cCux2NfljNhD3kYWeVztdctwZfNDc2JnpO1
n66/eZgyxBWbVtxxkjDSZqPvUSAMn2o3kZs1nQptIxQYJNVwaONfL897rh4Q/h5/RR2B1grWFQi+
Qt0BUACrv7Vu1wR9f2d+ZyF8YtrouBUM8JNaOc4frWuf9Lyh5R6K3T4Kp2wyZX+jvlA46hpW+8p4
iDlklkSbj7O3LTlqB+H3Y/nkSO0Vnp0iLHPAHj+/4Q5ud7K79bckNQiCz084AvIIqq/AgMbJUrY9
EFmzdn9g3Z3xf2koDplQ7HTiqTxlFfvc4MmnypPGYH+MG1Euhr2tgwphQwK2koQrCOB691Y9/ld8
pqlYUepbOrW6wl02E8JYPsrNA1ixyDRD396+bTn0RGu7f+ai0n/HO/kbEVio8L2Zvbc9drTSBdPv
iej3DcS6ok1pXdqAcCsHkllI+yuuWWywUOlIzdVrawQfLFGK24tNbaoRsS4QuxLsxklkLswpVdXx
qapyLVSVXbC+N376211GumvB6lngPR/nuk4eW0iAc0OUqEYm0J5DlApADf56soYsiKnuBJtgz7n9
o7J4wKlEV9MIF7x9ZLfNGwuQ4aq8H3sAJ4LFSxp7A1eLcj8EEwqXvkgNWdKhMSeRh84HLMxvGzmP
aUuOQh5ZnG/OR50t+GbDBL2tzInbJVh94oCgtR0fkW53ZAsI1H+hOIdHCrR3yb2hu0/GIsAvlEe0
ZcL6gPSL3La94tdr2AbhAIxdSkQhBDp4ddwa/TepbQM+HQ/XUfv5h8CwokG8G8QldygUOS8ta6HR
/l03AxWp3+49nHWHfnXeN8gxTIUhutrERzYsR9F4SRvu3dRIzb23oJ9RRVzvFtVzaR34deutJLl5
F2Af4njYjNPiaU/jACYfUGqmKhrrOt9lZjLya76gRjvpzuosqspklvFKlAZCVcRB2iCLuGt6JB8+
gxD4GX5XYhEa2SaPNVJrOJfckA56Yl/LzH/DjAkagxtbO8Fk1FxbBZjoaJRFZGWLhpn1aIOzsdcJ
j8B1H5u0knEiXXJ6i1fhU0d3ir+zD192ACKxx8cbGNx+VbLsTGhLPHg34pglSAcJFWMotY2ul+QL
alRxZ3Xx2e/ZlF0r3G2snfZEq8xV4s9es4nEoOplr8+QDxMMGILppxHQ1H+HmC2mm/GdSxLJgtA/
OIiJBAwH3xbP4oExc13o8/I6mbcCIaZ+9hvfz0dTdU9jA/QDDaOr2LtszqlnBGOaSbwoocNI/5e5
HsOPFcTJ9I7FQqzyB1S2Fyimv61bJZTmC3h1LgYLctcQrkOKRWlmZIcrVzbPThd4HrRADI0OSuDj
CmJ0d6suZC/6cm2Ww9wN//cZ78OLN7HU7cZAnYy1+GeFr3bocjVaamd5Wt6A0GTHtNNfYITwWbRF
yMQowcEYfj1MgR1iEUlZxY4UqnNMwn32BHdBzNlirz5YghRnzcISJ2rCFQ77q0Mdslpem0q/OcZ9
XPmV+rpZ8cjrLo4dRS1ukuUdhxTOj/kVsZWzgB5fSYwnHzlTarn4uvdE/agLAcSMYlkutbfrmQtk
TTveSAAlYEJMOM/V8Qf31SBS4Z/q5230nRwx1x8/ncgxmqXo8ab7PVq9z4s87d9hVDwxuj4VuujA
Orer4xsYtis5Su7+buxajj2MtqVA5HBdaN3H8dF+hDzgxDEv6SIy1iQe8GepFxPWGUbyVsvKevcf
mXcD+l9EhPzJybDhggehx/02PbPkcdyywTGtcb5j0Z8o+y9nKCaCic7Ia88nF6qDTJ5mQoFitRPF
/eZ/3S8hwOFgCpQYoVb2pQ7Dl/iQ+mek4wH8qxDo6dbnfGruAyrJf/GEe3e52u75kg8QakRnPUn4
/8hGJScznFnc/+OpHZKL25WsaPJWwJLF6gzVZX9FZAMkr/ipv42ZcKQ4TBt55F6ZiYZEcOvtA2Q6
GZzzjIGM/XKHeJm4PX03THbhjZs3br05XnANzA2opqfuOC69DMmxZYX/fcdkkFkkdSyFylRdiVfr
M5VMRrqYsTD21+jFqp+8bAMM/lrsOj1DA21c0Q6OZ/ixdzSPGzAYHmZ3tHKgzttm4dkf/Irhjbqj
/IbmlyMPDQV+Np8D26+qpPGLNQx2yM4jbQ9awLQlD/veNJjJ+AatUL50wgiy4kJi36LMuqGseUus
/iYfwfZ5uEs7nouUKHXJbi6rS9sItmIe/DNbOYgZ3rMr9zmGNhs9s8Tzrb/Gx22bFsMErcVtHWGq
aegekA1sooZKSf3XXT4lsBiQpWyBQt2pSf2UXo43OpDZLN2f79yN2O3LHOykw7gqgZd+K3Ms6zUb
IIa3HVN/gVazZslqGaa/iTRGhnfNy1UiknvQGCUpYNr/Nw/54Jk2z28RSo2gtXW+uqyKeq3I1aif
HuuQgIf9eEG3beDaTMlYshOzwx3S4xGEYkttE3xG3t2SC1IvwHnqaPcvxHn0TIXjuYo/5hFUhgjm
dFxMqRMlBuzKsQ5Rqj8f5fQlOCGCuzAJwM9pGmOmvsyWVT2ZkJdrjTxgNzohebz2gC1b8YnJxFZi
VOdV/QIfsswPrP2ZDSqML1inKp/MrMgag9oG3OAub0jPGDLUO+X9cC/RqriDUOoB/Na+38BL4rhf
wLzCm0dxI4dP5+qAL23eDsazUlUY6CDiTlMQ+QCqQwDHBYT0LQroTxatqtMHEv5yvc4zYSZkbxVY
1KEcSxVq9Ou5tvlj8q+i2ayKZgnmN4hN/tbmFn3lC2QpSjd2HpHqaax5TtX6FlXPELycx3PQUjXT
r2one+MP/jRrPaZsVaLUu4ECuDLeDFQgidCLn4Gn+VNqZsC/+1GYs2NOjZT+eqg1ucZUe9pLYZx1
sMsFZTYo6Pr4XvuVJMFRzG2oY7MoOTjddbdhiJDBhMhhnWOyCfWnXFyws1RsIlCpxjrum/+VlROW
yhAlmQzXEzhQK2vrRtyJACEJO82OxBVHCnmG+a/Gm8s6v+8bUiV+VOcX11IqSCkUp46ypog1uJQV
6tQu13rLX/YACOCJTMHIklLUuj3rIjnHd5L2RDYsO/cMV/vSpuYgcXcPgdsqukhsEWjvOCocJsha
8PVUG3sh1vD4sKtuBlaHEGuH9fvY/qRb+Q1guMe4k71ca35njdihhiI1f1svsLhWm5CbhQHdnO1r
WDXZ0qkjcUkA0BL6vNV5N2kVNixLJcLqJBFYaQw08Hso1WhfVGDQHlQ47lvepZRgiBC6jPdNlU0/
N57nUD9RrxJveYwJ3Kt4BAs6sr3FjwIyeoAfR0PRtMwAICHZ2F+n5LsfhRbgBTJdKll2Hch7v4LI
gQGzt61MDvbcrUjGcMSXRtu05Yc1DDH75mKqhoHvbjwTbnXGGB/BdiOGrIFvJokD16zACcJpS0PW
MG+YaQYsbyRfwSHClkXD7lfgU1Q+c9oR7sGOMsZHr7Wdu/91ndH33omuzuQcg9JYf1EoyQ/xmrr3
YwLChMLXL0iacrYstLoswtpq2loP+DHu2D5I1RQdTdlTd0M3Wd1+bCY/sULdWBn7tUHYODHi6krR
i5jVzjlaONPZDn/BUiQjmoVPayIzXspGhJXcMuAIdBdUTMn0f0hwa02oKhE1pRIV+3a9mDZnfg9I
gKPcvBo8JrS/+iIeVS9HMg6+XotZUHwLMuo6Y1AWqBcS6yvNq2UUKURgI2FdON7849eH9aIT6JnT
iLv1fqoXGhMgcALOPlpJRMlfDL4730XKbvFI5UHFxyOzJUV0C4jTz4BigCZAommIYEHunaGXHTUe
NpZ7s7cEgOcwIREFYPBZk2faByx+sgXP8cPQxU0YwvT+qeOv+/gRjoSfbvKBzO5JVcjttCxy1d2L
sPB/fbfjnby40WX8QAReoCNw37BfA6stj2mIKFLx67YdVfpgiXMXQyQymD66RolaEsTnI/JEES1H
30hGPvYZcmY68U3TbFQjjEiulB7OesK4OH8knwWUr75FUhq9oR/mPJBweVpV7SSJNd4bxwQmw4GX
2q3NRcTN4N1OhU5PzQWJ0lTup2Dr3IEXdPAbX1O+4tsChwVM3qreRv5/WOy7M3RJAqac0XsQSahA
KkAvTRjLx4z6/7tb04LfRJvPF+jerAFvR+PjNKbQdSkteThT5D1jFPwWZHKJSCiJtuWFcMvrpEUC
jBPf1tcewiKGR46nxVErNlp7p7RLVO5w+ZAF76ek2k8aizUMX1QaePNBpLwIVnOjpjxuWEQj6xzz
IEwnSKkvOV0LHNEug29cSarCmjiz3xGNHoCD4sclMbCRbFKQUzlrxX7ybRGfZZsn2rEVvIY/Vm3Z
PaB5vnl0EchH190SQYkJF/Sr6Z88HwC2qPxD6z9RWxMLRMKersRO8T9b77/VMUx/CYOuK345sUJi
xfUmLqorAU2ieiIJgxYVeBVskLKLdt14CsUUwNIOlOb14fIcPE5cSCZwBGyRfqxn7q6mcmzRXzsB
dtbNNIhYEkWeLmLvzRto4XhOJWTOIHg3XG6ni8uDSmnaR3GSd7aLtZg84nab3dnmjlocywl0Zsjt
p3GtDvbhw+i0Q3iOMhjoUWHD/QqJ93pM1IpMTjX8KXbrqqLWUHMjjsVqKj8oKA7XMw43YnDcahYu
NiTMqXMX6dWxVCcx3qwTGw/iUfrKo7UDYu2fHOyraeUxUJ8tkq3jDpoKWSh+HPOPSKCBJ61Ir0Qe
/Ydem3P9HUlY4dIOMUQaDWNdNFFIatG9Ta8zbtodGjuQQPE4+A0+AUjW/x43LGuNv7DYMkbFAGXX
+XvtIv7HZArkYgjhmOHuJzpGU++NGVYYMpYqRjtQIDPcFph/0hIOLUm7GxxrryqmWs6E47sTHqio
AamhGsbmbbJ7tMa8BmYm8jJJryGvsAmtY8kx4WyR82vJsw8J/a1Ue6i2U5ZMJWNlvkRXySkHIvrL
A1x304w84kOvsZHlu1NokwT7e+k8bovO07AYFrm8taWxV1+uNcxdbtbod7XDKa345CmE1WJsTJgI
HhZlGaHMPkJ43qJyFkubd4Ujp+4Nk3UK7DQlOH4t+MpJbGQak+L4eIIRnZjOvOKWQ63PamHYG+Ej
/+klN5KZgC/DgZTWj02WdQUlysFkbB+oK4mF+Ev4dVlJTaKBS/jRMfORBvPivYWHPay5SYTA5fq4
wBVIEpKxjt7IcehjUHiRMtu0uZvvfIRxWME1Ns2DDgL5eIVm56kK4Gh2bvmnRMyAZv2VYE1jaXyw
J+tY2obMVWSvLVygFK8hKlRkeRFZOLzxKGMVy9XMcOuPWPhgu6MscNDyxNgZKgQN5lTTzc49n32U
tweWCCNYlYSfwsYzFjbKKRzxVTQcE4SsT3LIvq6GZoPvVslMa0HhBuNWD70qCfGLZy1z+lSwEE1R
hPJuXWtispyjzLy5DsRj6EB+8DutDgKhpQ8wdf6SQasOTrQtwkj0aSyq5fTB7UWDOaiMnrimisJS
wuwV6vKslAp8B882NHDevyHXsDS/ETVQiEb2F8y2DzHuH5BzWbOE9MT2ZgReZBrO/HahfxVN16Tr
3cRPkbQs8s9EEKcpIozXxppeoGYRocIrHh+1zzan2BUmQOuBEJisyUtjFH9dXkuKzG+svUtNdgyd
p7H71UIKk478jTYe7cNOn2Gf/dJSbgktx+uDTXXYOflx7YKxHTErVI3TIi567H3TiFu8zVpOAAEo
3BtSMfQiZ8ijZq3vd+ui9Os7GckYb9tS4ZWzg2LWknGkgAKOqywMADse/uqZ2yp5IpUAAIETJ57L
Jefk0NkWrQmO8+Lkx21kYRWRk/vy0xR+1ddX9nJPvLqD8E45TyUMlc6eAdi7z3TbCLxgJWZxaEHE
ayVyG1ZyJK/1F52WfXniFQ8YFJeD9EEZwgSZpeV2MODqa+vSaR0vgWer5+2vKq1FvQ5/YnEmzhW8
9OMvd2wyqRU1XQF2J8eV9bcFr8WfuC/o16iww+4JaWoRray2NtmHhRY5bN1RW1OO9WlVtSoy1jHa
nZXNI9h4lr/Ovr5Mldmylz70PwZYXAI58AqtLKo+NJ9TG1KD1Iuot0QCQhzGCJF6k4RlsqrR2oCe
BODnBg5FpWsB5GnbqZ/B7F066hrm3oHI1p4ZN3ywZ+zEOYOQj20NhtyV7BkxE1ZUkBn9+sMVkVzl
FIOByGx2k+4xX99tRL+A9JVPjXOEdyHk5EbL49I4qD4SrTEzZONTNwRQWOeBwELf5bsYQlkvMVPy
dXOuopLhetGy43F90m5arBQvoHDd5v9kUe9CrNjOtbl3OxvQGjCg+ybjdExepLlTtVKHBypCXAMM
P8FqtWvfXWYhe5Kjo6WLgZG0JvacYPfciQhmyQbn8caWNlxWdkDfTtrnUGJDxF9lKuP7rooa/bXo
2INL5oDXs6KQYX1oNGsZm81WEKxd6nnxxs9Z3/FvLNt4/Z8s3xY2rBEsPKd+HszDpp5kYoAwvmkN
8eXW8zJ16ZHSu7Dts7zcqxpLY6+GOtqi9HE1zffpxZ9Kz3nZPubjl2lug57sipHjnx/1hodxcEBV
1/X6Kk80yqYvE2BZdBo21dtrAN/0af378BeoJr1k+Gych3C6OxoG7Kkgokq1B29OZEHdNfC6mOuQ
RZ6EbudsQZVVQjT8oUv67KLtXzlS5yFIKIljW1NmSr7+VN3X06wbnUNPIaXlgi5gRTT3IOmby6Hf
pzSlpQ+n6z92rC9r5hUlu5eHoe9HU+DdiVLYd6YAOG2CXPuihq72S3IIspF3htZ/nlCdAC2lYZYw
xoPOe0rGLPm2hasfcRWHVWubP59y1THrrmeDcrkOXoK+zizhHO01o76DAGpZLcXcWHGAbCY1IRaq
PJo4GS6go50cEogJIt+yRqfvi1v/WRW0fbJkSPNz3kbZYbYi1f/QdFh1xyTWSBYeQoJkoQiDUwZx
MIewimJDTgUdlWoANiXuCZQnSzjDEJvCRufsLiqFqHhQUy70NlIoKZDLrRSDYI0pIN8HIM24aDka
G7nZLfUg0TOlG4lEw8/Mb2V0DGtwCicd6PFWyeW7J+BZtfwvCCUdOMdODqW7yqS8/i5oy7E0o0eH
dCFkpdIDWOu5O8BqLnrvVyn3Ycs5rP6WbtLBIjTrEafbnY5iBLUQWHWLlFlG/kFKWLpSIfahEQUx
XXe0A4n/C4qaL+3dLhznbDERxCukWQ3V7f6VvaF97Kr1e2BkW3PUnOXZ8q+jWjvT8hi8hWcWqbty
fA+nHtJvhOeRxOQJndD6zQwe8kJ5W1s0hGLfwH9VsVQak2U1DUfPqgenCtqaRKTS08BNGa193cGY
IH+o3YIknxcGy1wUVUKdrvqza3l0VO2Et3MGKHj0tOq936gAXNCinu6a5guzZkYFmHjSE5uLxH4F
8COcpOmYWq75571701PPfN5pc38bwP3b8pZDreZSyNycF8NyqdnWuDxMMEbwuE4Oc6D1VTZBknF8
M2TMh+9oXKB+CA5xHZrGRHz2+alBzYaEz/49ACqRdfXCT6OePyMKWD8tSgv42y77QY92t63C7jBI
9Mt9spkRZMHVmb8wwh41duuajWKCbM9e6rX9DPM1LE736Cfag38adkQW569z83yyA4AI0GIOsmRn
J8uPBrTQI7lhh2cmD362T1UGOTf+XNyMMtKRx45U9K3WZKpiqVi+37x6y4vL9pEMFqjX5LnI1P2i
4KexvkjZS2YXDkA4ywaUgIIUONgXQemwe5L3X6YIYbJtZXXEyskeTzWsy0Z44fIjA9bq3HsCuyO4
QU2O7RFTpV97R249Hw+jwiPISe18AkPGAdL00QSi8o0g8DgQiRX/ZAaalmd0LkgdB4BR7soG/AKF
EdeKoE+XQGOF/9hhFG2/uV5fQhWjdBX8BEj5wsz1pjoXRM0N4q+J4F5PE0/9CzpslJ2Bj2X4BU7c
KDYNDY41X/FlAFrw0oFxTufsXElPlvvXA39WXQ+4f09y0XEbq8oAGJDmKVCw3Q20hD/m0h5bI/aO
VIr/U3Mctx0TEMlqWBh3ZYkTr+TATA96CnWDivlm9wv52z8DPXK39eUtRfiC2FifVDSIPjU+77cF
BlvmZXqbKDNutWkCYC1t4GTm6sRVC8anYr2bmWkwETmNAPJdVp5N3C6ou24iwOjdWg+jar78pVqE
s8tADI7k5LuOMzz8chqZGoMNugLjVchNF7bgoXvEzjP/U6AZFyvr5bLZ8AngfsOoWSq3VFMIvqrz
byzYuNUYAWPIdiCL1txFJOwKCQChSS6R4TG01Av6kQF072blDdEMlaXgd6E3d97F+zoUOUBGEcAL
0UvPX4cmMS6EzUu+0pj0YuyHpuPH2TeReZnRZ1X8Kg9/XY8DvieC8A/3JTfhYI1+QeiyQUaduQc/
OBszf1p75Tyv4pL65k+21Pck8ZG5kB2qaer5SKHll6KtNTF+bTOxscMr0chhYw4qcF2JP6QJJwPg
DZCoQF1UqtqgYbnibPfR4q4XxIvrY4sZK+hWwlcmw2kI5SPSWnMjl4jyFL5XbS++wvTH/67y3pp8
64EC8ICs+NM9exQfT4k91MzwS0xnpsvL8mLZKGgjfM3FXGan9sHNrM/xgpmIOAramC0O1tYbk7LS
qOpKrBRa/o07Gq7QgOeSA+JbR/j3AF5tUsxdj4WFiPkP44iYtVsmh8nZZpilc3/8L+BAmvxrecxN
oecflOHr1UGGRf7MNNAlA1HTPUG98otsGEiBOmRjaNwIz8KMLNbsVI+NDGdPlVvnHl2a+MZro6wW
LfUlw6VQmUA7UohKtgpgpCBrzxZWf7leRBa1GA9iIw6n35D0HMtllJpE0+2jV7gJ1V+MYhdLXKRO
EqhYaPica/qakJAQogvAaLzdtwg/BhtnwC7wUDTRx3lZIQn2zBZ9zvmclNmwf6l7ETQS4w8Tjq4r
yHW5A8D6CshVpl+mf/9p/R/3fbqiFtEi7FiCYDPHlCQyH055irjrFf8+eltsURJ440KFUGkLJmvv
5LrFGEtZEwkQgdg30/4TLsrIv7TSSHkf8vazzEuHxYzvYPzMlrkiSJ5ErTLH5rDpy+rZ6cRpxmV/
rbLodi6LLoF7DR8us2ttM28Xgc4q75+IV+1C6v4ZpQCrsUyTlsM7Gx8ilE+1BdvRaBaoMawSufXj
i8nA+JbMBS97z6+pE8RsFJTQX9I0JWSfbsvPwtBuOiab5cw572iqhL3Op/V3mDAcY31WAzZVSVEA
4s7m8BJSUCw5k3oLQD8Ga1Gs7vxLt5F3cyY85eUhTNPmbJQdDrKTGEi5qAc+nsDR6hRXJcd6Rxec
QegXcLORUPoTkiDKoqr+b4YFZ2qfpzGDzPL7LjnG5mhtYgu8tdYFF84+nelKIfKbClrDAhAhHyZr
L+fVKWSUvcwc+JGeS3Ja0KtTRZAw4WzSAMXfzWU0c6uVIag6Vxk8YSGJ3IyhJi+mQTz+KxN5TEEf
j2a0UynRvTqjdhJR0wX41uXUVPmMwd0h+IYIISVMSUoY9rI3lbQwfdnXKqodI856FVTz1Ec8V9JR
+8t77SKk1viF+Y+JiyNE2xayFhqMn6U9nMo8ni5GCkjCqomcapjEpr2AhjHGgOuB+5PN4O2Eaghl
1GAv17hgQrGAl4FMQV6ZBklYvKlarEVww0giE4TrTKUbSNpH2IK1SjyXBprVnKLwylx7BdjP3MxI
NUT/kaDkupYvbpmxx0GIuJeZaSbyX+qwGCM1aIa1hvfWSQxsnNYEPPd7lhDTNwzLJNg8xBGBOe1g
Z6utc4XBlIdgoBftcQJ2z93G905dpfII1Sl+WZO4WgP6fCG0LBRSrLF516wv9EqtCgCHIjSI02Ec
QNfQ/Aw3KjgLpgnt6z8QGZ8qDSppHS3EzKkiZ3Lg+YQMEvDSJ1JbGdHZ/Lu3cSEwXgyFIbr6nzVh
WfWhtdeiKF4OTEUeet9NWZCvmH3yzXmOrHj7IegFXldz3qGs0Gu/S9ZhvUIAMr/ZoIQcnmwh1kcL
DZzjWVblCKRJ4KCJTsqn159pYlQtjQ9gqOkEQKZCF/xRJ/WxgjnwS65/JHuEg8FcswC82AZr7Ima
vnQynOiEy2x5uerQSeFvKQfe9VUDkDvkWKKCBLWm9Z+UCOPRHRriXTnk+hYiqRfXfmUe4pS3PyiB
cevXReaSoIgYAcJogEFx0L6aDUUpA8w/+RSSQfrHbZTzSjoY3lPpxE+ae1MNwuQgZiR84MYU73ET
4OtMQa0V3t7aSoGslQOUqna1vVWeD+H3zcLGfsKxgS3i3k1TT0jTPgo3U2KX1/OmOcK8fUOkxHgN
VBj9xn30hg7EAwsCZIRljVVkeCtcciGQlCV8RKGtw01KJLgoCqRfuBIQYN7t2ctqHiHZeceHpZvD
vm89TwqeZwh3D0tFJ08v6CtwbR4v+QzE1b1inynwaE1W2rW+qOSA3B8iqN0F9ILksFdfCQ6ARaFV
1fUAtZa+wT6lkIEw0z8ABQiyo/Vxor3PGQ5m9ShvRcsIQi1gbhzm57b9L5P19BJSJIQhlF1f5ZK2
NKn8nQvmD2Q4IoUhPFSff0wE3DNefK2GbJTbUA6W5/qCrjrnri1/ISgnLRSjcoB2ePeLMA29L+tq
XzqSKOo9ksVVngkPjl1YrUtIAawnQQMmTOf1Dw/lo4GMexS0o4LxhsJV8DvCchYtvMsmpKqAtaLr
tcWDwCe85op32HtoA89MZ/o8QmsYji8398yrEtT1aLGw6+du1pXbFebuosIVE+YozhVnXcIG2K6G
4OkMvHNmPa2RfAyf6P682NGg/JPdLnsSKNcPtDgSy+6xv3It2C3RnCOPx7NK0McYeQRDBx/z5/Kz
JZCUMwmh4UfT6XQ6iUpzhGfv411kOENqSXSdSJ6NZQp+br1fe/n91IZnSU6ewc/xsLYdhnFx7Peu
NlCZtx/7La0GA/uNEDvX7RyG/0ghTGM8JW9rOFkNKHwAAMl/DxQboSHS/Mrsd9dpZzF0qcQ7LVzo
yFnyCOiAgslRSlYCz6ujIO8XfWmVea+evnRB3zH6d/U0WfHERJmPMBWAaNcTV9SBCSLMC3lttONv
lvKzrLMoFMnfctl4qbs9nz7p4kZBFjMj8wEShMaVLJuFf7aAS4FVlvJpTzs8OI0a/kDpodwbFYwC
jukjZFqfMw9Ieh6Q+4htsZXU4+FEWvBY7r+0Gq7wvCmMcO9VlVYvlBEeHBPXAilrsHk1zE/GoC21
9/dBksfgrM7tmN28DJLmLYO/Kzoz8o3ZoEKwO69uTaGDBUyXVaOtUVv5KolVse2AKfFClZQ7EDYn
D0dJkvqcaMEEJ3uX8DmpsgZhGMHE7yGfpTmC9pk8XlBBRIKSZ5UQop4jWbYlKmoe4uWBoxl9a5Ii
7u402HBf7/dI0pPoYxOq318G9v2Sfp0L7ASNqJQUQHmtlnZD4E6dyXH4X5QuxvFHeLZ0/4kxF4VQ
A/e9960X9YlMRWQd+uI/F27octY9cvD9bPwjhDHAdFZ7UWtjLnpo1ian6b4UdJWUZ6T/XoG/D2Qg
v02/FLlkm4NCUH/3MH9LoLA0JHTGrlcXkW763bSOsiELnGps+9fCc3MymxcBhnjhhCJdezHI4lRm
oQeT+2uz1bK3fEyDJ0lBXlbEstG+RNmvxhG4mEBXqRVeKs2OPCqYSZ0DE1qs3qg8omGG3L93mnbS
+eV8FA1DeIgHK0T7LECw5TdcVI8OG+JeUxiM/FIyZMJ6FOgrtLWuOdSMx0IWLBuNdGDO6H6MJUR+
6XKKoyiuZqgh1QHnbvkMDStoPv36/xGjjbcOJ/iDbZJ/rvVxKaZPqt+ztT0HL6fsRGQAzaHNereg
zfEV6DwzgwTQCEaC6yXMpYwfbnnLZolzYd0/MG5r+Y2SI/BHsaapVczkhNUIxmToJjMb2AxrY3Ca
3ZXQ8aT4uKR3L6X+BSbXjE9rs0u82rhBGfA7JObdrDE+1rNJk79YRX89cOPRSFtSK+qojPq5Jx6p
Q/zWAAd8Cx4XMKrRH9llqZuzIMP4DOS6TWY6+vNeDoy4sw6sx0GEoU1qtt56uwy91rrClm6F6WDF
ZxTci+XD/zILYXwRHUqJt/0ZJihTKPJX6okHQ7h5S20gH+REfMCRS5hwIRP7jI4oOl0AfFRynagN
05P3EZ8OPr4JbH137cCVYJtymB3Rrhg6DcbI/W9iNitFkDMCNRojLmXlGxJPsq2yxplrOjm6HXsv
2hCevOOTuzMRKphW3BR66/nuLnV/vyBeNNEjU3ksj/zFYUoose+zFHzG8Rsvpq6A15wwZwImutQp
4RiZP9JwXKwYeNJZVEsb2GICioAk0hVyqzM8pIZuJXBdADo2VajnYWBfRMntAfGE9nxz5SsB8tUM
8bLJ5uJp0t+PbfAsoBsoAzCrBlV3zSwtBkj0rnZkPPQf6hznbBVQu/aLhiI1RdLI8bfATg93BJ5b
XM8dA+T6COvArTsZvfTSYkWOyirZ8pRwGNG9iB8oBlhMoYnBvNJJP5lDjZNd2OkNedhejeKrZhFc
6hM4ksz8rlcq7rAD5iZ+vezEUBdNvlGpdhuVpVCvFlRSXmHbz007+9+fT3fXvofR405EBHU7UHXp
oXU4K/m/+1NFKZsy/KDe7XS4XZYlFz3MzPDSUyZYNp80hFt1Yczv/Wk8XrTX+vn3Aupw90omw4+g
qRWjNUem9en/FPHLotPxbKgnn8taWEnc1N1rW74B8ds809Sy0/r9PMvXq/Ln/2KH8rFgLdcgaAFJ
XzheYgft3ty7bTHG2nwFVDcQjgphcPTwLOExYwkPUB5zZ7wCUF5E9qOBds+hdxl37AKKdQgvz7bL
PemwCB9/h97JfonQv4suaNyAZhIl12vv6zoiwPf9JI9euiW2IHZYEqZv/uH3SMjXwofR82pRAqD9
LkMKt+0yxDMTVy1mPb/ChpWDtFiRAcvZ20KaWqDxow1mDkFmueE/Dglqw4/+fkmBwfQ/fBTloEEo
bz4s/eEgIIxVRzH8qcETP/Zu6N15h7CQ1wtKpjZuioyS36y7tSU+pzWaqaLv/JrB2Zrwbi74rR2R
oz+c0zlGpFZRI3xt/tuZakxmmduao9RhyHSh4MA0vEMn0mXcdwu1kXfFhxI9zALHt/1t5QkvTFaA
+S8xFilHvs9/JglT0N6eZY9V8noiLGSDSBhMpYUE3S4xfjrv1+6LYIGMJqQLnouElSH4AcEb6O+b
bAAlL/CrJ9Gn9Wbndm2i7RqiOiIkFxu6+XXQatFe4u3fY9GlERKZdtXULG04ddty17TjsTDfsrjp
q7oG/eS3S0TFnfh7sMuQbF/X4kQHX3qIsLm4DRXdEkQ+vm6ZkqnzMpqkHA7lptosbgPjaqUInpI7
OCim1LWkR0C5oJogoyenRfQS3nhheQuFkeNaWw/Eja4UGdU3EBNiz+W9daWp/KwAFotKgIBLLGV7
6Ty7oWm1fU00l39Kfe3EvYxGzC1oF1J3+I+1E6zSv1X+v158ivsP5o6wBzMwGf+woUNWhvuXiW1z
5DB1NpaFSx1qwG6BY/DsG51OnzG5QKutFXmbV3DIFU+kEtPg3KxCmqjWVLrXJzOULo1VT3jTMKeJ
WI5eoZqGPFpPqYf9osXAZV5eCdKX515LGVuuQKaUyOOBZrPDI5oV2wzXnUeyCe0K6JDZvsFSvrk/
QWOAQweTdBzIlmrDk7NTBCaW9qTlmMcgmieJaHbjbPeDj0sKpnEq4T7x+1hUiLaiyXfajEgA5hFN
JEfmOxhpSSiu5BK1jemvMQobn5heaNreKBTx3lsWXENXIAX7ebVwk5DsVBEDACmA/ngW4fd2Xv3y
yHKr3QYqNqBgouk4VmUENQDcCAiC8/VxZyA641d1jP2LbXj6IteSDB7zHGPaarKnrI2sGH60FlBs
v4cBo3pHZZ213FQ+SSVyavWc3L9dmv5fb5VT81flfZTFvI4okz2Sp73a5aQYWfTYvNmDS1egtryH
3Dr9edZUS4AVPORiVB/wZG9vXC6ZaoWNbU8C4rcZzGx4GCvNTHT4ktUkc97VAfOJi6/BNjl7/Ru2
Y8Jc9voFN1G/I6NDQTrzxooqg/p9YwqdFKGPoL3O5zfDUJNdkI8ur3UtWMFTu2B3lG96kRqmXJu+
QKIwqye+yxF0KyZXqmHqd5vorXLYmxmXRFde0UKVBnMkD5zdoE9ViI+M6KA2DbilCiWFOLRetvL3
FYdEcNj1R/t/RtVfCZq7GNrsy5WBc0PIkRm/2gNG0tXXKZtdLJZfL12UduXVPyealhl6OGLbwEVg
J/uPQ00Cn1O8CEJaLzq88hkrWohPAEHETlRU07CBGDj2fMZkookqiJQmoKT6qlizvzXUUNhJmJFZ
XCSpSDUW/0h4UcAH6VSS8QXvz7SFbh798QHP2ODwa6hYIpKIyWC8z4gr8hOOKn07wWWxwPSJCGJp
ge/KXJxm3cNhKCx2w+pql7Z+l1U2lQH/t6/5PLl0Jta4bxa3PSQCpDT+c+pbAHRGlMcjfa57+g/v
cN05j6zjGT4ZMYqgFAIhSSmRvsI5B6xqmj10ixUGX4qUYbJffM+b157hWf1BOrB5nW6rhgjsDnee
1VvvUHe3ZwOQnniZVsa59tH7rFJpggh9ZiQVoKFcPSFmmu4AjZgC5zHHW+kvfQTQcLVnyFabpthN
jAI2Czl+Pwv6vq2xuML+At7ROafp8OIuqmlRSscLJ71YUmwlASd1TmOfBm2kz0eWJW7dKg+vt9F+
xZj5JL8n1IAolqy7cOs07Tnvt5VE1aTkLJrHzOrW4pq7JFfXCx3jHm3cSSWICEcAKP2w2plTDPC3
wCeLj1rbz9FKbTlP4ES2tAnV3hOkAHTnN/aSpBl+xeYhHnXd8wLzHNo7odxr///bEvQ8VvI3t5Zl
5Dgeyf9rzpL/ihS5WBwv+Z1Rv+JgFpL7j3gjdD5Tz2nb5dNzf+hDrNCFK9blQBfWfl6wF4qylTpC
OaiWUx+WVwI/YMXsSYPkOZOjJalYsV+7F+14XGJbx0qOx89X8rCHQ3J1/7kYFq62n3AnH/7EZ2va
haGdB5ryqsoCu7F05BFl4aSc10pfceNelOENV+p9BKYNvMmCO1S+TvobAVhM+E4IEO4O7rj6ymKP
FrmKOFm5HxEXPctKWMqOCSweuwqrzi8BTYFttOTJxC97Ueaa+tjpQo7RmNDB7Z5bYa9Ct+J3Yxp+
yEGQhcVnbiYjm4y7ddfTSqzc+lXEnZNhBoL8X3u3YuuEHglbye2Dt9AkEfab+ztJ5tL+CUfvWAbO
yCN0VbUW13oN8TPt2O0X720uYXajpfE2CJfVNa/Lt8N8UpIREAJiyOILflU+Wu+66baVqQTVF5Um
1Ti5iWbZNypjyqXI5peE0bYV70CD3bPbZY2u9zS5S0sGa3yYrgnuT6ZScXiLQioh0B7ZSf/0vAni
W0yMVgwWKlbGcZl8r0hoB2mhDX4uluxbU4om4KSC7pTzdis1WfaH65UykTX6k9XOFaGnHKFhGUsv
kb/OMcOrooBPOBKX+rrfmgIz9nwH70wcZ/J4k1/QX8gM4zXmA9AlyLwgrW2JjGJsm/Eg9p7n8OoJ
69mmXYmqtt36+P6gN3H2VF78CXcokqNXfBz1OMLeJyuv7KrhKYh0EMG/NLx/fGGjYUBlqWuq4uW/
gAkZePpvSoMvHqVfkF2loQVENWgiGT2P7CU+C1zhhSWK4OJrXb4vH+1wqUzyi1uoT5sbdywWbOSG
lRhCUAeAFpP0oDSDU6/eYQycVrdkVg1Lk4jiqAUnGZGwh3sRyDtyYg+8wvm5PGTxG2Q5HfJ68WWd
QbUf7zMZd1JP6oVzjrQeqJU5qAKckafOxV0IWjcttQTaUNkm7FB2WTdcrQ/LOVnofyFHF8ZOK1Tb
nIm4pl0a9C0qWsKVufcaLy3mXuwIJ7RHTZwRc5xtZTTlYpx4p/4HK2TDs+BYWX1ikhb8xlG1MfC6
wOMKifPt8FjGXHCQRkFfDcq5eqI+U6qPKtwJIZw3i7GVyExaqq542LX+23m6YNdVbw32qziZvb0N
F3IIoqu58GLFm6oSXQf0RWVPhyJNL6M4QNwqwaa1pykkagWWJZcOdfQKwvZ9s1RBaFxeExnKrKLv
8jVXkwniFKyf2lTn5iQ/mYRMz/zk/5c/NgsZr+eNVuYgdr/J4rVqWIfLSuHy1kn3T6njfNQDQhoq
quOkWUo/DpAMtN556WDglGG0P2QwXBSULteV4C1iwAG/a0XPU7jYANvKHj4hrYBbbvnD1qZOflvu
a5nFGMZEv3ebBRT3/Z8MqrU9CNp/tu49xR9E4Y0YV6MKhEU6etcnQxG+jFsDwXh+C34Ro04ulJ1a
HcyCRFFR/M3PWik3AjCPo1xrtugPsS4hx8RXXzFg+/wB5IboYL82W/mnHhxpRKd+L2xS2U+c23Nn
GfcmMyi7PUhZXRpP+xh6DqkuVcnbu+E7DUgtjHOCqUq38I33B8TcFpZhthqnOlVxUf3inhHx83on
6eqm78E8/eq0hUkeqZzrsYvk+S6KRjs2nbr9SYKMVFLcF0H7lEZybr1+uvhZO2GcNki9LmCCvyrD
3m8v46xpowgaLk/reCZ+iyBlzYtYXVgtExKGOe1iZNlAlJadVB0JHm+q9YNWTEw1yl+wnBhWMZDB
tX3oxpxE9xGF3C04qFh1n8zoaxIH1cDGswoqtMIuXRKe8aN21ODy4cHobz6wmnfTsct7tTucSD1/
yDrtBbAV8DXTDBGpOzcMpJXfs2VHZPRU4+XE4TSZWzRwaveOKd9Bjge+nx65lQup1evb76Iil2iI
k7J0XBvoipHu4HlpI0Gt626g3/W/vQqu4Xbehs8n1IB/bDFqpUhpE/19r3sCTSrn5cDLyche2gi7
Cy8AiS75BUcrH3XO4Gb0jRbd6zUWkNDeWQO5SOFjjPKXnWs/G9Mwzc8ZbQ4i/zOoT/M5hoRSg3x1
RoPlUW8zDifLcaYRnD9Vszabtp9X8q0R257yjyxZuEqxNkkXsSjn6HSCTpA6KSpQvg0tlA6/AVpY
6+0IlbLEOLHmKkdsOJxaWAWyd4Gz4kvrBFNs6z0XEQSWBOSj8ui7miMlFNLbmSrfEGoz9dbwb6Xe
y26FXpGBJ99d4bQyvIIEolZ+hJqPtD6I32Hd+EOQs9tECDaNLBe8bJ3ScsBTABg8L6piw8kFEpjO
5AtUVZOn612zYyRAdFLnQWe5RslIjGS4RQUBktWHCbWLwjtzCHhcr57zOwFS+kn9ITpoo0B7GbRP
OdrftOIz5AwpuTyRh4qhjTyZbWCgG/FlQgygQXJM8u4ngkN1WIPFGCOD+LRrf8xg9wNXDAQifSOP
1n/KgbwmYeNf3JnRcRARU0/hsRO2iQKhRHVW+pUVx1B9QdK0QzufSVDk8IuLUf+1BZQ9W8Zf/blT
xPVS+xeDv3SKRGOsDAOggcbEu7fyB0KiPFeoRDSQm+pVPF5dINiYrhACMkhZH18zvzHOTUoEkcVa
BGxr1ZDFhCm0U/n8JlGqklu6oPzBQETjLAb0QoRy4j/tNdEjSZAosKYahyd7Ywtz39K+e7ZOUjQN
hehpxC/1X8lWTHmRgUe0opzOhhQZqm48/sxqneOwemYcKGjzfqpnTGFjbHwxzlIDhgBGupvGl+rE
c4n0LDgYG2zbaQYtVKwCyidGQCldWEdUcnQwbRtSMNxbLD6b8MaM5NpWOoKglyez7hqlU7uUxxhS
8kdMFh6n5Rqdb+cKDGGnnqUqBHWWc7LS10RGJklX84imv4m0iXYksWlldMzNjrzaRZrRQaCJyGY3
DGjJbPlKAwLBBmLv6CrldudGexstYJX5n2kjpu7mSuq15oeehjA5wwQx845hC38UjrELosd/IHl6
mA62pNInbKrXA1mbILpR1inRMWZaHkX2wTlbGgxWUkMDBSwJnlt+5cuJKGLUSMSUK8UnWo7IbwbL
HL2zzaHKVVALcWSNEybOgA/g01lHBeYDHJUDib5zWFdfeK5WUyM2HT7otsULKQ0+xS1HV9z9z3sY
QDMvlPEgONe+5kz4gFwaXgwQlCdny09UdCbYeXbdE5VH9xhdPpnrDG/e+8FoDM+zR7+zzmlz2FMg
sC0kBNOExCoNGqFkWZZm4kate+T+/Ks9Kr9bfELMBwP/p+2IgsVA4GPAh35qwuXoS7sTc7iSBtl8
8ERb2QQqKw0zSQ1vfz6lGnuwW7hciZn9lqekV/FMNwV3bIs3Eaex7LJoCj+coDvQUTsa2QqPYJZ+
0XS8tl2f5oIBmrpsey0jKRz7gUjodF9+H4nzmmz7EKFteQiuqn+ksFtvAkdtIlZdqieCyKyL9AaD
5kFzDCHn2oT9kDsMQdsP9Zs31P2m+3K8TzgKQ1AmSWn1fmIlhzQ1yvNerGKUB/hxLJegl2MqhC3E
3uDN/fERFiEiojVXKUxBrqG+U9f5kIa52tX8w3iS8y3RTIslpHo1npSAbNrwbXG07nYiHOKW4vdB
lpc0IIjL8s6ob0JZ6vzNhJITm9oMGOCiC/h0+goXlXNnVW6977VBd8p+1d23jXqeiubetT/IWCoH
ATGImjqgtEVhnILMu1xrdobU5PVnaYOzs78GpCBIYIKW/3Nv1xULgYDhhOQVBAX4eBB+CHfNOFMN
2XOBSTLs7dl0d1jtOzAJMHYj3liYp3zqoX66hjiOSy91UWIJ0j0EvAEBDkbzZLDw901x1hChFhbM
2Esu71koru0CMCB5egrNU1K9KR+TIetO1esOgFRugkiFp72Tsm+YNjdYp2POQlHhXMXcwGlyVldn
SsZhlC/WeQkM3ud03T+tfU1vF2Umny91KjGow9BNT+IZk6Om5PNmfZ+QPJEoAIS8IqB52mEugosE
52uiVDEzfGqyiESRi1obTQ+ckPI3ZOCC3Xrhe3TVP84bThevc0Wae7vXNWcMKuQYD6J6psw8EDng
IBm4BkDkQNLyj1gU7wCkzwgEBkEQEAZzvZvY3jjxupH6lI6y9zqz9eilen7fX37YgQRubWf9O19N
9QewXSI3/Zl/B8G7TZGyRLrVhh3CJH8DszrYU8fYJ2Db36VdLeqBQmV9dIh7+I1MgvF9/jGpz9iS
Cbu7ClIW2b36MTpLUCt59JivTgeJt2tBRw2LLrPzd/MKkeyyP8B28xj10iuLGL8CmbfVdgmWd/Ji
1aYUP4jxgoOIH1JbwE5q7eaT1wZmI2nozOgKNpVVTJapHOPgRvDlqTA6GpuDd7vHxR7pRH2Cim2w
5B1MiZzO8d1r2JWSLi5XMrgIMFehQ0d21ZgPeWX+s1IP7Ysh7yppE6u9pw8RaJYFAnQH6QR3rhuV
b5g2XQEwE+g6Fl+YD4u4UOZpbjiLrBniRy1x0Q2HCSwryfXR8SBNigu10dvHQc38XhVEcCKdZnn4
dTL7o0DVHRghd+LYeKJntl6C+AuK9+u4UegwEIc/ec6+8VKzDdu+yaaa6j+FSCEV/Mg+cU3LwyMH
GxZfP7uaAYGhktgBYH/PVlsrPLpsu2E82cIT5ANR6JD9CKnY7enne35+iB0T9vy59bPg09Wfv8qE
fgN3Hyszme1QGALbMucuraI1BY7U2g5ki8cb8TZMxXf0POas9f/PTbpij+LJvB3UjapETJmtD0ze
EArbsvnTl/dyorY2yLsEVWGASWqfi/Q1RzPILR49FJUOon+jO1VMzV5lPhzHgyzA39ZEZaaSBUy4
Ls8SKSiLVa84L/Hlbf7a29LDqbjfDUOvF0y1LSUvLwXxqQwqrGFnok+RHx8KZm1Q8Ztc4fRLK+PJ
lPTj51fkqM4Hdpsmgdmy4RzriatOhTml4G+KmdA5HnmJL4TUE58ty6Z2RTkC+Fx+yjA8UwlZSP5W
ZguVl7kdYvPqOnQcH4/0hIbuA96KkOD+ePuhdI97zvCawvD9NsHilc8Rij8JkPzqcEP1mJ2J2y5L
mlSPCoeb6em1y3StasXo+eaF/OFsgxJCV9Lw8b/CRyPT3tzhYe6IhKhHNNnWidcamNMJZT7PvFv0
60wIOEVEUq5hJU22HT8qi++V3+I3SPmn0x6uGn3wAKq9NWa/zMTnzxC2LrGBjLVLP9CQRluE8jZl
SjIViqHrvG0s1z6e17fgPCPQChFXqu3rmwJ4EL1x3gjdM5NOaJo2WVwqOkNvi3tpkq8OLbI6tWXQ
9IkeVzI/KBu5cJc++Z2Vq/bnOfbZmdlo/pGN9QSSrCvnqh2oPpnk2P8qz2dpkAAM5PNf4vdybLiE
IyTBm4odOZzTzsAL6U5RMgqOz4PkNImBKmncSnl+/hw3vagtmmHoLcI2QhobtTDZIi7r3nW+em6u
7Zg1rbaMGdm8scq5MyCbj180zeRA/g78z+czpRqSCQaqNyfnw4R2Z19t5O+Gh0CPj6fm4VGDHXhP
lzFeMXtvLsIy8XpICUUTY9iBeMTQ6ncKP0f5rdgD72J5dVTKlUaCugRiTl/azXjsmQqneP1Ejv/s
zLI+uBHJD3ojmUcRvWOQaV2dVVF7dxuP2s9Rprbo5+MCtu2RC8KTJCbAhqJAwOsgsc2UyWfNE7A1
aQ4Ssiz6tFYBDR503s1+o29VSj9DUbdGqMhEmxWJ3airmikYmMe6uDmm/j+vbf7otBLtgPvOxobs
/4ngjp0wmlxdW917aHqvS8yeto0Q3szkRq89BSS0TmcuX5mPf7xuK9H2KDJeuuMiwWIsfg8EIl35
5V1tHjOrmhBKFOAF64APH4dceB99QEfhpb2xfYlz1umSO2y24RteIa/9JBRgRO4xf8W2XmjAfWmG
aYJFenHjaCtEtlmYxoqcUlyENSdK84ipa9PPTu4Wll+kJHeVC9iKQEiBYPP8J35ZCZYaYaFobWcg
SltWo2rTJ4k0zPmFOlK7NuloebxzOSfShI26xxzeDUBqt0Y5P7ceIe0pEyOla3Pc8dVY+uXoD8QS
wpeDC6hQm5eYcCj73tpx/UdA6KqBuWD/TR3m9b+DfOEzJUIQDOUuN9kOv0xBz2u2wD1iXGhgEI8o
99l+VjR75otb6QBTYI4x1qnr/DfOUrTV+iRBQgIUA5kchXqKWTJ4OfSkZWVkwAH7JjutqvLH+VXV
7uucHHmG/oYJhJfbrYCUegWe69FXXbnEjElawPRjlDgJubMkPceEshNE0EkcDkUSsYUdHnbeTuja
T1GeigyETlXN1ZgT7frsaeckvHnib7O8ySPA7bUQce4UXj9CNLBiHnuj+DQ7Qr9I9JcOr+mNk6Av
K4dHecJfQA3L/G3hqNQOqEHoiKo5qpERLAWjb0p5YmL7ZbVIlTnOYj5eDLg8VigvcFiOR045MFpS
/9KirWqH3GuSI2gWjXHhvqNQWAB7gFdczLDpOUZYFtTlfXw5b9zKBgNqkVXhX6Du5pkRjOIRtKGX
NKIrdvZTGfOP9Ja/vj1kvGFwEhs83y28uYHBuWU/WQ2H5Hp12t/mEw/CO4Zydrkd2VeUlsqopHBZ
LdP3dWxR0HZvDhiK0gnqQO4g7y23sSVsv3L4AF14Zyp1pThUOO1rAuzVLOoth4BbOtzdKK1LBzR8
C15TISDSLTZlnao3jOoal3vju7Vw3Z1rxjMpDOEHmEWUsJVuUkww5J0fo4MeJ5IIbWwsIAWnGIKL
FMUneHFsYlj/GUxbuxBfV+5mei83Q2/V+X8JW5SDu4TmpYL3EIKomc3fAu9SLCrEgS5z/4huqnGU
9Nswb7oaLRxX2CW029c2/CbBoJABAez6kZkMpSYjZ16h4o6qEUxclVmgoL+Kn6lGIcKu3FRvpLE7
iDcmW2sHLc6Pg82zB0mf414VWTmeaD1/8WlRFbkvaW22G8pRENwz9JRw2pQCSx6UGhJJVi5oXhR8
g/tNvA+lAIDT/eXf1dPmGxsXapu/VLazvhJz+ecinsaJUvKNgP7AcbEwzrK3VEgBFlPZjxE8FV4k
JdbX8vL+q4bWHgl9O/yjidQUu9F6LTtWl4OpOvkP/wwVqh4kLc1ZKFyf7rOkIWuMVQh4R+ud0lBT
aRVsrKentrfZVVUAt4SgPlTzWHwkOtss8FBCBy1Jvee6E6fKlwH1ixAKdHJwurpyc+KheAJYaGEX
zfpLBGdqvsDNqXDQ+pQLo13vm8e+pzDjmuFiPt+xSSUTC8FCgZDA7MRi3J6mXIW28kWDHNlVQhHH
VqWmbvczi5lhyk2KHNasSIITsH1EAdBtFEJZxXss2Z6OLreAkujgcPeJsyBMXQwW7I7rSmyO0+Mx
tGgMSJltgjYrr5AmWgwsCZh1wbqwwwESEitzaHh6rdgplaGM8hV5Zx5nHTazYkd8GIN7G8QunnMF
TAms4fI62IRVhaWuhwpW/wIET50rFFV2aQyP5MIT2HSpYfSAb/wyhz2KLksBl0NdxHsSHUOuArL/
R8JSmPFZb5TV9v4x0idcH+M8/VteojcMz+05fHTZS4tipqWVg8QbYzAjJ6nCdTL6smjZ49f0IIgb
Xl0cPO37E/ef91GbWfDtx65Rh5NdkKMBmLatDHQSpr7S4PlDkdaVvrNTlBx9Qp/NkGcTp/CFXzOA
qZyAE1yhdJocX7m2M2weFFFyjGupJYcEiCXuE7YdYgLTqV4NFx8G3NCSUiyKKmzDhc0vYpCpDtKj
UABnH2EVrMh+hOdku9MRqCAI+R2VKXw1G5+99UTKIqNk8d81DD7NgLsB4iKFdifp6HHUS+EtwCqW
dinOMWVUOzR9rXOJ67jmck1m8da1Sj2yJD9vNU7Q12a+qGXBTPxNKCbMSfARHH4Qzx+LxhIIiEbJ
bpYrsbkwavWjTt82YfT1iZUgQUGh+2xCgHyk39yMttTKvPECmv0ZFQofjmKswlZFsyNWxhCpC8va
/PxaqRr6rRmaBXb1PKyCES64bJp8bVrI6BZQ9ov/pC/ecYiVI3WI++ulzKMtvDAOQ7WGSxaeVImS
JEm3YXT7aUNYFExS6Q+VQnrngi/+qFsZeQf+Q/jJAAZqsVW8D/xzbl/Fy1WHknm5I1lbqfniG+S9
VH7zfz1kf0T5OcrjDh4kwh7QSw8pZ8uQgLSyIR5SAm01DkbwYkeKEnY48kBnMM7B406NVyNBk/Gl
X+vQo7ebHiBN2ccffu71FUBVnWZNWCo1eMfviryPXRhVDais5+eOXVWXMcs1srI6z527Xzw/vxL8
bUDVsiRPwRZ26zroYrJTmPG3KPdrN0VL58KnxjYyQ5sv8OgESGGwRQKX6IUVRyrdtzwN/Moo7aRu
D0vvDYsSCc0rE2bJAA4c62bqKWlEswZkwZkqfAh9EV55nzpc+jiTKmx4A9dkoRM6BqLLptpDB0t7
FOoQln9d3KovV+NOaas5RDhhMIL8wpnqMI3AheOIRUNF1Snk5Jf5TEs83iYExfB1Y30zwsa94JDD
a4WdMt13WRvLuGw4oU2sg+Jjzagx8xtWrYilnG4fQX3l0nlHgoW1VWPUPpLHGn5JpbrADk/nIJAk
NYV954+t2CpuPAlKdb7cO7OTN7rbYxsNY8A3kLHkRQnTC+fTUpS1PFJ8W57bLC9J6Ck5/cL8WXM3
N2r9dcBMFJIljltp0lrBmdDWhVY1llxo+9h52+mNqnevWHEGt+m//kLqNw0XJW3CWGqqNayZOt1T
pkg/7Bg7sk/NhBCsb3HJ8HOkqHAt936TL4nPKpPyIt5RyYLOt2IbKSXIPOt848fqVwjNv636qgRi
WL4nXOFG1a+6dkOsNhab+P0Lg8X0zObT22KD+NmM3Sz4FT4nuwYgHJH1Jm1M/iObGdFaw7v2KuRT
iTg2IGQncxmXmzpS1j9Ksq472wDAAJc+KKt63riu7/+yCTSS//eb7jmQEU8yc2Wa/osRMSz6bT/Z
NBaFg5xR3OfinWrUZk6lcCFXluTGM7sOm1NUQA/R6lM++juZ2aLGyKCPOnQ63qfmn+rb7gT7D0A6
uWgqaSY/6wtHzwBTTcqD7dJ6291QXiYZQEfZ7YI4wkXMlxCz4+O/sE7tgiZgtZFNftHzog82Wopa
06Bo5CiqePoZSoCQ7y3H5aPreAkKDoXHo74lmUbQRqyegPeCY3X9mSSqECW+TgGVs/rpFQaCa4X+
IZl7j2P6gt13tdvpz6PmoUWnjTspp3mkbj/SlpmSlledPLccKAg6ChsOSb5h0ncFo38vnEP8t5H8
myhMZPQtcfuG14Umo6bNRdRibSM+RNjb2cJ8X7dLXBw9QRQuldefaQOuxqGt7qE7HrIL73O9jshF
gCgXrS7nLKUV2GwPhmbqWPLdOVvEI40izTG4d7+Mve/ivpZCJUuQmomypY9QMf2eYzVW4wG6TRDB
Zn8m0BJDQlhL93M5w/nnQw7moAcJj42BNr6OV1Wf0jEtgvZ5YvVakgy3HpBZ4TZz82Y4FzuEHa+/
rbgeDUKEBj43uPRADvtv0reKxvpRMnQDvdue5XIuFKGKCX6oFh064oWRaegVvRsjFka4xasNYlhD
2MjMUhWFETWFnjLaNLBBC/SQdZq0d/1+GkE/wOb6OFwq1fqqw7RizJepzxqirzPHCHgfTr+JXb0F
EaJ6fs6SQux0ohqhmbzIkzcvUY6JVojT80E/d3RJ/me88SDpPli4l1KgFSLYab0BAI7pBnie6VjP
3U9uYTbp3BEW8/S14uul+1FjiS50PtCNM/JfoK+Ledp994BsUDOg2KlVDnjN4ZXbgGZe+SJu/yS0
AwiZNjT8OPOwzvbZGleenR1GuXEIZWgCqD7LfoYsVDTZeqF253EO8PuPB8LII9Dlx5HpspqV3GXB
C2c0IveKXi/PT4/WGcq4gxFJD4mYeQF2gWU6FLykMMufzLPvYPjzLPzeGE+VBURtbhnH5XKU0y3F
oxIAItwnAR/rPhgvwmjG+pcLQoSLwEof7fyvAt637QPFslxpGdi9Cst1nnp1pIMJaqbxIspUAN45
C7aitgN7BrvHd/KC3L0El3mKsq9rtnnUeC3/RJIXffYe2TmeuUY4aDn4Focp7khq4cfVNaLiJYN2
EqKmusOaMTQJ+aCARcxglh+QjFsVWoQqn5sGwiRTqCgW4MJjgpMnTyr2AckNrSuVVfmBlSHYoOBx
S74Sc9Dt6GCbr/VrmcvS1RYxZ/b9f/0Ym/98KltMJQqPXiblEZpYvgaPs4zYxZI4T1wElVOwHimz
gjzv4zNNKeknBLokAGZzVhGjP9I2T2Eh6U51YM4UdCxKYfhQfy24Ajbr1xYl1Mj1Oga6GFRnxe7G
u02yl8FcIKmNIRPGLV+XZHrpA9u0e0KzlA+3xGThrbqXhXdy1558sMmuFL9C8IYISei9ni1f4g2E
JaFjyqovBd5PQf8WPIXsvdbxQ8O1qTnzRcoeHUcr3Urcmiq/Fy7Ago/64uNzQrfjy9dfPe0gArfZ
vVswEQSuSXUVO2tZV3x+fDvPIzju5k8ZFVAbFkfySAEOAHBInLwwIZJ2wiWgvv72CvQo5t2uhH0F
w+qrpesUcEc+xHMR/kJqX2DEB1ov/cipDBETpvMjzMOdcy/G+e3B9r+Hotl92p0sIgJqYAZ3jL1x
n8AVRGHaLDbH+vPf9RZMw5kCjjaevuD6ZdVE5Pow+KRSV3+axfYdJ2B8L9lMjBxNcrOMInwLO0lg
l1UiyaZqr4XH2OUqN27GlXW/Nc3SMyLCaH+Ksn87CneXJWGy/0QVA+0VkNz+0G+Ps0aQ3K+XbvD+
eubt5Uil8agdAXrKtR91W1PB+cb4BV09/uK+K6Qt7Y7Garu33v+R2zdHBnhNrGBp7P7nDobEcnUr
ZTOhORnhKkkVb2NkVLVkmhqN29onFG6i5/1N4BxblwxRBqrMzkWuO6DwrnKvJR8/nszrw/D1rzs0
df1Gu+wIcUX+jNBLLM6WO3U6nFlVAEAGV3sWAIwbMvgA8RQLR9YVDkjAqNsnJpyMqodYW3tDpUyy
5k3+HAGeyfV59N6fYAKNEUtJWFviNrmpr8LUt2JIQoEQhJNk/X/OlKc82WxMZPiQQUifR5Bt2e/x
gcE1mPjiLiR5b2KWGbXAmKXv9EfUs0faykXvrh9OuuB9Mvod3DHXAl7AYRgGc1rLmeJWCmTiwzoz
cqn8oiXKQ22VOGlO1j3IHA437QEta8T6mKSwLBPqTBkxaJgAlaWQQmqcVOkqc6+zwOd8pFgpfsj3
Vgl6FuwGtQcL6xqwqsb3e2COUhciQd//Z5vLvXbk2mQBSrsn+dxbv9urbh95Vy9V7vgbjTfPWk9E
HUmj6+drGmOiNtY8gubvbSmOHNlr4oW9t2wvleoenknJ/xd1Rk/VtAUV/74tKftO39qCaOMXQWcw
+J8cajlzqynP+b4IBRzCoM7v00ub4u4qmHKJqV+aGA1BoQqDasWKSop/uBJ9KqilBeynFhZaG7PW
KE8skNfBFt3iACinuPh22kGeyRd7eX38Fy60uriJ5XstVsDvKM8TQJV+rJ23Yh/seUBNXsWsjzLP
yZ7iOMqjd8wUdr2UQW6ptY58I41//aq5pEAWC293gayBDE8po2uSDvkyHnhcBXYLOkl6hyKBhm2e
wM12sB7FuR0dCTZzqgddSzA0z1Kuo68ersv6XbTV+o0a/j9co+Fn+sIcYnQ9elh9Jp9FiI94/Lkq
wO0kehCxu/TLsXxznb82FcEEATgWgWOf+irXFXlMXR2K2CTcCDgi52kTn9davd6qJ2WLXjEM7Amo
Lbzxr+B5CyGECcaYrKdISHa216s5RW61F+F9w0xDdTc8mw67tZoH3ezXrB756iyLBcduvmaeSwsR
gRq91zjmW+Mc4VhGqJKC5wdZZWVUpcsgKgKmjYwU81/tzklRSjzo4j6kruWbncukrENeAzAcmu0N
rgW+XEDu6NMPGElx426oLbKsGPUblUORUewPhiqiSh/i7Bg59+FJjnS6aVw2sVqlr/lqyEFP5bSC
aYQvu873iXh5qYX4Dr8lo8lxuJnkoGSCwAxoGSqyyWd5Tpf7lstwAVqdecTLGfT44s/WY96fIEyH
fUeqxTf53hW56F/RS74GlP8fy/Ru4/mWiM2BiXVbBsf9vPeaTVbFxN+zLvqvO4zllfWgy9P6K/fW
bHqzH9gxCMC/sQdwl6qfsatMdO1g0US/jSZBz28SF1EVKgB6uaue2uLQ4/bWaH4fQiUaUmG1QOny
UmD/lROCqG/XhETIDLZIcGpZHeNHvSUr+PM6rUB/XgLyB+ko7bP+t3tEyWtZPEl+Lxf+nDPJsEbB
K0Me3e58lvsondjcUP6hlU4S99yRS9RiN15aotNH1EQIsd9yBcB4efBKqvdtMJB8TESeKNN/TzY5
Ehgq7xAb2v/No2KAF3CQk3M9Hyhu7RCYf6jhfB7aUqdcpndT8JHjSfL2H8W7rHKOsoxwMUXV2jMG
yxD/6xgpXE5RkV6uxgNRU3E9VGvZGWhZkqLMMJoNB6AJ44rBhTJ3WzxZRuQbNLO07OX95GcSrKeo
dfOjPYZCIcGJi2nllKLwqJMrdGhGuINyxtZ9mQ4pQxBc9jnvMgcyhXu3AZ8mj39eRaXG2PqfitLD
rPHE5HTb9qZE2gZaMn/Iw79b/kF4E0L3TSmnmG7+zVqunpJ5bP5B0iaXDYTMFi8ZPoiZVwUHWNIz
7IxiOdVcAKiMC90PzPYuHuBhiEYvQdk7Wtk+3q+Nflx6xj9hETYY32gpumNb+I/lxOr/i8axwQ3L
Sv3ff1y7+b6u8pgVYiADTdz6SZVc747W0FMWFiJzMqF++56cBpWw+7NLM2PJdYdN2I6E6CEp5Eep
ch5tKPmxfR2xAg05v+iJCATUi7KveBnfx5sMdjhaYnRX2F23YAgLT2mf3LEYfq4IkY64Ch9K9rGv
+XCfwTZq96U80/RRYn5cRoGO4EBwr8Y8Xu8rdmgoNwI8179LWKO58K/ErtDxl3RMK5N8obCRDyX2
yxuNQb1VmDrydr/ZW8ujGFCY6NdtqsEfhsKAl7KyikUAoh3ZzQqipqQpy9tvsIrBrhJgurUzI3UW
8fQqb4eBo6sAEQV6udgw3d9sZ27rTlTZovnOP467CExVzRFoeAloFIQu7+Dj/VBSsqB1JyA+xtky
Zwezi3NUARTfvuNO1pRVGLNZuqhA+qFD9si/c9zW9pkqGuAkgn9r3Ttan21vYK9dihNZYTcDQU/1
2UYTIazaGaNS8Y7Hq/hsjxMpjfGFI7vJKWF+up+NcPmLGgJGHNN++zHLZ1QL4t5i8NuXo7yO9pjb
DKHjA1fZs7CqO/tH+7QBzonrViD1maXJtx99bdUlR1cOby4CXhVbY+jlkkUR3214FGAXyIXiZtWd
KUVLcjuNZXpKNjUHnE9BhmSiyReIeq+SVjKo1Eavwa+vo1MxS/vwPgaZuDvfnHffKb3Mm4kaH3PY
UZiv2cJRCzmOwLooG089ddT1MIEhMMQF8HhZUxo/rjJ628BNHIZ4PHlP+mtOYqvakpdB4ZeQ2oL7
u3kX+Go0h5GuGSZ3AMscffCm2ExHw3D+MACETYUNwxWSpi2r2t1n7VQssMTtmhp5UMEMNoSL7oU/
GA6YIEe6NPlYtpu3STydj/83Ntc7+KuU2lAg8ZTyOvtthsmqOpP4wFsLYSW5cXj4MrklBWQj9mB7
vay/MUQtIcjkH5fq6kEDDPfpAfrI7Jvawhr25USfl7n2lOhKeW9Mn/vst9/RFx3knCdKoX4MJoPP
j6fhK68M7SUIyHhxM29dIvtxCiEVyhnDXvTc9HPmVjTSpDFHK2bd5IuA1WXWucapOYFKtYccU+8g
OYsSHMAtwY1RpAM5/mFRR5aQmWdxQnz1RfhVedKAkW0AC+HropwTM9rKKZhiH4sdEy6wuXjjLOt/
3ULo/QjW5hBLRASl+LAFvpjjtBm4YS8w9nZ/Fl3YhIhMjV7009zY6REvvn1meXfODERaikfodWkz
WdXeCRjipgVGIpZVB3qdfQppQNEFKphwrG+wbopF1jNJsFhjpra5xCuILL/tLFP+huN+mJraOT9e
nH42NmXtoKjmy/2TxoXatJ8I9tr0fmKwvnWq7h++Zso14xObz5kTtjI0gK+iMn4vzbFxzA++I/Oc
KXbMsPfP39pJvc3NvRJy+P7JLfn4kxVvhYoQB/eGvKOisodNteqYfhCD+sNWvKxv5J0jSI8Gx+KQ
ZUbTiD88MIfPpofnoWi+OA4Za7JyHa5prX5LWjak+YNOzlopy1OHD+lxdLCy70tmci0mIhZpDD0y
0pcKCmc8MmEbGUqYAn1CemmInxa5hiD+TJw4W6hGxerTyVjpitKHmPcHHgh6PcKeek3Dwzw1nEoP
cRe8z3wfyZYqkNCz5nhV2rIckOQlYopkHRxIyp6We38TE0rZlxWmkxVVMQdRfChc+k/PNIMvKrar
jcwHkkIIYM1kKz4o3PlxKkaFW2hav621QjtHEQt8bAeAJX+mZ90qkLL8H+LEP0EoRWhavNLaYlCg
3FKh+wSprqi9h98U1awfeibMZ4s8b300440PjygdDc43qwZaOz9z/vti4H5KiN4+2eCXBpu2DCWy
/4j7TThWfo72v2jtHY2GG8HpjRPx+9E8hSWBKZFy2yUWSN3zHWH7f81N3waE6QqdKumDytISOhKA
r0g7m6AOC+E+UcSgoWUMV/Wt4XLXUgcz+EZyfjLQW8nXD1dDZDgdqMYATsrBNN+ZzUJB5OvLNjkx
sW2tWfdz6bMz2UfCAf5xZSfj22hdbwVGfCjL51mSkJaw/K+O3IT0+BioBWIP42biQ3wdOgViIOr/
ULd6RFIqhejY0GqoTYRrB8NZ9n7A+AmS3o126Ps9Z5X0t6RltMF9w9lcKGimHbteNC21sf22WxUz
iygxFizEU5ThHpvWKlHD0NJf6FG5R27JgJKwX0UawFd6iIls2XEw5Wwaj1HIF/9SVmhjKNVTNhNA
1EueGvc1CgO/I8QoJmN+I5gCUVmRruYYANoROq9TNr45SiMvqaou2MXdzVVnJgzU7IIGPfiE7Qld
x771UGfMyqH3ytm13LZ3rOogT0AZ+qW8GGdrhC2H4eR5SpaC/T9VfNFZUiTkHMJXiag0bFQ/C3Ax
w9pxGQkRoi2sivIRkKFagtUbvbAVeLgm6r9Fcj4SYnw6QSbuV7ZUBTeqCCflQx54qZYmoGeTHvtG
UL4XEwQtfhMZ0kCxqZY9Zb79skamMFGTeFVTNWD8N2ZcAMgBPRCbFEsMrBvT0autRfFrH8i38ddi
dymCvOSWno9N7mSeJJx2gDHIbcVoBdZyKwCCgoSHzx9g7CwKTlVkYIdq/IN8DAhdmv4rXCTSMgRt
YeOyWLGB+7DsmEPv1xm3vD7gSQ/N/B4pHoxZ4d05ksxbQmT0LMYJGh/e0z7FnU55+UKLSupBZHLU
rYB50H+W84Hyd974hUE4mD1IrHHhPj529V4876MAm2dzWjiNore00JdyzbyGUprRsQOdrSACuxPQ
b4+7Gj2hqMzitWM4ioDCYts8/yQupCrkk7CGLDOhh9dvpSK+WCddhkLYCO4XWQUPJxSQ305bQxO7
XiYpgrm16TZlFMnBsvoUhgtwHf8+zHJbk0uWjpfkftA5ecLFMwx8W377G2X0M+UpLBQ26ImvIpAL
qvd8qCYOcaZIDqALmclS8yIggkaMaA/zXq8I4MxQdxbl9RUzCjPBlZWRrUcJenIn4Pvq8uTkXWvw
w8a3YTbQwjOlf+/51O0htp0HaSnU/hvIAcE9L6LAn32KkUTs20BJrsY8EU3hCZBERl/Mt9ldDqmg
dHASgD8+CuqEeELhKnGmdcCP0MCnaNaeiFKAi84zFpxOtLQ+5QYe8hAUZu234W5iyTCgGn6i2kEX
FHdpTO1rBa7Dw+svkYB7cr7lcHVxLKch0Jy5YWY1+IR9qm9raAC464/LpmKwC+mCWaXiEJdeADqg
b/x5nAkhFlEO00UKu2fg0SEndS6HtbXEHPjp5KeHmmun981it+3J+QoGW/9tqSs3sJvlYbGA6i40
540n7tun2TtMg9Yqt2H1dVIL1oh4rc8VXuPXW35/Cr6dF4b/LRwid0L0CaDYjv/4CbXXcyZkReEI
O/tydibE3SyKRLAPcJvpcJ0JuglA9kXxDvsexl7hhCsuPspBtKyWqnu0NTnQeA5d9WsCYRbdDiJ5
YQ8BxBgRerWZRECKog8XvjWvuzKzIMbEyiovKDshRl7c5oqeg7kR+6esLLOmUUuNPR6gFjoRZ1Uj
KHTr9eiFzy0ybAPSpUQ0yOISKwZNgE6pcJ3rY+WQINUQ/2fNTyTTcf2CROjLstGcB66lldNeMBW7
H5AJ1vvq5e9indjK9rFEgIuvQoZmZ9av4zeR3rfXd9ZzenaFuv0KJm9MCNQ6XmQrcZ9ympK8SO5B
mHsAylOy8Daomo31g1oLEJE1E71rnriXGjExjNQWq+yotkagblN7pnuKcp2GfAQ2mUYqTf3Fwil+
tnOT+QX3HIqkaW+5nvXhlNinxyyTtBcJgemXpb2geXWALKjvtPG725JxC5B0Rp3fL4LwTK0iEsjJ
k6My83jra1/f3TE5ZFxqCmIlq6CCo8KkaTNnidI/0mpjJJfVccG8aIXd9rTYat1HL0s696H1qOvj
1Q2eduO4BGShevKWQhLlzAsAwlDmxjTU8EXTEQFaffMTKkYHzXYq6CrMyIgL4Bvb84GI1r8aqgRY
zxiErs06AwQa5Pq43jOrc5iBsWTVEEOtGFWzb9Sct1/IfS3zWPu8wG2zUNI8HY37K+kFQBdUthUQ
3YxDZpKoX/vP7z3hnYWS1/t5b3CxbYH4fCoomKq78Bc5zE0kctqYMV+iTvkgMGTvjkOeiGdcFkZX
9EgEM6L+EWOqI48Rvbh4LwmmXE2sbX86ilKuLy4saLCAc66APTT+5xzwwbvTFa0J76Ri9PyZJPWf
qaMAurPPsppgZxCGu8ihVl/bcx6q5Wr8gdfhY3y7/7KDUcpq3nIlBE4XEbD2l2Z6W9RnegLD+oom
cDeDWPilz34ZNfIciukGSmP8mtJezxW0x+giWZfZiuumjK8ZpaU9g/D9v40TyjZtYSohxLphnyuM
NlMuMxkJ++E7lPfuwAlP0rcKfsOTOTcXpH2guhUYR/dTKPIQh4myJjyo8gb7ByoJG8jTB2Hz9Tnk
w+GjCb3JnNBFvDePsJCRv3yemW2fqEuqVo1ACxld1on0tBQ2gO0Rw8+U+QxmD5RtZI+R6kApAyag
+olr8HZRVHrYkDACGiTBSJdx5Zw6H1mRc7UwZhSGVcUhlFhXYxWGsBR4wE8lVZd0n3Z9BRtoT6Kb
aHpudFCKWyy5X4JoU7prYGaekbzTWF3JXlaav/CT1OwJhDtbvOo017G7UZ3QJvz54IwVOTAaxYD+
fmRTT2AGgBU+GwDkPEJYjKoSYei7QnFIKlqeaGJuOrP8/1RSOvqCsXGt9KIZxi1dB3eiScm7k6cA
l62l0U3Lxkn7gl0vp9Ovk/kcFxvzcvdwL0CDoLl4LJHARCTMUc+IT0EpwMZ7F+NElik2gCMSQa2K
axZisaoma9L+SOidqyAFUNx3oF0WfIFYQCekwJ3Y8zjCAoVK5Q0j1OcrPFH+vjny99/5yYXRfHy6
dpbqGHrvmNgqF0qPUrEtdXdu9y/urUXwJVXqzhR3bLRFzLaMz0I9Od1lELzq66+ZFHu7Mv0wHf5z
FASpbiGykNEymxYNDzsjPBf4VxFH55csQcp14Q8m5xJgfWzcfrej4qS6w5+Oz0tSCgCpg6HzDYm2
QBEBIFnBQX7FmhyaaUZTmAJkxwHt8bWi8C8xLoKcWOWe9OCdB2dZ4spRWkw/bPg9zmPSLwHruDmZ
HG5azfw+9xWRn4pOPTwrUJWK395p+vD1woRTUw4RsGAlSwTEO/YzQGpSEXAJxnqf5P/knYh8T48a
467OMb/Ol+fF/bJFdFXiBkAbBUMZI1yeTr4lpQ4d8czympnbxBiaCriJP9ozVUm/+qjN6tcpgBIL
Jwop/JhFVjO2wYJwHBDSqY1H5zQTmK89MewB3P3K8IBsnOXaUcj2Fm2E41AuP5sDVSlWTgngAXER
wPHOj+4rMEaElCE8wr1ZizrzPW+wbOQ2rZtMQKT0yZDnkV1arzk60wpgdwjdgJVuqDsgsQfCjMxw
PMLUN2RCptS2mS0+IoorUNOyp3WjPkJFCZ2W4Tm7XFb0pt4WrUR2ypOSNzqTG7hJt4WcuHY8B1RA
b9TVUjVhim6Ws0MhSp2kyK0Dr+R17vG6k4PnM1DuXRWrtzeqbuBmlzFktHiqVCNSIl71m0KU/arg
cxQLHZvmsTlpHPUxT+jkW9QlUW4ZMYcG+8DxegochqTNk+Wy+y3+mfOYbUL9Rew14AfCc6fU0An8
7Q1EXhwDjzDT2BWa+yDFmjP2QGay49iSBb2V9VsMIsCwoRodU8P3exQJnGpGlHu7F5gZOhgb0+gS
4rCF0BrGM6vBAW3cqKSZH3pMNC9K4FpsK4pzd4nTdODBnhkZ/5ShS17kTeVyi0UES6KlPpPZCKBy
9Kvb56Dunb5ws/8mRbcnR+OXIXIQK6q/FawEIG6lpmlWDg55RUu1j4WAia5zyn6rb0sJ5S0MMKD7
MpSb4wbcV8y5XHpLPl910GA//nnZXeI0oLFC41v5/6RE3av6hz21XA1/Nm5v3hhed9PLU7nk4bPi
mGg0dyDjdF+nRvNVT+uw3uhxSbYkWyYaWrjL6c/iWdv8sQUCK5UGAFh4zffWBJYJX/iTHi7x1MYs
ZbU+uXy7ixNLvWgYTI1dr8qbjqzNbHWX4SyJNwDDecX17lgtiFnrZjvC0oRXY4I5W0RKURcxS7yn
nLjKjmpADdjBf9a+q2CIpIre9ZjzHqtarXLvixJtaU9//dvtVDIZ7q8CIUYsHHSzwESYaJNj5Fqn
LBnoz1oI0TAzaRCN8s3niWTlsen+GyyiSL6DPZiEw98CVUEb4Omy6v3SaOQYQ06O/heMkSt7NiSr
aLZLOKoT5HVh1Wfhvlph95DsRdjeMM/p7Im6eDQelK7cANPVg2989GG2KO72cCaVvKMWMrkJwvfe
u7luYSXj9FRuM3ObD2jFqLT/d0BRViE7//8sVFPP8O/l1AQHBK+lxvGb/x2qXWqiRM85OTJH2ks6
5HwKgt/dHsx1nPT9pyEbw7tuIvJUYD8472f1Z+6goO11k6DN2616bKilHqquHIvF9VIXrussYOnT
hA5hsTfq4Xjc0GEMgcJfzpYIve/OZQYdrAdRsgU1LL5sQDgEfZTwSN7yhbk18xbXSjREzg6bouAj
jJZG3IPA6cO7oZ/A/goQeDJuML6UKOjw3n6jdXOImP0K8ufyP+uweJBQPnVM2meyqfIl+sdCcpUY
YndoSkaj4i+1ucW2FQBRwtXctrFB7FBoiy71VrzlwHZGEqLHJGWxRvk/dt2vfv1gqzst3TjOO4hu
xPUZ3KtA+ZjT9If5BNn8wCgzWhTKAYAtbumPdPRGiTtg5fz5jgwJJFLChXh409JG5G1ne7iV8nDm
W0B6NQklb45i/zaQSvHKRO49LNUKxLXIACUrz7IgYmE4u1wCmYGLE/tfaWNVbG3WoUBkqbver72b
SdUflE6Pi354HC8jDfhwHCikdFXRJGcafVvva5otLX3uHLU0hwihNVDxSvkMw428Icm8fqiBOGjZ
dDsQFSt/86m8b9yXEb0Z0oLFb+1GSsmNA7XrocNHzxcrIfQgr/z+V9obQs16jkX0MeKKM0id5p2k
cW7byDxtEZsVRqe8C1unFaOLbAs9DVAY0H1i+TLZgYtZHkq1Jvfrep31I78DXmuF6xdcbXqDQt+E
NF0sTNn4qlgP5Io8tt9Y+BGE2Axa1TSJ0NyQRFPP9dt/Y1lzbC/+ySlIbOUMajAIGPZOrZyXIdo8
UCQPmWOLJThLuKZ3rjFdJiUI/Cg+2R/28skQjMqCh4FekEBQj4zJAxXQh9mGMqP/E/scQvUq5F/b
ObUzoiowMBUxFZ6Omp/+g9iCVTv2BNHQFKn2mzdmnz0x9wu+PGizki35vNU6IuzZKekZ0T3yuoxE
qMbXClXLzXLVCPObcMG6QD0jWmZNw1Vf4MwgG7xXfS3nGqp6APZrnBxkod1gvmhdgvg/PRt3HbVb
iHcpUzoopPpzzCqQJabsHmZHPGBtL5pr0S+HNibC2JU3iBiB+Zod/wKec7no2aFwVBKiV1XD83yl
812tud4bPKo8AXv8/Zv9DPCbxUcI+Me0SkbcQZHXScEU3FCSekIiII30MK7h8tPGXxcqWnLAeeAh
+gdgiV/t4WkPYnNLOgbZHznYRozPXYyd/VS8faGYaFr32YK4c65creJmT9lV00xqXa2pA4guzWt8
7jjblzn5MdemXpqghDhT95lHxQwB4F1CDq6ij4q6rSspe3qvuJ0yGFvxlwqIk1Kee5dGS6WN9oXs
21SDVQ/ygJK/65DEKzDxJUdteUTv1p6QEoSILBMLU+s/U5XsDuywcKVVuclavXgRgb7Ac0k8Fuy+
QyviXM/jxQMvHx1LyiVsrGQeYUJV11KfqK8mSzGO3rtYS3jiWoZBIIq0efOyxHjzUT33jlAaCsRD
+zLWD4EwaJvnH0cCPQ8y7TND+xf3n5BQbAsiwB08/1zOlyqDDE88vgWDVv+m6Ph8w1lyEBAfe7P1
brXW4Hp5BmHe7kSGgrt/tDN1NIvsgdGaGdbuQLJo9nhtJQhHVusO8mEVSntbpnz/AQ2OclyQpF1T
tHyO1PRI+4qfgQIxT2qMOwU77huQDXXCZyvv1Fgf5dsc0KqFTVA0AtaEekNOl5UA4jtHjBLZf5cM
P5qcQNBezPHS0vnb4Eo/NO//DmMW6zyb2VhytzpBKvdM9PnVrRTNm6if8FoN/ixhtYIakg9qRIgk
+J1tzvlnGaWaBCsbqgrHsysEOEP5L7O7C37R6SZhACPgKNoZlx/QhVFRDH2QsiCBWIkGnOZG3qqA
vixmi9YpqAwGnEolLKi6hcCVDb4ywOWNjgB0LlTo/i7EdR3kI7N99Aypof3ah0KKecD9WWXUs1bS
CJpgjll5uY1PHYrazyFw38Lwp0xVvyFzvxnoYD4LvJCbbCn6RoRSgxxsLEykx8tTKzhtWKAM6bYE
S5wXm21pr/zqtibeA2qxf4HH2JFw12lRm45no8OySMui1m3gqTe7+5MZIsPoHGod13ICu/ckl92o
N1kbwZauNDekFVmDETOkG4wPySxeNzKHWUeHIIvfjP0d+PTT5uEqnuMVFbVpHRcPQjnttRrtsA/U
kihx8FRnWqSRtf04/AwRtYc6S3NRK97kX1B9YfgpjMi7qqizOhpiyf+swreSW9zfxYNhp/k2gXd/
z4o6tPUBrzaiq586iZYntH6B0cHxOzpkpe7fJ8h7QtF75UreXqBY7IKK0NnDxhI+79DpcuxvQKht
1Lj8uyBpAgWNpnmKh/2gXgXg5I47AryDUZdvyChnaSUfesL6Xr6wcGL6tH0QAS7HaX6s0BeEh3eb
82lllJ2ORo6f8O3Wr8eoHB3QLwLGda2uXglIgkp/56J7AnMAk5fgBdq+YjtFKWGeHJEySTuXwnNQ
oV2k96kCWs9Y0zosEsFYoDQ7oL7go5VGEWJOi6hDSkotE+ILBh+4m54ko7FnUU2ZqDEAR3VECmQN
tCr1L8rGCaNEnVD3BNEH9e89dwI/PxcJaCDT7ZkUZW6obYpZDgLqwAopt2M0s0zRhuOoYPNXTo4j
wL6mUVMMQYRD6SDVx3iayjk6gQ3MFTW++Fbf9DGLUXzFqaOTRrLuSryZebPbdaivCGosOjmOTc6E
7HUaccd8Kca1STKDn8zAi642UMWs6ZGftBXzv5HlKbWKGDYD+9FiWql4NSQRDgrs1juE6vTCxXae
7CaVmq9JKND8aiPjw/WYidUfBRsZ9dCer3/ao9NbQ6eXac/A+lMO+NQ/bT8rtNUVVFyJ4a+NCCkM
eOfK6qrFgyMVi72kwEQncu+rw0VDufVpZoDoduhz6XDMNCVbRAcssuT1tr3R4KrApNyuU/DSBhRX
RIj4IReAcUfJo1Riigo/Vyz68KOim+ZVFbjwPoyFGbpJH5Kme6qztsM4lmBccBYDMrx5rHfB7t/b
KE8CPndZUE/IASaUY8Nu5HFYQ7u3B1Z0O2bm6qfyDV7BwIMAJNg37FOzSHLb8qXokquisErqwT++
RT8xQuEeEZIVcOJdG3QLxUczv5S3J1KQUYydnpuOaXiPQulXJPzq8LVCeJtk8/jWUj0d4Rj+8+P9
GYyVdrQo8Vx1ZEErkMmgNsvBG8yUq/JV2U527NEa+U6PEiQEaF5F1lmRYxuwdzf7BbCbWpyb5Lte
2SWWNVFmcqhYbNZJReqRfmXFYXUxJcN7YhN/RdjXHvqiUl7sWU2N9uvNUmU0bC3+MttkA7Tt6RsH
zAuuUxoUWthYaxMXuBsrPCFDiYxT+BGk0T404i9SWgh9SYhgwH3Bo4nSViB0tCSENv6N3THToX5B
L6IX4QXVYAbjYDpCidsielxxUSi8RHlg/FwqWQnCUnZh9jzG7TUQXl/nzLlMt5VWfXnDHZFEQBEZ
1aBbUUDZuCQ/kcOR84fxuEJAz9SjZYwpg05acUCy9ByGbSbXCEoJVWGjOjxsI9CPVZhlcRJbGhyg
slHZaPxzEOHyQSk6PwYuORioCRPpIDY8iH8qnLSlmQ/OEdqeMRTZuG3KiMLXBuot2nBD54dquXUc
ao36eelDVRyKiz2VCqEVWxnTNOK8YXhQtspaG+OQsbsBAzSbqPTXa0rTtcSz6xxwgGiGIMqu4/Wc
HyyAXyTf99RJn3AYMsrQxoU3ncFpb7F2gDJg8uEvKTPnn1vRlxTXHMMi/qr3x+pu4eyMfiLMmTL0
agfq+SWXBloNJmncRQclIxnUARiFWGmYWSN1j1aNxx2Jy6n7gwV9Ei6xIQvFXFMxkitOV4Dzvq8l
V5S90JlnJdQ/3l6wzgOcHdyqJN/V9bp1brZXHI/srXuR4/sLAgKMZiy9yt7xLHJR39rSJCiNZr+z
Hm1ImTeBUDiQg5xT+a4vBSKpDfRD+bAKadrUUC14vKmDkKW6J5VdP/2erRxXMfcsRL3uEGJyMoBl
fyEu559Le8OFukQ9or+bOh/VVfMI+WkaUoxlpq/iUETNeoKcEGeuLs3WbBxRWh1mKeRJuNrpf6cX
dF7PS7X/inCCmTZsMTC3jYvw+X+pufzYAmKa3PzTQrARVXdeH2YkUTzyX0y6tFIM934H2oqLvSyr
qOJuzHUua3Xs8sDcTYAKNf9tbrHLsZvWqOtM/CMpKxZXLRjgZmd3pvM/3eEB0mHPdeSzboMa+fmK
sFDNEqiHg1PXUW4GnbNNqXs4uDBHPhxXnLaIp3XENJsTODXoMzvjKWnZlaJDuk3tLkZEoM7cJUHv
L8IMDPOiXQMr2l0euupbzyZ7P9PgBnHuf3Tg8tuAWMBulFHfeOht9D7bvxvgtnFPvWHe4iFk8bFb
7ePeJbdHa0v4tz+UNv6tHRq1iprFaZuq9Lq3yGPuJyMnSB9Q2hL8fE6HbZyw1+z1Rh43NafgxxNs
HLs+RGdNMB7dKXvN1goTii+qhcSKd6dcaTUDvrqVp1CvQ07m7WcgSiyFWIwoJSKEWdZdLIO5mR5D
D37OcnRlO+TZR1481JZnCEFhiT93umEn01mbS9IW7fl0Am5dfTXqx03qH+MsTqRatEuPLId6/P1q
NB9haiBhnDz/2YfBb7/Md2TScndnN9huYl3U7+moTnfwBwlT47/gxHpHrEyf+5nkCBEfLeHNpTfy
c0fm8XCWhnO7M6mSlSnTK3Ji47VknI7YocfttLCli/gXMAQnpvgtMgoI75IFQWypygGJ8+GwOjKA
Dw9elLm2OIemOcUSkFA5dHPPBuKJKx9oMN+SUd1lCf64qM9Pj/xmpFJwFi929VHGv5uyA3NUS/Yi
RjlMaURhE+PiTrJ27n092StsQMiK1KzfFFAq7L4lar5lxbEjG4D4F1V5ucClQS6GxFCnU+wLDmX3
K7TYBo2VZa8tE7bgc24UFNvBkMQrdRWctwCv3iqjZedvnM/6JWZE0BGuqapZXZxGj8P3Ud5oijhk
GgvQwXC8KmRQe+pMVtN2TvhJ0cxiIvlxo40ltvG5hg1qDKDFHEbn53S36kaklyin0OW55PC1LFW1
u70jBvQNEoGjpZB8xKNDMjD+bs9A3OUvvaMoPhcVW51AM5zmJwXv67t7JcAGG0CAHW0QlpeA8dGL
ARjUWk73zXUKTgOj2s3CguNFw6CCnHRNOXXnCMdIsZq7aA0PcxQf2QpTC6Z88lMwicLa+oWob6FR
F9LSNqiiHMnZ2Slmm35EeP3ahgzfixL32xW7A37eJmABjzVWJ1iFfeggDkU6o7wkhf/A8rVrLOBH
DS8C9NL9aqHM3s+W6STFkFeqJ4dy6thFwUH8KQVYoUogcBlsl4ZyLurlFoC+ReTVk05rxq5aogMn
71KO2RP2LSKRlF1wWqPb5bLjSCsaXtPqF7qKWOYJrDEZkorEL2WRR0x2A/P6O4SKCBOuU+Dmo/3v
kKq9ZqZp1bSdMdpKf+LRykcDheJlib8sgkOL8arMFQNtZ5zuso8AC998HmdhsUzgMSMLqKt4i5GU
YSoZfTg69uIXbV7uvShvCDiiGFlpDu6rGlR9ZfksPsUwVGb/fENfU8RELqKyvIzQWBFBKPTX5bJF
xP/rEyEZE+3XyurPoTmeGJI5QKFus8To0Fnx93Dr/rj4o00+DN4kAoDXryHe4CsPZrzhbqhKaBUu
yXqRymfo4ETJp1ttk9rWJporI7resA4SwlkARxlWJryGLHg9Riq6Oj0ZOr0dy9LXTf+qoX+i6nuD
+t6aLNKiQXFmXge1IFuQF9FPjy/nza36r2AHuvvVBBj0hPuQLcUCNYVJWQJeogp2k8HI7o2oeS/8
zcKvkPRaazzgqoE/POU5+Y8RDipWpn1S/YVgzT4phzN1w9+1kaEt0laQrZngTJtZot34XyiTbOwE
CKUK+41LCA54iOjZSVVhbS/IVXylTjfMOlFvpb/AaiB6VHwLpTxKDrg+X++3niS59Tm+oLax1s+t
1gQ5n3sdM90jXLYvy9lejuxnQR5n8/xoq136zlLQsEx6ukQYSvAjzLoMspjgB1gbBJfi4EgqKAe7
oRkJvqfgIMk/+D2G8ZhI2CwZP3fU3RSbvIvofWqZ+GELEVP2YG/RxVd7POggQTJi7pOYRTHtxWfa
GjucxZvqJcHdE1HcM8b6MOauttIMMMFOyb755mkuqRSUPFUdGnBrlUQhmGGEEml2YEfckWY0R/OE
rXAORB9Xwuz3+5tDFCGBTGaADN/ar64PJK4gZ2CvPERa0j4RhmVempiXl6beb7rN/ntjH/Qn4H0Z
L9Ouu6kdmED7RpqnnDky6Ar/zAV/hOBnxS7WblcI+mEJHMdmG8y72lGPBzmBfhMrI9hr4TKR8y6C
rdlvi4npGbal74RW18Sl2xAdmKqcPuA3ZTxDVlWezW2mkKwmqQ7POSOEMrlk/DDTwxWztXa6lyGj
Y5b5GEkblBLrwrHgNig0NLOdNfGwx1v1fLTs+tSlZvnShKAtekpPUw7OsYiZUF36QfgP6YTXCaUK
kPTGscIlWMkwMgtiehfTxeRUxscvUOsRcjlgRJUDKH4B9meCeCqkV2ZHJZVkLjQ1TeD07TOKfR+A
E8Q6wRg4BVGmlqVAvuY++GGSs9LV0a4YOEkHeLMlPJINKnX5SASwl/94LK7ydNoLSM0lN25uK3cU
BsPbyZF+NLYvONWukAhjrapGRKERnm4swh9tf62xP0GCxvV/hE6iHCIByHMweyz/fBEbI+Kffk3w
bTPNiDfKp7vS2Skvq0Xwsn7z9HfYkSScU2rjWb0HsNyA+OFAoi0SJIcsmYDTKw2muVUe26guJXl3
8wukvBbV5fSb5YcDACOH1DZ8rE5GKBVagzgduUQ1hWiIok9h/FNKx6e5lptQ4ci6uFaBCYOqM1+k
VGXpO3LWlrOn/mvCxHpjUADzDoJm5xe3ZX+9d5g18sboqZYI3+Y89vvXDhMqBHEyEVUUXxagtxhC
K/8YhHlWCiA/Rkcg5J3vpme8jGGEfcvDmHY7dfSuyEAJM/8zMJUrUpPCqkgwncltyJjQTsPrikE/
PqMZzugDUyDpVe1jEletWQvTzCvha3hcfRQvoicDEDVuWPGoMjYafzSIga/caHZpDh2gbbdl7mjW
QUkyMozYXZcqYGetciXm2mUR7B9E4ZgvrEXNdNZZtkHVxy3FobswcMflprBBylL/zWCE9+JrqoZS
AmsOCEJKdRtPozc9kAxAeiaRoGDtmdzPO3NJJm2iyFmLytHHOs062uWI65MrFHywT4EIaP+S8nMJ
GZSrdR6QGpJfIQc53hghLuK0wE5AKEZEINGD6Luiy9uL/DmpAeXzzwjXzKCjPHZlSJGn9R/HQb4T
blmfGrjkBQgKvDbrTfRuTLVjf2/gVtXwdnT9a+22q5G4tR6fOW78DdOolTFviO1PgDRuCGb3+waU
qYnFpuVsMbeuSf9S/BkhpTAZREMnr1oyZKWA/J1FL5XDebU1qa63t6OGBAKkGqnWyNzOpWik5OFM
WVUZghVW9EZu6XmJNv0Pq82nV9HF1TrUvVrsh8O/VKyOnPBFncEPVARvGP1Peo5K6mtTQwn0V9Jg
mqB3dzAkWVXu/ltYTot7bBd6Zb9hVBIZJZCe12s/FFLABVybGo1d4dilOJpw6eUkklONuw7ICLed
jheDvvDVGWR0MIWKsA6q3Y3VPwIaGad+SmjBRXdI1Bwe11cgxbhee2xcEGEpjrF/e5XaQrf1c3aY
mZqveVOSFNzYRQ06vXnT+tsScLpLWTsIEhJwzLK6c0cz8aOrOy90oCeksksWw2IuNjVh3CaW/C2A
leLYUnb8Ga/Ehdl6o+FHfUkr1JV9/ieVPLgyjRn7+0X9ZM7B2bzhAY+HUb8lstISl2ZzkzpE6GbD
j4r/Ey6Bl2DtwDXaT2oOD1A3MOCcIxspNK+903pGEFNVa6G/m+W1HFdaSC2xHzM5T0xUxPclzvUA
6HKKKehPAJU7Y2MEV1zezzqr/16hMVmFmKPwg9h5qWaEcICYU0TkLcbNcer8X9W42ddCfhKsv552
LLMalzpcRD0dY3Ya7Ab194K96/ypt2Wips2Ph5ROcg926A3FKsMIuW6G1/8eIuHIfIqunsqypFgy
6sLeRJEK6lDvZaVboh+LCzhLRTXcYIMTYPFMv3AK8JVULowDBhIRpj4z0l6BVFgG+6gVRWmkB7wF
zGfln6ecJ5jXmFFuibE0SSGbjpGxCBBhPRacdKqr2qBhKO2SsbruSraRpXNoT/kVp0UnAXcCp0mI
XiwUXzQIYPCdEz9izttuxn1TOSlAEMEV1VIetG8iBiYEN0XgT0JgkNjaztUeCgBJPIFv/SH3HO24
fTwOTpDljMMs2CjTk2VxJlMw028Kz9RboB3IUMHNdzJTVGwguuUS8Edmn0p0moCH3cH16ZtHa+ZT
D2AfoaVczH8JOPFR6y/w/gjnsdBySFwKE5fPDfWGIn7K3HlpaBO/LyBD/O/8CjT+WovEwK/dYSbt
j+cOKXm5+Uek+741em93nhi5iw6CywKZRLaQ+2bCRfrNYio73PAKGBnGHQC4e7QnXz6Hh6vTfV7S
HQwThfqo6tHXjlbGToGHWwGR2uMF9aYwrj0WpREMPWfyOwa0GslcK3TfBl+rqBOScO/nEum3HnLG
GfvqiQXVcADHKsOg/fzbPyVquySkUHT8rW4FLgIkHo+kFLqnBgDN8YsdhSkbIoSkx7JIQfQSerhD
Woo+fONgBV8QalSi/vRmXuAD7UR0pY4jQ3GpW7Gcam8ZQcbwMKP2VLALk65MWFIs9CsGs8ib1h8y
RqB07KlyGLVO9BAgRszIAPScl/AYtK4EwYneBXn9Y+VGU65eK35916inGXZ1rnJSytZeDmJzVn0Y
gdNDxDfX4bVjNufuTRzq4mepUN8sZG7XGvigXyTlJNsielHbnw7vKSoLX7BS+OGjW5zJHlOZirba
EUy30bkWohYfyGnlroEkXj780TvQnNf4ZcPJhytrLG602z6LILBpX78VfX+RXATsVhGdGszJMo8z
ac42BTGB7Egsq7UhgosCq5rxe759wwwk0FZnipuaT4Qy4fpwUNkYRhMW8MSi8PzBwhdU1MlKSky/
ztjrIlZv23xxMADfoZlV6STR8pz50Gi8xgA+5aZ8jG5djWztJNI65TL+coubLhhrOZKgcZvpoNn3
WQbtOyfDd6SxpvC1U5Sq3t2NQDtVlC8paW4ZQOANmW6YRiLi6AmE9Lo7gHDtESyZ0hF2iHdhUZkK
RrgeDvTkD6g+7iLTJ9rK3WEsYvKScTAXg9xnzbLgUtkHnv7XXW2R9AkmlJBX60YFVN5yB+ks/CQe
8JamZi/gWn6fQYHCdbCnTklZ2RLUr0E8xlB8AqhLsssKE6ULkQFnNMy+WUNK6pVHq+ujRZP7ahWH
LpJYDbvKKIYL8/Kj/A2tReyTORSvo1pk+ab5UmqNj849s1SKaSzNuzW2TusSu6lcSg927A6pzZBA
Pv8IDwrn7OhGY73kxESf4QKLPt+iaXaXH62E3YNCO9Ody5C01g1sDEgtpIDVaRwNdHUAwhG6ywux
3kmLihQSotKEcNhGoLiithMWtl77UOKbcLy4dPfqix2DuE+9Xo4fpQqdNRDnHiHKvX2DWJ6NQut6
/UgWQKJnvdoxv+I3flyHX+jYyozwp6CHcnFgbQ6F5xIOUD3tdRD8pcBfud+KEOS33xkKk/Q2quOg
Mwra3uwr4AFknJ77wLaGo6SH+G6sC6qg+V3v/bfrqIgYvUcn6tYUiSNUwAU5+5TcCVIlAstG1G+d
tTSVz7FJTR3cgNQOQQ7u/0oJq/aCbh3+N1bwyCscf5InkxyVf9Vn7GjSegdv0YWsTHFlXha8unC1
BK8RxTzB3yxlWaw/bK0J87LmkmhKRXwdqW3qoFGjU3PeMJXdNp+ABGkdw6sL7BE0wauYww8bvqbd
73KCKb5vilzkQyXN3kffPcl/5HNtVyTLgXopRn6w9ZlNYVXVpo6uJYq8gjUoPOoaFVRV1WHrmppD
icWHSN9ePcgeWHaZ/JYi9OscWC9WEmEZapog2o7ZbIB02Ysy/IKqDYRPabKDrzl4/VzQDypCutPc
oF3ZWZolQiWoz27bRYd3Fktr5fUVQ1DSsbiI9OXUTdjCOZHyHC14mavjHB9z8dNaFgmWGmy8Tv3h
NSbhJ22JP/QhLv7L7HAhpzFjcwbFsKYhelgy/mdDIg35adID96seXosH+GjuTFlqQy8Rl/aXc+YZ
4rxl1OFrs/IjW2nMuucf4Jo36ROAbAz0YWSxJn8Ic2/hIeI0dZZTbYlS76co0TKqji5MEKUyvEjh
Qk/9oqFQHTEOJ11+D8dsSFtJg3Os+CyJQdT8+v0iU6Vy/YzH9s359dOD8Znbnw80UcGBOaQkuhNh
icjOc15bMNKSvi15+4vLD1lpP6RtoVJw5k5Acv5MXWQ8ONJTmdp6v89eTzH5p4/GxVpJuh2IBzI0
OgStjNnL9iHmQYY6X/OdB8JSwZD35g33LSOMjxr/UdZuVSCzIlyZEyWP5O2agIbCAeee+oa6BaDr
0KZ0Ud6rOfNyNIVejVDLc/QCHGMfNTC/h3U4ZVehX95M8q2r6IpvgesmHv6rxzWiEuSu2Etl+3mm
YNEiscFSimafLhqEbM4J6H0UfqxapoGVo8n0re7+0HbH7STDUB7y87NcN1sP09prq0+lHdI7dewi
Mgyk/AZYNlyWBvXsTH53KKiYZ+tIAu36bUYiWX4lsLoFcnmHC8koh0+ylLr8Ht/dmpZgAT/YPoKL
YiwpcapJpkUAyvALGxwyUDLfafj2F6E+erJfPwOlYFl1ueaKIucKzxR1zHERY/q0+k2YDmXoAUCr
ZsMTasMQK6W8RgzQdp3ThPdtkw0QViZJVm4gBuZGqbOnoaqC065ro4SwzUaR2wAS7tNDnmnaYuM4
WlFRn/8HOlFgIkyVdMuxIxvVNTMmDAsu78PgvnMb1p6pRDDTCQYca0f7uSPPqHwONlNjN6cQcQGI
aQUKa4WPETs56w9RRYYZV235A5Q+I7tvypcIN9uXgoDT9TeOUnY1G6GqMIT8H2loXVIfjdmch/aw
m2zBD4WA/8Uu5/ODT1bPUHWh38IqlLxq3ShqR2suYLiZvQGfqXvEQnZh9MJpJ6KNM6277brvX/gl
u7E36ap8/FwOSp7MOFGVbyG6nc0mkpnuXMv7GXYIiF8Rim6sN+A8ItBmka7IowRb4HEC+XstRXdh
3HaUMglDmXErGCVsunnpYk4OsY2d8ObzKO1jm2RAlAQKw3H6PAJP8IF7xg1QCFQ90UnUMp6vm4aI
0zJi05PbOPiFDnSDtcp5keuTkqKbL2eIHGoS3NVzmxjzpTE6u9DeIAcBD/+4YK9E9yoE0nEWEuri
zJzLnyfTt+dHhqQrQl91bI+VXZlxlLD8cBU1x1PWR8TAytjjOPtG6Ibu/HePedBk7wbs7qw1xBdZ
HHxTNpjPa6aYPUszyJQ/rs07l46eGA2NHwgupXt8hnGvAn8E5EUImCi0vv/Qe1kz2IAsje+DprU/
+32GbECNZJNo/NmwyMtNzcuDkYRhWrQ3joCZD+gh7EZoRNEXK3Vp+TJNUvqzgWUr9ULSR+jy5e+1
/yY9XZejTVFxKpf5rUmuKGgG5sjtEauYbouyifr8RWZEWMQCJ3vL4/PL2o4PfpX78NKhxfgozFpv
xvqzUklfuBt+VKeRV4ax5cRenyrA3titzkDfgXeBVAD27cmLW/55stfibf4/gknT9Eu07lnps2jg
Nohbz+3vxE7p7o0JOxhMlago5foOHEHtIm85eZrOTtj2ahRL2ZpqKDZ2p07otBCDPNDXGI0Eehvu
XdYI9MuMxktydURkXTGfc3XeyOXiLPJub2sEsoIfEG8mznA+EYgD0WhdxmeD+EBRvDKxAQxopyUJ
/nv2SGIgl02gIGbuRjVMui5wW2uPFgWNyukhAJNRSQDdHm4W8UF2iVC9nmKWH8ICVoOlFM2FuNhe
mRDbnJ42WZJGZHDTBAnHuaqF8bEMrHYVJCPdG6Yx6xM0Ms+nBpHVDyIflXc2sUZrXlm5PZyzmK8r
f5H7QMm8xgu1FA3YqrAnCfBKaMP6sQ0QL2J2voMGD5/F169xi7ex05EbNSCGXN+C79fGKcxACnnD
V9rufkGpdAQi3OwmZAtvbiOQeiJOImPm40l1dLSreNXqVvWSqgUp1e7A1vcgbIrmfzyGaMGFCVG8
O8Fuq1evWcvc+HwsGe9TRth3wULEJwG9SZKEtDoifpIJaFcIyqufTbpuoH7czjDJqiksEWYegiJg
Iv0dZUEHp7No3bWsnjt6QNiFDp6zqme3WlBeyLn4U9gQDbKuZswhDxf7N6pUXYpPLiH95ooZkX7h
luY2lAH7n9UY7UkeGzbZk2dcLll0OmJXllSrI+HiknWiO3lNcRm+aXDrGjpOJ9EEUBMPxv0XMD9o
HVi0otwb5ZM1ef5Hhvke77Rx8Sh5NBwkU+rNPUg4C6h6g8S8WSoKbgqY5BulWXjop+EiddJexJtN
L1r9HA3GOgD0p5TCyZ/aHaejyDxCivniWeZ9Tb4wCpBDGhl4/h2Ty0LsfODVpoJjH2PpfX9dms7J
PZn58HgJrA6dRWGYC4wDXl3REo3+zigN2svrNGsj7kuYeMQxDcgB8gz09b4GyIV1VxAC1m/ZkFbp
JW8U00ExYvCefm0vIMqTuouSzEHdT5DP3Hpx+lrAAJMR6SXuqy/IzIOD6D8ZIebJ2ctDAr5nJK0s
fkI0scF2jWObEpmGsPHtlDatUaXTLWji7u01FsJUfW7QMi/TDYIt8kbe9w+Ogqo5qGb3BT2rU1Z8
Gtf8xxKdI/oFYIVA13AMbkHFMgVnsLA4Uf4LIJZ8dknIrdQ+EmRNsnxASBcCumAJRtktsA7b5Qz3
vu9l5JW2HHg8lqkQ9vlFwehl5Le9AnOtt6g/yu7zq8naqDdcUMlw/lGARRmuds7uuHaQwdEXlnLo
zTvaAzxy4o4bxigOVkhS/MVO/WqHnNVM434S5aKHpbaV15TXmx9Y7PBBdGADVNMt1/S7g0HKoTcr
FRuSaHgJBhB8ZBPoCY/mujb81/lnlg2cH4x08ISLiQSyeLJaghj1zJqzgUJ+JmbD43Kq1qiL0fcB
0lNMTOu3FVgnW/QAOoZuKiATYtiS6R8a3oc/Wme3lmlF/P8NDi7r47fTDIsJnfAs4ypf3sZpg950
Gcwcv0vZ9tEcKo/etSL4rLdZS3tXhCq+adAQo/UACGxoezhTBpfC73/JtmoHfwVdIsumdES4xwVO
bsOla3DgifAuCnvRhXTJwesq6jox3LeMprT2cvLZwRoOMaoRfaiCpX9BAOwGgmiEXMznrcD+3aTM
DC63UwLF6o133361NGCnKKBvaVbMaAwTH5NTb9fDBixK7/oRtrpkv8Zwf32fcRdXB4Z6jVfkQEST
KkV1JeDNidR+3Gq0jhJeRG6ROVs5wUB/gDJ4o1lATAE89IRwH/7AtbjtwEVfgUZz0J3bUxqUXaoh
Lk7ENCdYup+NCwA2lfYDELSOT5nRvOUTEGih04iREkZNID9YzwNcmi9eN1jjKl7OH5FOuB+0IJIH
nZCjb1KgUu9MT+WcxHRYqImfXZ/BOdA4KO0+9prqH0Jh6C/PLvp1s1u2c/EX0BnRm/QcNlUGBbLA
Sh6+BDr6wLhtV1+v0TKy0HLLfA3Bi/vqKnDKaELNDupAYv6f2HMRkNo11gMZwt4UIH5GrCngGi7J
XlaKuZ8sYM31HDdR9reywJXBsEd8tKOymNLypUWjnXQy2vk7PRJKysblS3tjWYhPH07hOY7W1A6I
3JrOusmTHuGbwHN/ks1qZFKWyMWYDCwp0zMBMQTFw+g2Z2Lg7ZocsdRpQWS4ypVtn98ajlnbBSiD
gRpwibQ7XYFktH3YrP9Q20KnX3JxIZHyelUplbX9JDbHr6aXlE64Sm8+EaCYa45TAJWK8j6tBwXj
wZgbN53BJecNIFbxz9xS+CpA2EQo8p2vTnZSUXzcz8qK+DqhKlHcr0Z4MyYbswHF9g8vaXHhK038
wTrGA4uOPo7N+tG8DZoreclX8xndHPfxH2Vfocgj/BC7zzn87JspLjX7cZUS9JkeR+wY91kxeDvr
e70qjS+HIuHLcNyYYLS6JF9/JE+9QaXvSl7fpu2AUwukPdNCIxqLz8BwcLKEVw4YTv2kQmp02zKx
JKrSCyA4DgZYN44uC00gWVSOnyBqP/KpZ0D3FlWhzvL+LQXtpRI5Q1cNwhDzHZmbLm/5YEpaso51
corsi7umq4RUGZYR2YNW8WQsONYtejIXm12cINLOvXsMxX4mJTEgKlrEpR2aHuU9UrxLZ0k9VOWa
0kU0bk5JWI77I/fUgA7g5kjMyBT6Zijm6Oz3WIk/lMXEI5LNX7GZjja15cOAhcT66ZtEwrJv30nB
t1exFDuLCyp6Ss0EkyU9BGJXu4D6N0aTea2LSBOveRaJwtyoaCG0tGOLpuWDg7/hgpi4559gE/74
HmEI/nRnpjuhnFjNrW3YpQbl9zH+UpGygA5cSQfFFHCqFM2790NkJkO7Slxp0ymz8gTL3pH+VpZC
ONj/trIT27ZK/GTy1ineBUgwNDBKgZnTLkh/GOpOoBzJmBlefWyTMAJbwEeU7oAcb71dXJ+S6d7n
FTCTLM0wyofQyPkxiQGglSThnyibr91tP/e9gPyLRaR2VVOpz6lD5rWxnWiG8IjeVBM/jLSJGbOl
4ygAp3KtCeBykvCpRZehvux09KJMkxtrVrvO+6yfgRGGQrlgTb25aLLfbMnJCgmAdD/1HI9tkcT9
J6y6Xqf7iseLJlLaqHTYkqT3ec2ri/S7ZxtABVepXmcF1CzzC36x3SSYCmKznD6u1NSQ9zRg8ysU
yFpoMfyOz8H8MsgEH+cb4PGztUAvGhMOJzdio/rFNnMiQVX1biLCejakaDnt8FCd8p5Zsr9Rophf
v4MUliEz6oMBdThonCGbykrZEOczAVqH2z9e2G9CzCHTu+ncuM1L8jILicar1K1OcS7t3DflmbdN
zbamuHnnyw60d73A287nLaYWYtzJvYhkxoYMiOVjPVMlPthCMIxeKFSClH8pInqCu94RN5wn16ux
RXgPnaW1FPpsn3K6jTS0QWJLjOvxjBopFJ8v18MBUTYIMuRxZJ4wiy1tLm+P56mtQhOEB3v45Z/A
gvFW4Q6/IGJe8VerOhB6rSpzS3YWGDmuPGpOR8DLUY/PbXEIp9rG2KPblJN9A3DEmK5B4xI5pijm
EOu8BE2ZG8WUs+AlYBec2m8EhOMr86agfLS5XH74hThLax012Bgesx/+pJFvK4coGps86+gXW11J
8w9A+aTnykWf1gl8EmNKX+wLuvJh1diKTXbcWIKM4t5o5Vr547BqQADGraXo2rnithf1kEuruzB8
E7lWQZcWhdgKTQmDAvbsI0z8MxTAgpuX4yg8dzjV0mGrwrp6W95i3nYOjyAhkMoEV93t1Hqv/MsC
Oo1eiMtlsBkeoBt09VeMPey+STkS5WcVt7WsPNfJ4eXy+k9FbVSG3BAEpkgmgrq013OEVVMqT9ok
65VO2l3M0cutmJIHYK7CW229pErdEHDvrzxODi4meqL8nVmuu2C6c+8a9tJtGzZHJwXbdcKq/s9P
xJwRA4TPU9PqEnqc8D8weMwELzT7MRvbQ/BTcHsUcDkAZRQMcqe9Bg86x/8h8ZMv9VY4yLBzSG95
Fg0s+S3HEWAWpfZTRNy2H77HCR9FOsZpl4Nk8WcldO6mLIOUfLlbv3W3015FY3AiL/S5Fj7u5sRQ
bOz0A6kp0Mkd7l17lsn7eTMXGmDKfkhs4KHl1sseOYY/vWLGKGY5QoUNULQL2usJvVuNgDBkVYrK
coGYRvsLtQagrOsh8BNJBTmP+r+IDMcz5UK3MD//VQyWnPFsmUdYY97T/hleVrjes5Q2paQ4svM8
T2bObUsTrmitlgvsksDZcU47oXvu/BbPxzWI/OFisw6NbKYNrUU0ev8enn84a+wC0RdNfnmdYEV7
27JJSzxBFYzggbDDCeBj9SgyPKGyIgqFepAk+Q1ujykMhjZmIOOlQSg0WttEvGptx1GYIq429vpF
1JB5LUYqhCrPriQpIK9u9kGOQZApUTcuKPQcFFJZ8lrWRp7Dz5SsNuJ2n5uzHIx4T3qkVfLB6VQU
tK4c2uxtmQG30F6dFklTb8jJeTK7MD73TCLfIlkk39Ajt8bzgTxeubUOIja5CmHvMdWqraADHjDQ
7O26+UZti9gzrxKlPNFLJtjo5cHN6zqYR/j/oRwe0xc/NMHNfLQchIw+ska3Ywjol9JWNXgj4s52
FbzFQS733+hq/eVJlFcmIl4yF1/S9qDdJvRWlyRQaTKK8XjygSeCW7O5eLOcCxlRizwPyOIN82nr
hS0dRWYJry165P5K/N7rjOkdqgRy73uaHZjuLgZ4isqMVc4sL9mTMFlE06O6sxc/cAKHm21AhQho
AnxdbXWcFJSMkKo/PecAi8gf/VoQjnTC6MzYTNhOwX47YN4lwxujdLS+OScRjFVZdVGUNWE19Yyt
WqeODlOA6DLp/k5Edio7A7eVheHXS5ac7LQjc1APCpf6GM+5yrw4yPesHsiX8bFCuJN1jVVPrZbX
xV24ltfK3hGegfsd69CF49ajew6gTiYEFkII5xOT5nKKGFF498EA8L8vS1HD0pDrjJeQ759+rubH
ov8rmJ7mIZGVMQ1b+SWz68lCpc5XXfXywKEg2tqrd/0vogVlX5llc4SeKguDACv+hiZ0H79Vq3MN
A7MhupTizx490nSFynmTD1A1Li42hkeMyO/VbDz3MwQ4h1MnW5VkC1qyD+zdsDd1AIFi2MaBWvnY
3E4td8gVMBoD26A6cO0bnFhgmAsCgE3EwYX8dBrGkgIgtB/wqWggZ7u91OiSL5vW/WWSeV1UfwAd
QAouujjQoBRl1LlVkVq0lsBTb/fj0aV3RzrI+rH9kqGAglCSyz/ltYwCO+JAjUArKQtKfOSkfUyb
rruY5xcQbyfbmV3MmApQz194zzJub94tEiFsbXy4ZJ0YxaNxH9PQubDB8nykuVuUIXqf/DV/yCu8
IQm+JiXQtkd95EucNCE2D/OE0DgmVkfkL4zoAUQo/lHooGJns8VbHd4yDy6y/WdkhkSYcT7/Ue8h
maVEmS5djlqQlHrriuhfG54vtm5XwgRRYOHXfZJ57Hh7n6lPkVrRVrkvYNbPNnYwzWg1Ee0zMP4Q
YBHkjVwHuie+mKtIJHoydE6GdqOEafg0wldnDh57gX+IVcM7J9E8CbjTR2a38D3usOeqk7wj7kNl
/Zu1wibDfQRs84l/kaB/ehUUFr1g2reDwfYRDKvlYpzmGfomU5KYLerGPuurvj1avEH99buNNrmm
LiVW9LbG5KQM7bc+YP3VB4gcNXHLVr7lJbW0raW0dokcsWqKzY2DiUNEr6Wm/B41eA8FFrNMth4G
IXG629rgaYa81RpWo9FyKwIP40Cq+IZG1mHYTTL2kgwrgtwrXHvnSAJKRNi0t0/frZ4fXiBPzoMd
pqb7u+6De8iKiTEw9MnbBR704Mo5kMoas9E+89L84CYqImOGXxlTYODOAK3wy84fWMgdIxXXIncy
J6mkq60NgrwJOZsyIsikERoL65jHyr7yVwvmr4JPWob3iZ82QnUsQGAVCuXeXxsTzLQjyrntN83N
BX2NQhH4XWEyKEJB3tdrsWT03l7wl1TkCJ5/ObQZILClPSalvF8B5H7lGZwMg6JtidMUzkFXuiy+
IYcWqGKBajB3gz76mD/t4aLMBNFNiQ2zEUTCoKeoQQ4YcxU9kW8Qs4aMScZzVnLK3tIboIcsWrmy
ej1CSeF6QBTQLuigsALL/ZYDVnem2w5hhISz11d6oOw09dvWBaR29hYh5r9RTtszgftOyy5AWQlC
Lt0CssqBsX7GmhtOEDxq2TO9+ZLoimVT3QVuEIQksp0r5rzhTAqzTNw0uqXX48XzWI0nD+YU2kcn
SXKvAnEZXHODC5rQnML3lB+IzI6IvMs6xIi6C/MRaN/cqcDIu1/0qNQWPNy5El3c20Ah0a/u4WQI
NiFF5CPn6t72Uxru7xSf3ZqDsgaYYskogHXuGHg5GArPBNz8QSGOrIIkrY0leO2FapnOaUYpVmTp
Svy9T/fiBXSHWiWyl27RV0bMxQmTkBV3+F187spnbc8m/ZGu/9KB12XVniHepImAvjVrCFsu43bn
0IQpCZKIMaIQnzEfZ7xml27GhOkEFrfUXuo99v42pespB5pVMV1cr2VbOQTMquoY7WSss1oLrOXz
6oG3ydINxenqmmFVozTOi1lkK6pbbsg4m6LXdCbJmKrYd5LafuBz7WwirLU4F31vNOjTxgFK55d5
JGJ12DmTTVpsP8f1M5nSigXZ86EcRaeXasyL4dOU12Jw30MiiNQeFNHhetxz3DHwWBRbXgbc7UEn
7/BJBjWKH9/L0eMVRq6ZcggAVfxytlsqk2kkyaopVqw+VeDFFxvAUydJVbbAh7p1tWfxBbodITtq
t+G+NebNdUYyGen2x0lfaZeFfzKixc2QjgLOV/wha3SPcW3DpmpgGSMUNTqHsrHbw4Aq2V2Mpn4H
1GFCaC09P+6UNLflhg8gFLKFQypHmDOJ0UeynrKYkagZZc9e8X6IaQruJdXfhfZcX8kVTeTNgFjZ
DCKU3Bkv8l61V25i8Zr5YpjzfeRaDwHIs5naEK19PFLybF2p+Dcn1S45AR/F7IF92Fu/B9C04giB
39KDMF65mSENbDALq7iooqaDsG6sG8XBXhuYu28hwYcvLQQOph4KtMvAN6cW/IGne3Ipz4kp41ic
silRfE0E1oguSIdTCLBqO24MO+DmNbABJ1fR9cTPJ89AoEpftjEJGuBOUqrxtOzQjjdDa5a2Pc6v
7Raw7IMzPCBnVEVGy2Gv4eZwLGigvPcMLFdFizapL39BVvrCTDelkbjBPM1eppdfr4i8vQjzAxGN
xxtG5ZOyVF5llpNXDuSFx9KEv48nFAj+cfBXzZc233aaHqh1LjTAexyKDm7DY6MQxUFQ3Gzyhtnm
vVCk3/YltK4xpMjC0BYw3a587Y+ona58mM9LuVjrrQJ6YRc5Z36NeI2XQIWxQEFJhc2sD/isP0U1
Q09D+NCSxyy+0sXr0h8V4mD4P/2KVlECSht7BAISSt1GsjIZ0yJXE8iXAzzclZFdmiDvGkectAX4
Lb+V9CKCtv4pv2QIKdX7MdHh/rlfyMvxwqH2A6s8HSqaMHhnBwiIARd/hmjNMsVDPFBIURdFNBAO
/INAOeDz3IC6HxaovarDf8Q3Bnw80oY9kKzLBvWZ9KNkugZnlw7BGaEWcuLRek7UypWF9utRNg3b
UObLY47HaHR9c3RHuprQ3eRKOtGHB8P4MKXx5w/+wP3biNvEzsNhuUNnN/oZPAbWkukV12M//ugT
/HBa8s2+7hEJnrO9vPyeFshAGJsVdlg28yNrH5Aug4ZP7ASyJ0aRPEZjsc1+AqHwMcbIWMy7ZkWT
aJP2+x0qwOUS2fdLMvwszK9YB5cm93h5QVEFcjYAla+ZN/WeNWAAmLzVCzQp4ohT9KTWSTnPPYko
taM3naNz1z8Kkqzfe0ZQpFXus0tlooqoNU7jza6ppVIMm3fAY3uIw3Pv3P9TtlrCcxx8/dAy0Agm
3CHPFr/MCfjtotI4UReDFAmSd8NkaSSkJEBSBgSukewvj5aT9nsCI7TaONP8lZvwfh9mb+NXQ+S1
+4/lSNiuh/D73b7WipHx6Yk6/IdBWOBujHNhd/w1q/F5RoC3efCfERHJDM7St5Ww/i1hF5RGZXaI
Lz1OOTfZ8aX8mZWPJ7uphfDD73IMRmuhKH4ItDaaBz4OACDapHvvohhAoutpOdX5ehMKOD+uaQ/x
qV77hwG649HEn7uxgptYQIFGChGypV1KC+qm2RWfbEsfbkNRpRpUSuExj5OjH3Ri/7F0oGFMoDCZ
FeDRn8PwtmQpxb4K8Pw6xsZPbSmbr/rsiDvHldbGgYcJTEQQLF2ZYzI60sQzAIJXqEucjrkxu0ht
HEiTO3YkCUN5xZbewPzB+TqfjnxlYAaJCXy6TVs6Nd088ZtSWSPGSJIGTieVIRm5of9mxuRDse6y
tCGSB6esrOD5vEYWXUZi7Nw5FeLIYyDgHN9gZnHI1lZwSIHivEP0qVIBP2mWWVonuWnsvuW/B8x8
o4q4QXsFPQHtECsBMaMwZbydY1AOAyBJb6O1wtZRLHy6PiOyzc0MFj+hBRV7yfArtu9pWmmALdFz
PeXvZN81sKvsNktnBhmGRU6v7iz+9ZI+nyn3skeSsKmQrNbMlJzQDpjA5nw7xQ98S4L0Hsc6yWtu
cDm1VVlek51JXvHIO3LBHd8iHl/Z8G7UuyvFwSptsT8/q1RfZ78go2/zY0+tyoQ0dURg3ad3QO+V
eeKbRxFcwCpjAnr9+1GHJ+6XIg/bu7EQva7kqQS/HfbElvaxT+FiY2N0gZiiw5cJbKsROU2IJgcX
1Hndh/JCgodddatxbi4dNeFli/y/uIvV853oESXkFcDB8Ifx8+LOYfjo/j16aZTWdZRLxweXWqk2
6lYOHEg9TPRQYnFglXaeBhDCEaLH/vrLWzGUVPwAGzc4Q+55Ylezux9IBdB55LVfR0ETCYHVDpeI
vvJkBKFS2J3LtcERlMiIDG7nt2tM4q7rHu60Q/jQwzwVtSzIm5rEg910TOR0z9A5edMycQhg0/sn
G1TWHMITSZm4U6CrqRvf8bjIm+2p/y0rnH4fmEvfXP4RK3WGYzLOIPLv/CkDO2ij2+DyTZEMpFpG
EPLReM5aXbb4TnMJR55vDqbH6fBWpI+wAnY0o+nl6PDfhoqRjA0hi8idbwR9cEjieK8H9ca2qohR
lst5FvN43NzkQbyp4e74Xo9HaVfuR68UW6k0NzaGPnNBbNb2zLHXUKqwy92Fl1goomNjFDhFU9jP
/xqciAnqTIOW/pDJzxfL2YBKEONvoOazYtll6JAWTzbXKmEjbBNrNOAWbhZxhQFjPSO75aSLbLZi
Z6kg9aed7cFBqnuDWBqKs7PStzRnRqHKcf/r+ZpNGf5SmyNwdeGj/KY8i4d0hIDMpaM/idrS6nhV
9HjzjxkTRnuX2P0p+nat6AuagsqMyZ09JJNFFalkw9bjE0NNxqZvoNxFo3YPFtwTvwdBwNXjbyG5
JGLGsYUAQWnu1mZbAs3A/GknwrEotn1bzUCSFOuBYbxP2FiPn9XTtaGjbMJ6M3Tegp1e+Po5sKj2
aPJOQb+Q3pZrWkc3OzqoAoO/RDV78qZy0+5g6v8JUpbgxbuNU5jjDKjMJ1xZQ9yz4WtoAkY+10vL
HmCxXQh/J3wtUKlKVx3IFTbDLDGAIJcvR2eFGE2GAuoMyA/AmggwL+Y+c7etq6ZSTnySb90ULtlW
3Zdb/snS9Bz0woVYf1+yrQ1NaCQDXdGQVSxOZeMgzW4bLt59/S0yOiSJpHKeCdV5+nA3b5ZoktPa
3giUkAiQDyACN1+Gc4tL11lMk9UW3CpiDrwFx3eO73/FIU/YmgVkJtgc3BxB4qf9OZUOlLnu4Crq
uJnW6cMA26HJ12kLHvvYU0h6fk2Umvm3jExpEW+Jf/brPPd83U2qECJ+PTbLQpwadKBPzD0GrS94
NZ09N8bYO+U2XZ4eZb8xpUUfD57X0FvLZHSVjY7sGJexeojctr3jCg3WLP/137hpTv0W58DXfqvD
dO372uG4rn4aj+UCgczCig5xlexgYi8SPnHtMDFqa6wZHnSyW4xgp6JuVOUPWhPIDdRryxNzsq4g
4D1j+2y1cI90GAguOD9X54AyBe4OSAeom5KYX+KjpiQuu7Gjnk0mOuQu9dBigi9Vi28GQNu8O2x6
p1vz9sz8GwIb3SmezkpyU6KSS2IX5aVLg7d2WmTbAqkfbaW2V0DM/SEZMfkUFLw9frDOD18o+9ze
JSN5+Ao6ZxmRAU6St75ftYmD1HbqUw3BclhFSmYYYwfde6t5R4ZI5eJeB8xCE26TUE0cu4ZgZKKo
QhZYD1CoiznIp7TR+hNXMDm7UqUvoFAMsWFexcXdbv44GNTc+4/U76A36hfNDksUH4RyXsLH8viL
IBpCsdSQRnS/nasgNI2DmhYkmJV89AacnA1JidksaXpGscEXIiVq/t5dJm6RYVGStP5why1lzvQh
gvVN0yM+0vXW1dzNV6RQcRoOCspYWlNpxoFgVSokzVJG4W0SDe/xboxKmmMciPMWmLKYw0Fv9Ztp
VpfVIJ1WM17/UgpxwTLqPMlWlpqTAydaFkAeAThrCo8jqoGseWR/IvjzhI6x30cW0JBTCJmYBcDA
RG9JdDewFdJSFSsjTnU+F5BABxmHzqijZuIz8IPiEGVO/gB450j9ATK5HO3+pWOl/NgsfSPKo1xV
GbJEzhjDwnBYQJRVKIozKVr+r3WZ4OqFQoVyB+cQ85D08Saytv9b0GIHS1KvbmQG0qSvoVVWb/Tz
xlGKn7vKf1tvUzf8zSEvxiAl6Rl4wzLy5XmoAnn+Fjz23ldXnWg/VFq53C/q0pB/Sr3shB/F+mVb
kZ7/n57wiygt/YOPK634Ii10A2FcYRVpUpRnpH0EAPllDWE12NPlaDi9YnOmtnu3HyW4GZziQZRD
YyzxvjmV4VB3vJ7Gg8Af1O1Kt6fCBFlcH7ZVlZW0wLHyRZUXS0fIZFqpk8Oy1ZraKJRqKIgOLp1n
6GuzoJhV7dTp0oGlJIOOieRqmzAqkg93CnjSa0D0AQWlGgUt7sN0TMtq1Z9djrQYLFkT5SY1ldOg
z8M5PowPde2tqWi6c9vBUhU74eqvnOuBv5f8aejsC1UAyY+jzjl6A2LHbIEpjRM2DzfQZXG1vIR5
8HZxrBcpHvoUl+6JS4YVn4J6lurh3TZCo5/1W+4FGQgLsU+gi1PQs2PBWkMAE8Fv6orerY51lbPT
1QSXxf01xWA/ALFZQgW3yM40hmjCcmcyj8QrkY6e2b3JQTbigarbvXzihi4nuxQYdkgbCgxoGN3M
1fct7MXETJgE4Ru8k4oueuKNzI4Hd85pW3bxehYUBd84eszCmKh+epW3i87A0vfVf3kiPohfjxID
quCmgZ6kRVA6yzwpliEcDbYI6M46c4S0y5RSVbkBr96ExIb1mJWaO1nxp9Qaf9V0GtGbdEDujQwo
52wc5/uJWdCCMnt6XpcnEo1DpoJ4odqoC3ICCxilayQ+9ox7FCjERjq/x+pBjGFXx5etsu76sijt
63+UwjR6YCDT+BLumOQd443O5ndUwUbhRkNZSjm9c0UaLio+QdFKl1KAlBfflKzkyOiEUN7IsDMk
aFDN8bIf3a3JGSfpWgmgzJbSnjwHb+s+PmDmbj+8UIehU7Ka6/YXGQKu863jdSzFsckTi7VCvDti
T+9ek7WdRmBLs05BRiIvhMYeybag4QaC7w5/la87vXj7oCwWYEb5lCtHwG0Etqau0RdNpX5W9G89
7iq57IOueSem1dwiM0S2lxzSmDTAeyU5L+S0pCwshfL/YzvGGhko0IMrNi7m6Lc+UjuOw5kSxmQs
SEq0OLZf9kyyPa3s2h6gG/pvQ0lQ/Vn7czHTl6ZHSQtRmL57rXFkFQNwzNeuMRo7fV11VK59xq87
tIAXM8bMy28X7KJDSv75LK53iS0SVzeKqHdFCgNKvPzxWCyimiWUHz0mBGwPvVlQVdwQwBRN/ydR
rgjuVDQF+VYkve9/FkfG0ZvKUvgPELVZSOxFDLlKpwVCqRTCdrDoOa1Vkyuw5S+29qtzbrOi5qTz
4vhKAIpKiHgdCOed7Inz4Hw/OPWlXhBVyygij//KQJXTpZsdlNoHif8oYHFxnRSfDPRspedqgSYJ
Pk77RhIPQcpanapZb3i7HHgIBRMaYEVz+Fy5jBkv8hnjrSOMrtrrxWhKduNcceKgoCp64DWTafMk
tSXfN/+djEdRRFk9D5OpDfZjOYOI04/ckjzrsfTdVH6IxiYsrBhUQp2nh5ETJT868g/wxFtckzEJ
7c+7uPsipNVThhQ+a+q4uiWj8D53HsxN0JP4frHM1uoc+aBXWiX6WObLcghIbxkt+fqxnvqN5hsX
dj/RkYSljDZnQLaxPOkfz7XTUyeGsnBayqf2zL94LOs3DLAxSDue874nAMGWVKNpHJCmScS9CV/N
n9tUuvJ9yATOT4lkEjlULwm9MkXP3IOwenn2/sJcko9cW7GY++ibHxYb78Va5Y1hucIMGYxkAxfP
NXo63OfCs4Ooqq6/s1fkuW12iQ02rUGwRxac4/DM7OuY25yooGDKxT5SYpSrnzGVPLbPmo3c3/Io
RW5MGdzO3YdifoceNa7aJTIZIDLxcI5sJF9Nm+EjUntwi7JkdKt+mNr8lI5Gt1nizg9JLHIfCMJO
heIXFP2bSqfaLtWPZJCpuZeM2QoklAdsIdn7/qFMVc6jleaFvfwfUKlq6guK/vTfRHRbsPItKnuu
+CGLDI5vri4oNmYW5NRkEwNcT4xOp6t/HyVwVt5OviuRznLBWwKzK3Drdak2ajolIBEL88/eYuID
Er0/tNT1Lv3vFYESTVq+fmhmbh58y5buVpocJRHMnpm9hj6rJJWAtTOznl9CEpQJE29fF9dTHR32
gjWDpgsdMExeOdloPfPUy0KuKQSAr8JiEJfPM0Q7CXq+yTtZlrJ2TSl3YTxWuuigm+J3LQO0drnj
FRR6Si9UP2QyMsiWvEFHdiuIha6v1UIma1Slo9TW9c4c9aRR+/RKgxpL1JBvpqIzgT5yHfLh6gCX
uw2sP1FWsLFO1hw6tkZCgtvjr5CB5Rke9V1A9MXnZIfKJePlaRMhauLhsu7J8W4JXlXHabrKk2ZX
ZiNVrShdpv5SI8bZiCY5HOhJiZ5e9nOrN09XALjyZfBK7N1NBEhnC4z1cQoueOYbz749yMc76lXK
kz8ajkhMldaNB9eNSzL7nnDZm9DOtNOq7CJ0ERuv7DX5mW/8Y+VgAlS27zkSzJ/5mQMUKubVxLd7
nFJHXggl+YyOIveCx1xBSYWWZlQQdnRhD6HiTenNuEP9IRojZIt2y+Googk55dD++snWv09nyE7D
zDtiG8pC+7RziPIsLPiAyqMgZDj3py8il+8Q6I/P4FTN1ucBpU5DJlWy/5vd0T2hlhaTSeuyTSLA
9RTPE0Z+nPzxP+UOX0l3BTQEhx1PJFEtDYOWC+9MK4U5VdnjOhWGddm9ezntkQzhQqugzXl+nQgQ
xnt7mMRq5ZOXZnVmY4gbGNsRTJPjHEFicHG/SqQXSSJS2FoUDYeLy568FMQjqqOrL/Ex8lVq9WPt
6YWblXMTNy/CEGw+c0DpONSSSy1F/H8+uoy/PdBT1FNxQyAZn829Sx4q3kyI59PNL+OGL/Hp4KYj
C/sdfPsoSSMAuIdmLi21tnZxlTq0jvzV9iMH1zTkRo/D2BMsvKWnJ+cJrKgXsV2ROYEsf7kU686e
m11sh02MD2NW2jmLOmfS6dFRkD2j2TYUGD+146efEpj3LHyuwKoDFx3DKZmCGOk8IH7j6B5lDDoB
KU0QazgOZtGt6IuB7+EVBYX/Ku1XSnD95M1WDcUcZG0UFGwyp82gH7AbifaN4k+vnk1KcQUXfrVD
3TkhTrJgk1zKO0zyDXb59eFlGXVd2AdEXQo+i+VO9hiNSp7y/YBQot/eLLbxlnwS2akFvFHocYVE
HONHll6KLsLRj6DwEfz3e8Cvxc0MM1/Lpu4xhrDd5P1M1Zph+yj/P031qIY5S8Pe2y3kuE6U7RTq
j9nmuSy5GgheYo4gnWJsvOyhsXVIviNDAs5Hs2ul2NiSM1DvEklwTCgHGr293QwVjXS+sEXMuo/t
7giORM1YH1ec3tAO7AtcSm4yM5Xw4CHtgnEv3fWAwsZZsjzGLip+cQiMzKJrrGw/6kSbI+e3cZY1
FNLiQpUH75QF1bZN+TbYkLPziaSoQWLFamtrlg+tfCRvbxVqzrTuNE/PJWLg6yJxMyQi+9TL/4/K
dhdApAR/m2Qst4AnvvjZ+EopTZTExYu5RM0JKeSuAZVLfPxXkDPIJNhikIoCAx1Xvgso539ATqUq
RBx7UhiKbbBT06JNn6vX3DN2CFfYX/7h1ZGqSaG9ol+B/kO6LusYpbePSKrBqlaqIKFxWUOUQ91I
cSaDQMkY2aiCYFHxybJ08cngoodi8gjxA9txRzqFZa0dtLhgTyl2kNu7B+vf3xbXZ7c9ghTmVswp
y/lGkbIa7YWzcMKF+QmxC3ifDs0SDavr9kIQCaUcmODNm3ceKMnd9rIuYzlAZkgtSlcUfzoiU+4o
QRK6bsM+5agzNMptgr+5r0b9KfyshBhLiLz71H2YdLEKkoco+j2CLY4+YaDNHQudcwe02gmVDEh6
41XL4L+jGEd5G4kvK+10aMfE9vPVKz3bRbI3gZWxDRaHMcR3+xI0yGcFCpEOx9usiADhd78NCHWu
87ka4/V6XbJV7m11CRz8fFp1yzPn6r1fID5G+o2TcmZXOTzrBSB1sxQydLwALGOq76mvGUmp/eTF
1J6fPS8VTS8yPMC8J/f+p8FLz2mBeU8kgFIRp8tnNiNE02QSQtjdWcGe3ywY5LEAJSEauCDqUxQn
/slp1IGZ9FsXrNKo+tyd0Aaf+u1lnWx6FNCmvMY5nWaiqNuHZUR3OfpWh1b3JQ+oTZgs2Ke2IKuC
q00cU0YWox9kTo/gu7b1++d83SEdTj2SFn9tJqZos9Xm6XJhJKexvBRbw16EKVqdNV5oHcZMFUbk
GgZmUf1s8teMaleWaUJrzlgwY/dtqI3ei5KYUUHMgNlRz2W+ocGTAHGacgXZmFS/Oj7Gc9EFEB6E
BqKc3SmGzTFM/VHTDlyqFWbiKVdxCBdkxwAvgCRC3Aow6u4UHfgHCLZIB14LBXdQb7Prxhb6oLnu
x2D9c2OE9Sj2Xl/M0xeL7i+UoMnmazQIljZIjNI7GBnlmxOHty+eEDE4b+qt4+dyKUwVmKfIKH/N
LzEogy+8GY9wIWB6+yBqvbmrMShTxYDEdwNBe0j5ky2hwIijoSHGsBsrfeoZKA5arEYSXtTt3+hi
R4HniMc8B+zabZnlXPe7xhOnY9N6YOEZFqWfJbnrSrrJt+VC4YSS7dcwk0jQ0Z5DBPvgr/N/0TZU
kyp/MFc+/G3qVkW0MZ5eoCPjA3h8nkvdQTHSNpt85dxdKYLvMyYdFFAsjA3sE5oSLw1IxlSb34Pa
UnAPhzPQbQ+9RopuJs51I2BZkLzTrr/tUhb7xuUTxV9aTSpBJkvfrAbTqMws3DsFeV0YCqNQ4LuS
S2BQMg0Y38CHIUbSS+ee+NER4NANp/jqPmvUv+eU6MoJt1VB58zUDBiDLrSgSUfye+/9hqPUlae2
brEX0uR8eZzNiu0r9M6De8olFs/44LzJFEUI1kJfDjI/E3OgpxmNFYsfhJ3diodtZbo1+D8/Yye/
ck6JE8C0vkjB7oOgbDWiEgZPhBaQ7NeVyoUP92T4xOTxKiejkqXGuxnkKpOawPCnvLR9EXru+ZKJ
sNdZpQyIpa1ezf+l3bDMrfnSN2mO4hrW1AK8rHrl2YAn0ERT0An9pu6icgHdxR+ZnNCy+2xTTXfZ
tUfzmeCMjROlEi7c9BWLBJl7Ld5mfYHcqbdTcjmsFoyPOveYM/CZXLre8UYeakz4gEuZ9Mb4XOW0
m99i0I40AuEC7yVYrtf3o0gAXGlZPCCIxWPijLFWTXsHIuUv+NFiIKbmxVCC45uQJF7ZLKI3pQLC
ADRS6DH7LCHk21MEQjJyfvDOc5MyrE9XBeGhwaaJbI/tl92QpVb3kuE/rOv/OmmfdE1tp1sUyBR+
/wJ/PAzW4OJjksEjYCoGuPlJOe5q2JeS3PUvPVdHrJaSNh/W5T0NNT+pc7GiE2IrUOj2wCSbZqgX
iQcmF7U8+k7nHb3spcxPfGZ72JWivhAemqMmNfS8bYdjxumM/XOoB0vDmlw0iQHBHRoQKoBIQ3gM
9hubF4P8XNDv58twet1fIlRLZx8QXQBjHThHCC6VGsCaHBb8tlgld3r0WUMYKJikROadjNgdIgXU
RDV+X/3HSTf2Bb746aN0Xys1Ms5DDko6poEgdDcwMTQG7/9xFc7vtctKSYasahBqwfV6c9Kt/qTJ
0qYoEEH/7wPjO13lDNBjp64JS8pTh/H27Uodp7EqqnqPqL/k40slxSXzH30UUv92KbnDzWiGqsZ9
9qTFWca0KXD9yLs36LclPMRC9ng7HxC6JqaGdMUM9eNxOvRzUXkr8ZtWoYI+TCT4uSRwpOVNAl3O
VEnQISf3H4ooF+KgRjLv96t+mRIJFaggCgcyQ4zYiX/CK4vE30Xqnh/I8CL3Nvh8equAg98Psu+j
8kvb8b5HO2HsQN32ACAHvQhUlWKey8Twe/BK03eFn9AKXsxcZp82qogxNEhjKAeFGHWpmi+ncVsV
K/et8QI/zn9afrGy2J5VQqUdN3qakez3xfDM7VKxBEoj2/xLSSu8fWkoi2k9VNEVdbqxqjvn0sOq
X/YWkpNJv+Mok7N1T81kmHKITiafahDVR0elBsILnBbZQQD6n2r4VMAfoncR86YsCFg5xUmD9xXn
VyoqzCaG+jPT8M0hKDb4joY07AHWi8aqIYnrN5AzuxvkDQV1O7W+IIU3MPeDEpRCw3TRUJmKoCSN
MtWEsmBK7/QNoPiw8lqz717Jpr4bpugGyVkVTZ86v/tMu9L1+2hnDn36pK+mZJUPS6b698TSX8+L
JnjKE3M2ZoDLV5ya155NEh2S1Jz7XwkHalqNvj7NQb/gNyDsfok5FnbgOV6oWdt8f0Iva528YkLz
2I48arXsn2rybheh7mvapTHX49yl9SGaogdjLKMWV/7M3iv2RFIuNHJ3it8SGYD3aG2IS5SYvj06
r+nXBobHllpQKxx1vpiOlfB0RwGBr5nBjwbOhSAiZu4c7cKwfqgSS/jHU5LW6Z3bw0hhstZcNFCZ
ZjWKfDAFpxmlK17WHmNB96OFkL8W+i7erNOakuzbnkFYyKfNyspJlhR0cubgytjyD2FpMSOXLtH6
qsxqY+dt2riM5wGpG4g3VxlXCKJDHurvyrHApWEs3u08SZ20mxJIl4Ghd2p0g9/u8tggkE7APR5R
Ob9R4QeaE+OHbm78VeU6dkaotFX5/x8i8LR1PoVhE4JmEc7l9ta2Kvp+Htk85XMMlMnh8x1Oq5jq
k7RgSkQ0I34tVt7j8EgNT924xyZOpCMRrX9sBe5rzVKBnZzDqnBZftJjmpFFRxGbhOawzjpJKsBn
GKF5w0ECWzICPTRkZF7vYcpnlGoIKjyhaRI8554r2NBHxkaspAJTaYFFrGdrm9VniQOSGuEE3XNI
sQ1pKnAALP8UVeL3uQoIG0pepvYCEyGlOiHlvWM1MYm/JZKbWwBsGDGo5G0V784E0793T54aMLBy
vG6tKHeHOj1lWy0dSosI0DboaeMdnp+1/jgEHuHQ346/r0qbvgRl2J0RAmosMNAECGPRd8WyIJtR
ltIzYkJ8C1rYpc0VvOqNDJ4JSNGCaOkziTxFrx01xUNmbgWFXBr5UyJv9MDXzeVZR5xj0IilCB8U
8241RU+3KhTkKt3lNDFngZsckGhL418AJUoxIZqRCP6Gvb7aDYmtsNa3m/6z4fzXDmO9YKRPLRd+
pSB+p+3Ii15RQHPKFsbHEr9twAgD5KCqN8NZ/cmDBeEntzRvaT58FbQt4nHsTiKN91wBiRy738Xa
l9kYGCOcigH5mCrlrKHxtozScbDoCBOML7u46SA98pbJYJeLK+Q1cALIdvT2RWaOTCuovtp9Q/Y4
8mNc5ySyd5TBZH6OyC0UV3DsMEsWwSFkesGscJ5qhOc558DcoCz+IXVu8GRkgT5UWsSlawY/mbVj
AsYGlZ8JaLVBRAcDgzLNjQqIBcLkQFP5YV406nsN54rcCEu/ZQWTnCvwgYTsoCYo6MdyEdDEFhU7
olnD0ysVVDtURL+n0QLLaZECgEz3/0EQYu9YhfdinOyaO9I/JyXIpQTPxfRrKi3po0418N6rSEdq
kRt1xAbU+wCbt1ufFDMsl4nzGgGpQO+EgsoQD1rCq5DcPu6d5HIvpcEKtEIPjc7yyi+4pZmLnoXd
35zlp6g0vq8/gfE0P6zXqE9Icl5t5uJYTEMLiDGO7mjFYZ371m2oXf4QCB/FTPGGGzr1x7J66sU8
DBSkK8DomW9wGZm263ClUpmIdX6Gl1YzHtbEPS4WdMTPU4SnCf9j1oc39T17dO6EZ4vdHH1Ahips
cbvTvtSYDspMQq975URDG5qsKPVTfie8cT+ezfDbVz7+CSwvuYHzR8q0M6VNJtfmBhhKxJuZ37TR
JSOrl2Laa9IwDqVrUJpmShkzE0d6xqdlz/VhQzoNfuv8tLxTTWO4Fj1dy6lqVyEFyWtm5isfyoYM
NyS3m9iCb8aclzWb295xGcQ4GfrYJj9gioBSA3t4YkjCI2y3pm2Idpyt5drqmos/RDpxSI7tJRmg
bsOgW8xIgEGHHno8WkpklWxob949XWZC+G4hfW5wFR9Ux8104jseB5u/rv5VU7mvQAzfzXWVTR1x
nd631ll5lJthSiFmoVjLDGRlSFMfIQHsEC5UzhSqInz3mczP0aIV6kx6m93gKsj+04lHL+YuYpKK
p+Vak33ivdzD+A57jeVZegsUjaY72pqHmS+TFaw2bLWV4ZX/VksH658JP3shPY+ucZC97zsZi08I
x1k4v31tuDLjEEzTMKpSG7FB+meUSf3A7zJG7nJ56y04RYPNVf2C4PFBFN5hujL90bdVxjhP9Ike
abnf6DEbVLjCNblfJN2L0OEWMLz0KHZn3a8q0kcu5VaU9sjtpxWqsO1/6erZdLckZZu+c1kZdA+9
CbiZz9jz5kr0VPJRXfhR9HurKog+QW3d2VR5agln2gYs4U6h6Pj8eev6hYILFtJUbrXhTUa7DRpQ
7+bkMm5vbNb1Hi8BAUlddrzF+hu4hXM2+taoUOa8oaQgCaDbvk1tgMFnHwqlp1ek6Xv7rmOjbfhr
p6mxAhFbRgh+Fv75kTPP77d+L3i4B98fkfMLp4qLW8ipl+33DqhGpqXuFmwSKqHV5WyrmMeHMliA
MtBBbRFXWzpcl0Xnnryo2L9hDmtpAW4cTK+kP861E6n1OwBRCr8vzbqhHcwG8frOwaOoO314JC8Q
GuD/8dSSJl2JEfAB5fWhYJKCmG1yr+5Mnu+tPCsbGHGob5zi1nrsF1GLA4fS5XKKhJt5AdMgCudb
SgZU3HTnX5F5CqrKTAsyginiBO80ZG9a0mBkpfKyeeW863w13D0l2xEzvJKQltkWGzrtnHpN7HFi
Q/smDZQXtJxaA4qVgIPnP6s/BhMn2lMNyMvddSeTJeCZRZk2UwTBv6cK6OTGRvBtAA4ka/6mfAje
DBlm3UGtYoOOZ7uHKtYIGHjNT7NoO4Rh6G05ffmS/GUzW4mz/s5ECnjmihFTP8yxBT2qbKYAxdiL
7FvpvVOgxJw2xjdifPCFMu+1IlTJK2yH50zkJayefFYgjI8T2ns2ARc0CgAM1h/EOckkk/CzAW+d
LXbBtqSJiLRFTuRvVbjgcnjyMdY9i5ksZBku1FZhEXLAxFUJDrHzyV/FN3Is8H+qSC/hUnf8kfCb
EWRGV/mOsZQPhmb4FicVnGchodOB4Z5XpKQqLqCRvMenSuerGFOYxdjBZ1nwT/E/mZFJPdGnMSE6
cnFkbtVCRLELcgz2e4hFvqe7bMsy1y6u2VfihGjR2vGDjMtY4DPB4ZmTPOfL5DwJBX4JhhnYnMDM
G5Wlwqg+s+fHSsGfRldoN8Q2BNP6tRaz012S5o6JKbMQBN8Wcf93vPTBNXVT7c+sLa8u/XEieT03
zRAwawvj2tQaSsdkAZHa37z9ekN2bX3ZREbNpz1c65PHKPhSvl/wHbaSzPnX97P2Czr15BL+F06S
n+N5MivsAsi2nvZVxjw/SIqs+r40Xbd9FibuZajkL4lNL75Sa/Hdh3fTwdZgdOATGvvQC72SCjdC
b/3ItCuJD2L4P0OkIV6u8rADTdJ6225P9s7x7H7vmNGK9maL5ML+DY1l9Djey0z1dKb18cM/jVkU
AtHYLKWto/USy1RoiqowspuLczxh3+M7pjvhjpg5eROtk3kMQ4yqpyISnRx7JpGFK9qJvfpxyCx0
/3wT80h6+65s25r6vwRnUX4Zfusp+wj3m/NF6CJvWYe8EhdwFHe+LVCXujluhJJ3I0UxCcNhIxJr
Jzu69rC5eUYJ727tjGtHZOpPojZHPLbxCCHkVchX0IgoyrpUPNUgFZQvZRZAGCuNHj4pQTuJR9d3
/VbEmEw232LczAsBaA08P1YJQgC149vnIY9rPqtxphTkf9DbP6ce1tLrdYGTqtTuUubV6saxDD9b
5kHl6zFlmzEafh1lgKaFrnzw6iJKuUI7GZ4HisBj42YObZ0J9Jom/P1crhkriCgmWeAPq20I1Tmf
1awXRBm8UMs/NPrwP5gHwfkA+EmaDkZhFmofoCnRFvSWrtkMfjtIh1c3SIOJ9ZJH5IuoWCEGxQAs
jJRG349Mci70ttOgggo+KHC4pHm+AXBmNspQtWSHwNHSIhBAFnhEZ+31m6decDxnqjT3zSf6zhE1
bfCV8IkfsmVZ33JS+mnkBaq1UjkkaIgcvHfVdEIc1pKqUxrX0XUiLmosbD7GkSGf8hbJR3TKMleb
rrwwnCOiUhkDpF1du2dhCPSCdCR6xnEqDrwbcKHKNoGalS3w3UbBmxPeHfuHRa0tgei/1DI32z/N
tZoRljEkSUqKF1srpG4I/Ssxpk8u3E+8I6ZHE32pgMgJHICC6T4sbRY9a4BNYJywsg4kpWDfaua6
RkwUjZ78EQVVRs2+8rPd9Qot7X8YQCctXQbF+dVrneLb3n5WMvT3fDk8uWJxpjiCpq7YHIK1KRZ0
bNvoIUImYJeF1P7lOAw8jelsFb8wOLkptxjlmkXcqbRgnGOp0wQCmJiBE9n8CyfiB/lva3u3px8G
V7TXi98Fxvs1Q/rkqM7ZOdRzQCh0AiL856a5PnPhn4ULVKZNBeGOwX7O2GTqv5Wa1lpIZwo72Grz
z7JI4XGP/JXDDHHOSsiNL4EaSrkvALORc6DmDc+MCaGYUYLOzGeqYUd/ujakskW+dVCBJUGpnC13
U40cSXvB/Mu3A7Yv2lMOF3wpKc+s+ZlxKGKGTSQxkEo16DHXorolDFSxdJ43tv9vDr4uVGVMbsvf
pC12EqnX1iJjgHkQBogDu4Tmm1pskSSnuYPqvqd4WDR1XI9Lz1qN2RuLvZn0TiiW+AI2yVcvROto
83/H42jgrljodprRHXaz5jeBwv0KWp2P26pNOQb/yztRbIyZY4bl2kspxnkSxndqUYOSXU3zKAfV
WrWxGlW10hwC3GtTUOPtGzDtO8ra+pljdXQDP1kQbn0ncJRZtm+UL/QITv1k6HOK8Ep4hsI1RSfZ
XXojP0yL2TH14uLvMjd0+/zdyRIA3MxMIT3tKIZZr8aB4zJeTbReO6isaBSz/mopG3zt+o8wXJzg
RSvayHmRaCUHRyC4nic6GDM8Wz0NqkfAV9A6Fbn01SqgYc9soJnEmIBcwDHcyrKD7Q8lNpCNqiLG
aRyfGnAZRMWKYMsTJ031juR9qBjrDZgqwhVraWTfsO5ylz8muNgE8Gs1BxermctP7qpjYhe66wIv
+JpTHUOW1A4N7jXVBPmxJwZpMsF9+e+hLipNCWjK1Nx2LRDxwGzN1IuutaSS0iF8ZV7YEErducpR
iPNPEizhDvXF7JhZQfHvNA1Ac54ZcN5r83lWra6lzxeUhgJFGkyK51oh2JI8JP+m+Gf5XSFCy1ky
C+7g1eHVBxduyLOh8RsO2ZXWITv8SJm+g0LcrNCoGc6z5GOS1NsnstFfPY+hbo9l7jQfDtg8GeRd
qKleSqQ30xpAAwD6K2FlJ8ca7Wwvk45OWDdQ3DKxr6xyCcCdxd5HkIH6p6Xm944RcjyomaNNljSD
IKiEvWxC92Je5s0xFAY6DGqTk09o4orepmdkFf2AHIz41DhECUZtsPebIEcXKNri7Qy1V9KlqMS/
UMPIGUusgKckhmgoluhH0eTYLmHBF1Q9c4TRwj/i0AvqhQsc49otvRLMEgaBchskLOZ4uHrc9dbc
KfevRh2qQSs0lAVIKOBJWHm1+tVL00vqk+CYuNJhNZKBMBFI9oNThIVQI8U1hE00nsfYckK9GruD
+pc4JkM47vcvVnZMYrBTneafJhIcwRV/D2Ukk8mMe+sXUcWxWtfqak4he5aBg82wTjnfx5Nvkm7O
gRPR6xC27B3S8SsLHFDmYBLW/U7VxXCOJXzfQX2qdjGV4WjpmmgoyC3qN2X5OVJ/2PYCN3oH7Nly
z6uTeNVErdUvH/8X6QP8PRdYzNjpT/BmrlpBpSA0xtFm+yE7Zds/xOGF9CzPtqpLa+bYzMTPyZdd
eAUARi+Uy8iB7jDZHEGVjGnbqZIRASsgn5mCuYPzOtyRi4J8phMlmobBSDbXfXF8LaxIVz2msVcY
qE8EFELhyOHtwqLINTIsUQviXARCN3wjv3NNGifFrJ7roVru7ciiMYU+aXFbIVb66rJw8Ez/jyno
OI35VTDZxdod3LfuW7weCDLSdlfbKADRRW6RSDo48XpIx4hmtTKnm4EzaBIh8M2Ie1HsuZVS6Vbz
Fk0bGH+zxpjyF9ObFVUAYeC8fz49tgn6RoxxsnccN5RALz5nRwy0UeuAWcNKfrRT/jHKHyymC0lV
FSoh9cLA3unDkh+s4QWMbtBj63dZGtd1yOsjqWf4ED+o3Y4eEW4Lu1FkPlFLtxboEFKP1d+oNQiv
xqS82zj+S/THrAcs534rYiI0xvVWwFP5orLplOYCEFMr4AD2gcLEOuXsfjARlrIGQDLtXA/fVs6q
l2KkDtGC2flPoCUXeJsZw5Avzx5puy+PM6RkrW11A93RW9BsMPw/dqNDlHO9fcI1oG4ds2tmKGlf
fDe5QQGFe4W9cV+6tDg5bUnOnYQmILMur7AahSW7ySoe57xpNP9zz/ge2j7IQr2hnNma44f2iDWc
svxBjCL+d0+8RsrSmQjpGr3EJaIaoRzVoNQ7a3nBk2/WYXqrvNfCvhQAnay3IdGXahB9BC115KZ+
5mCsX8V6fato7qI7MC3b2YCtiMRd/6UN5FxDBrOP/nTm5uKk0kMCz18QZLIconnIXmQB2/pPLbLx
EaKT+r1jRfEu2MzAlor9tQ9NPWmtQPBs9Ptd2kE6Q5DJ3rPx3bzlIkD2vmIHPdHFwmYeZDQctAuM
7jpRVsoGyZ1uYaN4t3PkvdLvKV2S9u4DJx80cTXRQucbCyzuINbOEYN9xyfN0FWoUWb3zg0AuiJk
Z93dFEK+yvevqvcMwqmvADsvUT5AQMQLzJTElZhfzPn12flydTcVb9T5SRfmvZnDPwtF/rhBNthb
1npvwblo8ft4Jsv536nkByOd0NZBV+bU2saySoqQjfOYNnBYbtmWDVItH7nOLQhoQlBFgQOEr0iL
V9fAWVpUIelS8IDq1Eu6P7nXuzrHW+0ubnFPTYsI1FLoJGinXvYW3tiee8eRCJQBN9r9k46J3II2
0xB0dFfwSg8y9tfkpEET3WqYX3llT5si3RpQ7hlgKAC5JYAIEgNeVFs7XIMPbPwt2Jokn4MRP0cV
14yDhRI/X6fbKBo7236PAZD34rxNTV70grlwxYw+z75Uf/WHd6Rdo8PbGqcI8c0gUXTPthVqqXAV
PhDmqzqAM6JQkxZnPXjMlRKrMGbT0hs+1zY0VT2ixC7IsAVyEmr7kf9aPAjTBjEruFrMktpgMQMo
GSPfxUE83YMtc//6aFPgRSTtZrmCERs5dGPpOWFmzlwCYqtg8B+M1OUP1ZVh4+QTlcAJMjp/+rtl
id2ei85QLhGN4ZW9GgATPgTSM1SpJs8OJYNjzjejBIs7OwhFq9+wTWjKV9DRMnlWKNk1fVCKmHmT
BXMP6uC1Dmhc3SKdnMBSjAQEZNOkPdhY2pqMXecu6NDdxQFjGQGQh34N6G5oI9qDmkpeiGIfeQzf
+Gf1nBWxUvstZrbHu7Y7kS4Vtjz+nNKIQCTGf73eoKFl4K4QBOIOrg7DNNxjl58cUa+henetObkF
1Hktg9VIIkmF4jK0feeRoYxr9xyUbjFsZqqE0uktR0RasoQYpGigs1zkosnKHTRcQC0GPs5L3QQQ
CJrmSt0GnujfoRfuqZaf77QiHaU1D5WD6TozSrn3BEuHN0ZyfkZeDoJIGeXZpzeyXILzgRnjgbGa
v+B0973zZKnQ8CQaNWHM++yMKiE6Uv5W5XEwC5U6UV425SilxDNX9mPdb4CSGcbfYYpXtL+StkIl
IpTxhKtLajOJMy6EGDbVFfoC4TGUp/PcFuvrL+nMptU6KeEZv+l9HBJ9q2EcZQ+CTuAe/CtQgC5B
figTXO+Mqj91O/U1A1lcY1Y7zdwzhxCTd2tRwu6o8FjJyJggpQi28itLxp2wgrot2yl9n5ynylB4
EU3uClLyOBj9JCayDkDlHXx+y9zZt4wBIcd5mlRnyzVN3E3A/eDhoSrbk3eTqpPOZ7PlB/Pnsi4S
KYDi4s2g26jUTOZl+6PACA93IOE37HwzV+ou7qnH0ZZdFJ99Otu2FsLdFwP4kyrbScQX53qXEqHn
FLBy3Slx7gKMQ7MTpT31aeotwZuP4y0bz650SKEg477XqnYGG+ek23Nqt54loydja3ULNIFGgvhv
OZt2iAPk3L5ZYEzXMZM+dvKMuQq4IIZfB40HIzrMJuh+q5od9sFZBXe1LMGKta8h5AKFeiytHCoq
rYq1XQAsZnXS+ErCKIFGoYLxSq8XOtIOnXOiBQCQaM1gzcnxVnpQtWUw7ajlWgivIavkBOJPEuj8
xSATwuUvU1XuEJS66c8dd7axRwhiCMhBB1z4nnEfvvc3YliycIy/SRjTDdb/MoNRjCTp8j0qPLIB
xKhLt5vAKRSYzhDvE7nBX1mArGwDjd5ko4EsQfZ7NDqA94JHHA4Wc3QFz45Iyt5yxhDsut6pVczw
ByRTSMnqrCt/zmjQ6/MDcKunQV/diYtwF44o1FLMHXYMWjuGpDiNDLxp6+gnX8Wrwrg696A0EcYE
IjY0DAvryimiUvBt6OeANYS0ToHk9NElO8rpOAiBO2+Xgr4bEhfcVATRPUpr0Tk7nNw9Xpu67l9Y
9X0tAz79hlwAMWwRddCMPVn/lUHsPSZWJSQOVAY3nsQqXlk1+aP2z6vYeqa15RzXMR+zFSOqJa15
UFKhkSYdBwYhGQlQZHPFzwuerm61PHE07It198vD2YVXK8VpWGWXd0nz1ErMuZM0Eb2wyD2/zjx7
qNoR+siu+MpmW2Vh6oZ0HDQih61rmyihs2sUlhqTpRxgTf20MHXELAbdIJ0X8cGTpRjrGxDB3jgg
1O4LmmeBleGeGc1XiS2nulBA95e9FWC5Gku8txTQC4u3fuZZX9bkTLp0U8PdH3A8CLwfuj3GUfql
exdOe3ySfBd//gOvBJSzDzaE1TyrsBE7pvhKTUBAJgv3CpnwolfsevKuymtF7mS2rhVFkMpP8ltc
uyrrtQfqJlrh4PCpn00rmBwWteMgIFj4DX6xHaWywGDaSvD+zGYvqD/+KN1u6iC2YOTfpH8UHU2L
M2GTkqCzhYfRToqKkxIP3QTVctKF8ow+t4a3USekMpprzgHn3XxFSGMMXNzB3d5o5h/fowWU3csA
jyMhbCVUG12p3mNSwEnJHRZhV9bc4Drwas6vOWxoWu2IxwloKUOQIKCMc9PBae/nkbaXYi8usvUA
/GvWHAJsjKoLk4xtYpHZXO0F7+m9mIKw5GN2mYJSo62J2inl6ZzeXDuxRhOCGBj4JhKNjjOgW8ft
BcLFl4kfTJDR6+4SEfepyc4I9jIE9tIjgTnFjQEfHq4ZhQoLFmfcgyCCi3t/8Gak6LA6R2J10+jh
ZhO5c7iUgnG2cC0Xiu0kcqkbQSdecjEu79i83/a3sXz2aRtGRDR/UePK5DI4LGylmLRh+7pgFpnf
mKrItPhsF0mlg4mt576H/YNK5j9KJvUtCz10PueR1NyhBuR4evrruqBywY28WCFWIpZvkUSVRNsK
xovqgUWzCXPvNWIJBng+YjkWM2CVpSlUY2xIl5xEABPM6Ioi4tAaNXzWsR7/m1NcLrSDYSQ8dJKN
li848s6pP3reMqZRF9mNWG+vZA6XjyiTNzOt9Djl5Q+/cslzjUGArqAmMUK2VDlVOQbCpbXT6YII
U0mgww3pPBcv/FDOkOsyiYAQa85shjbwrBWPcT8GSUhDvgIjeLrwEjwIZxlzKUFtsDlMqydb3fYM
IYh5gGc6gVQs6OdtSSa/KSQs9IWkoR2qFsHayQOU8HZwIs2Cp56l6jR7MG/Goc+8EqkyHpAH992u
I02jM2v6tWRcESpJHV1w59z7HwaBSe3flUllqvahnBBwMnhIsmlC+W8igCY1iZEvFmVTwjIVBPFU
IZZMsMiTGLsrwktkLMVqJqXZVijzvAMEpLeqMwVG/+e9LBOzVNjS08m7VhfPgw5r2vlUSLaEfUti
Ms7/UbcPWDdxhM4I2Y8vL2Hfu+v2iocb2aSj+aaSeshXU070nkdpRBWqOipg1rqArikDr3jByNJN
zwK1waLuNqP2XboB3cnxfFDaYgmzLts6KmB/8gSo12HFUcItkVO9+xOxyjpye+iTlrdDbxekmNHV
hXLm9kQAALnsa+fDf9olLdu4k3Pb6jepXbc72R9K1K5RNf2uVpXMHICm0LcR/9FlfOOPKP9nFfK4
kS1EFnKC4Jp8jSLLI3FO9xEve1gkEVA7WqA+3R5Wc4cZxOrtUw2eEa8+acnzX6XxMn3tjuGLin+S
Mb6h7x1//3r9ejHBwtUb8KiAOK53VcfNSUxP1gyePaSqRAegQePeapt/dzdg7PHaz81yyLRmEQ0T
jE3sdsdj55MnTy8evfw4V0dsi56VtexTAE8LPQjvN6Y2lkuHaSezAHwiil6jTCqHHXy9sD8Fc+JD
VCngXG+bmiraFqy7AlLBqsyL76cllbEZyQNxeMHwbNkrXMXNyz+aFbQd63Zc/bQHoTqilNgaaHOm
dAzfHqDVrcMrW2I3++0s4HPeHP/TNH5yo4hBylBJQ2h1FjOXDWLF3/y53koaEA0nhdKmlwcQ7gbF
1FoAmbIlPyHlYwUsJxRwiR5cvwybfrM6i2uZcnxrDBjMYIbFne4/JF+tKK0phFcvJlVhEUluNH1t
YZmrj0Pz9+TbvoHepM+CDYAsHkZevw+ulfi3q1AVMDT+djM0r+eBKB0G7sTxlgoTCapjbCinm07k
VukA6u9tTBCk2r++vRLUUMNkGOdYJiwlLCcE9tZyld54BpxLqeUXC1zNw0/0B3/py69TeDidsD35
H0RUYW4z2CPUDqCo1k9xxWPEJzM7kx2H1glPIw0jexW0zPWn/wFTe//XqaK4myeyvQzUW1vBPuW+
Zw6oMvvOZwrWrnoyglE+WTIotuWu89mddnA1rsfhNbsPLW+3BPL3R6wfTozcP0poJruWfd6Xj6sF
XrCrOKeFGqJ+O9zLorCMjRhKVjED1Mmou0hBPvuhG1jrSvmLgWiu/HuWnRO0tGZ3fpnIsZdPuRuU
6kEwiS6nb093dnRwHlg0ZQJBZMhfMg0ccc0EMUcYl57e4sGhcShnaHBb0VwqfvZFIy1U75Q5Ksan
WoxurmxWc/+6wwz55Zv9ndDZYwLpAsb2NdaExjdNqDRmPi8hdjSbu/iUns1LhstFbeYMUfe++6GC
fS6MJwwVqxrORFDxMXsYSMiBjqIbB7rUT6B0sq+x5k2KU4u7rfROhVY71CfkNNeVjy+hCQCIgxGY
SP3JRdSWtj6B4cCvv2AHKQDfwSosmaMXXCuRXVcEFdWgM7FgxzNLAHgA1pkcSpIUF+dC63GOoztu
+4Y5D8xiB5q9KvHBzbO1Ste/r9nRuHFDm6bg0uEGN8LaLn47IkZVVb1wkKoRvqftx2NBFblh5G/q
OtUdHhetjfnJ8KnJ+ItSLZRRFr2eLXCnFrskrhxR55oxlZAanp5j6ZpK92uzQ3ECWfGAU9lF9MH5
vys7s1OJmhQM/5SftZ2j6IDf+/4J5DNiU8QpbVPlGijcsZoJ++Z/Oo0Vi6mMQUACu5c6hM4Q0E47
LI8h50TBYrG/foB5xR+7leRmg9FYD5C7D1EO7sRcsSKb7ckB5CkXT24jkHeEcgsCnYKg1568vall
I538cVnDsLgbtF17PuhmCM1I+6MRE5SK/4VoLizozKs+VvAEdk84jNRuILtr3qPN6zBtCWXXhgSe
8liIY2oli1Ctu6Ph3Ngebo2/YmmgdeO4zYqy+a/mD/287W1DxPomNZufS7Nc7NNMSwwCB0LIugV1
YdEA1EbLeqoWpSwa9MDsbZLXqa+la+M2V+53wBq+QmVbtq6wdVoXO4E7fmnMMyMmf9x4V0SL9+6S
9yTWTw6wAvCJ7/4ol98PEa0onS1mstseDMNJo8HSaEIgjMv2538b/GWK7+rSh0i5a6N77BGEwwsR
ZQRLNRKi/kduj2YNR0TuYwuVHlCYaU18o5HaBFYlCdIuxc/kG4rD9pkfbw6kosNed/k3Kh0b19As
ElExMtl3SHD2chDenylQu34xDYXpg7xiLSwaYm7jLANsyi2TXG1pPnLuNNaZRLzFZCxn3vXcqoo9
5L4+fbyjhBhqx/KqukirknibtRuRP355g670BGWhGu5VCJfu57e17IcJc7dt60XzmKZlWiKv350Z
CWzurcXagDJiAac/ZntZxppLZhXfb/jxHm4CM5u1pMs5k0pwYf2sazxLSQBuMyLaxtCTeyMKp+vu
WnqdqmyHbY1TV/hbd6BodwDev0qRVg7dPbbsQg/XsZ5yo/gPL9rq+0VAWTTRu7Fz0YMT9dXt3EZZ
oAWwRSbClH2kiO4Aho+C3zykCcR5s46zwUYiQKycEG9sGmCE+7MFHq/3YvJKz7T3FoZdFCYCPA72
f5eKCgxxQq7iJAykgfA0GbKc1KXgybz0Rotgqq/SLJZvukUwMWzbEaMa82zpsjDIfTmpxPjBCLVI
h+NSbjf1G7Z5ZFurbEt0cm4Ri9UJp90o/chaS5C9aqpdguekDdzfS2TmDkrjcSO3WvWDlvUXd+6Y
39Qoi3gZr2tR+ksUixEC3+hfc8dIH73vRSKB7ganfCD8atNaNaaF2mD7CG5iVUWnM+GAvGp9FJWI
koVh3z3RsfsfhxL1AR1D0lB02fVTFY1qcnR9odHUtooyyrUtVmgg/N1p9PYE6odE9lg4baET00fZ
l1BNWfFPrBL/Xg73CBnBfSCuKmtpXfTY8Oh3W4B+BjUPR0NaCFiGWOQwK+ycOfO4cnOZ5Ct2oCgO
6gw4l53uEwMBc3p4c3FRQYHf52ljJDxkaMuHLwmVrL7bANy8V5p45+KzFdExspPCqPFp4gFsFekQ
drra1UHMgjngMo3XAuVFTjvIzx8HaRHXVkVftst3/j++tSGaeoqnu8ZFlOtSJM40/1Ze92jri5QQ
ExHdgfxrRcwGpp2o3Y9zWe935xCOwrGl4QkohLNDSH2FUvVZCf1B0Q0fQQAuunEUzUT1Y5Tu23I2
DXxk075PJtJjZZyfvVG3UyqAP8u2jzQ9R7v5mA6ocgE0Oq+fnxSA/obGaE0Oi2MGxd+DeQ/3VJIH
c2gvW9A8uSTSVRKDK1+KLA5BGAPA65CpEzM354I242eB1JXRhAke1pTCOcnc2zlpeyMTifVfS+6R
Xv1ZeGqeMzGzmkqMxwthZg1GiAfEwIKtg/ypNbZxjpq/TKXDLatAGBfok0fVkL1VALbgtyiMXBkA
A9/N4S7fUV0zJHJMxOcL+uBOvctcuuKFcfRLLYmq0Nvhs2I513o2tCPQpG1iSiv8ywyXjg8Y1IDb
Moi5mBpYhX9xcCoiIrEArxJ77jNXbnr+Ddfwm73Sjv8OMBQl4YBojqhbygtZlXtOPxDvp+DayARv
CwF0rwn43xwHDWi/6Ud5y8Cz33NoBEm8RsdLsDWGKtvE4bc/75/0E8HSlz+wm+U9/nuDxlRCM2rF
cl/RnBqPdfbg0HXV/pCge0OWY7+ADh+lVhmj/0Bq/JdaD1Rd6uoHF80eRZsANgIWeMYvsiAauGcY
PuNL25ZDnBtABiATQvo3YkqLyeO0JglR4KKGHftDnKg2y5G3iwM4GZsKMZ/v5QU/UD62KbsTBWhy
EzSmdKukSrlEUgzH87nyPz2JvJcw/3Kz1E845lCR4U47fkcUB+BPvRR5380fZAaVtGzY4jq3Fplb
1HzNTq1ObvZ3LDxuIZpYxBv58pTMNGuEAU9/oOtUcsx5ogOJ7yVUlKpROoxTAUnjG5DG34E9JAqt
aN9jZKHm8/J4M8ZdeqVOYsMsJG6HpjxGAv8ZQei/Q120Swmq5kQBdwJiIfHJKE3AlpG/I3fQB9IC
Ai/adZ3bytRUUXuWaYwAu9sdb6OG+fDp3i2y4K3qxXbBGqJh1mPVasuPvNvfzAH8ktSaObg+a4/3
Krqjdd/x1DMVL1l7BlgETR6I0tA5gXVlid1yaihRMCUH/TapuNgEm37LiFm3jShKkzp81QC4wPpK
ps1sp7nbNTx/DCEFr0vZyh4wkpUD+l6h7pMS5sc3zuewo3ameHonLdzBWLe8SbhtcCtHrIpWDgaT
Sc4ih4DqxIc1FlTgx5jeJuWXWUWqgZUJBdrXqHTdTmIUhVZk0E1pf7//MO0ATopqFX9yyGC/jcg+
/Uire2MFKlMZDxPCmsRFzyf4gLkRf3mAHwdN7+mEViWgjeTYF9G7EHmUbzzy/9y5svqmnQTg+dgP
ksoUAD3c/0MB7rTQgqCjz8Zka4CT2dbga5aZ75lBQBRlTa3m62G/GOvthIgdmapXA/nKBaeaT0xq
VNaHTxrg3iJwWP4Rbt9mbTiNARtiaVofzyiqGBfSyLAI4iroRBo4aiOhbREETxA/fcOGeqR0QYKS
m58eaEjCxdzkaaG/K7NHX0bUzT4C5SfkdZ/4Zq5AMkElJ5UZq6+H3KvJWNkj8I7woWKZ9Z6UVKuW
mgMMzs5sGI10aj6mgw4u5dXCNiUhqvHegkZAc6uw4BLxCS1bQNU2Gs4kzaW9v/Fa7gMIFhK/CNCc
wuTyWPCbCQUG2dRt0FVwkj+0kvHw0kkXHsxd7IZCJtRbB0kBb3fg0WDlC2hWb/duOaIOTluwH3lG
XnOr6XyxprlRWqAAmPLMI3wIAdCRKejnJyHVaX69rHmii+TDrcf8goZnaVGwM9QF+y/2513lfyl/
uCFLM0JZwowJjaKpADFZwzIaVlPcDwS8o1hcjCFUEV5ayXI6RExdDXyQAT5bj/vNTT8A1IhAHYoT
2xOcyVI9ZLBRFyHEg+Y4IxFyX58PtZHqPeXI3lMc5cJOzZe850k0xjqikh+rOkA+hP/hQ05APQcd
xvl3pLVKt9dl23ySJuax0Z9P8A2+b4/WaaeQSBA38Mcv5bgFVCUH3/E6YodqQFO0KK7PZ+2DUO4k
BdP9Z1+eDadY69DuOhGSDdfkWz7vUg0pVVUbhLIgEfquDfK1kpiDLxocN+5z6gxhkS4EnpHH32xH
7hfN3q+H//Yvzk9mybQ9MexhBQSFBOnIsDErapxlavbB7/2QNV8brkxsi9Sk1mNx3Z3ad9xj645M
kLK63s79N41clEwBr7q9l7dKCZoNzcDJjL8yC43BhhDBLd3RTUAyF1boLG676IKp7k4pzq+cHTE5
3f6XIko7FJsrsSQ4pmICwqnEQGh1cURBHjdkPQiS33SuM2gZ0TFTaQqwMsFv4MJvTCdJ5Jvg7WbL
l5Vce9VR9rsTSIQVSt1kQoGLxNY+oFJGXpeNuLjrhYh0Nju4IKprnOHD6mn/ILpzEvZ1BTYTZto2
UwrzT1DUIzMiP9PbEgp8JDsWllJOnMfdMxCZarzqQPqJ8TqL0a84ozgUYyy/cBNQAZJmF54kumqL
gxZoacK35Ic03HbX2IrgLtUPhOTebhZuWCQByBIAtSoP/zjK+gilJpisT2FjEmvfmK3PDn5mGEti
NKLpGoVMjldISVxnu1eEDu+PPoKbwN/MaNpBDyzsGBqH+eDwGb4/ee0+uwRqSRvvO7SOnlfC3DF8
D3gt+6bHLmrVlnMSfqfTg/Ql2LuT0QpC4F8KgQhWJEFVPLRpU7jWVBvlU3fpx5npa8MtA68zaXT3
e4EMSi6Y4dUOkR5Jtnl7CWi5rdWtxOKoGlc37P4nCCgLwSN+a0g/UaGN1UncXbfRge61Ldw5f7CZ
6VzrDwCUesqGIPaDpy4U2Vq592tjNO/2bHKw/PphhJiYiB6GwSllvrn7JItG9GyEAxhB8to8XmlV
Ich4DhXwV/12bH4q7LohoMGzQGMEnToXU7K9qI2NtWKTOax51PmSnCPMeWMf1SnQzDFLKRzT8rDy
b/4LsADwiCHEm3zLoy2I8swe7TQ1GZbvJsj3in0xYZZxmAkKbJ0H/Pm2GUVNI4KNXFoivrmFkEQt
vHfkiutz3A/XkZDQ3NhzSskBEFFIy41g053yhZKhLTJPOYXwi9K21ACXZJzsO/EGIr3FerKVvAlk
FtE16zzFwnBcV9YizVH5cNowKZbPK0tF2y6wZ2rn7tyOWHbYPE+aX0Jo4rnizdqVCs0EAibk9GHO
IX6aVLnooqmTVrYssntmeW2dWcyfT9ny7GqniDK9HGlR1gHKKgq4xZbQV/vSO0xxGe4BjBSwYseF
HL844eAHwBhj8R57QXo7sbGQxJtMFj87SVQXlqin7mM8U2a/T2rn9hCjoRCVw/puZhezUtccOeQ3
H6kuzG2vR9+B29a5dcRwPR08LC2+Ty27F5W+Fuee2R4Rgh6z4hNDw9DhrgRpZivYVv9qupMpX71H
3hGQJm+RCFp2uRmdxy5k5DAsQQh3TzoCyDGgdrodm2q3yjiyLea7qRzJn0JgN72masDRRcrOyYXh
im2z0j1V7/jdwsdg3SGWhHP5oAbTSwFgMA14xTSNcOtI53C/HDR0YY5iZd/knsLQZyzWf6h64Pem
6uaXazCHtlVvPT02yi3Ciu+IQG5083iAh2veIWqKTSIijJ1QNFiaOHrnItE0ggegdqWD9UTzKR2q
mYxpCoysOTFmKoJym8uqlz+E4Vy82veof+WRicExtuBEQQMOMr1+zzQZoeoOAHXdfW/M54x1w11Y
WAwuVlOl+N+XIiDfGO946KH730970e7AhJZx+ZvOe3IrFBFwYbOZvSMUfRYr/4m99KUMlKKweQmS
dlAMekt00WErk0s4qNXLDd1MqpHpwSroxE4QpZmBRi85nHiCmaOxjyFr4y8RJzqhNsSsQcQOTjry
+JE3Bn+SHuIUTzHqxSW0JOmtpCQsV6bH/+0F+7b9dPxbnIBPSecwdGjv97UMKijUVnDwpVW6CCnZ
Qei2Il5/wshWu4ptstALkKu734f54jSDA49VFJGP2Trc3z8unmvMmFCrfcnget/kfOOTR99CDjqN
oR4uD/m8CkwixLNSmmLW6B7gPzma3B8L/06Y6KAIpiGx7VPDiK+Wthi5x83x2/iOwmcY5lGgzXwD
p9GTRmj/zSIryhDtI+SGJIgoAfFwVtKQZC2r3lKJS3xvpsFPpWX242RYLBEE6anjH2CLpq9TsyzH
YVdfFZnG90deaYPt9xTVH/k/l/b6bWGYC5gZhBYLNi0IG7pZumFmGccSbM6eKLjih0RzHCL3Vua/
uTx+w9bi0t7PDxNAk6achx3HdSCZbRO/oM8xQUK1kBEY/35qV1WWHoyaS198bXlaINGymx6pl6Yv
0C/vLQ6CuVJOMSGpe3lo5SylG7VPFzAB7JeIXT8GmPkMBvtjrLOgQIkfH6CcOBTgFTfsx8zLghkU
LGlVIagi78az2DenUF6Haiu04RhMU4GoiHoql9z0iSa9rYYSVbicI2zmnhGeV7KPXdzucgEnsipF
VnhtvokMbRbCap1idwPS4fSwGAzECtiFJF4pH+NiztgXiw+usGHlLQDtqsaG/ITIloShcNcy931/
K+uO99lHubGw6UjmZhJ3Wv/k7R7aBFCGT/O/PUSEBSaP54hkfog9hhT9KpO64OmaMAE49L8Enaxq
y5Qx+HrccqvmQc6llBdRgP+ewpYohyOLqKC4fAhJCEQi33okX2zBdx/IkKgK31Xhv75CIx+3outx
uoFoSDAHaKLxlIb06XIVpdiCMg6/D6qWmGh81p7WS2Rs6dqubWxCFpWOzLEyfflEDonFepwtzaIq
9ETGD3hJc1Sb2KQ0Q1H6B8MhE9Ycm+6kN4Gfqy783MWhp0ygxhL2XCi6v/8ii94hNjz6Jl26VgxI
HlbCz1MJSn3Vd3qufEEIPAAelr8hSQzreAgidYG9hP7Xb77ERJGhfV/gJPet7weg99uwUDlkWgvc
/TyGqjfYvP6o6UoHvD9QXD1uCp0GhKKj8n8rebBBe5+GaoU0+eHSLW+8I23hvbSvzxFO7+4kJkV0
VbRGDVjwsEvHY4QQGlFU8VnIBhm+Ggfd2whx+7YfPSsZPcmIHICb97h75wafAL2BRjMRUOkj2+HV
EMnMNLkI6Gk+GSdVqvpdGEcA1NIQdGsIqARWozZlNQvv6W+ZrOH98g54QoB3iwo/NbqZ1e8Wpn6O
HFMikz2naFe9riIt2Lio0hNxvXCE8qmYIHGWwD4bOQk65jjiNkL3qUMqB26TJmf1g/1tBLCDCvD9
ZA8p6c6+SwQP2DOhANRglVw3Jgf0VvUaaNV/2hyVKnln4g6eTYtyNPszznN3PMFD3gZcFX+VBdYQ
mMbTfKrOMIL++T/aRR+hH7IF7uxboYkD0yo/8cc0lAfPtE8BvcaqFb0YHs/2OhgEb3UvZ8lv5zCN
xquGTAb/dV5pYkjFN/EoB6VAqnz+gkcpD2Xpxt2IPyBXZQ3AYaps52I3SMjV1fWgVL5Hu2eP5Vse
w8GUoKpGQx/RRG/fcSWVQSxFUvnG5nYvvyPQ1eMkkfJu5hpjz3+sAQCeWlh+RpPwD+A6jedki3cu
X85TYDGNgxWcREFr6p1kEw3KV1ZrPqqakqwj3LFtl2mCabyapUinDclXxNNwrG3Mhykqp2wwjNPo
cvIqaJU0XKOUd3cx9r3YZWwEk8aOfHxo+Grr9yVLh0lMIwY4H06TzQchfxC21bB+ELunv2bknYUZ
KBHQnUmcgW7fLzWHjdHK5sw4AUEPBDeXCBAxLT38hCdwAyfX0SxuTocD3XBxOKbbPlJC9TwMae+a
MDhzsUfpW5KZCOoCG+IynP2gDLSg2lKw9s31sT2+RaVoXvHueUvC8XZU+UENjBrmsmZ3WkbsfuxA
GvYWYyE6hDTZXtdDCw3lq2HO5vElawrzq5QdpXeEha6AtWEy6wjlJ9SWXO1Q0ISTtCa8zi2YfcH/
GIfnQLH1MPjYC94/ivRJsN6POt7MAOBCkKAoLDV6x9rN/8BMBJKkUSGAsj9VQxEyX3Se0CpO2xeH
TFCMRZR5tps/QxJHD30PrlYUQp/YwiVa7m2RHgEPYtuEhystTL/4iy8jyJT2XS0MeHnygXH1/xsz
RqoXUYjtuYNRbVskvlPJbt/275gWflDLaUYNf9/69I1u7G2+p+wII8rXtKAmnpRofK/qnl8yCD0o
XZLajjWVGDtnNqrAA2w0ZBvAx3ycS8HA9XZDzKJ635jDnCli1KAVFWz0mFU6vjo/8rR+/7L0X4el
EjFvDa8tCP+jU3hlgW4J82Hu2eTqdB6TirpruI4jD51IQhGP9l5u3fqzNnsp89yiYZhM46jkojRw
8tyuF1TRE0/oEUG+b/mwKyiGLoPsbDo+1ht7B1wN6bfESkXKO70kdJfI8WlMLB2pjDO1GQqg0ep8
Xnmjd3tbTsCaMdicqiQar4w0Nj2T8QT5UWnLDmSB6eGHD5RhtK7kA4oKxr3iQPvT1YYrJfQAwxWt
qkwcW54nV1h6RzV6dC+YFJYBYnaT8ud1gb9X85KlTbh/3X4mk7ei4zm0xR95d4jBivZGNoNEw9T6
qZLVGsd65H7PnymPVD3VvDbPLO4HgDvre35b0tUn6ahJxCD89ObRTqvDpzyuYKJd6Yggj4+7hFLQ
UEbd5MbqDEnmCNqppSbQOzAP0Gi6C7yNGwSo72FDuUrBP1SCCwsyUTjS5jBym0CbA0db5XuTOi5h
vUj/rWBp0xZwT1Cto5Jlg4KaLr9z1QtSntyAoIke8cq0R5Ktnd19Etqd560EaTD2DjTyY7vUcshN
gT6lnRdxmVY6gvIsZCUzzgoaQmHZYW2/vF7z2axceQK/0WsT1nQoS42JAdfbR9SxyiL8RTkiHgaS
HPQ1yqLhwtMS4G/P+iowNy2B4GUmKhMgeD1pjxgRwnJqz63Xh/1seR3kdYgRcucBiUSpxEVF9HV0
q/NaI5cdGkfrfUD1oly8QnukrhnCrZQF7SqhR1lykPy4M3mnD9srHMR7194n2noQ0j2oeFoZ3ITq
58kluemBn4rlP8twp03iLHgmvI0pL+9rOKM0xuYmSUO7jlakDKuhHwDkcCgC9u4ntHo1WtdL6Cge
nGte24AoVLOgn7vibfi9Pg9Tvd/uS4ynZpiMPmUyXBg5xcwmaVTKLi2ejsLvH7XajZspJtEypMD3
MUYHyj5rG9RFvTaC/VLOLQRXGKpCYmCChTkwg/V5IVqaC8DuCaJD0OU1OkCUwG1wiyg3b7MiXKoS
2yAXAGXGK5Wj4T86ZAH9xOY5NRbF+8bHy0NCEYnY5YGoxsWFqalhc3DGESlE3oeQY9ndAYtd+oyx
bdoNCw/93P0fCM/iS3PltZjNxmtK6dH8fYeG2sEY7U6acREQFp15Rv9N+lpAjdBD/X6fk8Om2gcH
HOKTJghG1wfXmUktUtGQlAjCaE0ZS2LlDVTyXKal+DWp3QxbiH9010k+YL5mDKHQ2B+2pvdzPO9R
2r5cRwCqOe45k0O85iTiGniw5Zv6G4dvo81rqm4oxfHLA9jyJxHeWSTtjI2wkVeKuKwNqzHecZUl
yY04SjYtsvXjGEJ6URwIprqpHFG/RgUmH2VAC7us0TzvHGYaGBk3iZZ59nPlIx/eK3SFz7aF0+Ep
1jd/SQrnwwOsjuHJo48UGm6GwxZgYhCyqrxDptatoq3iku4UmZ4w5K3GYOKViRrQbkmWEjsz0fmt
oPwn/hWP/u2n05FCLwVv0E65Hwcg7uteLETjKvGG2HXzYjBNSe+dO+c87lYx3aEwg7t9ylZVpFze
mqf5y0MjOliPaYOYQ4OvnTiGW9nmjEBYGzjy0x2rLPBgbwDWK4wajduLRmuNI32hePK7bJe8X4uZ
fcssyHlqd4P4xaY4JXObBjBVKRCGeANtmPhNmKY1LTA8Z3w+kwj3I28ivWUkz3ZCN4xwSiTIuiu0
JZBAJB0rsz8Urjq8sZ5gMFUNHyGu8R+OBsZTIs+fp1zGm6W2/D2nWYegi1TP8OWFjEBCwDxBeLBn
B7WkQEiGfSRdkrlbUUF3muWzXM/kVggEzlhD3WqKH2kYRB7xeJ/IBLg31n9KeVJGGFtJc/LIlMob
D+BBMjHYKxaa9M4lJj2w0HxUhx6szS16RuQKaQlSi/xNU89WyZvrZaZKMee9Ade5XYLuZQhf9p52
QjpMdCAHWXkVtzFM//oTZ3sWOdgwXVjlNZ/Tnl2fkjWlsG83U1SiXkDdWT1vMHSZJ+0dOIbzKUFG
jBKVAjT2vlgOuEghTD/S9h9H/E3f5LSO5z0WU+DzRaEIhrJJyZDobPXhvOStLq9WAgFAc13TQnHs
vRus3eNRR4EVrgPwEAi9UUNjfpnA1qNUFVeg4LtUQA79lArGQn9qlkTWRKgaHWElxHjF3GFHQbh7
12nPPJcqVddDNzPc8B6sU/8/GcAM42qY7tlGOE0uFGCpaALHea8YtO9U1/GgjbvTQdSNyK4m0Twn
s0nr9a+JDb3/Hs/49qKmPtM5JGhmDUbK4rfrkPGCjdasKRxE4qWFYXB8AXa0RLAykNLW1KGeu8pf
iV2zrCnZflkbCmhe5EBD5AWnD0pp66963pm6hbW6spjkjM/AQ+XdbvbMoJvximTfMb13RVLk7WKy
9hME2kTxxcH9D1FUoj98JvV012/QyZWN5rlBcUyoz1Zm/E/oy2KiziJxBSap/b0mAXuVnrASOrx9
Xf5ImUb2/36EyVfiv2q41tNNOB/7xTFDHTzC3TdnJaghVupRtfndRu5U3fjEHHt3IYRKdKwtDqxM
qRmlbIQuG2pZI+7SYOdzXpM1o7prCNh06wBiy09RFqbnXMQ3aj1PcIo+GRAlYud35mTiBhTktZp2
758k0SkgJv2b4O6xDaL2oUcUUse+wAx+pDWDP8ektVbgWK4VMPdnu/hidsixIxAUXGMoXAHuftPh
vfEzFk8vphylBAauvFI9NGcfrUpVbXrQaymwsAHuqrbPTCfhlciE/3EGwpTH0xD+jpWogVPw4U0A
GjbyFIekcqUOP47NWkOeUec5LV3V5Gol5a+VqwclNJkga86OC3oPjauYpFyfcQ6iwX2idhSs7hLL
iqmB0vjwmzJAQxuRCtt1jcZO4nuyKRrEjeiy+uZHv1HyvJ+AfUF8atPmUsvC6cmPo+aFi6jxL7rs
XrgrGxd0dY37Qui1dn78IIkfvCaMT+sC6DeavwWHJD18gtyhmM3Yc20X1shp00WiEuQJoonePOjq
nR6drRYb8GsR7KcKVICwEU1eKPApNWxL0UfATUNw0jnfaz+kXhC9YLWKJRoodW6gLus3Hh6Q8IT1
Kpq70MvHKDadzvRHl/A9DEx9a9jZxmli6PBCVJYqyaUyO85P5MGWOYw9uxFEHmmVBNgiCJ3ifYgv
wRt6gyJYZm3N4mUT0KvsQvUZnMSVlSVoDxmDEk0dv3eO5TW1HsV7c9cvFnN+m8KgttYfGpwFllgK
zf3sJuXOXdoKwl26lfBrk7K6NNUp0jH6E5CbwGO5mVHD3OnwebLlgK3Cj3tPDEohmRIW5qPLeD0X
x35e+VrMamx5yUSefjLG0hJ73K7C3MD4sH5bCtOPF1EdWtvImbGT0nXURUghYobw9yjMHc6RhsWG
/qhEF4mKL2ZwaKxPGQYi1JTBD4dNKsH+8IDmljbAe7JlfrjJvu/PKJSo18rCE/V0aLDS2wLTpR2x
krMSneFudYV8tdIas7iOb1WLPz/2nRyeN4uVQ+Xb13XfW0Z6wMsM7N5nRDbUOjPQ+L3jPvZOWG8P
amT14UYSuEEJL4UWR0xPAr5bLwhzJ5jQ3kbSrWBmw5q9D5VaQf7J1eRqnuwRj6PDnIrTMG4U2XGt
alGxIaFs2gVBtrzLWIv0cA7hMIbDbX6/BgppRIplNJkEhz0BN7gGEjgSLEfixnRySTcKc6bDhYVB
d/8V+p7IO2w91EmQSJZ++zzPO4zQ5RiGN9x2XGQslIKrWANkcLxYI16COcZVxsWnAqxmWuvt80qe
18n2yFSQU0tL+Grb7serMgn1+TuKAZNN/I1i4PAob/PHRTGKo3DbEkOz9SqJBc0PZ/+iCWI+zE73
eGb67VXyZBVUn2lyBA5DgzUxqG3lVXODUWysFDgQB5S9aDwOymlJ4OBMLAFuu0Z7nlIP8Xz9dZyv
8FGYosmSbPYH2PZAUDnbzVjwrTh1nebSx01vnKIzPbMmbHZYkacTBs8i6diwROXpXYY1NmD0BWlX
4OPLiwjmI4sDOISQmLwPEQxW0FJOgFPmKC2zlvPGS3w9OHDPSQOJ0ggGHj12lv/NH/k8QSovyhR4
wYLyTIXg8b+kS/u0sAtzPg7SgRyevC5YVNGYojD/WtiF5eNB+SUS6pOtgq9tns9eWC5l7m6jPgVU
p9Jx8N/IJLkhY5BkDIcCXCVVYz34YAp6MTYLlll9VzE+cmg956Hp7krIwVNDj3USzTBn9h2xPvqZ
/PMwKc1LwIEzuSJW0sMgUvogdDGH70XN4+kQwQZGXJQ1JDQb1UlqclnQ902BFTTr/ECRTJhOFSrh
92FOu/Pd48cbYTELlTrBeOzwE4wlfIRxeoWfOcHpTwDwosg5LBghZrTk6nKG73sHf7NxvNcCJz35
2QrVu2GU0tbzrYgRAGzFs8Q/T+LK5Hp8np4JnvlF3xGDy0rNDKwNAXpQCjLfgF7JA/2CUw1QwAyE
9JAVTqWImvttmkJhTILbU+OlHWjmgCiWFmKV9jo1px/DjoYEwzPoUbfNK3l3LvQsl+sF/PQy4/W1
CAJeB34gxYPfQq4kXYSffe/4h4l3EvNE4pMXxVRxpLJ300uhqh5bO/nsIXNTh0+yOhH1R0eeOtiw
Yi27WpYcCwC55d5LX6lsuxyhCbHw601ePdHqDKCUVwafW4nfRaWRcaEAIgNOdHbEeI5FEDl6x3PZ
gALasozlxNWKGyNwRfEk0FaYCb/iQNP59NAS8kd1nw89DAR9r6apEIzwseSFNFvWnjZbGITLWJfw
oN3q9JSomohGaqxQqfYh6EXBUcH1QbKvmcuHSzEIsaiBheoqRc/Jcy3/kqNiEXTxbOrQF+N6Sq5i
bTiil7gWy1vU3Df9VjBb42q978vOa6T3QVFZmgKFfrPFiwvo41ddOZhqaRHuVERCnGjW480LeQuY
L5WiXRm7+x8QN08VkgLwZ58CQZMVPkGu/nqhif3dlCY8UZaGxiT9TS996SR+/lfEo5p6yyUxUZhE
/xkdFSqITgigcTOF1w+unZcfManmS+VDEpMCEfU4rDc36iGetgbX++qKUmm+50gYX9uXfvq2zmpX
RcJeqw5+GlGL1ff7DZCAwE67Bj5B8me9Hl8fusLW2kQtC+1TiAkhBN3mfQyxtTdApJXNpIuyer4g
RWIDrTB698NXjNjrgHm7uSS6uG4tLqkrldCZcjehvenk72qdZuPchJMgu+TBstlHF4tOWHf4D6T8
pECf9LTGnQmpcyvhnyYSrEmWDtHJ9hv0R5AKOzVlxl8ZevnANNjXo9+Lx7tAH/uktqEX/8U3ZrUv
urlMGduFr2plZX3YZd06Lc0aSmixmcDPa8uqTjRq+g9+jLQD1TcURzCHxhxoas2saL2woFe4WFnf
yryl/kbLHJnSim1vdwRTcOBB1hnyEHjGHwXwGEERYH8up92NOwveSY8Yyfjr1Tp1DVc+tGUz47lY
uL3Lpiyx/ydyZlCo9q/SEEyPDCE9GiEiQUuZNJzInKpPCYhyjCpCVdaWftqoO313/c3BbCvoIGPU
7/nbXNeqUyDpUQ28mTIkJVYVW1rPP4qF1mpe9jeEEsl1nmcGUztYeY8sqGRJ9cDXwEfqu14QKmuQ
9ybDukLUP292rpBYXXmKGei3wfnVIvtf5gBdAikAExOwpCkicQakbdZ7BSmSG7n8wAG4pch30bKn
9axnTLyDpgLmVrWLtla9v/Jd399g7It4uWvztAPCcg+g+fF3nhuwzwkyLQgHfYF1ZGxPC2GfNu6q
m17OUczGj+jKa70zyceYPN8Rx37Z9VhFojA5coWrBtXojtI4si1pLJmBr3qWiIskpi1jlqhXVQth
P9AbXjRDkvN8866azDQMRec5FGE/OWw0rdswsTW6KHC4dOqzkOM3BZq47ioFSYR2ADJoBzkJrKOU
D75k1Y5ToNrva/s4hqlHzy/6/rrQvGVnxJT4ft+FhwIdiD9DUqSo1Nl5zFFHRQQppolKQyz4bFkw
NxlBNxkPmlDyXBQqvK4EFOh7NOk6jWkPF6MUgAP/6xvP0dycKSzGCzVrzBmWpWi6wQ3Ltdh9AIs7
I26GPQOfvBeCaGKCSU1YhvOs6tY+ssM4pCk7IQFm6n3Q0INVMEmV1ONaxrgvmJ74oLEa2AawqmTj
ILSXgOu8nqcxQJRP2KyB1wqR+Zjl/pv1YJlWCqI+m4ZWZUYfLDXD/i5iiKN4GFYdlOIUSYRfy8Mm
6ZiTEvjWVuDkK/6HT9E6Fy0Q2GdkwSG+oLbiUQSujskla/heraxWnB7LOjkoWgnjIHNQxPQBB4gC
kwgGZw9e34CZTHhkz9PqmN6/CGeABoU9xIzLqq+wzxCHdVjOxHwrjDqXHu7+xKUkoEHEaP73QwQO
CMk7Ov7MkkVZjiNKMpyKWkGBe0b0t8P4hkY0Lf1QTpVnXBBSIwKoyr0+4jdJCv7hUFMlRNHYxg8z
3UmofCA7yN0ic2VzONvVqNCh/WngVHTVEZiIqMxfhffAmA+bHhsAE/gXCuFCiHyor0H19bpcapM6
o/RbNrm0avldtA6rqe0bCMVD1sQsEL6Z0YM0zV6zEmk2oGVBIm1GeLVN9/BVz1RB8an88mH6bh3H
YQvSned6moIMF2tyqSYrih/rBua8TOfyCnDs1cD50F8ibFjeh/ywCZvPVhoOZtURH8PDiIPcAdxk
mApZY41TvaRwQNHD2dnjrJn6zshx/r+BKlyhAi6oT+hEM4c9+lo6sVrtqa08XKGYUW5wMncUCJAV
JmtodWaU/q7dH3uLuo4eT5G4+YS4CuyfbOczMUdcomNwiQsz6lQB9yBoUL/cJ3ADEp9YJs+zJ0YQ
lY2HzttLSvgkuZ2ZB0megmN+P9V9jLM7fxSC8cK3fsetPCy/H+7i/nYinxGW1mdpex3lzqOWpdsh
pd4F21VnwUBRMqx+xtYjXFmZs+qIn9OHi462R2uwphjOkgOzf16hfkaSRU2KKIGAybVYvBQWc80/
/otRS8jjjWa/mhbzxvSd4vdx7uKEc/R8ytq7j4IeIcg6x6xnBZ0NcwrTxixZiT2lG/7te87+MTPc
Esd7KQo6l5v8eI7kY9R7uscS8TtE4fF7C/ix4M6jHcfi8OcsOm+wXqXg+0F4QjTmSS+dshRqFMXT
yyVlE6EKIFhCJo8fBeqtHNsuOEh/mTdcOLIuJFzR3KOabxAI45r2DodQzJgFcsaB61Sp+RGSt+nv
fkVVcWi/13epUjox1RfqADEN5jpNeTR9eOfx/VdeLZoRcJrJsG3aOLFiN4bPQRyNK9yctgZyF9cX
/IkSFR3g8RpykUHIGJJdcNo0fkwMgF4QloYvykD/H9RygqKLQO4+Fs0egifUhiKOhinYouDn5UCE
t0/QeYpajuIfLevK/q26tdnBhr8m3qch1nGuLqQ7T9e4sHsRnKfxUMzShVdCo2+YjxZg083gRW+J
4xCWR9Wl0miL5SRQXrBoGb4wJGdpmFlcVm8XKpuIePT38CWbg2vUIdigs1oQI4P1Lhe8veUlg6Sd
SwCm0aNpKd84TL/DRLizw2bt2mPPtSmGMlvLIaWyx5d7cihMZ5o/VVG0znWxzWE86RLx9tIrjt+i
7qCEFSZCGO5KAqaLu+Bo/AmRTXc7TgjJwF/MwYnXE38tZ1xxxwX7xGVyM8URe7pMIcRthQcuKlfQ
imEl62yoyC19/oMoV7rTn8PYhhTDR/Th428vmQ0BxERh5b59ahYvf/tvBXCOJUejE902aR440yX7
xUvCO7MGjHYlSVa47Gg82LxYDuaQW2akyQgPcptvT6uNmA3ExK2yebXhiI/iMNS1U+CwvpG7BfQY
JurGGaNiiFgKVnkSyOWpGFoENq6ee/PUwJ5pdjh+B0s38SiA3JPZisck/NzJXb3nrWtvKVPRfJbs
JHoqzGtZCJeiVPO3+mgW7EINRHlhi3AC16Ky1FZMTJqvvXA123IYl9pPU+hksdEIDE3YKWNWI8eW
MAcAkcBToa6VU7wunYiJDeYpnCMSs+Hmmv4NGpaqeASfvPPE8wdSfV7DzTo5MMgY7NP25fMEVnrp
bmbFlXP1O0II9O8D8uOIfFQb3wIub/yJ3wFMorICKHH9qFXPlbElo6uiHj86NnYr7eJ4DYPCVaBW
yFT29mol2uzxm7BSLNvj4Pu/LtNz34xR4i6rZN9jrMSLyND6ZsJCfztJpC6gYoZAXbl4vpNl1KQT
28lYkay5GQbUDROSknhZF9eVMM8K6aIQMEW1ptlw8eRVxujYgXoqMkfduvWaZmsujw4w2LQXqY2m
NSqQMdJlHv0mo6iljHfBIEXy8bpwx6LVDHVZmjuXK+9sQ/B9Ri8O76Er+9/GGo/rwDz6JJQRcF/4
tdaBQyYwoLfUQxHkJxn2wwx+d4AUhBglxr/ql823xC6Z9CtRdHMs9OzMqlLK2OHj3Oe1s0fOBsFH
W4VO42QQOXHzDxab9vlBn5IrJqlFE5BhDbBhM6v/DEzbAinn6LQs8tRkRXnTQ976eiNvOhOHOsYj
NaJcmkxD8UqEX5OVgBJfGAyFWg1MlAAyzg/whEe0wYif3pNIWaLXL4k+6/Pyd63Nb8bSnl4qHpkz
f6WF0bTLCQX4KeZlEzO/QCrupRXQfS/iaPgNiXIKAqhYMNf16Xcrg/2n/dBahIQLz9fDgI28b2Tu
72qVZpCkAAVJ6/9yXj0XvKHJ9Myul63vpzKkfv6aIz2cBb//kL+CS2Q3VGaV1R9FtR4fkYAVgOzc
bQMa2wuTTxMlygFuOPj0AxAikyfbWS9VHkEhicBYMvb501J8FW5knH0VCm2lUPa/1J4yW/LmiCow
a6EW51m6vNvAPl1MeZd7ggKqSGbVRVviVtpJkL1YieVzyfKZjeFvolFunZiumFtBNvtlFOEz+INb
0BW9SkJz8AL9qooDITd+rRM0TnpVe8jRoQQz24Jo+tNAUdkOrHSxCT9ekDxYm+dlpD5f5RnNNneH
/IbGFSllJPU4tFz/ncsM0W64TVJdorkMjk/TO7mEg8IoVQF0d9lD8Snfrb39j76Jn4ZW1gcIUXl+
i5BXxQiLmuf3lvx/dDPfAkve0dE+T7gmrpuAIXJ/g04/h8d+mH6l52SXcgx7SPm+KAV0G4W28JKj
e90tx/Hc4pOOsgvRp+vGeqWmWgBixcLYrn7D768fP9zHGkcgB+s2WEYm71kh64LvchUUCNhW8VcK
2VOGij6+pubOSIOWaydO1ZTRGMpmuuac2Rhn0PM7glBRMcJugMu/qYzFqOyxkVa8b2a9YQS0Zqoh
jJJPZvZ+9zs1UQYU2YFdwqomBlDAppj6UFFovmyfiEY7MBmaIMmAJW2CVl2UreZileyC0b8G8R5B
b71QNat2SCN++UfXAxFOlCK2+w2/+IXUpIPWeus0nXs8spGqM6okgQebeEVeCCsQxZBIRMmplIIw
h40m0NKQNrwWVusDjv9Rv452LN5lxf1yjyp3K4+HK7XejPwRnX8VVqce8k+9WXj0YtlO/VnQwe5/
1U8OYVSMZ8ZMHaQFqvNR004D+uG4sdYBox/QYqkcKWvFAE76xJeINNZ9wSu0PgPrl3w0mrfQDsFO
AZDxvTCeH9y70w6HOB6Q7XZ4xfouYYIddo0Jqx8ZqgAXMIPT7O36kE/5DxTqs6+b8kEvVY7pEQ9Z
NLxLzvfkqJAIkM9v86QQ4vN5ou/fmD9nm4amxntcz6mwCWf632DtSR+Ub2Z/jkG9Wfc+Q4MgYhdG
nTNwDfyJq7g8q6Xay0VhD6qMskAWrkyZ1Uyq0IUM31rqy0Khi8XoCBuJqhITZFDVjhmSuu1i6PxM
ao3KoY1v9lKxJhDYgWWtNOcHx/vxTuOSF6QJOxZ53qv/Dceo/rYehl33RNIHh1oCmtbetpt14SD6
kurMdGgK9s//93ZlfRJk5S0Rx5rD3+45kPZAj30BAH9iJf6DFvIBjindyjIxYWyopEj4Rck8iT8D
0W4e0NPRUx3i2iADvPkbKV6IDKVCp0mdtp0zP7lXMOtdydI8rnM5n4qibpDcEEv6Ei0GbolYKMZc
Jpvx7emB/vCJTcqWzDSoCgWO6QZXs5yn+22Q07LznddPl2s0uVdcrQ1OdXNd72Hl/hhkDxHgRZRr
r5GeCpCo6Y93JRo511ntcD9YxH054Lm9S1LziW9jtP0fIidiWam0cN3HhBg0JTeQin4dN10aiOEC
+1KMsh1ivBLLNSNnJp1M7eZ0mNVpHTXym0SsOm/joJgG5DIhbeCXCFgsjwSu1I6kHmNW2dW9F/kS
8VmZoXx+19VuFRzY7zF13bUIQ6vD5WWANZUffP50jU946EsytQi4cIT3s4cA7/XUJd4s7Q0vlTGY
IJOe6AQGz39Xi/muwAhE/sjmzYLFnpZmkQZZ0cb7uorsNQIUq4UTQOGQwU/sQWi3UfQo/00U6J79
psvuIs98sWGjqcVvQhmDKJNQKSOQNrnPTSD+NpiuIlC32zek8HeCPlLGOPpUwOPEF/APYPjk/mrJ
1x9CD86PaBqmw9jcmm9RUlp2O6zVWIPzH+3pXWJSi0D920JDH62LepUm9DVGWxqVjjg8zRCvMfS0
GY24fNtCWVfKrs5g1t3EX7+rqXpYmWtFe5IMFIlcZPA3sjI3y9cu7dRWarTN1aenuktzE6CGqTC9
RLt2bzgLSUWJ3C1qwnf8sMhFpqr3TZ+JFt9YsxM8KOE8Vua+DeOTczetMcqNOFnBDGxJGmKIYvbn
3RzO00iv7KhNGNrRg6lwhQWNuWKrQLQTNYp1/785PWPXba5z/HarscIKrofQasuSAnpK8Gd/OFPX
yi61ulkh0F8MonjIUpE6a5BUIhCEyyv6BsCzkzHDFYOmjYv3Q/6ZBeWfML8uZDoIKiEFYEbWvATW
uUcfPdrLlZUa3LIfRBbmCyoXSNc186sBm9SF6Sq5MOJcvZFqLImsTVMqI4PZfZ+aB0+hbzQXwCwx
eDsgNzjSHUcRyr0dS7CidIx5+cXYfpsaiq/0qdSn4A9aPdWbhHz7q+MZfgUvyAtUbKEHjwE3Ta2W
a/ABCMy7P2nsAalYm7oCMMHOdFAs5DD3H/3sjBILP1hj6mTEEeilP8auy5NfFT849pyXIZBACtTO
s3VmamVo3wg5zFRTQIxuv2HExI8p+wxOKjkPdCnUONjt1JjqAHYQDaK/3ZWehkp7OQzrVbpMI0LB
JZFagVQzP2Embjy0Bajoua/rEkPKAvrfPwg2yVx2o1LEzINjuFMsnzdVO6rE+auTZO1vPgnRc44F
Tt2OYHcPjFaUZZG5zSCmrGEehGUBaBG6YKb3Qul19CGZDqTbf6BNz5IawO4Wp9ID0DCpkrrzkhfE
QhwQVoU+CyXBdHGL+Am8cHpTRX33p9eJZpchtxVe6OatUpq6FFroZTIaG+y/oFvpwTBgTpAD9Z8A
hmlU3Xq0SG+GAMcqu/myYij9UYJJHRczW5Zk8eDKozMt+HrV4oG927tgVJq7J6fpjrYRpY2/I02p
c3c4dPdcySi30orGDFNkZOB48NAkn++KdUCwVit1GeDxBsaRnWeVjs3Uhl2YWjCDVDZ9EKlKukyt
TxqvBoGy4CXcq0Wqtfla2ZrUYaUk9JNb/gkx0mVKnbq72O5U0C4eZ372emdGGAf9C5m/P0JMhwsV
AQjkaCFY1wR6MUbYn1XyeUO6e8YrldhFb3fZ5YTsn/NJFln237Psjfn/Tfz0rRmJFRRZsd3apzgX
mjS2bsYR/d1tAGeuNmUTrGbXW+EKSbOM9wH0vTecniRxayaHFC3yW1MYheSmJWHnTwTkjbHlvlRu
A/9g6m3u3XyBjCgQ78zkRJcHzy9TKZI9B0ClTdqPhzWR6LPsn3sdvj91694VY8gWjie22MWyJEmo
8+oHpxA2imLZz6CiF5Uzh7BZZa7JA+DZvQDPbSbpXq1LMV+7UtZVC3g2FO/Y7d1r/Mm8DOoQX8l+
lmZlNZMrBICEpyDDN+h0+INYixp4vLhLwT3qaKfs+BSh+WMqLjsA52oSgmG01CdJdk5r1eGJy7wg
3dxn3irPKlEZyWZteJK8GflIr7fB8vz+8cPrgRdmh/GoV21j78c+ggMsuyUrEpRW4js/ANuUGVCy
VsLSViPWuQANi0KglvWfHZ/4EIgTC7NUojlKhEKSsZYQFWSZNOVp/q8sqoZOSy7/x7WsUbmTsYOS
MJq8fBr+aRh/s9pyCUVdrpUZpuGP5s9cvgQAQtbt38uVNyUdigrtyL7AZAqoiE5qEOIawLzeywhe
r/ivfad6y3l6lAWuzT65EadwsoWYBD8p8lMsbI3nRiaNK6O8ROqiLP74FilyrrLJsPE5sN+18qMT
++Ac1W9ryGPSZyHjP769KNgSL5pTDoGfr7MCYguFFmZuth90q4FZrCrluVGILx+OVc4u7n+07BZi
7BS1/k7pO5AtuK2hRDAuiAJdNuM2iwC6AzZ1zKm069lfJxhhCFNlFdsjazKDgvX3FGQuoyObF9Ic
5sTJNsKL9306gd5gxvSkV4ea/I/bURnja8j4zevh2SZHK5kLeaDIG9+M9u74Vlv0yvowBUWO4uWw
vLhTRzhKCLeI2mTj5zQr90IbnYplTA+R5napZUZFnp9tz070ajG2He14XaApT5QctVwhoTk0Nwug
QKdRJoRUzrtX+HnaDKPxJX9eIklm92gw5xYJCo1kIdDtlOOYFL8zY+6NaRmy68vhjwMqubcCoMqS
P5UsjrpXf4WeLZKDGaFLVrvsuodnPlj5oI64F1p+2ldhhADaLm7T1LLQqWkZcv5LI1sadV9wuIa5
wYhdTa/HtvQrOQ9+smFDLrJcz8qgLX9P2kPbVElrcKrHPo643dNRxgWakMJeFZTtT51p796JXesY
Iz9gOMQDK9rg/AnzdeCAdzhvSzUQ8RB0IWjj2ls52gTm4Nr+QbJkcWxQRIv335JdIkF4z8nAEmCn
ph99OvoGtmDeLQWQtUqUo04gQmcmg5BhRtig6SlD0KYHQhf1A1TNwCJoXJTbOtnHt/rmQfPPm6Zw
nbhaZiecSXvw6A/dx8XotCoIrqeWGGs/6nJLbuUa+RSNPuD9ypkTV92WkX5T7iiq7/jvExB8Gbt9
2JELym0RHbGe7T71U5JGoFE1Th+ytfZte457N9eQ6U7d1YoUY57O5d//MNYFBNHzwFgrBtbLnC/E
7GX1RMa6RcltbeTZXzExQ13ecJxfpyqimTWFj0guJB+Rmpqbm3yd730xUpWnws1RRZemo/zFTac3
0auxmYRkP7sQsyZcjHFAr1YGbflKEh7vAaymX1Qp122QmRE19QId5/Lmk497jVgPyIBrfYIAnjeF
huFpJo87qNv+SxHuM9IOTM/aWNhNiY6PyGHm0USF6hrebg6QO5LbxRcfACZBaecIPMMTXMdhlUZO
up4PjZHt03FtRxra4PaMTOhBIeRFZBHSQ5SgXofwJncim6EnGraOSyAj/uthp5SaaeFSDEcwZ0Mf
vlZkjw4MoUOvSsQ8nkonkauo97bPuzC9X6/f01eqBqLA6yWXK9nfH2qIXk9dE2DToyp1keqHJBWW
LnhC+4aU2SOESfWCKVKTRGdzzjSglM3y7CZD7AaFonBY4UTwfoXBh4tC9uBABKB/IXEXRONynoFQ
Gm8xo5ZOAf63kuedis8erffhJfGmvQ4FTcwqzqz8QRdaI9+rlFc3B0oyHhXnvVTTL1RLmq8pBKP2
WeyrAGn0x3bZbq9rKDecpTk5qhyCB0qmf3yizYy1BaNAWkKTIy3DCd4VDwYWlaYUkYms+qNwCC0r
3TVcQxfnbdcci4Ku+kcRg45DsNYzTfgIEVy5uUUeeN64roOUcEUU3cYpnnXSEFswY9oSj1bqJ6r4
WYUiZ2dWP3XG/f/jeqWw/HNaj/4FKlKrFU42o5eLJydYmHrrW+MPmfBXRaZo3M6DonXgWqS4i1n2
cQLDu8KsmDDQq3DSjihmI5FZG8WDoleUxeHALLOCJqbwVq7HN0KApPazhMHfRBpwZD1oVbL5RbJs
eClUvXk5OxbGDdKGdTN4E6v5PthY6n4S1PnON/tC7TLvDIWr8QsiFnGOtCN3MSa/g6AL+1mYRM8h
w/D9qSHWmmSHu/8w4vRHOxGEVXW6ombAar03InqzNzdxvjf9KZi1A+lsMVbTFe8s38513cnfg2nT
XLpZam8rqVhFiGf1qfb4N+aZXbliwQqmACHEBJAlZGmn0EpH/hEcDAfSQTQi+bx/R/eAaEWr6ycP
O3/SaBaWnAFIuUpEG1NUWJIE2MBumRP30xCj2K+h7fgYRWiZpLr5Sp8VQ7ZE5Cb4/Qs8ZLdXp5A0
nzcNz9PW2Y0vT2mIRqErGSs0Hw9V+4+If2G4CiL7uAekQZKRz9ePkrhR1SMsj+cwiBdL7rIaanTk
Nn7NrbQEI/nQ6/qskRUIU028Ra5iHwwqm6zGyLEbkHRUBTYQcyVyTeCSN+QaoQsnSwm2N5RMDcV4
CIA0ag+R8TajBwtU8i0dK8f/2ytUfsvsv8XgMuU+QkKub9XaGeTkf3gcYWxKjkiXFuxQVj11kLy2
ZR+lP7D13K8ROdF+JLftjuZ7WLWiN4yZtOvH/jUhJC5K1Ct4vClMjG6oJk+Sw6yHIowsR+ieVNHh
Yye651bV1y5gFxuOPM7htKrMMi3ALoQwsUE6N3M0dx4EBi2/q60e3xdvvXGQbYv2uznxBRtOyTzo
hyNb0uXBxUYnVNIve5yW8A3y7liuglsflOpeygCDnPvY2nfSoS05ZLJmhpPGj5Evvz30QUdHiM5o
YDPK9sS/FHkNakP/6lWZHdotEaSJJNu700yRzTiaKE2UY4cVSkB2sFInjKfanQ1FncYwE8ep8U7Y
VYDLhpAU8IPHAJ5M1hrim9fg0yknkxRd89mwW5jr0EXwIz9fJJmVpbbYp6gATv2XWGJSQJXQ2fXP
VBaSnnTKAXbwao4STi6FYQy9DOGrqUbjMzRJUw3mKSvexbNPgSHijqWJrawy2dC1qsFdN3JxZifU
TDFWVhUA6m+OPalSK4bv0mEKRW0AGoqwFEpiditKNa3AeTUIbAAOUGtGZiqiWwdzsYr4XYgGhCWr
kgggi7GYeS+4dIhIu/oRR2yth4JUMJnwSi2z69dj0WEdaTSPGjhfKEf28cbD8nniqBMuV7PEQCw3
AnbiF8XBT1qBIbs7yP8patGXMT5WeY9mLx0MJgdqbKRcFTEIaAPHvcMXDp8Bg5nEILP2qKRQ/EnL
P5N+H/xPhKqAg1DgrbakEya8pWPErOMotMkCwVzBsbUsP83YxWDElmYZ/tajlC4weeiNDlItrTyI
HJw+5i3NgksrPIKqJSNcq4bNUQ0r2fVuaCobXk6Ue9dySzV/PVDaPDDdYBvc8UvvsF0tvFdPRIa/
k90lddgvUefISNeOyzEfCNJSvU1vgAK9TkYGf51b8l/jR+g6hNNVuAv4V0wdSZA3QZdz94hoQRsb
DHNDWa9aeMIpVHPnNghfCyGe1eBtBxyfuFvGOejomrG5PVwbRRlc8K7b19JM1fZXTe2uvaSHYHte
7jGoaa5H0EASWqcMuTGiySiHr5foYEWq/s6PfI5qB7N+JdiHJczbrm/Xif5fMXw9DgFnXNuMiXZu
xdI0Q7FzO408sPUE4HzUp6s6iAp03c0ytrmC3yDUN9H29tCUtIn0YIVoZUTW/91U33eLV2XH+Ath
fLv2PoWCiMrOl1j0hvbrECmSMtiZ1h/7yn6232EQz6uxYR60l6DOcVyfxGyQgUU+9qX0wMxi1afO
68HHNH+iSuuO2FVHegvXgtBGwgssQKyBCv5mCP3D6RzJwJT6VLYKktNdskI0NiWv/5EAgDxTT44u
EjQ2JRFaxiXnq8+IC2kOh1SiRbBNvg3KYkiQqknIVBeLYh6vCdtPTqdbwcAmS7WlGA740iXsbS7C
B9j8dDzk35+eRgWDxH5gaRWy9RkxzbqI+OSNYEEaqRUHrX3lW3YcsjIT5jKadcnap53DZt1jjzt1
oBC4o2wNZkt8PT2J3y6Pz3r+Uxd0r7bMPfy+k4khlcVfbF+KVL4BNB0lPTlZ358BxY7HRqs8WblQ
mg1HQdJy+7h6o8hnI+t+T3y6RUzYZOlls3QpbeMY36d9NVczHqasI/u8tfvzzbQaJzxUGkepGiHj
NK28AcsAO+f8eqfjO2KIgv+Xu+LC7ICP9Vo+S4cI5AW61bV6E7/POQUliQ0+IkZhzIH4asvCDKWO
BPl/MkWcgyZucIx21qslZ0lwjhcfDI0lPPRJzJRWklQvPQGbZfUkjxWyzaODYD47VWLrOl1UECk8
sbTYQZe5nBzDkLb+YnM8d1KTh8aiaZMvRroltqayDbwfxvcKPfgWgyxisQJWC2XP2LVYTINckYCz
uqomX1VmEoFy0UXw0tnSKKvi80lrrEuMFprCX38hglsJSiDA0yhcvkBtihMrObuqDlUrCqXCI9wl
cnNHhtdvC+bNdpg5udM6Z617lXmwXGwjWQGk5pDWU529lYwxrrVGfPIXA7iXs4pN3heBwYXbOvrF
EVT/2vzoYIdNPTeoLGu7/1w427maWC6Aaon6AyYukPNza+aQeaP/iao/pLibfbP/lfyaQVU/f0Ew
hjd4yGGaN1i8eS25hriLscmzRLI95qH3haFI5oUBKt29yMLwNQTBgb1fpQ3s+b8n0s2D/iq5QCXy
KrebFabdPD/oOGMZaSBprS10HErtNaA8xI9UkphS5lMP0m6ZWzGP7gD+gzlUBG2ExpINkHRxDEwL
YV3XsiPLnxqttD/QbnJXJlhTvjVzQHf0LLDb3FXSsoDMEOXz/92/hQt/PxR8ej839iy1gyRuJjDj
Adr8BZ+idqXbNDAdoTArYnQrvCsgkVarks1dzodQg91tpdTL3Tv8VE3yDcbV+TpqFP/NTGRxZhV8
kh/ksb/rrNXMAAU1fuS1yDA6VRLCVy7lcclu6//2v3LCsXgGIFPaC8GyvVnDS3UUpxH/NU/7HfPN
s88fJOvVEV36hyrURhvb2+xwW7xnAJh6TzGlAxuJLGiLprHous4yTnUVISGZfsVcDXvAPu6keihv
JgdTrdpFm74y8UPAy+7VEYP/0DiJ/CXx1Lgrax7wcWDMGs1lE6lZDNB+BQdYQSZDTqX7BxaBX/mn
Jy85fXsL9Nz2lrzrd4ts6PFSMY1PfSYCOCcQUFWUSP7S/ra1m2IzVAru4mhRnDUox/3iNTNk66Q0
FjdEAroOELeVHIfBoxlDhmt6Wm0BfC1ZhkDBAYp/0TP0OZe1aVBJntyye2V6DH5ePs1TCM11bheK
l6sve8ANoS5x+26wqcz3gNbwd+1koGWAZtNkEPa/Rcr/4v8PNvUECcARQwHvusNjMCdqos5jsv4m
Gx/ti8WUeWXe6p5VrDqiHSXPdN7pw6bXBuxf5fYm/jF7fl33DRaqSXgeFGyY62qhTt1XIqgDkCyU
TWTKbOWXnvYUR0IVsKgv/Adab8xxkx+Q9icb0L1UQzWtAfNOhAp1Fxdzx1itnuOQ+LiAZR+G0U7Z
4DSivOsHsHP7r6ASjw1M04Kt9309Tt6haF6tlHHbeJG6/yNh/D+pwJvh0XPTmk1S4rUaxoeuodx2
ENfIjsZeFjY679pn0KnCJSsnmecLMwQAu8gO8jr3x3zGigi3oj8voOs29xHQinJVmjYnN3hpNKFn
9iNCthjlk//1EwNRyBJw1IwLMBWVdB6jvP5gFzkmh0Sl6JWgH8wfLCEey7rTP0Cecejcd/sKPzXo
jD7CJitxzWsOdy6FrBYQIL1xoqYUKGv+SrIFG2x/dbxoqGVfnBALhdsh/gNVfc3wgHbr1zgENqMe
4TsEt8RHW2vM0i0JtAXYV3AAD/moW2U5DN/BvUJE2Ccqg0UGnI0WfZm1KF2W3sYi6BSvDo/3kGzs
QcD+joheeZUmGwOPojCeh3NShYkm3tl90G1tEaFbEUALfTqymRjdgjNiEQwGaAtzakrpsehfnAuj
Ln4DP8TTxQ5k+xZdN3Lwmkic4ckovufZ4Bwn59xpxGgnEamJLWeL3eVDT05+ivZH71jP6vAcKlQ5
0ULhrQfUI3V9M4jHcqRnGmgpUPAiRZFmYjopeBovNBcVVdMcY+DMOHJeOsq7Sh9X4yiQiwHPusXd
oYhcbvZkH5yDUITmIVNKwep+UeoNV2/zh/hIDRNW533AJB0mt0bcGvKqTmYQdHJ+CzSsc5nARMuC
48/rZzKVOs1w7CtVN+2fbnL0eAGY1hT4302WPd62RkpfKWFQQrGns40KMdrFmfXfY0SDAUHTo7ls
sc6sZmfGiGqjq8ZOVA5pQ0rmBbJGDqbs06G0kDPOnHo/EFyi1yl80lzQ4ccgAib4KQIgfgD896Zt
TtO8KW0fy2tbtkeAqagY3dKX3ZdKRCr6A9JLTyKrpc4HnuI6Qy1JJKXkALiKWyqrgRCSCY+AlZLL
PbiXg2c0balewfiwCQZNqSePa0CdZeH1YwzxnOSeNu57y1P4SRLmBSqvSPOx61hNPfjYgDy5HYWh
XeT95bQRagJ0a8joNBxEFLFXXLF5auxoh9DBJ9bBQ74EsMWv6zbEri7XDAfw0HtiTaXuwdT0TGKE
hb5dC/dirEXBY2XrXOjDILX6ZzU9uxvKpLkjNuXdBJXdiMaYFyCVAMTICqheY4Fxc3FinNTalKCm
I8q1WPP0ASr7seK1/LWpTzOMjObVYCCT3RPOuMUR/iNGUGeFWKa7TexWJn97CNkemlGyhvF1vU8H
5Vd0ABr6Hhqha5lXDEPI7W5IG1Ll9xUkatpifs+4OmF+5fFGKbqVgOBCKP4KWNYco3nkEACKr3Lq
ynkL8q/NiFZJYjv2t212Df9jBVAnsnLyICikZ/b7PYtIOmZiR6Egf7FBmGgCXWqMYxKN2nSAqoqj
gqp3Q2URazKWL7kASUKI6x7DrUfCAJz/qigpCB+YS+kGiK3xh0eKW3RHzTfkgn6IF8AVYnU/bCgH
LnodwXaickg5X65NedcmAZ4dy2p6Cd8gK1WqP2ClwiEXHklFFA7AfVNnx5x5Kizbd+TkKwNQUj15
H6LtZ5PesTLy4yz6ZITrTzPPx0E2ZtoJ9qxn7J5eUjew8yc+FS6eGSlEgj1pYKo6LMjpVw6UrTrN
dthR9+amZITehKl/eTNgEzC00/MI8Gc3wxlSZS+U9dRU+xuHCz6wREagxDRiM/VmWVUJA1D8UHb6
gO8OoRoh9+JQBvw/69iW0B2HidYlj/u4yfMQz6qwRmwP3dHICGR930xth6IVgXzWrEpfefbcZLem
BOMASTCLZwlYNON+PLk2yft8qIpsISUQz3wxO0sJFuFffmL/lOLF23cASS7GyuUzwnbVPfY0dZGO
EnMtwgSDT8/KwCQzMNaUzgl2mQzXxpaqoedPGfQUAViTG//Kjty0w0esHG3pD5Cd8hy3snuh+k2I
OQxbZPv3ceVKIHsru4n0FTuNy6u3IN9XfDwZSenj0ZBvp9Lj3nue4USE+iKd3Qlkl93t6K2M4kQ3
wdFJNzqnDL094GmaE3v9P9MvKGyA/VHv7iqpWjCI3QB6Ymr/dvT5lctZxglJqqIjirgDaPX7Z/g3
93RAfYeZes3NuOCYjETZagKbJOnY8Atcq7alomH6KY+/KDWJgs9zW0wo+g/fFEb5jUqAkPm8Qfnr
Gw51a15Rg+J9qUbsQ5Xbtka6N0k5ZckuAgPTmLbmA6/6cwVkNGVpt6K/LtDZw02WarJu5WixgnFe
Sj7l4kowLqsi9FvETVEIuH02jH2qKM0zzhf7ligIkEqa8XVdWto8bUoqPGFux7iYny51E1G3KfwT
gi2myK0oyVYcMIiXtv+n3eIhIzxVWpwEjcHyZ9+aYnAesyuedL8ziaMW3ThH9qndbl4Bozr6g24O
cRQukGtrmoiIvL4p1SBlXZwAsJfFBo00RCHn/C9zQ5pPYbOe+yWIQSJKmiCVETzncUH42QdpLbSh
/W/X2OZj5d+UVPumQcDr2WJgp42kkrw2CP6yK0BGyoRPDnWxlJJB/qfPbPh0z6a3ymCMgywdffEe
d7kCWxHtAs4FnpT8o/fbvH0l8vTNW7XfHSzYxNEl0lnG8TAQKaTTjdMQjhkoZOmAsZDBX/uvTJ1/
4YBJKnWm5y+iuyLnuZhqo7vgu9mOzwxtfiSRxVEyXeWHM4tXcz1zoFiN/YEiNXoV+FQ+sojFL97O
oo7XykmosjcQzILsmVFmEEZ0Fb6DpkXLa206/KHTkBv0+u+TDo/oM6vCfgVhHWx5cujmGJadKicb
jqW0aTa3cgJ0hGDF6Y/GXVXNtWl1H7b3o1+b0uzH+fhYct4idwO2CEVVjQcYT/MLojGbPQ3iHoQU
siiAvgW5AKHbPYJ8eDoN5lb6lJNXmCe4zxnYhVVKvZYLfl5o1NYks8tzN7+wRSq6pBGXoqbRRxxu
HT8xGftaT6Uod0HsXZaAU5Cy21o3bl5gOQpIN2JNOcNWoHJX4N1aQ1K0PrKmduScuv27pOC1A+zX
CiP9oiTyxGAfHeNPigdpMv+WOLJIKXh6R3FDO9Q+17O+l3y4p2WROvWTbKWyFVx6iiPrwQd8Fpsf
VLfPa29JQR2/D1kXUtiCg0CKYGsB2DavBN+15IfRGH8rx4SyDOOegGh6xuw+C82XdDL4hN3IMjoj
ojyL7j6hGfYUrepyBR9YyUZpYi9559LWGCbsOVofucHTD61ZxeK5F8ivVXkoOqq8fLAzR6DyAWd8
JpwWhTBGHjDil5PB9nzUauE/PCgxRt4r+43bgFRgGxHAw3xh8oDIOpPBWBfxh0xMROONmbmTmpMZ
7ihMe/QD3oCjw+7SSE4vXFMePh4sofUsTK34k6mbtJF0qatpk4O+l/5WkDsyu7dfvCGqMmjvmKNS
fJTveVFz0ZHp41LwLlRZ7nfy56VOKqoKFJCLlvQuKWcr741/onTnmcdwTwt6Enzff77y25d3qne+
D0dnebcQmHPwfcMqCUHH3frLAZ+mneWIvSypUAvaKNdpWPQALbXaMjgF5ynUzBtJgHA9cu9S/SSN
1PhUSZMaNglmW2YEi6vBVnT9Bq653CfvtXJ//m3CI9UeK2YUN4iYP7K5vsjNjqu53AI/+w6UeP4b
+g+srM0MvROi3iAGofgyP1EYQ0yn5UcTvYb4178Vcz0q5p4FVqw1hyfjFCL1QwCf6GlWeeVD2pQ2
CPIBPJbH6tiu6vLvd98NPZs4yzIdPFerZtN1pqUXqZFoJji5Z7hYYUOojV5BGSeXMnNYNnzSjvLF
hsy2p8VF/+TBeKYg0XwKLr65rSSNyEzmcQpR959vdkwaRSFZLdQfymBcWcJHNIQMOXE1dLEoyezM
nMcxIT1ATcduFy7KghYl46aSwJp+SLuxPYZAqj3bTUBJbNNEidipmtaEjpCJo8Zy/FxTYPDL0yHo
wDA0cj8es99GCOVyZoNcekcc36VEODxSgt81ExNVVuuK7gb0oEEjUW8Uoamp+NrDzYoguu9Zdc9o
JdMutF2qLDyp2TZRzniH/zY1ADiOg6jc6NBuUExDQZsQka8m5kzCSN4H9Dw1D51odwWZc325ZyQH
ISYLxNe0aapJ4CQ6u+zDX4Rrrpr0i0IkuDh2Zuy6w2Jq6mamffwLpNpJ22lxfZQlGHpDYRFzhG+1
TaeiOZK3Q53J7Ljn7wgVcq4N77QCn1rggXj6GKQk91HpXx7fHb2uFVEtafCmaqTu3pItTAG+KBrZ
8z7cnR8Wx4iyp4NJ9kS9C2PwcBUnqjRXiQRlHtIWydzTq/BSvK0lYWWB4acnKgjsnJMgYNOT1dOz
x2sFDaGwree2WurCVW3fXDs8NUfZPqKc9sYyp6ayy8wCgtY5SBVc1c0kOeDtziET2ltMjuSUzhbo
ZGAhJ6+cGtt5OJBIl2VIp8lV3ZoXOu7pNnpJ5uWst2CzZ03LYxdvHXD5n9yPEzm3ri9g6Xdoiq17
jz3W6Yq/fXCFqJlsWfHeJm1gvjBcwgfvB6vGF77rqWf/36NrjbqnbCUyyNNRu7olbEg33rt18IvG
4aFSREW/JliYZtHvujejCpWTXPIY9o45D160D/CwS0HlTU54V33IO9+aeru+Sl2mhRA0eYpvabl+
vmAcV3huDMs1ito5aaz4Gg3zD+SMJ8R/pEHmZi6GC5HjkMSJh472Jwr9h+DW3/TUBGVTh2M7eQav
9VUb8o4RxzrpYdSnQLKbEMdND9QHa62B3pkxHxnbcyptbfi3fDUrG8xWlix3HndoHhDhLKBmYRgu
CDVepkn32/SixWm4iZmrdsj4hJWmrn5vqR5RT9jns+Znx0+qvbkMcj3ch96v+RpD2fMtxUnNokev
58rkBOlKKZ2/gWHCMFmgAnQVIPSCwk1a9b89myz3QvMCBuxHca00FkhjatMS2VQ/aQ07kuOhxKOg
nVBgoM2i3Od9rIXZi5QqnVj/DzJ7ny0ttL+DC381n/sDG1zwaCLh5oG9dNgDNvtnXdFc+GNvV1rR
ATFKwF2TdpqW1BrLy7iyarU3ZAK9DzH2QbsEWUEVOFuMBkNx0ogpz4mHCvoKzyLjySiU4PLamUxB
M+DkkRWoLrJic6Eq8zXBxXAYGUhVvhd72UE+g8D+och1D4iP7d7zpFQuG5f4dXsDBTGpEC0mnFFr
P3SjRpX0iCXQtL11GFYr4KUtR1O/6DjRie/YOD48Er24AjM9GH4Lagl/RscUfrzdimJy+sdoEs6d
O5cuebbLV0SI311G29LCBZM/MmKgEHoLU8PmuYLq5/kEDyfOYKxr9hDepMLAOBXcFi18obCul3Sc
ieQ28/dqNtK/mwhlmvI67L2sYmw2kkA8Po0GvUlTlwNhTrNwQ249UnirTy4DMk0OsTvRMOrR0/vF
imQrprA4z308EMmP1D06pRJOxcE2hSOgIa1Jo2Osl7HLmFRb1cqr3dplRLidjNE+iBqObQTTYS9W
jvq5jm25i9oSpUX+7lvMGBVDXv+lW02WSglxkqUoAuBYD1d1r7HhHxVyjFdtAwTUV2QHNksVPXv/
aoM7vJHz6AcbCuLJkdofDDZo0wQG8BxtXMye+XVzpe1gYbCy3oyDvTFrYLnABtgJOAOW3yrhRH1D
n9CmdBber4fwh1Pi2ohGUUTiNyPho5w236rLNz1o3E724/GcMtDW5LGlnHvqp4J9Qz5km6RGIWci
M3hhlhGuWjsBkzfNzR+B6DYWAxzpD9fywKxvp1UFCnmkezpc593tr6Rw3Yq6kce/80PQXSTcSpbD
xThG+fwin2WLiZ4gHoomfqTHtlD2Z371WOdXU/Wtvnim5oKAkZc+vDK0/ErmypypQgvaIBIGFTnV
KWgvVVdZ/2RAmlJlL7+TD7BnHqRJYBcaQRM0SrBwmztMoymEIyg/8do6xP3eAhxI7mLpM1lt8geR
CWo1R/N2Fvitv+LLXzTAWpVIl9pudU6C0bBrT4E8zQ+Ea8zI5M7YIQSM8FLgpTw+ptv6bDgINUWk
YzzF1bhdr27nLu/SlVRcNIyqpMqHN5mA1SYLtAmloy1ZWtVPjrhwJYrseUHm1X2M0MKcdKHChyQS
Jx71cPDT2Dt6M9z2SJpjjqowNowwfybbO7hDw+ndjFOPylT6Cq/tlv1LgGLZY4KBQ9x6wc657H5M
X1T5dSGCFwkR27e4UVh/G3Bmt59o5cfgFayJcsLAURNJhc42GmdvIWZQwMURZixcHNfUK715IaIT
uQLGqLUZFeYrzCHcL0f1Osc+7wn/1PwCYsgBYlkVRMehTVMainEceQlPsWlnxXXNtcYCf48x/fjm
tDkNXCpOqHUdbtOrzTXdbFLJh6QPffYTtIdifX8MAXnFRK34vGcG1ccELi66t3jUM/R+yboxHdgc
O7TzlUDN9cEv2jCO1bu7KIdoRNYGU7oR1mhkSdAoN09gNANe68O+roZjX/qSuKh8bKIYaA0X9FUo
N7bcQ6ZgqJCqOrRN43ir9B0+YGmUiCImXbGnCsjWzMHCoGUEA4yx1LMLtnOuOuBv/s35A76ApKwV
PfnpBmMWkqwWoYnTMhKjMFIxJ1Id4Irpl6Yp9SwS0NZaqCSVcJXoMGrquwm2j1Uwqnn91CgaWzrD
XlkmDc5oVX5gLDHGEOZcTfBrd8ctZRKiiZEebm5pAxOzr9jACMHO+6DjwspfLKL0F+koTWbaaFYG
o0j+1ioulhnU+Lo5vMAKgXRTOw8wF/JozRIDkyUgPLqf+qolnw/Edx694Z7ZNhcTy0/q6Er2NUJ/
ja9nppkZBuF5YMSttTSQmSTn7nHduV/nsHCsNDxWw1kRbGi8ZlSGOnFlIoyHLyyQomiZPd9cVgU8
7bNIpXfBZFeVpIjiwB0WMBzqRCM3EOYZgHBkGiZ7t3T9+bojXKj9h0te5xcWgWZmVBapIy65/3az
aQcea/oUKqbjRG7om8i67RSBkx4a37oAfyC6W34Swhpz4SyklwzRbECGqq9wvnmslZXVqcAGdVeG
ACRLUUQozl2yiecUdbo7qC7sxadad7XwXqNln5CtV+/e5NymPHcKyZOKSGmu2B2tYbkQjQXHDOyB
HBawVEU+dfIPvm5qN6l1H0dCazTeDJczjfqBpfT2oB3bYZZrFk9H96qUFzY7dRSe1q4+xQ5O9fDY
qVujxlY8hhghUfGTSB5Jbq/u7KRbLd8NoAbNC0NJlOrRDWD7hAIc0BR8vSHDBqELSvMr14i7MVWr
glVWAihMTXMfUC6E83LUxTOFYoiILjLIpUDmPopioQypUBCfm74CCmsTinXzKQHGf9R2UcQejuXq
aCRJeMfmalhan4TOjE886aE1+/eD5aD+YHmT1ZxeEkPP6yTXDErInwVdqTdMukpf9wVonhxJhyh0
3mAq/d9f54RafUul48burwk5/OEMs2wMrI7Wdd6ikkdLSP9wFPdOWaeJ2PsXkXQgh7bZRF2fURXB
uyxatqd0g/yjR7mT+Ieovflejq3olkJ7Ig0vjKQ1md1DeFsrGQZJRor+i+s+i8coqFqPGdItuQCL
sZTXYDxrnoX7yGwAZJ+oLkiQeMGUIOYNZTdX4rSNQNSrMLvwB4wjIvqlxVbuqFyzTUv2dWSsU/N1
m9PlwH00nj9OgPhYHjoXxVqgw980ao1yvHiv06luDFCxhuHVPa8eM17IvwaSjK3VroUTNUQT1s6e
40E4L1KsDTykNQ0Lzu9zw/iY7DkKsrZzAS4eXGtJpltZfNu6t9kl9HeAjlAGJAayNa/OT4KDaLN5
zUiglMhE1wjrPLceprJihRiOkJxTzEPGGQiTvkUQSQoBp4O0Kl7285TAQ8wiZf9y0RpgHI+IHmeY
GnDSCyNCScmA0lPSJnj3Bew6ZDziHrmAiInLk4U6W2CeLub5sN+qD7z1hx1dHp2g3JFmHxb3SUsn
IjLQi9iD9dv952rQhyaCB6lD0zTkf0XcD6idnS+BoO5EpTBJDdvXYB2rMyHngZqnzA9O0ONt9vve
NX5ubipof1qTQblcv65OuaEzCobs40pBRjozT0pg1ZSrNSG/bGl0knrXyeYvLjvYGKAtkWi34BCm
fZOm8kWUKtdOh5V7LMBrsxbMKIEHzG+Gsgsa1d6lsDRu3lesYksjXScQCNbdueI5YAAG2g2EW/av
fwjXG6Xu0qfnialoswYjnb5qB2ppXjNpsDh6ytgLr2cS1PKL1sCaRfKlv5wwdkrwjFgdYnijaC07
sSftx3VsP5LBx8o4R/bkQltuzA1FQVOLdcMQmVneH8aIkV7hVU6NyLJnth5PJ4XORCEjDk7Fx9kJ
dRd2Z5BLk1eNcGaew37XCJ1DHcH3uOADn8AR/zs9Xes1cEjNarS3I6tQhkgCdufZvGHE8fTaQGCm
orYJEetmL4WWO6wEEJ9hTBxFUuJkuHRq8zWxeCj93sBF+iekFovw2elAbfTXoDMZ+CzVPp9nVT4w
uHu9crgTzNuINRhXFvRG7biCsOEkG3hjMwjFEF3Ms8gRJXYjJQnPH9DebxC8013EG7NDi73B9+sA
GA89cvWwNmYY0DoGoKbUW5q2QmH5A7EfvdYAFom8YaajtNXDhKarFpM5v+SBWHgDhlp6xVukwooM
tWI6G92bSuKfxHXo2QCRNZ3i4Jm/WzDbGpSFPcd5uB7Ptfry3Wi2DNm92fwv4EykuFIaqZdxGQt/
EXrirVRjA3O97PVUTMOXDG1VikRthgcbpSO+b1khAskE5Bsvnxv4y+amKjUcH8lFDQvJwcLr0aTg
ALez/sgz2bXcqVdDcBnacRPZCT5A1SqHUchay2z/v63cIbtIlsLJ+QO9E+mnWWRTE9PPUPvejNO2
9lCSMyxnLTlFRinYG0Ff85vahNPcTTRc1JINla0IOVmiVS8q/xyZBLRzo0UdlscZcXUPcBqjA9bU
2zA1r1AzLmXDFqktzkzolsACtBmdKbIFEMYkq83VQ5hT9SWUoS7qJ02sD6VuxisrCpp86CXmexGK
rK6M/ZHgyUbsR+RtUBJ9IVq1sOIXm8GYCajOuObpceHcrmUwMXH99hlrpOJg3QsTog/Z8D6f0/yQ
WGI7jiF9tZuZ+GJbPRXM9uDKYsrIQGLmqfhjK+fjC02J5W6eOAFPAdDcFTXCjy5WCnP+OSnOgv6n
/DXAot/SIt5//DYTjE9XEW1JzvwIBzlF58a/F74vtn1CpKKpy/Xj8NT3pAC9+qiG3lyrAq4BmTcr
blHRjzfkboHdqYqHnRS+Rme5v0Yy3+H16ugVu0atoaYpMMmjVKjIFqPtC+4tIJRvSuImVIlYAzYu
u5fzxXYf8tXeUqSFqblKkA4WwEkF/7FboR1AYs+Qbws/FQEEFUjNAS55UxQ7zR/z1FSSppn3zeCq
K4jNNGbLTMyTWFJ/irou8ibUcM4YJzzmuAdh5Pe1GhtslBs5n+V0PMbCZ+OiD6S+mnvNFLedX/MM
u1q1FTebkJ4myZlLvwLFkf38QKG3HQHCSZsxrcD9af0M9TluMHbPvXdxoWEhmTaZqKtih/Sa/7Qd
5yqjlNjYm/9nwlSJ/4F9MFTjTud0lcS3Yn4Gy6nhtXEMUBh3h3tW/C5R0CuL40hH6WLclievSffL
WRTa4t37k/hS8z+9VVYpNGoDiO40l/3GAgvebhGWZKll/2ebP/qoSUIbPT4fP34aRHAcc5B8x/aE
VOrs2ikXsbvX5FehiWc1H8snnEr8rZhUkNg9NoaT8+Uz6D9laYZeCdNCj/F+HuNdnz2xo7OcssYx
oPXaehtJNLoGBp91ca6IziGgynPOx79RfagMhA5HiT6eRJw5/8yrCK3p2wUbjqQUgJjQ65M+h4SS
DSYKsmeE4bq6q4Fgu0/3eVV8ux/fOq8oPzZeyasM0+HW3usEDSxVBR3OKbyhXbxForTKAUe5aHr4
bMpFZ3228+9h2khjuIBnotg0pwMTckH2AGHXcYIhQU4w5MAVjDC9s1s7RgbmZCGXPlL18C6gnPuv
gEkthIr+heINvt0PFdAgENN4XKpiiodHDXTotMbvkraIdjUTbtTD53x05jWB3WS6a536HU8FUYFd
pHNHnKycBdOxtdA5bMuUdoOrA64hxsnskXPrRfTAd//IX8enuxcjohfToQC9Dew+iVeWtLeFV69X
bchI+kGVmsVmL7TYWMdtJ3HRUIYfSObOEI71C05zimfJ6deF4GkJoPkQ/CyH2Il+wV2kqde5GfrL
CCPiMUzaBR86PrnWImqXoMN36tmZqONkOrOsvsWxoQsQapkM1lYKaYoqrEMUxnsIajrBjHbj7w2L
HPIWtEbzFjKi8LPhJnpFHSBjAwVFgwYT3Z1eOtHZ3/3kQiYH3e3gBud8EIGG3xw0YJrii89OVZ5K
ltNpZDyM1sR9KXemt49GXNJY3FOeJfwEIoPy06wR+TdCPO7UqGQ6y6WHudi1YERnHjVK0bs5sRUZ
sNbEqnn08agANFVAA/2rcAwwFH3HodSTWOoEzrc21ucsYOMRPAsePRkm0wmXlUTlY27WyYCjClzy
O1pbf5aTj9zsXdM6AJAlOIw80RDnySUzrnaIS4m/AwM6lvq/KPzAYE0hjt2tG/BPQLgKQnUtlNMK
7J+XC51PUSab0WPOAZvxyAAN869vBIU3TIDvmIOAUgaAtOJtRff5W4Anugha8oBqAuSYHdhbqBqR
8jcGjLBypksWtVPNZ3w2FO1vMb4dtO+2BA3zMJP2RzsKSyXoLTvpULHt3INrIR4LTVCVFEXyJ274
IKMHLM2AvSDyDSM0TEcdC9VZ9q6HXeECUsQ2vB5Uk9rEIVoRN4a6h95H23OfoABwqgVC3/Zv3/Xn
ozm55dX8lN3m1alzij0Y9pIPT3CbfTQ/OkTrJA0jG8/ECIOcxaQuubvQfM8RikLlENzZHY9ojp7C
dx3WRiNCOhdhG+onXB7fVpCHTuHIuk0ZKDeIF7/r2RVBo4nl645vGD1KffkzjdY1X41KDWBWshnW
Jte8DxCfIjKy1A1eKayRpTtCHQJ0AHJD0EADQ22D9klRb6Ik51yLlLFl2rZdyVg2tOPIl0iaJ5X/
I7aQyptiKESGAVKf/bDYAoJ/2MLYqcjAXHvLUEE/YYXzBrjZw6jh5BDVsh74bDzTKzYuZ9mQTpnZ
g1erAZjwsOKtwla4t+5uippWMl2tkOjFuqEo4uDHT+V//dmMNnyszKl6KQKgFrA6ggceHnwiTkS4
BumjTJrchjhy94nSUM4snxqxV0APPVCMyW/M2/6z4mZI4rkgnGXltcf8/c5ZMbelAqhsqqyRuB6U
Mh6bC7zMwyC+nJvp1mAKP+3vGIYzoQYmuDcaonRuwRTI+TkY5/wr9LV/Q6UJexgBx4G1rqyFQ0e7
/g2cX/hX36waJBHBICjZ0MZi3B7/C4oRBV3FWZma0Ikt2nmic/tLLYRIrbZilPlzZK0S8mdGlVmx
v8dPhjzb2LFq8ZF+ChVuYW3buWMz2EoK5DKtE//5cIi+3asRormdblb1f+aEjGGyH4/JOa0Qy1ru
MdWqZnuGf+zpxiruAakX2ymKw280FtD32K3yYd3Av8qEOLTkSGYGnoJWyMw5z9tasy7yyV37F4XT
R3GlJhq6TFYz35R39XKL9IIwJF0ZwmZQSaLu9zqp7fetkCLGyuaBt6V+uek5NXR/RwIzCKG0eUrn
oqqNGDMwQQ+5hrkX4/mYPQYU5fX7egm0ih8kH7eIwt10O12yZmSjXKnyriVTaWvK/jieelI+WOMA
vj/W9vCC63S8z6UuHvSfvVg7yykFxtcFJxhdfZFbI4GaGizvel+aJiKy8zzPOsoRy/4WATiPlMWq
Lk0kgYW9JbEkUC4jIzMAzL97qB4UWCEJEpvKo54Jq1iZA/bAbDfZU7NMm3E+bDAtZl2s7XaDVCdE
65sTTJA5OsGE2hY0QXsj46gModWPLGuMwFlkvRINNZuOoYF8Ser20Hhd3jn6GoVOpv6MO1L+XtwL
dhCCaSi0L8+iK6crzIIbdf8rLiznVhDYuCxX3OGPfM2KeilXZQNAgDjEKe3e8I7MSXlWnUPBJMBy
yBq5TcAp+UlWeBLUOLfn5qSOGdT7ynriBu4S6MALL1AWn9cdYU+Ez9xbVEHDo5z1lEfG/cwxfyir
L6UsIK7eLjkc3XMmi+p0eemSyOqoSOXtyLRofnprYh/QHbbp0ANT7Vy3zYSs4CamU1RIblmYapTu
UcW3/1EKvsMiwJKaCg/e5fODAzNB+DFsAvOagUS4kqub6alLswoYytBfzxuZoSWqhf6dgOqb6JHp
3UIFmkesJ7SrXKz/Ts3z1DUKgHFvEy3KFkhjBqHYeE/2a28ZV3OijJp9yPDfgG3hHu/Clj3PUrjT
StyLFEh9F0qLwDQLPG33LdHlYFQMPb8S/cahNKyh9+vLJdXzXUiVn1PC27RgR4kJrDXFrDRgk9Jg
bcmT9+Ul55tzHt+KgGH/WaVXsZNo7Xxw8DZcKRRavHMe99mHTO0QwBG0nrcyE8MoiCMZcjtbhBar
x1mROTkt53WQV6Orzt7Z7uip5TIvJm30gwcac7X3vHGz7edIg1R5cmMWGgb/GL66U5aURlgnlS8B
mztKshZc9/EugDXVwcT4KM3g9eUES2X38Ftw4KCf5LGpZtM0JaNQk3bMOlrhfROLmFoVbRCwcHSu
kxdSy3PqxGEWgIdlH0qFGoNXRbh8+95FAgUvKNoF3HGOxLGMnv5TtHX99HNHqzKMLMxgkUlvcWoc
5iXiLNZ4EAj8dQOBuS1qFZg5zX1hmYRhQUaYzAf8dhY57uW0EhYMx+c52/H8oh0KZKpmynYHnTUT
qUXWj4uascYnWU1kOlQhwqggxNMxyJ7LocdpZoQOOgF05gqcuhfbpBpKuQNPmGbS8pwUbLu2x17i
GuDI9vV6At4gGJf7lH4QFCSfyUklr8WCW0kFfNlbRm1PPmY404Z2W5IreLa8JPILlqjZGX4Bj5NF
mscY/cxrS72P2/3TtvtVriuBaovFi+vd4szAIzM0lumEIlRWpj6sXyOLdiBw4JJ8VIBDehtlZ6MA
ugqMzdSlHean8g+pnJhgP6nrf4iqjZt2IEr/ReDqPbzedvdXQp2D36PgQ9yHymardxjDv5jZfEe3
nUP0Rc6iYIxp1u5frNsJOWXIVQmqZNVPl1NbgPinqTNw+sv8dVzC2QuX7mk4Xy8wc20/xcwz/o3n
tolHPStAW9E4ww3CLskDqrESxztiISfyH5Fpp3RaNuenzfwXcaP8EdokoiNkbL8zguxQOUTG9sqT
SYc7fE/RP8HQJnV03MLg5uoAC0Yd2SHF+RlKGE6lLQxSXZF/lioATXiilA2VFBJhJQtfzwZommUd
zK74vJu7Y7d6ljTACZTFLmGgZVo9ijfbEh6h9JnfehGlmnzC4BYhUOd1/zDyhjqsJyhmWKtK+Ryk
qtPyxwZox6T2RYIN/sICAL2jHACTKq0OArwjtQnWz7tUYzFZwChya2hLC6FQOovgG3EeN2MVgSWi
Z/rIkUaMI+59HPUZaE5emhtXiw3wlOjOIofijYlmDP19BH0YqIWSwYwgNY/mMtMGvYtx8xydMWW6
5LO1ywqfwUb9d5v4fXsDdsNfZmYg8nqHojon19Oooe0Y9l6vBxLHumZ8M4NAGK8Z0mUaq7rOP+Uu
7hXeNklXxmZYbMSqu1IbkDvuiR1W84YrbyRRUDtM3zZ63nn/VMU7glkMK7u+gznNsc4ZZaYcpYIu
pBZc2HVqtUBDxxd/1LItvgyt78ST9PXin6BTq5OXY/DTK1BOLQBAqDhQL7GsaKaK7jpNPyElcwZe
RM7VdMb4yOjnrKueOhXSR4vFECQFa9wnKlCnaCK+plMyVe+uxKpeZitHs73f9ZDwYWShGxeT/dDx
iiAqOdIlFAorxwVNsUh1zpNnX6T3xMpMRG5b9OZnAGe1HwfsR0Djctwz/P/0lkiintYbd+sBBEyl
iahW05l8Bvz1Ru/LcKHBz2AaDWxl8YrLCKTo0Az+dnpgv6gIqZ+/5rfo1uPXc3n+2DnL3yR3Vz82
D37ytgngh/kIzih2fnX/0LWFOhz2F5OCdy9Bb8OQ4EAPneWW4PN6iMc3x5WIdWwyPXKw+umslIf5
M0eKo/Ay3jZLn35cD1AVjBCt2CY58KbLvDdAqvD9KTiIHSRAqcz4JV3Dyfz+mg+e86HirXWqQLZe
bc4uP8AJ26Zl49oXc5RBDPnQ9g//WDXkbtKUU2Ks0FNA7J7GYZhMXRzmOcEsTGugYa6lRYingdmT
xdMW0zwIpn+02x2vanQ1hlWZIidamWpPscePzHgfVQoWAR2SXzcLqPr04n7Ima9kubT+PMI0dUyp
hJA7pg1acjLkFBcE+MpNGFs37CqV5vcfFYqhmGIjwSlV64qqgaY0iEY14qAUWKpr2/MO9IpmMEw4
gSK/27w6TZ9toVH49LnJ/h67LD4ig27LUrd0DSlMy5Dvv5qOKJEpQxTUog0NCWSedvm4tjCXxXH1
1RAtz0KnIZ6STjCv2PPNfEP2e1t9NSRnqlNqC+XdJeCVxYzQ6FdMbwbiA+qeqDzGUUBEr1ILFvZe
PIXThuUDBuoIkix4hfnSq25E0tnAhdI59dRWxflBPj5eVV8ZnQ+gqqYiUeolWxQTSZ8wZrBP9eni
Eh4/jMIcmZvf1DJjd/DE9NrO/u9j77ah37iLvyqvp9/+TXavdvNOJyG5Dys1Dj3GtTKRkniLWYX8
YQ80NwPYcGbcImglp3DGcRtKnHwT5qdCe5/yOO/JQcFwJsTDXKwhqkQLo/LOoCmaOnOE0YyN+cwx
LjNa5zRT9yE0ASVx3Ms3Kv4zjufuJQ+67aVRMCg2MRxZD0YXurXj0nFFD9UZCxSMp9WiUQosNx2L
yfxPO6pe5ZegM4Q4rTR7Udn9sbEt0zGMUE94Qi2EXt38/lJf8MBDDm5gEE53EUC/9qfQL8J6NNOi
yYC4Yzk6yFxxVl4fzLyOG3/bC1X75jXhPa7UvZDk3+WGhm8wYwGKIb7lgstpM62k+A7fLLzKHXeT
406+bFzDUnM66gwbDULFqkiNd/HI+zjnZHJvVfHTd7CWOlLbwBK3bpPPur8KN1AyERlbLNJjOPuQ
qhfC0X+wLGeN0XB8QgyXUEIKLYrT/ckU4P0xPzwi3Ld/00Ioz8pqb/yTjETom7osOB4oAMjBuB8Q
xjyojGpSO4p9cVvEjFBc7EoPa+kpdmr9++bE2z3u76We9PSgwAa3sesxwtBt7hIfNHKx2Il3ITvu
BkB/Bv5I3Mo8cIOuWHfkgH+BCgWFOLIJG8ZoXF3g+gymZcp2f7luPHuSP47PdIScunzmLrDX0XuZ
rer3LU0j95JWb2cShnyLOAMJRK8Ja9RtPx2VPI6o85WAo+kdGsPCvZ4PUd8wzHYPWlhXWymeq5kH
imJ2OjcYOHQi89GZ0trShwQYFfDmFvjpYN/B4vTipvVnwa0bLRBfK77Vv4FdnAxzHK473bA0MotR
9xNgvCd49YWlG6Vqrx317Oy9j/5lwSKA3/8ZSD5jPYvb9HpyklpW3UNTKTtczttRz1MDLULs4eMu
xoLED4N//bXL6ori26cfnmSxqlwLo6FBfmksQk7mGfCgMx13vhxcor3netX6nPPHGEejRhMrs7Qt
jkqxrbvQbmd+xUDUqBzKgDp+rkASJtb5FKPQoqr/moiLl8IPT4fNMfKIL2Nuu7PaMYn9wKHhzG0v
MvSMeXrnAxG3nIVeEPh7YFk5/1LLUHgULfWEAl0qWdGxNbsNsXhTIc0+VN0e5RFSEopTC1B7X//v
Kd8zY6dJa5vNk981/gpgboWNtvXsv7Oa1eeLEgO5z+Ef2+Irce7ZXwaO62m4Qv/f6LOxB7bMqhtD
1gwLaW+OyWVrsVO5Gf3Pt6wwwqlvHeH/oPbbn/jD9ZN7WR50yDF1bgmuhLVqWWieZ6nnhzdRnDmf
wbYBytebH+vhlG48hIJfQj7ociB9bAkJvq3tF8E4cAynm4SpKrqVdPl8xcMVU5DZcYN7nzdIv86R
+rQZ57q9HPVs/KGhHekhZocLX3Mbb1zoi0pbmZo5lQy+K6P8RyvW9kwfo9IXxw9NYglduc5adWDh
fFy5VhATTDAqOhysuGxuv+QmXF48u5I1b5l6eq7QgYfmQ+3h9MIpUiGruA2v+rKhgA4M9BfrbLSv
61CR/IcH7A7OpvYUrajyhfUddFaSovFt60WBoLcyJ3TXjwwFVNsVHw9+GI3rN+mD4mP2ihEf6MgW
1azLDxBkljtFFJO0UWPnQu7urby3bowX+cEpD/WHzWpYEUaIylEAVGfKKfRRVbxm6/6WvDuexsN8
QG8lCAe7yGVfRxcVcU5X2illl1pVXOSzKSZPN0btSqVQQzpgPIXOYgYE7d3u2C8o2//1mrMrbIpZ
kNgRWmN5vqIVyD/0cAMiQDPfW9KnV+km02DYnVFY1FxvjSYUxHA1T6SUA7d1MvFsRiwPtVJJybpN
m2MgveNGAWuoskkJe7J/u5a08FYD452LJs0dy09Sjuw7cgxLAUIcng+GAkyUxN/UiYr9opWhqv9u
2tNsX0yzZC9GX1W/fIQPvZ9EcQ9p1cL/hjIT4e8V7PPrxP95lp+Pg4o+svw5eGtPuQ/vRulMQc2m
zN7g/3e6cyC6bIg39MXKKP6In4m7yCvuNhkJHW6w0ihFMja68+fE5WSW4Jcvj9jr5TVShCe22GjY
hhgbsGxK5NfBlLs6PEz03xWbZGUBsSXfQB+PIBLIFi+AUOxET321nYRUjn9KixyxuyeizGoJeNkt
nApV4lBYuYdRaTUz6dqSIw0s3rKEzErrbrYXiPeCT5o1Rzk96XO0hr9E/8r5V4KUZU9AcLAOTp7Z
dUFQfI/SjgQLnv1KenLOsyopGH4OAHJF5jMYmZV/UKYLc3LlHqPnMSZ5dm+77E1ozay9qCXTwyCh
K7j5egAuGcbVgi4DHRRUqfVFm//7s44kJPqCp1KOTnJa0IaLFCfcd6TEFAMAnS35fPTOwdavAXzk
M3vkb1o7T8wQNpJUPkBh6vd8G3ik2cvjueDn+LUfbIY/s4DbaSY31iSXDk5RiCTQs30/pgElWlQi
RSbDkxzCDO9+uhUK65e6JMHv0z7x2UT3Z8X15NDJY4dqYG+XuTPV3hVaFHK3uPTCHOX6eSLgEq4c
+W6NrvPkZ3ia6vM3QZ3wEPP/E3DYPQYuce3KtoXvmQ8NMljtsIRoIXhtUHLSlzuANxKpL5Ez78IO
DdaP5C9/sz5O/xCKweIdktJxCJNuj9gdwWjjU6/BS175yWf1eaHjGtbWJXysaTOP1TYB+xZpDmEI
MP8t8IOU/eXQ4sHrVk5HiWZLdPQZXF5L1Ki84E9ZGW1fa/ciJxZkJpKiJCACK7JpHjjsOXewSsr3
RCFp4REfYsHdkeXCbau98S5yCJCnNF0LSSozjBTjckzJgPoC6JQcnd85pTPEPTfiIYVbpkTiGHOU
RAkc0ZCXAksTkoXShMEsgXcmlkTn2cNaMMolmHOnPIE8oiRnDQyW0at7WyF3GUiV7SO9/s8eYe36
4n7KNRNiTd/X6L5gcT+6Ut8BCdRYQA4mpnjCch2CF+R0OE7AfjAq+EDuuxfv9RnwJ/ruEwwz1zGz
/NNP2JgekccqCeeRtyykRNQ1j5xxHBYHK1/fTGLKnzAwLlC/cbBZUseW12TcU0mAZC5CMI7hxPH/
2NuFsbqItu+rlSHwX1Pc/L17gEuei+aEGOca1wUKButfLxeHjyKkjds+S2OG4N+JXc87hzHjhQ4n
zxIRisQvSTdf2Wo2Bweb8YoDSIJUoQaX4TMwxaGJciLQszSlD++qdFazgOLBEsyTaPpnv0mLXOA4
zdCQzvNvoMUShpS9J8KH2bsTwf97xyojD6WkTMhoAhd7JV09SdVYiz4T2Hs9M/k367aclHs/G87S
sjtBY+4cdqLI2r4IKfNfY8H45ZIWMlhjtZy2uhcE57RiIAzn+kgEf4Z27mxDFtVIo/x15jvP3kWE
K0enQoFcME2s96QkLQ27BbKiD9A5n8BSknFm42qzUzZ7KK2uNYx4efr06EcuaugWQbhgKFi1yWol
4nyjMzVCWY+VWqDu/6s4+pR+fEkt8s/SOWrDh1bgQrG+UeszTnnqaueh0jkswgUNDdn4rnAKdz2M
gmLWQszEsgs9UJ5/v2Cw194vrgc7W/r/VS3Op3vvww1B6gN6zlp96kfwt6EjqNhCahMuqQmc8vXx
oeFZ9H1tZtXdcowK8DLAoUV2ec7oy/Tj/kwwp2pjlLiDT7/bPnp4IUkJLccpZcw9n56bJgqEO+r7
/VROT3Dfoly+XsMatHw/WJMxIFxFeZKQuwKmfFUbnaRcmJKsflDP986psDoMt6NFmyeh2/bRCWk0
F1sdZq/4tN80rlVMTfYs7eznnR4pYoRHhXkLGaYtZ1VmP++Q3wIL71MnF4EvXjOrgisgoa9Gl4mu
3x8LotKPmDDUiBtccQ3hYchtbU9m0/AqKqvkmVHp3jm6XmZulRX46VrmTzPRe5t6sXaz9MgrNINn
dEQvIeUfXjZDq7l8I7ZJJUjUmIJckDYN+48JmxrTnkaNuWby4NeuJPJ1B5dP1RZvB2rSZVPSaiv/
5bhqzx4eKGlO6doK32GCSdoBwbuAiN7TdBR0Sqj7IzxufXWEKaU9xXi01jHPEraQ1XgYb3q9J2kn
yr4nzysmGJ4prNqIcO81i7d/8x3Dk3MaYMvkSnoTe+eR2eT8BJTT8By4P9SGn228ylvpLQtminlc
/ZMe23dM8S2swVduS8vaUstCChV+Ovh3aFtycLNmGlhUIqbJZRMaVleB6R6EDF79dLonp5YHLjgX
mb7RmJ91QZOvcbXYUHwYB+ULL74frph4I+86UlFgCK39+hWUHhV4JVJJpnxge3LHuRFvVZqjBTev
GoJ38VeLiK4FzFqtZNFl12upeAcB8SI6OxQZJkXgpH8Ot5eVQEtbziI52PJzLwRwHPuH6WRI1Eml
P1DuCQZmxs5XoGSZ+UE3w/VC5U3VY/y6Ze8wEG0whrOnbPvaBeZZCySNTO+02Hx981APQMb6Ugor
25bdmRkziGWdqcmPX21VMEym8CLRKMttKUX7ZL1pWS+8YT6Gezx9mBrdTbHoLilinBoe3sHpDbKz
Ry3VIfqj3Vl0AhFhL80UJUyMs1GwScLR7GqNZ8rlIqYqriulz/5C5ShsMqLkhqIPQsIgph5anEfk
4iLxJcbmX/khpbNheKSTsVEMFXAcOzK9+XDagbm5XnePhGIknLzZkEZ2tseT5TvBy1y7HAnfSWlw
S5HRp2vmxtkTJtk+e+P1yR6+ZsaOmG5rI6xKsr0nLvRh0kWgimRHM9vfwMMhh4UDqcd4KxVWbCl9
fOIeSqfuSVMKndhL8picQN2NfsYP0jh4olQZcIw0r9Veh182F7lVpTLZGzSJFOo+XyY/AhGmOQE3
4Xphiblc0mK+DjDvAHOc+ww4N+8sbp5Xv2ow6z/8nAaCmqVJVITnvsy+NCIEYgdJiPyMG5UD8IzN
Q/WpUWfDLxChusrhBOg07cgbVh88mVIgVJHNTDR0ZOykwxGRVpuWx4nx8pf78EEOLDEfTPqF0/8C
tcknXdmU2jvnJhIp6+V/S/3r12Kg6hjvB+begw9eWOtQV/35rC67IY3smfW9+c/6hwOVpk5iMhIT
fanYP0cpDDtejjh6pgMUQAiWPWdWehtOUZ5IZ90quL2bSgApkPEbarVXU6lS2eVe5br45epGZkUt
z6Y+pmYTlwjobuptKhu9f+RXw6tooF9it6uZjZfC39T7n2JXh4AYQ/bTCcCSwyMiZCjJlUQ8qqbU
2eUnZCvGwCDwSEX5UAZpty5Xjnb0iXAJ/GMjyOLeJX7dVoGfs5M740r+i5YJCBTbMbdJfK2RknwF
JX2qy+bEZqAjfy1lSosFs0E7ZDJ5dVbpsGzzDsIoHGlAR8dVNRn382MIFuE+QrmUZbtbHAXmfjlV
ibTcQysTWSmyDPkmRh9HczWSvIp31d625U703+l9YEIbuuMRQdBULMjT3KATaLmVH9aXzBsCp2HC
QQePir0M5f/gjlsWBxhnaUkYOiW4+89pqn3LIyNxlSs+3+kGuyIjB0cQUd0jnuiL+6AgCaif/KKf
AcQWZki8DVQWFdHYPu8ooS7RHtJQA7uPxJAgwijW+9+mpj3zGREBXxs8a6TnEj6ggTd33owF8Wgi
p5czIgmyaDWrZ3nGc3+gUCDemrK9v3o2KV3/Em6VU2rgFaUonX3KqfzNppnH3j9Jp7kRgI5POqTA
RUMaafMH546Tor63a6bV45PM4a/R4uXVHCjPHR/lsYMGlQG3ybEOKRd+kwvToIYg7Cdxj4KpcfUo
LaWpYvp7uoXerKf+EAHxcvovVOjJMV/BiVUQQ7PdO0OwdpnGT3Es4RyexPZVJP+XOr866pKeZr2+
sfQFeRh+My6umzW6o0g85ZQgR40znngLVKnG2EtgJWLCVY3csKAS12tBpBSDc8exew6WtpQ2ndgn
kRrS1ldQ4WVqXPYBxQOawLLwO4SmfKZZD7VqIE0V9Xg3oDp5pfHm07rIzLLy5E2HClOdYkS1l3k4
objquZSf3A+yAuWgY1WxW0Majg1ze9crgT2YbRxqnBYtqFUw8y7CASCAtgscNPHtTbaRWucz+mdv
yALGwNxxoEbceo/Xqq2T2Tp46YwRUz+AoXJ0mYl387VT1corFT1ndwkoigDSejsLJ7xeNtwShtwf
ygEX1nbBh+gSNsO6qDkV1X6CmyvOiKD4pnOdRVU0ORu9LnN7/f6TvnSKPpzVDsiflgOQEr3tdas9
SZTXRdoWt9H/n2Zp9wfG38rmFwYljgiXuEldD0qFnA3qexf8s5UZ5xxAQOFOzHeFzx9C/Y5cZe07
ZFJJaDfJf1TL7pE01xFJxFwVhHiLrLCzJKsk6hxGudXKJYdMvb484IzFY7iHEgL4yxS8wKegjipr
46JrUKSf7rB1fdTpn2VMlLuGvIqaAxfcqYid3V5q86TLwyWtbUX9GaB6Lj7F2C4ElzZOPy4nemDP
hOliyYpzmOvUOdyASvHk56gZr4M4BFbLjeBUTGesCVWRc0IjEFbU5JqxJQ4BtGgs8+tvTonSYHAi
9AqAnFcvi19wn/hTfRq2BFKeGXhEgnjgLWuTBpNN3djep3kClTnyvCZzLYESEEpvynj+Itcu0tMD
LzYFDBj3T5mBLEePsJoqQJQxQTYtW++cQxvAVlKbJdQ2U4Dht5q71VMo8z1ZdYg/e/AkXGxuAi6T
xXA1MeYMJkqnriD6oL5FhuvF0TLyLF+bHtx506zfRZrKGpEx8YU8sHwuHzDQ3CikFQ3Rb+ba5+aB
L32IIrcqyFxDhNRSZ06b7Ldx7onNpivwo7CnMw0GT/gI4AINmqYu8MqktI3H2R5kJlhsQ5EKpUTg
O8Y/WcpDytu8QgstD+j0HRHyxL4qx9kIW9KEML2ouWr4B418CioZJIA3esIRbo4zePGvn+aTIUCc
ppx/acQAXYiGmDzujgc+7vyEFAuCzfPSKSx2aFsjOlSp3TI6BvC1p7t+Ul4Pn2hp3lfgGtjHv0+T
JZO52U3wooahMW4tPJIgC/R16iU/N3n7yY2taHkTf1a7Fjz7wsQGKQ297taUiozkDEJJC5vG83KR
Wy30Kx3uGB0UmiKB7naGFWE2k+hLKOpeH/f0bjk5316ccc0Lo17CFJ8RbsIzRwDSI1/wBkZGH454
VGg24xI2lspRdP0I2j1MrVFcJYECm6tWY+P/zlQu4tv3bt1CQh+J6FGISHkV5MrvU96LavnQcRt+
3TOQ/IO0W4xhWeskKG+eHBWMQJedLVN5Xh9TPlvQNnt4BkkouIBj7zfbDIqGanNpT5yi/UeK0COb
H/BKDmzZ3GgskHe1ETHspGnBIVhln3ZMR8dC5/dbjuOIzGXbpcKx6XFyIKoNh5tDY6Vivb2bCoZU
dAHqp1qSpQg6teNiwd6i0dOqHHXG4Nfobo9+E1UWlWVihTwdX+89oh6Tjk9kEI+Swd5Vl4Ezu4N8
2/052BMkj9Q1TuosnLlJ6kYAjFt+Y8+WnWsagQ5ITEPF5xJ1sV3CS0Udd7mXNxWzz2AfBVpMrz9/
M1lDJeNYVj21LeA9ktBUGBDhcZgfeDV1MEykqI86qEl9SShvXt/obdZSd0kz/Uknggbm8GDIkUH1
RmLbtcqsG5J7+3NzdMDfScDgYExbu4alcQXHWzmuZVFqQRW2BCbLr4LymWkBkVqv9yWCB/Mi0SEO
uHLAp9wGcQ2rEO2dBgoa/28hJxNdbOLqxDe3K945bh3qFhAbKMpgIHHVcybBUMKh7aWziGBG8FHC
sGyH20/2jDdbdUBDF3pEl7lY8ODynbV/sfAzOea6Bw7bk3KVm8B9EncUvpgRiPk2oVrRzGeJmBPg
WbKL78u+ST1n4fWJC6UkDbTMkkz+hhrgvatI1pnq1z1MW3PnSP6m+mgSUkg+eIKIGvKJYsF0kWN6
KmHl3aVoLR3EkSGymp1Wy9s1g8uovXDEsX260Rqldhbtm6jcSda9kUbg5pq3po3PUAa9UqjxOOAV
xrRD2/8vZW7wPUmcaY2v4wvh/unj+z2DGgHPDUDjC2HKVj386jNqCz+u8bYN0Vvuj/mfU6wmaBP2
QYMmBUMnk304Isq0AF+cW3FuK2Q/3gz17JSbFOvsFKM/PrqggLWlmclyCQrdLx3yqHHHQ9PdIMXj
qBj3tDQGuDONwXt5P9mR/7VaTdKfMXe3UBpyYtpYCtIwFcMFbmrBjZHQv4x6XyNhld6d767uaxPN
c2fvzDb4Hd7vLeOvryO2oRf1ozacNAaEjuWCXS0+1H0r2p7OAco0eIBeSOmMKoDxAnCK9NAOZAiB
auG+XNZY5mVlO0c+qrjybH2CTxkyzva0jlp1B9QfJvAZkipxqdUVA5ZOnQq2b02Plj5FFl7MJqq3
5Km8cN32qIBJbm/LNPKPlhsN79XX70lrX0OTY8ecytbQrB8FyGam6AwyQmzd7hAem247Px0TeTn8
96eMn8Z5o03XiGjeH+s7nUdmqur7io6BbWt7Wzmr/H07YJF76gXNtW7EmlrZZzyxjPr++ByJDTIN
sWFayIxcYp0xV8zh+VFvfb3gM0oVhymsR9ts0LNATwEDRfkkA9cbC2QNMOnlQWYegX6rzcnjX7U8
StyAn6FRovw4Jpn1d/CB4kiyzR9tJyo/bP06IFqKrxWIHdTPyaATVzkJgQMmlH+V74kx6wU71Ftw
t2DxO+T35BToCJ2PKNizJurmmU9Fb2/hUl+EGseHVnui2ykSHSYUp0bPn7q3zSWzuaiwPLItMNqE
/geUaAOcunNNCUF0pWf9sbBSkGEPB3XpGtKVrMFUlRZXUrYMkjKZVvh7QPN8yRdTXkVt0vu6CiGl
TCTalUumcixcergpnQAZx3cpad1ELrJ0CiabVD8GMQzHvdR2R5BPW0pxCn0g8dCNL7zrccqTpmIf
HAAz0Czp5FqHJUEhi3VYMxB/3SDO6R/B5nRYPueGJaSS8rSpZL1g1WQ2w97sVd8cBN/bgV9KhtFp
qLUS5a0hOA+KiGsyF83vLZ91woYzoraYDSgTpoOitQ91c0HDYbkzlSbgOwwAOlrgsj+aI1vRsxfV
adN5XE/ZtdRpM4Hu0SHA8QWKqtTdGo6wlhUU+Mg4agNCb8ucq5roYU4/A8WAZ6gSx7NVCrJzRk+M
TN9qHKgiiiHLmEPzRY71xWG5EtCdhXbQYNIGwJsk+U4qGM+qHA3MlSX1TBlNLseLX8ZhPpsIUKo5
ffOg08C/rVpevUXSjl282gPBqbRmoLATVPMMsaAu5JnF3I/mg5w5Gjt7KA/6OnrG6MfcwI1sQevv
FZAE8MZ9Pa/VmfydNt/wCOw1VNAB/hrQvujfEuBVa2WzuvTUeiU7tftozymLHhYAwZ9YQOgm7N53
dDgExBoOH0+7Z91QLqzVrlSCCHT09fAXpAOB74Hxu9pJbf0POoRZMceXGkw4OeVuZg1bMVrIj48l
cNnSTVa56MlGv46qfmkZMWmdbFxCIMQOIjEc506/a1UfVA9ZwLD28B+4qzJJ8iP7eS75IvrqrK9j
zhBzOPzKqNgZdyJ/UifGgZKC7lBqwGrWjZnb33anF/yR8Poh/o5p3J/qz2DW02rFRUtKgqYOvtI8
NjmTOrwcvs1JOZ9fZKiF3Y2iyVMMnji36Ph7FWHKa99XafoizK1/QS35fL/x651D0KzSOUtPKSEN
PCOgDYtw+9dOVYizwUY27uGNJ4ARyc4gZxmvx3OgXEMzh8R558wS9gsNFieecbkbbINPaAyTtbjs
zgFP5lAeHZki4ao/PuqEu3qXPVVmGGS9eUcJWPUexxl/BB0mooURiE8wwpOqsM32RpGF0xbEC8e6
/ornd01/MeS0AAdYelm/cVRW5vlL9Apuy9XzG3d9rEcObklC4povH1GpBcDLOY6j12mpu06xu76y
27AiaK0PNXoL+stwGNYyjis6LAQctIYAZwebiCg7ZL09/yzUh8i32cuH6H1rKT3gfvZxCU3GiaSh
Pfvmpa+sqs5EI1Qh+trcDu6erJTYhKirACBMO9MKHFeoXAp/yySyBP/RSSEAnJLLzpfs+Fv0kY0d
CUhTVeON3pKH9fSXhvvvviXg6VK+pNxXGIAseEqRWo5Sd06lncsGs5x1hJakpYELxfoKsYjMs7n1
+X0oorj6qOdFBYW4W9Pn9216tJ/HG0Fo8UfHBJuvP/xWKdDaHWPpM2tgz8eXqHMJBOkEvzKLSJcw
e1bQUzJ/Os93GjmRaNnK7e+nAs5pH0MwioLT17z7aefKgRs6oCB87+UX6zfySatuvOV0zgoYh2HQ
Q1pPNbOP6Ug0/87OQZTllkeCRLsBf+ec0WgrqSOcCZ094+7jh6wUn0B/7v0u5HNGWQEc1dTL4W6N
KKxs1WPc/SRZSAlj+EU9zpWGlmWtHy4SkOBH62f84vv/vQs+CsMe2ciw7O41CXJRxjlu8KXgwMqG
Wacj0esLD+cxN6coBkiHYiei36vmGXqJnhDUJ+acIXgf/4Lf4o04MaUlQqVyBEyd0JKR9yZigKyr
VXZ6tAR3nNzwKSHp1ZlZQ66Doj/FNx5GMCHY39cE+TQrGtbQQLHno+l3qSHBBK2SY8XSoBKuvDQf
Kgo3BhHf0SBijhOLK8+25iUlUh+US5PNAYoyl7/xt3SnLcZkPJgeI4sZ9mhqWwVanKq0BGm6xa8t
S359k7bSg8IQTraa5gwYcc9vD/mCSFL/49ayCYn9TBjm+7Yv28kmEqB4cDTTMu4K3QABHl2VT0LK
IbQmzb4Up19wP/c49JoFqBqMUb9g4BHNB1BYHw9FQupMytyp5uOUfyPJUMJSdU+7yKrg7njDzIGV
HiuOeVhTwj2Iu0+dJnJM3nTLs+87Y2v7U7EbVoG446C+uqT9UM+ROs2DQJnFS8T37GlH9SMP02Uv
uV2kqjNwq1DKr+RKrf8dy4/kXCYERPKfGtKkf/AfhZPmEKwEPtAoUgNKH2XpMYjSlBoPFbEOdhZP
T/OemWlk5zukWB5+PJ2Pa+3ZtFoBSHpGSRevgDc+0VflffZnf70vu7s75B6Whqp0EBQhaGpgg3az
s2RRYSDZxGKobAFCDe4rRiOrhQhbn2+0017r6RqU6AHWAUuXpXQTGWNyfdsXPdW42R/fsIJ2K1iZ
CVtWRMd5KRohcfPou2ueDp23thMd0njDwG2Fdx9CHBWWYynanqQGRAPLKSEL3CxxG9VJ5eGII2s5
6SQ384mRLTXlkOq++vVPkY/rlfHQnQzRnQ0Ez7cb1+FwCnWJDctmGzhxEIMkJ/croOXEGhJpr4Ej
jIWWGsDVabWIMFxWrhwUFaB6MDEpC4FvsKF0pJthT7anTFI8xNzpMwFEBAgDNcXPtdD8eRgJBjbd
VGfAMjjCahdsn1AIGLxvRERD0UqYKLMMRilHfrCpxqM+YpJnBx6sWKbA8Gckf3Sl0iaEulD1Oj3J
VFc7/R0jeBKBGZ+mnEp3XidQaTXHlzPgEjH/zWgjzeiEalGqCs/b128vwSA2M20tiXjhc6U1sKR/
/CFoJ+v4Kh2gDWUccFF9Z5BaPHGA9lAEIjw0RwovYkVRcf73YlmVxURJU3sQmXNHN95PNg+Bsp0r
MUtypRAbE3R+juvaC/OPBtJU9gAo19OFfLWMOfU8IibCJmvsHD9HS5M9T/yFkjUN+tuHgeUBEvER
TVVswUVcn4zQwlTpXUOj2OR8f5cYYH1Ip/KkF9s4CBcZT11z14przWkh6yZfh2G4+4xuX+JTu8wZ
8tnXT2JzXDQonf1bG9lIWSLeCHOlWmz/3boNbXv+mv2NYGadMUA8w+IbLj+osUD172SJcLAw2+pT
u6MyaQMSVxY+Rlx6ufNODNOHK5nbh5ydk2R07bpvgnU3V6ED5fev8bEzkO3ehMV3y93qq0BNNqDk
fK7gXuyeMwTzgBW3bJ4V9wEMVRtQcOyZAq8P5/hQMEJMHJIrqYXIcG4A4iYCK+qf+sKQcQG5ODsy
9Zhe33kfkz0R28xYof+D3Vfg66fNM5yIkfEF21PJwU49zWugK9E/XlJ2nxBqa9lRuciNNMuYXFwL
6ZNdG15dTsB1KaVAA/8GWlrAShgwJRsjaQBZFGq4r5zHcXcnERx86VJNPW319K0NiGwc+LMbgyUO
PqVX+v43mRomDYTXrVh81GLk1Ex1kgIN+cEBAB5h/q2EMyaXOeDK1EOYSzlcc0E4yPfoZ8z9hfLp
r25rhgbs4glEsSamdnT1ulVPAFEb6Gss1n2X0b3HDg9jCqe4zzzqlS8v/Ao/k1D+N5icw+JVum5c
uHUptjHTilh8apBsOZuWe5+N6idex/6z/EVOYAVThYugk58ZvhfqnLSZoWCJ9IWI4VsxTm4wCYRO
tm7HNmewnfw3JX72fBeX1s1NDmndPfrtw8ZLMCsoZiHm+gDqzn0fv+TKRHVbyaCIBBcCwmALyROM
6/akfTIkJj1HVqZ3BEgFU/spFU49dMrB4VY7cHta91QO+KS5baeXf0DB3ux+d3EaXfxJeIuR0CZT
8ZmnLddqXGRT0bnA5WA8cm89DCs6U49REr2xmpxh/mzcG6ifYzJ6+3BhtHPFCxtAxl/p60xt8Rc4
CQeH9s7j6fB7z9Kr3wOsy+s3SF1OZUEPaOafWzkZC3TqP4xzyS9Y646K/UNTwdE4S4iO9wKRlkk4
V3nQhtw3JDe86rCUZYhNobyNtkVjOY3j1SpUCODVN2uahuzGBxDd+OhF1m1XZioaxU8tiu3p44Vr
DWZuosDp5LWvmHuH2I2gvDAsJMO78gABXRREOQiUtBzRYrjc+ndyRE0mghgsk+weEJiMLNLy93d6
+0Cgte5qHw3FODVVvh3Z8vKZX7fvbeTLJ49xmiyeWzeVipb+vU4jj6a9nDd9jh0gc5iS4c9SOvuN
JCm4GL68HchZRFIUI6rIkvKzexqyYY3+L4ujL4YtGYj+sm1UVsu9FchifdpmwP3wXoc3dOC9TIbF
6fd18NAQ47R3fTpmUyX6OswWqN7C14FAY20lGkr4Cf7CmlcMEYmSAEMW1iMCiCUsvrQfjAqmsb8Z
grEA93Ql35mdmX35VQbMPBNGJMZ8LV1nVUtrhP0I5RSDvtfFZjxSzuLkYvzvKdlK+7rkqVLRKOCr
Vp/QqDqLj/7YB4qlTcdq0dZMAunDdZaeFumJ0kS7MTLvFEMakCzYKoDr1S9BrxvC4Co0RAQ5VNeQ
oD6zSv2ayqg5kytyZwQYWR/HVHrWRJUqPAPHI/9H7MZEdHLiucvfVb8+AqdMKVKUILZveXmK4Bb0
MW7bKMJeerXV4Hdnn1b/I3tAhq14qhe0U3wU9w8tbpyL78wI2NoJqJxUhpsswAJxqK1gbyp9kU4+
aV9p6O2BzB8DsjbmHeZhWkoyzoJKOWwiXt9Imj5Td9Oz3oFfCgF90dk3EoPCqF+S9EgNp5CPY7U3
qyZAwYQafbB5UOtjAzBpQPUx8xJPTu3rmt2xASDuPgPBvDhTLCcCu8LdSnYID3+d4LfHo7dUUmKi
MXvcLdMC9r2xCYfmoBQBOZqr9MKGAqv+WtU6wzLdoU8uqsj7HrCsiLbCUuKb6vjmWWW5Bc1V0HsO
2Vp10w2UG27khflJzkrS39K6lthYaDYDrHB8tZnDxdJi2CkskTjyygXgWLsAThqTqbBD6ECeIvap
eKNFF2uhnRPtKw8E/3BVDTROJIXmOyfMn0viIngdY7K9126mOcrzs1+QpNLwRTalacy1QBf35OTa
+QRTtN4RxjC82xOownEvQV1EBOKxlKMOQM0bNXIXYZEmGXTglseEefpxCjOEYsqby4P0AU8A6rZh
zK0U7H0niLPfKHjrrKZv2X+cDYOt3LuaKG2GwtSVzyRpZkA0CbiFhts69wQhgOvikZxEMIdKz0L/
jrEqOSEbJ8Qk1ZiBOiZjP3z98Lgo8zyZ9LW3LJ5g77B+tQAjkyb9iZZn5Lu0JpQAPtJc8fm8O6lu
MieQbiTx13XLs0R0wtXGOehoWf4nBDiksEx3j5G+Srmq2YUUm3YGBjHtRxI4tRP9RsK8BeJzFCaK
wq5DDusfxOc2sXCr2Ab0j6gJgzHmE0bkvIlt0i2bUk8slfG4tZe9NKhTS4UOcbzgO1YtW93Q34zi
88lbWW9VlJ4OMGo4SfVDU3gJtDTMSOodtmiRhwqTcFqcs25jFw8Oyp2ZJEh2fzll3DAQDtVMwwfC
2I1OJn5M2mcT1lHDpgcFZRweoapB7cFRhru6gXmg2gGnsMJbBGNCUCd5hMNco99Sy+QIi3xtjgYz
YM5wasEXt388fL5b0AAhy0zpIJFixdiA+PZZx5Von4YTgtqL1KIRopGBdvgTu7O/LXRqPL2VOn7e
5UWsPEmcD9+pH0MrqoIT6BlA7JI/KYg5RzXra+wwuRngUOi0XuIOmckSyXm5B8kZ8uUyB2x3Tqd3
//qWCyyzFfPSCOxjvDHOM44e/DTf1jmkyayzSpm9ri/vu/7MIdGIF6Wi+fqn1u7bM5ww0aRRtwvo
bPPWjgvmvPaFOsD7vtVOw0wzBQnZXeA2ARozVfxQIPJh6i6zm6D2tBqMV5Gy1m+PjrmWnby7oBwN
O9KcoEbwz0MzqtABjC+zNL9P7wU3KdPFQVpEBvPcSwvp4fuH48xTiZuQeTCiWTV8TX1oH7CzHtbB
9zLZ2xpAVzGkRRWss4Ey2tQ+CjJbnu+smbd1uEHINU2dC4wIvXKAswlQtQ4oi9OMPsf4lg/j54Jq
vidAVZt1zA89U7LX2GyMfqzzvJ6JtaZJisOV6k641sFMCNbBuLhbnyMilVU1xvbl4SLsxlky4+dI
12kt69psZaYJMHvQ9dAceldCv6e8MjGhcmH/wbRmqpvGon/0NEVuOX5h71wEgG8UFrgeVH8SsTPY
XeGb/8KP8QJHNwaWWv+W7TQNg5qkZncAeT9QChx0HrSUWjZq2RxS69yi2IwaVzJqW4XfqWEY9zUf
Py3QiDGzef7PivOTuZJk6xbsCGEsU4XJB/RSXruzsS7X0ui+9n1zFkggFB306MT9h0fJVuNjo83f
a9pMEsbjYqAPVR8bR+SzCfDApWQALviq9YlkTlcYwrQPCmUBDAXTFZbpC2D2XKc6Nj1FOBZCiBuf
EaPeLqwxTYWDeK5i0hxU1fYf1xP7ZxFzzurFIydHb8gS4chsf7dBIfJsU/1CgjrKY8BxEKLv5GJB
5aK2ug+OUegJ1TQkHovQzj3ucKvcI19hXbcNGYAzu0U5rHYWhmJ3ODcGTvx2QqWFtQwKQ47ujQRV
cWbnwKKFklw+pJYBsp0Z6t0kVvA9aGLdMJncI6cgtwZVOvgM9mkHgpb/BYI0r45H9bztYi+pm6iI
kmdCV+We0yPPih094wkDvW2behjTp2bxYSHX4lZrzC3eJjmBEaGLdnMWYyKbEvaK7m6sOacl6j3l
Da+FXce7wOkkGURY6Z13I/y3pfMfT0wMJY/bZ+zR3ifVU2F0AQ78RbCLVdjKmOYYD9RDi6V9OAus
PYFJC+5A5Uhhd9MjpsMf/O3rpOOIZZgpccqNqyuQ8+kA4dKMV5HIdoxi3+7hDcagVDML1j8gDVMr
Gn2gtZdfR37MSDjI4eOUPulMGUWBkqyo0s5aKJoNN5V+w0oij2btZfkZUZh/utzwX0j2ANvvW1kg
Pt+GNE8q1qO9klNAP3j0ah0Sn5zXmVFToOVAcuGy2oIL4jSbPN7dbAVyAJZIWgfLfucOUGgnFog7
kQljR+EOR/6CopJyTz5P0Yv4j+V6kTouUUTUi1fid8PGF76wm65PlKzqQr1kafQqh/5yi9G4hnd+
x+X1+i2bHIbp4Xdm9cxPDL7YoGyocke0xLhd0VKVAuF3LHBIZ//a330m4I/MKW0suTroEQglBtah
PsCsSnLy2ACbt7CbA3ViDmw103TnYM0+N9JzDbl0CMNO5AfJEgR0ntwbeGrzHbDMs6RpcLxUJwcp
SUbf7baGMXHUhmjyaO1CjBdQUVlf3VI5VePnSSCuDvOiYAvJ8oMjQG/sYiF3kquuagxoYAltx/Wi
Wrpvm6UCVGBHbwnM+mcCKyy0ryu+VQRAJMCRvFAEvrvFUkobJ4OoxxQ1I0yserHeREaBB+2ZCOmZ
mLa+QX1EcX2MlzkKQDAG5MCIT9jGWPV65ibrBm7Tbgs9cU/IAFqLjBYNjKngQpuFlBhqUrGm10sH
KbnHgt4i/LVSVluxm/+W0RpbR7Jt2onyem0taI+ZbfdkDeN0djAeWC1+SQ+cis3uJk+TJF1X5A35
1klqI6pLB8hEL0mJAYG09tVcRZmP0wxzC5/cp71K8EjQ+xmlh8SkXFruo6Sf+5/5i5/OvCAZ9E0U
i1ZmwXsXy6dyqSphDWy+H5YvMHNyRV0aIFiEBp+x2WMEukMNG9T9frt0fUoKCPJwgfyK7ZX9RdIc
xOX0WInJ+UzWRYnz1tqZm+6ECHy42jwUvJjENN9MMV7Vn9VsuAnJ8jwaCmKu6/YInhwoiSFNpGXC
HPIzCHi5f78hCarvxDeoFm7FJgM+DHKors/21C2hjFA3kLOzQvUR/HoW2dPXQV11HKD5X+SgqFdq
AuwWU6xyB8mfufIgsHzZzbTGTrV8d2oqxaRRQlOTtdRwoiXlGqm8mABSdWJbtLN+NoyaLQ8Cpvzi
mnvGhRRgBy1CbVBA2q9nw5v57f5T12sDLvkKHVVh9d16uhElsKmXSKHr+t3A+pn7Skuf1FyO9RsF
h02EAwZLTRw1Z5DvlggjELyryQnhVFCBOZJyP+4afTLzFfGNJL8zHA8fBmWI6kpwCLnHKMeXufbI
9yRdwiU3G0+NjJtzaclKTn6zLP9AEiKRhvltRDcte7nWaDN6mIxk9MFhlyGBoBqJwt6Z9uhWbmhH
DM7oi1DHXnEGrTJLh3dIljegG2dhfHajTlrxV7eRnUZgv6y1j7QdwAOu/M3sUe7IQ6C7sD4+T68z
n1ZOEJFR0Bp6eUGjOLjQO4f+u0WVbBcCJbzjfAZmaR9jEXIeOtn/Tq1SmSpeA4Yyz8Err/mvW5MB
Gwv2Jk/UnoxOHdJF4IV4OaPQ6izLekMQyJDJNyPtDRvI5REMWZzyr9TidNKP7GFa00CKn4Ye+64Z
bJreR0aSPxi//kWbGdr8N1NRz/ZZ5C7K+CMiMWbH2Ntj5JKIa5xbieV/psve1UAtMu6KyluvHF/Y
Ql/IW3tp1UBs77FLp6vhE31FO96T5ETnF2SdZGM/XGMmC2skr1uhvRFx+b2BV9VCcxP63H/zupzS
KvrOZG6jaH0/2+95lmiTcSwO4qWYMKLIAYzHP8fVzBPbTBobna8Y2pSwbs3CDB2gZPeViochk7nT
tDskJ4BEwiGD0lvBK8k2YqPnXMsnBUCdC8rI1zU0/cYXew3/AMBjDkA6428lmpJKUX6YexZVLXSS
ZxeN62KJepqpucceBDWzQyaxUxrQhEbZ8NWspWNKDGLPGeEsYrzeXww3D6Bbb1hpgaLbtA1chL89
+e5xf+enVnADV+UROYNiu6ovZ1APCTINUTzODawNiLvYrUQg3Fd48cImlDfusIntuEEnYj6hC/VK
JSX2h3Xt+UYHzK1BC11MawFkgXRZfS+ljD3GVn4xrskBatOtgZfmfMJrpXsP2x2F2+V7GSMmuQ/B
J3ojbbkp4d9q0RKUfqHGACIkzHSRn5pk0rYA0dnH/4N+qJ20QTfAWHxLyITprDwhYhI4+spVUxBM
jpqm+ga4Q11ThQ3/plnEKBKIIZ5sNIw3zZi1FusE49mFbPBCp1tN1zWcMyzJ0A7LCbfUVWibOwxM
FEAKjQ8BlZbkqaZQDxg0nwn/89Xl5VvuCqf7RwXcI7ecKJdVsKBq+dJXusWvDht8UQ80ylZHp0jT
WhJcMxGqCYec5/eakzEA/uUAst/Qg80dcUon8URFhUD5VQ0CQAbad991JQxnF9+x4Z5whnLjzF3J
TwTawTuV0sEEphNtVo26Y9A2kPWYmOJj27CSor2+UDTPfaukcEf19nq9A1F+bGxo8RFZ3euduInB
3SylkQjLMfw5jt/ud1CyMxO7JGjnplexI/o9pp2DDLHGly9YjwhNP7Lt/cZf2NNG4MbzB6k4QNDH
2FMZmT6duU7xYP2NXyXteheLcCT2ESyoUem/W8Y/+P2GcqxhW7AhdimXx17OCUJsy3cmCMX7xDNK
uYubC7MhKN45wAGcgJ5vAqBnp+7hntUnDRwGcaQ8SISXGxtYZXoFVBJkLEoqrjNIVt1nx5Hn7/nD
6Z+J0wGO8FzbZVADPs6/z4j7fk0hAvtcc0H5wX7g+Ops+d/9/+MSpl84T9g5p5yM7aAlgGvqxbi6
sW37kq2salS/VnwieHkg8PMtueZo8ZgKdBqDUrIgZYvSb1MsqZoxT/DGpLXUx99ZyMybSjpxnfk1
9VMC8u7G0YDd2qxbOOOdoqE7U0iP9vnaNJjvrZ34m09oHXuPxyE1ljvmgOhNg9h4ogsGcx4j8sXV
7xQV7K+L7ftf9xWImQRoMQhsqPGBJP6mtO6lPB6/6Z6oZpENMfEaD3+dWbgEF5BMGSsoEyT+gTlO
h+mKv4LFOurraf5eJqBW5NAdSmVHakf+MAz9+rWike83gQAFpL/SBtHy5k7Yjb54xGMiTroM9EcW
awS82uSmdu+bxTrV1/pDHXQtZLhh6MTNHIsqH9T6X/N8xnI1LCUauui6Qjt77UJUsyxFIKKtFWce
d7689U4OzsvT/oLBMxp9AQC+mUQtod4fCL7s4mSbv/r0ystTCHEHQpjME/3iHi2WMYaCrGeQ+zA4
J9zYgNqpvqT59PaXcikp3Lo75FFH4RGhAN4L1PBnZ+t1beV7rVl4pMhHHpBU5vs29XIxIrFT3wTs
8AGuNzopJxVX1uewTi3cWEUWWVZQsc5vR9NpmyQ9WPR2oIy7cF3ZaIB+jRLYiAqV8pMvKc38ACj2
8/dZYOTvjWtsNA1cGmLqlK+drCv54x/R+sTwiC+WDDSJDwhHqs3hvmeS/B/z6OzUjRGRQgCrNmhy
ixxJ9vwPUaGzG0/2/Vx+sACWDXVl4h2jO6Q2BwOz94HADRU7YJl43Myex0j7C2EmyGvsWrEvx4Mh
B2ykeQ2ZFattkolvtmA201u67ZWLmuvxDE09MbgjXTR/bqTKM2KRxXdaimBWEfhqXkEfmAwcXIbD
yiiMckKROAAmFJ30F+VinNhOvPyYgnSJuhCbK5wMDM7sPMO5BXEqyMTUDe+TlbZ6rYClQQh9hoC1
5LMj7VLl5DcDrQfNSUC3yeZwtpDpQI21FEiC5mRSyRX4skvHX7gMESfghabdmRNXMUY34NFDmoYT
ZjO+GHqMK0HpqoDJBxZC0I6F2CcqklNPJM813sV150a6pOB4eArmLuciBQ1ErC6Ap0bBSTYBA1mV
7579Tl4EnF4RrOjw15oNoZ3wV7812KGx01Bjda8HY1OG8iIubHktuTd5wrHLnkA/70HjKCikBEue
OzuYjOYABHQ/nTr3WW/tnSAiMYmKZFzJnk0GJCBl7hmkykhcBSGlFnUip8WgvGHO6AZzgfhHk+iF
7RXzQijayn9DQtWGjg9h95kCFE7811Ha3HvBb77b/eswIZYe77jiUebjN2x4m4uaiWi0cYdX91Fm
xnZoG/Mcd05v1XaravDQXU+8KJX8C+xv5ji29akiEw1IIrCbfYRgnMXqu+m4NKZt/r/nQjnqsigL
cjVyHXxkDzyajZ7bn91ZqlJIaGwSzNyO55V0bzB/ICRlpqFFqBTbbeFfz2EY2Mm1wv7xOFFNiB5+
oZoi1SFnFNe88MmzF/idqnlT40VzOfM7jMJTOi4yUhIAl9FWOnClRJY1RCZkid8X4QzQZBIvq5tg
7rwLIL9p83K3sOmwwEpbgcrgjTxv7u+wYqcmvxexC1va3/nwUgG73jK7iYUv3duNdc2+e61ffM1o
S2SaDBZDQbMo5v/4C18VZo6hFnEjG//o77uGeMOg8m9917OPrLejPJH2hbfGJcbBheDL5ic0NnYC
XVNFAmMEjLDkJWIBvEDvAWa9QWDzWeddmZldlUelcuHlQrc9lmi5cueJlGIaqb399nTGXZXkasd+
g3k4f5RXwjeNLczn4z2DqW8QlWA2JCjt2huigMMRqPCovvlZ565ZSSBl2CxmErkcLH8/de/EoImC
F4IWi3MZuZv4T08tz5sqCuHiiEamgctTCEooWErWHMMZqfqtG/1v0owUHsyRA/qFtic/AP/aZWG2
N8+3Wef8GogG4tgLj2th5IsEYwhTsyKuwAd/ne+UYDdCiq7SEykxjPD08QQTtbUt+La4kI01RONq
INfay69KXd23A79BowsMNEhtEX9nY5Qe4Ngivx/d6r2A1gOL9VoY4GxToVDE8eluQxJ6I7IXR4Kv
d3/zrL2MajilWaNhF+BOj+tp0pkrPITptvgXmE5mOoWshCQHRGpXeBQPUPAJoy/3TABsghSXY8Zj
X5VwfGbn/RYvHy2A74htSDHO507Xi6gr7rIGl4/kHI6pmwtGUztlQ4njPprgjc8+YhTU+sXOx/1B
40o4SFIRA7FkzfDSobO66P0ftAZY6hust/4+7vYIEIm28Q8t8j9Ij1TFEk3Aajnj+51h9T9j3LQn
qct+4Y5abZMGsfv6YWOhk+vxrB8A6r8bkXoKui4Bm0CnrN6hoW5fWE11kiRBHY/ZWknnz9535+su
hOy9tgAPYnVPE4A2aK5IQplVDbCsY6VbxspSwo/VTwuu4+lNJ4MlQ7dQVul4KgT8fWUV/Rj/GLZY
h3UATbStziMxteINh3KvdAnjB2SqvFj5s40EdtUKrr7v2mOBvDflmEPYZONKeIaPcaZOBhHj+iAb
EGa4Shp9HubXKOxY1aHLBHh4SKOWTeSLhr0o88IkEOzrK919QI/vB+zDTAqEIPBwGZ0aRKRpTLWU
E3oDmo7MqcbseFSp1qgs6YHmsY2yBmuyonCHipEZCRJbP79HauvUbNY+qB9DNZx7GmdPygtA6z1F
a1QXLZdikU1H7KwCR2G7T2X7DX4sD1fP8s1W6CZae0KICyVz11ieRPw/BIOtSQEO3jqiEjw12ntq
hBHJuBxGSbCxh9ow6FbvyHLEb22vVuhBVMgfmfAB9itb3oz6eevYpnvo0uoNvZdAKk5pk0OoJ6NG
s1s07rnCdx+eDhKkweAOGRIuAtMOBSenEw5416QXQSO0OTrmOjDGRqKFCjfnvpEBkzyHBgVnB0Kr
NBWIpV1pGt57tZjaQgHzxovH4SQq2i5XCMFkTTNGSsxadA3Qj8vnUAIjLaVetF8MJy4jqz/PMJxi
7xB3xRYkIlQyWnl5mS9J47EZdPxsNqMC0T56ZM0leoQcdv7qoJjvi9rd/RXkIdpxABHNZrsWLZXM
efWoNKHzGg3e9UDxXmXeBksKwOc3+5JWRClzuwSNcpTaAD9aJZAXr5ZhFfJMksHFR2fA1rPGT7hr
D4APypPtTSHP+lz68wRzU3KvdP01sZi+BronMHKzYnFohxOj6O2h+euyl3LaNX4pRRKtyVCljIP+
KZjVI/3uVJ980Z2GkRutB65pO+ug+Zayq56l9A9LdbvNG/UcGaZO9ErWOLm2uz3kelu0vufIGzEV
UuhCwcVR38sd+kLqM1NfJWdhTLPkIGPovcWE3YqWrWOCCaDj/PkymKBMbG9cjb/9SHqOp8N8m7t4
guiWF7ZmKawVErCa+2cfpaboK6AI6Se0Wlc/dQziDb/7KomFsquF9P2+muzpbZjjawCAiQx1lOkk
yDGNHHtoF2BfuH+ZFNqeKcM0a5U+rZzkN9rNUQTiq6m5q1nRdVY1sXPzPgqAs/bCqfC0KwrVanVI
xFS4dn8byPCrp2HlOGwRjhgcDBfhdjSV1XTImrn4NSa275XGE0smHmvrnuEGdiJY/LhUZ9YaJZmg
YGpHoxAsJmkPec0nYAURgeYYEbqgGQIKv7akzoe03FIo9Xq6XHJC/sbLQLbZjTJzU1iM+qcO38xp
aXhM/n3iw+EiURcvWGY7ZSt2ggUHPllbQXAERkSFz9oIM1R8XUN7C9nq1xD7yFUU781uM8Wwv9l/
/q75yL2ZrST5lFRx2iXc0rdf7xOhuv34l6GZJW1T1x0bfUWPaytbEIJGG6O/JsOYXAKeuX+mKaD5
n4ZIqb2NMwUd0IE254bZvTa9eQ+8zLIP0S/rfPfrrnP1QPWOGrrvAmJvXpQPPxly3kmrpRl729bO
geAeAQWKLQQAlZR7rt2ZqWgV89xyCIB88QxUuLtIx0uM/QgwH3Ii20/RycW85UE5OhO8OyJpZtF8
FbWKYBIL58CoagrjkDDqETSBCm25ANAqOaLS7SQsOjMdnKMkb7iJoZYpMj4Jdn9Qrq2SAoLtpn51
9Zna9Yfpc0IuH3/PBWhXHfrmCdfBaioTJLlQfT0dHIdP4mebxoqbj0XWE4aiG0YpaBWC476kbeFI
PXQH6fmWmKGavgbPohiL4QmiknDehdwPkyz47FV+FlENsvKuBR/a5L1OQiK2MBamhD423Udk0maB
MUiobT3rjaDXPMqe1dIwQFyKMzNpCbLH9xgIxXDYRp4q9XfEr+4dInxvKS3c5FEBERipFblSiBjC
YPtdwOxdblfX5iEipjDyNKo7dlgNlEpCWFmbMFvz4zYY6jErxN0wrIQ3bMQKf1OTulh4YoNPZdrI
Wp1fk0ylvUbUqqHXx++ij44Ri5IC+KrC31mZUICmwrhL2uVpHdrkvjsEf7lKQwvUkJxCyuS/xIJ3
FYFkS0WabRrrHJXfe7oNjSEbvAfbbQ2WaZyfbk/xEbJoEFoupCdPUYcmpZ/xKhqSxxn/PHOHbplU
NopC3ZFZHrPbJ919ASflCLItelzHV4tFAKtDuP2wujjX8xQbJlIa6jduMHeTe+SPc/qGty8s/W2s
pbF8MxTsg4k5kYwotouRNHMt6CrPxSHL7JVrKCGDIQFROTsX+T8xe2V9D0FrYmdUV9Hos4lLjEb/
JeHy1GGVpjvIMilJ7mEdaLCZ3F+UTdWY/QgymHvV7zeel2LbiChfreG/6Svzwe770u7WGQpNInlg
ym9WP1bn5HpWAy30UcGedJapuSEhUH8HUPMV6tF3S7OGgYCsCJKC+HyOcKDTee5o82JzoMishmEG
PRAs4OnBx7oj3w+CkJrPqGyZGT7qO0coAp7Mu5QKbjZl1TZ0eHLXgNeelfi3268i3M6Ubb+ceNK/
uSU90YUPQVHPXOOvVpblzZSJBz+xKL6s8/W/wTumvQ0KtIa8CtdFnQBbOwegOVn+QYxkCAxeSH9V
Pb4nImLjDMth+R5xDACkQYgYG0Zg9Uf8byDFadnLo9v2HzZFFFkESpz51q6t0Hd7ngaDjPfPHLn7
ETaxw27E0gehFzbhcKhQ8G204B594bdIaEJ31CCaecJCuPikLYVgZUyqcxzXELYLNDe/mbUCjHEV
H5nRL8O/OT0N2uCyUDggQnA/FjC/vgzzFViHesJJPhwMwaDEHngR3UGedZJ9J533PrAfk8qJwM9D
bmN7XjEeS44VGimLgWrcBgDy4kCY6y41sP3V/xJxMkTZLlvEJv29gPL/kqzZyder0HOF3wNYd0uH
ju323S0ohq3Jr2cLHq+Bv2pWKB1yvkwWYcHeHIDP5kIxw4xyx7U9EuICuxsbcYXrSdI3StJJImox
hLpl6GqXOcaPxd9sncMtfdnZKjad8J2Hlt954WBBJijS6XWed8+Q/6V6c7r9kABBElcqihTg6rkj
3vAJqiIUCsC6PG/hpvIjVfaBeglNjg4qlJfcmjIz+6EKK76F93ZaEikbVxgjTS3ZZXOSzhoDcalw
oAQgXxsDDeU0Zsfcbnd64B+rFidaiHvpI4V4lyarBQcLVmfIgQGlFqypPDbf5l2SCXMHfAByJS+p
BLwHcYTwco0PmCb4dRw2acvunQfDTJ5y7gqxPmYlRaqW8zdNlhNirZHBuzmo1Lii4vF0CLVgoPwt
HVg7EJMLlCkUpAYTEQvR8TaR8eb2QmV/nUSbfqvhKt0gLIYuz449XaxIFbvA1Mn0NEKeMQKYE+p/
ybw67yZixC8v+7hMGg9qqY3dW6zI1JnQP02oAea7K+uzOx2crMDffevg9GiQfNf6WI5DGlR8Un5b
x2xGbGWHTFtoHxNK+tbXgauL3Fhr7bA2JBs7OTQ68ibF9w+S296FdAfa+oGTI9OJJ1426KaeOAxj
wYaGbCc+ZypKFWrU3S8bMb1/VZLHTYP0OUrPEByTmb8xqlNBfHMSMO9hRQUluLV9CRtiUcCOMsHV
My83UzxUbrwAlj9RNci2FqcQ0l9jHSCKChsB3hm/BF8TuVH2KoKJz+DxyKG6NwX963WRzqk8AJQM
ExTpi9MrgGIwi3CW4Cv5qMDs1cVamIs5qd13HES5JOFEuWXjf6c4NrDJADqxg27riXHjQ2V+aPlN
gjsTxMstLjVu2qAeZm0IH0NMwlRL1baHO/qqrZ2xdvQRWSJLT0HbFIGS79UmYMFI+twGVnr58d0d
rPGZXEJAgUgRJzzwJoA8seqIAmWl1vgpRzx9V3H3RJegQa26zk4Okzs2XlWwr0o+abu5ppSU1fCd
cThpahrjGyFXzn+wYr2p2x/h5vxr7iduIepTUSTCDxbPCX5S/0neLuMG1GsfF3CEc06nv4RzeIv1
qVvbXhqvGnChJpv3c1VwrhwcyAO9+LfeCC8oBDVr/bsjKpjguzFWqGxtMwAfNXf+IsiHe+NvDr7U
L94a0Gl3Vy9eJb1bhT4DbVmv+sqR8SYewYPDqJaB8o3w3mIu0CNtQwz+wEMkREJnKhY+dzpVKMqc
Guey7njISxggL5esSBiI7eBx498V7ydVgFKMZ++IngxstU2v7QggpqCOxJUGXsBZyXJDvVxfMNar
bysJYY23J8qQiGKxCyO1dic5qdrxeX/96c1FjygCBjmq2KXUFqhOUbf3zqKjwhF5U7f5RYQjg07h
dMG1Rm1xFX07pVLdnbb/DGuvoI8XocPKypqHv+p8HVSThSt9wTX106AsQfrcEmod+c6FmVubEGTP
brlSqLsr/9gQ2SmvDtwYoOH2Bpe4rmQdhD+EqMxSsQecP/0/tsaKeY4FZ6iQQbhYnZCstaOHsLrf
VZfIo7GBPVem7m1k69c0cnkIhdl7rPpjK/1r+Pua39eCGmSuvrauwzddnHN4Nh3G9pSc0fgfmzAa
TiUjKZuPSJy2FcKIGVvoxjE201RjA/cVnrOdlGLe0vGkxLIlBUEwcvPzEQbm8yaO5q6/JnoFMZ/a
VozhTmvn7fJ/8VjgqM6FjTfSktSImyk9k185LgCt1ba4DTkpvrQ5ggFJlQ4dv0Nz/gj3S2z9tN7p
bQKivRyDC2yS2uGPop2RKzORHbooN23uDPhQGW1jOP+y+qtkw+V6Y0hcPKgOTihjjQmZcgrat2u2
ytLEMvvhG1RtpSXmwKOLeJyeB7EmFUi1jpXzfbOXUnPNyBatfMfC5X0s+0Nap29sDRpd4ubg9kxK
nuLI2kaaAaTu+0NPCBahTQhBY1H/GaFr6s2dqEYLW2uyLG45GCt7oSRkLI8MnjdunqpifNx0DDIe
+hQILZSkb19nIevbAipx54QpsFr6e+f/iFpKWI3RNv9uybl727/INr5YVNcjCPSKNIty50Z53OTx
kbcRdn2MOdylkWJ4kmW91J7AdI9m22eAVTdgT7V/dcjgmw5TCocyZvdKYJTlemJf/sUH9l+qcr5J
YEOkno87T6Cq+DeYHga0PvELhR97M688S7MX/0OHazzeOZel2O7u8c6B5wZnG8KpGnl87gSPw4EI
oXOCCGGB7B2S3A2r1XGW/Rd053dJKrZmTqCQh75UrKsJmPFg3uyQIPe/fouQKSl8lnCNzzegOsk1
FGnxve70rbqTfO8UW+MNKoq8MoUT5h4u91UL4qvlClRLsYOpUYriKO+JccT13aWpZlg3/xp9Keej
wgTNFRzVH0Fy4PAD1nZDgFGzFxanrE0RunQn5D/f4kMa9NZl1k+ukulkVIq1NzaqXn60bF/Yr4Jw
UKiWH1i4YqJfxCjysHikK2UjktRTbZlAqTzhXpOoadrsYC4ciX9di4LqkTiD/NL9kJ+eNXXxF8QT
fNkM52gfgC5LYI0lpgOwGhK1kJ3YFYQKQkvNLT+KsEmzemJPzq9LVLsyjktMidF3uaLuGxQP50H5
G71KbyLTusWsex0VtnBRbPshatmo5RrKrxMkSPYbl1kAWNfH+eWby72+eyev+QoXJlcgADgEXzPC
vY1rIjb899svYdgW/6HnzggndMyssp4kyTxeXF0vlr3Jbb/r1MsQZ/WdCo+sNv9eeqIzCJibtlpM
FE/V37XiDqawmpavTqbfc/m/dD02jyun0o9wCIELkfWeSEWP5kITmGW8QBoIePk2IugplhO+dl7x
tVJSZN00WizTRoMsfjlbacF0f4NujEkFyKN4daou3cewD6sd0zpl3IaPlVX/RCjhqsimc5LyiPNC
EzFAcJLF/RFkKQ9si6cSA6cDspskC4NqUs28uYZqkYou7BGiXJ+eKaQM35ErxZlsZwCfoI1PBwMj
KqxQOOh2BsWyF73n7hkPkB45a9UjAJzFnVB5t8+BeespmtEjrLlK1V3BSxPmByDROx9z5S4PBjfD
glz0ha4m4/CrAdUpuQ3zLtyF6zGEfbHwNZylzrX2z5S19cnBFwP0v2A2jc31XNSxddBzuZAYzGF4
xQ6ct6QZ2uM5ra/lvE4e/+L2X4nsg+dblDtcEItZILXTtiavjrrWh8exXFFiM+Ck8x4ST5Z8BpL7
SWAcZylr2b2+h5Oi9qqKIrk1UFOsSuB9qg8atccARan0o1Pt2MWXwAedp8H3cCdb4d/Z/3qO3/Ea
2h0sbRX980GrT6afZCQmPxD7hFcGKL/Ob7TjCU+VdajRcDO/8VLFZg9w0rRjWUUU4dTG4POlclbL
OvI0HquyLrIl8ISQAOKM4/5EZc0lDGqX6sbP66hANwaiWq19WA8XlpzGFPdrZ5/3RccT4c7fVK0m
+Rj9tOe5h8YV/1EBLxOGYfH8n+zmJC8cIuwf/2egkE04G9mYj6O+363JVC07pc9Jn0ySUUZS8ajQ
Q63dgRH9cPDehLFSLw42yHXLW65lUx0vg18NtuYuDOeW8+KhSDp5/PmHCzx5mcuHE0PgnljMIiL3
wHzuA4s23yZdifnc/tdOsH24z5NpoafVmvQ63MukWKRxtp0sm9fN/bnv9PV43BKzzyFQLyBrJx5t
NxUPImdBetxn3Iy30u2HJiN0VHVqNnIkTW/ajGHdWcykKHWJ/1t0pK0YPLFvUx5ffVzcvWCZqBK+
067QTz6cyacHlYEQ/rgbz+F7t8cEFzk2/xq42hqa/r4BBOoeS/zdLao8rtsFlRfL7JJ8iL8SCQOr
D4dgWDAf7Qrtnx+8L+MlYPezSSPv1qnqy9UyV1YzKDpp4DV1Is8HU4MWMEhwmjrg6LOU9fTYO0kH
aL/1WB0HN1nCb0GaNWQgqPfo+ulEYSF2x576Dvd0uhyrQYeE8xitto2nQRwyRlZmtFQjutmySkiP
jzp6KYemOJd/fB7h0dzwylCZ/TfNeZCmoYo764KKboBopUCo+PEDSFU6n7Y/G+3OpEznMG8G3L7W
88r8YwBcgz9w9NAiua9dCARXRh/gbZ5M9H4maZ52hZjzYF42fe+nzYhIT9qfpYndB/wJyUx33Z8L
o3z03jPY0ZQ40+fpNqLJJ1FAa2xllpZw/TfEpD5oT6s/kFyIUVIM3L+tg3c3A0/hTJ6GEohHxTIH
NRTOdBYxkKDYsZioXcT9pbNVQFtXYnLudzh/85RmqUyplXRI/gy2GeAyeQ1qB4lXhvnYY4Tx7SXe
6hCJU8IuOd38YKqQGxAfQWs2yLCIv/DZSi7x/cBnD+kTlPhZ3QSJFOo79AxS7j5fc5lII3i0X9ke
4zM9Kd1q152J6JeUJU38F/ZQMcr/9j/niTPq5EZhy+4Rxtm2TjNSOAo9NUM5zKHHOxmg7SGE2iSW
PP3zoeCT6LFxuLwK2AAXh9ZxFAib/8eX1A/FxxVjtfO/w55KtpKKvLGaUrhh2+5B3j/pymtxN0Hh
iRR+JKXAc6heJBrRg6UKp3wCnlY/+M+lQMos6Rh53mhg7mr1WN4OC0OdJKTv0EMKgvx16+sE0VwO
41Wmw5KyKP7LfsAKy+gBL0EWmH3s5AWNQs5s7u4g/3dlbyEM2vKNBZaE7o/OC+WPLQqS9rirRJAp
jHHaxboNQC59UelPKigQqLbU15vSbWzpK4CKuRqmH+u3tlQjGFz//ZZR0tMCEo82iTvNyOTbHcz1
7DBqWZw9U1rLvDdozRwA+XKJkZk4DwF8J02wRlPlU4wmK5/XBKRZdT8v/nYPpE4s0uNsxan6UE6r
MZ2lTbY3dqXD7SYDVBTUgUWkgM4mXyOcqofBNeBsSruyS6NCQP4YgPAJDqml9ds1ho94YC49f/US
1B18Ok+hzYG4w1iqQov48d5jfJrvOZuy+z648xBDYEssqdu40pu8Xd77lfSbTpoCAGFhOmDtR1po
3Y+mRTecmR+kiWJRliD5b9Yym49oaIQjipTqhznyMAWpK+2ZYi3pWlcl6Y4A2loJzHaP30s2C4vi
LU4DyDK8MEfttLlfeeGM64FsBf5sqB0gB1FjMbuYjpWKHesw79pG4rg+hfjTyAK3D5zPHWjlIXqz
beAJq8ihIxkTRlqgmuIKhEhwlMgB5awTPYG6V+l5q9UdD2oi+vyWMjOItCwgJArtDvUSDiGJ8aRt
xy3yoy05BNrtFwhe4RoYI4J98hQYyOaBBI12PhbWREorE5jnuYYd/Qtk4t1v27IbEcvBo+Sp4Q8b
Rw74n1HVyl24YjJvt+hOdl6iJi2/nY5aUFRnJJNA53P6/wmevr2JlwNhg3/MIPRQwmYsoPbZV0dW
rgOkpATKGguZag96m+4TR63QE+CCv1qMnd8cgS9DzEfhNo8CW399mDo/1Fuz8xy0kg+w+zi6m+ul
BDns8Jpa4b8BvdbwlQv/tec3yaVpLvhq+chJSo5KdzuxcDj1TUli6MWasNcCNk56E60AB/MHVcU5
xv6b82YeqYQnSGnpPK6AmoOkCSQvbBCBadViVTTXT6ZPspSb1G4uUnz7gp6pVFRPSE77iUvorB7Q
VQCAQN3Pdrpk4zJZ/fg5eyLr3UGd8LItu6E0CzdiR+Jxnqb779feEMS9+gpjvA4K3z1GZJ/pRcAa
HoxONLMk8DgLmzWtve8eCX/+kEqqIiLrc+DJrVk9mYA5JQ8YCAbGIlrAdfOeaKcRusRZyeVAofXM
DdulmHpebjpTlRloPJg2VIW3klZBo2enKQLY7BCYtkNNtvU1ApukUt72rMpBE2DABexAdCJj6K0k
To0+VNYf7UvEqMOX/o5HM86x3HBdTJrPR98KMKk8jCtyAXWO9dBCSLgnl1eCjO+MbGovoPGqO/lG
Lgf6oO2moD9VdQtGqiZwmHYqmZjDswQXwoh/EQkEuOPiWHZcBHiOpV3KXoHojrT8YMV8LCc9uErf
1ylVIRwf3Y9Tsj86Y7q6556ZvcnTdGTXZ2cUZg/1kJwEr1YFmb/lzSo2Hw6WvX1U6+eIYfvP3GCd
ifhymoKNTKlIg0mmZJ8HcH1BtS0HGO6dIMCNSRiIHy0YEdoGaCbzIWYT3IVTuQczJCrdSwXd2IAW
+IHuNOm39IzQpiEmEC3Ck0c1189rH7SPaWadMFvX03SZqqWYX1ymr4e14TgUNPeatfQ09RPl4XSi
eenLgxiSGVbTSfaQck7SCG3gFDd82AUjepUWmv75IU6ufLjhklqn20bALvmfksFzmcBj5sPNEAgf
XqX1lULZ8SBqWosbkLUvtzVL6FCk8wm1E4y1RduU+l8ZgGP0xCu9owOBxr2WsPQADNRJc6CU0/sD
FWV4IdbchDUXfrs3HSFAOvgN9e11tiyyr1+LQsn/f2jf4F4wpI1PgU+ndvwYYAPatGYmO0WZosta
XhOPnM2k1Wp4WMSexMOQbrbbVx7TIxnsAL1feT6YaOAfdAnfV3OJOLrXfyPAcKlovLh4NgDKu+zD
S3C3UwnFxRyhETpVQFQ65BEGNxTHL/mSUpH9QuFb7QhjPEGrAT+/HHVx+SbrCG52CG17AgGOb1Ag
0V1gMTubkDVWPAJG6yeXzYFBI+HUzSJxmOxFz+Noenbxh1owZ3xvsEb5+cdoJ2fAJFAWDEpcMSzJ
o4av93d6WBCxAOBqVfLIdLe4cl7XGUwGdmkjxldJZ1U7msBrnUYG2yS8R5mkTN8uJi/HYqK6nYTS
jctbzjB1XtGk85FYkhIFxGlhtWL7k6nW1wCyXYyjPnNwYrOVvOs9ZinzELAgjyk9ayLf4/am2QLC
tuWk69LVZLL7zl69pfh3zwotXhHQMwiDTIrvmZKTe6GC2bFD7itD5Ce9OveZHQ9uBteFeBnna1RR
LZbJPv5ZkiXtt7MhLuf6C7FSRegEHRpV24E3+RE0UUWXDOyvEFqfk7t6KYShh212FqZMFcyK4BcU
xr8I6w8C/iSt9SXTerCq+9QhxKOmccdFVn8SdLjaAgdRH2EgBiI06pWGGBr1c/5n2byNiE5spH0e
xIxb1aHFV6xQCli37Zh9TNiOAAYDeRTN8OUXa1RkPhZm/mr1J2WIRfIMCemyyc84z+dU/hdellHR
rUGKpzbdcMNT8LRWWYvdElJ6IlfQzPlRpKfoO6isAA7R1Lnb2z12NM0eou6wQBaOYhYGGg68h8EH
vTdJJ2Sp8xe8nWCoV8Bhjs+bJ1sSNpHfDq6D81sozfsMADAlYGPYPwk+p8rTaPkJA0x69EhWtOCJ
kFC0bK7ITFu9BbszhSLfZbDizxrjsN5Uu03YgPeWNevUbft9z2qFJzUhzJaVW0le7K1nFb3atPlt
ZxvSX1DRJmAiD0Exyg1aYcsmW+ItmbElGW1mgNs7ujCqgKQO7Q8smutz4nDGd08hze/BlOp1Wv/o
dHWAXp760o47evT1ZSZi61YKjdHdnqPa92XtAayAg8vIH5dxtVufXTymc5n/9o+7RfGCe4RXGPYk
GnTL3W4t8vWXqVrrL0AV5BECIEXiOBqM1f1uvmWbEBEXMYc44LvV7xOF6QTgV2nZOMbM3S4jBnsE
Z1h/7/lZavJKWH4mhlzOHcim6gXA8m+2eEFy99tefHVXzzHW23HPT0Ku02n++tlbVVtPgR9SuFyt
3+LOQmZlsmtZp/zEwoJji7o0KREPg1yJnCr0f/hPkn8z9nykqNZ82o5ntG4JTIXsW/ZdqRxk30ux
KVbGPSNwGfZOCqaERUrIAIJjMsqZsxsWgz0hcpFxqaYpm5lpHF+vV8EElDobD7IOYxakIkc75tck
ZQwMSb6FZRu10MuPTAXwoSdP2L6TBb4ucrkKdnJhnpGycq8FjL8c8BF2aKiBsbBNxlIVyup02LMo
PMzYJS8i2zvowGJjEiictBO1+UVkNAav8FU3J/y54tQUiS5B9DAgL/Q776OhyJ2w8216MpW7b8yn
zVdVJilVzMIR/QtlAzjqz/F7wljhmzV8kf8xb/m5HCDrNI9ZsY6SQPhOf4SbGiPIDnt+AjL81NUW
AZ2uds9prlwKYP4Oo20wLby6ugLYlobHeaRim8x5hqnFzpGVqDKC6sLQ0wkmYhtJCsUcMv4lpgk2
H+9xiuR7Ka+qADgl/icTcKfeOr9V1plgp18ck5+NzhfP8eaeY7GsmoKrCSc79lI/N3Re4bYCyqh3
Q0zW0YtjoI9pCoqsh4L+Q2sR7Aes9wS4hfeBLO4z0cvl6+PUaG2kPSBFt91LOvUvzZ+TMwZrwSJS
xKW8jWTdO+83KxaAZ14IQXqrbCRIa3h2YOOG3t5G9uxQs3ZpwA5NqjidFfym60AR5T02XS5T+ZxI
rEfz7LoL7fxb0DyOUOWogoQKFmHx9d6PSmyj2naYoctyERiuWp90tB71dd/G6JtfZ+gnMsX6Nycy
2CU0/wWnQxuJa2py3jLdq8ITZOMr0Nsin59rvH4tluEMmfR7Gp+IywwFSGrcnylDwNB1WtzGAht+
r4Ff59Ch30MWqRnk6uWAq/BD/m/FS7/zU6Q54eciZKNIIQD4E6h2NApPU00a4+pB9x0xzBGZ55Yp
Ajm7469rW6RKRb70Eikx/bYqds33uA/beC6f7AtHapHFkgv/7S5tpjcl8vClh9JSVyTxRwLM7zrc
iPvJPHt6fgYuvwZ2B5788AJukjNaVMiGrqr9zszEysKnmu0+AwotX+4tg22UNYp3pgLSe8DV5jOV
5Thh2Uyeq+GOkSe91IvI1SmAMSjNwoncgSt8JH2MY2YAfAOi/2c1u0BVTB6Fr9fZPhW8t7RGebm4
zgYEFmS/ADcRaXzFTfd754SG6Gy6iVORvCYCumEXhpL5Au0pBIOs2dbKfzo/wtPH8HXnW9HMA8NV
3UTx4pXYzsphyuKDxT//SLNfYm7BzRJ39z1Hph+QnUzPuem+M4X1frUw7mfR6vCZkubq3l8EFx3P
r/C5HBe+qJGu9l7NbsQI7QMIhr0efzzxtcrMOtKiKPic9kXcDoUTRLtKg5JBg1eKBiE0jDITVhWA
zCTwTzJ05nKKu5c9S1pNdImZT+a5HQmZryuQwLVHCCcQPXo3/4RBpt/DRamAQTZMVP/Tar3VRWq8
UREPVNOonLRxWnWXqAW0nPYR1zlL3UwU25PSN405/EVTkgXcHrfR2GHZcJOr11P2PyTmb4/1/7NZ
3luQcSl24a7ophT7c9kbx2dr4NappdAzDtc/2DF1dmQ4XE8kpQLXYJ2Kwk+sHSYQGto5/zAAuw5w
JTZ7U7cYTNevr15rAtcnamcp/7Dqvpop4+smyHMs1mOMuaJBqONUqfIUOaSGB0NmqAVhHBPAD5z2
fY/6mjHyjQo6RpBEzAW+7U4NzbMGXtaF62OrglC+6rUQnrrHY3XP0uTjMZQg5eeXEWf8Bz3h9GCe
y8T1EkHXt9bAlv/LBupPE2hvEqXvSuRtShqU+IyOnl5Nk8DI08x/6+oM1zifTf92mFgUFrosQ0XI
SDxjmvhvOxs2PckZK3VPzWBvZN9MAl/cfUCdhI0ZCCJ7oBkFo4lfIXM5JpvUgsx5hx3AaIl7u6UT
zexvSYkobr3Qgietcgd0PZ533hWbw2JPeBRP3InShjbOWr/E/QiAfMx6xbzC/0TSUjBp8J6j3tmV
7ijynKpOJ0bZ/5iuy2P9YqOHJcmP3x4QopET184vY9UZzBSHrhsCJ22tm4oN3gFFktRXKb9WxYgE
PjI4ZcrdwepPFnfuRKWUIWPWfY0kbPIIowQNJeSUDX8apgZvNSZcpf9qZf4ibQ8hKfbc0U0QVoyu
/+57rLSJJPpV25C+uXQHRhEDVctUMRjv+jgWP6xi/nJd+OrFZ0ds4WS5iyaosdh/VcE70gwLqNko
SUSbrJdL5FRh+IT8F2/GNcbWv8Gm1r/mF1vuNcx131Z/e7wbKQLyxd8KQidlrC8vfXeiMz0RNB/V
UgleDagAIlTzAft5ZYAUnNXwYjpPxUFEYomSGTJker3mRLef3QmZogjotqOwxffo4I203XViE0g0
savbF742JjbxXltr6KwpXcsPRAeZkUZR0AwfeOzFPqLhobRM92WkYuCGOhQUqpUZNP1p+RLlQCT4
shd/Wv81sQdCjTH1xOOQsC3w0D8IARFsRkyreLsgacbTMSVI6SuSyrxXtgE4m65fMtQhej/JYAJO
GS8Sdq1hcMOnvHNFntVMY1ZSRVvVjx6h5xxDUJWjDKzoruH4P1n78oZuN4k0EimVu0xYafkT+W6w
FvCP3V0JWKU38MGK7q51TrES1DYFqyZzQv9zrtoJlOy1rRAKIqgKhF4y7ogHYRwkPvYuTfgsUG5D
dj17DkgRQ+tW5sIsMRWQKdB12yRZAYKMNtdBHfKHl8UmEgl4ZxLM5qiT82oBetrwLdNdhI6lTD85
8z/6TW1bmKEZBDDJ2FRGx5LexVrljbedvGAO57qRjUz++lAdU0afSkQLIUiTMdXMxir9ahIwdLtk
1EzQyWeDTATXGfUP2+snnSvbNKzIdgGORQNNb0JyASFNYn4L2iqFe0EB6JI2SbXryq/f2DmANdNh
S8err+VV/qc2kV4zTUjptiwz4HbC0dhf8mHdVuwho0W2PraiC8GuXC/G3MmKeYjJxPNNeYDXzdEq
dgVcS8xX6bFmRzi7LQ7DjeYMcQUxPsLP8Fuf6dhbrblcEG72/Z68iKoee75azhRl8aOXR6GL7H4u
5bc3ku7qtFZv8UNZsxs6rFw3hm6qfl3MEkb1nh4EYTsY2LOznrQMvoQm3rNFjrRgPELsRzMzhnJT
ye6YXZzehmXUlUkHqE00iJquvV+1QfRtElRSc+wVKiEROWHv7awejH4RFAy4JFJCFjbKLNRdmkMB
ilt/4UKMv6CycFG5K1AjKw4uWHaEBhKXXEFNNPn+MAzxu7GkFFBEsrrmlFebPV0Zq0Nzl9GPWvrT
cX76SJJHbUfgQEn8OMjc42Liblh28MJO5ZNfHQVkieMLf6LBQVkzrHG0Ref04002+bv8zUUNi0FV
9uRcVW82DCCeonr4EkH5A+QwNpTq4Rde266QKOqKVGtLjR0Fter1qTGG5I9lyCgIbKep96hFbODj
UJy3xYYCEFetAaiI8c769iWi1Q3GYaPYxjGs0pCfAaMZdI+g/fs8Zkgons2GYcSluWGCo6Qi6IVI
Ibd111RRSWI1+BiTCWcU+fnvB07wiGOmdQ9uupcEBUvQ5+SYcgAWRqjs5kPNJ4Mt1ysWfcviBp7H
bc6O6Sczvf1XDQgbor6FY54GRGi4iY6FsG6x19CZeiZrtyjkp2RNzxEc83LTQ/O3weqXB6mC6hje
PNSNaHU1odP0GNXdSLSo7tIepIx1JMo5ng+LthNbbiXwyJtV3euO0x3Veaj7PwunMDU7baXe89JD
7M5/6IvZLOhQQ3IgsKcS/FKpPsLUwlYYTDLM2dyyR4Etl+5p5DsoqrfkoeNyMrjgpciQHEwZ9pzZ
EV5Hgwb+J2G+XNoPRx9DpUlxN1xgMX6XVvlf0Rzt9zEZppLj/ecOCYXShJcJMuAnRn7u9Qokfal0
cFLg9J3w7GV8kjAlJiD20NpiAfnacnK8JCPGgUNKWkfdQNHyKqKGnQtF2OVhc7ylTBjnjKLoiPH8
8Dbn7zc7KlqqSaCMVbVNavoV5XfD9kS2t8HECG7wx0n/kgjRioood9ihAbPwxEM5k+PuA2mldhQH
L9ttfR3JmL0ky4uXN4mmtHjUWcpQrAsGt4CpOnJHCM1F4ykqSNCeXC7pdSBoZDEufWbtoE95wL47
9kcl2dKLdDkwOD230gsNQt6F7dNTrCaK8dTZY/4qtmVidAnF56uQPqnKKbB99yjJZiPET54isMpf
BcMFO0RRvulES02/G/G4I1rEaDqIecr5Ujf+x7GnjPiU0LvgDKwASyGwiplt0AeR77ORrOpnns3X
BHXJvWge+/3ZFVURaassW4ziFz7BhGWzCpMlUamR/nBoL8Q4KYGCUcHxPo76Ldz2RXbn3aagUj/B
DWQfQ8dppMAMXoQZXkC3sc+nmvs+TGrAlvh38TfacwnvicsU5SC60h67J/5IZ0VUGYBufZlllzx/
RqDIPdrBaMdNbAd82I2BD0MTbo1al6o06N5DDolH99Z711bDEydW/yDopHNWvL+7xn5KOqKUTthe
8bTYebk7xh00/MUPycSGw2aKmhCYA+bUPWMMg33JBvNe4yTkQ0H9poqmbMIkEbzH05dJmbl30ipX
waGTXOYQpWLrudK4FCUgEc6wdjxy/KdOMDSTHaWPteSv61lVhTEbOj4MM3GLiC5Q7CnEnc11fG9s
FJC42o+vuBIvtJRyHp5A64aykRKyNfuQL2I/U9WsI+FlUyqjKbrds7XakC8dIyhoVxWbQiU6HGnt
gix1un5Om1kT8ELU5+8Z9KXs7DYo6sJIk/FtXIu3yz6Sjo+qOPj1XM8ZrsJAZ2wigQOvZ8vz78nV
0VFHZlDNYFsULDugNJTIuZ80goYIhg7oekWPqMxoWzlDyjaiYgf1isNp+e22mKuT+qDbwWe0YuNO
m56wnVoFKJdQsfCeaJpUTz4+E9R3Z0MuDBc4G+Z0OXflb/cL5Ewh7Onl9r5DtTgMoPVBFiiMAEop
vU7qICapEZudpwKYsGI+66xu5dMHTg6gX+U+RajpptqDDcXo6eORW0hp715atfTlCpcfToSPR491
mrwgMdLk11hU8+7zb+al9op48QOrkHErMY31aAJl9Mjc83n17RY+XS3LkbsNbmuBO6jWJlxnjjZz
+JACVZND6J6jhggNh9alJ1CGRPPHsb5NVCV+cwVjwyGa0vM/K8HF4tQa3VRGDRilDYFPu6CVbTtU
hO0eU6h28bm84FS3sqt63ERbJWp1yNEjiP3eZxwOh4UAC5U5gwtw3m9lj+DWnz4kbOKKCifrZVVN
L6037cb8uwKzw5ryTj5x/zmaOhohhbX2ZSMf0yP4VSl6KY9WzPRFl9BE3B1pBm+b83W7X6w4IHNl
fec9uC7eqSKHkq8dn9AXOEAD7sqxtGRrGRIDu9k0bJVGNLyXIYhTw74BRv1LBiNwJ2WDq1/tp5Xq
XcmCQRDRNVp3kIKJ0xksasMMwJ/5st3PbxWlMzq3dWKBpEmhdA/Vwp01AdB4aNmot9DmetnVwwsY
XlV2oy4B1OJDVAAElMXBWXWpC7NEDebjKDO1GiJ+F9cofWvibSmhZ7f4Im7Xa/9QufXLk5583gxH
E9MIyOPCqlij0BfPDvmCIzyTHSBLjuq8yIUWL79VJwOHg3rfISZYtaZ7bnM7zaWFIBp38fP2/P/H
UVwbDi9Z3gZcKFUlelcErKB2oNc4adqAj6Y3cFDuVzo1mjkaB2WU6Wg79MzPGTf3/cFeGNojOq9z
OPVAVyzQ9Yw3qdpu5/5ZfP6Y5ZseGxk5pKannMUqiXpFoiJa1+srK8HLOv/0U3zwodhSe0KD7zYf
WYXGY4zsEdrajDNW9CNO/4A5wb8YkfZHJmjJaXwizVNd12OAK2fc4j/zXq+ciFFWAuURF+xNWZ3K
rip9bv8+/mDeIi1MH9a8qDP1ileWUxNhFzW9VMLW9EA0F95wPYlNTsm6DQmyCJK0qaYSw6b4wKfn
MTYDA8JxVveIxWSt1ANubpcC4o+ZKJTsfdU0wf/BYigGEuD4oUg6UAj5BpZE6ptEN54rJ7FcpB2R
6gxtShVp1yUt/Nbw/TPjY7Re6vz3boITud3ue8hpgVf2vjnhjDJ/s/OF/Ey2hwm56LcAkLKk/QbH
oh8WPHIPdKqxVb8lVRKqZGMfbBMXqCdE1DSIfAPPqs1j9JTclVpfuoRA6S2t+vh/OsQ4hbUD+uL8
x9OA48S8S+ShA7Fsb7AfPl2AUk5koV3nmApoW5DWgPkaLUKZd7VGDZVuSU3cFSQtLhmGXet5oPrf
s3a7lEDYPASlyYz1coXqmHmwVQUhK8AcEMx08rJ9vPwnXAeF+NxH/efIldpL1rtRdhbQZgEMLZQe
iN3E9m4t0Zbqc3/Fxc0JgBtTap3fRZ8eQ8dNV2puUAUSGtvNvimDJu+64qZhjy69lFdym08/h6BB
osrXB4f5klZUaxZaoCS47i6OU40xHBO3LH/nvks98FAfXftKZy9P2bI0w52hxePyV/ZRPmfa0DZg
Tz96CiUqYedOztexsn3KZ7ChS8BR3gt0XvPKFed+R9RXFF6eIdv6gqJ3Vp78z2CYNKG3w4RlRO7t
1KptRnIbrLIFiFHwHU4HIP2MsTznx8V5R3+UtWuQ2CwGP9kvenoViy46UtIxdt5Y6xitwiPclF6K
vfqXV1jQHWRBznPBhHAKJi63bhwwh4oM4v4Yf2o2L3gPd5rdh1bcbtThhkNYyLRd+49374ak1MbT
QgUX8+i0Be8Z7JHJfQD7xydxU0TqWRKJRMzMJ72ldOoOz91OLVQ2XjSR8yQlBZSIna/QAkkTmlmV
QkudJsjWtmALd6wHGMftD1n/s7ogdc1d6vDF+bT3FbgjIhRkrFh9rDOZRdehflhIOlpXho+GXZXl
OxSgXP+BbBmllyp3C6+MXDcyJNFOHmOQI3ETi2VFsQ+pe7noN1ktIzFcZATBcJ7cxlvNWBIJ9clt
R3py431eXGkCdCKbYkdEXwOZKTgmsdhlZ/+mOLIqIBRJIqDqsJQrXI39PvxNxk0dSWFvfxREXoV9
0Md1sIz8KxviT4ef+ujRNUfK6modKIrZh/f/y1XxorrEzngpB1KKEbmxEjL60VY56m7eDRbJKusC
7r1xWcrgMKG/+LUnaI3wR/9dvjKr+LJ2UNh5B7AExUxK+JDHM2dp8laO9bz7djvuXEQK7QlU1k+q
eaPDdFXQMI32RoYa7yyDwJnL9XiC6z8qWsJU4pHwNjx/vesoWhXPkVKxYay4qdqPt4kZt6xzY/7v
BoraBGI49vQogfU7KhEBcUdH11fnXhzaelumaxW6ZbrvGB2m81aXRdLUATZaUWPTaJFGrhN7D8bb
VDHXgBPOB5WyzA6KPkVtX3wPWtY0IHkYVFwyRlLBue0dqaZEfCdcZZcfi10ZKolT8ndXuFf01VHs
Q/OYX0uKz80VJIfzMRq//4g4SfLh+oTaj2gElPJpLiNZVheMR/wNl4/jPqIFyYy0duyXkrdV3icM
mu5I2c/2crYmfPPv9qeP5r23B0txZDZSKIoNNPsuBoZ03WctPbxtmipb/KHOKuPeeYvUxhUtqo1v
d73CVxMkjQ5SleQpwzWxp9y1WyzcTZDqQYE2CEnPwUOz4D8ok/uFbit9P9qgfu8EDtUu9BISQRH/
Id1U0erT4hha68XS6bW8f2juy6Z5yCJj0Ms/PhpbhX6TVrqBFGoxTGOZtfVxaAsUvpc3cgxSFM4q
18rYzrE88JP1x2JnCeD+6aW0Ex89K7+4H65gPg+osA87bYzz9ziQqnAZ4ZT52On9idn6+4cFWcWf
Zn3b4SqDWiDsiwphLivXbGUTb5AV6Xn5OANbEVXH6ReAMDX20r+tiQCM30sAt/VVc6ya3LvIrXq5
ZZoClNJ8cIehaMrj0ruF4/2tqqbuTgGjOca4oVAXcuCegittFfHXKNmNdFywterMEd0NuGs8wcbL
mpwDHoIqHyc1ppgN8Mb4YdQC+K2v8gM4eghaRJUOVEhX3Tntj1wHtx3Q5fhcC1Loh5xSejJDNzef
zIvnSnpj7lwnJxcCxugxGhKhDp6cvnKxLiiJBuTBYcsuKVd9J5Vn10xF8/2beVhn131szYMFFjBT
dL2y7hTWN2YUV3wD/AhKrLNKoKAsKRkAlENDTEwxxVYtWAXXKySmmDFew1nWbfhK4JKgUBGrZJ+w
cb7I3Kd1NZHxOGsgqvkD8av+KP4Ln40vlTtH0w42x0vJS95noxNtHRZ4iVmmF8WBLF/kEqR07QMx
U7jg3AtN6flOgAeJYjMlEHOQdO4V288Pc/Zm0kanJsbZ7O5csh9QiQ4R0QrNfrGieEmopPpS9S7C
amMYh5k7PtBleexBhJaNODrNy/3r6lZJqhHMK4vn49GICz0U2qw1bcnr06WMCibwwU2HUXxqxlkN
AZsIzehpQ7x6L5izi62umZDBCcC6bhpTFVWo5bKMXkIJwojk3YIKOd12k6PFY22nKQM6vVVH0OgS
WT1GF0R2VJCwn1R+mno/fPoTjFvl8uXHs5wqaslj69WPwGU5z+A8AGZi7rzarP+ahX6aay3sWzM6
ekfm85WLeI5W7tdv+DvJiRAevLsg/rbW3J/TgiLJHkiSlMIx7zP2i4FI6ot34+oPOwq7dzTh8wqf
IcwLbsJ5I9g+kEYUBS/oxd4yc+WvYJqns8DCakyjQGQSmp5J+zUtzBgyIxAdj6h0wDv20CWTuNBV
LUEy1e3RZgJKgC+6JLkuemeGQqwvgHeodOjoM/HaX4NGRPr7FLCddqycpMDph4T4RR5ODSkDKcPX
SLF9RKmdNX/zl2nziAzi43CXKuBRLDHBFj8VufPlcg0AdHolWUnT+6kzGU2nwnHb8qXo7u6Fd+WH
v/wFkpMTVbpJCI66J+YhKTPtTrFwX6JI+Fr+JDiolMAopf3bJIOIk6IB3218Lt2yedV/b/1g7439
howJ14+5Q0ZlvMYgCZw5KoGtgflmbrWlCp/0cXYvrEwqN0st/5gJa623/wqIxCPurizVwSqxAPcm
chH2rwWMVdeUgfJZn5SxB/GXOMT0FSFsQ6HFqQ9HpX5sB7UJgO1yILjDuALghp6a5FmI4fuBGM3s
UisMxscBjFkVI8yrMS93qKbMi5aKbFZtiZGQOHQJUVINtmjnm0CgVhS0CJJ658u9fUakU+4uHMSG
De+6TrMU8HLtIRSE1vjsNWrl0tdll2eJthuqAsHL/M8In9+f24DgIJ8STx4vGCG6bAsBRyfZjXxu
HXpaYPH4nszgg8Hqs8YbTNvdxACH886VZb20/SkjPi5ZZSioNX9fFLygzhpcZonNVMqr2EYDOEKd
FuasoAdx7ngXOMHE4rcqSqelSm0I0Kyuhg96AnrlKGyvo4hhwczWCuYfOor61mdqMni7vrk9qwZ7
umnbIWmJXB1oVkr8/zIx+34ap+XAdwwrYgy0ydvx5dVMpn2KTxHqPO+tNNFFAyCV5vmRnd4a+xN3
lb/CoUrv7RQFeeHXFI37fZPhFJAdXEO6YWPtp7w6BOBiHbsLqN9r89ozVeaXoBVSwS/+dPysytLI
iNmv9FA2AQAxHNoEhcefkgH8sgtamC66T+vKn4B5LBXrf9ovSBZyElH4SQJ1Unr5jvN/lYaRp1ns
+X9PepG3hPr57ESyWNs6NYlB6ya4qfH3Txa/UVNpFl8rDPlLpq3owgfpzI3oyvp6tt7l2IBhP/Gt
n5MjUlvA+A6DrKdx8vmOhpuNXq9DoPtoOkACVOKwxN48tYbDq8fo0dFb9oG/BJAY4bSr6Z7vtKKf
r3c4FJwhBxoRm1QHL0syo2OyuyMP5UZaikosV6+r/2IIVEm57JUOLL/anVcxSUSotyo9gPYcLn1P
SrKPRH7Dg1ZRU9+X2GxgiL3hzTWdEWmurivCT5pL4lRsIr506cwx5a+vsjNKbBXZIGKWdDpd5a4Z
am6NDoHF+P5wdsD78BJXS/2NP+N1Lj7g/wJK7NRp/3OdK0NEhQnzOshRAGIW05+hpnKxb9IBx0WW
+Cnx1wz7+nay2cADgpVT5Y2EiOX3WOenKknQt3rZTVORk7jNIAolo/5nGNoEF8Y0+E1kS7cmtpL2
NBOSAk3+ID2L4PxTDO6LIV7HLRwm8tj9Tk2cFo58TpFrnpGp7XYhHlk0Geh6OSwjBXZvm4jW++JJ
WEUMJI3SRE2yYird/acn4+6C0UScGtdtQ5/5fbBKlFYM41f3OtGKLq44+HbEM5dgS8RJ1r5W1hRO
rj1WugpZlw4652rBVwHGzSYR0Oq/7cvJacDUCcvisyMETgxcEtUS90UQPCU5/HSNpmMD0M1yIA7G
PiptjD23h3MYhNzuf0K7Qvl6Igw/u39pa/fhgqJo1nqCZfe2CMXdjTLxpwayuy8kVNe+GoGlXBqs
Fe2yrdIhbbHmDtMXVu3CY5/4Tt+HGDfTLIMkfhXrLrfsy3gmBvJHF35Vxi0vz2YMuGSvXSyiOFs/
4q9vgM/Ry15V1uYgD/vqT7wno07ifPDpTQrzew0XW/jCfVj2f9ux5Z2VCKKRh+7ApsJRcZizX1LH
QvijeH3FBeBTkksiHQJ23VL7JnNAcMGUviy06BEFBDkYD0HcsvIDkoO/7cjgi1WUB5eBu0q7YugZ
64TPnxshLm+C5RnDETCSGMgQ+h0qu9rPVRslLvz2JnMf+zwEI7BR9EoP2JJgIFQQqEk3+NUr0DRi
5aPic86WAa2Y3mjxxa3bz1YjVCXbGvIcpFTrQXLO60kexAuvGqLdu1qRHe6j2YePcev6ILdM7vY4
p8iEyyNcGyo3uGLOnZub31EYcagLqCslNFz8v9l52skb16Udo7rxcR61Ik148F43M3GZi60cn9n0
sg5DEmDZSZPCCdOcenXxFVVjeXQIP7Mqhxf9FuindPSJInmZczS9RcjnRcgj1vncqTOth/dsJhlr
N7z+4SdvGsQeqxTqlZCa1c8ujymMx2VbFuDGcRw7Oek423aYVpN/YT6kMGZY6Utlv64pjVR293Pr
maBKLUUsl2Q8p83+us+hGGRPOYI8Nwgn5gD2Z6t3C1jgIctMHBJbfhpAQOiJNwFJck9Sxdln2mXQ
raVTkrj+OeRV5oUTKIpnp96n4rABGd2mBNWLX/bLdoA03JMi9s5sHyxX8nZF7E5md3v9wZI7uNgT
qTyFg+JfrBsoZgoOQtaBm0sUgLUWhcun6YyB6ZmkOus9LUX75E5ecUwblcVCp+YjmoctYM9fzY64
zv/IMVHViDGgtw3xXKBuPz1D5ZzVz9Bce7a2iXtJW6yoZdZ+SbGn88f55a4O+vv39YBiTbFW5L8x
wW1eNO9fZiiwbTp7JlWT/cb3w6hiK3UGs78gFG7OukDsbuXeuCt1I5hrV6NRnaxFrWBzJGqhIxmW
5PmGo1o6t4plLrQk3C6tvjEkDYFrI1D9R8REnaLmgs2s2dPtwJqmOBDL4Xzri+wtgv292AZkJN7p
EYliUcZT5OJ2d336CqiW/at45HnqYGEMKddvAjyYXU+5ty4Lul2EqK6zXKYiiY1t0Q4xpGKJDCmh
prEQ9Ef1ZBBSOu+8GCoxz/hj++4rjqAN2pSu0IJPn3NYaxUdx2y/x0OTffOAwUkPtmwidwl8zpfY
xTOsQWtJ9M9ZPg85WJagtY4zOhangIic5ZTDehMFEgjSOhK9/yh3vSYE8lBb2kyUKOHNahimWjCm
/gXYwlwz/1Yp+BPx3g7VagJIhBX7h4d1kr0AcstL2mgHQpLHPjat13mz5I+CSNqRA/P0dh8xSZti
o7qZj5VjJu7mR6RWMfOfPZriyVtjjZRelt+asfrD8qXwOCWUqNp0DgVtegu99CmJ7Y9hHISten4s
fdv5TyGVspTXS25GLXRZoGcbIPVnboo6EQOQwEFfqgGkm1xMekItT+u5Cv+TBUB8nFACqBN4NPja
IOyQqTi9QX5lzpfYmtmSLCy0SpFZhqz9rI43z/u1y3IIHPYV4ht4QtTLtCh9hwj9GGhDqdxRn3Jo
BSN49vn8uwyPlRJkJfqBjrAChahcQjnUKxAuERcdaUe2Nf2Hr8SY6tz8kDIN6p3QB/aZqK7rGdAQ
eSSTWD7nNE6NaEPkyW8MxlB+cT1ID7chXVkmaL+7Vd2Z+IPey7ns8ALC7EV4wuiTjDQASKOQWQdq
ZPXBR8EOaEh+MneOt8A4Q7J7T2HQeriZqxHf32lsV8IB/miMeuvxvQad+JUxryQGnzoiua/QHp7o
em+kI2tC2i2gI5DrMVBJfPSIa+swD4P+h/ccj/r1KMuS2aGOfRETD4xECUq9YXjc/J85ytM1C49p
kS60D6YTdZg1kWvnhW8lF+jnn3j+FiWwsTMLuUtv4ClE4Wg4+CCg1ZhaVS6kchtIuMdxDzGQLbac
D3BYt8+fm9P7VfkaS4GVVjvtGeJ3zEjvYplOn6yE569PVGa7cLAtsYpFALdfHr7ZxtsfKwlNq0v4
Y8Qtj0k5Zvpvy5WGFI10a5TMewlO5X/IIJHXaP6mGV5fp4da88hBRcxzPpT0CcrssII+GaXJkIC+
tkFuNbQSlUrV2Cy/bLy/sJJXjS8gxJf6R8k3OgJBAwPOBeYvPW0NS3/u6g8m/x86UpAPU2XLIdG4
ierC3vanhUkYbQlzKg5m0AIkFUOkTTkqawxBu4SvriZWvKMOUxpCc56u3gLCxMz4Si61+e6xFiUg
Yrl1SyKB7wBDH73Fe7PU5at7dkr2dJRbQN0nnzqevZJ051ne0EG8AdEMPxvhL6Gwhfyecn8xpQUO
EpKtGn/LnZS4/FnG9ETxjBiO/Vyip3jKYWDVJ3Uzqd1OxcdSaCI/sbFHQVmXAOmCoQNRITjPnpRZ
ZFb6Aqm4vrL68Ps1Z4+492xVLhbgF8AWNRiV1q5n94YBKxIZqs8GFmMIabIerj665UK32y+RY8bs
pZQVeNZfYjXpzyqi+/IRmOVEEmTSMLOldc6/iQ9VtSYJi3ASsevf5Kr4iXBfBsPjAVcjVaPGzB9s
c1Yr884kYpAc4nS+eEsnJBwORdzzrHB0jDRByx1gmpsiP3jmj/6IevYng87Kg+Gs5zO/n+m+QNqT
FSh0gqZUmJFNzSEWVPpAYbFxcMMJauq8qbraGhY0tn0Y4NqcwRazXk73Kr6gxmzT4/X+sYvs8MjH
d11EFVVMwl0IttwHhlYlSgXMhS1NIKSA9LhXSkbhheRpwL51xho8p41DzJCzckvjSLVJ2hiUm8U/
xhZF+aJpLuoIhhALS507QxGlbrLoL5ihk6T/pJTqAMSaXKoAWKGf/tE9EGhW+M7JXei+YtV2Qkt4
kwOxrT//VZhs8/kTC7pW7X06BQSjlkVD7ZfgWoTlswcyJS16GQbN9e/cD5u5HGCfwpBLA920e2Vn
BBPMXa8sY903g1eVOhrWNR/UDnFVaSPGLUSQEO8KCY84iO1aoHW2j4W8+KQwFaIVF66RH/odSA8u
Xklmq+0ea8AHodXbONkXzDNJ/DR2WDcuUbXem0BJ/FEom6GupcJR5B7UpIikDh5LNNC5SPDN1+5M
AzxU4aS2k36M2FUtz5L9Tn9sscTjls+KQ1LW9m1h6cZraIoS56GLMCWsbUe8W8O0A6kjt+iFhX+4
MrVfCM6vHbGUtuziDT9OYjjYefw4Zp7jQRwVrViEc1BC90XXc6vvGl1/okTzZ7+tGVDS+yT0P7B3
NJ8mUiiGOCOogbm4ayc52a/t6o4Ie9YPeEuz7RjZvgRXApddA17Z4xuoObCLhJw9KVgoBmJKtPhQ
rEZFJfSS53gm1m2vxabbIgcstLv2cb9HZBsdQ0GcpqEYzxuvKDGAS13VOPzQvR4uX0Sow97Ar9jD
fUWxx2duBOxLYvf5z9lLDPczEgl/QFlTvegPx5IuaWF1MLYCnnqaX6NWLbGkZHkplqkLHXoKyNal
UzO6pEc5QIPr8KEKXk7D7HJq0anuAa2rO6iZsR+pHM2hRV2rhRA4miHbw/JAOizsuZko6E8xYbWQ
daO+wsh6pPm/x8cKxq/RH6Pif2ueHjv7KxdgxqYnydz/8hqM+f1Si42+ZJrDhe8OT/Dqd+zbG6oP
1is9goOp3XquXzl/TTq8Wr21tKp1LRXnHSgv5OVEubtCCerOKfqsugZNG2/QkCVXG4B1IhcEioyh
+uWTCBKlU/7vqeDuUuXEEkmVY+qdKYuu6e2+womks0zZwi21AyVpYY1zun5JMKQPAUnv1QNMPDLz
SaEeXfMp2/gFgQ5PSbwAWsk43i1Zhl1RoYz9yiDBRY085/4/d6C7geYfPS46hU7aVSdhAUdXqtHj
GuXrt9MevZGGhzft9/FqxnKlYFDlOhrWeg3hzHVm/bDQPyVa85BEVsTaUWN+0svPBHrdAN9D/sZG
Ri643PJyxUVW1v8K9wVn0JJpdthqA1X7dgs8KhEUEq7G6Zb52ga12VImk8rVKkaaA9X+da+Y7C6I
GwUcoQmzIvC0hf8VsRPALcOUF60IQFybaIZ7v6199Y7V0zUlLp8VOQ/o5OJEBzTr3pCi4cDSFgVD
2NGJUZx5YGiFgCcLby/5BjFYPHei83OgfksW+9IBvkP6UO0PjiDeJFwXwQGEBr9vFsr65ka55P8u
hvD+VHu0DeLTvgqg+YD7KzmZWWEqsnlZ1MRxL6tAUeKgz7FQDpqTH9WFASEWnsaKsOmIeFbej8Y2
AIjhAA6Y1MOCWb9jBlsplCEe3y04r0lDQOkcjdhIna356Pv/MOjKr4slCI7X56JPTOsLPRb/eIzi
5sKF42Yqt1j9idTkUaHcnVzKflwx9nnmzsGPQvmOudpXf3DNQ+ot4Ib53bGOdhic/Nye5gW0aFUb
zSBFvqGTVtDLZxLH8iakBcjYBMX7G7pK+BB9hf50aiGNRHq4hMmtJedf/NNzCLLX1kmn2MKNid7e
EN79z68Dez+UGtF2CPgaq33KkK1FJSfn6CVM92Oq5ZTKHjVS0Tbhy1Zra6bgpeM8y2izP40rFk3h
YV37euY9ucY+iSCN6abGmN+ZAfAjKwaPLn1/Tsc1oulnmwckLIkxNAOW+mKgKkWQpAXEgUg4WjrF
1tQtOGwPcBQqY+ImprLJoZpxZ4ULomMZ/ckOi5agbYt1v8sg/P/j93J5GThsYX9bYUHtFY93yQgz
fO3TXjGI7EPXckO3QVZnyQ6ldnL1bvPdcJpwag9NB0aZoy7EPn0KXSPw1afeChlNclrRxCofXZjJ
0tEK49K4CI2Mrymg0h17mGgfP5/M5A4CT/vn8Wg6pnXNiTDuiQV4kJ+uqPGuYEurJBm8PzCr4Tgf
DHG7VySNwrSIdOLUnoiqzi0r7wTSibDBCEjUT2aBdqov4EtNAXf4M9CFA4/PhYAqu98H9CgrGjvs
ZnfDEhNdrAIm0RGomRVmkYR2tOMfdvXWwSaSJ6ST/dvVeE3dahbBVQu9rVk7gD9jWHzK0+/VWMge
AvFCT92DTdVtSwLyeqjWqcpKgR/KFMts2aXWJsx012gdDZW1GVlwuIFiU9teGtBYo521dl17DJm4
wV6j8iepF1PsIK1oAHU2T8ZNq5sh4msedjxG5qZ3ftf+RhCOPTbwXe5gUY/hGtxru03QyfJhAtix
d381+XoolbTDR+G8eOBqoNFgrcrHVglj00Qq9oFDCnHi/WgJFGJ6zagD3nCDJDY9LTXpsYxJRCSX
2+bTQ7AHOakSttOySvcMSrQsT2ujSqvB7BYEB8JakNigLhXArc6obJ7iX8oc16MG43VkvtDSIkOW
H5d76qC0iHaQBNRHw+jVjW9eJnM6ieu3hcKAR7DStJ04pE+S3C5DVv1DpyQySAczl6tYIwjOgJSW
btLHT0KhCe31ouXYtPv/xrno3utFZlW0VQMZW7PW3svDTphMBObDBPmamrEpHnCIAWwnEFNLNleU
l/6v7mB2Kn4SK4Nmo9tF9ijCQkF0e4OzHE2NhDzEiS5J9MwIWUYeR04mBhRCYvtLByLu8rWxbRhr
momUF9o8C7DD1obH1JKNgCBtu2lZclScR1D5IX8bWgg7DcWWx5XwknjVyIyWG223AEiyjPpaj0Q5
Yl8Yi/7+RdjJuuqmeSDOVQ5P6aiuIaMWITbkkkTWx+uQ9QlfJlifGw0diYbXjazKEP4mF14CePlT
lUqiKLvpMaQRlnGmr50qXzeOdTcUiEijtm8DL1YxSQ/7eAsjLimqDw85Yz7V9B/FL5uLKwI/n/4V
H/XIK9zKo/ftizejkDKKHj+tZTlqMcIOTceV1tXkoW3H2sUl1A74Yz0BSJHt1OdUQbPdwCRuQ4kt
UAWhqQEAdE/g6Hg18HS68wwTROZWyFvkTttbLNFd5doyGHz1lsFuTAy9ZdEPcY4RsIN91jKSMmIz
BshpGUuO61zCE5TyNQ0JRMo7qCohm8NSr1ZsEnkbUy0RCzhYw2usnSTv9d++jIL1h1T8Q/I6qovA
ZRvtWSqZje7VRwD+CIc9S1fFs3xavpSA+ABUjllTutmUBh3N0qyDBsNLoFjGhY5SaKwonf+6cNDT
yv3AYJAb9LRmQH4N80tUoqCCrW1Qca/JoYr2Dd/RgwnpBbhqHb0SEqkdef/RGMBVNMcH2uTWb4Vl
p4aW4gVhnaD0iUErxOqWR7t3Wk9nB66NnisZ4huQDrwrVcroIjPujxR9IpWtiRJqF+ZPuG33mGjW
XOgWXGslWvzYORoYK2W9U/lX3FglbFsOXuIZ2dFaSa+ufaXMC6MFuvSsbUOHSVyPpu+sqP0ld3WX
XsyJV4/Hq/yDCSYQj9dUTh6X5AW2RcQKpe19K+DyEwrtIIuHnyXBQtkSQYIxSG9qgiw+lgYrCvm/
8KG2ZLTIm4vRPtswn/KtQndhvfo1utE1L/jf1MAA2m5oRWR9YjAR0PgP0rZakty4IPH/42zxBMot
kZsBoV6m0oBUoFvid7AlpCyxcbXke6JGB3PaTxonlgvC6SujClmpwBHlxJrMhINsJXQTJu+CwtMT
GGxmO11ukca1s2g0NLuByDaP1YXYj0qVG+k/r+Lvil6jOPhxtVJQVOjYuY5SUYDDNeDHEPnhoNvI
be5fHEEQhXlL9hBBUcd40JITgLWk3nfg4Ja0ctv4EDA/QnQGBiyJsAqXYcTAZEg8eSKrJjUHWICJ
PRvZBhzDg8FJLlfH7aCRh88NCZtj6HDoZn2Orpr95YW01VIXTPZkP+XZli4R0v2N61lJMDQwL8VR
SsU2ih8+4E4g4+sUflc14XOlhfV7WseelfbM0gIaM5ItaPCc+vccmdl0nb++WYR28l/nppc0srbH
ovRfxqIqi8vcAgliNICiP5S7d+algZSE58U29gtfpaUOwYS9KmrskhOrLTJ+SicBfWOR/xaf8c6w
dnhmNwmWxzl6XV3KG5VhM0IFqTlRvSQBVmWLlWYq5Swu6gDx1yKqBqNyTFEsOz8ew1bsvcoYiZ1Z
WzQgQc4+RBkkG+jfzRyEbB8DHg+Hyxu34XMo0QvksDrCaod7rBIw4sU8vnqtM2HHxy0Q69S+KQqv
yrmyDIiy5Q6iaVQYeSE46fwnQJ/pfSUyNW2U4Tua5tBLPHwIA+JMoFDqMZqhQT8MKEgAh3Y8gOoE
0Iu0Eu4Y8JFlyOimzDox6WoBUgLLIbNk6jfBllwdtQu4Np7ltf458yG59FV7fpLzVREt/CdVrM/s
/1FxFwRsb322bS7COK4GgnqiWdd8pjuDwi2OU7M37P3JRVzGiZokvO66AADDY6hfnxNeKh5ziJc3
8yvashg9/tP6PeabxLgKCIrtrWhp9BBX7hZ34586RUFfKBX5jClc1PXH7JMFqh/H2pCMoXjIRNNc
r4iaDM/9j3GxJsxAyd2inaZmGP0UOilzduOK/AnaZGGQYCRvY7m51Vjm3rRxoBkr6QRm4YwpOpKt
BXbVZwPtxYUM6Rz1nGTqLSqkAUgTYjsPc8fyIS4Lnfiao6PXrgf76crzrLAJerFBQPXwPOm2NDbJ
gQuXgyRYNC/a+KENhr4FY281WlflvVm3bqKnC/Prp6XZc7ZRG/HWYZb0ksgVOspXQPW2nLZE4Mf5
uGgZvPEPC/Px+3OJta104FiHOFSnKglJf4xYhvR6ivTZNsoCKh5tF2ez+zxbJEfAZ30HNp0lWcpg
1O+BVeSgFWpODPMOgq6PPeBmufumg5EGzXq6bm5VvH7KIiZXFRd5Dz5xHA9QzwkoFF4gbRC8c73i
uRgJFo8VC9S5sYDmC8I2TRidLL61JkGmDZJTwBgNHQLJGsIsxmY1er7yZvBIWBeYfyItLnMvCclv
ZTAf1YiXc2n+hgjqc1OX1P83Bf+zG8/epfVXXTmNR/l92bgALOUgRN/3GoMNOjQhw9XKN6YqRiYN
XTo2ZRTPV4psIIeCRryPbIEZbx5aYjbOJdcnq2FHxQZ1QFhrF9jvQG+yQkND4t7CI27uMXHALH3t
cj/UQlyt1CIAJlm93Ev9UYbJtbP104w7l8YcCAZAsbxwMh9vJ9a3MYlnU/eBskB+LlEQsQ3Bi8ez
ECXeLe+ZqntcmRPPlMPHNgY5ESwjRMjJ1aOW30Cm1Os0Z3iS9dHsiP8b+jQ+D9qTw/Q2OUfjtXei
LhnQycfIAa0b4to9DNmWwrXlBDlJL/PDq8tK/OVoOrwbGcVkiFu1uqK9NAWt/WSRmeE0MYO2ubqM
ULFO+DQq1ViPSD4atYAnmQhSdaQOTE2Wf2en4o5barPpNK0wCtLaNXNouYv5Il9nj1heGVxuJ4Re
ECeNwT6QbmmKWYXQqo/DmUkHx5nkUfjGLhT1EupCTZOoA2J/LRJveuG2iPfLDz8hT0K7DhIpWGn6
6vYUaBvJzX8olJTqI16vSR9/V2Ra2JThuTyjlUiiX4SJFIkhoJYp4ABXqdfH75xTDDUB+jL/dYlS
0/3QbH5A+O9/YY34a1DdICyQBJrdCqULxURxJn4bbaaDa+ClRpsgGFHiwQj5+wehdwz3UGfhTddM
oa48RBsYNF2RRcFPoxkEnb2r3/trrompmJagMObLv30BcM7ey9F3YUvsyy8CtIv4I76vvtpMFvx9
1S+1Hso90tc6Xz+csZsME/MsAovnmmhGSkhjo3wkcm/o0Zp9X4n6/CnMQW0l4CC0WxA7eAaWTqml
ERwMBQ2AZ+q8goD5AVVuIuP7PFVhvgNBoNzOK7m1yG/9wdgERMIFhm2ovr/fy6gU1Oe8/Q1xkdEn
Ez7ld8PxfAhlb0cAUt4oAKJJXhJWXBvUmIm6laLHbfhSG2PSvWNWplv37i2PQmaSzI8Fwfdn75LP
8Yun4MQaUdf8dqxTQ70nz4MyA6YtL8fgMCNYsNdrDCUCjj7BgdxL8NiMJ3ZU1QJKMikn5j6VsKCg
cutkhVJD80y29FGqPCvgE+Bq32h6B58uEDq7Eg93upFMva9aXE92xAvcBzpSH136H3kc71gwWQNr
Er0MUCJ1RM8s6xSYKkBoiONRAJZIs9PmrTgJZixcDlCZrZm2LeZK3U1EmX8UUKL3hBlVGR08V/Mv
kGJw1X8FEMD3dpI2W7rZ3ofuEwjopfLVCII0QCAe+IrCVHg0kH+kdufv6XyNMoKWFFiJWyqMFOGn
owJDeHwMSmLUQRAWCyPS8IJ2+oHD7QRZEy2Pji0HG0TbpzVAY9g10ykjge0iQ77eQIj7SwEPyytc
BvJdJ0hVbcc01J971I9MjP1NRE7x+BJ1w6QBR2UGeCWZtFwRs3SV5F9QiES/yJfm3DezBiYopDAt
4yKX8WHOzINcPTzk812NzBLBPr0rpeBANXX4lXs7Rr66xTSTp7UeQUD/PPKtI6myEGLM+NPmluvr
tN091nzWKD2QPv+prdAEjVXWDxQCZIpZ1y6IMOgRhMsNau6nbOVJ1aFrKzFjpbE3z1LVjmelJVTn
SxqNpkCWjAZUFUiU08TjRlsMF9r5x41MFlCskhV7YQlCEyTqFBaTfm2KvNDtQtld4iRZyrPdJfAD
KVkQ75EiIEyImhGf1J8px504e8F4aPXp1tekHVDlcYRJpU93W8tpdoGRcG1PEd+xtEwcpKQnRel1
3IsRVPz729BpkP1CZmk0BcX+VkDjQOrP+JiR77AQu4PijqaeNCQDAXU4zuffqvaQBAj9eGHSnY2e
+Dx+tOYZ+CknFns8D8+DVXeKvumRQz7T6qiR+NaYvrMgbXDS+JjKYp32UmcrcMwrXciuyNnSkgnp
RTigiGh4hKhEkMuKmwoVflzLoeDGpGm9XZvwZ6k1aLNpmegNKwZe7a3pnrdJghqaqo5VxWp04Mxy
Z3aXbfcrYId9DfnSWzYzpzRst+eikIRsYEKCkcAu3sBorHNJJrKkIYtoRa2s1XWT2+S/iXpilqO2
mdzwEtBgygducTgn6LD5rk7KlUchL++nImfTzlCxyyP6zJZDMYSSgyNnM5MKhMQQ/tVngbbQVGd+
VONevBsRpK+sN+FH//Z8bZmlTUwgY4d9ZhboJHQioFgY9sQq1AsgGFUtyzDdYcfhu9tUgmiZRpTH
AZHDuuEaGXzVQmqo7Wu0GwlkyuAi3shhQHmw9FQL7wiNFmT0S7n22uw3A6os9TfpZgOzO4nnxiLl
GeBP4MF3V7+wuezHsjOYP3orDc313O2BKJzVtQvZNRbOaRkvaetTSFt3VQfmJpk0GK4ECxEiQgtD
mwSrpdU+k1SGaGZPopVl0E8ypVabiEKGQkJwUWcUVXYBCjQW3E9ErHCYTlQVUat931MMXj5qenyW
hvMdALwglHWk4AOTpO4VbP5tumS5k6HFTHLxzN8hJ6uzDKc1qYPNrt4tv2JlBlmJOXouW1rXT7yA
jAA9YIVXDo5dnf3lMZencD8bcDXk6Ikw/0SMBTQ/f4KkUzjqXUWlHZJRJdBG9FWuU+i+Oqq/0Nhi
vyLo0T1PJs37QEhY3EKU6L88E/4JXrurZyGdFMBVPwdBWV+d8FXo/34cRc0zwjiExm4BEm2nfpR3
troV8lWOmwtI+nLSsw5psYOvwCTQYt3GfT5M19V9yDGnvGT5W2ISspP1reiOZDDd7eTNSzyeKpmu
V4DcpQfuAONV4Cs6YWs0cH2/Vh/xE37OxZVyPr0TYTayE6t3uoT6ScwjkXIr2hQjiAW6AjMsYYvy
qs5jS/NaSQyJN6HrwE+/wWuRaQQhre/WCqg1yd4mcLKBeouVoCWp0QeOKHEn2wcCB0hTvyP/45Y/
0/VZsynuF6TzKQSFvhB8iEuEZUR8MLmIJkYENZQmIA7y0soqLNvZ9epGJqk5GObiDzhMWDfYYz1w
ypu9B7ooCK5Ny16i1sWUzhk54CCQWty68sapyvuLU0jtPCOKiKwmfHnpPV3xd4xuZmzsnRGnWFJ0
zViL0nVYxD6+S/hjiIEThd9EHt+PjimUsytub7f5qIZTjSagXBVMFdVz2VR/WP7X2uRWWu2j+rOv
/fywS04ppQB08hxXzxBnIUcugxhp5eihGESO4kfM726NsHsI/BEVOMdShLnvNZ5Q5g6d9skDmKB6
TQChvtMxCbi456swAem+kx/RrPOJ1f+G2IX86gM2+0hDXf+kmu/3LxFUe8zRUqmdp58kTs2BkJf7
9Y8YMjZ9gAFMhZ4VOZdrstsToYtPX6ocJ6C1scgalD4HDk/3AhNcglPpnUzITFXxrmJdlH+wB3Wk
pgnyDn5M9fBed5NhpWlPbW4cDaQ0qn0dfx5La4QTHGCWlVZi0FiziXdgtHsWRzIOwlbWEZblwpUZ
MGU11ih6QJIZ3SBfCL+JApWOII9vOWsoDqjB+erYEpGoddg80m9fZVxdts5qzNKpqt5I+Iv7LXkb
9AvfXDlZ9F67OGpk0O/39yABT71KTox2fPCPbEvysYYbG2daDqNW2iLohshO/YRJNxoILWYNmMPT
EYjLld+M1qcaUdrE4LtY5wBgEsXYmAkpuaCcXF6TzvErOR7K88Np7Fbc9b4hsk/lb/oScQFUWlg4
EU8EF2DFUA9NZS71m0fL96d/f5PKa1muo25XmsjOz9IfZdbNYyM8vafsG4s81ClAuuEHrybHxk6X
w+cYARmOpaSnf3VaJPJWv2dgWaRVCNhBEGs1ZX8NkzE5y4p0qEmSYR1u9X/CmmpYKbuuLpOCwWrS
kPwaBgtXCZYJoW/F+Tt6LHt7vFf2lfcKNrZSHI4pCVUPiV9tmfqfQdLe7hTCPeHPoLubD/sMNRRC
CYfxfgBklbBwbH3z7mMaNl7K5nI4NIs9AgrU9JCgeX0wNE8DGy6dKV0W9Be98NcGaZLvcjLupLpJ
1jBuyTix3DGNiWrVJi6esOkWrTuQFYS/E33Df9VWKh4JQTgA24iYe0vw1TXmBNuCWv7C5TWSvqUF
Q1nTFhzz+CtVmgE+hSDKRtlVMT4eRktvy6QmxwdNE/E36yREEmTGJswO/+naKE/2061nN3O+KTR+
YBZYCcMshK6iXzowv2YL2XvWtQC6eL/WaWLG6ms4LhnOTOGjY/jOCb7MOcGh8ryycr7ou42gXJGP
dF9nOglM6OCv9dD4Bk7batSecT+1OkHDXOqazzvZoUFM04YUaGTAUn76T0yfg5bhckx5PXxjgWkT
mtYTDZ48bjLLxWooAxYBBmy0ftXpwfTMMItnPegMLLX7fUM1g0NKdy13SWjIVEcSli4QhD1CWqIn
gmrCtsUb4hGe89yaC5EEjn2561MhM3QGsAz45i8mETepuuleANZs3E7iwIHHB2YGJf70ZGEoPiAJ
X9WoTuiAdmPlqiehWTtMMwYmGrxDLExfTlBS+U8jiLUDj8qzk0INm329BS90pMqv79A790KCxH/Z
Mn+ZQqICdC8AcR/KA44E/05XHnciwODRj6AQ6wPVdXdKX5IIo1/5YDlsDVze12OFLw3OKNwoM3cP
fUtr4eyeR2XR5LTFgriu/UZQCbi7SHnDwDysPwkOGqzXJhjbpQe6uh8IF8HKgWtDGFM5rP+tyxIO
bxNxncDyGfI8X3yZd/xNHPgTs1gws8LEcJNUfWYTpFe9DkYVC3GOjbxbFRfFlB97r79iRwAbFWhj
4jYU1qNbF/JAMw3cxDf52fzqyc9BZN/3x/L1jyI1fHYKlzCdYxd/svarRzW6EmqrgABY7DozZ7nZ
aKyQrnH4UJGgBwFXMsLeNkSyCd5Rw3eBXv4crHHmny/a33lWP+9D2q2WyjK9z/DnU9uWwu5CFuES
NLMyyKqujEiKyiSEhYjfS3XxRCl8j5vp+IT8SPK2NsLXSh/7DiE5a0HjWwjIKBwA2DKRmR02C3s0
Mi5nK+PzyCQzFvolpJZNR1J0o8kE46OxJ7sGDnqALFTsammWpVdoKOSN5GH11IK2k4YiUeuTQT15
PoCKzfz0fAL1CeSa58XTFmgWLzbL2Mv8qoz6s+H5gpzBDTwVj09WVCrs3N65IWj5T7bbGpO7gbCT
pynRf6q2NlDf/tj2Cf6TarsteFDL70W6GziMiobuaoFp8efLVJqUOmvkOkIBs9cCzXtCCLS3MLQf
inF3kxJ5bmMgJYYOODby3lPl93Bh0yG2MhUhgkP3fgzmgUCAaz8V4E3Ywc6qNhVQEsSECILRDxB5
MPkVOiqmIUv/vuGpPM+NQ7clgqVSjNGjnB3T8dRK6kF9wb8VGTT22TNxJvj+vF58PQFd2hOPB97Z
c2o29D2vJEqfVxJFQkdrPAC73hBU09SF9dQ+2BdQeDs8J65Bj9gofbRQAYRNHsXtfDIPRdx0kXzT
dcz5z3+MjEyk6i3Kqmg3PJZivzYbd500/2t2I52Hh/kq4ts0QFTzelV8EnEnjPG+f+3A9H63hPNL
7VYQyaf3kpJ61wquV1oH6JpjBMaTp7O2br01jn2zZHb6iNP4DuWCsld/FAibLfFToLej6tlwAgnU
Upl+CTtxIx7TkuawRiUXKTaF8v+dwIU0klFycsHA7GS6yaAwjAW3I11du9va1nxFeaUHvyZZwRn8
n9l7Ms3d+AXXtTvS7rcJPgzrfzuIwxsoqiT/cgm3RCoU6FSf7qHgVkbVCSh4K5z1Zd3bLsyP9YWD
KKbCErUS9AhVEaFMVH7SNU7iovye9izhQbJnBJtXZRKWiL043/TRWRTN6FXAHpvuyumbX7YiFGWY
zB7eZ5BFwe5z2dSlm1BCSrE7pWWWiYw+YeTLA8vsv98Z/ELrad440kMzNwHGGigsiF8IAash/N/E
ZFA8LMM3iLxgzDR6ZEqEkCi/Fw+XEqIqRA7AmReTkEfqshHN7KTLhWEAzDy7d6C5D/U00CwmFrgi
atJtomdTHAboHXOM0a0SnnQZonfLPvd6OhNmBrw0Q0I2nQ6KitemebFBBMbaKrbeGobXgl+TIFVR
X8KWDqqxdx16QS29x56bI6czy+opXbWGYGklK9cFHRzoQg9ATYsMq5FAohbStHIYI3ShqzYAxaF/
cHeK+cyGwJyGh1UF/57H6v5IDfLLdMmCCpVN1D94fVj7AWEA2tPyiwuENsKsKaDUBqu/jcOY8ltN
bosJNoDmePcgAdhxrS4C/3m7JK++gNHPlfZjh0zr1hKqezfNq/N3BkRRw2OL6CE+uEBkN2UAz0lU
Fq+EH84ndPyxZlgG8giRVqls82QP9EMDLWoU3fc0T4u3DBQlSMKh/fe0s1nSFTBo77eY04RwemIt
//T65DsNONCRd5nUNAtGlNuhJaH7mF52RijewS/orlCbbkFCHnNInYeiVh/YMVfk2v96yNjcixps
zZ7hvuQd6uwufMpNcPyWMiir/6/dEDibF1oPrqvzuMSi3Yr5hC1521Lv1Sn9ZjZyMflGRVderXFv
oSsuHhmJ8/HagjtoIF16z3+h4e1nQWs0XDAyldofhh4Bog+I4AxlmsL4ZnBOXpNRNFh4Nr2nDAw5
jF8mUVnAMZRFE/CUlsmQnwamU358u5iD7fuNoLVJfwHg90r7a9ZZNr+BhbKTB9YgNw7p5hJ93u0g
ycgAfftQ7x8MzsfyJrm0C6n+A03M22oBSvTTSDnt2sryH8c5u9SBAlWUDjZD57eFxLKoG0J0ouXT
SvLxpKuCZt0aBoUYAtvnLdtxiQ2FzwoamGDsoWGSx6/9y6/QTfDQOCb9GiZeDMM3y1nyfxdNWbVL
OKLwO9w+vWI7clRTvfT7YiolDflotxPSvUbJE+egRwKiRTu7Efn3lVuZHWgDdBcr6mfm3d2bnDtE
qg/Ibv9DpDOxR9ddpYU5UAu6IyLnBGiieZ94QiG8IT5pHk2obW587o1eUyYa125Lr+DYVV2BLO+L
8sAyeJYqfvBpRCRmp5zk1CwpXVnUgZLgsBWPgNnKg50AprXecSaNpe/KbVOhoFheAGxFbCKrAsQW
2L1AumQ4g83fiC7cojYUlh4OTH8aSF13RiH3wudhhnfy3DSGuMcRTOB7k5WMMsG7tpknnLChWp+/
OckQHw7RXNnBkOuWi75oJdh6HubR7XUN9kb2kh+kBdBs6n24eYKudrk0Cjyj6fzCRvOMwNzNm1tJ
X8s7x9p6WQu0j8R4/UTT42RZPEnnUERMW2OdS8qpgog5mKlxyTyodd534jO4xYusOqc58apCBii0
ROSRcJyO0NV4/4v1OVT9ydb7dtwnJvOuIttIvgKX1oT3GykVVVVcKTW7n5asDr9UmRa1PTT3XMz5
lVDuADur6yfQI7LD4qCmIul3ShVfcyWTCnM2TmsfFELNJhficvbNp1TXizBmxH4CSOPymQgDmMmv
G6Hs1C1oi8obgeEaT7yg/vFxinrOqJJwk0VKKxq/1117XQ3IWQF5Id6LXXM9zsmWRLjcH2X0TGEm
13CCtQ0k4kEFKM1fkkv+im71MfMIAVVCuNPXw7K6WtCNWcngNKe4UPFNTBi3ScnYAFo/JuTRPDd3
EveS1Q38kP00+LNpLOxtJAAyiFuew+fTy/UbnbXW/Bjke0tgp8RHwSr7kU/ECmO3D/JMfMXwuarR
22JPJeeVWB4WkXXM0iBOz9UnDF9M3KuQNkcNiyjw7lY2sXVUFD4MMlvs1o2scRGzaYhzrsApVpJ1
hPLL21/dm5eF1CnWEamCOayiWuz8ipmU0IwhwXEocez8FpEtyOabjhq2XerzkdUZ2u2sjDVx5+nV
WE7Q3Xth2YKQ2nf9QxyycDVxOewkd+jUY0YE8M2mCrWr0iNgXWivLDm/1iElkzHsr6RjzdIbYGLA
WjdbRb05UbRQl+EWIqv/El7eITR51diOLaCccPhlfArOVArSP4rpuBDriif26x2BZofcoTEedypH
rE4VqVOoySUJ6szIjA2UD6Lyd/ORV3kcrb5DegN5t/Yao8IalKj6hgWWkc0ekP1EnsSjyJgAyswB
qSN4cycStSdw2dh7V+DaptZaLo8HSb6+9zgiNAJ77SRstBMEY369B5FNRA0FTA6PJS5L1WDD/mVl
NHfLZ8fNwornzCw5Trz1RE9yP9sRReGKY8MiEljG+tAqxe0OH7pZOZkholTnj13kkLPfIUnNxjDH
JPLTHsHx+D+9VJtN7bwKfXTCWr/uZoI7iXsxCvPNHfhsdodmsGa/5LwJDj8l3eUNGBiYhHz2D3K2
R2Kr7XJkZPuHL+LPv+yqBt4jKscNpH/3cGgi+Dglm/QRdbjK0up4dFK6VOppHy3YEmxgWxY8hQk2
a+vjjg1nw7LZ0Rrpeb0PTZOVP3W4MxvPsx2+2xFVerqBbCPITcJbtrFN7ajfwRWf7Be6bjUP4IHF
GdBVB/ApnQUUrXAyA96/NICSdLszzc1SXVL0/UJ5KAyIETDqZ2CKBTz85WvFmylOzwaMPwAKHsVN
XnLUtpd5o8ZHjjnHPJCr/tFMGDmO+QJHgbq7bscwwv1lQDJCAWk4xXA0xpQXbhNgbJl6XVT0uYXC
2MOAckqLzd5GRtGfbq6oJeK5Uwxh4gsSWOaptR0usJ1kqyol1Dmsl4rLUirW9dajm8OBl5Z5Hkaq
+7JueA8KLdc0+5dw8CNcl8CBk22xZDP/c+hM3gE5PgTmB5QK+Dhz+k8zRK8lpw2moscEUHmSobQQ
Vt7VAOOwxxA3ZuiL44eJXxMwvRwEHZGXDg3709i/yhr5VCZFyOdMMjhGxZ7YuqjfivPjK4JdnzrR
BPnGUaaj0cCOD/XUqGmDUwYeb/NuIt9BtIR0AE/O+JuxnlJkPk51CIt8TEcab6Qt+TIsUBBrivRQ
kZxtuxA9h10iB+ngnbo15qX4yh9yN3u8AWYbICUzyo6pZCKudDW3ELEltM/Jugap7Tbh1Mes6ZqI
KoC3tqMnBwLFbFgWOkmyoF8f+TgTyTnC9lG4TXEkRd2GU4YK04T6JWXzjvHAtkb4LBs7XEL7BgNJ
wnp1LNPrZnL/xu7nQm45/jkroNJxWoSXGby2Z3y1MnQNKjMksJP8zPNH2WoS/4zzb1VSQm5wiRC1
LfKNqeHEiic3VkwBS01yHrXpi+hvRhmQhDY7Ft+Cspsg3C8j2DmcpaOSwSqoq/m9q++hVbueqUTU
b9ZGx2+B1i/OA76SUSHJpTpc2mktWc4rzbLfenhIDvlxM5Aea26pd6RuSturrH1N5QynIvyH/CKQ
dI6lsT3R3QoPT5xDgy1w+gtuhw155BNOzqtLG3A0s0ifrdcPMfVUW3ZE1kvIhOsiTB1iDEH+YZeS
eg2fvAPTL7iZ8wmy68XuaoHCth4BJrsrpJuGo+DyRJKBdhY7Q8Q69XeGpqBhTEcWE6vGH5eZ5+o6
7GO0RkoX2wjya4IY58cip37p1vATAMCRlrk6pvoICMC0oZX9PV3+YjRsYJeQIVlEmfaUfxvmVxW8
LweXfAZjuBK45A/pEGbO8baNU3esmXqZQnlW8dCIdA2o7RurA61BWpJpROTB8nNY/DLcwI3+RD4P
W9Hf1RC3u1Y1PyG7XKVQp3m/Rqe8zW52olUi/0xQvU9hYbC9sqV7qKP5PzMMcnCk5FTiafkX8jNQ
7dXFEOlD/xjGqw83aLqEq7aoZ/kobI3OEr8Iwj3acQw+zbOYDYGhlGF8WE6ZThW/jUcGw5nOynys
quURSYnuX+q84qCUQIc6eqOgt5S7DOzUSE7xf1+vNRSej1RFpU+vRj8tNQrfGUM4o5aKsBhv8h8Q
PN0OPocDXehubPW1ntxWF22yHO4E9M/n4BXGgQeihVnckJBmKkVFfrvfhUFs46gplNRcYaCbhZJV
fobR3iyqEH0Kw/VU+kmlFgNoV+Wwojm4DAnXtZDW2cfdfWxdckH9uWTEsymt1mt+OhmVxn4jfg/z
DmhzAQwOXhhSH3eMPKSoJKPdbNNqNQEPx3b2ikJMSCLy++nJE1EBF+JCHmfI6dD6xBr6Aa/LcKCY
cUi20y2zzD6KNipSsG93OHmeIWXzMyQVGV3VK1IzUu5ThJDBfIZTwzHgp/jDZXmXG//Y1OjDMKBX
+P4QVLZ6Fwyp0zcEZyOHDQ39oqfJ3Mj3wkoZY2G0N+EaN1g9ogFDjodAuyA2BdhVX7d4phTFl9wq
XNMucA3VOvOjWdrY9cHiRbitCV3kk9TBOrz5THkTf4/lOArEjHGNMyUVM6Wf+VHQtC8B0qAgcsIx
RQEVpG07EahyWWUaTQW7aiStmFVUqxij1PTrdu5kVOCEnIW4wD0N1XyTy7S3rev6cx2Rs1j9f997
ihjp9u3Q9DO/DEb4B/KbLDkXbs2U5/xDAokt576BQ6hoWbjtlP5a+AXp3F6w4PHM9vGH1WNP8wgN
wvlYOQjL5H33/YGG5gt+66jTKTW/h+iO3UPGYaTpFbaDwG+s+EMMUVNkEgsA14/e3r/85Wy3nQCV
Wg8baVzPcVVhsIGwSZqh1llxRxCs7SFHDtmat6tBT2njoRAM4GMxpZmu3yGicrjjLvQW2sslz71Z
MB+SMHrvl1hz53MJda+BBbrfPng0gpKepz6EiCDo4GpWyDtRe47RUD3EI+1FL+YqXZvPGoG6rard
3ZzpUNZAo59euOlQKfYmJqI+eDHt+U1bbHqdAjEIGAdsrWBRjc9VRKobwy7Gru8B2YHIetf7SISO
6ElCw0WNjg/DXZr0j/HImCP+ED9TVeNEvx/lHqpaJ0hvX+2HqEH+5DC7srVB1bmUI4OzlO9ZQn/o
2eQgTTUPh0aA4hwTWCfFYPQMo6lF7JTtv6Rj2b+RhyLQdARKwqWIrvxAH07+DnC0/OuYGslwZ3jh
nGx7At0YDgfE+nTCnniH+jcpOb6Ubs1ulwkLLYnqygLnji3pPqA2JVP9oFX+YnPG/S/VMiDONfwY
GZfWNaOeRf5X7mWkp2Xmc2IyiqYm5fd3aLvdKyMjb2zyPVZth9RV8mUrtliPw4h7Hg5+rWW1I7vA
KxP6nZtjnXY8iguwbAWdvVkxa2InNU9oliFhVj7H0mbqAmNX8SWkpDrN+JVgtnww1E4CXK6gc0FP
byCAd141TmyROlA5EPWR8oMMD+tbpOPn5QOvMgaopYMclE1PvSmQX7nwGgzcsHg6JwfgHItGvVjG
TLA0wct967FqKygtZU5z+1ajEmrOHgaoFpHqa/g4CZTTotjPbsgLifFDMf0Tv864Cs1bAS5C9FVF
4Kfm0SbdEHSee1Tkkea/hg67JB/hO9zw24whZssU/7pjUqD2xGOJcvePkx/BZwSrNACJmTzvAKd7
vvkDygQgoOROOXjzAEr/rkuCSxDtAFriuNGKhNihaAzdXGmRx9+LSxrlCzFQecB6mh9EplKBluAG
suSsBoAO8rfFUe1wJqgbona9d1pHM3BhU4uKr4jtoFxLU/88MOGAO5MyhU+XoyL9VcYxtZE4QP/8
6RYzam6DyKHG74FbBehhXJfNcwknKcVwQcyba1GKWvDRlI39R/WujWiwU1hC6dGfpz8sQWb+Tk13
mBFJH5shqhAfT+hYhMXwiG3soJlamzmPZY2+6MLrsH0tnbTnIT/jdKXs+5P97hKu0feFjhL55a75
mso8w0cg9SSH78wkPRGBGtLLxG7luFnb3+CKuejQdX0nU2Me3Egu9K5eWSgqoi0TG8N74jsxvx2C
2QuL+2sHCTVEDPzLaSa8iAhbjTCGUMWH7C3IKojBg5smKtPjeIbL9LUsEKepMyl+Tlx7tS3rqAja
Dzo2wLS0/3IVeqf8upeOo6zROdfawR9UhVSdzvTPo3mKrKTCboy7BDnagVexjlXB8btnck+rPXJV
yKsdDtt//9rXbp1yGV27OEbYddxLtetrX+YhWLHzD3FYwe/9yxxoR/AcnCwRLAOFNqGFLtBRC/5U
xtrN3G8MCAl7HpGHsR2wilfeHCGVc9HKhA1SuYGhXT8Zjidq1KQUa1IuLqPZrLiFSwGhe2n1GA3h
GuSpL6kL+NHuMvVaUj30cOSVlLLjCmWPCWUW0f5tpgZEeCp/W3hnpWTeHcyFFZQKUzxswMFxGFNO
ahgP9JkLaVhp7+hMHG9haCGnDMCW4+IY45W/6jRf5ptqQV2abo2hiPusOL/FmRzPWyqVoMdeesQT
dvq3e8IOSx625RxOhso0TTJkoGtP5cagDraX7DvGic3k+ktuic6UqqLYxOlPN8C5ehc0NK/f7ujx
cBcKU60HufG2+lXzY2hO9N7BhVC5HNCJ6ZvtmQ7QpDzgqshYq2yO1z2QudmXZ6XacWrYMtLAQJJV
6u6n5sZlnSMCu45kgLIeP5/ouQWrlZTo3RCdfMVRvQG4nzJzDE3wMURMRvbDiWp4gH17OU7dfZCP
U2Im82TQ8tT1kufydTfiClR0+XJ6wOcFHG3QHggf+aoXZ38cH1v4waui2T5/MaHZQkoKrc/ugczZ
fwcvm3V0A1l5DiANmh9uAUzjvTnF/HkwluYB5MMC94SPPP7JK0PcdlnNko3J8O5oETElW2nAli6p
6i6+Qe71E+gRKiG0qxhOBonsqe1U6atHvNpO0D8hPhTN07YtGf4RXoW0vU5hthiJj3xVY1zgYD1N
DoybWX3kw45tWMbwXDn3qUsndCrlWWQLeV36GjJgkUY+Rvnx5NAaWaYBeryI4ORVe/h4iHgFwK13
8fYr6+blnm8u/DmBiy4ASw4O8MrUcO9vdDYeAB7td+batvIEG5wsGXJGJvv4socmxGnf+tzkhpjY
7b0UTKw2esVB3/cHmxv/FV8bSQjxrMVapYfZdpql/ndkzzOGGCSG0sESP2xAZRWcDf9vOMYQ2cHK
BOPAShEtxyVmRig1UsYGyiKZOSb+7hFiOPgzMpCU/fY5vIBhOgqBY9y2wj+1ElIh2jCcUooYqGee
gx+/FKlcxdJO1adyOjtzV1hqrsWFSLYGk2lyDyL3WaGRPi1K4mSqa9eIQgxSIcNzL9/xUJ/foQd7
seV9Z9N+QZv027QSFM6Up4QlC98BX8lhucibgzIsbmFfALhzfv5ghjF1a3pA9SjIH470PsGZ8RyD
CwLw4XBXQTp3H+J4F8ErPgkeNOgmLKA1Mwdpm2UA5tgnNUPnh3+FlPcz1ZFDpuTZwgcndT2zTz5U
+NvVqoUoajFyupNZoKHQbHXaRGnFu5NUdzZa6j7y7CIjWoQcX/KdkUaTnBxatbyfXvfOXnu/uF+6
aNS29E3dTiyqjue1mg5061JDfH2xNyN9rprGTd+9d5fA/ZKISahXAN3t1mdjKoge3lbU7Vqe4BE0
tqvI8PxPjFgARKX0hI3NT6HEqg/0/0BDRd9VS35qEemZMsUE0eybqYGEbvhNgh2nloFFSlV3cioz
lYsA9EXZIqRvgQKPihSVY4SNb4sQPsBM0kSacjqxEIJPK5x0NwSVxIXQGVHB6f2i2lUzumJXQQKX
aJmJvmvRl9l1U6jM73RK079w9bgpAkWocBzToeZ5IR7JX40lHkg8S5/Dmg3y+FKsTUGzEbKBNKUw
hTdNJUjbW1vcsz4wpGKGbbTL1S3zNXlsy0rCNFonnqEELnhP1Q/+0SbufvaOqDdqqsi5GqQL1BgO
zHSf5JjD8Sx/+SpvpyLU0Rh1Qpq49Lni4gJ3YT0klStmdRdzbAZZKGvOiaNF8a5oRcJ6VQS8kIpC
KhkTPM+r36AgU2IxQ8fvTCnzpu8D4VXhz1Nz+Kg3xFmSEZQCdINlFIx419/zZQwcwW9W6P3ECHkc
gUyJH7bdIEXbDfNtqhrlc4HoseigJVfcObTCMqwHzSLm5fbc1Xo4Ptna7XZjR69xw1+94hS7V+Bd
i+4MSqlpZVO8qgS5QwkX5TkhclOhiegiX/8FhoDPboU7m2xazQHS9FzYPZ+BZESg9gfVKQl1KU2y
lmoR5Bu0Aw1n+WmljRxHXDb5oCjC6MNmtwUtQ/aj9mTNH756TxWIz/VNWjD/G3Qf7lIvjs07npQi
SPEakNYIkcQHnUYd8oBAwBJ+DvW9ukTcrEcp4o+9CZ7iSYq9r3RypWmxbCMihh3k0sBq/KWRDWN3
dJ19CPgpzCW1m7k233/ll9WAtbeoTrHGiLt5SMz4cQCD/7OjhKLtSuwcm18MVGMl+xoNhpwRr8QZ
YOMS+0GkpCPVxNz1VN+ofocnjlj+sWUkXWGUVpIYSD088+5HPqZHv+CagXCJ7GszRxv44SEFS4qO
xWdDhmA5tM0/Vd6ilYr8nQH22d8b2cBun15jrY4+eQi4lfs40+GSdGmrRRmhcl20ySk5kWbUMvjm
Og43V0pnh0BkVumjrcVda5FxQ10FsAdhT1LQlWAEQs3+M5GVKq9/RyF2d+GZ0QWHPliKqdzj4XZO
sv3yGWqA0Fe0Lvkjxszm/177Ze3/tAgAVhO/SsTNsVfqCCW2sfXCSFVb2rX90R651VTdYPajWCqr
uD+0S6i6yLGXzIvsjiW5+v9Ae0y8EC8rWCfWOVS8v3NcIh/E7ZJOWMMJ8/Bzz6GIw8OhX8ktu55u
fv2qogmTFXNus7HG2Y+eoZ8h1hEvS2URRlPzJurTwpuU5Jkvq1juqozRt+Cmx2hfejX59iRuzN0F
/sdPP1/PyAvcFANmMX3apb/zr8ThBJN7BljXeEzQ/ejVfqmF0bB1I9GGh6t3m87acgah1GyF1lgi
o71G0ECnyEB8U1k6odLAxQqpCdJL0fw+t1N+V68R11xf2S86QSerbbKwtX3H/NY5/EP6tGn+Ghvg
FZ6Cb53rEVBktk4j0O0cFIcjP2zJH8d4KPFDWCjtXOk5MGZRJSUnS43mpVC0dZaYf58LwSOLuXVy
UDvxqs2natYNFY+BH+spWgLnw4y34kGM42NIZ+AGf7S3oOHk7I0YyK4aAqMLoUqPDrm4Yu0bgOGj
EkyN+LOKFXgjFoLFZjAaa4Z0r7TPZqDApODcZSw2d7f0EKHq4KXHSyFd10hu0vBYKIp2vF4pncBw
luENkDef/5t2W3Qk6aEIVRb3psu26wWOpdHCXCPKD0NJxIpzSWqTUd4lD6cBd3pKxLeUyYYVablk
F0nbF/o24C/vVfXzvye+YS8dfiCA3397b0A3Klt9zoLvYzAhIyc9U19TxPkCcD/1ibxwcROOSKQf
JP7gd1KqniwBhNjwLuv9ri5SpSRT9HFww7FMItHzmLgLY1zeKv//EpUqxcrQEpev4zYmkK8Ge2XM
PSZR/yeYZvSkN7GvQCWze71iFGVXd3VbHdLL//qWZnInSu3o63mnSXTfQRT6HNRlh1uDG4w8LQSp
za4ZSFUTICvyAWu0biLULVMUBq6GMaN38zG/2c/lMgl0yKiJQeCQGOESHYS7RW7AMZIfmCV3uf3B
DSc7qWwI7wWHRh3p4gFmpmuvz5TinSyRx379KhhcPt5APYJSzgFdc+U/+L16BdHDo5lzNAI1TIQp
EZJHG4SvzdtR9LoIj1CjS55R7Ci1usgDaQwq9OPpFaGSmDXLYz9tOQN5ksvgzhnolBc2PmS3FgH1
at8nh840peSa9ZAiWQgQry0dKfNPEi5P/uGyOqG41q1eHRYFdaVlGycsA3yXJjffHh8OOgr1xf7H
gw5IjAPidDivt8ArCL4N23K3bDC3zMoEDP2gp5e9lwGZfwmh6OwbmBY2cQ79ubg6msmcj4VQiY4r
+1DKqyTbBJk97vGQb4Ln9mDjPcm7iPE3MDEPS1GFEEXysZpNl71M6443tmpZaS6le66BoCbv0w4H
/vZIgNxwzdvZUfK9iVX2FcS7gcVLw8Qu654JXwKErn+Gt4i6K3NDazApFhlBEgogBXUtMgY8khBn
tf4XIKeeXD1j6CMbuZhrcml2P550ZqRw55EKxuT5dmWTEsNPqzwneG6MahA9ajs8cfxCFDxcFtWX
6+v5gx/WpSaBagzF+yjBHvhxoH8MnWyqa3lGGEjQf4oGW/qSSMLFGa+mvwLftrYVVCTX3vC9TWFX
o3K+MnFR1flR71a0LH6mKJqXzOwT5uMO7lpEusBV1DnahOmXjxrDisHhlNqLaOIZX5WYMdi9Gxjh
2bebYlmy0t/5eHBcC3REboTX7Tg80uQWSR2VhhRPH/p116aQwnUqyQG1sKXLUtEO34BPu8zxlohZ
Iz+qHyll4uoxfqLnKZJlRhYYTj2EGSF21zos+1sINwbnJnES7Tg8YDwpTBUv8UUFQbRi9zsvYaiA
/lukmTMm7t+Ie+fff29ePk9Qm45mvGMy+GzXs6TPqFV0QrJv1Ypk8JAU+3d213Lf9LWg5Ea8Ia20
evViK51vGq11QqrprfwZj+bzgVvGDgcsKSujM+SMkZBZ5CbOtrH/D2EEjcobTf88AY2xe3dwShe0
28IraVf1gXNSfS22ZVl3DE+JzmeRCc9s2cArXjgvHZ9Bp4MxISq+tZIO2vuV+NvyysWoXYoRT+Vp
3m1yySC/t1xic5f0rB4Y4SZlQIzpJffEfGnbnKy2MVh5gtinKZsZpIwex1k6mpKQewQXRW68dY+n
aiIYzmsDB3XrQdpjWhaYIYhHWDnL1340FZSX/Wa9IAXCpQpTf3M2kkJGqCNQHhYs9eRsb44ohL2t
tSJSb3N25JfvjpWqKYLimDhzXaytcsbMBZUHe90+6QwMKaUcCNiUGT+SFvWqR1kBGtUACSG6WmpY
wcdVj9lIykPpfeRQDVJ5NBv9crBkdTjQcT37R6VATw9we4TPzIlXpMQ+K7znPxwdtD8gxP5pacBk
uzJXuFZCGeTQ1JSR34vp6/CvuwxC+hPt2yDD5Lqe9PbrR1ikkvl4/YL6hnLZqsV/qOYP7+o5E7tG
yswg7qNHbClY7TGMLVFkRFzzmkyzJso+Je1ZlhKMz3nrrS/Iv4PZbtHjoqDcClDDIgWo4yt1AokR
t2S+kGN2VK83DcFw6gcHOj+XKrsFgwsdHU1UksD8ALE767KiSeocjxRYR2SxDXe5X4vk/36qbpUF
V8d2B8/W5Rt2VXsB6KTn/U4Tn0cnYgJJLC/RYvioCftrTTXSVoCjeAW3s9kh2eEn6LcDd3PIpojv
+xUne0Ac/XrrEEdrBxIu0JtfPw9eOkZgHb8nwZDeoye1weOH4LtPH/OnxRhuAoVFVYk8j1VSQ0ZD
wWiyS1on8R/kKhpY5TCUlqZHrc++o64IBYEdFSFFbqCARnIw5mgdDkUrAyFgue2y+/zRF9bHaqed
/9jaZtQiNiBS3Ufi36CQFuY7bXbY1OxUAVsCB0Is8ZObjkVPL+GetQT+gqYzjc+hgFiA000KPPOL
gaiP3Bwob5oB/GdJqT9/Of0lH5KpGHJ09qFFcOu/W682DgUjFqEDWGpkfqWVPW/8rtxR52dzXgo5
RK+roiN13tSvCaCqYAMkJz1a5vfMHCj4H4EgFtTZamNA9qowhBNb78NDsq0oLoiY+XlXjjxZMc90
jc/l+qMiqV+EiOUhp/6Ksg6rX2OEqT8rqI3DPZE44tCekodIYZAChabbNfYqAGB1c2wwU5MGVnA0
6lOBMmMqOioHvf5+XkXU+WF9FWlWskwKJUtJFnvTAFFzdZpqXPodqJMAnqxdwfW0QAMmh4SUUgwO
EMhOymcoO8sFy0Z+B49hAqjRVd4bYB+6onwOyXbTC5LnuPDUXzrZ8THLPkaWc9+VblRYWZemEH2C
77Kv5RlGfRgc9D9S/sn9sdtgDIzpg0dteX5w/didDPU7B2PSVMDD4FREFi2kMiqFaduIdqjMsBpd
LNQY/KpmE2bVd6i/zeWeXnJgwG8pIAIlWAYjuHw+yPLwzrGwKWNObqWjapCz1PEzhSKNv4+jOHX/
U8gp/Aydx6y1Pn7FO0849i5uug+D54ykTfuVwkEnjh6xgEWwgHGKOWxZZqP0DY4tltegkbcTP3zg
kG66ndylqudLLSdcOqqbtnQSgEkLl/kP6RMTfmHWSSh/fEdtFLjXIEXEZuI636TOgECbFtNRB/4b
ecVcmvaczGQMWSikbmnHj/QlKTx677q2Wv5xWC9uDEKB6ZW9mUYnNglblkvmn9wSO/TlyujMbl2L
h+K7c8JW9X2HcSta0ij3NQgLsKfRbiF958cDlHGnCYP2/mHH9a89SbKuHgX8jrqj9vlMW8hRHd6D
aw1VggBxLLwbHN6zWHRwQXSGDIWDt6BOvVDXDyeBq7Tz9Gt7r+I6PL+XGW5rfmErkAD0WZeTDyOY
3yTyTh57siC+vIqeDVeEM5LLzg0fXonE3LLt7CMGdBgfH3fC1OA4Q7lrsYZP4lLIUcWQ6G3u2eIq
Nvjx3/v7eUSLRps1+YuKHpx4EWJBWH8NpPbKgnoewyTgf8f9pAS5fb6q2BaMLQ6Gg49SdkQmkrFR
TyDflh+8LD+zB2cWklEXMPHVHl3VX9OheNr74R4WtB+NJLKNh1vkST/Ykgl0xEWiOfMYo/u/BQqi
/lfDCODy/T4ZdJJUBXVKc3ybFFMxJZ1Pv6/cz5s9CXSS95tkYzo0piyl7RUvNSGmMIkuqrLAmLPo
VHehzCCcxywSL5ZMIhBuz6ZviuPQR2G1N/7jLaIu0v5Up2DP/+ixZuKm465MlU9CznhTJzwHLT7C
Yw/fxTlAQyMGrV0AnmYRCNv4jl+QdpUsNoKkzvwOo0DwULrAidFIWw58E/NQuTBzJ7h88uaIZ/gH
NCSA61/Y3py36qHPbnGj5RPeiEDA/fAWIxJChAwY+sF3jCNGO/rd1KOm3inrcvyCcnJrmp5W7PhI
hmRoTmzLsmZNZYjoDq+oszOJ8mHGljUyhtutyLDQ1vtXTHEYowUeAYvB3x0+v9+k8z160hGB3DXZ
uztrcikCnnsBOQK4ZbCRFQTdjhq1d1D6KhDl+TryofSQb5BytCLOrv/EGIXX/IsJIqhKsozd6zhq
O3MGirFJW6ykg+VBG9fLSqASyoMwpbtOpXeIx7TDVV8cAt8pm2rlS1yDY7E8OUYeiJttZlNkXmMD
GilCyMybSwFpCjyB1hiXxF/6c4anndPG37gzoQiuiaX5wUa1Fcuml+9xl2vB3GpZAG8Ebl2uJhh4
Dcc81aC1ZmNYKfkzCHxNTAFA9XW0RVFiQtZ6+WTJidFKtOxomkQseVOy4/PRi0mmtIaXugDLBUhZ
V/4BGbz0rkt2gU/28Ixn3hTmT5z0ExpVaBu6nc51MeN++xZpcrxK4nku8in2pWEKrw8VWU/GG9fI
ziw2GPpWp5eaATBd7+O6OLLkThrC8bFPdsjC/z5yWT8O2Fc7KHwop9IN5yTj33iTKt57OiYAAuP+
++vnvLfVG7eZb4CqwXy9ci9gxMsD3HMdmhQyHTU20ZelZH08wj3LruuTI4QEOSQHHbdzt+THEBY1
8zk6pafJ0rcSUXB8SpEYJoWH0ztQ4KjAOC5u+pvwbiYxGyrfazgchsc/4Bc46qK2TDENppy/gFlY
vCRojvcttp/5tHWM54JsY/3LZT8V4jGZ0AmMWjdAhU7dEceqkp3Fi3gas5xK0xZSwEHYxikNhbH0
H44+tFsXTQacf53Zns5GpRsaq2uP1rhHsUF3C1cEVQzYLel2rJ1dExy2hjbdCEtfdHuXYn9IEsle
LP7wmYMiyy4H9/t6yxrfn+ld1CF0RwTY6jjYXJcLIEFPPBcTOhSJZSAqtapSqoQWrz4TfHyeFJeU
odZ2HZ7QvN9NA/OKRdQXYkIrVnP+GQjuovd75d2V7hfUln8nXNQG+NN1Aw9+4EcvfabQxviANfy8
3qPDBRpWmXgmwi9R/X48X9IXRAGQjgZt/BBKuh7x13hZyg+UyZ1JYuGf69wAkfExVsWWGwgfFHA1
OkLxt3ocdBttFZwkrC2Fd+jOQxKfQK853R1aNadLrK4V85ECQMw5xl4Ey2PWj2nt04Z8JU9yCQ4o
VPxUnfDRB7gEFqBSA1yIvnGXcYstCAxYhrVYJyreqXlvKpV/FThRsb+s5dJ4umoLUuCjmiOP4UAf
f79HVrpkxfInALXtaXUf490UUwiZEdX3DsJSQ0QgIcrYCabFJQrjb1GvkxSwkNIOnw3R3+JX9b1j
RXbM2TqlV1xnLzt3z79yD5zoVfVL84aCHYqrEQMErdKRhXIZylAeb/ntpMcdW1PqAieofyI4pnow
B8Xs/e9zOS5mBYgCey/xVYfUAVzj/6HtcDP/FZ+o+eoPfzYl5yx2TGZp0lfNr7Bf+IV4vDOPb9pk
LAxEShEJNzLeUZB4tOB+iR5vWMcodQW07ayycSbTV3B6mSKO9VuMOUaoRgFtVv4K/ULaau5N8HL4
mNAgpHdCC1CV8L/nG4xnYzOcO/rgzhumSnESNCiX2kIvwxcgs1YNdTzxxp1UZ2isvqa/DCC64Rqu
dn5LtqYXmAG3wUXnHgO/gEXE5Vrb4/OLPnkV8Fskob6AvUSY+9gUYmaU5jlGDYe8O8VCRmOQIKBC
SM04lvunZChaHuDIJ3nd3SS/eNxMM30pZqpxEaePrA+tVpT9vQ0Eqiq6sDlRc6T9pzy/RZhec3IN
3UA4yQiHAxMa4CeEhYfBp1Ab/V1VLAm8iJyGSRo65f9uHaeDigXDE54CaCD8z++KqLlNZdNCTCLN
PR2C9Lf8H27p/thux/a9IoM9FRyFkcVR56bytNZqyStFXmzIj6PoRkv12roefvx2eblEaIfKNlqZ
w07mh+h0eIDkKKo6zgUGNY7/FwWACD+jyCpGmufcE2PL/zV01ACIHLJeQqEhIw/kQxc+QZBrMVJQ
lkdqCpIUihtzgcn19Zz0arh8+2Nzp4BweUgBjLkaGFwgFwar7DxswhhHjDF5Q9jlGBv7Jc40/W9p
RNili+M0y7otCo6D2rUQgtsiXsl6w3kS84eQrDTVwmKs6ChApTh5ktASHMKH/v6sB3laKGLOkU64
vzvwxNhFrT9trVTD9UiCkKainqqVMS4oV4y7BTS3peheMK5Bh8g1jXPgsOVvCTd+2aXUbULBo1BX
GkG/ec6RYahuW6i1S9+WUla2dud946elQI7UIbmI7LEJdQju0ChPd3uBUAP8Z1NuWouiwuy8hgLB
pCLBPXQfR72WA2gfL6QjOjZGN8cToBStJc954n3VDmc3gaPpeVvO/UO+J/6CJ39V4017real+Y1y
mWxlrWqKSkTHsVPyHnHLPcgONl/wQvZkHLQTEVAPqrHMe8AK9WnkzC/DIiRdLDmI0TDtahBl+g4t
o3TOugsW+7R2INqcGYiiupcUqOBxWhCwGiwv3DxdDih1yDDE6uwPXkPkRtNT3QmiVKlCQyXnDG7D
ObAwJZdTYQOsg3eRSe5WjAIeLhMhnstK91906XunGA+pZgmKrGYANIDsj9PEWr1ilCCYIiVZ6UUS
e4pgOnrZMNzp7fYNlaihapoRJoe8+nILnG243Z9BF2eSLVY0Aldp4K1L2jXRNgwUy4AJWHAlUBKl
o1Sr7hWNgEieg8sNx9UkoSkKTRBnNuz8ljE7cLq3ILgXwkVFSSmvfIWMGVKRnRg+TYoIgg7as8fP
HUnWg4Q61/oerTmQfvlJQiuvhF6kT6e/hFJVQtW6vZK84dqUo2jjU1VRS55Q2f/2Zn7tJy1TdCzH
pME53PZ2PWYbxn1kZ2ZO7CdjuYG5xh34VZjtKNRJF+VLNRzxPr4xt0jQorYabzZfZz8R3mWEmloX
yNzsROTOUedASM4sLVsMpYREgAtW6R441PaHMagTB+t0H0Sh7Of19unKLpRaorH69BDLTL3ujtxD
Q5s2Vkq9SJvMrRp7/1XKoBssuGbpqzAgUoOHLDV9Pd1h5tX4Y7HUPsf7KkSYIQVOoi4Nxp+Yb8g1
Nd/zZWWDwlO37Fqdv3ErL3XZRLia4jm0pKbYHCXMM1oh8tDX/hh19j9lrIuJgbB053JaZ5oX4K8W
cJIkU6GR7oNzkIXQd3NcLZvWdPLUd/ROc05ars2ELfAken9EIcof7aUupwODX6bemTq8e3owIqfG
Dyiud4Wx7GoAhTkphhMekV9svOz3v7v1WAhdEkANnBztyndukFpUwdpqU7fSZx1gpPhWOzr2RTa2
EdmRATkZ1tN5GsNve4Y2G64AMDqW7IbbzAndDKjkc/Xm36UNSeck5fWdm8ZWTHclPDoDqmMbqYN+
WQxt4lkhaa4eOGuoR2XOPff3Cibk5tWmGATBJkWV1GNoULk8KprMC72Q9r0T5/Q2hO7673IE6cwY
0WiGVUME3IS1Zd/e6tREpfddDbQ/o651+JgSoVYHvK9z1AWilXy3QBWv0SS0McSqpdpIaxnbBRyd
wBnSPzGuxtIEGFVc0Vb9tvq5BzeunHAgHMa7HBTJ5jAl1/tqsXcSij59nH32qJ3eDYFTJUAlxzCF
tqAB7Giuxc07zHtWQDx1nme4MNwgENO6zwSI3Tu4w+V8sSIsNFfJPp/hK8iPDTF6D6dIZqnqpWiI
E1AwQvhIn35iiacb40eIewAR3LNl0ILSCg/kAnNOViH5G/7AcxWSWfCYFpEHQa0BKnGejWGJmLIc
2rtHnsA+pdMHXFgsc/uytPD1VqjzgaxzwO5WtJdhYek4QJntZyXWTcmYhFBC5l1yYd90xpS0Zpen
2ssE7ks6qFHSjwvrjNE5ykCTGU6ObDqSuR89LLYHgAXdgvS/WB8H2Yh6AlVfYMLQ3BEHHrlUo1QE
4+jkEfd9SSEw42X2xsDxPR+vXgTQCAcK420s//woy6g7qF8Qgg6UxnO8mlx0T4OvK3+onokQxeey
+OrE3cJI6ZBtCk7csgvR7XDYvNg6oFA2x6K99JygUW3EqdxTmT1qcDwFp4S1bFfJwUF7WaPpUz6u
tct6SJaHp8FQ1y/rnfbYYXMO8K0tOgh8Y0/aAQBfJ6ofZmI+Z+8IKj0+KEezNbqh62NdqBFPJ3pn
AIsGMRF/zxs+fnbr+Q1mSqMwNWzxEA8Xpf6TTgx/7d0oVzMT9MoJpKsE+cRKBvLI2/iJuweZurwe
eoW6y9qJS0krWPeFcKU2vUgEaX1jom9ExX2oGiFH2rDroJmqFrXJ99EH2RdZty8saaiouSzetkuH
um0n1/WBvxatYDc1s9eq2SRjqurRexzQLwHighcM7z6AnpugIDiUUGMUcnoE+6ZZBHyTNONSLbFZ
R8pp5ac5EdMVwkDzeG5Jdmg56bECoembmPfDxZ8WuFj4k99VgxmJct5HIiWlMBSFK+CfhJlnN1Ko
NwcZbSql8GOoNTS/aLyv5nXGbq2zOQCsmy6hiHMCYVUrhgxXuNUgIkv0QkITqLcVtbiIRaX4fyf7
ewjykhkMQCeMK+jmUwVqWC15zm2MhFnKG7Q+bFbGz4fuzC36fadE3UU/HUY2PimFAArP50hYWDCi
X1ZSAX/dUoXFSzhEIxu2oYln+NoAv+NV8vsTkyorSe287muRGLZ53HSIXOodTnxZYzpBSgNP/BOa
tkxr4lUgY/lDg/J50d9YSAmjHOmf4QWoqxtg2Vv9/85lknmGOUK51iiKrxje2yglnwJ1EOXWx2QL
4VN9hFXRrfccHnaLFojWm8d2x+BIhqaEh5PoSv8emv3tsdqmQdQ5JdL960dk6fSsTwz7gCNN67ev
/eXYIWdWHmHlBJ+3/2bAlT6DQmm+qctB0CrC1p+YBF+Y3t/iysWGI4Ep/fPd13G1AIC4kKkTak1T
ooVgoiKcsx0Yo9aq8Qo9k+Jr7TmOitcdaX462KBKoXMoaoTvd983B9kIflXw36llqH4cAAEpYGrB
Bg7sKSXGIYLF5xm4BbFnBY+3FT1V9j9PW0Iuet2FnMQopWCkpQ4F2UB1HzbYvNpkijDfN3W8se3j
qxnCkUhM3H/SJUd7RvrhQ+qIWNo0EO2O+BACYGsU5u+qFU44MVlOxYaGYhD0fHst4XsIwTbEPGsQ
77w6i2mhsfYuXEg1qJ7NBIoek525eG7wrePDTTFQXTskkUQzfjG5g6FC1img0ps8OwtzQHA1kZqb
v/Bs/m4Q6g/v/Y7qDJ8ldnlKnGt1jIm0IaIQKNdKxLPGXpzr9z0CYsaA67X+E8edASSpqJkuAZ6f
f26XG3Rzvub2H9RuQ3ec+3BogBIgdM1RzW6EppJfnKMw0jWxCsmqXuKLmfpCRBom10y5Bv5Te+bg
kp9qqAh60qPVhA0rK9pYfQEAZdMdifPr4UVV63AxSYckbX7Mrdp5ARRvWHvp62lXVahoXBlHQ+Gh
oQzztSAvH1pfZJU8/t8PXtdMdF3+Y5l6o2W3BNf8noce21fpErWqZqef7vVILFzqJHpllP7vlu2Q
O4Zbp9yZ0rmxG2obEgEd/NZnuT3DM0Na6FwGPxSUUUqiMN+JnAn9greVeHadl1rUuk8JTvWSG/gZ
GcbjuvT9VAn0YeFyumAxS/7zf9EU1VYrtwc59rt0UmNx+3/bAWcaNaWUb7wfQrCM2/iyb43/YATN
u5GdJGZ9V2dXF7VFAmSUdpTjbntsMiw/IwzzzlBnzwpvVNs1OipzyZ8Di/DWo7fNGN4orKVNrm7x
X2g5vFuZ6qikCHYa/ioOr/IhRiBuijlp3e2V66Ro5rjN4zMoBTHq6AV6J0OjNnX2F/QPkEusceCg
CbTAvgjB7IKcUl5v6A8/jDpZkBwG4EnzWAiJxQ1zuCJ6fu6DpgWkrBOmxgFFz1/YdX7B1zBNFPZw
iOOFnkQ00yfW6gjaQuB3Ybw9PAloUJPTjQ4pt50NZkEjWrZxOeR46qYKM0UOAyDWU8dyvtNLO2t9
uAXAkyat9GZR9MHOwfqzAzBIK/gwoJ8IlQcYJsVtZ3EpaRMAJqdIk49C6VrR/B220vYmqsolLTlU
Ac/ypWQlH6+rc+0ifnmI26KD9LsT/L9K0ovzO/AX/LwcHRToSfhSLbw8Q9lp4HBm+6MFmOmn5jKQ
0aOv0/QrjrzIMfZ3fe3y8/FPv7Rt2dkJh+Cxag4U1lLFUw8qAGJ+u5FAzurvutL6L9TyjAdVbjVI
GiclIkTBqdG4rYIrpTpNdgHN8UgN1QoKMP9pxf01BoYLGwIQ9UyPz9G0fNj0xUrijZKNRh9gvjWI
tp9cbSiFwnBLpunUDkt33xyt6DpQm3t2hsgPoavIuIOly//b44T4yykTrabmHczRohCJ+aX4FaKi
QX8kpaPIkGktwp2KWBvgteqQfgyRy1SLKgE2Ll5KwQetcMxWp3xVyYgXvNDzQzJccuayqm5b1ODp
DZLJSdRIYNwHBfcbkKRxPZEQ/coyvDGUJClFpYaU1B67lVpfYWoBk/RoKv8XfqQofbuHS5EDUO3R
19MetMi8ovBH9sEkRhjLOHK4AIKrYnAHmQTRJC5y/J++qiF6zRqLDHZ2JAQijq0W3TR29EdGlLjs
tjz8rewEdrxah8L+EzNpifO5CjD9UlUn3dQggaVP0x8eYpXsX3UPOHFzGNNfOuk2e8rN79dV3/gj
8CzQS3deEvLQu3GlEShd0ZVQfbrgGjWmX/kwUSbsEwgzF0rWWvq3KStnzHXfNQNqCeUeefDlw+8H
utVEOn8bjGQJaC4faePbJaDibgWmeY41jHgRtABUsxYuSTRE6wE9gJK5H57/BIn9G0fFyvWIgt6H
L85etT8JqAAjYcwzNh5PVJhYBVdpmQjQwYzWClzJFCqdU5imaqD7slKi2OXRFlRQi+iOJuSuN2NO
G+YCXUDSClFLAaFB9sMygzigPGG8V/DektC9K5+MhlG1LEMGBrYXous/sk80Dc+qUdidn4qU7ehC
+Q2uSjpkmBaquSsAQe+dXkvcQON/D+mSULF3RJ6brcnwU7LvGFVnZXT8RlTc+oUb54vWVXAe+BUM
mbEYiAYMZA5Uzzz9wEKqy+K1dauuo3n8dbxndvU0dE91YKlK3xHAQNn0gd7p8RsonKVeV3nszo4M
/8Q+QSohuSlj6kxgUg+qHRJiGQk7UV1Q9++U5VqsM5HAG7kdq5dzXxsJwmOEB3jetW7EvzkznpYC
jSlyW7DCeFBXxFt1iVqD+qXUs4hHiF0b1SxvHfav1wN+96jmxRnZd017GW7babp1bIN/erl/JGZn
FFmHWxysFX/lHMPUCSVtAZqav5qWZzi+SOs3FNbQ8LPRlpB0C6FIu9Jr3gkRafWGtiNA8qIlZNaE
yUyXNT2bMwAZW2HsFslxV9U5tX+533xcKF+eU5Pxvwr5hDrj5w9JFTx9kdZWBEeMxlDEtbcK0LPu
C4b0eO88VAb8zmuV2xnXE/vajB2RwMvrteqqsRCT3XBHv9Jhc4kl8fvO16KOJU7IAyZL4mhJS1zw
kfQUGpns2ogdPI1dLkHjpPUXowRGwJChosKBsRvxc2IASZI/YdBVbVxM7YtMEO5rM4qdXpp5AWjf
H6Z6qMtRGQCUsHPYtwx/H+HW7dE9KAHrGg84ciwjax2ayj2QK28q7BJS/M9PD+AU3i/RoVJDhDeh
NsQsF0kYv/1nxHBFjKJliYRCkIKlsaIedPbUgdtST/NXb40NbgSwOL82luXoI3zCTeuQABisQtGg
nltacOVrcMOByEfqixVGIRLWeIPTwnwdmq2W915onyA7RWcR5hQ98bUr8jHfPjCvy4ePiHm1neHW
iM5SIiZ9V8L/4NOor8iDvXSjJSrLSIdnpPrug7OlEbfack5rmXucsmjzBrvfKutVz9p15mhtqpuC
bnQHhEPbRJfXABVndWP4HGkcLDhWrIKgooUm55/nuNR8HufogI3D9AKxirY6E9m31K0FVC5KqkwB
yRlSfmZajopl4cGaGltZJ7sD03bfXC1tejJWRCtPT6ZbuJ6gY0YIMZsrfZr2JL+eZnD8OlScVv8O
hm/4jZnh1aLBn2kMpb+q8Utv+XSiXPJc9799SmQqsPyxyh3beVTfs/4gDDIFCTLF17A2Y5POqQgm
eqy6Lm62qkT/DQIaDLJR+t9DI9PUJRnHkA8wYQz98MK3QQPl2vbBLtV9dj1N4YLl2+32LRSuS6/f
iAs7obz8yiqn03EO0soL2IqhReGjlKVaSLXBYgWpA5cWxkEg03a+CgoD74NlO1mKqPgDDt6RT/If
pYeW6LmrYmkDXbES5SN10ow9rJueureu1nv4y3d3qcCsKycJjSBHKJXolQVDjLSmNgXIYQ/b2MK+
C+X7xjUUsMpIQm5VYKvg5iw2SVVw2zBCZ1X+a5vUq5TXZXbLvVWou5Ybq3WnH2Wp1VunhPINvD9U
56e8Q+gR6d3nimpzqQjNUR1DkVdiID2gMDBLQGVzsfO8cJdZg4FB1GvskywMv1oRjodTFvTT5rEV
XBeA6n4O00woxVafB+VjWhWgzybw7vcCc/BFK+lFN8Gm4mvI+Qqizx0eyORG3UWSiszE4LpcX+/g
JzscDSmY54NVU8oOC0+IlMFJoj3++iknWJD8DYuK5DeUNojf20bxjN98+oy4sB7nn2+ukZbm+fkJ
0GahaDTdtiOy4JWftxhfqTx5oy3YCm5X22SZewhq3wDJUYIEdy0mCmL0t9HrbrJPedaD3t4MRNgW
tOaRBd8s1+3tr/qgozSVMVQ9iic1aj7fVeMPsbG1RthWHu8oBwcmnBZuVyFiJ9GAnRL0oHsHGNaA
idoqNUBjMvJ8gOHstVY1szSQyXH9QiI9TbYMBB1qogOlsWDcC9EDn+FqyB1hmN9i+9dDSigP02OL
JR2MSHMjr+XxkUcw/eaJvQj+zw/WZAlGk7KInjXAXVEKQL1eK/qVjoBAaQqDngCKmqkInOEpNQ/H
NPwe7uMbyHra3JPq6PCHWcbWo86mLI9aP6aDUDVbJBHZ8gMJWvXnLj70qpxKFZkeIRn18wZbY/eu
7V+i3HmQwaR1nHujWa8R6Zqv2y1P9fqBrGSh/Y70abrFzVqSu2oGBTvRDDTZPLCGXoWRu+J5yf+a
ej/ua4Y4dhM6v57eoMYXF4OZoJDjzhMkYknoYGqmTxz2QtYllz6x2Hn4BiFZBa1TpkfCfNKRIlxG
/OwfVlgdIs4RDefKvH7LQWbtqlCEAwolV+4b6Awzc5lC6u76I9MWckB/Z8hwu/bmA+CrFQ2qM++1
Vf0UfxC5C3VeUANxnaHM0vVVie7cHNKOahZtX2SQNogQfcVlu1OyPVKDYBhp6Eqh/qUfuslXGnn+
vzvm3sCNPxXRO/cc2vAr88T6wLxSmP28Qy7Cs88Hh0ErAUsg8DfuOUDTjBXwrxqBXcoi4A6KE7lB
+cIzBxrfz1jkgPtC2KYcOLIMAEJmIuoblFNsG+Et1f5iE2xNNqAxxdRfnsrrVEaDNx+SmqtpAHGc
or++H7a85/UY7cGvNEsA8130cURa2zD6FB9ss4CTtBu4L6pgZRfyTNMmVQKURpO7j9YO1kqoZwoZ
ata3QXEmvGQ0nG3iTQYYaOZM7F8KM7l2N53WB9BEniGxQEXPHVNg8kp7hMsUphoo4Rkcuv/6auFE
2OzcM9iq6BcUwtlaoUgtoCTW2haOoxrHwpdEM4F8Pi0Pbb9dkyhnaVFHUlD7HS28Vv4bpmctnhVi
Idwc25n8wnnULjRV0G5wTkKh/2H29ES+Kb4F6+GbdH4eWFQnvsrXxdgUddZ1GdXqSxjEbT8/yMHQ
cce2ik2foOCX/DfJEJE6GVz3AajZqeE7bK+DVM2HaSXH6xzeGVONTKI3GAdsssNpffqeRMBKrQN1
dbbxziC3YzMbd/EOQw6pJEbAbIm6QZCwGVpc5NAnXzTb0Ug3KyWZFhLZGMLCKcETZcenLZNO9vEs
3bvMV+Bkz/ZHDCziI+GkvYRGx9V4YfSCDS9IZyPWu/QmEQ+fhJXBUvBm+03uJoMGDQxgrl5rNFaQ
2+eDQEHpuZO3g7yQbEXQfREP5Y7Ex089fpmTin0nii6hmdIeEX48x7RdpwaTSVjjegXG08352v69
JpepaqW1bKeA1oa6q1PI7jRSa2jCFJGOJZY4mr/czF7Om4b49g1WdDNzmhnT6dfaHwURfFRcghXr
u9Ssv7WXXxV+kOb1k6ze4YPD216N+J3KoDjt1jAkN0A95muEIuHid3gYlAFC7mSFAUTetrTsf/ga
mzOM8GzAoQIJ/GxS0FsT2tqx/rKbqSgJaGgXQj+fAJLcgMd4nmYbl79xyUwLhO3koh4OUt+bUNos
p5juLg0jGhhW9kbAICKqtkBTxBj4bbmF43ernt5nnQu/3+USEC3ND8Y6Gjxgehi7RfNKtScbT7VK
AVquK1BvyxZYW4xZvcWLUR5/0D/OKXG3kU82AqQn9Ig4/dqEGgJJApREmeWu4T8zIO1bU1Z4u77S
aGgHivw2c+8oWdfUVyukqkvfZ8ZykPe634xZQr10vkLjzJu7h2IuIRJIi1dYFy8xVL+W5HFSqDJU
wRGRKaSWdTxjQzyhmi6IAVjc3rv4ta3wd0wecJZtxym8HXTTU3lJZ7KLzV0ju24U9E2XEMhruI2w
PS3RUrm0KK6rVoOFAW7cNsIrgkKF2mLn2Js+tEhd6y0T7Ezraf5SexbYIdBd3lgfCMicMdHT9FqN
27sGUkF1uEsJU0pziHrJNqlCCpPdprpSMHYVWlVaM03XwB8BDiaU3qX0e+UiBxaK6UeIizM9Gvh/
B2CIsoPmtg1ihYbdRthTFAdE7cXtJ0SDy/T7XMnRhE16+1RavI9ejsL7AM/KsTLpb6lLa0o8Eo2k
A3OXYPysiZfF7siiyoNTOVv7Cnzte67VXSSafurHuNpeVpFFEUjZQqVGKe4IBjkAUrD+LvfOVL9H
o/iiL1hXLf/Jnpt4Y7BBS+koIhF/cINMFD/lbavrbkQMKixX6jNu7b6RD6B802iDOkoCKGPV709a
doyeZwtZUOWLX2k2mebJxOd/LGkqXftkCR5da/WiHat48zIXRqCbgCp7PbmQF1QKql0GIK5WcEyH
Y6o55+3VYhoh66Wz8/f7YfIouYPDZoTV4Aw6jR5YFU/8xY6PkrzopABAcR4bRbNvWsH7TsovBDni
dlZwg7Lr4HCa0IOj1moujsj8lnSNoHLnUOQsgb28nunC9PPTkcJe/lb/H0buIb3XcVOkUdUW5Z6O
UzsYhJzyvRJ3cd38+tIZrL0fIdG79HnxRwOhTRnic7ubkPriVO1W2jYXOh3Nqe95zHsUWJ/CsQ+X
aNa0s74CEbc/4cmLGWBQQRLv4ALAhSheJz+hBMTgcISlmzq4E+toK0r3nhLC4hiVKI5CnuHOtcz6
I5cdoUbO3FXOD/KMjGCZVACuf7L0RfKcTW2aQU/CBmoH/j+NRPtCFtaCCTrDqYXDv7kbSKEQrYOa
VT5T+tqa83IVaxi5G7m1Qw+jkWKdU7/AOEcQCcC8NCEyDDn+S0V1I7rxH/5Wca8+qr7Yp6UYCUNr
FybTyXA3zHGt0hHQ//sGmFj5u4+oDj0W8SPT6kYnJ0wkwAKJk7ArZtGnkVZy/ExZQi3DlB5nLBu5
Yxxsl02idq19X6H15Fq5/lZ0ar1yCEYRwFdXGNVc45B3kydqLxtq9x/V7CKQF66rf3+x8KfS75ZS
NYahbat4p8WwyVEJpOt5CSlk2Tl1QDL2nSMzP24fNjsdVDrqvEAxFs51uGpCowgp6SHpC+XO2M3I
/o0q46e1AzmPyYphjEYvvV3J+WMq0xmCGejwAFpr80JH8d2IcgFR7seH2EpU/C+GWwhEekzxiwIn
EencESDys5gWYGEYFsY/5pPisTMQ2zKypyojKa16YGsZoOYxyEbz5MmRWhMO1Tf1rAKPhzVBzBAK
18D2bOtn1w57K+i6ZhMUqFLfxlQzTQ9Nkwz3dyMYJn6u3cXfuhfxSUR9unyEEwT99ym9o6B4Ry/R
3v4UIIO+RJQ9W3lL869/IaL2gSV5NUHn9aAeGphCMqbLvoE9qKNDT+p6/WW6CedboIPme//7NN5w
zsFPepbK6krDY/U6pkVtAP2RFiPTqPAARHUUBS78JU2/9uwjkFn7a+Utwyv4LFtLYCxXRbg1ytZM
8fXmSe8rFAeqg8C/rRs3EM853auQQpiR/LNJfuy37qiLGrbrA53NSkpE0J0Jc/GBqGWd/SmHCGG0
hPyYhPhU7Sv7VvW8R09tREhcJoH3XmawV+d+h7ZoIXo+2Sk3lU6p4fZfxx3vi1WRitTY4FI169KS
xEFIDx+t/+ag3vVILzQahsCrWlhk9pd1Mz0IqlLMn0wzKczBEwJElI88TpeZ8sG0dQgNgiOY+Qm2
iC+qfPp/wGhV+iny6LBizAE+fl2w4SToauByQfahih3AFUmeiNiXMWH0NbkzkE8AThftuVocIc6a
jf81ZAC92n8gFQyvwBaFnRy5npx8j9wnS1Wy7/U2ZOUjNylIgM3lr14Xo70v2gMKzWCroFTjwGUc
R2vzjrFdqLCjtsmMjyxn5CHsZb7VG8/YHfTV87uy/5gu6HR+AWyZdV9tViqxk/HhoiTihXaaH84B
4k/7lXMp3UuIaLzXxyFvgnfwvBTz9XHEOuZwI3aGPrQ6ppXwh3hTGFx5SlUqNzxYwuatmQAVnfW+
IDr1I+WgZ4fyskVz28uhiulux/uD2LKBxezkmooZCYYGdnBmiyEv5OBO4KAvdzK1zhMArLjZizCI
PMdDOpWGIJcKBP4vjeHWSg+CqETHtFSZLvPMBOspMf/px21ZnQuhMwnqezTSHbVbfvQXJZW0pf0a
iJaonVPlYwMuPB0uUf7jwDvOU1frj0ikL23ikmFw58LC59LuKbojTO5qLgPZ/7QlOBT1zzWx3WOF
h/EaK37FxhQq+7x0iY0BEDqWoeTIsU7EOtqfXyU4XvzGHPaJBrFCpdHjGVqZFqPtt+HKKz6QOqQF
LglLUUAXw7RcpkIVI9SmVxuA/YaB0tsXYEvPLlpP3AvQfq/XBLix5V041Bnu1/YOnhdTWk4omcn9
uxY1NZN/EoR6jVjqsxg3BTcsn+V2652wC/tuoG7ugwfOblfmQ7YJ+RKfSNUIIAqjM9o4Q644Zn1Q
BlPpeBV+rEH6qNN30nGo8b9RaEEUvFlmcnzUQ3SrCy9mcOQKpPvUe3kuKMWgOzwgIBTo2rVJ+ebA
J7/ZB8Uba+YMCc3xe1C9Ivlv+cUR3YOFuMzzP6cB5zgkafaDmalwNpIsD92tiWv1hDOKxJPbOhZq
jLN6/2C5XTZIeNWnvahn1ZFupt5VIspwnIn3nnyYFtvQtd4LfKfcw38e0eEosUeMNUAfLeA6uYBC
ZjJOsRd/uF7Wn6Audh+wSoV7ZqL+pTVmhzBp7AgfZZB7a0/Ojotb69fzU5+H+w9Z/D21kFLEVXDM
xW81xkJKsx1X/yzeP/i6u1FLki6DMplDJRxYGPaqUk3DjUUqfBMgi39yXKRF3QqDm2M9cvPAyYzj
1/x1oBhkFaessDAkyH55yD5FmpVe0V+dJmBEFyKb9CH4gz2lT0DPmICum7T6Lwkq1Kp+Lk38Lyye
78PHcGfdntp5dmWWqrWWiwSQGxniZvDgMTEesbsvh8U4Xpo5gFN0Mm3fll8BU82tkp0LvXrjjOS7
0jMLRgVfXg/3sjNQjw1fSByoXVKRMW8S8XjDIz7qbdGkisTZCimWZI/BltXTT29AbFkKIj6qsTFv
ppyMgExjVceNRttPMi8Gq4NHxDcJZ+XHKkmKcO2vU3WvLGOo1xliHYYo4spTUZNINQ90lYbbNxdU
2GNAQIYvA/Z0rcTbxxHkX4kk5/uANydkeXgv7XjTjlqR+YxmtgBBsKLtH+CX++PhWw2N4KDrjlpf
bJysMedr+U9BKSDwnLt8TT5UG7ElBkTMBmcflsS+cT0GqQRgn3cKVxpYZKe3RR1k61ywDn16MbNX
x02TSWbAud2uW+Eze4uhbHy7G6nsPZLo527IgmkgOGnxULMwtH1XLsVd+ZfJ5utOWorA46yhWbjK
MJRDoWtV/nejFV7duMcdCPYZ9o5w3d0j34ZD0NPogB2n0oEJ8OCqu69TtP+FDa8CxX9zq2lBKD2o
8QJQ3F/Ib9t40/GN+szG4XKrPFRv8FHy3fraO3D0zi+dBstsRAdN03Dcqhb4RWZQzantDjGCXMCi
tQQY6pMTu1dpJ1QRG50YPT+r24/9fi+cQf08/boCWaYiYbUQh6A6G+mAwXnbur3RYNtaUCD3wuu+
ionN3AYos61F+b/IE+uggcqJFHiASR52Jn2Z7ccf0XDWtBQCbWeWesInjaE1ecttw1n0z8QsszRT
tnj/acpqMD+GOU2m7XQsH6dYX01o23K5LpSD+KvgCWnmNW+SuKcYZweYTH0GpsCYffrqrU1/v0n3
Q8ufP/8B8XswZVgtkmzRKWkfF8T/4M3J0j3KDg3T2kOEB/vw3bPjKfg/LvYPo22tcR3vhPajq/rS
UBlPx3HHoAKc/oB5e0YVr9IR+/RynKcvum6VM3M/h/herHbJw2QT/X7dwS8n8ik0pYQwizLxz86O
JnbvZOp5qBVR6c+7FLNxuSw1abDdjFRwPVJYeekAz6pS6jIosBU/ERwkl26f0TgSb9g0ZyOxY2CH
tq4xIB+4mFAbGZ/5wraCXnKEx1XIobEwyUM/KiuZxS8x7DFIGaHyzbD6nZY1oTfhr5yk+jAOD9HP
1/j2cuW18O9mkYZ9kJYP4HSp1yCGV/x9lcUbLmUj7IG3An+FU1zC6LE2ObIRDCgK9Gznk3dBtn61
fUhZRARr5UsNivIEWI3RIncaz+95Cm66i9gTILII32YBF+1i7aweaHO1DkQZucNIBILqMs3wVadG
C2uXKtIC5fAWxCFW8SEZldMM2cE1gnwhJrsZArKRH2vJJhvL+sWt4bVGCwgfiN2C8CUOF4AZsVWy
dE9o5idj5N/uTpI1alZfovWX7nobQFXQ2bAKhUeuiL+gQ5WzIie2sgsCaiP+OFiQVpKRg+mEOeev
FxAtKj47tktw0T2bQuL7MsMDB6KDtX4S216e0UbzrYUaIN6oBrIp+e+7nBxMg+CeF2SbX4j3bxQh
g/l+vSWI6fp2TsNDnIeFyWVs+HKGxEHr7gOqVo7MLcZNP81aBeIDppkaheJ3KjV7vKSaRy7v/iu9
fNklU6anulv8xa6TJr4z09Rq8aJR+f/+6c+zu2iSqVz2eppFubTULW9YGV/biZc38JPWB/638qNj
rex58jCyx8pf/FcdDVFxwOXo2GpG4gszplsbMvqXnezTg9yHdGMl+nELdCxnbX1gNRQhC/ruPrnB
StsSbsO1unFSQKHqSprUTP4vFaILqgqwu+b042zyctAwDpcjQQYLiTToByWIPs0qaRJx4KsApkKA
BO/yO5YglY7wMz1Itmu2MHLlA1QGX++RFwU6Ou6dsoSq7ixf36ToCQnHeLEDJoDIiOSL+B/fU3KJ
fYvPoesdQaxFiIuncBtJ333K7p8gGY9xWQvLtAZjJ5vcdG6+oLNCVFd9TYHc73HqJoMbNTHQYapE
uq9QQh5PTnLUT9zQQ5duzhiI4407Y1I6MGej5Mhojo1unRnJgdEteB6msLHC44rAc0qSev21FaNT
+O7YL3he9LEX8+ph36VTz0NpT1rtW76ZhWxF03bzSCAqS+0UUypqCMSVKtXvMNS99VeaX8lf2j4P
YvzyhHcrult0CPBHXp5plnmVYKdMgZnZa7qn8tWpoRcHPwqsp6puftg2dVVoqKxWaPT5/vUCBy83
KQFluT8RsWjuAaEaOOPFJCwq0HaJlH9J93CDuZfBeUTUlTedLayiwXVjC/5WIQ6MYRbH1GkMUOLV
RmIFsztfEDGSiIwWhJOhBVawyyoqFLox6CcxopK3knYFTKIFHQryq25/cM09H3E8V2ssiro2oLF8
Lexp0jFhZ0CjzJaTVxA3C58buMaFewSW9seaJatQmubq/tqzCNPq6v3a8lJKIET8CBAY3TxsZaOq
u2FJsopl3APkrhfC4n//KOcw0W7Wp37xP8GicWlZrK0j1XQuL3T42uWmknb14HITiCwDpFDaW+aK
8b4Cw7xFw4XajULGVgmzocJFhblTkVybXbhDPuhEZZ1ghBhWb7J9VVE3q2WoJ25X8s/2uYe9g+av
YA1yc1LvDOxOJNzvOeVosVQHwPlqG/sUWqeRGmbV7M0193491SITGB1oYSYsFoDtwkcLMLpBX00e
QjvjTYypxghGMnaCrUWGCseYI6iXAXx7vmz/K261cIy9SRKy4st5CI6Dor9D2VdhejsbpEbmebeE
JaJ47GXwe0apLZu2556PZzIFgvCZLsVP7WsZgyHLZ22INHuBvGF/w7dApCJQ23Q4tUeY8GFdBrwN
6o49mzT80KEbEcVUv83oO5bQ2Nu/W1fMCWLd6sWu6erMGjc77kZoH5tL6qPRdr9kyXw2BenOodVP
4wHA+1xOoU3L42ZHhqOgf+O6IAb12AHmqZTUX2aC/TDnedvYHEgCURBNic8/4uEE9m6aiIr4ibmi
dqwOVIqWJYwOAKP3atEtT+I7DKo6S++Iw4OKHaZbK9E1PL0e77dbZCu3kirS+cz3xkXA777fa4ll
gsM/+RJbW4+i639Pxja1NfrdZ9xnQYTJn0NH2/yOga4yDD7C/tCXHbwRcKDJ2T1TqDGtjXQhYDn/
LVQ1i+agin/HiV3mV+XQFAxe+NKThEN3Igz6gVN8XVkNPKqjH4US6UDV27FtPmE+MG5z0U9rvsns
J1AV2Bapd+S+bDzwqQ4WvBQJ1wEnPVQLkYJn7rRUih7TRSv1eBus91/AiwiIavAk7BrO5YjZh4qT
xlJAXEffDfSOyCDnEzEhDu8DyZU4AAttlScOHGQRB5B+ipE9DXBC4SKGE5GMc1P1X25wwXprcPCq
4ETez89bipqvAp5rK64WSOsg/JzEi+UrLI3uwcWfQIzxb3QAt5gjJm64/uZJeBvqttYCiILtzwQU
t13G7HBABh0C2otqnRxLgMQUO/Ugj0kz+Kq/e07Hl4xHZ9bfWlvwj21M/dEhYhIt4N8bRnm05GKR
Eac9FEMQ0tUd4jy+So73x6062lQjUSYEQ0PalZJtuOdaQJLYMSwc3u1CUhg4tK71nUK5waa39sY6
VCXBWQw7KcH/ISV/uJt8VRH3ouX1Km19kjLkydwpuBnr4dKCCB5rSDKZQziQAJKAHszDkE/4ieYa
sd2fsBr6EI+JOXvWFrj3STIC6yo687XEJD3VEdr53hi2sQURRuNbdxm/SOJI7aOFwY/wbxam7QT5
6THYi0k+Me16jrZQ/c96QvDS1hTyYzbcQTYTNbKJk1l+Pt85AxMhTGkG6iuBSQIOk7FVDZNYEybx
rh+Agrlv7MwEYG5DDzY6VaA3V5DnoG5XFF0ull3DuIiAG5gVRMSV2BXEGnbjuATBISn5lMlBTAz5
07naofXm6R5+zue/iDSP8pIFs5ewswucs7uGy5s9pjp+SJdKcDvldYFBCSwgPZsDNydWO1mCYqUA
hl0oQN59QPPcej9YuU70NbHxQhZoW6ToeXeaYj6LFh6CNcRTD9JHhXPGBrUss5FZlj9oGBRbQ+lT
39jn11kcb8IFiKnA2BgV1nVijcXYrq3hqoxJ+w0nLgn50l2a9Z5SPuYFYJIEvnV9pw+YDvE9nglS
8RhOSuHOhnEeLzorM2E+LjflGDQl46QTekzL5sC4wk+oscUzdP6FV7NL+9QE1U7fTCfYgrleQFCg
Q0dq/sR9Y7MbG6nzGcb0c/CEvYMSUv6OTCTxcrcNSQWM8eEQEYC4W8yVc9eSqHYkFyTvqpRuZAD2
1/xfvTLIseI7h64qK2uhvP5fF7yJKSqf2owgb1/s5iTULM3uDEr3GDCrx/XOOBIjaSvnvYcssE0W
fnm8JjNaJfe1MT56bFIfhO63U8XDbTSwrdKr9+rIpJMMvLtc+ZhOzlfiG+DmqLNyOjuarVkHf4Ei
OCDiRVZv/5cGZEXUZ86FGWQ3AI1x31RmcNqgqbItLJj7KmBX6De3BZV/LaESRZufplQolwOue1xu
fYfXhDJpE/5rxOVl5qv+H9lgOf/RBd3NxWK1zwDbJnmK5Jtg4kY+yjWjJw1ODQqB3qv28cN/xzCf
jT920aiGgy1lhh+Jk3ZW4Wh4anh7YFi2FByrmqoUM2yUvoSlus3WXKTVXeUIEkgMAKnd4gGu6cxA
1UpUiM1kmYqpVZzuFxo4Z7BFiIY/So6PEK9VaCC4sVONlQ9+86YpMZOlN4MpqPfW/1euJcjQUD1r
Zu2V0ixr8WESbG/kLDEpHK5pwv2cubvO25450iB8BtK3OdNZZVmtrLSEN1HfLC7y47RRM1rDQkbp
1L00ZwnBMorKm/zdjYx00OfXQJDUSlHQu6MU/s6Hm5eHlR8M9SUOCbxhaSuDTzwqSVqIzAAbG5dL
ir4vYDhAPe1RWZkca7vR3ABbRWl8GwvAe9hF+Rexed1ZSCQXqQY3oVQPPjqDWnDz86SmeebYN/y+
bRiWTRiHKWEHNg4L93U2k1iNSOlknte0OnUcTRxxohP5D1OVB18qIOSUdF179Kp/+lRtnIb3QRhQ
Pvg/jdyxTgL/lnBb9zehXH6UGrR5icLtE6ET+ohWJhlor+L3SRCZPtag35T5fl7sjOhPLUcutmaR
tCrTMPMeasZYFYsfEYWW4I82nXYEp4RsH9iS3rKxMdmdXHv0d0c/OVnt3BHResGEuH4q0Qv4VuQy
SIvRZEZVp/5SBy4aUvFXr4baCNCG1jYjT1VaMWcpl/0G5S5PG8GeT2vOwXTWzq44pG7k38oBC1QP
OEPblZgaRDDex+foKqLnYdSPY6F9yKc4ogtkqIyaHazTqUZcT7v4aWIa3AGj3ZjB8/N+k1grta8i
kmFB5DyhaOeWmmDqYutGFEHf6gLECH0lCl5G4TLFmxFj4NVs2+OZXm8p/NXd+2Pjy2INtSksC+bd
JelzBj7iJ5sFzl+xmohyQKGGF/Zm2KFA+nV5NjNIgNu5aqGH9ojojcJsSCuV9BFOEVTToDuaG8Sq
1W+uR+uIqMVxir2km/fzEdk1MtnTNdVSO1PMx/SaoH5XGe10BTQddDXyk3FolXdADoQas6IBw2K7
Oq1iYMc4FYFrybrSdNz6AEktHADmmK0PX2UEUCky1fsoz6jVFPH60eM9cqr+ZlX99NwabWyYMlhv
rmu3GrgX3AewUUm/G7iAoKFElOvXqoZNenI+sSu44dnxRTBUGVjyc98kv/6qy90X51D/7PY0ZINU
JUfqMw8HAt9HUKXcvz+1c7Z5/LHHj7XAsOCb3GV6DXjGkKzCaHDgFIxLf8/UQ1f4kVsKZfDxmPWa
E3BS44HkRYt/BSmX7LEv5Ut1cLjoBFcR34O57lDY19bhsiSfSjOKeduSDoMUwNxZjDy4cfKo9yZX
0idRyk/1QPY0T6dRePka4w46sF7b2G2xbDf3JtJzdiDScxAouGrvdAV4/2C9Zhd/AxpVJba8bIYk
8X3QryXZYw5VHOHpKE2CMfMxo1hBVvNgxQUm/NtuJJAr8XlO+yhUwnTxSb/YLFOv+I+PSD9zyXaG
dTyNZVU4RD74hQYwcPGhAbb6bbOQCiohxqyP12KGBMU5md3CWeYl0wxNvt9oKW0EuwuGZLVTjM/B
Wdl0oGqxbavehjwilX2ExldTFJHKa4+e4CZu5DoeGU5qL2onPksiTWXYEJmLGfP9uYgNFaUqGYFH
aLeSP8e1k8f8xLG3imQbInvVOqC3SUy5FliU5Ma5uA5f3EFhSRgQN/GKiQzai7wr8KZpdfsDkVF/
fhhjSC2ZcyM1f0AIN78WbW7RO4kjv2V+rsXbgrWmrnKkm9jEnPcJbE1fNInYzAbqZWdLRPGnA06z
/ZkChraxjlo8eJWYVAOKNgMpHHt1nO9kgX/BIpmUQaciYdSExioiK0XGDGDCQGyP/SkqTw7gJzV3
GLuhYx52CdQpTvJWwN15ASrEKBvxkLcdrWhEV2Jl9xnVpaxpcsyEBYvpdJ34A7vRD8t0U1zrTxI0
EIlh9HO7ku+4u3kqvuSnVvfagATpW28OuqeKvuMj9WCKY6qFY/345jozf6LZiwOQ+hnqFFTSQVRb
qVglSShQh57TqpfoU7oOf/8ZEcVsJ0gMiu2bM1Gip+e+UPu6JHNs/nBS+5pInY2flmbyejwMkCzw
oGRdsytI4Ww9paoOXtkBHsnXR5z/F/qasZWbUs5bEDhbAqEFxug+r/dF1ij5dfEAtiZEuJvJW9xI
MFIc9lCwOZmEctSxi+lSShpWVf+TqJvTiNltRoXy2CEGfPELPMuyInuj0zVvPlabEuvhP0WyvjE3
0nuADUTqbwcUsvHI+bejp+3jBF3Vuu7po7xYQb2CfwFnTotJLoRbZQtPNLOpMMrVTHzCGxGzicAm
CfyEQFJlQ5gk/nTq/NpB0rL9Bt2+QQrfI5HelAUBn/6ecNyFe+Q2Im2DJ2wIiEF4lQFLs7LRBkrX
F4PWyVo27zTzvt+BDk/kJZFUL7S1oSaOIrZHOa92zoHGs+MpGVgYpYbe6z5gRL50+uynEHI1Ys3I
nxGJo5oyYuVfNVEJFkRp1ijGDcwspgy5uc/Inv1u5R3u04n46EQzXImMm6dEqjesFoZ2gOCa8vWB
yPmsLmuEEbzJbHW6bOTxFQkvKqbDsmfbbF2tRY0nUz4KTtz2B6RLMH04icIc6EdasbmVfUOp95lp
vT+BcEeo2VBXYWrIB6pd07ebFtWyk0qqcyXVq9MY9+Ow0l4cry3n1cCNtFdhSx/7EyUjtlUVs1aM
GM1TgvlfU9P9O+/2TZ3snlRY0AJuyhHgZLQdQfnoMABgU8KhjIBqUr1IgnrNluYTFnyv2kUh0jyL
/G9G4B4mrgXhdl90KK+VYYPcx4PI6z5VxPfwygEp+E2iX3SkswtWK9MV4kupVnmQZ7hc4xprYcqp
0YPjZRVRpLkFits30+XA6Dl2U6m5tGai7QTUt2T4eNyZQVRYrOSS5LNQW/WcpSPEyMpB4+CpdQtp
7vHcdtBJpmR/iX9Q4Tz+mgZ5F3upWuuqorMeddMeMBhp4AyFOaRBt0N3OI8TrFvlTc+viCjpS2/3
eh0HeDd4g1Vu4h5Jmv3sL5RavEisvnnyOWNW0aVqJCQJkqB4JllEo5Zio3r8GEBdGZmAEGNrw+94
3P1cxPwCVxH2KJkN3F6l3v/nYxKdBayy12fi62TYCkUhS3zt9BVun2rei9w08UMjxeGgtGtNA8m4
dFa/3nhL5uu9Pbm+BTfdbCszPZOyes5QbWgI6mRcdV5BCAEU90c1hBwbyEglyiK/2lso0Jjkq9m1
esd6vi+PxIkVSK836fqjEZDOoB6YUlclfzUQd1Sf8jKkzV5DeJF1+9kZCD6y7+JYXOPwhyx4jvtz
MVGl8JrSsx5Zbp5+/CAu8WZtv7muosPXhuJhAqNsaRp6/Nn8QWPzQVSFNW20KUxxLglq54trM8gz
kqFCtKTycZqa3tf9VanPdOQ5Oxii85YqhGfwG11a+NJQ368rQ5MIU8jvybxNDZfsyuNK7MXCflHg
vF64/oQ+uDzulaWJ1KNrWOr1h89EkTXwNg6hHcgirgA8pR8bwY9+ztTbVSvMRF6Iyw4FRQF0076d
/R4LQ7awxMFQSfqp5uz22LsThNluj4jCxAvS0jdL+VBAqwb2BnciYleASRsCpFLvRN604a7FFgNC
A3i1F0I6xHT3v2dmTrATgMHcS6eKhTUd/bUiJ/6MWummxOeG0w7Vf/k6+bqzxTOB7w3mhI4XFA29
VvyqoG4eCotEqDnqYMvrqLblcn1n1F7deedNmAxdKh68G3s/CxVWLO4l+RafuO1fc3nMQABoCR4D
Xb096LdjiprBVZLL3WIixRxoLrs//ZbMAEhBvCKM2xVJMsgNsN9juCng6mWltnF+MeBW4vSXV2Ay
rQXWStAZ5p0808RBh1u6vRl2qgreFAtPI9C57DTX8xDcc8bdRdMkjop4avNUvrSW45p51NSrkTXB
tkt8cSHIlw5y4IJjZJq/OIihDlUWTEdVyqJ+YBLH9d9RHWhaLixg1emPNk4eb/hmH98OJ9Caez9X
0iSG0q6oY4HA2CxMHrvm0MiqtFmpjw+Ja+paxcEEJml93gZqlUtaWwy2lzMMANsnEju+T95WZRw1
4aNB9VIbLLbLgFJYiimECTA3l6i8R2PnCvkXPHscnQt02Ah8OZSi/XQwTNScgupsS0iZxTcLsJmc
cqDZt4pndDgWOaQl35Q1uU5HjFwdNRa6dF2rGwFrW0oEp9mWLywfQ7/FigVGTTo6A8perUSVL5u4
0+yaHySNv0/3rMXo3l7GSN6tfKX6TlRDNl1XRbTniFl53Us77OHxavYK25loZbd3sBVebaKGv57a
0M21UiuwthlZrBUqVC0n/4CsNVwI1XD0hXR8/uA8HwOTsLOLktu3vIF7zmNwJWAtkg6/mhcpKS99
tMJ3BqZYQlcH6PBFsxKPZ0MZtFMlGN8jmqqVBlL4nh7yYFr+wntRYP9CKGZT+J8tW0VBn6c8Dh5K
j64Rj0ckaCgT0rL6xv/9L7mP1AKHPzssHlRAIf3rPfnnSHd0yu+xE7sT0gyDiE0JIrEqIt0mdHeO
ws+CXmBIeYtNoYgKFRFsxhWkCNKTiWbHvuxMf6eumw0mS6U2XeiVOspEUbWz58Lei2U40dzLppIC
8U7B6pMNA/KZ9xxh2X6bL7R4PsPytOkS03QaTDAg18BlM8f94QA6cbCaugM0eIxaSHd382lLPJ3L
CaH6KYNpC05mntfRjtMSuP5nSQ2iUR9LyZUVVQ3/jw32mr9NVcAVPWHIL0lYOVRUP4LYMo7Lvay1
2EsmD/ezBsqJgezwlVT6y5tw9fXWiZ+J0g+RX7mLeJXJ5AwVK+vCW2O2awY4UWYUrv7K4pbkKz5B
G170qOXiSSxD7JzqeTEzcnEAuFu6elr0+7NYfHnmwjby9H7xhfvWnAtRV5NWAH+K1ZxbLxi4ciPP
jD6JlNk4cdPYrXvxOjZRqV1yE/APAjOSSbCITAxNtvPmTgTv61JfaU2UUrNGisxzpEFxE/hKi7CW
9+2sQ8PAKLg9sKwVQWlTMLAOh+p0zyLjwG34j5UezKigigLSSuzHGg75d0V7SuI2OZOs8PumOqBr
CUjoTeIf553+eEJ6RzzcvQqGEzHEVwzWRRG4rUFX/5w1AYRkyjNrswau71vFE/UHoU4RyyShSJhQ
ALoQC8OpfHIzH+E/NzNNThqG0BHWgl5sIJspY3ZnuZh+yMQ/w8CT/xUeznVY3yDH5WYRMLK3Hzpo
qylaMyby2hrwAvoM2XtEoLYxdYWCEaeIgZFtOZBRa/fV8Ofw3Yfy3Bf3VHrahFA+Q4E9vnMEt6eK
z6QOb/0CWDd9317Fb29I/Jpy/aI57k9QQw81LD/OQMbdKXblfQVAPXHcptDGr7Q0aUz/NTrdfadU
o/QMAIQyxVlnlAeI9r1pASTcTY7B042Hzn2lxseAzDjSBrwm0iihlizLrMmvg8y4K6rgtEORbEmK
zubStIaVvmmW90RlXoYUHsFp+e9MwKOTEx7xcfsW6MVENM0IEW1InsEKuIFWKuOqVWHkxtOE7yBX
e9Xk6EtyznfMBA03DyGeANSffncgNAXKSGI+7sstR+pAq2ewtgTk1PoqqlD4g/g0s/NdCZ+6/XXf
MLQMRbQLXByLx1kEe9e88ez2MEcuCupos0Fbk5RGI47Cs+d+sjGsAv7yDslX1B0EhEMlu3RsJt9L
YQDckqxwEGYrltinAiJyYp9I4/sGbx14OFJgncdvt6Lcg9TxlREBcJL7TJXzqQNcjSLJvYeGBAhK
tpyzdm0KgUKZSbXuqEm0X5DL+HLAcgz5UtY0dKcdnhYkx3kQkhxm3cQPnJ25WY/R/f3fln3Il95W
s7Jb+H3OlJfFw2Q0FuQW7XB9kKZkHMnvtw5hkd/SOq1Go+LunLGXsS9uwKsqC4kH3RgUuSYuINzX
QkTvV7GogPwpPL1XkASPbPbu3C6PuvlCzWJ2em096gx7QGCIzKnnxmR+h6dQupibJ/VV+q7O/mNm
XVVAZEl7IVA2s5tdvZmhvFGM8fCVkxLeL38FnPwtMqZyLD5KaywXkjSTL+E5slYWfH4R9H5GyRxT
CvUQ0311XvNvdgV9sDkdHlANXUyEwcZQBbPDxgzomIbggCZR5kGcTE9vF5Acf0NA2KU7vZvT4amq
WoXu4KKMq+YIZ5F3L9SWbr78rb0KtJsa/TEZDx+bQQSztfagoa+znzt0aBtA7KznnZTSy8TmJjWs
ac2PFG65ZVSJLuu+eYHIdURL/Va23CdRN1fss6DRb8lLCk47ZVIsjlBLAAqBH3g0jR8xTq7M3p5G
RoSXVj0yxvJD4R2KCjTOZpeA5434Zi6yK+iwjUIR++5Na/yYLJ8hx6FDN9O/0vOQcp8t8VvxrpFb
X661yCR6tzbPNUeDfeU0nvDRpLXeYUM9KtqVIpiaNtX7J0nhobOblG5j2tUNr0ceptTpD2/3bQh4
XgCpgCZjVvoVkYcA67LoZSOvue9W7hNpsycK6muPTERW6ihEBNcf+dWM7uBHRwG2Vu1p/aCjHRgO
8/2+Zs3m/8Vqvkf8FF0WV032fQvGVblYVEttmax7UZapbt3HoL+qNuoQM+oMUJ73lZAU+AVJfs88
CqyQ2NGtn+KGq6ScZ4Qbc7eVo6WW5cKzHFGbrR1qitarS6Jw9cWUSagTo+a7C5B4Bxkjk+0dv1mC
YxvzFb6Lodh5vwLMhVO/VKcIBLux+xuEH//GVyx08gthCddKdy0gyxdJeIa15MlwR6RlGOePn1IE
W95zKZZcy0LHsABCf/5f+Q17ahtJXxgV/oGjNEuQExzsyB9XxNg0zwyzSpTBsmjxGzpWDbarGjxs
9Qku2FfeQqVRAoI3Hcirx2Vq5d+w/dHdUH3BbqkY/DI6ilpwx3nqTzNno/PS3H5ZJT0n8/W1vOdE
FTnxyeLjkbBzHnJF4w8QUqQnDzWso0ZXhK+AUaS9QWzYdIIOVHOEkweLfmHA2F+yFcGzYhQJi0M5
H5yOYKWe+NxXQhHppdHiSYb1JQGjwdiUHgmFillOlbEuEwoC/kFm3hTp7p0qRb5QuNdZ5QrF4Nzr
YPhDf5+KCyGamwkAUUsDFi4kXNhONNZTpy1goKWgqScLqGh+Qn8j60X0BQ37AosiXY6GNlOgztrw
Nr6IzBOh7serOEWijOyU36gcL5KKfUsL3GTl41dhqXVzRRF8ytTGYVhNiFhP0TwGhS/VBlXAaH4f
ycA1bvFN79bCLvq3ifUYALaq9AfAVBwmH2fm1IpFtGRBrBYKNt2AMv+lPSN2W0cl0GhWbIqdWmf7
JCbjpzlEc1sliCOSugvJgljCjnJx9Utv0qXnrJGagaHy8ce/W3mv4V8xBpT3Qc2jrDqv599yVGJ0
R2t5cTUYzFEOD++AAXQEmRfzcKi+0JMa+WH984yCzNPOo9kgZuxq8vyjRqeTWAOLS67If8bYihd7
Pkzm+hxLhefoHbGggddJYDDQZ0ehZZc4CXrhemByLBu41iUof0NdkhRSNmLF2XJoWTg3e2SuMEbq
qHeUk97/lratU3WSyQ4B7WEBDMqrqY0eK78NLoLWq0GzK5zaEI+PORRUJ6lgUv/0TPpjdELNyvir
SBi5FTvps+GxAGDg23xyB5GtB1L/+kLNkc/D1dF2ah0XPrVv/TO1RzCaAY+srIr3i8dj1sow1M0C
n6M1p691o2zbGl33T+DOkey+PNsmUVSXf+/axyQzuYC1TeHB+ns7vJAGMHrYl566r4T+KcN9mpyt
I0N1vqWqUr+YR9RfISKsa3HUl+LCgh56AGiGGxKVWAjzi8XssRoD9Wf6irxSuaUBj3b94Q/Afsbl
FXiXlRI9Qjjjqkd46Su3Lour6Krn5mq8sNSIxMbobIRXgDWhJdc8yxjpeM0KE5vk51mCHajSK3kJ
x4mnlrKSoflT64ir8BfAc5dosYsrRIOq2/hB1S01fK1IwuWaJZ1BVorKeSyCtztgp2NSoGJ+2IOc
kH4ujOJ1Yyx5TkdSFaoTW8+hnAnXpAQfNI0V5dfsd+ci0owR8JigpYX413i5GiCrhu88llHuCKcM
HDb2EbhTIZmJnMBsw+EGNimGDI7QPLd2VIudGrgvL7JHPAL56MFH/ST7vR/a6uZVlY2MR66UrI3t
CYnMVjuRJ6x6zTdnryj82EdAk9pYV/Vg8pjKt9TdPrk31eivv6vuXxf7R146k5SPUsiWBJInSzwK
Xpfh/pmUKYxau4r/RGvfx4SqRq4ant0JomDKZXIeFyHHiP8wuiuU8BZwrz3kcQXkZdo7OUIhcui0
Pf1be5mbAt4Em1IiA8GRxZnZ3MM27Egf64TZv88/a+izK0Kjx5PBJXhbybDoLQqsBaRgVTd7lD7a
HZI6JdbrDOQLw1oLK/JZW4S5k7xuHmZqPqv9n22LfAbASz5z/CWKsChM2Um2cj7WHtkxUazz5EjE
TGb8tjy7RsBa7FEG3BB1Au3tXyJnLBfw6fTuN0xeN/OBAW64hh197rbSWEEp/YPURpEg8Rbb2nxz
HVeV5cQ7/71o7k2DxvePRzu220xhtIZGi+xtpPqGbZGv1SdVMprDbsXIuB/jANkMLJRR2e4E6Pef
bYlD8WlHNNvW2eQrCb7VtNoRkd59+GrgNHyk69FqG53Fr81ocZ5TAYBbGDu+y/jcY579NanfIEVE
+IFpgGODgfW8pKPhP6UfdJf1INjDXp0BClu3DYbafX/aRIN17xhYe2TYJ9lFoCFIP9iRc4vdmWWl
Lbkh1cNWycKxp6cmCtwgavUS+VigJtukzYGCNwsgTrDCqqrcwlTP9kky/yDyFbFpC0OwecLNXnzi
PNrJrxMKZj260syLmvaY8fpcaIvuIiW+Qtpfhs5Pp9TUc+GIx1caYmFzt2uBOTgWd7pxBNjUF6uz
ndwE0j2tHOrrUoVDT9cfxa60hGdqnDqUsBw2s2iCSim1ezQ6d0PmphHxM5FRzyhHxwMCFTFG1DnH
Ex5I2dGg9qp3/sO9qdMVys4gSFvkHy59WpAnFfTfW7hojdkZKeXR1Zd8N94IFDMxwcNdXG25jswa
9m9JiBA8d6zsvHuCIX0EcEAzy6MGly4SjRMUK59bGNotOPW8sYxEUk2DcdJsvmIXjpmrXFnIqUZ/
VT58ZTYS+2QVDRD6zxW4fnXBeBC/CUsSUUYpPLOfYvA7fYwsouu53fpgi/X6Ah+F2bVFcMBml5UW
x1fQ22q2asuQPpklRVygPq4YzS1jJTPfJb2UBlqOwM4gGSrtOALbN0kbR2lIdNtmtbkHh29Lb1VC
tY1gOMMROo6WthVh73Zb54c/xNPgLF4y4pUJ00pOVXgNV+xkc79UXLgdekC1ObunHA0WfKbeV8BS
kKpkMulz5ysLZOsF4K/GpyW5Yo0vXnOeD7S5bgcd5JWHg19q9GJXNr0e3CW06OP8rYApRlfp4NZH
FEzEWrhUnft+3McJdRsq+vYJk1PJepSbf9pDxeAQmXQbbztB9Iolj2F7k+95evPMYYVKIRAEFKGo
iNq0yyfGIfy2bAwcUhG+WXMXITOwKbNeUVpXOvG+GdCYIooSJnNDegmcGRZ7N0CN90IHpEYsYBHA
Gahn3bmBQSbGHv5pEdH9OZfEckn5c+HL+KNk9VZGVpz1FcF6YL8CxIXR5uuZ0X/c7aOZ4lKQqcBf
2eXzs1JwfIAWQ5bxJfUPgj8QKH1tVuJviiXYgl5xiNXqH3efdKX5APaJ01fXqBGPzyzBRhhC78VP
sdwZTFuQjtzs2MWbnA63Tu6IxIuLqB/9WKJEBVxGv9Gu0zVUYwU0eC6LZxsIx8g8SGnEvXBsmN21
8MIu+LBMBwb6TOuu9nAbtcXmuYkq6pbbG4cwW975glPLOGnCNtR3hpETFq5vlgyef4UqUDJ3X63u
SMf92rTUZoD+DWRVg+NBsnPLWv2esfunnz3IiG3WavCK7wFGnM1pxd/wqCxuncJSz0jRwFuMcc7r
irl7bKhNGbSugoXZa/uWoxhjfG9bHnnDtTKPAw92A4jw4KjIeiMq2cTUe9Bxh9jQfIMzPy2vJBXl
cvA8rKS5m1NpVWsFc7cWt3xaW2BryBFPmOr2wJedsSB+Hd12fMTIHqZzeGdZ/E8i6LPTXqRwqnKs
I3pdPZwUHZ9O9G4YNAIjrXvS8bmCO3Gu5GqOBwRheVdjn5b/AcO8QRoJI2hTk5klhTId/X/9xaj/
5tIvefqGlK3+hJMCF17mL2BzFaglnnxBdacXnJheyw4R7dAOl9nFgk9mTq79sgRnfAKi4uljOsFt
oZzY7Y7CndzkHCQFIJPZ8pva8PIlUMwxUW2TuCbvN8WKoE6kTr8lFiYbAULSFk4sRzLET7q2Vnci
aOvbj62a4+N0qkkKP60Oruw9r4gYYhK5sew65pXGF5yBZ5KXlK9bi7RdP/IgUmB+O90WvcEcH7wt
Y7kQj1eVE1MgErMiO+vffkGzFqoM3QkIQAu3OH2UVkehCWKvelLUog/Ng7MbTQghqqWiKyxvLbLP
FkIN5qSBtrl65Xw7C5Ta8mXZo0FH1h99gaMI4UbEXi/vVzzxz8t3uA/wQjF80N2wLmv77bgR+MSy
LHJuU0SRcntJvpUVZ8+R+Lq7VQWT/tvK3Z9RWlMRC4+KbLHvu2umS+23h65eCcoYBFSo85GtaD4G
HBVJr41MnJtgpfn9lI7+n18140iGuLR9uPZd6NWP1V8wesCQF6gazzI6xs/bxBacZ6MND2ySqqCF
/mieo8LxVlsAEmbpt8OuWXissS85mcnYJpTIH/8kXhnhykLoC/YjnMSTlfkRgFEA+dxkZmMkMru7
pU2GdheUZkU/BdD1dZD8QkS4yvJyMG3sk7OWvQfbgkuKI6JdFBkGi24JytAsq2mLCTvE4bM4WyOY
dJ7OBcCdhEv0bjhJoOsm+yTnLmBJFRUvsso8kX99QnGqiSdqr6g8ZdMLFXJIFEXJ4+TNnT9fnioa
4Xwt4/4c6ypDv3ViddBNCyZ92RWFTKIwZ+yQBz1rrGreTNfM9hXMAuG6tNPo51KeF5CBiAxlizP5
b/rF5cQ3J3m1seOy24VrI0pRzXYuwglqtz9RLmCBGgohw8mLsAkavcheLqrutdAHPGLxlFU6axQT
pEHOewBqzGCB8/pUOdp9dXx3ZoZGl30ICms7L/GFXJltJ+mZnIZUfugMPzznQdl7NTtYVMxnL+AL
xJZxATsx26Ehwh3FIqtFe0Kccb1oIpJYnhsa8A1MA4e5UbBxgT6/GCuBYjpXqk0SQqLiLiKQ6zu8
pP2rn9OKPKKELyIKQu3vInecZAB/UT6RDdsYrI0Ttjlp/xFBqbBZUkv/PuurDIDlRveadj1wAOyU
yzr5ZyYYX4t4iyhL+zYBPevBnL6nMN3BPjoPgfk4TbSDBJCnCeXm+6PvRCurwHqniVqjcg/Cg5oD
Ut3URdY3lqLBzWMFK5lv0dBMtnZUGO+dIR69b+xFYSZGvGYkQq/sDK8/T+/6ZOIlFQkxcHbGyGU6
TKuc1ABABMDQ6H36kZYpPZ4q5a6+KB/mqxB6/J/SWw2DV0yA7mZorLOKLMKVGq7NRIvdNLCTeslO
5NMqPbezFSLQXQvBAGHhgsiM2Vlt5le1tDMeaeZ7KMkus48kCP0t+sKwZLyFa+Qp5JG9hbbHgYny
+Iwi1sfhwsI2E/4teBIblq+m0Tmg2tdaeEmC9rFFd7lFYIzGITWvTkm0XOLuafVOo2hotwoUtA7H
EDYP8c+fzvTjvsazuA/XrcEhOnNMhLwLPhwwca599oAoUV7MyK3na1/eafiwKrRSmI9ORdUKhXug
QA2SY9owOGApRin2MH2IvM8Aim8oY3vupLvFwAoR3r1MhhpVrjMCskh/EURNLjuU1V4Wffhvl1dX
9juxxExEWtl6dcNkN3r/0KDSE15zwyaUe14Y5pf9cjkpjf+uQgzEv/w4nwNFvTRNxN83yJZfrxRE
dh24p9bkYFYNia3j/pLOXqycgJOHInQSs1/x+m2LdQV4YI3ZgD/ul+QWlAycRNO/cw2HQuOYWzBX
UTUGaDj8AklKQ+FucV1lo3/pTg7uaxJ4+YbnKa1cCchkxQwVMZXDBKxluF8Gnqs8Spr0yo9LH9Os
SjOiNwxQMt1SwUizGrdcMCLg/NhRecGymKSKYkb1DJJVmwwwUZnerW37R5jI2QG9eQvf3LnQkzZt
h52lwmZJuF56einseg0akLSNzrSk2WAy1Fuklf+c1rXXYH+V82ZSsWNh98Z5MryaNeTezlkH1OFu
9wluW7YxjEhbYtbWkXspKJvcPVImHIgSpQB5ux6z1jqcIUGewwqdkUdCMMVCbeNzvPsTDPaCw1A+
u2YLkcFb76hDIfPtcC4EQz8eMWdOjahvw91gQKUV6lhpddi3mLbStBT6JWEXb6TjEgaOhSHTn9CL
MzSE+72Dp7CHRdzNxJitim4du7Zm9SS0KqQ2KcCULVFfa1if9tqEPDlt9hQxOYAvY3UJ38+Hwbge
CbHSGrk3iraLOBloZlYKCqZkKJLs9M4cfdrq+9jqZ6gLbFiBDaD1QQYbD8VMejRcf98ZdnS4xVHm
sREbpZlSH4FDfNk4+FXGfx8n/t72apIIUdyk2n4lVt9tu5HPxwzoOsmoTl6RKizD4BjShTwRSPGn
+SozVDY/bBcKaz8SmLAQYetCPm4xC89+IS/SQPktpW46tdgDRKOHrKCDrS4L+3At2sy6qYzRaHdc
F4IUrg7svnydNKLn6neM2u9weYdMQn6zumdJvXxjbVpUNzMmNEFeqQGp62QX+zDc409xQhTXu5KY
lh4UgyDx0k02MTAM/TBKOzBlojQAhTwvqhRjNj89e5c6pxVQ3c5QWPjhr4s4BtldsPdakpxGcUS/
54BuKTuKpEvhdQeIhx3cUUzGwWXU5BvAvmFtLiT7xsFcDF/lJCR9b3/6hYKY3EltzKmeyQaDdEzd
Qzv7YTeQiyJxf5WCzd+JmM6Op6cNS8q2yISvKgNKqQMQozLdCl7hh+RkLKFDLlduec94pkFlUHKu
kHkseivhlnXgCLvi0+O4TUu7iiX9wx7pVCiBiUGXMqd/uK+VCxugzYFSwsReBZzQhQyGBVSi6ol0
990yD2mFhPreVxlb2Cr9sEvyatV4ccIOYmlWEz8EXxg+yqi7bun8QTkPuY2SgFkisSRQwVcyumdp
pWBJCqiSviFRUr2BuA5bJQl+B5XU8HjxVg3y1cpgJBcd1r+f7WJbmfvstbMxdlYYc8k9+TQ9UksR
jxaDHonTuwDMODLOlWCxpYliQnear2W69kAXTG/SUQq3wxJqmvcbwW51U8TxnubKBPH0mOeDdVhI
7I9z5K09jMlp6+m095w/d8hfYp9ecU1wm01E63Ebzrnkrhpv1ojajyHuXkhpmHDdo+o/bSTdBAze
AjBDu8oFvnC1zKfHpLoL+23++1lz6u6XQUuwA2b2zIDZnEcW+QJQcTL4+2L2me/iV9n2DDO56dC3
FU7AXx4gFotXYzgC/LL7NuplYSzOlNctaKL2DnLzpmGQXOJZp+fejloUJX7bnSkHfz44m1wzW+Ak
WidcKkudjTYe2c8ir3xYPFRDZI7uW+9e+o020uqgrn7xx+t4FJg2gctlHyPaITeeECLG/sc9kImT
JB04g2RBoENY62guk2wLqtzUWtKVZr1+PoVXYnkXC9s2th3qVdpPiNCcRXGubbGPmRwKctANI+No
Mdpc1ozWhafCCEeU3f1RcBL1ahlAjQjNtWaMVsAKe4t7p5wnqDIW0HwtnYBT08iyCeAezbtj611n
BfXbWxvy2C/zSlC8Fm29rX6ZHdVfODihy5uI7nIkFpq+CbjmIjPQLAtQca7slSLvUHFcUaw6XmWL
CHXuALSxpMDY94pf/pGF4ruzOgCFCEVGxBVJ1QjR9seKHc3P/nxpek8FllyRccQzPDBfvw9LSk0a
H3qDE1xuNJplbNF3hMesjDa/+cH0qeLaOpwKNRncC3PTaOynJkRJfwWRjjegls7nIx0LMoaFw8EY
iiwVHhPPA2h8+WazwAoUe4naoLSeGGc5L2uNx/S456hv7eCt89p7X3qjZmam9engnM+8XVpNvX8r
cWj+BElRjgVya7piBwsmgudloJ9mMnGJkeqMyokoFkHzBt0pHvSai+PjDSADO4TMriRNBsAXdySF
AR7rbFixtg7SlZk5ojvml+37DGO7r8+LKMg2UshjKWuVMfCuTEYMkQMe+ZPfQ4VZNGSPve3Je3iF
wJmFvTUf3r7OcwVFpsK/cq+g8Y5fA7bHnPQi8j5kla8T1b0pEG6FaeELc+2BOuXat+tevALivlIP
7bjz71bloNBRQxxjGtZH4hgANDeIDDB4+FyGbm0Jdzk3M9rAnlSzvKyoyhyBdAoi07kUtcXHz7zO
QkTFIX8ED+psMC9PId2hgrSVTu5TlhqleW1sXgPdUdt1Rn6fPnxTWqgadx8jR3+uaQHNqwS7SKkw
Llt+RVykIRwNjFAZgH0mULAe0LNikNpNd//JDRKqr9n4Sr+Hd85lgFg1iIJzyueI8Vrd/Mg/IRhX
f6IsFjrThaFU03P0w96Xh525cdAG7qFvecAAtTxLIHNOImKvo9Bz9BQu81y7SQw0UBwSVGkM1A1v
xx4vFEbjcF9XzXakSQET8PBXkHIzLdyd0bekq4KoEaW8EUQl+pbVmmLDDJdKznVKmBaSqWS2T4qb
+AW6w4pWiiJnpeZuVAny0K9lnLK+gUfUSGDfgcCYsW8QTxSCbIbV2IEY5dC388QQf1i/7QJnnssQ
zaSAfVDwYD6PxsyVRCXHYBTEilrovdzftARZ3osMSxcp9rIUK6kTJgFXgPtXfVul3SRI8GwkahBg
0WPMDApb7X9AziytW/V1YAEnVYGyIf/ChkiNhUqjokekMTSM4h2wsyhr2U0fVKAHNtXVunOWmutk
tvohW9Nu5NecrKoDAMeihG2bnnhOTO/JZ9PkJgGt2Cgil40wJ3Lyh8iOCiQrrZjF98zcCJFyZddS
DIL69VLZ99nI4LSTskIOy7aNmLytBz9layWJJBcsrQVaiGoR5NCXc8I8oTGcG4/BxwpvK/SCO9NM
qnIyetkt5P2iMv0sIe1YrDzPtxpPzjOsNyLtpEB1Cxq3/sUz7S1D6wIPHaBXXVTNOdlJVosiP7dc
CySZKhhEwZTmU04oUoJje880QGG7+9dhSF68W52d5NSsQHUPNxviL7Q69eLsyjRh+H3FB+P2gjc7
VK/Fka6YA9KyzfdO5VSezsYBYrbTy4/BpsmBb4amCmOoWjQyClpH/dCXLgx6OzbW1yH9lvDemolN
rH7YQBXf1zVdQQ/UiencSMAWh/o9FDNjZm3aRknmtEffdkUopQPe2rGL7P07kfOnqKc8JnBWmQxx
uXw0O9pH6ffcH7xp79xc7Y3rDGrrFMjd85VMRpU0ZDaArDKJqTL9OUe01y1ISxyWXLszs07dmVFz
A8EGTYJzoi4DocaWbOx4rCgABJjl4NRvYedexg1QfuXDkY7rASm+KTx0RMeLDIhTuzM2iZU/IOH/
FDqpOeqflFBjsL41SfnYIwbvvp7SipRTWC+Le38JWU48oeh7F7nifZAQxrISUzE/S7bAmZV6xHrX
y6KrfpjJMFS4/m9ofc/cS/r2wprzjjfZavlF3AOoVqVd3muV7x5n21vo3k0sEnmHCwzHqLQvx3DB
t1Fwh1Fh+u1a9KTyH27iiIKztPJzIEo36x2C97jvgXidH2ktgMYOT63qFl0oHFw/PjJYh3hBWWIs
cFeAjhQK8JaEcVnCOMu4vuLloobc3RiOAdlJfU7reInyHqxZLdbySuez9xA79qmIRoH8TkyB7QWp
Y4qPTA8q/meAhfEPWYtj1ybhntoakeB3EQ/FNzcYoGQPjco/7RcRv3QmRb6rPzBhx8PDa7a4e6DG
yCD2rhROBon9VjkWeTEz4dE2FaOgiVgqnv0xocM7XmDlwqKffSrWR+1FFea1hPHt3v0W3JbUyHfO
A52c1e8xw64JGFtN/bPdbwcslj8ntIDB6SlE91PHdZARUT+HoxnwDNVjPh9TMhZQic1KGHvvhm0Q
ptx+2yPwBS928IAKkXqJrFyxb6rAJusKevvGgGnkBic7PnZyON3gm448Up7wsgfsFqYnXoF4Dghc
aCUDliZBjoYQa8M05y954BTjr9YZVtd6qZiSJUy0PQALFEOXZSSaNdWI+l8/Io3kHYO5fauIOhKP
zXYXqmcHjgbA7NwCnoieZPNwcYeYUzttGAtkSSwa3kZwWX9hB51KXDAwrQFYuGYzXVZ/ZYv2tW/q
wUUK5LyYGnvCl5u8cmEtTZj3PLkxCzEGZfJqfKbaVpao1cb+r9LbejqbhvNPgZYdlOr0wG51ozpK
7vVytoR95tnLYCEHn2gqDFO76uqFstxpOYeKzm1bg1jNCBDF7VDqSG0X1XfF21gMHl2KLWrEUijs
jR0JPeb+VTKNrIYGNB2xamaYxhmJtTjN501JTpzLzzLYwNO6d7cFU5nDj48FgX8l0BWx91CIio49
aVTK+qR2OHjMksE9kWSomDfjzAdTu79rTn76oZPGYfPG0J6hArIyjqq+GroptEFawVDq+IbJCgTg
Vm7rbGSrPUpsb1nWjTzxNrkf1BTLxWSgGUFZh+GpeX0nvyntBRxEWUvlk9u2a9ED6+naCcdhC66G
ycRpeJUJxrmjsgwvdT7MH6igKu2og8JLLuqsfP1awjufNwL9/zXrtzPu3GvjdZ9UyZNIB+Q3p8qD
fWqMHeHMwnOgIakX1CPQT9aybGstNOYds2zObmASYtHN6Z5QBtIxebHd5Pxey9wzRu0mugNtb36e
M/rY9Weeqso0S5eofNPPjyjrzV7Ces87bFf9kqMrAJzr+EQTW+iGgkRl9CMWiYw27mYGEU+DYyj0
EX7gAWQmWyeINpLyaiO07hnF4X07IMQXO1/uN2OgGycO9Sj/rD9E2RwslMMx0PUbrTuHKlq3lnHA
22fZrc+KjMyDlVjfNIcLS9nMAMX8TClKT1fpGAhPCb/3NN8Cik76JNSkBeYzbSjLBrameWHOSDeI
JZEPvAp08VuQkg+lmubxFO8/nhgnQBYsaO+3Kijp+Q5CMXwUjx+H4uezpQ4X7qYHx7e78jUFDYR+
LaWo3Iv4vlx5tqg0WbyC03hhQ9K4Whz4mn8oxQvRSCMeRsURXeVAxpMBAUIIBVnWN2fNREVg0fHq
qG/30g5DyhqqMkGfkZmP1XBLFEdw/EJr8yTkDDTSQh4ohr2SoTriqYpxgkmb66BsNgCrz97KhQjY
rYaxHqZ6vuyCIE7M8a5lpgAqvahpJKVHa47rrbAwGoKf3UjBdGt0qDbSJuRsZ0Rv86hYvq+ICS5g
PhFIrBbr4z9+eF+agE/Q6xSD6So2XfJioztUlZOEs7NvPYKadkOjhkmCHu2mo5z1NSQWlgG/iKEv
yaw0kBMoVdz+kMstg6Uuo0jgJA5NE7AMmhbSQO0/Q3pm2P1mihWvzttARgNjr9FSA5uTMpAkCYYt
O3/9RlBDlbdBJtwo7jjak8q3USHZQmPFr1jGcXsDvdea/pFI2h8jR3JSU2fP6kPNxRJucNB2UAW0
sjYUmHkgtt1jUd5ZzINB+Mdy/vu/jY/JE+0x65669B0B8lkcPT0VLVSD+n1dpRJQp2oP5T1mAF4n
FsmAariw4KAdmCYZcDZ8c5xtGnICnTIlCt/ZKo/kF/19kbbqAgx9xl9OAiDF0flYOrAyuorxl6fL
d9uJizrbpnc2Wv7kCwZqaZL5EOhIsUvmUlkDxXSUkeuZ4BzaP4ghQB3lVm0Oo2UziVEM1AnxjASD
Sm7hqwEiaqd3VNhke7UonuZS+NclX/4q2A3wXttDtw5yEAckPaQmPt1SKGtTtlCU4Oiw1bn0fUE1
JIQ/scAZP2jw5qsY3yEGO7w73IqKYJle7njQv/Z1tKojwfawSh1H+pnnKVKKIbL4BkSZzbSSVp9M
Nj/ZeMzsAMJQiDiTu7cSkdq6Le4Yh0w7U5vBY+SZE6uWFrRnRozrSkmp2b9tkiWxjFENE2MXVRQD
krEUr2yYk36SwIxxriihEwMdnsBsSwc3Qc42j2E/i6e1xtKw5O7+X5CVyWkCj+HrVPBAiV93CowY
qIDrr5ey0u8GNWicprnFdj1fazZ8/K2Tuu/KUixkfW1JmSGFkiQnWaG8wPc6vwvyWPiE11rGuE4V
/F4J1UXIPCflYL9sDXzK8kLfFkBBZoy1NyhyN6i9LkT5Gq6z2QW7b330wTwRv4uhuVBvlfdoprpS
WkpVbGs0zX3ceTfasmph8Y/CPyE0XzRCMvqHznw6yIjlyHm0RS9ne8uEHQKh9Iv6wGe9/hznxscn
vGPepMNz/zlgjJdHRB6sjqMi2ozv2OIzeQqRDXNnLAWKX6ZQF1x0td2PGR585R24kKDPI6Hakh/q
bkSB5V435v7cW5rkEQTUK3X5rDewTRRLZ9J8jO7ny2Xgwx0nzei6r8bJmxYQyr8RxVouMQpeV7Ei
JvX0kozFL1OJUld/xIgQbr6Uyhlv+KC5JX471KDxCJW0/1cFqK7V1j2TWItDo5Qet4usoD6/EBmx
uZbXxfdN5jvus9A+b4EJJOa5OyJPxvIjhSaOno8ZuVmOfdwkZXXDJvC7dqPWxa9nnVUG7AYd3i4K
MnUm+yXwJn+OIRhf4o4eqgvLQE87t743EJ7xHiRqsezv0XTOZte2fkWzZB/Q3NalNHWmtpY+7fbq
XOXdiOtdr+KhOFPJuT5T0uaaskQ6XkbdtaC6of1NwYL/Sl50BJK4XkQoMhlXyajor+LNCPxpHJWK
FNC/16s7HQPG4sVMfG1cFph+MO6IsPjAlBZ0PaBzUViiaBAXT0eUP0nLjEzFAQyTrW4opMI2ru/n
4o3XpVL4bf5EmagpS7Ynuv383wkJbL7AzinRLgWAnPcKKpEym6D41/hxd/9U4vs6k/pcH8KolwEg
SdgrxwMR2aw7uDUwtioPYxpaBL2edbJn10kABnpbX9pMWvjARLEnV+gowXNgfnrQ70AV7lLeHGo8
zIsTaW9doD+MLiQCWEsGDJ8GIK4/8UYWGJ/Hv+TqcXOiOg+YMbLrZdP87Zs0TAdWlNEgNbLg0XHT
iupKJB6LpySC0KzpIubVUtc1zi3FXBgIv3Uo8SUSxQDWphrHwrIxdFnPOd/pxj2k9FMS5Q+CIOll
hb45KU/w08DBFiufOzxlIpoGmfRwsOihvdbLvuu9yX549/xohkM8GglKOdro2kY0Ovl6xIIGH/bS
QuQAN3eT/xH9IZ5AnHEDFqWi05gw5tfj4NxwDIq5vu1li8f65K6rii4IFHkFYCkZcq0EKI06Ehre
P2Up+8Ft8BBsPIUF5vbQyyPMsMZySLzXIjr2Aw+UPIyk9nKNJm/V6ReKjZ16wuLhf5iroGbxlhaM
LMYRisK8M5RFFogo0yLwCScH0PO/50pHjli8wlVE2t7LmzhkuMCqEANSLeyErfRYE2m1ynS1/Wno
rNn5SicZJ4tIHgrssN7sFdJAdG/vcQ9Hb3AEBSjr07HU6B2KrWDKHuqXdunXFwqtDwRCPxXOOaJo
UlisgDZ1FRL8LXGUohwN/5OS9qVVRFSSo9lCpdfsJn0Kl89seLNUIUdUfB6X6epUpteK6H3ltvis
svQqUokuYTaYM35jrZ0HyrvuEdUKm1MT2pJxvpaarHdKYCsDLF24oyRK7fk6/9sdfya4Z7y21SHC
Eb3qLdjZ0XIB4IR2iIWe1Uoyp2BKGj+jXZxZdcQG/61rlUvv7SKGrPUk3hLfGEMD3jBeVLCIT4w+
HHUlzPhjUHEaApFcsZR2ElCK/Vw9X3ehA9Y8Y8Bp2Vcl/Iap1RVaIGV2SmgoE+Ejf1cp022Q6O6x
fQ2XRv8xcS5eRcJ6/7+jlL+Fyg3VIytH2eW9y5WkZOci/wy63yteTSMDbLn53YF+RU/NgzhKJPYs
fF5KRHvqZCneHIfcZPTUfZxpf8dbtdkDPHs001CXVkpxdj/mdHWqHuuKtWYYsYR8DPBQNWIxXtOE
LdwHcOasebSDQ+zNNcRB8B+XSpwWbsnebMfiqmNfgv1s2b1uxOvveZKOk7bI/e70+IZ5CKGx9/WJ
DvaasxFRvUQND2uO7Y/MDPR7cg0GgPJmv9ojhszH1V6IkpF9pUJW28VSHBketgkund+nK5eLmGRz
wR+W8XPOz/0DHgbNLiw78LPNM0bUHIHrP+nlROyjEUXaqAUTxgoAvuI9LsUQToCFlJw2W6SScmlQ
FRwatmOJ1K9qbPZEmMYnn0opAxnWERStS3bFxHYwJLbfOvMpzOzQuH+h/HzgzohfNiyQ7Q3EJyj0
AEkGtbbxiq6O6muqsUn3rq8G29WAd3pTPZtqb03l3XANe6oJ6H+jLZeM6euE0yjjaJ6oCnBFIGqu
FfLAJNfvfs2aJUVuzRcgu5qR39R5g+zLd8p2FxKJd5ZQTuCeSkVw+ibKmy5S48Vc0idHlS7qgvwQ
S2vVQh4hnZkoSOV3S4oC0YTo6wN7IynAhD1S2XpzidEKUCUhj9mcbOBaP81AswUUPqmwD38oNGFk
e1y5Lmdw1vbyoIvN30kDoP5D+ROPQa1l6PZWtXniGB0wBlah9doqFlIbJiuyotRte+bXujY/Y2vE
PpaKwGWkgMbrodYlw22b0PP3+m62A+0Oy9goRfSXOtTllxocJMJAIzz05tvBRJy3n9oth42rSuG6
cTSXIfTvVs6AFcSd4B/UkS+HJ8BGruYGVqh+fG+keBUJotfuGQYpb1nqKmnA/3/VliL1awjLy5Us
al7BuS3xL1divV92CblkJy5phrq70zY4BVROpkXos5X3m0BCIyAbH94Q98amgO9IxqkzS3umpmgh
Q/yt8WbmdoBbkcUClT1vL8YOIcSxk0kuKQhodEI0C18tPgcmSQ8gOQIdJl1YUVMqzwovRbB7A5MA
HQZ4aJFOTUBTX8frfzWIyJQqf/nQONx5eF3t6IRC3KBWLZlw54kuETNb9IomFvA4gscZaqWQNF7g
JGHFTWs8R0wWvmOJ7A7TNG9ccwbj2W8RzFnzojloXNmUCSr8bhVhUCqvNMyJgs9N/zaVLvm95sX+
s580JczscM8DgfucHYtLYHm4sh5s0h7RpGoek4TcgDMyumDO3Go+IrKyH9C18253ExIyV2ovN38n
j3ytY95BG06PjUaaaDHwG3+BNxP01eyHK1+ZtaWgLBdq0GpuodqaOTbc+i82KXKgp0Wfn7AEHtK5
LfGansyeZ+TgIXwqWhBWbKH1nCCdLI+azds11P1a0anqysIczsW/vDtZlkylWqp3yVLyz9WoCvEt
vytv6DqQMwErCtBf4dQqVVnsXq8T5QVzzOj3UPF1xWLkbv60Jm7JFUyPeZkxftJtIyMr0aMSXAZv
EidSzMsbjTmBwCRaSS1KkCKi85eLnU4dP4cWJLcAPMYjYsxjxeiRD93Aph/LsaOHbHyzwrh9twui
dd1GPpivZOyYBTaCC7mY6f4I2d1kKRWZKRNPS86OPBVnAF8I8jsfjC5zdD5qhq738EUKlpUXmBxG
ldDCjCutfPDgXglDUu61+yk9+tgJupW0zCxwDxy27FunCfCRA/KMm8fIVufjJ8g8AlxOEhFKYStH
ASS0aJiZO59bGkDV8OsuDMoOJlFsunoQ7fDMzHIVD0SfwgU90Sbjc8SFYqJN5HMEFZ3scSA2A7nj
uAEEPEJJpDr4RgZtSlPAY6+lTatTny6vUd4FTkVqh/4kr6PTRHB1TtocMky1rH8jaNtpQt3x8LRs
wiLF6dzVSQO3fYjL3gkIF21yQ60fpcV32lJD/suyMY2sSdufSexs6X3izSdOEI2UM35gtTpKdFaG
Oegje2eB6F3IxrqLEz71ABrDM2Dglq/jvr8qkL9Tji0u7R/aHnTf5I+NlzmxA8dcZ5f3N9B4RD9+
mnTkU2F5H+TaiP9VOyuszE8te/Xx0iLxY2IThn+6UVslgtCHQ3zNGQHvsmhiIiEZlEvTNA/bPiEg
KFoDdCCrnOkG5TG8jLZZA+WDFt+3npCurtBhAkPZmVpxMQykSB59SkvOOewCfxVDN5sEe1GQauc0
LiOPvuWEJTUeooS1zCMXe6fe3n2+x8X4PUciwlsf4MIvxDI808rvp3GndCNo0nk58YtyODskKxeE
RaVe0Ojg2+SDSH1uawCkukOQrUPGMYL5RuugNAZrcZcnL0dNe1OuRXsngBJqQhliNj9D0dH/XPpi
bf8PgjA1rfzWL9uIrtIMILKXJ28nY69niLXQM96DTAhpXsuIfv2d8VanSnfOYF/NLNt6M0lc21MK
0hWLTNOEzThbwDDnOQG7aSvLfez+KTke/wqZKGBaZq9W6U//+/nUSHU9sVmzEP/hfo4n1Aj2slyE
/lTUPEFpX+6Rgxq6tsk4PE1In1bsfvnIxfeYcTs5bz9/whvo9kGdslkHa4SzS/gpDPie3I4SPsf4
YDB6cxuruk5H22m6Ua2AXurioMtxha3hX7tfwLv2SvUwXBuI3q/KgYXCjj3hHTTwxfqhnJthV9ok
8ArnRucZGXZ/fcZKns34ha51NJlWi5c7kandu7xHwlsHxWF6YOocOC+jrMRfbWHCjTcnoDNZCZ0U
Mc3hXp6ozLa1HODU3HOE8uVvxJlG+hjEGTbsc+Cpamc3KeF+gc7LEAV24gAAZoFoq88gTinSYEXs
dnFZSZkdk2Yre//heR4Q88lOkYvFX7FddglHACwpLrSd21H/lIeKnvwla80ktiT+XxU7jl9Ft5Ed
TZ3Fn5D8184oTTzm2d/UwigdBX9PG1vu9Y5qYfBdL5jKr5uOEbPdq6fjh9izjfVeq4vuCejIqQHD
z9GScnhcWR4PFZwkfjnK7qhrG4UtBIOZ+zcCI1jsNRwtJtET/tWct/vMcMbVvuQ2csYiQ5VwLmPi
/izjTHzqhjehaQzZthomOe1xj9sSBZulre+eBpjDFzQuJFP6KBwuR9/c/y0QR3Be5dwUWR5goJpn
7BXE8LgOO+SHiu/EVqJsnm8ECh0HiMQZX9jF6loPxvNXScAF87C+seNKSC48KrIdbyspuO1TihPo
SGM2usHS38jP+4T/k24q0eECdnNfWEMkoCcB0shvfMG/kw9FxbnJs8A1M78BlNaZj7tm1LoafhWJ
Uv+pY6oLrxoLmGpOpcltxi0odWMvESRR1EJ40fdJZyPfCFjaXm08Lr1IBrx4wp8RHtvTlgcJPYmi
ZsYPIMteX9A5eQXNBkiN1S6HSBWbOd9jVpfbU5wZysFpgPA8neBJqewzhIwiJ1D+cwJGuiyfa6CE
x7iddcCA469jA21cerz0OjlS8eXn3Lc2YLxlDE2BewiIiNISGFwsZByuH4vNKyB2M5gYZZYcNDGW
swbU898ccqN9H4S2WMl/Lc98WpAA4CakNCoZ7FEwSUB4quv2STPJZPXr/qPuXbsa+tjrukU/CMoi
hAJDFMS/pEbLFN6XJYCE3DarcdU1JGNEXUE/S+xKlIafhv4/M4wq90H+aRw5Ud59oqNavGqqZLCa
9DYTFNFd8BWhooLDFcDZXA/uCgUq/tq9BW3XFUWkKpSWbHQwlbJFEHbqUkxHbKm/BOqrKvTEHglO
sQirx4fitqC49Eu0b3WSDrjAQAv5OgUJAKw8wqJvr0llWincvkEzp8rtYAJH+0e2jIDmL84vf2Ti
uE6tAjQ5jNF4hr0BVAWIy7DS0zLpikM7pTtifnjchL+EqJWkP7RT1RC7DUrjxxnRHfcfyEf6102t
comUinGJQcqOhR0v5vTsg8tc3ZIvwjtA7JHOYWkrEMfwt/9OLV6ZIl/xEwHUol4SwmVGC5NSjkqv
calMtbvuxN4jNv9yr7iP6tdP64yMQok+noaf5ATbyRyJzoi4s7yfbKFHD35g7jKbgWQYPe9cJ/I8
P5HZoL5V6GZRP5MAxqZYeSM+lGrD5zP3Wo0Mo8A0TyGTQbUKlBQ0cKZr5g3Kr9OxBUQBLjXx2Zu6
vL+iF4KzquXYsXuxoa8xiOoF6Fg5EL5IBm9O5yqoTraS3/tH9sGfocWCrTFQ5KINN4nLF0qm6Mn5
10j+fTMucNc60EZHGnidK8/GPqM0jqqF65GWv3o/s7tHcn1nq0egtdHNlv0iu01Ua/YiH9GnEyid
GHaLTQQ5vMvO3EjhDIn4XgA+rS0RxHEqhT64RWUQugiMVF4W4c9hsVdJDOP3A7GSDBNeHFOJxZBA
k4JQgjHjaQzBQxZ1r9/iBxy2TUrSnsFaCrv0Dh6rAYzysrQBOZTn2B8MO/Nbam2RwfsA83idgfQ0
cvWdo+zzoG2DSsHzxCW5gposi06V70x3foyZIxLYW6SUb34hZ1JZ7yD4tw++FM8pEWYrdC1WqvKI
5y/wQi8Nd/DLuZhIIu4no5qlM13aIl/0PnFZU8p9Sxt8F8AqdJe169OvTlsEpJ6aIxy8qjghhKiQ
+E7LELDqxVLaCDWx+kJK0oNgYMNuCSvQ7TlVtf15nhXdBQhbhPY3peEzft9ZXG/koaCzM0YNhmw8
s2vQNuM2ggpAuo+RsWG6xtutPYJouBOY1Kp6ne3fDkc1k4WnprfqaORw/YNe3uFi1pFHR9Zi4rrR
WSH/fHBPWzBA6vvjRbM6JYBp32+UVHw7qEFsC5neDh0GMt2jrx6hftdlzv8KMPkstXZiHkUPbqMB
9AGKkXv9uEgOD+NhuMOfbuZWhPgMjp/CGztdICDAFt4rz5fbozAe1OXOi9bQPrvW7YwXE5OubB2b
JRRM7NbPuq8F6bXea3k4E8frI4KmSGy5OqoX1SNw1BbIZ1LUNEeWW3n4GJuhXguBBBMWZTdChhlZ
4NPCBFShlOmoNYeb8GhnJQbpQuITCLZcIFNzr4QEMGVhOZ25P3o0nunlpqrbA+QjeEU42xOxuilm
RfxA/e3vztvFeSubodrCDj97IOBHzYkA/nxX9cCg1IuoH5VmLVVWtpeevXKUKMqiiz5/GYj/UlT9
UYImUEyBpkuVupADPuGjArmVQStBia7jCj8y0DXMNxLwiqlWLYI731+OsqFUoAj41fcIeO5p32qy
7NernpsQhcNhYKOgXVD73KjMbru2dYDutVflCuvhEwxTqieSYd5FK2twEc+Ev+eSeaJgG29jkZCj
1uwdb+abmXsk1T4WQgPGvMiIhKiah9VORi2PYdwChkPQp1/WOPkfO2L5aoUl1hl3T772soGheO10
orVgi/E+VAoj8xEX/Nv28lq7Yt0C+ljA3bPbhjUyT+T1UA0UPmx4Mo5PrmrpIy2E27sje6VSeu0Q
m2apIvYYUtAb2OcLf+qvVg1sUzM/Aeq/6h6mO5mxJcwe1JEFlfYmvGDQ6QWBi3ndsLRlmWrAlCP1
VLB/Tnj//0Hc3yRo7JINkzYTw/S1W06O19+u2sLBbpnXbgkpBf7RucNyP+wHcKCS2Wx9FXAKEMn0
ZxWcXU6iT39KHWI6TdlVQknmcs1tnQ4zvk75ZOqJ6n9VxKJKX6xWciAA3jcdumTUwfz0A7RDwSsm
SVjugYTJvGGPsN+v6Y65KeBopHw3iefaEPGvH3gYecRycn8V/aRy9o+xpg0pf3V/J/Xf9aPdmmB3
2Z0dY+vr/wRE015Lov5bVvP4RPiF3+LvULTal89eoaI+BF0NjLQ0e3bRuhFycjnFjGTpdGK34cKx
Henn0fnicoGI02QQPuupFPyqdl4OwN6b+eieki9zhFSfj7UH9K9UA7AifNrFYRh1e/cwL2cmqtcq
hxD+xBquU5N0h1igEZ6gTQCrNxbte03JHRe0A/Gm9c2uwWS8bN7SR+QJwvB329vdh7tI6NHpD+zS
g9U0nkvS0Zqcf1bOcqGXkqlEWKs5u3DkEHKxNnnaa2anAb71tEeaQkTa+q5x3aaFllMXcWGuqNo8
3kPT0mErKBIGnKhiG3kWmjpgrd7bFpI573EFGfg5ru9h4HRXSETYDf3h6jUFb71focdF2IgSBXfS
mANJub0gU6rX7kSZR8wfqzvJMaDSc9GMmrfAC3LhdCw/wMTk8CgV9VIv0TvT5oJKVWWoi/I5UrTV
myYx62hvQ181BNrZJKKwPSiE6OdwL/SgAiijd323Pd9eqozg56gRQfRPAatuqlcIKb/xutjDUMBe
bcdxUDvIapHfqy41aj/80YIdwdGrz+8KffxgMBHhdpocxxS9ar4C5TO9WnkKoTixxnXEoJTiVOW0
PpChgzwmPSafsdy9iLR+lVB9s1FhuQwNOtS0sXqQX1hMgWI7iDs6ECGnITt9WSvqTS/7TOyVENB7
oRmUG6PmgTkRIauoNipsEHt+soiOUOgNzYSQRC6EBtd0v0pjucP27h3Kq1qqf91DipaZX7KuqJQG
aHI0uyZaFRqKHz3rUr0gKOgpIfaTzkvjPOKh+iONrCt8UvV0d69wjr1U5gKYGoGxfGbP9xTc14oN
HIAy2/bcwUQBEV0rtBeW5gXkH0cOKLMN6mZujvzH7rcjI3wQNsKQO6Tt03NGyCZmZeAqKetMEctc
SSQj0kihGwT4Ux3X7hnUwmq4nZFlZLedy5qCIXQk2dtBN6zQDCQDmNcdvNS+HuodbOiG8LRzIC/0
g6p0S4rc+7nDyVhSp1xfAJpKr1diJCPdVpxq2xBFUXLCk8rXBLhebwt4RVlj78vM1kx01auclCJN
YFru/3hK3cxIN3+GHig+48mQpCo1d2nD6UPhg1DnqshkybN4qBo8A/uc+ILQ33ojz6GtGbdiydNf
ucxt5ZFbeDFxeTQ4cb2EfNR9lHn8DYqz9IKV46UuI773UJMBJ3Xo8uschDFltLJybuolvjgj0srQ
svudEE+ZZZQE7TmS7uMpOP9jTwVHDwyJpQMLfKrRTpvL2joQWmF3LRsgjFaffdR6uyWyLOwnt0Kp
7OMZT+6ip4ihXQsN9KSdeFTUrF9qLmIE2EMyQ2nH8PVV4PCBXcetbAWUJ0m8xhzGDxRCyVw4jg+h
AEvSrce8lbyL0rVBySSRcyfoEWQxt/g48jVCfeYgTtN2B1IaP4t/9TcKZRp569PgwAUZgcGgBDEv
hTc6kbAx8AQpADwmg0tBZmyEJaTQcQDBv+fFz3baFk/rsCkNsYWi+TkBSqK3gbIF91S7kXyQCxQa
0NNcT2QTiY8YHGBuP/7vGGgP3+O+wSHuIdO4gqtGqkAqv+3v1XhDwimkKYUSUyINEBhRsAYoozZp
jpabY+jPD019FRAEP0o84Ax+u+SHr3U8V2w4xJ6DZj2pR+Vb6YVuduh4F5dEDMv5gVKjxPBbfqgN
4W9gc3ZmVEEktUYKySHkcGsdo+ZAdXQQVoaitTVsmZWl0U4x5IGC2E9t2z+CTwUsi5//Cn//+r+7
P8fFoY00dXqZLdVnLU9jmh9Fr6eMMZpwJtge6w+pvWiXKYxhPYEAv22aH9U9/Yx6nn92Noh3Jwti
FjnY8Gw59Nh6PPkjzT160DZMwVHgmb4MMCn6qY8E0GIk07BQAAy4vJ92vbhzquEqtd/jKYrKEh1q
z4Ukj4ggzOZKaaHUmKbAPM/0RzY5twzzSuDWJiZC2Dcr/1RJYukCGfhm3vQJwd3HO9x2UzhImntv
sj2jWTk8CDHi9J8YJLZsZ9fbh532ieNfFghL3QGuBcLIpxd+t2xkWlZ2WC09TYeyDonrtAjWwkNV
xAyR1n7ii6AEAL2pLwOCpwZh0ImEFx1q10CEuAfUl4OJEX2cyrzdGgm0cVqigA7JFKrGr17Vy/55
xjKZHV60uz4rISn8ze4Q7UqdlvyPlDqZggJ4yiMcSS6GZIqFQcqRZVTYeEIp2HzpKQeVzt6DYXXr
v7YqG2qqz5Xce93d6jYSVRblfIDm6akA7HWFr3C+ZMlvqilhI2nGPKsU2B1p6k1kZF7+0ICAz+CL
w1MudJflZnnDix4NOxMBJYhus2zhcmPXlRdwJgXZGgrBnZve5myBYlWdMgEmjUq9f9ZQAXCHMLVP
u5EKLJVD2QItbR+9Szq2NylHFoSTRJA4JW7atUY7YfUveQQrNLPJPz7NAJlG0lDk93hndYg0rTWr
bRYS+X2eUzeY1cYM5qTiSRflJrN5qeCJlSmEsINO2f7skbf4YIrIOAHJbAM/rkvMvUlgYxfGWlGp
WwISWR7q4VwBmisdcMYRU3DX+I9BXJPht4fTi9IzG0hajpuDD/Ao/WlxeJAgcBoaqATsqL9R02zl
iV3BDeqlrie0gkIlll3Bv2KBhSq5353tip2HKN88a2kxsyWbFSA20Vj7kkJYungLdZQ62uARd17E
HcTwRqYTVAm4GI59uM+sMlwPAKrAw1nXezI0xyj8QaeEO8TA3JIc/pE+ku2Hw64q0wBtQtP5TsfI
FrWuLw91dIWREDVaVs24ZvtQ9P5iIS9uXcT2sP+/QolNPXcz1W+yB7L6zHhWPmoZDGD9fwx0aTxY
AExxWPCBKScsBebkgu80R4UAi/2CEVdp1wbMEZBHqeN6EkZCL02i6t5omWEXu9RNtEt4GokciE3Z
VkkgdRh9z+Cvm8mooSMReLdTv2bwAvG83M4SPjSYyvH39k+sevsoSKbiA9KqsiqoetrVOpiJ8Okd
tgdUooOby1huFu0v/z5P8Bm53mrxN/bJ9YhJ598jWLdOI54loFG/txzWzUzfF2Pmw3UssdfoCLNf
M2gXdoGmoJoaC1vbT6zbNiHeZbY6b/++z7PtbH/ivw6tTYJOIVFQTrCfxfOhk22c2//F+37ht+pC
oBGRgA/7FrjSdeYr8tX/ZdC+i31DfCa32nl0iw47/FDiI8Rvl/KVGIUu42FLF4CT11RS/0M70x6W
+2NKYVDTkAt2TcBXSx5OFqmuUeyfhFm6LXO2i9M/D3/hMuHUL6N3+MVmgYZElWkcWmV1al8Ob0zH
rqQBlLSyXMgthPsyfJ80M++iz2n6GcpMzKZLmWiJVFfBMh6VgE0URC1WcyiOew2sm1c05BRokYhh
0J61ILnqCBczYKHHe/YGlmStDxx+SfASIR0/RWxJeJFEWc4n5imhPKbwrUJRXi2gxjaj4Ep32FLB
Zdj3+0IG0ja2bXJ6CqmOCEVSypR7VyuXGyrGCfBgQeOZtj4pBgAv4XnCl6R9QiHGwH+7xMdP7SYK
Vl1lxTAso9i+zZyChStm0nKP06j8mMKxy5ah2ko0FYNbxl30ADtk5rBkX3xJht4UzFQIa2kSjawl
sgri6xhjwWnFaiiYpKCAHbkFfUQZU8zW0Be3yJDUZZEahAFVTxDti0rbZm/SohSdLtO65B7wE9tS
0dLJAgZBDKG0z7jByCzthSF++8kHqsxQ+oOnqnlQgH9izx+IM9DmvANIp001rQD40FhoyghGD0m9
6kFg/hfIBzx8mPw5UQP1zzAyPn7rg1mWmLRPBFy/x2o1NItXnQEG3xPoaDL1zmpskSMEtbHY2KOw
OkPQWPmxkLT7e5qPc0XA+EeKNjgxFxdGf3rW8dcYz068PhrieW+V8HwGGb1AXbYuAx6uhn47BBe+
i2gCc94TO9VAApq3IutuQFjRH1p+Fo137JekKPf/eOPRC+2rcotEiPQx+czj7LZN7ZFZQos3WaQe
DrsNDBW5ICjM9biKog2koo2x9PQKD7x+DoxDxtTNvfdqFODoPRi6b3fkeKK3MhB8ldJHLtlfSCWN
qIxPhRQ1QQdKsxGa6AY9D+p0pIIDFbVjCS5pI+WlpJPzmFpYoboFvQ2Gv6wKCX1jbMmh1CRctL0/
rf9IGOo8AcM8IoZbXs8c9obGRzcxJlotstCQb0ba4dbkMhw+xI7WQYH/8umrUDofie9q2br3Px+7
GTptsX0Av3ZTEjAV0wbiEhpCXsFxX47rADKihWyq/m8GvmHNi240TLzfBa2GnGApltcITDtsv39m
4vZUgGmm4b/ii3+yIxNstcFNTYSa+Sgoz6fybCldVomx9J1b/T2EensN3D+917euEko+jRPTVhun
Q9dFerEUmrzAz5B/bLKmEELHMZEQpwTVJV3RroVs4Asi2jWdDtEy9Wpl9bcChMlrqGqvO3xWOfRh
L6si0U4o+q4XfNjEI4Z5DfZ4GX+03vFqSosWkDze4hZpUf318UnUSCYklA39LtLsE0swAQbUu+l5
IoAMN/zTR0u05bUR+xe3bLaRRfufwwEFSDtxHs1ZeEtysnvpJmSpOi6Kg9a6BIkncdqU4aOfm0CZ
xYndTJvecBkNRUXV2iDMUfx4pY7PgAHyjX4Wnd06W6VPl4NulHhsqs7x7FnG4Xv9dtjf+xX/aW4f
y81koRHPkYww9uB+ufnzOzYkXutKUrQ2Km5gm0ZkybwZoefXK09OtBesPLuFVrgg3U6lcMOt3qUg
WVAstPujWQg+bicXe66y5Yjsh4vQGDkNB/G/6vguzZOqh38Ezx3UZFcKTG9RY/4AN0UJJu17tyg1
/+NlFKt2Xolyz1CXRkDjld+UBJriBlCZS6jrRPQXLBHhy20gFnxgWwgKQWg/EvewNmSgj+6VqISA
9HSI9rkV8kDjxzSsi9dFXJddMEzJkkWx27CMH4kqDgYc3WngMeKrY6rnZ2uC92o4nYdvyByA0Zz7
+Dtgjx+AHb692abdVB4SEIdVWjst0P0IMcFETZHXpvcagcXDyou/fKV/DGojAAS/Sw/cKyJfFMQp
nCOtgcVTWdxsHZIUQHXM3jwV6mG88YQ6BgMEmE8Uqo8p2UT63dL1JE/fQjkIkrQ+ZxBI3SJo/h0+
z9cxR1XnYtulH9Im6g2SYVj1Z3I0HsOvRZ3xKu/xixVe+HzvmJOZALNurJdAMBIgO1w6R4hIXHZs
qSpAnmyONYqVihwZwpPvpFAARJ0z4rTs1ycpCWzAxo6ZO0m73veHWlAiOEyEFZTbFZlhOIsU0faN
Kob/8HCvwnD9rvndYdy0fyuJgm9HXrSbWXx9phR2dNLAhwJa0+8TTMKfny+DOLTgqUXEUh/LPvdp
i2d4HFjqLKY1X+lLAcVI4dSTXN2GgTaektHMkpC5e3lJ5LPODqoq4P0oA+jxXGeRk0h8EBRJvN5s
Nm5TdfGppVk495grWabFvTS0sdEqSMhmQd8bm9wHueAohiSn7zn7vtmS5415foXLc1ulDk7vlg/c
K7Igiwz7Ue35+vFdaecayKJ24DTdnplkxu3udtyHzlxHKkg5rlLzGifQ1aaDUOtVQ8hFWcvsnG2Z
BXBCFaB1el/eQI5eRvIKjtIcbfvIQjiZ7y5kyf9RLo671kDa/ExyyiI8Ied4IbWkhI4HFpn3fe+N
STVRZ0bXGgxlQevKj78PNgDnZtK2lrmdsdbeRn3m49wjgN6ApwkyXlTG5s63o6R2sgREYYmOj7dv
q8fE+ITdYW9jj20bbeCkoNnqWuSrwZ65oHFFeol0VDCYvYqcRiGTmuM3+v3fpsEHX0CxSUTmop8S
NrVug6SRFNbCgyM9iq65n20BFU8jEoj821rmvafMgMfw4LHocmFwR7wYN5bXwYSxQio1Tpoa0V36
d86//4vD8o9TdPhb3lcHth+4eP9vvyQfsJ6ROHK6ikIZPnSAeWyj4S/S5G7CjJ4mEYJHvzpUnVkh
O32pCcAhfs8mu+yjRz5GeEfWKBsRCfHipdBIJDGx5N20lW/I3pfi4RiphwkPx3CeHh0ah9GGxW8U
PmZTFOEdxxdACrqSsv6fqrUpoMZc9Uy6Qsw6U4ZvIWNuEIJes6Lxl1xGnhXIq2cSdcBNzB0ZOsvg
ffRM+LwfUM/X3ssWfjMJigSnu4gCFbdIj+BCTgm7bOcKMJz7TZYZlBQ179LWVNQ1ujEhgBuO7w+V
aHtiBmjPsjCmiwT8b4tyGBYQxNj2dmzGN2D5X6TFfZf19FcZ06cgPPYz4xOMvMWxyHypADAXI8jL
JgcaTe0WGU4GwsyTmi4xD+4aR19Z56RVrp/ytXfZdf43WVosP2yM9+afjZSSFRzKDID+Td8b7T1g
j6HdMjx14pyv3na2AQPMpTALgRw9URv9FyvdUhL2YBJU3QXuZ+mHqAhNM1mdioTEnw05B8+qGeK7
Ad3EoJNxXajejOofGm5p+NYvAoT4eucvNUsq+rnxywSuIn/rvK2CMNaV1OEqJ2GGy4mcMR9xHPxD
3SglKiZmdIxkKgfMyoBSsRgP5WHf6/NW0cJSir4FX08rYvh4x9Bbn5Z0mx8hx6FAI0qJmyGHvb1E
WM4aOW4au0UoAEnHhB+nz+gz7LQg3dTgBhCpmC5/dFp4XVGRODA4q8vb6DbULYTz7SvILPf+Nqcb
ATMshMgmiSo2uTBymCzAFyhoG4JO2UrBeNmh662qyhHwGkwtEogelfu266BbBbiRRAdqYQ0K7NZ+
Ids0+ChD+Kl7eufwJb6gXGIBGJMk8xdD7iSH9lNzNtV6Z41Ur3qra4/lXdmye4DpQNK1MYkePzLk
6dtaucO05co+lSqHLjtl7Ky8ojhc0jbxm1nUkxMSRfLcnXr86dFI8R9Ddnnz1M9nQvlnaY+k8Tmb
nKygqbUmYuZ1NPL1IgKkcB/dFQD5TwVvM/Q58n9hxHCl56LOKt97Uf3CVgZi2iCWFvPqFWKUf6HT
/rQAgujpQ8ICTDhVK2vIASyDuRWg83/pHTsDrUhOLdjpH1WQQKDb6O4TXZeFVjcqUs2Z8zP/L2ja
ayGrrEBEs59e48G0GkRQMgndgdsOYJrEcfcqIusFWMcsHAtJUcOSSsiCb+csRDy8np3Y9Z2Ji9UL
sFqKz6pv7RorEQpdOGU6xFQssH4XEF0DADqMCpBHOzRtmd52J8+NjBDMzgRPOk7+d5wVpQ2dhVIq
oKpOSL6ZdwGHt/huMmB6pYxP26uMTEqixFcRAhDvmw0WFXlvyCjFms7UpfhuEF3vOHskLV0h0aYL
1rShX29mR2pVR54NZ4n3nH2/z19+QMk+K5YnVNN4b5HRWjwwTedbcB+yp50IGbvXmxHcQjKpRg9O
ihtVGaCVLaeQRC60OJ++f5fmF7PYmdNJkFsWVNGajQ2sUHGKiZNmHDeHsoIslDVFjgcSQF8BzbBI
R9cN+rBOzKT0JmB4Cvse0FfvrVNO+NtvJGHb+gYHsSJiMO42URcAPnWRsTDO4Qky+1ZPCPElMD+b
NNxSa7BOkD3JBK/lmdHGHcG3emfvUcyfrBdplqF3LRFyiHv9sguY8ge9XIkxnD6xdCvygGq8FWXK
D5sgP5hVXX7ARLpAGdPNDzy/SThzHTh1rvOr6Wpd4qKzgnkF8X7ZFuaJmetcwaZrjmxuu+YJ1y4f
1RFbaafWILHuCRd3PyNwX3z24VcDjgvulVSLUbRHflgnZ/7Np9kjPTka9d4FOrikFzeQSsne+gHE
fKpXg2EP5gtIGLbw0pP9DHl1u19ce7LO+bN4bAnT6HDxgnACGJPfkolY4DdKtyqrC4HqP+tc630m
MHUmLWhZF6OW9Jv80PdYkFnqfBzTBiv652NeG8C5PhsksoT1CM2SuO4PaiR3obolVLQXGn41wSwB
6AZIVgH9bV8s9GvoLbdlgoYdk0HwFIuo63Ax2OmLBBrWKxpFsyif8aUvCs3Xtk5bMeqX1FqdRBFO
C4OnRF0iUqS8C3T6jSFyog5t9Qj8NTFVpRgbLNyjfmz2azs+HnaW2/sz25bzrAO24IMxjkVOUMZV
gjNaXx98NZyVQr2BCMPlNfegbFIPEXZXUs+Wc2z+Eo7/zcAmd+JMKaDWtF5bJ5mTs2c1L8OQT2gu
wzntztBCcMwkU+VCUU1XP5+KhMpro6t8YELMhrsZHGJmK9hQD1Xp3rTv4+a7SzRghVrbOfrpaCoh
Ashngaako1o23MruTURog2eybLwvOG3sLbmKXaSQNlCRDLwxB/EFMJml0NKtsqPiB5lkWhodeA5e
HeQgfMSnO0Qcxid48/ESqSq0N0pFw7+qxJVpU4G9sDK3n0HOPPi50rg2RiBV6SNJ4108MkLVyZZm
uzOlzImOl2AjbOQBO1vZ3H3HTXFFciyW+EFCDCx5FqaDfz/dCkeLzSBjILrPa0c7SkI5x/afgzUM
lga7H0yR6M0RCOL50hg11/snVNCBFirTlNTlx3/B6FDs4KTX7AMgCYMHWuflbXnjMIYBTC7yLVUF
RnhR7GE1B62ELT9WV63YtWdS3g3lLx1yFTHcIdhWGb03NJQKlsn7N9o0EcgB9OyAEuaJf6kL0t5x
i1cu8lYEAk85/Znd/zYLXCVUwYDkGHXYYtMXn6jB9nnM4Tiw0umGPuVvyCDYCIXziwfxtOPE8vIy
BQYZzIh5yt75aiuxQODcfOb8C5f+TeTCewk1Hi7iCy5FBrFQlg+UykBf57noCCPeTsIib26CSjbR
U3TxeGYNnGzHZhf7vLJ4eMmsYSKaCxO6Yd/AFXQ/hzKbm1SZPSXddu0YiCTgRTP8JgXcmqeXlWkv
x2tU9S/L9c0s75c4N/4pftZPBDqXlh6Ks10dM4dJUADQU2efVAL4hDtmIloOghzuzDcMBUW/Lrdw
Q11OEsW1BXjsYLJHSei+atMGqRhu+RNQjyh0t5Ftv+XEsReSrr4pptomm4KXXqtZqisZJ/rlWLGW
VXNI//cwtRzDvuFWJkOBW7EzvoArD1hvqtvwFlQFjChq2Q21CnaHg/xrDna2iJi1g/Z3zSffK1oG
bdoX7gsGKJQ9cfuEmesKJQ+brCtdDNOiS6x6idbD0wmC4cf7x9CqceugrfZJJZDdtUqNwTEofxN5
LyWZMOV/ltMo98nJet7X1mnOoftDJrBH5+CAPex6OiX8k5GirlCnORCSo7Ccq3AfPlcIOp/e6idZ
1gZbuG0P5mJYNpkaUYjzAvvUl+Dmtn36KYl5wBV6FYCcJEW4D6Oy2Idt4qRwXGL0CFKk17xoXH7e
cWvMTUmgz75xVescPAt9tGSO9uD5FAmMpwCyD8iyJo0Uv68X3Pbx1vaZ9ezls+TiBxVJjbuqkS3E
N09q7jaTVHjZbQ3G9i1395xiQeNtOLj55mPwWV7q9Rz0uMRBTp9zNCDO9x54+U/N+BJxHaf+MH9H
HImbb5m/80W2flam2qOYU+sebgCnpH2run6zgfKM9CGWU+mApAuNI6Cb9EMWYWhvhv7EIWtxjpJb
/FtZadZenzYQkBpyVpqTYXdak+uHCwKBdPvA/ZcX/NCi9tgCkFtPH8BB2PiEM6V+TZJZF+He4aly
MJJ6tZdyVFPheMkfYInFwqwBH57iWS0f9lGhCY/Lh5ZQcYmJLtXk2QfeI6I13xv8YFa7TKQgR1dL
9MYVSVLKKMSnJXD4llIwxvFLAkwlggowh2SII0l+mp070lUxWQoNYNw7ee7xl0iDStigVD6vY8uU
tzFbBllEvBoZ9b3aHDGI3xmuHBbOrhxkHQk7vkqbMI5j6JDd+4yUtlmVDIKZ3eSQT+GcMrdKmyC9
SRoBHKot7KN8BPqlhEKerovUrUUURi0FexQCVIWizoMjoyL3gE6wm8v4EDvbrcQmrqXplvV2/4gV
Qj7aDUH8lM6CV3qc9qu+xBs+7dXN7lE2aXzheEnAagzbNINCxHlrf10bHxFn0uDxjuleQZfN737m
llViY2Xx0UDK6PGQICWuLPdg93QJPiMefSr+OJ3H48Fd5hglRJAHFnJyHBk0jqLRY0D/JM8nfBUh
wbX/CsBfZwKW1/9/QBpRGYHdZygdq2Tuqngw5VyIvDIjAhxyPJef+SxflfUy5DJLKxIl0gfvkC6P
1CJmDq+Si6Zm/cVyOoLuWo08VhQYlwSNYs1aiFO9nz14SP0cLa0HhGRodT+k0Yp+NQDtRRq/Mifl
PRRq8w6LC0vDXwZMban/pSDGeZGqh0MEtfV/2JraN14xrX0nYVU/cfiwM1c0siKSz/InmEDJ8Dej
VuPB3LGmtXjsC5K1TKuKCECUGGCi1UAkoPFqH5l/u0t3v7F7lu+lXKX04zMZk69MnIavLvpJAViO
+VgY7SJ0pEDusbaH8crRqcXU5TVTUbVLNRrQNIsLrHLogDl4En7SDcV6h8i9Imdpp+a8FyU0BNpy
aUHXmwY3aqkq4E9dWE52IYUca3UdQ3spGtYB/bzEEvWDVH/ENdX4xHUFr2RUttIIesisExavdmNG
CoOffEga4MGjhVVm3ibTOTu4hX29FnxcuCS3UmuxkW+1HwUxtIlTuqfAor1/ebPBaw0/WR2qGfYY
L6DhjJpwhQpUdPQf/NwxxtjNZX0tfDVMK5HdqCq4n1buqcDCZZ9bg8j6N2+E0B+9PzPvvCdoKQ1W
GZNmDyeprOwqMhVwuIc1fn6eRGnkXfA2XWyk3CgxAI7HU/j2m8tpOjOGA2cxSf2H2emXC+YL8nwf
JFXoRrGeAoAN/il5Yz+ykzxl3w7fBEZs22t116TNnDCyZ7xU3mtFCaAZDNQFW0UdObvxrWq8I6tS
Dghd1g7MG65UOLsyTCvUk2WZ/Z/XG/nWgCb9bORql8KOzEtCHUqae2EPJX+y5kmYy8Nn/EoJj/8q
626sdi7v8EDCXaejPWKfD64AcmgrfGytYI5UQwq3VUC4AkFRlRx+rBjzNaLoRilH2LyunIGYksF4
G0kzUu6p45o2RKngFjQAxA7cop91pOvUeBqpnA1G7BbFHoXT/iYHYsCINK0EgC2CA/R0iZrPExZ8
X0RTg3LQYiDe4UC54L5K7KMx85Hffml/JCQJEs+jkdhewz2hvaJ2x9RXXn7ML8klIZwBgmdXthIh
reHjTClFhBQW+PB8bVt3DHv7wJKXLWUeUD9MMjZqaklLoqmqip3AJKLtFQa6ZFUiNQxLJ5Ys5enV
2YpLC18LiU2rudBp5lRywn5vqLF8tFMz9vFZFmKX6QgFNUUx7XsW4YfddcOWW7RaiQkdOqYyvGcx
UssC2cXC41V5gze5FEh9kllPpFSrmdDlPLWqm13UuHc56Lj8XwI/u0+GDe9S/hY7GaWsJ7LHI6Pk
c5FqQ5SEYb7SuqdK70Y6vTycChbx9reMmdXzLlrStdxhkHpNpfwP+EMA3D4+Z8qNF8g6goXOGfBO
yHdbkz5gk7X0awLWOXTFg5oZxE1HwnF9ssdOoCSOX0dW48E5emxZGNY0XzE5D7TRjKnfI7CCax4l
uCIC7kswvTeVCFuWfKp4bOtanAboejOh/63lSeiEK3DKA4QDNHW4h0FSC8qnvzoTjDRXd74rxpbL
pIrDxn+w0A8mKOO6cmFltb2w5+vIEpLhxxRTQPKCNVpBecqKf7cmwDbL2TOTsiOQ7jduSRtCY0m1
Zp2iMiSpwa2FBDzYKYCRzAOoXSV1FBo3sK66S8IHlp/SjZ3p0UvEdDatyJFaVMNsiTZGK7RUwQR2
jvIxkmEtIhfE1AMd0YSrox9HVNopmcEOC46p7j7K+4nByQY4zgUwvIN++a2EUt0hkP1g34bXnYfy
hkqCg7oJUU3t0zBLhR+rMpTTLgMqBjz11jZEaUeIyOSs9JoHGzsD+wRABr9Zn52OMQG4g4zgXFVI
tB/8T+RaXLZWTIu0gHfDAEp74uHVrNA6g6GQun7XDzuwPzPx1Hj9/sZmAXzHEIIwXYe3SZeLwJYX
aM2vlZneSqwT6DaCAS1LvoJur7Np6S6NXWJbzGY4hEvGkagpNf3BngkUEpAoXwSIY9FHG50IXLgj
Nvp71wfNOvVVvkOsw65n3V3ssBf/GIEpw4CDMvRNtAMX4qGsCjicldfrkLL/T8/OggjHKiittI+6
pDkKqluaq2g//kdvHjXptoldg1GZFvqhtvrXqCPgxuO55wBdqluC6EF3jaV7d2pBD7H46rNylywB
6dxSGx1XpIzN17hw0mXeFMbgbeeGrOFwef7Cp1q9qD/Ay2Q6l6hK/MigM7v8YyBLs0i7wIjhhGQ3
99/hAnPcZO8dgNeHK4iOL2K3WO4eCGDNmzzN/ZZ3GdYHxE0xF6Zor1+K/ulMmZ12iwmjP9bQ9ykI
UAmlTfAeb+F41U38NtBauPkfe5gbubakgnuepmERhYbsKk/X4Q3crR7BhamV59murSHTZu/4f2+P
VhZP7w3SoeU+x4kBbJEYFl+bN+077IKe05Atnw8DwRGMXDRlTkHGcH6pNG7MH3KXpJHF/ShfXnlM
LvoozDBRnnsYvUmCEIrFJaFzwMm7gp3+JDmTB/QE7mw00YJ5a+okTEZBcDeWAbv/v0F7mEfNW9aP
MiMEX9XYF/8uk3JQoCWiBp/AQUtFUwNID/2aeL0pu98C/zUPbRFFpwNL5WEkcfJKOj9C2mOb/h0Z
BfMElt1pA8XU6D3wkGf70t3Ix9qb6XH5ktPrCQW4rGJ08BNS0IxyCeRT7egmA0HbK6Dx7oOH6IfO
+vJVkBDixNPbNxWtS43bm0/T1ajtUSJz8MFIdlUeuUruKyqU12WNND6qZnLD7iNOfE/JR4BTvEF5
VtIORD7ftw7e0+oq0YyR2mkChwUA3aBxqCptFj7qegpIRhgTaWHovnmKln7HzKELVxmc3iBBjZMF
5oBPEW6bF8q9vB0aAVy8V2eGvDooG8wCmuAfGL/G5Tl2cxnI7nBFRBs/zhpBYGfjAtAly+DedK3X
TH0H7dVqEFFQiWglNaStSTGwo3tds3l9p3oNCWRblWBEdT/7I0KUcjb8sHtlgwOsKxomHbnEddII
v+gqNMy5eFXDvqnM8TgzUglt8H0HWN6udYUHp/P0+jBSVqY9EgIHNJYtqI+owlFrMX0T5Vulf/5J
0oqjXmM4/QZBXBqfr90LbIAwrqxvxF7FNMSXJpR5Q/K45Dfsm5QJACBRBshrnH4V1u9UHh4+lp+4
mR00tuYCljwLFWEKzwnQuu8Mf8h2pDGCsKtLI3HorsXlqFrDaocPjQh10Avi9zJBUFmIa7wIG97u
f0AYvmIJaJN6ed2H3yuJa4LeyvSD3YY0RCGDU+4n5UYZVOBUDBZk7BSjTH4srUEd+G5efU16C7xW
jGIPi3GcNOcLNJWQw0B94jlhXbOyjodxSIWmqarksWOCfclL6/14wreYR3zPFKWeNiO5bD27/vv9
9HSbgRIAZDPBiPUlVh4hd6VyhkA81wN6z97/tGPZc7AGO3jbfdMGrHY+pRSfa9hYgBmNvZRndShr
cFdvfBU4kEcrDUtbEGFPeT8am/N/5c/pVDkK2wxyMbM4wcomlHvXN4yBhpiW/tlepCn+L39pRZyE
cFw+l2U4CKXKxD+T8fCGhgRGVTw7Jm04NI4pkJaxfA2LkE6IWrCL503g4+Amo9aZhVG1/XP4FfI3
sqvHWF9Em+gKCvX7IqlR5D2jmp9/FyVDWoXKyVIs6Se7O+dFOydgde7Y3t6HlWPXGKXC1i2TepJP
gsL/zF0aQvAVrpdGIk9NsjEZpcATTWvmRczQacLlNOs8slKtSlki2TpTEZuCk4C7DEJ51jz/DLqQ
xDl7W3lXqjJz351zMwcj5QZ6aJf9ONNMvN6CPBUafNB68VmlLL2WVmqcs+V5kU7UC8jtDg8Mutfk
siQLPCIPhSwyp5jCkxRpyDE017jSziTdseJuWiZeJinxuiRT4wlLJ+ibcEcXM9kt/xjWeO2jJWoL
PKGvilLe0BVmLIK5WMJjMoe9FF8AKTSSTVyZ8rNp+vVzGZOFk73hvrvUHiyuo4wb2Xajf4XNJY7K
w403r+80nUVDwChBPaHUZAjJqUzrMGk5F7Pcqm+F6zFwsxdTB2/o1UIiC0ZX8apevwbmXPG2KjTy
ffYgJb+AY5f4VVEx2//0VIYQ+WvJFz9vGctMqfhwA6jfdFO6vmJS6rHpE6dYtRopIeJlOCM3Sv4s
Ol27rQMthxFi8C9cDw4YZNqIi7ZssAB8qOIkAhKbcD7a3aM6Ce/QdFoTSuJDyG5lvrE+afUvbyZP
am7WRIWwZY2HIh7niyEEb9WeSj65Ws/u3HRx1WjmMfIbDiwNBvOuZTqpUPzCupGmUi2KZPnNVQUF
MDuGMJAKC+jh7QK3/Ikt7yYzNODF+1m+iTRpq+ezTx3mDKS3LljxiAjEo9laFCU1vMlFa6RFRpqv
NvygLztn2bfN2ejfhNwtmfSx2Am4jakPrdl+xr22PN8sogLH+jA3Jno+sdhtp1qRjglwdrU+PzPN
5hJCOkUcWjyznHHd11VuLV47xtfm5rVdwJwHox827EWuIx98B5KYeN98wKIb44UFJy7aCVQYVCuo
8Aaogke0YCNtvKfOnvkWUKjnPJiPASUeBzdMylgJ3qN1DugGzYxb/tcxyZ+9rpEM/7PdEgyd1S6T
W3F2tpZ2Hl9V4qr31h0bg90zA87u/9/wnOYTlUSLW49jBZi8SC9GWS2YshbM/oja0pRRpQfChmGn
QwyhnrNqFbA357UIHfF35wFh7vI5hfP/6i8VkS5iKr7nQLAFcywNmmJMgu3mgg0y9nunWxJXH0+D
w79RQ1xWEmxYGn2kMj+MR8Tr6WhMwQXLxVo/bjMbPn+A+8Yb6H1WZ1oOLvQJbdQOnEfq8WVdV7mN
D/Tb4HEQdRIf4KUzEue7zNp7eSwSBxn3l6k2S8wHxgksS2mlR14aerZiBJspcs81RxSL7WjjPo57
vbgg36LhIBt38AFzD4fM2QG+BlxlrpnawffwAn4r9I5NFMKLK4lWOrLRGOujsz0QIA/z9m+8+Fbp
pv0cWrCbvN3U8nIRxFHoKHhJtUwiNwObnJrYi90FMEN3H3wpDDfF80C3M4Ks01ouxiwQ43VnhDic
sqFsf96CxY/dXcBZehYUp08gfUj4XvcpEJ308p8Y9V7vj2/SNSR8Vg93KUrBc7Re118lm1NoHqdk
ER2Lyslv282UQmlqi41hvT0SdRVw47TfP6p0ObeIlwVdUtBlIthoqaUZpnjRJJmvf+mG/Pcx8e3a
RzbKugxfCs/EotarmiLHdTN6KQUq+4lXqhO2iGrQ2TGssVzxOrHe7E/dY1oY+MYP6PJkTfFWicUa
ow65q7pXNtgI4D71yyVbKuwhIwbZpQ01P29fsNaFSoJy+Nm9nfy18349gdOSbg2Y++/ymoiijJ9K
I1xmRTgA3HHYtHCO0POZ3jGrg1pdfxCAZLbRfkD4d8KAcqDSDwViFcTTXs66JdL5lzI4lRyDPKiE
o8/OlD5KOcVlWrfDrvyxtfkaFMd78yaVrp4Fv1oOy5kZYCcAJggyyPRzjnJWfPhJnhefkeS+BbNG
rNbVG+23YuYcbbrFtTaovykzq/Txn2YGK3QwSZ1e3BHL32A1vkbitA2pQfKLhUFL7zPyiY/Qdiez
2m918Lw0ZMoGHyMav4ntR/pNXJbH+fko4zEQcjBdVqQCVcrAiz5YsCFvxOGp3VW1FaiQzREe2GXP
CYF2Fvd3eQvC75xqY/i44ITZj6l8EL/Lt4C/plg6nbgQPI4R9LWLCIPaK7CXgwDttdDAyLu8ujxJ
sUeY+0oOWlMuj9wGapYQCrHkOWwVtt8/PZmS8E55Rd29diElACLiGf+TIFLA0XXUJ2lXrGbCQPG2
wSGheSSl7uXYeZRCAtqvUeaW21Bl1u8rKW6k+0FX1gTIUOQ/uk+qut0Q5kYTlPs6gdjUZPL6lySv
bS7O2gtz4njwsw7beZMDDCUtkWOWBZw06wwb2WbsD6HGTUttxBcoGz5jX/p2gAzoy5SFbdSSQHfs
a0AA8ngysnf6Cw+wwhNYly/Os4m/+rOp33amWywlYrQkwtKZPC6XOUQwEToOYoxipbXkBndHHv9A
btbt5UNeVlvaww3eia89Hfb7vRicLNIt76YYIfR1QkzY/XmXMovK4/6k1nCl0KAo38gYLl8SSIEd
PIh+t48A42fNqNP7xmjnH8bIsH7W5pyvtcr0nNN/Yr4jX2nmVIrOuA9pSr0AkAP9+xRYnb9TvXzv
x6//kxA/lyDSkl8SP3u87QyxJnBXMw+fUolpkaOeLqkzTU00wtNU4JNZ1L0/Wr15EZvHyGbHwyla
MSu2tNSr226UnaVQYKsdSJbQ8qTbxUAZn5vMpnpvQdGVnuCIyELjN/JD9CoYBMR+whvT6sEcstu/
+NLmG2MtBebc6Zwp5yV/2kyqFJgM2wBNj9dVuJ34DQkgi0cRsoTGxoJw4ptD6uIqi+LUhLVZwUfX
Bj9EdM+zMhBApU5pA4lBwGgjW+TMBDrsLNgKd6lWI71nvjdA2q4oI1rFKvwlb6XVz1ul1DF0O8zt
ng11RId2TZP3Y5MgIZ10Guk243Fdx6Fddnmw998u8jsHNC2V8DZ1nJhly1mnYf7BxfdNpFIRcGv/
jbgOR84RetQrzsLOCe9BmMF4oVviip/IzUDLJOGBQYLWTbdxBEKDPdhky8I3+aetTeia1EkNEfB7
1rRSAweCoqV/Yp70Tbeh+SAhR5l0+RNVgzu2HbupmK4TjyKxfIF75yOf2bFpxcG1AurFuZGVCeJY
2dMxKd2XKrEqEf8K3lduXUGrAr/SmhviQBO8qs/eKBTIb82kSn1t9peaUYVU33afAjgI53RvP5Ai
SOxoq9R5CSGqp+qUDFsmYeMMoiO1q2TTAT3EO98K4VYA/CmCinz3Zkc07YlAx1fBGNUUDhCysEQp
m3NlFTUPRWbc2AHxP3i2C0R+pGrh1DTLeB0M5ZdtWiR3ew/TePRZCnqWeL2pmJ3RaJ9e/41xnzz1
wTqqvHM3zsZyiJ9iRY6tkmKPAQhNOmlINmHXZW0JL5mVtcAKZmSLV4eHBzWiCZjbok8trDE/BS9M
zxxQlOq1CTAUiQ/RfskKJuIKbU4b53CwbLFGJgnMw3cxsqSYaQT98GCIuqbCHRy75WVnugQus7u0
ZC8Yr7PSMsFld99izhpuEVRoqIKka6VdpW46Nw+lRIILUVYLA8OvkPRyQAJ9tMGw4ewn7M47aVjv
dExAwc2DCy7q0N8LF32ku6Bff/89diUtWHLpx/aXNjEsYc7yA2sByNKPXBUBH2Pu6PGtAeuamd6S
rtKuTDlM6hj/Ar32yld9wWvX1nMgVPm6BD4uY15vkq7reGmfF3agDhDffW3Wkrf7wtRJ86LgdZqX
Rs/e2TilOTPTeRa9xJd2PbKhFe5eNP4sPTBb4+Nwb+WogwaiaXYEWdLRBWPJpfYhH01y3G983Kyq
APHhBFY2i1jOyPxZ+2osbag4fBd4lM5pSBxGu6r0X4rfdQEZDCznDJA+/G2X/JG+z3OHcusaqnSH
ex48eLqGw6Zfbg9m8lmBWcuBjkS5DqYhM91tpS1fkJdLglcrzvEeyGNiV0PrIqrMqHfu/S3hsF/E
hDlyXA3LByMv+7qhWwQwZkuWsT8DOajMRUl9fL6i7sQfsnsGdSXyFX/fVJNP9wPVkOWY+0ebpTw/
uBi1xbUdXW7IoDodnTnQBAWoxtTBmKy5Wmpsa1CntVq7emnuIyHUa7x1nCk2s0m/pQ7gDs6F4tCy
aUA62G3gUCq9amNbW0kYYKpAj/ybggGzJ7HSd/ZPTLfmihlNaeaW8+rag5NAAFcnosVlzfljibGI
9ShCiVChY8lhl24ailKShXsT0xLjL01NqOoR99R3bXbzeKCyLjEe0swjIDaFrMKpgVu2kcW3I1pE
FJ2xgtbxvf73KTC+X++KLHqrfpHdYDzfs+wRPD4ZYvi0phJPJRRr7yMQsD5CScRfTlRrUmU1K2Ol
p4frWljJ0BbIPdXOX9YP/cgR76p1R5a0PzUlX56O9SU5IypDbiNqcHUuj5WlmCqJsXQt5DTM6t3u
W10CXU9kuEmVQEr+QNUoSlKo2bU7HOGxnz4xxvsOvz1mH0WcqqJCr+EP7V4uBrhcrmopP/ZB+cr3
V1kVheHibh5YjjuzvXGgZD/tZTbPPx3tEvAuvA5CbRLbb7f4TT5dEYTS9OekvJUWG9h7cqcCVJyz
F5IsWFTmC3WXejJZ3zwa0vA8ZkBnCAmK80iUppmkIdE5/58gAFRN84R9dUlKO07UdqrIPjeDU0iS
6+Ra/YhIH4O5y1/gHxJ1xUkts+8oSxdvPjt37dxQgx/ZrA2/+OGnozTw8/cqrXb0ASahYsQspeUo
V56Qp/HRLiwvooOI+Sr9yLwOSHJhheRVBm8CzkBHWkgBgcW86835cWP9VBUfGLNRJgQmfI0g/Ynu
YcX3oskYpnSOoS9ND9Q1oXkW9Cv21jHWvEQGuJljd0Y2uZIcb6qpgfdwalKaoMnZCNGLJz6KmPzs
cxG4t/4q68nkFDrI6H9g3YMcZiktO3ahDl+xrb6BlVqSdhwJRPJNuUEkEbkN9O0JR0kuiPIuoF8X
IEFcFSWGZvPZkDBfaRjS77hq1ZVf1Eo6eF4J1J6Du4oajS4wDsbpyTfkTkTYjDsRxyj1f3gpFPAv
6QywhrG6H3nFcWa/hfjamq6NfJVNpCxsOzwdgeZlE2VGUTzGZRaQpdEr42Tq2Jz3qdoXTFXOLqM1
kqQ3H5FinXJ8r5h/6evoou6i1JnKsUdfkirH1b8GG0fCn0ScRzvbMDHnG3xZqEbSuVfxkoW6yiai
xROsc4Q47c5AbuEKUTqjmlxlUsNQoUjX9YKY8ymK5BYySW38dwRiy16NBTSvG2Xiupr0A9w953AK
/oRy/FPY80N7SmK9JqFPwosPKbQVSfM1uXwVcR7X1ycgH+ygaeS7v7bZWbdHUg2gNHCS12mXOoaY
P3mzCxr5Czci7GsNuinCohlIgL6dZucM4Rq/fNNosK/pFyj3xaldvMceXWqVomUaySDsubpBOX7v
CEPvEbYbur9WcLTG72nBBPgskDawZqtIzKUx2WcQXpT6kvmrAbS7xoq18BzSOH9HzRGiPp2xIfgo
TwJZhkhReJiBJphJ8jZA7dirFxYeWk2rCBbMXgIH8vZRUalPBbbi52iGVD60d+SiyApwFv88ASS3
duwa6IFSpBhRcGdNAOVpij3n7zUJlsfeqemB9L9oxk3B8wj3v1PgJ8cIFdBSiOkzwJ7t26kKiAC8
uvjcM7UZ7ig4daZpSl0uAvINzoyvkjInX1z1PkGcSaPl9NXFKs2zP4LG3Gva6keRogHlEUYYV5+Z
xv7wDUqIo/Bq0qNBMerdsXD9Lv2+KsoQH0qBz7O5gMDUIEwftIR28rEYYV/HN8IiXMchJgtFjE9O
2O0JHqrYnzAFsyL+u4nH8/E0zU7TrydqwLqW2bt8M8sT7KrL7iv0wQau5fncw3/zMPcCFy63k5Da
TZqEMvTi4wltbh3F1HD5HHsuWenA1SP1k6R3g6M/4MbFhFF7f79ZiwN2yuZk9NXORnE4qQDCayPi
Nqa6UfPFxncTU9EwAnSJ1Apx3x0ApDa4mKQ4a+NxxTzhYZK9Tj9LtBHIPhcm6vvlN7URLSeOboZL
2fSmxdndJT5zHwsxBSgb/ft49wKXKpI0w/TlmFFpUZq/91xcCfF/p+Jwgak6pRh13THBsxPBmjzS
pkKdd7xlPIMcl4EVarcgXmCDgWQw4pckblKEpWj4wba5RotNuyPci69oLb6brxNZEUzdLWqtrAlS
vuG5XmtfT6coSHUZkFdwb9uUNFhbn3B+v+BXjHxGYlLUx6J6e4u+IE4cRMTW5+Vpf8FFntQNlfoB
ZWSsO4tH6YJZSQgUQ3Als6ieWE4/MDRUDaCEYsJYjc/k2+zeE1dX8kkH7ZYsxBcU10BXo0onp1u0
L0e7XaySs1WystfNqWAJvk4aCLBL8Hj3se6OTaSRtKva2c9bOEJVAwLi+LM4Q+ycZ6a1x8UGaTaH
4M9OyFeQ7bs0ePpZOE0aqQkIsq4kFy6NU5Dggyb2XWWjO8/oQFEbmivBQZyAk/iQU5dGiOMSQ5CI
vJGagZJYBTbOTlhHUw1sc4MyLTX14QXDBdg7b4hHYIdz202PVTxok1WeLax18SFswJQQMzmgzbrD
2jKw4lyCVmHUECXkp4Y1crH+XweFpd19KJ7TfuUfNg1vHVwXNJpDRsqCcijwttCohiNPIslJjWUh
vatlh3FpSlbWEMVHhR3d9dTDqt6PZZljKM5NOChk8VSlesg9qRQkhiy4YqL0ykKd9v+ChGs/xhsT
0QTnueeKzQZMSOs7U3tQtCM7U0+Yvdj3eWHmsuFD+7rC97iFH5PZvrd2HUfUPfURh3kf6YsniVJe
GnFTgJbuSojz3jxXgkwv1Kv+82Zbko4SEJ1JyYblGZQc0CpvDJyV7vBURXXLRb63XSep2feny7p3
u1bJbOKblkt0BGRIUb+35vuqUEH7U3rcDNXgHyV2KMixJQunsU9dkI9eScErenSbBcDMmx6k2E/m
+8UsNfoWFSpqeeiIxWgNBi3/Bdx93hs3+qAxgg7s2dF3KILXuywdKlwUHoX4MAwstf5WDceo+1Yf
TcPjW5fleNfqxlgodtSflzt+ymYZG2z3U0zv3nDCXi/WvvdMhm/W3t63tTgm5x7nAGgTTRB4yYx9
7GsKX9NoSE1akf5/MGHLORTzUOlGzIWXjK3ZmruV6V0svAP9lMa34yAtmfyAdHWJIga1dBKkegNl
LAnJuNbjIK6J4PjKAkagRtmf/WV1lFqeCrbGyn4gousTDeDqxWa6TwWa5Jmc8nzWSOFZUt9zhtbg
ZgRcnWMP2b39385ygz7iPSQ+4jWeYqMhn/3dFP2bRrXa7twi0piO2Ec4xXc3Fl+XkrBHTOxOnaPY
+TuytmzzYvtCyc49yPykrlgmV3ICF4mk90GH4+BU78KAQQDC+kgv3bJrvJF1ncUxLUtL/OkCM8LP
hl2O+cTFOnS7q3p4WeH5KQ3rz5hcSVZvW8FDYLTD3sIoFX10yFsOp+lG7mZZrDoSMGxFEh2Xbm9b
fNNYGv+csuoZi/s4g53/CMy1aajSpHtC48xRVWfHc+Njiwe4oVrgwNtcwhDGaWTScLKI7LFRqj2S
uizcw4MM4UTcV98yUdNV4Z8aetkCVd93KufscUMmDMt2LUHF1SqJEIZQ2xi7Xtinmm3fjxkOiy7O
Za46dQiPN0W+Xlyj7JNJlslF+9oMgJDBDVXtwM5A67+juH7pN87/oTSQ5+X9X04lYOmM+XpCPtEj
53yLYAaSY5eMnIQELbO8f9raBWgB/T/yE+iLdKWfVU5XBBEP8vilQml7SynC4w1og3prLh4g6ero
tZZVLlh8oh1Bcqz7OUOijdxTnF63Y78p/E6rFTQ4P9VpBBgWtGJZ0NnyK0Q34lPHcwml4D5mVx6h
y8ZPCbRiYA4nCCqN8cvdgUnPYFbKdVFW/0wwVxRyRlXN5BuGynum5wWQbcTt66n7vj9XgRZuTVmi
xD2zMI01QmJ7Q/ChE1x3ggO23Qb2QrrtJLtbh1mxE4BSr0JFkmR3hPtDukUa0k3c7/lYSbQr1Vqc
k6RQ3qf9xoq2Zy+3Lt4I1xckC2OKdONaHxbn6flLX3hzfas7RcgoC878fG4QCq8yjsQwdT4KlP0B
lsZ1sKXogdtOfCM6VAjdxYPR70G3BNam1ZElADyBkk+WjV6solNtFgTR9aAukrzy9c2Y8OosCBRm
f2UQgVzLceve2ObZidTvdTp3FOGuJVJKPfJ10C1IW18lHbE+z4wMurCTVQZp8oQSXfjz7YclLiL3
yx/aCQIVJ5Bf/4x4jdbkqNuB1L2R3YioApoQm6dQhxgElSYEjJSoaCup8ukFgpob1ROQWH3oLHml
rQTdcQG7degS3it6DxSc9qSfhbA8KiwrJ6wG8IJl1lv0edpATf9ZcCoaHyuPkFgG6CgAaPTBTXqw
fGVyYjxGHlh2r1ejXogtRSKoW6K+lnYUuvY5xI1rDSrlCWKV7RieZLO9+FnJj0c4WrqQ6E6waYAR
j5RFARZ7H1hQH3cxGA7oSjaDmwoMAxUIUg6CCCAphBUn11On3lo0/RyUmvAPgScse20vhqb5aUck
IR6QuSN07Pbf9tU5BQF3sFWvc+0I+qKn/lGWm75pFdUmk9lWsjGaxrfI5TDQulKuA6Y8njeJ5esL
1Ql/sMF//Ac99iGWLGLu0xdau/t5tI8hL7joq1O2rSY9kwAs/NDaL+avU0Enk6rTsjgV2VV59qwU
PugyMAoz9hzbp61QQRelvog0KeRboKAQiR/srpqilYa1aMfwTNPmqmUm/+/HZZ/2m3P6ExOnQAUD
3fj6zD5Ogf807mC2Z/Di+1b/VuQN8JhYqzPET3ctM0A17tT5aMCNtiz7Mx6R1E5BoU/n7DzdZ8L1
MZQieJiprqpmL8IVyYEg04p6FfKC/Z2sRFxso49pGfo+ea+y/QLLGgETi6TF7RxOfcI1r2KcRWqG
x/dyBczixe/KHUfM80PxIm3sFO2tLy0fP9uPsI5ikiEokZ6rO6PCoYfYJALw61TFi4dWxdkvHI5U
c4+y4fJogMIAFUcvmEQ15u39m240y9fP2TVYx0gqeBcdHpEh+Gysx99WMPlogspUvQftVxZl6ZT7
0n801JVu9LL9krF6RP/vs4sNynNBBHDBG3Qj1p9QgJ1LluyFCMteOSnBbUjYdW+gC3qxC90b/M1k
M+xeb0YhDrgDuQ4XpVOQROZrU0wwfsV1V4m9uXKMpB8Nf5bdxmdhyWEWIvtuNBT3CkuoKt4oK7cl
pmVqniF5W/RGv3gSC5wOtT9a/4SN79OaUF8zZR7XaUh59+IqRztZD8DMki7SHUdcAqiTl6TMvKgI
buauUNuE0lrzFgcWGaTTe9U5Yl1oTCbAfKGrdAUX8qkiqkDd3XtZC1pLJBrNJK+KtCWAJenHqGyf
JjUY0FlXJA1UtmqqHrd3/PpDyEy9DCONTDL9/di8kVVCwSlhQjDWQ54j8ESNCtL67a9QD6p3z+xw
PHOcJzMLP9p7oaZw2dkOpRL4fWtiTItPWzh/r8d6taxoJqmNTUdMjAVyoELVg73WKewWACd0ORz4
lhy0v/aKrZ6JYY/XT5dT4roYFI1seCcTEQq1YtpJ0WDICdxIbE4LqTDmxwcS4ahJN+cHmPYD/d8x
4X9LxpSt/MaCiB47bgx+L3qAMOtLa6vNWVsw1ytwRtjJx8J4VGrxI96tGdW/4mP2Jg+vxbnBzQrZ
52p4f+Ocyi2wiXKMiErz/fdagQmM/AQNx8Z9AuIZ/YNAeUl6TsM7x7fNUSSxCD1GblG/bZ0mfTrK
bnAoGIk0YszVaH4eZqAx9SeasUp0Ux1FMYClRjp/AyFqxWY2iqMfk5TanXn6rj36xiY3a/3kexg1
Tszl9deyd/NAlOsxvsQKvLEfzfxdCw6CcorU94NNpoEN3NUgavlLyEAF4sIkLUwHKkum1M4aorQl
AC6XaD8eWHC1YJdajh55E3oKaVAopdEpxq3qExe0rmV/yMwGQHoGSPfnmfCAHQ2tjRnB//LcjfEF
tLC48vAv1gn9yL/HRRjuDt+WUKstUU+QvSyH2XjbNhPSFk0OB+SheqSAdi5DvoQ1eCrbK48AL0Iu
3j1I2QjLy7UMiUKFoegyr82/bjR5Z6HuOS+8NC6rxunXWvLb9ytTgYKTthJYSsw9Ksjucea0nSzm
5O2LcG6WRRQpQKj8uzvzletD7bopPLC64gsi2A5vM8lEMJCT1A1uYBIDxHP1l6Ix6RTITZx8qfQE
n9tQNxifZwJTC+4RkXWbtF3tq/p4Xlg913yclHDELAYFE/izSyN2IQyZjOfOTNDfzj7IeppZZGrs
ryz+PwA2r6lReBGfCq3+Rs1D7V/+ezRcZnQAoAV/nCa0n8imsaqT6VWsgrZlOpngJ2cxOVdDV6iK
c4QKvNP0RvghpUi8/O31aBmX3LIhWkHZeXyxSi5JkHDPNvq7buz0c9LDgRbyB69DcC9IkzdYUwdD
oM5++CdScAz+dCo4/KVk6VCu8rjzTICVLwutM9bTIkH8WtsUy/MS7LCZ01oSpwYt/CAHdsQuHi6u
kx1XorPgNxvoi5i5t1fBU5c7+KV/ZfaBHj/OdbLTUUd2O6rm07u1a0dZbd0fodt4djX5LBV24gRb
D+D1CqQo2lXuKOZTuL5b5DJPB+uSsgp188crGyPtDOYZCki+0oddjEMZullkh/lCCghlJBPaAeHK
bCcveAhTDtohmo8lvtAjsPVCbMTq919gS0kDn8DPQd6pnzzPWQQX3Y5qVZ4qQGm9N6sfpD51bksR
MoHV8HBQm4Lp1w0lOMDqGkdsNaqkGbBlkmZvsbtyXbXlaezyqNjq60k0e/7s5GGOJxnavLQ//7Vf
+kVC8BzQM0gGtRBFKMUt7pO5qi4+4KVC1hJdyJHQUlLrYDlzV1nIp5yIOTffVF6mybcGWfiDWkDT
PhzY1Nr+uGIBzUmiOAJKRyS0KfGWQM1U+UsYNQ5+g1+NDDspvWbfYVbHaQnfXDwaZNIgZicyOGbs
4p/qnjP8fZY80/hAInNxXqRhyb19ruu30Kgk0iBgSm1l88F+ffpnEuAicVw8l6yaxpaQyQ0lFQnA
4ItPMMIdBW3UalQYyLLpjeuw/ZSAcpIofsQ0Dy5NjMU74QPWwJFW1JpuyMcDn61zEXB6HLdERo/Q
3JOvDXpDRaHwE/1xIFbVYFiv5OEM+Qdjb00W08FBnr0ZqKHlr2FyaYg7c6+unlu8ROaNBpFHeiNO
185fpDlVZyMJoJ2wVOLaZlv25nWwCNXPeuIEcgfykLedFJTFSieLLYSoayKUcsmMM4TNzvd7JkTf
XdYoTpSA8+rOmFkeNvuQw5CDyoUrdej4gsR4YBIdnmwOw0ymhItCuT8DINeG9Cs5ZxtZDN06Cn6P
XZ8d6wOOca79I4ZXL+JS5goRj23Udfb87MG1GPCDzeTxyI9N+BgiGh603MeMn57GJD2N9mEyPuuA
4V/+vYFLusESZebaZNP4ianj2Hayob7w6KuZlu7Qw5k1eAAoHMYDKZENWKKU/tFqlTttWbRccQM+
YpD4NlRhJB5EuC1EVsZGPZUP2M4nTwdal+zCwXD8IXBugAlYNriVXP7oISxOl5hPe5i1VgbPuYXA
7kQICKFOSaaHM0vtdWARiuXjRMc6YxDy60iJNf28RWaEHZE0T0s24ga+c+3VmHMki5oadfcrlHCX
Mutzxv7AVO3JCt5qZwcSTI7wDPmNPZ4B+RMBjzobSfVWhsPZzc+MhMbkmYF501CZwKaLRP41ETVM
NJYkkiKXSsu27bjK3qhDreH352Nlkr5uey7TDpCQw1/IL4gcpXDIdwOPTzUWvxML6o48Z/jzIQiO
qvyV/uryeUJQZHfC23SGZIT6ThXtzqjDpByFMyBv6KVKuOHze9nfKc9i1qEIH3GCof/RSXQAtCqj
Z6CyMgketp9buOhth3N454Gxjb41fHZkRT2w2KyzcJxjC9Agzl1lnLdZg6f4fIINdL5AO7fgAGte
gDXr6eSqgf5bBzX9IKjcnknNN4XPgfhySzsRXj+QsCzyiGSLGgHhXymOJWwl11WVjw0lHVy6+ww+
xlakK6vOHlKc7iptKJsI+BNLXM3/5jigkYuFRPMYrMEduVSkVXqjdiR/IlHg8XaxYTEkxjguJuca
yFqq5IehbkAcS5azrGXIW/f7aGYskuaCE5V8RGqGvqHNeCSQDhS3uYyt8RWmiPOcepZroJkQBSKD
yfX49oQy8VeeXz0MGR4tYi3KniRnZIrWdFGchrUi6d66Y5s1T6V9XAH/0pW0dmI8+nhcnldXu0Vq
eeezCYpueJUJlRoROnuQlRZmlFcd4dgILdQiohzkKWi1tdam7jsiEgLr+aodSs38i9npgsd3nvhv
5bI9bZ3YZPcH1F1VPRb05KMlraw/Qj4W0Allpra2lDsPpWWI1nbqnGo0jmMJJgvZqfvLNiBkTHlm
3JsZNKRbm46rz1o8YqesKjQqIJXnjBPRgR8wL7ZObPnHBxPm3ySo8zeS6Jeuoz8AX8GtHA5S/PNg
lWimTvBas8RLqmIf2H+zdqA+DskRhYih1pj2ce7SyUPwEKF/0S7ye/Iu843ZsdIub47n3fyP3CPZ
VyKx+Dcv9UvW18ibN8VrUnvOFCKpQSiq680QY0Wsmt+oGfyx1lX1rDgGMO0VMzEh2ZW4/UYaUP1c
EKzROd1zBT67bIAn6NdXmmpnsBelRIG6YZc0r1s8VSCv2Q1uSH08+FHcY4NA7Q5ByadZk8XLrIij
Us8Fm6OJAuWyzdnfsDFfuK08FEhRY60TwJ7q3D+euFnZ7MGO+F5Xejb8F9YQ6zWP5H4ool/oLMAS
lGYagn2Yje+L7ISLkFKJNH7mE7EpoqXmE5helLrIdzsSw9jcMlgBTPZHSnHexy5ybQvx9rgWs6sE
S6CJVaUPGh6K/hq2L9CeXq8qqIibiwh0J1fvgYJEOC9E5+4CCdn0LvsCwn/sLE0sXpWJIfhBpjNr
rdN5wnyNWjzqqx6+/H/yMM5njgosL95H3mtjmvar7O85/gu1NUzgcWuASemcElrNlBCmTOvt10u2
+n0ETu7wEpzJHgxPXhb94dWHtgr3TVO6eKgi4hBfr8sb/BgU3jvX0DzADRcW9KeleiGRzaIMqMIh
+U6SmoC4KFuLyWfPB8bFALslK9k/EzyN7vexUEwIKERn1/Heg+4JE4Rg+pWPUi0xJ2MFRAdYZlAk
1bmBwxIu1iIibKkGRpB/q0WmK4OjxVKdO3lWnr0UHN2h0STl+k27E8NdF0Cebx5qQqavrQ1gIhIm
g2qnZ46Ml7E7tgUYpNIFVCqABXT7L6kww+zsvULi3K2oelCVxpEUyZiCjxirBgu/OYv7ONnfbm6g
juk5wPXSx2HYHuhgZZLW0rIXp/r4F08Y+m0sIFhg5T5VbuxY9pqNcJwruwEekFpZBkTUa2hEd/C6
ghynmnABJpUNipWiEkS5YibQ+781cDNdT1l0adUXI8S+2Dxs9VjnLQAmlHs4iSJpk3nemazZ57EG
KeT+RFndnifeYAubqpwl5i+X6mD7mZSMWZtp9MuflAll0hTtAC6Ns8j+kG9Rris/eyCTtzeXTaYL
VS9VZ1zzyVA88NWa3TTax0uJHVb5Aoe4Oky5ZU7cYIfUG82fk8sA9D901ralQqbWHiJ1W135lTAY
jTxfZdQWECVeSv3Nyrsy7CuRHTkulc4llMpZiedIA7LLFk0+L94aPJRHFuzzqpfmIaY0RB4mfJp2
ljSVEePEbjhsryxN+jGoYJSuzf6XFJMOe9uW2yEdFOBlgcRMLdLugShntdea1pccM7N0P1I8x2sm
IUl9Kvkvc41Ej95i0881z47smPPkXxqAf2oZikpKZqgjBjcoAM1qgQlbKK/Mnt2VKJykWWofKeLP
ZqaTwSrkIS154WQa+Mox0GpE7bVrTfxvwNFcXT9ThHBzVS1Zqz2hhgz92+wr+sxbjiO64Mlkk0Uw
f43qyxt+8KHqmwG+97z8JCTpCfxqOIxNB4i9RW4gaEENUoe8HXyr49HQJCHsTznc585BJx1zz7R3
Rc+kXqHqgZCFy+YikVvmQOpbDJ2vArvmvI3tW7cNsLFyIeggrSoM1Ch0TsxMf85D2yvtFal+RkPd
re52wnd8NQGsgpptm6jI16LSMwN8c9CoRv8rE5keZ27T4biQCskdUjsFU76fePb8NrW2XESnssnb
dMdw1GDEnkTlR2EVv3zJA81BW9T8pvCwMtDQiEigsJNbRiUNcz9xJYb47PF6p9nqVLggy4OYW2Dz
mMbUM10P4kOV6t+w5OzTqai8s1kuuvNB02hnbakLV16HcllI7KAtEKAGNYlwUux1tZsw+9wrhguE
0yhk5i9CVyN9NcQmpddrwUzzzZGf9a4GUrkPRtfRmfU9UBP3EefWUIRkGeXMi/UK6pZ1ObwI8K01
wR5eunE9aeTyLAsnjYu5dRFFHZkHF3cfNw/PqWwA1dV37VqpK69a8GmekHLh2F8x1OfELyHW0h/m
0L5tcDUV/jEXPgPRm5n7RLMyXgEkDy6XnLImrCWaUqSfc5ta55po4i8VNH9CqSZ605cGCT2hU3UQ
1KFMFURitQReRnfeGY4s1UNw/0o+Dvq+QwKf8DR5g5QH71kyZinus8PZ3feVDZn59VtmkW6xCfyk
nH8FEOwGsan6ZYzbpWpAV3guqeAJ1iD/nQzPNMppU+d8M6rF/iD7D3oAefZT7Xh93TA6k9TEZWq0
wPCjr1AOoN2itBF0KmAffuR/wQzuOlG62nTNhcsh5VJc+JcyZzvRs7zBg44oUNfLJjP10rsLFK95
p45ZbdCP2TLe8/m8tIJ9ag0xx6/EeWUQJbMmxz+mu26qHF8RFWtEcQ0NAO3QHwPf/JUBmnh9TMSZ
G6SM46HxDNoUezWcbtOA1VYPFs5ahjOTy+S+sHvAGvCQknLPfTl6P9h0nYJ3k21t66Te1GbJfhOD
I2/b6jKxJ85XIZpSNMrmbEDdMOV1/wg/94AjuLSNLq5fMg4I9PK1tsIqeNTgzOQ6Zt8NuiGD3lEl
HljpA3CIp/XiCLPeGteieHMjlGLi43be6jmf2vekfU53NFXZ4/1UmnrF84P9mnqRoMLezk8vuFdW
qmxGovuicuYVjBZD6LTZ5VA9qRW8NqmgQfVEu76AxSkAdSBcWYrbmV6izo8R7FCybHiOb1I8W072
K5M3KqYiuzOw5hoCrWGMG4i2ojPCcaDcrVu8x8XKc9kLdWa8E6VM7o4tLOS4/O8VVUBVwOlS//Oz
U6pJuSiuNw/dSVl5X0FHAwtkLMo93sJi455xPPLitFQ6ACiwiFXPo3PhYkiTjwoI7gm9RwmGR1CZ
Hw3hEVfbyvBjrvkmKEeEDCaanPITeboA5DG+Qoiju37Dc+x4M9ZJkDDRqeFwzY1sf/46KQ3YqqC7
ofxAUt1S4wmJpLtInS/ut9WFAlVvzHHDAFRk3OBsLnU3TglWa8/sQW/ChmikO4kJBQk97PqghGQg
8eOik1okQH9+aRIzXjNpLpPBKR/lOsEW67w3EOxsLSUMss2NVCoR7gVqZZgrK/iOFJJzJBZhDpqT
HO1RZ3XTTFjvI/aK56Rk87xT9d6gYEZ8fDa1RdmxQ8BzToP4IzQ+0tMjV/HmRgnSEn5EVH7MNd3J
w8owLrQHwX92ZqbkQ+ecW9GhfvHEmLs3o6Pp3dwV8xDlvtAMpr4XOCZRb8GUHKB2A0DQWtptuBa5
KrQ++/ZZe3phV+7tafBLPms1D2b9xYo85sADSlVw/8neU3sNYOqF3vfDpp1V7OE6Yucv/tSTZB+3
lONGvuzR+HSU937e0lglg0WUhRX/NnvzZVVIoTFVWbcH+DYXkYWu+0m988XhhT1BEUky8ouX3P9p
ATzaHA3+6oqLCF+Ts6KADsmYgGPf2ML1QBt+F9WXZ9V993t9pxfaV0BtipIP9ZQVxYImHu8x3mla
zHFKC7SAIr/gh+ewVuJk+XtXvlxexMY3bRReYKj98ROQqm5yWfMpaYNfg1Am5n5AOoHjpSZcgiEi
QvXNu2XqwKQGyBtmgEV4v2HMzLgGA0nbyAQ7uTzoPT/o3mHJaydBMz59ixOansZ3p273V8DQgbgD
WWtGKrFAa473aTVsOySxaeexxfPFOp8Ow2ezEo3elUi2AlYbzf2x12ajP4tthusAuVJnJueIDBht
zsAqwVycDz15ryx7Lm5Kx06Era3qM2XvrlrVhTvywRPD+q2h+q56Yc83955pmvdywKzbte17Xv72
hUHdkV3X1tKr38n/hJo7qr620JuM4ntxYqEju7N2PL1i4cpr7jYSo99zV4QASEWSIJQF3TPbhU/2
UVl6NJrZik5x4mhVCpBSSo4PexqeijYQVRzUO8MGqyW/4i5pHlapLh+JMq9+uYZFpHEPrvRJNcY0
lqG/mtOeCtI45KZnitidUTPen5DWXefs2XyGaYon4U0sMLAyls6qONyI9/LBW5XErn8GeGwPY6s0
JrUeZ71jVY7BGGtF7tTCEnzEl8YDBMtsonh1yuRJbdvKDzgN1c24fGFZpIydh8sfZK0zsfIpnceU
D+0q5SO2q74PBw73iQBSSt97u517Z1ErlFqjntvTO01H4s8MKvO1ZdqlopG24Ih1DZ8jYvO4oSNE
AOJp2jeAtaKWrqG2v9kka61vLLvq5X+KfTz2PP2bZwdxhCj3oGus9WxoU3HzXlLT7KQBu2TVGdO8
3CdvYSR7Dp4D4n56dWpZlBKioPpV2EjCH5QT7eaoPCDwkmeDkeSRsaomcJIbi3hcVelunLEhRn0v
ISCsD4jFX35ykqMUd+TCND81ljiifT0+0uQ3/43w2sFQs9Sw/pn2LbZGyXik0VCA3xCg+lV7iTba
gkrH2MUg2O6Tb41VOxWC77AyloKgSXXO56q2qBEeCv2dnZEKsOoVkIXAS89XfYVSkrVHxCkGPNCw
DuMgxRPXXE0fV2ARz1r2X2Ya7N07BO31hQGahnLQDkVau7WENQkvg7OImmJYqwOZlLxhPtAVaG01
npQCR7eOHtepNI9z2ijPqoxlV45i5u7ES171nlraj6lCj6Mav6gLoABE3Qsl7VBP4fi0GIJR6fGr
eZt+qvdDqSl/TZWVowoKYPRMrD/3OD74aqJCAfQlrs1Ros8RSBCAr2o6oBO4RSY2ZBk/3t1emqHA
DRU2Llt5VWGBFy5v8n2qX4U603zPwom59ZBqqfQ3GucJ1YtKQt9DVosD65MP+vydF7YGC1g0hMlj
nbWP3Iy5Cr52aojnMLrln51hJAJ8BZwuQY2/O6hyGe8zkxfY4112nG4yUU4W8L37esidUaT4TAnb
tFccwJuHRV71zHg+RQyAKE6duuvZHWhmHwaVko8J4WVQqvYMAWrI3X6b8mFIxPmhUPa2Ms5613Eq
kz+lEqUYkgqrsGppweS5dtBezb2ORs/Pijrk9nbdIxKa4jIjCOzWegj0wU/mCL9YvJG7VrlkHZNm
u6jN8u6+ZGe4GFXrEoNwDwTecIdt83f8xLbjrZdkd3GkdUdErBZkhkuH0FlT+yL1Wp/VecYbQAFO
bLD1O82cS/QEv+4kJT7ywHKGsOM28XMKq2k8pUBytsiECk9vO1K71ywQ2ue9o4lB00Rajr+F+jS6
gDiOYaGMgXTDH81Iew19Xl3nFhIao5LY9Y/gVDjTMdSVXGyDNRLH0iLLthqYum5LYKBuAWCtM9Sr
2ea+KxGvDmtzdtl3zGbloZMuUUcRpv+/PutjDiHnBeeOdjsiwU9wASQLbBVyIUP/azS8oJJAEvb7
tiD1LVIz5dSHUQIdHTEIM1Ih4ugWqxa/r5TfXQbvYncaJ5FlubghC4yEEy9y5Y17RaicotAGr8Cm
5LXjSbPORxOVk0xEpztAH8zP8rFWMwuMrX7PtRdLil4D8sw9zPyOUDomw4obGppX6Rc8aXdwq/ct
2gXJvbSbvlB0xNGNvfiL7CNelCOmNkJmz6h5l+vKDO3t6j1n+WW7wCKXs5xd/L0yNHfB/u3GTCws
Wuuo4vSYNKI7CFY+RbHUYM2U2zXyG83PtUoFxWfg2E+unHsu5lQZ9Rwkly05PFP8Uz4SO7EVv0L+
4fglLjqf86M0vpBc7rHoZjx4of9gEkf9D/Xyf7kL2r1cFiKpImd62VqxucuJK36vi+gGZyps9tXe
K1xdzTjN+24CcT28Y3Dq4FJKpo6zaPdbmuM6uYGh/ea2Cn5iXAIOykvhe8TGN1NrbejVFfBPP1BT
50bNwWtTpeji+Hk+cDUSOZuU3zlplsvGRnKzyMNfO9al5ep8V61xn3vvWokVgK4ds1RTVO+H5Z6I
AhzT9X03No4GuvV1bu+drFs0rULYuiS0nuO5OHMNiynraHG32NmsM7tMqEauV5lJht3tjCkjC7qZ
Txqn8c/0xzN4PrgYNX8DCua/Fbk2mH6YspO3YrqfRBCmpvhYvR2ctBNaWjWr/tTd8C72Ab5+dH3E
rHeeWszsPGzl0EvC8qS4HfHdCi5p8GT0Yk5ztlZ/J1M0/P48SlPLgm69XOTgd1s4kJuJbsx2MqI5
6grT9Z0OkVyuXvp/owUZ4Pd2mOIA0cdp/PMCTyLMzAxdydtgAdkBjGXeChzBe9K6Nc6vBYcg7qBU
EjO4F2zkv7pSYBbkMwwOndkXXu0BjWQvFqOwxhteTh+FmvbiKc0WdVt/hG/hDYqChuOIduu+ZJ0V
3cl7OA+mzcP2q2ezEV6XxU5Fnti0TyKHbzThnUrFKCFcTIAjvkgafH70ypRxgxUy32OzNH62pbX5
zlAFLN2Zgu1+iy1ma5Vts0KWdKjUBdiesAl4osNHnMfWbiKs6Uq0oLmI5dtqV5o9UH3yvOaWWuh+
IiwTj8s8fx2pMVAg8RHDogmsWfW1kHFvXR+3URqPEos2LesvQ8yKL4Bje81s275l4pZoFqeihbYD
iJqF2W503BRcxqLk+nn6JvuCfRcxCDgYykTyMdQBA7SMocIG7vxDMj0jP62P1Egw2YSckzGRJ69u
CVo+YeNx4rFvI5Ng7vMIO80TfwAiphDw/QHWNkbKrfHX1SIwi3Emb/VlRLU85BpKUAc+uCGBBKb3
MIh88nEgPC2cm2wS7vIhYbk8X+01lEq9d58lJAXiNJwjapxAzj9fhGkkj0iNvLh48CVeI2XDTzCR
E6qM0+DW37PEdQYpZW6P5+bbJQBjJaI0M6iZZqb0z0cnBBIPC86XXM3l4RrAlLTnkF2vgdS9a4Ms
fITFZb4gLdHhak6wA7Y0jvQ3+P+rdb+PgWspwIUtmhAEyqUoV2KEh3DFtALGx0CL3QElI8p+zgAC
RtCuw9nJ4NSoH5VO2Lg5WYSt/2wiHUQ3rjToYFxiVbott02i++cjcgjUtJBfI5KumOUqYH9hVovn
V2I3KwQvpdaQFzpkIV+q1oCo+UmmJCO6AtSqNZVx6QPMwW2x3wwlZtsZPThh6OfSSvYDEY7oc5Uv
MZBT8Xz4RAJDF51+Xy6skbUW4hht9U2uyAsFA3V+rHoIspysJChfvuUO4+1ffgfUzPPVJKRksLeg
GI38GzYPG6Sjwz9fenxC+9r9oUm3Y0K6MjO4BkXwVXkAg2ISZQ3DNOS0OiC8QwMw2S58fRFnYhKh
dXlpx6lIVgwbrWzbODwEB8cruIf6FpT9XR/eqabLawzfSNw3vHPzHyvwERYd7WhUbpflMSNoVh1O
TPsUsHHzxLcFx4MLNVXO8Rx0xwCc5vNqluMYn+RYfyBnfPeRmN22I2J1aKtxU+w3wIJwru2haOYX
XvnQfmixgdN598f6t34YYy49Vuh4cGAevIbN8j7a62i1bDm4QlIoBWlqFkd+KTXiUiKK2Rn/Td8q
FklElTZS/u8P+zbYXYiWTuPMajsEJbgqh4Dm6itUd1kcj2xoXK2LaoBltlxZVTzpLjzmV9xCRuwa
OvMrKyG4kzywgn4720Zsjdi+Z7t6e8JBRBXCgokOE6+TDXKpEfm0jxZFOprMmjzZnHk+Wh3pdGA2
ZUFY951SC7DGAY0tmWbSPFxvLBEavir/OjO5apzhMX2IP0buuzp1GeQONiOVdESFYnUQk7Xelgdv
wEx/RNTlRoNl/jI4h6U8reG/TYy7UZx0YDNLzsE++G1djk+H2A1/lvvPVmS0txlp8r5J3mcLPwcv
pMZ1m3rcZFLd3irLf/62PF3iPKvRJghpaV5Qzugj7oqnEKu5qtY2QD/WlulAldijXc/52bqPgU3K
tpHHYyn9T+wlfNuvPDMs3U2dGd5ScgYfBhofNSuuRfJcCH5fbsCk/LmKJAS2o1uSI8KidkVxG7No
aqHt+jHv4GBCEwFVkffXcBJFozAzqAJdUKKs/RCUK8kDXuk5AKcUo/MUZkeJ7eOv78U1H6MPV7Z3
shVkiS0DZh+F3QW69aGcnEVK0cBMfdiyappQ4xnUG4hCpeRGM7IavGdgYj4UNuulhPouj25X//SP
tjjG3wknzlnE9ftHcUuBAqz6BE0BrM04nplt7JV9IpTLG8ckul64L+mOjUfm+wd8Q+h1La2C1BYb
mAiYLVkfR4R7ByG0s9JWorrPjgogJ4hWd3zMBHO6QPxwPb6S65JQYIqY2IMgQPzyQjb1Zu+v93nK
y0N0LW+U97pDyipFOMRtsVz4YJFGWuX99BGO98oLKNu68klsvGWkg0BKbfuk7hLZ2siAHx4+0avz
8CVWEAlQBQn7Bgr/dvYkbyDl444zOYhV2lgILlNB5XBTABDkPMDvhYCzC6mcImEJAgDsy+po/zef
zjk59mwT1COEGUqnt7tyTl7IH+Ux97/jP6LvAL+KOOYyRWodyV3REh6wb07oF9MhOkkwnnhC/M+g
xjHqNz/5bPAeK+C5ikxA/Lo1LVTqK+LYHhoXufqWZ9SDrl76G6jq2fBQqeGtst8uHVAduDFvNTKt
3NO5vIOiFYf2HB9R9ORulg26z03p/hWk4SVL/N0tpqgw0RB4AbtIpaq18tMt3BF1pf10EGFgiMhB
47M8C9F4fNKsMDUYJoGIri9eeS83ZxAQVf8Pb3bwKIKpcdvKfU5nL16g1sQsyldn3IVQgNdUVISm
3roFZk+J4Z6KT2pLkThG5o2sC5wf3TPan52xEfvdARX5dZYa4iDd3sGrC/lJ7eDu8csYcB+z2iHY
7OsTJ8JxqD8lTxEF+L6V47wRkQuwgpDwCfn53bRTqyGBPFpZesGu2rVJTrOvIAZXAwdv2ZXKRGw+
sCYu+SdyWvajwuu+ZHLBgZVTBbVRM23kq+0Jk6U0x8ppK83tSOHPlorWtvpqir5RG/UCpompQfCT
I+TETequl86V+/GredWbXDgYUTzF7UK/miCLgXvAHlvnB3vTpNiDJsXmu5XnMal+3v1LUaTax6t6
+UEed9yHmqKmMETON7OVnvtd6ipcO+VylPgfCUZNwG9FOTVTlyEdkQyHX9Ar/s9RsXyDF9C5gGzM
S0cAsf+wT9TgRUDSDcuhKVP4HxjEh2I600pJmVjsRwOZjkwcDBseN5M65lbW9AJtFJ0BSDeTCGWa
IYXPUYI4ztJ8a5MH7xOG4Ely4Zl5k5uRVxQEO5RPBSCcJKd4vCfKkBr0xdW1KuoY3WJIodq7P4S2
HPOUpXKYRgWVUxIa3GzXtWKuLpx8BQZP3v/MqjrxMyOuHymLPkU7YYx/sS3b3xl1t6R5U/G1Qx5r
oLnEjSLN5bEtKClgd4gLkkzJEhq2BPT0RblIU+vR75aciKcgCG75XVcToI+oHvPxMwr/xmeEIYNn
bo5GTWyEnBOUIlViC/CPb2IK89/v6ARg1Gt2Lz5qhx0Ia12sy8YVuXShwtA+Voe06lqDhDcxFXBE
TW02FFC4GiP3thGBqKIErqmOMNaCZt7PdddrSuGUifn3PzW9wVt6RZkyQewvYWP+E9wGcEygY5Vk
iDiDv8f4XByVmdOaRHsS4kuhFiKaLMxfEAeaMx/W4GRxRF5dDSFxxE5IbhVwdnDORb2/zIZ37NXn
nBu5GmWqrNfVN1nLrSvcB9wfFAkulC5/P1IE8qblcYaOnWJSb1CEoTZG2+tilr78FSEGwy1YjOGe
ANu5FjF+/OO3WsuwAJABTxuMraSGGs9V0QjD6fSHkKMH1uuigwvQsvTZooCf1UdSYxI+huGfSVn1
G4kiJxyGWvsjoHZ3NJXiu8/2xYu8T8NYPhXpXqlMz624bTcom7TK8w/2xJgxuw4ad3JFmGOdgVit
TPP8zGKAidC8d99coAYaRcCbRSguPa5/ZtqrdwlydtaaM4OWLLBV1xCqXk/ThRQaBj+YHIQQOWTw
q4g9sO4xV+F8PJH1fTNdWicWhUeyG99S6utb8s4rR1I/8Zq1MCAjqcA5gxNqYmdMxgg8B/lpqBEt
5S5FuBLUK5j5IWijyiAnj20txav9JZdyj0n6iytsyNVuViUUmrXWm0AfAsymGIc0QDHCJvFAHIvj
95rxnjCFGJc8s7Ss7Rdh7Tw1FuFyhaqqvDXNgDBe3WwFw2rqQeRX072CFFVt143cPS90iNoyHGlD
+6mNn7Kz3EdljscOtnIYMd3g7u11poIw3hAYJ7qPovIPJvzYRLDgv69V6e3E3iDA5nYbQGj1hK23
MyOSihsF/OJEzIEGq9yJQdFVwclGH9oGeHUQMksjWlpYOu4UWOebx+S3okhwvgUA0rYxGLACF52v
066HhLjgRTc8AuXchXvhtMhlgEdRUrLK2c1+eLQT+lqZ24R8S61tGNZByrtXfBDoJUU3mrGnb2p5
e/N7chNC4N8PgkRoHhFR8qlJ3xSXaE/BL6MM9PikOHS94BtRNjmVJLA2/9S6mnqbSpQF66P2aTDw
Uwgwh46b3lbytD2ChZW8c0g2Myt5xCRH1EM0oalNad2M0BISpPASNkjY4tfgxbw3+Uyu9MltyGT4
N7QSMIH1jH539M98u28F0zTnmfs+o/49gnTU+VZWCBM1W6Qdyz/EzAPa209pZJ1DgYglF4gSxDb2
a+H9SuaqJ0wS3rbPYW+2AnY6OqNeWHKQS5M0BZNq6jI49BSSEBhiIsjtTvXzFs+aE4qN1Fw+xgGj
MGH0KaQwDLfj0Qq/iVUckc/HtnjGoHVvh/rb7vhYKkLEQ2ILYkKNtNnzOOv3/ysmeFBJJBHoqzeF
2q/8hIwhgEnu15Q6sVJ5NxKxXas/mVCIdKRBPCLnkqg7JfYnxzEsk8Cd0v7nOWMlhv9Zn6vLBpB+
XCUR5ha1GyCqQy0nQe6X+NP8uWeYc2ccIHZM0J2MeS/Za4/NeeG3I9qbeYjs+2MKtyI8jOGdf0aB
HpfaF15RMst4tQ+5LTSirf/BCQhP89qScjFbe1A615MzTtUQq4omZLPX1nJKoKR2L6/CziQewzIT
dzMT6KauZVeJJhxfAOw0FQ+E2ywVuJfCUZDlTrEANviPKhUv08UU2tf/nAwqtl2pOOK9E3N9QgZr
4wG6O+hRyEkdg82B+5ZckwBBcLUHxeURDFEnT79py5aOmH+9rOc0cSyUbmWJ/ZKC20heXYwDXcuE
oUFvQXjLA48GfI2EkmnAlzufmvBUu4h63KTz8N6dKd2VTpAHFD9KokzhmpgGj/876iWWrRtqFU+J
QkhqYFEulQIL7+LBDYZk85HJACA5/JUzU2lQzf598ZwjtLKJEmXa9kBFtihI0ZEbw+AOQEtx3Baq
YQXRCzPC0xes5QgAmb42JdpT/CX21ewpucKBSKok3QPL2Yb7nedkH+WzvwvhdPm9n/HKMxUtGa+J
8d8xMr5tcrCMsbumfNGIdiWEb+biNsILS0yAzwcmZfZkGmgYdEQRdZBkZyub0ptdrvLKWk5Y/uZ5
l5QvzR8maef9W6VArDqNjmh4v2DwkD7ZX+d1fCG+bHjnA8E+l0YQaMkSfUILmYmoCqKbUtIQCooI
c8S4EyWm/tQipvfAOc/LmWNbPwqXm8o8I4Ks3Cwc93b9za43Ghp2LhXUW+QG1+VtPbQCfXsBIEO5
LEdZ5L9W9AkkR7kk0bJy68w+DAQzcCO4lb6WFkFYcjjKyOGTbqTh85wn85SKaMbPdRJgbmForkbY
NeH0tZF9JeG/OB/wlJrYWszDDrfJ6ex2yoG/PtbcV7A4XPcqUi7OCINjXzd92l3gf9qhTeBmgBL2
12VSACHERPhsrECYUbkO1VyVVikeGFH3ByGQnyxT+rhQjcfH9fwJQo/PlvynIdiGP9wUeostrIxV
z0er3+BElQ5XVTbG4QiADtUaQzyxbt2gt9TfcJ6V3T6jEmhtOcSkA2dremXR8WzdBBNfAefHVHwJ
oBQVYGNDNwfAqNikxGKll8NAsNGlUTzZrWfIwBFePGMYUrpOOXd1vIv6WwR3RCULUCdhejZvYIZY
Dea94PmdJCRdBANOWwWrM7oFbMfAxVImfknaSnSiJcQv+TtPtgAvCESfskrZFpEJRfkyAbCsagQR
3oKsBoSGohZxJLr1a5wXpBJPADWqdyLvscskMIuAfHLjYXDOhZt7nwoKbl581Y8S3xzosAX7O1Qk
Y3uSBstHnNM4k/MJgzuKf9djZiKwunqMOtC5wEXFcSQ9J6cZbixrEQaqyqh7Z+3AUtEtIB2o+Uhv
2pTe1cEMJuGvOFytOAkOvtN1oF2+Hrz/rRHFHwD1IoZ4qrpk7/yEDT0aAXvCi+xi4kCLRE2+x/K3
ICHWWm1GnF9XiuYLoUn8AWoxjCGBMst0H/+EQzcKIic/on5TRId/KE7xvFXDOMhY3os+hizTfDLR
ESj+FTub/P/Vu6oUmipnl7MQNzsWKu898wByV1uFkMd3d2v55nqqkFKeMHVDJRgO8K+gaC4LyAFt
2Qf+i29oGTk8lVUEqXQ7NoyiV+0oCEawY09iblbdzv5FJ1rFsSrJWDLMZMva9z9VJq6vQjwySutu
rMlLPBEzVK0lyPDil23LFUW15vdhK14d5dsNmcpwxZsEAdi/2gIKH3MvE32UzV2cd5q0fefOyfT/
expGgt9EP04FOA2SuASIxLth+leLadft+9WgO+5ebPbUec92/9DqYW4HkJKBNvscfYHWxDlL09e3
d8YtP5HO249hxN1QiStU4SBpGYVnIzbcRgWT3EPIanMjDVBdfzAu7miF8ybEA2DRn0U1R8DsFI6k
R85PpcZ/EhlJxZNiJsQgd1B80Rp5Vf/URc4CK4rWUei9WopJTEl5vjnk6LGjzK9ogu2e3rlfbpxN
dDPkTexSSXWdV3R1qJ3El5/uLMnPBqaNi3uwA9KtMXrR0/JwgIULpmw3u4ALoDMxbqtgn6dtl468
JRGVpg5E3arcPqIPKg1tTIEUzuD1XxTn0gGBugU9gvjLIZTGppSwSRxXDjarx93XBg+k7vypGoXw
VLsKtRIy+7EPDkildN0xQw1Y7L5ySYQxobCwCEOzbQUF1CVp6OKlo3oODsc9sDFBKYnq/VcJAh6y
8cmAElhupZAoGsJLH9MWqVYjewY9UUbgiRsIUPCeoMq6DHR+ULDKY6WHjCZKh+WcoOIV57Asy/jN
1AlvimGFhYmuVNV9Fj9gv4M6C07m79iy1c8TZQ1oknYlz5wUUdKv6C4NJZFV0iL9JqmHzlBphgMV
wGh+4PXzzpP6XNG8gKFdfP7CQNPSZ2/faCRVkO0jzPlaV25nTGnAFOX41sbK4t0w+f3H29nXYhlC
CbJIYd+LOGv5Zkkt9i/eSSNTXKUEZ4mFDT+C978mfa7YmAPTJxvJmWBsoLUHDVAQn58gbL77ULpN
H8+l/W+YWGGvPnJLahZswbZtw2ITccvvADiMEHrUK+ptGM0O114oov6cu6+f/lEG1mJe0461duh3
rSWmEv86zF8H0WCof3Wh+qMx//dKrITuQYA8unIH0lA2xM7pgj4pOS4PO428yFfrZ2J7xQfxgJDJ
vH/gvWyRFNhKmp99K4dI5aJpFoi7ndVvuN8eK1K/BvkKY6MJRS6OSVfHDYSkAnMG8bmvW2gQk92J
FpuUFNDVTgGo020I3R0KYpZmMDv+1KnreotDqs7vxHotSNf0iEUkXPfqV+lR6BvNOF+I9pe1Y7VT
ikSUdmUBAh3kh/0aAz6WS/4UsQ8P3SeN8NHsKFBsSnXoeCwu5XR5TWP8OzFJIQhr4Vvwue1s3RRa
MrHefrERqNoRApG1YMGuv/Uj3K3i8mpwhC+D4hbVT7vtPcZrT5zeKTly15JcDu+SQgM6MfiGvJwN
8nsdCk5acXvuIiyZiaXmclwLNWq3ye8Zrv9DyukCJxrfETLXxjiZURm/rfpzkHMCyrtSSYGYzLsu
QOouJSIYSQ7WRMsAHkqQ2r4vuqsOVWubGc2GlaLqQqkeAQ9VlLyBhS9kA/L0FzeWbYOfDtzHMYfX
IBsRmwfZrfPeJNccJ6VdpVUBaRWI7lc1nrj1OZDtOtpl/Qj+LqKcgsY7uoYHuQUvP+ncyum7ktVI
Z0ZKOsi8iwJyEbwg6buUHEZohQIaAMoC//zXgL2B2w72e0EDJOLU8JuG9Qpbgbj+52TAax8P1lU7
3dLJf/CLhVygnrALfTWU68aa9UzkTA7nPl8tO0Gfo5sA8whv6IKbbPf35jPnKJVnFUWOkiJvDVZW
cDXeQX95Iqw/APyPtNxSdLZNLguNq6bZosG5VSByXdytCpui7sxEoJU+Atze0C3RiPicOp0VkdUu
SSboG+ZAVb74u7ky6tKOK0AEWQapOXvSTv9E/CuQTLl0pWP7QTlPIIvGpjfUClemL71YogPxDGdz
+G6W+SeNpa6hn1GSnO7MGH+o92zbJgruRzrQwKDUpA4yN4Msu2F/6I+sdhGFy78apKpsExXSZ2uE
+RCN83Q6v02kfqAz3wAGObP4dMlMra8eW9/Xu9ld36Avoo8AcurfNT6ZTM5XG5o72ifAFO6BORnU
kUiWCF+zb605pPEEpuP4vDGhhSAmLLd0braZNpcoDJ1IWhJVEiHiFtUbEYhGy9NyDLkhjgBxLOt5
V8TyTB0i1Rmnzs/q97kD7eKRo99xNP9F34Ae+7xv3/rPsElsHSGC6FDfqyovmwuDINw4RCWOWRmQ
GdkyykwlKkOMahRzmOyNGQ5UYb31bysEhlyTsqD2xA2kHnD+Z+X1aYQqPyl1quLalEIIaHksBVTv
2SKJ2H5CUuFpTbyFob/eBWQaIcXwfCY2uZ8ytLqHHwp6Qbb9+4DR5JE6vGsQTLlVL/DjnPQEA9hw
Hd5CO9mrVfXUwObZ/G8/zJiM47m1gx/o33cejl7h+udx4TC5oVhQXMP6S+QLszaZkPZhtHxhLhsq
VOR5ni2C/NYemlnQ6GsYFTmRZvrq3ioi4XU/uWDQ3Qg0IeO+hNj+Mr6Tn0d67Y+d2TwGwsw8dLR3
r8ga7pFt6Oi5pjSgnXEIEhjIVPH7Ta0DVuouzoL6SC9sU2/3Q8jKh2/puQ5uu68B0iX4zE8cIp/y
g5/wAdiS//Ep03F5hcnDhm+hic9m0gV8+AM5KZpHOTqPTeAT2A/IR8/R3+i/24wbVq+ZboGIyjLf
t2fu8BjAcnfWmddLGsa8s9pvXIDApwSKNa1fn3y6oVGu5fYELr6toCbJWytmtuAB7hkWBd8hNLvI
ZWd940Ys7a2PgZRT4PeEgNEHJAXJ/oktg4Tvk57/gUkuNT+CmY7wtt4aEpFWqpr/LmwJeZE85BOt
x16RCihaytbM+ZsE1LV3Th5qCM7eT6oIe3H+cqCFVDbSebZDGpZWScv2sFPssg2bDZ7hcGWbwJ4t
NjoOqWMmKeC5U9r/IXToQo+zPeynTYUAbu+yZpNf7jEPDTZochYeMbZBkVxogqcG6ez4gL4CLg+H
awKSHGAN9Vxgjmy+UhJCX5tjxRfKjI9LkS0y67ByjfI9RnxOrO6kuc0L8ugN1r066ArYFKgVK4xG
mn9Z9hDftnOgDh3ubrp2sJkl4xOr+Kr4HXEhS+4/jQfZkpWfY2I8bTytPz+lCTiHet7dmN4Bze9F
ekWvwdr9KjaDtHwOnNvRUcE9QgjQbALsCRae5MlfdYmk8HqLMHd36imhUBHmL+QzLNbseNitdSrE
S9Es0anCN7q7efsBZBnUVMaOI5QsJAySwTHkwtEuvzJXJ0sv8ssefQoPZyKIkPXeywwrddXIxitk
hn79MxVRt+Uwvq7gmuxVGTIaJ9emarRrgyE/unRPk0PousZD0/r8zFnQxSLZBKaq6W1fPURa0jTQ
E0Cl01hQcJhgjTLMRXCIiVPXNncT69ip2WV4A5Se0jeHi4YmGFMPmFe3fpVNHyOPpeWDOVtpzVSf
I3BKnp4dTB+TpaJfPOTfTIamYyQ2j+nqMLVBMCF16gKaSXVAfFCHst3ZjMJ1iJjXQrCCF0eBk+vq
kryc5QTDl28K3Kzf0hxIQfre+WmNd8R4HnUNARoJsrIxaA7v7x+2jCJ5TAumbYcLR+yqE+fORPbw
5iyUYNzyCOz8ci8/PdfAJ9yAhh4SJdhf0qnWgDJ1vVbq+ha2B8VkkqO6xVhydieioWdqPiebg59J
Ig8OrwxdUtvQN/Ed8K733z7jPDv5Tyo0mJw4v+pSP/NTl61/ZDpThNNpLnqW98UBv5jIBPxIS41a
mAGsy8MTsdkK0X1hjmWmTCmGw8TB3t41bRh/cxkac6rCgR9pNgMnZfNhh1voUaZjj0hnh83nHEZc
ZHlsL3GcZw+b5zVmdRyEDWf/TrPG+qOH6+3+4UzC60yLOfedjAQt7im2il/NziQfoxzQIa6VqH6D
dcWZPsC+JtVY9tl3AcVpK8i0MqLrUmTRqhcSi6/839DipISLKOL+rcJJC2xjn6xgYSsU9Kl8iXCj
4jHB1QXa2G0KncL5KFcHcLuBTChr6ykVzvT60QmAYaFlhaSsZzE/5avDibhAIn31iM+kdvqxrn/y
P+ZveOzRErjt/iMXTPpsH8BmY/+ndtP3fzaLEflhfBkSVBZ8GFeUgT1H0KPtwreI9GUTMzMOo4bX
LMJ13bzljWvcc0MQ+ZqhULVo/Rl876bYePMkuzKMWE6yAChMhE+MVyQ+XaUhqJQh0xrOyualWDge
a5yFoWpJjUToyZJdgwErB0sUYmLpXCJVeu/0nQ7R8wFDIOHhwuf7sif18eAPrTotvKA6FRpqbPSV
M7SrZKzO8q/6KJtrhyDHOZaELrMSfrtEcA49x+xUAxNgNq9AqArJ1EFu7driAEaG2Yq6kQy4jE0u
8pKgwj8ZbAvmEph3upeerlbLE0bcGWJRv263dgrZuR6diatwC1+LzDEbePNYf/Dp+mRi9aiQfY1y
BbwWBtiZMyY9fR8sE1Tax9yUAy7VQMsXoIxw/mBORi6kcTfOjcH16MJr0Cao2fMKkgHHHAfeWVc+
NPJr/C+vb/Hof7cCGjVybdEMnnYJmRL957YcyfToP4GoVp8vHS/lH6LFR8Ew96rU6PC9Ns1dC0wN
+bpzlQTl20jwUzxXxLnba4pNxSM8xF+BZwGRue87u+LU4s0dViXNN93/nesCbOoaeQIdEhnehR+r
xE48RdZozFRPYmBSLTfo8NxugArCb0aXm3pcrm6c5NuhZZhoVSrlrXYvXPsdGuuvQFsSBxqpCEVo
kkyJUSQ+qYSm3WkDI3KSIoIG5nfM9wOkBPSwMZzk7ZIhM0o28UWQ+y6vAINyZ5mjdzRH+aEenCaY
spmmUyxNr7bh/N9CR4Co8cAwR3fzqkEHi7+Bp7sG+xImspEpConvmcTCUYuneha/R4wIxhKx3IQn
OPCRr/oHzpDF1RA6Gut5w2kcuhBwKBMSche3wHUy6zlPZKAYQklglwP89XVEzO0tKsSufT0gv2+V
787KK/Gr0KkcDRPydwO3KL4UZyToE4K4EOeoYryHls/IzWjDCcuWcsyDKDO4p75zVWGey3H0Za53
I+hMxaTp3YcsM+Y9DKOxvmaZx/KVNX5/PJBpk5Z83hdRsiWjHSxoGdDcAQ5Q/ULpMM2QMBoX1vkL
rAz/AKbqLMySLdaBbmn/dgWNjQzowbggwRgvfKxTz0CJO891IfdxkKd/neBzNSltHJKH1ir4qgoj
qj2wPLK8eBJyyzSdU1Z0tYVi+YfdPqGsd36p1peG6F79i1vBnmbiGgeJlywxJ+43+O87w9BbQtCO
UMHHS/ormFQoYeJiO+sXCBvOV31/6bVsS7IWfNhtVohppIoU21sCHU3Uw/Xd+7RyVeny9rAb/yTy
Yy/nHAlD7hm8yboHJyEgYCyafFprk2C7wlzed8HwNK34MGZu+UGAQSW7a2G40wD4bsLGDAABRMIr
zbc/VOLo0tSP0AxF/t3ro0Jc1Yp+kfdoZUYLCAQLa/9Oc0qEfnXFf+nOs4FXEe+hdtltWEQNjTw9
Ycodlnwd9SSzFI/qVYISjQp9npAu5r+ucfio/IXdMTWDYAKDeGzxp4KvVb5JQucbtoE98/NmaP6j
iTLLEXZqKQivfb1y15lwXcNp4yKblmk3Y6sjnuMHIwNR7YblrEZuh4Uf+cmaTjmtRY/TWZuE1i4A
Bmg2S7//+Rq9S9bTi6ZabrFrTnMlCtgavYwhGd0ToYI/2mwtgs6POYr6N+0xlltiNZohjgUNqy67
4dCYB/6e6IXwJlIJXJZEc0GiRjhnxozR1syG3Vu12Wf0iEa+vcAxdrUuYeHBBpncWt4/ymIJVEmP
4vFNQzS6Fcj0pD+ScV5VQbJxYPNpkslFGAkjSoapSJTRB+7hftHWjWHW2NJUgrA//uGeoYHzmwj0
GVKH6xOTPpHMdCM9syG6FzFibtqhC3uyVeDk8w6pbN0xs/JWxhRjsCZziJFIiISIn7rC/Noe3uyB
w9xuPCSO9l5OMM/f80U/ioB8Qotm3Dj9MykSMZzeczcItNn+a3zMmhHNU+vc0vWuvDA1g9253GBK
JyXeOqIdX7mfbltQPXx0KxaKWdPhNyzEE2xszgWWjFlfhiMpzYUgGDKwH7C2LllmYVUFS2qFDDyK
nfEej+3qiIwoOOL3I5se9WKHB8hBH/zjKs/tkuET2epJ0TCSGkQsMmf59/8onYepfktvUgNEdNG0
zl3EYAqQZlAqyzjDpaVKS7982SsuJAp2auUJjaHXmcQiQj0WmJzD1vPOsJXCs7fXWeHUCF0ROLiM
86A0ANIiWXn1u25kbicTJEoO7rQ8bCOxda10XY5g7ucFdNW9wuc/EMLDXbxLVvCisQ+DTopEV1dC
6sQn6gtdJsRWsWVaTuP/f8DBWZRGbWGjWJ87lZedAy8JVLcOyNbgZBHXuhoROWrAyLDuID2O5do6
FRBOOXvAaisH5ldi3uiWdLEgPhItVpMc10IdzY+B0YHNk4oAc2Q8gd7uap1XCt2lWeanvap1SqUV
AjCSQnOt2HFywxi873O+TfohCEHhJGRrW+Pp1VwMxy1XeNjzqtI47iobLlytwGZsH3cgh0MHEbvH
/n67s8fjy0lysNBbMW3mfiBRQsn8YOfyUJvDBuV7mCLLG4EVtbyvrSZZO0XIREgioVbeV3FR3yi6
7JHF6WLiPx8T7uH7gPun5Tl9fsHHxkbjluOHcs0J+duLR8VzFTDWNWfhlBDgfbxS8z62MpITl3dt
QmiJsZ6uw/FKrea5QvT9NZoJvQm9yZ/D1CPSjlGYJUIjig03+U04a7joILLfDUm+QFrvQIhJ4Jc7
NyJhKY4nqeQDs/TfLHR61a+dySEUYRWceRMpmOIz9y1W4ik1n3KVC2i6ybyLdJ/CXvGCQdxZqtK7
HdAXYV+BEC4R4n5D5tbryVqoRToF2XN23dzQgDqhN4crSoL4KAmdiLu+BrRR8kx+u0ePMijKNSSS
G+tWqpsjkfDyNK1Nio1i/zcjYHf8OtTkvbBJcS2MXbe0WFNG27sJtYlCnR8RibcdqPLkG1Hh32l6
fy/kJ0nbCuDzmkGmuafAQbzvroZkCoMec/7aVZDRlO+Zzb65BZAvAXiskZ4gRFytVI0oa1HqrfO/
R0IUGCrf5TjyHAVntUbnECL6rLrQQjuXKAhUzkmlzF81zYAavq6UZ9cENc7JnWt7YvkICKHXeHt6
PI7WSsaH1pOsLg9SX+qW6L8ZMz34Z9diZVTFFyBjTyB7AKst3ABSpovdBYWwlz0WO59c7D2wszWv
Ir5mj1oVs7eWa+qT7HNlIc4XPafHR0JOmvj54+R+ozNdAcUak5Hjfjed6V2csKxneDV4vPbOGDbx
MRsym5NTknRtOVYYbXJA8G2YjyJ7oZRdc5xc+DNTf5VS2hRSAdACdSuIjnk5jSL+IZeoMjA0n8Tr
iWsmnAe7l7jbgCYbfLvdgnwUXRC5OGqoiZovnwgzWhtfjM1lQFzg80pKpkfqRQo9NtH8nz7jBt1E
BbxCFYgamYMFLhUB0ZTdPLZcEr9qMngAYO9kDjrng93JXkGqdZPz8puyWkmYzX895u1eU6mrZ323
2+eTBJLNopQz9a2xdjsTL45v8cBxj1Q8rD+bupfojMyiWkl7kzQHCW9+ZkAF/fedvaSvYdZOayyL
xmG6S9HPX/gAg/aLxonrpdFGjhNA/RojLKlfZu+/RmMIGOfKlgG5I/lOG4mOzfqYluqryCITYPUY
+lIG7rREkdI8U9SUuOrXwttVyJdH9dquP9VJ1jsfn//OnEXaS+87Zl+vG+VgEsBdO30RVFZl4iA+
Aq4+VNf0NodwXMAk1g1yTRBwiONvfOnRKDavsV/1USeRvDPFy5zyrlkEofApIrNT4oiImS95BVmi
hl/iaKA+V/RILvnTvq4Wx51MGI99ZpKzHDjxk2vC/4EW+d9DMdhr0M2gNDbRz/MeaiFNueID5zsz
MYk06Ij+crCqM2+u4AgOLxcGXhSnhTn/SLTbUOKTf7yDOnnNalDBIsuA/XREP/+QP3auutHs0uMX
zbh8fMBO5/ENY89qF5cJ1SmdtOOEw46pBhbPSwLxW+CnTzehpZkiIJXRhfHYgSXpla6COZoiR/tK
P182gw6TyAcRUUhYSh+HL+j3Q6Qrb8q659SKgupdD5nArEZE2L94K/1LdZgF6+m7e0T//rRONsJ9
PPBaPe0g9BGkT8813FRCqGmhmWaOEGtJT3PjuUir/cqsGVnh0PsPYDlDlQuUBJbdETqUI2CslUCY
Dh9xzB3x3gD56LkAqnvsu6gE4feAiNnJqV/XG/vKea0MZbs5zChco/jEZ8pGSB1DTDSjTGpSwkTP
BWzqCqmrWSrMrLkZCXr+oY9mPbJm0TFcvPf/9k5i+WbPftvfE7UfyHvDwzcsEH6gUzltObU09Prl
TbOQq3MM/Y4qVfXyVrwtYmrnZOzPwbiZvLU/UGOzw4cvNy+dqNYBYe6uYdWaIXwcl9U6r4rhPPeH
l39UDZARh9NCFzNd9urWzDqdwspPsIIYmt0z8zZlDYnlFHW6rji/XK7VLtcPwmaPc3aad3WZxI8Y
/efBoqGERLEImN8aB8X7C1jDHzRTGydrXqjWl3cRubR21VM0vEp0e6XVN7SmJDTlpEPnzcjIAlf/
itvFnjGbF/ij0KgTyJ5ecJ/dYRi8Qd4nSgdrXL8OfGU6ilTdQdnDJte9TdhWwgsAObILINxvzeCz
XmgpSp+yKsmsC6gJQgHBaB5KslPRURHsjw/S0VDuQVtoZe+0MzzFzvvTD8P3VS3Ra+jNF6aInTqD
iu/j8kMG/91dFjbku/C7nTkrXG+0oA3DW265uCgZaRGD0wXvv9r51rKtnqiqCK/D4PNCSge/hSXu
F0rBUHn9GeqGd/aX11NVJtrb6kDjbBbEheQmfsucA9N5EsYBNtkxFaaAQhUEV8SA8BRfb2gWIyFv
hRl3xow2078LB/qoujRec4SJnzyBW04RyAh31kW/lCbh0Kz0CC+FngzukmtX8wz44qW9NBlIzN9B
Wgvpj9PNJhfE9YB5rf1fhMEuF0+vEfqpQrP2Kbrn8HfaxiQ8GeBMGH8Zie2YzFgx/navm8t1tHz5
zdkXprYE+c5R2aqGk2WnyczUyvA3yO77JbqJw5N73zt3toltxwLHvGgQykqPuz+khMDCatrV+KTD
A/AxN88Zmw56pX7q3N3UZ+yr69pUxa4uwTfT6nlDW0BPeAxg5Xv0uQOwqyoQGgV9Y6W8KbkbwOL/
msNjsIoh/I0dFz5L1GtVhLJ9lDHTOoQ/MEmzqfnXUZVVUCSNVBPfPb2Rah7xK6lfA1XAxduP6gl/
zmqi1fbNzbDH9g+Z1PnXApHKDRAnlpD43X1GOzio/arA5urM0HfbZ7VkokTOplT1OKCJXJopgQLQ
lXIQ6jyn60U7NmMKCSZyCAYGYoO+761nolF3uLXEOpnP1ESxmHUQngkgXt8Yk5ePOTkMTqzDxuzo
RwGsC1KgdPKa7EU0kdN7pxy1td2GIEUPRSIABMprOEB3utYwtYEYL5AVgqwKd1xa2F44f87Dfewx
MMnGnUhHEFOB9j+FY6Wz8JwtERnhY9LNura8AboGq3ImFuQixI9VDMyZgP9DjIA1/4uWeUr56rao
FHDWrv2UvVnQQGM7wmrM0uSEZP/vqNiEPbX1qTRyL87uNri56bVcBO6ypIcVJJ89v9Y0ITLTouvy
upPplcjedrk8HDIxAk3Sh0D8cwQQ5fu3xS3nOstUBJZxB1jQuKAymQdKnrW5lMyNraJLD4fkBb/4
+AiAPNEc3/Iwy449lzlcHBWYdO/BlGsAAfhd2pNE3aLjVwjGrd6WOQ797zPHSnUwmEcld+0xgRI9
aPEti0iH4yNkq3/9kSBQDSRwIIXHGxGDOoybvxFDW9YFsrvgSk7qXUeL468VQyVInNKE/6lcyVKI
ubxPkr7YXhZKuoN1YDdmTVkKxDXy4/YT6Ape1BzG4hcGRvVnW1yMIoRjxzSG/jsKhTXXqyHw1ait
+oVCylxJIXlgEMpfn7z7chCfODg3TKuiZPpcpPYJO0olph/Tz57cdFhCXKSY3wUXSwuye4SaHD2w
bESp+OGRf7HhXMqNlPwE59TvwR1ZmK86qICVAo0AeOq6Dcjycct9YieNcAG6DN2yWtLdaK6+BovV
tK5IB1t7jNjjahluVkUxLlUnR26R7E2FYVqviKVG6TinpusT+5p4jkPNggfmBW0b1Mowh5j/qp6P
ayJBkDsVm8GkwdZnHqquhqsOIf/NeF5pNOOyKIT1OofFOpHaG62HsEen9Ox/o82Hd9ZcyYmf/ZZ/
eW5rkpjfli8lTcodL6eNfmT0A5GIKe3xE4RBw/rMSamV+62joWH0lmnH60Iz3oIed6laOyNR+n3j
Bcxgt96kTCgypWvJjKzHuDr5hQSC5wbcl6Ta3fQy85wdAKKAJVRIl5Zl9OPEBLggPOb9YQT7vCyV
yHcKa6Rq8QV/Xms+2AjDyauVSJJ43czFCvZ7Qqmes3II2ApnBqmV6p/fLZGUpdUIlE27v3JyUngT
vGmqtmCB1pj+yjNxZVxvzTMIWbTxf02e7kv36AGVdeG9YZ1QvXHzKCr9PpBtmYkB+2HsPwg/bywP
63BfJ9zUfwOnQxyIPak312wBEPouu/iF3LdBSbOjcGl+2cQZEndzfiFgrmOOx/0mIgjM7TgAqWvl
DFWEazn117UeMeecGsruMnmCXbWDpp/pdWp3+AHsrkiqrMm5TK7UYQwR+WdFj1KNNCTnehi/PgNn
LUAFP3fDPIW3unKmUncl70ceCCdE27AwXygi6ek1A02qnnEzy58jkr73XRd9Oe92TiBPsXvkK/tA
yptPrVNCge0C/972gVm/I3FwJhQxS5HTVYMxrUVdQdpJ1DkJIMlTlmzgHDxGLJjJg3RD57V24fLi
GZxDPUHnLmkg2NTG+48JNvatQwDRFR0NsfU/SL70ILFqPjBFlYUANLJSNbF6np2jBR+mKq3vZf6z
gzfCfdUVRNsK1djuqJof6BzvFxWpSsXCOOgRhJ7hpCt9fnB8ZPxDkVTPiGuuwvZR5PJDWGnaCGno
DDHcgZT8NVXrwvNb+W04Q0in5Hxa74NRb4P0UDw1vRT60Zd6cToQnO98LyLdXGL8EddR4pdMPHe7
pb/D6mRl14crKTgD7r8nAzZP2YJWSo7GGMmQMVwPAMFdMIzmbK6gsUesMVaYAdrb4M9rrUPm08mv
DtIBcQpR0zr171f+QhhehFApHZn81RQCCyEXBIC4CYsioUw9mpIYT1mavbx018Cy6DCvLlx7jEWf
t3bIuOUCi452Cdz31VobCKuXoQ7wr05s6G97Y0qy9P4Bra9tbuLIrGdlGl9FHd0ORvkgZuayZPeq
h93QMMwh/KkfcuVzS2DBARVn7byOQNuomFmNUIAM2okPxbWouEZW2aVbWCzHCfT8YTnn2ucx9wTG
tNPrNHVhuVOPtM8FrpNtJGPW/wI2pW3WNUdZ52ysb/0YpayMKoo9GXhXud7w/z+7os3IuXZfF2vS
vvxWs8INCoWiXdCVC0Ko/6fPVXTkL4WAHpL0vj4PqvjYD0uvtrmYHhmGDh28jY4MoBnHMbzBkw2h
dAEaoP2Ul2e0UY6tVq5D6tw2d8XCAhL0Rg2ToZDZqVrNpgVIvTvtZx//DpnpMuzQNfu8TWW5K0Z/
n9p5WRhTDwOh9DLjUdHNM7tUPW9b2KIU6O3LZhpO+TQNnuuvK8CzwskifZ26g7ZDYIXSxpXa4ydr
63IEuh4wjzu6E1QF9ldAO/WupL2nJ5VhrbQd+2vtLLZPal/8iOddFq3+qdaFe9+AW/jajvlXTo9M
FlmOQL+KMMl8qmXfGxoP7GQlhT2jBYHMWJDciw87xIjedpDo4/xZ1yEjBAFU6i1LmPXQHneNPM++
j/67NRWFBlAaS0MUgtF799oUVreltMqH3iNI3U7Nv9ZA7o+NlTEHmjjgymnLgDbpyXSjFlFDFku6
+rFs4zqFKNwEDVvF8UbgcyeOTB6DY8Y+FkU7p0Rv/b8sztCR3fU9UZn/lruyDJ07V1ZncqEhQ+C1
HoC3FacLMwr3muwr4oz+WCz7StCcnbAd8gUxOIHzGK2yEyoHuH0E5f9eVStYWZq0RD/HqBhSEAl5
G2S5ErT5UOyZ5gtFL4erPNXXnTpPwkTv8s1V9IqsLIRo+nV8k4DoPb3yDts8EXFPtLhL4ebHzNV0
O/r3Kh/2ezHW3MxQXNdLsTYPnOHPtEPL2We1JiXvogNmg/udiKoGMheV5o93tNacFwjKajxs8zZT
8UsSVywymdPAhGshFhvQVMBEuPXRtZ02bqsx0iexDLt2RXU2PAWGHEV7QQcsSlKakxKuJy8uQ/XH
fVOzT4c/UChloWel+K/DSF207mL6Byu/OF3aBqU1zdAb0pvIRJlY+KYARmRYQ3zp0GyuWl5jrHw4
kRV/zqb/SkdfERN+X2gZl4zI+Va14CoSyYA2dlm1HMmHLK2J0NH44MI8KXlqMzwlXHNYhHqHMGm7
a/Q146YATP5rT0DMsVgzJZMRl+xyTkwsPxQc7t86lhrC6pQ+VEkQXWYBP77cJm2fMYNVngQJLuf9
ofW7PTNTMfF7libJ+RG89qqymET8LHhoDnOZnZB73APmzmTFakZ/5BD+JZvPpBta+vEEYUOg1DrV
v9gibIcGC1N+V4kYozxULHv0qnkOJGkrkRTq0l6HcH79mWufvHTWB02C6k6AIsW7NQjBxV6AKAqk
+uWS2JbFgW2DrV4A2WOXMLQpI7MhXsXaRZXoTpd1Je7K97oujcxt/t+jXMTMIsY+VQ4fXwSDhGNC
oIibn/FWUrT1jcB93NGpWZITXF2uaBRXhSitU6AKy8HhAq44AahYk4eR6Y9OW1/rGpH5X+02LsHs
4OtXmXXtpFgZbqRoXO3sK0cnHQ5kOrzYlmtxip4tDevaEGbYcdrfamjRMOfKpDSPEVUAMftVzkhX
0QTcf3M3VdJQ8t1/VHR5DM2NgegcobdAvRecI5GotnX4SqzhX/nGn+BN3zh2uvsdzVfOguwmRfkB
Ha45nl/86b0dO5uAjVz93Qe450kuXg9jgRIT72In/FOCkp0mPt9GIJ+yx9F1h56duk/GUpaTsWo0
48qvqBXFgi/FEcMHk3ht9/ssUnjY5JgA8WE7TnLEFc4Crgccg7EkOeBU0cybUjkHqJbW+/wcPfxd
pXPO+8fw73uPT6ERwgXzP9lQZ0Ovi1Z2iVrQ8Lm0atYLfS0SplZUaeIa/2t1MXR6YeKWwhyg0W8E
JwbsjzCZ1cVinINn/iLPWCxrZNXYVywnunpjxzIrSh6zJbDS4DZdGBo9zMBjowq2rN3v8vg1DKJy
QuHBGucOA2NAYNpUf7znrCMMwC0XnpH7fQ0kfJ/ZDNWn5rapBwOQPhD9bu+apvY5941JeXsabo6p
2dzRsE2EeU5gLuXFnVdF8FCfeNUOuOmEABoeGlSwx5eMsxVFaJDYMo9kmUS6N8eI1qOzHh3VJZ8d
F23pfjhp/NKz7b17eYqBEwMBkKhl/FZDAT0ULu6bsmefvAbsSzGWoNPEGyIT7/QsXzY/98VDL2Jh
kRCu7bCRsbDsgEFV4sp7yueQ+oPim4WhP0DW1ZDuW9tenfmq40nhDj9UtR+9TyzTft53Vt23ihC1
0To+TXCz2inK76tDJek5qQJEQKKFPGngdO9/3fLiyI5AeHDYDeugnTykCGQCFVhs8GhnkPH17EZy
/qcej4fSmTlsyX1O+DeALy4k3InoeMfIuDgDmHnHDzq8qTSTpM+vWrJXDVehoXsf7vzv6ZKvZFqt
4nicCNJpa1+gUBHTp/wK/ptxKaHgGhvanAQd7Gcw26q1pOR8lXhHki52TLaYll31bJqxqSXwoYs/
RqcGIahH95BGWr2obnQJ12qVwisJl1rGoflD5AG5rn3hi37AkyDEznTfJsgQnxYmCChnbuaJUx10
2dIO+ZTDmMly0S5z2IjHnnQSaL9/T3GDDGlGQ1oCqZ9qrwyte7ptJMCZgBGz5xdmdfIVU3hWjJkt
K+kiDpsPp2eXbqf9JbSdVCVU3TfBirg278zHNe1wRfgNlGrBBozWVutIpi8lvo17SX37XO8k78Zu
sU8os5lLSyjVNX/TV/tP4wwQRclxcc07eBsNitI98ST+cnnT/91wfV9pGtwBb4I2jC7SqSDMjfX3
xfFLNyLqd8n7RWgFskqoVF8RfS2PiaB7HMmmdk3PnZuUD53fNXmbyVcH3qSo5rehpBA1tY72WkT/
rNydxyN3jbkEQtFFbByvXEmEkKFgFbAP60u75/jbTFx6McS9fbnkc069c9+gy0eYjhrTcKIXpLmr
jmF9UXCetmO2YTEIJk+WJb6VrkqhRiSWUc7EX+ll5yyRaeG68l3SO63mmYuW8RkRE02ixy80v3Po
Q9C5LSaZBNOgJKifJnSOw68UjxPDGfTqlrzjqfccxAfXwH73mut5O/aGpAFK4plc0jlVTG2kBFKU
9IheWe3tCzPyrx479s4I5KeuZxdaRBqJJGAg5mJscazQvyfi+0547maM3l9bcCeKshIl59wDCa1C
A2o1rfB3KWSkYDmkH2ijB9cypkDzwJ63IQvD+Qrk9zsR9qY1ZgWTbSJXUI2e1+9LU3NmNIWjpFMF
N0R+Wh4pSTRdW1kcNyhh4ejg9/43LTlhfT0JlI53hsw98/KYsYrrJoE0A1kmOHCGeJjLPY52cA+n
guv7StXsmpi71PszWjHga7ipkrjImjZFoMuIp3EP8dOTZ3bC5SZaqBdUJfBJoFR5h1eXqnXRSFUM
F3Fl7nDGTGuYsnjaU+d7Gb3H/mVjfEX/SK3fHK9QncnRVTNdv7BNFAXh/YZJ99VNsCLJ9rPFr37p
jrjVnyy5h+fZiz6VWw9vW7EnTGfxa/MygueReSk8iNJV5ss/JqEW3VNQvict3whP3CxOgHVJmVmp
pXCb+6g8BYkHaPlzmGKUnOxx+jtZXtlJvgWfr7i1nUiaCiF7vZvUH67hLWi1FoaoMXF3cn4FLX2L
2MRVkLHN7lv4KT5cBgC6ZwDe1vShKzUFuivbWgnddNP26jFCEcclQsrG9HSla3wycDX9e07YzSAG
5vwu9Ud+bbsV4fS8WzTicxZHhxIV7W8vQ/eliMkZU6oIm1ze8wxY5ov3CHnx1qcwfSanNZ3/NZQm
8egaUSdJXlulwpVaC6mjl6buu+yZMryHD8UwN4HzehLe4Amad3Wu8FaRIjw8cjLUQB/xVXeWarM4
sOiF1GAHEJMt2Mnx0z7YZuK6XmQ+scZ90NXwi9IIFOuX9udrP5i+4XMg0VjVjBOsQzMu4q3R1dGf
kawmyBCzi/ObG6hvG0fChDxmSy0t6J6XWBjOeegUId1IqsZ3uSqgkFwhrh0hq6ttaESbBgAbVhAf
ZLOcmGut85igS6Os+zSPopk40MFIj/sZMvQphPJCAbbLudtH/O8sqkEW8NXmNpSph/SC6a3ILHAd
uT2TK0LPsxCW548XjCjt+7ilcKc4AW5uRU7oXKEmxZWVrExmrDsZW5zKWqiHxQZbelD+ppOxJaGG
cfMBbzEiLWuGcI2eJnXqRY9tdkN56E8Xh27US2dIqMfSI2VznRY5SOaJI79JoLKv1ZqJ9X5Hwa1F
5dZDP0XJT2mGs8IUOWoghsYR0wcu82Ge4+L9NitXCWImhJtnjVMKGpFGRox4jhEAyoESPH2pnfVx
5yk5s2x844lep+4UvjPZ4GA5MHUxF2/vZdmSAUd2I1IH/A8rVrKo0qYFovC1zPlVjcxFs7TbeRuf
Sde+Cz1n80rJEa+gg+GbSrRb6PAmSOafsOF7a/9Qf4ON2liUyAppNwFrkBxPPZNRCBlOzfdOIkyy
wwi+Yh2HX82zAyqkqGOmfd0wD9s3CEwzb1EA4wMisXTC+BoZzSf0lCsZ1A0u04xNTmycqWD9cqOJ
2mQv6NqiR7M+B3G09NhZNPgUvPA0ZllHbDcTTxag/fGtpAxr9HdYDgRJBt1zsIJ5iRBJw/0DZYMs
MVg5bvQUReDnnlZw5h3kbolBT2AthoWLd+41fGbi8hdVUH3ryV2nzmT4bBqIbWCUr16QIoVIDfAf
f1rBVBPmRtQ5HUi1IyFnZG8HnOUpmMU0rQUN5k7UXafdplaVzMWRRqSmusCjnY1pP6nHNepbK1Qo
iRKJ1EK/gKnLMQtLz7MHWVARJvHrUv77V9LX2iLlAB0xHbdp1GazX9PAzB9KOj7M+bIhRYwUHbD4
2erbxzNXJHzer8eA1EC6akphSCWx7KSQAwimAshF4sw/uEZBErwn2vvmkyLrDNFtIOJRs7/mV+wP
5UdHVoe4MROjiTFr720Bp4BdZe348bZO7R+3z6QsvWrYcdxdGyGqLo3GwUKJ1dd3Ny54k5/OZjGs
c2VmAK8ObI+zDS5Jie1QN1OfWmkRKkB70gqoY6aHdtp8hFDzi1iG5AXlzDVXX2XwQDaY7CS9xqvK
z4w9PNn68t0VeT+zsf1bsDZDsrnsfooMPCYBvtwTI8UZoitj46kf0W8X7U9D1VJp5MVkF1VXIBBl
W/6g9snHufy/8+vzwRUHroGOoxTpmFmvboHa0K1NakjWh8swEDEbdzeRCQd1GEprWk7NIdCYe2aY
QE/wHk8U2Ax0mgOMSXq6KIePi//Ki/fsFMuXeCxoMdavBcJ91YP57UYMlRmsNKWIT0l9AsaLWGxq
8p5b7LSm4DfmwWKZ3Vj2HFVRkNYv7QnNg93B9uGculdzFiuokN9mngdh8ChXy48mvNleHfsm3Oxl
tVhInqBvIcbYIjXDtBLh/pwArd+JEtDOofntz4dEgflsdne7jnLqFiV9WQUkcyK4AiN4H3CV249a
5pzsamh98c2XXq5aX+lvACDMhxWKHssiFkbiah6H4fPYErpkTT85eWhGuYzDJIFtauxJIoEvQCfw
KUdm7aPif6+BDCxw8/bnKY7PIGsoh9HojujVeVLiSxIHCkGIVvq8DgLYbNmPuRtZgs0viYcGUItQ
rWeYOvKJs8LFobnbIHCwNf+/dsT61qOfiGVbNakRoXvAb2BKbpWZOfmeuzOV+8L7ajf/UDljmvkQ
h5gPCE/kv5m3q03qcE8BHMVzRZEfiWXeBt00Bmfh00xoOhVaHZ8NQ05kO0IV65GRpffm6sf2MlmC
+UMTePpU0WtaRdAn0CC0Pczq3nHUAox8/tv9sAGDciAZjZItZ+CJLya00lntUHoDLcVvrO3zAWNW
nssezlLAV4GvSJ63d8nu9TBjzGr0J+vDtDWRy+YVPF4MBwFhcP/VlapT7zKVKz/c/9QHfRbHbjep
uxnkXqVpxGKgj0k/uBJEXKQBpAR8XKjR2KQ2LjP+ztudMfKkVjs0OlB3GtsC5vSQqv7EKdqd1CLa
QxeHVRiSaTtuwJGIAJieQc7JytpzieEEaAlr5nvfuTd7C93J32oUJvbwgQeZ6OKHsSUCwTVHTuiB
xEhd3TQJBw6yTclGDaEUoO+2F3pmjNz5DcVmHekDhB09lqAGNjP4E26Vqq8DJyRt/t52QlOlTUJF
nHRKjb0WFhIPZ3KKm78lw0PMs1CdkivhRrrgCFx1NdBEwyTZCHarT8egFFY9FAs8+gBmSspW1SGR
c2AvXppyO/XIU/b1Tq4fEvBR3GU6q8W2v0qeuA1L2xDEGYrexo9VpGEdsOXpRozA/vc+lntc2wKF
SxB0syA3pXyTuwFZd+d3Clf7dxhuE8PA+KIAofjHtmoM/4do1mNXH37O622/PI60LwQ2G/swVU9+
g0rEyH1Yov9anhjwqc8z8YjsBEkEeVgU5devxMGVEQ7W++p+ShSFaX/Z9TDf83gOsFpRuKu/ubec
5yFczXKZpR/Snjd95VLzjJyp73rjDQDSdUSdkTHUz+TLjNmD6hUyNyTfsOGItIVTlvRtp0Ghu6dD
LXGReDSTgGpXR3evEa/xWzqLMdJ/s52gOetIxQLpr2YjKlup704Bokk1LYnCHimQ9nrIU5krE+Hk
Hlnq5t6D6S3yVfbT2GWDqaIqN3jlfagvOQdXLkAZqHdz3PrzIuDgDqTAZFIZaTl76yc24CgTeae+
tZduppfTMdo3FKs+0viIyayg30wMgWtxepAZ5jouhMRs6/ngFhlgiDQe/l1teqPyb9dNRY7V+qBy
pIAZb863FmwztBv/rsf4y6stxRZuJx/s4oQIzbGCbuygIw9gQGhsB5lRhj6pVroosYNfmIEzFV+1
01/m58yTTp1pqrIFnTwAuGMRnTp//j8yPqPUEead05aRd7AVJSe3GN7RX9tFlGV+5haEDQkOmWZc
l53QOwnjRroMmI+txzfwWR2GHg+I4DM2G439AXFK3GKBQmRRtentNECSqE5xC8lLx0gwPMrfs1eC
GsDVq4AKMyKpxXBc2wWtj0LQOL/CQaYvvm4OPkfbcS/9qVylZ2LcBR6qWR42e8NlGmPr+FAdd/Lu
LDSCRncS01EG/dkReBeMzMeJFr2jN1lqGTqLknQCtnj7WLJ/Q0/41ScFmoRyflJLJrKxgUIIQniX
K6+vQ0dplWhT+vM/NJFM3nqmVuukJpaQeefa4jfZBE1iFo0d6/KjBCJbMQ8J01jJDQCunWH5AzAm
uBQEBLbXbu2bGZNpPlZRBPNIWiLAjuVSasPVhiTDsYbGS8aDExjy1kfPjw4ur0eDbNuwq4RwQIH8
lELX4IJ7Zamriojl8I44xTSHnQcozu6D6/+U7SZMPib3ip/kQJWQsdd8Upp+GygfjeRaNG36/qus
wIm6YV/mOckgRGLp+FGjTkPTIMgwy7/nn2pkqmzKETHuVKeNKUvJVJwvxx3gQhhtqvMfsWWLNEdk
ttu9xR+1s5XfzdcvZsCNZLzmnz9Me//O9zWcuNk8XMCGfZse11k8pBf0j3ywxJC/xwmi41Rytejf
aIgd2XNAf3HSgmZpBJMWXVeRkkKrTZR1c1H1G/bBhFumOLvfOvQ8L7nPnvliYE6k56v0Vhl3anEX
0NDJ79fRmftT9rJToMJ27l+1yMYKatotXZBsntEFKRNrseS9+4CcqFrzc2krqOmMy2s7A4cxEdRS
XJUzEiazj+1Wkbch09YHS7YNfKg35W+dWRf59YVcElWnURDDjjXvhd5uT3IE5IMC+NdFe0gIWBdF
CVuG1bpS8lbQ0W/F9pz+BgNfD01IRJ7GDHefydU+VEXIkKKEsv1omnvuxABHuP2AUsxQxYcJd8Wc
NpB5XMasTDll8ByxwzfzTu/E6cKTWQW8GndXwDVX+brFz2SatAYFGoeQp0bVUdejB6Di5GXdnlGn
cxk79QoS2Bt4BI5f1yX5+WwE/XrBfyxkLzB+OGYBjT+fb7BL1H7/CVnR5dLlqMJWIa1PqFd1aD+x
kqLTd5tcukDZoZ74OJ7+rte/rVFsb02WeZ5X4ODzSIh51RS+JCauOKDQFMNTYAb7OTbvaYd0GDaJ
Stv4f/gHVD8VE5sPJJicjBnzAwM4avQ5ExBhAReNEQuJAUrZVoQhEOV2UyarhrgFYtgRKvTAh9+/
Iuw3IAhXCAS0MMpmzQa+l0oABLtZ1sarTZWHzR8B4RRKBn1LqWmkItTttlIG2mVFSE2DLwSA5yqW
k+8YaTZQPelwmqTZBGgwBNYzWq9y5JP6AZiwP4YoTiPjjbF0zIRP1LNDUfwGeJlFO3IWwesmgMqV
HTLdSz3gDik0nVaF5D4RAhbEpgF4JX+n/1zvKe7wdH4QXqdidmX3kfgIi1GDuqbalg+q/OAOYtvM
Lwn+670299n0KEa7Ihkrn6gMN/Cwrek+5sRV56FCz6JUmfNjP3ReIJnIH7vt9ztWnJJ0yGb0IdNK
SLYoxaZfuMvKndBeb9TWFnJwIBw3Y7BTpAfTB/dC5MDdXqay1mX+1mAz9xHja9LNKdPv8MZikf6X
PQzE+4JtYwwAkWwdT/ufXpBZLQsw9B+cVK5wWHiRInSnGrT39UHd9ADPsKzniIW2ogTzA/NLgKPY
jSoXZzEndKiwRak7Cfz545upc23GevbYQ3OUXrU/pLSFmoMkJ7ynmmmChQYc9Cj6YXpL0CcU9+Bn
MPOHRfggzEE3VXEGyJ7CVtwUJmLAVWY5GVDhkY8FPYUXRVohhchLjhghiaih2t9wU9N3gv8JidpL
eRd9lZHGQV/Iv166h97a3HGFgF9Wqwxk0YUDRm8jGM47LoTreTsqatk7Qg2Zu/yZlS1GRJzxzkAV
9UORsx6SKzicMEoWVAtVWRWCQ3SbLmkf5QAbZ/FRj0YuM4zRpMkuM5Lb3/PNkYtMrKCWUfgtPyHr
9c7YH41Bj61UX6VJ4ebWCKq4gOVLj0EVn+fOUoCstizBBQqkpkZdao6VwrIN9lLUEfHtkejgGjex
3fC5NW0hldSKunx5plezRZ7N22Nu9/8HjmrZ5zz+cCaUJj6NHc6GsFxH6p/Vtb1HPqi2pRxK7JLE
4b5WZDuP7roVoef7qTkQIGDK1p1rjaXEutIUYh62kOk3RJE/9VriaTm5/ZY+x7R2cxzFkqrJyLwM
fiwZU2INHWmmPK2zhgU6Q0ZxgNjLTbNWIca2DoER4YJ00izXKmoBiGgTQPf8Ju2pgXXf/yVoHnjI
8yBTw3NQr0M/AW7yQJCvbgJactfR8jWkKFD2eXFrBoUWSmcAYwjCMhbzPJV4EK6SOXx3sDu65sIQ
EF2MyYs0HBW3rsXo3tiQIuVGFqF0btkbc8qnAvuhPhLvdjSnT1UFj/GKX0nQarY0B+NMIAi83hNo
RxTEmdWQm9ked70pLkgjwlhFMlyGW92Yi9D9Li+OCwLZqg/4OptVvoi0rz9J92mnm/Fdiw63epL9
cE8cPhjhNNBo0wsnMMWGhIdycJmDWBPtAZaVo2DLfo2cJJWtm7RPXpkfETjaGg9SknwcFCUilwMq
p1vZrTTfZorLitl9yHwhlx6CMIPcaEEpXtJYvRjdbD2dp2kKBGSW2XkNbw4d53f1+V/U3hyWXQUf
Ykd+e6m2/X7aJhe6j6BmDHHbCR37ZJnABkqio6R6Pz2JTUWEVky7MZKpyil+KM+2AfrNGRHBxlzG
Y2I4HU0sACqdAHxXYCpNcCvwrfPcPUoIk4Mdrqdh2yslXFZt1EOPBicPG32apWIIlNdssLBhvR/0
wFzwcWl0xdUKu2VISrmWYjLW3jkcTCs8NcOSpM42k6Cy46yVgoCWOQCRZ1FmcFct32xHw2BnWtOF
Djb/3uKCgDwVrV3CRNyoTPGR6fPywlPkM1f7Wm/wg8/NHyFLn3k+vfBbIUwxabSEPMO5Az2+0Ucv
obWNQnoMwQLXTPqvy/dXB0UQj00OLHI+3pomnRs1LDYw8HqAQmedfxm1dnKBwY73mieSxU6YWzQl
G7CF2wiKkCSBxDdCql6uzzQEPkO40FEAuwsmQ1ogW9tuXeGGmNXRGGBQGqFkNxrUd4ELfnOkNZAT
zxHbcvxAt8GmqiW5XLhyfEzHxNWqKqysyaOi8cNljYImivuCu2TJ/TcZ0hHlJODVlnep18FpxA1p
SRCSQoEWjbOxAUWcFNTnFnvkJX5LRlkf4FctTY9wFrYA3l9PJxfd3+G8FEKIERWDssF8z8u81QBl
hPv4SKdxhsr1HQ08WwCPxOjWKiQ0v7DORLUcsDH1+UvK04IWMmjvZAxeTdH3yng6d/xNwO544cMK
kcaVBf9J/JQkHvAAJ2VhaKlKGOjl2mPC/omnq4sV70BpQuY3zsv54QtthWLLJ4VAjepEh49E7Xsp
WnROWKGRxsGKUSvrNEFr0qL+lJqFWsh0clcQ2Que7B7gWnRYJ73xrtLwdRSBOTeIypMtBERiPt3K
NKTDMcTPO4d0VudQ8JDtbmSFfIlidorqefm8zP6NqHEWRnvAZTOg0bI4PNW7GhyPiV3vVBhUTvel
IW1aXQKnn5pDnWfgQvwaHY+19xeE17O5DJg1y1EJmezaNKuO7Sv8n0u781m+BPX3MTUUtvLKbYAr
X/HI96qkFDdglFi7YIiuNqSEPwf+Rgc4PARXqplsP2v2HAiasMUkW61cbzmiwk4X5CA0XE5/0t+G
7Hf+pg0C7m2VXP5apy7I3lt1cjLofFW1SRp0JLsO6GKaeNMZf6e+LiDzPScaCB0gsncoTXxAmpHB
cRKDCy4PYDQHOdlxs3099kX+5zJtGsbKDphcvfCfnEpA6K8TSaOl937/DTHX5DhFwu7LN5vXXsDY
WE/rOO3xGAHQ/uOZnIS8bvyKBPCs2c67ciLHmKI3vmP2fA4BfT6QxryWKDQdB8UnTvse3j88+ca2
vTttTEkkoVonxb7eeR6RFcCO6q+iKoDCLd9pFWDAiewg7nPu/xFDP6p134lun/IZnELJbo2titpW
IU8B/Jc8QOZqXviGVucizlwLUQOHzb5VdwyUsmRiYTCKOyQ8btFPYn4Z6MWzKo5GTl8nxRvuWQmn
2FcQ5tGzdDM4x51b8q+XxD25FbbLqSOc+qU9N/oziaEtvZaUm8/jlyi1ToMMLkMM1WZSBKSqqDvq
Q/oOgSK+lhN67TfZMfHtkIK3NHRbvSy9WpAgV7io+b4XGAw0Ar+iUztserhS/KZiKQobCLZl6x5q
KDBqxTKLUpnlTEv6rL9SjnBk0OLkLMiMZMjCFIlcmMfgb0EssVKTdaFrjlKaA99dBWHJCxVs2VQ8
1Oy0IPyMYcGhNdTeNP6UeKSH2BMta60rvbJb1tSqt8zlUeiC42PDnx7ZT4a6cgTB12U1yEKg899i
aKFOGhYMRcqbrYjW69wO/I04LSF9zpvYjaHHjrkVqtEmJqfYEfZjd9sH/p/111kswcIdFiM20zKq
kRVsqceMS26T2pabb7t1W2y2JNLzX9Yr+FyIVhS4ve5Xa1fdpiP6GqckqIXGtIQq2UCRTA9uy4CU
vqhFMBE3IiGhN+pdjwWheSvk7eXGOK3+pwR6Q0VtW+UFFML9z+HYWOe6CNMNu60Fkb49+HNkAkDJ
oMfKkcBYPrbjNJ6UcMXdLnzeOOpMsU//m83h92KNZdipg9nOejMscRUdszRgS8Vkf8qffBO+PTIg
PkQHHmbzugwXPkzmQf1leW4rjda78+tif1yswPhqumc8DerH8mrsgVxJBjaEtM+6qXluACME6DEN
YG2kkJF5Zc5iRzMoCGWMfBq2gSMyPtBovgVL+TpFxfw0EMCOkRfddWIhZDEq5oA28VAEp2jZ60oT
65KNpKYv1JOon28RMflw26940Vma+cwBD7uAI7N48zxlRJPgzd5ro1zdFSjWtiAB/LN0Gdn4Zeqg
N4W5yifnatp2G3hIVzPL5BYVLoENlBEOrUwaeiNFK5FKjvUpg2VaIzy5XP3Y+IIb3d/Yb2LpqD50
TcZi/4rRAUsnQhDISnTNRjfm60nZhby1KcEbKFoXmuzzh24I87wMZcrByhNE/pv0xFVjiGZEVOs1
6sscTnI4ryFYz02d5225+7Vsfh7rhU45O6kaf8CGWYPeuxEDb7AnDTFYYYKVUXdcxua/O2K2Iejt
gABHfCUl6q2r13pSDCZyWd7QqSQbJ+VVFNaYtMJ9dGaXoV+bxDfb7OZabfmUpWcfsJw23dUv3wbO
p1zxjSyf0sOgZ/cLUPVYsig6rULlGwBuC8lPqPM0S6GzMnB3MZIBI2KkdduYymelIoaJyIZSirkY
UMphmhATljbIZoRrkHCmxDhHBuF3oxlR5x9187kGUIL1NNSVL9JLenFSoJMA9RmKmlKG/oCxdBGp
qrwpU/BVmgrgSYndZh02uNyLMTUmB9AZoRsH3eBLEUJwrvt8M0bsNuFImO0DAdJiNJXLUYCd12YL
g2GKGPa0J9cDx/B3V+MlEeRSC7Ds9b12AXUZc9dbIwQc1hQsAhd3XtLbAQQmS9MlMtiE/5lXbNCR
UleLOfb367tRREx0uDoqjbNXqT/KPiQfSbuAI8l9FTSKbSBLoL1vrELkEYwD6UzG5kQ46c68tqH3
0qpkeU5Um39qGOmjXAysgdw/J57UXSeM6osDuYNg2pHPTOLCCyg9RWKBK5Y3ZpbP8CmyP6kj1m1T
EnOOM8FL1adiv1r5a20uHplUhftW9LuhkEb+71Q643Ye5wPjNT5DSWYl9dNRil2HDMVNHmlZROBw
UAeWBcaho6h6tqkDsSQezfeWsimNi6nTOjH2WGEM/OGguTHfYql88pYoMdjqLsFIWYDgItFT01pO
VNqC6irvb/IJ+rFpgUNAW9b1iKUQyluJ1kDXaNeIrQYU5nqQGyNVO367S6wvbLBtxwKTPYWCSYdE
5tRClDOtzpXBltbt5qUdQOg75lSEH1DeowQWhW782X5xDF/YRBas4mL+qt8vfYJxZFSKrG0cYFHX
2thLtZ82Z/DRftZVNN3v/arM9sOIEaG2KMhpWCBpVxahuKfKGWP+mZxlCHJf2NpGxTQvk4YgLU07
PT5pF3WNWCsskZNXKNpXZayjo7eYtZvyX0dchF73jKHNeqy94e7WrVj8V2+OawhKLDkMLoV2rA+d
QIykZOvX57YWWXii7UcUQQ6lYKxa8dIJfNMow0tWo6X+4mNBWiCVrjNeRMGRxuuQ09BNlCWlJT8m
LYSVid3GHYoYqJ4nAa/Q6LO61bGQRsXQPbsoyXqEqYz59ioT93pofEf/aUej1BQFuTx36WOlAiqX
YWZghbHvHb3OPa/5tV0xJr5a/CkeBCyG8+mVG6blGdXY5rET06mZmzyW+UWgOKC0Cd6tdNLdSADM
DSqmUOj0YNjHFONhoKV4MefLPLZIDTPmXuOQ+FCdabORxURAdteji1scTyKEzHhSUVcnupjD6kQk
Xkf7pgKanyWG7PrdnL+42CkB6RxxQV3Fd/M2xodm/SY06X4n9JyDJCZi9EaTSvF+QaYovpzMHCDp
h+vg0UcUSvgbXcrwGER+3tYVaDt3vAfZJR3qeiUUDclhjfqHqkjYL50KX0Xh6ppCOw9P6Zm8/vUb
Hn6dMzIQcRgaD7GMo4IyXCqIxOZX2OF7NpA3QS1sjmPt6MTPTa2U0JuTMN2pL6Vmad/BN/D9YkZu
qr7xOT2XDmFY83a9QPBS6RkokCxJBRc+9FoCjqneZUr/60EGknfkVx4nn0Am8Ul6Ga3JymdLvp1I
Bxw1zxPTaSPfQTf5niQQexTJ0E5vtmV5xU0fFpZK2Li69w72/mOvv8tGtCwveLR09O7tKCYvox6l
mqZ9LbJQTIyxTdx00o2mS9OD+ua0pqyFc1ORuFFtY+J/TAhQXefmMjxhY7Bfdlg5nWLaMfyRC5//
PTVayas4je8ZmiVrRgRkGul6A2ruTAydfpHXm3aLFV8kqNR/XjUXX6tvwy/hsD+Bp4yecS+PjhBp
UXQgY/9iP/xMIaAunIzFQBCT8KyXPOVLe2Q8nEi0Fll9TI4BpycG0KbBU9BNnQZkx+ZP8ECIra/X
BdRGKpoQRoSfYRUdrKiEhjvtr96Jcp0P6FeoCx7v8EGujSW0FC1Rq23QLxGCOSKaTQT6pwlpiTxU
NywZGYfsWU4+Iw+jeISjgyIVWf1VXRjM1WfteEUnKZx9ON7SiGXlGYEvbpCMOn2WJdRkp+CzQc2U
nJbNO5ypRj43BdEwCB1uA0lTm7M/D3DU9fS+YsuZGWxjtmEcYShajZ41k89z3Ya0o/Xkkz7KqX5s
91FzFZU/DnWXZcKtG/lYqtUU1GhUcRLG8lUHwWTJZnqzVE3RjjB3SrZoq8v/YO5UvwDdi3D70Rc/
SkMjK7EG9jOas8NQGTA70e6ZIa0mzM6kmIXXn6dAQdp0V65Lrf9XkK+6Zkps2tYD0FdYDhG26xSM
r/2X2DXhj6bHW7iCUxjpn9YbFxdCH6R8qtwwfktM12OWqcrsAOzsNMVCil1JaZdPpVrWubXS5PzK
FbDosXtBwCnH29MvW9QtOh8W59Rqai7TkUezQBugwQv60v42fw9KrFe6pqYv9/0bNX58uT7BmFuq
aayfWmaBVfZX1nRo/jPNpfx2FtfPDM6JkFzRnbg97ST/f+pkwIk0s02Bby+GspjkmPiAuMtJ9QjF
ByrhVIrgWCEhzI6eM9rv78G0eQOw2mel2HF28syVBbExBQHbxEqg2gDHorSr2NWdIw02jjdjofXz
JKGYVRWpMJCn8ZMhRzc6bZ0dwcSHrEK8w8ZqXHfQ0eSMOGh1xkDNYL1iouVXmnrsJdOiqE7NHhLg
2tWz2vRT77ODHFntSWjvJHJF3rkRbHskV4NileYEZpzs7iClUdF31A7L0q0p6KNVopSS5+4vSVC4
PvkkZ5yq8OxqfXdQCgDXu4zgwVXXN5cJXXzuZBLSCu+jjHS7VG4u80bbfc/X0NiXWGMktBpnlslV
EaOEFCceyxn58XZBbcLwY7BWihCvDJzDSb1T1E8dHtxuhus3AdGIKrk7aeFpXyCfdF5G/+jlXZ+4
jzQFX3lu0xJRzEXf0jeC38IKYbE66OQsdSugP9OUjYUCLJXsdoFXeUu2Lxsef4cpAXJSNY3a3ei+
TAiw4hVj6hl5DAtFKi0z0nN1AbcuslnSTXV2aC9TJregfQhhTCAiGLqctV6mrhqtwttff2uyriGd
bZh2hAcW6jTFrMEJnopmFTFC/Fz1Xi0GdP5LnBnbxWb+cUG5nucaFDJrZsAGiEeWRsOMtzEmLM1j
f9gtOmGk0IyqfFkoES8bPvElZxH/cQ+P/uJsT8lP0sB2lqbPStBJagnBhI5nsPDaVoN9nPTomabU
t7CkPoFuY4uAH0e7DPDw6lpHJgrEjfwhV/R4nKY2ccQUW58jV2tEQ8SD00qxHPFU1JugOADARoD8
+zztS6x0wmSDMsVSz9Htxr9O63Xh3pUIlpOvKqbMGmdEzFkoKGfnG6BaIOrbGlmFsRAekp2MfgZ7
uF9bNVfNBMtY407CveYck4ft9dXQfGcMJuD1HZhTfn2DFWTHnZn/gUmM7gyLVjSUJpLkrTEmRiFK
7ETbf1nfV9quXjDn9heZD0WbNCN9qoFaKjX41Yt3OvJRxujpgUCWJQiBk7rE68OX2o3QJgvUw1fh
V1M3WUjYupdHVI9ryd8xzO9Sk6eqIV7Vh1x0JJt3rOkiu4WksazJX11AHgZEcfxSrjZbfpzWBrfC
j5ByxQVYlF9WsqmVNPQxNPFn5KKUrHu+NYFg7rcAkF3q8MNEKCIOcDqvrD2iL5Eo+WR1W0H7ZZv6
WzU+RCTPUUDiF/nzGUYV85DEeaHRetZMex6417pb4mCgyz6CWAx/OHiAfVpXdUnvFDndUFG006Ka
X441hqt3dpqB0iibtRNroPsitkqsVCIqWWaPluQtsGzBp69fOrCOa86pMG4srt6HMM3ZElqflIL1
69x8MpmYCsZH3MAZcE1ExmNt/LtsyA0QCwATcsPcDeClofJvM3O9sGAE6AEtBeVC4+ftmC9N2VXI
Gs0Vpb7vktgN0VCn6i9hx8ZuutBbbFbue+XL67/DOu3zvfEins68ruYi5r4Gk0bc0qcoD7wAf0aB
ZdSUiIKrshj5uMwdKq8foO/7qOkPAR4Ct5qpgpXcsS+WLTLjP9a0Hth94NnNk/lDzuFYnCwXRPQj
PkKjGoJvQNIQcyb8qild7W/r57EVmQk9RNtTQLqy6seNcv83d2ZZUHIHbA/GxdDmbTVDJyVAUo4H
kJ4l4uYBAhh2ywu2KA0yz560l5oyhYHqUOqef7epUHToM47FctXbUoaeHDOYOzU/wrtvwXcOg+jA
wnzq/NWVo3lR98NkpjVGMdttB5pUcsdUrIDwJSBPf5WC7qi+khGpjo3GDagMVeMXKLZ7AXECNEg8
FlAQGHXflhfcxDJFN9wcB+FL9mDaffRJAQS/lVn6WjwsgIewq17v5s705q75DfuMmqM/wiH7PBqT
QS6CjSJc+uC4fxp1mI/BFGxoOl4DpjgU5ga6xfWogARw5EAdqeu0FCM6VVFWBL1m2Uv7rjNrwCdN
uSbkCZUi49wLgxaN6QD9vn/LXmgGO1NyBD7pmopBUOtAB2ilyXZ/q6SZUUzKLLPA7li+jKqLiUYp
9ZxQxWiPpaw43Vt+5eKd8fkWB/h1iUoHiIn9k00RQTTDAjT0gDUuyUGRinlQf6mwCMwz1ysV3+1B
q6G6oqHyfXBpdgOKKKbSDpxij3TO4LIrC2APu3zYuPJjE0GP+hK6aujx8N8yK9UmNeyLZDMl7AUT
2YschInvU3GPIjSFxx0nKTEKde4ou0pOFmpcHuNw9AEYrZZpsQwdF5exzrrLsIQxaYGn0474PmIL
1MdePgh+BvTKxoWc332IirM9BKuNvEiEldlcBDouCba7zUI0aIB1na+izstBTeN73+D0/AMtjDht
a3DJSiE/4OQxK4PM4Hyf6IuqXJO//vjormIaBmMoC5k5xYdsHsWYnoZ5N+wIqa7o2spXGB6+O7Eg
LdoEJJHc9sV8oQQOgllkPeCvcU1dz6egRwmfBRd7sCVxz/Vva+Wc0wqBDHx68HlXImluXMuzultY
pDFFA2pBwIUX4ropIm9DyXMKEdLVOAs69Fqh7p/sQGPtTyFNENNCshnxOWcC3KAFlcHZ8GtICaEC
ecYfVW0xUo4RIwB2n9dE0FMMGLwOum6iF24hXt7jjy5We75S2zRxO+K9gzNzilQxO3HJSmXe9Qa2
orN8iTkXEbSwKUI5rrl2sjl/2Tgj20noQ7xjEO7kh3TbyOAAUdpNpJrsWe1FivDr4GzWuOkS1L06
YY+TTGa91q7IlZKc1+ZhwbF65rk9qlzMNRb1+jgmJMYo6p+ElNmKzNx1fARfMRZpTSi8G8lC8lsd
SxO8X3DhxbVqgxBc+XpdORYcAF7KevsJHSw96N7+9AGfDpXQqiRrzfVS0HvuoYo5tmBmOxMiUZFz
SWBnxp1ojCzJk4GJ0IufJ57fjOBpibS6z9QODiyMJBhp0eSjHUh91Qa7rnV173yTJ3fsP3dkEQmX
JBYjjC0yau1AwrptUnH5oVAsYWS2vMhh4RAJq/ymAoK4WAybXojttxbcTogp9WwzTfrvSljNQePz
TGRGhjwwHv0cFyA/Syc8SENnpSiVqkUIHrS5tccSpsUmQKAdEsxjlpugUSRIdCgz22Sw2/3boTM4
dmLqh2PY5xtWZ5DntNG1THHpmPj85BAWvyBqFMJwpQCa1vabHrPT5GGodUJOz3NW99p35ldoyRkm
Y9thzTmlKuCszqCk8BhdLk45+czhZn/zTIu7eJlLS2DdnBGlHljaPhB5wxOYL9eFjxGH1P1JTRit
FNhNTbqfw5bHlb4MsUbR/5CsVXqtrNCtzAYovOVNY2abL6u3X5O4BCB2p2Koy86XfqTsb5JqBE+2
YhCT9n8q+Hf4N+NV8tPyF3El6BEfrMRznwcyhlihCH+fLPCzAztyxGPkpO59OVoSLQKR4mXzu6GZ
uosIQdHGozbmT1KlO2FVypCqkdDDO0b/xrg8ateUlztHIAeU8eqHQCpZDWvxpiUpZGIa0MEKcIEl
anhgh1SX6dP19eLobI+jgl6+FFPAGl9PM7bi1VjwWJ+yIQUaaK0RYniKpnvUdBysvnDNOzaEZQ5d
99B5bARWjzde3v9x1/kQoey4L4UduMTlEBZL9atjqOcQEXxrUWaHMV0CPOidwVyFXXCWaca0Yg7D
eu+JyJLYRW3Nz7+NsWoo6JHZKfyzNWOPlL/z9hl6AXo+JPDpdyI2CNNvSdJT5Jj7KcoWO/MhOGoh
fqiuf0fuQGUFa/XH7d+BG7LjU1/c5bfE33AcmL0Iig6NKo2fEA4u40CtwDzt1nG0Ez+/NcQfyxrn
dD8wzNGdhyjTCf7Hbetuj+UITkbi/nNRCr4I/C+xbLRW2vZtUwJ6xUYAdcMPBTInI+ITxQVymi0h
NVGOgEfX9rSHSXRqQNdESz8rlhUmt9MRYMpdYfMbHbVpowQg8ydywOA6zBHCbUmHbc5AJkUQI6qk
hebDUlSFyH6oAQ0z/KxlR05fyr3bnXWiNXyZIxHdbAEm1j7smwde2iMks585QFEU0x2lFXlKPvLC
3QCNMhe5NkhgIcaFET3mvv+DmX1TBEP3f4KyuVsKUtYWV0aPWFn7ISrJE9GDmc1V1+IrrIBhevfM
HCP5iQxcczSMg5ksyewdIydhIHk9B3ACys9seExRlQYUFHCp3Fwcpn73F/1TjxGQ6GpPinPt3yD7
AMy3hyWme2NhJf9tkFHr+9ets2hYDA5RQPa/cuhQpdHIHfHiK2WhXRHDnrZ8Hp1yLd7W1Ah6CEbF
lo+LCkzNQw/e0KN7Jr/BdEObQsA5zjOveH3ziTyHg3ZMgQGCeUgJPTyOeyJL+mvXrPTSCMAL71eS
4l6dMyFLWTATpowSiDjIUI7aNOcW6IlpaBcCL9YN7v5M83qvbScJCPDJgBE7EP12VGYCw7f1j6/E
IWYnKqcY+OyiwqOi81ls6DFkhPPCDt5KWN1fg3rY9xeIi5IvOWd6EAXuz6eE749ZM6a8Bpb4uyj9
UpLw71EkiXA7fRXPESOJlac5/Lq5+J4F9f4qM0r9uses6n9DrlQfYg90cCJHIq5szIdZTka3XkSb
/fHIgk6dYf4NcJJE1VdKoY/VB0oXAnPiz/1BX+ZxJfCIQynqUkYBmUPJRbgtpxo0SCbMxA9cm6mF
69f5p16F73V6Y/6mebQTMKhKSG3GT/3fH4Cc5dj6jCGzkEliZzF/euzjzkv3VJcj7TP15c9CYWSZ
NlrUkCNV0BzkY6x701u5vkqdusi5MFcUfPf8Q3h/ZmRf3yFdRj8TrPmc0Ju4nvpX3AOzpXD4nVz5
3OHrqIn7I9nKUIR56AuKR0xWMea2Dq7qjD5T9G5s8WTzUx1+DMrYb2j7FFv5llmz1ibSh6Rm2ClH
CdMb+jldZ64YFbQRg2Ud+s25ec7UzA8wANhr6yV5o2fzs92tsgCm6nSxeCO/QkuwLCeuD/gP3ZMb
OiDD8jzCNH81/X9J/HKOsXHp2NXRm/6QmodukU8s7gZXDS7PZrsnXIO8/rAaEQhE+BX1AlxfZUk8
1Ul1vT/1+Qa5JWq8+wEAGG1aAmRUWUxak7kV0ELhuYI/tXL/JPauhNq6Nje0bekuh7tfsWX+C9Ve
p+Fqad58ed1tNsFOnXIkvDyc28qZC+7RHRnyedI2TxAjPPKtgebdfn36SJCNrSCMi8JsLCo1uENe
n39uiXkqposXlTJedOQhM0qX6Tz0MkEanZh4FvZWGFCJAHYcSxGb0iRBKzRbs8P7Y/p6Nb9xlAcw
k5NYSxeNvN7cUcB9iLIEMFytvq75pZD2O841fWbgLG1VokYjOLiNHoOBVLZm+nMQWP25YbikjMnJ
Nd/662GFTe+8Rnq3Tx5rM1Jthi48ixDbAA7yyrkCbT/UTeDKLgxwJzHQZzJ2x7PCBSpyh87KELgG
YFA1ZjrDE75n8QGTpzYBoMMu+ug1SxAZANrKIMcGbEYKzNjEc91A/4AxuetY4/2LReTloyIpVz7p
QbrqNGgtWZgQvXl1JJhTUd9ZPo1Cj0BVi9DNBJ9Dq+oNeEMVaBIy6JheRCDVA7B4c8HHsNMnWhjP
c/oVjrGwks5DnEjF1k2EeUVQTmBghvGD9WZ2hba/Vdbh9UvnJS/zRuDN7blZgzWweGia+dgbeYVs
fxJ25zc2G7AwrLMAn0d8RcOXP7Wa8A7Zn8RXeOfeSEk1e1gtTBCEFw/zw1JSrisWFKVqzSya2245
ZVANjB9+AyiPkdnjWVKHrXRNJB+GsudVv/wEdkLx9IBZQ8Mlcan7xDKkzxhKJbmrtn80TFKPBUVY
NAgtBFN+iy1/3YR5rA4JG9wtrkE9Bf0HC0/iJahTyCVVGBE05EOWF08MRxAnguN1D4osL1aI+8v3
gPgQmnKIBSBxFzbDu2r8E8ER6/xjjv5XjGEybjzkI0AZ8+9FdG+gUeFW8Hp5iNDiTBviAHH/fwat
iXtYdF6KIpq5yjqApb4QBPvbHVsZcyH8JHZdas/cJeNAf93GkylnJZ9CztPVx6Ka1g79QSPqv6pt
ylUtOPVEAXvlmB/xQEPlwX3RZxc6lp9GhSjO4U0pqMKKOd9CeiNTLxiWXJREh5EAjrPXJaifetDq
N92HRXlboecMsvxFVxm/Ax3XdUzTX3v+MNqsoNqt3224LtI7cHhrDdd1e9s7Lmb3Dt6lpTPujVne
1gP/SsnaHME04oJFdHzm2D/Rh5X44azaEWG61R7ItUeDPHD1291sEHfKSzfJZIEB8Sp5QWZOTQGm
Ty8EI5iSk3ZNOaCTOeSBRBFcVi13uD+7f8yaQRgGCTFg9jymPFOBjQhsRxjAN7Ce/9YyrGk199Yt
rtEYZZQIylTIAz9AQM/uJRuyG50tXa5DePjAbCtzxXYkQHPzRmte4XWdL7JFxUXDMi+AsDGr9qPY
i4H2VnWYlg/rRF00CASB/JLXqaJlJp0ADXHokLDkHzgLrozDmA2V4cxsSR6/+bdnuMq/UVIvKssc
HHEGitsNV1R4jgBggtWG0LJKqHrp+r+HJyLi+DnjulYGBQi7CbMswyttqiv34mk0s/NkR7StKhzH
RHep6+vlCzdX0ZuU/tNTsv1xj5NTH0+KN4GgYLrqYw6x69ejlmfM+9rT4+DAiuvmbWMtGM+RFzjq
eFAPwRXbKrCDVJbpXoh52madoflnOmtrixB/PqehDGBc0Mb3U076GqH0SkW9d2XnzCfCWMfo9ZYA
94HvG+1baWUbCguMz8eOfzBhIsHwXI1ixdcC2MHfXsQ6Z9yGq7pPFPTvi44G0884ce1xcq2fCqIa
B0lyeo0CKsI7Xp2J8GwQYlwU5kUpteldP371gt5+bp76BRmRz+3pnHg4gLl8659CRfvD6/fhTmD7
lwi6gLNlehl/tTTAW5Vg9wvurCUcY/3nU/OPPbOprybYfySykEMSYAExM1AbEps+USxSnsEVWosj
RinUvxSYz+ObQihCL8ZPRqnfK1+tUamz9j0xL3mIoZ46BDpOH+HrlqtbpFpiIsF7aL/y6WBgLKrL
CdL+I5eQZ8EDsTlfuY206EOgOCHiKsb/1QEhX/1q6qRtc8AwYy3e9Jx4J95mghYFgOc4Ojrwx5KH
7cqRgAuvmIXc2LDfvvIwNLqsWI5bpZeLX5gIxXyOZQbC3Ehc+KtQUi1bSSJQ8pWNqStSXA5E6Kdp
GAcyXXKSu7H11o6exRcFEH8dHROOpCGR0K9msvKG57gJLPKS4bjsYKFFsHg1M1jTYZZ35yKQp+F7
dHGIN+1JBmBiKTQafswklLs7gS1WzATQm7o5YNwfO4B/8k7toNdXiVZkEzKY+WrdIgwKkRE3kfla
RQRwMO0+LDeoUL1Ff6MlD4gotxjXp8mbq1bNRXGUuCqiAYX6id5drlWvzmCOhZobOqg9BsWGIuDJ
zM7FnO6CIGGopx7SYR3mruytLM0/S3sIC5AtCtIsCIuRUk3UYaqjzqFtDsMewTAUxKGFgLARpygG
wZ1cXrj2azBFd0kCFt6XOiO9ca2wPhxLioUUaOQkZ5SINhX5dQ/QZ1bNnp9QBwPwUaLrr45uLW6j
XNBbPLJ4SJg6Md+feD1eCaMRG0X5++toftst9drMtfQQTl79MsmUr2XAnbIHv3n6Vi+ohSSRa4nA
CV6k5JdiLgncmEy509cfdmwKq28nH5J6FRzf90tHu0zGJdAhXc7HvQ6MHXYDqeuL5nmK/p8B5U13
Qx6K3RKjrMo1oYLvRwHsmj+MvgTuVIV3T0B/krOOPu+kRbeCdg1lerWl15T5C4zfD02TCQ+DPTs+
PMB6g7P/SpLEAWvWOckodg41HY6nSpKdXGyB9bhgipj11KqXgdMhhNwcN4en/SFFcSv/DwmRb6uP
uC2btMiynNkLXHdH67vZvCtT3z5e5dGfxnys4f61Z1lcBjJoCUSfEfENRiyzE8J/ZWA/IEqw6AfG
HgyHRgzaiWdMTacdl+xT7muffg/u+gmgZ8+Xzl3ooV7wqXPJVpL9SeGo5kCZyT71lmX864VrSfhr
V9Va2I2yxcRbuN4KlyxFgHmH6IhlnNbIyvJs06yutG03/fcBc907TfIUvkCsRVo+1hs4f2AuidTH
ZCwlg+FBHAS8zLvy4+KbwCd8jJF+bfQ7ytbbDcy9AdPmP6S+eAZHbYKWezD7rUfQ2XM++qeS9aJE
3RezChFowtKTe1F6FQoWCBtFAeU/OfcfkRzqX8MK8M5DhqdToUT/x9tU4HwOG+Rd1xIV+ejxbumh
2w/tOd9bwmc8IGNKKbrmaczPLiV0KBqIVkrdEZeMFIC4rBH2EVmbSnOAklxpt++dOVy4LiDNrTYe
Lwd7YBltEWLaflWJNe7I8D5svByBt1zxMw5JpJjXx3yCpXMZMDj2d10Qdmw+2VGMkaP2R4msV9co
PSV8rZ+1/v2OGPY6oCyJ0q9KDh44+t+4+he9DC7HQiEAozZqmdzsVduM8+q5BPJacFXvkBQtkGIB
vGb2VX7zhRzxsZQfAPVeRMjuowWXcQyGWyPjb3fXQ5tgg5+JafOUMYfcyMFmlbTkvN+6p7gD8X+u
KnxLIVcukV65Uw1Ko63QlF7Bry0MlPoKQyuxHt4KynIp+MpVJiLGKkNVNxgahONLI/Kzgc023Mor
lqhO8hb+qe8OIuUKudqcJ6j213VZF6iwJPEMFHvc8aBU2CRn7mnQoUNSbC7iOx0z/ouRFUaxrOeo
Om75xIN8z3yjoZqBs9TjqIxaZJKNo3hGsNCjwMiQI1tT2Lr5n7kamEEO9HWD/RISZndsLAuStXAG
brWEjEQbD18jJ9FoTdEcwk6q/3vAUaz+rZBWo+WTrYbW4tSAGVWK4OJ9Jr+JNfNhKPHzgUQgVpDO
SZaHiEFkB5e6YrT8msWL0+YZKsG9WSww3pcdR+Uy+r535GX246w2bLmoAhw6mCEWteqOYbCz6Yel
NxAxBJZ4zHxb5eURL1azxIivHhDbAIgqbEVkdfMhFqhqpXAqNhWhm5kzE+KdFsvK0x7nAi61jtBl
bN3cdBavB61A5SegY6TUQPiM6hmMu4/oNGaVnLv45y8JRRU/9YBf5406AjBIpxvbkAygIN2aQpvX
Sfr79aCrRQY3bow0kAYSco2YkOajwH/7SWIdzDQSXOD77nmmqMa6SjmaecZ9zdnT8WdNytVzLrvA
ti/VYgvVYCZvMgJoKgiOQy8WVokRe/HuMIFQtG4cP6jttGg9iqgkmeX7Jii/ZzCggYxlGkrc5rVT
68jQO/ixDLm08w62CssisCSx06jS+Ft1nVnpR4M3SYRBWbytWxgPZ7jnAAQkClD5ZrcI7WebC0YR
xAYIget74UCQNY89F7v9TprmPWJCReFS3sGqWmHR7PsCLl9uKB7ZtdPe2fzN0hnwxz5gDB+93K4X
/53JUOGfrnyL+OKeGrvBJ/Es/IJ/bQy3kZlb77m0iNWiX4IX1oJoGUdgrEZqrf83EzmFjX75PIz6
oVEA7Ntu7nqk/EJ2Zwj05w8N+yBPfQoyXlDFbDiMe2wDw7kKyvNXBHBweN7MWupqTBijsgbD6E7e
jwabvKSFJEV46AjVCLwzsGc/GKBZIdRb/rzLElKk3exdJoBov7yfd2geq5m5wSJZCo+V9VJY2Nqz
dWigVcKmhScmPwIpa1iGqQxsbDQrzwAKsCwzUszs5MAlGV6oIWkwvEhYohmCU3Toy1ZAjsKTGl87
REcH/b7LxVnr0iVpAQY2m1O0CeBmvKTRjfpa/g4Vz2pmjtTSu7l0OVpge7zIJOTtnSSDvkIMYxxy
fEw6zKKW1gwHTlAj9pQOyx+tNrlpKSLkSq89SBlRQuJz7DCW7ExoI6xdN860o6j1kKAz+p6NwdRZ
sbtwGo8XnBeIzy9oOpQGS/anBUuI5/BvcwR3QSZS4hGnbR3eHEoGs1yjR5WSjGdVK9DLs+ySZxh1
T2qsTPWM8C5bhlgWnZpEwP9GM6YLeE+LmWlRogjMVYk1yc/WQ02MKD1vW7pE5JLPYPxeRFyUCcZU
W0GJD+GBUJFPcEt/KsyOTTiScfoa0IV2OxXHNxepSktqx4oesdVykWt22RO99l1Phc0bWkEk3CsX
dOyYJAB+eka/k5OoJEJ85253YuoB5BaBBDtFKqGcO8eeg6c8NaPpB5YH9ixzsJt85lprnuDPXHgR
P+sGdgvkjUEhbhGHHIaHTXaOi9WNF+hYXO7CGZ8l94W2B2yv2kdXTAmKFd1RvScP/saEFJEDifyj
P4QI+z4Av05aaTledOHf8wJWcA5xuLeZWEKxxo9phLvRcs6yevIM/1RaomPjrWVR0R7W7NzuUB7B
cfK6n7XgytCh7SCZlfkQNHQHOkdc8g+IK2fn5TdCjdFxVSysgurvgLIsgolDegxa4nKcPngN+9vV
1D+7VgALvq6Gwa5Bgv+Ss39dCSKqM2EPPjlWkDDlMMiRbl7EtiY/F+q64eSKchDSThjTWIpMzgBY
djgFlp+9pzpxvaNNln0KbKavhH0E01HXuEfapKyQDkELpR99fGkIyCk0a7jk6S2J4j8c13rqSxPp
ibMuXwBfhN9qoIzQ8TnccGHrDbohTXWgt9NUHH4tXI/0Hnx+naI0Mz3RAi2K3hRJxBTJ+giv5bns
GnEOnCqaUePk0vLLwXYQwGCvnnJzUcwRluKnUFCeXRA/rNSY6HXsaK6t2lvwRXsXHFtesB8a4VZX
FPgMvu0oKVtCc/J+b14xwuo733B8XbAgMZ7MVJcKnSbdCKYn37lCtUZ26HHkJjdp0D5z9RJ4KbO3
nsBGvIAdn6mvwnr4uUSRKgVGDNpm2uBl6vIeiVrFxfu0d90pJ67VS5SfhvWrM53BIMGmMlwRWNJD
WDK9L4Mnf5+RfrBrVNEHOkLsy7j0Lik24HJQiq8Mnmcj5kmnDBHcXXjlL163mXCZ5ZHOrtbAqnuZ
uFF6rB+1/LnTgPOjQb83JsdR8PXdDs9Jnw6vaeB37vlTafR5dhHsq6TOHmnH7pe8+ynDxXyfPZ5i
SyT1EiOrdYjY8jko2TGLbxvPTnsf3LsmeYlfTRmoxy2txH025V3O9n46zg6N63WvPLYnT4L+s8fL
4kMUsL6u9/6tV1jeTo8hrpaUsj/63kYQLvFbvV1ACKKbkRwXxlN+zFIBeh4S3k5/cQRLyhZKDBSc
7XHfndjro76RSnVs5JjCKYfFP7Et6A5SNyNwkHmnhmLlxpivo+XzSrojQFUHIIMrhLoMvCMaKiLX
T+q4TmEU+fBKVm6o/WU8ahlvJt5iNClpwrm57x6zWqH9ujYSL+WoNJu6pVDnvoDJqXibTnSUMeUW
xsJhCsSzbwWXmp2wKo2qInS5RgpSEcfUHH3ZO3SJ6AJRJI8D9XmYH0pJR463+Vx7H1TV7yJgw1CE
AHFDJl0xKr1msq4+ZurHx3U9pTmx487VNI/SSJGhNISEOOki8zaO6iZo0ARJYEZ8J++c0pkU8mCw
zE2VgXzJdbK/Ep8CVL/DOAJRdnMhD4j3rRT22MHFi3JmUY6CVcI4rZ5Y5NEQ52GpMa4ZsGUydysT
+hvJ+fJNo4nOhej1vrKmXHpEdtYYYDE5o3g80caBmmXH1hFTWcTHT/qTeqkmVSWnt7J6D73fQhKf
e8l5pQSgvWiXq/sZcnPL/iCnz1DFksNZIa3Cjyjr5LKeB3PTm3jrrczxddi82iEPB2M6Ud0LuyJU
Y5tAiay1xGtSAKESi3IhA05U/WdMI0h460E/jXO8TmRtnfBnRWE7iFD4kGDfleHlABODfWGKEttz
uyykpSLW2Ci4xDqu6uKlm+jP5CqMFjvKVsEwqEn6g20tqm38wZ6gzWJhhg9pawPWL3sT1ZzOW0we
nC78ZI95NcGzzf3NE4jdFQglGBtnBMqUiwpTZRsxf0/TFTx/yYtuyAqu7b9bIZgBd+lYICB7JOT7
TxXeSKt9a82YQxzkjv4MMssIdAmSoB7AFOuA/Zspks35R8TVlxkOzL3p0JPqp8Ru9IlcIErksBXu
+nGgKuP4ro7uXlGnLvfw6tGow4V57G/w4pkYzGoenDPA8QtEgWH0hQjHkOIAcRb0itIaHKgu0kxB
F+p646ahbJvbq1DrNTUqEIvwOlLv7hXmXRMRVq/NPFylC51TmN1TahoTHMVtrrNIJGz0GvS6BN64
JO+NxaG2KkscASQ70jOkcTgMO/0NhtNn0pXwXFeFLG0BP+rIXplbHLGxwe+0lmdmPn6FkKWb0x+/
lWsSEgxMxtpHlSEh5zjvlMApUkr8qV4q6UknoPh2yF5Jf509fCsLsYTl9SPu0QKNKatZr091XM0d
u81Y6oa1Y1y9mCMEoDiE2WHgHSaUANl03gLjK++yjGpB9lk7vrOljLHMql+irNInh2iU3Vyuz9l2
ymOJVjDFYE0EfbZQAr+OQNNLxaGknKUoIr2NK2umX4kNdcro9TXpAjhJWRMC0JQ7JuGv95lASjWI
/kMx45gUQFQXThc7FhhXXDOowdwz5N4AsrBc/EG586eNRvrOvpZuDq/3mp/sVJ5BP8b6OvZmfKaI
I6jyeaV6fbtTUdDtaohgTjMXFnoKgijZHcvZEJ4dHDsDlT9VpFB1qUl/DnLfYlyKyFdGSD4F5y/D
WUu9+sFev0FnAKkfOTEHzyK2au9HSz5Mofxu22A3o1tVt76MQzMvxA4h2ksxTklPgSj7966dtB1U
8e0uaZmqu7v4eDaCo55UvD0nSLgiTFj4Ujttvaks1LToXEo9gTJjrqEcqYU7jBlmlF0lfdJeiVI5
EJOZuB0E2u2EcUIDebUuuALNxQLJfNUVVEtcsL8U0RIZ483NlzIK4n6x1OQSYBT+uE6ODvu4uHK1
6ppTZ72q1hl5GGEtg0JZuqJ7HUpPXJLXPLYivFxfeOME9s3YIMAI2PTf9EPeXsu4gGeNhoHPXcjk
7BrMgSIz/9FbPTHv/NKQm43kSojPvbgI5jeVDooSrKHipeJENoNsmeFImvZmY9pCfpXpkjqNPaWn
vwYE9ZR141rdspdp7g77w6qhJ7TYDj84M2y/2M97/yZIXJhvzgaotPNEqsTxH7lCIvZSC/o70tVS
Zcx6OHZ4qoV6oIuYraxiAmMhJAcsNhcvjjogWAfdFgMjyAAVvrkYrPlSWv/1uUxZ+jT0tBKUJx6y
lhM5qS2lQVgVE0KLoAnywMcYg/dWTMJ33IWQf8T7mKmi1GOtP6Lx+XAWvFOBar7W/Tb9Mezzk4xc
OM2losTZkqqpTNmw2mzPy2rbO8g3zCtpSBFYnJiDJe1SZtM3MutRx8f8qRIW/WRj9ehqBiTzXfkZ
r7vnMTRD+K1hO+pjAPMtnQvpc4Zsb92fkNKTo+NtGX82Y5CyUBZjWnJSuoQvJ0QY6kF+Q1RoREN1
gS96IFsJ/pAL9tatan5JQIt3I4oUg1JSoET0smVTKOyzW0kwxX6GuVkTocuiXxrTA1xWTB+dnSgS
6zTkJp9fbINPsk1xw3phj6nKRTgws7cGJx4bnExblKlI5GWujF7dqMpbDMk4YDZN0DAMQUSaQWJd
WyDCqFCzNf6MgW4cwgzLrlMbbJHVL8ITdM9jaPof94P1fALAuAimVgBLDPP7DRtVneqPOPV61r74
xKxtxFssx95P+IjkAR63PO9HgqCTCvyhz7RXGlP5Gng1WS1JV/HvAHiXygyx71ooAwg6gdP3FkYH
IUJnyqJbeSom/M9Agqogeqh7TzR6EA3824DDS/K9IOw09lXUtD5bsH0bAlC4SgHLYdhyyRvHkYzC
fl2hYdb8cw0y94fp4yatpMPv4LGUkjV1pyoih7wtjHUGhH/k4pgTkG2I1+W1iy3RX9Yw4bc4UID+
ZDvtsLWo5maei8TSWI/ZnMdhacQKTuDlBmmHP3MDY35f76Oxd/8o8N4cwohGKVdzcPZjDYTIGcrW
f4uZnskDbtuSgtcOeQ3ENo2Cd4nQ+KgqarqSEBwX/qKn/GQ6uiGvzsaL1OkfaVPLw2gj8klUPh4C
hdG3bSj6G0hKj33cu39ARzwR9gUbK9w0HY0hd6VGEbRpiuyDEyKiQyfbN8qa5jgbdj2lJpNnz5nW
z+xYl/553UFmLsYbLfAXQ+lixy+0zRG/0RrZkxTwH1qSpkmvaDwqiYUqpeIO1+XX6TR25GVwNIJr
V+t+8A7rZxs9u4xPvmPGw9/1sGxaB04YE2TDJbwfq3bBQ4sS/qy5iTqQier8ucr7LijQdkVYF3qn
knwncyDbhGPpUq7dw1PD7G1/LbUsuf1NZNCYm4uMmSEHE+y6cVtggbInZ/Ceik2MdM8qvtOPKPHk
gALjSklHLIkLktwrXx7ik5V6C0jX+sB7ISyszjoz63Bnmg2ZzXPTw4+uuBWMIIu3pkhFFrHblz2z
nrjeKi3YKAFpEPduXJUld10kIJM9ayME6yhYpjbwKHkBpjnCScUPPcDZioGZ0TKg/PqpW3Em98Ll
TwKuaJ2s8jKSnI0rTxUnyYM668mswtPwpb6rMZNzsZZOP6m9NGTmqR3MtCy2pC5eFletq+cyfl2L
vOkedeyGtOfosscw3jbQkN2cculkvmozdLNktkuF2C/2gUYM1Lw871q1+JH9FmeoHccB/R6GBVwD
e/3adi1A+njre2yOrHus7JCDG3AJ58JsVyPIThJ83rznB4rzblupHgjfJVsj3wqGhbmYEGQ+ZFcs
HX+RdvojrOKYKFMurQuj2q2DhfFYG/F/sJQ1A+8GtUYctg673s2ZhFvhSxs0IZAZJmtm5IPG9HK6
CyKgNRGK8c88DAN9jD/JoE8/a9SZP9VczkFrO7YkByvOJZESTlzD67kILNeD+ezYgwG5JE+Zre7u
i/mIsJixV5wNKndqyg45IBQGL1PkS0Q3Km3D7efcrJtzMNptrr8juNhmineYpKMnEIKYol/ZtdTw
xrI5ZBW7Bxdy7wDtrdZam7jibADBHMLMFwcppfQWXn+XnhtzE0yxRdp2dzRjat3mrP0X6UJ8J4cW
3CWa9AmwnPw+iYWfECRCgOqfgPrKZbkJzLjUVIvhJDHIhPJgBsYZtuaA6nVUDTD9lQCwFaQZKdaO
wn+Rtj9XE6i/yE6DGjw3Lae4LP3NxHZD7c/G6/rf+2dNX3mcxfDCyHZo23tX7LLyrZ3b5P4QYAcu
kxnrSfJKeE40vJy9bOj2TQYcrPpkErVgF8LNnbl4P62P7s31vQAJhzWJNPJcQqrtnFK0QmDkQDDx
EWHKQe96b+M+dxgpSLdHDNEJwum896TpzD8//mMGfhvKQ9kuGb8pq2Lq0Z6bmvMGRd5VIiFGzkaf
JxLWHdzb2zEB4L+KLvIVVSc/YnIx8apcB1Z2cst2zVwQ8N9VaiRvjs+127PEFKA9cyPWv+SuHCkS
fMXoTGlR9JaXebgmEI5/VfL/4a2TsxHH0nRFn3wPMmq2pyfIsE2xcLc/PwOfqlWEHPkdygaN3+8R
Wk94dm1wbSgMW+dsYK+w4entinrfWP++q6KYmK42iainc3Vdd9PBgjxN1Y6k2mvch88HAJVlyIlq
7oyqk7H4CzizIv51I8EVWflI19z126S2QsYatMoHg+tKbBDPHMI/yV011NHu1Nfq7HH+m49N/AnO
rnm8SQbc1NOSQFcU9rWSLOj/jkY1qMsq76Yxjsr0tWGkDwYxwu0fGoOKg49NEAyBm+AwnUU9STmx
k++P9Ch1Q70afOF7dSozccIHZ35II6bE5U/+YVsp542DXlLFq2sWdvZS/IlofyI1RymeZkSdBF17
181VuvY956FgO2Xbtb1AKJBhS3vKyruxoMZ1gLN3ZbyO6leP27D4qDjhnAI1RYJlvc9BpFmPhdAq
GPpwMB9ye0GeYRWMie2oLABrzF3MK6xDyFdXzpZcKnyfjP2Rxpntyg6u+xTXLnzkUTD5119311Ho
9fT6GfqiLgOsfCU9EA0ImdAk5NonH/h22bw9UfdiF1wu1IdxfIv65m9AZYXvp8Iuo4Q6PPX/C2cT
kKzbR23OiQozmeKhNg5eIXDW59yzQ3NT+zDuV4xp30hWeks5DubVet9U9Y9FC9RTA+ZOosxilg4A
Z54GZf/iGCADHWiaqnHgLAWbaH+cYJNbLBaL/ti0l6sxw+ON5pmwdvQQfYXTSll3iRp4hbYcTqyK
BEQiN+HaouN4mmjOjau71LNX/XdnDsJVj49DLEghii0+P15fYrcI6s0iEhHEDcWg0sYlhbD7+k7E
J3sRZ94qkyFNXczDb1S9j62UMcloukg1QTWMSysNB0Bs3BXCN5EfEpkrdaeKhQMHO3GEJ9iFwhXV
9I5nGYCSsjKK5bvQOyJQOTB4iGuQECkFLL1rmHnTUobX6TC5vD5I5s9FrXdkzORECipQDMoMvI6n
YR8r4wkQcwb1mMAPvVYM8gwhL0ldIP5OuD64MO7vs2WLQZLICxYhIDMEo1GiwdVS6AjcoZqMXkDx
TqYLzkMkAfJ9isYWxZSWGsbQA2VXh5HyUOydMThbIUwMSF22XQDBRiLNO7SZ1goZlnXHZFaSCNFd
KK+jINDCroLNyuL93AL3rqOKUkR8X/DVRMvDJlx15hFnxrghR/I0lQkVIMW/ngGQFC+MhSQKPj62
gBQMx1bgSs5UID2kN36Fh1/9Hd9NMDkM8xJ5eXES+dGvOBrl52BmajRHYkpwgf7qcSaL1jHC2bM5
3w9q6Zxu4Dk3Y1Uuij3RVJncxFkZPxsr0FJ5P8PRtY+UVkKAnm5Y08GDu/qAcK/IYZzdIpm0gTg+
QXWilC0ykH1mwSYl95g5J0mJlQ04rDHsrc9zyFowyv5R7YzrzOkFOZ6rrVVletgFCX/aTBiKrTDC
PLW1GIiBKFyZfqTEbb60GqFPFER6EPI6O6JcujAmGRYEtcrMG+tdhuFNFGBqH1ner0rFRyB4J7CB
hkLQIOuaHBQelw1kBhglpCzwLlMV1SF4SmhGaOkkGM5JjrlDqk7OVJG9jL79IElUN5AAPniPNiTo
aZTgFYHfwAlI4BkcgVca7xK3VHCHN/SQhGIirUlHne1fiNVC4+9+rO53m/cyC1jI4lIziGZl1OCa
5HrHHURVhTfHa5gZoAYryy68IXCKYhQDiSfQUhepvgZIYP3mM3mlo2vsU23pMPJ3T4LbgZn73MLX
O+Du9CFdIS7kYhIMX24eKKj+rqVw0I5ZY7UbGxaETUEeKiWyYCCXBx3V5dZClJof+OTl43f4s+x0
KgJsqXkVToacQuUEBA4yEH4YfRgEMJ7qWguzhDNmQ6lej14NkqFg+QTOB5GRTm0++DVNDpRagIHh
FLg+0VgufCHfmJux7egZP1SuYGWnXYr40KE9OHCsJWWozBZc6mdSXCOqy+DysOBrSTaZ9uOBl2qI
bp8mNPT1nbOrm+Svn50ejjdvxdapXCGUJ/TijQlB1ZtnGp6NaZ9uBzE9Bt2M4qksbIhFSRS2oi7S
lqucOp/gEWY9U2kaKYho5Z31fQiPFk9aMEiRNtYtR8D4iFtmVuQCdzkctP1DHoomqeosdJZM+IjK
VKpFfJkI9WPQdNngLoFb4pE62P2YGjiP3SSyDsIHusc/OFzT8nAE3VMmXNxfc8yk6dl2ER08MRWb
xFqJE/Ft61odjPw+HeKMpi7kkUPQURBNSs1EY7S0VRWjuf3v+tn8skCYlyjMlJC7MWJwf85LVZzc
etT5/gql/qTZ7N0w+5GRUouTIua187ODqXazIbq0JNR3pyCfe1Ml5WnMJTiVwYASSAk4q4H94y6M
kYGur0WfvT+yNazB20mv3bF5la/T0oZhQFFudqoe2yXHfe6UhMex5OCP6ywClV+XU+bj0RUZO01/
69HbuVSHjBxusZ5rlqalDoD4Mnz/75TySSeP5wPznWoUv+2xh6uYBeS2k4EufuQvXXeIYvskS0ZT
j/Hd7BAskz0LdLWckd/2qBwLZ8+KQHkVz50QzcpZYSM6TQM4lJpJwwMDyYR8/faK+iwExxY1mije
Xt6ilrrbkMPPf71Y119V+bKUIH+k8yt6w0OP6EGXmcoNa7fpOR2qAp81zpbTDWKSb4lyUV4vAceJ
/mSqDNcVMTKGi77crY4+Jll8NZol3+T/tDDPauE9719IxpZJG99ZxMEiC1hlWx+chcwAemfXXnt8
I29ieGk1cBDFJdKJfhNA67W1Moe9U7/GBnZM8k69J+PRaoIXPZF/Bq0Fw/pyOhnCZP/MMeDFO3WS
oMhMFjxRWp5LHnbr8KGKVl4irbZmpXkZfCwzjA0IDZLUZR3zY/esC0zBnChHQ63693LbsrGJ9xwy
ZlllWZf8pR/efJPFh7ESAWjwVaezt/WKskVcS1lEpYehre8Tn7/FAWpny1jeXpS9uM5tlnygThdj
d5ttzK4+b46PyBuN5DkHAQJKP1IOIJeciOxs4Ch04FK1SzEW2naIYpdXXXwopjQkR+akL6NW6FvE
mGvy8IODuA5bFLpvGUfAIwWDAZe/UnSMMwiWOK3c6c7xWb0mg++fvcKJglznh4cW1JwzWSGfrj6O
O4l/c0OZLYTvc0lrwR9L2YbAoc1sfwnZplq3l/FAh/1rXybPZmSLFnH2qfIcxgPyKXFb+TOyHTZq
DMuvDGhpMizZ3zPflQLY4jjPKzoQVW3B54yge3t8uKFwSVEiQ84ORqSGphrAjGBs636tA9WF5Z9I
g+HxHQNvYrr4gxYrRg1iyO01u1EawWCgwfwhTAblKkXXx3WWKQHz2gJdvepj95PGib3oJYlyeh/N
hPOELda9JQRQZkFTD4jvtcAZfL30ak2uy8i3NSVTNOrzay1nFXWTzBocVfmM3FiTDVk5AaJxmMcT
Te0VXHt1ZNIEOvvAFoXn6iEJKbD4kBaIgaj+D4rutjw9ZdN/kNCvcjBQUCR63jpiMDNUQsGLRAC6
fpoC931oOh8muZyxIyZzPRmlygGq/USkApfO89jgH8WnQmOP8CRKneiLuvLeR7fuUX+/UU42Ks12
hxsro4XtJaz+gpAwedsMuJU5d1oThWev6M71J45Ali97dl7mC/Zzv2d5XzJLx17NwqwZ9haZb08J
kiDqxatL7bGuPXQn/xlGT+TKelVpExB5qiiura//Ja858qlmvL0gTuGacJcxWP3eiOaM9ZerC0xN
z4DZYLyTvwUEXCSBC5a3XQPf+ZtHT7+r1ssGKmNgihl7GXtpxMrvDYc8RPqp9XsK4GMr3l0I3tYt
8efAffPEA2U5rc5bdbyuYQzu5LhQ4jOcvNzZAo4R4KZ1bgl9X2ACUHnyxw17Z5TZTWUEAB295Hde
PxAAWlJD5G0umKrUmE52i83ufvCBG11/LofsYOuIcqrXISuVysiuzjrI+lvNLYCGlje6HllU4WJK
WSsvhHpKvYw7yFeKUQPq8ua820BFajY6by8bI5e3hwW0V1i264i7sduU9kbmGy+h7OBoKWVAZX5W
ZAzJKvOgrVNQVCU+Ulx6j2F456O7bUySBgwMqn/8xa+bB/Cc60uefFocrZFOKuvwitIr4kaYvOH/
oIIgWXIgoY4cm9qJzDXyphj81wIQ7E1rYkr1busFboEfDK9lIUFH2LSnRaQysskgyMmIIfN2xiWn
maEg3qDoJqLbdNnRTTa0JkzuI6LgMhjSKuF0NtQTCdF3h2fZODetSXma2Gywoh2GtObRedt3IavS
dcHA1DOTsTSO9gk14RzHntIAJhzCGBai0FKOeZLEPYu5RArWDhG56Zi9Eu1SslJHGcaZYEckQOCL
uGXU7KDqzYGsLooMJ7gagIjy+RaoSQ34G6WI9CTu5MaAQzEkWknyTv6sa7l/ARhdMQrSZIxblamh
SF/DqEF0tlte80uclR4PMJB9EhRd+YtpMIZ8Hpu5XkOWOXCeu9f60ubvlOFdzoXkb+lfYgqHTcWO
v0BXICqXit1wCy9CMUVZJUk6nc+IZRLkbkDkBssodKwso7i3o2RDrkZLKiKBtQjubXvxOOjVD0vf
qql1Mj9+hXd3A7tAPouBqSC/4HUOVHgCKhpMH0IzXkfJSLWbpGsKjG6MGc72cZeZPfd+VmljooXT
lVVzL70PFnzyr1B1I0q6K6kMcU+TwBiei1Z+/sZzgcwC2bi6dvxpltigL75/tnEZAq9d4ENO5sPO
OtvB5bqQ9Iqf751BK0jz8xd9g1hw6De1mo8ubLgiMWIIQ64lM/6Gro4ETN/1tu/N8EWXNuPCYIxC
/Ad+4NcTOlLxVESgrV4YBcg0+3lJA5YG47ihqQd5jWcNsffJIs+a6hgmgT3lIQ/WTSvb5dhxC89w
QMj34T2qrr4pBoCe9vz4lbYNJmjmKfMEVEhWszGl+mMsIS5tc1uuchFuzeo2ZHp6FeaAoUIl1OIQ
/0zqBKLYkJnowOkQ8gMiBMJTTmyLlQrk9YVSXn/cWis+WJ2D09mjEIG33uEP/XuZjsIbK42bDWlS
d/XQM/B2v2XsU+bWDKrT5f9ZTfai4pe29d7ABTtpWZ/Hv6JYs4hOOa4Lkl2p9maNCf8POmPE426y
mTLOOeTR48FC5kpBMxVhi4nTRD16HlxfN6ipN1A5ZgFLOsTT/MUXiVc0b56534YlfD8ilJjLr9ey
EpUX3y/Juvuye6XB6ZqzPnonfHL/wNhzPLxVOha3mAwC7PGtQ55yaswLw+0JbuBbP/KYh0xZ8Wca
w+ZFAM2pgVeM2LH+N0isrusDCBGPyR/3HYfAkJb3DRui1b9PCevsPOAl9Kw+KUfDD9sERDNy/DvP
CliYt5A0Qxwtq5sItCthjslmg9RSUKewz9tJWifERmTq8P+9yn89Y0hymidVa1EOAUAg1oUWl6Kf
2FhJ6Leq1R8CkxBLFfCHAWLR/QecEkiemHAsErP2DvC8KTHqEv2IOMkdKlSocM/BUnCfredDD3nW
Qfpgflh8jn6QmjYED2uGI7lOIlsC4IZ+zlASbzrX8viUXKasIkXt9eMcT6sy27LSrtgIPRa2lIry
s+ezAVT2cnt0FpRs9R5q57DrLzNF5FtgzxTvAUrXfPf4SOOFXTr0CPBNX4nNzWMKTJCgKtcKtzje
ehZPMCv5JaUNQqGeSY+EDzIo9fpAjP68M+Z75xBImkkA8kI0CydfWm28hprX0TEZYfMuJHcMwc6K
eA5ea/UQ3J38VMMeC2Ee9Rt17loURQyGm6NvxTjQw71N9m+M9Yebe6ZFcqaHCFdgViVd7HrbI0kp
/RKe9OSvMgfAKrzWwIMggMy1gZDNdG8CGV7jZ5sWaIuPv/Hpy3yNV0Zz/iuB7ni2QNmD0nV7A9EB
GngtqJvJsvkF9xgBQHfQ5p+Sa5ZrOrNrvPf83HXLOKHhIwuVrVQf2rcsBT+bYbe5UotmycEn9uEy
p+qsNhEwRi45ewxo28b/0zl2kxyciyjSWFi74n/GLe4Dsdlt5KLco4qFSokO9gvtJVHHhgDUy81V
m+LGImKcndN81PMR7p3geflT9XVCr6hcdZmjArXqSibtOL2cC92QKiuwsv1WhJk+75iYoV00Ljbw
wPjxSRKAHhLyebEjo/Mbohpt/0lbce7dNoPrhEgv7yPQ7Yo+KgSr6AgUw1W693prkLtetO2lVfpn
Y/WRPGJozS/FX5ha0BqpIK1x+FkG6hKPuoU7UHJ+WDccivtjAi7PbZBPvY5XS+6pl0+zYfh64U35
dQfAFIFwv2B9LPH967PfzF5IXtdNMKyHspl8KSgz8M51xAO/74iuTNVT1ijt+JYUjMEraThcnzPP
Bfn5DrMDq2IghNJtzAlr8CphCN6bPaQ3TvoI+j89lSKfjeCLcNCRiA68sSkQXuVdg/vNd+Iz3vHe
Golwl2zOxOe/sDWbNxf9tHNzMBSrM3iXUgaS8H4qQO42RXytOx9ChKkh8gwBHKb9fR8KMxgctHPo
ZZ3uhpQ22A3vI7kGuS+LmRJ3V+uTzxlVFuGJ/ws78WOSQZVD3xNoWK9U6IkIn13waMLJqep0v1xA
N8Wi5Dbu3s1XHWofJ/FKHl9XYO/VNXNZpVG8SrIZuRFaAA3IhluzJxg313Xm++lOtMLqq8UdwLDs
1lm8tfs7pAnx/FpFc7P+sjtiAdNv0g8/oMIM30Jj+M75bdoNSjcZYZU07XkQ5DMN4ZZKfpb97QA/
Yg5hqfXGBM+sxNOPAnnrG5RdmBqyKBQKgImpUFxrOZyvbMlbWTGlRlX023Ofze0K8GjxI68y/E78
2e3Iu5iCHhoyv4iOLk4OuUBr5G7FuO4VZZf/WwbVs43GDUYDtjyjSn46xFO3VPqu1TQeNIV88uSE
wXK6LgemE62vp63Jjppkgwjj9i2luzInLKxC+QEnnEULgdbXG4KFQFvVzT+CRJ/Ohq9NxEt7CXGi
/Bb7zlbIumskF/2ktxPCOx2EO+dkxKUTi18n/AIz8qnCFjlQRA15+nHBdibEzaCmXx8epzAYq0F3
2Z2qHa8ez2EqC4CI5dwgGRyyUl54cKrA4u6oRm1jLhE5Fpf9bBCMV9DoMQRpZPBEv7A/2fX9pT4m
K4+r9Mu8jsftdyV1PwX0vZiJDopmEDvzFZQ8ewivo7Mlk7pmUndbV/pFkUhLPQqt5xQb/Imawz3D
ZmVx90NqMO3c+3LIODTKl38nb/cuzJdpEAYWiS4yUWAPJ75wnFiFGsgoz4yldwpMQH3CyAHzXjXW
aS+zkMgEdNgYYM12QWxWXLvpBkqSYD7YKPCHlVovou4Cll1fIhXQ26wcwCOMaws5M7XkZjaZcS/+
r71H5A0DAg528/Gec6RGqx+ax7y4V+ZzyOw5pbibvbQcLCc9U15cpdx81fSOub4yxeYRA7XvHvdg
VXcDHIHw/DgjVlquSmkTnhABBuTGnwsWoq4LbMQ7UWdgMpqk33l+vpEAMlj3otvQmTlzHDzaWNe6
O0fFXOjE8HcyGyUr3f5Ho2TMEWIuKofFSmAn1QbO+SCChwop23qWtiSFSznymedJBFIZ3GmYI4SN
YShPG2afZgzNtW8py5BIzG7tNbTE2HKmIVOxoAnAnL4yTppZ4zPQaows1t5xisoPQKYJyeUIE1Ki
8coQTGa8L3gxmhQiGPcrHKFvTdiVpqHtPY5b1N9sRb+tY3ue4J9OMJHqINIlkc+9wCoseYTg8dJF
jmNWEt/N5p480KhFEl+WeD2dajJ47p0NLJPvpMr1x1GHUcv++2lsBI6EcHfeE84IuGRMvXVnXy16
qpBskcl0L/Pi4FccBD7H1eVpDRyvR6b9e9CH7Oojldj2O3qr0Cw9IfJb7V3htgGk1Uk34Jj5v4nq
ZcihRKMo/80qSnnGbpiqrOpd5pRbxeynKYQGpA5hZvm6IPYGoVaLlkLPvWE8NeJZKpq3uZ+ZJR5P
CmFylh2IVYftKUFEXYHCI+eCZ9bVPZUUkCu41QzgTS5lIu8L7CRlEvNjVzEP+jFB+0B/0N+mNCmq
JnNxa0LVQX3Cwei5ozU0nhweUrHyU50wmdEdOrV6wDMZ6O207niOeqW0QoKIi6/iMt5MKhaNuHw7
cyOFcT/fiB+n09iTyILVjuB6iEHmnq92YL74h9eW1PhFosTT1DJt+MMIx7JMI4LcMqAGha9bBUs6
EyLTwKJ33AfqsHjk+Re21kxDRBMFHmmoLOCar5UKE2W4oZfeKfUNkfIVGXhF/IkdUR9Vwvirq7DM
c/1jACOwsOwO7hdI9uGJT42Mbj+OxMsCdtVlgvxvRyX1PtFcZjf/kFqJrUvtftXG731WXgTlgZi8
VITQK5TToByy7THaPRMoGGzMulxzDqPhRqCbaGAGBxyMD2qQirL/I4Iz2y5ygF+I2wCo3hIopFGB
bcLP72SVaIs3AnC8g6ciNVnM71kT8mRNm5lewMNa1C4U+IqoH+H+DbkHX8KgSxS3MEZZgI/a0E8Y
ZCWccIMLbJNpvodcrIqt1O8TR6Y55gHVzcjjWsn57F2/+aFdMY/hwdYRMdEyil7XXX4o9YrRYS/u
WErCS4V56uOdi9TkIcdBlnIegndAaviFQlGiPHv5FZzr7BYIleSuygZSAgg9lJvCy8TCfRgxAkF4
6lZE56Fdaoc+Lsnb4tKmfEtuEUv1bbAigMdpKvwNP4veDHtUmyZHm1ZvaeVlnaEw3Z8WcLb3yMhk
eGCMJkDl8x+8rvalwVaEGdtQ0cdQGrc8ecPWnMFKaQNYm+8jwwF4rAJ6lgZrZ319VSydqT9RqgOm
Ucq//+73nAZXItL6N7gS55VidC3TtQxEsxoXW2OmV9Y32/wZPOzrQXcPVN6N2IGFSvWNC3Btk/r5
AYxUGwG3fV6N7xUzd6hI3evrzIdz3uCUHJ+mRa4Q24/dfwzTw0a+vYEV7NenBiVKFo1NeKeU07Wn
fzkJMbja+crVrrFJ0O0NwJ7mEJHCKWqSNSMN+TJV06p3eCKXq3x2CmTIzXglg+7q6EAJdo31AAQj
8NEjZIDCq2Ajj+Md4yKKvSn9a6zMYV3eE/Bo39GJZ6OQESq+vxQWB7xh+uEuFCDefh1ic0L39etp
M4kZuT7jkW4qEV8GQ6jWQLLx19LoFim1cJjVbMVHepSfyBO8v0TMmSVWA7aftdYT3tmrdIOU/zQW
rgmzAfmDyW/05wVOHoz9rYcR1qBc3Lb81r9O7y1EghYu42lBQBFUGN8QnmVQ88FQ/mei+OueHjyD
q4r/x26VcfWmJc/pKCZqFE6pen98b6TH0mD5CJ+Tz0+KNDLyU4AftParVBZnWopsOD7xU+KRFNf4
Lxm6T4h34K7XMJsDZiXyjj2JQleHqTHK26gLHMimEYgbyHxJ5YbkRs+aTtG5MQ0rjwztdg4JQtE2
tNibgWbN4dI91GbHJ2LnVgjH36SDMeyJOonX054HUmttEDNNEO2SF79TPNKloLtfovaQeNx/U4bR
O6oycYUEbR1y2q3bMePTbSfmqXsNA1tmFZX90Rjuw8t6QGOVjprANSRjdF6UghXs71GPUrMfclZx
7N+0p/owU7sBaxdONhUGjapM0CWHDBjgTwspyjPp8aGZvmwaME6IfDVtS8m1wxtBN/fEcX4m+Xfw
IPFRe9zhRtvM6Ddk7hYc+lc/9rHP245amIVe5JpqXtJzYwOZXW1xE47gC2wZi1gLGm/1dSbzd0JC
rdCyT+lx5Q4/dQcQEfJMwwAkCoX47pyv5U8Y259TuF5RyXW8RNZW860CdOjF8EN7AcTBsAGZrxs2
7XXgKVfgsesNJtNKHnmZbdQ9ER6ZSyYOeQl46YFWaZF9sfF8hFQfCkIL1o8qKNwTHwZbjBatQzfb
WMiRqgKqkfqdg1vxcdkrKl7z/ZdaiuEQKHlWnDddfPvVfnQs4N+jMVUaqUBIsuCwWBi4AXvXirzv
Ox6Bt77TPjWqHWqk4WkY3v0skratoqUg4BkGQo5yOoc+/W43HjeMWv3DIgvkv83KSqGCfQhAfCZj
iPCNB9CQznQG7KgO6yv86DG5lvIRVKfJoUaxQ7qgzI39khQEDFtopoPED9MIUzydzNgCN0l/QiGG
wRAsB1QPGgTEra9wH9FX9SenEPNNmaw5VWG0m4NCNiglULF1/46frRIMMttth84Q/LlRFEYA65RK
PKHEaCMk3B5PCwRn+IO9reDMt/ZnWREC5fRRb6toB57OQCf5QX3igu3VjdkyWzHmjiMjfLFt5XHj
8eiDtffWt3kl9Uftu1AoYtodBBWSlW6caphG+wSlRKiT6E9WGhVn57+UCEeNbwTYTqwQcEgyRliS
vdX3nzhl4zeQt8/Ptm2MWOj40hWEYqaDCzErCA3GlTLu1vkTwN2zmCGyH579INjaGtxJN5Wcl5N5
YYysakeRE7wmUI5KcY2xLUkPXhhp2gre4l8hOGpBupFKd7/259ljN7qY5Wed6Z59/q1d9J/sAIvP
FbnatGr7+q79heryfUdT2GFzoAtA44Kyb6WDAjAIF5ONI1AkI7Dy9hwcCBDYN2l7pfOJwIkYgfwj
Cy1ungDlJIonPfsIAhHevR4OEftrFeqQQaZvJfoZVW7eNctqpiExPOehA+sWyrYEnoHp7u1wqNRN
2swHgQXcAPrBWXK+0ZOjUNreylZRQlkhecKrZNSV0G0tiotvZeiSrP57bTT0xSMu1B82VxIum+Fe
YDlh1JqRb2NS3xu4xRzROKOtMAWZv4TK+zvcQdXiJGk4MG0xFz2nH3d4FM9IX9qSFMx6fRrIMqDw
YL7BthmM9YG+Db5WZeKKhq6XnqAKu8qVS4N+css5b1sIGDJFO0j9PuTh2k8bv+XsdpW7ggapwDPl
v1XEdVLTcw5FmeU44POuOglM8VAZivz8SBW8ZmSX6114DFg9+MkfcMgTwQYvT/R6PXoX+9zlpFpx
m5j3mMuduff/3VTElY0KZbDozwICL9UhXcKRUeBuFxBTakJ4tvZmwNii/SYFkTNYJc+1ukL4fKh0
pLrTfm1rGK4b0MHrRDNe07EnbjT7FNdw8Ix7LjjKFoOGY0sPRJTSEmaOva8Qc6tQfUZ83MNaZ+rC
mNzCb/Pg6N3mH5s2lW/Ka3mnsHiO8ALFVtmO+61w7fkW87rajs919WLZoMW+XGO6YzTUoPnvltZk
SRL/zLKZe4VV/TC2zzZKqSUaqUJihHDzjCLhMSB2qIusRiaxu5ZCyXAtELzK3i6YwrfL1hgWW4XF
wvSM1Rst7ANej95CXpyGPkOcdscGfUU6IwfbfRTQh7nR+GMORCG9qLIImJo5oemuaNtaQQj6Le5F
04q80jQvJjPsNIHGO6QFZNeyfzZ4NBBlF6syU/zkmeyYBChJIce9VwJWagacKQUGwc1xCcGCmxWx
iJ697SZ0Bs7RpFQsI6i2MHtr2mtvPVgfCvRGgWOv2jKiKuOyQvmR4a3oa9J4B+rRMlUZwY6XxMLg
kBH9cYhp+H8Ju3FQsQ9vO4ItKPwzClJ7qVcNJ0xYQwCkmGpVXxzm6ILI5yB7oLmhKaWLqMbHBbGs
tipYNN3KYpyDbx5hYTlxv96QBYX+0ZPcj+kFHnbvEyDgb4QcNwdwWWd6VAtDwWN8PyWOkc9xga0v
iIcoUxkV5JYE5VBZKo2FgRHMi5uyERjgUYSf9yGImcp3xsFlPJs8l6ddoNtvqPcUVzew/jZCLTcl
b6ry2IcouwfpgBkpAQRhe9aDxKjF2Ad8TE65xHtiBi2xS+YhLR8MsnzGaiuCtjCOsa+4iqJJCAlM
zGxsfNn6zhGIqONLSXLlMS43ZQx8T4ChmwdgO/7xPKTEVQbMTbaUPOUXWumnxDrJTbbi5kUOM051
qhh/ebzd6P5Yr2PyWQAn+hlb4rwIgwVBMkbNAAlrGyQQUKlDpMbSJAZTudKth/UK7Afl24eflfVG
Psm7lrbNhqELsGRoJoJI0q95ffZ1atD32xmxJNbRubj4JDsv8J/8xaSxlg+Iic3wVEMUKmKAc9rG
ORLePiTQejCltoklCzmW+7NajlUOtJSHgBdEWqEuhP3FRyBo8wIFKiapDcgholdfmtBOyXQR2OKx
KNX2BFY4GA0ypiW93paPzMHeXiuKFBdVU59zSZ2Z9PRS24qvOeNCfQmiuAfny2uSJY8R6mF74Im3
It51vLwRkYNHfTQj4aLg1kf9viTtOL21HXovcsW1siDaVqq9HoBrjJcJWC1otjZNACqEth/W3Ydh
bgSHauszPWq+dGbiwMZ93vcKhX7akJmZ+TH7sVKt25HkvbURTIB/P+mWqdqgMn35Uug4uXTTMxva
agmcZjUYr0Te0tyParkO8vJnaEg+uUWBt0TLm6Jh08seaQ4RYk1Wu5IphfroWqjSS9+nbMOFzYEE
dZt/ujhVk2abK6vrP0ft1nDCAw7zE5DOPB1VNA8lIEEGNbQdlO8B7MlevdwUtrjP8wCqXQWn/B8G
XMxOtQGcnrBZ0WPbhqfQZwQKdLWLsZeNxPrUKq+jWzyRPV8XUMt9liIcmDHHa35DXvf7cMgZo/ej
X4Cy8EgSGS9ole5qxd2WSQFOSKbS3LwqmX8dUr8jfPiq8V0OHQQsPHCfpx02JmEUaLktztI7Eq+x
S1r2Q7d8yc6ueOa8O+i/Zx0RzDt2LafF2qMKfnluXglddbvshr2rXyKd1Mxpjpfdy8QvpnE+w4BS
b/VnKA8ZhRwpHedRX4H7xMNfOuc6f6a4EmVOD9fy/GVRPCFzmu3WYciz83Ba3MNjfwhV9nztHDxe
RH3pvb7WpaUB+fyQfykodbpMN8qhnvbSvPlLeDF/TBDsGsJA4JvIgSn3WGKXI+AmZNurL8Ct0yui
W91tGRm4wwCfqsEaZDEK+46ZPsKqrtJGbXPAdXWMmrKw8yJkiFB0xS773IV95glvsi4SF21fa/dg
XA6U+2KI4iHKrIpntiX8f0YBtOFh6OiSadILovEPOaKFlgSrbREqXXuQBXpzgP7Mz8LOG/QcwhjP
FXBU+/bPuV3HSvptB9uyKObkIxNGe5Wb7ITKBN5TgPE6Q61Co5RVP8hbK1Lxf6Q8J4tL+gcZ0ChQ
OHpjeHyGT775GVUdFScpswD9AqTyLj4JnirFwBLtlL+lvBTwNy5l9JqdRzAgJj0xMsHeWehJn2n4
97+7PsNFKLgitnxK80lrgLFWoXaVTNpSj5Z14sCkgHuUJyIeYDYEzEdSlE8mrsn+Gq24mQLqTLWO
IsTzWu7LU8CBdZKRf36qpmpSTrNBvxJQxbb3Vp0ZtS6J/yZwIwhexe/rd0v8Bwn9r/sElwJcqNDp
WPdsQmiFU+9ncBPPHW8UMpzE3+Yp+ZH+MbsrsNvf3/9YOVRoyR0U9KQpWz4f4ZH6OYndjy1tMsZ9
oSmu7i9Vg4CvtbDzJHRzJPD2ZtmZ9+i37Eiu67EuGFT3BwAHKuXJmwPCJ/cm/jJDeOIYjxq+HbIs
9xv4fgs7+ehIS5h/phPpAW98EmPZKE+pmSMDhlrrDpJ1iLcttj/3iMy2TtwZMb7dOJDpdxBqVHf0
eOK6dRcK8bwE/93KVlHytg8DOJL+DwAeseCf22K4/+QOb0c3975ZlbHZaqX9SmuzzmTnMkUpkuno
54RTwT+xDr2MdcjcSBEMyf9Afc9CfVrAik+m77dzqqoGfSq4+UhVoWko4tDBmPsUxen6a3t4fbY+
5Xoltcwys8gwaU5Uv3R3RCG6RM8J66jgRDEmOfWX2rdEr0SExPBnqdqFb4zBjDsXtb39V01HQJj2
nkCBmCij2CBcNuUXBh8JcjCZejMbORbEANlOmZtD3a/nKgFnpYqLBd5A6ZMeaUamYU1zxrciK6Ht
ETQnbQirahfCU4CsrBw+uyW7H7FxgiF4hBwzKlhbAytLmLYGXQScDJQiHhcqpgcMFmhMi8K1ieUQ
kVwvq8RxD30TVEmJE1i1gLt8z5MapK/sRrt6AvsWgzfi27W/5wCxabYXjsMg4hf8UPINvpaCHmm9
oz0uHbiAvRO2ZWb/9tyfYscmfVXMAPKqRLZPSkMxedrF1L4sru/is+X5Mr/c4IFGkbnyJ9/Q5fm7
41lbeFMrWResmkBnMMqUu563Laik2NUp7BcKPskNxfdBP3RoA/isNBnYTRfDtJ5NNGgYjOOt9YVs
8o56QRhKIMzFMIVGGGfQZI+QN1rBh87OtTOBrNH42T76sBhhqcATNpZucnfsvwHbLRyTfUorwvya
fzJFUljHLFvQwNidWySBZPKMj76xi6vrWG/2qlr3Jk59cI5F5tPVFXeou5sZhcJlW6OJaP8R/cj4
iW6QS12XU6zNVidCI5bavez3MIbdAdp+6KIen0bM36inwITYd6phyqwtdSLtpQQYGDERsHRoDbVL
2MEp+H/6E+zizprtE0I/nWqMl/RYemHkfgAxaoEMduab8fYxPNEaz7M1vF41m6vE/tY8VjZziP4K
H22ALL1qDINXIGSbZdMi3LBScX4yHESush5bPvuY/PWGpo2/Qll3Bd0D3JCq+SYhH0+0FLSFmaAY
t4Rgl3hreeLz7BSty6Cl8HHfl2MI3/U+7rYogbVlCFeDBl3kW1U+4FKvGEkVHBGVThn6IfA5VpVb
c30Qxj2jZyokepp+UXNO5BPL9y3weh5rKnxN8nfetaH3fqNoG6bz9Hp8AiS1YUZjowgHrCNuExvA
WyvPHcQeaTi0/toUH+DOQJVXMLGV2oBYEZ+Xf0xGIY89ZJR4xkyiKB/BsuwIZvFt7O7x8V3/iT6g
ru19RtrCFHvYQJpUwl8k7JwMeVkP2MsQMqA4WEPUKQ1wiA9WKDYOVd/bzqTDPw8rCl+6Yy1DlEf2
NJ4aO3h0TKSQZpC2RB1ydThPEwxBjNktR6bgDr5DiTBNuRmTmTICw+/eMkoXSNTvIYTKIO24UkzZ
w7QnICo2StN8Dgq0HvvMEhPkKfUrFGdV38+//b3PvAoGuMKDDY+JbtOGYrsiOEdxNvSKeGYY6MJc
TvKjO44tUFP9LHpre5UUpvjklRQCoY6LXT3z23JhniLFTZJOtQdtrJQ6yYQQ5bnmfQAMNqpzRF9n
LyoLkTnzloBB91G2ERREP5a/kQkPvUJjLcnHAnnqAgQIQjL8hMq3iHKXL8ItPNKLubkkYHyZ7zk6
YLrwtHgGb8tvI89OFI+2Ki9jFEGHGLEO9KWVC6ZmmiYTnswMH2+MbWn0ZuIoT1dOi9tUE2DloLjX
xLIZLmNSKutrIAi9/IqZxJNQzcep3SyZOZUj6jziDcQl2fTAtTamr7I+IF/Vn17jsuNdekw7S8HI
SYlRCH8toBEl8GSqDj7OqW5/lvxhprGquhjSntwhy/b2L90eH2BmfjwDS1pZ1iGGNAGUt82z95lt
Y9PD0lOJxMMN7n02ASjEeXmNN+u3J+cuLgGfw997O8+M+jEL+AfbJTJ8JShSGfjPpLLyBIkLdhQo
lbjl/a6t9xU9DQpnw2tm2rdYzS+ItsM6IDtVxoqT2d4yHq/xDIsn/zcfZ3dYT0XyI9cxvndQ7H/U
NQi/+Kr44yXxi89dGfZs5SSxJV4rjLKOuGVAC6kvQyj/oN8xXex4d4Ghx1xifOZd9kgAnXBgVxSc
PPO0P+Y/KEpEx4eWizvDILMniCzdctvX5CqTo6s1S0nBeD/OR6hCLgQZo8ntP9d38iNlvJSU3Y+F
2NQ7RYGV4DyVhyjJh1EHANtMyL1idjCsiYbQ/jGx0TqJSu5nrJQIKQ/uE9q8f5iwZnnQ/y2nDhBd
xnNHzaRns/cZHZVOtkj0P3v5JiDHBen3kX/0FlM+5RitBu/e0QG+H14r0gu8Ak+1lqjpj/G9dXcc
oMco8ZHT8UhPW83075tgrN0F+qf04Mzlu6tzF1HtuJPp71LEgXhCx1vBwL8lEIb2nB1NxBpC6xEq
LkWuVMeSrgkf1YIrBLSGuEO8BxcDOQrwPLPR56kn3MqwDtQXGAh9Qo9INZkwjNUVRWK03Ad5nkYE
HMDawaZlB/r4cbbn8FrXeZHSb4AAIoJaL0byAU6bBSfszT00kZeTDqHOoaMw599yRouBe7frN+op
C9YWCFoDMqRGCnZyJOMcSE81mcqMCbxO8YdG/H2NxnyO4ZYonlCpSom12Y+vj/ZcqJSeWgSV9B+3
0LgijIGdhfhVw1N12tBBC7evIuIzV6kK8VF/J8kaUGHqbzZ5SOLoBnFrRlH/0rfqA88+4EVIimXn
yReIueERQtUOYLYMiSp+WJHv2HHHIB3q4qkvhDiFCcoGw8kRfcd35DpZSl5MN5blL/PPJaJUgHIU
eVnYmIZxosdYlawNBoW0jMqVeOk2Evx7DcdpnvDXE69TBRfm1UFzn0zxUHKYgZKT/8rUXIV9eLtV
GDh9ihOs3GjOV2512tM4+3kLJ1/gkAKRwL0Q2N3J3Ny6Z/UUI2QGjA4DWJw8vYF4YrA/YtXSUlcv
vCtWMk9i1K9Y8l9DLYLx0jPff2auamVVqZYqwfLRvA2AJdsvR0evElvZX3UTnzA/618kk444AEOe
IE+ogNQRq0hRrtxpgmnUwg0VWusM4PetIq1nk6r6jrCpBqAui39BkqgbxBUwWCx07BTcCwgPPNlf
Eo6qznP3atDGYxWM6dCbRwz+wJN4r8eufxeA7ZpWeyf5XRKT0ah+8qedQIZ4xa8tl/bBMS/50uXA
vApE5gxUDOHvt+vwVopd8xGYVN+Rd+GaROAtzRzHa9GSgZlKPoduX6XxCprmoZmmE2kVsJ3VvtPo
fWs4kUEyLJ4CuLPuyrhx2AS3b/WbAhGnaEH2KSisacjUyKJ7pUPYawNinx7RykboKxyaz1tjUdbY
p5qm85qL5/3J4Ruw7evrOjdrHY+u7+UPtb/ofB1BTo8paNBnO6OMgvwmp7PSAhd0x9AgLmFtk6MA
out7rrnEmiLMS7M7zxn5iPbt0U872yQxG7egVMSt3STgZKw+CGhE5sfmTiV7wRYpHYqDA3TpYznh
TUXHAZ4fKcW1BqY74ENZErUmfSz/KEGg1V1B0yt0Ah8HbytlONt3nXS2Q/H8pDs1OUIPNffDtFHt
Icyl5X5BWN4HxaQ48tsK3oaMzmI49gHz2YDtoDFluKp/DGtZH0igfuZUbfbyoAGubSczcu/n2WBk
j3kdp5uWUWmELAJHT/5nXxM8Rn99v8miE2KuPgiJri3iIqe72XWqhsa2knTegOt5aQUPTH35vrO4
fP9mGwfhBXNOLK49EqsJmg5V3g5i5mIL8s5eCPO2yDyhJyymclNmFb7Qjhk4U9oYJ38aTtMtiMhY
TqlAE/s0GcVyGnZ51RMm4Fsi0swY1G3F9T1VmuYLvFpW2rW4/w2tLJl/3Qao3RW5Wf7tyHwkmxxi
75muu6XU0Y2d39sAdwqWPk99Cn9eOby+pvmCM6SGO5ti7xlKoydP2uQqgUw7hai4+kMwSDFpoUKf
03T/kCWkp0C3XKEJEmi5Q7z2uUoQD9JXL09FBen7hmWb1jNRxmiXUapG4A6s+qjE4Zy7JaF/u5GC
MFRWZIjwZm/QDHZ98HQWYTYIbrqvdenSmaCSWh2vO8LOTinC2X0ofxy9neeu/073YGeyy5mdbnfq
7smdsy6CLVFQ9K8l5WjrfD+oiisId6yJ9FC2qGYkuhZvjplcRZzi1lbp2xz07vKXu8by49HUMPDL
V0NqYpqq2dNxAw0DIgOcH8nktpFBbyCeikfQ0qZ53dHBUzGYG4bqJXwshvJFVIwvuDhiSCCl+MTo
+Mef/c1lCwnkj+FtZ/oHEw8JSTpP3q0B86cSRB6TQgTjUr68uETo/x0GBpQnnuwgb4qFxFqKlPmF
GlLZTrIFfOXn8Sfjo/NHyUTG0M40qBOW7V65hY2kdVmgbDVXIkqimwQWUyYqdnXd473Sn2Sl3Yhd
NWsdWSIPy805N0xp91vxi8Ky13DARZmc6+RKqxzE5zT3VwzwBGicC3AKU/6MCAWXbmmvbtho+vtN
9eG166ttEBzLqP1Ti/pZ1JGo55fpteFjs8AGYMbyI/fFLJOf+UhuSz22OLlPClTeA9vcHQ0A2avm
FL/ivKAZcMP/4mP5OKSHbTY2ow0QZQde9/OHffU/ZCvpDP9xIqnyfhhq8i3bhX+J6QgKyBFJfznz
JL0xEhaRKWg4nhCwPA/mUPlG+DYyiXAb+ItZYIdx8XYjmk2NoifNGTVOfsvTzvMqPODK8XHygGbF
dqCPXs/hUyhwqdqMklFuEOMZKszRwe0MfBYOWFZBo4tYhg8ILKtpLCPSA9j6fPu9Uy3uy70RFvu8
BAL5tF98EdDxep+m+sncyyLV3SMG+H+CO1WxXdrLAgXuS/9CqPxuiOzCx4/8QwmJaBOqNDJ2zsqp
i1Z4M53BNIDoVhGA+kEZ2vahAmYRN5SBy/iFzg6/c8ODx9x49bxDIvmwLk9qh/6hVw0eT2U754XH
0FZXSf5q5aQMy7APa1mwomuiOYpEvseam8MMsGDx61AC4BfkukGT2LLCv8bvdYKWOQoi//QNA/fM
Wh1oKn2CZnqDnMcd1kTd5NefszG30uawsuTP0h4vTKStOrBoxJDNye/EZ3l287t/5R9AySn2v/7m
5ZNtwHBKUMb8vNXlFV/BrjWoj2q4HwSAUWtUQ7CXQAc4NpK61pWw+syx2rP3uL9hCKbip6+YnEUR
N9Vezu8r6zl3F5k7wutPdjPA6kxZ5gGO9aZIEgoLx99CC112wwJwgoBNdKYTawZIAN3N6g8+gEFY
W2/YfGxnVGJD8dDOt76UTJdNTjNAVmeBshFPg+0/vSWm8cAm5JFZ0309+MtQ17D0PRB9sf0uy2oW
hHoJOBhZIe1txw5DqEmHl393O/JA5jdp4uWE9FoRcgS/YobB7GVHrPQPbXH68k1/yPROT6FxVFXy
YnNr4Wdi/JWUz8/37LV1UfYm9gpUtHsG5lynFpv1yaMXmhuq5Smpd73ZcYtVjzzU49ffQzY1uQVx
KNniZXJZtfmmN297uE6+YGoESUD+fu6E109hlcPJdEMVnB9tqV8TkmpwjzBWkmfLeHbYBpeHRP/r
RcDgZZ0nKAJGUAxdxHbP+IsMRheoekS8Ss4mjuKIcEssWPX0uz6Yi+xR4NhA+OTGmOttX5Oftmea
UQEn6NmR+xFKFEoUVMCAAT/MZYGMSU9pLPP06y5vZodjFme3WX2VD0xekqViH7Z61pkKeByudmTs
d8qhhDI4l+jvecP+nltw8tE2UKSF3a34LhrGagnOLB7wkmG4uFB8eGelIZrlV+BTaDMkQ80E1I4q
cm0NM4UhmxqDAhWrdf7o8x/ndoRwwRVnodnFE7UxcwSfmskidc2d10SyAElrY5bLxNz7iHCaXDAx
/TXBS0kODneAZjNLTXsWQxIIjIGHLDICocdmoTdQy/omWEeh3G2zer54xEjj69MdHHHNSrbAHP2n
GU93fnUtu7uQInLpTlccHdvOXqkrrG5zmggLxPubbvsjvztnq/BmlRU/lB1FX+mVn+clDR6khHVd
5zKbBJxRv+PsXjkV2E64s/1c3lLFiWSS29avUD4new6thExxcoDmKsuCs94Mx+OSexzef01L+aCq
4S54FYkRM40Oe/BdHNl8wtendSjBsLu0vmfQwbBQLeZcTHfgW41akAPD1NHLuKZwfRQ0J1rl7rpc
ZYbBmLdwLpLUr+/lzJ+Wqc0xO/bc6mvEc1CViiIuNeqQMFUVQ70ersVEbHARFj+qsr0VftVw0kJU
8GZfOqaFqyjG8OmWYfMJkzSNwSDLCSPQrFFMhGiqMfyeOzUotq1uCf8dxV/8qQnVsG5UrJLVcd7B
V6WzGeDzdoptiS8UVJ/a0VgcAqPRg6sbrPNU3EqUMGjYOkrYoSuFVaOuhR/9r0vaaRUByhhT3rjm
D+ygeGH8X2KWnReMk9kehJ3D9aPyc9H4E5S6sROq/AIu2KEij7og7HAtHSqvb/N9res1zw3ov6+B
lUgBobl7VX6rlb+EtuoLAQkvgDjRBXYNVV9jp/AYovrslnwGieyExJgr8pxvtb+RnRB6SFssmZ5r
jQqBvJnH/DZjd1d1TwBQCYsENO1AsAnD1iWR2xwue7fVhv+qsoyM8qvxAvQ6CsyIOPES8Ad3oi3I
k8z5laBJICpxxtN6u30YtLkFC7CXz7E16yDptJzOF3qfGYl9E2yGtKa4Oy6FKpgo9Xt4XRAIidg5
vt+LiOkhdGEjiF9XKK/c1XYC+/ueThAdK6whHHaNuLc5aKHlPMJ0t+Dm+YHkiUPOgWyUKg2m3gYh
UwXpg+0VznZG13J1YxxKqZf5KGNXfixwCsNNXen4lROka7EtHABeSBMjJeldphKS47pHxlkukupW
uQtaTtKL8o/rogtedh2JC00uy42e+tzHIhfl7GKwjEJFvcfwWWvNlgmw7lwYa2ooD6XFNHmsXnMt
68G46WYyaTB0vFc5I7hQbutkN5QSYo7CSmcHMNrk+tbmAbIvq0vlmrBIiZGArYXYmJPMcBQk+kRo
jq/7IaPKm7B57pm5lu0JRezUNq9w56EkCaddl7TqmkqVlbrpLltTrZR+IqRqs1dja7Qbz2l91UJS
GdRDj4zacLYXiNUDRWei/EHtNfT1377h1K+FzfiKoYyKAbRR7CZiffRUtPF7ap14bjNRrOVbi/8/
GCYOHtEtXtfgimKNOnXNs+0dL4ccJJOv2UQPhFzkZCPYAJ9f6HgOnl71/Gr1O1JaS4FV4lDxBL4T
KjWr+Jof9fSK3MeT8jYHeghueWdNaEjdseV2lvQoTOkRsta7kAoeyfEijGR1Z+YsK6bQ97s+hmFr
boBmU98IReO9il3YnHqarVB44HB8WVYfhqvHwkNeBPX5wZDhsg82ZXugIasa5x6nQ7CV7WWcTQDX
QyUxSE7eOfiEx3ZcE7fwoYWBWys142DnJgCa3yGA0CigV3Vn7udsTQBPAueM15KMaYwUtu3Rfe5L
bL8cwAxzhVdeavtVOl/6gOlSGAmCgxiYHrdzm3xSYI3qv2/3Tci3th1xJ6/XYdEGSu8IzfatPtWj
1lyx+5uDf6Cf7jutoPvfM9GOR/Fi6eA8LrXxHxf29Ge/qYPqS8NdpkYu0abSc081wR7J1IQjnkkz
qSoO2RXUkghgt4A1YjCcDW9Em/5IsaglgIUqAqVlXIS+j8EUVJlzZXnlVbzmQ+0NLT9RkJpPgyDa
idRMgcBT0xr/IujbTDllncWuuezxUpjihJF0dmJ8lhSJqLZpjGZtR4toJoAAAs3LJ4tDxw62WobA
qiK4O1T2WUY7W/GIE8ykgrtCbsT3tSzkfAt23b0QICtav1YGVdkqXDA5i3laCUUj8glQvowF5fET
bQO0ACQQKCSduw9KqKnvDOKbJWsPyfSCVEv8EVtELk0T0lh1mxJpS1UGX29L/GJl3KsswsIlQ/2O
E3hWc9lFFdDq334gn0QZZsmkHcAn1o5agUDrInQPyzacLNCrxOEzAszCDFLYhDOljrKHgjRqB5VJ
Abjbni23PT25e6HgaHhjxxzdk6RkFVVGYFLnemWfqpH8hXxwcmBwQlAsYU6sCAy8ua3TBf6SCcyQ
fVziNuJbj7Q7LvQv9FQarozEJc39pfWKqk6FkKSPvyw0eXP1uqtjvBii4cDvkzyJVfVbnDHaipf+
9Eodpf4/SN4cLGOqkKWyoHu0R7EixgQRGc+aaDI0gMLGwy0rdOV+A3ZUppoMsbZiRlwNjdzs9Jfd
8SiWRgt+xNo9yl3J1XBy7Xx020Q12LaP5N/VBUOk637OA99FPteSsFQ6NTmNNmL4IgWLm+x379AO
uFwKYfeJlbknIymbJNOF8GUiZZs+esQwYPiL3qcXHMzwTwa3w0qSuBOT742o1I6wSb0u2+eO2/b7
RsV/isdfqK8+9gcIeiMNDFm22Sex7dNJSgNUwLQearstG/K/XyRycgxgAjboXuzQoFdudxSByukf
2xqMAi+DcIpUknn9RtE0yaL94+JQjsDPrO9R7xCvAsRLyYAaUpz2Vf0uQiRENThrBOACC+nMbsb2
ff+HR5Iu2dmRaXmjGzqte8UsDvQ3n1DMT17sLPpmjQBtnzMhtkSJyTh9UDQuRH5gJqjWJfcMS589
gcpsnE+fUaKNRppMST6UD+svt9XSOrnyIaleovOSRueotHmK2ngLnTt5oATZ3HK2Kf341WAXbxG5
HJle6WDpu7P5gRSuAvtcCmsVguuNvaIpGvsjQLf+X27dqpK4LGfD1jDTs2KWmEbyV662h4FS9/gJ
tsYyS4QXVo/o5CzckQfTqsdJQppHHIOoz0795bpBLYKBwBVZv09rpI4KAVuYUGHEC4aXDAR1Iwtp
o3dJDVOpE2JKKxICDF4Z7jsjIPwZm8dBjSV05DUmJ6IKG+o1HHKTvwyd7itDI4D4ni1u4lR+lVdA
TLc91W41SMOgRhvQBB+pqlG0T1JeolAMof3JItabI7PJegpc7vwdtBWamHj4lOub2hzMn/0D3qha
/XjFHAOQ2f0onyXpkejUzmF5cMiIZtr65OLMPeubQJLrSrz3Bzozo/nC6Pso13+TeNjVzXHx4VmG
mjRWhA52Enl6psgSc+T//oxH8QDNlqsm2G7md1Pa2wcRA2pkx1NRsdld3H/AsDXffNtcmvqMp7Hq
og4mC6QJVWdtfKHe5UtbgHM3kkweErZGPjZ5Y5t96iHc70C61JNUl+Jsyt+Ts8JH5hHwLG64TDWu
f9kds+bBNSrKs+OXFrNaGjZbbMkcn+qvrRPQRTWfSYnocXHGY2jCmzy4CDOpxQLSj36uz/GxGBN4
ZHbOyUgBJ9jyAGZacZACAT+SC4rsDor1AjZvhLD9MgTMyjpWVehUKrRYt1S3VexgdA0hzgZcPMFV
4ArsTdEaS6DIvjnDO3Msnuf4DeAVEBEWEzUjCNwicW+eWhNYtVcFRI1Pj3WpPpuvBbA35p7l+Pxh
we1pC0dQpW2MxGABSKAS8z79naB3RRpv7cKU6FEbAAMOZn/T26eT0sxy1A6VX5xGXsizC78pYAVf
XhFBs5XgsWLw8R/r9Mb+z4ux3XjilPpJLKF97L70PDX0z8x3Otbqjqv4tAM1ogdgTJI0mqdoU4Z9
9DjbkOItUBnwlBZmb3KJvJpVeze/UY+xMzAs1MxHMoaZWGtV3Cb9HhPhET32i/YdsPLd3qxYSyXv
m+Sns55CZ3u1v+F4A2EWJjID7fQSLUMbgxXaCZz/96ar6yn8jDhFCjquGHjQI3hNsOPylcU/rnSn
wdze9DgweoKJKlSD9v2DgG8FbFAbw8u0njDHfYg493n9Ii+Yg35YO/Mk5sBf+qdDvEPXb7yGSXAC
c0DYm3DGRHaq8mo0p+Ce7P5D/DAbJjr/8ADgyrrG0+I4F9E20H+aRtjYO3swDWKlril1FmV48t1t
1CtftpCCWae4hYxguAF+/p3yldpXh18apLXnqEghsGcsGnZsDmod6GVPJywqylYeCUoQTG/wC0ne
SP7TnwLcwbhpYC5+TuuibPIiBpnr1oR686D7LDWMZRjDIddMCAOYa+akTgfQXMonlby8720DD9G9
r8jpRTMaYtKy4mBWIZJOAZzI9kVKntpK/KOnmD5FfPxk5Wc0Y/i7AW+VFSdPgUgcv5Q2x5BiK30u
lh+d7thYfi7lbfbWZsrFkLohzFFFnNiixKgBGlQP3Zohz+opVLmH+TY7m4voeNj1/6FFhuNmGzxf
sQVQHdRcRCBv4PuYolDj32ZsXhhH0AWsdmw8OkhbGsHsekNjrm/h3EXkcEAl+HNz7K1/pTIWvofc
LdjMHrGXen1EzgVOBGvzhTw9lS/SghqhJ7TdQKrEg401l8HGUZHZ7DGQ0OVGwoesrMYeoZ3eqfWR
jhgwD6XLhjjxZTx/o/ZqiXsJv/9F0dgU64+LbzMakGK8eXn4tljZnhSjED31+BoBO33kpW8BU8vJ
Z4zysvoEHrpVnSWXT8Gv2yBmTTZkVLtyWhqjvTAYUfQ8hP/V2ZX6G+ecl7FW7udwALIYEsaPCgk2
b3fyYmw6asPYdcTKIxkZ/eVI4KEq4CrGVFQtmv0kQ2c38plWvrjFAiL6b6eAkLkJ3CwjK2UplVAy
RsGUYe42bJkRHQdswygqv1mf1tUXBqdNGCotwdO0htjMzG81QNtSWUypGMXagwmc7uhNo+QBKrLI
WYoHH7v+CQqOH9zwLcMrpVbFJJk220SK4eMMAir5ATU8p6q4Kv+skeHfhSFthUb6mTIqzHgseDzF
c+bMwOSjrkVu8BwgYSwaP+LxV4JZxPLcEB1xck+DnIBEPU6S6+8ByU8hwNl4kKVziZn5rxEPz9xb
kGwuOdNfvFkn6UlEIM5w7NuAsPF2fyyqMzQZBKTojNCiH3RbrORdodCFbBYGXfGsaPb96GXdmvzq
dh42PczcnGtbn8LkkB+fuaLS3+tsw4ZBKnTCayOLqacpxLYjJVFvhfIv5LPaFHyDk671LPQe5rlt
V8wTQccZgOAl3P3iLyqWxrRS09x1CRBCqrrGa7Z+7cAm5WU3At/FpaFt3htw/2xx6drYAa8sky2X
qkA9q3BouROhbN9JXaiAIIZaW6UsRfRXj4O9OQkQMGEGHx95q5XPktrvQnTs65BPTnMMDG/Rw438
fe7G71kFJkMTsBrs23KBByLlxKQUmL/+G48q9Qbkm5tEY2Y22pJAvLYl/vBCe0K3Z/cJNMtYQQtb
01ay0toFdn9kdHATu9onTzazBlIZvOj6q5JgXg0db9KU6QL32+6hVJmQIcoeJIeYB33JRdixiNcC
s1pTpVRe4vbyeNIp8DrZQVltdiWfBMc/iS8yMDWX1S7i2sNAdQVF2LXc1i+kwSlJmHQRZJ/0Ytdz
t4Nma/1qKd9hWH0u6E5rswLut5LRQUJzRTwM4yU4nSHKYXFMCpo627NIPSj1SuAbnLgERgjNSN8J
ly0Fc41U+2ckjK6QD3TSDfxJ1M6BKwxw3Ff5hIlOwEklY3xCqx6ZGA5l+RKWOc3BBr8H2yuv3D6N
Kn5iYfja4gixYW50FkB1jKjLd34lrVBg0sQMshyaZ6nCKFe79W2fvS4hUQVXmLD6/lvAEhSdi5GQ
HqQMowNA65XXOf6HoEQUwsVRM+GWMuHzQGaLzXwVXiLKfX8mrWzRaMkZhw+6jFAaDAd98wuPtOFv
MK+KSHmVZuTZ8B4q77RCZjKiPxksA2a9B/psG5nOo3MwGfx3gCC9v386+XysZ7skWNy/tVzWNuWL
kD4UvCc0FPheUz8iV4Gi4urGCce9y7G84k++wRpZAj3hU0zS3UDWpjnjVV6aleeIVKpEZAgvCv6x
RXL1sTJ4DL9tkOHYWDvOgKDy/op16eUiJglkIb2P6z1tXFII9ktSnl65dH4Kae5LEA+wcfp2fflj
dO/lhucAjsnt3ympEEwcTgII9sj8C6kDfOTjzTtyikhue2nOLzfkYC4ZgHUf45ru7OvxgJAouNO/
jZZfmjIc877XQMMnKSNZSZzFrJwM7yI6RSvjorvRhvjKI+6Ct4RHkgiB2vwh+YN8LZI+MfWOggNd
ba48+qMCOn/qh2WuF7JrUP2Kl1ZKeSheaQeFVvaK4YJIf7RnL118WyImbM9QXExd3dpe7hKNbWpW
FseUbUcailZKhqWBU1qZVeaXj8jNXHKLiSw8wjkyOLmvWMSxaS3YREKFwf1T6Xr598aJdwoZlOHO
MlXyTqSk5dgTiTASfh9Iuc9HQ0rWF4TH29WZOVZr7BB3/9iqbAR1B0wqoU1XHHQU7oTWTS1tWdtg
ouGhabm07swqHTy1HTo/gp0wfeZajX6i5CcBdIHxFIAdfkRIk3Pv7qAaKLqOHkRSmDNk4D5ctCHB
bGi0so3F6phbfeR5ehLSGQ3ZIehzDzgy9NLKcKrBZiFeSoof6w4tSKtRteBSHEcqlyxU43TDkmgr
x7jmhMiAWOOqOgREFg4liUZ4XOKiiDyHhmlGxLgkFIi5vwipWTHIC90Fr4BvlFmzUX6nRasmgegU
4aBGTwmappTGzQAcihYm84SZceYEhkwH0KK4p3/0CXJ3dg+w1bqQ3xLTlAQnhfppKHUgOcqSnHqA
/yrF8yxT7xrvro0Hovv6xGf8wV9KllC3vVMEP36oy90C3Pc4BDzfgCZ9sRYEZ3DXuapXdELM0Y/P
mvgrF2WBuhSx+B1MHy9FQzwwPZ/1I17GJf0kcP3CaiY6ViusW4PH/YJXNnrzKmwfyL6BKSh4u9Xd
RHY0bWz5V2vuUj2mt0CkD9XQUXrwXXTZe25gZ3voXrEOVRj++AMUKz89S5BMEc239H9c5nrCrN6t
G8emJgiRxYSnemiSH7bbA/u5+axDw/6DUkVIHAWVFUNwbc7JiiWKdtEdponLOon3Ob7spCDRAjk0
7VtreI7bVyBHNuYeZRuZdiojDHdSnkNxJZRQ8TQCQRZD7Ah7xEJu0Vvr24o/Js885gnT+WuM15Lv
M9rj8onpSXDWy74X6OuxFQ9lgjv6Pg3F+/o5xIQJZEgODhpaD8XtDCQ85CDQzgWui1EQf/7sn4S1
cDPfvRbOwZErDPkUzS4jMg3JGos0YP/qCtA0YqLheQ/qV2umrcsfY9jjHgElcCkafBdSkm/WErN6
mlAGktjH68nBzg0f8sJOJtjHIaylqFOz7LYuyvSa8fLexKzprVf8vZcdyjmdNyWDvGEhgzqezUGS
JZ54uZZmlzsHOQRSlWsdugEMJIBAfbMvECD1HYcJDF0zqr0i9qjY+DRbQG1eXM3tt6Qznz6tY9xN
b6mF63Icla0YXJa96xiE+Q7ubEw9kcpYXb341B/2cU9X27Ql7HXI5jLEJD2nJA20wE5pTDrRn4q4
iFD9v6mnfp0s4pCZbBbp7efp8pk0zZDRKSDdvprCl0EKK55wtZvfwMiwuJJCY8WyaDVFcYbZA7T4
B9KrHLm9skVeT3O1FNAXGQDKp2Qh0hxAS/+YNtdXlCQBM/VREvkN0H2IXAycEjheJaNYQ6JsvNE4
BAiAE6etfkTr0rk4RQlOY65VOHWfYjcmOnL+orROzMdtLHufE0nS6KhRekhWcsa806PS6YMnJ7h6
IDw2vFHY+4B5bzdrm/e4oIQk5UPMczWXEGLw17ONMa6cEGOY7KQeMHVa1Eaatr963rNvOemSfSfR
KkY6Sj6PW02G5LRSqcz0yOgIjddad3S1A2SU8foBNx9/yzWLnZ4yKARaioZAh1xziPpnmzUiaPwk
bfeA+Xv39CSc6IgcJdh346mdEk0EaIsx/fg/l6z/OrVSrZRCjxmgGZkLFOes9YOj9YZVSHW8fZqo
WyHbje74FD3fhieHG+5q6cvvAFJiY04onX5FVTCE+CEDOU3+vZS3TjC2QtWJcKK+Ry2NEbjU0CIw
+RPXsOnpe4Nphb8ANvLLkOtqYh8Ntb8p9uLVsrtnWTKYFXVSmLdT+iEoNJk0r0eS/18/2f9zxr5m
/eTnruMbNnBtKH6/dbY5Cp5OKfnd1Y+IyenXdnAviTdi0pJ2Zps+Zqx9+n3W2bpYHJjAmFh4cQqm
1Y37xg3klyo93j55DX/BBgtdS8H8Bqn68dp68jTOkIWgWUWH999W7to6+qD2MHXPV6JSLkpmWRNQ
oqGjPo/TP3ew/khWzKeExYGKwoiX1mrFm4ayWVigVm3looVLsLdSZvnVN1L8SJ5d6z6qSSvycETm
LcprIp+yamvb9i16unTBl9jM7AcxdiGMglgDw6oasKIjdeOMeqdiWWDGoVOnDxUTuZXdYKhhoNUj
4pfAD7nnvuI4jIlBd6F1argAZ0DGjLf2oLJGHykb+ASz0PzaWlrfIxHxHD0RaITzlBR7Kp6beH+N
jh/bTf4vKx8X5k+Ok/bGTauERugj97F2Md+qSYucAqcLG6gItJwKeNPLAlswNfAN/XDbI0UIGjKG
wd6ZH3R4Rnalfz4OjIA9u8VE+6SBojptl1XEFR7m6hPPYHZbFG0Ld+AbKasNYNqH4AY56AcuUG/T
pyf3+aWaEblhvAaUtTbK8aFidRKEw8tCz3SoWJMLMaJqxuB9oUaGcWcl3iHzTaqInQ98B/ZZxyIl
2Ttgd2dUhXPnqt0E4SFaZjbZQElzIeZZozr7wibKMrK6csOO42/wft0vQvYPuJ+5WVcGOHISX6oJ
XpzihPHOqD+4snt4J4vY6NaAIqQt47vEnURRTte1oP3kq8G8ZlkTL8NtagTdvHDFgjHAfWFIpNuU
VmMaPREq6GDiiAsf9SBZ/vKHF6uBjPVdjXon+TRS+r2CG0Bi9pkkOag0SH347ifgPzc48Ftqcv0i
tFN4f7IiGNRh3D0LgkJ1pZ1IQznmzRDujFbWhGkjXlAF5O9DnUuc88ozgXb2VdEJ+IONunrG8u45
BDRjtIhVQm+RelasolB5tltqMJ6WwH7/zZyr9V23zD4iKJwWFs+FaO78WDvs4wOMs0QVWyopbef5
sgM0FoXAIho3x6R6C78huvIb48fGt82U+DlQQNvnZ8L8CZMfa/DOb0mDueJyHpDmjhwvwmx9ZBMr
eAdwvKp/eeIkD0KEcBrNPJFP+vYBu/6NcdOeYDftGEBPvlWuXTF/Xn4imNF6yRtmu6Cb0R5jyFuK
A1sDLEln/keG/TORgPkga4giS8qHEigqEsRnQ2fH0PoVlOVGurNnEZ1jPbLouTXVinKPN15d/E8R
tcKN0i171fmTK6gVPY/SDkJOMj631CfRLBixcC4K56ZLdEA88fvrfeWOcGnO2eLk4tDJo/3AWOiR
A/wwqnf9s23GfPm1joNZiPZ8oblrukW6i/g9YwKFDkceyUmFtuetBcOedPoTII1iRkk6xiy95Rdi
nCCOTpYHS5lXIi6zBdGUJVczzBrk0Nfl4u5JT3ECI4BNfR4mU3PAZwjRtCLgOEN2wdit0j2tMTJk
hnRC5doiLkEKpCsXGvkxCE+9R4+srDLgCjW2YEDYoeiJgWyLS0HBww732uLjZ9YcjeWgAk51TE9K
tWo9W8+gquebGcCcyNZ62wrHfrboXqvaDQRXxfvm9O/etLaPOgW6EZP0XY5ViYerR6ZwMfALA6y2
xPFj9KW1RHai7Yhhw1SCI8rRLkeEoYK+eT5/GyHIV3mmdD1bN3/ZZHaY+w5S1FyhAgyR9ITrHAII
+46QExvwnRciRM0jstHm8I4CfwLY1FB6NotZHvZJeaeajHtqT1B9nKzG/dvBcB5o2Y642rOd57c5
pH3rXlq18INME0MiGFOsPCp200cwZ2QV4Yh4kalovtL0Xfp+waAH9uOE4DcQ5Iq5Kv0GV0gzFoEd
vh+lLVpx054K8aPIu0fX41qZde9Za44fHfw11ovzqwC/AtHRYnG3/AbhZWAmRIi2dj1C0/AIOSNG
5trd5dEIlX9086gKXdcB3TEvGfL1TNDJpbHuvaCbQ+PPSQ8hU8nUJIVFuHtiRETw4cudydBybzY5
4FZFuMkJLuBKt5N5MCKLYaAqS9iO+SAAqwnv4jkyI6Oaro9Bx/WtYjvmNffEME+kgUlwhH+BQd3m
PptysQ9XRtWuabtomaNQxoNO0JiNV/vNVpFCY28ZPlSHvYe2jaQGYJtx7jqBlfy6BQ5NxUTEJbFz
kYpwdbkqtcq3MXXqMSlt6cI+WTbrF2yKpWgHzT5j2sT+ay0274ncBau/gg8ePs/i7tfqBZT4qHTX
rUmGnQdO+KHqcYluPUsfJq0GXPkZiPvsSrywki5wo2qGGYA7uUcQWf02eVcv/T7ZQor7sAxDlvvT
8WATSELW8IaUA3bOdc3vH28iAx8KI602QZiiYVzJlUm2Fo06kyMF2+L6vhKPzy+peJfN8d2AW6LI
VzoCp89qzLRLfroC/PjnGJ/VHkwx1PmzIkWbti4KrnRFlHPRoCQpuZDubrKyBOO0V3b5ArZirc+1
EHUNFqHqK8nTCs8SIvs1Ikg+J8dwVChPdIvQvRe4NdsLzYrUux0JY3DjIKOtf5um/e89avjfFU/P
zGpi295VvRpB6Wxal809ZmJxxP0BwTALc3CZaWsVfo2wq24KOUl7PbCSOTUcyoY/HDlvJBfUNJ0+
6lYiu9xeubDg0HuCETaO9Y3aMxn1VH7S5BlF0S4hFxegvdQfTqtBdUl68xfrQV54H559/z12zSza
YF7kMym/mg2uBYs0kSjJrjNeFxJ1e6DfXbl3ifWR8KKQITtsjHGIaxXzXJ4IHFgl7WmNS3ayh6Ze
8f2IOgyBc7ghOAECHpe6TJuSW/S5U8YP45nRi/lUqm4Hp86WTp0NN/ee+PikVHMkRnT+xUd+reZX
TY9TlormZHZ7gpwTj7eFMSkwL2NLTLQqU4on+rzdLc/g9HScZz5Nb7u0UTrjDkKG4aeDe7KTUpxN
S9STvq3bmOVstsQ9NEuSc7siobJZpUXNFx7iMT4EeNYMydTWLHdtEkreBNHvO8QCgs9oQgCW91WB
jzrva4v1tyXnU7co3mfVZtAcho42Ups2imEpsrbBvufDY6WQvnrD9ioGLo4Lva67BH9b8mExGxlR
t/gwJorS1MLO3hqg8Z8VZEA+hcXbcKhkPspr1CIC4PYivx9c0XhDOxNSTLTUyChjOjRkgsoYsNrE
tuAH9wixKXkdrLc6HcR5V+UZO3C14kDzTM1yHMagmQQRf8Hc/xUGLZTWja/vt/U+SwwUM1p3WNQO
1qtXujpA0Oj8fxZBNl6ii99reeSWT7e5b6yUi+wbtsxaXNQEE0Iv1CYE22AWxRc/M8b4lb66BtLC
D+EMaGEfyfgfjWFFRNIyxR1zSDSUYbNneRX1CIhbtTkBJEuRJ4nfWNu6H6p5FNqh81fBc7qFrCd/
2Yer1AfIGornkRdYKFRJUWyuqO9A3A+j7FDxmJ0zxG18lFoHF38tnFC6WzzM/6q6dJ11GBYspWGN
g/mosNIJLhMo2DnoFOGHHx4j/asXwdr2EpBBOLuQ/4lHXvuLJZXnrqDqpCgUI462Ijf/3XbOE6Vp
XdSMg3sSqeNq/tng7aqvFv33MVtGOrJZFWtI7MmtETX7okN1kUq9BnCHfnE1+SZGFk7VltGodEjI
/0x4eVfmwh8rtxJKH9zCMedsh2JkAifMgLCWXpk8TvSEykYjJRXBy1U/X/jsosWfL1k0ftZ2LLj9
lGFGrHQI1751D6QmNqc0Bo1evFqzQ+bh6dXAeRtl1Df1pFNcZ10+O+T1SshZyTOkMb2BYxLs0iif
OR6iA7G1i2COWYKfJaYYUvL6nku8bzKrsuQh3AAtCwFMBch4kU8nKIRfQtPElntucXx/csO0Tpft
ejG85wy0xQ38amvKDoIgR2ufUyWDAHl8WLWRvbmA7gDpjlTnpDJj1jxLDCigWgUbgZ1SMkn5HtAP
uhxNt8V7h5izMJQuijpVCNfdnIGelXjf7FROI12oYLO5z6pxP+Qne1JyddwN4riyt/8A0Onltxak
Ao9D4SfJZLS+M0FE91lem9lhQXvxVa1/xTixWYNM6KH7vxz4eNfIow/pA0KnXNKTiBD8qZ5J/2vy
a/hzzc29uAmIpxJ6atOTyEnU1t6bfdBKhq3aJAffW4XrpWjQC3NuK56ri4venrgtwOWQbCjLZ5cO
NTBLIxCHUbUN1S2BCMkCpLfEF72nq2bVwuvl8r7FOlmMxv1SwPp6nHGTQCwu+vfpmEHoMxeRSpgH
kdku043bsAsIDg7pMhGowDEmOzLFSB13CRcPQs/lcLQqD9YzuAocb4r/W9J8G+lexbQa6aH+hX2J
i6pRtvmBI3Zxsi96ErM+cjmOtzxJwQQqhVtkEtEjC4jMipPvFdtFZfvWQKblyvGTRi4hbeLsvgll
YIgxstCPbT+TlmWpBkGB5rJxzmWx5r19rC/0DO3lkZjYgIqn3TBms4zIXHaF+tGQRSv7g/m++FGm
BGlvcAgZxfVn1MmtAZJekTaZWvh8qTBqwRDrTFG7Iti0BIcMcUbyxoUxEhd3XdTOWK8TpZR9KhAh
MugzsFwcnhfcp2jfdjEBxpuxuXFvd72aHmNrg7SQ2dl2/6b2m3DzYL/2qgz3dSurmOBWMNgw/7tY
M63PAgBqShZN2HZplFJMsBIgE2vXT0bBfJTWeKLH9G8zyPQ0wyr0YffS2rdy6cA1D42TiBo4JdAC
1WGwxvOzeXVLgAxNR8J1hiveD85mAWG/pUl/p4shobR/FhC4s9ViYVIIrMN91O6beMWouzMVPm1N
oLCi48IySanF1P3gkFhTwftmN9HSPWs716hI7LaR/NW2xmdz7vrcd9XNGSthJd0TfU8AeSfshxnG
7jpuqdmkouZrliWzvlDMp9UDYWI9uIMfNWLz+4PeQAp3VOO830XnqtemQtIuuv8J/djb7p1vnyow
kFxKV5CrIwIwQ09T6NPwS0lo5Eu5uMzuQEjyvK2Az9ngQEFVjuHgBc4Lp6T6pZlOu2iUcRpansVA
P7lOxhAYB2URrgnOw/s0ytGEet21h6TYBLQoF9JpWFoYSOhcY+vnipBQyKiu6CN1SsmPKajPFAkp
ia9v/SKMewwiXGm0YleigtPapOZeqWl1Ko8AhGs/Oy3ZcblpXpR7TdMSf4wwNC5/gwDdg/5IZKTq
XBsDkzKnXzxAgYxBcyM2RuNgSHcncV0GP8gXHSrE7CCREVg8A8eGipV3NKOub0ORkxPA/rkDyyu1
dmTPhlEPg2aNdvUZiSgRYDis9zNnhZ6d/xHTyGpSlfdZY/98YlhrLKvvb3Dwm2X9uggOslGBCGPK
S7mAx5qDM2zw5Ps2oizXs++KZlYe6cnQu43ETHHjXNB6ZSpXjeW6G2lfsjd8D5S56o67mrqylwLG
J9lWD01+aU/J5f3GpDrDcF87i5jOHEYJTihoMq1j9YK71fWt8u3ujvHvy5K0VZiUx6Yr614W7Qa7
ecjWWNwbebRhw7JeWZdPtix3DwSYJYkfHcC9nkysSCxsXl/hEO5XByuOoFuHwXwXFGZxEnNNqKSR
ZPGrzK5DOyR0HMWwkyQOrcy7mxRXOdD3nHcghmTCEtQsTpZeB5hfj2t6JViNDUMuxPyoQuVxUXDW
P2I6zORyZKAQiVkc0VpSuHgwLPNbaXhPF21zZgAmWd9ukvxVzm7S3wlT1wFV1bC+wGKiItbXYtbH
NISyd6e5XTQZfBgChi0j5QZzpv3p+BZCd4rwaPc06CUFH45DN/D4ha40ZOpwcGFeRWcGTC+rrwhI
waTVDJmxSUpJt3/OVBnRlTuriT3psxQEiQSk6KLTOyP+4pcnJz+SMSY3xdsy+50UEYpkIm0NrM4G
iJjkbS0wvCy9vIrNjaroN24Z3LK/gNItD2BMOeBzBy8txWNBZK0WoJzvrZooJWH43itWcrOZc8YL
qog63knXt0UtmOZkvvU0YOJJ/gbfeZ6YYtT41wewwLbohzJ4lp/phR6l5Uu0MapqLbHW+DN/xA7L
+MwDGczk4dX10sDxjT1XS030BQfQ/d9Bwnbyzn1EifGDzAr29Z0406fpklo4ESxkZHK6WUMCeJHi
jS/o62XnvkBe2MiCaCVWhTa0GTbTiz0Q2Obdc1+NjRWlITIQ5XQ3yTQ8ZdqVy4XbFzZ5R/PXzM2S
c1zdc51YWWN7oqrhv33UjQEi9/WEv1b+A3QR0YHQt++4r9pUnCOqwXr6h1c70fCFcoszEQK4KM9B
pOuCwRnuOVWQq/cBjhOefhrc2uKQA/9OHGo4OvkLIhAv9jRCk24oEQDSzhJQVzG2rhWioZlikBQo
Dy9+fxpTvYOtLKc2DqGSauz/y2nAmBZyyz9tkLc8hkMWTkn9CvSW0csXm5CGol6rI7MFfTqnWGGh
taCJszhy62H3YK/yv3SFVvnTKlopqscdMkl+ecJWYtBTkmdK7L22R2/WFhw5v9l6hZWL9+Rkkf3a
8V+HfPgvFV5h+veHn3WJBOa62GABj/hBoOrCPEPL0jYoLSsBLYYql+j7jOMKso+Xhfh+kNqdBe2C
HVeWL71MsZzhzgrVdtufWkH3UFNgugcoeN5Dym1D++x2QUgXg+sK9kZO2jJjzY3HNYaZCwb/34Va
uT4XbsQlhtTrj7ySS71Zxk45iGHoom9kRhT2Pbat8rxYGzpNbJWOkk5jnBnGoTMFXawJ/X6LX2bk
CwZIrluUURwh9Ubzwj+asBrrNRt7q33J7xltwMyT8/iGF2V6Aag0F6KTnU1O3QgqTKap6ulRLy1w
+AINSnwQd38fyz+HLmD3F+fHh8V0Q0N5dOx01bpx2hKYo5bBaJiZyneQkdkLCRSxVr0WqWWvFK3K
zuMHH2vk9RF4StLI7n1ZYF0q62kNvrAr7WnTf7+bhqkIOWEPSRWeG8W5gWWHXtfnHu+toZR1Rh6e
Vyx3Kpzktv2ypIfazBTq7HdhNXT8etDTT+C2sgBVIiibD8OprYju9Bpa64Aq8uinNUnBpsoreTGy
0M/4SP+SRZRihKdLfJXJol8YamIXTdis4Own69QUih4yTgqthRnoBgssJn0X1ZTvBanjjQQUdYNz
pRtOAWNTtM1OdJGY9DhnXLeqvVAM7lZKSzH+2MYpau8qFxFJWpXCYI3d7ME0G+LUnSAsVNbjNNX7
x2jCABPLsAKMECycn8KF93MX/vfven2kkQUMuweQ/TkDfPD0bWdiV1LkV9KdqdMTh4s8I3huDlP6
oC0wKWIPDWgy0w89Sqrq4Lqldi/90w4iwUmUgkiNK6UJMU3SJs/FEogJ7yDPlsuCzG/4ntrcUs/j
HY5cPE8R9AHXTdJ8ntxd9mMhwfkGGVGJr7lUhqceFyp9lyg1Hy/TCrCuThQ2oXsA/9kmE0EPjeWd
JObhC9vkJZ2NbFRaJIPzkTCWiapsKx38NzLVYcrsFKNYnpu3s9UlSF21oUUikMOo/ohAceqDn4KJ
53ohx+W811ceKm2DrfmwuUadK3DtYvl1HhPmlVjua40s6ZM1TXr0ncn4eTykDjJAO81ZQEp5c11t
222HPNLtjnu83v2oa7q+JikOiEue/iMRlc1jehc1BFAPF64NRyUMDLiMSljoQHHMEGYKXe79TCwJ
qWKtPI/rLo/YLUdWp6HNxv01wPTfYxVG3oCnEi331AAO3jdNxZqe5dJTBAdyqPCHMitaDzRhQykw
pAnbgmJq+vLTfPgP+TtO3g2Rt2yPfxnaI/ZM19JFyA8qf5NYahSW4+ntqJooJOenpRnoZDVxKMn9
36PX7mxKN4KBV07a3F+pFRgk90uCWM6l8odsG9c9MXNhfvWfwWSIW4/zqXkBGiWmkzn5O/48ajPm
oPh1NabYuxpiG6ra6IYKm3hHh2OglUAAGP6KI7/EmWhAhHfGY8t1K5k77TMHTKcGXG+NmaXUhLhE
nQ5aZtj8mv7qQ2icK5ArjAFHekoRKm8Vd9slvgpQI5FLgsqj5HGCkbCOBXSF1IalhxZnvB1vFwfl
Z4jD836R1Gwmldh2hdT8cYP3A6aw3NSwj/gzM6N45Vryq52l6/sy0T6f04XGkECZImx75cEQcUxf
mYGgFZ6xviyk2x3YDVltqm2kaz+B/ZXquQH+FeMfEwJ5LiMZ904S3DAJxx9tpCLuvg6XoSXosz8R
vCvc8eOfTzAIU3wqkkyLZ7leKj5+CABdQ4v0MmiXZG0BdSzDEFKN0WNOuvGXCo9Z6W8tiHds4fqg
S7AhNyazzawfaBpPAmhBdykGDTOjG5ncnlMnCfzgl7aUojoozUwNFy3UIBq00+BtwNgwUlamsFrU
UAXnYu3Xugvcw72MEvRn+aZDlLDDn5EfoThxp5yu74DENZRIpQOxP9qjE0qK/5f617jrN9btNdXG
4QLMPtO2A9tLmjsYC8p5N3TvKcpbWfDF0Tv25WxgxiONeHZP8wbN0MSoFUnOXSKTLXSRE3xZwrfh
AC7c7li95kMTzgEiPHVSRQR4WNR+JTki6K8Ecwz1tSDFU8jO8MdKbXt3zSxFwnqKXFT4c5PrtlYd
YjnOCrfF+Ww02o2FgQzWb77oIKQqk+iRTvffaS3T5qNhgzIxmwZbNt+d0LH9Yc6gz7fpb2V8GBeC
aiFUP6ZPVAWJOCYbm2277DenjJ9ThFhs+TPYNoV4PCHqlWZVpleCV0GjRFDjjBo75cN/VO5zySW3
DeDHxEVYxG9elD72By1TWdyyF6Oh8+Gc/HUKrA5yU3Sv0IW3vFuq/tpXpDH89bCbivY5VWlHw7Gu
bN5BuXSzUrponu7ewHtBXck9b30Ahdc+RW9+u6MKWkkkNvIc6m2o9qv+o0vnSu72kSvvFoP9I/s1
Ugs/EHKQg4CrW0o5yhlCXDoDZt7CCyFpo+6AIu820SM8xcCjQwlBo00/Ev6c6a7k/UZJLgqQ+BXi
63omdAZ3OazyUQhpw7473FBlHbv1a56OoInEW1/RiEd+UPD3R24YLM/dP1YaqjWkAL1+gJ+Umeah
nKOPu1y5t4PlOO9D3J2Q+0FCXCvNlDW5cp9WD3BLtPPVTq0psVJfoFzfNNGlv21Ru9Zyc+kwzNsr
I+IH7Z0LsbSAN+FaAhapDAInMzzk3M7GpwpUmMeh3n1NuYPU2wsxbQCQ/NWc3wNqJbBVeC/2zqli
eQCW0MiQemS4SZ5k20MiEfYpldtgu0smQDUWLBU17vYnKzcBBbr/qfXjOIERcyZEva749E02YNwd
bg0wSSGKNbLvpe66lUd41CytgoWpUk9L5SAumO8PwurFTPLc8NKAr4GHpHQN0N7JcFt/A2CNyhyz
MIEE+tFFEcXqUL5ewKwGeSZecAjtaCrs67SeauIEL3gOKHt8QGrSY2YU+79mqY915xIjm0heVuwC
2N3tEk3rr9nUgpKBewmz5lgjSDp6Rr7Q3ktYfmYld4F6VtwlJsoOahHyLDU+Gu4QTOK/PW5BCaTb
zSYt5cMcaNl2Cl+bjBdBQc98piOxXP1SXcaGzoyW5fYhA91shWfxst2pUzI0HBx2j6J/J6IYhMUC
7sRFsXUSfjiKLZ0PoOmaDPR1WZQC1jBxwXUNTd0g6RbwY+dOlKgcuDziXYxq2RpLN6Bh6SapKo0R
riYfC1ihWO33aWp+CXG7pX8VqK/BUuzyznwmfclTqQpgMk2UPDaOCviXb8m4rNaNM5bSTCDI9sfh
NJ4EIzogUZ5Tskj0Mljn0cK40zgwIj7PW0B5o9wuEQXhEY7q/BfYcpIV/AN0laoPtxQkQSZjJwzw
CfkwZyxdsla8fNfjyKEDVprVfDbHoE07lntBayEwYBYZV4rUbEireYhm3EfPPWKpB5GCyxmPZd8H
2vA1RW4LVzvOV0NMrQUGTjc4Kj5T52f05FVNNuHwLcPFO/XM/J4aKSMB0yYiS+SG70MPYWHv2g6e
Y7p7WI21Gm+TbbpTd6TLLOdmX7xytSdhhXkBGE2sh8hyphac8FmnYNdsMNs6SNru6Zc3NEqz9nns
NrctkUfozb3bMXi/BRClnrkDP6iq1Zrc6X+NXDOSWM9rB36/XjhbTxHZKGak9ZjGR3r0lgai0GJi
zOOWVBxKb0cpVY0lokCDQ3FOK0JPJeVJgPY0Ws4uuQv+hSWxNGRpr9KC6Hhw84eCq05uwJgQaHw5
AKjnsifOt+eL23Nje+MiDYDmU+VaTAdOLiLfJo4jQNRAVQUMPAergw5nb3xjr1yC4JHs/UiHh/oU
MnpK+Thm8C3fsE4yBpyTrhAnggLGvca/DplIz33yC+Z8G4LntNiEJLStORUY818RyfJBTR2CkOeu
XWa2SZSS6iDatJA9vyavPPlri6QkJo4OSrJ06vgBWD4XpkxdmbF/dAuJgC8jfpxPNrjyzYZ/6YuH
QJw9HzhR51OnTZOQvNTj+cuZjF0+ggMIWvr6yTEgKkEgbDtxKA5JiL+jud6cEKXY1RtxSL7OEHRd
g1N7WWTIvI0KH+qRUW42aAaESenTSFBQwcjerFmBVmC9lX+74sfg9imZIlc/2EZ0YRxg5BKoGv+w
11ECJAHbc7xtmdpABadMr3McMPzNf7Qh75bQFFzqCcMviA51rgkIxoLRvwVuAsbOiqkdoDG2zxNg
SKzw818kwAN0vaqcrBhhCpZ99y8y5//Pvpdnvfz6OkTz9mDmFnjEfn8EWy3REXrOVuHKbSbxcxpY
UuuJua/fJJ3Nh7P+iFoJRkmN/pj9LfeKMO51bjKnwoNc97/KrytrvLLWH+3+aMu87WNuWnr1IaKF
PDN3Vfx5lpk7lUtHrv5klsCBd1fN+5HA1VF3ieEQC9d/+H7sQZx63ipc4m1zKhJ0ZCFnrQU4cdjw
FAXax92a7x2BtqjCOqgvyK+d6N8MMi6r9akml2HDxZSKhkqLrDUvCSG7VOHPqM0YRLpVYwGl1EV8
u+vLtxLQWALholQyX6Rp7FNIzSU9zY+IFRVD690mMj7e8JeO46zY7vMSA24AbWd5p0cVd1En0Syw
T4on7sQpwutS22OEWC5DjWCc9NKHev+h4BFhZGDUnNfZAVi6fL7LwLndtKTayropp4Tqdg5eR06D
ddmENupH9vS2mupT4aBQl2E+yuIp+BaPYebuPfzKZi7Dz6sV05tWTmh+PENKbB6jlvmA1ZePGltU
hquOBxdocjR1s6MfJbzjOuHfGv14NY3P9mdR/SSy43ZGB1Y+a/KExRt7RDeU6k5PF9mwK6cyNZAl
yxSbqTnb5O9c1a1Tfde4YJjMVv5E8G4Z/eIBxHxYT23j/ou1idnzko80MKjsnXI+4adIPzy5s45M
6xArp3GyTGl+j6jR+e3zmSGuJIUPNWP3hKA0UsKGV1iHygamkgT6NsJkoUljQl3rWPGqRQK3Of1K
/0mS24Rj6d3OWl+G2DZJwsJzr1KD3OTlPjW3D3zVV/N+LifGuO+YhHEJUvX94lv0nn6Th4hnuqFr
+hNUM/sd1cXCEPhGMKDMGokk+mmAV7zkzEam005FlDkQNZ4kBheqiK6oWQr5iuKChO648PLoBi7e
z2nM0UhWGA4AqYN1HExSqFcWtJ1nfijLBOv4gQ7PznxnmQgomWhWqDukiWZBye3mXhFr70873O3b
Ty2c5By5XAUFk/xfmX8aqbey+gzi11NYsD2NUIEEovDFk8bbxWGT5e0TKaqZSxBfPwVlajY8l3PR
OodVrX+xJIy2rMPMjt/SAeeOeHHpBLiTzLY55emw5MLPpJVBJrIf0zmgm3opdxV/KlXvbsWvSBdn
/y2hw7B+cLNFGjng15OG47VzO2cW9OCN+Jssmzoj8oN3X3IZwICloSbpgG5cojuDEcj3iY3do2e7
OsO+r6ZxYNZMDbNLH3gR8n2AA5i4FB1525p3ZwSa2IygBgKeNDUGnNX6PM74uXvXyiJ9YQLPngBm
I8P9WiqcXRoBEodyHTMjpQgLHuz7xQ8RsptwltQcTi0NG8XdMYxGqjEHZk7vivtYxwoCzKyOIPXe
boWQhiH7o63z5pk6RbvWfUikp6oeWXyU0LYA31rQGgqn8B05RKbiuPuXiCQ5J7moBHT2I4Z6MNKz
fu9O5VZVMQ50XTu9m8/jzfeufpFrE73Cdtgz9n1mjDYWrv0ngg1NnYTjZutZhOzrurUdHn338+cB
D6HsJLrhH+G0HdDb4UcEUL1hA8qAs9QnHaj37xh5NOol+uxSOg5LScnaqh+AMpjJ0fuAozHBfCKw
mGPRhvTCZhjhrRWaSJaSeBKihtAHx17CWp2UpSc+mnmB4xsro0V4/qQqBb9hRu7QTrUPRyZfxv0S
bj5jK1+ffrZ+17MWMdPtIHyBXzVrUxNMRQ50710x+oNVYILdhUpAHe2mQny4WhswW4aLVsbJyzLr
t9uqAzbsT2iA7LS/mApJiKZpIDvSYJxeslhoNBtKBBZ44eWOvExe1nUPio9AeqeRuFgI5PSf8pJY
supqR109ljWimKSdXYmp8qhCS32S4jZ36duRiIHhRepR++skUx7b9l3dbDBm0qI1uSWat6Xfqxmd
XXEA82tnGN/cyIrEQkLGjml9+7MmyxZ0lQHQmPEeHJdfz/yIvQdhUAZ4+pDRQpWITeaY1O2tagGx
5aMV04P4eMcc5NgGdLUAVQWodqiEEDHlDOoWuvJyf4pIuiCcZlgy7D9tYLLaU3zgYpAXd3tpVw4d
+qsufvE0QLN8UaYVKnSxLLfEv5EW7Sn9UwYtPdFHfWWLtIthPvdDtiK+zLfVXL0RMk4IYlt2tz5/
bc5DcvYEoPjb3G8JcFzOTazf2SKfjVaDO8WlKsTC2iAAaWg8Nz1xIMHblBggMRc3l0mgr7Y6MiyO
DE1C/Nyd4QKeaixNvURJ1G2NGPiOcpOnpDUx4IybGnlIveiFQOdZplXITgfeNVl0CYCBlfoHUN4J
EUZlKv2FBvgHP6AzbtJjYUq+rZT1IUq62XD1HWDjOOfyrtVh1U5DyzoizhKsBiehtbGFD1DN77WP
jBKdPJn3yB8PWa5hOI0NaPPLvuedcPxa1qjcGluHK64h5IpfwisKWxz0Bbt7+MROvi2e056yEH0D
+wC30Zro9+gs4WxjIj/H/EJLrx/WBkD1DNO1CoIpPMbj6SgiFT8b65+GlOlfEKyIcviVtKMJlkeb
rCvuzB/HopaadiAGXhnst8bF6jeaU9/7UezwhhQekoRSt6D3CCxATp1a2FN9oqMDNdPnDujRXXFE
6bdBFa8MXf4QDUc7zP73rgEZ56VR5IFrvhmBKRZiB+gSXXPBekrhhJQh2o58ReD22nPMtxdFqJ2q
O7itSrzuBz4ULDbmUStmQq4YeTrc2GVs5hDWrLnK4hvt5YtJbGGeTIV78QAGGB4Q9y4ZOmLGa8ct
J7yKyLtySWFKd4bd+W7NCHi57mU5c3uq7QpIW3L/41bZTY2Ldn8Q/Xsi2IoVzG3+bZbaHdJjo4Zo
YMHDt6dHxToZJ0UwYyFz6uMkm87q1r4fIggAr8G66xZfDzv4ll/EItX6nzBSYsc2QlBs3og6g6dW
I69TnSy/WXX85twKFpwaFtzjikh8jGlx9tEm6bflbCKbkSjcHN1T94AYoW9SdZKD5SRw0aplZP/c
BMkgzvOtl4tmaZc+575DTyejrM8pag6QGkMQGN3oe0gypduE/EaA6QMy4xzU4Td44mUrwsz22irX
Cae5z3XfMgxk/6HCFvCSgaFb44s/K2inLzKkbLv85Ny+q16TyrlOFbwgiauBDdg0fqCDyiBRenco
BaOtOmdNaXuoxWxeCnidOcA0wpmGVOOoV0w16b3GT4GPPor742vfRznwZDHm0cE5W6fy4l7dUD6j
oHC1/yVjAwAPDmyc8dpQwP79klgP83GTDDdHTDyEJYesbZ3E8hAID2JmzMFYM3cCdFFeU+RDg3aW
/fzcgO7yJRTH150CxhrxasBILKUlVFnwjJm+O4roWKnM+VMVRNE/6R5tMDBkzU7FeWRjJQC+cmAA
WHnRq/72ERkr9hV545CCNDvpbpq++D0wubMKpvLHCcySu4RUltqgTvvK5uSpfdSJ4dy3sigbhYm7
2G7mV/B1rFycmR/4cQ/h43X4yKeOf+3rum2NrOLS+6KSfds/oMHLC7J2FC6wyUMdXAfVWneMEcxP
OacYO/VJco2H0/wDiiUbRiximye9JBqicaN3x2bfIy6Q+os54m4YQwXVrHjiPPmPxL8vm3Ei5+Ep
SRW1enSvzUGQbDwGvmcnBRyWMRBv4ttQWmaB3jya4ArNw7x9/U1kpIHEDF6nA7CRUrDp0sdD1MS6
b+s+d/OFOOlXW0cOIVxtuZRXTgVABT9uUR/jRuMipsVoNjlwMAhNf0ueVQ6cB/9s+rk9ex59aqKB
N9x9WOQv02MH9Kv6ihN9FXiIhGp2P2fZfeJsTKdErIzF1tWKnqLu8fko+CSqBe86dcnw5M6c3kz6
/saXUcuu+bGpUOYpt0nRgPdnsNgL5pvdRx9+B4mMlD0N6TnBX/dY9Nc2tqr2qIhPvD9FBXc6Tunv
isNkSeROYJ+T5x9gaetdR0osclAr/U3soA32pUEMOVS6P1ApkS4UftjczvrDp7HZwkQakKPPSbWt
FsjPDDz7LDHlat1mTFsJvymMBjyn+5uYRfTwODHVdvGtZjtktGl3KK3Ta7beZF2Fk8DaCntuDoHk
EGJLhmUmVWqEOUrIXgtOl7zicR5AmUgcvt5Csxt9llmfGgTT3cK/6Auon/YgrlyG/6uRchDfPfZZ
y3/91zgCe6hBoOIKzPUdWk2iKYcotPFsnVjILYfVkqgaPbPBrv/Y9PYA/ahDU8sp4b59ewy3+6A8
qGlD5QM1PhvglVeLv0IHXDtx4EUMRk2YtnNVYrLUwktG3e0JCmrsQEBOcoUh4VN+F5anNXmyuzjy
aOBERGy9zc4uuh6Z/qWPBK0773wKnYjaMqa+oCaZRQva7D8LCK2c1pL2+N6c/uNBJGp8RAw4tnBL
XWuagSPCr6D4da6WPH59GmoYXAQ58ITTxQOXShsXxNajjUio1asWoppioPxRIsOO+0qknbNLiuXB
3bUxysIJPFj7IHBhIAsZYypimFhTKXs2xGvG1eg54rZyoRYu0IuGHnwlZITcCfCgz5Msm43jF4lm
L4I0HsOjICcCVvr0Hm3zy9bTolksiaHlQjyLQtB9SKaxLVab+itRx0TcdPDJy1YigQrOI9uSocGd
gv9G/7U2BVv2HXGxaf1NXG4PIgnz20oeGnUngUrUNP2Hrv5SVO7SkX7pqCCTeZr4yocuZ1kZ94ib
vmCzUg6JaUIRcr7MY61JjnY8mqMgj0QraKeHqeMPoqbVnmWEFGJrRPvxoSqiN4puJLwO6uw4LtFZ
6MTJmR9a5j2pQf6rhpocafpd5UcTs/wGPG2v3ZO0Odgba2m3zsAwjP0ptf7IhcE4/7HCKPVSjmZb
Hm/pC3snvmnrdFS371VogqcZhHvl5Rpilddh+Cmoz/gefE/vn6xYfR+9isyf2ONMBdfG9JtiFGvS
tcJAmMIlOeMkfn+QTtHQYIRJom4syXlyqesDGZixxPQsAS2dJDuPL5aBih37ZiUMRzc8FMEuCXsX
4U+VbJI5tRz2eMLVx9rx7zLkkSM7EOt5Xp3Xmx51CSiLMG+VzmvK4FM9kQZJOSJ6k7vZIBhLT+1+
/xAL+Da3VQL3YxTaEx+CQq43vcBakJaGrfBybvGcnCaSX2KaV7vdsiiyBji1jnHKFMcSHHprjcZK
ASJ+jyX0Sd1GWsbgfHGi4BaB5i+GmhOJl2fM+w1yIxO8U1PmsVfHyziV5RHWtUfyxaPBcDO7a8Eo
vNvcP9tA8QTLs2b0bQgGaf46m+/czvSpqtNSr/oUMosrpZWxqTdraZsLBCE5wddPoc3c2bGvcEAm
wN6H87IoxZ27I6C3a7Osb8IjZsN7KUG8QyX9muaGIcVrC+EVy7P1D/QImW/alO59GqdbouGhwlFz
gEeJmadjuHFYddpQ9obpTe1j2/H+n8rhKNVJL1emtSn2n5Q1ENRCv17WBdLph2k82/C2zgzGS9o2
XiHc634WtM2EeeqedvSOIkte3NoH/RheQQ5SFTlyxA5iM1OJO2Oya71TaU9f07uyjwGOYsgJlPRd
npp0juVc7rf3WhZt0Ythx9ndYmX/yUnMlOb3MCECNdIv8bOixHG7MA1tqKLND6BePVOBzqeBdcYY
TsXNvKEAE0kML1YDdCDeV+pA3wtzhKd4DzePCRYFGY/Eiae0f0qCBKBGCj/nJ9h4jEdQ6lyXYaS9
dDqw7pLfE2PJVsNzCFzAlb2afBK1wDdVoiYlXi76A62BVNY2uL7fB6eZdCdYLbh4IVTvq8pHSXW3
wMqwNKV9Af8kL2GXCFAYFK6gC7KG+hAUCYgp90Y2om3OURg2qPFCAqks/nGutdVAD7sQ2GGESDyT
LFP1Ari+3vmXU+KTY6Uq20vviJDoGBnQZd59kFKTrxB9hn2DjEujVbpIj1AMihWpWYozCBxtB8BG
HpVllS/L+I6AjiM/W3NvoUgSqzkv+8xwZNcBt6FWSncMA/XDKUp+htYjQYpCLh9E8HwOPDydSHyZ
WGhiIktrcTbUv8+fV3RNbVZQhBKG6Kd6sMGT45xzRHAGQdrtSLqu3csbcS+Q0Y+r93+jHRK021XT
QXmbJAHRPzCiLE3LReO3E2N1bIUr5TDAzT/NUQb8eeFcLYtPdPmW/xR8HPKG7WFDZWZFG/G2AlT+
MTi4Aoh3P2x4XqrhY8GBv7xB2LLXUYhLh1GCQIzQNoFNQC82bVh1Racz+rvys/XRIMRuFIxpinYW
5lGk6ggpFIvEehFPhH4ZDPnVappXLYGRXgouGLbkyp1vFV/KWyO64GsYkuqVVwJJAluUcHp1sjIn
GldAbmItgAvl7puS9v0gE7t++b2g3E32x/XXHGSZQuXpF7ExG5RWigLODQWoHWnmIkvilukDZU3j
X7649Kg/PdP/3os2zEQgQt5JvENozJHhpgzVUCLRUr71rOwNK1FmL1Owx3D+oMrOQU1EU0x7muLw
+zdQn9nZwLVzXrPmyYBlHZWW1n5zgEU6HJbl1JmEojqcoCOvRRBG+vyc1R2TGf0kepd53+hOtgph
B6B3Cuwnx7xOvEc5euPgndemAClMku/mIGPt5uTC/uIpyhrubLFvQdW+97v3QcaWe/IEAkB05wp+
+ZC2jdaiY1PrN3+06pxnXNqa73itp0SwQjLiW5HAIkk+yLjRRtd7BTDzLVYRmm2MlvcMQBmPIP9z
7xJI49Hev/q51H4g8crBR0KmU44A62MuG4MI80/WKMtSvbHozaEN2onB1QEzwwatvMIO7JLdy0TF
1YPwXGjNZw+oxQg86LhKsqGRO8AVpKMqgGO24OoethhVgLdr2sWEtJPSb3o3moqLfDVV0SmoQYHw
qnb55+gCNV+CI/b0fbW4CG39v+4jMHmsS1x/d/H0gycVD7YAtvIqVG6nAiGRCl8BnWGE3IoSfm0M
jMe3noZ7E9cXm9czK7HuDKmVAmGiaJnAHNsSamsDF5FDIT46IjsGhOpcayAX9+P50WV27Yir/DKm
OPCzjBq5GvFzoy1wIrLLAUH4y0EhQMIFriTokE1mPaks6nLdsc0jn4oS1fXWA6XwEkyJX/YRtsO5
tE1KEE31XdHupqv2Rw+a2RIC8AUr5tZSmLUef7444eoyRdh+JqMpSthBGna7vofhCsZfjKttY/7B
+owcBcUwfUGyHhgKSZW6e6OSEUH+hIinGUZZ5cgM4yHPtIfK8pZVm7Mxo8jjzcFJSdXTEO6hJ9Jf
Ebut4wbqCO2w+y2tc7854ITMEy0OS6WJgKZFZaHLOqg8qu+5BvEhHtiq0YkLvipqHm2YfDemnzUA
6vl66u9JMXhlGy0WcCEJVDh4agBpcOsI5EE56HbHgE5pjIhs0lAGPqkV2QP4b6bUzB1x++wwsiUY
VTk4UFcG1J+6qbYoUtixXj8bzsj3uGkuztKx2xAEzpGOApP/g1d6YGmr/ge+FCuWGxSRct8hV50p
I40T2SwMDzdYTB173GBi1XnkJPzFqCA+FkMNfDO3LOp0rHiLCxi68ltKBBHA9BygTEov4bJiXoJH
kqWSBQ+EpjPbSCeslKkEix3N3DPf8voreBaIJUmhZ6LdRQy49NhhJtwEGqvnRvhYzvDsXreHlHcY
1ShbYxX9UHh9Ileku18owQyhMnVtL9fu2V2PHFlY3NEr7BXJdYsb3hHysJfy4o2ywCgvjkfz6UnS
YMnwE7tZRoZ0Q4+qKBbXyBgP4eMF39+TzE2fVhbCG1kdNR0nUuVY4n+gVVWZ16EFebms4jqq7FY3
UDCHakd+Jr8SpXaoqu8H3W9j8GImrozWQ1kbeLr0pyOZG6R4SfC4CIlO5EknaxYlJZW7ABiRuO8o
FXI9NTBQ3gU4/yz4feZybtKCp9Tnqr//hBIXFhmwvdDa9G0TJcjsG4+wGKJYISWJyWImkMYyQ+bv
ZpVWYD5Vx0PF2RwI8vfXKZGFsiJLSDlZWIOGmmp0eVDrVL+UiLsKJI8FFjolrsZhbBm6pmjUFDXN
bObdjt/mzRxi55NypueuBfD+uwJSqNGI2paJNz2Kxwum0tU3W6aHBrZDyM0ZXx14DTn3bJgskzwf
dLXSq4olF96uuIYKq2D2bxC3/XV9aPTFuTMzdWoXZOeH7bJHY2cJfZFw/aYAg6RDwcijS2GL//JB
cREIDtunE2QsgvSCX36x5rR9+O+1mWohN/Opdi5eWm3xLo86IR6LqhDB/GEniNmZUNecSDXSqU4X
gSmn3ceZt19nla3j7UDWAEz0Lu8qQPmzOpyrKnH2t/u6Q/Gj0lnIT9iVqhvMtlIvpnDpPLSpoRtC
HCkuzKKYYmekYFS3bhA1vjhFfctqvEmrv4LG4ukNpCs5Iu+k7zdWZOG22UY6NK0NuVPQ3TV5Ed0I
erd/cm2+QeQrFU6A4cAY3Sx4xbW1TADU4dmZ3a6LVtSXzujyWHayGvEau5/neu+rY6kiWKShHAkx
Iv5HRAmcRsZaSQzqAwzgPLX/rxI2p2nnTkW+zuC7Q8hSYs9r7hfYk6U+nanvt3hPZOATmUnL3d8n
9fGn2zMmzAmG68007wFKNptADMVbOwwiDr4oy4OHSO2X3swQ49iuZ9ZO9uh/MmQLEj8D1KR9Z/Xq
Pb0r21oJKB66EmZc8EzoALmeponPydI/xc/OBMU0dxlCiNmYo8wbQoCO/i2zbkl7vqg6mGkw2zO3
HlIV2VHNMuxT2B5LYuiV7wACt7MMfclVJZl/kGKVo4ZTn5CzZ3ecsA06akO+90Husa+xDAG07+Zy
Ub+WjZLu9y/MnUq+Zop5yN2NhF1gpdGyqrc96SgiU1tC8ambO2whZdl/7q3w212iR1nw6I0d0VUt
Xe0lIzbY6KmvGxpqd7R5w/AmoeNZAOZ0OlovJhbsu2cjKewMxgRhrUYHpIG21NPP0h2XL2f/dLIF
w+CByv0nEAjeDDmBdVj+4nIj/UstVnP3zwwO5AsdluzTmdplkmdrvnWpdorrAxUMjtDSiHEzc4dM
v97RI/i0mj3S9b5NMqiVCyoqzhIBVuDaIvaZ85r0noKYZfRuPFfzjpdhGtTBQj0RWW+fDYDSKE0Y
A/Sf7/4QWmynVH+EZ0kLGJ0oK503UEPArE3rCzfOODpYFR5Xh1I0K+mH+rEIiQYyV3djXjBzjrzJ
aEdrqtgrg0XH8taSqIrZ1EbJAefHpca8nCMZbX5DKQsB2FQa780lSaw5+y2ADQ89FCc24xWwOuSQ
FcvjTaZUAu43BwZx/DyV61omxEsCoasz5VQgehB2hg/ZfPWAPqI7dU3/wEzQHzdm07dkpZxfF3Vq
qSA+CmTjyhXYlsZKHIzdFN9ZONA6exhhvhELAv3/YIsDaouj7QXDKkqm7WhmN9wpyIXdLUg3Z+Pj
8Vi/dQ/DuXcJoxiWiNJz86H+kEI5iaSA96yOeRt5bMiA9EJyHWJIPnz/Ca0TkctWIYTo8V2IxRXr
wdJskv/5J9wHuROUMCtN4zy0iF2p3nXCd6PtTarB8Wj+s8q+lY8BBgyFw3+KgYxif+xHZuozbd6U
qr3TQMpJgT+hfPI1GaVzza6Hq38XPKCnUS+1zo07GcQYoOelsgPbHvZaGu4WVWcJjdXvhSEjJWq4
x/2fJpAIb8bCZKAfHC8xG6BHEEboSYbon8QmOxqI1qbbWlHQbw+yGSJQWSn1261S+TqFiQIUwDM3
f3l765cEYcnOOZE6imhdbJ4gs1an/QVxnSsjJZtema5u5+tFT28XiwjPaTlXcYxEmRiHlo3mOS8i
p1u99BHYEApIR7OA4XIt1917U81MBBx+lfeVsdB26zf8qufU+84dDhLSye53345jXBca2U60JAPj
F/JsOgA0ROUalx2JL/HhxIvNxVb4JdQISHxdlxqUU5wNRATUTQ6LC0o6QqmMh11n0AgsIhhWjuHq
wHjyZKy8ZKZget47Px6fXiDhyCtXaUdnp3kGKAesAXM/WqOnGi22EPkYY24d2PAACbJIIABOY0Q+
tIJ5uhfWGAqpcHfw401bVfF/vsmdYyz9JkaWoVmfIDGxf6Pnuf8bpMHkl7LlPM5qAaxR5LasaXMU
RHJheGDavuI82RXxAf58UF2ntIc2+mhFmX9dKoxCpEfKEdGUcCedSF068xMNKESkYiBRx6NMpUL9
33Bd8ayOnVZft9qRmmbMJ8gLx8wlROdmKerk5/hn0xJMNWMCHX2jgTSvCzmWi01jYJ4K08ULFrBp
/JT3KSeRE/EOEYg5EsLZyxxvOqHu3/13ttMxP3QYOZhZgdroq1d0ePEmhJtr8NtJDaqn9eCb2RRa
QpgIiX7R8bs2hexSXQ8Cp1PEMbEbq5PW0hSK92EXKJyh7FWseseyII+5/AAKXpeF5MkVa7O/hM7f
082/0y9E5Yf5MiBqmAsSg2LAbvJmyhNl2aW6jvaEmqEpE1j+2vjllREYSWvJaGA7ANfRrFYkElaw
yYLDiPpo4b4FgFYZ3XXtlCH7ZnOO5Iye8vQz4iuWAdYLqB0WJfH4frnjCzvciq/95M+62wcH9PZY
VJiwG3lB7HaHx7GkIdtCk6EIis5/s/VNmRkIEl2ifL7UVVLF0oq7eEvB6kVar56SXaB+xRdwB5BT
ns3caM267tYf+czQyklZ5pMs2ySuF4DiDwjRLy2er4GfmzMSjcOLDWvPgH72xbr7gb5qK4IQ0xN2
tRIr1l48GCdDYedNhY6cEfA32YUjdpcINF6cW3vV+RsZksW3Tnh0jKG6/J4SYJdUCfAquJP0XAYN
g6XXqaf7ZipRVJVEbBbPbiuMTavnCflPntoB8IJUMrk2Zfx6rfBz47BxuxCud1/VH3PsezmtKT2j
X205/C+jXlvA2LBXuuxxj+SymHFTI81jmfG/dLG9Jx2euPhaCpJRCu3aKvgI2IHgyCBjo0391L6N
nIzqIox0wdIqXP+40ptw7NmRDKvtOfS+at5jloeI2/sS6kQKwgj3NHqC9RwLZ9Kv4E1F+KBOEpnx
QVGZtE41L8xBOZ6QCC0pAUH865LSHweBZZbw5Wst45odRf++yZtOOW4DS++28xmOseBsARjCLSFH
aIldQTmp2PnQuPeJHwq3ciBc4Zs01mxxt5BTwyHznO50yl/U8YAWpAtosyNQ4kWon7IdGXRWwNwn
1XupyjFugazKrOx/DHmwZ3fSMtPjKThWVPcKriMTBzXc0YLcinGAU0Ppd225O1fsJVktxA97f1hc
eTsrRSbeKCz2RI8zEJ+ll13bAs28iplPDMtUvpQc6rumObk+ex47kuS7H8tv1YltDSUnroM8IAM9
LUTJM9Gj85P83Fg+42qYznNBeI+4owS48QC/f7w8yeHJf6/e0sfnbc5cy+Xoyz0KD4Qazvmehpq8
gYnmJFMjZi7dqSPUKhtuVVTia+6K0e+bdBTfZHf9cSgE4exadGPJlRwjvM2Xp+ChJpWDXTNG9lKi
ZqISj+mDnWAtQ8JzouaGwXw1XxzgKy9CCX+uu0y110INVyVHrEyth2/DG/7Hnk2Ymgeapicyl3oX
mH534Iwn966Of3TWuw4ibeQFer8gV+juqQsgx96Mr9DgQENekwFIXL/ByrSm3HbgYE7NojBopxK9
69sMOK4Biz/WJejM5Q49g1tL6MB/OzUhe3T46yKHjugYOT+agaTyr77awNihhzHy1Xwziivzrdww
AONNfi++Bi2nxapst/qL8v3d0xuaEwOT4R7kIbmKJovIv8i8S527BcWJ/JgJnnSlzKZIQHWoGlEt
9W4qJ6K+UEq5MU/okTWa4SEAwhku20rALI5nXjh5P/2Flye1z410tXP2EnZNr2BKItwfBkwBt/rH
uhm3TYAgy0W9cgYZpMqUgGzfoXg2+GSCqwgf134lOMmOvQsfVDyhRPbO75UPbBXABvK8Sg8dEYYh
9IAsR8kaMQIoZuAbtyGK5lUeJEtDEkt1cNp7H5vikNY1PvzOrOl6sAmUwnCZfPhd/rHJVV2v5+2/
IXNCfEn+XV2iqmeX2J4kFt97tQPZF8k2lp2IxrECEnYThvdexYO4Dc7U08RnCWwco8cpPZxbcFlq
qOkUT2ARI7uALTFVT+wq7O0aixwPZk5ANo0lHhFnJcCC3bR2BXHwgxmFZxffYBrUOfK/WY3eNS+Y
+dR7B8d135LBrFpgM3jdsgfsUc1dLi4Auhtj/B/7RTLzPoGZ2lZqK3mzh8zSYlp5NwUwqrqel28E
7KXdzKnGY2Iwhk/8I30auwNWPkbgIqpQeCObrW6Igr2+49/XcXmtwIUmcHmP0WRFMOe5RoaMFBHk
2b/sR8y8mSao30wef9LRUJs33q1/rQJgQTEVpdDyp2ahtHgYhG7f+JAknckhzNXKd5LhGHwLiLoe
SsnZzIV+TSkEeC9a2c+REgGv+d/Ru1C2lOgij4PtEptkmBAWsafR0lHkfX4BaSFssjQp3sDhxmlX
tYeCjtr4QD1Z2MqjQf8SNqCrGF6XRwh8ov398pvNjE8NYd+EUUwahI01od2z2k1mpuC4p0NGJOIo
PdapYUm9CiSTY3IDbetk7cjZiAIofOLZ8A8uPVrql5JwSOctG9UFi98rWhjJEcOox/XQ/gXyc3sG
QgU1J2ui3JN8c6Ruo9fT229PAtPniV5jHcE5OKMis9ZtZJXwP11CGORL4yCE+KE6YrtI7Q+q61FX
v7eABPS+UPzcjJOG9HxAXZWOpjYBaLi7peU99KJUgmglA2XbeQaa5P94TjbHnnGUJVzk62+ylLXc
MTV4zGFkSrXw1KKUe46tXEq+LvZ679xUYcl4W2v7WyrDIkKryiWIkmR6u789hc5GJ0JZZIHgGZTn
RiPlWunzUIYdkwYbRbYNZL++gnEJNiJdsCPTxWOq1JVf+7YBIlxaoAhYnhNAaNJ0irO0jFjpxBxX
Eg8cIK/691Bbp/994DDXgsYZQiWTsRO3YPav5QwORUinuIDdbhF+MQ5jbxof4P0JreNLrgKxd8XR
fDXyxejwlOJUJ2DasD+JiYzKSUeKoGh3WJYUinPvs5OxB7R/KLeWpE7uDYvR00i9miCX9DH26nXe
6vD/cK1lFFJj/CNuDmXBI2XS1Yrfm5qv7+ow0jG++KbSjMzIp5vXtcuy1GFteowx60ZGID8DNEIN
sGj1cLamBH0ZpZRVBDkYbcMRuSbfACzvS7Hko+v4NiQLSWB28odDwEF0ZWbJt0gXonsQhfJ/4HHX
vfqw5dsIw7nOhNDsk43Xwt6CoeVm/IRot6b3+ZFMytvS3F9kCiZcitzuvjzFfdN2lXyypdr/P+m4
oQv9L9TgQcQD4rIzHCua2o50TUILjE6iOkSOHW7Fu565pmB4OUGrtP3pQKbmDiHc0rIeUCA/fdKt
8I4sP7XTdbsVu5TZmVHHH4GBBlI6KTpeiYq1akJlsoGH+caSsIeG1vsmLwpzpC0xBLgzkIg11XRE
LvXiyE1l6+Ww8vMYFJuIChqefEHva1hn+uE/8sbnvDwwn6fOdUdZLf9IA6GBpa1NWy+Vdcv60oyl
brcYMutTfdW5NEAUVZspKPJ28woMSZh6VurLipHnq+hu+VNzmYUfR7dQKC6aYImqME1lM8JvSzKw
bqYNF+REPSC9mhdRy+RF8onVd00QvRin1Nj6Fx8N9btFtyuGb9jHS8+68REQ5S/4XRIufFJ3rzmf
wlDFmD1ruRVbzSZ3koolfnK/GzhMDVbQ2um4gGAo5omBtFvX6pZdhCZPsWWBXVNOpt76Q+aFrW8h
8UxaUlkADjKQvTRHOdZK7cEk+6k9gBMAz1m9qiLk3B+8VGPLvcwjrCtCAF6p4OYjL2fN3bVhhUG4
viBJbs1CUcCxmLzAg0ujLy+dtnlyZdacJ2VgEZiHTGg8a/1TDTPSsRSy+WZXNByfVXsmZ7S7HHhy
GgDBjVsJkWB4+O+pkk/fBJeB1gOf3qzn6EK6L+cEpivFqQimbvMND4TzYRSUyqhhkoFQNmQETIo7
6w5X/QGVkyOrv2v83sO7EKnfljj5/dx2FGYStJfmBiAYwvZTCpFKYTJj922WDwdhXu6WqKGtqdD8
agEx7wBYijvbMQrO+21aRbY1Nb5+hDv/pybQ952TXSOf4dodawTSIm7VpSaeP1It1nqkr81TjYhE
sc9lhx6XL1FhHp3Ski+UQewNMUPbs4H1dpL40NPxcZL+xG9NeKGjeVWVjpCgnHwcBTpD5IyQxeq2
L9SYWBvCTWGlOehoYZlBTNfhHNICy5dK5jKwOW8PHfpLyfgj9J0DlHqT0WADAf5LCmaHeB/CjWyd
Vw8dJhEPNMQqNwz/uct2CuHjqTmcqomes4dnkwpj8YCCWRVnUtza52/T46QXho1Z00UVDpj9/wje
891K2w6wNbZZttUhy8qoBIuVxO90kYdWZayv1kT6+lWR8L5GJCR47LmAUUI1VzOl7P9+4Vhc7Alk
0NNLmiNvkQwkHnBizSXYR0vFuDsdPD4BiS3m9vVlx0QQjoLS2VkjCQaVgqmYnAWCcR0DCi4gAmJ3
/LgyCjxaBuUy4B384QyzJR1wG8bzs9JLmH/Hbl1Wa73ZeDgzBty8yPqq4R042Ni62HqXAbjfSo+B
PqszZCCmqhi0UqgZGMqPpVrYNvDhvLR03hgpVClfinT5XMj7JzDb38xpgD0al5HZ/8dc9JB5tA/d
+Sw0Mp3Vgyya3s1O+qNfH6DpMrqe3jB5yVVRPCCl8U7beQrUjBPeDqAG/JmiXqFtTBVyEGxB7UUx
PUxjitTdFMb6PyHTcblIWQmx43Bu46XDbTbNyCDwTYq7MvoVnEZzmk8oVB1khCWxrQloumjFVv8+
MM76V/qpkzzwI/dWXDqaZIeaIfT3wX0sQjc0QzmCloOXI87qagWTJMsafWR1NYB5XHYYuZwEJBUy
9srYX1YW0GhtI1s2LEyicOIK2Ssqv4ziyeHQ0AItc7ZnxSG4UNmVEgcngao2qnwIUkBTNbAWJe3u
2Zyoc/UO/d73Q4Qc7FlZZlJ80bmVIJ1C6q4faSyUSn8wUFCJiQ0PoVK5KEqI+St1CIjCdmZrDaEB
RfN57FOnUOT7lKoDKVBK/dK9n9cX4T8aIBpm4iM70yAKP5dpfw4eMMFH7ZDayOiHPkAk62mZ2rYu
vKeQ9cyHubP/pgl5Tq9dIfLfVC3Av6TV3GOmSvI2PQr5iQ338xkYAkbxUcHFf00UeTzApoQC3RUO
c97R/YxFgqTXpyTNHNP0KUPBcTgHypdrwN9MUhS0KRzvXQU0SoqSB8TSOrTjWHFb47AlnnVlm8uA
WSzo/9h3nHT4YZD4x5U4VD2H1vHLIhE3jv3Hgoqy794QJoS1AzjPAd7AbFJ5zBfNj2ZCcjRV6OQS
3DsMg+A9+UztX3dOgj9MJbJ5f2mW52402/QeOX4RZPsoTl8sW8U1vkSITpgPbJys3axTcNKkxsh8
q6xgXr71/OjfHgnTAgsepseFHiAifSAdbZOBcBVE85I/fAyGT+00RhDHvs3RGL/72tWQ3KqB4sgC
6Tbouj1zqCYtnZ15xZc0F57EGt4P6U8wvnudpbFt81CJwHp3USw1vH9srMH9XURpBl4daqRZxNwD
luvo4AG5cVQ9zdn7DyINFgrcBOsZJQNOBht7gmTHmRpdSeIKvVkGU3pRvgQVtD/BjhE3TtgA2GrW
+oGGd4IrVOPushKGKYOzCtr6gVBzAlXdu0inCFD4kDx8AsTXx/FbTupA8NMxIiE2tFxFLDe1QylA
+LFY0yYofuAnzr1OD/xEug5ToEBIdICksKZOmnPQ1D2/aaIlqrwmOWXZyO3Bw3MK2q7ErGW1QlAR
N4sx+LL+eQtoq8MIOHVbkr3JLkPHlbpDEmIPeQxHPgCkYOY0fI4YeMAVU4nzBRkx2iW1x20oFugL
vodlrPD0YKdAPM9k1kaydTT1E6JjRa2ALihFVZHVi4I10CryhYJp+ddGzwWaqy5azckkDvDpDlKI
HKHF8nMWBj0KiP9kt1s1DxhJ6zESrjIrKtAmj4VmLO1NE+yuIBCyri00wFxrurq9WH8SE+Loz9kZ
rJPnDgda1Pl/VofHm7yD04okivSBxLzfeQ5jSgNeMvO5qfQ0VuAXQzOhy0VZoqTF5ZLskVrkJQ/M
sgggGoxMCmlimfvUx5/bx6HkPlvqe/EwnFkV52eaSrVu0IcK8vScgEEAku/ALRFvIbWRnmiRb4n9
5WcjoNSJHtC9M3wKyDh7605nMI4zY7CZ+I8kyMGp1/aUSv+Kcfo1S4QbGRpD63osHbyLEduvgWzA
M/OuNTXnmTuJTAm8ODocn2eZkwcIV08qOuQslUfT2xaWWZgRdadLpH+tAEVBjXa2+xBJpc6cfSt6
ygb0TgSrussF0TOUmC+n8DEKZFZp8gQ4e5wzxrObSmL7QTgyG2eiUJfTcKFP622Ew1t1DAEiSpDk
ABSARkNzJJkhFBXjfS7ApTQyO/8Scpmq6Y2Pe/R5VR3mtaUuJ6prqe/YW6D9et/OyGq5laxhl12D
xxOmaM/QAVA6CO44s+bRvQzRv8n3loADMsI2W5BJBcyshax/Z7sSsi0BU5WBSdQxhZvurkJSWjCY
RJJMGc8zvTecbi/qKI/mmVY6gxo7125rKFg68xqdqsndDUOzQVzsalhJvCe5zylG0cDg8jC6iZqA
cvQnRVaKE9dNEBJhta7E3uYVokTtFawVagmCovwShwBpoEGpb0bMBhmklIdQFpRit5MrBuh2emMq
eYpP+k2hSjQuk97RBmR55M2e8UMsnM/fuwz4cOW5qi1bqbwGJYlMuCFjfBBD0dDfGcs84Zz19L1P
+YUgcNxa2+0La5DHcF3Dbcf55PvlAe2C5zzZMUf515V0dIFdKRy+pejw1zylc7gt0jDdK/+R3pLc
mNiuhADldqdM8jJc5sVT752l561N4W8MoqtUyNhUR8uPIxppFE5fo4AqWKHCDqDb0DjvW9HYg1GG
VHjtTGUpMV+t8656CB1WezvcxmBFW+7+N8Dpq4e0GLzDWdUPq4Fn1yHREFTRkEKSfJubfTBbqWuN
tAq6gd1iZ4SADZI+nIUbAKRwBEHy9lmqRVFoXOXoxZO+JL4gjIahkhkddKfNDfcaFZEMMWaS3TeC
qXthrmfqowscd6KNW3MlqTEUcZa7fBdinWIQH5bY+YQwa+DOgMbWNoCL0cIFoR5XkeWIDEQsHGbB
dqLjmD060uG4ncTtMzXUu0xhDQOaEWzhfDlzCpY7sT/eSR+pOgRee5+UPs9e+H8kJqx/Fn6CR6Vp
FpBxJEwk9F6vgceXqs0d29ZBJeDTIkSIO3fX8XGu64jAIXRky8/UtwRb9oKA6ybqRpPI7M7qOho3
vEhvxWDviv2dlvudBTgWVgH2GfYt5Y/IaZVZQkP5Q/WeCkOehiCY37ErlFm3Y4P3lJ7jU1geuMf2
YMoAy25GE9+nJGFSAeyIoNn8v0t7+lAqd+FKJqZ1nBwiN+qX5s/wcGkEz51pSrN2ASmF408tyJJH
BueNs5n4w9O+kap/o5gWCEiv6ylsZlDbJPZugkpscZQrHVHWYR+xy5NbPeeVtrpMOpHWXQmiVUKg
p2DGozn7gieQ1ZZCsH+Ol4S/MXq5mWcyhbp0PVDp00Y6PEIibYI9PttBHqs1z3IrWy+A8P0v5NrU
fmkFktYjwNeAQwF7s4ENocLSFn+ouqEPu2KNwBwgflTbDQgzBZlHMl0bc1L8dABVLXxShjtpzp3S
gVnKBF5wDQ1NZ6emEjY2K+mbC8XIYzEA0Gs9xxzdB3QNmg8LXiKHyVbiHIMbxDvGGAscjYp8suaR
dSirg5QLCDlHXYkqMiAomaOZM5hqYsiraFJO8it6xsHCu9o5NTpxGn6HQANMnDHYFCFTlidWZ/F5
ryuSGLIJEdgiqQRBPhwKQKG77IX/V3vWKgnx/lEjNvh8idHPWTEVzshEb0Ij7tWjwCE50dQun20E
QaluwCxaYtAQyRgvWCK6tuqD2/C74POmrM/fHbLNZFGbjckTyu5AvcNnPpXiuCtVP2cWUZHher1r
6+PoYa3YIuIHl6ybZ9FhYX+x6vhBm3RYaDVUGaaSnxWViM981zF2XNfg0reItadHOMPF/py0Aj2L
W/cI39sGHW0+roH47sOqtGRe38c4tR3z4xPGUB0QyJFp8T6Vx6VegPySkwcmVetWFxBfcDuV1YZd
dGNRAnUOeRs3HMaa+qB4P2ufj08mnhMB1fS4Vz/WFFy4Saw3YSy/yWrQG473HzMCcZIy0jCCXiFe
KbYnsbOojTK/LB4BwfpVmoFEXp9dO30gM479mQAJu6cxL3dpCG7GS++HQth3Q94TVyPiOlUBLoAi
z4PIaikosgagLP+0JNZYP/d50VJngDXCzaiiwsivMXhq6OTftd+J0w0Ji9Id1MN7dfevI1m4cRr/
9m+qxTV0vJeiuJk06RBzsGZBXa+ttH3eREz+h+ufIGwelNuuI+DMf9Qx7hm4ZmOMD1hCzLiGDPXh
EVXl8XLrXZTFqLgrtAIUi9NYxD7zxd8Jv5n0RI29KEkiBIwTWdWHO/Y/ncNkqYy9FzObp6wvjpNR
M2HNFZPfKXCqQkRuveRbfVDaCZh+NA2kK+gNy2KJLeyTtn3jqRWDg9TegMIirInM3TVoGeif0rjI
LKgERUxRBmGAyQmS1n1XRBLOE82BPcoUE8qo7kL4woIOEhzZ5DNTf4WfaK+Tz87YyTQ47MAqqk8t
NCEoAToVUerZKryB2a6Kfcfmgl3GycwDkd8Y+0s673L1AtH9+gxkjPjenZg41zrfvlCr3Ktn3FWj
zs/B3Qqx1dvpm07tjoNVSsHDrKu2+zPIrRXJNjGCFMrTN8AEk2mKvuqekwyIi9Vv+/kz0IpxWYSV
Qcx3OnrFfOLKlJBehiBzsny3YVZcrffvPbmawIHDkBCet6tbfzYpWVMgtpqPy0/0Z8rKBBj0OKLD
+iNX5FYDqtdtoV7/xpMaxBb6EhEeO4Ps40Yier/r2/B96my99qp/Qy6Jh1pBP7Uh6SJ6kmnFYb7q
xJIAKOxS+cupHbxxy947Nj40UVe4JQzUkoUP/E97Xr+k9GJEHXL90hEHDZoNe0IAjZgiEcg8q2or
ySWn883g6DEw2Q+VbRCTyOoz5woJ5Hw520MQnRBWAo3XBxeqqQyx0btVp3bDJOEXGS/rNW9ygttD
mgfAt3s8478xeR5p85JiFhyDIN6DUYhKosTZwAcn8sT43VBCTGj/R1FHuPYUgNqHQa4hUfJhdwLx
KR6OvTI8+pLp+FhgdKcwZL7kf5PhYNt9MVBKQpcka1O0TpWyFG1pTkSsi6JhL/xSRnoW0l2m1bfW
Pq+Ydl2muApPOu2kVj4E4luqNh/d2BSz6SK8eXXrtsZwNzlqfvzA1pKfyjPS/uPyM+WaPCB2SKL8
oqyVfexdRzPk6e0vQcNPslPFlxC0yEb/k7Xy2O3eL+i59VNIHJ+o8d2QZaldHLgIqKlg9QkgVzh3
7CYSFnsK+a2uJ7TndvLrxnUw+HDrm4c1/9EerS6IIb7soWzGPgzN5P/3oKnPPOaRPk8Rq9cpgtVt
SjeggTOTEUjK9kHrkIXKIvsuixSnwZKH1aNjPkZlIFw1BNoE6mLKGuLB0NDohyWNkLdhLdR0bLsC
EPFN8LCxOx15Qvx2u7kzC5AcTY/wBpAKxnmYZcb7admCD+W1bUEohWMFd9nOjuJYQadV2AvfB8nC
+MSGkG0mjnogkXz2KKkZbZPODq2OFZ4m5+EKgpdGEbzcJcD1QWB6y2E/zOqH4JOHlAK6XXZl58R3
Wm5XIFgcOMdzoeoewLA2SyNKJUgN2QI5dSKRAnBixSANPVjlT32XFjbkmSbZvOQnKXDA/9V25MHG
v9RC/Asur4sjQ/0yQSSDWxFcPZGeDtEsK0aOC3YdPc9bT/F7ClDOasu+Zo6ah+W2EOJH0+aoUO1N
uP1hDm+yNM07sAY32s55F7mQJRBi2B/vf1sfW7SK3GEfaFyiXFyfb4TrunGWM9NsTbPI5f/WLIP2
QTrLtZeIjLsriQFxUu8LYnxPo//nFfLiu0vXejquBayFVahv9VULagSlOSG9FMsh4vYjfXfxiYBE
ElzsAP8IXJRyro3Z/hqeWiq7hg5aoKP1n3CjPRpKgiwh9QLLF8vYtFBV6doCTdPXTc+PkILprSFT
mhgKt6ocOdueKdv0McmgAvP26C0aKsoy0GvGsrzQXO0YB5OBbp50xDz2OQGpLzm/oQl7jeTkNh8w
Kh/vOOJlBepBGGlNkNsCeXMoolME1tkdtaUoQuGkXTwln5TjVxmr7sG0d4tsiUbTl8Vfx0nlOc+i
HVW0fNqTaUx3ACpEXFUXJaZVooaZ8bMWG15dPQyIYNddOuHpA3K3M9L7aHGauplal/wqU57knUWd
A9q7ccg6M5YvWSCqr9NO6tezvtZDjCfNW2F7NkSgVf7976MMoW3WzmlgvfKWnaSS7PExKF6BRTYP
JMA+Oz+R9UdIPvv9A6lC17wWlIoIZz3ebhGPJdAOs1oNg7WUoyQk9qnp5VpjkHS9q8pvWttrTwx5
eF2A3/JQXVCm6vQHzzddskskfxIP0/jBbejPWb53DgxowIIqfikrAUWMBNpRNbISuXWveBKevDMD
e/cQib8lfQxpbt0Y5+qTX7oq6ILliAPJMaKzIQvb4hXmHzBLwJoeyBcqM2IjF/KI+2ZrFLMnM+8f
ljZTaB5pxq5uPCBp89pX4HCYWr3f83CBCBFPKKX77ZxDfTq4wvVyMb1Lx7GAqxyjbNuNxHfrv+DM
UssIyKUtKLX9fCyuvitiYQrf6Zkodtjm+YR1ab55iySBFFrcpevp9QXesZmiSHvOsAg24nK0/aB4
+p1W6RIES2/OecTAYUi0gIoIS8R1Tcw3Z6Q9+goyiBByfX2LjAkx89gaO/nX5bcaBOn0Qbh8kxef
1EAHSSjB/TPtnoPpYaib4I/CVJyx6DDkB9dbP2npeyvy9JfOWl7skZmaS0tFBDK9pNMog5MHul0D
GHluyZx75INU4ab9HtdSLVRBKnySmRFHHXruAxBI1S1BnuGxVFVFQw+MGTjscG+xlDer8jFOQ8AI
2iTJGwJlzFKdefFssXtDk7SrGL6uLUR8/UgLr5h0eqZ2OH/k1lwp34m1Y+yywH6CWpWDUBLQsGrT
7qeeM2Basd2KitpCTSeYaPU+n1nKyWkjSvDOyZpolq/4xGCSa2X+bkcd9TcOU0KktEHvWD0ZuRIm
2KkhQ4SXFox0hPTNYKEe4wMY0PUUMGN6KRtp6srQEkt545yQSrsrBofojR/UaoGyLPvkH9rYaURo
QSkDg0aPpWkzX6AFkJVZm8md6cu5BO14dEifY5cY0/iddazUyeZO7SETWa3/mboDmD1pg/pDVchI
gtbdhCQ40pM4IRobT50jPH/CYJXos46uAHdbTrdulDzF+aO+REOPjDDrMYIiyn/yOt/kHyjlmL+p
1vE8NTjGa4MNlfq7DBg5QFkByAH2njDpa/qdw0K3KhJ6MI4usMSHSP/GBSMg6u6oix7KpKndx1bR
UG0Lo9QyNaAif2N1zzpBSw79e5Dg9dU0rqd26Ykowti+BbRVS2m5F2DxGB2yd9TU6DZugUlZ9GP6
oU/Wg5QtGBn9N32fOWM9tIOyNJUc9N+GCJbh6bh2Vts5o9WvYVG1xNxUi/Uo0Nrip1eAa36LEhuZ
R2mkez4kOxjp4K3xSRThxRxo8gjXYdL4J5+RniwPvA5k2nS0Ej/BlnsifsuVpDyv6saWXEnAznJh
MS2EQbCruubH+i/RHAq6KzIlVUIWxM1KHkXUxD2FYLPmVG9t2SggixbubLZdtedbDuL9tAwkQAzC
AdZwQec3NNmma23yOZ9jiKSwEPnzZq8d5w5rds8d8xAyOdiTh5fHWsa69qpTafHbaUJbTDuadBfB
JUOVMaCFOzwtv8nBUMGbUV1/jrF4FrKZQ4HFISEkVhLJeielZr7DVL10KCqZB8h2da2DtLw2Y1aV
sJlLjKk+iRGxBaHiF0YA2pNCUWi8X1vv036IOkflq6ciMRdB85poV1DVbQwbImaYxWt6zP6U8CJ/
cSnhPB7P45KvNRMeFzc4sDkl1pYN4rhWku8ZF/+03UuGP+SnHxjybYzbIekb4mOkCRZM7kgeMDXj
oC5VvWe8sV3E7MO4BkxEAxDCwpJtiNo3qCsBLpuchk46PIxWKDmwvDxPkDbKzhZcHy+sFYI8IXJy
bCSS/B59p4dbtQh56TZTZP2X51Y0qeg4UmXGJWnk9wZsGeIX8+s3Q+xEywfkHZewnKHGXIKS2ta4
VCGrmwzL+7MeCdkJsAyq1ERy/0Y+wSukMKLlE5g/+hSCVtia/1ulxSse01KD+gHoxBsQimcLrmyt
NM4u9loNU27tY/0wJl9/MasgajTMccnR/NjxwAlMD/7GVUmC8ryoCOTVVKbMzPxbveq9IfTD4vn7
/l52TeyG15nyS8K1FflFksW0ZYv+vgwtIWKbE4qT9MJscvNLp+FEzIbn7sSyzH05y/gjZ1zgApgN
mfw6ibVraR4ok/MVoLNPsOnoT1eNrpuHjJqM1iMfX8YMON0Sh5jtoQvDNqf6z6V73ZQkCLAHbcs7
qX1SbAnGUAB6O29eyMHqYrbpnogYqRpx2MMTQ1v+Cxc3OZ3g/E+yxASGsKNcX+JWa4SgenEHqvtB
llzywSVrHHBnx0/VNTNLhh/1usPIY0fL8W1btmO4zWJkPNeEelU3cTuOaKV3qT6ti0P4p3mwtFyN
7KZM2HNCgonk52aYbQxrHLo2EO7dfnx8zrdlXfxsyOMwhFhhOI94cUizgV97dbFLNwrLRkd915fI
Ldk1Etd9MPzkd8Ri7eP/QkkBTY14Zx7fhDs4sklzeAN0fyQamJBSggdlgmDsKpCmKIsgDQdKd4Eq
d3KKLJ/DtD/vmaLLRriVtC1/YE4S/PAVnO01u+9KKnOUEvBFoGd0ea6ENolNyZ7NpaTDa4lUMKMa
XuiXQYdD0kNP45OQ+AK2+cKVcw/82quqatfHb9hKDxwSQ2QXxvF9vHVsbAitgOetaAkN4I/Y8IeA
gAvVn/g3UDaz3NLKVMVxVmJewwQet9UX5fH8iF/g6XUl557fteANk8NXsbUrC0gF62VSGD8edgjH
VUef22jcn6ZNKRm1MP5nJRtURlIr4R/CSKiZD4ss5QUlJg5AdB1dReS1wk5csq1yCmgK72jRnzSR
ik1ugDIM9hmzfiMBHJ+lio9A0Hoi81wINLleojrC48HGlsasxI73EG0jpcHhvtYIcYIVk7aaTjt9
VkCU6cJwVmikVKLBIPbALtvKStCgMyFsL/TWcNH4zkZgIiLuRGGfBSfWwSFdpEyN0F7uRj6CsLNG
oWnQqCiuWg0ASj/QQAkb8W7D3h0gEayMTFcf13UOlZDgh4Nj027WebtUjSPOdx35CR2Kx9naar71
/oaaFGS7nSvQ9pk5KjiSvffiJUiMYWQnSy6U4nnLensl5wndyzc4UnMqFOIKPKTCEz6y2jkzBynM
JpFXsxfyA7+ByQEtiDheYLhLqG1AR1L5vLr5yqwPirTyH57FwOT+gY8w+FAlmxPN6xw46GPEZuCN
9bJdkDvuyJ+Lnw7KPlCRJ0rS5UwAaVC+MlSS+zxILGYduwd1JBfVop8epwY6lN/NjoSGGJ9bcIOm
4RxWEVoM+lPqi72udvFRw7NOwd0ya3KOJgm3UXTVRlQXyKG7s8baeYo4h7GZLMObuxcfQhOzCLHu
4tAVhZco/deZxNa6i/wtB2LCXurRJ10GYv4nfVOzx+Q/8280Fn37LHZZdIMMqXnnQHCDaRToyMuz
k1wb8Hi4nAgVxPqYzsu1/6IkEKcELSx+A60T+++PtoakAX4HJHtdAtuZ+2k4HB/nnWFY3AluFKLK
leHeML+Lcm8Shls34ah5PpJdYwLizgxs0juefZOxUGErfdGxMxsajZ9KinyL63NfuoOmgVuyGi4d
x++lnpAE+rlPigxCMOBy9E+7PC64svyR9J1KFrsyfAHzg6RlSiN5CBhJLfDfzehh5NK8dBSf0xBB
AR6Gfl4AFMV94O5ZxQNyc/9tEmxgAh26z3HkbF4QpDVwawhdVW08EnWv0Zk9GvXd8ldrpCOZZ6ME
Wwk39U/iFLd2nwy1Hwp6+bIFa9+3Ld5x5BjJp0rEUSIPaPsZXvlgDK0cWN13UPD+kQrf6YSDxP9W
o2qHolbJf3wLztme//QbeeGQs+a5bwbMswv7H2DERTAWfsuBWFHGN67+SqY2CcJ1Rok02zA/NuQN
bp1vsmHQhGdS23Dj8UsfK5phnjUCSoI6m6WSb1d1HFY1Txxt1uiD+gSQxY806BzWPrXiEcjIONvV
esgQXf7Mfjb0yTZitFpsVbMRTw57DP/zmeEyGgb3RfdyJLRdhETxVNyD2EYhR28cE50TSJ8SNp2l
Gkj/HEGIMHnoV68KTW6qsRA6LtHjApn580eWrjqCrymU5e8JJ5z4CMh2T3IR7zXOEXysAd4EPrnA
FRooza8X5JM2pzDZHD4nvVVKzn6zeLSv21DUoWVnFyP+Xvib3IpY/Rx+pr7LfgqBRJlk2UInMxiO
LRxX84FlIOoHvEzamQhWPSPCQGLvY9AOYZshbthTS2qDOfjCIvNRjdj5Fn3TLqmY3v5JB0XJ24/O
lDUh2uuEPZ5o1kIi/Zp1EDsvU1A58p5Q9D693wc157yj85hDmmWXgTPgKfY3J6YJCPzncRJe8916
Usuz7V1hir1Ij4VQ3k+ws7Gvps5uMXpziLqj61ARj+nJACv1NrGo9fRArvq+ecZja3mB/UHm89vo
8ra/sgNXZvat0tF7f4QfYzn2iPaWyp9f8enmYG4H02XN3ILDHtJUAeBI8yTwt/kofnytHcKBIOxO
Jszzc94XM17rjyYvGJQr/Nlvxzz1RIwnwd7UgNhLXLT5uzPJHDekioBtCxRyNma2qwOD/El7jqUz
Vqze70YCmnl09A8wxfn/c17ycVG5iDrmSKK3u2Mrn3JUG9KEKMwzMvRuDJorhaGSDse+zBHAitxR
3HyoP76NNG6SbzI5hXDwW4hJKBp8DrOQsfpLj5SSBYHaOq28DWHj050lwkCpqa/c5DMM6ET9Fn8x
5to7cXnPsddhpLYIL10WEwbGiIPRmafzVovNh9ERLuDCEtYdzZbQYa0KcaOuUDfb9DSoR8cioJNm
deFkRWlXCGaumvtBxtR85px++rNd873ET2dOos22nq43a4PkJsR0s+cE1XSHBaXwrPhac3sTW/Om
x6+h3np0aTqD8GIymYiiPF0h3a8Mv6aywWO+U78rAzTD/JENZns0uS7ypQaJ1nK9cWDJ1vrK9G2N
RG+3xa+aG8cM+pjPSzJBCJhffzyOn2CP7TmXfirLo0XOXy3cITqjGliTMDeTYUJFsksBfoj4AWoY
vK6fR6ICecb/TSNFRGr55edjDrxUT/sYQUq+sW40v34p4DuXukpEFbXAshJPVDWTi6KYvejPuBuL
5W+PWX88AoQ4TWtkUjtrJfwv7HD41VWyN20DJmW+lfzJlx5+4ZMBJymecb0zCqVTMgfMRzmaGLA/
+GVnQAE4DrMCFnQGbF9y5Y2mwTI2bGnnXrfvPVMlQKdFNwy/htBgW0uDWdBrQ1m2zz4uuhb8UsS3
E4FiaFZzEttnoTGP70f3G/a219uMfsWuhaNwJkrnm/7I8FJTSw0BKsKeMq3n5H/6k3riXU8Ak10K
TmIWHMpLiJMjnZDBHxcbccjw9vs1CU8dx9dGqgf2b9mtU0He4e23UL8YK3gNCEQCRHqd0hxUu/oO
NIInqn5exFjVUQPx+Ahk6IeIKESDVwikWmI6J0FeSwpiAOUsxsRa97iK/s6rOLas9DBdtH9ap6Bz
BZ6w2f8aTilqshq2vN3g/5rivMl1vSYrm301WIwSHTSLYrN4RUYq9yxpr421IkGUemvcpLwvkDSp
G/phuruj6sMXwnUR5RSAL0aZ3axBYl619xVHnRK3fTP/HlR05PZD08JFnqE7dqnmtwe5VX22g2ge
CS6K9f0j7v5n4b8Z6Vd7flE1LwfDrAocPNhnpvhQ02aMRu8jFgNg9i+UIQdC2q0d+E5x+imHDAke
mlauTuU7Rhs6Cg14FOCThdCBbyiLm68+mr3tdFec53W/bltCIA/581mElZVyKC95bScss4UF2+fH
OLl39qrvNscCGUfh/ymRWAJr4c9v5OGgPjBVxlKsFgvsGCMWC0Btfcq/YJVGo1FlbwEb1wMMDBAA
62vEdkDvbd1rMSk1vZQtMhD56omHYf5NNPyW4Cgsi+4PECfRPVo0TOzdWnbNlT1vTyaklyaf8U5H
mkt2CPcjHkxltfHGqT+77Qp1JfZe1GU0o5bAY2WCiExeK7ahxVJppNt7yq75UWWXRU6xe84ullj3
KfcDDyP+jUJvGln/gwNv2oWNTvy7Yfk7EIZw95Y1iXWujmhH7m/eGoNqIXsLkDsFQhy2jZrzvTKw
cg2iYgeKvlTBTqZgJ7M/n6kl3408hs7Y6zUgC3KKLv1SOljzWU+X8we5XRso+O+SB7vyu6xZmTvf
AYHt+heawnF9TJQ2BCUth6H9GOQv3pzphPBlpkUR6gX8G6SN/m7RErNokyoffeOsmPKyySO50sFI
xWP1JIKGqLkCjjuAfiuIWepgI0v0tBOpBqvGO+4ov2xWHu2vsPZTsJEsVuCmKv8+P46Rll2YVzxl
gCUSnAxUWEv0ij9zqyTRSgWP/TzTrYMicgTCezv/Z+QrzuxFupp++dVIZsoAJEZSoBkW4Gr8mqql
mTV4wRhz4AG8E4nAPARU8MCesNCYiE9O70xlvi4JKrCkmgVmHYqeGBXrr5PuBH+sWv4FM7K5mtWY
UbqWaPGyWub10COP0DPCcuLrjGS0ye9hOIHLoJKsBLLT0aLHVO6bH3lu2hZizUEpvHkTC9ZraTDu
f3nHczraK9Y88it62PrOPykkidw5Lczpd68gI7/qLOoiMPn02Y1LoCMjxSWDPd1mN0FTZXv7CthF
oQAN1CxA2urHKb4htWsGyo/FGbDWLzFKssznNw3fJcyZPoUqa1SWQd5DNJopSblIYofdz34SQBtJ
Y5JCCtpABQH4JNdTJEWSa48JywHc4b5mz8l2iOqLVCWruEvLrnrlLCWG184AEaK/c7UcgyQ74c/q
ad+Lz6J7aMkkxkzjd5NrwdV3L0GgKI913Kn/5Di6vGLAbLqV7UzTnZbCzkfpKVWtZg2ogQyEX8Bh
jSwQb/hyWiAdEA2ZsgxoXFzD6k84RDMI7SYS2o88HGBqgw1pBUBGE/CMHG9prl/cKdx+R8g87vWl
sD/sO0A6JFK/ZvhSiDIKu6ZnZHajT4/f3wzAECDvuX8h9uvIf7bbxIFQ7gqliIHTu1IKozwDQ0mg
pqtuHLjWylpFECAr+Hl5to5yDB4KimT24ke2/Qt/aDHYmSphUp3qq1bl7GSD8u790qGjd57f9klh
4VEqwhj2Drkij5izbmx9Oh2RgpdJFYjfPqrT6CnB4HIW6Q845Ebgxp8l2BTJLiSWgEWvzLQ+QXSo
FN9wMclwIxfgQ1UCMLZfoCozuhJnTqd/M1xEfksy+P72Qcq/vnZdVat/V/+Qev6kt9YhpomfhnJn
bQSAudl4Cu5QRdFpW/p/fRvq7M84/34mS4Bxn3B03CVjZamFB/HrZ6Bl6Ma2k1TV/DxlXPFw318O
66s0MgsBAQZY0a/mezrTPU+vKHlgTR8w2QP7dLrzfGFWj54smdVWwcB9+OAfqBeA05/2OsVE5ZiC
FIWt4lA/KRyuOybTMBrHOcAuptWoQEGzfxvu0NQRovTuP9y1djn6ai4wpigqpfhcGADodrF7jnvB
mjLGerK5XDVKKtJtKndq1iEzQU6BGWBhQiN30MkaNqucF/XJ3E/aEK80Z3KBigs5+RDL/N0OnueV
HM1mOzbRMac2oBmYlSyHDCnGbXKqDwoB7G8NpFV0yDqUHwq0xl5nBO94/av6gx70SsYd1D6IRBnZ
2y0KiQvX7JngTTMyENN0AkVsryAmS+ohi0HPd1JUzjagWhfEeYhWBW/rAejmxblKyN9sx/onXkiA
0xiCF94Kp1cjx6gfmNT/T57L/XruDq52hM1tqFAt5Y5XO7+1RouKsTiPtGBMua/JIBgRzCM6I5mZ
FkPSiGYvfsloWPGznqJR7zWBNGNsZzJl1HRYKEjZ3BbKwutKJKvOX+VbwEVwhJqEZkp7Mk4XiNch
VHO0ncVQcWFoeTuDIQ6Kg9AHoyDfJxoohMUYtH9Va1ZyM8Ozazkp3FNnw9G21zesF4rKuPRA0CHD
fgDKclFr8sZhC2nj6HCLxO/zI3lPY1Nmz89l5hpucwzHjyfVhO+DSzKvrFrqr7GuzFdOhU88Yefr
/VLyKSmBLJgNd6JBf8lQAvjc+ZUYzl4pPZ54VxwwraTB3tmcAwG7FHC7Y6tZt8SsYxm03f4Kpf4W
920rKiCHfi0iBP/DyB9COY6hQy+3nWYGKAtt36e/2CZaulwzrMT+9TCW3VZY8ek98TYu3vEqPLAF
ociHuPCKmXzRozPy81MPO/NmKi5ooU4mmsMHxOtWc9IwZ++cC2Rfh3jBQ4QWAvRV4ra2FJAirXFk
sRCjzoubs/UZJbphT7DiMF9XTiLFBP8KnggjEcMd3iANHFXT8o35ABBUUGdpPes34TcSMpuF2VmR
NyfS8RLnp9ZTjeEurYQh3KNt6Wjc8HaX/1T0MToPe8UjVze7PZtLeBnebkYAMWoupTfqq+DipJHc
K7ywC6oOK2caX30QFCc2M3JlmGJZOr/6K0Gz+EcJ8t/0th3pNJJrCREVn+3if7tqdd5UqAPNFANM
1eUiux/mWagZsKr1NHwii6kcod4vlgfinNkhR0VXmfbgcFrUdgWUZaDXs8DzLmWgWHl6uMIkoDrc
046rs0/Eqac9kvHc2NIo8FFmjb1M1HldkFu27EAdAtbCwJBmysjuyT5J1/VZTv0M2Vwql8z3AwKU
EVnFntIp0IeU9di1oo/RY3U7XfkuQHFabfmQz54dg5dZ0Z+yNAUwF0iNqLQP/GG7HbUSN5Ji03LT
ht8ahhK90J/j053M/Ow+1z2X2D1tjENFW8D1uWHDiOb+9Kp0+Rwm0oLFtj6PuGakptnEbB9ZCP4Q
ozhEzyM9tUnPfi+dTAoMtX+o9CS+Rli0QAmQpivr8YZY+w8iOknM/fss5JR5uB+if/CgCbN9lJQj
wY3JDjw6+jV5roRtyiG8gOvBGVUFt+yI4zyNQE7/jBZC/gpDRDaKy7A1GXwUynBYTu9g1Z6IhKRP
woRGivrWC9wHmahVLEgayaZhV+SJg20T0na/azxwHDgtnjym8H/bhQ4SMaO5OqjzVyZxBJgXUI7x
1Ezyju90rISLiYPS8ZtpzIdn/WIjIE9IMGP2WxDMCMcKz4RqROdUXn63xw9o+gShXjKyW1J8kVsr
nYQM2Y2dLmm9g39R5aFZMHSbFHJQ8bxMtnEERbKsqzR8gIm86PAhrJRomQGrTGTrZZI4ZeOf/yHA
szRamWqnQsQWrYOEv49BzS9TGLmNoFAGKg9gpYHAmR7Afu0z+DsnUC5B4JyG2Gx/IAJC7Pp1+aay
HpilqnBeZGCMETdId9rCeo1NKbt6clUs4BMsM0evs4BS44WoUvXl8xwCY27+IuwhOXbrlLGmw9l4
mBX5Mj1gF4VOcdwipy843QSsb8O+X+cfAdpwMma4R4jWDGmzpvLVkkObY5oaDAf/V3XqcZIz+Vs2
8WHIcmwPwTdDvb36WlhAbwgkYlZtP/0eiMcG6Jxj70zMTgboNGwC0bh/zL0fDMZIdIYuKAXUwbdx
6eOnykIhdpHMhcJn53wBqwrhQKiYOY7eUrSgPd33URD/Y7yWPGgGlg7JLiUnyFt9A63gYkdnylRC
Er7iFHs/h5LHDpPlqwk6OAMZBM0wxjXaRKjEf5/XKbV9a1G9v1XYgym3G02Nna57JG6c/aW7TfYK
dHwWH27tO3RBjDv4uwH39SrMZY9PstERmwvNQILiUXDduokJjLVbT/yj5o6IB4Ei0tJzzbSFrbXX
94WL+XvoqECSJ61itQYy5Vrel5EAYIWR4tgXjGGOgbNOcePCfMkGjm9plpM7VsPUXbNon9qn25FZ
3QApmryhmvb+t4I1kZRP+Pl10jrdrD6DnuucLgJVfBHxtEGNknDguckDTt6f5aTh7bXreGFKmb8h
jIf+DEFeZlvjDCjVWgwHUmEPvc837vl7vCyCRqbGmvQBnvyiyybS7F7Wm+uzB2iTphtwKi6OZ+ZO
bvHnigmIKyab2bg7I//i16kCxSax499CCl8DbnBYy54TI0WLQJIpF8g1+7N6/nv5UKB9mhHsNYaV
20jkm5aN3+j8imMaoWstwcNQQIfE6+hMYFSeVBBpmwyYrcus+dk3E5tjtxkBfxjAg5Tf5OJqNyEs
OmsWxhnbvjZQheBTbaQm58P10pQc6bj+ICMy4Yo/2+FTauzuK9pckWc7mfq6Jd8p4o4kAO/+fquC
EBeb7vd+ele9iyMtsuC1WJRB6nVTMiwmdB8QAAQZCwnXDU0DQApU50feGtYNV22RIYCsTGsm7A25
bTXkug6w5idTuq1IU4zXUszKY95b1onOQAi+xINnYrxo48hjagwC1ILpYeqfY13uIH7k5qakCFcC
Dd/x7eRKnvMLDJqMRhran4B2ObOjUDmN+NWyBkshexf2hRur6ZQuip6q6QBlLCIVFTV/NAwL2lCt
3YlOrU5sHnUX5RYiwolXco80j1O+z+au+CNuDljIeoi/hr7Ae++oaHeDlkO3MPSvC+MPcdfbMdBh
fUB+2y39+RFbFynMAq7xJ3kFWLVfHQiTOe/EL5rk/CyNBJ9zxN7UIWxMckGL94S5sZAXZT6bvAg/
PIlKxmnMhbb2+dHFGacEwE0/Kpa/786GCFt6sgYm1kwR5yJbLwhxvvED2k05pIscJSbvj+l/C1uj
5wc2FthPqFeDQU8gKF6vLBAE+ISY3JXAmQBRT11FHoCV2twHSqI2fUZbWrF5nidftgqEKq6f8741
Kat5tPUW+KW7Rt4v7mLq3hcUhlB1bdxKrcolQH5UtGN8X6Ev2NUFdiwBIEIv3kwsuAlFD7pWUPS/
ykQJ0mGE9SGjO9YOaE+rAwTV+d2sh++rwBZ6PPd07drbr/3XOk4A8007dLV51K1gQooBlisNum+f
Rx2SLFxuY+PXQzvkOwW6uaFxmd4OAER1Jm6EDGcNuDpww1yD6i7gsANJa/8agTiVXmE+n/H/gLqN
pRb9jkPE6XmoJQdHbjxaA+Vh4nDDRMpe2fiTQ7na6wH9IqQ+x4o/3pcsLHH/d3m6DO0P9JZmM+H9
/hiEsJk4eUHIoRt+VJkxn0yH4y+EnSZN7f8Jv/QdNOxlcp6dbRMjnHv0VaHEaxnEDF6T43SJhuLP
EzXdOz8kcFscrRK6iwJJwVpcl3e6/O8k5rIWse6KPfD4Dy9OEaylorr4rHsrOPCO/IjvCbgzsrB5
9vkwBb/FUimJsN1a4By57Fl7WF3FNLDQDIeHpNVLzC3yPtLcyHnuPjvBmFd5ILPXHa75FT/yH2OJ
nsjj/nIpYTWb5CMpC7q+9l7uF4FZuGssw0sK2f0LphwU1gt3Tw7Egr8Qcwy0ko8vQ+pSNcwnx8Iv
dNZteT0KZRnoeLnresRhL8I9nDRlyWtCx+B7tiObR/8y4+J7LKu1C9AFEsAFll3VBMSTeiw86lRG
nokikchAi9GHYcFRJhdigYPerQHoRSCMcNzuQFnA9FeC7FYKM9GibS4wyrLTQP4WiX2v9zdSsoTz
5FKssrOKRZ9cc8j9d6x4g1xlofeDf7R+bJ27WUZ5VX+kIx7GOdwkc28uARp8vdGxRkFQyXkUFeq6
Kv56Iy1ob+l0sH/Va+mUoV4M7n3+F+F1tv1FQK8y8pug06IYKOrx2sNbn24qbDWoQBCiQyGxbutL
XQbnLtWF7iD2ErunTlzpyt0LZq3HtOv6/BBO1D11ZG22wi2Q0zgpdJZejD/BcF7p+k+e7iOZDr0T
Vum3wM+0cyHJn7kzai8HBUjLwXIm9kfgLpIoszyZXrwvAM9FBfqOtecZa11VtTzZ9NZEVmD7Vcfk
v2K+7Al3IPIZHLGluZ6hUM0sxMdN27cp/DK7F545wySl6WZ8nsNymHAGVZavFjJIpCkfeU756zYv
FUiSXZ2CNqkbEgidhVJAZZvWCfpcn+fhI6bWhJcHa2jjjSmQ9bE2UDoXEaa7HGOMdQ8cjcPhM2zr
CnNUhk5hpYk8KSZzwW4SiUTZsSiR3jw3mW52RJlopaQWachKKI2Q/PgPyrxn9L6ThMuKP5FKeJZV
wWF41o148ZW580Lb8zjjlkXWEJ7gulJed/jHG+8+NEEBtoG/bJT4PO97/TYtdgh+qCHO4yVoT8Y1
n/5Lg/TPmeRRVJ4fWDh0Fcr3nJS6HFZlXRWJLa4aJLjLHiNULQOqGf9bd7cjxi8xP6yBsDXc4Zpw
sd/yRM3K4tNz8rTOnoWNwOtzyLcgile4ACIocTDc9tcV/ZAHQWiS33fGQWNfB9+QkMlEUAHqeTsv
Yu1yO+x84GNJYDw57W589nybEjjRxlCZaiZxWYT9OY/T+YC2OYDu4ZmiJVgGia1Xre52Z0GdBl5t
4NMToXHQdY1pyQYmYL6U55CcPFjiFdVEfPBdam0Sm+1p81wK7MbOSagJALhdmlO/7ASIEQJLcVgj
TKCAHcI3AurNyc9FvMwrRw4L6KxZ2pHjFTGWO6fbrY3LU35b9Rf7OfmvOlxwYKsTKu1/OX8rX/0G
9WpSjuHmjlg7cjf84HbZxNGN8dzkMzOKetOH+KWf4flyRTwibxSk32Re6FNCaD5M+4G0I55QMdWF
jGcgqJtSUbYLMK7jdnAr9vG115LfSYlHl4L0keurSWEmrjYbAXAIQLgcVHxYm+3jvWhGVOJqIPWG
r24wkPe7KwTl9Qwv1k+eFiIg6Fu/Ih2EA3NwXjgkjuh7DmFIU1g5RN7IuoFdvdRYoAv97RU5N/O4
yBECaf2QZE8t29aWy53vsm6HPoevXQN2u3todwLc2BAOycZyYLxoI/tlvaAoPNeOo9UnWfapLdOW
C/EbpWCO+yHx0hzBLNsjBPlAG6MAm3uO6ckasjS4HSOlJRanmdCJQ841lgvc26BD/QkfGoPy8UJg
FK/osCvvOb2jzJzdkLlvLhSJg8FgUkC2SK4B/szqkb2PuHHE7MJz1BxVpecxDB0xMO2zddy9ivDz
OXaMMA4gn0X6khv/I18ZgoAWv7kAbwA4hAfIDXGBzmIfDgBDCeb43FQLfyZllt/g32yBN/uM8LNi
KLaX+KWoN7oR60AqBkt182Z74wtGU0Q7txx1ZELL58ID30bDu+zcYRC4/t0k7DPsuO+6Xf+y6gCQ
fA/1Orx4H+EzOguAIL+B8eAh/6P6qYk65OayZeDSaiZHBTJMDeGt7gHhZ3XBIIslA+Ef3sdchZcM
SP2gljAkow6JbF6C7kUNGl6DSG9ZMmGNQ+e6+ysqZq14WiU74k2FlhpZXbmGe3TgePinKdfbxRJB
pKrUWxMusv5SxP6sF81z5NNjOYULB42aqokaRulvd3Xye3VU2aw6f+igmyn3JA8u5iaA9nhgTHGo
DWxF1HIfMDAYyIqWCRPBFlXdf+V9VsCtSdhlVE2vcVVTRIXGP6tatqWDXdECR4A+qFXvzs9OfAHX
imcE+XAFGVh6Tm4Y9iLByaG0BDasyWbxl5/ZSTUKglswn5mpSM7ztU7td+st5OYSh4AjBORs2tlu
ot45Eg+NGKNfTXZojLapkai2AKleT9s82ok/kpWUpUt/fDgDhtk698/DRA0NMSpWZuUi8tIRKXhO
7fwINWttF0uhbeasGTFEgkftDdVR6kmSo7hOCAFT4JrzZfp9F0kUZc+zCyKoE4ISy25gtAxp3Wul
E0fgY0RIM7nqy8tWQjrue+GlvVQ4CpWETK+Jc6fZwC1p0Gnl3ZXoumKO8/r4tEOpx4MmRZWNY85d
5kH8DXa4YDM1ymHjPbYRf/ujGE/35TmD3riu8GZ3ZqFUa9l/TgMHbglpxKVEGzolMhdqkcOfO4k3
qCW3zC8QtydRh1ahjDstJfZBRlBUbKjnKjO2LLghfWQdXkW+k8+DSiKZS0l33QTr5dyL/GL7a075
1Y3XFwfj9CV8DnCqYJ3SdpwYQFl3DFTR3SDkzJkYidyNx/KD3pCKVdBailR37Ta3M1ZXsMSyA19u
RvB2AJj0wHrIXeEOWJibqAbRtJhNMT+cuGIWc9vjfDEg5/Tmk2zMLvX6n1xFj+dWOYmuS49jPY0G
SElysDpLoJt/JqgM1S2ZzorTSvyj+9K8FeN4gI8YSj2bnLFTsAT0oYdtYxjisFpRkff3NvE+fXLp
dqMh+TsK0rgID/TSlpcicUbgyfmdKctdtranBoxqv7uBnE7lS+46t6zHKG5tCoeabjOYNklDYkVm
i+I3s9qgczcSgAF5pI14d05V0pxI1Eye+254zaaKMD/QXnasVQsBQVA80g9phyuv4frhunfQqygi
DHW75YOK6qh+3MeifNXFhunOJJEDgffQ2P+SCfbO8EIy2rWgmYpci3c3MdARdwDqYRUsxnzDG6UT
KwzWZZ3bmAxmNoJ8kMXsjVwmWGgRntwO3z2EPzxi0y+ddTXeVSaxPZMKO7Q1MAdk30FFCvUoyYiz
VByDo25f1EDq48rKCEry75LfTCWdHbhzrA9Y77BYgtjxIsWIZ9NKkoDTPP4WtzTKUgoN0qliqP7B
ZCyVXP1tOJlTOb2kq41bkicsO/UlzTLPQhuqBmcvTZxtpkXxZcyEkzusMiFXfKVig6ZGIVRWjfc4
N+x4+ZiojGbbeEYR521FKhlcpngbGsXqMyrbEXxqc+69RYcD6RwWMCgg/yDL4mfrsI3GEp/quwcD
BDlo/2uDDGn/KHx1cglWJ5ZEtQemP5WkUNwqnOp29DAxC9jRg+nW5m2p2fmUzwQBUJ+FObfy7eDP
WKClSNxdxnso8hbIURmbnCA4UJRl5W088E5He1aqjAEUc1wKHoJDR37GHjlLi9Y3UNI1qvH+AlHf
gKz0CX29J3IX+NmchGq96CKwMpaJfco3U3PL+FyWxM5R3dMSr/cW9n7cM+Xpx01HU3tVyS9wNDCG
JQ/SZlQ6GVkSlvl6xgfVKZKoUq+VKDzL7zCT304vV4Vh8mu8RAQfEKpYYMQCHIxw6ObEGiaPbIKG
zNOGZB6brYIr63WEw7vbNeLZiVTwN4kqPexSUJtgKZz0Aqn97rIgh8QFNzM8yhY8QhZNyMRxcWtM
4WpVXvGfd6SOpBd6kfaoBUPZMU4KrwyTZ4cPdcxR56M9I2zl9AEwWpB0HifclAtFLs9JPB1zNgpF
iMvLOetxyMtGW1BT0iPF5lNFNo8cT1hqxuGiNsGyTYbTRrxPRk+YaiqpkaukBmtw0qeoCkSmURTc
+IFNeCCYXjnR+3Lcbpx/OFm/EAza5Hsno9KjqRNDPvBPj/tUovP/cCy2JroQkLYSLmlsVbXQmMri
aJbKWTLe86PiYSIYQXLuM8sKwFCtX1ePa2Cvwfpd5DJVmHEs0Xed0kNCmTxp45eBt1JfzV9JIhJK
wRJSIMS1JrfM73Xt/AGv2y9bu6Hsnia5BysxtWMEJgPZIBQpsgVemxvaC0QTpskKU01X331L1UO/
nR9Iug9yq+KSgQSliIQbhua+B06f8MWBgt0jW1ZQVgomXQrZkDNc4yYStEHucj2zUbLb/bfYdj1l
ovWIrx7hWHYcZjiM4tPc2JLw1p+V1PcFVySKa7UGEa5ISWmvjyxwpkaq8hxDyyEfpaGpH7mE8GYd
pCRC7aVXOii4Hkz4bR77+Js/kfb7QQP1JXf6UgLKbt0z7LrL7ZGS6ZOAAG3llBBUZ7238KJNIp9E
synlgNlbXrnWIv+gQUPesAFvpTtEp7q1RvrcqIcs0cwAeZ3ZV3SHd1BQqc2X0k6xYkUp7frqjPcC
7z6knsXnd0s5w/+tAV4W0Qy/zTouUjJhavz0EIGtNUNJHsY9nkBXyt6D0hhT6ylt6MD9XSjvz/sn
R0FPEbkTw08IppFlP264HmEgT5zKGz+ClCqQ70yOxknMuKx+6ik5leHgJxy8HFOlzTqMB64YAuCH
713CO16J7znhy5Sr/tbZMs0CwRsEX/AJH0AfSv6lt5dzhHYOGZmaccLbVao5WrzlF47wugHCrJnF
N88vEaZtppPVjWU3M9VIvNBXJRjHU5+qAaudnu29+QX8+foz7XaXJLF3IUIuvR/QL0k0ggmP0iNT
f90Peip5HVW7zn85+QUumAE4nu48VnLVtDnY5ZJzgS17HQSDbR6BYiIvl8bsCoorCaTl89dJXfgo
3VnRqp5fiRqsOzoX0odXAwtexKKGH+nPU9i+mYZHXLal8quK/VtVw5pgIvFnojVn4KhHFacWWgQS
KrzD/QPBxkk2eKU3PJAPQL1fVL1L6MAdzww5RF2CNeS0pBvK4s91wXbJ8/W9mOujvgAnwcIE4qfW
CYZ39eluNDhV6RWkjnKBcAnI1ib4tatgotDmhv40R0feFkuI2exBTNTKP10NT4fKHqZs1ADWf00K
Lx+7wK2MfPjA2/qIw87W/vgDr2zui4L+xf1TI77csqlb9HJaHlSxCq85fQgDugySzaw0rSLzmlkA
855YZypE/LWJfTzyHILTcuv56HbrX0Uw35Xj+uh4SitJdaUQJRVM0zTgTVdDef9pjK5j2CIoijn/
qpsid+HBrcKEXuuCNCX4/U2RI2D7eAmc/J1ay61q5fDvEt/toQOfNElj5b+VuXtpVCr8GDzPH+7B
XkIDPT4+vQD5CZP8cTxZUWH7gMY3fwtOx38Weu1d464cPPfdhMXqYjAXH5wYRifePgc6mmaFUDG/
iaf3Et+Wxrr+9/zTX4VOgPQ1tQKVN6mwZ/FUHva+9+H/yaSbKkiIroDrpQZa34mLBQcAy4a6KPSb
vifPRgWtYKZP5P3tKDf3CmvkazkvMQPzHsU4cOGL24+mcpO73plkqH6QIwEsBIpc7EE+ZCwYt6Me
cJyFqVWsev3xCRni2Db0A7Oet4XalCHrXmuhRqvphtk2CBXmSfoPpaMNBiRQj/u3RLi8McFbQQqC
tVSitEfCOuyFGLcsJ4TGYtqkoYgvUrNaI31oflojBfhmyo5r6EB+JKF1ZWRUiPeVSQH/YfFuORpH
o5ZcKrSvVxlNm3o46sCW2qbS/zO3vxE1F9Rd4+wblVxP0thNBir6ZTGJsXQpgD5XRZqCDbyBbkqX
QbBqOS6lRTDawcijDo98qfqIvCEXyQEdHoi0QffVF04VWp1I2AbrE2swStalerW8rV4RjDj6tBh0
I0LD+kplki+f5aUABPHHEh0S002WO9i645wHycbgFfCEjLap4lbEdqySouMpAqwbHBFpSMuh3pVP
NaXXez2djoGe1mfxUzxGa9H8kZ6tO88bH4VoZEaLcHqQxhkwShmyxVV5UJHHIffRqPpIP+xVRIXW
QCESnObqIypFg+nDUwfrUGhyVSo9+wMnGaa3qfOG72Sl8D0DbOjz0mgOJBBzjJByDvGlO2zOZpVi
+eZlw+Oixc32AYA9v2Vfoifn+ZIHCyaSiqHtvnjFbiAXAviXYwUdZ60vFfLaVSpA+Hrodaj/xKLD
DLwhDo4kiab4uCmSaCiF5urRSN2rguL6egXaNneTFfmisbOe/3RTYcH69aPKvoh0MyODkAOq68Yr
+qRt3PpGYfths6fZ9a1OihXmguUWY9rsSXW2glpXcvYnu5U6BezQ3oRBMSQDQLdPXHMaLhUPA+vN
zIB6/b9s0pwOwQAT7+HHD360/RKQo+60AjWp2mAB9UNrTyT9665qNYF8JHE/h6Yd4I5zcFC9zQTE
AhspzPs3GGZElgGRrPjgATKt2BzfHxk4swVzQeEA6dzhPFIPPB8au4VZOibp1ftgXsHSrWf/H8Iw
zvPjbBHurk0fD0oxUvtr6ZkOtEXgq8tIBjPa89XdWO5oWRi8nClGX7XxxvAvdBNezF11HrLC1H7H
pBHn5Y+aClyXj9Eu4sviWBWVY4El0fallx1KmHOoWgFMPe0g24I9aQIerMN2n9cf7CTCV1UybTJ6
W25JpYiIWaKMRiwuIKCTZqayAdAm8YTWxyOe3/PdWIp0i9SDUwxTSV3gm1Lt/wDw0dHt9A51UDYl
MYxut5+GXJo2mLV8a8Nc0yxsUNoaDXjzNL6R5OYBhkEWUAaGuY76log0mt6YIXnlijMvPA/ug6lp
4xzfu1hxr6uodvCzSrkp2PAOclCq9Xtruj/itcHnMyA83PtuO/jS+CAOOocfZlYCoqnjbuEkXLuL
Az5fd9wSVX0OS73MZ69tdjaPMGWPFSuPCeNRRkdNbx0qaWvQAUACGLOIu6qOXFXRPNBochobMTNB
yL1FqYNJQOzSTnU6hvgGxiC7KBYrX2TMzw9rtmR2t92mMUW/uyrW16A9GqBDp5wTc8hYrLWfL8KG
fTYX8C/VZlg4eDQHQ/qi4qvcVDFqOXo/t4aMqLK5+0rCrUs561qntU8tF+DKQQXVjHr/VTwkG8ru
Ws8zPzBw2zmQhQJil9Y3ClNIdWsWCDj5po9E+wbbkhJePVMiVnzdKZ38Zl2SizGn2f9tpA0V38NF
YV9UR0gvKwlhKXwJjcST09t1Qp+tQQUwaGcmPQByKF6wlBpBJ2N0nYv5diO4u/ZBfLUI6GT29JJ2
OefWEmkQ6VQbqOgDaC3gU0Qmna6l9uMlArqaOQZ6xyk6iuHckzPor5KTKLyHgwzNe2WvLitbYVQu
AS1FyxgHYW38Q47F5VhTKAObEqIigzD5yfWteoqW5aYXfi7/+LCatsDISvszrbJNhztKAeUmLN5J
fp9NhFZ0OQ5Jl0eU8XyVBdbs3iahyf2L6/RXL/cmu0qhU+3RUXtFzqA4JtL1ANJt2RRqCr/Zziu1
2OfxfURDcP6LHb0paxEXND0Ag2oIRhQixJjl7DyRaPBPM906M9meB1awNyu2pabblDu8h0eUvSWE
Krk7QF6rQJLowjEQBszRhjHDGRFYW7IIR9Rk76fKlgNJhRaM4KqiIYa2nQw07RHtRoJtzb4fpbl7
KMXAVP80Bjfj/WaMbbQ8eqa0nWl3HaVFCiSeIsiHSyKxU5OJV/IGrxXmuOG5l7GWcZxQDD+Cnu3D
i1SAwr9iLB5vwmkWoqpcShu1+RkZPJVuORr6R1Ib6tDBE4k+t5hshFqPQSpBPPQUmtlofzF7QmLe
KdHomrRUpVou1AUCJAz0Dj8/UTwJQk1JcBNBIt2YJ69OtQOu8nVm5eyRcwWp/XNXwby6nJmtCZOZ
uN47T3b03zwbUecLd7iBZcLM3kiephtgk3CRHvV3S3sM2TTDgvt2WmwVduVoLxM4z+AZpnbkqx7K
hs1Acl0T8cQVULbGD9xQ2nvJY5MN1XwiKPTEIpvc3IkTFadPxu8U3IuyL7axwVUjuN1+7PDWoW5Z
R4dDvvRv/31BD8bi542pwUyww77CtOtFVUT7nmnD13RvaDxaNtA3vZDWDKON/6pv6oFvSaVKZcPo
wiZph7Ysqp2ldrhBbHii3oOLMm03az+JoznRkKwWSp5ZtEv5Ohnw2KDorIwzkz9l/BWYIMLGkW38
mkljwZlFt37ycrrOKhbcweu4gtqyA2HBY3oQGyAvTtPZTEpigRO97VmJ1aRerjjQJ0/M9IhI3hwD
Y1NZdOt8+ASpS+cc0cWJKC/4UMcqSWdtWBTz5gge68cLukAUyMPon4oK9EZVKNqpuQAPVY0W1faa
8UFUgjPLiVoqUfvmbOYkdfCYvDYpKCJARyj9sBlrSYf/m0WCm73JJAWNTn1phI+fXC5IHToE9+RM
715VbbAZ3edybuLqMYm2eJQhfKZUgDxLhVNheAu+dcSHPzGp9CS/peICV1oUaMYH+nqMBTa/EKtv
XkDVHCZkgVBSclGMXAbSlj4Hg+e3SoX4bPuTYH8tQ6VHU4oUd3uBE8T2bjx4sqlpLICAJjZc1fQl
1TQztmG+oygAEB+waMIPY7pVr3lEGvW9po4EaoODwP11J1Bg/YiSsY6c4OmqUWrxO99sibd4KHba
xRLQ57j79cdPDHwtNisGnvh9MJ8seuJzG0MGtye1idU1Mwe+LfhYMXeute4Twh2Q3s7r7uyYTcvP
TvBRVuHh7s86/7jRLKqz9k61Fmm//gNyqmIeSCnT7hNhx2iPJpEPncDSd4g0jmA7CMpUwyJl1Bkw
G1f+aEBOJVG5yBlBDDp3YitQVrGmqxm/nLITGukL9KbmZ11F3M6Uwo/BWSgq0dwtrjnEXqcii7R6
5nU5o5EjKYz8SA/BiOsOP689ZTSvxV4IOagFa1GgFK/7W0UlkKrE3cEyQbGuBGoBfXxvaw1jKABr
PuhEzDBfEiFCAcOH1lmHqxfkusVXZDaA6tF+yd51tZQPwm83NceL69iSELjUo2tODWnP0SZRgzh6
nqwR7osbTRMqLw88EyKYX9A3rMcC8FQyYA0dD9dTgCveGOQP/FwiZMxd1fNEZXqWhvq58MAhpNp4
XC2PfnyVhTnjtGHNeybbocI4DnPQGX5woxCVl63Tk3gJyqFNM4cQqzIiu35a8Zz+EiAonSwlAvTA
Ot6u/c46XhUVFWMX/VSGluSyGyB5I28+tPVPgMD+vts872MmfTZQvfS/684Qr4QyZZs5l3eBvLN6
KnGMMpg9LXgnNQjv9TL8i+guKyB3QFIGxRxtTq1+ItsrICkU1juyPl17/QgCi47aXmAFTwRvo6bI
qTsBzyz6fdokbgmc6e0ctXQboh8mFhZgQa/Q8eU+O1tIIWWyL/i0f0fI29cBZxNKeV2UNsIps1iT
zVlp5Lc7q3+KFhpcJV7M6exg87E9fbg9JXUL7sVwgDdBC0bEI29hyxBbwTCnlIOjkSH+lbze9dwo
Vx8XZyk69nPAE82H6jpI/b8ljoVLMbIc7XvoFXxEiPTgTjwbP/j4xp16yIZWEC5p6oQ1s+bJ+zxE
nZo/SU2p8VT+Y0FRmUkBAzgwS4hfkfe1YHkfFvyRBUKpxIaMbiWJApKH5e+TL6mzGXkbEkH5shSq
wp3iV1nascvkfy4uU0Dj7m1csvyv2aGVO5eBN/wn78IrPDhgRSy2PXvG8ZByf7rR8PxjvzwymidA
+SvK476RveIJmjSSiXqEQvoKVm8gTDXJqhKQtvDw61I966WWFgMBRu+9XHhK/mpCBrF+UjFw+xFF
aAi2SQUcdYcObP1sN0sW8KHMvJWIvU4v3RBu8GOS+TQa3x3fJ4vw991a1aa3BGEodOh9b6mkiGd/
MFlWNmpiGvASfd1sbSBn2d3oTqAs0DKEsfkPrlB/rApLS4wraFOSP6uLgpCbw+8M5df+pG5bFYUo
W+BRqZAd7CDgT1J3FI7f/QqGOXJ4lTwf1KdF9MW/5GfV3W/bAlu9olSyGAfY9qUyiYZyHeQg+QtZ
O0jw15i/gY+CPDAz3Of096QF/GkeIZWldbMBuyHo3ZKr5qb6PaY3po6Ph9smhemAgoEnT0R0OVlN
75r9hkHe7cVOMX1Sw9AvqneWC1uRh+Vby4LBRBNjjuVA73DZNdYf0jrytp5MyiZfwJWjcAq9IKZQ
mh6iZh3E1fS/VlibWmcyLbsFvkfHy82CkYKSG7jK2N/8O+GTUBXbyRAdKcHwj/Z5K9AtP4Ksz9AA
BS8GXf2q5FxBZMZSIWtypmcuNmqzBJf9uL0V4I+gMNlTvpngmvcdZr7vuK6mVqhKinc0L6xamB3M
vgKC8AQr8OboSllhHrgu/pA45LNFwvuwMVXye8rK3idBHlLVyXsLPdldCnKZZbK5eHSpMtg1M4Qp
JrBMC4kZUNaZMmk0dTQ7Xa/GU+Wtdu2ZF75BqXm5P4xVgFuk/MT12eNOFdiCRUTF1rDZM2F62uuA
9Mkov6CpCB251c0MV5SuV95ABSW0bJv9tCChHzvJrq0iklfMU8wJju8i3pwV26s1jA0BQ20nJ6Mw
6EiN3DqCyDDlKdKbEbZvPBCOmhMWp6KVj+Zy8w6uDVyZDJaYqAau/t2m86xwLcyD47E1992TnpIn
FXtvvpXkMdXHSzFGZE8uoEJ2LF71s2T/2fjneyScHbK1LVFEGfsOaYA53Jom2UxixrDJRC/h+P4k
Yrn8tcIFiJu6XfSyQn5xVzIKwJO7I+Y0GrCGayqzl3oTpjqnnlhJiVWpMFx5yS6s+oivbt5ciN/c
mQR0tGAJvJjR1RVCTI6WmQ8lL4dp8O7zW6Iq1dd0vWdBhnFr6dIRK+KOzzNAT503m6dZUpSaUmNn
APzsVTRuzwYVHNJlCyEuSkdJzBlIeazgi78oPT+vJ1m3SIGbzO1sT5l/8yDFPIx2I2oIpInHs2q1
E9A0W1EQO6Nmd7SofENCLdU9ELGtky87jobkQaic91w+ouLoT/6Fubf24Whn+Qx2lwYaGNNbeGaY
z2Z/x6OJBPg4IaBDWtJVdNiBFgUlyG732M/xuEyRlUOAxGpib/Dvv8RrL6v8XsC+5pyIIvZ5PaeZ
kcjuB7ZuPtpe7nNVrdakOPoJW6GPFnq86gRoSJiJGCr5yRF1LZ7HYKNfMbg+UlMulFRFhLwGSma/
Gpl+lXbGfL+2v2vrK6BbOEgKH09aq6e3xBxfpAdHdWLBSBROh5gKAehQz0PBaKswcDr1/DJjnE1g
Jf7zn5s0Bn8NWliEK0eJ8j3WxLkr59jyY8ZgLkcJ3bnoub71JD85uJysxDfoaW4lA8SzxT/5fKPW
hN32Md/jDx5ej312zuAOGGO4sthFavTSka91PlqIA6bGH5tY11d08rnwFne4qtfnSNheYQ19lbtM
pxPUOsUZwN7kwQCEGThPG+iZbgQoTBRRFiTBR8lNM/epp44/7hlJiDDvb42v5CM1RgW74smPuRjD
at07o1hztXoZBM1PLUjkoi4HoIFb1pCrmf6/UU1WuB0OEh1JPX1Zc+CQWeU0BWrANFTFMWEq9s4a
tC7N8A1xyvlx5Plws+yZ9OFUnQGZsLeDysSdVX9U24aNI/azRIRlXzfeqtAmKAe1e5y2HqUUqm8U
Fk3yIHfhC2N9hbWRyYeAiH7Z2hjsWt3nG4UoU0cHcMmrQEnRzXcemacPmDHJKVqCHGU8w2WnaZcx
NxaI/ZoxIxgRxcNxJJPMLay7fiEAJekk9EchNzfl1eJghbT4Lbu5W7qp2AjhFYxkRJWsm2ubt6Xl
6NxwD19t/M7fgzmf7f+ZII/AwwTDk6WdkvArUb7YyNQwDePw5aMLXG2Phff7gUUwDqvuESfCKlRx
IXjy/7IUXF7guZBqNduWUhypkoSKFBLA+2bHLpw7oA2iRP7fAKz9Iq9CRz3UQa8Ku3AXrgr7w2dX
A7iZO2ux9tITzPr26ObAo2OFQwbu2URDOOr8WiamrNwaPZlxPHgaXP09QBIbgZ/BPPsXwsFtpleu
KPhIO3UuYWjXXn5U0DwvHCX1heo2AiHUQ848FMVDFqPlxGS//M05q0Api5bCFIt42IulTv9hpo7A
JOxXWHYdxV/GFqC5YdukeTShG61I5PZ22+WbTadb2h+iVtpukDJB36Npie+tSAShwRg3ewenlet5
gbzWwr/0bBItTC+sHytquwAn4kNssUuNYJiCDQrG/O3TngOnOhW8eDQFOORyBBds+pk3qd6jvK0L
fK9KlfNnE0Uznw5Dfk32QPNtv0hAPtOFxwhFQsEPwHO0IAFm9/XeCDoXXrIIu2LWjntdkM/olft2
ssxbC53r4fSvv28DADoa6vtSPeHLpdOaL633JYUkbKpKH/HYxhIwmmzy34LnY6Ld00KHmQ8SWt/P
kSKYGeO5mQvcS6UlQfT+7cKLgqJ1J9C5ucEngRrzqdjCe8hJ+AOHXvDwn1HHLNTuu8CPM4qTYoWo
nCKpV2c/zeCGwKD9WGtNiSlUZKUNndVNqAgI+U2viOaUDt9jo/d72ISgF9499Xa4dByRhcykV4ja
wpPNkT+5IkbmjIibNSFRheAHBnxBPPF5SHs22RZiEs4KoRR823CZ/MIIV5dkPJZ+1+e8/EEePd1q
hBdVSQ4QIZ/5qtakGAJfk7tCxT7+dmam1dB3dphhlp2GLng2W9QvEmoF54cW21lBZdl9wVby1UkS
0BHrmxv86Foxi141PYP+vIAPhVcvS98i6Fxc6RCRmOO3e/zSc8aOUJxdZD4tdlq8ipHxwfDSW1Kl
y9WvGmsWlGl0JUukVvgR3zsLqp2gf4qnDadhVbZUwa2A3FWoVw9KFVDPWgYw7voyEIZOyZvkKvI2
fZ2tagNZqsC7ab2VlxMcHxnPKnIUoIhF7ai4ZPUaFgcqtKVvWPhsNyXMdvESt5aFDLqgGKRNSdFU
lz1ERHHQ2Wg9ToaTInbIDtrDNWbtojeGgVbXlu11qPQNjR0zQlTCoaLc6LmG5Viog9NOGk+nMmqs
wpP1M/CtQsIyMl6lSBnkj/C4B3S6OIKbh41Pfd1I4rk8ftjHHh3woMrFBaMhmlSZhUl17bIgn5rM
Y7QCf37s+t7qUV5yRNzxqK1qSBB0nJhYSoFgPiodLo21wNCXVBFAY29LbWyK1lK/x/tBMOteeYae
gImhghOhoEr1TgEzw9b94Qc4uYM/MnUtpzpRuoSMngsb5asQCdivEtcE6iGCDrC9NpgSIAEqwsMT
YfFUC6cEyB4Scb9Dx5JzL+q3NRy+hP6uPh4Tg0xVNKka2E7t3BMHekh2zS33btzMKZ1K9tpU+Ztb
WYi15SBbq8y7emWURCwdmrhYQDwS1KmrEzavJXRGrR1zKifUo6MISab8GW76ltOUOQW2U1R9hxqm
AoSLGHF7S1K7i3kAuN/6Ec+v02rxaxzj0pIPGy1V5mTgikjzK5SHw1mrrbmghEBzOYNW4ohGVq/G
aljshTXtZ5ey6roHXAGLREMOdTVlsQvml1dfp/IKD83ap9F8dOPPfCloYYnhUT6RbycO60EXXCps
2TmDkhQdWqYBZZbyBJoTkfk24lbr8UlptHJ9ZCjaR5WIfj7xlE9IT/Nm7lJuA4OcgdXj0GqrRj47
qsO/G5MWlQNyFwwN5sretj/tMv4SrphJcZ8q66gHeoGuftqm2z4n/tzkEuyrcihWIpLnRAUzoszE
DPxeiZ7fcrC8/R5H024aO39O80BSJV2wFKpz1MkWgDxQDvHqdiIsGeJYU1zhu6PNusZRtbvrgCps
DIuXD1lenWlhgOKhFGGIIXX7e2//joVSX6wJ2nVetpjsldIYCYlsnX//cWSFpXLG5nV6Dt1OEhTp
FynX8ZaWJzrHRXn/+KrdoVx71g0A/C3HPqX7faoC0Sb5m9mWuyrmqYJZWXSTjOXdfh1MdpmJak2X
nSR/sFRfaSe4EXTVp5SHCTXPBppoRAH34yqaMgI/93+0Vrp7Ra42KsfoY+XBa8bj2QkHT07EYBzG
8aPaz0+zNRxhYAHCN3zJ0rCPY1ImDO2o8j35yyUZQXXRr6Js+QXL9bWg0UgqajTS9X0cWZ9Uh9gC
YaHuUxQMjiY+rOpNn1NJIMzVeIR8/WJbZoQel1CQtxWjEB1BH8uEK/evJMFBGgqT85ZlVSHyjTzf
huWDaKNcrTFIx4Us887Prsl322wTM9oq5DDC7LAWshYupj3F9UJNZA5uzyPrkn9WRqLnDJgnu/HX
ZSZUPkVEfRFRHW/BQ5OGkiIHYpDdo/5w92Ik5aXxv0i7mAedHoZ3uhD41r4eQ3S/9RxmHfks8B7K
TIbOx4ezihaYAnnXoD3t1R7SudQQq+O8LjOJoBHbOMOWg+q3tVO7hiQQnYaBK9oR6twTGmhaKtZL
R4P2x2b5VGF8FKDjiXI7NHmJUaR5kXEKhqgnvR8bmeWmSbHssj+hY3Jr9qTcSaYcKR4g/kxMdsBF
WEvEkR9e/TWcNbOJK6WEkFOZ1oMK+1IGlGLvGhGfNLhPmowzOaUmQyDChCcJNpf9Uxl4jgn5zf/j
9OsiaIVG5w0Gg9bvGGi22Pd2h41pFVWYcMCJGDbgXi3WjoEUSyEkCT4OJvcCAWrJHJu03a6GnyEB
uxu5NOuFoxZBDichVmufNaw6G3n5WO1Hff8UTZqOopF3luh5kwajHX8cgn4TFj7/LhfpxJj8Zw3O
cfTdZv0Ync636QGoyqJvYvbvBFdRtb3gjD0oQ2ijrKSivhTmTuem6dwqETBDzERfDo+fnmhNBxTt
MQmZFeYDMHp0tJU7HVCQVGCVYz7hcAR9aeftzbcE38MdWuWsWDyMJO2I5IjypmmEQDAAoZ3gvEJ7
2CSRSXTA1j8foutMK+fOsks+lpklafrrLtKUMbSDRU00GuMQm7ETG75HIddOzY58ffZcN/IxBtmy
I49iPMy2cjvtK7S9egvOtC9Kc+/sBmDEyFOk5SmHJjewayklzMRLsJliqV2imO0IGo6tsxiBfUIg
JKZcytBQDlXL+CI1dcsdbRhU4n3H+HA2kWUROMTtBSR5XMXal3KCt+l+IDGRlT2KQHpkDoB3x8Az
9qELnqFw7GQWZkxv3kM1eMdFC46GuHFfRYT7Ljd/Ak32UFBt1VahvHGInIjvoh0SotU9/9SCCftn
r/xzCdmgNHGLrYxgzHnHdGTzRW1/GVyE9w6eSwatmjp3dWza5j7jJqlF4/P6kDPL1d41TUjJes/B
MGRWhYt71VFx+ngfb6b8QHYKbhMMNaxbuXFExRyeFOjRdE7l9GSi9Q4L0Vvk+v1LjdOnq7eOtOVf
y0PQdbkmjWVe70rNKbgg/RAMvcGhWzs0Codmy2ftXqxIjBYfy68WZDhol1wJmWMwm4jY1YgVg+Pt
gE5yOwO5sydSz0sUfBrbwsSxmawLbQMF7B5m87A3OBsoORFGh8aYCfHb05AI/dSO2atKeN5at7KV
js1AyGnjliiop6NnF+Zhjs1+xkmDfPyvmDO/KXEyeim9fTahxu7mwaICNl5YqFOrEgFESBQvob3/
+LSl7wGxToCc/s1d29pa/x7914R1WcInYFhrzWK/CxSltgDiO2HYxoW9fH4gmbJjpG4YzbRDYSsY
/RtdWFxn+iWcXk8hiWLzLA5woERThq3dWrJheMclw6hYy+kL7kaTKAqm2IBQNSBSZBoIjcMhC/dy
wUgsIHmAQNjoK490EwylTBvsLa9jF8kLdTpZd05BnoO7F2efm4OMUiLq+iMMw5NsAMnrMfcW2mD0
BEwMoowG6bgy+7kBg6kfnX6m4KM3D67R2A+9wXlsAkrbvcxQQW3AFT6sGFKz4sq5ONZIneZAP1tJ
VXSLVUSqoHE83GemzxomfaGOMAAG7CcBs9fBOKARKo4ofYIuY1p78ZEJPqUGD9ggxGAWCpOFj9Qo
0EGt3If2dls0a3W7qVuFLR8v1hmOrTiTG0OYWk7E/n1rqMD/a+5rPgPDkEl+4SViirJqd1kd1THp
Gdz8VMM769svj6O1/mfu5lGZ3pujc/UJRZyzsUTSW8+v5qY6JBwHe4PQZDW53knNizds7yJe1ivQ
aYBfy2KV+ryzxtk9FinlVxWIxuFpdarHbXmfFqfvES9+8MkXc+EQD8Ah7jesc+0+SRBa3KiWD/PT
kyqHOLIfHh84A+ufQJJB+QXOHtBZXYCM62fZ86jZGHe8zHx8UiPC7Yfr/YM8p+De96PcD/M5jPd5
D0g1H9V4xoZ2w+B9gommSQ9r80Q5L/2zOEMCUMoHmDcK/BRnjFAO847Jza+wYeNOVV0Jbs3Dt+Ae
anZABenoUiplRHGD4hW1W9A/FoXhK8yFVsL7uMNFh1fLqKd+uRtLKw1N/ocvMUA1uhFtICpQe00F
SVtokoUt3SJg0tUbcyuJc9p5u1ux/qakCqAQyRRETsPv3VU/JgCMSxqTwJwuNBotZLflSzaivg+4
mLXQuzyzQfdGDrvBEw0K0qHpMr/1GJYA+TSIavblwtukte4I728r+XZxKuPU7WphDyPMXZehAeOA
heFVkPCBTCx1JsORz+gPjYzVtUC/jz0oRI4jfzYBon/KSqEZCjXsypYrwQYunUWIdGHJI9VhwTpt
MYp4Io/omV3u2yE+lWL75VDbh+e5QNXdbuQp9zlwiAqWEO1LEftrWyF6Uw9YeMXnjuS0vPVrWkYL
Qr4qltPVMv2gSbl4ej5BctopllvmM8zZnzpVAUH/TwX5TP2M6SrnRel7W63Y2uXKLo34N9R+Me9+
aXNqHRtAcTgWsTecfsGKLNwArYlP85qRgQ4lUwAVNxyc4MinJTyQ/JNlAvL9SfJlm7VqTsaKCfvR
Y+z/lJ+cUIZyd/SYlzScj5U1ok6cBm3LAD6dw18V34S0LKEIe3NZL7jrpwnbdELMbco7iqDZ5Yht
vxF+e2++1O7OZkxNR2VEowx9XLwh4fY6pMAfuXxJ9sfBC2QJw9ZypiW8MToRrAql1KvLm1755BX5
4GB4qfK5Te+fQBTtj2oXRge7wxLEb4vGwMW0duzkNeFfRu2FJ5up64S0slbIY/TlaeRKzkkeBuQt
iZtT66+sv9tTGrTNxiqcL0dpQEz20ckYYzRNBe8hgq7DuPchUYt8UlIE0v1CbPYaQktrg38fUQzS
tnfHxy/XfO6+4tjU/7Dm0YnOkkkGsCRFBTSFXY1Fd2y7oErtQ9SXzKosRktTvRbUFDnl+BVYh1CE
TNYac/GGmB7A0cSO0eBzIgylSLjGD4q9w13ZXzyiXz6edgtQNJHgJXzZsXiFFH4/63quymUAQ4gL
zPzvX/3vPPLR6XzMpyLE4PRQoSY4mokGrYsfG+jScADt2Nfywte6X3TS2YD8t1w6osREB9N8eFN5
lZeCWmTw/ogIw5jtWSiioevIOCNKZQkb8fcubJKIZmpg693qIaYxhQDa+/PYe0/FxdGV0XwV190T
t+XTnb5HKXpgMevBe2Zzi0HYs7BVnnYNR8WSFo2DkZKedkWFj7e6ytFV0t1h2OXIO/HRPUxMSLtk
q5u87oCiwGgN8oD9TWFDGeP3xwhZdaXtUUsULuUbwV/ISctL4STe9OOmLQEJ/6hGD+PqDziqFZRH
Pj4Mr6S0CoDAInuW3qtzLAYw0kr9nH6iw6ZwRKAIlOlmwbVpU/dbnowIhOKCHnqAdOXCUmmL5Bxj
kuqoPPw4usQOkvOfmKw7GXDDpLhy8loHGjTDRf9fdqXeZ+Esb2yFdxK8HTw4kwq4Opiq7CwNDWRq
QGolfOXGrpHsEYmjaOmXj65Yuxk5yLE4Wzf/cCi1Aai4/R1TUGLhQhqITi/8JrxuaU/K/YWM2WLn
Tt2D2lvDwNk6/ZUAU6LFHk4Qne3ZCY8ykMvPOt8dSMqSTrKYL1CmfAt+P4UrCEmJwARZoWbCL1bd
fNpd6NAFHA2NW5eMpNW1ldQtBS/kA8Ij+WZ6pseTq3pxfzPWOMjKEvnRClAOTTkkfMxUSp3//BkB
vgWcvdql4iGWEQt+if32s/y8ezXtzFy+wBHILQabx7cAcbDBJaL/m4OGb60Zumgv0Q9RtyKO0CGB
2yr8SAKkNrhwNe0kOCl4gn3sO4hpaRGbBdYtJe7SJ8+WnG64/i4MTvzq7flLOClSj1ET0scwowtV
tW6BabrmTGZWxHup37wNB4h4Tuh4fYeP4Wkn3swxgs4cVl7N3OakX9uZIcTcFB++TBDfmKe19B7j
+Yk0w1K4cvdHeWcDDbSmaE+iLuxGz9dfn4r0s9S349dhLAeK8ABpa+yR8cxun3msGqW2EIODOeuT
YJwDFoYSEz/3ToxJ6SAq4RBI7sR3G/LKzs68JH8ERM/l10oXkhUEKlAh/cfrG0qiF0ek4IDtBvt1
AiavaNJZFFhEVisszyvgnfRp/Eie/J5cxHuhjvUCMuNqXUFfDebguLex/QuszQDga0LRpE2WG2m7
MBJJT69WlisUQIofe+CCivFyXhOofjZ8LYMuJ5gu8N5+M3kEuZYdhZq611MaE3T9o4ue4PZtret5
d7EmOEq7BIc1S7f3wRD+zL6/eW+C7fpPRBHkq7iinYvgFbk81Rot383lzXkooDRXlFw+HE2EN9q2
nJKp4b8ORVDM9cv3xwRGqvz8OV7qnfTwaT13h8F6N8RTcU3wVFIR44YfpD26hQLLU3oLR8lxPcHr
6zIalhFOHOwQmFDztyA47udflwsch1hI+njqZIOOdEJEa3uY4++1Bs2M7OukwxhSj3JRrj42Dpdx
MLepp1kXMntRHSkUroPOKEWYvECCWkll/s0mBGbap0aIV9w6aLAbK0ykYEBZSsGjCtaeTdRW7+rG
urTeq30oV2avA072N75dm2ZnB0qM9xOD9LbCzYoVA1lpQ2Gu1ZCFY5+78DMSyIbsD62zMWbIIH7C
xD9BywCEUV6tKpl3XGHzqH4KXZIRT1YTH8m5G2N91S+REgS0In7w+CASWfXZKIVhDHR07L4kHQqs
kZcKADdqT7iDd6Q7Jd7dm1VAidRPoIIRBcqtnuvui4iRSMpbQJo8+6SUOuPsp4/qneDvrZziQd3D
/bCeN86N3kXiyNyH54ELyomzDuf4tIOQFdoaym0i0HGb1IA7YjP67/9Ed1TXkUJ8nLoVv4mmT1u4
qWZp5iL34vWOVqAHwGUuWy8UAmaVwQcQm4nAzQLxzPzxYP7TOlLcoCtJZoGWh99TrNHaH+aebFxQ
cUZpMu2q2D2m7JR0ATVsd3slJC2DLANgzbcDdDgBCH3A49AXHAzIejzGp0qNjoo4RUNl/8AkGkjW
LLzoVYATOmWQc1JmDjAllsYkexPNIIWc8kDNH2agpRTdeVi32fEAGJOoVRpra7TLLCzi8Xo+HpFn
aJgS8GN4tKK9gQBOfGO/YWQxgHwHeTm/NN2N1fCVqC2eizxyhxbqHyqaCJlYOpriM4OVjoDsspmY
tF0DXX2G0KH3RiMj7R26x6TH6PH4i2tCyjUzL226ppAUMtujuUiziXKhRafObrbqmuIQGyF/8wLa
qouAQ/Wt27cThteDJU8DrGhQIjBDoCfvDTSMFxQ1qB+BCEaUCBWtFcU1Wa+Nmp9yVExHraRerHTx
sPw6UTYQlv7tio+mXkjzJruj80g4IgfYPSfiIoMQ4qHAcZAZKDeC1MQ5JulYLwInKD9A0HgPsEON
DTEwt6VsZYe1QyoGKOJ5GatvoJfjNe1WqPODd7+QlbOdoBJNwDXO0pc/gqw1xExDKlhGY3FaCpuv
pAnFwHHQHdfjK/N/rAPav5dmCaPHDDskGchS1ARQFoRcOYiV6iR0wf12LftFSYXZBhgg8nsX4tZ5
TA2IKNBz0W2nrlIiDiyDxL6Yow5nh5iJXrwaqql3cK+e6gWF6O5kv9S380iWIZcMZGS0CdTlbJcf
31+wfVgrVh1TaavAtJOR5oTK2pp0KLhpk5lcmxVP0Lljotl20ZBLq0UBdCpWKRx73X/dREPW9L+H
ndL/kvqRibchuUgVk9TvMfceP6x4gNy2PRDmSq7Gj0a5X88QiqChooIbrt8lPS6gpY0x5xiYl3yo
b1iU18opPI+uPQy86su3b9Ykr2xdvvjjMbMbLSScOu+JV5uMOdM+ZxgiiQZZfDrWELSHmJNgfczW
GLaShWhSm2KdLErWw1Li3+onUlld1Zh5/I3Zbqe3DQK292UErwAfRvjJMKDb5cwVX0A76uowwYGL
sNbBqY94IYVM4qz0kaohGGyhJLblEV31o/oYb54VyOpa7lEWJ9ZrKTb/S2BvdJdb/Fj0B9JtSKzw
hMocoeRyqZGyBmpBdyZlZkosmtu4q1C6wWFurT7Ty6H/qOfL8QJa26c1SdWEdYDsxidbBg70qBUv
/8r0LlavfvED9S2gherRD7JUmU8DfBKZjvR7s2/8pcA8lpLoxyvp2TZkvDLdimrRS6GJfLSJZnMl
9yoMo+7mmwFEs+U6UobOfFF3BAG1U8XGqs3UrU72LRED6LUymtpkiwmNSUXo0H+6q+3H9md5imSX
B7uoz/2nm4hBHwdpKIjpoYafPP4n4jB9nFHMUbWDl9dPGTabpHp4Wf8I2JdtSHqwcA5wfoKvqy9G
gBffADEWBYs1FfL4KtbQHP/h3McV0rc884Aywr4eHeptQntddFhSFcncnKak8r2dD5d6tzmgMpVx
IVDaXaXoQzY2HnIumZlb7WqxE5AzjWWy0oTELrKgdaowgfdPWNassH/GWREeaX0z5McLEMTNCyH0
NYXznCFORwblx2Xh+7hEAByh95PmcW9otpNhB6gt3zeZCo6Ex1MZrVCZSQCAlhPVqoPg3vuKqw0L
VsdsAKEhksFYdNTuvpFAOE+Z2oqFxpbP7JL41jdUMLNcGg3+C/g9XeS43kUfvWPULBZhDsnJ0jgb
KiaBfc/uDlvJTaNZLpreR2j7bui2REP4oDKGSDRzgLRewu9oRnxYbeGibxPpKFoq9KBWslcr4cHU
bpUy38SKfdrxqO5o8V+x6Vew1gVNBeh84N7Nh4pkOL94tj+s/FfvJljwvKS0yjmWSaMlSjnmYB2R
RlHMVPhlmAQ37lfTNcu8LBgiWglEa6hl5WSCzOUY8SNygRD1AqsuQernJlxovsGRxts5ZO4oIcWE
MhYS/LVDQ5Z0aPckeGtrseFLKvxK4cLZx1kF/FozCRJqJcd3wHIuwwxbxwQ5t2D55nmBkDh+HfMF
fXm1MhWuebQ5VevxeQPH0JhrWRE4GCqmpqWN9zIN58SuHWmBX4wknDqi5guZp6jcB4KJntRY/4+F
wDAACkQOQhyy9slguGoycAPpD8ErV3vl+/iPWtqYffuDJ5fup7vh8tVCOoaWpBx70R7b6Es6VTry
uaKcf8idiMhjZ+TCYMY4yL9XGMfFvflLWBFKbVbFpj4r+47onunbV/bl4mE6bSGUAdh/SWnKC0Xe
wbrtUUXDIwpbAc422OOwLukMt9w8LlaIHq2BRCNSCxzzGU8HCRqIUJX/7ERTvAjgNxLD+TowNDb/
1kos6RmnJuyOKTHGLRzcwKJgBRIgt1z+xYYYHvOmyW6DILYfkYNl52qtL0/aOfLpvk+qtCdsvnvo
usRDImItmlCtDWM7t9fm0V0pSSzBMdrlee+l+k64NGyKrvqNJGqUrIOCmu5sYWpQyCiAhLLlU7Nd
DpcZgOnwTR57V5gAQ4agy7qmzzVscag4b8jNDL2n2glTN2A6n/JtXyZqQTBhudk2cf316DgFLHAE
JzeQEuvcuL2+1BtI5EdkhmpbJmvfnSpr7mn+X5jLHqwhrPFfLJBk4pNRqssRsVfpz88sx5+eXezq
C/Ema/Zqk5vsbuqVXF1DxI1+ZFXNeuyydlPR7/Sr/7ppdRiyzaewH8V/MU9tEU5JfMv6dZEieVh1
x8zlPld3uSg85bDmJ5W0aofXvnijAJPuBKL6lttIKgM0+Ln/EGuEdvigBhzv+2jXGbSevHfw7QBU
+Uwav0F0oN2ONYNu4ehHLtUcc4i5WapuB3XyAXianDnkXze4VeeO1sj+fy//nshbIvH++6708f+6
iLa5oqYGbHD4cy1NYvi0zDfsfEkfLxTXHh2PxxocT1Dtms5s9YTxzSQT8U8f0OiUd6NhufZ3v12K
nwuQL1zj+WqNcUSalJ9syM/ZQB4ypC/h0Em7XCv7F3JIIHOrBQ3k4DGjL0fqtegMTxG75T/Z807W
c4278ref3s+E6oovtHscA+WG7GDfYXQlUEil5JbmQKIgOE+sv6eR5vy4FCk0Gxn2ZKenrirMrD7a
RKwVl5AQSCt5fGAzkbYUFIH/hS4ytDBa5IZvLfg6aBQaeOZZEq4cc3Bkq4jGJEuG/7s9Dmsy6fb5
4yoZBfSBc7RaVssQn2VT1dGbIXWYoz5GA47y4BnS8v1xTFqVVrjG5dYUYDWFvd+0urk1aDBO7Zqb
QSTdxb9SOfJv8nOh+Z7I3cjgitbr10xZK+RsfwI7NxX/QVAx4wj566I+ndfLuelUKJBDHBzHUMfT
O0VAk60qhmL6cyN3xtLJBLVmCZ35wqt/jc9YZlWiBXSa57wwuBNiIfx5tVQtk/GGGcHHSxKck9aq
x1oqNdmIhr6g9lUq1UJeORS7SeTb2cfj7vgr1UZy0cfKPB9brGA6wAwViiin6jUQWWjWlYY1C9wz
8fzHQKDR81Iu/TOC2Zk5iu3Hf+vXeCTQMCQmv/yhgqLGydgM+S7ipZHqCTrSircPaxPbJuKmabwj
J+u6MH4P1nFd+0HI4d5KHkowZWltIUM9B0+54LWWvqUkyDlbfL4VDfEk2AglUQN8wk5BNHpJUJXu
NCqgaFfAzg4BDoP0R2nrn2fYOthgjLwuKkNeKi4yX2X6Ro8SJwsC47rocvTf4ccdntxc2Jx31pzH
JozWjOZNW+ze7iT5CtHVlHK/5qQQ2qY/UZT7B1qub/yDKhX/ZWtItPdvDviZ8OsFY7ejrU261MQZ
eGiAnuFGpz9rRvwmKgPzIunaDx/bLuE1N6sGL4fnAO6RCFJ69IVwkCypCoL4Cmr0eehsRL1t5T69
EnfBbhckWChUWbR7zDVUXoBapN/iNIS7MKFa8gsHQ9If5olEPWWsmjt59jg5IdsmaBS3vWG4ndBt
p6EPJ6+IynoHk9fLMaihnMqpx5ijYB/9gqdoDpeww1XIaOYlDdbQ8T4xobtOvXP7Wcf19aCwsazT
3sjX+uXa71HAsjnu6LYIvGBuClUHDctlAEnTUSHIFQBLAl1oMIcvu6C/yRoEj6XTG8MF1E3gMUyQ
R9VesoEsKQjYfDDEwzuNOUzqAMsPkzpl9yCuyxanapzPSMXi5ZBVCnOCuB12i6Hewpek1NyhKtnX
ASralqOK4I1bGq9ul7P5uWqwgtFJsBBUfGwznUO05mSC0Lq3tQNoa8IgcHcMqEJuNl8g9mUvfvTM
0YeH/tGYNz8HGmOgy/zLmXgjN0rJfoglgp/lHHw9VK3+u7tER2m0lDmz4uvPkcpNAiVYqaCln/Zf
BBxeyDjH97x3VgAUCzRDdAD3tjuQZxw5EfiR5TfVSFDN7Re7smZMUyssKEBrkdNE1Ip+FIRWtv5u
Wyh9gbfreiasn70YdlviJuUaIVNdPM/Yf1b5QY84/+Vgu7NXnClbA5A1mlog1b3A7u8KiwIFio85
iBVvGj60xu+NtblE1wYu0iuPMvhInp54izhG/7mwrkRY6+3VsRFgaQg6uM9OVwzFrfBaNP4iHLs9
6vkDznCnbxjPIpkXgxunzHT4dyNvUwSn9MwcumdoE+l8j8YXabxkq8AwmLjhuUZh4Y0ToogcRo68
hjUqFv/Hmw+nCrWQcooxZTLadeH/Warx51e6zsHSpkGe+0DPPMRElI8qxiEWeHJTFr1GBnh7K8UQ
bg9KgZKb4bmMxXllZ12pbLihIQbGgLSUlka5ct0/BFZcD1JGd8FKaKN7IoFUIK0Ri5K/IFi1C1mU
gmYtsOEpEomS6xeMDF77+kqn3jehE8rEfQ55C9prgbjJYPG+2mWWfz75Z5vp9PIi4DqQn9G4s5IY
zIhGyZ02VLXbWRGh84N+j9ri+DOCL1cEVGCUEXUR4Sn+doIZmLHQiiPXRoQ/3EBAOSl4z9tzH4Zd
7bCUT1dikfvsvEdTmHV74OMVtzX2lheXm+vk35/UWOF8gdCE8Oac5USa77yW9tn5VHyyqoRxGuzA
S/kBBpiUNKJykCW4450ztl8zJYxqJxTOASyj9nY0xGsH3iGdsdE2EcAmFXSftOtSOPERGRgbAVpq
QYR2IGfkX35vzJR/7nOkoWQfqNEQJZe6b2mLNEv0MK9JhyUyuM9pqe/4REyX6W0F6hAusn0CCYXC
Yr6HJNW068NH8PoIiuU8gKc8mJcXV5shjHW4ouObiL8Pi2LLfA5NT33QT5Xm1HvqyQIAaOj6/hcq
2hdZ1JZX+RO/givqg1vYJs8krxE28DDK1npzYjkZl2MRI4/BPjNb/D0OYiYf8MeUmaRbwB6GYfwm
JxdwpWDFXTnOi7/5UT9cmnlfBWmH6HxpKWGEGrJKYxki+wMhrB0OjfeoBzE7iLah7odwh7KmVRyC
vOyyHgVi866aFUrUoeJFiXeQwGqScT0I5wLOpMDN785AhghoxzAKFDQofozP9kd0P795v5cDX6dH
4FTut93akWTTp75WukHKKivUkkuc+VssVijuN1qcZCy75jGMF2Nd5e96/ULZBNpS8uThSj8oJs26
uBZLX1jnQhInSPsTTm589I8Bzr2TumcOHQzfsIO4Ijv5ys3XLZcGy7xjiyM9+wDly+HyPa8T/xUu
1ST9rTKOBnhFb6LOx8bjnXcX3WM3k1MgVFsBa5HIowGCGyMMqVVRbDxFMyw6CoSSRV1qiPnVxkv5
1jvBcIMAda3GGQ0JMaNsi1U9OkZemZjXyz/2uiVFIo8xZwkItDoRKelkWrCQc/2EHD8y/eAcrjGu
+1SwOBBbOau6gLuzK+HDv3JhMg3g75LsedOKDdkZfj1Ji3sOZ0hB4+DxKF3nnw1Fes0Q0LFXeqdt
eocQQFfZHV+WLAvJwWX39StDxP3sZKooZBTK8Ut2E67Fd8Td2BCxppI/razJFb2C2Bp1wIVd8Hz2
kiu4C98Kzfh6Em5RlOk9s3lZwswq81T7INPKHTzY03f4yOR+5MaMvYnbQxwbJCCK/F6Mp7U9hcUG
3p7oRgCYHQj17jlyr1hy7BFpYO1csQxuiy1x8QhhndtizvtvFTYZnAnUSrHYAR45+FyS/wi8dCP6
HNJhfanpEHGNWxYnvtLlmV/9jH6lZWwsGQphb34MuCQxHmgX7whWqAu8XxySfAJE3C2Z8F28qGs+
5cBDpi4/lF3mA09g09U9cFPYYydjT1Fs1lNe0XNiN3qZ3zIB/l+Q2Ab9Iv+EUurW/mTOg63EXh9G
D9RK1xcdD/TbBc2REb6cukhrFwYSx1pIkgnXtV3p3bU/WQS1gwmJxJuA5c6S5BhBipUTSQRY+cnc
bZvNwH3t0l+67NHd/5jSan4DgQ30reJFf8RLF9YsMN4imukJ3IIM9OJ4lx7D24Lu2HVipQISyMLK
1ydD+wjP9NlJWWZplhOBf5s+F6NxNPemNAr0b/HpFshsOD+Gp9Ab5YmCQMa7n8QM3umIbpY3OEN9
DCeATIAz/0pMZnXwhf5OKusibqYFUVkg7culqz6m1CuWf6Ss8hMdVbGuvAhpyLzbpGnwl9xt7Bfa
nOiIIAH5yagSCxtFqjZsdUTBnw0DIykHC/i+INcGKASIrgSoxteXTCu5SZc7ZvBmdYtjDPtcZJXe
99n2vl6BRMCYZkzSOdi6bSK/gz+9J3hoWI1itagLhVasRv8nxIdwJcbxxsSWJlCBGQpzrCFS2mS8
mG1gK9EWRQbMx0QFevoQ3OZqEi5W+vCs25ENQ0WW8zb32xms2B7iTKGHvkuOn75WlRpNOci4/lpc
tE54SAlIXCyDnv+n5sqM8agF0KJ9fIwLMjNXf6EHomuBGFR2F6Mnv/mObZfP0CrTs9IbrJHyZDx/
fPYsR5FYlTCtBldISazlX0dgYNksR2e15nG5D0e0ab/NtAdd34rtXO8KOarz/pN4t6W2SdqtnKeY
VAicYwz7o9v/xqSdl3dcIV8UfggQ44BfFB2foTJJeRaEmfb6e9jUmh6BzwdZXBqNJ/nvluN3PZxa
bSDN9v4Sz5fnsl47hwcywyyTQa6VzjGawEa17JqZWHO9HxFF4v+JJmoEDmEuqjfW+pHAhf4q0gsR
bcIdzC6jEQKOUuJhHlTkUj4dRfawnHRLsLdaVWoDfi3jukckvBHOdGIdYOg1V/30OgseB0YSjbPr
gP5zmfOtQR6y4dEmlzkwDw4AlPjdK1sufk7t7qEBKjHpNywoKEySAeEOm3xS7k4ou5s6dEDBwaVI
/sjB4NHXMqndRWKIqt5fRAL1u1f+43jf0p/I/aIxkn7OFReOhDqGodjHBtIcpuAldWASdKt+Pgj2
O3xlBmhW0sAis76ZP/OOBjE4zSYHdzfdMTIAMCvdw/H55QVL2WCRhY1rTKuPdJxvzwlJd7BXg3e/
FJYMjuDex8GEkfXPaGigCn+8E+eHWrScJJib7yJm6uApYlk5qE/MDxkuuNbeMymOOIX+EBDJzkIe
WlzBzhd9VeGEgsJrQ3/PJIQwbS0pIYEXaucPiqC8xzBAPy5dA8XDkToGyU+zBzCUuT2cnZyTmztx
BL+u8z3XdMs5pnHDpvwgwNuLGQeUvi5Xx/VY18bg/1VxXOtJDqEiFROWP33qZCoJnzufUAN7gE4N
6Bj33407vdxecBGEQdqxPiAil/PyovoK0c/eq1QEVh3YBO61aLPFcnY3G1/IS6BySCQ6Yq6hL7aq
aqGXWKUi98IF9anwWnRCfvBcS2c92/Gn/icTVcVYzSZMbSgYcHVRinyM3OGVcb48BrgjFrT5hHqR
RN4WsRyX/7N70HWfrouWVo9Sx0C9KPiM6BW4dHOOy0Syq2eeAy/JB51t+PPRz4BjVW70EPAGjAJY
SRqYE56pc0i+62r1fhbk8tsYlTAt+uTpCyzKcByyWk97aB/cR1pIYc7r+dLaK1pwNSka7KiSA3/j
dMCSw81NMVB8V4hq4CgCKYgWcY4OuTCt+0YWCB/Ksp6AabsudKVv1up0kSE8xzuKdrYJpnFAMUag
BbipaNPZauggT40+35LRJ2ynnFEy7qa12olwUfUeyh2pb31qVBMIBXD99YUJ+cfxWYH3wYR0cQKQ
J8FOGUCpwzuKxgMjj3Znhbod+bsjuOh2mCB06uP3+lHFPF4JgJLyZ0RxIjcTMzDYXFuApUmeIrU7
Y86aWBDh0MQXiG+vihKp56r+8OTDkdUmv6f2WA6ungeQwMa4itEpHQMA1AqwTSWZ+KXirYw1htNV
G7CQQ7F+vkt6FHCliVaCCvWX0nomp/l6+ymSvWhlAfaqGB/FuGQCae/JJWfvSaBEJsSkxzNHz1ny
1Gv4ywN1DwhqdOTViiie6rfUPNit4DyL0ZZ2BA1jM5pj8ns1W+200gGz1LwBfyVtnYffWa5j7biK
gIzvCQ74zKbGLuaSEeX+O/kY00yCAfeQh/BGjg9xuDY6dN+y11gADVz9MOhmbL32SyDnaBjCGeF8
AxKaWRnMBFrO4psq/rvWmsjH6ti5wiE2ENeyMmojEynYOzzc6Q9Yh1A1XqogNa6xM5XZIS0aySc+
IvJyVR9lJ3qS3oqFRDny3lQ1aZk/W56ay4CiNlh9UWvXI8Xp820imA0ZyYRnSLdFFb5Tu4Hqe3gB
czHXHH5AzhscogE/laO5wIHMqAjzrfPvWAveuH1Ga/Z8wVykoSmrb3rb9D+CaROV0PFaQpwUwx8U
lb+L1TTbPTolXtmKlGKKGkEqyWhkiMH6TZ6aMRSWR7fgfhtc8BzlmO+qIbz3nkRbJLE3DfEg6nud
W5ZNDcn4UdpucfC6Itok6mvpUP3oUx90sttjIFpsvr1ZoGRmQS1kzqf9IizWvBqXN+/tTYV74PAP
IYQu4kBRKEy9PQ8zpepvyejoxXGeq2Ylgikp+b48biBM2w1r6bwIvmy7sWPQwI4NK32QLMnoBh4T
7rR9F/RUYkyOJEhz+qBCBGP4+LLqJ9MoXrqvKdj5UEkIKONJwfbtYLEGhVfstqV+1OfFApHYr/pn
u9saRCbihW3G+5AJ8gb5kzmBVbU6cNtcJTIy70NP2em1dqwr2UX7rSb/ZIavtJ40t63v5+qxii2c
dooSCBoXNLd1TVzjyqXsAbW8hj5MeCFdGDYCw3coXgT077k2XPVhCax4gJ4fG1c7z333GHo340BI
/7oOuQRXaE9HONoWlP/MMFYmp/l+eKeckQJ4nvAtFhuZpymgasY024JBkBwj4vHMm+OGlbGlKUaL
ABkkzN5K3R7EfjmiZHnKZ2ehkrzGjSSaIUuRvs9JDHBXYfdr83fxFBCe7KzJ1DJ+7d/7+SUyUFWm
bzBjS9RG3ndi0p5woZ79+l8JR17JAKa9sIJkTdqfjbRPnajdzM0ysf3dbzMwv60p0k3vU8Vssza+
IPzVMz96vNez80fpVQYLYIfg3+X1wntqnB0Z8lfqUvqXc8+FrMSuyaTGnkTc4WVbni2MaN4mny88
q4tOdhJaMDbmdtzG18nxLSs8647dVslETdzbCDdHYIl2Jck90gOxxkjL23OCelg9Agfviqt+mUSm
DhOikEAqFv5XCDyFXqB8gorA4op1eytljW3JT25qLNJbrANUWBBXCcVFQwBIGQLIDqZ39RJ1A4ud
22zeKImaz2vSgLLUYGWiGxrBSJaovU4X9DWXkzizdgQGA//UieMVHJc+IgkhnsxWnG6ZywfG56b1
C+RWmDG8ooxmUZq+Uw+fzAPKOIj7TwB111ax20eOgjNl4k422le0aUtgjQBTshueRbzpRRVoZ+n4
Dk15/gST36Z1MlYMvdCx0eBnTmudfusZOUOjPoLaLiBitcNsI1wn/h9h/BUeUbF3KneJ2ZKswaIr
LBmd/DD+xxML9MsKqMbjgZPCrw7BeosOEcjvH/rZaNOhiR6nmJtAIPk5H/D4FP6IEi5HYwU+PMDf
nF9IuQs0cg26nEykpXhEH+mVgZsS2dagJQnZBLSDpebvUgiB3ki2EWDntI7H3U40vRur2e8Gt1UB
czXXnyI3ibQ07moHs1HF9HXoSBQTKKZZIT23eHfjLrkCPCPnD7+pVIf4X5sOOOOAqFi059eJ8SFH
ZeR3O56XATXIG5+tgG/u4wHOBNj8JqimPnhUfG0ThPjGSt/5lNOQBTnFoIIqDRaUZRi+Lwiw55oh
khdAb+9Ad1ZnKVFQBEQhvatChO1U2nJFPztBkWKNpbRZNd5ly/ZUpoNP9ey22ufe4DDvjalJMHXj
URD7Oy1ARKWVm0pke4Bb00PzVBlWMPo7rSPDo0JUO39OwvHENax5CEEo7gj7C5A3U/MnPgw4j1ct
w0FHzIbgs4PEkN0QJCu5ROqoxGQbHmWmLXycxgg3+75BcFcWTAyQuoRTXaUR/z8tptM0LQaoI5yr
IvvHu5i++VTjn1OQNnU/4/aclghCw3XxvERCw2DzNPmAvTvSO1JeiQtVUBiA3aHTVtrH6ylfv10k
LxNqfuKqcD3VL74lPDJSBlhesJ0h/lAksVPDdRebeA4tY0ZelVd2/z4J0OumQ5JpKvMw/A6x29x6
spl7bwVOjK3kypX07eGWyjdjwXvyEjfwpMuxNjDrA9a4KIepg4fqoBaCmcYQW4VcpkGF7uRuLgvT
DkPtEn9CVbKdAk3QowZBIRsCnifYwMFHpFzrxq+HmwYUUdd+C+FA03g+Ypi2uDGPVk0VRHveWMhJ
0m57XnfN5pJ896yvdQsu/Ng+jtlQagDAKyDCOonQ+rZz+U7xtJigeBQscho5o6itqaOP21J4Vuny
0JGeYUZISwd0AteRkA4lNSEDf5EeOnX/PrUTt1dOKqA0+YXKg5rCqSERyuyTX8iVX2DjdDOOY3ZM
LUNhMjAmRUMfyRj5vMiusRbkXNjdOEiZNhrf9J/mb0+lWNqXbcBh/zzxAfvM8ZiXzxvqsbmNfrCw
Gg91O3muAq5sueej58f7mwtV3kol4gPQVSLExSgjCGqMF9j5aeBg1jrZgi5wz3LVwWDLCF6DrUSv
e9JRnKfbI8GhXT5InplQ0EgsbOqAVzDEZ17WlauhqQg944LVHomqCrT8D5lgsEe0Kzr5fkoE/eUX
mtsSDUa4VU6LZVxpkRresjlcTblB2JYw2z74hMdmPoTP1ck163O+iozYmNWhUe8v+O1dyq500SF1
ENdNaU4fxMg3kMN9SDgCR/j1nwMYgqqfUVwPU2kH+mftMBzBxvgSLDk1n4T2UfoIoGnaTft2fCFN
xLXSBBxL6UqFhC39Ec/JxdHKuqucP+wtf2+17YYFOfD2QpLOwlX2mLBvaOcfft4RsJnTYVIKiqJk
pIIikopqNmaCNOXJwyPN2pH+nxpc/+/72MB1Ak86DWBaQK2WsZdLzws5A4ygL1SzI2EfO/tsRtK9
NWq/wDXclhUrWp4qWDvM+huyahL06OpjXA+MVp7DLMDfil4xeF5JYOJrJTmXxw+1wneeNN1OO+ym
6QxrJQfA1587v3DZOsAmdQPDz9K6zdPBVam8+jjL30+4hcVYTksqBToPKD87gAXBgRmfHEUqvpN8
/B/2XMTyrhOdK2v0LH+oFvB0ds/9m8mzZopOE66xGZpHOL/Ij8G5sDh99KgN19juUyR7Ql6eAy1O
1HWAtdGopCGEb4/m/P3UdBLrF7h0fKQkxJ3Ha8/a6yX9WIWgyaTJ/D5XH3huIrq2lRsKcC+B8LDu
i2Ezom76Jn8rTj8eoNuntflw2zDC6S3T2nS4+zIQt0sOqpK5t0k5CxTxjyOgBYLkZRS4UmNDUwBY
b0OgFi7E9LtM5yVaDyaquP2quDLJGO22UB+o0qHHCU5VWfKKkQ61xVuYe1ShW312IjwkxRtLUg10
Ck8dHDUMoxvMuN8JkNbQn8MeQDy7SIKL3tYLCJHrYlOgzMahqbWkDswsWrmSSmtqDD8ec++F+P1N
4UwOqJ+HYBihV0Zb4ouR1eLN0wggM5/1zNo6DJDnFXFNNk5iPAJ/QoQ6s+DssxafDQnRbaRqjJP6
yXTN7/hBFWefEDEvY+fIjGUtq8PpSmHYnzmz2dYVE3pDQ2bSI5wBZ7VE0Oxcr0jdXsvJngyOYt4Z
U9RjSJ3QTbJZ+i44++l0GE+FVDz5xUHL70cqSBCc5GTuqxf+CIq6i3pFYmLdnpYsbIgONGpgiFTw
9jOMJgSae/Bz6UzkVROiSdrNOvE+f5diyoZxX4g+FfYQ+G1IljqeITbBUftJBMvApc0dpuycLzmG
zvwE6p2wOL/N9VNWQgFPrI0qTR8VFMQHYnT5jrTL3WN7Nj/tJbaQPFkOcy01f6Alaq+ZKuxuQkEF
7zoN360W1MbIeuGdmHX74Oh/K9x59rRO2YvRJi12h8yzrmUESg5t8mo8D3WcrAxhy9ERThKqIEx7
X79sbaOMt124aC9WcnGmuJkjPL/11+obEqAvwd44FHwsw+hG5l+uYDqwsdixQZD2B5Uy5TwhK6pv
Td1JwkFS+xhuNgcAetABcjIGAGkDc0vw+qy2plB+La0BzgPQMoV4RsP0UGX/FAqNUqykQvXZZPIp
r0AAQloXcOk2f4M4HtylHGJeV2bTUJXE62JR6MA8IOjnQjIbhCa6Pk0nDut3mvuBKYYEJFU2vPxT
sfM6NaKnZ+eSRJeY/US4s2zGgFBpj0TLM3xNVHaTbeeTD1OfWz0WMaSWcKIuEyZklD4Wq59tFJk7
DU0MkRHvp49fsWetdfK+3dG22mMRUXHs3I41Ux6RnSsuJ+vpbywc66k4r4PQstkC5OZJKgJp1h6u
EC7/z7PkfmoMwARBRzG0bdoGv5h63NJXxK1gQLCfQx5KGNyPB52sxdMtJiXL/4o49qZ3FhaAXOnh
9cWtcKg2DbnCUiSPoZWlV//eb1Lx2H9KDJfXSZqlUaIkGTCHa9qO3f9JDwPX7yHf++HCA9qeJGnc
W0hLTsfJu0hpKi7dSBdOEpY4t9/MbmDM+ls1TpfV7qOYuixr14sDGe5CDoQPnGUmoQEgsGDHavmS
HfPte2fqEdmLu2nVW75aEMcBsB0yLobtrKrClOQuchpaLGL67MfXE0/2QaZ/utuopKozzXfr97kn
6H1S8FLfGPPo3gQxbX4fWV7JCF+bydyRMt4A689fY9qm5uCA21A2gE8tZY2b+typruFmBmrlVngX
hhnZq1nkktWaMSi9Frbyow/ZAjNzjVDh6SjmFNAFUAxkWY5wY7uoIEPqxSZUK+Q86Nf96Nq0awoV
87hOeuWKfhkLgh4v83MRaHgN7aX3z9JXPL7+y0MKtnyFBqmLfeVnE1jTiVhlwM+bkPcv9A112EUd
0fA82MQCdlm+UCZf6+sxFuFCGri8j2CeBFIGNuVhT/cu65Xgt6WJim8zgsi+r524+g3EpQG14WMn
75zx6n1iL12dbiZXiw/phucc0YWpxZDxsV8VJE8pDm7Oa5s5QNJZJIrVuiUw4/Bslt0eQpcVYCRw
w3azziujfpssfxwWl3+6eYci8Jk+pYbez15ask3CFOIn7kyrbEy06NExpCq1lNKGzgp959drioVC
QGQVCvbyIzLEFsSmdjzTm4IGwDBW2s8lckT4mV+GaVQu1dVt0zvotcwZpC4E6LkM27aLSX8ePm+W
M0J+CjzwpWe5T4fmgteOwpfjj1DCvEcE30k+PzQEKzVwuxVSp6WUZSgQUIJaL/dBttngA9xUAtC4
S2Tm0f38u3BZD/bIiMdoj8Y2J1WGSBerATcy6cHI/5pR1mtqd0flgPDRKn6ybU/UizVQZUtsN18V
0HZ+bs4siHHzbLRpz8ZYXwmYTKSMyVsPTlF+4bWwQaoUDgPMgKFNs8QifVrKdj7jS4FQMVU+LLUh
nmY4aykUM2BPY/lMwhMzuLNfXNhpcvdR5TjgDrKhdNZNDcu3dlKr2qitq0H/zW7rPsHq9vg6awBM
xG0Tgjyhr3acu6WoSRqzTzcD2oHDp8a07+4hF2FKQRvuQLKaMBQDG6Fp+0is5aKJo5D0UeWId3sY
hjAfANljdpaokZYZ0K/BX2d+b5Txi9l0TPwrOBdYbAkngqlXv9z1LgKSj4rJufO4xudUW+F2b+gE
wUjvZKQZ2BxKW5jw2uMkcBQziB4jpp3nF28Yx+yLv/hv9wbrxnJdiFALajZ1z7QYu7rnClML2Y9V
t/fTJwgNOywqV7Wdsc4zjhlHIS/7/1xAkxjdyoqcMEz2VGgjSzPFrEbX9NBYxP5seDcEu5+AbXJx
kYow3ZOtSu0U+vRsCX8HjEIJkuC0HTC+E0blfQUOTSMGXdKQJfD9Ojsg1jEf2Xba+StFvzvOT967
4kDG1+DpMAROE+YUdYEj1/2i+Q0jw2ufZkMKdiVJgRHSDnvbYRPMTnPQNMfLkNpuCv66gMY3+s/Z
bCJEoFPMfsQ2sawOksWWXn2quZSp5l/8Ma/oBePkbrTjcxXiZTLO0zx/U4AiA/GW4pGpWHKBVnlo
cOB0xQqbE7EjeocPW/O08ST+BgRZbE+T9DmhpjNxuWYcyKORhvfbfKd6isTf+/Fkk/Pb75P3+Y8J
LyR3e4i3fCTxTzc22vvwhtiJ/YHNs269LPHiUTm1hHHqc7matJ8viSs2JNXu370hdvjlO+esOWHt
6ZSlLdfexY8tdEyWQh6qvwZZbN8J6xCS6NBLal7ywFVLt58RIQpBg97UKrUkjxzqsHgQ3zC308UJ
bVMOQMBgznhwhmG4Yr+qvdmUKJFUANmH1LBWYp1Iva3TkU8STmRS9A+VMoe33D/KXZVlxy7/WEEL
m3y5/EOuMJ6xpReMZZI0z7ZI/bx8xBbRisFzoy5KPS+BrNYRgjancfVBS9iPdy2w6m2o/iLGj9p6
tRZK+omfLHl6aP9XSF4NaS4iIywMiLoVz6ZjozxkKFdmaqD57OIpn8y2dBIdtgdjOT2dDnDNGNka
6NtpQSkp8Fq2WW5cU4hJ1nVtJkw5kL7TPIEYq9DrMLMsiD5l3tuzWJSvqA9IxMmfZBPE/RmM0loY
6gWN+EviGwHAjC7mrgyqN92zqSGEhT5No2vyEluMZ5V/JlHb/w/UZgHG3M1XsaLggLUIebtXdUvy
dZbTriPgwFfvLNLpSuYXBiIHI1V5f+o1/wrqmNMuvIP0eNab5XkyjVKzS3vYoHT4ZIduMOykn4w7
VKy0Zp/9PIrQlvv84Ie1v8zQyi+JUPlUWUdn8RRx96/8KERg+xhM5Lb7irtdQd/mER52Bk7vhpfI
FNIpMB+i6RyT3q7qNsEIjeDu2oTKfZc76IFpZt5z/zoNLZSzWZAYHYl5K8QOzbxMT+u/0eqvfzfu
xMsFI6DEy97cd1efSqj+vUI/eouiXTSS5DMuxCjfuRPY4w02makhRL8oG/HGeO7kmnbaTCDBDc/+
avUnrMdcz0Pw6ybxjh4pj7bL47AmR4vcxxldiFGJkEf5lifmD31B+3BK7hUjh6WlpH1NRjFWZwu0
nTPH0Vd5hDvKlJNvKkNjhe3Ue+oxDh3qAPgAEHAbFSa7IfPvVM+FkjtzBayPA5UKZhLk5JxDgbil
2JDkMMnQST7as4zX25iGJCC0Hn6PmWfLqzKinVGJAGczFnQp6Fu9+WnQUi7wtKu863PtAKejRTwJ
WYP3Rf7OF6DMUhLbR0Jda0dYiGqciFyL3SKCJkmaLBhUpITtwDpIF86UNHBnZOqA9zsTf2tqLTae
TxVyWmfxnq1xwHKabFIWYl4NOVxpI7LkrujA/wZkTwBjEvUnUZoOuANOvPW2gR+BND27WUIwUZ8g
VrD0zoLAjFUvxJ3xMGJEHCBQ6rggz6vRq+PTNPbgkv5I1clmrBchtMOm3Qz7s2s+Ugarg3wf8e+h
fAdG17350mOFi7GJQnfjFsmjtFAu2HGrHxeqXC6sO5H+7vPy3yxRuDBF/8w0oYN3OUUSlEiz6zxY
J8OeeojfJ9tIF0yAat1X1fp+t7Xzr74aqLeagKjti71hOTqz4VQ7qAhTyxM2VGQgiXOav/okhW1t
1u/gZsIs8moAaQZZg8lbPOR5cCtpdF7KxL4+F9KuSS5wR3g0wVOCgQ76378HjaYW4da4RYk3WJju
4xWivw8j6K231aaXTAx5Rd1nLFRoiAWQCAkcSD7VJXTNRaW3ZNFAr4HL+z+R559iBZ0d3tzEG/ar
/r05J0u7bLUOj0q6guAilNeY/UMHSr0aK+fPb9x64k9aZyZHkQQS82SsUWeEb3ZQEjfz9MqIhxU3
6OsEn7T+Vt+UkuWDOLM4zO2OUWSqbfDGcRWnm9I6JRrwiV+aS+17HsUEULwNjnaEiVv0l+c1KP9h
nyrqwCkuc6A2wBmu5HTJyix9BDg3tXJN4laQLKCI7fQc6JPOswYyRadb8B2pTqZSHB8IWKUNc2+S
uzDI78cOsh0IWlLjtNAmE7YzrZihwYmTd/AU6fRNwb/U1jkzobx5WVTTI/o4l6C6D8rjObAD7Yf9
1dtkJ535WNbuhbIaGwspF//Wte2vt2UgaQnm7KLtY5Ve11sF1nx1n5TzVBzEEKchCQEyOky02AX8
PaNQshaVZRd3kZhISQcFxr9YA28cmZiIozFRdKFbL90zKcYYZsC3osofSv4mhaL7vmBtRrYYqwgA
TLGgzm5XSJP60Y5PTDwqIANXY9CwO820ngtFLfd+dcjERzsLt8ta/45VWQDvOAOSOf/4aYGyC6tI
GHwcxSpy63xTPJaljmdzVMemQAoP3abB9gZV3BVmYIxO9tXmK5grbjnsTKpCCIQT0rkdAx0m5Nbg
jEQuKC81tOilBtWfsGPWVU6L0jVx+cglrD0aEgnkNzQr/iApZNt39UZ2JLT8kGlHY6o5AlZDP1kG
9hNuERTPdfJ8LlCmhFRPXnNs0GkUJjbM1QgCAB2d+UfWc/H4ivMlX74Dry/BqxAaIx6Hjo1UPsg5
llwtzyLhjwxOblxSrEcAwflC++kbrVIoBdxetntNbZi2zbysQzk7I9tQ8om9AsLpc4OD6z+TWd5r
tRGB4D1Q7iFUIYaA/J1SjED/+1RKyLgXSmnLD4SIXwogS2/nEEzuYMbuU0ZO7qkNVGuRSri9uAH9
IOn/1V4lwsbHqVzPJirlEykPQjV9/i33AfCOeH2RmmcxVoFM2luPO8wXCKk6BWy2+ZGDi2ky6Z3J
/gF3nmtN2MSwMkVMCPUDQxDTA5/ZdCLZWktAVlA5UjLlkMs8qmPu4i1OKLsE2d346kizSR5CGKy8
9JtzUhIuukAp9uWEfbWgNKy2L82ujFfPWR35Yi05ykvNf/1EF1mwPxmmVcJ2U2c2jZ+eu0lxcASM
w153kjHMJTYL21H/6pfNExoOJIscNiouBRjjgP6EnK5dKevNHlwWlzACg++RFzKwZrPMn2XF98yE
cKBrEe2sFmlbjZqmM3DXVXl+9TQJmKquw10qJyLvqTZ1MJ30Ru0VNNBqpzdTopI3qrK0EaCnfBrz
wVTL5IEfeVeGtfA5TIqhD+5VJ7cnOupYLU2zMd2kGytWdhci3UWWbRoVBS96OJZh5wTFFh11Yv2T
2QdrO51HbyRWsbz83HqdylvoI1gOv5qM15/aR8UnvfydDR9D+e+/AamAFXflU9hkJpI2O0+EaCVG
KUkeSMuX/8btq5/gpDl33EK4X03VZqgK8Tdlh1lVSAucm82Et27UA2ZGPcAJNruUMON8iOdFUV3Y
B9/nwVmkn0kL2Wq1lDrp3LmQu/8ufhmOCeKBQg5redavblLllpv5hpJ9gqkhowOOGcn6Er6Fq8+Z
olr0j+5pVZvSbfJ33vqY2SJXHePCqDQ2q8oqM6u9IH2vcIz3YOImRJqUy3vGN/pYoG6ai5+2GlHT
OWNdcJlFmwJvvSf8nbb31IHCi0uiFS8GWU164SybhAaD1ZPsQ/uasv6I7cT2lQbJ/vrXVMy4o/Jo
IxytoydFZm6GqgGtCLzsCaePDebS0oRr3HanZ0SJ2qvNqtfenDCHoyEal4gokNN2KrkVlGjKH79C
gdPfxypBNF20GxUzblTKRP+4JehuVDbCsLtCnZHPCYBjK1uC08hEd0bMUmAsKlEi0eDll8AsQBzP
vPXQFzjO2j3AfHwIuT5bt/ueBSw+PvMVcJFvnSw5zyTz6Xee3lZsd9GSpfCI2YEtpHEcbHvTkFzK
ZFcdyUaXZZc/ySQ0FuqDYMwQkGboU/inGWusUVOApc6xkEs3pz7Sn8qh72Ot5kZvk8xQirRy3Q75
mWYZj8Ufr0bFS2DUww96pFITy33BX3tw/BEvS/lC1jLrkiUMhiMjcCda4zHwn3moZwQZk+Fv3vMM
28yMp1F7BXiIaxfvlPICcaNvE7UvtWEnxWb6xcMONAlzPgJitBBIdGOy+TwRctpzP/g5AiRRCq6W
T/f0opjT3mBCnxCpnmIXH7QCh1mV9JQk4/9D/UvFqYVLgMC86U+qKuoJcFTzuqHZ5ftzLo1fm6gK
kmyZESjsgbyJC3zKpOlHUFHGQU9ifDol8CsTBVwxHPEVA0/hqvwunVpHFOKWR3jaaW/G5Is6VJVS
c6G3eRrsohOHa9Nd3YYwxdKH/s8EX9lR8mkDyC/x+bX5V/ani0qiLj0CrE3SQ10XNQZXi0bQWNba
e/DJkPuHyWNLyz+NViOZaDvlhEtr4DdJ50lNDMDEj7Dj4bTUNe6POZHEHEmN77AsSjwTWma7GbKM
dYfMF7c3/TznynFDhrEuc70tnovCOxGDtEOFXUGpYVZF33mBNgV6Mvhg+jBgoku/e6mxpKKU7Rxb
W8e1CwtFdtVCMdiiHAjVHovUWcTcdFYDgIM7mMa73rKm/QqKj2KRzE4c4XjmZrquggzJJwGA1CZj
esWNHZ6eXPZybkUtuNivtitpj2u8O64AwtWquzm5I0gnkTcVlzYV7zVLx86k5JECQm3zZ47gozqY
+x2rXrTCynv02lFMTs0WcAzfDasJk+nx+KA+oGQwX1pzB2+VzCGAtLGYrfiaAjsbwpao67i+JZke
3BXJyoZprLt/8NNK98+DWfdrJiIVOm+jNIL/K8YAJWp7VYgzrLt7WjOXvgQtijOTAllwbB2T8AeZ
/ZTkDZikwz0CerXnoWOIreEtmTUcMVLhyGV1Fe2llR6SGnb/+nqCdkmFaz/GkuKIXaC6dRLLZAxc
u5DUuvdjMyeREkuSt7NmHQxm3f9L6SDN3dhiXUjcWHSZ/67jeCKFMKwpYecsVCEpDGvMv/wyotyu
Apy7kL60cn/EZgGdly+Ys5YMh62c7Kfzn8eoh6hsDEjL/CcvlICtJffmZGyFJuECK7bhP9hwcGWZ
CP8CU/gmAMm3ltnA4Mlsa02K3i3fm8foEqi1yYPMHicoAUC0FBbBHuG7Mar6P5wwcj0zWNf2AGaD
5gvLukDJ1/1qRX/z7Mpx6qJQpH3n91fq41l5Y3krBV9aU0KRjC9uNMXjTAjAzpf6hCva5vqlA95y
1khemFJfnuNgqtawD4ZNdSX0qPk8ZoKYXtmHPWJ0c3dM5KndZcHkVkBpcpe4LIka9Q5HUeFVR2ml
Kg6+xE1SiGT3qMh63Y/rj2dnvPSumSZ4G/cZfs81U5d16t/elAZIj3yMc4Y8YLtAvjvOh7A6SrI7
/WobECsTVPLeyoG58R6Fls/PmQoAKuUjAa5iXkS9aayAaaqzmiXo2934HWNfuF8dnwF7hGQI0bpU
XjdtVGpgqfvgkvIKZn/l2fIRke591f7MvrEtQTlVlHe8gNt67kOnWVB2YdL1lmrZe1P+SNxDj+Jj
edJAyrDYsAkq9GU2qilvoqjtwW1WvVkSbzoHphvOKOBlsy9szqvQMgjazLhBbkqVQYT5iiF4hx0B
+bP05Jlsp98EKWUyU/BYm+aBLzOgTzRRTCgk4aHKYsk6D4Su8yUcCGMTxsoH0l5w2evKj9aK0pV6
BatxTtNZJ+fvbee+c6+u9Rtkg0PUTRw71VLogxK8XST1j8vgLgFki4P3l2AEsoLViByx7ZJGIXPf
WPqARVDpHNrHm+fVSRVwxzEKs1IROKXcz3NQl+Qgg6lKYRh5FAQoDpvoR+kOsWUeFskUrNGi/aBv
xKFj3GORLt6LoeucgzINfU3JblR1xcBDYNG+p5GK9JOkbox3lvv8kzWVkr488x3Ci4d1iT3NFykc
NLk8uSUtA9ZKTmKNiL8/wubaSkqWRdm9y5XMfxHYXvT8VjWHL/oen2F0juF+HUGASxLXR6MIadOh
Og27Hpi1cRYAryqu/otiY8wvxLSSm5OTedK1v9YZAMeVsQzjgy44b/fXfSqIeuiKTtQDpPi60BOh
RKz27boCwH3XVO+amKUNPXN0/jVbMzTM5OiH+LN59sdqY1x7VDRA1OMQKx2vVDxzHgdVr8EBE1o9
VseQK0dTxqiw4tUpl1ifDNBJ1RGgOefMMeRo7uLzYAGDk+FjlRQEzFVC0wwuC9iF/t9kSx+tVcU2
F3ImIFqY0Cb7zdqvmkQv64+rHtipBtxfzyx3WsdpS6bAouYLAgkmoe8UYF2/zcyjJpdAXPqT4Qec
0pE12qNklz2tsT4eY0JFnAWbdOkkT/ArmwTQSh8twwq1YZKR8s073XScWGno549iviBIQIo8sSYQ
qzJ2I7oJMf4bqljEdptHdJUohVmrG2J4/TtH87nH9XxAFqG5r1A/jEi4bYD4KfUAwo8U/MZscpJw
P8RELhOjkRgPMcx8iKRKs+Qa6ggdqgoWQwt9YwnWWeo7jkyhReHT0F7rIPcn4vgO0pMEijTJsuu9
FSfhXI/5q1lKrYq6V1z9GvLXhYAX8PHzFdUmQs27d3nVw5268V55L84cRcNDQRoQXrKNN1oMDzNs
5qkQHTs5ZQmbGAcwtuOMlJu6pZfV0dCJd2wcEPEnWK2y1/cFUsgIJFhXPOgu2y97/kepSlAvD2PN
SypgEpj6XZm1ZNTRArAjVmXNrtDjUp4O6Z8bd2gHY3+Ap0BkeQAfnup4BYVbjMkgBpED1Gqnn3KR
K2A5g8fDhmAPMFpcWakWQZZDukzPnbLSq2sweI08jmCL6MKgsrWvOpsU8uw0n8IkhX8VeQPN5L6/
ok8bAK/l1mHZ5hY8UEJZNE3myWme13L3hLn10jO0JjQqABGZQ9M3WV/4WN4SteRhcofBHlAeccDE
sKbjWbMohAT/UQcL7cgNryd0Lh7R8+tdlVSWZkb7CKffH4PU3AqQCPcadUf+VF3OzyryCmClkjkt
b3nqRqq/tGy4WzMo7BNJTwijPWTeEzsJCaqlzxmrygkkM4yOTkPWStln2jKTuERneFiQV9W4ZzBO
sOMWk+Pd9DnuCfY0qfjTM3X5V8BKZzVW4kfp0ZD4U+00if4Pl7XcHy3V07aR1SFE4YwYc81Zbxyh
ZAjmZO384D6MC7NbxrQjYdvXrGUv4aZNtrVHASF+qWOS0EIR/DnmSZ0nD7c/rmR2L9psnOq7q0X6
Bi4gkbcEpASv4NWUSM4Ds9inJ0MJ3FrxGXmTNP159Y8dtJvyfJBNfSc9mAfrF26k4rdbNmCN1keH
S7/vr9NCaqOfu/px24u/a4BNTdqbdyLegti0BWycmgjE/jntPgupZR0U1vbJuJpwULpOwgEWmY42
HqhXDPsZ2ZVqqYS8TRDsOXcA9eemLNwY8wLES/wqh+mamzAEgTWsexiqIRbBfYVURsarABzx9YjY
B4j9BK6pgF9qU93a5GhzjAOghkV5kxBdICEsWF0Btu2U1saXcknuqgibVDN+xmAK/Gp7o+/0L9tX
yAyfIefmYdixA2COOC9BHeFHnBQ5MCam3d1pl08Vpzrekxf/E+8y5eHE2bPVmBCA5GsPia72snN6
rCfbPKCob1H3Szd2qKVJqvPhKK9oHNZ0S4tMtiIpM0eOzI7pQdGc8zleY8dvAfP6k1SKPmyA5lPb
ilZBs8bXe93hazIJRox8K6jgrjovlp7ubymDgaZHgRaLozbWKzVkQGdA2jt/b+Wd2oHdYDL1CsPi
iLuXDl9a/PwBm+qbJ2PspMQdSo9zXEaDEi/N3R499iQVVaA+yX+ToT7h/uIgSzj6pRW8L5r//dI2
ZuxDgjKNf4leBT7A4Q1dx60br84L94SDvLuc91We57Q76bIt7BDIA2LafGDRTKLto6dt0BDn/KpF
hb9oCstHkqkP9IUm3gewGtC1k6leTKQeyu7TKxhvZu8unIEmjp3lPtfrvsuh/z+XaR9fRfIAq4c0
6r9zXpRjtgIogf7OVgsQpUijFQ9z0El4oqcKYhyOsxlTk1AU1aM8HH7GnwU1t1iw47uGKzLnuKMK
TcziyE3ARi21vJ0fQoFGT6a+uv8pIQ99n7D3iPgGmCDKDYVrBRvnJ7giUgDTZFZD+jqRdbzqOvNm
yhZ4vZV4iOor9l1in8AEC8UAHcojM3muhyLB6F8VGR7Ffc9Xk3tNFUJc+vlrmZF4iGhVlWOjGyzK
y5zM6hQr+At+k6KUUlDu0nXoSwW64qtLtfzVcCmsbzPAE4gC49PbqN5OckxF8s/t55LoY9a/JWDY
brumc+EN6CeLmzLkO20aQhPcHT8HJF11KellmdvK/bk8CpREWxwCZvgSG+Jowu34tLnMoFQTfB1P
5+i5jsNaIs+gIIFJHbYLg+xCk6ILuNwoDtt6JmMNa+XZVM9Amne46104CoJrZdWEb7Tgqr02WP17
M6u1pKFdJ6Ovjhpiwl9Zdfo3rIUxFNerntXmxT3YikCaufw8XCYJWhniZ3MBoiDdluNYUjuLiOBD
voqdA3n02NOYaBk3RengsgB4T5dc0xxaHVb3TW0MhPmexXNhNmlZzb6lEf7QQvlfNI7KxTZiWrfq
LExKwRVV+POIhoY6M4ti20WUFi6qCuuq/6Mgn1IXOJlmmVGGzZFDsm19KgkXUPWU5/Zi1oRsIvpP
Cto2ZsicvCgbDg4WuPlu7u+W5VbgHSOnKJeeN5yAfEr5yqNkAIYtwLVJXvtoEkwwTrf23ge0ta8F
r9l5NUKSGiv3qSvdWd7Izzp16GE9s2E73/1lZF/NXsOAf0vz1YYauhZ6+OIzVWVBRmwpJf5FU7sm
S5LixxHohS+6spJGoj6DsxFMUIh2GHglKX3HR3NJgO9Tvv+OiycSgZVZdJ2l3Vl3LGCILO3JQVuC
EKjK1UA1DNp0MvhQ2WoAyMDkf4wBDKFzcmJQRFRNHXgCY+wJWH7hqnUZwjZ9CFNp2CTcvZwKOLKN
UXYxRWdRnFIXRn40ak2t/Jds1LT99Sf4d9ofkIPheL4dCLHYlUnuBea4WXA6RYHw2FPQ+V+YXUJ6
RFb+ofHRv6soR4rB+aqZ06+835/KiEtxT5Ur2j3lepY3ldpeSm2fbIrFsivR3O576qZIpaGOvCYC
wguH77nwXvbzHEayamP56Vjs1zbf0kntwq8P8VfUiDrN7jcqPbWvxpQ3qlKmSjrB1zmM2G8Mgtib
KbcxaO0IjJunGg5jkbUyn+T6CrkOX9juHCsD3RVwLy1BwuEG0W2ABynyR2GtN0lqvHe0j8SMb+AX
jgn17EJRtj7pF+SxTzExXJ7mbHTl3QHotB1bnXJQbLoepg9myjGzXN1PdEFuHwGDz1Khn3xbjkbg
riV1nFhrZO0lNO+CpRWg4f99tDXiP2KmSEgLj1+JXirrcEcuIQczLDtlBAvjSI1gfkkmwyw5uZaY
4lzpMuTuLuOBaNJnOM/6JN0qeDTb05cTKC6wycETJDxN72SsyvTwdNRviWa8HAoze00p5WBuHjx2
aanAM0yet/nAuDnma7aWwMr6hInnSR/tzPd7L23iULuQxwYXTzWatYVKtjB+R6FouYdzkQdrMX08
+nO0wAcX26BCYA0N7bQHYmH6VjSL1ggRxAbR8q0s4sOKFD09ISwiVLKn6fbr5dKYSZAGSq+LYd0l
kiBhOAxOdSkRXft4YxA38Cl9lAfD7Dhgb/eQ288iK5yiqBTYlyNjoruUnaeJEIhLFkRG2wQ+eMEZ
zZNaRJGcYYGFou2Lrn3qaD+OgMaVonMXGQIJaMopAv93olFcPOiysgmSSUF5e8WHMfv/27FuiWS2
bF8Lk+jnolsgCJtD7/VGQgCmOz5VmKROi97ANvB6c1uq3UixdxwF238KVb5xtqu+keNFh6vbzOpv
f4IwOY5D8C5JtDBstwoWojnk6RGUHro3r1MuL8EnRmyO/wgtuugCzZOYEQljf/wg1Q7WpZtYkJ4U
yeCYA+4BQ8svnP7Pgp65OejcUv3dLpCmydEQXNu0VStA1ILo6m7aiQhC99xnlsLuS1dPf4/L2VHq
YXikAR2WIVCRtnZQGwrYChPIK2V5lDjkPgLqa/h/ce4dqQ9WowdmIhoNaa+s5LNJxkziIQXhtsdL
prB/SN1ICxy2/83zr0h6nP9f2KOUeBX57sRi7aPf78nC/XVD+HWHJisnFUTS349VO0R3tV3OgXu5
9TkUeSyFG/Qh95QQIjKaOkwwvruOnrPaCggJ2fNCWJJEl2COGtAKCL0chJfKL5hfH0w124u4FfkS
H3xZDf6fbVUDHn/BUU8/EgrxeCw8/npqzXY0FxJu8CUCQGtaN3McxEvRTdUx3+Qhn813VaGGrdHp
i/StQOAW61eKLkl4zehHO1eMT6WT6MIyLrz0PWyUWgFQMfYtcdqEHKoLQaORyc4t4FC1sJBQI+t3
Hn5qNCFL9pZexyPQ1R+o/QJlQWvuKDi78hwcGKXQashKoZ5Fjjfo5Jp/J4KstHYMjzArBU4680r6
mFGik6zvhtHvkm/ms0PKkH4xwoIs6p2ZZJ53qhbYZJ0dXpioR+vTvg27x/A/7tFC356Vk1pc3J/a
woOwuKoq8JgfUeoCZ7vrFeKsrrRLCd0xFQTd4gENeoSa8VRcgSfILz/DE+KpCpYFZqdkVUx2yczO
43ne8E73WgDv3hawb6EZDZ8s1kGgv2ldtGzPrW9m8k+gjXcj+fV+jZw1lmzbs62PUJtsx5WBqTk0
YI+1jAUyUW87i7+u9VgJsCTgIsvCMLzGCB4DPSe9UqseYRsc1PtiaCm/dSBUXZ6mWD2/RYbnA537
KQ7nq2/tivD/5+0eFRv9IgnGKyMMmJjJZW0u1B5wTJrCwWwvPR53W9IsVGMvCsmY2ktsKjngjE+q
uZzalSbnRYAkGThNtlUDOQTPg5eKVuV/ybCYSeX2dYQ0b2749vyvmvyuHn7xFMcqdke763nqA9Y9
hqHtCQVtQ3blNucMYp+0+evQ5FH+AHLoGKW7wIzPMJB1He4/nxEGKUL6JQHBd6YljoYfwL3sDuCo
Jn5U9XNMgUV5lbtaZC64PebdXa8fiI9EP0/bHTyRQbWoNJs9ZxuKNKYdni4xtID+FiMZ4/P63SPa
PlBrTOLh+PELoEqbK8Ib7si42RWUvicpRJZ9I4YxjZrvFh7gS+Q2UmyGog7aQ69uFU92+qZtaQ2h
nL+NA1hjwV+o3utVBdMLON1tmIhi2aFCtMRr3XqgL6MUfS2G9HW+46h69sw1L5Eo3MDO31w5ozDT
x4zvHDq5vz8Fz5nlz3EvbztyOqSBJtGMrD+bpBgL0gTDj5SMOn5GtXTqiobtyorBDdMioWfSWkC0
+ii9lyVOVTJq9pbA2/JsOn3mcpFU913cG90YNH9XALV2TTF/4Wp0A5zTAW6jADNOf/kRqMDSemVM
iL+dAGYs/QoyMdJ0BH87cRpEao8INh4XyCT9ScfQYX1T93XGatneLoXga0yNKW+D4/65eEpDCiUi
DMhxCgwRzvC5mm/zaPje1waeeeu4wDND1tF7qLmF7rMxWbw52Hfw1XgXmjsbbPQ7Q4IyCnP4O26o
xtHwl7DJNuzyFqzyiO5fjTpvDmjo9lMatm503xZZA6O0QdgrR1IdpYHIewbqMw2SlRmXe62jo7Av
SXNKY/X9rO2p/clukoOfpZre4yfs8yIYBJiUsD/ozqA18OvWQNRCbf3KbrlDlRl+SFPOEJV4ReiE
SEOvv0+OPtff0syb07WdEGhvGCyPPWhTfufpjS5GFwK43No3Xv0mP9dHVKc4z2MnXyB2DYP6cxx8
/TX23mppamxoEzDH6ZwU4FZHMWvh7dcc/rVR8O4938eKnmigjs3ipk2dWnNEx07oopYUPZ+H6T0W
sXsicpB15nzDYPirBfDhMEXnF95t0tLk51qaeTBLkvC1fVY+vgLwK0tzrtIFSzeBy10dAWf78Nnn
15QB+/ARBUHvHhpStPOk3lzEkUipBWYvoHZcF7uylOG6Wb5uhHbkEdhhslMg0T1ZHDARxmQ5O2Of
RIvefsfKIkP09PBgAg+h/lKDe2EMXP+yVVCjCcUUg4P3oTTpY+55PvtrYLxjwMCTtLGhJOcdFluo
9pTpa9uR2HSYHXxLQvGY2AGPIqt/D+VI4qCNLKkK9N3qXcnI4NiRtNb6mVnj48oZxL3fiPwXPNZL
7XFIP3rrBkFwfDb5kuBYr6mvM1a+oTp8weNmus2+VOGL+7AePRULHn2tyPrnLYX/WEVV2SldVN+A
3Mp9DHrn0cFcqqrADMTqchen0VgiJm4aGMfa5wHWY/RzbP9bRP4k/wi1DfO9j1JmL22KnIAbCM+K
yPnHdz9BxwNZqMMZNYh2Yuot4hHCxY1rDlDdvTjDwBkhGuE8Cc9rbe5HpfW+/xe7BblbNHpF4qAa
hW6uvHHG89T6KOn1TxkQYXASUFSojsC+LlB/4uOJYCntrJ71lxoyJaNqE6QbunfCHQEj3FfaHVB9
PNa7RsH2v0mj6g+9m5W0v4/pOQOyjF/1k2xBO1e/0JNZ8BpfGAHvW8TquhHAraWGzkvSBMwWsahH
u+Ggs5tNr0d2hgn+aaQsdicUkPRceH9CF7B+7gReDnnkwxLRpHdjq0yEfueO4PiTjyxVo3aFXjzu
5Hk8scviANlMys1Q1NAlE3NfS4fDfKy2RuaCfKPppPx3KhMi6TN0R9WfM3URqFhW2jtwX1yfwTXT
jeSZwMkLPxKMIkip4rfAMlTOttlVBhPOa0PttXbQULa3ncCLRs9zPf5+SPiSIwtivED9L69P0Bsv
Q15NrauB+x/8Bot40lp2UQvLzK9bYuMNwQ+56SECNqW8RnNYGzK8n8aMixaahIA+pmvlC3VALfjJ
/DNlXHO431rApCUOWVilkBimqeYzcgyab1Ze7Uuualtf2MNPE7vpGhlQ+nL9EtjcFFiQx4mveRLp
fMGwIF1nwXY6pLkSg9lHVbPGvzzPJfphgAZty6oPeZ9OsVdgwilftJJGww6LSaTjDfWecLz6Y4OW
qd/Yo5oavPupO9RA7UBMTpEV4U9IZxz+OuT2H5SwNrOzkP1MR9sqZbWK3RVsrD8gtgV0Kb2pHKO6
lhLa4+kVIZIde997Q1SbxhKDvaI19XS7xtLOSVd7rki4xiHrCuOJCjatU+EUmOWW9uT/heAS0ZQ3
2efAV4KJJFwiH0rh7dZ7n2eerMi8igSHGl4DBvzF85YvPnXEyTOtWgd0psg9XDnflr+3O1TmM4NK
bFewnMEXXMV90M1Jzpt84WjuTdmffNmWl8QIG18rh4IhwzWWsCLBayQKzMcdVqWHTbDbUA3K6M6b
/oKGyBzvXJjyWJymYkP0QxVlPZsSQlzA8lKP5Opx7hl2br96lMWzi66HLCZDKAS3x+tiJz/3m7dj
uRQkOJ04oFmNHxvJCYNAgikwZfNSF1FbZ5Pug0HACiFs8V2XlXvHfYN3KC4vgSwQ3iOvLYDC+Zhb
Bn+lG3s6TqZMhFbU0yiTEn2DLl1PboE8Q2CgF+mpCJW5+6MxEqF1dV8D06JK8/qUhGwsbxjL6pn2
C4ReBR78lxxcKK91NilGff08gk8d5gJR1FX9TcoDHtFNtgmACDjEdAyvk+nUdr2tTWjXnxlhqMSV
LR6ysuLg5pqjS9h/9dAzXsQtjEMfW7eJkcj8hHYmIlfgixv1JQuKJRbqA2tJbc7og4SlJV+7Viis
FjP9WGM6He54vDc5rieHx74DT8fV3iKDycCbjg8jnFD7vyceXbMuWYwaQphw4d0dFHhc/eDXHCM2
nyja/b6T/np/CI5pRFCvwXClq2woBXwkD70c986E8qoN/DCWqERSPcqsYJRu/sWEBrpzrLOz8fpR
hUgyszV3AG920td2FF+rsYK/zTjBtPF4CsYCOBD635czGXZ7tY4ASgAnp9v8c5xSrhqOwqBIPROE
nOJ3MdhbjVShAQUqyP/HdIleS0Kvg4QVk8PfBe9jbeLtphTl9zWOj6NxSngAkCiElGsl5pNC4aeH
4mSPdhQWTNx1jTpUIUXsJHqfzJeNazbGLER3zoGVvzwqD6Gzw0U5Qy3jdzyzz9xMmzvLziawpFBq
lOQSQ/gWEWrnycqD8Icn3w2GW+Ww6oQ2FIL6RSwQZcv9CJ4BeLJkmzH/C0Ym+VK0y43onsQKCK8Q
MTjYTAf3q+DAevvUqicDL40LgGcr2wKBO2+oRZk5db0mXOkqI2YQsfurAgF5X1woKa4q/JC5tj1M
RI2eTcsYH3GEjFt+r1KJ+Kk03lTkWTJ+d2vK5j6v8wfjc6FYUOLCT1NszGWN2kCTl2vfLA6OkY0y
fegpq3i/T8cH0pCQc82x2qexVeqs2rhXJ4rG2jA6SlKdYMmaG0BTnrawueIN4CM1Vj7C9R2Ka844
q0duKXuzuv2y6Ohk0nDm6bBB+r9/gMKTBGg40xzXkjib7MNGpaLybl1UQiWIOdo9ghgvIXjvHEhp
RdtKdVkZ6hLkIYw8eULEGBOxJX0pKndeSCovxNlsqvfDUxLaiuezn1ZuUoZTdYGKHPezAROcjml/
+YbVHwgzIpACREuo+6JiNqZQ0zrbD3ACQzEHCfjCD8AxlTQXB3E8i5Q7fLWFGapolvi0HPXbezow
GhOvt9HX+pqO0Dud0XTScy/ThkysYVcjuJzdhLUitW9RhhuRHhbX3CaEOvqaLrzQJ8y0v6i2Tzkx
w1tA4aL5+QBRyTFcNSHPHSb5dMexuDY8PbtMpKUfmCZYcj+Gaz779Cs0AVwWpmwAnqP6mLR0NY6I
0A7OO80p7rZvPeK83jaYK0ycmYfSPFdlycNILl7twxSkpWEdnihxzTWbCdElGZq6c/cpyENPVLVj
V727ax1WmK4uv3PiiX6774t3iMv3Z4VUkKH7b5wndTe8/qsmsa7YIno/Trq2cI31/Cl2PmCgfXro
C1IvAaVkhR42Cdwm/y2Eg/woaxkHHYsbT8oM/PXSFHt83FX2YL06n4VpzWDT7NdhemSEQWiLGIh9
QolYFpr+wncyyTlxPfuMKhz5KV0Cok3ItK+tSjOB67FOeUEKRZ6Tp19Pr7CF2ZuyuuHFgmdvU26T
hpc2sL4v8YIBd/4keh0kLZOq3yali0YDthv3Uv97f+GAxD+jL4JSwypGSHlHxkhSjHjTUIyaypw/
yPy1OHkB6FLQwHa6nvTfBmFIt3tJIxxW4uZeCGshzNjGHUvpa7/ezjhEdUVlVmqlvD2n865avp9G
Mu9Yp5tCqe0LimQ7qji3iYGbE9vZojpxu5vbv7fmQekpqcY3BBUkS1ONnRivZEX7xIP8rZfPqHuk
vA4/ZZWHah+C+XTBE3P2aIWuCVkDka/BhZcS7N5HJ0HrieWNeX+U1+mnMQL4snK5r2t/n+CyolKa
iWcyw3O1BHTdFXBR5LsR3nG/bkODvM2XIhWre4HRqTRyn216TeJG384C9z54itZe8RfobNjXyv8n
rok5l8P5IJ74kRPBC6kAvLeD8aANm0qOdynTBKpBmonnkJW2WJQfFydZesOimXXdqtK6GxigXTvW
Uy72k0S5Gj1RGdRuZDISY9MVBjHPqUplpSQp+6X4+quUzd6kdUr/jKyf5ZiiRtyeCB7H2IgVo8Ip
RP5ZVBhiXYIWEG3ktz5zD/VlSPeu7ISfBICs81C+bUtr6eJB+J3KrhXQgWxuXJtCmE0KGRP56nN9
A9DLrb9dHPi2sgdB7bpzBBXBZACR1b70k6Q+rvzIjQRSim4YV6bGivDOGpkMbI/0m7auSybDbpCX
KGn2WVobhwHC+MdU7ZQ/dACSv5tRvA/4aB62DreMClkdHoIrRmlLGEAXym7O2coVZ1ojnM8c+sMp
1tI1QpX+RHX8l+sLTNqNp5IZq3JnfS+KYRfn80BXOprGV+iwS4ibtReOKnyXxUEQHszm2zhp5CLS
GOjJS2DbuXquVMuwsh+Dqe45W795Syz68JLBIjml9BrN9zaKzgJ52ezYrx/hEV6K8z0cVbJDw5d4
yab1BqqT7CcqKnZec3dxXS3UmBBAbT3kgzH8e8J1kj7ZTvIvJdB++JwKAIp9Ih6FmAi6YjT+OD0f
OvgPUmMlHKi1jBAFJZ0et5XjMAuPNNjIGz0ecF8aoGjZ+mjqCyQ4WmjGvK4V2eSiMjUw00zWo/AE
fwyYOJg92yYKa+0WEpnlv+ZCi7Npk2dysPtYXC01pOLAXGbgwvkSPVg4uMjP1wKQLyX7/HK4UBB9
OoQyMGMOOwjwuhh913ULEug3OMVHp0gF2Th+8MQfHwFx8zYvtWURVVGtePv3tIcSp74fK0kyeII5
TBMe3bkonaTWEqK0t3SzjPolornph7C4D3SmU0QGuzGFWhlzjA6YCSb2g3tRwlG2A/Oup8Nqt0rh
m+P241Zt6lJJI58F9NAK6Pc11iO05lR23AAB/k0M0CYbMvjYbVbojWxqNKjZZ+1xZxZfYJGHoR4Z
X3a64BaIoV0sFexgW+Q+Sayu75MZT7lOrE2k63DN0xj68HnG73rL1oegDf7pH9zKBUnDGVZizqp9
EZwfCK8pnhwAi1FMeFj1XcdCj+O6ZGC73YHpLPzCWOnIQ0EdFw7cxDsgDpKzOWcHCHWAaQLaJTiQ
XGVVjp7tEbJlxFiZrrfe1Gy2mHH8mTISvEZifi3dls5vhuZ8aCIy4NgcTEmKXW6iXMbEk29hWLIW
OYBhYGA8RDOCcqBxB4DzCT88ZP3mUIEgVtG9RoDa9ugLW1spwwhBb+5eAmOZjrtsZxNeluZOrRJR
XD+XcTn7wOA2O3Xy4ZDGjaLMwymrUNk8Wi2IFEGCTyFCP97X/Fq84Hs72a70ogmLaZEWjBgQ1Dug
L/HWpYZtqljMmi3tSFK2iN3GgVHcz+ImYVkzPnF2p1WubVgMtE2g5KM38OClQamvU9v+SRUWpHjo
5I2CwP/zMyCOQCnZ1Gg7Q+/g5EiFiO2QwHZyWRyzIIeUbkjHR/P0vjvYILI+45m5tHmShJJ8ggl+
Gh6gYnA8AAHmkfox5r975bn3omYCZ7rx76hYm3c20Z+fvNmgIEsFCWTYzZZZx5cuixMfZmFpaOVU
MKt+B1LxNMUb1v6AOOQ5PSGWpCcNUTqwUYBnfJDlCPoPhRaGD7wpLoQonKw5R3fgHykjukVcy1yk
YYB6JmRji4F4K262ic4zSXv2kFyCnPflqsvWZZcxyPvNx+mcNP+D+9dViy/ozZwiuWd+TUaFobHM
iQaY6Z62jmUTR+0cstsK7DRe6yIKNDB2krYwaN/wmtYmVlGa14veI0AEp7bQhjAk5f76+H81/3Ri
ZcG9GAjafmfRJlTAP/L0VyT5KsIpZIhd4dKJ7klqlffFebQVuCDcHWngTkt+WkPx8a4YK/FeJ3mP
KZ08ui0n9c9khhOA+BTYIOevjvE/1iA9irxYxttWwMaOF8Nqf9c7MIB1IYSLMi7Oza4TURWzpZ4h
b5T5PTvATYILfGqc8KDSL3dHuXnqIxzLH0AYa5B//Ig6T3NQr/aTf1BuJkGxPESbDkHVqYVS5Acs
lWSktZz+gJVLYKktCxPhzY0efBukS/amRh7sW5Adcxb+wIN3Ajm6Z2dmWtV8eTBazo4vjXi+qrqB
sUcMJ+89J3NmHbjHipuk0g4pt8gctkTUeamP8ukCo05ec/aWTyBuIb6+FleRRZD3yFaBkJxwGtR4
KnsMjx1gNVEqC32itSJOL+HgwYkK5D0hFO/elR6e7eVKCRH5j4O3EkJTKkhJEYxP8CJJm/akTvxN
gaG2KPbS2zITmKadRKHI/GyHP1HSOflLntwMD88b9zVtm9hqp9YE4t/u2Hj65hUXnIEZ3r8ebgO/
dJV9/RbHY8oSoA6H2U0jZHwy1QisIUcUbJgtGROKTs0rqAe26HCldP+/oOefEb+0HN28GBlpdjfZ
QGYBC1IRGuUaKkNp+40Mg5oHbLWm8NrLiyog1smxEoGnIzvePK4EAPn8PMSZrMjpudGh9naoWqoO
2+N891k7Ud2/xRr5Wk85FsdevDWIZnu9aLONGIQRBMiPbmRgkJWkp7/VjzVu149j8T74kcqszKbU
SREt+JkvAGmt+xUtHHwYE72+nZsqkpBjOuQ6MAg+POkx8lWOFGV7H+WwEFtpTtr23l8OKLlEw541
/HRPnNO1rd8YEtA7ULz4Sa+c4kOwRyyM2/tg+VPK1XUe2l3SmPniOEgRSM+p8svZt9UQVzbPje7n
9KPJWNkXhrMQ2wHPuAauK/3HQZounxWV5ISrXt3w5McrzVZwiTzYh4A0Xaw1UVHHak01M+i/1mI8
abeoyqrMuRYImc87iztsi+uU4VDLVlp7uz08lgASNlHPGx9vwprzA7p8rg/xmnDRn3Bxa1wVDuw2
4DAqFh1kLzO1uXJsaEp9V45KFFRPba9MsEMLc0LXqOcS5TjYyYd3uuw5cwgXG2qTpyVNDOQNCOZm
jtNDfjwpaqUPH7CXj8I4S1cyNZ+u3JMz7oW33gm/DHxeZAZ3Oqkjk5FtX/dqI+4a25BIqbv0IzrA
3U/Sgv0C6ZJTOBVpI4ZpSDSg7LZMcf42400a41aVgla9PdtS1r9xfesDUQmwSUs7mDG7ghL9u3wQ
2Lmn7rkUsYvLduc+kYO80A/gggFJKxKeQ8fGm9eJOF7B42pyAfgvMraWcFOsDliG6qNO538DL4Mp
Lxu4WjOOC2R7vBBYMyPLLYNxX9LTu+C8SOSBxKkZPjAfSo7HXXw6XWqpVb9f9RyxpcPhET05MR8p
ToGghujoY7Zgb2jJvRgjXMxcaBdomG57QjOlOwGhSpFVXwT35nq+/HMjPEBrymVdXwYcsP8WKEkE
2OmLibxZTqAgEcIeiuNH2nUF5ci2jubc6DdU1alliOFsi2u41tB61kC/4rW/Lu8OU5C8uBAtb3vD
DjnPMGRrQwHERFc7w2N8Ej1CZUcLiLRuQwwkvZVHJK43s5FKTEyJde7MUn4Y2egg//kxUEdzIuEq
G6FYlsX50shVrvaho7EHaU8OtlZ+vv4B+LwuPlTBefZBku9PPzHRQCkzr8MNTXYQuJJjQj1vQpF7
WSulToP0Y3Le+9nl9V2rt9nglNeYGxHP3hDvaiiJdAFik41os36YHs/KoSVgAWQA6p2KQNPymKay
mnuMr7Ukr0xZXzE6z9phuB8YYttcdRV8KSC/DtbY59Wp6JwBRZ/ru+TCyVsZ+7eVMMve8xpW5mn+
OeQekZzQP78Qq+J1hODS1GVTJ1cAAJJAwVHo3vD8cyWKAY354aC0XkbKNbyHIXPIJtOyRQQKCvu/
zQGbmdqhL3SZPIT+y/arqtqEqyePz4NTKiKeUyYqirn6eU0VkxPUpgNJA0uPDEr6PnZaLhXd1EOy
6eMSAGlsF31Q039sbEiMmwPsdudd2+YPRamAPiazt27IpNnVHvlLrqcBrR/2OXljCsmbBxRY5+DS
CPRoqY2Id00Sy/luWbzPpNlK5R+jyq4JI2LVzA1hje6B2YaNQfruSfCXO9800QVhAf2XZMwOdiMY
4FWftJZBqdwKBo7EJcJ1vRYGsBVN4mDD5sZfRDiNJh8BvV1YHXfdh7wneAqPl4wpRpKi+dCuhhKl
YnjDjuS9RtUqaafIfPEreuGGuSTWWCCvzohAABy82NFQUNh881sYSDOfiMxEtaYpZEKu/R/sq6/n
EMubJdb+ueRgfT78zBpJgBQsEdMaGW3m+dZbIeywmkP8X4P/widiJeyqY1IRUHVeNRhPqk9xCVVY
9crSP2qHk1mCajnrTlk7yJs6gyctlRbO+A2Hf5wMUZMBZGcfxCMNrPcjIIfZXJblwHm7PutWfbCU
DPZxUuaWGbbO+WDdXcyJlqq0SnhqKKMl03sv1Xqs5VUEPwzVT8bOJXpVtugjIJe7m2oWdQdyr8pT
yXgDCNLuQ93cH2vJOSSpHpFqkjQMBhN9H3scVjLdBYWlIGRzMaMTol2CyFJWQVx38Xm+7WDMfqoh
EpjZ70MTIkWEPENd/JQY9Qd4O0dbIPQ74ONI+WDfJE+PpZ30C4HfNpXthsStVBheWRB+aD+10HAx
6CD3OxVO2ICL3LSbIXpPO0qxv95S1486/JM61gizO7FLMtZAOgVFfz/ORXhIRVQfP+VrGFSx82bC
s2ntTO/g5WAeRdC113iZK5nPyrF1Ay4CUIflJ5YUK8IdGnpRLCaKD6PGsoqcq6xfjJJoB7TCUibu
3j3cJ6sOgj2Ms+yI4GF7i4wZyaM4SlQulNJSPHaeMuvpi6uz2djPBHyuX60gH1a/LA90oCQf00TI
0yhUYw8XruiRn8f4aQuScKbuJAWWwv40GqEzW+gETniMNlHWvFG8j8x3qNcqX6qgefLrmxM6cBUo
Dkdxp/r9ye5MchgelzRCR4rEtuiALEiXHFLlzxcA+Htvm3TfMLefQ2xS4724gMBFqXq1Y0vW40C6
Yn57a6utpG45XQ0V6n3j4UUm0NUd3S5Xw9QLIZISA468o2QkqvhjbwFtbvkheGlbwr2wsRwvDg48
3Js3omr3G0LvMYf1URZyiJOTJ42jIc3o76HfSUjYAlvn0l4oIal+lvVvfQWX6wN0ubyg5Wr8h9+d
bN24ceW0nM4CJ6JbiJqCkABNSBspKLVe4Maz+0+9C1Cs5W54rsziez6h7mLlCnyF1jOKjor8FdkY
S6KyB/u5B3JUMJsbgI7ZvA4BF8JzFzWz6Aqx4alDCavtsiQqtUvn7hpb+qhwc2JC6rkZJIA9OeYW
6WyX0zzY+/5RO/HVJXeCxatnaKEDqGKT/rSswKqYcg+k8i4+4ZR7vm6pj4TR6ozfJKSOeMHQ1p/b
ZeA2yBSGm/joo3WLoLYZskMUuO5ND4JT5UIMywWeD5wxS0aSMr9zmy4fQ0OVm2hwoVaZnYO+8iWe
CyVsQl7mFyQ2EHWHBMfciSK3VlmAhrDF1tj+5ALgungu+zZNm1NCGmkg8Ulm4Qck7YMb/0HSdsFD
rDUVQfT/2S9jy72w8CuTuN8II/pH41msvwOqnnKGkSCEpseTXjnZMivex8ilMOalTsqyP6inC8L3
sxcGhQP7Yv4NdRKm/fxxzVUtTJ35E66WL1msqn9bnkSXDADJ72Uo1EUwZikFh+cxmHUjCU75fUdD
L4EMwwx7NBAN280MaA3pvDSd1REyWnD7JOXkaQmxTNYqieJqRSIdQwe++9IDB50lLAXD0lWVSMQN
JeG8uqwakO4xU9CfUH8XKECWTHSvRwD1yiXttYlPqSrBtNYpsYGMy4Nr4N4dKUCQANZlIVgcSrg4
6hqrL+QeH7BXZNCPQdHB4mgIeajFj2QC/jNAidr4DeqezOfE8S6VPkDg8cbf2DFEkxFApa7OFOKI
bs+Tpg5h8Bi6+ZP8Qe7qKW9w9ZNaKioOsTzKYruwAQeR+lTOi2YdkWUXGrkGwRZHJUBZ3JCtTI6B
1JYOD+Vn7LeuLS2XHQZYksx/fBolbalryFY7cp32YgkiJvA0rvJv+X8Ka982IV+N5di80YauF3ou
YfLVngkTHqn371iBIORmY14kDviDCYcd4Lvd2/zCq6eVKh6QHsBckeQ1lVF73lnKwMJ64qMfLB91
COx6RVuKNMm1dglb74L3VJX1y7oQRg5G5ul331uhkUnhhDa031rvHrNDB+XdG0HEosbnTaEuRwn4
eZfi85aXEdOZKHLBgp/y3ZIn8CIJ9dVLOpIsBYEDP9XO4CO7CG9YCObgg237OgJjGPOioEkhIQp2
7bYy8oK5t+Z6wCjCq/Mh77jqJEumeeyooRTjGijFKvDfZz8NTfg23AD3Bf82MwX3OeJylvMdHaaB
p34SnQaxJwoWHFvPhJ4rcbcIIc9M5CWAYCN3JzRI8MBmbx2nfprJB4EZ/ofaqGKMCjFJ2FCnYVFI
Nu921UlJgjcfiEJz7tD0zjDsD8eGxhwQEcCPJYHcpYm+yfd+OdcSKziDeFtqiQVpvpwdPgRmLLKD
h8CC/xttz3/+VIXCNNwGdJhHsSzEBvbj1LwU1SXaH3VxOyRCNyqYWHFRk5lNWxGpFiMsRch90IJZ
OE7WaZykE21RfGcrgb42iXdXh2iwME7mYMZSFF2/c10GvPqxMd6ALc3R7FaTgH2PD5QVlYK/uX3Q
Iqc9OAucU7gxPqL6Nw4O4PfxAIwwCgpg1baEztmT4oXrKE/w/hUe0t2u6bLYh6yr5kKOpYYxKEeC
sNlQ0BK6VNNIATastoI2uazjf33etLuLECpIGY7v7QEDoi+4teQ/BWcPqTAbteM+ru387MOogsgO
2cmAxNpMHURkIvyvCg3S26P7JZFRgoZVdcE+/OssfhoKhNUeKxd9tOs/LD/TRJGFVahXkMUCm2dt
2Iq0pH4jqFajs7FiKLOuMWC2APMLIKsIMwH9leVhjHmYVdQa5ZO1uJjezd6GCdaevU3tsPluLcrq
4/IhRj7h3zjRTSzFa0FWA4lgFg8Odq3GoS3ILMaERkatdyu8qnVQNxWIDjH7B9duLpYdeLxhn49A
mW6duCTy3u1kTifRUCWB437z47Bi2y5DP3Y2i3ylkQjwCWbA6eE8RAvVa6JNYkpNYlUJ8FbYg8Gp
k3HkwqTz4NN7IXCYrv1D1Mvcz3pbhYMDk+NmxdGttIvuoRnxqaDrwhWWMLK7SoazX4iJTzawWIGp
C1RuZxZ86h5tkq3WjmQtLETfc1vno16o4iOU8+hYN7h8ZJuZaCzBfdTwqbq7MvuG655Yz21TDd3W
L8/0i+7qqLAwPqYryr5Ryc1Y+1hfiGfyChwBCHg45plqmlHGD1Mlq9WC7di+pXV6tDsb0+dANovN
xIfyGLzjpI1cX7cuH5w5T6KMn38LbC99YqbVsrm4reg+AAjgU+id2QKTYPoNijIEc61S16Qjj5n5
8blYHlxB9uGalWntG6IvZKdqNNbSWqh3tFzOyxjERb8fM6VKIzgbOnsvuD+hj3m7Iri+bRuv1ALs
qx8XwRhXzQX9GNAcygXi+w7nB5LZ6NgVDP7nSo2ndzXPsDn7roz/5gWV5Ub1TwxhCcNuU0kSzJw6
+j8plHuPr0hu0mwojCIEAZr2bRizPM/WPkVxLpStKEfkumBsgA37Cg1MuFVFhvrkFLa1zV1qCQe8
JjDkXMYygb13Lsbz/+LdQcAe+oTZgn8J14gw+sSx5vGH5MMS6deTHs9AXmi2J/vkd9Eb2/7WN0wW
pp8vybZ1z/hNDs95sO/8CMsu6yo1yfpQEV4oBTd+tpTP9npSPTebjdpiSW3UG/5p1TdBxANPtQU1
+SToFhrnhSCXmpTOPt07ZO+n2eth1DUk2Wt/JQP7hItGrSln1pBs1hyDlDsQGXswkGtgHZKibmDc
Vd3gJQ177wKy/MNPWyzoIFMrHG4iSgft1q3BOUitzPt0NnMhai3HPE+JNCh9MSkRxBb05iHBpMu1
7yHu1cNTmSqT0NQt9a6R6HZqizN7Oxkj7glglEsFhvuYfXoAzrGvujEcI5mA/BXwbP4Zs9++j9IT
3zVgCVL3WtqNnsK4kWGA0HdU4vq4eUd/ZS90ggBHchlXWT2NzkPXZ+Q8VPTmZhHXweRYQyWCqYM6
rmaL3gEW6ct3apzHWjiTXJzCxKJ94l1KR2ktOv31yIWF01weLKw9gnePXBKSyGwy2cdNXB2l9vs3
JbqG5UqlrSlTrKwE8hDJhVPcuheY/3SIejK5VfQL8rxpGMiu3oRblU0g7HUJYobq1D9bpsTQbgQo
ExF4pnXSPnTHAEt/oeu3m+aarhiaa0SlN7J3oSJwjIHa1QnzyQcVyWzd6Iy3UXru2iMG1/yKT72d
lmhLIr8RxIc06bs3qeS+a4sQ4fgLFgTLBH94/47bajHr78Uphv3MvCBWnMP3p5oLwXKM53m99gvM
AD8T0lZBAZluMcSQkFZcVcV5i+91ZMNemVqVeDEkcNUZzw9zNwnBTKDjZfraRPqCEqKHW0w+yKZc
lsV2Tk8WbBAO96EO9QeQ4ZVz0ArY+unjpIqx+uLmQOE1AoAmemXCMjtJqdy1B7wqmKd76nQ992si
0jN7a+tx70fauFrY8QJ+eBhnes3sfTHDyb2KDD72ez4HoKKDedMSKiYTW8ErleDeb+1cb7sM7Mse
Hklq2Ik7dDlafs1LnmvLh8PSg1n8vYBBB89iS+Kd0VjZyZAkRjsFB/Ptb0i+b5LAO+pdYF2E1UCP
4kcQhNGQlOEDS8UhpDc0FMvtJRya3D52lUyyMTFnTuz+Elg9HGoXeBbl0w6IQEoby7EnkwXcCqNq
plD5xI0ynGANMMzhLBXBd+H1JjJ9BtR3BRr3np2JDE+c11C/ySuXgjXfjP+HPI8E0eWDwM1+Yjti
DSslBs0SCzOanuuCt3KYvA97N0dCi201BAPWg0hmKckqYsqJ8Ew+DDgAnnMrprqw0nOTClI6UwRw
twIf1SHfjjzbFv7IFHVqP3nN5eNUUyf6r9cWGSyzB47ZwQu94HyXhDJTpI6Hx+we0u3tRNcwVHff
LOmyS2el3oZC5zdnXfQCtoUNS+f0jFfywWBDfmsr/5sW4xa0kCllMRPfg+u8wBXB2H8lxh8T7oZG
anfAlC2OHU/EanpqVY6PVOmcN6cFWT+c6FS5LcgkFDSLNffrgwtE/WAbrn33T8VHpT8QvfRVJD9p
augbT8ZPCrZU7xniII2FdTKDpSGX4DWNrmfDizPt8MYw4m52QRvRk422sz201vLAITjqNNigyPe7
6i9EdGcANrJNrZOMY/FGLeeMvFc7W8uoSCCehb7vO0vbQBWFZnp+NEp/gnshw0KuyHEwjjxikWKZ
v/HX4Yg6OrA+tVGPosYBtZD/wRL5jzqlJw2yclcU4znm7yhTm9jA2cEjE9DOf033RnRnFfMkboNF
SOk/MFIg4sbkNwPQtEnnWU1wEL+68c9eRKIu/vTz4L+OyxnLLdZ37OyKl0j/Dq5punpwJ7vndDo3
IXxtgLQ1ql2Ud4dCTqhRRIYfKJqC8GmXOlF8nFVxEklIVDmSB4N2MO3eUHSujL664iEuTDhBsDpl
CChG1U9cRmYBy7y0uDLXMwU/p2bW73vxNAKuUfgTuEEtf9b/ov2tiYFW47vsFj6grwzml30IE3rD
ZJ0nkoAuDq/0F2/lRNTat+bYOdUhCQwaj/LXDqcxhnk9EkYRgJZAB/SSuIU/3Y41yYHiW50bSnvB
3C8KbBkgGQ+1QBglQ7QTxa/wn2ZfjgTXzLiDTv6hJO1Vlcqa4QsGkYaFVn2nUmBt1mWk6ep24/x7
fx1zQFYKjak2jlxhQr3H4/B6vENyHVjCGQ8JAR5IMvCvLfHqmriJS2mIQ8JELRBh1WGctS3d37Cl
l8O7so4c2iW6717he/0e0ThBeSjKU5eHbWGY2NXvV+muzb9e/bSslpbmMIjtitGYWVUkFgk5V3Pa
jpqDixV9U0h0DEI1klHXFlzcCYrIP674S0L2Heym+81urW4h+oTno55gCsvqVrhQTL4pwqiUgEEI
02jGBQNeE+2fxTCMncxXXu2UgK25EmA/xcAgAh7XzU337c5P+2kA9vmwdUi553jNeTM4/anlztOe
wwMJKwSNPg4UX3B0kTpcJuQuOeP0zHuLooTtwS+VU8ZaBBfx/Is585JCjXXHwsUYgIkOzzmfEGH4
OIVCZ70pZCmdGGkGgW58L9zouFAP2rCa9IMq34OGJNea+wA0H7ro1pbQrZn6jkw1lHO6ZsOEBevq
b+KdeCBg7ZHnT8TYt7h1FiY5lLHvPq8tk9w+ev5zdyYcoiwGExJWlCOPTLeT/XgUvL44+RYCd9Sr
Ehjp0RE1GidFdWbCVVYtMazDI2qRbt+FvBjUvVLYzaHj66KejUGkWsRx16Pp8p5D8eW9/ObN8bfm
rl6TKBfSeRpWUM+tTr3+8LUCSzFD0/XI+wtiNW1D8y67PW51VcQdgLrHJ5tKLbaiwCJ6TU4YrHX9
u74CIR6qY/HxSkvI9LCqKCtCc2cDj2udA1sLku5BnJAEFyq9jpfY4LmaYwVsw8u1+LK9Nk60DXOV
joCScQlizdn4wV5wI3+is2F3amHXh7Z6jyeT+nQPk5NQFK5mDvGpbNpJ9OcO3x5yFqzpmhc895UF
Z/JLiAis8cuKxW4dLxQ0WWRIfwBxDQOhrzGwp7Ufb9aOiT0bItwMpP5XOkpKnK1n4oeAdrhirI9k
OVQHCZPZMDfuOYKExuUl8Fn9IL1hbP+4iD6zisZ5B1BXN7b0OgQFnDLUZOsTatQShNFN/LUyzWzK
ihFbucBHMZ+ihRjvEB90poRoD4eyKjHqpJTz0gYO90VnYM25PiQsif90OPIZtnpH26UUydm53O9F
oFg3Jg3w++0XdwRpfLBDwT1/sRl85K/r1XhCLj3DGBKkbLTHsmOAA9n6FisQKngRotZS978hkQUS
uBuTA/khumLC6rf/YbyAwrgDv3WKTUC6oXig7u0PZ4XgM0afnmQdz1jyWqPr398HGEruuumKl8mw
jUt+1k6/c0clbWFC6LFmQtKNLx4pfWHdszKMcCk1qP0ZTIiKlJvhO870EkHCZKg/HjuptB5OtusQ
la4nueoz97V9XjXIOGozu2EAmE1zvgghbgKYD1ygy/eAslYHxxjXM6/DneAG3+QZoAp/+IhCXx/t
eOj/QaHiyOYUXdjz42TimhUdflCnePGd3GeCmkazyxIAMe9ovok2jrK+0YCSG6sRyqUcE5UwaDNz
fFuchjJXcEz1skw7UBg6rpnJ8XXCd/GdQ3SBFCdTNdLu9ZlJw8Ax4l6bxlUIhxhhY13OqhC7yTD/
laxBLwrMlA/2qJeDMGA7tsHEgHcRzoArb2Cmc7YkeO7+D/ex/nb7h+U1irEdT9mX61Ve7kTooxug
3p+NPpe3w5T5FTuf0q+iFvP0e7qglWyKfX+wD6ilKsDameId8qR9k66NVdY7gP3TvdPndbArQrDt
VQoa1qHubeVV4Cp1feWsZNEIqEAFZ9WgHVafbxf+f67bqdiA6n93B+d16Jbk9nDjr/a+41nIiHzI
b/Tn0Jk/qq4Fuxi3lhS4p6Lc9edAaoThrKtsGyJmwMoNSgduYfN/XLYKO35cAwARSFCP1E63jUT9
UMNjwr4x+lDvyALp+w4zoqfdUt2QoIF9EjauWYvQsXhx6eGJ9VmnLYNi07sKEj9ydxKwC/JtP59i
GusBxvxV5zpdiNzRLYrfZoQgZdbfyiP1na7kutVNmBP3HNSybSN1GihG2CTFrRWs/gfcMY95Hwpb
MIVeXM/+Zy+OaghY9oKEyTrPzWnvdDIVx60C139DIH1wRCynjRjkyGkQKiEgn64KVpJmoM2kQ//F
3+BTQuE8I5BgbI/2Yl/nub5qCFtzZQTEET/wR0pXdjZZaal+J4wSRxduCiwu6rhouH0NfcjvdxMo
cZ3WErg+avBEzta9fyj2Utxm3r0bVFT7GC38dq+DjnCUBQCZQ8ErxZtHvrTWbJvn7tEMPI6riR8q
y3XNIqp/IvNT4yqvh2Gmi7jVbX0lOsS5mYU2DlNiLN8rav8UNg7c+4CAafqktU9fL6Z4gxKOufCa
XsdEKpP1J45sCBfiskLDfHnqB2EJIEuxqzzRQGtoUdyRGCtFxBBLgrW8TDxknhHzmF4CfduEA8me
S4RcGLqyOuQL70u0QVwdJS9sx03rGHwVp32uX0ZGWZ6KkikLDpARSXs+pJCPqNEcrJBFAfKG5AFK
bbpnT/AQYLmRwGtZMdi09YqPzDGPjZSM3vliMMO0itJfw3MHmUD6a7YnY55jGUpVSP239YYZmQoB
GNVJ8rGnQBytiqG9xjVzn2CeodbGvYhyPvUvXPBqUHTPvhvVRA59xdJU3JMQsysQYIiiwa6Jp3Pq
QuFkLi6q9UxzjJGT27l72VIhDARZ89MtC+r87nAgBH9Iso6Qi2/tOqF+4l2tzWUamRFzx5Ra+s1W
rqzMUnEbsV+wOteAqqZp1PYwsdGDESws/i5Joo0VMIFUOqULS+cRfZZDBeGn4mYriHv5Lo49s3xZ
f25GTd3hMgfO8aV0mnb6g8YoAcZ16QiwuttNGyTgva8CrDO7VKJOAxohk+6TZqp719l+KSuqiXMN
K1kAX+5ljGBRpiNEkI19kORA9sqIRTSzDkk/dMyn1UJLB6cOQp7CAp7TpsMDrtZWtFYtSSobHcOt
k9mlAx9ptxU0gCQtZGaIbMWlQqmri2c/dXJoymk7vRVTc13k0j/6szsAVL4CUgMvsvxTEj/YNHwW
ii833LhHfaHK2yZbs8BUJEhnpgcdP/dFkEhh96M/euuDysmwBjlF/pWOy6YLifMUI0ImIL5Ez9Bt
1bWygeNoSkh/ADRQAMfYiuL9VhSO45zURyqYe4jS7RO7RmJm+fnNIGIChmr1e3fEkx5MBEDN2S5H
nl1LvmHZQVrLycdEAeAmfggALHVLeYSzhEwnqsEV6b9nQvKYnqc5n7ahs2y7NCGWJKeHjN0aj2QY
urMsKZcuGImekGhQE0G6z2xaSr+j+4kG+7+NQqh8eKR4bvStQpF78F7+rgl4BW0WZGNwlwC65Xur
e0SnjEP0KPxG52LGKr8w9sZn1Bv458tsp6zdv2DXu4VJCQv9TECxYXOCRIyazXaVsq0O3UapcBP0
MxAZozcj3GdqyYvv+HBsTXzSpQuwf6GU/hxyJoqVG8Qt0mxzs4uR+mccnI3FsO8FZoozbhL1p8ne
TkR+wU0N6PUaSkNf9IrzGCgQSLIgIWui+OtxCCxU8bYY7nXy3CF7mYxUXRyEyq/UhuOH4VXTZ5rn
/LzeuaU9Tc5NkPRdhgTcXj9Nj+l+dbhDoGzajSlPw6HaqtBokicjXlV28a9TE9oU6o5hOSVgs59E
wB9SpenwDkSaCtmbq7tYNDBrm/rsrfdW8csq5zo/hccaks6qL5PDASplnddZTcBMR+qT8t7BvZt7
344yvNufaUCnxZVyh5TdlJyzuATZGsuLE7E+Dcx7T9Tep5DLqelIfH8yhZvDh9xPKKfIHa+HCDXF
HlJ8GYBpXs/aANxmxCYVa4tvSDvaKydFskkFCgunEBiLT7/I5knUfr5Zuysz/VY8qcPg+xL64veT
AlFM7L1cVQW2nxf+MFpw1UipAt5r7LxUCaBgesYA7XLSmTCU/uDEhjt812FNyRlDqGT2P+rH9nsi
jU+xlRVq18MnOs45PctIiBzLx+76vjFm5cc0fe93dHeTsk965PQClWeZ2hd0sotzag4bLzDe0hG1
fOKd5iuW9ZBzqwXuRt4jUMSLitQdFI7q5xRuGZXt7/sQ5vr9KSUpKTOFhKtf3FIWfuEGnIef91LB
mkkStNkWCA5Q7ANW+faj5n0FyIg3PmcZq9yi1IbBdWsCAzCOHMXxyM7kMxVZKvS1bG/JQT+Shatk
56SH1ZD8BEJteMQzQwo3ft1Si2u/yNQI64fCtZsJ0RU8/9j+Z80G+hq7DaI34P4qMV/6oU+bQQ4e
6RdFpeofYIsKpm5FjVS7PMYKdxjF4VyfxWS1WHqNDWDq087xOWd/5M6BSGNOnzayrNDXwLTEVHEi
Sv7ZXmEDvdwYITvkkpF9WzS+Q2c4+9nO7NfEg/8WB+Jxg662BS6AJWiOD9D47Ltdg8yGwIS97RrT
LNK2AZnlLOz9XqQ0/g715OUWowNYSPiAW8Qevji8xAaRquOcPE9BRtQG89X3+c7GE4iXs+G30inw
0SctD9gEVpXt4lDyke1oamOqFOtg7MWQ48QMm9WMnTeQ3WwmVLkPW7gIvXY+QoyEhX9V6jsmwtSU
qstVP6oPJlhSvXFGxcCaaSECPkeofrjaZYm68OKqt/oeDdKw3JR0TPikAkSrjUjzUKbGK8Ky1Ee5
FxT50tKi8Ldz0MtTSea199MOaPt0+fCEpoz9Ak/fS5zA4bm0KwYBv0zNYeCmpJJSuN1539O2sgai
C5j12LaqxLvVrt8zAjTUG15QoIwG98ROE6ey7jolyj1q3ua5zwd9WDkS9fGKjzK8Zb3jW8/HOlGd
x63HrcvPFF0pAJu2W2oSC/4d4r2xZQjBb/KX0ssT4871qs5r8dil9OWPPjWRW3P/l15xMRbF7uGt
xzueWKMUjuso+sh8V4tYPAQBvNU4vfDjrn9wwwKnPUfxRgIOAYoo/R1fP5MvuaGLnhUz3YmGpqci
jsORTKngpuuJ87O8QZz0JVIT5F173GCUJzSDM/0k+KzyPfkcFphJMtPHK/6rKkIaL2/vzDRw2UX5
7N+8Wu10CauCjxykuEY/nkM40PqjCShseOoKjFeMocK6+7LZRf6+AIdy0nrEGIPxCU2Eh6CUO/Ll
zGYlVTGCZOYQ4RBEwZ8xse/YmypkaZCBLd5tHDW4KPEzlpvi5352FFjL9sHmLYarPOgePX+5oyBJ
6VA8nccYKVfCBFbnMz0dy5jDHxEGCDgNTslj1+z/txLdAGMVETNugTf9O7yoocHBn03cnNX2uhUv
U1jlzLRj+DQmWfQ8SXmFOsLVgXFOIYQJ0n+qymGNoOrCRZYPwhE++lAlmE5KnpSfZ3UwjMLT9kB+
kAELJ89V1Wg8oYQoBgt5SLyJyhdsMGYbZ909N6XSdlq0OQ5K53ovPbu6nnqe0gVLsdw7Ts8o0oB3
hn2BYRc9Er8EaoomQxDPLzr+XyBQ5H7ZsazJLKx/RAqalz+nb0/c4bVYSxzGCHjOj/LxF5GDks8Y
EKYu75e+KTImEO+17ojblZjRu5B8LE8UhbabSNsAZ8ZeI8LWUWM/W9p/fC0NAGixMcRFL7QJrkgp
Br4g99ahajk5KkDfeJp7HXP7kgtgr6bZ66x2X5PS5UeRzH0yXOO57KFEpxNsKi7x+9jZ9Ufl64E+
uCVcMu7xNd7upr/mv6WSvGKQdc/EhfTHK5wIhsNGFaMB9d34gLGBPHj49HGaLkmkbwHrpJfinzM1
olB6fr1QIh08zaU/UEPbatwqOBmM4VyufEXDpuromowi/bKwfadTAa/WsfyH2DW40L5wR5E+Mip/
wVzedof5+axGVv48EQzifyh33Xz07WMbryQJzREs/2GrC36l9awdGTdlXVBIN2T/W832O3mjShV1
bkxYluOEGYweeDXMlF+3hSr/1Upvbv4+SeWDTht3DtcXwT8D+C1wMkBb2vfx0K5Q27JybZzbuKmU
snNbVHE8exlkZhbywaI+E0EZJIhJK5zxbSr8yGMT9a/hMzT+K+TUe5nl+2qbhnQzMgfiaIVh0pZ3
pps7NxEavxpHRt0cO8Qi8fSMpOzWT+TQwv/8zQzItLcXVRVRL4HwSjAEmfmDJVBlXYPsVmBuWfbY
9EpgjK2OdsG85T5igJD/q1RwUcoD2cLm7dhtvWZP6zt1Gna47vCaLSmxTfISfozhPBVcdrKwVtev
lqs0UEvLlX5yJMOztrbZuitc6En6fry/a5Z7xR5tsM9d1Mp3CMDAQarlBb26qXpjo2Xzhri6Lyo1
h9qKyq0Qj8Fqb/CFlzwjZwNQ0zOPA1EGgqXw+cPbT96JLHRe0Es0ahp3ZwZVUY0eNK9LrStQQ6E8
sBcCQ/0RhHYZ+hoVeMp2+e27E5vxoShbBvWJCypZG6Ez8sa75LL5ThEm94Nxn/bNKWJPeYCQQUN9
3jyba9p0BBTZ4zuo5mI7jqb/7TVcbqI/tBfI//VYbNaPdLWrPfyMiAZOVmJs05scjurAWAbJGAQB
KR7kceJYuRHXWMEjrrije+znsGk84VF0lx+TBY6jBkLXh9oO/DWJ9Z2bmvaiTrCFwAN8oDJxJe/M
6L4U/Esk94bsn0XSUY99vxr6QQHBbxC2mz/J0JEd4VThBod93ZC9UyZJc4MmVIHzB9i+nuuWqSN7
4LNUGiaIeO0PEsRegJoSVUVk6yRC0MzTCwSrRjBp/4FXEpJoHJZbZQFwnTqK35LaHMYaWgigJqEL
YloCswt1bhsWbbRdQh0h5QYoZJsUkwjhOzWddI44QcFWf0pMiJYwVB0VeloLYMO0zYGaAHZd4i6Q
X4VuD00RJzyzRFpm1eJHhI9JuYqaSlsViM7vsUarh7tO7aEhbyHPziTSenk4VDB+D5OzgE6RWdvj
CZopiqv+pRBiRvb9xjfhe4tt/l2dObyjPnuEVGxzKj7ZLXRzToQmxNnFhGWku58KIyrLWPqPeQUG
6E3KxjoEJNPIUSaj9x1b57nd0iXBAGhdNW+GxMB6PxQG2CRAV0UBi5rWH5+YRTIzI3zGdrPj11oP
j5O4Z7RR00UjQR6SdpYwvgcT0T/6aInHUKBZe/j0NZ8MKEc0faKdots1p9Fh7YaTXJGQp4ktXwA4
4/JpbZrG/Os7nIFZ0BgdQgGrD78mTvVjjVDAfdPfCqbAlFD3Dw6L/hHdRa8jvagAoX63tPIfeVRA
rXkhp+UlnkEl7FqLTvoU95ujrzFrbg9JGzIT7QOxwhqPhjF3CEh5un0znmlQYlaSYySVfK4u8OaP
iMfO0Zu51GxX185EBgKOpzcRIJO2XqyTuNcx4RDesnw0uRj+/Etz3Ry4/7dqPR/DmOpS9t82WJGY
hOhaWiaE/Bn84xHncTg4uicj+TTtaoGezZmJs8QnvSUCmJP8xdF3TA29Dzq7ElfR8i1gHm8urng3
cm0zvWZMsWDYlRG1DM9GGT7Q7A7VBpFvRQpTAHxWapXgqyipq7p4TkGbvc7NYNBbdeLrt6f7P5Hj
fAkI7Y1wjlqyzYW/P0zHfGuQdGLvmjQ88Qd9Jgf+XmDK3pJOAo8xkdQLkZW8SrZzMjRfQq9v4cjX
uctMIv7RF7awBJiN54o++SnjxJVPzuSD1meiNKR7PEUOyImgqz0Tl5TGdV9Shisl0QJjuwzH63RT
UyLrBLWrgdipP16Te7CCSoN+e7ywz9UJq5LSn3fkg+pfVpjHlo5CmKCL5ibuz30m1jciNlOk1R3G
cTvvDB6SIggsE0A178Et23QceRTi/k4r//GN6yGxdaJtZiPhQGIQ4m6K4DyAR5OnspGvbmwrIunn
mQ/jW1Fz6BidJZ9I0CPKF6aCzqN+KtUCXruZ0FcEzAafeZWqIrAHjnSED0BSvxSEVTe9Hs1WNdqF
5iZwlfPwjawbmygMQK8060h5dYDANXldpeqiKUcz5R26CWE7Wclnjp0PD57Vg+jLv8FISv/78S6A
wZlfDySc9zH+LspI6TS4B/3iDW7akWWbDIAHNZ6wvmPYOg14T8cxeVFi5gO8U6bA1WTBtEYHuqOB
1XlIest8T53wR+rBL6xFTpE2mkDC/c5FE/S5tFGU2W+d+Ax/O3VxubNMERCPzZu+wFtPKkNBs8/h
78faHVqjHj/VYpKB3KDNGOlGyLRq25vyBS78LjqGxKx3WKLoBIscT2cX0IX/R1+Z6N25JljTvNVO
kCIovd2ff3ZIUA6vRTQkqiG3Frdo5bsju9bI8apZ4lYvBV6o4gSppVBSymRj+K7wxhTgFxntq96k
LZoC0YhMaQyt/f+kxiX/23J3Vi5KipcNyo6ny9Jr3N/O++N1uiiqMz0L0q5PPWW2r7IY1pgNg0Iv
/p6ky/+AJBkn1Q+jlXTQPA1SWBHhiC7CtjIsxVIPogAtyYeOCLeoLY4CvNsYoR6XRZj+tRs3d1Vb
/BjW5ScQ+8Ty+XzL48nW5G1GXlWkrFCEvb1KK223FXtHqMoLyj6Aa5Evoy2kF30P05A63OIytE6W
lbCmarbpAAtSfrJ66ET08Oal51z+zn0TB2MOLdMib/Mm4vJiyEx+kdrcOSsh+u4fMbD/FUyRxmjV
7t2Uy9jGx0s5jltwvxYHu/YxEyL5BtDyshQn/xWgCCLR4F9OOuEJnhY4VNy0obfYAqStyyw7+ipm
clr4gMnLIbH3Uo++P+0c3Yq1Xby/PIS0uS85iUeG1zRMXYu5jdUFHczL92Bn5aYbsNLbcmPDuapN
jndoRwr7bpiaQ3sB29S4jnqZo0Ev1khI6YgZaK1cY2UHfxKSWMKdTJCrLWnU9Hpu/iiGyWt3flsX
iXL69GaTpYETWQ8lp3BR7Pd0cmfB+szUQ0AHeSMaCAaA/GXwMKfLQwY0hXwyqzjypth5FTjUes0z
InvMLTgeWJZ7UL4wbpXJPwO9rjQ0kEeGuOXsNO8p0w282aTBDx5Wt4RWxuK8IAYiz+dWasVtNCT5
o+wFpYul1Jrylo97opFm4O/RfSL74njTxaFN9pJYKRcc4huKJDiAuKUvRsfOIOVe/WwJx2Dtnnig
wLJFiERTMs8vI8PiORaANvQ0x+qJ9nJByyJRPm7J+sARoJCT+2DfJbVZLUfANJmdQNQe7QMp9PXF
n+jE1XZ98VURbsIEiaatQ6pTmevPSz/i/9PBn44F6mOqjkW3lDyBArERK3c1DgmbVQ/FouyiT2xB
6w0/pcwt3mcOaAJ5KmWP8hesku7eX1ZXhy426c2EuJPhv7uNCHK6LevmwX1OT4716WwGm5cnQ7Fn
j2BQufDUpCVCHiWO9F7367swVOP7KNW3UwU1zseLmN+bisURRknP60ACbStL5chlS5zAC6HYZ6B+
Oj6SHOwBYsGUXNGMcgWmw34AARL2P0fEGmyxGPz5FmKsW9SAOok9+nG8nvrUgaSXlu7/BQ74Gz91
hcolWI+mV6EhKV3aZuk44K1hVChnAMc7478UQs1Fvq7DFzhQ3IRFgQD1WurL5R/WL3yxEuggp1yt
pFU+zblXhEghRFlfW4mXn6Bh9ngb9GG3q1LyX5UxdPHiJvXl7lsvQwgak4G6T9k9hlfe+khoQHoX
YRafBA8ooAesJ8fK3u+bXrXjf4N5jA+lgPrwIJbf28is0V4bHae+xCCwrtEZOs28ysn7rM4MzzHo
BV/dxdncLCTydl65Gc4ZZpX2sv+yfEHj+r+rBtMOD0+m7FRfqwKvArTz5p4X0mzscDTt4pUT5ERh
d3F4hYHs+/1tTcOcrZQTgEMWBIDILIC7HgSHJIxLbdPX/r+lc3c/OsbOWK3ckU7eFNiAijOX81L9
7b/KvaPXDTjuz9kRYuQYj8QNHzOAz/8gGrv4w+me0xB4LL60kIAWBl+uMN0IYcCocIYppQfJhtHl
5I24f7i95uXp2t495QCGbwDAkJjV9aIBKe4RyE7SwgxHoK7DvsGgXPclV51bMF2TavdCIbnVy+A2
LILEbP6JeE4GL7fnW2GvMe1q/7OfKN2p4hnATb583Bp0SWgXtibicPzrhuA7Wlzy7nLiiaPE2BKN
+zKgZIpmKdqYFrwDsXloNCm9psK9ulQzn24ujfKyBu5mqvE9nYCOXJEPhB1QStGKsXwtNCOKql8e
gIOU0FY+q7Pqtx1B/bUbHTA0Y9DDEfk0XHkxhH+JOhJ3rCfgoczieFenzuA86djQAImx64W4RFfK
NCHvBse/JGPn9gLZwUuhIaBPdk2zD0348XTQQ5vcRtXyEJErqcNVUox7yXmloo+TArGW09no5SSG
TRrs6WhBYdIyx++236rJnuuyJmwCxPtl0stIsL/wAu85DHmVkmu4XtxTwVboR17CePziADTImlbz
PkLVpGdIp61VPT/5wmPpro6Q25IFYfhba+8QC/XH4riNXWx7+/8CSvLnUQ0dF+0jPazjBwtFMPFN
QXHcnvdRvGYCkx1m3CilVYjbylJF7DP3iJmaV9J0JIVVvej+tJUta66M2kiGuihQWIivsVP34X3t
CbWAzXLByGiL7dfe8tfsHV4q5paBcVrcaXmdUl11wJLLoWuOHH/F1DfIet3BWiQxr/oN1tnfkzca
eYU/fd++sScfjlpcZOf/R6F2N0obPdRTrvW3owzKcmklEJ3t0ucKxwQSqqk4jDWWYhXPrsIqqhTR
1nVnd+RVqTMuTAhWaBhT6eYo1g7JbyJy6WbJQvca2d5VxICxngmdL5rcFDR761JXfVJi8kFppTv+
fCFip8L0ev42j8AmLdqLTQSE3ZMKvQtUURpPgQJg4h/hi9PcF2P+bXSGEmeFf5BncjRnOpWywRMv
g0S6T+AB9j31JccxMmTj9GRK5QkC88TcYpQWwl9L1G9eeBrSojz/GV8M0vidVg3SYTxnq4vLILmf
kMQc1EWYJzWVrDAnLv7N9MajD39m3tJIa587glty380i9ie++Kqi52OB525KJ/EaKWO71zHHbfl0
HIvCsotRNPmZ5L0UmuvdHDQAcnTIAHQsdFvoc+m3akBbhWEvWBPPu2v5ZEiERbRwmz0HuaWfnWt4
n28aN9whQc1DuL/loscAuy7UJ6JPiAjmPFgH+9JfUBSWZQ7gX699ut10kusUKLZWwjgGjH4m64x0
MktQaXDJEgLC2YNw5Up0L2DHo4k8voY+wjQ7/FL8y9pw/LVg2USVqk9cdRkAwqGp9aNE4ZUQuVDL
tSv/HCUpbGmonBvwt4lcz8vVGM9tSBvVjBFVlzmZ+ZFjKzF7bUiwN7u/w5VZ2dbnUmgV+v2bft7W
ZHM+fzjsqHKVr0WfvG1lcPSPlI9F1bacwkFWCTX3TuQLj6LrgmvyRpOUjEJEl0FjE+AH4J58QmXi
mi40Zo1+BKmPmRmg54R8sx9Ff6xKHz22u6TeZGSGkeE7kwj68e6tLCFoDPykFEINXhE6EhJ4mGnk
MhMuc/HKUwWlrEE8TL56wmCffWIX+1Jrd0LUyLX4I+Ajwtz6UB+ufjbIOgrVxG3JoEdegtwwXno0
RnODXhA7l7vE/NmDtbf4tFRrlYFptl4GRze+q86V3PVXb9D+fwOz1OVKiL7s8UhnJGyrQGckappS
2CqYcW4uoW1NeAEX+oUIqFkkxD4dgWaIWFkj9II6xQ88T9EtbpYvHwAW5Gpnpi/BO2u6kdegLDrx
OES7AezoglpQ92JFf0MkRCZ5Tgpv0TJdxsb41wgN9F7tWfQMVuZfF57T0NncH6c9sFsIVhhH8t2w
5wHmmrfS4PTJSZrBA6H4zBUzNxSK0ojVDfcZVjEwsxbXgLKI3slI0er84GsD5op/PjeWYbialjns
E03lyyxM4Ls3jaQmbjDJwaEEM8O45UQw1xNpIYd8bupDkpZ0SmJL5AwKCcMaImNbQsoHZi7h/za8
b9zzgHt+SXAgfJ8Dp/prkE74lLgBCLCehbfKnUED6hMh17QPU21ahhv3Bx4XZe6uHjIkvwyLMlO4
ns4BX+2QnewP2gCR3C7JakcrrCzsRqEjVVeqt0S/5zha59Ih4mgOc2GiSxdN52BivPXUiaC2qm6y
lH6rOpl5oKqfxNyA4NnuceNH+NGIf6tgMIKJNfwrEVHnhGQwwxdmLgFqVlSlm5EQNGX6VUzpUib/
m77IRTuNtcGYMyRrDuNd8OUZe5tLZI+GfDzsUhb/vFYzLBD8tB3zHt970ppKI/AEmBjbL0PhLNww
74bo2QDv0eXEn2zVcKAR8jh4VoHD5an5W6Bf8N6F/rJhlIq1UWKWE0m1ABJOU/RV7ZZQTOz8dXuG
3jbzNLnAOek4QcLV/gVys1ql+1NATmybLVNckm/JhJJrwHX4KHP2qQBezAMxn8nDG/0Dc3JRVAjJ
fKNIVfmtaXdmtVAjtgou6MeAEpg74z2Rweb5oOuCOrZtMoASMGo3b9I9+i+XTL4frX4XXQ7v6kR3
YAbw08nKvbfH8qtGvbW6j2fYAqjGbvJfd/MlWQgzWXVAhAFIwaey2ZgFbVXn+29hGHbXP+6sRMTG
DbCZw7zfKP6WruO8Kkkk0HFrP5xH3Rn9CGJdATvCv3g6SvRahRIvDks0s1Uj4/wL+reS6P9xesJh
pR6TqvPw6p+oT/TA5hRSgxXVVNmu0NHW84GYIOAOpazWL98CnW8ei6dMCOiFaRw1GGTTfe8BCL+H
VheGDHT5IhfdEmHpA9/1M0E5MMOUKu6m4U5jhU9C+hwYvR55RS3ts6Lz0urOpuniX1Da2B/5/4RG
dF1cIFubfrB4NL55UAwYaSDaM87u/U7jXvD6wyy9xSE/eRrMkB/cbVP9SqEIJbFXU3rSJLZW4PvM
KxpGcvmlM4DJNYtj96rcL+k9rWQqamRKyorhnbPe84bGU6nTP5faV8AZjvVJlGNR/2fArwNPaBvV
jsHiYiF8Xgct7sCiLettNLuk0VX7ifDqA3mXdhGqoz0FZpH08iQ1ZERYCtDJxd/3Neye3SpUQmk7
3mP43/Y2eW67Ge7O2I4OZS98pqyxTrFFsgzw/Af8/Mguh690Dt0TVRp4Ov5n6JQaboViKGzthKSE
9AgOGZoXGRyVhSYW3IFv6IEZYZFIzdJhtmhGroO/Qffe22tbkOJdlH5pAHSVvj1SNQRMIzJerE5f
eTmVUou+whznRJnttCiuaeoc7Oydd1RDh+1VhMnR80VvXEiLBXhE47tLZhMvMPuRWLmFdTLriyTw
OvvGj2Z1uzIxyWDx/6yxgK6HQ5OJtjNjA+vHFOktCMq52PSM4RD0/AOH3uI7xOA+3Mjre0Ft7MZ/
OIl5rDdMmiRCy2sjJ3rhC24vPxGmaREd5roKFVMkqa0P9n2qKNSDXdpSjx0ShU7C2fpzvdgUvQeI
bTfkJBwGN5aj2g4SHm7XNjgb6tIElHE++beurXh2+J0HpDMzZzKu/lfdf14hcERZUlU9r/0Vr6Ju
JRpdxvZXyzdTeOBd8otQxapzpn+XlxFd1dabq2crB3A/bLKP+0IvT3YQXlXf2vNENCTg0r1Yj3nr
r2pDnkzd53scrTx3qd4HO1uJ4V883AUeL18MCNzo2O2t3+0gPvYGKptQodr2N60/oXUVbGvBFtqv
LkqsST4wUh+C54MYvTji3tvslmglfgczfXCiRjD0zegrbon4U3AFE3Df5nVmBBkieYz5vR/o+utL
+aCtteR5CuejDnJkS7XQWu7GasHUdqmRQ2c1SVsY3p78blj/W9DY8SaQIQeTUxbeFZUXP+6SQqUL
Qz7ftFaloQ7Cr7cxoyovzkz6euDVWyR0xXuiYjFUfF/NVcLIDUl2Nqo72vJ/BZN+RC+rdv6jLHxB
MYaUx8KA5ohKQCJB9Kc1un1c+V+96vGkaS6w3xfHI93cigr7KPIesn8f/d04kKmHblRyKeq5lEO2
LuWFBaNFcgbiL23LaLXhXRN/M1yzWAHWZYwSlz9OMJj9GdvEgcWEk6amBYxh8Dkd/Ml4ftCMyqme
83EM6dMHki7V8bELnoQyMY7C1USJOJYzDzIjGPLYbyLPGywS9m4PeEje3RjEDhR59cNSPmd+Xbg1
Y02pamtMmDqpXBjLt4a1dTYLPDnmFKlZBx9vh6b6bgIz6tRLi0gbaW7NRlu+rYpi+xc/QabmRh8b
6HuPonWJ/xhlpUePnTkesI8yPByoMb+0ikVtD6KdnTY57MRIecxXJ/zLnVMJAQKozNO8GrHJBXOt
TLD7rE/muVYeDJpaYXU0yx4zd+EQRNXH3hqA8JjMBuHhnXkRhS4ay7c8Xtq9nj38BsORR/U4p7J2
pmtshGBqhTzF7K7v2iHEmt7/BVK/sHoc0uz2UYCz2ugjykQrQwO74xa89inX+QzeKLRsqFBFN0I/
MqcZuX4+1YtOOhK4pt5McX6mUh5/vLKti4J91JHEa0Qe6BchjbRFVPJEbiBA6ppniU8wDkERUqQD
L1+amC8HBIo1J8NFTPfZD/VZemxWc5bBM0DGFvFTvbDfI7YmdjD5zjNHiGMq9q3KrGM97YqMwoY+
C7O4ROrnWa5irpnd/DU14mCH8JIFNYVkLyyizrtnYvdDip/zqGPYUa8m93arJoAjCrTK0iBF475q
h5kR7oxgGoi7Zigf1tpBvKlIQfbNMcMi0kVkyt7RwxUsWAaN8wI+ne/B74jAfWhTQALQRaYsnQTR
Oj+mzM7TygpzBt+sH7CzmJKSDcc/1bmIsNhQJ/yzbPvriDfvONwGjK1O8eIvTv/9WLqlK8jtNopO
MmmrpX8HRbpWBJbizAr87DoHNAuuJKGiXMA1HCuxZebxYMQDz6h65W0AhyonVKnWT9UJhwUVdm3T
bUeVDMllUK9908AnnqHOfAFTEDEIr64IIm1M7W+PUbjMyjim43OXAyn0PzKgpm+xk8PVAlMx9a6t
r3cTkWA0VcNBS/85JAWvaD7mAECqrkU66jnerbksUlud+QbqpR3QjRbupYTK7euoHeNlIu4OVXY+
P1/vmRvGh7ZlMLKyKslUGExphC1QVohTwVO4snDVilFUhyoq8GS1WGLNBoqkIxgihTlue0Igmm1b
Qlu5j+rWmRTYQzCiVmJFKUt5nV8vHJrv+XDdkaAKyZIf5qtX8H2btZ1sOmDH0Y1OYexU9NkU+R1P
5nxc2bnfeirQ6rNGkgVcF9pChOEUOhvP5Bh9UfMMMpGNYS03edYCyjx5aUqOsqOIwbhmzo/j6jrC
tHARZzLq5Lorr/aRQ5CehIfCqs//vTkut3ty8o9reWaGQUzX9wLJWqYZMhWbhG+ANVve67XsXz+s
nkP6NxyAsV3/pVpQWro7dpkuPXI4Qp4hOvEqewE7bNp41uRBEmHHsDemY7ct/aSoS74iThNgxF/v
/ubSJGDbwJPrt3Xq7t42EM4wgDUHIGyuu3m+WAGPo9kcml3Y2jcZN6LMtghICd5sc8fH8r814DQ6
CYXZpxczgGlGQ6kmIoC6qnxoCteddwRDgLN+ksQZevnSXefUv1p1Q7xonqk1Wms3LjoHLbVZTDdT
PwuER8hj1Y/QkPjUY8S1gv/jIARQVdpnx3flJIl5SwixFQv7iXJvVEc3vganiyhynw/YQytVHuTi
Zzvi4+AmiSTtZnRg9VDUSKS8dGGn2sYUoWYJwo/TRVo8PgXp6MDB30AMSWkIyUi0S7oNaxXVqt3p
QeCxLWtwF26w+idWdjXJSAhvKMmXISb24Pe8buHYfX1Ged27RVgMiTIy/kMmxD4D2UQGWwXDIQF4
sbgFuV8rb3t3w6yJV4p9peDeQNZC0PglaWMJMAPRA5b1tyaH/l2pZgVj3LCsbqeP/fBW+fS3gADK
lDAkXg5fVx1lzuoTamNjo+vqhbhHpFDfGQS68PJ+/xipQXS0ZlggkxXqBUHiaJWWCR/LuYIFadOe
cLR+tz+8xiwIG/PPqUQty/eCLvgRr+PFK9UUu+AifvG3D1VoXBgxl6/o+GBfbZdLaGhfN3Vx8++0
jubckOdehmDZadjs5Y3JCooPRwVd5Xm2baUhDxsbRNp0E/zCx5dCXE9AcAEvJvLBiR5Dy0GGLfaG
DEIB0+MSzrSoXrzNK17/mharkMDXG5OljLgnDmZzFoB+peZtkMW/pQJpmBE+8u4SXguVizN3QU3t
BFMLxA+lrWplUDEj7fcjFcykvkdJLYy/h9aKLH2cTz4OlH0SUJUhMwNW5oA9MoP2r14fDbivPiOm
viKpYjYzjBDJ1kcDPo3T4VXqvZ9tM0rjpve41Vkdxo9yUj+uXSC5PUSdlPJ7MwsHeaSccKWGF9bi
/jsuQufs3e8LMlTy/njGde/lGf/0v4Zi8Uj7FY8tu2axYKoe6Zsiz/m4KL0RfIVnJmh4+C4gx8r5
Mok6vhZofJCcoMhk+mt3wwH43Lg1tzhkTTGu1ZAYDG+VvyDYSkpP7OFAzqi9fqw0CcxbsJLHRg5S
OfU53IH/+skFU5Im4Cei3zgu8BfuGA0Pr2yc5yEiQ5bcBAQOYASn8zCug2HIoN30V/iykI3M2FaL
bEGbDQ7/zWcGddsr/0UB9js47Gs3zHT7trG257fRq2Jr8rUbl/QYi/C2hl4QMD79wRP3Kv2FvR2l
XshwwpG6qibEHRbtzZQH6CYtoRw53izoGIbUkmzxBfHLDymr5qjZjqI4AW8k21IsQ8Jz0WMIE/mT
uJw5lqa9UC9eR+JPVFeT+lW18LqzBK8C3LUbyVhyUjyQbtsMGuHbhrP4LR+FjBYVEcdlVfTWOZTp
AuW5A0myps3hvkQ7CfaXQ67C6rOpVkB1AJSS7p9B0uOaeO3iUZwdVcFKQ1hkpO+fv6vswEl1Xnno
iuc8shaO2ZFaViWgb8Dl3CoheWKmQZknUNuM1REvGeYStcrw4yVv/7H5LfoCXHZZZP5q79t46Edm
A2QyLPqnjwtW4Zg/X1Zxl4SIqpVfQoK4fj8jGigybyGEBf3HkXK0JyMqtFltYyq/+DZ5/sbu7WZF
CbKpijjRweflDN+Yu1RJTxn/GaDIyzD7qCoH7RMfygtxXuoHjUC1mQ5tLiHK6wkdIlGfIZwoDcQr
T8Bmqplqw7BG8P7oh+5EvPL2Ln5sR/9s7kzjGqwOfW+UTaogbpzEtC7SPe9vfJWakoLql2tUdBGe
GngsYnjN62yZW3LnsxGk0HX0XyQSTA6IYXxnOzO32ofbQNVD1PCG075dxZQ1ZvAFhzu2BqtDsZOy
wOSx0Wbw5O/3mbP1VAaFEo2nF8o081hdLLzIURAaLxbld0IHBpm9pb51CE2khVlNg47yA457Zres
I5gIvJiAojEvbYGe43K85Mtvq1dOsrRQNglFotyEoBPY2D236w8bDrTCsyWB7bYt8pDOV76SKkEV
62pkdW+bhjjGBKPQq3FjRpBpKjx+U/yF/+gU2d31BOodVbBFBY/DEMhUy0NvEIVpOOX8CjSEKVum
rL7K1CoByAFdr29JyuYn7KPACZCJlEEh3QqJ6lPiuWL9ROaEw8zoFwao0PkkqmEPtQSV7hlxRi3t
oCScRg+5WBll5FMz6RzhVEdDi8Hy7JELLltglSNbV8yWobvt/Y9WytHcZv/9ZU8xOGBcXg0NAgx7
3mMU/XtVwvbDNXETlJnrscAwkptgCqrkLXlakxHNHk6PbX7mW0gUpWRUu2T87LOSL6qduqiwEpgd
kyQAHcoZTHr3U4DSNRXGp7PK6cpKt3gG7lITO8bSEXeSeHsxB8I78Nk297FDvtwOJIjpsHX74Uod
Lekw5CPAXIr4gNPdu/TIHvtPl+QsYyJwwfbBswo9nwSVKj9uj7ieOece5JUGutBrHENNTFGlnJtr
nCidEasJnj+UlBBY09WEBfua0riARAeTbFH54UIdQtDNdhH0JOoZCfNNuOrYpWFB7HDvNh0wCDCF
3pSy6nasY2+p7IPeeEygXTW645i+nd5GnTN59W7qy3gf0HrTIDTIcWSfoZXFcXU5/cBYVP4qiKz1
ZwQQzN5nnw4cQQIoJhr7Wc4CPUpEORrkME1IvO5OG1sigM9yk4OFTUziY9dIoOgx3wI+eI2J77Ck
/ffkymuCFpgJKTKaHjGD2zaRh+Hd7Q1FzWU6FOWJn4oHV5TeTvurOVGgTk82du7CHk2lmHURfUy8
o1ACtevoGCaPaMlNSv8x8sRUjr3dt0I0wui9SdGia32uygYdK4KSXitG1/KHoaiAUgBxjZdhVGin
8+1KQ/+TcVs98r+K+uRhFOQ7VRhM7584qagyQkOVfITUfZD/sxz4jo9zjdL7VV2rzdXv3rdv9jRV
Ttij8qRj7gfKdUbIndVKrsogq0uYIWv8p1jW2yoR+dU7Du0U16AuCDzX95Qjnm/2kvbD4bvYAQXA
qzb6y6cQyskGTJjI8IRDDLrJFCa9F2E6ycutKkGXRxIpFyOZL8ZuiHgwyIIrql685hcSipiEU6t1
hxVx3zSgTMhvhCQGA0gUmscrfYL5AjyH6FzYh5qY35dkXKg5bVHCpjMyIggbW5FfB7SLp+8CgP3v
LMzxbmIy7VeQ/q4DHdyUdcTO/DSDqY+ZZlnydJ2RpfQql55+gX//wH54isB7L9BTe3RMf/VztKxj
k6icRnr+O01ZC/V4B8qh9BrZE4Q5rD2WBXaw6+oPnjbOm8tdmoHN55DIIYUyrbs2eFoC66s/6nyE
qNddl1g5qfMh/uy4VPH+92+Ah8DYwoL12/5iGLhF3PotIujxyREUvl66ynxENoGKBo019fS6XOIm
NtkDOynFNRqSQ6IeBlP60Qz5qazLb9s/GrrE0KJThdkfu+9D1u8zE5xSP/PX3Vv6u5c4v2KO7eBG
HqnsaicIDSHib6/gNGd9Rl5jlEKEx8uFkDnxkqn137fwTs8bzY/snENDIA9ZJRqoOG8N4G/GvgZc
Yb4sSGq1f/4okFdVM/4MxXLoNdoW67iblzLLq8EGRp2Ca3L4rmjIWOfVw0KLBDV8cs2qH5/n/HGA
33tzhjz0/AIDGbPvuez+H6LM3F0ZKQasVuVr/L7f+NCPIzqo5SZKmNTcLS9ExrV5hJouYePFn1Fz
pLDcDFsdyWmruW/FWUk6yrjmQyELyO+7P1wQMh8z4jAplbxowklbQ7um7WwaRnmF4FqMzzQmoOE8
ewLzNzpcyyRpx66zVYRA+a/wyHZJfoWHY2Uj3meH7p2a7Ln4mEr1KqTRMlEe3eI4SvkwydwqC3DB
MSavPtMb+tPU2V13fVxQs1aeWT8jthUx3c28hSQP4u3JyGNyQNDod/HOwro/mHygfZhJoYy8B1Xw
vgO69vjN+jnJEc4LXk0bEzWaa1HJMzN7aRDHMSOpUNiMVAmGsFRqSjVHNg1aaAhBex9sQSkGl8Fl
G+1cdgepOlKfL34SWcp/1vA3GFvJp5STL7zurlRHPF51DZA27VUQeSDWw2f/PYQbIISGYtflKV4i
MNaVer3C7nQENv6vMlL8WGuRqnf/U5MdAGk7I/Mx64LcGbmhRYtSK6LTEVl5XkvIb1WF907PrpBG
Lc3TTgvHYdZWrSrLkMch8eyCle5203IjyB1u2RrU6h1D3YE/d8cW+02yGUzmXSFINyRQKiRZH+Cb
1oN7uV0RfdM5EXJFIlrUFRct+k24Eb2Rs7LDQQzeVRG4J6hQPMuxll0HJRt/Jo2bmqdJiZOiD9MG
IVlH8QXiHrCnkRnFgClx8T6GNiclxTiXnWfMdaaPX/PIYqfMgEy+foIM3y/GRXSKWbdWhfagZmIc
k3vJm2GefsDBksWsCaj6G5BPyhgnzJvQ8rto0Ozzi030OAIb7GWZY/+gBxAOiLuCwp7+zApsgdQt
NO90HepJB8Mj72zFOjTfcY14CbsEt8RiR1EeKz+XPWHjdYc0umXoBIpR4QHvBn8JLzks/I1hHe/h
suD4yQdExAcyXvbfCA447tbIzR+k7vsIVXRSOY+RUAzM+8enZywVi+v1sIukkc2+wHjY+Nh+zkn2
JotaU3z3VHnItPNICdLWzke/sMnmtfRsPe8UrclJf09B0lg6UXL2iaqWAv64P1/qlJklnoiYaJfz
ZCJEDov04nkV3pctl56cjURF9uBT+xENu3acSCLoEw9Ui6ecbPmJwcGGvp4BU6XYCtEl/z0XTcV9
480y9UdJq9pxfnSgIdqJuXhTARhWwoelKAbJYS/+JLOczF25dDAD3lHlxaNVxzoFzTcjbZWNzvjL
v2rP24zPNHQxrPsO3LBNyEBcLGYe6OtquTCIH9Jet2gRv5ICWJ2zt4E28CUa948fKGR+5TIvlb/M
uquCB+eneuwYaEClYgkxPnPo48vqQPLoBnrPO57oG/3krk3umi9zcOcf2NKkfbnb4/MlTVr0Sn2X
min1v75xLqskHlAhWa5yTP/nbaYJuBJOnT8j5vH3WzBhkq7ce6rhfbL++ay6qLMtesISPXwJgHye
injIivUOt2QBH6WOpwBy3TQgJCSRKUgMgGig6aAfn3YivX4tVCBFtkpujQWXNc/Ne9UOOoaeKV1E
/sJpEj+z61vOoKAx0y7U4KxnPv1XoByvHZXHgoUSSVlZAH9EhVnoovBpBiX/BE3QG9zlxjAoJAjF
y5jkM6sjsZ0gGqi2FcmOSoTYmT5ZBbSgUdcxq80keqeqXf/GFgbvZD7FKmZusJsblnJprniczlOA
3aoItBlCRBaAqdwtAWo1zz0+OBna/p7vWILDpS9t/UB5KV5cT9JB8vp8FEF3UerSt7dFGw8t6YMN
zFp70FN/fDl9nBkAwmGQUwQAJmQ1g2FglK+ttA7wDVFIL72LFCpNHZs+u0xccSsO33FMZvZUiRg2
zlK5wnwUaR58CH3FKg/gP28Me+2SNYx+MEv75ER8qm7skOqS70aYnNxindWMbJ8BuMUbcttXRzF5
9O+/7NYpzPx2gMwLpQCMIBZWawypquwq9sy8imAP6uWGEngEw0DSz5uueqCudxrmhrxujgpd7PBp
z4t2kXgmKPCceuG9beLZsYJOENBQKnx0Pp+2ECP9PlRLvoyYdbwWiisR6VEVrQfzoHR8zOo+dO9r
/mYCzMObVfhbT11wkGwqvPVBA7MUtAXTQHh8X+fJl68QNkcOGhZuL/DMeyN+plZJsj4QP6LnE8Mv
yuBKPBlGRUYQqEKknGsCqooOIRsQRB8+W+R+FUXw7oI6cjcUR+DWkDH0fyH2eWWwNx+FWvfbhqqH
9Q4iWs3vBilDpuq2jl6JD5tSpVPaOskiKcKeS3Oi37fDugEj1bS8V0nVLu2Gqg4FWSJxvWPo5n8u
UxQ0+/AJ+hcq7k+yJhShmnqebgAkNGKpZeb/0fe6wAqYOqnsSPmotX1+8dutIZRJd3SJo/xVt/So
NysMSU55DJTtkaA/t4CMpggVZi9eUqNmNViDvqt7TQG26fHfDFSPSLgmpRMDUBor1xRcif4sTUlo
CgLn6j457O9o/xdp8aj+RfTrdH56CskCL7skHZWBvlZiJwWE8SyiyoOOjDFMm5zIfWnBcg1gpE3e
11oBX4qhACWRs4wmRrtkWxHTyQ5l1s0J/7EK9eZL0nlTcV0DbW0PTm2oDFhOsrSm22oXJSF1pZUH
ZfOS5KR57+9Jx94e9pquok0/K3lu/nBCh9wxLucp7t/alQBsMmB9P7CGjRmSD/RDR2el0qhGVBTo
f9uY39SUcXKbPFgJ7YLW8UukLssX8FP3q+bs6+F03+n55v5DJQL2hYyYrVrQOF1SJchHf8lD83RE
MMt4cpF02UF7cfIX/Y+JbR8IAqMeECCNx/FYSuCE7JCE3deXgAcAhpoXL2ZPg70kIzCvi9MisQ4U
ySOpk/GHU6Ox6BWh8HGL5Y5lefDW8iODIjG/gOAQ9zk+KZ4ATs4J5JnitGrZxp4ZxOCYdMBwAqLR
raOfuLIxehJAafxU/rVRHBdNOu7E1LqGLdIXghMO6irP7z7etzF332De3gkrl/0YLKAwYPBf/hcy
DMAaBvoMYnbM9UIGu8Ze05zP4bSVzBC//UvmUf5skY5PIejPwS1HahlM/IHU1t8KCZ42BtkXg567
fBfIwUhoN37I4MKLW6bJJ0HfQ5uqMzpzoGxOSatreLZ4I7CzzxUOM0fgLaTFkTKg0MZ9bLRdQdcu
nKAWNXajJjkNLtOeWuZtKE8INhU0y6i0/6vpzFwC6F5zt6Wy8ddkG4ZALv6eg7DZvV/8sfJGFLJG
spVpw4WyhHMl5b3sM3QMaFB7JVND03Zz1v5XYQC7zfqOa7hYyhv6k+I7lS9B/iX8NbpuFOzAqNVx
M8vlzUmGl55/UvKQQcMsqgEOveuvI3GsJJDzjQWlTABfFksZl33/rGfQgKDBO82f7bVoF6ZwNOrU
UQRppz5UWatxQIrrCjo/9dg2dUIOOK31dAZ66OXj6Cx9Zt4F+LxpaRe/r4gv5tjPL3pzpLG6jb8O
qWDVRmvGGOYmGRuLg+3p4c948PIbNVfNIyrblwubvqUasOWiu9VaeEKkpUuzAOz/7qLELlS7zv41
sShtw8KhxyQ/rz1ud1+evlKvVDZGmARZAJjSC+eTlHuLYXiFVaU8o2zuKzM/YLf4MiaaUoWSaGmV
Zx2QSACocSDRpCdcac7F6S2g44RCpB9DautGsEcAMrTJ67Ks2BW/VVTczQspDtEgiLUa+UQx65Lk
yaoBIz6TMg/0ucoy65bB9t4/Mn2P7IFfJk1TxelMIfpgy+1qU+IRWQvj3Bei3Qrt9mUTfDm253Zm
rcTilaUtnjw/w45R0tMMB0X/D/sP3MHmzQKFgKmqfF9a9H6Z9RiYdtC6w+Y727TLskiLtaJzCOFG
0LEPQ9I/Bvkh4XmJ3OxjgWcEcoHjqraq/BA5YvoaE5P/Oik2pupte9dbvnxP5sjvP5p10znvetIp
MY9AXWG7xFjt/5yP8Xg1GwhCzVk2Ghn3S/KDdHcWw3NpQrd2MlAP7xqgOGSbkeVERGGfsA1U1FPt
z4zScGfGeM7fL0v1V4jLyqTBQfN3xmFiN0P6Zt+pF89CVdPMJkvT932leZo5rFqEaN79/GQb2t3i
L3hcS2bojxANxLIw+cF0+zeAGNKchwzI09WwE/303gUDKPFKzN+8GXuykaYsjQfjCWJmjNMHJbS7
7uPDOGGzP/NvxoQC9AqVJE/ZrhtRPMAs0SM6C6l5u675ACrsGZ0MrKscGmVm1v93/kuOdp0IFvOI
PZiV/d2qz/i65IV34mqMCsGHQLteJGVTu6kgd7jk+xLvlEIIpNkwRtjsmZOks2ASO9+sy2Cu7Ik/
qPwCA2dvPzrd2kkhfG8LKaSyc7fFkIKyQhUhfyINFp9Lbn4oamYwA6uJnTwUZ3eg83s/lpE8yx9a
UAOArfdicyDf7E4nlDg4gRUe4BnFkPP4IlhBqoiEVfjYd4SVhpAy66DGNcyByj11RUCVjimj4VhW
o77LiO29rx9eck6mHGli9FTJdETwRPJGqoxn+aIS5y9bjfYG4YPNL5tPQf4qVd3mmGnviySSYU2Q
fKBPNX/VlG2Nd+tY8bygQ08tmr/ryTAZwKwcIEkAy/CVoZY/VPtf4nRCHm5+EIYQnPVu3nSn6MIM
07grO5cDvMl9wYfv33bFBTr3tKubMBBjjVmPfyDyuSJ1MP8E9fdnSjxLJprrvFUnY4jw62iAhc1A
g/4PKtS10ftmc6PG64z/EE1oQkPK1+mODx0y1RNSy69KTYcjglc9VNE+hLmB1S6U9xZqs3hpWx10
hkPIfZxmwhgxQRZ6NU7fbpYQt234rJ+S99YXhuicD5aLFC07QrNVuq/0gL7YwZdHS2s8jXaDJGOB
ihVG4bPxzzI07MmVWZKknhiXpppfK92vfLRNumehJXl40DUaEDokFIMz/FEoNg65RLoJWglszkqO
57AkL6C7pmENLdmgLMXO5QSj7/jg47XZn1465tGEtlfskAUtw7qtovBQNvVGEvM4rU22fxLNhXYe
tnyVCM2+43kKKtGWb7kjyT05a3HAaBp5l+1PtiSyHpG36TS7v7FCtMuKmR9zzCkWIbKpZGcHRLFa
o54mb6b2tWWEDifdaEkGd7HvCNEhmQqWOiufRvOycR6huwbnXbLQezrHgqPjFolF/LYGed3gS5oZ
uLKdExxEJIISios6E0CV7IfJxMbMh0XasyY6QRtHWUu2oTvx0B6oiYpNrV9PJJhpqQuJYFtk7r00
JbyA1YnITHSIxLpAg3NO1GVTD6qZUGnTyoMvUheONmzD3QBu7QYcwwKm0jpZPrZ0jLng7yteNmp4
w1irC6oQ4WibDjkF7hbPJZcETFh5Eba3kiavCFooyqfysMEbT3f4U3FIoKK0ep1G04B747WnfSjh
jwjo+HHH4PmEyy0rcdcUfBTdlFMdMULmGMGLIYxulkzTeQQQdkjB9Yylzz8hKyZkwiSjyCYyxsa0
PTD8qnn5QT9y96vj0spiaYc04PjreRJRV3W4UQ3HwOm6RMRb6VsrpkQP0GsD9OFy9ovzg+pPjaf9
ZB6ZlR/vj0YyUzjgnrjWl0EFcliYUuN+yE9klDe/87TdxlluYyxg6lseMig/yzoiEYLpOr9GaX6i
HYHqXovJeDyuf+o/MlODyuZ/p6xSRaPmpzHgef54exaADQ2Dur0BDLsua8QjNRrRz/wE8VwgbzVb
ewiRoazbD1EujHCB1LdFJbepooZHtAT7SuY3zKkvX5v6nCZuPBWbqpX558PBw1zGb5DERqGfJg+F
81giS/wcHPSwe6gWbZqeARXWUkqOQU/X+XRSH/A0nkNWNROBgZM7Z74T89mZdcFoIxyS9+x731/N
Y1rwUa8i1WNZ7AWfA1Wg1n7BQajbfYOzhHUSSLOTAG9lDohkQLFfVXNBXlI4Cy47dIWgZyt5j7XJ
t+lzjwKOCiJwNAWHkOB84+iUSd5aneuDFER6NqLDL2K7PgoHdsXPkBGecBTeIIFJtG8PJM2DknJG
CfzZwoNYopj1c/LHWzeJIVhpbYoqPE/h7ecR/50VdXgY1Un+ID86hv3D2eHCd7i6+JcoRge2gFQL
q3vTqN8jEEzt0HCLge6GOGOntPlR6ZgQtF69/7453H1fOGDb2YFxpbVJ0cUJYY6Do7efbzu/GwMU
1Rp7IP9oeSAbDzWsbgW3znqYZiLXIYeMXsXFNdmwPxsHnBIEF7qJXtJWntRKTVqdc1lgzNpbFnLU
M8xRTvsWtJZY9O3HbgG1qYHGgM1aCaleSrmz+Dm7tVi5cwjFXXzdrAKbC7ewrHI60vGBcHmmKWYH
eZJhLu+Qbp3Na/UmBnaFjaspA1t6nAJwpjxRqCuw9bxfwZMLYsEbEjQIm/Orm0VxtNZd4CYZCqbM
aTTUqabgVSHWnZs7AJnlKjV0RIvJwCDv1bZ6JiqO4FUjTTC37slCKDzj7+tOkQLQLsuQvqAHkTjI
Vb+7stDEHLYsfd81gFLTctRc0hzlhv3Noz88+zHcQXfWOS+g4DFD70VAQStsWOfB6uboB43euwl1
jyu/cIMZtTeNmwMBPTr8JJCjr2H0Oq+rh+3uMMF5oZdyq5cEgi+4FXjxX1c9m3ws7NsRwDqbvQ42
lx0QmXoWMPhDv/FWdq4ZxuuRaC30kzseXbQakBuJq/NhMTYGDz5e9yhyt/scqo0ehnFrjxebqa2j
A9GpG21vneP7GesPEH3cHGGPMK7PhHxb+v9dr4JAveB3iSFLs1hQCukJsf/93BPU1tNLNh9wvpZp
EvMzzDW8g9MpnHw+m+nilHdAYlIHsbqyAza+6R3e9ehPBDfLUBXKwsjyvSo9gVJ64tUpahlfsIys
jvvkKKLMaZJpLxMvTMs6Q54Bq2f+Kyk3SfVMC/U3NPO94THMXu9WmBpLsa4mPnKaHXCihLgmX8Ji
7DQjW+pQzmbzQoCnHlXM+Wc8DbXCe6qQNeBVvBYswL6PhML357KqNqEYW3LjA35x43M7tMqKguzL
MJp6I+Nmn05bVevnS4TgnLKi4ygtAauylCcaqUHfAcbdNP6uYeDM7eFq0VaExWFlaTa9KyRsiI27
HIXPaopIBYwcm2UPKFxmDEAGuMDaZwLEbgI8/ycZdkw67PgcswcuYFHEYH6bSu+SIvkifejv3Blj
BWiZuy3l6+Npd5cSw6Fhrer+4NuhGo4YU8XZIGNPv3RTB49NFPUOC5FpR+51wSi2xgeb1wkUdVug
yf59ABncBZt4zEnfWjqwzOvBAJcRl3ZO3+ldwlgu+CG3HrVnO3CE1VjsWZYRdgJZeQRCNwruZI1F
vfjZmmKFjMzgXhdX36PocL3AA5k9JMjvQ0/JLmSfOWh7NJVmPXMw2qLckwjN9T/uovAi6o97ZAdT
w8xiDgwBwFpIAgBrym+HbDhMngH41zGh6ZsemA842nNm45eu1+1Ead+4j7O18Sfak6Z2DXZFCwdA
ziA7MLVg9kD1HCduF04K06OisA/sDm0lhkUsssclGl33as+JboEMd2IYXDxCZpAztvoyLG5TEtrm
7vYpv6WepmnhSE7BfxhDXBoem8Nc0KGTa2Q9xjFnJJtIhChSFf1CJ5Nw+2vD+PpZIveuy7smHGMg
0MkNb1NKsVOUtXO56Di5uxdz6e382zaV30Rfk6B2PNy2T/lS6hOsLLk0SkuARx1cgaTrZh/JfKwm
ostOpGL5BgkJLAn18FUJMXPwi/qoKlHbqbrOi1U3UavLLnytHJpOQXh5YHEwucdmdQftJkdVT+Xo
HouZTOy7rqgbNeSXkgulNlJbPEtGfR0bj1CYWpAX3wWHvyLKysj5JV9+gwI7ipTWtwsNBrU3CO6V
h2dMwwWyLZKo0Wdz9uEiDvXC5+q28JaaG5+HVdE/2pHQRdDtn3ZtEGMmSjdN0ZT6Bgxyyu2ay3ml
gRkO5M3nJKeZiJ4KnKSwp8Bp1wiKdrEckERFTn12ueEYB0cHDEFtlhrGFDDM8Z3WNTo50pnbydIY
nG++vbhVJFRpBGPH6gZtbFyxcNm5UQBdtSDONDmA/debdDTUAQLn7jrRII7RaPijwEAYNUW93K4v
GQKTYRc9XeVfVLb8IprMgz4I8cBRDhMZQuZRH+Jt8j8uMA5OEqwExtyvF3u30uxK4xwydUjRhMdA
+VYr9wMM+5d64Hx5t+3hqErganSV+DS7ICuqy+qLeF5VqEF6lUE8ALJ8PK38cqFTHqOxeriCuHEd
ATuQThy9FheUP2h3kZ23zXq+LppCeyCwcrfrCF+omYNbVkQI7yhLT9gwFvkL3TxP2p6x94Y2bFaF
kL/h66erB0ZiDobAKFqmctYIkk+gDlatN4JXs4z5o3eQSN3JQZ0hkQb7IpiqzhJbzyRByIqJXscl
cB4A8sVcY5aXo+gOilEohOcWycXCVFH50HBViPL9iSLFmsmykR3P9JO041M9vkO0lrHXPbOPodiw
hYfQw9/wiD9+8dDe7/xbq9nzcDDNoK/QNszO2tvEtMTj6DctZesEnegUKtl1nXChqfdEmBpeCDZ4
ehmE20RuWA6PmY3e7BQJg9xpnxCgVuo4TGeCqM3BWSVmURktcJSJUh74HTV/8/114gW0L8AsZdTE
J8Ld7TMV6DYrfTEUUj9N9roxQtGGMxR9GPr6QODaGZ6SLtkXE+JMk9hFIF9TaahgmjK4O/ZoaWGk
0o7oq5H5Ik132LdYElVJ9psfvYkOgtbjPlG5iT3UYPZObFTSpjDSo5bcXdxvnhAtjRKYamuQkJiK
PfWFyf39skoKYKx7ji5IPX+zqxdWbf9n2Fsv0L1EA3qXkWXPToDe2cbr2SGlRgbgwf1ui4kk9Qde
NfWbVbFnVi7R1RVWCbTvAkG1IIdcEY5+vOwupwDtim6JeIbdJ5Msl4PsqkyN4KNlPAz1ZeM3tupy
v2A5roYNVE8GL8T8OsJxwMCK8NBfDjxXyL6db1qWGGuBOUcL+eAH1xp+tFPY0Zcx28twHnJXaoPx
0Ie0Qcfp2h7GIrNgHaYUOUqGb0pl+mAQUHjxb/ubd7ExauLJ1kFNEPbrLNpXeQMRRpNsMVDySJAL
etMsmfKlLgXfiDQIkJivdhC/HeIT9G9EuGP9n6z84ja4/0VrMfPTMNDrSHjOI2oy2XJk8tbuAmAa
Qyw5D292LzHxtx4fR+XMpDD8QV7y3vnu4SyLE0CN6jJKzSJDmpzn+UJJyODCyLZdWnsiAkQw905n
wsiHzGRZS9IgdK3kndFMA3vPpMzzXK8l7hEzLx8OETMgVE9O4AOl2O98pAJD2vXSKkxwGkgrASrM
KkPw90Gi354T3gsExrXJaaa1oSgt2tWarFEEw1tH5AVfNW3xX9mPanmaBrzBaYUcBESwr69fqeem
r/l+v+UBds+ZgabKHFrRnpPuvhmSh7rXUZWe5tZGgh3eQzZNzkPOUyKq743g0kly5ShFMogzutaC
nO+6H2DvOxm43Kmq5JqzltKt71dFeuxT4XoSfZsPNR16phD+M+y+Yy89YFXdLt3+nbfxr9cKf003
TeFmas0pZn4OOQ9oRMS88BA0h/eBf6Ua80dNhclateutSSzUzH0P4wskUOP+2XNBGhWMM1/wREo0
1zCl2fhLcdk1CLn8nK8EcI9vMr8hTqze3sk7iovifDksUqKf43JxIxPjWbITRZqsulnqnCR2zQbM
f9akRCCr0s9L6qQ1U17AzyGbsZhrk+XYSFfqSaIYSwd47OWzRjU/qvU0EEdM7JGW2TzvzCsaO01X
BdsMQkUdmwR8aRI+GNsMRsMgjULXGgVLk2F3riWf7cutFO88q123dkqn9eOoYKgugcXMIQgy6Qlk
n1Vl2FUj2Yi2sIeCJuaw882k1QAXI8kHA6bRB9wpwoc7yzK8+vHul8tMzIAMfD/wSFiEvz/B12qK
IthwedZy51iB3G/XwVQZPDub+YSqQtuQDfPCVzrF5Yl13+0/O9Xs9OAZpvtdF0/nyyjhJn2yNc0d
9lffhj5sqb0C1JTrcq1Te9s/c8zNoP9mmJ1rUqGcCdis1srKbzBdVmUCj+GN+gqgwBtzgRmnvPhL
/s7snz0Y5eRoB0qN/vC4wLXN2hO+QXKL7fTGIFuarme767N2mLpozbnK3Ayr420KgKFZl5Z3VMX/
oh5OfEv8Pn40oUpJAzKr1+GkLDiX4YUBhRVlkb41eAUWdy1fPI6x2Zpa8FysVPoieNg4iPM62+zL
DnfzEzVyuhcgemOiNSRZrBBmfd442JKNqSfmb1MM0z3hReiYFw+VMTNCnA1/NTXcOP7ug+ZsSNIZ
AJNwSZDkc6dCdyqppspTiBa5xdwu5OcW/MrdR4cpT4bkB6h8VFMf04QKIEOyfDAy2ZdUPc1QWGsM
br9mekWL6V+EoazPOcatYzW5xeARly2bLbb5rVcJz1RZ4aumY6N2hfJy/0CyR2cMcPF30EA9kMPm
vji46I0fRsbyceUAj2zxiCfAMdUQHUCxQB6+CBdkEWv7KbZHHHi6jxbW5uNrWckeNoF7VrV2SCqg
hQm+Cnq8fxVV2iXp3arFo71/kws3A4zgDRVTjf7gxI2JmaeNadOj7qvA8rnlJwNPtrXaGnoQrSOu
BneLfwMJUt5eg926ZtQ9LVLgEb+PQB0c75W0y9mlJm1J3Wydge0BtTfYh64N3Oc0H7MH4usSCvHp
SJTu6mVs+Dg6uorqyEUCZPX0+9YZsf2Z61YTvEmtJ1L0uv+ZGgbv1sWQWAWYy8lQHNzpJezOrZ0Y
vj88DRShhEtytn3uLzmjfufZZShNJOdhzuY0sP2MjtOsyCKmj/o+D/lJBT4AYVVvWntE4XDaUmJB
S0jIu+uSgTJxi/kuz0Qfgrt8qlrGvDODvlGYuU8g8YqCuBqvNNqKOFWEayISmBK0SvymhfgAYr/z
vBBt53T08u3/8JH4DzjZYB/RhPIeOYP6CFEyAwopRQZ1Rz172FS32YGsA3LdCk9wZI4A6UTOMJUX
70YSgpCLw522k6SBE5vhM/OuekUukxoaga6hB1ramRYEtjSa57gja4gmdlyQ19LyEZUmpvCGwQ48
l6EhO4UPS5LCK5ou9I2HdEC5NcileAQXVNIrRTRemTWdB22WcEdvsq+EjcEFPTllE00ie/BF5Tc1
NSNqo3NbcVa5QcX/LlpL9qzsNLb84YC8Q4miZe/VG4SuX8kI7jUu0AjhxujJmJc9Lokhawf1wLwA
7GUOaowckWWJNJJqp4jaI7cKJ0FDLVfN83LvL1yDsMyk7dOlo6+s7mtKDvi6pNWj6tMsmXdHTWYR
cbFJ6rLnd/I5C7Eq1DaHSVkXCFTxJfYd3L8B1p15kF2rrcOcK404pFIFH1o8DldugJLgOxvisFT9
gpLlsEqbQfBUxKO8dnrY6cgNDwPq/qujO462iuW8bOfNaKsRGe7UQJUOWBzbIgSikd3AwKG/OzpE
VUsMtit4FVFP9iidhRsNs+ONfy0sqed7SSUwa2dxloRKuy0oLJO7nER9DcVy2cit+PZ8+mD2KvpR
euN0d3uIcteMaSUyQPUB8VzVP4CtHoQsP6klZqRJnQv7ZuSipTmlWLsGzve4trm807aSljWE6NIh
dlMC710dGPuiOm2tX78a87PCKqEgw//dvE1I7U+pEd+k4Wd2vw0Y8DyEGhi58va9NWR/XVvOr/vr
uHznizc/8sxk8DRJWpEmZKwRSHVGUmYwT+t/vBI6FQGv0/LFJOvBJE1CGg8VisU8IcU1q4eqOgkO
onkPnMNbx1bwV8bEhsalhA8ChyVAW0goi+GqK6u/ncFeTwdPDBxrEiaBXsYTuVwcMo1g3CuL8kg6
6toJNNHSrIM6F7IImvORv6QoSyygbOZiv3LQVuR4QzoeafJZ2Sv3t+LCcEEWKSLkkCuWIqiYWZsC
xkGeuJnx8DWBqLZXHll46Ph0GLUxuSx1tO1aJGAkd6qod+rsnqgvwqOj5JYQjOCpJLgWSXrNXWTn
XnIvO1DacqACcgRINYku2dkDIClG5G8Aq8fDtl8BT6ViJJp/1I7TYV7XkcEyWWEqz8JXqfBRGc7F
Xn+BJ6VvtOhNzVv3ExU01zD9HGUauGsdtRvvNq4e9jXkTJXxCLEj1w4PbhoMGSFgeRnpdsBYLhyt
joNopH15kJ18rLin+QXVBkzNtVXRXD4A8cG3PBjSvdA2Bzl3u70txKDYa1VhmUzkjpf3Yhy5sNBn
i8XLBdD38L7jz91twzkacyYKsSoqk22HzslhdCN5UNZwerEYJ1T8vJ89bEHV1VTESsr5cqBZ7Amh
nslhj/Eb2JvHlcIg2N/goooJvnLdSKXFND8rhYZrTfAAK9+oSIKKXmJBFJqQBN9D2xpq1ICvHmln
Gudwd0aCS0+ye89QTOh1ca7V+OLf7UGvBC2tHIgbLc/WlKtrXjkPoAhO2++IYSjfo2BeYXU4RM7W
0WySrzmISc0+bNZ3aTmPvqglV+dJdPSUTiz3NHT9V0PWFOjqAaI4iE/82IhQfZNspyIToXh6P5SH
1+UjqK7h1p3jXq51xuPTmp6X3hOn5/qy85vIT2LQ3zMw40N2W5bDd6WgLM33vJmkxFrKe3IhJZ2g
KJ1s21OQgkPnONObNNw3bwwNdujSdT/xg21oPd+bsth80ugV3M9lkPvBB7uts9k0ZXOnsjlCSPjo
CeDq+vwE5H7Lq7Tr0HI8up51wljVnnAULzUgNubQsdc07fCVzKQu1LNYwV5gX9aitCGPiwNfB9PI
Bogsu1xkeTCOQLSSWEx7jqeam2WW+tiS9bw0NYDvmeejhMEiPPySkVfl5ZVp7tPmAd8SYwBjWO9S
dM9rv43a2QKtXR8Qfvyna3s79ffbDKgobLsxs6HD5YQF9Kdl7wNABZUSiTFV6v14W3Vpsg52Vi2w
Y/E3HYbw4OZe/1BUYnSUcCV7ECqfDJcJTTX1QTiPOcS8YscihzgZjg5lgSwYnexgNSJPoqF+S2kV
Uiuc9lLHcMWkqbYIKCl4g66RWV951CVcmSHgszl8V/h361/J2UE3ABt7BmgrygyDAIZnLJobM/g3
xPV7z++l/1BdFjIcqfIqV/rJhVoaNrV7Ch8n/DmyKSmDD3e1UrlByEyKbUuwtFzTzCdsk42cXAKt
FmFCmyuFTQicNmbAMcBFZu90GHv1I7k+rTY7Wp93EYf0zseYhKNfK425n6DoNy690+37AAcqfZdj
4ykTjziN0htwnrW31UIuk0EgJMJzcq8ePxsUlfYGa4bHeFMoSK5V0FCGJ1s3Rf0J6U8kyKj6Bted
TJRUGwvTKBjoO1vQMYp5N4o9SjzvodaWonNnAG19MNku8lpsfede9j9nnTWUoxfKrrSn54FGCWC2
e1XNFE/Infe/KeeW9c0IUQThN4hDhC58rwQ3iNuzstU40VsHHtsR9ZwlAVT7PORfBNcnsFoOMcyw
MF0x/vy8XlqIZjs9Wcx/6nx+tFEex+W6ws7MtmIl9MZduBmIQOrclCgfpu4I/Ag4oCLPB2fnjMwG
eVQF5RimEQlB80ONTRvfE5RjP6MqkAGaNv5AsvPmmKXG/lUjudaBMrd0m6bqQmledFVij6F4+BHD
3ZJ4yiBYR1U0s2M1j6VFi080K8/WBIONKppmFGQv0qrXnAVD4HpAB2indbLHF/xrImx/umKlmyNw
Iupfc6Y1sR/t9sdw8UmcCvwtbDjZPWI8BHshhdY4DzMlj7NFP7ftPQtfUa6LAaB9CYxwzI/3H84v
q+Swb3bYJiVN+HnC9mlMIZc00MndAs6GmHFOLSZWGHU2fqA/cmUyZxFemq0d06AJcvPrw2KtNDC+
+r3Ak3ylH/RXjNdlaZlcmBfqAijkdqsBUUoSx45T663HewQ9bVLzCpJKvuahmkfyYwXpaEBPgIlR
4hW1t2Pj2oAXQ69J6aENrcUBMdh1oBuGGWIUdh8QMB5orw4hyNSNIaynWTUYIdxJ73X/fX/Jt0YI
J0ynQJvEtVvhxhnfDKjlnKn9wJHnzLsth+twK/5mco44j6lkbWdJHdSM5AabRKRSZq5CRLabZqbc
rwQC/LAGLUQB1qfP4x7nLbMV7dhFIQM7kgwFwdVNhqm8kw8xifhMGUzxpQuAFrG+EOPvwO2QEgpJ
4J6lwrBdHSPJxdPLzvb5STJN8cKC9RDSjD976yV27p/nxa/X4VHYHHvLkomRGELAtGRcr7Zt6bDx
3WYBc3mRi89rfcOnprJnDoZkBnGhc8HmR8PVDqw7fEilOdnVWp9ymlofC5BZrLohKxDT94+rTQy2
mBtfc3uZAo4JCwS+2BPA3f5ULV8JrdRveT/7SlEJ54rK8i3s37GfIsPy2lHlsuftCHDSrnT/gHIM
ICR1mllr7fNAeWykrqQM0hNc/ysdRKqcji+93BGLsnKvXBiPA8E+Z8tKXCKXF6Am1fM25ZGlF0cV
bFyGktep4isowtSIvPs4Bi5Qe8CuD38jXYex6QGvX2J5+EmF4Cuh2Z8kXYMJMbN6FI3kVLbilRtt
hTjH2V6UazKtRk+vsApBGObGPypjhpVFjmYk/9tZMpSO9K8/24F7tdZlt2fAkwhplPQcfZYRV8K4
LFKrUvZiR/usXKs8YDvUtP83Z5zQcBDZXH/26Q92z/Bawd193XiLwfyVkdUeoVUC0JDq/WJSKqHy
FHIh2NnK+plJ9pVRw8PkKYtYESVQPCBxv+5fUvIOVhNBY+oKXI8FSpuWwQkgNli2j4masAqKuwci
91XHbPkbYBb4KVVOPJxR6oIgHBUMr3LCd8hBg8Z4wiEyHso1Joe5U0Qwe2tByXz2c5GpDNoUkCwL
XPwydA3DnTjrwsp6491c/naHdqTGcusB03Ctu35zR7iC8Tv+sJNiOvpQy/qxxBgVW9WhnWlPY21t
HIJt6xzCrD9IE8yyIORrCiElWyloNkkO7/lbrzPDLuftURB8kb8yR3zduLFMw6Gpr37iZJekB0gt
d3ATADUxMy010Cwx8/NcKgK466t+zwaJGFkgcY04Zuk2P9F5dKU3EgC+72ewpjpnEo/v8Rk4EPHB
Jy6pKIL9k5NIwazxcAys+x3DdHqE8h5Dm8I6F8/bX5IOtlukYR7b4KLKPbHtbnoe/axydr8li7u0
OMcq8hwojQbC0qTbYOlWGXpUHBVLle3JsU1zRnkpsylnATt/NbwLl9noH8Wr/QG/D1y+6E/9NR3R
ski7BUVRR4B6lc3LwSwwrd3A0Zs/NWP/++bL2nZezTjvInWlqFUtrNNiIRLkh2rKjHcGz/LObG9t
1gnQ87b5c6An5pN9BcVMKCoCbUVczftVB4dK/4rAekAgb5KCnrgAk1S2GWqJ4KfAWyxdGYo7o3Xg
gMceFQuUWl44QiM0Mjv0aN7BGHcws2CbYOGPIskIdH8FMKMIaWrDJKJKw4oZCkYUyK496ojpj5h5
MsdAVat9+Ii2ChMerpr57yl3Mfkmbw4ujJXOSQH4ZzUd6v34k0MmxAJ/eEDmfNfhJ2eiqpHe1eyo
ujpUOf6r85ezCKJA93dgaYqSIy0YBrDuYqn1qrJIOLV6DAje/v8LSO6kE/AfKOsgKsaRWKyLClvr
U5e4WEbghySy4DWU75MQjl1d/uFNbmFM8ADidBcU9qAZUbMB4nJ6sDWTnU7XOQFY0UGX9thxIzQT
hClANl50MrVNYhsKQoKcHYC+SR+MBFGreGPn7JEbzlp/rwAouzPHtcrZCweLqqT7+DifJHuC2lZ5
hfaZmbKzxJLStekGCYisGB0eeH9s4B0m2ba4TAxzH16CtF/9lJt49WzGQ6XvfZp/vCzZAvVwIZI+
xXP4Or9kYszCiL5XPIBnR8qSsI0NGkqQblWndaABzbZFGUiR4hG2f4yh4bd82mYNdzjSgGM4WjsV
Cxh2kcP840Z1+4pjscPFgK9NSKPtzMtEIvb2PXuLVNqDu9//b5+Q6IJIAfMWVW1MeCwU12o+oiCe
0aMFmZJECQCbhzRoSh4Bk38AOdUttlltmi2mGhGZ+MHYonZvKRBfDXSWTfQxnNcotvO6PVGzNAj8
InoEm9F+iGIQ9Iw+7gPeel92xtZgpvwDdrGYGXjrWJVi9vYw1ZADUp36iDe5Pj0Y+1/8D6u0Q3qG
ztV1IUjcfJLXrucOIjuG1xgXC9qpxaV+CEeQCUntCON8+eoxltOdkxrJ0Wm69pihvT5Artzyjqhg
XuhM1WZi2SSZ4LNaT3lAEfqHWNgrVCN7EF2IyWFo1VIkV5bRa05fIQZD+iJgn3UTVmKUYajqZhl7
llrnMV/lmR4DJH5uO2SIrCMyUIhzLRU/n1nerjSPpbgO7q1zdyxwD39SEjzdCpt+WsdhTkWTGC+i
2o6DZ6xDPCJMIDFw3yvLksAzb4kR1yslsD99/4eKFmbQmuG6mOHR14ZJuqTBy1b9N5nXN0KfJh/c
KpQNUTNtwFOyh1Ew5qRGm1HRgyB9LsOYZXYRAIfZgk06LvYvQPEZB+Qu58C3zPysB6Qi6xNsIppT
OApaUY/AgII8ZbYGZwH7mTip4WwHNcWIxdztvwz/ZP/yh4oop86D7XDD+Bmqxq559ku/S+/yYIof
ESuy8MYobnyoIseqmQ7H5i4IPVC1ooQC0OzpkD9ZakzBS4LDDnKEbj4fIfX7t1GuyxxOBXTI/rAW
tcgXA2fAm+U0Xy2gGKWgij221A9CkjOeicF3o4+UZOt3UGs01ac76y+nHy8tWzt5eQVV+gM8ocOU
8cmFcHQwDjmcjpLCfr49M73y/027RW1pNj2JUzgQDbwzM/BEukVoAoUL8Gfj/RwX9hS8d0BicP0W
Arv1MYmV4fAZaSqY/3YyC1IfY64Ul/xw3Uq9af6m5cW8NXFhgSFDFksZ1o98ffXbbZeoS0+uS+kJ
Us68IqhrwCPd2FfLAhHVFa46WqrDuaOvRKyiqot6NXhVm+E2ydWQKGQfe9lFLz1CxOuuGd/K03GI
c7DlG2vE+fA9BwEj1kLKGuZyfiSg8tOwObAuMZyVGJn6AHKjILz9BAliS1TS7mG+6048zLgh2pd3
41mA5YIiin4K4s28vE6TV4akOFP7K/he6+wXLoBkJAavSULwH3giChwgkwxdoKG2GuwR6g8nOvjf
+2IRQUJmr7OZcndvEbr0xPCjLCIwvyQpTNzUcI3QK6m1WbpD7ITu+nkhdEPktgDFWqAVOVI2/QOY
or1U2RcltGm9BOo373K9g6bjmddI+P/NgFH9tvMjQCqcRwFb/zqO3dF7p9zKNN87F0i5RcBhzSSG
QNZxVJRi3lbdJMC72M0OlvKa3JUNmmdoau2ZfEe6nGMGsJu7U7apHjx5Fk5JrJF3cf3oLKIc/B5o
WTorJLQ6D2YwUEDJtlsnZ43ZwLjndwNphguDjfNR3+jbr4Mnahe1ttY6wrrZahNnvr5f4EWkiKYH
LVn9qt7qQ4i6CgLDcbs6uSrpvgPN5JKzRQnnplX6m46NjCUcNvIL2mAAnaiBH8RCuYuhzSMlAYAh
gcvNNkkBgsb9NIx6N7E267oBkBixydfv9NkVJ+Qh7wSHu5Vjz9mtjXLa/gbXK1LZU47gw6NPbqSP
Pqx62X9DywxEvu5/dkT0y4f4lNMdhmBpOHpvdU18Myf4UmUeri3UECpEwMWcPaIe8n2XdGSFN2t5
3W0TPT8KaQAR42JY67ilj4cItnMkkCg1uVtFLmU/K9Ul/8Zbr/hlVGVT0GY5Jc8KbM+NIN3p/Z1U
14Vve8u8RsDD0ZRqmO/AIrkHmU6lEWH+mqqAdKvw+eU5/KqfBqZHdmEP/XGwRft68BOApeFvoQnu
CBfUUKH5f5OYGyMZmO+WeKTPpxIcIB7imBJIpIzxITmwBhZOdqEypNSXdvyTxA/bQmIfrpm/IIIM
CxakWBqGNlhfa+Wv6Lg2q7P7+XiCgdnqw537YkMfIz6fLrz6GmScoWfb42EJ1HeuJMx9HYr+FxLW
KkAkscInI9P+2RNQcFXcHHef02zN+OK4RikQN9QfbjjoTP0zdgKbjW5l0CQGFq0vwk4avxvs9o8V
bdu9qBjyPN7IjBJ0iRWmMhsIEJ0pUAUevm1PdAxZwLGH7tlUnhkeKMCQke66NRe6wc7jz2l3RgmT
UzB/zioRVOn9SUEp435feuRi9+NXW4JhEjELihtJv3lxusVUxT5e20LKzarAlZrQIQ8JrIAbnLu+
eEqmIeIZG5qlhUTfDmaBXLM9X3qQClAPxK9MNBxT+zjpYfHR+hHyJ/OOlTx5anN0w0oMEKD/W5DP
BUyez8KVzad4EkwA8mEs8douF7CM/lW2K95AjYsQhFN/FhxWSmShBjrDgEd4TvV/SoeFcb2RHEj2
9LlEzTfCxh4/oVySx6PKC8lQ+T3/0fvdK1UjWmrzvarpvGHHTRaGLuJJL/SlgBrwXM3BG4Td3rFH
+z5EcSPp/hJNFnENfFZcPGYDv1ENIxnKkkRO/Eb5MkqHq6RQ2OKu5CnBchg7/FvaJi9bLowiCVfI
PRy1A43S9qkV7a2mEJ3LFf13Ag4MLy/GbeG/lLmjfwXRCbLGyPqDYE0wLrdIXrL60tbSvIwtcXeR
7BxO5HBUD7Zsrh0Da0zObjRm8wzIzYBESdAipoYuw4DWqzaacqrdwsRMvIxxsPx/uphMRVE5+som
uz8VX7oYYeR9ZTtjq8JhYL0FIxbHnOX8QUqsMI+dMhpA1jTJvdFcEI03chjIaUZbS0EEPMn+e+is
KLSHYMUiMIVFIg0mPdDTCKZZM0gTmOs1uVFgrLYIAM3BUsjPETNODfaXAkCSOHZ1UVSmutpMmaWU
Gf6dPsvzOjTnnQxM5b+wLStPxEaVoq5EZlRuuhh3nfI7UudHK9DrR4kLga0IIZfTkpQv1L2UaN8p
sbeuPgznZHT6cVuG3W/Z+rlaQfb0WJqao9GLaSKGfcDSrpEMj+tkWZhJurpwRgz/gt/PwytjfWJP
I20eVLjBwS3FX4PJVRk1zxhoW76UEst2l3Yh0KBpCXJU82qISFN/T8vS5KExTTXmR2eoAaEDlHGE
0pHbsWIU8V2BQn9bMmTLpkSqqyKDPSlybmLJZcdn7taxi38qTe+ToDRiN/ALPX5wbcLWdzOpYnQG
aR5wVpiAwV9jo0oD0im1Q50waN/zqWbLHbCpdFvVNGRq6jAyr5E2zUAS/WWlgaFo41vd7X/GSVZ8
aiHP2FBdtputVAGe6yqZXalslm+HkIPpL7swhcVXplRbB1BwtPMdUbDPl4pcBv0nhxpnHDceSUQ3
zD/3Ws/PNWtG9/d1LbNmCn2wBLR7rqSTGuDi6ZsetXhX4FUP2PufHttZy9wnAi/KeNUJ4i3Q762V
9D+j3kTugfGLDo0R/Tm2NTijsWpps4f9WCRWfxryrd4Fm2y/QWsEs+1COCOkG+4vPo8GpG3aeJIO
A9kQx1Yk1GM0V0fja/35PuXs0t52aqQCp6SCjUiooXvUzVJPVOBg7isoY8iJltLDK/5CuYadPZZM
PCpvTAUo9rRO0CL8H93Psk9pCKMMMvhTEB4GzCIYgQAltjlTIDZBXXcvGaUtrOubfAELMjluOPQI
yKEVInSGVnape0Fk23EPxfPEW8bgikJfyxJ5w7b4mGufrBjrPcSxPlomM2FfI+dRY8tWUGK6zJoW
qv+QSxCui9qNAmAxFKVPc9WbgR3TGcVQCVraS8SmPV5ffBdW9Q+jvKzq4zW7AA2CMyP8dzWJqukO
8KyUIr33kgpTV04OyBaCZ+lBYQ5jds6U34WsBRFThg7Wye/UU33i25ol2kG7gSAwCAn92KX7rzK8
h7AmJVKXmnTM+h9OW+CxvKihWJRh+z290wRZYf9va8hXjgUEcxrr46PqQsh5sFIyTL3Vf8JvTc7c
g7qrXeBSjHZqA8xRtjVDG+TV/d3l4/JLJ3JwXvK1SiujChlrmVHXQ/6sW0ajFbil2idedyy+m8CU
n1+baqphz1vyp3zCn70T2aOwOH11uF9KulXPtRVnOXkuUgxRfo8kqoVbiKOhvpY3bp3W5bjg8/6P
7PAP18+BGIzUkBTLBDEHHNUr6yIuqmOthheXV0fmQvVrluKsKXyIG8CkiYUSuadLR1FGZ9QGkrxk
MMQCBwvY1hBHcUTbVKaz7FQ3KroO5aUPt5Mcml8d3VD+eIDoJkSc4upbOp65J5ws+0okhitew/of
3RvcQwMxDHddG5YRLrOKSA/v+ZrJmAypuTQoHWt2vvxE8KWfMrC6E7Z2bQmeH+pnEYeWSMF7x7d/
4UUxOsU6qqcVvDaUFbliBGVZx2oBFlq5Brcqf+VOfPtRHpG318bLpXHiFcQap6BfEOM6HBetK2mb
PfcQj8ISSMbbSFbXRHD1J2FQpujzoyD+9WIdZ2V/beJiWfhdD9MjcnxYSvnyNw1EWvAN1gfjzocV
7a4aj3lyoc/eoOJGj7oXBrRoj1LKXxHlF07yqg2V6UHo3gFePeyB1k5/U35U3aet8IqwXKRl5Zx9
Xt1GMR6R+ZBsibLhceHuebOpDWiWFAx0soSG/FYAU6z5VvliWydhfm/GfE1rva68Dcn3j7X5
`protect end_protected
